module aes_aes_die_0 ( clk, key, ld, rst, text_in, done, text_out, sa00_sr_0, sa00_sr_1, 
       sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, 
       sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, 
       sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, 
       sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, 
       sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, 
       sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, 
       sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa20_sr_0, 
       sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_0, sa21_sr_1, 
       sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, 
       sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, 
       sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, 
       sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, 
       sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, 
       sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, 
       u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_16, 
       u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_3, 
       u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa01_0, 
        sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, sa02_1, 
        sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, sa03_2, 
        sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, sa10_3, 
        sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, 
        sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, 
        sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, 
        sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, 
        sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa22_0, 
        sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa23_0, sa23_1, 
        sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
        sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, sa31_3, 
        sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, 
        sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, sa33_5, 
        sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_0, w3_1, w3_10, 
        w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, 
        w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9 );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;
  input sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_sr_0, 
        sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, sa02_sr_1, 
        sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, 
        sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, 
        sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, 
        sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, 
        sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, 
        sa13_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, 
        sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa22_sr_0, 
        sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, 
        sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, 
        sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, 
        sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, 
        sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, 
        sa33_sr_6, sa33_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, 
        u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, u0_subword_21, u0_subword_22, 
        u0_subword_23, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9;
  output sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa01_0, 
        sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, sa02_1, 
        sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, sa03_2, 
        sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, sa10_3, 
        sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, 
        sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, 
        sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, 
        sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, sa20_7, 
        sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa22_0, 
        sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa23_0, sa23_1, 
        sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
        sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, sa31_2, sa31_3, 
        sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, 
        sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, sa33_5, 
        sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_0, w3_1, w3_10, 
        w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, 
        w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9;
  wire N100, N101, N102, N103, N104, N105, N114, N115, N116, 
       N117, N118, N119, N120, N121, N130, N131, N132, N133, 
       N134, N135, N136, N137, N146, N147, N148, N149, N150, 
       N151, N152, N153, N162, N163, N164, N165, N166, N167, 
       N168, N169, N178, N179, N180, N181, N182, N183, N184, 
       N185, N194, N195, N196, N197, N198, N199, N200, N201, 
       N210, N211, N212, N213, N214, N215, N216, N217, N226, 
       N227, N228, N229, N23, N230, N231, N232, N233, N242, 
       N243, N244, N245, N246, N247, N248, N249, N258, N259, 
       N260, N261, N262, N263, N264, N265, N274, N275, N276, 
       N277, N278, N279, N280, N281, N34, N35, N36, N37, 
       N378, N379, N38, N380, N381, N382, N383, N384, N385, 
       N386, N387, N388, N389, N39, N390, N391, N392, N393, 
       N394, N395, N396, N397, N398, N399, N40, N400, N401, 
       N402, N403, N404, N405, N406, N407, N408, N409, N41, 
       N410, N411, N412, N413, N414, N415, N416, N417, N418, 
       N419, N420, N421, N422, N423, N424, N425, N426, N427, 
       N428, N429, N430, N431, N432, N433, N434, N435, N436, 
       N437, N438, N439, N440, N441, N442, N443, N444, N445, 
       N446, N447, N448, N449, N450, N451, N452, N453, N454, 
       N455, N456, N457, N458, N459, N460, N461, N462, N463, 
       N464, N465, N466, N467, N468, N469, N470, N471, N472, 
       N473, N474, N475, N476, N477, N478, N479, N480, N481, 
       N482, N483, N484, N485, N486, N487, N488, N489, N490, 
       N491, N492, N493, N494, N495, N496, N497, N498, N499, 
       N50, N500, N501, N502, N503, N504, N505, N51, N52, 
       N53, N54, N55, N56, N57, N66, N67, N68, N69, 
       N70, N71, N72, N73, N82, N83, N84, N85, N86, 
       N87, N88, N89, N98, N99, n1, n10, n100, n1000, 
       n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
       n101, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
       n1018, n1019, n102, n1020, n1021, n1022, n1023, n1024, n1025, 
       n1026, n1027, n1028, n1029, n103, n1030, n1031, n1032, n1033, 
       n1034, n1035, n1036, n1037, n1038, n1039, n104, n1040, n1041, 
       n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n105, 
       n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
       n1059, n106, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
       n1067, n1068, n1069, n107, n1070, n1071, n1072, n1073, n1074, 
       n1075, n1076, n1077, n1078, n1079, n108, n1080, n1081, n1082, 
       n1083, n1084, n1085, n1086, n1087, n1088, n1089, n109, n1090, 
       n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
       n11, n110, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
       n1107, n1108, n1109, n111, n1110, n1111, n1112, n1113, n1114, 
       n1115, n1116, n1117, n1118, n1119, n112, n1120, n1121, n1122, 
       n1123, n1124, n1125, n1126, n1127, n1128, n1129, n113, n1130, 
       n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
       n114, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
       n1148, n1149, n115, n1150, n1151, n1152, n1153, n1154, n1155, 
       n1156, n1157, n1158, n1159, n116, n1160, n1161, n1162, n1163, 
       n1164, n1165, n1166, n1167, n1168, n1169, n117, n1170, n1171, 
       n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n118, 
       n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
       n1189, n119, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
       n1197, n1198, n1199, n12, n120, n1200, n1201, n1202, n1203, 
       n1204, n1205, n1206, n1207, n1208, n1209, n121, n1210, n1211, 
       n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n122, 
       n1220, n1221, n1222, n123, n124, n125, n126, n127, n128, 
       n129, n13, n130, n131, n132, n133, n134, n135, n136, 
       n137, n138, n139, n14, n140, n141, n142, n143, n144, 
       n145, n146, n147, n148, n149, n15, n150, n151, n152, 
       n153, n154, n155, n156, n157, n158, n159, n16, n160, 
       n161, n162, n163, n164, n165, n166, n167, n168, n169, 
       n17, n170, n171, n172, n173, n174, n175, n176, n177, 
       n178, n179, n18, n180, n181, n182, n183, n184, n185, 
       n186, n187, n188, n189, n19, n190, n191, n192, n193, 
       n194, n195, n196, n197, n198, n199, n2, n20, n200, 
       n201, n202, n203, n204, n205, n206, n207, n208, n209, 
       n21, n210, n211, n212, n213, n214, n215, n216, n217, 
       n218, n219, n22, n220, n221, n222, n223, n224, n225, 
       n226, n227, n228, n229, n23, n230, n231, n232, n233, 
       n234, n235, n236, n237, n238, n239, n24, n240, n241, 
       n242, n243, n244, n245, n246, n247, n248, n249, n25, 
       n250, n251, n252, n253, n254, n255, n256, n258, n259, 
       n26, n260, n261, n262, n263, n264, n265, n266, n267, 
       n268, n269, n27, n270, n271, n272, n275, n276, n277, 
       n278, n279, n28, n280, n281, n283, n284, n285, n286, 
       n288, n289, n29, n290, n291, n292, n294, n295, n296, 
       n297, n298, n3, n30, n300, n301, n302, n303, n304, 
       n305, n306, n307, n308, n309, n31, n310, n311, n312, 
       n314, n315, n316, n317, n318, n319, n32, n321, n322, 
       n323, n324, n325, n327, n328, n329, n33, n330, n331, 
       n332, n334, n335, n336, n337, n338, n339, n34, n341, 
       n342, n343, n345, n347, n348, n349, n35, n350, n351, 
       n352, n353, n354, n355, n356, n357, n358, n359, n36, 
       n360, n361, n362, n363, n365, n366, n367, n368, n369, 
       n37, n370, n372, n373, n374, n375, n376, n378, n379, 
       n38, n380, n381, n382, n384, n385, n386, n387, n388, 
       n39, n390, n391, n392, n394, n395, n396, n398, n399, 
       n4, n40, n400, n401, n402, n403, n404, n405, n407, 
       n408, n409, n41, n410, n412, n413, n414, n416, n417, 
       n418, n419, n42, n421, n422, n423, n424, n425, n426, 
       n427, n428, n429, n43, n431, n432, n433, n434, n436, 
       n437, n438, n439, n44, n440, n441, n442, n443, n444, 
       n445, n446, n448, n449, n45, n450, n451, n452, n453, 
       n454, n455, n456, n457, n459, n46, n460, n461, n462, 
       n464, n465, n466, n468, n469, n47, n470, n471, n472, 
       n473, n475, n476, n477, n478, n479, n48, n481, n482, 
       n483, n484, n485, n486, n487, n488, n489, n49, n490, 
       n491, n492, n493, n495, n496, n497, n498, n499, n5, 
       n50, n500, n502, n503, n504, n505, n506, n508, n509, 
       n51, n510, n511, n512, n513, n515, n516, n517, n518, 
       n519, n52, n520, n521, n522, n523, n524, n526, n528, 
       n529, n53, n530, n531, n532, n533, n534, n535, n536, 
       n537, n538, n539, n54, n540, n541, n542, n543, n544, 
       n546, n547, n548, n55, n550, n551, n552, n554, n555, 
       n556, n557, n558, n56, n560, n561, n562, n564, n565, 
       n566, n568, n569, n57, n570, n571, n572, n573, n574, 
       n575, n576, n577, n578, n579, n58, n581, n582, n583, 
       n584, n586, n587, n588, n59, n590, n591, n592, n593, 
       n595, n596, n597, n598, n599, n6, n60, n600, n601, 
       n602, n603, n605, n606, n607, n608, n609, n61, n610, 
       n611, n612, n613, n614, n615, n616, n617, n618, n619, 
       n62, n620, n622, n623, n624, n625, n626, n628, n629, 
       n63, n630, n632, n633, n634, n635, n636, n638, n639, 
       n64, n640, n642, n643, n644, n645, n646, n647, n649, 
       n65, n650, n651, n652, n653, n655, n656, n657, n658, 
       n659, n66, n660, n661, n662, n663, n664, n665, n666, 
       n667, n669, n67, n670, n671, n672, n673, n674, n676, 
       n677, n678, n679, n68, n680, n682, n683, n684, n685, 
       n686, n687, n689, n69, n690, n691, n692, n693, n694, 
       n696, n697, n698, n7, n70, n700, n702, n703, n704, 
       n705, n706, n707, n708, n709, n71, n710, n711, n712, 
       n713, n714, n715, n716, n718, n719, n72, n720, n721, 
       n722, n724, n725, n726, n728, n729, n73, n730, n731, 
       n732, n734, n735, n736, n738, n739, n74, n740, n742, 
       n743, n744, n745, n746, n747, n748, n749, n75, n750, 
       n751, n752, n753, n755, n756, n757, n758, n76, n760, 
       n761, n762, n764, n765, n766, n767, n769, n77, n770, 
       n771, n772, n773, n774, n775, n776, n777, n778, n779, 
       n78, n780, n781, n782, n783, n784, n785, n786, n787, 
       n788, n789, n79, n790, n791, n792, n793, n794, n796, 
       n797, n798, n799, n8, n80, n800, n801, n802, n803, 
       n804, n806, n807, n808, n809, n81, n810, n812, n813, 
       n814, n816, n817, n818, n819, n82, n820, n821, n823, 
       n824, n825, n826, n827, n828, n829, n83, n830, n831, 
       n832, n833, n834, n835, n836, n837, n838, n839, n84, 
       n840, n841, n843, n844, n845, n846, n847, n848, n85, 
       n850, n851, n852, n853, n854, n856, n857, n858, n859, 
       n86, n861, n862, n863, n864, n865, n866, n867, n868, 
       n869, n87, n870, n872, n874, n875, n876, n877, n878, 
       n879, n88, n880, n881, n882, n883, n884, n885, n886, 
       n887, n888, n889, n89, n890, n892, n893, n894, n896, 
       n898, n899, n9, n90, n900, n901, n902, n903, n904, 
       n905, n907, n908, n909, n91, n911, n912, n913, n915, 
       n916, n917, n918, n919, n92, n920, n921, n922, n923, 
       n924, n925, n926, n927, n929, n93, n930, n931, n932, 
       n933, n935, n936, n937, n939, n94, n940, n941, n942, 
       n944, n945, n946, n947, n948, n949, n95, n950, n951, 
       n952, n954, n955, n956, n957, n958, n959, n96, n960, 
       n961, n962, n964, n965, n966, n967, n969, n97, n970, 
       n971, n972, n973, n974, n975, n976, n977, n978, n979, 
       n98, n980, n981, n982, n983, n984, n985, n986, n987, 
       n988, n989, n99, n990, n991, n992, n993, n994, n995, 
       n996, n997, n998, n999, u0_N108, u0_N109, u0_N110, u0_N111, u0_N112, 
       u0_N113, u0_N114, u0_N115, u0_N116, u0_N117, u0_N118, u0_N119, u0_N120, u0_N121, 
       u0_N122, u0_N123, u0_N124, u0_N125, u0_N126, u0_N127, u0_N128, u0_N129, u0_N130, 
       u0_N131, u0_N132, u0_N133, u0_N134, u0_N135, u0_N136, u0_N137, u0_N138, u0_N139, 
       u0_N174, u0_N175, u0_N176, u0_N177, u0_N178, u0_N179, u0_N180, u0_N181, u0_N182, 
       u0_N183, u0_N184, u0_N185, u0_N186, u0_N187, u0_N188, u0_N189, u0_N190, u0_N191, 
       u0_N192, u0_N193, u0_N194, u0_N195, u0_N196, u0_N197, u0_N198, u0_N199, u0_N200, 
       u0_N201, u0_N202, u0_N203, u0_N204, u0_N205, u0_N240, u0_N241, u0_N242, u0_N243, 
       u0_N244, u0_N245, u0_N246, u0_N247, u0_N248, u0_N249, u0_N250, u0_N251, u0_N252, 
       u0_N253, u0_N254, u0_N255, u0_N256, u0_N257, u0_N258, u0_N259, u0_N260, u0_N261, 
       u0_N262, u0_N263, u0_N264, u0_N265, u0_N266, u0_N267, u0_N268, u0_N269, u0_N270, 
       u0_N271, u0_N42, u0_N43, u0_N44, u0_N45, u0_N46, u0_N47, u0_N48, u0_N49, 
       u0_N50, u0_N51, u0_N52, u0_N53, u0_N54, u0_N55, u0_N56, u0_N57, u0_N58, 
       u0_N59, u0_N60, u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, u0_N66, u0_N67, 
       u0_N68, u0_N69, u0_N70, u0_N71, u0_N72, u0_N73, u0_n1, u0_n10, u0_n100, 
       u0_n101, u0_n102, u0_n103, u0_n104, u0_n105, u0_n106, u0_n107, u0_n108, u0_n109, 
       u0_n11, u0_n110, u0_n111, u0_n112, u0_n113, u0_n114, u0_n115, u0_n116, u0_n117, 
       u0_n118, u0_n119, u0_n12, u0_n120, u0_n121, u0_n122, u0_n123, u0_n124, u0_n125, 
       u0_n126, u0_n127, u0_n128, u0_n129, u0_n13, u0_n130, u0_n131, u0_n132, u0_n133, 
       u0_n134, u0_n135, u0_n136, u0_n137, u0_n138, u0_n139, u0_n14, u0_n140, u0_n141, 
       u0_n142, u0_n143, u0_n144, u0_n145, u0_n146, u0_n147, u0_n148, u0_n149, u0_n15, 
       u0_n150, u0_n151, u0_n152, u0_n153, u0_n154, u0_n155, u0_n156, u0_n157, u0_n158, 
       u0_n159, u0_n16, u0_n160, u0_n161, u0_n162, u0_n163, u0_n164, u0_n165, u0_n166, 
       u0_n167, u0_n168, u0_n169, u0_n17, u0_n170, u0_n171, u0_n172, u0_n173, u0_n174, 
       u0_n175, u0_n176, u0_n177, u0_n178, u0_n179, u0_n18, u0_n180, u0_n181, u0_n182, 
       u0_n183, u0_n184, u0_n185, u0_n186, u0_n187, u0_n188, u0_n189, u0_n19, u0_n190, 
       u0_n191, u0_n192, u0_n193, u0_n194, u0_n195, u0_n196, u0_n197, u0_n198, u0_n199, 
       u0_n2, u0_n20, u0_n200, u0_n201, u0_n202, u0_n203, u0_n204, u0_n205, u0_n206, 
       u0_n207, u0_n208, u0_n209, u0_n21, u0_n210, u0_n211, u0_n212, u0_n213, u0_n214, 
       u0_n215, u0_n216, u0_n217, u0_n218, u0_n219, u0_n22, u0_n220, u0_n221, u0_n222, 
       u0_n223, u0_n224, u0_n225, u0_n226, u0_n227, u0_n228, u0_n229, u0_n23, u0_n230, 
       u0_n231, u0_n232, u0_n233, u0_n234, u0_n235, u0_n236, u0_n237, u0_n238, u0_n239, 
       u0_n24, u0_n240, u0_n241, u0_n242, u0_n243, u0_n244, u0_n245, u0_n246, u0_n247, 
       u0_n248, u0_n249, u0_n25, u0_n250, u0_n251, u0_n253, u0_n254, u0_n255, u0_n257, 
       u0_n258, u0_n259, u0_n26, u0_n261, u0_n262, u0_n263, u0_n264, u0_n265, u0_n267, 
       u0_n269, u0_n27, u0_n271, u0_n273, u0_n275, u0_n277, u0_n279, u0_n28, u0_n281, 
       u0_n283, u0_n285, u0_n287, u0_n29, u0_n3, u0_n30, u0_n31, u0_n32, u0_n33, 
       u0_n34, u0_n35, u0_n36, u0_n37, u0_n38, u0_n39, u0_n4, u0_n40, u0_n41, 
       u0_n42, u0_n43, u0_n44, u0_n45, u0_n46, u0_n47, u0_n48, u0_n49, u0_n5, 
       u0_n50, u0_n51, u0_n52, u0_n53, u0_n54, u0_n55, u0_n56, u0_n57, u0_n58, 
       u0_n59, u0_n6, u0_n60, u0_n61, u0_n62, u0_n63, u0_n64, u0_n65, u0_n66, 
       u0_n67, u0_n68, u0_n69, u0_n7, u0_n70, u0_n71, u0_n72, u0_n73, u0_n74, 
       u0_n75, u0_n76, u0_n77, u0_n78, u0_n79, u0_n8, u0_n80, u0_n81, u0_n82, 
       u0_n83, u0_n84, u0_n85, u0_n86, u0_n87, u0_n88, u0_n89, u0_n9, u0_n90, 
       u0_n91, u0_n92, u0_n93, u0_n94, u0_n95, u0_n96, u0_n97, u0_n98, u0_n99, 
       u0_r0_N70, u0_r0_N71, u0_r0_N72, u0_r0_N73, u0_r0_N74, u0_r0_N75, u0_r0_N76, u0_r0_N77, u0_r0_N78, 
       u0_r0_N79, u0_r0_N80, u0_r0_N81, u0_r0_n1, u0_r0_n10, u0_r0_n11, u0_r0_n12, u0_r0_n13, u0_r0_n14, 
       u0_r0_n15, u0_r0_n16, u0_r0_n17, u0_r0_n18, u0_r0_n19, u0_r0_n2, u0_r0_n20, u0_r0_n21, u0_r0_n22, 
       u0_r0_n23, u0_r0_n24, u0_r0_n25, u0_r0_n3, u0_r0_n4, u0_r0_n5, u0_r0_n6, u0_r0_n7, u0_r0_n8, 
       u0_r0_n9, u0_r0_rcnt_0, u0_r0_rcnt_1, u0_r0_rcnt_2, u0_rcon_24, u0_rcon_25, u0_rcon_26, u0_rcon_27, u0_rcon_28, 
       u0_rcon_29, u0_rcon_30, u0_rcon_31, u0_subword_24, u0_subword_25, u0_subword_26, u0_subword_27, u0_subword_28, u0_subword_29, 
       u0_subword_30, u0_subword_31, u0_u0_n1, u0_u0_n171, u0_u0_n22, u0_u0_n438, u0_u0_n439, u0_u0_n440, u0_u0_n441, 
       u0_u0_n442, u0_u0_n443, u0_u0_n444, u0_u0_n445, u0_u0_n446, u0_u0_n447, u0_u0_n448, u0_u0_n449, u0_u0_n450, 
       u0_u0_n451, u0_u0_n452, u0_u0_n453, u0_u0_n454, u0_u0_n455, u0_u0_n456, u0_u0_n457, u0_u0_n458, u0_u0_n459, 
       u0_u0_n460, u0_u0_n461, u0_u0_n462, u0_u0_n463, u0_u0_n464, u0_u0_n465, u0_u0_n466, u0_u0_n467, u0_u0_n468, 
       u0_u0_n469, u0_u0_n470, u0_u0_n471, u0_u0_n472, u0_u0_n473, u0_u0_n474, u0_u0_n475, u0_u0_n476, u0_u0_n477, 
       u0_u0_n478, u0_u0_n479, u0_u0_n480, u0_u0_n481, u0_u0_n482, u0_u0_n483, u0_u0_n484, u0_u0_n485, u0_u0_n486, 
       u0_u0_n487, u0_u0_n488, u0_u0_n489, u0_u0_n490, u0_u0_n491, u0_u0_n492, u0_u0_n493, u0_u0_n494, u0_u0_n495, 
       u0_u0_n496, u0_u0_n497, u0_u0_n498, u0_u0_n499, u0_u0_n500, u0_u0_n501, u0_u0_n502, u0_u0_n503, u0_u0_n504, 
       u0_u0_n505, u0_u0_n506, u0_u0_n507, u0_u0_n508, u0_u0_n509, u0_u0_n510, u0_u0_n511, u0_u0_n512, u0_u0_n513, 
       u0_u0_n514, u0_u0_n515, u0_u0_n516, u0_u0_n517, u0_u0_n518, u0_u0_n519, u0_u0_n520, u0_u0_n521, u0_u0_n522, 
       u0_u0_n523, u0_u0_n524, u0_u0_n525, u0_u0_n526, u0_u0_n527, u0_u0_n528, u0_u0_n529, u0_u0_n530, u0_u0_n531, 
       u0_u0_n532, u0_u0_n533, u0_u0_n534, u0_u0_n535, u0_u0_n536, u0_u0_n537, u0_u0_n538, u0_u0_n539, u0_u0_n540, 
       u0_u0_n541, u0_u0_n542, u0_u0_n543, u0_u0_n544, u0_u0_n545, u0_u0_n546, u0_u0_n547, u0_u0_n548, u0_u0_n549, 
       u0_u0_n550, u0_u0_n551, u0_u0_n552, u0_u0_n553, u0_u0_n554, u0_u0_n555, u0_u0_n556, u0_u0_n557, u0_u0_n558, 
       u0_u0_n559, u0_u0_n560, u0_u0_n561, u0_u0_n562, u0_u0_n563, u0_u0_n564, u0_u0_n565, u0_u0_n566, u0_u0_n567, 
       u0_u0_n568, u0_u0_n569, u0_u0_n570, u0_u0_n571, u0_u0_n572, u0_u0_n573, u0_u0_n574, u0_u0_n575, u0_u0_n576, 
       u0_u0_n577, u0_u0_n578, u0_u0_n579, u0_u0_n580, u0_u0_n581, u0_u0_n582, u0_u0_n583, u0_u0_n584, u0_u0_n585, 
       u0_u0_n586, u0_u0_n587, u0_u0_n588, u0_u0_n589, u0_u0_n590, u0_u0_n591, u0_u0_n592, u0_u0_n593, u0_u0_n594, 
       u0_u0_n595, u0_u0_n596, u0_u0_n597, u0_u0_n598, u0_u0_n599, u0_u0_n600, u0_u0_n601, u0_u0_n602, u0_u0_n603, 
       u0_u0_n604, u0_u0_n605, u0_u0_n606, u0_u0_n607, u0_u0_n608, u0_u0_n609, u0_u0_n610, u0_u0_n611, u0_u0_n612, 
       u0_u0_n613, u0_u0_n614, u0_u0_n615, u0_u0_n616, u0_u0_n617, u0_u0_n618, u0_u0_n619, u0_u0_n620, u0_u0_n621, 
       u0_u0_n622, u0_u0_n623, u0_u0_n624, u0_u0_n625, u0_u0_n626, u0_u0_n627, u0_u0_n628, u0_u0_n629, u0_u0_n630, 
       u0_u0_n631, u0_u0_n632, u0_u0_n633, u0_u0_n634, u0_u0_n635, u0_u0_n636, u0_u0_n637, u0_u0_n638, u0_u0_n639, 
       u0_u0_n640, u0_u0_n641, u0_u0_n642, u0_u0_n643, u0_u0_n644, u0_u0_n645, u0_u0_n646, u0_u0_n647, u0_u0_n648, 
       u0_u0_n649, u0_u0_n650, u0_u0_n651, u0_u0_n652, u0_u0_n653, u0_u0_n654, u0_u0_n655, u0_u0_n656, u0_u0_n657, 
       u0_u0_n658, u0_u0_n659, u0_u0_n660, u0_u0_n661, u0_u0_n662, u0_u0_n663, u0_u0_n664, u0_u0_n665, u0_u0_n666, 
       u0_u0_n667, u0_u0_n668, u0_u0_n669, u0_u0_n670, u0_u0_n671, u0_u0_n672, u0_u0_n673, u0_u0_n674, u0_u0_n675, 
       u0_u0_n676, u0_u0_n677, u0_u0_n678, u0_u0_n679, u0_u0_n680, u0_u0_n681, u0_u0_n682, u0_u0_n683, u0_u0_n684, 
       u0_u0_n685, u0_u0_n686, u0_u0_n687, u0_u0_n688, u0_u0_n689, u0_u0_n690, u0_u0_n691, u0_u0_n692, u0_u0_n693, 
       u0_u0_n694, u0_u0_n695, u0_u0_n696, u0_u0_n697, u0_u0_n698, u0_u0_n699, u0_u0_n700, u0_u0_n701, u0_u0_n702, 
       u0_u0_n703, u0_u0_n704, u0_u0_n705, u0_u0_n706, u0_u0_n707, u0_u0_n708, u0_u0_n709, u0_u0_n710, u0_u0_n711, 
       u0_u0_n712, u0_u0_n713, u0_u0_n714, u0_u0_n715, u0_u0_n716, u0_u0_n717, u0_u0_n718, u0_u0_n719, u0_u0_n720, 
       u0_u0_n721, u0_u0_n722, u0_u0_n723, u0_u0_n724, u0_u0_n725, u0_u0_n726, u0_u0_n727, u0_u0_n728, u0_u0_n729, 
       u0_u0_n730, u0_u0_n731, u0_u0_n732, u0_u0_n733, u0_u0_n734, u0_u0_n735, u0_u0_n736, u0_u0_n737, u0_u0_n738, 
       u0_u0_n739, u0_u0_n740, u0_u0_n741, u0_u0_n742, u0_u0_n743, u0_u0_n744, u0_u0_n745, u0_u0_n746, u0_u0_n747, 
       u0_u0_n748, u0_u0_n749, u0_u0_n750, u0_u0_n751, u0_u0_n752, u0_u0_n753, u0_u0_n754, u0_u0_n755, u0_u0_n756, 
       u0_u0_n757, u0_u0_n758, u0_u0_n759, u0_u0_n760, u0_u0_n761, u0_u0_n762, u0_u0_n763, u0_u0_n764, u0_u0_n765, 
       u0_u0_n766, u0_u0_n767, u0_u0_n768, u0_u0_n769, u0_u0_n770, u0_u0_n771, u0_u0_n772, u0_u0_n773, u0_u0_n774, 
       u0_u0_n775, u0_u0_n776, u0_u0_n777, u0_u0_n778, u0_u0_n779, u0_u0_n780, u0_u0_n781, u0_u0_n782, u0_u0_n783, 
       u0_u0_n784, u0_u0_n785, u0_u0_n786, u0_u0_n787, u0_u0_n788, u0_u0_n789, u0_u0_n790, u0_u0_n791, u0_u0_n792, 
       u0_u0_n793, u0_u0_n794, u0_u0_n795, u0_u0_n796, u0_u0_n797, u0_u0_n798, u0_u0_n799, u0_u0_n800, u0_u0_n801, 
       u0_u0_n802, u0_u0_n803, u0_u0_n804, u0_u0_n805, u0_u0_n806, u0_u0_n807, u0_u0_n808, u0_u0_n809, u0_u0_n810, 
       u0_u0_n811, u0_u0_n812, u0_u0_n813, u0_u0_n814, u0_u0_n815, u0_u0_n816, u0_u0_n817, u0_u0_n818, u0_u0_n819, 
       u0_u0_n820, u0_u0_n821, u0_u0_n822, u0_u0_n823, u0_u0_n824, u0_u0_n825, u0_u0_n826, u0_u0_n827, u0_u0_n828, 
       u0_u0_n829, u0_u0_n830, u0_u0_n831, u0_u0_n832, u0_u0_n833, u0_u0_n834, u0_u0_n835, u0_u0_n836, u0_u0_n837, 
       u0_u0_n838, u0_u0_n839, u0_u0_n840, u0_u0_n841, u0_u0_n842, u0_u0_n843, u0_u0_n844, u0_u0_n845, u0_u0_n846, 
       u0_u0_n847, u0_u0_n848, u0_u0_n849, u0_u0_n850, u0_u0_n851, u0_u0_n852, u0_u0_n853, u0_u0_n854, u0_u0_n855, 
       u0_u0_n856, u0_u0_n857, u0_u0_n858, u0_u0_n859, u0_u0_n860, u0_u0_n861, u0_u0_n862, u0_u0_n863, u0_u0_n864, 
       u0_u0_n865, u0_u0_n866, u0_u0_n867, u0_u0_n868, u0_u0_n869, u0_u0_n870, u0_u0_n871, u0_u0_n872, u0_u0_n873, 
       u0_u0_n874, u0_u0_n875, u0_u0_n876, u0_u0_n877, u0_u0_n878, u0_u0_n879, w0_0, w0_1, w0_10, 
       w0_11, w0_12, w0_13, w0_14, w0_15, w0_16, w0_17, w0_18, w0_19, 
       w0_2, w0_20, w0_21, w0_22, w0_23, w0_24, w0_25, w0_26, w0_27, 
       w0_28, w0_29, w0_3, w0_30, w0_31, w0_4, w0_5, w0_6, w0_7, 
       w0_8, w0_9, w1_0, w1_1, w1_10, w1_11, w1_12, w1_13, w1_14, 
       w1_15, w1_16, w1_17, w1_18, w1_19, w1_2, w1_20, w1_21, w1_22, 
       w1_23, w1_24, w1_25, w1_26, w1_27, w1_28, w1_29, w1_3, w1_30, 
       w1_31, w1_4, w1_5, w1_6, w1_7, w1_8, w1_9, w2_0, w2_1, 
       w2_10, w2_11, w2_12, w2_13, w2_14, w2_15, w2_16, w2_17, w2_18, 
       w2_19, w2_2, w2_20, w2_21, w2_22, w2_23, w2_24, w2_25, w2_26, 
       w2_27, w2_28, w2_29, w2_3, w2_30, w2_31, w2_4, w2_5, w2_6, 
       w2_7, w2_8, w2_9, w3_12, w3_13, w3_14, w3_15, w3_16, w3_17, 
       w3_18, w3_19, w3_20, w3_21, w3_22,  w3_23;
  NAND2_X1 U10 (.A2( ld ) , .ZN( n8 ) , .A1( text_in[3] ) );
  NAND2_X1 U100 (.A2( ld ) , .ZN( n98 ) , .A1( text_in[48] ) );
  XOR2_X1 U1001 (.Z( n728 ) , .B( n729 ) , .A( sa11_sr_0 ) );
  XOR2_X1 U1002 (.Z( n729 ) , .B( sa21_sr_0 ) , .A( w1_17 ) );
  XNOR2_X1 U1004 (.B( n683 ) , .ZN( n730 ) , .A( sa01_sr_1 ) );
  XOR2_X1 U1005 (.A( n163 ) , .Z( n725 ) , .B( w1_17 ) );
  OAI22_X1 U1007 (.ZN( N194 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n731 ) , .B1( n732 ) );
  XOR2_X1 U1009 (.A( n690 ) , .B( n713 ) , .Z( n734 ) );
  OAI21_X1 U101 (.B1( ld ) , .A( n100 ) , .ZN( n1027 ) , .B2( n99 ) );
  XOR2_X1 U1010 (.Z( n713 ) , .A( sa11_sr_7 ) , .B( sa21_sr_7 ) );
  XOR2_X1 U1012 (.A( n161 ) , .Z( n731 ) , .B( w1_16 ) );
  OAI22_X1 U1014 (.ZN( N185 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n735 ) , .B1( n736 ) );
  XOR2_X1 U1016 (.A( n650 ) , .B( n665 ) , .Z( n738 ) );
  XOR2_X1 U1017 (.Z( n650 ) , .A( sa21_sr_6 ) , .B( sa31_sr_6 ) );
  XOR2_X1 U1019 (.A( n159 ) , .Z( n735 ) , .B( w1_15 ) );
  NAND2_X1 U102 (.A2( ld ) , .ZN( n100 ) , .A1( text_in[49] ) );
  OAI22_X1 U1021 (.ZN( N184 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n739 ) , .B1( n740 ) );
  XOR2_X1 U1023 (.A( n644 ) , .B( n656 ) , .Z( n742 ) );
  XOR2_X1 U1024 (.Z( n656 ) , .A( sa21_sr_5 ) , .B( sa31_sr_5 ) );
  XOR2_X1 U1026 (.A( n157 ) , .Z( n739 ) , .B( w1_14 ) );
  OAI22_X1 U1028 (.ZN( N183 ) , .A1( n1109 ) , .B2( n1221 ) , .A2( n743 ) , .B1( n744 ) );
  XOR2_X1 U1029 (.Z( n744 ) , .A( n745 ) , .B( n746 ) );
  OAI21_X1 U103 (.B1( ld ) , .B2( n101 ) , .A( n102 ) , .ZN( n1028 ) );
  XOR2_X1 U1030 (.A( n651 ) , .B( n663 ) , .Z( n746 ) );
  XOR2_X1 U1031 (.Z( n663 ) , .A( sa21_sr_4 ) , .B( sa31_sr_4 ) );
  XNOR2_X1 U1032 (.ZN( n745 ) , .B( sa31_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U1033 (.A( n155 ) , .Z( n743 ) , .B( w1_13 ) );
  OAI22_X1 U1035 (.ZN( N182 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n747 ) , .B1( n748 ) );
  XOR2_X1 U1036 (.Z( n748 ) , .A( n749 ) , .B( n750 ) );
  XOR2_X1 U1037 (.A( n657 ) , .B( n670 ) , .Z( n750 ) );
  XOR2_X1 U1038 (.Z( n670 ) , .A( sa21_sr_3 ) , .B( sa31_sr_3 ) );
  XOR2_X1 U1039 (.B( n643 ) , .Z( n749 ) , .A( n751 ) );
  NAND2_X1 U104 (.A2( ld ) , .ZN( n102 ) , .A1( text_in[50] ) );
  XNOR2_X1 U1040 (.ZN( n751 ) , .B( sa31_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U1041 (.A( n153 ) , .Z( n747 ) , .B( w1_12 ) );
  OAI22_X1 U1043 (.ZN( N181 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n752 ) , .B1( n753 ) );
  XOR2_X1 U1045 (.A( n662 ) , .B( n677 ) , .Z( n755 ) );
  XOR2_X1 U1046 (.Z( n677 ) , .A( sa21_sr_2 ) , .B( sa31_sr_2 ) );
  XNOR2_X1 U1048 (.ZN( n756 ) , .B( sa31_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U1049 (.A( n151 ) , .Z( n752 ) , .B( w1_11 ) );
  OAI21_X1 U105 (.B1( ld ) , .ZN( n1029 ) , .B2( n103 ) , .A( n104 ) );
  OAI22_X1 U1051 (.ZN( N180 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n757 ) , .B1( n758 ) );
  XOR2_X1 U1053 (.A( n671 ) , .B( n683 ) , .Z( n760 ) );
  XOR2_X1 U1054 (.Z( n683 ) , .A( sa21_sr_1 ) , .B( sa31_sr_1 ) );
  XOR2_X1 U1056 (.A( n149 ) , .Z( n757 ) , .B( w1_10 ) );
  OAI22_X1 U1058 (.ZN( N179 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n761 ) , .B1( n762 ) );
  NAND2_X1 U106 (.A2( ld ) , .ZN( n104 ) , .A1( text_in[51] ) );
  XOR2_X1 U1060 (.A( n678 ) , .B( n690 ) , .Z( n764 ) );
  XOR2_X1 U1061 (.Z( n690 ) , .A( sa21_sr_0 ) , .B( sa31_sr_0 ) );
  XNOR2_X1 U1063 (.ZN( n765 ) , .B( sa31_sr_1 ) , .A( w1_9 ) );
  XOR2_X1 U1064 (.A( n147 ) , .Z( n761 ) , .B( w1_9 ) );
  OAI22_X1 U1066 (.ZN( N178 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n766 ) , .B1( n767 ) );
  XOR2_X1 U1068 (.A( n643 ) , .B( n684 ) , .Z( n769 ) );
  XOR2_X1 U1069 (.Z( n643 ) , .A( sa21_sr_7 ) , .B( sa31_sr_7 ) );
  OAI21_X1 U107 (.B1( ld ) , .ZN( n1030 ) , .B2( n105 ) , .A( n106 ) );
  XOR2_X1 U1071 (.A( n145 ) , .Z( n766 ) , .B( w1_8 ) );
  OAI22_X1 U1073 (.ZN( N169 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n770 ) , .B1( n771 ) );
  XOR2_X1 U1074 (.Z( n771 ) , .A( n772 ) , .B( n773 ) );
  XOR2_X1 U1075 (.B( n665 ) , .Z( n773 ) , .A( sa01_sr_6 ) );
  XOR2_X1 U1076 (.Z( n665 ) , .A( sa01_sr_7 ) , .B( sa11_sr_7 ) );
  XNOR2_X1 U1077 (.ZN( n772 ) , .B( n774 ) , .A( sa21_sr_7 ) );
  XOR2_X1 U1078 (.Z( n774 ) , .B( sa31_sr_6 ) , .A( w1_7 ) );
  XOR2_X1 U1079 (.A( n143 ) , .Z( n770 ) , .B( w1_7 ) );
  NAND2_X1 U108 (.A2( ld ) , .ZN( n106 ) , .A1( text_in[52] ) );
  OAI22_X1 U1081 (.ZN( N168 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n775 ) , .B1( n776 ) );
  XOR2_X1 U1082 (.Z( n776 ) , .A( n777 ) , .B( n778 ) );
  XOR2_X1 U1083 (.Z( n778 ) , .B( n779 ) , .A( sa21_sr_6 ) );
  XOR2_X1 U1084 (.Z( n779 ) , .B( sa31_sr_5 ) , .A( w1_6 ) );
  XNOR2_X1 U1085 (.B( n644 ) , .ZN( n777 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U1086 (.Z( n644 ) , .A( sa01_sr_6 ) , .B( sa11_sr_6 ) );
  XOR2_X1 U1087 (.A( n141 ) , .Z( n775 ) , .B( w1_6 ) );
  OAI22_X1 U1089 (.ZN( N167 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n780 ) , .B1( n781 ) );
  OAI21_X1 U109 (.B1( ld ) , .ZN( n1031 ) , .B2( n107 ) , .A( n108 ) );
  XOR2_X1 U1090 (.Z( n781 ) , .A( n782 ) , .B( n783 ) );
  XOR2_X1 U1091 (.Z( n783 ) , .B( n784 ) , .A( sa21_sr_5 ) );
  XOR2_X1 U1092 (.Z( n784 ) , .B( sa31_sr_4 ) , .A( w1_5 ) );
  XNOR2_X1 U1093 (.B( n651 ) , .ZN( n782 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U1094 (.Z( n651 ) , .A( sa01_sr_5 ) , .B( sa11_sr_5 ) );
  XOR2_X1 U1095 (.A( n139 ) , .Z( n780 ) , .B( w1_5 ) );
  OAI22_X1 U1097 (.ZN( N166 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n785 ) , .B1( n786 ) );
  XOR2_X1 U1098 (.Z( n786 ) , .A( n787 ) , .B( n788 ) );
  XOR2_X1 U1099 (.Z( n788 ) , .B( n789 ) , .A( sa21_sr_4 ) );
  OAI21_X1 U11 (.B1( ld ) , .A( n10 ) , .B2( n9 ) , .ZN( n982 ) );
  NAND2_X1 U110 (.A2( ld ) , .ZN( n108 ) , .A1( text_in[53] ) );
  XOR2_X1 U1100 (.Z( n789 ) , .B( sa31_sr_3 ) , .A( w1_4 ) );
  XOR2_X1 U1101 (.Z( n787 ) , .A( n790 ) , .B( n791 ) );
  XNOR2_X1 U1102 (.B( n657 ) , .ZN( n790 ) , .A( sa01_sr_3 ) );
  XOR2_X1 U1103 (.Z( n657 ) , .A( sa01_sr_4 ) , .B( sa11_sr_4 ) );
  XOR2_X1 U1104 (.A( n137 ) , .Z( n785 ) , .B( w1_4 ) );
  OAI22_X1 U1106 (.ZN( N165 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n792 ) , .B1( n793 ) );
  XOR2_X1 U1109 (.Z( n796 ) , .B( sa31_sr_2 ) , .A( w1_3 ) );
  OAI21_X1 U111 (.B1( ld ) , .ZN( n1032 ) , .B2( n109 ) , .A( n110 ) );
  XOR2_X1 U1110 (.B( n791 ) , .Z( n794 ) , .A( n797 ) );
  XNOR2_X1 U1111 (.B( n662 ) , .ZN( n797 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U1112 (.Z( n662 ) , .A( sa01_sr_3 ) , .B( sa11_sr_3 ) );
  XOR2_X1 U1113 (.A( n135 ) , .Z( n792 ) , .B( w1_3 ) );
  OAI22_X1 U1115 (.ZN( N164 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n798 ) , .B1( n799 ) );
  XOR2_X1 U1116 (.Z( n799 ) , .A( n800 ) , .B( n801 ) );
  XOR2_X1 U1117 (.Z( n801 ) , .B( n802 ) , .A( sa21_sr_2 ) );
  XOR2_X1 U1118 (.Z( n802 ) , .B( sa31_sr_1 ) , .A( w1_2 ) );
  XNOR2_X1 U1119 (.B( n671 ) , .ZN( n800 ) , .A( sa01_sr_1 ) );
  NAND2_X1 U112 (.A2( ld ) , .ZN( n110 ) , .A1( text_in[54] ) );
  XOR2_X1 U1120 (.Z( n671 ) , .A( sa01_sr_2 ) , .B( sa11_sr_2 ) );
  XOR2_X1 U1121 (.A( n133 ) , .Z( n798 ) , .B( w1_2 ) );
  OAI22_X1 U1123 (.ZN( N163 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n803 ) , .B1( n804 ) );
  XOR2_X1 U1125 (.Z( n806 ) , .B( n807 ) , .A( sa21_sr_1 ) );
  XOR2_X1 U1126 (.Z( n807 ) , .B( sa31_sr_0 ) , .A( w1_1 ) );
  XNOR2_X1 U1128 (.B( n678 ) , .ZN( n808 ) , .A( sa01_sr_0 ) );
  XOR2_X1 U1129 (.Z( n678 ) , .A( sa01_sr_1 ) , .B( sa11_sr_1 ) );
  OAI21_X1 U113 (.B1( ld ) , .ZN( n1033 ) , .B2( n111 ) , .A( n112 ) );
  XOR2_X1 U1130 (.A( n131 ) , .Z( n803 ) , .B( w1_1 ) );
  OAI22_X1 U1132 (.ZN( N162 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n809 ) , .B1( n810 ) );
  XOR2_X1 U1134 (.A( n684 ) , .B( n791 ) , .Z( n812 ) );
  XOR2_X1 U1135 (.Z( n791 ) , .A( sa01_sr_7 ) , .B( sa31_sr_7 ) );
  XOR2_X1 U1136 (.Z( n684 ) , .A( sa01_sr_0 ) , .B( sa11_sr_0 ) );
  XOR2_X1 U1138 (.A( n129 ) , .Z( n809 ) , .B( w1_0 ) );
  NAND2_X1 U114 (.A2( ld ) , .ZN( n112 ) , .A1( text_in[55] ) );
  OAI22_X1 U1140 (.ZN( N153 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n813 ) , .B1( n814 ) );
  XOR2_X1 U1142 (.Z( n816 ) , .A( n817 ) , .B( n818 ) );
  INV_X1 U1144 (.ZN( n819 ) , .A( sa12_sr_7 ) );
  XOR2_X1 U1145 (.A( n127 ) , .Z( n813 ) , .B( w2_31 ) );
  OAI22_X1 U1147 (.ZN( N152 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n820 ) , .B1( n821 ) );
  XOR2_X1 U1149 (.Z( n823 ) , .A( n824 ) , .B( n825 ) );
  OAI21_X1 U115 (.B1( ld ) , .ZN( n1034 ) , .B2( n113 ) , .A( n114 ) );
  XOR2_X1 U1151 (.A( n125 ) , .Z( n820 ) , .B( w2_30 ) );
  OAI22_X1 U1153 (.ZN( N151 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n826 ) , .B1( n827 ) );
  XOR2_X1 U1154 (.Z( n827 ) , .A( n828 ) , .B( n829 ) );
  XOR2_X1 U1155 (.Z( n829 ) , .A( n830 ) , .B( n831 ) );
  XNOR2_X1 U1156 (.ZN( n828 ) , .B( sa12_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U1157 (.A( n123 ) , .Z( n826 ) , .B( w2_29 ) );
  OAI22_X1 U1159 (.ZN( N150 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n832 ) , .B1( n833 ) );
  NAND2_X1 U116 (.A2( ld ) , .ZN( n114 ) , .A1( text_in[56] ) );
  XOR2_X1 U1160 (.Z( n833 ) , .A( n834 ) , .B( n835 ) );
  XOR2_X1 U1161 (.Z( n835 ) , .A( n836 ) , .B( n837 ) );
  XOR2_X1 U1162 (.Z( n834 ) , .A( n838 ) , .B( n839 ) );
  XNOR2_X1 U1163 (.ZN( n838 ) , .B( sa12_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U1164 (.A( n121 ) , .Z( n832 ) , .B( w2_28 ) );
  OAI22_X1 U1166 (.ZN( N149 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n840 ) , .B1( n841 ) );
  XOR2_X1 U1168 (.Z( n843 ) , .B( n844 ) , .A( n845 ) );
  OAI21_X1 U117 (.B1( ld ) , .ZN( n1035 ) , .B2( n115 ) , .A( n116 ) );
  XNOR2_X1 U1170 (.ZN( n846 ) , .B( sa12_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U1171 (.A( n119 ) , .Z( n840 ) , .B( w2_27 ) );
  OAI22_X1 U1173 (.ZN( N148 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n847 ) , .B1( n848 ) );
  XOR2_X1 U1175 (.A( n277 ) , .Z( n850 ) , .B( n851 ) );
  XOR2_X1 U1177 (.A( n117 ) , .Z( n847 ) , .B( w2_26 ) );
  OAI22_X1 U1179 (.ZN( N147 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n852 ) , .B1( n853 ) );
  NAND2_X1 U118 (.A2( ld ) , .ZN( n116 ) , .A1( text_in[57] ) );
  XOR2_X1 U1182 (.B( n284 ) , .Z( n854 ) , .A( n857 ) );
  XNOR2_X1 U1183 (.ZN( n857 ) , .B( sa12_sr_1 ) , .A( w2_25 ) );
  XOR2_X1 U1184 (.A( n115 ) , .Z( n852 ) , .B( w2_25 ) );
  OAI22_X1 U1186 (.ZN( N146 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n858 ) , .B1( n859 ) );
  XOR2_X1 U1188 (.A( n836 ) , .Z( n861 ) , .B( n862 ) );
  OAI21_X1 U119 (.B1( ld ) , .ZN( n1036 ) , .B2( n117 ) , .A( n118 ) );
  XOR2_X1 U1190 (.A( n113 ) , .Z( n858 ) , .B( w2_24 ) );
  OAI22_X1 U1192 (.ZN( N137 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n863 ) , .B1( n864 ) );
  XOR2_X1 U1193 (.Z( n864 ) , .A( n865 ) , .B( n866 ) );
  XOR2_X1 U1194 (.B( n817 ) , .Z( n866 ) , .A( sa02_sr_7 ) );
  XNOR2_X1 U1195 (.ZN( n865 ) , .B( n867 ) , .A( sa12_sr_6 ) );
  XOR2_X1 U1196 (.Z( n867 ) , .B( sa22_sr_6 ) , .A( w2_23 ) );
  XOR2_X1 U1197 (.A( n111 ) , .Z( n863 ) , .B( w2_23 ) );
  OAI22_X1 U1199 (.ZN( N136 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n868 ) , .B1( n869 ) );
  NAND2_X1 U12 (.A2( ld ) , .ZN( n10 ) , .A1( text_in[4] ) );
  NAND2_X1 U120 (.A2( ld ) , .ZN( n118 ) , .A1( text_in[58] ) );
  XOR2_X1 U1202 (.Z( n872 ) , .B( sa22_sr_5 ) , .A( w2_22 ) );
  XOR2_X1 U1205 (.A( n109 ) , .Z( n868 ) , .B( w2_22 ) );
  OAI22_X1 U1207 (.ZN( N135 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n874 ) , .B1( n875 ) );
  XOR2_X1 U1208 (.Z( n875 ) , .A( n876 ) , .B( n877 ) );
  XOR2_X1 U1209 (.Z( n877 ) , .B( n878 ) , .A( sa12_sr_4 ) );
  OAI21_X1 U121 (.B1( ld ) , .ZN( n1037 ) , .B2( n119 ) , .A( n120 ) );
  XOR2_X1 U1210 (.Z( n878 ) , .B( sa22_sr_4 ) , .A( w2_21 ) );
  XNOR2_X1 U1211 (.B( n831 ) , .ZN( n876 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1212 (.A( n107 ) , .Z( n874 ) , .B( w2_21 ) );
  OAI22_X1 U1214 (.ZN( N134 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n879 ) , .B1( n880 ) );
  XOR2_X1 U1215 (.Z( n880 ) , .A( n881 ) , .B( n882 ) );
  XOR2_X1 U1216 (.Z( n882 ) , .B( n883 ) , .A( sa12_sr_3 ) );
  XOR2_X1 U1217 (.Z( n883 ) , .B( sa22_sr_3 ) , .A( w2_20 ) );
  XOR2_X1 U1218 (.Z( n881 ) , .A( n884 ) , .B( n885 ) );
  XNOR2_X1 U1219 (.B( n839 ) , .ZN( n884 ) , .A( sa02_sr_4 ) );
  NAND2_X1 U122 (.A2( ld ) , .ZN( n120 ) , .A1( text_in[59] ) );
  XOR2_X1 U1220 (.A( n105 ) , .Z( n879 ) , .B( w2_20 ) );
  OAI22_X1 U1222 (.ZN( N133 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n886 ) , .B1( n887 ) );
  XOR2_X1 U1223 (.Z( n887 ) , .A( n888 ) , .B( n889 ) );
  XOR2_X1 U1224 (.Z( n889 ) , .B( n890 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1225 (.Z( n890 ) , .B( sa22_sr_2 ) , .A( w2_19 ) );
  XOR2_X1 U1228 (.A( n103 ) , .Z( n886 ) , .B( w2_19 ) );
  OAI21_X1 U123 (.B1( ld ) , .ZN( n1038 ) , .B2( n121 ) , .A( n122 ) );
  OAI22_X1 U1230 (.ZN( N132 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n892 ) , .B1( n893 ) );
  XOR2_X1 U1233 (.Z( n896 ) , .B( sa22_sr_1 ) , .A( w2_18 ) );
  XOR2_X1 U1236 (.A( n101 ) , .Z( n892 ) , .B( w2_18 ) );
  OAI22_X1 U1238 (.ZN( N131 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n898 ) , .B1( n899 ) );
  XOR2_X1 U1239 (.Z( n899 ) , .A( n900 ) , .B( n901 ) );
  NAND2_X1 U124 (.A2( ld ) , .ZN( n122 ) , .A1( text_in[60] ) );
  XOR2_X1 U1240 (.Z( n901 ) , .B( n902 ) , .A( sa12_sr_0 ) );
  XOR2_X1 U1241 (.Z( n902 ) , .B( sa22_sr_0 ) , .A( w2_17 ) );
  XOR2_X1 U1242 (.B( n885 ) , .Z( n900 ) , .A( n903 ) );
  XNOR2_X1 U1243 (.B( n856 ) , .ZN( n903 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1244 (.Z( n898 ) , .A( n99 ) , .B( w2_17 ) );
  OAI22_X1 U1246 (.ZN( N130 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n904 ) , .B1( n905 ) );
  XOR2_X1 U1248 (.A( n862 ) , .B( n885 ) , .Z( n907 ) );
  XOR2_X1 U1249 (.Z( n885 ) , .A( sa12_sr_7 ) , .B( sa22_sr_7 ) );
  OAI21_X1 U125 (.B1( ld ) , .ZN( n1039 ) , .B2( n123 ) , .A( n124 ) );
  XOR2_X1 U1251 (.Z( n904 ) , .A( n97 ) , .B( w2_16 ) );
  OAI22_X1 U1253 (.ZN( N121 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n908 ) , .B1( n909 ) );
  XOR2_X1 U1255 (.A( n824 ) , .B( n836 ) , .Z( n911 ) );
  XOR2_X1 U1256 (.Z( n824 ) , .A( sa22_sr_6 ) , .B( sa32_sr_6 ) );
  XOR2_X1 U1258 (.Z( n908 ) , .A( n95 ) , .B( w2_15 ) );
  NAND2_X1 U126 (.A2( ld ) , .ZN( n124 ) , .A1( text_in[61] ) );
  OAI22_X1 U1260 (.ZN( N120 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n912 ) , .B1( n913 ) );
  XOR2_X1 U1262 (.A( n818 ) , .B( n831 ) , .Z( n915 ) );
  XOR2_X1 U1263 (.Z( n831 ) , .A( sa22_sr_5 ) , .B( sa32_sr_5 ) );
  XOR2_X1 U1265 (.Z( n912 ) , .A( n93 ) , .B( w2_14 ) );
  OAI22_X1 U1267 (.ZN( N119 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n916 ) , .B1( n917 ) );
  XOR2_X1 U1268 (.Z( n917 ) , .A( n918 ) , .B( n919 ) );
  XOR2_X1 U1269 (.A( n825 ) , .B( n839 ) , .Z( n919 ) );
  OAI21_X1 U127 (.B1( ld ) , .ZN( n1040 ) , .B2( n125 ) , .A( n126 ) );
  XOR2_X1 U1270 (.Z( n839 ) , .A( sa22_sr_4 ) , .B( sa32_sr_4 ) );
  XNOR2_X1 U1271 (.ZN( n918 ) , .B( sa32_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U1272 (.A( n91 ) , .Z( n916 ) , .B( w2_13 ) );
  OAI22_X1 U1274 (.ZN( N118 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n920 ) , .B1( n921 ) );
  XOR2_X1 U1275 (.Z( n921 ) , .A( n922 ) , .B( n923 ) );
  XOR2_X1 U1276 (.A( n830 ) , .B( n844 ) , .Z( n923 ) );
  XOR2_X1 U1277 (.Z( n844 ) , .A( sa22_sr_3 ) , .B( sa32_sr_3 ) );
  INV_X1 U1278 (.ZN( n830 ) , .A( n924 ) );
  XOR2_X1 U1279 (.B( n817 ) , .Z( n922 ) , .A( n925 ) );
  NAND2_X1 U128 (.A2( ld ) , .ZN( n126 ) , .A1( text_in[62] ) );
  XNOR2_X1 U1280 (.ZN( n925 ) , .B( sa32_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U1281 (.A( n89 ) , .Z( n920 ) , .B( w2_12 ) );
  OAI22_X1 U1283 (.ZN( N117 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n926 ) , .B1( n927 ) );
  XOR2_X1 U1285 (.A( n837 ) , .B( n851 ) , .Z( n929 ) );
  INV_X1 U1287 (.ZN( n837 ) , .A( n930 ) );
  XNOR2_X1 U1289 (.ZN( n931 ) , .B( sa32_sr_3 ) , .A( w2_11 ) );
  OAI21_X1 U129 (.B1( ld ) , .ZN( n1041 ) , .B2( n127 ) , .A( n128 ) );
  XOR2_X1 U1290 (.A( n87 ) , .Z( n926 ) , .B( w2_11 ) );
  OAI22_X1 U1292 (.ZN( N116 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n932 ) , .B1( n933 ) );
  XOR2_X1 U1294 (.A( n845 ) , .B( n856 ) , .Z( n935 ) );
  XOR2_X1 U1295 (.Z( n856 ) , .A( sa22_sr_1 ) , .B( sa32_sr_1 ) );
  XOR2_X1 U1297 (.A( n85 ) , .Z( n932 ) , .B( w2_10 ) );
  OAI22_X1 U1299 (.ZN( N115 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n936 ) , .B1( n937 ) );
  OAI21_X1 U13 (.B1( ld ) , .B2( n11 ) , .A( n12 ) , .ZN( n983 ) );
  NAND2_X1 U130 (.A2( ld ) , .ZN( n128 ) , .A1( text_in[63] ) );
  XOR2_X1 U1301 (.A( n817 ) , .B( n862 ) , .Z( n939 ) );
  XOR2_X1 U1302 (.Z( n862 ) , .A( sa22_sr_0 ) , .B( sa32_sr_0 ) );
  XOR2_X1 U1304 (.Z( n277 ) , .A( sa02_sr_1 ) , .B( sa12_sr_1 ) );
  XNOR2_X1 U1305 (.ZN( n940 ) , .B( sa32_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U1306 (.A( n83 ) , .Z( n936 ) , .B( w2_9 ) );
  OAI22_X1 U1308 (.ZN( N114 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n941 ) , .B1( n942 ) );
  OAI21_X1 U131 (.B1( ld ) , .ZN( n1042 ) , .B2( n129 ) , .A( n130 ) );
  XOR2_X1 U1310 (.A( n284 ) , .B( n817 ) , .Z( n944 ) );
  XOR2_X1 U1311 (.Z( n817 ) , .A( sa22_sr_7 ) , .B( sa32_sr_7 ) );
  XOR2_X1 U1312 (.Z( n284 ) , .A( sa02_sr_0 ) , .B( sa12_sr_0 ) );
  XOR2_X1 U1314 (.A( n81 ) , .Z( n941 ) , .B( w2_8 ) );
  OAI22_X1 U1316 (.ZN( N105 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n945 ) , .B1( n946 ) );
  XOR2_X1 U1317 (.Z( n946 ) , .A( n947 ) , .B( n948 ) );
  XOR2_X1 U1318 (.B( n836 ) , .Z( n948 ) , .A( sa02_sr_6 ) );
  XOR2_X1 U1319 (.Z( n836 ) , .A( sa02_sr_7 ) , .B( sa12_sr_7 ) );
  NAND2_X1 U132 (.A2( ld ) , .ZN( n130 ) , .A1( text_in[64] ) );
  XNOR2_X1 U1320 (.ZN( n947 ) , .B( n949 ) , .A( sa22_sr_7 ) );
  XOR2_X1 U1321 (.Z( n949 ) , .B( sa32_sr_6 ) , .A( w2_7 ) );
  XOR2_X1 U1322 (.A( n79 ) , .Z( n945 ) , .B( w2_7 ) );
  OAI22_X1 U1324 (.ZN( N104 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n950 ) , .B1( n951 ) );
  XOR2_X1 U1327 (.Z( n954 ) , .B( sa32_sr_5 ) , .A( w2_6 ) );
  XNOR2_X1 U1328 (.B( n818 ) , .ZN( n952 ) , .A( sa02_sr_5 ) );
  XOR2_X1 U1329 (.Z( n818 ) , .A( sa02_sr_6 ) , .B( sa12_sr_6 ) );
  OAI21_X1 U133 (.B1( ld ) , .ZN( n1043 ) , .B2( n131 ) , .A( n132 ) );
  XOR2_X1 U1330 (.A( n77 ) , .Z( n950 ) , .B( w2_6 ) );
  OAI22_X1 U1332 (.ZN( N103 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n955 ) , .B1( n956 ) );
  XOR2_X1 U1333 (.Z( n956 ) , .A( n957 ) , .B( n958 ) );
  XOR2_X1 U1334 (.Z( n958 ) , .B( n959 ) , .A( sa22_sr_5 ) );
  XOR2_X1 U1335 (.Z( n959 ) , .B( sa32_sr_4 ) , .A( w2_5 ) );
  XNOR2_X1 U1336 (.B( n825 ) , .ZN( n957 ) , .A( sa02_sr_4 ) );
  XOR2_X1 U1337 (.Z( n825 ) , .A( sa02_sr_5 ) , .B( sa12_sr_5 ) );
  XOR2_X1 U1338 (.A( n75 ) , .Z( n955 ) , .B( w2_5 ) );
  NAND2_X1 U134 (.A2( ld ) , .ZN( n132 ) , .A1( text_in[65] ) );
  OAI22_X1 U1340 (.ZN( N102 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n960 ) , .B1( n961 ) );
  XOR2_X1 U1343 (.Z( n964 ) , .B( sa32_sr_3 ) , .A( w2_4 ) );
  XOR2_X1 U1344 (.A( n924 ) , .Z( n962 ) , .B( n965 ) );
  XOR2_X1 U1345 (.B( n279 ) , .Z( n965 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1346 (.ZN( n924 ) , .A( sa02_sr_4 ) , .B( sa12_sr_4 ) );
  XOR2_X1 U1347 (.A( n73 ) , .Z( n960 ) , .B( w2_4 ) );
  OAI22_X1 U1349 (.ZN( N101 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n966 ) , .B1( n967 ) );
  OAI21_X1 U135 (.B1( ld ) , .ZN( n1044 ) , .B2( n133 ) , .A( n134 ) );
  XOR2_X1 U1351 (.Z( n969 ) , .B( n970 ) , .A( sa22_sr_3 ) );
  XOR2_X1 U1352 (.Z( n970 ) , .B( sa32_sr_2 ) , .A( w2_3 ) );
  XOR2_X1 U1354 (.B( n279 ) , .Z( n971 ) , .A( sa02_sr_2 ) );
  XOR2_X1 U1355 (.Z( n279 ) , .A( sa02_sr_7 ) , .B( sa32_sr_7 ) );
  XNOR2_X1 U1356 (.ZN( n930 ) , .A( sa02_sr_3 ) , .B( sa12_sr_3 ) );
  XOR2_X1 U1357 (.A( n71 ) , .Z( n966 ) , .B( w2_3 ) );
  OAI22_X1 U1359 (.ZN( N100 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n972 ) , .B1( n973 ) );
  NAND2_X1 U136 (.A2( ld ) , .ZN( n134 ) , .A1( text_in[66] ) );
  XOR2_X1 U1361 (.Z( n973 ) , .A( n974 ) , .B( n975 ) );
  XOR2_X1 U1362 (.Z( n975 ) , .B( n976 ) , .A( sa22_sr_2 ) );
  XOR2_X1 U1363 (.Z( n976 ) , .B( sa32_sr_1 ) , .A( w2_2 ) );
  XNOR2_X1 U1364 (.B( n845 ) , .ZN( n974 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1365 (.Z( n845 ) , .B( sa02_sr_2 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1366 (.A( n69 ) , .Z( n972 ) , .B( w2_2 ) );
  CLKBUF_X1 U1368 (.Z( n1219 ) , .A( n1220 ) );
  CLKBUF_X1 U1369 (.A( n1109 ) , .Z( n1212 ) );
  OAI21_X1 U137 (.B1( ld ) , .ZN( n1045 ) , .B2( n135 ) , .A( n136 ) );
  XOR2_X1 U1370 (.A( n1115 ) , .Z( n382 ) , .B( n384 ) );
  XOR2_X1 U1371 (.Z( n1115 ) , .B( n386 ) , .A( w3_16 ) );
  XNOR2_X1 U1372 (.B( n1116 ) , .ZN( n338 ) , .A( sa13_sr_6 ) );
  XOR2_X1 U1373 (.Z( n1116 ) , .B( sa23_sr_6 ) , .A( w3_23 ) );
  XOR2_X1 U1374 (.Z( N495 ) , .B( sa32_sr_2 ) , .A( w2_2 ) );
  XNOR2_X1 U1375 (.A( n1117 ) , .B( n885 ) , .ZN( n888 ) );
  XOR2_X1 U1376 (.Z( n1117 ) , .B( n844 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1377 (.A( n1118 ) , .B( n539 ) , .ZN( n542 ) );
  XOR2_X1 U1378 (.Z( n1118 ) , .B( n496 ) , .A( sa00_sr_3 ) );
  XNOR2_X1 U1379 (.B( n476 ) , .ZN( n524 ) , .A( sa00_sr_6 ) );
  NAND2_X1 U138 (.A2( ld ) , .ZN( n136 ) , .A1( text_in[67] ) );
  XNOR2_X1 U1380 (.B( n824 ) , .ZN( n870 ) , .A( sa02_sr_6 ) );
  XNOR2_X1 U1381 (.B( n650 ) , .ZN( n698 ) , .A( sa01_sr_6 ) );
  XNOR2_X1 U1382 (.B( n295 ) , .ZN( n343 ) , .A( sa03_sr_6 ) );
  XNOR2_X1 U1383 (.B( n851 ) , .ZN( n894 ) , .A( sa02_sr_2 ) );
  INV_X1 U1384 (.A( n1114 ) , .ZN( n1214 ) );
  BUF_X1 U1385 (.Z( n1217 ) , .A( n1221 ) );
  BUF_X1 U1386 (.Z( n1218 ) , .A( n1221 ) );
  XNOR2_X1 U1387 (.A( n1119 ) , .ZN( n405 ) , .B( n407 ) );
  XNOR2_X1 U1388 (.ZN( n1119 ) , .B( n289 ) , .A( n408 ) );
  XNOR2_X1 U1389 (.A( n1120 ) , .ZN( n312 ) , .B( n314 ) );
  OAI21_X1 U139 (.B1( ld ) , .ZN( n1046 ) , .B2( n137 ) , .A( n138 ) );
  XNOR2_X1 U1390 (.ZN( n1120 ) , .B( n307 ) , .A( n317 ) );
  XNOR2_X1 U1391 (.A( n1121 ) , .ZN( n392 ) , .B( n394 ) );
  XOR2_X1 U1392 (.Z( n1121 ) , .B( sa33_sr_6 ) , .A( w3_14 ) );
  XNOR2_X1 U1393 (.B( n1122 ) , .ZN( n428 ) , .A( n429 ) );
  XNOR2_X1 U1394 (.ZN( n1122 ) , .B( n431 ) , .A( sa23_sr_6 ) );
  XNOR2_X1 U1395 (.A( n1123 ) , .ZN( n388 ) , .B( n390 ) );
  XOR2_X1 U1396 (.Z( n1123 ) , .B( sa33_sr_7 ) , .A( w3_15 ) );
  XNOR2_X1 U1397 (.A( n1124 ) , .ZN( n396 ) , .B( n398 ) );
  XOR2_X1 U1398 (.Z( n1124 ) , .B( sa33_sr_5 ) , .A( w3_13 ) );
  INV_X1 U1399 (.A( n1213 ) , .ZN( n1221 ) );
  NAND2_X1 U14 (.A2( ld ) , .ZN( n12 ) , .A1( text_in[5] ) );
  NAND2_X1 U140 (.A2( ld ) , .ZN( n138 ) , .A1( text_in[68] ) );
  INV_X1 U1400 (.A( n1212 ) , .ZN( n1220 ) );
  XNOR2_X1 U1401 (.A( n1125 ) , .ZN( n753 ) , .B( n755 ) );
  XNOR2_X1 U1402 (.ZN( n1125 ) , .B( n643 ) , .A( n756 ) );
  XNOR2_X1 U1403 (.A( n1126 ) , .ZN( n493 ) , .B( n495 ) );
  XNOR2_X1 U1404 (.ZN( n1126 ) , .B( n488 ) , .A( n498 ) );
  XNOR2_X1 U1405 (.A( n1127 ) , .ZN( n841 ) , .B( n843 ) );
  XNOR2_X1 U1406 (.ZN( n1127 ) , .B( n836 ) , .A( n846 ) );
  XNOR2_X1 U1407 (.A( n1128 ) , .ZN( n933 ) , .B( n935 ) );
  XOR2_X1 U1408 (.Z( n1128 ) , .B( sa32_sr_2 ) , .A( w2_10 ) );
  XNOR2_X1 U1409 (.A( n1129 ) , .ZN( n667 ) , .B( n669 ) );
  OAI21_X1 U141 (.B1( ld ) , .ZN( n1047 ) , .B2( n139 ) , .A( n140 ) );
  XNOR2_X1 U1410 (.ZN( n1129 ) , .B( n665 ) , .A( n672 ) );
  XNOR2_X1 U1411 (.A( n1130 ) , .ZN( n848 ) , .B( n850 ) );
  XOR2_X1 U1412 (.Z( n1130 ) , .B( sa12_sr_2 ) , .A( w2_26 ) );
  XNOR2_X1 U1413 (.B( n1131 ) , .ZN( n602 ) , .A( n603 ) );
  XNOR2_X1 U1414 (.ZN( n1131 ) , .B( n605 ) , .A( sa20_sr_6 ) );
  XNOR2_X1 U1415 (.A( n1132 ) , .ZN( n479 ) , .B( n481 ) );
  XOR2_X1 U1416 (.Z( n1132 ) , .B( sa10_sr_5 ) , .A( w0_29 ) );
  XNOR2_X1 U1417 (.A( n1133 ) , .ZN( n272 ) , .B( n275 ) );
  XOR2_X1 U1418 (.Z( n1133 ) , .A( n277 ) , .B( n278 ) );
  XNOR2_X1 U1419 (.B( n1134 ) , .ZN( n433 ) , .A( n434 ) );
  NAND2_X1 U142 (.A2( ld ) , .ZN( n140 ) , .A1( text_in[69] ) );
  XNOR2_X1 U1420 (.ZN( n1134 ) , .B( n436 ) , .A( sa23_sr_5 ) );
  XNOR2_X1 U1421 (.A( n1135 ) , .ZN( n579 ) , .B( n581 ) );
  XNOR2_X1 U1422 (.ZN( n1135 ) , .B( n469 ) , .A( n582 ) );
  XNOR2_X1 U1423 (.A( n1136 ) , .ZN( n814 ) , .B( n816 ) );
  XNOR2_X1 U1424 (.ZN( n1136 ) , .B( n819 ) , .A( w2_31 ) );
  XNOR2_X1 U1425 (.A( n1137 ) , .ZN( n325 ) , .B( n327 ) );
  XNOR2_X1 U1426 (.ZN( n1137 ) , .B( n307 ) , .A( n330 ) );
  XNOR2_X1 U1427 (.A( n1138 ) , .ZN( n927 ) , .B( n929 ) );
  XNOR2_X1 U1428 (.ZN( n1138 ) , .B( n817 ) , .A( n931 ) );
  XNOR2_X1 U1429 (.B( n1139 ) , .ZN( n893 ) , .A( n894 ) );
  OAI21_X1 U143 (.B1( ld ) , .ZN( n1048 ) , .B2( n141 ) , .A( n142 ) );
  XNOR2_X1 U1430 (.ZN( n1139 ) , .B( n896 ) , .A( sa12_sr_1 ) );
  XNOR2_X1 U1431 (.B( n1140 ) , .ZN( n445 ) , .A( n446 ) );
  XNOR2_X1 U1432 (.ZN( n1140 ) , .B( n448 ) , .A( sa23_sr_3 ) );
  XNOR2_X1 U1433 (.B( n1141 ) , .ZN( n362 ) , .A( n363 ) );
  XNOR2_X1 U1434 (.ZN( n1141 ) , .B( n365 ) , .A( sa13_sr_2 ) );
  XNOR2_X1 U1435 (.B( n1142 ) , .ZN( n369 ) , .A( n370 ) );
  XNOR2_X1 U1436 (.ZN( n1142 ) , .B( n372 ) , .A( sa13_sr_1 ) );
  XNOR2_X1 U1437 (.B( n1143 ) , .ZN( n715 ) , .A( n716 ) );
  XNOR2_X1 U1438 (.ZN( n1143 ) , .B( n718 ) , .A( sa11_sr_2 ) );
  XNOR2_X1 U1439 (.A( n1144 ) , .ZN( n500 ) , .B( n502 ) );
  NAND2_X1 U144 (.A2( ld ) , .ZN( n142 ) , .A1( text_in[70] ) );
  XOR2_X1 U1440 (.Z( n1144 ) , .B( sa10_sr_2 ) , .A( w0_26 ) );
  XNOR2_X1 U1441 (.A( n1145 ) , .ZN( n967 ) , .B( n969 ) );
  XNOR2_X1 U1442 (.ZN( n1145 ) , .A( n930 ) , .B( n971 ) );
  XNOR2_X1 U1443 (.A( n1146 ) , .ZN( n640 ) , .B( n642 ) );
  XNOR2_X1 U1444 (.ZN( n1146 ) , .B( n645 ) , .A( w1_31 ) );
  XNOR2_X1 U1445 (.A( n1147 ) , .ZN( n687 ) , .B( n689 ) );
  XOR2_X1 U1446 (.Z( n1147 ) , .B( sa11_sr_0 ) , .A( w1_24 ) );
  XNOR2_X1 U1447 (.A( n1148 ) , .ZN( n281 ) , .B( n283 ) );
  XOR2_X1 U1448 (.Z( n1148 ) , .B( sa22_sr_0 ) , .A( w2_0 ) );
  XNOR2_X1 U1449 (.B( n1149 ) , .ZN( n619 ) , .A( n620 ) );
  OAI21_X1 U145 (.B1( ld ) , .ZN( n1049 ) , .B2( n143 ) , .A( n144 ) );
  XNOR2_X1 U1450 (.ZN( n1149 ) , .B( n622 ) , .A( sa20_sr_3 ) );
  XNOR2_X1 U1451 (.A( n1150 ) , .ZN( n937 ) , .B( n939 ) );
  XNOR2_X1 U1452 (.ZN( n1150 ) , .B( n277 ) , .A( n940 ) );
  XNOR2_X1 U1453 (.A( n1151 ) , .ZN( n859 ) , .B( n861 ) );
  XOR2_X1 U1454 (.Z( n1151 ) , .B( sa12_sr_0 ) , .A( w2_24 ) );
  XNOR2_X1 U1455 (.A( n1152 ) , .ZN( n736 ) , .B( n738 ) );
  XOR2_X1 U1456 (.Z( n1152 ) , .B( sa31_sr_7 ) , .A( w1_15 ) );
  XNOR2_X1 U1457 (.A( n1153 ) , .ZN( n562 ) , .B( n564 ) );
  XOR2_X1 U1458 (.Z( n1153 ) , .B( sa30_sr_7 ) , .A( w0_15 ) );
  XNOR2_X1 U1459 (.A( n1154 ) , .ZN( n909 ) , .B( n911 ) );
  NAND2_X1 U146 (.A2( ld ) , .ZN( n144 ) , .A1( text_in[71] ) );
  XOR2_X1 U1460 (.Z( n1154 ) , .B( sa32_sr_7 ) , .A( w2_15 ) );
  XNOR2_X1 U1461 (.A( n1155 ) , .ZN( n473 ) , .B( n475 ) );
  XOR2_X1 U1462 (.Z( n1155 ) , .B( sa10_sr_6 ) , .A( w0_30 ) );
  XNOR2_X1 U1463 (.A( n1156 ) , .ZN( n821 ) , .B( n823 ) );
  XOR2_X1 U1464 (.Z( n1156 ) , .B( sa12_sr_6 ) , .A( w2_30 ) );
  XNOR2_X1 U1465 (.A( n1157 ) , .ZN( n647 ) , .B( n649 ) );
  XOR2_X1 U1466 (.Z( n1157 ) , .B( sa11_sr_6 ) , .A( w1_30 ) );
  XNOR2_X1 U1467 (.A( n1158 ) , .ZN( n588 ) , .B( n590 ) );
  XNOR2_X1 U1468 (.ZN( n1158 ) , .B( n469 ) , .A( n591 ) );
  XNOR2_X1 U1469 (.A( n1159 ) , .ZN( n762 ) , .B( n764 ) );
  OAI21_X1 U147 (.B1( ld ) , .ZN( n1050 ) , .B2( n145 ) , .A( n146 ) );
  XNOR2_X1 U1470 (.ZN( n1159 ) , .B( n643 ) , .A( n765 ) );
  XNOR2_X1 U1471 (.B( n1160 ) , .ZN( n523 ) , .A( n524 ) );
  XNOR2_X1 U1472 (.ZN( n1160 ) , .B( n526 ) , .A( sa10_sr_5 ) );
  XNOR2_X1 U1473 (.B( n1161 ) , .ZN( n869 ) , .A( n870 ) );
  XNOR2_X1 U1474 (.ZN( n1161 ) , .B( n872 ) , .A( sa12_sr_5 ) );
  XNOR2_X1 U1475 (.B( n1162 ) , .ZN( n697 ) , .A( n698 ) );
  XNOR2_X1 U1476 (.ZN( n1162 ) , .B( n700 ) , .A( sa11_sr_5 ) );
  XNOR2_X1 U1477 (.A( n1163 ) , .ZN( n740 ) , .B( n742 ) );
  XOR2_X1 U1478 (.Z( n1163 ) , .B( sa31_sr_6 ) , .A( w1_14 ) );
  XNOR2_X1 U1479 (.A( n1164 ) , .ZN( n913 ) , .B( n915 ) );
  NAND2_X1 U148 (.A2( ld ) , .ZN( n146 ) , .A1( text_in[72] ) );
  XOR2_X1 U1480 (.Z( n1164 ) , .B( sa32_sr_6 ) , .A( w2_14 ) );
  XNOR2_X1 U1481 (.A( n1165 ) , .ZN( n414 ) , .B( n416 ) );
  XNOR2_X1 U1482 (.ZN( n1165 ) , .B( n289 ) , .A( n417 ) );
  XNOR2_X1 U1483 (.A( n1166 ) , .ZN( n506 ) , .B( n508 ) );
  XNOR2_X1 U1484 (.ZN( n1166 ) , .B( n488 ) , .A( n511 ) );
  XNOR2_X1 U1485 (.B( n1167 ) , .ZN( n793 ) , .A( n794 ) );
  XNOR2_X1 U1486 (.ZN( n1167 ) , .B( n796 ) , .A( sa21_sr_3 ) );
  XNOR2_X1 U1487 (.A( n1168 ) , .ZN( n942 ) , .B( n944 ) );
  XOR2_X1 U1488 (.Z( n1168 ) , .B( sa32_sr_0 ) , .A( w2_8 ) );
  XNOR2_X1 U1489 (.A( n1169 ) , .ZN( n566 ) , .B( n568 ) );
  OAI21_X1 U149 (.B1( ld ) , .ZN( n1051 ) , .B2( n147 ) , .A( n148 ) );
  XOR2_X1 U1490 (.Z( n1169 ) , .B( sa30_sr_6 ) , .A( w0_14 ) );
  XNOR2_X1 U1491 (.A( n1170 ) , .ZN( n767 ) , .B( n769 ) );
  XOR2_X1 U1492 (.Z( n1170 ) , .B( sa31_sr_0 ) , .A( w1_8 ) );
  XNOR2_X1 U1493 (.A( n1171 ) , .ZN( n732 ) , .B( n734 ) );
  XOR2_X1 U1494 (.Z( n1171 ) , .B( sa01_sr_0 ) , .A( w1_16 ) );
  XNOR2_X1 U1495 (.B( n1172 ) , .ZN( n853 ) , .A( n854 ) );
  XNOR2_X1 U1496 (.ZN( n1172 ) , .A( n836 ) , .B( n856 ) );
  XNOR2_X1 U1497 (.A( n1173 ) , .ZN( n905 ) , .B( n907 ) );
  XOR2_X1 U1498 (.Z( n1173 ) , .B( sa02_sr_0 ) , .A( w2_16 ) );
  XNOR2_X1 U1499 (.A( n1174 ) , .ZN( n653 ) , .B( n655 ) );
  OAI21_X1 U15 (.B1( ld ) , .B2( n13 ) , .A( n14 ) , .ZN( n984 ) );
  NAND2_X1 U150 (.A2( ld ) , .ZN( n148 ) , .A1( text_in[73] ) );
  XOR2_X1 U1500 (.Z( n1174 ) , .B( sa11_sr_5 ) , .A( w1_29 ) );
  XNOR2_X1 U1501 (.B( n1175 ) , .ZN( n456 ) , .A( n457 ) );
  XNOR2_X1 U1502 (.ZN( n1175 ) , .B( n459 ) , .A( sa23_sr_1 ) );
  XNOR2_X1 U1503 (.B( n1176 ) , .ZN( n721 ) , .A( n722 ) );
  XNOR2_X1 U1504 (.ZN( n1176 ) , .B( n724 ) , .A( sa11_sr_1 ) );
  XNOR2_X1 U1505 (.A( n1177 ) , .ZN( n680 ) , .B( n682 ) );
  XNOR2_X1 U1506 (.ZN( n1177 ) , .B( n665 ) , .A( n685 ) );
  XNOR2_X1 U1507 (.B( n1178 ) , .ZN( n625 ) , .A( n626 ) );
  XNOR2_X1 U1508 (.ZN( n1178 ) , .B( n628 ) , .A( sa20_sr_2 ) );
  XNOR2_X1 U1509 (.B( n1179 ) , .ZN( n547 ) , .A( n548 ) );
  OAI21_X1 U151 (.B1( ld ) , .ZN( n1052 ) , .B2( n149 ) , .A( n150 ) );
  XNOR2_X1 U1510 (.ZN( n1179 ) , .B( n550 ) , .A( sa10_sr_1 ) );
  XNOR2_X1 U1511 (.B( n1180 ) , .ZN( n375 ) , .A( n376 ) );
  XNOR2_X1 U1512 (.ZN( n1180 ) , .B( n378 ) , .A( sa13_sr_0 ) );
  XNOR2_X1 U1513 (.B( n1181 ) , .ZN( n961 ) , .A( n962 ) );
  XNOR2_X1 U1514 (.ZN( n1181 ) , .B( n964 ) , .A( sa22_sr_4 ) );
  XNOR2_X1 U1515 (.B( n1182 ) , .ZN( n342 ) , .A( n343 ) );
  XNOR2_X1 U1516 (.ZN( n1182 ) , .B( n345 ) , .A( sa13_sr_5 ) );
  XNOR2_X1 U1517 (.A( n1183 ) , .ZN( n552 ) , .B( n554 ) );
  XNOR2_X1 U1518 (.ZN( n1183 ) , .B( n539 ) , .A( n556 ) );
  XNOR2_X1 U1519 (.A( n1184 ) , .ZN( n810 ) , .B( n812 ) );
  NAND2_X1 U152 (.A2( ld ) , .ZN( n150 ) , .A1( text_in[74] ) );
  XOR2_X1 U1520 (.Z( n1184 ) , .B( sa21_sr_0 ) , .A( w1_0 ) );
  XNOR2_X1 U1521 (.A( n1185 ) , .ZN( n726 ) , .B( n728 ) );
  XNOR2_X1 U1522 (.ZN( n1185 ) , .B( n713 ) , .A( n730 ) );
  XNOR2_X1 U1523 (.B( n1186 ) , .ZN( n951 ) , .A( n952 ) );
  XNOR2_X1 U1524 (.ZN( n1186 ) , .B( n954 ) , .A( sa22_sr_6 ) );
  XNOR2_X1 U1525 (.A( n1187 ) , .ZN( n804 ) , .B( n806 ) );
  XNOR2_X1 U1526 (.ZN( n1187 ) , .B( n791 ) , .A( n808 ) );
  XNOR2_X1 U1527 (.A( n1188 ) , .ZN( n630 ) , .B( n632 ) );
  XNOR2_X1 U1528 (.ZN( n1188 ) , .B( n617 ) , .A( n634 ) );
  XOR2_X1 U1529 (.B( n1189 ) , .Z( n693 ) , .A( sa11_sr_6 ) );
  OAI21_X1 U153 (.B1( ld ) , .ZN( n1053 ) , .B2( n151 ) , .A( n152 ) );
  XNOR2_X1 U1530 (.ZN( n1189 ) , .B( sa21_sr_6 ) , .A( w1_23 ) );
  XNOR2_X1 U1531 (.A( n1190 ) , .ZN( n419 ) , .B( n421 ) );
  XOR2_X1 U1532 (.Z( n1190 ) , .B( sa33_sr_0 ) , .A( w3_8 ) );
  XNOR2_X1 U1533 (.A( n1191 ) , .ZN( n466 ) , .B( n468 ) );
  XNOR2_X1 U1534 (.ZN( n1191 ) , .B( n471 ) , .A( w0_31 ) );
  XNOR2_X1 U1535 (.A( n1192 ) , .ZN( n513 ) , .B( n515 ) );
  XOR2_X1 U1536 (.Z( n1192 ) , .B( sa10_sr_0 ) , .A( w0_24 ) );
  XNOR2_X1 U1537 (.A( n1193 ) , .ZN( n332 ) , .B( n334 ) );
  XOR2_X1 U1538 (.Z( n1193 ) , .B( sa13_sr_0 ) , .A( w3_24 ) );
  XNOR2_X1 U1539 (.A( n1194 ) , .ZN( n593 ) , .B( n595 ) );
  NAND2_X1 U154 (.A2( ld ) , .ZN( n152 ) , .A1( text_in[75] ) );
  XOR2_X1 U1540 (.Z( n1194 ) , .B( sa30_sr_0 ) , .A( w0_8 ) );
  XNOR2_X1 U1541 (.A( n1195 ) , .ZN( n286 ) , .B( n288 ) );
  XOR2_X1 U1542 (.Z( n1195 ) , .B( sa13_sr_7 ) , .A( w3_31 ) );
  XNOR2_X1 U1543 (.A( n1196 ) , .ZN( n584 ) , .B( n586 ) );
  XOR2_X1 U1544 (.Z( n1196 ) , .B( sa30_sr_2 ) , .A( w0_10 ) );
  XNOR2_X1 U1545 (.A( n1197 ) , .ZN( n674 ) , .B( n676 ) );
  XOR2_X1 U1546 (.Z( n1197 ) , .B( sa11_sr_2 ) , .A( w1_26 ) );
  XNOR2_X1 U1547 (.A( n1198 ) , .ZN( n758 ) , .B( n760 ) );
  XOR2_X1 U1548 (.Z( n1198 ) , .B( sa31_sr_2 ) , .A( w1_10 ) );
  XNOR2_X1 U1549 (.A( n1199 ) , .ZN( n298 ) , .B( n300 ) );
  OAI21_X1 U155 (.B1( ld ) , .ZN( n1054 ) , .B2( n153 ) , .A( n154 ) );
  XOR2_X1 U1550 (.Z( n1199 ) , .B( sa13_sr_5 ) , .A( w3_29 ) );
  XNOR2_X1 U1551 (.A( n1200 ) , .ZN( n319 ) , .B( n321 ) );
  XOR2_X1 U1552 (.Z( n1200 ) , .B( sa13_sr_2 ) , .A( w3_26 ) );
  XNOR2_X1 U1553 (.A( n1201 ) , .ZN( n410 ) , .B( n412 ) );
  XOR2_X1 U1554 (.Z( n1201 ) , .B( sa33_sr_2 ) , .A( w3_10 ) );
  XNOR2_X1 U1555 (.A( n1202 ) , .ZN( n462 ) , .B( n464 ) );
  XOR2_X1 U1556 (.Z( n1202 ) , .B( sa23_sr_0 ) , .A( w3_0 ) );
  XNOR2_X1 U1557 (.A( n1203 ) , .ZN( n558 ) , .B( n560 ) );
  XOR2_X1 U1558 (.Z( n1203 ) , .B( sa00_sr_0 ) , .A( w0_16 ) );
  XNOR2_X1 U1559 (.A( n1204 ) , .ZN( n636 ) , .B( n638 ) );
  NAND2_X1 U156 (.A2( ld ) , .ZN( n154 ) , .A1( text_in[76] ) );
  XOR2_X1 U1560 (.Z( n1204 ) , .B( sa20_sr_0 ) , .A( w0_0 ) );
  XNOR2_X1 U1561 (.A( n1205 ) , .ZN( n292 ) , .B( n294 ) );
  XOR2_X1 U1562 (.Z( n1205 ) , .B( sa13_sr_6 ) , .A( w3_30 ) );
  XNOR2_X1 U1563 (.ZN( N415 ) , .B( n1206 ) , .A( w0_18 ) );
  XNOR2_X1 U1564 (.ZN( N463 ) , .B( n1208 ) , .A( w2_10 ) );
  BUF_X1 U1565 (.A( n1109 ) , .Z( n1213 ) );
  XNOR2_X1 U1566 (.ZN( N423 ) , .B( n1207 ) , .A( w1_18 ) );
  INV_X1 U1567 (.ZN( n1206 ) , .A( sa10_sr_2 ) );
  INV_X1 U1568 (.ZN( n1207 ) , .A( sa11_sr_2 ) );
  NAND2_X1 U1569 (.A2( n1209 ) , .ZN( n1210 ) , .A1( sa22_sr_2 ) );
  OAI21_X1 U157 (.B1( ld ) , .ZN( n1055 ) , .B2( n155 ) , .A( n156 ) );
  NAND2_X1 U1570 (.A1( n1208 ) , .ZN( n1211 ) , .A2( sa32_sr_2 ) );
  NAND2_X1 U1571 (.A1( n1210 ) , .A2( n1211 ) , .ZN( n851 ) );
  INV_X1 U1572 (.ZN( n1208 ) , .A( sa22_sr_2 ) );
  INV_X1 U1573 (.ZN( n1209 ) , .A( sa32_sr_2 ) );
  INV_X1 U1574 (.ZN( n1215 ) , .A( n1221 ) );
  INV_X1 U1575 (.ZN( n1216 ) , .A( n1221 ) );
  INV_X1 U1576 (.A( ld ) , .ZN( n1222 ) );
  NAND2_X1 U158 (.A2( ld ) , .ZN( n156 ) , .A1( text_in[77] ) );
  OAI21_X1 U159 (.B1( ld ) , .ZN( n1056 ) , .B2( n157 ) , .A( n158 ) );
  NAND2_X1 U16 (.A2( ld ) , .ZN( n14 ) , .A1( text_in[6] ) );
  NAND2_X1 U160 (.A2( ld ) , .ZN( n158 ) , .A1( text_in[78] ) );
  OAI21_X1 U161 (.B1( ld ) , .ZN( n1057 ) , .B2( n159 ) , .A( n160 ) );
  NAND2_X1 U162 (.A2( ld ) , .ZN( n160 ) , .A1( text_in[79] ) );
  OAI21_X1 U163 (.B1( ld ) , .ZN( n1058 ) , .B2( n161 ) , .A( n162 ) );
  NAND2_X1 U164 (.A2( ld ) , .ZN( n162 ) , .A1( text_in[80] ) );
  OAI21_X1 U165 (.B1( ld ) , .ZN( n1059 ) , .B2( n163 ) , .A( n164 ) );
  NAND2_X1 U166 (.A2( ld ) , .ZN( n164 ) , .A1( text_in[81] ) );
  OAI21_X1 U167 (.B1( ld ) , .ZN( n1060 ) , .B2( n165 ) , .A( n166 ) );
  NAND2_X1 U168 (.A2( ld ) , .ZN( n166 ) , .A1( text_in[82] ) );
  OAI21_X1 U169 (.B1( ld ) , .ZN( n1061 ) , .B2( n167 ) , .A( n168 ) );
  OAI21_X1 U17 (.B1( ld ) , .B2( n15 ) , .A( n16 ) , .ZN( n985 ) );
  NAND2_X1 U170 (.A2( ld ) , .ZN( n168 ) , .A1( text_in[83] ) );
  OAI21_X1 U171 (.B1( ld ) , .ZN( n1062 ) , .B2( n169 ) , .A( n170 ) );
  NAND2_X1 U172 (.A2( ld ) , .ZN( n170 ) , .A1( text_in[84] ) );
  OAI21_X1 U173 (.B1( ld ) , .ZN( n1063 ) , .B2( n171 ) , .A( n172 ) );
  NAND2_X1 U174 (.A2( ld ) , .ZN( n172 ) , .A1( text_in[85] ) );
  OAI21_X1 U175 (.B1( ld ) , .ZN( n1064 ) , .B2( n173 ) , .A( n174 ) );
  NAND2_X1 U176 (.A2( ld ) , .ZN( n174 ) , .A1( text_in[86] ) );
  OAI21_X1 U177 (.B1( ld ) , .ZN( n1065 ) , .B2( n175 ) , .A( n176 ) );
  NAND2_X1 U178 (.A2( ld ) , .ZN( n176 ) , .A1( text_in[87] ) );
  OAI21_X1 U179 (.B1( ld ) , .ZN( n1066 ) , .B2( n177 ) , .A( n178 ) );
  NAND2_X1 U18 (.A2( ld ) , .ZN( n16 ) , .A1( text_in[7] ) );
  NAND2_X1 U180 (.A2( ld ) , .ZN( n178 ) , .A1( text_in[88] ) );
  OAI21_X1 U181 (.B1( ld ) , .ZN( n1067 ) , .B2( n179 ) , .A( n180 ) );
  NAND2_X1 U182 (.A2( ld ) , .ZN( n180 ) , .A1( text_in[89] ) );
  OAI21_X1 U183 (.B1( ld ) , .ZN( n1068 ) , .B2( n181 ) , .A( n182 ) );
  NAND2_X1 U184 (.A2( ld ) , .ZN( n182 ) , .A1( text_in[90] ) );
  OAI21_X1 U185 (.B1( ld ) , .ZN( n1069 ) , .B2( n183 ) , .A( n184 ) );
  NAND2_X1 U186 (.A2( ld ) , .ZN( n184 ) , .A1( text_in[91] ) );
  OAI21_X1 U187 (.B1( ld ) , .ZN( n1070 ) , .B2( n185 ) , .A( n186 ) );
  NAND2_X1 U188 (.A2( ld ) , .ZN( n186 ) , .A1( text_in[92] ) );
  OAI21_X1 U189 (.B1( ld ) , .ZN( n1071 ) , .B2( n187 ) , .A( n188 ) );
  OAI21_X1 U19 (.B1( ld ) , .B2( n17 ) , .A( n18 ) , .ZN( n986 ) );
  NAND2_X1 U190 (.A2( ld ) , .ZN( n188 ) , .A1( text_in[93] ) );
  OAI21_X1 U191 (.B1( ld ) , .ZN( n1072 ) , .B2( n189 ) , .A( n190 ) );
  NAND2_X1 U192 (.A2( ld ) , .ZN( n190 ) , .A1( text_in[94] ) );
  OAI21_X1 U193 (.B1( ld ) , .ZN( n1073 ) , .B2( n191 ) , .A( n192 ) );
  NAND2_X1 U194 (.A2( ld ) , .ZN( n192 ) , .A1( text_in[95] ) );
  OAI21_X1 U195 (.B1( ld ) , .ZN( n1074 ) , .B2( n193 ) , .A( n194 ) );
  NAND2_X1 U196 (.A2( ld ) , .ZN( n194 ) , .A1( text_in[96] ) );
  OAI21_X1 U197 (.B1( ld ) , .ZN( n1075 ) , .B2( n195 ) , .A( n196 ) );
  NAND2_X1 U198 (.A2( ld ) , .ZN( n196 ) , .A1( text_in[97] ) );
  OAI21_X1 U199 (.B1( ld ) , .ZN( n1076 ) , .B2( n197 ) , .A( n198 ) );
  NAND2_X1 U20 (.A2( ld ) , .ZN( n18 ) , .A1( text_in[8] ) );
  NAND2_X1 U200 (.A2( ld ) , .ZN( n198 ) , .A1( text_in[98] ) );
  OAI21_X1 U201 (.B1( ld ) , .ZN( n1077 ) , .B2( n199 ) , .A( n200 ) );
  NAND2_X1 U202 (.A2( ld ) , .ZN( n200 ) , .A1( text_in[99] ) );
  OAI21_X1 U203 (.B1( ld ) , .ZN( n1078 ) , .B2( n201 ) , .A( n202 ) );
  NAND2_X1 U204 (.A2( ld ) , .ZN( n202 ) , .A1( text_in[100] ) );
  OAI21_X1 U205 (.B1( ld ) , .ZN( n1079 ) , .B2( n203 ) , .A( n204 ) );
  NAND2_X1 U206 (.A2( ld ) , .ZN( n204 ) , .A1( text_in[101] ) );
  OAI21_X1 U207 (.B1( ld ) , .ZN( n1080 ) , .B2( n205 ) , .A( n206 ) );
  NAND2_X1 U208 (.A2( ld ) , .ZN( n206 ) , .A1( text_in[102] ) );
  OAI21_X1 U209 (.B1( ld ) , .ZN( n1081 ) , .B2( n207 ) , .A( n208 ) );
  OAI21_X1 U21 (.B1( ld ) , .B2( n19 ) , .A( n20 ) , .ZN( n987 ) );
  NAND2_X1 U210 (.A2( ld ) , .ZN( n208 ) , .A1( text_in[103] ) );
  OAI21_X1 U211 (.B1( ld ) , .ZN( n1082 ) , .B2( n209 ) , .A( n210 ) );
  NAND2_X1 U212 (.A2( ld ) , .ZN( n210 ) , .A1( text_in[104] ) );
  OAI21_X1 U213 (.B1( ld ) , .ZN( n1083 ) , .B2( n211 ) , .A( n212 ) );
  NAND2_X1 U214 (.A2( ld ) , .ZN( n212 ) , .A1( text_in[105] ) );
  OAI21_X1 U215 (.B1( ld ) , .ZN( n1084 ) , .B2( n213 ) , .A( n214 ) );
  NAND2_X1 U216 (.A2( ld ) , .ZN( n214 ) , .A1( text_in[106] ) );
  OAI21_X1 U217 (.B1( ld ) , .ZN( n1085 ) , .B2( n215 ) , .A( n216 ) );
  NAND2_X1 U218 (.A2( ld ) , .ZN( n216 ) , .A1( text_in[107] ) );
  OAI21_X1 U219 (.B1( ld ) , .ZN( n1086 ) , .B2( n217 ) , .A( n218 ) );
  NAND2_X1 U22 (.A2( ld ) , .ZN( n20 ) , .A1( text_in[9] ) );
  NAND2_X1 U220 (.A2( ld ) , .ZN( n218 ) , .A1( text_in[108] ) );
  OAI21_X1 U221 (.B1( ld ) , .ZN( n1087 ) , .B2( n219 ) , .A( n220 ) );
  NAND2_X1 U222 (.A2( ld ) , .ZN( n220 ) , .A1( text_in[109] ) );
  OAI21_X1 U223 (.B1( ld ) , .ZN( n1088 ) , .B2( n221 ) , .A( n222 ) );
  NAND2_X1 U224 (.A2( ld ) , .ZN( n222 ) , .A1( text_in[110] ) );
  OAI21_X1 U225 (.B1( ld ) , .ZN( n1089 ) , .B2( n223 ) , .A( n224 ) );
  NAND2_X1 U226 (.A2( ld ) , .ZN( n224 ) , .A1( text_in[111] ) );
  OAI21_X1 U227 (.B1( ld ) , .ZN( n1090 ) , .B2( n225 ) , .A( n226 ) );
  NAND2_X1 U228 (.A2( ld ) , .ZN( n226 ) , .A1( text_in[112] ) );
  OAI21_X1 U229 (.B1( ld ) , .ZN( n1091 ) , .B2( n227 ) , .A( n228 ) );
  OAI21_X1 U23 (.B1( ld ) , .B2( n21 ) , .A( n22 ) , .ZN( n988 ) );
  NAND2_X1 U230 (.A2( ld ) , .ZN( n228 ) , .A1( text_in[113] ) );
  OAI21_X1 U231 (.B1( ld ) , .ZN( n1092 ) , .B2( n229 ) , .A( n230 ) );
  NAND2_X1 U232 (.A2( ld ) , .ZN( n230 ) , .A1( text_in[114] ) );
  OAI21_X1 U233 (.B1( ld ) , .ZN( n1093 ) , .B2( n231 ) , .A( n232 ) );
  NAND2_X1 U234 (.A2( ld ) , .ZN( n232 ) , .A1( text_in[115] ) );
  OAI21_X1 U235 (.B1( ld ) , .ZN( n1094 ) , .B2( n233 ) , .A( n234 ) );
  NAND2_X1 U236 (.A2( ld ) , .ZN( n234 ) , .A1( text_in[116] ) );
  OAI21_X1 U237 (.B1( ld ) , .ZN( n1095 ) , .B2( n235 ) , .A( n236 ) );
  NAND2_X1 U238 (.A2( ld ) , .ZN( n236 ) , .A1( text_in[117] ) );
  OAI21_X1 U239 (.B1( ld ) , .ZN( n1096 ) , .B2( n237 ) , .A( n238 ) );
  NAND2_X1 U24 (.A2( ld ) , .ZN( n22 ) , .A1( text_in[10] ) );
  NAND2_X1 U240 (.A2( ld ) , .ZN( n238 ) , .A1( text_in[118] ) );
  OAI21_X1 U241 (.B1( ld ) , .ZN( n1097 ) , .B2( n239 ) , .A( n240 ) );
  NAND2_X1 U242 (.A2( ld ) , .ZN( n240 ) , .A1( text_in[119] ) );
  OAI21_X1 U243 (.B1( ld ) , .ZN( n1098 ) , .B2( n241 ) , .A( n242 ) );
  NAND2_X1 U244 (.A2( ld ) , .ZN( n242 ) , .A1( text_in[120] ) );
  OAI21_X1 U245 (.B1( ld ) , .ZN( n1099 ) , .B2( n243 ) , .A( n244 ) );
  NAND2_X1 U246 (.A2( ld ) , .ZN( n244 ) , .A1( text_in[121] ) );
  OAI21_X1 U247 (.B1( ld ) , .ZN( n1100 ) , .B2( n245 ) , .A( n246 ) );
  NAND2_X1 U248 (.A2( ld ) , .ZN( n246 ) , .A1( text_in[122] ) );
  OAI21_X1 U249 (.B1( ld ) , .ZN( n1101 ) , .B2( n247 ) , .A( n248 ) );
  OAI21_X1 U25 (.B1( ld ) , .B2( n23 ) , .A( n24 ) , .ZN( n989 ) );
  NAND2_X1 U250 (.A2( ld ) , .ZN( n248 ) , .A1( text_in[123] ) );
  OAI21_X1 U251 (.B1( ld ) , .ZN( n1102 ) , .B2( n249 ) , .A( n250 ) );
  NAND2_X1 U252 (.A2( ld ) , .ZN( n250 ) , .A1( text_in[124] ) );
  OAI21_X1 U253 (.B1( ld ) , .ZN( n1103 ) , .B2( n251 ) , .A( n252 ) );
  NAND2_X1 U254 (.A2( ld ) , .ZN( n252 ) , .A1( text_in[125] ) );
  OAI21_X1 U255 (.B1( ld ) , .ZN( n1104 ) , .B2( n253 ) , .A( n254 ) );
  NAND2_X1 U256 (.A2( ld ) , .ZN( n254 ) , .A1( text_in[126] ) );
  OAI21_X1 U257 (.B1( ld ) , .ZN( n1105 ) , .B2( n255 ) , .A( n256 ) );
  NAND2_X1 U258 (.A2( ld ) , .ZN( n256 ) , .A1( text_in[127] ) );
  AOI21_X1 U259 (.ZN( n1110 ) , .B1( n1222 ) , .B2( n258 ) , .A( n259 ) );
  NAND2_X1 U26 (.A2( ld ) , .ZN( n24 ) , .A1( text_in[11] ) );
  OAI21_X1 U260 (.ZN( n258 ) , .B1( n260 ) , .B2( n261 ) , .A( n262 ) );
  NOR3_X1 U261 (.A2( ld ) , .ZN( n1111 ) , .A1( n259 ) , .A3( n263 ) );
  AOI22_X1 U262 (.ZN( n263 ) , .A1( n264 ) , .A2( n265 ) , .B1( n266 ) , .B2( n267 ) );
  NOR2_X1 U263 (.A1( n1106 ) , .ZN( n264 ) , .A2( n267 ) );
  INV_X1 U265 (.ZN( n1112 ) , .A( n268 ) );
  OAI21_X1 U266 (.B1( ld ) , .ZN( n268 ) , .B2( n269 ) , .A( rst ) );
  AOI21_X1 U267 (.A( n1106 ) , .B1( n1107 ) , .B2( n265 ) , .ZN( n269 ) );
  INV_X1 U268 (.ZN( n265 ) , .A( n266 ) );
  NAND2_X1 U269 (.A1( n1108 ) , .A2( n262 ) , .ZN( n266 ) );
  OAI21_X1 U27 (.B1( ld ) , .B2( n25 ) , .A( n26 ) , .ZN( n990 ) );
  XNOR2_X1 U270 (.B( n261 ) , .ZN( n262 ) , .A( n977 ) );
  AOI21_X1 U272 (.ZN( n1113 ) , .B1( n1222 ) , .A( n259 ) , .B2( n270 ) );
  INV_X1 U273 (.ZN( n259 ) , .A( rst ) );
  OAI21_X1 U274 (.A( n1108 ) , .B2( n260 ) , .ZN( n270 ) , .B1( n977 ) );
  OAI22_X1 U276 (.ZN( N99 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n271 ) , .B1( n272 ) );
  XOR2_X1 U278 (.Z( n275 ) , .B( n276 ) , .A( sa22_sr_1 ) );
  XOR2_X1 U279 (.Z( n276 ) , .B( sa32_sr_0 ) , .A( w2_1 ) );
  NAND2_X1 U28 (.A2( ld ) , .ZN( n26 ) , .A1( text_in[12] ) );
  XOR2_X1 U281 (.Z( n278 ) , .B( n279 ) , .A( sa02_sr_0 ) );
  XOR2_X1 U282 (.Z( n271 ) , .A( n67 ) , .B( w2_1 ) );
  OAI22_X1 U284 (.ZN( N98 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n280 ) , .B1( n281 ) );
  XOR2_X1 U286 (.A( n279 ) , .Z( n283 ) , .B( n284 ) );
  XOR2_X1 U288 (.Z( n280 ) , .A( n65 ) , .B( w2_0 ) );
  OAI21_X1 U29 (.B1( ld ) , .B2( n27 ) , .A( n28 ) , .ZN( n991 ) );
  OAI22_X1 U290 (.ZN( N89 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n285 ) , .B1( n286 ) );
  XOR2_X1 U292 (.Z( n288 ) , .A( n289 ) , .B( n290 ) );
  XOR2_X1 U294 (.Z( n285 ) , .A( n63 ) , .B( w3_31 ) );
  OAI22_X1 U296 (.ZN( N88 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n291 ) , .B1( n292 ) );
  XOR2_X1 U298 (.Z( n294 ) , .A( n295 ) , .B( n296 ) );
  OAI21_X1 U3 (.B1( ld ) , .B2( n1 ) , .A( n2 ) , .ZN( n978 ) );
  NAND2_X1 U30 (.A2( ld ) , .ZN( n28 ) , .A1( text_in[13] ) );
  XOR2_X1 U300 (.Z( n291 ) , .A( n61 ) , .B( w3_30 ) );
  OAI22_X1 U302 (.ZN( N87 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n297 ) , .B1( n298 ) );
  XOR2_X1 U304 (.Z( n300 ) , .A( n301 ) , .B( n302 ) );
  XOR2_X1 U306 (.Z( n297 ) , .A( n59 ) , .B( w3_29 ) );
  OAI22_X1 U308 (.ZN( N86 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n303 ) , .B1( n304 ) );
  XOR2_X1 U309 (.Z( n304 ) , .A( n305 ) , .B( n306 ) );
  OAI21_X1 U31 (.B1( ld ) , .B2( n29 ) , .A( n30 ) , .ZN( n992 ) );
  XOR2_X1 U310 (.Z( n306 ) , .A( n307 ) , .B( n308 ) );
  XOR2_X1 U311 (.Z( n305 ) , .A( n309 ) , .B( n310 ) );
  XNOR2_X1 U312 (.ZN( n309 ) , .B( sa13_sr_4 ) , .A( w3_28 ) );
  XOR2_X1 U313 (.Z( n303 ) , .A( n57 ) , .B( w3_28 ) );
  OAI22_X1 U315 (.ZN( N85 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n311 ) , .B1( n312 ) );
  XOR2_X1 U317 (.Z( n314 ) , .A( n315 ) , .B( n316 ) );
  XNOR2_X1 U319 (.ZN( n317 ) , .B( sa13_sr_3 ) , .A( w3_27 ) );
  NAND2_X1 U32 (.A2( ld ) , .ZN( n30 ) , .A1( text_in[14] ) );
  XOR2_X1 U320 (.Z( n311 ) , .A( n55 ) , .B( w3_27 ) );
  OAI22_X1 U322 (.ZN( N84 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n318 ) , .B1( n319 ) );
  XOR2_X1 U324 (.Z( n321 ) , .A( n322 ) , .B( n323 ) );
  XOR2_X1 U326 (.Z( n318 ) , .A( n53 ) , .B( w3_26 ) );
  OAI22_X1 U328 (.ZN( N83 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n324 ) , .B1( n325 ) );
  OAI21_X1 U33 (.B1( ld ) , .B2( n31 ) , .A( n32 ) , .ZN( n993 ) );
  XOR2_X1 U330 (.Z( n327 ) , .A( n328 ) , .B( n329 ) );
  XNOR2_X1 U332 (.ZN( n330 ) , .B( sa13_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U333 (.Z( n324 ) , .A( n51 ) , .B( w3_25 ) );
  OAI22_X1 U335 (.ZN( N82 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n331 ) , .B1( n332 ) );
  XOR2_X1 U337 (.A( n307 ) , .Z( n334 ) , .B( n335 ) );
  XOR2_X1 U339 (.Z( n331 ) , .A( n49 ) , .B( w3_24 ) );
  NAND2_X1 U34 (.A2( ld ) , .ZN( n32 ) , .A1( text_in[15] ) );
  OAI22_X1 U341 (.ZN( N73 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n336 ) , .B1( n337 ) );
  XOR2_X1 U342 (.Z( n337 ) , .A( n338 ) , .B( n339 ) );
  XOR2_X1 U343 (.B( n289 ) , .Z( n339 ) , .A( sa03_sr_7 ) );
  XOR2_X1 U346 (.Z( n336 ) , .A( n47 ) , .B( w3_23 ) );
  OAI22_X1 U348 (.ZN( N72 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n341 ) , .B1( n342 ) );
  OAI21_X1 U35 (.B1( ld ) , .B2( n33 ) , .A( n34 ) , .ZN( n994 ) );
  XOR2_X1 U351 (.Z( n345 ) , .B( sa23_sr_5 ) , .A( w3_22 ) );
  XOR2_X1 U354 (.Z( n341 ) , .A( n45 ) , .B( w3_22 ) );
  OAI22_X1 U356 (.ZN( N71 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n347 ) , .B1( n348 ) );
  XOR2_X1 U357 (.Z( n348 ) , .A( n349 ) , .B( n350 ) );
  XOR2_X1 U358 (.Z( n350 ) , .B( n351 ) , .A( sa13_sr_4 ) );
  XOR2_X1 U359 (.Z( n351 ) , .B( sa23_sr_4 ) , .A( w3_21 ) );
  NAND2_X1 U36 (.A2( ld ) , .ZN( n34 ) , .A1( text_in[16] ) );
  XOR2_X1 U360 (.B( n301 ) , .Z( n349 ) , .A( n352 ) );
  XOR2_X1 U361 (.Z( n347 ) , .A( n43 ) , .B( w3_21 ) );
  OAI22_X1 U363 (.ZN( N70 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n353 ) , .B1( n354 ) );
  XOR2_X1 U364 (.Z( n354 ) , .A( n355 ) , .B( n356 ) );
  XOR2_X1 U365 (.Z( n356 ) , .B( n357 ) , .A( sa13_sr_3 ) );
  XOR2_X1 U366 (.Z( n357 ) , .B( sa23_sr_3 ) , .A( w3_20 ) );
  XOR2_X1 U367 (.Z( n355 ) , .A( n358 ) , .B( n359 ) );
  XOR2_X1 U368 (.B( n310 ) , .Z( n358 ) , .A( n360 ) );
  XOR2_X1 U369 (.Z( n353 ) , .A( n41 ) , .B( w3_20 ) );
  OAI21_X1 U37 (.B1( ld ) , .B2( n35 ) , .A( n36 ) , .ZN( n995 ) );
  OAI22_X1 U371 (.ZN( N69 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n361 ) , .B1( n362 ) );
  XOR2_X1 U374 (.Z( n365 ) , .B( sa23_sr_2 ) , .A( w3_19 ) );
  XOR2_X1 U375 (.B( n359 ) , .Z( n363 ) , .A( n366 ) );
  XOR2_X1 U376 (.B( n315 ) , .Z( n366 ) , .A( n367 ) );
  XOR2_X1 U377 (.Z( n361 ) , .A( n39 ) , .B( w3_19 ) );
  OAI22_X1 U379 (.ZN( N68 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n368 ) , .B1( n369 ) );
  NAND2_X1 U38 (.A2( ld ) , .ZN( n36 ) , .A1( text_in[17] ) );
  XOR2_X1 U382 (.Z( n372 ) , .B( sa23_sr_1 ) , .A( w3_18 ) );
  XOR2_X1 U383 (.B( n322 ) , .Z( n370 ) , .A( n373 ) );
  XOR2_X1 U384 (.Z( n368 ) , .A( n37 ) , .B( w3_18 ) );
  OAI22_X1 U386 (.ZN( N67 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n374 ) , .B1( n375 ) );
  XOR2_X1 U389 (.Z( n378 ) , .B( sa23_sr_0 ) , .A( w3_17 ) );
  OAI21_X1 U39 (.B1( ld ) , .B2( n37 ) , .A( n38 ) , .ZN( n996 ) );
  XOR2_X1 U390 (.B( n359 ) , .Z( n376 ) , .A( n379 ) );
  XOR2_X1 U391 (.B( n328 ) , .Z( n379 ) , .A( n380 ) );
  XOR2_X1 U392 (.A( n35 ) , .Z( n374 ) , .B( w3_17 ) );
  OAI22_X1 U394 (.ZN( N66 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n381 ) , .B1( n382 ) );
  XOR2_X1 U396 (.A( n335 ) , .B( n359 ) , .Z( n384 ) );
  XNOR2_X1 U397 (.ZN( n359 ) , .B( n385 ) , .A( sa13_sr_7 ) );
  XOR2_X1 U399 (.A( n33 ) , .Z( n381 ) , .B( w3_16 ) );
  NAND2_X1 U4 (.A2( ld ) , .ZN( n2 ) , .A1( text_in[0] ) );
  NAND2_X1 U40 (.A2( ld ) , .ZN( n38 ) , .A1( text_in[18] ) );
  OAI22_X1 U401 (.ZN( N57 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n387 ) , .B1( n388 ) );
  XOR2_X1 U403 (.A( n295 ) , .B( n307 ) , .Z( n390 ) );
  XOR2_X1 U404 (.Z( n295 ) , .A( sa23_sr_6 ) , .B( sa33_sr_6 ) );
  XOR2_X1 U406 (.A( n31 ) , .Z( n387 ) , .B( w3_15 ) );
  OAI22_X1 U408 (.ZN( N56 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n391 ) , .B1( n392 ) );
  OAI21_X1 U41 (.B1( ld ) , .B2( n39 ) , .A( n40 ) , .ZN( n997 ) );
  XOR2_X1 U410 (.A( n290 ) , .B( n301 ) , .Z( n394 ) );
  XOR2_X1 U411 (.Z( n301 ) , .A( sa23_sr_5 ) , .B( sa33_sr_5 ) );
  XOR2_X1 U413 (.A( n29 ) , .Z( n391 ) , .B( w3_14 ) );
  OAI22_X1 U415 (.ZN( N55 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n395 ) , .B1( n396 ) );
  XOR2_X1 U417 (.A( n296 ) , .B( n310 ) , .Z( n398 ) );
  XOR2_X1 U418 (.Z( n310 ) , .A( sa23_sr_4 ) , .B( sa33_sr_4 ) );
  NAND2_X1 U42 (.A2( ld ) , .ZN( n40 ) , .A1( text_in[19] ) );
  XOR2_X1 U420 (.A( n27 ) , .Z( n395 ) , .B( w3_13 ) );
  OAI22_X1 U422 (.ZN( N54 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n399 ) , .B1( n400 ) );
  XOR2_X1 U423 (.Z( n400 ) , .A( n401 ) , .B( n402 ) );
  XOR2_X1 U424 (.A( n302 ) , .B( n315 ) , .Z( n402 ) );
  XOR2_X1 U425 (.Z( n315 ) , .A( sa23_sr_3 ) , .B( sa33_sr_3 ) );
  XOR2_X1 U426 (.B( n289 ) , .Z( n401 ) , .A( n403 ) );
  XNOR2_X1 U427 (.ZN( n403 ) , .B( sa33_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U428 (.A( n25 ) , .Z( n399 ) , .B( w3_12 ) );
  OAI21_X1 U43 (.B1( ld ) , .B2( n41 ) , .A( n42 ) , .ZN( n998 ) );
  OAI22_X1 U430 (.ZN( N53 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n404 ) , .B1( n405 ) );
  XOR2_X1 U432 (.A( n308 ) , .B( n322 ) , .Z( n407 ) );
  XOR2_X1 U433 (.Z( n322 ) , .A( sa23_sr_2 ) , .B( sa33_sr_2 ) );
  XNOR2_X1 U435 (.ZN( n408 ) , .B( sa33_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U436 (.A( n23 ) , .Z( n404 ) , .B( w3_11 ) );
  OAI22_X1 U438 (.ZN( N52 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n409 ) , .B1( n410 ) );
  NAND2_X1 U44 (.A2( ld ) , .ZN( n42 ) , .A1( text_in[20] ) );
  XOR2_X1 U440 (.A( n316 ) , .B( n328 ) , .Z( n412 ) );
  XOR2_X1 U441 (.Z( n328 ) , .A( sa23_sr_1 ) , .B( sa33_sr_1 ) );
  XOR2_X1 U443 (.A( n21 ) , .Z( n409 ) , .B( w3_10 ) );
  OAI22_X1 U445 (.ZN( N51 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n413 ) , .B1( n414 ) );
  XOR2_X1 U447 (.A( n323 ) , .B( n335 ) , .Z( n416 ) );
  XOR2_X1 U448 (.Z( n335 ) , .A( sa23_sr_0 ) , .B( sa33_sr_0 ) );
  OAI21_X1 U45 (.B1( ld ) , .B2( n43 ) , .A( n44 ) , .ZN( n999 ) );
  XNOR2_X1 U450 (.ZN( n417 ) , .B( sa33_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U451 (.A( n19 ) , .Z( n413 ) , .B( w3_9 ) );
  XOR2_X1 U453 (.Z( N505 ) , .B( sa33_sr_0 ) , .A( w3_0 ) );
  XOR2_X1 U454 (.Z( N504 ) , .B( sa33_sr_1 ) , .A( w3_1 ) );
  XOR2_X1 U455 (.Z( N503 ) , .B( sa33_sr_2 ) , .A( w3_2 ) );
  XOR2_X1 U456 (.Z( N502 ) , .B( sa33_sr_3 ) , .A( w3_3 ) );
  XOR2_X1 U457 (.Z( N501 ) , .B( sa33_sr_4 ) , .A( w3_4 ) );
  XOR2_X1 U458 (.Z( N500 ) , .B( sa33_sr_5 ) , .A( w3_5 ) );
  OAI22_X1 U459 (.ZN( N50 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n418 ) , .B1( n419 ) );
  NAND2_X1 U46 (.A2( ld ) , .ZN( n44 ) , .A1( text_in[21] ) );
  XOR2_X1 U461 (.A( n289 ) , .B( n329 ) , .Z( n421 ) );
  XOR2_X1 U462 (.Z( n289 ) , .A( sa23_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U464 (.A( n17 ) , .Z( n418 ) , .B( w3_8 ) );
  XOR2_X1 U466 (.Z( N499 ) , .B( sa33_sr_6 ) , .A( w3_6 ) );
  XOR2_X1 U467 (.Z( N498 ) , .B( sa33_sr_7 ) , .A( w3_7 ) );
  XOR2_X1 U468 (.Z( N497 ) , .B( sa32_sr_0 ) , .A( w2_0 ) );
  XOR2_X1 U469 (.Z( N496 ) , .B( sa32_sr_1 ) , .A( w2_1 ) );
  OAI21_X1 U47 (.B1( ld ) , .ZN( n1000 ) , .B2( n45 ) , .A( n46 ) );
  XOR2_X1 U471 (.Z( N494 ) , .B( sa32_sr_3 ) , .A( w2_3 ) );
  XOR2_X1 U472 (.Z( N493 ) , .B( sa32_sr_4 ) , .A( w2_4 ) );
  XOR2_X1 U473 (.Z( N492 ) , .B( sa32_sr_5 ) , .A( w2_5 ) );
  XOR2_X1 U474 (.Z( N491 ) , .B( sa32_sr_6 ) , .A( w2_6 ) );
  XOR2_X1 U475 (.Z( N490 ) , .B( sa32_sr_7 ) , .A( w2_7 ) );
  XOR2_X1 U476 (.Z( N489 ) , .B( sa31_sr_0 ) , .A( w1_0 ) );
  XOR2_X1 U477 (.Z( N488 ) , .B( sa31_sr_1 ) , .A( w1_1 ) );
  XOR2_X1 U478 (.Z( N487 ) , .B( sa31_sr_2 ) , .A( w1_2 ) );
  XOR2_X1 U479 (.Z( N486 ) , .B( sa31_sr_3 ) , .A( w1_3 ) );
  NAND2_X1 U48 (.A2( ld ) , .ZN( n46 ) , .A1( text_in[22] ) );
  XOR2_X1 U480 (.Z( N485 ) , .B( sa31_sr_4 ) , .A( w1_4 ) );
  XOR2_X1 U481 (.Z( N484 ) , .B( sa31_sr_5 ) , .A( w1_5 ) );
  XOR2_X1 U482 (.Z( N483 ) , .B( sa31_sr_6 ) , .A( w1_6 ) );
  XOR2_X1 U483 (.Z( N482 ) , .B( sa31_sr_7 ) , .A( w1_7 ) );
  XOR2_X1 U484 (.Z( N481 ) , .B( sa30_sr_0 ) , .A( w0_0 ) );
  XOR2_X1 U485 (.Z( N480 ) , .B( sa30_sr_1 ) , .A( w0_1 ) );
  XOR2_X1 U486 (.Z( N479 ) , .B( sa30_sr_2 ) , .A( w0_2 ) );
  XOR2_X1 U487 (.Z( N478 ) , .B( sa30_sr_3 ) , .A( w0_3 ) );
  XOR2_X1 U488 (.Z( N477 ) , .B( sa30_sr_4 ) , .A( w0_4 ) );
  XOR2_X1 U489 (.Z( N476 ) , .B( sa30_sr_5 ) , .A( w0_5 ) );
  OAI21_X1 U49 (.B1( ld ) , .ZN( n1001 ) , .B2( n47 ) , .A( n48 ) );
  XOR2_X1 U490 (.Z( N475 ) , .B( sa30_sr_6 ) , .A( w0_6 ) );
  XOR2_X1 U491 (.Z( N474 ) , .B( sa30_sr_7 ) , .A( w0_7 ) );
  XOR2_X1 U492 (.Z( N473 ) , .B( sa23_sr_0 ) , .A( w3_8 ) );
  XOR2_X1 U493 (.Z( N472 ) , .B( sa23_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U494 (.Z( N471 ) , .B( sa23_sr_2 ) , .A( w3_10 ) );
  XOR2_X1 U495 (.Z( N470 ) , .B( sa23_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U496 (.Z( N469 ) , .B( sa23_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U497 (.Z( N468 ) , .B( sa23_sr_5 ) , .A( w3_13 ) );
  XOR2_X1 U498 (.Z( N467 ) , .B( sa23_sr_6 ) , .A( w3_14 ) );
  XOR2_X1 U499 (.Z( N466 ) , .B( sa23_sr_7 ) , .A( w3_15 ) );
  OAI21_X1 U5 (.B1( ld ) , .B2( n3 ) , .A( n4 ) , .ZN( n979 ) );
  NAND2_X1 U50 (.A2( ld ) , .ZN( n48 ) , .A1( text_in[23] ) );
  XOR2_X1 U500 (.Z( N465 ) , .B( sa22_sr_0 ) , .A( w2_8 ) );
  XOR2_X1 U501 (.Z( N464 ) , .B( sa22_sr_1 ) , .A( w2_9 ) );
  XOR2_X1 U503 (.Z( N462 ) , .B( sa22_sr_3 ) , .A( w2_11 ) );
  XOR2_X1 U504 (.Z( N461 ) , .B( sa22_sr_4 ) , .A( w2_12 ) );
  XOR2_X1 U505 (.Z( N460 ) , .B( sa22_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U506 (.Z( N459 ) , .B( sa22_sr_6 ) , .A( w2_14 ) );
  XOR2_X1 U507 (.Z( N458 ) , .B( sa22_sr_7 ) , .A( w2_15 ) );
  XOR2_X1 U508 (.Z( N457 ) , .B( sa21_sr_0 ) , .A( w1_8 ) );
  XOR2_X1 U509 (.Z( N456 ) , .B( sa21_sr_1 ) , .A( w1_9 ) );
  OAI21_X1 U51 (.B1( ld ) , .ZN( n1002 ) , .B2( n49 ) , .A( n50 ) );
  XOR2_X1 U510 (.Z( N455 ) , .B( sa21_sr_2 ) , .A( w1_10 ) );
  XOR2_X1 U511 (.Z( N454 ) , .B( sa21_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U512 (.Z( N453 ) , .B( sa21_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U513 (.Z( N452 ) , .B( sa21_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U514 (.Z( N451 ) , .B( sa21_sr_6 ) , .A( w1_14 ) );
  XOR2_X1 U515 (.Z( N450 ) , .B( sa21_sr_7 ) , .A( w1_15 ) );
  XOR2_X1 U516 (.Z( N449 ) , .B( sa20_sr_0 ) , .A( w0_8 ) );
  XOR2_X1 U517 (.Z( N448 ) , .B( sa20_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U518 (.Z( N447 ) , .B( sa20_sr_2 ) , .A( w0_10 ) );
  XOR2_X1 U519 (.Z( N446 ) , .B( sa20_sr_3 ) , .A( w0_11 ) );
  NAND2_X1 U52 (.A2( ld ) , .ZN( n50 ) , .A1( text_in[24] ) );
  XOR2_X1 U520 (.Z( N445 ) , .B( sa20_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U521 (.Z( N444 ) , .B( sa20_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U522 (.Z( N443 ) , .B( sa20_sr_6 ) , .A( w0_14 ) );
  XOR2_X1 U523 (.Z( N442 ) , .B( sa20_sr_7 ) , .A( w0_15 ) );
  XOR2_X1 U524 (.Z( N441 ) , .B( sa13_sr_0 ) , .A( w3_16 ) );
  XOR2_X1 U525 (.Z( N440 ) , .B( sa13_sr_1 ) , .A( w3_17 ) );
  XOR2_X1 U526 (.Z( N439 ) , .B( sa13_sr_2 ) , .A( w3_18 ) );
  XOR2_X1 U527 (.Z( N438 ) , .B( sa13_sr_3 ) , .A( w3_19 ) );
  XOR2_X1 U528 (.Z( N437 ) , .B( sa13_sr_4 ) , .A( w3_20 ) );
  XOR2_X1 U529 (.Z( N436 ) , .B( sa13_sr_5 ) , .A( w3_21 ) );
  OAI21_X1 U53 (.B1( ld ) , .ZN( n1003 ) , .B2( n51 ) , .A( n52 ) );
  XOR2_X1 U530 (.Z( N435 ) , .B( sa13_sr_6 ) , .A( w3_22 ) );
  XOR2_X1 U531 (.Z( N434 ) , .B( sa13_sr_7 ) , .A( w3_23 ) );
  XOR2_X1 U532 (.Z( N433 ) , .B( sa12_sr_0 ) , .A( w2_16 ) );
  XOR2_X1 U533 (.Z( N432 ) , .B( sa12_sr_1 ) , .A( w2_17 ) );
  XOR2_X1 U534 (.Z( N431 ) , .B( sa12_sr_2 ) , .A( w2_18 ) );
  XOR2_X1 U535 (.Z( N430 ) , .B( sa12_sr_3 ) , .A( w2_19 ) );
  XOR2_X1 U536 (.Z( N429 ) , .B( sa12_sr_4 ) , .A( w2_20 ) );
  XOR2_X1 U537 (.Z( N428 ) , .B( sa12_sr_5 ) , .A( w2_21 ) );
  XOR2_X1 U538 (.Z( N427 ) , .B( sa12_sr_6 ) , .A( w2_22 ) );
  XOR2_X1 U539 (.Z( N426 ) , .B( sa12_sr_7 ) , .A( w2_23 ) );
  NAND2_X1 U54 (.A2( ld ) , .ZN( n52 ) , .A1( text_in[25] ) );
  XOR2_X1 U540 (.Z( N425 ) , .B( sa11_sr_0 ) , .A( w1_16 ) );
  XOR2_X1 U541 (.Z( N424 ) , .B( sa11_sr_1 ) , .A( w1_17 ) );
  XOR2_X1 U543 (.Z( N422 ) , .B( sa11_sr_3 ) , .A( w1_19 ) );
  XOR2_X1 U544 (.Z( N421 ) , .B( sa11_sr_4 ) , .A( w1_20 ) );
  XOR2_X1 U545 (.Z( N420 ) , .B( sa11_sr_5 ) , .A( w1_21 ) );
  XOR2_X1 U546 (.Z( N419 ) , .B( sa11_sr_6 ) , .A( w1_22 ) );
  XOR2_X1 U547 (.Z( N418 ) , .B( sa11_sr_7 ) , .A( w1_23 ) );
  XOR2_X1 U548 (.Z( N417 ) , .B( sa10_sr_0 ) , .A( w0_16 ) );
  XOR2_X1 U549 (.Z( N416 ) , .B( sa10_sr_1 ) , .A( w0_17 ) );
  OAI21_X1 U55 (.B1( ld ) , .ZN( n1004 ) , .B2( n53 ) , .A( n54 ) );
  XOR2_X1 U551 (.Z( N414 ) , .B( sa10_sr_3 ) , .A( w0_19 ) );
  XOR2_X1 U552 (.Z( N413 ) , .B( sa10_sr_4 ) , .A( w0_20 ) );
  XOR2_X1 U553 (.Z( N412 ) , .B( sa10_sr_5 ) , .A( w0_21 ) );
  XOR2_X1 U554 (.Z( N411 ) , .B( sa10_sr_6 ) , .A( w0_22 ) );
  XOR2_X1 U555 (.Z( N410 ) , .B( sa10_sr_7 ) , .A( w0_23 ) );
  OAI22_X1 U556 (.ZN( N41 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n422 ) , .B1( n423 ) );
  XOR2_X1 U557 (.Z( n423 ) , .A( n424 ) , .B( n425 ) );
  XOR2_X1 U558 (.B( n307 ) , .Z( n425 ) , .A( sa03_sr_6 ) );
  XOR2_X1 U559 (.Z( n307 ) , .A( sa03_sr_7 ) , .B( sa13_sr_7 ) );
  NAND2_X1 U56 (.A2( ld ) , .ZN( n54 ) , .A1( text_in[26] ) );
  XOR2_X1 U560 (.A( n385 ) , .Z( n424 ) , .B( n426 ) );
  XOR2_X1 U561 (.Z( n426 ) , .B( sa33_sr_6 ) , .A( w3_7 ) );
  INV_X1 U562 (.ZN( n385 ) , .A( sa23_sr_7 ) );
  XOR2_X1 U563 (.A( n15 ) , .Z( n422 ) , .B( w3_7 ) );
  XOR2_X1 U565 (.Z( N409 ) , .B( sa03_sr_0 ) , .A( w3_24 ) );
  XOR2_X1 U566 (.Z( N408 ) , .B( sa03_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U567 (.Z( N407 ) , .B( sa03_sr_2 ) , .A( w3_26 ) );
  XOR2_X1 U568 (.Z( N406 ) , .B( sa03_sr_3 ) , .A( w3_27 ) );
  XOR2_X1 U569 (.Z( N405 ) , .B( sa03_sr_4 ) , .A( w3_28 ) );
  OAI21_X1 U57 (.B1( ld ) , .ZN( n1005 ) , .B2( n55 ) , .A( n56 ) );
  XOR2_X1 U570 (.Z( N404 ) , .B( sa03_sr_5 ) , .A( w3_29 ) );
  XOR2_X1 U571 (.Z( N403 ) , .B( sa03_sr_6 ) , .A( w3_30 ) );
  XOR2_X1 U572 (.Z( N402 ) , .B( sa03_sr_7 ) , .A( w3_31 ) );
  XOR2_X1 U573 (.Z( N401 ) , .B( sa02_sr_0 ) , .A( w2_24 ) );
  XOR2_X1 U574 (.Z( N400 ) , .B( sa02_sr_1 ) , .A( w2_25 ) );
  OAI22_X1 U575 (.ZN( N40 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n427 ) , .B1( n428 ) );
  XOR2_X1 U578 (.Z( n431 ) , .B( sa33_sr_5 ) , .A( w3_6 ) );
  XOR2_X1 U579 (.B( n290 ) , .A( n352 ) , .Z( n429 ) );
  NAND2_X1 U58 (.A2( ld ) , .ZN( n56 ) , .A1( text_in[27] ) );
  XOR2_X1 U580 (.Z( n290 ) , .A( sa03_sr_6 ) , .B( sa13_sr_6 ) );
  INV_X1 U581 (.ZN( n352 ) , .A( sa03_sr_5 ) );
  XOR2_X1 U582 (.A( n13 ) , .Z( n427 ) , .B( w3_6 ) );
  XOR2_X1 U584 (.Z( N399 ) , .B( sa02_sr_2 ) , .A( w2_26 ) );
  XOR2_X1 U585 (.Z( N398 ) , .B( sa02_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U586 (.Z( N397 ) , .B( sa02_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U587 (.Z( N396 ) , .B( sa02_sr_5 ) , .A( w2_29 ) );
  XOR2_X1 U588 (.Z( N395 ) , .B( sa02_sr_6 ) , .A( w2_30 ) );
  XOR2_X1 U589 (.Z( N394 ) , .B( sa02_sr_7 ) , .A( w2_31 ) );
  OAI21_X1 U59 (.B1( ld ) , .ZN( n1006 ) , .B2( n57 ) , .A( n58 ) );
  XOR2_X1 U590 (.Z( N393 ) , .B( sa01_sr_0 ) , .A( w1_24 ) );
  XOR2_X1 U591 (.Z( N392 ) , .B( sa01_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U592 (.Z( N391 ) , .B( sa01_sr_2 ) , .A( w1_26 ) );
  XOR2_X1 U593 (.Z( N390 ) , .B( sa01_sr_3 ) , .A( w1_27 ) );
  OAI22_X1 U594 (.ZN( N39 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n432 ) , .B1( n433 ) );
  XOR2_X1 U597 (.Z( n436 ) , .B( sa33_sr_4 ) , .A( w3_5 ) );
  XOR2_X1 U598 (.B( n296 ) , .A( n360 ) , .Z( n434 ) );
  XOR2_X1 U599 (.Z( n296 ) , .A( sa03_sr_5 ) , .B( sa13_sr_5 ) );
  NAND2_X1 U6 (.A2( ld ) , .ZN( n4 ) , .A1( text_in[1] ) );
  NAND2_X1 U60 (.A2( ld ) , .ZN( n58 ) , .A1( text_in[28] ) );
  INV_X1 U600 (.ZN( n360 ) , .A( sa03_sr_4 ) );
  XOR2_X1 U601 (.A( n11 ) , .Z( n432 ) , .B( w3_5 ) );
  XOR2_X1 U603 (.Z( N389 ) , .B( sa01_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U604 (.Z( N388 ) , .B( sa01_sr_5 ) , .A( w1_29 ) );
  XOR2_X1 U605 (.Z( N387 ) , .B( sa01_sr_6 ) , .A( w1_30 ) );
  XOR2_X1 U606 (.Z( N386 ) , .B( sa01_sr_7 ) , .A( w1_31 ) );
  XOR2_X1 U607 (.Z( N385 ) , .B( sa00_sr_0 ) , .A( w0_24 ) );
  XOR2_X1 U608 (.Z( N384 ) , .B( sa00_sr_1 ) , .A( w0_25 ) );
  XOR2_X1 U609 (.Z( N383 ) , .B( sa00_sr_2 ) , .A( w0_26 ) );
  OAI21_X1 U61 (.B1( ld ) , .ZN( n1007 ) , .B2( n59 ) , .A( n60 ) );
  XOR2_X1 U610 (.Z( N382 ) , .B( sa00_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U611 (.Z( N381 ) , .B( sa00_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U612 (.Z( N380 ) , .B( sa00_sr_5 ) , .A( w0_29 ) );
  OAI22_X1 U613 (.ZN( N38 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n437 ) , .B1( n438 ) );
  XOR2_X1 U614 (.Z( n438 ) , .A( n439 ) , .B( n440 ) );
  XOR2_X1 U615 (.Z( n440 ) , .B( n441 ) , .A( sa23_sr_4 ) );
  XOR2_X1 U616 (.Z( n441 ) , .B( sa33_sr_3 ) , .A( w3_4 ) );
  XOR2_X1 U617 (.Z( n439 ) , .A( n442 ) , .B( n443 ) );
  XOR2_X1 U618 (.B( n302 ) , .A( n367 ) , .Z( n442 ) );
  XOR2_X1 U619 (.Z( n302 ) , .A( sa03_sr_4 ) , .B( sa13_sr_4 ) );
  NAND2_X1 U62 (.A2( ld ) , .ZN( n60 ) , .A1( text_in[29] ) );
  INV_X1 U620 (.ZN( n367 ) , .A( sa03_sr_3 ) );
  XOR2_X1 U621 (.Z( n437 ) , .A( n9 ) , .B( w3_4 ) );
  XOR2_X1 U623 (.Z( N379 ) , .B( sa00_sr_6 ) , .A( w0_30 ) );
  XOR2_X1 U624 (.Z( N378 ) , .B( sa00_sr_7 ) , .A( w0_31 ) );
  OAI22_X1 U625 (.ZN( N37 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n444 ) , .B1( n445 ) );
  XOR2_X1 U628 (.Z( n448 ) , .B( sa33_sr_2 ) , .A( w3_3 ) );
  XOR2_X1 U629 (.B( n443 ) , .Z( n446 ) , .A( n449 ) );
  OAI21_X1 U63 (.B1( ld ) , .ZN( n1008 ) , .B2( n61 ) , .A( n62 ) );
  XOR2_X1 U630 (.B( n308 ) , .A( n373 ) , .Z( n449 ) );
  XOR2_X1 U631 (.Z( n308 ) , .A( sa03_sr_3 ) , .B( sa13_sr_3 ) );
  INV_X1 U632 (.ZN( n373 ) , .A( sa03_sr_2 ) );
  XOR2_X1 U633 (.Z( n444 ) , .A( n7 ) , .B( w3_3 ) );
  OAI22_X1 U635 (.ZN( N36 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n450 ) , .B1( n451 ) );
  XOR2_X1 U636 (.Z( n451 ) , .A( n452 ) , .B( n453 ) );
  XOR2_X1 U637 (.Z( n453 ) , .B( n454 ) , .A( sa23_sr_2 ) );
  XOR2_X1 U638 (.Z( n454 ) , .B( sa33_sr_1 ) , .A( w3_2 ) );
  XOR2_X1 U639 (.B( n316 ) , .A( n380 ) , .Z( n452 ) );
  NAND2_X1 U64 (.A2( ld ) , .ZN( n62 ) , .A1( text_in[30] ) );
  XOR2_X1 U640 (.Z( n316 ) , .A( sa03_sr_2 ) , .B( sa13_sr_2 ) );
  INV_X1 U641 (.ZN( n380 ) , .A( sa03_sr_1 ) );
  XOR2_X1 U642 (.Z( n450 ) , .A( n5 ) , .B( w3_2 ) );
  OAI22_X1 U644 (.ZN( N35 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n455 ) , .B1( n456 ) );
  XOR2_X1 U647 (.Z( n459 ) , .B( sa33_sr_0 ) , .A( w3_1 ) );
  XOR2_X1 U648 (.B( n443 ) , .Z( n457 ) , .A( n460 ) );
  XOR2_X1 U649 (.B( n323 ) , .A( n386 ) , .Z( n460 ) );
  OAI21_X1 U65 (.B1( ld ) , .ZN( n1009 ) , .B2( n63 ) , .A( n64 ) );
  XOR2_X1 U650 (.Z( n323 ) , .A( sa03_sr_1 ) , .B( sa13_sr_1 ) );
  INV_X1 U651 (.ZN( n386 ) , .A( sa03_sr_0 ) );
  XOR2_X1 U652 (.A( n3 ) , .Z( n455 ) , .B( w3_1 ) );
  OAI22_X1 U654 (.ZN( N34 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n461 ) , .B1( n462 ) );
  XOR2_X1 U656 (.A( n329 ) , .B( n443 ) , .Z( n464 ) );
  XOR2_X1 U657 (.Z( n443 ) , .A( sa03_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U658 (.Z( n329 ) , .A( sa03_sr_0 ) , .B( sa13_sr_0 ) );
  NAND2_X1 U66 (.A2( ld ) , .ZN( n64 ) , .A1( text_in[31] ) );
  XOR2_X1 U660 (.A( n1 ) , .Z( n461 ) , .B( w3_0 ) );
  OAI22_X1 U662 (.ZN( N281 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n465 ) , .B1( n466 ) );
  XOR2_X1 U664 (.Z( n468 ) , .A( n469 ) , .B( n470 ) );
  INV_X1 U666 (.ZN( n471 ) , .A( sa10_sr_7 ) );
  XOR2_X1 U667 (.A( n255 ) , .Z( n465 ) , .B( w0_31 ) );
  OAI22_X1 U669 (.ZN( N280 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n472 ) , .B1( n473 ) );
  OAI21_X1 U67 (.B1( ld ) , .ZN( n1010 ) , .B2( n65 ) , .A( n66 ) );
  XOR2_X1 U671 (.Z( n475 ) , .A( n476 ) , .B( n477 ) );
  XOR2_X1 U673 (.A( n253 ) , .Z( n472 ) , .B( w0_30 ) );
  OAI22_X1 U675 (.ZN( N279 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n478 ) , .B1( n479 ) );
  XOR2_X1 U677 (.Z( n481 ) , .A( n482 ) , .B( n483 ) );
  XOR2_X1 U679 (.A( n251 ) , .Z( n478 ) , .B( w0_29 ) );
  NAND2_X1 U68 (.A2( ld ) , .ZN( n66 ) , .A1( text_in[32] ) );
  OAI22_X1 U681 (.ZN( N278 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n484 ) , .B1( n485 ) );
  XOR2_X1 U682 (.Z( n485 ) , .A( n486 ) , .B( n487 ) );
  XOR2_X1 U683 (.Z( n487 ) , .A( n488 ) , .B( n489 ) );
  XOR2_X1 U684 (.Z( n486 ) , .A( n490 ) , .B( n491 ) );
  XNOR2_X1 U685 (.ZN( n490 ) , .B( sa10_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U686 (.A( n249 ) , .Z( n484 ) , .B( w0_28 ) );
  OAI22_X1 U688 (.ZN( N277 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n492 ) , .B1( n493 ) );
  OAI21_X1 U69 (.B1( ld ) , .ZN( n1011 ) , .B2( n67 ) , .A( n68 ) );
  XOR2_X1 U690 (.Z( n495 ) , .A( n496 ) , .B( n497 ) );
  XNOR2_X1 U692 (.ZN( n498 ) , .B( sa10_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U693 (.A( n247 ) , .Z( n492 ) , .B( w0_27 ) );
  OAI22_X1 U695 (.ZN( N276 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n499 ) , .B1( n500 ) );
  XOR2_X1 U697 (.Z( n502 ) , .A( n503 ) , .B( n504 ) );
  XOR2_X1 U699 (.A( n245 ) , .Z( n499 ) , .B( w0_26 ) );
  OAI21_X1 U7 (.B1( ld ) , .B2( n5 ) , .A( n6 ) , .ZN( n980 ) );
  NAND2_X1 U70 (.A2( ld ) , .ZN( n68 ) , .A1( text_in[33] ) );
  OAI22_X1 U701 (.ZN( N275 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n505 ) , .B1( n506 ) );
  XOR2_X1 U703 (.Z( n508 ) , .A( n509 ) , .B( n510 ) );
  XNOR2_X1 U705 (.ZN( n511 ) , .B( sa10_sr_1 ) , .A( w0_25 ) );
  XOR2_X1 U706 (.A( n243 ) , .Z( n505 ) , .B( w0_25 ) );
  OAI22_X1 U708 (.ZN( N274 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n512 ) , .B1( n513 ) );
  OAI21_X1 U71 (.B1( ld ) , .ZN( n1012 ) , .B2( n69 ) , .A( n70 ) );
  XOR2_X1 U710 (.A( n488 ) , .Z( n515 ) , .B( n516 ) );
  XOR2_X1 U712 (.A( n241 ) , .Z( n512 ) , .B( w0_24 ) );
  OAI22_X1 U714 (.ZN( N265 ) , .B2( n1114 ) , .A1( n1215 ) , .A2( n517 ) , .B1( n518 ) );
  XOR2_X1 U715 (.Z( n518 ) , .A( n519 ) , .B( n520 ) );
  XOR2_X1 U716 (.B( n469 ) , .Z( n520 ) , .A( sa00_sr_7 ) );
  XNOR2_X1 U717 (.ZN( n519 ) , .B( n521 ) , .A( sa10_sr_6 ) );
  XOR2_X1 U718 (.Z( n521 ) , .B( sa20_sr_6 ) , .A( w0_23 ) );
  XOR2_X1 U719 (.A( n239 ) , .Z( n517 ) , .B( w0_23 ) );
  NAND2_X1 U72 (.A2( ld ) , .ZN( n70 ) , .A1( text_in[34] ) );
  OAI22_X1 U721 (.ZN( N264 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n522 ) , .B1( n523 ) );
  XOR2_X1 U724 (.Z( n526 ) , .B( sa20_sr_5 ) , .A( w0_22 ) );
  XOR2_X1 U727 (.A( n237 ) , .Z( n522 ) , .B( w0_22 ) );
  OAI22_X1 U729 (.ZN( N263 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n528 ) , .B1( n529 ) );
  OAI21_X1 U73 (.B1( ld ) , .ZN( n1013 ) , .B2( n71 ) , .A( n72 ) );
  XOR2_X1 U730 (.Z( n529 ) , .A( n530 ) , .B( n531 ) );
  XOR2_X1 U731 (.Z( n531 ) , .B( n532 ) , .A( sa10_sr_4 ) );
  XOR2_X1 U732 (.Z( n532 ) , .B( sa20_sr_4 ) , .A( w0_21 ) );
  XNOR2_X1 U733 (.B( n482 ) , .ZN( n530 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U734 (.A( n235 ) , .Z( n528 ) , .B( w0_21 ) );
  OAI22_X1 U736 (.ZN( N262 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n533 ) , .B1( n534 ) );
  XOR2_X1 U737 (.Z( n534 ) , .A( n535 ) , .B( n536 ) );
  XOR2_X1 U738 (.Z( n536 ) , .B( n537 ) , .A( sa10_sr_3 ) );
  XOR2_X1 U739 (.Z( n537 ) , .B( sa20_sr_3 ) , .A( w0_20 ) );
  NAND2_X1 U74 (.A2( ld ) , .ZN( n72 ) , .A1( text_in[35] ) );
  XOR2_X1 U740 (.Z( n535 ) , .A( n538 ) , .B( n539 ) );
  XNOR2_X1 U741 (.B( n491 ) , .ZN( n538 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U742 (.A( n233 ) , .Z( n533 ) , .B( w0_20 ) );
  OAI22_X1 U744 (.ZN( N261 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n540 ) , .B1( n541 ) );
  XOR2_X1 U745 (.Z( n541 ) , .A( n542 ) , .B( n543 ) );
  XOR2_X1 U746 (.Z( n543 ) , .B( n544 ) , .A( sa10_sr_2 ) );
  XOR2_X1 U747 (.Z( n544 ) , .B( sa20_sr_2 ) , .A( w0_19 ) );
  OAI21_X1 U75 (.B1( ld ) , .ZN( n1014 ) , .B2( n73 ) , .A( n74 ) );
  XOR2_X1 U750 (.A( n231 ) , .Z( n540 ) , .B( w0_19 ) );
  OAI22_X1 U752 (.ZN( N260 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n546 ) , .B1( n547 ) );
  XOR2_X1 U755 (.Z( n550 ) , .B( sa20_sr_1 ) , .A( w0_18 ) );
  XNOR2_X1 U756 (.B( n503 ) , .ZN( n548 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U757 (.A( n229 ) , .Z( n546 ) , .B( w0_18 ) );
  OAI22_X1 U759 (.ZN( N259 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n551 ) , .B1( n552 ) );
  NAND2_X1 U76 (.A2( ld ) , .ZN( n74 ) , .A1( text_in[36] ) );
  XOR2_X1 U761 (.Z( n554 ) , .B( n555 ) , .A( sa10_sr_0 ) );
  XOR2_X1 U762 (.Z( n555 ) , .B( sa20_sr_0 ) , .A( w0_17 ) );
  XNOR2_X1 U764 (.B( n509 ) , .ZN( n556 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U765 (.A( n227 ) , .Z( n551 ) , .B( w0_17 ) );
  OAI22_X1 U767 (.ZN( N258 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n557 ) , .B1( n558 ) );
  XOR2_X1 U769 (.A( n516 ) , .B( n539 ) , .Z( n560 ) );
  OAI21_X1 U77 (.B1( ld ) , .ZN( n1015 ) , .B2( n75 ) , .A( n76 ) );
  XOR2_X1 U770 (.Z( n539 ) , .A( sa10_sr_7 ) , .B( sa20_sr_7 ) );
  XOR2_X1 U772 (.A( n225 ) , .Z( n557 ) , .B( w0_16 ) );
  OAI22_X1 U774 (.ZN( N249 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n561 ) , .B1( n562 ) );
  XOR2_X1 U776 (.A( n476 ) , .B( n488 ) , .Z( n564 ) );
  XOR2_X1 U777 (.Z( n476 ) , .A( sa20_sr_6 ) , .B( sa30_sr_6 ) );
  XOR2_X1 U779 (.A( n223 ) , .Z( n561 ) , .B( w0_15 ) );
  NAND2_X1 U78 (.A2( ld ) , .ZN( n76 ) , .A1( text_in[37] ) );
  OAI22_X1 U781 (.ZN( N248 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n565 ) , .B1( n566 ) );
  XOR2_X1 U783 (.A( n470 ) , .B( n482 ) , .Z( n568 ) );
  XOR2_X1 U784 (.Z( n482 ) , .A( sa20_sr_5 ) , .B( sa30_sr_5 ) );
  XOR2_X1 U786 (.A( n221 ) , .Z( n565 ) , .B( w0_14 ) );
  OAI22_X1 U788 (.ZN( N247 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n569 ) , .B1( n570 ) );
  XOR2_X1 U789 (.Z( n570 ) , .A( n571 ) , .B( n572 ) );
  OAI21_X1 U79 (.B1( ld ) , .ZN( n1016 ) , .B2( n77 ) , .A( n78 ) );
  XOR2_X1 U790 (.A( n477 ) , .B( n491 ) , .Z( n572 ) );
  XOR2_X1 U791 (.Z( n491 ) , .A( sa20_sr_4 ) , .B( sa30_sr_4 ) );
  XNOR2_X1 U792 (.ZN( n571 ) , .B( sa30_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U793 (.A( n219 ) , .Z( n569 ) , .B( w0_13 ) );
  OAI22_X1 U795 (.ZN( N246 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n573 ) , .B1( n574 ) );
  XOR2_X1 U796 (.Z( n574 ) , .A( n575 ) , .B( n576 ) );
  XOR2_X1 U797 (.A( n483 ) , .B( n496 ) , .Z( n576 ) );
  XOR2_X1 U798 (.Z( n496 ) , .A( sa20_sr_3 ) , .B( sa30_sr_3 ) );
  XOR2_X1 U799 (.B( n469 ) , .Z( n575 ) , .A( n577 ) );
  NAND2_X1 U8 (.A2( ld ) , .ZN( n6 ) , .A1( text_in[2] ) );
  NAND2_X1 U80 (.A2( ld ) , .ZN( n78 ) , .A1( text_in[38] ) );
  XNOR2_X1 U800 (.ZN( n577 ) , .B( sa30_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U801 (.A( n217 ) , .Z( n573 ) , .B( w0_12 ) );
  OAI22_X1 U803 (.ZN( N245 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n578 ) , .B1( n579 ) );
  XOR2_X1 U805 (.A( n489 ) , .B( n503 ) , .Z( n581 ) );
  XOR2_X1 U806 (.Z( n503 ) , .A( sa20_sr_2 ) , .B( sa30_sr_2 ) );
  XNOR2_X1 U808 (.ZN( n582 ) , .B( sa30_sr_3 ) , .A( w0_11 ) );
  XOR2_X1 U809 (.A( n215 ) , .Z( n578 ) , .B( w0_11 ) );
  OAI21_X1 U81 (.B1( ld ) , .ZN( n1017 ) , .B2( n79 ) , .A( n80 ) );
  OAI22_X1 U811 (.ZN( N244 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n583 ) , .B1( n584 ) );
  XOR2_X1 U813 (.A( n497 ) , .B( n509 ) , .Z( n586 ) );
  XOR2_X1 U814 (.Z( n509 ) , .A( sa20_sr_1 ) , .B( sa30_sr_1 ) );
  XOR2_X1 U816 (.A( n213 ) , .Z( n583 ) , .B( w0_10 ) );
  OAI22_X1 U818 (.ZN( N243 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n587 ) , .B1( n588 ) );
  NAND2_X1 U82 (.A2( ld ) , .ZN( n80 ) , .A1( text_in[39] ) );
  XOR2_X1 U820 (.A( n504 ) , .B( n516 ) , .Z( n590 ) );
  XOR2_X1 U821 (.Z( n516 ) , .A( sa20_sr_0 ) , .B( sa30_sr_0 ) );
  XNOR2_X1 U823 (.ZN( n591 ) , .B( sa30_sr_1 ) , .A( w0_9 ) );
  XOR2_X1 U824 (.A( n211 ) , .Z( n587 ) , .B( w0_9 ) );
  OAI22_X1 U826 (.ZN( N242 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n592 ) , .B1( n593 ) );
  XOR2_X1 U828 (.A( n469 ) , .B( n510 ) , .Z( n595 ) );
  XOR2_X1 U829 (.Z( n469 ) , .A( sa20_sr_7 ) , .B( sa30_sr_7 ) );
  OAI21_X1 U83 (.B1( ld ) , .ZN( n1018 ) , .B2( n81 ) , .A( n82 ) );
  XOR2_X1 U831 (.A( n209 ) , .Z( n592 ) , .B( w0_8 ) );
  OAI22_X1 U833 (.ZN( N233 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n596 ) , .B1( n597 ) );
  XOR2_X1 U834 (.Z( n597 ) , .A( n598 ) , .B( n599 ) );
  XOR2_X1 U835 (.B( n488 ) , .Z( n599 ) , .A( sa00_sr_6 ) );
  XOR2_X1 U836 (.Z( n488 ) , .A( sa00_sr_7 ) , .B( sa10_sr_7 ) );
  XNOR2_X1 U837 (.ZN( n598 ) , .B( n600 ) , .A( sa20_sr_7 ) );
  XOR2_X1 U838 (.Z( n600 ) , .B( sa30_sr_6 ) , .A( w0_7 ) );
  XOR2_X1 U839 (.A( n207 ) , .Z( n596 ) , .B( w0_7 ) );
  NAND2_X1 U84 (.A2( ld ) , .ZN( n82 ) , .A1( text_in[40] ) );
  OAI22_X1 U841 (.ZN( N232 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n601 ) , .B1( n602 ) );
  XOR2_X1 U844 (.Z( n605 ) , .B( sa30_sr_5 ) , .A( w0_6 ) );
  XNOR2_X1 U845 (.B( n470 ) , .ZN( n603 ) , .A( sa00_sr_5 ) );
  XOR2_X1 U846 (.Z( n470 ) , .A( sa00_sr_6 ) , .B( sa10_sr_6 ) );
  XOR2_X1 U847 (.A( n205 ) , .Z( n601 ) , .B( w0_6 ) );
  OAI22_X1 U849 (.ZN( N231 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n606 ) , .B1( n607 ) );
  OAI21_X1 U85 (.B1( ld ) , .ZN( n1019 ) , .B2( n83 ) , .A( n84 ) );
  XOR2_X1 U850 (.Z( n607 ) , .A( n608 ) , .B( n609 ) );
  XOR2_X1 U851 (.Z( n609 ) , .B( n610 ) , .A( sa20_sr_5 ) );
  XOR2_X1 U852 (.Z( n610 ) , .B( sa30_sr_4 ) , .A( w0_5 ) );
  XNOR2_X1 U853 (.B( n477 ) , .ZN( n608 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U854 (.Z( n477 ) , .A( sa00_sr_5 ) , .B( sa10_sr_5 ) );
  XOR2_X1 U855 (.A( n203 ) , .Z( n606 ) , .B( w0_5 ) );
  OAI22_X1 U857 (.ZN( N230 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n611 ) , .B1( n612 ) );
  XOR2_X1 U858 (.Z( n612 ) , .A( n613 ) , .B( n614 ) );
  XOR2_X1 U859 (.Z( n614 ) , .B( n615 ) , .A( sa20_sr_4 ) );
  NAND2_X1 U86 (.A2( ld ) , .ZN( n84 ) , .A1( text_in[41] ) );
  XOR2_X1 U860 (.Z( n615 ) , .B( sa30_sr_3 ) , .A( w0_4 ) );
  XOR2_X1 U861 (.Z( n613 ) , .A( n616 ) , .B( n617 ) );
  XNOR2_X1 U862 (.B( n483 ) , .ZN( n616 ) , .A( sa00_sr_3 ) );
  XOR2_X1 U863 (.Z( n483 ) , .A( sa00_sr_4 ) , .B( sa10_sr_4 ) );
  XOR2_X1 U864 (.A( n201 ) , .Z( n611 ) , .B( w0_4 ) );
  NOR4_X1 U866 (.ZN( N23 ) , .A3( ld ) , .A2( n1108 ) , .A4( n260 ) , .A1( n977 ) );
  NAND2_X1 U867 (.A1( n1106 ) , .A2( n1107 ) , .ZN( n260 ) );
  OAI22_X1 U868 (.ZN( N229 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n618 ) , .B1( n619 ) );
  OAI21_X1 U87 (.B1( ld ) , .ZN( n1020 ) , .B2( n85 ) , .A( n86 ) );
  XOR2_X1 U871 (.Z( n622 ) , .B( sa30_sr_2 ) , .A( w0_3 ) );
  XOR2_X1 U872 (.B( n617 ) , .Z( n620 ) , .A( n623 ) );
  XNOR2_X1 U873 (.B( n489 ) , .ZN( n623 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U874 (.Z( n489 ) , .A( sa00_sr_3 ) , .B( sa10_sr_3 ) );
  XOR2_X1 U875 (.A( n199 ) , .Z( n618 ) , .B( w0_3 ) );
  OAI22_X1 U877 (.ZN( N228 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n624 ) , .B1( n625 ) );
  NAND2_X1 U88 (.A2( ld ) , .ZN( n86 ) , .A1( text_in[42] ) );
  XOR2_X1 U880 (.Z( n628 ) , .B( sa30_sr_1 ) , .A( w0_2 ) );
  XNOR2_X1 U881 (.B( n497 ) , .ZN( n626 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U882 (.Z( n497 ) , .A( sa00_sr_2 ) , .B( sa10_sr_2 ) );
  XOR2_X1 U883 (.A( n197 ) , .Z( n624 ) , .B( w0_2 ) );
  OAI22_X1 U885 (.ZN( N227 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n629 ) , .B1( n630 ) );
  XOR2_X1 U887 (.Z( n632 ) , .B( n633 ) , .A( sa20_sr_1 ) );
  XOR2_X1 U888 (.Z( n633 ) , .B( sa30_sr_0 ) , .A( w0_1 ) );
  OAI21_X1 U89 (.B1( ld ) , .ZN( n1021 ) , .B2( n87 ) , .A( n88 ) );
  XNOR2_X1 U890 (.B( n504 ) , .ZN( n634 ) , .A( sa00_sr_0 ) );
  XOR2_X1 U891 (.Z( n504 ) , .A( sa00_sr_1 ) , .B( sa10_sr_1 ) );
  XOR2_X1 U892 (.A( n195 ) , .Z( n629 ) , .B( w0_1 ) );
  OAI22_X1 U894 (.ZN( N226 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n635 ) , .B1( n636 ) );
  XOR2_X1 U896 (.A( n510 ) , .B( n617 ) , .Z( n638 ) );
  XOR2_X1 U897 (.Z( n617 ) , .A( sa00_sr_7 ) , .B( sa30_sr_7 ) );
  XOR2_X1 U898 (.Z( n510 ) , .A( sa00_sr_0 ) , .B( sa10_sr_0 ) );
  OAI21_X1 U9 (.B1( ld ) , .B2( n7 ) , .A( n8 ) , .ZN( n981 ) );
  NAND2_X1 U90 (.A2( ld ) , .ZN( n88 ) , .A1( text_in[43] ) );
  XOR2_X1 U900 (.A( n193 ) , .Z( n635 ) , .B( w0_0 ) );
  OAI22_X1 U902 (.ZN( N217 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n639 ) , .B1( n640 ) );
  XOR2_X1 U904 (.Z( n642 ) , .A( n643 ) , .B( n644 ) );
  INV_X1 U906 (.ZN( n645 ) , .A( sa11_sr_7 ) );
  XOR2_X1 U907 (.A( n191 ) , .Z( n639 ) , .B( w1_31 ) );
  OAI22_X1 U909 (.ZN( N216 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n646 ) , .B1( n647 ) );
  OAI21_X1 U91 (.B1( ld ) , .ZN( n1022 ) , .B2( n89 ) , .A( n90 ) );
  XOR2_X1 U911 (.Z( n649 ) , .A( n650 ) , .B( n651 ) );
  XOR2_X1 U913 (.A( n189 ) , .Z( n646 ) , .B( w1_30 ) );
  OAI22_X1 U915 (.ZN( N215 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n652 ) , .B1( n653 ) );
  XOR2_X1 U917 (.Z( n655 ) , .A( n656 ) , .B( n657 ) );
  XOR2_X1 U919 (.A( n187 ) , .Z( n652 ) , .B( w1_29 ) );
  NAND2_X1 U92 (.A2( ld ) , .ZN( n90 ) , .A1( text_in[44] ) );
  OAI22_X1 U921 (.ZN( N214 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n658 ) , .B1( n659 ) );
  XOR2_X1 U922 (.Z( n659 ) , .A( n660 ) , .B( n661 ) );
  XOR2_X1 U923 (.Z( n661 ) , .A( n662 ) , .B( n663 ) );
  XOR2_X1 U924 (.Z( n660 ) , .A( n664 ) , .B( n665 ) );
  XNOR2_X1 U925 (.ZN( n664 ) , .B( sa11_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U926 (.A( n185 ) , .Z( n658 ) , .B( w1_28 ) );
  OAI22_X1 U928 (.ZN( N213 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n666 ) , .B1( n667 ) );
  OAI21_X1 U93 (.B1( ld ) , .ZN( n1023 ) , .B2( n91 ) , .A( n92 ) );
  XOR2_X1 U930 (.Z( n669 ) , .A( n670 ) , .B( n671 ) );
  XNOR2_X1 U932 (.ZN( n672 ) , .B( sa11_sr_3 ) , .A( w1_27 ) );
  XOR2_X1 U933 (.A( n183 ) , .Z( n666 ) , .B( w1_27 ) );
  OAI22_X1 U935 (.ZN( N212 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n673 ) , .B1( n674 ) );
  XOR2_X1 U937 (.Z( n676 ) , .A( n677 ) , .B( n678 ) );
  XOR2_X1 U939 (.A( n181 ) , .Z( n673 ) , .B( w1_26 ) );
  NAND2_X1 U94 (.A2( ld ) , .ZN( n92 ) , .A1( text_in[45] ) );
  OAI22_X1 U941 (.ZN( N211 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n679 ) , .B1( n680 ) );
  XOR2_X1 U943 (.Z( n682 ) , .A( n683 ) , .B( n684 ) );
  XNOR2_X1 U945 (.ZN( n685 ) , .B( sa11_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U946 (.A( n179 ) , .Z( n679 ) , .B( w1_25 ) );
  OAI22_X1 U948 (.ZN( N210 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n686 ) , .B1( n687 ) );
  OAI21_X1 U95 (.B1( ld ) , .ZN( n1024 ) , .B2( n93 ) , .A( n94 ) );
  XOR2_X1 U950 (.A( n665 ) , .Z( n689 ) , .B( n690 ) );
  XOR2_X1 U952 (.A( n177 ) , .Z( n686 ) , .B( w1_24 ) );
  OAI22_X1 U954 (.ZN( N201 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n691 ) , .B1( n692 ) );
  XOR2_X1 U955 (.Z( n692 ) , .A( n693 ) , .B( n694 ) );
  XOR2_X1 U956 (.B( n643 ) , .Z( n694 ) , .A( sa01_sr_7 ) );
  XOR2_X1 U959 (.A( n175 ) , .Z( n691 ) , .B( w1_23 ) );
  NAND2_X1 U96 (.A2( ld ) , .ZN( n94 ) , .A1( text_in[46] ) );
  OAI22_X1 U961 (.ZN( N200 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n696 ) , .B1( n697 ) );
  XOR2_X1 U964 (.Z( n700 ) , .B( sa21_sr_5 ) , .A( w1_22 ) );
  XOR2_X1 U967 (.A( n173 ) , .Z( n696 ) , .B( w1_22 ) );
  OAI22_X1 U969 (.ZN( N199 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n702 ) , .B1( n703 ) );
  OAI21_X1 U97 (.B1( ld ) , .ZN( n1025 ) , .B2( n95 ) , .A( n96 ) );
  XOR2_X1 U970 (.Z( n703 ) , .A( n704 ) , .B( n705 ) );
  XOR2_X1 U971 (.Z( n705 ) , .B( n706 ) , .A( sa11_sr_4 ) );
  XOR2_X1 U972 (.Z( n706 ) , .B( sa21_sr_4 ) , .A( w1_21 ) );
  XNOR2_X1 U973 (.B( n656 ) , .ZN( n704 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U974 (.A( n171 ) , .Z( n702 ) , .B( w1_21 ) );
  OAI22_X1 U976 (.ZN( N198 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n707 ) , .B1( n708 ) );
  XOR2_X1 U977 (.Z( n708 ) , .A( n709 ) , .B( n710 ) );
  XOR2_X1 U978 (.Z( n710 ) , .B( n711 ) , .A( sa11_sr_3 ) );
  XOR2_X1 U979 (.Z( n711 ) , .B( sa21_sr_3 ) , .A( w1_20 ) );
  NAND2_X1 U98 (.A2( ld ) , .ZN( n96 ) , .A1( text_in[47] ) );
  XOR2_X1 U980 (.Z( n709 ) , .A( n712 ) , .B( n713 ) );
  XNOR2_X1 U981 (.B( n663 ) , .ZN( n712 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U982 (.A( n169 ) , .Z( n707 ) , .B( w1_20 ) );
  OAI22_X1 U984 (.ZN( N197 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n714 ) , .B1( n715 ) );
  XOR2_X1 U987 (.Z( n718 ) , .B( sa21_sr_2 ) , .A( w1_19 ) );
  XOR2_X1 U988 (.B( n713 ) , .Z( n716 ) , .A( n719 ) );
  XNOR2_X1 U989 (.B( n670 ) , .ZN( n719 ) , .A( sa01_sr_3 ) );
  OAI21_X1 U99 (.B1( ld ) , .ZN( n1026 ) , .B2( n97 ) , .A( n98 ) );
  XOR2_X1 U990 (.A( n167 ) , .Z( n714 ) , .B( w1_19 ) );
  OAI22_X1 U992 (.ZN( N196 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n720 ) , .B1( n721 ) );
  XOR2_X1 U995 (.Z( n724 ) , .B( sa21_sr_1 ) , .A( w1_18 ) );
  XNOR2_X1 U996 (.B( n677 ) , .ZN( n722 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U997 (.A( n165 ) , .Z( n720 ) , .B( w1_18 ) );
  OAI22_X1 U999 (.ZN( N195 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n725 ) , .B1( n726 ) );
  DFF_X1 dcnt_reg_0 (.CK( clk ) , .QN( n1108 ) , .D( n1113 ) , .Q( n261 ) );
  DFF_X1 dcnt_reg_1 (.CK( clk ) , .D( n1110 ) , .Q( n977 ) );
  DFF_X1 dcnt_reg_2 (.CK( clk ) , .QN( n1107 ) , .D( n1111 ) , .Q( n267 ) );
  DFF_X1 dcnt_reg_3 (.CK( clk ) , .QN( n1106 ) , .D( n1112 ) );
  DFF_X1 done_reg (.D( N23 ) , .CK( clk ) , .Q( done ) );
  DFF_X1 ld_r_reg (.CK( clk ) , .D( ld ) , .QN( n1109 ) , .Q( n1114 ) );
  DFF_X1 sa00_reg_0 (.D( N274 ) , .CK( clk ) , .Q( sa00_0 ) );
  DFF_X1 sa00_reg_1 (.D( N275 ) , .CK( clk ) , .Q( sa00_1 ) );
  DFF_X1 sa00_reg_2 (.D( N276 ) , .CK( clk ) , .Q( sa00_2 ) );
  DFF_X1 sa00_reg_3 (.D( N277 ) , .CK( clk ) , .Q( sa00_3 ) );
  DFF_X1 sa00_reg_4 (.D( N278 ) , .CK( clk ) , .Q( sa00_4 ) );
  DFF_X1 sa00_reg_5 (.D( N279 ) , .CK( clk ) , .Q( sa00_5 ) );
  DFF_X1 sa00_reg_6 (.D( N280 ) , .CK( clk ) , .Q( sa00_6 ) );
  DFF_X1 sa00_reg_7 (.D( N281 ) , .CK( clk ) , .Q( sa00_7 ) );
  DFF_X1 sa01_reg_0 (.D( N210 ) , .CK( clk ) , .Q( sa01_0 ) );
  DFF_X1 sa01_reg_1 (.D( N211 ) , .CK( clk ) , .Q( sa01_1 ) );
  DFF_X1 sa01_reg_2 (.D( N212 ) , .CK( clk ) , .Q( sa01_2 ) );
  DFF_X1 sa01_reg_3 (.D( N213 ) , .CK( clk ) , .Q( sa01_3 ) );
  DFF_X1 sa01_reg_4 (.D( N214 ) , .CK( clk ) , .Q( sa01_4 ) );
  DFF_X1 sa01_reg_5 (.D( N215 ) , .CK( clk ) , .Q( sa01_5 ) );
  DFF_X1 sa01_reg_6 (.D( N216 ) , .CK( clk ) , .Q( sa01_6 ) );
  DFF_X1 sa01_reg_7 (.D( N217 ) , .CK( clk ) , .Q( sa01_7 ) );
  DFF_X1 sa02_reg_0 (.D( N146 ) , .CK( clk ) , .Q( sa02_0 ) );
  DFF_X1 sa02_reg_1 (.D( N147 ) , .CK( clk ) , .Q( sa02_1 ) );
  DFF_X1 sa02_reg_2 (.D( N148 ) , .CK( clk ) , .Q( sa02_2 ) );
  DFF_X1 sa02_reg_3 (.D( N149 ) , .CK( clk ) , .Q( sa02_3 ) );
  DFF_X1 sa02_reg_4 (.D( N150 ) , .CK( clk ) , .Q( sa02_4 ) );
  DFF_X1 sa02_reg_5 (.D( N151 ) , .CK( clk ) , .Q( sa02_5 ) );
  DFF_X1 sa02_reg_6 (.D( N152 ) , .CK( clk ) , .Q( sa02_6 ) );
  DFF_X1 sa02_reg_7 (.D( N153 ) , .CK( clk ) , .Q( sa02_7 ) );
  DFF_X1 sa03_reg_0 (.D( N82 ) , .CK( clk ) , .Q( sa03_0 ) );
  DFF_X1 sa03_reg_1 (.D( N83 ) , .CK( clk ) , .Q( sa03_1 ) );
  DFF_X1 sa03_reg_2 (.D( N84 ) , .CK( clk ) , .Q( sa03_2 ) );
  DFF_X1 sa03_reg_3 (.D( N85 ) , .CK( clk ) , .Q( sa03_3 ) );
  DFF_X1 sa03_reg_4 (.D( N86 ) , .CK( clk ) , .Q( sa03_4 ) );
  DFF_X1 sa03_reg_5 (.D( N87 ) , .CK( clk ) , .Q( sa03_5 ) );
  DFF_X1 sa03_reg_6 (.D( N88 ) , .CK( clk ) , .Q( sa03_6 ) );
  DFF_X1 sa03_reg_7 (.D( N89 ) , .CK( clk ) , .Q( sa03_7 ) );
  DFF_X1 sa10_reg_0 (.D( N258 ) , .CK( clk ) , .Q( sa10_0 ) );
  DFF_X1 sa10_reg_1 (.D( N259 ) , .CK( clk ) , .Q( sa10_1 ) );
  DFF_X1 sa10_reg_2 (.D( N260 ) , .CK( clk ) , .Q( sa10_2 ) );
  DFF_X1 sa10_reg_3 (.D( N261 ) , .CK( clk ) , .Q( sa10_3 ) );
  DFF_X1 sa10_reg_4 (.D( N262 ) , .CK( clk ) , .Q( sa10_4 ) );
  DFF_X1 sa10_reg_5 (.D( N263 ) , .CK( clk ) , .Q( sa10_5 ) );
  DFF_X1 sa10_reg_6 (.D( N264 ) , .CK( clk ) , .Q( sa10_6 ) );
  DFF_X1 sa10_reg_7 (.D( N265 ) , .CK( clk ) , .Q( sa10_7 ) );
  DFF_X1 sa11_reg_0 (.D( N194 ) , .CK( clk ) , .Q( sa11_0 ) );
  DFF_X1 sa11_reg_1 (.D( N195 ) , .CK( clk ) , .Q( sa11_1 ) );
  DFF_X1 sa11_reg_2 (.D( N196 ) , .CK( clk ) , .Q( sa11_2 ) );
  DFF_X1 sa11_reg_3 (.D( N197 ) , .CK( clk ) , .Q( sa11_3 ) );
  DFF_X1 sa11_reg_4 (.D( N198 ) , .CK( clk ) , .Q( sa11_4 ) );
  DFF_X1 sa11_reg_5 (.D( N199 ) , .CK( clk ) , .Q( sa11_5 ) );
  DFF_X1 sa11_reg_6 (.D( N200 ) , .CK( clk ) , .Q( sa11_6 ) );
  DFF_X1 sa11_reg_7 (.D( N201 ) , .CK( clk ) , .Q( sa11_7 ) );
  DFF_X1 sa12_reg_0 (.D( N130 ) , .CK( clk ) , .Q( sa12_0 ) );
  DFF_X1 sa12_reg_1 (.D( N131 ) , .CK( clk ) , .Q( sa12_1 ) );
  DFF_X1 sa12_reg_2 (.D( N132 ) , .CK( clk ) , .Q( sa12_2 ) );
  DFF_X1 sa12_reg_3 (.D( N133 ) , .CK( clk ) , .Q( sa12_3 ) );
  DFF_X1 sa12_reg_4 (.D( N134 ) , .CK( clk ) , .Q( sa12_4 ) );
  DFF_X1 sa12_reg_5 (.D( N135 ) , .CK( clk ) , .Q( sa12_5 ) );
  DFF_X1 sa12_reg_6 (.D( N136 ) , .CK( clk ) , .Q( sa12_6 ) );
  DFF_X1 sa12_reg_7 (.D( N137 ) , .CK( clk ) , .Q( sa12_7 ) );
  DFF_X1 sa13_reg_0 (.D( N66 ) , .CK( clk ) , .Q( sa13_0 ) );
  DFF_X1 sa13_reg_1 (.D( N67 ) , .CK( clk ) , .Q( sa13_1 ) );
  DFF_X1 sa13_reg_2 (.D( N68 ) , .CK( clk ) , .Q( sa13_2 ) );
  DFF_X1 sa13_reg_3 (.D( N69 ) , .CK( clk ) , .Q( sa13_3 ) );
  DFF_X1 sa13_reg_4 (.D( N70 ) , .CK( clk ) , .Q( sa13_4 ) );
  DFF_X1 sa13_reg_5 (.D( N71 ) , .CK( clk ) , .Q( sa13_5 ) );
  DFF_X1 sa13_reg_6 (.D( N72 ) , .CK( clk ) , .Q( sa13_6 ) );
  DFF_X1 sa13_reg_7 (.D( N73 ) , .CK( clk ) , .Q( sa13_7 ) );
  DFF_X1 sa20_reg_0 (.D( N242 ) , .CK( clk ) , .Q( sa20_0 ) );
  DFF_X1 sa20_reg_1 (.D( N243 ) , .CK( clk ) , .Q( sa20_1 ) );
  DFF_X1 sa20_reg_2 (.D( N244 ) , .CK( clk ) , .Q( sa20_2 ) );
  DFF_X1 sa20_reg_3 (.D( N245 ) , .CK( clk ) , .Q( sa20_3 ) );
  DFF_X1 sa20_reg_4 (.D( N246 ) , .CK( clk ) , .Q( sa20_4 ) );
  DFF_X1 sa20_reg_5 (.D( N247 ) , .CK( clk ) , .Q( sa20_5 ) );
  DFF_X1 sa20_reg_6 (.D( N248 ) , .CK( clk ) , .Q( sa20_6 ) );
  DFF_X1 sa20_reg_7 (.D( N249 ) , .CK( clk ) , .Q( sa20_7 ) );
  DFF_X1 sa21_reg_0 (.D( N178 ) , .CK( clk ) , .Q( sa21_0 ) );
  DFF_X1 sa21_reg_1 (.D( N179 ) , .CK( clk ) , .Q( sa21_1 ) );
  DFF_X1 sa21_reg_2 (.D( N180 ) , .CK( clk ) , .Q( sa21_2 ) );
  DFF_X1 sa21_reg_3 (.D( N181 ) , .CK( clk ) , .Q( sa21_3 ) );
  DFF_X1 sa21_reg_4 (.D( N182 ) , .CK( clk ) , .Q( sa21_4 ) );
  DFF_X1 sa21_reg_5 (.D( N183 ) , .CK( clk ) , .Q( sa21_5 ) );
  DFF_X1 sa21_reg_6 (.D( N184 ) , .CK( clk ) , .Q( sa21_6 ) );
  DFF_X1 sa21_reg_7 (.D( N185 ) , .CK( clk ) , .Q( sa21_7 ) );
  DFF_X1 sa22_reg_0 (.D( N114 ) , .CK( clk ) , .Q( sa22_0 ) );
  DFF_X1 sa22_reg_1 (.D( N115 ) , .CK( clk ) , .Q( sa22_1 ) );
  DFF_X1 sa22_reg_2 (.D( N116 ) , .CK( clk ) , .Q( sa22_2 ) );
  DFF_X1 sa22_reg_3 (.D( N117 ) , .CK( clk ) , .Q( sa22_3 ) );
  DFF_X1 sa22_reg_4 (.D( N118 ) , .CK( clk ) , .Q( sa22_4 ) );
  DFF_X1 sa22_reg_5 (.D( N119 ) , .CK( clk ) , .Q( sa22_5 ) );
  DFF_X1 sa22_reg_6 (.D( N120 ) , .CK( clk ) , .Q( sa22_6 ) );
  DFF_X1 sa22_reg_7 (.D( N121 ) , .CK( clk ) , .Q( sa22_7 ) );
  DFF_X1 sa23_reg_0 (.D( N50 ) , .CK( clk ) , .Q( sa23_0 ) );
  DFF_X1 sa23_reg_1 (.D( N51 ) , .CK( clk ) , .Q( sa23_1 ) );
  DFF_X1 sa23_reg_2 (.D( N52 ) , .CK( clk ) , .Q( sa23_2 ) );
  DFF_X1 sa23_reg_3 (.D( N53 ) , .CK( clk ) , .Q( sa23_3 ) );
  DFF_X1 sa23_reg_4 (.D( N54 ) , .CK( clk ) , .Q( sa23_4 ) );
  DFF_X1 sa23_reg_5 (.D( N55 ) , .CK( clk ) , .Q( sa23_5 ) );
  DFF_X1 sa23_reg_6 (.D( N56 ) , .CK( clk ) , .Q( sa23_6 ) );
  DFF_X1 sa23_reg_7 (.D( N57 ) , .CK( clk ) , .Q( sa23_7 ) );
  DFF_X1 sa30_reg_0 (.D( N226 ) , .CK( clk ) , .Q( sa30_0 ) );
  DFF_X1 sa30_reg_1 (.D( N227 ) , .CK( clk ) , .Q( sa30_1 ) );
  DFF_X1 sa30_reg_2 (.D( N228 ) , .CK( clk ) , .Q( sa30_2 ) );
  DFF_X1 sa30_reg_3 (.D( N229 ) , .CK( clk ) , .Q( sa30_3 ) );
  DFF_X1 sa30_reg_4 (.D( N230 ) , .CK( clk ) , .Q( sa30_4 ) );
  DFF_X1 sa30_reg_5 (.D( N231 ) , .CK( clk ) , .Q( sa30_5 ) );
  DFF_X1 sa30_reg_6 (.D( N232 ) , .CK( clk ) , .Q( sa30_6 ) );
  DFF_X1 sa30_reg_7 (.D( N233 ) , .CK( clk ) , .Q( sa30_7 ) );
  DFF_X1 sa31_reg_0 (.D( N162 ) , .CK( clk ) , .Q( sa31_0 ) );
  DFF_X1 sa31_reg_1 (.D( N163 ) , .CK( clk ) , .Q( sa31_1 ) );
  DFF_X1 sa31_reg_2 (.D( N164 ) , .CK( clk ) , .Q( sa31_2 ) );
  DFF_X1 sa31_reg_3 (.D( N165 ) , .CK( clk ) , .Q( sa31_3 ) );
  DFF_X1 sa31_reg_4 (.D( N166 ) , .CK( clk ) , .Q( sa31_4 ) );
  DFF_X1 sa31_reg_5 (.D( N167 ) , .CK( clk ) , .Q( sa31_5 ) );
  DFF_X1 sa31_reg_6 (.D( N168 ) , .CK( clk ) , .Q( sa31_6 ) );
  DFF_X1 sa31_reg_7 (.D( N169 ) , .CK( clk ) , .Q( sa31_7 ) );
  DFF_X1 sa32_reg_0 (.D( N98 ) , .CK( clk ) , .Q( sa32_0 ) );
  DFF_X1 sa32_reg_1 (.D( N99 ) , .CK( clk ) , .Q( sa32_1 ) );
  DFF_X1 sa32_reg_2 (.D( N100 ) , .CK( clk ) , .Q( sa32_2 ) );
  DFF_X1 sa32_reg_3 (.D( N101 ) , .CK( clk ) , .Q( sa32_3 ) );
  DFF_X1 sa32_reg_4 (.D( N102 ) , .CK( clk ) , .Q( sa32_4 ) );
  DFF_X1 sa32_reg_5 (.D( N103 ) , .CK( clk ) , .Q( sa32_5 ) );
  DFF_X1 sa32_reg_6 (.D( N104 ) , .CK( clk ) , .Q( sa32_6 ) );
  DFF_X1 sa32_reg_7 (.D( N105 ) , .CK( clk ) , .Q( sa32_7 ) );
  DFF_X1 sa33_reg_0 (.D( N34 ) , .CK( clk ) , .Q( sa33_0 ) );
  DFF_X1 sa33_reg_1 (.D( N35 ) , .CK( clk ) , .Q( sa33_1 ) );
  DFF_X1 sa33_reg_2 (.D( N36 ) , .CK( clk ) , .Q( sa33_2 ) );
  DFF_X1 sa33_reg_3 (.D( N37 ) , .CK( clk ) , .Q( sa33_3 ) );
  DFF_X1 sa33_reg_4 (.D( N38 ) , .CK( clk ) , .Q( sa33_4 ) );
  DFF_X1 sa33_reg_5 (.D( N39 ) , .CK( clk ) , .Q( sa33_5 ) );
  DFF_X1 sa33_reg_6 (.D( N40 ) , .CK( clk ) , .Q( sa33_6 ) );
  DFF_X1 sa33_reg_7 (.D( N41 ) , .CK( clk ) , .Q( sa33_7 ) );
  DFF_X1 text_in_r_reg_0 (.CK( clk ) , .QN( n1 ) , .D( n978 ) );
  DFF_X1 text_in_r_reg_1 (.CK( clk ) , .QN( n3 ) , .D( n979 ) );
  DFF_X1 text_in_r_reg_10 (.CK( clk ) , .QN( n21 ) , .D( n988 ) );
  DFF_X1 text_in_r_reg_100 (.CK( clk ) , .D( n1078 ) , .QN( n201 ) );
  DFF_X1 text_in_r_reg_101 (.CK( clk ) , .D( n1079 ) , .QN( n203 ) );
  DFF_X1 text_in_r_reg_102 (.CK( clk ) , .D( n1080 ) , .QN( n205 ) );
  DFF_X1 text_in_r_reg_103 (.CK( clk ) , .D( n1081 ) , .QN( n207 ) );
  DFF_X1 text_in_r_reg_104 (.CK( clk ) , .D( n1082 ) , .QN( n209 ) );
  DFF_X1 text_in_r_reg_105 (.CK( clk ) , .D( n1083 ) , .QN( n211 ) );
  DFF_X1 text_in_r_reg_106 (.CK( clk ) , .D( n1084 ) , .QN( n213 ) );
  DFF_X1 text_in_r_reg_107 (.CK( clk ) , .D( n1085 ) , .QN( n215 ) );
  DFF_X1 text_in_r_reg_108 (.CK( clk ) , .D( n1086 ) , .QN( n217 ) );
  DFF_X1 text_in_r_reg_109 (.CK( clk ) , .D( n1087 ) , .QN( n219 ) );
  DFF_X1 text_in_r_reg_11 (.CK( clk ) , .QN( n23 ) , .D( n989 ) );
  DFF_X1 text_in_r_reg_110 (.CK( clk ) , .D( n1088 ) , .QN( n221 ) );
  DFF_X1 text_in_r_reg_111 (.CK( clk ) , .D( n1089 ) , .QN( n223 ) );
  DFF_X1 text_in_r_reg_112 (.CK( clk ) , .D( n1090 ) , .QN( n225 ) );
  DFF_X1 text_in_r_reg_113 (.CK( clk ) , .D( n1091 ) , .QN( n227 ) );
  DFF_X1 text_in_r_reg_114 (.CK( clk ) , .D( n1092 ) , .QN( n229 ) );
  DFF_X1 text_in_r_reg_115 (.CK( clk ) , .D( n1093 ) , .QN( n231 ) );
  DFF_X1 text_in_r_reg_116 (.CK( clk ) , .D( n1094 ) , .QN( n233 ) );
  DFF_X1 text_in_r_reg_117 (.CK( clk ) , .D( n1095 ) , .QN( n235 ) );
  DFF_X1 text_in_r_reg_118 (.CK( clk ) , .D( n1096 ) , .QN( n237 ) );
  DFF_X1 text_in_r_reg_119 (.CK( clk ) , .D( n1097 ) , .QN( n239 ) );
  DFF_X1 text_in_r_reg_12 (.CK( clk ) , .QN( n25 ) , .D( n990 ) );
  DFF_X1 text_in_r_reg_120 (.CK( clk ) , .D( n1098 ) , .QN( n241 ) );
  DFF_X1 text_in_r_reg_121 (.CK( clk ) , .D( n1099 ) , .QN( n243 ) );
  DFF_X1 text_in_r_reg_122 (.CK( clk ) , .D( n1100 ) , .QN( n245 ) );
  DFF_X1 text_in_r_reg_123 (.CK( clk ) , .D( n1101 ) , .QN( n247 ) );
  DFF_X1 text_in_r_reg_124 (.CK( clk ) , .D( n1102 ) , .QN( n249 ) );
  DFF_X1 text_in_r_reg_125 (.CK( clk ) , .D( n1103 ) , .QN( n251 ) );
  DFF_X1 text_in_r_reg_126 (.CK( clk ) , .D( n1104 ) , .QN( n253 ) );
  DFF_X1 text_in_r_reg_127 (.CK( clk ) , .D( n1105 ) , .QN( n255 ) );
  DFF_X1 text_in_r_reg_13 (.CK( clk ) , .QN( n27 ) , .D( n991 ) );
  DFF_X1 text_in_r_reg_14 (.CK( clk ) , .QN( n29 ) , .D( n992 ) );
  DFF_X1 text_in_r_reg_15 (.CK( clk ) , .QN( n31 ) , .D( n993 ) );
  DFF_X1 text_in_r_reg_16 (.CK( clk ) , .QN( n33 ) , .D( n994 ) );
  DFF_X1 text_in_r_reg_17 (.CK( clk ) , .QN( n35 ) , .D( n995 ) );
  DFF_X1 text_in_r_reg_18 (.CK( clk ) , .QN( n37 ) , .D( n996 ) );
  DFF_X1 text_in_r_reg_19 (.CK( clk ) , .QN( n39 ) , .D( n997 ) );
  DFF_X1 text_in_r_reg_2 (.CK( clk ) , .QN( n5 ) , .D( n980 ) );
  DFF_X1 text_in_r_reg_20 (.CK( clk ) , .QN( n41 ) , .D( n998 ) );
  DFF_X1 text_in_r_reg_21 (.CK( clk ) , .QN( n43 ) , .D( n999 ) );
  DFF_X1 text_in_r_reg_22 (.CK( clk ) , .D( n1000 ) , .QN( n45 ) );
  DFF_X1 text_in_r_reg_23 (.CK( clk ) , .D( n1001 ) , .QN( n47 ) );
  DFF_X1 text_in_r_reg_24 (.CK( clk ) , .D( n1002 ) , .QN( n49 ) );
  DFF_X1 text_in_r_reg_25 (.CK( clk ) , .D( n1003 ) , .QN( n51 ) );
  DFF_X1 text_in_r_reg_26 (.CK( clk ) , .D( n1004 ) , .QN( n53 ) );
  DFF_X1 text_in_r_reg_27 (.CK( clk ) , .D( n1005 ) , .QN( n55 ) );
  DFF_X1 text_in_r_reg_28 (.CK( clk ) , .D( n1006 ) , .QN( n57 ) );
  DFF_X1 text_in_r_reg_29 (.CK( clk ) , .D( n1007 ) , .QN( n59 ) );
  DFF_X1 text_in_r_reg_3 (.CK( clk ) , .QN( n7 ) , .D( n981 ) );
  DFF_X1 text_in_r_reg_30 (.CK( clk ) , .D( n1008 ) , .QN( n61 ) );
  DFF_X1 text_in_r_reg_31 (.CK( clk ) , .D( n1009 ) , .QN( n63 ) );
  DFF_X1 text_in_r_reg_32 (.CK( clk ) , .D( n1010 ) , .QN( n65 ) );
  DFF_X1 text_in_r_reg_33 (.CK( clk ) , .D( n1011 ) , .QN( n67 ) );
  DFF_X1 text_in_r_reg_34 (.CK( clk ) , .D( n1012 ) , .QN( n69 ) );
  DFF_X1 text_in_r_reg_35 (.CK( clk ) , .D( n1013 ) , .QN( n71 ) );
  DFF_X1 text_in_r_reg_36 (.CK( clk ) , .D( n1014 ) , .QN( n73 ) );
  DFF_X1 text_in_r_reg_37 (.CK( clk ) , .D( n1015 ) , .QN( n75 ) );
  DFF_X1 text_in_r_reg_38 (.CK( clk ) , .D( n1016 ) , .QN( n77 ) );
  DFF_X1 text_in_r_reg_39 (.CK( clk ) , .D( n1017 ) , .QN( n79 ) );
  DFF_X1 text_in_r_reg_4 (.CK( clk ) , .QN( n9 ) , .D( n982 ) );
  DFF_X1 text_in_r_reg_40 (.CK( clk ) , .D( n1018 ) , .QN( n81 ) );
  DFF_X1 text_in_r_reg_41 (.CK( clk ) , .D( n1019 ) , .QN( n83 ) );
  DFF_X1 text_in_r_reg_42 (.CK( clk ) , .D( n1020 ) , .QN( n85 ) );
  DFF_X1 text_in_r_reg_43 (.CK( clk ) , .D( n1021 ) , .QN( n87 ) );
  DFF_X1 text_in_r_reg_44 (.CK( clk ) , .D( n1022 ) , .QN( n89 ) );
  DFF_X1 text_in_r_reg_45 (.CK( clk ) , .D( n1023 ) , .QN( n91 ) );
  DFF_X1 text_in_r_reg_46 (.CK( clk ) , .D( n1024 ) , .QN( n93 ) );
  DFF_X1 text_in_r_reg_47 (.CK( clk ) , .D( n1025 ) , .QN( n95 ) );
  DFF_X1 text_in_r_reg_48 (.CK( clk ) , .D( n1026 ) , .QN( n97 ) );
  DFF_X1 text_in_r_reg_49 (.CK( clk ) , .D( n1027 ) , .QN( n99 ) );
  DFF_X1 text_in_r_reg_5 (.CK( clk ) , .QN( n11 ) , .D( n983 ) );
  DFF_X1 text_in_r_reg_50 (.CK( clk ) , .QN( n101 ) , .D( n1028 ) );
  DFF_X1 text_in_r_reg_51 (.CK( clk ) , .D( n1029 ) , .QN( n103 ) );
  DFF_X1 text_in_r_reg_52 (.CK( clk ) , .D( n1030 ) , .QN( n105 ) );
  DFF_X1 text_in_r_reg_53 (.CK( clk ) , .D( n1031 ) , .QN( n107 ) );
  DFF_X1 text_in_r_reg_54 (.CK( clk ) , .D( n1032 ) , .QN( n109 ) );
  DFF_X1 text_in_r_reg_55 (.CK( clk ) , .D( n1033 ) , .QN( n111 ) );
  DFF_X1 text_in_r_reg_56 (.CK( clk ) , .D( n1034 ) , .QN( n113 ) );
  DFF_X1 text_in_r_reg_57 (.CK( clk ) , .D( n1035 ) , .QN( n115 ) );
  DFF_X1 text_in_r_reg_58 (.CK( clk ) , .D( n1036 ) , .QN( n117 ) );
  DFF_X1 text_in_r_reg_59 (.CK( clk ) , .D( n1037 ) , .QN( n119 ) );
  DFF_X1 text_in_r_reg_6 (.CK( clk ) , .QN( n13 ) , .D( n984 ) );
  DFF_X1 text_in_r_reg_60 (.CK( clk ) , .D( n1038 ) , .QN( n121 ) );
  DFF_X1 text_in_r_reg_61 (.CK( clk ) , .D( n1039 ) , .QN( n123 ) );
  DFF_X1 text_in_r_reg_62 (.CK( clk ) , .D( n1040 ) , .QN( n125 ) );
  DFF_X1 text_in_r_reg_63 (.CK( clk ) , .D( n1041 ) , .QN( n127 ) );
  DFF_X1 text_in_r_reg_64 (.CK( clk ) , .D( n1042 ) , .QN( n129 ) );
  DFF_X1 text_in_r_reg_65 (.CK( clk ) , .D( n1043 ) , .QN( n131 ) );
  DFF_X1 text_in_r_reg_66 (.CK( clk ) , .D( n1044 ) , .QN( n133 ) );
  DFF_X1 text_in_r_reg_67 (.CK( clk ) , .D( n1045 ) , .QN( n135 ) );
  DFF_X1 text_in_r_reg_68 (.CK( clk ) , .D( n1046 ) , .QN( n137 ) );
  DFF_X1 text_in_r_reg_69 (.CK( clk ) , .D( n1047 ) , .QN( n139 ) );
  DFF_X1 text_in_r_reg_7 (.CK( clk ) , .QN( n15 ) , .D( n985 ) );
  DFF_X1 text_in_r_reg_70 (.CK( clk ) , .D( n1048 ) , .QN( n141 ) );
  DFF_X1 text_in_r_reg_71 (.CK( clk ) , .D( n1049 ) , .QN( n143 ) );
  DFF_X1 text_in_r_reg_72 (.CK( clk ) , .D( n1050 ) , .QN( n145 ) );
  DFF_X1 text_in_r_reg_73 (.CK( clk ) , .D( n1051 ) , .QN( n147 ) );
  DFF_X1 text_in_r_reg_74 (.CK( clk ) , .D( n1052 ) , .QN( n149 ) );
  DFF_X1 text_in_r_reg_75 (.CK( clk ) , .D( n1053 ) , .QN( n151 ) );
  DFF_X1 text_in_r_reg_76 (.CK( clk ) , .D( n1054 ) , .QN( n153 ) );
  DFF_X1 text_in_r_reg_77 (.CK( clk ) , .D( n1055 ) , .QN( n155 ) );
  DFF_X1 text_in_r_reg_78 (.CK( clk ) , .D( n1056 ) , .QN( n157 ) );
  DFF_X1 text_in_r_reg_79 (.CK( clk ) , .D( n1057 ) , .QN( n159 ) );
  DFF_X1 text_in_r_reg_8 (.CK( clk ) , .QN( n17 ) , .D( n986 ) );
  DFF_X1 text_in_r_reg_80 (.CK( clk ) , .D( n1058 ) , .QN( n161 ) );
  DFF_X1 text_in_r_reg_81 (.CK( clk ) , .D( n1059 ) , .QN( n163 ) );
  DFF_X1 text_in_r_reg_82 (.CK( clk ) , .D( n1060 ) , .QN( n165 ) );
  DFF_X1 text_in_r_reg_83 (.CK( clk ) , .D( n1061 ) , .QN( n167 ) );
  DFF_X1 text_in_r_reg_84 (.CK( clk ) , .D( n1062 ) , .QN( n169 ) );
  DFF_X1 text_in_r_reg_85 (.CK( clk ) , .D( n1063 ) , .QN( n171 ) );
  DFF_X1 text_in_r_reg_86 (.CK( clk ) , .D( n1064 ) , .QN( n173 ) );
  DFF_X1 text_in_r_reg_87 (.CK( clk ) , .D( n1065 ) , .QN( n175 ) );
  DFF_X1 text_in_r_reg_88 (.CK( clk ) , .D( n1066 ) , .QN( n177 ) );
  DFF_X1 text_in_r_reg_89 (.CK( clk ) , .D( n1067 ) , .QN( n179 ) );
  DFF_X1 text_in_r_reg_9 (.CK( clk ) , .QN( n19 ) , .D( n987 ) );
  DFF_X1 text_in_r_reg_90 (.CK( clk ) , .D( n1068 ) , .QN( n181 ) );
  DFF_X1 text_in_r_reg_91 (.CK( clk ) , .D( n1069 ) , .QN( n183 ) );
  DFF_X1 text_in_r_reg_92 (.CK( clk ) , .D( n1070 ) , .QN( n185 ) );
  DFF_X1 text_in_r_reg_93 (.CK( clk ) , .D( n1071 ) , .QN( n187 ) );
  DFF_X1 text_in_r_reg_94 (.CK( clk ) , .D( n1072 ) , .QN( n189 ) );
  DFF_X1 text_in_r_reg_95 (.CK( clk ) , .D( n1073 ) , .QN( n191 ) );
  DFF_X1 text_in_r_reg_96 (.CK( clk ) , .D( n1074 ) , .QN( n193 ) );
  DFF_X1 text_in_r_reg_97 (.CK( clk ) , .D( n1075 ) , .QN( n195 ) );
  DFF_X1 text_in_r_reg_98 (.CK( clk ) , .D( n1076 ) , .QN( n197 ) );
  DFF_X1 text_in_r_reg_99 (.CK( clk ) , .D( n1077 ) , .QN( n199 ) );
  DFF_X1 text_out_reg_0 (.D( N505 ) , .CK( clk ) , .Q( text_out[0] ) );
  DFF_X1 text_out_reg_1 (.D( N504 ) , .CK( clk ) , .Q( text_out[1] ) );
  DFF_X1 text_out_reg_10 (.D( N471 ) , .CK( clk ) , .Q( text_out[10] ) );
  DFF_X1 text_out_reg_100 (.D( N477 ) , .CK( clk ) , .Q( text_out[100] ) );
  DFF_X1 text_out_reg_101 (.D( N476 ) , .CK( clk ) , .Q( text_out[101] ) );
  DFF_X1 text_out_reg_102 (.D( N475 ) , .CK( clk ) , .Q( text_out[102] ) );
  DFF_X1 text_out_reg_103 (.D( N474 ) , .CK( clk ) , .Q( text_out[103] ) );
  DFF_X1 text_out_reg_104 (.D( N449 ) , .CK( clk ) , .Q( text_out[104] ) );
  DFF_X1 text_out_reg_105 (.D( N448 ) , .CK( clk ) , .Q( text_out[105] ) );
  DFF_X1 text_out_reg_106 (.D( N447 ) , .CK( clk ) , .Q( text_out[106] ) );
  DFF_X1 text_out_reg_107 (.D( N446 ) , .CK( clk ) , .Q( text_out[107] ) );
  DFF_X1 text_out_reg_108 (.D( N445 ) , .CK( clk ) , .Q( text_out[108] ) );
  DFF_X1 text_out_reg_109 (.D( N444 ) , .CK( clk ) , .Q( text_out[109] ) );
  DFF_X1 text_out_reg_11 (.D( N470 ) , .CK( clk ) , .Q( text_out[11] ) );
  DFF_X1 text_out_reg_110 (.D( N443 ) , .CK( clk ) , .Q( text_out[110] ) );
  DFF_X1 text_out_reg_111 (.D( N442 ) , .CK( clk ) , .Q( text_out[111] ) );
  DFF_X1 text_out_reg_112 (.D( N417 ) , .CK( clk ) , .Q( text_out[112] ) );
  DFF_X1 text_out_reg_113 (.D( N416 ) , .CK( clk ) , .Q( text_out[113] ) );
  DFF_X1 text_out_reg_114 (.D( N415 ) , .CK( clk ) , .Q( text_out[114] ) );
  DFF_X1 text_out_reg_115 (.D( N414 ) , .CK( clk ) , .Q( text_out[115] ) );
  DFF_X1 text_out_reg_116 (.D( N413 ) , .CK( clk ) , .Q( text_out[116] ) );
  DFF_X1 text_out_reg_117 (.D( N412 ) , .CK( clk ) , .Q( text_out[117] ) );
  DFF_X1 text_out_reg_118 (.D( N411 ) , .CK( clk ) , .Q( text_out[118] ) );
  DFF_X1 text_out_reg_119 (.D( N410 ) , .CK( clk ) , .Q( text_out[119] ) );
  DFF_X1 text_out_reg_12 (.D( N469 ) , .CK( clk ) , .Q( text_out[12] ) );
  DFF_X1 text_out_reg_120 (.D( N385 ) , .CK( clk ) , .Q( text_out[120] ) );
  DFF_X1 text_out_reg_121 (.D( N384 ) , .CK( clk ) , .Q( text_out[121] ) );
  DFF_X1 text_out_reg_122 (.D( N383 ) , .CK( clk ) , .Q( text_out[122] ) );
  DFF_X1 text_out_reg_123 (.D( N382 ) , .CK( clk ) , .Q( text_out[123] ) );
  DFF_X1 text_out_reg_124 (.D( N381 ) , .CK( clk ) , .Q( text_out[124] ) );
  DFF_X1 text_out_reg_125 (.D( N380 ) , .CK( clk ) , .Q( text_out[125] ) );
  DFF_X1 text_out_reg_126 (.D( N379 ) , .CK( clk ) , .Q( text_out[126] ) );
  DFF_X1 text_out_reg_127 (.D( N378 ) , .CK( clk ) , .Q( text_out[127] ) );
  DFF_X1 text_out_reg_13 (.D( N468 ) , .CK( clk ) , .Q( text_out[13] ) );
  DFF_X1 text_out_reg_14 (.D( N467 ) , .CK( clk ) , .Q( text_out[14] ) );
  DFF_X1 text_out_reg_15 (.D( N466 ) , .CK( clk ) , .Q( text_out[15] ) );
  DFF_X1 text_out_reg_16 (.D( N441 ) , .CK( clk ) , .Q( text_out[16] ) );
  DFF_X1 text_out_reg_17 (.D( N440 ) , .CK( clk ) , .Q( text_out[17] ) );
  DFF_X1 text_out_reg_18 (.D( N439 ) , .CK( clk ) , .Q( text_out[18] ) );
  DFF_X1 text_out_reg_19 (.D( N438 ) , .CK( clk ) , .Q( text_out[19] ) );
  DFF_X1 text_out_reg_2 (.D( N503 ) , .CK( clk ) , .Q( text_out[2] ) );
  DFF_X1 text_out_reg_20 (.D( N437 ) , .CK( clk ) , .Q( text_out[20] ) );
  DFF_X1 text_out_reg_21 (.D( N436 ) , .CK( clk ) , .Q( text_out[21] ) );
  DFF_X1 text_out_reg_22 (.D( N435 ) , .CK( clk ) , .Q( text_out[22] ) );
  DFF_X1 text_out_reg_23 (.D( N434 ) , .CK( clk ) , .Q( text_out[23] ) );
  DFF_X1 text_out_reg_24 (.D( N409 ) , .CK( clk ) , .Q( text_out[24] ) );
  DFF_X1 text_out_reg_25 (.D( N408 ) , .CK( clk ) , .Q( text_out[25] ) );
  DFF_X1 text_out_reg_26 (.D( N407 ) , .CK( clk ) , .Q( text_out[26] ) );
  DFF_X1 text_out_reg_27 (.D( N406 ) , .CK( clk ) , .Q( text_out[27] ) );
  DFF_X1 text_out_reg_28 (.D( N405 ) , .CK( clk ) , .Q( text_out[28] ) );
  DFF_X1 text_out_reg_29 (.D( N404 ) , .CK( clk ) , .Q( text_out[29] ) );
  DFF_X1 text_out_reg_3 (.D( N502 ) , .CK( clk ) , .Q( text_out[3] ) );
  DFF_X1 text_out_reg_30 (.D( N403 ) , .CK( clk ) , .Q( text_out[30] ) );
  DFF_X1 text_out_reg_31 (.D( N402 ) , .CK( clk ) , .Q( text_out[31] ) );
  DFF_X1 text_out_reg_32 (.D( N497 ) , .CK( clk ) , .Q( text_out[32] ) );
  DFF_X1 text_out_reg_33 (.D( N496 ) , .CK( clk ) , .Q( text_out[33] ) );
  DFF_X1 text_out_reg_34 (.D( N495 ) , .CK( clk ) , .Q( text_out[34] ) );
  DFF_X1 text_out_reg_35 (.D( N494 ) , .CK( clk ) , .Q( text_out[35] ) );
  DFF_X1 text_out_reg_36 (.D( N493 ) , .CK( clk ) , .Q( text_out[36] ) );
  DFF_X1 text_out_reg_37 (.D( N492 ) , .CK( clk ) , .Q( text_out[37] ) );
  DFF_X1 text_out_reg_38 (.D( N491 ) , .CK( clk ) , .Q( text_out[38] ) );
  DFF_X1 text_out_reg_39 (.D( N490 ) , .CK( clk ) , .Q( text_out[39] ) );
  DFF_X1 text_out_reg_4 (.D( N501 ) , .CK( clk ) , .Q( text_out[4] ) );
  DFF_X1 text_out_reg_40 (.D( N465 ) , .CK( clk ) , .Q( text_out[40] ) );
  DFF_X1 text_out_reg_41 (.D( N464 ) , .CK( clk ) , .Q( text_out[41] ) );
  DFF_X1 text_out_reg_42 (.D( N463 ) , .CK( clk ) , .Q( text_out[42] ) );
  DFF_X1 text_out_reg_43 (.D( N462 ) , .CK( clk ) , .Q( text_out[43] ) );
  DFF_X1 text_out_reg_44 (.D( N461 ) , .CK( clk ) , .Q( text_out[44] ) );
  DFF_X1 text_out_reg_45 (.D( N460 ) , .CK( clk ) , .Q( text_out[45] ) );
  DFF_X1 text_out_reg_46 (.D( N459 ) , .CK( clk ) , .Q( text_out[46] ) );
  DFF_X1 text_out_reg_47 (.D( N458 ) , .CK( clk ) , .Q( text_out[47] ) );
  DFF_X1 text_out_reg_48 (.D( N433 ) , .CK( clk ) , .Q( text_out[48] ) );
  DFF_X1 text_out_reg_49 (.D( N432 ) , .CK( clk ) , .Q( text_out[49] ) );
  DFF_X1 text_out_reg_5 (.D( N500 ) , .CK( clk ) , .Q( text_out[5] ) );
  DFF_X1 text_out_reg_50 (.D( N431 ) , .CK( clk ) , .Q( text_out[50] ) );
  DFF_X1 text_out_reg_51 (.D( N430 ) , .CK( clk ) , .Q( text_out[51] ) );
  DFF_X1 text_out_reg_52 (.D( N429 ) , .CK( clk ) , .Q( text_out[52] ) );
  DFF_X1 text_out_reg_53 (.D( N428 ) , .CK( clk ) , .Q( text_out[53] ) );
  DFF_X1 text_out_reg_54 (.D( N427 ) , .CK( clk ) , .Q( text_out[54] ) );
  DFF_X1 text_out_reg_55 (.D( N426 ) , .CK( clk ) , .Q( text_out[55] ) );
  DFF_X1 text_out_reg_56 (.D( N401 ) , .CK( clk ) , .Q( text_out[56] ) );
  DFF_X1 text_out_reg_57 (.D( N400 ) , .CK( clk ) , .Q( text_out[57] ) );
  DFF_X1 text_out_reg_58 (.D( N399 ) , .CK( clk ) , .Q( text_out[58] ) );
  DFF_X1 text_out_reg_59 (.D( N398 ) , .CK( clk ) , .Q( text_out[59] ) );
  DFF_X1 text_out_reg_6 (.D( N499 ) , .CK( clk ) , .Q( text_out[6] ) );
  DFF_X1 text_out_reg_60 (.D( N397 ) , .CK( clk ) , .Q( text_out[60] ) );
  DFF_X1 text_out_reg_61 (.D( N396 ) , .CK( clk ) , .Q( text_out[61] ) );
  DFF_X1 text_out_reg_62 (.D( N395 ) , .CK( clk ) , .Q( text_out[62] ) );
  DFF_X1 text_out_reg_63 (.D( N394 ) , .CK( clk ) , .Q( text_out[63] ) );
  DFF_X1 text_out_reg_64 (.D( N489 ) , .CK( clk ) , .Q( text_out[64] ) );
  DFF_X1 text_out_reg_65 (.D( N488 ) , .CK( clk ) , .Q( text_out[65] ) );
  DFF_X1 text_out_reg_66 (.D( N487 ) , .CK( clk ) , .Q( text_out[66] ) );
  DFF_X1 text_out_reg_67 (.D( N486 ) , .CK( clk ) , .Q( text_out[67] ) );
  DFF_X1 text_out_reg_68 (.D( N485 ) , .CK( clk ) , .Q( text_out[68] ) );
  DFF_X1 text_out_reg_69 (.D( N484 ) , .CK( clk ) , .Q( text_out[69] ) );
  DFF_X1 text_out_reg_7 (.D( N498 ) , .CK( clk ) , .Q( text_out[7] ) );
  DFF_X1 text_out_reg_70 (.D( N483 ) , .CK( clk ) , .Q( text_out[70] ) );
  DFF_X1 text_out_reg_71 (.D( N482 ) , .CK( clk ) , .Q( text_out[71] ) );
  DFF_X1 text_out_reg_72 (.D( N457 ) , .CK( clk ) , .Q( text_out[72] ) );
  DFF_X1 text_out_reg_73 (.D( N456 ) , .CK( clk ) , .Q( text_out[73] ) );
  DFF_X1 text_out_reg_74 (.D( N455 ) , .CK( clk ) , .Q( text_out[74] ) );
  DFF_X1 text_out_reg_75 (.D( N454 ) , .CK( clk ) , .Q( text_out[75] ) );
  DFF_X1 text_out_reg_76 (.D( N453 ) , .CK( clk ) , .Q( text_out[76] ) );
  DFF_X1 text_out_reg_77 (.D( N452 ) , .CK( clk ) , .Q( text_out[77] ) );
  DFF_X1 text_out_reg_78 (.D( N451 ) , .CK( clk ) , .Q( text_out[78] ) );
  DFF_X1 text_out_reg_79 (.D( N450 ) , .CK( clk ) , .Q( text_out[79] ) );
  DFF_X1 text_out_reg_8 (.D( N473 ) , .CK( clk ) , .Q( text_out[8] ) );
  DFF_X1 text_out_reg_80 (.D( N425 ) , .CK( clk ) , .Q( text_out[80] ) );
  DFF_X1 text_out_reg_81 (.D( N424 ) , .CK( clk ) , .Q( text_out[81] ) );
  DFF_X1 text_out_reg_82 (.D( N423 ) , .CK( clk ) , .Q( text_out[82] ) );
  DFF_X1 text_out_reg_83 (.D( N422 ) , .CK( clk ) , .Q( text_out[83] ) );
  DFF_X1 text_out_reg_84 (.D( N421 ) , .CK( clk ) , .Q( text_out[84] ) );
  DFF_X1 text_out_reg_85 (.D( N420 ) , .CK( clk ) , .Q( text_out[85] ) );
  DFF_X1 text_out_reg_86 (.D( N419 ) , .CK( clk ) , .Q( text_out[86] ) );
  DFF_X1 text_out_reg_87 (.D( N418 ) , .CK( clk ) , .Q( text_out[87] ) );
  DFF_X1 text_out_reg_88 (.D( N393 ) , .CK( clk ) , .Q( text_out[88] ) );
  DFF_X1 text_out_reg_89 (.D( N392 ) , .CK( clk ) , .Q( text_out[89] ) );
  DFF_X1 text_out_reg_9 (.D( N472 ) , .CK( clk ) , .Q( text_out[9] ) );
  DFF_X1 text_out_reg_90 (.D( N391 ) , .CK( clk ) , .Q( text_out[90] ) );
  DFF_X1 text_out_reg_91 (.D( N390 ) , .CK( clk ) , .Q( text_out[91] ) );
  DFF_X1 text_out_reg_92 (.D( N389 ) , .CK( clk ) , .Q( text_out[92] ) );
  DFF_X1 text_out_reg_93 (.D( N388 ) , .CK( clk ) , .Q( text_out[93] ) );
  DFF_X1 text_out_reg_94 (.D( N387 ) , .CK( clk ) , .Q( text_out[94] ) );
  DFF_X1 text_out_reg_95 (.D( N386 ) , .CK( clk ) , .Q( text_out[95] ) );
  DFF_X1 text_out_reg_96 (.D( N481 ) , .CK( clk ) , .Q( text_out[96] ) );
  DFF_X1 text_out_reg_97 (.D( N480 ) , .CK( clk ) , .Q( text_out[97] ) );
  DFF_X1 text_out_reg_98 (.D( N479 ) , .CK( clk ) , .Q( text_out[98] ) );
  DFF_X1 text_out_reg_99 (.D( N478 ) , .CK( clk ) , .Q( text_out[99] ) );
  XNOR2_X1 u0_U10 (.ZN( u0_n57 ) , .B( u0_subword_3 ) , .A( w0_3 ) );
  NAND2_X1 u0_U100 (.A1( key[62] ) , .A2( ld ) , .ZN( u0_n163 ) );
  NAND2_X1 u0_U101 (.A1( key[15] ) , .A2( ld ) , .ZN( u0_n114 ) );
  NAND2_X1 u0_U102 (.A1( key[74] ) , .A2( ld ) , .ZN( u0_n267 ) );
  NAND2_X1 u0_U103 (.A1( key[10] ) , .A2( ld ) , .ZN( u0_n129 ) );
  NAND2_X1 u0_U104 (.A1( key[72] ) , .A2( ld ) , .ZN( u0_n271 ) );
  NAND2_X1 u0_U105 (.A2( key[127] ) , .A1( ld ) , .ZN( u0_n2 ) );
  NAND2_X1 u0_U106 (.A1( key[6] ) , .A2( ld ) , .ZN( u0_n141 ) );
  NAND2_X1 u0_U107 (.A1( key[2] ) , .A2( ld ) , .ZN( u0_n153 ) );
  NAND2_X1 u0_U108 (.A1( key[73] ) , .A2( ld ) , .ZN( u0_n269 ) );
  NAND2_X1 u0_U109 (.A1( key[30] ) , .A2( ld ) , .ZN( u0_n69 ) );
  XNOR2_X1 u0_U11 (.ZN( u0_n41 ) , .B( u0_subword_11 ) , .A( w0_11 ) );
  NAND2_X1 u0_U110 (.A1( key[29] ) , .A2( ld ) , .ZN( u0_n72 ) );
  NAND2_X1 u0_U111 (.A1( key[17] ) , .A2( ld ) , .ZN( u0_n108 ) );
  NAND2_X1 u0_U112 (.A1( key[18] ) , .A2( ld ) , .ZN( u0_n105 ) );
  NAND2_X1 u0_U113 (.A1( key[16] ) , .A2( ld ) , .ZN( u0_n111 ) );
  NAND2_X1 u0_U114 (.A1( key[9] ) , .A2( ld ) , .ZN( u0_n132 ) );
  NAND2_X1 u0_U115 (.A1( key[19] ) , .A2( ld ) , .ZN( u0_n102 ) );
  NAND2_X1 u0_U116 (.A1( key[8] ) , .A2( ld ) , .ZN( u0_n135 ) );
  NAND2_X1 u0_U117 (.A1( key[3] ) , .A2( ld ) , .ZN( u0_n150 ) );
  NAND2_X1 u0_U118 (.A1( key[0] ) , .A2( ld ) , .ZN( u0_n159 ) );
  NAND2_X1 u0_U119 (.A1( key[5] ) , .A2( ld ) , .ZN( u0_n144 ) );
  XNOR2_X1 u0_U12 (.ZN( u0_n33 ) , .B( u0_subword_15 ) , .A( w0_15 ) );
  NAND2_X1 u0_U120 (.A1( key[1] ) , .A2( ld ) , .ZN( u0_n156 ) );
  OAI21_X1 u0_U121 (.B1( ld ) , .ZN( u0_N181 ) , .B2( u0_n139 ) , .A( u0_n209 ) );
  NAND2_X1 u0_U122 (.A1( key[39] ) , .A2( ld ) , .ZN( u0_n209 ) );
  OAI21_X1 u0_U123 (.B1( ld ) , .ZN( u0_N135 ) , .B2( u0_n170 ) , .A( u0_n233 ) );
  NAND2_X1 u0_U124 (.A1( key[91] ) , .A2( ld ) , .ZN( u0_n233 ) );
  OAI21_X1 u0_U125 (.B1( ld ) , .ZN( u0_N57 ) , .B2( u0_n33 ) , .A( u0_n34 ) );
  NAND2_X1 u0_U126 (.A1( key[111] ) , .A2( ld ) , .ZN( u0_n34 ) );
  OAI21_X1 u0_U127 (.B1( ld ) , .ZN( u0_N46 ) , .B2( u0_n55 ) , .A( u0_n56 ) );
  NAND2_X1 u0_U128 (.A1( key[100] ) , .A2( ld ) , .ZN( u0_n56 ) );
  OAI21_X1 u0_U129 (.B1( ld ) , .ZN( u0_N45 ) , .B2( u0_n57 ) , .A( u0_n58 ) );
  XNOR2_X1 u0_U13 (.ZN( u0_n17 ) , .B( u0_subword_23 ) , .A( w0_23 ) );
  NAND2_X1 u0_U130 (.A1( key[99] ) , .A2( ld ) , .ZN( u0_n58 ) );
  OAI21_X1 u0_U131 (.B1( ld ) , .ZN( u0_N43 ) , .B2( u0_n61 ) , .A( u0_n62 ) );
  NAND2_X1 u0_U132 (.A1( key[97] ) , .A2( ld ) , .ZN( u0_n62 ) );
  OAI21_X1 u0_U133 (.B1( ld ) , .ZN( u0_N54 ) , .B2( u0_n39 ) , .A( u0_n40 ) );
  NAND2_X1 u0_U134 (.A1( key[108] ) , .A2( ld ) , .ZN( u0_n40 ) );
  OAI21_X1 u0_U135 (.B1( ld ) , .ZN( u0_N51 ) , .B2( u0_n45 ) , .A( u0_n46 ) );
  NAND2_X1 u0_U136 (.A1( key[105] ) , .A2( ld ) , .ZN( u0_n46 ) );
  OAI21_X1 u0_U137 (.B1( ld ) , .ZN( u0_N65 ) , .B2( u0_n17 ) , .A( u0_n18 ) );
  NAND2_X1 u0_U138 (.A1( key[119] ) , .A2( ld ) , .ZN( u0_n18 ) );
  OAI21_X1 u0_U139 (.B1( ld ) , .ZN( u0_N71 ) , .B2( u0_n5 ) , .A( u0_n6 ) );
  XNOR2_X1 u0_U14 (.ZN( u0_n45 ) , .B( u0_subword_9 ) , .A( w0_9 ) );
  NAND2_X1 u0_U140 (.A1( key[125] ) , .A2( ld ) , .ZN( u0_n6 ) );
  OAI21_X1 u0_U141 (.B1( ld ) , .ZN( u0_N70 ) , .B2( u0_n7 ) , .A( u0_n8 ) );
  NAND2_X1 u0_U142 (.A1( key[124] ) , .A2( ld ) , .ZN( u0_n8 ) );
  OAI21_X1 u0_U143 (.B1( ld ) , .ZN( u0_N69 ) , .A( u0_n10 ) , .B2( u0_n9 ) );
  NAND2_X1 u0_U144 (.A1( key[123] ) , .A2( ld ) , .ZN( u0_n10 ) );
  OAI21_X1 u0_U145 (.B1( ld ) , .ZN( u0_N123 ) , .B2( u0_n194 ) , .A( u0_n257 ) );
  NAND2_X1 u0_U146 (.A1( key[79] ) , .A2( ld ) , .ZN( u0_n257 ) );
  OAI21_X1 u0_U147 (.B1( ld ) , .ZN( u0_N131 ) , .B2( u0_n178 ) , .A( u0_n241 ) );
  NAND2_X1 u0_U148 (.A1( key[87] ) , .A2( ld ) , .ZN( u0_n241 ) );
  OAI21_X1 u0_U149 (.B1( ld ) , .ZN( u0_N121 ) , .B2( u0_n198 ) , .A( u0_n261 ) );
  XNOR2_X1 u0_U15 (.ZN( u0_n23 ) , .B( u0_subword_20 ) , .A( w0_20 ) );
  NAND2_X1 u0_U150 (.A1( key[77] ) , .A2( ld ) , .ZN( u0_n261 ) );
  OAI21_X1 u0_U151 (.B1( ld ) , .ZN( u0_N47 ) , .B2( u0_n53 ) , .A( u0_n54 ) );
  NAND2_X1 u0_U152 (.A1( key[101] ) , .A2( ld ) , .ZN( u0_n54 ) );
  OAI21_X1 u0_U153 (.B1( ld ) , .ZN( u0_N63 ) , .B2( u0_n21 ) , .A( u0_n22 ) );
  NAND2_X1 u0_U154 (.A1( key[117] ) , .A2( ld ) , .ZN( u0_n22 ) );
  OAI21_X1 u0_U155 (.B1( ld ) , .ZN( u0_N129 ) , .B2( u0_n182 ) , .A( u0_n245 ) );
  NAND2_X1 u0_U156 (.A1( key[85] ) , .A2( ld ) , .ZN( u0_n245 ) );
  OAI21_X1 u0_U157 (.B1( ld ) , .ZN( u0_N62 ) , .B2( u0_n23 ) , .A( u0_n24 ) );
  NAND2_X1 u0_U158 (.A1( key[116] ) , .A2( ld ) , .ZN( u0_n24 ) );
  OAI21_X1 u0_U159 (.B1( ld ) , .ZN( u0_N55 ) , .B2( u0_n37 ) , .A( u0_n38 ) );
  XNOR2_X1 u0_U16 (.ZN( u0_n37 ) , .B( u0_subword_13 ) , .A( w0_13 ) );
  NAND2_X1 u0_U160 (.A1( key[109] ) , .A2( ld ) , .ZN( u0_n38 ) );
  OAI21_X1 u0_U161 (.B1( ld ) , .ZN( u0_N120 ) , .B2( u0_n200 ) , .A( u0_n263 ) );
  NAND2_X1 u0_U162 (.A1( key[76] ) , .A2( ld ) , .ZN( u0_n263 ) );
  OAI21_X1 u0_U163 (.B1( ld ) , .ZN( u0_N53 ) , .B2( u0_n41 ) , .A( u0_n42 ) );
  NAND2_X1 u0_U164 (.A1( key[107] ) , .A2( ld ) , .ZN( u0_n42 ) );
  OAI21_X1 u0_U165 (.B1( ld ) , .ZN( u0_N268 ) , .B2( u0_n74 ) , .A( u0_n75 ) );
  NAND2_X1 u0_U166 (.A1( key[28] ) , .A2( ld ) , .ZN( u0_n75 ) );
  OAI21_X1 u0_U167 (.B1( ld ) , .ZN( u0_N271 ) , .B2( u0_n65 ) , .A( u0_n66 ) );
  NAND2_X1 u0_U168 (.A1( key[31] ) , .A2( ld ) , .ZN( u0_n66 ) );
  OAI21_X1 u0_U169 (.B1( ld ) , .ZN( u0_N260 ) , .B2( u0_n98 ) , .A( u0_n99 ) );
  XNOR2_X1 u0_U17 (.ZN( u0_n53 ) , .B( u0_subword_5 ) , .A( w0_5 ) );
  NAND2_X1 u0_U170 (.A1( key[20] ) , .A2( ld ) , .ZN( u0_n99 ) );
  OAI21_X1 u0_U171 (.B1( ld ) , .ZN( u0_N251 ) , .B2( u0_n125 ) , .A( u0_n126 ) );
  NAND2_X1 u0_U172 (.A1( key[11] ) , .A2( ld ) , .ZN( u0_n126 ) );
  OAI21_X1 u0_U173 (.B1( ld ) , .ZN( u0_N244 ) , .B2( u0_n146 ) , .A( u0_n147 ) );
  NAND2_X1 u0_U174 (.A1( key[4] ) , .A2( ld ) , .ZN( u0_n147 ) );
  OAI21_X1 u0_U175 (.B1( ld ) , .ZN( u0_N115 ) , .B2( u0_n210 ) , .A( u0_n273 ) );
  NAND2_X1 u0_U176 (.A1( key[71] ) , .A2( ld ) , .ZN( u0_n273 ) );
  OAI21_X1 u0_U177 (.B1( ld ) , .ZN( u0_N113 ) , .B2( u0_n214 ) , .A( u0_n277 ) );
  NAND2_X1 u0_U178 (.A1( key[69] ) , .A2( ld ) , .ZN( u0_n277 ) );
  OAI21_X1 u0_U179 (.B1( ld ) , .ZN( u0_N111 ) , .B2( u0_n218 ) , .A( u0_n281 ) );
  XNOR2_X1 u0_U18 (.ZN( u0_n21 ) , .B( u0_subword_21 ) , .A( w0_21 ) );
  NAND2_X1 u0_U180 (.A1( key[67] ) , .A2( ld ) , .ZN( u0_n281 ) );
  XNOR2_X1 u0_U181 (.ZN( u0_n226 ) , .B( u0_subword_31 ) , .A( w0_31 ) );
  OAI21_X1 u0_U182 (.B1( ld ) , .ZN( u0_N42 ) , .B2( u0_n63 ) , .A( u0_n64 ) );
  XNOR2_X1 u0_U183 (.ZN( u0_n61 ) , .B( u0_subword_1 ) , .A( w0_1 ) );
  OAI21_X1 u0_U184 (.B1( ld ) , .ZN( u0_N50 ) , .B2( u0_n47 ) , .A( u0_n48 ) );
  XNOR2_X1 u0_U185 (.ZN( u0_n55 ) , .B( u0_subword_4 ) , .A( w0_4 ) );
  OAI21_X1 u0_U186 (.B1( ld ) , .ZN( u0_N44 ) , .B2( u0_n59 ) , .A( u0_n60 ) );
  OAI21_X1 u0_U187 (.B1( ld ) , .ZN( u0_N59 ) , .B2( u0_n29 ) , .A( u0_n30 ) );
  OAI21_X1 u0_U188 (.B1( ld ) , .ZN( u0_N247 ) , .B2( u0_n137 ) , .A( u0_n138 ) );
  OAI21_X1 u0_U189 (.B1( ld ) , .ZN( u0_N67 ) , .B2( u0_n13 ) , .A( u0_n14 ) );
  NAND2_X1 u0_U19 (.A1( key[22] ) , .A2( ld ) , .ZN( u0_n93 ) );
  OAI21_X1 u0_U190 (.B1( ld ) , .ZN( u0_N252 ) , .B2( u0_n122 ) , .A( u0_n123 ) );
  OAI21_X1 u0_U191 (.B1( ld ) , .ZN( u0_N186 ) , .B2( u0_n124 ) , .A( u0_n199 ) );
  OAI21_X1 u0_U192 (.B1( ld ) , .ZN( u0_N269 ) , .B2( u0_n71 ) , .A( u0_n72 ) );
  OAI21_X1 u0_U193 (.B1( ld ) , .ZN( u0_N73 ) , .B2( u0_n1 ) , .A( u0_n2 ) );
  XNOR2_X1 u0_U194 (.ZN( u0_n15 ) , .A( u0_n240 ) , .B( u0_n246 ) );
  XNOR2_X1 u0_U195 (.B( u0_n248 ) , .ZN( u0_n86 ) , .A( u0_n88 ) );
  OAI21_X1 u0_U196 (.B1( ld ) , .ZN( u0_N254 ) , .B2( u0_n116 ) , .A( u0_n117 ) );
  OAI21_X1 u0_U197 (.B1( ld ) , .ZN( u0_N109 ) , .B2( u0_n222 ) , .A( u0_n285 ) );
  OAI21_X1 u0_U198 (.B1( ld ) , .ZN( u0_N119 ) , .B2( u0_n202 ) , .A( u0_n265 ) );
  OAI21_X1 u0_U199 (.B1( ld ) , .ZN( u0_N185 ) , .B2( u0_n127 ) , .A( u0_n201 ) );
  XNOR2_X1 u0_U20 (.ZN( u0_n25 ) , .B( u0_subword_19 ) , .A( w0_19 ) );
  OAI21_X1 u0_U200 (.B1( ld ) , .ZN( u0_N136 ) , .B2( u0_n168 ) , .A( u0_n231 ) );
  OAI21_X1 u0_U201 (.B1( ld ) , .ZN( u0_N202 ) , .A( u0_n167 ) , .B2( u0_n76 ) );
  XNOR2_X1 u0_U202 (.ZN( u0_n31 ) , .B( u0_subword_16 ) , .A( w0_16 ) );
  INV_X1 u0_U203 (.A( u0_n250 ) , .ZN( w3_13 ) );
  OAI21_X1 u0_U204 (.B1( ld ) , .ZN( u0_N128 ) , .B2( u0_n184 ) , .A( u0_n247 ) );
  OAI21_X1 u0_U205 (.B1( ld ) , .ZN( u0_N194 ) , .B2( u0_n100 ) , .A( u0_n183 ) );
  INV_X1 u0_U206 (.A( u0_n254 ) , .ZN( w3_14 ) );
  OAI21_X1 u0_U207 (.B1( ld ) , .ZN( u0_N245 ) , .B2( u0_n143 ) , .A( u0_n144 ) );
  OAI21_X1 u0_U208 (.B1( ld ) , .ZN( u0_N179 ) , .B2( u0_n145 ) , .A( u0_n213 ) );
  OAI21_X1 u0_U209 (.B1( ld ) , .ZN( u0_N249 ) , .B2( u0_n131 ) , .A( u0_n132 ) );
  XNOR2_X1 u0_U21 (.ZN( u0_n49 ) , .B( u0_subword_7 ) , .A( w0_7 ) );
  INV_X1 u0_U210 (.A( u0_n258 ) , .ZN( w3_12 ) );
  XNOR2_X1 u0_U211 (.ZN( u0_n43 ) , .B( u0_subword_10 ) , .A( w0_10 ) );
  XNOR2_X1 u0_U212 (.ZN( u0_n59 ) , .A( u0_subword_2 ) , .B( w0_2 ) );
  OAI21_X1 u0_U213 (.B1( ld ) , .ZN( u0_N49 ) , .B2( u0_n49 ) , .A( u0_n50 ) );
  OAI21_X1 u0_U214 (.B1( ld ) , .ZN( u0_N125 ) , .B2( u0_n190 ) , .A( u0_n253 ) );
  XNOR2_X1 u0_U215 (.ZN( u0_n164 ) , .B( u0_n262 ) , .A( u0_n3 ) );
  OAI21_X1 u0_U216 (.B1( ld ) , .ZN( u0_N262 ) , .B2( u0_n92 ) , .A( u0_n93 ) );
  XNOR2_X1 u0_U217 (.ZN( u0_n27 ) , .B( u0_subword_18 ) , .A( w0_18 ) );
  OAI21_X1 u0_U218 (.B1( ld ) , .ZN( u0_N139 ) , .B2( u0_n162 ) , .A( u0_n225 ) );
  OAI21_X1 u0_U219 (.B1( ld ) , .ZN( u0_N205 ) , .A( u0_n161 ) , .B2( u0_n67 ) );
  XNOR2_X1 u0_U22 (.ZN( u0_n29 ) , .B( u0_subword_17 ) , .A( w0_17 ) );
  OAI21_X1 u0_U220 (.B1( ld ) , .ZN( u0_N112 ) , .B2( u0_n216 ) , .A( u0_n279 ) );
  OAI21_X1 u0_U221 (.B1( ld ) , .ZN( u0_N178 ) , .B2( u0_n148 ) , .A( u0_n215 ) );
  OAI21_X1 u0_U222 (.B1( ld ) , .ZN( u0_N246 ) , .B2( u0_n140 ) , .A( u0_n141 ) );
  OAI21_X1 u0_U223 (.B1( ld ) , .ZN( u0_N243 ) , .B2( u0_n149 ) , .A( u0_n150 ) );
  OAI21_X1 u0_U224 (.B1( ld ) , .ZN( u0_N177 ) , .B2( u0_n151 ) , .A( u0_n217 ) );
  OAI21_X1 u0_U225 (.B1( ld ) , .ZN( u0_N133 ) , .B2( u0_n174 ) , .A( u0_n237 ) );
  OAI21_X1 u0_U226 (.B1( ld ) , .ZN( u0_N259 ) , .B2( u0_n101 ) , .A( u0_n102 ) );
  OAI21_X1 u0_U227 (.B1( ld ) , .ZN( u0_N61 ) , .B2( u0_n25 ) , .A( u0_n26 ) );
  OAI21_X1 u0_U228 (.B1( ld ) , .ZN( u0_N255 ) , .B2( u0_n113 ) , .A( u0_n114 ) );
  OAI21_X1 u0_U229 (.B1( ld ) , .ZN( u0_N189 ) , .B2( u0_n115 ) , .A( u0_n193 ) );
  XNOR2_X1 u0_U23 (.ZN( u0_n39 ) , .B( u0_subword_12 ) , .A( w0_12 ) );
  INV_X1 u0_U230 (.A( u0_n264 ) , .ZN( w3_15 ) );
  OAI21_X1 u0_U231 (.B1( ld ) , .ZN( u0_N263 ) , .B2( u0_n89 ) , .A( u0_n90 ) );
  OAI21_X1 u0_U232 (.B1( ld ) , .ZN( u0_N197 ) , .A( u0_n177 ) , .B2( u0_n91 ) );
  OAI21_X1 u0_U233 (.B1( ld ) , .ZN( u0_N117 ) , .B2( u0_n206 ) , .A( u0_n269 ) );
  OAI21_X1 u0_U234 (.B1( ld ) , .ZN( u0_N183 ) , .B2( u0_n133 ) , .A( u0_n205 ) );
  XNOR2_X1 u0_U235 (.ZN( u0_n47 ) , .B( u0_subword_8 ) , .A( w0_8 ) );
  OAI21_X1 u0_U236 (.B1( ld ) , .ZN( u0_N127 ) , .B2( u0_n186 ) , .A( u0_n249 ) );
  OAI21_X1 u0_U237 (.B1( ld ) , .ZN( u0_N193 ) , .B2( u0_n103 ) , .A( u0_n185 ) );
  OAI21_X1 u0_U238 (.B1( ld ) , .ZN( u0_N241 ) , .B2( u0_n155 ) , .A( u0_n156 ) );
  OAI21_X1 u0_U239 (.B1( ld ) , .ZN( u0_N175 ) , .B2( u0_n157 ) , .A( u0_n221 ) );
  NAND2_X1 u0_U24 (.A1( key[47] ) , .A2( ld ) , .ZN( u0_n193 ) );
  XNOR2_X1 u0_U240 (.ZN( u0_n35 ) , .B( u0_subword_14 ) , .A( w0_14 ) );
  OAI21_X1 u0_U241 (.B1( ld ) , .ZN( u0_N257 ) , .B2( u0_n107 ) , .A( u0_n108 ) );
  OAI21_X1 u0_U242 (.B1( ld ) , .ZN( u0_N191 ) , .B2( u0_n109 ) , .A( u0_n189 ) );
  OAI21_X1 u0_U243 (.B1( ld ) , .ZN( u0_N48 ) , .B2( u0_n51 ) , .A( u0_n52 ) );
  OAI21_X1 u0_U244 (.B1( ld ) , .ZN( u0_N116 ) , .B2( u0_n208 ) , .A( u0_n271 ) );
  OAI21_X1 u0_U245 (.B1( ld ) , .ZN( u0_N264 ) , .B2( u0_n86 ) , .A( u0_n87 ) );
  OAI21_X1 u0_U246 (.B1( ld ) , .ZN( u0_N66 ) , .B2( u0_n15 ) , .A( u0_n16 ) );
  OAI21_X1 u0_U247 (.B1( ld ) , .ZN( u0_N64 ) , .B2( u0_n19 ) , .A( u0_n20 ) );
  XNOR2_X1 u0_U248 (.ZN( u0_n63 ) , .B( u0_subword_0 ) , .A( w0_0 ) );
  OAI21_X1 u0_U249 (.B1( ld ) , .ZN( u0_N265 ) , .B2( u0_n83 ) , .A( u0_n84 ) );
  NAND2_X1 u0_U25 (.A1( key[55] ) , .A2( ld ) , .ZN( u0_n177 ) );
  OAI21_X1 u0_U250 (.B1( ld ) , .ZN( u0_N199 ) , .A( u0_n173 ) , .B2( u0_n85 ) );
  OAI21_X1 u0_U251 (.B1( ld ) , .ZN( u0_N108 ) , .B2( u0_n224 ) , .A( u0_n287 ) );
  OAI21_X1 u0_U252 (.B1( ld ) , .ZN( u0_N256 ) , .B2( u0_n110 ) , .A( u0_n111 ) );
  OAI21_X1 u0_U253 (.B1( ld ) , .ZN( u0_N58 ) , .B2( u0_n31 ) , .A( u0_n32 ) );
  XNOR2_X1 u0_U254 (.ZN( u0_n240 ) , .B( u0_subword_24 ) , .A( w0_24 ) );
  OAI21_X1 u0_U255 (.B1( ld ) , .ZN( u0_N267 ) , .B2( u0_n77 ) , .A( u0_n78 ) );
  OAI21_X1 u0_U256 (.B1( ld ) , .ZN( u0_N201 ) , .A( u0_n169 ) , .B2( u0_n79 ) );
  OAI21_X1 u0_U257 (.B1( ld ) , .ZN( u0_N72 ) , .B2( u0_n3 ) , .A( u0_n4 ) );
  OAI21_X1 u0_U258 (.B1( ld ) , .ZN( u0_N138 ) , .B2( u0_n164 ) , .A( u0_n227 ) );
  XNOR2_X1 u0_U259 (.ZN( u0_n51 ) , .B( u0_subword_6 ) , .A( w0_6 ) );
  NAND2_X1 u0_U26 (.A1( key[37] ) , .A2( ld ) , .ZN( u0_n213 ) );
  XNOR2_X1 u0_U260 (.ZN( u0_n230 ) , .B( u0_subword_29 ) , .A( w0_29 ) );
  OAI21_X1 u0_U261 (.B1( ld ) , .ZN( u0_N56 ) , .B2( u0_n35 ) , .A( u0_n36 ) );
  XNOR2_X1 u0_U262 (.ZN( u0_n19 ) , .B( u0_subword_22 ) , .A( w0_22 ) );
  OAI21_X1 u0_U263 (.B1( ld ) , .ZN( u0_N261 ) , .B2( u0_n95 ) , .A( u0_n96 ) );
  OAI21_X1 u0_U264 (.B1( ld ) , .ZN( u0_N195 ) , .A( u0_n181 ) , .B2( u0_n97 ) );
  OAI21_X1 u0_U265 (.B1( ld ) , .ZN( u0_N137 ) , .B2( u0_n166 ) , .A( u0_n229 ) );
  OAI21_X1 u0_U266 (.B1( ld ) , .ZN( u0_N203 ) , .A( u0_n165 ) , .B2( u0_n73 ) );
  OAI21_X1 u0_U267 (.B1( ld ) , .ZN( u0_N266 ) , .B2( u0_n80 ) , .A( u0_n81 ) );
  OAI21_X1 u0_U268 (.B1( ld ) , .ZN( u0_N114 ) , .B2( u0_n212 ) , .A( u0_n275 ) );
  OAI21_X1 u0_U269 (.B1( ld ) , .ZN( u0_N180 ) , .B2( u0_n142 ) , .A( u0_n211 ) );
  NAND2_X1 u0_U27 (.A1( key[35] ) , .A2( ld ) , .ZN( u0_n217 ) );
  OAI21_X1 u0_U270 (.B1( ld ) , .ZN( u0_N130 ) , .B2( u0_n180 ) , .A( u0_n243 ) );
  OAI21_X1 u0_U271 (.B1( ld ) , .ZN( u0_N196 ) , .A( u0_n179 ) , .B2( u0_n94 ) );
  OAI21_X1 u0_U272 (.B1( ld ) , .ZN( u0_N242 ) , .B2( u0_n152 ) , .A( u0_n153 ) );
  OAI21_X1 u0_U273 (.B1( ld ) , .ZN( u0_N122 ) , .B2( u0_n196 ) , .A( u0_n259 ) );
  OAI21_X1 u0_U274 (.B1( ld ) , .ZN( u0_N188 ) , .B2( u0_n118 ) , .A( u0_n195 ) );
  OAI21_X1 u0_U275 (.B1( ld ) , .ZN( u0_N253 ) , .B2( u0_n119 ) , .A( u0_n120 ) );
  OAI21_X1 u0_U276 (.B1( ld ) , .ZN( u0_N187 ) , .B2( u0_n121 ) , .A( u0_n197 ) );
  OAI21_X1 u0_U277 (.B1( ld ) , .ZN( u0_N270 ) , .B2( u0_n68 ) , .A( u0_n69 ) );
  OAI21_X1 u0_U278 (.B1( ld ) , .ZN( u0_N204 ) , .A( u0_n163 ) , .B2( u0_n70 ) );
  OAI21_X1 u0_U279 (.B1( ld ) , .ZN( u0_N124 ) , .B2( u0_n192 ) , .A( u0_n255 ) );
  NAND2_X1 u0_U28 (.A1( key[93] ) , .A2( ld ) , .ZN( u0_n229 ) );
  OAI21_X1 u0_U280 (.B1( ld ) , .ZN( u0_N190 ) , .B2( u0_n112 ) , .A( u0_n191 ) );
  OAI21_X1 u0_U281 (.B1( ld ) , .ZN( u0_N248 ) , .B2( u0_n134 ) , .A( u0_n135 ) );
  OAI21_X1 u0_U282 (.B1( ld ) , .ZN( u0_N182 ) , .B2( u0_n136 ) , .A( u0_n207 ) );
  OAI21_X1 u0_U283 (.B1( ld ) , .ZN( u0_N132 ) , .B2( u0_n176 ) , .A( u0_n239 ) );
  OAI21_X1 u0_U284 (.B1( ld ) , .ZN( u0_N198 ) , .A( u0_n175 ) , .B2( u0_n88 ) );
  OAI21_X1 u0_U285 (.B1( ld ) , .ZN( u0_N240 ) , .B2( u0_n158 ) , .A( u0_n159 ) );
  OAI21_X1 u0_U286 (.B1( ld ) , .ZN( u0_N174 ) , .B2( u0_n160 ) , .A( u0_n223 ) );
  XNOR2_X1 u0_U287 (.ZN( u0_n236 ) , .A( u0_subword_26 ) , .B( w0_26 ) );
  OAI21_X1 u0_U288 (.B1( ld ) , .ZN( u0_N52 ) , .B2( u0_n43 ) , .A( u0_n44 ) );
  OAI21_X1 u0_U289 (.B1( ld ) , .ZN( u0_N118 ) , .B2( u0_n204 ) , .A( u0_n267 ) );
  NAND2_X1 u0_U29 (.A1( key[92] ) , .A2( ld ) , .ZN( u0_n231 ) );
  OAI21_X1 u0_U290 (.B1( ld ) , .ZN( u0_N60 ) , .B2( u0_n27 ) , .A( u0_n28 ) );
  XOR2_X1 u0_U291 (.Z( u0_n65 ) , .A( u0_n67 ) , .B( w3_31 ) );
  XOR2_X1 u0_U292 (.Z( u0_n68 ) , .A( u0_n70 ) , .B( w3_30 ) );
  XOR2_X1 u0_U293 (.Z( u0_n71 ) , .A( u0_n73 ) , .B( w3_29 ) );
  XOR2_X1 u0_U294 (.Z( u0_n74 ) , .A( u0_n76 ) , .B( w3_28 ) );
  XOR2_X1 u0_U295 (.Z( u0_n77 ) , .A( u0_n79 ) , .B( w3_27 ) );
  XOR2_X1 u0_U296 (.Z( u0_n80 ) , .A( u0_n82 ) , .B( w3_26 ) );
  XOR2_X1 u0_U297 (.Z( u0_n83 ) , .A( u0_n85 ) , .B( w3_25 ) );
  OAI21_X1 u0_U298 (.B1( ld ) , .ZN( u0_N126 ) , .B2( u0_n188 ) , .A( u0_n251 ) );
  XOR2_X1 u0_U299 (.Z( u0_n89 ) , .A( u0_n91 ) , .B( w3_23 ) );
  XNOR2_X1 u0_U3 (.A( u0_n11 ) , .ZN( u0_n172 ) , .B( u0_n242 ) );
  NAND2_X1 u0_U30 (.A1( key[59] ) , .A2( ld ) , .ZN( u0_n169 ) );
  XOR2_X1 u0_U300 (.Z( u0_n92 ) , .A( u0_n94 ) , .B( w3_22 ) );
  XOR2_X1 u0_U301 (.Z( u0_n95 ) , .A( u0_n97 ) , .B( w3_21 ) );
  XOR2_X1 u0_U302 (.A( u0_n100 ) , .Z( u0_n98 ) , .B( w3_20 ) );
  XOR2_X1 u0_U303 (.Z( u0_n101 ) , .A( u0_n103 ) , .B( w3_19 ) );
  XOR2_X1 u0_U304 (.Z( u0_n104 ) , .A( u0_n106 ) , .B( w3_18 ) );
  XOR2_X1 u0_U305 (.Z( u0_n107 ) , .A( u0_n109 ) , .B( w3_17 ) );
  XOR2_X1 u0_U306 (.Z( u0_n110 ) , .A( u0_n112 ) , .B( w3_16 ) );
  XOR2_X1 u0_U307 (.Z( u0_n113 ) , .A( u0_n115 ) , .B( w3_15 ) );
  XOR2_X1 u0_U308 (.Z( u0_n116 ) , .A( u0_n118 ) , .B( w3_14 ) );
  XOR2_X1 u0_U309 (.Z( u0_n119 ) , .A( u0_n121 ) , .B( w3_13 ) );
  NAND2_X1 u0_U31 (.A1( key[53] ) , .A2( ld ) , .ZN( u0_n181 ) );
  XOR2_X1 u0_U310 (.Z( u0_n122 ) , .A( u0_n124 ) , .B( w3_12 ) );
  XOR2_X1 u0_U311 (.Z( u0_n125 ) , .A( u0_n127 ) , .B( w3_11 ) );
  XOR2_X1 u0_U312 (.Z( u0_n128 ) , .A( u0_n130 ) , .B( w3_10 ) );
  XOR2_X1 u0_U313 (.Z( u0_n131 ) , .A( u0_n133 ) , .B( w3_9 ) );
  XOR2_X1 u0_U314 (.Z( u0_n134 ) , .A( u0_n136 ) , .B( w3_8 ) );
  XOR2_X1 u0_U315 (.Z( u0_n137 ) , .A( u0_n139 ) , .B( w3_7 ) );
  XOR2_X1 u0_U316 (.Z( u0_n140 ) , .A( u0_n142 ) , .B( w3_6 ) );
  XOR2_X1 u0_U317 (.Z( u0_n143 ) , .A( u0_n145 ) , .B( w3_5 ) );
  XOR2_X1 u0_U318 (.Z( u0_n146 ) , .A( u0_n148 ) , .B( w3_4 ) );
  XOR2_X1 u0_U319 (.Z( u0_n149 ) , .A( u0_n151 ) , .B( w3_3 ) );
  NAND2_X1 u0_U32 (.A1( key[45] ) , .A2( ld ) , .ZN( u0_n197 ) );
  XOR2_X1 u0_U320 (.Z( u0_n152 ) , .A( u0_n154 ) , .B( w3_2 ) );
  XOR2_X1 u0_U321 (.Z( u0_n155 ) , .A( u0_n157 ) , .B( w3_1 ) );
  XOR2_X1 u0_U322 (.Z( u0_n158 ) , .A( u0_n160 ) , .B( w3_0 ) );
  XOR2_X1 u0_U323 (.A( u0_n162 ) , .Z( u0_n67 ) , .B( w2_31 ) );
  XOR2_X1 u0_U324 (.A( u0_n164 ) , .Z( u0_n70 ) , .B( w2_30 ) );
  XOR2_X1 u0_U325 (.A( u0_n166 ) , .Z( u0_n73 ) , .B( w2_29 ) );
  XOR2_X1 u0_U326 (.A( u0_n168 ) , .Z( u0_n76 ) , .B( w2_28 ) );
  XOR2_X1 u0_U327 (.A( u0_n170 ) , .Z( u0_n79 ) , .B( w2_27 ) );
  OAI21_X1 u0_U328 (.B1( ld ) , .ZN( u0_N68 ) , .B2( u0_n11 ) , .A( u0_n12 ) );
  XOR2_X1 u0_U329 (.A( u0_n174 ) , .Z( u0_n85 ) , .B( w2_25 ) );
  NAND2_X1 u0_U33 (.A1( key[44] ) , .A2( ld ) , .ZN( u0_n199 ) );
  XOR2_X1 u0_U330 (.A( u0_n176 ) , .Z( u0_n88 ) , .B( w2_24 ) );
  XOR2_X1 u0_U331 (.A( u0_n178 ) , .Z( u0_n91 ) , .B( w2_23 ) );
  XOR2_X1 u0_U332 (.A( u0_n180 ) , .Z( u0_n94 ) , .B( w2_22 ) );
  XOR2_X1 u0_U333 (.A( u0_n182 ) , .Z( u0_n97 ) , .B( w2_21 ) );
  XOR2_X1 u0_U334 (.Z( u0_n100 ) , .A( u0_n184 ) , .B( w2_20 ) );
  XOR2_X1 u0_U335 (.Z( u0_n103 ) , .A( u0_n186 ) , .B( w2_19 ) );
  XOR2_X1 u0_U336 (.Z( u0_n106 ) , .A( u0_n188 ) , .B( w2_18 ) );
  XOR2_X1 u0_U337 (.Z( u0_n109 ) , .A( u0_n190 ) , .B( w2_17 ) );
  XOR2_X1 u0_U338 (.Z( u0_n112 ) , .A( u0_n192 ) , .B( w2_16 ) );
  XOR2_X1 u0_U339 (.Z( u0_n115 ) , .A( u0_n194 ) , .B( w2_15 ) );
  NAND2_X1 u0_U34 (.A1( key[65] ) , .A2( ld ) , .ZN( u0_n285 ) );
  XOR2_X1 u0_U340 (.Z( u0_n118 ) , .A( u0_n196 ) , .B( w2_14 ) );
  XOR2_X1 u0_U341 (.Z( u0_n121 ) , .A( u0_n198 ) , .B( w2_13 ) );
  XOR2_X1 u0_U342 (.Z( u0_n124 ) , .A( u0_n200 ) , .B( w2_12 ) );
  XOR2_X1 u0_U343 (.Z( u0_n127 ) , .A( u0_n202 ) , .B( w2_11 ) );
  XOR2_X1 u0_U344 (.Z( u0_n130 ) , .A( u0_n204 ) , .B( w2_10 ) );
  XOR2_X1 u0_U345 (.Z( u0_n133 ) , .A( u0_n206 ) , .B( w2_9 ) );
  XOR2_X1 u0_U346 (.Z( u0_n136 ) , .A( u0_n208 ) , .B( w2_8 ) );
  XOR2_X1 u0_U347 (.Z( u0_n139 ) , .A( u0_n210 ) , .B( w2_7 ) );
  XOR2_X1 u0_U348 (.Z( u0_n142 ) , .A( u0_n212 ) , .B( w2_6 ) );
  XOR2_X1 u0_U349 (.Z( u0_n145 ) , .A( u0_n214 ) , .B( w2_5 ) );
  NAND2_X1 u0_U35 (.A1( key[68] ) , .A2( ld ) , .ZN( u0_n279 ) );
  XOR2_X1 u0_U350 (.Z( u0_n148 ) , .A( u0_n216 ) , .B( w2_4 ) );
  XOR2_X1 u0_U351 (.Z( u0_n151 ) , .A( u0_n218 ) , .B( w2_3 ) );
  XOR2_X1 u0_U352 (.Z( u0_n154 ) , .A( u0_n220 ) , .B( w2_2 ) );
  XOR2_X1 u0_U353 (.Z( u0_n157 ) , .A( u0_n222 ) , .B( w2_1 ) );
  XOR2_X1 u0_U354 (.Z( u0_n160 ) , .A( u0_n224 ) , .B( w2_0 ) );
  XOR2_X1 u0_U355 (.A( u0_n1 ) , .Z( u0_n162 ) , .B( w1_31 ) );
  XOR2_X1 u0_U356 (.Z( u0_n1 ) , .A( u0_n226 ) , .B( u0_rcon_31 ) );
  OAI21_X1 u0_U357 (.B1( ld ) , .ZN( u0_N258 ) , .B2( u0_n104 ) , .A( u0_n105 ) );
  XOR2_X1 u0_U358 (.A( u0_n228 ) , .Z( u0_n3 ) , .B( u0_rcon_30 ) );
  XOR2_X1 u0_U359 (.Z( u0_n166 ) , .A( u0_n5 ) , .B( w1_29 ) );
  NAND2_X1 u0_U36 (.A1( key[103] ) , .A2( ld ) , .ZN( u0_n50 ) );
  XOR2_X1 u0_U360 (.A( u0_n230 ) , .Z( u0_n5 ) , .B( u0_rcon_29 ) );
  XOR2_X1 u0_U361 (.Z( u0_n168 ) , .A( u0_n7 ) , .B( w1_28 ) );
  XOR2_X1 u0_U362 (.A( u0_n232 ) , .Z( u0_n7 ) , .B( u0_rcon_28 ) );
  XOR2_X1 u0_U363 (.Z( u0_n170 ) , .A( u0_n9 ) , .B( w1_27 ) );
  XOR2_X1 u0_U364 (.A( u0_n234 ) , .Z( u0_n9 ) , .B( u0_rcon_27 ) );
  OAI21_X1 u0_U365 (.B1( ld ) , .ZN( u0_N192 ) , .B2( u0_n106 ) , .A( u0_n187 ) );
  XOR2_X1 u0_U366 (.Z( u0_n11 ) , .A( u0_n236 ) , .B( u0_rcon_26 ) );
  XOR2_X1 u0_U367 (.A( u0_n13 ) , .Z( u0_n174 ) , .B( w1_25 ) );
  XOR2_X1 u0_U368 (.Z( u0_n13 ) , .A( u0_n238 ) , .B( u0_rcon_25 ) );
  XOR2_X1 u0_U369 (.A( u0_n15 ) , .Z( u0_n176 ) , .B( w1_24 ) );
  NAND2_X1 u0_U37 (.A1( key[102] ) , .A2( ld ) , .ZN( u0_n52 ) );
  OAI21_X1 u0_U370 (.B1( ld ) , .ZN( u0_N110 ) , .B2( u0_n220 ) , .A( u0_n283 ) );
  XOR2_X1 u0_U371 (.A( u0_n17 ) , .Z( u0_n178 ) , .B( w1_23 ) );
  OAI21_X1 u0_U372 (.B1( ld ) , .ZN( u0_N176 ) , .B2( u0_n154 ) , .A( u0_n219 ) );
  XOR2_X1 u0_U373 (.Z( u0_n180 ) , .A( u0_n19 ) , .B( w1_22 ) );
  OAI21_X1 u0_U374 (.B1( ld ) , .ZN( u0_N250 ) , .B2( u0_n128 ) , .A( u0_n129 ) );
  XOR2_X1 u0_U375 (.Z( u0_n182 ) , .A( u0_n21 ) , .B( w1_21 ) );
  OAI21_X1 u0_U376 (.B1( ld ) , .ZN( u0_N184 ) , .B2( u0_n130 ) , .A( u0_n203 ) );
  XOR2_X1 u0_U377 (.Z( u0_n184 ) , .A( u0_n23 ) , .B( w1_20 ) );
  OAI21_X1 u0_U378 (.B1( ld ) , .ZN( u0_N134 ) , .B2( u0_n172 ) , .A( u0_n235 ) );
  XOR2_X1 u0_U379 (.Z( u0_n186 ) , .A( u0_n25 ) , .B( w1_19 ) );
  NAND2_X1 u0_U38 (.A1( key[96] ) , .A2( ld ) , .ZN( u0_n64 ) );
  OAI21_X1 u0_U380 (.B1( ld ) , .ZN( u0_N200 ) , .A( u0_n171 ) , .B2( u0_n82 ) );
  XOR2_X1 u0_U381 (.Z( u0_n188 ) , .A( u0_n27 ) , .B( w1_18 ) );
  XOR2_X1 u0_U383 (.Z( u0_n190 ) , .A( u0_n29 ) , .B( w1_17 ) );
  XOR2_X1 u0_U385 (.Z( u0_n192 ) , .A( u0_n31 ) , .B( w1_16 ) );
  XOR2_X1 u0_U387 (.Z( u0_n194 ) , .A( u0_n33 ) , .B( w1_15 ) );
  XOR2_X1 u0_U389 (.Z( u0_n196 ) , .A( u0_n35 ) , .B( w1_14 ) );
  NAND2_X1 u0_U39 (.A1( key[115] ) , .A2( ld ) , .ZN( u0_n26 ) );
  XOR2_X1 u0_U391 (.Z( u0_n198 ) , .A( u0_n37 ) , .B( w1_13 ) );
  XOR2_X1 u0_U393 (.Z( u0_n200 ) , .A( u0_n39 ) , .B( w1_12 ) );
  XOR2_X1 u0_U395 (.Z( u0_n202 ) , .A( u0_n41 ) , .B( w1_11 ) );
  XOR2_X1 u0_U397 (.Z( u0_n204 ) , .A( u0_n43 ) , .B( w1_10 ) );
  XOR2_X1 u0_U399 (.Z( u0_n206 ) , .A( u0_n45 ) , .B( w1_9 ) );
  XNOR2_X1 u0_U4 (.A( u0_n172 ) , .B( u0_n244 ) , .ZN( u0_n82 ) );
  NAND2_X1 u0_U40 (.A1( key[114] ) , .A2( ld ) , .ZN( u0_n28 ) );
  XOR2_X1 u0_U401 (.Z( u0_n208 ) , .A( u0_n47 ) , .B( w1_8 ) );
  XOR2_X1 u0_U403 (.Z( u0_n210 ) , .A( u0_n49 ) , .B( w1_7 ) );
  XOR2_X1 u0_U405 (.Z( u0_n212 ) , .A( u0_n51 ) , .B( w1_6 ) );
  XOR2_X1 u0_U407 (.Z( u0_n214 ) , .A( u0_n53 ) , .B( w1_5 ) );
  XOR2_X1 u0_U409 (.Z( u0_n216 ) , .A( u0_n55 ) , .B( w1_4 ) );
  NAND2_X1 u0_U41 (.A1( key[112] ) , .A2( ld ) , .ZN( u0_n32 ) );
  XOR2_X1 u0_U411 (.Z( u0_n218 ) , .A( u0_n57 ) , .B( w1_3 ) );
  XOR2_X1 u0_U413 (.Z( u0_n220 ) , .A( u0_n59 ) , .B( w1_2 ) );
  XOR2_X1 u0_U415 (.Z( u0_n222 ) , .A( u0_n61 ) , .B( w1_1 ) );
  XOR2_X1 u0_U417 (.Z( u0_n224 ) , .A( u0_n63 ) , .B( w1_0 ) );
  NAND2_X1 u0_U42 (.A1( key[106] ) , .A2( ld ) , .ZN( u0_n44 ) );
  NAND2_X1 u0_U43 (.A1( key[64] ) , .A2( ld ) , .ZN( u0_n287 ) );
  NAND2_X1 u0_U44 (.A1( key[126] ) , .A2( ld ) , .ZN( u0_n4 ) );
  NAND2_X1 u0_U45 (.A1( key[23] ) , .A2( ld ) , .ZN( u0_n90 ) );
  NAND2_X1 u0_U46 (.A1( key[21] ) , .A2( ld ) , .ZN( u0_n96 ) );
  NAND2_X1 u0_U47 (.A1( key[24] ) , .A2( ld ) , .ZN( u0_n87 ) );
  NAND2_X1 u0_U48 (.A1( key[25] ) , .A2( ld ) , .ZN( u0_n84 ) );
  NAND2_X1 u0_U49 (.A1( key[122] ) , .A2( ld ) , .ZN( u0_n12 ) );
  XNOR2_X1 u0_U5 (.ZN( u0_n232 ) , .B( u0_subword_28 ) , .A( w0_28 ) );
  NAND2_X1 u0_U50 (.A1( key[118] ) , .A2( ld ) , .ZN( u0_n20 ) );
  NAND2_X1 u0_U51 (.A1( key[89] ) , .A2( ld ) , .ZN( u0_n237 ) );
  NAND2_X1 u0_U52 (.A1( key[120] ) , .A2( ld ) , .ZN( u0_n16 ) );
  NAND2_X1 u0_U53 (.A1( key[88] ) , .A2( ld ) , .ZN( u0_n239 ) );
  NAND2_X1 u0_U54 (.A1( key[86] ) , .A2( ld ) , .ZN( u0_n243 ) );
  NAND2_X1 u0_U55 (.A1( key[82] ) , .A2( ld ) , .ZN( u0_n251 ) );
  NAND2_X1 u0_U56 (.A1( key[80] ) , .A2( ld ) , .ZN( u0_n255 ) );
  NAND2_X1 u0_U57 (.A1( key[78] ) , .A2( ld ) , .ZN( u0_n259 ) );
  NAND2_X1 u0_U58 (.A1( key[26] ) , .A2( ld ) , .ZN( u0_n81 ) );
  NAND2_X1 u0_U59 (.A1( key[27] ) , .A2( ld ) , .ZN( u0_n78 ) );
  XNOR2_X1 u0_U6 (.ZN( u0_n234 ) , .B( u0_subword_27 ) , .A( w0_27 ) );
  NAND2_X1 u0_U60 (.A1( key[98] ) , .A2( ld ) , .ZN( u0_n60 ) );
  NAND2_X1 u0_U61 (.A1( key[121] ) , .A2( ld ) , .ZN( u0_n14 ) );
  NAND2_X1 u0_U62 (.A1( key[84] ) , .A2( ld ) , .ZN( u0_n247 ) );
  NAND2_X1 u0_U63 (.A1( key[83] ) , .A2( ld ) , .ZN( u0_n249 ) );
  NAND2_X1 u0_U64 (.A1( key[113] ) , .A2( ld ) , .ZN( u0_n30 ) );
  NAND2_X1 u0_U65 (.A1( key[81] ) , .A2( ld ) , .ZN( u0_n253 ) );
  NAND2_X1 u0_U66 (.A1( key[110] ) , .A2( ld ) , .ZN( u0_n36 ) );
  NAND2_X1 u0_U67 (.A1( key[75] ) , .A2( ld ) , .ZN( u0_n265 ) );
  NAND2_X1 u0_U68 (.A1( key[104] ) , .A2( ld ) , .ZN( u0_n48 ) );
  NAND2_X1 u0_U69 (.A1( key[95] ) , .A2( ld ) , .ZN( u0_n225 ) );
  XNOR2_X1 u0_U7 (.ZN( u0_n228 ) , .B( u0_subword_30 ) , .A( w0_30 ) );
  NAND2_X1 u0_U70 (.A1( key[63] ) , .A2( ld ) , .ZN( u0_n161 ) );
  NAND2_X1 u0_U71 (.A1( key[38] ) , .A2( ld ) , .ZN( u0_n211 ) );
  NAND2_X1 u0_U72 (.A1( key[36] ) , .A2( ld ) , .ZN( u0_n215 ) );
  NAND2_X1 u0_U73 (.A1( key[34] ) , .A2( ld ) , .ZN( u0_n219 ) );
  NAND2_X1 u0_U74 (.A1( key[33] ) , .A2( ld ) , .ZN( u0_n221 ) );
  NAND2_X1 u0_U75 (.A1( key[32] ) , .A2( ld ) , .ZN( u0_n223 ) );
  NAND2_X1 u0_U76 (.A1( key[94] ) , .A2( ld ) , .ZN( u0_n227 ) );
  NAND2_X1 u0_U77 (.A1( key[61] ) , .A2( ld ) , .ZN( u0_n165 ) );
  NAND2_X1 u0_U78 (.A1( key[60] ) , .A2( ld ) , .ZN( u0_n167 ) );
  NAND2_X1 u0_U79 (.A1( key[90] ) , .A2( ld ) , .ZN( u0_n235 ) );
  XNOR2_X1 u0_U8 (.ZN( u0_n238 ) , .B( u0_subword_25 ) , .A( w0_25 ) );
  NAND2_X1 u0_U80 (.A1( key[58] ) , .A2( ld ) , .ZN( u0_n171 ) );
  NAND2_X1 u0_U81 (.A1( key[57] ) , .A2( ld ) , .ZN( u0_n173 ) );
  NAND2_X1 u0_U82 (.A1( key[56] ) , .A2( ld ) , .ZN( u0_n175 ) );
  NAND2_X1 u0_U83 (.A1( key[54] ) , .A2( ld ) , .ZN( u0_n179 ) );
  NAND2_X1 u0_U84 (.A1( key[52] ) , .A2( ld ) , .ZN( u0_n183 ) );
  NAND2_X1 u0_U85 (.A1( key[51] ) , .A2( ld ) , .ZN( u0_n185 ) );
  NAND2_X1 u0_U86 (.A1( key[50] ) , .A2( ld ) , .ZN( u0_n187 ) );
  NAND2_X1 u0_U87 (.A1( key[49] ) , .A2( ld ) , .ZN( u0_n189 ) );
  NAND2_X1 u0_U88 (.A1( key[48] ) , .A2( ld ) , .ZN( u0_n191 ) );
  NAND2_X1 u0_U89 (.A1( key[46] ) , .A2( ld ) , .ZN( u0_n195 ) );
  INV_X1 u0_U9 (.ZN( u0_n246 ) , .A( u0_rcon_24 ) );
  NAND2_X1 u0_U90 (.A1( key[43] ) , .A2( ld ) , .ZN( u0_n201 ) );
  NAND2_X1 u0_U91 (.A1( key[42] ) , .A2( ld ) , .ZN( u0_n203 ) );
  NAND2_X1 u0_U92 (.A1( key[41] ) , .A2( ld ) , .ZN( u0_n205 ) );
  NAND2_X1 u0_U93 (.A1( key[40] ) , .A2( ld ) , .ZN( u0_n207 ) );
  NAND2_X1 u0_U94 (.A1( key[13] ) , .A2( ld ) , .ZN( u0_n120 ) );
  NAND2_X1 u0_U95 (.A1( key[14] ) , .A2( ld ) , .ZN( u0_n117 ) );
  NAND2_X1 u0_U96 (.A1( key[12] ) , .A2( ld ) , .ZN( u0_n123 ) );
  NAND2_X1 u0_U97 (.A1( key[7] ) , .A2( ld ) , .ZN( u0_n138 ) );
  NAND2_X1 u0_U98 (.A1( key[70] ) , .A2( ld ) , .ZN( u0_n275 ) );
  NAND2_X1 u0_U99 (.A1( key[66] ) , .A2( ld ) , .ZN( u0_n283 ) );
  OAI21_X1 u0_r0_U27 (.ZN( u0_r0_N70 ) , .B1( u0_r0_n4 ) , .B2( u0_r0_n5 ) , .A( u0_r0_n9 ) );
  NAND4_X1 u0_r0_U28 (.A3( u0_r0_N78 ) , .A2( u0_r0_n12 ) , .ZN( u0_r0_n14 ) , .A1( u0_r0_n18 ) , .A4( u0_r0_n2 ) );
  NAND2_X1 u0_r0_U29 (.A1( u0_r0_N80 ) , .ZN( u0_r0_n11 ) , .A2( u0_r0_n17 ) );
  NOR2_X1 u0_r0_U30 (.A2( ld ) , .ZN( u0_r0_N79 ) , .A1( u0_r0_n12 ) );
  NOR2_X1 u0_r0_U31 (.A2( ld ) , .ZN( u0_r0_N80 ) , .A1( u0_r0_n18 ) );
  NAND2_X1 u0_r0_U32 (.ZN( u0_r0_N71 ) , .A1( u0_r0_n10 ) , .A2( u0_r0_n23 ) );
  INV_X1 u0_r0_U33 (.A( u0_r0_n17 ) , .ZN( u0_r0_n2 ) );
  INV_X1 u0_r0_U34 (.A( u0_r0_n24 ) , .ZN( u0_r0_n5 ) );
  INV_X1 u0_r0_U35 (.A( u0_r0_n25 ) , .ZN( u0_r0_n4 ) );
  XNOR2_X1 u0_r0_U36 (.ZN( u0_r0_n12 ) , .B( u0_r0_rcnt_0 ) , .A( u0_r0_rcnt_1 ) );
  OAI21_X1 u0_r0_U37 (.B1( u0_r0_n12 ) , .A( u0_r0_n21 ) , .ZN( u0_r0_n25 ) , .B2( u0_r0_n6 ) );
  NAND4_X1 u0_r0_U38 (.ZN( u0_r0_n10 ) , .A1( u0_r0_n24 ) , .A2( u0_r0_n25 ) , .A4( u0_r0_n3 ) , .A3( u0_r0_n9 ) );
  OAI22_X1 u0_r0_U39 (.ZN( u0_r0_N73 ) , .B1( u0_r0_n16 ) , .A2( u0_r0_n19 ) , .B2( u0_r0_n20 ) , .A1( u0_r0_rcnt_0 ) );
  NAND2_X1 u0_r0_U40 (.A1( u0_r0_n12 ) , .ZN( u0_r0_n20 ) , .A2( u0_r0_rcnt_0 ) );
  NOR3_X1 u0_r0_U41 (.ZN( u0_r0_N76 ) , .A1( u0_r0_n11 ) , .A2( u0_r0_n12 ) , .A3( u0_r0_n8 ) );
  NOR3_X1 u0_r0_U42 (.ZN( u0_r0_N77 ) , .A1( u0_r0_n11 ) , .A3( u0_r0_n12 ) , .A2( u0_r0_rcnt_0 ) );
  NAND2_X1 u0_r0_U43 (.ZN( u0_r0_n21 ) , .A1( u0_r0_rcnt_0 ) , .A2( u0_r0_rcnt_1 ) );
  NOR2_X1 u0_r0_U44 (.A2( ld ) , .ZN( u0_r0_N78 ) , .A1( u0_r0_rcnt_0 ) );
  OAI21_X1 u0_r0_U45 (.ZN( u0_r0_N72 ) , .A( u0_r0_n14 ) , .B2( u0_r0_n19 ) , .B1( u0_r0_n8 ) );
  OAI21_X1 u0_r0_U46 (.ZN( u0_r0_N75 ) , .B1( u0_r0_n11 ) , .B2( u0_r0_n13 ) , .A( u0_r0_n14 ) );
  NAND2_X1 u0_r0_U47 (.A1( u0_r0_n12 ) , .ZN( u0_r0_n13 ) , .A2( u0_r0_n8 ) );
  NOR2_X1 u0_r0_U48 (.A2( u0_r0_n21 ) , .ZN( u0_r0_n22 ) , .A1( u0_r0_n6 ) );
  OAI21_X1 u0_r0_U49 (.B1( u0_r0_N70 ) , .ZN( u0_r0_N81 ) , .A( u0_r0_n10 ) , .B2( u0_r0_n3 ) );
  NAND2_X1 u0_r0_U50 (.ZN( u0_r0_N74 ) , .A2( u0_r0_n1 ) , .A1( u0_r0_n14 ) );
  INV_X1 u0_r0_U51 (.ZN( u0_r0_n1 ) , .A( u0_r0_n15 ) );
  AOI211_X1 u0_r0_U52 (.C2( u0_r0_n11 ) , .ZN( u0_r0_n15 ) , .C1( u0_r0_n16 ) , .B( u0_r0_n7 ) , .A( u0_r0_n8 ) );
  INV_X1 u0_r0_U53 (.A( u0_r0_n12 ) , .ZN( u0_r0_n7 ) );
  INV_X1 u0_r0_U54 (.A( ld ) , .ZN( u0_r0_n9 ) );
  NAND3_X1 u0_r0_U55 (.ZN( u0_r0_n16 ) , .A3( u0_r0_n18 ) , .A1( u0_r0_n2 ) , .A2( u0_r0_n9 ) );
  NAND3_X1 u0_r0_U56 (.A3( u0_r0_N79 ) , .A1( u0_r0_n17 ) , .A2( u0_r0_n18 ) , .ZN( u0_r0_n19 ) );
  XOR2_X1 u0_r0_U57 (.Z( u0_r0_n18 ) , .A( u0_r0_n21 ) , .B( u0_r0_rcnt_2 ) );
  XOR2_X1 u0_r0_U58 (.Z( u0_r0_n17 ) , .B( u0_r0_n22 ) , .A( u0_r0_n3 ) );
  NAND3_X1 u0_r0_U59 (.ZN( u0_r0_n23 ) , .A3( u0_r0_n4 ) , .A1( u0_r0_n5 ) , .A2( u0_r0_n9 ) );
  XOR2_X1 u0_r0_U60 (.B( u0_r0_n12 ) , .Z( u0_r0_n24 ) , .A( u0_r0_n6 ) );
  DFF_X1 u0_r0_out_reg_24 (.CK( clk ) , .D( u0_r0_N70 ) , .Q( u0_rcon_24 ) );
  DFF_X1 u0_r0_out_reg_25 (.CK( clk ) , .D( u0_r0_N71 ) , .Q( u0_rcon_25 ) );
  DFF_X1 u0_r0_out_reg_26 (.CK( clk ) , .D( u0_r0_N72 ) , .Q( u0_rcon_26 ) );
  DFF_X1 u0_r0_out_reg_27 (.CK( clk ) , .D( u0_r0_N73 ) , .Q( u0_rcon_27 ) );
  DFF_X1 u0_r0_out_reg_28 (.CK( clk ) , .D( u0_r0_N74 ) , .Q( u0_rcon_28 ) );
  DFF_X1 u0_r0_out_reg_29 (.CK( clk ) , .D( u0_r0_N75 ) , .Q( u0_rcon_29 ) );
  DFF_X1 u0_r0_out_reg_30 (.CK( clk ) , .D( u0_r0_N76 ) , .Q( u0_rcon_30 ) );
  DFF_X1 u0_r0_out_reg_31 (.CK( clk ) , .D( u0_r0_N77 ) , .Q( u0_rcon_31 ) );
  DFF_X1 u0_r0_rcnt_reg_0 (.CK( clk ) , .D( u0_r0_N78 ) , .QN( u0_r0_n8 ) , .Q( u0_r0_rcnt_0 ) );
  DFF_X1 u0_r0_rcnt_reg_1 (.CK( clk ) , .D( u0_r0_N79 ) , .Q( u0_r0_rcnt_1 ) );
  DFF_X1 u0_r0_rcnt_reg_2 (.CK( clk ) , .D( u0_r0_N80 ) , .QN( u0_r0_n6 ) , .Q( u0_r0_rcnt_2 ) );
  DFF_X1 u0_r0_rcnt_reg_3 (.CK( clk ) , .D( u0_r0_N81 ) , .QN( u0_r0_n3 ) );
  INV_X1 u0_u0_U10 (.A( u0_u0_n1 ) , .ZN( u0_u0_n440 ) );
  AOI22_X1 u0_u0_U100 (.A2( u0_u0_n787 ) , .ZN( u0_u0_n788 ) , .B2( u0_u0_n836 ) , .A1( u0_u0_n839 ) , .B1( u0_u0_n867 ) );
  INV_X1 u0_u0_U101 (.A( u0_u0_n767 ) , .ZN( u0_u0_n835 ) );
  NOR2_X1 u0_u0_U102 (.ZN( u0_u0_n653 ) , .A1( u0_u0_n859 ) , .A2( u0_u0_n872 ) );
  INV_X1 u0_u0_U103 (.A( u0_u0_n759 ) , .ZN( u0_u0_n873 ) );
  OAI21_X1 u0_u0_U104 (.A( u0_u0_n439 ) , .B1( u0_u0_n758 ) , .ZN( u0_u0_n759 ) , .B2( u0_u0_n872 ) );
  NOR4_X1 u0_u0_U105 (.A4( u0_u0_n671 ) , .A3( u0_u0_n672 ) , .A2( u0_u0_n673 ) , .A1( u0_u0_n674 ) , .ZN( u0_u0_n682 ) );
  NOR4_X1 u0_u0_U106 (.A4( u0_u0_n667 ) , .A3( u0_u0_n668 ) , .A2( u0_u0_n669 ) , .A1( u0_u0_n670 ) , .ZN( u0_u0_n683 ) );
  NOR2_X1 u0_u0_U107 (.ZN( u0_u0_n738 ) , .A2( u0_u0_n837 ) , .A1( u0_u0_n850 ) );
  OR4_X1 u0_u0_U108 (.ZN( u0_u0_n472 ) , .A4( u0_u0_n524 ) , .A3( u0_u0_n535 ) , .A2( u0_u0_n584 ) , .A1( u0_u0_n717 ) );
  OR4_X1 u0_u0_U109 (.A4( u0_u0_n524 ) , .A2( u0_u0_n525 ) , .A1( u0_u0_n526 ) , .ZN( u0_u0_n528 ) , .A3( u0_u0_n826 ) );
  NAND2_X2 u0_u0_U11 (.A1( u0_u0_n455 ) , .A2( u0_u0_n466 ) , .ZN( u0_u0_n797 ) );
  OR4_X1 u0_u0_U110 (.A4( u0_u0_n688 ) , .A3( u0_u0_n689 ) , .A2( u0_u0_n690 ) , .A1( u0_u0_n691 ) , .ZN( u0_u0_n696 ) );
  OR4_X1 u0_u0_U111 (.A4( u0_u0_n572 ) , .A3( u0_u0_n573 ) , .A2( u0_u0_n574 ) , .ZN( u0_u0_n578 ) , .A1( u0_u0_n671 ) );
  OR4_X1 u0_u0_U112 (.ZN( u0_u0_n498 ) , .A4( u0_u0_n540 ) , .A2( u0_u0_n553 ) , .A1( u0_u0_n565 ) , .A3( u0_u0_n638 ) );
  INV_X1 u0_u0_U113 (.A( u0_u0_n442 ) , .ZN( u0_u0_n843 ) );
  OR3_X1 u0_u0_U114 (.A3( u0_u0_n512 ) , .A2( u0_u0_n513 ) , .A1( u0_u0_n514 ) , .ZN( u0_u0_n517 ) );
  INV_X1 u0_u0_U115 (.A( u0_u0_n469 ) , .ZN( u0_u0_n868 ) );
  OAI21_X1 u0_u0_U116 (.ZN( u0_u0_n469 ) , .B1( u0_u0_n814 ) , .A( u0_u0_n839 ) , .B2( u0_u0_n856 ) );
  AOI221_X1 u0_u0_U117 (.A( u0_u0_n718 ) , .B2( u0_u0_n719 ) , .ZN( u0_u0_n725 ) , .C1( u0_u0_n837 ) , .B1( u0_u0_n844 ) , .C2( u0_u0_n867 ) );
  OR2_X1 u0_u0_U118 (.A2( u0_u0_n716 ) , .A1( u0_u0_n717 ) , .ZN( u0_u0_n718 ) );
  NOR4_X1 u0_u0_U119 (.A4( u0_u0_n504 ) , .A3( u0_u0_n505 ) , .A2( u0_u0_n506 ) , .ZN( u0_u0_n507 ) , .A1( u0_u0_n533 ) );
  NAND2_X1 u0_u0_U12 (.A1( u0_u0_n457 ) , .A2( u0_u0_n477 ) , .ZN( u0_u0_n821 ) );
  NOR4_X1 u0_u0_U120 (.A4( u0_u0_n823 ) , .A3( u0_u0_n824 ) , .A2( u0_u0_n825 ) , .A1( u0_u0_n826 ) , .ZN( u0_u0_n827 ) );
  INV_X1 u0_u0_U121 (.A( u0_u0_n754 ) , .ZN( u0_u0_n867 ) );
  AOI221_X1 u0_u0_U122 (.C1( u0_u0_n444 ) , .A( u0_u0_n769 ) , .ZN( u0_u0_n779 ) , .C2( u0_u0_n815 ) , .B2( u0_u0_n840 ) , .B1( u0_u0_n870 ) );
  INV_X1 u0_u0_U123 (.A( u0_u0_n766 ) , .ZN( u0_u0_n840 ) );
  INV_X1 u0_u0_U124 (.A( u0_u0_n735 ) , .ZN( u0_u0_n844 ) );
  INV_X1 u0_u0_U125 (.A( u0_u0_n795 ) , .ZN( u0_u0_n837 ) );
  AOI211_X1 u0_u0_U126 (.B( u0_u0_n595 ) , .A( u0_u0_n596 ) , .ZN( u0_u0_n602 ) , .C2( u0_u0_n816 ) , .C1( u0_u0_n838 ) );
  AOI211_X1 u0_u0_U127 (.A( u0_u0_n502 ) , .ZN( u0_u0_n509 ) , .B( u0_u0_n807 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n856 ) );
  OAI221_X1 u0_u0_U128 (.A( u0_u0_n732 ) , .C2( u0_u0_n733 ) , .B2( u0_u0_n734 ) , .B1( u0_u0_n735 ) , .ZN( u0_u0_n742 ) , .C1( u0_u0_n822 ) );
  AOI22_X1 u0_u0_U129 (.ZN( u0_u0_n732 ) , .B1( u0_u0_n837 ) , .A2( u0_u0_n843 ) , .A1( u0_u0_n867 ) , .B2( u0_u0_n870 ) );
  NAND2_X1 u0_u0_U13 (.A2( u0_u0_n459 ) , .A1( u0_u0_n461 ) , .ZN( u0_u0_n811 ) );
  NOR4_X1 u0_u0_U130 (.A4( u0_u0_n645 ) , .A3( u0_u0_n646 ) , .A2( u0_u0_n647 ) , .A1( u0_u0_n648 ) , .ZN( u0_u0_n649 ) );
  AOI21_X1 u0_u0_U131 (.ZN( u0_u0_n645 ) , .B2( u0_u0_n754 ) , .A( u0_u0_n793 ) , .B1( u0_u0_n817 ) );
  NOR4_X1 u0_u0_U132 (.A4( u0_u0_n798 ) , .A3( u0_u0_n799 ) , .A2( u0_u0_n800 ) , .A1( u0_u0_n801 ) , .ZN( u0_u0_n802 ) );
  OAI21_X1 u0_u0_U133 (.A( u0_u0_n792 ) , .B2( u0_u0_n793 ) , .B1( u0_u0_n794 ) , .ZN( u0_u0_n800 ) );
  OAI221_X1 u0_u0_U134 (.A( u0_u0_n788 ) , .C2( u0_u0_n789 ) , .B2( u0_u0_n790 ) , .B1( u0_u0_n791 ) , .ZN( u0_u0_n801 ) , .C1( u0_u0_n818 ) );
  NOR3_X1 u0_u0_U135 (.ZN( u0_u0_n496 ) , .A1( u0_u0_n787 ) , .A2( u0_u0_n855 ) , .A3( u0_u0_n867 ) );
  AOI211_X1 u0_u0_U136 (.B( u0_u0_n750 ) , .A( u0_u0_n751 ) , .ZN( u0_u0_n764 ) , .C1( u0_u0_n837 ) , .C2( u0_u0_n858 ) );
  AOI211_X1 u0_u0_U137 (.B( u0_u0_n700 ) , .A( u0_u0_n701 ) , .ZN( u0_u0_n711 ) , .C2( u0_u0_n836 ) , .C1( u0_u0_n856 ) );
  AOI211_X1 u0_u0_U138 (.C2( u0_u0_n444 ) , .B( u0_u0_n730 ) , .A( u0_u0_n731 ) , .ZN( u0_u0_n744 ) , .C1( u0_u0_n848 ) );
  INV_X1 u0_u0_U139 (.A( u0_u0_n793 ) , .ZN( u0_u0_n850 ) );
  NOR3_X1 u0_u0_U14 (.A3( u0_u0_n171 ) , .A1( u0_u0_n622 ) , .A2( u0_u0_n623 ) , .ZN( u0_u0_n624 ) );
  NOR2_X1 u0_u0_U140 (.ZN( u0_u0_n672 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U141 (.ZN( u0_u0_n576 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U142 (.ZN( u0_u0_n538 ) , .A2( u0_u0_n754 ) , .A1( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U143 (.ZN( u0_u0_n512 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n767 ) );
  BUF_X2 u0_u0_U144 (.Z( u0_u0_n441 ) , .A( u0_u0_n796 ) );
  CLKBUF_X3 u0_u0_U145 (.Z( u0_u0_n442 ) , .A( u0_u0_n703 ) );
  NOR2_X1 u0_u0_U146 (.ZN( u0_u0_n667 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n795 ) );
  NOR2_X1 u0_u0_U147 (.ZN( u0_u0_n515 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U148 (.ZN( u0_u0_n673 ) , .A1( u0_u0_n755 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U149 (.A( u0_u0_n819 ) , .ZN( u0_u0_n838 ) );
  NOR3_X1 u0_u0_U15 (.A3( u0_u0_n438 ) , .A1( u0_u0_n781 ) , .ZN( u0_u0_n804 ) , .A2( u0_u0_n806 ) );
  NOR2_X1 u0_u0_U150 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n668 ) , .A1( u0_u0_n734 ) );
  NOR2_X1 u0_u0_U151 (.ZN( u0_u0_n669 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U152 (.ZN( u0_u0_n513 ) , .A1( u0_u0_n817 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U153 (.ZN( u0_u0_n661 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U154 (.ZN( u0_u0_n551 ) , .A1( u0_u0_n754 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U155 (.ZN( u0_u0_n636 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U156 (.A1( u0_u0_n754 ) , .ZN( u0_u0_n772 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U157 (.A1( u0_u0_n442 ) , .ZN( u0_u0_n775 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U158 (.A( u0_u0_n752 ) , .ZN( u0_u0_n839 ) );
  INV_X1 u0_u0_U159 (.A( u0_u0_n755 ) , .ZN( u0_u0_n847 ) );
  OR4_X1 u0_u0_U16 (.A4( u0_u0_n586 ) , .A3( u0_u0_n587 ) , .A2( u0_u0_n588 ) , .A1( u0_u0_n589 ) , .ZN( u0_u0_n590 ) );
  NOR2_X1 u0_u0_U160 (.ZN( u0_u0_n621 ) , .A1( u0_u0_n790 ) , .A2( u0_u0_n820 ) );
  NOR2_X1 u0_u0_U161 (.ZN( u0_u0_n635 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U162 (.ZN( u0_u0_n716 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n768 ) );
  NOR2_X1 u0_u0_U163 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n600 ) , .A1( u0_u0_n733 ) );
  NOR2_X1 u0_u0_U164 (.ZN( u0_u0_n620 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U165 (.B1( u0_u0_n631 ) , .ZN( u0_u0_n633 ) , .A( u0_u0_n768 ) , .B2( u0_u0_n819 ) );
  AOI21_X1 u0_u0_U166 (.ZN( u0_u0_n597 ) , .B2( u0_u0_n768 ) , .A( u0_u0_n790 ) , .B1( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U167 (.ZN( u0_u0_n521 ) , .A( u0_u0_n734 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n808 ) );
  AOI21_X1 u0_u0_U168 (.ZN( u0_u0_n545 ) , .B2( u0_u0_n817 ) , .A( u0_u0_n819 ) , .B1( u0_u0_n820 ) );
  INV_X1 u0_u0_U169 (.A( u0_u0_n808 ) , .ZN( u0_u0_n848 ) );
  NOR2_X1 u0_u0_U17 (.A2( u0_u0_n22 ) , .A1( u0_u0_n590 ) , .ZN( u0_u0_n591 ) );
  AOI21_X1 u0_u0_U170 (.ZN( u0_u0_n546 ) , .A( u0_u0_n768 ) , .B2( u0_u0_n784 ) , .B1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U171 (.ZN( u0_u0_n574 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n767 ) );
  AOI21_X1 u0_u0_U172 (.B1( u0_u0_n692 ) , .ZN( u0_u0_n693 ) , .A( u0_u0_n733 ) , .B2( u0_u0_n766 ) );
  NOR2_X1 u0_u0_U173 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n572 ) , .A1( u0_u0_n768 ) );
  INV_X1 u0_u0_U174 (.A( u0_u0_n733 ) , .ZN( u0_u0_n857 ) );
  INV_X1 u0_u0_U175 (.A( u0_u0_n734 ) , .ZN( u0_u0_n872 ) );
  AOI21_X1 u0_u0_U176 (.B2( u0_u0_n442 ) , .ZN( u0_u0_n577 ) , .B1( u0_u0_n811 ) , .A( u0_u0_n817 ) );
  NOR2_X1 u0_u0_U177 (.ZN( u0_u0_n527 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U178 (.ZN( u0_u0_n695 ) , .B2( u0_u0_n754 ) , .B1( u0_u0_n768 ) , .A( u0_u0_n811 ) );
  AOI21_X1 u0_u0_U179 (.B2( u0_u0_n442 ) , .ZN( u0_u0_n484 ) , .A( u0_u0_n754 ) , .B1( u0_u0_n784 ) );
  NOR3_X1 u0_u0_U18 (.A3( u0_u0_n805 ) , .A2( u0_u0_n806 ) , .A1( u0_u0_n807 ) , .ZN( u0_u0_n830 ) );
  INV_X1 u0_u0_U180 (.A( u0_u0_n817 ) , .ZN( u0_u0_n859 ) );
  INV_X1 u0_u0_U181 (.A( u0_u0_n811 ) , .ZN( u0_u0_n846 ) );
  INV_X1 u0_u0_U182 (.A( u0_u0_n768 ) , .ZN( u0_u0_n870 ) );
  OAI21_X1 u0_u0_U183 (.A( u0_u0_n704 ) , .ZN( u0_u0_n708 ) , .B2( u0_u0_n755 ) , .B1( u0_u0_n809 ) );
  OAI21_X1 u0_u0_U184 (.ZN( u0_u0_n704 ) , .B2( u0_u0_n838 ) , .B1( u0_u0_n843 ) , .A( u0_u0_n864 ) );
  NOR2_X1 u0_u0_U185 (.ZN( u0_u0_n476 ) , .A2( u0_u0_n784 ) , .A1( u0_u0_n820 ) );
  NAND2_X1 u0_u0_U186 (.A2( u0_u0_n767 ) , .A1( u0_u0_n811 ) , .ZN( u0_u0_n815 ) );
  BUF_X1 u0_u0_U187 (.Z( u0_u0_n443 ) , .A( u0_u0_n818 ) );
  INV_X1 u0_u0_U188 (.A( u0_u0_n790 ) , .ZN( u0_u0_n851 ) );
  INV_X1 u0_u0_U189 (.A( u0_u0_n822 ) , .ZN( u0_u0_n849 ) );
  NOR3_X1 u0_u0_U19 (.ZN( u0_u0_n604 ) , .A1( u0_u0_n614 ) , .A3( u0_u0_n728 ) , .A2( u0_u0_n747 ) );
  OAI22_X1 u0_u0_U190 (.B2( u0_u0_n755 ) , .B1( u0_u0_n756 ) , .A1( u0_u0_n757 ) , .ZN( u0_u0_n761 ) , .A2( u0_u0_n811 ) );
  NOR3_X1 u0_u0_U191 (.ZN( u0_u0_n757 ) , .A2( u0_u0_n858 ) , .A1( u0_u0_n867 ) , .A3( u0_u0_n869 ) );
  NOR2_X1 u0_u0_U192 (.ZN( u0_u0_n756 ) , .A2( u0_u0_n857 ) , .A1( u0_u0_n864 ) );
  AND2_X1 u0_u0_U193 (.ZN( u0_u0_n753 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n791 ) );
  AND2_X1 u0_u0_U194 (.ZN( u0_u0_n737 ) , .A1( u0_u0_n784 ) , .A2( u0_u0_n790 ) );
  AOI221_X1 u0_u0_U195 (.A( u0_u0_n503 ) , .ZN( u0_u0_n508 ) , .B2( u0_u0_n848 ) , .C1( u0_u0_n851 ) , .C2( u0_u0_n864 ) , .B1( u0_u0_n866 ) );
  AOI221_X1 u0_u0_U196 (.A( u0_u0_n687 ) , .ZN( u0_u0_n698 ) , .B2( u0_u0_n845 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n866 ) , .B1( u0_u0_n869 ) );
  INV_X1 u0_u0_U197 (.A( u0_u0_n686 ) , .ZN( u0_u0_n845 ) );
  OAI221_X1 u0_u0_U198 (.A( u0_u0_n702 ) , .ZN( u0_u0_n709 ) , .C2( u0_u0_n789 ) , .C1( u0_u0_n790 ) , .B1( u0_u0_n791 ) , .B2( u0_u0_n811 ) );
  AOI22_X1 u0_u0_U199 (.ZN( u0_u0_n702 ) , .A1( u0_u0_n835 ) , .B2( u0_u0_n848 ) , .A2( u0_u0_n869 ) , .B1( u0_u0_n872 ) );
  NOR3_X1 u0_u0_U20 (.A1( u0_u0_n1 ) , .ZN( u0_u0_n510 ) , .A2( u0_u0_n685 ) , .A3( u0_u0_n782 ) );
  OAI222_X1 u0_u0_U200 (.A2( u0_u0_n675 ) , .ZN( u0_u0_n680 ) , .B1( u0_u0_n752 ) , .B2( u0_u0_n789 ) , .C2( u0_u0_n793 ) , .C1( u0_u0_n820 ) , .A1( u0_u0_n822 ) );
  NAND2_X1 u0_u0_U201 (.A2( u0_u0_n454 ) , .A1( u0_u0_n466 ) , .ZN( u0_u0_n733 ) );
  NAND2_X1 u0_u0_U202 (.A2( u0_u0_n454 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n734 ) );
  NAND2_X1 u0_u0_U203 (.A2( u0_u0_n455 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n768 ) );
  NAND2_X1 u0_u0_U204 (.A2( u0_u0_n454 ) , .A1( u0_u0_n470 ) , .ZN( u0_u0_n820 ) );
  NAND2_X1 u0_u0_U205 (.A2( u0_u0_n466 ) , .A1( u0_u0_n471 ) , .ZN( u0_u0_n785 ) );
  NAND2_X1 u0_u0_U206 (.A1( u0_u0_n453 ) , .A2( u0_u0_n471 ) , .ZN( u0_u0_n754 ) );
  NOR2_X1 u0_u0_U207 (.ZN( u0_u0_n471 ) , .A2( u0_u0_n852 ) , .A1( u0_u0_n853 ) );
  NAND2_X1 u0_u0_U208 (.A2( u0_u0_n467 ) , .A1( u0_u0_n468 ) , .ZN( u0_u0_n752 ) );
  NAND2_X1 u0_u0_U209 (.A1( u0_u0_n468 ) , .A2( u0_u0_n478 ) , .ZN( u0_u0_n793 ) );
  NOR3_X1 u0_u0_U21 (.A2( u0_u0_n613 ) , .A1( u0_u0_n614 ) , .ZN( u0_u0_n652 ) , .A3( u0_u0_n727 ) );
  NOR4_X1 u0_u0_U210 (.A4( u0_u0_n739 ) , .A3( u0_u0_n740 ) , .A2( u0_u0_n741 ) , .A1( u0_u0_n742 ) , .ZN( u0_u0_n743 ) );
  NOR4_X1 u0_u0_U211 (.A4( u0_u0_n706 ) , .A3( u0_u0_n707 ) , .A2( u0_u0_n708 ) , .A1( u0_u0_n709 ) , .ZN( u0_u0_n710 ) );
  NOR4_X1 u0_u0_U212 (.A3( u0_u0_n760 ) , .A2( u0_u0_n761 ) , .A1( u0_u0_n762 ) , .ZN( u0_u0_n763 ) , .A4( u0_u0_n873 ) );
  NOR2_X1 u0_u0_U213 (.ZN( u0_u0_n477 ) , .A1( u0_u0_n831 ) , .A2( w3_17 ) );
  AOI221_X1 u0_u0_U214 (.A( u0_u0_n786 ) , .ZN( u0_u0_n803 ) , .C2( u0_u0_n842 ) , .B2( u0_u0_n843 ) , .B1( u0_u0_n869 ) , .C1( u0_u0_n870 ) );
  NAND4_X1 u0_u0_U215 (.ZN( u0_subword_25 ) , .A4( u0_u0_n601 ) , .A3( u0_u0_n602 ) , .A2( u0_u0_n603 ) , .A1( u0_u0_n604 ) );
  NOR4_X1 u0_u0_U216 (.A4( u0_u0_n597 ) , .A3( u0_u0_n598 ) , .A2( u0_u0_n599 ) , .A1( u0_u0_n600 ) , .ZN( u0_u0_n601 ) );
  NAND4_X1 u0_u0_U217 (.ZN( u0_subword_24 ) , .A4( u0_u0_n507 ) , .A3( u0_u0_n508 ) , .A2( u0_u0_n509 ) , .A1( u0_u0_n510 ) );
  AOI222_X1 u0_u0_U218 (.B2( u0_u0_n644 ) , .ZN( u0_u0_n650 ) , .B1( u0_u0_n846 ) , .A1( u0_u0_n847 ) , .C2( u0_u0_n851 ) , .C1( u0_u0_n867 ) , .A2( u0_u0_n869 ) );
  AND2_X1 u0_u0_U219 (.ZN( u0_u0_n453 ) , .A2( w3_22 ) , .A1( w3_23 ) );
  NOR3_X1 u0_u0_U22 (.A3( u0_u0_n746 ) , .A2( u0_u0_n747 ) , .A1( u0_u0_n748 ) , .ZN( u0_u0_n765 ) );
  NAND4_X1 u0_u0_U220 (.ZN( u0_subword_31 ) , .A4( u0_u0_n827 ) , .A3( u0_u0_n828 ) , .A2( u0_u0_n829 ) , .A1( u0_u0_n830 ) );
  AOI222_X1 u0_u0_U221 (.C2( u0_u0_n814 ) , .B2( u0_u0_n815 ) , .A2( u0_u0_n816 ) , .ZN( u0_u0_n828 ) , .C1( u0_u0_n837 ) , .A1( u0_u0_n844 ) , .B1( u0_u0_n858 ) );
  INV_X1 u0_u0_U222 (.ZN( u0_u0_n853 ) , .A( w3_21 ) );
  NAND4_X1 u0_u0_U223 (.A4( u0_u0_n697 ) , .A3( u0_u0_n698 ) , .A1( u0_u0_n699 ) , .ZN( u0_u0_n781 ) , .A2( u0_u0_n876 ) );
  NAND2_X2 u0_u0_U224 (.A2( u0_u0_n470 ) , .A1( u0_u0_n471 ) , .ZN( u0_u0_n817 ) );
  NAND2_X1 u0_u0_U225 (.A2( u0_u0_n447 ) , .A1( u0_u0_n458 ) , .ZN( u0_u0_n796 ) );
  AOI222_X1 u0_u0_U226 (.ZN( u0_u0_n780 ) , .A1( u0_u0_n835 ) , .C1( u0_u0_n839 ) , .B2( u0_u0_n846 ) , .A2( u0_u0_n855 ) , .B1( u0_u0_n865 ) , .C2( u0_u0_n877 ) );
  OAI21_X1 u0_u0_U227 (.ZN( u0_u0_n736 ) , .A( u0_u0_n838 ) , .B2( u0_u0_n857 ) , .B1( u0_u0_n877 ) );
  AOI222_X1 u0_u0_U228 (.ZN( u0_u0_n569 ) , .B1( u0_u0_n835 ) , .C1( u0_u0_n846 ) , .A2( u0_u0_n848 ) , .A1( u0_u0_n859 ) , .B2( u0_u0_n867 ) , .C2( u0_u0_n877 ) );
  OAI21_X1 u0_u0_U229 (.ZN( u0_u0_n792 ) , .A( u0_u0_n844 ) , .B1( u0_u0_n867 ) , .B2( u0_u0_n877 ) );
  NOR3_X1 u0_u0_U23 (.A3( u0_u0_n727 ) , .A1( u0_u0_n728 ) , .ZN( u0_u0_n745 ) , .A2( u0_u0_n746 ) );
  NAND4_X1 u0_u0_U230 (.A4( u0_u0_n479 ) , .A3( u0_u0_n480 ) , .A2( u0_u0_n481 ) , .A1( u0_u0_n482 ) , .ZN( u0_u0_n684 ) );
  NOR4_X1 u0_u0_U231 (.ZN( u0_u0_n479 ) , .A2( u0_u0_n527 ) , .A4( u0_u0_n600 ) , .A1( u0_u0_n615 ) , .A3( u0_u0_n635 ) );
  NAND2_X1 u0_u0_U232 (.A2( u0_u0_n467 ) , .A1( u0_u0_n477 ) , .ZN( u0_u0_n703 ) );
  NAND2_X1 u0_u0_U233 (.A2( u0_u0_n460 ) , .A1( u0_u0_n461 ) , .ZN( u0_u0_n735 ) );
  NAND2_X1 u0_u0_U234 (.A1( u0_u0_n460 ) , .A2( u0_u0_n467 ) , .ZN( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U235 (.ZN( u0_u0_n461 ) , .A1( u0_u0_n833 ) , .A2( w3_19 ) );
  NAND2_X2 u0_u0_U236 (.A1( u0_u0_n457 ) , .A2( u0_u0_n460 ) , .ZN( u0_u0_n819 ) );
  AOI211_X1 u0_u0_U237 (.B( u0_u0_n812 ) , .A( u0_u0_n813 ) , .ZN( u0_u0_n829 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n855 ) );
  NOR2_X1 u0_u0_U238 (.A1( u0_u0_n684 ) , .ZN( u0_u0_n699 ) , .A2( u0_u0_n812 ) );
  OAI222_X1 u0_u0_U239 (.B1( u0_u0_n442 ) , .ZN( u0_u0_n623 ) , .C1( u0_u0_n729 ) , .C2( u0_u0_n752 ) , .B2( u0_u0_n791 ) , .A2( u0_u0_n797 ) , .A1( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U24 (.ZN( u0_u0_n581 ) , .A1( u0_u0_n628 ) , .A2( u0_u0_n750 ) );
  AOI21_X1 u0_u0_U240 (.A( u0_u0_n676 ) , .B1( u0_u0_n677 ) , .ZN( u0_u0_n678 ) , .B2( u0_u0_n860 ) );
  AOI21_X1 u0_u0_U241 (.B1( u0_u0_n445 ) , .ZN( u0_u0_n516 ) , .B2( u0_u0_n675 ) , .A( u0_u0_n735 ) );
  INV_X1 u0_u0_U242 (.A( u0_u0_n675 ) , .ZN( u0_u0_n869 ) );
  NOR2_X1 u0_u0_U243 (.ZN( u0_u0_n658 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U244 (.ZN( u0_u0_n533 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n784 ) );
  AOI21_X1 u0_u0_U245 (.ZN( u0_u0_n483 ) , .A( u0_u0_n675 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U246 (.ZN( u0_u0_n608 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U247 (.ZN( u0_u0_n634 ) , .A2( u0_u0_n675 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U248 (.ZN( u0_u0_n587 ) , .A1( u0_u0_n675 ) , .A2( u0_u0_n793 ) );
  NAND2_X2 u0_u0_U249 (.A1( u0_u0_n458 ) , .A2( u0_u0_n471 ) , .ZN( u0_u0_n675 ) );
  NOR2_X1 u0_u0_U25 (.ZN( u0_u0_n501 ) , .A1( u0_u0_n684 ) , .A2( u0_u0_n700 ) );
  NAND4_X1 u0_u0_U250 (.A4( u0_u0_n541 ) , .A3( u0_u0_n542 ) , .A2( u0_u0_n543 ) , .A1( u0_u0_n544 ) , .ZN( u0_u0_n628 ) );
  OAI222_X1 u0_u0_U251 (.A2( u0_u0_n445 ) , .B2( u0_u0_n713 ) , .ZN( u0_u0_n714 ) , .C2( u0_u0_n729 ) , .B1( u0_u0_n752 ) , .A1( u0_u0_n811 ) , .C1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U252 (.ZN( u0_u0_n524 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n793 ) );
  NOR2_X1 u0_u0_U253 (.ZN( u0_u0_n526 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U254 (.A2( u0_u0_n713 ) , .A1( u0_u0_n767 ) , .ZN( u0_u0_n799 ) );
  NOR2_X1 u0_u0_U255 (.A2( u0_u0_n713 ) , .A1( u0_u0_n755 ) , .ZN( u0_u0_n776 ) );
  NOR2_X1 u0_u0_U256 (.ZN( u0_u0_n523 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U257 (.ZN( u0_u0_n688 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n822 ) );
  OAI22_X1 u0_u0_U258 (.ZN( u0_u0_n489 ) , .A1( u0_u0_n713 ) , .B2( u0_u0_n790 ) , .A2( u0_u0_n811 ) , .B1( u0_u0_n817 ) );
  NOR2_X1 u0_u0_U259 (.ZN( u0_u0_n549 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U26 (.ZN( u0_u0_n712 ) , .A2( u0_u0_n781 ) , .A1( u0_u0_n805 ) );
  NOR2_X1 u0_u0_U260 (.ZN( u0_u0_n585 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n735 ) );
  NOR2_X1 u0_u0_U261 (.ZN( u0_u0_n535 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U262 (.ZN( u0_u0_n674 ) , .A2( u0_u0_n713 ) , .A1( u0_u0_n795 ) );
  AOI222_X1 u0_u0_U263 (.ZN( u0_u0_n531 ) , .A1( u0_u0_n839 ) , .B2( u0_u0_n842 ) , .C1( u0_u0_n849 ) , .C2( u0_u0_n855 ) , .A2( u0_u0_n857 ) , .B1( u0_u0_n870 ) );
  AOI222_X1 u0_u0_U264 (.ZN( u0_u0_n612 ) , .A1( u0_u0_n835 ) , .C2( u0_u0_n842 ) , .B1( u0_u0_n847 ) , .A2( u0_u0_n860 ) , .B2( u0_u0_n865 ) , .C1( u0_u0_n872 ) );
  NOR3_X1 u0_u0_U265 (.ZN( u0_u0_n446 ) , .A2( u0_u0_n841 ) , .A3( u0_u0_n842 ) , .A1( u0_u0_n851 ) );
  NAND2_X1 u0_u0_U266 (.ZN( u0_u0_n619 ) , .A2( u0_u0_n842 ) , .A1( u0_u0_n877 ) );
  OAI22_X1 u0_u0_U267 (.A1( u0_u0_n445 ) , .B2( u0_u0_n784 ) , .B1( u0_u0_n785 ) , .ZN( u0_u0_n786 ) , .A2( u0_u0_n819 ) );
  NAND4_X1 u0_u0_U268 (.A4( u0_u0_n499 ) , .A3( u0_u0_n500 ) , .A1( u0_u0_n501 ) , .ZN( u0_u0_n807 ) , .A2( u0_u0_n871 ) );
  AOI21_X1 u0_u0_U269 (.ZN( u0_u0_n575 ) , .B1( u0_u0_n755 ) , .B2( u0_u0_n767 ) , .A( u0_u0_n785 ) );
  AOI222_X1 u0_u0_U27 (.ZN( u0_u0_n666 ) , .A2( u0_u0_n844 ) , .B1( u0_u0_n846 ) , .C2( u0_u0_n850 ) , .A1( u0_u0_n864 ) , .C1( u0_u0_n867 ) , .B2( u0_u0_n874 ) );
  NAND2_X1 u0_u0_U270 (.ZN( u0_u0_n719 ) , .A1( u0_u0_n733 ) , .A2( u0_u0_n785 ) );
  OAI22_X1 u0_u0_U271 (.B1( u0_u0_n496 ) , .ZN( u0_u0_n497 ) , .A1( u0_u0_n692 ) , .A2( u0_u0_n768 ) , .B2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U272 (.ZN( u0_u0_n662 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n785 ) );
  NOR2_X1 u0_u0_U273 (.A2( u0_u0_n442 ) , .A1( u0_u0_n785 ) , .ZN( u0_u0_n825 ) );
  NOR2_X1 u0_u0_U274 (.ZN( u0_u0_n514 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U275 (.ZN( u0_u0_n607 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U276 (.ZN( u0_u0_n617 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U277 (.ZN( u0_u0_n552 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n819 ) );
  INV_X1 u0_u0_U278 (.A( u0_u0_n785 ) , .ZN( u0_u0_n855 ) );
  AOI21_X1 u0_u0_U279 (.ZN( u0_u0_n646 ) , .B2( u0_u0_n752 ) , .A( u0_u0_n797 ) , .B1( u0_u0_n808 ) );
  INV_X1 u0_u0_U28 (.A( u0_u0_n653 ) , .ZN( u0_u0_n874 ) );
  AOI21_X1 u0_u0_U280 (.A( u0_u0_n738 ) , .ZN( u0_u0_n739 ) , .B2( u0_u0_n785 ) , .B1( u0_u0_n797 ) );
  NAND4_X1 u0_u0_U281 (.A4( u0_u0_n554 ) , .A3( u0_u0_n555 ) , .A2( u0_u0_n556 ) , .A1( u0_u0_n557 ) , .ZN( u0_u0_n750 ) );
  AOI21_X1 u0_u0_U282 (.ZN( u0_u0_n520 ) , .A( u0_u0_n784 ) , .B2( u0_u0_n797 ) , .B1( u0_u0_n817 ) );
  AOI21_X1 u0_u0_U283 (.B2( u0_u0_n768 ) , .ZN( u0_u0_n769 ) , .A( u0_u0_n793 ) , .B1( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U284 (.ZN( u0_u0_n456 ) , .B2( u0_u0_n797 ) , .A( u0_u0_n808 ) , .B1( u0_u0_n820 ) );
  INV_X1 u0_u0_U285 (.A( u0_u0_n797 ) , .ZN( u0_u0_n856 ) );
  NOR2_X1 u0_u0_U286 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n721 ) , .A1( u0_u0_n797 ) );
  NOR2_X1 u0_u0_U287 (.ZN( u0_u0_n563 ) , .A1( u0_u0_n797 ) , .A2( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U288 (.ZN( u0_u0_n589 ) , .A1( u0_u0_n797 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U289 (.ZN( u0_u0_n550 ) , .A2( u0_u0_n790 ) , .A1( u0_u0_n797 ) );
  NOR4_X1 u0_u0_U29 (.ZN( u0_u0_n491 ) , .A2( u0_u0_n539 ) , .A1( u0_u0_n564 ) , .A3( u0_u0_n637 ) , .A4( u0_u0_n723 ) );
  INV_X1 u0_u0_U290 (.ZN( u0_u0_n444 ) , .A( u0_u0_n820 ) );
  INV_X1 u0_u0_U291 (.A( u0_u0_n444 ) , .ZN( u0_u0_n445 ) );
  NOR4_X1 u0_u0_U292 (.A2( u0_u0_n497 ) , .A1( u0_u0_n498 ) , .ZN( u0_u0_n499 ) , .A3( u0_u0_n586 ) , .A4( u0_u0_n618 ) );
  INV_X1 u0_u0_U293 (.ZN( u0_u0_n832 ) , .A( w3_17 ) );
  AOI21_X1 u0_u0_U294 (.B1( u0_u0_n445 ) , .ZN( u0_u0_n595 ) , .B2( u0_u0_n705 ) , .A( u0_u0_n822 ) );
  AOI21_X1 u0_u0_U295 (.B1( u0_u0_n705 ) , .ZN( u0_u0_n706 ) , .A( u0_u0_n737 ) , .B2( u0_u0_n768 ) );
  INV_X1 u0_u0_U296 (.A( u0_u0_n705 ) , .ZN( u0_u0_n858 ) );
  AOI21_X1 u0_u0_U297 (.ZN( u0_u0_n448 ) , .A( u0_u0_n705 ) , .B1( u0_u0_n738 ) , .B2( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U298 (.ZN( u0_u0_n583 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U299 (.ZN( u0_u0_n689 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n808 ) );
  OR4_X1 u0_u0_U3 (.ZN( u0_u0_n1 ) , .A4( u0_u0_n451 ) , .A3( u0_u0_n452 ) , .A2( u0_u0_n522 ) , .A1( u0_u0_n547 ) );
  NOR4_X1 u0_u0_U30 (.ZN( u0_u0_n485 ) , .A1( u0_u0_n526 ) , .A4( u0_u0_n563 ) , .A3( u0_u0_n588 ) , .A2( u0_u0_n636 ) );
  NOR2_X1 u0_u0_U300 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n547 ) , .A1( u0_u0_n705 ) );
  NAND2_X1 u0_u0_U301 (.A1( u0_u0_n705 ) , .A2( u0_u0_n734 ) , .ZN( u0_u0_n787 ) );
  NAND2_X2 u0_u0_U302 (.A1( u0_u0_n447 ) , .A2( u0_u0_n466 ) , .ZN( u0_u0_n705 ) );
  NOR4_X1 u0_u0_U303 (.A3( u0_u0_n679 ) , .A1( u0_u0_n680 ) , .ZN( u0_u0_n681 ) , .A4( u0_u0_n720 ) , .A2( u0_u0_n863 ) );
  INV_X1 u0_u0_U304 (.A( u0_u0_n678 ) , .ZN( u0_u0_n863 ) );
  NOR2_X1 u0_u0_U305 (.ZN( u0_u0_n459 ) , .A1( u0_u0_n831 ) , .A2( u0_u0_n832 ) );
  AOI21_X1 u0_u0_U306 (.ZN( u0_u0_n504 ) , .A( u0_u0_n729 ) , .B2( u0_u0_n767 ) , .B1( u0_u0_n819 ) );
  OAI22_X1 u0_u0_U307 (.ZN( u0_u0_n495 ) , .A1( u0_u0_n729 ) , .B2( u0_u0_n733 ) , .B1( u0_u0_n735 ) , .A2( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U308 (.ZN( u0_u0_n717 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n795 ) );
  NOR2_X1 u0_u0_U309 (.ZN( u0_u0_n534 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n808 ) );
  NOR4_X1 u0_u0_U31 (.ZN( u0_u0_n462 ) , .A2( u0_u0_n523 ) , .A1( u0_u0_n549 ) , .A3( u0_u0_n585 ) , .A4( u0_u0_n621 ) );
  NOR2_X1 u0_u0_U310 (.ZN( u0_u0_n532 ) , .A1( u0_u0_n729 ) , .A2( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U311 (.ZN( u0_u0_n615 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U312 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n638 ) , .A1( u0_u0_n729 ) );
  NOR2_X1 u0_u0_U313 (.ZN( u0_u0_n540 ) , .A1( u0_u0_n729 ) , .A2( u0_u0_n793 ) );
  NOR2_X1 u0_u0_U314 (.ZN( u0_u0_n539 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n735 ) );
  INV_X1 u0_u0_U315 (.A( u0_u0_n729 ) , .ZN( u0_u0_n860 ) );
  NAND2_X2 u0_u0_U316 (.A1( u0_u0_n447 ) , .A2( u0_u0_n470 ) , .ZN( u0_u0_n713 ) );
  NAND2_X2 u0_u0_U317 (.A1( u0_u0_n455 ) , .A2( u0_u0_n470 ) , .ZN( u0_u0_n729 ) );
  AOI211_X1 u0_u0_U318 (.C1( u0_u0_n439 ) , .C2( u0_u0_n444 ) , .A( u0_u0_n594 ) , .ZN( u0_u0_n603 ) , .B( u0_u0_n627 ) );
  NOR3_X1 u0_u0_U319 (.A2( u0_u0_n627 ) , .A3( u0_u0_n628 ) , .ZN( u0_u0_n642 ) , .A1( u0_u0_n730 ) );
  OR3_X1 u0_u0_U32 (.ZN( u0_u0_n452 ) , .A1( u0_u0_n534 ) , .A3( u0_u0_n583 ) , .A2( u0_u0_n879 ) );
  AOI21_X1 u0_u0_U320 (.B2( u0_u0_n443 ) , .ZN( u0_u0_n599 ) , .B1( u0_u0_n755 ) , .A( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U321 (.A( u0_u0_n817 ) , .B2( u0_u0_n818 ) , .B1( u0_u0_n819 ) , .ZN( u0_u0_n824 ) );
  AOI21_X1 u0_u0_U322 (.A( u0_u0_n443 ) , .ZN( u0_u0_n655 ) , .B1( u0_u0_n734 ) , .B2( u0_u0_n768 ) );
  NOR2_X1 u0_u0_U323 (.A2( u0_u0_n818 ) , .A1( u0_u0_n820 ) , .ZN( u0_u0_n826 ) );
  NOR2_X1 u0_u0_U324 (.A2( u0_u0_n443 ) , .A1( u0_u0_n675 ) , .ZN( u0_u0_n771 ) );
  NOR2_X1 u0_u0_U325 (.ZN( u0_u0_n584 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U326 (.ZN( u0_u0_n671 ) , .A1( u0_u0_n785 ) , .A2( u0_u0_n818 ) );
  NAND2_X2 u0_u0_U327 (.A2( u0_u0_n460 ) , .A1( u0_u0_n478 ) , .ZN( u0_u0_n784 ) );
  NOR2_X1 u0_u0_U328 (.A1( u0_u0_n705 ) , .ZN( u0_u0_n773 ) , .A2( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U329 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n660 ) , .A1( u0_u0_n733 ) );
  INV_X1 u0_u0_U33 (.A( u0_u0_n619 ) , .ZN( u0_u0_n879 ) );
  NOR2_X1 u0_u0_U330 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n637 ) , .A1( u0_u0_n729 ) );
  INV_X1 u0_u0_U331 (.A( u0_u0_n818 ) , .ZN( u0_u0_n841 ) );
  NAND2_X2 u0_u0_U332 (.A1( u0_u0_n457 ) , .A2( u0_u0_n459 ) , .ZN( u0_u0_n767 ) );
  NOR2_X1 u0_u0_U333 (.ZN( u0_u0_n478 ) , .A1( w3_18 ) , .A2( w3_19 ) );
  AOI21_X1 u0_u0_U334 (.A( u0_u0_n441 ) , .ZN( u0_u0_n647 ) , .B1( u0_u0_n686 ) , .B2( u0_u0_n822 ) );
  NAND2_X2 u0_u0_U335 (.A1( u0_u0_n453 ) , .A2( u0_u0_n455 ) , .ZN( u0_u0_n810 ) );
  AOI21_X1 u0_u0_U336 (.B2( u0_u0_n441 ) , .A( u0_u0_n795 ) , .B1( u0_u0_n797 ) , .ZN( u0_u0_n798 ) );
  OAI22_X1 u0_u0_U337 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n701 ) , .A2( u0_u0_n735 ) , .A1( u0_u0_n785 ) , .B2( u0_u0_n822 ) );
  AOI21_X1 u0_u0_U338 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n503 ) , .A( u0_u0_n784 ) , .B1( u0_u0_n809 ) );
  AOI21_X1 u0_u0_U339 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n632 ) , .B2( u0_u0_n675 ) , .A( u0_u0_n795 ) );
  NOR4_X1 u0_u0_U34 (.A1( u0_u0_n537 ) , .ZN( u0_u0_n542 ) , .A2( u0_u0_n660 ) , .A4( u0_u0_n674 ) , .A3( u0_u0_n770 ) );
  NAND2_X2 u0_u0_U340 (.A1( u0_u0_n461 ) , .A2( u0_u0_n468 ) , .ZN( u0_u0_n755 ) );
  AOI21_X1 u0_u0_U341 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n570 ) , .B1( u0_u0_n729 ) , .A( u0_u0_n784 ) );
  NAND2_X2 u0_u0_U342 (.A1( u0_u0_n457 ) , .A2( u0_u0_n468 ) , .ZN( u0_u0_n795 ) );
  AOI21_X1 u0_u0_U343 (.B2( u0_u0_n441 ) , .ZN( u0_u0_n449 ) , .B1( u0_u0_n794 ) , .A( u0_u0_n819 ) );
  NOR2_X1 u0_u0_U344 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n670 ) , .A1( u0_u0_n790 ) );
  NOR2_X1 u0_u0_U345 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n561 ) , .A1( u0_u0_n755 ) );
  NOR2_X1 u0_u0_U346 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n565 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U347 (.A1( u0_u0_n441 ) , .A2( u0_u0_n443 ) , .ZN( u0_u0_n690 ) );
  NOR2_X1 u0_u0_U348 (.A1( u0_u0_n441 ) , .ZN( u0_u0_n648 ) , .A2( u0_u0_n793 ) );
  NAND2_X2 u0_u0_U349 (.A1( u0_u0_n453 ) , .A2( u0_u0_n454 ) , .ZN( u0_u0_n791 ) );
  NOR4_X1 u0_u0_U35 (.A4( u0_u0_n547 ) , .A3( u0_u0_n548 ) , .A2( u0_u0_n549 ) , .ZN( u0_u0_n556 ) , .A1( u0_u0_n694 ) );
  NOR2_X1 u0_u0_U350 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n548 ) , .A1( u0_u0_n767 ) );
  INV_X1 u0_u0_U351 (.A( u0_u0_n796 ) , .ZN( u0_u0_n877 ) );
  NOR2_X1 u0_u0_U352 (.ZN( u0_u0_n586 ) , .A2( u0_u0_n703 ) , .A1( u0_u0_n796 ) );
  NOR2_X1 u0_u0_U353 (.ZN( u0_u0_n467 ) , .A1( u0_u0_n834 ) , .A2( w3_18 ) );
  AOI221_X1 u0_u0_U354 (.A( u0_u0_n582 ) , .ZN( u0_u0_n593 ) , .B2( u0_u0_n836 ) , .C2( u0_u0_n848 ) , .B1( u0_u0_n859 ) , .C1( u0_u0_n865 ) );
  NOR2_X1 u0_u0_U355 (.ZN( u0_u0_n457 ) , .A1( u0_u0_n833 ) , .A2( u0_u0_n834 ) );
  INV_X1 u0_u0_U356 (.ZN( u0_u0_n834 ) , .A( w3_19 ) );
  NAND2_X2 u0_u0_U357 (.A1( u0_u0_n459 ) , .A2( u0_u0_n478 ) , .ZN( u0_u0_n790 ) );
  INV_X1 u0_u0_U358 (.ZN( u0_u0_n833 ) , .A( w3_18 ) );
  AOI222_X1 u0_u0_U359 (.ZN( u0_u0_n611 ) , .B2( u0_u0_n677 ) , .B1( u0_u0_n758 ) , .C2( u0_u0_n836 ) , .A1( u0_u0_n838 ) , .A2( u0_u0_n866 ) , .C1( u0_u0_n867 ) );
  NOR4_X1 u0_u0_U36 (.A4( u0_u0_n583 ) , .A3( u0_u0_n584 ) , .A2( u0_u0_n585 ) , .ZN( u0_u0_n592 ) , .A1( u0_u0_n689 ) );
  AOI222_X1 u0_u0_U360 (.ZN( u0_u0_n519 ) , .C1( u0_u0_n837 ) , .B2( u0_u0_n842 ) , .A2( u0_u0_n848 ) , .C2( u0_u0_n866 ) , .B1( u0_u0_n867 ) , .A1( u0_u0_n870 ) );
  AOI221_X1 u0_u0_U361 (.A( u0_u0_n489 ) , .ZN( u0_u0_n494 ) , .B1( u0_u0_n836 ) , .C2( u0_u0_n849 ) , .C1( u0_u0_n857 ) , .B2( u0_u0_n866 ) );
  NOR2_X1 u0_u0_U362 (.ZN( u0_u0_n794 ) , .A2( u0_u0_n866 ) , .A1( u0_u0_n872 ) );
  INV_X1 u0_u0_U363 (.A( u0_u0_n791 ) , .ZN( u0_u0_n866 ) );
  OAI22_X1 u0_u0_U364 (.ZN( u0_u0_n643 ) , .A1( u0_u0_n705 ) , .B2( u0_u0_n733 ) , .A2( u0_u0_n767 ) , .B1( u0_u0_n821 ) );
  OAI22_X1 u0_u0_U365 (.A1( u0_u0_n729 ) , .ZN( u0_u0_n731 ) , .B2( u0_u0_n755 ) , .B1( u0_u0_n817 ) , .A2( u0_u0_n821 ) );
  AOI21_X1 u0_u0_U366 (.ZN( u0_u0_n505 ) , .B1( u0_u0_n686 ) , .A( u0_u0_n817 ) , .B2( u0_u0_n821 ) );
  AOI21_X1 u0_u0_U367 (.A( u0_u0_n445 ) , .B2( u0_u0_n821 ) , .B1( u0_u0_n822 ) , .ZN( u0_u0_n823 ) );
  OAI22_X1 u0_u0_U368 (.A1( u0_u0_n445 ) , .ZN( u0_u0_n630 ) , .B1( u0_u0_n675 ) , .B2( u0_u0_n752 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U369 (.A2( u0_u0_n441 ) , .ZN( u0_u0_n605 ) , .A1( u0_u0_n821 ) );
  NOR3_X1 u0_u0_U37 (.ZN( u0_u0_n555 ) , .A2( u0_u0_n657 ) , .A1( u0_u0_n673 ) , .A3( u0_u0_n776 ) );
  NOR2_X1 u0_u0_U370 (.ZN( u0_u0_n537 ) , .A2( u0_u0_n785 ) , .A1( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U371 (.ZN( u0_u0_n525 ) , .A2( u0_u0_n705 ) , .A1( u0_u0_n821 ) );
  NAND2_X2 u0_u0_U372 (.A1( u0_u0_n461 ) , .A2( u0_u0_n477 ) , .ZN( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U373 (.A1( u0_u0_n675 ) , .ZN( u0_u0_n694 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U374 (.ZN( u0_u0_n564 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n821 ) );
  NAND2_X2 u0_u0_U375 (.A1( u0_u0_n459 ) , .A2( u0_u0_n467 ) , .ZN( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U376 (.ZN( u0_u0_n691 ) , .A1( u0_u0_n734 ) , .A2( u0_u0_n821 ) );
  INV_X1 u0_u0_U377 (.A( u0_u0_n821 ) , .ZN( u0_u0_n836 ) );
  NAND2_X1 u0_u0_U378 (.ZN( u0_u0_n677 ) , .A1( u0_u0_n811 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U379 (.ZN( u0_u0_n460 ) , .A1( u0_u0_n832 ) , .A2( w3_16 ) );
  AOI211_X1 u0_u0_U38 (.B( u0_u0_n545 ) , .A( u0_u0_n546 ) , .ZN( u0_u0_n557 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n856 ) );
  NOR2_X1 u0_u0_U380 (.ZN( u0_u0_n468 ) , .A2( w3_16 ) , .A1( w3_17 ) );
  INV_X1 u0_u0_U381 (.ZN( u0_u0_n831 ) , .A( w3_16 ) );
  AOI211_X1 u0_u0_U382 (.A( u0_u0_n643 ) , .ZN( u0_u0_n651 ) , .B( u0_u0_n748 ) , .C2( u0_u0_n844 ) , .C1( u0_u0_n859 ) );
  NAND4_X1 u0_u0_U383 (.A4( u0_u0_n639 ) , .A3( u0_u0_n640 ) , .A2( u0_u0_n641 ) , .A1( u0_u0_n642 ) , .ZN( u0_u0_n748 ) );
  AOI21_X1 u0_u0_U384 (.ZN( u0_u0_n582 ) , .B2( u0_u0_n729 ) , .B1( u0_u0_n753 ) , .A( u0_u0_n790 ) );
  NAND2_X2 u0_u0_U385 (.A2( u0_u0_n447 ) , .A1( u0_u0_n453 ) , .ZN( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U386 (.ZN( u0_u0_n466 ) , .A1( u0_u0_n854 ) , .A2( w3_23 ) );
  INV_X1 u0_u0_U387 (.ZN( u0_u0_n862 ) , .A( w3_23 ) );
  NOR2_X1 u0_u0_U388 (.ZN( u0_u0_n447 ) , .A2( w3_20 ) , .A1( w3_21 ) );
  NOR2_X1 u0_u0_U389 (.ZN( u0_u0_n454 ) , .A1( u0_u0_n852 ) , .A2( w3_21 ) );
  NOR4_X1 u0_u0_U39 (.A4( u0_u0_n550 ) , .A3( u0_u0_n551 ) , .A2( u0_u0_n552 ) , .A1( u0_u0_n553 ) , .ZN( u0_u0_n554 ) );
  OAI21_X1 u0_u0_U390 (.A( u0_u0_n736 ) , .B1( u0_u0_n737 ) , .ZN( u0_u0_n741 ) , .B2( u0_u0_n810 ) );
  OAI222_X1 u0_u0_U391 (.B2( u0_u0_n752 ) , .B1( u0_u0_n753 ) , .A2( u0_u0_n754 ) , .ZN( u0_u0_n762 ) , .C2( u0_u0_n810 ) , .C1( u0_u0_n819 ) , .A1( u0_u0_n822 ) );
  OAI22_X1 u0_u0_U392 (.B2( u0_u0_n808 ) , .B1( u0_u0_n809 ) , .A2( u0_u0_n810 ) , .A1( u0_u0_n811 ) , .ZN( u0_u0_n813 ) );
  OAI222_X1 u0_u0_U393 (.ZN( u0_u0_n511 ) , .C2( u0_u0_n631 ) , .B2( u0_u0_n653 ) , .B1( u0_u0_n752 ) , .A2( u0_u0_n753 ) , .C1( u0_u0_n810 ) , .A1( u0_u0_n811 ) );
  AOI21_X1 u0_u0_U394 (.ZN( u0_u0_n656 ) , .A( u0_u0_n784 ) , .B1( u0_u0_n797 ) , .B2( u0_u0_n810 ) );
  INV_X1 u0_u0_U395 (.A( u0_u0_n810 ) , .ZN( u0_u0_n864 ) );
  NOR2_X1 u0_u0_U396 (.ZN( u0_u0_n740 ) , .A2( u0_u0_n808 ) , .A1( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U397 (.ZN( u0_u0_n490 ) , .A1( u0_u0_n793 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U398 (.ZN( u0_u0_n573 ) , .A1( u0_u0_n752 ) , .A2( u0_u0_n810 ) );
  AOI21_X1 u0_u0_U399 (.A( u0_u0_n442 ) , .ZN( u0_u0_n558 ) , .B1( u0_u0_n675 ) , .B2( u0_u0_n810 ) );
  OR4_X1 u0_u0_U4 (.A4( u0_u0_n448 ) , .A2( u0_u0_n449 ) , .A1( u0_u0_n450 ) , .ZN( u0_u0_n451 ) , .A3( u0_u0_n559 ) );
  AOI221_X1 u0_u0_U40 (.A( u0_u0_n495 ) , .ZN( u0_u0_n500 ) , .B2( u0_u0_n841 ) , .C2( u0_u0_n846 ) , .C1( u0_u0_n856 ) , .B1( u0_u0_n864 ) );
  NAND2_X1 u0_u0_U400 (.ZN( u0_u0_n758 ) , .A1( u0_u0_n768 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U401 (.ZN( u0_u0_n720 ) , .A1( u0_u0_n810 ) , .A2( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U402 (.ZN( u0_u0_n562 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U403 (.ZN( u0_u0_n676 ) , .A1( u0_u0_n795 ) , .A2( u0_u0_n810 ) );
  NAND4_X1 u0_u0_U404 (.ZN( u0_subword_27 ) , .A2( u0_u0_n440 ) , .A4( u0_u0_n710 ) , .A3( u0_u0_n711 ) , .A1( u0_u0_n712 ) );
  OAI22_X1 u0_u0_U405 (.B2( u0_u0_n749 ) , .ZN( u0_u0_n751 ) , .A2( u0_u0_n767 ) , .B1( u0_u0_n785 ) , .A1( u0_u0_n797 ) );
  OAI22_X1 u0_u0_U406 (.B1( u0_u0_n441 ) , .ZN( u0_u0_n502 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n785 ) , .B2( u0_u0_n811 ) );
  NOR2_X1 u0_u0_U407 (.ZN( u0_u0_n522 ) , .A1( u0_u0_n713 ) , .A2( u0_u0_n749 ) );
  OAI22_X1 u0_u0_U408 (.ZN( u0_u0_n715 ) , .A2( u0_u0_n733 ) , .B2( u0_u0_n734 ) , .A1( u0_u0_n749 ) , .B1( u0_u0_n818 ) );
  NOR2_X1 u0_u0_U409 (.A2( u0_u0_n749 ) , .ZN( u0_u0_n774 ) , .A1( u0_u0_n817 ) );
  INV_X1 u0_u0_U41 (.A( u0_u0_n783 ) , .ZN( u0_u0_n871 ) );
  OAI22_X1 u0_u0_U410 (.B1( u0_u0_n446 ) , .ZN( u0_u0_n450 ) , .A2( u0_u0_n733 ) , .A1( u0_u0_n749 ) , .B2( u0_u0_n754 ) );
  NOR2_X1 u0_u0_U411 (.ZN( u0_u0_n553 ) , .A1( u0_u0_n705 ) , .A2( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U412 (.ZN( u0_u0_n536 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n797 ) );
  NOR2_X1 u0_u0_U413 (.A2( u0_u0_n749 ) , .ZN( u0_u0_n760 ) , .A1( u0_u0_n810 ) );
  NOR2_X1 u0_u0_U414 (.A1( u0_u0_n675 ) , .ZN( u0_u0_n679 ) , .A2( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U415 (.ZN( u0_u0_n723 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n749 ) );
  NOR2_X1 u0_u0_U416 (.ZN( u0_u0_n588 ) , .A1( u0_u0_n749 ) , .A2( u0_u0_n820 ) );
  INV_X1 u0_u0_U417 (.A( u0_u0_n749 ) , .ZN( u0_u0_n842 ) );
  NAND4_X1 u0_u0_U418 (.ZN( u0_subword_26 ) , .A4( u0_u0_n649 ) , .A3( u0_u0_n650 ) , .A1( u0_u0_n651 ) , .A2( u0_u0_n652 ) );
  OAI22_X1 u0_u0_U419 (.ZN( u0_u0_n594 ) , .A2( u0_u0_n752 ) , .B2( u0_u0_n767 ) , .A1( u0_u0_n768 ) , .B1( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U42 (.ZN( u0_u0_n686 ) , .A2( u0_u0_n839 ) , .A1( u0_u0_n844 ) );
  NAND2_X1 u0_u0_U420 (.A1( u0_u0_n734 ) , .A2( u0_u0_n789 ) , .ZN( u0_u0_n816 ) );
  AOI21_X1 u0_u0_U421 (.ZN( u0_u0_n598 ) , .B1( u0_u0_n733 ) , .B2( u0_u0_n789 ) , .A( u0_u0_n795 ) );
  AOI21_X1 u0_u0_U422 (.ZN( u0_u0_n654 ) , .A( u0_u0_n767 ) , .B2( u0_u0_n789 ) , .B1( u0_u0_n797 ) );
  AOI21_X1 u0_u0_U423 (.ZN( u0_u0_n629 ) , .B1( u0_u0_n705 ) , .A( u0_u0_n784 ) , .B2( u0_u0_n789 ) );
  OAI22_X1 u0_u0_U424 (.ZN( u0_u0_n687 ) , .A1( u0_u0_n705 ) , .A2( u0_u0_n735 ) , .B2( u0_u0_n789 ) , .B1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U425 (.ZN( u0_u0_n657 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n793 ) );
  OAI21_X1 u0_u0_U426 (.A( u0_u0_n619 ) , .ZN( u0_u0_n622 ) , .B1( u0_u0_n631 ) , .B2( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U427 (.ZN( u0_u0_n559 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n789 ) );
  NOR2_X1 u0_u0_U428 (.ZN( u0_u0_n616 ) , .A1( u0_u0_n789 ) , .A2( u0_u0_n821 ) );
  NOR2_X1 u0_u0_U429 (.A2( u0_u0_n442 ) , .ZN( u0_u0_n606 ) , .A1( u0_u0_n789 ) );
  NAND4_X1 u0_u0_U43 (.A4( u0_u0_n609 ) , .A3( u0_u0_n610 ) , .A2( u0_u0_n611 ) , .A1( u0_u0_n612 ) , .ZN( u0_u0_n727 ) );
  INV_X1 u0_u0_U430 (.A( u0_u0_n789 ) , .ZN( u0_u0_n865 ) );
  NOR2_X1 u0_u0_U431 (.ZN( u0_u0_n470 ) , .A2( w3_22 ) , .A1( w3_23 ) );
  NOR2_X1 u0_u0_U432 (.ZN( u0_u0_n458 ) , .A1( u0_u0_n862 ) , .A2( w3_22 ) );
  INV_X1 u0_u0_U433 (.ZN( u0_u0_n854 ) , .A( w3_22 ) );
  AOI21_X1 u0_u0_U434 (.A( u0_u0_n442 ) , .ZN( u0_u0_n506 ) , .B1( u0_u0_n713 ) , .B2( u0_u0_n791 ) );
  OAI22_X1 u0_u0_U435 (.ZN( u0_u0_n596 ) , .B1( u0_u0_n735 ) , .B2( u0_u0_n754 ) , .A2( u0_u0_n791 ) , .A1( u0_u0_n808 ) );
  NOR2_X1 u0_u0_U436 (.ZN( u0_u0_n659 ) , .A1( u0_u0_n767 ) , .A2( u0_u0_n791 ) );
  NAND3_X1 u0_u0_U437 (.ZN( u0_subword_30 ) , .A3( u0_u0_n802 ) , .A2( u0_u0_n803 ) , .A1( u0_u0_n804 ) );
  NAND3_X1 u0_u0_U438 (.ZN( u0_subword_29 ) , .A3( u0_u0_n763 ) , .A2( u0_u0_n764 ) , .A1( u0_u0_n765 ) );
  NAND3_X1 u0_u0_U439 (.ZN( u0_subword_28 ) , .A3( u0_u0_n743 ) , .A2( u0_u0_n744 ) , .A1( u0_u0_n745 ) );
  NOR4_X1 u0_u0_U44 (.A3( u0_u0_n606 ) , .A2( u0_u0_n607 ) , .A1( u0_u0_n608 ) , .ZN( u0_u0_n609 ) , .A4( u0_u0_n661 ) );
  NAND3_X1 u0_u0_U440 (.A3( u0_u0_n681 ) , .A2( u0_u0_n682 ) , .A1( u0_u0_n683 ) , .ZN( u0_u0_n812 ) );
  NAND3_X1 u0_u0_U441 (.ZN( u0_u0_n644 ) , .A3( u0_u0_n713 ) , .A2( u0_u0_n729 ) , .A1( u0_u0_n797 ) );
  NAND3_X1 u0_u0_U442 (.A3( u0_u0_n624 ) , .A2( u0_u0_n625 ) , .A1( u0_u0_n626 ) , .ZN( u0_u0_n730 ) );
  NAND3_X1 u0_u0_U443 (.A1( u0_u0_n591 ) , .A2( u0_u0_n592 ) , .A3( u0_u0_n593 ) , .ZN( u0_u0_n627 ) );
  NAND3_X1 u0_u0_U444 (.ZN( u0_u0_n571 ) , .A3( u0_u0_n686 ) , .A2( u0_u0_n755 ) , .A1( u0_u0_n790 ) );
  NAND3_X1 u0_u0_U445 (.A3( u0_u0_n529 ) , .A2( u0_u0_n530 ) , .A1( u0_u0_n531 ) , .ZN( u0_u0_n747 ) );
  NAND3_X1 u0_u0_U446 (.A3( u0_u0_n518 ) , .A1( u0_u0_n519 ) , .ZN( u0_u0_n614 ) , .A2( u0_u0_n875 ) );
  NAND3_X1 u0_u0_U447 (.A3( u0_u0_n473 ) , .A2( u0_u0_n474 ) , .A1( u0_u0_n475 ) , .ZN( u0_u0_n782 ) );
  NAND2_X1 u0_u0_U448 (.A2( u0_u0_n754 ) , .A1( u0_u0_n791 ) , .ZN( u0_u0_n814 ) );
  NOR2_X1 u0_u0_U449 (.A2( u0_u0_n443 ) , .ZN( u0_u0_n560 ) , .A1( u0_u0_n791 ) );
  NOR3_X1 u0_u0_U45 (.A1( u0_u0_n605 ) , .ZN( u0_u0_n610 ) , .A3( u0_u0_n669 ) , .A2( u0_u0_n775 ) );
  NOR2_X1 u0_u0_U450 (.ZN( u0_u0_n618 ) , .A1( u0_u0_n784 ) , .A2( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U451 (.ZN( u0_u0_n722 ) , .A2( u0_u0_n749 ) , .A1( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U452 (.ZN( u0_u0_n707 ) , .A2( u0_u0_n791 ) , .A1( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U453 (.A1( u0_u0_n735 ) , .ZN( u0_u0_n770 ) , .A2( u0_u0_n791 ) );
  NOR2_X1 u0_u0_U454 (.ZN( u0_u0_n455 ) , .A1( u0_u0_n853 ) , .A2( w3_20 ) );
  INV_X1 u0_u0_U455 (.ZN( u0_u0_n852 ) , .A( w3_20 ) );
  NAND4_X1 u0_u0_U46 (.A4( u0_u0_n566 ) , .A3( u0_u0_n567 ) , .A2( u0_u0_n568 ) , .A1( u0_u0_n569 ) , .ZN( u0_u0_n613 ) );
  NOR4_X1 u0_u0_U47 (.ZN( u0_u0_n567 ) , .A1( u0_u0_n659 ) , .A3( u0_u0_n667 ) , .A4( u0_u0_n691 ) , .A2( u0_u0_n773 ) );
  NOR4_X1 u0_u0_U48 (.A4( u0_u0_n558 ) , .A3( u0_u0_n559 ) , .A2( u0_u0_n560 ) , .A1( u0_u0_n561 ) , .ZN( u0_u0_n568 ) );
  NOR4_X1 u0_u0_U49 (.A4( u0_u0_n562 ) , .A3( u0_u0_n563 ) , .A2( u0_u0_n564 ) , .A1( u0_u0_n565 ) , .ZN( u0_u0_n566 ) );
  OR3_X1 u0_u0_U5 (.ZN( u0_u0_n22 ) , .A3( u0_u0_n658 ) , .A1( u0_u0_n668 ) , .A2( u0_u0_n772 ) );
  NOR4_X1 u0_u0_U50 (.A4( u0_u0_n693 ) , .A3( u0_u0_n694 ) , .A2( u0_u0_n695 ) , .A1( u0_u0_n696 ) , .ZN( u0_u0_n697 ) );
  INV_X1 u0_u0_U51 (.A( u0_u0_n685 ) , .ZN( u0_u0_n876 ) );
  NOR4_X1 u0_u0_U52 (.A4( u0_u0_n532 ) , .A2( u0_u0_n533 ) , .A1( u0_u0_n534 ) , .ZN( u0_u0_n544 ) , .A3( u0_u0_n707 ) );
  NOR4_X1 u0_u0_U53 (.A4( u0_u0_n535 ) , .A3( u0_u0_n536 ) , .ZN( u0_u0_n543 ) , .A2( u0_u0_n690 ) , .A1( u0_u0_n799 ) );
  NOR4_X1 u0_u0_U54 (.A4( u0_u0_n538 ) , .A3( u0_u0_n539 ) , .A2( u0_u0_n540 ) , .ZN( u0_u0_n541 ) , .A1( u0_u0_n825 ) );
  NOR4_X1 u0_u0_U55 (.A4( u0_u0_n520 ) , .A3( u0_u0_n521 ) , .A2( u0_u0_n522 ) , .A1( u0_u0_n523 ) , .ZN( u0_u0_n530 ) );
  NOR4_X1 u0_u0_U56 (.A3( u0_u0_n527 ) , .A1( u0_u0_n528 ) , .ZN( u0_u0_n529 ) , .A2( u0_u0_n679 ) , .A4( u0_u0_n774 ) );
  NOR4_X1 u0_u0_U57 (.A4( u0_u0_n476 ) , .ZN( u0_u0_n482 ) , .A3( u0_u0_n562 ) , .A1( u0_u0_n740 ) , .A2( u0_u0_n760 ) );
  NOR4_X1 u0_u0_U58 (.ZN( u0_u0_n481 ) , .A1( u0_u0_n537 ) , .A3( u0_u0_n574 ) , .A4( u0_u0_n606 ) , .A2( u0_u0_n648 ) );
  NOR4_X1 u0_u0_U59 (.ZN( u0_u0_n480 ) , .A1( u0_u0_n512 ) , .A3( u0_u0_n550 ) , .A2( u0_u0_n589 ) , .A4( u0_u0_n721 ) );
  OR2_X1 u0_u0_U6 (.ZN( u0_u0_n171 ) , .A2( u0_u0_n620 ) , .A1( u0_u0_n621 ) );
  NOR4_X1 u0_u0_U60 (.A4( u0_u0_n635 ) , .A3( u0_u0_n636 ) , .A2( u0_u0_n637 ) , .A1( u0_u0_n638 ) , .ZN( u0_u0_n639 ) );
  NOR4_X1 u0_u0_U61 (.A4( u0_u0_n632 ) , .A3( u0_u0_n633 ) , .A2( u0_u0_n634 ) , .ZN( u0_u0_n640 ) , .A1( u0_u0_n670 ) );
  AOI211_X1 u0_u0_U62 (.B( u0_u0_n629 ) , .A( u0_u0_n630 ) , .ZN( u0_u0_n641 ) , .C2( u0_u0_n841 ) , .C1( u0_u0_n867 ) );
  NAND4_X1 u0_u0_U63 (.A4( u0_u0_n777 ) , .A3( u0_u0_n778 ) , .A2( u0_u0_n779 ) , .A1( u0_u0_n780 ) , .ZN( u0_u0_n806 ) );
  NOR3_X1 u0_u0_U64 (.A3( u0_u0_n770 ) , .A2( u0_u0_n771 ) , .A1( u0_u0_n772 ) , .ZN( u0_u0_n778 ) );
  NOR4_X1 u0_u0_U65 (.A4( u0_u0_n773 ) , .A3( u0_u0_n774 ) , .A2( u0_u0_n775 ) , .A1( u0_u0_n776 ) , .ZN( u0_u0_n777 ) );
  NAND4_X1 u0_u0_U66 (.A4( u0_u0_n663 ) , .A3( u0_u0_n664 ) , .A2( u0_u0_n665 ) , .A1( u0_u0_n666 ) , .ZN( u0_u0_n805 ) );
  NOR3_X1 u0_u0_U67 (.A3( u0_u0_n654 ) , .A2( u0_u0_n655 ) , .A1( u0_u0_n656 ) , .ZN( u0_u0_n665 ) );
  NOR3_X1 u0_u0_U68 (.A3( u0_u0_n657 ) , .A2( u0_u0_n658 ) , .A1( u0_u0_n659 ) , .ZN( u0_u0_n664 ) );
  NOR3_X1 u0_u0_U69 (.A3( u0_u0_n660 ) , .A2( u0_u0_n661 ) , .A1( u0_u0_n662 ) , .ZN( u0_u0_n663 ) );
  OR2_X1 u0_u0_U7 (.ZN( u0_u0_n438 ) , .A1( u0_u0_n782 ) , .A2( u0_u0_n783 ) );
  NOR4_X1 u0_u0_U70 (.A4( u0_u0_n515 ) , .A2( u0_u0_n516 ) , .A1( u0_u0_n517 ) , .ZN( u0_u0_n518 ) , .A3( u0_u0_n676 ) );
  INV_X1 u0_u0_U71 (.A( u0_u0_n511 ) , .ZN( u0_u0_n875 ) );
  NOR2_X1 u0_u0_U72 (.ZN( u0_u0_n809 ) , .A1( u0_u0_n859 ) , .A2( u0_u0_n865 ) );
  NAND4_X1 u0_u0_U73 (.A4( u0_u0_n491 ) , .A3( u0_u0_n492 ) , .A2( u0_u0_n493 ) , .A1( u0_u0_n494 ) , .ZN( u0_u0_n783 ) );
  NOR4_X1 u0_u0_U74 (.A4( u0_u0_n490 ) , .ZN( u0_u0_n493 ) , .A1( u0_u0_n572 ) , .A2( u0_u0_n587 ) , .A3( u0_u0_n608 ) );
  NOR4_X1 u0_u0_U75 (.ZN( u0_u0_n492 ) , .A1( u0_u0_n513 ) , .A2( u0_u0_n525 ) , .A4( u0_u0_n552 ) , .A3( u0_u0_n617 ) );
  NAND4_X1 u0_u0_U76 (.A4( u0_u0_n462 ) , .A3( u0_u0_n463 ) , .A2( u0_u0_n464 ) , .A1( u0_u0_n465 ) , .ZN( u0_u0_n685 ) );
  NOR3_X1 u0_u0_U77 (.ZN( u0_u0_n463 ) , .A3( u0_u0_n536 ) , .A1( u0_u0_n561 ) , .A2( u0_u0_n576 ) );
  AOI221_X1 u0_u0_U78 (.A( u0_u0_n456 ) , .ZN( u0_u0_n465 ) , .C2( u0_u0_n758 ) , .B1( u0_u0_n837 ) , .C1( u0_u0_n847 ) , .B2( u0_u0_n865 ) );
  NOR4_X1 u0_u0_U79 (.ZN( u0_u0_n464 ) , .A2( u0_u0_n515 ) , .A1( u0_u0_n605 ) , .A4( u0_u0_n634 ) , .A3( u0_u0_n716 ) );
  NAND2_X2 u0_u0_U8 (.A2( u0_u0_n477 ) , .A1( u0_u0_n478 ) , .ZN( u0_u0_n822 ) );
  NOR2_X1 u0_u0_U80 (.ZN( u0_u0_n766 ) , .A1( u0_u0_n838 ) , .A2( u0_u0_n839 ) );
  NOR2_X1 u0_u0_U81 (.ZN( u0_u0_n631 ) , .A2( u0_u0_n841 ) , .A1( u0_u0_n844 ) );
  NAND4_X1 u0_u0_U82 (.A4( u0_u0_n485 ) , .A3( u0_u0_n486 ) , .A2( u0_u0_n487 ) , .A1( u0_u0_n488 ) , .ZN( u0_u0_n700 ) );
  NOR3_X1 u0_u0_U83 (.ZN( u0_u0_n486 ) , .A2( u0_u0_n514 ) , .A3( u0_u0_n607 ) , .A1( u0_u0_n616 ) );
  NOR4_X1 u0_u0_U84 (.ZN( u0_u0_n487 ) , .A3( u0_u0_n538 ) , .A4( u0_u0_n551 ) , .A2( u0_u0_n573 ) , .A1( u0_u0_n722 ) );
  AOI211_X1 u0_u0_U85 (.B( u0_u0_n483 ) , .A( u0_u0_n484 ) , .ZN( u0_u0_n488 ) , .C2( u0_u0_n838 ) , .C1( u0_u0_n865 ) );
  AOI222_X1 u0_u0_U86 (.A2( u0_u0_n444 ) , .ZN( u0_u0_n475 ) , .B1( u0_u0_n837 ) , .A1( u0_u0_n844 ) , .C1( u0_u0_n847 ) , .C2( u0_u0_n856 ) , .B2( u0_u0_n869 ) );
  NOR4_X1 u0_u0_U87 (.A1( u0_u0_n472 ) , .ZN( u0_u0_n473 ) , .A4( u0_u0_n548 ) , .A2( u0_u0_n560 ) , .A3( u0_u0_n620 ) );
  AOI221_X1 u0_u0_U88 (.ZN( u0_u0_n474 ) , .C2( u0_u0_n719 ) , .B2( u0_u0_n836 ) , .C1( u0_u0_n850 ) , .B1( u0_u0_n864 ) , .A( u0_u0_n868 ) );
  NAND4_X1 u0_u0_U89 (.A4( u0_u0_n724 ) , .A3( u0_u0_n725 ) , .A2( u0_u0_n726 ) , .ZN( u0_u0_n746 ) , .A1( u0_u0_n861 ) );
  CLKBUF_X1 u0_u0_U9 (.Z( u0_u0_n439 ) , .A( u0_u0_n850 ) );
  INV_X1 u0_u0_U90 (.A( u0_u0_n714 ) , .ZN( u0_u0_n861 ) );
  NOR4_X1 u0_u0_U91 (.A4( u0_u0_n720 ) , .A3( u0_u0_n721 ) , .A2( u0_u0_n722 ) , .A1( u0_u0_n723 ) , .ZN( u0_u0_n724 ) );
  AOI221_X1 u0_u0_U92 (.B2( u0_u0_n439 ) , .A( u0_u0_n715 ) , .ZN( u0_u0_n726 ) , .C2( u0_u0_n849 ) , .C1( u0_u0_n865 ) , .B1( u0_u0_n866 ) );
  NAND4_X1 u0_u0_U93 (.A4( u0_u0_n579 ) , .A3( u0_u0_n580 ) , .A1( u0_u0_n581 ) , .ZN( u0_u0_n728 ) , .A2( u0_u0_n878 ) );
  AOI221_X1 u0_u0_U94 (.A( u0_u0_n570 ) , .C2( u0_u0_n571 ) , .ZN( u0_u0_n580 ) , .B2( u0_u0_n850 ) , .B1( u0_u0_n857 ) , .C1( u0_u0_n858 ) );
  NOR4_X1 u0_u0_U95 (.A4( u0_u0_n575 ) , .A3( u0_u0_n576 ) , .A2( u0_u0_n577 ) , .A1( u0_u0_n578 ) , .ZN( u0_u0_n579 ) );
  INV_X1 u0_u0_U96 (.A( u0_u0_n613 ) , .ZN( u0_u0_n878 ) );
  NOR4_X1 u0_u0_U97 (.A4( u0_u0_n615 ) , .A3( u0_u0_n616 ) , .A2( u0_u0_n617 ) , .A1( u0_u0_n618 ) , .ZN( u0_u0_n625 ) );
  NOR4_X1 u0_u0_U98 (.ZN( u0_u0_n626 ) , .A1( u0_u0_n662 ) , .A3( u0_u0_n672 ) , .A4( u0_u0_n688 ) , .A2( u0_u0_n771 ) );
  NOR2_X1 u0_u0_U99 (.ZN( u0_u0_n692 ) , .A1( u0_u0_n836 ) , .A2( u0_u0_n837 ) );
  DFF_X1 u0_w_reg_0_0 (.CK( clk ) , .D( u0_N42 ) , .Q( w0_0 ) );
  DFF_X1 u0_w_reg_0_1 (.CK( clk ) , .D( u0_N43 ) , .Q( w0_1 ) );
  DFF_X1 u0_w_reg_0_10 (.CK( clk ) , .D( u0_N52 ) , .Q( w0_10 ) );
  DFF_X1 u0_w_reg_0_11 (.CK( clk ) , .D( u0_N53 ) , .Q( w0_11 ) );
  DFF_X1 u0_w_reg_0_12 (.CK( clk ) , .D( u0_N54 ) , .Q( w0_12 ) );
  DFF_X1 u0_w_reg_0_13 (.CK( clk ) , .D( u0_N55 ) , .Q( w0_13 ) );
  DFF_X1 u0_w_reg_0_14 (.CK( clk ) , .D( u0_N56 ) , .Q( w0_14 ) );
  DFF_X1 u0_w_reg_0_15 (.CK( clk ) , .D( u0_N57 ) , .Q( w0_15 ) );
  DFF_X1 u0_w_reg_0_16 (.CK( clk ) , .D( u0_N58 ) , .Q( w0_16 ) );
  DFF_X1 u0_w_reg_0_17 (.CK( clk ) , .D( u0_N59 ) , .Q( w0_17 ) );
  DFF_X1 u0_w_reg_0_18 (.CK( clk ) , .D( u0_N60 ) , .Q( w0_18 ) );
  DFF_X1 u0_w_reg_0_19 (.CK( clk ) , .D( u0_N61 ) , .Q( w0_19 ) );
  DFF_X1 u0_w_reg_0_2 (.CK( clk ) , .D( u0_N44 ) , .Q( w0_2 ) );
  DFF_X1 u0_w_reg_0_20 (.CK( clk ) , .D( u0_N62 ) , .Q( w0_20 ) );
  DFF_X1 u0_w_reg_0_21 (.CK( clk ) , .D( u0_N63 ) , .Q( w0_21 ) );
  DFF_X1 u0_w_reg_0_22 (.CK( clk ) , .D( u0_N64 ) , .Q( w0_22 ) );
  DFF_X1 u0_w_reg_0_23 (.CK( clk ) , .D( u0_N65 ) , .Q( w0_23 ) );
  DFF_X1 u0_w_reg_0_24 (.CK( clk ) , .D( u0_N66 ) , .Q( w0_24 ) );
  DFF_X1 u0_w_reg_0_25 (.CK( clk ) , .D( u0_N67 ) , .Q( w0_25 ) );
  DFF_X1 u0_w_reg_0_26 (.CK( clk ) , .D( u0_N68 ) , .Q( w0_26 ) );
  DFF_X1 u0_w_reg_0_27 (.CK( clk ) , .D( u0_N69 ) , .Q( w0_27 ) );
  DFF_X1 u0_w_reg_0_28 (.CK( clk ) , .D( u0_N70 ) , .Q( w0_28 ) );
  DFF_X1 u0_w_reg_0_29 (.CK( clk ) , .D( u0_N71 ) , .Q( w0_29 ) );
  DFF_X1 u0_w_reg_0_3 (.CK( clk ) , .D( u0_N45 ) , .Q( w0_3 ) );
  DFF_X1 u0_w_reg_0_30 (.CK( clk ) , .D( u0_N72 ) , .Q( w0_30 ) );
  DFF_X1 u0_w_reg_0_31 (.CK( clk ) , .D( u0_N73 ) , .Q( w0_31 ) );
  DFF_X1 u0_w_reg_0_4 (.CK( clk ) , .D( u0_N46 ) , .Q( w0_4 ) );
  DFF_X1 u0_w_reg_0_5 (.CK( clk ) , .D( u0_N47 ) , .Q( w0_5 ) );
  DFF_X1 u0_w_reg_0_6 (.CK( clk ) , .D( u0_N48 ) , .Q( w0_6 ) );
  DFF_X1 u0_w_reg_0_7 (.CK( clk ) , .D( u0_N49 ) , .Q( w0_7 ) );
  DFF_X1 u0_w_reg_0_8 (.CK( clk ) , .D( u0_N50 ) , .Q( w0_8 ) );
  DFF_X1 u0_w_reg_0_9 (.CK( clk ) , .D( u0_N51 ) , .Q( w0_9 ) );
  DFF_X1 u0_w_reg_1_0 (.CK( clk ) , .D( u0_N108 ) , .Q( w1_0 ) );
  DFF_X1 u0_w_reg_1_1 (.CK( clk ) , .D( u0_N109 ) , .Q( w1_1 ) );
  DFF_X1 u0_w_reg_1_10 (.CK( clk ) , .D( u0_N118 ) , .Q( w1_10 ) );
  DFF_X1 u0_w_reg_1_11 (.CK( clk ) , .D( u0_N119 ) , .Q( w1_11 ) );
  DFF_X1 u0_w_reg_1_12 (.CK( clk ) , .D( u0_N120 ) , .Q( w1_12 ) );
  DFF_X1 u0_w_reg_1_13 (.CK( clk ) , .D( u0_N121 ) , .Q( w1_13 ) );
  DFF_X1 u0_w_reg_1_14 (.CK( clk ) , .D( u0_N122 ) , .Q( w1_14 ) );
  DFF_X1 u0_w_reg_1_15 (.CK( clk ) , .D( u0_N123 ) , .Q( w1_15 ) );
  DFF_X1 u0_w_reg_1_16 (.CK( clk ) , .D( u0_N124 ) , .Q( w1_16 ) );
  DFF_X1 u0_w_reg_1_17 (.CK( clk ) , .D( u0_N125 ) , .Q( w1_17 ) );
  DFF_X1 u0_w_reg_1_18 (.CK( clk ) , .D( u0_N126 ) , .Q( w1_18 ) );
  DFF_X1 u0_w_reg_1_19 (.CK( clk ) , .D( u0_N127 ) , .Q( w1_19 ) );
  DFF_X1 u0_w_reg_1_2 (.CK( clk ) , .D( u0_N110 ) , .Q( w1_2 ) );
  DFF_X1 u0_w_reg_1_20 (.CK( clk ) , .D( u0_N128 ) , .Q( w1_20 ) );
  DFF_X1 u0_w_reg_1_21 (.CK( clk ) , .D( u0_N129 ) , .Q( w1_21 ) );
  DFF_X1 u0_w_reg_1_22 (.CK( clk ) , .D( u0_N130 ) , .Q( w1_22 ) );
  DFF_X1 u0_w_reg_1_23 (.CK( clk ) , .D( u0_N131 ) , .Q( w1_23 ) );
  DFF_X1 u0_w_reg_1_24 (.CK( clk ) , .D( u0_N132 ) , .Q( w1_24 ) );
  DFF_X1 u0_w_reg_1_25 (.CK( clk ) , .D( u0_N133 ) , .Q( w1_25 ) );
  DFF_X1 u0_w_reg_1_26 (.CK( clk ) , .D( u0_N134 ) , .QN( u0_n242 ) , .Q( w1_26 ) );
  DFF_X1 u0_w_reg_1_27 (.CK( clk ) , .D( u0_N135 ) , .Q( w1_27 ) );
  DFF_X1 u0_w_reg_1_28 (.CK( clk ) , .D( u0_N136 ) , .Q( w1_28 ) );
  DFF_X1 u0_w_reg_1_29 (.CK( clk ) , .D( u0_N137 ) , .Q( w1_29 ) );
  DFF_X1 u0_w_reg_1_3 (.CK( clk ) , .D( u0_N111 ) , .Q( w1_3 ) );
  DFF_X1 u0_w_reg_1_30 (.CK( clk ) , .D( u0_N138 ) , .QN( u0_n262 ) , .Q( w1_30 ) );
  DFF_X1 u0_w_reg_1_31 (.CK( clk ) , .D( u0_N139 ) , .Q( w1_31 ) );
  DFF_X1 u0_w_reg_1_4 (.CK( clk ) , .D( u0_N112 ) , .Q( w1_4 ) );
  DFF_X1 u0_w_reg_1_5 (.CK( clk ) , .D( u0_N113 ) , .Q( w1_5 ) );
  DFF_X1 u0_w_reg_1_6 (.CK( clk ) , .D( u0_N114 ) , .Q( w1_6 ) );
  DFF_X1 u0_w_reg_1_7 (.CK( clk ) , .D( u0_N115 ) , .Q( w1_7 ) );
  DFF_X1 u0_w_reg_1_8 (.CK( clk ) , .D( u0_N116 ) , .Q( w1_8 ) );
  DFF_X1 u0_w_reg_1_9 (.CK( clk ) , .D( u0_N117 ) , .Q( w1_9 ) );
  DFF_X1 u0_w_reg_2_0 (.CK( clk ) , .D( u0_N174 ) , .Q( w2_0 ) );
  DFF_X1 u0_w_reg_2_1 (.CK( clk ) , .D( u0_N175 ) , .Q( w2_1 ) );
  DFF_X1 u0_w_reg_2_10 (.CK( clk ) , .D( u0_N184 ) , .Q( w2_10 ) );
  DFF_X1 u0_w_reg_2_11 (.CK( clk ) , .D( u0_N185 ) , .Q( w2_11 ) );
  DFF_X1 u0_w_reg_2_12 (.CK( clk ) , .D( u0_N186 ) , .Q( w2_12 ) );
  DFF_X1 u0_w_reg_2_13 (.CK( clk ) , .D( u0_N187 ) , .Q( w2_13 ) );
  DFF_X1 u0_w_reg_2_14 (.CK( clk ) , .D( u0_N188 ) , .Q( w2_14 ) );
  DFF_X1 u0_w_reg_2_15 (.CK( clk ) , .D( u0_N189 ) , .Q( w2_15 ) );
  DFF_X1 u0_w_reg_2_16 (.CK( clk ) , .D( u0_N190 ) , .Q( w2_16 ) );
  DFF_X1 u0_w_reg_2_17 (.CK( clk ) , .D( u0_N191 ) , .Q( w2_17 ) );
  DFF_X1 u0_w_reg_2_18 (.CK( clk ) , .D( u0_N192 ) , .Q( w2_18 ) );
  DFF_X1 u0_w_reg_2_19 (.CK( clk ) , .D( u0_N193 ) , .Q( w2_19 ) );
  DFF_X1 u0_w_reg_2_2 (.CK( clk ) , .D( u0_N176 ) , .Q( w2_2 ) );
  DFF_X1 u0_w_reg_2_20 (.CK( clk ) , .D( u0_N194 ) , .Q( w2_20 ) );
  DFF_X1 u0_w_reg_2_21 (.CK( clk ) , .D( u0_N195 ) , .Q( w2_21 ) );
  DFF_X1 u0_w_reg_2_22 (.CK( clk ) , .D( u0_N196 ) , .Q( w2_22 ) );
  DFF_X1 u0_w_reg_2_23 (.CK( clk ) , .D( u0_N197 ) , .Q( w2_23 ) );
  DFF_X1 u0_w_reg_2_24 (.CK( clk ) , .D( u0_N198 ) , .Q( w2_24 ) );
  DFF_X1 u0_w_reg_2_25 (.CK( clk ) , .D( u0_N199 ) , .Q( w2_25 ) );
  DFF_X1 u0_w_reg_2_26 (.CK( clk ) , .D( u0_N200 ) , .QN( u0_n244 ) , .Q( w2_26 ) );
  DFF_X1 u0_w_reg_2_27 (.CK( clk ) , .D( u0_N201 ) , .Q( w2_27 ) );
  DFF_X1 u0_w_reg_2_28 (.CK( clk ) , .D( u0_N202 ) , .Q( w2_28 ) );
  DFF_X1 u0_w_reg_2_29 (.CK( clk ) , .D( u0_N203 ) , .Q( w2_29 ) );
  DFF_X1 u0_w_reg_2_3 (.CK( clk ) , .D( u0_N177 ) , .Q( w2_3 ) );
  DFF_X1 u0_w_reg_2_30 (.CK( clk ) , .D( u0_N204 ) , .Q( w2_30 ) );
  DFF_X1 u0_w_reg_2_31 (.CK( clk ) , .D( u0_N205 ) , .Q( w2_31 ) );
  DFF_X1 u0_w_reg_2_4 (.CK( clk ) , .D( u0_N178 ) , .Q( w2_4 ) );
  DFF_X1 u0_w_reg_2_5 (.CK( clk ) , .D( u0_N179 ) , .Q( w2_5 ) );
  DFF_X1 u0_w_reg_2_6 (.CK( clk ) , .D( u0_N180 ) , .Q( w2_6 ) );
  DFF_X1 u0_w_reg_2_7 (.CK( clk ) , .D( u0_N181 ) , .Q( w2_7 ) );
  DFF_X1 u0_w_reg_2_8 (.CK( clk ) , .D( u0_N182 ) , .Q( w2_8 ) );
  DFF_X1 u0_w_reg_2_9 (.CK( clk ) , .D( u0_N183 ) , .Q( w2_9 ) );
  DFF_X1 u0_w_reg_3_0 (.CK( clk ) , .D( u0_N240 ) , .Q( w3_0 ) );
  DFF_X1 u0_w_reg_3_1 (.CK( clk ) , .D( u0_N241 ) , .Q( w3_1 ) );
  DFF_X1 u0_w_reg_3_10 (.CK( clk ) , .D( u0_N250 ) , .Q( w3_10 ) );
  DFF_X1 u0_w_reg_3_11 (.CK( clk ) , .D( u0_N251 ) , .Q( w3_11 ) );
  DFF_X1 u0_w_reg_3_12 (.CK( clk ) , .D( u0_N252 ) , .QN( u0_n258 ) , .Q( u0_n274 ) );
  DFF_X1 u0_w_reg_3_13 (.CK( clk ) , .D( u0_N253 ) , .QN( u0_n250 ) , .Q( u0_n272 ) );
  DFF_X1 u0_w_reg_3_14 (.CK( clk ) , .D( u0_N254 ) , .QN( u0_n254 ) , .Q( u0_n270 ) );
  DFF_X1 u0_w_reg_3_15 (.CK( clk ) , .D( u0_N255 ) , .QN( u0_n264 ) , .Q( u0_n268 ) );
  DFF_X1 u0_w_reg_3_16 (.CK( clk ) , .D( u0_N256 ) , .Q( w3_16 ) );
  DFF_X1 u0_w_reg_3_17 (.CK( clk ) , .D( u0_N257 ) , .Q( w3_17 ) );
  DFF_X1 u0_w_reg_3_18 (.CK( clk ) , .D( u0_N258 ) , .Q( w3_18 ) );
  DFF_X1 u0_w_reg_3_19 (.CK( clk ) , .D( u0_N259 ) , .Q( w3_19 ) );
  DFF_X1 u0_w_reg_3_2 (.CK( clk ) , .D( u0_N242 ) , .Q( w3_2 ) );
  DFF_X1 u0_w_reg_3_20 (.CK( clk ) , .D( u0_N260 ) , .Q( w3_20 ) );
  DFF_X1 u0_w_reg_3_21 (.CK( clk ) , .D( u0_N261 ) , .Q( w3_21 ) );
  DFF_X1 u0_w_reg_3_22 (.CK( clk ) , .D( u0_N262 ) , .Q( w3_22 ) );
  DFF_X1 u0_w_reg_3_23 (.CK( clk ) , .D( u0_N263 ) , .Q( w3_23 ) );
  DFF_X1 u0_w_reg_3_24 (.CK( clk ) , .D( u0_N264 ) , .QN( u0_n248 ) , .Q( w3_24 ) );
  DFF_X1 u0_w_reg_3_25 (.CK( clk ) , .D( u0_N265 ) , .Q( w3_25 ) );
  DFF_X1 u0_w_reg_3_26 (.CK( clk ) , .D( u0_N266 ) , .Q( w3_26 ) );
  DFF_X1 u0_w_reg_3_27 (.CK( clk ) , .D( u0_N267 ) , .Q( w3_27 ) );
  DFF_X1 u0_w_reg_3_28 (.CK( clk ) , .D( u0_N268 ) , .Q( w3_28 ) );
  DFF_X1 u0_w_reg_3_29 (.CK( clk ) , .D( u0_N269 ) , .Q( w3_29 ) );
  DFF_X1 u0_w_reg_3_3 (.CK( clk ) , .D( u0_N243 ) , .Q( w3_3 ) );
  DFF_X1 u0_w_reg_3_30 (.CK( clk ) , .D( u0_N270 ) , .Q( w3_30 ) );
  DFF_X1 u0_w_reg_3_31 (.CK( clk ) , .D( u0_N271 ) , .Q( w3_31 ) );
  DFF_X1 u0_w_reg_3_4 (.CK( clk ) , .D( u0_N244 ) , .Q( w3_4 ) );
  DFF_X1 u0_w_reg_3_5 (.CK( clk ) , .D( u0_N245 ) , .Q( w3_5 ) );
  DFF_X1 u0_w_reg_3_6 (.CK( clk ) , .D( u0_N246 ) , .Q( w3_6 ) );
  DFF_X1 u0_w_reg_3_7 (.CK( clk ) , .D( u0_N247 ) , .Q( w3_7 ) );
  DFF_X1 u0_w_reg_3_8 (.CK( clk ) , .D( u0_N248 ) , .Q( w3_8 ) );
  DFF_X1 u0_w_reg_3_9 (.CK( clk ) , .D( u0_N249 ) , .Q( w3_9 ) );
endmodule
