module des_des_die_15 ( u0_FP_33, u0_FP_34, u0_FP_35, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, u0_FP_41, 
       u0_FP_64, u0_K16_4, u0_K16_8, u0_K4_43, u0_K4_48, u0_K6_11, u0_K6_13, u0_K6_16, u0_K8_1, 
       u0_K8_11, u0_L14_13, u0_L14_17, u0_L14_18, u0_L14_2, u0_L14_23, u0_L14_28, u0_L14_31, u0_L14_9, 
       u0_L2_12, u0_L2_15, u0_L2_21, u0_L2_22, u0_L2_27, u0_L2_32, u0_L2_5, u0_L2_7, u0_L4_13, 
       u0_L4_16, u0_L4_17, u0_L4_18, u0_L4_2, u0_L4_23, u0_L4_24, u0_L4_28, u0_L4_30, u0_L4_31, 
       u0_L4_6, u0_L4_9, u0_L6_13, u0_L6_17, u0_L6_18, u0_L6_2, u0_L6_23, u0_L6_28, u0_L6_31, 
       u0_L6_9, u0_R2_1, u0_R2_24, u0_R2_25, u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_30, 
       u0_R2_31, u0_R2_32, u0_R4_1, u0_R4_10, u0_R4_11, u0_R4_12, u0_R4_13, u0_R4_2, u0_R4_3, 
       u0_R4_32, u0_R4_4, u0_R4_5, u0_R4_6, u0_R4_7, u0_R4_8, u0_R4_9, u0_R6_1, u0_R6_2, 
       u0_R6_3, u0_R6_32, u0_R6_4, u0_R6_5, u0_R6_6, u0_R6_7, u0_R6_8, u0_R6_9, u0_key_r_44, 
       u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_39, u0_uk_K_r2_50, u0_uk_K_r4_3, u0_uk_K_r4_33, u0_uk_K_r4_4, u0_uk_K_r4_41, u0_uk_K_r4_47, 
       u0_uk_K_r4_54, u0_uk_K_r4_55, u0_uk_K_r6_10, u0_uk_K_r6_19, u0_uk_K_r6_27, u0_uk_K_r6_3, u0_uk_K_r6_53, u0_uk_n10, u0_uk_n100, 
       u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n141, u0_uk_n142, u0_uk_n145, 
       u0_uk_n146, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, 
       u0_uk_n202, u0_uk_n207, u0_uk_n223, u0_uk_n240, u0_uk_n242, u0_uk_n251, u0_uk_n252, u0_uk_n257, u0_uk_n27, 
       u0_uk_n31, u0_uk_n318, u0_uk_n324, u0_uk_n330, u0_uk_n337, u0_uk_n339, u0_uk_n343, u0_uk_n344, u0_uk_n350, 
       u0_uk_n351, u0_uk_n352, u0_uk_n356, u0_uk_n358, u0_uk_n410, u0_uk_n414, u0_uk_n423, u0_uk_n426, u0_uk_n427, 
       u0_uk_n432, u0_uk_n435, u0_uk_n436, u0_uk_n441, u0_uk_n442, u0_uk_n448, u0_uk_n498, u0_uk_n499, u0_uk_n505, 
       u0_uk_n506, u0_uk_n508, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n521, u0_uk_n522, u0_uk_n527, u0_uk_n528, 
       u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n60, u0_uk_n63, u0_uk_n630, u0_uk_n636, u0_uk_n637, u0_uk_n639, 
       u0_uk_n640, u0_uk_n644, u0_uk_n646, u0_uk_n651, u0_uk_n652, u0_uk_n659, u0_uk_n660, u0_uk_n664, u0_uk_n667, 
       u0_uk_n668, u0_uk_n785, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n83, u0_uk_n92, u0_uk_n93, u1_L0_15, 
       u1_L0_21, u1_L0_27, u1_L0_5, u1_L5_1, u1_L5_10, u1_L5_20, u1_L5_26, u1_R0_1, u1_R0_28, 
       u1_R0_29, u1_R0_30, u1_R0_31, u1_R0_32, u1_R5_12, u1_R5_13, u1_R5_14, u1_R5_15, u1_R5_16, 
       u1_R5_17, u1_uk_K_r0_2, u1_uk_K_r0_52, u1_uk_K_r5_13, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_40, u1_uk_K_r5_5, u1_uk_K_r5_53, 
       u1_uk_n10, u1_uk_n11, u1_uk_n1266, u1_uk_n1271, u1_uk_n1276, u1_uk_n1281, u1_uk_n1282, u1_uk_n1286, u1_uk_n1293, 
       u1_uk_n1303, u1_uk_n1304, u1_uk_n145, u1_uk_n1483, u1_uk_n1495, u1_uk_n1498, u1_uk_n1505, u1_uk_n1526, u1_uk_n155, 
       u1_uk_n162, u1_uk_n17, u1_uk_n187, u1_uk_n191, u1_uk_n207, u1_uk_n217, u1_uk_n222, u1_uk_n231, u1_uk_n240, 
       u1_uk_n271, u1_uk_n297, u1_uk_n298, u1_uk_n60, u1_uk_n92, u2_K11_45, u2_K11_48, u2_K14_10, u2_K14_11, 
       u2_K14_12, u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_3, u2_K14_39, u2_K14_42, 
       u2_K14_6, u2_K14_8, u2_K15_28, u2_K15_29, u2_K15_31, u2_K15_34, u2_K15_35, u2_K15_39, u2_K3_7, 
       u2_K4_14, u2_K4_21, u2_K4_22, u2_K8_8, u2_K9_15, u2_K9_3, u2_K9_5, u2_L12_11, u2_L12_12, 
       u2_L12_13, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_19, u2_L12_2, u2_L12_22, u2_L12_23, u2_L12_24, 
       u2_L12_28, u2_L12_29, u2_L12_30, u2_L12_31, u2_L12_32, u2_L12_4, u2_L12_6, u2_L12_7, u2_L12_9, 
       u2_L13_11, u2_L13_12, u2_L13_14, u2_L13_15, u2_L13_19, u2_L13_21, u2_L13_22, u2_L13_25, u2_L13_27, 
       u2_L13_29, u2_L13_3, u2_L13_32, u2_L13_4, u2_L13_5, u2_L13_7, u2_L13_8, u2_L1_13, u2_L1_18, 
       u2_L1_2, u2_L1_28, u2_L2_1, u2_L2_10, u2_L2_16, u2_L2_20, u2_L2_24, u2_L2_26, u2_L2_30, 
       u2_L2_6, u2_L6_13, u2_L6_18, u2_L6_2, u2_L6_28, u2_L7_13, u2_L7_16, u2_L7_17, u2_L7_18, 
       u2_L7_2, u2_L7_23, u2_L7_24, u2_L7_28, u2_L7_30, u2_L7_31, u2_L7_6, u2_L7_9, u2_L9_15, 
       u2_L9_21, u2_L9_27, u2_L9_5, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_2, 
       u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R12_26, u2_R12_27, u2_R12_28, 
       u2_R12_29, u2_R12_3, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, 
       u2_R13_1, u2_R13_16, u2_R13_17, u2_R13_18, u2_R13_19, u2_R13_20, u2_R13_21, u2_R13_22, u2_R13_23, 
       u2_R13_24, u2_R13_25, u2_R13_26, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_30, u2_R13_31, u2_R13_32, 
       u2_R1_4, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_10, u2_R2_11, u2_R2_12, 
       u2_R2_13, u2_R2_14, u2_R2_15, u2_R2_16, u2_R2_17, u2_R2_8, u2_R2_9, u2_R6_4, u2_R6_5, 
       u2_R6_6, u2_R6_7, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_10, u2_R7_11, u2_R7_12, u2_R7_13, 
       u2_R7_2, u2_R7_3, u2_R7_32, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, 
       u2_R9_1, u2_R9_28, u2_R9_29, u2_R9_30, u2_R9_31, u2_R9_32, u2_key_r_1, u2_key_r_49, u2_uk_K_r11_33, 
       u2_uk_K_r12_1, u2_uk_K_r12_10, u2_uk_K_r12_30, u2_uk_K_r12_36, u2_uk_K_r12_7, u2_uk_K_r13_0, u2_uk_K_r13_22, u2_uk_K_r13_38, u2_uk_K_r1_18, 
       u2_uk_K_r2_18, u2_uk_K_r2_27, u2_uk_K_r2_50, u2_uk_K_r2_55, u2_uk_K_r6_3, u2_uk_K_r6_53, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, 
       u2_uk_K_r7_39, u2_uk_K_r7_46, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r9_15, u2_uk_K_r9_23, u2_uk_n1022, u2_uk_n1024, u2_uk_n1097, 
       u2_uk_n11, u2_uk_n110, u2_uk_n1119, u2_uk_n1120, u2_uk_n1121, u2_uk_n1125, u2_uk_n1130, u2_uk_n1141, u2_uk_n118, 
       u2_uk_n1280, u2_uk_n1285, u2_uk_n1286, u2_uk_n129, u2_uk_n1291, u2_uk_n1295, u2_uk_n1296, u2_uk_n1306, u2_uk_n1311, 
       u2_uk_n1322, u2_uk_n1324, u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1335, u2_uk_n1339, u2_uk_n1347, u2_uk_n1348, 
       u2_uk_n1356, u2_uk_n1363, u2_uk_n147, u2_uk_n1500, u2_uk_n1502, u2_uk_n1506, u2_uk_n1508, u2_uk_n1519, u2_uk_n1521, 
       u2_uk_n1535, u2_uk_n1543, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n155, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, 
       u2_uk_n1568, u2_uk_n1573, u2_uk_n1574, u2_uk_n1580, u2_uk_n163, u2_uk_n1632, u2_uk_n164, u2_uk_n1653, u2_uk_n1673, 
       u2_uk_n1674, u2_uk_n1769, u2_uk_n1770, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1781, u2_uk_n1783, 
       u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1791, u2_uk_n1793, u2_uk_n1794, u2_uk_n1796, u2_uk_n1797, u2_uk_n1801, 
       u2_uk_n1803, u2_uk_n1805, u2_uk_n1807, u2_uk_n1808, u2_uk_n1811, u2_uk_n1817, u2_uk_n1818, u2_uk_n1819, u2_uk_n182, 
       u2_uk_n1824, u2_uk_n1825, u2_uk_n1826, u2_uk_n1835, u2_uk_n1836, u2_uk_n1837, u2_uk_n1840, u2_uk_n1845, u2_uk_n1846, 
       u2_uk_n1849, u2_uk_n1853, u2_uk_n1854, u2_uk_n1855, u2_uk_n1856, u2_uk_n187, u2_uk_n191, u2_uk_n202, u2_uk_n207, 
       u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n230, u2_uk_n231, u2_uk_n31, u2_uk_n385, 
       u2_uk_n702, u2_uk_n92, u2_uk_n93, u2_uk_n933, u2_uk_n939, u2_uk_n941, u2_uk_n942, u2_uk_n943, u2_uk_n944, 
       u2_uk_n945, u0_FP_13, u0_FP_17, u0_FP_18, u0_FP_2, u0_FP_23, u0_FP_28, u0_FP_31, u0_FP_9, u0_N100, 
        u0_N102, u0_N107, u0_N110, u0_N116, u0_N117, u0_N122, u0_N127, u0_N161, u0_N165, 
        u0_N168, u0_N172, u0_N175, u0_N176, u0_N177, u0_N182, u0_N183, u0_N187, u0_N189, 
        u0_N190, u0_N225, u0_N232, u0_N236, u0_N240, u0_N241, u0_N246, u0_N251, u0_N254, 
        u0_uk_n680, u1_N192, u1_N201, u1_N211, u1_N217, u1_N36, u1_N46, u1_N52, u1_N58, 
        u2_N101, u2_N105, u2_N111, u2_N115, u2_N119, u2_N121, u2_N125, u2_N225, u2_N236, 
        u2_N241, u2_N251, u2_N257, u2_N261, u2_N264, u2_N268, u2_N271, u2_N272, u2_N273, 
        u2_N278, u2_N279, u2_N283, u2_N285, u2_N286, u2_N324, u2_N334, u2_N340, u2_N346, 
        u2_N417, u2_N419, u2_N421, u2_N422, u2_N424, u2_N426, u2_N427, u2_N428, u2_N431, 
        u2_N432, u2_N433, u2_N434, u2_N437, u2_N438, u2_N439, u2_N443, u2_N444, u2_N445, 
        u2_N446, u2_N447, u2_N450, u2_N451, u2_N452, u2_N454, u2_N455, u2_N458, u2_N459, 
        u2_N461, u2_N462, u2_N466, u2_N468, u2_N469, u2_N472, u2_N474, u2_N476, u2_N479, 
        u2_N65, u2_N76, u2_N81, u2_N91, u2_N96, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n1034, 
        u2_uk_n109, u2_uk_n1143, u2_uk_n117, u2_uk_n128, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n161, 
        u2_uk_n162, u2_uk_n17, u2_uk_n203, u2_uk_n222, u2_uk_n223, u2_uk_n605, u2_uk_n63, u2_uk_n83, u2_uk_n94, 
        u2_uk_n988, u2_uk_n99 );
  input u0_FP_33, u0_FP_34, u0_FP_35, u0_FP_36, u0_FP_37, u0_FP_38, u0_FP_39, u0_FP_40, u0_FP_41, 
        u0_FP_64, u0_K16_4, u0_K16_8, u0_K4_43, u0_K4_48, u0_K6_11, u0_K6_13, u0_K6_16, u0_K8_1, 
        u0_K8_11, u0_L14_13, u0_L14_17, u0_L14_18, u0_L14_2, u0_L14_23, u0_L14_28, u0_L14_31, u0_L14_9, 
        u0_L2_12, u0_L2_15, u0_L2_21, u0_L2_22, u0_L2_27, u0_L2_32, u0_L2_5, u0_L2_7, u0_L4_13, 
        u0_L4_16, u0_L4_17, u0_L4_18, u0_L4_2, u0_L4_23, u0_L4_24, u0_L4_28, u0_L4_30, u0_L4_31, 
        u0_L4_6, u0_L4_9, u0_L6_13, u0_L6_17, u0_L6_18, u0_L6_2, u0_L6_23, u0_L6_28, u0_L6_31, 
        u0_L6_9, u0_R2_1, u0_R2_24, u0_R2_25, u0_R2_26, u0_R2_27, u0_R2_28, u0_R2_29, u0_R2_30, 
        u0_R2_31, u0_R2_32, u0_R4_1, u0_R4_10, u0_R4_11, u0_R4_12, u0_R4_13, u0_R4_2, u0_R4_3, 
        u0_R4_32, u0_R4_4, u0_R4_5, u0_R4_6, u0_R4_7, u0_R4_8, u0_R4_9, u0_R6_1, u0_R6_2, 
        u0_R6_3, u0_R6_32, u0_R6_4, u0_R6_5, u0_R6_6, u0_R6_7, u0_R6_8, u0_R6_9, u0_key_r_44, 
        u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_39, u0_uk_K_r2_50, u0_uk_K_r4_3, u0_uk_K_r4_33, u0_uk_K_r4_4, u0_uk_K_r4_41, u0_uk_K_r4_47, 
        u0_uk_K_r4_54, u0_uk_K_r4_55, u0_uk_K_r6_10, u0_uk_K_r6_19, u0_uk_K_r6_27, u0_uk_K_r6_3, u0_uk_K_r6_53, u0_uk_n10, u0_uk_n100, 
        u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n141, u0_uk_n142, u0_uk_n145, 
        u0_uk_n146, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, 
        u0_uk_n202, u0_uk_n207, u0_uk_n223, u0_uk_n240, u0_uk_n242, u0_uk_n251, u0_uk_n252, u0_uk_n257, u0_uk_n27, 
        u0_uk_n31, u0_uk_n318, u0_uk_n324, u0_uk_n330, u0_uk_n337, u0_uk_n339, u0_uk_n343, u0_uk_n344, u0_uk_n350, 
        u0_uk_n351, u0_uk_n352, u0_uk_n356, u0_uk_n358, u0_uk_n410, u0_uk_n414, u0_uk_n423, u0_uk_n426, u0_uk_n427, 
        u0_uk_n432, u0_uk_n435, u0_uk_n436, u0_uk_n441, u0_uk_n442, u0_uk_n448, u0_uk_n498, u0_uk_n499, u0_uk_n505, 
        u0_uk_n506, u0_uk_n508, u0_uk_n513, u0_uk_n514, u0_uk_n516, u0_uk_n521, u0_uk_n522, u0_uk_n527, u0_uk_n528, 
        u0_uk_n537, u0_uk_n538, u0_uk_n539, u0_uk_n60, u0_uk_n63, u0_uk_n630, u0_uk_n636, u0_uk_n637, u0_uk_n639, 
        u0_uk_n640, u0_uk_n644, u0_uk_n646, u0_uk_n651, u0_uk_n652, u0_uk_n659, u0_uk_n660, u0_uk_n664, u0_uk_n667, 
        u0_uk_n668, u0_uk_n785, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n83, u0_uk_n92, u0_uk_n93, u1_L0_15, 
        u1_L0_21, u1_L0_27, u1_L0_5, u1_L5_1, u1_L5_10, u1_L5_20, u1_L5_26, u1_R0_1, u1_R0_28, 
        u1_R0_29, u1_R0_30, u1_R0_31, u1_R0_32, u1_R5_12, u1_R5_13, u1_R5_14, u1_R5_15, u1_R5_16, 
        u1_R5_17, u1_uk_K_r0_2, u1_uk_K_r0_52, u1_uk_K_r5_13, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_40, u1_uk_K_r5_5, u1_uk_K_r5_53, 
        u1_uk_n10, u1_uk_n11, u1_uk_n1266, u1_uk_n1271, u1_uk_n1276, u1_uk_n1281, u1_uk_n1282, u1_uk_n1286, u1_uk_n1293, 
        u1_uk_n1303, u1_uk_n1304, u1_uk_n145, u1_uk_n1483, u1_uk_n1495, u1_uk_n1498, u1_uk_n1505, u1_uk_n1526, u1_uk_n155, 
        u1_uk_n162, u1_uk_n17, u1_uk_n187, u1_uk_n191, u1_uk_n207, u1_uk_n217, u1_uk_n222, u1_uk_n231, u1_uk_n240, 
        u1_uk_n271, u1_uk_n297, u1_uk_n298, u1_uk_n60, u1_uk_n92, u2_K11_45, u2_K11_48, u2_K14_10, u2_K14_11, 
        u2_K14_12, u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_3, u2_K14_39, u2_K14_42, 
        u2_K14_6, u2_K14_8, u2_K15_28, u2_K15_29, u2_K15_31, u2_K15_34, u2_K15_35, u2_K15_39, u2_K3_7, 
        u2_K4_14, u2_K4_21, u2_K4_22, u2_K8_8, u2_K9_15, u2_K9_3, u2_K9_5, u2_L12_11, u2_L12_12, 
        u2_L12_13, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_19, u2_L12_2, u2_L12_22, u2_L12_23, u2_L12_24, 
        u2_L12_28, u2_L12_29, u2_L12_30, u2_L12_31, u2_L12_32, u2_L12_4, u2_L12_6, u2_L12_7, u2_L12_9, 
        u2_L13_11, u2_L13_12, u2_L13_14, u2_L13_15, u2_L13_19, u2_L13_21, u2_L13_22, u2_L13_25, u2_L13_27, 
        u2_L13_29, u2_L13_3, u2_L13_32, u2_L13_4, u2_L13_5, u2_L13_7, u2_L13_8, u2_L1_13, u2_L1_18, 
        u2_L1_2, u2_L1_28, u2_L2_1, u2_L2_10, u2_L2_16, u2_L2_20, u2_L2_24, u2_L2_26, u2_L2_30, 
        u2_L2_6, u2_L6_13, u2_L6_18, u2_L6_2, u2_L6_28, u2_L7_13, u2_L7_16, u2_L7_17, u2_L7_18, 
        u2_L7_2, u2_L7_23, u2_L7_24, u2_L7_28, u2_L7_30, u2_L7_31, u2_L7_6, u2_L7_9, u2_L9_15, 
        u2_L9_21, u2_L9_27, u2_L9_5, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_2, 
        u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_23, u2_R12_24, u2_R12_25, u2_R12_26, u2_R12_27, u2_R12_28, 
        u2_R12_29, u2_R12_3, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, 
        u2_R13_1, u2_R13_16, u2_R13_17, u2_R13_18, u2_R13_19, u2_R13_20, u2_R13_21, u2_R13_22, u2_R13_23, 
        u2_R13_24, u2_R13_25, u2_R13_26, u2_R13_27, u2_R13_28, u2_R13_29, u2_R13_30, u2_R13_31, u2_R13_32, 
        u2_R1_4, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_10, u2_R2_11, u2_R2_12, 
        u2_R2_13, u2_R2_14, u2_R2_15, u2_R2_16, u2_R2_17, u2_R2_8, u2_R2_9, u2_R6_4, u2_R6_5, 
        u2_R6_6, u2_R6_7, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_10, u2_R7_11, u2_R7_12, u2_R7_13, 
        u2_R7_2, u2_R7_3, u2_R7_32, u2_R7_4, u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, 
        u2_R9_1, u2_R9_28, u2_R9_29, u2_R9_30, u2_R9_31, u2_R9_32, u2_key_r_1, u2_key_r_49, u2_uk_K_r11_33, 
        u2_uk_K_r12_1, u2_uk_K_r12_10, u2_uk_K_r12_30, u2_uk_K_r12_36, u2_uk_K_r12_7, u2_uk_K_r13_0, u2_uk_K_r13_22, u2_uk_K_r13_38, u2_uk_K_r1_18, 
        u2_uk_K_r2_18, u2_uk_K_r2_27, u2_uk_K_r2_50, u2_uk_K_r2_55, u2_uk_K_r6_3, u2_uk_K_r6_53, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_32, 
        u2_uk_K_r7_39, u2_uk_K_r7_46, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r9_15, u2_uk_K_r9_23, u2_uk_n1022, u2_uk_n1024, u2_uk_n1097, 
        u2_uk_n11, u2_uk_n110, u2_uk_n1119, u2_uk_n1120, u2_uk_n1121, u2_uk_n1125, u2_uk_n1130, u2_uk_n1141, u2_uk_n118, 
        u2_uk_n1280, u2_uk_n1285, u2_uk_n1286, u2_uk_n129, u2_uk_n1291, u2_uk_n1295, u2_uk_n1296, u2_uk_n1306, u2_uk_n1311, 
        u2_uk_n1322, u2_uk_n1324, u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1335, u2_uk_n1339, u2_uk_n1347, u2_uk_n1348, 
        u2_uk_n1356, u2_uk_n1363, u2_uk_n147, u2_uk_n1500, u2_uk_n1502, u2_uk_n1506, u2_uk_n1508, u2_uk_n1519, u2_uk_n1521, 
        u2_uk_n1535, u2_uk_n1543, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n155, u2_uk_n1555, u2_uk_n1556, u2_uk_n1563, 
        u2_uk_n1568, u2_uk_n1573, u2_uk_n1574, u2_uk_n1580, u2_uk_n163, u2_uk_n1632, u2_uk_n164, u2_uk_n1653, u2_uk_n1673, 
        u2_uk_n1674, u2_uk_n1769, u2_uk_n1770, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1781, u2_uk_n1783, 
        u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1791, u2_uk_n1793, u2_uk_n1794, u2_uk_n1796, u2_uk_n1797, u2_uk_n1801, 
        u2_uk_n1803, u2_uk_n1805, u2_uk_n1807, u2_uk_n1808, u2_uk_n1811, u2_uk_n1817, u2_uk_n1818, u2_uk_n1819, u2_uk_n182, 
        u2_uk_n1824, u2_uk_n1825, u2_uk_n1826, u2_uk_n1835, u2_uk_n1836, u2_uk_n1837, u2_uk_n1840, u2_uk_n1845, u2_uk_n1846, 
        u2_uk_n1849, u2_uk_n1853, u2_uk_n1854, u2_uk_n1855, u2_uk_n1856, u2_uk_n187, u2_uk_n191, u2_uk_n202, u2_uk_n207, 
        u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n230, u2_uk_n231, u2_uk_n31, u2_uk_n385, 
        u2_uk_n702, u2_uk_n92, u2_uk_n93, u2_uk_n933, u2_uk_n939, u2_uk_n941, u2_uk_n942, u2_uk_n943, u2_uk_n944, 
        u2_uk_n945;
  output u0_FP_13, u0_FP_17, u0_FP_18, u0_FP_2, u0_FP_23, u0_FP_28, u0_FP_31, u0_FP_9, u0_N100, 
        u0_N102, u0_N107, u0_N110, u0_N116, u0_N117, u0_N122, u0_N127, u0_N161, u0_N165, 
        u0_N168, u0_N172, u0_N175, u0_N176, u0_N177, u0_N182, u0_N183, u0_N187, u0_N189, 
        u0_N190, u0_N225, u0_N232, u0_N236, u0_N240, u0_N241, u0_N246, u0_N251, u0_N254, 
        u0_uk_n680, u1_N192, u1_N201, u1_N211, u1_N217, u1_N36, u1_N46, u1_N52, u1_N58, 
        u2_N101, u2_N105, u2_N111, u2_N115, u2_N119, u2_N121, u2_N125, u2_N225, u2_N236, 
        u2_N241, u2_N251, u2_N257, u2_N261, u2_N264, u2_N268, u2_N271, u2_N272, u2_N273, 
        u2_N278, u2_N279, u2_N283, u2_N285, u2_N286, u2_N324, u2_N334, u2_N340, u2_N346, 
        u2_N417, u2_N419, u2_N421, u2_N422, u2_N424, u2_N426, u2_N427, u2_N428, u2_N431, 
        u2_N432, u2_N433, u2_N434, u2_N437, u2_N438, u2_N439, u2_N443, u2_N444, u2_N445, 
        u2_N446, u2_N447, u2_N450, u2_N451, u2_N452, u2_N454, u2_N455, u2_N458, u2_N459, 
        u2_N461, u2_N462, u2_N466, u2_N468, u2_N469, u2_N472, u2_N474, u2_N476, u2_N479, 
        u2_N65, u2_N76, u2_N81, u2_N91, u2_N96, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n1034, 
        u2_uk_n109, u2_uk_n1143, u2_uk_n117, u2_uk_n128, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n161, 
        u2_uk_n162, u2_uk_n17, u2_uk_n203, u2_uk_n222, u2_uk_n223, u2_uk_n605, u2_uk_n63, u2_uk_n83, u2_uk_n94, 
        u2_uk_n988, u2_uk_n99;
  wire u0_K16_1, u0_K16_10, u0_K16_11, u0_K16_12, u0_K16_2, u0_K16_3, u0_K16_5, u0_K16_6, u0_K16_7, 
       u0_K16_9, u0_K4_37, u0_K4_38, u0_K4_39, u0_K4_40, u0_K4_41, u0_K4_42, u0_K4_44, u0_K4_45, 
       u0_K4_46, u0_K4_47, u0_K6_1, u0_K6_10, u0_K6_12, u0_K6_14, u0_K6_15, u0_K6_17, u0_K6_18, 
       u0_K6_2, u0_K6_3, u0_K6_4, u0_K6_5, u0_K6_6, u0_K6_7, u0_K6_8, u0_K6_9, u0_K8_10, 
       u0_K8_12, u0_K8_2, u0_K8_3, u0_K8_4, u0_K8_5, u0_K8_6, u0_K8_7, u0_K8_8, u0_K8_9, 
       u0_out15_13, u0_out15_17, u0_out15_18, u0_out15_2, u0_out15_23, u0_out15_28, u0_out15_31, u0_out15_9, u0_out3_12, 
       u0_out3_15, u0_out3_21, u0_out3_22, u0_out3_27, u0_out3_32, u0_out3_5, u0_out3_7, u0_out5_13, u0_out5_16, 
       u0_out5_17, u0_out5_18, u0_out5_2, u0_out5_23, u0_out5_24, u0_out5_28, u0_out5_30, u0_out5_31, u0_out5_6, 
       u0_out5_9, u0_out7_13, u0_out7_17, u0_out7_18, u0_out7_2, u0_out7_23, u0_out7_28, u0_out7_31, u0_out7_9, 
       u0_u15_X_1, u0_u15_X_10, u0_u15_X_11, u0_u15_X_12, u0_u15_X_2, u0_u15_X_3, u0_u15_X_4, u0_u15_X_5, u0_u15_X_6, 
       u0_u15_X_7, u0_u15_X_8, u0_u15_X_9, u0_u15_u0_n100, u0_u15_u0_n101, u0_u15_u0_n102, u0_u15_u0_n103, u0_u15_u0_n104, u0_u15_u0_n105, 
       u0_u15_u0_n106, u0_u15_u0_n107, u0_u15_u0_n108, u0_u15_u0_n109, u0_u15_u0_n110, u0_u15_u0_n111, u0_u15_u0_n112, u0_u15_u0_n113, u0_u15_u0_n114, 
       u0_u15_u0_n115, u0_u15_u0_n116, u0_u15_u0_n117, u0_u15_u0_n118, u0_u15_u0_n119, u0_u15_u0_n120, u0_u15_u0_n121, u0_u15_u0_n122, u0_u15_u0_n123, 
       u0_u15_u0_n124, u0_u15_u0_n125, u0_u15_u0_n126, u0_u15_u0_n127, u0_u15_u0_n128, u0_u15_u0_n129, u0_u15_u0_n130, u0_u15_u0_n131, u0_u15_u0_n132, 
       u0_u15_u0_n133, u0_u15_u0_n134, u0_u15_u0_n135, u0_u15_u0_n136, u0_u15_u0_n137, u0_u15_u0_n138, u0_u15_u0_n139, u0_u15_u0_n140, u0_u15_u0_n141, 
       u0_u15_u0_n142, u0_u15_u0_n143, u0_u15_u0_n144, u0_u15_u0_n145, u0_u15_u0_n146, u0_u15_u0_n147, u0_u15_u0_n148, u0_u15_u0_n149, u0_u15_u0_n150, 
       u0_u15_u0_n151, u0_u15_u0_n152, u0_u15_u0_n153, u0_u15_u0_n154, u0_u15_u0_n155, u0_u15_u0_n156, u0_u15_u0_n157, u0_u15_u0_n158, u0_u15_u0_n159, 
       u0_u15_u0_n160, u0_u15_u0_n161, u0_u15_u0_n162, u0_u15_u0_n163, u0_u15_u0_n164, u0_u15_u0_n165, u0_u15_u0_n166, u0_u15_u0_n167, u0_u15_u0_n168, 
       u0_u15_u0_n169, u0_u15_u0_n170, u0_u15_u0_n171, u0_u15_u0_n172, u0_u15_u0_n173, u0_u15_u0_n174, u0_u15_u0_n88, u0_u15_u0_n89, u0_u15_u0_n90, 
       u0_u15_u0_n91, u0_u15_u0_n92, u0_u15_u0_n93, u0_u15_u0_n94, u0_u15_u0_n95, u0_u15_u0_n96, u0_u15_u0_n97, u0_u15_u0_n98, u0_u15_u0_n99, 
       u0_u15_u1_n100, u0_u15_u1_n101, u0_u15_u1_n102, u0_u15_u1_n103, u0_u15_u1_n104, u0_u15_u1_n105, u0_u15_u1_n106, u0_u15_u1_n107, u0_u15_u1_n108, 
       u0_u15_u1_n109, u0_u15_u1_n110, u0_u15_u1_n111, u0_u15_u1_n112, u0_u15_u1_n113, u0_u15_u1_n114, u0_u15_u1_n115, u0_u15_u1_n116, u0_u15_u1_n117, 
       u0_u15_u1_n118, u0_u15_u1_n119, u0_u15_u1_n120, u0_u15_u1_n121, u0_u15_u1_n122, u0_u15_u1_n123, u0_u15_u1_n124, u0_u15_u1_n125, u0_u15_u1_n126, 
       u0_u15_u1_n127, u0_u15_u1_n128, u0_u15_u1_n129, u0_u15_u1_n130, u0_u15_u1_n131, u0_u15_u1_n132, u0_u15_u1_n133, u0_u15_u1_n134, u0_u15_u1_n135, 
       u0_u15_u1_n136, u0_u15_u1_n137, u0_u15_u1_n138, u0_u15_u1_n139, u0_u15_u1_n140, u0_u15_u1_n141, u0_u15_u1_n142, u0_u15_u1_n143, u0_u15_u1_n144, 
       u0_u15_u1_n145, u0_u15_u1_n146, u0_u15_u1_n147, u0_u15_u1_n148, u0_u15_u1_n149, u0_u15_u1_n150, u0_u15_u1_n151, u0_u15_u1_n152, u0_u15_u1_n153, 
       u0_u15_u1_n154, u0_u15_u1_n155, u0_u15_u1_n156, u0_u15_u1_n157, u0_u15_u1_n158, u0_u15_u1_n159, u0_u15_u1_n160, u0_u15_u1_n161, u0_u15_u1_n162, 
       u0_u15_u1_n163, u0_u15_u1_n164, u0_u15_u1_n165, u0_u15_u1_n166, u0_u15_u1_n167, u0_u15_u1_n168, u0_u15_u1_n169, u0_u15_u1_n170, u0_u15_u1_n171, 
       u0_u15_u1_n172, u0_u15_u1_n173, u0_u15_u1_n174, u0_u15_u1_n175, u0_u15_u1_n176, u0_u15_u1_n177, u0_u15_u1_n178, u0_u15_u1_n179, u0_u15_u1_n180, 
       u0_u15_u1_n181, u0_u15_u1_n182, u0_u15_u1_n183, u0_u15_u1_n184, u0_u15_u1_n185, u0_u15_u1_n186, u0_u15_u1_n187, u0_u15_u1_n188, u0_u15_u1_n95, 
       u0_u15_u1_n96, u0_u15_u1_n97, u0_u15_u1_n98, u0_u15_u1_n99, u0_u3_X_37, u0_u3_X_38, u0_u3_X_39, u0_u3_X_40, u0_u3_X_41, 
       u0_u3_X_42, u0_u3_X_43, u0_u3_X_44, u0_u3_X_45, u0_u3_X_46, u0_u3_X_47, u0_u3_X_48, u0_u3_u6_n100, u0_u3_u6_n101, 
       u0_u3_u6_n102, u0_u3_u6_n103, u0_u3_u6_n104, u0_u3_u6_n105, u0_u3_u6_n106, u0_u3_u6_n107, u0_u3_u6_n108, u0_u3_u6_n109, u0_u3_u6_n110, 
       u0_u3_u6_n111, u0_u3_u6_n112, u0_u3_u6_n113, u0_u3_u6_n114, u0_u3_u6_n115, u0_u3_u6_n116, u0_u3_u6_n117, u0_u3_u6_n118, u0_u3_u6_n119, 
       u0_u3_u6_n120, u0_u3_u6_n121, u0_u3_u6_n122, u0_u3_u6_n123, u0_u3_u6_n124, u0_u3_u6_n125, u0_u3_u6_n126, u0_u3_u6_n127, u0_u3_u6_n128, 
       u0_u3_u6_n129, u0_u3_u6_n130, u0_u3_u6_n131, u0_u3_u6_n132, u0_u3_u6_n133, u0_u3_u6_n134, u0_u3_u6_n135, u0_u3_u6_n136, u0_u3_u6_n137, 
       u0_u3_u6_n138, u0_u3_u6_n139, u0_u3_u6_n140, u0_u3_u6_n141, u0_u3_u6_n142, u0_u3_u6_n143, u0_u3_u6_n144, u0_u3_u6_n145, u0_u3_u6_n146, 
       u0_u3_u6_n147, u0_u3_u6_n148, u0_u3_u6_n149, u0_u3_u6_n150, u0_u3_u6_n151, u0_u3_u6_n152, u0_u3_u6_n153, u0_u3_u6_n154, u0_u3_u6_n155, 
       u0_u3_u6_n156, u0_u3_u6_n157, u0_u3_u6_n158, u0_u3_u6_n159, u0_u3_u6_n160, u0_u3_u6_n161, u0_u3_u6_n162, u0_u3_u6_n163, u0_u3_u6_n164, 
       u0_u3_u6_n165, u0_u3_u6_n166, u0_u3_u6_n167, u0_u3_u6_n168, u0_u3_u6_n169, u0_u3_u6_n170, u0_u3_u6_n171, u0_u3_u6_n172, u0_u3_u6_n173, 
       u0_u3_u6_n174, u0_u3_u6_n88, u0_u3_u6_n89, u0_u3_u6_n90, u0_u3_u6_n91, u0_u3_u6_n92, u0_u3_u6_n93, u0_u3_u6_n94, u0_u3_u6_n95, 
       u0_u3_u6_n96, u0_u3_u6_n97, u0_u3_u6_n98, u0_u3_u6_n99, u0_u3_u7_n100, u0_u3_u7_n101, u0_u3_u7_n102, u0_u3_u7_n103, u0_u3_u7_n104, 
       u0_u3_u7_n105, u0_u3_u7_n106, u0_u3_u7_n107, u0_u3_u7_n108, u0_u3_u7_n109, u0_u3_u7_n110, u0_u3_u7_n111, u0_u3_u7_n112, u0_u3_u7_n113, 
       u0_u3_u7_n114, u0_u3_u7_n115, u0_u3_u7_n116, u0_u3_u7_n117, u0_u3_u7_n118, u0_u3_u7_n119, u0_u3_u7_n120, u0_u3_u7_n121, u0_u3_u7_n122, 
       u0_u3_u7_n123, u0_u3_u7_n124, u0_u3_u7_n125, u0_u3_u7_n126, u0_u3_u7_n127, u0_u3_u7_n128, u0_u3_u7_n129, u0_u3_u7_n130, u0_u3_u7_n131, 
       u0_u3_u7_n132, u0_u3_u7_n133, u0_u3_u7_n134, u0_u3_u7_n135, u0_u3_u7_n136, u0_u3_u7_n137, u0_u3_u7_n138, u0_u3_u7_n139, u0_u3_u7_n140, 
       u0_u3_u7_n141, u0_u3_u7_n142, u0_u3_u7_n143, u0_u3_u7_n144, u0_u3_u7_n145, u0_u3_u7_n146, u0_u3_u7_n147, u0_u3_u7_n148, u0_u3_u7_n149, 
       u0_u3_u7_n150, u0_u3_u7_n151, u0_u3_u7_n152, u0_u3_u7_n153, u0_u3_u7_n154, u0_u3_u7_n155, u0_u3_u7_n156, u0_u3_u7_n157, u0_u3_u7_n158, 
       u0_u3_u7_n159, u0_u3_u7_n160, u0_u3_u7_n161, u0_u3_u7_n162, u0_u3_u7_n163, u0_u3_u7_n164, u0_u3_u7_n165, u0_u3_u7_n166, u0_u3_u7_n167, 
       u0_u3_u7_n168, u0_u3_u7_n169, u0_u3_u7_n170, u0_u3_u7_n171, u0_u3_u7_n172, u0_u3_u7_n173, u0_u3_u7_n174, u0_u3_u7_n175, u0_u3_u7_n176, 
       u0_u3_u7_n177, u0_u3_u7_n178, u0_u3_u7_n179, u0_u3_u7_n180, u0_u3_u7_n91, u0_u3_u7_n92, u0_u3_u7_n93, u0_u3_u7_n94, u0_u3_u7_n95, 
       u0_u3_u7_n96, u0_u3_u7_n97, u0_u3_u7_n98, u0_u3_u7_n99, u0_u5_X_1, u0_u5_X_10, u0_u5_X_11, u0_u5_X_12, u0_u5_X_13, 
       u0_u5_X_14, u0_u5_X_15, u0_u5_X_16, u0_u5_X_17, u0_u5_X_18, u0_u5_X_2, u0_u5_X_3, u0_u5_X_4, u0_u5_X_5, 
       u0_u5_X_6, u0_u5_X_7, u0_u5_X_8, u0_u5_X_9, u0_u5_u0_n100, u0_u5_u0_n101, u0_u5_u0_n102, u0_u5_u0_n103, u0_u5_u0_n104, 
       u0_u5_u0_n105, u0_u5_u0_n106, u0_u5_u0_n107, u0_u5_u0_n108, u0_u5_u0_n109, u0_u5_u0_n110, u0_u5_u0_n111, u0_u5_u0_n112, u0_u5_u0_n113, 
       u0_u5_u0_n114, u0_u5_u0_n115, u0_u5_u0_n116, u0_u5_u0_n117, u0_u5_u0_n118, u0_u5_u0_n119, u0_u5_u0_n120, u0_u5_u0_n121, u0_u5_u0_n122, 
       u0_u5_u0_n123, u0_u5_u0_n124, u0_u5_u0_n125, u0_u5_u0_n126, u0_u5_u0_n127, u0_u5_u0_n128, u0_u5_u0_n129, u0_u5_u0_n130, u0_u5_u0_n131, 
       u0_u5_u0_n132, u0_u5_u0_n133, u0_u5_u0_n134, u0_u5_u0_n135, u0_u5_u0_n136, u0_u5_u0_n137, u0_u5_u0_n138, u0_u5_u0_n139, u0_u5_u0_n140, 
       u0_u5_u0_n141, u0_u5_u0_n142, u0_u5_u0_n143, u0_u5_u0_n144, u0_u5_u0_n145, u0_u5_u0_n146, u0_u5_u0_n147, u0_u5_u0_n148, u0_u5_u0_n149, 
       u0_u5_u0_n150, u0_u5_u0_n151, u0_u5_u0_n152, u0_u5_u0_n153, u0_u5_u0_n154, u0_u5_u0_n155, u0_u5_u0_n156, u0_u5_u0_n157, u0_u5_u0_n158, 
       u0_u5_u0_n159, u0_u5_u0_n160, u0_u5_u0_n161, u0_u5_u0_n162, u0_u5_u0_n163, u0_u5_u0_n164, u0_u5_u0_n165, u0_u5_u0_n166, u0_u5_u0_n167, 
       u0_u5_u0_n168, u0_u5_u0_n169, u0_u5_u0_n170, u0_u5_u0_n171, u0_u5_u0_n172, u0_u5_u0_n173, u0_u5_u0_n174, u0_u5_u0_n88, u0_u5_u0_n89, 
       u0_u5_u0_n90, u0_u5_u0_n91, u0_u5_u0_n92, u0_u5_u0_n93, u0_u5_u0_n94, u0_u5_u0_n95, u0_u5_u0_n96, u0_u5_u0_n97, u0_u5_u0_n98, 
       u0_u5_u0_n99, u0_u5_u1_n100, u0_u5_u1_n101, u0_u5_u1_n102, u0_u5_u1_n103, u0_u5_u1_n104, u0_u5_u1_n105, u0_u5_u1_n106, u0_u5_u1_n107, 
       u0_u5_u1_n108, u0_u5_u1_n109, u0_u5_u1_n110, u0_u5_u1_n111, u0_u5_u1_n112, u0_u5_u1_n113, u0_u5_u1_n114, u0_u5_u1_n115, u0_u5_u1_n116, 
       u0_u5_u1_n117, u0_u5_u1_n118, u0_u5_u1_n119, u0_u5_u1_n120, u0_u5_u1_n121, u0_u5_u1_n122, u0_u5_u1_n123, u0_u5_u1_n124, u0_u5_u1_n125, 
       u0_u5_u1_n126, u0_u5_u1_n127, u0_u5_u1_n128, u0_u5_u1_n129, u0_u5_u1_n130, u0_u5_u1_n131, u0_u5_u1_n132, u0_u5_u1_n133, u0_u5_u1_n134, 
       u0_u5_u1_n135, u0_u5_u1_n136, u0_u5_u1_n137, u0_u5_u1_n138, u0_u5_u1_n139, u0_u5_u1_n140, u0_u5_u1_n141, u0_u5_u1_n142, u0_u5_u1_n143, 
       u0_u5_u1_n144, u0_u5_u1_n145, u0_u5_u1_n146, u0_u5_u1_n147, u0_u5_u1_n148, u0_u5_u1_n149, u0_u5_u1_n150, u0_u5_u1_n151, u0_u5_u1_n152, 
       u0_u5_u1_n153, u0_u5_u1_n154, u0_u5_u1_n155, u0_u5_u1_n156, u0_u5_u1_n157, u0_u5_u1_n158, u0_u5_u1_n159, u0_u5_u1_n160, u0_u5_u1_n161, 
       u0_u5_u1_n162, u0_u5_u1_n163, u0_u5_u1_n164, u0_u5_u1_n165, u0_u5_u1_n166, u0_u5_u1_n167, u0_u5_u1_n168, u0_u5_u1_n169, u0_u5_u1_n170, 
       u0_u5_u1_n171, u0_u5_u1_n172, u0_u5_u1_n173, u0_u5_u1_n174, u0_u5_u1_n175, u0_u5_u1_n176, u0_u5_u1_n177, u0_u5_u1_n178, u0_u5_u1_n179, 
       u0_u5_u1_n180, u0_u5_u1_n181, u0_u5_u1_n182, u0_u5_u1_n183, u0_u5_u1_n184, u0_u5_u1_n185, u0_u5_u1_n186, u0_u5_u1_n187, u0_u5_u1_n188, 
       u0_u5_u1_n95, u0_u5_u1_n96, u0_u5_u1_n97, u0_u5_u1_n98, u0_u5_u1_n99, u0_u5_u2_n100, u0_u5_u2_n101, u0_u5_u2_n102, u0_u5_u2_n103, 
       u0_u5_u2_n104, u0_u5_u2_n105, u0_u5_u2_n106, u0_u5_u2_n107, u0_u5_u2_n108, u0_u5_u2_n109, u0_u5_u2_n110, u0_u5_u2_n111, u0_u5_u2_n112, 
       u0_u5_u2_n113, u0_u5_u2_n114, u0_u5_u2_n115, u0_u5_u2_n116, u0_u5_u2_n117, u0_u5_u2_n118, u0_u5_u2_n119, u0_u5_u2_n120, u0_u5_u2_n121, 
       u0_u5_u2_n122, u0_u5_u2_n123, u0_u5_u2_n124, u0_u5_u2_n125, u0_u5_u2_n126, u0_u5_u2_n127, u0_u5_u2_n128, u0_u5_u2_n129, u0_u5_u2_n130, 
       u0_u5_u2_n131, u0_u5_u2_n132, u0_u5_u2_n133, u0_u5_u2_n134, u0_u5_u2_n135, u0_u5_u2_n136, u0_u5_u2_n137, u0_u5_u2_n138, u0_u5_u2_n139, 
       u0_u5_u2_n140, u0_u5_u2_n141, u0_u5_u2_n142, u0_u5_u2_n143, u0_u5_u2_n144, u0_u5_u2_n145, u0_u5_u2_n146, u0_u5_u2_n147, u0_u5_u2_n148, 
       u0_u5_u2_n149, u0_u5_u2_n150, u0_u5_u2_n151, u0_u5_u2_n152, u0_u5_u2_n153, u0_u5_u2_n154, u0_u5_u2_n155, u0_u5_u2_n156, u0_u5_u2_n157, 
       u0_u5_u2_n158, u0_u5_u2_n159, u0_u5_u2_n160, u0_u5_u2_n161, u0_u5_u2_n162, u0_u5_u2_n163, u0_u5_u2_n164, u0_u5_u2_n165, u0_u5_u2_n166, 
       u0_u5_u2_n167, u0_u5_u2_n168, u0_u5_u2_n169, u0_u5_u2_n170, u0_u5_u2_n171, u0_u5_u2_n172, u0_u5_u2_n173, u0_u5_u2_n174, u0_u5_u2_n175, 
       u0_u5_u2_n176, u0_u5_u2_n177, u0_u5_u2_n178, u0_u5_u2_n179, u0_u5_u2_n180, u0_u5_u2_n181, u0_u5_u2_n182, u0_u5_u2_n183, u0_u5_u2_n184, 
       u0_u5_u2_n185, u0_u5_u2_n186, u0_u5_u2_n187, u0_u5_u2_n188, u0_u5_u2_n95, u0_u5_u2_n96, u0_u5_u2_n97, u0_u5_u2_n98, u0_u5_u2_n99, 
       u0_u7_X_1, u0_u7_X_10, u0_u7_X_11, u0_u7_X_12, u0_u7_X_2, u0_u7_X_3, u0_u7_X_4, u0_u7_X_5, u0_u7_X_6, 
       u0_u7_X_7, u0_u7_X_8, u0_u7_X_9, u0_u7_u0_n100, u0_u7_u0_n101, u0_u7_u0_n102, u0_u7_u0_n103, u0_u7_u0_n104, u0_u7_u0_n105, 
       u0_u7_u0_n106, u0_u7_u0_n107, u0_u7_u0_n108, u0_u7_u0_n109, u0_u7_u0_n110, u0_u7_u0_n111, u0_u7_u0_n112, u0_u7_u0_n113, u0_u7_u0_n114, 
       u0_u7_u0_n115, u0_u7_u0_n116, u0_u7_u0_n117, u0_u7_u0_n118, u0_u7_u0_n119, u0_u7_u0_n120, u0_u7_u0_n121, u0_u7_u0_n122, u0_u7_u0_n123, 
       u0_u7_u0_n124, u0_u7_u0_n125, u0_u7_u0_n126, u0_u7_u0_n127, u0_u7_u0_n128, u0_u7_u0_n129, u0_u7_u0_n130, u0_u7_u0_n131, u0_u7_u0_n132, 
       u0_u7_u0_n133, u0_u7_u0_n134, u0_u7_u0_n135, u0_u7_u0_n136, u0_u7_u0_n137, u0_u7_u0_n138, u0_u7_u0_n139, u0_u7_u0_n140, u0_u7_u0_n141, 
       u0_u7_u0_n142, u0_u7_u0_n143, u0_u7_u0_n144, u0_u7_u0_n145, u0_u7_u0_n146, u0_u7_u0_n147, u0_u7_u0_n148, u0_u7_u0_n149, u0_u7_u0_n150, 
       u0_u7_u0_n151, u0_u7_u0_n152, u0_u7_u0_n153, u0_u7_u0_n154, u0_u7_u0_n155, u0_u7_u0_n156, u0_u7_u0_n157, u0_u7_u0_n158, u0_u7_u0_n159, 
       u0_u7_u0_n160, u0_u7_u0_n161, u0_u7_u0_n162, u0_u7_u0_n163, u0_u7_u0_n164, u0_u7_u0_n165, u0_u7_u0_n166, u0_u7_u0_n167, u0_u7_u0_n168, 
       u0_u7_u0_n169, u0_u7_u0_n170, u0_u7_u0_n171, u0_u7_u0_n172, u0_u7_u0_n173, u0_u7_u0_n174, u0_u7_u0_n88, u0_u7_u0_n89, u0_u7_u0_n90, 
       u0_u7_u0_n91, u0_u7_u0_n92, u0_u7_u0_n93, u0_u7_u0_n94, u0_u7_u0_n95, u0_u7_u0_n96, u0_u7_u0_n97, u0_u7_u0_n98, u0_u7_u0_n99, 
       u0_u7_u1_n100, u0_u7_u1_n101, u0_u7_u1_n102, u0_u7_u1_n103, u0_u7_u1_n104, u0_u7_u1_n105, u0_u7_u1_n106, u0_u7_u1_n107, u0_u7_u1_n108, 
       u0_u7_u1_n109, u0_u7_u1_n110, u0_u7_u1_n111, u0_u7_u1_n112, u0_u7_u1_n113, u0_u7_u1_n114, u0_u7_u1_n115, u0_u7_u1_n116, u0_u7_u1_n117, 
       u0_u7_u1_n118, u0_u7_u1_n119, u0_u7_u1_n120, u0_u7_u1_n121, u0_u7_u1_n122, u0_u7_u1_n123, u0_u7_u1_n124, u0_u7_u1_n125, u0_u7_u1_n126, 
       u0_u7_u1_n127, u0_u7_u1_n128, u0_u7_u1_n129, u0_u7_u1_n130, u0_u7_u1_n131, u0_u7_u1_n132, u0_u7_u1_n133, u0_u7_u1_n134, u0_u7_u1_n135, 
       u0_u7_u1_n136, u0_u7_u1_n137, u0_u7_u1_n138, u0_u7_u1_n139, u0_u7_u1_n140, u0_u7_u1_n141, u0_u7_u1_n142, u0_u7_u1_n143, u0_u7_u1_n144, 
       u0_u7_u1_n145, u0_u7_u1_n146, u0_u7_u1_n147, u0_u7_u1_n148, u0_u7_u1_n149, u0_u7_u1_n150, u0_u7_u1_n151, u0_u7_u1_n152, u0_u7_u1_n153, 
       u0_u7_u1_n154, u0_u7_u1_n155, u0_u7_u1_n156, u0_u7_u1_n157, u0_u7_u1_n158, u0_u7_u1_n159, u0_u7_u1_n160, u0_u7_u1_n161, u0_u7_u1_n162, 
       u0_u7_u1_n163, u0_u7_u1_n164, u0_u7_u1_n165, u0_u7_u1_n166, u0_u7_u1_n167, u0_u7_u1_n168, u0_u7_u1_n169, u0_u7_u1_n170, u0_u7_u1_n171, 
       u0_u7_u1_n172, u0_u7_u1_n173, u0_u7_u1_n174, u0_u7_u1_n175, u0_u7_u1_n176, u0_u7_u1_n177, u0_u7_u1_n178, u0_u7_u1_n179, u0_u7_u1_n180, 
       u0_u7_u1_n181, u0_u7_u1_n182, u0_u7_u1_n183, u0_u7_u1_n184, u0_u7_u1_n185, u0_u7_u1_n186, u0_u7_u1_n187, u0_u7_u1_n188, u0_u7_u1_n95, 
       u0_u7_u1_n96, u0_u7_u1_n97, u0_u7_u1_n98, u0_u7_u1_n99, u0_uk_n743, u0_uk_n749, u0_uk_n754, u0_uk_n761, u0_uk_n787, 
       u0_uk_n788, u0_uk_n800, u0_uk_n801, u0_uk_n825, u0_uk_n903, u0_uk_n910, u0_uk_n911, u1_K2_43, u1_K2_44, 
       u1_K2_45, u1_K2_46, u1_K2_47, u1_K2_48, u1_K7_19, u1_K7_20, u1_K7_21, u1_K7_22, u1_K7_23, 
       u1_K7_24, u1_out1_15, u1_out1_21, u1_out1_27, u1_out1_5, u1_out6_1, u1_out6_10, u1_out6_20, u1_out6_26, 
       u1_u1_X_43, u1_u1_X_44, u1_u1_X_45, u1_u1_X_46, u1_u1_X_47, u1_u1_X_48, u1_u1_u7_n100, u1_u1_u7_n101, u1_u1_u7_n102, 
       u1_u1_u7_n103, u1_u1_u7_n104, u1_u1_u7_n105, u1_u1_u7_n106, u1_u1_u7_n107, u1_u1_u7_n108, u1_u1_u7_n109, u1_u1_u7_n110, u1_u1_u7_n111, 
       u1_u1_u7_n112, u1_u1_u7_n113, u1_u1_u7_n114, u1_u1_u7_n115, u1_u1_u7_n116, u1_u1_u7_n117, u1_u1_u7_n118, u1_u1_u7_n119, u1_u1_u7_n120, 
       u1_u1_u7_n121, u1_u1_u7_n122, u1_u1_u7_n123, u1_u1_u7_n124, u1_u1_u7_n125, u1_u1_u7_n126, u1_u1_u7_n127, u1_u1_u7_n128, u1_u1_u7_n129, 
       u1_u1_u7_n130, u1_u1_u7_n131, u1_u1_u7_n132, u1_u1_u7_n133, u1_u1_u7_n134, u1_u1_u7_n135, u1_u1_u7_n136, u1_u1_u7_n137, u1_u1_u7_n138, 
       u1_u1_u7_n139, u1_u1_u7_n140, u1_u1_u7_n141, u1_u1_u7_n142, u1_u1_u7_n143, u1_u1_u7_n144, u1_u1_u7_n145, u1_u1_u7_n146, u1_u1_u7_n147, 
       u1_u1_u7_n148, u1_u1_u7_n149, u1_u1_u7_n150, u1_u1_u7_n151, u1_u1_u7_n152, u1_u1_u7_n153, u1_u1_u7_n154, u1_u1_u7_n155, u1_u1_u7_n156, 
       u1_u1_u7_n157, u1_u1_u7_n158, u1_u1_u7_n159, u1_u1_u7_n160, u1_u1_u7_n161, u1_u1_u7_n162, u1_u1_u7_n163, u1_u1_u7_n164, u1_u1_u7_n165, 
       u1_u1_u7_n166, u1_u1_u7_n167, u1_u1_u7_n168, u1_u1_u7_n169, u1_u1_u7_n170, u1_u1_u7_n171, u1_u1_u7_n172, u1_u1_u7_n173, u1_u1_u7_n174, 
       u1_u1_u7_n175, u1_u1_u7_n176, u1_u1_u7_n177, u1_u1_u7_n178, u1_u1_u7_n179, u1_u1_u7_n180, u1_u1_u7_n91, u1_u1_u7_n92, u1_u1_u7_n93, 
       u1_u1_u7_n94, u1_u1_u7_n95, u1_u1_u7_n96, u1_u1_u7_n97, u1_u1_u7_n98, u1_u1_u7_n99, u1_u6_X_19, u1_u6_X_20, u1_u6_X_21, 
       u1_u6_X_22, u1_u6_X_23, u1_u6_X_24, u1_u6_u3_n100, u1_u6_u3_n101, u1_u6_u3_n102, u1_u6_u3_n103, u1_u6_u3_n104, u1_u6_u3_n105, 
       u1_u6_u3_n106, u1_u6_u3_n107, u1_u6_u3_n108, u1_u6_u3_n109, u1_u6_u3_n110, u1_u6_u3_n111, u1_u6_u3_n112, u1_u6_u3_n113, u1_u6_u3_n114, 
       u1_u6_u3_n115, u1_u6_u3_n116, u1_u6_u3_n117, u1_u6_u3_n118, u1_u6_u3_n119, u1_u6_u3_n120, u1_u6_u3_n121, u1_u6_u3_n122, u1_u6_u3_n123, 
       u1_u6_u3_n124, u1_u6_u3_n125, u1_u6_u3_n126, u1_u6_u3_n127, u1_u6_u3_n128, u1_u6_u3_n129, u1_u6_u3_n130, u1_u6_u3_n131, u1_u6_u3_n132, 
       u1_u6_u3_n133, u1_u6_u3_n134, u1_u6_u3_n135, u1_u6_u3_n136, u1_u6_u3_n137, u1_u6_u3_n138, u1_u6_u3_n139, u1_u6_u3_n140, u1_u6_u3_n141, 
       u1_u6_u3_n142, u1_u6_u3_n143, u1_u6_u3_n144, u1_u6_u3_n145, u1_u6_u3_n146, u1_u6_u3_n147, u1_u6_u3_n148, u1_u6_u3_n149, u1_u6_u3_n150, 
       u1_u6_u3_n151, u1_u6_u3_n152, u1_u6_u3_n153, u1_u6_u3_n154, u1_u6_u3_n155, u1_u6_u3_n156, u1_u6_u3_n157, u1_u6_u3_n158, u1_u6_u3_n159, 
       u1_u6_u3_n160, u1_u6_u3_n161, u1_u6_u3_n162, u1_u6_u3_n163, u1_u6_u3_n164, u1_u6_u3_n165, u1_u6_u3_n166, u1_u6_u3_n167, u1_u6_u3_n168, 
       u1_u6_u3_n169, u1_u6_u3_n170, u1_u6_u3_n171, u1_u6_u3_n172, u1_u6_u3_n173, u1_u6_u3_n174, u1_u6_u3_n175, u1_u6_u3_n176, u1_u6_u3_n177, 
       u1_u6_u3_n178, u1_u6_u3_n179, u1_u6_u3_n180, u1_u6_u3_n181, u1_u6_u3_n182, u1_u6_u3_n183, u1_u6_u3_n184, u1_u6_u3_n185, u1_u6_u3_n186, 
       u1_u6_u3_n94, u1_u6_u3_n95, u1_u6_u3_n96, u1_u6_u3_n97, u1_u6_u3_n98, u1_u6_u3_n99, u1_uk_n1032, u1_uk_n1033, u1_uk_n1109, 
       u1_uk_n1110, u1_uk_n1111, u1_uk_n1112, u1_uk_n1113, u2_K11_43, u2_K11_44, u2_K11_46, u2_K11_47, u2_K14_1, 
       u2_K14_15, u2_K14_2, u2_K14_31, u2_K14_32, u2_K14_33, u2_K14_34, u2_K14_35, u2_K14_36, u2_K14_37, 
       u2_K14_38, u2_K14_4, u2_K14_40, u2_K14_41, u2_K14_5, u2_K14_7, u2_K14_9, u2_K15_25, u2_K15_26, 
       u2_K15_27, u2_K15_30, u2_K15_32, u2_K15_33, u2_K15_36, u2_K15_37, u2_K15_38, u2_K15_40, u2_K15_41, 
       u2_K15_42, u2_K15_43, u2_K15_44, u2_K15_45, u2_K15_46, u2_K15_47, u2_K15_48, u2_K3_10, u2_K3_11, 
       u2_K3_12, u2_K3_8, u2_K3_9, u2_K4_13, u2_K4_15, u2_K4_16, u2_K4_17, u2_K4_18, u2_K4_19, 
       u2_K4_20, u2_K4_23, u2_K4_24, u2_K8_10, u2_K8_11, u2_K8_12, u2_K8_7, u2_K8_9, u2_K9_1, 
       u2_K9_10, u2_K9_11, u2_K9_12, u2_K9_13, u2_K9_14, u2_K9_16, u2_K9_17, u2_K9_18, u2_K9_2, 
       u2_K9_4, u2_K9_6, u2_K9_7, u2_K9_8, u2_K9_9, u2_out10_15, u2_out10_21, u2_out10_27, u2_out10_5, 
       u2_out13_11, u2_out13_12, u2_out13_13, u2_out13_16, u2_out13_17, u2_out13_18, u2_out13_19, u2_out13_2, u2_out13_22, 
       u2_out13_23, u2_out13_24, u2_out13_28, u2_out13_29, u2_out13_30, u2_out13_31, u2_out13_32, u2_out13_4, u2_out13_6, 
       u2_out13_7, u2_out13_9, u2_out14_11, u2_out14_12, u2_out14_14, u2_out14_15, u2_out14_19, u2_out14_21, u2_out14_22, 
       u2_out14_25, u2_out14_27, u2_out14_29, u2_out14_3, u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_7, u2_out14_8, 
       u2_out2_13, u2_out2_18, u2_out2_2, u2_out2_28, u2_out3_1, u2_out3_10, u2_out3_16, u2_out3_20, u2_out3_24, 
       u2_out3_26, u2_out3_30, u2_out3_6, u2_out7_13, u2_out7_18, u2_out7_2, u2_out7_28, u2_out8_13, u2_out8_16, 
       u2_out8_17, u2_out8_18, u2_out8_2, u2_out8_23, u2_out8_24, u2_out8_28, u2_out8_30, u2_out8_31, u2_out8_6, 
       u2_out8_9, u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_47, u2_u10_X_48, u2_u10_u7_n100, u2_u10_u7_n101, 
       u2_u10_u7_n102, u2_u10_u7_n103, u2_u10_u7_n104, u2_u10_u7_n105, u2_u10_u7_n106, u2_u10_u7_n107, u2_u10_u7_n108, u2_u10_u7_n109, u2_u10_u7_n110, 
       u2_u10_u7_n111, u2_u10_u7_n112, u2_u10_u7_n113, u2_u10_u7_n114, u2_u10_u7_n115, u2_u10_u7_n116, u2_u10_u7_n117, u2_u10_u7_n118, u2_u10_u7_n119, 
       u2_u10_u7_n120, u2_u10_u7_n121, u2_u10_u7_n122, u2_u10_u7_n123, u2_u10_u7_n124, u2_u10_u7_n125, u2_u10_u7_n126, u2_u10_u7_n127, u2_u10_u7_n128, 
       u2_u10_u7_n129, u2_u10_u7_n130, u2_u10_u7_n131, u2_u10_u7_n132, u2_u10_u7_n133, u2_u10_u7_n134, u2_u10_u7_n135, u2_u10_u7_n136, u2_u10_u7_n137, 
       u2_u10_u7_n138, u2_u10_u7_n139, u2_u10_u7_n140, u2_u10_u7_n141, u2_u10_u7_n142, u2_u10_u7_n143, u2_u10_u7_n144, u2_u10_u7_n145, u2_u10_u7_n146, 
       u2_u10_u7_n147, u2_u10_u7_n148, u2_u10_u7_n149, u2_u10_u7_n150, u2_u10_u7_n151, u2_u10_u7_n152, u2_u10_u7_n153, u2_u10_u7_n154, u2_u10_u7_n155, 
       u2_u10_u7_n156, u2_u10_u7_n157, u2_u10_u7_n158, u2_u10_u7_n159, u2_u10_u7_n160, u2_u10_u7_n161, u2_u10_u7_n162, u2_u10_u7_n163, u2_u10_u7_n164, 
       u2_u10_u7_n165, u2_u10_u7_n166, u2_u10_u7_n167, u2_u10_u7_n168, u2_u10_u7_n169, u2_u10_u7_n170, u2_u10_u7_n171, u2_u10_u7_n172, u2_u10_u7_n173, 
       u2_u10_u7_n174, u2_u10_u7_n175, u2_u10_u7_n176, u2_u10_u7_n177, u2_u10_u7_n178, u2_u10_u7_n179, u2_u10_u7_n180, u2_u10_u7_n91, u2_u10_u7_n92, 
       u2_u10_u7_n93, u2_u10_u7_n94, u2_u10_u7_n95, u2_u10_u7_n96, u2_u10_u7_n97, u2_u10_u7_n98, u2_u10_u7_n99, u2_u13_X_1, u2_u13_X_10, 
       u2_u13_X_11, u2_u13_X_12, u2_u13_X_13, u2_u13_X_14, u2_u13_X_15, u2_u13_X_16, u2_u13_X_17, u2_u13_X_18, u2_u13_X_2, 
       u2_u13_X_3, u2_u13_X_31, u2_u13_X_32, u2_u13_X_33, u2_u13_X_34, u2_u13_X_35, u2_u13_X_36, u2_u13_X_37, u2_u13_X_38, 
       u2_u13_X_39, u2_u13_X_4, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, u2_u13_X_5, u2_u13_X_6, u2_u13_X_7, u2_u13_X_8, 
       u2_u13_X_9, u2_u13_u0_n100, u2_u13_u0_n101, u2_u13_u0_n102, u2_u13_u0_n103, u2_u13_u0_n104, u2_u13_u0_n105, u2_u13_u0_n106, u2_u13_u0_n107, 
       u2_u13_u0_n108, u2_u13_u0_n109, u2_u13_u0_n110, u2_u13_u0_n111, u2_u13_u0_n112, u2_u13_u0_n113, u2_u13_u0_n114, u2_u13_u0_n115, u2_u13_u0_n116, 
       u2_u13_u0_n117, u2_u13_u0_n118, u2_u13_u0_n119, u2_u13_u0_n120, u2_u13_u0_n121, u2_u13_u0_n122, u2_u13_u0_n123, u2_u13_u0_n124, u2_u13_u0_n125, 
       u2_u13_u0_n126, u2_u13_u0_n127, u2_u13_u0_n128, u2_u13_u0_n129, u2_u13_u0_n130, u2_u13_u0_n131, u2_u13_u0_n132, u2_u13_u0_n133, u2_u13_u0_n134, 
       u2_u13_u0_n135, u2_u13_u0_n136, u2_u13_u0_n137, u2_u13_u0_n138, u2_u13_u0_n139, u2_u13_u0_n140, u2_u13_u0_n141, u2_u13_u0_n142, u2_u13_u0_n143, 
       u2_u13_u0_n144, u2_u13_u0_n145, u2_u13_u0_n146, u2_u13_u0_n147, u2_u13_u0_n148, u2_u13_u0_n149, u2_u13_u0_n150, u2_u13_u0_n151, u2_u13_u0_n152, 
       u2_u13_u0_n153, u2_u13_u0_n154, u2_u13_u0_n155, u2_u13_u0_n156, u2_u13_u0_n157, u2_u13_u0_n158, u2_u13_u0_n159, u2_u13_u0_n160, u2_u13_u0_n161, 
       u2_u13_u0_n162, u2_u13_u0_n163, u2_u13_u0_n164, u2_u13_u0_n165, u2_u13_u0_n166, u2_u13_u0_n167, u2_u13_u0_n168, u2_u13_u0_n169, u2_u13_u0_n170, 
       u2_u13_u0_n171, u2_u13_u0_n172, u2_u13_u0_n173, u2_u13_u0_n174, u2_u13_u0_n88, u2_u13_u0_n89, u2_u13_u0_n90, u2_u13_u0_n91, u2_u13_u0_n92, 
       u2_u13_u0_n93, u2_u13_u0_n94, u2_u13_u0_n95, u2_u13_u0_n96, u2_u13_u0_n97, u2_u13_u0_n98, u2_u13_u0_n99, u2_u13_u1_n100, u2_u13_u1_n101, 
       u2_u13_u1_n102, u2_u13_u1_n103, u2_u13_u1_n104, u2_u13_u1_n105, u2_u13_u1_n106, u2_u13_u1_n107, u2_u13_u1_n108, u2_u13_u1_n109, u2_u13_u1_n110, 
       u2_u13_u1_n111, u2_u13_u1_n112, u2_u13_u1_n113, u2_u13_u1_n114, u2_u13_u1_n115, u2_u13_u1_n116, u2_u13_u1_n117, u2_u13_u1_n118, u2_u13_u1_n119, 
       u2_u13_u1_n120, u2_u13_u1_n121, u2_u13_u1_n122, u2_u13_u1_n123, u2_u13_u1_n124, u2_u13_u1_n125, u2_u13_u1_n126, u2_u13_u1_n127, u2_u13_u1_n128, 
       u2_u13_u1_n129, u2_u13_u1_n130, u2_u13_u1_n131, u2_u13_u1_n132, u2_u13_u1_n133, u2_u13_u1_n134, u2_u13_u1_n135, u2_u13_u1_n136, u2_u13_u1_n137, 
       u2_u13_u1_n138, u2_u13_u1_n139, u2_u13_u1_n140, u2_u13_u1_n141, u2_u13_u1_n142, u2_u13_u1_n143, u2_u13_u1_n144, u2_u13_u1_n145, u2_u13_u1_n146, 
       u2_u13_u1_n147, u2_u13_u1_n148, u2_u13_u1_n149, u2_u13_u1_n150, u2_u13_u1_n151, u2_u13_u1_n152, u2_u13_u1_n153, u2_u13_u1_n154, u2_u13_u1_n155, 
       u2_u13_u1_n156, u2_u13_u1_n157, u2_u13_u1_n158, u2_u13_u1_n159, u2_u13_u1_n160, u2_u13_u1_n161, u2_u13_u1_n162, u2_u13_u1_n163, u2_u13_u1_n164, 
       u2_u13_u1_n165, u2_u13_u1_n166, u2_u13_u1_n167, u2_u13_u1_n168, u2_u13_u1_n169, u2_u13_u1_n170, u2_u13_u1_n171, u2_u13_u1_n172, u2_u13_u1_n173, 
       u2_u13_u1_n174, u2_u13_u1_n175, u2_u13_u1_n176, u2_u13_u1_n177, u2_u13_u1_n178, u2_u13_u1_n179, u2_u13_u1_n180, u2_u13_u1_n181, u2_u13_u1_n182, 
       u2_u13_u1_n183, u2_u13_u1_n184, u2_u13_u1_n185, u2_u13_u1_n186, u2_u13_u1_n187, u2_u13_u1_n188, u2_u13_u1_n95, u2_u13_u1_n96, u2_u13_u1_n97, 
       u2_u13_u1_n98, u2_u13_u1_n99, u2_u13_u2_n100, u2_u13_u2_n101, u2_u13_u2_n102, u2_u13_u2_n103, u2_u13_u2_n104, u2_u13_u2_n105, u2_u13_u2_n106, 
       u2_u13_u2_n107, u2_u13_u2_n108, u2_u13_u2_n109, u2_u13_u2_n110, u2_u13_u2_n111, u2_u13_u2_n112, u2_u13_u2_n113, u2_u13_u2_n114, u2_u13_u2_n115, 
       u2_u13_u2_n116, u2_u13_u2_n117, u2_u13_u2_n118, u2_u13_u2_n119, u2_u13_u2_n120, u2_u13_u2_n121, u2_u13_u2_n122, u2_u13_u2_n123, u2_u13_u2_n124, 
       u2_u13_u2_n125, u2_u13_u2_n126, u2_u13_u2_n127, u2_u13_u2_n128, u2_u13_u2_n129, u2_u13_u2_n130, u2_u13_u2_n131, u2_u13_u2_n132, u2_u13_u2_n133, 
       u2_u13_u2_n134, u2_u13_u2_n135, u2_u13_u2_n136, u2_u13_u2_n137, u2_u13_u2_n138, u2_u13_u2_n139, u2_u13_u2_n140, u2_u13_u2_n141, u2_u13_u2_n142, 
       u2_u13_u2_n143, u2_u13_u2_n144, u2_u13_u2_n145, u2_u13_u2_n146, u2_u13_u2_n147, u2_u13_u2_n148, u2_u13_u2_n149, u2_u13_u2_n150, u2_u13_u2_n151, 
       u2_u13_u2_n152, u2_u13_u2_n153, u2_u13_u2_n154, u2_u13_u2_n155, u2_u13_u2_n156, u2_u13_u2_n157, u2_u13_u2_n158, u2_u13_u2_n159, u2_u13_u2_n160, 
       u2_u13_u2_n161, u2_u13_u2_n162, u2_u13_u2_n163, u2_u13_u2_n164, u2_u13_u2_n165, u2_u13_u2_n166, u2_u13_u2_n167, u2_u13_u2_n168, u2_u13_u2_n169, 
       u2_u13_u2_n170, u2_u13_u2_n171, u2_u13_u2_n172, u2_u13_u2_n173, u2_u13_u2_n174, u2_u13_u2_n175, u2_u13_u2_n176, u2_u13_u2_n177, u2_u13_u2_n178, 
       u2_u13_u2_n179, u2_u13_u2_n180, u2_u13_u2_n181, u2_u13_u2_n182, u2_u13_u2_n183, u2_u13_u2_n184, u2_u13_u2_n185, u2_u13_u2_n186, u2_u13_u2_n187, 
       u2_u13_u2_n188, u2_u13_u2_n95, u2_u13_u2_n96, u2_u13_u2_n97, u2_u13_u2_n98, u2_u13_u2_n99, u2_u13_u5_n100, u2_u13_u5_n101, u2_u13_u5_n102, 
       u2_u13_u5_n103, u2_u13_u5_n104, u2_u13_u5_n105, u2_u13_u5_n106, u2_u13_u5_n107, u2_u13_u5_n108, u2_u13_u5_n109, u2_u13_u5_n110, u2_u13_u5_n111, 
       u2_u13_u5_n112, u2_u13_u5_n113, u2_u13_u5_n114, u2_u13_u5_n115, u2_u13_u5_n116, u2_u13_u5_n117, u2_u13_u5_n118, u2_u13_u5_n119, u2_u13_u5_n120, 
       u2_u13_u5_n121, u2_u13_u5_n122, u2_u13_u5_n123, u2_u13_u5_n124, u2_u13_u5_n125, u2_u13_u5_n126, u2_u13_u5_n127, u2_u13_u5_n128, u2_u13_u5_n129, 
       u2_u13_u5_n130, u2_u13_u5_n131, u2_u13_u5_n132, u2_u13_u5_n133, u2_u13_u5_n134, u2_u13_u5_n135, u2_u13_u5_n136, u2_u13_u5_n137, u2_u13_u5_n138, 
       u2_u13_u5_n139, u2_u13_u5_n140, u2_u13_u5_n141, u2_u13_u5_n142, u2_u13_u5_n143, u2_u13_u5_n144, u2_u13_u5_n145, u2_u13_u5_n146, u2_u13_u5_n147, 
       u2_u13_u5_n148, u2_u13_u5_n149, u2_u13_u5_n150, u2_u13_u5_n151, u2_u13_u5_n152, u2_u13_u5_n153, u2_u13_u5_n154, u2_u13_u5_n155, u2_u13_u5_n156, 
       u2_u13_u5_n157, u2_u13_u5_n158, u2_u13_u5_n159, u2_u13_u5_n160, u2_u13_u5_n161, u2_u13_u5_n162, u2_u13_u5_n163, u2_u13_u5_n164, u2_u13_u5_n165, 
       u2_u13_u5_n166, u2_u13_u5_n167, u2_u13_u5_n168, u2_u13_u5_n169, u2_u13_u5_n170, u2_u13_u5_n171, u2_u13_u5_n172, u2_u13_u5_n173, u2_u13_u5_n174, 
       u2_u13_u5_n175, u2_u13_u5_n176, u2_u13_u5_n177, u2_u13_u5_n178, u2_u13_u5_n179, u2_u13_u5_n180, u2_u13_u5_n181, u2_u13_u5_n182, u2_u13_u5_n183, 
       u2_u13_u5_n184, u2_u13_u5_n185, u2_u13_u5_n186, u2_u13_u5_n187, u2_u13_u5_n188, u2_u13_u5_n189, u2_u13_u5_n190, u2_u13_u5_n191, u2_u13_u5_n192, 
       u2_u13_u5_n193, u2_u13_u5_n194, u2_u13_u5_n195, u2_u13_u5_n196, u2_u13_u5_n99, u2_u13_u6_n100, u2_u13_u6_n101, u2_u13_u6_n102, u2_u13_u6_n103, 
       u2_u13_u6_n104, u2_u13_u6_n105, u2_u13_u6_n106, u2_u13_u6_n107, u2_u13_u6_n108, u2_u13_u6_n109, u2_u13_u6_n110, u2_u13_u6_n111, u2_u13_u6_n112, 
       u2_u13_u6_n113, u2_u13_u6_n114, u2_u13_u6_n115, u2_u13_u6_n116, u2_u13_u6_n117, u2_u13_u6_n118, u2_u13_u6_n119, u2_u13_u6_n120, u2_u13_u6_n121, 
       u2_u13_u6_n122, u2_u13_u6_n123, u2_u13_u6_n124, u2_u13_u6_n125, u2_u13_u6_n126, u2_u13_u6_n127, u2_u13_u6_n128, u2_u13_u6_n129, u2_u13_u6_n130, 
       u2_u13_u6_n131, u2_u13_u6_n132, u2_u13_u6_n133, u2_u13_u6_n134, u2_u13_u6_n135, u2_u13_u6_n136, u2_u13_u6_n137, u2_u13_u6_n138, u2_u13_u6_n139, 
       u2_u13_u6_n140, u2_u13_u6_n141, u2_u13_u6_n142, u2_u13_u6_n143, u2_u13_u6_n144, u2_u13_u6_n145, u2_u13_u6_n146, u2_u13_u6_n147, u2_u13_u6_n148, 
       u2_u13_u6_n149, u2_u13_u6_n150, u2_u13_u6_n151, u2_u13_u6_n152, u2_u13_u6_n153, u2_u13_u6_n154, u2_u13_u6_n155, u2_u13_u6_n156, u2_u13_u6_n157, 
       u2_u13_u6_n158, u2_u13_u6_n159, u2_u13_u6_n160, u2_u13_u6_n161, u2_u13_u6_n162, u2_u13_u6_n163, u2_u13_u6_n164, u2_u13_u6_n165, u2_u13_u6_n166, 
       u2_u13_u6_n167, u2_u13_u6_n168, u2_u13_u6_n169, u2_u13_u6_n170, u2_u13_u6_n171, u2_u13_u6_n172, u2_u13_u6_n173, u2_u13_u6_n174, u2_u13_u6_n88, 
       u2_u13_u6_n89, u2_u13_u6_n90, u2_u13_u6_n91, u2_u13_u6_n92, u2_u13_u6_n93, u2_u13_u6_n94, u2_u13_u6_n95, u2_u13_u6_n96, u2_u13_u6_n97, 
       u2_u13_u6_n98, u2_u13_u6_n99, u2_u14_X_25, u2_u14_X_26, u2_u14_X_27, u2_u14_X_28, u2_u14_X_29, u2_u14_X_30, u2_u14_X_31, 
       u2_u14_X_32, u2_u14_X_33, u2_u14_X_34, u2_u14_X_35, u2_u14_X_36, u2_u14_X_37, u2_u14_X_38, u2_u14_X_39, u2_u14_X_40, 
       u2_u14_X_41, u2_u14_X_42, u2_u14_X_43, u2_u14_X_44, u2_u14_X_45, u2_u14_X_46, u2_u14_X_47, u2_u14_X_48, u2_u14_u4_n100, 
       u2_u14_u4_n101, u2_u14_u4_n102, u2_u14_u4_n103, u2_u14_u4_n104, u2_u14_u4_n105, u2_u14_u4_n106, u2_u14_u4_n107, u2_u14_u4_n108, u2_u14_u4_n109, 
       u2_u14_u4_n110, u2_u14_u4_n111, u2_u14_u4_n112, u2_u14_u4_n113, u2_u14_u4_n114, u2_u14_u4_n115, u2_u14_u4_n116, u2_u14_u4_n117, u2_u14_u4_n118, 
       u2_u14_u4_n119, u2_u14_u4_n120, u2_u14_u4_n121, u2_u14_u4_n122, u2_u14_u4_n123, u2_u14_u4_n124, u2_u14_u4_n125, u2_u14_u4_n126, u2_u14_u4_n127, 
       u2_u14_u4_n128, u2_u14_u4_n129, u2_u14_u4_n130, u2_u14_u4_n131, u2_u14_u4_n132, u2_u14_u4_n133, u2_u14_u4_n134, u2_u14_u4_n135, u2_u14_u4_n136, 
       u2_u14_u4_n137, u2_u14_u4_n138, u2_u14_u4_n139, u2_u14_u4_n140, u2_u14_u4_n141, u2_u14_u4_n142, u2_u14_u4_n143, u2_u14_u4_n144, u2_u14_u4_n145, 
       u2_u14_u4_n146, u2_u14_u4_n147, u2_u14_u4_n148, u2_u14_u4_n149, u2_u14_u4_n150, u2_u14_u4_n151, u2_u14_u4_n152, u2_u14_u4_n153, u2_u14_u4_n154, 
       u2_u14_u4_n155, u2_u14_u4_n156, u2_u14_u4_n157, u2_u14_u4_n158, u2_u14_u4_n159, u2_u14_u4_n160, u2_u14_u4_n161, u2_u14_u4_n162, u2_u14_u4_n163, 
       u2_u14_u4_n164, u2_u14_u4_n165, u2_u14_u4_n166, u2_u14_u4_n167, u2_u14_u4_n168, u2_u14_u4_n169, u2_u14_u4_n170, u2_u14_u4_n171, u2_u14_u4_n172, 
       u2_u14_u4_n173, u2_u14_u4_n174, u2_u14_u4_n175, u2_u14_u4_n176, u2_u14_u4_n177, u2_u14_u4_n178, u2_u14_u4_n179, u2_u14_u4_n180, u2_u14_u4_n181, 
       u2_u14_u4_n182, u2_u14_u4_n183, u2_u14_u4_n184, u2_u14_u4_n185, u2_u14_u4_n186, u2_u14_u4_n94, u2_u14_u4_n95, u2_u14_u4_n96, u2_u14_u4_n97, 
       u2_u14_u4_n98, u2_u14_u4_n99, u2_u14_u5_n100, u2_u14_u5_n101, u2_u14_u5_n102, u2_u14_u5_n103, u2_u14_u5_n104, u2_u14_u5_n105, u2_u14_u5_n106, 
       u2_u14_u5_n107, u2_u14_u5_n108, u2_u14_u5_n109, u2_u14_u5_n110, u2_u14_u5_n111, u2_u14_u5_n112, u2_u14_u5_n113, u2_u14_u5_n114, u2_u14_u5_n115, 
       u2_u14_u5_n116, u2_u14_u5_n117, u2_u14_u5_n118, u2_u14_u5_n119, u2_u14_u5_n120, u2_u14_u5_n121, u2_u14_u5_n122, u2_u14_u5_n123, u2_u14_u5_n124, 
       u2_u14_u5_n125, u2_u14_u5_n126, u2_u14_u5_n127, u2_u14_u5_n128, u2_u14_u5_n129, u2_u14_u5_n130, u2_u14_u5_n131, u2_u14_u5_n132, u2_u14_u5_n133, 
       u2_u14_u5_n134, u2_u14_u5_n135, u2_u14_u5_n136, u2_u14_u5_n137, u2_u14_u5_n138, u2_u14_u5_n139, u2_u14_u5_n140, u2_u14_u5_n141, u2_u14_u5_n142, 
       u2_u14_u5_n143, u2_u14_u5_n144, u2_u14_u5_n145, u2_u14_u5_n146, u2_u14_u5_n147, u2_u14_u5_n148, u2_u14_u5_n149, u2_u14_u5_n150, u2_u14_u5_n151, 
       u2_u14_u5_n152, u2_u14_u5_n153, u2_u14_u5_n154, u2_u14_u5_n155, u2_u14_u5_n156, u2_u14_u5_n157, u2_u14_u5_n158, u2_u14_u5_n159, u2_u14_u5_n160, 
       u2_u14_u5_n161, u2_u14_u5_n162, u2_u14_u5_n163, u2_u14_u5_n164, u2_u14_u5_n165, u2_u14_u5_n166, u2_u14_u5_n167, u2_u14_u5_n168, u2_u14_u5_n169, 
       u2_u14_u5_n170, u2_u14_u5_n171, u2_u14_u5_n172, u2_u14_u5_n173, u2_u14_u5_n174, u2_u14_u5_n175, u2_u14_u5_n176, u2_u14_u5_n177, u2_u14_u5_n178, 
       u2_u14_u5_n179, u2_u14_u5_n180, u2_u14_u5_n181, u2_u14_u5_n182, u2_u14_u5_n183, u2_u14_u5_n184, u2_u14_u5_n185, u2_u14_u5_n186, u2_u14_u5_n187, 
       u2_u14_u5_n188, u2_u14_u5_n189, u2_u14_u5_n190, u2_u14_u5_n191, u2_u14_u5_n192, u2_u14_u5_n193, u2_u14_u5_n194, u2_u14_u5_n195, u2_u14_u5_n196, 
       u2_u14_u5_n99, u2_u14_u6_n100, u2_u14_u6_n101, u2_u14_u6_n102, u2_u14_u6_n103, u2_u14_u6_n104, u2_u14_u6_n105, u2_u14_u6_n106, u2_u14_u6_n107, 
       u2_u14_u6_n108, u2_u14_u6_n109, u2_u14_u6_n110, u2_u14_u6_n111, u2_u14_u6_n112, u2_u14_u6_n113, u2_u14_u6_n114, u2_u14_u6_n115, u2_u14_u6_n116, 
       u2_u14_u6_n117, u2_u14_u6_n118, u2_u14_u6_n119, u2_u14_u6_n120, u2_u14_u6_n121, u2_u14_u6_n122, u2_u14_u6_n123, u2_u14_u6_n124, u2_u14_u6_n125, 
       u2_u14_u6_n126, u2_u14_u6_n127, u2_u14_u6_n128, u2_u14_u6_n129, u2_u14_u6_n130, u2_u14_u6_n131, u2_u14_u6_n132, u2_u14_u6_n133, u2_u14_u6_n134, 
       u2_u14_u6_n135, u2_u14_u6_n136, u2_u14_u6_n137, u2_u14_u6_n138, u2_u14_u6_n139, u2_u14_u6_n140, u2_u14_u6_n141, u2_u14_u6_n142, u2_u14_u6_n143, 
       u2_u14_u6_n144, u2_u14_u6_n145, u2_u14_u6_n146, u2_u14_u6_n147, u2_u14_u6_n148, u2_u14_u6_n149, u2_u14_u6_n150, u2_u14_u6_n151, u2_u14_u6_n152, 
       u2_u14_u6_n153, u2_u14_u6_n154, u2_u14_u6_n155, u2_u14_u6_n156, u2_u14_u6_n157, u2_u14_u6_n158, u2_u14_u6_n159, u2_u14_u6_n160, u2_u14_u6_n161, 
       u2_u14_u6_n162, u2_u14_u6_n163, u2_u14_u6_n164, u2_u14_u6_n165, u2_u14_u6_n166, u2_u14_u6_n167, u2_u14_u6_n168, u2_u14_u6_n169, u2_u14_u6_n170, 
       u2_u14_u6_n171, u2_u14_u6_n172, u2_u14_u6_n173, u2_u14_u6_n174, u2_u14_u6_n88, u2_u14_u6_n89, u2_u14_u6_n90, u2_u14_u6_n91, u2_u14_u6_n92, 
       u2_u14_u6_n93, u2_u14_u6_n94, u2_u14_u6_n95, u2_u14_u6_n96, u2_u14_u6_n97, u2_u14_u6_n98, u2_u14_u6_n99, u2_u14_u7_n100, u2_u14_u7_n101, 
       u2_u14_u7_n102, u2_u14_u7_n103, u2_u14_u7_n104, u2_u14_u7_n105, u2_u14_u7_n106, u2_u14_u7_n107, u2_u14_u7_n108, u2_u14_u7_n109, u2_u14_u7_n110, 
       u2_u14_u7_n111, u2_u14_u7_n112, u2_u14_u7_n113, u2_u14_u7_n114, u2_u14_u7_n115, u2_u14_u7_n116, u2_u14_u7_n117, u2_u14_u7_n118, u2_u14_u7_n119, 
       u2_u14_u7_n120, u2_u14_u7_n121, u2_u14_u7_n122, u2_u14_u7_n123, u2_u14_u7_n124, u2_u14_u7_n125, u2_u14_u7_n126, u2_u14_u7_n127, u2_u14_u7_n128, 
       u2_u14_u7_n129, u2_u14_u7_n130, u2_u14_u7_n131, u2_u14_u7_n132, u2_u14_u7_n133, u2_u14_u7_n134, u2_u14_u7_n135, u2_u14_u7_n136, u2_u14_u7_n137, 
       u2_u14_u7_n138, u2_u14_u7_n139, u2_u14_u7_n140, u2_u14_u7_n141, u2_u14_u7_n142, u2_u14_u7_n143, u2_u14_u7_n144, u2_u14_u7_n145, u2_u14_u7_n146, 
       u2_u14_u7_n147, u2_u14_u7_n148, u2_u14_u7_n149, u2_u14_u7_n150, u2_u14_u7_n151, u2_u14_u7_n152, u2_u14_u7_n153, u2_u14_u7_n154, u2_u14_u7_n155, 
       u2_u14_u7_n156, u2_u14_u7_n157, u2_u14_u7_n158, u2_u14_u7_n159, u2_u14_u7_n160, u2_u14_u7_n161, u2_u14_u7_n162, u2_u14_u7_n163, u2_u14_u7_n164, 
       u2_u14_u7_n165, u2_u14_u7_n166, u2_u14_u7_n167, u2_u14_u7_n168, u2_u14_u7_n169, u2_u14_u7_n170, u2_u14_u7_n171, u2_u14_u7_n172, u2_u14_u7_n173, 
       u2_u14_u7_n174, u2_u14_u7_n175, u2_u14_u7_n176, u2_u14_u7_n177, u2_u14_u7_n178, u2_u14_u7_n179, u2_u14_u7_n180, u2_u14_u7_n91, u2_u14_u7_n92, 
       u2_u14_u7_n93, u2_u14_u7_n94, u2_u14_u7_n95, u2_u14_u7_n96, u2_u14_u7_n97, u2_u14_u7_n98, u2_u14_u7_n99, u2_u2_X_10, u2_u2_X_11, 
       u2_u2_X_12, u2_u2_X_7, u2_u2_X_8, u2_u2_X_9, u2_u2_u1_n100, u2_u2_u1_n101, u2_u2_u1_n102, u2_u2_u1_n103, u2_u2_u1_n104, 
       u2_u2_u1_n105, u2_u2_u1_n106, u2_u2_u1_n107, u2_u2_u1_n108, u2_u2_u1_n109, u2_u2_u1_n110, u2_u2_u1_n111, u2_u2_u1_n112, u2_u2_u1_n113, 
       u2_u2_u1_n114, u2_u2_u1_n115, u2_u2_u1_n116, u2_u2_u1_n117, u2_u2_u1_n118, u2_u2_u1_n119, u2_u2_u1_n120, u2_u2_u1_n121, u2_u2_u1_n122, 
       u2_u2_u1_n123, u2_u2_u1_n124, u2_u2_u1_n125, u2_u2_u1_n126, u2_u2_u1_n127, u2_u2_u1_n128, u2_u2_u1_n129, u2_u2_u1_n130, u2_u2_u1_n131, 
       u2_u2_u1_n132, u2_u2_u1_n133, u2_u2_u1_n134, u2_u2_u1_n135, u2_u2_u1_n136, u2_u2_u1_n137, u2_u2_u1_n138, u2_u2_u1_n139, u2_u2_u1_n140, 
       u2_u2_u1_n141, u2_u2_u1_n142, u2_u2_u1_n143, u2_u2_u1_n144, u2_u2_u1_n145, u2_u2_u1_n146, u2_u2_u1_n147, u2_u2_u1_n148, u2_u2_u1_n149, 
       u2_u2_u1_n150, u2_u2_u1_n151, u2_u2_u1_n152, u2_u2_u1_n153, u2_u2_u1_n154, u2_u2_u1_n155, u2_u2_u1_n156, u2_u2_u1_n157, u2_u2_u1_n158, 
       u2_u2_u1_n159, u2_u2_u1_n160, u2_u2_u1_n161, u2_u2_u1_n162, u2_u2_u1_n163, u2_u2_u1_n164, u2_u2_u1_n165, u2_u2_u1_n166, u2_u2_u1_n167, 
       u2_u2_u1_n168, u2_u2_u1_n169, u2_u2_u1_n170, u2_u2_u1_n171, u2_u2_u1_n172, u2_u2_u1_n173, u2_u2_u1_n174, u2_u2_u1_n175, u2_u2_u1_n176, 
       u2_u2_u1_n177, u2_u2_u1_n178, u2_u2_u1_n179, u2_u2_u1_n180, u2_u2_u1_n181, u2_u2_u1_n182, u2_u2_u1_n183, u2_u2_u1_n184, u2_u2_u1_n185, 
       u2_u2_u1_n186, u2_u2_u1_n187, u2_u2_u1_n188, u2_u2_u1_n95, u2_u2_u1_n96, u2_u2_u1_n97, u2_u2_u1_n98, u2_u2_u1_n99, u2_u3_X_13, 
       u2_u3_X_14, u2_u3_X_15, u2_u3_X_16, u2_u3_X_17, u2_u3_X_18, u2_u3_X_19, u2_u3_X_20, u2_u3_X_21, u2_u3_X_22, 
       u2_u3_X_23, u2_u3_X_24, u2_u3_u2_n100, u2_u3_u2_n101, u2_u3_u2_n102, u2_u3_u2_n103, u2_u3_u2_n104, u2_u3_u2_n105, u2_u3_u2_n106, 
       u2_u3_u2_n107, u2_u3_u2_n108, u2_u3_u2_n109, u2_u3_u2_n110, u2_u3_u2_n111, u2_u3_u2_n112, u2_u3_u2_n113, u2_u3_u2_n114, u2_u3_u2_n115, 
       u2_u3_u2_n116, u2_u3_u2_n117, u2_u3_u2_n118, u2_u3_u2_n119, u2_u3_u2_n120, u2_u3_u2_n121, u2_u3_u2_n122, u2_u3_u2_n123, u2_u3_u2_n124, 
       u2_u3_u2_n125, u2_u3_u2_n126, u2_u3_u2_n127, u2_u3_u2_n128, u2_u3_u2_n129, u2_u3_u2_n130, u2_u3_u2_n131, u2_u3_u2_n132, u2_u3_u2_n133, 
       u2_u3_u2_n134, u2_u3_u2_n135, u2_u3_u2_n136, u2_u3_u2_n137, u2_u3_u2_n138, u2_u3_u2_n139, u2_u3_u2_n140, u2_u3_u2_n141, u2_u3_u2_n142, 
       u2_u3_u2_n143, u2_u3_u2_n144, u2_u3_u2_n145, u2_u3_u2_n146, u2_u3_u2_n147, u2_u3_u2_n148, u2_u3_u2_n149, u2_u3_u2_n150, u2_u3_u2_n151, 
       u2_u3_u2_n152, u2_u3_u2_n153, u2_u3_u2_n154, u2_u3_u2_n155, u2_u3_u2_n156, u2_u3_u2_n157, u2_u3_u2_n158, u2_u3_u2_n159, u2_u3_u2_n160, 
       u2_u3_u2_n161, u2_u3_u2_n162, u2_u3_u2_n163, u2_u3_u2_n164, u2_u3_u2_n165, u2_u3_u2_n166, u2_u3_u2_n167, u2_u3_u2_n168, u2_u3_u2_n169, 
       u2_u3_u2_n170, u2_u3_u2_n171, u2_u3_u2_n172, u2_u3_u2_n173, u2_u3_u2_n174, u2_u3_u2_n175, u2_u3_u2_n176, u2_u3_u2_n177, u2_u3_u2_n178, 
       u2_u3_u2_n179, u2_u3_u2_n180, u2_u3_u2_n181, u2_u3_u2_n182, u2_u3_u2_n183, u2_u3_u2_n184, u2_u3_u2_n185, u2_u3_u2_n186, u2_u3_u2_n187, 
       u2_u3_u2_n188, u2_u3_u2_n95, u2_u3_u2_n96, u2_u3_u2_n97, u2_u3_u2_n98, u2_u3_u2_n99, u2_u3_u3_n100, u2_u3_u3_n101, u2_u3_u3_n102, 
       u2_u3_u3_n103, u2_u3_u3_n104, u2_u3_u3_n105, u2_u3_u3_n106, u2_u3_u3_n107, u2_u3_u3_n108, u2_u3_u3_n109, u2_u3_u3_n110, u2_u3_u3_n111, 
       u2_u3_u3_n112, u2_u3_u3_n113, u2_u3_u3_n114, u2_u3_u3_n115, u2_u3_u3_n116, u2_u3_u3_n117, u2_u3_u3_n118, u2_u3_u3_n119, u2_u3_u3_n120, 
       u2_u3_u3_n121, u2_u3_u3_n122, u2_u3_u3_n123, u2_u3_u3_n124, u2_u3_u3_n125, u2_u3_u3_n126, u2_u3_u3_n127, u2_u3_u3_n128, u2_u3_u3_n129, 
       u2_u3_u3_n130, u2_u3_u3_n131, u2_u3_u3_n132, u2_u3_u3_n133, u2_u3_u3_n134, u2_u3_u3_n135, u2_u3_u3_n136, u2_u3_u3_n137, u2_u3_u3_n138, 
       u2_u3_u3_n139, u2_u3_u3_n140, u2_u3_u3_n141, u2_u3_u3_n142, u2_u3_u3_n143, u2_u3_u3_n144, u2_u3_u3_n145, u2_u3_u3_n146, u2_u3_u3_n147, 
       u2_u3_u3_n148, u2_u3_u3_n149, u2_u3_u3_n150, u2_u3_u3_n151, u2_u3_u3_n152, u2_u3_u3_n153, u2_u3_u3_n154, u2_u3_u3_n155, u2_u3_u3_n156, 
       u2_u3_u3_n157, u2_u3_u3_n158, u2_u3_u3_n159, u2_u3_u3_n160, u2_u3_u3_n161, u2_u3_u3_n162, u2_u3_u3_n163, u2_u3_u3_n164, u2_u3_u3_n165, 
       u2_u3_u3_n166, u2_u3_u3_n167, u2_u3_u3_n168, u2_u3_u3_n169, u2_u3_u3_n170, u2_u3_u3_n171, u2_u3_u3_n172, u2_u3_u3_n173, u2_u3_u3_n174, 
       u2_u3_u3_n175, u2_u3_u3_n176, u2_u3_u3_n177, u2_u3_u3_n178, u2_u3_u3_n179, u2_u3_u3_n180, u2_u3_u3_n181, u2_u3_u3_n182, u2_u3_u3_n183, 
       u2_u3_u3_n184, u2_u3_u3_n185, u2_u3_u3_n186, u2_u3_u3_n94, u2_u3_u3_n95, u2_u3_u3_n96, u2_u3_u3_n97, u2_u3_u3_n98, u2_u3_u3_n99, 
       u2_u7_X_10, u2_u7_X_11, u2_u7_X_12, u2_u7_X_7, u2_u7_X_8, u2_u7_X_9, u2_u7_u1_n100, u2_u7_u1_n101, u2_u7_u1_n102, 
       u2_u7_u1_n103, u2_u7_u1_n104, u2_u7_u1_n105, u2_u7_u1_n106, u2_u7_u1_n107, u2_u7_u1_n108, u2_u7_u1_n109, u2_u7_u1_n110, u2_u7_u1_n111, 
       u2_u7_u1_n112, u2_u7_u1_n113, u2_u7_u1_n114, u2_u7_u1_n115, u2_u7_u1_n116, u2_u7_u1_n117, u2_u7_u1_n118, u2_u7_u1_n119, u2_u7_u1_n120, 
       u2_u7_u1_n121, u2_u7_u1_n122, u2_u7_u1_n123, u2_u7_u1_n124, u2_u7_u1_n125, u2_u7_u1_n126, u2_u7_u1_n127, u2_u7_u1_n128, u2_u7_u1_n129, 
       u2_u7_u1_n130, u2_u7_u1_n131, u2_u7_u1_n132, u2_u7_u1_n133, u2_u7_u1_n134, u2_u7_u1_n135, u2_u7_u1_n136, u2_u7_u1_n137, u2_u7_u1_n138, 
       u2_u7_u1_n139, u2_u7_u1_n140, u2_u7_u1_n141, u2_u7_u1_n142, u2_u7_u1_n143, u2_u7_u1_n144, u2_u7_u1_n145, u2_u7_u1_n146, u2_u7_u1_n147, 
       u2_u7_u1_n148, u2_u7_u1_n149, u2_u7_u1_n150, u2_u7_u1_n151, u2_u7_u1_n152, u2_u7_u1_n153, u2_u7_u1_n154, u2_u7_u1_n155, u2_u7_u1_n156, 
       u2_u7_u1_n157, u2_u7_u1_n158, u2_u7_u1_n159, u2_u7_u1_n160, u2_u7_u1_n161, u2_u7_u1_n162, u2_u7_u1_n163, u2_u7_u1_n164, u2_u7_u1_n165, 
       u2_u7_u1_n166, u2_u7_u1_n167, u2_u7_u1_n168, u2_u7_u1_n169, u2_u7_u1_n170, u2_u7_u1_n171, u2_u7_u1_n172, u2_u7_u1_n173, u2_u7_u1_n174, 
       u2_u7_u1_n175, u2_u7_u1_n176, u2_u7_u1_n177, u2_u7_u1_n178, u2_u7_u1_n179, u2_u7_u1_n180, u2_u7_u1_n181, u2_u7_u1_n182, u2_u7_u1_n183, 
       u2_u7_u1_n184, u2_u7_u1_n185, u2_u7_u1_n186, u2_u7_u1_n187, u2_u7_u1_n188, u2_u7_u1_n95, u2_u7_u1_n96, u2_u7_u1_n97, u2_u7_u1_n98, 
       u2_u7_u1_n99, u2_u8_X_1, u2_u8_X_10, u2_u8_X_11, u2_u8_X_12, u2_u8_X_13, u2_u8_X_14, u2_u8_X_15, u2_u8_X_16, 
       u2_u8_X_17, u2_u8_X_18, u2_u8_X_2, u2_u8_X_3, u2_u8_X_4, u2_u8_X_5, u2_u8_X_6, u2_u8_X_7, u2_u8_X_8, 
       u2_u8_X_9, u2_u8_u0_n100, u2_u8_u0_n101, u2_u8_u0_n102, u2_u8_u0_n103, u2_u8_u0_n104, u2_u8_u0_n105, u2_u8_u0_n106, u2_u8_u0_n107, 
       u2_u8_u0_n108, u2_u8_u0_n109, u2_u8_u0_n110, u2_u8_u0_n111, u2_u8_u0_n112, u2_u8_u0_n113, u2_u8_u0_n114, u2_u8_u0_n115, u2_u8_u0_n116, 
       u2_u8_u0_n117, u2_u8_u0_n118, u2_u8_u0_n119, u2_u8_u0_n120, u2_u8_u0_n121, u2_u8_u0_n122, u2_u8_u0_n123, u2_u8_u0_n124, u2_u8_u0_n125, 
       u2_u8_u0_n126, u2_u8_u0_n127, u2_u8_u0_n128, u2_u8_u0_n129, u2_u8_u0_n130, u2_u8_u0_n131, u2_u8_u0_n132, u2_u8_u0_n133, u2_u8_u0_n134, 
       u2_u8_u0_n135, u2_u8_u0_n136, u2_u8_u0_n137, u2_u8_u0_n138, u2_u8_u0_n139, u2_u8_u0_n140, u2_u8_u0_n141, u2_u8_u0_n142, u2_u8_u0_n143, 
       u2_u8_u0_n144, u2_u8_u0_n145, u2_u8_u0_n146, u2_u8_u0_n147, u2_u8_u0_n148, u2_u8_u0_n149, u2_u8_u0_n150, u2_u8_u0_n151, u2_u8_u0_n152, 
       u2_u8_u0_n153, u2_u8_u0_n154, u2_u8_u0_n155, u2_u8_u0_n156, u2_u8_u0_n157, u2_u8_u0_n158, u2_u8_u0_n159, u2_u8_u0_n160, u2_u8_u0_n161, 
       u2_u8_u0_n162, u2_u8_u0_n163, u2_u8_u0_n164, u2_u8_u0_n165, u2_u8_u0_n166, u2_u8_u0_n167, u2_u8_u0_n168, u2_u8_u0_n169, u2_u8_u0_n170, 
       u2_u8_u0_n171, u2_u8_u0_n172, u2_u8_u0_n173, u2_u8_u0_n174, u2_u8_u0_n88, u2_u8_u0_n89, u2_u8_u0_n90, u2_u8_u0_n91, u2_u8_u0_n92, 
       u2_u8_u0_n93, u2_u8_u0_n94, u2_u8_u0_n95, u2_u8_u0_n96, u2_u8_u0_n97, u2_u8_u0_n98, u2_u8_u0_n99, u2_u8_u1_n100, u2_u8_u1_n101, 
       u2_u8_u1_n102, u2_u8_u1_n103, u2_u8_u1_n104, u2_u8_u1_n105, u2_u8_u1_n106, u2_u8_u1_n107, u2_u8_u1_n108, u2_u8_u1_n109, u2_u8_u1_n110, 
       u2_u8_u1_n111, u2_u8_u1_n112, u2_u8_u1_n113, u2_u8_u1_n114, u2_u8_u1_n115, u2_u8_u1_n116, u2_u8_u1_n117, u2_u8_u1_n118, u2_u8_u1_n119, 
       u2_u8_u1_n120, u2_u8_u1_n121, u2_u8_u1_n122, u2_u8_u1_n123, u2_u8_u1_n124, u2_u8_u1_n125, u2_u8_u1_n126, u2_u8_u1_n127, u2_u8_u1_n128, 
       u2_u8_u1_n129, u2_u8_u1_n130, u2_u8_u1_n131, u2_u8_u1_n132, u2_u8_u1_n133, u2_u8_u1_n134, u2_u8_u1_n135, u2_u8_u1_n136, u2_u8_u1_n137, 
       u2_u8_u1_n138, u2_u8_u1_n139, u2_u8_u1_n140, u2_u8_u1_n141, u2_u8_u1_n142, u2_u8_u1_n143, u2_u8_u1_n144, u2_u8_u1_n145, u2_u8_u1_n146, 
       u2_u8_u1_n147, u2_u8_u1_n148, u2_u8_u1_n149, u2_u8_u1_n150, u2_u8_u1_n151, u2_u8_u1_n152, u2_u8_u1_n153, u2_u8_u1_n154, u2_u8_u1_n155, 
       u2_u8_u1_n156, u2_u8_u1_n157, u2_u8_u1_n158, u2_u8_u1_n159, u2_u8_u1_n160, u2_u8_u1_n161, u2_u8_u1_n162, u2_u8_u1_n163, u2_u8_u1_n164, 
       u2_u8_u1_n165, u2_u8_u1_n166, u2_u8_u1_n167, u2_u8_u1_n168, u2_u8_u1_n169, u2_u8_u1_n170, u2_u8_u1_n171, u2_u8_u1_n172, u2_u8_u1_n173, 
       u2_u8_u1_n174, u2_u8_u1_n175, u2_u8_u1_n176, u2_u8_u1_n177, u2_u8_u1_n178, u2_u8_u1_n179, u2_u8_u1_n180, u2_u8_u1_n181, u2_u8_u1_n182, 
       u2_u8_u1_n183, u2_u8_u1_n184, u2_u8_u1_n185, u2_u8_u1_n186, u2_u8_u1_n187, u2_u8_u1_n188, u2_u8_u1_n95, u2_u8_u1_n96, u2_u8_u1_n97, 
       u2_u8_u1_n98, u2_u8_u1_n99, u2_u8_u2_n100, u2_u8_u2_n101, u2_u8_u2_n102, u2_u8_u2_n103, u2_u8_u2_n104, u2_u8_u2_n105, u2_u8_u2_n106, 
       u2_u8_u2_n107, u2_u8_u2_n108, u2_u8_u2_n109, u2_u8_u2_n110, u2_u8_u2_n111, u2_u8_u2_n112, u2_u8_u2_n113, u2_u8_u2_n114, u2_u8_u2_n115, 
       u2_u8_u2_n116, u2_u8_u2_n117, u2_u8_u2_n118, u2_u8_u2_n119, u2_u8_u2_n120, u2_u8_u2_n121, u2_u8_u2_n122, u2_u8_u2_n123, u2_u8_u2_n124, 
       u2_u8_u2_n125, u2_u8_u2_n126, u2_u8_u2_n127, u2_u8_u2_n128, u2_u8_u2_n129, u2_u8_u2_n130, u2_u8_u2_n131, u2_u8_u2_n132, u2_u8_u2_n133, 
       u2_u8_u2_n134, u2_u8_u2_n135, u2_u8_u2_n136, u2_u8_u2_n137, u2_u8_u2_n138, u2_u8_u2_n139, u2_u8_u2_n140, u2_u8_u2_n141, u2_u8_u2_n142, 
       u2_u8_u2_n143, u2_u8_u2_n144, u2_u8_u2_n145, u2_u8_u2_n146, u2_u8_u2_n147, u2_u8_u2_n148, u2_u8_u2_n149, u2_u8_u2_n150, u2_u8_u2_n151, 
       u2_u8_u2_n152, u2_u8_u2_n153, u2_u8_u2_n154, u2_u8_u2_n155, u2_u8_u2_n156, u2_u8_u2_n157, u2_u8_u2_n158, u2_u8_u2_n159, u2_u8_u2_n160, 
       u2_u8_u2_n161, u2_u8_u2_n162, u2_u8_u2_n163, u2_u8_u2_n164, u2_u8_u2_n165, u2_u8_u2_n166, u2_u8_u2_n167, u2_u8_u2_n168, u2_u8_u2_n169, 
       u2_u8_u2_n170, u2_u8_u2_n171, u2_u8_u2_n172, u2_u8_u2_n173, u2_u8_u2_n174, u2_u8_u2_n175, u2_u8_u2_n176, u2_u8_u2_n177, u2_u8_u2_n178, 
       u2_u8_u2_n179, u2_u8_u2_n180, u2_u8_u2_n181, u2_u8_u2_n182, u2_u8_u2_n183, u2_u8_u2_n184, u2_u8_u2_n185, u2_u8_u2_n186, u2_u8_u2_n187, 
       u2_u8_u2_n188, u2_u8_u2_n95, u2_u8_u2_n96, u2_u8_u2_n97, u2_u8_u2_n98, u2_u8_u2_n99, u2_uk_n1019, u2_uk_n1021, u2_uk_n1026, 
       u2_uk_n1098, u2_uk_n1117, u2_uk_n1118, u2_uk_n1122, u2_uk_n1123, u2_uk_n386, u2_uk_n692, u2_uk_n694, u2_uk_n932, 
       u2_uk_n938,  u2_uk_n940;
  XOR2_X1 u0_U309 (.B( u0_L6_31 ) , .Z( u0_N254 ) , .A( u0_out7_31 ) );
  XOR2_X1 u0_U312 (.B( u0_L6_28 ) , .Z( u0_N251 ) , .A( u0_out7_28 ) );
  XOR2_X1 u0_U318 (.B( u0_L6_23 ) , .Z( u0_N246 ) , .A( u0_out7_23 ) );
  XOR2_X1 u0_U323 (.B( u0_L6_18 ) , .Z( u0_N241 ) , .A( u0_out7_18 ) );
  XOR2_X1 u0_U324 (.B( u0_L6_17 ) , .Z( u0_N240 ) , .A( u0_out7_17 ) );
  XOR2_X1 u0_U329 (.B( u0_L6_13 ) , .Z( u0_N236 ) , .A( u0_out7_13 ) );
  XOR2_X1 u0_U333 (.B( u0_L6_9 ) , .Z( u0_N232 ) , .A( u0_out7_9 ) );
  XOR2_X1 u0_U341 (.B( u0_L6_2 ) , .Z( u0_N225 ) , .A( u0_out7_2 ) );
  XOR2_X1 u0_U380 (.B( u0_L4_31 ) , .Z( u0_N190 ) , .A( u0_out5_31 ) );
  XOR2_X1 u0_U382 (.B( u0_L4_30 ) , .Z( u0_N189 ) , .A( u0_out5_30 ) );
  XOR2_X1 u0_U384 (.B( u0_L4_28 ) , .Z( u0_N187 ) , .A( u0_out5_28 ) );
  XOR2_X1 u0_U388 (.B( u0_L4_24 ) , .Z( u0_N183 ) , .A( u0_out5_24 ) );
  XOR2_X1 u0_U389 (.B( u0_L4_23 ) , .Z( u0_N182 ) , .A( u0_out5_23 ) );
  XOR2_X1 u0_U395 (.B( u0_L4_18 ) , .Z( u0_N177 ) , .A( u0_out5_18 ) );
  XOR2_X1 u0_U396 (.B( u0_L4_17 ) , .Z( u0_N176 ) , .A( u0_out5_17 ) );
  XOR2_X1 u0_U397 (.B( u0_L4_16 ) , .Z( u0_N175 ) , .A( u0_out5_16 ) );
  XOR2_X1 u0_U400 (.B( u0_L4_13 ) , .Z( u0_N172 ) , .A( u0_out5_13 ) );
  XOR2_X1 u0_U405 (.B( u0_L4_9 ) , .Z( u0_N168 ) , .A( u0_out5_9 ) );
  XOR2_X1 u0_U408 (.B( u0_L4_6 ) , .Z( u0_N165 ) , .A( u0_out5_6 ) );
  XOR2_X1 u0_U412 (.B( u0_L4_2 ) , .Z( u0_N161 ) , .A( u0_out5_2 ) );
  XOR2_X1 u0_U450 (.B( u0_L2_32 ) , .Z( u0_N127 ) , .A( u0_out3_32 ) );
  XOR2_X1 u0_U455 (.B( u0_L2_27 ) , .Z( u0_N122 ) , .A( u0_out3_27 ) );
  XOR2_X1 u0_U461 (.B( u0_L2_22 ) , .Z( u0_N117 ) , .A( u0_out3_22 ) );
  XOR2_X1 u0_U462 (.B( u0_L2_21 ) , .Z( u0_N116 ) , .A( u0_out3_21 ) );
  XOR2_X1 u0_U468 (.B( u0_L2_15 ) , .Z( u0_N110 ) , .A( u0_out3_15 ) );
  XOR2_X1 u0_U472 (.B( u0_L2_12 ) , .Z( u0_N107 ) , .A( u0_out3_12 ) );
  XOR2_X1 u0_U477 (.B( u0_L2_7 ) , .Z( u0_N102 ) , .A( u0_out3_7 ) );
  XOR2_X1 u0_U479 (.B( u0_L2_5 ) , .Z( u0_N100 ) , .A( u0_out3_5 ) );
  XOR2_X1 u0_U483 (.Z( u0_FP_9 ) , .B( u0_L14_9 ) , .A( u0_out15_9 ) );
  XOR2_X1 u0_U491 (.Z( u0_FP_31 ) , .B( u0_L14_31 ) , .A( u0_out15_31 ) );
  XOR2_X1 u0_U493 (.Z( u0_FP_2 ) , .B( u0_L14_2 ) , .A( u0_out15_2 ) );
  XOR2_X1 u0_U495 (.Z( u0_FP_28 ) , .B( u0_L14_28 ) , .A( u0_out15_28 ) );
  XOR2_X1 u0_U500 (.Z( u0_FP_23 ) , .B( u0_L14_23 ) , .A( u0_out15_23 ) );
  XOR2_X1 u0_U506 (.Z( u0_FP_18 ) , .B( u0_L14_18 ) , .A( u0_out15_18 ) );
  XOR2_X1 u0_U507 (.Z( u0_FP_17 ) , .B( u0_L14_17 ) , .A( u0_out15_17 ) );
  XOR2_X1 u0_U511 (.Z( u0_FP_13 ) , .B( u0_L14_13 ) , .A( u0_out15_13 ) );
  XOR2_X1 u0_u15_U1 (.A( u0_FP_38 ) , .B( u0_K16_9 ) , .Z( u0_u15_X_9 ) );
  XOR2_X1 u0_u15_U16 (.A( u0_FP_34 ) , .B( u0_K16_3 ) , .Z( u0_u15_X_3 ) );
  XOR2_X1 u0_u15_U2 (.A( u0_FP_37 ) , .B( u0_K16_8 ) , .Z( u0_u15_X_8 ) );
  XOR2_X1 u0_u15_U27 (.A( u0_FP_33 ) , .B( u0_K16_2 ) , .Z( u0_u15_X_2 ) );
  XOR2_X1 u0_u15_U3 (.A( u0_FP_36 ) , .B( u0_K16_7 ) , .Z( u0_u15_X_7 ) );
  XOR2_X1 u0_u15_U38 (.A( u0_FP_64 ) , .B( u0_K16_1 ) , .Z( u0_u15_X_1 ) );
  XOR2_X1 u0_u15_U4 (.A( u0_FP_37 ) , .B( u0_K16_6 ) , .Z( u0_u15_X_6 ) );
  XOR2_X1 u0_u15_U46 (.A( u0_FP_41 ) , .B( u0_K16_12 ) , .Z( u0_u15_X_12 ) );
  XOR2_X1 u0_u15_U47 (.A( u0_FP_40 ) , .B( u0_K16_11 ) , .Z( u0_u15_X_11 ) );
  XOR2_X1 u0_u15_U48 (.A( u0_FP_39 ) , .B( u0_K16_10 ) , .Z( u0_u15_X_10 ) );
  XOR2_X1 u0_u15_U5 (.A( u0_FP_36 ) , .B( u0_K16_5 ) , .Z( u0_u15_X_5 ) );
  XOR2_X1 u0_u15_U6 (.A( u0_FP_35 ) , .B( u0_K16_4 ) , .Z( u0_u15_X_4 ) );
  AND3_X1 u0_u15_u0_U10 (.A2( u0_u15_u0_n112 ) , .ZN( u0_u15_u0_n127 ) , .A3( u0_u15_u0_n130 ) , .A1( u0_u15_u0_n148 ) );
  NAND2_X1 u0_u15_u0_U11 (.ZN( u0_u15_u0_n113 ) , .A1( u0_u15_u0_n139 ) , .A2( u0_u15_u0_n149 ) );
  AND2_X1 u0_u15_u0_U12 (.ZN( u0_u15_u0_n107 ) , .A1( u0_u15_u0_n130 ) , .A2( u0_u15_u0_n140 ) );
  AND2_X1 u0_u15_u0_U13 (.A2( u0_u15_u0_n129 ) , .A1( u0_u15_u0_n130 ) , .ZN( u0_u15_u0_n151 ) );
  AND2_X1 u0_u15_u0_U14 (.A1( u0_u15_u0_n108 ) , .A2( u0_u15_u0_n125 ) , .ZN( u0_u15_u0_n145 ) );
  INV_X1 u0_u15_u0_U15 (.A( u0_u15_u0_n143 ) , .ZN( u0_u15_u0_n173 ) );
  NOR2_X1 u0_u15_u0_U16 (.A2( u0_u15_u0_n136 ) , .ZN( u0_u15_u0_n147 ) , .A1( u0_u15_u0_n160 ) );
  AOI21_X1 u0_u15_u0_U17 (.B1( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n132 ) , .A( u0_u15_u0_n165 ) , .B2( u0_u15_u0_n93 ) );
  INV_X1 u0_u15_u0_U18 (.A( u0_u15_u0_n142 ) , .ZN( u0_u15_u0_n165 ) );
  OAI221_X1 u0_u15_u0_U19 (.C1( u0_u15_u0_n121 ) , .ZN( u0_u15_u0_n122 ) , .B2( u0_u15_u0_n127 ) , .A( u0_u15_u0_n143 ) , .B1( u0_u15_u0_n144 ) , .C2( u0_u15_u0_n147 ) );
  OAI22_X1 u0_u15_u0_U20 (.B1( u0_u15_u0_n131 ) , .A1( u0_u15_u0_n144 ) , .B2( u0_u15_u0_n147 ) , .A2( u0_u15_u0_n90 ) , .ZN( u0_u15_u0_n91 ) );
  AND3_X1 u0_u15_u0_U21 (.A3( u0_u15_u0_n121 ) , .A2( u0_u15_u0_n125 ) , .A1( u0_u15_u0_n148 ) , .ZN( u0_u15_u0_n90 ) );
  OAI22_X1 u0_u15_u0_U22 (.B1( u0_u15_u0_n125 ) , .ZN( u0_u15_u0_n126 ) , .A1( u0_u15_u0_n138 ) , .A2( u0_u15_u0_n146 ) , .B2( u0_u15_u0_n147 ) );
  NOR2_X1 u0_u15_u0_U23 (.A1( u0_u15_u0_n163 ) , .A2( u0_u15_u0_n164 ) , .ZN( u0_u15_u0_n95 ) );
  INV_X1 u0_u15_u0_U24 (.A( u0_u15_u0_n136 ) , .ZN( u0_u15_u0_n161 ) );
  NOR2_X1 u0_u15_u0_U25 (.A1( u0_u15_u0_n120 ) , .ZN( u0_u15_u0_n143 ) , .A2( u0_u15_u0_n167 ) );
  OAI221_X1 u0_u15_u0_U26 (.C1( u0_u15_u0_n112 ) , .ZN( u0_u15_u0_n120 ) , .B1( u0_u15_u0_n138 ) , .B2( u0_u15_u0_n141 ) , .C2( u0_u15_u0_n147 ) , .A( u0_u15_u0_n172 ) );
  AOI211_X1 u0_u15_u0_U27 (.B( u0_u15_u0_n115 ) , .A( u0_u15_u0_n116 ) , .C2( u0_u15_u0_n117 ) , .C1( u0_u15_u0_n118 ) , .ZN( u0_u15_u0_n119 ) );
  AOI22_X1 u0_u15_u0_U28 (.B2( u0_u15_u0_n109 ) , .A2( u0_u15_u0_n110 ) , .ZN( u0_u15_u0_n111 ) , .B1( u0_u15_u0_n118 ) , .A1( u0_u15_u0_n160 ) );
  NAND2_X1 u0_u15_u0_U29 (.A2( u0_u15_u0_n102 ) , .A1( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n149 ) );
  INV_X1 u0_u15_u0_U3 (.A( u0_u15_u0_n113 ) , .ZN( u0_u15_u0_n166 ) );
  INV_X1 u0_u15_u0_U30 (.A( u0_u15_u0_n118 ) , .ZN( u0_u15_u0_n158 ) );
  NAND2_X1 u0_u15_u0_U31 (.A2( u0_u15_u0_n100 ) , .ZN( u0_u15_u0_n131 ) , .A1( u0_u15_u0_n92 ) );
  NAND2_X1 u0_u15_u0_U32 (.ZN( u0_u15_u0_n108 ) , .A1( u0_u15_u0_n92 ) , .A2( u0_u15_u0_n94 ) );
  AOI21_X1 u0_u15_u0_U33 (.ZN( u0_u15_u0_n104 ) , .B1( u0_u15_u0_n107 ) , .B2( u0_u15_u0_n141 ) , .A( u0_u15_u0_n144 ) );
  AOI21_X1 u0_u15_u0_U34 (.B1( u0_u15_u0_n127 ) , .B2( u0_u15_u0_n129 ) , .A( u0_u15_u0_n138 ) , .ZN( u0_u15_u0_n96 ) );
  NAND2_X1 u0_u15_u0_U35 (.A2( u0_u15_u0_n102 ) , .ZN( u0_u15_u0_n114 ) , .A1( u0_u15_u0_n92 ) );
  AOI21_X1 u0_u15_u0_U36 (.ZN( u0_u15_u0_n116 ) , .B2( u0_u15_u0_n142 ) , .A( u0_u15_u0_n144 ) , .B1( u0_u15_u0_n166 ) );
  NAND2_X1 u0_u15_u0_U37 (.A2( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n140 ) , .A1( u0_u15_u0_n94 ) );
  NAND2_X1 u0_u15_u0_U38 (.A1( u0_u15_u0_n100 ) , .A2( u0_u15_u0_n103 ) , .ZN( u0_u15_u0_n125 ) );
  NAND2_X1 u0_u15_u0_U39 (.A1( u0_u15_u0_n101 ) , .A2( u0_u15_u0_n102 ) , .ZN( u0_u15_u0_n150 ) );
  AOI21_X1 u0_u15_u0_U4 (.B1( u0_u15_u0_n114 ) , .ZN( u0_u15_u0_n115 ) , .B2( u0_u15_u0_n129 ) , .A( u0_u15_u0_n161 ) );
  INV_X1 u0_u15_u0_U40 (.A( u0_u15_u0_n138 ) , .ZN( u0_u15_u0_n160 ) );
  NAND2_X1 u0_u15_u0_U41 (.A2( u0_u15_u0_n100 ) , .A1( u0_u15_u0_n101 ) , .ZN( u0_u15_u0_n139 ) );
  NAND2_X1 u0_u15_u0_U42 (.ZN( u0_u15_u0_n112 ) , .A2( u0_u15_u0_n92 ) , .A1( u0_u15_u0_n93 ) );
  NAND2_X1 u0_u15_u0_U43 (.A1( u0_u15_u0_n101 ) , .ZN( u0_u15_u0_n130 ) , .A2( u0_u15_u0_n94 ) );
  NAND2_X1 u0_u15_u0_U44 (.A2( u0_u15_u0_n101 ) , .ZN( u0_u15_u0_n121 ) , .A1( u0_u15_u0_n93 ) );
  INV_X1 u0_u15_u0_U45 (.ZN( u0_u15_u0_n172 ) , .A( u0_u15_u0_n88 ) );
  OAI222_X1 u0_u15_u0_U46 (.C1( u0_u15_u0_n108 ) , .A1( u0_u15_u0_n125 ) , .B2( u0_u15_u0_n128 ) , .B1( u0_u15_u0_n144 ) , .A2( u0_u15_u0_n158 ) , .C2( u0_u15_u0_n161 ) , .ZN( u0_u15_u0_n88 ) );
  OR3_X1 u0_u15_u0_U47 (.A3( u0_u15_u0_n152 ) , .A2( u0_u15_u0_n153 ) , .A1( u0_u15_u0_n154 ) , .ZN( u0_u15_u0_n155 ) );
  AOI21_X1 u0_u15_u0_U48 (.B2( u0_u15_u0_n150 ) , .B1( u0_u15_u0_n151 ) , .ZN( u0_u15_u0_n152 ) , .A( u0_u15_u0_n158 ) );
  AOI21_X1 u0_u15_u0_U49 (.A( u0_u15_u0_n144 ) , .B2( u0_u15_u0_n145 ) , .B1( u0_u15_u0_n146 ) , .ZN( u0_u15_u0_n154 ) );
  AOI21_X1 u0_u15_u0_U5 (.B2( u0_u15_u0_n131 ) , .ZN( u0_u15_u0_n134 ) , .B1( u0_u15_u0_n151 ) , .A( u0_u15_u0_n158 ) );
  AOI21_X1 u0_u15_u0_U50 (.A( u0_u15_u0_n147 ) , .B2( u0_u15_u0_n148 ) , .B1( u0_u15_u0_n149 ) , .ZN( u0_u15_u0_n153 ) );
  INV_X1 u0_u15_u0_U51 (.ZN( u0_u15_u0_n171 ) , .A( u0_u15_u0_n99 ) );
  OAI211_X1 u0_u15_u0_U52 (.C2( u0_u15_u0_n140 ) , .C1( u0_u15_u0_n161 ) , .A( u0_u15_u0_n169 ) , .B( u0_u15_u0_n98 ) , .ZN( u0_u15_u0_n99 ) );
  AOI211_X1 u0_u15_u0_U53 (.C1( u0_u15_u0_n118 ) , .A( u0_u15_u0_n123 ) , .B( u0_u15_u0_n96 ) , .C2( u0_u15_u0_n97 ) , .ZN( u0_u15_u0_n98 ) );
  INV_X1 u0_u15_u0_U54 (.ZN( u0_u15_u0_n169 ) , .A( u0_u15_u0_n91 ) );
  NOR2_X1 u0_u15_u0_U55 (.A2( u0_u15_X_4 ) , .A1( u0_u15_X_5 ) , .ZN( u0_u15_u0_n118 ) );
  NOR2_X1 u0_u15_u0_U56 (.A2( u0_u15_X_1 ) , .ZN( u0_u15_u0_n101 ) , .A1( u0_u15_u0_n163 ) );
  NOR2_X1 u0_u15_u0_U57 (.A2( u0_u15_X_3 ) , .A1( u0_u15_X_6 ) , .ZN( u0_u15_u0_n94 ) );
  NOR2_X1 u0_u15_u0_U58 (.A2( u0_u15_X_6 ) , .ZN( u0_u15_u0_n100 ) , .A1( u0_u15_u0_n162 ) );
  NAND2_X1 u0_u15_u0_U59 (.A2( u0_u15_X_4 ) , .A1( u0_u15_X_5 ) , .ZN( u0_u15_u0_n144 ) );
  NOR2_X1 u0_u15_u0_U6 (.A1( u0_u15_u0_n108 ) , .ZN( u0_u15_u0_n123 ) , .A2( u0_u15_u0_n158 ) );
  NOR2_X1 u0_u15_u0_U60 (.A2( u0_u15_X_5 ) , .ZN( u0_u15_u0_n136 ) , .A1( u0_u15_u0_n159 ) );
  NAND2_X1 u0_u15_u0_U61 (.A1( u0_u15_X_5 ) , .ZN( u0_u15_u0_n138 ) , .A2( u0_u15_u0_n159 ) );
  AND2_X1 u0_u15_u0_U62 (.A2( u0_u15_X_3 ) , .A1( u0_u15_X_6 ) , .ZN( u0_u15_u0_n102 ) );
  AND2_X1 u0_u15_u0_U63 (.A1( u0_u15_X_6 ) , .A2( u0_u15_u0_n162 ) , .ZN( u0_u15_u0_n93 ) );
  INV_X1 u0_u15_u0_U64 (.A( u0_u15_X_4 ) , .ZN( u0_u15_u0_n159 ) );
  INV_X1 u0_u15_u0_U65 (.A( u0_u15_X_1 ) , .ZN( u0_u15_u0_n164 ) );
  INV_X1 u0_u15_u0_U66 (.A( u0_u15_X_3 ) , .ZN( u0_u15_u0_n162 ) );
  INV_X1 u0_u15_u0_U67 (.A( u0_u15_u0_n126 ) , .ZN( u0_u15_u0_n168 ) );
  AOI211_X1 u0_u15_u0_U68 (.B( u0_u15_u0_n133 ) , .A( u0_u15_u0_n134 ) , .C2( u0_u15_u0_n135 ) , .C1( u0_u15_u0_n136 ) , .ZN( u0_u15_u0_n137 ) );
  INV_X1 u0_u15_u0_U69 (.ZN( u0_u15_u0_n174 ) , .A( u0_u15_u0_n89 ) );
  OAI21_X1 u0_u15_u0_U7 (.B1( u0_u15_u0_n150 ) , .B2( u0_u15_u0_n158 ) , .A( u0_u15_u0_n172 ) , .ZN( u0_u15_u0_n89 ) );
  AOI211_X1 u0_u15_u0_U70 (.B( u0_u15_u0_n104 ) , .A( u0_u15_u0_n105 ) , .ZN( u0_u15_u0_n106 ) , .C2( u0_u15_u0_n113 ) , .C1( u0_u15_u0_n160 ) );
  OR4_X1 u0_u15_u0_U71 (.ZN( u0_out15_17 ) , .A4( u0_u15_u0_n122 ) , .A2( u0_u15_u0_n123 ) , .A1( u0_u15_u0_n124 ) , .A3( u0_u15_u0_n170 ) );
  AOI21_X1 u0_u15_u0_U72 (.B2( u0_u15_u0_n107 ) , .ZN( u0_u15_u0_n124 ) , .B1( u0_u15_u0_n128 ) , .A( u0_u15_u0_n161 ) );
  INV_X1 u0_u15_u0_U73 (.A( u0_u15_u0_n111 ) , .ZN( u0_u15_u0_n170 ) );
  OR4_X1 u0_u15_u0_U74 (.ZN( u0_out15_31 ) , .A4( u0_u15_u0_n155 ) , .A2( u0_u15_u0_n156 ) , .A1( u0_u15_u0_n157 ) , .A3( u0_u15_u0_n173 ) );
  AOI21_X1 u0_u15_u0_U75 (.A( u0_u15_u0_n138 ) , .B2( u0_u15_u0_n139 ) , .B1( u0_u15_u0_n140 ) , .ZN( u0_u15_u0_n157 ) );
  AOI21_X1 u0_u15_u0_U76 (.B2( u0_u15_u0_n141 ) , .B1( u0_u15_u0_n142 ) , .ZN( u0_u15_u0_n156 ) , .A( u0_u15_u0_n161 ) );
  AOI21_X1 u0_u15_u0_U77 (.B1( u0_u15_u0_n132 ) , .ZN( u0_u15_u0_n133 ) , .A( u0_u15_u0_n144 ) , .B2( u0_u15_u0_n166 ) );
  OAI22_X1 u0_u15_u0_U78 (.ZN( u0_u15_u0_n105 ) , .A2( u0_u15_u0_n132 ) , .B1( u0_u15_u0_n146 ) , .A1( u0_u15_u0_n147 ) , .B2( u0_u15_u0_n161 ) );
  NAND2_X1 u0_u15_u0_U79 (.ZN( u0_u15_u0_n110 ) , .A2( u0_u15_u0_n132 ) , .A1( u0_u15_u0_n145 ) );
  AND2_X1 u0_u15_u0_U8 (.A1( u0_u15_u0_n114 ) , .A2( u0_u15_u0_n121 ) , .ZN( u0_u15_u0_n146 ) );
  INV_X1 u0_u15_u0_U80 (.A( u0_u15_u0_n119 ) , .ZN( u0_u15_u0_n167 ) );
  NAND2_X1 u0_u15_u0_U81 (.ZN( u0_u15_u0_n148 ) , .A1( u0_u15_u0_n93 ) , .A2( u0_u15_u0_n95 ) );
  NAND2_X1 u0_u15_u0_U82 (.A1( u0_u15_u0_n100 ) , .ZN( u0_u15_u0_n129 ) , .A2( u0_u15_u0_n95 ) );
  NAND2_X1 u0_u15_u0_U83 (.A1( u0_u15_u0_n102 ) , .ZN( u0_u15_u0_n128 ) , .A2( u0_u15_u0_n95 ) );
  NOR2_X1 u0_u15_u0_U84 (.A2( u0_u15_X_1 ) , .A1( u0_u15_X_2 ) , .ZN( u0_u15_u0_n92 ) );
  NAND2_X1 u0_u15_u0_U85 (.ZN( u0_u15_u0_n142 ) , .A1( u0_u15_u0_n94 ) , .A2( u0_u15_u0_n95 ) );
  NOR2_X1 u0_u15_u0_U86 (.A2( u0_u15_X_2 ) , .ZN( u0_u15_u0_n103 ) , .A1( u0_u15_u0_n164 ) );
  INV_X1 u0_u15_u0_U87 (.A( u0_u15_X_2 ) , .ZN( u0_u15_u0_n163 ) );
  NAND3_X1 u0_u15_u0_U88 (.ZN( u0_out15_23 ) , .A3( u0_u15_u0_n137 ) , .A1( u0_u15_u0_n168 ) , .A2( u0_u15_u0_n171 ) );
  NAND3_X1 u0_u15_u0_U89 (.A3( u0_u15_u0_n127 ) , .A2( u0_u15_u0_n128 ) , .ZN( u0_u15_u0_n135 ) , .A1( u0_u15_u0_n150 ) );
  AND2_X1 u0_u15_u0_U9 (.A1( u0_u15_u0_n131 ) , .ZN( u0_u15_u0_n141 ) , .A2( u0_u15_u0_n150 ) );
  NAND3_X1 u0_u15_u0_U90 (.ZN( u0_u15_u0_n117 ) , .A3( u0_u15_u0_n132 ) , .A2( u0_u15_u0_n139 ) , .A1( u0_u15_u0_n148 ) );
  NAND3_X1 u0_u15_u0_U91 (.ZN( u0_u15_u0_n109 ) , .A2( u0_u15_u0_n114 ) , .A3( u0_u15_u0_n140 ) , .A1( u0_u15_u0_n149 ) );
  NAND3_X1 u0_u15_u0_U92 (.ZN( u0_out15_9 ) , .A3( u0_u15_u0_n106 ) , .A2( u0_u15_u0_n171 ) , .A1( u0_u15_u0_n174 ) );
  NAND3_X1 u0_u15_u0_U93 (.A2( u0_u15_u0_n128 ) , .A1( u0_u15_u0_n132 ) , .A3( u0_u15_u0_n146 ) , .ZN( u0_u15_u0_n97 ) );
  NOR2_X1 u0_u15_u1_U10 (.A1( u0_u15_u1_n112 ) , .A2( u0_u15_u1_n116 ) , .ZN( u0_u15_u1_n118 ) );
  NAND3_X1 u0_u15_u1_U100 (.ZN( u0_u15_u1_n113 ) , .A1( u0_u15_u1_n120 ) , .A3( u0_u15_u1_n133 ) , .A2( u0_u15_u1_n155 ) );
  OAI21_X1 u0_u15_u1_U11 (.ZN( u0_u15_u1_n101 ) , .B1( u0_u15_u1_n141 ) , .A( u0_u15_u1_n146 ) , .B2( u0_u15_u1_n183 ) );
  AOI21_X1 u0_u15_u1_U12 (.B2( u0_u15_u1_n155 ) , .B1( u0_u15_u1_n156 ) , .ZN( u0_u15_u1_n157 ) , .A( u0_u15_u1_n174 ) );
  NAND2_X1 u0_u15_u1_U13 (.ZN( u0_u15_u1_n140 ) , .A2( u0_u15_u1_n150 ) , .A1( u0_u15_u1_n155 ) );
  NAND2_X1 u0_u15_u1_U14 (.A1( u0_u15_u1_n131 ) , .ZN( u0_u15_u1_n147 ) , .A2( u0_u15_u1_n153 ) );
  INV_X1 u0_u15_u1_U15 (.A( u0_u15_u1_n139 ) , .ZN( u0_u15_u1_n174 ) );
  OR4_X1 u0_u15_u1_U16 (.A4( u0_u15_u1_n106 ) , .A3( u0_u15_u1_n107 ) , .ZN( u0_u15_u1_n108 ) , .A1( u0_u15_u1_n117 ) , .A2( u0_u15_u1_n184 ) );
  AOI21_X1 u0_u15_u1_U17 (.ZN( u0_u15_u1_n106 ) , .A( u0_u15_u1_n112 ) , .B1( u0_u15_u1_n154 ) , .B2( u0_u15_u1_n156 ) );
  AOI21_X1 u0_u15_u1_U18 (.ZN( u0_u15_u1_n107 ) , .B1( u0_u15_u1_n134 ) , .B2( u0_u15_u1_n149 ) , .A( u0_u15_u1_n174 ) );
  INV_X1 u0_u15_u1_U19 (.A( u0_u15_u1_n101 ) , .ZN( u0_u15_u1_n184 ) );
  INV_X1 u0_u15_u1_U20 (.A( u0_u15_u1_n112 ) , .ZN( u0_u15_u1_n171 ) );
  NAND2_X1 u0_u15_u1_U21 (.ZN( u0_u15_u1_n141 ) , .A1( u0_u15_u1_n153 ) , .A2( u0_u15_u1_n156 ) );
  AND2_X1 u0_u15_u1_U22 (.A1( u0_u15_u1_n123 ) , .ZN( u0_u15_u1_n134 ) , .A2( u0_u15_u1_n161 ) );
  NAND2_X1 u0_u15_u1_U23 (.A2( u0_u15_u1_n115 ) , .A1( u0_u15_u1_n116 ) , .ZN( u0_u15_u1_n148 ) );
  NAND2_X1 u0_u15_u1_U24 (.A2( u0_u15_u1_n133 ) , .A1( u0_u15_u1_n135 ) , .ZN( u0_u15_u1_n159 ) );
  NAND2_X1 u0_u15_u1_U25 (.A2( u0_u15_u1_n115 ) , .A1( u0_u15_u1_n120 ) , .ZN( u0_u15_u1_n132 ) );
  INV_X1 u0_u15_u1_U26 (.A( u0_u15_u1_n154 ) , .ZN( u0_u15_u1_n178 ) );
  INV_X1 u0_u15_u1_U27 (.A( u0_u15_u1_n151 ) , .ZN( u0_u15_u1_n183 ) );
  AND2_X1 u0_u15_u1_U28 (.A1( u0_u15_u1_n129 ) , .A2( u0_u15_u1_n133 ) , .ZN( u0_u15_u1_n149 ) );
  INV_X1 u0_u15_u1_U29 (.A( u0_u15_u1_n131 ) , .ZN( u0_u15_u1_n180 ) );
  INV_X1 u0_u15_u1_U3 (.A( u0_u15_u1_n159 ) , .ZN( u0_u15_u1_n182 ) );
  OAI221_X1 u0_u15_u1_U30 (.A( u0_u15_u1_n119 ) , .C2( u0_u15_u1_n129 ) , .ZN( u0_u15_u1_n138 ) , .B2( u0_u15_u1_n152 ) , .C1( u0_u15_u1_n174 ) , .B1( u0_u15_u1_n187 ) );
  INV_X1 u0_u15_u1_U31 (.A( u0_u15_u1_n148 ) , .ZN( u0_u15_u1_n187 ) );
  AOI211_X1 u0_u15_u1_U32 (.B( u0_u15_u1_n117 ) , .A( u0_u15_u1_n118 ) , .ZN( u0_u15_u1_n119 ) , .C2( u0_u15_u1_n146 ) , .C1( u0_u15_u1_n159 ) );
  NOR2_X1 u0_u15_u1_U33 (.A1( u0_u15_u1_n168 ) , .A2( u0_u15_u1_n176 ) , .ZN( u0_u15_u1_n98 ) );
  AOI211_X1 u0_u15_u1_U34 (.B( u0_u15_u1_n162 ) , .A( u0_u15_u1_n163 ) , .C2( u0_u15_u1_n164 ) , .ZN( u0_u15_u1_n165 ) , .C1( u0_u15_u1_n171 ) );
  AOI21_X1 u0_u15_u1_U35 (.A( u0_u15_u1_n160 ) , .B2( u0_u15_u1_n161 ) , .ZN( u0_u15_u1_n162 ) , .B1( u0_u15_u1_n182 ) );
  OR2_X1 u0_u15_u1_U36 (.A2( u0_u15_u1_n157 ) , .A1( u0_u15_u1_n158 ) , .ZN( u0_u15_u1_n163 ) );
  NAND2_X1 u0_u15_u1_U37 (.A1( u0_u15_u1_n128 ) , .ZN( u0_u15_u1_n146 ) , .A2( u0_u15_u1_n160 ) );
  NAND2_X1 u0_u15_u1_U38 (.A2( u0_u15_u1_n112 ) , .ZN( u0_u15_u1_n139 ) , .A1( u0_u15_u1_n152 ) );
  NAND2_X1 u0_u15_u1_U39 (.A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n156 ) , .A2( u0_u15_u1_n99 ) );
  AOI221_X1 u0_u15_u1_U4 (.A( u0_u15_u1_n138 ) , .C2( u0_u15_u1_n139 ) , .C1( u0_u15_u1_n140 ) , .B2( u0_u15_u1_n141 ) , .ZN( u0_u15_u1_n142 ) , .B1( u0_u15_u1_n175 ) );
  AOI221_X1 u0_u15_u1_U40 (.B1( u0_u15_u1_n140 ) , .ZN( u0_u15_u1_n167 ) , .B2( u0_u15_u1_n172 ) , .C2( u0_u15_u1_n175 ) , .C1( u0_u15_u1_n178 ) , .A( u0_u15_u1_n188 ) );
  INV_X1 u0_u15_u1_U41 (.ZN( u0_u15_u1_n188 ) , .A( u0_u15_u1_n97 ) );
  AOI211_X1 u0_u15_u1_U42 (.A( u0_u15_u1_n118 ) , .C1( u0_u15_u1_n132 ) , .C2( u0_u15_u1_n139 ) , .B( u0_u15_u1_n96 ) , .ZN( u0_u15_u1_n97 ) );
  AOI21_X1 u0_u15_u1_U43 (.B2( u0_u15_u1_n121 ) , .B1( u0_u15_u1_n135 ) , .A( u0_u15_u1_n152 ) , .ZN( u0_u15_u1_n96 ) );
  NOR2_X1 u0_u15_u1_U44 (.ZN( u0_u15_u1_n117 ) , .A1( u0_u15_u1_n121 ) , .A2( u0_u15_u1_n160 ) );
  AOI21_X1 u0_u15_u1_U45 (.A( u0_u15_u1_n128 ) , .B2( u0_u15_u1_n129 ) , .ZN( u0_u15_u1_n130 ) , .B1( u0_u15_u1_n150 ) );
  OAI21_X1 u0_u15_u1_U46 (.B2( u0_u15_u1_n123 ) , .ZN( u0_u15_u1_n145 ) , .B1( u0_u15_u1_n160 ) , .A( u0_u15_u1_n185 ) );
  INV_X1 u0_u15_u1_U47 (.A( u0_u15_u1_n122 ) , .ZN( u0_u15_u1_n185 ) );
  AOI21_X1 u0_u15_u1_U48 (.B2( u0_u15_u1_n120 ) , .B1( u0_u15_u1_n121 ) , .ZN( u0_u15_u1_n122 ) , .A( u0_u15_u1_n128 ) );
  NAND2_X1 u0_u15_u1_U49 (.ZN( u0_u15_u1_n112 ) , .A1( u0_u15_u1_n169 ) , .A2( u0_u15_u1_n170 ) );
  AOI211_X1 u0_u15_u1_U5 (.ZN( u0_u15_u1_n124 ) , .A( u0_u15_u1_n138 ) , .C2( u0_u15_u1_n139 ) , .B( u0_u15_u1_n145 ) , .C1( u0_u15_u1_n147 ) );
  NAND2_X1 u0_u15_u1_U50 (.ZN( u0_u15_u1_n129 ) , .A2( u0_u15_u1_n95 ) , .A1( u0_u15_u1_n98 ) );
  NAND2_X1 u0_u15_u1_U51 (.A1( u0_u15_u1_n102 ) , .ZN( u0_u15_u1_n154 ) , .A2( u0_u15_u1_n99 ) );
  NAND2_X1 u0_u15_u1_U52 (.A2( u0_u15_u1_n100 ) , .ZN( u0_u15_u1_n135 ) , .A1( u0_u15_u1_n99 ) );
  AOI21_X1 u0_u15_u1_U53 (.A( u0_u15_u1_n152 ) , .B2( u0_u15_u1_n153 ) , .B1( u0_u15_u1_n154 ) , .ZN( u0_u15_u1_n158 ) );
  INV_X1 u0_u15_u1_U54 (.A( u0_u15_u1_n160 ) , .ZN( u0_u15_u1_n175 ) );
  NAND2_X1 u0_u15_u1_U55 (.A1( u0_u15_u1_n100 ) , .ZN( u0_u15_u1_n116 ) , .A2( u0_u15_u1_n95 ) );
  NAND2_X1 u0_u15_u1_U56 (.A1( u0_u15_u1_n102 ) , .ZN( u0_u15_u1_n131 ) , .A2( u0_u15_u1_n95 ) );
  NAND2_X1 u0_u15_u1_U57 (.A2( u0_u15_u1_n104 ) , .ZN( u0_u15_u1_n121 ) , .A1( u0_u15_u1_n98 ) );
  NAND2_X1 u0_u15_u1_U58 (.A1( u0_u15_u1_n103 ) , .ZN( u0_u15_u1_n153 ) , .A2( u0_u15_u1_n98 ) );
  NAND2_X1 u0_u15_u1_U59 (.A2( u0_u15_u1_n104 ) , .A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n133 ) );
  AOI22_X1 u0_u15_u1_U6 (.B2( u0_u15_u1_n136 ) , .A2( u0_u15_u1_n137 ) , .ZN( u0_u15_u1_n143 ) , .A1( u0_u15_u1_n171 ) , .B1( u0_u15_u1_n173 ) );
  NAND2_X1 u0_u15_u1_U60 (.ZN( u0_u15_u1_n150 ) , .A2( u0_u15_u1_n98 ) , .A1( u0_u15_u1_n99 ) );
  NAND2_X1 u0_u15_u1_U61 (.A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n155 ) , .A2( u0_u15_u1_n95 ) );
  OAI21_X1 u0_u15_u1_U62 (.ZN( u0_u15_u1_n109 ) , .B1( u0_u15_u1_n129 ) , .B2( u0_u15_u1_n160 ) , .A( u0_u15_u1_n167 ) );
  NAND2_X1 u0_u15_u1_U63 (.A2( u0_u15_u1_n100 ) , .A1( u0_u15_u1_n103 ) , .ZN( u0_u15_u1_n120 ) );
  NAND2_X1 u0_u15_u1_U64 (.A1( u0_u15_u1_n102 ) , .A2( u0_u15_u1_n104 ) , .ZN( u0_u15_u1_n115 ) );
  NAND2_X1 u0_u15_u1_U65 (.A2( u0_u15_u1_n100 ) , .A1( u0_u15_u1_n104 ) , .ZN( u0_u15_u1_n151 ) );
  NAND2_X1 u0_u15_u1_U66 (.A2( u0_u15_u1_n103 ) , .A1( u0_u15_u1_n105 ) , .ZN( u0_u15_u1_n161 ) );
  INV_X1 u0_u15_u1_U67 (.A( u0_u15_u1_n152 ) , .ZN( u0_u15_u1_n173 ) );
  INV_X1 u0_u15_u1_U68 (.A( u0_u15_u1_n128 ) , .ZN( u0_u15_u1_n172 ) );
  NAND2_X1 u0_u15_u1_U69 (.A2( u0_u15_u1_n102 ) , .A1( u0_u15_u1_n103 ) , .ZN( u0_u15_u1_n123 ) );
  INV_X1 u0_u15_u1_U7 (.A( u0_u15_u1_n147 ) , .ZN( u0_u15_u1_n181 ) );
  NOR2_X1 u0_u15_u1_U70 (.A2( u0_u15_X_7 ) , .A1( u0_u15_X_8 ) , .ZN( u0_u15_u1_n95 ) );
  NOR2_X1 u0_u15_u1_U71 (.A1( u0_u15_X_12 ) , .A2( u0_u15_X_9 ) , .ZN( u0_u15_u1_n100 ) );
  NOR2_X1 u0_u15_u1_U72 (.A2( u0_u15_X_8 ) , .A1( u0_u15_u1_n177 ) , .ZN( u0_u15_u1_n99 ) );
  NOR2_X1 u0_u15_u1_U73 (.A2( u0_u15_X_12 ) , .ZN( u0_u15_u1_n102 ) , .A1( u0_u15_u1_n176 ) );
  NOR2_X1 u0_u15_u1_U74 (.A2( u0_u15_X_9 ) , .ZN( u0_u15_u1_n105 ) , .A1( u0_u15_u1_n168 ) );
  NAND2_X1 u0_u15_u1_U75 (.A1( u0_u15_X_10 ) , .ZN( u0_u15_u1_n160 ) , .A2( u0_u15_u1_n169 ) );
  NAND2_X1 u0_u15_u1_U76 (.A2( u0_u15_X_10 ) , .A1( u0_u15_X_11 ) , .ZN( u0_u15_u1_n152 ) );
  NAND2_X1 u0_u15_u1_U77 (.A1( u0_u15_X_11 ) , .ZN( u0_u15_u1_n128 ) , .A2( u0_u15_u1_n170 ) );
  AND2_X1 u0_u15_u1_U78 (.A2( u0_u15_X_7 ) , .A1( u0_u15_X_8 ) , .ZN( u0_u15_u1_n104 ) );
  AND2_X1 u0_u15_u1_U79 (.A1( u0_u15_X_8 ) , .ZN( u0_u15_u1_n103 ) , .A2( u0_u15_u1_n177 ) );
  AOI22_X1 u0_u15_u1_U8 (.B2( u0_u15_u1_n113 ) , .A2( u0_u15_u1_n114 ) , .ZN( u0_u15_u1_n125 ) , .A1( u0_u15_u1_n171 ) , .B1( u0_u15_u1_n173 ) );
  INV_X1 u0_u15_u1_U80 (.A( u0_u15_X_10 ) , .ZN( u0_u15_u1_n170 ) );
  INV_X1 u0_u15_u1_U81 (.A( u0_u15_X_9 ) , .ZN( u0_u15_u1_n176 ) );
  INV_X1 u0_u15_u1_U82 (.A( u0_u15_X_11 ) , .ZN( u0_u15_u1_n169 ) );
  INV_X1 u0_u15_u1_U83 (.A( u0_u15_X_12 ) , .ZN( u0_u15_u1_n168 ) );
  INV_X1 u0_u15_u1_U84 (.A( u0_u15_X_7 ) , .ZN( u0_u15_u1_n177 ) );
  NAND4_X1 u0_u15_u1_U85 (.ZN( u0_out15_18 ) , .A4( u0_u15_u1_n165 ) , .A3( u0_u15_u1_n166 ) , .A1( u0_u15_u1_n167 ) , .A2( u0_u15_u1_n186 ) );
  AOI22_X1 u0_u15_u1_U86 (.B2( u0_u15_u1_n146 ) , .B1( u0_u15_u1_n147 ) , .A2( u0_u15_u1_n148 ) , .ZN( u0_u15_u1_n166 ) , .A1( u0_u15_u1_n172 ) );
  INV_X1 u0_u15_u1_U87 (.A( u0_u15_u1_n145 ) , .ZN( u0_u15_u1_n186 ) );
  NAND4_X1 u0_u15_u1_U88 (.ZN( u0_out15_2 ) , .A4( u0_u15_u1_n142 ) , .A3( u0_u15_u1_n143 ) , .A2( u0_u15_u1_n144 ) , .A1( u0_u15_u1_n179 ) );
  OAI21_X1 u0_u15_u1_U89 (.B2( u0_u15_u1_n132 ) , .ZN( u0_u15_u1_n144 ) , .A( u0_u15_u1_n146 ) , .B1( u0_u15_u1_n180 ) );
  NAND2_X1 u0_u15_u1_U9 (.ZN( u0_u15_u1_n114 ) , .A1( u0_u15_u1_n134 ) , .A2( u0_u15_u1_n156 ) );
  INV_X1 u0_u15_u1_U90 (.A( u0_u15_u1_n130 ) , .ZN( u0_u15_u1_n179 ) );
  NAND4_X1 u0_u15_u1_U91 (.ZN( u0_out15_28 ) , .A4( u0_u15_u1_n124 ) , .A3( u0_u15_u1_n125 ) , .A2( u0_u15_u1_n126 ) , .A1( u0_u15_u1_n127 ) );
  OAI21_X1 u0_u15_u1_U92 (.ZN( u0_u15_u1_n127 ) , .B2( u0_u15_u1_n139 ) , .B1( u0_u15_u1_n175 ) , .A( u0_u15_u1_n183 ) );
  OAI21_X1 u0_u15_u1_U93 (.ZN( u0_u15_u1_n126 ) , .B2( u0_u15_u1_n140 ) , .A( u0_u15_u1_n146 ) , .B1( u0_u15_u1_n178 ) );
  OR4_X1 u0_u15_u1_U94 (.ZN( u0_out15_13 ) , .A4( u0_u15_u1_n108 ) , .A3( u0_u15_u1_n109 ) , .A2( u0_u15_u1_n110 ) , .A1( u0_u15_u1_n111 ) );
  AOI21_X1 u0_u15_u1_U95 (.ZN( u0_u15_u1_n111 ) , .A( u0_u15_u1_n128 ) , .B2( u0_u15_u1_n131 ) , .B1( u0_u15_u1_n135 ) );
  AOI21_X1 u0_u15_u1_U96 (.ZN( u0_u15_u1_n110 ) , .A( u0_u15_u1_n116 ) , .B1( u0_u15_u1_n152 ) , .B2( u0_u15_u1_n160 ) );
  NAND3_X1 u0_u15_u1_U97 (.A3( u0_u15_u1_n149 ) , .A2( u0_u15_u1_n150 ) , .A1( u0_u15_u1_n151 ) , .ZN( u0_u15_u1_n164 ) );
  NAND3_X1 u0_u15_u1_U98 (.A3( u0_u15_u1_n134 ) , .A2( u0_u15_u1_n135 ) , .ZN( u0_u15_u1_n136 ) , .A1( u0_u15_u1_n151 ) );
  NAND3_X1 u0_u15_u1_U99 (.A1( u0_u15_u1_n133 ) , .ZN( u0_u15_u1_n137 ) , .A2( u0_u15_u1_n154 ) , .A3( u0_u15_u1_n181 ) );
  XOR2_X1 u0_u3_U10 (.B( u0_K4_45 ) , .A( u0_R2_30 ) , .Z( u0_u3_X_45 ) );
  XOR2_X1 u0_u3_U11 (.B( u0_K4_44 ) , .A( u0_R2_29 ) , .Z( u0_u3_X_44 ) );
  XOR2_X1 u0_u3_U12 (.B( u0_K4_43 ) , .A( u0_R2_28 ) , .Z( u0_u3_X_43 ) );
  XOR2_X1 u0_u3_U13 (.B( u0_K4_42 ) , .A( u0_R2_29 ) , .Z( u0_u3_X_42 ) );
  XOR2_X1 u0_u3_U14 (.B( u0_K4_41 ) , .A( u0_R2_28 ) , .Z( u0_u3_X_41 ) );
  XOR2_X1 u0_u3_U15 (.B( u0_K4_40 ) , .A( u0_R2_27 ) , .Z( u0_u3_X_40 ) );
  XOR2_X1 u0_u3_U17 (.B( u0_K4_39 ) , .A( u0_R2_26 ) , .Z( u0_u3_X_39 ) );
  XOR2_X1 u0_u3_U18 (.B( u0_K4_38 ) , .A( u0_R2_25 ) , .Z( u0_u3_X_38 ) );
  XOR2_X1 u0_u3_U19 (.B( u0_K4_37 ) , .A( u0_R2_24 ) , .Z( u0_u3_X_37 ) );
  XOR2_X1 u0_u3_U7 (.B( u0_K4_48 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_48 ) );
  XOR2_X1 u0_u3_U8 (.B( u0_K4_47 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_47 ) );
  XOR2_X1 u0_u3_U9 (.B( u0_K4_46 ) , .A( u0_R2_31 ) , .Z( u0_u3_X_46 ) );
  INV_X1 u0_u3_u6_U10 (.ZN( u0_u3_u6_n172 ) , .A( u0_u3_u6_n88 ) );
  OAI21_X1 u0_u3_u6_U11 (.A( u0_u3_u6_n159 ) , .B1( u0_u3_u6_n169 ) , .B2( u0_u3_u6_n173 ) , .ZN( u0_u3_u6_n90 ) );
  AOI22_X1 u0_u3_u6_U12 (.A2( u0_u3_u6_n151 ) , .B2( u0_u3_u6_n161 ) , .A1( u0_u3_u6_n167 ) , .B1( u0_u3_u6_n170 ) , .ZN( u0_u3_u6_n89 ) );
  AOI21_X1 u0_u3_u6_U13 (.ZN( u0_u3_u6_n106 ) , .A( u0_u3_u6_n142 ) , .B2( u0_u3_u6_n159 ) , .B1( u0_u3_u6_n164 ) );
  INV_X1 u0_u3_u6_U14 (.A( u0_u3_u6_n155 ) , .ZN( u0_u3_u6_n161 ) );
  INV_X1 u0_u3_u6_U15 (.A( u0_u3_u6_n128 ) , .ZN( u0_u3_u6_n164 ) );
  NAND2_X1 u0_u3_u6_U16 (.ZN( u0_u3_u6_n110 ) , .A1( u0_u3_u6_n122 ) , .A2( u0_u3_u6_n129 ) );
  NAND2_X1 u0_u3_u6_U17 (.ZN( u0_u3_u6_n124 ) , .A2( u0_u3_u6_n146 ) , .A1( u0_u3_u6_n148 ) );
  INV_X1 u0_u3_u6_U18 (.A( u0_u3_u6_n132 ) , .ZN( u0_u3_u6_n171 ) );
  AND2_X1 u0_u3_u6_U19 (.A1( u0_u3_u6_n100 ) , .ZN( u0_u3_u6_n130 ) , .A2( u0_u3_u6_n147 ) );
  INV_X1 u0_u3_u6_U20 (.A( u0_u3_u6_n127 ) , .ZN( u0_u3_u6_n173 ) );
  INV_X1 u0_u3_u6_U21 (.A( u0_u3_u6_n121 ) , .ZN( u0_u3_u6_n167 ) );
  INV_X1 u0_u3_u6_U22 (.A( u0_u3_u6_n100 ) , .ZN( u0_u3_u6_n169 ) );
  INV_X1 u0_u3_u6_U23 (.A( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n170 ) );
  INV_X1 u0_u3_u6_U24 (.A( u0_u3_u6_n113 ) , .ZN( u0_u3_u6_n168 ) );
  AND2_X1 u0_u3_u6_U25 (.A1( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n119 ) , .ZN( u0_u3_u6_n133 ) );
  AND2_X1 u0_u3_u6_U26 (.A2( u0_u3_u6_n121 ) , .A1( u0_u3_u6_n122 ) , .ZN( u0_u3_u6_n131 ) );
  AND3_X1 u0_u3_u6_U27 (.ZN( u0_u3_u6_n120 ) , .A2( u0_u3_u6_n127 ) , .A1( u0_u3_u6_n132 ) , .A3( u0_u3_u6_n145 ) );
  INV_X1 u0_u3_u6_U28 (.A( u0_u3_u6_n146 ) , .ZN( u0_u3_u6_n163 ) );
  AOI222_X1 u0_u3_u6_U29 (.ZN( u0_u3_u6_n114 ) , .A1( u0_u3_u6_n118 ) , .A2( u0_u3_u6_n126 ) , .B2( u0_u3_u6_n151 ) , .C2( u0_u3_u6_n159 ) , .C1( u0_u3_u6_n168 ) , .B1( u0_u3_u6_n169 ) );
  INV_X1 u0_u3_u6_U3 (.A( u0_u3_u6_n110 ) , .ZN( u0_u3_u6_n166 ) );
  NOR2_X1 u0_u3_u6_U30 (.A1( u0_u3_u6_n162 ) , .A2( u0_u3_u6_n165 ) , .ZN( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U31 (.A1( u0_u3_u6_n144 ) , .ZN( u0_u3_u6_n151 ) , .A2( u0_u3_u6_n158 ) );
  NAND2_X1 u0_u3_u6_U32 (.ZN( u0_u3_u6_n132 ) , .A1( u0_u3_u6_n91 ) , .A2( u0_u3_u6_n97 ) );
  AOI22_X1 u0_u3_u6_U33 (.B2( u0_u3_u6_n110 ) , .B1( u0_u3_u6_n111 ) , .A1( u0_u3_u6_n112 ) , .ZN( u0_u3_u6_n115 ) , .A2( u0_u3_u6_n161 ) );
  NAND4_X1 u0_u3_u6_U34 (.A3( u0_u3_u6_n109 ) , .ZN( u0_u3_u6_n112 ) , .A4( u0_u3_u6_n132 ) , .A2( u0_u3_u6_n147 ) , .A1( u0_u3_u6_n166 ) );
  NOR2_X1 u0_u3_u6_U35 (.ZN( u0_u3_u6_n109 ) , .A1( u0_u3_u6_n170 ) , .A2( u0_u3_u6_n173 ) );
  NOR2_X1 u0_u3_u6_U36 (.A2( u0_u3_u6_n126 ) , .ZN( u0_u3_u6_n155 ) , .A1( u0_u3_u6_n160 ) );
  NAND2_X1 u0_u3_u6_U37 (.ZN( u0_u3_u6_n146 ) , .A2( u0_u3_u6_n94 ) , .A1( u0_u3_u6_n99 ) );
  AOI21_X1 u0_u3_u6_U38 (.A( u0_u3_u6_n144 ) , .B2( u0_u3_u6_n145 ) , .B1( u0_u3_u6_n146 ) , .ZN( u0_u3_u6_n150 ) );
  AOI211_X1 u0_u3_u6_U39 (.B( u0_u3_u6_n134 ) , .A( u0_u3_u6_n135 ) , .C1( u0_u3_u6_n136 ) , .ZN( u0_u3_u6_n137 ) , .C2( u0_u3_u6_n151 ) );
  INV_X1 u0_u3_u6_U4 (.A( u0_u3_u6_n142 ) , .ZN( u0_u3_u6_n174 ) );
  AOI21_X1 u0_u3_u6_U40 (.B2( u0_u3_u6_n132 ) , .B1( u0_u3_u6_n133 ) , .ZN( u0_u3_u6_n134 ) , .A( u0_u3_u6_n158 ) );
  NAND4_X1 u0_u3_u6_U41 (.A4( u0_u3_u6_n127 ) , .A3( u0_u3_u6_n128 ) , .A2( u0_u3_u6_n129 ) , .A1( u0_u3_u6_n130 ) , .ZN( u0_u3_u6_n136 ) );
  AOI21_X1 u0_u3_u6_U42 (.B1( u0_u3_u6_n131 ) , .ZN( u0_u3_u6_n135 ) , .A( u0_u3_u6_n144 ) , .B2( u0_u3_u6_n146 ) );
  INV_X1 u0_u3_u6_U43 (.A( u0_u3_u6_n111 ) , .ZN( u0_u3_u6_n158 ) );
  NAND2_X1 u0_u3_u6_U44 (.ZN( u0_u3_u6_n127 ) , .A1( u0_u3_u6_n91 ) , .A2( u0_u3_u6_n92 ) );
  NAND2_X1 u0_u3_u6_U45 (.ZN( u0_u3_u6_n129 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n96 ) );
  INV_X1 u0_u3_u6_U46 (.A( u0_u3_u6_n144 ) , .ZN( u0_u3_u6_n159 ) );
  NAND2_X1 u0_u3_u6_U47 (.ZN( u0_u3_u6_n145 ) , .A2( u0_u3_u6_n97 ) , .A1( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U48 (.ZN( u0_u3_u6_n148 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n94 ) );
  NAND2_X1 u0_u3_u6_U49 (.ZN( u0_u3_u6_n108 ) , .A2( u0_u3_u6_n139 ) , .A1( u0_u3_u6_n144 ) );
  NAND2_X1 u0_u3_u6_U5 (.A2( u0_u3_u6_n143 ) , .ZN( u0_u3_u6_n152 ) , .A1( u0_u3_u6_n166 ) );
  NAND2_X1 u0_u3_u6_U50 (.ZN( u0_u3_u6_n121 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n97 ) );
  NAND2_X1 u0_u3_u6_U51 (.ZN( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n95 ) );
  AND2_X1 u0_u3_u6_U52 (.ZN( u0_u3_u6_n118 ) , .A2( u0_u3_u6_n91 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U53 (.ZN( u0_u3_u6_n147 ) , .A2( u0_u3_u6_n98 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U54 (.ZN( u0_u3_u6_n128 ) , .A1( u0_u3_u6_n94 ) , .A2( u0_u3_u6_n96 ) );
  NAND2_X1 u0_u3_u6_U55 (.ZN( u0_u3_u6_n119 ) , .A2( u0_u3_u6_n95 ) , .A1( u0_u3_u6_n99 ) );
  NAND2_X1 u0_u3_u6_U56 (.ZN( u0_u3_u6_n123 ) , .A2( u0_u3_u6_n91 ) , .A1( u0_u3_u6_n96 ) );
  NAND2_X1 u0_u3_u6_U57 (.ZN( u0_u3_u6_n100 ) , .A2( u0_u3_u6_n92 ) , .A1( u0_u3_u6_n98 ) );
  NAND2_X1 u0_u3_u6_U58 (.ZN( u0_u3_u6_n122 ) , .A1( u0_u3_u6_n94 ) , .A2( u0_u3_u6_n97 ) );
  INV_X1 u0_u3_u6_U59 (.A( u0_u3_u6_n139 ) , .ZN( u0_u3_u6_n160 ) );
  AOI22_X1 u0_u3_u6_U6 (.B2( u0_u3_u6_n101 ) , .A1( u0_u3_u6_n102 ) , .ZN( u0_u3_u6_n103 ) , .B1( u0_u3_u6_n160 ) , .A2( u0_u3_u6_n161 ) );
  NAND2_X1 u0_u3_u6_U60 (.ZN( u0_u3_u6_n113 ) , .A1( u0_u3_u6_n96 ) , .A2( u0_u3_u6_n98 ) );
  NOR2_X1 u0_u3_u6_U61 (.A2( u0_u3_X_40 ) , .A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n126 ) );
  NOR2_X1 u0_u3_u6_U62 (.A2( u0_u3_X_39 ) , .A1( u0_u3_X_42 ) , .ZN( u0_u3_u6_n92 ) );
  NOR2_X1 u0_u3_u6_U63 (.A2( u0_u3_X_39 ) , .A1( u0_u3_u6_n156 ) , .ZN( u0_u3_u6_n97 ) );
  NOR2_X1 u0_u3_u6_U64 (.A2( u0_u3_X_38 ) , .A1( u0_u3_u6_n165 ) , .ZN( u0_u3_u6_n95 ) );
  NOR2_X1 u0_u3_u6_U65 (.A2( u0_u3_X_41 ) , .ZN( u0_u3_u6_n111 ) , .A1( u0_u3_u6_n157 ) );
  NOR2_X1 u0_u3_u6_U66 (.A2( u0_u3_X_37 ) , .A1( u0_u3_u6_n162 ) , .ZN( u0_u3_u6_n94 ) );
  NOR2_X1 u0_u3_u6_U67 (.A2( u0_u3_X_37 ) , .A1( u0_u3_X_38 ) , .ZN( u0_u3_u6_n91 ) );
  NAND2_X1 u0_u3_u6_U68 (.A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n144 ) , .A2( u0_u3_u6_n157 ) );
  NAND2_X1 u0_u3_u6_U69 (.A2( u0_u3_X_40 ) , .A1( u0_u3_X_41 ) , .ZN( u0_u3_u6_n139 ) );
  NOR2_X1 u0_u3_u6_U7 (.A1( u0_u3_u6_n118 ) , .ZN( u0_u3_u6_n143 ) , .A2( u0_u3_u6_n168 ) );
  AND2_X1 u0_u3_u6_U70 (.A1( u0_u3_X_39 ) , .A2( u0_u3_u6_n156 ) , .ZN( u0_u3_u6_n96 ) );
  AND2_X1 u0_u3_u6_U71 (.A1( u0_u3_X_39 ) , .A2( u0_u3_X_42 ) , .ZN( u0_u3_u6_n99 ) );
  INV_X1 u0_u3_u6_U72 (.A( u0_u3_X_40 ) , .ZN( u0_u3_u6_n157 ) );
  INV_X1 u0_u3_u6_U73 (.A( u0_u3_X_37 ) , .ZN( u0_u3_u6_n165 ) );
  INV_X1 u0_u3_u6_U74 (.A( u0_u3_X_38 ) , .ZN( u0_u3_u6_n162 ) );
  INV_X1 u0_u3_u6_U75 (.A( u0_u3_X_42 ) , .ZN( u0_u3_u6_n156 ) );
  NAND4_X1 u0_u3_u6_U76 (.ZN( u0_out3_32 ) , .A4( u0_u3_u6_n103 ) , .A3( u0_u3_u6_n104 ) , .A2( u0_u3_u6_n105 ) , .A1( u0_u3_u6_n106 ) );
  AOI22_X1 u0_u3_u6_U77 (.ZN( u0_u3_u6_n105 ) , .A2( u0_u3_u6_n108 ) , .A1( u0_u3_u6_n118 ) , .B2( u0_u3_u6_n126 ) , .B1( u0_u3_u6_n171 ) );
  AOI22_X1 u0_u3_u6_U78 (.ZN( u0_u3_u6_n104 ) , .A1( u0_u3_u6_n111 ) , .B1( u0_u3_u6_n124 ) , .B2( u0_u3_u6_n151 ) , .A2( u0_u3_u6_n93 ) );
  NAND4_X1 u0_u3_u6_U79 (.ZN( u0_out3_12 ) , .A4( u0_u3_u6_n114 ) , .A3( u0_u3_u6_n115 ) , .A2( u0_u3_u6_n116 ) , .A1( u0_u3_u6_n117 ) );
  AOI21_X1 u0_u3_u6_U8 (.B1( u0_u3_u6_n107 ) , .B2( u0_u3_u6_n132 ) , .A( u0_u3_u6_n158 ) , .ZN( u0_u3_u6_n88 ) );
  OAI22_X1 u0_u3_u6_U80 (.B2( u0_u3_u6_n111 ) , .ZN( u0_u3_u6_n116 ) , .B1( u0_u3_u6_n126 ) , .A2( u0_u3_u6_n164 ) , .A1( u0_u3_u6_n167 ) );
  OAI21_X1 u0_u3_u6_U81 (.A( u0_u3_u6_n108 ) , .ZN( u0_u3_u6_n117 ) , .B2( u0_u3_u6_n141 ) , .B1( u0_u3_u6_n163 ) );
  OAI211_X1 u0_u3_u6_U82 (.ZN( u0_out3_22 ) , .B( u0_u3_u6_n137 ) , .A( u0_u3_u6_n138 ) , .C2( u0_u3_u6_n139 ) , .C1( u0_u3_u6_n140 ) );
  AOI22_X1 u0_u3_u6_U83 (.B1( u0_u3_u6_n124 ) , .A2( u0_u3_u6_n125 ) , .A1( u0_u3_u6_n126 ) , .ZN( u0_u3_u6_n138 ) , .B2( u0_u3_u6_n161 ) );
  AND4_X1 u0_u3_u6_U84 (.A3( u0_u3_u6_n119 ) , .A1( u0_u3_u6_n120 ) , .A4( u0_u3_u6_n129 ) , .ZN( u0_u3_u6_n140 ) , .A2( u0_u3_u6_n143 ) );
  OAI211_X1 u0_u3_u6_U85 (.ZN( u0_out3_7 ) , .B( u0_u3_u6_n153 ) , .C2( u0_u3_u6_n154 ) , .C1( u0_u3_u6_n155 ) , .A( u0_u3_u6_n174 ) );
  NOR3_X1 u0_u3_u6_U86 (.A1( u0_u3_u6_n141 ) , .ZN( u0_u3_u6_n154 ) , .A3( u0_u3_u6_n164 ) , .A2( u0_u3_u6_n171 ) );
  AOI211_X1 u0_u3_u6_U87 (.B( u0_u3_u6_n149 ) , .A( u0_u3_u6_n150 ) , .C2( u0_u3_u6_n151 ) , .C1( u0_u3_u6_n152 ) , .ZN( u0_u3_u6_n153 ) );
  NAND3_X1 u0_u3_u6_U88 (.A2( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n125 ) , .A1( u0_u3_u6_n130 ) , .A3( u0_u3_u6_n131 ) );
  NAND3_X1 u0_u3_u6_U89 (.A3( u0_u3_u6_n133 ) , .ZN( u0_u3_u6_n141 ) , .A1( u0_u3_u6_n145 ) , .A2( u0_u3_u6_n148 ) );
  AOI21_X1 u0_u3_u6_U9 (.B2( u0_u3_u6_n147 ) , .B1( u0_u3_u6_n148 ) , .ZN( u0_u3_u6_n149 ) , .A( u0_u3_u6_n158 ) );
  NAND3_X1 u0_u3_u6_U90 (.ZN( u0_u3_u6_n101 ) , .A3( u0_u3_u6_n107 ) , .A2( u0_u3_u6_n121 ) , .A1( u0_u3_u6_n127 ) );
  NAND3_X1 u0_u3_u6_U91 (.ZN( u0_u3_u6_n102 ) , .A3( u0_u3_u6_n130 ) , .A2( u0_u3_u6_n145 ) , .A1( u0_u3_u6_n166 ) );
  NAND3_X1 u0_u3_u6_U92 (.A3( u0_u3_u6_n113 ) , .A1( u0_u3_u6_n119 ) , .A2( u0_u3_u6_n123 ) , .ZN( u0_u3_u6_n93 ) );
  NAND3_X1 u0_u3_u6_U93 (.ZN( u0_u3_u6_n142 ) , .A2( u0_u3_u6_n172 ) , .A3( u0_u3_u6_n89 ) , .A1( u0_u3_u6_n90 ) );
  AND3_X1 u0_u3_u7_U10 (.A3( u0_u3_u7_n110 ) , .A2( u0_u3_u7_n127 ) , .A1( u0_u3_u7_n132 ) , .ZN( u0_u3_u7_n92 ) );
  OAI21_X1 u0_u3_u7_U11 (.A( u0_u3_u7_n161 ) , .B1( u0_u3_u7_n168 ) , .B2( u0_u3_u7_n173 ) , .ZN( u0_u3_u7_n91 ) );
  AOI211_X1 u0_u3_u7_U12 (.A( u0_u3_u7_n117 ) , .ZN( u0_u3_u7_n118 ) , .C2( u0_u3_u7_n126 ) , .C1( u0_u3_u7_n177 ) , .B( u0_u3_u7_n180 ) );
  OAI22_X1 u0_u3_u7_U13 (.B1( u0_u3_u7_n115 ) , .ZN( u0_u3_u7_n117 ) , .A2( u0_u3_u7_n133 ) , .A1( u0_u3_u7_n137 ) , .B2( u0_u3_u7_n162 ) );
  INV_X1 u0_u3_u7_U14 (.A( u0_u3_u7_n116 ) , .ZN( u0_u3_u7_n180 ) );
  NOR3_X1 u0_u3_u7_U15 (.ZN( u0_u3_u7_n115 ) , .A3( u0_u3_u7_n145 ) , .A2( u0_u3_u7_n168 ) , .A1( u0_u3_u7_n169 ) );
  OAI211_X1 u0_u3_u7_U16 (.B( u0_u3_u7_n122 ) , .A( u0_u3_u7_n123 ) , .C2( u0_u3_u7_n124 ) , .ZN( u0_u3_u7_n154 ) , .C1( u0_u3_u7_n162 ) );
  AOI222_X1 u0_u3_u7_U17 (.ZN( u0_u3_u7_n122 ) , .C2( u0_u3_u7_n126 ) , .C1( u0_u3_u7_n145 ) , .B1( u0_u3_u7_n161 ) , .A2( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n170 ) , .A1( u0_u3_u7_n176 ) );
  INV_X1 u0_u3_u7_U18 (.A( u0_u3_u7_n133 ) , .ZN( u0_u3_u7_n176 ) );
  NOR3_X1 u0_u3_u7_U19 (.A2( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n135 ) , .ZN( u0_u3_u7_n136 ) , .A3( u0_u3_u7_n171 ) );
  NOR2_X1 u0_u3_u7_U20 (.A1( u0_u3_u7_n130 ) , .A2( u0_u3_u7_n134 ) , .ZN( u0_u3_u7_n153 ) );
  INV_X1 u0_u3_u7_U21 (.A( u0_u3_u7_n101 ) , .ZN( u0_u3_u7_n165 ) );
  NOR2_X1 u0_u3_u7_U22 (.ZN( u0_u3_u7_n111 ) , .A2( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n169 ) );
  AOI21_X1 u0_u3_u7_U23 (.ZN( u0_u3_u7_n104 ) , .B2( u0_u3_u7_n112 ) , .B1( u0_u3_u7_n127 ) , .A( u0_u3_u7_n164 ) );
  AOI21_X1 u0_u3_u7_U24 (.ZN( u0_u3_u7_n106 ) , .B1( u0_u3_u7_n133 ) , .B2( u0_u3_u7_n146 ) , .A( u0_u3_u7_n162 ) );
  AOI21_X1 u0_u3_u7_U25 (.A( u0_u3_u7_n101 ) , .ZN( u0_u3_u7_n107 ) , .B2( u0_u3_u7_n128 ) , .B1( u0_u3_u7_n175 ) );
  INV_X1 u0_u3_u7_U26 (.A( u0_u3_u7_n138 ) , .ZN( u0_u3_u7_n171 ) );
  INV_X1 u0_u3_u7_U27 (.A( u0_u3_u7_n131 ) , .ZN( u0_u3_u7_n177 ) );
  INV_X1 u0_u3_u7_U28 (.A( u0_u3_u7_n110 ) , .ZN( u0_u3_u7_n174 ) );
  NAND2_X1 u0_u3_u7_U29 (.A1( u0_u3_u7_n129 ) , .A2( u0_u3_u7_n132 ) , .ZN( u0_u3_u7_n149 ) );
  OAI21_X1 u0_u3_u7_U3 (.ZN( u0_u3_u7_n159 ) , .A( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n171 ) , .B1( u0_u3_u7_n174 ) );
  NAND2_X1 u0_u3_u7_U30 (.A1( u0_u3_u7_n113 ) , .A2( u0_u3_u7_n124 ) , .ZN( u0_u3_u7_n130 ) );
  INV_X1 u0_u3_u7_U31 (.A( u0_u3_u7_n112 ) , .ZN( u0_u3_u7_n173 ) );
  INV_X1 u0_u3_u7_U32 (.A( u0_u3_u7_n128 ) , .ZN( u0_u3_u7_n168 ) );
  INV_X1 u0_u3_u7_U33 (.A( u0_u3_u7_n148 ) , .ZN( u0_u3_u7_n169 ) );
  INV_X1 u0_u3_u7_U34 (.A( u0_u3_u7_n127 ) , .ZN( u0_u3_u7_n179 ) );
  NOR2_X1 u0_u3_u7_U35 (.ZN( u0_u3_u7_n101 ) , .A2( u0_u3_u7_n150 ) , .A1( u0_u3_u7_n156 ) );
  AOI211_X1 u0_u3_u7_U36 (.B( u0_u3_u7_n154 ) , .A( u0_u3_u7_n155 ) , .C1( u0_u3_u7_n156 ) , .ZN( u0_u3_u7_n157 ) , .C2( u0_u3_u7_n172 ) );
  INV_X1 u0_u3_u7_U37 (.A( u0_u3_u7_n153 ) , .ZN( u0_u3_u7_n172 ) );
  AOI211_X1 u0_u3_u7_U38 (.B( u0_u3_u7_n139 ) , .A( u0_u3_u7_n140 ) , .C2( u0_u3_u7_n141 ) , .ZN( u0_u3_u7_n142 ) , .C1( u0_u3_u7_n156 ) );
  NAND4_X1 u0_u3_u7_U39 (.A3( u0_u3_u7_n127 ) , .A2( u0_u3_u7_n128 ) , .A1( u0_u3_u7_n129 ) , .ZN( u0_u3_u7_n141 ) , .A4( u0_u3_u7_n147 ) );
  INV_X1 u0_u3_u7_U4 (.A( u0_u3_u7_n111 ) , .ZN( u0_u3_u7_n170 ) );
  AOI21_X1 u0_u3_u7_U40 (.A( u0_u3_u7_n137 ) , .B1( u0_u3_u7_n138 ) , .ZN( u0_u3_u7_n139 ) , .B2( u0_u3_u7_n146 ) );
  OAI22_X1 u0_u3_u7_U41 (.B1( u0_u3_u7_n136 ) , .ZN( u0_u3_u7_n140 ) , .A1( u0_u3_u7_n153 ) , .B2( u0_u3_u7_n162 ) , .A2( u0_u3_u7_n164 ) );
  AOI21_X1 u0_u3_u7_U42 (.ZN( u0_u3_u7_n123 ) , .B1( u0_u3_u7_n165 ) , .B2( u0_u3_u7_n177 ) , .A( u0_u3_u7_n97 ) );
  AOI21_X1 u0_u3_u7_U43 (.B2( u0_u3_u7_n113 ) , .B1( u0_u3_u7_n124 ) , .A( u0_u3_u7_n125 ) , .ZN( u0_u3_u7_n97 ) );
  INV_X1 u0_u3_u7_U44 (.A( u0_u3_u7_n125 ) , .ZN( u0_u3_u7_n161 ) );
  INV_X1 u0_u3_u7_U45 (.A( u0_u3_u7_n152 ) , .ZN( u0_u3_u7_n162 ) );
  AOI22_X1 u0_u3_u7_U46 (.A2( u0_u3_u7_n114 ) , .ZN( u0_u3_u7_n119 ) , .B1( u0_u3_u7_n130 ) , .A1( u0_u3_u7_n156 ) , .B2( u0_u3_u7_n165 ) );
  NAND2_X1 u0_u3_u7_U47 (.A2( u0_u3_u7_n112 ) , .ZN( u0_u3_u7_n114 ) , .A1( u0_u3_u7_n175 ) );
  AND2_X1 u0_u3_u7_U48 (.ZN( u0_u3_u7_n145 ) , .A2( u0_u3_u7_n98 ) , .A1( u0_u3_u7_n99 ) );
  NOR2_X1 u0_u3_u7_U49 (.ZN( u0_u3_u7_n137 ) , .A1( u0_u3_u7_n150 ) , .A2( u0_u3_u7_n161 ) );
  INV_X1 u0_u3_u7_U5 (.A( u0_u3_u7_n149 ) , .ZN( u0_u3_u7_n175 ) );
  AOI21_X1 u0_u3_u7_U50 (.ZN( u0_u3_u7_n105 ) , .B2( u0_u3_u7_n110 ) , .A( u0_u3_u7_n125 ) , .B1( u0_u3_u7_n147 ) );
  NAND2_X1 u0_u3_u7_U51 (.ZN( u0_u3_u7_n146 ) , .A1( u0_u3_u7_n95 ) , .A2( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U52 (.A2( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n147 ) , .A1( u0_u3_u7_n93 ) );
  NAND2_X1 u0_u3_u7_U53 (.A1( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n127 ) , .A2( u0_u3_u7_n99 ) );
  OR2_X1 u0_u3_u7_U54 (.ZN( u0_u3_u7_n126 ) , .A2( u0_u3_u7_n152 ) , .A1( u0_u3_u7_n156 ) );
  NAND2_X1 u0_u3_u7_U55 (.A2( u0_u3_u7_n102 ) , .A1( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n133 ) );
  NAND2_X1 u0_u3_u7_U56 (.ZN( u0_u3_u7_n112 ) , .A2( u0_u3_u7_n96 ) , .A1( u0_u3_u7_n99 ) );
  NAND2_X1 u0_u3_u7_U57 (.A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n128 ) , .A1( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U58 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n113 ) , .A2( u0_u3_u7_n93 ) );
  NAND2_X1 u0_u3_u7_U59 (.A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n124 ) , .A1( u0_u3_u7_n96 ) );
  INV_X1 u0_u3_u7_U6 (.A( u0_u3_u7_n154 ) , .ZN( u0_u3_u7_n178 ) );
  NAND2_X1 u0_u3_u7_U60 (.ZN( u0_u3_u7_n110 ) , .A1( u0_u3_u7_n95 ) , .A2( u0_u3_u7_n96 ) );
  INV_X1 u0_u3_u7_U61 (.A( u0_u3_u7_n150 ) , .ZN( u0_u3_u7_n164 ) );
  AND2_X1 u0_u3_u7_U62 (.ZN( u0_u3_u7_n134 ) , .A1( u0_u3_u7_n93 ) , .A2( u0_u3_u7_n98 ) );
  NAND2_X1 u0_u3_u7_U63 (.A1( u0_u3_u7_n100 ) , .A2( u0_u3_u7_n102 ) , .ZN( u0_u3_u7_n129 ) );
  NAND2_X1 u0_u3_u7_U64 (.A2( u0_u3_u7_n103 ) , .ZN( u0_u3_u7_n131 ) , .A1( u0_u3_u7_n95 ) );
  NAND2_X1 u0_u3_u7_U65 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n138 ) , .A2( u0_u3_u7_n99 ) );
  NAND2_X1 u0_u3_u7_U66 (.ZN( u0_u3_u7_n132 ) , .A1( u0_u3_u7_n93 ) , .A2( u0_u3_u7_n96 ) );
  NAND2_X1 u0_u3_u7_U67 (.A1( u0_u3_u7_n100 ) , .ZN( u0_u3_u7_n148 ) , .A2( u0_u3_u7_n95 ) );
  NOR2_X1 u0_u3_u7_U68 (.A2( u0_u3_X_47 ) , .ZN( u0_u3_u7_n150 ) , .A1( u0_u3_u7_n163 ) );
  NOR2_X1 u0_u3_u7_U69 (.A2( u0_u3_X_43 ) , .A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n103 ) );
  AOI211_X1 u0_u3_u7_U7 (.ZN( u0_u3_u7_n116 ) , .A( u0_u3_u7_n155 ) , .C1( u0_u3_u7_n161 ) , .C2( u0_u3_u7_n171 ) , .B( u0_u3_u7_n94 ) );
  NOR2_X1 u0_u3_u7_U70 (.A2( u0_u3_X_48 ) , .A1( u0_u3_u7_n166 ) , .ZN( u0_u3_u7_n95 ) );
  NOR2_X1 u0_u3_u7_U71 (.A2( u0_u3_X_45 ) , .A1( u0_u3_X_48 ) , .ZN( u0_u3_u7_n99 ) );
  NOR2_X1 u0_u3_u7_U72 (.A2( u0_u3_X_44 ) , .A1( u0_u3_u7_n167 ) , .ZN( u0_u3_u7_n98 ) );
  NOR2_X1 u0_u3_u7_U73 (.A2( u0_u3_X_46 ) , .A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n152 ) );
  AND2_X1 u0_u3_u7_U74 (.A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n156 ) , .A2( u0_u3_u7_n163 ) );
  NAND2_X1 u0_u3_u7_U75 (.A2( u0_u3_X_46 ) , .A1( u0_u3_X_47 ) , .ZN( u0_u3_u7_n125 ) );
  AND2_X1 u0_u3_u7_U76 (.A2( u0_u3_X_45 ) , .A1( u0_u3_X_48 ) , .ZN( u0_u3_u7_n102 ) );
  AND2_X1 u0_u3_u7_U77 (.A2( u0_u3_X_43 ) , .A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n96 ) );
  AND2_X1 u0_u3_u7_U78 (.A1( u0_u3_X_44 ) , .ZN( u0_u3_u7_n100 ) , .A2( u0_u3_u7_n167 ) );
  AND2_X1 u0_u3_u7_U79 (.A1( u0_u3_X_48 ) , .A2( u0_u3_u7_n166 ) , .ZN( u0_u3_u7_n93 ) );
  OAI222_X1 u0_u3_u7_U8 (.C2( u0_u3_u7_n101 ) , .B2( u0_u3_u7_n111 ) , .A1( u0_u3_u7_n113 ) , .C1( u0_u3_u7_n146 ) , .A2( u0_u3_u7_n162 ) , .B1( u0_u3_u7_n164 ) , .ZN( u0_u3_u7_n94 ) );
  INV_X1 u0_u3_u7_U80 (.A( u0_u3_X_46 ) , .ZN( u0_u3_u7_n163 ) );
  INV_X1 u0_u3_u7_U81 (.A( u0_u3_X_43 ) , .ZN( u0_u3_u7_n167 ) );
  INV_X1 u0_u3_u7_U82 (.A( u0_u3_X_45 ) , .ZN( u0_u3_u7_n166 ) );
  NAND4_X1 u0_u3_u7_U83 (.ZN( u0_out3_5 ) , .A4( u0_u3_u7_n108 ) , .A3( u0_u3_u7_n109 ) , .A1( u0_u3_u7_n116 ) , .A2( u0_u3_u7_n123 ) );
  AOI22_X1 u0_u3_u7_U84 (.ZN( u0_u3_u7_n109 ) , .A2( u0_u3_u7_n126 ) , .B2( u0_u3_u7_n145 ) , .B1( u0_u3_u7_n156 ) , .A1( u0_u3_u7_n171 ) );
  NOR4_X1 u0_u3_u7_U85 (.A4( u0_u3_u7_n104 ) , .A3( u0_u3_u7_n105 ) , .A2( u0_u3_u7_n106 ) , .A1( u0_u3_u7_n107 ) , .ZN( u0_u3_u7_n108 ) );
  NAND4_X1 u0_u3_u7_U86 (.ZN( u0_out3_27 ) , .A4( u0_u3_u7_n118 ) , .A3( u0_u3_u7_n119 ) , .A2( u0_u3_u7_n120 ) , .A1( u0_u3_u7_n121 ) );
  OAI21_X1 u0_u3_u7_U87 (.ZN( u0_u3_u7_n121 ) , .B2( u0_u3_u7_n145 ) , .A( u0_u3_u7_n150 ) , .B1( u0_u3_u7_n174 ) );
  OAI21_X1 u0_u3_u7_U88 (.ZN( u0_u3_u7_n120 ) , .A( u0_u3_u7_n161 ) , .B2( u0_u3_u7_n170 ) , .B1( u0_u3_u7_n179 ) );
  NAND4_X1 u0_u3_u7_U89 (.ZN( u0_out3_21 ) , .A4( u0_u3_u7_n157 ) , .A3( u0_u3_u7_n158 ) , .A2( u0_u3_u7_n159 ) , .A1( u0_u3_u7_n160 ) );
  OAI221_X1 u0_u3_u7_U9 (.C1( u0_u3_u7_n101 ) , .C2( u0_u3_u7_n147 ) , .ZN( u0_u3_u7_n155 ) , .B2( u0_u3_u7_n162 ) , .A( u0_u3_u7_n91 ) , .B1( u0_u3_u7_n92 ) );
  OAI21_X1 u0_u3_u7_U90 (.B1( u0_u3_u7_n145 ) , .ZN( u0_u3_u7_n160 ) , .A( u0_u3_u7_n161 ) , .B2( u0_u3_u7_n177 ) );
  AOI22_X1 u0_u3_u7_U91 (.B2( u0_u3_u7_n149 ) , .B1( u0_u3_u7_n150 ) , .A2( u0_u3_u7_n151 ) , .A1( u0_u3_u7_n152 ) , .ZN( u0_u3_u7_n158 ) );
  NAND4_X1 u0_u3_u7_U92 (.ZN( u0_out3_15 ) , .A4( u0_u3_u7_n142 ) , .A3( u0_u3_u7_n143 ) , .A2( u0_u3_u7_n144 ) , .A1( u0_u3_u7_n178 ) );
  OR2_X1 u0_u3_u7_U93 (.A2( u0_u3_u7_n125 ) , .A1( u0_u3_u7_n129 ) , .ZN( u0_u3_u7_n144 ) );
  AOI22_X1 u0_u3_u7_U94 (.A2( u0_u3_u7_n126 ) , .ZN( u0_u3_u7_n143 ) , .B2( u0_u3_u7_n165 ) , .B1( u0_u3_u7_n173 ) , .A1( u0_u3_u7_n174 ) );
  NAND3_X1 u0_u3_u7_U95 (.A3( u0_u3_u7_n146 ) , .A2( u0_u3_u7_n147 ) , .A1( u0_u3_u7_n148 ) , .ZN( u0_u3_u7_n151 ) );
  NAND3_X1 u0_u3_u7_U96 (.A3( u0_u3_u7_n131 ) , .A2( u0_u3_u7_n132 ) , .A1( u0_u3_u7_n133 ) , .ZN( u0_u3_u7_n135 ) );
  XOR2_X1 u0_u5_U1 (.B( u0_K6_9 ) , .A( u0_R4_6 ) , .Z( u0_u5_X_9 ) );
  XOR2_X1 u0_u5_U16 (.B( u0_K6_3 ) , .A( u0_R4_2 ) , .Z( u0_u5_X_3 ) );
  XOR2_X1 u0_u5_U2 (.B( u0_K6_8 ) , .A( u0_R4_5 ) , .Z( u0_u5_X_8 ) );
  XOR2_X1 u0_u5_U27 (.B( u0_K6_2 ) , .A( u0_R4_1 ) , .Z( u0_u5_X_2 ) );
  XOR2_X1 u0_u5_U3 (.B( u0_K6_7 ) , .A( u0_R4_4 ) , .Z( u0_u5_X_7 ) );
  XOR2_X1 u0_u5_U38 (.B( u0_K6_1 ) , .A( u0_R4_32 ) , .Z( u0_u5_X_1 ) );
  XOR2_X1 u0_u5_U4 (.B( u0_K6_6 ) , .A( u0_R4_5 ) , .Z( u0_u5_X_6 ) );
  XOR2_X1 u0_u5_U40 (.B( u0_K6_18 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_18 ) );
  XOR2_X1 u0_u5_U41 (.B( u0_K6_17 ) , .A( u0_R4_12 ) , .Z( u0_u5_X_17 ) );
  XOR2_X1 u0_u5_U42 (.B( u0_K6_16 ) , .A( u0_R4_11 ) , .Z( u0_u5_X_16 ) );
  XOR2_X1 u0_u5_U43 (.B( u0_K6_15 ) , .A( u0_R4_10 ) , .Z( u0_u5_X_15 ) );
  XOR2_X1 u0_u5_U44 (.B( u0_K6_14 ) , .A( u0_R4_9 ) , .Z( u0_u5_X_14 ) );
  XOR2_X1 u0_u5_U45 (.B( u0_K6_13 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_13 ) );
  XOR2_X1 u0_u5_U46 (.B( u0_K6_12 ) , .A( u0_R4_9 ) , .Z( u0_u5_X_12 ) );
  XOR2_X1 u0_u5_U47 (.B( u0_K6_11 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_11 ) );
  XOR2_X1 u0_u5_U48 (.B( u0_K6_10 ) , .A( u0_R4_7 ) , .Z( u0_u5_X_10 ) );
  XOR2_X1 u0_u5_U5 (.B( u0_K6_5 ) , .A( u0_R4_4 ) , .Z( u0_u5_X_5 ) );
  XOR2_X1 u0_u5_U6 (.B( u0_K6_4 ) , .A( u0_R4_3 ) , .Z( u0_u5_X_4 ) );
  AND2_X1 u0_u5_u0_U10 (.A1( u0_u5_u0_n131 ) , .ZN( u0_u5_u0_n141 ) , .A2( u0_u5_u0_n150 ) );
  AND3_X1 u0_u5_u0_U11 (.A2( u0_u5_u0_n112 ) , .ZN( u0_u5_u0_n127 ) , .A3( u0_u5_u0_n130 ) , .A1( u0_u5_u0_n148 ) );
  AND2_X1 u0_u5_u0_U12 (.ZN( u0_u5_u0_n107 ) , .A1( u0_u5_u0_n130 ) , .A2( u0_u5_u0_n140 ) );
  AND2_X1 u0_u5_u0_U13 (.A2( u0_u5_u0_n129 ) , .A1( u0_u5_u0_n130 ) , .ZN( u0_u5_u0_n151 ) );
  AND2_X1 u0_u5_u0_U14 (.A1( u0_u5_u0_n108 ) , .A2( u0_u5_u0_n125 ) , .ZN( u0_u5_u0_n145 ) );
  INV_X1 u0_u5_u0_U15 (.A( u0_u5_u0_n143 ) , .ZN( u0_u5_u0_n173 ) );
  NOR2_X1 u0_u5_u0_U16 (.A2( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n147 ) , .A1( u0_u5_u0_n160 ) );
  AOI21_X1 u0_u5_u0_U17 (.B1( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n132 ) , .A( u0_u5_u0_n165 ) , .B2( u0_u5_u0_n93 ) );
  OAI22_X1 u0_u5_u0_U18 (.B1( u0_u5_u0_n131 ) , .A1( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n147 ) , .A2( u0_u5_u0_n90 ) , .ZN( u0_u5_u0_n91 ) );
  AND3_X1 u0_u5_u0_U19 (.A3( u0_u5_u0_n121 ) , .A2( u0_u5_u0_n125 ) , .A1( u0_u5_u0_n148 ) , .ZN( u0_u5_u0_n90 ) );
  OAI22_X1 u0_u5_u0_U20 (.B1( u0_u5_u0_n125 ) , .ZN( u0_u5_u0_n126 ) , .A1( u0_u5_u0_n138 ) , .A2( u0_u5_u0_n146 ) , .B2( u0_u5_u0_n147 ) );
  NOR2_X1 u0_u5_u0_U21 (.A1( u0_u5_u0_n163 ) , .A2( u0_u5_u0_n164 ) , .ZN( u0_u5_u0_n95 ) );
  AOI22_X1 u0_u5_u0_U22 (.B2( u0_u5_u0_n109 ) , .A2( u0_u5_u0_n110 ) , .ZN( u0_u5_u0_n111 ) , .B1( u0_u5_u0_n118 ) , .A1( u0_u5_u0_n160 ) );
  NAND2_X1 u0_u5_u0_U23 (.A2( u0_u5_u0_n102 ) , .A1( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n149 ) );
  INV_X1 u0_u5_u0_U24 (.A( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n161 ) );
  INV_X1 u0_u5_u0_U25 (.A( u0_u5_u0_n118 ) , .ZN( u0_u5_u0_n158 ) );
  NAND2_X1 u0_u5_u0_U26 (.A2( u0_u5_u0_n100 ) , .ZN( u0_u5_u0_n131 ) , .A1( u0_u5_u0_n92 ) );
  NAND2_X1 u0_u5_u0_U27 (.ZN( u0_u5_u0_n108 ) , .A1( u0_u5_u0_n92 ) , .A2( u0_u5_u0_n94 ) );
  AOI21_X1 u0_u5_u0_U28 (.ZN( u0_u5_u0_n104 ) , .B1( u0_u5_u0_n107 ) , .B2( u0_u5_u0_n141 ) , .A( u0_u5_u0_n144 ) );
  AOI21_X1 u0_u5_u0_U29 (.B1( u0_u5_u0_n127 ) , .B2( u0_u5_u0_n129 ) , .A( u0_u5_u0_n138 ) , .ZN( u0_u5_u0_n96 ) );
  INV_X1 u0_u5_u0_U3 (.A( u0_u5_u0_n113 ) , .ZN( u0_u5_u0_n166 ) );
  NAND2_X1 u0_u5_u0_U30 (.A2( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n114 ) , .A1( u0_u5_u0_n92 ) );
  NOR2_X1 u0_u5_u0_U31 (.A1( u0_u5_u0_n120 ) , .ZN( u0_u5_u0_n143 ) , .A2( u0_u5_u0_n167 ) );
  OAI221_X1 u0_u5_u0_U32 (.C1( u0_u5_u0_n112 ) , .ZN( u0_u5_u0_n120 ) , .B1( u0_u5_u0_n138 ) , .B2( u0_u5_u0_n141 ) , .C2( u0_u5_u0_n147 ) , .A( u0_u5_u0_n172 ) );
  AOI211_X1 u0_u5_u0_U33 (.B( u0_u5_u0_n115 ) , .A( u0_u5_u0_n116 ) , .C2( u0_u5_u0_n117 ) , .C1( u0_u5_u0_n118 ) , .ZN( u0_u5_u0_n119 ) );
  NAND2_X1 u0_u5_u0_U34 (.A2( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n140 ) , .A1( u0_u5_u0_n94 ) );
  NAND2_X1 u0_u5_u0_U35 (.A1( u0_u5_u0_n100 ) , .A2( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n125 ) );
  NAND2_X1 u0_u5_u0_U36 (.A1( u0_u5_u0_n101 ) , .A2( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n150 ) );
  INV_X1 u0_u5_u0_U37 (.A( u0_u5_u0_n138 ) , .ZN( u0_u5_u0_n160 ) );
  NAND2_X1 u0_u5_u0_U38 (.A2( u0_u5_u0_n100 ) , .A1( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n139 ) );
  NAND2_X1 u0_u5_u0_U39 (.ZN( u0_u5_u0_n112 ) , .A2( u0_u5_u0_n92 ) , .A1( u0_u5_u0_n93 ) );
  AOI21_X1 u0_u5_u0_U4 (.B1( u0_u5_u0_n114 ) , .ZN( u0_u5_u0_n115 ) , .B2( u0_u5_u0_n129 ) , .A( u0_u5_u0_n161 ) );
  NAND2_X1 u0_u5_u0_U40 (.A1( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n130 ) , .A2( u0_u5_u0_n94 ) );
  INV_X1 u0_u5_u0_U41 (.ZN( u0_u5_u0_n172 ) , .A( u0_u5_u0_n88 ) );
  OAI222_X1 u0_u5_u0_U42 (.C1( u0_u5_u0_n108 ) , .A1( u0_u5_u0_n125 ) , .B2( u0_u5_u0_n128 ) , .B1( u0_u5_u0_n144 ) , .A2( u0_u5_u0_n158 ) , .C2( u0_u5_u0_n161 ) , .ZN( u0_u5_u0_n88 ) );
  NAND2_X1 u0_u5_u0_U43 (.A2( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n121 ) , .A1( u0_u5_u0_n93 ) );
  OR3_X1 u0_u5_u0_U44 (.A3( u0_u5_u0_n152 ) , .A2( u0_u5_u0_n153 ) , .A1( u0_u5_u0_n154 ) , .ZN( u0_u5_u0_n155 ) );
  AOI21_X1 u0_u5_u0_U45 (.A( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n145 ) , .B1( u0_u5_u0_n146 ) , .ZN( u0_u5_u0_n154 ) );
  AOI21_X1 u0_u5_u0_U46 (.B2( u0_u5_u0_n150 ) , .B1( u0_u5_u0_n151 ) , .ZN( u0_u5_u0_n152 ) , .A( u0_u5_u0_n158 ) );
  AOI21_X1 u0_u5_u0_U47 (.A( u0_u5_u0_n147 ) , .B2( u0_u5_u0_n148 ) , .B1( u0_u5_u0_n149 ) , .ZN( u0_u5_u0_n153 ) );
  INV_X1 u0_u5_u0_U48 (.ZN( u0_u5_u0_n171 ) , .A( u0_u5_u0_n99 ) );
  OAI211_X1 u0_u5_u0_U49 (.C2( u0_u5_u0_n140 ) , .C1( u0_u5_u0_n161 ) , .A( u0_u5_u0_n169 ) , .B( u0_u5_u0_n98 ) , .ZN( u0_u5_u0_n99 ) );
  AOI21_X1 u0_u5_u0_U5 (.B2( u0_u5_u0_n131 ) , .ZN( u0_u5_u0_n134 ) , .B1( u0_u5_u0_n151 ) , .A( u0_u5_u0_n158 ) );
  AOI211_X1 u0_u5_u0_U50 (.C1( u0_u5_u0_n118 ) , .A( u0_u5_u0_n123 ) , .B( u0_u5_u0_n96 ) , .C2( u0_u5_u0_n97 ) , .ZN( u0_u5_u0_n98 ) );
  INV_X1 u0_u5_u0_U51 (.ZN( u0_u5_u0_n169 ) , .A( u0_u5_u0_n91 ) );
  NOR2_X1 u0_u5_u0_U52 (.A2( u0_u5_X_4 ) , .A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n118 ) );
  NOR2_X1 u0_u5_u0_U53 (.A2( u0_u5_X_1 ) , .ZN( u0_u5_u0_n101 ) , .A1( u0_u5_u0_n163 ) );
  NOR2_X1 u0_u5_u0_U54 (.A2( u0_u5_X_3 ) , .A1( u0_u5_X_6 ) , .ZN( u0_u5_u0_n94 ) );
  NOR2_X1 u0_u5_u0_U55 (.A2( u0_u5_X_6 ) , .ZN( u0_u5_u0_n100 ) , .A1( u0_u5_u0_n162 ) );
  NAND2_X1 u0_u5_u0_U56 (.A2( u0_u5_X_4 ) , .A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n144 ) );
  NOR2_X1 u0_u5_u0_U57 (.A2( u0_u5_X_5 ) , .ZN( u0_u5_u0_n136 ) , .A1( u0_u5_u0_n159 ) );
  NAND2_X1 u0_u5_u0_U58 (.A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n138 ) , .A2( u0_u5_u0_n159 ) );
  AND2_X1 u0_u5_u0_U59 (.A2( u0_u5_X_3 ) , .A1( u0_u5_X_6 ) , .ZN( u0_u5_u0_n102 ) );
  NOR2_X1 u0_u5_u0_U6 (.A1( u0_u5_u0_n108 ) , .ZN( u0_u5_u0_n123 ) , .A2( u0_u5_u0_n158 ) );
  AND2_X1 u0_u5_u0_U60 (.A1( u0_u5_X_6 ) , .A2( u0_u5_u0_n162 ) , .ZN( u0_u5_u0_n93 ) );
  INV_X1 u0_u5_u0_U61 (.A( u0_u5_X_4 ) , .ZN( u0_u5_u0_n159 ) );
  INV_X1 u0_u5_u0_U62 (.A( u0_u5_X_1 ) , .ZN( u0_u5_u0_n164 ) );
  INV_X1 u0_u5_u0_U63 (.A( u0_u5_X_3 ) , .ZN( u0_u5_u0_n162 ) );
  AOI211_X1 u0_u5_u0_U64 (.B( u0_u5_u0_n133 ) , .A( u0_u5_u0_n134 ) , .C2( u0_u5_u0_n135 ) , .C1( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n137 ) );
  INV_X1 u0_u5_u0_U65 (.A( u0_u5_u0_n126 ) , .ZN( u0_u5_u0_n168 ) );
  OR4_X1 u0_u5_u0_U66 (.ZN( u0_out5_17 ) , .A4( u0_u5_u0_n122 ) , .A2( u0_u5_u0_n123 ) , .A1( u0_u5_u0_n124 ) , .A3( u0_u5_u0_n170 ) );
  AOI21_X1 u0_u5_u0_U67 (.B2( u0_u5_u0_n107 ) , .ZN( u0_u5_u0_n124 ) , .B1( u0_u5_u0_n128 ) , .A( u0_u5_u0_n161 ) );
  INV_X1 u0_u5_u0_U68 (.A( u0_u5_u0_n111 ) , .ZN( u0_u5_u0_n170 ) );
  OR4_X1 u0_u5_u0_U69 (.ZN( u0_out5_31 ) , .A4( u0_u5_u0_n155 ) , .A2( u0_u5_u0_n156 ) , .A1( u0_u5_u0_n157 ) , .A3( u0_u5_u0_n173 ) );
  OAI21_X1 u0_u5_u0_U7 (.B1( u0_u5_u0_n150 ) , .B2( u0_u5_u0_n158 ) , .A( u0_u5_u0_n172 ) , .ZN( u0_u5_u0_n89 ) );
  AOI21_X1 u0_u5_u0_U70 (.A( u0_u5_u0_n138 ) , .B2( u0_u5_u0_n139 ) , .B1( u0_u5_u0_n140 ) , .ZN( u0_u5_u0_n157 ) );
  INV_X1 u0_u5_u0_U71 (.ZN( u0_u5_u0_n174 ) , .A( u0_u5_u0_n89 ) );
  AOI211_X1 u0_u5_u0_U72 (.B( u0_u5_u0_n104 ) , .A( u0_u5_u0_n105 ) , .ZN( u0_u5_u0_n106 ) , .C2( u0_u5_u0_n113 ) , .C1( u0_u5_u0_n160 ) );
  INV_X1 u0_u5_u0_U73 (.A( u0_u5_u0_n142 ) , .ZN( u0_u5_u0_n165 ) );
  AOI21_X1 u0_u5_u0_U74 (.ZN( u0_u5_u0_n116 ) , .B2( u0_u5_u0_n142 ) , .A( u0_u5_u0_n144 ) , .B1( u0_u5_u0_n166 ) );
  AOI21_X1 u0_u5_u0_U75 (.B2( u0_u5_u0_n141 ) , .B1( u0_u5_u0_n142 ) , .ZN( u0_u5_u0_n156 ) , .A( u0_u5_u0_n161 ) );
  OAI221_X1 u0_u5_u0_U76 (.C1( u0_u5_u0_n121 ) , .ZN( u0_u5_u0_n122 ) , .B2( u0_u5_u0_n127 ) , .A( u0_u5_u0_n143 ) , .B1( u0_u5_u0_n144 ) , .C2( u0_u5_u0_n147 ) );
  AOI21_X1 u0_u5_u0_U77 (.B1( u0_u5_u0_n132 ) , .ZN( u0_u5_u0_n133 ) , .A( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n166 ) );
  OAI22_X1 u0_u5_u0_U78 (.ZN( u0_u5_u0_n105 ) , .A2( u0_u5_u0_n132 ) , .B1( u0_u5_u0_n146 ) , .A1( u0_u5_u0_n147 ) , .B2( u0_u5_u0_n161 ) );
  NAND2_X1 u0_u5_u0_U79 (.ZN( u0_u5_u0_n110 ) , .A2( u0_u5_u0_n132 ) , .A1( u0_u5_u0_n145 ) );
  AND2_X1 u0_u5_u0_U8 (.A1( u0_u5_u0_n114 ) , .A2( u0_u5_u0_n121 ) , .ZN( u0_u5_u0_n146 ) );
  INV_X1 u0_u5_u0_U80 (.A( u0_u5_u0_n119 ) , .ZN( u0_u5_u0_n167 ) );
  NAND2_X1 u0_u5_u0_U81 (.ZN( u0_u5_u0_n148 ) , .A1( u0_u5_u0_n93 ) , .A2( u0_u5_u0_n95 ) );
  NAND2_X1 u0_u5_u0_U82 (.A1( u0_u5_u0_n100 ) , .ZN( u0_u5_u0_n129 ) , .A2( u0_u5_u0_n95 ) );
  NAND2_X1 u0_u5_u0_U83 (.A1( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n128 ) , .A2( u0_u5_u0_n95 ) );
  NOR2_X1 u0_u5_u0_U84 (.A2( u0_u5_X_1 ) , .A1( u0_u5_X_2 ) , .ZN( u0_u5_u0_n92 ) );
  NAND2_X1 u0_u5_u0_U85 (.ZN( u0_u5_u0_n142 ) , .A1( u0_u5_u0_n94 ) , .A2( u0_u5_u0_n95 ) );
  NOR2_X1 u0_u5_u0_U86 (.A2( u0_u5_X_2 ) , .ZN( u0_u5_u0_n103 ) , .A1( u0_u5_u0_n164 ) );
  INV_X1 u0_u5_u0_U87 (.A( u0_u5_X_2 ) , .ZN( u0_u5_u0_n163 ) );
  NAND3_X1 u0_u5_u0_U88 (.ZN( u0_out5_23 ) , .A3( u0_u5_u0_n137 ) , .A1( u0_u5_u0_n168 ) , .A2( u0_u5_u0_n171 ) );
  NAND3_X1 u0_u5_u0_U89 (.A3( u0_u5_u0_n127 ) , .A2( u0_u5_u0_n128 ) , .ZN( u0_u5_u0_n135 ) , .A1( u0_u5_u0_n150 ) );
  NAND2_X1 u0_u5_u0_U9 (.ZN( u0_u5_u0_n113 ) , .A1( u0_u5_u0_n139 ) , .A2( u0_u5_u0_n149 ) );
  NAND3_X1 u0_u5_u0_U90 (.ZN( u0_u5_u0_n117 ) , .A3( u0_u5_u0_n132 ) , .A2( u0_u5_u0_n139 ) , .A1( u0_u5_u0_n148 ) );
  NAND3_X1 u0_u5_u0_U91 (.ZN( u0_u5_u0_n109 ) , .A2( u0_u5_u0_n114 ) , .A3( u0_u5_u0_n140 ) , .A1( u0_u5_u0_n149 ) );
  NAND3_X1 u0_u5_u0_U92 (.ZN( u0_out5_9 ) , .A3( u0_u5_u0_n106 ) , .A2( u0_u5_u0_n171 ) , .A1( u0_u5_u0_n174 ) );
  NAND3_X1 u0_u5_u0_U93 (.A2( u0_u5_u0_n128 ) , .A1( u0_u5_u0_n132 ) , .A3( u0_u5_u0_n146 ) , .ZN( u0_u5_u0_n97 ) );
  NOR2_X1 u0_u5_u1_U10 (.A1( u0_u5_u1_n112 ) , .A2( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n118 ) );
  NAND3_X1 u0_u5_u1_U100 (.ZN( u0_u5_u1_n113 ) , .A1( u0_u5_u1_n120 ) , .A3( u0_u5_u1_n133 ) , .A2( u0_u5_u1_n155 ) );
  OAI21_X1 u0_u5_u1_U11 (.ZN( u0_u5_u1_n101 ) , .B1( u0_u5_u1_n141 ) , .A( u0_u5_u1_n146 ) , .B2( u0_u5_u1_n183 ) );
  AOI21_X1 u0_u5_u1_U12 (.B2( u0_u5_u1_n155 ) , .B1( u0_u5_u1_n156 ) , .ZN( u0_u5_u1_n157 ) , .A( u0_u5_u1_n174 ) );
  NAND2_X1 u0_u5_u1_U13 (.ZN( u0_u5_u1_n140 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n155 ) );
  NAND2_X1 u0_u5_u1_U14 (.A1( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n153 ) );
  INV_X1 u0_u5_u1_U15 (.A( u0_u5_u1_n139 ) , .ZN( u0_u5_u1_n174 ) );
  OR4_X1 u0_u5_u1_U16 (.A4( u0_u5_u1_n106 ) , .A3( u0_u5_u1_n107 ) , .ZN( u0_u5_u1_n108 ) , .A1( u0_u5_u1_n117 ) , .A2( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U17 (.ZN( u0_u5_u1_n106 ) , .A( u0_u5_u1_n112 ) , .B1( u0_u5_u1_n154 ) , .B2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U18 (.A( u0_u5_u1_n101 ) , .ZN( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U19 (.ZN( u0_u5_u1_n107 ) , .B1( u0_u5_u1_n134 ) , .B2( u0_u5_u1_n149 ) , .A( u0_u5_u1_n174 ) );
  INV_X1 u0_u5_u1_U20 (.A( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n171 ) );
  NAND2_X1 u0_u5_u1_U21 (.ZN( u0_u5_u1_n141 ) , .A1( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n156 ) );
  AND2_X1 u0_u5_u1_U22 (.A1( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n161 ) );
  NAND2_X1 u0_u5_u1_U23 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n148 ) );
  NAND2_X1 u0_u5_u1_U24 (.A2( u0_u5_u1_n133 ) , .A1( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n159 ) );
  NAND2_X1 u0_u5_u1_U25 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n120 ) , .ZN( u0_u5_u1_n132 ) );
  INV_X1 u0_u5_u1_U26 (.A( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n178 ) );
  INV_X1 u0_u5_u1_U27 (.A( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n183 ) );
  AND2_X1 u0_u5_u1_U28 (.A1( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n149 ) );
  INV_X1 u0_u5_u1_U29 (.A( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U3 (.A( u0_u5_u1_n159 ) , .ZN( u0_u5_u1_n182 ) );
  OAI221_X1 u0_u5_u1_U30 (.A( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n138 ) , .B2( u0_u5_u1_n152 ) , .C1( u0_u5_u1_n174 ) , .B1( u0_u5_u1_n187 ) );
  INV_X1 u0_u5_u1_U31 (.A( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n187 ) );
  AOI211_X1 u0_u5_u1_U32 (.B( u0_u5_u1_n117 ) , .A( u0_u5_u1_n118 ) , .ZN( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n146 ) , .C1( u0_u5_u1_n159 ) );
  NOR2_X1 u0_u5_u1_U33 (.A1( u0_u5_u1_n168 ) , .A2( u0_u5_u1_n176 ) , .ZN( u0_u5_u1_n98 ) );
  OAI21_X1 u0_u5_u1_U34 (.B2( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n145 ) , .B1( u0_u5_u1_n160 ) , .A( u0_u5_u1_n185 ) );
  INV_X1 u0_u5_u1_U35 (.A( u0_u5_u1_n122 ) , .ZN( u0_u5_u1_n185 ) );
  AOI21_X1 u0_u5_u1_U36 (.B2( u0_u5_u1_n120 ) , .B1( u0_u5_u1_n121 ) , .ZN( u0_u5_u1_n122 ) , .A( u0_u5_u1_n128 ) );
  NAND2_X1 u0_u5_u1_U37 (.A1( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n146 ) , .A2( u0_u5_u1_n160 ) );
  NAND2_X1 u0_u5_u1_U38 (.A2( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n139 ) , .A1( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U39 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n156 ) , .A2( u0_u5_u1_n99 ) );
  AOI221_X1 u0_u5_u1_U4 (.A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .C1( u0_u5_u1_n140 ) , .B2( u0_u5_u1_n141 ) , .ZN( u0_u5_u1_n142 ) , .B1( u0_u5_u1_n175 ) );
  AOI221_X1 u0_u5_u1_U40 (.B1( u0_u5_u1_n140 ) , .ZN( u0_u5_u1_n167 ) , .B2( u0_u5_u1_n172 ) , .C2( u0_u5_u1_n175 ) , .C1( u0_u5_u1_n178 ) , .A( u0_u5_u1_n188 ) );
  INV_X1 u0_u5_u1_U41 (.ZN( u0_u5_u1_n188 ) , .A( u0_u5_u1_n97 ) );
  AOI211_X1 u0_u5_u1_U42 (.A( u0_u5_u1_n118 ) , .C1( u0_u5_u1_n132 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n96 ) , .ZN( u0_u5_u1_n97 ) );
  AOI21_X1 u0_u5_u1_U43 (.B2( u0_u5_u1_n121 ) , .B1( u0_u5_u1_n135 ) , .A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n96 ) );
  NOR2_X1 u0_u5_u1_U44 (.ZN( u0_u5_u1_n117 ) , .A1( u0_u5_u1_n121 ) , .A2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U45 (.A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n130 ) , .B1( u0_u5_u1_n150 ) );
  NAND2_X1 u0_u5_u1_U46 (.ZN( u0_u5_u1_n112 ) , .A1( u0_u5_u1_n169 ) , .A2( u0_u5_u1_n170 ) );
  NAND2_X1 u0_u5_u1_U47 (.ZN( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n95 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U48 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n154 ) , .A2( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U49 (.A2( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n135 ) , .A1( u0_u5_u1_n99 ) );
  AOI211_X1 u0_u5_u1_U5 (.ZN( u0_u5_u1_n124 ) , .A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n145 ) , .C1( u0_u5_u1_n147 ) );
  AOI21_X1 u0_u5_u1_U50 (.A( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n153 ) , .B1( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n158 ) );
  INV_X1 u0_u5_u1_U51 (.A( u0_u5_u1_n160 ) , .ZN( u0_u5_u1_n175 ) );
  NAND2_X1 u0_u5_u1_U52 (.A1( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n116 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U53 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n131 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U54 (.A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n121 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U55 (.A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U56 (.A2( u0_u5_u1_n104 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n133 ) );
  NAND2_X1 u0_u5_u1_U57 (.ZN( u0_u5_u1_n150 ) , .A2( u0_u5_u1_n98 ) , .A1( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U58 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n155 ) , .A2( u0_u5_u1_n95 ) );
  OAI21_X1 u0_u5_u1_U59 (.ZN( u0_u5_u1_n109 ) , .B1( u0_u5_u1_n129 ) , .B2( u0_u5_u1_n160 ) , .A( u0_u5_u1_n167 ) );
  AOI22_X1 u0_u5_u1_U6 (.B2( u0_u5_u1_n136 ) , .A2( u0_u5_u1_n137 ) , .ZN( u0_u5_u1_n143 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  NAND2_X1 u0_u5_u1_U60 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n120 ) );
  NAND2_X1 u0_u5_u1_U61 (.A1( u0_u5_u1_n102 ) , .A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n115 ) );
  NAND2_X1 u0_u5_u1_U62 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n151 ) );
  NAND2_X1 u0_u5_u1_U63 (.A2( u0_u5_u1_n103 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n161 ) );
  INV_X1 u0_u5_u1_U64 (.A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U65 (.A( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U66 (.A2( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n123 ) );
  AOI211_X1 u0_u5_u1_U67 (.B( u0_u5_u1_n162 ) , .A( u0_u5_u1_n163 ) , .C2( u0_u5_u1_n164 ) , .ZN( u0_u5_u1_n165 ) , .C1( u0_u5_u1_n171 ) );
  AOI21_X1 u0_u5_u1_U68 (.A( u0_u5_u1_n160 ) , .B2( u0_u5_u1_n161 ) , .ZN( u0_u5_u1_n162 ) , .B1( u0_u5_u1_n182 ) );
  OR2_X1 u0_u5_u1_U69 (.A2( u0_u5_u1_n157 ) , .A1( u0_u5_u1_n158 ) , .ZN( u0_u5_u1_n163 ) );
  INV_X1 u0_u5_u1_U7 (.A( u0_u5_u1_n147 ) , .ZN( u0_u5_u1_n181 ) );
  NOR2_X1 u0_u5_u1_U70 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n95 ) );
  NOR2_X1 u0_u5_u1_U71 (.A1( u0_u5_X_12 ) , .A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n100 ) );
  NOR2_X1 u0_u5_u1_U72 (.A2( u0_u5_X_8 ) , .A1( u0_u5_u1_n177 ) , .ZN( u0_u5_u1_n99 ) );
  NOR2_X1 u0_u5_u1_U73 (.A2( u0_u5_X_12 ) , .ZN( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n176 ) );
  NOR2_X1 u0_u5_u1_U74 (.A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n105 ) , .A1( u0_u5_u1_n168 ) );
  NAND2_X1 u0_u5_u1_U75 (.A1( u0_u5_X_10 ) , .ZN( u0_u5_u1_n160 ) , .A2( u0_u5_u1_n169 ) );
  NAND2_X1 u0_u5_u1_U76 (.A2( u0_u5_X_10 ) , .A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U77 (.A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n128 ) , .A2( u0_u5_u1_n170 ) );
  AND2_X1 u0_u5_u1_U78 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n104 ) );
  AND2_X1 u0_u5_u1_U79 (.A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n103 ) , .A2( u0_u5_u1_n177 ) );
  AOI22_X1 u0_u5_u1_U8 (.B2( u0_u5_u1_n113 ) , .A2( u0_u5_u1_n114 ) , .ZN( u0_u5_u1_n125 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U80 (.A( u0_u5_X_10 ) , .ZN( u0_u5_u1_n170 ) );
  INV_X1 u0_u5_u1_U81 (.A( u0_u5_X_9 ) , .ZN( u0_u5_u1_n176 ) );
  INV_X1 u0_u5_u1_U82 (.A( u0_u5_X_11 ) , .ZN( u0_u5_u1_n169 ) );
  INV_X1 u0_u5_u1_U83 (.A( u0_u5_X_12 ) , .ZN( u0_u5_u1_n168 ) );
  INV_X1 u0_u5_u1_U84 (.A( u0_u5_X_7 ) , .ZN( u0_u5_u1_n177 ) );
  NAND4_X1 u0_u5_u1_U85 (.ZN( u0_out5_28 ) , .A4( u0_u5_u1_n124 ) , .A3( u0_u5_u1_n125 ) , .A2( u0_u5_u1_n126 ) , .A1( u0_u5_u1_n127 ) );
  OAI21_X1 u0_u5_u1_U86 (.ZN( u0_u5_u1_n127 ) , .B2( u0_u5_u1_n139 ) , .B1( u0_u5_u1_n175 ) , .A( u0_u5_u1_n183 ) );
  OAI21_X1 u0_u5_u1_U87 (.ZN( u0_u5_u1_n126 ) , .B2( u0_u5_u1_n140 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n178 ) );
  NAND4_X1 u0_u5_u1_U88 (.ZN( u0_out5_18 ) , .A4( u0_u5_u1_n165 ) , .A3( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n167 ) , .A2( u0_u5_u1_n186 ) );
  AOI22_X1 u0_u5_u1_U89 (.B2( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U9 (.ZN( u0_u5_u1_n114 ) , .A1( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U90 (.A( u0_u5_u1_n145 ) , .ZN( u0_u5_u1_n186 ) );
  NAND4_X1 u0_u5_u1_U91 (.ZN( u0_out5_2 ) , .A4( u0_u5_u1_n142 ) , .A3( u0_u5_u1_n143 ) , .A2( u0_u5_u1_n144 ) , .A1( u0_u5_u1_n179 ) );
  OAI21_X1 u0_u5_u1_U92 (.B2( u0_u5_u1_n132 ) , .ZN( u0_u5_u1_n144 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U93 (.A( u0_u5_u1_n130 ) , .ZN( u0_u5_u1_n179 ) );
  OR4_X1 u0_u5_u1_U94 (.ZN( u0_out5_13 ) , .A4( u0_u5_u1_n108 ) , .A3( u0_u5_u1_n109 ) , .A2( u0_u5_u1_n110 ) , .A1( u0_u5_u1_n111 ) );
  AOI21_X1 u0_u5_u1_U95 (.ZN( u0_u5_u1_n110 ) , .A( u0_u5_u1_n116 ) , .B1( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U96 (.ZN( u0_u5_u1_n111 ) , .A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n131 ) , .B1( u0_u5_u1_n135 ) );
  NAND3_X1 u0_u5_u1_U97 (.A3( u0_u5_u1_n149 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n164 ) );
  NAND3_X1 u0_u5_u1_U98 (.A3( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n136 ) , .A1( u0_u5_u1_n151 ) );
  NAND3_X1 u0_u5_u1_U99 (.A1( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n137 ) , .A2( u0_u5_u1_n154 ) , .A3( u0_u5_u1_n181 ) );
  OAI22_X1 u0_u5_u2_U10 (.ZN( u0_u5_u2_n109 ) , .A2( u0_u5_u2_n113 ) , .B2( u0_u5_u2_n133 ) , .B1( u0_u5_u2_n167 ) , .A1( u0_u5_u2_n168 ) );
  NAND3_X1 u0_u5_u2_U100 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n98 ) );
  OAI22_X1 u0_u5_u2_U11 (.B1( u0_u5_u2_n151 ) , .A2( u0_u5_u2_n152 ) , .A1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n160 ) , .B2( u0_u5_u2_n168 ) );
  NOR3_X1 u0_u5_u2_U12 (.A1( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n151 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U13 (.ZN( u0_u5_u2_n144 ) , .B2( u0_u5_u2_n155 ) , .A( u0_u5_u2_n172 ) , .B1( u0_u5_u2_n185 ) );
  AOI21_X1 u0_u5_u2_U14 (.B2( u0_u5_u2_n143 ) , .ZN( u0_u5_u2_n145 ) , .B1( u0_u5_u2_n152 ) , .A( u0_u5_u2_n171 ) );
  AOI21_X1 u0_u5_u2_U15 (.B2( u0_u5_u2_n120 ) , .B1( u0_u5_u2_n121 ) , .ZN( u0_u5_u2_n126 ) , .A( u0_u5_u2_n167 ) );
  INV_X1 u0_u5_u2_U16 (.A( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n171 ) );
  INV_X1 u0_u5_u2_U17 (.A( u0_u5_u2_n120 ) , .ZN( u0_u5_u2_n188 ) );
  NAND2_X1 u0_u5_u2_U18 (.A2( u0_u5_u2_n122 ) , .ZN( u0_u5_u2_n150 ) , .A1( u0_u5_u2_n152 ) );
  INV_X1 u0_u5_u2_U19 (.A( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U20 (.A( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n173 ) );
  NAND2_X1 u0_u5_u2_U21 (.A1( u0_u5_u2_n132 ) , .A2( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n157 ) );
  INV_X1 u0_u5_u2_U22 (.A( u0_u5_u2_n113 ) , .ZN( u0_u5_u2_n178 ) );
  INV_X1 u0_u5_u2_U23 (.A( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n175 ) );
  INV_X1 u0_u5_u2_U24 (.A( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n181 ) );
  INV_X1 u0_u5_u2_U25 (.A( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n177 ) );
  INV_X1 u0_u5_u2_U26 (.A( u0_u5_u2_n116 ) , .ZN( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U27 (.A( u0_u5_u2_n131 ) , .ZN( u0_u5_u2_n179 ) );
  INV_X1 u0_u5_u2_U28 (.A( u0_u5_u2_n154 ) , .ZN( u0_u5_u2_n176 ) );
  NAND2_X1 u0_u5_u2_U29 (.A2( u0_u5_u2_n116 ) , .A1( u0_u5_u2_n117 ) , .ZN( u0_u5_u2_n118 ) );
  NOR2_X1 u0_u5_u2_U3 (.ZN( u0_u5_u2_n121 ) , .A2( u0_u5_u2_n177 ) , .A1( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U30 (.A( u0_u5_u2_n132 ) , .ZN( u0_u5_u2_n182 ) );
  INV_X1 u0_u5_u2_U31 (.A( u0_u5_u2_n158 ) , .ZN( u0_u5_u2_n183 ) );
  OAI21_X1 u0_u5_u2_U32 (.A( u0_u5_u2_n156 ) , .B1( u0_u5_u2_n157 ) , .ZN( u0_u5_u2_n158 ) , .B2( u0_u5_u2_n179 ) );
  NOR2_X1 u0_u5_u2_U33 (.ZN( u0_u5_u2_n156 ) , .A1( u0_u5_u2_n166 ) , .A2( u0_u5_u2_n169 ) );
  NOR2_X1 u0_u5_u2_U34 (.A2( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n140 ) );
  NOR2_X1 u0_u5_u2_U35 (.A2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n153 ) , .A1( u0_u5_u2_n156 ) );
  AOI211_X1 u0_u5_u2_U36 (.ZN( u0_u5_u2_n130 ) , .C1( u0_u5_u2_n138 ) , .C2( u0_u5_u2_n179 ) , .B( u0_u5_u2_n96 ) , .A( u0_u5_u2_n97 ) );
  OAI22_X1 u0_u5_u2_U37 (.B1( u0_u5_u2_n133 ) , .A2( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n152 ) , .B2( u0_u5_u2_n168 ) , .ZN( u0_u5_u2_n97 ) );
  OAI221_X1 u0_u5_u2_U38 (.B1( u0_u5_u2_n113 ) , .C1( u0_u5_u2_n132 ) , .A( u0_u5_u2_n149 ) , .B2( u0_u5_u2_n171 ) , .C2( u0_u5_u2_n172 ) , .ZN( u0_u5_u2_n96 ) );
  OAI221_X1 u0_u5_u2_U39 (.A( u0_u5_u2_n115 ) , .C2( u0_u5_u2_n123 ) , .B2( u0_u5_u2_n143 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n163 ) , .C1( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U4 (.A( u0_u5_u2_n134 ) , .ZN( u0_u5_u2_n185 ) );
  OAI21_X1 u0_u5_u2_U40 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n115 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n178 ) );
  OAI221_X1 u0_u5_u2_U41 (.A( u0_u5_u2_n135 ) , .B2( u0_u5_u2_n136 ) , .B1( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n162 ) , .C2( u0_u5_u2_n167 ) , .C1( u0_u5_u2_n185 ) );
  AND3_X1 u0_u5_u2_U42 (.A3( u0_u5_u2_n131 ) , .A2( u0_u5_u2_n132 ) , .A1( u0_u5_u2_n133 ) , .ZN( u0_u5_u2_n136 ) );
  AOI22_X1 u0_u5_u2_U43 (.ZN( u0_u5_u2_n135 ) , .B1( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n156 ) , .B2( u0_u5_u2_n180 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U44 (.ZN( u0_u5_u2_n149 ) , .B1( u0_u5_u2_n173 ) , .B2( u0_u5_u2_n188 ) , .A( u0_u5_u2_n95 ) );
  AND3_X1 u0_u5_u2_U45 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n95 ) );
  OAI21_X1 u0_u5_u2_U46 (.A( u0_u5_u2_n141 ) , .B2( u0_u5_u2_n142 ) , .ZN( u0_u5_u2_n146 ) , .B1( u0_u5_u2_n153 ) );
  OAI21_X1 u0_u5_u2_U47 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n141 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n177 ) );
  NOR3_X1 u0_u5_u2_U48 (.ZN( u0_u5_u2_n142 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n178 ) , .A1( u0_u5_u2_n181 ) );
  OAI21_X1 u0_u5_u2_U49 (.A( u0_u5_u2_n101 ) , .B2( u0_u5_u2_n121 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n164 ) );
  INV_X1 u0_u5_u2_U5 (.A( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n184 ) );
  NAND2_X1 u0_u5_u2_U50 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n155 ) );
  NAND2_X1 u0_u5_u2_U51 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n143 ) );
  NAND2_X1 u0_u5_u2_U52 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n152 ) );
  NAND2_X1 u0_u5_u2_U53 (.A1( u0_u5_u2_n100 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n132 ) );
  INV_X1 u0_u5_u2_U54 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U55 (.A( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n167 ) );
  NAND2_X1 u0_u5_u2_U56 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n113 ) );
  NAND2_X1 u0_u5_u2_U57 (.A1( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n131 ) );
  NAND2_X1 u0_u5_u2_U58 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n139 ) );
  NAND2_X1 u0_u5_u2_U59 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n133 ) );
  NOR4_X1 u0_u5_u2_U6 (.A4( u0_u5_u2_n124 ) , .A3( u0_u5_u2_n125 ) , .A2( u0_u5_u2_n126 ) , .A1( u0_u5_u2_n127 ) , .ZN( u0_u5_u2_n128 ) );
  NAND2_X1 u0_u5_u2_U60 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n103 ) , .ZN( u0_u5_u2_n154 ) );
  NAND2_X1 u0_u5_u2_U61 (.A2( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n104 ) , .ZN( u0_u5_u2_n119 ) );
  NAND2_X1 u0_u5_u2_U62 (.A2( u0_u5_u2_n107 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n123 ) );
  NAND2_X1 u0_u5_u2_U63 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n122 ) );
  INV_X1 u0_u5_u2_U64 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n172 ) );
  NAND2_X1 u0_u5_u2_U65 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n102 ) , .ZN( u0_u5_u2_n116 ) );
  NAND2_X1 u0_u5_u2_U66 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n120 ) );
  NAND2_X1 u0_u5_u2_U67 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n117 ) );
  INV_X1 u0_u5_u2_U68 (.ZN( u0_u5_u2_n187 ) , .A( u0_u5_u2_n99 ) );
  OAI21_X1 u0_u5_u2_U69 (.B1( u0_u5_u2_n137 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n98 ) , .ZN( u0_u5_u2_n99 ) );
  AOI21_X1 u0_u5_u2_U7 (.B2( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n127 ) , .A( u0_u5_u2_n137 ) , .B1( u0_u5_u2_n155 ) );
  NOR2_X1 u0_u5_u2_U70 (.A2( u0_u5_X_16 ) , .ZN( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n166 ) );
  NOR2_X1 u0_u5_u2_U71 (.A2( u0_u5_X_13 ) , .A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n100 ) );
  NOR2_X1 u0_u5_u2_U72 (.A2( u0_u5_X_16 ) , .A1( u0_u5_X_17 ) , .ZN( u0_u5_u2_n138 ) );
  NOR2_X1 u0_u5_u2_U73 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n104 ) );
  NOR2_X1 u0_u5_u2_U74 (.A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n174 ) );
  NOR2_X1 u0_u5_u2_U75 (.A2( u0_u5_X_15 ) , .ZN( u0_u5_u2_n102 ) , .A1( u0_u5_u2_n165 ) );
  NOR2_X1 u0_u5_u2_U76 (.A2( u0_u5_X_17 ) , .ZN( u0_u5_u2_n114 ) , .A1( u0_u5_u2_n169 ) );
  AND2_X1 u0_u5_u2_U77 (.A1( u0_u5_X_15 ) , .ZN( u0_u5_u2_n105 ) , .A2( u0_u5_u2_n165 ) );
  AND2_X1 u0_u5_u2_U78 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n107 ) );
  AND2_X1 u0_u5_u2_U79 (.A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n174 ) );
  AOI21_X1 u0_u5_u2_U8 (.ZN( u0_u5_u2_n124 ) , .B1( u0_u5_u2_n131 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n172 ) );
  AND2_X1 u0_u5_u2_U80 (.A1( u0_u5_X_13 ) , .A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n108 ) );
  INV_X1 u0_u5_u2_U81 (.A( u0_u5_X_16 ) , .ZN( u0_u5_u2_n169 ) );
  INV_X1 u0_u5_u2_U82 (.A( u0_u5_X_17 ) , .ZN( u0_u5_u2_n166 ) );
  INV_X1 u0_u5_u2_U83 (.A( u0_u5_X_13 ) , .ZN( u0_u5_u2_n174 ) );
  INV_X1 u0_u5_u2_U84 (.A( u0_u5_X_18 ) , .ZN( u0_u5_u2_n165 ) );
  NAND4_X1 u0_u5_u2_U85 (.ZN( u0_out5_30 ) , .A4( u0_u5_u2_n147 ) , .A3( u0_u5_u2_n148 ) , .A2( u0_u5_u2_n149 ) , .A1( u0_u5_u2_n187 ) );
  NOR3_X1 u0_u5_u2_U86 (.A3( u0_u5_u2_n144 ) , .A2( u0_u5_u2_n145 ) , .A1( u0_u5_u2_n146 ) , .ZN( u0_u5_u2_n147 ) );
  AOI21_X1 u0_u5_u2_U87 (.B2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n148 ) , .A( u0_u5_u2_n162 ) , .B1( u0_u5_u2_n182 ) );
  NAND4_X1 u0_u5_u2_U88 (.ZN( u0_out5_24 ) , .A4( u0_u5_u2_n111 ) , .A3( u0_u5_u2_n112 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n187 ) );
  AOI221_X1 u0_u5_u2_U89 (.A( u0_u5_u2_n109 ) , .B1( u0_u5_u2_n110 ) , .ZN( u0_u5_u2_n111 ) , .C1( u0_u5_u2_n134 ) , .C2( u0_u5_u2_n170 ) , .B2( u0_u5_u2_n173 ) );
  AOI21_X1 u0_u5_u2_U9 (.B2( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n125 ) , .A( u0_u5_u2_n171 ) , .B1( u0_u5_u2_n184 ) );
  AOI21_X1 u0_u5_u2_U90 (.ZN( u0_u5_u2_n112 ) , .B2( u0_u5_u2_n156 ) , .A( u0_u5_u2_n164 ) , .B1( u0_u5_u2_n181 ) );
  NAND4_X1 u0_u5_u2_U91 (.ZN( u0_out5_16 ) , .A4( u0_u5_u2_n128 ) , .A3( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n186 ) );
  AOI22_X1 u0_u5_u2_U92 (.A2( u0_u5_u2_n118 ) , .ZN( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n140 ) , .B1( u0_u5_u2_n157 ) , .B2( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U93 (.A( u0_u5_u2_n163 ) , .ZN( u0_u5_u2_n186 ) );
  OR4_X1 u0_u5_u2_U94 (.ZN( u0_out5_6 ) , .A4( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n162 ) , .A2( u0_u5_u2_n163 ) , .A1( u0_u5_u2_n164 ) );
  OR3_X1 u0_u5_u2_U95 (.A2( u0_u5_u2_n159 ) , .A1( u0_u5_u2_n160 ) , .ZN( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n183 ) );
  AOI21_X1 u0_u5_u2_U96 (.B2( u0_u5_u2_n154 ) , .B1( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n159 ) , .A( u0_u5_u2_n167 ) );
  NAND3_X1 u0_u5_u2_U97 (.A2( u0_u5_u2_n117 ) , .A1( u0_u5_u2_n122 ) , .A3( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n134 ) );
  NAND3_X1 u0_u5_u2_U98 (.ZN( u0_u5_u2_n110 ) , .A2( u0_u5_u2_n131 ) , .A3( u0_u5_u2_n139 ) , .A1( u0_u5_u2_n154 ) );
  NAND3_X1 u0_u5_u2_U99 (.A2( u0_u5_u2_n100 ) , .ZN( u0_u5_u2_n101 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n114 ) );
  XOR2_X1 u0_u7_U1 (.B( u0_K8_9 ) , .A( u0_R6_6 ) , .Z( u0_u7_X_9 ) );
  XOR2_X1 u0_u7_U16 (.B( u0_K8_3 ) , .A( u0_R6_2 ) , .Z( u0_u7_X_3 ) );
  XOR2_X1 u0_u7_U2 (.B( u0_K8_8 ) , .A( u0_R6_5 ) , .Z( u0_u7_X_8 ) );
  XOR2_X1 u0_u7_U27 (.B( u0_K8_2 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_2 ) );
  XOR2_X1 u0_u7_U3 (.B( u0_K8_7 ) , .A( u0_R6_4 ) , .Z( u0_u7_X_7 ) );
  XOR2_X1 u0_u7_U38 (.B( u0_K8_1 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_1 ) );
  XOR2_X1 u0_u7_U4 (.B( u0_K8_6 ) , .A( u0_R6_5 ) , .Z( u0_u7_X_6 ) );
  XOR2_X1 u0_u7_U46 (.B( u0_K8_12 ) , .A( u0_R6_9 ) , .Z( u0_u7_X_12 ) );
  XOR2_X1 u0_u7_U47 (.B( u0_K8_11 ) , .A( u0_R6_8 ) , .Z( u0_u7_X_11 ) );
  XOR2_X1 u0_u7_U48 (.B( u0_K8_10 ) , .A( u0_R6_7 ) , .Z( u0_u7_X_10 ) );
  XOR2_X1 u0_u7_U5 (.B( u0_K8_5 ) , .A( u0_R6_4 ) , .Z( u0_u7_X_5 ) );
  XOR2_X1 u0_u7_U6 (.B( u0_K8_4 ) , .A( u0_R6_3 ) , .Z( u0_u7_X_4 ) );
  AND3_X1 u0_u7_u0_U10 (.A2( u0_u7_u0_n112 ) , .ZN( u0_u7_u0_n127 ) , .A3( u0_u7_u0_n130 ) , .A1( u0_u7_u0_n148 ) );
  NAND2_X1 u0_u7_u0_U11 (.ZN( u0_u7_u0_n113 ) , .A1( u0_u7_u0_n139 ) , .A2( u0_u7_u0_n149 ) );
  AND2_X1 u0_u7_u0_U12 (.ZN( u0_u7_u0_n107 ) , .A1( u0_u7_u0_n130 ) , .A2( u0_u7_u0_n140 ) );
  AND2_X1 u0_u7_u0_U13 (.A2( u0_u7_u0_n129 ) , .A1( u0_u7_u0_n130 ) , .ZN( u0_u7_u0_n151 ) );
  AND2_X1 u0_u7_u0_U14 (.A1( u0_u7_u0_n108 ) , .A2( u0_u7_u0_n125 ) , .ZN( u0_u7_u0_n145 ) );
  INV_X1 u0_u7_u0_U15 (.A( u0_u7_u0_n143 ) , .ZN( u0_u7_u0_n173 ) );
  NOR2_X1 u0_u7_u0_U16 (.A2( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n147 ) , .A1( u0_u7_u0_n160 ) );
  INV_X1 u0_u7_u0_U17 (.ZN( u0_u7_u0_n172 ) , .A( u0_u7_u0_n88 ) );
  OAI222_X1 u0_u7_u0_U18 (.C1( u0_u7_u0_n108 ) , .A1( u0_u7_u0_n125 ) , .B2( u0_u7_u0_n128 ) , .B1( u0_u7_u0_n144 ) , .A2( u0_u7_u0_n158 ) , .C2( u0_u7_u0_n161 ) , .ZN( u0_u7_u0_n88 ) );
  NOR2_X1 u0_u7_u0_U19 (.A1( u0_u7_u0_n163 ) , .A2( u0_u7_u0_n164 ) , .ZN( u0_u7_u0_n95 ) );
  AOI21_X1 u0_u7_u0_U20 (.B1( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n132 ) , .A( u0_u7_u0_n165 ) , .B2( u0_u7_u0_n93 ) );
  INV_X1 u0_u7_u0_U21 (.A( u0_u7_u0_n142 ) , .ZN( u0_u7_u0_n165 ) );
  OAI22_X1 u0_u7_u0_U22 (.B1( u0_u7_u0_n125 ) , .ZN( u0_u7_u0_n126 ) , .A1( u0_u7_u0_n138 ) , .A2( u0_u7_u0_n146 ) , .B2( u0_u7_u0_n147 ) );
  OAI22_X1 u0_u7_u0_U23 (.B1( u0_u7_u0_n131 ) , .A1( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n147 ) , .A2( u0_u7_u0_n90 ) , .ZN( u0_u7_u0_n91 ) );
  AND3_X1 u0_u7_u0_U24 (.A3( u0_u7_u0_n121 ) , .A2( u0_u7_u0_n125 ) , .A1( u0_u7_u0_n148 ) , .ZN( u0_u7_u0_n90 ) );
  NAND2_X1 u0_u7_u0_U25 (.A1( u0_u7_u0_n100 ) , .A2( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n125 ) );
  INV_X1 u0_u7_u0_U26 (.A( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n161 ) );
  AOI22_X1 u0_u7_u0_U27 (.B2( u0_u7_u0_n109 ) , .A2( u0_u7_u0_n110 ) , .ZN( u0_u7_u0_n111 ) , .B1( u0_u7_u0_n118 ) , .A1( u0_u7_u0_n160 ) );
  NAND2_X1 u0_u7_u0_U28 (.A1( u0_u7_u0_n100 ) , .ZN( u0_u7_u0_n129 ) , .A2( u0_u7_u0_n95 ) );
  INV_X1 u0_u7_u0_U29 (.A( u0_u7_u0_n118 ) , .ZN( u0_u7_u0_n158 ) );
  INV_X1 u0_u7_u0_U3 (.A( u0_u7_u0_n113 ) , .ZN( u0_u7_u0_n166 ) );
  AOI21_X1 u0_u7_u0_U30 (.ZN( u0_u7_u0_n104 ) , .B1( u0_u7_u0_n107 ) , .B2( u0_u7_u0_n141 ) , .A( u0_u7_u0_n144 ) );
  AOI21_X1 u0_u7_u0_U31 (.B1( u0_u7_u0_n127 ) , .B2( u0_u7_u0_n129 ) , .A( u0_u7_u0_n138 ) , .ZN( u0_u7_u0_n96 ) );
  AOI21_X1 u0_u7_u0_U32 (.ZN( u0_u7_u0_n116 ) , .B2( u0_u7_u0_n142 ) , .A( u0_u7_u0_n144 ) , .B1( u0_u7_u0_n166 ) );
  NOR2_X1 u0_u7_u0_U33 (.A1( u0_u7_u0_n120 ) , .ZN( u0_u7_u0_n143 ) , .A2( u0_u7_u0_n167 ) );
  OAI221_X1 u0_u7_u0_U34 (.C1( u0_u7_u0_n112 ) , .ZN( u0_u7_u0_n120 ) , .B1( u0_u7_u0_n138 ) , .B2( u0_u7_u0_n141 ) , .C2( u0_u7_u0_n147 ) , .A( u0_u7_u0_n172 ) );
  AOI211_X1 u0_u7_u0_U35 (.B( u0_u7_u0_n115 ) , .A( u0_u7_u0_n116 ) , .C2( u0_u7_u0_n117 ) , .C1( u0_u7_u0_n118 ) , .ZN( u0_u7_u0_n119 ) );
  NAND2_X1 u0_u7_u0_U36 (.A2( u0_u7_u0_n100 ) , .A1( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n139 ) );
  NAND2_X1 u0_u7_u0_U37 (.A2( u0_u7_u0_n100 ) , .ZN( u0_u7_u0_n131 ) , .A1( u0_u7_u0_n92 ) );
  NAND2_X1 u0_u7_u0_U38 (.A1( u0_u7_u0_n101 ) , .A2( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n150 ) );
  INV_X1 u0_u7_u0_U39 (.A( u0_u7_u0_n138 ) , .ZN( u0_u7_u0_n160 ) );
  AOI21_X1 u0_u7_u0_U4 (.B1( u0_u7_u0_n114 ) , .ZN( u0_u7_u0_n115 ) , .B2( u0_u7_u0_n129 ) , .A( u0_u7_u0_n161 ) );
  NAND2_X1 u0_u7_u0_U40 (.A1( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n128 ) , .A2( u0_u7_u0_n95 ) );
  NAND2_X1 u0_u7_u0_U41 (.ZN( u0_u7_u0_n148 ) , .A1( u0_u7_u0_n93 ) , .A2( u0_u7_u0_n95 ) );
  NAND2_X1 u0_u7_u0_U42 (.A2( u0_u7_u0_n102 ) , .A1( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n149 ) );
  NAND2_X1 u0_u7_u0_U43 (.A2( u0_u7_u0_n102 ) , .ZN( u0_u7_u0_n114 ) , .A1( u0_u7_u0_n92 ) );
  NAND2_X1 u0_u7_u0_U44 (.A2( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n121 ) , .A1( u0_u7_u0_n93 ) );
  NAND2_X1 u0_u7_u0_U45 (.ZN( u0_u7_u0_n112 ) , .A2( u0_u7_u0_n92 ) , .A1( u0_u7_u0_n93 ) );
  OR3_X1 u0_u7_u0_U46 (.A3( u0_u7_u0_n152 ) , .A2( u0_u7_u0_n153 ) , .A1( u0_u7_u0_n154 ) , .ZN( u0_u7_u0_n155 ) );
  AOI21_X1 u0_u7_u0_U47 (.A( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n145 ) , .B1( u0_u7_u0_n146 ) , .ZN( u0_u7_u0_n154 ) );
  AOI21_X1 u0_u7_u0_U48 (.B2( u0_u7_u0_n150 ) , .B1( u0_u7_u0_n151 ) , .ZN( u0_u7_u0_n152 ) , .A( u0_u7_u0_n158 ) );
  AOI21_X1 u0_u7_u0_U49 (.A( u0_u7_u0_n147 ) , .B2( u0_u7_u0_n148 ) , .B1( u0_u7_u0_n149 ) , .ZN( u0_u7_u0_n153 ) );
  AOI21_X1 u0_u7_u0_U5 (.B2( u0_u7_u0_n131 ) , .ZN( u0_u7_u0_n134 ) , .B1( u0_u7_u0_n151 ) , .A( u0_u7_u0_n158 ) );
  INV_X1 u0_u7_u0_U50 (.ZN( u0_u7_u0_n171 ) , .A( u0_u7_u0_n99 ) );
  OAI211_X1 u0_u7_u0_U51 (.C2( u0_u7_u0_n140 ) , .C1( u0_u7_u0_n161 ) , .A( u0_u7_u0_n169 ) , .B( u0_u7_u0_n98 ) , .ZN( u0_u7_u0_n99 ) );
  INV_X1 u0_u7_u0_U52 (.ZN( u0_u7_u0_n169 ) , .A( u0_u7_u0_n91 ) );
  AOI211_X1 u0_u7_u0_U53 (.C1( u0_u7_u0_n118 ) , .A( u0_u7_u0_n123 ) , .B( u0_u7_u0_n96 ) , .C2( u0_u7_u0_n97 ) , .ZN( u0_u7_u0_n98 ) );
  NOR2_X1 u0_u7_u0_U54 (.A2( u0_u7_X_4 ) , .A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n118 ) );
  NOR2_X1 u0_u7_u0_U55 (.A2( u0_u7_X_2 ) , .ZN( u0_u7_u0_n103 ) , .A1( u0_u7_u0_n164 ) );
  NOR2_X1 u0_u7_u0_U56 (.A2( u0_u7_X_1 ) , .A1( u0_u7_X_2 ) , .ZN( u0_u7_u0_n92 ) );
  NOR2_X1 u0_u7_u0_U57 (.A2( u0_u7_X_1 ) , .ZN( u0_u7_u0_n101 ) , .A1( u0_u7_u0_n163 ) );
  NAND2_X1 u0_u7_u0_U58 (.A2( u0_u7_X_4 ) , .A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n144 ) );
  NOR2_X1 u0_u7_u0_U59 (.A2( u0_u7_X_5 ) , .ZN( u0_u7_u0_n136 ) , .A1( u0_u7_u0_n159 ) );
  NOR2_X1 u0_u7_u0_U6 (.A1( u0_u7_u0_n108 ) , .ZN( u0_u7_u0_n123 ) , .A2( u0_u7_u0_n158 ) );
  NAND2_X1 u0_u7_u0_U60 (.A1( u0_u7_X_5 ) , .ZN( u0_u7_u0_n138 ) , .A2( u0_u7_u0_n159 ) );
  NOR2_X1 u0_u7_u0_U61 (.A2( u0_u7_X_3 ) , .A1( u0_u7_X_6 ) , .ZN( u0_u7_u0_n94 ) );
  AND2_X1 u0_u7_u0_U62 (.A2( u0_u7_X_3 ) , .A1( u0_u7_X_6 ) , .ZN( u0_u7_u0_n102 ) );
  AND2_X1 u0_u7_u0_U63 (.A1( u0_u7_X_6 ) , .A2( u0_u7_u0_n162 ) , .ZN( u0_u7_u0_n93 ) );
  INV_X1 u0_u7_u0_U64 (.A( u0_u7_X_4 ) , .ZN( u0_u7_u0_n159 ) );
  INV_X1 u0_u7_u0_U65 (.A( u0_u7_X_1 ) , .ZN( u0_u7_u0_n164 ) );
  INV_X1 u0_u7_u0_U66 (.A( u0_u7_X_2 ) , .ZN( u0_u7_u0_n163 ) );
  INV_X1 u0_u7_u0_U67 (.A( u0_u7_u0_n126 ) , .ZN( u0_u7_u0_n168 ) );
  AOI211_X1 u0_u7_u0_U68 (.B( u0_u7_u0_n133 ) , .A( u0_u7_u0_n134 ) , .C2( u0_u7_u0_n135 ) , .C1( u0_u7_u0_n136 ) , .ZN( u0_u7_u0_n137 ) );
  OR4_X1 u0_u7_u0_U69 (.ZN( u0_out7_17 ) , .A4( u0_u7_u0_n122 ) , .A2( u0_u7_u0_n123 ) , .A1( u0_u7_u0_n124 ) , .A3( u0_u7_u0_n170 ) );
  OAI21_X1 u0_u7_u0_U7 (.B1( u0_u7_u0_n150 ) , .B2( u0_u7_u0_n158 ) , .A( u0_u7_u0_n172 ) , .ZN( u0_u7_u0_n89 ) );
  AOI21_X1 u0_u7_u0_U70 (.B2( u0_u7_u0_n107 ) , .ZN( u0_u7_u0_n124 ) , .B1( u0_u7_u0_n128 ) , .A( u0_u7_u0_n161 ) );
  INV_X1 u0_u7_u0_U71 (.A( u0_u7_u0_n111 ) , .ZN( u0_u7_u0_n170 ) );
  OR4_X1 u0_u7_u0_U72 (.ZN( u0_out7_31 ) , .A4( u0_u7_u0_n155 ) , .A2( u0_u7_u0_n156 ) , .A1( u0_u7_u0_n157 ) , .A3( u0_u7_u0_n173 ) );
  AOI21_X1 u0_u7_u0_U73 (.A( u0_u7_u0_n138 ) , .B2( u0_u7_u0_n139 ) , .B1( u0_u7_u0_n140 ) , .ZN( u0_u7_u0_n157 ) );
  AOI21_X1 u0_u7_u0_U74 (.B2( u0_u7_u0_n141 ) , .B1( u0_u7_u0_n142 ) , .ZN( u0_u7_u0_n156 ) , .A( u0_u7_u0_n161 ) );
  INV_X1 u0_u7_u0_U75 (.ZN( u0_u7_u0_n174 ) , .A( u0_u7_u0_n89 ) );
  AOI211_X1 u0_u7_u0_U76 (.B( u0_u7_u0_n104 ) , .A( u0_u7_u0_n105 ) , .ZN( u0_u7_u0_n106 ) , .C2( u0_u7_u0_n113 ) , .C1( u0_u7_u0_n160 ) );
  OAI221_X1 u0_u7_u0_U77 (.C1( u0_u7_u0_n121 ) , .ZN( u0_u7_u0_n122 ) , .B2( u0_u7_u0_n127 ) , .A( u0_u7_u0_n143 ) , .B1( u0_u7_u0_n144 ) , .C2( u0_u7_u0_n147 ) );
  NOR2_X1 u0_u7_u0_U78 (.A2( u0_u7_X_6 ) , .ZN( u0_u7_u0_n100 ) , .A1( u0_u7_u0_n162 ) );
  INV_X1 u0_u7_u0_U79 (.A( u0_u7_X_3 ) , .ZN( u0_u7_u0_n162 ) );
  AND2_X1 u0_u7_u0_U8 (.A1( u0_u7_u0_n114 ) , .A2( u0_u7_u0_n121 ) , .ZN( u0_u7_u0_n146 ) );
  AOI21_X1 u0_u7_u0_U80 (.B1( u0_u7_u0_n132 ) , .ZN( u0_u7_u0_n133 ) , .A( u0_u7_u0_n144 ) , .B2( u0_u7_u0_n166 ) );
  OAI22_X1 u0_u7_u0_U81 (.ZN( u0_u7_u0_n105 ) , .A2( u0_u7_u0_n132 ) , .B1( u0_u7_u0_n146 ) , .A1( u0_u7_u0_n147 ) , .B2( u0_u7_u0_n161 ) );
  NAND2_X1 u0_u7_u0_U82 (.ZN( u0_u7_u0_n110 ) , .A2( u0_u7_u0_n132 ) , .A1( u0_u7_u0_n145 ) );
  INV_X1 u0_u7_u0_U83 (.A( u0_u7_u0_n119 ) , .ZN( u0_u7_u0_n167 ) );
  NAND2_X1 u0_u7_u0_U84 (.A2( u0_u7_u0_n103 ) , .ZN( u0_u7_u0_n140 ) , .A1( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U85 (.A1( u0_u7_u0_n101 ) , .ZN( u0_u7_u0_n130 ) , .A2( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U86 (.ZN( u0_u7_u0_n108 ) , .A1( u0_u7_u0_n92 ) , .A2( u0_u7_u0_n94 ) );
  NAND2_X1 u0_u7_u0_U87 (.ZN( u0_u7_u0_n142 ) , .A1( u0_u7_u0_n94 ) , .A2( u0_u7_u0_n95 ) );
  NAND3_X1 u0_u7_u0_U88 (.ZN( u0_out7_23 ) , .A3( u0_u7_u0_n137 ) , .A1( u0_u7_u0_n168 ) , .A2( u0_u7_u0_n171 ) );
  NAND3_X1 u0_u7_u0_U89 (.A3( u0_u7_u0_n127 ) , .A2( u0_u7_u0_n128 ) , .ZN( u0_u7_u0_n135 ) , .A1( u0_u7_u0_n150 ) );
  AND2_X1 u0_u7_u0_U9 (.A1( u0_u7_u0_n131 ) , .ZN( u0_u7_u0_n141 ) , .A2( u0_u7_u0_n150 ) );
  NAND3_X1 u0_u7_u0_U90 (.ZN( u0_u7_u0_n117 ) , .A3( u0_u7_u0_n132 ) , .A2( u0_u7_u0_n139 ) , .A1( u0_u7_u0_n148 ) );
  NAND3_X1 u0_u7_u0_U91 (.ZN( u0_u7_u0_n109 ) , .A2( u0_u7_u0_n114 ) , .A3( u0_u7_u0_n140 ) , .A1( u0_u7_u0_n149 ) );
  NAND3_X1 u0_u7_u0_U92 (.ZN( u0_out7_9 ) , .A3( u0_u7_u0_n106 ) , .A2( u0_u7_u0_n171 ) , .A1( u0_u7_u0_n174 ) );
  NAND3_X1 u0_u7_u0_U93 (.A2( u0_u7_u0_n128 ) , .A1( u0_u7_u0_n132 ) , .A3( u0_u7_u0_n146 ) , .ZN( u0_u7_u0_n97 ) );
  AOI21_X1 u0_u7_u1_U10 (.B2( u0_u7_u1_n155 ) , .B1( u0_u7_u1_n156 ) , .ZN( u0_u7_u1_n157 ) , .A( u0_u7_u1_n174 ) );
  NAND3_X1 u0_u7_u1_U100 (.ZN( u0_u7_u1_n113 ) , .A1( u0_u7_u1_n120 ) , .A3( u0_u7_u1_n133 ) , .A2( u0_u7_u1_n155 ) );
  NAND2_X1 u0_u7_u1_U11 (.ZN( u0_u7_u1_n140 ) , .A2( u0_u7_u1_n150 ) , .A1( u0_u7_u1_n155 ) );
  NAND2_X1 u0_u7_u1_U12 (.A1( u0_u7_u1_n131 ) , .ZN( u0_u7_u1_n147 ) , .A2( u0_u7_u1_n153 ) );
  AOI22_X1 u0_u7_u1_U13 (.B2( u0_u7_u1_n136 ) , .A2( u0_u7_u1_n137 ) , .ZN( u0_u7_u1_n143 ) , .A1( u0_u7_u1_n171 ) , .B1( u0_u7_u1_n173 ) );
  INV_X1 u0_u7_u1_U14 (.A( u0_u7_u1_n147 ) , .ZN( u0_u7_u1_n181 ) );
  INV_X1 u0_u7_u1_U15 (.A( u0_u7_u1_n139 ) , .ZN( u0_u7_u1_n174 ) );
  OR4_X1 u0_u7_u1_U16 (.A4( u0_u7_u1_n106 ) , .A3( u0_u7_u1_n107 ) , .ZN( u0_u7_u1_n108 ) , .A1( u0_u7_u1_n117 ) , .A2( u0_u7_u1_n184 ) );
  AOI21_X1 u0_u7_u1_U17 (.ZN( u0_u7_u1_n106 ) , .A( u0_u7_u1_n112 ) , .B1( u0_u7_u1_n154 ) , .B2( u0_u7_u1_n156 ) );
  AOI21_X1 u0_u7_u1_U18 (.ZN( u0_u7_u1_n107 ) , .B1( u0_u7_u1_n134 ) , .B2( u0_u7_u1_n149 ) , .A( u0_u7_u1_n174 ) );
  INV_X1 u0_u7_u1_U19 (.A( u0_u7_u1_n101 ) , .ZN( u0_u7_u1_n184 ) );
  INV_X1 u0_u7_u1_U20 (.A( u0_u7_u1_n112 ) , .ZN( u0_u7_u1_n171 ) );
  NAND2_X1 u0_u7_u1_U21 (.ZN( u0_u7_u1_n141 ) , .A1( u0_u7_u1_n153 ) , .A2( u0_u7_u1_n156 ) );
  AND2_X1 u0_u7_u1_U22 (.A1( u0_u7_u1_n123 ) , .ZN( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n161 ) );
  NAND2_X1 u0_u7_u1_U23 (.A2( u0_u7_u1_n115 ) , .A1( u0_u7_u1_n116 ) , .ZN( u0_u7_u1_n148 ) );
  NAND2_X1 u0_u7_u1_U24 (.A2( u0_u7_u1_n133 ) , .A1( u0_u7_u1_n135 ) , .ZN( u0_u7_u1_n159 ) );
  NAND2_X1 u0_u7_u1_U25 (.A2( u0_u7_u1_n115 ) , .A1( u0_u7_u1_n120 ) , .ZN( u0_u7_u1_n132 ) );
  INV_X1 u0_u7_u1_U26 (.A( u0_u7_u1_n154 ) , .ZN( u0_u7_u1_n178 ) );
  INV_X1 u0_u7_u1_U27 (.A( u0_u7_u1_n151 ) , .ZN( u0_u7_u1_n183 ) );
  AND2_X1 u0_u7_u1_U28 (.A1( u0_u7_u1_n129 ) , .A2( u0_u7_u1_n133 ) , .ZN( u0_u7_u1_n149 ) );
  INV_X1 u0_u7_u1_U29 (.A( u0_u7_u1_n131 ) , .ZN( u0_u7_u1_n180 ) );
  INV_X1 u0_u7_u1_U3 (.A( u0_u7_u1_n159 ) , .ZN( u0_u7_u1_n182 ) );
  OAI221_X1 u0_u7_u1_U30 (.A( u0_u7_u1_n119 ) , .C2( u0_u7_u1_n129 ) , .ZN( u0_u7_u1_n138 ) , .B2( u0_u7_u1_n152 ) , .C1( u0_u7_u1_n174 ) , .B1( u0_u7_u1_n187 ) );
  INV_X1 u0_u7_u1_U31 (.A( u0_u7_u1_n148 ) , .ZN( u0_u7_u1_n187 ) );
  AOI211_X1 u0_u7_u1_U32 (.B( u0_u7_u1_n117 ) , .A( u0_u7_u1_n118 ) , .ZN( u0_u7_u1_n119 ) , .C2( u0_u7_u1_n146 ) , .C1( u0_u7_u1_n159 ) );
  NOR2_X1 u0_u7_u1_U33 (.A1( u0_u7_u1_n168 ) , .A2( u0_u7_u1_n176 ) , .ZN( u0_u7_u1_n98 ) );
  AOI211_X1 u0_u7_u1_U34 (.B( u0_u7_u1_n162 ) , .A( u0_u7_u1_n163 ) , .C2( u0_u7_u1_n164 ) , .ZN( u0_u7_u1_n165 ) , .C1( u0_u7_u1_n171 ) );
  AOI21_X1 u0_u7_u1_U35 (.A( u0_u7_u1_n160 ) , .B2( u0_u7_u1_n161 ) , .ZN( u0_u7_u1_n162 ) , .B1( u0_u7_u1_n182 ) );
  OR2_X1 u0_u7_u1_U36 (.A2( u0_u7_u1_n157 ) , .A1( u0_u7_u1_n158 ) , .ZN( u0_u7_u1_n163 ) );
  NAND2_X1 u0_u7_u1_U37 (.A1( u0_u7_u1_n128 ) , .ZN( u0_u7_u1_n146 ) , .A2( u0_u7_u1_n160 ) );
  NAND2_X1 u0_u7_u1_U38 (.A2( u0_u7_u1_n112 ) , .ZN( u0_u7_u1_n139 ) , .A1( u0_u7_u1_n152 ) );
  NAND2_X1 u0_u7_u1_U39 (.A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n156 ) , .A2( u0_u7_u1_n99 ) );
  AOI221_X1 u0_u7_u1_U4 (.A( u0_u7_u1_n138 ) , .C2( u0_u7_u1_n139 ) , .C1( u0_u7_u1_n140 ) , .B2( u0_u7_u1_n141 ) , .ZN( u0_u7_u1_n142 ) , .B1( u0_u7_u1_n175 ) );
  AOI221_X1 u0_u7_u1_U40 (.B1( u0_u7_u1_n140 ) , .ZN( u0_u7_u1_n167 ) , .B2( u0_u7_u1_n172 ) , .C2( u0_u7_u1_n175 ) , .C1( u0_u7_u1_n178 ) , .A( u0_u7_u1_n188 ) );
  INV_X1 u0_u7_u1_U41 (.ZN( u0_u7_u1_n188 ) , .A( u0_u7_u1_n97 ) );
  AOI211_X1 u0_u7_u1_U42 (.A( u0_u7_u1_n118 ) , .C1( u0_u7_u1_n132 ) , .C2( u0_u7_u1_n139 ) , .B( u0_u7_u1_n96 ) , .ZN( u0_u7_u1_n97 ) );
  AOI21_X1 u0_u7_u1_U43 (.B2( u0_u7_u1_n121 ) , .B1( u0_u7_u1_n135 ) , .A( u0_u7_u1_n152 ) , .ZN( u0_u7_u1_n96 ) );
  NOR2_X1 u0_u7_u1_U44 (.ZN( u0_u7_u1_n117 ) , .A1( u0_u7_u1_n121 ) , .A2( u0_u7_u1_n160 ) );
  OAI21_X1 u0_u7_u1_U45 (.B2( u0_u7_u1_n123 ) , .ZN( u0_u7_u1_n145 ) , .B1( u0_u7_u1_n160 ) , .A( u0_u7_u1_n185 ) );
  INV_X1 u0_u7_u1_U46 (.A( u0_u7_u1_n122 ) , .ZN( u0_u7_u1_n185 ) );
  AOI21_X1 u0_u7_u1_U47 (.B2( u0_u7_u1_n120 ) , .B1( u0_u7_u1_n121 ) , .ZN( u0_u7_u1_n122 ) , .A( u0_u7_u1_n128 ) );
  AOI21_X1 u0_u7_u1_U48 (.A( u0_u7_u1_n128 ) , .B2( u0_u7_u1_n129 ) , .ZN( u0_u7_u1_n130 ) , .B1( u0_u7_u1_n150 ) );
  NAND2_X1 u0_u7_u1_U49 (.ZN( u0_u7_u1_n112 ) , .A1( u0_u7_u1_n169 ) , .A2( u0_u7_u1_n170 ) );
  AOI211_X1 u0_u7_u1_U5 (.ZN( u0_u7_u1_n124 ) , .A( u0_u7_u1_n138 ) , .C2( u0_u7_u1_n139 ) , .B( u0_u7_u1_n145 ) , .C1( u0_u7_u1_n147 ) );
  NAND2_X1 u0_u7_u1_U50 (.ZN( u0_u7_u1_n129 ) , .A2( u0_u7_u1_n95 ) , .A1( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U51 (.A1( u0_u7_u1_n102 ) , .ZN( u0_u7_u1_n154 ) , .A2( u0_u7_u1_n99 ) );
  NAND2_X1 u0_u7_u1_U52 (.A2( u0_u7_u1_n100 ) , .ZN( u0_u7_u1_n135 ) , .A1( u0_u7_u1_n99 ) );
  AOI21_X1 u0_u7_u1_U53 (.A( u0_u7_u1_n152 ) , .B2( u0_u7_u1_n153 ) , .B1( u0_u7_u1_n154 ) , .ZN( u0_u7_u1_n158 ) );
  INV_X1 u0_u7_u1_U54 (.A( u0_u7_u1_n160 ) , .ZN( u0_u7_u1_n175 ) );
  NAND2_X1 u0_u7_u1_U55 (.A1( u0_u7_u1_n100 ) , .ZN( u0_u7_u1_n116 ) , .A2( u0_u7_u1_n95 ) );
  NAND2_X1 u0_u7_u1_U56 (.A1( u0_u7_u1_n102 ) , .ZN( u0_u7_u1_n131 ) , .A2( u0_u7_u1_n95 ) );
  NAND2_X1 u0_u7_u1_U57 (.A2( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n121 ) , .A1( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U58 (.A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n153 ) , .A2( u0_u7_u1_n98 ) );
  NAND2_X1 u0_u7_u1_U59 (.A2( u0_u7_u1_n104 ) , .A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n133 ) );
  AOI22_X1 u0_u7_u1_U6 (.B2( u0_u7_u1_n113 ) , .A2( u0_u7_u1_n114 ) , .ZN( u0_u7_u1_n125 ) , .A1( u0_u7_u1_n171 ) , .B1( u0_u7_u1_n173 ) );
  NAND2_X1 u0_u7_u1_U60 (.ZN( u0_u7_u1_n150 ) , .A2( u0_u7_u1_n98 ) , .A1( u0_u7_u1_n99 ) );
  NAND2_X1 u0_u7_u1_U61 (.A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n155 ) , .A2( u0_u7_u1_n95 ) );
  OAI21_X1 u0_u7_u1_U62 (.ZN( u0_u7_u1_n109 ) , .B1( u0_u7_u1_n129 ) , .B2( u0_u7_u1_n160 ) , .A( u0_u7_u1_n167 ) );
  NAND2_X1 u0_u7_u1_U63 (.A2( u0_u7_u1_n100 ) , .A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n120 ) );
  NAND2_X1 u0_u7_u1_U64 (.A1( u0_u7_u1_n102 ) , .A2( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n115 ) );
  NAND2_X1 u0_u7_u1_U65 (.A2( u0_u7_u1_n100 ) , .A1( u0_u7_u1_n104 ) , .ZN( u0_u7_u1_n151 ) );
  NAND2_X1 u0_u7_u1_U66 (.A2( u0_u7_u1_n103 ) , .A1( u0_u7_u1_n105 ) , .ZN( u0_u7_u1_n161 ) );
  INV_X1 u0_u7_u1_U67 (.A( u0_u7_u1_n152 ) , .ZN( u0_u7_u1_n173 ) );
  INV_X1 u0_u7_u1_U68 (.A( u0_u7_u1_n128 ) , .ZN( u0_u7_u1_n172 ) );
  NAND2_X1 u0_u7_u1_U69 (.A2( u0_u7_u1_n102 ) , .A1( u0_u7_u1_n103 ) , .ZN( u0_u7_u1_n123 ) );
  NAND2_X1 u0_u7_u1_U7 (.ZN( u0_u7_u1_n114 ) , .A1( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n156 ) );
  NOR2_X1 u0_u7_u1_U70 (.A2( u0_u7_X_7 ) , .A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n95 ) );
  NOR2_X1 u0_u7_u1_U71 (.A1( u0_u7_X_12 ) , .A2( u0_u7_X_9 ) , .ZN( u0_u7_u1_n100 ) );
  NOR2_X1 u0_u7_u1_U72 (.A2( u0_u7_X_8 ) , .A1( u0_u7_u1_n177 ) , .ZN( u0_u7_u1_n99 ) );
  NOR2_X1 u0_u7_u1_U73 (.A2( u0_u7_X_12 ) , .ZN( u0_u7_u1_n102 ) , .A1( u0_u7_u1_n176 ) );
  NOR2_X1 u0_u7_u1_U74 (.A2( u0_u7_X_9 ) , .ZN( u0_u7_u1_n105 ) , .A1( u0_u7_u1_n168 ) );
  NAND2_X1 u0_u7_u1_U75 (.A1( u0_u7_X_10 ) , .ZN( u0_u7_u1_n160 ) , .A2( u0_u7_u1_n169 ) );
  NAND2_X1 u0_u7_u1_U76 (.A2( u0_u7_X_10 ) , .A1( u0_u7_X_11 ) , .ZN( u0_u7_u1_n152 ) );
  NAND2_X1 u0_u7_u1_U77 (.A1( u0_u7_X_11 ) , .ZN( u0_u7_u1_n128 ) , .A2( u0_u7_u1_n170 ) );
  AND2_X1 u0_u7_u1_U78 (.A2( u0_u7_X_7 ) , .A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n104 ) );
  AND2_X1 u0_u7_u1_U79 (.A1( u0_u7_X_8 ) , .ZN( u0_u7_u1_n103 ) , .A2( u0_u7_u1_n177 ) );
  NOR2_X1 u0_u7_u1_U8 (.A1( u0_u7_u1_n112 ) , .A2( u0_u7_u1_n116 ) , .ZN( u0_u7_u1_n118 ) );
  INV_X1 u0_u7_u1_U80 (.A( u0_u7_X_10 ) , .ZN( u0_u7_u1_n170 ) );
  INV_X1 u0_u7_u1_U81 (.A( u0_u7_X_9 ) , .ZN( u0_u7_u1_n176 ) );
  INV_X1 u0_u7_u1_U82 (.A( u0_u7_X_11 ) , .ZN( u0_u7_u1_n169 ) );
  INV_X1 u0_u7_u1_U83 (.A( u0_u7_X_12 ) , .ZN( u0_u7_u1_n168 ) );
  INV_X1 u0_u7_u1_U84 (.A( u0_u7_X_7 ) , .ZN( u0_u7_u1_n177 ) );
  NAND4_X1 u0_u7_u1_U85 (.ZN( u0_out7_28 ) , .A4( u0_u7_u1_n124 ) , .A3( u0_u7_u1_n125 ) , .A2( u0_u7_u1_n126 ) , .A1( u0_u7_u1_n127 ) );
  OAI21_X1 u0_u7_u1_U86 (.ZN( u0_u7_u1_n127 ) , .B2( u0_u7_u1_n139 ) , .B1( u0_u7_u1_n175 ) , .A( u0_u7_u1_n183 ) );
  OAI21_X1 u0_u7_u1_U87 (.ZN( u0_u7_u1_n126 ) , .B2( u0_u7_u1_n140 ) , .A( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n178 ) );
  NAND4_X1 u0_u7_u1_U88 (.ZN( u0_out7_18 ) , .A4( u0_u7_u1_n165 ) , .A3( u0_u7_u1_n166 ) , .A1( u0_u7_u1_n167 ) , .A2( u0_u7_u1_n186 ) );
  AOI22_X1 u0_u7_u1_U89 (.B2( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n147 ) , .A2( u0_u7_u1_n148 ) , .ZN( u0_u7_u1_n166 ) , .A1( u0_u7_u1_n172 ) );
  OAI21_X1 u0_u7_u1_U9 (.ZN( u0_u7_u1_n101 ) , .B1( u0_u7_u1_n141 ) , .A( u0_u7_u1_n146 ) , .B2( u0_u7_u1_n183 ) );
  INV_X1 u0_u7_u1_U90 (.A( u0_u7_u1_n145 ) , .ZN( u0_u7_u1_n186 ) );
  NAND4_X1 u0_u7_u1_U91 (.ZN( u0_out7_2 ) , .A4( u0_u7_u1_n142 ) , .A3( u0_u7_u1_n143 ) , .A2( u0_u7_u1_n144 ) , .A1( u0_u7_u1_n179 ) );
  OAI21_X1 u0_u7_u1_U92 (.B2( u0_u7_u1_n132 ) , .ZN( u0_u7_u1_n144 ) , .A( u0_u7_u1_n146 ) , .B1( u0_u7_u1_n180 ) );
  INV_X1 u0_u7_u1_U93 (.A( u0_u7_u1_n130 ) , .ZN( u0_u7_u1_n179 ) );
  OR4_X1 u0_u7_u1_U94 (.ZN( u0_out7_13 ) , .A4( u0_u7_u1_n108 ) , .A3( u0_u7_u1_n109 ) , .A2( u0_u7_u1_n110 ) , .A1( u0_u7_u1_n111 ) );
  AOI21_X1 u0_u7_u1_U95 (.ZN( u0_u7_u1_n111 ) , .A( u0_u7_u1_n128 ) , .B2( u0_u7_u1_n131 ) , .B1( u0_u7_u1_n135 ) );
  AOI21_X1 u0_u7_u1_U96 (.ZN( u0_u7_u1_n110 ) , .A( u0_u7_u1_n116 ) , .B1( u0_u7_u1_n152 ) , .B2( u0_u7_u1_n160 ) );
  NAND3_X1 u0_u7_u1_U97 (.A3( u0_u7_u1_n149 ) , .A2( u0_u7_u1_n150 ) , .A1( u0_u7_u1_n151 ) , .ZN( u0_u7_u1_n164 ) );
  NAND3_X1 u0_u7_u1_U98 (.A3( u0_u7_u1_n134 ) , .A2( u0_u7_u1_n135 ) , .ZN( u0_u7_u1_n136 ) , .A1( u0_u7_u1_n151 ) );
  NAND3_X1 u0_u7_u1_U99 (.A1( u0_u7_u1_n133 ) , .ZN( u0_u7_u1_n137 ) , .A2( u0_u7_u1_n154 ) , .A3( u0_u7_u1_n181 ) );
  OAI21_X1 u0_uk_U1002 (.ZN( u0_K8_4 ) , .B2( u0_uk_n351 ) , .A( u0_uk_n743 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U1003 (.A1( u0_uk_K_r6_19 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n743 ) );
  OAI21_X1 u0_uk_U1058 (.ZN( u0_K4_38 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n505 ) , .A( u0_uk_n825 ) );
  NAND2_X1 u0_uk_U1059 (.A1( u0_uk_K_r2_50 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n825 ) );
  INV_X1 u0_uk_U1113 (.ZN( u0_K8_12 ) , .A( u0_uk_n761 ) );
  AOI22_X1 u0_uk_U1114 (.B2( u0_uk_K_r6_3 ) , .A2( u0_uk_K_r6_53 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n761 ) );
  INV_X1 u0_uk_U1156 (.ZN( u0_K6_2 ) , .A( u0_uk_n793 ) );
  INV_X1 u0_uk_U1158 (.ZN( u0_K8_3 ) , .A( u0_uk_n749 ) );
  OAI22_X1 u0_uk_U123 (.ZN( u0_K4_47 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n499 ) , .B2( u0_uk_n508 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U186 (.ZN( u0_K6_14 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n442 ) , .A2( u0_uk_n448 ) );
  OAI22_X1 u0_uk_U272 (.ZN( u0_K4_44 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .A2( u0_uk_n521 ) , .B2( u0_uk_n538 ) );
  OAI22_X1 u0_uk_U277 (.ZN( u0_K16_6 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n639 ) , .B2( u0_uk_n644 ) );
  OAI22_X1 u0_uk_U279 (.ZN( u0_K6_6 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n410 ) , .B2( u0_uk_n414 ) , .B1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U280 (.ZN( u0_K6_8 ) , .B2( u0_uk_n442 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n786 ) );
  OAI22_X1 u0_uk_U287 (.ZN( u0_K8_8 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n324 ) , .B2( u0_uk_n330 ) );
  OAI22_X1 u0_uk_U326 (.ZN( u0_K4_46 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n514 ) , .B2( u0_uk_n528 ) );
  INV_X1 u0_uk_U341 (.ZN( u0_K6_4 ) , .A( u0_uk_n788 ) );
  AOI22_X1 u0_uk_U342 (.B2( u0_uk_K_r4_41 ) , .A2( u0_uk_K_r4_47 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n788 ) );
  OAI22_X1 u0_uk_U365 (.ZN( u0_K4_40 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n506 ) , .B2( u0_uk_n516 ) );
  OAI22_X1 u0_uk_U409 (.ZN( u0_K8_9 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n162 ) , .B2( u0_uk_n350 ) , .A2( u0_uk_n356 ) );
  OAI22_X1 u0_uk_U429 (.ZN( u0_K16_9 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n630 ) , .B2( u0_uk_n637 ) );
  OAI22_X1 u0_uk_U463 (.ZN( u0_K4_37 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n251 ) , .A2( u0_uk_n513 ) , .B2( u0_uk_n527 ) );
  INV_X1 u0_uk_U464 (.ZN( u0_K6_9 ) , .A( u0_uk_n785 ) );
  OAI21_X1 u0_uk_U493 (.ZN( u0_K8_2 ) , .B2( u0_uk_n343 ) , .A( u0_uk_n754 ) , .B1( u0_uk_n83 ) );
  NAND2_X1 u0_uk_U494 (.A1( u0_uk_K_r6_27 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n754 ) );
  OAI21_X1 u0_uk_U532 (.ZN( u0_K16_12 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n660 ) , .A( u0_uk_n910 ) );
  NAND2_X1 u0_uk_U533 (.A1( u0_uk_K_r14_12 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n910 ) );
  INV_X1 u0_uk_U542 (.ZN( u0_K6_17 ) , .A( u0_uk_n800 ) );
  AOI22_X1 u0_uk_U543 (.B2( u0_uk_K_r4_4 ) , .A2( u0_uk_K_r4_55 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n800 ) );
  OAI22_X1 u0_uk_U571 (.ZN( u0_K16_10 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n636 ) , .B2( u0_uk_n639 ) );
  OAI22_X1 u0_uk_U581 (.ZN( u0_K8_10 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n337 ) , .B2( u0_uk_n339 ) );
  INV_X1 u0_uk_U582 (.ZN( u0_K6_10 ) , .A( u0_uk_n801 ) );
  AOI22_X1 u0_uk_U583 (.B2( u0_uk_K_r4_3 ) , .A2( u0_uk_K_r4_54 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n801 ) );
  OAI21_X1 u0_uk_U622 (.ZN( u0_K16_11 ) , .B1( u0_uk_n146 ) , .B2( u0_uk_n646 ) , .A( u0_uk_n911 ) );
  NAND2_X1 u0_uk_U623 (.A1( u0_uk_K_r14_39 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n911 ) );
  INV_X1 u0_uk_U649 (.A( u0_key_r_44 ) , .ZN( u0_uk_n680 ) );
  OAI22_X1 u0_uk_U677 (.ZN( u0_K16_3 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n652 ) , .B2( u0_uk_n660 ) );
  OAI22_X1 u0_uk_U685 (.ZN( u0_K16_7 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n651 ) , .B2( u0_uk_n659 ) );
  OAI21_X1 u0_uk_U699 (.ZN( u0_K6_7 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n423 ) , .A( u0_uk_n787 ) );
  NAND2_X1 u0_uk_U700 (.A1( u0_uk_K_r4_33 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n787 ) );
  OAI22_X1 u0_uk_U733 (.ZN( u0_K4_42 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n521 ) , .B2( u0_uk_n528 ) );
  OAI22_X1 u0_uk_U798 (.ZN( u0_K16_1 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n637 ) , .B2( u0_uk_n640 ) );
  OAI22_X1 u0_uk_U799 (.ZN( u0_K6_1 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n410 ) , .B2( u0_uk_n426 ) );
  INV_X1 u0_uk_U827 (.ZN( u0_K6_18 ) , .A( u0_uk_n799 ) );
  AOI22_X1 u0_uk_U846 (.B2( u0_uk_K_r6_10 ) , .A2( u0_uk_K_r6_3 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n749 ) );
  OAI21_X1 u0_uk_U860 (.ZN( u0_K16_2 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n668 ) , .A( u0_uk_n903 ) );
  NAND2_X1 u0_uk_U861 (.A1( u0_uk_K_r14_11 ) , .A2( u0_uk_n118 ) , .ZN( u0_uk_n903 ) );
  OAI22_X1 u0_uk_U879 (.ZN( u0_K8_5 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n318 ) , .B2( u0_uk_n324 ) );
  OAI22_X1 u0_uk_U880 (.ZN( u0_K6_5 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n432 ) , .B2( u0_uk_n436 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U891 (.ZN( u0_K8_6 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n339 ) , .B2( u0_uk_n344 ) );
  OAI22_X1 u0_uk_U897 (.ZN( u0_K6_12 ) , .A1( u0_uk_n257 ) , .B2( u0_uk_n432 ) , .A2( u0_uk_n448 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U91 (.ZN( u0_K4_41 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n522 ) , .B2( u0_uk_n539 ) );
  OAI22_X1 u0_uk_U925 (.ZN( u0_K4_39 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n516 ) , .B2( u0_uk_n537 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U94 (.ZN( u0_K16_5 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n187 ) , .B2( u0_uk_n664 ) , .A2( u0_uk_n667 ) );
  OAI22_X1 u0_uk_U978 (.ZN( u0_K4_45 ) , .B1( u0_uk_n163 ) , .A1( u0_uk_n27 ) , .A2( u0_uk_n498 ) , .B2( u0_uk_n537 ) );
  OAI22_X1 u0_uk_U981 (.ZN( u0_K6_3 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n427 ) , .B2( u0_uk_n441 ) );
  OAI22_X1 u0_uk_U983 (.ZN( u0_K8_7 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n257 ) , .B2( u0_uk_n352 ) , .A2( u0_uk_n358 ) );
  OAI22_X1 u0_uk_U987 (.ZN( u0_K6_15 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n423 ) , .B2( u0_uk_n435 ) );
  XOR2_X1 u1_U192 (.B( u1_L0_5 ) , .Z( u1_N36 ) , .A( u1_out1_5 ) );
  XOR2_X1 u1_U350 (.B( u1_L5_26 ) , .Z( u1_N217 ) , .A( u1_out6_26 ) );
  XOR2_X1 u1_U356 (.B( u1_L5_20 ) , .Z( u1_N211 ) , .A( u1_out6_20 ) );
  XOR2_X1 u1_U367 (.B( u1_L5_10 ) , .Z( u1_N201 ) , .A( u1_out6_10 ) );
  XOR2_X1 u1_U378 (.B( u1_L5_1 ) , .Z( u1_N192 ) , .A( u1_out6_1 ) );
  XOR2_X1 u1_U48 (.B( u1_L0_27 ) , .Z( u1_N58 ) , .A( u1_out1_27 ) );
  XOR2_X1 u1_U54 (.B( u1_L0_21 ) , .Z( u1_N52 ) , .A( u1_out1_21 ) );
  XOR2_X1 u1_U81 (.B( u1_L0_15 ) , .Z( u1_N46 ) , .A( u1_out1_15 ) );
  XOR2_X1 u1_u1_U10 (.B( u1_K2_45 ) , .A( u1_R0_30 ) , .Z( u1_u1_X_45 ) );
  XOR2_X1 u1_u1_U11 (.B( u1_K2_44 ) , .A( u1_R0_29 ) , .Z( u1_u1_X_44 ) );
  XOR2_X1 u1_u1_U12 (.B( u1_K2_43 ) , .A( u1_R0_28 ) , .Z( u1_u1_X_43 ) );
  XOR2_X1 u1_u1_U7 (.B( u1_K2_48 ) , .A( u1_R0_1 ) , .Z( u1_u1_X_48 ) );
  XOR2_X1 u1_u1_U8 (.B( u1_K2_47 ) , .A( u1_R0_32 ) , .Z( u1_u1_X_47 ) );
  XOR2_X1 u1_u1_U9 (.B( u1_K2_46 ) , .A( u1_R0_31 ) , .Z( u1_u1_X_46 ) );
  AND3_X1 u1_u1_u7_U10 (.A3( u1_u1_u7_n110 ) , .A2( u1_u1_u7_n127 ) , .A1( u1_u1_u7_n132 ) , .ZN( u1_u1_u7_n92 ) );
  OAI21_X1 u1_u1_u7_U11 (.A( u1_u1_u7_n161 ) , .B1( u1_u1_u7_n168 ) , .B2( u1_u1_u7_n173 ) , .ZN( u1_u1_u7_n91 ) );
  AOI211_X1 u1_u1_u7_U12 (.A( u1_u1_u7_n117 ) , .ZN( u1_u1_u7_n118 ) , .C2( u1_u1_u7_n126 ) , .C1( u1_u1_u7_n177 ) , .B( u1_u1_u7_n180 ) );
  OAI22_X1 u1_u1_u7_U13 (.B1( u1_u1_u7_n115 ) , .ZN( u1_u1_u7_n117 ) , .A2( u1_u1_u7_n133 ) , .A1( u1_u1_u7_n137 ) , .B2( u1_u1_u7_n162 ) );
  INV_X1 u1_u1_u7_U14 (.A( u1_u1_u7_n116 ) , .ZN( u1_u1_u7_n180 ) );
  NOR3_X1 u1_u1_u7_U15 (.ZN( u1_u1_u7_n115 ) , .A3( u1_u1_u7_n145 ) , .A2( u1_u1_u7_n168 ) , .A1( u1_u1_u7_n169 ) );
  OAI211_X1 u1_u1_u7_U16 (.B( u1_u1_u7_n122 ) , .A( u1_u1_u7_n123 ) , .C2( u1_u1_u7_n124 ) , .ZN( u1_u1_u7_n154 ) , .C1( u1_u1_u7_n162 ) );
  AOI222_X1 u1_u1_u7_U17 (.ZN( u1_u1_u7_n122 ) , .C2( u1_u1_u7_n126 ) , .C1( u1_u1_u7_n145 ) , .B1( u1_u1_u7_n161 ) , .A2( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n170 ) , .A1( u1_u1_u7_n176 ) );
  INV_X1 u1_u1_u7_U18 (.A( u1_u1_u7_n133 ) , .ZN( u1_u1_u7_n176 ) );
  NOR3_X1 u1_u1_u7_U19 (.A2( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n135 ) , .ZN( u1_u1_u7_n136 ) , .A3( u1_u1_u7_n171 ) );
  NOR2_X1 u1_u1_u7_U20 (.A1( u1_u1_u7_n130 ) , .A2( u1_u1_u7_n134 ) , .ZN( u1_u1_u7_n153 ) );
  INV_X1 u1_u1_u7_U21 (.A( u1_u1_u7_n101 ) , .ZN( u1_u1_u7_n165 ) );
  NOR2_X1 u1_u1_u7_U22 (.ZN( u1_u1_u7_n111 ) , .A2( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n169 ) );
  AOI21_X1 u1_u1_u7_U23 (.ZN( u1_u1_u7_n104 ) , .B2( u1_u1_u7_n112 ) , .B1( u1_u1_u7_n127 ) , .A( u1_u1_u7_n164 ) );
  AOI21_X1 u1_u1_u7_U24 (.ZN( u1_u1_u7_n106 ) , .B1( u1_u1_u7_n133 ) , .B2( u1_u1_u7_n146 ) , .A( u1_u1_u7_n162 ) );
  AOI21_X1 u1_u1_u7_U25 (.A( u1_u1_u7_n101 ) , .ZN( u1_u1_u7_n107 ) , .B2( u1_u1_u7_n128 ) , .B1( u1_u1_u7_n175 ) );
  INV_X1 u1_u1_u7_U26 (.A( u1_u1_u7_n138 ) , .ZN( u1_u1_u7_n171 ) );
  INV_X1 u1_u1_u7_U27 (.A( u1_u1_u7_n131 ) , .ZN( u1_u1_u7_n177 ) );
  INV_X1 u1_u1_u7_U28 (.A( u1_u1_u7_n110 ) , .ZN( u1_u1_u7_n174 ) );
  NAND2_X1 u1_u1_u7_U29 (.A1( u1_u1_u7_n129 ) , .A2( u1_u1_u7_n132 ) , .ZN( u1_u1_u7_n149 ) );
  OAI21_X1 u1_u1_u7_U3 (.ZN( u1_u1_u7_n159 ) , .A( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n171 ) , .B1( u1_u1_u7_n174 ) );
  NAND2_X1 u1_u1_u7_U30 (.A1( u1_u1_u7_n113 ) , .A2( u1_u1_u7_n124 ) , .ZN( u1_u1_u7_n130 ) );
  INV_X1 u1_u1_u7_U31 (.A( u1_u1_u7_n112 ) , .ZN( u1_u1_u7_n173 ) );
  INV_X1 u1_u1_u7_U32 (.A( u1_u1_u7_n128 ) , .ZN( u1_u1_u7_n168 ) );
  INV_X1 u1_u1_u7_U33 (.A( u1_u1_u7_n148 ) , .ZN( u1_u1_u7_n169 ) );
  INV_X1 u1_u1_u7_U34 (.A( u1_u1_u7_n127 ) , .ZN( u1_u1_u7_n179 ) );
  NOR2_X1 u1_u1_u7_U35 (.ZN( u1_u1_u7_n101 ) , .A2( u1_u1_u7_n150 ) , .A1( u1_u1_u7_n156 ) );
  AOI211_X1 u1_u1_u7_U36 (.B( u1_u1_u7_n154 ) , .A( u1_u1_u7_n155 ) , .C1( u1_u1_u7_n156 ) , .ZN( u1_u1_u7_n157 ) , .C2( u1_u1_u7_n172 ) );
  INV_X1 u1_u1_u7_U37 (.A( u1_u1_u7_n153 ) , .ZN( u1_u1_u7_n172 ) );
  AOI211_X1 u1_u1_u7_U38 (.B( u1_u1_u7_n139 ) , .A( u1_u1_u7_n140 ) , .C2( u1_u1_u7_n141 ) , .ZN( u1_u1_u7_n142 ) , .C1( u1_u1_u7_n156 ) );
  NAND4_X1 u1_u1_u7_U39 (.A3( u1_u1_u7_n127 ) , .A2( u1_u1_u7_n128 ) , .A1( u1_u1_u7_n129 ) , .ZN( u1_u1_u7_n141 ) , .A4( u1_u1_u7_n147 ) );
  INV_X1 u1_u1_u7_U4 (.A( u1_u1_u7_n111 ) , .ZN( u1_u1_u7_n170 ) );
  AOI21_X1 u1_u1_u7_U40 (.A( u1_u1_u7_n137 ) , .B1( u1_u1_u7_n138 ) , .ZN( u1_u1_u7_n139 ) , .B2( u1_u1_u7_n146 ) );
  OAI22_X1 u1_u1_u7_U41 (.B1( u1_u1_u7_n136 ) , .ZN( u1_u1_u7_n140 ) , .A1( u1_u1_u7_n153 ) , .B2( u1_u1_u7_n162 ) , .A2( u1_u1_u7_n164 ) );
  AOI21_X1 u1_u1_u7_U42 (.ZN( u1_u1_u7_n123 ) , .B1( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n177 ) , .A( u1_u1_u7_n97 ) );
  AOI21_X1 u1_u1_u7_U43 (.B2( u1_u1_u7_n113 ) , .B1( u1_u1_u7_n124 ) , .A( u1_u1_u7_n125 ) , .ZN( u1_u1_u7_n97 ) );
  INV_X1 u1_u1_u7_U44 (.A( u1_u1_u7_n125 ) , .ZN( u1_u1_u7_n161 ) );
  INV_X1 u1_u1_u7_U45 (.A( u1_u1_u7_n152 ) , .ZN( u1_u1_u7_n162 ) );
  AOI22_X1 u1_u1_u7_U46 (.A2( u1_u1_u7_n114 ) , .ZN( u1_u1_u7_n119 ) , .B1( u1_u1_u7_n130 ) , .A1( u1_u1_u7_n156 ) , .B2( u1_u1_u7_n165 ) );
  NAND2_X1 u1_u1_u7_U47 (.A2( u1_u1_u7_n112 ) , .ZN( u1_u1_u7_n114 ) , .A1( u1_u1_u7_n175 ) );
  AND2_X1 u1_u1_u7_U48 (.ZN( u1_u1_u7_n145 ) , .A2( u1_u1_u7_n98 ) , .A1( u1_u1_u7_n99 ) );
  NOR2_X1 u1_u1_u7_U49 (.ZN( u1_u1_u7_n137 ) , .A1( u1_u1_u7_n150 ) , .A2( u1_u1_u7_n161 ) );
  INV_X1 u1_u1_u7_U5 (.A( u1_u1_u7_n149 ) , .ZN( u1_u1_u7_n175 ) );
  AOI21_X1 u1_u1_u7_U50 (.ZN( u1_u1_u7_n105 ) , .B2( u1_u1_u7_n110 ) , .A( u1_u1_u7_n125 ) , .B1( u1_u1_u7_n147 ) );
  NAND2_X1 u1_u1_u7_U51 (.ZN( u1_u1_u7_n146 ) , .A1( u1_u1_u7_n95 ) , .A2( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U52 (.A2( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n147 ) , .A1( u1_u1_u7_n93 ) );
  NAND2_X1 u1_u1_u7_U53 (.A1( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n127 ) , .A2( u1_u1_u7_n99 ) );
  OR2_X1 u1_u1_u7_U54 (.ZN( u1_u1_u7_n126 ) , .A2( u1_u1_u7_n152 ) , .A1( u1_u1_u7_n156 ) );
  NAND2_X1 u1_u1_u7_U55 (.A2( u1_u1_u7_n102 ) , .A1( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n133 ) );
  NAND2_X1 u1_u1_u7_U56 (.ZN( u1_u1_u7_n112 ) , .A2( u1_u1_u7_n96 ) , .A1( u1_u1_u7_n99 ) );
  NAND2_X1 u1_u1_u7_U57 (.A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n128 ) , .A1( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U58 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n113 ) , .A2( u1_u1_u7_n93 ) );
  NAND2_X1 u1_u1_u7_U59 (.A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n124 ) , .A1( u1_u1_u7_n96 ) );
  INV_X1 u1_u1_u7_U6 (.A( u1_u1_u7_n154 ) , .ZN( u1_u1_u7_n178 ) );
  NAND2_X1 u1_u1_u7_U60 (.ZN( u1_u1_u7_n110 ) , .A1( u1_u1_u7_n95 ) , .A2( u1_u1_u7_n96 ) );
  INV_X1 u1_u1_u7_U61 (.A( u1_u1_u7_n150 ) , .ZN( u1_u1_u7_n164 ) );
  AND2_X1 u1_u1_u7_U62 (.ZN( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n93 ) , .A2( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U63 (.A1( u1_u1_u7_n100 ) , .A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n129 ) );
  NAND2_X1 u1_u1_u7_U64 (.A2( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n131 ) , .A1( u1_u1_u7_n95 ) );
  NAND2_X1 u1_u1_u7_U65 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n138 ) , .A2( u1_u1_u7_n99 ) );
  NAND2_X1 u1_u1_u7_U66 (.ZN( u1_u1_u7_n132 ) , .A1( u1_u1_u7_n93 ) , .A2( u1_u1_u7_n96 ) );
  NAND2_X1 u1_u1_u7_U67 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n148 ) , .A2( u1_u1_u7_n95 ) );
  NOR2_X1 u1_u1_u7_U68 (.A2( u1_u1_X_47 ) , .ZN( u1_u1_u7_n150 ) , .A1( u1_u1_u7_n163 ) );
  NOR2_X1 u1_u1_u7_U69 (.A2( u1_u1_X_43 ) , .A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n103 ) );
  AOI211_X1 u1_u1_u7_U7 (.ZN( u1_u1_u7_n116 ) , .A( u1_u1_u7_n155 ) , .C1( u1_u1_u7_n161 ) , .C2( u1_u1_u7_n171 ) , .B( u1_u1_u7_n94 ) );
  NOR2_X1 u1_u1_u7_U70 (.A2( u1_u1_X_48 ) , .A1( u1_u1_u7_n166 ) , .ZN( u1_u1_u7_n95 ) );
  NOR2_X1 u1_u1_u7_U71 (.A2( u1_u1_X_45 ) , .A1( u1_u1_X_48 ) , .ZN( u1_u1_u7_n99 ) );
  NOR2_X1 u1_u1_u7_U72 (.A2( u1_u1_X_44 ) , .A1( u1_u1_u7_n167 ) , .ZN( u1_u1_u7_n98 ) );
  NOR2_X1 u1_u1_u7_U73 (.A2( u1_u1_X_46 ) , .A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n152 ) );
  AND2_X1 u1_u1_u7_U74 (.A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n156 ) , .A2( u1_u1_u7_n163 ) );
  NAND2_X1 u1_u1_u7_U75 (.A2( u1_u1_X_46 ) , .A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n125 ) );
  AND2_X1 u1_u1_u7_U76 (.A2( u1_u1_X_45 ) , .A1( u1_u1_X_48 ) , .ZN( u1_u1_u7_n102 ) );
  AND2_X1 u1_u1_u7_U77 (.A2( u1_u1_X_43 ) , .A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n96 ) );
  AND2_X1 u1_u1_u7_U78 (.A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n100 ) , .A2( u1_u1_u7_n167 ) );
  AND2_X1 u1_u1_u7_U79 (.A1( u1_u1_X_48 ) , .A2( u1_u1_u7_n166 ) , .ZN( u1_u1_u7_n93 ) );
  OAI222_X1 u1_u1_u7_U8 (.C2( u1_u1_u7_n101 ) , .B2( u1_u1_u7_n111 ) , .A1( u1_u1_u7_n113 ) , .C1( u1_u1_u7_n146 ) , .A2( u1_u1_u7_n162 ) , .B1( u1_u1_u7_n164 ) , .ZN( u1_u1_u7_n94 ) );
  INV_X1 u1_u1_u7_U80 (.A( u1_u1_X_46 ) , .ZN( u1_u1_u7_n163 ) );
  INV_X1 u1_u1_u7_U81 (.A( u1_u1_X_43 ) , .ZN( u1_u1_u7_n167 ) );
  INV_X1 u1_u1_u7_U82 (.A( u1_u1_X_45 ) , .ZN( u1_u1_u7_n166 ) );
  NAND4_X1 u1_u1_u7_U83 (.ZN( u1_out1_5 ) , .A4( u1_u1_u7_n108 ) , .A3( u1_u1_u7_n109 ) , .A1( u1_u1_u7_n116 ) , .A2( u1_u1_u7_n123 ) );
  AOI22_X1 u1_u1_u7_U84 (.ZN( u1_u1_u7_n109 ) , .A2( u1_u1_u7_n126 ) , .B2( u1_u1_u7_n145 ) , .B1( u1_u1_u7_n156 ) , .A1( u1_u1_u7_n171 ) );
  NOR4_X1 u1_u1_u7_U85 (.A4( u1_u1_u7_n104 ) , .A3( u1_u1_u7_n105 ) , .A2( u1_u1_u7_n106 ) , .A1( u1_u1_u7_n107 ) , .ZN( u1_u1_u7_n108 ) );
  NAND4_X1 u1_u1_u7_U86 (.ZN( u1_out1_27 ) , .A4( u1_u1_u7_n118 ) , .A3( u1_u1_u7_n119 ) , .A2( u1_u1_u7_n120 ) , .A1( u1_u1_u7_n121 ) );
  OAI21_X1 u1_u1_u7_U87 (.ZN( u1_u1_u7_n121 ) , .B2( u1_u1_u7_n145 ) , .A( u1_u1_u7_n150 ) , .B1( u1_u1_u7_n174 ) );
  OAI21_X1 u1_u1_u7_U88 (.ZN( u1_u1_u7_n120 ) , .A( u1_u1_u7_n161 ) , .B2( u1_u1_u7_n170 ) , .B1( u1_u1_u7_n179 ) );
  NAND4_X1 u1_u1_u7_U89 (.ZN( u1_out1_21 ) , .A4( u1_u1_u7_n157 ) , .A3( u1_u1_u7_n158 ) , .A2( u1_u1_u7_n159 ) , .A1( u1_u1_u7_n160 ) );
  OAI221_X1 u1_u1_u7_U9 (.C1( u1_u1_u7_n101 ) , .C2( u1_u1_u7_n147 ) , .ZN( u1_u1_u7_n155 ) , .B2( u1_u1_u7_n162 ) , .A( u1_u1_u7_n91 ) , .B1( u1_u1_u7_n92 ) );
  OAI21_X1 u1_u1_u7_U90 (.B1( u1_u1_u7_n145 ) , .ZN( u1_u1_u7_n160 ) , .A( u1_u1_u7_n161 ) , .B2( u1_u1_u7_n177 ) );
  AOI22_X1 u1_u1_u7_U91 (.B2( u1_u1_u7_n149 ) , .B1( u1_u1_u7_n150 ) , .A2( u1_u1_u7_n151 ) , .A1( u1_u1_u7_n152 ) , .ZN( u1_u1_u7_n158 ) );
  NAND4_X1 u1_u1_u7_U92 (.ZN( u1_out1_15 ) , .A4( u1_u1_u7_n142 ) , .A3( u1_u1_u7_n143 ) , .A2( u1_u1_u7_n144 ) , .A1( u1_u1_u7_n178 ) );
  OR2_X1 u1_u1_u7_U93 (.A2( u1_u1_u7_n125 ) , .A1( u1_u1_u7_n129 ) , .ZN( u1_u1_u7_n144 ) );
  AOI22_X1 u1_u1_u7_U94 (.A2( u1_u1_u7_n126 ) , .ZN( u1_u1_u7_n143 ) , .B2( u1_u1_u7_n165 ) , .B1( u1_u1_u7_n173 ) , .A1( u1_u1_u7_n174 ) );
  NAND3_X1 u1_u1_u7_U95 (.A3( u1_u1_u7_n146 ) , .A2( u1_u1_u7_n147 ) , .A1( u1_u1_u7_n148 ) , .ZN( u1_u1_u7_n151 ) );
  NAND3_X1 u1_u1_u7_U96 (.A3( u1_u1_u7_n131 ) , .A2( u1_u1_u7_n132 ) , .A1( u1_u1_u7_n133 ) , .ZN( u1_u1_u7_n135 ) );
  XOR2_X1 u1_u6_U33 (.B( u1_K7_24 ) , .A( u1_R5_17 ) , .Z( u1_u6_X_24 ) );
  XOR2_X1 u1_u6_U34 (.B( u1_K7_23 ) , .A( u1_R5_16 ) , .Z( u1_u6_X_23 ) );
  XOR2_X1 u1_u6_U35 (.B( u1_K7_22 ) , .A( u1_R5_15 ) , .Z( u1_u6_X_22 ) );
  XOR2_X1 u1_u6_U36 (.B( u1_K7_21 ) , .A( u1_R5_14 ) , .Z( u1_u6_X_21 ) );
  XOR2_X1 u1_u6_U37 (.B( u1_K7_20 ) , .A( u1_R5_13 ) , .Z( u1_u6_X_20 ) );
  XOR2_X1 u1_u6_U39 (.B( u1_K7_19 ) , .A( u1_R5_12 ) , .Z( u1_u6_X_19 ) );
  OAI22_X1 u1_u6_u3_U10 (.B1( u1_u6_u3_n113 ) , .A2( u1_u6_u3_n135 ) , .A1( u1_u6_u3_n150 ) , .B2( u1_u6_u3_n164 ) , .ZN( u1_u6_u3_n98 ) );
  OAI211_X1 u1_u6_u3_U11 (.B( u1_u6_u3_n106 ) , .ZN( u1_u6_u3_n119 ) , .C2( u1_u6_u3_n128 ) , .C1( u1_u6_u3_n167 ) , .A( u1_u6_u3_n181 ) );
  AOI221_X1 u1_u6_u3_U12 (.C1( u1_u6_u3_n105 ) , .ZN( u1_u6_u3_n106 ) , .A( u1_u6_u3_n131 ) , .B2( u1_u6_u3_n132 ) , .C2( u1_u6_u3_n133 ) , .B1( u1_u6_u3_n169 ) );
  INV_X1 u1_u6_u3_U13 (.ZN( u1_u6_u3_n181 ) , .A( u1_u6_u3_n98 ) );
  NAND2_X1 u1_u6_u3_U14 (.ZN( u1_u6_u3_n105 ) , .A2( u1_u6_u3_n130 ) , .A1( u1_u6_u3_n155 ) );
  AOI22_X1 u1_u6_u3_U15 (.B1( u1_u6_u3_n115 ) , .A2( u1_u6_u3_n116 ) , .ZN( u1_u6_u3_n123 ) , .B2( u1_u6_u3_n133 ) , .A1( u1_u6_u3_n169 ) );
  NAND2_X1 u1_u6_u3_U16 (.ZN( u1_u6_u3_n116 ) , .A2( u1_u6_u3_n151 ) , .A1( u1_u6_u3_n182 ) );
  NOR2_X1 u1_u6_u3_U17 (.ZN( u1_u6_u3_n126 ) , .A2( u1_u6_u3_n150 ) , .A1( u1_u6_u3_n164 ) );
  AOI21_X1 u1_u6_u3_U18 (.ZN( u1_u6_u3_n112 ) , .B2( u1_u6_u3_n146 ) , .B1( u1_u6_u3_n155 ) , .A( u1_u6_u3_n167 ) );
  NAND2_X1 u1_u6_u3_U19 (.A1( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n142 ) , .A2( u1_u6_u3_n164 ) );
  NAND2_X1 u1_u6_u3_U20 (.ZN( u1_u6_u3_n132 ) , .A2( u1_u6_u3_n152 ) , .A1( u1_u6_u3_n156 ) );
  AND2_X1 u1_u6_u3_U21 (.A2( u1_u6_u3_n113 ) , .A1( u1_u6_u3_n114 ) , .ZN( u1_u6_u3_n151 ) );
  INV_X1 u1_u6_u3_U22 (.A( u1_u6_u3_n133 ) , .ZN( u1_u6_u3_n165 ) );
  INV_X1 u1_u6_u3_U23 (.A( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n170 ) );
  NAND2_X1 u1_u6_u3_U24 (.A1( u1_u6_u3_n107 ) , .A2( u1_u6_u3_n108 ) , .ZN( u1_u6_u3_n140 ) );
  NAND2_X1 u1_u6_u3_U25 (.ZN( u1_u6_u3_n117 ) , .A1( u1_u6_u3_n124 ) , .A2( u1_u6_u3_n148 ) );
  NAND2_X1 u1_u6_u3_U26 (.ZN( u1_u6_u3_n143 ) , .A1( u1_u6_u3_n165 ) , .A2( u1_u6_u3_n167 ) );
  INV_X1 u1_u6_u3_U27 (.A( u1_u6_u3_n130 ) , .ZN( u1_u6_u3_n177 ) );
  INV_X1 u1_u6_u3_U28 (.A( u1_u6_u3_n128 ) , .ZN( u1_u6_u3_n176 ) );
  INV_X1 u1_u6_u3_U29 (.A( u1_u6_u3_n155 ) , .ZN( u1_u6_u3_n174 ) );
  INV_X1 u1_u6_u3_U3 (.A( u1_u6_u3_n129 ) , .ZN( u1_u6_u3_n183 ) );
  INV_X1 u1_u6_u3_U30 (.A( u1_u6_u3_n139 ) , .ZN( u1_u6_u3_n185 ) );
  NOR2_X1 u1_u6_u3_U31 (.ZN( u1_u6_u3_n135 ) , .A2( u1_u6_u3_n141 ) , .A1( u1_u6_u3_n169 ) );
  OAI222_X1 u1_u6_u3_U32 (.C2( u1_u6_u3_n107 ) , .A2( u1_u6_u3_n108 ) , .B1( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n138 ) , .B2( u1_u6_u3_n146 ) , .C1( u1_u6_u3_n154 ) , .A1( u1_u6_u3_n164 ) );
  NOR4_X1 u1_u6_u3_U33 (.A4( u1_u6_u3_n157 ) , .A3( u1_u6_u3_n158 ) , .A2( u1_u6_u3_n159 ) , .A1( u1_u6_u3_n160 ) , .ZN( u1_u6_u3_n161 ) );
  AOI21_X1 u1_u6_u3_U34 (.B2( u1_u6_u3_n152 ) , .B1( u1_u6_u3_n153 ) , .ZN( u1_u6_u3_n158 ) , .A( u1_u6_u3_n164 ) );
  AOI21_X1 u1_u6_u3_U35 (.A( u1_u6_u3_n154 ) , .B2( u1_u6_u3_n155 ) , .B1( u1_u6_u3_n156 ) , .ZN( u1_u6_u3_n157 ) );
  AOI21_X1 u1_u6_u3_U36 (.A( u1_u6_u3_n149 ) , .B2( u1_u6_u3_n150 ) , .B1( u1_u6_u3_n151 ) , .ZN( u1_u6_u3_n159 ) );
  AOI211_X1 u1_u6_u3_U37 (.ZN( u1_u6_u3_n109 ) , .A( u1_u6_u3_n119 ) , .C2( u1_u6_u3_n129 ) , .B( u1_u6_u3_n138 ) , .C1( u1_u6_u3_n141 ) );
  AOI211_X1 u1_u6_u3_U38 (.B( u1_u6_u3_n119 ) , .A( u1_u6_u3_n120 ) , .C2( u1_u6_u3_n121 ) , .ZN( u1_u6_u3_n122 ) , .C1( u1_u6_u3_n179 ) );
  INV_X1 u1_u6_u3_U39 (.A( u1_u6_u3_n156 ) , .ZN( u1_u6_u3_n179 ) );
  INV_X1 u1_u6_u3_U4 (.A( u1_u6_u3_n140 ) , .ZN( u1_u6_u3_n182 ) );
  OAI22_X1 u1_u6_u3_U40 (.B1( u1_u6_u3_n118 ) , .ZN( u1_u6_u3_n120 ) , .A1( u1_u6_u3_n135 ) , .B2( u1_u6_u3_n154 ) , .A2( u1_u6_u3_n178 ) );
  AND3_X1 u1_u6_u3_U41 (.ZN( u1_u6_u3_n118 ) , .A2( u1_u6_u3_n124 ) , .A1( u1_u6_u3_n144 ) , .A3( u1_u6_u3_n152 ) );
  INV_X1 u1_u6_u3_U42 (.A( u1_u6_u3_n121 ) , .ZN( u1_u6_u3_n164 ) );
  NAND2_X1 u1_u6_u3_U43 (.ZN( u1_u6_u3_n133 ) , .A1( u1_u6_u3_n154 ) , .A2( u1_u6_u3_n164 ) );
  OAI211_X1 u1_u6_u3_U44 (.B( u1_u6_u3_n127 ) , .ZN( u1_u6_u3_n139 ) , .C1( u1_u6_u3_n150 ) , .C2( u1_u6_u3_n154 ) , .A( u1_u6_u3_n184 ) );
  INV_X1 u1_u6_u3_U45 (.A( u1_u6_u3_n125 ) , .ZN( u1_u6_u3_n184 ) );
  AOI221_X1 u1_u6_u3_U46 (.A( u1_u6_u3_n126 ) , .ZN( u1_u6_u3_n127 ) , .C2( u1_u6_u3_n132 ) , .C1( u1_u6_u3_n169 ) , .B2( u1_u6_u3_n170 ) , .B1( u1_u6_u3_n174 ) );
  OAI22_X1 u1_u6_u3_U47 (.A1( u1_u6_u3_n124 ) , .ZN( u1_u6_u3_n125 ) , .B2( u1_u6_u3_n145 ) , .A2( u1_u6_u3_n165 ) , .B1( u1_u6_u3_n167 ) );
  NOR2_X1 u1_u6_u3_U48 (.A1( u1_u6_u3_n113 ) , .ZN( u1_u6_u3_n131 ) , .A2( u1_u6_u3_n154 ) );
  NAND2_X1 u1_u6_u3_U49 (.A1( u1_u6_u3_n103 ) , .ZN( u1_u6_u3_n150 ) , .A2( u1_u6_u3_n99 ) );
  INV_X1 u1_u6_u3_U5 (.A( u1_u6_u3_n117 ) , .ZN( u1_u6_u3_n178 ) );
  NAND2_X1 u1_u6_u3_U50 (.A2( u1_u6_u3_n102 ) , .ZN( u1_u6_u3_n155 ) , .A1( u1_u6_u3_n97 ) );
  INV_X1 u1_u6_u3_U51 (.A( u1_u6_u3_n141 ) , .ZN( u1_u6_u3_n167 ) );
  AOI21_X1 u1_u6_u3_U52 (.B2( u1_u6_u3_n114 ) , .B1( u1_u6_u3_n146 ) , .A( u1_u6_u3_n154 ) , .ZN( u1_u6_u3_n94 ) );
  AOI21_X1 u1_u6_u3_U53 (.ZN( u1_u6_u3_n110 ) , .B2( u1_u6_u3_n142 ) , .B1( u1_u6_u3_n186 ) , .A( u1_u6_u3_n95 ) );
  INV_X1 u1_u6_u3_U54 (.A( u1_u6_u3_n145 ) , .ZN( u1_u6_u3_n186 ) );
  AOI21_X1 u1_u6_u3_U55 (.B1( u1_u6_u3_n124 ) , .A( u1_u6_u3_n149 ) , .B2( u1_u6_u3_n155 ) , .ZN( u1_u6_u3_n95 ) );
  INV_X1 u1_u6_u3_U56 (.A( u1_u6_u3_n149 ) , .ZN( u1_u6_u3_n169 ) );
  NAND2_X1 u1_u6_u3_U57 (.ZN( u1_u6_u3_n124 ) , .A1( u1_u6_u3_n96 ) , .A2( u1_u6_u3_n97 ) );
  NAND2_X1 u1_u6_u3_U58 (.A2( u1_u6_u3_n100 ) , .ZN( u1_u6_u3_n146 ) , .A1( u1_u6_u3_n96 ) );
  NAND2_X1 u1_u6_u3_U59 (.A1( u1_u6_u3_n101 ) , .ZN( u1_u6_u3_n145 ) , .A2( u1_u6_u3_n99 ) );
  AOI221_X1 u1_u6_u3_U6 (.A( u1_u6_u3_n131 ) , .C2( u1_u6_u3_n132 ) , .C1( u1_u6_u3_n133 ) , .ZN( u1_u6_u3_n134 ) , .B1( u1_u6_u3_n143 ) , .B2( u1_u6_u3_n177 ) );
  NAND2_X1 u1_u6_u3_U60 (.A1( u1_u6_u3_n100 ) , .ZN( u1_u6_u3_n156 ) , .A2( u1_u6_u3_n99 ) );
  NAND2_X1 u1_u6_u3_U61 (.A2( u1_u6_u3_n101 ) , .A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n148 ) );
  NAND2_X1 u1_u6_u3_U62 (.A1( u1_u6_u3_n100 ) , .A2( u1_u6_u3_n102 ) , .ZN( u1_u6_u3_n128 ) );
  NAND2_X1 u1_u6_u3_U63 (.A2( u1_u6_u3_n101 ) , .A1( u1_u6_u3_n102 ) , .ZN( u1_u6_u3_n152 ) );
  NAND2_X1 u1_u6_u3_U64 (.A2( u1_u6_u3_n101 ) , .ZN( u1_u6_u3_n114 ) , .A1( u1_u6_u3_n96 ) );
  NAND2_X1 u1_u6_u3_U65 (.ZN( u1_u6_u3_n107 ) , .A1( u1_u6_u3_n97 ) , .A2( u1_u6_u3_n99 ) );
  NAND2_X1 u1_u6_u3_U66 (.A2( u1_u6_u3_n100 ) , .A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n113 ) );
  NAND2_X1 u1_u6_u3_U67 (.A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n153 ) , .A2( u1_u6_u3_n97 ) );
  NAND2_X1 u1_u6_u3_U68 (.A2( u1_u6_u3_n103 ) , .A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n130 ) );
  NAND2_X1 u1_u6_u3_U69 (.A2( u1_u6_u3_n103 ) , .ZN( u1_u6_u3_n144 ) , .A1( u1_u6_u3_n96 ) );
  OAI22_X1 u1_u6_u3_U7 (.B2( u1_u6_u3_n147 ) , .A2( u1_u6_u3_n148 ) , .ZN( u1_u6_u3_n160 ) , .B1( u1_u6_u3_n165 ) , .A1( u1_u6_u3_n168 ) );
  NAND2_X1 u1_u6_u3_U70 (.A1( u1_u6_u3_n102 ) , .A2( u1_u6_u3_n103 ) , .ZN( u1_u6_u3_n108 ) );
  NOR2_X1 u1_u6_u3_U71 (.A2( u1_u6_X_19 ) , .A1( u1_u6_X_20 ) , .ZN( u1_u6_u3_n99 ) );
  NOR2_X1 u1_u6_u3_U72 (.A2( u1_u6_X_21 ) , .A1( u1_u6_X_24 ) , .ZN( u1_u6_u3_n103 ) );
  NOR2_X1 u1_u6_u3_U73 (.A2( u1_u6_X_24 ) , .A1( u1_u6_u3_n171 ) , .ZN( u1_u6_u3_n97 ) );
  NOR2_X1 u1_u6_u3_U74 (.A2( u1_u6_X_23 ) , .ZN( u1_u6_u3_n141 ) , .A1( u1_u6_u3_n166 ) );
  NOR2_X1 u1_u6_u3_U75 (.A2( u1_u6_X_19 ) , .A1( u1_u6_u3_n172 ) , .ZN( u1_u6_u3_n96 ) );
  NAND2_X1 u1_u6_u3_U76 (.A1( u1_u6_X_22 ) , .A2( u1_u6_X_23 ) , .ZN( u1_u6_u3_n154 ) );
  NAND2_X1 u1_u6_u3_U77 (.A1( u1_u6_X_23 ) , .ZN( u1_u6_u3_n149 ) , .A2( u1_u6_u3_n166 ) );
  NOR2_X1 u1_u6_u3_U78 (.A2( u1_u6_X_22 ) , .A1( u1_u6_X_23 ) , .ZN( u1_u6_u3_n121 ) );
  AND2_X1 u1_u6_u3_U79 (.A1( u1_u6_X_24 ) , .ZN( u1_u6_u3_n101 ) , .A2( u1_u6_u3_n171 ) );
  AND3_X1 u1_u6_u3_U8 (.A3( u1_u6_u3_n144 ) , .A2( u1_u6_u3_n145 ) , .A1( u1_u6_u3_n146 ) , .ZN( u1_u6_u3_n147 ) );
  AND2_X1 u1_u6_u3_U80 (.A1( u1_u6_X_19 ) , .ZN( u1_u6_u3_n102 ) , .A2( u1_u6_u3_n172 ) );
  AND2_X1 u1_u6_u3_U81 (.A1( u1_u6_X_21 ) , .A2( u1_u6_X_24 ) , .ZN( u1_u6_u3_n100 ) );
  AND2_X1 u1_u6_u3_U82 (.A2( u1_u6_X_19 ) , .A1( u1_u6_X_20 ) , .ZN( u1_u6_u3_n104 ) );
  INV_X1 u1_u6_u3_U83 (.A( u1_u6_X_22 ) , .ZN( u1_u6_u3_n166 ) );
  INV_X1 u1_u6_u3_U84 (.A( u1_u6_X_21 ) , .ZN( u1_u6_u3_n171 ) );
  INV_X1 u1_u6_u3_U85 (.A( u1_u6_X_20 ) , .ZN( u1_u6_u3_n172 ) );
  NAND4_X1 u1_u6_u3_U86 (.ZN( u1_out6_20 ) , .A4( u1_u6_u3_n122 ) , .A3( u1_u6_u3_n123 ) , .A1( u1_u6_u3_n175 ) , .A2( u1_u6_u3_n180 ) );
  INV_X1 u1_u6_u3_U87 (.A( u1_u6_u3_n126 ) , .ZN( u1_u6_u3_n180 ) );
  INV_X1 u1_u6_u3_U88 (.A( u1_u6_u3_n112 ) , .ZN( u1_u6_u3_n175 ) );
  NAND4_X1 u1_u6_u3_U89 (.ZN( u1_out6_26 ) , .A4( u1_u6_u3_n109 ) , .A3( u1_u6_u3_n110 ) , .A2( u1_u6_u3_n111 ) , .A1( u1_u6_u3_n173 ) );
  INV_X1 u1_u6_u3_U9 (.A( u1_u6_u3_n143 ) , .ZN( u1_u6_u3_n168 ) );
  INV_X1 u1_u6_u3_U90 (.ZN( u1_u6_u3_n173 ) , .A( u1_u6_u3_n94 ) );
  OAI21_X1 u1_u6_u3_U91 (.ZN( u1_u6_u3_n111 ) , .B2( u1_u6_u3_n117 ) , .A( u1_u6_u3_n133 ) , .B1( u1_u6_u3_n176 ) );
  NAND4_X1 u1_u6_u3_U92 (.ZN( u1_out6_1 ) , .A4( u1_u6_u3_n161 ) , .A3( u1_u6_u3_n162 ) , .A2( u1_u6_u3_n163 ) , .A1( u1_u6_u3_n185 ) );
  NAND2_X1 u1_u6_u3_U93 (.ZN( u1_u6_u3_n163 ) , .A2( u1_u6_u3_n170 ) , .A1( u1_u6_u3_n176 ) );
  AOI22_X1 u1_u6_u3_U94 (.B2( u1_u6_u3_n140 ) , .B1( u1_u6_u3_n141 ) , .A2( u1_u6_u3_n142 ) , .ZN( u1_u6_u3_n162 ) , .A1( u1_u6_u3_n177 ) );
  OR4_X1 u1_u6_u3_U95 (.ZN( u1_out6_10 ) , .A4( u1_u6_u3_n136 ) , .A3( u1_u6_u3_n137 ) , .A1( u1_u6_u3_n138 ) , .A2( u1_u6_u3_n139 ) );
  OAI222_X1 u1_u6_u3_U96 (.C1( u1_u6_u3_n128 ) , .ZN( u1_u6_u3_n137 ) , .B1( u1_u6_u3_n148 ) , .A2( u1_u6_u3_n150 ) , .B2( u1_u6_u3_n154 ) , .C2( u1_u6_u3_n164 ) , .A1( u1_u6_u3_n167 ) );
  OAI221_X1 u1_u6_u3_U97 (.A( u1_u6_u3_n134 ) , .B2( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n136 ) , .C1( u1_u6_u3_n149 ) , .B1( u1_u6_u3_n151 ) , .C2( u1_u6_u3_n183 ) );
  NAND3_X1 u1_u6_u3_U98 (.A1( u1_u6_u3_n114 ) , .ZN( u1_u6_u3_n115 ) , .A2( u1_u6_u3_n145 ) , .A3( u1_u6_u3_n153 ) );
  NAND3_X1 u1_u6_u3_U99 (.ZN( u1_u6_u3_n129 ) , .A2( u1_u6_u3_n144 ) , .A1( u1_u6_u3_n153 ) , .A3( u1_u6_u3_n182 ) );
  OAI21_X1 u1_uk_U135 (.ZN( u1_K2_47 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1033 ) , .B2( u1_uk_n1271 ) );
  NAND2_X1 u1_uk_U136 (.A1( u1_uk_K_r0_52 ) , .ZN( u1_uk_n1033 ) , .A2( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U165 (.ZN( u1_K7_19 ) , .B2( u1_uk_n1495 ) , .A2( u1_uk_n1505 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n92 ) );
  INV_X1 u1_uk_U203 (.ZN( u1_K7_24 ) , .A( u1_uk_n1113 ) );
  AOI22_X1 u1_uk_U204 (.B2( u1_uk_K_r5_18 ) , .A2( u1_uk_K_r5_40 ) , .ZN( u1_uk_n1113 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U286 (.ZN( u1_K2_44 ) , .B2( u1_uk_n1281 ) , .A2( u1_uk_n1303 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U342 (.ZN( u1_K2_46 ) , .A2( u1_uk_n1266 ) , .B2( u1_uk_n1293 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U659 (.ZN( u1_K2_43 ) , .A( u1_uk_n1032 ) , .B2( u1_uk_n1276 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U660 (.A1( u1_uk_K_r0_2 ) , .ZN( u1_uk_n1032 ) , .A2( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U771 (.ZN( u1_K7_21 ) , .A( u1_uk_n1110 ) , .B2( u1_uk_n1526 ) , .B1( u1_uk_n271 ) );
  NAND2_X1 u1_uk_U772 (.A1( u1_uk_K_r5_19 ) , .ZN( u1_uk_n1110 ) , .A2( u1_uk_n217 ) );
  INV_X1 u1_uk_U837 (.ZN( u1_K7_20 ) , .A( u1_uk_n1109 ) );
  AOI22_X1 u1_uk_U838 (.B2( u1_uk_K_r5_18 ) , .A2( u1_uk_K_r5_53 ) , .A1( u1_uk_n11 ) , .ZN( u1_uk_n1109 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U954 (.ZN( u1_K2_48 ) , .B2( u1_uk_n1271 ) , .A2( u1_uk_n1286 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U979 (.ZN( u1_K2_45 ) , .B2( u1_uk_n1282 ) , .A2( u1_uk_n1304 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U996 (.ZN( u1_K7_22 ) , .A( u1_uk_n1111 ) , .B2( u1_uk_n1498 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U997 (.A1( u1_uk_K_r5_5 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1111 ) );
  OAI21_X1 u1_uk_U998 (.ZN( u1_K7_23 ) , .A( u1_uk_n1112 ) , .B2( u1_uk_n1483 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U999 (.A1( u1_uk_K_r5_13 ) , .ZN( u1_uk_n1112 ) , .A2( u1_uk_n17 ) );
  XOR2_X1 u2_U104 (.B( u2_L12_24 ) , .Z( u2_N439 ) , .A( u2_out13_24 ) );
  XOR2_X1 u2_U105 (.B( u2_L12_23 ) , .Z( u2_N438 ) , .A( u2_out13_23 ) );
  XOR2_X1 u2_U106 (.B( u2_L12_22 ) , .Z( u2_N437 ) , .A( u2_out13_22 ) );
  XOR2_X1 u2_U109 (.B( u2_L12_19 ) , .Z( u2_N434 ) , .A( u2_out13_19 ) );
  XOR2_X1 u2_U11 (.B( u2_L1_28 ) , .Z( u2_N91 ) , .A( u2_out2_28 ) );
  XOR2_X1 u2_U110 (.B( u2_L12_18 ) , .Z( u2_N433 ) , .A( u2_out13_18 ) );
  XOR2_X1 u2_U111 (.B( u2_L12_17 ) , .Z( u2_N432 ) , .A( u2_out13_17 ) );
  XOR2_X1 u2_U112 (.B( u2_L12_16 ) , .Z( u2_N431 ) , .A( u2_out13_16 ) );
  XOR2_X1 u2_U116 (.B( u2_L12_13 ) , .Z( u2_N428 ) , .A( u2_out13_13 ) );
  XOR2_X1 u2_U117 (.B( u2_L12_12 ) , .Z( u2_N427 ) , .A( u2_out13_12 ) );
  XOR2_X1 u2_U118 (.B( u2_L12_11 ) , .Z( u2_N426 ) , .A( u2_out13_11 ) );
  XOR2_X1 u2_U120 (.B( u2_L12_9 ) , .Z( u2_N424 ) , .A( u2_out13_9 ) );
  XOR2_X1 u2_U122 (.B( u2_L12_7 ) , .Z( u2_N422 ) , .A( u2_out13_7 ) );
  XOR2_X1 u2_U123 (.B( u2_L12_6 ) , .Z( u2_N421 ) , .A( u2_out13_6 ) );
  XOR2_X1 u2_U126 (.B( u2_L12_4 ) , .Z( u2_N419 ) , .A( u2_out13_4 ) );
  XOR2_X1 u2_U128 (.B( u2_L12_2 ) , .Z( u2_N417 ) , .A( u2_out13_2 ) );
  XOR2_X1 u2_U207 (.B( u2_L9_27 ) , .Z( u2_N346 ) , .A( u2_out10_27 ) );
  XOR2_X1 u2_U213 (.B( u2_L9_21 ) , .Z( u2_N340 ) , .A( u2_out10_21 ) );
  XOR2_X1 u2_U22 (.B( u2_L1_18 ) , .Z( u2_N81 ) , .A( u2_out2_18 ) );
  XOR2_X1 u2_U220 (.B( u2_L9_15 ) , .Z( u2_N334 ) , .A( u2_out10_15 ) );
  XOR2_X1 u2_U231 (.B( u2_L9_5 ) , .Z( u2_N324 ) , .A( u2_out10_5 ) );
  XOR2_X1 u2_U274 (.B( u2_L7_31 ) , .Z( u2_N286 ) , .A( u2_out8_31 ) );
  XOR2_X1 u2_U275 (.B( u2_L7_30 ) , .Z( u2_N285 ) , .A( u2_out8_30 ) );
  XOR2_X1 u2_U277 (.B( u2_L7_28 ) , .Z( u2_N283 ) , .A( u2_out8_28 ) );
  XOR2_X1 u2_U28 (.B( u2_L1_13 ) , .Z( u2_N76 ) , .A( u2_out2_13 ) );
  XOR2_X1 u2_U282 (.B( u2_L7_24 ) , .Z( u2_N279 ) , .A( u2_out8_24 ) );
  XOR2_X1 u2_U283 (.B( u2_L7_23 ) , .Z( u2_N278 ) , .A( u2_out8_23 ) );
  XOR2_X1 u2_U288 (.B( u2_L7_18 ) , .Z( u2_N273 ) , .A( u2_out8_18 ) );
  XOR2_X1 u2_U289 (.B( u2_L7_17 ) , .Z( u2_N272 ) , .A( u2_out8_17 ) );
  XOR2_X1 u2_U290 (.B( u2_L7_16 ) , .Z( u2_N271 ) , .A( u2_out8_16 ) );
  XOR2_X1 u2_U294 (.B( u2_L7_13 ) , .Z( u2_N268 ) , .A( u2_out8_13 ) );
  XOR2_X1 u2_U298 (.B( u2_L7_9 ) , .Z( u2_N264 ) , .A( u2_out8_9 ) );
  XOR2_X1 u2_U301 (.B( u2_L7_6 ) , .Z( u2_N261 ) , .A( u2_out8_6 ) );
  XOR2_X1 u2_U306 (.B( u2_L7_2 ) , .Z( u2_N257 ) , .A( u2_out8_2 ) );
  XOR2_X1 u2_U312 (.B( u2_L6_28 ) , .Z( u2_N251 ) , .A( u2_out7_28 ) );
  XOR2_X1 u2_U323 (.B( u2_L6_18 ) , .Z( u2_N241 ) , .A( u2_out7_18 ) );
  XOR2_X1 u2_U329 (.B( u2_L6_13 ) , .Z( u2_N236 ) , .A( u2_out7_13 ) );
  XOR2_X1 u2_U341 (.B( u2_L6_2 ) , .Z( u2_N225 ) , .A( u2_out7_2 ) );
  XOR2_X1 u2_U40 (.B( u2_L1_2 ) , .Z( u2_N65 ) , .A( u2_out2_2 ) );
  XOR2_X1 u2_U452 (.B( u2_L2_30 ) , .Z( u2_N125 ) , .A( u2_out3_30 ) );
  XOR2_X1 u2_U456 (.B( u2_L2_26 ) , .Z( u2_N121 ) , .A( u2_out3_26 ) );
  XOR2_X1 u2_U459 (.B( u2_L2_24 ) , .Z( u2_N119 ) , .A( u2_out3_24 ) );
  XOR2_X1 u2_U463 (.B( u2_L2_20 ) , .Z( u2_N115 ) , .A( u2_out3_20 ) );
  XOR2_X1 u2_U467 (.B( u2_L2_16 ) , .Z( u2_N111 ) , .A( u2_out3_16 ) );
  XOR2_X1 u2_U474 (.B( u2_L2_10 ) , .Z( u2_N105 ) , .A( u2_out3_10 ) );
  XOR2_X1 u2_U478 (.B( u2_L2_6 ) , .Z( u2_N101 ) , .A( u2_out3_6 ) );
  XOR2_X1 u2_U6 (.B( u2_L2_1 ) , .Z( u2_N96 ) , .A( u2_out3_1 ) );
  XOR2_X1 u2_U60 (.B( u2_L13_32 ) , .Z( u2_N479 ) , .A( u2_out14_32 ) );
  XOR2_X1 u2_U63 (.B( u2_L13_29 ) , .Z( u2_N476 ) , .A( u2_out14_29 ) );
  XOR2_X1 u2_U65 (.B( u2_L13_27 ) , .Z( u2_N474 ) , .A( u2_out14_27 ) );
  XOR2_X1 u2_U67 (.B( u2_L13_25 ) , .Z( u2_N472 ) , .A( u2_out14_25 ) );
  XOR2_X1 u2_U71 (.B( u2_L13_22 ) , .Z( u2_N469 ) , .A( u2_out14_22 ) );
  XOR2_X1 u2_U72 (.B( u2_L13_21 ) , .Z( u2_N468 ) , .A( u2_out14_21 ) );
  XOR2_X1 u2_U74 (.B( u2_L13_19 ) , .Z( u2_N466 ) , .A( u2_out14_19 ) );
  XOR2_X1 u2_U78 (.B( u2_L13_15 ) , .Z( u2_N462 ) , .A( u2_out14_15 ) );
  XOR2_X1 u2_U79 (.B( u2_L13_14 ) , .Z( u2_N461 ) , .A( u2_out14_14 ) );
  XOR2_X1 u2_U82 (.B( u2_L13_12 ) , .Z( u2_N459 ) , .A( u2_out14_12 ) );
  XOR2_X1 u2_U83 (.B( u2_L13_11 ) , .Z( u2_N458 ) , .A( u2_out14_11 ) );
  XOR2_X1 u2_U86 (.B( u2_L13_8 ) , .Z( u2_N455 ) , .A( u2_out14_8 ) );
  XOR2_X1 u2_U87 (.B( u2_L13_7 ) , .Z( u2_N454 ) , .A( u2_out14_7 ) );
  XOR2_X1 u2_U89 (.B( u2_L13_5 ) , .Z( u2_N452 ) , .A( u2_out14_5 ) );
  XOR2_X1 u2_U90 (.B( u2_L13_4 ) , .Z( u2_N451 ) , .A( u2_out14_4 ) );
  XOR2_X1 u2_U91 (.B( u2_L13_3 ) , .Z( u2_N450 ) , .A( u2_out14_3 ) );
  XOR2_X1 u2_U95 (.B( u2_L12_32 ) , .Z( u2_N447 ) , .A( u2_out13_32 ) );
  XOR2_X1 u2_U96 (.B( u2_L12_31 ) , .Z( u2_N446 ) , .A( u2_out13_31 ) );
  XOR2_X1 u2_U97 (.B( u2_L12_30 ) , .Z( u2_N445 ) , .A( u2_out13_30 ) );
  XOR2_X1 u2_U98 (.B( u2_L12_29 ) , .Z( u2_N444 ) , .A( u2_out13_29 ) );
  XOR2_X1 u2_U99 (.B( u2_L12_28 ) , .Z( u2_N443 ) , .A( u2_out13_28 ) );
  XOR2_X1 u2_u10_U10 (.B( u2_K11_45 ) , .A( u2_R9_30 ) , .Z( u2_u10_X_45 ) );
  XOR2_X1 u2_u10_U11 (.B( u2_K11_44 ) , .A( u2_R9_29 ) , .Z( u2_u10_X_44 ) );
  XOR2_X1 u2_u10_U12 (.B( u2_K11_43 ) , .A( u2_R9_28 ) , .Z( u2_u10_X_43 ) );
  XOR2_X1 u2_u10_U7 (.B( u2_K11_48 ) , .A( u2_R9_1 ) , .Z( u2_u10_X_48 ) );
  XOR2_X1 u2_u10_U8 (.B( u2_K11_47 ) , .A( u2_R9_32 ) , .Z( u2_u10_X_47 ) );
  XOR2_X1 u2_u10_U9 (.B( u2_K11_46 ) , .A( u2_R9_31 ) , .Z( u2_u10_X_46 ) );
  AND3_X1 u2_u10_u7_U10 (.A3( u2_u10_u7_n110 ) , .A2( u2_u10_u7_n127 ) , .A1( u2_u10_u7_n132 ) , .ZN( u2_u10_u7_n92 ) );
  OAI21_X1 u2_u10_u7_U11 (.A( u2_u10_u7_n161 ) , .B1( u2_u10_u7_n168 ) , .B2( u2_u10_u7_n173 ) , .ZN( u2_u10_u7_n91 ) );
  AOI211_X1 u2_u10_u7_U12 (.A( u2_u10_u7_n117 ) , .ZN( u2_u10_u7_n118 ) , .C2( u2_u10_u7_n126 ) , .C1( u2_u10_u7_n177 ) , .B( u2_u10_u7_n180 ) );
  OAI22_X1 u2_u10_u7_U13 (.B1( u2_u10_u7_n115 ) , .ZN( u2_u10_u7_n117 ) , .A2( u2_u10_u7_n133 ) , .A1( u2_u10_u7_n137 ) , .B2( u2_u10_u7_n162 ) );
  INV_X1 u2_u10_u7_U14 (.A( u2_u10_u7_n116 ) , .ZN( u2_u10_u7_n180 ) );
  NOR3_X1 u2_u10_u7_U15 (.ZN( u2_u10_u7_n115 ) , .A3( u2_u10_u7_n145 ) , .A2( u2_u10_u7_n168 ) , .A1( u2_u10_u7_n169 ) );
  OAI211_X1 u2_u10_u7_U16 (.B( u2_u10_u7_n122 ) , .A( u2_u10_u7_n123 ) , .C2( u2_u10_u7_n124 ) , .ZN( u2_u10_u7_n154 ) , .C1( u2_u10_u7_n162 ) );
  AOI222_X1 u2_u10_u7_U17 (.ZN( u2_u10_u7_n122 ) , .C2( u2_u10_u7_n126 ) , .C1( u2_u10_u7_n145 ) , .B1( u2_u10_u7_n161 ) , .A2( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n170 ) , .A1( u2_u10_u7_n176 ) );
  INV_X1 u2_u10_u7_U18 (.A( u2_u10_u7_n133 ) , .ZN( u2_u10_u7_n176 ) );
  NOR3_X1 u2_u10_u7_U19 (.A2( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n135 ) , .ZN( u2_u10_u7_n136 ) , .A3( u2_u10_u7_n171 ) );
  NOR2_X1 u2_u10_u7_U20 (.A1( u2_u10_u7_n130 ) , .A2( u2_u10_u7_n134 ) , .ZN( u2_u10_u7_n153 ) );
  INV_X1 u2_u10_u7_U21 (.A( u2_u10_u7_n101 ) , .ZN( u2_u10_u7_n165 ) );
  NOR2_X1 u2_u10_u7_U22 (.ZN( u2_u10_u7_n111 ) , .A2( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n169 ) );
  AOI21_X1 u2_u10_u7_U23 (.ZN( u2_u10_u7_n104 ) , .B2( u2_u10_u7_n112 ) , .B1( u2_u10_u7_n127 ) , .A( u2_u10_u7_n164 ) );
  AOI21_X1 u2_u10_u7_U24 (.ZN( u2_u10_u7_n106 ) , .B1( u2_u10_u7_n133 ) , .B2( u2_u10_u7_n146 ) , .A( u2_u10_u7_n162 ) );
  AOI21_X1 u2_u10_u7_U25 (.A( u2_u10_u7_n101 ) , .ZN( u2_u10_u7_n107 ) , .B2( u2_u10_u7_n128 ) , .B1( u2_u10_u7_n175 ) );
  INV_X1 u2_u10_u7_U26 (.A( u2_u10_u7_n138 ) , .ZN( u2_u10_u7_n171 ) );
  INV_X1 u2_u10_u7_U27 (.A( u2_u10_u7_n131 ) , .ZN( u2_u10_u7_n177 ) );
  INV_X1 u2_u10_u7_U28 (.A( u2_u10_u7_n110 ) , .ZN( u2_u10_u7_n174 ) );
  NAND2_X1 u2_u10_u7_U29 (.A1( u2_u10_u7_n129 ) , .A2( u2_u10_u7_n132 ) , .ZN( u2_u10_u7_n149 ) );
  OAI21_X1 u2_u10_u7_U3 (.ZN( u2_u10_u7_n159 ) , .A( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n171 ) , .B1( u2_u10_u7_n174 ) );
  NAND2_X1 u2_u10_u7_U30 (.A1( u2_u10_u7_n113 ) , .A2( u2_u10_u7_n124 ) , .ZN( u2_u10_u7_n130 ) );
  INV_X1 u2_u10_u7_U31 (.A( u2_u10_u7_n112 ) , .ZN( u2_u10_u7_n173 ) );
  INV_X1 u2_u10_u7_U32 (.A( u2_u10_u7_n128 ) , .ZN( u2_u10_u7_n168 ) );
  INV_X1 u2_u10_u7_U33 (.A( u2_u10_u7_n148 ) , .ZN( u2_u10_u7_n169 ) );
  INV_X1 u2_u10_u7_U34 (.A( u2_u10_u7_n127 ) , .ZN( u2_u10_u7_n179 ) );
  NOR2_X1 u2_u10_u7_U35 (.ZN( u2_u10_u7_n101 ) , .A2( u2_u10_u7_n150 ) , .A1( u2_u10_u7_n156 ) );
  AOI211_X1 u2_u10_u7_U36 (.B( u2_u10_u7_n154 ) , .A( u2_u10_u7_n155 ) , .C1( u2_u10_u7_n156 ) , .ZN( u2_u10_u7_n157 ) , .C2( u2_u10_u7_n172 ) );
  INV_X1 u2_u10_u7_U37 (.A( u2_u10_u7_n153 ) , .ZN( u2_u10_u7_n172 ) );
  AOI211_X1 u2_u10_u7_U38 (.B( u2_u10_u7_n139 ) , .A( u2_u10_u7_n140 ) , .C2( u2_u10_u7_n141 ) , .ZN( u2_u10_u7_n142 ) , .C1( u2_u10_u7_n156 ) );
  NAND4_X1 u2_u10_u7_U39 (.A3( u2_u10_u7_n127 ) , .A2( u2_u10_u7_n128 ) , .A1( u2_u10_u7_n129 ) , .ZN( u2_u10_u7_n141 ) , .A4( u2_u10_u7_n147 ) );
  INV_X1 u2_u10_u7_U4 (.A( u2_u10_u7_n111 ) , .ZN( u2_u10_u7_n170 ) );
  AOI21_X1 u2_u10_u7_U40 (.A( u2_u10_u7_n137 ) , .B1( u2_u10_u7_n138 ) , .ZN( u2_u10_u7_n139 ) , .B2( u2_u10_u7_n146 ) );
  OAI22_X1 u2_u10_u7_U41 (.B1( u2_u10_u7_n136 ) , .ZN( u2_u10_u7_n140 ) , .A1( u2_u10_u7_n153 ) , .B2( u2_u10_u7_n162 ) , .A2( u2_u10_u7_n164 ) );
  AOI21_X1 u2_u10_u7_U42 (.ZN( u2_u10_u7_n123 ) , .B1( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n177 ) , .A( u2_u10_u7_n97 ) );
  AOI21_X1 u2_u10_u7_U43 (.B2( u2_u10_u7_n113 ) , .B1( u2_u10_u7_n124 ) , .A( u2_u10_u7_n125 ) , .ZN( u2_u10_u7_n97 ) );
  INV_X1 u2_u10_u7_U44 (.A( u2_u10_u7_n125 ) , .ZN( u2_u10_u7_n161 ) );
  INV_X1 u2_u10_u7_U45 (.A( u2_u10_u7_n152 ) , .ZN( u2_u10_u7_n162 ) );
  AOI22_X1 u2_u10_u7_U46 (.A2( u2_u10_u7_n114 ) , .ZN( u2_u10_u7_n119 ) , .B1( u2_u10_u7_n130 ) , .A1( u2_u10_u7_n156 ) , .B2( u2_u10_u7_n165 ) );
  NAND2_X1 u2_u10_u7_U47 (.A2( u2_u10_u7_n112 ) , .ZN( u2_u10_u7_n114 ) , .A1( u2_u10_u7_n175 ) );
  AND2_X1 u2_u10_u7_U48 (.ZN( u2_u10_u7_n145 ) , .A2( u2_u10_u7_n98 ) , .A1( u2_u10_u7_n99 ) );
  NOR2_X1 u2_u10_u7_U49 (.ZN( u2_u10_u7_n137 ) , .A1( u2_u10_u7_n150 ) , .A2( u2_u10_u7_n161 ) );
  INV_X1 u2_u10_u7_U5 (.A( u2_u10_u7_n149 ) , .ZN( u2_u10_u7_n175 ) );
  AOI21_X1 u2_u10_u7_U50 (.ZN( u2_u10_u7_n105 ) , .B2( u2_u10_u7_n110 ) , .A( u2_u10_u7_n125 ) , .B1( u2_u10_u7_n147 ) );
  NAND2_X1 u2_u10_u7_U51 (.ZN( u2_u10_u7_n146 ) , .A1( u2_u10_u7_n95 ) , .A2( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U52 (.A2( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n147 ) , .A1( u2_u10_u7_n93 ) );
  NAND2_X1 u2_u10_u7_U53 (.A1( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n127 ) , .A2( u2_u10_u7_n99 ) );
  OR2_X1 u2_u10_u7_U54 (.ZN( u2_u10_u7_n126 ) , .A2( u2_u10_u7_n152 ) , .A1( u2_u10_u7_n156 ) );
  NAND2_X1 u2_u10_u7_U55 (.A2( u2_u10_u7_n102 ) , .A1( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n133 ) );
  NAND2_X1 u2_u10_u7_U56 (.ZN( u2_u10_u7_n112 ) , .A2( u2_u10_u7_n96 ) , .A1( u2_u10_u7_n99 ) );
  NAND2_X1 u2_u10_u7_U57 (.A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n128 ) , .A1( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U58 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n113 ) , .A2( u2_u10_u7_n93 ) );
  NAND2_X1 u2_u10_u7_U59 (.A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n124 ) , .A1( u2_u10_u7_n96 ) );
  INV_X1 u2_u10_u7_U6 (.A( u2_u10_u7_n154 ) , .ZN( u2_u10_u7_n178 ) );
  NAND2_X1 u2_u10_u7_U60 (.ZN( u2_u10_u7_n110 ) , .A1( u2_u10_u7_n95 ) , .A2( u2_u10_u7_n96 ) );
  INV_X1 u2_u10_u7_U61 (.A( u2_u10_u7_n150 ) , .ZN( u2_u10_u7_n164 ) );
  AND2_X1 u2_u10_u7_U62 (.ZN( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n93 ) , .A2( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U63 (.A1( u2_u10_u7_n100 ) , .A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n129 ) );
  NAND2_X1 u2_u10_u7_U64 (.A2( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n131 ) , .A1( u2_u10_u7_n95 ) );
  NAND2_X1 u2_u10_u7_U65 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n138 ) , .A2( u2_u10_u7_n99 ) );
  NAND2_X1 u2_u10_u7_U66 (.ZN( u2_u10_u7_n132 ) , .A1( u2_u10_u7_n93 ) , .A2( u2_u10_u7_n96 ) );
  NAND2_X1 u2_u10_u7_U67 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n148 ) , .A2( u2_u10_u7_n95 ) );
  NOR2_X1 u2_u10_u7_U68 (.A2( u2_u10_X_47 ) , .ZN( u2_u10_u7_n150 ) , .A1( u2_u10_u7_n163 ) );
  NOR2_X1 u2_u10_u7_U69 (.A2( u2_u10_X_43 ) , .A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n103 ) );
  AOI211_X1 u2_u10_u7_U7 (.ZN( u2_u10_u7_n116 ) , .A( u2_u10_u7_n155 ) , .C1( u2_u10_u7_n161 ) , .C2( u2_u10_u7_n171 ) , .B( u2_u10_u7_n94 ) );
  NOR2_X1 u2_u10_u7_U70 (.A2( u2_u10_X_48 ) , .A1( u2_u10_u7_n166 ) , .ZN( u2_u10_u7_n95 ) );
  NOR2_X1 u2_u10_u7_U71 (.A2( u2_u10_X_45 ) , .A1( u2_u10_X_48 ) , .ZN( u2_u10_u7_n99 ) );
  NOR2_X1 u2_u10_u7_U72 (.A2( u2_u10_X_44 ) , .A1( u2_u10_u7_n167 ) , .ZN( u2_u10_u7_n98 ) );
  NOR2_X1 u2_u10_u7_U73 (.A2( u2_u10_X_46 ) , .A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n152 ) );
  AND2_X1 u2_u10_u7_U74 (.A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n156 ) , .A2( u2_u10_u7_n163 ) );
  NAND2_X1 u2_u10_u7_U75 (.A2( u2_u10_X_46 ) , .A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n125 ) );
  AND2_X1 u2_u10_u7_U76 (.A2( u2_u10_X_45 ) , .A1( u2_u10_X_48 ) , .ZN( u2_u10_u7_n102 ) );
  AND2_X1 u2_u10_u7_U77 (.A2( u2_u10_X_43 ) , .A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n96 ) );
  AND2_X1 u2_u10_u7_U78 (.A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n100 ) , .A2( u2_u10_u7_n167 ) );
  AND2_X1 u2_u10_u7_U79 (.A1( u2_u10_X_48 ) , .A2( u2_u10_u7_n166 ) , .ZN( u2_u10_u7_n93 ) );
  OAI222_X1 u2_u10_u7_U8 (.C2( u2_u10_u7_n101 ) , .B2( u2_u10_u7_n111 ) , .A1( u2_u10_u7_n113 ) , .C1( u2_u10_u7_n146 ) , .A2( u2_u10_u7_n162 ) , .B1( u2_u10_u7_n164 ) , .ZN( u2_u10_u7_n94 ) );
  INV_X1 u2_u10_u7_U80 (.A( u2_u10_X_46 ) , .ZN( u2_u10_u7_n163 ) );
  INV_X1 u2_u10_u7_U81 (.A( u2_u10_X_43 ) , .ZN( u2_u10_u7_n167 ) );
  INV_X1 u2_u10_u7_U82 (.A( u2_u10_X_45 ) , .ZN( u2_u10_u7_n166 ) );
  NAND4_X1 u2_u10_u7_U83 (.ZN( u2_out10_27 ) , .A4( u2_u10_u7_n118 ) , .A3( u2_u10_u7_n119 ) , .A2( u2_u10_u7_n120 ) , .A1( u2_u10_u7_n121 ) );
  OAI21_X1 u2_u10_u7_U84 (.ZN( u2_u10_u7_n121 ) , .B2( u2_u10_u7_n145 ) , .A( u2_u10_u7_n150 ) , .B1( u2_u10_u7_n174 ) );
  OAI21_X1 u2_u10_u7_U85 (.ZN( u2_u10_u7_n120 ) , .A( u2_u10_u7_n161 ) , .B2( u2_u10_u7_n170 ) , .B1( u2_u10_u7_n179 ) );
  NAND4_X1 u2_u10_u7_U86 (.ZN( u2_out10_21 ) , .A4( u2_u10_u7_n157 ) , .A3( u2_u10_u7_n158 ) , .A2( u2_u10_u7_n159 ) , .A1( u2_u10_u7_n160 ) );
  OAI21_X1 u2_u10_u7_U87 (.B1( u2_u10_u7_n145 ) , .ZN( u2_u10_u7_n160 ) , .A( u2_u10_u7_n161 ) , .B2( u2_u10_u7_n177 ) );
  AOI22_X1 u2_u10_u7_U88 (.B2( u2_u10_u7_n149 ) , .B1( u2_u10_u7_n150 ) , .A2( u2_u10_u7_n151 ) , .A1( u2_u10_u7_n152 ) , .ZN( u2_u10_u7_n158 ) );
  NAND4_X1 u2_u10_u7_U89 (.ZN( u2_out10_15 ) , .A4( u2_u10_u7_n142 ) , .A3( u2_u10_u7_n143 ) , .A2( u2_u10_u7_n144 ) , .A1( u2_u10_u7_n178 ) );
  OAI221_X1 u2_u10_u7_U9 (.C1( u2_u10_u7_n101 ) , .C2( u2_u10_u7_n147 ) , .ZN( u2_u10_u7_n155 ) , .B2( u2_u10_u7_n162 ) , .A( u2_u10_u7_n91 ) , .B1( u2_u10_u7_n92 ) );
  OR2_X1 u2_u10_u7_U90 (.A2( u2_u10_u7_n125 ) , .A1( u2_u10_u7_n129 ) , .ZN( u2_u10_u7_n144 ) );
  AOI22_X1 u2_u10_u7_U91 (.A2( u2_u10_u7_n126 ) , .ZN( u2_u10_u7_n143 ) , .B2( u2_u10_u7_n165 ) , .B1( u2_u10_u7_n173 ) , .A1( u2_u10_u7_n174 ) );
  NAND4_X1 u2_u10_u7_U92 (.ZN( u2_out10_5 ) , .A4( u2_u10_u7_n108 ) , .A3( u2_u10_u7_n109 ) , .A1( u2_u10_u7_n116 ) , .A2( u2_u10_u7_n123 ) );
  AOI22_X1 u2_u10_u7_U93 (.ZN( u2_u10_u7_n109 ) , .A2( u2_u10_u7_n126 ) , .B2( u2_u10_u7_n145 ) , .B1( u2_u10_u7_n156 ) , .A1( u2_u10_u7_n171 ) );
  NOR4_X1 u2_u10_u7_U94 (.A4( u2_u10_u7_n104 ) , .A3( u2_u10_u7_n105 ) , .A2( u2_u10_u7_n106 ) , .A1( u2_u10_u7_n107 ) , .ZN( u2_u10_u7_n108 ) );
  NAND3_X1 u2_u10_u7_U95 (.A3( u2_u10_u7_n146 ) , .A2( u2_u10_u7_n147 ) , .A1( u2_u10_u7_n148 ) , .ZN( u2_u10_u7_n151 ) );
  NAND3_X1 u2_u10_u7_U96 (.A3( u2_u10_u7_n131 ) , .A2( u2_u10_u7_n132 ) , .A1( u2_u10_u7_n133 ) , .ZN( u2_u10_u7_n135 ) );
  XOR2_X1 u2_u13_U1 (.B( u2_K14_9 ) , .A( u2_R12_6 ) , .Z( u2_u13_X_9 ) );
  XOR2_X1 u2_u13_U13 (.B( u2_K14_42 ) , .A( u2_R12_29 ) , .Z( u2_u13_X_42 ) );
  XOR2_X1 u2_u13_U14 (.B( u2_K14_41 ) , .A( u2_R12_28 ) , .Z( u2_u13_X_41 ) );
  XOR2_X1 u2_u13_U15 (.B( u2_K14_40 ) , .A( u2_R12_27 ) , .Z( u2_u13_X_40 ) );
  XOR2_X1 u2_u13_U16 (.B( u2_K14_3 ) , .A( u2_R12_2 ) , .Z( u2_u13_X_3 ) );
  XOR2_X1 u2_u13_U17 (.B( u2_K14_39 ) , .A( u2_R12_26 ) , .Z( u2_u13_X_39 ) );
  XOR2_X1 u2_u13_U18 (.B( u2_K14_38 ) , .A( u2_R12_25 ) , .Z( u2_u13_X_38 ) );
  XOR2_X1 u2_u13_U19 (.B( u2_K14_37 ) , .A( u2_R12_24 ) , .Z( u2_u13_X_37 ) );
  XOR2_X1 u2_u13_U2 (.B( u2_K14_8 ) , .A( u2_R12_5 ) , .Z( u2_u13_X_8 ) );
  XOR2_X1 u2_u13_U20 (.B( u2_K14_36 ) , .A( u2_R12_25 ) , .Z( u2_u13_X_36 ) );
  XOR2_X1 u2_u13_U21 (.B( u2_K14_35 ) , .A( u2_R12_24 ) , .Z( u2_u13_X_35 ) );
  XOR2_X1 u2_u13_U22 (.B( u2_K14_34 ) , .A( u2_R12_23 ) , .Z( u2_u13_X_34 ) );
  XOR2_X1 u2_u13_U23 (.B( u2_K14_33 ) , .A( u2_R12_22 ) , .Z( u2_u13_X_33 ) );
  XOR2_X1 u2_u13_U24 (.B( u2_K14_32 ) , .A( u2_R12_21 ) , .Z( u2_u13_X_32 ) );
  XOR2_X1 u2_u13_U25 (.B( u2_K14_31 ) , .A( u2_R12_20 ) , .Z( u2_u13_X_31 ) );
  XOR2_X1 u2_u13_U27 (.B( u2_K14_2 ) , .A( u2_R12_1 ) , .Z( u2_u13_X_2 ) );
  XOR2_X1 u2_u13_U3 (.B( u2_K14_7 ) , .A( u2_R12_4 ) , .Z( u2_u13_X_7 ) );
  XOR2_X1 u2_u13_U38 (.B( u2_K14_1 ) , .A( u2_R12_32 ) , .Z( u2_u13_X_1 ) );
  XOR2_X1 u2_u13_U4 (.B( u2_K14_6 ) , .A( u2_R12_5 ) , .Z( u2_u13_X_6 ) );
  XOR2_X1 u2_u13_U40 (.B( u2_K14_18 ) , .A( u2_R12_13 ) , .Z( u2_u13_X_18 ) );
  XOR2_X1 u2_u13_U41 (.B( u2_K14_17 ) , .A( u2_R12_12 ) , .Z( u2_u13_X_17 ) );
  XOR2_X1 u2_u13_U42 (.B( u2_K14_16 ) , .A( u2_R12_11 ) , .Z( u2_u13_X_16 ) );
  XOR2_X1 u2_u13_U43 (.B( u2_K14_15 ) , .A( u2_R12_10 ) , .Z( u2_u13_X_15 ) );
  XOR2_X1 u2_u13_U44 (.B( u2_K14_14 ) , .A( u2_R12_9 ) , .Z( u2_u13_X_14 ) );
  XOR2_X1 u2_u13_U45 (.B( u2_K14_13 ) , .A( u2_R12_8 ) , .Z( u2_u13_X_13 ) );
  XOR2_X1 u2_u13_U46 (.B( u2_K14_12 ) , .A( u2_R12_9 ) , .Z( u2_u13_X_12 ) );
  XOR2_X1 u2_u13_U47 (.B( u2_K14_11 ) , .A( u2_R12_8 ) , .Z( u2_u13_X_11 ) );
  XOR2_X1 u2_u13_U48 (.B( u2_K14_10 ) , .A( u2_R12_7 ) , .Z( u2_u13_X_10 ) );
  XOR2_X1 u2_u13_U5 (.B( u2_K14_5 ) , .A( u2_R12_4 ) , .Z( u2_u13_X_5 ) );
  XOR2_X1 u2_u13_U6 (.B( u2_K14_4 ) , .A( u2_R12_3 ) , .Z( u2_u13_X_4 ) );
  AND3_X1 u2_u13_u0_U10 (.A2( u2_u13_u0_n112 ) , .ZN( u2_u13_u0_n127 ) , .A3( u2_u13_u0_n130 ) , .A1( u2_u13_u0_n148 ) );
  NAND2_X1 u2_u13_u0_U11 (.ZN( u2_u13_u0_n113 ) , .A1( u2_u13_u0_n139 ) , .A2( u2_u13_u0_n149 ) );
  AND2_X1 u2_u13_u0_U12 (.ZN( u2_u13_u0_n107 ) , .A1( u2_u13_u0_n130 ) , .A2( u2_u13_u0_n140 ) );
  AND2_X1 u2_u13_u0_U13 (.A2( u2_u13_u0_n129 ) , .A1( u2_u13_u0_n130 ) , .ZN( u2_u13_u0_n151 ) );
  AND2_X1 u2_u13_u0_U14 (.A1( u2_u13_u0_n108 ) , .A2( u2_u13_u0_n125 ) , .ZN( u2_u13_u0_n145 ) );
  INV_X1 u2_u13_u0_U15 (.A( u2_u13_u0_n143 ) , .ZN( u2_u13_u0_n173 ) );
  NOR2_X1 u2_u13_u0_U16 (.A2( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n147 ) , .A1( u2_u13_u0_n160 ) );
  INV_X1 u2_u13_u0_U17 (.ZN( u2_u13_u0_n172 ) , .A( u2_u13_u0_n88 ) );
  OAI222_X1 u2_u13_u0_U18 (.C1( u2_u13_u0_n108 ) , .A1( u2_u13_u0_n125 ) , .B2( u2_u13_u0_n128 ) , .B1( u2_u13_u0_n144 ) , .A2( u2_u13_u0_n158 ) , .C2( u2_u13_u0_n161 ) , .ZN( u2_u13_u0_n88 ) );
  NOR2_X1 u2_u13_u0_U19 (.A1( u2_u13_u0_n163 ) , .A2( u2_u13_u0_n164 ) , .ZN( u2_u13_u0_n95 ) );
  AOI21_X1 u2_u13_u0_U20 (.B1( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n132 ) , .A( u2_u13_u0_n165 ) , .B2( u2_u13_u0_n93 ) );
  INV_X1 u2_u13_u0_U21 (.A( u2_u13_u0_n142 ) , .ZN( u2_u13_u0_n165 ) );
  OAI221_X1 u2_u13_u0_U22 (.C1( u2_u13_u0_n121 ) , .ZN( u2_u13_u0_n122 ) , .B2( u2_u13_u0_n127 ) , .A( u2_u13_u0_n143 ) , .B1( u2_u13_u0_n144 ) , .C2( u2_u13_u0_n147 ) );
  OAI22_X1 u2_u13_u0_U23 (.B1( u2_u13_u0_n125 ) , .ZN( u2_u13_u0_n126 ) , .A1( u2_u13_u0_n138 ) , .A2( u2_u13_u0_n146 ) , .B2( u2_u13_u0_n147 ) );
  OAI22_X1 u2_u13_u0_U24 (.B1( u2_u13_u0_n131 ) , .A1( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n147 ) , .A2( u2_u13_u0_n90 ) , .ZN( u2_u13_u0_n91 ) );
  AND3_X1 u2_u13_u0_U25 (.A3( u2_u13_u0_n121 ) , .A2( u2_u13_u0_n125 ) , .A1( u2_u13_u0_n148 ) , .ZN( u2_u13_u0_n90 ) );
  INV_X1 u2_u13_u0_U26 (.A( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n161 ) );
  NOR2_X1 u2_u13_u0_U27 (.A1( u2_u13_u0_n120 ) , .ZN( u2_u13_u0_n143 ) , .A2( u2_u13_u0_n167 ) );
  OAI221_X1 u2_u13_u0_U28 (.C1( u2_u13_u0_n112 ) , .ZN( u2_u13_u0_n120 ) , .B1( u2_u13_u0_n138 ) , .B2( u2_u13_u0_n141 ) , .C2( u2_u13_u0_n147 ) , .A( u2_u13_u0_n172 ) );
  AOI211_X1 u2_u13_u0_U29 (.B( u2_u13_u0_n115 ) , .A( u2_u13_u0_n116 ) , .C2( u2_u13_u0_n117 ) , .C1( u2_u13_u0_n118 ) , .ZN( u2_u13_u0_n119 ) );
  INV_X1 u2_u13_u0_U3 (.A( u2_u13_u0_n113 ) , .ZN( u2_u13_u0_n166 ) );
  AOI22_X1 u2_u13_u0_U30 (.B2( u2_u13_u0_n109 ) , .A2( u2_u13_u0_n110 ) , .ZN( u2_u13_u0_n111 ) , .B1( u2_u13_u0_n118 ) , .A1( u2_u13_u0_n160 ) );
  INV_X1 u2_u13_u0_U31 (.A( u2_u13_u0_n118 ) , .ZN( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U32 (.ZN( u2_u13_u0_n104 ) , .B1( u2_u13_u0_n107 ) , .B2( u2_u13_u0_n141 ) , .A( u2_u13_u0_n144 ) );
  AOI21_X1 u2_u13_u0_U33 (.B1( u2_u13_u0_n127 ) , .B2( u2_u13_u0_n129 ) , .A( u2_u13_u0_n138 ) , .ZN( u2_u13_u0_n96 ) );
  AOI21_X1 u2_u13_u0_U34 (.ZN( u2_u13_u0_n116 ) , .B2( u2_u13_u0_n142 ) , .A( u2_u13_u0_n144 ) , .B1( u2_u13_u0_n166 ) );
  NAND2_X1 u2_u13_u0_U35 (.A1( u2_u13_u0_n100 ) , .A2( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n125 ) );
  NAND2_X1 u2_u13_u0_U36 (.A1( u2_u13_u0_n101 ) , .A2( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n150 ) );
  INV_X1 u2_u13_u0_U37 (.A( u2_u13_u0_n138 ) , .ZN( u2_u13_u0_n160 ) );
  NAND2_X1 u2_u13_u0_U38 (.A1( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n128 ) , .A2( u2_u13_u0_n95 ) );
  NAND2_X1 u2_u13_u0_U39 (.A1( u2_u13_u0_n100 ) , .ZN( u2_u13_u0_n129 ) , .A2( u2_u13_u0_n95 ) );
  AOI21_X1 u2_u13_u0_U4 (.B1( u2_u13_u0_n114 ) , .ZN( u2_u13_u0_n115 ) , .B2( u2_u13_u0_n129 ) , .A( u2_u13_u0_n161 ) );
  NAND2_X1 u2_u13_u0_U40 (.A2( u2_u13_u0_n100 ) , .ZN( u2_u13_u0_n131 ) , .A1( u2_u13_u0_n92 ) );
  NAND2_X1 u2_u13_u0_U41 (.A2( u2_u13_u0_n100 ) , .A1( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n139 ) );
  NAND2_X1 u2_u13_u0_U42 (.ZN( u2_u13_u0_n148 ) , .A1( u2_u13_u0_n93 ) , .A2( u2_u13_u0_n95 ) );
  NAND2_X1 u2_u13_u0_U43 (.A2( u2_u13_u0_n102 ) , .A1( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n149 ) );
  NAND2_X1 u2_u13_u0_U44 (.A2( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n114 ) , .A1( u2_u13_u0_n92 ) );
  NAND2_X1 u2_u13_u0_U45 (.A2( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n121 ) , .A1( u2_u13_u0_n93 ) );
  NAND2_X1 u2_u13_u0_U46 (.ZN( u2_u13_u0_n112 ) , .A2( u2_u13_u0_n92 ) , .A1( u2_u13_u0_n93 ) );
  OR3_X1 u2_u13_u0_U47 (.A3( u2_u13_u0_n152 ) , .A2( u2_u13_u0_n153 ) , .A1( u2_u13_u0_n154 ) , .ZN( u2_u13_u0_n155 ) );
  AOI21_X1 u2_u13_u0_U48 (.B2( u2_u13_u0_n150 ) , .B1( u2_u13_u0_n151 ) , .ZN( u2_u13_u0_n152 ) , .A( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U49 (.A( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n145 ) , .B1( u2_u13_u0_n146 ) , .ZN( u2_u13_u0_n154 ) );
  AOI21_X1 u2_u13_u0_U5 (.B2( u2_u13_u0_n131 ) , .ZN( u2_u13_u0_n134 ) , .B1( u2_u13_u0_n151 ) , .A( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U50 (.A( u2_u13_u0_n147 ) , .B2( u2_u13_u0_n148 ) , .B1( u2_u13_u0_n149 ) , .ZN( u2_u13_u0_n153 ) );
  INV_X1 u2_u13_u0_U51 (.ZN( u2_u13_u0_n171 ) , .A( u2_u13_u0_n99 ) );
  OAI211_X1 u2_u13_u0_U52 (.C2( u2_u13_u0_n140 ) , .C1( u2_u13_u0_n161 ) , .A( u2_u13_u0_n169 ) , .B( u2_u13_u0_n98 ) , .ZN( u2_u13_u0_n99 ) );
  INV_X1 u2_u13_u0_U53 (.ZN( u2_u13_u0_n169 ) , .A( u2_u13_u0_n91 ) );
  AOI211_X1 u2_u13_u0_U54 (.C1( u2_u13_u0_n118 ) , .A( u2_u13_u0_n123 ) , .B( u2_u13_u0_n96 ) , .C2( u2_u13_u0_n97 ) , .ZN( u2_u13_u0_n98 ) );
  NOR2_X1 u2_u13_u0_U55 (.A2( u2_u13_X_6 ) , .ZN( u2_u13_u0_n100 ) , .A1( u2_u13_u0_n162 ) );
  NOR2_X1 u2_u13_u0_U56 (.A2( u2_u13_X_4 ) , .A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n118 ) );
  NOR2_X1 u2_u13_u0_U57 (.A2( u2_u13_X_2 ) , .ZN( u2_u13_u0_n103 ) , .A1( u2_u13_u0_n164 ) );
  NOR2_X1 u2_u13_u0_U58 (.A2( u2_u13_X_1 ) , .A1( u2_u13_X_2 ) , .ZN( u2_u13_u0_n92 ) );
  NOR2_X1 u2_u13_u0_U59 (.A2( u2_u13_X_1 ) , .ZN( u2_u13_u0_n101 ) , .A1( u2_u13_u0_n163 ) );
  NOR2_X1 u2_u13_u0_U6 (.A1( u2_u13_u0_n108 ) , .ZN( u2_u13_u0_n123 ) , .A2( u2_u13_u0_n158 ) );
  NAND2_X1 u2_u13_u0_U60 (.A2( u2_u13_X_4 ) , .A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n144 ) );
  NOR2_X1 u2_u13_u0_U61 (.A2( u2_u13_X_5 ) , .ZN( u2_u13_u0_n136 ) , .A1( u2_u13_u0_n159 ) );
  NAND2_X1 u2_u13_u0_U62 (.A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n138 ) , .A2( u2_u13_u0_n159 ) );
  NOR2_X1 u2_u13_u0_U63 (.A2( u2_u13_X_3 ) , .A1( u2_u13_X_6 ) , .ZN( u2_u13_u0_n94 ) );
  AND2_X1 u2_u13_u0_U64 (.A2( u2_u13_X_3 ) , .A1( u2_u13_X_6 ) , .ZN( u2_u13_u0_n102 ) );
  AND2_X1 u2_u13_u0_U65 (.A1( u2_u13_X_6 ) , .A2( u2_u13_u0_n162 ) , .ZN( u2_u13_u0_n93 ) );
  INV_X1 u2_u13_u0_U66 (.A( u2_u13_X_4 ) , .ZN( u2_u13_u0_n159 ) );
  INV_X1 u2_u13_u0_U67 (.A( u2_u13_X_1 ) , .ZN( u2_u13_u0_n164 ) );
  INV_X1 u2_u13_u0_U68 (.A( u2_u13_X_2 ) , .ZN( u2_u13_u0_n163 ) );
  INV_X1 u2_u13_u0_U69 (.A( u2_u13_X_3 ) , .ZN( u2_u13_u0_n162 ) );
  OAI21_X1 u2_u13_u0_U7 (.B1( u2_u13_u0_n150 ) , .B2( u2_u13_u0_n158 ) , .A( u2_u13_u0_n172 ) , .ZN( u2_u13_u0_n89 ) );
  INV_X1 u2_u13_u0_U70 (.A( u2_u13_u0_n126 ) , .ZN( u2_u13_u0_n168 ) );
  AOI211_X1 u2_u13_u0_U71 (.B( u2_u13_u0_n133 ) , .A( u2_u13_u0_n134 ) , .C2( u2_u13_u0_n135 ) , .C1( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n137 ) );
  INV_X1 u2_u13_u0_U72 (.ZN( u2_u13_u0_n174 ) , .A( u2_u13_u0_n89 ) );
  AOI211_X1 u2_u13_u0_U73 (.B( u2_u13_u0_n104 ) , .A( u2_u13_u0_n105 ) , .ZN( u2_u13_u0_n106 ) , .C2( u2_u13_u0_n113 ) , .C1( u2_u13_u0_n160 ) );
  OR4_X1 u2_u13_u0_U74 (.ZN( u2_out13_17 ) , .A4( u2_u13_u0_n122 ) , .A2( u2_u13_u0_n123 ) , .A1( u2_u13_u0_n124 ) , .A3( u2_u13_u0_n170 ) );
  AOI21_X1 u2_u13_u0_U75 (.B2( u2_u13_u0_n107 ) , .ZN( u2_u13_u0_n124 ) , .B1( u2_u13_u0_n128 ) , .A( u2_u13_u0_n161 ) );
  INV_X1 u2_u13_u0_U76 (.A( u2_u13_u0_n111 ) , .ZN( u2_u13_u0_n170 ) );
  OR4_X1 u2_u13_u0_U77 (.ZN( u2_out13_31 ) , .A4( u2_u13_u0_n155 ) , .A2( u2_u13_u0_n156 ) , .A1( u2_u13_u0_n157 ) , .A3( u2_u13_u0_n173 ) );
  AOI21_X1 u2_u13_u0_U78 (.A( u2_u13_u0_n138 ) , .B2( u2_u13_u0_n139 ) , .B1( u2_u13_u0_n140 ) , .ZN( u2_u13_u0_n157 ) );
  AOI21_X1 u2_u13_u0_U79 (.B2( u2_u13_u0_n141 ) , .B1( u2_u13_u0_n142 ) , .ZN( u2_u13_u0_n156 ) , .A( u2_u13_u0_n161 ) );
  AND2_X1 u2_u13_u0_U8 (.A1( u2_u13_u0_n114 ) , .A2( u2_u13_u0_n121 ) , .ZN( u2_u13_u0_n146 ) );
  AOI21_X1 u2_u13_u0_U80 (.B1( u2_u13_u0_n132 ) , .ZN( u2_u13_u0_n133 ) , .A( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n166 ) );
  OAI22_X1 u2_u13_u0_U81 (.ZN( u2_u13_u0_n105 ) , .A2( u2_u13_u0_n132 ) , .B1( u2_u13_u0_n146 ) , .A1( u2_u13_u0_n147 ) , .B2( u2_u13_u0_n161 ) );
  NAND2_X1 u2_u13_u0_U82 (.ZN( u2_u13_u0_n110 ) , .A2( u2_u13_u0_n132 ) , .A1( u2_u13_u0_n145 ) );
  INV_X1 u2_u13_u0_U83 (.A( u2_u13_u0_n119 ) , .ZN( u2_u13_u0_n167 ) );
  NAND2_X1 u2_u13_u0_U84 (.A2( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n140 ) , .A1( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U85 (.A1( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n130 ) , .A2( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U86 (.ZN( u2_u13_u0_n108 ) , .A1( u2_u13_u0_n92 ) , .A2( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U87 (.ZN( u2_u13_u0_n142 ) , .A1( u2_u13_u0_n94 ) , .A2( u2_u13_u0_n95 ) );
  NAND3_X1 u2_u13_u0_U88 (.ZN( u2_out13_23 ) , .A3( u2_u13_u0_n137 ) , .A1( u2_u13_u0_n168 ) , .A2( u2_u13_u0_n171 ) );
  NAND3_X1 u2_u13_u0_U89 (.A3( u2_u13_u0_n127 ) , .A2( u2_u13_u0_n128 ) , .ZN( u2_u13_u0_n135 ) , .A1( u2_u13_u0_n150 ) );
  AND2_X1 u2_u13_u0_U9 (.A1( u2_u13_u0_n131 ) , .ZN( u2_u13_u0_n141 ) , .A2( u2_u13_u0_n150 ) );
  NAND3_X1 u2_u13_u0_U90 (.ZN( u2_u13_u0_n117 ) , .A3( u2_u13_u0_n132 ) , .A2( u2_u13_u0_n139 ) , .A1( u2_u13_u0_n148 ) );
  NAND3_X1 u2_u13_u0_U91 (.ZN( u2_u13_u0_n109 ) , .A2( u2_u13_u0_n114 ) , .A3( u2_u13_u0_n140 ) , .A1( u2_u13_u0_n149 ) );
  NAND3_X1 u2_u13_u0_U92 (.ZN( u2_out13_9 ) , .A3( u2_u13_u0_n106 ) , .A2( u2_u13_u0_n171 ) , .A1( u2_u13_u0_n174 ) );
  NAND3_X1 u2_u13_u0_U93 (.A2( u2_u13_u0_n128 ) , .A1( u2_u13_u0_n132 ) , .A3( u2_u13_u0_n146 ) , .ZN( u2_u13_u0_n97 ) );
  AOI21_X1 u2_u13_u1_U10 (.B2( u2_u13_u1_n155 ) , .B1( u2_u13_u1_n156 ) , .ZN( u2_u13_u1_n157 ) , .A( u2_u13_u1_n174 ) );
  NAND3_X1 u2_u13_u1_U100 (.ZN( u2_u13_u1_n113 ) , .A1( u2_u13_u1_n120 ) , .A3( u2_u13_u1_n133 ) , .A2( u2_u13_u1_n155 ) );
  NAND2_X1 u2_u13_u1_U11 (.ZN( u2_u13_u1_n140 ) , .A2( u2_u13_u1_n150 ) , .A1( u2_u13_u1_n155 ) );
  NAND2_X1 u2_u13_u1_U12 (.A1( u2_u13_u1_n131 ) , .ZN( u2_u13_u1_n147 ) , .A2( u2_u13_u1_n153 ) );
  INV_X1 u2_u13_u1_U13 (.A( u2_u13_u1_n139 ) , .ZN( u2_u13_u1_n174 ) );
  OR4_X1 u2_u13_u1_U14 (.A4( u2_u13_u1_n106 ) , .A3( u2_u13_u1_n107 ) , .ZN( u2_u13_u1_n108 ) , .A1( u2_u13_u1_n117 ) , .A2( u2_u13_u1_n184 ) );
  AOI21_X1 u2_u13_u1_U15 (.ZN( u2_u13_u1_n106 ) , .A( u2_u13_u1_n112 ) , .B1( u2_u13_u1_n154 ) , .B2( u2_u13_u1_n156 ) );
  AOI21_X1 u2_u13_u1_U16 (.ZN( u2_u13_u1_n107 ) , .B1( u2_u13_u1_n134 ) , .B2( u2_u13_u1_n149 ) , .A( u2_u13_u1_n174 ) );
  INV_X1 u2_u13_u1_U17 (.A( u2_u13_u1_n101 ) , .ZN( u2_u13_u1_n184 ) );
  INV_X1 u2_u13_u1_U18 (.A( u2_u13_u1_n112 ) , .ZN( u2_u13_u1_n171 ) );
  NAND2_X1 u2_u13_u1_U19 (.ZN( u2_u13_u1_n141 ) , .A1( u2_u13_u1_n153 ) , .A2( u2_u13_u1_n156 ) );
  AND2_X1 u2_u13_u1_U20 (.A1( u2_u13_u1_n123 ) , .ZN( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n161 ) );
  NAND2_X1 u2_u13_u1_U21 (.A2( u2_u13_u1_n115 ) , .A1( u2_u13_u1_n116 ) , .ZN( u2_u13_u1_n148 ) );
  NAND2_X1 u2_u13_u1_U22 (.A2( u2_u13_u1_n133 ) , .A1( u2_u13_u1_n135 ) , .ZN( u2_u13_u1_n159 ) );
  NAND2_X1 u2_u13_u1_U23 (.A2( u2_u13_u1_n115 ) , .A1( u2_u13_u1_n120 ) , .ZN( u2_u13_u1_n132 ) );
  INV_X1 u2_u13_u1_U24 (.A( u2_u13_u1_n154 ) , .ZN( u2_u13_u1_n178 ) );
  AOI22_X1 u2_u13_u1_U25 (.B2( u2_u13_u1_n113 ) , .A2( u2_u13_u1_n114 ) , .ZN( u2_u13_u1_n125 ) , .A1( u2_u13_u1_n171 ) , .B1( u2_u13_u1_n173 ) );
  NAND2_X1 u2_u13_u1_U26 (.ZN( u2_u13_u1_n114 ) , .A1( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n156 ) );
  INV_X1 u2_u13_u1_U27 (.A( u2_u13_u1_n151 ) , .ZN( u2_u13_u1_n183 ) );
  AND2_X1 u2_u13_u1_U28 (.A1( u2_u13_u1_n129 ) , .A2( u2_u13_u1_n133 ) , .ZN( u2_u13_u1_n149 ) );
  INV_X1 u2_u13_u1_U29 (.A( u2_u13_u1_n131 ) , .ZN( u2_u13_u1_n180 ) );
  INV_X1 u2_u13_u1_U3 (.A( u2_u13_u1_n159 ) , .ZN( u2_u13_u1_n182 ) );
  OAI221_X1 u2_u13_u1_U30 (.A( u2_u13_u1_n119 ) , .C2( u2_u13_u1_n129 ) , .ZN( u2_u13_u1_n138 ) , .B2( u2_u13_u1_n152 ) , .C1( u2_u13_u1_n174 ) , .B1( u2_u13_u1_n187 ) );
  INV_X1 u2_u13_u1_U31 (.A( u2_u13_u1_n148 ) , .ZN( u2_u13_u1_n187 ) );
  AOI211_X1 u2_u13_u1_U32 (.B( u2_u13_u1_n117 ) , .A( u2_u13_u1_n118 ) , .ZN( u2_u13_u1_n119 ) , .C2( u2_u13_u1_n146 ) , .C1( u2_u13_u1_n159 ) );
  NOR2_X1 u2_u13_u1_U33 (.A1( u2_u13_u1_n168 ) , .A2( u2_u13_u1_n176 ) , .ZN( u2_u13_u1_n98 ) );
  AOI211_X1 u2_u13_u1_U34 (.B( u2_u13_u1_n162 ) , .A( u2_u13_u1_n163 ) , .C2( u2_u13_u1_n164 ) , .ZN( u2_u13_u1_n165 ) , .C1( u2_u13_u1_n171 ) );
  AOI21_X1 u2_u13_u1_U35 (.A( u2_u13_u1_n160 ) , .B2( u2_u13_u1_n161 ) , .ZN( u2_u13_u1_n162 ) , .B1( u2_u13_u1_n182 ) );
  OR2_X1 u2_u13_u1_U36 (.A2( u2_u13_u1_n157 ) , .A1( u2_u13_u1_n158 ) , .ZN( u2_u13_u1_n163 ) );
  OAI21_X1 u2_u13_u1_U37 (.B2( u2_u13_u1_n123 ) , .ZN( u2_u13_u1_n145 ) , .B1( u2_u13_u1_n160 ) , .A( u2_u13_u1_n185 ) );
  INV_X1 u2_u13_u1_U38 (.A( u2_u13_u1_n122 ) , .ZN( u2_u13_u1_n185 ) );
  AOI21_X1 u2_u13_u1_U39 (.B2( u2_u13_u1_n120 ) , .B1( u2_u13_u1_n121 ) , .ZN( u2_u13_u1_n122 ) , .A( u2_u13_u1_n128 ) );
  AOI221_X1 u2_u13_u1_U4 (.A( u2_u13_u1_n138 ) , .C2( u2_u13_u1_n139 ) , .C1( u2_u13_u1_n140 ) , .B2( u2_u13_u1_n141 ) , .ZN( u2_u13_u1_n142 ) , .B1( u2_u13_u1_n175 ) );
  NAND2_X1 u2_u13_u1_U40 (.A1( u2_u13_u1_n128 ) , .ZN( u2_u13_u1_n146 ) , .A2( u2_u13_u1_n160 ) );
  NAND2_X1 u2_u13_u1_U41 (.A2( u2_u13_u1_n112 ) , .ZN( u2_u13_u1_n139 ) , .A1( u2_u13_u1_n152 ) );
  NAND2_X1 u2_u13_u1_U42 (.A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n156 ) , .A2( u2_u13_u1_n99 ) );
  AOI221_X1 u2_u13_u1_U43 (.B1( u2_u13_u1_n140 ) , .ZN( u2_u13_u1_n167 ) , .B2( u2_u13_u1_n172 ) , .C2( u2_u13_u1_n175 ) , .C1( u2_u13_u1_n178 ) , .A( u2_u13_u1_n188 ) );
  INV_X1 u2_u13_u1_U44 (.ZN( u2_u13_u1_n188 ) , .A( u2_u13_u1_n97 ) );
  AOI211_X1 u2_u13_u1_U45 (.A( u2_u13_u1_n118 ) , .C1( u2_u13_u1_n132 ) , .C2( u2_u13_u1_n139 ) , .B( u2_u13_u1_n96 ) , .ZN( u2_u13_u1_n97 ) );
  AOI21_X1 u2_u13_u1_U46 (.B2( u2_u13_u1_n121 ) , .B1( u2_u13_u1_n135 ) , .A( u2_u13_u1_n152 ) , .ZN( u2_u13_u1_n96 ) );
  NOR2_X1 u2_u13_u1_U47 (.ZN( u2_u13_u1_n117 ) , .A1( u2_u13_u1_n121 ) , .A2( u2_u13_u1_n160 ) );
  AOI21_X1 u2_u13_u1_U48 (.A( u2_u13_u1_n128 ) , .B2( u2_u13_u1_n129 ) , .ZN( u2_u13_u1_n130 ) , .B1( u2_u13_u1_n150 ) );
  NAND2_X1 u2_u13_u1_U49 (.ZN( u2_u13_u1_n112 ) , .A1( u2_u13_u1_n169 ) , .A2( u2_u13_u1_n170 ) );
  AOI211_X1 u2_u13_u1_U5 (.ZN( u2_u13_u1_n124 ) , .A( u2_u13_u1_n138 ) , .C2( u2_u13_u1_n139 ) , .B( u2_u13_u1_n145 ) , .C1( u2_u13_u1_n147 ) );
  NAND2_X1 u2_u13_u1_U50 (.ZN( u2_u13_u1_n129 ) , .A2( u2_u13_u1_n95 ) , .A1( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U51 (.A1( u2_u13_u1_n102 ) , .ZN( u2_u13_u1_n154 ) , .A2( u2_u13_u1_n99 ) );
  NAND2_X1 u2_u13_u1_U52 (.A2( u2_u13_u1_n100 ) , .ZN( u2_u13_u1_n135 ) , .A1( u2_u13_u1_n99 ) );
  AOI21_X1 u2_u13_u1_U53 (.A( u2_u13_u1_n152 ) , .B2( u2_u13_u1_n153 ) , .B1( u2_u13_u1_n154 ) , .ZN( u2_u13_u1_n158 ) );
  INV_X1 u2_u13_u1_U54 (.A( u2_u13_u1_n160 ) , .ZN( u2_u13_u1_n175 ) );
  NAND2_X1 u2_u13_u1_U55 (.A1( u2_u13_u1_n100 ) , .ZN( u2_u13_u1_n116 ) , .A2( u2_u13_u1_n95 ) );
  NAND2_X1 u2_u13_u1_U56 (.A1( u2_u13_u1_n102 ) , .ZN( u2_u13_u1_n131 ) , .A2( u2_u13_u1_n95 ) );
  NAND2_X1 u2_u13_u1_U57 (.A2( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n121 ) , .A1( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U58 (.A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n153 ) , .A2( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U59 (.A2( u2_u13_u1_n104 ) , .A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n133 ) );
  AOI22_X1 u2_u13_u1_U6 (.B2( u2_u13_u1_n136 ) , .A2( u2_u13_u1_n137 ) , .ZN( u2_u13_u1_n143 ) , .A1( u2_u13_u1_n171 ) , .B1( u2_u13_u1_n173 ) );
  NAND2_X1 u2_u13_u1_U60 (.ZN( u2_u13_u1_n150 ) , .A2( u2_u13_u1_n98 ) , .A1( u2_u13_u1_n99 ) );
  NAND2_X1 u2_u13_u1_U61 (.A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n155 ) , .A2( u2_u13_u1_n95 ) );
  OAI21_X1 u2_u13_u1_U62 (.ZN( u2_u13_u1_n109 ) , .B1( u2_u13_u1_n129 ) , .B2( u2_u13_u1_n160 ) , .A( u2_u13_u1_n167 ) );
  NAND2_X1 u2_u13_u1_U63 (.A2( u2_u13_u1_n100 ) , .A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n120 ) );
  NAND2_X1 u2_u13_u1_U64 (.A1( u2_u13_u1_n102 ) , .A2( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n115 ) );
  NAND2_X1 u2_u13_u1_U65 (.A2( u2_u13_u1_n100 ) , .A1( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n151 ) );
  NAND2_X1 u2_u13_u1_U66 (.A2( u2_u13_u1_n103 ) , .A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n161 ) );
  INV_X1 u2_u13_u1_U67 (.A( u2_u13_u1_n152 ) , .ZN( u2_u13_u1_n173 ) );
  INV_X1 u2_u13_u1_U68 (.A( u2_u13_u1_n128 ) , .ZN( u2_u13_u1_n172 ) );
  NAND2_X1 u2_u13_u1_U69 (.A2( u2_u13_u1_n102 ) , .A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n123 ) );
  INV_X1 u2_u13_u1_U7 (.A( u2_u13_u1_n147 ) , .ZN( u2_u13_u1_n181 ) );
  NOR2_X1 u2_u13_u1_U70 (.A2( u2_u13_X_7 ) , .A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n95 ) );
  NOR2_X1 u2_u13_u1_U71 (.A1( u2_u13_X_12 ) , .A2( u2_u13_X_9 ) , .ZN( u2_u13_u1_n100 ) );
  NOR2_X1 u2_u13_u1_U72 (.A2( u2_u13_X_8 ) , .A1( u2_u13_u1_n177 ) , .ZN( u2_u13_u1_n99 ) );
  NOR2_X1 u2_u13_u1_U73 (.A2( u2_u13_X_12 ) , .ZN( u2_u13_u1_n102 ) , .A1( u2_u13_u1_n176 ) );
  NOR2_X1 u2_u13_u1_U74 (.A2( u2_u13_X_9 ) , .ZN( u2_u13_u1_n105 ) , .A1( u2_u13_u1_n168 ) );
  NAND2_X1 u2_u13_u1_U75 (.A1( u2_u13_X_10 ) , .ZN( u2_u13_u1_n160 ) , .A2( u2_u13_u1_n169 ) );
  NAND2_X1 u2_u13_u1_U76 (.A2( u2_u13_X_10 ) , .A1( u2_u13_X_11 ) , .ZN( u2_u13_u1_n152 ) );
  NAND2_X1 u2_u13_u1_U77 (.A1( u2_u13_X_11 ) , .ZN( u2_u13_u1_n128 ) , .A2( u2_u13_u1_n170 ) );
  AND2_X1 u2_u13_u1_U78 (.A2( u2_u13_X_7 ) , .A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n104 ) );
  AND2_X1 u2_u13_u1_U79 (.A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n103 ) , .A2( u2_u13_u1_n177 ) );
  NOR2_X1 u2_u13_u1_U8 (.A1( u2_u13_u1_n112 ) , .A2( u2_u13_u1_n116 ) , .ZN( u2_u13_u1_n118 ) );
  INV_X1 u2_u13_u1_U80 (.A( u2_u13_X_10 ) , .ZN( u2_u13_u1_n170 ) );
  INV_X1 u2_u13_u1_U81 (.A( u2_u13_X_9 ) , .ZN( u2_u13_u1_n176 ) );
  INV_X1 u2_u13_u1_U82 (.A( u2_u13_X_11 ) , .ZN( u2_u13_u1_n169 ) );
  INV_X1 u2_u13_u1_U83 (.A( u2_u13_X_12 ) , .ZN( u2_u13_u1_n168 ) );
  INV_X1 u2_u13_u1_U84 (.A( u2_u13_X_7 ) , .ZN( u2_u13_u1_n177 ) );
  NAND4_X1 u2_u13_u1_U85 (.ZN( u2_out13_28 ) , .A4( u2_u13_u1_n124 ) , .A3( u2_u13_u1_n125 ) , .A2( u2_u13_u1_n126 ) , .A1( u2_u13_u1_n127 ) );
  OAI21_X1 u2_u13_u1_U86 (.ZN( u2_u13_u1_n127 ) , .B2( u2_u13_u1_n139 ) , .B1( u2_u13_u1_n175 ) , .A( u2_u13_u1_n183 ) );
  OAI21_X1 u2_u13_u1_U87 (.ZN( u2_u13_u1_n126 ) , .B2( u2_u13_u1_n140 ) , .A( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n178 ) );
  NAND4_X1 u2_u13_u1_U88 (.ZN( u2_out13_18 ) , .A4( u2_u13_u1_n165 ) , .A3( u2_u13_u1_n166 ) , .A1( u2_u13_u1_n167 ) , .A2( u2_u13_u1_n186 ) );
  AOI22_X1 u2_u13_u1_U89 (.B2( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n147 ) , .A2( u2_u13_u1_n148 ) , .ZN( u2_u13_u1_n166 ) , .A1( u2_u13_u1_n172 ) );
  OAI21_X1 u2_u13_u1_U9 (.ZN( u2_u13_u1_n101 ) , .B1( u2_u13_u1_n141 ) , .A( u2_u13_u1_n146 ) , .B2( u2_u13_u1_n183 ) );
  INV_X1 u2_u13_u1_U90 (.A( u2_u13_u1_n145 ) , .ZN( u2_u13_u1_n186 ) );
  NAND4_X1 u2_u13_u1_U91 (.ZN( u2_out13_2 ) , .A4( u2_u13_u1_n142 ) , .A3( u2_u13_u1_n143 ) , .A2( u2_u13_u1_n144 ) , .A1( u2_u13_u1_n179 ) );
  OAI21_X1 u2_u13_u1_U92 (.B2( u2_u13_u1_n132 ) , .ZN( u2_u13_u1_n144 ) , .A( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n180 ) );
  INV_X1 u2_u13_u1_U93 (.A( u2_u13_u1_n130 ) , .ZN( u2_u13_u1_n179 ) );
  OR4_X1 u2_u13_u1_U94 (.ZN( u2_out13_13 ) , .A4( u2_u13_u1_n108 ) , .A3( u2_u13_u1_n109 ) , .A2( u2_u13_u1_n110 ) , .A1( u2_u13_u1_n111 ) );
  AOI21_X1 u2_u13_u1_U95 (.ZN( u2_u13_u1_n111 ) , .A( u2_u13_u1_n128 ) , .B2( u2_u13_u1_n131 ) , .B1( u2_u13_u1_n135 ) );
  AOI21_X1 u2_u13_u1_U96 (.ZN( u2_u13_u1_n110 ) , .A( u2_u13_u1_n116 ) , .B1( u2_u13_u1_n152 ) , .B2( u2_u13_u1_n160 ) );
  NAND3_X1 u2_u13_u1_U97 (.A3( u2_u13_u1_n149 ) , .A2( u2_u13_u1_n150 ) , .A1( u2_u13_u1_n151 ) , .ZN( u2_u13_u1_n164 ) );
  NAND3_X1 u2_u13_u1_U98 (.A3( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n135 ) , .ZN( u2_u13_u1_n136 ) , .A1( u2_u13_u1_n151 ) );
  NAND3_X1 u2_u13_u1_U99 (.A1( u2_u13_u1_n133 ) , .ZN( u2_u13_u1_n137 ) , .A2( u2_u13_u1_n154 ) , .A3( u2_u13_u1_n181 ) );
  OAI22_X1 u2_u13_u2_U10 (.B1( u2_u13_u2_n151 ) , .A2( u2_u13_u2_n152 ) , .A1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n160 ) , .B2( u2_u13_u2_n168 ) );
  NAND3_X1 u2_u13_u2_U100 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n98 ) );
  NOR3_X1 u2_u13_u2_U11 (.A1( u2_u13_u2_n150 ) , .ZN( u2_u13_u2_n151 ) , .A3( u2_u13_u2_n175 ) , .A2( u2_u13_u2_n188 ) );
  AOI21_X1 u2_u13_u2_U12 (.B2( u2_u13_u2_n123 ) , .ZN( u2_u13_u2_n125 ) , .A( u2_u13_u2_n171 ) , .B1( u2_u13_u2_n184 ) );
  INV_X1 u2_u13_u2_U13 (.A( u2_u13_u2_n150 ) , .ZN( u2_u13_u2_n184 ) );
  AOI21_X1 u2_u13_u2_U14 (.ZN( u2_u13_u2_n144 ) , .B2( u2_u13_u2_n155 ) , .A( u2_u13_u2_n172 ) , .B1( u2_u13_u2_n185 ) );
  AOI21_X1 u2_u13_u2_U15 (.B2( u2_u13_u2_n143 ) , .ZN( u2_u13_u2_n145 ) , .B1( u2_u13_u2_n152 ) , .A( u2_u13_u2_n171 ) );
  INV_X1 u2_u13_u2_U16 (.A( u2_u13_u2_n156 ) , .ZN( u2_u13_u2_n171 ) );
  INV_X1 u2_u13_u2_U17 (.A( u2_u13_u2_n120 ) , .ZN( u2_u13_u2_n188 ) );
  NAND2_X1 u2_u13_u2_U18 (.A2( u2_u13_u2_n122 ) , .ZN( u2_u13_u2_n150 ) , .A1( u2_u13_u2_n152 ) );
  INV_X1 u2_u13_u2_U19 (.A( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n170 ) );
  INV_X1 u2_u13_u2_U20 (.A( u2_u13_u2_n137 ) , .ZN( u2_u13_u2_n173 ) );
  NAND2_X1 u2_u13_u2_U21 (.A1( u2_u13_u2_n132 ) , .A2( u2_u13_u2_n139 ) , .ZN( u2_u13_u2_n157 ) );
  INV_X1 u2_u13_u2_U22 (.A( u2_u13_u2_n113 ) , .ZN( u2_u13_u2_n178 ) );
  INV_X1 u2_u13_u2_U23 (.A( u2_u13_u2_n139 ) , .ZN( u2_u13_u2_n175 ) );
  INV_X1 u2_u13_u2_U24 (.A( u2_u13_u2_n155 ) , .ZN( u2_u13_u2_n181 ) );
  INV_X1 u2_u13_u2_U25 (.A( u2_u13_u2_n119 ) , .ZN( u2_u13_u2_n177 ) );
  INV_X1 u2_u13_u2_U26 (.A( u2_u13_u2_n116 ) , .ZN( u2_u13_u2_n180 ) );
  INV_X1 u2_u13_u2_U27 (.A( u2_u13_u2_n131 ) , .ZN( u2_u13_u2_n179 ) );
  INV_X1 u2_u13_u2_U28 (.A( u2_u13_u2_n154 ) , .ZN( u2_u13_u2_n176 ) );
  NAND2_X1 u2_u13_u2_U29 (.A2( u2_u13_u2_n116 ) , .A1( u2_u13_u2_n117 ) , .ZN( u2_u13_u2_n118 ) );
  NOR2_X1 u2_u13_u2_U3 (.ZN( u2_u13_u2_n121 ) , .A2( u2_u13_u2_n177 ) , .A1( u2_u13_u2_n180 ) );
  INV_X1 u2_u13_u2_U30 (.A( u2_u13_u2_n132 ) , .ZN( u2_u13_u2_n182 ) );
  INV_X1 u2_u13_u2_U31 (.A( u2_u13_u2_n158 ) , .ZN( u2_u13_u2_n183 ) );
  OAI21_X1 u2_u13_u2_U32 (.A( u2_u13_u2_n156 ) , .B1( u2_u13_u2_n157 ) , .ZN( u2_u13_u2_n158 ) , .B2( u2_u13_u2_n179 ) );
  NOR2_X1 u2_u13_u2_U33 (.ZN( u2_u13_u2_n156 ) , .A1( u2_u13_u2_n166 ) , .A2( u2_u13_u2_n169 ) );
  NOR2_X1 u2_u13_u2_U34 (.A2( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n137 ) , .A1( u2_u13_u2_n140 ) );
  NOR2_X1 u2_u13_u2_U35 (.A2( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n153 ) , .A1( u2_u13_u2_n156 ) );
  AOI211_X1 u2_u13_u2_U36 (.ZN( u2_u13_u2_n130 ) , .C1( u2_u13_u2_n138 ) , .C2( u2_u13_u2_n179 ) , .B( u2_u13_u2_n96 ) , .A( u2_u13_u2_n97 ) );
  OAI22_X1 u2_u13_u2_U37 (.B1( u2_u13_u2_n133 ) , .A2( u2_u13_u2_n137 ) , .A1( u2_u13_u2_n152 ) , .B2( u2_u13_u2_n168 ) , .ZN( u2_u13_u2_n97 ) );
  OAI221_X1 u2_u13_u2_U38 (.B1( u2_u13_u2_n113 ) , .C1( u2_u13_u2_n132 ) , .A( u2_u13_u2_n149 ) , .B2( u2_u13_u2_n171 ) , .C2( u2_u13_u2_n172 ) , .ZN( u2_u13_u2_n96 ) );
  OAI221_X1 u2_u13_u2_U39 (.A( u2_u13_u2_n115 ) , .C2( u2_u13_u2_n123 ) , .B2( u2_u13_u2_n143 ) , .B1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n163 ) , .C1( u2_u13_u2_n168 ) );
  INV_X1 u2_u13_u2_U4 (.A( u2_u13_u2_n134 ) , .ZN( u2_u13_u2_n185 ) );
  OAI21_X1 u2_u13_u2_U40 (.A( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n115 ) , .B1( u2_u13_u2_n176 ) , .B2( u2_u13_u2_n178 ) );
  OAI221_X1 u2_u13_u2_U41 (.A( u2_u13_u2_n135 ) , .B2( u2_u13_u2_n136 ) , .B1( u2_u13_u2_n137 ) , .ZN( u2_u13_u2_n162 ) , .C2( u2_u13_u2_n167 ) , .C1( u2_u13_u2_n185 ) );
  AND3_X1 u2_u13_u2_U42 (.A3( u2_u13_u2_n131 ) , .A2( u2_u13_u2_n132 ) , .A1( u2_u13_u2_n133 ) , .ZN( u2_u13_u2_n136 ) );
  AOI22_X1 u2_u13_u2_U43 (.ZN( u2_u13_u2_n135 ) , .B1( u2_u13_u2_n140 ) , .A1( u2_u13_u2_n156 ) , .B2( u2_u13_u2_n180 ) , .A2( u2_u13_u2_n188 ) );
  AOI21_X1 u2_u13_u2_U44 (.ZN( u2_u13_u2_n149 ) , .B1( u2_u13_u2_n173 ) , .B2( u2_u13_u2_n188 ) , .A( u2_u13_u2_n95 ) );
  AND3_X1 u2_u13_u2_U45 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n156 ) , .ZN( u2_u13_u2_n95 ) );
  OAI21_X1 u2_u13_u2_U46 (.A( u2_u13_u2_n141 ) , .B2( u2_u13_u2_n142 ) , .ZN( u2_u13_u2_n146 ) , .B1( u2_u13_u2_n153 ) );
  OAI21_X1 u2_u13_u2_U47 (.A( u2_u13_u2_n140 ) , .ZN( u2_u13_u2_n141 ) , .B1( u2_u13_u2_n176 ) , .B2( u2_u13_u2_n177 ) );
  NOR3_X1 u2_u13_u2_U48 (.ZN( u2_u13_u2_n142 ) , .A3( u2_u13_u2_n175 ) , .A2( u2_u13_u2_n178 ) , .A1( u2_u13_u2_n181 ) );
  OAI21_X1 u2_u13_u2_U49 (.A( u2_u13_u2_n101 ) , .B2( u2_u13_u2_n121 ) , .B1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n164 ) );
  NOR4_X1 u2_u13_u2_U5 (.A4( u2_u13_u2_n124 ) , .A3( u2_u13_u2_n125 ) , .A2( u2_u13_u2_n126 ) , .A1( u2_u13_u2_n127 ) , .ZN( u2_u13_u2_n128 ) );
  NAND2_X1 u2_u13_u2_U50 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n155 ) );
  NAND2_X1 u2_u13_u2_U51 (.A2( u2_u13_u2_n105 ) , .A1( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n143 ) );
  NAND2_X1 u2_u13_u2_U52 (.A1( u2_u13_u2_n104 ) , .A2( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n152 ) );
  NAND2_X1 u2_u13_u2_U53 (.A1( u2_u13_u2_n100 ) , .A2( u2_u13_u2_n105 ) , .ZN( u2_u13_u2_n132 ) );
  INV_X1 u2_u13_u2_U54 (.A( u2_u13_u2_n140 ) , .ZN( u2_u13_u2_n168 ) );
  INV_X1 u2_u13_u2_U55 (.A( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n167 ) );
  NAND2_X1 u2_u13_u2_U56 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n113 ) );
  NAND2_X1 u2_u13_u2_U57 (.A1( u2_u13_u2_n106 ) , .A2( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n131 ) );
  NAND2_X1 u2_u13_u2_U58 (.A1( u2_u13_u2_n103 ) , .A2( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n139 ) );
  NAND2_X1 u2_u13_u2_U59 (.A1( u2_u13_u2_n103 ) , .A2( u2_u13_u2_n105 ) , .ZN( u2_u13_u2_n133 ) );
  AOI21_X1 u2_u13_u2_U6 (.B2( u2_u13_u2_n119 ) , .ZN( u2_u13_u2_n127 ) , .A( u2_u13_u2_n137 ) , .B1( u2_u13_u2_n155 ) );
  NAND2_X1 u2_u13_u2_U60 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n103 ) , .ZN( u2_u13_u2_n154 ) );
  NAND2_X1 u2_u13_u2_U61 (.A2( u2_u13_u2_n103 ) , .A1( u2_u13_u2_n104 ) , .ZN( u2_u13_u2_n119 ) );
  NAND2_X1 u2_u13_u2_U62 (.A2( u2_u13_u2_n107 ) , .A1( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n123 ) );
  NAND2_X1 u2_u13_u2_U63 (.A1( u2_u13_u2_n104 ) , .A2( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n122 ) );
  INV_X1 u2_u13_u2_U64 (.A( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n172 ) );
  NAND2_X1 u2_u13_u2_U65 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n102 ) , .ZN( u2_u13_u2_n116 ) );
  NAND2_X1 u2_u13_u2_U66 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n120 ) );
  NAND2_X1 u2_u13_u2_U67 (.A2( u2_u13_u2_n105 ) , .A1( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n117 ) );
  INV_X1 u2_u13_u2_U68 (.ZN( u2_u13_u2_n187 ) , .A( u2_u13_u2_n99 ) );
  OAI21_X1 u2_u13_u2_U69 (.B1( u2_u13_u2_n137 ) , .B2( u2_u13_u2_n143 ) , .A( u2_u13_u2_n98 ) , .ZN( u2_u13_u2_n99 ) );
  AOI21_X1 u2_u13_u2_U7 (.ZN( u2_u13_u2_n124 ) , .B1( u2_u13_u2_n131 ) , .B2( u2_u13_u2_n143 ) , .A( u2_u13_u2_n172 ) );
  NOR2_X1 u2_u13_u2_U70 (.A2( u2_u13_X_16 ) , .ZN( u2_u13_u2_n140 ) , .A1( u2_u13_u2_n166 ) );
  NOR2_X1 u2_u13_u2_U71 (.A2( u2_u13_X_13 ) , .A1( u2_u13_X_14 ) , .ZN( u2_u13_u2_n100 ) );
  NOR2_X1 u2_u13_u2_U72 (.A2( u2_u13_X_16 ) , .A1( u2_u13_X_17 ) , .ZN( u2_u13_u2_n138 ) );
  NOR2_X1 u2_u13_u2_U73 (.A2( u2_u13_X_15 ) , .A1( u2_u13_X_18 ) , .ZN( u2_u13_u2_n104 ) );
  NOR2_X1 u2_u13_u2_U74 (.A2( u2_u13_X_14 ) , .ZN( u2_u13_u2_n103 ) , .A1( u2_u13_u2_n174 ) );
  NOR2_X1 u2_u13_u2_U75 (.A2( u2_u13_X_15 ) , .ZN( u2_u13_u2_n102 ) , .A1( u2_u13_u2_n165 ) );
  NOR2_X1 u2_u13_u2_U76 (.A2( u2_u13_X_17 ) , .ZN( u2_u13_u2_n114 ) , .A1( u2_u13_u2_n169 ) );
  AND2_X1 u2_u13_u2_U77 (.A1( u2_u13_X_15 ) , .ZN( u2_u13_u2_n105 ) , .A2( u2_u13_u2_n165 ) );
  AND2_X1 u2_u13_u2_U78 (.A2( u2_u13_X_15 ) , .A1( u2_u13_X_18 ) , .ZN( u2_u13_u2_n107 ) );
  AND2_X1 u2_u13_u2_U79 (.A1( u2_u13_X_14 ) , .ZN( u2_u13_u2_n106 ) , .A2( u2_u13_u2_n174 ) );
  AOI21_X1 u2_u13_u2_U8 (.B2( u2_u13_u2_n120 ) , .B1( u2_u13_u2_n121 ) , .ZN( u2_u13_u2_n126 ) , .A( u2_u13_u2_n167 ) );
  AND2_X1 u2_u13_u2_U80 (.A1( u2_u13_X_13 ) , .A2( u2_u13_X_14 ) , .ZN( u2_u13_u2_n108 ) );
  INV_X1 u2_u13_u2_U81 (.A( u2_u13_X_16 ) , .ZN( u2_u13_u2_n169 ) );
  INV_X1 u2_u13_u2_U82 (.A( u2_u13_X_17 ) , .ZN( u2_u13_u2_n166 ) );
  INV_X1 u2_u13_u2_U83 (.A( u2_u13_X_13 ) , .ZN( u2_u13_u2_n174 ) );
  INV_X1 u2_u13_u2_U84 (.A( u2_u13_X_18 ) , .ZN( u2_u13_u2_n165 ) );
  NAND4_X1 u2_u13_u2_U85 (.ZN( u2_out13_30 ) , .A4( u2_u13_u2_n147 ) , .A3( u2_u13_u2_n148 ) , .A2( u2_u13_u2_n149 ) , .A1( u2_u13_u2_n187 ) );
  AOI21_X1 u2_u13_u2_U86 (.B2( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n148 ) , .A( u2_u13_u2_n162 ) , .B1( u2_u13_u2_n182 ) );
  NOR3_X1 u2_u13_u2_U87 (.A3( u2_u13_u2_n144 ) , .A2( u2_u13_u2_n145 ) , .A1( u2_u13_u2_n146 ) , .ZN( u2_u13_u2_n147 ) );
  NAND4_X1 u2_u13_u2_U88 (.ZN( u2_out13_24 ) , .A4( u2_u13_u2_n111 ) , .A3( u2_u13_u2_n112 ) , .A1( u2_u13_u2_n130 ) , .A2( u2_u13_u2_n187 ) );
  AOI221_X1 u2_u13_u2_U89 (.A( u2_u13_u2_n109 ) , .B1( u2_u13_u2_n110 ) , .ZN( u2_u13_u2_n111 ) , .C1( u2_u13_u2_n134 ) , .C2( u2_u13_u2_n170 ) , .B2( u2_u13_u2_n173 ) );
  OAI22_X1 u2_u13_u2_U9 (.ZN( u2_u13_u2_n109 ) , .A2( u2_u13_u2_n113 ) , .B2( u2_u13_u2_n133 ) , .B1( u2_u13_u2_n167 ) , .A1( u2_u13_u2_n168 ) );
  AOI21_X1 u2_u13_u2_U90 (.ZN( u2_u13_u2_n112 ) , .B2( u2_u13_u2_n156 ) , .A( u2_u13_u2_n164 ) , .B1( u2_u13_u2_n181 ) );
  NAND4_X1 u2_u13_u2_U91 (.ZN( u2_out13_16 ) , .A4( u2_u13_u2_n128 ) , .A3( u2_u13_u2_n129 ) , .A1( u2_u13_u2_n130 ) , .A2( u2_u13_u2_n186 ) );
  AOI22_X1 u2_u13_u2_U92 (.A2( u2_u13_u2_n118 ) , .ZN( u2_u13_u2_n129 ) , .A1( u2_u13_u2_n140 ) , .B1( u2_u13_u2_n157 ) , .B2( u2_u13_u2_n170 ) );
  INV_X1 u2_u13_u2_U93 (.A( u2_u13_u2_n163 ) , .ZN( u2_u13_u2_n186 ) );
  OR4_X1 u2_u13_u2_U94 (.ZN( u2_out13_6 ) , .A4( u2_u13_u2_n161 ) , .A3( u2_u13_u2_n162 ) , .A2( u2_u13_u2_n163 ) , .A1( u2_u13_u2_n164 ) );
  OR3_X1 u2_u13_u2_U95 (.A2( u2_u13_u2_n159 ) , .A1( u2_u13_u2_n160 ) , .ZN( u2_u13_u2_n161 ) , .A3( u2_u13_u2_n183 ) );
  AOI21_X1 u2_u13_u2_U96 (.B2( u2_u13_u2_n154 ) , .B1( u2_u13_u2_n155 ) , .ZN( u2_u13_u2_n159 ) , .A( u2_u13_u2_n167 ) );
  NAND3_X1 u2_u13_u2_U97 (.A2( u2_u13_u2_n117 ) , .A1( u2_u13_u2_n122 ) , .A3( u2_u13_u2_n123 ) , .ZN( u2_u13_u2_n134 ) );
  NAND3_X1 u2_u13_u2_U98 (.ZN( u2_u13_u2_n110 ) , .A2( u2_u13_u2_n131 ) , .A3( u2_u13_u2_n139 ) , .A1( u2_u13_u2_n154 ) );
  NAND3_X1 u2_u13_u2_U99 (.A2( u2_u13_u2_n100 ) , .ZN( u2_u13_u2_n101 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n114 ) );
  INV_X1 u2_u13_u5_U10 (.A( u2_u13_u5_n121 ) , .ZN( u2_u13_u5_n177 ) );
  NOR3_X1 u2_u13_u5_U100 (.A3( u2_u13_u5_n141 ) , .A1( u2_u13_u5_n142 ) , .ZN( u2_u13_u5_n143 ) , .A2( u2_u13_u5_n191 ) );
  NAND4_X1 u2_u13_u5_U101 (.ZN( u2_out13_4 ) , .A4( u2_u13_u5_n112 ) , .A2( u2_u13_u5_n113 ) , .A1( u2_u13_u5_n114 ) , .A3( u2_u13_u5_n195 ) );
  AOI211_X1 u2_u13_u5_U102 (.A( u2_u13_u5_n110 ) , .C1( u2_u13_u5_n111 ) , .ZN( u2_u13_u5_n112 ) , .B( u2_u13_u5_n118 ) , .C2( u2_u13_u5_n177 ) );
  AOI222_X1 u2_u13_u5_U103 (.ZN( u2_u13_u5_n113 ) , .A1( u2_u13_u5_n131 ) , .C1( u2_u13_u5_n148 ) , .B2( u2_u13_u5_n174 ) , .C2( u2_u13_u5_n178 ) , .A2( u2_u13_u5_n179 ) , .B1( u2_u13_u5_n99 ) );
  NAND3_X1 u2_u13_u5_U104 (.A2( u2_u13_u5_n154 ) , .A3( u2_u13_u5_n158 ) , .A1( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n99 ) );
  NOR2_X1 u2_u13_u5_U11 (.ZN( u2_u13_u5_n160 ) , .A2( u2_u13_u5_n173 ) , .A1( u2_u13_u5_n177 ) );
  INV_X1 u2_u13_u5_U12 (.A( u2_u13_u5_n150 ) , .ZN( u2_u13_u5_n174 ) );
  AOI21_X1 u2_u13_u5_U13 (.A( u2_u13_u5_n160 ) , .B2( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n162 ) , .B1( u2_u13_u5_n192 ) );
  INV_X1 u2_u13_u5_U14 (.A( u2_u13_u5_n159 ) , .ZN( u2_u13_u5_n192 ) );
  AOI21_X1 u2_u13_u5_U15 (.A( u2_u13_u5_n156 ) , .B2( u2_u13_u5_n157 ) , .B1( u2_u13_u5_n158 ) , .ZN( u2_u13_u5_n163 ) );
  AOI21_X1 u2_u13_u5_U16 (.B2( u2_u13_u5_n139 ) , .B1( u2_u13_u5_n140 ) , .ZN( u2_u13_u5_n141 ) , .A( u2_u13_u5_n150 ) );
  OAI21_X1 u2_u13_u5_U17 (.A( u2_u13_u5_n133 ) , .B2( u2_u13_u5_n134 ) , .B1( u2_u13_u5_n135 ) , .ZN( u2_u13_u5_n142 ) );
  OAI21_X1 u2_u13_u5_U18 (.ZN( u2_u13_u5_n133 ) , .B2( u2_u13_u5_n147 ) , .A( u2_u13_u5_n173 ) , .B1( u2_u13_u5_n188 ) );
  NAND2_X1 u2_u13_u5_U19 (.A2( u2_u13_u5_n119 ) , .A1( u2_u13_u5_n123 ) , .ZN( u2_u13_u5_n137 ) );
  INV_X1 u2_u13_u5_U20 (.A( u2_u13_u5_n155 ) , .ZN( u2_u13_u5_n194 ) );
  NAND2_X1 u2_u13_u5_U21 (.A1( u2_u13_u5_n121 ) , .ZN( u2_u13_u5_n132 ) , .A2( u2_u13_u5_n172 ) );
  NAND2_X1 u2_u13_u5_U22 (.A2( u2_u13_u5_n122 ) , .ZN( u2_u13_u5_n136 ) , .A1( u2_u13_u5_n154 ) );
  NAND2_X1 u2_u13_u5_U23 (.A2( u2_u13_u5_n119 ) , .A1( u2_u13_u5_n120 ) , .ZN( u2_u13_u5_n159 ) );
  INV_X1 u2_u13_u5_U24 (.A( u2_u13_u5_n156 ) , .ZN( u2_u13_u5_n175 ) );
  INV_X1 u2_u13_u5_U25 (.A( u2_u13_u5_n158 ) , .ZN( u2_u13_u5_n188 ) );
  INV_X1 u2_u13_u5_U26 (.A( u2_u13_u5_n152 ) , .ZN( u2_u13_u5_n179 ) );
  INV_X1 u2_u13_u5_U27 (.A( u2_u13_u5_n140 ) , .ZN( u2_u13_u5_n182 ) );
  INV_X1 u2_u13_u5_U28 (.A( u2_u13_u5_n151 ) , .ZN( u2_u13_u5_n183 ) );
  INV_X1 u2_u13_u5_U29 (.A( u2_u13_u5_n123 ) , .ZN( u2_u13_u5_n185 ) );
  NOR2_X1 u2_u13_u5_U3 (.ZN( u2_u13_u5_n134 ) , .A1( u2_u13_u5_n183 ) , .A2( u2_u13_u5_n190 ) );
  INV_X1 u2_u13_u5_U30 (.A( u2_u13_u5_n161 ) , .ZN( u2_u13_u5_n184 ) );
  INV_X1 u2_u13_u5_U31 (.A( u2_u13_u5_n139 ) , .ZN( u2_u13_u5_n189 ) );
  INV_X1 u2_u13_u5_U32 (.A( u2_u13_u5_n157 ) , .ZN( u2_u13_u5_n190 ) );
  INV_X1 u2_u13_u5_U33 (.A( u2_u13_u5_n120 ) , .ZN( u2_u13_u5_n193 ) );
  NAND2_X1 u2_u13_u5_U34 (.ZN( u2_u13_u5_n111 ) , .A1( u2_u13_u5_n140 ) , .A2( u2_u13_u5_n155 ) );
  NOR2_X1 u2_u13_u5_U35 (.ZN( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n170 ) , .A2( u2_u13_u5_n180 ) );
  INV_X1 u2_u13_u5_U36 (.A( u2_u13_u5_n117 ) , .ZN( u2_u13_u5_n196 ) );
  OAI221_X1 u2_u13_u5_U37 (.A( u2_u13_u5_n116 ) , .ZN( u2_u13_u5_n117 ) , .B2( u2_u13_u5_n119 ) , .C1( u2_u13_u5_n153 ) , .C2( u2_u13_u5_n158 ) , .B1( u2_u13_u5_n172 ) );
  AOI222_X1 u2_u13_u5_U38 (.ZN( u2_u13_u5_n116 ) , .B2( u2_u13_u5_n145 ) , .C1( u2_u13_u5_n148 ) , .A2( u2_u13_u5_n174 ) , .C2( u2_u13_u5_n177 ) , .B1( u2_u13_u5_n187 ) , .A1( u2_u13_u5_n193 ) );
  INV_X1 u2_u13_u5_U39 (.A( u2_u13_u5_n115 ) , .ZN( u2_u13_u5_n187 ) );
  INV_X1 u2_u13_u5_U4 (.A( u2_u13_u5_n138 ) , .ZN( u2_u13_u5_n191 ) );
  AOI22_X1 u2_u13_u5_U40 (.B2( u2_u13_u5_n131 ) , .A2( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n169 ) , .B1( u2_u13_u5_n174 ) , .A1( u2_u13_u5_n185 ) );
  NOR2_X1 u2_u13_u5_U41 (.A1( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n150 ) , .A2( u2_u13_u5_n173 ) );
  AOI21_X1 u2_u13_u5_U42 (.A( u2_u13_u5_n118 ) , .B2( u2_u13_u5_n145 ) , .ZN( u2_u13_u5_n168 ) , .B1( u2_u13_u5_n186 ) );
  INV_X1 u2_u13_u5_U43 (.A( u2_u13_u5_n122 ) , .ZN( u2_u13_u5_n186 ) );
  NOR2_X1 u2_u13_u5_U44 (.A1( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n152 ) , .A2( u2_u13_u5_n176 ) );
  NOR2_X1 u2_u13_u5_U45 (.A1( u2_u13_u5_n115 ) , .ZN( u2_u13_u5_n118 ) , .A2( u2_u13_u5_n153 ) );
  NOR2_X1 u2_u13_u5_U46 (.A2( u2_u13_u5_n145 ) , .ZN( u2_u13_u5_n156 ) , .A1( u2_u13_u5_n174 ) );
  NOR2_X1 u2_u13_u5_U47 (.ZN( u2_u13_u5_n121 ) , .A2( u2_u13_u5_n145 ) , .A1( u2_u13_u5_n176 ) );
  AOI22_X1 u2_u13_u5_U48 (.ZN( u2_u13_u5_n114 ) , .A2( u2_u13_u5_n137 ) , .A1( u2_u13_u5_n145 ) , .B2( u2_u13_u5_n175 ) , .B1( u2_u13_u5_n193 ) );
  OAI211_X1 u2_u13_u5_U49 (.B( u2_u13_u5_n124 ) , .A( u2_u13_u5_n125 ) , .C2( u2_u13_u5_n126 ) , .C1( u2_u13_u5_n127 ) , .ZN( u2_u13_u5_n128 ) );
  OAI21_X1 u2_u13_u5_U5 (.B2( u2_u13_u5_n136 ) , .B1( u2_u13_u5_n137 ) , .ZN( u2_u13_u5_n138 ) , .A( u2_u13_u5_n177 ) );
  NOR3_X1 u2_u13_u5_U50 (.ZN( u2_u13_u5_n127 ) , .A1( u2_u13_u5_n136 ) , .A3( u2_u13_u5_n148 ) , .A2( u2_u13_u5_n182 ) );
  OAI21_X1 u2_u13_u5_U51 (.ZN( u2_u13_u5_n124 ) , .A( u2_u13_u5_n177 ) , .B2( u2_u13_u5_n183 ) , .B1( u2_u13_u5_n189 ) );
  OAI21_X1 u2_u13_u5_U52 (.ZN( u2_u13_u5_n125 ) , .A( u2_u13_u5_n174 ) , .B2( u2_u13_u5_n185 ) , .B1( u2_u13_u5_n190 ) );
  AOI21_X1 u2_u13_u5_U53 (.A( u2_u13_u5_n153 ) , .B2( u2_u13_u5_n154 ) , .B1( u2_u13_u5_n155 ) , .ZN( u2_u13_u5_n164 ) );
  AOI21_X1 u2_u13_u5_U54 (.ZN( u2_u13_u5_n110 ) , .B1( u2_u13_u5_n122 ) , .B2( u2_u13_u5_n139 ) , .A( u2_u13_u5_n153 ) );
  INV_X1 u2_u13_u5_U55 (.A( u2_u13_u5_n153 ) , .ZN( u2_u13_u5_n176 ) );
  INV_X1 u2_u13_u5_U56 (.A( u2_u13_u5_n126 ) , .ZN( u2_u13_u5_n173 ) );
  AND2_X1 u2_u13_u5_U57 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n147 ) );
  AND2_X1 u2_u13_u5_U58 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n148 ) );
  NAND2_X1 u2_u13_u5_U59 (.A1( u2_u13_u5_n105 ) , .A2( u2_u13_u5_n106 ) , .ZN( u2_u13_u5_n158 ) );
  INV_X1 u2_u13_u5_U6 (.A( u2_u13_u5_n135 ) , .ZN( u2_u13_u5_n178 ) );
  NAND2_X1 u2_u13_u5_U60 (.A2( u2_u13_u5_n108 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n139 ) );
  NAND2_X1 u2_u13_u5_U61 (.A1( u2_u13_u5_n106 ) , .A2( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n119 ) );
  NAND2_X1 u2_u13_u5_U62 (.A2( u2_u13_u5_n103 ) , .A1( u2_u13_u5_n105 ) , .ZN( u2_u13_u5_n140 ) );
  NAND2_X1 u2_u13_u5_U63 (.A2( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n105 ) , .ZN( u2_u13_u5_n155 ) );
  NAND2_X1 u2_u13_u5_U64 (.A2( u2_u13_u5_n106 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n122 ) );
  NAND2_X1 u2_u13_u5_U65 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n106 ) , .ZN( u2_u13_u5_n115 ) );
  NAND2_X1 u2_u13_u5_U66 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n103 ) , .ZN( u2_u13_u5_n161 ) );
  NAND2_X1 u2_u13_u5_U67 (.A1( u2_u13_u5_n105 ) , .A2( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n154 ) );
  INV_X1 u2_u13_u5_U68 (.A( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n172 ) );
  NAND2_X1 u2_u13_u5_U69 (.A1( u2_u13_u5_n103 ) , .A2( u2_u13_u5_n108 ) , .ZN( u2_u13_u5_n123 ) );
  OAI22_X1 u2_u13_u5_U7 (.B2( u2_u13_u5_n149 ) , .B1( u2_u13_u5_n150 ) , .A2( u2_u13_u5_n151 ) , .A1( u2_u13_u5_n152 ) , .ZN( u2_u13_u5_n165 ) );
  NAND2_X1 u2_u13_u5_U70 (.A2( u2_u13_u5_n103 ) , .A1( u2_u13_u5_n107 ) , .ZN( u2_u13_u5_n151 ) );
  NAND2_X1 u2_u13_u5_U71 (.A2( u2_u13_u5_n107 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n120 ) );
  NAND2_X1 u2_u13_u5_U72 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n109 ) , .ZN( u2_u13_u5_n157 ) );
  AND2_X1 u2_u13_u5_U73 (.A2( u2_u13_u5_n100 ) , .A1( u2_u13_u5_n104 ) , .ZN( u2_u13_u5_n131 ) );
  INV_X1 u2_u13_u5_U74 (.A( u2_u13_u5_n102 ) , .ZN( u2_u13_u5_n195 ) );
  OAI221_X1 u2_u13_u5_U75 (.A( u2_u13_u5_n101 ) , .ZN( u2_u13_u5_n102 ) , .C2( u2_u13_u5_n115 ) , .C1( u2_u13_u5_n126 ) , .B1( u2_u13_u5_n134 ) , .B2( u2_u13_u5_n160 ) );
  OAI21_X1 u2_u13_u5_U76 (.ZN( u2_u13_u5_n101 ) , .B1( u2_u13_u5_n137 ) , .A( u2_u13_u5_n146 ) , .B2( u2_u13_u5_n147 ) );
  NOR2_X1 u2_u13_u5_U77 (.A2( u2_u13_X_34 ) , .A1( u2_u13_X_35 ) , .ZN( u2_u13_u5_n145 ) );
  NOR2_X1 u2_u13_u5_U78 (.A2( u2_u13_X_34 ) , .ZN( u2_u13_u5_n146 ) , .A1( u2_u13_u5_n171 ) );
  NOR2_X1 u2_u13_u5_U79 (.A2( u2_u13_X_31 ) , .A1( u2_u13_X_32 ) , .ZN( u2_u13_u5_n103 ) );
  NOR3_X1 u2_u13_u5_U8 (.A2( u2_u13_u5_n147 ) , .A1( u2_u13_u5_n148 ) , .ZN( u2_u13_u5_n149 ) , .A3( u2_u13_u5_n194 ) );
  NOR2_X1 u2_u13_u5_U80 (.A2( u2_u13_X_36 ) , .ZN( u2_u13_u5_n105 ) , .A1( u2_u13_u5_n180 ) );
  NOR2_X1 u2_u13_u5_U81 (.A2( u2_u13_X_33 ) , .ZN( u2_u13_u5_n108 ) , .A1( u2_u13_u5_n170 ) );
  NOR2_X1 u2_u13_u5_U82 (.A2( u2_u13_X_33 ) , .A1( u2_u13_X_36 ) , .ZN( u2_u13_u5_n107 ) );
  NOR2_X1 u2_u13_u5_U83 (.A2( u2_u13_X_31 ) , .ZN( u2_u13_u5_n104 ) , .A1( u2_u13_u5_n181 ) );
  NAND2_X1 u2_u13_u5_U84 (.A2( u2_u13_X_34 ) , .A1( u2_u13_X_35 ) , .ZN( u2_u13_u5_n153 ) );
  NAND2_X1 u2_u13_u5_U85 (.A1( u2_u13_X_34 ) , .ZN( u2_u13_u5_n126 ) , .A2( u2_u13_u5_n171 ) );
  AND2_X1 u2_u13_u5_U86 (.A1( u2_u13_X_31 ) , .A2( u2_u13_X_32 ) , .ZN( u2_u13_u5_n106 ) );
  AND2_X1 u2_u13_u5_U87 (.A1( u2_u13_X_31 ) , .ZN( u2_u13_u5_n109 ) , .A2( u2_u13_u5_n181 ) );
  INV_X1 u2_u13_u5_U88 (.A( u2_u13_X_33 ) , .ZN( u2_u13_u5_n180 ) );
  INV_X1 u2_u13_u5_U89 (.A( u2_u13_X_35 ) , .ZN( u2_u13_u5_n171 ) );
  NOR2_X1 u2_u13_u5_U9 (.ZN( u2_u13_u5_n135 ) , .A1( u2_u13_u5_n173 ) , .A2( u2_u13_u5_n176 ) );
  INV_X1 u2_u13_u5_U90 (.A( u2_u13_X_36 ) , .ZN( u2_u13_u5_n170 ) );
  INV_X1 u2_u13_u5_U91 (.A( u2_u13_X_32 ) , .ZN( u2_u13_u5_n181 ) );
  NAND4_X1 u2_u13_u5_U92 (.ZN( u2_out13_29 ) , .A4( u2_u13_u5_n129 ) , .A3( u2_u13_u5_n130 ) , .A2( u2_u13_u5_n168 ) , .A1( u2_u13_u5_n196 ) );
  AOI221_X1 u2_u13_u5_U93 (.A( u2_u13_u5_n128 ) , .ZN( u2_u13_u5_n129 ) , .C2( u2_u13_u5_n132 ) , .B2( u2_u13_u5_n159 ) , .B1( u2_u13_u5_n176 ) , .C1( u2_u13_u5_n184 ) );
  AOI222_X1 u2_u13_u5_U94 (.ZN( u2_u13_u5_n130 ) , .A2( u2_u13_u5_n146 ) , .B1( u2_u13_u5_n147 ) , .C2( u2_u13_u5_n175 ) , .B2( u2_u13_u5_n179 ) , .A1( u2_u13_u5_n188 ) , .C1( u2_u13_u5_n194 ) );
  NAND4_X1 u2_u13_u5_U95 (.ZN( u2_out13_19 ) , .A4( u2_u13_u5_n166 ) , .A3( u2_u13_u5_n167 ) , .A2( u2_u13_u5_n168 ) , .A1( u2_u13_u5_n169 ) );
  AOI22_X1 u2_u13_u5_U96 (.B2( u2_u13_u5_n145 ) , .A2( u2_u13_u5_n146 ) , .ZN( u2_u13_u5_n167 ) , .B1( u2_u13_u5_n182 ) , .A1( u2_u13_u5_n189 ) );
  NOR4_X1 u2_u13_u5_U97 (.A4( u2_u13_u5_n162 ) , .A3( u2_u13_u5_n163 ) , .A2( u2_u13_u5_n164 ) , .A1( u2_u13_u5_n165 ) , .ZN( u2_u13_u5_n166 ) );
  NAND4_X1 u2_u13_u5_U98 (.ZN( u2_out13_11 ) , .A4( u2_u13_u5_n143 ) , .A3( u2_u13_u5_n144 ) , .A2( u2_u13_u5_n169 ) , .A1( u2_u13_u5_n196 ) );
  AOI22_X1 u2_u13_u5_U99 (.A2( u2_u13_u5_n132 ) , .ZN( u2_u13_u5_n144 ) , .B2( u2_u13_u5_n145 ) , .B1( u2_u13_u5_n184 ) , .A1( u2_u13_u5_n194 ) );
  AOI22_X1 u2_u13_u6_U10 (.A2( u2_u13_u6_n151 ) , .B2( u2_u13_u6_n161 ) , .A1( u2_u13_u6_n167 ) , .B1( u2_u13_u6_n170 ) , .ZN( u2_u13_u6_n89 ) );
  AOI21_X1 u2_u13_u6_U11 (.B1( u2_u13_u6_n107 ) , .B2( u2_u13_u6_n132 ) , .A( u2_u13_u6_n158 ) , .ZN( u2_u13_u6_n88 ) );
  AOI21_X1 u2_u13_u6_U12 (.B2( u2_u13_u6_n147 ) , .B1( u2_u13_u6_n148 ) , .ZN( u2_u13_u6_n149 ) , .A( u2_u13_u6_n158 ) );
  AOI21_X1 u2_u13_u6_U13 (.ZN( u2_u13_u6_n106 ) , .A( u2_u13_u6_n142 ) , .B2( u2_u13_u6_n159 ) , .B1( u2_u13_u6_n164 ) );
  INV_X1 u2_u13_u6_U14 (.A( u2_u13_u6_n155 ) , .ZN( u2_u13_u6_n161 ) );
  INV_X1 u2_u13_u6_U15 (.A( u2_u13_u6_n128 ) , .ZN( u2_u13_u6_n164 ) );
  NAND2_X1 u2_u13_u6_U16 (.ZN( u2_u13_u6_n110 ) , .A1( u2_u13_u6_n122 ) , .A2( u2_u13_u6_n129 ) );
  NAND2_X1 u2_u13_u6_U17 (.ZN( u2_u13_u6_n124 ) , .A2( u2_u13_u6_n146 ) , .A1( u2_u13_u6_n148 ) );
  INV_X1 u2_u13_u6_U18 (.A( u2_u13_u6_n132 ) , .ZN( u2_u13_u6_n171 ) );
  AND2_X1 u2_u13_u6_U19 (.A1( u2_u13_u6_n100 ) , .ZN( u2_u13_u6_n130 ) , .A2( u2_u13_u6_n147 ) );
  INV_X1 u2_u13_u6_U20 (.A( u2_u13_u6_n127 ) , .ZN( u2_u13_u6_n173 ) );
  INV_X1 u2_u13_u6_U21 (.A( u2_u13_u6_n121 ) , .ZN( u2_u13_u6_n167 ) );
  INV_X1 u2_u13_u6_U22 (.A( u2_u13_u6_n100 ) , .ZN( u2_u13_u6_n169 ) );
  INV_X1 u2_u13_u6_U23 (.A( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n170 ) );
  INV_X1 u2_u13_u6_U24 (.A( u2_u13_u6_n113 ) , .ZN( u2_u13_u6_n168 ) );
  AND2_X1 u2_u13_u6_U25 (.A1( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n119 ) , .ZN( u2_u13_u6_n133 ) );
  AND2_X1 u2_u13_u6_U26 (.A2( u2_u13_u6_n121 ) , .A1( u2_u13_u6_n122 ) , .ZN( u2_u13_u6_n131 ) );
  AND3_X1 u2_u13_u6_U27 (.ZN( u2_u13_u6_n120 ) , .A2( u2_u13_u6_n127 ) , .A1( u2_u13_u6_n132 ) , .A3( u2_u13_u6_n145 ) );
  INV_X1 u2_u13_u6_U28 (.A( u2_u13_u6_n146 ) , .ZN( u2_u13_u6_n163 ) );
  AOI222_X1 u2_u13_u6_U29 (.ZN( u2_u13_u6_n114 ) , .A1( u2_u13_u6_n118 ) , .A2( u2_u13_u6_n126 ) , .B2( u2_u13_u6_n151 ) , .C2( u2_u13_u6_n159 ) , .C1( u2_u13_u6_n168 ) , .B1( u2_u13_u6_n169 ) );
  INV_X1 u2_u13_u6_U3 (.A( u2_u13_u6_n110 ) , .ZN( u2_u13_u6_n166 ) );
  NOR2_X1 u2_u13_u6_U30 (.A1( u2_u13_u6_n162 ) , .A2( u2_u13_u6_n165 ) , .ZN( u2_u13_u6_n98 ) );
  AOI211_X1 u2_u13_u6_U31 (.B( u2_u13_u6_n134 ) , .A( u2_u13_u6_n135 ) , .C1( u2_u13_u6_n136 ) , .ZN( u2_u13_u6_n137 ) , .C2( u2_u13_u6_n151 ) );
  AOI21_X1 u2_u13_u6_U32 (.B2( u2_u13_u6_n132 ) , .B1( u2_u13_u6_n133 ) , .ZN( u2_u13_u6_n134 ) , .A( u2_u13_u6_n158 ) );
  AOI21_X1 u2_u13_u6_U33 (.B1( u2_u13_u6_n131 ) , .ZN( u2_u13_u6_n135 ) , .A( u2_u13_u6_n144 ) , .B2( u2_u13_u6_n146 ) );
  NAND4_X1 u2_u13_u6_U34 (.A4( u2_u13_u6_n127 ) , .A3( u2_u13_u6_n128 ) , .A2( u2_u13_u6_n129 ) , .A1( u2_u13_u6_n130 ) , .ZN( u2_u13_u6_n136 ) );
  NAND2_X1 u2_u13_u6_U35 (.A1( u2_u13_u6_n144 ) , .ZN( u2_u13_u6_n151 ) , .A2( u2_u13_u6_n158 ) );
  NAND2_X1 u2_u13_u6_U36 (.ZN( u2_u13_u6_n132 ) , .A1( u2_u13_u6_n91 ) , .A2( u2_u13_u6_n97 ) );
  AOI22_X1 u2_u13_u6_U37 (.B2( u2_u13_u6_n110 ) , .B1( u2_u13_u6_n111 ) , .A1( u2_u13_u6_n112 ) , .ZN( u2_u13_u6_n115 ) , .A2( u2_u13_u6_n161 ) );
  NAND4_X1 u2_u13_u6_U38 (.A3( u2_u13_u6_n109 ) , .ZN( u2_u13_u6_n112 ) , .A4( u2_u13_u6_n132 ) , .A2( u2_u13_u6_n147 ) , .A1( u2_u13_u6_n166 ) );
  NOR2_X1 u2_u13_u6_U39 (.ZN( u2_u13_u6_n109 ) , .A1( u2_u13_u6_n170 ) , .A2( u2_u13_u6_n173 ) );
  INV_X1 u2_u13_u6_U4 (.A( u2_u13_u6_n142 ) , .ZN( u2_u13_u6_n174 ) );
  NOR2_X1 u2_u13_u6_U40 (.A2( u2_u13_u6_n126 ) , .ZN( u2_u13_u6_n155 ) , .A1( u2_u13_u6_n160 ) );
  NAND2_X1 u2_u13_u6_U41 (.ZN( u2_u13_u6_n146 ) , .A2( u2_u13_u6_n94 ) , .A1( u2_u13_u6_n99 ) );
  AOI21_X1 u2_u13_u6_U42 (.A( u2_u13_u6_n144 ) , .B2( u2_u13_u6_n145 ) , .B1( u2_u13_u6_n146 ) , .ZN( u2_u13_u6_n150 ) );
  INV_X1 u2_u13_u6_U43 (.A( u2_u13_u6_n111 ) , .ZN( u2_u13_u6_n158 ) );
  NAND2_X1 u2_u13_u6_U44 (.ZN( u2_u13_u6_n127 ) , .A1( u2_u13_u6_n91 ) , .A2( u2_u13_u6_n92 ) );
  NAND2_X1 u2_u13_u6_U45 (.ZN( u2_u13_u6_n129 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n96 ) );
  INV_X1 u2_u13_u6_U46 (.A( u2_u13_u6_n144 ) , .ZN( u2_u13_u6_n159 ) );
  NAND2_X1 u2_u13_u6_U47 (.ZN( u2_u13_u6_n145 ) , .A2( u2_u13_u6_n97 ) , .A1( u2_u13_u6_n98 ) );
  NAND2_X1 u2_u13_u6_U48 (.ZN( u2_u13_u6_n148 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n94 ) );
  NAND2_X1 u2_u13_u6_U49 (.ZN( u2_u13_u6_n108 ) , .A2( u2_u13_u6_n139 ) , .A1( u2_u13_u6_n144 ) );
  NAND2_X1 u2_u13_u6_U5 (.A2( u2_u13_u6_n143 ) , .ZN( u2_u13_u6_n152 ) , .A1( u2_u13_u6_n166 ) );
  NAND2_X1 u2_u13_u6_U50 (.ZN( u2_u13_u6_n121 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n97 ) );
  NAND2_X1 u2_u13_u6_U51 (.ZN( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n95 ) );
  AND2_X1 u2_u13_u6_U52 (.ZN( u2_u13_u6_n118 ) , .A2( u2_u13_u6_n91 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U53 (.ZN( u2_u13_u6_n147 ) , .A2( u2_u13_u6_n98 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U54 (.ZN( u2_u13_u6_n128 ) , .A1( u2_u13_u6_n94 ) , .A2( u2_u13_u6_n96 ) );
  NAND2_X1 u2_u13_u6_U55 (.ZN( u2_u13_u6_n119 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U56 (.ZN( u2_u13_u6_n123 ) , .A2( u2_u13_u6_n91 ) , .A1( u2_u13_u6_n96 ) );
  NAND2_X1 u2_u13_u6_U57 (.ZN( u2_u13_u6_n100 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n98 ) );
  NAND2_X1 u2_u13_u6_U58 (.ZN( u2_u13_u6_n122 ) , .A1( u2_u13_u6_n94 ) , .A2( u2_u13_u6_n97 ) );
  INV_X1 u2_u13_u6_U59 (.A( u2_u13_u6_n139 ) , .ZN( u2_u13_u6_n160 ) );
  AOI22_X1 u2_u13_u6_U6 (.B2( u2_u13_u6_n101 ) , .A1( u2_u13_u6_n102 ) , .ZN( u2_u13_u6_n103 ) , .B1( u2_u13_u6_n160 ) , .A2( u2_u13_u6_n161 ) );
  NAND2_X1 u2_u13_u6_U60 (.ZN( u2_u13_u6_n113 ) , .A1( u2_u13_u6_n96 ) , .A2( u2_u13_u6_n98 ) );
  NOR2_X1 u2_u13_u6_U61 (.A2( u2_u13_X_40 ) , .A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n126 ) );
  NOR2_X1 u2_u13_u6_U62 (.A2( u2_u13_X_39 ) , .A1( u2_u13_X_42 ) , .ZN( u2_u13_u6_n92 ) );
  NOR2_X1 u2_u13_u6_U63 (.A2( u2_u13_X_39 ) , .A1( u2_u13_u6_n156 ) , .ZN( u2_u13_u6_n97 ) );
  NOR2_X1 u2_u13_u6_U64 (.A2( u2_u13_X_38 ) , .A1( u2_u13_u6_n165 ) , .ZN( u2_u13_u6_n95 ) );
  NOR2_X1 u2_u13_u6_U65 (.A2( u2_u13_X_41 ) , .ZN( u2_u13_u6_n111 ) , .A1( u2_u13_u6_n157 ) );
  NOR2_X1 u2_u13_u6_U66 (.A2( u2_u13_X_37 ) , .A1( u2_u13_u6_n162 ) , .ZN( u2_u13_u6_n94 ) );
  NOR2_X1 u2_u13_u6_U67 (.A2( u2_u13_X_37 ) , .A1( u2_u13_X_38 ) , .ZN( u2_u13_u6_n91 ) );
  NAND2_X1 u2_u13_u6_U68 (.A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n144 ) , .A2( u2_u13_u6_n157 ) );
  NAND2_X1 u2_u13_u6_U69 (.A2( u2_u13_X_40 ) , .A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n139 ) );
  NOR2_X1 u2_u13_u6_U7 (.A1( u2_u13_u6_n118 ) , .ZN( u2_u13_u6_n143 ) , .A2( u2_u13_u6_n168 ) );
  AND2_X1 u2_u13_u6_U70 (.A1( u2_u13_X_39 ) , .A2( u2_u13_u6_n156 ) , .ZN( u2_u13_u6_n96 ) );
  AND2_X1 u2_u13_u6_U71 (.A1( u2_u13_X_39 ) , .A2( u2_u13_X_42 ) , .ZN( u2_u13_u6_n99 ) );
  INV_X1 u2_u13_u6_U72 (.A( u2_u13_X_40 ) , .ZN( u2_u13_u6_n157 ) );
  INV_X1 u2_u13_u6_U73 (.A( u2_u13_X_37 ) , .ZN( u2_u13_u6_n165 ) );
  INV_X1 u2_u13_u6_U74 (.A( u2_u13_X_38 ) , .ZN( u2_u13_u6_n162 ) );
  INV_X1 u2_u13_u6_U75 (.A( u2_u13_X_42 ) , .ZN( u2_u13_u6_n156 ) );
  NAND4_X1 u2_u13_u6_U76 (.ZN( u2_out13_32 ) , .A4( u2_u13_u6_n103 ) , .A3( u2_u13_u6_n104 ) , .A2( u2_u13_u6_n105 ) , .A1( u2_u13_u6_n106 ) );
  AOI22_X1 u2_u13_u6_U77 (.ZN( u2_u13_u6_n105 ) , .A2( u2_u13_u6_n108 ) , .A1( u2_u13_u6_n118 ) , .B2( u2_u13_u6_n126 ) , .B1( u2_u13_u6_n171 ) );
  AOI22_X1 u2_u13_u6_U78 (.ZN( u2_u13_u6_n104 ) , .A1( u2_u13_u6_n111 ) , .B1( u2_u13_u6_n124 ) , .B2( u2_u13_u6_n151 ) , .A2( u2_u13_u6_n93 ) );
  NAND4_X1 u2_u13_u6_U79 (.ZN( u2_out13_12 ) , .A4( u2_u13_u6_n114 ) , .A3( u2_u13_u6_n115 ) , .A2( u2_u13_u6_n116 ) , .A1( u2_u13_u6_n117 ) );
  OAI21_X1 u2_u13_u6_U8 (.A( u2_u13_u6_n159 ) , .B1( u2_u13_u6_n169 ) , .B2( u2_u13_u6_n173 ) , .ZN( u2_u13_u6_n90 ) );
  OAI22_X1 u2_u13_u6_U80 (.B2( u2_u13_u6_n111 ) , .ZN( u2_u13_u6_n116 ) , .B1( u2_u13_u6_n126 ) , .A2( u2_u13_u6_n164 ) , .A1( u2_u13_u6_n167 ) );
  OAI21_X1 u2_u13_u6_U81 (.A( u2_u13_u6_n108 ) , .ZN( u2_u13_u6_n117 ) , .B2( u2_u13_u6_n141 ) , .B1( u2_u13_u6_n163 ) );
  OAI211_X1 u2_u13_u6_U82 (.ZN( u2_out13_7 ) , .B( u2_u13_u6_n153 ) , .C2( u2_u13_u6_n154 ) , .C1( u2_u13_u6_n155 ) , .A( u2_u13_u6_n174 ) );
  NOR3_X1 u2_u13_u6_U83 (.A1( u2_u13_u6_n141 ) , .ZN( u2_u13_u6_n154 ) , .A3( u2_u13_u6_n164 ) , .A2( u2_u13_u6_n171 ) );
  AOI211_X1 u2_u13_u6_U84 (.B( u2_u13_u6_n149 ) , .A( u2_u13_u6_n150 ) , .C2( u2_u13_u6_n151 ) , .C1( u2_u13_u6_n152 ) , .ZN( u2_u13_u6_n153 ) );
  OAI211_X1 u2_u13_u6_U85 (.ZN( u2_out13_22 ) , .B( u2_u13_u6_n137 ) , .A( u2_u13_u6_n138 ) , .C2( u2_u13_u6_n139 ) , .C1( u2_u13_u6_n140 ) );
  AOI22_X1 u2_u13_u6_U86 (.B1( u2_u13_u6_n124 ) , .A2( u2_u13_u6_n125 ) , .A1( u2_u13_u6_n126 ) , .ZN( u2_u13_u6_n138 ) , .B2( u2_u13_u6_n161 ) );
  AND4_X1 u2_u13_u6_U87 (.A3( u2_u13_u6_n119 ) , .A1( u2_u13_u6_n120 ) , .A4( u2_u13_u6_n129 ) , .ZN( u2_u13_u6_n140 ) , .A2( u2_u13_u6_n143 ) );
  NAND3_X1 u2_u13_u6_U88 (.A2( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n125 ) , .A1( u2_u13_u6_n130 ) , .A3( u2_u13_u6_n131 ) );
  NAND3_X1 u2_u13_u6_U89 (.A3( u2_u13_u6_n133 ) , .ZN( u2_u13_u6_n141 ) , .A1( u2_u13_u6_n145 ) , .A2( u2_u13_u6_n148 ) );
  INV_X1 u2_u13_u6_U9 (.ZN( u2_u13_u6_n172 ) , .A( u2_u13_u6_n88 ) );
  NAND3_X1 u2_u13_u6_U90 (.ZN( u2_u13_u6_n101 ) , .A3( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n121 ) , .A1( u2_u13_u6_n127 ) );
  NAND3_X1 u2_u13_u6_U91 (.ZN( u2_u13_u6_n102 ) , .A3( u2_u13_u6_n130 ) , .A2( u2_u13_u6_n145 ) , .A1( u2_u13_u6_n166 ) );
  NAND3_X1 u2_u13_u6_U92 (.A3( u2_u13_u6_n113 ) , .A1( u2_u13_u6_n119 ) , .A2( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n93 ) );
  NAND3_X1 u2_u13_u6_U93 (.ZN( u2_u13_u6_n142 ) , .A2( u2_u13_u6_n172 ) , .A3( u2_u13_u6_n89 ) , .A1( u2_u13_u6_n90 ) );
  XOR2_X1 u2_u14_U10 (.B( u2_K15_45 ) , .A( u2_R13_30 ) , .Z( u2_u14_X_45 ) );
  XOR2_X1 u2_u14_U11 (.B( u2_K15_44 ) , .A( u2_R13_29 ) , .Z( u2_u14_X_44 ) );
  XOR2_X1 u2_u14_U12 (.B( u2_K15_43 ) , .A( u2_R13_28 ) , .Z( u2_u14_X_43 ) );
  XOR2_X1 u2_u14_U13 (.B( u2_K15_42 ) , .A( u2_R13_29 ) , .Z( u2_u14_X_42 ) );
  XOR2_X1 u2_u14_U14 (.B( u2_K15_41 ) , .A( u2_R13_28 ) , .Z( u2_u14_X_41 ) );
  XOR2_X1 u2_u14_U15 (.B( u2_K15_40 ) , .A( u2_R13_27 ) , .Z( u2_u14_X_40 ) );
  XOR2_X1 u2_u14_U17 (.B( u2_K15_39 ) , .A( u2_R13_26 ) , .Z( u2_u14_X_39 ) );
  XOR2_X1 u2_u14_U18 (.B( u2_K15_38 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_38 ) );
  XOR2_X1 u2_u14_U19 (.B( u2_K15_37 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_37 ) );
  XOR2_X1 u2_u14_U20 (.B( u2_K15_36 ) , .A( u2_R13_25 ) , .Z( u2_u14_X_36 ) );
  XOR2_X1 u2_u14_U21 (.B( u2_K15_35 ) , .A( u2_R13_24 ) , .Z( u2_u14_X_35 ) );
  XOR2_X1 u2_u14_U22 (.B( u2_K15_34 ) , .A( u2_R13_23 ) , .Z( u2_u14_X_34 ) );
  XOR2_X1 u2_u14_U23 (.B( u2_K15_33 ) , .A( u2_R13_22 ) , .Z( u2_u14_X_33 ) );
  XOR2_X1 u2_u14_U24 (.B( u2_K15_32 ) , .A( u2_R13_21 ) , .Z( u2_u14_X_32 ) );
  XOR2_X1 u2_u14_U25 (.B( u2_K15_31 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_31 ) );
  XOR2_X1 u2_u14_U26 (.B( u2_K15_30 ) , .A( u2_R13_21 ) , .Z( u2_u14_X_30 ) );
  XOR2_X1 u2_u14_U28 (.B( u2_K15_29 ) , .A( u2_R13_20 ) , .Z( u2_u14_X_29 ) );
  XOR2_X1 u2_u14_U29 (.B( u2_K15_28 ) , .A( u2_R13_19 ) , .Z( u2_u14_X_28 ) );
  XOR2_X1 u2_u14_U30 (.B( u2_K15_27 ) , .A( u2_R13_18 ) , .Z( u2_u14_X_27 ) );
  XOR2_X1 u2_u14_U31 (.B( u2_K15_26 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_26 ) );
  XOR2_X1 u2_u14_U32 (.B( u2_K15_25 ) , .A( u2_R13_16 ) , .Z( u2_u14_X_25 ) );
  XOR2_X1 u2_u14_U7 (.B( u2_K15_48 ) , .A( u2_R13_1 ) , .Z( u2_u14_X_48 ) );
  XOR2_X1 u2_u14_U8 (.B( u2_K15_47 ) , .A( u2_R13_32 ) , .Z( u2_u14_X_47 ) );
  XOR2_X1 u2_u14_U9 (.B( u2_K15_46 ) , .A( u2_R13_31 ) , .Z( u2_u14_X_46 ) );
  OAI22_X1 u2_u14_u4_U10 (.B2( u2_u14_u4_n135 ) , .ZN( u2_u14_u4_n137 ) , .B1( u2_u14_u4_n153 ) , .A1( u2_u14_u4_n155 ) , .A2( u2_u14_u4_n171 ) );
  AND3_X1 u2_u14_u4_U11 (.A2( u2_u14_u4_n134 ) , .ZN( u2_u14_u4_n135 ) , .A3( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n157 ) );
  NAND2_X1 u2_u14_u4_U12 (.ZN( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n173 ) );
  AOI21_X1 u2_u14_u4_U13 (.B2( u2_u14_u4_n160 ) , .B1( u2_u14_u4_n161 ) , .ZN( u2_u14_u4_n162 ) , .A( u2_u14_u4_n170 ) );
  AOI21_X1 u2_u14_u4_U14 (.ZN( u2_u14_u4_n107 ) , .B2( u2_u14_u4_n143 ) , .A( u2_u14_u4_n174 ) , .B1( u2_u14_u4_n184 ) );
  AOI21_X1 u2_u14_u4_U15 (.B2( u2_u14_u4_n158 ) , .B1( u2_u14_u4_n159 ) , .ZN( u2_u14_u4_n163 ) , .A( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U16 (.A( u2_u14_u4_n153 ) , .B2( u2_u14_u4_n154 ) , .B1( u2_u14_u4_n155 ) , .ZN( u2_u14_u4_n165 ) );
  AOI21_X1 u2_u14_u4_U17 (.A( u2_u14_u4_n156 ) , .B2( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n164 ) , .B1( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U18 (.A( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n170 ) );
  AND2_X1 u2_u14_u4_U19 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n155 ) , .A1( u2_u14_u4_n160 ) );
  INV_X1 u2_u14_u4_U20 (.A( u2_u14_u4_n156 ) , .ZN( u2_u14_u4_n175 ) );
  NAND2_X1 u2_u14_u4_U21 (.A2( u2_u14_u4_n118 ) , .ZN( u2_u14_u4_n131 ) , .A1( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U22 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n130 ) );
  NAND2_X1 u2_u14_u4_U23 (.ZN( u2_u14_u4_n117 ) , .A2( u2_u14_u4_n118 ) , .A1( u2_u14_u4_n148 ) );
  NAND2_X1 u2_u14_u4_U24 (.ZN( u2_u14_u4_n129 ) , .A1( u2_u14_u4_n134 ) , .A2( u2_u14_u4_n148 ) );
  AND3_X1 u2_u14_u4_U25 (.A1( u2_u14_u4_n119 ) , .A2( u2_u14_u4_n143 ) , .A3( u2_u14_u4_n154 ) , .ZN( u2_u14_u4_n161 ) );
  AND2_X1 u2_u14_u4_U26 (.A1( u2_u14_u4_n145 ) , .A2( u2_u14_u4_n147 ) , .ZN( u2_u14_u4_n159 ) );
  OR3_X1 u2_u14_u4_U27 (.A3( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n115 ) , .A1( u2_u14_u4_n116 ) , .ZN( u2_u14_u4_n136 ) );
  AOI21_X1 u2_u14_u4_U28 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n116 ) , .B2( u2_u14_u4_n173 ) , .B1( u2_u14_u4_n174 ) );
  AOI21_X1 u2_u14_u4_U29 (.ZN( u2_u14_u4_n115 ) , .B2( u2_u14_u4_n145 ) , .B1( u2_u14_u4_n146 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U3 (.ZN( u2_u14_u4_n121 ) , .A1( u2_u14_u4_n181 ) , .A2( u2_u14_u4_n182 ) );
  OAI22_X1 u2_u14_u4_U30 (.ZN( u2_u14_u4_n114 ) , .A2( u2_u14_u4_n121 ) , .B1( u2_u14_u4_n160 ) , .B2( u2_u14_u4_n170 ) , .A1( u2_u14_u4_n171 ) );
  INV_X1 u2_u14_u4_U31 (.A( u2_u14_u4_n158 ) , .ZN( u2_u14_u4_n182 ) );
  INV_X1 u2_u14_u4_U32 (.ZN( u2_u14_u4_n181 ) , .A( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U33 (.A( u2_u14_u4_n144 ) , .ZN( u2_u14_u4_n179 ) );
  INV_X1 u2_u14_u4_U34 (.A( u2_u14_u4_n157 ) , .ZN( u2_u14_u4_n178 ) );
  NAND2_X1 u2_u14_u4_U35 (.A2( u2_u14_u4_n154 ) , .A1( u2_u14_u4_n96 ) , .ZN( u2_u14_u4_n97 ) );
  INV_X1 u2_u14_u4_U36 (.ZN( u2_u14_u4_n186 ) , .A( u2_u14_u4_n95 ) );
  OAI221_X1 u2_u14_u4_U37 (.C1( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n158 ) , .B2( u2_u14_u4_n171 ) , .C2( u2_u14_u4_n173 ) , .A( u2_u14_u4_n94 ) , .ZN( u2_u14_u4_n95 ) );
  AOI222_X1 u2_u14_u4_U38 (.B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n138 ) , .C2( u2_u14_u4_n175 ) , .A2( u2_u14_u4_n179 ) , .C1( u2_u14_u4_n181 ) , .B1( u2_u14_u4_n185 ) , .ZN( u2_u14_u4_n94 ) );
  INV_X1 u2_u14_u4_U39 (.A( u2_u14_u4_n113 ) , .ZN( u2_u14_u4_n185 ) );
  INV_X1 u2_u14_u4_U4 (.A( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n184 ) );
  INV_X1 u2_u14_u4_U40 (.A( u2_u14_u4_n143 ) , .ZN( u2_u14_u4_n183 ) );
  NOR2_X1 u2_u14_u4_U41 (.ZN( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n168 ) , .A2( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U42 (.A1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n153 ) );
  NOR2_X1 u2_u14_u4_U43 (.A2( u2_u14_u4_n128 ) , .A1( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n156 ) );
  AOI22_X1 u2_u14_u4_U44 (.B2( u2_u14_u4_n122 ) , .A1( u2_u14_u4_n123 ) , .ZN( u2_u14_u4_n124 ) , .B1( u2_u14_u4_n128 ) , .A2( u2_u14_u4_n172 ) );
  INV_X1 u2_u14_u4_U45 (.A( u2_u14_u4_n153 ) , .ZN( u2_u14_u4_n172 ) );
  NAND2_X1 u2_u14_u4_U46 (.A2( u2_u14_u4_n120 ) , .ZN( u2_u14_u4_n123 ) , .A1( u2_u14_u4_n161 ) );
  AOI22_X1 u2_u14_u4_U47 (.B2( u2_u14_u4_n132 ) , .A2( u2_u14_u4_n133 ) , .ZN( u2_u14_u4_n140 ) , .A1( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n179 ) );
  NAND2_X1 u2_u14_u4_U48 (.ZN( u2_u14_u4_n133 ) , .A2( u2_u14_u4_n146 ) , .A1( u2_u14_u4_n154 ) );
  NAND2_X1 u2_u14_u4_U49 (.A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n154 ) , .A2( u2_u14_u4_n98 ) );
  NOR4_X1 u2_u14_u4_U5 (.A4( u2_u14_u4_n106 ) , .A3( u2_u14_u4_n107 ) , .A2( u2_u14_u4_n108 ) , .A1( u2_u14_u4_n109 ) , .ZN( u2_u14_u4_n110 ) );
  NAND2_X1 u2_u14_u4_U50 (.A1( u2_u14_u4_n101 ) , .ZN( u2_u14_u4_n158 ) , .A2( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U51 (.ZN( u2_u14_u4_n127 ) , .A( u2_u14_u4_n136 ) , .B2( u2_u14_u4_n150 ) , .B1( u2_u14_u4_n180 ) );
  INV_X1 u2_u14_u4_U52 (.A( u2_u14_u4_n160 ) , .ZN( u2_u14_u4_n180 ) );
  NAND2_X1 u2_u14_u4_U53 (.A2( u2_u14_u4_n104 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n146 ) );
  NAND2_X1 u2_u14_u4_U54 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n160 ) );
  NAND2_X1 u2_u14_u4_U55 (.ZN( u2_u14_u4_n134 ) , .A1( u2_u14_u4_n98 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U56 (.A1( u2_u14_u4_n103 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n143 ) );
  NAND2_X1 u2_u14_u4_U57 (.A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n145 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U58 (.A1( u2_u14_u4_n100 ) , .A2( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n120 ) );
  NAND2_X1 u2_u14_u4_U59 (.A1( u2_u14_u4_n102 ) , .A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n148 ) );
  AOI21_X1 u2_u14_u4_U6 (.ZN( u2_u14_u4_n106 ) , .B2( u2_u14_u4_n146 ) , .B1( u2_u14_u4_n158 ) , .A( u2_u14_u4_n170 ) );
  NAND2_X1 u2_u14_u4_U60 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n157 ) );
  INV_X1 u2_u14_u4_U61 (.A( u2_u14_u4_n150 ) , .ZN( u2_u14_u4_n173 ) );
  INV_X1 u2_u14_u4_U62 (.A( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n171 ) );
  NAND2_X1 u2_u14_u4_U63 (.A1( u2_u14_u4_n100 ) , .ZN( u2_u14_u4_n118 ) , .A2( u2_u14_u4_n99 ) );
  NAND2_X1 u2_u14_u4_U64 (.A2( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n144 ) );
  NAND2_X1 u2_u14_u4_U65 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n105 ) , .ZN( u2_u14_u4_n96 ) );
  INV_X1 u2_u14_u4_U66 (.A( u2_u14_u4_n128 ) , .ZN( u2_u14_u4_n174 ) );
  NAND2_X1 u2_u14_u4_U67 (.A2( u2_u14_u4_n102 ) , .ZN( u2_u14_u4_n119 ) , .A1( u2_u14_u4_n98 ) );
  NAND2_X1 u2_u14_u4_U68 (.A2( u2_u14_u4_n101 ) , .A1( u2_u14_u4_n103 ) , .ZN( u2_u14_u4_n147 ) );
  NAND2_X1 u2_u14_u4_U69 (.A2( u2_u14_u4_n104 ) , .ZN( u2_u14_u4_n113 ) , .A1( u2_u14_u4_n99 ) );
  AOI21_X1 u2_u14_u4_U7 (.ZN( u2_u14_u4_n108 ) , .B2( u2_u14_u4_n134 ) , .B1( u2_u14_u4_n155 ) , .A( u2_u14_u4_n156 ) );
  NOR2_X1 u2_u14_u4_U70 (.A2( u2_u14_X_28 ) , .ZN( u2_u14_u4_n150 ) , .A1( u2_u14_u4_n168 ) );
  NOR2_X1 u2_u14_u4_U71 (.A2( u2_u14_X_29 ) , .ZN( u2_u14_u4_n152 ) , .A1( u2_u14_u4_n169 ) );
  NOR2_X1 u2_u14_u4_U72 (.A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n105 ) , .A1( u2_u14_u4_n176 ) );
  NOR2_X1 u2_u14_u4_U73 (.A2( u2_u14_X_26 ) , .ZN( u2_u14_u4_n100 ) , .A1( u2_u14_u4_n177 ) );
  NOR2_X1 u2_u14_u4_U74 (.A2( u2_u14_X_28 ) , .A1( u2_u14_X_29 ) , .ZN( u2_u14_u4_n128 ) );
  NOR2_X1 u2_u14_u4_U75 (.A2( u2_u14_X_27 ) , .A1( u2_u14_X_30 ) , .ZN( u2_u14_u4_n102 ) );
  NOR2_X1 u2_u14_u4_U76 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n98 ) );
  AND2_X1 u2_u14_u4_U77 (.A2( u2_u14_X_25 ) , .A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n104 ) );
  AND2_X1 u2_u14_u4_U78 (.A1( u2_u14_X_30 ) , .A2( u2_u14_u4_n176 ) , .ZN( u2_u14_u4_n99 ) );
  AND2_X1 u2_u14_u4_U79 (.A1( u2_u14_X_26 ) , .ZN( u2_u14_u4_n101 ) , .A2( u2_u14_u4_n177 ) );
  AOI21_X1 u2_u14_u4_U8 (.ZN( u2_u14_u4_n109 ) , .A( u2_u14_u4_n153 ) , .B1( u2_u14_u4_n159 ) , .B2( u2_u14_u4_n184 ) );
  AND2_X1 u2_u14_u4_U80 (.A1( u2_u14_X_27 ) , .A2( u2_u14_X_30 ) , .ZN( u2_u14_u4_n103 ) );
  INV_X1 u2_u14_u4_U81 (.A( u2_u14_X_28 ) , .ZN( u2_u14_u4_n169 ) );
  INV_X1 u2_u14_u4_U82 (.A( u2_u14_X_29 ) , .ZN( u2_u14_u4_n168 ) );
  INV_X1 u2_u14_u4_U83 (.A( u2_u14_X_25 ) , .ZN( u2_u14_u4_n177 ) );
  INV_X1 u2_u14_u4_U84 (.A( u2_u14_X_27 ) , .ZN( u2_u14_u4_n176 ) );
  NAND4_X1 u2_u14_u4_U85 (.ZN( u2_out14_25 ) , .A4( u2_u14_u4_n139 ) , .A3( u2_u14_u4_n140 ) , .A2( u2_u14_u4_n141 ) , .A1( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U86 (.A( u2_u14_u4_n128 ) , .B2( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n130 ) , .ZN( u2_u14_u4_n142 ) );
  OAI21_X1 u2_u14_u4_U87 (.B2( u2_u14_u4_n131 ) , .ZN( u2_u14_u4_n141 ) , .A( u2_u14_u4_n175 ) , .B1( u2_u14_u4_n183 ) );
  NAND4_X1 u2_u14_u4_U88 (.ZN( u2_out14_14 ) , .A4( u2_u14_u4_n124 ) , .A3( u2_u14_u4_n125 ) , .A2( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n127 ) );
  AOI22_X1 u2_u14_u4_U89 (.B2( u2_u14_u4_n117 ) , .ZN( u2_u14_u4_n126 ) , .A1( u2_u14_u4_n129 ) , .B1( u2_u14_u4_n152 ) , .A2( u2_u14_u4_n175 ) );
  AOI211_X1 u2_u14_u4_U9 (.B( u2_u14_u4_n136 ) , .A( u2_u14_u4_n137 ) , .C2( u2_u14_u4_n138 ) , .ZN( u2_u14_u4_n139 ) , .C1( u2_u14_u4_n182 ) );
  AOI22_X1 u2_u14_u4_U90 (.ZN( u2_u14_u4_n125 ) , .B2( u2_u14_u4_n131 ) , .A2( u2_u14_u4_n132 ) , .B1( u2_u14_u4_n138 ) , .A1( u2_u14_u4_n178 ) );
  NAND4_X1 u2_u14_u4_U91 (.ZN( u2_out14_8 ) , .A4( u2_u14_u4_n110 ) , .A3( u2_u14_u4_n111 ) , .A2( u2_u14_u4_n112 ) , .A1( u2_u14_u4_n186 ) );
  NAND2_X1 u2_u14_u4_U92 (.ZN( u2_u14_u4_n112 ) , .A2( u2_u14_u4_n130 ) , .A1( u2_u14_u4_n150 ) );
  AOI22_X1 u2_u14_u4_U93 (.ZN( u2_u14_u4_n111 ) , .B2( u2_u14_u4_n132 ) , .A1( u2_u14_u4_n152 ) , .B1( u2_u14_u4_n178 ) , .A2( u2_u14_u4_n97 ) );
  AOI22_X1 u2_u14_u4_U94 (.B2( u2_u14_u4_n149 ) , .B1( u2_u14_u4_n150 ) , .A2( u2_u14_u4_n151 ) , .A1( u2_u14_u4_n152 ) , .ZN( u2_u14_u4_n167 ) );
  NOR4_X1 u2_u14_u4_U95 (.A4( u2_u14_u4_n162 ) , .A3( u2_u14_u4_n163 ) , .A2( u2_u14_u4_n164 ) , .A1( u2_u14_u4_n165 ) , .ZN( u2_u14_u4_n166 ) );
  NAND3_X1 u2_u14_u4_U96 (.ZN( u2_out14_3 ) , .A3( u2_u14_u4_n166 ) , .A1( u2_u14_u4_n167 ) , .A2( u2_u14_u4_n186 ) );
  NAND3_X1 u2_u14_u4_U97 (.A3( u2_u14_u4_n146 ) , .A2( u2_u14_u4_n147 ) , .A1( u2_u14_u4_n148 ) , .ZN( u2_u14_u4_n149 ) );
  NAND3_X1 u2_u14_u4_U98 (.A3( u2_u14_u4_n143 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n145 ) , .ZN( u2_u14_u4_n151 ) );
  NAND3_X1 u2_u14_u4_U99 (.A3( u2_u14_u4_n121 ) , .ZN( u2_u14_u4_n122 ) , .A2( u2_u14_u4_n144 ) , .A1( u2_u14_u4_n154 ) );
  INV_X1 u2_u14_u5_U10 (.A( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U100 (.A3( u2_u14_u5_n141 ) , .A1( u2_u14_u5_n142 ) , .ZN( u2_u14_u5_n143 ) , .A2( u2_u14_u5_n191 ) );
  NAND4_X1 u2_u14_u5_U101 (.ZN( u2_out14_4 ) , .A4( u2_u14_u5_n112 ) , .A2( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n114 ) , .A3( u2_u14_u5_n195 ) );
  AOI211_X1 u2_u14_u5_U102 (.A( u2_u14_u5_n110 ) , .C1( u2_u14_u5_n111 ) , .ZN( u2_u14_u5_n112 ) , .B( u2_u14_u5_n118 ) , .C2( u2_u14_u5_n177 ) );
  AOI222_X1 u2_u14_u5_U103 (.ZN( u2_u14_u5_n113 ) , .A1( u2_u14_u5_n131 ) , .C1( u2_u14_u5_n148 ) , .B2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n178 ) , .A2( u2_u14_u5_n179 ) , .B1( u2_u14_u5_n99 ) );
  NAND3_X1 u2_u14_u5_U104 (.A2( u2_u14_u5_n154 ) , .A3( u2_u14_u5_n158 ) , .A1( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n99 ) );
  NOR2_X1 u2_u14_u5_U11 (.ZN( u2_u14_u5_n160 ) , .A2( u2_u14_u5_n173 ) , .A1( u2_u14_u5_n177 ) );
  INV_X1 u2_u14_u5_U12 (.A( u2_u14_u5_n150 ) , .ZN( u2_u14_u5_n174 ) );
  AOI21_X1 u2_u14_u5_U13 (.A( u2_u14_u5_n160 ) , .B2( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n162 ) , .B1( u2_u14_u5_n192 ) );
  INV_X1 u2_u14_u5_U14 (.A( u2_u14_u5_n159 ) , .ZN( u2_u14_u5_n192 ) );
  AOI21_X1 u2_u14_u5_U15 (.A( u2_u14_u5_n156 ) , .B2( u2_u14_u5_n157 ) , .B1( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n163 ) );
  AOI21_X1 u2_u14_u5_U16 (.B2( u2_u14_u5_n139 ) , .B1( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n141 ) , .A( u2_u14_u5_n150 ) );
  OAI21_X1 u2_u14_u5_U17 (.A( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n134 ) , .B1( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n142 ) );
  OAI21_X1 u2_u14_u5_U18 (.ZN( u2_u14_u5_n133 ) , .B2( u2_u14_u5_n147 ) , .A( u2_u14_u5_n173 ) , .B1( u2_u14_u5_n188 ) );
  NAND2_X1 u2_u14_u5_U19 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n137 ) );
  INV_X1 u2_u14_u5_U20 (.A( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n194 ) );
  NAND2_X1 u2_u14_u5_U21 (.A1( u2_u14_u5_n121 ) , .ZN( u2_u14_u5_n132 ) , .A2( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U22 (.A2( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n136 ) , .A1( u2_u14_u5_n154 ) );
  NAND2_X1 u2_u14_u5_U23 (.A2( u2_u14_u5_n119 ) , .A1( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n159 ) );
  INV_X1 u2_u14_u5_U24 (.A( u2_u14_u5_n156 ) , .ZN( u2_u14_u5_n175 ) );
  INV_X1 u2_u14_u5_U25 (.A( u2_u14_u5_n158 ) , .ZN( u2_u14_u5_n188 ) );
  INV_X1 u2_u14_u5_U26 (.A( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n179 ) );
  INV_X1 u2_u14_u5_U27 (.A( u2_u14_u5_n140 ) , .ZN( u2_u14_u5_n182 ) );
  INV_X1 u2_u14_u5_U28 (.A( u2_u14_u5_n151 ) , .ZN( u2_u14_u5_n183 ) );
  INV_X1 u2_u14_u5_U29 (.A( u2_u14_u5_n123 ) , .ZN( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U3 (.ZN( u2_u14_u5_n134 ) , .A1( u2_u14_u5_n183 ) , .A2( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U30 (.A( u2_u14_u5_n161 ) , .ZN( u2_u14_u5_n184 ) );
  INV_X1 u2_u14_u5_U31 (.A( u2_u14_u5_n139 ) , .ZN( u2_u14_u5_n189 ) );
  INV_X1 u2_u14_u5_U32 (.A( u2_u14_u5_n157 ) , .ZN( u2_u14_u5_n190 ) );
  INV_X1 u2_u14_u5_U33 (.A( u2_u14_u5_n120 ) , .ZN( u2_u14_u5_n193 ) );
  NAND2_X1 u2_u14_u5_U34 (.ZN( u2_u14_u5_n111 ) , .A1( u2_u14_u5_n140 ) , .A2( u2_u14_u5_n155 ) );
  INV_X1 u2_u14_u5_U35 (.A( u2_u14_u5_n117 ) , .ZN( u2_u14_u5_n196 ) );
  OAI221_X1 u2_u14_u5_U36 (.A( u2_u14_u5_n116 ) , .ZN( u2_u14_u5_n117 ) , .B2( u2_u14_u5_n119 ) , .C1( u2_u14_u5_n153 ) , .C2( u2_u14_u5_n158 ) , .B1( u2_u14_u5_n172 ) );
  AOI222_X1 u2_u14_u5_U37 (.ZN( u2_u14_u5_n116 ) , .B2( u2_u14_u5_n145 ) , .C1( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n174 ) , .C2( u2_u14_u5_n177 ) , .B1( u2_u14_u5_n187 ) , .A1( u2_u14_u5_n193 ) );
  INV_X1 u2_u14_u5_U38 (.A( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n187 ) );
  NOR2_X1 u2_u14_u5_U39 (.ZN( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n170 ) , .A2( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U4 (.A( u2_u14_u5_n138 ) , .ZN( u2_u14_u5_n191 ) );
  AOI22_X1 u2_u14_u5_U40 (.B2( u2_u14_u5_n131 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n169 ) , .B1( u2_u14_u5_n174 ) , .A1( u2_u14_u5_n185 ) );
  NOR2_X1 u2_u14_u5_U41 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n173 ) );
  AOI21_X1 u2_u14_u5_U42 (.A( u2_u14_u5_n118 ) , .B2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n168 ) , .B1( u2_u14_u5_n186 ) );
  INV_X1 u2_u14_u5_U43 (.A( u2_u14_u5_n122 ) , .ZN( u2_u14_u5_n186 ) );
  NOR2_X1 u2_u14_u5_U44 (.A1( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n152 ) , .A2( u2_u14_u5_n176 ) );
  NOR2_X1 u2_u14_u5_U45 (.A1( u2_u14_u5_n115 ) , .ZN( u2_u14_u5_n118 ) , .A2( u2_u14_u5_n153 ) );
  NOR2_X1 u2_u14_u5_U46 (.A2( u2_u14_u5_n145 ) , .ZN( u2_u14_u5_n156 ) , .A1( u2_u14_u5_n174 ) );
  NOR2_X1 u2_u14_u5_U47 (.ZN( u2_u14_u5_n121 ) , .A2( u2_u14_u5_n145 ) , .A1( u2_u14_u5_n176 ) );
  AOI22_X1 u2_u14_u5_U48 (.ZN( u2_u14_u5_n114 ) , .A2( u2_u14_u5_n137 ) , .A1( u2_u14_u5_n145 ) , .B2( u2_u14_u5_n175 ) , .B1( u2_u14_u5_n193 ) );
  OAI211_X1 u2_u14_u5_U49 (.B( u2_u14_u5_n124 ) , .A( u2_u14_u5_n125 ) , .C2( u2_u14_u5_n126 ) , .C1( u2_u14_u5_n127 ) , .ZN( u2_u14_u5_n128 ) );
  OAI21_X1 u2_u14_u5_U5 (.B2( u2_u14_u5_n136 ) , .B1( u2_u14_u5_n137 ) , .ZN( u2_u14_u5_n138 ) , .A( u2_u14_u5_n177 ) );
  NOR3_X1 u2_u14_u5_U50 (.ZN( u2_u14_u5_n127 ) , .A1( u2_u14_u5_n136 ) , .A3( u2_u14_u5_n148 ) , .A2( u2_u14_u5_n182 ) );
  OAI21_X1 u2_u14_u5_U51 (.ZN( u2_u14_u5_n124 ) , .A( u2_u14_u5_n177 ) , .B2( u2_u14_u5_n183 ) , .B1( u2_u14_u5_n189 ) );
  OAI21_X1 u2_u14_u5_U52 (.ZN( u2_u14_u5_n125 ) , .A( u2_u14_u5_n174 ) , .B2( u2_u14_u5_n185 ) , .B1( u2_u14_u5_n190 ) );
  AOI21_X1 u2_u14_u5_U53 (.A( u2_u14_u5_n153 ) , .B2( u2_u14_u5_n154 ) , .B1( u2_u14_u5_n155 ) , .ZN( u2_u14_u5_n164 ) );
  AOI21_X1 u2_u14_u5_U54 (.ZN( u2_u14_u5_n110 ) , .B1( u2_u14_u5_n122 ) , .B2( u2_u14_u5_n139 ) , .A( u2_u14_u5_n153 ) );
  INV_X1 u2_u14_u5_U55 (.A( u2_u14_u5_n153 ) , .ZN( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U56 (.A( u2_u14_u5_n126 ) , .ZN( u2_u14_u5_n173 ) );
  AND2_X1 u2_u14_u5_U57 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n147 ) );
  AND2_X1 u2_u14_u5_U58 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n148 ) );
  NAND2_X1 u2_u14_u5_U59 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n158 ) );
  INV_X1 u2_u14_u5_U6 (.A( u2_u14_u5_n135 ) , .ZN( u2_u14_u5_n178 ) );
  NAND2_X1 u2_u14_u5_U60 (.A2( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n139 ) );
  NAND2_X1 u2_u14_u5_U61 (.A1( u2_u14_u5_n106 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n119 ) );
  NAND2_X1 u2_u14_u5_U62 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n140 ) );
  NAND2_X1 u2_u14_u5_U63 (.A2( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n105 ) , .ZN( u2_u14_u5_n155 ) );
  NAND2_X1 u2_u14_u5_U64 (.A2( u2_u14_u5_n106 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n122 ) );
  NAND2_X1 u2_u14_u5_U65 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n106 ) , .ZN( u2_u14_u5_n115 ) );
  NAND2_X1 u2_u14_u5_U66 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n103 ) , .ZN( u2_u14_u5_n161 ) );
  NAND2_X1 u2_u14_u5_U67 (.A1( u2_u14_u5_n105 ) , .A2( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n154 ) );
  INV_X1 u2_u14_u5_U68 (.A( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n172 ) );
  NAND2_X1 u2_u14_u5_U69 (.A1( u2_u14_u5_n103 ) , .A2( u2_u14_u5_n108 ) , .ZN( u2_u14_u5_n123 ) );
  OAI22_X1 u2_u14_u5_U7 (.B2( u2_u14_u5_n149 ) , .B1( u2_u14_u5_n150 ) , .A2( u2_u14_u5_n151 ) , .A1( u2_u14_u5_n152 ) , .ZN( u2_u14_u5_n165 ) );
  NAND2_X1 u2_u14_u5_U70 (.A2( u2_u14_u5_n103 ) , .A1( u2_u14_u5_n107 ) , .ZN( u2_u14_u5_n151 ) );
  NAND2_X1 u2_u14_u5_U71 (.A2( u2_u14_u5_n107 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n120 ) );
  NAND2_X1 u2_u14_u5_U72 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n109 ) , .ZN( u2_u14_u5_n157 ) );
  AND2_X1 u2_u14_u5_U73 (.A2( u2_u14_u5_n100 ) , .A1( u2_u14_u5_n104 ) , .ZN( u2_u14_u5_n131 ) );
  INV_X1 u2_u14_u5_U74 (.A( u2_u14_u5_n102 ) , .ZN( u2_u14_u5_n195 ) );
  OAI221_X1 u2_u14_u5_U75 (.A( u2_u14_u5_n101 ) , .ZN( u2_u14_u5_n102 ) , .C2( u2_u14_u5_n115 ) , .C1( u2_u14_u5_n126 ) , .B1( u2_u14_u5_n134 ) , .B2( u2_u14_u5_n160 ) );
  OAI21_X1 u2_u14_u5_U76 (.ZN( u2_u14_u5_n101 ) , .B1( u2_u14_u5_n137 ) , .A( u2_u14_u5_n146 ) , .B2( u2_u14_u5_n147 ) );
  NOR2_X1 u2_u14_u5_U77 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n145 ) );
  NOR2_X1 u2_u14_u5_U78 (.A2( u2_u14_X_34 ) , .ZN( u2_u14_u5_n146 ) , .A1( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U79 (.A2( u2_u14_X_31 ) , .A1( u2_u14_X_32 ) , .ZN( u2_u14_u5_n103 ) );
  NOR3_X1 u2_u14_u5_U8 (.A2( u2_u14_u5_n147 ) , .A1( u2_u14_u5_n148 ) , .ZN( u2_u14_u5_n149 ) , .A3( u2_u14_u5_n194 ) );
  NOR2_X1 u2_u14_u5_U80 (.A2( u2_u14_X_36 ) , .ZN( u2_u14_u5_n105 ) , .A1( u2_u14_u5_n180 ) );
  NOR2_X1 u2_u14_u5_U81 (.A2( u2_u14_X_33 ) , .ZN( u2_u14_u5_n108 ) , .A1( u2_u14_u5_n170 ) );
  NOR2_X1 u2_u14_u5_U82 (.A2( u2_u14_X_33 ) , .A1( u2_u14_X_36 ) , .ZN( u2_u14_u5_n107 ) );
  NOR2_X1 u2_u14_u5_U83 (.A2( u2_u14_X_31 ) , .ZN( u2_u14_u5_n104 ) , .A1( u2_u14_u5_n181 ) );
  NAND2_X1 u2_u14_u5_U84 (.A2( u2_u14_X_34 ) , .A1( u2_u14_X_35 ) , .ZN( u2_u14_u5_n153 ) );
  NAND2_X1 u2_u14_u5_U85 (.A1( u2_u14_X_34 ) , .ZN( u2_u14_u5_n126 ) , .A2( u2_u14_u5_n171 ) );
  AND2_X1 u2_u14_u5_U86 (.A1( u2_u14_X_31 ) , .A2( u2_u14_X_32 ) , .ZN( u2_u14_u5_n106 ) );
  AND2_X1 u2_u14_u5_U87 (.A1( u2_u14_X_31 ) , .ZN( u2_u14_u5_n109 ) , .A2( u2_u14_u5_n181 ) );
  INV_X1 u2_u14_u5_U88 (.A( u2_u14_X_33 ) , .ZN( u2_u14_u5_n180 ) );
  INV_X1 u2_u14_u5_U89 (.A( u2_u14_X_35 ) , .ZN( u2_u14_u5_n171 ) );
  NOR2_X1 u2_u14_u5_U9 (.ZN( u2_u14_u5_n135 ) , .A1( u2_u14_u5_n173 ) , .A2( u2_u14_u5_n176 ) );
  INV_X1 u2_u14_u5_U90 (.A( u2_u14_X_36 ) , .ZN( u2_u14_u5_n170 ) );
  INV_X1 u2_u14_u5_U91 (.A( u2_u14_X_32 ) , .ZN( u2_u14_u5_n181 ) );
  NAND4_X1 u2_u14_u5_U92 (.ZN( u2_out14_29 ) , .A4( u2_u14_u5_n129 ) , .A3( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n196 ) );
  AOI221_X1 u2_u14_u5_U93 (.A( u2_u14_u5_n128 ) , .ZN( u2_u14_u5_n129 ) , .C2( u2_u14_u5_n132 ) , .B2( u2_u14_u5_n159 ) , .B1( u2_u14_u5_n176 ) , .C1( u2_u14_u5_n184 ) );
  AOI222_X1 u2_u14_u5_U94 (.ZN( u2_u14_u5_n130 ) , .A2( u2_u14_u5_n146 ) , .B1( u2_u14_u5_n147 ) , .C2( u2_u14_u5_n175 ) , .B2( u2_u14_u5_n179 ) , .A1( u2_u14_u5_n188 ) , .C1( u2_u14_u5_n194 ) );
  NAND4_X1 u2_u14_u5_U95 (.ZN( u2_out14_19 ) , .A4( u2_u14_u5_n166 ) , .A3( u2_u14_u5_n167 ) , .A2( u2_u14_u5_n168 ) , .A1( u2_u14_u5_n169 ) );
  AOI22_X1 u2_u14_u5_U96 (.B2( u2_u14_u5_n145 ) , .A2( u2_u14_u5_n146 ) , .ZN( u2_u14_u5_n167 ) , .B1( u2_u14_u5_n182 ) , .A1( u2_u14_u5_n189 ) );
  NOR4_X1 u2_u14_u5_U97 (.A4( u2_u14_u5_n162 ) , .A3( u2_u14_u5_n163 ) , .A2( u2_u14_u5_n164 ) , .A1( u2_u14_u5_n165 ) , .ZN( u2_u14_u5_n166 ) );
  NAND4_X1 u2_u14_u5_U98 (.ZN( u2_out14_11 ) , .A4( u2_u14_u5_n143 ) , .A3( u2_u14_u5_n144 ) , .A2( u2_u14_u5_n169 ) , .A1( u2_u14_u5_n196 ) );
  AOI22_X1 u2_u14_u5_U99 (.A2( u2_u14_u5_n132 ) , .ZN( u2_u14_u5_n144 ) , .B2( u2_u14_u5_n145 ) , .B1( u2_u14_u5_n184 ) , .A1( u2_u14_u5_n194 ) );
  AOI22_X1 u2_u14_u6_U10 (.A2( u2_u14_u6_n151 ) , .B2( u2_u14_u6_n161 ) , .A1( u2_u14_u6_n167 ) , .B1( u2_u14_u6_n170 ) , .ZN( u2_u14_u6_n89 ) );
  AOI21_X1 u2_u14_u6_U11 (.B1( u2_u14_u6_n107 ) , .B2( u2_u14_u6_n132 ) , .A( u2_u14_u6_n158 ) , .ZN( u2_u14_u6_n88 ) );
  AOI21_X1 u2_u14_u6_U12 (.B2( u2_u14_u6_n147 ) , .B1( u2_u14_u6_n148 ) , .ZN( u2_u14_u6_n149 ) , .A( u2_u14_u6_n158 ) );
  AOI21_X1 u2_u14_u6_U13 (.ZN( u2_u14_u6_n106 ) , .A( u2_u14_u6_n142 ) , .B2( u2_u14_u6_n159 ) , .B1( u2_u14_u6_n164 ) );
  INV_X1 u2_u14_u6_U14 (.A( u2_u14_u6_n155 ) , .ZN( u2_u14_u6_n161 ) );
  INV_X1 u2_u14_u6_U15 (.A( u2_u14_u6_n128 ) , .ZN( u2_u14_u6_n164 ) );
  NAND2_X1 u2_u14_u6_U16 (.ZN( u2_u14_u6_n110 ) , .A1( u2_u14_u6_n122 ) , .A2( u2_u14_u6_n129 ) );
  NAND2_X1 u2_u14_u6_U17 (.ZN( u2_u14_u6_n124 ) , .A2( u2_u14_u6_n146 ) , .A1( u2_u14_u6_n148 ) );
  INV_X1 u2_u14_u6_U18 (.A( u2_u14_u6_n132 ) , .ZN( u2_u14_u6_n171 ) );
  AND2_X1 u2_u14_u6_U19 (.A1( u2_u14_u6_n100 ) , .ZN( u2_u14_u6_n130 ) , .A2( u2_u14_u6_n147 ) );
  INV_X1 u2_u14_u6_U20 (.A( u2_u14_u6_n127 ) , .ZN( u2_u14_u6_n173 ) );
  INV_X1 u2_u14_u6_U21 (.A( u2_u14_u6_n121 ) , .ZN( u2_u14_u6_n167 ) );
  INV_X1 u2_u14_u6_U22 (.A( u2_u14_u6_n100 ) , .ZN( u2_u14_u6_n169 ) );
  INV_X1 u2_u14_u6_U23 (.A( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n170 ) );
  INV_X1 u2_u14_u6_U24 (.A( u2_u14_u6_n113 ) , .ZN( u2_u14_u6_n168 ) );
  AND2_X1 u2_u14_u6_U25 (.A1( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n119 ) , .ZN( u2_u14_u6_n133 ) );
  AND2_X1 u2_u14_u6_U26 (.A2( u2_u14_u6_n121 ) , .A1( u2_u14_u6_n122 ) , .ZN( u2_u14_u6_n131 ) );
  AND3_X1 u2_u14_u6_U27 (.ZN( u2_u14_u6_n120 ) , .A2( u2_u14_u6_n127 ) , .A1( u2_u14_u6_n132 ) , .A3( u2_u14_u6_n145 ) );
  INV_X1 u2_u14_u6_U28 (.A( u2_u14_u6_n146 ) , .ZN( u2_u14_u6_n163 ) );
  AOI222_X1 u2_u14_u6_U29 (.ZN( u2_u14_u6_n114 ) , .A1( u2_u14_u6_n118 ) , .A2( u2_u14_u6_n126 ) , .B2( u2_u14_u6_n151 ) , .C2( u2_u14_u6_n159 ) , .C1( u2_u14_u6_n168 ) , .B1( u2_u14_u6_n169 ) );
  INV_X1 u2_u14_u6_U3 (.A( u2_u14_u6_n110 ) , .ZN( u2_u14_u6_n166 ) );
  NOR2_X1 u2_u14_u6_U30 (.A1( u2_u14_u6_n162 ) , .A2( u2_u14_u6_n165 ) , .ZN( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U31 (.A1( u2_u14_u6_n144 ) , .ZN( u2_u14_u6_n151 ) , .A2( u2_u14_u6_n158 ) );
  NAND2_X1 u2_u14_u6_U32 (.ZN( u2_u14_u6_n132 ) , .A1( u2_u14_u6_n91 ) , .A2( u2_u14_u6_n97 ) );
  AOI22_X1 u2_u14_u6_U33 (.B2( u2_u14_u6_n110 ) , .B1( u2_u14_u6_n111 ) , .A1( u2_u14_u6_n112 ) , .ZN( u2_u14_u6_n115 ) , .A2( u2_u14_u6_n161 ) );
  NAND4_X1 u2_u14_u6_U34 (.A3( u2_u14_u6_n109 ) , .ZN( u2_u14_u6_n112 ) , .A4( u2_u14_u6_n132 ) , .A2( u2_u14_u6_n147 ) , .A1( u2_u14_u6_n166 ) );
  NOR2_X1 u2_u14_u6_U35 (.ZN( u2_u14_u6_n109 ) , .A1( u2_u14_u6_n170 ) , .A2( u2_u14_u6_n173 ) );
  NOR2_X1 u2_u14_u6_U36 (.A2( u2_u14_u6_n126 ) , .ZN( u2_u14_u6_n155 ) , .A1( u2_u14_u6_n160 ) );
  NAND2_X1 u2_u14_u6_U37 (.ZN( u2_u14_u6_n146 ) , .A2( u2_u14_u6_n94 ) , .A1( u2_u14_u6_n99 ) );
  AOI21_X1 u2_u14_u6_U38 (.A( u2_u14_u6_n144 ) , .B2( u2_u14_u6_n145 ) , .B1( u2_u14_u6_n146 ) , .ZN( u2_u14_u6_n150 ) );
  AOI211_X1 u2_u14_u6_U39 (.B( u2_u14_u6_n134 ) , .A( u2_u14_u6_n135 ) , .C1( u2_u14_u6_n136 ) , .ZN( u2_u14_u6_n137 ) , .C2( u2_u14_u6_n151 ) );
  INV_X1 u2_u14_u6_U4 (.A( u2_u14_u6_n142 ) , .ZN( u2_u14_u6_n174 ) );
  AOI21_X1 u2_u14_u6_U40 (.B2( u2_u14_u6_n132 ) , .B1( u2_u14_u6_n133 ) , .ZN( u2_u14_u6_n134 ) , .A( u2_u14_u6_n158 ) );
  NAND4_X1 u2_u14_u6_U41 (.A4( u2_u14_u6_n127 ) , .A3( u2_u14_u6_n128 ) , .A2( u2_u14_u6_n129 ) , .A1( u2_u14_u6_n130 ) , .ZN( u2_u14_u6_n136 ) );
  AOI21_X1 u2_u14_u6_U42 (.B1( u2_u14_u6_n131 ) , .ZN( u2_u14_u6_n135 ) , .A( u2_u14_u6_n144 ) , .B2( u2_u14_u6_n146 ) );
  INV_X1 u2_u14_u6_U43 (.A( u2_u14_u6_n111 ) , .ZN( u2_u14_u6_n158 ) );
  NAND2_X1 u2_u14_u6_U44 (.ZN( u2_u14_u6_n127 ) , .A1( u2_u14_u6_n91 ) , .A2( u2_u14_u6_n92 ) );
  NAND2_X1 u2_u14_u6_U45 (.ZN( u2_u14_u6_n129 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n96 ) );
  INV_X1 u2_u14_u6_U46 (.A( u2_u14_u6_n144 ) , .ZN( u2_u14_u6_n159 ) );
  NAND2_X1 u2_u14_u6_U47 (.ZN( u2_u14_u6_n145 ) , .A2( u2_u14_u6_n97 ) , .A1( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U48 (.ZN( u2_u14_u6_n148 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n94 ) );
  NAND2_X1 u2_u14_u6_U49 (.ZN( u2_u14_u6_n108 ) , .A2( u2_u14_u6_n139 ) , .A1( u2_u14_u6_n144 ) );
  NAND2_X1 u2_u14_u6_U5 (.A2( u2_u14_u6_n143 ) , .ZN( u2_u14_u6_n152 ) , .A1( u2_u14_u6_n166 ) );
  NAND2_X1 u2_u14_u6_U50 (.ZN( u2_u14_u6_n121 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n97 ) );
  NAND2_X1 u2_u14_u6_U51 (.ZN( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n95 ) );
  AND2_X1 u2_u14_u6_U52 (.ZN( u2_u14_u6_n118 ) , .A2( u2_u14_u6_n91 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U53 (.ZN( u2_u14_u6_n147 ) , .A2( u2_u14_u6_n98 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U54 (.ZN( u2_u14_u6_n128 ) , .A1( u2_u14_u6_n94 ) , .A2( u2_u14_u6_n96 ) );
  NAND2_X1 u2_u14_u6_U55 (.ZN( u2_u14_u6_n119 ) , .A2( u2_u14_u6_n95 ) , .A1( u2_u14_u6_n99 ) );
  NAND2_X1 u2_u14_u6_U56 (.ZN( u2_u14_u6_n123 ) , .A2( u2_u14_u6_n91 ) , .A1( u2_u14_u6_n96 ) );
  NAND2_X1 u2_u14_u6_U57 (.ZN( u2_u14_u6_n100 ) , .A2( u2_u14_u6_n92 ) , .A1( u2_u14_u6_n98 ) );
  NAND2_X1 u2_u14_u6_U58 (.ZN( u2_u14_u6_n122 ) , .A1( u2_u14_u6_n94 ) , .A2( u2_u14_u6_n97 ) );
  INV_X1 u2_u14_u6_U59 (.A( u2_u14_u6_n139 ) , .ZN( u2_u14_u6_n160 ) );
  AOI22_X1 u2_u14_u6_U6 (.B2( u2_u14_u6_n101 ) , .A1( u2_u14_u6_n102 ) , .ZN( u2_u14_u6_n103 ) , .B1( u2_u14_u6_n160 ) , .A2( u2_u14_u6_n161 ) );
  NAND2_X1 u2_u14_u6_U60 (.ZN( u2_u14_u6_n113 ) , .A1( u2_u14_u6_n96 ) , .A2( u2_u14_u6_n98 ) );
  NOR2_X1 u2_u14_u6_U61 (.A2( u2_u14_X_40 ) , .A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n126 ) );
  NOR2_X1 u2_u14_u6_U62 (.A2( u2_u14_X_39 ) , .A1( u2_u14_X_42 ) , .ZN( u2_u14_u6_n92 ) );
  NOR2_X1 u2_u14_u6_U63 (.A2( u2_u14_X_39 ) , .A1( u2_u14_u6_n156 ) , .ZN( u2_u14_u6_n97 ) );
  NOR2_X1 u2_u14_u6_U64 (.A2( u2_u14_X_38 ) , .A1( u2_u14_u6_n165 ) , .ZN( u2_u14_u6_n95 ) );
  NOR2_X1 u2_u14_u6_U65 (.A2( u2_u14_X_41 ) , .ZN( u2_u14_u6_n111 ) , .A1( u2_u14_u6_n157 ) );
  NOR2_X1 u2_u14_u6_U66 (.A2( u2_u14_X_37 ) , .A1( u2_u14_u6_n162 ) , .ZN( u2_u14_u6_n94 ) );
  NOR2_X1 u2_u14_u6_U67 (.A2( u2_u14_X_37 ) , .A1( u2_u14_X_38 ) , .ZN( u2_u14_u6_n91 ) );
  NAND2_X1 u2_u14_u6_U68 (.A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n144 ) , .A2( u2_u14_u6_n157 ) );
  NAND2_X1 u2_u14_u6_U69 (.A2( u2_u14_X_40 ) , .A1( u2_u14_X_41 ) , .ZN( u2_u14_u6_n139 ) );
  NOR2_X1 u2_u14_u6_U7 (.A1( u2_u14_u6_n118 ) , .ZN( u2_u14_u6_n143 ) , .A2( u2_u14_u6_n168 ) );
  AND2_X1 u2_u14_u6_U70 (.A1( u2_u14_X_39 ) , .A2( u2_u14_u6_n156 ) , .ZN( u2_u14_u6_n96 ) );
  AND2_X1 u2_u14_u6_U71 (.A1( u2_u14_X_39 ) , .A2( u2_u14_X_42 ) , .ZN( u2_u14_u6_n99 ) );
  INV_X1 u2_u14_u6_U72 (.A( u2_u14_X_40 ) , .ZN( u2_u14_u6_n157 ) );
  INV_X1 u2_u14_u6_U73 (.A( u2_u14_X_37 ) , .ZN( u2_u14_u6_n165 ) );
  INV_X1 u2_u14_u6_U74 (.A( u2_u14_X_38 ) , .ZN( u2_u14_u6_n162 ) );
  INV_X1 u2_u14_u6_U75 (.A( u2_u14_X_42 ) , .ZN( u2_u14_u6_n156 ) );
  NAND4_X1 u2_u14_u6_U76 (.ZN( u2_out14_32 ) , .A4( u2_u14_u6_n103 ) , .A3( u2_u14_u6_n104 ) , .A2( u2_u14_u6_n105 ) , .A1( u2_u14_u6_n106 ) );
  AOI22_X1 u2_u14_u6_U77 (.ZN( u2_u14_u6_n105 ) , .A2( u2_u14_u6_n108 ) , .A1( u2_u14_u6_n118 ) , .B2( u2_u14_u6_n126 ) , .B1( u2_u14_u6_n171 ) );
  AOI22_X1 u2_u14_u6_U78 (.ZN( u2_u14_u6_n104 ) , .A1( u2_u14_u6_n111 ) , .B1( u2_u14_u6_n124 ) , .B2( u2_u14_u6_n151 ) , .A2( u2_u14_u6_n93 ) );
  NAND4_X1 u2_u14_u6_U79 (.ZN( u2_out14_12 ) , .A4( u2_u14_u6_n114 ) , .A3( u2_u14_u6_n115 ) , .A2( u2_u14_u6_n116 ) , .A1( u2_u14_u6_n117 ) );
  INV_X1 u2_u14_u6_U8 (.ZN( u2_u14_u6_n172 ) , .A( u2_u14_u6_n88 ) );
  OAI22_X1 u2_u14_u6_U80 (.B2( u2_u14_u6_n111 ) , .ZN( u2_u14_u6_n116 ) , .B1( u2_u14_u6_n126 ) , .A2( u2_u14_u6_n164 ) , .A1( u2_u14_u6_n167 ) );
  OAI21_X1 u2_u14_u6_U81 (.A( u2_u14_u6_n108 ) , .ZN( u2_u14_u6_n117 ) , .B2( u2_u14_u6_n141 ) , .B1( u2_u14_u6_n163 ) );
  OAI211_X1 u2_u14_u6_U82 (.ZN( u2_out14_22 ) , .B( u2_u14_u6_n137 ) , .A( u2_u14_u6_n138 ) , .C2( u2_u14_u6_n139 ) , .C1( u2_u14_u6_n140 ) );
  AOI22_X1 u2_u14_u6_U83 (.B1( u2_u14_u6_n124 ) , .A2( u2_u14_u6_n125 ) , .A1( u2_u14_u6_n126 ) , .ZN( u2_u14_u6_n138 ) , .B2( u2_u14_u6_n161 ) );
  AND4_X1 u2_u14_u6_U84 (.A3( u2_u14_u6_n119 ) , .A1( u2_u14_u6_n120 ) , .A4( u2_u14_u6_n129 ) , .ZN( u2_u14_u6_n140 ) , .A2( u2_u14_u6_n143 ) );
  OAI211_X1 u2_u14_u6_U85 (.ZN( u2_out14_7 ) , .B( u2_u14_u6_n153 ) , .C2( u2_u14_u6_n154 ) , .C1( u2_u14_u6_n155 ) , .A( u2_u14_u6_n174 ) );
  NOR3_X1 u2_u14_u6_U86 (.A1( u2_u14_u6_n141 ) , .ZN( u2_u14_u6_n154 ) , .A3( u2_u14_u6_n164 ) , .A2( u2_u14_u6_n171 ) );
  AOI211_X1 u2_u14_u6_U87 (.B( u2_u14_u6_n149 ) , .A( u2_u14_u6_n150 ) , .C2( u2_u14_u6_n151 ) , .C1( u2_u14_u6_n152 ) , .ZN( u2_u14_u6_n153 ) );
  NAND3_X1 u2_u14_u6_U88 (.A2( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n125 ) , .A1( u2_u14_u6_n130 ) , .A3( u2_u14_u6_n131 ) );
  NAND3_X1 u2_u14_u6_U89 (.A3( u2_u14_u6_n133 ) , .ZN( u2_u14_u6_n141 ) , .A1( u2_u14_u6_n145 ) , .A2( u2_u14_u6_n148 ) );
  OAI21_X1 u2_u14_u6_U9 (.A( u2_u14_u6_n159 ) , .B1( u2_u14_u6_n169 ) , .B2( u2_u14_u6_n173 ) , .ZN( u2_u14_u6_n90 ) );
  NAND3_X1 u2_u14_u6_U90 (.ZN( u2_u14_u6_n101 ) , .A3( u2_u14_u6_n107 ) , .A2( u2_u14_u6_n121 ) , .A1( u2_u14_u6_n127 ) );
  NAND3_X1 u2_u14_u6_U91 (.ZN( u2_u14_u6_n102 ) , .A3( u2_u14_u6_n130 ) , .A2( u2_u14_u6_n145 ) , .A1( u2_u14_u6_n166 ) );
  NAND3_X1 u2_u14_u6_U92 (.A3( u2_u14_u6_n113 ) , .A1( u2_u14_u6_n119 ) , .A2( u2_u14_u6_n123 ) , .ZN( u2_u14_u6_n93 ) );
  NAND3_X1 u2_u14_u6_U93 (.ZN( u2_u14_u6_n142 ) , .A2( u2_u14_u6_n172 ) , .A3( u2_u14_u6_n89 ) , .A1( u2_u14_u6_n90 ) );
  OAI21_X1 u2_u14_u7_U10 (.A( u2_u14_u7_n161 ) , .B1( u2_u14_u7_n168 ) , .B2( u2_u14_u7_n173 ) , .ZN( u2_u14_u7_n91 ) );
  AOI211_X1 u2_u14_u7_U11 (.A( u2_u14_u7_n117 ) , .ZN( u2_u14_u7_n118 ) , .C2( u2_u14_u7_n126 ) , .C1( u2_u14_u7_n177 ) , .B( u2_u14_u7_n180 ) );
  OAI22_X1 u2_u14_u7_U12 (.B1( u2_u14_u7_n115 ) , .ZN( u2_u14_u7_n117 ) , .A2( u2_u14_u7_n133 ) , .A1( u2_u14_u7_n137 ) , .B2( u2_u14_u7_n162 ) );
  INV_X1 u2_u14_u7_U13 (.A( u2_u14_u7_n116 ) , .ZN( u2_u14_u7_n180 ) );
  NOR3_X1 u2_u14_u7_U14 (.ZN( u2_u14_u7_n115 ) , .A3( u2_u14_u7_n145 ) , .A2( u2_u14_u7_n168 ) , .A1( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U15 (.A( u2_u14_u7_n133 ) , .ZN( u2_u14_u7_n176 ) );
  NOR3_X1 u2_u14_u7_U16 (.A2( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n135 ) , .ZN( u2_u14_u7_n136 ) , .A3( u2_u14_u7_n171 ) );
  NOR2_X1 u2_u14_u7_U17 (.A1( u2_u14_u7_n130 ) , .A2( u2_u14_u7_n134 ) , .ZN( u2_u14_u7_n153 ) );
  AOI21_X1 u2_u14_u7_U18 (.ZN( u2_u14_u7_n104 ) , .B2( u2_u14_u7_n112 ) , .B1( u2_u14_u7_n127 ) , .A( u2_u14_u7_n164 ) );
  AOI21_X1 u2_u14_u7_U19 (.ZN( u2_u14_u7_n106 ) , .B1( u2_u14_u7_n133 ) , .B2( u2_u14_u7_n146 ) , .A( u2_u14_u7_n162 ) );
  AOI21_X1 u2_u14_u7_U20 (.A( u2_u14_u7_n101 ) , .ZN( u2_u14_u7_n107 ) , .B2( u2_u14_u7_n128 ) , .B1( u2_u14_u7_n175 ) );
  INV_X1 u2_u14_u7_U21 (.A( u2_u14_u7_n101 ) , .ZN( u2_u14_u7_n165 ) );
  NOR2_X1 u2_u14_u7_U22 (.ZN( u2_u14_u7_n111 ) , .A2( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U23 (.A( u2_u14_u7_n138 ) , .ZN( u2_u14_u7_n171 ) );
  INV_X1 u2_u14_u7_U24 (.A( u2_u14_u7_n131 ) , .ZN( u2_u14_u7_n177 ) );
  INV_X1 u2_u14_u7_U25 (.A( u2_u14_u7_n110 ) , .ZN( u2_u14_u7_n174 ) );
  NAND2_X1 u2_u14_u7_U26 (.A1( u2_u14_u7_n129 ) , .A2( u2_u14_u7_n132 ) , .ZN( u2_u14_u7_n149 ) );
  NAND2_X1 u2_u14_u7_U27 (.A1( u2_u14_u7_n113 ) , .A2( u2_u14_u7_n124 ) , .ZN( u2_u14_u7_n130 ) );
  INV_X1 u2_u14_u7_U28 (.A( u2_u14_u7_n112 ) , .ZN( u2_u14_u7_n173 ) );
  INV_X1 u2_u14_u7_U29 (.A( u2_u14_u7_n128 ) , .ZN( u2_u14_u7_n168 ) );
  OAI21_X1 u2_u14_u7_U3 (.ZN( u2_u14_u7_n159 ) , .A( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n171 ) , .B1( u2_u14_u7_n174 ) );
  INV_X1 u2_u14_u7_U30 (.A( u2_u14_u7_n148 ) , .ZN( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U31 (.A( u2_u14_u7_n127 ) , .ZN( u2_u14_u7_n179 ) );
  NOR2_X1 u2_u14_u7_U32 (.ZN( u2_u14_u7_n101 ) , .A2( u2_u14_u7_n150 ) , .A1( u2_u14_u7_n156 ) );
  AOI211_X1 u2_u14_u7_U33 (.B( u2_u14_u7_n139 ) , .A( u2_u14_u7_n140 ) , .C2( u2_u14_u7_n141 ) , .ZN( u2_u14_u7_n142 ) , .C1( u2_u14_u7_n156 ) );
  NAND4_X1 u2_u14_u7_U34 (.A3( u2_u14_u7_n127 ) , .A2( u2_u14_u7_n128 ) , .A1( u2_u14_u7_n129 ) , .ZN( u2_u14_u7_n141 ) , .A4( u2_u14_u7_n147 ) );
  AOI21_X1 u2_u14_u7_U35 (.A( u2_u14_u7_n137 ) , .B1( u2_u14_u7_n138 ) , .ZN( u2_u14_u7_n139 ) , .B2( u2_u14_u7_n146 ) );
  OAI22_X1 u2_u14_u7_U36 (.B1( u2_u14_u7_n136 ) , .ZN( u2_u14_u7_n140 ) , .A1( u2_u14_u7_n153 ) , .B2( u2_u14_u7_n162 ) , .A2( u2_u14_u7_n164 ) );
  INV_X1 u2_u14_u7_U37 (.A( u2_u14_u7_n125 ) , .ZN( u2_u14_u7_n161 ) );
  AOI21_X1 u2_u14_u7_U38 (.ZN( u2_u14_u7_n123 ) , .B1( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n177 ) , .A( u2_u14_u7_n97 ) );
  AOI21_X1 u2_u14_u7_U39 (.B2( u2_u14_u7_n113 ) , .B1( u2_u14_u7_n124 ) , .A( u2_u14_u7_n125 ) , .ZN( u2_u14_u7_n97 ) );
  INV_X1 u2_u14_u7_U4 (.A( u2_u14_u7_n149 ) , .ZN( u2_u14_u7_n175 ) );
  INV_X1 u2_u14_u7_U40 (.A( u2_u14_u7_n152 ) , .ZN( u2_u14_u7_n162 ) );
  AOI22_X1 u2_u14_u7_U41 (.A2( u2_u14_u7_n114 ) , .ZN( u2_u14_u7_n119 ) , .B1( u2_u14_u7_n130 ) , .A1( u2_u14_u7_n156 ) , .B2( u2_u14_u7_n165 ) );
  NAND2_X1 u2_u14_u7_U42 (.A2( u2_u14_u7_n112 ) , .ZN( u2_u14_u7_n114 ) , .A1( u2_u14_u7_n175 ) );
  NOR2_X1 u2_u14_u7_U43 (.ZN( u2_u14_u7_n137 ) , .A1( u2_u14_u7_n150 ) , .A2( u2_u14_u7_n161 ) );
  AND2_X1 u2_u14_u7_U44 (.ZN( u2_u14_u7_n145 ) , .A2( u2_u14_u7_n98 ) , .A1( u2_u14_u7_n99 ) );
  AOI21_X1 u2_u14_u7_U45 (.ZN( u2_u14_u7_n105 ) , .B2( u2_u14_u7_n110 ) , .A( u2_u14_u7_n125 ) , .B1( u2_u14_u7_n147 ) );
  NAND2_X1 u2_u14_u7_U46 (.ZN( u2_u14_u7_n146 ) , .A1( u2_u14_u7_n95 ) , .A2( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U47 (.A2( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n147 ) , .A1( u2_u14_u7_n93 ) );
  NAND2_X1 u2_u14_u7_U48 (.A1( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n127 ) , .A2( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U49 (.A2( u2_u14_u7_n102 ) , .A1( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n133 ) );
  INV_X1 u2_u14_u7_U5 (.A( u2_u14_u7_n154 ) , .ZN( u2_u14_u7_n178 ) );
  OR2_X1 u2_u14_u7_U50 (.ZN( u2_u14_u7_n126 ) , .A2( u2_u14_u7_n152 ) , .A1( u2_u14_u7_n156 ) );
  NAND2_X1 u2_u14_u7_U51 (.ZN( u2_u14_u7_n112 ) , .A2( u2_u14_u7_n96 ) , .A1( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U52 (.A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n128 ) , .A1( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U53 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n113 ) , .A2( u2_u14_u7_n93 ) );
  NAND2_X1 u2_u14_u7_U54 (.ZN( u2_u14_u7_n110 ) , .A1( u2_u14_u7_n95 ) , .A2( u2_u14_u7_n96 ) );
  INV_X1 u2_u14_u7_U55 (.A( u2_u14_u7_n150 ) , .ZN( u2_u14_u7_n164 ) );
  AND2_X1 u2_u14_u7_U56 (.ZN( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n93 ) , .A2( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U57 (.A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n124 ) , .A1( u2_u14_u7_n96 ) );
  NAND2_X1 u2_u14_u7_U58 (.A1( u2_u14_u7_n100 ) , .A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n129 ) );
  NAND2_X1 u2_u14_u7_U59 (.A2( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n131 ) , .A1( u2_u14_u7_n95 ) );
  AOI211_X1 u2_u14_u7_U6 (.ZN( u2_u14_u7_n116 ) , .A( u2_u14_u7_n155 ) , .C1( u2_u14_u7_n161 ) , .C2( u2_u14_u7_n171 ) , .B( u2_u14_u7_n94 ) );
  NAND2_X1 u2_u14_u7_U60 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n138 ) , .A2( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U61 (.ZN( u2_u14_u7_n132 ) , .A1( u2_u14_u7_n93 ) , .A2( u2_u14_u7_n96 ) );
  NAND2_X1 u2_u14_u7_U62 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n148 ) , .A2( u2_u14_u7_n95 ) );
  AOI211_X1 u2_u14_u7_U63 (.B( u2_u14_u7_n154 ) , .A( u2_u14_u7_n155 ) , .C1( u2_u14_u7_n156 ) , .ZN( u2_u14_u7_n157 ) , .C2( u2_u14_u7_n172 ) );
  INV_X1 u2_u14_u7_U64 (.A( u2_u14_u7_n153 ) , .ZN( u2_u14_u7_n172 ) );
  NOR2_X1 u2_u14_u7_U65 (.A2( u2_u14_X_47 ) , .ZN( u2_u14_u7_n150 ) , .A1( u2_u14_u7_n163 ) );
  NOR2_X1 u2_u14_u7_U66 (.A2( u2_u14_X_43 ) , .A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n103 ) );
  NOR2_X1 u2_u14_u7_U67 (.A2( u2_u14_X_48 ) , .A1( u2_u14_u7_n166 ) , .ZN( u2_u14_u7_n95 ) );
  NOR2_X1 u2_u14_u7_U68 (.A2( u2_u14_X_45 ) , .A1( u2_u14_X_48 ) , .ZN( u2_u14_u7_n99 ) );
  NOR2_X1 u2_u14_u7_U69 (.A2( u2_u14_X_44 ) , .A1( u2_u14_u7_n167 ) , .ZN( u2_u14_u7_n98 ) );
  OAI222_X1 u2_u14_u7_U7 (.C2( u2_u14_u7_n101 ) , .B2( u2_u14_u7_n111 ) , .A1( u2_u14_u7_n113 ) , .C1( u2_u14_u7_n146 ) , .A2( u2_u14_u7_n162 ) , .B1( u2_u14_u7_n164 ) , .ZN( u2_u14_u7_n94 ) );
  NOR2_X1 u2_u14_u7_U70 (.A2( u2_u14_X_46 ) , .A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n152 ) );
  NAND2_X1 u2_u14_u7_U71 (.A2( u2_u14_X_46 ) , .A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n125 ) );
  AND2_X1 u2_u14_u7_U72 (.A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n156 ) , .A2( u2_u14_u7_n163 ) );
  AND2_X1 u2_u14_u7_U73 (.A2( u2_u14_X_45 ) , .A1( u2_u14_X_48 ) , .ZN( u2_u14_u7_n102 ) );
  AND2_X1 u2_u14_u7_U74 (.A2( u2_u14_X_43 ) , .A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n96 ) );
  AND2_X1 u2_u14_u7_U75 (.A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n100 ) , .A2( u2_u14_u7_n167 ) );
  AND2_X1 u2_u14_u7_U76 (.A1( u2_u14_X_48 ) , .A2( u2_u14_u7_n166 ) , .ZN( u2_u14_u7_n93 ) );
  INV_X1 u2_u14_u7_U77 (.A( u2_u14_X_46 ) , .ZN( u2_u14_u7_n163 ) );
  INV_X1 u2_u14_u7_U78 (.A( u2_u14_X_45 ) , .ZN( u2_u14_u7_n166 ) );
  INV_X1 u2_u14_u7_U79 (.A( u2_u14_X_43 ) , .ZN( u2_u14_u7_n167 ) );
  OAI221_X1 u2_u14_u7_U8 (.C1( u2_u14_u7_n101 ) , .C2( u2_u14_u7_n147 ) , .ZN( u2_u14_u7_n155 ) , .B2( u2_u14_u7_n162 ) , .A( u2_u14_u7_n91 ) , .B1( u2_u14_u7_n92 ) );
  NAND4_X1 u2_u14_u7_U80 (.ZN( u2_out14_27 ) , .A4( u2_u14_u7_n118 ) , .A3( u2_u14_u7_n119 ) , .A2( u2_u14_u7_n120 ) , .A1( u2_u14_u7_n121 ) );
  OAI21_X1 u2_u14_u7_U81 (.ZN( u2_u14_u7_n121 ) , .B2( u2_u14_u7_n145 ) , .A( u2_u14_u7_n150 ) , .B1( u2_u14_u7_n174 ) );
  OAI21_X1 u2_u14_u7_U82 (.ZN( u2_u14_u7_n120 ) , .A( u2_u14_u7_n161 ) , .B2( u2_u14_u7_n170 ) , .B1( u2_u14_u7_n179 ) );
  NAND4_X1 u2_u14_u7_U83 (.ZN( u2_out14_21 ) , .A4( u2_u14_u7_n157 ) , .A3( u2_u14_u7_n158 ) , .A2( u2_u14_u7_n159 ) , .A1( u2_u14_u7_n160 ) );
  OAI21_X1 u2_u14_u7_U84 (.B1( u2_u14_u7_n145 ) , .ZN( u2_u14_u7_n160 ) , .A( u2_u14_u7_n161 ) , .B2( u2_u14_u7_n177 ) );
  AOI22_X1 u2_u14_u7_U85 (.B2( u2_u14_u7_n149 ) , .B1( u2_u14_u7_n150 ) , .A2( u2_u14_u7_n151 ) , .A1( u2_u14_u7_n152 ) , .ZN( u2_u14_u7_n158 ) );
  NAND4_X1 u2_u14_u7_U86 (.ZN( u2_out14_15 ) , .A4( u2_u14_u7_n142 ) , .A3( u2_u14_u7_n143 ) , .A2( u2_u14_u7_n144 ) , .A1( u2_u14_u7_n178 ) );
  OR2_X1 u2_u14_u7_U87 (.A2( u2_u14_u7_n125 ) , .A1( u2_u14_u7_n129 ) , .ZN( u2_u14_u7_n144 ) );
  AOI22_X1 u2_u14_u7_U88 (.A2( u2_u14_u7_n126 ) , .ZN( u2_u14_u7_n143 ) , .B2( u2_u14_u7_n165 ) , .B1( u2_u14_u7_n173 ) , .A1( u2_u14_u7_n174 ) );
  NAND4_X1 u2_u14_u7_U89 (.ZN( u2_out14_5 ) , .A4( u2_u14_u7_n108 ) , .A3( u2_u14_u7_n109 ) , .A1( u2_u14_u7_n116 ) , .A2( u2_u14_u7_n123 ) );
  AND3_X1 u2_u14_u7_U9 (.A3( u2_u14_u7_n110 ) , .A2( u2_u14_u7_n127 ) , .A1( u2_u14_u7_n132 ) , .ZN( u2_u14_u7_n92 ) );
  AOI22_X1 u2_u14_u7_U90 (.ZN( u2_u14_u7_n109 ) , .A2( u2_u14_u7_n126 ) , .B2( u2_u14_u7_n145 ) , .B1( u2_u14_u7_n156 ) , .A1( u2_u14_u7_n171 ) );
  NOR4_X1 u2_u14_u7_U91 (.A4( u2_u14_u7_n104 ) , .A3( u2_u14_u7_n105 ) , .A2( u2_u14_u7_n106 ) , .A1( u2_u14_u7_n107 ) , .ZN( u2_u14_u7_n108 ) );
  OAI211_X1 u2_u14_u7_U92 (.B( u2_u14_u7_n122 ) , .A( u2_u14_u7_n123 ) , .C2( u2_u14_u7_n124 ) , .ZN( u2_u14_u7_n154 ) , .C1( u2_u14_u7_n162 ) );
  AOI222_X1 u2_u14_u7_U93 (.ZN( u2_u14_u7_n122 ) , .C2( u2_u14_u7_n126 ) , .C1( u2_u14_u7_n145 ) , .B1( u2_u14_u7_n161 ) , .A2( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n170 ) , .A1( u2_u14_u7_n176 ) );
  INV_X1 u2_u14_u7_U94 (.A( u2_u14_u7_n111 ) , .ZN( u2_u14_u7_n170 ) );
  NAND3_X1 u2_u14_u7_U95 (.A3( u2_u14_u7_n146 ) , .A2( u2_u14_u7_n147 ) , .A1( u2_u14_u7_n148 ) , .ZN( u2_u14_u7_n151 ) );
  NAND3_X1 u2_u14_u7_U96 (.A3( u2_u14_u7_n131 ) , .A2( u2_u14_u7_n132 ) , .A1( u2_u14_u7_n133 ) , .ZN( u2_u14_u7_n135 ) );
  XOR2_X1 u2_u2_U1 (.B( u2_K3_9 ) , .A( u2_R1_6 ) , .Z( u2_u2_X_9 ) );
  XOR2_X1 u2_u2_U2 (.B( u2_K3_8 ) , .A( u2_R1_5 ) , .Z( u2_u2_X_8 ) );
  XOR2_X1 u2_u2_U3 (.B( u2_K3_7 ) , .A( u2_R1_4 ) , .Z( u2_u2_X_7 ) );
  XOR2_X1 u2_u2_U46 (.B( u2_K3_12 ) , .A( u2_R1_9 ) , .Z( u2_u2_X_12 ) );
  XOR2_X1 u2_u2_U47 (.B( u2_K3_11 ) , .A( u2_R1_8 ) , .Z( u2_u2_X_11 ) );
  XOR2_X1 u2_u2_U48 (.B( u2_K3_10 ) , .A( u2_R1_7 ) , .Z( u2_u2_X_10 ) );
  NOR2_X1 u2_u2_u1_U10 (.A1( u2_u2_u1_n112 ) , .A2( u2_u2_u1_n116 ) , .ZN( u2_u2_u1_n118 ) );
  NAND3_X1 u2_u2_u1_U100 (.ZN( u2_u2_u1_n113 ) , .A1( u2_u2_u1_n120 ) , .A3( u2_u2_u1_n133 ) , .A2( u2_u2_u1_n155 ) );
  OAI21_X1 u2_u2_u1_U11 (.ZN( u2_u2_u1_n101 ) , .B1( u2_u2_u1_n141 ) , .A( u2_u2_u1_n146 ) , .B2( u2_u2_u1_n183 ) );
  AOI21_X1 u2_u2_u1_U12 (.B2( u2_u2_u1_n155 ) , .B1( u2_u2_u1_n156 ) , .ZN( u2_u2_u1_n157 ) , .A( u2_u2_u1_n174 ) );
  OR4_X1 u2_u2_u1_U13 (.A4( u2_u2_u1_n106 ) , .A3( u2_u2_u1_n107 ) , .ZN( u2_u2_u1_n108 ) , .A1( u2_u2_u1_n117 ) , .A2( u2_u2_u1_n184 ) );
  AOI21_X1 u2_u2_u1_U14 (.ZN( u2_u2_u1_n106 ) , .A( u2_u2_u1_n112 ) , .B1( u2_u2_u1_n154 ) , .B2( u2_u2_u1_n156 ) );
  INV_X1 u2_u2_u1_U15 (.A( u2_u2_u1_n101 ) , .ZN( u2_u2_u1_n184 ) );
  AOI21_X1 u2_u2_u1_U16 (.ZN( u2_u2_u1_n107 ) , .B1( u2_u2_u1_n134 ) , .B2( u2_u2_u1_n149 ) , .A( u2_u2_u1_n174 ) );
  NAND2_X1 u2_u2_u1_U17 (.ZN( u2_u2_u1_n140 ) , .A2( u2_u2_u1_n150 ) , .A1( u2_u2_u1_n155 ) );
  NAND2_X1 u2_u2_u1_U18 (.A1( u2_u2_u1_n131 ) , .ZN( u2_u2_u1_n147 ) , .A2( u2_u2_u1_n153 ) );
  INV_X1 u2_u2_u1_U19 (.A( u2_u2_u1_n139 ) , .ZN( u2_u2_u1_n174 ) );
  INV_X1 u2_u2_u1_U20 (.A( u2_u2_u1_n112 ) , .ZN( u2_u2_u1_n171 ) );
  NAND2_X1 u2_u2_u1_U21 (.ZN( u2_u2_u1_n141 ) , .A1( u2_u2_u1_n153 ) , .A2( u2_u2_u1_n156 ) );
  AND2_X1 u2_u2_u1_U22 (.A1( u2_u2_u1_n123 ) , .ZN( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n161 ) );
  NAND2_X1 u2_u2_u1_U23 (.A2( u2_u2_u1_n115 ) , .A1( u2_u2_u1_n116 ) , .ZN( u2_u2_u1_n148 ) );
  NAND2_X1 u2_u2_u1_U24 (.A2( u2_u2_u1_n133 ) , .A1( u2_u2_u1_n135 ) , .ZN( u2_u2_u1_n159 ) );
  NAND2_X1 u2_u2_u1_U25 (.A2( u2_u2_u1_n115 ) , .A1( u2_u2_u1_n120 ) , .ZN( u2_u2_u1_n132 ) );
  INV_X1 u2_u2_u1_U26 (.A( u2_u2_u1_n154 ) , .ZN( u2_u2_u1_n178 ) );
  INV_X1 u2_u2_u1_U27 (.A( u2_u2_u1_n151 ) , .ZN( u2_u2_u1_n183 ) );
  AND2_X1 u2_u2_u1_U28 (.A1( u2_u2_u1_n129 ) , .A2( u2_u2_u1_n133 ) , .ZN( u2_u2_u1_n149 ) );
  INV_X1 u2_u2_u1_U29 (.A( u2_u2_u1_n131 ) , .ZN( u2_u2_u1_n180 ) );
  INV_X1 u2_u2_u1_U3 (.A( u2_u2_u1_n159 ) , .ZN( u2_u2_u1_n182 ) );
  OAI221_X1 u2_u2_u1_U30 (.A( u2_u2_u1_n119 ) , .C2( u2_u2_u1_n129 ) , .ZN( u2_u2_u1_n138 ) , .B2( u2_u2_u1_n152 ) , .C1( u2_u2_u1_n174 ) , .B1( u2_u2_u1_n187 ) );
  INV_X1 u2_u2_u1_U31 (.A( u2_u2_u1_n148 ) , .ZN( u2_u2_u1_n187 ) );
  AOI211_X1 u2_u2_u1_U32 (.B( u2_u2_u1_n117 ) , .A( u2_u2_u1_n118 ) , .ZN( u2_u2_u1_n119 ) , .C2( u2_u2_u1_n146 ) , .C1( u2_u2_u1_n159 ) );
  NOR2_X1 u2_u2_u1_U33 (.A1( u2_u2_u1_n168 ) , .A2( u2_u2_u1_n176 ) , .ZN( u2_u2_u1_n98 ) );
  AOI211_X1 u2_u2_u1_U34 (.B( u2_u2_u1_n162 ) , .A( u2_u2_u1_n163 ) , .C2( u2_u2_u1_n164 ) , .ZN( u2_u2_u1_n165 ) , .C1( u2_u2_u1_n171 ) );
  AOI21_X1 u2_u2_u1_U35 (.A( u2_u2_u1_n160 ) , .B2( u2_u2_u1_n161 ) , .ZN( u2_u2_u1_n162 ) , .B1( u2_u2_u1_n182 ) );
  OR2_X1 u2_u2_u1_U36 (.A2( u2_u2_u1_n157 ) , .A1( u2_u2_u1_n158 ) , .ZN( u2_u2_u1_n163 ) );
  OAI21_X1 u2_u2_u1_U37 (.B2( u2_u2_u1_n123 ) , .ZN( u2_u2_u1_n145 ) , .B1( u2_u2_u1_n160 ) , .A( u2_u2_u1_n185 ) );
  INV_X1 u2_u2_u1_U38 (.A( u2_u2_u1_n122 ) , .ZN( u2_u2_u1_n185 ) );
  AOI21_X1 u2_u2_u1_U39 (.B2( u2_u2_u1_n120 ) , .B1( u2_u2_u1_n121 ) , .ZN( u2_u2_u1_n122 ) , .A( u2_u2_u1_n128 ) );
  AOI221_X1 u2_u2_u1_U4 (.A( u2_u2_u1_n138 ) , .C2( u2_u2_u1_n139 ) , .C1( u2_u2_u1_n140 ) , .B2( u2_u2_u1_n141 ) , .ZN( u2_u2_u1_n142 ) , .B1( u2_u2_u1_n175 ) );
  NAND2_X1 u2_u2_u1_U40 (.A1( u2_u2_u1_n128 ) , .ZN( u2_u2_u1_n146 ) , .A2( u2_u2_u1_n160 ) );
  NAND2_X1 u2_u2_u1_U41 (.A2( u2_u2_u1_n112 ) , .ZN( u2_u2_u1_n139 ) , .A1( u2_u2_u1_n152 ) );
  NAND2_X1 u2_u2_u1_U42 (.A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n156 ) , .A2( u2_u2_u1_n99 ) );
  AOI221_X1 u2_u2_u1_U43 (.B1( u2_u2_u1_n140 ) , .ZN( u2_u2_u1_n167 ) , .B2( u2_u2_u1_n172 ) , .C2( u2_u2_u1_n175 ) , .C1( u2_u2_u1_n178 ) , .A( u2_u2_u1_n188 ) );
  INV_X1 u2_u2_u1_U44 (.ZN( u2_u2_u1_n188 ) , .A( u2_u2_u1_n97 ) );
  AOI211_X1 u2_u2_u1_U45 (.A( u2_u2_u1_n118 ) , .C1( u2_u2_u1_n132 ) , .C2( u2_u2_u1_n139 ) , .B( u2_u2_u1_n96 ) , .ZN( u2_u2_u1_n97 ) );
  AOI21_X1 u2_u2_u1_U46 (.B2( u2_u2_u1_n121 ) , .B1( u2_u2_u1_n135 ) , .A( u2_u2_u1_n152 ) , .ZN( u2_u2_u1_n96 ) );
  NOR2_X1 u2_u2_u1_U47 (.ZN( u2_u2_u1_n117 ) , .A1( u2_u2_u1_n121 ) , .A2( u2_u2_u1_n160 ) );
  AOI21_X1 u2_u2_u1_U48 (.A( u2_u2_u1_n128 ) , .B2( u2_u2_u1_n129 ) , .ZN( u2_u2_u1_n130 ) , .B1( u2_u2_u1_n150 ) );
  NAND2_X1 u2_u2_u1_U49 (.ZN( u2_u2_u1_n112 ) , .A1( u2_u2_u1_n169 ) , .A2( u2_u2_u1_n170 ) );
  AOI211_X1 u2_u2_u1_U5 (.ZN( u2_u2_u1_n124 ) , .A( u2_u2_u1_n138 ) , .C2( u2_u2_u1_n139 ) , .B( u2_u2_u1_n145 ) , .C1( u2_u2_u1_n147 ) );
  NAND2_X1 u2_u2_u1_U50 (.ZN( u2_u2_u1_n129 ) , .A2( u2_u2_u1_n95 ) , .A1( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U51 (.A1( u2_u2_u1_n102 ) , .ZN( u2_u2_u1_n154 ) , .A2( u2_u2_u1_n99 ) );
  NAND2_X1 u2_u2_u1_U52 (.A2( u2_u2_u1_n100 ) , .ZN( u2_u2_u1_n135 ) , .A1( u2_u2_u1_n99 ) );
  AOI21_X1 u2_u2_u1_U53 (.A( u2_u2_u1_n152 ) , .B2( u2_u2_u1_n153 ) , .B1( u2_u2_u1_n154 ) , .ZN( u2_u2_u1_n158 ) );
  INV_X1 u2_u2_u1_U54 (.A( u2_u2_u1_n160 ) , .ZN( u2_u2_u1_n175 ) );
  NAND2_X1 u2_u2_u1_U55 (.A1( u2_u2_u1_n100 ) , .ZN( u2_u2_u1_n116 ) , .A2( u2_u2_u1_n95 ) );
  NAND2_X1 u2_u2_u1_U56 (.A1( u2_u2_u1_n102 ) , .ZN( u2_u2_u1_n131 ) , .A2( u2_u2_u1_n95 ) );
  NAND2_X1 u2_u2_u1_U57 (.A2( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n121 ) , .A1( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U58 (.A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n153 ) , .A2( u2_u2_u1_n98 ) );
  NAND2_X1 u2_u2_u1_U59 (.A2( u2_u2_u1_n104 ) , .A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n133 ) );
  AOI22_X1 u2_u2_u1_U6 (.B2( u2_u2_u1_n113 ) , .A2( u2_u2_u1_n114 ) , .ZN( u2_u2_u1_n125 ) , .A1( u2_u2_u1_n171 ) , .B1( u2_u2_u1_n173 ) );
  NAND2_X1 u2_u2_u1_U60 (.ZN( u2_u2_u1_n150 ) , .A2( u2_u2_u1_n98 ) , .A1( u2_u2_u1_n99 ) );
  NAND2_X1 u2_u2_u1_U61 (.A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n155 ) , .A2( u2_u2_u1_n95 ) );
  OAI21_X1 u2_u2_u1_U62 (.ZN( u2_u2_u1_n109 ) , .B1( u2_u2_u1_n129 ) , .B2( u2_u2_u1_n160 ) , .A( u2_u2_u1_n167 ) );
  NAND2_X1 u2_u2_u1_U63 (.A2( u2_u2_u1_n100 ) , .A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n120 ) );
  NAND2_X1 u2_u2_u1_U64 (.A1( u2_u2_u1_n102 ) , .A2( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n115 ) );
  NAND2_X1 u2_u2_u1_U65 (.A2( u2_u2_u1_n100 ) , .A1( u2_u2_u1_n104 ) , .ZN( u2_u2_u1_n151 ) );
  NAND2_X1 u2_u2_u1_U66 (.A2( u2_u2_u1_n103 ) , .A1( u2_u2_u1_n105 ) , .ZN( u2_u2_u1_n161 ) );
  INV_X1 u2_u2_u1_U67 (.A( u2_u2_u1_n152 ) , .ZN( u2_u2_u1_n173 ) );
  INV_X1 u2_u2_u1_U68 (.A( u2_u2_u1_n128 ) , .ZN( u2_u2_u1_n172 ) );
  NAND2_X1 u2_u2_u1_U69 (.A2( u2_u2_u1_n102 ) , .A1( u2_u2_u1_n103 ) , .ZN( u2_u2_u1_n123 ) );
  NAND2_X1 u2_u2_u1_U7 (.ZN( u2_u2_u1_n114 ) , .A1( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n156 ) );
  NOR2_X1 u2_u2_u1_U70 (.A2( u2_u2_X_7 ) , .A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n95 ) );
  NOR2_X1 u2_u2_u1_U71 (.A1( u2_u2_X_12 ) , .A2( u2_u2_X_9 ) , .ZN( u2_u2_u1_n100 ) );
  NOR2_X1 u2_u2_u1_U72 (.A2( u2_u2_X_8 ) , .A1( u2_u2_u1_n177 ) , .ZN( u2_u2_u1_n99 ) );
  NOR2_X1 u2_u2_u1_U73 (.A2( u2_u2_X_12 ) , .ZN( u2_u2_u1_n102 ) , .A1( u2_u2_u1_n176 ) );
  NOR2_X1 u2_u2_u1_U74 (.A2( u2_u2_X_9 ) , .ZN( u2_u2_u1_n105 ) , .A1( u2_u2_u1_n168 ) );
  NAND2_X1 u2_u2_u1_U75 (.A1( u2_u2_X_10 ) , .ZN( u2_u2_u1_n160 ) , .A2( u2_u2_u1_n169 ) );
  NAND2_X1 u2_u2_u1_U76 (.A2( u2_u2_X_10 ) , .A1( u2_u2_X_11 ) , .ZN( u2_u2_u1_n152 ) );
  NAND2_X1 u2_u2_u1_U77 (.A1( u2_u2_X_11 ) , .ZN( u2_u2_u1_n128 ) , .A2( u2_u2_u1_n170 ) );
  AND2_X1 u2_u2_u1_U78 (.A2( u2_u2_X_7 ) , .A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n104 ) );
  AND2_X1 u2_u2_u1_U79 (.A1( u2_u2_X_8 ) , .ZN( u2_u2_u1_n103 ) , .A2( u2_u2_u1_n177 ) );
  AOI22_X1 u2_u2_u1_U8 (.B2( u2_u2_u1_n136 ) , .A2( u2_u2_u1_n137 ) , .ZN( u2_u2_u1_n143 ) , .A1( u2_u2_u1_n171 ) , .B1( u2_u2_u1_n173 ) );
  INV_X1 u2_u2_u1_U80 (.A( u2_u2_X_10 ) , .ZN( u2_u2_u1_n170 ) );
  INV_X1 u2_u2_u1_U81 (.A( u2_u2_X_9 ) , .ZN( u2_u2_u1_n176 ) );
  INV_X1 u2_u2_u1_U82 (.A( u2_u2_X_11 ) , .ZN( u2_u2_u1_n169 ) );
  INV_X1 u2_u2_u1_U83 (.A( u2_u2_X_12 ) , .ZN( u2_u2_u1_n168 ) );
  INV_X1 u2_u2_u1_U84 (.A( u2_u2_X_7 ) , .ZN( u2_u2_u1_n177 ) );
  NAND4_X1 u2_u2_u1_U85 (.ZN( u2_out2_28 ) , .A4( u2_u2_u1_n124 ) , .A3( u2_u2_u1_n125 ) , .A2( u2_u2_u1_n126 ) , .A1( u2_u2_u1_n127 ) );
  OAI21_X1 u2_u2_u1_U86 (.ZN( u2_u2_u1_n127 ) , .B2( u2_u2_u1_n139 ) , .B1( u2_u2_u1_n175 ) , .A( u2_u2_u1_n183 ) );
  OAI21_X1 u2_u2_u1_U87 (.ZN( u2_u2_u1_n126 ) , .B2( u2_u2_u1_n140 ) , .A( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n178 ) );
  NAND4_X1 u2_u2_u1_U88 (.ZN( u2_out2_18 ) , .A4( u2_u2_u1_n165 ) , .A3( u2_u2_u1_n166 ) , .A1( u2_u2_u1_n167 ) , .A2( u2_u2_u1_n186 ) );
  AOI22_X1 u2_u2_u1_U89 (.B2( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n147 ) , .A2( u2_u2_u1_n148 ) , .ZN( u2_u2_u1_n166 ) , .A1( u2_u2_u1_n172 ) );
  INV_X1 u2_u2_u1_U9 (.A( u2_u2_u1_n147 ) , .ZN( u2_u2_u1_n181 ) );
  INV_X1 u2_u2_u1_U90 (.A( u2_u2_u1_n145 ) , .ZN( u2_u2_u1_n186 ) );
  NAND4_X1 u2_u2_u1_U91 (.ZN( u2_out2_2 ) , .A4( u2_u2_u1_n142 ) , .A3( u2_u2_u1_n143 ) , .A2( u2_u2_u1_n144 ) , .A1( u2_u2_u1_n179 ) );
  OAI21_X1 u2_u2_u1_U92 (.B2( u2_u2_u1_n132 ) , .ZN( u2_u2_u1_n144 ) , .A( u2_u2_u1_n146 ) , .B1( u2_u2_u1_n180 ) );
  INV_X1 u2_u2_u1_U93 (.A( u2_u2_u1_n130 ) , .ZN( u2_u2_u1_n179 ) );
  OR4_X1 u2_u2_u1_U94 (.ZN( u2_out2_13 ) , .A4( u2_u2_u1_n108 ) , .A3( u2_u2_u1_n109 ) , .A2( u2_u2_u1_n110 ) , .A1( u2_u2_u1_n111 ) );
  AOI21_X1 u2_u2_u1_U95 (.ZN( u2_u2_u1_n111 ) , .A( u2_u2_u1_n128 ) , .B2( u2_u2_u1_n131 ) , .B1( u2_u2_u1_n135 ) );
  AOI21_X1 u2_u2_u1_U96 (.ZN( u2_u2_u1_n110 ) , .A( u2_u2_u1_n116 ) , .B1( u2_u2_u1_n152 ) , .B2( u2_u2_u1_n160 ) );
  NAND3_X1 u2_u2_u1_U97 (.A3( u2_u2_u1_n149 ) , .A2( u2_u2_u1_n150 ) , .A1( u2_u2_u1_n151 ) , .ZN( u2_u2_u1_n164 ) );
  NAND3_X1 u2_u2_u1_U98 (.A3( u2_u2_u1_n134 ) , .A2( u2_u2_u1_n135 ) , .ZN( u2_u2_u1_n136 ) , .A1( u2_u2_u1_n151 ) );
  NAND3_X1 u2_u2_u1_U99 (.A1( u2_u2_u1_n133 ) , .ZN( u2_u2_u1_n137 ) , .A2( u2_u2_u1_n154 ) , .A3( u2_u2_u1_n181 ) );
  XOR2_X1 u2_u3_U33 (.B( u2_K4_24 ) , .A( u2_R2_17 ) , .Z( u2_u3_X_24 ) );
  XOR2_X1 u2_u3_U34 (.B( u2_K4_23 ) , .A( u2_R2_16 ) , .Z( u2_u3_X_23 ) );
  XOR2_X1 u2_u3_U35 (.B( u2_K4_22 ) , .A( u2_R2_15 ) , .Z( u2_u3_X_22 ) );
  XOR2_X1 u2_u3_U36 (.B( u2_K4_21 ) , .A( u2_R2_14 ) , .Z( u2_u3_X_21 ) );
  XOR2_X1 u2_u3_U37 (.B( u2_K4_20 ) , .A( u2_R2_13 ) , .Z( u2_u3_X_20 ) );
  XOR2_X1 u2_u3_U39 (.B( u2_K4_19 ) , .A( u2_R2_12 ) , .Z( u2_u3_X_19 ) );
  XOR2_X1 u2_u3_U40 (.B( u2_K4_18 ) , .A( u2_R2_13 ) , .Z( u2_u3_X_18 ) );
  XOR2_X1 u2_u3_U41 (.B( u2_K4_17 ) , .A( u2_R2_12 ) , .Z( u2_u3_X_17 ) );
  XOR2_X1 u2_u3_U42 (.B( u2_K4_16 ) , .A( u2_R2_11 ) , .Z( u2_u3_X_16 ) );
  XOR2_X1 u2_u3_U43 (.B( u2_K4_15 ) , .A( u2_R2_10 ) , .Z( u2_u3_X_15 ) );
  XOR2_X1 u2_u3_U44 (.B( u2_K4_14 ) , .A( u2_R2_9 ) , .Z( u2_u3_X_14 ) );
  XOR2_X1 u2_u3_U45 (.B( u2_K4_13 ) , .A( u2_R2_8 ) , .Z( u2_u3_X_13 ) );
  OAI22_X1 u2_u3_u2_U10 (.B1( u2_u3_u2_n151 ) , .A2( u2_u3_u2_n152 ) , .A1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n160 ) , .B2( u2_u3_u2_n168 ) );
  NAND3_X1 u2_u3_u2_U100 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n98 ) );
  NOR3_X1 u2_u3_u2_U11 (.A1( u2_u3_u2_n150 ) , .ZN( u2_u3_u2_n151 ) , .A3( u2_u3_u2_n175 ) , .A2( u2_u3_u2_n188 ) );
  AOI21_X1 u2_u3_u2_U12 (.B2( u2_u3_u2_n123 ) , .ZN( u2_u3_u2_n125 ) , .A( u2_u3_u2_n171 ) , .B1( u2_u3_u2_n184 ) );
  INV_X1 u2_u3_u2_U13 (.A( u2_u3_u2_n150 ) , .ZN( u2_u3_u2_n184 ) );
  AOI21_X1 u2_u3_u2_U14 (.ZN( u2_u3_u2_n144 ) , .B2( u2_u3_u2_n155 ) , .A( u2_u3_u2_n172 ) , .B1( u2_u3_u2_n185 ) );
  AOI21_X1 u2_u3_u2_U15 (.B2( u2_u3_u2_n143 ) , .ZN( u2_u3_u2_n145 ) , .B1( u2_u3_u2_n152 ) , .A( u2_u3_u2_n171 ) );
  INV_X1 u2_u3_u2_U16 (.A( u2_u3_u2_n156 ) , .ZN( u2_u3_u2_n171 ) );
  INV_X1 u2_u3_u2_U17 (.A( u2_u3_u2_n120 ) , .ZN( u2_u3_u2_n188 ) );
  NAND2_X1 u2_u3_u2_U18 (.A2( u2_u3_u2_n122 ) , .ZN( u2_u3_u2_n150 ) , .A1( u2_u3_u2_n152 ) );
  INV_X1 u2_u3_u2_U19 (.A( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n170 ) );
  INV_X1 u2_u3_u2_U20 (.A( u2_u3_u2_n137 ) , .ZN( u2_u3_u2_n173 ) );
  NAND2_X1 u2_u3_u2_U21 (.A1( u2_u3_u2_n132 ) , .A2( u2_u3_u2_n139 ) , .ZN( u2_u3_u2_n157 ) );
  INV_X1 u2_u3_u2_U22 (.A( u2_u3_u2_n113 ) , .ZN( u2_u3_u2_n178 ) );
  INV_X1 u2_u3_u2_U23 (.A( u2_u3_u2_n139 ) , .ZN( u2_u3_u2_n175 ) );
  INV_X1 u2_u3_u2_U24 (.A( u2_u3_u2_n155 ) , .ZN( u2_u3_u2_n181 ) );
  INV_X1 u2_u3_u2_U25 (.A( u2_u3_u2_n119 ) , .ZN( u2_u3_u2_n177 ) );
  INV_X1 u2_u3_u2_U26 (.A( u2_u3_u2_n116 ) , .ZN( u2_u3_u2_n180 ) );
  INV_X1 u2_u3_u2_U27 (.A( u2_u3_u2_n131 ) , .ZN( u2_u3_u2_n179 ) );
  INV_X1 u2_u3_u2_U28 (.A( u2_u3_u2_n154 ) , .ZN( u2_u3_u2_n176 ) );
  NAND2_X1 u2_u3_u2_U29 (.A2( u2_u3_u2_n116 ) , .A1( u2_u3_u2_n117 ) , .ZN( u2_u3_u2_n118 ) );
  NOR2_X1 u2_u3_u2_U3 (.ZN( u2_u3_u2_n121 ) , .A2( u2_u3_u2_n177 ) , .A1( u2_u3_u2_n180 ) );
  INV_X1 u2_u3_u2_U30 (.A( u2_u3_u2_n132 ) , .ZN( u2_u3_u2_n182 ) );
  INV_X1 u2_u3_u2_U31 (.A( u2_u3_u2_n158 ) , .ZN( u2_u3_u2_n183 ) );
  OAI21_X1 u2_u3_u2_U32 (.A( u2_u3_u2_n156 ) , .B1( u2_u3_u2_n157 ) , .ZN( u2_u3_u2_n158 ) , .B2( u2_u3_u2_n179 ) );
  NOR2_X1 u2_u3_u2_U33 (.ZN( u2_u3_u2_n156 ) , .A1( u2_u3_u2_n166 ) , .A2( u2_u3_u2_n169 ) );
  NOR2_X1 u2_u3_u2_U34 (.A2( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n137 ) , .A1( u2_u3_u2_n140 ) );
  NOR2_X1 u2_u3_u2_U35 (.A2( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n153 ) , .A1( u2_u3_u2_n156 ) );
  AOI211_X1 u2_u3_u2_U36 (.ZN( u2_u3_u2_n130 ) , .C1( u2_u3_u2_n138 ) , .C2( u2_u3_u2_n179 ) , .B( u2_u3_u2_n96 ) , .A( u2_u3_u2_n97 ) );
  OAI22_X1 u2_u3_u2_U37 (.B1( u2_u3_u2_n133 ) , .A2( u2_u3_u2_n137 ) , .A1( u2_u3_u2_n152 ) , .B2( u2_u3_u2_n168 ) , .ZN( u2_u3_u2_n97 ) );
  OAI221_X1 u2_u3_u2_U38 (.B1( u2_u3_u2_n113 ) , .C1( u2_u3_u2_n132 ) , .A( u2_u3_u2_n149 ) , .B2( u2_u3_u2_n171 ) , .C2( u2_u3_u2_n172 ) , .ZN( u2_u3_u2_n96 ) );
  OAI221_X1 u2_u3_u2_U39 (.A( u2_u3_u2_n115 ) , .C2( u2_u3_u2_n123 ) , .B2( u2_u3_u2_n143 ) , .B1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n163 ) , .C1( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U4 (.A( u2_u3_u2_n134 ) , .ZN( u2_u3_u2_n185 ) );
  OAI21_X1 u2_u3_u2_U40 (.A( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n115 ) , .B1( u2_u3_u2_n176 ) , .B2( u2_u3_u2_n178 ) );
  OAI221_X1 u2_u3_u2_U41 (.A( u2_u3_u2_n135 ) , .B2( u2_u3_u2_n136 ) , .B1( u2_u3_u2_n137 ) , .ZN( u2_u3_u2_n162 ) , .C2( u2_u3_u2_n167 ) , .C1( u2_u3_u2_n185 ) );
  AND3_X1 u2_u3_u2_U42 (.A3( u2_u3_u2_n131 ) , .A2( u2_u3_u2_n132 ) , .A1( u2_u3_u2_n133 ) , .ZN( u2_u3_u2_n136 ) );
  AOI22_X1 u2_u3_u2_U43 (.ZN( u2_u3_u2_n135 ) , .B1( u2_u3_u2_n140 ) , .A1( u2_u3_u2_n156 ) , .B2( u2_u3_u2_n180 ) , .A2( u2_u3_u2_n188 ) );
  AOI21_X1 u2_u3_u2_U44 (.ZN( u2_u3_u2_n149 ) , .B1( u2_u3_u2_n173 ) , .B2( u2_u3_u2_n188 ) , .A( u2_u3_u2_n95 ) );
  AND3_X1 u2_u3_u2_U45 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n156 ) , .ZN( u2_u3_u2_n95 ) );
  OAI21_X1 u2_u3_u2_U46 (.A( u2_u3_u2_n141 ) , .B2( u2_u3_u2_n142 ) , .ZN( u2_u3_u2_n146 ) , .B1( u2_u3_u2_n153 ) );
  OAI21_X1 u2_u3_u2_U47 (.A( u2_u3_u2_n140 ) , .ZN( u2_u3_u2_n141 ) , .B1( u2_u3_u2_n176 ) , .B2( u2_u3_u2_n177 ) );
  NOR3_X1 u2_u3_u2_U48 (.ZN( u2_u3_u2_n142 ) , .A3( u2_u3_u2_n175 ) , .A2( u2_u3_u2_n178 ) , .A1( u2_u3_u2_n181 ) );
  OAI21_X1 u2_u3_u2_U49 (.A( u2_u3_u2_n101 ) , .B2( u2_u3_u2_n121 ) , .B1( u2_u3_u2_n153 ) , .ZN( u2_u3_u2_n164 ) );
  NOR4_X1 u2_u3_u2_U5 (.A4( u2_u3_u2_n124 ) , .A3( u2_u3_u2_n125 ) , .A2( u2_u3_u2_n126 ) , .A1( u2_u3_u2_n127 ) , .ZN( u2_u3_u2_n128 ) );
  NAND2_X1 u2_u3_u2_U50 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n155 ) );
  NAND2_X1 u2_u3_u2_U51 (.A2( u2_u3_u2_n105 ) , .A1( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n143 ) );
  NAND2_X1 u2_u3_u2_U52 (.A1( u2_u3_u2_n104 ) , .A2( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n152 ) );
  NAND2_X1 u2_u3_u2_U53 (.A1( u2_u3_u2_n100 ) , .A2( u2_u3_u2_n105 ) , .ZN( u2_u3_u2_n132 ) );
  INV_X1 u2_u3_u2_U54 (.A( u2_u3_u2_n140 ) , .ZN( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U55 (.A( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n167 ) );
  INV_X1 u2_u3_u2_U56 (.ZN( u2_u3_u2_n187 ) , .A( u2_u3_u2_n99 ) );
  OAI21_X1 u2_u3_u2_U57 (.B1( u2_u3_u2_n137 ) , .B2( u2_u3_u2_n143 ) , .A( u2_u3_u2_n98 ) , .ZN( u2_u3_u2_n99 ) );
  NAND2_X1 u2_u3_u2_U58 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n113 ) );
  NAND2_X1 u2_u3_u2_U59 (.A1( u2_u3_u2_n106 ) , .A2( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n131 ) );
  AOI21_X1 u2_u3_u2_U6 (.B2( u2_u3_u2_n119 ) , .ZN( u2_u3_u2_n127 ) , .A( u2_u3_u2_n137 ) , .B1( u2_u3_u2_n155 ) );
  NAND2_X1 u2_u3_u2_U60 (.A1( u2_u3_u2_n103 ) , .A2( u2_u3_u2_n107 ) , .ZN( u2_u3_u2_n139 ) );
  NAND2_X1 u2_u3_u2_U61 (.A1( u2_u3_u2_n103 ) , .A2( u2_u3_u2_n105 ) , .ZN( u2_u3_u2_n133 ) );
  NAND2_X1 u2_u3_u2_U62 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n103 ) , .ZN( u2_u3_u2_n154 ) );
  NAND2_X1 u2_u3_u2_U63 (.A2( u2_u3_u2_n103 ) , .A1( u2_u3_u2_n104 ) , .ZN( u2_u3_u2_n119 ) );
  NAND2_X1 u2_u3_u2_U64 (.A2( u2_u3_u2_n107 ) , .A1( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n123 ) );
  NAND2_X1 u2_u3_u2_U65 (.A1( u2_u3_u2_n104 ) , .A2( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n122 ) );
  INV_X1 u2_u3_u2_U66 (.A( u2_u3_u2_n114 ) , .ZN( u2_u3_u2_n172 ) );
  NAND2_X1 u2_u3_u2_U67 (.A2( u2_u3_u2_n100 ) , .A1( u2_u3_u2_n102 ) , .ZN( u2_u3_u2_n116 ) );
  NAND2_X1 u2_u3_u2_U68 (.A1( u2_u3_u2_n102 ) , .A2( u2_u3_u2_n108 ) , .ZN( u2_u3_u2_n120 ) );
  NAND2_X1 u2_u3_u2_U69 (.A2( u2_u3_u2_n105 ) , .A1( u2_u3_u2_n106 ) , .ZN( u2_u3_u2_n117 ) );
  AOI21_X1 u2_u3_u2_U7 (.ZN( u2_u3_u2_n124 ) , .B1( u2_u3_u2_n131 ) , .B2( u2_u3_u2_n143 ) , .A( u2_u3_u2_n172 ) );
  NOR2_X1 u2_u3_u2_U70 (.A2( u2_u3_X_16 ) , .ZN( u2_u3_u2_n140 ) , .A1( u2_u3_u2_n166 ) );
  NOR2_X1 u2_u3_u2_U71 (.A2( u2_u3_X_13 ) , .A1( u2_u3_X_14 ) , .ZN( u2_u3_u2_n100 ) );
  NOR2_X1 u2_u3_u2_U72 (.A2( u2_u3_X_16 ) , .A1( u2_u3_X_17 ) , .ZN( u2_u3_u2_n138 ) );
  NOR2_X1 u2_u3_u2_U73 (.A2( u2_u3_X_15 ) , .A1( u2_u3_X_18 ) , .ZN( u2_u3_u2_n104 ) );
  NOR2_X1 u2_u3_u2_U74 (.A2( u2_u3_X_14 ) , .ZN( u2_u3_u2_n103 ) , .A1( u2_u3_u2_n174 ) );
  NOR2_X1 u2_u3_u2_U75 (.A2( u2_u3_X_15 ) , .ZN( u2_u3_u2_n102 ) , .A1( u2_u3_u2_n165 ) );
  NOR2_X1 u2_u3_u2_U76 (.A2( u2_u3_X_17 ) , .ZN( u2_u3_u2_n114 ) , .A1( u2_u3_u2_n169 ) );
  AND2_X1 u2_u3_u2_U77 (.A1( u2_u3_X_15 ) , .ZN( u2_u3_u2_n105 ) , .A2( u2_u3_u2_n165 ) );
  AND2_X1 u2_u3_u2_U78 (.A2( u2_u3_X_15 ) , .A1( u2_u3_X_18 ) , .ZN( u2_u3_u2_n107 ) );
  AND2_X1 u2_u3_u2_U79 (.A1( u2_u3_X_14 ) , .ZN( u2_u3_u2_n106 ) , .A2( u2_u3_u2_n174 ) );
  AOI21_X1 u2_u3_u2_U8 (.B2( u2_u3_u2_n120 ) , .B1( u2_u3_u2_n121 ) , .ZN( u2_u3_u2_n126 ) , .A( u2_u3_u2_n167 ) );
  AND2_X1 u2_u3_u2_U80 (.A1( u2_u3_X_13 ) , .A2( u2_u3_X_14 ) , .ZN( u2_u3_u2_n108 ) );
  INV_X1 u2_u3_u2_U81 (.A( u2_u3_X_16 ) , .ZN( u2_u3_u2_n169 ) );
  INV_X1 u2_u3_u2_U82 (.A( u2_u3_X_17 ) , .ZN( u2_u3_u2_n166 ) );
  INV_X1 u2_u3_u2_U83 (.A( u2_u3_X_13 ) , .ZN( u2_u3_u2_n174 ) );
  INV_X1 u2_u3_u2_U84 (.A( u2_u3_X_18 ) , .ZN( u2_u3_u2_n165 ) );
  NAND4_X1 u2_u3_u2_U85 (.ZN( u2_out3_24 ) , .A4( u2_u3_u2_n111 ) , .A3( u2_u3_u2_n112 ) , .A1( u2_u3_u2_n130 ) , .A2( u2_u3_u2_n187 ) );
  AOI221_X1 u2_u3_u2_U86 (.A( u2_u3_u2_n109 ) , .B1( u2_u3_u2_n110 ) , .ZN( u2_u3_u2_n111 ) , .C1( u2_u3_u2_n134 ) , .C2( u2_u3_u2_n170 ) , .B2( u2_u3_u2_n173 ) );
  AOI21_X1 u2_u3_u2_U87 (.ZN( u2_u3_u2_n112 ) , .B2( u2_u3_u2_n156 ) , .A( u2_u3_u2_n164 ) , .B1( u2_u3_u2_n181 ) );
  NAND4_X1 u2_u3_u2_U88 (.ZN( u2_out3_16 ) , .A4( u2_u3_u2_n128 ) , .A3( u2_u3_u2_n129 ) , .A1( u2_u3_u2_n130 ) , .A2( u2_u3_u2_n186 ) );
  AOI22_X1 u2_u3_u2_U89 (.A2( u2_u3_u2_n118 ) , .ZN( u2_u3_u2_n129 ) , .A1( u2_u3_u2_n140 ) , .B1( u2_u3_u2_n157 ) , .B2( u2_u3_u2_n170 ) );
  OAI22_X1 u2_u3_u2_U9 (.ZN( u2_u3_u2_n109 ) , .A2( u2_u3_u2_n113 ) , .B2( u2_u3_u2_n133 ) , .B1( u2_u3_u2_n167 ) , .A1( u2_u3_u2_n168 ) );
  INV_X1 u2_u3_u2_U90 (.A( u2_u3_u2_n163 ) , .ZN( u2_u3_u2_n186 ) );
  NAND4_X1 u2_u3_u2_U91 (.ZN( u2_out3_30 ) , .A4( u2_u3_u2_n147 ) , .A3( u2_u3_u2_n148 ) , .A2( u2_u3_u2_n149 ) , .A1( u2_u3_u2_n187 ) );
  AOI21_X1 u2_u3_u2_U92 (.B2( u2_u3_u2_n138 ) , .ZN( u2_u3_u2_n148 ) , .A( u2_u3_u2_n162 ) , .B1( u2_u3_u2_n182 ) );
  NOR3_X1 u2_u3_u2_U93 (.A3( u2_u3_u2_n144 ) , .A2( u2_u3_u2_n145 ) , .A1( u2_u3_u2_n146 ) , .ZN( u2_u3_u2_n147 ) );
  OR4_X1 u2_u3_u2_U94 (.ZN( u2_out3_6 ) , .A4( u2_u3_u2_n161 ) , .A3( u2_u3_u2_n162 ) , .A2( u2_u3_u2_n163 ) , .A1( u2_u3_u2_n164 ) );
  OR3_X1 u2_u3_u2_U95 (.A2( u2_u3_u2_n159 ) , .A1( u2_u3_u2_n160 ) , .ZN( u2_u3_u2_n161 ) , .A3( u2_u3_u2_n183 ) );
  AOI21_X1 u2_u3_u2_U96 (.B2( u2_u3_u2_n154 ) , .B1( u2_u3_u2_n155 ) , .ZN( u2_u3_u2_n159 ) , .A( u2_u3_u2_n167 ) );
  NAND3_X1 u2_u3_u2_U97 (.A2( u2_u3_u2_n117 ) , .A1( u2_u3_u2_n122 ) , .A3( u2_u3_u2_n123 ) , .ZN( u2_u3_u2_n134 ) );
  NAND3_X1 u2_u3_u2_U98 (.ZN( u2_u3_u2_n110 ) , .A2( u2_u3_u2_n131 ) , .A3( u2_u3_u2_n139 ) , .A1( u2_u3_u2_n154 ) );
  NAND3_X1 u2_u3_u2_U99 (.A2( u2_u3_u2_n100 ) , .ZN( u2_u3_u2_n101 ) , .A1( u2_u3_u2_n104 ) , .A3( u2_u3_u2_n114 ) );
  OAI22_X1 u2_u3_u3_U10 (.B1( u2_u3_u3_n113 ) , .A2( u2_u3_u3_n135 ) , .A1( u2_u3_u3_n150 ) , .B2( u2_u3_u3_n164 ) , .ZN( u2_u3_u3_n98 ) );
  OAI211_X1 u2_u3_u3_U11 (.B( u2_u3_u3_n106 ) , .ZN( u2_u3_u3_n119 ) , .C2( u2_u3_u3_n128 ) , .C1( u2_u3_u3_n167 ) , .A( u2_u3_u3_n181 ) );
  AOI221_X1 u2_u3_u3_U12 (.C1( u2_u3_u3_n105 ) , .ZN( u2_u3_u3_n106 ) , .A( u2_u3_u3_n131 ) , .B2( u2_u3_u3_n132 ) , .C2( u2_u3_u3_n133 ) , .B1( u2_u3_u3_n169 ) );
  INV_X1 u2_u3_u3_U13 (.ZN( u2_u3_u3_n181 ) , .A( u2_u3_u3_n98 ) );
  NAND2_X1 u2_u3_u3_U14 (.ZN( u2_u3_u3_n105 ) , .A2( u2_u3_u3_n130 ) , .A1( u2_u3_u3_n155 ) );
  AOI22_X1 u2_u3_u3_U15 (.B1( u2_u3_u3_n115 ) , .A2( u2_u3_u3_n116 ) , .ZN( u2_u3_u3_n123 ) , .B2( u2_u3_u3_n133 ) , .A1( u2_u3_u3_n169 ) );
  NAND2_X1 u2_u3_u3_U16 (.ZN( u2_u3_u3_n116 ) , .A2( u2_u3_u3_n151 ) , .A1( u2_u3_u3_n182 ) );
  NOR2_X1 u2_u3_u3_U17 (.ZN( u2_u3_u3_n126 ) , .A2( u2_u3_u3_n150 ) , .A1( u2_u3_u3_n164 ) );
  AOI21_X1 u2_u3_u3_U18 (.ZN( u2_u3_u3_n112 ) , .B2( u2_u3_u3_n146 ) , .B1( u2_u3_u3_n155 ) , .A( u2_u3_u3_n167 ) );
  NAND2_X1 u2_u3_u3_U19 (.A1( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n142 ) , .A2( u2_u3_u3_n164 ) );
  NAND2_X1 u2_u3_u3_U20 (.ZN( u2_u3_u3_n132 ) , .A2( u2_u3_u3_n152 ) , .A1( u2_u3_u3_n156 ) );
  INV_X1 u2_u3_u3_U21 (.A( u2_u3_u3_n133 ) , .ZN( u2_u3_u3_n165 ) );
  AND2_X1 u2_u3_u3_U22 (.A2( u2_u3_u3_n113 ) , .A1( u2_u3_u3_n114 ) , .ZN( u2_u3_u3_n151 ) );
  INV_X1 u2_u3_u3_U23 (.A( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n170 ) );
  NAND2_X1 u2_u3_u3_U24 (.A1( u2_u3_u3_n107 ) , .A2( u2_u3_u3_n108 ) , .ZN( u2_u3_u3_n140 ) );
  NAND2_X1 u2_u3_u3_U25 (.ZN( u2_u3_u3_n117 ) , .A1( u2_u3_u3_n124 ) , .A2( u2_u3_u3_n148 ) );
  NAND2_X1 u2_u3_u3_U26 (.ZN( u2_u3_u3_n143 ) , .A1( u2_u3_u3_n165 ) , .A2( u2_u3_u3_n167 ) );
  INV_X1 u2_u3_u3_U27 (.A( u2_u3_u3_n130 ) , .ZN( u2_u3_u3_n177 ) );
  INV_X1 u2_u3_u3_U28 (.A( u2_u3_u3_n128 ) , .ZN( u2_u3_u3_n176 ) );
  INV_X1 u2_u3_u3_U29 (.A( u2_u3_u3_n155 ) , .ZN( u2_u3_u3_n174 ) );
  INV_X1 u2_u3_u3_U3 (.A( u2_u3_u3_n140 ) , .ZN( u2_u3_u3_n182 ) );
  INV_X1 u2_u3_u3_U30 (.A( u2_u3_u3_n139 ) , .ZN( u2_u3_u3_n185 ) );
  NOR2_X1 u2_u3_u3_U31 (.ZN( u2_u3_u3_n135 ) , .A2( u2_u3_u3_n141 ) , .A1( u2_u3_u3_n169 ) );
  OAI222_X1 u2_u3_u3_U32 (.C2( u2_u3_u3_n107 ) , .A2( u2_u3_u3_n108 ) , .B1( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n138 ) , .B2( u2_u3_u3_n146 ) , .C1( u2_u3_u3_n154 ) , .A1( u2_u3_u3_n164 ) );
  NOR4_X1 u2_u3_u3_U33 (.A4( u2_u3_u3_n157 ) , .A3( u2_u3_u3_n158 ) , .A2( u2_u3_u3_n159 ) , .A1( u2_u3_u3_n160 ) , .ZN( u2_u3_u3_n161 ) );
  AOI21_X1 u2_u3_u3_U34 (.B2( u2_u3_u3_n152 ) , .B1( u2_u3_u3_n153 ) , .ZN( u2_u3_u3_n158 ) , .A( u2_u3_u3_n164 ) );
  AOI21_X1 u2_u3_u3_U35 (.A( u2_u3_u3_n149 ) , .B2( u2_u3_u3_n150 ) , .B1( u2_u3_u3_n151 ) , .ZN( u2_u3_u3_n159 ) );
  AOI21_X1 u2_u3_u3_U36 (.A( u2_u3_u3_n154 ) , .B2( u2_u3_u3_n155 ) , .B1( u2_u3_u3_n156 ) , .ZN( u2_u3_u3_n157 ) );
  AOI211_X1 u2_u3_u3_U37 (.ZN( u2_u3_u3_n109 ) , .A( u2_u3_u3_n119 ) , .C2( u2_u3_u3_n129 ) , .B( u2_u3_u3_n138 ) , .C1( u2_u3_u3_n141 ) );
  AOI211_X1 u2_u3_u3_U38 (.B( u2_u3_u3_n119 ) , .A( u2_u3_u3_n120 ) , .C2( u2_u3_u3_n121 ) , .ZN( u2_u3_u3_n122 ) , .C1( u2_u3_u3_n179 ) );
  INV_X1 u2_u3_u3_U39 (.A( u2_u3_u3_n156 ) , .ZN( u2_u3_u3_n179 ) );
  INV_X1 u2_u3_u3_U4 (.A( u2_u3_u3_n129 ) , .ZN( u2_u3_u3_n183 ) );
  OAI22_X1 u2_u3_u3_U40 (.B1( u2_u3_u3_n118 ) , .ZN( u2_u3_u3_n120 ) , .A1( u2_u3_u3_n135 ) , .B2( u2_u3_u3_n154 ) , .A2( u2_u3_u3_n178 ) );
  AND3_X1 u2_u3_u3_U41 (.ZN( u2_u3_u3_n118 ) , .A2( u2_u3_u3_n124 ) , .A1( u2_u3_u3_n144 ) , .A3( u2_u3_u3_n152 ) );
  INV_X1 u2_u3_u3_U42 (.A( u2_u3_u3_n121 ) , .ZN( u2_u3_u3_n164 ) );
  NAND2_X1 u2_u3_u3_U43 (.ZN( u2_u3_u3_n133 ) , .A1( u2_u3_u3_n154 ) , .A2( u2_u3_u3_n164 ) );
  NOR2_X1 u2_u3_u3_U44 (.A1( u2_u3_u3_n113 ) , .ZN( u2_u3_u3_n131 ) , .A2( u2_u3_u3_n154 ) );
  NAND2_X1 u2_u3_u3_U45 (.A1( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n150 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U46 (.A2( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n155 ) , .A1( u2_u3_u3_n97 ) );
  OAI211_X1 u2_u3_u3_U47 (.B( u2_u3_u3_n127 ) , .ZN( u2_u3_u3_n139 ) , .C1( u2_u3_u3_n150 ) , .C2( u2_u3_u3_n154 ) , .A( u2_u3_u3_n184 ) );
  INV_X1 u2_u3_u3_U48 (.A( u2_u3_u3_n125 ) , .ZN( u2_u3_u3_n184 ) );
  AOI221_X1 u2_u3_u3_U49 (.A( u2_u3_u3_n126 ) , .ZN( u2_u3_u3_n127 ) , .C2( u2_u3_u3_n132 ) , .C1( u2_u3_u3_n169 ) , .B2( u2_u3_u3_n170 ) , .B1( u2_u3_u3_n174 ) );
  INV_X1 u2_u3_u3_U5 (.A( u2_u3_u3_n117 ) , .ZN( u2_u3_u3_n178 ) );
  OAI22_X1 u2_u3_u3_U50 (.A1( u2_u3_u3_n124 ) , .ZN( u2_u3_u3_n125 ) , .B2( u2_u3_u3_n145 ) , .A2( u2_u3_u3_n165 ) , .B1( u2_u3_u3_n167 ) );
  INV_X1 u2_u3_u3_U51 (.A( u2_u3_u3_n141 ) , .ZN( u2_u3_u3_n167 ) );
  AOI21_X1 u2_u3_u3_U52 (.B2( u2_u3_u3_n114 ) , .B1( u2_u3_u3_n146 ) , .A( u2_u3_u3_n154 ) , .ZN( u2_u3_u3_n94 ) );
  AOI21_X1 u2_u3_u3_U53 (.ZN( u2_u3_u3_n110 ) , .B2( u2_u3_u3_n142 ) , .B1( u2_u3_u3_n186 ) , .A( u2_u3_u3_n95 ) );
  INV_X1 u2_u3_u3_U54 (.A( u2_u3_u3_n145 ) , .ZN( u2_u3_u3_n186 ) );
  AOI21_X1 u2_u3_u3_U55 (.B1( u2_u3_u3_n124 ) , .A( u2_u3_u3_n149 ) , .B2( u2_u3_u3_n155 ) , .ZN( u2_u3_u3_n95 ) );
  INV_X1 u2_u3_u3_U56 (.A( u2_u3_u3_n149 ) , .ZN( u2_u3_u3_n169 ) );
  NAND2_X1 u2_u3_u3_U57 (.ZN( u2_u3_u3_n124 ) , .A1( u2_u3_u3_n96 ) , .A2( u2_u3_u3_n97 ) );
  NAND2_X1 u2_u3_u3_U58 (.A2( u2_u3_u3_n100 ) , .ZN( u2_u3_u3_n146 ) , .A1( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U59 (.A1( u2_u3_u3_n101 ) , .ZN( u2_u3_u3_n145 ) , .A2( u2_u3_u3_n99 ) );
  AOI221_X1 u2_u3_u3_U6 (.A( u2_u3_u3_n131 ) , .C2( u2_u3_u3_n132 ) , .C1( u2_u3_u3_n133 ) , .ZN( u2_u3_u3_n134 ) , .B1( u2_u3_u3_n143 ) , .B2( u2_u3_u3_n177 ) );
  NAND2_X1 u2_u3_u3_U60 (.A1( u2_u3_u3_n100 ) , .ZN( u2_u3_u3_n156 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U61 (.A2( u2_u3_u3_n101 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n148 ) );
  NAND2_X1 u2_u3_u3_U62 (.A1( u2_u3_u3_n100 ) , .A2( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n128 ) );
  NAND2_X1 u2_u3_u3_U63 (.A2( u2_u3_u3_n101 ) , .A1( u2_u3_u3_n102 ) , .ZN( u2_u3_u3_n152 ) );
  NAND2_X1 u2_u3_u3_U64 (.A2( u2_u3_u3_n101 ) , .ZN( u2_u3_u3_n114 ) , .A1( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U65 (.ZN( u2_u3_u3_n107 ) , .A1( u2_u3_u3_n97 ) , .A2( u2_u3_u3_n99 ) );
  NAND2_X1 u2_u3_u3_U66 (.A2( u2_u3_u3_n100 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n113 ) );
  NAND2_X1 u2_u3_u3_U67 (.A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n153 ) , .A2( u2_u3_u3_n97 ) );
  NAND2_X1 u2_u3_u3_U68 (.A2( u2_u3_u3_n103 ) , .A1( u2_u3_u3_n104 ) , .ZN( u2_u3_u3_n130 ) );
  NAND2_X1 u2_u3_u3_U69 (.A2( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n144 ) , .A1( u2_u3_u3_n96 ) );
  OAI22_X1 u2_u3_u3_U7 (.B2( u2_u3_u3_n147 ) , .A2( u2_u3_u3_n148 ) , .ZN( u2_u3_u3_n160 ) , .B1( u2_u3_u3_n165 ) , .A1( u2_u3_u3_n168 ) );
  NAND2_X1 u2_u3_u3_U70 (.A1( u2_u3_u3_n102 ) , .A2( u2_u3_u3_n103 ) , .ZN( u2_u3_u3_n108 ) );
  NOR2_X1 u2_u3_u3_U71 (.A2( u2_u3_X_19 ) , .A1( u2_u3_X_20 ) , .ZN( u2_u3_u3_n99 ) );
  NOR2_X1 u2_u3_u3_U72 (.A2( u2_u3_X_21 ) , .A1( u2_u3_X_24 ) , .ZN( u2_u3_u3_n103 ) );
  NOR2_X1 u2_u3_u3_U73 (.A2( u2_u3_X_24 ) , .A1( u2_u3_u3_n171 ) , .ZN( u2_u3_u3_n97 ) );
  NOR2_X1 u2_u3_u3_U74 (.A2( u2_u3_X_23 ) , .ZN( u2_u3_u3_n141 ) , .A1( u2_u3_u3_n166 ) );
  NOR2_X1 u2_u3_u3_U75 (.A2( u2_u3_X_19 ) , .A1( u2_u3_u3_n172 ) , .ZN( u2_u3_u3_n96 ) );
  NAND2_X1 u2_u3_u3_U76 (.A1( u2_u3_X_22 ) , .A2( u2_u3_X_23 ) , .ZN( u2_u3_u3_n154 ) );
  NAND2_X1 u2_u3_u3_U77 (.A1( u2_u3_X_23 ) , .ZN( u2_u3_u3_n149 ) , .A2( u2_u3_u3_n166 ) );
  NOR2_X1 u2_u3_u3_U78 (.A2( u2_u3_X_22 ) , .A1( u2_u3_X_23 ) , .ZN( u2_u3_u3_n121 ) );
  AND2_X1 u2_u3_u3_U79 (.A1( u2_u3_X_24 ) , .ZN( u2_u3_u3_n101 ) , .A2( u2_u3_u3_n171 ) );
  AND3_X1 u2_u3_u3_U8 (.A3( u2_u3_u3_n144 ) , .A2( u2_u3_u3_n145 ) , .A1( u2_u3_u3_n146 ) , .ZN( u2_u3_u3_n147 ) );
  AND2_X1 u2_u3_u3_U80 (.A1( u2_u3_X_19 ) , .ZN( u2_u3_u3_n102 ) , .A2( u2_u3_u3_n172 ) );
  AND2_X1 u2_u3_u3_U81 (.A1( u2_u3_X_21 ) , .A2( u2_u3_X_24 ) , .ZN( u2_u3_u3_n100 ) );
  AND2_X1 u2_u3_u3_U82 (.A2( u2_u3_X_19 ) , .A1( u2_u3_X_20 ) , .ZN( u2_u3_u3_n104 ) );
  INV_X1 u2_u3_u3_U83 (.A( u2_u3_X_22 ) , .ZN( u2_u3_u3_n166 ) );
  INV_X1 u2_u3_u3_U84 (.A( u2_u3_X_21 ) , .ZN( u2_u3_u3_n171 ) );
  INV_X1 u2_u3_u3_U85 (.A( u2_u3_X_20 ) , .ZN( u2_u3_u3_n172 ) );
  NAND4_X1 u2_u3_u3_U86 (.ZN( u2_out3_26 ) , .A4( u2_u3_u3_n109 ) , .A3( u2_u3_u3_n110 ) , .A2( u2_u3_u3_n111 ) , .A1( u2_u3_u3_n173 ) );
  INV_X1 u2_u3_u3_U87 (.ZN( u2_u3_u3_n173 ) , .A( u2_u3_u3_n94 ) );
  OAI21_X1 u2_u3_u3_U88 (.ZN( u2_u3_u3_n111 ) , .B2( u2_u3_u3_n117 ) , .A( u2_u3_u3_n133 ) , .B1( u2_u3_u3_n176 ) );
  NAND4_X1 u2_u3_u3_U89 (.ZN( u2_out3_20 ) , .A4( u2_u3_u3_n122 ) , .A3( u2_u3_u3_n123 ) , .A1( u2_u3_u3_n175 ) , .A2( u2_u3_u3_n180 ) );
  INV_X1 u2_u3_u3_U9 (.A( u2_u3_u3_n143 ) , .ZN( u2_u3_u3_n168 ) );
  INV_X1 u2_u3_u3_U90 (.A( u2_u3_u3_n126 ) , .ZN( u2_u3_u3_n180 ) );
  INV_X1 u2_u3_u3_U91 (.A( u2_u3_u3_n112 ) , .ZN( u2_u3_u3_n175 ) );
  NAND4_X1 u2_u3_u3_U92 (.ZN( u2_out3_1 ) , .A4( u2_u3_u3_n161 ) , .A3( u2_u3_u3_n162 ) , .A2( u2_u3_u3_n163 ) , .A1( u2_u3_u3_n185 ) );
  NAND2_X1 u2_u3_u3_U93 (.ZN( u2_u3_u3_n163 ) , .A2( u2_u3_u3_n170 ) , .A1( u2_u3_u3_n176 ) );
  AOI22_X1 u2_u3_u3_U94 (.B2( u2_u3_u3_n140 ) , .B1( u2_u3_u3_n141 ) , .A2( u2_u3_u3_n142 ) , .ZN( u2_u3_u3_n162 ) , .A1( u2_u3_u3_n177 ) );
  OAI222_X1 u2_u3_u3_U95 (.C1( u2_u3_u3_n128 ) , .ZN( u2_u3_u3_n137 ) , .B1( u2_u3_u3_n148 ) , .A2( u2_u3_u3_n150 ) , .B2( u2_u3_u3_n154 ) , .C2( u2_u3_u3_n164 ) , .A1( u2_u3_u3_n167 ) );
  OR4_X1 u2_u3_u3_U96 (.ZN( u2_out3_10 ) , .A4( u2_u3_u3_n136 ) , .A3( u2_u3_u3_n137 ) , .A1( u2_u3_u3_n138 ) , .A2( u2_u3_u3_n139 ) );
  OAI221_X1 u2_u3_u3_U97 (.A( u2_u3_u3_n134 ) , .B2( u2_u3_u3_n135 ) , .ZN( u2_u3_u3_n136 ) , .C1( u2_u3_u3_n149 ) , .B1( u2_u3_u3_n151 ) , .C2( u2_u3_u3_n183 ) );
  NAND3_X1 u2_u3_u3_U98 (.A1( u2_u3_u3_n114 ) , .ZN( u2_u3_u3_n115 ) , .A2( u2_u3_u3_n145 ) , .A3( u2_u3_u3_n153 ) );
  NAND3_X1 u2_u3_u3_U99 (.ZN( u2_u3_u3_n129 ) , .A2( u2_u3_u3_n144 ) , .A1( u2_u3_u3_n153 ) , .A3( u2_u3_u3_n182 ) );
  XOR2_X1 u2_u7_U1 (.B( u2_K8_9 ) , .A( u2_R6_6 ) , .Z( u2_u7_X_9 ) );
  XOR2_X1 u2_u7_U2 (.B( u2_K8_8 ) , .A( u2_R6_5 ) , .Z( u2_u7_X_8 ) );
  XOR2_X1 u2_u7_U3 (.B( u2_K8_7 ) , .A( u2_R6_4 ) , .Z( u2_u7_X_7 ) );
  XOR2_X1 u2_u7_U46 (.B( u2_K8_12 ) , .A( u2_R6_9 ) , .Z( u2_u7_X_12 ) );
  XOR2_X1 u2_u7_U47 (.B( u2_K8_11 ) , .A( u2_R6_8 ) , .Z( u2_u7_X_11 ) );
  XOR2_X1 u2_u7_U48 (.B( u2_K8_10 ) , .A( u2_R6_7 ) , .Z( u2_u7_X_10 ) );
  AOI21_X1 u2_u7_u1_U10 (.B2( u2_u7_u1_n155 ) , .B1( u2_u7_u1_n156 ) , .ZN( u2_u7_u1_n157 ) , .A( u2_u7_u1_n174 ) );
  NAND3_X1 u2_u7_u1_U100 (.ZN( u2_u7_u1_n113 ) , .A1( u2_u7_u1_n120 ) , .A3( u2_u7_u1_n133 ) , .A2( u2_u7_u1_n155 ) );
  NAND2_X1 u2_u7_u1_U11 (.ZN( u2_u7_u1_n140 ) , .A2( u2_u7_u1_n150 ) , .A1( u2_u7_u1_n155 ) );
  NAND2_X1 u2_u7_u1_U12 (.A1( u2_u7_u1_n131 ) , .ZN( u2_u7_u1_n147 ) , .A2( u2_u7_u1_n153 ) );
  AOI22_X1 u2_u7_u1_U13 (.B2( u2_u7_u1_n136 ) , .A2( u2_u7_u1_n137 ) , .ZN( u2_u7_u1_n143 ) , .A1( u2_u7_u1_n171 ) , .B1( u2_u7_u1_n173 ) );
  INV_X1 u2_u7_u1_U14 (.A( u2_u7_u1_n147 ) , .ZN( u2_u7_u1_n181 ) );
  INV_X1 u2_u7_u1_U15 (.A( u2_u7_u1_n139 ) , .ZN( u2_u7_u1_n174 ) );
  OR4_X1 u2_u7_u1_U16 (.A4( u2_u7_u1_n106 ) , .A3( u2_u7_u1_n107 ) , .ZN( u2_u7_u1_n108 ) , .A1( u2_u7_u1_n117 ) , .A2( u2_u7_u1_n184 ) );
  AOI21_X1 u2_u7_u1_U17 (.ZN( u2_u7_u1_n106 ) , .A( u2_u7_u1_n112 ) , .B1( u2_u7_u1_n154 ) , .B2( u2_u7_u1_n156 ) );
  AOI21_X1 u2_u7_u1_U18 (.ZN( u2_u7_u1_n107 ) , .B1( u2_u7_u1_n134 ) , .B2( u2_u7_u1_n149 ) , .A( u2_u7_u1_n174 ) );
  INV_X1 u2_u7_u1_U19 (.A( u2_u7_u1_n101 ) , .ZN( u2_u7_u1_n184 ) );
  INV_X1 u2_u7_u1_U20 (.A( u2_u7_u1_n112 ) , .ZN( u2_u7_u1_n171 ) );
  NAND2_X1 u2_u7_u1_U21 (.ZN( u2_u7_u1_n141 ) , .A1( u2_u7_u1_n153 ) , .A2( u2_u7_u1_n156 ) );
  AND2_X1 u2_u7_u1_U22 (.A1( u2_u7_u1_n123 ) , .ZN( u2_u7_u1_n134 ) , .A2( u2_u7_u1_n161 ) );
  NAND2_X1 u2_u7_u1_U23 (.A2( u2_u7_u1_n115 ) , .A1( u2_u7_u1_n116 ) , .ZN( u2_u7_u1_n148 ) );
  NAND2_X1 u2_u7_u1_U24 (.A2( u2_u7_u1_n133 ) , .A1( u2_u7_u1_n135 ) , .ZN( u2_u7_u1_n159 ) );
  NAND2_X1 u2_u7_u1_U25 (.A2( u2_u7_u1_n115 ) , .A1( u2_u7_u1_n120 ) , .ZN( u2_u7_u1_n132 ) );
  INV_X1 u2_u7_u1_U26 (.A( u2_u7_u1_n154 ) , .ZN( u2_u7_u1_n178 ) );
  INV_X1 u2_u7_u1_U27 (.A( u2_u7_u1_n151 ) , .ZN( u2_u7_u1_n183 ) );
  AND2_X1 u2_u7_u1_U28 (.A1( u2_u7_u1_n129 ) , .A2( u2_u7_u1_n133 ) , .ZN( u2_u7_u1_n149 ) );
  INV_X1 u2_u7_u1_U29 (.A( u2_u7_u1_n131 ) , .ZN( u2_u7_u1_n180 ) );
  INV_X1 u2_u7_u1_U3 (.A( u2_u7_u1_n159 ) , .ZN( u2_u7_u1_n182 ) );
  OAI221_X1 u2_u7_u1_U30 (.A( u2_u7_u1_n119 ) , .C2( u2_u7_u1_n129 ) , .ZN( u2_u7_u1_n138 ) , .B2( u2_u7_u1_n152 ) , .C1( u2_u7_u1_n174 ) , .B1( u2_u7_u1_n187 ) );
  INV_X1 u2_u7_u1_U31 (.A( u2_u7_u1_n148 ) , .ZN( u2_u7_u1_n187 ) );
  AOI211_X1 u2_u7_u1_U32 (.B( u2_u7_u1_n117 ) , .A( u2_u7_u1_n118 ) , .ZN( u2_u7_u1_n119 ) , .C2( u2_u7_u1_n146 ) , .C1( u2_u7_u1_n159 ) );
  NOR2_X1 u2_u7_u1_U33 (.A1( u2_u7_u1_n168 ) , .A2( u2_u7_u1_n176 ) , .ZN( u2_u7_u1_n98 ) );
  AOI211_X1 u2_u7_u1_U34 (.B( u2_u7_u1_n162 ) , .A( u2_u7_u1_n163 ) , .C2( u2_u7_u1_n164 ) , .ZN( u2_u7_u1_n165 ) , .C1( u2_u7_u1_n171 ) );
  AOI21_X1 u2_u7_u1_U35 (.A( u2_u7_u1_n160 ) , .B2( u2_u7_u1_n161 ) , .ZN( u2_u7_u1_n162 ) , .B1( u2_u7_u1_n182 ) );
  OR2_X1 u2_u7_u1_U36 (.A2( u2_u7_u1_n157 ) , .A1( u2_u7_u1_n158 ) , .ZN( u2_u7_u1_n163 ) );
  NAND2_X1 u2_u7_u1_U37 (.A1( u2_u7_u1_n128 ) , .ZN( u2_u7_u1_n146 ) , .A2( u2_u7_u1_n160 ) );
  NAND2_X1 u2_u7_u1_U38 (.A2( u2_u7_u1_n112 ) , .ZN( u2_u7_u1_n139 ) , .A1( u2_u7_u1_n152 ) );
  NAND2_X1 u2_u7_u1_U39 (.A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n156 ) , .A2( u2_u7_u1_n99 ) );
  AOI221_X1 u2_u7_u1_U4 (.A( u2_u7_u1_n138 ) , .C2( u2_u7_u1_n139 ) , .C1( u2_u7_u1_n140 ) , .B2( u2_u7_u1_n141 ) , .ZN( u2_u7_u1_n142 ) , .B1( u2_u7_u1_n175 ) );
  AOI221_X1 u2_u7_u1_U40 (.B1( u2_u7_u1_n140 ) , .ZN( u2_u7_u1_n167 ) , .B2( u2_u7_u1_n172 ) , .C2( u2_u7_u1_n175 ) , .C1( u2_u7_u1_n178 ) , .A( u2_u7_u1_n188 ) );
  INV_X1 u2_u7_u1_U41 (.ZN( u2_u7_u1_n188 ) , .A( u2_u7_u1_n97 ) );
  AOI211_X1 u2_u7_u1_U42 (.A( u2_u7_u1_n118 ) , .C1( u2_u7_u1_n132 ) , .C2( u2_u7_u1_n139 ) , .B( u2_u7_u1_n96 ) , .ZN( u2_u7_u1_n97 ) );
  AOI21_X1 u2_u7_u1_U43 (.B2( u2_u7_u1_n121 ) , .B1( u2_u7_u1_n135 ) , .A( u2_u7_u1_n152 ) , .ZN( u2_u7_u1_n96 ) );
  NOR2_X1 u2_u7_u1_U44 (.ZN( u2_u7_u1_n117 ) , .A1( u2_u7_u1_n121 ) , .A2( u2_u7_u1_n160 ) );
  OAI21_X1 u2_u7_u1_U45 (.B2( u2_u7_u1_n123 ) , .ZN( u2_u7_u1_n145 ) , .B1( u2_u7_u1_n160 ) , .A( u2_u7_u1_n185 ) );
  INV_X1 u2_u7_u1_U46 (.A( u2_u7_u1_n122 ) , .ZN( u2_u7_u1_n185 ) );
  AOI21_X1 u2_u7_u1_U47 (.B2( u2_u7_u1_n120 ) , .B1( u2_u7_u1_n121 ) , .ZN( u2_u7_u1_n122 ) , .A( u2_u7_u1_n128 ) );
  AOI21_X1 u2_u7_u1_U48 (.A( u2_u7_u1_n128 ) , .B2( u2_u7_u1_n129 ) , .ZN( u2_u7_u1_n130 ) , .B1( u2_u7_u1_n150 ) );
  NAND2_X1 u2_u7_u1_U49 (.ZN( u2_u7_u1_n112 ) , .A1( u2_u7_u1_n169 ) , .A2( u2_u7_u1_n170 ) );
  AOI211_X1 u2_u7_u1_U5 (.ZN( u2_u7_u1_n124 ) , .A( u2_u7_u1_n138 ) , .C2( u2_u7_u1_n139 ) , .B( u2_u7_u1_n145 ) , .C1( u2_u7_u1_n147 ) );
  NAND2_X1 u2_u7_u1_U50 (.ZN( u2_u7_u1_n129 ) , .A2( u2_u7_u1_n95 ) , .A1( u2_u7_u1_n98 ) );
  NAND2_X1 u2_u7_u1_U51 (.A1( u2_u7_u1_n102 ) , .ZN( u2_u7_u1_n154 ) , .A2( u2_u7_u1_n99 ) );
  NAND2_X1 u2_u7_u1_U52 (.A2( u2_u7_u1_n100 ) , .ZN( u2_u7_u1_n135 ) , .A1( u2_u7_u1_n99 ) );
  AOI21_X1 u2_u7_u1_U53 (.A( u2_u7_u1_n152 ) , .B2( u2_u7_u1_n153 ) , .B1( u2_u7_u1_n154 ) , .ZN( u2_u7_u1_n158 ) );
  INV_X1 u2_u7_u1_U54 (.A( u2_u7_u1_n160 ) , .ZN( u2_u7_u1_n175 ) );
  NAND2_X1 u2_u7_u1_U55 (.A1( u2_u7_u1_n100 ) , .ZN( u2_u7_u1_n116 ) , .A2( u2_u7_u1_n95 ) );
  NAND2_X1 u2_u7_u1_U56 (.A1( u2_u7_u1_n102 ) , .ZN( u2_u7_u1_n131 ) , .A2( u2_u7_u1_n95 ) );
  NAND2_X1 u2_u7_u1_U57 (.A2( u2_u7_u1_n104 ) , .ZN( u2_u7_u1_n121 ) , .A1( u2_u7_u1_n98 ) );
  NAND2_X1 u2_u7_u1_U58 (.A1( u2_u7_u1_n103 ) , .ZN( u2_u7_u1_n153 ) , .A2( u2_u7_u1_n98 ) );
  NAND2_X1 u2_u7_u1_U59 (.A2( u2_u7_u1_n104 ) , .A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n133 ) );
  AOI22_X1 u2_u7_u1_U6 (.B2( u2_u7_u1_n113 ) , .A2( u2_u7_u1_n114 ) , .ZN( u2_u7_u1_n125 ) , .A1( u2_u7_u1_n171 ) , .B1( u2_u7_u1_n173 ) );
  NAND2_X1 u2_u7_u1_U60 (.ZN( u2_u7_u1_n150 ) , .A2( u2_u7_u1_n98 ) , .A1( u2_u7_u1_n99 ) );
  NAND2_X1 u2_u7_u1_U61 (.A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n155 ) , .A2( u2_u7_u1_n95 ) );
  OAI21_X1 u2_u7_u1_U62 (.ZN( u2_u7_u1_n109 ) , .B1( u2_u7_u1_n129 ) , .B2( u2_u7_u1_n160 ) , .A( u2_u7_u1_n167 ) );
  NAND2_X1 u2_u7_u1_U63 (.A2( u2_u7_u1_n100 ) , .A1( u2_u7_u1_n103 ) , .ZN( u2_u7_u1_n120 ) );
  NAND2_X1 u2_u7_u1_U64 (.A1( u2_u7_u1_n102 ) , .A2( u2_u7_u1_n104 ) , .ZN( u2_u7_u1_n115 ) );
  NAND2_X1 u2_u7_u1_U65 (.A2( u2_u7_u1_n100 ) , .A1( u2_u7_u1_n104 ) , .ZN( u2_u7_u1_n151 ) );
  NAND2_X1 u2_u7_u1_U66 (.A2( u2_u7_u1_n103 ) , .A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n161 ) );
  INV_X1 u2_u7_u1_U67 (.A( u2_u7_u1_n152 ) , .ZN( u2_u7_u1_n173 ) );
  INV_X1 u2_u7_u1_U68 (.A( u2_u7_u1_n128 ) , .ZN( u2_u7_u1_n172 ) );
  NAND2_X1 u2_u7_u1_U69 (.A2( u2_u7_u1_n102 ) , .A1( u2_u7_u1_n103 ) , .ZN( u2_u7_u1_n123 ) );
  NAND2_X1 u2_u7_u1_U7 (.ZN( u2_u7_u1_n114 ) , .A1( u2_u7_u1_n134 ) , .A2( u2_u7_u1_n156 ) );
  NOR2_X1 u2_u7_u1_U70 (.A2( u2_u7_X_7 ) , .A1( u2_u7_X_8 ) , .ZN( u2_u7_u1_n95 ) );
  NOR2_X1 u2_u7_u1_U71 (.A1( u2_u7_X_12 ) , .A2( u2_u7_X_9 ) , .ZN( u2_u7_u1_n100 ) );
  NOR2_X1 u2_u7_u1_U72 (.A2( u2_u7_X_8 ) , .A1( u2_u7_u1_n177 ) , .ZN( u2_u7_u1_n99 ) );
  NOR2_X1 u2_u7_u1_U73 (.A2( u2_u7_X_12 ) , .ZN( u2_u7_u1_n102 ) , .A1( u2_u7_u1_n176 ) );
  NOR2_X1 u2_u7_u1_U74 (.A2( u2_u7_X_9 ) , .ZN( u2_u7_u1_n105 ) , .A1( u2_u7_u1_n168 ) );
  NAND2_X1 u2_u7_u1_U75 (.A1( u2_u7_X_10 ) , .ZN( u2_u7_u1_n160 ) , .A2( u2_u7_u1_n169 ) );
  NAND2_X1 u2_u7_u1_U76 (.A2( u2_u7_X_10 ) , .A1( u2_u7_X_11 ) , .ZN( u2_u7_u1_n152 ) );
  NAND2_X1 u2_u7_u1_U77 (.A1( u2_u7_X_11 ) , .ZN( u2_u7_u1_n128 ) , .A2( u2_u7_u1_n170 ) );
  AND2_X1 u2_u7_u1_U78 (.A2( u2_u7_X_7 ) , .A1( u2_u7_X_8 ) , .ZN( u2_u7_u1_n104 ) );
  AND2_X1 u2_u7_u1_U79 (.A1( u2_u7_X_8 ) , .ZN( u2_u7_u1_n103 ) , .A2( u2_u7_u1_n177 ) );
  NOR2_X1 u2_u7_u1_U8 (.A1( u2_u7_u1_n112 ) , .A2( u2_u7_u1_n116 ) , .ZN( u2_u7_u1_n118 ) );
  INV_X1 u2_u7_u1_U80 (.A( u2_u7_X_10 ) , .ZN( u2_u7_u1_n170 ) );
  INV_X1 u2_u7_u1_U81 (.A( u2_u7_X_9 ) , .ZN( u2_u7_u1_n176 ) );
  INV_X1 u2_u7_u1_U82 (.A( u2_u7_X_11 ) , .ZN( u2_u7_u1_n169 ) );
  INV_X1 u2_u7_u1_U83 (.A( u2_u7_X_12 ) , .ZN( u2_u7_u1_n168 ) );
  INV_X1 u2_u7_u1_U84 (.A( u2_u7_X_7 ) , .ZN( u2_u7_u1_n177 ) );
  NAND4_X1 u2_u7_u1_U85 (.ZN( u2_out7_28 ) , .A4( u2_u7_u1_n124 ) , .A3( u2_u7_u1_n125 ) , .A2( u2_u7_u1_n126 ) , .A1( u2_u7_u1_n127 ) );
  OAI21_X1 u2_u7_u1_U86 (.ZN( u2_u7_u1_n127 ) , .B2( u2_u7_u1_n139 ) , .B1( u2_u7_u1_n175 ) , .A( u2_u7_u1_n183 ) );
  OAI21_X1 u2_u7_u1_U87 (.ZN( u2_u7_u1_n126 ) , .B2( u2_u7_u1_n140 ) , .A( u2_u7_u1_n146 ) , .B1( u2_u7_u1_n178 ) );
  NAND4_X1 u2_u7_u1_U88 (.ZN( u2_out7_18 ) , .A4( u2_u7_u1_n165 ) , .A3( u2_u7_u1_n166 ) , .A1( u2_u7_u1_n167 ) , .A2( u2_u7_u1_n186 ) );
  AOI22_X1 u2_u7_u1_U89 (.B2( u2_u7_u1_n146 ) , .B1( u2_u7_u1_n147 ) , .A2( u2_u7_u1_n148 ) , .ZN( u2_u7_u1_n166 ) , .A1( u2_u7_u1_n172 ) );
  OAI21_X1 u2_u7_u1_U9 (.ZN( u2_u7_u1_n101 ) , .B1( u2_u7_u1_n141 ) , .A( u2_u7_u1_n146 ) , .B2( u2_u7_u1_n183 ) );
  INV_X1 u2_u7_u1_U90 (.A( u2_u7_u1_n145 ) , .ZN( u2_u7_u1_n186 ) );
  NAND4_X1 u2_u7_u1_U91 (.ZN( u2_out7_2 ) , .A4( u2_u7_u1_n142 ) , .A3( u2_u7_u1_n143 ) , .A2( u2_u7_u1_n144 ) , .A1( u2_u7_u1_n179 ) );
  OAI21_X1 u2_u7_u1_U92 (.B2( u2_u7_u1_n132 ) , .ZN( u2_u7_u1_n144 ) , .A( u2_u7_u1_n146 ) , .B1( u2_u7_u1_n180 ) );
  INV_X1 u2_u7_u1_U93 (.A( u2_u7_u1_n130 ) , .ZN( u2_u7_u1_n179 ) );
  OR4_X1 u2_u7_u1_U94 (.ZN( u2_out7_13 ) , .A4( u2_u7_u1_n108 ) , .A3( u2_u7_u1_n109 ) , .A2( u2_u7_u1_n110 ) , .A1( u2_u7_u1_n111 ) );
  AOI21_X1 u2_u7_u1_U95 (.ZN( u2_u7_u1_n111 ) , .A( u2_u7_u1_n128 ) , .B2( u2_u7_u1_n131 ) , .B1( u2_u7_u1_n135 ) );
  AOI21_X1 u2_u7_u1_U96 (.ZN( u2_u7_u1_n110 ) , .A( u2_u7_u1_n116 ) , .B1( u2_u7_u1_n152 ) , .B2( u2_u7_u1_n160 ) );
  NAND3_X1 u2_u7_u1_U97 (.A3( u2_u7_u1_n149 ) , .A2( u2_u7_u1_n150 ) , .A1( u2_u7_u1_n151 ) , .ZN( u2_u7_u1_n164 ) );
  NAND3_X1 u2_u7_u1_U98 (.A3( u2_u7_u1_n134 ) , .A2( u2_u7_u1_n135 ) , .ZN( u2_u7_u1_n136 ) , .A1( u2_u7_u1_n151 ) );
  NAND3_X1 u2_u7_u1_U99 (.A1( u2_u7_u1_n133 ) , .ZN( u2_u7_u1_n137 ) , .A2( u2_u7_u1_n154 ) , .A3( u2_u7_u1_n181 ) );
  XOR2_X1 u2_u8_U1 (.B( u2_K9_9 ) , .A( u2_R7_6 ) , .Z( u2_u8_X_9 ) );
  XOR2_X1 u2_u8_U16 (.B( u2_K9_3 ) , .A( u2_R7_2 ) , .Z( u2_u8_X_3 ) );
  XOR2_X1 u2_u8_U2 (.B( u2_K9_8 ) , .A( u2_R7_5 ) , .Z( u2_u8_X_8 ) );
  XOR2_X1 u2_u8_U27 (.B( u2_K9_2 ) , .A( u2_R7_1 ) , .Z( u2_u8_X_2 ) );
  XOR2_X1 u2_u8_U3 (.B( u2_K9_7 ) , .A( u2_R7_4 ) , .Z( u2_u8_X_7 ) );
  XOR2_X1 u2_u8_U38 (.B( u2_K9_1 ) , .A( u2_R7_32 ) , .Z( u2_u8_X_1 ) );
  XOR2_X1 u2_u8_U4 (.B( u2_K9_6 ) , .A( u2_R7_5 ) , .Z( u2_u8_X_6 ) );
  XOR2_X1 u2_u8_U40 (.B( u2_K9_18 ) , .A( u2_R7_13 ) , .Z( u2_u8_X_18 ) );
  XOR2_X1 u2_u8_U41 (.B( u2_K9_17 ) , .A( u2_R7_12 ) , .Z( u2_u8_X_17 ) );
  XOR2_X1 u2_u8_U42 (.B( u2_K9_16 ) , .A( u2_R7_11 ) , .Z( u2_u8_X_16 ) );
  XOR2_X1 u2_u8_U43 (.B( u2_K9_15 ) , .A( u2_R7_10 ) , .Z( u2_u8_X_15 ) );
  XOR2_X1 u2_u8_U44 (.B( u2_K9_14 ) , .A( u2_R7_9 ) , .Z( u2_u8_X_14 ) );
  XOR2_X1 u2_u8_U45 (.B( u2_K9_13 ) , .A( u2_R7_8 ) , .Z( u2_u8_X_13 ) );
  XOR2_X1 u2_u8_U46 (.B( u2_K9_12 ) , .A( u2_R7_9 ) , .Z( u2_u8_X_12 ) );
  XOR2_X1 u2_u8_U47 (.B( u2_K9_11 ) , .A( u2_R7_8 ) , .Z( u2_u8_X_11 ) );
  XOR2_X1 u2_u8_U48 (.B( u2_K9_10 ) , .A( u2_R7_7 ) , .Z( u2_u8_X_10 ) );
  XOR2_X1 u2_u8_U5 (.B( u2_K9_5 ) , .A( u2_R7_4 ) , .Z( u2_u8_X_5 ) );
  XOR2_X1 u2_u8_U6 (.B( u2_K9_4 ) , .A( u2_R7_3 ) , .Z( u2_u8_X_4 ) );
  AND2_X1 u2_u8_u0_U10 (.A1( u2_u8_u0_n131 ) , .ZN( u2_u8_u0_n141 ) , .A2( u2_u8_u0_n150 ) );
  AND3_X1 u2_u8_u0_U11 (.A2( u2_u8_u0_n112 ) , .ZN( u2_u8_u0_n127 ) , .A3( u2_u8_u0_n130 ) , .A1( u2_u8_u0_n148 ) );
  AND2_X1 u2_u8_u0_U12 (.ZN( u2_u8_u0_n107 ) , .A1( u2_u8_u0_n130 ) , .A2( u2_u8_u0_n140 ) );
  AND2_X1 u2_u8_u0_U13 (.A2( u2_u8_u0_n129 ) , .A1( u2_u8_u0_n130 ) , .ZN( u2_u8_u0_n151 ) );
  AND2_X1 u2_u8_u0_U14 (.A1( u2_u8_u0_n108 ) , .A2( u2_u8_u0_n125 ) , .ZN( u2_u8_u0_n145 ) );
  INV_X1 u2_u8_u0_U15 (.A( u2_u8_u0_n143 ) , .ZN( u2_u8_u0_n173 ) );
  NOR2_X1 u2_u8_u0_U16 (.A2( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n147 ) , .A1( u2_u8_u0_n160 ) );
  AOI21_X1 u2_u8_u0_U17 (.B1( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n132 ) , .A( u2_u8_u0_n165 ) , .B2( u2_u8_u0_n93 ) );
  OAI22_X1 u2_u8_u0_U18 (.B1( u2_u8_u0_n131 ) , .A1( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n147 ) , .A2( u2_u8_u0_n90 ) , .ZN( u2_u8_u0_n91 ) );
  AND3_X1 u2_u8_u0_U19 (.A3( u2_u8_u0_n121 ) , .A2( u2_u8_u0_n125 ) , .A1( u2_u8_u0_n148 ) , .ZN( u2_u8_u0_n90 ) );
  OAI22_X1 u2_u8_u0_U20 (.B1( u2_u8_u0_n125 ) , .ZN( u2_u8_u0_n126 ) , .A1( u2_u8_u0_n138 ) , .A2( u2_u8_u0_n146 ) , .B2( u2_u8_u0_n147 ) );
  NOR2_X1 u2_u8_u0_U21 (.A1( u2_u8_u0_n163 ) , .A2( u2_u8_u0_n164 ) , .ZN( u2_u8_u0_n95 ) );
  AOI22_X1 u2_u8_u0_U22 (.B2( u2_u8_u0_n109 ) , .A2( u2_u8_u0_n110 ) , .ZN( u2_u8_u0_n111 ) , .B1( u2_u8_u0_n118 ) , .A1( u2_u8_u0_n160 ) );
  NAND2_X1 u2_u8_u0_U23 (.A2( u2_u8_u0_n102 ) , .A1( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n149 ) );
  INV_X1 u2_u8_u0_U24 (.A( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n161 ) );
  INV_X1 u2_u8_u0_U25 (.A( u2_u8_u0_n118 ) , .ZN( u2_u8_u0_n158 ) );
  NAND2_X1 u2_u8_u0_U26 (.A2( u2_u8_u0_n100 ) , .ZN( u2_u8_u0_n131 ) , .A1( u2_u8_u0_n92 ) );
  NAND2_X1 u2_u8_u0_U27 (.ZN( u2_u8_u0_n108 ) , .A1( u2_u8_u0_n92 ) , .A2( u2_u8_u0_n94 ) );
  AOI21_X1 u2_u8_u0_U28 (.ZN( u2_u8_u0_n104 ) , .B1( u2_u8_u0_n107 ) , .B2( u2_u8_u0_n141 ) , .A( u2_u8_u0_n144 ) );
  AOI21_X1 u2_u8_u0_U29 (.B1( u2_u8_u0_n127 ) , .B2( u2_u8_u0_n129 ) , .A( u2_u8_u0_n138 ) , .ZN( u2_u8_u0_n96 ) );
  INV_X1 u2_u8_u0_U3 (.A( u2_u8_u0_n113 ) , .ZN( u2_u8_u0_n166 ) );
  NAND2_X1 u2_u8_u0_U30 (.A2( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n114 ) , .A1( u2_u8_u0_n92 ) );
  NOR2_X1 u2_u8_u0_U31 (.A1( u2_u8_u0_n120 ) , .ZN( u2_u8_u0_n143 ) , .A2( u2_u8_u0_n167 ) );
  OAI221_X1 u2_u8_u0_U32 (.C1( u2_u8_u0_n112 ) , .ZN( u2_u8_u0_n120 ) , .B1( u2_u8_u0_n138 ) , .B2( u2_u8_u0_n141 ) , .C2( u2_u8_u0_n147 ) , .A( u2_u8_u0_n172 ) );
  AOI211_X1 u2_u8_u0_U33 (.B( u2_u8_u0_n115 ) , .A( u2_u8_u0_n116 ) , .C2( u2_u8_u0_n117 ) , .C1( u2_u8_u0_n118 ) , .ZN( u2_u8_u0_n119 ) );
  NAND2_X1 u2_u8_u0_U34 (.A2( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n140 ) , .A1( u2_u8_u0_n94 ) );
  NAND2_X1 u2_u8_u0_U35 (.A1( u2_u8_u0_n100 ) , .A2( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n125 ) );
  NAND2_X1 u2_u8_u0_U36 (.A1( u2_u8_u0_n101 ) , .A2( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n150 ) );
  INV_X1 u2_u8_u0_U37 (.A( u2_u8_u0_n138 ) , .ZN( u2_u8_u0_n160 ) );
  NAND2_X1 u2_u8_u0_U38 (.A2( u2_u8_u0_n100 ) , .A1( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n139 ) );
  NAND2_X1 u2_u8_u0_U39 (.ZN( u2_u8_u0_n112 ) , .A2( u2_u8_u0_n92 ) , .A1( u2_u8_u0_n93 ) );
  AOI21_X1 u2_u8_u0_U4 (.B1( u2_u8_u0_n114 ) , .ZN( u2_u8_u0_n115 ) , .B2( u2_u8_u0_n129 ) , .A( u2_u8_u0_n161 ) );
  NAND2_X1 u2_u8_u0_U40 (.A1( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n130 ) , .A2( u2_u8_u0_n94 ) );
  INV_X1 u2_u8_u0_U41 (.ZN( u2_u8_u0_n172 ) , .A( u2_u8_u0_n88 ) );
  OAI222_X1 u2_u8_u0_U42 (.C1( u2_u8_u0_n108 ) , .A1( u2_u8_u0_n125 ) , .B2( u2_u8_u0_n128 ) , .B1( u2_u8_u0_n144 ) , .A2( u2_u8_u0_n158 ) , .C2( u2_u8_u0_n161 ) , .ZN( u2_u8_u0_n88 ) );
  NAND2_X1 u2_u8_u0_U43 (.A2( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n121 ) , .A1( u2_u8_u0_n93 ) );
  OR3_X1 u2_u8_u0_U44 (.A3( u2_u8_u0_n152 ) , .A2( u2_u8_u0_n153 ) , .A1( u2_u8_u0_n154 ) , .ZN( u2_u8_u0_n155 ) );
  AOI21_X1 u2_u8_u0_U45 (.A( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n145 ) , .B1( u2_u8_u0_n146 ) , .ZN( u2_u8_u0_n154 ) );
  AOI21_X1 u2_u8_u0_U46 (.B2( u2_u8_u0_n150 ) , .B1( u2_u8_u0_n151 ) , .ZN( u2_u8_u0_n152 ) , .A( u2_u8_u0_n158 ) );
  AOI21_X1 u2_u8_u0_U47 (.A( u2_u8_u0_n147 ) , .B2( u2_u8_u0_n148 ) , .B1( u2_u8_u0_n149 ) , .ZN( u2_u8_u0_n153 ) );
  INV_X1 u2_u8_u0_U48 (.ZN( u2_u8_u0_n171 ) , .A( u2_u8_u0_n99 ) );
  OAI211_X1 u2_u8_u0_U49 (.C2( u2_u8_u0_n140 ) , .C1( u2_u8_u0_n161 ) , .A( u2_u8_u0_n169 ) , .B( u2_u8_u0_n98 ) , .ZN( u2_u8_u0_n99 ) );
  AOI21_X1 u2_u8_u0_U5 (.B2( u2_u8_u0_n131 ) , .ZN( u2_u8_u0_n134 ) , .B1( u2_u8_u0_n151 ) , .A( u2_u8_u0_n158 ) );
  INV_X1 u2_u8_u0_U50 (.ZN( u2_u8_u0_n169 ) , .A( u2_u8_u0_n91 ) );
  AOI211_X1 u2_u8_u0_U51 (.C1( u2_u8_u0_n118 ) , .A( u2_u8_u0_n123 ) , .B( u2_u8_u0_n96 ) , .C2( u2_u8_u0_n97 ) , .ZN( u2_u8_u0_n98 ) );
  NOR2_X1 u2_u8_u0_U52 (.A2( u2_u8_X_4 ) , .A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n118 ) );
  NOR2_X1 u2_u8_u0_U53 (.A2( u2_u8_X_1 ) , .ZN( u2_u8_u0_n101 ) , .A1( u2_u8_u0_n163 ) );
  NOR2_X1 u2_u8_u0_U54 (.A2( u2_u8_X_3 ) , .A1( u2_u8_X_6 ) , .ZN( u2_u8_u0_n94 ) );
  NOR2_X1 u2_u8_u0_U55 (.A2( u2_u8_X_6 ) , .ZN( u2_u8_u0_n100 ) , .A1( u2_u8_u0_n162 ) );
  NAND2_X1 u2_u8_u0_U56 (.A2( u2_u8_X_4 ) , .A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n144 ) );
  NOR2_X1 u2_u8_u0_U57 (.A2( u2_u8_X_5 ) , .ZN( u2_u8_u0_n136 ) , .A1( u2_u8_u0_n159 ) );
  NAND2_X1 u2_u8_u0_U58 (.A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n138 ) , .A2( u2_u8_u0_n159 ) );
  AND2_X1 u2_u8_u0_U59 (.A2( u2_u8_X_3 ) , .A1( u2_u8_X_6 ) , .ZN( u2_u8_u0_n102 ) );
  NOR2_X1 u2_u8_u0_U6 (.A1( u2_u8_u0_n108 ) , .ZN( u2_u8_u0_n123 ) , .A2( u2_u8_u0_n158 ) );
  AND2_X1 u2_u8_u0_U60 (.A1( u2_u8_X_6 ) , .A2( u2_u8_u0_n162 ) , .ZN( u2_u8_u0_n93 ) );
  INV_X1 u2_u8_u0_U61 (.A( u2_u8_X_4 ) , .ZN( u2_u8_u0_n159 ) );
  INV_X1 u2_u8_u0_U62 (.A( u2_u8_X_1 ) , .ZN( u2_u8_u0_n164 ) );
  INV_X1 u2_u8_u0_U63 (.A( u2_u8_X_3 ) , .ZN( u2_u8_u0_n162 ) );
  INV_X1 u2_u8_u0_U64 (.A( u2_u8_u0_n126 ) , .ZN( u2_u8_u0_n168 ) );
  AOI211_X1 u2_u8_u0_U65 (.B( u2_u8_u0_n133 ) , .A( u2_u8_u0_n134 ) , .C2( u2_u8_u0_n135 ) , .C1( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n137 ) );
  OR4_X1 u2_u8_u0_U66 (.ZN( u2_out8_17 ) , .A4( u2_u8_u0_n122 ) , .A2( u2_u8_u0_n123 ) , .A1( u2_u8_u0_n124 ) , .A3( u2_u8_u0_n170 ) );
  AOI21_X1 u2_u8_u0_U67 (.B2( u2_u8_u0_n107 ) , .ZN( u2_u8_u0_n124 ) , .B1( u2_u8_u0_n128 ) , .A( u2_u8_u0_n161 ) );
  INV_X1 u2_u8_u0_U68 (.A( u2_u8_u0_n111 ) , .ZN( u2_u8_u0_n170 ) );
  OR4_X1 u2_u8_u0_U69 (.ZN( u2_out8_31 ) , .A4( u2_u8_u0_n155 ) , .A2( u2_u8_u0_n156 ) , .A1( u2_u8_u0_n157 ) , .A3( u2_u8_u0_n173 ) );
  OAI21_X1 u2_u8_u0_U7 (.B1( u2_u8_u0_n150 ) , .B2( u2_u8_u0_n158 ) , .A( u2_u8_u0_n172 ) , .ZN( u2_u8_u0_n89 ) );
  AOI21_X1 u2_u8_u0_U70 (.A( u2_u8_u0_n138 ) , .B2( u2_u8_u0_n139 ) , .B1( u2_u8_u0_n140 ) , .ZN( u2_u8_u0_n157 ) );
  AOI211_X1 u2_u8_u0_U71 (.B( u2_u8_u0_n104 ) , .A( u2_u8_u0_n105 ) , .ZN( u2_u8_u0_n106 ) , .C2( u2_u8_u0_n113 ) , .C1( u2_u8_u0_n160 ) );
  INV_X1 u2_u8_u0_U72 (.ZN( u2_u8_u0_n174 ) , .A( u2_u8_u0_n89 ) );
  INV_X1 u2_u8_u0_U73 (.A( u2_u8_u0_n142 ) , .ZN( u2_u8_u0_n165 ) );
  AOI21_X1 u2_u8_u0_U74 (.ZN( u2_u8_u0_n116 ) , .B2( u2_u8_u0_n142 ) , .A( u2_u8_u0_n144 ) , .B1( u2_u8_u0_n166 ) );
  AOI21_X1 u2_u8_u0_U75 (.B2( u2_u8_u0_n141 ) , .B1( u2_u8_u0_n142 ) , .ZN( u2_u8_u0_n156 ) , .A( u2_u8_u0_n161 ) );
  OAI221_X1 u2_u8_u0_U76 (.C1( u2_u8_u0_n121 ) , .ZN( u2_u8_u0_n122 ) , .B2( u2_u8_u0_n127 ) , .A( u2_u8_u0_n143 ) , .B1( u2_u8_u0_n144 ) , .C2( u2_u8_u0_n147 ) );
  AOI21_X1 u2_u8_u0_U77 (.B1( u2_u8_u0_n132 ) , .ZN( u2_u8_u0_n133 ) , .A( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n166 ) );
  OAI22_X1 u2_u8_u0_U78 (.ZN( u2_u8_u0_n105 ) , .A2( u2_u8_u0_n132 ) , .B1( u2_u8_u0_n146 ) , .A1( u2_u8_u0_n147 ) , .B2( u2_u8_u0_n161 ) );
  NAND2_X1 u2_u8_u0_U79 (.ZN( u2_u8_u0_n110 ) , .A2( u2_u8_u0_n132 ) , .A1( u2_u8_u0_n145 ) );
  AND2_X1 u2_u8_u0_U8 (.A1( u2_u8_u0_n114 ) , .A2( u2_u8_u0_n121 ) , .ZN( u2_u8_u0_n146 ) );
  INV_X1 u2_u8_u0_U80 (.A( u2_u8_u0_n119 ) , .ZN( u2_u8_u0_n167 ) );
  NAND2_X1 u2_u8_u0_U81 (.ZN( u2_u8_u0_n148 ) , .A1( u2_u8_u0_n93 ) , .A2( u2_u8_u0_n95 ) );
  NAND2_X1 u2_u8_u0_U82 (.A1( u2_u8_u0_n100 ) , .ZN( u2_u8_u0_n129 ) , .A2( u2_u8_u0_n95 ) );
  NAND2_X1 u2_u8_u0_U83 (.A1( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n128 ) , .A2( u2_u8_u0_n95 ) );
  NOR2_X1 u2_u8_u0_U84 (.A2( u2_u8_X_1 ) , .A1( u2_u8_X_2 ) , .ZN( u2_u8_u0_n92 ) );
  NAND2_X1 u2_u8_u0_U85 (.ZN( u2_u8_u0_n142 ) , .A1( u2_u8_u0_n94 ) , .A2( u2_u8_u0_n95 ) );
  NOR2_X1 u2_u8_u0_U86 (.A2( u2_u8_X_2 ) , .ZN( u2_u8_u0_n103 ) , .A1( u2_u8_u0_n164 ) );
  INV_X1 u2_u8_u0_U87 (.A( u2_u8_X_2 ) , .ZN( u2_u8_u0_n163 ) );
  NAND3_X1 u2_u8_u0_U88 (.ZN( u2_out8_23 ) , .A3( u2_u8_u0_n137 ) , .A1( u2_u8_u0_n168 ) , .A2( u2_u8_u0_n171 ) );
  NAND3_X1 u2_u8_u0_U89 (.A3( u2_u8_u0_n127 ) , .A2( u2_u8_u0_n128 ) , .ZN( u2_u8_u0_n135 ) , .A1( u2_u8_u0_n150 ) );
  NAND2_X1 u2_u8_u0_U9 (.ZN( u2_u8_u0_n113 ) , .A1( u2_u8_u0_n139 ) , .A2( u2_u8_u0_n149 ) );
  NAND3_X1 u2_u8_u0_U90 (.ZN( u2_u8_u0_n117 ) , .A3( u2_u8_u0_n132 ) , .A2( u2_u8_u0_n139 ) , .A1( u2_u8_u0_n148 ) );
  NAND3_X1 u2_u8_u0_U91 (.ZN( u2_u8_u0_n109 ) , .A2( u2_u8_u0_n114 ) , .A3( u2_u8_u0_n140 ) , .A1( u2_u8_u0_n149 ) );
  NAND3_X1 u2_u8_u0_U92 (.ZN( u2_out8_9 ) , .A3( u2_u8_u0_n106 ) , .A2( u2_u8_u0_n171 ) , .A1( u2_u8_u0_n174 ) );
  NAND3_X1 u2_u8_u0_U93 (.A2( u2_u8_u0_n128 ) , .A1( u2_u8_u0_n132 ) , .A3( u2_u8_u0_n146 ) , .ZN( u2_u8_u0_n97 ) );
  AOI21_X1 u2_u8_u1_U10 (.B2( u2_u8_u1_n155 ) , .B1( u2_u8_u1_n156 ) , .ZN( u2_u8_u1_n157 ) , .A( u2_u8_u1_n174 ) );
  NAND3_X1 u2_u8_u1_U100 (.ZN( u2_u8_u1_n113 ) , .A1( u2_u8_u1_n120 ) , .A3( u2_u8_u1_n133 ) , .A2( u2_u8_u1_n155 ) );
  NAND2_X1 u2_u8_u1_U11 (.ZN( u2_u8_u1_n140 ) , .A2( u2_u8_u1_n150 ) , .A1( u2_u8_u1_n155 ) );
  NAND2_X1 u2_u8_u1_U12 (.A1( u2_u8_u1_n131 ) , .ZN( u2_u8_u1_n147 ) , .A2( u2_u8_u1_n153 ) );
  AOI22_X1 u2_u8_u1_U13 (.B2( u2_u8_u1_n136 ) , .A2( u2_u8_u1_n137 ) , .ZN( u2_u8_u1_n143 ) , .A1( u2_u8_u1_n171 ) , .B1( u2_u8_u1_n173 ) );
  INV_X1 u2_u8_u1_U14 (.A( u2_u8_u1_n147 ) , .ZN( u2_u8_u1_n181 ) );
  INV_X1 u2_u8_u1_U15 (.A( u2_u8_u1_n139 ) , .ZN( u2_u8_u1_n174 ) );
  OR4_X1 u2_u8_u1_U16 (.A4( u2_u8_u1_n106 ) , .A3( u2_u8_u1_n107 ) , .ZN( u2_u8_u1_n108 ) , .A1( u2_u8_u1_n117 ) , .A2( u2_u8_u1_n184 ) );
  AOI21_X1 u2_u8_u1_U17 (.ZN( u2_u8_u1_n106 ) , .A( u2_u8_u1_n112 ) , .B1( u2_u8_u1_n154 ) , .B2( u2_u8_u1_n156 ) );
  AOI21_X1 u2_u8_u1_U18 (.ZN( u2_u8_u1_n107 ) , .B1( u2_u8_u1_n134 ) , .B2( u2_u8_u1_n149 ) , .A( u2_u8_u1_n174 ) );
  INV_X1 u2_u8_u1_U19 (.A( u2_u8_u1_n101 ) , .ZN( u2_u8_u1_n184 ) );
  INV_X1 u2_u8_u1_U20 (.A( u2_u8_u1_n112 ) , .ZN( u2_u8_u1_n171 ) );
  NAND2_X1 u2_u8_u1_U21 (.ZN( u2_u8_u1_n141 ) , .A1( u2_u8_u1_n153 ) , .A2( u2_u8_u1_n156 ) );
  AND2_X1 u2_u8_u1_U22 (.A1( u2_u8_u1_n123 ) , .ZN( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n161 ) );
  NAND2_X1 u2_u8_u1_U23 (.A2( u2_u8_u1_n115 ) , .A1( u2_u8_u1_n116 ) , .ZN( u2_u8_u1_n148 ) );
  NAND2_X1 u2_u8_u1_U24 (.A2( u2_u8_u1_n133 ) , .A1( u2_u8_u1_n135 ) , .ZN( u2_u8_u1_n159 ) );
  NAND2_X1 u2_u8_u1_U25 (.A2( u2_u8_u1_n115 ) , .A1( u2_u8_u1_n120 ) , .ZN( u2_u8_u1_n132 ) );
  INV_X1 u2_u8_u1_U26 (.A( u2_u8_u1_n154 ) , .ZN( u2_u8_u1_n178 ) );
  INV_X1 u2_u8_u1_U27 (.A( u2_u8_u1_n151 ) , .ZN( u2_u8_u1_n183 ) );
  AND2_X1 u2_u8_u1_U28 (.A1( u2_u8_u1_n129 ) , .A2( u2_u8_u1_n133 ) , .ZN( u2_u8_u1_n149 ) );
  INV_X1 u2_u8_u1_U29 (.A( u2_u8_u1_n131 ) , .ZN( u2_u8_u1_n180 ) );
  INV_X1 u2_u8_u1_U3 (.A( u2_u8_u1_n159 ) , .ZN( u2_u8_u1_n182 ) );
  AOI221_X1 u2_u8_u1_U30 (.B1( u2_u8_u1_n140 ) , .ZN( u2_u8_u1_n167 ) , .B2( u2_u8_u1_n172 ) , .C2( u2_u8_u1_n175 ) , .C1( u2_u8_u1_n178 ) , .A( u2_u8_u1_n188 ) );
  INV_X1 u2_u8_u1_U31 (.ZN( u2_u8_u1_n188 ) , .A( u2_u8_u1_n97 ) );
  AOI211_X1 u2_u8_u1_U32 (.A( u2_u8_u1_n118 ) , .C1( u2_u8_u1_n132 ) , .C2( u2_u8_u1_n139 ) , .B( u2_u8_u1_n96 ) , .ZN( u2_u8_u1_n97 ) );
  AOI21_X1 u2_u8_u1_U33 (.B2( u2_u8_u1_n121 ) , .B1( u2_u8_u1_n135 ) , .A( u2_u8_u1_n152 ) , .ZN( u2_u8_u1_n96 ) );
  OAI221_X1 u2_u8_u1_U34 (.A( u2_u8_u1_n119 ) , .C2( u2_u8_u1_n129 ) , .ZN( u2_u8_u1_n138 ) , .B2( u2_u8_u1_n152 ) , .C1( u2_u8_u1_n174 ) , .B1( u2_u8_u1_n187 ) );
  INV_X1 u2_u8_u1_U35 (.A( u2_u8_u1_n148 ) , .ZN( u2_u8_u1_n187 ) );
  AOI211_X1 u2_u8_u1_U36 (.B( u2_u8_u1_n117 ) , .A( u2_u8_u1_n118 ) , .ZN( u2_u8_u1_n119 ) , .C2( u2_u8_u1_n146 ) , .C1( u2_u8_u1_n159 ) );
  NOR2_X1 u2_u8_u1_U37 (.A1( u2_u8_u1_n168 ) , .A2( u2_u8_u1_n176 ) , .ZN( u2_u8_u1_n98 ) );
  AOI211_X1 u2_u8_u1_U38 (.B( u2_u8_u1_n162 ) , .A( u2_u8_u1_n163 ) , .C2( u2_u8_u1_n164 ) , .ZN( u2_u8_u1_n165 ) , .C1( u2_u8_u1_n171 ) );
  AOI21_X1 u2_u8_u1_U39 (.A( u2_u8_u1_n160 ) , .B2( u2_u8_u1_n161 ) , .ZN( u2_u8_u1_n162 ) , .B1( u2_u8_u1_n182 ) );
  AOI221_X1 u2_u8_u1_U4 (.A( u2_u8_u1_n138 ) , .C2( u2_u8_u1_n139 ) , .C1( u2_u8_u1_n140 ) , .B2( u2_u8_u1_n141 ) , .ZN( u2_u8_u1_n142 ) , .B1( u2_u8_u1_n175 ) );
  OR2_X1 u2_u8_u1_U40 (.A2( u2_u8_u1_n157 ) , .A1( u2_u8_u1_n158 ) , .ZN( u2_u8_u1_n163 ) );
  NAND2_X1 u2_u8_u1_U41 (.A1( u2_u8_u1_n128 ) , .ZN( u2_u8_u1_n146 ) , .A2( u2_u8_u1_n160 ) );
  NAND2_X1 u2_u8_u1_U42 (.A2( u2_u8_u1_n112 ) , .ZN( u2_u8_u1_n139 ) , .A1( u2_u8_u1_n152 ) );
  NAND2_X1 u2_u8_u1_U43 (.A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n156 ) , .A2( u2_u8_u1_n99 ) );
  NOR2_X1 u2_u8_u1_U44 (.ZN( u2_u8_u1_n117 ) , .A1( u2_u8_u1_n121 ) , .A2( u2_u8_u1_n160 ) );
  OAI21_X1 u2_u8_u1_U45 (.B2( u2_u8_u1_n123 ) , .ZN( u2_u8_u1_n145 ) , .B1( u2_u8_u1_n160 ) , .A( u2_u8_u1_n185 ) );
  INV_X1 u2_u8_u1_U46 (.A( u2_u8_u1_n122 ) , .ZN( u2_u8_u1_n185 ) );
  AOI21_X1 u2_u8_u1_U47 (.B2( u2_u8_u1_n120 ) , .B1( u2_u8_u1_n121 ) , .ZN( u2_u8_u1_n122 ) , .A( u2_u8_u1_n128 ) );
  AOI21_X1 u2_u8_u1_U48 (.A( u2_u8_u1_n128 ) , .B2( u2_u8_u1_n129 ) , .ZN( u2_u8_u1_n130 ) , .B1( u2_u8_u1_n150 ) );
  NAND2_X1 u2_u8_u1_U49 (.ZN( u2_u8_u1_n112 ) , .A1( u2_u8_u1_n169 ) , .A2( u2_u8_u1_n170 ) );
  AOI211_X1 u2_u8_u1_U5 (.ZN( u2_u8_u1_n124 ) , .A( u2_u8_u1_n138 ) , .C2( u2_u8_u1_n139 ) , .B( u2_u8_u1_n145 ) , .C1( u2_u8_u1_n147 ) );
  NAND2_X1 u2_u8_u1_U50 (.ZN( u2_u8_u1_n129 ) , .A2( u2_u8_u1_n95 ) , .A1( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U51 (.A1( u2_u8_u1_n102 ) , .ZN( u2_u8_u1_n154 ) , .A2( u2_u8_u1_n99 ) );
  NAND2_X1 u2_u8_u1_U52 (.A2( u2_u8_u1_n100 ) , .ZN( u2_u8_u1_n135 ) , .A1( u2_u8_u1_n99 ) );
  AOI21_X1 u2_u8_u1_U53 (.A( u2_u8_u1_n152 ) , .B2( u2_u8_u1_n153 ) , .B1( u2_u8_u1_n154 ) , .ZN( u2_u8_u1_n158 ) );
  INV_X1 u2_u8_u1_U54 (.A( u2_u8_u1_n160 ) , .ZN( u2_u8_u1_n175 ) );
  NAND2_X1 u2_u8_u1_U55 (.A1( u2_u8_u1_n100 ) , .ZN( u2_u8_u1_n116 ) , .A2( u2_u8_u1_n95 ) );
  NAND2_X1 u2_u8_u1_U56 (.A1( u2_u8_u1_n102 ) , .ZN( u2_u8_u1_n131 ) , .A2( u2_u8_u1_n95 ) );
  NAND2_X1 u2_u8_u1_U57 (.A2( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n121 ) , .A1( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U58 (.A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n153 ) , .A2( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U59 (.A2( u2_u8_u1_n104 ) , .A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n133 ) );
  AOI22_X1 u2_u8_u1_U6 (.B2( u2_u8_u1_n113 ) , .A2( u2_u8_u1_n114 ) , .ZN( u2_u8_u1_n125 ) , .A1( u2_u8_u1_n171 ) , .B1( u2_u8_u1_n173 ) );
  NAND2_X1 u2_u8_u1_U60 (.ZN( u2_u8_u1_n150 ) , .A2( u2_u8_u1_n98 ) , .A1( u2_u8_u1_n99 ) );
  NAND2_X1 u2_u8_u1_U61 (.A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n155 ) , .A2( u2_u8_u1_n95 ) );
  OAI21_X1 u2_u8_u1_U62 (.ZN( u2_u8_u1_n109 ) , .B1( u2_u8_u1_n129 ) , .B2( u2_u8_u1_n160 ) , .A( u2_u8_u1_n167 ) );
  NAND2_X1 u2_u8_u1_U63 (.A2( u2_u8_u1_n100 ) , .A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n120 ) );
  NAND2_X1 u2_u8_u1_U64 (.A1( u2_u8_u1_n102 ) , .A2( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n115 ) );
  NAND2_X1 u2_u8_u1_U65 (.A2( u2_u8_u1_n100 ) , .A1( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n151 ) );
  NAND2_X1 u2_u8_u1_U66 (.A2( u2_u8_u1_n103 ) , .A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n161 ) );
  INV_X1 u2_u8_u1_U67 (.A( u2_u8_u1_n152 ) , .ZN( u2_u8_u1_n173 ) );
  INV_X1 u2_u8_u1_U68 (.A( u2_u8_u1_n128 ) , .ZN( u2_u8_u1_n172 ) );
  NAND2_X1 u2_u8_u1_U69 (.A2( u2_u8_u1_n102 ) , .A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n123 ) );
  NAND2_X1 u2_u8_u1_U7 (.ZN( u2_u8_u1_n114 ) , .A1( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n156 ) );
  NOR2_X1 u2_u8_u1_U70 (.A2( u2_u8_X_7 ) , .A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n95 ) );
  NOR2_X1 u2_u8_u1_U71 (.A1( u2_u8_X_12 ) , .A2( u2_u8_X_9 ) , .ZN( u2_u8_u1_n100 ) );
  NOR2_X1 u2_u8_u1_U72 (.A2( u2_u8_X_8 ) , .A1( u2_u8_u1_n177 ) , .ZN( u2_u8_u1_n99 ) );
  NOR2_X1 u2_u8_u1_U73 (.A2( u2_u8_X_12 ) , .ZN( u2_u8_u1_n102 ) , .A1( u2_u8_u1_n176 ) );
  NOR2_X1 u2_u8_u1_U74 (.A2( u2_u8_X_9 ) , .ZN( u2_u8_u1_n105 ) , .A1( u2_u8_u1_n168 ) );
  NAND2_X1 u2_u8_u1_U75 (.A1( u2_u8_X_10 ) , .ZN( u2_u8_u1_n160 ) , .A2( u2_u8_u1_n169 ) );
  NAND2_X1 u2_u8_u1_U76 (.A2( u2_u8_X_10 ) , .A1( u2_u8_X_11 ) , .ZN( u2_u8_u1_n152 ) );
  NAND2_X1 u2_u8_u1_U77 (.A1( u2_u8_X_11 ) , .ZN( u2_u8_u1_n128 ) , .A2( u2_u8_u1_n170 ) );
  AND2_X1 u2_u8_u1_U78 (.A2( u2_u8_X_7 ) , .A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n104 ) );
  AND2_X1 u2_u8_u1_U79 (.A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n103 ) , .A2( u2_u8_u1_n177 ) );
  NOR2_X1 u2_u8_u1_U8 (.A1( u2_u8_u1_n112 ) , .A2( u2_u8_u1_n116 ) , .ZN( u2_u8_u1_n118 ) );
  INV_X1 u2_u8_u1_U80 (.A( u2_u8_X_10 ) , .ZN( u2_u8_u1_n170 ) );
  INV_X1 u2_u8_u1_U81 (.A( u2_u8_X_9 ) , .ZN( u2_u8_u1_n176 ) );
  INV_X1 u2_u8_u1_U82 (.A( u2_u8_X_11 ) , .ZN( u2_u8_u1_n169 ) );
  INV_X1 u2_u8_u1_U83 (.A( u2_u8_X_12 ) , .ZN( u2_u8_u1_n168 ) );
  INV_X1 u2_u8_u1_U84 (.A( u2_u8_X_7 ) , .ZN( u2_u8_u1_n177 ) );
  NAND4_X1 u2_u8_u1_U85 (.ZN( u2_out8_28 ) , .A4( u2_u8_u1_n124 ) , .A3( u2_u8_u1_n125 ) , .A2( u2_u8_u1_n126 ) , .A1( u2_u8_u1_n127 ) );
  OAI21_X1 u2_u8_u1_U86 (.ZN( u2_u8_u1_n127 ) , .B2( u2_u8_u1_n139 ) , .B1( u2_u8_u1_n175 ) , .A( u2_u8_u1_n183 ) );
  OAI21_X1 u2_u8_u1_U87 (.ZN( u2_u8_u1_n126 ) , .B2( u2_u8_u1_n140 ) , .A( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n178 ) );
  NAND4_X1 u2_u8_u1_U88 (.ZN( u2_out8_18 ) , .A4( u2_u8_u1_n165 ) , .A3( u2_u8_u1_n166 ) , .A1( u2_u8_u1_n167 ) , .A2( u2_u8_u1_n186 ) );
  AOI22_X1 u2_u8_u1_U89 (.B2( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n147 ) , .A2( u2_u8_u1_n148 ) , .ZN( u2_u8_u1_n166 ) , .A1( u2_u8_u1_n172 ) );
  OAI21_X1 u2_u8_u1_U9 (.ZN( u2_u8_u1_n101 ) , .B1( u2_u8_u1_n141 ) , .A( u2_u8_u1_n146 ) , .B2( u2_u8_u1_n183 ) );
  INV_X1 u2_u8_u1_U90 (.A( u2_u8_u1_n145 ) , .ZN( u2_u8_u1_n186 ) );
  NAND4_X1 u2_u8_u1_U91 (.ZN( u2_out8_2 ) , .A4( u2_u8_u1_n142 ) , .A3( u2_u8_u1_n143 ) , .A2( u2_u8_u1_n144 ) , .A1( u2_u8_u1_n179 ) );
  OAI21_X1 u2_u8_u1_U92 (.B2( u2_u8_u1_n132 ) , .ZN( u2_u8_u1_n144 ) , .A( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n180 ) );
  INV_X1 u2_u8_u1_U93 (.A( u2_u8_u1_n130 ) , .ZN( u2_u8_u1_n179 ) );
  OR4_X1 u2_u8_u1_U94 (.ZN( u2_out8_13 ) , .A4( u2_u8_u1_n108 ) , .A3( u2_u8_u1_n109 ) , .A2( u2_u8_u1_n110 ) , .A1( u2_u8_u1_n111 ) );
  AOI21_X1 u2_u8_u1_U95 (.ZN( u2_u8_u1_n111 ) , .A( u2_u8_u1_n128 ) , .B2( u2_u8_u1_n131 ) , .B1( u2_u8_u1_n135 ) );
  AOI21_X1 u2_u8_u1_U96 (.ZN( u2_u8_u1_n110 ) , .A( u2_u8_u1_n116 ) , .B1( u2_u8_u1_n152 ) , .B2( u2_u8_u1_n160 ) );
  NAND3_X1 u2_u8_u1_U97 (.A3( u2_u8_u1_n149 ) , .A2( u2_u8_u1_n150 ) , .A1( u2_u8_u1_n151 ) , .ZN( u2_u8_u1_n164 ) );
  NAND3_X1 u2_u8_u1_U98 (.A3( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n135 ) , .ZN( u2_u8_u1_n136 ) , .A1( u2_u8_u1_n151 ) );
  NAND3_X1 u2_u8_u1_U99 (.A1( u2_u8_u1_n133 ) , .ZN( u2_u8_u1_n137 ) , .A2( u2_u8_u1_n154 ) , .A3( u2_u8_u1_n181 ) );
  OAI22_X1 u2_u8_u2_U10 (.B1( u2_u8_u2_n151 ) , .A2( u2_u8_u2_n152 ) , .A1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n160 ) , .B2( u2_u8_u2_n168 ) );
  NAND3_X1 u2_u8_u2_U100 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n98 ) );
  NOR3_X1 u2_u8_u2_U11 (.A1( u2_u8_u2_n150 ) , .ZN( u2_u8_u2_n151 ) , .A3( u2_u8_u2_n175 ) , .A2( u2_u8_u2_n188 ) );
  AOI21_X1 u2_u8_u2_U12 (.B2( u2_u8_u2_n123 ) , .ZN( u2_u8_u2_n125 ) , .A( u2_u8_u2_n171 ) , .B1( u2_u8_u2_n184 ) );
  INV_X1 u2_u8_u2_U13 (.A( u2_u8_u2_n150 ) , .ZN( u2_u8_u2_n184 ) );
  AOI21_X1 u2_u8_u2_U14 (.ZN( u2_u8_u2_n144 ) , .B2( u2_u8_u2_n155 ) , .A( u2_u8_u2_n172 ) , .B1( u2_u8_u2_n185 ) );
  AOI21_X1 u2_u8_u2_U15 (.B2( u2_u8_u2_n143 ) , .ZN( u2_u8_u2_n145 ) , .B1( u2_u8_u2_n152 ) , .A( u2_u8_u2_n171 ) );
  INV_X1 u2_u8_u2_U16 (.A( u2_u8_u2_n156 ) , .ZN( u2_u8_u2_n171 ) );
  INV_X1 u2_u8_u2_U17 (.A( u2_u8_u2_n120 ) , .ZN( u2_u8_u2_n188 ) );
  NAND2_X1 u2_u8_u2_U18 (.A2( u2_u8_u2_n122 ) , .ZN( u2_u8_u2_n150 ) , .A1( u2_u8_u2_n152 ) );
  INV_X1 u2_u8_u2_U19 (.A( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n170 ) );
  INV_X1 u2_u8_u2_U20 (.A( u2_u8_u2_n137 ) , .ZN( u2_u8_u2_n173 ) );
  NAND2_X1 u2_u8_u2_U21 (.A1( u2_u8_u2_n132 ) , .A2( u2_u8_u2_n139 ) , .ZN( u2_u8_u2_n157 ) );
  INV_X1 u2_u8_u2_U22 (.A( u2_u8_u2_n113 ) , .ZN( u2_u8_u2_n178 ) );
  INV_X1 u2_u8_u2_U23 (.A( u2_u8_u2_n139 ) , .ZN( u2_u8_u2_n175 ) );
  INV_X1 u2_u8_u2_U24 (.A( u2_u8_u2_n155 ) , .ZN( u2_u8_u2_n181 ) );
  INV_X1 u2_u8_u2_U25 (.A( u2_u8_u2_n119 ) , .ZN( u2_u8_u2_n177 ) );
  INV_X1 u2_u8_u2_U26 (.A( u2_u8_u2_n116 ) , .ZN( u2_u8_u2_n180 ) );
  INV_X1 u2_u8_u2_U27 (.A( u2_u8_u2_n131 ) , .ZN( u2_u8_u2_n179 ) );
  INV_X1 u2_u8_u2_U28 (.A( u2_u8_u2_n154 ) , .ZN( u2_u8_u2_n176 ) );
  NAND2_X1 u2_u8_u2_U29 (.A2( u2_u8_u2_n116 ) , .A1( u2_u8_u2_n117 ) , .ZN( u2_u8_u2_n118 ) );
  NOR2_X1 u2_u8_u2_U3 (.ZN( u2_u8_u2_n121 ) , .A2( u2_u8_u2_n177 ) , .A1( u2_u8_u2_n180 ) );
  INV_X1 u2_u8_u2_U30 (.A( u2_u8_u2_n132 ) , .ZN( u2_u8_u2_n182 ) );
  INV_X1 u2_u8_u2_U31 (.A( u2_u8_u2_n158 ) , .ZN( u2_u8_u2_n183 ) );
  OAI21_X1 u2_u8_u2_U32 (.A( u2_u8_u2_n156 ) , .B1( u2_u8_u2_n157 ) , .ZN( u2_u8_u2_n158 ) , .B2( u2_u8_u2_n179 ) );
  NOR2_X1 u2_u8_u2_U33 (.ZN( u2_u8_u2_n156 ) , .A1( u2_u8_u2_n166 ) , .A2( u2_u8_u2_n169 ) );
  NOR2_X1 u2_u8_u2_U34 (.A2( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n137 ) , .A1( u2_u8_u2_n140 ) );
  NOR2_X1 u2_u8_u2_U35 (.A2( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n153 ) , .A1( u2_u8_u2_n156 ) );
  AOI211_X1 u2_u8_u2_U36 (.ZN( u2_u8_u2_n130 ) , .C1( u2_u8_u2_n138 ) , .C2( u2_u8_u2_n179 ) , .B( u2_u8_u2_n96 ) , .A( u2_u8_u2_n97 ) );
  OAI22_X1 u2_u8_u2_U37 (.B1( u2_u8_u2_n133 ) , .A2( u2_u8_u2_n137 ) , .A1( u2_u8_u2_n152 ) , .B2( u2_u8_u2_n168 ) , .ZN( u2_u8_u2_n97 ) );
  OAI221_X1 u2_u8_u2_U38 (.B1( u2_u8_u2_n113 ) , .C1( u2_u8_u2_n132 ) , .A( u2_u8_u2_n149 ) , .B2( u2_u8_u2_n171 ) , .C2( u2_u8_u2_n172 ) , .ZN( u2_u8_u2_n96 ) );
  OAI221_X1 u2_u8_u2_U39 (.A( u2_u8_u2_n115 ) , .C2( u2_u8_u2_n123 ) , .B2( u2_u8_u2_n143 ) , .B1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n163 ) , .C1( u2_u8_u2_n168 ) );
  INV_X1 u2_u8_u2_U4 (.A( u2_u8_u2_n134 ) , .ZN( u2_u8_u2_n185 ) );
  OAI21_X1 u2_u8_u2_U40 (.A( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n115 ) , .B1( u2_u8_u2_n176 ) , .B2( u2_u8_u2_n178 ) );
  OAI221_X1 u2_u8_u2_U41 (.A( u2_u8_u2_n135 ) , .B2( u2_u8_u2_n136 ) , .B1( u2_u8_u2_n137 ) , .ZN( u2_u8_u2_n162 ) , .C2( u2_u8_u2_n167 ) , .C1( u2_u8_u2_n185 ) );
  AND3_X1 u2_u8_u2_U42 (.A3( u2_u8_u2_n131 ) , .A2( u2_u8_u2_n132 ) , .A1( u2_u8_u2_n133 ) , .ZN( u2_u8_u2_n136 ) );
  AOI22_X1 u2_u8_u2_U43 (.ZN( u2_u8_u2_n135 ) , .B1( u2_u8_u2_n140 ) , .A1( u2_u8_u2_n156 ) , .B2( u2_u8_u2_n180 ) , .A2( u2_u8_u2_n188 ) );
  AOI21_X1 u2_u8_u2_U44 (.ZN( u2_u8_u2_n149 ) , .B1( u2_u8_u2_n173 ) , .B2( u2_u8_u2_n188 ) , .A( u2_u8_u2_n95 ) );
  AND3_X1 u2_u8_u2_U45 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n156 ) , .ZN( u2_u8_u2_n95 ) );
  OAI21_X1 u2_u8_u2_U46 (.A( u2_u8_u2_n141 ) , .B2( u2_u8_u2_n142 ) , .ZN( u2_u8_u2_n146 ) , .B1( u2_u8_u2_n153 ) );
  OAI21_X1 u2_u8_u2_U47 (.A( u2_u8_u2_n140 ) , .ZN( u2_u8_u2_n141 ) , .B1( u2_u8_u2_n176 ) , .B2( u2_u8_u2_n177 ) );
  NOR3_X1 u2_u8_u2_U48 (.ZN( u2_u8_u2_n142 ) , .A3( u2_u8_u2_n175 ) , .A2( u2_u8_u2_n178 ) , .A1( u2_u8_u2_n181 ) );
  OAI21_X1 u2_u8_u2_U49 (.A( u2_u8_u2_n101 ) , .B2( u2_u8_u2_n121 ) , .B1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n164 ) );
  NOR4_X1 u2_u8_u2_U5 (.A4( u2_u8_u2_n124 ) , .A3( u2_u8_u2_n125 ) , .A2( u2_u8_u2_n126 ) , .A1( u2_u8_u2_n127 ) , .ZN( u2_u8_u2_n128 ) );
  NAND2_X1 u2_u8_u2_U50 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n155 ) );
  NAND2_X1 u2_u8_u2_U51 (.A2( u2_u8_u2_n105 ) , .A1( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n143 ) );
  NAND2_X1 u2_u8_u2_U52 (.A1( u2_u8_u2_n104 ) , .A2( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n152 ) );
  NAND2_X1 u2_u8_u2_U53 (.A1( u2_u8_u2_n100 ) , .A2( u2_u8_u2_n105 ) , .ZN( u2_u8_u2_n132 ) );
  INV_X1 u2_u8_u2_U54 (.A( u2_u8_u2_n140 ) , .ZN( u2_u8_u2_n168 ) );
  INV_X1 u2_u8_u2_U55 (.A( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n167 ) );
  NAND2_X1 u2_u8_u2_U56 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n113 ) );
  NAND2_X1 u2_u8_u2_U57 (.A1( u2_u8_u2_n106 ) , .A2( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n131 ) );
  NAND2_X1 u2_u8_u2_U58 (.A1( u2_u8_u2_n103 ) , .A2( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n139 ) );
  NAND2_X1 u2_u8_u2_U59 (.A1( u2_u8_u2_n103 ) , .A2( u2_u8_u2_n105 ) , .ZN( u2_u8_u2_n133 ) );
  AOI21_X1 u2_u8_u2_U6 (.B2( u2_u8_u2_n119 ) , .ZN( u2_u8_u2_n127 ) , .A( u2_u8_u2_n137 ) , .B1( u2_u8_u2_n155 ) );
  NAND2_X1 u2_u8_u2_U60 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n103 ) , .ZN( u2_u8_u2_n154 ) );
  NAND2_X1 u2_u8_u2_U61 (.A2( u2_u8_u2_n103 ) , .A1( u2_u8_u2_n104 ) , .ZN( u2_u8_u2_n119 ) );
  NAND2_X1 u2_u8_u2_U62 (.A2( u2_u8_u2_n107 ) , .A1( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n123 ) );
  NAND2_X1 u2_u8_u2_U63 (.A1( u2_u8_u2_n104 ) , .A2( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n122 ) );
  INV_X1 u2_u8_u2_U64 (.A( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n172 ) );
  NAND2_X1 u2_u8_u2_U65 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n102 ) , .ZN( u2_u8_u2_n116 ) );
  NAND2_X1 u2_u8_u2_U66 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n120 ) );
  NAND2_X1 u2_u8_u2_U67 (.A2( u2_u8_u2_n105 ) , .A1( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n117 ) );
  INV_X1 u2_u8_u2_U68 (.ZN( u2_u8_u2_n187 ) , .A( u2_u8_u2_n99 ) );
  OAI21_X1 u2_u8_u2_U69 (.B1( u2_u8_u2_n137 ) , .B2( u2_u8_u2_n143 ) , .A( u2_u8_u2_n98 ) , .ZN( u2_u8_u2_n99 ) );
  AOI21_X1 u2_u8_u2_U7 (.ZN( u2_u8_u2_n124 ) , .B1( u2_u8_u2_n131 ) , .B2( u2_u8_u2_n143 ) , .A( u2_u8_u2_n172 ) );
  NOR2_X1 u2_u8_u2_U70 (.A2( u2_u8_X_16 ) , .ZN( u2_u8_u2_n140 ) , .A1( u2_u8_u2_n166 ) );
  NOR2_X1 u2_u8_u2_U71 (.A2( u2_u8_X_13 ) , .A1( u2_u8_X_14 ) , .ZN( u2_u8_u2_n100 ) );
  NOR2_X1 u2_u8_u2_U72 (.A2( u2_u8_X_16 ) , .A1( u2_u8_X_17 ) , .ZN( u2_u8_u2_n138 ) );
  NOR2_X1 u2_u8_u2_U73 (.A2( u2_u8_X_15 ) , .A1( u2_u8_X_18 ) , .ZN( u2_u8_u2_n104 ) );
  NOR2_X1 u2_u8_u2_U74 (.A2( u2_u8_X_14 ) , .ZN( u2_u8_u2_n103 ) , .A1( u2_u8_u2_n174 ) );
  NOR2_X1 u2_u8_u2_U75 (.A2( u2_u8_X_15 ) , .ZN( u2_u8_u2_n102 ) , .A1( u2_u8_u2_n165 ) );
  NOR2_X1 u2_u8_u2_U76 (.A2( u2_u8_X_17 ) , .ZN( u2_u8_u2_n114 ) , .A1( u2_u8_u2_n169 ) );
  AND2_X1 u2_u8_u2_U77 (.A1( u2_u8_X_15 ) , .ZN( u2_u8_u2_n105 ) , .A2( u2_u8_u2_n165 ) );
  AND2_X1 u2_u8_u2_U78 (.A2( u2_u8_X_15 ) , .A1( u2_u8_X_18 ) , .ZN( u2_u8_u2_n107 ) );
  AND2_X1 u2_u8_u2_U79 (.A1( u2_u8_X_14 ) , .ZN( u2_u8_u2_n106 ) , .A2( u2_u8_u2_n174 ) );
  AOI21_X1 u2_u8_u2_U8 (.B2( u2_u8_u2_n120 ) , .B1( u2_u8_u2_n121 ) , .ZN( u2_u8_u2_n126 ) , .A( u2_u8_u2_n167 ) );
  AND2_X1 u2_u8_u2_U80 (.A1( u2_u8_X_13 ) , .A2( u2_u8_X_14 ) , .ZN( u2_u8_u2_n108 ) );
  INV_X1 u2_u8_u2_U81 (.A( u2_u8_X_16 ) , .ZN( u2_u8_u2_n169 ) );
  INV_X1 u2_u8_u2_U82 (.A( u2_u8_X_17 ) , .ZN( u2_u8_u2_n166 ) );
  INV_X1 u2_u8_u2_U83 (.A( u2_u8_X_13 ) , .ZN( u2_u8_u2_n174 ) );
  INV_X1 u2_u8_u2_U84 (.A( u2_u8_X_18 ) , .ZN( u2_u8_u2_n165 ) );
  NAND4_X1 u2_u8_u2_U85 (.ZN( u2_out8_30 ) , .A4( u2_u8_u2_n147 ) , .A3( u2_u8_u2_n148 ) , .A2( u2_u8_u2_n149 ) , .A1( u2_u8_u2_n187 ) );
  NOR3_X1 u2_u8_u2_U86 (.A3( u2_u8_u2_n144 ) , .A2( u2_u8_u2_n145 ) , .A1( u2_u8_u2_n146 ) , .ZN( u2_u8_u2_n147 ) );
  AOI21_X1 u2_u8_u2_U87 (.B2( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n148 ) , .A( u2_u8_u2_n162 ) , .B1( u2_u8_u2_n182 ) );
  NAND4_X1 u2_u8_u2_U88 (.ZN( u2_out8_24 ) , .A4( u2_u8_u2_n111 ) , .A3( u2_u8_u2_n112 ) , .A1( u2_u8_u2_n130 ) , .A2( u2_u8_u2_n187 ) );
  AOI221_X1 u2_u8_u2_U89 (.A( u2_u8_u2_n109 ) , .B1( u2_u8_u2_n110 ) , .ZN( u2_u8_u2_n111 ) , .C1( u2_u8_u2_n134 ) , .C2( u2_u8_u2_n170 ) , .B2( u2_u8_u2_n173 ) );
  OAI22_X1 u2_u8_u2_U9 (.ZN( u2_u8_u2_n109 ) , .A2( u2_u8_u2_n113 ) , .B2( u2_u8_u2_n133 ) , .B1( u2_u8_u2_n167 ) , .A1( u2_u8_u2_n168 ) );
  AOI21_X1 u2_u8_u2_U90 (.ZN( u2_u8_u2_n112 ) , .B2( u2_u8_u2_n156 ) , .A( u2_u8_u2_n164 ) , .B1( u2_u8_u2_n181 ) );
  NAND4_X1 u2_u8_u2_U91 (.ZN( u2_out8_16 ) , .A4( u2_u8_u2_n128 ) , .A3( u2_u8_u2_n129 ) , .A1( u2_u8_u2_n130 ) , .A2( u2_u8_u2_n186 ) );
  AOI22_X1 u2_u8_u2_U92 (.A2( u2_u8_u2_n118 ) , .ZN( u2_u8_u2_n129 ) , .A1( u2_u8_u2_n140 ) , .B1( u2_u8_u2_n157 ) , .B2( u2_u8_u2_n170 ) );
  INV_X1 u2_u8_u2_U93 (.A( u2_u8_u2_n163 ) , .ZN( u2_u8_u2_n186 ) );
  OR4_X1 u2_u8_u2_U94 (.ZN( u2_out8_6 ) , .A4( u2_u8_u2_n161 ) , .A3( u2_u8_u2_n162 ) , .A2( u2_u8_u2_n163 ) , .A1( u2_u8_u2_n164 ) );
  OR3_X1 u2_u8_u2_U95 (.A2( u2_u8_u2_n159 ) , .A1( u2_u8_u2_n160 ) , .ZN( u2_u8_u2_n161 ) , .A3( u2_u8_u2_n183 ) );
  AOI21_X1 u2_u8_u2_U96 (.B2( u2_u8_u2_n154 ) , .B1( u2_u8_u2_n155 ) , .ZN( u2_u8_u2_n159 ) , .A( u2_u8_u2_n167 ) );
  NAND3_X1 u2_u8_u2_U97 (.A2( u2_u8_u2_n117 ) , .A1( u2_u8_u2_n122 ) , .A3( u2_u8_u2_n123 ) , .ZN( u2_u8_u2_n134 ) );
  NAND3_X1 u2_u8_u2_U98 (.ZN( u2_u8_u2_n110 ) , .A2( u2_u8_u2_n131 ) , .A3( u2_u8_u2_n139 ) , .A1( u2_u8_u2_n154 ) );
  NAND3_X1 u2_u8_u2_U99 (.A2( u2_u8_u2_n100 ) , .ZN( u2_u8_u2_n101 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n114 ) );
  OAI21_X1 u2_uk_U1033 (.ZN( u2_K15_32 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1825 ) , .A( u2_uk_n941 ) );
  NAND2_X1 u2_uk_U1040 (.A1( u2_uk_K_r2_50 ) , .A2( u2_uk_n102 ) , .ZN( u2_uk_n1034 ) );
  INV_X1 u2_uk_U1060 (.A( u2_key_r_1 ) , .ZN( u2_uk_n1143 ) );
  OAI22_X1 u2_uk_U107 (.ZN( u2_K14_41 ) , .A1( u2_uk_n147 ) , .A2( u2_uk_n1776 ) , .B2( u2_uk_n1781 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1098 (.ZN( u2_K8_12 ) , .A( u2_uk_n1098 ) );
  AOI22_X1 u2_uk_U1099 (.B2( u2_uk_K_r6_3 ) , .A2( u2_uk_K_r6_53 ) , .ZN( u2_uk_n1098 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n220 ) );
  INV_X1 u2_uk_U1122 (.ZN( u2_K4_20 ) , .A( u2_uk_n1024 ) );
  INV_X1 u2_uk_U113 (.ZN( u2_K11_47 ) , .A( u2_uk_n386 ) );
  AOI22_X1 u2_uk_U114 (.B2( u2_uk_K_r9_15 ) , .A2( u2_uk_K_r9_23 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n223 ) , .ZN( u2_uk_n386 ) );
  INV_X1 u2_uk_U1143 (.ZN( u2_K15_43 ) , .A( u2_uk_n944 ) );
  INV_X1 u2_uk_U1153 (.ZN( u2_K9_2 ) , .A( u2_uk_n1130 ) );
  INV_X1 u2_uk_U12 (.A( u2_uk_n145 ) , .ZN( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U125 (.ZN( u2_K4_15 ) , .B2( u2_uk_n1328 ) , .A2( u2_uk_n1356 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U14 (.A( u2_uk_n145 ) , .ZN( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U146 (.ZN( u2_K14_15 ) , .A2( u2_uk_n1773 ) , .B2( u2_uk_n1811 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U16 (.A( u2_uk_n146 ) , .ZN( u2_uk_n99 ) );
  INV_X1 u2_uk_U17 (.ZN( u2_uk_n109 ) , .A( u2_uk_n146 ) );
  OAI21_X1 u2_uk_U181 (.ZN( u2_K9_14 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1121 ) , .B2( u2_uk_n1574 ) );
  INV_X1 u2_uk_U19 (.ZN( u2_uk_n100 ) , .A( u2_uk_n146 ) );
  OAI22_X1 u2_uk_U196 (.ZN( u2_K4_24 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1322 ) , .A2( u2_uk_n1363 ) , .B1( u2_uk_n142 ) );
  INV_X1 u2_uk_U20 (.ZN( u2_uk_n102 ) , .A( u2_uk_n146 ) );
  INV_X1 u2_uk_U206 (.ZN( u2_K15_30 ) , .A( u2_uk_n940 ) );
  AOI22_X1 u2_uk_U207 (.B2( u2_uk_K_r13_0 ) , .A2( u2_uk_K_r13_38 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n940 ) );
  INV_X1 u2_uk_U21 (.ZN( u2_uk_n128 ) , .A( u2_uk_n223 ) );
  BUF_X1 u2_uk_U22 (.Z( u2_uk_n141 ) , .A( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U235 (.ZN( u2_K14_31 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1797 ) , .A2( u2_uk_n1803 ) , .A1( u2_uk_n94 ) );
  BUF_X1 u2_uk_U24 (.Z( u2_uk_n145 ) , .A( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U249 (.ZN( u2_K15_44 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1836 ) , .A2( u2_uk_n1854 ) , .A1( u2_uk_n230 ) );
  BUF_X1 u2_uk_U25 (.Z( u2_uk_n142 ) , .A( u2_uk_n222 ) );
  OAI21_X1 u2_uk_U250 (.ZN( u2_K15_48 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1824 ) , .A( u2_uk_n945 ) );
  OAI22_X1 u2_uk_U259 (.ZN( u2_K11_44 ) , .A1( u2_uk_n142 ) , .B2( u2_uk_n1653 ) , .A2( u2_uk_n1673 ) , .B1( u2_uk_n63 ) );
  BUF_X1 u2_uk_U28 (.Z( u2_uk_n146 ) , .A( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U294 (.ZN( u2_K3_8 ) , .A2( u2_uk_n1280 ) , .B2( u2_uk_n1296 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U3 (.ZN( u2_uk_n10 ) , .A( u2_uk_n141 ) );
  BUF_X1 u2_uk_U30 (.Z( u2_uk_n161 ) , .A( u2_uk_n213 ) );
  INV_X1 u2_uk_U305 (.ZN( u2_K15_26 ) , .A( u2_uk_n939 ) );
  BUF_X1 u2_uk_U32 (.Z( u2_uk_n162 ) , .A( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U322 (.ZN( u2_K15_46 ) , .B1( u2_uk_n17 ) , .A2( u2_uk_n1818 ) , .B2( u2_uk_n1845 ) , .A1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U330 (.A1( u2_key_r_49 ) , .A2( u2_uk_n94 ) , .ZN( u2_uk_n988 ) );
  OAI22_X1 u2_uk_U332 (.ZN( u2_K14_4 ) , .B2( u2_uk_n1786 ) , .A2( u2_uk_n1794 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U334 (.ZN( u2_K11_46 ) , .A( u2_uk_n385 ) );
  OAI21_X1 u2_uk_U352 (.ZN( u2_K14_40 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1793 ) , .A( u2_uk_n702 ) );
  OAI22_X1 u2_uk_U355 (.ZN( u2_K15_40 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n17 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1849 ) );
  OAI21_X1 u2_uk_U362 (.ZN( u2_K15_33 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1840 ) , .A( u2_uk_n942 ) );
  OAI22_X1 u2_uk_U383 (.ZN( u2_K14_1 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1778 ) , .A2( u2_uk_n1783 ) );
  OAI22_X1 u2_uk_U398 (.ZN( u2_K9_16 ) , .B2( u2_uk_n1548 ) , .A2( u2_uk_n1555 ) , .B1( u2_uk_n220 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U403 (.ZN( u2_K4_16 ) , .B2( u2_uk_n1329 ) , .A2( u2_uk_n1333 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U409 (.ZN( u2_K14_9 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1788 ) , .A( u2_uk_n933 ) );
  BUF_X1 u2_uk_U41 (.Z( u2_uk_n203 ) , .A( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U414 (.ZN( u2_K8_9 ) , .A2( u2_uk_n1502 ) , .B2( u2_uk_n1508 ) , .B1( u2_uk_n161 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U422 (.ZN( u2_K9_9 ) , .A( u2_uk_n1141 ) );
  OAI21_X1 u2_uk_U428 (.ZN( u2_K3_9 ) , .A( u2_uk_n1019 ) , .B2( u2_uk_n1295 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U429 (.A1( u2_uk_K_r1_18 ) , .ZN( u2_uk_n1019 ) , .A2( u2_uk_n217 ) );
  BUF_X1 u2_uk_U43 (.A( u2_uk_n141 ) , .Z( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U453 (.ZN( u2_K14_33 ) , .A1( u2_uk_n155 ) , .B2( u2_uk_n1785 ) , .A2( u2_uk_n1803 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U460 (.ZN( u2_K15_37 ) , .A2( u2_uk_n1819 ) , .B2( u2_uk_n1846 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U461 (.ZN( u2_K14_37 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1785 ) , .A2( u2_uk_n1791 ) , .A1( u2_uk_n94 ) );
  BUF_X1 u2_uk_U47 (.Z( u2_uk_n223 ) , .A( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U496 (.ZN( u2_K14_2 ) , .B2( u2_uk_n1794 ) , .A2( u2_uk_n1801 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U5 (.ZN( u2_uk_n117 ) , .A( u2_uk_n161 ) );
  OAI21_X1 u2_uk_U505 (.ZN( u2_K9_12 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1119 ) , .B2( u2_uk_n1543 ) );
  OAI21_X1 u2_uk_U512 (.ZN( u2_K9_17 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1122 ) , .B2( u2_uk_n1568 ) );
  NAND2_X1 u2_uk_U513 (.A1( u2_uk_K_r7_26 ) , .ZN( u2_uk_n1122 ) , .A2( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U517 (.ZN( u2_K4_17 ) , .A( u2_uk_n1021 ) , .B2( u2_uk_n1339 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U518 (.A1( u2_uk_K_r2_27 ) , .ZN( u2_uk_n1021 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U530 (.ZN( u2_K3_12 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1306 ) , .A2( u2_uk_n1311 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U548 (.ZN( u2_K15_36 ) , .B2( u2_uk_n1826 ) , .A2( u2_uk_n1840 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U549 (.ZN( u2_K14_36 ) , .A1( u2_uk_n141 ) , .B2( u2_uk_n1770 ) , .A2( u2_uk_n1808 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U564 (.ZN( u2_K15_38 ) , .A( u2_uk_n943 ) );
  INV_X1 u2_uk_U579 (.ZN( u2_K9_10 ) , .A( u2_uk_n1117 ) );
  AOI22_X1 u2_uk_U580 (.B2( u2_uk_K_r7_25 ) , .A2( u2_uk_K_r7_32 ) , .B1( u2_uk_n110 ) , .ZN( u2_uk_n1117 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U581 (.ZN( u2_K8_10 ) , .B2( u2_uk_n1519 ) , .A2( u2_uk_n1521 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U6 (.A( u2_uk_n146 ) , .ZN( u2_uk_n17 ) );
  INV_X1 u2_uk_U61 (.ZN( u2_K14_34 ) , .A( u2_uk_n692 ) );
  INV_X1 u2_uk_U612 (.ZN( u2_K14_35 ) , .A( u2_uk_n694 ) );
  AOI22_X1 u2_uk_U613 (.B2( u2_uk_K_r12_1 ) , .A2( u2_uk_K_r12_7 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n694 ) );
  AOI22_X1 u2_uk_U62 (.B2( u2_uk_K_r12_30 ) , .A2( u2_uk_K_r12_36 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n692 ) );
  OAI21_X1 u2_uk_U633 (.ZN( u2_K8_11 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1097 ) , .B2( u2_uk_n1535 ) );
  INV_X1 u2_uk_U635 (.ZN( u2_K9_11 ) , .A( u2_uk_n1118 ) );
  AOI22_X1 u2_uk_U636 (.B2( u2_uk_K_r7_48 ) , .A2( u2_uk_K_r7_55 ) , .B1( u2_uk_n100 ) , .ZN( u2_uk_n1118 ) , .A1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U639 (.ZN( u2_K3_11 ) , .A2( u2_uk_n1280 ) , .B2( u2_uk_n1285 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U671 (.ZN( u2_K11_43 ) , .A1( u2_uk_n161 ) , .B2( u2_uk_n1632 ) , .A2( u2_uk_n1674 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U707 (.ZN( u2_K15_25 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1846 ) , .A( u2_uk_n938 ) );
  NAND2_X1 u2_uk_U708 (.A1( u2_uk_K_r13_22 ) , .A2( u2_uk_n214 ) , .ZN( u2_uk_n938 ) );
  OAI22_X1 u2_uk_U723 (.ZN( u2_K14_32 ) , .A1( u2_uk_n155 ) , .B2( u2_uk_n1769 ) , .A2( u2_uk_n1807 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U727 (.ZN( u2_K15_42 ) , .B1( u2_uk_n161 ) , .B2( u2_uk_n1849 ) , .A2( u2_uk_n1855 ) , .A1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U754 (.ZN( u2_K9_13 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1120 ) , .B2( u2_uk_n1549 ) );
  INV_X1 u2_uk_U76 (.ZN( u2_K4_23 ) , .A( u2_uk_n1026 ) );
  OAI22_X1 u2_uk_U767 (.ZN( u2_K15_27 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1835 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  AOI22_X1 u2_uk_U77 (.B2( u2_uk_K_r2_18 ) , .A2( u2_uk_K_r2_55 ) , .ZN( u2_uk_n1026 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U775 (.ZN( u2_K4_13 ) , .A1( u2_uk_n102 ) , .A2( u2_uk_n1324 ) , .B2( u2_uk_n1328 ) , .B1( u2_uk_n230 ) );
  INV_X1 u2_uk_U797 (.ZN( u2_K9_1 ) , .A( u2_uk_n1125 ) );
  OAI21_X1 u2_uk_U799 (.ZN( u2_K4_18 ) , .B1( u2_uk_n10 ) , .A( u2_uk_n1022 ) , .B2( u2_uk_n1348 ) );
  INV_X1 u2_uk_U8 (.A( u2_uk_n145 ) , .ZN( u2_uk_n63 ) );
  NAND2_X1 u2_uk_U804 (.A1( u2_uk_K_r11_33 ) , .ZN( u2_uk_n605 ) , .A2( u2_uk_n99 ) );
  INV_X1 u2_uk_U820 (.ZN( u2_K9_18 ) , .A( u2_uk_n1123 ) );
  AOI22_X1 u2_uk_U821 (.B2( u2_uk_K_r7_39 ) , .A2( u2_uk_K_r7_46 ) , .B1( u2_uk_n110 ) , .ZN( u2_uk_n1123 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U863 (.ZN( u2_K3_10 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1286 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1291 ) );
  OAI22_X1 u2_uk_U864 (.ZN( u2_K15_45 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1837 ) , .A2( u2_uk_n1855 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U873 (.ZN( u2_K9_7 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1544 ) , .B2( u2_uk_n1548 ) );
  OAI22_X1 u2_uk_U876 (.ZN( u2_K14_7 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1786 ) , .A2( u2_uk_n1805 ) );
  OAI22_X1 u2_uk_U88 (.ZN( u2_K15_41 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1835 ) , .A2( u2_uk_n1853 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U913 (.ZN( u2_K9_6 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1555 ) , .A2( u2_uk_n1563 ) , .B1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U914 (.ZN( u2_K9_8 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1573 ) , .A2( u2_uk_n1580 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U923 (.ZN( u2_K15_47 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1824 ) , .A2( u2_uk_n1856 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U930 (.ZN( u2_K9_4 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1549 ) , .A2( u2_uk_n1556 ) , .B1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U937 (.ZN( u2_K4_19 ) , .B2( u2_uk_n1335 ) , .A2( u2_uk_n1347 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U94 (.ZN( u2_K14_5 ) , .B2( u2_uk_n1796 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n932 ) );
  OAI22_X1 u2_uk_U943 (.ZN( u2_K14_38 ) , .B1( u2_uk_n145 ) , .A2( u2_uk_n1777 ) , .B2( u2_uk_n1793 ) , .A1( u2_uk_n93 ) );
  NAND2_X1 u2_uk_U95 (.A1( u2_uk_K_r12_10 ) , .A2( u2_uk_n223 ) , .ZN( u2_uk_n932 ) );
  OAI22_X1 u2_uk_U958 (.ZN( u2_K8_7 ) , .A2( u2_uk_n1500 ) , .B2( u2_uk_n1506 ) , .B1( u2_uk_n164 ) , .A1( u2_uk_n92 ) );
endmodule

