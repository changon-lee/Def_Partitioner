module aes_aes_die_5 ( n101, n103, n105, n1109, n1114, n115, n117, n119, n121, 
       n13, n143, n15, n195, n197, n199, n201, n203, n207, 
       n209, n21, n213, n215, n217, n219, n225, n23, n231, 
       n247, n249, n25, n253, n3, n31, n33, n35, n37, 
       n47, n49, n5, n51, n53, n55, n57, n59, n61, 
       n63, n65, n665, n67, n69, n7, n73, n79, n81, 
       n85, n9, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, 
       sa00_sr_7, sa01_sr_6, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
       sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, 
       sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa10_sr_0, 
       sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa12_sr_0, sa12_sr_1, 
       sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, 
       sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
       sa22_sr_4, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, 
       sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, 
       sa30_sr_7, sa31_sr_6, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, 
       sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, 
       w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_15, w0_16, w0_18, 
       w0_19, w0_2, w0_20, w0_25, w0_26, w0_27, w0_28, w0_3, w0_30, 
       w0_4, w0_5, w0_7, w0_8, w1_7, w2_0, w2_1, w2_10, w2_11, 
       w2_13, w2_16, w2_18, w2_19, w2_2, w2_20, w2_25, w2_26, w2_27, 
       w2_28, w2_4, w2_7, w2_8, w2_9, w3_0, w3_1, w3_10, w3_11, 
       w3_12, w3_13, w3_15, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, 
       w3_21, w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, 
       w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9, N100, N102, N105, N114, N116, N132, N133, N134, N147, 
        N148, N149, N150, N169, N227, N228, N229, N230, N231, 
        N233, N242, N244, N245, N246, N247, N258, N261, N277, 
        N278, N280, N35, N36, N37, N38, N40, N41, N430, 
        N434, N435, N436, N437, N438, N439, N440, N441, N463, 
        N52, N53, N54, N57, N66, N67, N68, N73, N82, 
        N83, N84, N85, N86, N87, N88, N89, N98, N99, 
        n1145, n1183, n1212, n1213, n1214, n1215, n1216, n1217, n1219, 
        n1220, n1221, n342, n348, n354, n362, n394, n396, n414, 
        n419, n433, n462, n469, n481, n482, n500, n506, n515, 
        n524, n534, n547, n562, n590, n636, n817, n823, n830, 
        n861, n870, n900, n905, n911, n917, n923, n927, n937, 
        n957, u0_n49, u0_n53, u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, u0_subword_6 );
  input n101, n103, n105, n1109, n1114, n115, n117, n119, n121, 
        n13, n143, n15, n195, n197, n199, n201, n203, n207, 
        n209, n21, n213, n215, n217, n219, n225, n23, n231, 
        n247, n249, n25, n253, n3, n31, n33, n35, n37, 
        n47, n49, n5, n51, n53, n55, n57, n59, n61, 
        n63, n65, n665, n67, n69, n7, n73, n79, n81, 
        n85, n9, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, 
        sa00_sr_7, sa01_sr_6, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, 
        sa02_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, 
        sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa10_sr_0, 
        sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa12_sr_0, sa12_sr_1, 
        sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_7, sa20_sr_0, sa20_sr_1, sa20_sr_2, sa20_sr_3, 
        sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, 
        sa22_sr_4, sa22_sr_6, sa22_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, 
        sa23_sr_6, sa23_sr_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, 
        sa30_sr_7, sa31_sr_6, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, 
        sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, 
        w0_0, w0_1, w0_10, w0_11, w0_12, w0_13, w0_15, w0_16, w0_18, 
        w0_19, w0_2, w0_20, w0_25, w0_26, w0_27, w0_28, w0_3, w0_30, 
        w0_4, w0_5, w0_7, w0_8, w1_7, w2_0, w2_1, w2_10, w2_11, 
        w2_13, w2_16, w2_18, w2_19, w2_2, w2_20, w2_25, w2_26, w2_27, 
        w2_28, w2_4, w2_7, w2_8, w2_9, w3_0, w3_1, w3_10, w3_11, 
        w3_12, w3_13, w3_15, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, 
        w3_21, w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, 
        w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9;
  output N100, N102, N105, N114, N116, N132, N133, N134, N147, 
        N148, N149, N150, N169, N227, N228, N229, N230, N231, 
        N233, N242, N244, N245, N246, N247, N258, N261, N277, 
        N278, N280, N35, N36, N37, N38, N40, N41, N430, 
        N434, N435, N436, N437, N438, N439, N440, N441, N463, 
        N52, N53, N54, N57, N66, N67, N68, N73, N82, 
        N83, N84, N85, N86, N87, N88, N89, N98, N99, 
        n1145, n1183, n1212, n1213, n1214, n1215, n1216, n1217, n1219, 
        n1220, n1221, n342, n348, n354, n362, n394, n396, n414, 
        n419, n433, n462, n469, n481, n482, n500, n506, n515, 
        n524, n534, n547, n562, n590, n636, n817, n823, n830, 
        n861, n870, n900, n905, n911, n917, n923, n927, n937, 
        n957, u0_n49, u0_n53, u0_n55, u0_n57, u0_n59, u0_n61, u0_n63, u0_subword_6;
  wire n1115, n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, 
       n1126, n1127, n1128, n1130, n1133, n1134, n1135, n1137, n1138, 
       n1139, n1140, n1141, n1142, n1144, n1148, n1149, n1150, n1153, 
       n1155, n1165, n1166, n1168, n1172, n1173, n1175, n1178, n1179, 
       n1180, n1181, n1182, n1188, n1190, n1193, n1194, n1195, n1196, 
       n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1208, n1209, 
       n1210, n1211, n271, n272, n275, n276, n277, n278, n279, 
       n280, n281, n283, n284, n285, n286, n288, n289, n290, 
       n291, n292, n294, n295, n296, n297, n298, n300, n301, 
       n302, n303, n304, n305, n306, n307, n308, n309, n310, 
       n311, n312, n314, n315, n316, n317, n318, n319, n321, 
       n322, n323, n324, n325, n327, n328, n329, n330, n331, 
       n332, n334, n335, n336, n337, n338, n339, n343, n345, 
       n349, n350, n351, n352, n355, n356, n357, n358, n359, 
       n360, n363, n365, n366, n367, n368, n369, n370, n372, 
       n373, n374, n375, n376, n378, n379, n380, n381, n382, 
       n384, n385, n386, n387, n388, n390, n398, n399, n400, 
       n401, n402, n403, n404, n405, n407, n408, n409, n410, 
       n412, n416, n417, n421, n422, n423, n424, n425, n426, 
       n427, n428, n429, n431, n434, n436, n437, n438, n439, 
       n440, n441, n442, n443, n444, n445, n446, n448, n449, 
       n450, n451, n452, n453, n454, n455, n456, n457, n459, 
       n460, n464, n472, n473, n475, n476, n477, n483, n484, 
       n485, n486, n487, n488, n489, n490, n491, n492, n493, 
       n495, n496, n497, n498, n502, n503, n504, n508, n509, 
       n510, n511, n516, n535, n536, n537, n538, n539, n540, 
       n541, n542, n543, n544, n548, n550, n556, n557, n558, 
       n560, n564, n569, n570, n571, n572, n573, n574, n575, 
       n576, n577, n578, n579, n581, n582, n583, n584, n586, 
       n592, n593, n595, n596, n597, n598, n599, n600, n606, 
       n607, n608, n609, n610, n611, n612, n613, n614, n615, 
       n616, n617, n618, n619, n620, n622, n623, n624, n625, 
       n626, n628, n629, n630, n632, n633, n634, n638, n770, 
       n771, n772, n773, n774, n824, n825, n832, n833, n834, 
       n835, n836, n837, n838, n839, n840, n841, n843, n844, 
       n845, n846, n847, n848, n850, n851, n852, n853, n854, 
       n856, n857, n862, n879, n880, n881, n882, n883, n884, 
       n885, n886, n887, n888, n889, n890, n892, n893, n894, 
       n896, n903, n907, n918, n919, n924, n929, n930, n931, 
       n932, n933, n935, n939, n940, n941, n942, n944, n945, 
       n946, n947, n948, n949, n960, n961, n962, n964, n965, 
       n971, n972, n973, n974, n975, n976, sa13_sr_0, sa13_sr_1, sa13_sr_2, 
       sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, u0_subword_0, u0_subword_1, u0_subword_2, u0_subword_3, 
       u0_subword_4, u0_subword_5, u0_subword_7, u0_u3_n41, u0_u3_n438, u0_u3_n439, u0_u3_n440, u0_u3_n441, u0_u3_n442, 
       u0_u3_n443, u0_u3_n444, u0_u3_n445, u0_u3_n446, u0_u3_n447, u0_u3_n448, u0_u3_n449, u0_u3_n450, u0_u3_n451, 
       u0_u3_n452, u0_u3_n453, u0_u3_n454, u0_u3_n455, u0_u3_n456, u0_u3_n457, u0_u3_n458, u0_u3_n459, u0_u3_n460, 
       u0_u3_n461, u0_u3_n462, u0_u3_n463, u0_u3_n464, u0_u3_n465, u0_u3_n466, u0_u3_n467, u0_u3_n468, u0_u3_n469, 
       u0_u3_n470, u0_u3_n471, u0_u3_n472, u0_u3_n473, u0_u3_n474, u0_u3_n475, u0_u3_n476, u0_u3_n477, u0_u3_n478, 
       u0_u3_n479, u0_u3_n480, u0_u3_n481, u0_u3_n482, u0_u3_n483, u0_u3_n484, u0_u3_n485, u0_u3_n486, u0_u3_n487, 
       u0_u3_n488, u0_u3_n489, u0_u3_n490, u0_u3_n491, u0_u3_n492, u0_u3_n493, u0_u3_n494, u0_u3_n495, u0_u3_n496, 
       u0_u3_n497, u0_u3_n498, u0_u3_n499, u0_u3_n500, u0_u3_n501, u0_u3_n502, u0_u3_n503, u0_u3_n504, u0_u3_n505, 
       u0_u3_n506, u0_u3_n507, u0_u3_n508, u0_u3_n509, u0_u3_n510, u0_u3_n511, u0_u3_n512, u0_u3_n513, u0_u3_n514, 
       u0_u3_n515, u0_u3_n516, u0_u3_n517, u0_u3_n518, u0_u3_n519, u0_u3_n520, u0_u3_n521, u0_u3_n522, u0_u3_n523, 
       u0_u3_n524, u0_u3_n525, u0_u3_n526, u0_u3_n527, u0_u3_n528, u0_u3_n529, u0_u3_n530, u0_u3_n531, u0_u3_n532, 
       u0_u3_n533, u0_u3_n534, u0_u3_n535, u0_u3_n536, u0_u3_n537, u0_u3_n538, u0_u3_n539, u0_u3_n540, u0_u3_n541, 
       u0_u3_n542, u0_u3_n543, u0_u3_n544, u0_u3_n545, u0_u3_n546, u0_u3_n547, u0_u3_n548, u0_u3_n549, u0_u3_n550, 
       u0_u3_n551, u0_u3_n552, u0_u3_n553, u0_u3_n554, u0_u3_n555, u0_u3_n556, u0_u3_n557, u0_u3_n558, u0_u3_n559, 
       u0_u3_n560, u0_u3_n561, u0_u3_n562, u0_u3_n563, u0_u3_n564, u0_u3_n565, u0_u3_n566, u0_u3_n567, u0_u3_n568, 
       u0_u3_n569, u0_u3_n570, u0_u3_n571, u0_u3_n572, u0_u3_n573, u0_u3_n574, u0_u3_n575, u0_u3_n576, u0_u3_n577, 
       u0_u3_n578, u0_u3_n579, u0_u3_n580, u0_u3_n581, u0_u3_n582, u0_u3_n583, u0_u3_n584, u0_u3_n585, u0_u3_n586, 
       u0_u3_n587, u0_u3_n588, u0_u3_n589, u0_u3_n590, u0_u3_n591, u0_u3_n592, u0_u3_n593, u0_u3_n594, u0_u3_n595, 
       u0_u3_n596, u0_u3_n597, u0_u3_n598, u0_u3_n599, u0_u3_n600, u0_u3_n601, u0_u3_n602, u0_u3_n603, u0_u3_n604, 
       u0_u3_n605, u0_u3_n606, u0_u3_n607, u0_u3_n608, u0_u3_n609, u0_u3_n610, u0_u3_n611, u0_u3_n612, u0_u3_n613, 
       u0_u3_n614, u0_u3_n615, u0_u3_n616, u0_u3_n617, u0_u3_n618, u0_u3_n619, u0_u3_n620, u0_u3_n621, u0_u3_n622, 
       u0_u3_n623, u0_u3_n624, u0_u3_n625, u0_u3_n626, u0_u3_n627, u0_u3_n628, u0_u3_n629, u0_u3_n630, u0_u3_n631, 
       u0_u3_n632, u0_u3_n633, u0_u3_n634, u0_u3_n635, u0_u3_n636, u0_u3_n637, u0_u3_n638, u0_u3_n639, u0_u3_n640, 
       u0_u3_n641, u0_u3_n642, u0_u3_n643, u0_u3_n644, u0_u3_n645, u0_u3_n646, u0_u3_n647, u0_u3_n648, u0_u3_n649, 
       u0_u3_n650, u0_u3_n651, u0_u3_n652, u0_u3_n653, u0_u3_n654, u0_u3_n655, u0_u3_n656, u0_u3_n657, u0_u3_n658, 
       u0_u3_n659, u0_u3_n660, u0_u3_n661, u0_u3_n662, u0_u3_n663, u0_u3_n664, u0_u3_n665, u0_u3_n666, u0_u3_n667, 
       u0_u3_n668, u0_u3_n669, u0_u3_n670, u0_u3_n671, u0_u3_n672, u0_u3_n673, u0_u3_n674, u0_u3_n675, u0_u3_n676, 
       u0_u3_n677, u0_u3_n678, u0_u3_n679, u0_u3_n680, u0_u3_n681, u0_u3_n682, u0_u3_n683, u0_u3_n684, u0_u3_n685, 
       u0_u3_n686, u0_u3_n687, u0_u3_n688, u0_u3_n689, u0_u3_n690, u0_u3_n691, u0_u3_n692, u0_u3_n693, u0_u3_n694, 
       u0_u3_n695, u0_u3_n696, u0_u3_n697, u0_u3_n698, u0_u3_n699, u0_u3_n700, u0_u3_n701, u0_u3_n702, u0_u3_n703, 
       u0_u3_n704, u0_u3_n705, u0_u3_n706, u0_u3_n707, u0_u3_n708, u0_u3_n709, u0_u3_n710, u0_u3_n711, u0_u3_n712, 
       u0_u3_n713, u0_u3_n714, u0_u3_n715, u0_u3_n716, u0_u3_n717, u0_u3_n718, u0_u3_n719, u0_u3_n720, u0_u3_n721, 
       u0_u3_n722, u0_u3_n723, u0_u3_n724, u0_u3_n725, u0_u3_n726, u0_u3_n727, u0_u3_n728, u0_u3_n729, u0_u3_n730, 
       u0_u3_n731, u0_u3_n732, u0_u3_n733, u0_u3_n734, u0_u3_n735, u0_u3_n736, u0_u3_n737, u0_u3_n738, u0_u3_n739, 
       u0_u3_n740, u0_u3_n741, u0_u3_n742, u0_u3_n743, u0_u3_n744, u0_u3_n745, u0_u3_n746, u0_u3_n747, u0_u3_n748, 
       u0_u3_n749, u0_u3_n750, u0_u3_n751, u0_u3_n752, u0_u3_n753, u0_u3_n754, u0_u3_n755, u0_u3_n756, u0_u3_n757, 
       u0_u3_n758, u0_u3_n759, u0_u3_n760, u0_u3_n761, u0_u3_n762, u0_u3_n763, u0_u3_n764, u0_u3_n765, u0_u3_n766, 
       u0_u3_n767, u0_u3_n768, u0_u3_n769, u0_u3_n770, u0_u3_n771, u0_u3_n772, u0_u3_n773, u0_u3_n774, u0_u3_n775, 
       u0_u3_n776, u0_u3_n777, u0_u3_n778, u0_u3_n779, u0_u3_n780, u0_u3_n781, u0_u3_n782, u0_u3_n783, u0_u3_n784, 
       u0_u3_n785, u0_u3_n786, u0_u3_n787, u0_u3_n788, u0_u3_n789, u0_u3_n790, u0_u3_n791, u0_u3_n792, u0_u3_n793, 
       u0_u3_n794, u0_u3_n795, u0_u3_n796, u0_u3_n797, u0_u3_n798, u0_u3_n799, u0_u3_n800, u0_u3_n801, u0_u3_n802, 
       u0_u3_n803, u0_u3_n804, u0_u3_n805, u0_u3_n806, u0_u3_n807, u0_u3_n808, u0_u3_n809, u0_u3_n810, u0_u3_n811, 
       u0_u3_n812, u0_u3_n813, u0_u3_n814, u0_u3_n815, u0_u3_n816, u0_u3_n817, u0_u3_n818, u0_u3_n819, u0_u3_n820, 
       u0_u3_n821, u0_u3_n822, u0_u3_n823, u0_u3_n824, u0_u3_n825, u0_u3_n826, u0_u3_n827, u0_u3_n828, u0_u3_n829, 
       u0_u3_n830, u0_u3_n831, u0_u3_n832, u0_u3_n833, u0_u3_n834, u0_u3_n835, u0_u3_n836, u0_u3_n837, u0_u3_n838, 
       u0_u3_n839, u0_u3_n840, u0_u3_n841, u0_u3_n842, u0_u3_n843, u0_u3_n844, u0_u3_n845, u0_u3_n846, u0_u3_n847, 
       u0_u3_n848, u0_u3_n849, u0_u3_n850, u0_u3_n851, u0_u3_n852, u0_u3_n853, u0_u3_n854, u0_u3_n855, u0_u3_n856, 
       u0_u3_n857, u0_u3_n858, u0_u3_n859, u0_u3_n860, u0_u3_n861, u0_u3_n862, u0_u3_n863, u0_u3_n864, u0_u3_n865, 
       u0_u3_n866, u0_u3_n867, u0_u3_n868, u0_u3_n869, u0_u3_n870, u0_u3_n871, u0_u3_n872, u0_u3_n873, u0_u3_n874, 
       u0_u3_n875, u0_u3_n876, u0_u3_n877, u0_u3_n878, us10_n438, us10_n439, us10_n440, us10_n441, us10_n442, 
       us10_n443, us10_n444, us10_n445, us10_n446, us10_n447, us10_n448, us10_n449, us10_n450, us10_n451, 
       us10_n452, us10_n453, us10_n454, us10_n455, us10_n456, us10_n457, us10_n458, us10_n459, us10_n460, 
       us10_n461, us10_n462, us10_n463, us10_n464, us10_n465, us10_n466, us10_n467, us10_n468, us10_n469, 
       us10_n470, us10_n471, us10_n472, us10_n473, us10_n474, us10_n475, us10_n476, us10_n477, us10_n478, 
       us10_n479, us10_n480, us10_n481, us10_n482, us10_n483, us10_n484, us10_n485, us10_n486, us10_n487, 
       us10_n488, us10_n489, us10_n490, us10_n491, us10_n492, us10_n493, us10_n494, us10_n495, us10_n496, 
       us10_n497, us10_n498, us10_n499, us10_n500, us10_n501, us10_n502, us10_n503, us10_n504, us10_n505, 
       us10_n506, us10_n507, us10_n508, us10_n509, us10_n510, us10_n511, us10_n512, us10_n513, us10_n514, 
       us10_n515, us10_n516, us10_n517, us10_n518, us10_n519, us10_n520, us10_n521, us10_n522, us10_n523, 
       us10_n524, us10_n525, us10_n526, us10_n527, us10_n528, us10_n529, us10_n530, us10_n531, us10_n532, 
       us10_n533, us10_n534, us10_n535, us10_n536, us10_n537, us10_n538, us10_n539, us10_n540, us10_n541, 
       us10_n542, us10_n543, us10_n544, us10_n545, us10_n546, us10_n547, us10_n548, us10_n549, us10_n550, 
       us10_n551, us10_n552, us10_n553, us10_n554, us10_n555, us10_n556, us10_n557, us10_n558, us10_n559, 
       us10_n560, us10_n561, us10_n562, us10_n563, us10_n564, us10_n565, us10_n566, us10_n567, us10_n568, 
       us10_n569, us10_n570, us10_n571, us10_n572, us10_n573, us10_n574, us10_n575, us10_n576, us10_n577, 
       us10_n578, us10_n579, us10_n580, us10_n581, us10_n582, us10_n583, us10_n584, us10_n585, us10_n586, 
       us10_n587, us10_n588, us10_n589, us10_n590, us10_n591, us10_n592, us10_n593, us10_n594, us10_n595, 
       us10_n596, us10_n597, us10_n598, us10_n599, us10_n600, us10_n601, us10_n602, us10_n603, us10_n604, 
       us10_n605, us10_n606, us10_n607, us10_n608, us10_n609, us10_n610, us10_n611, us10_n612, us10_n613, 
       us10_n614, us10_n615, us10_n616, us10_n617, us10_n618, us10_n619, us10_n620, us10_n621, us10_n622, 
       us10_n623, us10_n624, us10_n625, us10_n626, us10_n627, us10_n628, us10_n629, us10_n630, us10_n631, 
       us10_n632, us10_n633, us10_n634, us10_n635, us10_n636, us10_n637, us10_n638, us10_n639, us10_n640, 
       us10_n641, us10_n642, us10_n643, us10_n644, us10_n645, us10_n646, us10_n647, us10_n648, us10_n649, 
       us10_n650, us10_n651, us10_n652, us10_n653, us10_n654, us10_n655, us10_n656, us10_n657, us10_n658, 
       us10_n659, us10_n660, us10_n661, us10_n662, us10_n663, us10_n664, us10_n665, us10_n666, us10_n667, 
       us10_n668, us10_n669, us10_n670, us10_n671, us10_n672, us10_n673, us10_n674, us10_n675, us10_n676, 
       us10_n677, us10_n678, us10_n679, us10_n680, us10_n681, us10_n682, us10_n683, us10_n684, us10_n685, 
       us10_n686, us10_n687, us10_n688, us10_n689, us10_n690, us10_n691, us10_n692, us10_n693, us10_n694, 
       us10_n695, us10_n696, us10_n697, us10_n698, us10_n699, us10_n700, us10_n701, us10_n702, us10_n703, 
       us10_n704, us10_n705, us10_n706, us10_n707, us10_n708, us10_n709, us10_n710, us10_n711, us10_n712, 
       us10_n713, us10_n714, us10_n715, us10_n716, us10_n717, us10_n718, us10_n719, us10_n720, us10_n721, 
       us10_n722, us10_n723, us10_n724, us10_n725, us10_n726, us10_n727, us10_n728, us10_n729, us10_n730, 
       us10_n731, us10_n732, us10_n733, us10_n734, us10_n735, us10_n736, us10_n737, us10_n738, us10_n739, 
       us10_n740, us10_n741, us10_n742, us10_n743, us10_n744, us10_n745, us10_n746, us10_n747, us10_n748, 
       us10_n749, us10_n750, us10_n751, us10_n752, us10_n753, us10_n754, us10_n755, us10_n756, us10_n757, 
       us10_n758, us10_n759, us10_n760, us10_n761, us10_n762, us10_n763, us10_n764, us10_n765, us10_n766, 
       us10_n767, us10_n768, us10_n769, us10_n770, us10_n771, us10_n772, us10_n773, us10_n774, us10_n775, 
       us10_n776, us10_n777, us10_n778, us10_n779, us10_n780, us10_n781, us10_n782, us10_n783, us10_n784, 
       us10_n785, us10_n786, us10_n787, us10_n788, us10_n789, us10_n790, us10_n791, us10_n792, us10_n793, 
       us10_n794, us10_n795, us10_n796, us10_n797, us10_n798, us10_n799, us10_n800, us10_n801, us10_n802, 
       us10_n803, us10_n804, us10_n805, us10_n806, us10_n807, us10_n808, us10_n809, us10_n810, us10_n811, 
       us10_n812, us10_n813, us10_n814, us10_n815, us10_n816, us10_n817, us10_n818, us10_n819, us10_n820, 
       us10_n821, us10_n822, us10_n823, us10_n824, us10_n825, us10_n826, us10_n827, us10_n828, us10_n829, 
       us10_n830, us10_n831, us10_n832, us10_n833, us10_n834, us10_n835, us10_n836, us10_n837, us10_n838, 
       us10_n839, us10_n840, us10_n841, us10_n842, us10_n843, us10_n844, us10_n845, us10_n846, us10_n847, 
       us10_n848, us10_n849, us10_n850, us10_n851, us10_n852, us10_n853, us10_n854, us10_n855, us10_n856, 
       us10_n857, us10_n858, us10_n859, us10_n860, us10_n861, us10_n862, us10_n863, us10_n864, us10_n865, 
       us10_n866, us10_n867, us10_n868, us10_n869, us10_n870, us10_n871, us10_n872, us10_n873, us10_n874, 
       us10_n875,  us10_n876;
  OAI22_X1 U1073 (.ZN( N169 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n770 ) , .B1( n771 ) );
  XOR2_X1 U1074 (.Z( n771 ) , .A( n772 ) , .B( n773 ) );
  XOR2_X1 U1075 (.B( n665 ) , .Z( n773 ) , .A( sa01_sr_6 ) );
  XNOR2_X1 U1077 (.ZN( n772 ) , .B( n774 ) , .A( sa21_sr_7 ) );
  XOR2_X1 U1078 (.Z( n774 ) , .B( sa31_sr_6 ) , .A( w1_7 ) );
  XOR2_X1 U1079 (.A( n143 ) , .Z( n770 ) , .B( w1_7 ) );
  XOR2_X1 U1149 (.Z( n823 ) , .A( n824 ) , .B( n825 ) );
  OAI22_X1 U1159 (.ZN( N150 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n832 ) , .B1( n833 ) );
  XOR2_X1 U1160 (.Z( n833 ) , .A( n834 ) , .B( n835 ) );
  XOR2_X1 U1161 (.Z( n835 ) , .A( n836 ) , .B( n837 ) );
  XOR2_X1 U1162 (.Z( n834 ) , .A( n838 ) , .B( n839 ) );
  XNOR2_X1 U1163 (.ZN( n838 ) , .B( sa12_sr_4 ) , .A( w2_28 ) );
  XOR2_X1 U1164 (.A( n121 ) , .Z( n832 ) , .B( w2_28 ) );
  OAI22_X1 U1166 (.ZN( N149 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n840 ) , .B1( n841 ) );
  XOR2_X1 U1168 (.Z( n843 ) , .B( n844 ) , .A( n845 ) );
  XNOR2_X1 U1170 (.ZN( n846 ) , .B( sa12_sr_3 ) , .A( w2_27 ) );
  XOR2_X1 U1171 (.A( n119 ) , .Z( n840 ) , .B( w2_27 ) );
  OAI22_X1 U1173 (.ZN( N148 ) , .A1( n1215 ) , .B2( n1219 ) , .A2( n847 ) , .B1( n848 ) );
  XOR2_X1 U1175 (.A( n277 ) , .Z( n850 ) , .B( n851 ) );
  XOR2_X1 U1177 (.A( n117 ) , .Z( n847 ) , .B( w2_26 ) );
  OAI22_X1 U1179 (.ZN( N147 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n852 ) , .B1( n853 ) );
  XOR2_X1 U1182 (.B( n284 ) , .Z( n854 ) , .A( n857 ) );
  XNOR2_X1 U1183 (.ZN( n857 ) , .B( sa12_sr_1 ) , .A( w2_25 ) );
  XOR2_X1 U1184 (.A( n115 ) , .Z( n852 ) , .B( w2_25 ) );
  XOR2_X1 U1188 (.A( n836 ) , .Z( n861 ) , .B( n862 ) );
  OAI22_X1 U1214 (.ZN( N134 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n879 ) , .B1( n880 ) );
  XOR2_X1 U1215 (.Z( n880 ) , .A( n881 ) , .B( n882 ) );
  XOR2_X1 U1216 (.Z( n882 ) , .B( n883 ) , .A( sa12_sr_3 ) );
  XOR2_X1 U1217 (.Z( n883 ) , .B( sa22_sr_3 ) , .A( w2_20 ) );
  XOR2_X1 U1218 (.Z( n881 ) , .A( n884 ) , .B( n885 ) );
  XNOR2_X1 U1219 (.B( n839 ) , .ZN( n884 ) , .A( sa02_sr_4 ) );
  XOR2_X1 U1220 (.A( n105 ) , .Z( n879 ) , .B( w2_20 ) );
  OAI22_X1 U1222 (.ZN( N133 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n886 ) , .B1( n887 ) );
  XOR2_X1 U1223 (.Z( n887 ) , .A( n888 ) , .B( n889 ) );
  XOR2_X1 U1224 (.Z( n889 ) , .B( n890 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1225 (.Z( n890 ) , .B( sa22_sr_2 ) , .A( w2_19 ) );
  XOR2_X1 U1228 (.A( n103 ) , .Z( n886 ) , .B( w2_19 ) );
  OAI22_X1 U1230 (.ZN( N132 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n892 ) , .B1( n893 ) );
  XOR2_X1 U1233 (.Z( n896 ) , .B( sa22_sr_1 ) , .A( w2_18 ) );
  XOR2_X1 U1236 (.A( n101 ) , .Z( n892 ) , .B( w2_18 ) );
  XOR2_X1 U1242 (.B( n885 ) , .Z( n900 ) , .A( n903 ) );
  XNOR2_X1 U1243 (.B( n856 ) , .ZN( n903 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1248 (.A( n862 ) , .B( n885 ) , .Z( n907 ) );
  XOR2_X1 U1249 (.Z( n885 ) , .A( sa12_sr_7 ) , .B( sa22_sr_7 ) );
  XOR2_X1 U1255 (.A( n824 ) , .B( n836 ) , .Z( n911 ) );
  XOR2_X1 U1256 (.Z( n824 ) , .A( sa22_sr_6 ) , .B( sa32_sr_6 ) );
  XOR2_X1 U1268 (.Z( n917 ) , .A( n918 ) , .B( n919 ) );
  XOR2_X1 U1269 (.A( n825 ) , .B( n839 ) , .Z( n919 ) );
  XOR2_X1 U1270 (.Z( n839 ) , .A( sa22_sr_4 ) , .B( sa32_sr_4 ) );
  XNOR2_X1 U1271 (.ZN( n918 ) , .B( sa32_sr_5 ) , .A( w2_13 ) );
  XOR2_X1 U1276 (.A( n830 ) , .B( n844 ) , .Z( n923 ) );
  XOR2_X1 U1277 (.Z( n844 ) , .A( sa22_sr_3 ) , .B( sa32_sr_3 ) );
  INV_X1 U1278 (.ZN( n830 ) , .A( n924 ) );
  XOR2_X1 U1285 (.A( n837 ) , .B( n851 ) , .Z( n929 ) );
  INV_X1 U1287 (.ZN( n837 ) , .A( n930 ) );
  XNOR2_X1 U1289 (.ZN( n931 ) , .B( sa32_sr_3 ) , .A( w2_11 ) );
  OAI22_X1 U1292 (.ZN( N116 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n932 ) , .B1( n933 ) );
  XOR2_X1 U1294 (.A( n845 ) , .B( n856 ) , .Z( n935 ) );
  XOR2_X1 U1295 (.Z( n856 ) , .A( sa22_sr_1 ) , .B( sa32_sr_1 ) );
  XOR2_X1 U1297 (.A( n85 ) , .Z( n932 ) , .B( w2_10 ) );
  XOR2_X1 U1301 (.A( n817 ) , .B( n862 ) , .Z( n939 ) );
  XOR2_X1 U1302 (.Z( n862 ) , .A( sa22_sr_0 ) , .B( sa32_sr_0 ) );
  XOR2_X1 U1304 (.Z( n277 ) , .A( sa02_sr_1 ) , .B( sa12_sr_1 ) );
  XNOR2_X1 U1305 (.ZN( n940 ) , .B( sa32_sr_1 ) , .A( w2_9 ) );
  OAI22_X1 U1308 (.ZN( N114 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n941 ) , .B1( n942 ) );
  XOR2_X1 U1310 (.A( n284 ) , .B( n817 ) , .Z( n944 ) );
  XOR2_X1 U1311 (.Z( n817 ) , .A( sa22_sr_7 ) , .B( sa32_sr_7 ) );
  XOR2_X1 U1312 (.Z( n284 ) , .A( sa02_sr_0 ) , .B( sa12_sr_0 ) );
  XOR2_X1 U1314 (.A( n81 ) , .Z( n941 ) , .B( w2_8 ) );
  OAI22_X1 U1316 (.ZN( N105 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n945 ) , .B1( n946 ) );
  XOR2_X1 U1317 (.Z( n946 ) , .A( n947 ) , .B( n948 ) );
  XOR2_X1 U1318 (.B( n836 ) , .Z( n948 ) , .A( sa02_sr_6 ) );
  XOR2_X1 U1319 (.Z( n836 ) , .A( sa02_sr_7 ) , .B( sa12_sr_7 ) );
  XNOR2_X1 U1320 (.ZN( n947 ) , .B( n949 ) , .A( sa22_sr_7 ) );
  XOR2_X1 U1321 (.Z( n949 ) , .B( sa32_sr_6 ) , .A( w2_7 ) );
  XOR2_X1 U1322 (.A( n79 ) , .Z( n945 ) , .B( w2_7 ) );
  XNOR2_X1 U1336 (.B( n825 ) , .ZN( n957 ) , .A( sa02_sr_4 ) );
  XOR2_X1 U1337 (.Z( n825 ) , .A( sa02_sr_5 ) , .B( sa12_sr_5 ) );
  OAI22_X1 U1340 (.ZN( N102 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n960 ) , .B1( n961 ) );
  XOR2_X1 U1343 (.Z( n964 ) , .B( sa32_sr_3 ) , .A( w2_4 ) );
  XOR2_X1 U1344 (.A( n924 ) , .Z( n962 ) , .B( n965 ) );
  XOR2_X1 U1345 (.B( n279 ) , .Z( n965 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1346 (.ZN( n924 ) , .A( sa02_sr_4 ) , .B( sa12_sr_4 ) );
  XOR2_X1 U1347 (.A( n73 ) , .Z( n960 ) , .B( w2_4 ) );
  XOR2_X1 U1354 (.B( n279 ) , .Z( n971 ) , .A( sa02_sr_2 ) );
  XOR2_X1 U1355 (.Z( n279 ) , .A( sa02_sr_7 ) , .B( sa32_sr_7 ) );
  XNOR2_X1 U1356 (.ZN( n930 ) , .A( sa02_sr_3 ) , .B( sa12_sr_3 ) );
  OAI22_X1 U1359 (.ZN( N100 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n972 ) , .B1( n973 ) );
  XOR2_X1 U1361 (.Z( n973 ) , .A( n974 ) , .B( n975 ) );
  XOR2_X1 U1362 (.Z( n975 ) , .B( n976 ) , .A( sa22_sr_2 ) );
  XOR2_X1 U1363 (.Z( n976 ) , .B( sa32_sr_1 ) , .A( w2_2 ) );
  XNOR2_X1 U1364 (.B( n845 ) , .ZN( n974 ) , .A( sa02_sr_1 ) );
  XOR2_X1 U1365 (.Z( n845 ) , .B( sa02_sr_2 ) , .A( sa12_sr_2 ) );
  XOR2_X1 U1366 (.A( n69 ) , .Z( n972 ) , .B( w2_2 ) );
  CLKBUF_X1 U1368 (.Z( n1219 ) , .A( n1220 ) );
  CLKBUF_X1 U1369 (.A( n1109 ) , .Z( n1212 ) );
  XOR2_X1 U1370 (.A( n1115 ) , .Z( n382 ) , .B( n384 ) );
  XOR2_X1 U1371 (.Z( n1115 ) , .B( n386 ) , .A( w3_16 ) );
  XNOR2_X1 U1372 (.B( n1116 ) , .ZN( n338 ) , .A( sa13_sr_6 ) );
  XOR2_X1 U1373 (.Z( n1116 ) , .B( sa23_sr_6 ) , .A( w3_23 ) );
  XNOR2_X1 U1375 (.A( n1117 ) , .B( n885 ) , .ZN( n888 ) );
  XOR2_X1 U1376 (.Z( n1117 ) , .B( n844 ) , .A( sa02_sr_3 ) );
  XNOR2_X1 U1377 (.A( n1118 ) , .B( n539 ) , .ZN( n542 ) );
  XOR2_X1 U1378 (.Z( n1118 ) , .B( n496 ) , .A( sa00_sr_3 ) );
  XNOR2_X1 U1379 (.B( n476 ) , .ZN( n524 ) , .A( sa00_sr_6 ) );
  XNOR2_X1 U1380 (.B( n824 ) , .ZN( n870 ) , .A( sa02_sr_6 ) );
  XNOR2_X1 U1382 (.B( n295 ) , .ZN( n343 ) , .A( sa03_sr_6 ) );
  XNOR2_X1 U1383 (.B( n851 ) , .ZN( n894 ) , .A( sa02_sr_2 ) );
  INV_X1 U1384 (.A( n1114 ) , .ZN( n1214 ) );
  BUF_X1 U1385 (.Z( n1217 ) , .A( n1221 ) );
  XNOR2_X1 U1387 (.A( n1119 ) , .ZN( n405 ) , .B( n407 ) );
  XNOR2_X1 U1388 (.ZN( n1119 ) , .B( n289 ) , .A( n408 ) );
  XNOR2_X1 U1389 (.A( n1120 ) , .ZN( n312 ) , .B( n314 ) );
  XNOR2_X1 U1390 (.ZN( n1120 ) , .B( n307 ) , .A( n317 ) );
  XNOR2_X1 U1393 (.B( n1122 ) , .ZN( n428 ) , .A( n429 ) );
  XNOR2_X1 U1394 (.ZN( n1122 ) , .B( n431 ) , .A( sa23_sr_6 ) );
  XNOR2_X1 U1395 (.A( n1123 ) , .ZN( n388 ) , .B( n390 ) );
  XOR2_X1 U1396 (.Z( n1123 ) , .B( sa33_sr_7 ) , .A( w3_15 ) );
  XNOR2_X1 U1397 (.A( n1124 ) , .ZN( n396 ) , .B( n398 ) );
  XOR2_X1 U1398 (.Z( n1124 ) , .B( sa33_sr_5 ) , .A( w3_13 ) );
  INV_X1 U1399 (.A( n1213 ) , .ZN( n1221 ) );
  INV_X1 U1400 (.A( n1212 ) , .ZN( n1220 ) );
  XNOR2_X1 U1403 (.A( n1126 ) , .ZN( n493 ) , .B( n495 ) );
  XNOR2_X1 U1404 (.ZN( n1126 ) , .B( n488 ) , .A( n498 ) );
  XNOR2_X1 U1405 (.A( n1127 ) , .ZN( n841 ) , .B( n843 ) );
  XNOR2_X1 U1406 (.ZN( n1127 ) , .B( n836 ) , .A( n846 ) );
  XNOR2_X1 U1407 (.A( n1128 ) , .ZN( n933 ) , .B( n935 ) );
  XOR2_X1 U1408 (.Z( n1128 ) , .B( sa32_sr_2 ) , .A( w2_10 ) );
  XNOR2_X1 U1411 (.A( n1130 ) , .ZN( n848 ) , .B( n850 ) );
  XOR2_X1 U1412 (.Z( n1130 ) , .B( sa12_sr_2 ) , .A( w2_26 ) );
  XNOR2_X1 U1417 (.A( n1133 ) , .ZN( n272 ) , .B( n275 ) );
  XOR2_X1 U1418 (.Z( n1133 ) , .A( n277 ) , .B( n278 ) );
  XNOR2_X1 U1419 (.B( n1134 ) , .ZN( n433 ) , .A( n434 ) );
  XNOR2_X1 U1420 (.ZN( n1134 ) , .B( n436 ) , .A( sa23_sr_5 ) );
  XNOR2_X1 U1421 (.A( n1135 ) , .ZN( n579 ) , .B( n581 ) );
  XNOR2_X1 U1422 (.ZN( n1135 ) , .B( n469 ) , .A( n582 ) );
  XNOR2_X1 U1425 (.A( n1137 ) , .ZN( n325 ) , .B( n327 ) );
  XNOR2_X1 U1426 (.ZN( n1137 ) , .B( n307 ) , .A( n330 ) );
  XNOR2_X1 U1427 (.A( n1138 ) , .ZN( n927 ) , .B( n929 ) );
  XNOR2_X1 U1428 (.ZN( n1138 ) , .B( n817 ) , .A( n931 ) );
  XNOR2_X1 U1429 (.B( n1139 ) , .ZN( n893 ) , .A( n894 ) );
  XNOR2_X1 U1430 (.ZN( n1139 ) , .B( n896 ) , .A( sa12_sr_1 ) );
  XNOR2_X1 U1431 (.B( n1140 ) , .ZN( n445 ) , .A( n446 ) );
  XNOR2_X1 U1432 (.ZN( n1140 ) , .B( n448 ) , .A( sa23_sr_3 ) );
  XNOR2_X1 U1433 (.B( n1141 ) , .ZN( n362 ) , .A( n363 ) );
  XNOR2_X1 U1434 (.ZN( n1141 ) , .B( n365 ) , .A( sa13_sr_2 ) );
  XNOR2_X1 U1435 (.B( n1142 ) , .ZN( n369 ) , .A( n370 ) );
  XNOR2_X1 U1436 (.ZN( n1142 ) , .B( n372 ) , .A( sa13_sr_1 ) );
  XNOR2_X1 U1439 (.A( n1144 ) , .ZN( n500 ) , .B( n502 ) );
  XOR2_X1 U1440 (.Z( n1144 ) , .B( sa10_sr_2 ) , .A( w0_26 ) );
  XNOR2_X1 U1442 (.ZN( n1145 ) , .A( n930 ) , .B( n971 ) );
  XNOR2_X1 U1447 (.A( n1148 ) , .ZN( n281 ) , .B( n283 ) );
  XOR2_X1 U1448 (.Z( n1148 ) , .B( sa22_sr_0 ) , .A( w2_0 ) );
  XNOR2_X1 U1449 (.B( n1149 ) , .ZN( n619 ) , .A( n620 ) );
  XNOR2_X1 U1450 (.ZN( n1149 ) , .B( n622 ) , .A( sa20_sr_3 ) );
  XNOR2_X1 U1451 (.A( n1150 ) , .ZN( n937 ) , .B( n939 ) );
  XNOR2_X1 U1452 (.ZN( n1150 ) , .B( n277 ) , .A( n940 ) );
  XNOR2_X1 U1457 (.A( n1153 ) , .ZN( n562 ) , .B( n564 ) );
  XOR2_X1 U1458 (.Z( n1153 ) , .B( sa30_sr_7 ) , .A( w0_15 ) );
  XNOR2_X1 U1461 (.A( n1155 ) , .ZN( n473 ) , .B( n475 ) );
  XOR2_X1 U1462 (.Z( n1155 ) , .B( sa10_sr_6 ) , .A( w0_30 ) );
  XNOR2_X1 U1481 (.A( n1165 ) , .ZN( n414 ) , .B( n416 ) );
  XNOR2_X1 U1482 (.ZN( n1165 ) , .B( n289 ) , .A( n417 ) );
  XNOR2_X1 U1483 (.A( n1166 ) , .ZN( n506 ) , .B( n508 ) );
  XNOR2_X1 U1484 (.ZN( n1166 ) , .B( n488 ) , .A( n511 ) );
  XNOR2_X1 U1487 (.A( n1168 ) , .ZN( n942 ) , .B( n944 ) );
  XOR2_X1 U1488 (.Z( n1168 ) , .B( sa32_sr_0 ) , .A( w2_8 ) );
  XNOR2_X1 U1495 (.B( n1172 ) , .ZN( n853 ) , .A( n854 ) );
  XNOR2_X1 U1496 (.ZN( n1172 ) , .A( n836 ) , .B( n856 ) );
  XNOR2_X1 U1497 (.A( n1173 ) , .ZN( n905 ) , .B( n907 ) );
  XOR2_X1 U1498 (.Z( n1173 ) , .B( sa02_sr_0 ) , .A( w2_16 ) );
  XNOR2_X1 U1501 (.B( n1175 ) , .ZN( n456 ) , .A( n457 ) );
  XNOR2_X1 U1502 (.ZN( n1175 ) , .B( n459 ) , .A( sa23_sr_1 ) );
  XNOR2_X1 U1507 (.B( n1178 ) , .ZN( n625 ) , .A( n626 ) );
  XNOR2_X1 U1508 (.ZN( n1178 ) , .B( n628 ) , .A( sa20_sr_2 ) );
  XNOR2_X1 U1509 (.B( n1179 ) , .ZN( n547 ) , .A( n548 ) );
  XNOR2_X1 U1510 (.ZN( n1179 ) , .B( n550 ) , .A( sa10_sr_1 ) );
  XNOR2_X1 U1511 (.B( n1180 ) , .ZN( n375 ) , .A( n376 ) );
  XNOR2_X1 U1512 (.ZN( n1180 ) , .B( n378 ) , .A( sa13_sr_0 ) );
  XNOR2_X1 U1513 (.B( n1181 ) , .ZN( n961 ) , .A( n962 ) );
  XNOR2_X1 U1514 (.ZN( n1181 ) , .B( n964 ) , .A( sa22_sr_4 ) );
  XNOR2_X1 U1515 (.B( n1182 ) , .ZN( n342 ) , .A( n343 ) );
  XNOR2_X1 U1516 (.ZN( n1182 ) , .B( n345 ) , .A( sa13_sr_5 ) );
  XNOR2_X1 U1518 (.ZN( n1183 ) , .B( n539 ) , .A( n556 ) );
  XNOR2_X1 U1527 (.A( n1188 ) , .ZN( n630 ) , .B( n632 ) );
  XNOR2_X1 U1528 (.ZN( n1188 ) , .B( n617 ) , .A( n634 ) );
  XNOR2_X1 U1531 (.A( n1190 ) , .ZN( n419 ) , .B( n421 ) );
  XOR2_X1 U1532 (.Z( n1190 ) , .B( sa33_sr_0 ) , .A( w3_8 ) );
  XNOR2_X1 U1537 (.A( n1193 ) , .ZN( n332 ) , .B( n334 ) );
  XOR2_X1 U1538 (.Z( n1193 ) , .B( sa13_sr_0 ) , .A( w3_24 ) );
  XNOR2_X1 U1539 (.A( n1194 ) , .ZN( n593 ) , .B( n595 ) );
  XOR2_X1 U1540 (.Z( n1194 ) , .B( sa30_sr_0 ) , .A( w0_8 ) );
  XNOR2_X1 U1541 (.A( n1195 ) , .ZN( n286 ) , .B( n288 ) );
  XOR2_X1 U1542 (.Z( n1195 ) , .B( sa13_sr_7 ) , .A( w3_31 ) );
  XNOR2_X1 U1543 (.A( n1196 ) , .ZN( n584 ) , .B( n586 ) );
  XOR2_X1 U1544 (.Z( n1196 ) , .B( sa30_sr_2 ) , .A( w0_10 ) );
  XNOR2_X1 U1549 (.A( n1199 ) , .ZN( n298 ) , .B( n300 ) );
  XOR2_X1 U1550 (.Z( n1199 ) , .B( sa13_sr_5 ) , .A( w3_29 ) );
  XNOR2_X1 U1551 (.A( n1200 ) , .ZN( n319 ) , .B( n321 ) );
  XOR2_X1 U1552 (.Z( n1200 ) , .B( sa13_sr_2 ) , .A( w3_26 ) );
  XNOR2_X1 U1553 (.A( n1201 ) , .ZN( n410 ) , .B( n412 ) );
  XOR2_X1 U1554 (.Z( n1201 ) , .B( sa33_sr_2 ) , .A( w3_10 ) );
  XNOR2_X1 U1555 (.A( n1202 ) , .ZN( n462 ) , .B( n464 ) );
  XOR2_X1 U1556 (.Z( n1202 ) , .B( sa23_sr_0 ) , .A( w3_0 ) );
  XNOR2_X1 U1557 (.A( n1203 ) , .ZN( n558 ) , .B( n560 ) );
  XOR2_X1 U1558 (.Z( n1203 ) , .B( sa00_sr_0 ) , .A( w0_16 ) );
  XNOR2_X1 U1559 (.A( n1204 ) , .ZN( n636 ) , .B( n638 ) );
  XOR2_X1 U1560 (.Z( n1204 ) , .B( sa20_sr_0 ) , .A( w0_0 ) );
  XNOR2_X1 U1561 (.A( n1205 ) , .ZN( n292 ) , .B( n294 ) );
  XOR2_X1 U1562 (.Z( n1205 ) , .B( sa13_sr_6 ) , .A( w3_30 ) );
  XNOR2_X1 U1564 (.ZN( N463 ) , .B( n1208 ) , .A( w2_10 ) );
  BUF_X1 U1565 (.A( n1109 ) , .Z( n1213 ) );
  NAND2_X1 U1569 (.A2( n1209 ) , .ZN( n1210 ) , .A1( sa22_sr_2 ) );
  NAND2_X1 U1570 (.A1( n1208 ) , .ZN( n1211 ) , .A2( sa32_sr_2 ) );
  NAND2_X1 U1571 (.A1( n1210 ) , .A2( n1211 ) , .ZN( n851 ) );
  INV_X1 U1572 (.ZN( n1208 ) , .A( sa22_sr_2 ) );
  INV_X1 U1573 (.ZN( n1209 ) , .A( sa32_sr_2 ) );
  INV_X1 U1574 (.ZN( n1215 ) , .A( n1221 ) );
  INV_X1 U1575 (.ZN( n1216 ) , .A( n1221 ) );
  OAI22_X1 U276 (.ZN( N99 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n271 ) , .B1( n272 ) );
  XOR2_X1 U278 (.Z( n275 ) , .B( n276 ) , .A( sa22_sr_1 ) );
  XOR2_X1 U279 (.Z( n276 ) , .B( sa32_sr_0 ) , .A( w2_1 ) );
  XOR2_X1 U281 (.Z( n278 ) , .B( n279 ) , .A( sa02_sr_0 ) );
  XOR2_X1 U282 (.Z( n271 ) , .A( n67 ) , .B( w2_1 ) );
  OAI22_X1 U284 (.ZN( N98 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n280 ) , .B1( n281 ) );
  XOR2_X1 U286 (.A( n279 ) , .Z( n283 ) , .B( n284 ) );
  XOR2_X1 U288 (.Z( n280 ) , .A( n65 ) , .B( w2_0 ) );
  OAI22_X1 U290 (.ZN( N89 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n285 ) , .B1( n286 ) );
  XOR2_X1 U292 (.Z( n288 ) , .A( n289 ) , .B( n290 ) );
  XOR2_X1 U294 (.Z( n285 ) , .A( n63 ) , .B( w3_31 ) );
  OAI22_X1 U296 (.ZN( N88 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n291 ) , .B1( n292 ) );
  XOR2_X1 U298 (.Z( n294 ) , .A( n295 ) , .B( n296 ) );
  XOR2_X1 U300 (.Z( n291 ) , .A( n61 ) , .B( w3_30 ) );
  OAI22_X1 U302 (.ZN( N87 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n297 ) , .B1( n298 ) );
  XOR2_X1 U304 (.Z( n300 ) , .A( n301 ) , .B( n302 ) );
  XOR2_X1 U306 (.Z( n297 ) , .A( n59 ) , .B( w3_29 ) );
  OAI22_X1 U308 (.ZN( N86 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n303 ) , .B1( n304 ) );
  XOR2_X1 U309 (.Z( n304 ) , .A( n305 ) , .B( n306 ) );
  XOR2_X1 U310 (.Z( n306 ) , .A( n307 ) , .B( n308 ) );
  XOR2_X1 U311 (.Z( n305 ) , .A( n309 ) , .B( n310 ) );
  XNOR2_X1 U312 (.ZN( n309 ) , .B( sa13_sr_4 ) , .A( w3_28 ) );
  XOR2_X1 U313 (.Z( n303 ) , .A( n57 ) , .B( w3_28 ) );
  OAI22_X1 U315 (.ZN( N85 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n311 ) , .B1( n312 ) );
  XOR2_X1 U317 (.Z( n314 ) , .A( n315 ) , .B( n316 ) );
  XNOR2_X1 U319 (.ZN( n317 ) , .B( sa13_sr_3 ) , .A( w3_27 ) );
  XOR2_X1 U320 (.Z( n311 ) , .A( n55 ) , .B( w3_27 ) );
  OAI22_X1 U322 (.ZN( N84 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n318 ) , .B1( n319 ) );
  XOR2_X1 U324 (.Z( n321 ) , .A( n322 ) , .B( n323 ) );
  XOR2_X1 U326 (.Z( n318 ) , .A( n53 ) , .B( w3_26 ) );
  OAI22_X1 U328 (.ZN( N83 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n324 ) , .B1( n325 ) );
  XOR2_X1 U330 (.Z( n327 ) , .A( n328 ) , .B( n329 ) );
  XNOR2_X1 U332 (.ZN( n330 ) , .B( sa13_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U333 (.Z( n324 ) , .A( n51 ) , .B( w3_25 ) );
  OAI22_X1 U335 (.ZN( N82 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n331 ) , .B1( n332 ) );
  XOR2_X1 U337 (.A( n307 ) , .Z( n334 ) , .B( n335 ) );
  XOR2_X1 U339 (.Z( n331 ) , .A( n49 ) , .B( w3_24 ) );
  OAI22_X1 U341 (.ZN( N73 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n336 ) , .B1( n337 ) );
  XOR2_X1 U342 (.Z( n337 ) , .A( n338 ) , .B( n339 ) );
  XOR2_X1 U343 (.B( n289 ) , .Z( n339 ) , .A( sa03_sr_7 ) );
  XOR2_X1 U346 (.Z( n336 ) , .A( n47 ) , .B( w3_23 ) );
  XOR2_X1 U351 (.Z( n345 ) , .B( sa23_sr_5 ) , .A( w3_22 ) );
  XOR2_X1 U357 (.Z( n348 ) , .A( n349 ) , .B( n350 ) );
  XOR2_X1 U358 (.Z( n350 ) , .B( n351 ) , .A( sa13_sr_4 ) );
  XOR2_X1 U359 (.Z( n351 ) , .B( sa23_sr_4 ) , .A( w3_21 ) );
  XOR2_X1 U360 (.B( n301 ) , .Z( n349 ) , .A( n352 ) );
  XOR2_X1 U364 (.Z( n354 ) , .A( n355 ) , .B( n356 ) );
  XOR2_X1 U365 (.Z( n356 ) , .B( n357 ) , .A( sa13_sr_3 ) );
  XOR2_X1 U366 (.Z( n357 ) , .B( sa23_sr_3 ) , .A( w3_20 ) );
  XOR2_X1 U367 (.Z( n355 ) , .A( n358 ) , .B( n359 ) );
  XOR2_X1 U368 (.B( n310 ) , .Z( n358 ) , .A( n360 ) );
  XOR2_X1 U374 (.Z( n365 ) , .B( sa23_sr_2 ) , .A( w3_19 ) );
  XOR2_X1 U375 (.B( n359 ) , .Z( n363 ) , .A( n366 ) );
  XOR2_X1 U376 (.B( n315 ) , .Z( n366 ) , .A( n367 ) );
  OAI22_X1 U379 (.ZN( N68 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n368 ) , .B1( n369 ) );
  XOR2_X1 U382 (.Z( n372 ) , .B( sa23_sr_1 ) , .A( w3_18 ) );
  XOR2_X1 U383 (.B( n322 ) , .Z( n370 ) , .A( n373 ) );
  XOR2_X1 U384 (.Z( n368 ) , .A( n37 ) , .B( w3_18 ) );
  OAI22_X1 U386 (.ZN( N67 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n374 ) , .B1( n375 ) );
  XOR2_X1 U389 (.Z( n378 ) , .B( sa23_sr_0 ) , .A( w3_17 ) );
  XOR2_X1 U390 (.B( n359 ) , .Z( n376 ) , .A( n379 ) );
  XOR2_X1 U391 (.B( n328 ) , .Z( n379 ) , .A( n380 ) );
  XOR2_X1 U392 (.A( n35 ) , .Z( n374 ) , .B( w3_17 ) );
  OAI22_X1 U394 (.ZN( N66 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n381 ) , .B1( n382 ) );
  XOR2_X1 U396 (.A( n335 ) , .B( n359 ) , .Z( n384 ) );
  XNOR2_X1 U397 (.ZN( n359 ) , .B( n385 ) , .A( sa13_sr_7 ) );
  XOR2_X1 U399 (.A( n33 ) , .Z( n381 ) , .B( w3_16 ) );
  OAI22_X1 U401 (.ZN( N57 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n387 ) , .B1( n388 ) );
  XOR2_X1 U403 (.A( n295 ) , .B( n307 ) , .Z( n390 ) );
  XOR2_X1 U404 (.Z( n295 ) , .A( sa23_sr_6 ) , .B( sa33_sr_6 ) );
  XOR2_X1 U406 (.A( n31 ) , .Z( n387 ) , .B( w3_15 ) );
  XOR2_X1 U410 (.A( n290 ) , .B( n301 ) , .Z( n394 ) );
  XOR2_X1 U411 (.Z( n301 ) , .A( sa23_sr_5 ) , .B( sa33_sr_5 ) );
  XOR2_X1 U417 (.A( n296 ) , .B( n310 ) , .Z( n398 ) );
  XOR2_X1 U418 (.Z( n310 ) , .A( sa23_sr_4 ) , .B( sa33_sr_4 ) );
  OAI22_X1 U422 (.ZN( N54 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n399 ) , .B1( n400 ) );
  XOR2_X1 U423 (.Z( n400 ) , .A( n401 ) , .B( n402 ) );
  XOR2_X1 U424 (.A( n302 ) , .B( n315 ) , .Z( n402 ) );
  XOR2_X1 U425 (.Z( n315 ) , .A( sa23_sr_3 ) , .B( sa33_sr_3 ) );
  XOR2_X1 U426 (.B( n289 ) , .Z( n401 ) , .A( n403 ) );
  XNOR2_X1 U427 (.ZN( n403 ) , .B( sa33_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U428 (.A( n25 ) , .Z( n399 ) , .B( w3_12 ) );
  OAI22_X1 U430 (.ZN( N53 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n404 ) , .B1( n405 ) );
  XOR2_X1 U432 (.A( n308 ) , .B( n322 ) , .Z( n407 ) );
  XOR2_X1 U433 (.Z( n322 ) , .A( sa23_sr_2 ) , .B( sa33_sr_2 ) );
  XNOR2_X1 U435 (.ZN( n408 ) , .B( sa33_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U436 (.A( n23 ) , .Z( n404 ) , .B( w3_11 ) );
  OAI22_X1 U438 (.ZN( N52 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n409 ) , .B1( n410 ) );
  XOR2_X1 U440 (.A( n316 ) , .B( n328 ) , .Z( n412 ) );
  XOR2_X1 U441 (.Z( n328 ) , .A( sa23_sr_1 ) , .B( sa33_sr_1 ) );
  XOR2_X1 U443 (.A( n21 ) , .Z( n409 ) , .B( w3_10 ) );
  XOR2_X1 U447 (.A( n323 ) , .B( n335 ) , .Z( n416 ) );
  XOR2_X1 U448 (.Z( n335 ) , .A( sa23_sr_0 ) , .B( sa33_sr_0 ) );
  XNOR2_X1 U450 (.ZN( n417 ) , .B( sa33_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U461 (.A( n289 ) , .B( n329 ) , .Z( n421 ) );
  XOR2_X1 U462 (.Z( n289 ) , .A( sa23_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U524 (.Z( N441 ) , .B( sa13_sr_0 ) , .A( w3_16 ) );
  XOR2_X1 U525 (.Z( N440 ) , .B( sa13_sr_1 ) , .A( w3_17 ) );
  XOR2_X1 U526 (.Z( N439 ) , .B( sa13_sr_2 ) , .A( w3_18 ) );
  XOR2_X1 U527 (.Z( N438 ) , .B( sa13_sr_3 ) , .A( w3_19 ) );
  XOR2_X1 U528 (.Z( N437 ) , .B( sa13_sr_4 ) , .A( w3_20 ) );
  XOR2_X1 U529 (.Z( N436 ) , .B( sa13_sr_5 ) , .A( w3_21 ) );
  XOR2_X1 U530 (.Z( N435 ) , .B( sa13_sr_6 ) , .A( w3_22 ) );
  XOR2_X1 U531 (.Z( N434 ) , .B( sa13_sr_7 ) , .A( w3_23 ) );
  XOR2_X1 U535 (.Z( N430 ) , .B( sa12_sr_3 ) , .A( w2_19 ) );
  OAI22_X1 U556 (.ZN( N41 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n422 ) , .B1( n423 ) );
  XOR2_X1 U557 (.Z( n423 ) , .A( n424 ) , .B( n425 ) );
  XOR2_X1 U558 (.B( n307 ) , .Z( n425 ) , .A( sa03_sr_6 ) );
  XOR2_X1 U559 (.Z( n307 ) , .A( sa03_sr_7 ) , .B( sa13_sr_7 ) );
  XOR2_X1 U560 (.A( n385 ) , .Z( n424 ) , .B( n426 ) );
  XOR2_X1 U561 (.Z( n426 ) , .B( sa33_sr_6 ) , .A( w3_7 ) );
  INV_X1 U562 (.ZN( n385 ) , .A( sa23_sr_7 ) );
  XOR2_X1 U563 (.A( n15 ) , .Z( n422 ) , .B( w3_7 ) );
  OAI22_X1 U575 (.ZN( N40 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n427 ) , .B1( n428 ) );
  XOR2_X1 U578 (.Z( n431 ) , .B( sa33_sr_5 ) , .A( w3_6 ) );
  XOR2_X1 U579 (.B( n290 ) , .A( n352 ) , .Z( n429 ) );
  XOR2_X1 U580 (.Z( n290 ) , .A( sa03_sr_6 ) , .B( sa13_sr_6 ) );
  INV_X1 U581 (.ZN( n352 ) , .A( sa03_sr_5 ) );
  XOR2_X1 U582 (.A( n13 ) , .Z( n427 ) , .B( w3_6 ) );
  XOR2_X1 U597 (.Z( n436 ) , .B( sa33_sr_4 ) , .A( w3_5 ) );
  XOR2_X1 U598 (.B( n296 ) , .A( n360 ) , .Z( n434 ) );
  XOR2_X1 U599 (.Z( n296 ) , .A( sa03_sr_5 ) , .B( sa13_sr_5 ) );
  INV_X1 U600 (.ZN( n360 ) , .A( sa03_sr_4 ) );
  OAI22_X1 U613 (.ZN( N38 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n437 ) , .B1( n438 ) );
  XOR2_X1 U614 (.Z( n438 ) , .A( n439 ) , .B( n440 ) );
  XOR2_X1 U615 (.Z( n440 ) , .B( n441 ) , .A( sa23_sr_4 ) );
  XOR2_X1 U616 (.Z( n441 ) , .B( sa33_sr_3 ) , .A( w3_4 ) );
  XOR2_X1 U617 (.Z( n439 ) , .A( n442 ) , .B( n443 ) );
  XOR2_X1 U618 (.B( n302 ) , .A( n367 ) , .Z( n442 ) );
  XOR2_X1 U619 (.Z( n302 ) , .A( sa03_sr_4 ) , .B( sa13_sr_4 ) );
  INV_X1 U620 (.ZN( n367 ) , .A( sa03_sr_3 ) );
  XOR2_X1 U621 (.Z( n437 ) , .A( n9 ) , .B( w3_4 ) );
  OAI22_X1 U625 (.ZN( N37 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n444 ) , .B1( n445 ) );
  XOR2_X1 U628 (.Z( n448 ) , .B( sa33_sr_2 ) , .A( w3_3 ) );
  XOR2_X1 U629 (.B( n443 ) , .Z( n446 ) , .A( n449 ) );
  XOR2_X1 U630 (.B( n308 ) , .A( n373 ) , .Z( n449 ) );
  XOR2_X1 U631 (.Z( n308 ) , .A( sa03_sr_3 ) , .B( sa13_sr_3 ) );
  INV_X1 U632 (.ZN( n373 ) , .A( sa03_sr_2 ) );
  XOR2_X1 U633 (.Z( n444 ) , .A( n7 ) , .B( w3_3 ) );
  OAI22_X1 U635 (.ZN( N36 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n450 ) , .B1( n451 ) );
  XOR2_X1 U636 (.Z( n451 ) , .A( n452 ) , .B( n453 ) );
  XOR2_X1 U637 (.Z( n453 ) , .B( n454 ) , .A( sa23_sr_2 ) );
  XOR2_X1 U638 (.Z( n454 ) , .B( sa33_sr_1 ) , .A( w3_2 ) );
  XOR2_X1 U639 (.B( n316 ) , .A( n380 ) , .Z( n452 ) );
  XOR2_X1 U640 (.Z( n316 ) , .A( sa03_sr_2 ) , .B( sa13_sr_2 ) );
  INV_X1 U641 (.ZN( n380 ) , .A( sa03_sr_1 ) );
  XOR2_X1 U642 (.Z( n450 ) , .A( n5 ) , .B( w3_2 ) );
  OAI22_X1 U644 (.ZN( N35 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n455 ) , .B1( n456 ) );
  XOR2_X1 U647 (.Z( n459 ) , .B( sa33_sr_0 ) , .A( w3_1 ) );
  XOR2_X1 U648 (.B( n443 ) , .Z( n457 ) , .A( n460 ) );
  XOR2_X1 U649 (.B( n323 ) , .A( n386 ) , .Z( n460 ) );
  XOR2_X1 U650 (.Z( n323 ) , .A( sa03_sr_1 ) , .B( sa13_sr_1 ) );
  INV_X1 U651 (.ZN( n386 ) , .A( sa03_sr_0 ) );
  XOR2_X1 U652 (.A( n3 ) , .Z( n455 ) , .B( w3_1 ) );
  XOR2_X1 U656 (.A( n329 ) , .B( n443 ) , .Z( n464 ) );
  XOR2_X1 U657 (.Z( n443 ) , .A( sa03_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U658 (.Z( n329 ) , .A( sa03_sr_0 ) , .B( sa13_sr_0 ) );
  OAI22_X1 U669 (.ZN( N280 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n472 ) , .B1( n473 ) );
  XOR2_X1 U671 (.Z( n475 ) , .A( n476 ) , .B( n477 ) );
  XOR2_X1 U673 (.A( n253 ) , .Z( n472 ) , .B( w0_30 ) );
  XOR2_X1 U677 (.Z( n481 ) , .A( n482 ) , .B( n483 ) );
  OAI22_X1 U681 (.ZN( N278 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n484 ) , .B1( n485 ) );
  XOR2_X1 U682 (.Z( n485 ) , .A( n486 ) , .B( n487 ) );
  XOR2_X1 U683 (.Z( n487 ) , .A( n488 ) , .B( n489 ) );
  XOR2_X1 U684 (.Z( n486 ) , .A( n490 ) , .B( n491 ) );
  XNOR2_X1 U685 (.ZN( n490 ) , .B( sa10_sr_4 ) , .A( w0_28 ) );
  XOR2_X1 U686 (.A( n249 ) , .Z( n484 ) , .B( w0_28 ) );
  OAI22_X1 U688 (.ZN( N277 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n492 ) , .B1( n493 ) );
  XOR2_X1 U690 (.Z( n495 ) , .A( n496 ) , .B( n497 ) );
  XNOR2_X1 U692 (.ZN( n498 ) , .B( sa10_sr_3 ) , .A( w0_27 ) );
  XOR2_X1 U693 (.A( n247 ) , .Z( n492 ) , .B( w0_27 ) );
  XOR2_X1 U697 (.Z( n502 ) , .A( n503 ) , .B( n504 ) );
  XOR2_X1 U703 (.Z( n508 ) , .A( n509 ) , .B( n510 ) );
  XNOR2_X1 U705 (.ZN( n511 ) , .B( sa10_sr_1 ) , .A( w0_25 ) );
  XOR2_X1 U710 (.A( n488 ) , .Z( n515 ) , .B( n516 ) );
  XOR2_X1 U737 (.Z( n534 ) , .A( n535 ) , .B( n536 ) );
  XOR2_X1 U738 (.Z( n536 ) , .B( n537 ) , .A( sa10_sr_3 ) );
  XOR2_X1 U739 (.Z( n537 ) , .B( sa20_sr_3 ) , .A( w0_20 ) );
  XOR2_X1 U740 (.Z( n535 ) , .A( n538 ) , .B( n539 ) );
  XNOR2_X1 U741 (.B( n491 ) , .ZN( n538 ) , .A( sa00_sr_4 ) );
  OAI22_X1 U744 (.ZN( N261 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n540 ) , .B1( n541 ) );
  XOR2_X1 U745 (.Z( n541 ) , .A( n542 ) , .B( n543 ) );
  XOR2_X1 U746 (.Z( n543 ) , .B( n544 ) , .A( sa10_sr_2 ) );
  XOR2_X1 U747 (.Z( n544 ) , .B( sa20_sr_2 ) , .A( w0_19 ) );
  XOR2_X1 U750 (.A( n231 ) , .Z( n540 ) , .B( w0_19 ) );
  XOR2_X1 U755 (.Z( n550 ) , .B( sa20_sr_1 ) , .A( w0_18 ) );
  XNOR2_X1 U756 (.B( n503 ) , .ZN( n548 ) , .A( sa00_sr_2 ) );
  XNOR2_X1 U764 (.B( n509 ) , .ZN( n556 ) , .A( sa00_sr_1 ) );
  OAI22_X1 U767 (.ZN( N258 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n557 ) , .B1( n558 ) );
  XOR2_X1 U769 (.A( n516 ) , .B( n539 ) , .Z( n560 ) );
  XOR2_X1 U770 (.Z( n539 ) , .A( sa10_sr_7 ) , .B( sa20_sr_7 ) );
  XOR2_X1 U772 (.A( n225 ) , .Z( n557 ) , .B( w0_16 ) );
  XOR2_X1 U776 (.A( n476 ) , .B( n488 ) , .Z( n564 ) );
  XOR2_X1 U777 (.Z( n476 ) , .A( sa20_sr_6 ) , .B( sa30_sr_6 ) );
  XOR2_X1 U784 (.Z( n482 ) , .A( sa20_sr_5 ) , .B( sa30_sr_5 ) );
  OAI22_X1 U788 (.ZN( N247 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n569 ) , .B1( n570 ) );
  XOR2_X1 U789 (.Z( n570 ) , .A( n571 ) , .B( n572 ) );
  XOR2_X1 U790 (.A( n477 ) , .B( n491 ) , .Z( n572 ) );
  XOR2_X1 U791 (.Z( n491 ) , .A( sa20_sr_4 ) , .B( sa30_sr_4 ) );
  XNOR2_X1 U792 (.ZN( n571 ) , .B( sa30_sr_5 ) , .A( w0_13 ) );
  XOR2_X1 U793 (.A( n219 ) , .Z( n569 ) , .B( w0_13 ) );
  OAI22_X1 U795 (.ZN( N246 ) , .A1( n1213 ) , .B2( n1217 ) , .A2( n573 ) , .B1( n574 ) );
  XOR2_X1 U796 (.Z( n574 ) , .A( n575 ) , .B( n576 ) );
  XOR2_X1 U797 (.A( n483 ) , .B( n496 ) , .Z( n576 ) );
  XOR2_X1 U798 (.Z( n496 ) , .A( sa20_sr_3 ) , .B( sa30_sr_3 ) );
  XOR2_X1 U799 (.B( n469 ) , .Z( n575 ) , .A( n577 ) );
  XNOR2_X1 U800 (.ZN( n577 ) , .B( sa30_sr_4 ) , .A( w0_12 ) );
  XOR2_X1 U801 (.A( n217 ) , .Z( n573 ) , .B( w0_12 ) );
  OAI22_X1 U803 (.ZN( N245 ) , .B2( n1114 ) , .A1( n1216 ) , .A2( n578 ) , .B1( n579 ) );
  XOR2_X1 U805 (.A( n489 ) , .B( n503 ) , .Z( n581 ) );
  XOR2_X1 U806 (.Z( n503 ) , .A( sa20_sr_2 ) , .B( sa30_sr_2 ) );
  XNOR2_X1 U808 (.ZN( n582 ) , .B( sa30_sr_3 ) , .A( w0_11 ) );
  XOR2_X1 U809 (.A( n215 ) , .Z( n578 ) , .B( w0_11 ) );
  OAI22_X1 U811 (.ZN( N244 ) , .A1( n1212 ) , .B2( n1220 ) , .A2( n583 ) , .B1( n584 ) );
  XOR2_X1 U813 (.A( n497 ) , .B( n509 ) , .Z( n586 ) );
  XOR2_X1 U814 (.Z( n509 ) , .A( sa20_sr_1 ) , .B( sa30_sr_1 ) );
  XOR2_X1 U816 (.A( n213 ) , .Z( n583 ) , .B( w0_10 ) );
  XOR2_X1 U820 (.A( n504 ) , .B( n516 ) , .Z( n590 ) );
  XOR2_X1 U821 (.Z( n516 ) , .A( sa20_sr_0 ) , .B( sa30_sr_0 ) );
  OAI22_X1 U826 (.ZN( N242 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n592 ) , .B1( n593 ) );
  XOR2_X1 U828 (.A( n469 ) , .B( n510 ) , .Z( n595 ) );
  XOR2_X1 U829 (.Z( n469 ) , .A( sa20_sr_7 ) , .B( sa30_sr_7 ) );
  XOR2_X1 U831 (.A( n209 ) , .Z( n592 ) , .B( w0_8 ) );
  OAI22_X1 U833 (.ZN( N233 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n596 ) , .B1( n597 ) );
  XOR2_X1 U834 (.Z( n597 ) , .A( n598 ) , .B( n599 ) );
  XOR2_X1 U835 (.B( n488 ) , .Z( n599 ) , .A( sa00_sr_6 ) );
  XOR2_X1 U836 (.Z( n488 ) , .A( sa00_sr_7 ) , .B( sa10_sr_7 ) );
  XNOR2_X1 U837 (.ZN( n598 ) , .B( n600 ) , .A( sa20_sr_7 ) );
  XOR2_X1 U838 (.Z( n600 ) , .B( sa30_sr_6 ) , .A( w0_7 ) );
  XOR2_X1 U839 (.A( n207 ) , .Z( n596 ) , .B( w0_7 ) );
  OAI22_X1 U849 (.ZN( N231 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n606 ) , .B1( n607 ) );
  XOR2_X1 U850 (.Z( n607 ) , .A( n608 ) , .B( n609 ) );
  XOR2_X1 U851 (.Z( n609 ) , .B( n610 ) , .A( sa20_sr_5 ) );
  XOR2_X1 U852 (.Z( n610 ) , .B( sa30_sr_4 ) , .A( w0_5 ) );
  XNOR2_X1 U853 (.B( n477 ) , .ZN( n608 ) , .A( sa00_sr_4 ) );
  XOR2_X1 U854 (.Z( n477 ) , .A( sa00_sr_5 ) , .B( sa10_sr_5 ) );
  XOR2_X1 U855 (.A( n203 ) , .Z( n606 ) , .B( w0_5 ) );
  OAI22_X1 U857 (.ZN( N230 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n611 ) , .B1( n612 ) );
  XOR2_X1 U858 (.Z( n612 ) , .A( n613 ) , .B( n614 ) );
  XOR2_X1 U859 (.Z( n614 ) , .B( n615 ) , .A( sa20_sr_4 ) );
  XOR2_X1 U860 (.Z( n615 ) , .B( sa30_sr_3 ) , .A( w0_4 ) );
  XOR2_X1 U861 (.Z( n613 ) , .A( n616 ) , .B( n617 ) );
  XNOR2_X1 U862 (.B( n483 ) , .ZN( n616 ) , .A( sa00_sr_3 ) );
  XOR2_X1 U863 (.Z( n483 ) , .A( sa00_sr_4 ) , .B( sa10_sr_4 ) );
  XOR2_X1 U864 (.A( n201 ) , .Z( n611 ) , .B( w0_4 ) );
  OAI22_X1 U868 (.ZN( N229 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n618 ) , .B1( n619 ) );
  XOR2_X1 U871 (.Z( n622 ) , .B( sa30_sr_2 ) , .A( w0_3 ) );
  XOR2_X1 U872 (.B( n617 ) , .Z( n620 ) , .A( n623 ) );
  XNOR2_X1 U873 (.B( n489 ) , .ZN( n623 ) , .A( sa00_sr_2 ) );
  XOR2_X1 U874 (.Z( n489 ) , .A( sa00_sr_3 ) , .B( sa10_sr_3 ) );
  XOR2_X1 U875 (.A( n199 ) , .Z( n618 ) , .B( w0_3 ) );
  OAI22_X1 U877 (.ZN( N228 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n624 ) , .B1( n625 ) );
  XOR2_X1 U880 (.Z( n628 ) , .B( sa30_sr_1 ) , .A( w0_2 ) );
  XNOR2_X1 U881 (.B( n497 ) , .ZN( n626 ) , .A( sa00_sr_1 ) );
  XOR2_X1 U882 (.Z( n497 ) , .A( sa00_sr_2 ) , .B( sa10_sr_2 ) );
  XOR2_X1 U883 (.A( n197 ) , .Z( n624 ) , .B( w0_2 ) );
  OAI22_X1 U885 (.ZN( N227 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n629 ) , .B1( n630 ) );
  XOR2_X1 U887 (.Z( n632 ) , .B( n633 ) , .A( sa20_sr_1 ) );
  XOR2_X1 U888 (.Z( n633 ) , .B( sa30_sr_0 ) , .A( w0_1 ) );
  XNOR2_X1 U890 (.B( n504 ) , .ZN( n634 ) , .A( sa00_sr_0 ) );
  XOR2_X1 U891 (.Z( n504 ) , .A( sa00_sr_1 ) , .B( sa10_sr_1 ) );
  XOR2_X1 U892 (.A( n195 ) , .Z( n629 ) , .B( w0_1 ) );
  XOR2_X1 U896 (.A( n510 ) , .B( n617 ) , .Z( n638 ) );
  XOR2_X1 U897 (.Z( n617 ) , .A( sa00_sr_7 ) , .B( sa30_sr_7 ) );
  XOR2_X1 U898 (.Z( n510 ) , .A( sa00_sr_0 ) , .B( sa10_sr_0 ) );
  XNOR2_X1 u0_U10 (.ZN( u0_n57 ) , .B( u0_subword_3 ) , .A( w0_3 ) );
  XNOR2_X1 u0_U17 (.ZN( u0_n53 ) , .B( u0_subword_5 ) , .A( w0_5 ) );
  XNOR2_X1 u0_U183 (.ZN( u0_n61 ) , .B( u0_subword_1 ) , .A( w0_1 ) );
  XNOR2_X1 u0_U185 (.ZN( u0_n55 ) , .B( u0_subword_4 ) , .A( w0_4 ) );
  XNOR2_X1 u0_U21 (.ZN( u0_n49 ) , .B( u0_subword_7 ) , .A( w0_7 ) );
  XNOR2_X1 u0_U212 (.ZN( u0_n59 ) , .A( u0_subword_2 ) , .B( w0_2 ) );
  XNOR2_X1 u0_U248 (.ZN( u0_n63 ) , .B( u0_subword_0 ) , .A( w0_0 ) );
  NOR2_X1 u0_u3_U10 (.ZN( u0_u3_n578 ) , .A1( u0_u3_n625 ) , .A2( u0_u3_n748 ) );
  NOR2_X1 u0_u3_U100 (.ZN( u0_u3_n669 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U101 (.ZN( u0_u3_n535 ) , .A2( u0_u3_n752 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U102 (.A2( u0_u3_n711 ) , .A1( u0_u3_n765 ) , .ZN( u0_u3_n797 ) );
  OAI22_X1 u0_u3_U103 (.B1( u0_u3_n493 ) , .ZN( u0_u3_n494 ) , .A1( u0_u3_n689 ) , .A2( u0_u3_n766 ) , .B2( u0_u3_n820 ) );
  NOR3_X1 u0_u3_U104 (.ZN( u0_u3_n493 ) , .A1( u0_u3_n785 ) , .A2( u0_u3_n852 ) , .A3( u0_u3_n865 ) );
  NOR2_X1 u0_u3_U105 (.ZN( u0_u3_n509 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n765 ) );
  NOR2_X1 u0_u3_U106 (.ZN( u0_u3_n520 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n806 ) );
  OAI21_X1 u0_u3_U107 (.ZN( u0_u3_n734 ) , .A( u0_u3_n836 ) , .B2( u0_u3_n854 ) , .B1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U108 (.ZN( u0_u3_n604 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U109 (.A2( u0_u3_n711 ) , .A1( u0_u3_n753 ) , .ZN( u0_u3_n774 ) );
  NOR2_X1 u0_u3_U11 (.A1( u0_u3_n681 ) , .ZN( u0_u3_n696 ) , .A2( u0_u3_n810 ) );
  NOR2_X1 u0_u3_U110 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n670 ) , .A1( u0_u3_n753 ) );
  BUF_X2 u0_u3_U111 (.Z( u0_u3_n439 ) , .A( u0_u3_n794 ) );
  OAI21_X1 u0_u3_U112 (.ZN( u0_u3_n790 ) , .A( u0_u3_n841 ) , .B1( u0_u3_n865 ) , .B2( u0_u3_n875 ) );
  BUF_X2 u0_u3_U113 (.Z( u0_u3_n41 ) , .A( u0_u3_n700 ) );
  NOR2_X1 u0_u3_U114 (.ZN( u0_u3_n632 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U115 (.ZN( u0_u3_n512 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U116 (.ZN( u0_u3_n510 ) , .A1( u0_u3_n815 ) , .A2( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U117 (.ZN( u0_u3_n666 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U118 (.ZN( u0_u3_n546 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U119 (.ZN( u0_u3_n511 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n788 ) );
  INV_X1 u0_u3_U12 (.A( u0_u3_n683 ) , .ZN( u0_u3_n842 ) );
  NOR2_X1 u0_u3_U120 (.ZN( u0_u3_n547 ) , .A2( u0_u3_n788 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U121 (.ZN( u0_u3_n685 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U122 (.ZN( u0_u3_n572 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n765 ) , .A( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U123 (.ZN( u0_u3_n714 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U124 (.ZN( u0_u3_n532 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U125 (.ZN( u0_u3_n518 ) , .A( u0_u3_n732 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U126 (.ZN( u0_u3_n617 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n815 ) );
  INV_X1 u0_u3_U127 (.A( u0_u3_n753 ) , .ZN( u0_u3_n844 ) );
  AOI21_X1 u0_u3_U128 (.ZN( u0_u3_n594 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n788 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U129 (.ZN( u0_u3_n517 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n795 ) , .B1( u0_u3_n815 ) );
  INV_X1 u0_u3_U13 (.A( u0_u3_n650 ) , .ZN( u0_u3_n872 ) );
  AOI21_X1 u0_u3_U130 (.B1( u0_u3_n689 ) , .ZN( u0_u3_n690 ) , .A( u0_u3_n731 ) , .B2( u0_u3_n764 ) );
  INV_X1 u0_u3_U131 (.A( u0_u3_n731 ) , .ZN( u0_u3_n854 ) );
  NOR2_X1 u0_u3_U132 (.ZN( u0_u3_n571 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n765 ) );
  INV_X1 u0_u3_U133 (.A( u0_u3_n795 ) , .ZN( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U134 (.A1( u0_u3_n752 ) , .ZN( u0_u3_n770 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U135 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n618 ) , .A1( u0_u3_n788 ) );
  AOI211_X1 u0_u3_U136 (.C2( u0_u3_n440 ) , .B( u0_u3_n626 ) , .A( u0_u3_n627 ) , .ZN( u0_u3_n638 ) , .C1( u0_u3_n865 ) );
  NOR4_X1 u0_u3_U137 (.A4( u0_u3_n632 ) , .A3( u0_u3_n633 ) , .A2( u0_u3_n634 ) , .A1( u0_u3_n635 ) , .ZN( u0_u3_n636 ) );
  NOR4_X1 u0_u3_U138 (.A4( u0_u3_n629 ) , .A3( u0_u3_n630 ) , .A2( u0_u3_n631 ) , .ZN( u0_u3_n637 ) , .A1( u0_u3_n667 ) );
  INV_X1 u0_u3_U139 (.A( u0_u3_n783 ) , .ZN( u0_u3_n852 ) );
  NOR4_X1 u0_u3_U14 (.A4( u0_u3_n547 ) , .A3( u0_u3_n548 ) , .A2( u0_u3_n549 ) , .A1( u0_u3_n550 ) , .ZN( u0_u3_n551 ) );
  OAI21_X1 u0_u3_U140 (.A( u0_u3_n701 ) , .ZN( u0_u3_n705 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n807 ) );
  OAI21_X1 u0_u3_U141 (.ZN( u0_u3_n701 ) , .B2( u0_u3_n836 ) , .B1( u0_u3_n840 ) , .A( u0_u3_n862 ) );
  INV_X1 u0_u3_U142 (.A( u0_u3_n732 ) , .ZN( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U143 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n628 ) , .A1( u0_u3_n841 ) );
  INV_X1 u0_u3_U144 (.A( u0_u3_n766 ) , .ZN( u0_u3_n868 ) );
  NOR2_X1 u0_u3_U145 (.ZN( u0_u3_n473 ) , .A2( u0_u3_n782 ) , .A1( u0_u3_n818 ) );
  INV_X1 u0_u3_U146 (.A( u0_u3_n440 ) , .ZN( u0_u3_n816 ) );
  INV_X1 u0_u3_U147 (.A( u0_u3_n820 ) , .ZN( u0_u3_n846 ) );
  NAND2_X1 u0_u3_U148 (.ZN( u0_u3_n717 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n783 ) );
  INV_X1 u0_u3_U149 (.A( u0_u3_n788 ) , .ZN( u0_u3_n848 ) );
  NOR4_X1 u0_u3_U15 (.A4( u0_u3_n448 ) , .A3( u0_u3_n449 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n544 ) , .ZN( u0_u3_n709 ) );
  AOI221_X1 u0_u3_U150 (.A( u0_u3_n767 ) , .ZN( u0_u3_n777 ) , .C2( u0_u3_n813 ) , .B2( u0_u3_n838 ) , .C1( u0_u3_n857 ) , .B1( u0_u3_n868 ) );
  INV_X1 u0_u3_U151 (.A( u0_u3_n764 ) , .ZN( u0_u3_n838 ) );
  AND2_X1 u0_u3_U152 (.ZN( u0_u3_n735 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n788 ) );
  AOI221_X1 u0_u3_U153 (.A( u0_u3_n453 ) , .ZN( u0_u3_n462 ) , .C2( u0_u3_n756 ) , .B1( u0_u3_n835 ) , .C1( u0_u3_n844 ) , .B2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U154 (.ZN( u0_u3_n453 ) , .B2( u0_u3_n795 ) , .A( u0_u3_n806 ) , .B1( u0_u3_n818 ) );
  AOI211_X1 u0_u3_U155 (.A( u0_u3_n591 ) , .ZN( u0_u3_n600 ) , .B( u0_u3_n624 ) , .C1( u0_u3_n847 ) , .C2( u0_u3_n857 ) );
  OAI221_X1 u0_u3_U156 (.A( u0_u3_n730 ) , .C2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .B1( u0_u3_n733 ) , .ZN( u0_u3_n740 ) , .C1( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U157 (.A1( u0_u3_n444 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n711 ) );
  NAND2_X1 u0_u3_U158 (.A2( u0_u3_n474 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U159 (.A2( u0_u3_n463 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n783 ) );
  OR3_X1 u0_u3_U16 (.ZN( u0_u3_n449 ) , .A1( u0_u3_n531 ) , .A3( u0_u3_n580 ) , .A2( u0_u3_n877 ) );
  NAND2_X1 u0_u3_U160 (.A1( u0_u3_n458 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n806 ) );
  NAND2_X1 u0_u3_U161 (.A2( u0_u3_n451 ) , .A1( u0_u3_n463 ) , .ZN( u0_u3_n731 ) );
  NAND2_X1 u0_u3_U162 (.A1( u0_u3_n452 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n727 ) );
  NAND2_X1 u0_u3_U163 (.A2( u0_u3_n457 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U164 (.ZN( u0_u3_n456 ) , .A1( u0_u3_n829 ) , .A2( u0_u3_n830 ) );
  NAND2_X1 u0_u3_U165 (.A2( u0_u3_n467 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n815 ) );
  NAND2_X1 u0_u3_U166 (.A2( u0_u3_n451 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n732 ) );
  NAND2_X1 u0_u3_U167 (.A2( u0_u3_n452 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n766 ) );
  NAND2_X1 u0_u3_U168 (.A1( u0_u3_n454 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U169 (.A1( u0_u3_n456 ) , .A2( u0_u3_n464 ) , .ZN( u0_u3_n747 ) );
  OR4_X1 u0_u3_U17 (.A4( u0_u3_n445 ) , .A2( u0_u3_n446 ) , .A1( u0_u3_n447 ) , .ZN( u0_u3_n448 ) , .A3( u0_u3_n556 ) );
  NAND2_X1 u0_u3_U170 (.A2( u0_u3_n444 ) , .A1( u0_u3_n450 ) , .ZN( u0_u3_n787 ) );
  NAND2_X1 u0_u3_U171 (.A1( u0_u3_n454 ) , .A2( u0_u3_n457 ) , .ZN( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U172 (.A1( u0_u3_n450 ) , .A2( u0_u3_n452 ) , .ZN( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U173 (.A2( u0_u3_n456 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U174 (.A1( u0_u3_n450 ) , .A2( u0_u3_n451 ) , .ZN( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U175 (.A2( u0_u3_n464 ) , .A1( u0_u3_n465 ) , .ZN( u0_u3_n750 ) );
  NAND2_X1 u0_u3_U176 (.A1( u0_u3_n465 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n791 ) );
  NAND2_X1 u0_u3_U177 (.A2( u0_u3_n457 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n733 ) );
  NAND2_X1 u0_u3_U178 (.A1( u0_u3_n454 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n793 ) );
  AND2_X1 u0_u3_U179 (.ZN( u0_u3_n440 ) , .A1( u0_u3_n457 ) , .A2( u0_u3_n464 ) );
  INV_X1 u0_u3_U18 (.A( u0_u3_n616 ) , .ZN( u0_u3_n877 ) );
  NOR2_X1 u0_u3_U180 (.ZN( u0_u3_n452 ) , .A1( u0_u3_n850 ) , .A2( w3_28 ) );
  NAND4_X1 u0_u3_U181 (.ZN( u0_subword_1 ) , .A4( u0_u3_n598 ) , .A3( u0_u3_n599 ) , .A2( u0_u3_n600 ) , .A1( u0_u3_n601 ) );
  AOI211_X1 u0_u3_U182 (.B( u0_u3_n592 ) , .A( u0_u3_n593 ) , .ZN( u0_u3_n599 ) , .C2( u0_u3_n814 ) , .C1( u0_u3_n836 ) );
  NOR4_X1 u0_u3_U183 (.A4( u0_u3_n594 ) , .A3( u0_u3_n595 ) , .A2( u0_u3_n596 ) , .A1( u0_u3_n597 ) , .ZN( u0_u3_n598 ) );
  NOR4_X1 u0_u3_U184 (.A4( u0_u3_n737 ) , .A3( u0_u3_n738 ) , .A2( u0_u3_n739 ) , .A1( u0_u3_n740 ) , .ZN( u0_u3_n741 ) );
  AOI211_X1 u0_u3_U185 (.B( u0_u3_n728 ) , .A( u0_u3_n729 ) , .ZN( u0_u3_n742 ) , .C1( u0_u3_n845 ) , .C2( u0_u3_n857 ) );
  AOI222_X1 u0_u3_U186 (.B2( u0_u3_n641 ) , .ZN( u0_u3_n647 ) , .B1( u0_u3_n843 ) , .A1( u0_u3_n844 ) , .C2( u0_u3_n848 ) , .C1( u0_u3_n865 ) , .A2( u0_u3_n867 ) );
  NOR4_X1 u0_u3_U187 (.A4( u0_u3_n642 ) , .A3( u0_u3_n643 ) , .A2( u0_u3_n644 ) , .A1( u0_u3_n645 ) , .ZN( u0_u3_n646 ) );
  AOI221_X1 u0_u3_U188 (.A( u0_u3_n784 ) , .ZN( u0_u3_n801 ) , .C2( u0_u3_n839 ) , .B2( u0_u3_n840 ) , .B1( u0_u3_n867 ) , .C1( u0_u3_n868 ) );
  NOR4_X1 u0_u3_U189 (.A4( u0_u3_n796 ) , .A3( u0_u3_n797 ) , .A2( u0_u3_n798 ) , .A1( u0_u3_n799 ) , .ZN( u0_u3_n800 ) );
  NOR4_X1 u0_u3_U19 (.ZN( u0_u3_n478 ) , .A1( u0_u3_n534 ) , .A3( u0_u3_n571 ) , .A4( u0_u3_n603 ) , .A2( u0_u3_n645 ) );
  NAND4_X1 u0_u3_U190 (.ZN( u0_subword_0 ) , .A4( u0_u3_n504 ) , .A3( u0_u3_n505 ) , .A2( u0_u3_n506 ) , .A1( u0_u3_n507 ) );
  NOR4_X1 u0_u3_U191 (.A4( u0_u3_n501 ) , .A3( u0_u3_n502 ) , .A2( u0_u3_n503 ) , .ZN( u0_u3_n504 ) , .A1( u0_u3_n530 ) );
  AOI221_X1 u0_u3_U192 (.A( u0_u3_n500 ) , .ZN( u0_u3_n505 ) , .B2( u0_u3_n845 ) , .C1( u0_u3_n848 ) , .C2( u0_u3_n862 ) , .B1( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U193 (.A4( u0_u3_n703 ) , .A3( u0_u3_n704 ) , .A2( u0_u3_n705 ) , .A1( u0_u3_n706 ) , .ZN( u0_u3_n707 ) );
  NOR4_X1 u0_u3_U194 (.A3( u0_u3_n758 ) , .A2( u0_u3_n759 ) , .A1( u0_u3_n760 ) , .ZN( u0_u3_n761 ) , .A4( u0_u3_n871 ) );
  AOI211_X1 u0_u3_U195 (.B( u0_u3_n748 ) , .A( u0_u3_n749 ) , .ZN( u0_u3_n762 ) , .C1( u0_u3_n835 ) , .C2( u0_u3_n855 ) );
  NAND4_X1 u0_u3_U196 (.ZN( u0_subword_7 ) , .A4( u0_u3_n825 ) , .A3( u0_u3_n826 ) , .A2( u0_u3_n827 ) , .A1( u0_u3_n828 ) );
  NOR4_X1 u0_u3_U197 (.A4( u0_u3_n821 ) , .A3( u0_u3_n822 ) , .A2( u0_u3_n823 ) , .A1( u0_u3_n824 ) , .ZN( u0_u3_n825 ) );
  NAND2_X1 u0_u3_U198 (.A2( u0_u3_n464 ) , .A1( u0_u3_n474 ) , .ZN( u0_u3_n700 ) );
  NAND2_X1 u0_u3_U199 (.A2( u0_u3_n451 ) , .A1( u0_u3_n467 ) , .ZN( u0_u3_n818 ) );
  INV_X1 u0_u3_U20 (.A( u0_u3_n752 ) , .ZN( u0_u3_n865 ) );
  OAI21_X1 u0_u3_U200 (.B1( u0_u3_n756 ) , .ZN( u0_u3_n757 ) , .A( u0_u3_n847 ) , .B2( u0_u3_n870 ) );
  AOI221_X1 u0_u3_U201 (.A( u0_u3_n567 ) , .C2( u0_u3_n568 ) , .ZN( u0_u3_n577 ) , .B2( u0_u3_n847 ) , .B1( u0_u3_n854 ) , .C1( u0_u3_n855 ) );
  AOI222_X1 u0_u3_U202 (.ZN( u0_u3_n663 ) , .A2( u0_u3_n841 ) , .B1( u0_u3_n843 ) , .C2( u0_u3_n847 ) , .A1( u0_u3_n862 ) , .C1( u0_u3_n865 ) , .B2( u0_u3_n872 ) );
  AOI221_X1 u0_u3_U203 (.A( u0_u3_n713 ) , .ZN( u0_u3_n724 ) , .C2( u0_u3_n846 ) , .B2( u0_u3_n847 ) , .C1( u0_u3_n863 ) , .B1( u0_u3_n864 ) );
  NAND4_X1 u0_u3_U204 (.A4( u0_u3_n538 ) , .A3( u0_u3_n539 ) , .A2( u0_u3_n540 ) , .A1( u0_u3_n541 ) , .ZN( u0_u3_n625 ) );
  NOR4_X1 u0_u3_U205 (.A1( u0_u3_n534 ) , .ZN( u0_u3_n539 ) , .A2( u0_u3_n657 ) , .A4( u0_u3_n671 ) , .A3( u0_u3_n768 ) );
  NAND4_X1 u0_u3_U206 (.A4( u0_u3_n496 ) , .A3( u0_u3_n497 ) , .A1( u0_u3_n498 ) , .ZN( u0_u3_n805 ) , .A2( u0_u3_n869 ) );
  NOR4_X1 u0_u3_U207 (.A2( u0_u3_n494 ) , .A1( u0_u3_n495 ) , .ZN( u0_u3_n496 ) , .A3( u0_u3_n583 ) , .A4( u0_u3_n615 ) );
  NAND2_X1 u0_u3_U208 (.A1( u0_u3_n444 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n702 ) );
  NAND2_X1 u0_u3_U209 (.A1( u0_u3_n455 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n672 ) );
  AOI222_X1 u0_u3_U21 (.ZN( u0_u3_n566 ) , .B1( u0_u3_n833 ) , .C1( u0_u3_n843 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n856 ) , .B2( u0_u3_n865 ) , .C2( u0_u3_n875 ) );
  NAND4_X1 u0_u3_U210 (.A4( u0_u3_n563 ) , .A3( u0_u3_n564 ) , .A2( u0_u3_n565 ) , .A1( u0_u3_n566 ) , .ZN( u0_u3_n610 ) );
  NOR4_X1 u0_u3_U211 (.ZN( u0_u3_n564 ) , .A1( u0_u3_n656 ) , .A3( u0_u3_n664 ) , .A4( u0_u3_n688 ) , .A2( u0_u3_n771 ) );
  NOR2_X1 u0_u3_U212 (.ZN( u0_u3_n454 ) , .A1( u0_u3_n831 ) , .A2( u0_u3_n832 ) );
  INV_X1 u0_u3_U213 (.ZN( u0_u3_n831 ) , .A( w3_26 ) );
  NOR2_X1 u0_u3_U214 (.ZN( u0_u3_n710 ) , .A2( u0_u3_n779 ) , .A1( u0_u3_n803 ) );
  OAI21_X1 u0_u3_U215 (.A( u0_u3_n734 ) , .B1( u0_u3_n735 ) , .ZN( u0_u3_n739 ) , .B2( u0_u3_n808 ) );
  AOI21_X1 u0_u3_U216 (.ZN( u0_u3_n653 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n795 ) , .B2( u0_u3_n808 ) );
  INV_X1 u0_u3_U217 (.A( u0_u3_n808 ) , .ZN( u0_u3_n862 ) );
  NOR2_X1 u0_u3_U218 (.ZN( u0_u3_n738 ) , .A2( u0_u3_n806 ) , .A1( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U219 (.ZN( u0_u3_n756 ) , .A1( u0_u3_n766 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U22 (.ZN( u0_u3_n482 ) , .A1( u0_u3_n523 ) , .A4( u0_u3_n560 ) , .A3( u0_u3_n585 ) , .A2( u0_u3_n633 ) );
  NOR2_X1 u0_u3_U220 (.ZN( u0_u3_n559 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n808 ) );
  OAI221_X1 u0_u3_U221 (.A( u0_u3_n699 ) , .ZN( u0_u3_n706 ) , .C2( u0_u3_n787 ) , .C1( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .B2( u0_u3_n809 ) );
  OAI222_X1 u0_u3_U222 (.B1( u0_u3_n41 ) , .ZN( u0_u3_n620 ) , .C1( u0_u3_n727 ) , .C2( u0_u3_n750 ) , .B2( u0_u3_n789 ) , .A2( u0_u3_n795 ) , .A1( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U223 (.A2( u0_u3_n444 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n794 ) );
  OAI222_X1 u0_u3_U224 (.B2( u0_u3_n711 ) , .ZN( u0_u3_n712 ) , .C2( u0_u3_n727 ) , .B1( u0_u3_n750 ) , .A1( u0_u3_n809 ) , .C1( u0_u3_n817 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U225 (.A( u0_u3_n675 ) , .ZN( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U226 (.ZN( u0_u3_n531 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U227 (.ZN( u0_u3_n529 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n753 ) );
  INV_X1 u0_u3_U228 (.A( u0_u3_n727 ) , .ZN( u0_u3_n858 ) );
  NOR2_X1 u0_u3_U229 (.ZN( u0_u3_n450 ) , .A2( u0_u3_n851 ) , .A1( u0_u3_n860 ) );
  NOR4_X1 u0_u3_U23 (.A4( u0_u3_n559 ) , .A3( u0_u3_n560 ) , .A2( u0_u3_n561 ) , .A1( u0_u3_n562 ) , .ZN( u0_u3_n563 ) );
  AOI222_X1 u0_u3_U230 (.ZN( u0_u3_n528 ) , .A1( u0_u3_n837 ) , .B2( u0_u3_n839 ) , .C1( u0_u3_n846 ) , .C2( u0_u3_n852 ) , .A2( u0_u3_n854 ) , .B1( u0_u3_n868 ) );
  NOR3_X1 u0_u3_U231 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n443 ) , .A3( u0_u3_n839 ) , .A1( u0_u3_n848 ) );
  NAND2_X1 u0_u3_U232 (.ZN( u0_u3_n616 ) , .A2( u0_u3_n839 ) , .A1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U233 (.ZN( u0_u3_n498 ) , .A1( u0_u3_n681 ) , .A2( u0_u3_n697 ) );
  AOI211_X1 u0_u3_U234 (.B( u0_u3_n697 ) , .A( u0_u3_n698 ) , .ZN( u0_u3_n708 ) , .C2( u0_u3_n834 ) , .C1( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U235 (.ZN( u0_u3_n586 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U236 (.ZN( u0_u3_n543 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n782 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U237 (.ZN( u0_u3_n612 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U238 (.ZN( u0_u3_n718 ) , .A1( u0_u3_n808 ) , .A2( u0_u3_n820 ) );
  OAI21_X1 u0_u3_U239 (.A( u0_u3_n790 ) , .B2( u0_u3_n791 ) , .B1( u0_u3_n792 ) , .ZN( u0_u3_n798 ) );
  NOR4_X1 u0_u3_U24 (.A4( u0_u3_n555 ) , .A3( u0_u3_n556 ) , .A2( u0_u3_n557 ) , .A1( u0_u3_n558 ) , .ZN( u0_u3_n565 ) );
  AOI21_X1 u0_u3_U240 (.ZN( u0_u3_n642 ) , .B2( u0_u3_n752 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U241 (.A( u0_u3_n736 ) , .ZN( u0_u3_n737 ) , .B2( u0_u3_n783 ) , .B1( u0_u3_n795 ) );
  AOI21_X1 u0_u3_U242 (.B2( u0_u3_n766 ) , .ZN( u0_u3_n767 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U243 (.ZN( u0_u3_n521 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U244 (.ZN( u0_u3_n487 ) , .A1( u0_u3_n791 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U245 (.ZN( u0_u3_n537 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n791 ) );
  INV_X1 u0_u3_U246 (.A( u0_u3_n791 ) , .ZN( u0_u3_n847 ) );
  OAI22_X1 u0_u3_U247 (.B2( u0_u3_n782 ) , .B1( u0_u3_n783 ) , .ZN( u0_u3_n784 ) , .A2( u0_u3_n817 ) , .A1( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U248 (.ZN( u0_u3_n501 ) , .A( u0_u3_n727 ) , .B2( u0_u3_n765 ) , .B1( u0_u3_n817 ) );
  NAND4_X1 u0_u3_U249 (.A4( u0_u3_n482 ) , .A3( u0_u3_n483 ) , .A2( u0_u3_n484 ) , .A1( u0_u3_n485 ) , .ZN( u0_u3_n697 ) );
  NOR4_X1 u0_u3_U25 (.A4( u0_u3_n771 ) , .A3( u0_u3_n772 ) , .A2( u0_u3_n773 ) , .A1( u0_u3_n774 ) , .ZN( u0_u3_n775 ) );
  AOI21_X1 u0_u3_U250 (.ZN( u0_u3_n542 ) , .B2( u0_u3_n815 ) , .A( u0_u3_n817 ) , .B1( u0_u3_n818 ) );
  NOR2_X1 u0_u3_U251 (.ZN( u0_u3_n523 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U252 (.ZN( u0_u3_n549 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n817 ) );
  INV_X1 u0_u3_U253 (.A( u0_u3_n817 ) , .ZN( u0_u3_n836 ) );
  NOR2_X1 u0_u3_U254 (.ZN( u0_u3_n548 ) , .A1( u0_u3_n752 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U255 (.ZN( u0_u3_n560 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U256 (.A( u0_u3_n673 ) , .B1( u0_u3_n674 ) , .ZN( u0_u3_n675 ) , .B2( u0_u3_n858 ) );
  AOI22_X1 u0_u3_U257 (.A2( u0_u3_n785 ) , .ZN( u0_u3_n786 ) , .B2( u0_u3_n834 ) , .A1( u0_u3_n837 ) , .B1( u0_u3_n865 ) );
  AOI21_X1 u0_u3_U258 (.ZN( u0_u3_n643 ) , .B2( u0_u3_n750 ) , .A( u0_u3_n795 ) , .B1( u0_u3_n806 ) );
  NAND4_X1 u0_u3_U259 (.A4( u0_u3_n775 ) , .A3( u0_u3_n776 ) , .A2( u0_u3_n777 ) , .A1( u0_u3_n778 ) , .ZN( u0_u3_n804 ) );
  NOR3_X1 u0_u3_U26 (.A3( u0_u3_n768 ) , .A2( u0_u3_n769 ) , .A1( u0_u3_n770 ) , .ZN( u0_u3_n776 ) );
  OAI21_X1 u0_u3_U260 (.ZN( u0_u3_n466 ) , .B1( u0_u3_n812 ) , .A( u0_u3_n837 ) , .B2( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U261 (.ZN( u0_u3_n659 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U262 (.ZN( u0_u3_n683 ) , .A2( u0_u3_n837 ) , .A1( u0_u3_n841 ) );
  NOR2_X1 u0_u3_U263 (.ZN( u0_u3_n764 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n837 ) );
  NOR2_X1 u0_u3_U264 (.ZN( u0_u3_n570 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U265 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n633 ) , .A1( u0_u3_n750 ) );
  INV_X1 u0_u3_U266 (.A( u0_u3_n750 ) , .ZN( u0_u3_n837 ) );
  NOR4_X1 u0_u3_U267 (.ZN( u0_u3_n488 ) , .A2( u0_u3_n536 ) , .A1( u0_u3_n561 ) , .A3( u0_u3_n634 ) , .A4( u0_u3_n721 ) );
  NAND4_X1 u0_u3_U268 (.A4( u0_u3_n488 ) , .A3( u0_u3_n489 ) , .A2( u0_u3_n490 ) , .A1( u0_u3_n491 ) , .ZN( u0_u3_n781 ) );
  AOI21_X1 u0_u3_U269 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n592 ) , .B2( u0_u3_n702 ) , .A( u0_u3_n820 ) );
  NAND4_X1 u0_u3_U27 (.A4( u0_u3_n606 ) , .A3( u0_u3_n607 ) , .A2( u0_u3_n608 ) , .A1( u0_u3_n609 ) , .ZN( u0_u3_n725 ) );
  AOI21_X1 u0_u3_U270 (.B1( u0_u3_n702 ) , .ZN( u0_u3_n703 ) , .A( u0_u3_n735 ) , .B2( u0_u3_n766 ) );
  INV_X1 u0_u3_U271 (.A( u0_u3_n702 ) , .ZN( u0_u3_n855 ) );
  AOI21_X1 u0_u3_U272 (.ZN( u0_u3_n445 ) , .A( u0_u3_n702 ) , .B1( u0_u3_n736 ) , .B2( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U273 (.ZN( u0_u3_n686 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U274 (.ZN( u0_u3_n580 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U275 (.A1( u0_u3_n702 ) , .A2( u0_u3_n732 ) , .ZN( u0_u3_n785 ) );
  NOR3_X1 u0_u3_U276 (.A3( u0_u3_n744 ) , .A2( u0_u3_n745 ) , .A1( u0_u3_n746 ) , .ZN( u0_u3_n763 ) );
  OAI22_X1 u0_u3_U277 (.ZN( u0_u3_n492 ) , .A1( u0_u3_n727 ) , .B2( u0_u3_n731 ) , .B1( u0_u3_n733 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U278 (.ZN( u0_u3_n582 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n733 ) );
  NOR2_X1 u0_u3_U279 (.ZN( u0_u3_n536 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n733 ) );
  NOR3_X1 u0_u3_U28 (.A1( u0_u3_n602 ) , .ZN( u0_u3_n607 ) , .A3( u0_u3_n666 ) , .A2( u0_u3_n773 ) );
  AOI222_X1 u0_u3_U280 (.ZN( u0_u3_n608 ) , .B2( u0_u3_n674 ) , .B1( u0_u3_n756 ) , .C2( u0_u3_n834 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n864 ) , .C1( u0_u3_n865 ) );
  AOI221_X1 u0_u3_U281 (.A( u0_u3_n486 ) , .ZN( u0_u3_n491 ) , .B1( u0_u3_n834 ) , .C2( u0_u3_n846 ) , .C1( u0_u3_n854 ) , .B2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U282 (.ZN( u0_u3_n792 ) , .A2( u0_u3_n864 ) , .A1( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U283 (.ZN( u0_u3_n464 ) , .A1( u0_u3_n832 ) , .A2( w3_26 ) );
  NOR2_X1 u0_u3_U284 (.ZN( u0_u3_n474 ) , .A1( u0_u3_n829 ) , .A2( w3_25 ) );
  AOI21_X1 u0_u3_U285 (.A( u0_u3_n439 ) , .ZN( u0_u3_n644 ) , .B1( u0_u3_n683 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U286 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n500 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n807 ) );
  OAI22_X1 u0_u3_U287 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n698 ) , .A2( u0_u3_n733 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U288 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n567 ) , .B1( u0_u3_n727 ) , .A( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U289 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n446 ) , .B1( u0_u3_n792 ) , .A( u0_u3_n817 ) );
  NOR4_X1 u0_u3_U29 (.A3( u0_u3_n603 ) , .A2( u0_u3_n604 ) , .A1( u0_u3_n605 ) , .ZN( u0_u3_n606 ) , .A4( u0_u3_n658 ) );
  NOR2_X1 u0_u3_U290 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n667 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U291 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n558 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U292 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n562 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U293 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n645 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U294 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n545 ) , .A1( u0_u3_n765 ) );
  INV_X1 u0_u3_U295 (.A( u0_u3_n794 ) , .ZN( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U296 (.ZN( u0_u3_n463 ) , .A1( u0_u3_n851 ) , .A2( w3_31 ) );
  AOI21_X1 u0_u3_U297 (.B2( u0_u3_n439 ) , .A( u0_u3_n793 ) , .B1( u0_u3_n795 ) , .ZN( u0_u3_n796 ) );
  AOI222_X1 u0_u3_U298 (.C2( u0_u3_n812 ) , .B2( u0_u3_n813 ) , .A2( u0_u3_n814 ) , .ZN( u0_u3_n826 ) , .C1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .B1( u0_u3_n855 ) );
  AOI22_X1 u0_u3_U299 (.ZN( u0_u3_n730 ) , .B1( u0_u3_n835 ) , .A2( u0_u3_n840 ) , .A1( u0_u3_n865 ) , .B2( u0_u3_n868 ) );
  BUF_X1 u0_u3_U3 (.Z( u0_u3_n438 ) , .A( u0_u3_n818 ) );
  NOR4_X1 u0_u3_U30 (.A4( u0_u3_n487 ) , .ZN( u0_u3_n490 ) , .A1( u0_u3_n569 ) , .A2( u0_u3_n584 ) , .A3( u0_u3_n605 ) );
  AOI222_X1 u0_u3_U300 (.ZN( u0_u3_n516 ) , .C1( u0_u3_n835 ) , .B2( u0_u3_n839 ) , .A2( u0_u3_n845 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n865 ) , .A1( u0_u3_n868 ) );
  AOI222_X1 u0_u3_U301 (.ZN( u0_u3_n472 ) , .B1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n853 ) , .A2( u0_u3_n857 ) , .B2( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U302 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n658 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U303 (.ZN( u0_u3_n715 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U304 (.ZN( u0_u3_n689 ) , .A1( u0_u3_n834 ) , .A2( u0_u3_n835 ) );
  NOR2_X1 u0_u3_U305 (.ZN( u0_u3_n524 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U306 (.ZN( u0_u3_n664 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U307 (.ZN( u0_u3_n736 ) , .A2( u0_u3_n835 ) , .A1( u0_u3_n847 ) );
  NOR2_X1 u0_u3_U308 (.ZN( u0_u3_n671 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U309 (.ZN( u0_u3_n673 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U31 (.ZN( u0_u3_n489 ) , .A1( u0_u3_n510 ) , .A2( u0_u3_n522 ) , .A4( u0_u3_n549 ) , .A3( u0_u3_n614 ) );
  INV_X1 u0_u3_U310 (.A( u0_u3_n793 ) , .ZN( u0_u3_n835 ) );
  AOI21_X1 u0_u3_U311 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n513 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n733 ) );
  AOI21_X1 u0_u3_U312 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n629 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n793 ) );
  INV_X1 u0_u3_U313 (.A( u0_u3_n672 ) , .ZN( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U314 (.ZN( u0_u3_n655 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U315 (.ZN( u0_u3_n631 ) , .A2( u0_u3_n672 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U316 (.ZN( u0_u3_n605 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U317 (.ZN( u0_u3_n530 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U318 (.ZN( u0_u3_n584 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U319 (.ZN( u0_u3_n444 ) , .A2( w3_28 ) , .A1( w3_29 ) );
  NOR4_X1 u0_u3_U32 (.A4( u0_u3_n529 ) , .A2( u0_u3_n530 ) , .A1( u0_u3_n531 ) , .ZN( u0_u3_n541 ) , .A3( u0_u3_n704 ) );
  NOR2_X1 u0_u3_U320 (.ZN( u0_u3_n468 ) , .A2( u0_u3_n849 ) , .A1( u0_u3_n850 ) );
  OAI222_X1 u0_u3_U321 (.B2( u0_u3_n750 ) , .B1( u0_u3_n751 ) , .A2( u0_u3_n752 ) , .ZN( u0_u3_n760 ) , .C2( u0_u3_n808 ) , .C1( u0_u3_n817 ) , .A1( u0_u3_n820 ) );
  INV_X1 u0_u3_U322 (.A( u0_u3_n789 ) , .ZN( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U323 (.A4( u0_u3_n617 ) , .A3( u0_u3_n618 ) , .A1( u0_u3_n619 ) , .A2( u0_u3_n620 ) , .ZN( u0_u3_n621 ) );
  INV_X1 u0_u3_U324 (.ZN( u0_u3_n830 ) , .A( w3_25 ) );
  OAI22_X1 u0_u3_U325 (.B2( u0_u3_n753 ) , .B1( u0_u3_n754 ) , .A1( u0_u3_n755 ) , .ZN( u0_u3_n759 ) , .A2( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U326 (.B2( u0_u3_n806 ) , .B1( u0_u3_n807 ) , .A2( u0_u3_n808 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n811 ) );
  AOI21_X1 u0_u3_U327 (.ZN( u0_u3_n692 ) , .B2( u0_u3_n752 ) , .B1( u0_u3_n766 ) , .A( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U328 (.A2( u0_u3_n765 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n813 ) );
  NOR2_X1 u0_u3_U329 (.ZN( u0_u3_n573 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n809 ) );
  NOR4_X1 u0_u3_U33 (.A4( u0_u3_n535 ) , .A3( u0_u3_n536 ) , .A2( u0_u3_n537 ) , .ZN( u0_u3_n538 ) , .A1( u0_u3_n823 ) );
  NOR2_X1 u0_u3_U330 (.ZN( u0_u3_n614 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U331 (.ZN( u0_u3_n486 ) , .A1( u0_u3_n711 ) , .B2( u0_u3_n788 ) , .A2( u0_u3_n809 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U332 (.ZN( u0_u3_n480 ) , .A( u0_u3_n672 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n809 ) );
  INV_X1 u0_u3_U333 (.A( u0_u3_n809 ) , .ZN( u0_u3_n843 ) );
  OAI221_X1 u0_u3_U334 (.A( u0_u3_n786 ) , .C2( u0_u3_n787 ) , .B2( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .ZN( u0_u3_n799 ) , .C1( u0_u3_n816 ) );
  NAND2_X1 u0_u3_U335 (.A1( u0_u3_n732 ) , .A2( u0_u3_n787 ) , .ZN( u0_u3_n814 ) );
  OAI22_X1 u0_u3_U336 (.ZN( u0_u3_n591 ) , .A2( u0_u3_n750 ) , .B2( u0_u3_n765 ) , .A1( u0_u3_n766 ) , .B1( u0_u3_n787 ) );
  AOI21_X1 u0_u3_U337 (.ZN( u0_u3_n595 ) , .B1( u0_u3_n731 ) , .B2( u0_u3_n787 ) , .A( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U338 (.ZN( u0_u3_n807 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U339 (.ZN( u0_u3_n626 ) , .B1( u0_u3_n702 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U34 (.A4( u0_u3_n532 ) , .A3( u0_u3_n533 ) , .ZN( u0_u3_n540 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n797 ) );
  NAND2_X2 u0_u3_U340 (.A1( u0_u3_n458 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n753 ) );
  AOI222_X1 u0_u3_U341 (.ZN( u0_u3_n778 ) , .A1( u0_u3_n833 ) , .C1( u0_u3_n837 ) , .B2( u0_u3_n843 ) , .A2( u0_u3_n852 ) , .B1( u0_u3_n863 ) , .C2( u0_u3_n875 ) );
  AOI222_X1 u0_u3_U342 (.ZN( u0_u3_n609 ) , .A1( u0_u3_n833 ) , .C2( u0_u3_n839 ) , .B1( u0_u3_n844 ) , .A2( u0_u3_n858 ) , .B2( u0_u3_n863 ) , .C1( u0_u3_n870 ) );
  AOI21_X1 u0_u3_U343 (.ZN( u0_u3_n651 ) , .A( u0_u3_n765 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n795 ) );
  OAI22_X1 u0_u3_U344 (.ZN( u0_u3_n684 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n733 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U345 (.ZN( u0_u3_n654 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U346 (.ZN( u0_u3_n751 ) , .A1( u0_u3_n863 ) , .A2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U347 (.ZN( u0_u3_n455 ) , .A1( u0_u3_n860 ) , .A2( w3_30 ) );
  NOR2_X1 u0_u3_U348 (.ZN( u0_u3_n467 ) , .A2( w3_30 ) , .A1( w3_31 ) );
  AND2_X1 u0_u3_U349 (.ZN( u0_u3_n441 ) , .A2( u0_u3_n834 ) , .A1( u0_u3_n856 ) );
  NOR3_X1 u0_u3_U35 (.A3( u0_u3_n803 ) , .A2( u0_u3_n804 ) , .A1( u0_u3_n805 ) , .ZN( u0_u3_n828 ) );
  AND2_X1 u0_u3_U350 (.ZN( u0_u3_n442 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U351 (.A3( u0_u3_n441 ) , .A2( u0_u3_n442 ) , .A1( u0_u3_n579 ) , .ZN( u0_u3_n590 ) );
  INV_X1 u0_u3_U352 (.A( u0_u3_n815 ) , .ZN( u0_u3_n856 ) );
  INV_X1 u0_u3_U353 (.A( u0_u3_n787 ) , .ZN( u0_u3_n863 ) );
  INV_X1 u0_u3_U354 (.A( u0_u3_n806 ) , .ZN( u0_u3_n845 ) );
  INV_X1 u0_u3_U355 (.A( u0_u3_n41 ) , .ZN( u0_u3_n840 ) );
  NOR2_X1 u0_u3_U356 (.A1( u0_u3_n41 ) , .ZN( u0_u3_n773 ) , .A2( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U357 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n574 ) , .B1( u0_u3_n809 ) , .A( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U358 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n665 ) , .A1( u0_u3_n732 ) );
  NOR2_X1 u0_u3_U359 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n635 ) , .A1( u0_u3_n727 ) );
  NAND4_X1 u0_u3_U36 (.A4( u0_u3_n660 ) , .A3( u0_u3_n661 ) , .A2( u0_u3_n662 ) , .A1( u0_u3_n663 ) , .ZN( u0_u3_n803 ) );
  NOR2_X1 u0_u3_U360 (.A2( u0_u3_n41 ) , .A1( u0_u3_n783 ) , .ZN( u0_u3_n823 ) );
  AOI21_X1 u0_u3_U361 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n481 ) , .A( u0_u3_n752 ) , .B1( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U362 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n569 ) , .A1( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U363 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n719 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U364 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n597 ) , .A1( u0_u3_n731 ) );
  AOI21_X1 u0_u3_U365 (.A( u0_u3_n41 ) , .ZN( u0_u3_n555 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U366 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n544 ) , .A1( u0_u3_n702 ) );
  NOR2_X1 u0_u3_U367 (.ZN( u0_u3_n583 ) , .A2( u0_u3_n700 ) , .A1( u0_u3_n794 ) );
  NOR4_X1 u0_u3_U368 (.A4( u0_u3_n779 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n781 ) , .ZN( u0_u3_n802 ) , .A2( u0_u3_n804 ) );
  NAND4_X1 u0_u3_U369 (.A4( u0_u3_n694 ) , .A3( u0_u3_n695 ) , .A1( u0_u3_n696 ) , .ZN( u0_u3_n779 ) , .A2( u0_u3_n874 ) );
  NOR3_X1 u0_u3_U37 (.A3( u0_u3_n654 ) , .A2( u0_u3_n655 ) , .A1( u0_u3_n656 ) , .ZN( u0_u3_n661 ) );
  AOI21_X1 u0_u3_U370 (.ZN( u0_u3_n596 ) , .B1( u0_u3_n753 ) , .A( u0_u3_n795 ) , .B2( u0_u3_n816 ) );
  AOI21_X1 u0_u3_U371 (.A( u0_u3_n815 ) , .B2( u0_u3_n816 ) , .B1( u0_u3_n817 ) , .ZN( u0_u3_n822 ) );
  OAI222_X1 u0_u3_U372 (.ZN( u0_u3_n508 ) , .C2( u0_u3_n628 ) , .B2( u0_u3_n650 ) , .B1( u0_u3_n750 ) , .A2( u0_u3_n751 ) , .C1( u0_u3_n808 ) , .A1( u0_u3_n809 ) );
  AOI21_X1 u0_u3_U373 (.B1( u0_u3_n628 ) , .ZN( u0_u3_n630 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U374 (.ZN( u0_u3_n652 ) , .B1( u0_u3_n732 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n816 ) );
  OAI21_X1 u0_u3_U375 (.A( u0_u3_n616 ) , .ZN( u0_u3_n619 ) , .B1( u0_u3_n628 ) , .B2( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U376 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n769 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U377 (.A2( u0_u3_n816 ) , .A1( u0_u3_n818 ) , .ZN( u0_u3_n824 ) );
  NOR2_X1 u0_u3_U378 (.ZN( u0_u3_n581 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U379 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n687 ) , .A2( u0_u3_n816 ) );
  NOR3_X1 u0_u3_U38 (.A3( u0_u3_n651 ) , .A2( u0_u3_n652 ) , .A1( u0_u3_n653 ) , .ZN( u0_u3_n662 ) );
  NOR2_X1 u0_u3_U380 (.ZN( u0_u3_n657 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U381 (.A1( u0_u3_n702 ) , .ZN( u0_u3_n771 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U382 (.ZN( u0_u3_n668 ) , .A1( u0_u3_n783 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U383 (.ZN( u0_u3_n634 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U384 (.ZN( u0_u3_n475 ) , .A2( w3_26 ) , .A1( w3_27 ) );
  NOR2_X1 u0_u3_U385 (.ZN( u0_u3_n458 ) , .A1( u0_u3_n831 ) , .A2( w3_27 ) );
  INV_X1 u0_u3_U386 (.ZN( u0_u3_n832 ) , .A( w3_27 ) );
  NOR3_X1 u0_u3_U387 (.A3( u0_u3_n624 ) , .A2( u0_u3_n625 ) , .ZN( u0_u3_n639 ) , .A1( u0_u3_n728 ) );
  NOR4_X1 u0_u3_U388 (.A1( u0_u3_n587 ) , .ZN( u0_u3_n588 ) , .A3( u0_u3_n655 ) , .A2( u0_u3_n665 ) , .A4( u0_u3_n770 ) );
  OAI22_X1 u0_u3_U389 (.ZN( u0_u3_n640 ) , .A1( u0_u3_n702 ) , .B2( u0_u3_n731 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n819 ) );
  NOR3_X1 u0_u3_U39 (.A3( u0_u3_n657 ) , .A2( u0_u3_n658 ) , .A1( u0_u3_n659 ) , .ZN( u0_u3_n660 ) );
  AOI21_X1 u0_u3_U390 (.ZN( u0_u3_n502 ) , .B1( u0_u3_n683 ) , .A( u0_u3_n815 ) , .B2( u0_u3_n819 ) );
  OAI22_X1 u0_u3_U391 (.A1( u0_u3_n727 ) , .ZN( u0_u3_n729 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n815 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U392 (.A( u0_u3_n438 ) , .B2( u0_u3_n819 ) , .B1( u0_u3_n820 ) , .ZN( u0_u3_n821 ) );
  OAI22_X1 u0_u3_U393 (.A1( u0_u3_n438 ) , .ZN( u0_u3_n627 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n750 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U394 (.ZN( u0_u3_n522 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U395 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n691 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U396 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n602 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U397 (.ZN( u0_u3_n534 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U398 (.ZN( u0_u3_n561 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U399 (.ZN( u0_u3_n688 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U4 (.A1( u0_u3_n452 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U40 (.A4( u0_u3_n664 ) , .A3( u0_u3_n665 ) , .A2( u0_u3_n666 ) , .A1( u0_u3_n667 ) , .ZN( u0_u3_n680 ) );
  INV_X1 u0_u3_U400 (.A( u0_u3_n819 ) , .ZN( u0_u3_n834 ) );
  NAND2_X1 u0_u3_U401 (.ZN( u0_u3_n674 ) , .A1( u0_u3_n809 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U402 (.ZN( u0_u3_n465 ) , .A2( w3_24 ) , .A1( w3_25 ) );
  NOR2_X1 u0_u3_U403 (.ZN( u0_u3_n457 ) , .A1( u0_u3_n830 ) , .A2( w3_24 ) );
  INV_X1 u0_u3_U404 (.ZN( u0_u3_n829 ) , .A( w3_24 ) );
  INV_X1 u0_u3_U405 (.ZN( u0_u3_n850 ) , .A( w3_29 ) );
  NOR2_X1 u0_u3_U406 (.ZN( u0_u3_n451 ) , .A1( u0_u3_n849 ) , .A2( w3_29 ) );
  NAND4_X1 u0_u3_U407 (.ZN( u0_subword_3 ) , .A4( u0_u3_n707 ) , .A3( u0_u3_n708 ) , .A2( u0_u3_n709 ) , .A1( u0_u3_n710 ) );
  INV_X1 u0_u3_U408 (.A( u0_u3_n709 ) , .ZN( u0_u3_n878 ) );
  OAI22_X1 u0_u3_U409 (.B2( u0_u3_n747 ) , .ZN( u0_u3_n749 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n783 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U41 (.A4( u0_u3_n668 ) , .A3( u0_u3_n669 ) , .A2( u0_u3_n670 ) , .A1( u0_u3_n671 ) , .ZN( u0_u3_n679 ) );
  OAI22_X1 u0_u3_U410 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n499 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n809 ) );
  NOR2_X1 u0_u3_U411 (.ZN( u0_u3_n519 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n747 ) );
  OAI22_X1 u0_u3_U412 (.ZN( u0_u3_n713 ) , .A2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .A1( u0_u3_n747 ) , .B1( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U413 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n772 ) , .A1( u0_u3_n815 ) );
  OAI22_X1 u0_u3_U414 (.B1( u0_u3_n443 ) , .ZN( u0_u3_n447 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n747 ) , .B2( u0_u3_n752 ) );
  NOR2_X1 u0_u3_U415 (.ZN( u0_u3_n550 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U416 (.ZN( u0_u3_n556 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U417 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n758 ) , .A1( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U418 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n676 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U419 (.ZN( u0_u3_n533 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U42 (.A3( u0_u3_n676 ) , .A1( u0_u3_n677 ) , .ZN( u0_u3_n678 ) , .A4( u0_u3_n718 ) , .A2( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U420 (.ZN( u0_u3_n721 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U421 (.ZN( u0_u3_n585 ) , .A1( u0_u3_n747 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U422 (.A( u0_u3_n747 ) , .ZN( u0_u3_n839 ) );
  AOI21_X1 u0_u3_U423 (.ZN( u0_u3_n579 ) , .B2( u0_u3_n727 ) , .B1( u0_u3_n751 ) , .A( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U424 (.A4( u0_u3_n636 ) , .A3( u0_u3_n637 ) , .A2( u0_u3_n638 ) , .A1( u0_u3_n639 ) , .ZN( u0_u3_n746 ) );
  INV_X1 u0_u3_U425 (.ZN( u0_u3_n851 ) , .A( w3_30 ) );
  INV_X1 u0_u3_U426 (.ZN( u0_u3_n860 ) , .A( w3_31 ) );
  NAND4_X1 u0_u3_U427 (.ZN( u0_subword_2 ) , .A4( u0_u3_n646 ) , .A3( u0_u3_n647 ) , .A2( u0_u3_n648 ) , .A1( u0_u3_n649 ) );
  AOI211_X1 u0_u3_U428 (.A( u0_u3_n640 ) , .ZN( u0_u3_n648 ) , .B( u0_u3_n746 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n856 ) );
  NOR2_X1 u0_u3_U429 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n603 ) , .A1( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U43 (.A1( u0_u3_n469 ) , .ZN( u0_u3_n470 ) , .A4( u0_u3_n545 ) , .A2( u0_u3_n557 ) , .A3( u0_u3_n617 ) );
  OAI222_X1 u0_u3_U430 (.A2( u0_u3_n672 ) , .ZN( u0_u3_n677 ) , .B1( u0_u3_n750 ) , .B2( u0_u3_n787 ) , .C2( u0_u3_n791 ) , .C1( u0_u3_n818 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U431 (.ZN( u0_u3_n613 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U432 (.A( u0_u3_n41 ) , .ZN( u0_u3_n503 ) , .B1( u0_u3_n711 ) , .B2( u0_u3_n789 ) );
  OAI22_X1 u0_u3_U433 (.ZN( u0_u3_n593 ) , .B1( u0_u3_n733 ) , .B2( u0_u3_n752 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U434 (.ZN( u0_u3_n656 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U435 (.A2( u0_u3_n752 ) , .A1( u0_u3_n789 ) , .ZN( u0_u3_n812 ) );
  NOR2_X1 u0_u3_U436 (.ZN( u0_u3_n557 ) , .A1( u0_u3_n789 ) , .A2( u0_u3_n816 ) );
  NAND3_X1 u0_u3_U437 (.ZN( u0_subword_6 ) , .A3( u0_u3_n800 ) , .A2( u0_u3_n801 ) , .A1( u0_u3_n802 ) );
  NAND3_X1 u0_u3_U438 (.ZN( u0_subword_5 ) , .A3( u0_u3_n761 ) , .A2( u0_u3_n762 ) , .A1( u0_u3_n763 ) );
  NAND3_X1 u0_u3_U439 (.ZN( u0_subword_4 ) , .A3( u0_u3_n741 ) , .A2( u0_u3_n742 ) , .A1( u0_u3_n743 ) );
  AOI221_X1 u0_u3_U44 (.ZN( u0_u3_n471 ) , .C2( u0_u3_n717 ) , .B2( u0_u3_n834 ) , .C1( u0_u3_n847 ) , .B1( u0_u3_n862 ) , .A( u0_u3_n866 ) );
  NAND3_X1 u0_u3_U440 (.A3( u0_u3_n678 ) , .A2( u0_u3_n679 ) , .A1( u0_u3_n680 ) , .ZN( u0_u3_n810 ) );
  NAND3_X1 u0_u3_U441 (.ZN( u0_u3_n641 ) , .A3( u0_u3_n711 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n795 ) );
  NAND3_X1 u0_u3_U442 (.A3( u0_u3_n621 ) , .A2( u0_u3_n622 ) , .A1( u0_u3_n623 ) , .ZN( u0_u3_n728 ) );
  NAND3_X1 u0_u3_U443 (.A3( u0_u3_n588 ) , .A2( u0_u3_n589 ) , .A1( u0_u3_n590 ) , .ZN( u0_u3_n624 ) );
  NAND3_X1 u0_u3_U444 (.ZN( u0_u3_n568 ) , .A3( u0_u3_n683 ) , .A2( u0_u3_n753 ) , .A1( u0_u3_n788 ) );
  NAND3_X1 u0_u3_U445 (.A3( u0_u3_n526 ) , .A2( u0_u3_n527 ) , .A1( u0_u3_n528 ) , .ZN( u0_u3_n745 ) );
  NAND3_X1 u0_u3_U446 (.A3( u0_u3_n515 ) , .A1( u0_u3_n516 ) , .ZN( u0_u3_n611 ) , .A2( u0_u3_n873 ) );
  NAND3_X1 u0_u3_U447 (.A3( u0_u3_n470 ) , .A2( u0_u3_n471 ) , .A1( u0_u3_n472 ) , .ZN( u0_u3_n780 ) );
  NOR2_X1 u0_u3_U448 (.ZN( u0_u3_n615 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n789 ) );
  NOR2_X1 u0_u3_U449 (.ZN( u0_u3_n720 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n789 ) );
  NOR4_X1 u0_u3_U45 (.A4( u0_u3_n517 ) , .A3( u0_u3_n518 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n520 ) , .ZN( u0_u3_n527 ) );
  NOR2_X1 u0_u3_U450 (.ZN( u0_u3_n704 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U451 (.A1( u0_u3_n733 ) , .ZN( u0_u3_n768 ) , .A2( u0_u3_n789 ) );
  INV_X1 u0_u3_U452 (.ZN( u0_u3_n849 ) , .A( w3_28 ) );
  NOR4_X1 u0_u3_U46 (.A3( u0_u3_n524 ) , .A1( u0_u3_n525 ) , .ZN( u0_u3_n526 ) , .A2( u0_u3_n676 ) , .A4( u0_u3_n772 ) );
  NAND4_X1 u0_u3_U47 (.A4( u0_u3_n576 ) , .A3( u0_u3_n577 ) , .A1( u0_u3_n578 ) , .ZN( u0_u3_n726 ) , .A2( u0_u3_n876 ) );
  NOR4_X1 u0_u3_U48 (.A4( u0_u3_n572 ) , .A3( u0_u3_n573 ) , .A2( u0_u3_n574 ) , .A1( u0_u3_n575 ) , .ZN( u0_u3_n576 ) );
  INV_X1 u0_u3_U49 (.A( u0_u3_n610 ) , .ZN( u0_u3_n876 ) );
  NAND2_X1 u0_u3_U5 (.A1( u0_u3_n456 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U50 (.A4( u0_u3_n459 ) , .A3( u0_u3_n460 ) , .A2( u0_u3_n461 ) , .A1( u0_u3_n462 ) , .ZN( u0_u3_n682 ) );
  NOR3_X1 u0_u3_U51 (.ZN( u0_u3_n460 ) , .A3( u0_u3_n533 ) , .A1( u0_u3_n558 ) , .A2( u0_u3_n573 ) );
  NOR4_X1 u0_u3_U52 (.ZN( u0_u3_n459 ) , .A2( u0_u3_n520 ) , .A1( u0_u3_n546 ) , .A3( u0_u3_n582 ) , .A4( u0_u3_n618 ) );
  NOR4_X1 u0_u3_U53 (.ZN( u0_u3_n461 ) , .A2( u0_u3_n512 ) , .A1( u0_u3_n602 ) , .A4( u0_u3_n631 ) , .A3( u0_u3_n714 ) );
  NAND4_X1 u0_u3_U54 (.A4( u0_u3_n722 ) , .A3( u0_u3_n723 ) , .A2( u0_u3_n724 ) , .ZN( u0_u3_n744 ) , .A1( u0_u3_n859 ) );
  INV_X1 u0_u3_U55 (.A( u0_u3_n712 ) , .ZN( u0_u3_n859 ) );
  NOR4_X1 u0_u3_U56 (.A4( u0_u3_n718 ) , .A3( u0_u3_n719 ) , .A2( u0_u3_n720 ) , .A1( u0_u3_n721 ) , .ZN( u0_u3_n722 ) );
  NOR3_X1 u0_u3_U57 (.ZN( u0_u3_n483 ) , .A2( u0_u3_n511 ) , .A3( u0_u3_n604 ) , .A1( u0_u3_n613 ) );
  NOR4_X1 u0_u3_U58 (.ZN( u0_u3_n484 ) , .A3( u0_u3_n535 ) , .A4( u0_u3_n548 ) , .A2( u0_u3_n570 ) , .A1( u0_u3_n720 ) );
  AOI211_X1 u0_u3_U59 (.B( u0_u3_n480 ) , .A( u0_u3_n481 ) , .ZN( u0_u3_n485 ) , .C2( u0_u3_n836 ) , .C1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U6 (.ZN( u0_u3_n601 ) , .A1( u0_u3_n611 ) , .A3( u0_u3_n726 ) , .A2( u0_u3_n745 ) );
  INV_X1 u0_u3_U60 (.A( u0_u3_n682 ) , .ZN( u0_u3_n874 ) );
  NOR4_X1 u0_u3_U61 (.A4( u0_u3_n690 ) , .A3( u0_u3_n691 ) , .A2( u0_u3_n692 ) , .A1( u0_u3_n693 ) , .ZN( u0_u3_n694 ) );
  AOI221_X1 u0_u3_U62 (.A( u0_u3_n684 ) , .ZN( u0_u3_n695 ) , .B2( u0_u3_n842 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n867 ) );
  NAND4_X1 u0_u3_U63 (.A4( u0_u3_n476 ) , .A3( u0_u3_n477 ) , .A2( u0_u3_n478 ) , .A1( u0_u3_n479 ) , .ZN( u0_u3_n681 ) );
  NOR4_X1 u0_u3_U64 (.A4( u0_u3_n473 ) , .ZN( u0_u3_n479 ) , .A3( u0_u3_n559 ) , .A1( u0_u3_n738 ) , .A2( u0_u3_n758 ) );
  NOR4_X1 u0_u3_U65 (.ZN( u0_u3_n477 ) , .A1( u0_u3_n509 ) , .A3( u0_u3_n547 ) , .A2( u0_u3_n586 ) , .A4( u0_u3_n719 ) );
  NOR4_X1 u0_u3_U66 (.ZN( u0_u3_n476 ) , .A2( u0_u3_n524 ) , .A4( u0_u3_n597 ) , .A1( u0_u3_n612 ) , .A3( u0_u3_n632 ) );
  NAND4_X1 u0_u3_U67 (.A4( u0_u3_n551 ) , .A3( u0_u3_n552 ) , .A2( u0_u3_n553 ) , .A1( u0_u3_n554 ) , .ZN( u0_u3_n748 ) );
  AOI211_X1 u0_u3_U68 (.B( u0_u3_n542 ) , .A( u0_u3_n543 ) , .ZN( u0_u3_n554 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  NOR3_X1 u0_u3_U69 (.ZN( u0_u3_n552 ) , .A2( u0_u3_n654 ) , .A1( u0_u3_n670 ) , .A3( u0_u3_n774 ) );
  NOR3_X1 u0_u3_U7 (.ZN( u0_u3_n507 ) , .A2( u0_u3_n682 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n878 ) );
  NOR4_X1 u0_u3_U70 (.A4( u0_u3_n544 ) , .A3( u0_u3_n545 ) , .A2( u0_u3_n546 ) , .ZN( u0_u3_n553 ) , .A1( u0_u3_n691 ) );
  NOR4_X1 u0_u3_U71 (.A4( u0_u3_n612 ) , .A3( u0_u3_n613 ) , .A2( u0_u3_n614 ) , .A1( u0_u3_n615 ) , .ZN( u0_u3_n622 ) );
  NOR4_X1 u0_u3_U72 (.ZN( u0_u3_n623 ) , .A1( u0_u3_n659 ) , .A3( u0_u3_n669 ) , .A4( u0_u3_n685 ) , .A2( u0_u3_n769 ) );
  INV_X1 u0_u3_U73 (.A( u0_u3_n765 ) , .ZN( u0_u3_n833 ) );
  NOR2_X1 u0_u3_U74 (.ZN( u0_u3_n650 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n870 ) );
  NOR4_X1 u0_u3_U75 (.A4( u0_u3_n580 ) , .A3( u0_u3_n581 ) , .A2( u0_u3_n582 ) , .ZN( u0_u3_n589 ) , .A1( u0_u3_n686 ) );
  INV_X1 u0_u3_U76 (.A( u0_u3_n818 ) , .ZN( u0_u3_n857 ) );
  OR4_X1 u0_u3_U77 (.A4( u0_u3_n685 ) , .A3( u0_u3_n686 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n688 ) , .ZN( u0_u3_n693 ) );
  OR4_X1 u0_u3_U78 (.ZN( u0_u3_n469 ) , .A4( u0_u3_n521 ) , .A3( u0_u3_n532 ) , .A2( u0_u3_n581 ) , .A1( u0_u3_n715 ) );
  OR4_X1 u0_u3_U79 (.A4( u0_u3_n569 ) , .A3( u0_u3_n570 ) , .A2( u0_u3_n571 ) , .ZN( u0_u3_n575 ) , .A1( u0_u3_n668 ) );
  NOR3_X1 u0_u3_U8 (.A2( u0_u3_n610 ) , .A1( u0_u3_n611 ) , .ZN( u0_u3_n649 ) , .A3( u0_u3_n725 ) );
  OR4_X1 u0_u3_U80 (.A4( u0_u3_n521 ) , .A2( u0_u3_n522 ) , .A1( u0_u3_n523 ) , .ZN( u0_u3_n525 ) , .A3( u0_u3_n824 ) );
  OR4_X1 u0_u3_U81 (.A4( u0_u3_n583 ) , .A3( u0_u3_n584 ) , .A2( u0_u3_n585 ) , .A1( u0_u3_n586 ) , .ZN( u0_u3_n587 ) );
  OR4_X1 u0_u3_U82 (.ZN( u0_u3_n495 ) , .A4( u0_u3_n537 ) , .A2( u0_u3_n550 ) , .A1( u0_u3_n562 ) , .A3( u0_u3_n635 ) );
  NOR4_X1 u0_u3_U83 (.A4( u0_u3_n512 ) , .A2( u0_u3_n513 ) , .A1( u0_u3_n514 ) , .ZN( u0_u3_n515 ) , .A3( u0_u3_n673 ) );
  INV_X1 u0_u3_U84 (.A( u0_u3_n508 ) , .ZN( u0_u3_n873 ) );
  OR3_X1 u0_u3_U85 (.A3( u0_u3_n509 ) , .A2( u0_u3_n510 ) , .A1( u0_u3_n511 ) , .ZN( u0_u3_n514 ) );
  INV_X1 u0_u3_U86 (.A( u0_u3_n757 ) , .ZN( u0_u3_n871 ) );
  AOI221_X1 u0_u3_U87 (.A( u0_u3_n716 ) , .B2( u0_u3_n717 ) , .ZN( u0_u3_n723 ) , .C1( u0_u3_n835 ) , .B1( u0_u3_n841 ) , .C2( u0_u3_n865 ) );
  OR2_X1 u0_u3_U88 (.A2( u0_u3_n714 ) , .A1( u0_u3_n715 ) , .ZN( u0_u3_n716 ) );
  INV_X1 u0_u3_U89 (.A( u0_u3_n466 ) , .ZN( u0_u3_n866 ) );
  NOR3_X1 u0_u3_U9 (.A3( u0_u3_n725 ) , .A1( u0_u3_n726 ) , .ZN( u0_u3_n743 ) , .A2( u0_u3_n744 ) );
  NAND2_X1 u0_u3_U90 (.A1( u0_u3_n454 ) , .A2( u0_u3_n456 ) , .ZN( u0_u3_n765 ) );
  AOI22_X1 u0_u3_U91 (.ZN( u0_u3_n699 ) , .A1( u0_u3_n833 ) , .B2( u0_u3_n845 ) , .A2( u0_u3_n867 ) , .B1( u0_u3_n870 ) );
  NOR3_X1 u0_u3_U92 (.ZN( u0_u3_n755 ) , .A2( u0_u3_n855 ) , .A1( u0_u3_n865 ) , .A3( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U93 (.ZN( u0_u3_n754 ) , .A2( u0_u3_n854 ) , .A1( u0_u3_n862 ) );
  AOI211_X1 u0_u3_U94 (.A( u0_u3_n499 ) , .ZN( u0_u3_n506 ) , .B( u0_u3_n805 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  AOI211_X1 u0_u3_U95 (.B( u0_u3_n810 ) , .A( u0_u3_n811 ) , .ZN( u0_u3_n827 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n852 ) );
  NAND2_X1 u0_u3_U96 (.A1( u0_u3_n450 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n752 ) );
  INV_X1 u0_u3_U97 (.A( u0_u3_n733 ) , .ZN( u0_u3_n841 ) );
  AOI221_X1 u0_u3_U98 (.B2( u0_u3_n440 ) , .A( u0_u3_n492 ) , .ZN( u0_u3_n497 ) , .C2( u0_u3_n843 ) , .C1( u0_u3_n853 ) , .B1( u0_u3_n862 ) );
  INV_X1 u0_u3_U99 (.A( u0_u3_n781 ) , .ZN( u0_u3_n869 ) );
  NOR2_X1 us10_U10 (.A1( us10_n678 ) , .ZN( us10_n693 ) , .A2( us10_n807 ) );
  NOR3_X1 us10_U100 (.ZN( us10_n549 ) , .A2( us10_n651 ) , .A1( us10_n667 ) , .A3( us10_n771 ) );
  AOI211_X1 us10_U101 (.B( us10_n539 ) , .A( us10_n540 ) , .ZN( us10_n551 ) , .C2( us10_n839 ) , .C1( us10_n851 ) );
  NOR4_X1 us10_U102 (.A4( us10_n544 ) , .A3( us10_n545 ) , .A2( us10_n546 ) , .A1( us10_n547 ) , .ZN( us10_n548 ) );
  NOR4_X1 us10_U103 (.ZN( us10_n620 ) , .A1( us10_n656 ) , .A3( us10_n666 ) , .A4( us10_n682 ) , .A2( us10_n766 ) );
  NOR4_X1 us10_U104 (.A4( us10_n609 ) , .A3( us10_n610 ) , .A2( us10_n611 ) , .A1( us10_n612 ) , .ZN( us10_n619 ) );
  NOR4_X1 us10_U105 (.A4( us10_n614 ) , .A3( us10_n615 ) , .A2( us10_n616 ) , .A1( us10_n617 ) , .ZN( us10_n618 ) );
  NAND4_X1 us10_U106 (.A4( us10_n485 ) , .A3( us10_n486 ) , .A2( us10_n487 ) , .A1( us10_n488 ) , .ZN( us10_n778 ) );
  NOR4_X1 us10_U107 (.A4( us10_n484 ) , .ZN( us10_n487 ) , .A1( us10_n566 ) , .A2( us10_n581 ) , .A3( us10_n602 ) );
  NOR4_X1 us10_U108 (.ZN( us10_n486 ) , .A1( us10_n507 ) , .A2( us10_n519 ) , .A4( us10_n546 ) , .A3( us10_n611 ) );
  NOR4_X1 us10_U109 (.ZN( us10_n485 ) , .A2( us10_n533 ) , .A1( us10_n558 ) , .A3( us10_n631 ) , .A4( us10_n718 ) );
  INV_X1 us10_U11 (.A( us10_n680 ) , .ZN( us10_n840 ) );
  NAND4_X1 us10_U110 (.A4( us10_n691 ) , .A3( us10_n692 ) , .A1( us10_n693 ) , .ZN( us10_n776 ) , .A2( us10_n872 ) );
  AOI221_X1 us10_U111 (.A( us10_n681 ) , .ZN( us10_n692 ) , .B2( us10_n840 ) , .C1( us10_n842 ) , .C2( us10_n862 ) , .B1( us10_n865 ) );
  INV_X1 us10_U112 (.A( us10_n679 ) , .ZN( us10_n872 ) );
  NOR4_X1 us10_U113 (.A4( us10_n687 ) , .A3( us10_n688 ) , .A2( us10_n689 ) , .A1( us10_n690 ) , .ZN( us10_n691 ) );
  NAND4_X1 us10_U114 (.A4( us10_n473 ) , .A3( us10_n474 ) , .A2( us10_n475 ) , .A1( us10_n476 ) , .ZN( us10_n678 ) );
  NOR4_X1 us10_U115 (.A4( us10_n470 ) , .ZN( us10_n476 ) , .A3( us10_n556 ) , .A1( us10_n735 ) , .A2( us10_n755 ) );
  NOR4_X1 us10_U116 (.ZN( us10_n475 ) , .A1( us10_n531 ) , .A3( us10_n568 ) , .A4( us10_n600 ) , .A2( us10_n642 ) );
  NOR4_X1 us10_U117 (.ZN( us10_n474 ) , .A1( us10_n506 ) , .A3( us10_n544 ) , .A2( us10_n583 ) , .A4( us10_n716 ) );
  NAND4_X1 us10_U118 (.A4( us10_n719 ) , .A3( us10_n720 ) , .A2( us10_n721 ) , .ZN( us10_n741 ) , .A1( us10_n857 ) );
  INV_X1 us10_U119 (.A( us10_n709 ) , .ZN( us10_n857 ) );
  NOR4_X1 us10_U12 (.A4( us10_n445 ) , .A3( us10_n446 ) , .A2( us10_n516 ) , .A1( us10_n541 ) , .ZN( us10_n706 ) );
  NOR4_X1 us10_U120 (.A4( us10_n715 ) , .A3( us10_n716 ) , .A2( us10_n717 ) , .A1( us10_n718 ) , .ZN( us10_n719 ) );
  AOI221_X1 us10_U121 (.A( us10_n710 ) , .ZN( us10_n721 ) , .C2( us10_n844 ) , .B2( us10_n845 ) , .C1( us10_n861 ) , .B1( us10_n862 ) );
  NOR2_X1 us10_U122 (.ZN( us10_n789 ) , .A2( us10_n862 ) , .A1( us10_n868 ) );
  NOR2_X1 us10_U123 (.ZN( us10_n733 ) , .A2( us10_n832 ) , .A1( us10_n845 ) );
  NAND4_X1 us10_U124 (.A4( us10_n573 ) , .A3( us10_n574 ) , .A1( us10_n575 ) , .ZN( us10_n723 ) , .A2( us10_n874 ) );
  NOR4_X1 us10_U125 (.A4( us10_n569 ) , .A3( us10_n570 ) , .A2( us10_n571 ) , .A1( us10_n572 ) , .ZN( us10_n573 ) );
  AOI221_X1 us10_U126 (.A( us10_n564 ) , .C2( us10_n565 ) , .ZN( us10_n574 ) , .B2( us10_n845 ) , .B1( us10_n852 ) , .C1( us10_n853 ) );
  INV_X1 us10_U127 (.A( us10_n607 ) , .ZN( us10_n874 ) );
  NAND4_X1 us10_U128 (.A4( us10_n633 ) , .A3( us10_n634 ) , .A2( us10_n635 ) , .A1( us10_n636 ) , .ZN( us10_n743 ) );
  AOI211_X1 us10_U129 (.B( us10_n623 ) , .A( us10_n624 ) , .ZN( us10_n635 ) , .C2( us10_n836 ) , .C1( us10_n863 ) );
  OR3_X1 us10_U13 (.ZN( us10_n446 ) , .A1( us10_n528 ) , .A3( us10_n577 ) , .A2( us10_n875 ) );
  NOR4_X1 us10_U130 (.A4( us10_n629 ) , .A3( us10_n630 ) , .A2( us10_n631 ) , .A1( us10_n632 ) , .ZN( us10_n633 ) );
  NOR4_X1 us10_U131 (.A4( us10_n626 ) , .A3( us10_n627 ) , .A2( us10_n628 ) , .ZN( us10_n634 ) , .A1( us10_n664 ) );
  NAND4_X1 us10_U132 (.A4( us10_n493 ) , .A3( us10_n494 ) , .A1( us10_n495 ) , .ZN( us10_n802 ) , .A2( us10_n867 ) );
  AOI221_X1 us10_U133 (.A( us10_n489 ) , .ZN( us10_n494 ) , .B2( us10_n836 ) , .C2( us10_n841 ) , .C1( us10_n851 ) , .B1( us10_n860 ) );
  INV_X1 us10_U134 (.A( us10_n778 ) , .ZN( us10_n867 ) );
  NOR2_X1 us10_U135 (.ZN( us10_n495 ) , .A1( us10_n678 ) , .A2( us10_n694 ) );
  NOR2_X1 us10_U136 (.ZN( us10_n748 ) , .A1( us10_n861 ) , .A2( us10_n862 ) );
  NOR2_X1 us10_U137 (.ZN( us10_n647 ) , .A1( us10_n854 ) , .A2( us10_n868 ) );
  INV_X1 us10_U138 (.A( us10_n762 ) , .ZN( us10_n830 ) );
  OR4_X1 us10_U139 (.ZN( us10_n466 ) , .A4( us10_n518 ) , .A3( us10_n529 ) , .A2( us10_n578 ) , .A1( us10_n712 ) );
  OR4_X1 us10_U14 (.A4( us10_n442 ) , .A2( us10_n443 ) , .A1( us10_n444 ) , .ZN( us10_n445 ) , .A3( us10_n553 ) );
  OR4_X1 us10_U140 (.A4( us10_n566 ) , .A3( us10_n567 ) , .A2( us10_n568 ) , .ZN( us10_n572 ) , .A1( us10_n665 ) );
  OR4_X1 us10_U141 (.A4( us10_n518 ) , .A2( us10_n519 ) , .A1( us10_n520 ) , .ZN( us10_n522 ) , .A3( us10_n821 ) );
  OR4_X1 us10_U142 (.A4( us10_n682 ) , .A3( us10_n683 ) , .A2( us10_n684 ) , .A1( us10_n685 ) , .ZN( us10_n690 ) );
  OR4_X1 us10_U143 (.A4( us10_n580 ) , .A3( us10_n581 ) , .A2( us10_n582 ) , .A1( us10_n583 ) , .ZN( us10_n584 ) );
  NAND2_X1 us10_U144 (.ZN( us10_n613 ) , .A2( us10_n837 ) , .A1( us10_n873 ) );
  OR3_X1 us10_U145 (.A3( us10_n506 ) , .A2( us10_n507 ) , .A1( us10_n508 ) , .ZN( us10_n511 ) );
  INV_X1 us10_U146 (.A( us10_n672 ) , .ZN( us10_n859 ) );
  AOI21_X1 us10_U147 (.A( us10_n670 ) , .B1( us10_n671 ) , .ZN( us10_n672 ) , .B2( us10_n856 ) );
  INV_X1 us10_U148 (.A( us10_n754 ) , .ZN( us10_n869 ) );
  OAI21_X1 us10_U149 (.B1( us10_n753 ) , .ZN( us10_n754 ) , .A( us10_n845 ) , .B2( us10_n868 ) );
  INV_X1 us10_U15 (.A( us10_n613 ) , .ZN( us10_n875 ) );
  INV_X1 us10_U150 (.A( us10_n463 ) , .ZN( us10_n864 ) );
  OAI21_X1 us10_U151 (.ZN( us10_n463 ) , .B1( us10_n809 ) , .A( us10_n834 ) , .B2( us10_n851 ) );
  AOI222_X1 us10_U152 (.ZN( us10_n660 ) , .A2( us10_n839 ) , .B1( us10_n841 ) , .C2( us10_n845 ) , .A1( us10_n860 ) , .C1( us10_n863 ) , .B2( us10_n870 ) );
  INV_X1 us10_U153 (.A( us10_n647 ) , .ZN( us10_n870 ) );
  NAND2_X1 us10_U154 (.A1( us10_n447 ) , .A2( us10_n465 ) , .ZN( us10_n749 ) );
  OAI222_X1 us10_U155 (.B2( us10_n708 ) , .ZN( us10_n709 ) , .C2( us10_n724 ) , .B1( us10_n747 ) , .A1( us10_n806 ) , .C1( us10_n814 ) , .A2( us10_n815 ) );
  OAI222_X1 us10_U156 (.A2( us10_n669 ) , .ZN( us10_n674 ) , .B1( us10_n747 ) , .B2( us10_n784 ) , .C2( us10_n788 ) , .C1( us10_n815 ) , .A1( us10_n817 ) );
  OAI222_X1 us10_U157 (.ZN( us10_n617 ) , .B1( us10_n697 ) , .C1( us10_n724 ) , .C2( us10_n747 ) , .B2( us10_n786 ) , .A2( us10_n792 ) , .A1( us10_n816 ) );
  NOR4_X1 us10_U158 (.A2( us10_n491 ) , .A1( us10_n492 ) , .ZN( us10_n493 ) , .A3( us10_n580 ) , .A4( us10_n612 ) );
  OR4_X1 us10_U159 (.ZN( us10_n492 ) , .A4( us10_n534 ) , .A2( us10_n547 ) , .A1( us10_n559 ) , .A3( us10_n632 ) );
  INV_X1 us10_U16 (.A( us10_n749 ) , .ZN( us10_n863 ) );
  OAI22_X1 us10_U160 (.B1( us10_n490 ) , .ZN( us10_n491 ) , .A1( us10_n686 ) , .A2( us10_n763 ) , .B2( us10_n817 ) );
  NOR3_X1 us10_U161 (.ZN( us10_n490 ) , .A1( us10_n782 ) , .A2( us10_n850 ) , .A3( us10_n863 ) );
  INV_X1 us10_U162 (.A( us10_n730 ) , .ZN( us10_n839 ) );
  AOI221_X1 us10_U163 (.A( us10_n450 ) , .ZN( us10_n459 ) , .C2( us10_n753 ) , .B1( us10_n832 ) , .C1( us10_n842 ) , .B2( us10_n861 ) );
  AOI21_X1 us10_U164 (.ZN( us10_n450 ) , .B2( us10_n792 ) , .A( us10_n803 ) , .B1( us10_n815 ) );
  AOI221_X1 us10_U165 (.A( us10_n483 ) , .ZN( us10_n488 ) , .B1( us10_n831 ) , .C2( us10_n844 ) , .C1( us10_n852 ) , .B2( us10_n862 ) );
  OAI22_X1 us10_U166 (.ZN( us10_n483 ) , .A1( us10_n708 ) , .B2( us10_n785 ) , .A2( us10_n806 ) , .B1( us10_n812 ) );
  INV_X1 us10_U167 (.A( us10_n790 ) , .ZN( us10_n832 ) );
  NAND2_X1 us10_U168 (.A1( us10_n451 ) , .A2( us10_n453 ) , .ZN( us10_n762 ) );
  INV_X1 us10_U169 (.A( us10_n786 ) , .ZN( us10_n862 ) );
  AOI222_X1 us10_U17 (.ZN( us10_n605 ) , .B2( us10_n671 ) , .B1( us10_n753 ) , .C2( us10_n831 ) , .A1( us10_n833 ) , .A2( us10_n862 ) , .C1( us10_n863 ) );
  OAI221_X1 us10_U170 (.A( us10_n783 ) , .C2( us10_n784 ) , .B2( us10_n785 ) , .B1( us10_n786 ) , .ZN( us10_n796 ) , .C1( us10_n813 ) );
  AOI22_X1 us10_U171 (.A2( us10_n782 ) , .ZN( us10_n783 ) , .B2( us10_n831 ) , .A1( us10_n834 ) , .B1( us10_n863 ) );
  OAI221_X1 us10_U172 (.A( us10_n696 ) , .ZN( us10_n703 ) , .C2( us10_n784 ) , .C1( us10_n785 ) , .B1( us10_n786 ) , .B2( us10_n806 ) );
  AOI22_X1 us10_U173 (.ZN( us10_n696 ) , .A1( us10_n830 ) , .B2( us10_n843 ) , .A2( us10_n865 ) , .B1( us10_n868 ) );
  OAI221_X1 us10_U174 (.A( us10_n727 ) , .C2( us10_n728 ) , .B2( us10_n729 ) , .B1( us10_n730 ) , .ZN( us10_n737 ) , .C1( us10_n817 ) );
  AOI22_X1 us10_U175 (.ZN( us10_n727 ) , .B1( us10_n832 ) , .A2( us10_n838 ) , .A1( us10_n863 ) , .B2( us10_n866 ) );
  INV_X1 us10_U176 (.A( us10_n784 ) , .ZN( us10_n861 ) );
  OAI22_X1 us10_U177 (.ZN( us10_n710 ) , .A2( us10_n728 ) , .B2( us10_n729 ) , .A1( us10_n744 ) , .B1( us10_n813 ) );
  INV_X1 us10_U178 (.A( us10_n816 ) , .ZN( us10_n831 ) );
  INV_X1 us10_U179 (.A( us10_n788 ) , .ZN( us10_n845 ) );
  AOI222_X1 us10_U18 (.ZN( us10_n563 ) , .B1( us10_n830 ) , .C1( us10_n841 ) , .A2( us10_n843 ) , .A1( us10_n854 ) , .B2( us10_n863 ) , .C2( us10_n873 ) );
  OAI22_X1 us10_U180 (.ZN( us10_n588 ) , .A2( us10_n747 ) , .B2( us10_n762 ) , .A1( us10_n763 ) , .B1( us10_n784 ) );
  OAI22_X1 us10_U181 (.ZN( us10_n489 ) , .A1( us10_n724 ) , .B2( us10_n728 ) , .B1( us10_n730 ) , .A2( us10_n779 ) );
  OAI22_X1 us10_U182 (.ZN( us10_n624 ) , .B1( us10_n669 ) , .B2( us10_n747 ) , .A1( us10_n815 ) , .A2( us10_n816 ) );
  INV_X1 us10_U183 (.A( us10_n744 ) , .ZN( us10_n837 ) );
  OAI22_X1 us10_U184 (.ZN( us10_n681 ) , .A1( us10_n699 ) , .A2( us10_n730 ) , .B2( us10_n784 ) , .B1( us10_n817 ) );
  OAI22_X1 us10_U185 (.B2( us10_n779 ) , .B1( us10_n780 ) , .ZN( us10_n781 ) , .A2( us10_n814 ) , .A1( us10_n815 ) );
  OAI22_X1 us10_U186 (.A1( us10_n724 ) , .ZN( us10_n726 ) , .B2( us10_n750 ) , .B1( us10_n812 ) , .A2( us10_n816 ) );
  INV_X1 us10_U187 (.A( us10_n814 ) , .ZN( us10_n833 ) );
  OAI22_X1 us10_U188 (.B2( us10_n744 ) , .ZN( us10_n746 ) , .A2( us10_n762 ) , .B1( us10_n780 ) , .A1( us10_n792 ) );
  INV_X1 us10_U189 (.A( us10_n669 ) , .ZN( us10_n865 ) );
  NOR4_X1 us10_U19 (.ZN( us10_n473 ) , .A2( us10_n521 ) , .A4( us10_n594 ) , .A1( us10_n609 ) , .A3( us10_n629 ) );
  OAI22_X1 us10_U190 (.ZN( us10_n496 ) , .A2( us10_n744 ) , .A1( us10_n780 ) , .B1( us10_n791 ) , .B2( us10_n806 ) );
  INV_X1 us10_U191 (.A( us10_n750 ) , .ZN( us10_n842 ) );
  AOI211_X1 us10_U192 (.A( us10_n637 ) , .ZN( us10_n645 ) , .B( us10_n743 ) , .C2( us10_n839 ) , .C1( us10_n854 ) );
  OAI22_X1 us10_U193 (.ZN( us10_n637 ) , .A1( us10_n699 ) , .B2( us10_n728 ) , .A2( us10_n762 ) , .B1( us10_n816 ) );
  OAI22_X1 us10_U194 (.ZN( us10_n590 ) , .B1( us10_n730 ) , .B2( us10_n749 ) , .A2( us10_n786 ) , .A1( us10_n803 ) );
  OAI22_X1 us10_U195 (.ZN( us10_n695 ) , .A2( us10_n730 ) , .A1( us10_n780 ) , .B1( us10_n791 ) , .B2( us10_n817 ) );
  INV_X1 us10_U196 (.A( us10_n747 ) , .ZN( us10_n834 ) );
  NOR2_X1 us10_U197 (.A1( us10_n697 ) , .ZN( us10_n770 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U198 (.ZN( us10_n666 ) , .A1( us10_n728 ) , .A2( us10_n803 ) );
  NOR2_X1 us10_U199 (.ZN( us10_n594 ) , .A2( us10_n697 ) , .A1( us10_n728 ) );
  NOR4_X1 us10_U20 (.ZN( us10_n479 ) , .A1( us10_n520 ) , .A4( us10_n557 ) , .A3( us10_n582 ) , .A2( us10_n630 ) );
  NOR2_X1 us10_U200 (.ZN( us10_n600 ) , .A2( us10_n697 ) , .A1( us10_n784 ) );
  NOR2_X1 us10_U201 (.ZN( us10_n570 ) , .A1( us10_n728 ) , .A2( us10_n806 ) );
  NOR2_X1 us10_U202 (.ZN( us10_n532 ) , .A2( us10_n749 ) , .A1( us10_n750 ) );
  NOR2_X1 us10_U203 (.ZN( us10_n615 ) , .A1( us10_n785 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U204 (.ZN( us10_n629 ) , .A2( us10_n728 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U205 (.ZN( us10_n654 ) , .A1( us10_n728 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U206 (.ZN( us10_n546 ) , .A2( us10_n780 ) , .A1( us10_n814 ) );
  NOR2_X1 us10_U207 (.ZN( us10_n718 ) , .A2( us10_n724 ) , .A1( us10_n744 ) );
  NOR2_X1 us10_U208 (.ZN( us10_n577 ) , .A2( us10_n699 ) , .A1( us10_n814 ) );
  NOR2_X1 us10_U209 (.ZN( us10_n612 ) , .A1( us10_n779 ) , .A2( us10_n786 ) );
  NOR4_X1 us10_U21 (.A4( us10_n532 ) , .A3( us10_n533 ) , .A2( us10_n534 ) , .ZN( us10_n535 ) , .A1( us10_n820 ) );
  NOR2_X1 us10_U210 (.ZN( us10_n628 ) , .A2( us10_n669 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U211 (.ZN( us10_n610 ) , .A1( us10_n784 ) , .A2( us10_n816 ) );
  NOR2_X1 us10_U212 (.ZN( us10_n651 ) , .A1( us10_n784 ) , .A2( us10_n788 ) );
  NOR2_X1 us10_U213 (.ZN( us10_n531 ) , .A2( us10_n780 ) , .A1( us10_n816 ) );
  NOR2_X1 us10_U214 (.ZN( us10_n599 ) , .A2( us10_n791 ) , .A1( us10_n816 ) );
  INV_X1 us10_U215 (.A( us10_n728 ) , .ZN( us10_n852 ) );
  NOR2_X1 us10_U216 (.A2( us10_n708 ) , .A1( us10_n750 ) , .ZN( us10_n771 ) );
  NOR2_X1 us10_U217 (.A1( us10_n699 ) , .ZN( us10_n768 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U218 (.ZN( us10_n667 ) , .A1( us10_n750 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U219 (.ZN( us10_n541 ) , .A2( us10_n697 ) , .A1( us10_n699 ) );
  NOR4_X1 us10_U22 (.A4( us10_n541 ) , .A3( us10_n542 ) , .A2( us10_n543 ) , .ZN( us10_n550 ) , .A1( us10_n688 ) );
  NOR2_X1 us10_U220 (.ZN( us10_n508 ) , .A2( us10_n780 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U221 (.ZN( us10_n543 ) , .A2( us10_n708 ) , .A1( us10_n785 ) );
  NOR2_X1 us10_U222 (.ZN( us10_n555 ) , .A1( us10_n750 ) , .A2( us10_n791 ) );
  NOR2_X1 us10_U223 (.ZN( us10_n611 ) , .A2( us10_n780 ) , .A1( us10_n806 ) );
  NOR2_X1 us10_U224 (.ZN( us10_n664 ) , .A1( us10_n785 ) , .A2( us10_n791 ) );
  NOR2_X1 us10_U225 (.ZN( us10_n652 ) , .A1( us10_n669 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U226 (.A1( us10_n669 ) , .ZN( us10_n673 ) , .A2( us10_n744 ) );
  NOR2_X1 us10_U227 (.ZN( us10_n602 ) , .A1( us10_n669 ) , .A2( us10_n803 ) );
  NOR2_X1 us10_U228 (.A1( us10_n669 ) , .ZN( us10_n688 ) , .A2( us10_n816 ) );
  NOR2_X1 us10_U229 (.A2( us10_n744 ) , .ZN( us10_n769 ) , .A1( us10_n812 ) );
  AOI221_X1 us10_U23 (.A( us10_n713 ) , .B2( us10_n714 ) , .ZN( us10_n720 ) , .C1( us10_n832 ) , .B1( us10_n839 ) , .C2( us10_n863 ) );
  INV_X1 us10_U230 (.A( us10_n792 ) , .ZN( us10_n851 ) );
  NOR2_X1 us10_U231 (.A1( us10_n669 ) , .ZN( us10_n766 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U232 (.ZN( us10_n527 ) , .A1( us10_n669 ) , .A2( us10_n779 ) );
  NOR2_X1 us10_U233 (.A2( us10_n697 ) , .ZN( us10_n716 ) , .A1( us10_n792 ) );
  OAI22_X1 us10_U234 (.B1( us10_n440 ) , .ZN( us10_n444 ) , .A2( us10_n728 ) , .A1( us10_n744 ) , .B2( us10_n749 ) );
  NOR3_X1 us10_U235 (.ZN( us10_n440 ) , .A2( us10_n836 ) , .A3( us10_n837 ) , .A1( us10_n846 ) );
  NOR2_X1 us10_U236 (.ZN( us10_n601 ) , .A2( us10_n780 ) , .A1( us10_n803 ) );
  NOR2_X1 us10_U237 (.ZN( us10_n661 ) , .A1( us10_n729 ) , .A2( us10_n790 ) );
  NOR2_X1 us10_U238 (.ZN( us10_n631 ) , .A1( us10_n724 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U239 (.ZN( us10_n528 ) , .A2( us10_n724 ) , .A1( us10_n803 ) );
  OR2_X1 us10_U24 (.A2( us10_n711 ) , .A1( us10_n712 ) , .ZN( us10_n713 ) );
  NOR2_X1 us10_U240 (.ZN( us10_n509 ) , .A1( us10_n729 ) , .A2( us10_n779 ) );
  NOR2_X1 us10_U241 (.ZN( us10_n507 ) , .A1( us10_n812 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U242 (.ZN( us10_n662 ) , .A2( us10_n697 ) , .A1( us10_n729 ) );
  NOR2_X1 us10_U243 (.ZN( us10_n630 ) , .A1( us10_n747 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U244 (.ZN( us10_n554 ) , .A1( us10_n786 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U245 (.ZN( us10_n545 ) , .A1( us10_n749 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U246 (.ZN( us10_n557 ) , .A1( us10_n792 ) , .A2( us10_n814 ) );
  NOR2_X1 us10_U247 (.ZN( us10_n717 ) , .A2( us10_n744 ) , .A1( us10_n786 ) );
  NOR2_X1 us10_U248 (.ZN( us10_n544 ) , .A2( us10_n785 ) , .A1( us10_n792 ) );
  INV_X1 us10_U249 (.A( us10_n806 ) , .ZN( us10_n841 ) );
  NOR2_X1 us10_U25 (.ZN( us10_n680 ) , .A2( us10_n834 ) , .A1( us10_n839 ) );
  OAI21_X1 us10_U250 (.ZN( us10_n731 ) , .A( us10_n833 ) , .B2( us10_n852 ) , .B1( us10_n873 ) );
  NOR2_X1 us10_U251 (.A2( us10_n697 ) , .A1( us10_n780 ) , .ZN( us10_n820 ) );
  NOR2_X1 us10_U252 (.ZN( us10_n663 ) , .A1( us10_n729 ) , .A2( us10_n785 ) );
  OAI22_X1 us10_U253 (.B2( us10_n750 ) , .B1( us10_n751 ) , .A1( us10_n752 ) , .ZN( us10_n756 ) , .A2( us10_n806 ) );
  NOR2_X1 us10_U254 (.ZN( us10_n751 ) , .A2( us10_n852 ) , .A1( us10_n860 ) );
  NOR3_X1 us10_U255 (.ZN( us10_n752 ) , .A2( us10_n853 ) , .A1( us10_n863 ) , .A3( us10_n865 ) );
  NOR2_X1 us10_U256 (.ZN( us10_n656 ) , .A1( us10_n747 ) , .A2( us10_n780 ) );
  NOR2_X1 us10_U257 (.ZN( us10_n530 ) , .A2( us10_n744 ) , .A1( us10_n792 ) );
  NOR2_X1 us10_U258 (.ZN( us10_n506 ) , .A2( us10_n728 ) , .A1( us10_n762 ) );
  NOR2_X1 us10_U259 (.ZN( us10_n558 ) , .A1( us10_n708 ) , .A2( us10_n816 ) );
  NOR4_X1 us10_U26 (.A4( us10_n514 ) , .A3( us10_n515 ) , .A2( us10_n516 ) , .A1( us10_n517 ) , .ZN( us10_n524 ) );
  NOR2_X1 us10_U260 (.ZN( us10_n516 ) , .A1( us10_n708 ) , .A2( us10_n744 ) );
  NOR2_X1 us10_U261 (.ZN( us10_n614 ) , .A1( us10_n762 ) , .A2( us10_n812 ) );
  AOI21_X1 us10_U262 (.A( us10_n812 ) , .B2( us10_n813 ) , .B1( us10_n814 ) , .ZN( us10_n819 ) );
  NOR2_X1 us10_U263 (.A1( us10_n749 ) , .ZN( us10_n767 ) , .A2( us10_n803 ) );
  AOI21_X1 us10_U264 (.ZN( us10_n593 ) , .B1( us10_n750 ) , .A( us10_n792 ) , .B2( us10_n813 ) );
  NOR2_X1 us10_U265 (.A1( us10_n730 ) , .ZN( us10_n765 ) , .A2( us10_n786 ) );
  NOR2_X1 us10_U266 (.ZN( us10_n655 ) , .A1( us10_n790 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U267 (.ZN( us10_n701 ) , .A2( us10_n786 ) , .A1( us10_n817 ) );
  NOR2_X1 us10_U268 (.ZN( us10_n579 ) , .A2( us10_n708 ) , .A1( us10_n730 ) );
  NOR2_X1 us10_U269 (.ZN( us10_n533 ) , .A2( us10_n724 ) , .A1( us10_n730 ) );
  AOI222_X1 us10_U27 (.ZN( us10_n525 ) , .A1( us10_n834 ) , .B2( us10_n837 ) , .C1( us10_n844 ) , .C2( us10_n850 ) , .A2( us10_n852 ) , .B1( us10_n866 ) );
  NOR2_X1 us10_U270 (.ZN( us10_n668 ) , .A2( us10_n708 ) , .A1( us10_n790 ) );
  INV_X1 us10_U271 (.A( us10_n813 ) , .ZN( us10_n836 ) );
  NOR2_X1 us10_U272 (.ZN( us10_n521 ) , .A1( us10_n790 ) , .A2( us10_n812 ) );
  AOI21_X1 us10_U273 (.ZN( us10_n571 ) , .B2( us10_n697 ) , .B1( us10_n806 ) , .A( us10_n812 ) );
  INV_X1 us10_U274 (.A( us10_n763 ) , .ZN( us10_n866 ) );
  NOR2_X1 us10_U275 (.ZN( us10_n517 ) , .A1( us10_n708 ) , .A2( us10_n803 ) );
  AOI21_X1 us10_U276 (.A( us10_n815 ) , .B2( us10_n816 ) , .B1( us10_n817 ) , .ZN( us10_n818 ) );
  INV_X1 us10_U277 (.A( us10_n729 ) , .ZN( us10_n868 ) );
  NOR2_X1 us10_U278 (.ZN( us10_n542 ) , .A1( us10_n762 ) , .A2( us10_n791 ) );
  AOI21_X1 us10_U279 (.ZN( us10_n499 ) , .B1( us10_n680 ) , .A( us10_n812 ) , .B2( us10_n816 ) );
  NOR4_X1 us10_U28 (.A3( us10_n521 ) , .A1( us10_n522 ) , .ZN( us10_n523 ) , .A2( us10_n673 ) , .A4( us10_n769 ) );
  NOR2_X1 us10_U280 (.ZN( us10_n609 ) , .A2( us10_n724 ) , .A1( us10_n817 ) );
  NOR2_X1 us10_U281 (.ZN( us10_n642 ) , .A2( us10_n788 ) , .A1( us10_n791 ) );
  AOI21_X1 us10_U282 (.ZN( us10_n592 ) , .B1( us10_n728 ) , .B2( us10_n784 ) , .A( us10_n790 ) );
  NOR2_X1 us10_U283 (.ZN( us10_n653 ) , .A1( us10_n762 ) , .A2( us10_n786 ) );
  AOI21_X1 us10_U284 (.B1( us10_n625 ) , .ZN( us10_n627 ) , .A( us10_n763 ) , .B2( us10_n814 ) );
  AOI21_X1 us10_U285 (.ZN( us10_n478 ) , .B2( us10_n697 ) , .A( us10_n749 ) , .B1( us10_n779 ) );
  AOI21_X1 us10_U286 (.ZN( us10_n648 ) , .A( us10_n762 ) , .B2( us10_n784 ) , .B1( us10_n792 ) );
  AOI21_X1 us10_U287 (.ZN( us10_n623 ) , .B1( us10_n699 ) , .A( us10_n779 ) , .B2( us10_n784 ) );
  NOR2_X1 us10_U288 (.ZN( us10_n582 ) , .A1( us10_n744 ) , .A2( us10_n815 ) );
  NOR2_X1 us10_U289 (.A2( us10_n708 ) , .A1( us10_n762 ) , .ZN( us10_n794 ) );
  AOI221_X1 us10_U29 (.A( us10_n781 ) , .ZN( us10_n798 ) , .C2( us10_n837 ) , .B2( us10_n838 ) , .B1( us10_n865 ) , .C1( us10_n866 ) );
  NOR2_X1 us10_U290 (.ZN( us10_n553 ) , .A2( us10_n744 ) , .A1( us10_n784 ) );
  NOR2_X1 us10_U291 (.ZN( us10_n519 ) , .A2( us10_n699 ) , .A1( us10_n816 ) );
  AOI21_X1 us10_U292 (.ZN( us10_n626 ) , .B2( us10_n669 ) , .A( us10_n790 ) , .B1( us10_n791 ) );
  NOR2_X1 us10_U293 (.ZN( us10_n520 ) , .A2( us10_n708 ) , .A1( us10_n814 ) );
  AOI21_X1 us10_U294 (.ZN( us10_n477 ) , .A( us10_n669 ) , .B1( us10_n750 ) , .B2( us10_n806 ) );
  AOI21_X1 us10_U295 (.ZN( us10_n589 ) , .B2( us10_n699 ) , .B1( us10_n815 ) , .A( us10_n817 ) );
  AOI21_X1 us10_U296 (.ZN( us10_n510 ) , .B2( us10_n669 ) , .A( us10_n730 ) , .B1( us10_n815 ) );
  AOI21_X1 us10_U297 (.ZN( us10_n540 ) , .A( us10_n763 ) , .B2( us10_n779 ) , .B1( us10_n817 ) );
  AOI21_X1 us10_U298 (.ZN( us10_n515 ) , .A( us10_n729 ) , .B1( us10_n750 ) , .B2( us10_n803 ) );
  NOR2_X1 us10_U299 (.ZN( us10_n547 ) , .A1( us10_n699 ) , .A2( us10_n744 ) );
  NAND4_X1 us10_U3 (.ZN( sa13_sr_0 ) , .A4( us10_n501 ) , .A3( us10_n502 ) , .A2( us10_n503 ) , .A1( us10_n504 ) );
  NOR4_X1 us10_U30 (.A4( us10_n793 ) , .A3( us10_n794 ) , .A2( us10_n795 ) , .A1( us10_n796 ) , .ZN( us10_n797 ) );
  NOR2_X1 us10_U300 (.ZN( us10_n581 ) , .A1( us10_n669 ) , .A2( us10_n788 ) );
  AOI21_X1 us10_U301 (.ZN( us10_n539 ) , .B2( us10_n812 ) , .A( us10_n814 ) , .B1( us10_n815 ) );
  NOR2_X1 us10_U302 (.ZN( us10_n559 ) , .A2( us10_n791 ) , .A1( us10_n803 ) );
  AOI21_X1 us10_U303 (.ZN( us10_n498 ) , .A( us10_n724 ) , .B2( us10_n762 ) , .B1( us10_n814 ) );
  NAND2_X2 us10_U304 (.A2( us10_n461 ) , .A1( us10_n462 ) , .ZN( us10_n747 ) );
  AOI21_X1 us10_U305 (.B1( us10_n699 ) , .ZN( us10_n700 ) , .A( us10_n732 ) , .B2( us10_n763 ) );
  AOI21_X1 us10_U306 (.ZN( us10_n591 ) , .B2( us10_n763 ) , .A( us10_n785 ) , .B1( us10_n812 ) );
  AOI21_X1 us10_U307 (.ZN( us10_n640 ) , .B2( us10_n747 ) , .A( us10_n792 ) , .B1( us10_n803 ) );
  AOI21_X1 us10_U308 (.ZN( us10_n569 ) , .B1( us10_n750 ) , .B2( us10_n762 ) , .A( us10_n780 ) );
  NOR2_X1 us10_U309 (.ZN( us10_n683 ) , .A2( us10_n699 ) , .A1( us10_n803 ) );
  NOR4_X1 us10_U31 (.A4( us10_n776 ) , .A3( us10_n777 ) , .A1( us10_n778 ) , .ZN( us10_n799 ) , .A2( us10_n801 ) );
  NOR2_X1 us10_U310 (.ZN( us10_n665 ) , .A1( us10_n780 ) , .A2( us10_n813 ) );
  AOI21_X1 us10_U311 (.ZN( us10_n500 ) , .A( us10_n697 ) , .B1( us10_n708 ) , .B2( us10_n786 ) );
  NOR2_X1 us10_U312 (.ZN( us10_n685 ) , .A1( us10_n729 ) , .A2( us10_n816 ) );
  INV_X1 us10_U313 (.A( us10_n791 ) , .ZN( us10_n873 ) );
  AOI21_X1 us10_U314 (.ZN( us10_n649 ) , .B1( us10_n729 ) , .B2( us10_n763 ) , .A( us10_n813 ) );
  AOI21_X1 us10_U315 (.B1( us10_n686 ) , .ZN( us10_n687 ) , .A( us10_n728 ) , .B2( us10_n761 ) );
  INV_X1 us10_U316 (.A( us10_n699 ) , .ZN( us10_n853 ) );
  NOR2_X1 us10_U317 (.ZN( us10_n568 ) , .A1( us10_n729 ) , .A2( us10_n762 ) );
  NOR2_X1 us10_U318 (.ZN( us10_n578 ) , .A1( us10_n708 ) , .A2( us10_n813 ) );
  AOI21_X1 us10_U319 (.ZN( us10_n514 ) , .A( us10_n779 ) , .B2( us10_n792 ) , .B1( us10_n812 ) );
  NOR4_X1 us10_U32 (.A4( us10_n734 ) , .A3( us10_n735 ) , .A2( us10_n736 ) , .A1( us10_n737 ) , .ZN( us10_n738 ) );
  NOR2_X1 us10_U320 (.ZN( us10_n684 ) , .A1( us10_n791 ) , .A2( us10_n813 ) );
  NOR2_X1 us10_U321 (.ZN( us10_n580 ) , .A2( us10_n697 ) , .A1( us10_n791 ) );
  NOR2_X1 us10_U322 (.A2( us10_n813 ) , .A1( us10_n815 ) , .ZN( us10_n821 ) );
  NOR2_X1 us10_U323 (.ZN( us10_n566 ) , .A2( us10_n697 ) , .A1( us10_n763 ) );
  AOI21_X1 us10_U324 (.ZN( us10_n497 ) , .A( us10_n779 ) , .B2( us10_n791 ) , .B1( us10_n804 ) );
  AOI21_X1 us10_U325 (.ZN( us10_n564 ) , .B1( us10_n724 ) , .A( us10_n779 ) , .B2( us10_n791 ) );
  NOR2_X1 us10_U326 (.ZN( us10_n632 ) , .A2( us10_n697 ) , .A1( us10_n724 ) );
  NAND2_X2 us10_U327 (.A2( us10_n454 ) , .A1( us10_n472 ) , .ZN( us10_n779 ) );
  NOR2_X1 us10_U328 (.ZN( us10_n529 ) , .A1( us10_n708 ) , .A2( us10_n779 ) );
  AOI21_X1 us10_U329 (.ZN( us10_n639 ) , .B2( us10_n749 ) , .A( us10_n788 ) , .B1( us10_n812 ) );
  AOI211_X1 us10_U33 (.B( us10_n725 ) , .A( us10_n726 ) , .ZN( us10_n739 ) , .C1( us10_n843 ) , .C2( us10_n855 ) );
  AOI21_X1 us10_U330 (.ZN( us10_n689 ) , .B2( us10_n749 ) , .B1( us10_n763 ) , .A( us10_n806 ) );
  AOI21_X1 us10_U331 (.A( us10_n790 ) , .B2( us10_n791 ) , .B1( us10_n792 ) , .ZN( us10_n793 ) );
  AOI21_X1 us10_U332 (.A( us10_n733 ) , .ZN( us10_n734 ) , .B2( us10_n780 ) , .B1( us10_n792 ) );
  AOI21_X1 us10_U333 (.ZN( us10_n641 ) , .B1( us10_n680 ) , .A( us10_n791 ) , .B2( us10_n817 ) );
  NOR2_X1 us10_U334 (.ZN( us10_n583 ) , .A1( us10_n792 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U335 (.ZN( us10_n711 ) , .A1( us10_n762 ) , .A2( us10_n763 ) );
  NOR2_X1 us10_U336 (.ZN( us10_n534 ) , .A1( us10_n724 ) , .A2( us10_n788 ) );
  NOR2_X1 us10_U337 (.ZN( us10_n682 ) , .A2( us10_n708 ) , .A1( us10_n817 ) );
  INV_X1 us10_U338 (.A( us10_n697 ) , .ZN( us10_n838 ) );
  AOI21_X1 us10_U339 (.ZN( us10_n442 ) , .A( us10_n699 ) , .B1( us10_n733 ) , .B2( us10_n750 ) );
  NOR3_X1 us10_U34 (.A3( us10_n722 ) , .A1( us10_n723 ) , .ZN( us10_n740 ) , .A2( us10_n741 ) );
  NAND2_X2 us10_U340 (.A1( us10_n455 ) , .A2( us10_n462 ) , .ZN( us10_n750 ) );
  INV_X1 us10_U341 (.A( us10_n815 ) , .ZN( us10_n855 ) );
  OAI21_X1 us10_U342 (.A( us10_n613 ) , .ZN( us10_n616 ) , .B1( us10_n625 ) , .B2( us10_n784 ) );
  NAND2_X2 us10_U343 (.A1( us10_n462 ) , .A2( us10_n472 ) , .ZN( us10_n788 ) );
  OAI21_X1 us10_U344 (.A( us10_n698 ) , .ZN( us10_n702 ) , .B2( us10_n750 ) , .B1( us10_n804 ) );
  OAI21_X1 us10_U345 (.ZN( us10_n698 ) , .B2( us10_n833 ) , .B1( us10_n838 ) , .A( us10_n860 ) );
  INV_X1 us10_U346 (.A( us10_n785 ) , .ZN( us10_n846 ) );
  INV_X1 us10_U347 (.A( us10_n780 ) , .ZN( us10_n850 ) );
  OAI21_X1 us10_U348 (.A( us10_n787 ) , .B2( us10_n788 ) , .B1( us10_n789 ) , .ZN( us10_n795 ) );
  OAI21_X1 us10_U349 (.ZN( us10_n787 ) , .A( us10_n839 ) , .B1( us10_n863 ) , .B2( us10_n873 ) );
  NOR4_X1 us10_U35 (.A3( us10_n755 ) , .A2( us10_n756 ) , .A1( us10_n757 ) , .ZN( us10_n758 ) , .A4( us10_n869 ) );
  NAND2_X1 us10_U350 (.A1( us10_n729 ) , .A2( us10_n784 ) , .ZN( us10_n811 ) );
  NAND2_X1 us10_U351 (.ZN( us10_n671 ) , .A1( us10_n806 ) , .A2( us10_n816 ) );
  NAND2_X1 us10_U352 (.ZN( us10_n714 ) , .A1( us10_n728 ) , .A2( us10_n780 ) );
  AOI21_X1 us10_U353 (.ZN( us10_n443 ) , .B1( us10_n789 ) , .B2( us10_n791 ) , .A( us10_n814 ) );
  NOR2_X1 us10_U354 (.ZN( us10_n712 ) , .A2( us10_n724 ) , .A1( us10_n790 ) );
  NAND2_X1 us10_U355 (.A2( us10_n762 ) , .A1( us10_n806 ) , .ZN( us10_n810 ) );
  NAND2_X2 us10_U356 (.A1( us10_n454 ) , .A2( us10_n461 ) , .ZN( us10_n813 ) );
  NOR2_X1 us10_U357 (.ZN( us10_n470 ) , .A2( us10_n779 ) , .A1( us10_n815 ) );
  NAND2_X1 us10_U358 (.A1( us10_n699 ) , .A2( us10_n729 ) , .ZN( us10_n782 ) );
  NOR2_X1 us10_U359 (.ZN( us10_n526 ) , .A1( us10_n724 ) , .A2( us10_n750 ) );
  AOI211_X1 us10_U36 (.B( us10_n745 ) , .A( us10_n746 ) , .ZN( us10_n759 ) , .C1( us10_n832 ) , .C2( us10_n853 ) );
  NOR2_X1 us10_U360 (.ZN( us10_n518 ) , .A1( us10_n708 ) , .A2( us10_n788 ) );
  NAND2_X1 us10_U361 (.A2( us10_n749 ) , .A1( us10_n786 ) , .ZN( us10_n809 ) );
  INV_X1 us10_U362 (.A( us10_n817 ) , .ZN( us10_n844 ) );
  NAND2_X2 us10_U363 (.A1( us10_n451 ) , .A2( us10_n454 ) , .ZN( us10_n814 ) );
  INV_X1 us10_U364 (.A( us10_n724 ) , .ZN( us10_n856 ) );
  AND2_X1 us10_U365 (.ZN( us10_n732 ) , .A1( us10_n779 ) , .A2( us10_n785 ) );
  AOI221_X1 us10_U366 (.A( us10_n764 ) , .ZN( us10_n774 ) , .C2( us10_n810 ) , .B2( us10_n835 ) , .C1( us10_n855 ) , .B1( us10_n866 ) );
  AOI21_X1 us10_U367 (.B2( us10_n763 ) , .ZN( us10_n764 ) , .A( us10_n788 ) , .B1( us10_n792 ) );
  INV_X1 us10_U368 (.A( us10_n761 ) , .ZN( us10_n835 ) );
  NAND2_X1 us10_U369 (.A1( us10_n451 ) , .A2( us10_n471 ) , .ZN( us10_n816 ) );
  NOR3_X1 us10_U37 (.A3( us10_n741 ) , .A2( us10_n742 ) , .A1( us10_n743 ) , .ZN( us10_n760 ) );
  NAND2_X1 us10_U370 (.A2( us10_n441 ) , .A1( us10_n447 ) , .ZN( us10_n784 ) );
  NAND2_X1 us10_U371 (.A2( us10_n448 ) , .A1( us10_n460 ) , .ZN( us10_n728 ) );
  NAND2_X1 us10_U372 (.A1( us10_n453 ) , .A2( us10_n472 ) , .ZN( us10_n785 ) );
  NAND2_X1 us10_U373 (.A1( us10_n453 ) , .A2( us10_n461 ) , .ZN( us10_n744 ) );
  NAND2_X1 us10_U374 (.A1( us10_n452 ) , .A2( us10_n465 ) , .ZN( us10_n669 ) );
  NAND2_X1 us10_U375 (.A2( us10_n453 ) , .A1( us10_n455 ) , .ZN( us10_n806 ) );
  NAND2_X1 us10_U376 (.A1( us10_n441 ) , .A2( us10_n460 ) , .ZN( us10_n699 ) );
  NAND2_X1 us10_U377 (.A1( us10_n455 ) , .A2( us10_n471 ) , .ZN( us10_n803 ) );
  NAND2_X1 us10_U378 (.A2( us10_n464 ) , .A1( us10_n465 ) , .ZN( us10_n812 ) );
  NAND2_X1 us10_U379 (.A1( us10_n447 ) , .A2( us10_n448 ) , .ZN( us10_n786 ) );
  NAND4_X1 us10_U38 (.ZN( sa13_sr_3 ) , .A4( us10_n704 ) , .A3( us10_n705 ) , .A2( us10_n706 ) , .A1( us10_n707 ) );
  NAND2_X2 us10_U380 (.A2( us10_n461 ) , .A1( us10_n471 ) , .ZN( us10_n697 ) );
  NAND2_X1 us10_U381 (.A2( us10_n448 ) , .A1( us10_n452 ) , .ZN( us10_n729 ) );
  NAND2_X1 us10_U382 (.A2( us10_n449 ) , .A1( us10_n452 ) , .ZN( us10_n763 ) );
  NAND2_X1 us10_U383 (.A2( us10_n454 ) , .A1( us10_n455 ) , .ZN( us10_n730 ) );
  NOR2_X1 us10_U384 (.ZN( us10_n465 ) , .A2( us10_n847 ) , .A1( us10_n848 ) );
  NOR2_X1 us10_U385 (.ZN( us10_n453 ) , .A1( us10_n826 ) , .A2( us10_n827 ) );
  NOR2_X1 us10_U386 (.ZN( us10_n451 ) , .A1( us10_n828 ) , .A2( us10_n829 ) );
  NAND2_X1 us10_U387 (.A1( us10_n451 ) , .A2( us10_n462 ) , .ZN( us10_n790 ) );
  NAND2_X2 us10_U388 (.A2( us10_n448 ) , .A1( us10_n464 ) , .ZN( us10_n815 ) );
  NAND2_X2 us10_U389 (.A2( us10_n441 ) , .A1( us10_n452 ) , .ZN( us10_n791 ) );
  NOR4_X1 us10_U39 (.A4( us10_n700 ) , .A3( us10_n701 ) , .A2( us10_n702 ) , .A1( us10_n703 ) , .ZN( us10_n704 ) );
  NAND2_X2 us10_U390 (.A1( us10_n449 ) , .A2( us10_n464 ) , .ZN( us10_n724 ) );
  NAND2_X1 us10_U391 (.A1( us10_n447 ) , .A2( us10_n449 ) , .ZN( us10_n805 ) );
  NAND2_X2 us10_U392 (.A1( us10_n449 ) , .A2( us10_n460 ) , .ZN( us10_n792 ) );
  NAND2_X2 us10_U393 (.A1( us10_n441 ) , .A2( us10_n464 ) , .ZN( us10_n708 ) );
  NAND2_X2 us10_U394 (.A2( us10_n471 ) , .A1( us10_n472 ) , .ZN( us10_n817 ) );
  NAND2_X2 us10_U395 (.A2( us10_n460 ) , .A1( us10_n465 ) , .ZN( us10_n780 ) );
  NOR2_X1 us10_U396 (.ZN( us10_n447 ) , .A2( us10_n849 ) , .A1( us10_n858 ) );
  NOR2_X1 us10_U397 (.A2( sa10_6 ) , .A1( sa10_7 ) , .ZN( us10_n464 ) );
  NOR2_X1 us10_U398 (.A2( sa10_7 ) , .ZN( us10_n460 ) , .A1( us10_n849 ) );
  NOR2_X1 us10_U399 (.A2( sa10_4 ) , .ZN( us10_n449 ) , .A1( us10_n848 ) );
  NOR3_X1 us10_U4 (.ZN( us10_n598 ) , .A1( us10_n608 ) , .A3( us10_n723 ) , .A2( us10_n742 ) );
  AOI211_X1 us10_U40 (.B( us10_n694 ) , .A( us10_n695 ) , .ZN( us10_n705 ) , .C2( us10_n831 ) , .C1( us10_n851 ) );
  NOR2_X1 us10_U400 (.A2( sa10_4 ) , .A1( sa10_5 ) , .ZN( us10_n441 ) );
  NOR2_X1 us10_U401 (.A2( sa10_5 ) , .ZN( us10_n448 ) , .A1( us10_n847 ) );
  NOR2_X1 us10_U402 (.A2( sa10_1 ) , .ZN( us10_n471 ) , .A1( us10_n826 ) );
  NOR2_X1 us10_U403 (.A2( sa10_2 ) , .A1( sa10_3 ) , .ZN( us10_n472 ) );
  NOR2_X1 us10_U404 (.A2( sa10_6 ) , .ZN( us10_n452 ) , .A1( us10_n858 ) );
  NOR2_X1 us10_U405 (.A2( sa10_2 ) , .ZN( us10_n461 ) , .A1( us10_n829 ) );
  NOR2_X1 us10_U406 (.A2( sa10_3 ) , .ZN( us10_n455 ) , .A1( us10_n828 ) );
  INV_X1 us10_U407 (.A( sa10_6 ) , .ZN( us10_n849 ) );
  INV_X1 us10_U408 (.A( sa10_4 ) , .ZN( us10_n847 ) );
  INV_X1 us10_U409 (.A( sa10_3 ) , .ZN( us10_n829 ) );
  NOR2_X1 us10_U41 (.ZN( us10_n707 ) , .A2( us10_n776 ) , .A1( us10_n800 ) );
  INV_X1 us10_U410 (.A( sa10_2 ) , .ZN( us10_n828 ) );
  INV_X1 us10_U411 (.A( sa10_7 ) , .ZN( us10_n858 ) );
  INV_X1 us10_U412 (.A( sa10_5 ) , .ZN( us10_n848 ) );
  INV_X1 us10_U413 (.A( sa10_1 ) , .ZN( us10_n827 ) );
  INV_X1 us10_U414 (.A( sa10_0 ) , .ZN( us10_n826 ) );
  NOR2_X1 us10_U415 (.A2( sa10_0 ) , .A1( sa10_1 ) , .ZN( us10_n462 ) );
  NOR2_X1 us10_U416 (.A2( sa10_0 ) , .ZN( us10_n454 ) , .A1( us10_n827 ) );
  OAI222_X1 us10_U417 (.B2( us10_n747 ) , .B1( us10_n748 ) , .A2( us10_n749 ) , .ZN( us10_n757 ) , .C2( us10_n805 ) , .C1( us10_n814 ) , .A1( us10_n817 ) );
  OAI22_X1 us10_U418 (.B2( us10_n803 ) , .B1( us10_n804 ) , .A2( us10_n805 ) , .A1( us10_n806 ) , .ZN( us10_n808 ) );
  OAI21_X1 us10_U419 (.A( us10_n731 ) , .B1( us10_n732 ) , .ZN( us10_n736 ) , .B2( us10_n805 ) );
  NAND4_X1 us10_U42 (.ZN( sa13_sr_7 ) , .A4( us10_n822 ) , .A3( us10_n823 ) , .A2( us10_n824 ) , .A1( us10_n825 ) );
  OAI222_X1 us10_U420 (.ZN( us10_n505 ) , .C2( us10_n625 ) , .B2( us10_n647 ) , .B1( us10_n747 ) , .A2( us10_n748 ) , .C1( us10_n805 ) , .A1( us10_n806 ) );
  AOI21_X1 us10_U421 (.ZN( us10_n650 ) , .A( us10_n779 ) , .B1( us10_n792 ) , .B2( us10_n805 ) );
  INV_X1 us10_U422 (.A( us10_n805 ) , .ZN( us10_n860 ) );
  NOR2_X1 us10_U423 (.ZN( us10_n735 ) , .A2( us10_n803 ) , .A1( us10_n805 ) );
  NOR2_X1 us10_U424 (.ZN( us10_n484 ) , .A1( us10_n788 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U425 (.A2( us10_n744 ) , .ZN( us10_n755 ) , .A1( us10_n805 ) );
  NAND2_X1 us10_U426 (.ZN( us10_n753 ) , .A1( us10_n763 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U427 (.ZN( us10_n715 ) , .A1( us10_n805 ) , .A2( us10_n817 ) );
  NOR2_X1 us10_U428 (.ZN( us10_n567 ) , .A1( us10_n747 ) , .A2( us10_n805 ) );
  AOI21_X1 us10_U429 (.ZN( us10_n552 ) , .B1( us10_n669 ) , .A( us10_n697 ) , .B2( us10_n805 ) );
  NOR4_X1 us10_U43 (.A4( us10_n818 ) , .A3( us10_n819 ) , .A2( us10_n820 ) , .A1( us10_n821 ) , .ZN( us10_n822 ) );
  NOR2_X1 us10_U430 (.ZN( us10_n556 ) , .A1( us10_n762 ) , .A2( us10_n805 ) );
  NOR2_X1 us10_U431 (.ZN( us10_n670 ) , .A1( us10_n790 ) , .A2( us10_n805 ) );
  AND2_X1 us10_U432 (.ZN( us10_n438 ) , .A2( us10_n831 ) , .A1( us10_n854 ) );
  AND2_X1 us10_U433 (.ZN( us10_n439 ) , .A2( us10_n843 ) , .A1( us10_n861 ) );
  NOR3_X1 us10_U434 (.A1( us10_n438 ) , .A2( us10_n439 ) , .A3( us10_n576 ) , .ZN( us10_n587 ) );
  NAND4_X1 us10_U435 (.ZN( sa13_sr_2 ) , .A4( us10_n643 ) , .A3( us10_n644 ) , .A2( us10_n645 ) , .A1( us10_n646 ) );
  INV_X1 us10_U436 (.A( us10_n812 ) , .ZN( us10_n854 ) );
  NAND3_X1 us10_U437 (.ZN( sa13_sr_6 ) , .A3( us10_n797 ) , .A2( us10_n798 ) , .A1( us10_n799 ) );
  NAND3_X1 us10_U438 (.ZN( sa13_sr_5 ) , .A3( us10_n758 ) , .A2( us10_n759 ) , .A1( us10_n760 ) );
  NAND3_X1 us10_U439 (.ZN( sa13_sr_4 ) , .A3( us10_n738 ) , .A2( us10_n739 ) , .A1( us10_n740 ) );
  AOI222_X1 us10_U44 (.C2( us10_n809 ) , .B2( us10_n810 ) , .A2( us10_n811 ) , .ZN( us10_n823 ) , .C1( us10_n832 ) , .A1( us10_n839 ) , .B1( us10_n853 ) );
  NAND3_X1 us10_U440 (.A3( us10_n675 ) , .A2( us10_n676 ) , .A1( us10_n677 ) , .ZN( us10_n807 ) );
  NAND3_X1 us10_U441 (.ZN( us10_n638 ) , .A3( us10_n708 ) , .A2( us10_n724 ) , .A1( us10_n792 ) );
  NAND3_X1 us10_U442 (.A3( us10_n618 ) , .A2( us10_n619 ) , .A1( us10_n620 ) , .ZN( us10_n725 ) );
  NAND3_X1 us10_U443 (.A3( us10_n585 ) , .A2( us10_n586 ) , .A1( us10_n587 ) , .ZN( us10_n621 ) );
  NAND3_X1 us10_U444 (.ZN( us10_n565 ) , .A3( us10_n680 ) , .A2( us10_n750 ) , .A1( us10_n785 ) );
  NAND3_X1 us10_U445 (.A3( us10_n523 ) , .A2( us10_n524 ) , .A1( us10_n525 ) , .ZN( us10_n742 ) );
  NAND3_X1 us10_U446 (.A3( us10_n512 ) , .A1( us10_n513 ) , .ZN( us10_n608 ) , .A2( us10_n871 ) );
  NAND3_X1 us10_U447 (.A3( us10_n467 ) , .A2( us10_n468 ) , .A1( us10_n469 ) , .ZN( us10_n777 ) );
  INV_X1 us10_U448 (.A( us10_n803 ) , .ZN( us10_n843 ) );
  AOI21_X1 us10_U449 (.ZN( us10_n576 ) , .B2( us10_n724 ) , .B1( us10_n748 ) , .A( us10_n785 ) );
  AOI211_X1 us10_U45 (.B( us10_n807 ) , .A( us10_n808 ) , .ZN( us10_n824 ) , .C1( us10_n842 ) , .C2( us10_n850 ) );
  NOR4_X1 us10_U46 (.A4( us10_n498 ) , .A3( us10_n499 ) , .A2( us10_n500 ) , .ZN( us10_n501 ) , .A1( us10_n527 ) );
  AOI221_X1 us10_U47 (.A( us10_n497 ) , .ZN( us10_n502 ) , .B2( us10_n843 ) , .C1( us10_n846 ) , .C2( us10_n860 ) , .B1( us10_n862 ) );
  AOI211_X1 us10_U48 (.A( us10_n496 ) , .ZN( us10_n503 ) , .B( us10_n802 ) , .C2( us10_n839 ) , .C1( us10_n851 ) );
  NAND4_X1 us10_U49 (.ZN( sa13_sr_1 ) , .A4( us10_n595 ) , .A3( us10_n596 ) , .A2( us10_n597 ) , .A1( us10_n598 ) );
  NOR3_X1 us10_U5 (.A3( us10_n800 ) , .A2( us10_n801 ) , .A1( us10_n802 ) , .ZN( us10_n825 ) );
  NOR4_X1 us10_U50 (.A4( us10_n591 ) , .A3( us10_n592 ) , .A2( us10_n593 ) , .A1( us10_n594 ) , .ZN( us10_n595 ) );
  AOI211_X1 us10_U51 (.B( us10_n589 ) , .A( us10_n590 ) , .ZN( us10_n596 ) , .C2( us10_n811 ) , .C1( us10_n833 ) );
  AOI211_X1 us10_U52 (.A( us10_n588 ) , .ZN( us10_n597 ) , .B( us10_n621 ) , .C1( us10_n845 ) , .C2( us10_n855 ) );
  NOR2_X1 us10_U53 (.ZN( us10_n804 ) , .A1( us10_n854 ) , .A2( us10_n861 ) );
  NOR2_X1 us10_U54 (.ZN( us10_n625 ) , .A2( us10_n836 ) , .A1( us10_n839 ) );
  AOI222_X1 us10_U55 (.ZN( us10_n469 ) , .B1( us10_n832 ) , .A1( us10_n839 ) , .C1( us10_n842 ) , .C2( us10_n851 ) , .A2( us10_n855 ) , .B2( us10_n865 ) );
  NOR4_X1 us10_U56 (.A1( us10_n466 ) , .ZN( us10_n467 ) , .A4( us10_n542 ) , .A2( us10_n554 ) , .A3( us10_n614 ) );
  AOI221_X1 us10_U57 (.ZN( us10_n468 ) , .C2( us10_n714 ) , .B2( us10_n831 ) , .C1( us10_n845 ) , .B1( us10_n860 ) , .A( us10_n864 ) );
  NAND4_X1 us10_U58 (.A4( us10_n603 ) , .A3( us10_n604 ) , .A2( us10_n605 ) , .A1( us10_n606 ) , .ZN( us10_n722 ) );
  NOR3_X1 us10_U59 (.A1( us10_n599 ) , .ZN( us10_n604 ) , .A3( us10_n663 ) , .A2( us10_n770 ) );
  NOR3_X1 us10_U6 (.ZN( us10_n504 ) , .A2( us10_n679 ) , .A3( us10_n777 ) , .A1( us10_n876 ) );
  NOR4_X1 us10_U60 (.A3( us10_n600 ) , .A2( us10_n601 ) , .A1( us10_n602 ) , .ZN( us10_n603 ) , .A4( us10_n655 ) );
  AOI222_X1 us10_U61 (.ZN( us10_n606 ) , .A1( us10_n830 ) , .C2( us10_n837 ) , .B1( us10_n842 ) , .A2( us10_n856 ) , .B2( us10_n861 ) , .C1( us10_n868 ) );
  AOI222_X1 us10_U62 (.B2( us10_n638 ) , .ZN( us10_n644 ) , .B1( us10_n841 ) , .A1( us10_n842 ) , .C2( us10_n846 ) , .C1( us10_n863 ) , .A2( us10_n865 ) );
  NOR4_X1 us10_U63 (.A4( us10_n639 ) , .A3( us10_n640 ) , .A2( us10_n641 ) , .A1( us10_n642 ) , .ZN( us10_n643 ) );
  NOR3_X1 us10_U64 (.A2( us10_n607 ) , .A1( us10_n608 ) , .ZN( us10_n646 ) , .A3( us10_n722 ) );
  NAND4_X1 us10_U65 (.A4( us10_n657 ) , .A3( us10_n658 ) , .A2( us10_n659 ) , .A1( us10_n660 ) , .ZN( us10_n800 ) );
  NOR3_X1 us10_U66 (.A3( us10_n648 ) , .A2( us10_n649 ) , .A1( us10_n650 ) , .ZN( us10_n659 ) );
  NOR3_X1 us10_U67 (.A3( us10_n651 ) , .A2( us10_n652 ) , .A1( us10_n653 ) , .ZN( us10_n658 ) );
  NOR3_X1 us10_U68 (.A3( us10_n654 ) , .A2( us10_n655 ) , .A1( us10_n656 ) , .ZN( us10_n657 ) );
  NAND4_X1 us10_U69 (.A4( us10_n560 ) , .A3( us10_n561 ) , .A2( us10_n562 ) , .A1( us10_n563 ) , .ZN( us10_n607 ) );
  INV_X1 us10_U7 (.A( us10_n706 ) , .ZN( us10_n876 ) );
  NOR4_X1 us10_U70 (.A4( us10_n552 ) , .A3( us10_n553 ) , .A2( us10_n554 ) , .A1( us10_n555 ) , .ZN( us10_n562 ) );
  NOR4_X1 us10_U71 (.A4( us10_n556 ) , .A3( us10_n557 ) , .A2( us10_n558 ) , .A1( us10_n559 ) , .ZN( us10_n560 ) );
  NOR4_X1 us10_U72 (.ZN( us10_n561 ) , .A1( us10_n653 ) , .A3( us10_n661 ) , .A4( us10_n685 ) , .A2( us10_n768 ) );
  NAND4_X1 us10_U73 (.A4( us10_n772 ) , .A3( us10_n773 ) , .A2( us10_n774 ) , .A1( us10_n775 ) , .ZN( us10_n801 ) );
  NOR3_X1 us10_U74 (.A3( us10_n765 ) , .A2( us10_n766 ) , .A1( us10_n767 ) , .ZN( us10_n773 ) );
  NOR4_X1 us10_U75 (.A4( us10_n768 ) , .A3( us10_n769 ) , .A2( us10_n770 ) , .A1( us10_n771 ) , .ZN( us10_n772 ) );
  AOI222_X1 us10_U76 (.ZN( us10_n775 ) , .A1( us10_n830 ) , .C1( us10_n834 ) , .B2( us10_n841 ) , .A2( us10_n850 ) , .B1( us10_n861 ) , .C2( us10_n873 ) );
  NOR4_X1 us10_U77 (.A4( us10_n665 ) , .A3( us10_n666 ) , .A2( us10_n667 ) , .A1( us10_n668 ) , .ZN( us10_n676 ) );
  NOR4_X1 us10_U78 (.A4( us10_n661 ) , .A3( us10_n662 ) , .A2( us10_n663 ) , .A1( us10_n664 ) , .ZN( us10_n677 ) );
  NOR4_X1 us10_U79 (.A3( us10_n673 ) , .A1( us10_n674 ) , .ZN( us10_n675 ) , .A4( us10_n715 ) , .A2( us10_n859 ) );
  NOR3_X1 us10_U8 (.A3( us10_n621 ) , .A2( us10_n622 ) , .ZN( us10_n636 ) , .A1( us10_n725 ) );
  NOR2_X1 us10_U80 (.ZN( us10_n761 ) , .A1( us10_n833 ) , .A2( us10_n834 ) );
  NOR4_X1 us10_U81 (.A4( us10_n577 ) , .A3( us10_n578 ) , .A2( us10_n579 ) , .ZN( us10_n586 ) , .A1( us10_n683 ) );
  NOR4_X1 us10_U82 (.A1( us10_n584 ) , .ZN( us10_n585 ) , .A3( us10_n652 ) , .A2( us10_n662 ) , .A4( us10_n767 ) );
  AOI222_X1 us10_U83 (.ZN( us10_n513 ) , .C1( us10_n832 ) , .B2( us10_n837 ) , .A2( us10_n843 ) , .C2( us10_n862 ) , .B1( us10_n863 ) , .A1( us10_n866 ) );
  NOR4_X1 us10_U84 (.A4( us10_n509 ) , .A2( us10_n510 ) , .A1( us10_n511 ) , .ZN( us10_n512 ) , .A3( us10_n670 ) );
  INV_X1 us10_U85 (.A( us10_n505 ) , .ZN( us10_n871 ) );
  NAND4_X1 us10_U86 (.A4( us10_n456 ) , .A3( us10_n457 ) , .A2( us10_n458 ) , .A1( us10_n459 ) , .ZN( us10_n679 ) );
  NOR3_X1 us10_U87 (.ZN( us10_n457 ) , .A3( us10_n530 ) , .A1( us10_n555 ) , .A2( us10_n570 ) );
  NOR4_X1 us10_U88 (.ZN( us10_n458 ) , .A2( us10_n509 ) , .A1( us10_n599 ) , .A4( us10_n628 ) , .A3( us10_n711 ) );
  NOR4_X1 us10_U89 (.ZN( us10_n456 ) , .A2( us10_n517 ) , .A1( us10_n543 ) , .A3( us10_n579 ) , .A4( us10_n615 ) );
  NOR2_X1 us10_U9 (.ZN( us10_n575 ) , .A1( us10_n622 ) , .A2( us10_n745 ) );
  NAND4_X1 us10_U90 (.A4( us10_n535 ) , .A3( us10_n536 ) , .A2( us10_n537 ) , .A1( us10_n538 ) , .ZN( us10_n622 ) );
  NOR4_X1 us10_U91 (.A4( us10_n526 ) , .A2( us10_n527 ) , .A1( us10_n528 ) , .ZN( us10_n538 ) , .A3( us10_n701 ) );
  NOR4_X1 us10_U92 (.A1( us10_n531 ) , .ZN( us10_n536 ) , .A2( us10_n654 ) , .A4( us10_n668 ) , .A3( us10_n765 ) );
  NOR4_X1 us10_U93 (.A4( us10_n529 ) , .A3( us10_n530 ) , .ZN( us10_n537 ) , .A2( us10_n684 ) , .A1( us10_n794 ) );
  NOR2_X1 us10_U94 (.ZN( us10_n686 ) , .A1( us10_n831 ) , .A2( us10_n832 ) );
  NAND4_X1 us10_U95 (.A4( us10_n479 ) , .A3( us10_n480 ) , .A2( us10_n481 ) , .A1( us10_n482 ) , .ZN( us10_n694 ) );
  NOR3_X1 us10_U96 (.ZN( us10_n480 ) , .A2( us10_n508 ) , .A3( us10_n601 ) , .A1( us10_n610 ) );
  AOI211_X1 us10_U97 (.B( us10_n477 ) , .A( us10_n478 ) , .ZN( us10_n482 ) , .C2( us10_n833 ) , .C1( us10_n861 ) );
  NOR4_X1 us10_U98 (.ZN( us10_n481 ) , .A3( us10_n532 ) , .A4( us10_n545 ) , .A2( us10_n567 ) , .A1( us10_n717 ) );
  NAND4_X1 us10_U99 (.A4( us10_n548 ) , .A3( us10_n549 ) , .A2( us10_n550 ) , .A1( us10_n551 ) , .ZN( us10_n745 ) );
endmodule

