module des_des_die_3 ( u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_K12_19, u0_K12_35, u0_K12_36, u0_K13_41, 
       u0_K15_13, u0_K16_38, u0_K1_13, u0_K1_14, u0_K1_17, u0_K2_29, u0_K2_30, u0_K2_31, u0_K3_12, 
       u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_5, u0_K3_6, u0_K6_11, u0_K6_13, u0_K6_19, 
       u0_K6_20, u0_K6_23, u0_K6_24, u0_K6_41, u0_R0_18, u0_R0_19, u0_R0_20, u0_R0_21, u0_R0_28, 
       u0_R10_12, u0_R10_14, u0_R10_16, u0_R10_17, u0_R10_20, u0_R10_21, u0_R10_24, u0_R10_25, u0_R10_28, 
       u0_R10_29, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_2, 
       u0_R11_28, u0_R11_3, u0_R11_32, u0_R11_5, u0_R11_6, u0_R12_30, u0_R13_8, u0_R1_1, u0_R1_12, 
       u0_R1_13, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R4_1, u0_R4_12, 
       u0_R4_13, u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_24, u0_R4_25, 
       u0_R4_26, u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, u0_R4_4, u0_R4_5, 
       u0_R4_8, u0_R4_9, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_4, 
       u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_15, u0_desIn_r_23, u0_desIn_r_29, u0_desIn_r_3, 
       u0_desIn_r_31, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_63, u0_desIn_r_7, 
       u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_19, u0_key_r_20, u0_key_r_4, u0_key_r_41, u0_key_r_47, u0_key_r_48, 
       u0_key_r_5, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, 
       u0_u10_X_21, u0_u10_X_22, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, u0_u11_X_18, u0_u11_X_20, u0_u11_X_22, 
       u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, 
       u0_u12_X_2, u0_u12_X_24, u0_u12_X_37, u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, 
       u0_u12_X_46, u0_u12_X_48, u0_u12_X_5, u0_u12_X_7, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, u0_u13_X_48, 
       u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, u0_u14_X_18, u0_u14_X_19, u0_u14_X_20, 
       u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_42, u0_u1_X_25, 
       u0_u1_X_26, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, u0_u1_X_36, u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_40, 
       u0_u1_X_42, u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_3, u0_u2_X_9, u0_u5_X_10, u0_u5_X_15, u0_u5_X_16, 
       u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, u0_u5_X_9, u0_uk_K_r0_15, u0_uk_K_r0_28, 
       u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_41, u0_uk_K_r10_44, 
       u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_39, 
       u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_25, u0_uk_K_r14_15, u0_uk_K_r14_2, u0_uk_K_r14_50, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, 
       u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_33, u0_uk_K_r9_6, u0_uk_n100, 
       u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n101, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n109, 
       u0_uk_n115, u0_uk_n118, u0_uk_n121, u0_uk_n122, u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n131, u0_uk_n139, 
       u0_uk_n143, u0_uk_n144, u0_uk_n146, u0_uk_n148, u0_uk_n153, u0_uk_n155, u0_uk_n161, u0_uk_n164, u0_uk_n172, 
       u0_uk_n173, u0_uk_n179, u0_uk_n180, u0_uk_n187, u0_uk_n188, u0_uk_n190, u0_uk_n191, u0_uk_n195, u0_uk_n196, 
       u0_uk_n197, u0_uk_n200, u0_uk_n201, u0_uk_n206, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, u0_uk_n221, 
       u0_uk_n225, u0_uk_n230, u0_uk_n240, u0_uk_n257, u0_uk_n410, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n414, 
       u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n428, u0_uk_n429, 
       u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, u0_uk_n439, u0_uk_n440, u0_uk_n442, 
       u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n450, u0_uk_n547, u0_uk_n552, u0_uk_n557, u0_uk_n562, 
       u0_uk_n565, u0_uk_n568, u0_uk_n573, u0_uk_n578, u0_uk_n58, u0_uk_n63, u0_uk_n632, u0_uk_n643, u0_uk_n657, 
       u0_uk_n670, u0_uk_n674, u0_uk_n684, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, u0_uk_n786, u0_uk_n793, 
       u0_uk_n799, u0_uk_n8, u0_uk_n800, u0_uk_n83, u0_uk_n869, u0_uk_n892, u0_uk_n898, u0_uk_n91, u0_uk_n92, 
       u0_uk_n93, u0_uk_n94, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n976, u0_uk_n982, u0_uk_n99, 
       u0_uk_n999, u1_FP_40, u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, 
       u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, u1_K10_44, u1_K10_47, u1_K10_48, 
       u1_K11_11, u1_K11_13, u1_K11_2, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, u1_K11_7, 
       u1_K13_14, u1_K13_17, u1_K13_18, u1_K13_20, u1_K13_48, u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_42, 
       u1_K14_44, u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, u1_K15_2, 
       u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, u1_K15_36, 
       u1_K15_37, u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, u1_K16_13, 
       u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_20, u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_35, 
       u1_K1_1, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_20, u1_K2_23, u1_K2_24, u1_K2_25, 
       u1_K2_26, u1_K2_29, u1_K2_30, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, u1_K2_48, u1_K3_1, 
       u1_K3_2, u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, 
       u1_K3_5, u1_K3_6, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_6, u1_K5_19, u1_K5_23, u1_K5_24, 
       u1_K6_25, u1_K6_26, u1_K6_29, u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K7_1, 
       u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_2, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, 
       u1_K7_44, u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_7, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_29, 
       u1_K9_31, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, u1_K9_6, 
       u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, u1_R0_21, u1_R0_28, u1_R0_29, 
       u1_R0_32, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, 
       u1_R12_1, u1_R12_29, u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, 
       u1_R13_24, u1_R13_25, u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, 
       u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_32, u1_R1_4, u1_R1_5, u1_R2_1, u1_R2_2, 
       u1_R2_32, u1_R2_5, u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, 
       u1_R3_17, u1_R4_16, u1_R4_17, u1_R4_20, u1_R4_21, u1_R4_24, u1_R4_25, u1_R5_1, u1_R5_12, 
       u1_R5_13, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, 
       u1_R5_8, u1_R5_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, 
       u1_R7_20, u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, u1_R8_1, 
       u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R9_1, 
       u1_R9_12, u1_R9_20, u1_R9_21, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, 
       u1_desIn_r_25, u1_desIn_r_39, u1_desIn_r_57, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_2, u1_u0_X_3, u1_u0_X_31, 
       u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, 
       u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, u1_u0_X_48, u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, 
       u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, u1_u10_X_18, u1_u10_X_3, u1_u10_X_33, u1_u10_X_39, u1_u10_X_4, 
       u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, u1_u10_X_47, u1_u10_X_6, 
       u1_u10_X_8, u1_u10_X_9, u1_u12_X_1, u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, 
       u1_u12_X_3, u1_u12_X_4, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, u1_u12_X_9, u1_u13_X_10, 
       u1_u13_X_11, u1_u13_X_12, u1_u13_X_3, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, u1_u13_X_4, u1_u13_X_40, u1_u13_X_41, 
       u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, u1_u14_X_1, 
       u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, u1_u14_X_22, u1_u14_X_27, u1_u14_X_28, 
       u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, 
       u1_u14_X_9, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, u1_u15_X_22, u1_u15_X_23, u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, 
       u1_u15_X_27, u1_u15_X_28, u1_u15_X_33, u1_u15_X_36, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_37, 
       u1_u1_X_38, u1_u1_X_39, u1_u1_X_40, u1_u1_X_45, u1_u1_X_46, u1_u2_X_3, u1_u2_X_39, u1_u2_X_4, u1_u2_X_40, 
       u1_u2_X_45, u1_u2_X_46, u1_u3_X_4, u1_u3_X_5, u1_u3_X_7, u1_u3_X_9, u1_u4_X_21, u1_u5_X_27, u1_u5_X_28, 
       u1_u5_X_33, u1_u5_X_34, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_3, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, 
       u1_u6_X_45, u1_u6_X_9, u1_u8_X_21, u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, 
       u1_u8_X_39, u1_u8_X_4, u1_u8_X_40, u1_u8_X_45, u1_u8_X_46, u1_u9_X_34, u1_u9_X_39, u1_u9_X_40, u1_u9_X_45, 
       u1_u9_X_46, u1_uk_n1015, u1_uk_n1025, u1_uk_n1031, u1_uk_n1050, u1_uk_n1061, u1_uk_n1065, u1_uk_n1070, u1_uk_n1073, 
       u1_uk_n1074, u1_uk_n1105, u1_uk_n1106, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1154, u1_uk_n1155, 
       u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, u1_uk_n1166, u1_uk_n1167, u1_uk_n1170, 
       u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n437, u1_uk_n443, 
       u1_uk_n454, u1_uk_n496, u1_uk_n672, u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, 
       u1_uk_n949, u1_uk_n950, u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, 
       u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, u2_FP_48, u2_FP_49, 
       u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, u2_FP_64, u2_K11_11, 
       u2_K11_13, u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, u2_K16_19, 
       u2_K16_2, u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, u2_K16_32, 
       u2_K16_35, u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, u2_K16_5, 
       u2_K16_6, u2_K16_7, u2_K16_8, u2_K8_1, u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, 
       u2_K8_19, u2_K8_2, u2_K8_20, u2_K8_47, u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, 
       u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, 
       u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_22, u2_R7_24, u2_R7_25, 
       u2_R7_28, u2_R7_29, u2_R9_12, u2_R9_8, u2_R9_9, u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, u2_u10_X_18, 
       u2_u10_X_7, u2_u10_X_8, u2_u10_X_9, u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, u2_u15_X_22, u2_u15_X_27, 
       u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, u2_u15_X_46, u2_u15_X_9, 
       u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, u2_u7_X_44, 
       u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, u2_u8_X_31, u2_u8_X_32, u2_u8_X_34, u2_u8_X_39, u2_u8_X_40, u2_u8_X_45, 
       u2_u8_X_46, u2_u8_X_47, u2_uk_K_r7_0, u2_uk_n1098, u2_uk_n1110, u2_uk_n1113, u2_uk_n1132, u2_uk_n1133, u2_uk_n1136, 
       u2_uk_n1137, u2_uk_n1140, u2_uk_n155, u2_uk_n1585, u2_uk_n214, u2_uk_n313, u2_uk_n319, u2_uk_n335, u2_uk_n955, 
       u2_uk_n958, u2_uk_n959, u2_uk_n963, u0_out0_1, u0_out0_10, u0_out0_13, u0_out0_16, u0_out0_17, u0_out0_18, u0_out0_2, u0_out0_20, u0_out0_23, 
        u0_out0_24, u0_out0_26, u0_out0_28, u0_out0_30, u0_out0_31, u0_out0_6, u0_out0_9, u0_out10_1, u0_out10_10, 
        u0_out10_13, u0_out10_16, u0_out10_18, u0_out10_2, u0_out10_20, u0_out10_24, u0_out10_26, u0_out10_28, u0_out10_30, 
        u0_out10_6, u0_out11_1, u0_out11_10, u0_out11_11, u0_out11_12, u0_out11_16, u0_out11_19, u0_out11_20, u0_out11_22, 
        u0_out11_24, u0_out11_26, u0_out11_29, u0_out11_30, u0_out11_32, u0_out11_4, u0_out11_6, u0_out11_7, u0_out12_1, 
        u0_out12_10, u0_out12_12, u0_out12_13, u0_out12_15, u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_2, u0_out12_20, 
        u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_26, u0_out12_27, u0_out12_28, u0_out12_30, u0_out12_31, 
        u0_out12_32, u0_out12_5, u0_out12_6, u0_out12_7, u0_out12_9, u0_out13_15, u0_out13_21, u0_out13_27, u0_out13_5, 
        u0_out14_1, u0_out14_10, u0_out14_13, u0_out14_16, u0_out14_18, u0_out14_2, u0_out14_20, u0_out14_24, u0_out14_26, 
        u0_out14_28, u0_out14_30, u0_out14_6, u0_out15_12, u0_out15_22, u0_out15_32, u0_out15_7, u0_out1_11, u0_out1_12, 
        u0_out1_14, u0_out1_19, u0_out1_22, u0_out1_25, u0_out1_29, u0_out1_3, u0_out1_32, u0_out1_4, u0_out1_7, 
        u0_out1_8, u0_out2_13, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_2, u0_out2_23, u0_out2_24, u0_out2_28, 
        u0_out2_30, u0_out2_31, u0_out2_6, u0_out2_9, u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, u0_out5_13, 
        u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, u0_out5_21, 
        u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_3, 
        u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, u0_out5_9, 
        u0_uk_n10, u0_uk_n102, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, 
        u0_uk_n147, u0_uk_n162, u0_uk_n163, u0_uk_n182, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n217, 
        u0_uk_n220, u0_uk_n222, u0_uk_n231, u0_uk_n238, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n31, 
        u0_uk_n60, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_15, u1_out0_17, u1_out0_18, u1_out0_19, u1_out0_2, 
        u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_27, u1_out0_28, u1_out0_29, u1_out0_31, u1_out0_32, u1_out0_4, 
        u1_out0_5, u1_out0_7, u1_out0_9, u1_out10_11, u1_out10_12, u1_out10_13, u1_out10_15, u1_out10_16, u1_out10_17, 
        u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_21, u1_out10_22, u1_out10_23, u1_out10_24, u1_out10_27, u1_out10_28, 
        u1_out10_29, u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_9, 
        u1_out12_1, u1_out12_10, u1_out12_13, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_2, u1_out12_20, 
        u1_out12_21, u1_out12_23, u1_out12_24, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_30, u1_out12_31, u1_out12_5, 
        u1_out12_6, u1_out12_9, u1_out13_12, u1_out13_13, u1_out13_15, u1_out13_17, u1_out13_18, u1_out13_2, u1_out13_21, 
        u1_out13_22, u1_out13_23, u1_out13_27, u1_out13_28, u1_out13_31, u1_out13_32, u1_out13_5, u1_out13_7, u1_out13_9, 
        u1_out14_1, u1_out14_10, u1_out14_11, u1_out14_12, u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, 
        u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_20, u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, 
        u1_out14_26, u1_out14_27, u1_out14_28, u1_out14_29, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, 
        u1_out14_5, u1_out14_6, u1_out14_7, u1_out14_8, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_14, 
        u1_out15_16, u1_out15_19, u1_out15_20, u1_out15_24, u1_out15_25, u1_out15_26, u1_out15_29, u1_out15_3, u1_out15_30, 
        u1_out15_4, u1_out15_6, u1_out15_8, u1_out1_1, u1_out1_10, u1_out1_12, u1_out1_14, u1_out1_15, u1_out1_20, 
        u1_out1_21, u1_out1_22, u1_out1_25, u1_out1_26, u1_out1_27, u1_out1_3, u1_out1_32, u1_out1_5, u1_out1_7, 
        u1_out1_8, u1_out2_12, u1_out2_15, u1_out2_17, u1_out2_21, u1_out2_22, u1_out2_23, u1_out2_27, u1_out2_31, 
        u1_out2_32, u1_out2_5, u1_out2_7, u1_out2_9, u1_out3_13, u1_out3_17, u1_out3_18, u1_out3_2, u1_out3_23, 
        u1_out3_28, u1_out3_31, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_20, u1_out4_26, u1_out5_11, u1_out5_14, 
        u1_out5_19, u1_out5_25, u1_out5_29, u1_out5_3, u1_out5_4, u1_out5_8, u1_out6_12, u1_out6_13, u1_out6_15, 
        u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_2, u1_out6_21, u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_27, 
        u1_out6_28, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_9, u1_out8_1, 
        u1_out8_10, u1_out8_11, u1_out8_12, u1_out8_14, u1_out8_15, u1_out8_17, u1_out8_19, u1_out8_20, u1_out8_21, 
        u1_out8_22, u1_out8_23, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_29, u1_out8_3, u1_out8_31, u1_out8_32, 
        u1_out8_4, u1_out8_5, u1_out8_7, u1_out8_8, u1_out8_9, u1_out9_11, u1_out9_12, u1_out9_15, u1_out9_19, 
        u1_out9_21, u1_out9_22, u1_out9_27, u1_out9_29, u1_out9_32, u1_out9_4, u1_out9_5, u1_out9_7, u2_out10_13, 
        u2_out10_16, u2_out10_18, u2_out10_2, u2_out10_24, u2_out10_28, u2_out10_30, u2_out10_6, u2_out15_1, u2_out15_10, 
        u2_out15_11, u2_out15_12, u2_out15_13, u2_out15_14, u2_out15_15, u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_19, 
        u2_out15_2, u2_out15_20, u2_out15_21, u2_out15_22, u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_27, 
        u2_out15_28, u2_out15_29, u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_6, 
        u2_out15_7, u2_out15_8, u2_out15_9, u2_out7_1, u2_out7_10, u2_out7_13, u2_out7_15, u2_out7_16, u2_out7_17, 
        u2_out7_18, u2_out7_2, u2_out7_20, u2_out7_21, u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_27, u2_out7_28, 
        u2_out7_30, u2_out7_31, u2_out7_5, u2_out7_6, u2_out7_9, u2_out8_11, u2_out8_12, u2_out8_15, u2_out8_19, 
        u2_out8_21, u2_out8_22, u2_out8_27, u2_out8_29, u2_out8_32, u2_out8_4, u2_out8_5, u2_out8_7 );
  input u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_K12_19, u0_K12_35, u0_K12_36, u0_K13_41, 
        u0_K15_13, u0_K16_38, u0_K1_13, u0_K1_14, u0_K1_17, u0_K2_29, u0_K2_30, u0_K2_31, u0_K3_12, 
        u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_5, u0_K3_6, u0_K6_11, u0_K6_13, u0_K6_19, 
        u0_K6_20, u0_K6_23, u0_K6_24, u0_K6_41, u0_R0_18, u0_R0_19, u0_R0_20, u0_R0_21, u0_R0_28, 
        u0_R10_12, u0_R10_14, u0_R10_16, u0_R10_17, u0_R10_20, u0_R10_21, u0_R10_24, u0_R10_25, u0_R10_28, 
        u0_R10_29, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_2, 
        u0_R11_28, u0_R11_3, u0_R11_32, u0_R11_5, u0_R11_6, u0_R12_30, u0_R13_8, u0_R1_1, u0_R1_12, 
        u0_R1_13, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R4_1, u0_R4_12, 
        u0_R4_13, u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_24, u0_R4_25, 
        u0_R4_26, u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, u0_R4_4, u0_R4_5, 
        u0_R4_8, u0_R4_9, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_4, 
        u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_15, u0_desIn_r_23, u0_desIn_r_29, u0_desIn_r_3, 
        u0_desIn_r_31, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_63, u0_desIn_r_7, 
        u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_19, u0_key_r_20, u0_key_r_4, u0_key_r_41, u0_key_r_47, u0_key_r_48, 
        u0_key_r_5, u0_key_r_54, u0_key_r_55, u0_key_r_6, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, 
        u0_u10_X_21, u0_u10_X_22, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, u0_u11_X_18, u0_u11_X_20, u0_u11_X_22, 
        u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, 
        u0_u12_X_2, u0_u12_X_24, u0_u12_X_37, u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, 
        u0_u12_X_46, u0_u12_X_48, u0_u12_X_5, u0_u12_X_7, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, u0_u13_X_48, 
        u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, u0_u14_X_18, u0_u14_X_19, u0_u14_X_20, 
        u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_42, u0_u1_X_25, 
        u0_u1_X_26, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, u0_u1_X_36, u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_40, 
        u0_u1_X_42, u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_3, u0_u2_X_9, u0_u5_X_10, u0_u5_X_15, u0_u5_X_16, 
        u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, u0_u5_X_9, u0_uk_K_r0_15, u0_uk_K_r0_28, 
        u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_7, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_41, u0_uk_K_r10_44, 
        u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, u0_uk_K_r11_33, u0_uk_K_r11_39, 
        u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_25, u0_uk_K_r14_15, u0_uk_K_r14_2, u0_uk_K_r14_50, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, 
        u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_33, u0_uk_K_r9_6, u0_uk_n100, 
        u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n101, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n109, 
        u0_uk_n115, u0_uk_n118, u0_uk_n121, u0_uk_n122, u0_uk_n126, u0_uk_n127, u0_uk_n128, u0_uk_n131, u0_uk_n139, 
        u0_uk_n143, u0_uk_n144, u0_uk_n146, u0_uk_n148, u0_uk_n153, u0_uk_n155, u0_uk_n161, u0_uk_n164, u0_uk_n172, 
        u0_uk_n173, u0_uk_n179, u0_uk_n180, u0_uk_n187, u0_uk_n188, u0_uk_n190, u0_uk_n191, u0_uk_n195, u0_uk_n196, 
        u0_uk_n197, u0_uk_n200, u0_uk_n201, u0_uk_n206, u0_uk_n212, u0_uk_n213, u0_uk_n214, u0_uk_n215, u0_uk_n221, 
        u0_uk_n225, u0_uk_n230, u0_uk_n240, u0_uk_n257, u0_uk_n410, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n414, 
        u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, u0_uk_n428, u0_uk_n429, 
        u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, u0_uk_n439, u0_uk_n440, u0_uk_n442, 
        u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n450, u0_uk_n547, u0_uk_n552, u0_uk_n557, u0_uk_n562, 
        u0_uk_n565, u0_uk_n568, u0_uk_n573, u0_uk_n578, u0_uk_n58, u0_uk_n63, u0_uk_n632, u0_uk_n643, u0_uk_n657, 
        u0_uk_n670, u0_uk_n674, u0_uk_n684, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, u0_uk_n786, u0_uk_n793, 
        u0_uk_n799, u0_uk_n8, u0_uk_n800, u0_uk_n83, u0_uk_n869, u0_uk_n892, u0_uk_n898, u0_uk_n91, u0_uk_n92, 
        u0_uk_n93, u0_uk_n94, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n976, u0_uk_n982, u0_uk_n99, 
        u0_uk_n999, u1_FP_40, u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, 
        u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, u1_K10_44, u1_K10_47, u1_K10_48, 
        u1_K11_11, u1_K11_13, u1_K11_2, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, u1_K11_7, 
        u1_K13_14, u1_K13_17, u1_K13_18, u1_K13_20, u1_K13_48, u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_42, 
        u1_K14_44, u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, u1_K15_2, 
        u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, u1_K15_36, 
        u1_K15_37, u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, u1_K16_13, 
        u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_20, u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_35, 
        u1_K1_1, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_20, u1_K2_23, u1_K2_24, u1_K2_25, 
        u1_K2_26, u1_K2_29, u1_K2_30, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, u1_K2_48, u1_K3_1, 
        u1_K3_2, u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, 
        u1_K3_5, u1_K3_6, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_6, u1_K5_19, u1_K5_23, u1_K5_24, 
        u1_K6_25, u1_K6_26, u1_K6_29, u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K7_1, 
        u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_2, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, 
        u1_K7_44, u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_7, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_29, 
        u1_K9_31, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, u1_K9_6, 
        u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, u1_R0_21, u1_R0_28, u1_R0_29, 
        u1_R0_32, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, 
        u1_R12_1, u1_R12_29, u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, 
        u1_R13_24, u1_R13_25, u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, 
        u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_32, u1_R1_4, u1_R1_5, u1_R2_1, u1_R2_2, 
        u1_R2_32, u1_R2_5, u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, 
        u1_R3_17, u1_R4_16, u1_R4_17, u1_R4_20, u1_R4_21, u1_R4_24, u1_R4_25, u1_R5_1, u1_R5_12, 
        u1_R5_13, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, u1_R5_32, u1_R5_4, u1_R5_5, 
        u1_R5_8, u1_R5_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_18, 
        u1_R7_20, u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, u1_R8_1, 
        u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R9_1, 
        u1_R9_12, u1_R9_20, u1_R9_21, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, 
        u1_desIn_r_25, u1_desIn_r_39, u1_desIn_r_57, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_2, u1_u0_X_3, u1_u0_X_31, 
        u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, 
        u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, u1_u0_X_48, u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, 
        u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, u1_u10_X_18, u1_u10_X_3, u1_u10_X_33, u1_u10_X_39, u1_u10_X_4, 
        u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, u1_u10_X_47, u1_u10_X_6, 
        u1_u10_X_8, u1_u10_X_9, u1_u12_X_1, u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, 
        u1_u12_X_3, u1_u12_X_4, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, u1_u12_X_9, u1_u13_X_10, 
        u1_u13_X_11, u1_u13_X_12, u1_u13_X_3, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, u1_u13_X_4, u1_u13_X_40, u1_u13_X_41, 
        u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, u1_u14_X_1, 
        u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, u1_u14_X_22, u1_u14_X_27, u1_u14_X_28, 
        u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, 
        u1_u14_X_9, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, u1_u15_X_22, u1_u15_X_23, u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, 
        u1_u15_X_27, u1_u15_X_28, u1_u15_X_33, u1_u15_X_36, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_37, 
        u1_u1_X_38, u1_u1_X_39, u1_u1_X_40, u1_u1_X_45, u1_u1_X_46, u1_u2_X_3, u1_u2_X_39, u1_u2_X_4, u1_u2_X_40, 
        u1_u2_X_45, u1_u2_X_46, u1_u3_X_4, u1_u3_X_5, u1_u3_X_7, u1_u3_X_9, u1_u4_X_21, u1_u5_X_27, u1_u5_X_28, 
        u1_u5_X_33, u1_u5_X_34, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_3, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, 
        u1_u6_X_45, u1_u6_X_9, u1_u8_X_21, u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, 
        u1_u8_X_39, u1_u8_X_4, u1_u8_X_40, u1_u8_X_45, u1_u8_X_46, u1_u9_X_34, u1_u9_X_39, u1_u9_X_40, u1_u9_X_45, 
        u1_u9_X_46, u1_uk_n1015, u1_uk_n1025, u1_uk_n1031, u1_uk_n1050, u1_uk_n1061, u1_uk_n1065, u1_uk_n1070, u1_uk_n1073, 
        u1_uk_n1074, u1_uk_n1105, u1_uk_n1106, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, u1_uk_n1126, u1_uk_n1154, u1_uk_n1155, 
        u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, u1_uk_n1166, u1_uk_n1167, u1_uk_n1170, 
        u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n437, u1_uk_n443, 
        u1_uk_n454, u1_uk_n496, u1_uk_n672, u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, 
        u1_uk_n949, u1_uk_n950, u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, 
        u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, u2_FP_48, u2_FP_49, 
        u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, u2_FP_64, u2_K11_11, 
        u2_K11_13, u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, u2_K16_19, 
        u2_K16_2, u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, u2_K16_32, 
        u2_K16_35, u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, u2_K16_5, 
        u2_K16_6, u2_K16_7, u2_K16_8, u2_K8_1, u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, 
        u2_K8_19, u2_K8_2, u2_K8_20, u2_K8_47, u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, 
        u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, 
        u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_22, u2_R7_24, u2_R7_25, 
        u2_R7_28, u2_R7_29, u2_R9_12, u2_R9_8, u2_R9_9, u2_u10_X_10, u2_u10_X_15, u2_u10_X_16, u2_u10_X_18, 
        u2_u10_X_7, u2_u10_X_8, u2_u10_X_9, u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, u2_u15_X_22, u2_u15_X_27, 
        u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, u2_u15_X_46, u2_u15_X_9, 
        u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, u2_u7_X_44, 
        u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, u2_u8_X_31, u2_u8_X_32, u2_u8_X_34, u2_u8_X_39, u2_u8_X_40, u2_u8_X_45, 
        u2_u8_X_46, u2_u8_X_47, u2_uk_K_r7_0, u2_uk_n1098, u2_uk_n1110, u2_uk_n1113, u2_uk_n1132, u2_uk_n1133, u2_uk_n1136, 
        u2_uk_n1137, u2_uk_n1140, u2_uk_n155, u2_uk_n1585, u2_uk_n214, u2_uk_n313, u2_uk_n319, u2_uk_n335, u2_uk_n955, 
        u2_uk_n958, u2_uk_n959, u2_uk_n963;
  output u0_out0_1, u0_out0_10, u0_out0_13, u0_out0_16, u0_out0_17, u0_out0_18, u0_out0_2, u0_out0_20, u0_out0_23, 
        u0_out0_24, u0_out0_26, u0_out0_28, u0_out0_30, u0_out0_31, u0_out0_6, u0_out0_9, u0_out10_1, u0_out10_10, 
        u0_out10_13, u0_out10_16, u0_out10_18, u0_out10_2, u0_out10_20, u0_out10_24, u0_out10_26, u0_out10_28, u0_out10_30, 
        u0_out10_6, u0_out11_1, u0_out11_10, u0_out11_11, u0_out11_12, u0_out11_16, u0_out11_19, u0_out11_20, u0_out11_22, 
        u0_out11_24, u0_out11_26, u0_out11_29, u0_out11_30, u0_out11_32, u0_out11_4, u0_out11_6, u0_out11_7, u0_out12_1, 
        u0_out12_10, u0_out12_12, u0_out12_13, u0_out12_15, u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_2, u0_out12_20, 
        u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_26, u0_out12_27, u0_out12_28, u0_out12_30, u0_out12_31, 
        u0_out12_32, u0_out12_5, u0_out12_6, u0_out12_7, u0_out12_9, u0_out13_15, u0_out13_21, u0_out13_27, u0_out13_5, 
        u0_out14_1, u0_out14_10, u0_out14_13, u0_out14_16, u0_out14_18, u0_out14_2, u0_out14_20, u0_out14_24, u0_out14_26, 
        u0_out14_28, u0_out14_30, u0_out14_6, u0_out15_12, u0_out15_22, u0_out15_32, u0_out15_7, u0_out1_11, u0_out1_12, 
        u0_out1_14, u0_out1_19, u0_out1_22, u0_out1_25, u0_out1_29, u0_out1_3, u0_out1_32, u0_out1_4, u0_out1_7, 
        u0_out1_8, u0_out2_13, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_2, u0_out2_23, u0_out2_24, u0_out2_28, 
        u0_out2_30, u0_out2_31, u0_out2_6, u0_out2_9, u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, u0_out5_13, 
        u0_out5_14, u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, u0_out5_21, 
        u0_out5_22, u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_3, 
        u0_out5_30, u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, u0_out5_9, 
        u0_uk_n10, u0_uk_n102, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, 
        u0_uk_n147, u0_uk_n162, u0_uk_n163, u0_uk_n182, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n217, 
        u0_uk_n220, u0_uk_n222, u0_uk_n231, u0_uk_n238, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n31, 
        u0_uk_n60, u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_15, u1_out0_17, u1_out0_18, u1_out0_19, u1_out0_2, 
        u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_27, u1_out0_28, u1_out0_29, u1_out0_31, u1_out0_32, u1_out0_4, 
        u1_out0_5, u1_out0_7, u1_out0_9, u1_out10_11, u1_out10_12, u1_out10_13, u1_out10_15, u1_out10_16, u1_out10_17, 
        u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_21, u1_out10_22, u1_out10_23, u1_out10_24, u1_out10_27, u1_out10_28, 
        u1_out10_29, u1_out10_30, u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_9, 
        u1_out12_1, u1_out12_10, u1_out12_13, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_2, u1_out12_20, 
        u1_out12_21, u1_out12_23, u1_out12_24, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_30, u1_out12_31, u1_out12_5, 
        u1_out12_6, u1_out12_9, u1_out13_12, u1_out13_13, u1_out13_15, u1_out13_17, u1_out13_18, u1_out13_2, u1_out13_21, 
        u1_out13_22, u1_out13_23, u1_out13_27, u1_out13_28, u1_out13_31, u1_out13_32, u1_out13_5, u1_out13_7, u1_out13_9, 
        u1_out14_1, u1_out14_10, u1_out14_11, u1_out14_12, u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, 
        u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_20, u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, 
        u1_out14_26, u1_out14_27, u1_out14_28, u1_out14_29, u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, 
        u1_out14_5, u1_out14_6, u1_out14_7, u1_out14_8, u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_14, 
        u1_out15_16, u1_out15_19, u1_out15_20, u1_out15_24, u1_out15_25, u1_out15_26, u1_out15_29, u1_out15_3, u1_out15_30, 
        u1_out15_4, u1_out15_6, u1_out15_8, u1_out1_1, u1_out1_10, u1_out1_12, u1_out1_14, u1_out1_15, u1_out1_20, 
        u1_out1_21, u1_out1_22, u1_out1_25, u1_out1_26, u1_out1_27, u1_out1_3, u1_out1_32, u1_out1_5, u1_out1_7, 
        u1_out1_8, u1_out2_12, u1_out2_15, u1_out2_17, u1_out2_21, u1_out2_22, u1_out2_23, u1_out2_27, u1_out2_31, 
        u1_out2_32, u1_out2_5, u1_out2_7, u1_out2_9, u1_out3_13, u1_out3_17, u1_out3_18, u1_out3_2, u1_out3_23, 
        u1_out3_28, u1_out3_31, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_20, u1_out4_26, u1_out5_11, u1_out5_14, 
        u1_out5_19, u1_out5_25, u1_out5_29, u1_out5_3, u1_out5_4, u1_out5_8, u1_out6_12, u1_out6_13, u1_out6_15, 
        u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_2, u1_out6_21, u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_27, 
        u1_out6_28, u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_9, u1_out8_1, 
        u1_out8_10, u1_out8_11, u1_out8_12, u1_out8_14, u1_out8_15, u1_out8_17, u1_out8_19, u1_out8_20, u1_out8_21, 
        u1_out8_22, u1_out8_23, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_29, u1_out8_3, u1_out8_31, u1_out8_32, 
        u1_out8_4, u1_out8_5, u1_out8_7, u1_out8_8, u1_out8_9, u1_out9_11, u1_out9_12, u1_out9_15, u1_out9_19, 
        u1_out9_21, u1_out9_22, u1_out9_27, u1_out9_29, u1_out9_32, u1_out9_4, u1_out9_5, u1_out9_7, u2_out10_13, 
        u2_out10_16, u2_out10_18, u2_out10_2, u2_out10_24, u2_out10_28, u2_out10_30, u2_out10_6, u2_out15_1, u2_out15_10, 
        u2_out15_11, u2_out15_12, u2_out15_13, u2_out15_14, u2_out15_15, u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_19, 
        u2_out15_2, u2_out15_20, u2_out15_21, u2_out15_22, u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_27, 
        u2_out15_28, u2_out15_29, u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_6, 
        u2_out15_7, u2_out15_8, u2_out15_9, u2_out7_1, u2_out7_10, u2_out7_13, u2_out7_15, u2_out7_16, u2_out7_17, 
        u2_out7_18, u2_out7_2, u2_out7_20, u2_out7_21, u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_27, u2_out7_28, 
        u2_out7_30, u2_out7_31, u2_out7_5, u2_out7_6, u2_out7_9, u2_out8_11, u2_out8_12, u2_out8_15, u2_out8_19, 
        u2_out8_21, u2_out8_22, u2_out8_27, u2_out8_29, u2_out8_32, u2_out8_4, u2_out8_5, u2_out8_7;
  wire u0_K11_10, u0_K11_11, u0_K11_12, u0_K11_13, u0_K11_14, u0_K11_15, u0_K11_16, u0_K11_17, u0_K11_18, 
       u0_K11_19, u0_K11_20, u0_K11_23, u0_K11_24, u0_K11_7, u0_K11_8, u0_K11_9, u0_K12_17, u0_K12_21, 
       u0_K12_23, u0_K12_24, u0_K12_31, u0_K12_32, u0_K12_37, u0_K12_38, u0_K12_41, u0_K12_42, u0_K13_1, 
       u0_K13_15, u0_K13_16, u0_K13_17, u0_K13_18, u0_K13_19, u0_K13_20, u0_K13_21, u0_K13_22, u0_K13_23, 
       u0_K13_3, u0_K13_4, u0_K13_43, u0_K13_47, u0_K13_6, u0_K13_8, u0_K13_9, u0_K14_45, u0_K15_11, 
       u0_K16_37, u0_K16_39, u0_K16_40, u0_K16_41, u0_K1_1, u0_K1_10, u0_K1_11, u0_K1_12, u0_K1_18, 
       u0_K1_19, u0_K1_2, u0_K1_20, u0_K1_24, u0_K1_3, u0_K1_4, u0_K1_5, u0_K1_6, u0_K1_7, 
       u0_K1_8, u0_K1_9, u0_K2_27, u0_K2_28, u0_K2_32, u0_K2_41, u0_K3_1, u0_K3_11, u0_K3_2, 
       u0_K3_4, u0_K3_7, u0_K3_8, u0_K6_1, u0_K6_12, u0_K6_14, u0_K6_17, u0_K6_18, u0_K6_2, 
       u0_K6_25, u0_K6_26, u0_K6_28, u0_K6_29, u0_K6_30, u0_K6_31, u0_K6_32, u0_K6_33, u0_K6_35, 
       u0_K6_36, u0_K6_37, u0_K6_38, u0_K6_39, u0_K6_4, u0_K6_40, u0_K6_42, u0_K6_43, u0_K6_44, 
       u0_K6_45, u0_K6_47, u0_K6_48, u0_K6_5, u0_K6_6, u0_K6_7, u0_K6_8, u0_u0_X_1, u0_u0_X_10, 
       u0_u0_X_11, u0_u0_X_12, u0_u0_X_13, u0_u0_X_14, u0_u0_X_17, u0_u0_X_18, u0_u0_X_19, u0_u0_X_2, u0_u0_X_20, 
       u0_u0_X_24, u0_u0_X_3, u0_u0_X_4, u0_u0_X_5, u0_u0_X_6, u0_u0_X_7, u0_u0_X_8, u0_u0_X_9, u0_u0_u0_n1, 
       u0_u0_u0_n10, u0_u0_u0_n11, u0_u0_u0_n12, u0_u0_u0_n13, u0_u0_u0_n14, u0_u0_u0_n15, u0_u0_u0_n16, u0_u0_u0_n17, u0_u0_u0_n18, 
       u0_u0_u0_n19, u0_u0_u0_n2, u0_u0_u0_n20, u0_u0_u0_n21, u0_u0_u0_n22, u0_u0_u0_n23, u0_u0_u0_n24, u0_u0_u0_n25, u0_u0_u0_n26, 
       u0_u0_u0_n27, u0_u0_u0_n28, u0_u0_u0_n29, u0_u0_u0_n3, u0_u0_u0_n30, u0_u0_u0_n31, u0_u0_u0_n32, u0_u0_u0_n33, u0_u0_u0_n34, 
       u0_u0_u0_n35, u0_u0_u0_n36, u0_u0_u0_n37, u0_u0_u0_n38, u0_u0_u0_n39, u0_u0_u0_n4, u0_u0_u0_n40, u0_u0_u0_n41, u0_u0_u0_n42, 
       u0_u0_u0_n43, u0_u0_u0_n44, u0_u0_u0_n45, u0_u0_u0_n46, u0_u0_u0_n47, u0_u0_u0_n48, u0_u0_u0_n49, u0_u0_u0_n5, u0_u0_u0_n50, 
       u0_u0_u0_n51, u0_u0_u0_n52, u0_u0_u0_n53, u0_u0_u0_n54, u0_u0_u0_n55, u0_u0_u0_n56, u0_u0_u0_n57, u0_u0_u0_n58, u0_u0_u0_n59, 
       u0_u0_u0_n6, u0_u0_u0_n60, u0_u0_u0_n61, u0_u0_u0_n62, u0_u0_u0_n63, u0_u0_u0_n64, u0_u0_u0_n65, u0_u0_u0_n66, u0_u0_u0_n67, 
       u0_u0_u0_n68, u0_u0_u0_n69, u0_u0_u0_n7, u0_u0_u0_n70, u0_u0_u0_n71, u0_u0_u0_n72, u0_u0_u0_n73, u0_u0_u0_n74, u0_u0_u0_n75, 
       u0_u0_u0_n76, u0_u0_u0_n77, u0_u0_u0_n78, u0_u0_u0_n79, u0_u0_u0_n8, u0_u0_u0_n80, u0_u0_u0_n81, u0_u0_u0_n82, u0_u0_u0_n83, 
       u0_u0_u0_n84, u0_u0_u0_n85, u0_u0_u0_n86, u0_u0_u0_n87, u0_u0_u0_n9, u0_u0_u1_n1, u0_u0_u1_n10, u0_u0_u1_n11, u0_u0_u1_n12, 
       u0_u0_u1_n13, u0_u0_u1_n14, u0_u0_u1_n15, u0_u0_u1_n16, u0_u0_u1_n17, u0_u0_u1_n18, u0_u0_u1_n19, u0_u0_u1_n2, u0_u0_u1_n20, 
       u0_u0_u1_n21, u0_u0_u1_n22, u0_u0_u1_n23, u0_u0_u1_n24, u0_u0_u1_n25, u0_u0_u1_n26, u0_u0_u1_n27, u0_u0_u1_n28, u0_u0_u1_n29, 
       u0_u0_u1_n3, u0_u0_u1_n30, u0_u0_u1_n31, u0_u0_u1_n32, u0_u0_u1_n33, u0_u0_u1_n34, u0_u0_u1_n35, u0_u0_u1_n36, u0_u0_u1_n37, 
       u0_u0_u1_n38, u0_u0_u1_n39, u0_u0_u1_n4, u0_u0_u1_n40, u0_u0_u1_n41, u0_u0_u1_n42, u0_u0_u1_n43, u0_u0_u1_n44, u0_u0_u1_n45, 
       u0_u0_u1_n46, u0_u0_u1_n47, u0_u0_u1_n48, u0_u0_u1_n49, u0_u0_u1_n5, u0_u0_u1_n50, u0_u0_u1_n51, u0_u0_u1_n52, u0_u0_u1_n53, 
       u0_u0_u1_n54, u0_u0_u1_n55, u0_u0_u1_n56, u0_u0_u1_n57, u0_u0_u1_n58, u0_u0_u1_n59, u0_u0_u1_n6, u0_u0_u1_n60, u0_u0_u1_n61, 
       u0_u0_u1_n62, u0_u0_u1_n63, u0_u0_u1_n64, u0_u0_u1_n65, u0_u0_u1_n66, u0_u0_u1_n67, u0_u0_u1_n68, u0_u0_u1_n69, u0_u0_u1_n7, 
       u0_u0_u1_n70, u0_u0_u1_n71, u0_u0_u1_n72, u0_u0_u1_n73, u0_u0_u1_n74, u0_u0_u1_n75, u0_u0_u1_n76, u0_u0_u1_n77, u0_u0_u1_n78, 
       u0_u0_u1_n79, u0_u0_u1_n8, u0_u0_u1_n80, u0_u0_u1_n81, u0_u0_u1_n82, u0_u0_u1_n83, u0_u0_u1_n84, u0_u0_u1_n85, u0_u0_u1_n86, 
       u0_u0_u1_n87, u0_u0_u1_n88, u0_u0_u1_n89, u0_u0_u1_n9, u0_u0_u1_n90, u0_u0_u1_n91, u0_u0_u1_n92, u0_u0_u1_n93, u0_u0_u1_n94, 
       u0_u0_u2_n1, u0_u0_u2_n10, u0_u0_u2_n11, u0_u0_u2_n12, u0_u0_u2_n13, u0_u0_u2_n14, u0_u0_u2_n15, u0_u0_u2_n16, u0_u0_u2_n17, 
       u0_u0_u2_n18, u0_u0_u2_n19, u0_u0_u2_n2, u0_u0_u2_n20, u0_u0_u2_n21, u0_u0_u2_n22, u0_u0_u2_n23, u0_u0_u2_n24, u0_u0_u2_n25, 
       u0_u0_u2_n26, u0_u0_u2_n27, u0_u0_u2_n28, u0_u0_u2_n29, u0_u0_u2_n3, u0_u0_u2_n30, u0_u0_u2_n31, u0_u0_u2_n32, u0_u0_u2_n33, 
       u0_u0_u2_n34, u0_u0_u2_n35, u0_u0_u2_n36, u0_u0_u2_n37, u0_u0_u2_n38, u0_u0_u2_n39, u0_u0_u2_n4, u0_u0_u2_n40, u0_u0_u2_n41, 
       u0_u0_u2_n42, u0_u0_u2_n43, u0_u0_u2_n44, u0_u0_u2_n45, u0_u0_u2_n46, u0_u0_u2_n47, u0_u0_u2_n48, u0_u0_u2_n49, u0_u0_u2_n5, 
       u0_u0_u2_n50, u0_u0_u2_n51, u0_u0_u2_n52, u0_u0_u2_n53, u0_u0_u2_n54, u0_u0_u2_n55, u0_u0_u2_n56, u0_u0_u2_n57, u0_u0_u2_n58, 
       u0_u0_u2_n59, u0_u0_u2_n6, u0_u0_u2_n60, u0_u0_u2_n61, u0_u0_u2_n62, u0_u0_u2_n63, u0_u0_u2_n64, u0_u0_u2_n65, u0_u0_u2_n66, 
       u0_u0_u2_n67, u0_u0_u2_n68, u0_u0_u2_n69, u0_u0_u2_n7, u0_u0_u2_n70, u0_u0_u2_n71, u0_u0_u2_n72, u0_u0_u2_n73, u0_u0_u2_n74, 
       u0_u0_u2_n75, u0_u0_u2_n76, u0_u0_u2_n77, u0_u0_u2_n78, u0_u0_u2_n79, u0_u0_u2_n8, u0_u0_u2_n80, u0_u0_u2_n81, u0_u0_u2_n82, 
       u0_u0_u2_n83, u0_u0_u2_n84, u0_u0_u2_n85, u0_u0_u2_n86, u0_u0_u2_n87, u0_u0_u2_n88, u0_u0_u2_n89, u0_u0_u2_n9, u0_u0_u2_n90, 
       u0_u0_u2_n91, u0_u0_u2_n92, u0_u0_u2_n93, u0_u0_u2_n94, u0_u0_u3_n1, u0_u0_u3_n10, u0_u0_u3_n11, u0_u0_u3_n12, u0_u0_u3_n13, 
       u0_u0_u3_n14, u0_u0_u3_n15, u0_u0_u3_n16, u0_u0_u3_n17, u0_u0_u3_n18, u0_u0_u3_n19, u0_u0_u3_n2, u0_u0_u3_n20, u0_u0_u3_n21, 
       u0_u0_u3_n22, u0_u0_u3_n23, u0_u0_u3_n24, u0_u0_u3_n25, u0_u0_u3_n26, u0_u0_u3_n27, u0_u0_u3_n28, u0_u0_u3_n29, u0_u0_u3_n3, 
       u0_u0_u3_n30, u0_u0_u3_n31, u0_u0_u3_n32, u0_u0_u3_n33, u0_u0_u3_n34, u0_u0_u3_n35, u0_u0_u3_n36, u0_u0_u3_n37, u0_u0_u3_n38, 
       u0_u0_u3_n39, u0_u0_u3_n4, u0_u0_u3_n40, u0_u0_u3_n41, u0_u0_u3_n42, u0_u0_u3_n43, u0_u0_u3_n44, u0_u0_u3_n45, u0_u0_u3_n46, 
       u0_u0_u3_n47, u0_u0_u3_n48, u0_u0_u3_n49, u0_u0_u3_n5, u0_u0_u3_n50, u0_u0_u3_n51, u0_u0_u3_n52, u0_u0_u3_n53, u0_u0_u3_n54, 
       u0_u0_u3_n55, u0_u0_u3_n56, u0_u0_u3_n57, u0_u0_u3_n58, u0_u0_u3_n59, u0_u0_u3_n6, u0_u0_u3_n60, u0_u0_u3_n61, u0_u0_u3_n62, 
       u0_u0_u3_n63, u0_u0_u3_n64, u0_u0_u3_n65, u0_u0_u3_n66, u0_u0_u3_n67, u0_u0_u3_n68, u0_u0_u3_n69, u0_u0_u3_n7, u0_u0_u3_n70, 
       u0_u0_u3_n71, u0_u0_u3_n72, u0_u0_u3_n73, u0_u0_u3_n74, u0_u0_u3_n75, u0_u0_u3_n76, u0_u0_u3_n77, u0_u0_u3_n78, u0_u0_u3_n79, 
       u0_u0_u3_n8, u0_u0_u3_n80, u0_u0_u3_n81, u0_u0_u3_n82, u0_u0_u3_n83, u0_u0_u3_n84, u0_u0_u3_n85, u0_u0_u3_n86, u0_u0_u3_n87, 
       u0_u0_u3_n88, u0_u0_u3_n89, u0_u0_u3_n9, u0_u0_u3_n90, u0_u0_u3_n91, u0_u0_u3_n92, u0_u0_u3_n93, u0_u10_X_10, u0_u10_X_11, 
       u0_u10_X_12, u0_u10_X_13, u0_u10_X_14, u0_u10_X_15, u0_u10_X_16, u0_u10_X_17, u0_u10_X_18, u0_u10_X_19, u0_u10_X_20, 
       u0_u10_X_23, u0_u10_X_24, u0_u10_X_7, u0_u10_X_8, u0_u10_X_9, u0_u10_u1_n100, u0_u10_u1_n101, u0_u10_u1_n102, u0_u10_u1_n103, 
       u0_u10_u1_n104, u0_u10_u1_n105, u0_u10_u1_n106, u0_u10_u1_n107, u0_u10_u1_n108, u0_u10_u1_n109, u0_u10_u1_n110, u0_u10_u1_n111, u0_u10_u1_n112, 
       u0_u10_u1_n113, u0_u10_u1_n114, u0_u10_u1_n115, u0_u10_u1_n116, u0_u10_u1_n117, u0_u10_u1_n118, u0_u10_u1_n119, u0_u10_u1_n120, u0_u10_u1_n121, 
       u0_u10_u1_n122, u0_u10_u1_n123, u0_u10_u1_n124, u0_u10_u1_n125, u0_u10_u1_n126, u0_u10_u1_n127, u0_u10_u1_n128, u0_u10_u1_n129, u0_u10_u1_n130, 
       u0_u10_u1_n131, u0_u10_u1_n132, u0_u10_u1_n133, u0_u10_u1_n134, u0_u10_u1_n135, u0_u10_u1_n136, u0_u10_u1_n137, u0_u10_u1_n138, u0_u10_u1_n139, 
       u0_u10_u1_n140, u0_u10_u1_n141, u0_u10_u1_n142, u0_u10_u1_n143, u0_u10_u1_n144, u0_u10_u1_n145, u0_u10_u1_n146, u0_u10_u1_n147, u0_u10_u1_n148, 
       u0_u10_u1_n149, u0_u10_u1_n150, u0_u10_u1_n151, u0_u10_u1_n152, u0_u10_u1_n153, u0_u10_u1_n154, u0_u10_u1_n155, u0_u10_u1_n156, u0_u10_u1_n157, 
       u0_u10_u1_n158, u0_u10_u1_n159, u0_u10_u1_n160, u0_u10_u1_n161, u0_u10_u1_n162, u0_u10_u1_n163, u0_u10_u1_n164, u0_u10_u1_n165, u0_u10_u1_n166, 
       u0_u10_u1_n167, u0_u10_u1_n168, u0_u10_u1_n169, u0_u10_u1_n170, u0_u10_u1_n171, u0_u10_u1_n172, u0_u10_u1_n173, u0_u10_u1_n174, u0_u10_u1_n175, 
       u0_u10_u1_n176, u0_u10_u1_n177, u0_u10_u1_n178, u0_u10_u1_n179, u0_u10_u1_n180, u0_u10_u1_n181, u0_u10_u1_n182, u0_u10_u1_n183, u0_u10_u1_n184, 
       u0_u10_u1_n185, u0_u10_u1_n186, u0_u10_u1_n187, u0_u10_u1_n188, u0_u10_u1_n95, u0_u10_u1_n96, u0_u10_u1_n97, u0_u10_u1_n98, u0_u10_u1_n99, 
       u0_u10_u2_n100, u0_u10_u2_n101, u0_u10_u2_n102, u0_u10_u2_n103, u0_u10_u2_n104, u0_u10_u2_n105, u0_u10_u2_n106, u0_u10_u2_n107, u0_u10_u2_n108, 
       u0_u10_u2_n109, u0_u10_u2_n110, u0_u10_u2_n111, u0_u10_u2_n112, u0_u10_u2_n113, u0_u10_u2_n114, u0_u10_u2_n115, u0_u10_u2_n116, u0_u10_u2_n117, 
       u0_u10_u2_n118, u0_u10_u2_n119, u0_u10_u2_n120, u0_u10_u2_n121, u0_u10_u2_n122, u0_u10_u2_n123, u0_u10_u2_n124, u0_u10_u2_n125, u0_u10_u2_n126, 
       u0_u10_u2_n127, u0_u10_u2_n128, u0_u10_u2_n129, u0_u10_u2_n130, u0_u10_u2_n131, u0_u10_u2_n132, u0_u10_u2_n133, u0_u10_u2_n134, u0_u10_u2_n135, 
       u0_u10_u2_n136, u0_u10_u2_n137, u0_u10_u2_n138, u0_u10_u2_n139, u0_u10_u2_n140, u0_u10_u2_n141, u0_u10_u2_n142, u0_u10_u2_n143, u0_u10_u2_n144, 
       u0_u10_u2_n145, u0_u10_u2_n146, u0_u10_u2_n147, u0_u10_u2_n148, u0_u10_u2_n149, u0_u10_u2_n150, u0_u10_u2_n151, u0_u10_u2_n152, u0_u10_u2_n153, 
       u0_u10_u2_n154, u0_u10_u2_n155, u0_u10_u2_n156, u0_u10_u2_n157, u0_u10_u2_n158, u0_u10_u2_n159, u0_u10_u2_n160, u0_u10_u2_n161, u0_u10_u2_n162, 
       u0_u10_u2_n163, u0_u10_u2_n164, u0_u10_u2_n165, u0_u10_u2_n166, u0_u10_u2_n167, u0_u10_u2_n168, u0_u10_u2_n169, u0_u10_u2_n170, u0_u10_u2_n171, 
       u0_u10_u2_n172, u0_u10_u2_n173, u0_u10_u2_n174, u0_u10_u2_n175, u0_u10_u2_n176, u0_u10_u2_n177, u0_u10_u2_n178, u0_u10_u2_n179, u0_u10_u2_n180, 
       u0_u10_u2_n181, u0_u10_u2_n182, u0_u10_u2_n183, u0_u10_u2_n184, u0_u10_u2_n185, u0_u10_u2_n186, u0_u10_u2_n187, u0_u10_u2_n188, u0_u10_u2_n95, 
       u0_u10_u2_n96, u0_u10_u2_n97, u0_u10_u2_n98, u0_u10_u2_n99, u0_u10_u3_n100, u0_u10_u3_n101, u0_u10_u3_n102, u0_u10_u3_n103, u0_u10_u3_n104, 
       u0_u10_u3_n105, u0_u10_u3_n106, u0_u10_u3_n107, u0_u10_u3_n108, u0_u10_u3_n109, u0_u10_u3_n110, u0_u10_u3_n111, u0_u10_u3_n112, u0_u10_u3_n113, 
       u0_u10_u3_n114, u0_u10_u3_n115, u0_u10_u3_n116, u0_u10_u3_n117, u0_u10_u3_n118, u0_u10_u3_n119, u0_u10_u3_n120, u0_u10_u3_n121, u0_u10_u3_n122, 
       u0_u10_u3_n123, u0_u10_u3_n124, u0_u10_u3_n125, u0_u10_u3_n126, u0_u10_u3_n127, u0_u10_u3_n128, u0_u10_u3_n129, u0_u10_u3_n130, u0_u10_u3_n131, 
       u0_u10_u3_n132, u0_u10_u3_n133, u0_u10_u3_n134, u0_u10_u3_n135, u0_u10_u3_n136, u0_u10_u3_n137, u0_u10_u3_n138, u0_u10_u3_n139, u0_u10_u3_n140, 
       u0_u10_u3_n141, u0_u10_u3_n142, u0_u10_u3_n143, u0_u10_u3_n144, u0_u10_u3_n145, u0_u10_u3_n146, u0_u10_u3_n147, u0_u10_u3_n148, u0_u10_u3_n149, 
       u0_u10_u3_n150, u0_u10_u3_n151, u0_u10_u3_n152, u0_u10_u3_n153, u0_u10_u3_n154, u0_u10_u3_n155, u0_u10_u3_n156, u0_u10_u3_n157, u0_u10_u3_n158, 
       u0_u10_u3_n159, u0_u10_u3_n160, u0_u10_u3_n161, u0_u10_u3_n162, u0_u10_u3_n163, u0_u10_u3_n164, u0_u10_u3_n165, u0_u10_u3_n166, u0_u10_u3_n167, 
       u0_u10_u3_n168, u0_u10_u3_n169, u0_u10_u3_n170, u0_u10_u3_n171, u0_u10_u3_n172, u0_u10_u3_n173, u0_u10_u3_n174, u0_u10_u3_n175, u0_u10_u3_n176, 
       u0_u10_u3_n177, u0_u10_u3_n178, u0_u10_u3_n179, u0_u10_u3_n180, u0_u10_u3_n181, u0_u10_u3_n182, u0_u10_u3_n183, u0_u10_u3_n184, u0_u10_u3_n185, 
       u0_u10_u3_n186, u0_u10_u3_n94, u0_u10_u3_n95, u0_u10_u3_n96, u0_u10_u3_n97, u0_u10_u3_n98, u0_u10_u3_n99, u0_u11_X_17, u0_u11_X_19, 
       u0_u11_X_21, u0_u11_X_23, u0_u11_X_24, u0_u11_X_31, u0_u11_X_32, u0_u11_X_35, u0_u11_X_36, u0_u11_X_37, u0_u11_X_38, 
       u0_u11_X_41, u0_u11_X_42, u0_u11_u2_n100, u0_u11_u2_n101, u0_u11_u2_n102, u0_u11_u2_n103, u0_u11_u2_n104, u0_u11_u2_n105, u0_u11_u2_n106, 
       u0_u11_u2_n107, u0_u11_u2_n108, u0_u11_u2_n109, u0_u11_u2_n110, u0_u11_u2_n111, u0_u11_u2_n112, u0_u11_u2_n113, u0_u11_u2_n114, u0_u11_u2_n115, 
       u0_u11_u2_n116, u0_u11_u2_n117, u0_u11_u2_n118, u0_u11_u2_n119, u0_u11_u2_n120, u0_u11_u2_n121, u0_u11_u2_n122, u0_u11_u2_n123, u0_u11_u2_n124, 
       u0_u11_u2_n125, u0_u11_u2_n126, u0_u11_u2_n127, u0_u11_u2_n128, u0_u11_u2_n129, u0_u11_u2_n130, u0_u11_u2_n131, u0_u11_u2_n132, u0_u11_u2_n133, 
       u0_u11_u2_n134, u0_u11_u2_n135, u0_u11_u2_n136, u0_u11_u2_n137, u0_u11_u2_n138, u0_u11_u2_n139, u0_u11_u2_n140, u0_u11_u2_n141, u0_u11_u2_n142, 
       u0_u11_u2_n143, u0_u11_u2_n144, u0_u11_u2_n145, u0_u11_u2_n146, u0_u11_u2_n147, u0_u11_u2_n148, u0_u11_u2_n149, u0_u11_u2_n150, u0_u11_u2_n151, 
       u0_u11_u2_n152, u0_u11_u2_n153, u0_u11_u2_n154, u0_u11_u2_n155, u0_u11_u2_n156, u0_u11_u2_n157, u0_u11_u2_n158, u0_u11_u2_n159, u0_u11_u2_n160, 
       u0_u11_u2_n161, u0_u11_u2_n162, u0_u11_u2_n163, u0_u11_u2_n164, u0_u11_u2_n165, u0_u11_u2_n166, u0_u11_u2_n167, u0_u11_u2_n168, u0_u11_u2_n169, 
       u0_u11_u2_n170, u0_u11_u2_n171, u0_u11_u2_n172, u0_u11_u2_n173, u0_u11_u2_n174, u0_u11_u2_n175, u0_u11_u2_n176, u0_u11_u2_n177, u0_u11_u2_n178, 
       u0_u11_u2_n179, u0_u11_u2_n180, u0_u11_u2_n181, u0_u11_u2_n182, u0_u11_u2_n183, u0_u11_u2_n184, u0_u11_u2_n185, u0_u11_u2_n186, u0_u11_u2_n187, 
       u0_u11_u2_n188, u0_u11_u2_n95, u0_u11_u2_n96, u0_u11_u2_n97, u0_u11_u2_n98, u0_u11_u2_n99, u0_u11_u3_n100, u0_u11_u3_n101, u0_u11_u3_n102, 
       u0_u11_u3_n103, u0_u11_u3_n104, u0_u11_u3_n105, u0_u11_u3_n106, u0_u11_u3_n107, u0_u11_u3_n108, u0_u11_u3_n109, u0_u11_u3_n110, u0_u11_u3_n111, 
       u0_u11_u3_n112, u0_u11_u3_n113, u0_u11_u3_n114, u0_u11_u3_n115, u0_u11_u3_n116, u0_u11_u3_n117, u0_u11_u3_n118, u0_u11_u3_n119, u0_u11_u3_n120, 
       u0_u11_u3_n121, u0_u11_u3_n122, u0_u11_u3_n123, u0_u11_u3_n124, u0_u11_u3_n125, u0_u11_u3_n126, u0_u11_u3_n127, u0_u11_u3_n128, u0_u11_u3_n129, 
       u0_u11_u3_n130, u0_u11_u3_n131, u0_u11_u3_n132, u0_u11_u3_n133, u0_u11_u3_n134, u0_u11_u3_n135, u0_u11_u3_n136, u0_u11_u3_n137, u0_u11_u3_n138, 
       u0_u11_u3_n139, u0_u11_u3_n140, u0_u11_u3_n141, u0_u11_u3_n142, u0_u11_u3_n143, u0_u11_u3_n144, u0_u11_u3_n145, u0_u11_u3_n146, u0_u11_u3_n147, 
       u0_u11_u3_n148, u0_u11_u3_n149, u0_u11_u3_n150, u0_u11_u3_n151, u0_u11_u3_n152, u0_u11_u3_n153, u0_u11_u3_n154, u0_u11_u3_n155, u0_u11_u3_n156, 
       u0_u11_u3_n157, u0_u11_u3_n158, u0_u11_u3_n159, u0_u11_u3_n160, u0_u11_u3_n161, u0_u11_u3_n162, u0_u11_u3_n163, u0_u11_u3_n164, u0_u11_u3_n165, 
       u0_u11_u3_n166, u0_u11_u3_n167, u0_u11_u3_n168, u0_u11_u3_n169, u0_u11_u3_n170, u0_u11_u3_n171, u0_u11_u3_n172, u0_u11_u3_n173, u0_u11_u3_n174, 
       u0_u11_u3_n175, u0_u11_u3_n176, u0_u11_u3_n177, u0_u11_u3_n178, u0_u11_u3_n179, u0_u11_u3_n180, u0_u11_u3_n181, u0_u11_u3_n182, u0_u11_u3_n183, 
       u0_u11_u3_n184, u0_u11_u3_n185, u0_u11_u3_n186, u0_u11_u3_n94, u0_u11_u3_n95, u0_u11_u3_n96, u0_u11_u3_n97, u0_u11_u3_n98, u0_u11_u3_n99, 
       u0_u11_u5_n100, u0_u11_u5_n101, u0_u11_u5_n102, u0_u11_u5_n103, u0_u11_u5_n104, u0_u11_u5_n105, u0_u11_u5_n106, u0_u11_u5_n107, u0_u11_u5_n108, 
       u0_u11_u5_n109, u0_u11_u5_n110, u0_u11_u5_n111, u0_u11_u5_n112, u0_u11_u5_n113, u0_u11_u5_n114, u0_u11_u5_n115, u0_u11_u5_n116, u0_u11_u5_n117, 
       u0_u11_u5_n118, u0_u11_u5_n119, u0_u11_u5_n120, u0_u11_u5_n121, u0_u11_u5_n122, u0_u11_u5_n123, u0_u11_u5_n124, u0_u11_u5_n125, u0_u11_u5_n126, 
       u0_u11_u5_n127, u0_u11_u5_n128, u0_u11_u5_n129, u0_u11_u5_n130, u0_u11_u5_n131, u0_u11_u5_n132, u0_u11_u5_n133, u0_u11_u5_n134, u0_u11_u5_n135, 
       u0_u11_u5_n136, u0_u11_u5_n137, u0_u11_u5_n138, u0_u11_u5_n139, u0_u11_u5_n140, u0_u11_u5_n141, u0_u11_u5_n142, u0_u11_u5_n143, u0_u11_u5_n144, 
       u0_u11_u5_n145, u0_u11_u5_n146, u0_u11_u5_n147, u0_u11_u5_n148, u0_u11_u5_n149, u0_u11_u5_n150, u0_u11_u5_n151, u0_u11_u5_n152, u0_u11_u5_n153, 
       u0_u11_u5_n154, u0_u11_u5_n155, u0_u11_u5_n156, u0_u11_u5_n157, u0_u11_u5_n158, u0_u11_u5_n159, u0_u11_u5_n160, u0_u11_u5_n161, u0_u11_u5_n162, 
       u0_u11_u5_n163, u0_u11_u5_n164, u0_u11_u5_n165, u0_u11_u5_n166, u0_u11_u5_n167, u0_u11_u5_n168, u0_u11_u5_n169, u0_u11_u5_n170, u0_u11_u5_n171, 
       u0_u11_u5_n172, u0_u11_u5_n173, u0_u11_u5_n174, u0_u11_u5_n175, u0_u11_u5_n176, u0_u11_u5_n177, u0_u11_u5_n178, u0_u11_u5_n179, u0_u11_u5_n180, 
       u0_u11_u5_n181, u0_u11_u5_n182, u0_u11_u5_n183, u0_u11_u5_n184, u0_u11_u5_n185, u0_u11_u5_n186, u0_u11_u5_n187, u0_u11_u5_n188, u0_u11_u5_n189, 
       u0_u11_u5_n190, u0_u11_u5_n191, u0_u11_u5_n192, u0_u11_u5_n193, u0_u11_u5_n194, u0_u11_u5_n195, u0_u11_u5_n196, u0_u11_u5_n99, u0_u11_u6_n100, 
       u0_u11_u6_n101, u0_u11_u6_n102, u0_u11_u6_n103, u0_u11_u6_n104, u0_u11_u6_n105, u0_u11_u6_n106, u0_u11_u6_n107, u0_u11_u6_n108, u0_u11_u6_n109, 
       u0_u11_u6_n110, u0_u11_u6_n111, u0_u11_u6_n112, u0_u11_u6_n113, u0_u11_u6_n114, u0_u11_u6_n115, u0_u11_u6_n116, u0_u11_u6_n117, u0_u11_u6_n118, 
       u0_u11_u6_n119, u0_u11_u6_n120, u0_u11_u6_n121, u0_u11_u6_n122, u0_u11_u6_n123, u0_u11_u6_n124, u0_u11_u6_n125, u0_u11_u6_n126, u0_u11_u6_n127, 
       u0_u11_u6_n128, u0_u11_u6_n129, u0_u11_u6_n130, u0_u11_u6_n131, u0_u11_u6_n132, u0_u11_u6_n133, u0_u11_u6_n134, u0_u11_u6_n135, u0_u11_u6_n136, 
       u0_u11_u6_n137, u0_u11_u6_n138, u0_u11_u6_n139, u0_u11_u6_n140, u0_u11_u6_n141, u0_u11_u6_n142, u0_u11_u6_n143, u0_u11_u6_n144, u0_u11_u6_n145, 
       u0_u11_u6_n146, u0_u11_u6_n147, u0_u11_u6_n148, u0_u11_u6_n149, u0_u11_u6_n150, u0_u11_u6_n151, u0_u11_u6_n152, u0_u11_u6_n153, u0_u11_u6_n154, 
       u0_u11_u6_n155, u0_u11_u6_n156, u0_u11_u6_n157, u0_u11_u6_n158, u0_u11_u6_n159, u0_u11_u6_n160, u0_u11_u6_n161, u0_u11_u6_n162, u0_u11_u6_n163, 
       u0_u11_u6_n164, u0_u11_u6_n165, u0_u11_u6_n166, u0_u11_u6_n167, u0_u11_u6_n168, u0_u11_u6_n169, u0_u11_u6_n170, u0_u11_u6_n171, u0_u11_u6_n172, 
       u0_u11_u6_n173, u0_u11_u6_n174, u0_u11_u6_n88, u0_u11_u6_n89, u0_u11_u6_n90, u0_u11_u6_n91, u0_u11_u6_n92, u0_u11_u6_n93, u0_u11_u6_n94, 
       u0_u11_u6_n95, u0_u11_u6_n96, u0_u11_u6_n97, u0_u11_u6_n98, u0_u11_u6_n99, u0_u12_X_1, u0_u12_X_15, u0_u12_X_16, u0_u12_X_17, 
       u0_u12_X_18, u0_u12_X_19, u0_u12_X_20, u0_u12_X_21, u0_u12_X_22, u0_u12_X_23, u0_u12_X_3, u0_u12_X_4, u0_u12_X_41, 
       u0_u12_X_43, u0_u12_X_47, u0_u12_X_6, u0_u12_X_8, u0_u12_X_9, u0_u12_u0_n100, u0_u12_u0_n101, u0_u12_u0_n102, u0_u12_u0_n103, 
       u0_u12_u0_n104, u0_u12_u0_n105, u0_u12_u0_n106, u0_u12_u0_n107, u0_u12_u0_n108, u0_u12_u0_n109, u0_u12_u0_n110, u0_u12_u0_n111, u0_u12_u0_n112, 
       u0_u12_u0_n113, u0_u12_u0_n114, u0_u12_u0_n115, u0_u12_u0_n116, u0_u12_u0_n117, u0_u12_u0_n118, u0_u12_u0_n119, u0_u12_u0_n120, u0_u12_u0_n121, 
       u0_u12_u0_n122, u0_u12_u0_n123, u0_u12_u0_n124, u0_u12_u0_n125, u0_u12_u0_n126, u0_u12_u0_n127, u0_u12_u0_n128, u0_u12_u0_n129, u0_u12_u0_n130, 
       u0_u12_u0_n131, u0_u12_u0_n132, u0_u12_u0_n133, u0_u12_u0_n134, u0_u12_u0_n135, u0_u12_u0_n136, u0_u12_u0_n137, u0_u12_u0_n138, u0_u12_u0_n139, 
       u0_u12_u0_n140, u0_u12_u0_n141, u0_u12_u0_n142, u0_u12_u0_n143, u0_u12_u0_n144, u0_u12_u0_n145, u0_u12_u0_n146, u0_u12_u0_n147, u0_u12_u0_n148, 
       u0_u12_u0_n149, u0_u12_u0_n150, u0_u12_u0_n151, u0_u12_u0_n152, u0_u12_u0_n153, u0_u12_u0_n154, u0_u12_u0_n155, u0_u12_u0_n156, u0_u12_u0_n157, 
       u0_u12_u0_n158, u0_u12_u0_n159, u0_u12_u0_n160, u0_u12_u0_n161, u0_u12_u0_n162, u0_u12_u0_n163, u0_u12_u0_n164, u0_u12_u0_n165, u0_u12_u0_n166, 
       u0_u12_u0_n167, u0_u12_u0_n168, u0_u12_u0_n169, u0_u12_u0_n170, u0_u12_u0_n171, u0_u12_u0_n172, u0_u12_u0_n173, u0_u12_u0_n174, u0_u12_u0_n88, 
       u0_u12_u0_n89, u0_u12_u0_n90, u0_u12_u0_n91, u0_u12_u0_n92, u0_u12_u0_n93, u0_u12_u0_n94, u0_u12_u0_n95, u0_u12_u0_n96, u0_u12_u0_n97, 
       u0_u12_u0_n98, u0_u12_u0_n99, u0_u12_u1_n100, u0_u12_u1_n101, u0_u12_u1_n102, u0_u12_u1_n103, u0_u12_u1_n104, u0_u12_u1_n105, u0_u12_u1_n106, 
       u0_u12_u1_n107, u0_u12_u1_n108, u0_u12_u1_n109, u0_u12_u1_n110, u0_u12_u1_n111, u0_u12_u1_n112, u0_u12_u1_n113, u0_u12_u1_n114, u0_u12_u1_n115, 
       u0_u12_u1_n116, u0_u12_u1_n117, u0_u12_u1_n118, u0_u12_u1_n119, u0_u12_u1_n120, u0_u12_u1_n121, u0_u12_u1_n122, u0_u12_u1_n123, u0_u12_u1_n124, 
       u0_u12_u1_n125, u0_u12_u1_n126, u0_u12_u1_n127, u0_u12_u1_n128, u0_u12_u1_n129, u0_u12_u1_n130, u0_u12_u1_n131, u0_u12_u1_n132, u0_u12_u1_n133, 
       u0_u12_u1_n134, u0_u12_u1_n135, u0_u12_u1_n136, u0_u12_u1_n137, u0_u12_u1_n138, u0_u12_u1_n139, u0_u12_u1_n140, u0_u12_u1_n141, u0_u12_u1_n142, 
       u0_u12_u1_n143, u0_u12_u1_n144, u0_u12_u1_n145, u0_u12_u1_n146, u0_u12_u1_n147, u0_u12_u1_n148, u0_u12_u1_n149, u0_u12_u1_n150, u0_u12_u1_n151, 
       u0_u12_u1_n152, u0_u12_u1_n153, u0_u12_u1_n154, u0_u12_u1_n155, u0_u12_u1_n156, u0_u12_u1_n157, u0_u12_u1_n158, u0_u12_u1_n159, u0_u12_u1_n160, 
       u0_u12_u1_n161, u0_u12_u1_n162, u0_u12_u1_n163, u0_u12_u1_n164, u0_u12_u1_n165, u0_u12_u1_n166, u0_u12_u1_n167, u0_u12_u1_n168, u0_u12_u1_n169, 
       u0_u12_u1_n170, u0_u12_u1_n171, u0_u12_u1_n172, u0_u12_u1_n173, u0_u12_u1_n174, u0_u12_u1_n175, u0_u12_u1_n176, u0_u12_u1_n177, u0_u12_u1_n178, 
       u0_u12_u1_n179, u0_u12_u1_n180, u0_u12_u1_n181, u0_u12_u1_n182, u0_u12_u1_n183, u0_u12_u1_n184, u0_u12_u1_n185, u0_u12_u1_n186, u0_u12_u1_n187, 
       u0_u12_u1_n188, u0_u12_u1_n95, u0_u12_u1_n96, u0_u12_u1_n97, u0_u12_u1_n98, u0_u12_u1_n99, u0_u12_u2_n100, u0_u12_u2_n101, u0_u12_u2_n102, 
       u0_u12_u2_n103, u0_u12_u2_n104, u0_u12_u2_n105, u0_u12_u2_n106, u0_u12_u2_n107, u0_u12_u2_n108, u0_u12_u2_n109, u0_u12_u2_n110, u0_u12_u2_n111, 
       u0_u12_u2_n112, u0_u12_u2_n113, u0_u12_u2_n114, u0_u12_u2_n115, u0_u12_u2_n116, u0_u12_u2_n117, u0_u12_u2_n118, u0_u12_u2_n119, u0_u12_u2_n120, 
       u0_u12_u2_n121, u0_u12_u2_n122, u0_u12_u2_n123, u0_u12_u2_n124, u0_u12_u2_n125, u0_u12_u2_n126, u0_u12_u2_n127, u0_u12_u2_n128, u0_u12_u2_n129, 
       u0_u12_u2_n130, u0_u12_u2_n131, u0_u12_u2_n132, u0_u12_u2_n133, u0_u12_u2_n134, u0_u12_u2_n135, u0_u12_u2_n136, u0_u12_u2_n137, u0_u12_u2_n138, 
       u0_u12_u2_n139, u0_u12_u2_n140, u0_u12_u2_n141, u0_u12_u2_n142, u0_u12_u2_n143, u0_u12_u2_n144, u0_u12_u2_n145, u0_u12_u2_n146, u0_u12_u2_n147, 
       u0_u12_u2_n148, u0_u12_u2_n149, u0_u12_u2_n150, u0_u12_u2_n151, u0_u12_u2_n152, u0_u12_u2_n153, u0_u12_u2_n154, u0_u12_u2_n155, u0_u12_u2_n156, 
       u0_u12_u2_n157, u0_u12_u2_n158, u0_u12_u2_n159, u0_u12_u2_n160, u0_u12_u2_n161, u0_u12_u2_n162, u0_u12_u2_n163, u0_u12_u2_n164, u0_u12_u2_n165, 
       u0_u12_u2_n166, u0_u12_u2_n167, u0_u12_u2_n168, u0_u12_u2_n169, u0_u12_u2_n170, u0_u12_u2_n171, u0_u12_u2_n172, u0_u12_u2_n173, u0_u12_u2_n174, 
       u0_u12_u2_n175, u0_u12_u2_n176, u0_u12_u2_n177, u0_u12_u2_n178, u0_u12_u2_n179, u0_u12_u2_n180, u0_u12_u2_n181, u0_u12_u2_n182, u0_u12_u2_n183, 
       u0_u12_u2_n184, u0_u12_u2_n185, u0_u12_u2_n186, u0_u12_u2_n187, u0_u12_u2_n188, u0_u12_u2_n95, u0_u12_u2_n96, u0_u12_u2_n97, u0_u12_u2_n98, 
       u0_u12_u2_n99, u0_u12_u3_n100, u0_u12_u3_n101, u0_u12_u3_n102, u0_u12_u3_n103, u0_u12_u3_n104, u0_u12_u3_n105, u0_u12_u3_n106, u0_u12_u3_n107, 
       u0_u12_u3_n108, u0_u12_u3_n109, u0_u12_u3_n110, u0_u12_u3_n111, u0_u12_u3_n112, u0_u12_u3_n113, u0_u12_u3_n114, u0_u12_u3_n115, u0_u12_u3_n116, 
       u0_u12_u3_n117, u0_u12_u3_n118, u0_u12_u3_n119, u0_u12_u3_n120, u0_u12_u3_n121, u0_u12_u3_n122, u0_u12_u3_n123, u0_u12_u3_n124, u0_u12_u3_n125, 
       u0_u12_u3_n126, u0_u12_u3_n127, u0_u12_u3_n128, u0_u12_u3_n129, u0_u12_u3_n130, u0_u12_u3_n131, u0_u12_u3_n132, u0_u12_u3_n133, u0_u12_u3_n134, 
       u0_u12_u3_n135, u0_u12_u3_n136, u0_u12_u3_n137, u0_u12_u3_n138, u0_u12_u3_n139, u0_u12_u3_n140, u0_u12_u3_n141, u0_u12_u3_n142, u0_u12_u3_n143, 
       u0_u12_u3_n144, u0_u12_u3_n145, u0_u12_u3_n146, u0_u12_u3_n147, u0_u12_u3_n148, u0_u12_u3_n149, u0_u12_u3_n150, u0_u12_u3_n151, u0_u12_u3_n152, 
       u0_u12_u3_n153, u0_u12_u3_n154, u0_u12_u3_n155, u0_u12_u3_n156, u0_u12_u3_n157, u0_u12_u3_n158, u0_u12_u3_n159, u0_u12_u3_n160, u0_u12_u3_n161, 
       u0_u12_u3_n162, u0_u12_u3_n163, u0_u12_u3_n164, u0_u12_u3_n165, u0_u12_u3_n166, u0_u12_u3_n167, u0_u12_u3_n168, u0_u12_u3_n169, u0_u12_u3_n170, 
       u0_u12_u3_n171, u0_u12_u3_n172, u0_u12_u3_n173, u0_u12_u3_n174, u0_u12_u3_n175, u0_u12_u3_n176, u0_u12_u3_n177, u0_u12_u3_n178, u0_u12_u3_n179, 
       u0_u12_u3_n180, u0_u12_u3_n181, u0_u12_u3_n182, u0_u12_u3_n183, u0_u12_u3_n184, u0_u12_u3_n185, u0_u12_u3_n186, u0_u12_u3_n94, u0_u12_u3_n95, 
       u0_u12_u3_n96, u0_u12_u3_n97, u0_u12_u3_n98, u0_u12_u3_n99, u0_u12_u6_n100, u0_u12_u6_n101, u0_u12_u6_n102, u0_u12_u6_n103, u0_u12_u6_n104, 
       u0_u12_u6_n105, u0_u12_u6_n106, u0_u12_u6_n107, u0_u12_u6_n108, u0_u12_u6_n109, u0_u12_u6_n110, u0_u12_u6_n111, u0_u12_u6_n112, u0_u12_u6_n113, 
       u0_u12_u6_n114, u0_u12_u6_n115, u0_u12_u6_n116, u0_u12_u6_n117, u0_u12_u6_n118, u0_u12_u6_n119, u0_u12_u6_n120, u0_u12_u6_n121, u0_u12_u6_n122, 
       u0_u12_u6_n123, u0_u12_u6_n124, u0_u12_u6_n125, u0_u12_u6_n126, u0_u12_u6_n127, u0_u12_u6_n128, u0_u12_u6_n129, u0_u12_u6_n130, u0_u12_u6_n131, 
       u0_u12_u6_n132, u0_u12_u6_n133, u0_u12_u6_n134, u0_u12_u6_n135, u0_u12_u6_n136, u0_u12_u6_n137, u0_u12_u6_n138, u0_u12_u6_n139, u0_u12_u6_n140, 
       u0_u12_u6_n141, u0_u12_u6_n142, u0_u12_u6_n143, u0_u12_u6_n144, u0_u12_u6_n145, u0_u12_u6_n146, u0_u12_u6_n147, u0_u12_u6_n148, u0_u12_u6_n149, 
       u0_u12_u6_n150, u0_u12_u6_n151, u0_u12_u6_n152, u0_u12_u6_n153, u0_u12_u6_n154, u0_u12_u6_n155, u0_u12_u6_n156, u0_u12_u6_n157, u0_u12_u6_n158, 
       u0_u12_u6_n159, u0_u12_u6_n160, u0_u12_u6_n161, u0_u12_u6_n162, u0_u12_u6_n163, u0_u12_u6_n164, u0_u12_u6_n165, u0_u12_u6_n166, u0_u12_u6_n167, 
       u0_u12_u6_n168, u0_u12_u6_n169, u0_u12_u6_n170, u0_u12_u6_n171, u0_u12_u6_n172, u0_u12_u6_n173, u0_u12_u6_n174, u0_u12_u6_n88, u0_u12_u6_n89, 
       u0_u12_u6_n90, u0_u12_u6_n91, u0_u12_u6_n92, u0_u12_u6_n93, u0_u12_u6_n94, u0_u12_u6_n95, u0_u12_u6_n96, u0_u12_u6_n97, u0_u12_u6_n98, 
       u0_u12_u6_n99, u0_u12_u7_n100, u0_u12_u7_n101, u0_u12_u7_n102, u0_u12_u7_n103, u0_u12_u7_n104, u0_u12_u7_n105, u0_u12_u7_n106, u0_u12_u7_n107, 
       u0_u12_u7_n108, u0_u12_u7_n109, u0_u12_u7_n110, u0_u12_u7_n111, u0_u12_u7_n112, u0_u12_u7_n113, u0_u12_u7_n114, u0_u12_u7_n115, u0_u12_u7_n116, 
       u0_u12_u7_n117, u0_u12_u7_n118, u0_u12_u7_n119, u0_u12_u7_n120, u0_u12_u7_n121, u0_u12_u7_n122, u0_u12_u7_n123, u0_u12_u7_n124, u0_u12_u7_n125, 
       u0_u12_u7_n126, u0_u12_u7_n127, u0_u12_u7_n128, u0_u12_u7_n129, u0_u12_u7_n130, u0_u12_u7_n131, u0_u12_u7_n132, u0_u12_u7_n133, u0_u12_u7_n134, 
       u0_u12_u7_n135, u0_u12_u7_n136, u0_u12_u7_n137, u0_u12_u7_n138, u0_u12_u7_n139, u0_u12_u7_n140, u0_u12_u7_n141, u0_u12_u7_n142, u0_u12_u7_n143, 
       u0_u12_u7_n144, u0_u12_u7_n145, u0_u12_u7_n146, u0_u12_u7_n147, u0_u12_u7_n148, u0_u12_u7_n149, u0_u12_u7_n150, u0_u12_u7_n151, u0_u12_u7_n152, 
       u0_u12_u7_n153, u0_u12_u7_n154, u0_u12_u7_n155, u0_u12_u7_n156, u0_u12_u7_n157, u0_u12_u7_n158, u0_u12_u7_n159, u0_u12_u7_n160, u0_u12_u7_n161, 
       u0_u12_u7_n162, u0_u12_u7_n163, u0_u12_u7_n164, u0_u12_u7_n165, u0_u12_u7_n166, u0_u12_u7_n167, u0_u12_u7_n168, u0_u12_u7_n169, u0_u12_u7_n170, 
       u0_u12_u7_n171, u0_u12_u7_n172, u0_u12_u7_n173, u0_u12_u7_n174, u0_u12_u7_n175, u0_u12_u7_n176, u0_u12_u7_n177, u0_u12_u7_n178, u0_u12_u7_n179, 
       u0_u12_u7_n180, u0_u12_u7_n91, u0_u12_u7_n92, u0_u12_u7_n93, u0_u12_u7_n94, u0_u12_u7_n95, u0_u12_u7_n96, u0_u12_u7_n97, u0_u12_u7_n98, 
       u0_u12_u7_n99, u0_u13_X_45, u0_u13_u7_n100, u0_u13_u7_n101, u0_u13_u7_n102, u0_u13_u7_n103, u0_u13_u7_n104, u0_u13_u7_n105, u0_u13_u7_n106, 
       u0_u13_u7_n107, u0_u13_u7_n108, u0_u13_u7_n109, u0_u13_u7_n110, u0_u13_u7_n111, u0_u13_u7_n112, u0_u13_u7_n113, u0_u13_u7_n114, u0_u13_u7_n115, 
       u0_u13_u7_n116, u0_u13_u7_n117, u0_u13_u7_n118, u0_u13_u7_n119, u0_u13_u7_n120, u0_u13_u7_n121, u0_u13_u7_n122, u0_u13_u7_n123, u0_u13_u7_n124, 
       u0_u13_u7_n125, u0_u13_u7_n126, u0_u13_u7_n127, u0_u13_u7_n128, u0_u13_u7_n129, u0_u13_u7_n130, u0_u13_u7_n131, u0_u13_u7_n132, u0_u13_u7_n133, 
       u0_u13_u7_n134, u0_u13_u7_n135, u0_u13_u7_n136, u0_u13_u7_n137, u0_u13_u7_n138, u0_u13_u7_n139, u0_u13_u7_n140, u0_u13_u7_n141, u0_u13_u7_n142, 
       u0_u13_u7_n143, u0_u13_u7_n144, u0_u13_u7_n145, u0_u13_u7_n146, u0_u13_u7_n147, u0_u13_u7_n148, u0_u13_u7_n149, u0_u13_u7_n150, u0_u13_u7_n151, 
       u0_u13_u7_n152, u0_u13_u7_n153, u0_u13_u7_n154, u0_u13_u7_n155, u0_u13_u7_n156, u0_u13_u7_n157, u0_u13_u7_n158, u0_u13_u7_n159, u0_u13_u7_n160, 
       u0_u13_u7_n161, u0_u13_u7_n162, u0_u13_u7_n163, u0_u13_u7_n164, u0_u13_u7_n165, u0_u13_u7_n166, u0_u13_u7_n167, u0_u13_u7_n168, u0_u13_u7_n169, 
       u0_u13_u7_n170, u0_u13_u7_n171, u0_u13_u7_n172, u0_u13_u7_n173, u0_u13_u7_n174, u0_u13_u7_n175, u0_u13_u7_n176, u0_u13_u7_n177, u0_u13_u7_n178, 
       u0_u13_u7_n179, u0_u13_u7_n180, u0_u13_u7_n91, u0_u13_u7_n92, u0_u13_u7_n93, u0_u13_u7_n94, u0_u13_u7_n95, u0_u13_u7_n96, u0_u13_u7_n97, 
       u0_u13_u7_n98, u0_u13_u7_n99, u0_u14_X_11, u0_u14_X_13, u0_u14_u1_n100, u0_u14_u1_n101, u0_u14_u1_n102, u0_u14_u1_n103, u0_u14_u1_n104, 
       u0_u14_u1_n105, u0_u14_u1_n106, u0_u14_u1_n107, u0_u14_u1_n108, u0_u14_u1_n109, u0_u14_u1_n110, u0_u14_u1_n111, u0_u14_u1_n112, u0_u14_u1_n113, 
       u0_u14_u1_n114, u0_u14_u1_n115, u0_u14_u1_n116, u0_u14_u1_n117, u0_u14_u1_n118, u0_u14_u1_n119, u0_u14_u1_n120, u0_u14_u1_n121, u0_u14_u1_n122, 
       u0_u14_u1_n123, u0_u14_u1_n124, u0_u14_u1_n125, u0_u14_u1_n126, u0_u14_u1_n127, u0_u14_u1_n128, u0_u14_u1_n129, u0_u14_u1_n130, u0_u14_u1_n131, 
       u0_u14_u1_n132, u0_u14_u1_n133, u0_u14_u1_n134, u0_u14_u1_n135, u0_u14_u1_n136, u0_u14_u1_n137, u0_u14_u1_n138, u0_u14_u1_n139, u0_u14_u1_n140, 
       u0_u14_u1_n141, u0_u14_u1_n142, u0_u14_u1_n143, u0_u14_u1_n144, u0_u14_u1_n145, u0_u14_u1_n146, u0_u14_u1_n147, u0_u14_u1_n148, u0_u14_u1_n149, 
       u0_u14_u1_n150, u0_u14_u1_n151, u0_u14_u1_n152, u0_u14_u1_n153, u0_u14_u1_n154, u0_u14_u1_n155, u0_u14_u1_n156, u0_u14_u1_n157, u0_u14_u1_n158, 
       u0_u14_u1_n159, u0_u14_u1_n160, u0_u14_u1_n161, u0_u14_u1_n162, u0_u14_u1_n163, u0_u14_u1_n164, u0_u14_u1_n165, u0_u14_u1_n166, u0_u14_u1_n167, 
       u0_u14_u1_n168, u0_u14_u1_n169, u0_u14_u1_n170, u0_u14_u1_n171, u0_u14_u1_n172, u0_u14_u1_n173, u0_u14_u1_n174, u0_u14_u1_n175, u0_u14_u1_n176, 
       u0_u14_u1_n177, u0_u14_u1_n178, u0_u14_u1_n179, u0_u14_u1_n180, u0_u14_u1_n181, u0_u14_u1_n182, u0_u14_u1_n183, u0_u14_u1_n184, u0_u14_u1_n185, 
       u0_u14_u1_n186, u0_u14_u1_n187, u0_u14_u1_n188, u0_u14_u1_n95, u0_u14_u1_n96, u0_u14_u1_n97, u0_u14_u1_n98, u0_u14_u1_n99, u0_u14_u2_n100, 
       u0_u14_u2_n101, u0_u14_u2_n102, u0_u14_u2_n103, u0_u14_u2_n104, u0_u14_u2_n105, u0_u14_u2_n106, u0_u14_u2_n107, u0_u14_u2_n108, u0_u14_u2_n109, 
       u0_u14_u2_n110, u0_u14_u2_n111, u0_u14_u2_n112, u0_u14_u2_n113, u0_u14_u2_n114, u0_u14_u2_n115, u0_u14_u2_n116, u0_u14_u2_n117, u0_u14_u2_n118, 
       u0_u14_u2_n119, u0_u14_u2_n120, u0_u14_u2_n121, u0_u14_u2_n122, u0_u14_u2_n123, u0_u14_u2_n124, u0_u14_u2_n125, u0_u14_u2_n126, u0_u14_u2_n127, 
       u0_u14_u2_n128, u0_u14_u2_n129, u0_u14_u2_n130, u0_u14_u2_n131, u0_u14_u2_n132, u0_u14_u2_n133, u0_u14_u2_n134, u0_u14_u2_n135, u0_u14_u2_n136, 
       u0_u14_u2_n137, u0_u14_u2_n138, u0_u14_u2_n139, u0_u14_u2_n140, u0_u14_u2_n141, u0_u14_u2_n142, u0_u14_u2_n143, u0_u14_u2_n144, u0_u14_u2_n145, 
       u0_u14_u2_n146, u0_u14_u2_n147, u0_u14_u2_n148, u0_u14_u2_n149, u0_u14_u2_n150, u0_u14_u2_n151, u0_u14_u2_n152, u0_u14_u2_n153, u0_u14_u2_n154, 
       u0_u14_u2_n155, u0_u14_u2_n156, u0_u14_u2_n157, u0_u14_u2_n158, u0_u14_u2_n159, u0_u14_u2_n160, u0_u14_u2_n161, u0_u14_u2_n162, u0_u14_u2_n163, 
       u0_u14_u2_n164, u0_u14_u2_n165, u0_u14_u2_n166, u0_u14_u2_n167, u0_u14_u2_n168, u0_u14_u2_n169, u0_u14_u2_n170, u0_u14_u2_n171, u0_u14_u2_n172, 
       u0_u14_u2_n173, u0_u14_u2_n174, u0_u14_u2_n175, u0_u14_u2_n176, u0_u14_u2_n177, u0_u14_u2_n178, u0_u14_u2_n179, u0_u14_u2_n180, u0_u14_u2_n181, 
       u0_u14_u2_n182, u0_u14_u2_n183, u0_u14_u2_n184, u0_u14_u2_n185, u0_u14_u2_n186, u0_u14_u2_n187, u0_u14_u2_n188, u0_u14_u2_n95, u0_u14_u2_n96, 
       u0_u14_u2_n97, u0_u14_u2_n98, u0_u14_u2_n99, u0_u14_u3_n100, u0_u14_u3_n101, u0_u14_u3_n102, u0_u14_u3_n103, u0_u14_u3_n104, u0_u14_u3_n105, 
       u0_u14_u3_n106, u0_u14_u3_n107, u0_u14_u3_n108, u0_u14_u3_n109, u0_u14_u3_n110, u0_u14_u3_n111, u0_u14_u3_n112, u0_u14_u3_n113, u0_u14_u3_n114, 
       u0_u14_u3_n115, u0_u14_u3_n116, u0_u14_u3_n117, u0_u14_u3_n118, u0_u14_u3_n119, u0_u14_u3_n120, u0_u14_u3_n121, u0_u14_u3_n122, u0_u14_u3_n123, 
       u0_u14_u3_n124, u0_u14_u3_n125, u0_u14_u3_n126, u0_u14_u3_n127, u0_u14_u3_n128, u0_u14_u3_n129, u0_u14_u3_n130, u0_u14_u3_n131, u0_u14_u3_n132, 
       u0_u14_u3_n133, u0_u14_u3_n134, u0_u14_u3_n135, u0_u14_u3_n136, u0_u14_u3_n137, u0_u14_u3_n138, u0_u14_u3_n139, u0_u14_u3_n140, u0_u14_u3_n141, 
       u0_u14_u3_n142, u0_u14_u3_n143, u0_u14_u3_n144, u0_u14_u3_n145, u0_u14_u3_n146, u0_u14_u3_n147, u0_u14_u3_n148, u0_u14_u3_n149, u0_u14_u3_n150, 
       u0_u14_u3_n151, u0_u14_u3_n152, u0_u14_u3_n153, u0_u14_u3_n154, u0_u14_u3_n155, u0_u14_u3_n156, u0_u14_u3_n157, u0_u14_u3_n158, u0_u14_u3_n159, 
       u0_u14_u3_n160, u0_u14_u3_n161, u0_u14_u3_n162, u0_u14_u3_n163, u0_u14_u3_n164, u0_u14_u3_n165, u0_u14_u3_n166, u0_u14_u3_n167, u0_u14_u3_n168, 
       u0_u14_u3_n169, u0_u14_u3_n170, u0_u14_u3_n171, u0_u14_u3_n172, u0_u14_u3_n173, u0_u14_u3_n174, u0_u14_u3_n175, u0_u14_u3_n176, u0_u14_u3_n177, 
       u0_u14_u3_n178, u0_u14_u3_n179, u0_u14_u3_n180, u0_u14_u3_n181, u0_u14_u3_n182, u0_u14_u3_n183, u0_u14_u3_n184, u0_u14_u3_n185, u0_u14_u3_n186, 
       u0_u14_u3_n94, u0_u14_u3_n95, u0_u14_u3_n96, u0_u14_u3_n97, u0_u14_u3_n98, u0_u14_u3_n99, u0_u15_X_37, u0_u15_X_38, u0_u15_X_39, 
       u0_u15_X_40, u0_u15_X_41, u0_u15_u6_n100, u0_u15_u6_n101, u0_u15_u6_n102, u0_u15_u6_n103, u0_u15_u6_n104, u0_u15_u6_n105, u0_u15_u6_n106, 
       u0_u15_u6_n107, u0_u15_u6_n108, u0_u15_u6_n109, u0_u15_u6_n110, u0_u15_u6_n111, u0_u15_u6_n112, u0_u15_u6_n113, u0_u15_u6_n114, u0_u15_u6_n115, 
       u0_u15_u6_n116, u0_u15_u6_n117, u0_u15_u6_n118, u0_u15_u6_n119, u0_u15_u6_n120, u0_u15_u6_n121, u0_u15_u6_n122, u0_u15_u6_n123, u0_u15_u6_n124, 
       u0_u15_u6_n125, u0_u15_u6_n126, u0_u15_u6_n127, u0_u15_u6_n128, u0_u15_u6_n129, u0_u15_u6_n130, u0_u15_u6_n131, u0_u15_u6_n132, u0_u15_u6_n133, 
       u0_u15_u6_n134, u0_u15_u6_n135, u0_u15_u6_n136, u0_u15_u6_n137, u0_u15_u6_n138, u0_u15_u6_n139, u0_u15_u6_n140, u0_u15_u6_n141, u0_u15_u6_n142, 
       u0_u15_u6_n143, u0_u15_u6_n144, u0_u15_u6_n145, u0_u15_u6_n146, u0_u15_u6_n147, u0_u15_u6_n148, u0_u15_u6_n149, u0_u15_u6_n150, u0_u15_u6_n151, 
       u0_u15_u6_n152, u0_u15_u6_n153, u0_u15_u6_n154, u0_u15_u6_n155, u0_u15_u6_n156, u0_u15_u6_n157, u0_u15_u6_n158, u0_u15_u6_n159, u0_u15_u6_n160, 
       u0_u15_u6_n161, u0_u15_u6_n162, u0_u15_u6_n163, u0_u15_u6_n164, u0_u15_u6_n165, u0_u15_u6_n166, u0_u15_u6_n167, u0_u15_u6_n168, u0_u15_u6_n169, 
       u0_u15_u6_n170, u0_u15_u6_n171, u0_u15_u6_n172, u0_u15_u6_n173, u0_u15_u6_n174, u0_u15_u6_n88, u0_u15_u6_n89, u0_u15_u6_n90, u0_u15_u6_n91, 
       u0_u15_u6_n92, u0_u15_u6_n93, u0_u15_u6_n94, u0_u15_u6_n95, u0_u15_u6_n96, u0_u15_u6_n97, u0_u15_u6_n98, u0_u15_u6_n99, u0_u1_X_27, 
       u0_u1_X_28, u0_u1_X_29, u0_u1_X_30, u0_u1_X_31, u0_u1_X_32, u0_u1_X_41, u0_u1_u4_n100, u0_u1_u4_n101, u0_u1_u4_n102, 
       u0_u1_u4_n103, u0_u1_u4_n104, u0_u1_u4_n105, u0_u1_u4_n106, u0_u1_u4_n107, u0_u1_u4_n108, u0_u1_u4_n109, u0_u1_u4_n110, u0_u1_u4_n111, 
       u0_u1_u4_n112, u0_u1_u4_n113, u0_u1_u4_n114, u0_u1_u4_n115, u0_u1_u4_n116, u0_u1_u4_n117, u0_u1_u4_n118, u0_u1_u4_n119, u0_u1_u4_n120, 
       u0_u1_u4_n121, u0_u1_u4_n122, u0_u1_u4_n123, u0_u1_u4_n124, u0_u1_u4_n125, u0_u1_u4_n126, u0_u1_u4_n127, u0_u1_u4_n128, u0_u1_u4_n129, 
       u0_u1_u4_n130, u0_u1_u4_n131, u0_u1_u4_n132, u0_u1_u4_n133, u0_u1_u4_n134, u0_u1_u4_n135, u0_u1_u4_n136, u0_u1_u4_n137, u0_u1_u4_n138, 
       u0_u1_u4_n139, u0_u1_u4_n140, u0_u1_u4_n141, u0_u1_u4_n142, u0_u1_u4_n143, u0_u1_u4_n144, u0_u1_u4_n145, u0_u1_u4_n146, u0_u1_u4_n147, 
       u0_u1_u4_n148, u0_u1_u4_n149, u0_u1_u4_n150, u0_u1_u4_n151, u0_u1_u4_n152, u0_u1_u4_n153, u0_u1_u4_n154, u0_u1_u4_n155, u0_u1_u4_n156, 
       u0_u1_u4_n157, u0_u1_u4_n158, u0_u1_u4_n159, u0_u1_u4_n160, u0_u1_u4_n161, u0_u1_u4_n162, u0_u1_u4_n163, u0_u1_u4_n164, u0_u1_u4_n165, 
       u0_u1_u4_n166, u0_u1_u4_n167, u0_u1_u4_n168, u0_u1_u4_n169, u0_u1_u4_n170, u0_u1_u4_n171, u0_u1_u4_n172, u0_u1_u4_n173, u0_u1_u4_n174, 
       u0_u1_u4_n175, u0_u1_u4_n176, u0_u1_u4_n177, u0_u1_u4_n178, u0_u1_u4_n179, u0_u1_u4_n180, u0_u1_u4_n181, u0_u1_u4_n182, u0_u1_u4_n183, 
       u0_u1_u4_n184, u0_u1_u4_n185, u0_u1_u4_n186, u0_u1_u4_n94, u0_u1_u4_n95, u0_u1_u4_n96, u0_u1_u4_n97, u0_u1_u4_n98, u0_u1_u4_n99, 
       u0_u1_u5_n100, u0_u1_u5_n101, u0_u1_u5_n102, u0_u1_u5_n103, u0_u1_u5_n104, u0_u1_u5_n105, u0_u1_u5_n106, u0_u1_u5_n107, u0_u1_u5_n108, 
       u0_u1_u5_n109, u0_u1_u5_n110, u0_u1_u5_n111, u0_u1_u5_n112, u0_u1_u5_n113, u0_u1_u5_n114, u0_u1_u5_n115, u0_u1_u5_n116, u0_u1_u5_n117, 
       u0_u1_u5_n118, u0_u1_u5_n119, u0_u1_u5_n120, u0_u1_u5_n121, u0_u1_u5_n122, u0_u1_u5_n123, u0_u1_u5_n124, u0_u1_u5_n125, u0_u1_u5_n126, 
       u0_u1_u5_n127, u0_u1_u5_n128, u0_u1_u5_n129, u0_u1_u5_n130, u0_u1_u5_n131, u0_u1_u5_n132, u0_u1_u5_n133, u0_u1_u5_n134, u0_u1_u5_n135, 
       u0_u1_u5_n136, u0_u1_u5_n137, u0_u1_u5_n138, u0_u1_u5_n139, u0_u1_u5_n140, u0_u1_u5_n141, u0_u1_u5_n142, u0_u1_u5_n143, u0_u1_u5_n144, 
       u0_u1_u5_n145, u0_u1_u5_n146, u0_u1_u5_n147, u0_u1_u5_n148, u0_u1_u5_n149, u0_u1_u5_n150, u0_u1_u5_n151, u0_u1_u5_n152, u0_u1_u5_n153, 
       u0_u1_u5_n154, u0_u1_u5_n155, u0_u1_u5_n156, u0_u1_u5_n157, u0_u1_u5_n158, u0_u1_u5_n159, u0_u1_u5_n160, u0_u1_u5_n161, u0_u1_u5_n162, 
       u0_u1_u5_n163, u0_u1_u5_n164, u0_u1_u5_n165, u0_u1_u5_n166, u0_u1_u5_n167, u0_u1_u5_n168, u0_u1_u5_n169, u0_u1_u5_n170, u0_u1_u5_n171, 
       u0_u1_u5_n172, u0_u1_u5_n173, u0_u1_u5_n174, u0_u1_u5_n175, u0_u1_u5_n176, u0_u1_u5_n177, u0_u1_u5_n178, u0_u1_u5_n179, u0_u1_u5_n180, 
       u0_u1_u5_n181, u0_u1_u5_n182, u0_u1_u5_n183, u0_u1_u5_n184, u0_u1_u5_n185, u0_u1_u5_n186, u0_u1_u5_n187, u0_u1_u5_n188, u0_u1_u5_n189, 
       u0_u1_u5_n190, u0_u1_u5_n191, u0_u1_u5_n192, u0_u1_u5_n193, u0_u1_u5_n194, u0_u1_u5_n195, u0_u1_u5_n196, u0_u1_u5_n99, u0_u1_u6_n100, 
       u0_u1_u6_n101, u0_u1_u6_n102, u0_u1_u6_n103, u0_u1_u6_n104, u0_u1_u6_n105, u0_u1_u6_n106, u0_u1_u6_n107, u0_u1_u6_n108, u0_u1_u6_n109, 
       u0_u1_u6_n110, u0_u1_u6_n111, u0_u1_u6_n112, u0_u1_u6_n113, u0_u1_u6_n114, u0_u1_u6_n115, u0_u1_u6_n116, u0_u1_u6_n117, u0_u1_u6_n118, 
       u0_u1_u6_n119, u0_u1_u6_n120, u0_u1_u6_n121, u0_u1_u6_n122, u0_u1_u6_n123, u0_u1_u6_n124, u0_u1_u6_n125, u0_u1_u6_n126, u0_u1_u6_n127, 
       u0_u1_u6_n128, u0_u1_u6_n129, u0_u1_u6_n130, u0_u1_u6_n131, u0_u1_u6_n132, u0_u1_u6_n133, u0_u1_u6_n134, u0_u1_u6_n135, u0_u1_u6_n136, 
       u0_u1_u6_n137, u0_u1_u6_n138, u0_u1_u6_n139, u0_u1_u6_n140, u0_u1_u6_n141, u0_u1_u6_n142, u0_u1_u6_n143, u0_u1_u6_n144, u0_u1_u6_n145, 
       u0_u1_u6_n146, u0_u1_u6_n147, u0_u1_u6_n148, u0_u1_u6_n149, u0_u1_u6_n150, u0_u1_u6_n151, u0_u1_u6_n152, u0_u1_u6_n153, u0_u1_u6_n154, 
       u0_u1_u6_n155, u0_u1_u6_n156, u0_u1_u6_n157, u0_u1_u6_n158, u0_u1_u6_n159, u0_u1_u6_n160, u0_u1_u6_n161, u0_u1_u6_n162, u0_u1_u6_n163, 
       u0_u1_u6_n164, u0_u1_u6_n165, u0_u1_u6_n166, u0_u1_u6_n167, u0_u1_u6_n168, u0_u1_u6_n169, u0_u1_u6_n170, u0_u1_u6_n171, u0_u1_u6_n172, 
       u0_u1_u6_n173, u0_u1_u6_n174, u0_u1_u6_n88, u0_u1_u6_n89, u0_u1_u6_n90, u0_u1_u6_n91, u0_u1_u6_n92, u0_u1_u6_n93, u0_u1_u6_n94, 
       u0_u1_u6_n95, u0_u1_u6_n96, u0_u1_u6_n97, u0_u1_u6_n98, u0_u1_u6_n99, u0_u2_X_1, u0_u2_X_11, u0_u2_X_12, u0_u2_X_13, 
       u0_u2_X_14, u0_u2_X_17, u0_u2_X_18, u0_u2_X_2, u0_u2_X_4, u0_u2_X_5, u0_u2_X_6, u0_u2_X_7, u0_u2_X_8, 
       u0_u2_u0_n100, u0_u2_u0_n101, u0_u2_u0_n102, u0_u2_u0_n103, u0_u2_u0_n104, u0_u2_u0_n105, u0_u2_u0_n106, u0_u2_u0_n107, u0_u2_u0_n108, 
       u0_u2_u0_n109, u0_u2_u0_n110, u0_u2_u0_n111, u0_u2_u0_n112, u0_u2_u0_n113, u0_u2_u0_n114, u0_u2_u0_n115, u0_u2_u0_n116, u0_u2_u0_n117, 
       u0_u2_u0_n118, u0_u2_u0_n119, u0_u2_u0_n120, u0_u2_u0_n121, u0_u2_u0_n122, u0_u2_u0_n123, u0_u2_u0_n124, u0_u2_u0_n125, u0_u2_u0_n126, 
       u0_u2_u0_n127, u0_u2_u0_n128, u0_u2_u0_n129, u0_u2_u0_n130, u0_u2_u0_n131, u0_u2_u0_n132, u0_u2_u0_n133, u0_u2_u0_n134, u0_u2_u0_n135, 
       u0_u2_u0_n136, u0_u2_u0_n137, u0_u2_u0_n138, u0_u2_u0_n139, u0_u2_u0_n140, u0_u2_u0_n141, u0_u2_u0_n142, u0_u2_u0_n143, u0_u2_u0_n144, 
       u0_u2_u0_n145, u0_u2_u0_n146, u0_u2_u0_n147, u0_u2_u0_n148, u0_u2_u0_n149, u0_u2_u0_n150, u0_u2_u0_n151, u0_u2_u0_n152, u0_u2_u0_n153, 
       u0_u2_u0_n154, u0_u2_u0_n155, u0_u2_u0_n156, u0_u2_u0_n157, u0_u2_u0_n158, u0_u2_u0_n159, u0_u2_u0_n160, u0_u2_u0_n161, u0_u2_u0_n162, 
       u0_u2_u0_n163, u0_u2_u0_n164, u0_u2_u0_n165, u0_u2_u0_n166, u0_u2_u0_n167, u0_u2_u0_n168, u0_u2_u0_n169, u0_u2_u0_n170, u0_u2_u0_n171, 
       u0_u2_u0_n172, u0_u2_u0_n173, u0_u2_u0_n174, u0_u2_u0_n88, u0_u2_u0_n89, u0_u2_u0_n90, u0_u2_u0_n91, u0_u2_u0_n92, u0_u2_u0_n93, 
       u0_u2_u0_n94, u0_u2_u0_n95, u0_u2_u0_n96, u0_u2_u0_n97, u0_u2_u0_n98, u0_u2_u0_n99, u0_u2_u1_n100, u0_u2_u1_n101, u0_u2_u1_n102, 
       u0_u2_u1_n103, u0_u2_u1_n104, u0_u2_u1_n105, u0_u2_u1_n106, u0_u2_u1_n107, u0_u2_u1_n108, u0_u2_u1_n109, u0_u2_u1_n110, u0_u2_u1_n111, 
       u0_u2_u1_n112, u0_u2_u1_n113, u0_u2_u1_n114, u0_u2_u1_n115, u0_u2_u1_n116, u0_u2_u1_n117, u0_u2_u1_n118, u0_u2_u1_n119, u0_u2_u1_n120, 
       u0_u2_u1_n121, u0_u2_u1_n122, u0_u2_u1_n123, u0_u2_u1_n124, u0_u2_u1_n125, u0_u2_u1_n126, u0_u2_u1_n127, u0_u2_u1_n128, u0_u2_u1_n129, 
       u0_u2_u1_n130, u0_u2_u1_n131, u0_u2_u1_n132, u0_u2_u1_n133, u0_u2_u1_n134, u0_u2_u1_n135, u0_u2_u1_n136, u0_u2_u1_n137, u0_u2_u1_n138, 
       u0_u2_u1_n139, u0_u2_u1_n140, u0_u2_u1_n141, u0_u2_u1_n142, u0_u2_u1_n143, u0_u2_u1_n144, u0_u2_u1_n145, u0_u2_u1_n146, u0_u2_u1_n147, 
       u0_u2_u1_n148, u0_u2_u1_n149, u0_u2_u1_n150, u0_u2_u1_n151, u0_u2_u1_n152, u0_u2_u1_n153, u0_u2_u1_n154, u0_u2_u1_n155, u0_u2_u1_n156, 
       u0_u2_u1_n157, u0_u2_u1_n158, u0_u2_u1_n159, u0_u2_u1_n160, u0_u2_u1_n161, u0_u2_u1_n162, u0_u2_u1_n163, u0_u2_u1_n164, u0_u2_u1_n165, 
       u0_u2_u1_n166, u0_u2_u1_n167, u0_u2_u1_n168, u0_u2_u1_n169, u0_u2_u1_n170, u0_u2_u1_n171, u0_u2_u1_n172, u0_u2_u1_n173, u0_u2_u1_n174, 
       u0_u2_u1_n175, u0_u2_u1_n176, u0_u2_u1_n177, u0_u2_u1_n178, u0_u2_u1_n179, u0_u2_u1_n180, u0_u2_u1_n181, u0_u2_u1_n182, u0_u2_u1_n183, 
       u0_u2_u1_n184, u0_u2_u1_n185, u0_u2_u1_n186, u0_u2_u1_n187, u0_u2_u1_n188, u0_u2_u1_n95, u0_u2_u1_n96, u0_u2_u1_n97, u0_u2_u1_n98, 
       u0_u2_u1_n99, u0_u2_u2_n100, u0_u2_u2_n101, u0_u2_u2_n102, u0_u2_u2_n103, u0_u2_u2_n104, u0_u2_u2_n105, u0_u2_u2_n106, u0_u2_u2_n107, 
       u0_u2_u2_n108, u0_u2_u2_n109, u0_u2_u2_n110, u0_u2_u2_n111, u0_u2_u2_n112, u0_u2_u2_n113, u0_u2_u2_n114, u0_u2_u2_n115, u0_u2_u2_n116, 
       u0_u2_u2_n117, u0_u2_u2_n118, u0_u2_u2_n119, u0_u2_u2_n120, u0_u2_u2_n121, u0_u2_u2_n122, u0_u2_u2_n123, u0_u2_u2_n124, u0_u2_u2_n125, 
       u0_u2_u2_n126, u0_u2_u2_n127, u0_u2_u2_n128, u0_u2_u2_n129, u0_u2_u2_n130, u0_u2_u2_n131, u0_u2_u2_n132, u0_u2_u2_n133, u0_u2_u2_n134, 
       u0_u2_u2_n135, u0_u2_u2_n136, u0_u2_u2_n137, u0_u2_u2_n138, u0_u2_u2_n139, u0_u2_u2_n140, u0_u2_u2_n141, u0_u2_u2_n142, u0_u2_u2_n143, 
       u0_u2_u2_n144, u0_u2_u2_n145, u0_u2_u2_n146, u0_u2_u2_n147, u0_u2_u2_n148, u0_u2_u2_n149, u0_u2_u2_n150, u0_u2_u2_n151, u0_u2_u2_n152, 
       u0_u2_u2_n153, u0_u2_u2_n154, u0_u2_u2_n155, u0_u2_u2_n156, u0_u2_u2_n157, u0_u2_u2_n158, u0_u2_u2_n159, u0_u2_u2_n160, u0_u2_u2_n161, 
       u0_u2_u2_n162, u0_u2_u2_n163, u0_u2_u2_n164, u0_u2_u2_n165, u0_u2_u2_n166, u0_u2_u2_n167, u0_u2_u2_n168, u0_u2_u2_n169, u0_u2_u2_n170, 
       u0_u2_u2_n171, u0_u2_u2_n172, u0_u2_u2_n173, u0_u2_u2_n174, u0_u2_u2_n175, u0_u2_u2_n176, u0_u2_u2_n177, u0_u2_u2_n178, u0_u2_u2_n179, 
       u0_u2_u2_n180, u0_u2_u2_n181, u0_u2_u2_n182, u0_u2_u2_n183, u0_u2_u2_n184, u0_u2_u2_n185, u0_u2_u2_n186, u0_u2_u2_n187, u0_u2_u2_n188, 
       u0_u2_u2_n95, u0_u2_u2_n96, u0_u2_u2_n97, u0_u2_u2_n98, u0_u2_u2_n99, u0_u5_X_1, u0_u5_X_11, u0_u5_X_12, u0_u5_X_13, 
       u0_u5_X_14, u0_u5_X_17, u0_u5_X_18, u0_u5_X_19, u0_u5_X_2, u0_u5_X_20, u0_u5_X_23, u0_u5_X_24, u0_u5_X_25, 
       u0_u5_X_26, u0_u5_X_28, u0_u5_X_29, u0_u5_X_30, u0_u5_X_31, u0_u5_X_32, u0_u5_X_33, u0_u5_X_35, u0_u5_X_36, 
       u0_u5_X_37, u0_u5_X_38, u0_u5_X_39, u0_u5_X_4, u0_u5_X_40, u0_u5_X_41, u0_u5_X_42, u0_u5_X_43, u0_u5_X_44, 
       u0_u5_X_45, u0_u5_X_47, u0_u5_X_48, u0_u5_X_5, u0_u5_X_6, u0_u5_X_7, u0_u5_X_8, u0_u5_u0_n100, u0_u5_u0_n101, 
       u0_u5_u0_n102, u0_u5_u0_n103, u0_u5_u0_n104, u0_u5_u0_n105, u0_u5_u0_n106, u0_u5_u0_n107, u0_u5_u0_n108, u0_u5_u0_n109, u0_u5_u0_n110, 
       u0_u5_u0_n111, u0_u5_u0_n112, u0_u5_u0_n113, u0_u5_u0_n114, u0_u5_u0_n115, u0_u5_u0_n116, u0_u5_u0_n117, u0_u5_u0_n118, u0_u5_u0_n119, 
       u0_u5_u0_n120, u0_u5_u0_n121, u0_u5_u0_n122, u0_u5_u0_n123, u0_u5_u0_n124, u0_u5_u0_n125, u0_u5_u0_n126, u0_u5_u0_n127, u0_u5_u0_n128, 
       u0_u5_u0_n129, u0_u5_u0_n130, u0_u5_u0_n131, u0_u5_u0_n132, u0_u5_u0_n133, u0_u5_u0_n134, u0_u5_u0_n135, u0_u5_u0_n136, u0_u5_u0_n137, 
       u0_u5_u0_n138, u0_u5_u0_n139, u0_u5_u0_n140, u0_u5_u0_n141, u0_u5_u0_n142, u0_u5_u0_n143, u0_u5_u0_n144, u0_u5_u0_n145, u0_u5_u0_n146, 
       u0_u5_u0_n147, u0_u5_u0_n148, u0_u5_u0_n149, u0_u5_u0_n150, u0_u5_u0_n151, u0_u5_u0_n152, u0_u5_u0_n153, u0_u5_u0_n154, u0_u5_u0_n155, 
       u0_u5_u0_n156, u0_u5_u0_n157, u0_u5_u0_n158, u0_u5_u0_n159, u0_u5_u0_n160, u0_u5_u0_n161, u0_u5_u0_n162, u0_u5_u0_n163, u0_u5_u0_n164, 
       u0_u5_u0_n165, u0_u5_u0_n166, u0_u5_u0_n167, u0_u5_u0_n168, u0_u5_u0_n169, u0_u5_u0_n170, u0_u5_u0_n171, u0_u5_u0_n172, u0_u5_u0_n173, 
       u0_u5_u0_n174, u0_u5_u0_n88, u0_u5_u0_n89, u0_u5_u0_n90, u0_u5_u0_n91, u0_u5_u0_n92, u0_u5_u0_n93, u0_u5_u0_n94, u0_u5_u0_n95, 
       u0_u5_u0_n96, u0_u5_u0_n97, u0_u5_u0_n98, u0_u5_u0_n99, u0_u5_u1_n100, u0_u5_u1_n101, u0_u5_u1_n102, u0_u5_u1_n103, u0_u5_u1_n104, 
       u0_u5_u1_n105, u0_u5_u1_n106, u0_u5_u1_n107, u0_u5_u1_n108, u0_u5_u1_n109, u0_u5_u1_n110, u0_u5_u1_n111, u0_u5_u1_n112, u0_u5_u1_n113, 
       u0_u5_u1_n114, u0_u5_u1_n115, u0_u5_u1_n116, u0_u5_u1_n117, u0_u5_u1_n118, u0_u5_u1_n119, u0_u5_u1_n120, u0_u5_u1_n121, u0_u5_u1_n122, 
       u0_u5_u1_n123, u0_u5_u1_n124, u0_u5_u1_n125, u0_u5_u1_n126, u0_u5_u1_n127, u0_u5_u1_n128, u0_u5_u1_n129, u0_u5_u1_n130, u0_u5_u1_n131, 
       u0_u5_u1_n132, u0_u5_u1_n133, u0_u5_u1_n134, u0_u5_u1_n135, u0_u5_u1_n136, u0_u5_u1_n137, u0_u5_u1_n138, u0_u5_u1_n139, u0_u5_u1_n140, 
       u0_u5_u1_n141, u0_u5_u1_n142, u0_u5_u1_n143, u0_u5_u1_n144, u0_u5_u1_n145, u0_u5_u1_n146, u0_u5_u1_n147, u0_u5_u1_n148, u0_u5_u1_n149, 
       u0_u5_u1_n150, u0_u5_u1_n151, u0_u5_u1_n152, u0_u5_u1_n153, u0_u5_u1_n154, u0_u5_u1_n155, u0_u5_u1_n156, u0_u5_u1_n157, u0_u5_u1_n158, 
       u0_u5_u1_n159, u0_u5_u1_n160, u0_u5_u1_n161, u0_u5_u1_n162, u0_u5_u1_n163, u0_u5_u1_n164, u0_u5_u1_n165, u0_u5_u1_n166, u0_u5_u1_n167, 
       u0_u5_u1_n168, u0_u5_u1_n169, u0_u5_u1_n170, u0_u5_u1_n171, u0_u5_u1_n172, u0_u5_u1_n173, u0_u5_u1_n174, u0_u5_u1_n175, u0_u5_u1_n176, 
       u0_u5_u1_n177, u0_u5_u1_n178, u0_u5_u1_n179, u0_u5_u1_n180, u0_u5_u1_n181, u0_u5_u1_n182, u0_u5_u1_n183, u0_u5_u1_n184, u0_u5_u1_n185, 
       u0_u5_u1_n186, u0_u5_u1_n187, u0_u5_u1_n188, u0_u5_u1_n95, u0_u5_u1_n96, u0_u5_u1_n97, u0_u5_u1_n98, u0_u5_u1_n99, u0_u5_u2_n100, 
       u0_u5_u2_n101, u0_u5_u2_n102, u0_u5_u2_n103, u0_u5_u2_n104, u0_u5_u2_n105, u0_u5_u2_n106, u0_u5_u2_n107, u0_u5_u2_n108, u0_u5_u2_n109, 
       u0_u5_u2_n110, u0_u5_u2_n111, u0_u5_u2_n112, u0_u5_u2_n113, u0_u5_u2_n114, u0_u5_u2_n115, u0_u5_u2_n116, u0_u5_u2_n117, u0_u5_u2_n118, 
       u0_u5_u2_n119, u0_u5_u2_n120, u0_u5_u2_n121, u0_u5_u2_n122, u0_u5_u2_n123, u0_u5_u2_n124, u0_u5_u2_n125, u0_u5_u2_n126, u0_u5_u2_n127, 
       u0_u5_u2_n128, u0_u5_u2_n129, u0_u5_u2_n130, u0_u5_u2_n131, u0_u5_u2_n132, u0_u5_u2_n133, u0_u5_u2_n134, u0_u5_u2_n135, u0_u5_u2_n136, 
       u0_u5_u2_n137, u0_u5_u2_n138, u0_u5_u2_n139, u0_u5_u2_n140, u0_u5_u2_n141, u0_u5_u2_n142, u0_u5_u2_n143, u0_u5_u2_n144, u0_u5_u2_n145, 
       u0_u5_u2_n146, u0_u5_u2_n147, u0_u5_u2_n148, u0_u5_u2_n149, u0_u5_u2_n150, u0_u5_u2_n151, u0_u5_u2_n152, u0_u5_u2_n153, u0_u5_u2_n154, 
       u0_u5_u2_n155, u0_u5_u2_n156, u0_u5_u2_n157, u0_u5_u2_n158, u0_u5_u2_n159, u0_u5_u2_n160, u0_u5_u2_n161, u0_u5_u2_n162, u0_u5_u2_n163, 
       u0_u5_u2_n164, u0_u5_u2_n165, u0_u5_u2_n166, u0_u5_u2_n167, u0_u5_u2_n168, u0_u5_u2_n169, u0_u5_u2_n170, u0_u5_u2_n171, u0_u5_u2_n172, 
       u0_u5_u2_n173, u0_u5_u2_n174, u0_u5_u2_n175, u0_u5_u2_n176, u0_u5_u2_n177, u0_u5_u2_n178, u0_u5_u2_n179, u0_u5_u2_n180, u0_u5_u2_n181, 
       u0_u5_u2_n182, u0_u5_u2_n183, u0_u5_u2_n184, u0_u5_u2_n185, u0_u5_u2_n186, u0_u5_u2_n187, u0_u5_u2_n188, u0_u5_u2_n95, u0_u5_u2_n96, 
       u0_u5_u2_n97, u0_u5_u2_n98, u0_u5_u2_n99, u0_u5_u3_n100, u0_u5_u3_n101, u0_u5_u3_n102, u0_u5_u3_n103, u0_u5_u3_n104, u0_u5_u3_n105, 
       u0_u5_u3_n106, u0_u5_u3_n107, u0_u5_u3_n108, u0_u5_u3_n109, u0_u5_u3_n110, u0_u5_u3_n111, u0_u5_u3_n112, u0_u5_u3_n113, u0_u5_u3_n114, 
       u0_u5_u3_n115, u0_u5_u3_n116, u0_u5_u3_n117, u0_u5_u3_n118, u0_u5_u3_n119, u0_u5_u3_n120, u0_u5_u3_n121, u0_u5_u3_n122, u0_u5_u3_n123, 
       u0_u5_u3_n124, u0_u5_u3_n125, u0_u5_u3_n126, u0_u5_u3_n127, u0_u5_u3_n128, u0_u5_u3_n129, u0_u5_u3_n130, u0_u5_u3_n131, u0_u5_u3_n132, 
       u0_u5_u3_n133, u0_u5_u3_n134, u0_u5_u3_n135, u0_u5_u3_n136, u0_u5_u3_n137, u0_u5_u3_n138, u0_u5_u3_n139, u0_u5_u3_n140, u0_u5_u3_n141, 
       u0_u5_u3_n142, u0_u5_u3_n143, u0_u5_u3_n144, u0_u5_u3_n145, u0_u5_u3_n146, u0_u5_u3_n147, u0_u5_u3_n148, u0_u5_u3_n149, u0_u5_u3_n150, 
       u0_u5_u3_n151, u0_u5_u3_n152, u0_u5_u3_n153, u0_u5_u3_n154, u0_u5_u3_n155, u0_u5_u3_n156, u0_u5_u3_n157, u0_u5_u3_n158, u0_u5_u3_n159, 
       u0_u5_u3_n160, u0_u5_u3_n161, u0_u5_u3_n162, u0_u5_u3_n163, u0_u5_u3_n164, u0_u5_u3_n165, u0_u5_u3_n166, u0_u5_u3_n167, u0_u5_u3_n168, 
       u0_u5_u3_n169, u0_u5_u3_n170, u0_u5_u3_n171, u0_u5_u3_n172, u0_u5_u3_n173, u0_u5_u3_n174, u0_u5_u3_n175, u0_u5_u3_n176, u0_u5_u3_n177, 
       u0_u5_u3_n178, u0_u5_u3_n179, u0_u5_u3_n180, u0_u5_u3_n181, u0_u5_u3_n182, u0_u5_u3_n183, u0_u5_u3_n184, u0_u5_u3_n185, u0_u5_u3_n186, 
       u0_u5_u3_n94, u0_u5_u3_n95, u0_u5_u3_n96, u0_u5_u3_n97, u0_u5_u3_n98, u0_u5_u3_n99, u0_u5_u4_n100, u0_u5_u4_n101, u0_u5_u4_n102, 
       u0_u5_u4_n103, u0_u5_u4_n104, u0_u5_u4_n105, u0_u5_u4_n106, u0_u5_u4_n107, u0_u5_u4_n108, u0_u5_u4_n109, u0_u5_u4_n110, u0_u5_u4_n111, 
       u0_u5_u4_n112, u0_u5_u4_n113, u0_u5_u4_n114, u0_u5_u4_n115, u0_u5_u4_n116, u0_u5_u4_n117, u0_u5_u4_n118, u0_u5_u4_n119, u0_u5_u4_n120, 
       u0_u5_u4_n121, u0_u5_u4_n122, u0_u5_u4_n123, u0_u5_u4_n124, u0_u5_u4_n125, u0_u5_u4_n126, u0_u5_u4_n127, u0_u5_u4_n128, u0_u5_u4_n129, 
       u0_u5_u4_n130, u0_u5_u4_n131, u0_u5_u4_n132, u0_u5_u4_n133, u0_u5_u4_n134, u0_u5_u4_n135, u0_u5_u4_n136, u0_u5_u4_n137, u0_u5_u4_n138, 
       u0_u5_u4_n139, u0_u5_u4_n140, u0_u5_u4_n141, u0_u5_u4_n142, u0_u5_u4_n143, u0_u5_u4_n144, u0_u5_u4_n145, u0_u5_u4_n146, u0_u5_u4_n147, 
       u0_u5_u4_n148, u0_u5_u4_n149, u0_u5_u4_n150, u0_u5_u4_n151, u0_u5_u4_n152, u0_u5_u4_n153, u0_u5_u4_n154, u0_u5_u4_n155, u0_u5_u4_n156, 
       u0_u5_u4_n157, u0_u5_u4_n158, u0_u5_u4_n159, u0_u5_u4_n160, u0_u5_u4_n161, u0_u5_u4_n162, u0_u5_u4_n163, u0_u5_u4_n164, u0_u5_u4_n165, 
       u0_u5_u4_n166, u0_u5_u4_n167, u0_u5_u4_n168, u0_u5_u4_n169, u0_u5_u4_n170, u0_u5_u4_n171, u0_u5_u4_n172, u0_u5_u4_n173, u0_u5_u4_n174, 
       u0_u5_u4_n175, u0_u5_u4_n176, u0_u5_u4_n177, u0_u5_u4_n178, u0_u5_u4_n179, u0_u5_u4_n180, u0_u5_u4_n181, u0_u5_u4_n182, u0_u5_u4_n183, 
       u0_u5_u4_n184, u0_u5_u4_n185, u0_u5_u4_n186, u0_u5_u4_n94, u0_u5_u4_n95, u0_u5_u4_n96, u0_u5_u4_n97, u0_u5_u4_n98, u0_u5_u4_n99, 
       u0_u5_u5_n100, u0_u5_u5_n101, u0_u5_u5_n102, u0_u5_u5_n103, u0_u5_u5_n104, u0_u5_u5_n105, u0_u5_u5_n106, u0_u5_u5_n107, u0_u5_u5_n108, 
       u0_u5_u5_n109, u0_u5_u5_n110, u0_u5_u5_n111, u0_u5_u5_n112, u0_u5_u5_n113, u0_u5_u5_n114, u0_u5_u5_n115, u0_u5_u5_n116, u0_u5_u5_n117, 
       u0_u5_u5_n118, u0_u5_u5_n119, u0_u5_u5_n120, u0_u5_u5_n121, u0_u5_u5_n122, u0_u5_u5_n123, u0_u5_u5_n124, u0_u5_u5_n125, u0_u5_u5_n126, 
       u0_u5_u5_n127, u0_u5_u5_n128, u0_u5_u5_n129, u0_u5_u5_n130, u0_u5_u5_n131, u0_u5_u5_n132, u0_u5_u5_n133, u0_u5_u5_n134, u0_u5_u5_n135, 
       u0_u5_u5_n136, u0_u5_u5_n137, u0_u5_u5_n138, u0_u5_u5_n139, u0_u5_u5_n140, u0_u5_u5_n141, u0_u5_u5_n142, u0_u5_u5_n143, u0_u5_u5_n144, 
       u0_u5_u5_n145, u0_u5_u5_n146, u0_u5_u5_n147, u0_u5_u5_n148, u0_u5_u5_n149, u0_u5_u5_n150, u0_u5_u5_n151, u0_u5_u5_n152, u0_u5_u5_n153, 
       u0_u5_u5_n154, u0_u5_u5_n155, u0_u5_u5_n156, u0_u5_u5_n157, u0_u5_u5_n158, u0_u5_u5_n159, u0_u5_u5_n160, u0_u5_u5_n161, u0_u5_u5_n162, 
       u0_u5_u5_n163, u0_u5_u5_n164, u0_u5_u5_n165, u0_u5_u5_n166, u0_u5_u5_n167, u0_u5_u5_n168, u0_u5_u5_n169, u0_u5_u5_n170, u0_u5_u5_n171, 
       u0_u5_u5_n172, u0_u5_u5_n173, u0_u5_u5_n174, u0_u5_u5_n175, u0_u5_u5_n176, u0_u5_u5_n177, u0_u5_u5_n178, u0_u5_u5_n179, u0_u5_u5_n180, 
       u0_u5_u5_n181, u0_u5_u5_n182, u0_u5_u5_n183, u0_u5_u5_n184, u0_u5_u5_n185, u0_u5_u5_n186, u0_u5_u5_n187, u0_u5_u5_n188, u0_u5_u5_n189, 
       u0_u5_u5_n190, u0_u5_u5_n191, u0_u5_u5_n192, u0_u5_u5_n193, u0_u5_u5_n194, u0_u5_u5_n195, u0_u5_u5_n196, u0_u5_u5_n99, u0_u5_u6_n100, 
       u0_u5_u6_n101, u0_u5_u6_n102, u0_u5_u6_n103, u0_u5_u6_n104, u0_u5_u6_n105, u0_u5_u6_n106, u0_u5_u6_n107, u0_u5_u6_n108, u0_u5_u6_n109, 
       u0_u5_u6_n110, u0_u5_u6_n111, u0_u5_u6_n112, u0_u5_u6_n113, u0_u5_u6_n114, u0_u5_u6_n115, u0_u5_u6_n116, u0_u5_u6_n117, u0_u5_u6_n118, 
       u0_u5_u6_n119, u0_u5_u6_n120, u0_u5_u6_n121, u0_u5_u6_n122, u0_u5_u6_n123, u0_u5_u6_n124, u0_u5_u6_n125, u0_u5_u6_n126, u0_u5_u6_n127, 
       u0_u5_u6_n128, u0_u5_u6_n129, u0_u5_u6_n130, u0_u5_u6_n131, u0_u5_u6_n132, u0_u5_u6_n133, u0_u5_u6_n134, u0_u5_u6_n135, u0_u5_u6_n136, 
       u0_u5_u6_n137, u0_u5_u6_n138, u0_u5_u6_n139, u0_u5_u6_n140, u0_u5_u6_n141, u0_u5_u6_n142, u0_u5_u6_n143, u0_u5_u6_n144, u0_u5_u6_n145, 
       u0_u5_u6_n146, u0_u5_u6_n147, u0_u5_u6_n148, u0_u5_u6_n149, u0_u5_u6_n150, u0_u5_u6_n151, u0_u5_u6_n152, u0_u5_u6_n153, u0_u5_u6_n154, 
       u0_u5_u6_n155, u0_u5_u6_n156, u0_u5_u6_n157, u0_u5_u6_n158, u0_u5_u6_n159, u0_u5_u6_n160, u0_u5_u6_n161, u0_u5_u6_n162, u0_u5_u6_n163, 
       u0_u5_u6_n164, u0_u5_u6_n165, u0_u5_u6_n166, u0_u5_u6_n167, u0_u5_u6_n168, u0_u5_u6_n169, u0_u5_u6_n170, u0_u5_u6_n171, u0_u5_u6_n172, 
       u0_u5_u6_n173, u0_u5_u6_n174, u0_u5_u6_n88, u0_u5_u6_n89, u0_u5_u6_n90, u0_u5_u6_n91, u0_u5_u6_n92, u0_u5_u6_n93, u0_u5_u6_n94, 
       u0_u5_u6_n95, u0_u5_u6_n96, u0_u5_u6_n97, u0_u5_u6_n98, u0_u5_u6_n99, u0_u5_u7_n100, u0_u5_u7_n101, u0_u5_u7_n102, u0_u5_u7_n103, 
       u0_u5_u7_n104, u0_u5_u7_n105, u0_u5_u7_n106, u0_u5_u7_n107, u0_u5_u7_n108, u0_u5_u7_n109, u0_u5_u7_n110, u0_u5_u7_n111, u0_u5_u7_n112, 
       u0_u5_u7_n113, u0_u5_u7_n114, u0_u5_u7_n115, u0_u5_u7_n116, u0_u5_u7_n117, u0_u5_u7_n118, u0_u5_u7_n119, u0_u5_u7_n120, u0_u5_u7_n121, 
       u0_u5_u7_n122, u0_u5_u7_n123, u0_u5_u7_n124, u0_u5_u7_n125, u0_u5_u7_n126, u0_u5_u7_n127, u0_u5_u7_n128, u0_u5_u7_n129, u0_u5_u7_n130, 
       u0_u5_u7_n131, u0_u5_u7_n132, u0_u5_u7_n133, u0_u5_u7_n134, u0_u5_u7_n135, u0_u5_u7_n136, u0_u5_u7_n137, u0_u5_u7_n138, u0_u5_u7_n139, 
       u0_u5_u7_n140, u0_u5_u7_n141, u0_u5_u7_n142, u0_u5_u7_n143, u0_u5_u7_n144, u0_u5_u7_n145, u0_u5_u7_n146, u0_u5_u7_n147, u0_u5_u7_n148, 
       u0_u5_u7_n149, u0_u5_u7_n150, u0_u5_u7_n151, u0_u5_u7_n152, u0_u5_u7_n153, u0_u5_u7_n154, u0_u5_u7_n155, u0_u5_u7_n156, u0_u5_u7_n157, 
       u0_u5_u7_n158, u0_u5_u7_n159, u0_u5_u7_n160, u0_u5_u7_n161, u0_u5_u7_n162, u0_u5_u7_n163, u0_u5_u7_n164, u0_u5_u7_n165, u0_u5_u7_n166, 
       u0_u5_u7_n167, u0_u5_u7_n168, u0_u5_u7_n169, u0_u5_u7_n170, u0_u5_u7_n171, u0_u5_u7_n172, u0_u5_u7_n173, u0_u5_u7_n174, u0_u5_u7_n175, 
       u0_u5_u7_n176, u0_u5_u7_n177, u0_u5_u7_n178, u0_u5_u7_n179, u0_u5_u7_n180, u0_u5_u7_n91, u0_u5_u7_n92, u0_u5_u7_n93, u0_u5_u7_n94, 
       u0_u5_u7_n95, u0_u5_u7_n96, u0_u5_u7_n97, u0_u5_u7_n98, u0_u5_u7_n99, u0_uk_n1003, u0_uk_n673, u0_uk_n679, u0_uk_n683, 
       u0_uk_n703, u0_uk_n704, u0_uk_n708, u0_uk_n712, u0_uk_n713, u0_uk_n787, u0_uk_n788, u0_uk_n789, u0_uk_n791, 
       u0_uk_n794, u0_uk_n795, u0_uk_n858, u0_uk_n860, u0_uk_n861, u0_uk_n862, u0_uk_n881, u0_uk_n886, u0_uk_n887, 
       u0_uk_n891, u0_uk_n893, u0_uk_n899, u0_uk_n900, u0_uk_n924, u0_uk_n929, u0_uk_n940, u0_uk_n943, u0_uk_n944, 
       u0_uk_n951, u0_uk_n952, u0_uk_n953, u0_uk_n954, u0_uk_n955, u0_uk_n966, u0_uk_n972, u0_uk_n973, u0_uk_n975, 
       u0_uk_n979, u0_uk_n983, u0_uk_n996, u1_K10_33, u1_K10_35, u1_K10_37, u1_K10_38, u1_K11_12, u1_K11_14, 
       u1_K11_17, u1_K11_31, u1_K11_34, u1_K11_36, u1_K11_5, u1_K13_11, u1_K13_12, u1_K13_13, u1_K13_15, 
       u1_K13_19, u1_K13_2, u1_K13_5, u1_K13_6, u1_K13_7, u1_K15_26, u1_K15_30, u1_K15_38, u1_K15_43, 
       u1_K15_8, u1_K16_29, u1_K16_34, u1_K1_41, u1_K2_19, u1_K2_41, u1_K4_10, u1_K4_2, u1_K4_3, 
       u1_K4_8, u1_K5_20, u1_K5_22, u1_K7_12, u1_K7_13, u1_K7_42, u1_K7_46, u1_K7_6, u1_K7_8, 
       u1_K9_1, u1_K9_19, u1_K9_2, u1_K9_20, u1_K9_22, u1_K9_26, u1_K9_27, u1_K9_35, u1_K9_41, 
       u1_K9_42, u1_K9_48, u1_u0_X_1, u1_u0_X_41, u1_u0_X_43, u1_u0_X_47, u1_u0_X_6, u1_u0_X_8, u1_u0_u0_n100, 
       u1_u0_u0_n101, u1_u0_u0_n102, u1_u0_u0_n103, u1_u0_u0_n104, u1_u0_u0_n105, u1_u0_u0_n106, u1_u0_u0_n107, u1_u0_u0_n108, u1_u0_u0_n109, 
       u1_u0_u0_n110, u1_u0_u0_n111, u1_u0_u0_n112, u1_u0_u0_n113, u1_u0_u0_n114, u1_u0_u0_n115, u1_u0_u0_n116, u1_u0_u0_n117, u1_u0_u0_n118, 
       u1_u0_u0_n119, u1_u0_u0_n120, u1_u0_u0_n121, u1_u0_u0_n122, u1_u0_u0_n123, u1_u0_u0_n124, u1_u0_u0_n125, u1_u0_u0_n126, u1_u0_u0_n127, 
       u1_u0_u0_n128, u1_u0_u0_n129, u1_u0_u0_n130, u1_u0_u0_n131, u1_u0_u0_n132, u1_u0_u0_n133, u1_u0_u0_n134, u1_u0_u0_n135, u1_u0_u0_n136, 
       u1_u0_u0_n137, u1_u0_u0_n138, u1_u0_u0_n139, u1_u0_u0_n140, u1_u0_u0_n141, u1_u0_u0_n142, u1_u0_u0_n143, u1_u0_u0_n144, u1_u0_u0_n145, 
       u1_u0_u0_n146, u1_u0_u0_n147, u1_u0_u0_n148, u1_u0_u0_n149, u1_u0_u0_n150, u1_u0_u0_n151, u1_u0_u0_n152, u1_u0_u0_n153, u1_u0_u0_n154, 
       u1_u0_u0_n155, u1_u0_u0_n156, u1_u0_u0_n157, u1_u0_u0_n158, u1_u0_u0_n159, u1_u0_u0_n160, u1_u0_u0_n161, u1_u0_u0_n162, u1_u0_u0_n163, 
       u1_u0_u0_n164, u1_u0_u0_n165, u1_u0_u0_n166, u1_u0_u0_n167, u1_u0_u0_n168, u1_u0_u0_n169, u1_u0_u0_n170, u1_u0_u0_n171, u1_u0_u0_n172, 
       u1_u0_u0_n173, u1_u0_u0_n174, u1_u0_u0_n88, u1_u0_u0_n89, u1_u0_u0_n90, u1_u0_u0_n91, u1_u0_u0_n92, u1_u0_u0_n93, u1_u0_u0_n94, 
       u1_u0_u0_n95, u1_u0_u0_n96, u1_u0_u0_n97, u1_u0_u0_n98, u1_u0_u0_n99, u1_u0_u1_n100, u1_u0_u1_n101, u1_u0_u1_n102, u1_u0_u1_n103, 
       u1_u0_u1_n104, u1_u0_u1_n105, u1_u0_u1_n106, u1_u0_u1_n107, u1_u0_u1_n108, u1_u0_u1_n109, u1_u0_u1_n110, u1_u0_u1_n111, u1_u0_u1_n112, 
       u1_u0_u1_n113, u1_u0_u1_n114, u1_u0_u1_n115, u1_u0_u1_n116, u1_u0_u1_n117, u1_u0_u1_n118, u1_u0_u1_n119, u1_u0_u1_n120, u1_u0_u1_n121, 
       u1_u0_u1_n122, u1_u0_u1_n123, u1_u0_u1_n124, u1_u0_u1_n125, u1_u0_u1_n126, u1_u0_u1_n127, u1_u0_u1_n128, u1_u0_u1_n129, u1_u0_u1_n130, 
       u1_u0_u1_n131, u1_u0_u1_n132, u1_u0_u1_n133, u1_u0_u1_n134, u1_u0_u1_n135, u1_u0_u1_n136, u1_u0_u1_n137, u1_u0_u1_n138, u1_u0_u1_n139, 
       u1_u0_u1_n140, u1_u0_u1_n141, u1_u0_u1_n142, u1_u0_u1_n143, u1_u0_u1_n144, u1_u0_u1_n145, u1_u0_u1_n146, u1_u0_u1_n147, u1_u0_u1_n148, 
       u1_u0_u1_n149, u1_u0_u1_n150, u1_u0_u1_n151, u1_u0_u1_n152, u1_u0_u1_n153, u1_u0_u1_n154, u1_u0_u1_n155, u1_u0_u1_n156, u1_u0_u1_n157, 
       u1_u0_u1_n158, u1_u0_u1_n159, u1_u0_u1_n160, u1_u0_u1_n161, u1_u0_u1_n162, u1_u0_u1_n163, u1_u0_u1_n164, u1_u0_u1_n165, u1_u0_u1_n166, 
       u1_u0_u1_n167, u1_u0_u1_n168, u1_u0_u1_n169, u1_u0_u1_n170, u1_u0_u1_n171, u1_u0_u1_n172, u1_u0_u1_n173, u1_u0_u1_n174, u1_u0_u1_n175, 
       u1_u0_u1_n176, u1_u0_u1_n177, u1_u0_u1_n178, u1_u0_u1_n179, u1_u0_u1_n180, u1_u0_u1_n181, u1_u0_u1_n182, u1_u0_u1_n183, u1_u0_u1_n184, 
       u1_u0_u1_n185, u1_u0_u1_n186, u1_u0_u1_n187, u1_u0_u1_n188, u1_u0_u1_n95, u1_u0_u1_n96, u1_u0_u1_n97, u1_u0_u1_n98, u1_u0_u1_n99, 
       u1_u0_u5_n100, u1_u0_u5_n101, u1_u0_u5_n102, u1_u0_u5_n103, u1_u0_u5_n104, u1_u0_u5_n105, u1_u0_u5_n106, u1_u0_u5_n107, u1_u0_u5_n108, 
       u1_u0_u5_n109, u1_u0_u5_n110, u1_u0_u5_n111, u1_u0_u5_n112, u1_u0_u5_n113, u1_u0_u5_n114, u1_u0_u5_n115, u1_u0_u5_n116, u1_u0_u5_n117, 
       u1_u0_u5_n118, u1_u0_u5_n119, u1_u0_u5_n120, u1_u0_u5_n121, u1_u0_u5_n122, u1_u0_u5_n123, u1_u0_u5_n124, u1_u0_u5_n125, u1_u0_u5_n126, 
       u1_u0_u5_n127, u1_u0_u5_n128, u1_u0_u5_n129, u1_u0_u5_n130, u1_u0_u5_n131, u1_u0_u5_n132, u1_u0_u5_n133, u1_u0_u5_n134, u1_u0_u5_n135, 
       u1_u0_u5_n136, u1_u0_u5_n137, u1_u0_u5_n138, u1_u0_u5_n139, u1_u0_u5_n140, u1_u0_u5_n141, u1_u0_u5_n142, u1_u0_u5_n143, u1_u0_u5_n144, 
       u1_u0_u5_n145, u1_u0_u5_n146, u1_u0_u5_n147, u1_u0_u5_n148, u1_u0_u5_n149, u1_u0_u5_n150, u1_u0_u5_n151, u1_u0_u5_n152, u1_u0_u5_n153, 
       u1_u0_u5_n154, u1_u0_u5_n155, u1_u0_u5_n156, u1_u0_u5_n157, u1_u0_u5_n158, u1_u0_u5_n159, u1_u0_u5_n160, u1_u0_u5_n161, u1_u0_u5_n162, 
       u1_u0_u5_n163, u1_u0_u5_n164, u1_u0_u5_n165, u1_u0_u5_n166, u1_u0_u5_n167, u1_u0_u5_n168, u1_u0_u5_n169, u1_u0_u5_n170, u1_u0_u5_n171, 
       u1_u0_u5_n172, u1_u0_u5_n173, u1_u0_u5_n174, u1_u0_u5_n175, u1_u0_u5_n176, u1_u0_u5_n177, u1_u0_u5_n178, u1_u0_u5_n179, u1_u0_u5_n180, 
       u1_u0_u5_n181, u1_u0_u5_n182, u1_u0_u5_n183, u1_u0_u5_n184, u1_u0_u5_n185, u1_u0_u5_n186, u1_u0_u5_n187, u1_u0_u5_n188, u1_u0_u5_n189, 
       u1_u0_u5_n190, u1_u0_u5_n191, u1_u0_u5_n192, u1_u0_u5_n193, u1_u0_u5_n194, u1_u0_u5_n195, u1_u0_u5_n196, u1_u0_u5_n99, u1_u0_u6_n100, 
       u1_u0_u6_n101, u1_u0_u6_n102, u1_u0_u6_n103, u1_u0_u6_n104, u1_u0_u6_n105, u1_u0_u6_n106, u1_u0_u6_n107, u1_u0_u6_n108, u1_u0_u6_n109, 
       u1_u0_u6_n110, u1_u0_u6_n111, u1_u0_u6_n112, u1_u0_u6_n113, u1_u0_u6_n114, u1_u0_u6_n115, u1_u0_u6_n116, u1_u0_u6_n117, u1_u0_u6_n118, 
       u1_u0_u6_n119, u1_u0_u6_n120, u1_u0_u6_n121, u1_u0_u6_n122, u1_u0_u6_n123, u1_u0_u6_n124, u1_u0_u6_n125, u1_u0_u6_n126, u1_u0_u6_n127, 
       u1_u0_u6_n128, u1_u0_u6_n129, u1_u0_u6_n130, u1_u0_u6_n131, u1_u0_u6_n132, u1_u0_u6_n133, u1_u0_u6_n134, u1_u0_u6_n135, u1_u0_u6_n136, 
       u1_u0_u6_n137, u1_u0_u6_n138, u1_u0_u6_n139, u1_u0_u6_n140, u1_u0_u6_n141, u1_u0_u6_n142, u1_u0_u6_n143, u1_u0_u6_n144, u1_u0_u6_n145, 
       u1_u0_u6_n146, u1_u0_u6_n147, u1_u0_u6_n148, u1_u0_u6_n149, u1_u0_u6_n150, u1_u0_u6_n151, u1_u0_u6_n152, u1_u0_u6_n153, u1_u0_u6_n154, 
       u1_u0_u6_n155, u1_u0_u6_n156, u1_u0_u6_n157, u1_u0_u6_n158, u1_u0_u6_n159, u1_u0_u6_n160, u1_u0_u6_n161, u1_u0_u6_n162, u1_u0_u6_n163, 
       u1_u0_u6_n164, u1_u0_u6_n165, u1_u0_u6_n166, u1_u0_u6_n167, u1_u0_u6_n168, u1_u0_u6_n169, u1_u0_u6_n170, u1_u0_u6_n171, u1_u0_u6_n172, 
       u1_u0_u6_n173, u1_u0_u6_n174, u1_u0_u6_n88, u1_u0_u6_n89, u1_u0_u6_n90, u1_u0_u6_n91, u1_u0_u6_n92, u1_u0_u6_n93, u1_u0_u6_n94, 
       u1_u0_u6_n95, u1_u0_u6_n96, u1_u0_u6_n97, u1_u0_u6_n98, u1_u0_u6_n99, u1_u0_u7_n100, u1_u0_u7_n101, u1_u0_u7_n102, u1_u0_u7_n103, 
       u1_u0_u7_n104, u1_u0_u7_n105, u1_u0_u7_n106, u1_u0_u7_n107, u1_u0_u7_n108, u1_u0_u7_n109, u1_u0_u7_n110, u1_u0_u7_n111, u1_u0_u7_n112, 
       u1_u0_u7_n113, u1_u0_u7_n114, u1_u0_u7_n115, u1_u0_u7_n116, u1_u0_u7_n117, u1_u0_u7_n118, u1_u0_u7_n119, u1_u0_u7_n120, u1_u0_u7_n121, 
       u1_u0_u7_n122, u1_u0_u7_n123, u1_u0_u7_n124, u1_u0_u7_n125, u1_u0_u7_n126, u1_u0_u7_n127, u1_u0_u7_n128, u1_u0_u7_n129, u1_u0_u7_n130, 
       u1_u0_u7_n131, u1_u0_u7_n132, u1_u0_u7_n133, u1_u0_u7_n134, u1_u0_u7_n135, u1_u0_u7_n136, u1_u0_u7_n137, u1_u0_u7_n138, u1_u0_u7_n139, 
       u1_u0_u7_n140, u1_u0_u7_n141, u1_u0_u7_n142, u1_u0_u7_n143, u1_u0_u7_n144, u1_u0_u7_n145, u1_u0_u7_n146, u1_u0_u7_n147, u1_u0_u7_n148, 
       u1_u0_u7_n149, u1_u0_u7_n150, u1_u0_u7_n151, u1_u0_u7_n152, u1_u0_u7_n153, u1_u0_u7_n154, u1_u0_u7_n155, u1_u0_u7_n156, u1_u0_u7_n157, 
       u1_u0_u7_n158, u1_u0_u7_n159, u1_u0_u7_n160, u1_u0_u7_n161, u1_u0_u7_n162, u1_u0_u7_n163, u1_u0_u7_n164, u1_u0_u7_n165, u1_u0_u7_n166, 
       u1_u0_u7_n167, u1_u0_u7_n168, u1_u0_u7_n169, u1_u0_u7_n170, u1_u0_u7_n171, u1_u0_u7_n172, u1_u0_u7_n173, u1_u0_u7_n174, u1_u0_u7_n175, 
       u1_u0_u7_n176, u1_u0_u7_n177, u1_u0_u7_n178, u1_u0_u7_n179, u1_u0_u7_n180, u1_u0_u7_n91, u1_u0_u7_n92, u1_u0_u7_n93, u1_u0_u7_n94, 
       u1_u0_u7_n95, u1_u0_u7_n96, u1_u0_u7_n97, u1_u0_u7_n98, u1_u0_u7_n99, u1_u10_X_11, u1_u10_X_12, u1_u10_X_13, u1_u10_X_14, 
       u1_u10_X_17, u1_u10_X_2, u1_u10_X_31, u1_u10_X_32, u1_u10_X_34, u1_u10_X_35, u1_u10_X_36, u1_u10_X_37, u1_u10_X_38, 
       u1_u10_X_48, u1_u10_X_5, u1_u10_X_7, u1_u10_u0_n100, u1_u10_u0_n101, u1_u10_u0_n102, u1_u10_u0_n103, u1_u10_u0_n104, u1_u10_u0_n105, 
       u1_u10_u0_n106, u1_u10_u0_n107, u1_u10_u0_n108, u1_u10_u0_n109, u1_u10_u0_n110, u1_u10_u0_n111, u1_u10_u0_n112, u1_u10_u0_n113, u1_u10_u0_n114, 
       u1_u10_u0_n115, u1_u10_u0_n116, u1_u10_u0_n117, u1_u10_u0_n118, u1_u10_u0_n119, u1_u10_u0_n120, u1_u10_u0_n121, u1_u10_u0_n122, u1_u10_u0_n123, 
       u1_u10_u0_n124, u1_u10_u0_n125, u1_u10_u0_n126, u1_u10_u0_n127, u1_u10_u0_n128, u1_u10_u0_n129, u1_u10_u0_n130, u1_u10_u0_n131, u1_u10_u0_n132, 
       u1_u10_u0_n133, u1_u10_u0_n134, u1_u10_u0_n135, u1_u10_u0_n136, u1_u10_u0_n137, u1_u10_u0_n138, u1_u10_u0_n139, u1_u10_u0_n140, u1_u10_u0_n141, 
       u1_u10_u0_n142, u1_u10_u0_n143, u1_u10_u0_n144, u1_u10_u0_n145, u1_u10_u0_n146, u1_u10_u0_n147, u1_u10_u0_n148, u1_u10_u0_n149, u1_u10_u0_n150, 
       u1_u10_u0_n151, u1_u10_u0_n152, u1_u10_u0_n153, u1_u10_u0_n154, u1_u10_u0_n155, u1_u10_u0_n156, u1_u10_u0_n157, u1_u10_u0_n158, u1_u10_u0_n159, 
       u1_u10_u0_n160, u1_u10_u0_n161, u1_u10_u0_n162, u1_u10_u0_n163, u1_u10_u0_n164, u1_u10_u0_n165, u1_u10_u0_n166, u1_u10_u0_n167, u1_u10_u0_n168, 
       u1_u10_u0_n169, u1_u10_u0_n170, u1_u10_u0_n171, u1_u10_u0_n172, u1_u10_u0_n173, u1_u10_u0_n174, u1_u10_u0_n88, u1_u10_u0_n89, u1_u10_u0_n90, 
       u1_u10_u0_n91, u1_u10_u0_n92, u1_u10_u0_n93, u1_u10_u0_n94, u1_u10_u0_n95, u1_u10_u0_n96, u1_u10_u0_n97, u1_u10_u0_n98, u1_u10_u0_n99, 
       u1_u10_u1_n100, u1_u10_u1_n101, u1_u10_u1_n102, u1_u10_u1_n103, u1_u10_u1_n104, u1_u10_u1_n105, u1_u10_u1_n106, u1_u10_u1_n107, u1_u10_u1_n108, 
       u1_u10_u1_n109, u1_u10_u1_n110, u1_u10_u1_n111, u1_u10_u1_n112, u1_u10_u1_n113, u1_u10_u1_n114, u1_u10_u1_n115, u1_u10_u1_n116, u1_u10_u1_n117, 
       u1_u10_u1_n118, u1_u10_u1_n119, u1_u10_u1_n120, u1_u10_u1_n121, u1_u10_u1_n122, u1_u10_u1_n123, u1_u10_u1_n124, u1_u10_u1_n125, u1_u10_u1_n126, 
       u1_u10_u1_n127, u1_u10_u1_n128, u1_u10_u1_n129, u1_u10_u1_n130, u1_u10_u1_n131, u1_u10_u1_n132, u1_u10_u1_n133, u1_u10_u1_n134, u1_u10_u1_n135, 
       u1_u10_u1_n136, u1_u10_u1_n137, u1_u10_u1_n138, u1_u10_u1_n139, u1_u10_u1_n140, u1_u10_u1_n141, u1_u10_u1_n142, u1_u10_u1_n143, u1_u10_u1_n144, 
       u1_u10_u1_n145, u1_u10_u1_n146, u1_u10_u1_n147, u1_u10_u1_n148, u1_u10_u1_n149, u1_u10_u1_n150, u1_u10_u1_n151, u1_u10_u1_n152, u1_u10_u1_n153, 
       u1_u10_u1_n154, u1_u10_u1_n155, u1_u10_u1_n156, u1_u10_u1_n157, u1_u10_u1_n158, u1_u10_u1_n159, u1_u10_u1_n160, u1_u10_u1_n161, u1_u10_u1_n162, 
       u1_u10_u1_n163, u1_u10_u1_n164, u1_u10_u1_n165, u1_u10_u1_n166, u1_u10_u1_n167, u1_u10_u1_n168, u1_u10_u1_n169, u1_u10_u1_n170, u1_u10_u1_n171, 
       u1_u10_u1_n172, u1_u10_u1_n173, u1_u10_u1_n174, u1_u10_u1_n175, u1_u10_u1_n176, u1_u10_u1_n177, u1_u10_u1_n178, u1_u10_u1_n179, u1_u10_u1_n180, 
       u1_u10_u1_n181, u1_u10_u1_n182, u1_u10_u1_n183, u1_u10_u1_n184, u1_u10_u1_n185, u1_u10_u1_n186, u1_u10_u1_n187, u1_u10_u1_n188, u1_u10_u1_n95, 
       u1_u10_u1_n96, u1_u10_u1_n97, u1_u10_u1_n98, u1_u10_u1_n99, u1_u10_u2_n100, u1_u10_u2_n101, u1_u10_u2_n102, u1_u10_u2_n103, u1_u10_u2_n104, 
       u1_u10_u2_n105, u1_u10_u2_n106, u1_u10_u2_n107, u1_u10_u2_n108, u1_u10_u2_n109, u1_u10_u2_n110, u1_u10_u2_n111, u1_u10_u2_n112, u1_u10_u2_n113, 
       u1_u10_u2_n114, u1_u10_u2_n115, u1_u10_u2_n116, u1_u10_u2_n117, u1_u10_u2_n118, u1_u10_u2_n119, u1_u10_u2_n120, u1_u10_u2_n121, u1_u10_u2_n122, 
       u1_u10_u2_n123, u1_u10_u2_n124, u1_u10_u2_n125, u1_u10_u2_n126, u1_u10_u2_n127, u1_u10_u2_n128, u1_u10_u2_n129, u1_u10_u2_n130, u1_u10_u2_n131, 
       u1_u10_u2_n132, u1_u10_u2_n133, u1_u10_u2_n134, u1_u10_u2_n135, u1_u10_u2_n136, u1_u10_u2_n137, u1_u10_u2_n138, u1_u10_u2_n139, u1_u10_u2_n140, 
       u1_u10_u2_n141, u1_u10_u2_n142, u1_u10_u2_n143, u1_u10_u2_n144, u1_u10_u2_n145, u1_u10_u2_n146, u1_u10_u2_n147, u1_u10_u2_n148, u1_u10_u2_n149, 
       u1_u10_u2_n150, u1_u10_u2_n151, u1_u10_u2_n152, u1_u10_u2_n153, u1_u10_u2_n154, u1_u10_u2_n155, u1_u10_u2_n156, u1_u10_u2_n157, u1_u10_u2_n158, 
       u1_u10_u2_n159, u1_u10_u2_n160, u1_u10_u2_n161, u1_u10_u2_n162, u1_u10_u2_n163, u1_u10_u2_n164, u1_u10_u2_n165, u1_u10_u2_n166, u1_u10_u2_n167, 
       u1_u10_u2_n168, u1_u10_u2_n169, u1_u10_u2_n170, u1_u10_u2_n171, u1_u10_u2_n172, u1_u10_u2_n173, u1_u10_u2_n174, u1_u10_u2_n175, u1_u10_u2_n176, 
       u1_u10_u2_n177, u1_u10_u2_n178, u1_u10_u2_n179, u1_u10_u2_n180, u1_u10_u2_n181, u1_u10_u2_n182, u1_u10_u2_n183, u1_u10_u2_n184, u1_u10_u2_n185, 
       u1_u10_u2_n186, u1_u10_u2_n187, u1_u10_u2_n188, u1_u10_u2_n95, u1_u10_u2_n96, u1_u10_u2_n97, u1_u10_u2_n98, u1_u10_u2_n99, u1_u10_u5_n100, 
       u1_u10_u5_n101, u1_u10_u5_n102, u1_u10_u5_n103, u1_u10_u5_n104, u1_u10_u5_n105, u1_u10_u5_n106, u1_u10_u5_n107, u1_u10_u5_n108, u1_u10_u5_n109, 
       u1_u10_u5_n110, u1_u10_u5_n111, u1_u10_u5_n112, u1_u10_u5_n113, u1_u10_u5_n114, u1_u10_u5_n115, u1_u10_u5_n116, u1_u10_u5_n117, u1_u10_u5_n118, 
       u1_u10_u5_n119, u1_u10_u5_n120, u1_u10_u5_n121, u1_u10_u5_n122, u1_u10_u5_n123, u1_u10_u5_n124, u1_u10_u5_n125, u1_u10_u5_n126, u1_u10_u5_n127, 
       u1_u10_u5_n128, u1_u10_u5_n129, u1_u10_u5_n130, u1_u10_u5_n131, u1_u10_u5_n132, u1_u10_u5_n133, u1_u10_u5_n134, u1_u10_u5_n135, u1_u10_u5_n136, 
       u1_u10_u5_n137, u1_u10_u5_n138, u1_u10_u5_n139, u1_u10_u5_n140, u1_u10_u5_n141, u1_u10_u5_n142, u1_u10_u5_n143, u1_u10_u5_n144, u1_u10_u5_n145, 
       u1_u10_u5_n146, u1_u10_u5_n147, u1_u10_u5_n148, u1_u10_u5_n149, u1_u10_u5_n150, u1_u10_u5_n151, u1_u10_u5_n152, u1_u10_u5_n153, u1_u10_u5_n154, 
       u1_u10_u5_n155, u1_u10_u5_n156, u1_u10_u5_n157, u1_u10_u5_n158, u1_u10_u5_n159, u1_u10_u5_n160, u1_u10_u5_n161, u1_u10_u5_n162, u1_u10_u5_n163, 
       u1_u10_u5_n164, u1_u10_u5_n165, u1_u10_u5_n166, u1_u10_u5_n167, u1_u10_u5_n168, u1_u10_u5_n169, u1_u10_u5_n170, u1_u10_u5_n171, u1_u10_u5_n172, 
       u1_u10_u5_n173, u1_u10_u5_n174, u1_u10_u5_n175, u1_u10_u5_n176, u1_u10_u5_n177, u1_u10_u5_n178, u1_u10_u5_n179, u1_u10_u5_n180, u1_u10_u5_n181, 
       u1_u10_u5_n182, u1_u10_u5_n183, u1_u10_u5_n184, u1_u10_u5_n185, u1_u10_u5_n186, u1_u10_u5_n187, u1_u10_u5_n188, u1_u10_u5_n189, u1_u10_u5_n190, 
       u1_u10_u5_n191, u1_u10_u5_n192, u1_u10_u5_n193, u1_u10_u5_n194, u1_u10_u5_n195, u1_u10_u5_n196, u1_u10_u5_n99, u1_u10_u6_n100, u1_u10_u6_n101, 
       u1_u10_u6_n102, u1_u10_u6_n103, u1_u10_u6_n104, u1_u10_u6_n105, u1_u10_u6_n106, u1_u10_u6_n107, u1_u10_u6_n108, u1_u10_u6_n109, u1_u10_u6_n110, 
       u1_u10_u6_n111, u1_u10_u6_n112, u1_u10_u6_n113, u1_u10_u6_n114, u1_u10_u6_n115, u1_u10_u6_n116, u1_u10_u6_n117, u1_u10_u6_n118, u1_u10_u6_n119, 
       u1_u10_u6_n120, u1_u10_u6_n121, u1_u10_u6_n122, u1_u10_u6_n123, u1_u10_u6_n124, u1_u10_u6_n125, u1_u10_u6_n126, u1_u10_u6_n127, u1_u10_u6_n128, 
       u1_u10_u6_n129, u1_u10_u6_n130, u1_u10_u6_n131, u1_u10_u6_n132, u1_u10_u6_n133, u1_u10_u6_n134, u1_u10_u6_n135, u1_u10_u6_n136, u1_u10_u6_n137, 
       u1_u10_u6_n138, u1_u10_u6_n139, u1_u10_u6_n140, u1_u10_u6_n141, u1_u10_u6_n142, u1_u10_u6_n143, u1_u10_u6_n144, u1_u10_u6_n145, u1_u10_u6_n146, 
       u1_u10_u6_n147, u1_u10_u6_n148, u1_u10_u6_n149, u1_u10_u6_n150, u1_u10_u6_n151, u1_u10_u6_n152, u1_u10_u6_n153, u1_u10_u6_n154, u1_u10_u6_n155, 
       u1_u10_u6_n156, u1_u10_u6_n157, u1_u10_u6_n158, u1_u10_u6_n159, u1_u10_u6_n160, u1_u10_u6_n161, u1_u10_u6_n162, u1_u10_u6_n163, u1_u10_u6_n164, 
       u1_u10_u6_n165, u1_u10_u6_n166, u1_u10_u6_n167, u1_u10_u6_n168, u1_u10_u6_n169, u1_u10_u6_n170, u1_u10_u6_n171, u1_u10_u6_n172, u1_u10_u6_n173, 
       u1_u10_u6_n174, u1_u10_u6_n88, u1_u10_u6_n89, u1_u10_u6_n90, u1_u10_u6_n91, u1_u10_u6_n92, u1_u10_u6_n93, u1_u10_u6_n94, u1_u10_u6_n95, 
       u1_u10_u6_n96, u1_u10_u6_n97, u1_u10_u6_n98, u1_u10_u6_n99, u1_u10_u7_n100, u1_u10_u7_n101, u1_u10_u7_n102, u1_u10_u7_n103, u1_u10_u7_n104, 
       u1_u10_u7_n105, u1_u10_u7_n106, u1_u10_u7_n107, u1_u10_u7_n108, u1_u10_u7_n109, u1_u10_u7_n110, u1_u10_u7_n111, u1_u10_u7_n112, u1_u10_u7_n113, 
       u1_u10_u7_n114, u1_u10_u7_n115, u1_u10_u7_n116, u1_u10_u7_n117, u1_u10_u7_n118, u1_u10_u7_n119, u1_u10_u7_n120, u1_u10_u7_n121, u1_u10_u7_n122, 
       u1_u10_u7_n123, u1_u10_u7_n124, u1_u10_u7_n125, u1_u10_u7_n126, u1_u10_u7_n127, u1_u10_u7_n128, u1_u10_u7_n129, u1_u10_u7_n130, u1_u10_u7_n131, 
       u1_u10_u7_n132, u1_u10_u7_n133, u1_u10_u7_n134, u1_u10_u7_n135, u1_u10_u7_n136, u1_u10_u7_n137, u1_u10_u7_n138, u1_u10_u7_n139, u1_u10_u7_n140, 
       u1_u10_u7_n141, u1_u10_u7_n142, u1_u10_u7_n143, u1_u10_u7_n144, u1_u10_u7_n145, u1_u10_u7_n146, u1_u10_u7_n147, u1_u10_u7_n148, u1_u10_u7_n149, 
       u1_u10_u7_n150, u1_u10_u7_n151, u1_u10_u7_n152, u1_u10_u7_n153, u1_u10_u7_n154, u1_u10_u7_n155, u1_u10_u7_n156, u1_u10_u7_n157, u1_u10_u7_n158, 
       u1_u10_u7_n159, u1_u10_u7_n160, u1_u10_u7_n161, u1_u10_u7_n162, u1_u10_u7_n163, u1_u10_u7_n164, u1_u10_u7_n165, u1_u10_u7_n166, u1_u10_u7_n167, 
       u1_u10_u7_n168, u1_u10_u7_n169, u1_u10_u7_n170, u1_u10_u7_n171, u1_u10_u7_n172, u1_u10_u7_n173, u1_u10_u7_n174, u1_u10_u7_n175, u1_u10_u7_n176, 
       u1_u10_u7_n177, u1_u10_u7_n178, u1_u10_u7_n179, u1_u10_u7_n180, u1_u10_u7_n91, u1_u10_u7_n92, u1_u10_u7_n93, u1_u10_u7_n94, u1_u10_u7_n95, 
       u1_u10_u7_n96, u1_u10_u7_n97, u1_u10_u7_n98, u1_u10_u7_n99, u1_u12_X_11, u1_u12_X_12, u1_u12_X_13, u1_u12_X_14, u1_u12_X_15, 
       u1_u12_X_17, u1_u12_X_18, u1_u12_X_19, u1_u12_X_2, u1_u12_X_20, u1_u12_X_48, u1_u12_X_5, u1_u12_X_6, u1_u12_X_7, 
       u1_u12_X_8, u1_u12_u0_n100, u1_u12_u0_n101, u1_u12_u0_n102, u1_u12_u0_n103, u1_u12_u0_n104, u1_u12_u0_n105, u1_u12_u0_n106, u1_u12_u0_n107, 
       u1_u12_u0_n108, u1_u12_u0_n109, u1_u12_u0_n110, u1_u12_u0_n111, u1_u12_u0_n112, u1_u12_u0_n113, u1_u12_u0_n114, u1_u12_u0_n115, u1_u12_u0_n116, 
       u1_u12_u0_n117, u1_u12_u0_n118, u1_u12_u0_n119, u1_u12_u0_n120, u1_u12_u0_n121, u1_u12_u0_n122, u1_u12_u0_n123, u1_u12_u0_n124, u1_u12_u0_n125, 
       u1_u12_u0_n126, u1_u12_u0_n127, u1_u12_u0_n128, u1_u12_u0_n129, u1_u12_u0_n130, u1_u12_u0_n131, u1_u12_u0_n132, u1_u12_u0_n133, u1_u12_u0_n134, 
       u1_u12_u0_n135, u1_u12_u0_n136, u1_u12_u0_n137, u1_u12_u0_n138, u1_u12_u0_n139, u1_u12_u0_n140, u1_u12_u0_n141, u1_u12_u0_n142, u1_u12_u0_n143, 
       u1_u12_u0_n144, u1_u12_u0_n145, u1_u12_u0_n146, u1_u12_u0_n147, u1_u12_u0_n148, u1_u12_u0_n149, u1_u12_u0_n150, u1_u12_u0_n151, u1_u12_u0_n152, 
       u1_u12_u0_n153, u1_u12_u0_n154, u1_u12_u0_n155, u1_u12_u0_n156, u1_u12_u0_n157, u1_u12_u0_n158, u1_u12_u0_n159, u1_u12_u0_n160, u1_u12_u0_n161, 
       u1_u12_u0_n162, u1_u12_u0_n163, u1_u12_u0_n164, u1_u12_u0_n165, u1_u12_u0_n166, u1_u12_u0_n167, u1_u12_u0_n168, u1_u12_u0_n169, u1_u12_u0_n170, 
       u1_u12_u0_n171, u1_u12_u0_n172, u1_u12_u0_n173, u1_u12_u0_n174, u1_u12_u0_n88, u1_u12_u0_n89, u1_u12_u0_n90, u1_u12_u0_n91, u1_u12_u0_n92, 
       u1_u12_u0_n93, u1_u12_u0_n94, u1_u12_u0_n95, u1_u12_u0_n96, u1_u12_u0_n97, u1_u12_u0_n98, u1_u12_u0_n99, u1_u12_u1_n100, u1_u12_u1_n101, 
       u1_u12_u1_n102, u1_u12_u1_n103, u1_u12_u1_n104, u1_u12_u1_n105, u1_u12_u1_n106, u1_u12_u1_n107, u1_u12_u1_n108, u1_u12_u1_n109, u1_u12_u1_n110, 
       u1_u12_u1_n111, u1_u12_u1_n112, u1_u12_u1_n113, u1_u12_u1_n114, u1_u12_u1_n115, u1_u12_u1_n116, u1_u12_u1_n117, u1_u12_u1_n118, u1_u12_u1_n119, 
       u1_u12_u1_n120, u1_u12_u1_n121, u1_u12_u1_n122, u1_u12_u1_n123, u1_u12_u1_n124, u1_u12_u1_n125, u1_u12_u1_n126, u1_u12_u1_n127, u1_u12_u1_n128, 
       u1_u12_u1_n129, u1_u12_u1_n130, u1_u12_u1_n131, u1_u12_u1_n132, u1_u12_u1_n133, u1_u12_u1_n134, u1_u12_u1_n135, u1_u12_u1_n136, u1_u12_u1_n137, 
       u1_u12_u1_n138, u1_u12_u1_n139, u1_u12_u1_n140, u1_u12_u1_n141, u1_u12_u1_n142, u1_u12_u1_n143, u1_u12_u1_n144, u1_u12_u1_n145, u1_u12_u1_n146, 
       u1_u12_u1_n147, u1_u12_u1_n148, u1_u12_u1_n149, u1_u12_u1_n150, u1_u12_u1_n151, u1_u12_u1_n152, u1_u12_u1_n153, u1_u12_u1_n154, u1_u12_u1_n155, 
       u1_u12_u1_n156, u1_u12_u1_n157, u1_u12_u1_n158, u1_u12_u1_n159, u1_u12_u1_n160, u1_u12_u1_n161, u1_u12_u1_n162, u1_u12_u1_n163, u1_u12_u1_n164, 
       u1_u12_u1_n165, u1_u12_u1_n166, u1_u12_u1_n167, u1_u12_u1_n168, u1_u12_u1_n169, u1_u12_u1_n170, u1_u12_u1_n171, u1_u12_u1_n172, u1_u12_u1_n173, 
       u1_u12_u1_n174, u1_u12_u1_n175, u1_u12_u1_n176, u1_u12_u1_n177, u1_u12_u1_n178, u1_u12_u1_n179, u1_u12_u1_n180, u1_u12_u1_n181, u1_u12_u1_n182, 
       u1_u12_u1_n183, u1_u12_u1_n184, u1_u12_u1_n185, u1_u12_u1_n186, u1_u12_u1_n187, u1_u12_u1_n188, u1_u12_u1_n95, u1_u12_u1_n96, u1_u12_u1_n97, 
       u1_u12_u1_n98, u1_u12_u1_n99, u1_u12_u2_n100, u1_u12_u2_n101, u1_u12_u2_n102, u1_u12_u2_n103, u1_u12_u2_n104, u1_u12_u2_n105, u1_u12_u2_n106, 
       u1_u12_u2_n107, u1_u12_u2_n108, u1_u12_u2_n109, u1_u12_u2_n110, u1_u12_u2_n111, u1_u12_u2_n112, u1_u12_u2_n113, u1_u12_u2_n114, u1_u12_u2_n115, 
       u1_u12_u2_n116, u1_u12_u2_n117, u1_u12_u2_n118, u1_u12_u2_n119, u1_u12_u2_n120, u1_u12_u2_n121, u1_u12_u2_n122, u1_u12_u2_n123, u1_u12_u2_n124, 
       u1_u12_u2_n125, u1_u12_u2_n126, u1_u12_u2_n127, u1_u12_u2_n128, u1_u12_u2_n129, u1_u12_u2_n130, u1_u12_u2_n131, u1_u12_u2_n132, u1_u12_u2_n133, 
       u1_u12_u2_n134, u1_u12_u2_n135, u1_u12_u2_n136, u1_u12_u2_n137, u1_u12_u2_n138, u1_u12_u2_n139, u1_u12_u2_n140, u1_u12_u2_n141, u1_u12_u2_n142, 
       u1_u12_u2_n143, u1_u12_u2_n144, u1_u12_u2_n145, u1_u12_u2_n146, u1_u12_u2_n147, u1_u12_u2_n148, u1_u12_u2_n149, u1_u12_u2_n150, u1_u12_u2_n151, 
       u1_u12_u2_n152, u1_u12_u2_n153, u1_u12_u2_n154, u1_u12_u2_n155, u1_u12_u2_n156, u1_u12_u2_n157, u1_u12_u2_n158, u1_u12_u2_n159, u1_u12_u2_n160, 
       u1_u12_u2_n161, u1_u12_u2_n162, u1_u12_u2_n163, u1_u12_u2_n164, u1_u12_u2_n165, u1_u12_u2_n166, u1_u12_u2_n167, u1_u12_u2_n168, u1_u12_u2_n169, 
       u1_u12_u2_n170, u1_u12_u2_n171, u1_u12_u2_n172, u1_u12_u2_n173, u1_u12_u2_n174, u1_u12_u2_n175, u1_u12_u2_n176, u1_u12_u2_n177, u1_u12_u2_n178, 
       u1_u12_u2_n179, u1_u12_u2_n180, u1_u12_u2_n181, u1_u12_u2_n182, u1_u12_u2_n183, u1_u12_u2_n184, u1_u12_u2_n185, u1_u12_u2_n186, u1_u12_u2_n187, 
       u1_u12_u2_n188, u1_u12_u2_n95, u1_u12_u2_n96, u1_u12_u2_n97, u1_u12_u2_n98, u1_u12_u2_n99, u1_u12_u3_n100, u1_u12_u3_n101, u1_u12_u3_n102, 
       u1_u12_u3_n103, u1_u12_u3_n104, u1_u12_u3_n105, u1_u12_u3_n106, u1_u12_u3_n107, u1_u12_u3_n108, u1_u12_u3_n109, u1_u12_u3_n110, u1_u12_u3_n111, 
       u1_u12_u3_n112, u1_u12_u3_n113, u1_u12_u3_n114, u1_u12_u3_n115, u1_u12_u3_n116, u1_u12_u3_n117, u1_u12_u3_n118, u1_u12_u3_n119, u1_u12_u3_n120, 
       u1_u12_u3_n121, u1_u12_u3_n122, u1_u12_u3_n123, u1_u12_u3_n124, u1_u12_u3_n125, u1_u12_u3_n126, u1_u12_u3_n127, u1_u12_u3_n128, u1_u12_u3_n129, 
       u1_u12_u3_n130, u1_u12_u3_n131, u1_u12_u3_n132, u1_u12_u3_n133, u1_u12_u3_n134, u1_u12_u3_n135, u1_u12_u3_n136, u1_u12_u3_n137, u1_u12_u3_n138, 
       u1_u12_u3_n139, u1_u12_u3_n140, u1_u12_u3_n141, u1_u12_u3_n142, u1_u12_u3_n143, u1_u12_u3_n144, u1_u12_u3_n145, u1_u12_u3_n146, u1_u12_u3_n147, 
       u1_u12_u3_n148, u1_u12_u3_n149, u1_u12_u3_n150, u1_u12_u3_n151, u1_u12_u3_n152, u1_u12_u3_n153, u1_u12_u3_n154, u1_u12_u3_n155, u1_u12_u3_n156, 
       u1_u12_u3_n157, u1_u12_u3_n158, u1_u12_u3_n159, u1_u12_u3_n160, u1_u12_u3_n161, u1_u12_u3_n162, u1_u12_u3_n163, u1_u12_u3_n164, u1_u12_u3_n165, 
       u1_u12_u3_n166, u1_u12_u3_n167, u1_u12_u3_n168, u1_u12_u3_n169, u1_u12_u3_n170, u1_u12_u3_n171, u1_u12_u3_n172, u1_u12_u3_n173, u1_u12_u3_n174, 
       u1_u12_u3_n175, u1_u12_u3_n176, u1_u12_u3_n177, u1_u12_u3_n178, u1_u12_u3_n179, u1_u12_u3_n180, u1_u12_u3_n181, u1_u12_u3_n182, u1_u12_u3_n183, 
       u1_u12_u3_n184, u1_u12_u3_n185, u1_u12_u3_n186, u1_u12_u3_n94, u1_u12_u3_n95, u1_u12_u3_n96, u1_u12_u3_n97, u1_u12_u3_n98, u1_u12_u3_n99, 
       u1_u12_u7_n100, u1_u12_u7_n101, u1_u12_u7_n102, u1_u12_u7_n103, u1_u12_u7_n104, u1_u12_u7_n105, u1_u12_u7_n106, u1_u12_u7_n107, u1_u12_u7_n108, 
       u1_u12_u7_n109, u1_u12_u7_n110, u1_u12_u7_n111, u1_u12_u7_n112, u1_u12_u7_n113, u1_u12_u7_n114, u1_u12_u7_n115, u1_u12_u7_n116, u1_u12_u7_n117, 
       u1_u12_u7_n118, u1_u12_u7_n119, u1_u12_u7_n120, u1_u12_u7_n121, u1_u12_u7_n122, u1_u12_u7_n123, u1_u12_u7_n124, u1_u12_u7_n125, u1_u12_u7_n126, 
       u1_u12_u7_n127, u1_u12_u7_n128, u1_u12_u7_n129, u1_u12_u7_n130, u1_u12_u7_n131, u1_u12_u7_n132, u1_u12_u7_n133, u1_u12_u7_n134, u1_u12_u7_n135, 
       u1_u12_u7_n136, u1_u12_u7_n137, u1_u12_u7_n138, u1_u12_u7_n139, u1_u12_u7_n140, u1_u12_u7_n141, u1_u12_u7_n142, u1_u12_u7_n143, u1_u12_u7_n144, 
       u1_u12_u7_n145, u1_u12_u7_n146, u1_u12_u7_n147, u1_u12_u7_n148, u1_u12_u7_n149, u1_u12_u7_n150, u1_u12_u7_n151, u1_u12_u7_n152, u1_u12_u7_n153, 
       u1_u12_u7_n154, u1_u12_u7_n155, u1_u12_u7_n156, u1_u12_u7_n157, u1_u12_u7_n158, u1_u12_u7_n159, u1_u12_u7_n160, u1_u12_u7_n161, u1_u12_u7_n162, 
       u1_u12_u7_n163, u1_u12_u7_n164, u1_u12_u7_n165, u1_u12_u7_n166, u1_u12_u7_n167, u1_u12_u7_n168, u1_u12_u7_n169, u1_u12_u7_n170, u1_u12_u7_n171, 
       u1_u12_u7_n172, u1_u12_u7_n173, u1_u12_u7_n174, u1_u12_u7_n175, u1_u12_u7_n176, u1_u12_u7_n177, u1_u12_u7_n178, u1_u12_u7_n179, u1_u12_u7_n180, 
       u1_u12_u7_n91, u1_u12_u7_n92, u1_u12_u7_n93, u1_u12_u7_n94, u1_u12_u7_n95, u1_u12_u7_n96, u1_u12_u7_n97, u1_u12_u7_n98, u1_u12_u7_n99, 
       u1_u13_X_1, u1_u13_X_2, u1_u13_X_42, u1_u13_X_44, u1_u13_X_47, u1_u13_X_48, u1_u13_u0_n100, u1_u13_u0_n101, u1_u13_u0_n102, 
       u1_u13_u0_n103, u1_u13_u0_n104, u1_u13_u0_n105, u1_u13_u0_n106, u1_u13_u0_n107, u1_u13_u0_n108, u1_u13_u0_n109, u1_u13_u0_n110, u1_u13_u0_n111, 
       u1_u13_u0_n112, u1_u13_u0_n113, u1_u13_u0_n114, u1_u13_u0_n115, u1_u13_u0_n116, u1_u13_u0_n117, u1_u13_u0_n118, u1_u13_u0_n119, u1_u13_u0_n120, 
       u1_u13_u0_n121, u1_u13_u0_n122, u1_u13_u0_n123, u1_u13_u0_n124, u1_u13_u0_n125, u1_u13_u0_n126, u1_u13_u0_n127, u1_u13_u0_n128, u1_u13_u0_n129, 
       u1_u13_u0_n130, u1_u13_u0_n131, u1_u13_u0_n132, u1_u13_u0_n133, u1_u13_u0_n134, u1_u13_u0_n135, u1_u13_u0_n136, u1_u13_u0_n137, u1_u13_u0_n138, 
       u1_u13_u0_n139, u1_u13_u0_n140, u1_u13_u0_n141, u1_u13_u0_n142, u1_u13_u0_n143, u1_u13_u0_n144, u1_u13_u0_n145, u1_u13_u0_n146, u1_u13_u0_n147, 
       u1_u13_u0_n148, u1_u13_u0_n149, u1_u13_u0_n150, u1_u13_u0_n151, u1_u13_u0_n152, u1_u13_u0_n153, u1_u13_u0_n154, u1_u13_u0_n155, u1_u13_u0_n156, 
       u1_u13_u0_n157, u1_u13_u0_n158, u1_u13_u0_n159, u1_u13_u0_n160, u1_u13_u0_n161, u1_u13_u0_n162, u1_u13_u0_n163, u1_u13_u0_n164, u1_u13_u0_n165, 
       u1_u13_u0_n166, u1_u13_u0_n167, u1_u13_u0_n168, u1_u13_u0_n169, u1_u13_u0_n170, u1_u13_u0_n171, u1_u13_u0_n172, u1_u13_u0_n173, u1_u13_u0_n174, 
       u1_u13_u0_n88, u1_u13_u0_n89, u1_u13_u0_n90, u1_u13_u0_n91, u1_u13_u0_n92, u1_u13_u0_n93, u1_u13_u0_n94, u1_u13_u0_n95, u1_u13_u0_n96, 
       u1_u13_u0_n97, u1_u13_u0_n98, u1_u13_u0_n99, u1_u13_u1_n100, u1_u13_u1_n101, u1_u13_u1_n102, u1_u13_u1_n103, u1_u13_u1_n104, u1_u13_u1_n105, 
       u1_u13_u1_n106, u1_u13_u1_n107, u1_u13_u1_n108, u1_u13_u1_n109, u1_u13_u1_n110, u1_u13_u1_n111, u1_u13_u1_n112, u1_u13_u1_n113, u1_u13_u1_n114, 
       u1_u13_u1_n115, u1_u13_u1_n116, u1_u13_u1_n117, u1_u13_u1_n118, u1_u13_u1_n119, u1_u13_u1_n120, u1_u13_u1_n121, u1_u13_u1_n122, u1_u13_u1_n123, 
       u1_u13_u1_n124, u1_u13_u1_n125, u1_u13_u1_n126, u1_u13_u1_n127, u1_u13_u1_n128, u1_u13_u1_n129, u1_u13_u1_n130, u1_u13_u1_n131, u1_u13_u1_n132, 
       u1_u13_u1_n133, u1_u13_u1_n134, u1_u13_u1_n135, u1_u13_u1_n136, u1_u13_u1_n137, u1_u13_u1_n138, u1_u13_u1_n139, u1_u13_u1_n140, u1_u13_u1_n141, 
       u1_u13_u1_n142, u1_u13_u1_n143, u1_u13_u1_n144, u1_u13_u1_n145, u1_u13_u1_n146, u1_u13_u1_n147, u1_u13_u1_n148, u1_u13_u1_n149, u1_u13_u1_n150, 
       u1_u13_u1_n151, u1_u13_u1_n152, u1_u13_u1_n153, u1_u13_u1_n154, u1_u13_u1_n155, u1_u13_u1_n156, u1_u13_u1_n157, u1_u13_u1_n158, u1_u13_u1_n159, 
       u1_u13_u1_n160, u1_u13_u1_n161, u1_u13_u1_n162, u1_u13_u1_n163, u1_u13_u1_n164, u1_u13_u1_n165, u1_u13_u1_n166, u1_u13_u1_n167, u1_u13_u1_n168, 
       u1_u13_u1_n169, u1_u13_u1_n170, u1_u13_u1_n171, u1_u13_u1_n172, u1_u13_u1_n173, u1_u13_u1_n174, u1_u13_u1_n175, u1_u13_u1_n176, u1_u13_u1_n177, 
       u1_u13_u1_n178, u1_u13_u1_n179, u1_u13_u1_n180, u1_u13_u1_n181, u1_u13_u1_n182, u1_u13_u1_n183, u1_u13_u1_n184, u1_u13_u1_n185, u1_u13_u1_n186, 
       u1_u13_u1_n187, u1_u13_u1_n188, u1_u13_u1_n95, u1_u13_u1_n96, u1_u13_u1_n97, u1_u13_u1_n98, u1_u13_u1_n99, u1_u13_u6_n100, u1_u13_u6_n101, 
       u1_u13_u6_n102, u1_u13_u6_n103, u1_u13_u6_n104, u1_u13_u6_n105, u1_u13_u6_n106, u1_u13_u6_n107, u1_u13_u6_n108, u1_u13_u6_n109, u1_u13_u6_n110, 
       u1_u13_u6_n111, u1_u13_u6_n112, u1_u13_u6_n113, u1_u13_u6_n114, u1_u13_u6_n115, u1_u13_u6_n116, u1_u13_u6_n117, u1_u13_u6_n118, u1_u13_u6_n119, 
       u1_u13_u6_n120, u1_u13_u6_n121, u1_u13_u6_n122, u1_u13_u6_n123, u1_u13_u6_n124, u1_u13_u6_n125, u1_u13_u6_n126, u1_u13_u6_n127, u1_u13_u6_n128, 
       u1_u13_u6_n129, u1_u13_u6_n130, u1_u13_u6_n131, u1_u13_u6_n132, u1_u13_u6_n133, u1_u13_u6_n134, u1_u13_u6_n135, u1_u13_u6_n136, u1_u13_u6_n137, 
       u1_u13_u6_n138, u1_u13_u6_n139, u1_u13_u6_n140, u1_u13_u6_n141, u1_u13_u6_n142, u1_u13_u6_n143, u1_u13_u6_n144, u1_u13_u6_n145, u1_u13_u6_n146, 
       u1_u13_u6_n147, u1_u13_u6_n148, u1_u13_u6_n149, u1_u13_u6_n150, u1_u13_u6_n151, u1_u13_u6_n152, u1_u13_u6_n153, u1_u13_u6_n154, u1_u13_u6_n155, 
       u1_u13_u6_n156, u1_u13_u6_n157, u1_u13_u6_n158, u1_u13_u6_n159, u1_u13_u6_n160, u1_u13_u6_n161, u1_u13_u6_n162, u1_u13_u6_n163, u1_u13_u6_n164, 
       u1_u13_u6_n165, u1_u13_u6_n166, u1_u13_u6_n167, u1_u13_u6_n168, u1_u13_u6_n169, u1_u13_u6_n170, u1_u13_u6_n171, u1_u13_u6_n172, u1_u13_u6_n173, 
       u1_u13_u6_n174, u1_u13_u6_n88, u1_u13_u6_n89, u1_u13_u6_n90, u1_u13_u6_n91, u1_u13_u6_n92, u1_u13_u6_n93, u1_u13_u6_n94, u1_u13_u6_n95, 
       u1_u13_u6_n96, u1_u13_u6_n97, u1_u13_u6_n98, u1_u13_u6_n99, u1_u13_u7_n100, u1_u13_u7_n101, u1_u13_u7_n102, u1_u13_u7_n103, u1_u13_u7_n104, 
       u1_u13_u7_n105, u1_u13_u7_n106, u1_u13_u7_n107, u1_u13_u7_n108, u1_u13_u7_n109, u1_u13_u7_n110, u1_u13_u7_n111, u1_u13_u7_n112, u1_u13_u7_n113, 
       u1_u13_u7_n114, u1_u13_u7_n115, u1_u13_u7_n116, u1_u13_u7_n117, u1_u13_u7_n118, u1_u13_u7_n119, u1_u13_u7_n120, u1_u13_u7_n121, u1_u13_u7_n122, 
       u1_u13_u7_n123, u1_u13_u7_n124, u1_u13_u7_n125, u1_u13_u7_n126, u1_u13_u7_n127, u1_u13_u7_n128, u1_u13_u7_n129, u1_u13_u7_n130, u1_u13_u7_n131, 
       u1_u13_u7_n132, u1_u13_u7_n133, u1_u13_u7_n134, u1_u13_u7_n135, u1_u13_u7_n136, u1_u13_u7_n137, u1_u13_u7_n138, u1_u13_u7_n139, u1_u13_u7_n140, 
       u1_u13_u7_n141, u1_u13_u7_n142, u1_u13_u7_n143, u1_u13_u7_n144, u1_u13_u7_n145, u1_u13_u7_n146, u1_u13_u7_n147, u1_u13_u7_n148, u1_u13_u7_n149, 
       u1_u13_u7_n150, u1_u13_u7_n151, u1_u13_u7_n152, u1_u13_u7_n153, u1_u13_u7_n154, u1_u13_u7_n155, u1_u13_u7_n156, u1_u13_u7_n157, u1_u13_u7_n158, 
       u1_u13_u7_n159, u1_u13_u7_n160, u1_u13_u7_n161, u1_u13_u7_n162, u1_u13_u7_n163, u1_u13_u7_n164, u1_u13_u7_n165, u1_u13_u7_n166, u1_u13_u7_n167, 
       u1_u13_u7_n168, u1_u13_u7_n169, u1_u13_u7_n170, u1_u13_u7_n171, u1_u13_u7_n172, u1_u13_u7_n173, u1_u13_u7_n174, u1_u13_u7_n175, u1_u13_u7_n176, 
       u1_u13_u7_n177, u1_u13_u7_n178, u1_u13_u7_n179, u1_u13_u7_n180, u1_u13_u7_n91, u1_u13_u7_n92, u1_u13_u7_n93, u1_u13_u7_n94, u1_u13_u7_n95, 
       u1_u13_u7_n96, u1_u13_u7_n97, u1_u13_u7_n98, u1_u13_u7_n99, u1_u14_X_11, u1_u14_X_12, u1_u14_X_13, u1_u14_X_14, u1_u14_X_18, 
       u1_u14_X_2, u1_u14_X_20, u1_u14_X_23, u1_u14_X_24, u1_u14_X_25, u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u14_X_31, 
       u1_u14_X_32, u1_u14_X_35, u1_u14_X_36, u1_u14_X_37, u1_u14_X_38, u1_u14_X_41, u1_u14_X_42, u1_u14_X_43, u1_u14_X_44, 
       u1_u14_X_48, u1_u14_X_5, u1_u14_X_6, u1_u14_X_7, u1_u14_X_8, u1_u14_u0_n100, u1_u14_u0_n101, u1_u14_u0_n102, u1_u14_u0_n103, 
       u1_u14_u0_n104, u1_u14_u0_n105, u1_u14_u0_n106, u1_u14_u0_n107, u1_u14_u0_n108, u1_u14_u0_n109, u1_u14_u0_n110, u1_u14_u0_n111, u1_u14_u0_n112, 
       u1_u14_u0_n113, u1_u14_u0_n114, u1_u14_u0_n115, u1_u14_u0_n116, u1_u14_u0_n117, u1_u14_u0_n118, u1_u14_u0_n119, u1_u14_u0_n120, u1_u14_u0_n121, 
       u1_u14_u0_n122, u1_u14_u0_n123, u1_u14_u0_n124, u1_u14_u0_n125, u1_u14_u0_n126, u1_u14_u0_n127, u1_u14_u0_n128, u1_u14_u0_n129, u1_u14_u0_n130, 
       u1_u14_u0_n131, u1_u14_u0_n132, u1_u14_u0_n133, u1_u14_u0_n134, u1_u14_u0_n135, u1_u14_u0_n136, u1_u14_u0_n137, u1_u14_u0_n138, u1_u14_u0_n139, 
       u1_u14_u0_n140, u1_u14_u0_n141, u1_u14_u0_n142, u1_u14_u0_n143, u1_u14_u0_n144, u1_u14_u0_n145, u1_u14_u0_n146, u1_u14_u0_n147, u1_u14_u0_n148, 
       u1_u14_u0_n149, u1_u14_u0_n150, u1_u14_u0_n151, u1_u14_u0_n152, u1_u14_u0_n153, u1_u14_u0_n154, u1_u14_u0_n155, u1_u14_u0_n156, u1_u14_u0_n157, 
       u1_u14_u0_n158, u1_u14_u0_n159, u1_u14_u0_n160, u1_u14_u0_n161, u1_u14_u0_n162, u1_u14_u0_n163, u1_u14_u0_n164, u1_u14_u0_n165, u1_u14_u0_n166, 
       u1_u14_u0_n167, u1_u14_u0_n168, u1_u14_u0_n169, u1_u14_u0_n170, u1_u14_u0_n171, u1_u14_u0_n172, u1_u14_u0_n173, u1_u14_u0_n174, u1_u14_u0_n88, 
       u1_u14_u0_n89, u1_u14_u0_n90, u1_u14_u0_n91, u1_u14_u0_n92, u1_u14_u0_n93, u1_u14_u0_n94, u1_u14_u0_n95, u1_u14_u0_n96, u1_u14_u0_n97, 
       u1_u14_u0_n98, u1_u14_u0_n99, u1_u14_u1_n100, u1_u14_u1_n101, u1_u14_u1_n102, u1_u14_u1_n103, u1_u14_u1_n104, u1_u14_u1_n105, u1_u14_u1_n106, 
       u1_u14_u1_n107, u1_u14_u1_n108, u1_u14_u1_n109, u1_u14_u1_n110, u1_u14_u1_n111, u1_u14_u1_n112, u1_u14_u1_n113, u1_u14_u1_n114, u1_u14_u1_n115, 
       u1_u14_u1_n116, u1_u14_u1_n117, u1_u14_u1_n118, u1_u14_u1_n119, u1_u14_u1_n120, u1_u14_u1_n121, u1_u14_u1_n122, u1_u14_u1_n123, u1_u14_u1_n124, 
       u1_u14_u1_n125, u1_u14_u1_n126, u1_u14_u1_n127, u1_u14_u1_n128, u1_u14_u1_n129, u1_u14_u1_n130, u1_u14_u1_n131, u1_u14_u1_n132, u1_u14_u1_n133, 
       u1_u14_u1_n134, u1_u14_u1_n135, u1_u14_u1_n136, u1_u14_u1_n137, u1_u14_u1_n138, u1_u14_u1_n139, u1_u14_u1_n140, u1_u14_u1_n141, u1_u14_u1_n142, 
       u1_u14_u1_n143, u1_u14_u1_n144, u1_u14_u1_n145, u1_u14_u1_n146, u1_u14_u1_n147, u1_u14_u1_n148, u1_u14_u1_n149, u1_u14_u1_n150, u1_u14_u1_n151, 
       u1_u14_u1_n152, u1_u14_u1_n153, u1_u14_u1_n154, u1_u14_u1_n155, u1_u14_u1_n156, u1_u14_u1_n157, u1_u14_u1_n158, u1_u14_u1_n159, u1_u14_u1_n160, 
       u1_u14_u1_n161, u1_u14_u1_n162, u1_u14_u1_n163, u1_u14_u1_n164, u1_u14_u1_n165, u1_u14_u1_n166, u1_u14_u1_n167, u1_u14_u1_n168, u1_u14_u1_n169, 
       u1_u14_u1_n170, u1_u14_u1_n171, u1_u14_u1_n172, u1_u14_u1_n173, u1_u14_u1_n174, u1_u14_u1_n175, u1_u14_u1_n176, u1_u14_u1_n177, u1_u14_u1_n178, 
       u1_u14_u1_n179, u1_u14_u1_n180, u1_u14_u1_n181, u1_u14_u1_n182, u1_u14_u1_n183, u1_u14_u1_n184, u1_u14_u1_n185, u1_u14_u1_n186, u1_u14_u1_n187, 
       u1_u14_u1_n188, u1_u14_u1_n95, u1_u14_u1_n96, u1_u14_u1_n97, u1_u14_u1_n98, u1_u14_u1_n99, u1_u14_u2_n100, u1_u14_u2_n101, u1_u14_u2_n102, 
       u1_u14_u2_n103, u1_u14_u2_n104, u1_u14_u2_n105, u1_u14_u2_n106, u1_u14_u2_n107, u1_u14_u2_n108, u1_u14_u2_n109, u1_u14_u2_n110, u1_u14_u2_n111, 
       u1_u14_u2_n112, u1_u14_u2_n113, u1_u14_u2_n114, u1_u14_u2_n115, u1_u14_u2_n116, u1_u14_u2_n117, u1_u14_u2_n118, u1_u14_u2_n119, u1_u14_u2_n120, 
       u1_u14_u2_n121, u1_u14_u2_n122, u1_u14_u2_n123, u1_u14_u2_n124, u1_u14_u2_n125, u1_u14_u2_n126, u1_u14_u2_n127, u1_u14_u2_n128, u1_u14_u2_n129, 
       u1_u14_u2_n130, u1_u14_u2_n131, u1_u14_u2_n132, u1_u14_u2_n133, u1_u14_u2_n134, u1_u14_u2_n135, u1_u14_u2_n136, u1_u14_u2_n137, u1_u14_u2_n138, 
       u1_u14_u2_n139, u1_u14_u2_n140, u1_u14_u2_n141, u1_u14_u2_n142, u1_u14_u2_n143, u1_u14_u2_n144, u1_u14_u2_n145, u1_u14_u2_n146, u1_u14_u2_n147, 
       u1_u14_u2_n148, u1_u14_u2_n149, u1_u14_u2_n150, u1_u14_u2_n151, u1_u14_u2_n152, u1_u14_u2_n153, u1_u14_u2_n154, u1_u14_u2_n155, u1_u14_u2_n156, 
       u1_u14_u2_n157, u1_u14_u2_n158, u1_u14_u2_n159, u1_u14_u2_n160, u1_u14_u2_n161, u1_u14_u2_n162, u1_u14_u2_n163, u1_u14_u2_n164, u1_u14_u2_n165, 
       u1_u14_u2_n166, u1_u14_u2_n167, u1_u14_u2_n168, u1_u14_u2_n169, u1_u14_u2_n170, u1_u14_u2_n171, u1_u14_u2_n172, u1_u14_u2_n173, u1_u14_u2_n174, 
       u1_u14_u2_n175, u1_u14_u2_n176, u1_u14_u2_n177, u1_u14_u2_n178, u1_u14_u2_n179, u1_u14_u2_n180, u1_u14_u2_n181, u1_u14_u2_n182, u1_u14_u2_n183, 
       u1_u14_u2_n184, u1_u14_u2_n185, u1_u14_u2_n186, u1_u14_u2_n187, u1_u14_u2_n188, u1_u14_u2_n95, u1_u14_u2_n96, u1_u14_u2_n97, u1_u14_u2_n98, 
       u1_u14_u2_n99, u1_u14_u3_n100, u1_u14_u3_n101, u1_u14_u3_n102, u1_u14_u3_n103, u1_u14_u3_n104, u1_u14_u3_n105, u1_u14_u3_n106, u1_u14_u3_n107, 
       u1_u14_u3_n108, u1_u14_u3_n109, u1_u14_u3_n110, u1_u14_u3_n111, u1_u14_u3_n112, u1_u14_u3_n113, u1_u14_u3_n114, u1_u14_u3_n115, u1_u14_u3_n116, 
       u1_u14_u3_n117, u1_u14_u3_n118, u1_u14_u3_n119, u1_u14_u3_n120, u1_u14_u3_n121, u1_u14_u3_n122, u1_u14_u3_n123, u1_u14_u3_n124, u1_u14_u3_n125, 
       u1_u14_u3_n126, u1_u14_u3_n127, u1_u14_u3_n128, u1_u14_u3_n129, u1_u14_u3_n130, u1_u14_u3_n131, u1_u14_u3_n132, u1_u14_u3_n133, u1_u14_u3_n134, 
       u1_u14_u3_n135, u1_u14_u3_n136, u1_u14_u3_n137, u1_u14_u3_n138, u1_u14_u3_n139, u1_u14_u3_n140, u1_u14_u3_n141, u1_u14_u3_n142, u1_u14_u3_n143, 
       u1_u14_u3_n144, u1_u14_u3_n145, u1_u14_u3_n146, u1_u14_u3_n147, u1_u14_u3_n148, u1_u14_u3_n149, u1_u14_u3_n150, u1_u14_u3_n151, u1_u14_u3_n152, 
       u1_u14_u3_n153, u1_u14_u3_n154, u1_u14_u3_n155, u1_u14_u3_n156, u1_u14_u3_n157, u1_u14_u3_n158, u1_u14_u3_n159, u1_u14_u3_n160, u1_u14_u3_n161, 
       u1_u14_u3_n162, u1_u14_u3_n163, u1_u14_u3_n164, u1_u14_u3_n165, u1_u14_u3_n166, u1_u14_u3_n167, u1_u14_u3_n168, u1_u14_u3_n169, u1_u14_u3_n170, 
       u1_u14_u3_n171, u1_u14_u3_n172, u1_u14_u3_n173, u1_u14_u3_n174, u1_u14_u3_n175, u1_u14_u3_n176, u1_u14_u3_n177, u1_u14_u3_n178, u1_u14_u3_n179, 
       u1_u14_u3_n180, u1_u14_u3_n181, u1_u14_u3_n182, u1_u14_u3_n183, u1_u14_u3_n184, u1_u14_u3_n185, u1_u14_u3_n186, u1_u14_u3_n94, u1_u14_u3_n95, 
       u1_u14_u3_n96, u1_u14_u3_n97, u1_u14_u3_n98, u1_u14_u3_n99, u1_u14_u4_n100, u1_u14_u4_n101, u1_u14_u4_n102, u1_u14_u4_n103, u1_u14_u4_n104, 
       u1_u14_u4_n105, u1_u14_u4_n106, u1_u14_u4_n107, u1_u14_u4_n108, u1_u14_u4_n109, u1_u14_u4_n110, u1_u14_u4_n111, u1_u14_u4_n112, u1_u14_u4_n113, 
       u1_u14_u4_n114, u1_u14_u4_n115, u1_u14_u4_n116, u1_u14_u4_n117, u1_u14_u4_n118, u1_u14_u4_n119, u1_u14_u4_n120, u1_u14_u4_n121, u1_u14_u4_n122, 
       u1_u14_u4_n123, u1_u14_u4_n124, u1_u14_u4_n125, u1_u14_u4_n126, u1_u14_u4_n127, u1_u14_u4_n128, u1_u14_u4_n129, u1_u14_u4_n130, u1_u14_u4_n131, 
       u1_u14_u4_n132, u1_u14_u4_n133, u1_u14_u4_n134, u1_u14_u4_n135, u1_u14_u4_n136, u1_u14_u4_n137, u1_u14_u4_n138, u1_u14_u4_n139, u1_u14_u4_n140, 
       u1_u14_u4_n141, u1_u14_u4_n142, u1_u14_u4_n143, u1_u14_u4_n144, u1_u14_u4_n145, u1_u14_u4_n146, u1_u14_u4_n147, u1_u14_u4_n148, u1_u14_u4_n149, 
       u1_u14_u4_n150, u1_u14_u4_n151, u1_u14_u4_n152, u1_u14_u4_n153, u1_u14_u4_n154, u1_u14_u4_n155, u1_u14_u4_n156, u1_u14_u4_n157, u1_u14_u4_n158, 
       u1_u14_u4_n159, u1_u14_u4_n160, u1_u14_u4_n161, u1_u14_u4_n162, u1_u14_u4_n163, u1_u14_u4_n164, u1_u14_u4_n165, u1_u14_u4_n166, u1_u14_u4_n167, 
       u1_u14_u4_n168, u1_u14_u4_n169, u1_u14_u4_n170, u1_u14_u4_n171, u1_u14_u4_n172, u1_u14_u4_n173, u1_u14_u4_n174, u1_u14_u4_n175, u1_u14_u4_n176, 
       u1_u14_u4_n177, u1_u14_u4_n178, u1_u14_u4_n179, u1_u14_u4_n180, u1_u14_u4_n181, u1_u14_u4_n182, u1_u14_u4_n183, u1_u14_u4_n184, u1_u14_u4_n185, 
       u1_u14_u4_n186, u1_u14_u4_n94, u1_u14_u4_n95, u1_u14_u4_n96, u1_u14_u4_n97, u1_u14_u4_n98, u1_u14_u4_n99, u1_u14_u5_n100, u1_u14_u5_n101, 
       u1_u14_u5_n102, u1_u14_u5_n103, u1_u14_u5_n104, u1_u14_u5_n105, u1_u14_u5_n106, u1_u14_u5_n107, u1_u14_u5_n108, u1_u14_u5_n109, u1_u14_u5_n110, 
       u1_u14_u5_n111, u1_u14_u5_n112, u1_u14_u5_n113, u1_u14_u5_n114, u1_u14_u5_n115, u1_u14_u5_n116, u1_u14_u5_n117, u1_u14_u5_n118, u1_u14_u5_n119, 
       u1_u14_u5_n120, u1_u14_u5_n121, u1_u14_u5_n122, u1_u14_u5_n123, u1_u14_u5_n124, u1_u14_u5_n125, u1_u14_u5_n126, u1_u14_u5_n127, u1_u14_u5_n128, 
       u1_u14_u5_n129, u1_u14_u5_n130, u1_u14_u5_n131, u1_u14_u5_n132, u1_u14_u5_n133, u1_u14_u5_n134, u1_u14_u5_n135, u1_u14_u5_n136, u1_u14_u5_n137, 
       u1_u14_u5_n138, u1_u14_u5_n139, u1_u14_u5_n140, u1_u14_u5_n141, u1_u14_u5_n142, u1_u14_u5_n143, u1_u14_u5_n144, u1_u14_u5_n145, u1_u14_u5_n146, 
       u1_u14_u5_n147, u1_u14_u5_n148, u1_u14_u5_n149, u1_u14_u5_n150, u1_u14_u5_n151, u1_u14_u5_n152, u1_u14_u5_n153, u1_u14_u5_n154, u1_u14_u5_n155, 
       u1_u14_u5_n156, u1_u14_u5_n157, u1_u14_u5_n158, u1_u14_u5_n159, u1_u14_u5_n160, u1_u14_u5_n161, u1_u14_u5_n162, u1_u14_u5_n163, u1_u14_u5_n164, 
       u1_u14_u5_n165, u1_u14_u5_n166, u1_u14_u5_n167, u1_u14_u5_n168, u1_u14_u5_n169, u1_u14_u5_n170, u1_u14_u5_n171, u1_u14_u5_n172, u1_u14_u5_n173, 
       u1_u14_u5_n174, u1_u14_u5_n175, u1_u14_u5_n176, u1_u14_u5_n177, u1_u14_u5_n178, u1_u14_u5_n179, u1_u14_u5_n180, u1_u14_u5_n181, u1_u14_u5_n182, 
       u1_u14_u5_n183, u1_u14_u5_n184, u1_u14_u5_n185, u1_u14_u5_n186, u1_u14_u5_n187, u1_u14_u5_n188, u1_u14_u5_n189, u1_u14_u5_n190, u1_u14_u5_n191, 
       u1_u14_u5_n192, u1_u14_u5_n193, u1_u14_u5_n194, u1_u14_u5_n195, u1_u14_u5_n196, u1_u14_u5_n99, u1_u14_u6_n100, u1_u14_u6_n101, u1_u14_u6_n102, 
       u1_u14_u6_n103, u1_u14_u6_n104, u1_u14_u6_n105, u1_u14_u6_n106, u1_u14_u6_n107, u1_u14_u6_n108, u1_u14_u6_n109, u1_u14_u6_n110, u1_u14_u6_n111, 
       u1_u14_u6_n112, u1_u14_u6_n113, u1_u14_u6_n114, u1_u14_u6_n115, u1_u14_u6_n116, u1_u14_u6_n117, u1_u14_u6_n118, u1_u14_u6_n119, u1_u14_u6_n120, 
       u1_u14_u6_n121, u1_u14_u6_n122, u1_u14_u6_n123, u1_u14_u6_n124, u1_u14_u6_n125, u1_u14_u6_n126, u1_u14_u6_n127, u1_u14_u6_n128, u1_u14_u6_n129, 
       u1_u14_u6_n130, u1_u14_u6_n131, u1_u14_u6_n132, u1_u14_u6_n133, u1_u14_u6_n134, u1_u14_u6_n135, u1_u14_u6_n136, u1_u14_u6_n137, u1_u14_u6_n138, 
       u1_u14_u6_n139, u1_u14_u6_n140, u1_u14_u6_n141, u1_u14_u6_n142, u1_u14_u6_n143, u1_u14_u6_n144, u1_u14_u6_n145, u1_u14_u6_n146, u1_u14_u6_n147, 
       u1_u14_u6_n148, u1_u14_u6_n149, u1_u14_u6_n150, u1_u14_u6_n151, u1_u14_u6_n152, u1_u14_u6_n153, u1_u14_u6_n154, u1_u14_u6_n155, u1_u14_u6_n156, 
       u1_u14_u6_n157, u1_u14_u6_n158, u1_u14_u6_n159, u1_u14_u6_n160, u1_u14_u6_n161, u1_u14_u6_n162, u1_u14_u6_n163, u1_u14_u6_n164, u1_u14_u6_n165, 
       u1_u14_u6_n166, u1_u14_u6_n167, u1_u14_u6_n168, u1_u14_u6_n169, u1_u14_u6_n170, u1_u14_u6_n171, u1_u14_u6_n172, u1_u14_u6_n173, u1_u14_u6_n174, 
       u1_u14_u6_n88, u1_u14_u6_n89, u1_u14_u6_n90, u1_u14_u6_n91, u1_u14_u6_n92, u1_u14_u6_n93, u1_u14_u6_n94, u1_u14_u6_n95, u1_u14_u6_n96, 
       u1_u14_u6_n97, u1_u14_u6_n98, u1_u14_u6_n99, u1_u14_u7_n100, u1_u14_u7_n101, u1_u14_u7_n102, u1_u14_u7_n103, u1_u14_u7_n104, u1_u14_u7_n105, 
       u1_u14_u7_n106, u1_u14_u7_n107, u1_u14_u7_n108, u1_u14_u7_n109, u1_u14_u7_n110, u1_u14_u7_n111, u1_u14_u7_n112, u1_u14_u7_n113, u1_u14_u7_n114, 
       u1_u14_u7_n115, u1_u14_u7_n116, u1_u14_u7_n117, u1_u14_u7_n118, u1_u14_u7_n119, u1_u14_u7_n120, u1_u14_u7_n121, u1_u14_u7_n122, u1_u14_u7_n123, 
       u1_u14_u7_n124, u1_u14_u7_n125, u1_u14_u7_n126, u1_u14_u7_n127, u1_u14_u7_n128, u1_u14_u7_n129, u1_u14_u7_n130, u1_u14_u7_n131, u1_u14_u7_n132, 
       u1_u14_u7_n133, u1_u14_u7_n134, u1_u14_u7_n135, u1_u14_u7_n136, u1_u14_u7_n137, u1_u14_u7_n138, u1_u14_u7_n139, u1_u14_u7_n140, u1_u14_u7_n141, 
       u1_u14_u7_n142, u1_u14_u7_n143, u1_u14_u7_n144, u1_u14_u7_n145, u1_u14_u7_n146, u1_u14_u7_n147, u1_u14_u7_n148, u1_u14_u7_n149, u1_u14_u7_n150, 
       u1_u14_u7_n151, u1_u14_u7_n152, u1_u14_u7_n153, u1_u14_u7_n154, u1_u14_u7_n155, u1_u14_u7_n156, u1_u14_u7_n157, u1_u14_u7_n158, u1_u14_u7_n159, 
       u1_u14_u7_n160, u1_u14_u7_n161, u1_u14_u7_n162, u1_u14_u7_n163, u1_u14_u7_n164, u1_u14_u7_n165, u1_u14_u7_n166, u1_u14_u7_n167, u1_u14_u7_n168, 
       u1_u14_u7_n169, u1_u14_u7_n170, u1_u14_u7_n171, u1_u14_u7_n172, u1_u14_u7_n173, u1_u14_u7_n174, u1_u14_u7_n175, u1_u14_u7_n176, u1_u14_u7_n177, 
       u1_u14_u7_n178, u1_u14_u7_n179, u1_u14_u7_n180, u1_u14_u7_n91, u1_u14_u7_n92, u1_u14_u7_n93, u1_u14_u7_n94, u1_u14_u7_n95, u1_u14_u7_n96, 
       u1_u14_u7_n97, u1_u14_u7_n98, u1_u14_u7_n99, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_19, u1_u15_X_20, 
       u1_u15_X_29, u1_u15_X_30, u1_u15_X_31, u1_u15_X_32, u1_u15_X_34, u1_u15_X_35, u1_u15_u2_n100, u1_u15_u2_n101, u1_u15_u2_n102, 
       u1_u15_u2_n103, u1_u15_u2_n104, u1_u15_u2_n105, u1_u15_u2_n106, u1_u15_u2_n107, u1_u15_u2_n108, u1_u15_u2_n109, u1_u15_u2_n110, u1_u15_u2_n111, 
       u1_u15_u2_n112, u1_u15_u2_n113, u1_u15_u2_n114, u1_u15_u2_n115, u1_u15_u2_n116, u1_u15_u2_n117, u1_u15_u2_n118, u1_u15_u2_n119, u1_u15_u2_n120, 
       u1_u15_u2_n121, u1_u15_u2_n122, u1_u15_u2_n123, u1_u15_u2_n124, u1_u15_u2_n125, u1_u15_u2_n126, u1_u15_u2_n127, u1_u15_u2_n128, u1_u15_u2_n129, 
       u1_u15_u2_n130, u1_u15_u2_n131, u1_u15_u2_n132, u1_u15_u2_n133, u1_u15_u2_n134, u1_u15_u2_n135, u1_u15_u2_n136, u1_u15_u2_n137, u1_u15_u2_n138, 
       u1_u15_u2_n139, u1_u15_u2_n140, u1_u15_u2_n141, u1_u15_u2_n142, u1_u15_u2_n143, u1_u15_u2_n144, u1_u15_u2_n145, u1_u15_u2_n146, u1_u15_u2_n147, 
       u1_u15_u2_n148, u1_u15_u2_n149, u1_u15_u2_n150, u1_u15_u2_n151, u1_u15_u2_n152, u1_u15_u2_n153, u1_u15_u2_n154, u1_u15_u2_n155, u1_u15_u2_n156, 
       u1_u15_u2_n157, u1_u15_u2_n158, u1_u15_u2_n159, u1_u15_u2_n160, u1_u15_u2_n161, u1_u15_u2_n162, u1_u15_u2_n163, u1_u15_u2_n164, u1_u15_u2_n165, 
       u1_u15_u2_n166, u1_u15_u2_n167, u1_u15_u2_n168, u1_u15_u2_n169, u1_u15_u2_n170, u1_u15_u2_n171, u1_u15_u2_n172, u1_u15_u2_n173, u1_u15_u2_n174, 
       u1_u15_u2_n175, u1_u15_u2_n176, u1_u15_u2_n177, u1_u15_u2_n178, u1_u15_u2_n179, u1_u15_u2_n180, u1_u15_u2_n181, u1_u15_u2_n182, u1_u15_u2_n183, 
       u1_u15_u2_n184, u1_u15_u2_n185, u1_u15_u2_n186, u1_u15_u2_n187, u1_u15_u2_n188, u1_u15_u2_n95, u1_u15_u2_n96, u1_u15_u2_n97, u1_u15_u2_n98, 
       u1_u15_u2_n99, u1_u15_u3_n100, u1_u15_u3_n101, u1_u15_u3_n102, u1_u15_u3_n103, u1_u15_u3_n104, u1_u15_u3_n105, u1_u15_u3_n106, u1_u15_u3_n107, 
       u1_u15_u3_n108, u1_u15_u3_n109, u1_u15_u3_n110, u1_u15_u3_n111, u1_u15_u3_n112, u1_u15_u3_n113, u1_u15_u3_n114, u1_u15_u3_n115, u1_u15_u3_n116, 
       u1_u15_u3_n117, u1_u15_u3_n118, u1_u15_u3_n119, u1_u15_u3_n120, u1_u15_u3_n121, u1_u15_u3_n122, u1_u15_u3_n123, u1_u15_u3_n124, u1_u15_u3_n125, 
       u1_u15_u3_n126, u1_u15_u3_n127, u1_u15_u3_n128, u1_u15_u3_n129, u1_u15_u3_n130, u1_u15_u3_n131, u1_u15_u3_n132, u1_u15_u3_n133, u1_u15_u3_n134, 
       u1_u15_u3_n135, u1_u15_u3_n136, u1_u15_u3_n137, u1_u15_u3_n138, u1_u15_u3_n139, u1_u15_u3_n140, u1_u15_u3_n141, u1_u15_u3_n142, u1_u15_u3_n143, 
       u1_u15_u3_n144, u1_u15_u3_n145, u1_u15_u3_n146, u1_u15_u3_n147, u1_u15_u3_n148, u1_u15_u3_n149, u1_u15_u3_n150, u1_u15_u3_n151, u1_u15_u3_n152, 
       u1_u15_u3_n153, u1_u15_u3_n154, u1_u15_u3_n155, u1_u15_u3_n156, u1_u15_u3_n157, u1_u15_u3_n158, u1_u15_u3_n159, u1_u15_u3_n160, u1_u15_u3_n161, 
       u1_u15_u3_n162, u1_u15_u3_n163, u1_u15_u3_n164, u1_u15_u3_n165, u1_u15_u3_n166, u1_u15_u3_n167, u1_u15_u3_n168, u1_u15_u3_n169, u1_u15_u3_n170, 
       u1_u15_u3_n171, u1_u15_u3_n172, u1_u15_u3_n173, u1_u15_u3_n174, u1_u15_u3_n175, u1_u15_u3_n176, u1_u15_u3_n177, u1_u15_u3_n178, u1_u15_u3_n179, 
       u1_u15_u3_n180, u1_u15_u3_n181, u1_u15_u3_n182, u1_u15_u3_n183, u1_u15_u3_n184, u1_u15_u3_n185, u1_u15_u3_n186, u1_u15_u3_n94, u1_u15_u3_n95, 
       u1_u15_u3_n96, u1_u15_u3_n97, u1_u15_u3_n98, u1_u15_u3_n99, u1_u15_u4_n100, u1_u15_u4_n101, u1_u15_u4_n102, u1_u15_u4_n103, u1_u15_u4_n104, 
       u1_u15_u4_n105, u1_u15_u4_n106, u1_u15_u4_n107, u1_u15_u4_n108, u1_u15_u4_n109, u1_u15_u4_n110, u1_u15_u4_n111, u1_u15_u4_n112, u1_u15_u4_n113, 
       u1_u15_u4_n114, u1_u15_u4_n115, u1_u15_u4_n116, u1_u15_u4_n117, u1_u15_u4_n118, u1_u15_u4_n119, u1_u15_u4_n120, u1_u15_u4_n121, u1_u15_u4_n122, 
       u1_u15_u4_n123, u1_u15_u4_n124, u1_u15_u4_n125, u1_u15_u4_n126, u1_u15_u4_n127, u1_u15_u4_n128, u1_u15_u4_n129, u1_u15_u4_n130, u1_u15_u4_n131, 
       u1_u15_u4_n132, u1_u15_u4_n133, u1_u15_u4_n134, u1_u15_u4_n135, u1_u15_u4_n136, u1_u15_u4_n137, u1_u15_u4_n138, u1_u15_u4_n139, u1_u15_u4_n140, 
       u1_u15_u4_n141, u1_u15_u4_n142, u1_u15_u4_n143, u1_u15_u4_n144, u1_u15_u4_n145, u1_u15_u4_n146, u1_u15_u4_n147, u1_u15_u4_n148, u1_u15_u4_n149, 
       u1_u15_u4_n150, u1_u15_u4_n151, u1_u15_u4_n152, u1_u15_u4_n153, u1_u15_u4_n154, u1_u15_u4_n155, u1_u15_u4_n156, u1_u15_u4_n157, u1_u15_u4_n158, 
       u1_u15_u4_n159, u1_u15_u4_n160, u1_u15_u4_n161, u1_u15_u4_n162, u1_u15_u4_n163, u1_u15_u4_n164, u1_u15_u4_n165, u1_u15_u4_n166, u1_u15_u4_n167, 
       u1_u15_u4_n168, u1_u15_u4_n169, u1_u15_u4_n170, u1_u15_u4_n171, u1_u15_u4_n172, u1_u15_u4_n173, u1_u15_u4_n174, u1_u15_u4_n175, u1_u15_u4_n176, 
       u1_u15_u4_n177, u1_u15_u4_n178, u1_u15_u4_n179, u1_u15_u4_n180, u1_u15_u4_n181, u1_u15_u4_n182, u1_u15_u4_n183, u1_u15_u4_n184, u1_u15_u4_n185, 
       u1_u15_u4_n186, u1_u15_u4_n94, u1_u15_u4_n95, u1_u15_u4_n96, u1_u15_u4_n97, u1_u15_u4_n98, u1_u15_u4_n99, u1_u15_u5_n100, u1_u15_u5_n101, 
       u1_u15_u5_n102, u1_u15_u5_n103, u1_u15_u5_n104, u1_u15_u5_n105, u1_u15_u5_n106, u1_u15_u5_n107, u1_u15_u5_n108, u1_u15_u5_n109, u1_u15_u5_n110, 
       u1_u15_u5_n111, u1_u15_u5_n112, u1_u15_u5_n113, u1_u15_u5_n114, u1_u15_u5_n115, u1_u15_u5_n116, u1_u15_u5_n117, u1_u15_u5_n118, u1_u15_u5_n119, 
       u1_u15_u5_n120, u1_u15_u5_n121, u1_u15_u5_n122, u1_u15_u5_n123, u1_u15_u5_n124, u1_u15_u5_n125, u1_u15_u5_n126, u1_u15_u5_n127, u1_u15_u5_n128, 
       u1_u15_u5_n129, u1_u15_u5_n130, u1_u15_u5_n131, u1_u15_u5_n132, u1_u15_u5_n133, u1_u15_u5_n134, u1_u15_u5_n135, u1_u15_u5_n136, u1_u15_u5_n137, 
       u1_u15_u5_n138, u1_u15_u5_n139, u1_u15_u5_n140, u1_u15_u5_n141, u1_u15_u5_n142, u1_u15_u5_n143, u1_u15_u5_n144, u1_u15_u5_n145, u1_u15_u5_n146, 
       u1_u15_u5_n147, u1_u15_u5_n148, u1_u15_u5_n149, u1_u15_u5_n150, u1_u15_u5_n151, u1_u15_u5_n152, u1_u15_u5_n153, u1_u15_u5_n154, u1_u15_u5_n155, 
       u1_u15_u5_n156, u1_u15_u5_n157, u1_u15_u5_n158, u1_u15_u5_n159, u1_u15_u5_n160, u1_u15_u5_n161, u1_u15_u5_n162, u1_u15_u5_n163, u1_u15_u5_n164, 
       u1_u15_u5_n165, u1_u15_u5_n166, u1_u15_u5_n167, u1_u15_u5_n168, u1_u15_u5_n169, u1_u15_u5_n170, u1_u15_u5_n171, u1_u15_u5_n172, u1_u15_u5_n173, 
       u1_u15_u5_n174, u1_u15_u5_n175, u1_u15_u5_n176, u1_u15_u5_n177, u1_u15_u5_n178, u1_u15_u5_n179, u1_u15_u5_n180, u1_u15_u5_n181, u1_u15_u5_n182, 
       u1_u15_u5_n183, u1_u15_u5_n184, u1_u15_u5_n185, u1_u15_u5_n186, u1_u15_u5_n187, u1_u15_u5_n188, u1_u15_u5_n189, u1_u15_u5_n190, u1_u15_u5_n191, 
       u1_u15_u5_n192, u1_u15_u5_n193, u1_u15_u5_n194, u1_u15_u5_n195, u1_u15_u5_n196, u1_u15_u5_n99, u1_u1_X_19, u1_u1_X_20, u1_u1_X_23, 
       u1_u1_X_24, u1_u1_X_25, u1_u1_X_26, u1_u1_X_29, u1_u1_X_30, u1_u1_X_41, u1_u1_X_42, u1_u1_X_43, u1_u1_X_44, 
       u1_u1_X_47, u1_u1_X_48, u1_u1_u3_n100, u1_u1_u3_n101, u1_u1_u3_n102, u1_u1_u3_n103, u1_u1_u3_n104, u1_u1_u3_n105, u1_u1_u3_n106, 
       u1_u1_u3_n107, u1_u1_u3_n108, u1_u1_u3_n109, u1_u1_u3_n110, u1_u1_u3_n111, u1_u1_u3_n112, u1_u1_u3_n113, u1_u1_u3_n114, u1_u1_u3_n115, 
       u1_u1_u3_n116, u1_u1_u3_n117, u1_u1_u3_n118, u1_u1_u3_n119, u1_u1_u3_n120, u1_u1_u3_n121, u1_u1_u3_n122, u1_u1_u3_n123, u1_u1_u3_n124, 
       u1_u1_u3_n125, u1_u1_u3_n126, u1_u1_u3_n127, u1_u1_u3_n128, u1_u1_u3_n129, u1_u1_u3_n130, u1_u1_u3_n131, u1_u1_u3_n132, u1_u1_u3_n133, 
       u1_u1_u3_n134, u1_u1_u3_n135, u1_u1_u3_n136, u1_u1_u3_n137, u1_u1_u3_n138, u1_u1_u3_n139, u1_u1_u3_n140, u1_u1_u3_n141, u1_u1_u3_n142, 
       u1_u1_u3_n143, u1_u1_u3_n144, u1_u1_u3_n145, u1_u1_u3_n146, u1_u1_u3_n147, u1_u1_u3_n148, u1_u1_u3_n149, u1_u1_u3_n150, u1_u1_u3_n151, 
       u1_u1_u3_n152, u1_u1_u3_n153, u1_u1_u3_n154, u1_u1_u3_n155, u1_u1_u3_n156, u1_u1_u3_n157, u1_u1_u3_n158, u1_u1_u3_n159, u1_u1_u3_n160, 
       u1_u1_u3_n161, u1_u1_u3_n162, u1_u1_u3_n163, u1_u1_u3_n164, u1_u1_u3_n165, u1_u1_u3_n166, u1_u1_u3_n167, u1_u1_u3_n168, u1_u1_u3_n169, 
       u1_u1_u3_n170, u1_u1_u3_n171, u1_u1_u3_n172, u1_u1_u3_n173, u1_u1_u3_n174, u1_u1_u3_n175, u1_u1_u3_n176, u1_u1_u3_n177, u1_u1_u3_n178, 
       u1_u1_u3_n179, u1_u1_u3_n180, u1_u1_u3_n181, u1_u1_u3_n182, u1_u1_u3_n183, u1_u1_u3_n184, u1_u1_u3_n185, u1_u1_u3_n186, u1_u1_u3_n94, 
       u1_u1_u3_n95, u1_u1_u3_n96, u1_u1_u3_n97, u1_u1_u3_n98, u1_u1_u3_n99, u1_u1_u4_n100, u1_u1_u4_n101, u1_u1_u4_n102, u1_u1_u4_n103, 
       u1_u1_u4_n104, u1_u1_u4_n105, u1_u1_u4_n106, u1_u1_u4_n107, u1_u1_u4_n108, u1_u1_u4_n109, u1_u1_u4_n110, u1_u1_u4_n111, u1_u1_u4_n112, 
       u1_u1_u4_n113, u1_u1_u4_n114, u1_u1_u4_n115, u1_u1_u4_n116, u1_u1_u4_n117, u1_u1_u4_n118, u1_u1_u4_n119, u1_u1_u4_n120, u1_u1_u4_n121, 
       u1_u1_u4_n122, u1_u1_u4_n123, u1_u1_u4_n124, u1_u1_u4_n125, u1_u1_u4_n126, u1_u1_u4_n127, u1_u1_u4_n128, u1_u1_u4_n129, u1_u1_u4_n130, 
       u1_u1_u4_n131, u1_u1_u4_n132, u1_u1_u4_n133, u1_u1_u4_n134, u1_u1_u4_n135, u1_u1_u4_n136, u1_u1_u4_n137, u1_u1_u4_n138, u1_u1_u4_n139, 
       u1_u1_u4_n140, u1_u1_u4_n141, u1_u1_u4_n142, u1_u1_u4_n143, u1_u1_u4_n144, u1_u1_u4_n145, u1_u1_u4_n146, u1_u1_u4_n147, u1_u1_u4_n148, 
       u1_u1_u4_n149, u1_u1_u4_n150, u1_u1_u4_n151, u1_u1_u4_n152, u1_u1_u4_n153, u1_u1_u4_n154, u1_u1_u4_n155, u1_u1_u4_n156, u1_u1_u4_n157, 
       u1_u1_u4_n158, u1_u1_u4_n159, u1_u1_u4_n160, u1_u1_u4_n161, u1_u1_u4_n162, u1_u1_u4_n163, u1_u1_u4_n164, u1_u1_u4_n165, u1_u1_u4_n166, 
       u1_u1_u4_n167, u1_u1_u4_n168, u1_u1_u4_n169, u1_u1_u4_n170, u1_u1_u4_n171, u1_u1_u4_n172, u1_u1_u4_n173, u1_u1_u4_n174, u1_u1_u4_n175, 
       u1_u1_u4_n176, u1_u1_u4_n177, u1_u1_u4_n178, u1_u1_u4_n179, u1_u1_u4_n180, u1_u1_u4_n181, u1_u1_u4_n182, u1_u1_u4_n183, u1_u1_u4_n184, 
       u1_u1_u4_n185, u1_u1_u4_n186, u1_u1_u4_n94, u1_u1_u4_n95, u1_u1_u4_n96, u1_u1_u4_n97, u1_u1_u4_n98, u1_u1_u4_n99, u1_u1_u6_n100, 
       u1_u1_u6_n101, u1_u1_u6_n102, u1_u1_u6_n103, u1_u1_u6_n104, u1_u1_u6_n105, u1_u1_u6_n106, u1_u1_u6_n107, u1_u1_u6_n108, u1_u1_u6_n109, 
       u1_u1_u6_n110, u1_u1_u6_n111, u1_u1_u6_n112, u1_u1_u6_n113, u1_u1_u6_n114, u1_u1_u6_n115, u1_u1_u6_n116, u1_u1_u6_n117, u1_u1_u6_n118, 
       u1_u1_u6_n119, u1_u1_u6_n120, u1_u1_u6_n121, u1_u1_u6_n122, u1_u1_u6_n123, u1_u1_u6_n124, u1_u1_u6_n125, u1_u1_u6_n126, u1_u1_u6_n127, 
       u1_u1_u6_n128, u1_u1_u6_n129, u1_u1_u6_n130, u1_u1_u6_n131, u1_u1_u6_n132, u1_u1_u6_n133, u1_u1_u6_n134, u1_u1_u6_n135, u1_u1_u6_n136, 
       u1_u1_u6_n137, u1_u1_u6_n138, u1_u1_u6_n139, u1_u1_u6_n140, u1_u1_u6_n141, u1_u1_u6_n142, u1_u1_u6_n143, u1_u1_u6_n144, u1_u1_u6_n145, 
       u1_u1_u6_n146, u1_u1_u6_n147, u1_u1_u6_n148, u1_u1_u6_n149, u1_u1_u6_n150, u1_u1_u6_n151, u1_u1_u6_n152, u1_u1_u6_n153, u1_u1_u6_n154, 
       u1_u1_u6_n155, u1_u1_u6_n156, u1_u1_u6_n157, u1_u1_u6_n158, u1_u1_u6_n159, u1_u1_u6_n160, u1_u1_u6_n161, u1_u1_u6_n162, u1_u1_u6_n163, 
       u1_u1_u6_n164, u1_u1_u6_n165, u1_u1_u6_n166, u1_u1_u6_n167, u1_u1_u6_n168, u1_u1_u6_n169, u1_u1_u6_n170, u1_u1_u6_n171, u1_u1_u6_n172, 
       u1_u1_u6_n173, u1_u1_u6_n174, u1_u1_u6_n88, u1_u1_u6_n89, u1_u1_u6_n90, u1_u1_u6_n91, u1_u1_u6_n92, u1_u1_u6_n93, u1_u1_u6_n94, 
       u1_u1_u6_n95, u1_u1_u6_n96, u1_u1_u6_n97, u1_u1_u6_n98, u1_u1_u6_n99, u1_u1_u7_n100, u1_u1_u7_n101, u1_u1_u7_n102, u1_u1_u7_n103, 
       u1_u1_u7_n104, u1_u1_u7_n105, u1_u1_u7_n106, u1_u1_u7_n107, u1_u1_u7_n108, u1_u1_u7_n109, u1_u1_u7_n110, u1_u1_u7_n111, u1_u1_u7_n112, 
       u1_u1_u7_n113, u1_u1_u7_n114, u1_u1_u7_n115, u1_u1_u7_n116, u1_u1_u7_n117, u1_u1_u7_n118, u1_u1_u7_n119, u1_u1_u7_n120, u1_u1_u7_n121, 
       u1_u1_u7_n122, u1_u1_u7_n123, u1_u1_u7_n124, u1_u1_u7_n125, u1_u1_u7_n126, u1_u1_u7_n127, u1_u1_u7_n128, u1_u1_u7_n129, u1_u1_u7_n130, 
       u1_u1_u7_n131, u1_u1_u7_n132, u1_u1_u7_n133, u1_u1_u7_n134, u1_u1_u7_n135, u1_u1_u7_n136, u1_u1_u7_n137, u1_u1_u7_n138, u1_u1_u7_n139, 
       u1_u1_u7_n140, u1_u1_u7_n141, u1_u1_u7_n142, u1_u1_u7_n143, u1_u1_u7_n144, u1_u1_u7_n145, u1_u1_u7_n146, u1_u1_u7_n147, u1_u1_u7_n148, 
       u1_u1_u7_n149, u1_u1_u7_n150, u1_u1_u7_n151, u1_u1_u7_n152, u1_u1_u7_n153, u1_u1_u7_n154, u1_u1_u7_n155, u1_u1_u7_n156, u1_u1_u7_n157, 
       u1_u1_u7_n158, u1_u1_u7_n159, u1_u1_u7_n160, u1_u1_u7_n161, u1_u1_u7_n162, u1_u1_u7_n163, u1_u1_u7_n164, u1_u1_u7_n165, u1_u1_u7_n166, 
       u1_u1_u7_n167, u1_u1_u7_n168, u1_u1_u7_n169, u1_u1_u7_n170, u1_u1_u7_n171, u1_u1_u7_n172, u1_u1_u7_n173, u1_u1_u7_n174, u1_u1_u7_n175, 
       u1_u1_u7_n176, u1_u1_u7_n177, u1_u1_u7_n178, u1_u1_u7_n179, u1_u1_u7_n180, u1_u1_u7_n91, u1_u1_u7_n92, u1_u1_u7_n93, u1_u1_u7_n94, 
       u1_u1_u7_n95, u1_u1_u7_n96, u1_u1_u7_n97, u1_u1_u7_n98, u1_u1_u7_n99, u1_u2_X_1, u1_u2_X_2, u1_u2_X_37, u1_u2_X_38, 
       u1_u2_X_41, u1_u2_X_42, u1_u2_X_43, u1_u2_X_44, u1_u2_X_47, u1_u2_X_48, u1_u2_X_5, u1_u2_X_6, u1_u2_u0_n100, 
       u1_u2_u0_n101, u1_u2_u0_n102, u1_u2_u0_n103, u1_u2_u0_n104, u1_u2_u0_n105, u1_u2_u0_n106, u1_u2_u0_n107, u1_u2_u0_n108, u1_u2_u0_n109, 
       u1_u2_u0_n110, u1_u2_u0_n111, u1_u2_u0_n112, u1_u2_u0_n113, u1_u2_u0_n114, u1_u2_u0_n115, u1_u2_u0_n116, u1_u2_u0_n117, u1_u2_u0_n118, 
       u1_u2_u0_n119, u1_u2_u0_n120, u1_u2_u0_n121, u1_u2_u0_n122, u1_u2_u0_n123, u1_u2_u0_n124, u1_u2_u0_n125, u1_u2_u0_n126, u1_u2_u0_n127, 
       u1_u2_u0_n128, u1_u2_u0_n129, u1_u2_u0_n130, u1_u2_u0_n131, u1_u2_u0_n132, u1_u2_u0_n133, u1_u2_u0_n134, u1_u2_u0_n135, u1_u2_u0_n136, 
       u1_u2_u0_n137, u1_u2_u0_n138, u1_u2_u0_n139, u1_u2_u0_n140, u1_u2_u0_n141, u1_u2_u0_n142, u1_u2_u0_n143, u1_u2_u0_n144, u1_u2_u0_n145, 
       u1_u2_u0_n146, u1_u2_u0_n147, u1_u2_u0_n148, u1_u2_u0_n149, u1_u2_u0_n150, u1_u2_u0_n151, u1_u2_u0_n152, u1_u2_u0_n153, u1_u2_u0_n154, 
       u1_u2_u0_n155, u1_u2_u0_n156, u1_u2_u0_n157, u1_u2_u0_n158, u1_u2_u0_n159, u1_u2_u0_n160, u1_u2_u0_n161, u1_u2_u0_n162, u1_u2_u0_n163, 
       u1_u2_u0_n164, u1_u2_u0_n165, u1_u2_u0_n166, u1_u2_u0_n167, u1_u2_u0_n168, u1_u2_u0_n169, u1_u2_u0_n170, u1_u2_u0_n171, u1_u2_u0_n172, 
       u1_u2_u0_n173, u1_u2_u0_n174, u1_u2_u0_n88, u1_u2_u0_n89, u1_u2_u0_n90, u1_u2_u0_n91, u1_u2_u0_n92, u1_u2_u0_n93, u1_u2_u0_n94, 
       u1_u2_u0_n95, u1_u2_u0_n96, u1_u2_u0_n97, u1_u2_u0_n98, u1_u2_u0_n99, u1_u2_u6_n100, u1_u2_u6_n101, u1_u2_u6_n102, u1_u2_u6_n103, 
       u1_u2_u6_n104, u1_u2_u6_n105, u1_u2_u6_n106, u1_u2_u6_n107, u1_u2_u6_n108, u1_u2_u6_n109, u1_u2_u6_n110, u1_u2_u6_n111, u1_u2_u6_n112, 
       u1_u2_u6_n113, u1_u2_u6_n114, u1_u2_u6_n115, u1_u2_u6_n116, u1_u2_u6_n117, u1_u2_u6_n118, u1_u2_u6_n119, u1_u2_u6_n120, u1_u2_u6_n121, 
       u1_u2_u6_n122, u1_u2_u6_n123, u1_u2_u6_n124, u1_u2_u6_n125, u1_u2_u6_n126, u1_u2_u6_n127, u1_u2_u6_n128, u1_u2_u6_n129, u1_u2_u6_n130, 
       u1_u2_u6_n131, u1_u2_u6_n132, u1_u2_u6_n133, u1_u2_u6_n134, u1_u2_u6_n135, u1_u2_u6_n136, u1_u2_u6_n137, u1_u2_u6_n138, u1_u2_u6_n139, 
       u1_u2_u6_n140, u1_u2_u6_n141, u1_u2_u6_n142, u1_u2_u6_n143, u1_u2_u6_n144, u1_u2_u6_n145, u1_u2_u6_n146, u1_u2_u6_n147, u1_u2_u6_n148, 
       u1_u2_u6_n149, u1_u2_u6_n150, u1_u2_u6_n151, u1_u2_u6_n152, u1_u2_u6_n153, u1_u2_u6_n154, u1_u2_u6_n155, u1_u2_u6_n156, u1_u2_u6_n157, 
       u1_u2_u6_n158, u1_u2_u6_n159, u1_u2_u6_n160, u1_u2_u6_n161, u1_u2_u6_n162, u1_u2_u6_n163, u1_u2_u6_n164, u1_u2_u6_n165, u1_u2_u6_n166, 
       u1_u2_u6_n167, u1_u2_u6_n168, u1_u2_u6_n169, u1_u2_u6_n170, u1_u2_u6_n171, u1_u2_u6_n172, u1_u2_u6_n173, u1_u2_u6_n174, u1_u2_u6_n88, 
       u1_u2_u6_n89, u1_u2_u6_n90, u1_u2_u6_n91, u1_u2_u6_n92, u1_u2_u6_n93, u1_u2_u6_n94, u1_u2_u6_n95, u1_u2_u6_n96, u1_u2_u6_n97, 
       u1_u2_u6_n98, u1_u2_u6_n99, u1_u2_u7_n100, u1_u2_u7_n101, u1_u2_u7_n102, u1_u2_u7_n103, u1_u2_u7_n104, u1_u2_u7_n105, u1_u2_u7_n106, 
       u1_u2_u7_n107, u1_u2_u7_n108, u1_u2_u7_n109, u1_u2_u7_n110, u1_u2_u7_n111, u1_u2_u7_n112, u1_u2_u7_n113, u1_u2_u7_n114, u1_u2_u7_n115, 
       u1_u2_u7_n116, u1_u2_u7_n117, u1_u2_u7_n118, u1_u2_u7_n119, u1_u2_u7_n120, u1_u2_u7_n121, u1_u2_u7_n122, u1_u2_u7_n123, u1_u2_u7_n124, 
       u1_u2_u7_n125, u1_u2_u7_n126, u1_u2_u7_n127, u1_u2_u7_n128, u1_u2_u7_n129, u1_u2_u7_n130, u1_u2_u7_n131, u1_u2_u7_n132, u1_u2_u7_n133, 
       u1_u2_u7_n134, u1_u2_u7_n135, u1_u2_u7_n136, u1_u2_u7_n137, u1_u2_u7_n138, u1_u2_u7_n139, u1_u2_u7_n140, u1_u2_u7_n141, u1_u2_u7_n142, 
       u1_u2_u7_n143, u1_u2_u7_n144, u1_u2_u7_n145, u1_u2_u7_n146, u1_u2_u7_n147, u1_u2_u7_n148, u1_u2_u7_n149, u1_u2_u7_n150, u1_u2_u7_n151, 
       u1_u2_u7_n152, u1_u2_u7_n153, u1_u2_u7_n154, u1_u2_u7_n155, u1_u2_u7_n156, u1_u2_u7_n157, u1_u2_u7_n158, u1_u2_u7_n159, u1_u2_u7_n160, 
       u1_u2_u7_n161, u1_u2_u7_n162, u1_u2_u7_n163, u1_u2_u7_n164, u1_u2_u7_n165, u1_u2_u7_n166, u1_u2_u7_n167, u1_u2_u7_n168, u1_u2_u7_n169, 
       u1_u2_u7_n170, u1_u2_u7_n171, u1_u2_u7_n172, u1_u2_u7_n173, u1_u2_u7_n174, u1_u2_u7_n175, u1_u2_u7_n176, u1_u2_u7_n177, u1_u2_u7_n178, 
       u1_u2_u7_n179, u1_u2_u7_n180, u1_u2_u7_n91, u1_u2_u7_n92, u1_u2_u7_n93, u1_u2_u7_n94, u1_u2_u7_n95, u1_u2_u7_n96, u1_u2_u7_n97, 
       u1_u2_u7_n98, u1_u2_u7_n99, u1_u3_X_1, u1_u3_X_10, u1_u3_X_11, u1_u3_X_12, u1_u3_X_2, u1_u3_X_3, u1_u3_X_6, 
       u1_u3_X_8, u1_u3_u0_n100, u1_u3_u0_n101, u1_u3_u0_n102, u1_u3_u0_n103, u1_u3_u0_n104, u1_u3_u0_n105, u1_u3_u0_n106, u1_u3_u0_n107, 
       u1_u3_u0_n108, u1_u3_u0_n109, u1_u3_u0_n110, u1_u3_u0_n111, u1_u3_u0_n112, u1_u3_u0_n113, u1_u3_u0_n114, u1_u3_u0_n115, u1_u3_u0_n116, 
       u1_u3_u0_n117, u1_u3_u0_n118, u1_u3_u0_n119, u1_u3_u0_n120, u1_u3_u0_n121, u1_u3_u0_n122, u1_u3_u0_n123, u1_u3_u0_n124, u1_u3_u0_n125, 
       u1_u3_u0_n126, u1_u3_u0_n127, u1_u3_u0_n128, u1_u3_u0_n129, u1_u3_u0_n130, u1_u3_u0_n131, u1_u3_u0_n132, u1_u3_u0_n133, u1_u3_u0_n134, 
       u1_u3_u0_n135, u1_u3_u0_n136, u1_u3_u0_n137, u1_u3_u0_n138, u1_u3_u0_n139, u1_u3_u0_n140, u1_u3_u0_n141, u1_u3_u0_n142, u1_u3_u0_n143, 
       u1_u3_u0_n144, u1_u3_u0_n145, u1_u3_u0_n146, u1_u3_u0_n147, u1_u3_u0_n148, u1_u3_u0_n149, u1_u3_u0_n150, u1_u3_u0_n151, u1_u3_u0_n152, 
       u1_u3_u0_n153, u1_u3_u0_n154, u1_u3_u0_n155, u1_u3_u0_n156, u1_u3_u0_n157, u1_u3_u0_n158, u1_u3_u0_n159, u1_u3_u0_n160, u1_u3_u0_n161, 
       u1_u3_u0_n162, u1_u3_u0_n163, u1_u3_u0_n164, u1_u3_u0_n165, u1_u3_u0_n166, u1_u3_u0_n167, u1_u3_u0_n168, u1_u3_u0_n169, u1_u3_u0_n170, 
       u1_u3_u0_n171, u1_u3_u0_n172, u1_u3_u0_n173, u1_u3_u0_n174, u1_u3_u0_n88, u1_u3_u0_n89, u1_u3_u0_n90, u1_u3_u0_n91, u1_u3_u0_n92, 
       u1_u3_u0_n93, u1_u3_u0_n94, u1_u3_u0_n95, u1_u3_u0_n96, u1_u3_u0_n97, u1_u3_u0_n98, u1_u3_u0_n99, u1_u3_u1_n100, u1_u3_u1_n101, 
       u1_u3_u1_n102, u1_u3_u1_n103, u1_u3_u1_n104, u1_u3_u1_n105, u1_u3_u1_n106, u1_u3_u1_n107, u1_u3_u1_n108, u1_u3_u1_n109, u1_u3_u1_n110, 
       u1_u3_u1_n111, u1_u3_u1_n112, u1_u3_u1_n113, u1_u3_u1_n114, u1_u3_u1_n115, u1_u3_u1_n116, u1_u3_u1_n117, u1_u3_u1_n118, u1_u3_u1_n119, 
       u1_u3_u1_n120, u1_u3_u1_n121, u1_u3_u1_n122, u1_u3_u1_n123, u1_u3_u1_n124, u1_u3_u1_n125, u1_u3_u1_n126, u1_u3_u1_n127, u1_u3_u1_n128, 
       u1_u3_u1_n129, u1_u3_u1_n130, u1_u3_u1_n131, u1_u3_u1_n132, u1_u3_u1_n133, u1_u3_u1_n134, u1_u3_u1_n135, u1_u3_u1_n136, u1_u3_u1_n137, 
       u1_u3_u1_n138, u1_u3_u1_n139, u1_u3_u1_n140, u1_u3_u1_n141, u1_u3_u1_n142, u1_u3_u1_n143, u1_u3_u1_n144, u1_u3_u1_n145, u1_u3_u1_n146, 
       u1_u3_u1_n147, u1_u3_u1_n148, u1_u3_u1_n149, u1_u3_u1_n150, u1_u3_u1_n151, u1_u3_u1_n152, u1_u3_u1_n153, u1_u3_u1_n154, u1_u3_u1_n155, 
       u1_u3_u1_n156, u1_u3_u1_n157, u1_u3_u1_n158, u1_u3_u1_n159, u1_u3_u1_n160, u1_u3_u1_n161, u1_u3_u1_n162, u1_u3_u1_n163, u1_u3_u1_n164, 
       u1_u3_u1_n165, u1_u3_u1_n166, u1_u3_u1_n167, u1_u3_u1_n168, u1_u3_u1_n169, u1_u3_u1_n170, u1_u3_u1_n171, u1_u3_u1_n172, u1_u3_u1_n173, 
       u1_u3_u1_n174, u1_u3_u1_n175, u1_u3_u1_n176, u1_u3_u1_n177, u1_u3_u1_n178, u1_u3_u1_n179, u1_u3_u1_n180, u1_u3_u1_n181, u1_u3_u1_n182, 
       u1_u3_u1_n183, u1_u3_u1_n184, u1_u3_u1_n185, u1_u3_u1_n186, u1_u3_u1_n187, u1_u3_u1_n188, u1_u3_u1_n95, u1_u3_u1_n96, u1_u3_u1_n97, 
       u1_u3_u1_n98, u1_u3_u1_n99, u1_u4_X_19, u1_u4_X_20, u1_u4_X_22, u1_u4_X_23, u1_u4_X_24, u1_u4_u3_n100, u1_u4_u3_n101, 
       u1_u4_u3_n102, u1_u4_u3_n103, u1_u4_u3_n104, u1_u4_u3_n105, u1_u4_u3_n106, u1_u4_u3_n107, u1_u4_u3_n108, u1_u4_u3_n109, u1_u4_u3_n110, 
       u1_u4_u3_n111, u1_u4_u3_n112, u1_u4_u3_n113, u1_u4_u3_n114, u1_u4_u3_n115, u1_u4_u3_n116, u1_u4_u3_n117, u1_u4_u3_n118, u1_u4_u3_n119, 
       u1_u4_u3_n120, u1_u4_u3_n121, u1_u4_u3_n122, u1_u4_u3_n123, u1_u4_u3_n124, u1_u4_u3_n125, u1_u4_u3_n126, u1_u4_u3_n127, u1_u4_u3_n128, 
       u1_u4_u3_n129, u1_u4_u3_n130, u1_u4_u3_n131, u1_u4_u3_n132, u1_u4_u3_n133, u1_u4_u3_n134, u1_u4_u3_n135, u1_u4_u3_n136, u1_u4_u3_n137, 
       u1_u4_u3_n138, u1_u4_u3_n139, u1_u4_u3_n140, u1_u4_u3_n141, u1_u4_u3_n142, u1_u4_u3_n143, u1_u4_u3_n144, u1_u4_u3_n145, u1_u4_u3_n146, 
       u1_u4_u3_n147, u1_u4_u3_n148, u1_u4_u3_n149, u1_u4_u3_n150, u1_u4_u3_n151, u1_u4_u3_n152, u1_u4_u3_n153, u1_u4_u3_n154, u1_u4_u3_n155, 
       u1_u4_u3_n156, u1_u4_u3_n157, u1_u4_u3_n158, u1_u4_u3_n159, u1_u4_u3_n160, u1_u4_u3_n161, u1_u4_u3_n162, u1_u4_u3_n163, u1_u4_u3_n164, 
       u1_u4_u3_n165, u1_u4_u3_n166, u1_u4_u3_n167, u1_u4_u3_n168, u1_u4_u3_n169, u1_u4_u3_n170, u1_u4_u3_n171, u1_u4_u3_n172, u1_u4_u3_n173, 
       u1_u4_u3_n174, u1_u4_u3_n175, u1_u4_u3_n176, u1_u4_u3_n177, u1_u4_u3_n178, u1_u4_u3_n179, u1_u4_u3_n180, u1_u4_u3_n181, u1_u4_u3_n182, 
       u1_u4_u3_n183, u1_u4_u3_n184, u1_u4_u3_n185, u1_u4_u3_n186, u1_u4_u3_n94, u1_u4_u3_n95, u1_u4_u3_n96, u1_u4_u3_n97, u1_u4_u3_n98, 
       u1_u4_u3_n99, u1_u5_X_25, u1_u5_X_26, u1_u5_X_29, u1_u5_X_30, u1_u5_X_31, u1_u5_X_32, u1_u5_X_35, u1_u5_X_36, 
       u1_u5_u4_n100, u1_u5_u4_n101, u1_u5_u4_n102, u1_u5_u4_n103, u1_u5_u4_n104, u1_u5_u4_n105, u1_u5_u4_n106, u1_u5_u4_n107, u1_u5_u4_n108, 
       u1_u5_u4_n109, u1_u5_u4_n110, u1_u5_u4_n111, u1_u5_u4_n112, u1_u5_u4_n113, u1_u5_u4_n114, u1_u5_u4_n115, u1_u5_u4_n116, u1_u5_u4_n117, 
       u1_u5_u4_n118, u1_u5_u4_n119, u1_u5_u4_n120, u1_u5_u4_n121, u1_u5_u4_n122, u1_u5_u4_n123, u1_u5_u4_n124, u1_u5_u4_n125, u1_u5_u4_n126, 
       u1_u5_u4_n127, u1_u5_u4_n128, u1_u5_u4_n129, u1_u5_u4_n130, u1_u5_u4_n131, u1_u5_u4_n132, u1_u5_u4_n133, u1_u5_u4_n134, u1_u5_u4_n135, 
       u1_u5_u4_n136, u1_u5_u4_n137, u1_u5_u4_n138, u1_u5_u4_n139, u1_u5_u4_n140, u1_u5_u4_n141, u1_u5_u4_n142, u1_u5_u4_n143, u1_u5_u4_n144, 
       u1_u5_u4_n145, u1_u5_u4_n146, u1_u5_u4_n147, u1_u5_u4_n148, u1_u5_u4_n149, u1_u5_u4_n150, u1_u5_u4_n151, u1_u5_u4_n152, u1_u5_u4_n153, 
       u1_u5_u4_n154, u1_u5_u4_n155, u1_u5_u4_n156, u1_u5_u4_n157, u1_u5_u4_n158, u1_u5_u4_n159, u1_u5_u4_n160, u1_u5_u4_n161, u1_u5_u4_n162, 
       u1_u5_u4_n163, u1_u5_u4_n164, u1_u5_u4_n165, u1_u5_u4_n166, u1_u5_u4_n167, u1_u5_u4_n168, u1_u5_u4_n169, u1_u5_u4_n170, u1_u5_u4_n171, 
       u1_u5_u4_n172, u1_u5_u4_n173, u1_u5_u4_n174, u1_u5_u4_n175, u1_u5_u4_n176, u1_u5_u4_n177, u1_u5_u4_n178, u1_u5_u4_n179, u1_u5_u4_n180, 
       u1_u5_u4_n181, u1_u5_u4_n182, u1_u5_u4_n183, u1_u5_u4_n184, u1_u5_u4_n185, u1_u5_u4_n186, u1_u5_u4_n94, u1_u5_u4_n95, u1_u5_u4_n96, 
       u1_u5_u4_n97, u1_u5_u4_n98, u1_u5_u4_n99, u1_u5_u5_n100, u1_u5_u5_n101, u1_u5_u5_n102, u1_u5_u5_n103, u1_u5_u5_n104, u1_u5_u5_n105, 
       u1_u5_u5_n106, u1_u5_u5_n107, u1_u5_u5_n108, u1_u5_u5_n109, u1_u5_u5_n110, u1_u5_u5_n111, u1_u5_u5_n112, u1_u5_u5_n113, u1_u5_u5_n114, 
       u1_u5_u5_n115, u1_u5_u5_n116, u1_u5_u5_n117, u1_u5_u5_n118, u1_u5_u5_n119, u1_u5_u5_n120, u1_u5_u5_n121, u1_u5_u5_n122, u1_u5_u5_n123, 
       u1_u5_u5_n124, u1_u5_u5_n125, u1_u5_u5_n126, u1_u5_u5_n127, u1_u5_u5_n128, u1_u5_u5_n129, u1_u5_u5_n130, u1_u5_u5_n131, u1_u5_u5_n132, 
       u1_u5_u5_n133, u1_u5_u5_n134, u1_u5_u5_n135, u1_u5_u5_n136, u1_u5_u5_n137, u1_u5_u5_n138, u1_u5_u5_n139, u1_u5_u5_n140, u1_u5_u5_n141, 
       u1_u5_u5_n142, u1_u5_u5_n143, u1_u5_u5_n144, u1_u5_u5_n145, u1_u5_u5_n146, u1_u5_u5_n147, u1_u5_u5_n148, u1_u5_u5_n149, u1_u5_u5_n150, 
       u1_u5_u5_n151, u1_u5_u5_n152, u1_u5_u5_n153, u1_u5_u5_n154, u1_u5_u5_n155, u1_u5_u5_n156, u1_u5_u5_n157, u1_u5_u5_n158, u1_u5_u5_n159, 
       u1_u5_u5_n160, u1_u5_u5_n161, u1_u5_u5_n162, u1_u5_u5_n163, u1_u5_u5_n164, u1_u5_u5_n165, u1_u5_u5_n166, u1_u5_u5_n167, u1_u5_u5_n168, 
       u1_u5_u5_n169, u1_u5_u5_n170, u1_u5_u5_n171, u1_u5_u5_n172, u1_u5_u5_n173, u1_u5_u5_n174, u1_u5_u5_n175, u1_u5_u5_n176, u1_u5_u5_n177, 
       u1_u5_u5_n178, u1_u5_u5_n179, u1_u5_u5_n180, u1_u5_u5_n181, u1_u5_u5_n182, u1_u5_u5_n183, u1_u5_u5_n184, u1_u5_u5_n185, u1_u5_u5_n186, 
       u1_u5_u5_n187, u1_u5_u5_n188, u1_u5_u5_n189, u1_u5_u5_n190, u1_u5_u5_n191, u1_u5_u5_n192, u1_u5_u5_n193, u1_u5_u5_n194, u1_u5_u5_n195, 
       u1_u5_u5_n196, u1_u5_u5_n99, u1_u6_X_1, u1_u6_X_11, u1_u6_X_12, u1_u6_X_13, u1_u6_X_14, u1_u6_X_17, u1_u6_X_18, 
       u1_u6_X_2, u1_u6_X_37, u1_u6_X_38, u1_u6_X_41, u1_u6_X_42, u1_u6_X_43, u1_u6_X_44, u1_u6_X_46, u1_u6_X_47, 
       u1_u6_X_48, u1_u6_X_5, u1_u6_X_6, u1_u6_X_7, u1_u6_X_8, u1_u6_u0_n100, u1_u6_u0_n101, u1_u6_u0_n102, u1_u6_u0_n103, 
       u1_u6_u0_n104, u1_u6_u0_n105, u1_u6_u0_n106, u1_u6_u0_n107, u1_u6_u0_n108, u1_u6_u0_n109, u1_u6_u0_n110, u1_u6_u0_n111, u1_u6_u0_n112, 
       u1_u6_u0_n113, u1_u6_u0_n114, u1_u6_u0_n115, u1_u6_u0_n116, u1_u6_u0_n117, u1_u6_u0_n118, u1_u6_u0_n119, u1_u6_u0_n120, u1_u6_u0_n121, 
       u1_u6_u0_n122, u1_u6_u0_n123, u1_u6_u0_n124, u1_u6_u0_n125, u1_u6_u0_n126, u1_u6_u0_n127, u1_u6_u0_n128, u1_u6_u0_n129, u1_u6_u0_n130, 
       u1_u6_u0_n131, u1_u6_u0_n132, u1_u6_u0_n133, u1_u6_u0_n134, u1_u6_u0_n135, u1_u6_u0_n136, u1_u6_u0_n137, u1_u6_u0_n138, u1_u6_u0_n139, 
       u1_u6_u0_n140, u1_u6_u0_n141, u1_u6_u0_n142, u1_u6_u0_n143, u1_u6_u0_n144, u1_u6_u0_n145, u1_u6_u0_n146, u1_u6_u0_n147, u1_u6_u0_n148, 
       u1_u6_u0_n149, u1_u6_u0_n150, u1_u6_u0_n151, u1_u6_u0_n152, u1_u6_u0_n153, u1_u6_u0_n154, u1_u6_u0_n155, u1_u6_u0_n156, u1_u6_u0_n157, 
       u1_u6_u0_n158, u1_u6_u0_n159, u1_u6_u0_n160, u1_u6_u0_n161, u1_u6_u0_n162, u1_u6_u0_n163, u1_u6_u0_n164, u1_u6_u0_n165, u1_u6_u0_n166, 
       u1_u6_u0_n167, u1_u6_u0_n168, u1_u6_u0_n169, u1_u6_u0_n170, u1_u6_u0_n171, u1_u6_u0_n172, u1_u6_u0_n173, u1_u6_u0_n174, u1_u6_u0_n88, 
       u1_u6_u0_n89, u1_u6_u0_n90, u1_u6_u0_n91, u1_u6_u0_n92, u1_u6_u0_n93, u1_u6_u0_n94, u1_u6_u0_n95, u1_u6_u0_n96, u1_u6_u0_n97, 
       u1_u6_u0_n98, u1_u6_u0_n99, u1_u6_u1_n100, u1_u6_u1_n101, u1_u6_u1_n102, u1_u6_u1_n103, u1_u6_u1_n104, u1_u6_u1_n105, u1_u6_u1_n106, 
       u1_u6_u1_n107, u1_u6_u1_n108, u1_u6_u1_n109, u1_u6_u1_n110, u1_u6_u1_n111, u1_u6_u1_n112, u1_u6_u1_n113, u1_u6_u1_n114, u1_u6_u1_n115, 
       u1_u6_u1_n116, u1_u6_u1_n117, u1_u6_u1_n118, u1_u6_u1_n119, u1_u6_u1_n120, u1_u6_u1_n121, u1_u6_u1_n122, u1_u6_u1_n123, u1_u6_u1_n124, 
       u1_u6_u1_n125, u1_u6_u1_n126, u1_u6_u1_n127, u1_u6_u1_n128, u1_u6_u1_n129, u1_u6_u1_n130, u1_u6_u1_n131, u1_u6_u1_n132, u1_u6_u1_n133, 
       u1_u6_u1_n134, u1_u6_u1_n135, u1_u6_u1_n136, u1_u6_u1_n137, u1_u6_u1_n138, u1_u6_u1_n139, u1_u6_u1_n140, u1_u6_u1_n141, u1_u6_u1_n142, 
       u1_u6_u1_n143, u1_u6_u1_n144, u1_u6_u1_n145, u1_u6_u1_n146, u1_u6_u1_n147, u1_u6_u1_n148, u1_u6_u1_n149, u1_u6_u1_n150, u1_u6_u1_n151, 
       u1_u6_u1_n152, u1_u6_u1_n153, u1_u6_u1_n154, u1_u6_u1_n155, u1_u6_u1_n156, u1_u6_u1_n157, u1_u6_u1_n158, u1_u6_u1_n159, u1_u6_u1_n160, 
       u1_u6_u1_n161, u1_u6_u1_n162, u1_u6_u1_n163, u1_u6_u1_n164, u1_u6_u1_n165, u1_u6_u1_n166, u1_u6_u1_n167, u1_u6_u1_n168, u1_u6_u1_n169, 
       u1_u6_u1_n170, u1_u6_u1_n171, u1_u6_u1_n172, u1_u6_u1_n173, u1_u6_u1_n174, u1_u6_u1_n175, u1_u6_u1_n176, u1_u6_u1_n177, u1_u6_u1_n178, 
       u1_u6_u1_n179, u1_u6_u1_n180, u1_u6_u1_n181, u1_u6_u1_n182, u1_u6_u1_n183, u1_u6_u1_n184, u1_u6_u1_n185, u1_u6_u1_n186, u1_u6_u1_n187, 
       u1_u6_u1_n188, u1_u6_u1_n95, u1_u6_u1_n96, u1_u6_u1_n97, u1_u6_u1_n98, u1_u6_u1_n99, u1_u6_u2_n100, u1_u6_u2_n101, u1_u6_u2_n102, 
       u1_u6_u2_n103, u1_u6_u2_n104, u1_u6_u2_n105, u1_u6_u2_n106, u1_u6_u2_n107, u1_u6_u2_n108, u1_u6_u2_n109, u1_u6_u2_n110, u1_u6_u2_n111, 
       u1_u6_u2_n112, u1_u6_u2_n113, u1_u6_u2_n114, u1_u6_u2_n115, u1_u6_u2_n116, u1_u6_u2_n117, u1_u6_u2_n118, u1_u6_u2_n119, u1_u6_u2_n120, 
       u1_u6_u2_n121, u1_u6_u2_n122, u1_u6_u2_n123, u1_u6_u2_n124, u1_u6_u2_n125, u1_u6_u2_n126, u1_u6_u2_n127, u1_u6_u2_n128, u1_u6_u2_n129, 
       u1_u6_u2_n130, u1_u6_u2_n131, u1_u6_u2_n132, u1_u6_u2_n133, u1_u6_u2_n134, u1_u6_u2_n135, u1_u6_u2_n136, u1_u6_u2_n137, u1_u6_u2_n138, 
       u1_u6_u2_n139, u1_u6_u2_n140, u1_u6_u2_n141, u1_u6_u2_n142, u1_u6_u2_n143, u1_u6_u2_n144, u1_u6_u2_n145, u1_u6_u2_n146, u1_u6_u2_n147, 
       u1_u6_u2_n148, u1_u6_u2_n149, u1_u6_u2_n150, u1_u6_u2_n151, u1_u6_u2_n152, u1_u6_u2_n153, u1_u6_u2_n154, u1_u6_u2_n155, u1_u6_u2_n156, 
       u1_u6_u2_n157, u1_u6_u2_n158, u1_u6_u2_n159, u1_u6_u2_n160, u1_u6_u2_n161, u1_u6_u2_n162, u1_u6_u2_n163, u1_u6_u2_n164, u1_u6_u2_n165, 
       u1_u6_u2_n166, u1_u6_u2_n167, u1_u6_u2_n168, u1_u6_u2_n169, u1_u6_u2_n170, u1_u6_u2_n171, u1_u6_u2_n172, u1_u6_u2_n173, u1_u6_u2_n174, 
       u1_u6_u2_n175, u1_u6_u2_n176, u1_u6_u2_n177, u1_u6_u2_n178, u1_u6_u2_n179, u1_u6_u2_n180, u1_u6_u2_n181, u1_u6_u2_n182, u1_u6_u2_n183, 
       u1_u6_u2_n184, u1_u6_u2_n185, u1_u6_u2_n186, u1_u6_u2_n187, u1_u6_u2_n188, u1_u6_u2_n95, u1_u6_u2_n96, u1_u6_u2_n97, u1_u6_u2_n98, 
       u1_u6_u2_n99, u1_u6_u6_n100, u1_u6_u6_n101, u1_u6_u6_n102, u1_u6_u6_n103, u1_u6_u6_n104, u1_u6_u6_n105, u1_u6_u6_n106, u1_u6_u6_n107, 
       u1_u6_u6_n108, u1_u6_u6_n109, u1_u6_u6_n110, u1_u6_u6_n111, u1_u6_u6_n112, u1_u6_u6_n113, u1_u6_u6_n114, u1_u6_u6_n115, u1_u6_u6_n116, 
       u1_u6_u6_n117, u1_u6_u6_n118, u1_u6_u6_n119, u1_u6_u6_n120, u1_u6_u6_n121, u1_u6_u6_n122, u1_u6_u6_n123, u1_u6_u6_n124, u1_u6_u6_n125, 
       u1_u6_u6_n126, u1_u6_u6_n127, u1_u6_u6_n128, u1_u6_u6_n129, u1_u6_u6_n130, u1_u6_u6_n131, u1_u6_u6_n132, u1_u6_u6_n133, u1_u6_u6_n134, 
       u1_u6_u6_n135, u1_u6_u6_n136, u1_u6_u6_n137, u1_u6_u6_n138, u1_u6_u6_n139, u1_u6_u6_n140, u1_u6_u6_n141, u1_u6_u6_n142, u1_u6_u6_n143, 
       u1_u6_u6_n144, u1_u6_u6_n145, u1_u6_u6_n146, u1_u6_u6_n147, u1_u6_u6_n148, u1_u6_u6_n149, u1_u6_u6_n150, u1_u6_u6_n151, u1_u6_u6_n152, 
       u1_u6_u6_n153, u1_u6_u6_n154, u1_u6_u6_n155, u1_u6_u6_n156, u1_u6_u6_n157, u1_u6_u6_n158, u1_u6_u6_n159, u1_u6_u6_n160, u1_u6_u6_n161, 
       u1_u6_u6_n162, u1_u6_u6_n163, u1_u6_u6_n164, u1_u6_u6_n165, u1_u6_u6_n166, u1_u6_u6_n167, u1_u6_u6_n168, u1_u6_u6_n169, u1_u6_u6_n170, 
       u1_u6_u6_n171, u1_u6_u6_n172, u1_u6_u6_n173, u1_u6_u6_n174, u1_u6_u6_n88, u1_u6_u6_n89, u1_u6_u6_n90, u1_u6_u6_n91, u1_u6_u6_n92, 
       u1_u6_u6_n93, u1_u6_u6_n94, u1_u6_u6_n95, u1_u6_u6_n96, u1_u6_u6_n97, u1_u6_u6_n98, u1_u6_u6_n99, u1_u6_u7_n100, u1_u6_u7_n101, 
       u1_u6_u7_n102, u1_u6_u7_n103, u1_u6_u7_n104, u1_u6_u7_n105, u1_u6_u7_n106, u1_u6_u7_n107, u1_u6_u7_n108, u1_u6_u7_n109, u1_u6_u7_n110, 
       u1_u6_u7_n111, u1_u6_u7_n112, u1_u6_u7_n113, u1_u6_u7_n114, u1_u6_u7_n115, u1_u6_u7_n116, u1_u6_u7_n117, u1_u6_u7_n118, u1_u6_u7_n119, 
       u1_u6_u7_n120, u1_u6_u7_n121, u1_u6_u7_n122, u1_u6_u7_n123, u1_u6_u7_n124, u1_u6_u7_n125, u1_u6_u7_n126, u1_u6_u7_n127, u1_u6_u7_n128, 
       u1_u6_u7_n129, u1_u6_u7_n130, u1_u6_u7_n131, u1_u6_u7_n132, u1_u6_u7_n133, u1_u6_u7_n134, u1_u6_u7_n135, u1_u6_u7_n136, u1_u6_u7_n137, 
       u1_u6_u7_n138, u1_u6_u7_n139, u1_u6_u7_n140, u1_u6_u7_n141, u1_u6_u7_n142, u1_u6_u7_n143, u1_u6_u7_n144, u1_u6_u7_n145, u1_u6_u7_n146, 
       u1_u6_u7_n147, u1_u6_u7_n148, u1_u6_u7_n149, u1_u6_u7_n150, u1_u6_u7_n151, u1_u6_u7_n152, u1_u6_u7_n153, u1_u6_u7_n154, u1_u6_u7_n155, 
       u1_u6_u7_n156, u1_u6_u7_n157, u1_u6_u7_n158, u1_u6_u7_n159, u1_u6_u7_n160, u1_u6_u7_n161, u1_u6_u7_n162, u1_u6_u7_n163, u1_u6_u7_n164, 
       u1_u6_u7_n165, u1_u6_u7_n166, u1_u6_u7_n167, u1_u6_u7_n168, u1_u6_u7_n169, u1_u6_u7_n170, u1_u6_u7_n171, u1_u6_u7_n172, u1_u6_u7_n173, 
       u1_u6_u7_n174, u1_u6_u7_n175, u1_u6_u7_n176, u1_u6_u7_n177, u1_u6_u7_n178, u1_u6_u7_n179, u1_u6_u7_n180, u1_u6_u7_n91, u1_u6_u7_n92, 
       u1_u6_u7_n93, u1_u6_u7_n94, u1_u6_u7_n95, u1_u6_u7_n96, u1_u6_u7_n97, u1_u6_u7_n98, u1_u6_u7_n99, u1_u8_X_1, u1_u8_X_19, 
       u1_u8_X_2, u1_u8_X_20, u1_u8_X_22, u1_u8_X_23, u1_u8_X_24, u1_u8_X_25, u1_u8_X_26, u1_u8_X_27, u1_u8_X_29, 
       u1_u8_X_31, u1_u8_X_35, u1_u8_X_36, u1_u8_X_37, u1_u8_X_38, u1_u8_X_41, u1_u8_X_42, u1_u8_X_43, u1_u8_X_44, 
       u1_u8_X_47, u1_u8_X_48, u1_u8_X_5, u1_u8_X_6, u1_u8_u0_n100, u1_u8_u0_n101, u1_u8_u0_n102, u1_u8_u0_n103, u1_u8_u0_n104, 
       u1_u8_u0_n105, u1_u8_u0_n106, u1_u8_u0_n107, u1_u8_u0_n108, u1_u8_u0_n109, u1_u8_u0_n110, u1_u8_u0_n111, u1_u8_u0_n112, u1_u8_u0_n113, 
       u1_u8_u0_n114, u1_u8_u0_n115, u1_u8_u0_n116, u1_u8_u0_n117, u1_u8_u0_n118, u1_u8_u0_n119, u1_u8_u0_n120, u1_u8_u0_n121, u1_u8_u0_n122, 
       u1_u8_u0_n123, u1_u8_u0_n124, u1_u8_u0_n125, u1_u8_u0_n126, u1_u8_u0_n127, u1_u8_u0_n128, u1_u8_u0_n129, u1_u8_u0_n130, u1_u8_u0_n131, 
       u1_u8_u0_n132, u1_u8_u0_n133, u1_u8_u0_n134, u1_u8_u0_n135, u1_u8_u0_n136, u1_u8_u0_n137, u1_u8_u0_n138, u1_u8_u0_n139, u1_u8_u0_n140, 
       u1_u8_u0_n141, u1_u8_u0_n142, u1_u8_u0_n143, u1_u8_u0_n144, u1_u8_u0_n145, u1_u8_u0_n146, u1_u8_u0_n147, u1_u8_u0_n148, u1_u8_u0_n149, 
       u1_u8_u0_n150, u1_u8_u0_n151, u1_u8_u0_n152, u1_u8_u0_n153, u1_u8_u0_n154, u1_u8_u0_n155, u1_u8_u0_n156, u1_u8_u0_n157, u1_u8_u0_n158, 
       u1_u8_u0_n159, u1_u8_u0_n160, u1_u8_u0_n161, u1_u8_u0_n162, u1_u8_u0_n163, u1_u8_u0_n164, u1_u8_u0_n165, u1_u8_u0_n166, u1_u8_u0_n167, 
       u1_u8_u0_n168, u1_u8_u0_n169, u1_u8_u0_n170, u1_u8_u0_n171, u1_u8_u0_n172, u1_u8_u0_n173, u1_u8_u0_n174, u1_u8_u0_n88, u1_u8_u0_n89, 
       u1_u8_u0_n90, u1_u8_u0_n91, u1_u8_u0_n92, u1_u8_u0_n93, u1_u8_u0_n94, u1_u8_u0_n95, u1_u8_u0_n96, u1_u8_u0_n97, u1_u8_u0_n98, 
       u1_u8_u0_n99, u1_u8_u3_n100, u1_u8_u3_n101, u1_u8_u3_n102, u1_u8_u3_n103, u1_u8_u3_n104, u1_u8_u3_n105, u1_u8_u3_n106, u1_u8_u3_n107, 
       u1_u8_u3_n108, u1_u8_u3_n109, u1_u8_u3_n110, u1_u8_u3_n111, u1_u8_u3_n112, u1_u8_u3_n113, u1_u8_u3_n114, u1_u8_u3_n115, u1_u8_u3_n116, 
       u1_u8_u3_n117, u1_u8_u3_n118, u1_u8_u3_n119, u1_u8_u3_n120, u1_u8_u3_n121, u1_u8_u3_n122, u1_u8_u3_n123, u1_u8_u3_n124, u1_u8_u3_n125, 
       u1_u8_u3_n126, u1_u8_u3_n127, u1_u8_u3_n128, u1_u8_u3_n129, u1_u8_u3_n130, u1_u8_u3_n131, u1_u8_u3_n132, u1_u8_u3_n133, u1_u8_u3_n134, 
       u1_u8_u3_n135, u1_u8_u3_n136, u1_u8_u3_n137, u1_u8_u3_n138, u1_u8_u3_n139, u1_u8_u3_n140, u1_u8_u3_n141, u1_u8_u3_n142, u1_u8_u3_n143, 
       u1_u8_u3_n144, u1_u8_u3_n145, u1_u8_u3_n146, u1_u8_u3_n147, u1_u8_u3_n148, u1_u8_u3_n149, u1_u8_u3_n150, u1_u8_u3_n151, u1_u8_u3_n152, 
       u1_u8_u3_n153, u1_u8_u3_n154, u1_u8_u3_n155, u1_u8_u3_n156, u1_u8_u3_n157, u1_u8_u3_n158, u1_u8_u3_n159, u1_u8_u3_n160, u1_u8_u3_n161, 
       u1_u8_u3_n162, u1_u8_u3_n163, u1_u8_u3_n164, u1_u8_u3_n165, u1_u8_u3_n166, u1_u8_u3_n167, u1_u8_u3_n168, u1_u8_u3_n169, u1_u8_u3_n170, 
       u1_u8_u3_n171, u1_u8_u3_n172, u1_u8_u3_n173, u1_u8_u3_n174, u1_u8_u3_n175, u1_u8_u3_n176, u1_u8_u3_n177, u1_u8_u3_n178, u1_u8_u3_n179, 
       u1_u8_u3_n180, u1_u8_u3_n181, u1_u8_u3_n182, u1_u8_u3_n183, u1_u8_u3_n184, u1_u8_u3_n185, u1_u8_u3_n186, u1_u8_u3_n94, u1_u8_u3_n95, 
       u1_u8_u3_n96, u1_u8_u3_n97, u1_u8_u3_n98, u1_u8_u3_n99, u1_u8_u4_n100, u1_u8_u4_n101, u1_u8_u4_n102, u1_u8_u4_n103, u1_u8_u4_n104, 
       u1_u8_u4_n105, u1_u8_u4_n106, u1_u8_u4_n107, u1_u8_u4_n108, u1_u8_u4_n109, u1_u8_u4_n110, u1_u8_u4_n111, u1_u8_u4_n112, u1_u8_u4_n113, 
       u1_u8_u4_n114, u1_u8_u4_n115, u1_u8_u4_n116, u1_u8_u4_n117, u1_u8_u4_n118, u1_u8_u4_n119, u1_u8_u4_n120, u1_u8_u4_n121, u1_u8_u4_n122, 
       u1_u8_u4_n123, u1_u8_u4_n124, u1_u8_u4_n125, u1_u8_u4_n126, u1_u8_u4_n127, u1_u8_u4_n128, u1_u8_u4_n129, u1_u8_u4_n130, u1_u8_u4_n131, 
       u1_u8_u4_n132, u1_u8_u4_n133, u1_u8_u4_n134, u1_u8_u4_n135, u1_u8_u4_n136, u1_u8_u4_n137, u1_u8_u4_n138, u1_u8_u4_n139, u1_u8_u4_n140, 
       u1_u8_u4_n141, u1_u8_u4_n142, u1_u8_u4_n143, u1_u8_u4_n144, u1_u8_u4_n145, u1_u8_u4_n146, u1_u8_u4_n147, u1_u8_u4_n148, u1_u8_u4_n149, 
       u1_u8_u4_n150, u1_u8_u4_n151, u1_u8_u4_n152, u1_u8_u4_n153, u1_u8_u4_n154, u1_u8_u4_n155, u1_u8_u4_n156, u1_u8_u4_n157, u1_u8_u4_n158, 
       u1_u8_u4_n159, u1_u8_u4_n160, u1_u8_u4_n161, u1_u8_u4_n162, u1_u8_u4_n163, u1_u8_u4_n164, u1_u8_u4_n165, u1_u8_u4_n166, u1_u8_u4_n167, 
       u1_u8_u4_n168, u1_u8_u4_n169, u1_u8_u4_n170, u1_u8_u4_n171, u1_u8_u4_n172, u1_u8_u4_n173, u1_u8_u4_n174, u1_u8_u4_n175, u1_u8_u4_n176, 
       u1_u8_u4_n177, u1_u8_u4_n178, u1_u8_u4_n179, u1_u8_u4_n180, u1_u8_u4_n181, u1_u8_u4_n182, u1_u8_u4_n183, u1_u8_u4_n184, u1_u8_u4_n185, 
       u1_u8_u4_n186, u1_u8_u4_n94, u1_u8_u4_n95, u1_u8_u4_n96, u1_u8_u4_n97, u1_u8_u4_n98, u1_u8_u4_n99, u1_u8_u5_n100, u1_u8_u5_n101, 
       u1_u8_u5_n102, u1_u8_u5_n103, u1_u8_u5_n104, u1_u8_u5_n105, u1_u8_u5_n106, u1_u8_u5_n107, u1_u8_u5_n108, u1_u8_u5_n109, u1_u8_u5_n110, 
       u1_u8_u5_n111, u1_u8_u5_n112, u1_u8_u5_n113, u1_u8_u5_n114, u1_u8_u5_n115, u1_u8_u5_n116, u1_u8_u5_n117, u1_u8_u5_n118, u1_u8_u5_n119, 
       u1_u8_u5_n120, u1_u8_u5_n121, u1_u8_u5_n122, u1_u8_u5_n123, u1_u8_u5_n124, u1_u8_u5_n125, u1_u8_u5_n126, u1_u8_u5_n127, u1_u8_u5_n128, 
       u1_u8_u5_n129, u1_u8_u5_n130, u1_u8_u5_n131, u1_u8_u5_n132, u1_u8_u5_n133, u1_u8_u5_n134, u1_u8_u5_n135, u1_u8_u5_n136, u1_u8_u5_n137, 
       u1_u8_u5_n138, u1_u8_u5_n139, u1_u8_u5_n140, u1_u8_u5_n141, u1_u8_u5_n142, u1_u8_u5_n143, u1_u8_u5_n144, u1_u8_u5_n145, u1_u8_u5_n146, 
       u1_u8_u5_n147, u1_u8_u5_n148, u1_u8_u5_n149, u1_u8_u5_n150, u1_u8_u5_n151, u1_u8_u5_n152, u1_u8_u5_n153, u1_u8_u5_n154, u1_u8_u5_n155, 
       u1_u8_u5_n156, u1_u8_u5_n157, u1_u8_u5_n158, u1_u8_u5_n159, u1_u8_u5_n160, u1_u8_u5_n161, u1_u8_u5_n162, u1_u8_u5_n163, u1_u8_u5_n164, 
       u1_u8_u5_n165, u1_u8_u5_n166, u1_u8_u5_n167, u1_u8_u5_n168, u1_u8_u5_n169, u1_u8_u5_n170, u1_u8_u5_n171, u1_u8_u5_n172, u1_u8_u5_n173, 
       u1_u8_u5_n174, u1_u8_u5_n175, u1_u8_u5_n176, u1_u8_u5_n177, u1_u8_u5_n178, u1_u8_u5_n179, u1_u8_u5_n180, u1_u8_u5_n181, u1_u8_u5_n182, 
       u1_u8_u5_n183, u1_u8_u5_n184, u1_u8_u5_n185, u1_u8_u5_n186, u1_u8_u5_n187, u1_u8_u5_n188, u1_u8_u5_n189, u1_u8_u5_n190, u1_u8_u5_n191, 
       u1_u8_u5_n192, u1_u8_u5_n193, u1_u8_u5_n194, u1_u8_u5_n195, u1_u8_u5_n196, u1_u8_u5_n99, u1_u8_u6_n100, u1_u8_u6_n101, u1_u8_u6_n102, 
       u1_u8_u6_n103, u1_u8_u6_n104, u1_u8_u6_n105, u1_u8_u6_n106, u1_u8_u6_n107, u1_u8_u6_n108, u1_u8_u6_n109, u1_u8_u6_n110, u1_u8_u6_n111, 
       u1_u8_u6_n112, u1_u8_u6_n113, u1_u8_u6_n114, u1_u8_u6_n115, u1_u8_u6_n116, u1_u8_u6_n117, u1_u8_u6_n118, u1_u8_u6_n119, u1_u8_u6_n120, 
       u1_u8_u6_n121, u1_u8_u6_n122, u1_u8_u6_n123, u1_u8_u6_n124, u1_u8_u6_n125, u1_u8_u6_n126, u1_u8_u6_n127, u1_u8_u6_n128, u1_u8_u6_n129, 
       u1_u8_u6_n130, u1_u8_u6_n131, u1_u8_u6_n132, u1_u8_u6_n133, u1_u8_u6_n134, u1_u8_u6_n135, u1_u8_u6_n136, u1_u8_u6_n137, u1_u8_u6_n138, 
       u1_u8_u6_n139, u1_u8_u6_n140, u1_u8_u6_n141, u1_u8_u6_n142, u1_u8_u6_n143, u1_u8_u6_n144, u1_u8_u6_n145, u1_u8_u6_n146, u1_u8_u6_n147, 
       u1_u8_u6_n148, u1_u8_u6_n149, u1_u8_u6_n150, u1_u8_u6_n151, u1_u8_u6_n152, u1_u8_u6_n153, u1_u8_u6_n154, u1_u8_u6_n155, u1_u8_u6_n156, 
       u1_u8_u6_n157, u1_u8_u6_n158, u1_u8_u6_n159, u1_u8_u6_n160, u1_u8_u6_n161, u1_u8_u6_n162, u1_u8_u6_n163, u1_u8_u6_n164, u1_u8_u6_n165, 
       u1_u8_u6_n166, u1_u8_u6_n167, u1_u8_u6_n168, u1_u8_u6_n169, u1_u8_u6_n170, u1_u8_u6_n171, u1_u8_u6_n172, u1_u8_u6_n173, u1_u8_u6_n174, 
       u1_u8_u6_n88, u1_u8_u6_n89, u1_u8_u6_n90, u1_u8_u6_n91, u1_u8_u6_n92, u1_u8_u6_n93, u1_u8_u6_n94, u1_u8_u6_n95, u1_u8_u6_n96, 
       u1_u8_u6_n97, u1_u8_u6_n98, u1_u8_u6_n99, u1_u8_u7_n100, u1_u8_u7_n101, u1_u8_u7_n102, u1_u8_u7_n103, u1_u8_u7_n104, u1_u8_u7_n105, 
       u1_u8_u7_n106, u1_u8_u7_n107, u1_u8_u7_n108, u1_u8_u7_n109, u1_u8_u7_n110, u1_u8_u7_n111, u1_u8_u7_n112, u1_u8_u7_n113, u1_u8_u7_n114, 
       u1_u8_u7_n115, u1_u8_u7_n116, u1_u8_u7_n117, u1_u8_u7_n118, u1_u8_u7_n119, u1_u8_u7_n120, u1_u8_u7_n121, u1_u8_u7_n122, u1_u8_u7_n123, 
       u1_u8_u7_n124, u1_u8_u7_n125, u1_u8_u7_n126, u1_u8_u7_n127, u1_u8_u7_n128, u1_u8_u7_n129, u1_u8_u7_n130, u1_u8_u7_n131, u1_u8_u7_n132, 
       u1_u8_u7_n133, u1_u8_u7_n134, u1_u8_u7_n135, u1_u8_u7_n136, u1_u8_u7_n137, u1_u8_u7_n138, u1_u8_u7_n139, u1_u8_u7_n140, u1_u8_u7_n141, 
       u1_u8_u7_n142, u1_u8_u7_n143, u1_u8_u7_n144, u1_u8_u7_n145, u1_u8_u7_n146, u1_u8_u7_n147, u1_u8_u7_n148, u1_u8_u7_n149, u1_u8_u7_n150, 
       u1_u8_u7_n151, u1_u8_u7_n152, u1_u8_u7_n153, u1_u8_u7_n154, u1_u8_u7_n155, u1_u8_u7_n156, u1_u8_u7_n157, u1_u8_u7_n158, u1_u8_u7_n159, 
       u1_u8_u7_n160, u1_u8_u7_n161, u1_u8_u7_n162, u1_u8_u7_n163, u1_u8_u7_n164, u1_u8_u7_n165, u1_u8_u7_n166, u1_u8_u7_n167, u1_u8_u7_n168, 
       u1_u8_u7_n169, u1_u8_u7_n170, u1_u8_u7_n171, u1_u8_u7_n172, u1_u8_u7_n173, u1_u8_u7_n174, u1_u8_u7_n175, u1_u8_u7_n176, u1_u8_u7_n177, 
       u1_u8_u7_n178, u1_u8_u7_n179, u1_u8_u7_n180, u1_u8_u7_n91, u1_u8_u7_n92, u1_u8_u7_n93, u1_u8_u7_n94, u1_u8_u7_n95, u1_u8_u7_n96, 
       u1_u8_u7_n97, u1_u8_u7_n98, u1_u8_u7_n99, u1_u9_X_31, u1_u9_X_32, u1_u9_X_33, u1_u9_X_35, u1_u9_X_36, u1_u9_X_37, 
       u1_u9_X_38, u1_u9_X_41, u1_u9_X_42, u1_u9_X_43, u1_u9_X_44, u1_u9_X_47, u1_u9_X_48, u1_u9_u5_n100, u1_u9_u5_n101, 
       u1_u9_u5_n102, u1_u9_u5_n103, u1_u9_u5_n104, u1_u9_u5_n105, u1_u9_u5_n106, u1_u9_u5_n107, u1_u9_u5_n108, u1_u9_u5_n109, u1_u9_u5_n110, 
       u1_u9_u5_n111, u1_u9_u5_n112, u1_u9_u5_n113, u1_u9_u5_n114, u1_u9_u5_n115, u1_u9_u5_n116, u1_u9_u5_n117, u1_u9_u5_n118, u1_u9_u5_n119, 
       u1_u9_u5_n120, u1_u9_u5_n121, u1_u9_u5_n122, u1_u9_u5_n123, u1_u9_u5_n124, u1_u9_u5_n125, u1_u9_u5_n126, u1_u9_u5_n127, u1_u9_u5_n128, 
       u1_u9_u5_n129, u1_u9_u5_n130, u1_u9_u5_n131, u1_u9_u5_n132, u1_u9_u5_n133, u1_u9_u5_n134, u1_u9_u5_n135, u1_u9_u5_n136, u1_u9_u5_n137, 
       u1_u9_u5_n138, u1_u9_u5_n139, u1_u9_u5_n140, u1_u9_u5_n141, u1_u9_u5_n142, u1_u9_u5_n143, u1_u9_u5_n144, u1_u9_u5_n145, u1_u9_u5_n146, 
       u1_u9_u5_n147, u1_u9_u5_n148, u1_u9_u5_n149, u1_u9_u5_n150, u1_u9_u5_n151, u1_u9_u5_n152, u1_u9_u5_n153, u1_u9_u5_n154, u1_u9_u5_n155, 
       u1_u9_u5_n156, u1_u9_u5_n157, u1_u9_u5_n158, u1_u9_u5_n159, u1_u9_u5_n160, u1_u9_u5_n161, u1_u9_u5_n162, u1_u9_u5_n163, u1_u9_u5_n164, 
       u1_u9_u5_n165, u1_u9_u5_n166, u1_u9_u5_n167, u1_u9_u5_n168, u1_u9_u5_n169, u1_u9_u5_n170, u1_u9_u5_n171, u1_u9_u5_n172, u1_u9_u5_n173, 
       u1_u9_u5_n174, u1_u9_u5_n175, u1_u9_u5_n176, u1_u9_u5_n177, u1_u9_u5_n178, u1_u9_u5_n179, u1_u9_u5_n180, u1_u9_u5_n181, u1_u9_u5_n182, 
       u1_u9_u5_n183, u1_u9_u5_n184, u1_u9_u5_n185, u1_u9_u5_n186, u1_u9_u5_n187, u1_u9_u5_n188, u1_u9_u5_n189, u1_u9_u5_n190, u1_u9_u5_n191, 
       u1_u9_u5_n192, u1_u9_u5_n193, u1_u9_u5_n194, u1_u9_u5_n195, u1_u9_u5_n196, u1_u9_u5_n99, u1_u9_u6_n100, u1_u9_u6_n101, u1_u9_u6_n102, 
       u1_u9_u6_n103, u1_u9_u6_n104, u1_u9_u6_n105, u1_u9_u6_n106, u1_u9_u6_n107, u1_u9_u6_n108, u1_u9_u6_n109, u1_u9_u6_n110, u1_u9_u6_n111, 
       u1_u9_u6_n112, u1_u9_u6_n113, u1_u9_u6_n114, u1_u9_u6_n115, u1_u9_u6_n116, u1_u9_u6_n117, u1_u9_u6_n118, u1_u9_u6_n119, u1_u9_u6_n120, 
       u1_u9_u6_n121, u1_u9_u6_n122, u1_u9_u6_n123, u1_u9_u6_n124, u1_u9_u6_n125, u1_u9_u6_n126, u1_u9_u6_n127, u1_u9_u6_n128, u1_u9_u6_n129, 
       u1_u9_u6_n130, u1_u9_u6_n131, u1_u9_u6_n132, u1_u9_u6_n133, u1_u9_u6_n134, u1_u9_u6_n135, u1_u9_u6_n136, u1_u9_u6_n137, u1_u9_u6_n138, 
       u1_u9_u6_n139, u1_u9_u6_n140, u1_u9_u6_n141, u1_u9_u6_n142, u1_u9_u6_n143, u1_u9_u6_n144, u1_u9_u6_n145, u1_u9_u6_n146, u1_u9_u6_n147, 
       u1_u9_u6_n148, u1_u9_u6_n149, u1_u9_u6_n150, u1_u9_u6_n151, u1_u9_u6_n152, u1_u9_u6_n153, u1_u9_u6_n154, u1_u9_u6_n155, u1_u9_u6_n156, 
       u1_u9_u6_n157, u1_u9_u6_n158, u1_u9_u6_n159, u1_u9_u6_n160, u1_u9_u6_n161, u1_u9_u6_n162, u1_u9_u6_n163, u1_u9_u6_n164, u1_u9_u6_n165, 
       u1_u9_u6_n166, u1_u9_u6_n167, u1_u9_u6_n168, u1_u9_u6_n169, u1_u9_u6_n170, u1_u9_u6_n171, u1_u9_u6_n172, u1_u9_u6_n173, u1_u9_u6_n174, 
       u1_u9_u6_n88, u1_u9_u6_n89, u1_u9_u6_n90, u1_u9_u6_n91, u1_u9_u6_n92, u1_u9_u6_n93, u1_u9_u6_n94, u1_u9_u6_n95, u1_u9_u6_n96, 
       u1_u9_u6_n97, u1_u9_u6_n98, u1_u9_u6_n99, u1_u9_u7_n100, u1_u9_u7_n101, u1_u9_u7_n102, u1_u9_u7_n103, u1_u9_u7_n104, u1_u9_u7_n105, 
       u1_u9_u7_n106, u1_u9_u7_n107, u1_u9_u7_n108, u1_u9_u7_n109, u1_u9_u7_n110, u1_u9_u7_n111, u1_u9_u7_n112, u1_u9_u7_n113, u1_u9_u7_n114, 
       u1_u9_u7_n115, u1_u9_u7_n116, u1_u9_u7_n117, u1_u9_u7_n118, u1_u9_u7_n119, u1_u9_u7_n120, u1_u9_u7_n121, u1_u9_u7_n122, u1_u9_u7_n123, 
       u1_u9_u7_n124, u1_u9_u7_n125, u1_u9_u7_n126, u1_u9_u7_n127, u1_u9_u7_n128, u1_u9_u7_n129, u1_u9_u7_n130, u1_u9_u7_n131, u1_u9_u7_n132, 
       u1_u9_u7_n133, u1_u9_u7_n134, u1_u9_u7_n135, u1_u9_u7_n136, u1_u9_u7_n137, u1_u9_u7_n138, u1_u9_u7_n139, u1_u9_u7_n140, u1_u9_u7_n141, 
       u1_u9_u7_n142, u1_u9_u7_n143, u1_u9_u7_n144, u1_u9_u7_n145, u1_u9_u7_n146, u1_u9_u7_n147, u1_u9_u7_n148, u1_u9_u7_n149, u1_u9_u7_n150, 
       u1_u9_u7_n151, u1_u9_u7_n152, u1_u9_u7_n153, u1_u9_u7_n154, u1_u9_u7_n155, u1_u9_u7_n156, u1_u9_u7_n157, u1_u9_u7_n158, u1_u9_u7_n159, 
       u1_u9_u7_n160, u1_u9_u7_n161, u1_u9_u7_n162, u1_u9_u7_n163, u1_u9_u7_n164, u1_u9_u7_n165, u1_u9_u7_n166, u1_u9_u7_n167, u1_u9_u7_n168, 
       u1_u9_u7_n169, u1_u9_u7_n170, u1_u9_u7_n171, u1_u9_u7_n172, u1_u9_u7_n173, u1_u9_u7_n174, u1_u9_u7_n175, u1_u9_u7_n176, u1_u9_u7_n177, 
       u1_u9_u7_n178, u1_u9_u7_n179, u1_u9_u7_n180, u1_u9_u7_n91, u1_u9_u7_n92, u1_u9_u7_n93, u1_u9_u7_n94, u1_u9_u7_n95, u1_u9_u7_n96, 
       u1_u9_u7_n97, u1_u9_u7_n98, u1_u9_u7_n99, u2_K11_12, u2_K11_14, u2_K11_17, u2_K16_29, u2_K16_34, u2_K16_37, 
       u2_K16_43, u2_K8_12, u2_K8_3, u2_K8_43, u2_K9_33, u2_K9_35, u2_K9_41, u2_K9_42, u2_K9_44, 
       u2_K9_48, u2_u10_X_11, u2_u10_X_12, u2_u10_X_13, u2_u10_X_14, u2_u10_X_17, u2_u10_u1_n100, u2_u10_u1_n101, u2_u10_u1_n102, 
       u2_u10_u1_n103, u2_u10_u1_n104, u2_u10_u1_n105, u2_u10_u1_n106, u2_u10_u1_n107, u2_u10_u1_n108, u2_u10_u1_n109, u2_u10_u1_n110, u2_u10_u1_n111, 
       u2_u10_u1_n112, u2_u10_u1_n113, u2_u10_u1_n114, u2_u10_u1_n115, u2_u10_u1_n116, u2_u10_u1_n117, u2_u10_u1_n118, u2_u10_u1_n119, u2_u10_u1_n120, 
       u2_u10_u1_n121, u2_u10_u1_n122, u2_u10_u1_n123, u2_u10_u1_n124, u2_u10_u1_n125, u2_u10_u1_n126, u2_u10_u1_n127, u2_u10_u1_n128, u2_u10_u1_n129, 
       u2_u10_u1_n130, u2_u10_u1_n131, u2_u10_u1_n132, u2_u10_u1_n133, u2_u10_u1_n134, u2_u10_u1_n135, u2_u10_u1_n136, u2_u10_u1_n137, u2_u10_u1_n138, 
       u2_u10_u1_n139, u2_u10_u1_n140, u2_u10_u1_n141, u2_u10_u1_n142, u2_u10_u1_n143, u2_u10_u1_n144, u2_u10_u1_n145, u2_u10_u1_n146, u2_u10_u1_n147, 
       u2_u10_u1_n148, u2_u10_u1_n149, u2_u10_u1_n150, u2_u10_u1_n151, u2_u10_u1_n152, u2_u10_u1_n153, u2_u10_u1_n154, u2_u10_u1_n155, u2_u10_u1_n156, 
       u2_u10_u1_n157, u2_u10_u1_n158, u2_u10_u1_n159, u2_u10_u1_n160, u2_u10_u1_n161, u2_u10_u1_n162, u2_u10_u1_n163, u2_u10_u1_n164, u2_u10_u1_n165, 
       u2_u10_u1_n166, u2_u10_u1_n167, u2_u10_u1_n168, u2_u10_u1_n169, u2_u10_u1_n170, u2_u10_u1_n171, u2_u10_u1_n172, u2_u10_u1_n173, u2_u10_u1_n174, 
       u2_u10_u1_n175, u2_u10_u1_n176, u2_u10_u1_n177, u2_u10_u1_n178, u2_u10_u1_n179, u2_u10_u1_n180, u2_u10_u1_n181, u2_u10_u1_n182, u2_u10_u1_n183, 
       u2_u10_u1_n184, u2_u10_u1_n185, u2_u10_u1_n186, u2_u10_u1_n187, u2_u10_u1_n188, u2_u10_u1_n95, u2_u10_u1_n96, u2_u10_u1_n97, u2_u10_u1_n98, 
       u2_u10_u1_n99, u2_u10_u2_n100, u2_u10_u2_n101, u2_u10_u2_n102, u2_u10_u2_n103, u2_u10_u2_n104, u2_u10_u2_n105, u2_u10_u2_n106, u2_u10_u2_n107, 
       u2_u10_u2_n108, u2_u10_u2_n109, u2_u10_u2_n110, u2_u10_u2_n111, u2_u10_u2_n112, u2_u10_u2_n113, u2_u10_u2_n114, u2_u10_u2_n115, u2_u10_u2_n116, 
       u2_u10_u2_n117, u2_u10_u2_n118, u2_u10_u2_n119, u2_u10_u2_n120, u2_u10_u2_n121, u2_u10_u2_n122, u2_u10_u2_n123, u2_u10_u2_n124, u2_u10_u2_n125, 
       u2_u10_u2_n126, u2_u10_u2_n127, u2_u10_u2_n128, u2_u10_u2_n129, u2_u10_u2_n130, u2_u10_u2_n131, u2_u10_u2_n132, u2_u10_u2_n133, u2_u10_u2_n134, 
       u2_u10_u2_n135, u2_u10_u2_n136, u2_u10_u2_n137, u2_u10_u2_n138, u2_u10_u2_n139, u2_u10_u2_n140, u2_u10_u2_n141, u2_u10_u2_n142, u2_u10_u2_n143, 
       u2_u10_u2_n144, u2_u10_u2_n145, u2_u10_u2_n146, u2_u10_u2_n147, u2_u10_u2_n148, u2_u10_u2_n149, u2_u10_u2_n150, u2_u10_u2_n151, u2_u10_u2_n152, 
       u2_u10_u2_n153, u2_u10_u2_n154, u2_u10_u2_n155, u2_u10_u2_n156, u2_u10_u2_n157, u2_u10_u2_n158, u2_u10_u2_n159, u2_u10_u2_n160, u2_u10_u2_n161, 
       u2_u10_u2_n162, u2_u10_u2_n163, u2_u10_u2_n164, u2_u10_u2_n165, u2_u10_u2_n166, u2_u10_u2_n167, u2_u10_u2_n168, u2_u10_u2_n169, u2_u10_u2_n170, 
       u2_u10_u2_n171, u2_u10_u2_n172, u2_u10_u2_n173, u2_u10_u2_n174, u2_u10_u2_n175, u2_u10_u2_n176, u2_u10_u2_n177, u2_u10_u2_n178, u2_u10_u2_n179, 
       u2_u10_u2_n180, u2_u10_u2_n181, u2_u10_u2_n182, u2_u10_u2_n183, u2_u10_u2_n184, u2_u10_u2_n185, u2_u10_u2_n186, u2_u10_u2_n187, u2_u10_u2_n188, 
       u2_u10_u2_n95, u2_u10_u2_n96, u2_u10_u2_n97, u2_u10_u2_n98, u2_u10_u2_n99, u2_u15_X_1, u2_u15_X_11, u2_u15_X_12, u2_u15_X_13, 
       u2_u15_X_14, u2_u15_X_17, u2_u15_X_18, u2_u15_X_19, u2_u15_X_2, u2_u15_X_20, u2_u15_X_23, u2_u15_X_24, u2_u15_X_25, 
       u2_u15_X_26, u2_u15_X_29, u2_u15_X_30, u2_u15_X_31, u2_u15_X_32, u2_u15_X_34, u2_u15_X_35, u2_u15_X_36, u2_u15_X_37, 
       u2_u15_X_38, u2_u15_X_41, u2_u15_X_42, u2_u15_X_43, u2_u15_X_44, u2_u15_X_47, u2_u15_X_48, u2_u15_X_5, u2_u15_X_6, 
       u2_u15_X_7, u2_u15_X_8, u2_u15_u0_n100, u2_u15_u0_n101, u2_u15_u0_n102, u2_u15_u0_n103, u2_u15_u0_n104, u2_u15_u0_n105, u2_u15_u0_n106, 
       u2_u15_u0_n107, u2_u15_u0_n108, u2_u15_u0_n109, u2_u15_u0_n110, u2_u15_u0_n111, u2_u15_u0_n112, u2_u15_u0_n113, u2_u15_u0_n114, u2_u15_u0_n115, 
       u2_u15_u0_n116, u2_u15_u0_n117, u2_u15_u0_n118, u2_u15_u0_n119, u2_u15_u0_n120, u2_u15_u0_n121, u2_u15_u0_n122, u2_u15_u0_n123, u2_u15_u0_n124, 
       u2_u15_u0_n125, u2_u15_u0_n126, u2_u15_u0_n127, u2_u15_u0_n128, u2_u15_u0_n129, u2_u15_u0_n130, u2_u15_u0_n131, u2_u15_u0_n132, u2_u15_u0_n133, 
       u2_u15_u0_n134, u2_u15_u0_n135, u2_u15_u0_n136, u2_u15_u0_n137, u2_u15_u0_n138, u2_u15_u0_n139, u2_u15_u0_n140, u2_u15_u0_n141, u2_u15_u0_n142, 
       u2_u15_u0_n143, u2_u15_u0_n144, u2_u15_u0_n145, u2_u15_u0_n146, u2_u15_u0_n147, u2_u15_u0_n148, u2_u15_u0_n149, u2_u15_u0_n150, u2_u15_u0_n151, 
       u2_u15_u0_n152, u2_u15_u0_n153, u2_u15_u0_n154, u2_u15_u0_n155, u2_u15_u0_n156, u2_u15_u0_n157, u2_u15_u0_n158, u2_u15_u0_n159, u2_u15_u0_n160, 
       u2_u15_u0_n161, u2_u15_u0_n162, u2_u15_u0_n163, u2_u15_u0_n164, u2_u15_u0_n165, u2_u15_u0_n166, u2_u15_u0_n167, u2_u15_u0_n168, u2_u15_u0_n169, 
       u2_u15_u0_n170, u2_u15_u0_n171, u2_u15_u0_n172, u2_u15_u0_n173, u2_u15_u0_n174, u2_u15_u0_n88, u2_u15_u0_n89, u2_u15_u0_n90, u2_u15_u0_n91, 
       u2_u15_u0_n92, u2_u15_u0_n93, u2_u15_u0_n94, u2_u15_u0_n95, u2_u15_u0_n96, u2_u15_u0_n97, u2_u15_u0_n98, u2_u15_u0_n99, u2_u15_u1_n100, 
       u2_u15_u1_n101, u2_u15_u1_n102, u2_u15_u1_n103, u2_u15_u1_n104, u2_u15_u1_n105, u2_u15_u1_n106, u2_u15_u1_n107, u2_u15_u1_n108, u2_u15_u1_n109, 
       u2_u15_u1_n110, u2_u15_u1_n111, u2_u15_u1_n112, u2_u15_u1_n113, u2_u15_u1_n114, u2_u15_u1_n115, u2_u15_u1_n116, u2_u15_u1_n117, u2_u15_u1_n118, 
       u2_u15_u1_n119, u2_u15_u1_n120, u2_u15_u1_n121, u2_u15_u1_n122, u2_u15_u1_n123, u2_u15_u1_n124, u2_u15_u1_n125, u2_u15_u1_n126, u2_u15_u1_n127, 
       u2_u15_u1_n128, u2_u15_u1_n129, u2_u15_u1_n130, u2_u15_u1_n131, u2_u15_u1_n132, u2_u15_u1_n133, u2_u15_u1_n134, u2_u15_u1_n135, u2_u15_u1_n136, 
       u2_u15_u1_n137, u2_u15_u1_n138, u2_u15_u1_n139, u2_u15_u1_n140, u2_u15_u1_n141, u2_u15_u1_n142, u2_u15_u1_n143, u2_u15_u1_n144, u2_u15_u1_n145, 
       u2_u15_u1_n146, u2_u15_u1_n147, u2_u15_u1_n148, u2_u15_u1_n149, u2_u15_u1_n150, u2_u15_u1_n151, u2_u15_u1_n152, u2_u15_u1_n153, u2_u15_u1_n154, 
       u2_u15_u1_n155, u2_u15_u1_n156, u2_u15_u1_n157, u2_u15_u1_n158, u2_u15_u1_n159, u2_u15_u1_n160, u2_u15_u1_n161, u2_u15_u1_n162, u2_u15_u1_n163, 
       u2_u15_u1_n164, u2_u15_u1_n165, u2_u15_u1_n166, u2_u15_u1_n167, u2_u15_u1_n168, u2_u15_u1_n169, u2_u15_u1_n170, u2_u15_u1_n171, u2_u15_u1_n172, 
       u2_u15_u1_n173, u2_u15_u1_n174, u2_u15_u1_n175, u2_u15_u1_n176, u2_u15_u1_n177, u2_u15_u1_n178, u2_u15_u1_n179, u2_u15_u1_n180, u2_u15_u1_n181, 
       u2_u15_u1_n182, u2_u15_u1_n183, u2_u15_u1_n184, u2_u15_u1_n185, u2_u15_u1_n186, u2_u15_u1_n187, u2_u15_u1_n188, u2_u15_u1_n95, u2_u15_u1_n96, 
       u2_u15_u1_n97, u2_u15_u1_n98, u2_u15_u1_n99, u2_u15_u2_n100, u2_u15_u2_n101, u2_u15_u2_n102, u2_u15_u2_n103, u2_u15_u2_n104, u2_u15_u2_n105, 
       u2_u15_u2_n106, u2_u15_u2_n107, u2_u15_u2_n108, u2_u15_u2_n109, u2_u15_u2_n110, u2_u15_u2_n111, u2_u15_u2_n112, u2_u15_u2_n113, u2_u15_u2_n114, 
       u2_u15_u2_n115, u2_u15_u2_n116, u2_u15_u2_n117, u2_u15_u2_n118, u2_u15_u2_n119, u2_u15_u2_n120, u2_u15_u2_n121, u2_u15_u2_n122, u2_u15_u2_n123, 
       u2_u15_u2_n124, u2_u15_u2_n125, u2_u15_u2_n126, u2_u15_u2_n127, u2_u15_u2_n128, u2_u15_u2_n129, u2_u15_u2_n130, u2_u15_u2_n131, u2_u15_u2_n132, 
       u2_u15_u2_n133, u2_u15_u2_n134, u2_u15_u2_n135, u2_u15_u2_n136, u2_u15_u2_n137, u2_u15_u2_n138, u2_u15_u2_n139, u2_u15_u2_n140, u2_u15_u2_n141, 
       u2_u15_u2_n142, u2_u15_u2_n143, u2_u15_u2_n144, u2_u15_u2_n145, u2_u15_u2_n146, u2_u15_u2_n147, u2_u15_u2_n148, u2_u15_u2_n149, u2_u15_u2_n150, 
       u2_u15_u2_n151, u2_u15_u2_n152, u2_u15_u2_n153, u2_u15_u2_n154, u2_u15_u2_n155, u2_u15_u2_n156, u2_u15_u2_n157, u2_u15_u2_n158, u2_u15_u2_n159, 
       u2_u15_u2_n160, u2_u15_u2_n161, u2_u15_u2_n162, u2_u15_u2_n163, u2_u15_u2_n164, u2_u15_u2_n165, u2_u15_u2_n166, u2_u15_u2_n167, u2_u15_u2_n168, 
       u2_u15_u2_n169, u2_u15_u2_n170, u2_u15_u2_n171, u2_u15_u2_n172, u2_u15_u2_n173, u2_u15_u2_n174, u2_u15_u2_n175, u2_u15_u2_n176, u2_u15_u2_n177, 
       u2_u15_u2_n178, u2_u15_u2_n179, u2_u15_u2_n180, u2_u15_u2_n181, u2_u15_u2_n182, u2_u15_u2_n183, u2_u15_u2_n184, u2_u15_u2_n185, u2_u15_u2_n186, 
       u2_u15_u2_n187, u2_u15_u2_n188, u2_u15_u2_n95, u2_u15_u2_n96, u2_u15_u2_n97, u2_u15_u2_n98, u2_u15_u2_n99, u2_u15_u3_n100, u2_u15_u3_n101, 
       u2_u15_u3_n102, u2_u15_u3_n103, u2_u15_u3_n104, u2_u15_u3_n105, u2_u15_u3_n106, u2_u15_u3_n107, u2_u15_u3_n108, u2_u15_u3_n109, u2_u15_u3_n110, 
       u2_u15_u3_n111, u2_u15_u3_n112, u2_u15_u3_n113, u2_u15_u3_n114, u2_u15_u3_n115, u2_u15_u3_n116, u2_u15_u3_n117, u2_u15_u3_n118, u2_u15_u3_n119, 
       u2_u15_u3_n120, u2_u15_u3_n121, u2_u15_u3_n122, u2_u15_u3_n123, u2_u15_u3_n124, u2_u15_u3_n125, u2_u15_u3_n126, u2_u15_u3_n127, u2_u15_u3_n128, 
       u2_u15_u3_n129, u2_u15_u3_n130, u2_u15_u3_n131, u2_u15_u3_n132, u2_u15_u3_n133, u2_u15_u3_n134, u2_u15_u3_n135, u2_u15_u3_n136, u2_u15_u3_n137, 
       u2_u15_u3_n138, u2_u15_u3_n139, u2_u15_u3_n140, u2_u15_u3_n141, u2_u15_u3_n142, u2_u15_u3_n143, u2_u15_u3_n144, u2_u15_u3_n145, u2_u15_u3_n146, 
       u2_u15_u3_n147, u2_u15_u3_n148, u2_u15_u3_n149, u2_u15_u3_n150, u2_u15_u3_n151, u2_u15_u3_n152, u2_u15_u3_n153, u2_u15_u3_n154, u2_u15_u3_n155, 
       u2_u15_u3_n156, u2_u15_u3_n157, u2_u15_u3_n158, u2_u15_u3_n159, u2_u15_u3_n160, u2_u15_u3_n161, u2_u15_u3_n162, u2_u15_u3_n163, u2_u15_u3_n164, 
       u2_u15_u3_n165, u2_u15_u3_n166, u2_u15_u3_n167, u2_u15_u3_n168, u2_u15_u3_n169, u2_u15_u3_n170, u2_u15_u3_n171, u2_u15_u3_n172, u2_u15_u3_n173, 
       u2_u15_u3_n174, u2_u15_u3_n175, u2_u15_u3_n176, u2_u15_u3_n177, u2_u15_u3_n178, u2_u15_u3_n179, u2_u15_u3_n180, u2_u15_u3_n181, u2_u15_u3_n182, 
       u2_u15_u3_n183, u2_u15_u3_n184, u2_u15_u3_n185, u2_u15_u3_n186, u2_u15_u3_n94, u2_u15_u3_n95, u2_u15_u3_n96, u2_u15_u3_n97, u2_u15_u3_n98, 
       u2_u15_u3_n99, u2_u15_u4_n100, u2_u15_u4_n101, u2_u15_u4_n102, u2_u15_u4_n103, u2_u15_u4_n104, u2_u15_u4_n105, u2_u15_u4_n106, u2_u15_u4_n107, 
       u2_u15_u4_n108, u2_u15_u4_n109, u2_u15_u4_n110, u2_u15_u4_n111, u2_u15_u4_n112, u2_u15_u4_n113, u2_u15_u4_n114, u2_u15_u4_n115, u2_u15_u4_n116, 
       u2_u15_u4_n117, u2_u15_u4_n118, u2_u15_u4_n119, u2_u15_u4_n120, u2_u15_u4_n121, u2_u15_u4_n122, u2_u15_u4_n123, u2_u15_u4_n124, u2_u15_u4_n125, 
       u2_u15_u4_n126, u2_u15_u4_n127, u2_u15_u4_n128, u2_u15_u4_n129, u2_u15_u4_n130, u2_u15_u4_n131, u2_u15_u4_n132, u2_u15_u4_n133, u2_u15_u4_n134, 
       u2_u15_u4_n135, u2_u15_u4_n136, u2_u15_u4_n137, u2_u15_u4_n138, u2_u15_u4_n139, u2_u15_u4_n140, u2_u15_u4_n141, u2_u15_u4_n142, u2_u15_u4_n143, 
       u2_u15_u4_n144, u2_u15_u4_n145, u2_u15_u4_n146, u2_u15_u4_n147, u2_u15_u4_n148, u2_u15_u4_n149, u2_u15_u4_n150, u2_u15_u4_n151, u2_u15_u4_n152, 
       u2_u15_u4_n153, u2_u15_u4_n154, u2_u15_u4_n155, u2_u15_u4_n156, u2_u15_u4_n157, u2_u15_u4_n158, u2_u15_u4_n159, u2_u15_u4_n160, u2_u15_u4_n161, 
       u2_u15_u4_n162, u2_u15_u4_n163, u2_u15_u4_n164, u2_u15_u4_n165, u2_u15_u4_n166, u2_u15_u4_n167, u2_u15_u4_n168, u2_u15_u4_n169, u2_u15_u4_n170, 
       u2_u15_u4_n171, u2_u15_u4_n172, u2_u15_u4_n173, u2_u15_u4_n174, u2_u15_u4_n175, u2_u15_u4_n176, u2_u15_u4_n177, u2_u15_u4_n178, u2_u15_u4_n179, 
       u2_u15_u4_n180, u2_u15_u4_n181, u2_u15_u4_n182, u2_u15_u4_n183, u2_u15_u4_n184, u2_u15_u4_n185, u2_u15_u4_n186, u2_u15_u4_n94, u2_u15_u4_n95, 
       u2_u15_u4_n96, u2_u15_u4_n97, u2_u15_u4_n98, u2_u15_u4_n99, u2_u15_u5_n100, u2_u15_u5_n101, u2_u15_u5_n102, u2_u15_u5_n103, u2_u15_u5_n104, 
       u2_u15_u5_n105, u2_u15_u5_n106, u2_u15_u5_n107, u2_u15_u5_n108, u2_u15_u5_n109, u2_u15_u5_n110, u2_u15_u5_n111, u2_u15_u5_n112, u2_u15_u5_n113, 
       u2_u15_u5_n114, u2_u15_u5_n115, u2_u15_u5_n116, u2_u15_u5_n117, u2_u15_u5_n118, u2_u15_u5_n119, u2_u15_u5_n120, u2_u15_u5_n121, u2_u15_u5_n122, 
       u2_u15_u5_n123, u2_u15_u5_n124, u2_u15_u5_n125, u2_u15_u5_n126, u2_u15_u5_n127, u2_u15_u5_n128, u2_u15_u5_n129, u2_u15_u5_n130, u2_u15_u5_n131, 
       u2_u15_u5_n132, u2_u15_u5_n133, u2_u15_u5_n134, u2_u15_u5_n135, u2_u15_u5_n136, u2_u15_u5_n137, u2_u15_u5_n138, u2_u15_u5_n139, u2_u15_u5_n140, 
       u2_u15_u5_n141, u2_u15_u5_n142, u2_u15_u5_n143, u2_u15_u5_n144, u2_u15_u5_n145, u2_u15_u5_n146, u2_u15_u5_n147, u2_u15_u5_n148, u2_u15_u5_n149, 
       u2_u15_u5_n150, u2_u15_u5_n151, u2_u15_u5_n152, u2_u15_u5_n153, u2_u15_u5_n154, u2_u15_u5_n155, u2_u15_u5_n156, u2_u15_u5_n157, u2_u15_u5_n158, 
       u2_u15_u5_n159, u2_u15_u5_n160, u2_u15_u5_n161, u2_u15_u5_n162, u2_u15_u5_n163, u2_u15_u5_n164, u2_u15_u5_n165, u2_u15_u5_n166, u2_u15_u5_n167, 
       u2_u15_u5_n168, u2_u15_u5_n169, u2_u15_u5_n170, u2_u15_u5_n171, u2_u15_u5_n172, u2_u15_u5_n173, u2_u15_u5_n174, u2_u15_u5_n175, u2_u15_u5_n176, 
       u2_u15_u5_n177, u2_u15_u5_n178, u2_u15_u5_n179, u2_u15_u5_n180, u2_u15_u5_n181, u2_u15_u5_n182, u2_u15_u5_n183, u2_u15_u5_n184, u2_u15_u5_n185, 
       u2_u15_u5_n186, u2_u15_u5_n187, u2_u15_u5_n188, u2_u15_u5_n189, u2_u15_u5_n190, u2_u15_u5_n191, u2_u15_u5_n192, u2_u15_u5_n193, u2_u15_u5_n194, 
       u2_u15_u5_n195, u2_u15_u5_n196, u2_u15_u5_n99, u2_u15_u6_n100, u2_u15_u6_n101, u2_u15_u6_n102, u2_u15_u6_n103, u2_u15_u6_n104, u2_u15_u6_n105, 
       u2_u15_u6_n106, u2_u15_u6_n107, u2_u15_u6_n108, u2_u15_u6_n109, u2_u15_u6_n110, u2_u15_u6_n111, u2_u15_u6_n112, u2_u15_u6_n113, u2_u15_u6_n114, 
       u2_u15_u6_n115, u2_u15_u6_n116, u2_u15_u6_n117, u2_u15_u6_n118, u2_u15_u6_n119, u2_u15_u6_n120, u2_u15_u6_n121, u2_u15_u6_n122, u2_u15_u6_n123, 
       u2_u15_u6_n124, u2_u15_u6_n125, u2_u15_u6_n126, u2_u15_u6_n127, u2_u15_u6_n128, u2_u15_u6_n129, u2_u15_u6_n130, u2_u15_u6_n131, u2_u15_u6_n132, 
       u2_u15_u6_n133, u2_u15_u6_n134, u2_u15_u6_n135, u2_u15_u6_n136, u2_u15_u6_n137, u2_u15_u6_n138, u2_u15_u6_n139, u2_u15_u6_n140, u2_u15_u6_n141, 
       u2_u15_u6_n142, u2_u15_u6_n143, u2_u15_u6_n144, u2_u15_u6_n145, u2_u15_u6_n146, u2_u15_u6_n147, u2_u15_u6_n148, u2_u15_u6_n149, u2_u15_u6_n150, 
       u2_u15_u6_n151, u2_u15_u6_n152, u2_u15_u6_n153, u2_u15_u6_n154, u2_u15_u6_n155, u2_u15_u6_n156, u2_u15_u6_n157, u2_u15_u6_n158, u2_u15_u6_n159, 
       u2_u15_u6_n160, u2_u15_u6_n161, u2_u15_u6_n162, u2_u15_u6_n163, u2_u15_u6_n164, u2_u15_u6_n165, u2_u15_u6_n166, u2_u15_u6_n167, u2_u15_u6_n168, 
       u2_u15_u6_n169, u2_u15_u6_n170, u2_u15_u6_n171, u2_u15_u6_n172, u2_u15_u6_n173, u2_u15_u6_n174, u2_u15_u6_n88, u2_u15_u6_n89, u2_u15_u6_n90, 
       u2_u15_u6_n91, u2_u15_u6_n92, u2_u15_u6_n93, u2_u15_u6_n94, u2_u15_u6_n95, u2_u15_u6_n96, u2_u15_u6_n97, u2_u15_u6_n98, u2_u15_u6_n99, 
       u2_u15_u7_n100, u2_u15_u7_n101, u2_u15_u7_n102, u2_u15_u7_n103, u2_u15_u7_n104, u2_u15_u7_n105, u2_u15_u7_n106, u2_u15_u7_n107, u2_u15_u7_n108, 
       u2_u15_u7_n109, u2_u15_u7_n110, u2_u15_u7_n111, u2_u15_u7_n112, u2_u15_u7_n113, u2_u15_u7_n114, u2_u15_u7_n115, u2_u15_u7_n116, u2_u15_u7_n117, 
       u2_u15_u7_n118, u2_u15_u7_n119, u2_u15_u7_n120, u2_u15_u7_n121, u2_u15_u7_n122, u2_u15_u7_n123, u2_u15_u7_n124, u2_u15_u7_n125, u2_u15_u7_n126, 
       u2_u15_u7_n127, u2_u15_u7_n128, u2_u15_u7_n129, u2_u15_u7_n130, u2_u15_u7_n131, u2_u15_u7_n132, u2_u15_u7_n133, u2_u15_u7_n134, u2_u15_u7_n135, 
       u2_u15_u7_n136, u2_u15_u7_n137, u2_u15_u7_n138, u2_u15_u7_n139, u2_u15_u7_n140, u2_u15_u7_n141, u2_u15_u7_n142, u2_u15_u7_n143, u2_u15_u7_n144, 
       u2_u15_u7_n145, u2_u15_u7_n146, u2_u15_u7_n147, u2_u15_u7_n148, u2_u15_u7_n149, u2_u15_u7_n150, u2_u15_u7_n151, u2_u15_u7_n152, u2_u15_u7_n153, 
       u2_u15_u7_n154, u2_u15_u7_n155, u2_u15_u7_n156, u2_u15_u7_n157, u2_u15_u7_n158, u2_u15_u7_n159, u2_u15_u7_n160, u2_u15_u7_n161, u2_u15_u7_n162, 
       u2_u15_u7_n163, u2_u15_u7_n164, u2_u15_u7_n165, u2_u15_u7_n166, u2_u15_u7_n167, u2_u15_u7_n168, u2_u15_u7_n169, u2_u15_u7_n170, u2_u15_u7_n171, 
       u2_u15_u7_n172, u2_u15_u7_n173, u2_u15_u7_n174, u2_u15_u7_n175, u2_u15_u7_n176, u2_u15_u7_n177, u2_u15_u7_n178, u2_u15_u7_n179, u2_u15_u7_n180, 
       u2_u15_u7_n91, u2_u15_u7_n92, u2_u15_u7_n93, u2_u15_u7_n94, u2_u15_u7_n95, u2_u15_u7_n96, u2_u15_u7_n97, u2_u15_u7_n98, u2_u15_u7_n99, 
       u2_u7_X_1, u2_u7_X_11, u2_u7_X_12, u2_u7_X_13, u2_u7_X_14, u2_u7_X_17, u2_u7_X_18, u2_u7_X_19, u2_u7_X_2, 
       u2_u7_X_20, u2_u7_X_3, u2_u7_X_43, u2_u7_X_47, u2_u7_X_48, u2_u7_X_5, u2_u7_X_6, u2_u7_X_7, u2_u7_X_8, 
       u2_u7_u0_n100, u2_u7_u0_n101, u2_u7_u0_n102, u2_u7_u0_n103, u2_u7_u0_n104, u2_u7_u0_n105, u2_u7_u0_n106, u2_u7_u0_n107, u2_u7_u0_n108, 
       u2_u7_u0_n109, u2_u7_u0_n110, u2_u7_u0_n111, u2_u7_u0_n112, u2_u7_u0_n113, u2_u7_u0_n114, u2_u7_u0_n115, u2_u7_u0_n116, u2_u7_u0_n117, 
       u2_u7_u0_n118, u2_u7_u0_n119, u2_u7_u0_n120, u2_u7_u0_n121, u2_u7_u0_n122, u2_u7_u0_n123, u2_u7_u0_n124, u2_u7_u0_n125, u2_u7_u0_n126, 
       u2_u7_u0_n127, u2_u7_u0_n128, u2_u7_u0_n129, u2_u7_u0_n130, u2_u7_u0_n131, u2_u7_u0_n132, u2_u7_u0_n133, u2_u7_u0_n134, u2_u7_u0_n135, 
       u2_u7_u0_n136, u2_u7_u0_n137, u2_u7_u0_n138, u2_u7_u0_n139, u2_u7_u0_n140, u2_u7_u0_n141, u2_u7_u0_n142, u2_u7_u0_n143, u2_u7_u0_n144, 
       u2_u7_u0_n145, u2_u7_u0_n146, u2_u7_u0_n147, u2_u7_u0_n148, u2_u7_u0_n149, u2_u7_u0_n150, u2_u7_u0_n151, u2_u7_u0_n152, u2_u7_u0_n153, 
       u2_u7_u0_n154, u2_u7_u0_n155, u2_u7_u0_n156, u2_u7_u0_n157, u2_u7_u0_n158, u2_u7_u0_n159, u2_u7_u0_n160, u2_u7_u0_n161, u2_u7_u0_n162, 
       u2_u7_u0_n163, u2_u7_u0_n164, u2_u7_u0_n165, u2_u7_u0_n166, u2_u7_u0_n167, u2_u7_u0_n168, u2_u7_u0_n169, u2_u7_u0_n170, u2_u7_u0_n171, 
       u2_u7_u0_n172, u2_u7_u0_n173, u2_u7_u0_n174, u2_u7_u0_n88, u2_u7_u0_n89, u2_u7_u0_n90, u2_u7_u0_n91, u2_u7_u0_n92, u2_u7_u0_n93, 
       u2_u7_u0_n94, u2_u7_u0_n95, u2_u7_u0_n96, u2_u7_u0_n97, u2_u7_u0_n98, u2_u7_u0_n99, u2_u7_u1_n100, u2_u7_u1_n101, u2_u7_u1_n102, 
       u2_u7_u1_n103, u2_u7_u1_n104, u2_u7_u1_n105, u2_u7_u1_n106, u2_u7_u1_n107, u2_u7_u1_n108, u2_u7_u1_n109, u2_u7_u1_n110, u2_u7_u1_n111, 
       u2_u7_u1_n112, u2_u7_u1_n113, u2_u7_u1_n114, u2_u7_u1_n115, u2_u7_u1_n116, u2_u7_u1_n117, u2_u7_u1_n118, u2_u7_u1_n119, u2_u7_u1_n120, 
       u2_u7_u1_n121, u2_u7_u1_n122, u2_u7_u1_n123, u2_u7_u1_n124, u2_u7_u1_n125, u2_u7_u1_n126, u2_u7_u1_n127, u2_u7_u1_n128, u2_u7_u1_n129, 
       u2_u7_u1_n130, u2_u7_u1_n131, u2_u7_u1_n132, u2_u7_u1_n133, u2_u7_u1_n134, u2_u7_u1_n135, u2_u7_u1_n136, u2_u7_u1_n137, u2_u7_u1_n138, 
       u2_u7_u1_n139, u2_u7_u1_n140, u2_u7_u1_n141, u2_u7_u1_n142, u2_u7_u1_n143, u2_u7_u1_n144, u2_u7_u1_n145, u2_u7_u1_n146, u2_u7_u1_n147, 
       u2_u7_u1_n148, u2_u7_u1_n149, u2_u7_u1_n150, u2_u7_u1_n151, u2_u7_u1_n152, u2_u7_u1_n153, u2_u7_u1_n154, u2_u7_u1_n155, u2_u7_u1_n156, 
       u2_u7_u1_n157, u2_u7_u1_n158, u2_u7_u1_n159, u2_u7_u1_n160, u2_u7_u1_n161, u2_u7_u1_n162, u2_u7_u1_n163, u2_u7_u1_n164, u2_u7_u1_n165, 
       u2_u7_u1_n166, u2_u7_u1_n167, u2_u7_u1_n168, u2_u7_u1_n169, u2_u7_u1_n170, u2_u7_u1_n171, u2_u7_u1_n172, u2_u7_u1_n173, u2_u7_u1_n174, 
       u2_u7_u1_n175, u2_u7_u1_n176, u2_u7_u1_n177, u2_u7_u1_n178, u2_u7_u1_n179, u2_u7_u1_n180, u2_u7_u1_n181, u2_u7_u1_n182, u2_u7_u1_n183, 
       u2_u7_u1_n184, u2_u7_u1_n185, u2_u7_u1_n186, u2_u7_u1_n187, u2_u7_u1_n188, u2_u7_u1_n95, u2_u7_u1_n96, u2_u7_u1_n97, u2_u7_u1_n98, 
       u2_u7_u1_n99, u2_u7_u2_n100, u2_u7_u2_n101, u2_u7_u2_n102, u2_u7_u2_n103, u2_u7_u2_n104, u2_u7_u2_n105, u2_u7_u2_n106, u2_u7_u2_n107, 
       u2_u7_u2_n108, u2_u7_u2_n109, u2_u7_u2_n110, u2_u7_u2_n111, u2_u7_u2_n112, u2_u7_u2_n113, u2_u7_u2_n114, u2_u7_u2_n115, u2_u7_u2_n116, 
       u2_u7_u2_n117, u2_u7_u2_n118, u2_u7_u2_n119, u2_u7_u2_n120, u2_u7_u2_n121, u2_u7_u2_n122, u2_u7_u2_n123, u2_u7_u2_n124, u2_u7_u2_n125, 
       u2_u7_u2_n126, u2_u7_u2_n127, u2_u7_u2_n128, u2_u7_u2_n129, u2_u7_u2_n130, u2_u7_u2_n131, u2_u7_u2_n132, u2_u7_u2_n133, u2_u7_u2_n134, 
       u2_u7_u2_n135, u2_u7_u2_n136, u2_u7_u2_n137, u2_u7_u2_n138, u2_u7_u2_n139, u2_u7_u2_n140, u2_u7_u2_n141, u2_u7_u2_n142, u2_u7_u2_n143, 
       u2_u7_u2_n144, u2_u7_u2_n145, u2_u7_u2_n146, u2_u7_u2_n147, u2_u7_u2_n148, u2_u7_u2_n149, u2_u7_u2_n150, u2_u7_u2_n151, u2_u7_u2_n152, 
       u2_u7_u2_n153, u2_u7_u2_n154, u2_u7_u2_n155, u2_u7_u2_n156, u2_u7_u2_n157, u2_u7_u2_n158, u2_u7_u2_n159, u2_u7_u2_n160, u2_u7_u2_n161, 
       u2_u7_u2_n162, u2_u7_u2_n163, u2_u7_u2_n164, u2_u7_u2_n165, u2_u7_u2_n166, u2_u7_u2_n167, u2_u7_u2_n168, u2_u7_u2_n169, u2_u7_u2_n170, 
       u2_u7_u2_n171, u2_u7_u2_n172, u2_u7_u2_n173, u2_u7_u2_n174, u2_u7_u2_n175, u2_u7_u2_n176, u2_u7_u2_n177, u2_u7_u2_n178, u2_u7_u2_n179, 
       u2_u7_u2_n180, u2_u7_u2_n181, u2_u7_u2_n182, u2_u7_u2_n183, u2_u7_u2_n184, u2_u7_u2_n185, u2_u7_u2_n186, u2_u7_u2_n187, u2_u7_u2_n188, 
       u2_u7_u2_n95, u2_u7_u2_n96, u2_u7_u2_n97, u2_u7_u2_n98, u2_u7_u2_n99, u2_u7_u3_n100, u2_u7_u3_n101, u2_u7_u3_n102, u2_u7_u3_n103, 
       u2_u7_u3_n104, u2_u7_u3_n105, u2_u7_u3_n106, u2_u7_u3_n107, u2_u7_u3_n108, u2_u7_u3_n109, u2_u7_u3_n110, u2_u7_u3_n111, u2_u7_u3_n112, 
       u2_u7_u3_n113, u2_u7_u3_n114, u2_u7_u3_n115, u2_u7_u3_n116, u2_u7_u3_n117, u2_u7_u3_n118, u2_u7_u3_n119, u2_u7_u3_n120, u2_u7_u3_n121, 
       u2_u7_u3_n122, u2_u7_u3_n123, u2_u7_u3_n124, u2_u7_u3_n125, u2_u7_u3_n126, u2_u7_u3_n127, u2_u7_u3_n128, u2_u7_u3_n129, u2_u7_u3_n130, 
       u2_u7_u3_n131, u2_u7_u3_n132, u2_u7_u3_n133, u2_u7_u3_n134, u2_u7_u3_n135, u2_u7_u3_n136, u2_u7_u3_n137, u2_u7_u3_n138, u2_u7_u3_n139, 
       u2_u7_u3_n140, u2_u7_u3_n141, u2_u7_u3_n142, u2_u7_u3_n143, u2_u7_u3_n144, u2_u7_u3_n145, u2_u7_u3_n146, u2_u7_u3_n147, u2_u7_u3_n148, 
       u2_u7_u3_n149, u2_u7_u3_n150, u2_u7_u3_n151, u2_u7_u3_n152, u2_u7_u3_n153, u2_u7_u3_n154, u2_u7_u3_n155, u2_u7_u3_n156, u2_u7_u3_n157, 
       u2_u7_u3_n158, u2_u7_u3_n159, u2_u7_u3_n160, u2_u7_u3_n161, u2_u7_u3_n162, u2_u7_u3_n163, u2_u7_u3_n164, u2_u7_u3_n165, u2_u7_u3_n166, 
       u2_u7_u3_n167, u2_u7_u3_n168, u2_u7_u3_n169, u2_u7_u3_n170, u2_u7_u3_n171, u2_u7_u3_n172, u2_u7_u3_n173, u2_u7_u3_n174, u2_u7_u3_n175, 
       u2_u7_u3_n176, u2_u7_u3_n177, u2_u7_u3_n178, u2_u7_u3_n179, u2_u7_u3_n180, u2_u7_u3_n181, u2_u7_u3_n182, u2_u7_u3_n183, u2_u7_u3_n184, 
       u2_u7_u3_n185, u2_u7_u3_n186, u2_u7_u3_n94, u2_u7_u3_n95, u2_u7_u3_n96, u2_u7_u3_n97, u2_u7_u3_n98, u2_u7_u3_n99, u2_u7_u7_n100, 
       u2_u7_u7_n101, u2_u7_u7_n102, u2_u7_u7_n103, u2_u7_u7_n104, u2_u7_u7_n105, u2_u7_u7_n106, u2_u7_u7_n107, u2_u7_u7_n108, u2_u7_u7_n109, 
       u2_u7_u7_n110, u2_u7_u7_n111, u2_u7_u7_n112, u2_u7_u7_n113, u2_u7_u7_n114, u2_u7_u7_n115, u2_u7_u7_n116, u2_u7_u7_n117, u2_u7_u7_n118, 
       u2_u7_u7_n119, u2_u7_u7_n120, u2_u7_u7_n121, u2_u7_u7_n122, u2_u7_u7_n123, u2_u7_u7_n124, u2_u7_u7_n125, u2_u7_u7_n126, u2_u7_u7_n127, 
       u2_u7_u7_n128, u2_u7_u7_n129, u2_u7_u7_n130, u2_u7_u7_n131, u2_u7_u7_n132, u2_u7_u7_n133, u2_u7_u7_n134, u2_u7_u7_n135, u2_u7_u7_n136, 
       u2_u7_u7_n137, u2_u7_u7_n138, u2_u7_u7_n139, u2_u7_u7_n140, u2_u7_u7_n141, u2_u7_u7_n142, u2_u7_u7_n143, u2_u7_u7_n144, u2_u7_u7_n145, 
       u2_u7_u7_n146, u2_u7_u7_n147, u2_u7_u7_n148, u2_u7_u7_n149, u2_u7_u7_n150, u2_u7_u7_n151, u2_u7_u7_n152, u2_u7_u7_n153, u2_u7_u7_n154, 
       u2_u7_u7_n155, u2_u7_u7_n156, u2_u7_u7_n157, u2_u7_u7_n158, u2_u7_u7_n159, u2_u7_u7_n160, u2_u7_u7_n161, u2_u7_u7_n162, u2_u7_u7_n163, 
       u2_u7_u7_n164, u2_u7_u7_n165, u2_u7_u7_n166, u2_u7_u7_n167, u2_u7_u7_n168, u2_u7_u7_n169, u2_u7_u7_n170, u2_u7_u7_n171, u2_u7_u7_n172, 
       u2_u7_u7_n173, u2_u7_u7_n174, u2_u7_u7_n175, u2_u7_u7_n176, u2_u7_u7_n177, u2_u7_u7_n178, u2_u7_u7_n179, u2_u7_u7_n180, u2_u7_u7_n91, 
       u2_u7_u7_n92, u2_u7_u7_n93, u2_u7_u7_n94, u2_u7_u7_n95, u2_u7_u7_n96, u2_u7_u7_n97, u2_u7_u7_n98, u2_u7_u7_n99, u2_u8_X_33, 
       u2_u8_X_35, u2_u8_X_36, u2_u8_X_37, u2_u8_X_38, u2_u8_X_41, u2_u8_X_42, u2_u8_X_43, u2_u8_X_44, u2_u8_X_48, 
       u2_u8_u5_n100, u2_u8_u5_n101, u2_u8_u5_n102, u2_u8_u5_n103, u2_u8_u5_n104, u2_u8_u5_n105, u2_u8_u5_n106, u2_u8_u5_n107, u2_u8_u5_n108, 
       u2_u8_u5_n109, u2_u8_u5_n110, u2_u8_u5_n111, u2_u8_u5_n112, u2_u8_u5_n113, u2_u8_u5_n114, u2_u8_u5_n115, u2_u8_u5_n116, u2_u8_u5_n117, 
       u2_u8_u5_n118, u2_u8_u5_n119, u2_u8_u5_n120, u2_u8_u5_n121, u2_u8_u5_n122, u2_u8_u5_n123, u2_u8_u5_n124, u2_u8_u5_n125, u2_u8_u5_n126, 
       u2_u8_u5_n127, u2_u8_u5_n128, u2_u8_u5_n129, u2_u8_u5_n130, u2_u8_u5_n131, u2_u8_u5_n132, u2_u8_u5_n133, u2_u8_u5_n134, u2_u8_u5_n135, 
       u2_u8_u5_n136, u2_u8_u5_n137, u2_u8_u5_n138, u2_u8_u5_n139, u2_u8_u5_n140, u2_u8_u5_n141, u2_u8_u5_n142, u2_u8_u5_n143, u2_u8_u5_n144, 
       u2_u8_u5_n145, u2_u8_u5_n146, u2_u8_u5_n147, u2_u8_u5_n148, u2_u8_u5_n149, u2_u8_u5_n150, u2_u8_u5_n151, u2_u8_u5_n152, u2_u8_u5_n153, 
       u2_u8_u5_n154, u2_u8_u5_n155, u2_u8_u5_n156, u2_u8_u5_n157, u2_u8_u5_n158, u2_u8_u5_n159, u2_u8_u5_n160, u2_u8_u5_n161, u2_u8_u5_n162, 
       u2_u8_u5_n163, u2_u8_u5_n164, u2_u8_u5_n165, u2_u8_u5_n166, u2_u8_u5_n167, u2_u8_u5_n168, u2_u8_u5_n169, u2_u8_u5_n170, u2_u8_u5_n171, 
       u2_u8_u5_n172, u2_u8_u5_n173, u2_u8_u5_n174, u2_u8_u5_n175, u2_u8_u5_n176, u2_u8_u5_n177, u2_u8_u5_n178, u2_u8_u5_n179, u2_u8_u5_n180, 
       u2_u8_u5_n181, u2_u8_u5_n182, u2_u8_u5_n183, u2_u8_u5_n184, u2_u8_u5_n185, u2_u8_u5_n186, u2_u8_u5_n187, u2_u8_u5_n188, u2_u8_u5_n189, 
       u2_u8_u5_n190, u2_u8_u5_n191, u2_u8_u5_n192, u2_u8_u5_n193, u2_u8_u5_n194, u2_u8_u5_n195, u2_u8_u5_n196, u2_u8_u5_n99, u2_u8_u6_n100, 
       u2_u8_u6_n101, u2_u8_u6_n102, u2_u8_u6_n103, u2_u8_u6_n104, u2_u8_u6_n105, u2_u8_u6_n106, u2_u8_u6_n107, u2_u8_u6_n108, u2_u8_u6_n109, 
       u2_u8_u6_n110, u2_u8_u6_n111, u2_u8_u6_n112, u2_u8_u6_n113, u2_u8_u6_n114, u2_u8_u6_n115, u2_u8_u6_n116, u2_u8_u6_n117, u2_u8_u6_n118, 
       u2_u8_u6_n119, u2_u8_u6_n120, u2_u8_u6_n121, u2_u8_u6_n122, u2_u8_u6_n123, u2_u8_u6_n124, u2_u8_u6_n125, u2_u8_u6_n126, u2_u8_u6_n127, 
       u2_u8_u6_n128, u2_u8_u6_n129, u2_u8_u6_n130, u2_u8_u6_n131, u2_u8_u6_n132, u2_u8_u6_n133, u2_u8_u6_n134, u2_u8_u6_n135, u2_u8_u6_n136, 
       u2_u8_u6_n137, u2_u8_u6_n138, u2_u8_u6_n139, u2_u8_u6_n140, u2_u8_u6_n141, u2_u8_u6_n142, u2_u8_u6_n143, u2_u8_u6_n144, u2_u8_u6_n145, 
       u2_u8_u6_n146, u2_u8_u6_n147, u2_u8_u6_n148, u2_u8_u6_n149, u2_u8_u6_n150, u2_u8_u6_n151, u2_u8_u6_n152, u2_u8_u6_n153, u2_u8_u6_n154, 
       u2_u8_u6_n155, u2_u8_u6_n156, u2_u8_u6_n157, u2_u8_u6_n158, u2_u8_u6_n159, u2_u8_u6_n160, u2_u8_u6_n161, u2_u8_u6_n162, u2_u8_u6_n163, 
       u2_u8_u6_n164, u2_u8_u6_n165, u2_u8_u6_n166, u2_u8_u6_n167, u2_u8_u6_n168, u2_u8_u6_n169, u2_u8_u6_n170, u2_u8_u6_n171, u2_u8_u6_n172, 
       u2_u8_u6_n173, u2_u8_u6_n174, u2_u8_u6_n88, u2_u8_u6_n89, u2_u8_u6_n90, u2_u8_u6_n91, u2_u8_u6_n92, u2_u8_u6_n93, u2_u8_u6_n94, 
       u2_u8_u6_n95, u2_u8_u6_n96, u2_u8_u6_n97, u2_u8_u6_n98, u2_u8_u6_n99, u2_u8_u7_n100, u2_u8_u7_n101, u2_u8_u7_n102, u2_u8_u7_n103, 
       u2_u8_u7_n104, u2_u8_u7_n105, u2_u8_u7_n106, u2_u8_u7_n107, u2_u8_u7_n108, u2_u8_u7_n109, u2_u8_u7_n110, u2_u8_u7_n111, u2_u8_u7_n112, 
       u2_u8_u7_n113, u2_u8_u7_n114, u2_u8_u7_n115, u2_u8_u7_n116, u2_u8_u7_n117, u2_u8_u7_n118, u2_u8_u7_n119, u2_u8_u7_n120, u2_u8_u7_n121, 
       u2_u8_u7_n122, u2_u8_u7_n123, u2_u8_u7_n124, u2_u8_u7_n125, u2_u8_u7_n126, u2_u8_u7_n127, u2_u8_u7_n128, u2_u8_u7_n129, u2_u8_u7_n130, 
       u2_u8_u7_n131, u2_u8_u7_n132, u2_u8_u7_n133, u2_u8_u7_n134, u2_u8_u7_n135, u2_u8_u7_n136, u2_u8_u7_n137, u2_u8_u7_n138, u2_u8_u7_n139, 
       u2_u8_u7_n140, u2_u8_u7_n141, u2_u8_u7_n142, u2_u8_u7_n143, u2_u8_u7_n144, u2_u8_u7_n145, u2_u8_u7_n146, u2_u8_u7_n147, u2_u8_u7_n148, 
       u2_u8_u7_n149, u2_u8_u7_n150, u2_u8_u7_n151, u2_u8_u7_n152, u2_u8_u7_n153, u2_u8_u7_n154, u2_u8_u7_n155, u2_u8_u7_n156, u2_u8_u7_n157, 
       u2_u8_u7_n158, u2_u8_u7_n159, u2_u8_u7_n160, u2_u8_u7_n161, u2_u8_u7_n162, u2_u8_u7_n163, u2_u8_u7_n164, u2_u8_u7_n165, u2_u8_u7_n166, 
       u2_u8_u7_n167, u2_u8_u7_n168, u2_u8_u7_n169, u2_u8_u7_n170, u2_u8_u7_n171, u2_u8_u7_n172, u2_u8_u7_n173, u2_u8_u7_n174, u2_u8_u7_n175, 
       u2_u8_u7_n176, u2_u8_u7_n177, u2_u8_u7_n178, u2_u8_u7_n179, u2_u8_u7_n180, u2_u8_u7_n91, u2_u8_u7_n92, u2_u8_u7_n93, u2_u8_u7_n94, 
       u2_u8_u7_n95, u2_u8_u7_n96, u2_u8_u7_n97, u2_u8_u7_n98, u2_u8_u7_n99,  u2_uk_n1138;
  XOR2_X1 u0_u0_U1 (.B( u0_K1_9 ) , .A( u0_desIn_r_47 ) , .Z( u0_u0_X_9 ) );
  XOR2_X1 u0_u0_U16 (.B( u0_K1_3 ) , .A( u0_desIn_r_15 ) , .Z( u0_u0_X_3 ) );
  XOR2_X1 u0_u0_U2 (.B( u0_K1_8 ) , .A( u0_desIn_r_39 ) , .Z( u0_u0_X_8 ) );
  XOR2_X1 u0_u0_U27 (.B( u0_K1_2 ) , .A( u0_desIn_r_7 ) , .Z( u0_u0_X_2 ) );
  XOR2_X1 u0_u0_U3 (.B( u0_K1_7 ) , .A( u0_desIn_r_31 ) , .Z( u0_u0_X_7 ) );
  XOR2_X1 u0_u0_U33 (.B( u0_K1_24 ) , .A( u0_desIn_r_3 ) , .Z( u0_u0_X_24 ) );
  XOR2_X1 u0_u0_U37 (.B( u0_K1_20 ) , .A( u0_desIn_r_37 ) , .Z( u0_u0_X_20 ) );
  XOR2_X1 u0_u0_U38 (.B( u0_K1_1 ) , .A( u0_desIn_r_57 ) , .Z( u0_u0_X_1 ) );
  XOR2_X1 u0_u0_U39 (.B( u0_K1_19 ) , .A( u0_desIn_r_29 ) , .Z( u0_u0_X_19 ) );
  XOR2_X1 u0_u0_U4 (.B( u0_K1_6 ) , .A( u0_desIn_r_39 ) , .Z( u0_u0_X_6 ) );
  XOR2_X1 u0_u0_U40 (.B( u0_K1_18 ) , .A( u0_desIn_r_37 ) , .Z( u0_u0_X_18 ) );
  XOR2_X1 u0_u0_U41 (.B( u0_K1_17 ) , .A( u0_desIn_r_29 ) , .Z( u0_u0_X_17 ) );
  XOR2_X1 u0_u0_U44 (.B( u0_K1_14 ) , .A( u0_desIn_r_5 ) , .Z( u0_u0_X_14 ) );
  XOR2_X1 u0_u0_U45 (.B( u0_K1_13 ) , .A( u0_desIn_r_63 ) , .Z( u0_u0_X_13 ) );
  XOR2_X1 u0_u0_U46 (.B( u0_K1_12 ) , .A( u0_desIn_r_5 ) , .Z( u0_u0_X_12 ) );
  XOR2_X1 u0_u0_U47 (.B( u0_K1_11 ) , .A( u0_desIn_r_63 ) , .Z( u0_u0_X_11 ) );
  XOR2_X1 u0_u0_U48 (.B( u0_K1_10 ) , .A( u0_desIn_r_55 ) , .Z( u0_u0_X_10 ) );
  XOR2_X1 u0_u0_U5 (.B( u0_K1_5 ) , .A( u0_desIn_r_31 ) , .Z( u0_u0_X_5 ) );
  XOR2_X1 u0_u0_U6 (.B( u0_K1_4 ) , .A( u0_desIn_r_23 ) , .Z( u0_u0_X_4 ) );
  AND3_X1 u0_u0_u0_U10 (.A1( u0_u0_u0_n27 ) , .A3( u0_u0_u0_n45 ) , .ZN( u0_u0_u0_n48 ) , .A2( u0_u0_u0_n63 ) );
  NAND2_X1 u0_u0_u0_U11 (.A2( u0_u0_u0_n26 ) , .A1( u0_u0_u0_n36 ) , .ZN( u0_u0_u0_n62 ) );
  AND2_X1 u0_u0_u0_U12 (.A2( u0_u0_u0_n35 ) , .A1( u0_u0_u0_n45 ) , .ZN( u0_u0_u0_n68 ) );
  AND2_X1 u0_u0_u0_U13 (.ZN( u0_u0_u0_n24 ) , .A1( u0_u0_u0_n45 ) , .A2( u0_u0_u0_n46 ) );
  AND2_X1 u0_u0_u0_U14 (.ZN( u0_u0_u0_n30 ) , .A2( u0_u0_u0_n50 ) , .A1( u0_u0_u0_n67 ) );
  INV_X1 u0_u0_u0_U15 (.ZN( u0_u0_u0_n2 ) , .A( u0_u0_u0_n32 ) );
  NOR2_X1 u0_u0_u0_U16 (.A1( u0_u0_u0_n15 ) , .ZN( u0_u0_u0_n28 ) , .A2( u0_u0_u0_n39 ) );
  AOI21_X1 u0_u0_u0_U17 (.A( u0_u0_u0_n10 ) , .ZN( u0_u0_u0_n43 ) , .B1( u0_u0_u0_n72 ) , .B2( u0_u0_u0_n82 ) );
  INV_X1 u0_u0_u0_U18 (.ZN( u0_u0_u0_n10 ) , .A( u0_u0_u0_n33 ) );
  OAI22_X1 u0_u0_u0_U19 (.B2( u0_u0_u0_n28 ) , .A2( u0_u0_u0_n29 ) , .A1( u0_u0_u0_n37 ) , .ZN( u0_u0_u0_n49 ) , .B1( u0_u0_u0_n50 ) );
  OAI22_X1 u0_u0_u0_U20 (.B2( u0_u0_u0_n28 ) , .A1( u0_u0_u0_n31 ) , .B1( u0_u0_u0_n44 ) , .ZN( u0_u0_u0_n84 ) , .A2( u0_u0_u0_n85 ) );
  AND3_X1 u0_u0_u0_U21 (.A1( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n50 ) , .A3( u0_u0_u0_n54 ) , .ZN( u0_u0_u0_n85 ) );
  NAND2_X1 u0_u0_u0_U22 (.ZN( u0_u0_u0_n50 ) , .A2( u0_u0_u0_n72 ) , .A1( u0_u0_u0_n75 ) );
  INV_X1 u0_u0_u0_U23 (.ZN( u0_u0_u0_n14 ) , .A( u0_u0_u0_n39 ) );
  AOI22_X1 u0_u0_u0_U24 (.A1( u0_u0_u0_n15 ) , .B1( u0_u0_u0_n57 ) , .ZN( u0_u0_u0_n64 ) , .A2( u0_u0_u0_n65 ) , .B2( u0_u0_u0_n66 ) );
  NAND2_X1 u0_u0_u0_U25 (.ZN( u0_u0_u0_n46 ) , .A1( u0_u0_u0_n75 ) , .A2( u0_u0_u0_n80 ) );
  INV_X1 u0_u0_u0_U26 (.ZN( u0_u0_u0_n17 ) , .A( u0_u0_u0_n57 ) );
  AOI21_X1 u0_u0_u0_U27 (.A( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n34 ) , .B1( u0_u0_u0_n68 ) , .ZN( u0_u0_u0_n71 ) );
  AOI21_X1 u0_u0_u0_U28 (.A( u0_u0_u0_n37 ) , .B2( u0_u0_u0_n46 ) , .B1( u0_u0_u0_n48 ) , .ZN( u0_u0_u0_n79 ) );
  AOI21_X1 u0_u0_u0_U29 (.A( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n33 ) , .ZN( u0_u0_u0_n59 ) , .B1( u0_u0_u0_n9 ) );
  INV_X1 u0_u0_u0_U3 (.A( u0_u0_u0_n62 ) , .ZN( u0_u0_u0_n9 ) );
  NOR2_X1 u0_u0_u0_U30 (.ZN( u0_u0_u0_n32 ) , .A1( u0_u0_u0_n55 ) , .A2( u0_u0_u0_n8 ) );
  OAI221_X1 u0_u0_u0_U31 (.C2( u0_u0_u0_n28 ) , .A( u0_u0_u0_n3 ) , .B2( u0_u0_u0_n34 ) , .B1( u0_u0_u0_n37 ) , .ZN( u0_u0_u0_n55 ) , .C1( u0_u0_u0_n63 ) );
  AOI211_X1 u0_u0_u0_U32 (.ZN( u0_u0_u0_n56 ) , .C1( u0_u0_u0_n57 ) , .C2( u0_u0_u0_n58 ) , .A( u0_u0_u0_n59 ) , .B( u0_u0_u0_n60 ) );
  NAND2_X1 u0_u0_u0_U33 (.ZN( u0_u0_u0_n47 ) , .A1( u0_u0_u0_n73 ) , .A2( u0_u0_u0_n80 ) );
  NAND2_X1 u0_u0_u0_U34 (.ZN( u0_u0_u0_n36 ) , .A1( u0_u0_u0_n74 ) , .A2( u0_u0_u0_n75 ) );
  NAND2_X1 u0_u0_u0_U35 (.ZN( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n80 ) , .A1( u0_u0_u0_n82 ) );
  NAND2_X1 u0_u0_u0_U36 (.ZN( u0_u0_u0_n44 ) , .A2( u0_u0_u0_n75 ) , .A1( u0_u0_u0_n83 ) );
  NAND2_X1 u0_u0_u0_U37 (.ZN( u0_u0_u0_n25 ) , .A2( u0_u0_u0_n73 ) , .A1( u0_u0_u0_n74 ) );
  INV_X1 u0_u0_u0_U38 (.ZN( u0_u0_u0_n15 ) , .A( u0_u0_u0_n37 ) );
  NAND2_X1 u0_u0_u0_U39 (.ZN( u0_u0_u0_n26 ) , .A1( u0_u0_u0_n72 ) , .A2( u0_u0_u0_n73 ) );
  AOI21_X1 u0_u0_u0_U4 (.A( u0_u0_u0_n14 ) , .B2( u0_u0_u0_n46 ) , .ZN( u0_u0_u0_n60 ) , .B1( u0_u0_u0_n61 ) );
  NAND2_X1 u0_u0_u0_U40 (.ZN( u0_u0_u0_n61 ) , .A2( u0_u0_u0_n73 ) , .A1( u0_u0_u0_n83 ) );
  INV_X1 u0_u0_u0_U41 (.ZN( u0_u0_u0_n3 ) , .A( u0_u0_u0_n87 ) );
  OAI222_X1 u0_u0_u0_U42 (.C2( u0_u0_u0_n14 ) , .A2( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n31 ) , .B2( u0_u0_u0_n47 ) , .A1( u0_u0_u0_n50 ) , .C1( u0_u0_u0_n67 ) , .ZN( u0_u0_u0_n87 ) );
  NAND2_X1 u0_u0_u0_U43 (.ZN( u0_u0_u0_n54 ) , .A2( u0_u0_u0_n74 ) , .A1( u0_u0_u0_n82 ) );
  NAND2_X1 u0_u0_u0_U44 (.ZN( u0_u0_u0_n63 ) , .A1( u0_u0_u0_n82 ) , .A2( u0_u0_u0_n83 ) );
  OR3_X1 u0_u0_u0_U45 (.ZN( u0_u0_u0_n20 ) , .A1( u0_u0_u0_n21 ) , .A2( u0_u0_u0_n22 ) , .A3( u0_u0_u0_n23 ) );
  AOI21_X1 u0_u0_u0_U46 (.A( u0_u0_u0_n17 ) , .ZN( u0_u0_u0_n23 ) , .B1( u0_u0_u0_n24 ) , .B2( u0_u0_u0_n25 ) );
  AOI21_X1 u0_u0_u0_U47 (.ZN( u0_u0_u0_n21 ) , .B1( u0_u0_u0_n29 ) , .B2( u0_u0_u0_n30 ) , .A( u0_u0_u0_n31 ) );
  AOI21_X1 u0_u0_u0_U48 (.ZN( u0_u0_u0_n22 ) , .B1( u0_u0_u0_n26 ) , .B2( u0_u0_u0_n27 ) , .A( u0_u0_u0_n28 ) );
  INV_X1 u0_u0_u0_U49 (.ZN( u0_u0_u0_n4 ) , .A( u0_u0_u0_n76 ) );
  AOI21_X1 u0_u0_u0_U5 (.A( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n24 ) , .ZN( u0_u0_u0_n41 ) , .B2( u0_u0_u0_n44 ) );
  OAI211_X1 u0_u0_u0_U50 (.C1( u0_u0_u0_n14 ) , .C2( u0_u0_u0_n35 ) , .A( u0_u0_u0_n6 ) , .ZN( u0_u0_u0_n76 ) , .B( u0_u0_u0_n77 ) );
  INV_X1 u0_u0_u0_U51 (.ZN( u0_u0_u0_n6 ) , .A( u0_u0_u0_n84 ) );
  AOI211_X1 u0_u0_u0_U52 (.A( u0_u0_u0_n52 ) , .C1( u0_u0_u0_n57 ) , .ZN( u0_u0_u0_n77 ) , .C2( u0_u0_u0_n78 ) , .B( u0_u0_u0_n79 ) );
  NOR2_X1 u0_u0_u0_U53 (.A2( u0_u0_X_4 ) , .A1( u0_u0_X_5 ) , .ZN( u0_u0_u0_n57 ) );
  NOR2_X1 u0_u0_u0_U54 (.A2( u0_u0_X_2 ) , .A1( u0_u0_u0_n11 ) , .ZN( u0_u0_u0_n72 ) );
  NOR2_X1 u0_u0_u0_U55 (.A2( u0_u0_X_1 ) , .A1( u0_u0_X_2 ) , .ZN( u0_u0_u0_n83 ) );
  NOR2_X1 u0_u0_u0_U56 (.A2( u0_u0_X_1 ) , .A1( u0_u0_u0_n12 ) , .ZN( u0_u0_u0_n74 ) );
  NAND2_X1 u0_u0_u0_U57 (.A2( u0_u0_X_4 ) , .A1( u0_u0_X_5 ) , .ZN( u0_u0_u0_n31 ) );
  NOR2_X1 u0_u0_u0_U58 (.A2( u0_u0_X_5 ) , .A1( u0_u0_u0_n16 ) , .ZN( u0_u0_u0_n39 ) );
  NAND2_X1 u0_u0_u0_U59 (.A1( u0_u0_X_5 ) , .A2( u0_u0_u0_n16 ) , .ZN( u0_u0_u0_n37 ) );
  NOR2_X1 u0_u0_u0_U6 (.A2( u0_u0_u0_n17 ) , .ZN( u0_u0_u0_n52 ) , .A1( u0_u0_u0_n67 ) );
  AND2_X1 u0_u0_u0_U60 (.A2( u0_u0_X_3 ) , .A1( u0_u0_X_6 ) , .ZN( u0_u0_u0_n73 ) );
  AND2_X1 u0_u0_u0_U61 (.A1( u0_u0_X_6 ) , .A2( u0_u0_u0_n13 ) , .ZN( u0_u0_u0_n82 ) );
  INV_X1 u0_u0_u0_U62 (.A( u0_u0_X_4 ) , .ZN( u0_u0_u0_n16 ) );
  INV_X1 u0_u0_u0_U63 (.A( u0_u0_X_2 ) , .ZN( u0_u0_u0_n12 ) );
  INV_X1 u0_u0_u0_U64 (.A( u0_u0_X_3 ) , .ZN( u0_u0_u0_n13 ) );
  AOI211_X1 u0_u0_u0_U65 (.C1( u0_u0_u0_n15 ) , .C2( u0_u0_u0_n62 ) , .ZN( u0_u0_u0_n69 ) , .A( u0_u0_u0_n70 ) , .B( u0_u0_u0_n71 ) );
  INV_X1 u0_u0_u0_U66 (.ZN( u0_u0_u0_n1 ) , .A( u0_u0_u0_n86 ) );
  OR4_X1 u0_u0_u0_U67 (.ZN( u0_out0_17 ) , .A3( u0_u0_u0_n5 ) , .A1( u0_u0_u0_n51 ) , .A2( u0_u0_u0_n52 ) , .A4( u0_u0_u0_n53 ) );
  AOI21_X1 u0_u0_u0_U68 (.A( u0_u0_u0_n14 ) , .B1( u0_u0_u0_n47 ) , .ZN( u0_u0_u0_n51 ) , .B2( u0_u0_u0_n68 ) );
  INV_X1 u0_u0_u0_U69 (.ZN( u0_u0_u0_n5 ) , .A( u0_u0_u0_n64 ) );
  OAI21_X1 u0_u0_u0_U7 (.B2( u0_u0_u0_n17 ) , .B1( u0_u0_u0_n25 ) , .A( u0_u0_u0_n3 ) , .ZN( u0_u0_u0_n86 ) );
  OR4_X1 u0_u0_u0_U70 (.ZN( u0_out0_31 ) , .A1( u0_u0_u0_n18 ) , .A2( u0_u0_u0_n19 ) , .A3( u0_u0_u0_n2 ) , .A4( u0_u0_u0_n20 ) );
  AOI21_X1 u0_u0_u0_U71 (.ZN( u0_u0_u0_n18 ) , .B1( u0_u0_u0_n35 ) , .B2( u0_u0_u0_n36 ) , .A( u0_u0_u0_n37 ) );
  AOI21_X1 u0_u0_u0_U72 (.A( u0_u0_u0_n14 ) , .ZN( u0_u0_u0_n19 ) , .B1( u0_u0_u0_n33 ) , .B2( u0_u0_u0_n34 ) );
  INV_X1 u0_u0_u0_U73 (.A( u0_u0_u0_n49 ) , .ZN( u0_u0_u0_n7 ) );
  AOI211_X1 u0_u0_u0_U74 (.ZN( u0_u0_u0_n38 ) , .C1( u0_u0_u0_n39 ) , .C2( u0_u0_u0_n40 ) , .A( u0_u0_u0_n41 ) , .B( u0_u0_u0_n42 ) );
  NOR2_X1 u0_u0_u0_U75 (.A2( u0_u0_u0_n11 ) , .A1( u0_u0_u0_n12 ) , .ZN( u0_u0_u0_n80 ) );
  OAI221_X1 u0_u0_u0_U76 (.C2( u0_u0_u0_n28 ) , .B1( u0_u0_u0_n31 ) , .A( u0_u0_u0_n32 ) , .B2( u0_u0_u0_n48 ) , .ZN( u0_u0_u0_n53 ) , .C1( u0_u0_u0_n54 ) );
  INV_X1 u0_u0_u0_U77 (.A( u0_u0_X_1 ) , .ZN( u0_u0_u0_n11 ) );
  AOI21_X1 u0_u0_u0_U78 (.A( u0_u0_u0_n31 ) , .ZN( u0_u0_u0_n42 ) , .B1( u0_u0_u0_n43 ) , .B2( u0_u0_u0_n9 ) );
  OAI22_X1 u0_u0_u0_U79 (.B2( u0_u0_u0_n14 ) , .A1( u0_u0_u0_n28 ) , .B1( u0_u0_u0_n29 ) , .A2( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n70 ) );
  AND2_X1 u0_u0_u0_U8 (.ZN( u0_u0_u0_n29 ) , .A2( u0_u0_u0_n54 ) , .A1( u0_u0_u0_n61 ) );
  NAND2_X1 u0_u0_u0_U80 (.A1( u0_u0_u0_n30 ) , .A2( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n65 ) );
  INV_X1 u0_u0_u0_U81 (.A( u0_u0_u0_n56 ) , .ZN( u0_u0_u0_n8 ) );
  NAND2_X1 u0_u0_u0_U82 (.ZN( u0_u0_u0_n35 ) , .A2( u0_u0_u0_n72 ) , .A1( u0_u0_u0_n81 ) );
  NAND2_X1 u0_u0_u0_U83 (.ZN( u0_u0_u0_n45 ) , .A1( u0_u0_u0_n74 ) , .A2( u0_u0_u0_n81 ) );
  NAND2_X1 u0_u0_u0_U84 (.ZN( u0_u0_u0_n67 ) , .A2( u0_u0_u0_n81 ) , .A1( u0_u0_u0_n83 ) );
  NAND2_X1 u0_u0_u0_U85 (.ZN( u0_u0_u0_n33 ) , .A2( u0_u0_u0_n80 ) , .A1( u0_u0_u0_n81 ) );
  NOR2_X1 u0_u0_u0_U86 (.A2( u0_u0_X_6 ) , .A1( u0_u0_u0_n13 ) , .ZN( u0_u0_u0_n75 ) );
  NOR2_X1 u0_u0_u0_U87 (.A2( u0_u0_X_3 ) , .A1( u0_u0_X_6 ) , .ZN( u0_u0_u0_n81 ) );
  NAND3_X1 u0_u0_u0_U88 (.ZN( u0_out0_23 ) , .A3( u0_u0_u0_n38 ) , .A2( u0_u0_u0_n4 ) , .A1( u0_u0_u0_n7 ) );
  NAND3_X1 u0_u0_u0_U89 (.A1( u0_u0_u0_n25 ) , .ZN( u0_u0_u0_n40 ) , .A2( u0_u0_u0_n47 ) , .A3( u0_u0_u0_n48 ) );
  AND2_X1 u0_u0_u0_U9 (.A2( u0_u0_u0_n25 ) , .ZN( u0_u0_u0_n34 ) , .A1( u0_u0_u0_n44 ) );
  NAND3_X1 u0_u0_u0_U90 (.A1( u0_u0_u0_n27 ) , .A2( u0_u0_u0_n36 ) , .A3( u0_u0_u0_n43 ) , .ZN( u0_u0_u0_n58 ) );
  NAND3_X1 u0_u0_u0_U91 (.A1( u0_u0_u0_n26 ) , .A3( u0_u0_u0_n35 ) , .A2( u0_u0_u0_n61 ) , .ZN( u0_u0_u0_n66 ) );
  NAND3_X1 u0_u0_u0_U92 (.ZN( u0_out0_9 ) , .A1( u0_u0_u0_n1 ) , .A2( u0_u0_u0_n4 ) , .A3( u0_u0_u0_n69 ) );
  NAND3_X1 u0_u0_u0_U93 (.A3( u0_u0_u0_n29 ) , .A1( u0_u0_u0_n43 ) , .A2( u0_u0_u0_n47 ) , .ZN( u0_u0_u0_n78 ) );
  AOI21_X1 u0_u0_u1_U10 (.A( u0_u0_u1_n15 ) , .ZN( u0_u0_u1_n32 ) , .B1( u0_u0_u1_n33 ) , .B2( u0_u0_u1_n34 ) );
  NAND3_X1 u0_u0_u1_U100 (.A2( u0_u0_u1_n34 ) , .A3( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n69 ) , .ZN( u0_u0_u1_n76 ) );
  NAND2_X1 u0_u0_u1_U11 (.A1( u0_u0_u1_n34 ) , .A2( u0_u0_u1_n39 ) , .ZN( u0_u0_u1_n49 ) );
  NAND2_X1 u0_u0_u1_U12 (.A2( u0_u0_u1_n36 ) , .ZN( u0_u0_u1_n42 ) , .A1( u0_u0_u1_n58 ) );
  AOI22_X1 u0_u0_u1_U13 (.B1( u0_u0_u1_n16 ) , .A1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n46 ) , .A2( u0_u0_u1_n52 ) , .B2( u0_u0_u1_n53 ) );
  INV_X1 u0_u0_u1_U14 (.A( u0_u0_u1_n42 ) , .ZN( u0_u0_u1_n8 ) );
  INV_X1 u0_u0_u1_U15 (.ZN( u0_u0_u1_n15 ) , .A( u0_u0_u1_n50 ) );
  OR4_X1 u0_u0_u1_U16 (.A2( u0_u0_u1_n5 ) , .A1( u0_u0_u1_n72 ) , .ZN( u0_u0_u1_n81 ) , .A3( u0_u0_u1_n82 ) , .A4( u0_u0_u1_n83 ) );
  AOI21_X1 u0_u0_u1_U17 (.B2( u0_u0_u1_n33 ) , .B1( u0_u0_u1_n35 ) , .A( u0_u0_u1_n77 ) , .ZN( u0_u0_u1_n83 ) );
  AOI21_X1 u0_u0_u1_U18 (.A( u0_u0_u1_n15 ) , .B2( u0_u0_u1_n40 ) , .B1( u0_u0_u1_n55 ) , .ZN( u0_u0_u1_n82 ) );
  INV_X1 u0_u0_u1_U19 (.ZN( u0_u0_u1_n5 ) , .A( u0_u0_u1_n88 ) );
  INV_X1 u0_u0_u1_U20 (.ZN( u0_u0_u1_n18 ) , .A( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U21 (.A2( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n36 ) , .ZN( u0_u0_u1_n48 ) );
  AND2_X1 u0_u0_u1_U22 (.A2( u0_u0_u1_n28 ) , .ZN( u0_u0_u1_n55 ) , .A1( u0_u0_u1_n66 ) );
  NAND2_X1 u0_u0_u1_U23 (.ZN( u0_u0_u1_n41 ) , .A1( u0_u0_u1_n73 ) , .A2( u0_u0_u1_n74 ) );
  NAND2_X1 u0_u0_u1_U24 (.ZN( u0_u0_u1_n30 ) , .A1( u0_u0_u1_n54 ) , .A2( u0_u0_u1_n56 ) );
  NAND2_X1 u0_u0_u1_U25 (.ZN( u0_u0_u1_n57 ) , .A1( u0_u0_u1_n69 ) , .A2( u0_u0_u1_n74 ) );
  INV_X1 u0_u0_u1_U26 (.ZN( u0_u0_u1_n11 ) , .A( u0_u0_u1_n35 ) );
  INV_X1 u0_u0_u1_U27 (.A( u0_u0_u1_n38 ) , .ZN( u0_u0_u1_n6 ) );
  AND2_X1 u0_u0_u1_U28 (.ZN( u0_u0_u1_n40 ) , .A2( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n60 ) );
  INV_X1 u0_u0_u1_U29 (.A( u0_u0_u1_n58 ) , .ZN( u0_u0_u1_n9 ) );
  INV_X1 u0_u0_u1_U3 (.A( u0_u0_u1_n30 ) , .ZN( u0_u0_u1_n7 ) );
  AOI221_X1 u0_u0_u1_U30 (.A( u0_u0_u1_n1 ) , .C1( u0_u0_u1_n11 ) , .C2( u0_u0_u1_n14 ) , .B2( u0_u0_u1_n17 ) , .ZN( u0_u0_u1_n22 ) , .B1( u0_u0_u1_n49 ) );
  INV_X1 u0_u0_u1_U31 (.ZN( u0_u0_u1_n1 ) , .A( u0_u0_u1_n92 ) );
  AOI211_X1 u0_u0_u1_U32 (.C2( u0_u0_u1_n50 ) , .C1( u0_u0_u1_n57 ) , .A( u0_u0_u1_n71 ) , .ZN( u0_u0_u1_n92 ) , .B( u0_u0_u1_n93 ) );
  AOI21_X1 u0_u0_u1_U33 (.A( u0_u0_u1_n37 ) , .B1( u0_u0_u1_n54 ) , .B2( u0_u0_u1_n68 ) , .ZN( u0_u0_u1_n93 ) );
  OAI221_X1 u0_u0_u1_U34 (.C1( u0_u0_u1_n15 ) , .B1( u0_u0_u1_n2 ) , .B2( u0_u0_u1_n37 ) , .ZN( u0_u0_u1_n51 ) , .C2( u0_u0_u1_n60 ) , .A( u0_u0_u1_n70 ) );
  INV_X1 u0_u0_u1_U35 (.ZN( u0_u0_u1_n2 ) , .A( u0_u0_u1_n41 ) );
  AOI211_X1 u0_u0_u1_U36 (.C1( u0_u0_u1_n30 ) , .C2( u0_u0_u1_n43 ) , .ZN( u0_u0_u1_n70 ) , .A( u0_u0_u1_n71 ) , .B( u0_u0_u1_n72 ) );
  NOR2_X1 u0_u0_u1_U37 (.A2( u0_u0_u1_n13 ) , .A1( u0_u0_u1_n21 ) , .ZN( u0_u0_u1_n91 ) );
  AOI211_X1 u0_u0_u1_U38 (.C1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n24 ) , .C2( u0_u0_u1_n25 ) , .A( u0_u0_u1_n26 ) , .B( u0_u0_u1_n27 ) );
  AOI21_X1 u0_u0_u1_U39 (.ZN( u0_u0_u1_n27 ) , .B2( u0_u0_u1_n28 ) , .A( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n7 ) );
  AOI221_X1 u0_u0_u1_U4 (.B1( u0_u0_u1_n14 ) , .ZN( u0_u0_u1_n47 ) , .B2( u0_u0_u1_n48 ) , .C1( u0_u0_u1_n49 ) , .C2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n51 ) );
  OR2_X1 u0_u0_u1_U40 (.ZN( u0_u0_u1_n26 ) , .A1( u0_u0_u1_n31 ) , .A2( u0_u0_u1_n32 ) );
  NAND2_X1 u0_u0_u1_U41 (.A2( u0_u0_u1_n29 ) , .ZN( u0_u0_u1_n43 ) , .A1( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U42 (.A1( u0_u0_u1_n37 ) , .ZN( u0_u0_u1_n50 ) , .A2( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U43 (.ZN( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n90 ) );
  NOR2_X1 u0_u0_u1_U44 (.A2( u0_u0_u1_n29 ) , .A1( u0_u0_u1_n68 ) , .ZN( u0_u0_u1_n72 ) );
  AOI21_X1 u0_u0_u1_U45 (.B1( u0_u0_u1_n39 ) , .ZN( u0_u0_u1_n59 ) , .B2( u0_u0_u1_n60 ) , .A( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U46 (.A2( u0_u0_u1_n19 ) , .A1( u0_u0_u1_n20 ) , .ZN( u0_u0_u1_n77 ) );
  NAND2_X1 u0_u0_u1_U47 (.ZN( u0_u0_u1_n60 ) , .A1( u0_u0_u1_n91 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U48 (.ZN( u0_u0_u1_n35 ) , .A1( u0_u0_u1_n87 ) , .A2( u0_u0_u1_n90 ) );
  NAND2_X1 u0_u0_u1_U49 (.ZN( u0_u0_u1_n54 ) , .A2( u0_u0_u1_n89 ) , .A1( u0_u0_u1_n90 ) );
  AOI211_X1 u0_u0_u1_U5 (.C1( u0_u0_u1_n42 ) , .B( u0_u0_u1_n44 ) , .C2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n51 ) , .ZN( u0_u0_u1_n65 ) );
  AOI21_X1 u0_u0_u1_U50 (.ZN( u0_u0_u1_n31 ) , .B1( u0_u0_u1_n35 ) , .B2( u0_u0_u1_n36 ) , .A( u0_u0_u1_n37 ) );
  INV_X1 u0_u0_u1_U51 (.ZN( u0_u0_u1_n14 ) , .A( u0_u0_u1_n29 ) );
  NAND2_X1 u0_u0_u1_U52 (.ZN( u0_u0_u1_n73 ) , .A1( u0_u0_u1_n89 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U53 (.ZN( u0_u0_u1_n58 ) , .A1( u0_u0_u1_n87 ) , .A2( u0_u0_u1_n94 ) );
  NAND2_X1 u0_u0_u1_U54 (.ZN( u0_u0_u1_n68 ) , .A2( u0_u0_u1_n85 ) , .A1( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U55 (.ZN( u0_u0_u1_n36 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U56 (.ZN( u0_u0_u1_n56 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n85 ) );
  NAND2_X1 u0_u0_u1_U57 (.ZN( u0_u0_u1_n39 ) , .A1( u0_u0_u1_n90 ) , .A2( u0_u0_u1_n91 ) );
  NAND2_X1 u0_u0_u1_U58 (.ZN( u0_u0_u1_n34 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n94 ) );
  OAI21_X1 u0_u0_u1_U59 (.A( u0_u0_u1_n22 ) , .B2( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n60 ) , .ZN( u0_u0_u1_n80 ) );
  AOI22_X1 u0_u0_u1_U6 (.B1( u0_u0_u1_n16 ) , .A1( u0_u0_u1_n18 ) , .ZN( u0_u0_u1_n64 ) , .A2( u0_u0_u1_n75 ) , .B2( u0_u0_u1_n76 ) );
  NAND2_X1 u0_u0_u1_U60 (.ZN( u0_u0_u1_n69 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n89 ) );
  NAND2_X1 u0_u0_u1_U61 (.ZN( u0_u0_u1_n74 ) , .A2( u0_u0_u1_n85 ) , .A1( u0_u0_u1_n87 ) );
  NAND2_X1 u0_u0_u1_U62 (.ZN( u0_u0_u1_n38 ) , .A1( u0_u0_u1_n85 ) , .A2( u0_u0_u1_n89 ) );
  NAND2_X1 u0_u0_u1_U63 (.ZN( u0_u0_u1_n28 ) , .A1( u0_u0_u1_n84 ) , .A2( u0_u0_u1_n86 ) );
  INV_X1 u0_u0_u1_U64 (.ZN( u0_u0_u1_n16 ) , .A( u0_u0_u1_n37 ) );
  INV_X1 u0_u0_u1_U65 (.ZN( u0_u0_u1_n17 ) , .A( u0_u0_u1_n61 ) );
  NAND2_X1 u0_u0_u1_U66 (.ZN( u0_u0_u1_n66 ) , .A1( u0_u0_u1_n86 ) , .A2( u0_u0_u1_n87 ) );
  OAI21_X1 u0_u0_u1_U67 (.B1( u0_u0_u1_n29 ) , .A( u0_u0_u1_n4 ) , .ZN( u0_u0_u1_n44 ) , .B2( u0_u0_u1_n66 ) );
  INV_X1 u0_u0_u1_U68 (.ZN( u0_u0_u1_n4 ) , .A( u0_u0_u1_n67 ) );
  AOI21_X1 u0_u0_u1_U69 (.A( u0_u0_u1_n61 ) , .ZN( u0_u0_u1_n67 ) , .B1( u0_u0_u1_n68 ) , .B2( u0_u0_u1_n69 ) );
  NAND2_X1 u0_u0_u1_U7 (.A2( u0_u0_u1_n33 ) , .A1( u0_u0_u1_n55 ) , .ZN( u0_u0_u1_n75 ) );
  NOR2_X1 u0_u0_u1_U70 (.A2( u0_u0_X_7 ) , .A1( u0_u0_X_8 ) , .ZN( u0_u0_u1_n94 ) );
  NOR2_X1 u0_u0_u1_U71 (.A1( u0_u0_X_12 ) , .A2( u0_u0_X_9 ) , .ZN( u0_u0_u1_n89 ) );
  NOR2_X1 u0_u0_u1_U72 (.A2( u0_u0_X_8 ) , .A1( u0_u0_u1_n12 ) , .ZN( u0_u0_u1_n90 ) );
  NOR2_X1 u0_u0_u1_U73 (.A2( u0_u0_X_12 ) , .A1( u0_u0_u1_n13 ) , .ZN( u0_u0_u1_n87 ) );
  NOR2_X1 u0_u0_u1_U74 (.A2( u0_u0_X_9 ) , .A1( u0_u0_u1_n21 ) , .ZN( u0_u0_u1_n84 ) );
  NAND2_X1 u0_u0_u1_U75 (.A1( u0_u0_X_10 ) , .A2( u0_u0_u1_n20 ) , .ZN( u0_u0_u1_n29 ) );
  NAND2_X1 u0_u0_u1_U76 (.A2( u0_u0_X_10 ) , .A1( u0_u0_X_11 ) , .ZN( u0_u0_u1_n37 ) );
  NAND2_X1 u0_u0_u1_U77 (.A1( u0_u0_X_11 ) , .A2( u0_u0_u1_n19 ) , .ZN( u0_u0_u1_n61 ) );
  AND2_X1 u0_u0_u1_U78 (.A2( u0_u0_X_7 ) , .A1( u0_u0_X_8 ) , .ZN( u0_u0_u1_n85 ) );
  AND2_X1 u0_u0_u1_U79 (.A1( u0_u0_X_8 ) , .A2( u0_u0_u1_n12 ) , .ZN( u0_u0_u1_n86 ) );
  NOR2_X1 u0_u0_u1_U8 (.ZN( u0_u0_u1_n71 ) , .A2( u0_u0_u1_n73 ) , .A1( u0_u0_u1_n77 ) );
  INV_X1 u0_u0_u1_U80 (.A( u0_u0_X_10 ) , .ZN( u0_u0_u1_n19 ) );
  INV_X1 u0_u0_u1_U81 (.A( u0_u0_X_9 ) , .ZN( u0_u0_u1_n13 ) );
  INV_X1 u0_u0_u1_U82 (.A( u0_u0_X_11 ) , .ZN( u0_u0_u1_n20 ) );
  INV_X1 u0_u0_u1_U83 (.A( u0_u0_X_12 ) , .ZN( u0_u0_u1_n21 ) );
  INV_X1 u0_u0_u1_U84 (.A( u0_u0_X_7 ) , .ZN( u0_u0_u1_n12 ) );
  NAND4_X1 u0_u0_u1_U85 (.ZN( u0_out0_18 ) , .A1( u0_u0_u1_n22 ) , .A3( u0_u0_u1_n23 ) , .A4( u0_u0_u1_n24 ) , .A2( u0_u0_u1_n3 ) );
  AOI22_X1 u0_u0_u1_U86 (.A1( u0_u0_u1_n17 ) , .ZN( u0_u0_u1_n23 ) , .A2( u0_u0_u1_n41 ) , .B1( u0_u0_u1_n42 ) , .B2( u0_u0_u1_n43 ) );
  INV_X1 u0_u0_u1_U87 (.ZN( u0_u0_u1_n3 ) , .A( u0_u0_u1_n44 ) );
  NAND4_X1 u0_u0_u1_U88 (.ZN( u0_out0_2 ) , .A1( u0_u0_u1_n10 ) , .A2( u0_u0_u1_n45 ) , .A3( u0_u0_u1_n46 ) , .A4( u0_u0_u1_n47 ) );
  OAI21_X1 u0_u0_u1_U89 (.A( u0_u0_u1_n43 ) , .ZN( u0_u0_u1_n45 ) , .B2( u0_u0_u1_n57 ) , .B1( u0_u0_u1_n9 ) );
  OAI21_X1 u0_u0_u1_U9 (.A( u0_u0_u1_n43 ) , .B1( u0_u0_u1_n48 ) , .B2( u0_u0_u1_n6 ) , .ZN( u0_u0_u1_n88 ) );
  INV_X1 u0_u0_u1_U90 (.ZN( u0_u0_u1_n10 ) , .A( u0_u0_u1_n59 ) );
  NAND4_X1 u0_u0_u1_U91 (.ZN( u0_out0_28 ) , .A1( u0_u0_u1_n62 ) , .A2( u0_u0_u1_n63 ) , .A3( u0_u0_u1_n64 ) , .A4( u0_u0_u1_n65 ) );
  OAI21_X1 u0_u0_u1_U92 (.B1( u0_u0_u1_n14 ) , .B2( u0_u0_u1_n50 ) , .A( u0_u0_u1_n6 ) , .ZN( u0_u0_u1_n62 ) );
  OAI21_X1 u0_u0_u1_U93 (.B1( u0_u0_u1_n11 ) , .A( u0_u0_u1_n43 ) , .B2( u0_u0_u1_n49 ) , .ZN( u0_u0_u1_n63 ) );
  OR4_X1 u0_u0_u1_U94 (.ZN( u0_out0_13 ) , .A1( u0_u0_u1_n78 ) , .A2( u0_u0_u1_n79 ) , .A3( u0_u0_u1_n80 ) , .A4( u0_u0_u1_n81 ) );
  AOI21_X1 u0_u0_u1_U95 (.B1( u0_u0_u1_n54 ) , .B2( u0_u0_u1_n58 ) , .A( u0_u0_u1_n61 ) , .ZN( u0_u0_u1_n78 ) );
  AOI21_X1 u0_u0_u1_U96 (.B2( u0_u0_u1_n29 ) , .B1( u0_u0_u1_n37 ) , .A( u0_u0_u1_n73 ) , .ZN( u0_u0_u1_n79 ) );
  NAND3_X1 u0_u0_u1_U97 (.ZN( u0_u0_u1_n25 ) , .A1( u0_u0_u1_n38 ) , .A2( u0_u0_u1_n39 ) , .A3( u0_u0_u1_n40 ) );
  NAND3_X1 u0_u0_u1_U98 (.A1( u0_u0_u1_n38 ) , .ZN( u0_u0_u1_n53 ) , .A2( u0_u0_u1_n54 ) , .A3( u0_u0_u1_n55 ) );
  NAND3_X1 u0_u0_u1_U99 (.A2( u0_u0_u1_n35 ) , .ZN( u0_u0_u1_n52 ) , .A1( u0_u0_u1_n56 ) , .A3( u0_u0_u1_n8 ) );
  OAI22_X1 u0_u0_u2_U10 (.B2( u0_u0_u2_n21 ) , .ZN( u0_u0_u2_n29 ) , .A1( u0_u0_u2_n36 ) , .A2( u0_u0_u2_n37 ) , .B1( u0_u0_u2_n38 ) );
  NAND3_X1 u0_u0_u2_U100 (.A3( u0_u0_u2_n51 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n89 ) , .ZN( u0_u0_u2_n91 ) );
  NOR3_X1 u0_u0_u2_U11 (.A2( u0_u0_u2_n1 ) , .A3( u0_u0_u2_n14 ) , .ZN( u0_u0_u2_n38 ) , .A1( u0_u0_u2_n39 ) );
  AOI21_X1 u0_u0_u2_U12 (.A( u0_u0_u2_n18 ) , .B1( u0_u0_u2_n5 ) , .ZN( u0_u0_u2_n64 ) , .B2( u0_u0_u2_n66 ) );
  INV_X1 u0_u0_u2_U13 (.A( u0_u0_u2_n39 ) , .ZN( u0_u0_u2_n5 ) );
  AOI21_X1 u0_u0_u2_U14 (.A( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n34 ) , .B1( u0_u0_u2_n4 ) , .ZN( u0_u0_u2_n45 ) );
  AOI21_X1 u0_u0_u2_U15 (.A( u0_u0_u2_n18 ) , .B1( u0_u0_u2_n37 ) , .ZN( u0_u0_u2_n44 ) , .B2( u0_u0_u2_n46 ) );
  INV_X1 u0_u0_u2_U16 (.ZN( u0_u0_u2_n18 ) , .A( u0_u0_u2_n33 ) );
  INV_X1 u0_u0_u2_U17 (.ZN( u0_u0_u2_n1 ) , .A( u0_u0_u2_n69 ) );
  NAND2_X1 u0_u0_u2_U18 (.A1( u0_u0_u2_n37 ) , .ZN( u0_u0_u2_n39 ) , .A2( u0_u0_u2_n67 ) );
  INV_X1 u0_u0_u2_U19 (.ZN( u0_u0_u2_n19 ) , .A( u0_u0_u2_n36 ) );
  INV_X1 u0_u0_u2_U20 (.ZN( u0_u0_u2_n16 ) , .A( u0_u0_u2_n52 ) );
  NAND2_X1 u0_u0_u2_U21 (.ZN( u0_u0_u2_n32 ) , .A2( u0_u0_u2_n50 ) , .A1( u0_u0_u2_n57 ) );
  INV_X1 u0_u0_u2_U22 (.ZN( u0_u0_u2_n11 ) , .A( u0_u0_u2_n76 ) );
  INV_X1 u0_u0_u2_U23 (.ZN( u0_u0_u2_n14 ) , .A( u0_u0_u2_n50 ) );
  INV_X1 u0_u0_u2_U24 (.A( u0_u0_u2_n34 ) , .ZN( u0_u0_u2_n8 ) );
  INV_X1 u0_u0_u2_U25 (.ZN( u0_u0_u2_n12 ) , .A( u0_u0_u2_n70 ) );
  INV_X1 u0_u0_u2_U26 (.A( u0_u0_u2_n73 ) , .ZN( u0_u0_u2_n9 ) );
  INV_X1 u0_u0_u2_U27 (.ZN( u0_u0_u2_n10 ) , .A( u0_u0_u2_n58 ) );
  INV_X1 u0_u0_u2_U28 (.ZN( u0_u0_u2_n13 ) , .A( u0_u0_u2_n35 ) );
  NAND2_X1 u0_u0_u2_U29 (.ZN( u0_u0_u2_n71 ) , .A1( u0_u0_u2_n72 ) , .A2( u0_u0_u2_n73 ) );
  NOR2_X1 u0_u0_u2_U3 (.A2( u0_u0_u2_n12 ) , .ZN( u0_u0_u2_n68 ) , .A1( u0_u0_u2_n9 ) );
  INV_X1 u0_u0_u2_U30 (.A( u0_u0_u2_n57 ) , .ZN( u0_u0_u2_n7 ) );
  INV_X1 u0_u0_u2_U31 (.A( u0_u0_u2_n31 ) , .ZN( u0_u0_u2_n6 ) );
  OAI21_X1 u0_u0_u2_U32 (.B2( u0_u0_u2_n10 ) , .ZN( u0_u0_u2_n31 ) , .B1( u0_u0_u2_n32 ) , .A( u0_u0_u2_n33 ) );
  NOR2_X1 u0_u0_u2_U33 (.A2( u0_u0_u2_n20 ) , .A1( u0_u0_u2_n23 ) , .ZN( u0_u0_u2_n33 ) );
  NOR2_X1 u0_u0_u2_U34 (.A1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n52 ) , .A2( u0_u0_u2_n75 ) );
  NOR2_X1 u0_u0_u2_U35 (.A1( u0_u0_u2_n33 ) , .ZN( u0_u0_u2_n36 ) , .A2( u0_u0_u2_n51 ) );
  AOI211_X1 u0_u0_u2_U36 (.C2( u0_u0_u2_n10 ) , .C1( u0_u0_u2_n51 ) , .ZN( u0_u0_u2_n59 ) , .A( u0_u0_u2_n92 ) , .B( u0_u0_u2_n93 ) );
  OAI22_X1 u0_u0_u2_U37 (.B2( u0_u0_u2_n21 ) , .A1( u0_u0_u2_n37 ) , .A2( u0_u0_u2_n52 ) , .B1( u0_u0_u2_n56 ) , .ZN( u0_u0_u2_n92 ) );
  OAI221_X1 u0_u0_u2_U38 (.C2( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n18 ) , .A( u0_u0_u2_n40 ) , .C1( u0_u0_u2_n57 ) , .B1( u0_u0_u2_n76 ) , .ZN( u0_u0_u2_n93 ) );
  OAI221_X1 u0_u0_u2_U39 (.C1( u0_u0_u2_n21 ) , .ZN( u0_u0_u2_n26 ) , .B1( u0_u0_u2_n36 ) , .B2( u0_u0_u2_n46 ) , .C2( u0_u0_u2_n66 ) , .A( u0_u0_u2_n74 ) );
  INV_X1 u0_u0_u2_U4 (.ZN( u0_u0_u2_n4 ) , .A( u0_u0_u2_n55 ) );
  OAI21_X1 u0_u0_u2_U40 (.B2( u0_u0_u2_n11 ) , .B1( u0_u0_u2_n13 ) , .ZN( u0_u0_u2_n74 ) , .A( u0_u0_u2_n75 ) );
  OAI221_X1 u0_u0_u2_U41 (.C2( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n27 ) , .C1( u0_u0_u2_n4 ) , .B1( u0_u0_u2_n52 ) , .B2( u0_u0_u2_n53 ) , .A( u0_u0_u2_n54 ) );
  AND3_X1 u0_u0_u2_U42 (.ZN( u0_u0_u2_n53 ) , .A1( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n57 ) , .A3( u0_u0_u2_n58 ) );
  AOI22_X1 u0_u0_u2_U43 (.A2( u0_u0_u2_n1 ) , .A1( u0_u0_u2_n33 ) , .B1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n54 ) , .B2( u0_u0_u2_n9 ) );
  AOI21_X1 u0_u0_u2_U44 (.B2( u0_u0_u2_n1 ) , .B1( u0_u0_u2_n16 ) , .ZN( u0_u0_u2_n40 ) , .A( u0_u0_u2_n94 ) );
  AND3_X1 u0_u0_u2_U45 (.A3( u0_u0_u2_n33 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n89 ) , .ZN( u0_u0_u2_n94 ) );
  OAI21_X1 u0_u0_u2_U46 (.B1( u0_u0_u2_n36 ) , .ZN( u0_u0_u2_n43 ) , .B2( u0_u0_u2_n47 ) , .A( u0_u0_u2_n48 ) );
  OAI21_X1 u0_u0_u2_U47 (.B2( u0_u0_u2_n12 ) , .B1( u0_u0_u2_n13 ) , .ZN( u0_u0_u2_n48 ) , .A( u0_u0_u2_n49 ) );
  NOR3_X1 u0_u0_u2_U48 (.A2( u0_u0_u2_n11 ) , .A3( u0_u0_u2_n14 ) , .ZN( u0_u0_u2_n47 ) , .A1( u0_u0_u2_n8 ) );
  OAI21_X1 u0_u0_u2_U49 (.ZN( u0_u0_u2_n25 ) , .B1( u0_u0_u2_n36 ) , .B2( u0_u0_u2_n68 ) , .A( u0_u0_u2_n88 ) );
  NOR4_X1 u0_u0_u2_U5 (.ZN( u0_u0_u2_n61 ) , .A1( u0_u0_u2_n62 ) , .A2( u0_u0_u2_n63 ) , .A3( u0_u0_u2_n64 ) , .A4( u0_u0_u2_n65 ) );
  NAND2_X1 u0_u0_u2_U50 (.ZN( u0_u0_u2_n34 ) , .A1( u0_u0_u2_n82 ) , .A2( u0_u0_u2_n89 ) );
  NAND2_X1 u0_u0_u2_U51 (.ZN( u0_u0_u2_n46 ) , .A1( u0_u0_u2_n81 ) , .A2( u0_u0_u2_n84 ) );
  NAND2_X1 u0_u0_u2_U52 (.ZN( u0_u0_u2_n37 ) , .A2( u0_u0_u2_n83 ) , .A1( u0_u0_u2_n85 ) );
  NAND2_X1 u0_u0_u2_U53 (.ZN( u0_u0_u2_n57 ) , .A2( u0_u0_u2_n84 ) , .A1( u0_u0_u2_n89 ) );
  INV_X1 u0_u0_u2_U54 (.ZN( u0_u0_u2_n21 ) , .A( u0_u0_u2_n49 ) );
  INV_X1 u0_u0_u2_U55 (.ZN( u0_u0_u2_n22 ) , .A( u0_u0_u2_n51 ) );
  NAND2_X1 u0_u0_u2_U56 (.ZN( u0_u0_u2_n76 ) , .A2( u0_u0_u2_n83 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U57 (.ZN( u0_u0_u2_n58 ) , .A2( u0_u0_u2_n82 ) , .A1( u0_u0_u2_n83 ) );
  NAND2_X1 u0_u0_u2_U58 (.ZN( u0_u0_u2_n50 ) , .A2( u0_u0_u2_n82 ) , .A1( u0_u0_u2_n86 ) );
  NAND2_X1 u0_u0_u2_U59 (.ZN( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n84 ) , .A1( u0_u0_u2_n86 ) );
  AOI21_X1 u0_u0_u2_U6 (.B1( u0_u0_u2_n34 ) , .A( u0_u0_u2_n52 ) , .ZN( u0_u0_u2_n62 ) , .B2( u0_u0_u2_n70 ) );
  NAND2_X1 u0_u0_u2_U60 (.ZN( u0_u0_u2_n35 ) , .A2( u0_u0_u2_n86 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U61 (.ZN( u0_u0_u2_n70 ) , .A1( u0_u0_u2_n85 ) , .A2( u0_u0_u2_n86 ) );
  NAND2_X1 u0_u0_u2_U62 (.ZN( u0_u0_u2_n66 ) , .A1( u0_u0_u2_n81 ) , .A2( u0_u0_u2_n82 ) );
  NAND2_X1 u0_u0_u2_U63 (.ZN( u0_u0_u2_n67 ) , .A2( u0_u0_u2_n81 ) , .A1( u0_u0_u2_n85 ) );
  INV_X1 u0_u0_u2_U64 (.ZN( u0_u0_u2_n17 ) , .A( u0_u0_u2_n75 ) );
  NAND2_X1 u0_u0_u2_U65 (.ZN( u0_u0_u2_n73 ) , .A1( u0_u0_u2_n87 ) , .A2( u0_u0_u2_n89 ) );
  NAND2_X1 u0_u0_u2_U66 (.ZN( u0_u0_u2_n69 ) , .A2( u0_u0_u2_n81 ) , .A1( u0_u0_u2_n87 ) );
  NAND2_X1 u0_u0_u2_U67 (.ZN( u0_u0_u2_n72 ) , .A1( u0_u0_u2_n83 ) , .A2( u0_u0_u2_n84 ) );
  INV_X1 u0_u0_u2_U68 (.ZN( u0_u0_u2_n2 ) , .A( u0_u0_u2_n90 ) );
  OAI21_X1 u0_u0_u2_U69 (.B2( u0_u0_u2_n46 ) , .B1( u0_u0_u2_n52 ) , .ZN( u0_u0_u2_n90 ) , .A( u0_u0_u2_n91 ) );
  AOI21_X1 u0_u0_u2_U7 (.A( u0_u0_u2_n17 ) , .B2( u0_u0_u2_n46 ) , .B1( u0_u0_u2_n58 ) , .ZN( u0_u0_u2_n65 ) );
  NOR2_X1 u0_u0_u2_U70 (.A2( u0_u0_X_16 ) , .A1( u0_u0_u2_n23 ) , .ZN( u0_u0_u2_n49 ) );
  NOR2_X1 u0_u0_u2_U71 (.A2( u0_u0_X_13 ) , .A1( u0_u0_X_14 ) , .ZN( u0_u0_u2_n89 ) );
  NOR2_X1 u0_u0_u2_U72 (.A2( u0_u0_X_16 ) , .A1( u0_u0_X_17 ) , .ZN( u0_u0_u2_n51 ) );
  NOR2_X1 u0_u0_u2_U73 (.A2( u0_u0_X_15 ) , .A1( u0_u0_X_18 ) , .ZN( u0_u0_u2_n85 ) );
  NOR2_X1 u0_u0_u2_U74 (.A2( u0_u0_X_14 ) , .A1( u0_u0_u2_n15 ) , .ZN( u0_u0_u2_n86 ) );
  NOR2_X1 u0_u0_u2_U75 (.A2( u0_u0_X_15 ) , .A1( u0_u0_u2_n24 ) , .ZN( u0_u0_u2_n87 ) );
  NOR2_X1 u0_u0_u2_U76 (.A2( u0_u0_X_17 ) , .A1( u0_u0_u2_n20 ) , .ZN( u0_u0_u2_n75 ) );
  AND2_X1 u0_u0_u2_U77 (.A1( u0_u0_X_15 ) , .A2( u0_u0_u2_n24 ) , .ZN( u0_u0_u2_n84 ) );
  AND2_X1 u0_u0_u2_U78 (.A2( u0_u0_X_15 ) , .A1( u0_u0_X_18 ) , .ZN( u0_u0_u2_n82 ) );
  AND2_X1 u0_u0_u2_U79 (.A1( u0_u0_X_14 ) , .A2( u0_u0_u2_n15 ) , .ZN( u0_u0_u2_n83 ) );
  AOI21_X1 u0_u0_u2_U8 (.A( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n63 ) , .B1( u0_u0_u2_n68 ) , .B2( u0_u0_u2_n69 ) );
  AND2_X1 u0_u0_u2_U80 (.A1( u0_u0_X_13 ) , .A2( u0_u0_X_14 ) , .ZN( u0_u0_u2_n81 ) );
  INV_X1 u0_u0_u2_U81 (.A( u0_u0_X_16 ) , .ZN( u0_u0_u2_n20 ) );
  INV_X1 u0_u0_u2_U82 (.A( u0_u0_X_17 ) , .ZN( u0_u0_u2_n23 ) );
  INV_X1 u0_u0_u2_U83 (.A( u0_u0_X_13 ) , .ZN( u0_u0_u2_n15 ) );
  INV_X1 u0_u0_u2_U84 (.A( u0_u0_X_18 ) , .ZN( u0_u0_u2_n24 ) );
  NAND4_X1 u0_u0_u2_U85 (.ZN( u0_out0_30 ) , .A1( u0_u0_u2_n2 ) , .A2( u0_u0_u2_n40 ) , .A3( u0_u0_u2_n41 ) , .A4( u0_u0_u2_n42 ) );
  NOR3_X1 u0_u0_u2_U86 (.ZN( u0_u0_u2_n42 ) , .A1( u0_u0_u2_n43 ) , .A2( u0_u0_u2_n44 ) , .A3( u0_u0_u2_n45 ) );
  AOI21_X1 u0_u0_u2_U87 (.A( u0_u0_u2_n27 ) , .ZN( u0_u0_u2_n41 ) , .B2( u0_u0_u2_n51 ) , .B1( u0_u0_u2_n7 ) );
  NAND4_X1 u0_u0_u2_U88 (.ZN( u0_out0_24 ) , .A2( u0_u0_u2_n2 ) , .A1( u0_u0_u2_n59 ) , .A3( u0_u0_u2_n77 ) , .A4( u0_u0_u2_n78 ) );
  AOI221_X1 u0_u0_u2_U89 (.B2( u0_u0_u2_n16 ) , .C2( u0_u0_u2_n19 ) , .C1( u0_u0_u2_n55 ) , .ZN( u0_u0_u2_n78 ) , .B1( u0_u0_u2_n79 ) , .A( u0_u0_u2_n80 ) );
  OAI22_X1 u0_u0_u2_U9 (.A1( u0_u0_u2_n21 ) , .B1( u0_u0_u2_n22 ) , .B2( u0_u0_u2_n56 ) , .A2( u0_u0_u2_n76 ) , .ZN( u0_u0_u2_n80 ) );
  AOI21_X1 u0_u0_u2_U90 (.A( u0_u0_u2_n25 ) , .B2( u0_u0_u2_n33 ) , .ZN( u0_u0_u2_n77 ) , .B1( u0_u0_u2_n8 ) );
  NAND4_X1 u0_u0_u2_U91 (.ZN( u0_out0_16 ) , .A2( u0_u0_u2_n3 ) , .A1( u0_u0_u2_n59 ) , .A3( u0_u0_u2_n60 ) , .A4( u0_u0_u2_n61 ) );
  AOI22_X1 u0_u0_u2_U92 (.B2( u0_u0_u2_n19 ) , .B1( u0_u0_u2_n32 ) , .A1( u0_u0_u2_n49 ) , .ZN( u0_u0_u2_n60 ) , .A2( u0_u0_u2_n71 ) );
  INV_X1 u0_u0_u2_U93 (.A( u0_u0_u2_n26 ) , .ZN( u0_u0_u2_n3 ) );
  OR4_X1 u0_u0_u2_U94 (.ZN( u0_out0_6 ) , .A1( u0_u0_u2_n25 ) , .A2( u0_u0_u2_n26 ) , .A3( u0_u0_u2_n27 ) , .A4( u0_u0_u2_n28 ) );
  OR3_X1 u0_u0_u2_U95 (.ZN( u0_u0_u2_n28 ) , .A1( u0_u0_u2_n29 ) , .A2( u0_u0_u2_n30 ) , .A3( u0_u0_u2_n6 ) );
  AOI21_X1 u0_u0_u2_U96 (.A( u0_u0_u2_n22 ) , .ZN( u0_u0_u2_n30 ) , .B1( u0_u0_u2_n34 ) , .B2( u0_u0_u2_n35 ) );
  NAND3_X1 u0_u0_u2_U97 (.ZN( u0_u0_u2_n55 ) , .A3( u0_u0_u2_n66 ) , .A1( u0_u0_u2_n67 ) , .A2( u0_u0_u2_n72 ) );
  NAND3_X1 u0_u0_u2_U98 (.A1( u0_u0_u2_n35 ) , .A3( u0_u0_u2_n50 ) , .A2( u0_u0_u2_n58 ) , .ZN( u0_u0_u2_n79 ) );
  NAND3_X1 u0_u0_u2_U99 (.A3( u0_u0_u2_n75 ) , .A1( u0_u0_u2_n85 ) , .ZN( u0_u0_u2_n88 ) , .A2( u0_u0_u2_n89 ) );
  OAI22_X1 u0_u0_u3_U10 (.B2( u0_u0_u3_n23 ) , .A1( u0_u0_u3_n37 ) , .A2( u0_u0_u3_n52 ) , .B1( u0_u0_u3_n74 ) , .ZN( u0_u0_u3_n89 ) );
  OAI211_X1 u0_u0_u3_U11 (.C1( u0_u0_u3_n20 ) , .C2( u0_u0_u3_n59 ) , .A( u0_u0_u3_n6 ) , .ZN( u0_u0_u3_n68 ) , .B( u0_u0_u3_n81 ) );
  AOI221_X1 u0_u0_u3_U12 (.B1( u0_u0_u3_n18 ) , .C2( u0_u0_u3_n54 ) , .B2( u0_u0_u3_n55 ) , .A( u0_u0_u3_n56 ) , .ZN( u0_u0_u3_n81 ) , .C1( u0_u0_u3_n82 ) );
  INV_X1 u0_u0_u3_U13 (.ZN( u0_u0_u3_n6 ) , .A( u0_u0_u3_n89 ) );
  NAND2_X1 u0_u0_u3_U14 (.A1( u0_u0_u3_n32 ) , .A2( u0_u0_u3_n57 ) , .ZN( u0_u0_u3_n82 ) );
  AOI22_X1 u0_u0_u3_U15 (.A1( u0_u0_u3_n18 ) , .B2( u0_u0_u3_n54 ) , .ZN( u0_u0_u3_n64 ) , .A2( u0_u0_u3_n71 ) , .B1( u0_u0_u3_n72 ) );
  NAND2_X1 u0_u0_u3_U16 (.A2( u0_u0_u3_n36 ) , .A1( u0_u0_u3_n5 ) , .ZN( u0_u0_u3_n71 ) );
  NOR2_X1 u0_u0_u3_U17 (.A1( u0_u0_u3_n23 ) , .A2( u0_u0_u3_n37 ) , .ZN( u0_u0_u3_n61 ) );
  AOI21_X1 u0_u0_u3_U18 (.A( u0_u0_u3_n20 ) , .B1( u0_u0_u3_n32 ) , .B2( u0_u0_u3_n41 ) , .ZN( u0_u0_u3_n75 ) );
  NAND2_X1 u0_u0_u3_U19 (.A2( u0_u0_u3_n23 ) , .ZN( u0_u0_u3_n45 ) , .A1( u0_u0_u3_n52 ) );
  NAND2_X1 u0_u0_u3_U20 (.A1( u0_u0_u3_n31 ) , .A2( u0_u0_u3_n35 ) , .ZN( u0_u0_u3_n55 ) );
  INV_X1 u0_u0_u3_U21 (.ZN( u0_u0_u3_n22 ) , .A( u0_u0_u3_n54 ) );
  AND2_X1 u0_u0_u3_U22 (.ZN( u0_u0_u3_n36 ) , .A1( u0_u0_u3_n73 ) , .A2( u0_u0_u3_n74 ) );
  INV_X1 u0_u0_u3_U23 (.ZN( u0_u0_u3_n17 ) , .A( u0_u0_u3_n52 ) );
  NAND2_X1 u0_u0_u3_U24 (.ZN( u0_u0_u3_n47 ) , .A2( u0_u0_u3_n79 ) , .A1( u0_u0_u3_n80 ) );
  NAND2_X1 u0_u0_u3_U25 (.A2( u0_u0_u3_n39 ) , .A1( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n70 ) );
  NAND2_X1 u0_u0_u3_U26 (.A2( u0_u0_u3_n20 ) , .A1( u0_u0_u3_n22 ) , .ZN( u0_u0_u3_n44 ) );
  INV_X1 u0_u0_u3_U27 (.ZN( u0_u0_u3_n10 ) , .A( u0_u0_u3_n57 ) );
  INV_X1 u0_u0_u3_U28 (.ZN( u0_u0_u3_n11 ) , .A( u0_u0_u3_n59 ) );
  INV_X1 u0_u0_u3_U29 (.ZN( u0_u0_u3_n13 ) , .A( u0_u0_u3_n32 ) );
  INV_X1 u0_u0_u3_U3 (.A( u0_u0_u3_n47 ) , .ZN( u0_u0_u3_n5 ) );
  INV_X1 u0_u0_u3_U30 (.ZN( u0_u0_u3_n2 ) , .A( u0_u0_u3_n48 ) );
  NOR2_X1 u0_u0_u3_U31 (.A1( u0_u0_u3_n18 ) , .A2( u0_u0_u3_n46 ) , .ZN( u0_u0_u3_n52 ) );
  OAI222_X1 u0_u0_u3_U32 (.A1( u0_u0_u3_n23 ) , .C1( u0_u0_u3_n33 ) , .B2( u0_u0_u3_n41 ) , .ZN( u0_u0_u3_n49 ) , .B1( u0_u0_u3_n52 ) , .A2( u0_u0_u3_n79 ) , .C2( u0_u0_u3_n80 ) );
  NOR4_X1 u0_u0_u3_U33 (.ZN( u0_u0_u3_n26 ) , .A1( u0_u0_u3_n27 ) , .A2( u0_u0_u3_n28 ) , .A3( u0_u0_u3_n29 ) , .A4( u0_u0_u3_n30 ) );
  AOI21_X1 u0_u0_u3_U34 (.A( u0_u0_u3_n23 ) , .ZN( u0_u0_u3_n29 ) , .B1( u0_u0_u3_n34 ) , .B2( u0_u0_u3_n35 ) );
  AOI21_X1 u0_u0_u3_U35 (.ZN( u0_u0_u3_n30 ) , .B1( u0_u0_u3_n31 ) , .B2( u0_u0_u3_n32 ) , .A( u0_u0_u3_n33 ) );
  AOI21_X1 u0_u0_u3_U36 (.ZN( u0_u0_u3_n28 ) , .B1( u0_u0_u3_n36 ) , .B2( u0_u0_u3_n37 ) , .A( u0_u0_u3_n38 ) );
  OAI211_X1 u0_u0_u3_U37 (.A( u0_u0_u3_n3 ) , .C2( u0_u0_u3_n33 ) , .C1( u0_u0_u3_n37 ) , .ZN( u0_u0_u3_n48 ) , .B( u0_u0_u3_n60 ) );
  INV_X1 u0_u0_u3_U38 (.ZN( u0_u0_u3_n3 ) , .A( u0_u0_u3_n62 ) );
  AOI221_X1 u0_u0_u3_U39 (.B1( u0_u0_u3_n13 ) , .B2( u0_u0_u3_n17 ) , .C1( u0_u0_u3_n18 ) , .C2( u0_u0_u3_n55 ) , .ZN( u0_u0_u3_n60 ) , .A( u0_u0_u3_n61 ) );
  INV_X1 u0_u0_u3_U4 (.ZN( u0_u0_u3_n4 ) , .A( u0_u0_u3_n58 ) );
  OAI22_X1 u0_u0_u3_U40 (.B1( u0_u0_u3_n20 ) , .A2( u0_u0_u3_n22 ) , .B2( u0_u0_u3_n42 ) , .ZN( u0_u0_u3_n62 ) , .A1( u0_u0_u3_n63 ) );
  AOI211_X1 u0_u0_u3_U41 (.C1( u0_u0_u3_n46 ) , .B( u0_u0_u3_n49 ) , .C2( u0_u0_u3_n58 ) , .A( u0_u0_u3_n68 ) , .ZN( u0_u0_u3_n78 ) );
  AOI211_X1 u0_u0_u3_U42 (.ZN( u0_u0_u3_n65 ) , .C2( u0_u0_u3_n66 ) , .A( u0_u0_u3_n67 ) , .B( u0_u0_u3_n68 ) , .C1( u0_u0_u3_n8 ) );
  INV_X1 u0_u0_u3_U43 (.A( u0_u0_u3_n31 ) , .ZN( u0_u0_u3_n8 ) );
  OAI22_X1 u0_u0_u3_U44 (.B2( u0_u0_u3_n33 ) , .A1( u0_u0_u3_n52 ) , .ZN( u0_u0_u3_n67 ) , .B1( u0_u0_u3_n69 ) , .A2( u0_u0_u3_n9 ) );
  AND3_X1 u0_u0_u3_U45 (.A3( u0_u0_u3_n35 ) , .A1( u0_u0_u3_n43 ) , .A2( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n69 ) );
  INV_X1 u0_u0_u3_U46 (.ZN( u0_u0_u3_n23 ) , .A( u0_u0_u3_n66 ) );
  NAND2_X1 u0_u0_u3_U47 (.A2( u0_u0_u3_n23 ) , .A1( u0_u0_u3_n33 ) , .ZN( u0_u0_u3_n54 ) );
  NOR2_X1 u0_u0_u3_U48 (.A2( u0_u0_u3_n33 ) , .ZN( u0_u0_u3_n56 ) , .A1( u0_u0_u3_n74 ) );
  NAND2_X1 u0_u0_u3_U49 (.ZN( u0_u0_u3_n37 ) , .A1( u0_u0_u3_n84 ) , .A2( u0_u0_u3_n88 ) );
  INV_X1 u0_u0_u3_U5 (.A( u0_u0_u3_n70 ) , .ZN( u0_u0_u3_n9 ) );
  NAND2_X1 u0_u0_u3_U50 (.ZN( u0_u0_u3_n32 ) , .A2( u0_u0_u3_n85 ) , .A1( u0_u0_u3_n90 ) );
  INV_X1 u0_u0_u3_U51 (.ZN( u0_u0_u3_n20 ) , .A( u0_u0_u3_n46 ) );
  AOI21_X1 u0_u0_u3_U52 (.A( u0_u0_u3_n33 ) , .B1( u0_u0_u3_n41 ) , .B2( u0_u0_u3_n73 ) , .ZN( u0_u0_u3_n93 ) );
  AOI21_X1 u0_u0_u3_U53 (.B1( u0_u0_u3_n1 ) , .B2( u0_u0_u3_n45 ) , .ZN( u0_u0_u3_n77 ) , .A( u0_u0_u3_n92 ) );
  INV_X1 u0_u0_u3_U54 (.ZN( u0_u0_u3_n1 ) , .A( u0_u0_u3_n42 ) );
  AOI21_X1 u0_u0_u3_U55 (.B2( u0_u0_u3_n32 ) , .A( u0_u0_u3_n38 ) , .B1( u0_u0_u3_n63 ) , .ZN( u0_u0_u3_n92 ) );
  INV_X1 u0_u0_u3_U56 (.ZN( u0_u0_u3_n18 ) , .A( u0_u0_u3_n38 ) );
  NAND2_X1 u0_u0_u3_U57 (.ZN( u0_u0_u3_n63 ) , .A2( u0_u0_u3_n90 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U58 (.ZN( u0_u0_u3_n41 ) , .A2( u0_u0_u3_n87 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U59 (.ZN( u0_u0_u3_n42 ) , .A1( u0_u0_u3_n86 ) , .A2( u0_u0_u3_n88 ) );
  AOI221_X1 u0_u0_u3_U6 (.B2( u0_u0_u3_n10 ) , .B1( u0_u0_u3_n44 ) , .ZN( u0_u0_u3_n53 ) , .C1( u0_u0_u3_n54 ) , .C2( u0_u0_u3_n55 ) , .A( u0_u0_u3_n56 ) );
  NAND2_X1 u0_u0_u3_U60 (.ZN( u0_u0_u3_n31 ) , .A1( u0_u0_u3_n87 ) , .A2( u0_u0_u3_n88 ) );
  NAND2_X1 u0_u0_u3_U61 (.ZN( u0_u0_u3_n39 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n86 ) );
  NAND2_X1 u0_u0_u3_U62 (.ZN( u0_u0_u3_n59 ) , .A2( u0_u0_u3_n85 ) , .A1( u0_u0_u3_n87 ) );
  NAND2_X1 u0_u0_u3_U63 (.ZN( u0_u0_u3_n35 ) , .A1( u0_u0_u3_n85 ) , .A2( u0_u0_u3_n86 ) );
  NAND2_X1 u0_u0_u3_U64 (.ZN( u0_u0_u3_n73 ) , .A2( u0_u0_u3_n86 ) , .A1( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U65 (.ZN( u0_u0_u3_n80 ) , .A2( u0_u0_u3_n88 ) , .A1( u0_u0_u3_n90 ) );
  NAND2_X1 u0_u0_u3_U66 (.ZN( u0_u0_u3_n74 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n87 ) );
  NAND2_X1 u0_u0_u3_U67 (.ZN( u0_u0_u3_n34 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n90 ) );
  NAND2_X1 u0_u0_u3_U68 (.ZN( u0_u0_u3_n57 ) , .A1( u0_u0_u3_n83 ) , .A2( u0_u0_u3_n84 ) );
  NAND2_X1 u0_u0_u3_U69 (.ZN( u0_u0_u3_n43 ) , .A2( u0_u0_u3_n84 ) , .A1( u0_u0_u3_n91 ) );
  OAI22_X1 u0_u0_u3_U7 (.A1( u0_u0_u3_n19 ) , .B1( u0_u0_u3_n22 ) , .ZN( u0_u0_u3_n27 ) , .A2( u0_u0_u3_n39 ) , .B2( u0_u0_u3_n40 ) );
  NAND2_X1 u0_u0_u3_U70 (.ZN( u0_u0_u3_n79 ) , .A2( u0_u0_u3_n84 ) , .A1( u0_u0_u3_n85 ) );
  NOR2_X1 u0_u0_u3_U71 (.A2( u0_u0_X_19 ) , .A1( u0_u0_X_20 ) , .ZN( u0_u0_u3_n88 ) );
  NOR2_X1 u0_u0_u3_U72 (.A2( u0_u0_X_21 ) , .A1( u0_u0_X_24 ) , .ZN( u0_u0_u3_n84 ) );
  NOR2_X1 u0_u0_u3_U73 (.A2( u0_u0_X_24 ) , .A1( u0_u0_u3_n16 ) , .ZN( u0_u0_u3_n90 ) );
  NOR2_X1 u0_u0_u3_U74 (.A2( u0_u0_X_23 ) , .A1( u0_u0_u3_n21 ) , .ZN( u0_u0_u3_n46 ) );
  NOR2_X1 u0_u0_u3_U75 (.A2( u0_u0_X_19 ) , .A1( u0_u0_u3_n15 ) , .ZN( u0_u0_u3_n91 ) );
  NAND2_X1 u0_u0_u3_U76 (.A1( u0_u0_X_22 ) , .A2( u0_u0_X_23 ) , .ZN( u0_u0_u3_n33 ) );
  NAND2_X1 u0_u0_u3_U77 (.A1( u0_u0_X_23 ) , .A2( u0_u0_u3_n21 ) , .ZN( u0_u0_u3_n38 ) );
  NOR2_X1 u0_u0_u3_U78 (.A2( u0_u0_X_22 ) , .A1( u0_u0_X_23 ) , .ZN( u0_u0_u3_n66 ) );
  AND2_X1 u0_u0_u3_U79 (.A1( u0_u0_X_24 ) , .A2( u0_u0_u3_n16 ) , .ZN( u0_u0_u3_n86 ) );
  AND3_X1 u0_u0_u3_U8 (.ZN( u0_u0_u3_n40 ) , .A1( u0_u0_u3_n41 ) , .A2( u0_u0_u3_n42 ) , .A3( u0_u0_u3_n43 ) );
  AND2_X1 u0_u0_u3_U80 (.A1( u0_u0_X_19 ) , .A2( u0_u0_u3_n15 ) , .ZN( u0_u0_u3_n85 ) );
  AND2_X1 u0_u0_u3_U81 (.A1( u0_u0_X_21 ) , .A2( u0_u0_X_24 ) , .ZN( u0_u0_u3_n87 ) );
  AND2_X1 u0_u0_u3_U82 (.A2( u0_u0_X_19 ) , .A1( u0_u0_X_20 ) , .ZN( u0_u0_u3_n83 ) );
  INV_X1 u0_u0_u3_U83 (.A( u0_u0_X_22 ) , .ZN( u0_u0_u3_n21 ) );
  INV_X1 u0_u0_u3_U84 (.A( u0_u0_X_21 ) , .ZN( u0_u0_u3_n16 ) );
  INV_X1 u0_u0_u3_U85 (.A( u0_u0_X_20 ) , .ZN( u0_u0_u3_n15 ) );
  NAND4_X1 u0_u0_u3_U86 (.ZN( u0_out0_26 ) , .A1( u0_u0_u3_n14 ) , .A2( u0_u0_u3_n76 ) , .A3( u0_u0_u3_n77 ) , .A4( u0_u0_u3_n78 ) );
  INV_X1 u0_u0_u3_U87 (.ZN( u0_u0_u3_n14 ) , .A( u0_u0_u3_n93 ) );
  OAI21_X1 u0_u0_u3_U88 (.B1( u0_u0_u3_n11 ) , .A( u0_u0_u3_n54 ) , .B2( u0_u0_u3_n70 ) , .ZN( u0_u0_u3_n76 ) );
  NAND4_X1 u0_u0_u3_U89 (.ZN( u0_out0_1 ) , .A1( u0_u0_u3_n2 ) , .A2( u0_u0_u3_n24 ) , .A3( u0_u0_u3_n25 ) , .A4( u0_u0_u3_n26 ) );
  INV_X1 u0_u0_u3_U9 (.ZN( u0_u0_u3_n19 ) , .A( u0_u0_u3_n44 ) );
  NAND2_X1 u0_u0_u3_U90 (.A1( u0_u0_u3_n11 ) , .A2( u0_u0_u3_n17 ) , .ZN( u0_u0_u3_n24 ) );
  AOI22_X1 u0_u0_u3_U91 (.A1( u0_u0_u3_n10 ) , .ZN( u0_u0_u3_n25 ) , .A2( u0_u0_u3_n45 ) , .B1( u0_u0_u3_n46 ) , .B2( u0_u0_u3_n47 ) );
  NAND4_X1 u0_u0_u3_U92 (.ZN( u0_out0_20 ) , .A1( u0_u0_u3_n12 ) , .A3( u0_u0_u3_n64 ) , .A4( u0_u0_u3_n65 ) , .A2( u0_u0_u3_n7 ) );
  INV_X1 u0_u0_u3_U93 (.A( u0_u0_u3_n61 ) , .ZN( u0_u0_u3_n7 ) );
  INV_X1 u0_u0_u3_U94 (.ZN( u0_u0_u3_n12 ) , .A( u0_u0_u3_n75 ) );
  OR4_X1 u0_u0_u3_U95 (.ZN( u0_out0_10 ) , .A2( u0_u0_u3_n48 ) , .A1( u0_u0_u3_n49 ) , .A3( u0_u0_u3_n50 ) , .A4( u0_u0_u3_n51 ) );
  OAI222_X1 u0_u0_u3_U96 (.A1( u0_u0_u3_n20 ) , .C2( u0_u0_u3_n23 ) , .B2( u0_u0_u3_n33 ) , .A2( u0_u0_u3_n37 ) , .B1( u0_u0_u3_n39 ) , .ZN( u0_u0_u3_n50 ) , .C1( u0_u0_u3_n59 ) );
  OAI221_X1 u0_u0_u3_U97 (.B1( u0_u0_u3_n36 ) , .C1( u0_u0_u3_n38 ) , .C2( u0_u0_u3_n4 ) , .ZN( u0_u0_u3_n51 ) , .B2( u0_u0_u3_n52 ) , .A( u0_u0_u3_n53 ) );
  NAND3_X1 u0_u0_u3_U98 (.A3( u0_u0_u3_n34 ) , .A2( u0_u0_u3_n42 ) , .ZN( u0_u0_u3_n72 ) , .A1( u0_u0_u3_n73 ) );
  NAND3_X1 u0_u0_u3_U99 (.A1( u0_u0_u3_n34 ) , .A2( u0_u0_u3_n43 ) , .A3( u0_u0_u3_n5 ) , .ZN( u0_u0_u3_n58 ) );
  XOR2_X1 u0_u10_U1 (.B( u0_K11_9 ) , .A( u0_R9_6 ) , .Z( u0_u10_X_9 ) );
  XOR2_X1 u0_u10_U2 (.B( u0_K11_8 ) , .A( u0_R9_5 ) , .Z( u0_u10_X_8 ) );
  XOR2_X1 u0_u10_U3 (.B( u0_K11_7 ) , .A( u0_R9_4 ) , .Z( u0_u10_X_7 ) );
  XOR2_X1 u0_u10_U33 (.B( u0_K11_24 ) , .A( u0_R9_17 ) , .Z( u0_u10_X_24 ) );
  XOR2_X1 u0_u10_U34 (.B( u0_K11_23 ) , .A( u0_R9_16 ) , .Z( u0_u10_X_23 ) );
  XOR2_X1 u0_u10_U37 (.B( u0_K11_20 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_20 ) );
  XOR2_X1 u0_u10_U39 (.B( u0_K11_19 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_19 ) );
  XOR2_X1 u0_u10_U40 (.B( u0_K11_18 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_18 ) );
  XOR2_X1 u0_u10_U41 (.B( u0_K11_17 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_17 ) );
  XOR2_X1 u0_u10_U42 (.B( u0_K11_16 ) , .A( u0_R9_11 ) , .Z( u0_u10_X_16 ) );
  XOR2_X1 u0_u10_U43 (.B( u0_K11_15 ) , .A( u0_R9_10 ) , .Z( u0_u10_X_15 ) );
  XOR2_X1 u0_u10_U44 (.B( u0_K11_14 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_14 ) );
  XOR2_X1 u0_u10_U45 (.B( u0_K11_13 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_13 ) );
  XOR2_X1 u0_u10_U46 (.B( u0_K11_12 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_12 ) );
  XOR2_X1 u0_u10_U47 (.B( u0_K11_11 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_11 ) );
  XOR2_X1 u0_u10_U48 (.B( u0_K11_10 ) , .A( u0_R9_7 ) , .Z( u0_u10_X_10 ) );
  AOI21_X1 u0_u10_u1_U10 (.B2( u0_u10_u1_n155 ) , .B1( u0_u10_u1_n156 ) , .ZN( u0_u10_u1_n157 ) , .A( u0_u10_u1_n174 ) );
  NAND3_X1 u0_u10_u1_U100 (.ZN( u0_u10_u1_n113 ) , .A1( u0_u10_u1_n120 ) , .A3( u0_u10_u1_n133 ) , .A2( u0_u10_u1_n155 ) );
  NAND2_X1 u0_u10_u1_U11 (.ZN( u0_u10_u1_n140 ) , .A2( u0_u10_u1_n150 ) , .A1( u0_u10_u1_n155 ) );
  NAND2_X1 u0_u10_u1_U12 (.A1( u0_u10_u1_n131 ) , .ZN( u0_u10_u1_n147 ) , .A2( u0_u10_u1_n153 ) );
  AOI22_X1 u0_u10_u1_U13 (.B2( u0_u10_u1_n136 ) , .A2( u0_u10_u1_n137 ) , .ZN( u0_u10_u1_n143 ) , .A1( u0_u10_u1_n171 ) , .B1( u0_u10_u1_n173 ) );
  INV_X1 u0_u10_u1_U14 (.A( u0_u10_u1_n147 ) , .ZN( u0_u10_u1_n181 ) );
  INV_X1 u0_u10_u1_U15 (.A( u0_u10_u1_n139 ) , .ZN( u0_u10_u1_n174 ) );
  OR4_X1 u0_u10_u1_U16 (.A4( u0_u10_u1_n106 ) , .A3( u0_u10_u1_n107 ) , .ZN( u0_u10_u1_n108 ) , .A1( u0_u10_u1_n117 ) , .A2( u0_u10_u1_n184 ) );
  AOI21_X1 u0_u10_u1_U17 (.ZN( u0_u10_u1_n106 ) , .A( u0_u10_u1_n112 ) , .B1( u0_u10_u1_n154 ) , .B2( u0_u10_u1_n156 ) );
  AOI21_X1 u0_u10_u1_U18 (.ZN( u0_u10_u1_n107 ) , .B1( u0_u10_u1_n134 ) , .B2( u0_u10_u1_n149 ) , .A( u0_u10_u1_n174 ) );
  INV_X1 u0_u10_u1_U19 (.A( u0_u10_u1_n101 ) , .ZN( u0_u10_u1_n184 ) );
  INV_X1 u0_u10_u1_U20 (.A( u0_u10_u1_n112 ) , .ZN( u0_u10_u1_n171 ) );
  NAND2_X1 u0_u10_u1_U21 (.ZN( u0_u10_u1_n141 ) , .A1( u0_u10_u1_n153 ) , .A2( u0_u10_u1_n156 ) );
  AND2_X1 u0_u10_u1_U22 (.A1( u0_u10_u1_n123 ) , .ZN( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n161 ) );
  NAND2_X1 u0_u10_u1_U23 (.A2( u0_u10_u1_n115 ) , .A1( u0_u10_u1_n116 ) , .ZN( u0_u10_u1_n148 ) );
  NAND2_X1 u0_u10_u1_U24 (.A2( u0_u10_u1_n133 ) , .A1( u0_u10_u1_n135 ) , .ZN( u0_u10_u1_n159 ) );
  NAND2_X1 u0_u10_u1_U25 (.A2( u0_u10_u1_n115 ) , .A1( u0_u10_u1_n120 ) , .ZN( u0_u10_u1_n132 ) );
  INV_X1 u0_u10_u1_U26 (.A( u0_u10_u1_n154 ) , .ZN( u0_u10_u1_n178 ) );
  INV_X1 u0_u10_u1_U27 (.A( u0_u10_u1_n151 ) , .ZN( u0_u10_u1_n183 ) );
  AND2_X1 u0_u10_u1_U28 (.A1( u0_u10_u1_n129 ) , .A2( u0_u10_u1_n133 ) , .ZN( u0_u10_u1_n149 ) );
  INV_X1 u0_u10_u1_U29 (.A( u0_u10_u1_n131 ) , .ZN( u0_u10_u1_n180 ) );
  INV_X1 u0_u10_u1_U3 (.A( u0_u10_u1_n159 ) , .ZN( u0_u10_u1_n182 ) );
  OAI221_X1 u0_u10_u1_U30 (.A( u0_u10_u1_n119 ) , .C2( u0_u10_u1_n129 ) , .ZN( u0_u10_u1_n138 ) , .B2( u0_u10_u1_n152 ) , .C1( u0_u10_u1_n174 ) , .B1( u0_u10_u1_n187 ) );
  INV_X1 u0_u10_u1_U31 (.A( u0_u10_u1_n148 ) , .ZN( u0_u10_u1_n187 ) );
  AOI211_X1 u0_u10_u1_U32 (.B( u0_u10_u1_n117 ) , .A( u0_u10_u1_n118 ) , .ZN( u0_u10_u1_n119 ) , .C2( u0_u10_u1_n146 ) , .C1( u0_u10_u1_n159 ) );
  NOR2_X1 u0_u10_u1_U33 (.A1( u0_u10_u1_n168 ) , .A2( u0_u10_u1_n176 ) , .ZN( u0_u10_u1_n98 ) );
  OAI21_X1 u0_u10_u1_U34 (.B2( u0_u10_u1_n123 ) , .ZN( u0_u10_u1_n145 ) , .B1( u0_u10_u1_n160 ) , .A( u0_u10_u1_n185 ) );
  INV_X1 u0_u10_u1_U35 (.A( u0_u10_u1_n122 ) , .ZN( u0_u10_u1_n185 ) );
  AOI21_X1 u0_u10_u1_U36 (.B2( u0_u10_u1_n120 ) , .B1( u0_u10_u1_n121 ) , .ZN( u0_u10_u1_n122 ) , .A( u0_u10_u1_n128 ) );
  NAND2_X1 u0_u10_u1_U37 (.A1( u0_u10_u1_n128 ) , .ZN( u0_u10_u1_n146 ) , .A2( u0_u10_u1_n160 ) );
  NAND2_X1 u0_u10_u1_U38 (.A2( u0_u10_u1_n112 ) , .ZN( u0_u10_u1_n139 ) , .A1( u0_u10_u1_n152 ) );
  NAND2_X1 u0_u10_u1_U39 (.A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n156 ) , .A2( u0_u10_u1_n99 ) );
  AOI221_X1 u0_u10_u1_U4 (.A( u0_u10_u1_n138 ) , .C2( u0_u10_u1_n139 ) , .C1( u0_u10_u1_n140 ) , .B2( u0_u10_u1_n141 ) , .ZN( u0_u10_u1_n142 ) , .B1( u0_u10_u1_n175 ) );
  AOI221_X1 u0_u10_u1_U40 (.B1( u0_u10_u1_n140 ) , .ZN( u0_u10_u1_n167 ) , .B2( u0_u10_u1_n172 ) , .C2( u0_u10_u1_n175 ) , .C1( u0_u10_u1_n178 ) , .A( u0_u10_u1_n188 ) );
  INV_X1 u0_u10_u1_U41 (.ZN( u0_u10_u1_n188 ) , .A( u0_u10_u1_n97 ) );
  AOI211_X1 u0_u10_u1_U42 (.A( u0_u10_u1_n118 ) , .C1( u0_u10_u1_n132 ) , .C2( u0_u10_u1_n139 ) , .B( u0_u10_u1_n96 ) , .ZN( u0_u10_u1_n97 ) );
  AOI21_X1 u0_u10_u1_U43 (.B2( u0_u10_u1_n121 ) , .B1( u0_u10_u1_n135 ) , .A( u0_u10_u1_n152 ) , .ZN( u0_u10_u1_n96 ) );
  NOR2_X1 u0_u10_u1_U44 (.ZN( u0_u10_u1_n117 ) , .A1( u0_u10_u1_n121 ) , .A2( u0_u10_u1_n160 ) );
  AOI21_X1 u0_u10_u1_U45 (.A( u0_u10_u1_n128 ) , .B2( u0_u10_u1_n129 ) , .ZN( u0_u10_u1_n130 ) , .B1( u0_u10_u1_n150 ) );
  NAND2_X1 u0_u10_u1_U46 (.ZN( u0_u10_u1_n112 ) , .A1( u0_u10_u1_n169 ) , .A2( u0_u10_u1_n170 ) );
  NAND2_X1 u0_u10_u1_U47 (.ZN( u0_u10_u1_n129 ) , .A2( u0_u10_u1_n95 ) , .A1( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U48 (.A1( u0_u10_u1_n102 ) , .ZN( u0_u10_u1_n154 ) , .A2( u0_u10_u1_n99 ) );
  NAND2_X1 u0_u10_u1_U49 (.A2( u0_u10_u1_n100 ) , .ZN( u0_u10_u1_n135 ) , .A1( u0_u10_u1_n99 ) );
  AOI211_X1 u0_u10_u1_U5 (.ZN( u0_u10_u1_n124 ) , .A( u0_u10_u1_n138 ) , .C2( u0_u10_u1_n139 ) , .B( u0_u10_u1_n145 ) , .C1( u0_u10_u1_n147 ) );
  AOI21_X1 u0_u10_u1_U50 (.A( u0_u10_u1_n152 ) , .B2( u0_u10_u1_n153 ) , .B1( u0_u10_u1_n154 ) , .ZN( u0_u10_u1_n158 ) );
  INV_X1 u0_u10_u1_U51 (.A( u0_u10_u1_n160 ) , .ZN( u0_u10_u1_n175 ) );
  NAND2_X1 u0_u10_u1_U52 (.A1( u0_u10_u1_n100 ) , .ZN( u0_u10_u1_n116 ) , .A2( u0_u10_u1_n95 ) );
  NAND2_X1 u0_u10_u1_U53 (.A1( u0_u10_u1_n102 ) , .ZN( u0_u10_u1_n131 ) , .A2( u0_u10_u1_n95 ) );
  NAND2_X1 u0_u10_u1_U54 (.A2( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n121 ) , .A1( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U55 (.A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n153 ) , .A2( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U56 (.A2( u0_u10_u1_n104 ) , .A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n133 ) );
  NAND2_X1 u0_u10_u1_U57 (.ZN( u0_u10_u1_n150 ) , .A2( u0_u10_u1_n98 ) , .A1( u0_u10_u1_n99 ) );
  NAND2_X1 u0_u10_u1_U58 (.A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n155 ) , .A2( u0_u10_u1_n95 ) );
  OAI21_X1 u0_u10_u1_U59 (.ZN( u0_u10_u1_n109 ) , .B1( u0_u10_u1_n129 ) , .B2( u0_u10_u1_n160 ) , .A( u0_u10_u1_n167 ) );
  AOI22_X1 u0_u10_u1_U6 (.B2( u0_u10_u1_n113 ) , .A2( u0_u10_u1_n114 ) , .ZN( u0_u10_u1_n125 ) , .A1( u0_u10_u1_n171 ) , .B1( u0_u10_u1_n173 ) );
  NAND2_X1 u0_u10_u1_U60 (.A2( u0_u10_u1_n100 ) , .A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n120 ) );
  NAND2_X1 u0_u10_u1_U61 (.A1( u0_u10_u1_n102 ) , .A2( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n115 ) );
  NAND2_X1 u0_u10_u1_U62 (.A2( u0_u10_u1_n100 ) , .A1( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n151 ) );
  NAND2_X1 u0_u10_u1_U63 (.A2( u0_u10_u1_n103 ) , .A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n161 ) );
  INV_X1 u0_u10_u1_U64 (.A( u0_u10_u1_n152 ) , .ZN( u0_u10_u1_n173 ) );
  INV_X1 u0_u10_u1_U65 (.A( u0_u10_u1_n128 ) , .ZN( u0_u10_u1_n172 ) );
  NAND2_X1 u0_u10_u1_U66 (.A2( u0_u10_u1_n102 ) , .A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n123 ) );
  AOI211_X1 u0_u10_u1_U67 (.B( u0_u10_u1_n162 ) , .A( u0_u10_u1_n163 ) , .C2( u0_u10_u1_n164 ) , .ZN( u0_u10_u1_n165 ) , .C1( u0_u10_u1_n171 ) );
  AOI21_X1 u0_u10_u1_U68 (.A( u0_u10_u1_n160 ) , .B2( u0_u10_u1_n161 ) , .ZN( u0_u10_u1_n162 ) , .B1( u0_u10_u1_n182 ) );
  OR2_X1 u0_u10_u1_U69 (.A2( u0_u10_u1_n157 ) , .A1( u0_u10_u1_n158 ) , .ZN( u0_u10_u1_n163 ) );
  NAND2_X1 u0_u10_u1_U7 (.ZN( u0_u10_u1_n114 ) , .A1( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n156 ) );
  NOR2_X1 u0_u10_u1_U70 (.A2( u0_u10_X_7 ) , .A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n95 ) );
  NOR2_X1 u0_u10_u1_U71 (.A1( u0_u10_X_12 ) , .A2( u0_u10_X_9 ) , .ZN( u0_u10_u1_n100 ) );
  NOR2_X1 u0_u10_u1_U72 (.A2( u0_u10_X_8 ) , .A1( u0_u10_u1_n177 ) , .ZN( u0_u10_u1_n99 ) );
  NOR2_X1 u0_u10_u1_U73 (.A2( u0_u10_X_12 ) , .ZN( u0_u10_u1_n102 ) , .A1( u0_u10_u1_n176 ) );
  NOR2_X1 u0_u10_u1_U74 (.A2( u0_u10_X_9 ) , .ZN( u0_u10_u1_n105 ) , .A1( u0_u10_u1_n168 ) );
  NAND2_X1 u0_u10_u1_U75 (.A1( u0_u10_X_10 ) , .ZN( u0_u10_u1_n160 ) , .A2( u0_u10_u1_n169 ) );
  NAND2_X1 u0_u10_u1_U76 (.A2( u0_u10_X_10 ) , .A1( u0_u10_X_11 ) , .ZN( u0_u10_u1_n152 ) );
  NAND2_X1 u0_u10_u1_U77 (.A1( u0_u10_X_11 ) , .ZN( u0_u10_u1_n128 ) , .A2( u0_u10_u1_n170 ) );
  AND2_X1 u0_u10_u1_U78 (.A2( u0_u10_X_7 ) , .A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n104 ) );
  AND2_X1 u0_u10_u1_U79 (.A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n103 ) , .A2( u0_u10_u1_n177 ) );
  NOR2_X1 u0_u10_u1_U8 (.A1( u0_u10_u1_n112 ) , .A2( u0_u10_u1_n116 ) , .ZN( u0_u10_u1_n118 ) );
  INV_X1 u0_u10_u1_U80 (.A( u0_u10_X_10 ) , .ZN( u0_u10_u1_n170 ) );
  INV_X1 u0_u10_u1_U81 (.A( u0_u10_X_9 ) , .ZN( u0_u10_u1_n176 ) );
  INV_X1 u0_u10_u1_U82 (.A( u0_u10_X_11 ) , .ZN( u0_u10_u1_n169 ) );
  INV_X1 u0_u10_u1_U83 (.A( u0_u10_X_12 ) , .ZN( u0_u10_u1_n168 ) );
  INV_X1 u0_u10_u1_U84 (.A( u0_u10_X_7 ) , .ZN( u0_u10_u1_n177 ) );
  NAND4_X1 u0_u10_u1_U85 (.ZN( u0_out10_28 ) , .A4( u0_u10_u1_n124 ) , .A3( u0_u10_u1_n125 ) , .A2( u0_u10_u1_n126 ) , .A1( u0_u10_u1_n127 ) );
  OAI21_X1 u0_u10_u1_U86 (.ZN( u0_u10_u1_n127 ) , .B2( u0_u10_u1_n139 ) , .B1( u0_u10_u1_n175 ) , .A( u0_u10_u1_n183 ) );
  OAI21_X1 u0_u10_u1_U87 (.ZN( u0_u10_u1_n126 ) , .B2( u0_u10_u1_n140 ) , .A( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n178 ) );
  NAND4_X1 u0_u10_u1_U88 (.ZN( u0_out10_18 ) , .A4( u0_u10_u1_n165 ) , .A3( u0_u10_u1_n166 ) , .A1( u0_u10_u1_n167 ) , .A2( u0_u10_u1_n186 ) );
  AOI22_X1 u0_u10_u1_U89 (.B2( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n147 ) , .A2( u0_u10_u1_n148 ) , .ZN( u0_u10_u1_n166 ) , .A1( u0_u10_u1_n172 ) );
  OAI21_X1 u0_u10_u1_U9 (.ZN( u0_u10_u1_n101 ) , .B1( u0_u10_u1_n141 ) , .A( u0_u10_u1_n146 ) , .B2( u0_u10_u1_n183 ) );
  INV_X1 u0_u10_u1_U90 (.A( u0_u10_u1_n145 ) , .ZN( u0_u10_u1_n186 ) );
  NAND4_X1 u0_u10_u1_U91 (.ZN( u0_out10_2 ) , .A4( u0_u10_u1_n142 ) , .A3( u0_u10_u1_n143 ) , .A2( u0_u10_u1_n144 ) , .A1( u0_u10_u1_n179 ) );
  OAI21_X1 u0_u10_u1_U92 (.B2( u0_u10_u1_n132 ) , .ZN( u0_u10_u1_n144 ) , .A( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n180 ) );
  INV_X1 u0_u10_u1_U93 (.A( u0_u10_u1_n130 ) , .ZN( u0_u10_u1_n179 ) );
  OR4_X1 u0_u10_u1_U94 (.ZN( u0_out10_13 ) , .A4( u0_u10_u1_n108 ) , .A3( u0_u10_u1_n109 ) , .A2( u0_u10_u1_n110 ) , .A1( u0_u10_u1_n111 ) );
  AOI21_X1 u0_u10_u1_U95 (.ZN( u0_u10_u1_n111 ) , .A( u0_u10_u1_n128 ) , .B2( u0_u10_u1_n131 ) , .B1( u0_u10_u1_n135 ) );
  AOI21_X1 u0_u10_u1_U96 (.ZN( u0_u10_u1_n110 ) , .A( u0_u10_u1_n116 ) , .B1( u0_u10_u1_n152 ) , .B2( u0_u10_u1_n160 ) );
  NAND3_X1 u0_u10_u1_U97 (.A3( u0_u10_u1_n149 ) , .A2( u0_u10_u1_n150 ) , .A1( u0_u10_u1_n151 ) , .ZN( u0_u10_u1_n164 ) );
  NAND3_X1 u0_u10_u1_U98 (.A3( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n135 ) , .ZN( u0_u10_u1_n136 ) , .A1( u0_u10_u1_n151 ) );
  NAND3_X1 u0_u10_u1_U99 (.A1( u0_u10_u1_n133 ) , .ZN( u0_u10_u1_n137 ) , .A2( u0_u10_u1_n154 ) , .A3( u0_u10_u1_n181 ) );
  OAI22_X1 u0_u10_u2_U10 (.ZN( u0_u10_u2_n109 ) , .A2( u0_u10_u2_n113 ) , .B2( u0_u10_u2_n133 ) , .B1( u0_u10_u2_n167 ) , .A1( u0_u10_u2_n168 ) );
  NAND3_X1 u0_u10_u2_U100 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n98 ) );
  OAI22_X1 u0_u10_u2_U11 (.B1( u0_u10_u2_n151 ) , .A2( u0_u10_u2_n152 ) , .A1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n160 ) , .B2( u0_u10_u2_n168 ) );
  NOR3_X1 u0_u10_u2_U12 (.A1( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n151 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U13 (.ZN( u0_u10_u2_n144 ) , .B2( u0_u10_u2_n155 ) , .A( u0_u10_u2_n172 ) , .B1( u0_u10_u2_n185 ) );
  AOI21_X1 u0_u10_u2_U14 (.B2( u0_u10_u2_n143 ) , .ZN( u0_u10_u2_n145 ) , .B1( u0_u10_u2_n152 ) , .A( u0_u10_u2_n171 ) );
  AOI21_X1 u0_u10_u2_U15 (.B2( u0_u10_u2_n120 ) , .B1( u0_u10_u2_n121 ) , .ZN( u0_u10_u2_n126 ) , .A( u0_u10_u2_n167 ) );
  INV_X1 u0_u10_u2_U16 (.A( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n171 ) );
  INV_X1 u0_u10_u2_U17 (.A( u0_u10_u2_n120 ) , .ZN( u0_u10_u2_n188 ) );
  NAND2_X1 u0_u10_u2_U18 (.A2( u0_u10_u2_n122 ) , .ZN( u0_u10_u2_n150 ) , .A1( u0_u10_u2_n152 ) );
  INV_X1 u0_u10_u2_U19 (.A( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U20 (.A( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n173 ) );
  NAND2_X1 u0_u10_u2_U21 (.A1( u0_u10_u2_n132 ) , .A2( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n157 ) );
  INV_X1 u0_u10_u2_U22 (.A( u0_u10_u2_n113 ) , .ZN( u0_u10_u2_n178 ) );
  INV_X1 u0_u10_u2_U23 (.A( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n175 ) );
  INV_X1 u0_u10_u2_U24 (.A( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n181 ) );
  INV_X1 u0_u10_u2_U25 (.A( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n177 ) );
  INV_X1 u0_u10_u2_U26 (.A( u0_u10_u2_n116 ) , .ZN( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U27 (.A( u0_u10_u2_n131 ) , .ZN( u0_u10_u2_n179 ) );
  INV_X1 u0_u10_u2_U28 (.A( u0_u10_u2_n154 ) , .ZN( u0_u10_u2_n176 ) );
  NAND2_X1 u0_u10_u2_U29 (.A2( u0_u10_u2_n116 ) , .A1( u0_u10_u2_n117 ) , .ZN( u0_u10_u2_n118 ) );
  NOR2_X1 u0_u10_u2_U3 (.ZN( u0_u10_u2_n121 ) , .A2( u0_u10_u2_n177 ) , .A1( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U30 (.A( u0_u10_u2_n132 ) , .ZN( u0_u10_u2_n182 ) );
  INV_X1 u0_u10_u2_U31 (.A( u0_u10_u2_n158 ) , .ZN( u0_u10_u2_n183 ) );
  OAI21_X1 u0_u10_u2_U32 (.A( u0_u10_u2_n156 ) , .B1( u0_u10_u2_n157 ) , .ZN( u0_u10_u2_n158 ) , .B2( u0_u10_u2_n179 ) );
  NOR2_X1 u0_u10_u2_U33 (.ZN( u0_u10_u2_n156 ) , .A1( u0_u10_u2_n166 ) , .A2( u0_u10_u2_n169 ) );
  NOR2_X1 u0_u10_u2_U34 (.A2( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n140 ) );
  NOR2_X1 u0_u10_u2_U35 (.A2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n153 ) , .A1( u0_u10_u2_n156 ) );
  AOI211_X1 u0_u10_u2_U36 (.ZN( u0_u10_u2_n130 ) , .C1( u0_u10_u2_n138 ) , .C2( u0_u10_u2_n179 ) , .B( u0_u10_u2_n96 ) , .A( u0_u10_u2_n97 ) );
  OAI22_X1 u0_u10_u2_U37 (.B1( u0_u10_u2_n133 ) , .A2( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n152 ) , .B2( u0_u10_u2_n168 ) , .ZN( u0_u10_u2_n97 ) );
  OAI221_X1 u0_u10_u2_U38 (.B1( u0_u10_u2_n113 ) , .C1( u0_u10_u2_n132 ) , .A( u0_u10_u2_n149 ) , .B2( u0_u10_u2_n171 ) , .C2( u0_u10_u2_n172 ) , .ZN( u0_u10_u2_n96 ) );
  OAI221_X1 u0_u10_u2_U39 (.A( u0_u10_u2_n115 ) , .C2( u0_u10_u2_n123 ) , .B2( u0_u10_u2_n143 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n163 ) , .C1( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U4 (.A( u0_u10_u2_n134 ) , .ZN( u0_u10_u2_n185 ) );
  OAI21_X1 u0_u10_u2_U40 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n115 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n178 ) );
  OAI221_X1 u0_u10_u2_U41 (.A( u0_u10_u2_n135 ) , .B2( u0_u10_u2_n136 ) , .B1( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n162 ) , .C2( u0_u10_u2_n167 ) , .C1( u0_u10_u2_n185 ) );
  AND3_X1 u0_u10_u2_U42 (.A3( u0_u10_u2_n131 ) , .A2( u0_u10_u2_n132 ) , .A1( u0_u10_u2_n133 ) , .ZN( u0_u10_u2_n136 ) );
  AOI22_X1 u0_u10_u2_U43 (.ZN( u0_u10_u2_n135 ) , .B1( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n156 ) , .B2( u0_u10_u2_n180 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U44 (.ZN( u0_u10_u2_n149 ) , .B1( u0_u10_u2_n173 ) , .B2( u0_u10_u2_n188 ) , .A( u0_u10_u2_n95 ) );
  AND3_X1 u0_u10_u2_U45 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n95 ) );
  OAI21_X1 u0_u10_u2_U46 (.A( u0_u10_u2_n141 ) , .B2( u0_u10_u2_n142 ) , .ZN( u0_u10_u2_n146 ) , .B1( u0_u10_u2_n153 ) );
  OAI21_X1 u0_u10_u2_U47 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n141 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n177 ) );
  NOR3_X1 u0_u10_u2_U48 (.ZN( u0_u10_u2_n142 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n178 ) , .A1( u0_u10_u2_n181 ) );
  OAI21_X1 u0_u10_u2_U49 (.A( u0_u10_u2_n101 ) , .B2( u0_u10_u2_n121 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n164 ) );
  INV_X1 u0_u10_u2_U5 (.A( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n184 ) );
  NAND2_X1 u0_u10_u2_U50 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n155 ) );
  NAND2_X1 u0_u10_u2_U51 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n143 ) );
  NAND2_X1 u0_u10_u2_U52 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n152 ) );
  NAND2_X1 u0_u10_u2_U53 (.A1( u0_u10_u2_n100 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n132 ) );
  INV_X1 u0_u10_u2_U54 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U55 (.A( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n167 ) );
  NAND2_X1 u0_u10_u2_U56 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n113 ) );
  NAND2_X1 u0_u10_u2_U57 (.A1( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n131 ) );
  NAND2_X1 u0_u10_u2_U58 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n139 ) );
  NAND2_X1 u0_u10_u2_U59 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n133 ) );
  NOR4_X1 u0_u10_u2_U6 (.A4( u0_u10_u2_n124 ) , .A3( u0_u10_u2_n125 ) , .A2( u0_u10_u2_n126 ) , .A1( u0_u10_u2_n127 ) , .ZN( u0_u10_u2_n128 ) );
  NAND2_X1 u0_u10_u2_U60 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n103 ) , .ZN( u0_u10_u2_n154 ) );
  NAND2_X1 u0_u10_u2_U61 (.A2( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n104 ) , .ZN( u0_u10_u2_n119 ) );
  NAND2_X1 u0_u10_u2_U62 (.A2( u0_u10_u2_n107 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n123 ) );
  NAND2_X1 u0_u10_u2_U63 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n122 ) );
  INV_X1 u0_u10_u2_U64 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n172 ) );
  NAND2_X1 u0_u10_u2_U65 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n102 ) , .ZN( u0_u10_u2_n116 ) );
  NAND2_X1 u0_u10_u2_U66 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n120 ) );
  NAND2_X1 u0_u10_u2_U67 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n117 ) );
  INV_X1 u0_u10_u2_U68 (.ZN( u0_u10_u2_n187 ) , .A( u0_u10_u2_n99 ) );
  OAI21_X1 u0_u10_u2_U69 (.B1( u0_u10_u2_n137 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n98 ) , .ZN( u0_u10_u2_n99 ) );
  AOI21_X1 u0_u10_u2_U7 (.ZN( u0_u10_u2_n124 ) , .B1( u0_u10_u2_n131 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n172 ) );
  NOR2_X1 u0_u10_u2_U70 (.A2( u0_u10_X_16 ) , .ZN( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n166 ) );
  NOR2_X1 u0_u10_u2_U71 (.A2( u0_u10_X_13 ) , .A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n100 ) );
  NOR2_X1 u0_u10_u2_U72 (.A2( u0_u10_X_16 ) , .A1( u0_u10_X_17 ) , .ZN( u0_u10_u2_n138 ) );
  NOR2_X1 u0_u10_u2_U73 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n104 ) );
  NOR2_X1 u0_u10_u2_U74 (.A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n174 ) );
  NOR2_X1 u0_u10_u2_U75 (.A2( u0_u10_X_15 ) , .ZN( u0_u10_u2_n102 ) , .A1( u0_u10_u2_n165 ) );
  NOR2_X1 u0_u10_u2_U76 (.A2( u0_u10_X_17 ) , .ZN( u0_u10_u2_n114 ) , .A1( u0_u10_u2_n169 ) );
  AND2_X1 u0_u10_u2_U77 (.A1( u0_u10_X_15 ) , .ZN( u0_u10_u2_n105 ) , .A2( u0_u10_u2_n165 ) );
  AND2_X1 u0_u10_u2_U78 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n107 ) );
  AND2_X1 u0_u10_u2_U79 (.A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n174 ) );
  AOI21_X1 u0_u10_u2_U8 (.B2( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n127 ) , .A( u0_u10_u2_n137 ) , .B1( u0_u10_u2_n155 ) );
  AND2_X1 u0_u10_u2_U80 (.A1( u0_u10_X_13 ) , .A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n108 ) );
  INV_X1 u0_u10_u2_U81 (.A( u0_u10_X_16 ) , .ZN( u0_u10_u2_n169 ) );
  INV_X1 u0_u10_u2_U82 (.A( u0_u10_X_17 ) , .ZN( u0_u10_u2_n166 ) );
  INV_X1 u0_u10_u2_U83 (.A( u0_u10_X_13 ) , .ZN( u0_u10_u2_n174 ) );
  INV_X1 u0_u10_u2_U84 (.A( u0_u10_X_18 ) , .ZN( u0_u10_u2_n165 ) );
  NAND4_X1 u0_u10_u2_U85 (.ZN( u0_out10_30 ) , .A4( u0_u10_u2_n147 ) , .A3( u0_u10_u2_n148 ) , .A2( u0_u10_u2_n149 ) , .A1( u0_u10_u2_n187 ) );
  NOR3_X1 u0_u10_u2_U86 (.A3( u0_u10_u2_n144 ) , .A2( u0_u10_u2_n145 ) , .A1( u0_u10_u2_n146 ) , .ZN( u0_u10_u2_n147 ) );
  AOI21_X1 u0_u10_u2_U87 (.B2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n148 ) , .A( u0_u10_u2_n162 ) , .B1( u0_u10_u2_n182 ) );
  NAND4_X1 u0_u10_u2_U88 (.ZN( u0_out10_24 ) , .A4( u0_u10_u2_n111 ) , .A3( u0_u10_u2_n112 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n187 ) );
  AOI221_X1 u0_u10_u2_U89 (.A( u0_u10_u2_n109 ) , .B1( u0_u10_u2_n110 ) , .ZN( u0_u10_u2_n111 ) , .C1( u0_u10_u2_n134 ) , .C2( u0_u10_u2_n170 ) , .B2( u0_u10_u2_n173 ) );
  AOI21_X1 u0_u10_u2_U9 (.B2( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n125 ) , .A( u0_u10_u2_n171 ) , .B1( u0_u10_u2_n184 ) );
  AOI21_X1 u0_u10_u2_U90 (.ZN( u0_u10_u2_n112 ) , .B2( u0_u10_u2_n156 ) , .A( u0_u10_u2_n164 ) , .B1( u0_u10_u2_n181 ) );
  NAND4_X1 u0_u10_u2_U91 (.ZN( u0_out10_16 ) , .A4( u0_u10_u2_n128 ) , .A3( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n186 ) );
  AOI22_X1 u0_u10_u2_U92 (.A2( u0_u10_u2_n118 ) , .ZN( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n140 ) , .B1( u0_u10_u2_n157 ) , .B2( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U93 (.A( u0_u10_u2_n163 ) , .ZN( u0_u10_u2_n186 ) );
  OR4_X1 u0_u10_u2_U94 (.ZN( u0_out10_6 ) , .A4( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n162 ) , .A2( u0_u10_u2_n163 ) , .A1( u0_u10_u2_n164 ) );
  OR3_X1 u0_u10_u2_U95 (.A2( u0_u10_u2_n159 ) , .A1( u0_u10_u2_n160 ) , .ZN( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n183 ) );
  AOI21_X1 u0_u10_u2_U96 (.B2( u0_u10_u2_n154 ) , .B1( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n159 ) , .A( u0_u10_u2_n167 ) );
  NAND3_X1 u0_u10_u2_U97 (.A2( u0_u10_u2_n117 ) , .A1( u0_u10_u2_n122 ) , .A3( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n134 ) );
  NAND3_X1 u0_u10_u2_U98 (.ZN( u0_u10_u2_n110 ) , .A2( u0_u10_u2_n131 ) , .A3( u0_u10_u2_n139 ) , .A1( u0_u10_u2_n154 ) );
  NAND3_X1 u0_u10_u2_U99 (.A2( u0_u10_u2_n100 ) , .ZN( u0_u10_u2_n101 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n114 ) );
  OAI22_X1 u0_u10_u3_U10 (.B1( u0_u10_u3_n113 ) , .A2( u0_u10_u3_n135 ) , .A1( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n164 ) , .ZN( u0_u10_u3_n98 ) );
  OAI211_X1 u0_u10_u3_U11 (.B( u0_u10_u3_n106 ) , .ZN( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n128 ) , .C1( u0_u10_u3_n167 ) , .A( u0_u10_u3_n181 ) );
  AOI221_X1 u0_u10_u3_U12 (.C1( u0_u10_u3_n105 ) , .ZN( u0_u10_u3_n106 ) , .A( u0_u10_u3_n131 ) , .B2( u0_u10_u3_n132 ) , .C2( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n169 ) );
  INV_X1 u0_u10_u3_U13 (.ZN( u0_u10_u3_n181 ) , .A( u0_u10_u3_n98 ) );
  NAND2_X1 u0_u10_u3_U14 (.ZN( u0_u10_u3_n105 ) , .A2( u0_u10_u3_n130 ) , .A1( u0_u10_u3_n155 ) );
  AOI22_X1 u0_u10_u3_U15 (.B1( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n116 ) , .ZN( u0_u10_u3_n123 ) , .B2( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U16 (.ZN( u0_u10_u3_n116 ) , .A2( u0_u10_u3_n151 ) , .A1( u0_u10_u3_n182 ) );
  NOR2_X1 u0_u10_u3_U17 (.ZN( u0_u10_u3_n126 ) , .A2( u0_u10_u3_n150 ) , .A1( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U18 (.ZN( u0_u10_u3_n112 ) , .B2( u0_u10_u3_n146 ) , .B1( u0_u10_u3_n155 ) , .A( u0_u10_u3_n167 ) );
  NAND2_X1 u0_u10_u3_U19 (.A1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n142 ) , .A2( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U20 (.ZN( u0_u10_u3_n132 ) , .A2( u0_u10_u3_n152 ) , .A1( u0_u10_u3_n156 ) );
  AND2_X1 u0_u10_u3_U21 (.A2( u0_u10_u3_n113 ) , .A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n151 ) );
  INV_X1 u0_u10_u3_U22 (.A( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n165 ) );
  INV_X1 u0_u10_u3_U23 (.A( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n170 ) );
  NAND2_X1 u0_u10_u3_U24 (.A1( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .ZN( u0_u10_u3_n140 ) );
  NAND2_X1 u0_u10_u3_U25 (.ZN( u0_u10_u3_n117 ) , .A1( u0_u10_u3_n124 ) , .A2( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U26 (.ZN( u0_u10_u3_n143 ) , .A1( u0_u10_u3_n165 ) , .A2( u0_u10_u3_n167 ) );
  INV_X1 u0_u10_u3_U27 (.A( u0_u10_u3_n130 ) , .ZN( u0_u10_u3_n177 ) );
  INV_X1 u0_u10_u3_U28 (.A( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n176 ) );
  INV_X1 u0_u10_u3_U29 (.A( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n174 ) );
  INV_X1 u0_u10_u3_U3 (.A( u0_u10_u3_n129 ) , .ZN( u0_u10_u3_n183 ) );
  INV_X1 u0_u10_u3_U30 (.A( u0_u10_u3_n139 ) , .ZN( u0_u10_u3_n185 ) );
  NOR2_X1 u0_u10_u3_U31 (.ZN( u0_u10_u3_n135 ) , .A2( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n169 ) );
  OAI222_X1 u0_u10_u3_U32 (.C2( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .B1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n138 ) , .B2( u0_u10_u3_n146 ) , .C1( u0_u10_u3_n154 ) , .A1( u0_u10_u3_n164 ) );
  NOR4_X1 u0_u10_u3_U33 (.A4( u0_u10_u3_n157 ) , .A3( u0_u10_u3_n158 ) , .A2( u0_u10_u3_n159 ) , .A1( u0_u10_u3_n160 ) , .ZN( u0_u10_u3_n161 ) );
  AOI21_X1 u0_u10_u3_U34 (.B2( u0_u10_u3_n152 ) , .B1( u0_u10_u3_n153 ) , .ZN( u0_u10_u3_n158 ) , .A( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U35 (.A( u0_u10_u3_n154 ) , .B2( u0_u10_u3_n155 ) , .B1( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n157 ) );
  AOI21_X1 u0_u10_u3_U36 (.A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n150 ) , .B1( u0_u10_u3_n151 ) , .ZN( u0_u10_u3_n159 ) );
  AOI211_X1 u0_u10_u3_U37 (.ZN( u0_u10_u3_n109 ) , .A( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n129 ) , .B( u0_u10_u3_n138 ) , .C1( u0_u10_u3_n141 ) );
  AOI211_X1 u0_u10_u3_U38 (.B( u0_u10_u3_n119 ) , .A( u0_u10_u3_n120 ) , .C2( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n122 ) , .C1( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U39 (.A( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U4 (.A( u0_u10_u3_n140 ) , .ZN( u0_u10_u3_n182 ) );
  OAI22_X1 u0_u10_u3_U40 (.B1( u0_u10_u3_n118 ) , .ZN( u0_u10_u3_n120 ) , .A1( u0_u10_u3_n135 ) , .B2( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n178 ) );
  AND3_X1 u0_u10_u3_U41 (.ZN( u0_u10_u3_n118 ) , .A2( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n144 ) , .A3( u0_u10_u3_n152 ) );
  INV_X1 u0_u10_u3_U42 (.A( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U43 (.ZN( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n164 ) );
  OAI211_X1 u0_u10_u3_U44 (.B( u0_u10_u3_n127 ) , .ZN( u0_u10_u3_n139 ) , .C1( u0_u10_u3_n150 ) , .C2( u0_u10_u3_n154 ) , .A( u0_u10_u3_n184 ) );
  INV_X1 u0_u10_u3_U45 (.A( u0_u10_u3_n125 ) , .ZN( u0_u10_u3_n184 ) );
  AOI221_X1 u0_u10_u3_U46 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n127 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n169 ) , .B2( u0_u10_u3_n170 ) , .B1( u0_u10_u3_n174 ) );
  OAI22_X1 u0_u10_u3_U47 (.A1( u0_u10_u3_n124 ) , .ZN( u0_u10_u3_n125 ) , .B2( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n165 ) , .B1( u0_u10_u3_n167 ) );
  NOR2_X1 u0_u10_u3_U48 (.A1( u0_u10_u3_n113 ) , .ZN( u0_u10_u3_n131 ) , .A2( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U49 (.A1( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n150 ) , .A2( u0_u10_u3_n99 ) );
  INV_X1 u0_u10_u3_U5 (.A( u0_u10_u3_n117 ) , .ZN( u0_u10_u3_n178 ) );
  NAND2_X1 u0_u10_u3_U50 (.A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n155 ) , .A1( u0_u10_u3_n97 ) );
  INV_X1 u0_u10_u3_U51 (.A( u0_u10_u3_n141 ) , .ZN( u0_u10_u3_n167 ) );
  AOI21_X1 u0_u10_u3_U52 (.B2( u0_u10_u3_n114 ) , .B1( u0_u10_u3_n146 ) , .A( u0_u10_u3_n154 ) , .ZN( u0_u10_u3_n94 ) );
  AOI21_X1 u0_u10_u3_U53 (.ZN( u0_u10_u3_n110 ) , .B2( u0_u10_u3_n142 ) , .B1( u0_u10_u3_n186 ) , .A( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U54 (.A( u0_u10_u3_n145 ) , .ZN( u0_u10_u3_n186 ) );
  AOI21_X1 u0_u10_u3_U55 (.B1( u0_u10_u3_n124 ) , .A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U56 (.A( u0_u10_u3_n149 ) , .ZN( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U57 (.ZN( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n96 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U58 (.A2( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n146 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U59 (.A1( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n99 ) );
  AOI221_X1 u0_u10_u3_U6 (.A( u0_u10_u3_n131 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n134 ) , .B1( u0_u10_u3_n143 ) , .B2( u0_u10_u3_n177 ) );
  NAND2_X1 u0_u10_u3_U60 (.A1( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n156 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U61 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U62 (.A1( u0_u10_u3_n100 ) , .A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n128 ) );
  NAND2_X1 u0_u10_u3_U63 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n152 ) );
  NAND2_X1 u0_u10_u3_U64 (.A2( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n114 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U65 (.ZN( u0_u10_u3_n107 ) , .A1( u0_u10_u3_n97 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U66 (.A2( u0_u10_u3_n100 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n113 ) );
  NAND2_X1 u0_u10_u3_U67 (.A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n153 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U68 (.A2( u0_u10_u3_n103 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n130 ) );
  NAND2_X1 u0_u10_u3_U69 (.A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n96 ) );
  OAI22_X1 u0_u10_u3_U7 (.B2( u0_u10_u3_n147 ) , .A2( u0_u10_u3_n148 ) , .ZN( u0_u10_u3_n160 ) , .B1( u0_u10_u3_n165 ) , .A1( u0_u10_u3_n168 ) );
  NAND2_X1 u0_u10_u3_U70 (.A1( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n108 ) );
  NOR2_X1 u0_u10_u3_U71 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n99 ) );
  NOR2_X1 u0_u10_u3_U72 (.A2( u0_u10_X_21 ) , .A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n103 ) );
  NOR2_X1 u0_u10_u3_U73 (.A2( u0_u10_X_24 ) , .A1( u0_u10_u3_n171 ) , .ZN( u0_u10_u3_n97 ) );
  NOR2_X1 u0_u10_u3_U74 (.A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U75 (.A2( u0_u10_X_19 ) , .A1( u0_u10_u3_n172 ) , .ZN( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U76 (.A1( u0_u10_X_22 ) , .A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U77 (.A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n149 ) , .A2( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U78 (.A2( u0_u10_X_22 ) , .A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n121 ) );
  AND2_X1 u0_u10_u3_U79 (.A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n101 ) , .A2( u0_u10_u3_n171 ) );
  AND3_X1 u0_u10_u3_U8 (.A3( u0_u10_u3_n144 ) , .A2( u0_u10_u3_n145 ) , .A1( u0_u10_u3_n146 ) , .ZN( u0_u10_u3_n147 ) );
  AND2_X1 u0_u10_u3_U80 (.A1( u0_u10_X_19 ) , .ZN( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n172 ) );
  AND2_X1 u0_u10_u3_U81 (.A1( u0_u10_X_21 ) , .A2( u0_u10_X_24 ) , .ZN( u0_u10_u3_n100 ) );
  AND2_X1 u0_u10_u3_U82 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n104 ) );
  INV_X1 u0_u10_u3_U83 (.A( u0_u10_X_22 ) , .ZN( u0_u10_u3_n166 ) );
  INV_X1 u0_u10_u3_U84 (.A( u0_u10_X_21 ) , .ZN( u0_u10_u3_n171 ) );
  INV_X1 u0_u10_u3_U85 (.A( u0_u10_X_20 ) , .ZN( u0_u10_u3_n172 ) );
  OR4_X1 u0_u10_u3_U86 (.ZN( u0_out10_10 ) , .A4( u0_u10_u3_n136 ) , .A3( u0_u10_u3_n137 ) , .A1( u0_u10_u3_n138 ) , .A2( u0_u10_u3_n139 ) );
  OAI222_X1 u0_u10_u3_U87 (.C1( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n137 ) , .B1( u0_u10_u3_n148 ) , .A2( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n154 ) , .C2( u0_u10_u3_n164 ) , .A1( u0_u10_u3_n167 ) );
  OAI221_X1 u0_u10_u3_U88 (.A( u0_u10_u3_n134 ) , .B2( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n136 ) , .C1( u0_u10_u3_n149 ) , .B1( u0_u10_u3_n151 ) , .C2( u0_u10_u3_n183 ) );
  NAND4_X1 u0_u10_u3_U89 (.ZN( u0_out10_26 ) , .A4( u0_u10_u3_n109 ) , .A3( u0_u10_u3_n110 ) , .A2( u0_u10_u3_n111 ) , .A1( u0_u10_u3_n173 ) );
  INV_X1 u0_u10_u3_U9 (.A( u0_u10_u3_n143 ) , .ZN( u0_u10_u3_n168 ) );
  INV_X1 u0_u10_u3_U90 (.ZN( u0_u10_u3_n173 ) , .A( u0_u10_u3_n94 ) );
  OAI21_X1 u0_u10_u3_U91 (.ZN( u0_u10_u3_n111 ) , .B2( u0_u10_u3_n117 ) , .A( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n176 ) );
  NAND4_X1 u0_u10_u3_U92 (.ZN( u0_out10_20 ) , .A4( u0_u10_u3_n122 ) , .A3( u0_u10_u3_n123 ) , .A1( u0_u10_u3_n175 ) , .A2( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U93 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U94 (.A( u0_u10_u3_n112 ) , .ZN( u0_u10_u3_n175 ) );
  NAND4_X1 u0_u10_u3_U95 (.ZN( u0_out10_1 ) , .A4( u0_u10_u3_n161 ) , .A3( u0_u10_u3_n162 ) , .A2( u0_u10_u3_n163 ) , .A1( u0_u10_u3_n185 ) );
  NAND2_X1 u0_u10_u3_U96 (.ZN( u0_u10_u3_n163 ) , .A2( u0_u10_u3_n170 ) , .A1( u0_u10_u3_n176 ) );
  AOI22_X1 u0_u10_u3_U97 (.B2( u0_u10_u3_n140 ) , .B1( u0_u10_u3_n141 ) , .A2( u0_u10_u3_n142 ) , .ZN( u0_u10_u3_n162 ) , .A1( u0_u10_u3_n177 ) );
  NAND3_X1 u0_u10_u3_U98 (.A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n145 ) , .A3( u0_u10_u3_n153 ) );
  NAND3_X1 u0_u10_u3_U99 (.ZN( u0_u10_u3_n129 ) , .A2( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n153 ) , .A3( u0_u10_u3_n182 ) );
  XOR2_X1 u0_u11_U13 (.B( u0_K12_42 ) , .A( u0_R10_29 ) , .Z( u0_u11_X_42 ) );
  XOR2_X1 u0_u11_U14 (.B( u0_K12_41 ) , .A( u0_R10_28 ) , .Z( u0_u11_X_41 ) );
  XOR2_X1 u0_u11_U18 (.B( u0_K12_38 ) , .A( u0_R10_25 ) , .Z( u0_u11_X_38 ) );
  XOR2_X1 u0_u11_U19 (.B( u0_K12_37 ) , .A( u0_R10_24 ) , .Z( u0_u11_X_37 ) );
  XOR2_X1 u0_u11_U20 (.B( u0_K12_36 ) , .A( u0_R10_25 ) , .Z( u0_u11_X_36 ) );
  XOR2_X1 u0_u11_U21 (.B( u0_K12_35 ) , .A( u0_R10_24 ) , .Z( u0_u11_X_35 ) );
  XOR2_X1 u0_u11_U24 (.B( u0_K12_32 ) , .A( u0_R10_21 ) , .Z( u0_u11_X_32 ) );
  XOR2_X1 u0_u11_U25 (.B( u0_K12_31 ) , .A( u0_R10_20 ) , .Z( u0_u11_X_31 ) );
  XOR2_X1 u0_u11_U33 (.B( u0_K12_24 ) , .A( u0_R10_17 ) , .Z( u0_u11_X_24 ) );
  XOR2_X1 u0_u11_U34 (.B( u0_K12_23 ) , .A( u0_R10_16 ) , .Z( u0_u11_X_23 ) );
  XOR2_X1 u0_u11_U36 (.B( u0_K12_21 ) , .A( u0_R10_14 ) , .Z( u0_u11_X_21 ) );
  XOR2_X1 u0_u11_U39 (.B( u0_K12_19 ) , .A( u0_R10_12 ) , .Z( u0_u11_X_19 ) );
  XOR2_X1 u0_u11_U41 (.B( u0_K12_17 ) , .A( u0_R10_12 ) , .Z( u0_u11_X_17 ) );
  OAI22_X1 u0_u11_u2_U10 (.ZN( u0_u11_u2_n109 ) , .A2( u0_u11_u2_n113 ) , .B2( u0_u11_u2_n133 ) , .B1( u0_u11_u2_n167 ) , .A1( u0_u11_u2_n168 ) );
  NAND3_X1 u0_u11_u2_U100 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n98 ) );
  OAI22_X1 u0_u11_u2_U11 (.B1( u0_u11_u2_n151 ) , .A2( u0_u11_u2_n152 ) , .A1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n160 ) , .B2( u0_u11_u2_n168 ) );
  NOR3_X1 u0_u11_u2_U12 (.A1( u0_u11_u2_n150 ) , .ZN( u0_u11_u2_n151 ) , .A3( u0_u11_u2_n175 ) , .A2( u0_u11_u2_n188 ) );
  AOI21_X1 u0_u11_u2_U13 (.ZN( u0_u11_u2_n144 ) , .B2( u0_u11_u2_n155 ) , .A( u0_u11_u2_n172 ) , .B1( u0_u11_u2_n185 ) );
  AOI21_X1 u0_u11_u2_U14 (.B2( u0_u11_u2_n143 ) , .ZN( u0_u11_u2_n145 ) , .B1( u0_u11_u2_n152 ) , .A( u0_u11_u2_n171 ) );
  AOI21_X1 u0_u11_u2_U15 (.B2( u0_u11_u2_n120 ) , .B1( u0_u11_u2_n121 ) , .ZN( u0_u11_u2_n126 ) , .A( u0_u11_u2_n167 ) );
  INV_X1 u0_u11_u2_U16 (.A( u0_u11_u2_n156 ) , .ZN( u0_u11_u2_n171 ) );
  INV_X1 u0_u11_u2_U17 (.A( u0_u11_u2_n120 ) , .ZN( u0_u11_u2_n188 ) );
  NAND2_X1 u0_u11_u2_U18 (.A2( u0_u11_u2_n122 ) , .ZN( u0_u11_u2_n150 ) , .A1( u0_u11_u2_n152 ) );
  INV_X1 u0_u11_u2_U19 (.A( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n170 ) );
  INV_X1 u0_u11_u2_U20 (.A( u0_u11_u2_n137 ) , .ZN( u0_u11_u2_n173 ) );
  NAND2_X1 u0_u11_u2_U21 (.A1( u0_u11_u2_n132 ) , .A2( u0_u11_u2_n139 ) , .ZN( u0_u11_u2_n157 ) );
  INV_X1 u0_u11_u2_U22 (.A( u0_u11_u2_n113 ) , .ZN( u0_u11_u2_n178 ) );
  INV_X1 u0_u11_u2_U23 (.A( u0_u11_u2_n139 ) , .ZN( u0_u11_u2_n175 ) );
  INV_X1 u0_u11_u2_U24 (.A( u0_u11_u2_n155 ) , .ZN( u0_u11_u2_n181 ) );
  INV_X1 u0_u11_u2_U25 (.A( u0_u11_u2_n119 ) , .ZN( u0_u11_u2_n177 ) );
  INV_X1 u0_u11_u2_U26 (.A( u0_u11_u2_n116 ) , .ZN( u0_u11_u2_n180 ) );
  INV_X1 u0_u11_u2_U27 (.A( u0_u11_u2_n131 ) , .ZN( u0_u11_u2_n179 ) );
  INV_X1 u0_u11_u2_U28 (.A( u0_u11_u2_n154 ) , .ZN( u0_u11_u2_n176 ) );
  NAND2_X1 u0_u11_u2_U29 (.A2( u0_u11_u2_n116 ) , .A1( u0_u11_u2_n117 ) , .ZN( u0_u11_u2_n118 ) );
  NOR2_X1 u0_u11_u2_U3 (.ZN( u0_u11_u2_n121 ) , .A2( u0_u11_u2_n177 ) , .A1( u0_u11_u2_n180 ) );
  INV_X1 u0_u11_u2_U30 (.A( u0_u11_u2_n132 ) , .ZN( u0_u11_u2_n182 ) );
  INV_X1 u0_u11_u2_U31 (.A( u0_u11_u2_n158 ) , .ZN( u0_u11_u2_n183 ) );
  OAI21_X1 u0_u11_u2_U32 (.A( u0_u11_u2_n156 ) , .B1( u0_u11_u2_n157 ) , .ZN( u0_u11_u2_n158 ) , .B2( u0_u11_u2_n179 ) );
  NOR2_X1 u0_u11_u2_U33 (.ZN( u0_u11_u2_n156 ) , .A1( u0_u11_u2_n166 ) , .A2( u0_u11_u2_n169 ) );
  NOR2_X1 u0_u11_u2_U34 (.A2( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n137 ) , .A1( u0_u11_u2_n140 ) );
  NOR2_X1 u0_u11_u2_U35 (.A2( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n153 ) , .A1( u0_u11_u2_n156 ) );
  AOI211_X1 u0_u11_u2_U36 (.ZN( u0_u11_u2_n130 ) , .C1( u0_u11_u2_n138 ) , .C2( u0_u11_u2_n179 ) , .B( u0_u11_u2_n96 ) , .A( u0_u11_u2_n97 ) );
  OAI22_X1 u0_u11_u2_U37 (.B1( u0_u11_u2_n133 ) , .A2( u0_u11_u2_n137 ) , .A1( u0_u11_u2_n152 ) , .B2( u0_u11_u2_n168 ) , .ZN( u0_u11_u2_n97 ) );
  OAI221_X1 u0_u11_u2_U38 (.B1( u0_u11_u2_n113 ) , .C1( u0_u11_u2_n132 ) , .A( u0_u11_u2_n149 ) , .B2( u0_u11_u2_n171 ) , .C2( u0_u11_u2_n172 ) , .ZN( u0_u11_u2_n96 ) );
  OAI221_X1 u0_u11_u2_U39 (.A( u0_u11_u2_n115 ) , .C2( u0_u11_u2_n123 ) , .B2( u0_u11_u2_n143 ) , .B1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n163 ) , .C1( u0_u11_u2_n168 ) );
  INV_X1 u0_u11_u2_U4 (.A( u0_u11_u2_n134 ) , .ZN( u0_u11_u2_n185 ) );
  OAI21_X1 u0_u11_u2_U40 (.A( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n115 ) , .B1( u0_u11_u2_n176 ) , .B2( u0_u11_u2_n178 ) );
  OAI221_X1 u0_u11_u2_U41 (.A( u0_u11_u2_n135 ) , .B2( u0_u11_u2_n136 ) , .B1( u0_u11_u2_n137 ) , .ZN( u0_u11_u2_n162 ) , .C2( u0_u11_u2_n167 ) , .C1( u0_u11_u2_n185 ) );
  AND3_X1 u0_u11_u2_U42 (.A3( u0_u11_u2_n131 ) , .A2( u0_u11_u2_n132 ) , .A1( u0_u11_u2_n133 ) , .ZN( u0_u11_u2_n136 ) );
  AOI22_X1 u0_u11_u2_U43 (.ZN( u0_u11_u2_n135 ) , .B1( u0_u11_u2_n140 ) , .A1( u0_u11_u2_n156 ) , .B2( u0_u11_u2_n180 ) , .A2( u0_u11_u2_n188 ) );
  AOI21_X1 u0_u11_u2_U44 (.ZN( u0_u11_u2_n149 ) , .B1( u0_u11_u2_n173 ) , .B2( u0_u11_u2_n188 ) , .A( u0_u11_u2_n95 ) );
  AND3_X1 u0_u11_u2_U45 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n156 ) , .ZN( u0_u11_u2_n95 ) );
  OAI21_X1 u0_u11_u2_U46 (.A( u0_u11_u2_n101 ) , .B2( u0_u11_u2_n121 ) , .B1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n164 ) );
  NAND2_X1 u0_u11_u2_U47 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n155 ) );
  NAND2_X1 u0_u11_u2_U48 (.A2( u0_u11_u2_n105 ) , .A1( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n143 ) );
  NAND2_X1 u0_u11_u2_U49 (.A1( u0_u11_u2_n104 ) , .A2( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n152 ) );
  INV_X1 u0_u11_u2_U5 (.A( u0_u11_u2_n150 ) , .ZN( u0_u11_u2_n184 ) );
  NAND2_X1 u0_u11_u2_U50 (.A1( u0_u11_u2_n100 ) , .A2( u0_u11_u2_n105 ) , .ZN( u0_u11_u2_n132 ) );
  INV_X1 u0_u11_u2_U51 (.A( u0_u11_u2_n140 ) , .ZN( u0_u11_u2_n168 ) );
  INV_X1 u0_u11_u2_U52 (.A( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n167 ) );
  OAI21_X1 u0_u11_u2_U53 (.A( u0_u11_u2_n141 ) , .B2( u0_u11_u2_n142 ) , .ZN( u0_u11_u2_n146 ) , .B1( u0_u11_u2_n153 ) );
  OAI21_X1 u0_u11_u2_U54 (.A( u0_u11_u2_n140 ) , .ZN( u0_u11_u2_n141 ) , .B1( u0_u11_u2_n176 ) , .B2( u0_u11_u2_n177 ) );
  NOR3_X1 u0_u11_u2_U55 (.ZN( u0_u11_u2_n142 ) , .A3( u0_u11_u2_n175 ) , .A2( u0_u11_u2_n178 ) , .A1( u0_u11_u2_n181 ) );
  NAND2_X1 u0_u11_u2_U56 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n113 ) );
  NAND2_X1 u0_u11_u2_U57 (.A1( u0_u11_u2_n106 ) , .A2( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n131 ) );
  NAND2_X1 u0_u11_u2_U58 (.A1( u0_u11_u2_n103 ) , .A2( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n139 ) );
  NAND2_X1 u0_u11_u2_U59 (.A1( u0_u11_u2_n103 ) , .A2( u0_u11_u2_n105 ) , .ZN( u0_u11_u2_n133 ) );
  NOR4_X1 u0_u11_u2_U6 (.A4( u0_u11_u2_n124 ) , .A3( u0_u11_u2_n125 ) , .A2( u0_u11_u2_n126 ) , .A1( u0_u11_u2_n127 ) , .ZN( u0_u11_u2_n128 ) );
  NAND2_X1 u0_u11_u2_U60 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n103 ) , .ZN( u0_u11_u2_n154 ) );
  NAND2_X1 u0_u11_u2_U61 (.A2( u0_u11_u2_n103 ) , .A1( u0_u11_u2_n104 ) , .ZN( u0_u11_u2_n119 ) );
  NAND2_X1 u0_u11_u2_U62 (.A2( u0_u11_u2_n107 ) , .A1( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n123 ) );
  NAND2_X1 u0_u11_u2_U63 (.A1( u0_u11_u2_n104 ) , .A2( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n122 ) );
  INV_X1 u0_u11_u2_U64 (.A( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n172 ) );
  NAND2_X1 u0_u11_u2_U65 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n102 ) , .ZN( u0_u11_u2_n116 ) );
  NAND2_X1 u0_u11_u2_U66 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n120 ) );
  NAND2_X1 u0_u11_u2_U67 (.A2( u0_u11_u2_n105 ) , .A1( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n117 ) );
  INV_X1 u0_u11_u2_U68 (.ZN( u0_u11_u2_n187 ) , .A( u0_u11_u2_n99 ) );
  OAI21_X1 u0_u11_u2_U69 (.B1( u0_u11_u2_n137 ) , .B2( u0_u11_u2_n143 ) , .A( u0_u11_u2_n98 ) , .ZN( u0_u11_u2_n99 ) );
  AOI21_X1 u0_u11_u2_U7 (.ZN( u0_u11_u2_n124 ) , .B1( u0_u11_u2_n131 ) , .B2( u0_u11_u2_n143 ) , .A( u0_u11_u2_n172 ) );
  NOR2_X1 u0_u11_u2_U70 (.A2( u0_u11_X_16 ) , .ZN( u0_u11_u2_n140 ) , .A1( u0_u11_u2_n166 ) );
  NOR2_X1 u0_u11_u2_U71 (.A2( u0_u11_X_13 ) , .A1( u0_u11_X_14 ) , .ZN( u0_u11_u2_n100 ) );
  NOR2_X1 u0_u11_u2_U72 (.A2( u0_u11_X_16 ) , .A1( u0_u11_X_17 ) , .ZN( u0_u11_u2_n138 ) );
  NOR2_X1 u0_u11_u2_U73 (.A2( u0_u11_X_15 ) , .A1( u0_u11_X_18 ) , .ZN( u0_u11_u2_n104 ) );
  NOR2_X1 u0_u11_u2_U74 (.A2( u0_u11_X_14 ) , .ZN( u0_u11_u2_n103 ) , .A1( u0_u11_u2_n174 ) );
  NOR2_X1 u0_u11_u2_U75 (.A2( u0_u11_X_15 ) , .ZN( u0_u11_u2_n102 ) , .A1( u0_u11_u2_n165 ) );
  NOR2_X1 u0_u11_u2_U76 (.A2( u0_u11_X_17 ) , .ZN( u0_u11_u2_n114 ) , .A1( u0_u11_u2_n169 ) );
  AND2_X1 u0_u11_u2_U77 (.A1( u0_u11_X_15 ) , .ZN( u0_u11_u2_n105 ) , .A2( u0_u11_u2_n165 ) );
  AND2_X1 u0_u11_u2_U78 (.A2( u0_u11_X_15 ) , .A1( u0_u11_X_18 ) , .ZN( u0_u11_u2_n107 ) );
  AND2_X1 u0_u11_u2_U79 (.A1( u0_u11_X_14 ) , .ZN( u0_u11_u2_n106 ) , .A2( u0_u11_u2_n174 ) );
  AOI21_X1 u0_u11_u2_U8 (.B2( u0_u11_u2_n119 ) , .ZN( u0_u11_u2_n127 ) , .A( u0_u11_u2_n137 ) , .B1( u0_u11_u2_n155 ) );
  AND2_X1 u0_u11_u2_U80 (.A1( u0_u11_X_13 ) , .A2( u0_u11_X_14 ) , .ZN( u0_u11_u2_n108 ) );
  INV_X1 u0_u11_u2_U81 (.A( u0_u11_X_16 ) , .ZN( u0_u11_u2_n169 ) );
  INV_X1 u0_u11_u2_U82 (.A( u0_u11_X_17 ) , .ZN( u0_u11_u2_n166 ) );
  INV_X1 u0_u11_u2_U83 (.A( u0_u11_X_13 ) , .ZN( u0_u11_u2_n174 ) );
  INV_X1 u0_u11_u2_U84 (.A( u0_u11_X_18 ) , .ZN( u0_u11_u2_n165 ) );
  NAND4_X1 u0_u11_u2_U85 (.ZN( u0_out11_30 ) , .A4( u0_u11_u2_n147 ) , .A3( u0_u11_u2_n148 ) , .A2( u0_u11_u2_n149 ) , .A1( u0_u11_u2_n187 ) );
  NOR3_X1 u0_u11_u2_U86 (.A3( u0_u11_u2_n144 ) , .A2( u0_u11_u2_n145 ) , .A1( u0_u11_u2_n146 ) , .ZN( u0_u11_u2_n147 ) );
  AOI21_X1 u0_u11_u2_U87 (.B2( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n148 ) , .A( u0_u11_u2_n162 ) , .B1( u0_u11_u2_n182 ) );
  NAND4_X1 u0_u11_u2_U88 (.ZN( u0_out11_24 ) , .A4( u0_u11_u2_n111 ) , .A3( u0_u11_u2_n112 ) , .A1( u0_u11_u2_n130 ) , .A2( u0_u11_u2_n187 ) );
  AOI221_X1 u0_u11_u2_U89 (.A( u0_u11_u2_n109 ) , .B1( u0_u11_u2_n110 ) , .ZN( u0_u11_u2_n111 ) , .C1( u0_u11_u2_n134 ) , .C2( u0_u11_u2_n170 ) , .B2( u0_u11_u2_n173 ) );
  AOI21_X1 u0_u11_u2_U9 (.B2( u0_u11_u2_n123 ) , .ZN( u0_u11_u2_n125 ) , .A( u0_u11_u2_n171 ) , .B1( u0_u11_u2_n184 ) );
  AOI21_X1 u0_u11_u2_U90 (.ZN( u0_u11_u2_n112 ) , .B2( u0_u11_u2_n156 ) , .A( u0_u11_u2_n164 ) , .B1( u0_u11_u2_n181 ) );
  NAND4_X1 u0_u11_u2_U91 (.ZN( u0_out11_16 ) , .A4( u0_u11_u2_n128 ) , .A3( u0_u11_u2_n129 ) , .A1( u0_u11_u2_n130 ) , .A2( u0_u11_u2_n186 ) );
  AOI22_X1 u0_u11_u2_U92 (.A2( u0_u11_u2_n118 ) , .ZN( u0_u11_u2_n129 ) , .A1( u0_u11_u2_n140 ) , .B1( u0_u11_u2_n157 ) , .B2( u0_u11_u2_n170 ) );
  INV_X1 u0_u11_u2_U93 (.A( u0_u11_u2_n163 ) , .ZN( u0_u11_u2_n186 ) );
  OR4_X1 u0_u11_u2_U94 (.ZN( u0_out11_6 ) , .A4( u0_u11_u2_n161 ) , .A3( u0_u11_u2_n162 ) , .A2( u0_u11_u2_n163 ) , .A1( u0_u11_u2_n164 ) );
  OR3_X1 u0_u11_u2_U95 (.A2( u0_u11_u2_n159 ) , .A1( u0_u11_u2_n160 ) , .ZN( u0_u11_u2_n161 ) , .A3( u0_u11_u2_n183 ) );
  AOI21_X1 u0_u11_u2_U96 (.B2( u0_u11_u2_n154 ) , .B1( u0_u11_u2_n155 ) , .ZN( u0_u11_u2_n159 ) , .A( u0_u11_u2_n167 ) );
  NAND3_X1 u0_u11_u2_U97 (.A2( u0_u11_u2_n117 ) , .A1( u0_u11_u2_n122 ) , .A3( u0_u11_u2_n123 ) , .ZN( u0_u11_u2_n134 ) );
  NAND3_X1 u0_u11_u2_U98 (.ZN( u0_u11_u2_n110 ) , .A2( u0_u11_u2_n131 ) , .A3( u0_u11_u2_n139 ) , .A1( u0_u11_u2_n154 ) );
  NAND3_X1 u0_u11_u2_U99 (.A2( u0_u11_u2_n100 ) , .ZN( u0_u11_u2_n101 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n114 ) );
  OAI211_X1 u0_u11_u3_U10 (.B( u0_u11_u3_n106 ) , .ZN( u0_u11_u3_n119 ) , .C2( u0_u11_u3_n128 ) , .C1( u0_u11_u3_n167 ) , .A( u0_u11_u3_n181 ) );
  INV_X1 u0_u11_u3_U11 (.ZN( u0_u11_u3_n181 ) , .A( u0_u11_u3_n98 ) );
  AOI221_X1 u0_u11_u3_U12 (.C1( u0_u11_u3_n105 ) , .ZN( u0_u11_u3_n106 ) , .A( u0_u11_u3_n131 ) , .B2( u0_u11_u3_n132 ) , .C2( u0_u11_u3_n133 ) , .B1( u0_u11_u3_n169 ) );
  OAI22_X1 u0_u11_u3_U13 (.B1( u0_u11_u3_n113 ) , .A2( u0_u11_u3_n135 ) , .A1( u0_u11_u3_n150 ) , .B2( u0_u11_u3_n164 ) , .ZN( u0_u11_u3_n98 ) );
  AOI22_X1 u0_u11_u3_U14 (.B1( u0_u11_u3_n115 ) , .A2( u0_u11_u3_n116 ) , .ZN( u0_u11_u3_n123 ) , .B2( u0_u11_u3_n133 ) , .A1( u0_u11_u3_n169 ) );
  NAND2_X1 u0_u11_u3_U15 (.ZN( u0_u11_u3_n116 ) , .A2( u0_u11_u3_n151 ) , .A1( u0_u11_u3_n182 ) );
  NOR2_X1 u0_u11_u3_U16 (.ZN( u0_u11_u3_n126 ) , .A2( u0_u11_u3_n150 ) , .A1( u0_u11_u3_n164 ) );
  AOI21_X1 u0_u11_u3_U17 (.ZN( u0_u11_u3_n112 ) , .B2( u0_u11_u3_n146 ) , .B1( u0_u11_u3_n155 ) , .A( u0_u11_u3_n167 ) );
  NAND2_X1 u0_u11_u3_U18 (.A1( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n142 ) , .A2( u0_u11_u3_n164 ) );
  NAND2_X1 u0_u11_u3_U19 (.ZN( u0_u11_u3_n132 ) , .A2( u0_u11_u3_n152 ) , .A1( u0_u11_u3_n156 ) );
  INV_X1 u0_u11_u3_U20 (.A( u0_u11_u3_n133 ) , .ZN( u0_u11_u3_n165 ) );
  NAND2_X1 u0_u11_u3_U21 (.ZN( u0_u11_u3_n143 ) , .A1( u0_u11_u3_n165 ) , .A2( u0_u11_u3_n167 ) );
  AND2_X1 u0_u11_u3_U22 (.A2( u0_u11_u3_n113 ) , .A1( u0_u11_u3_n114 ) , .ZN( u0_u11_u3_n151 ) );
  INV_X1 u0_u11_u3_U23 (.A( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n170 ) );
  NAND2_X1 u0_u11_u3_U24 (.A1( u0_u11_u3_n107 ) , .A2( u0_u11_u3_n108 ) , .ZN( u0_u11_u3_n140 ) );
  NAND2_X1 u0_u11_u3_U25 (.ZN( u0_u11_u3_n117 ) , .A1( u0_u11_u3_n124 ) , .A2( u0_u11_u3_n148 ) );
  INV_X1 u0_u11_u3_U26 (.A( u0_u11_u3_n130 ) , .ZN( u0_u11_u3_n177 ) );
  INV_X1 u0_u11_u3_U27 (.A( u0_u11_u3_n128 ) , .ZN( u0_u11_u3_n176 ) );
  NAND2_X1 u0_u11_u3_U28 (.ZN( u0_u11_u3_n105 ) , .A2( u0_u11_u3_n130 ) , .A1( u0_u11_u3_n155 ) );
  INV_X1 u0_u11_u3_U29 (.A( u0_u11_u3_n155 ) , .ZN( u0_u11_u3_n174 ) );
  INV_X1 u0_u11_u3_U3 (.A( u0_u11_u3_n140 ) , .ZN( u0_u11_u3_n182 ) );
  INV_X1 u0_u11_u3_U30 (.A( u0_u11_u3_n139 ) , .ZN( u0_u11_u3_n185 ) );
  NOR2_X1 u0_u11_u3_U31 (.ZN( u0_u11_u3_n135 ) , .A2( u0_u11_u3_n141 ) , .A1( u0_u11_u3_n169 ) );
  INV_X1 u0_u11_u3_U32 (.A( u0_u11_u3_n156 ) , .ZN( u0_u11_u3_n179 ) );
  OAI22_X1 u0_u11_u3_U33 (.B1( u0_u11_u3_n118 ) , .ZN( u0_u11_u3_n120 ) , .A1( u0_u11_u3_n135 ) , .B2( u0_u11_u3_n154 ) , .A2( u0_u11_u3_n178 ) );
  AND3_X1 u0_u11_u3_U34 (.ZN( u0_u11_u3_n118 ) , .A2( u0_u11_u3_n124 ) , .A1( u0_u11_u3_n144 ) , .A3( u0_u11_u3_n152 ) );
  OAI222_X1 u0_u11_u3_U35 (.C2( u0_u11_u3_n107 ) , .A2( u0_u11_u3_n108 ) , .B1( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n138 ) , .B2( u0_u11_u3_n146 ) , .C1( u0_u11_u3_n154 ) , .A1( u0_u11_u3_n164 ) );
  NOR4_X1 u0_u11_u3_U36 (.A4( u0_u11_u3_n157 ) , .A3( u0_u11_u3_n158 ) , .A2( u0_u11_u3_n159 ) , .A1( u0_u11_u3_n160 ) , .ZN( u0_u11_u3_n161 ) );
  AOI21_X1 u0_u11_u3_U37 (.B2( u0_u11_u3_n152 ) , .B1( u0_u11_u3_n153 ) , .ZN( u0_u11_u3_n158 ) , .A( u0_u11_u3_n164 ) );
  AOI21_X1 u0_u11_u3_U38 (.A( u0_u11_u3_n154 ) , .B2( u0_u11_u3_n155 ) , .B1( u0_u11_u3_n156 ) , .ZN( u0_u11_u3_n157 ) );
  AOI21_X1 u0_u11_u3_U39 (.A( u0_u11_u3_n149 ) , .B2( u0_u11_u3_n150 ) , .B1( u0_u11_u3_n151 ) , .ZN( u0_u11_u3_n159 ) );
  INV_X1 u0_u11_u3_U4 (.A( u0_u11_u3_n129 ) , .ZN( u0_u11_u3_n183 ) );
  AOI211_X1 u0_u11_u3_U40 (.ZN( u0_u11_u3_n109 ) , .A( u0_u11_u3_n119 ) , .C2( u0_u11_u3_n129 ) , .B( u0_u11_u3_n138 ) , .C1( u0_u11_u3_n141 ) );
  INV_X1 u0_u11_u3_U41 (.A( u0_u11_u3_n121 ) , .ZN( u0_u11_u3_n164 ) );
  NAND2_X1 u0_u11_u3_U42 (.ZN( u0_u11_u3_n133 ) , .A1( u0_u11_u3_n154 ) , .A2( u0_u11_u3_n164 ) );
  OAI211_X1 u0_u11_u3_U43 (.B( u0_u11_u3_n127 ) , .ZN( u0_u11_u3_n139 ) , .C1( u0_u11_u3_n150 ) , .C2( u0_u11_u3_n154 ) , .A( u0_u11_u3_n184 ) );
  INV_X1 u0_u11_u3_U44 (.A( u0_u11_u3_n125 ) , .ZN( u0_u11_u3_n184 ) );
  AOI221_X1 u0_u11_u3_U45 (.A( u0_u11_u3_n126 ) , .ZN( u0_u11_u3_n127 ) , .C2( u0_u11_u3_n132 ) , .C1( u0_u11_u3_n169 ) , .B2( u0_u11_u3_n170 ) , .B1( u0_u11_u3_n174 ) );
  OAI22_X1 u0_u11_u3_U46 (.A1( u0_u11_u3_n124 ) , .ZN( u0_u11_u3_n125 ) , .B2( u0_u11_u3_n145 ) , .A2( u0_u11_u3_n165 ) , .B1( u0_u11_u3_n167 ) );
  NOR2_X1 u0_u11_u3_U47 (.A1( u0_u11_u3_n113 ) , .ZN( u0_u11_u3_n131 ) , .A2( u0_u11_u3_n154 ) );
  NAND2_X1 u0_u11_u3_U48 (.A1( u0_u11_u3_n103 ) , .ZN( u0_u11_u3_n150 ) , .A2( u0_u11_u3_n99 ) );
  NAND2_X1 u0_u11_u3_U49 (.A2( u0_u11_u3_n102 ) , .ZN( u0_u11_u3_n155 ) , .A1( u0_u11_u3_n97 ) );
  INV_X1 u0_u11_u3_U5 (.A( u0_u11_u3_n117 ) , .ZN( u0_u11_u3_n178 ) );
  INV_X1 u0_u11_u3_U50 (.A( u0_u11_u3_n141 ) , .ZN( u0_u11_u3_n167 ) );
  AOI21_X1 u0_u11_u3_U51 (.B2( u0_u11_u3_n114 ) , .B1( u0_u11_u3_n146 ) , .A( u0_u11_u3_n154 ) , .ZN( u0_u11_u3_n94 ) );
  AOI21_X1 u0_u11_u3_U52 (.ZN( u0_u11_u3_n110 ) , .B2( u0_u11_u3_n142 ) , .B1( u0_u11_u3_n186 ) , .A( u0_u11_u3_n95 ) );
  INV_X1 u0_u11_u3_U53 (.A( u0_u11_u3_n145 ) , .ZN( u0_u11_u3_n186 ) );
  AOI21_X1 u0_u11_u3_U54 (.B1( u0_u11_u3_n124 ) , .A( u0_u11_u3_n149 ) , .B2( u0_u11_u3_n155 ) , .ZN( u0_u11_u3_n95 ) );
  INV_X1 u0_u11_u3_U55 (.A( u0_u11_u3_n149 ) , .ZN( u0_u11_u3_n169 ) );
  NAND2_X1 u0_u11_u3_U56 (.ZN( u0_u11_u3_n124 ) , .A1( u0_u11_u3_n96 ) , .A2( u0_u11_u3_n97 ) );
  NAND2_X1 u0_u11_u3_U57 (.A2( u0_u11_u3_n100 ) , .ZN( u0_u11_u3_n146 ) , .A1( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U58 (.A1( u0_u11_u3_n101 ) , .ZN( u0_u11_u3_n145 ) , .A2( u0_u11_u3_n99 ) );
  NAND2_X1 u0_u11_u3_U59 (.A1( u0_u11_u3_n100 ) , .ZN( u0_u11_u3_n156 ) , .A2( u0_u11_u3_n99 ) );
  AOI221_X1 u0_u11_u3_U6 (.A( u0_u11_u3_n131 ) , .C2( u0_u11_u3_n132 ) , .C1( u0_u11_u3_n133 ) , .ZN( u0_u11_u3_n134 ) , .B1( u0_u11_u3_n143 ) , .B2( u0_u11_u3_n177 ) );
  NAND2_X1 u0_u11_u3_U60 (.A2( u0_u11_u3_n101 ) , .A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n148 ) );
  NAND2_X1 u0_u11_u3_U61 (.A1( u0_u11_u3_n100 ) , .A2( u0_u11_u3_n102 ) , .ZN( u0_u11_u3_n128 ) );
  NAND2_X1 u0_u11_u3_U62 (.A2( u0_u11_u3_n101 ) , .A1( u0_u11_u3_n102 ) , .ZN( u0_u11_u3_n152 ) );
  NAND2_X1 u0_u11_u3_U63 (.A2( u0_u11_u3_n101 ) , .ZN( u0_u11_u3_n114 ) , .A1( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U64 (.ZN( u0_u11_u3_n107 ) , .A1( u0_u11_u3_n97 ) , .A2( u0_u11_u3_n99 ) );
  NAND2_X1 u0_u11_u3_U65 (.A2( u0_u11_u3_n100 ) , .A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n113 ) );
  NAND2_X1 u0_u11_u3_U66 (.A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n153 ) , .A2( u0_u11_u3_n97 ) );
  NAND2_X1 u0_u11_u3_U67 (.A2( u0_u11_u3_n103 ) , .A1( u0_u11_u3_n104 ) , .ZN( u0_u11_u3_n130 ) );
  NAND2_X1 u0_u11_u3_U68 (.A2( u0_u11_u3_n103 ) , .ZN( u0_u11_u3_n144 ) , .A1( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U69 (.A1( u0_u11_u3_n102 ) , .A2( u0_u11_u3_n103 ) , .ZN( u0_u11_u3_n108 ) );
  OAI22_X1 u0_u11_u3_U7 (.B2( u0_u11_u3_n147 ) , .A2( u0_u11_u3_n148 ) , .ZN( u0_u11_u3_n160 ) , .B1( u0_u11_u3_n165 ) , .A1( u0_u11_u3_n168 ) );
  NOR2_X1 u0_u11_u3_U70 (.A2( u0_u11_X_19 ) , .A1( u0_u11_X_20 ) , .ZN( u0_u11_u3_n99 ) );
  NOR2_X1 u0_u11_u3_U71 (.A2( u0_u11_X_21 ) , .A1( u0_u11_X_24 ) , .ZN( u0_u11_u3_n103 ) );
  NOR2_X1 u0_u11_u3_U72 (.A2( u0_u11_X_24 ) , .A1( u0_u11_u3_n171 ) , .ZN( u0_u11_u3_n97 ) );
  NOR2_X1 u0_u11_u3_U73 (.A2( u0_u11_X_19 ) , .A1( u0_u11_u3_n172 ) , .ZN( u0_u11_u3_n96 ) );
  NAND2_X1 u0_u11_u3_U74 (.A1( u0_u11_X_22 ) , .A2( u0_u11_X_23 ) , .ZN( u0_u11_u3_n154 ) );
  AND2_X1 u0_u11_u3_U75 (.A1( u0_u11_X_24 ) , .ZN( u0_u11_u3_n101 ) , .A2( u0_u11_u3_n171 ) );
  AND2_X1 u0_u11_u3_U76 (.A1( u0_u11_X_19 ) , .ZN( u0_u11_u3_n102 ) , .A2( u0_u11_u3_n172 ) );
  AND2_X1 u0_u11_u3_U77 (.A1( u0_u11_X_21 ) , .A2( u0_u11_X_24 ) , .ZN( u0_u11_u3_n100 ) );
  AND2_X1 u0_u11_u3_U78 (.A2( u0_u11_X_19 ) , .A1( u0_u11_X_20 ) , .ZN( u0_u11_u3_n104 ) );
  INV_X1 u0_u11_u3_U79 (.A( u0_u11_X_21 ) , .ZN( u0_u11_u3_n171 ) );
  AND3_X1 u0_u11_u3_U8 (.A3( u0_u11_u3_n144 ) , .A2( u0_u11_u3_n145 ) , .A1( u0_u11_u3_n146 ) , .ZN( u0_u11_u3_n147 ) );
  INV_X1 u0_u11_u3_U80 (.A( u0_u11_X_20 ) , .ZN( u0_u11_u3_n172 ) );
  INV_X1 u0_u11_u3_U81 (.A( u0_u11_X_22 ) , .ZN( u0_u11_u3_n166 ) );
  NAND4_X1 u0_u11_u3_U82 (.ZN( u0_out11_26 ) , .A4( u0_u11_u3_n109 ) , .A3( u0_u11_u3_n110 ) , .A2( u0_u11_u3_n111 ) , .A1( u0_u11_u3_n173 ) );
  INV_X1 u0_u11_u3_U83 (.ZN( u0_u11_u3_n173 ) , .A( u0_u11_u3_n94 ) );
  OAI21_X1 u0_u11_u3_U84 (.ZN( u0_u11_u3_n111 ) , .B2( u0_u11_u3_n117 ) , .A( u0_u11_u3_n133 ) , .B1( u0_u11_u3_n176 ) );
  NAND4_X1 u0_u11_u3_U85 (.ZN( u0_out11_1 ) , .A4( u0_u11_u3_n161 ) , .A3( u0_u11_u3_n162 ) , .A2( u0_u11_u3_n163 ) , .A1( u0_u11_u3_n185 ) );
  NAND2_X1 u0_u11_u3_U86 (.ZN( u0_u11_u3_n163 ) , .A2( u0_u11_u3_n170 ) , .A1( u0_u11_u3_n176 ) );
  AOI22_X1 u0_u11_u3_U87 (.B2( u0_u11_u3_n140 ) , .B1( u0_u11_u3_n141 ) , .A2( u0_u11_u3_n142 ) , .ZN( u0_u11_u3_n162 ) , .A1( u0_u11_u3_n177 ) );
  NAND4_X1 u0_u11_u3_U88 (.ZN( u0_out11_20 ) , .A4( u0_u11_u3_n122 ) , .A3( u0_u11_u3_n123 ) , .A1( u0_u11_u3_n175 ) , .A2( u0_u11_u3_n180 ) );
  INV_X1 u0_u11_u3_U89 (.A( u0_u11_u3_n126 ) , .ZN( u0_u11_u3_n180 ) );
  INV_X1 u0_u11_u3_U9 (.A( u0_u11_u3_n143 ) , .ZN( u0_u11_u3_n168 ) );
  INV_X1 u0_u11_u3_U90 (.A( u0_u11_u3_n112 ) , .ZN( u0_u11_u3_n175 ) );
  OR4_X1 u0_u11_u3_U91 (.ZN( u0_out11_10 ) , .A4( u0_u11_u3_n136 ) , .A3( u0_u11_u3_n137 ) , .A1( u0_u11_u3_n138 ) , .A2( u0_u11_u3_n139 ) );
  OAI222_X1 u0_u11_u3_U92 (.C1( u0_u11_u3_n128 ) , .ZN( u0_u11_u3_n137 ) , .B1( u0_u11_u3_n148 ) , .A2( u0_u11_u3_n150 ) , .B2( u0_u11_u3_n154 ) , .C2( u0_u11_u3_n164 ) , .A1( u0_u11_u3_n167 ) );
  AOI211_X1 u0_u11_u3_U93 (.B( u0_u11_u3_n119 ) , .A( u0_u11_u3_n120 ) , .C2( u0_u11_u3_n121 ) , .ZN( u0_u11_u3_n122 ) , .C1( u0_u11_u3_n179 ) );
  OAI221_X1 u0_u11_u3_U94 (.A( u0_u11_u3_n134 ) , .B2( u0_u11_u3_n135 ) , .ZN( u0_u11_u3_n136 ) , .C1( u0_u11_u3_n149 ) , .B1( u0_u11_u3_n151 ) , .C2( u0_u11_u3_n183 ) );
  NOR2_X1 u0_u11_u3_U95 (.A2( u0_u11_X_23 ) , .ZN( u0_u11_u3_n141 ) , .A1( u0_u11_u3_n166 ) );
  NAND2_X1 u0_u11_u3_U96 (.A1( u0_u11_X_23 ) , .ZN( u0_u11_u3_n149 ) , .A2( u0_u11_u3_n166 ) );
  NOR2_X1 u0_u11_u3_U97 (.A2( u0_u11_X_22 ) , .A1( u0_u11_X_23 ) , .ZN( u0_u11_u3_n121 ) );
  NAND3_X1 u0_u11_u3_U98 (.A1( u0_u11_u3_n114 ) , .ZN( u0_u11_u3_n115 ) , .A2( u0_u11_u3_n145 ) , .A3( u0_u11_u3_n153 ) );
  NAND3_X1 u0_u11_u3_U99 (.ZN( u0_u11_u3_n129 ) , .A2( u0_u11_u3_n144 ) , .A1( u0_u11_u3_n153 ) , .A3( u0_u11_u3_n182 ) );
  INV_X1 u0_u11_u5_U10 (.A( u0_u11_u5_n121 ) , .ZN( u0_u11_u5_n177 ) );
  NOR3_X1 u0_u11_u5_U100 (.A3( u0_u11_u5_n141 ) , .A1( u0_u11_u5_n142 ) , .ZN( u0_u11_u5_n143 ) , .A2( u0_u11_u5_n191 ) );
  NAND4_X1 u0_u11_u5_U101 (.ZN( u0_out11_4 ) , .A4( u0_u11_u5_n112 ) , .A2( u0_u11_u5_n113 ) , .A1( u0_u11_u5_n114 ) , .A3( u0_u11_u5_n195 ) );
  AOI211_X1 u0_u11_u5_U102 (.A( u0_u11_u5_n110 ) , .C1( u0_u11_u5_n111 ) , .ZN( u0_u11_u5_n112 ) , .B( u0_u11_u5_n118 ) , .C2( u0_u11_u5_n177 ) );
  AOI222_X1 u0_u11_u5_U103 (.ZN( u0_u11_u5_n113 ) , .A1( u0_u11_u5_n131 ) , .C1( u0_u11_u5_n148 ) , .B2( u0_u11_u5_n174 ) , .C2( u0_u11_u5_n178 ) , .A2( u0_u11_u5_n179 ) , .B1( u0_u11_u5_n99 ) );
  NAND3_X1 u0_u11_u5_U104 (.A2( u0_u11_u5_n154 ) , .A3( u0_u11_u5_n158 ) , .A1( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n99 ) );
  NOR2_X1 u0_u11_u5_U11 (.ZN( u0_u11_u5_n160 ) , .A2( u0_u11_u5_n173 ) , .A1( u0_u11_u5_n177 ) );
  INV_X1 u0_u11_u5_U12 (.A( u0_u11_u5_n150 ) , .ZN( u0_u11_u5_n174 ) );
  AOI21_X1 u0_u11_u5_U13 (.A( u0_u11_u5_n160 ) , .B2( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n162 ) , .B1( u0_u11_u5_n192 ) );
  INV_X1 u0_u11_u5_U14 (.A( u0_u11_u5_n159 ) , .ZN( u0_u11_u5_n192 ) );
  AOI21_X1 u0_u11_u5_U15 (.A( u0_u11_u5_n156 ) , .B2( u0_u11_u5_n157 ) , .B1( u0_u11_u5_n158 ) , .ZN( u0_u11_u5_n163 ) );
  AOI21_X1 u0_u11_u5_U16 (.B2( u0_u11_u5_n139 ) , .B1( u0_u11_u5_n140 ) , .ZN( u0_u11_u5_n141 ) , .A( u0_u11_u5_n150 ) );
  OAI21_X1 u0_u11_u5_U17 (.A( u0_u11_u5_n133 ) , .B2( u0_u11_u5_n134 ) , .B1( u0_u11_u5_n135 ) , .ZN( u0_u11_u5_n142 ) );
  OAI21_X1 u0_u11_u5_U18 (.ZN( u0_u11_u5_n133 ) , .B2( u0_u11_u5_n147 ) , .A( u0_u11_u5_n173 ) , .B1( u0_u11_u5_n188 ) );
  NAND2_X1 u0_u11_u5_U19 (.A2( u0_u11_u5_n119 ) , .A1( u0_u11_u5_n123 ) , .ZN( u0_u11_u5_n137 ) );
  INV_X1 u0_u11_u5_U20 (.A( u0_u11_u5_n155 ) , .ZN( u0_u11_u5_n194 ) );
  NAND2_X1 u0_u11_u5_U21 (.A1( u0_u11_u5_n121 ) , .ZN( u0_u11_u5_n132 ) , .A2( u0_u11_u5_n172 ) );
  NAND2_X1 u0_u11_u5_U22 (.A2( u0_u11_u5_n122 ) , .ZN( u0_u11_u5_n136 ) , .A1( u0_u11_u5_n154 ) );
  NAND2_X1 u0_u11_u5_U23 (.A2( u0_u11_u5_n119 ) , .A1( u0_u11_u5_n120 ) , .ZN( u0_u11_u5_n159 ) );
  INV_X1 u0_u11_u5_U24 (.A( u0_u11_u5_n156 ) , .ZN( u0_u11_u5_n175 ) );
  INV_X1 u0_u11_u5_U25 (.A( u0_u11_u5_n158 ) , .ZN( u0_u11_u5_n188 ) );
  INV_X1 u0_u11_u5_U26 (.A( u0_u11_u5_n152 ) , .ZN( u0_u11_u5_n179 ) );
  INV_X1 u0_u11_u5_U27 (.A( u0_u11_u5_n140 ) , .ZN( u0_u11_u5_n182 ) );
  INV_X1 u0_u11_u5_U28 (.A( u0_u11_u5_n151 ) , .ZN( u0_u11_u5_n183 ) );
  INV_X1 u0_u11_u5_U29 (.A( u0_u11_u5_n123 ) , .ZN( u0_u11_u5_n185 ) );
  NOR2_X1 u0_u11_u5_U3 (.ZN( u0_u11_u5_n134 ) , .A1( u0_u11_u5_n183 ) , .A2( u0_u11_u5_n190 ) );
  INV_X1 u0_u11_u5_U30 (.A( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n184 ) );
  INV_X1 u0_u11_u5_U31 (.A( u0_u11_u5_n139 ) , .ZN( u0_u11_u5_n189 ) );
  INV_X1 u0_u11_u5_U32 (.A( u0_u11_u5_n157 ) , .ZN( u0_u11_u5_n190 ) );
  INV_X1 u0_u11_u5_U33 (.A( u0_u11_u5_n120 ) , .ZN( u0_u11_u5_n193 ) );
  NAND2_X1 u0_u11_u5_U34 (.ZN( u0_u11_u5_n111 ) , .A1( u0_u11_u5_n140 ) , .A2( u0_u11_u5_n155 ) );
  NOR2_X1 u0_u11_u5_U35 (.ZN( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n170 ) , .A2( u0_u11_u5_n180 ) );
  INV_X1 u0_u11_u5_U36 (.A( u0_u11_u5_n117 ) , .ZN( u0_u11_u5_n196 ) );
  OAI221_X1 u0_u11_u5_U37 (.A( u0_u11_u5_n116 ) , .ZN( u0_u11_u5_n117 ) , .B2( u0_u11_u5_n119 ) , .C1( u0_u11_u5_n153 ) , .C2( u0_u11_u5_n158 ) , .B1( u0_u11_u5_n172 ) );
  AOI222_X1 u0_u11_u5_U38 (.ZN( u0_u11_u5_n116 ) , .B2( u0_u11_u5_n145 ) , .C1( u0_u11_u5_n148 ) , .A2( u0_u11_u5_n174 ) , .C2( u0_u11_u5_n177 ) , .B1( u0_u11_u5_n187 ) , .A1( u0_u11_u5_n193 ) );
  INV_X1 u0_u11_u5_U39 (.A( u0_u11_u5_n115 ) , .ZN( u0_u11_u5_n187 ) );
  INV_X1 u0_u11_u5_U4 (.A( u0_u11_u5_n138 ) , .ZN( u0_u11_u5_n191 ) );
  AOI22_X1 u0_u11_u5_U40 (.B2( u0_u11_u5_n131 ) , .A2( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n169 ) , .B1( u0_u11_u5_n174 ) , .A1( u0_u11_u5_n185 ) );
  NOR2_X1 u0_u11_u5_U41 (.A1( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n150 ) , .A2( u0_u11_u5_n173 ) );
  AOI21_X1 u0_u11_u5_U42 (.A( u0_u11_u5_n118 ) , .B2( u0_u11_u5_n145 ) , .ZN( u0_u11_u5_n168 ) , .B1( u0_u11_u5_n186 ) );
  INV_X1 u0_u11_u5_U43 (.A( u0_u11_u5_n122 ) , .ZN( u0_u11_u5_n186 ) );
  NOR2_X1 u0_u11_u5_U44 (.A1( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n152 ) , .A2( u0_u11_u5_n176 ) );
  NOR2_X1 u0_u11_u5_U45 (.A1( u0_u11_u5_n115 ) , .ZN( u0_u11_u5_n118 ) , .A2( u0_u11_u5_n153 ) );
  NOR2_X1 u0_u11_u5_U46 (.A2( u0_u11_u5_n145 ) , .ZN( u0_u11_u5_n156 ) , .A1( u0_u11_u5_n174 ) );
  NOR2_X1 u0_u11_u5_U47 (.ZN( u0_u11_u5_n121 ) , .A2( u0_u11_u5_n145 ) , .A1( u0_u11_u5_n176 ) );
  AOI22_X1 u0_u11_u5_U48 (.ZN( u0_u11_u5_n114 ) , .A2( u0_u11_u5_n137 ) , .A1( u0_u11_u5_n145 ) , .B2( u0_u11_u5_n175 ) , .B1( u0_u11_u5_n193 ) );
  OAI211_X1 u0_u11_u5_U49 (.B( u0_u11_u5_n124 ) , .A( u0_u11_u5_n125 ) , .C2( u0_u11_u5_n126 ) , .C1( u0_u11_u5_n127 ) , .ZN( u0_u11_u5_n128 ) );
  OAI21_X1 u0_u11_u5_U5 (.B2( u0_u11_u5_n136 ) , .B1( u0_u11_u5_n137 ) , .ZN( u0_u11_u5_n138 ) , .A( u0_u11_u5_n177 ) );
  OAI21_X1 u0_u11_u5_U50 (.ZN( u0_u11_u5_n124 ) , .A( u0_u11_u5_n177 ) , .B2( u0_u11_u5_n183 ) , .B1( u0_u11_u5_n189 ) );
  NOR3_X1 u0_u11_u5_U51 (.ZN( u0_u11_u5_n127 ) , .A1( u0_u11_u5_n136 ) , .A3( u0_u11_u5_n148 ) , .A2( u0_u11_u5_n182 ) );
  OAI21_X1 u0_u11_u5_U52 (.ZN( u0_u11_u5_n125 ) , .A( u0_u11_u5_n174 ) , .B2( u0_u11_u5_n185 ) , .B1( u0_u11_u5_n190 ) );
  AOI21_X1 u0_u11_u5_U53 (.A( u0_u11_u5_n153 ) , .B2( u0_u11_u5_n154 ) , .B1( u0_u11_u5_n155 ) , .ZN( u0_u11_u5_n164 ) );
  AOI21_X1 u0_u11_u5_U54 (.ZN( u0_u11_u5_n110 ) , .B1( u0_u11_u5_n122 ) , .B2( u0_u11_u5_n139 ) , .A( u0_u11_u5_n153 ) );
  INV_X1 u0_u11_u5_U55 (.A( u0_u11_u5_n153 ) , .ZN( u0_u11_u5_n176 ) );
  INV_X1 u0_u11_u5_U56 (.A( u0_u11_u5_n126 ) , .ZN( u0_u11_u5_n173 ) );
  AND2_X1 u0_u11_u5_U57 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n147 ) );
  AND2_X1 u0_u11_u5_U58 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n148 ) );
  NAND2_X1 u0_u11_u5_U59 (.A1( u0_u11_u5_n105 ) , .A2( u0_u11_u5_n106 ) , .ZN( u0_u11_u5_n158 ) );
  INV_X1 u0_u11_u5_U6 (.A( u0_u11_u5_n135 ) , .ZN( u0_u11_u5_n178 ) );
  NAND2_X1 u0_u11_u5_U60 (.A2( u0_u11_u5_n108 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n139 ) );
  NAND2_X1 u0_u11_u5_U61 (.A1( u0_u11_u5_n106 ) , .A2( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n119 ) );
  NAND2_X1 u0_u11_u5_U62 (.A2( u0_u11_u5_n103 ) , .A1( u0_u11_u5_n105 ) , .ZN( u0_u11_u5_n140 ) );
  NAND2_X1 u0_u11_u5_U63 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n105 ) , .ZN( u0_u11_u5_n155 ) );
  NAND2_X1 u0_u11_u5_U64 (.A2( u0_u11_u5_n106 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n122 ) );
  NAND2_X1 u0_u11_u5_U65 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n106 ) , .ZN( u0_u11_u5_n115 ) );
  NAND2_X1 u0_u11_u5_U66 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n103 ) , .ZN( u0_u11_u5_n161 ) );
  NAND2_X1 u0_u11_u5_U67 (.A1( u0_u11_u5_n105 ) , .A2( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n154 ) );
  INV_X1 u0_u11_u5_U68 (.A( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n172 ) );
  NAND2_X1 u0_u11_u5_U69 (.A1( u0_u11_u5_n103 ) , .A2( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n123 ) );
  OAI22_X1 u0_u11_u5_U7 (.B2( u0_u11_u5_n149 ) , .B1( u0_u11_u5_n150 ) , .A2( u0_u11_u5_n151 ) , .A1( u0_u11_u5_n152 ) , .ZN( u0_u11_u5_n165 ) );
  NAND2_X1 u0_u11_u5_U70 (.A2( u0_u11_u5_n103 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n151 ) );
  NAND2_X1 u0_u11_u5_U71 (.A2( u0_u11_u5_n107 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n120 ) );
  NAND2_X1 u0_u11_u5_U72 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n157 ) );
  AND2_X1 u0_u11_u5_U73 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n104 ) , .ZN( u0_u11_u5_n131 ) );
  INV_X1 u0_u11_u5_U74 (.A( u0_u11_u5_n102 ) , .ZN( u0_u11_u5_n195 ) );
  OAI221_X1 u0_u11_u5_U75 (.A( u0_u11_u5_n101 ) , .ZN( u0_u11_u5_n102 ) , .C2( u0_u11_u5_n115 ) , .C1( u0_u11_u5_n126 ) , .B1( u0_u11_u5_n134 ) , .B2( u0_u11_u5_n160 ) );
  OAI21_X1 u0_u11_u5_U76 (.ZN( u0_u11_u5_n101 ) , .B1( u0_u11_u5_n137 ) , .A( u0_u11_u5_n146 ) , .B2( u0_u11_u5_n147 ) );
  NOR2_X1 u0_u11_u5_U77 (.A2( u0_u11_X_34 ) , .A1( u0_u11_X_35 ) , .ZN( u0_u11_u5_n145 ) );
  NOR2_X1 u0_u11_u5_U78 (.A2( u0_u11_X_34 ) , .ZN( u0_u11_u5_n146 ) , .A1( u0_u11_u5_n171 ) );
  NOR2_X1 u0_u11_u5_U79 (.A2( u0_u11_X_31 ) , .A1( u0_u11_X_32 ) , .ZN( u0_u11_u5_n103 ) );
  NOR3_X1 u0_u11_u5_U8 (.A2( u0_u11_u5_n147 ) , .A1( u0_u11_u5_n148 ) , .ZN( u0_u11_u5_n149 ) , .A3( u0_u11_u5_n194 ) );
  NOR2_X1 u0_u11_u5_U80 (.A2( u0_u11_X_36 ) , .ZN( u0_u11_u5_n105 ) , .A1( u0_u11_u5_n180 ) );
  NOR2_X1 u0_u11_u5_U81 (.A2( u0_u11_X_33 ) , .ZN( u0_u11_u5_n108 ) , .A1( u0_u11_u5_n170 ) );
  NOR2_X1 u0_u11_u5_U82 (.A2( u0_u11_X_33 ) , .A1( u0_u11_X_36 ) , .ZN( u0_u11_u5_n107 ) );
  NOR2_X1 u0_u11_u5_U83 (.A2( u0_u11_X_31 ) , .ZN( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n181 ) );
  NAND2_X1 u0_u11_u5_U84 (.A2( u0_u11_X_34 ) , .A1( u0_u11_X_35 ) , .ZN( u0_u11_u5_n153 ) );
  NAND2_X1 u0_u11_u5_U85 (.A1( u0_u11_X_34 ) , .ZN( u0_u11_u5_n126 ) , .A2( u0_u11_u5_n171 ) );
  AND2_X1 u0_u11_u5_U86 (.A1( u0_u11_X_31 ) , .A2( u0_u11_X_32 ) , .ZN( u0_u11_u5_n106 ) );
  AND2_X1 u0_u11_u5_U87 (.A1( u0_u11_X_31 ) , .ZN( u0_u11_u5_n109 ) , .A2( u0_u11_u5_n181 ) );
  INV_X1 u0_u11_u5_U88 (.A( u0_u11_X_33 ) , .ZN( u0_u11_u5_n180 ) );
  INV_X1 u0_u11_u5_U89 (.A( u0_u11_X_35 ) , .ZN( u0_u11_u5_n171 ) );
  NOR2_X1 u0_u11_u5_U9 (.ZN( u0_u11_u5_n135 ) , .A1( u0_u11_u5_n173 ) , .A2( u0_u11_u5_n176 ) );
  INV_X1 u0_u11_u5_U90 (.A( u0_u11_X_36 ) , .ZN( u0_u11_u5_n170 ) );
  INV_X1 u0_u11_u5_U91 (.A( u0_u11_X_32 ) , .ZN( u0_u11_u5_n181 ) );
  NAND4_X1 u0_u11_u5_U92 (.ZN( u0_out11_29 ) , .A4( u0_u11_u5_n129 ) , .A3( u0_u11_u5_n130 ) , .A2( u0_u11_u5_n168 ) , .A1( u0_u11_u5_n196 ) );
  AOI221_X1 u0_u11_u5_U93 (.A( u0_u11_u5_n128 ) , .ZN( u0_u11_u5_n129 ) , .C2( u0_u11_u5_n132 ) , .B2( u0_u11_u5_n159 ) , .B1( u0_u11_u5_n176 ) , .C1( u0_u11_u5_n184 ) );
  AOI222_X1 u0_u11_u5_U94 (.ZN( u0_u11_u5_n130 ) , .A2( u0_u11_u5_n146 ) , .B1( u0_u11_u5_n147 ) , .C2( u0_u11_u5_n175 ) , .B2( u0_u11_u5_n179 ) , .A1( u0_u11_u5_n188 ) , .C1( u0_u11_u5_n194 ) );
  NAND4_X1 u0_u11_u5_U95 (.ZN( u0_out11_19 ) , .A4( u0_u11_u5_n166 ) , .A3( u0_u11_u5_n167 ) , .A2( u0_u11_u5_n168 ) , .A1( u0_u11_u5_n169 ) );
  AOI22_X1 u0_u11_u5_U96 (.B2( u0_u11_u5_n145 ) , .A2( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n167 ) , .B1( u0_u11_u5_n182 ) , .A1( u0_u11_u5_n189 ) );
  NOR4_X1 u0_u11_u5_U97 (.A4( u0_u11_u5_n162 ) , .A3( u0_u11_u5_n163 ) , .A2( u0_u11_u5_n164 ) , .A1( u0_u11_u5_n165 ) , .ZN( u0_u11_u5_n166 ) );
  NAND4_X1 u0_u11_u5_U98 (.ZN( u0_out11_11 ) , .A4( u0_u11_u5_n143 ) , .A3( u0_u11_u5_n144 ) , .A2( u0_u11_u5_n169 ) , .A1( u0_u11_u5_n196 ) );
  AOI22_X1 u0_u11_u5_U99 (.A2( u0_u11_u5_n132 ) , .ZN( u0_u11_u5_n144 ) , .B2( u0_u11_u5_n145 ) , .B1( u0_u11_u5_n184 ) , .A1( u0_u11_u5_n194 ) );
  OAI21_X1 u0_u11_u6_U10 (.A( u0_u11_u6_n159 ) , .B1( u0_u11_u6_n169 ) , .B2( u0_u11_u6_n173 ) , .ZN( u0_u11_u6_n90 ) );
  INV_X1 u0_u11_u6_U11 (.ZN( u0_u11_u6_n172 ) , .A( u0_u11_u6_n88 ) );
  AOI22_X1 u0_u11_u6_U12 (.A2( u0_u11_u6_n151 ) , .B2( u0_u11_u6_n161 ) , .A1( u0_u11_u6_n167 ) , .B1( u0_u11_u6_n170 ) , .ZN( u0_u11_u6_n89 ) );
  AOI21_X1 u0_u11_u6_U13 (.ZN( u0_u11_u6_n106 ) , .A( u0_u11_u6_n142 ) , .B2( u0_u11_u6_n159 ) , .B1( u0_u11_u6_n164 ) );
  INV_X1 u0_u11_u6_U14 (.A( u0_u11_u6_n155 ) , .ZN( u0_u11_u6_n161 ) );
  INV_X1 u0_u11_u6_U15 (.A( u0_u11_u6_n128 ) , .ZN( u0_u11_u6_n164 ) );
  NAND2_X1 u0_u11_u6_U16 (.ZN( u0_u11_u6_n110 ) , .A1( u0_u11_u6_n122 ) , .A2( u0_u11_u6_n129 ) );
  NAND2_X1 u0_u11_u6_U17 (.ZN( u0_u11_u6_n124 ) , .A2( u0_u11_u6_n146 ) , .A1( u0_u11_u6_n148 ) );
  INV_X1 u0_u11_u6_U18 (.A( u0_u11_u6_n132 ) , .ZN( u0_u11_u6_n171 ) );
  AND2_X1 u0_u11_u6_U19 (.A1( u0_u11_u6_n100 ) , .ZN( u0_u11_u6_n130 ) , .A2( u0_u11_u6_n147 ) );
  INV_X1 u0_u11_u6_U20 (.A( u0_u11_u6_n127 ) , .ZN( u0_u11_u6_n173 ) );
  INV_X1 u0_u11_u6_U21 (.A( u0_u11_u6_n121 ) , .ZN( u0_u11_u6_n167 ) );
  INV_X1 u0_u11_u6_U22 (.A( u0_u11_u6_n100 ) , .ZN( u0_u11_u6_n169 ) );
  INV_X1 u0_u11_u6_U23 (.A( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n170 ) );
  INV_X1 u0_u11_u6_U24 (.A( u0_u11_u6_n113 ) , .ZN( u0_u11_u6_n168 ) );
  AND2_X1 u0_u11_u6_U25 (.A1( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n119 ) , .ZN( u0_u11_u6_n133 ) );
  AND2_X1 u0_u11_u6_U26 (.A2( u0_u11_u6_n121 ) , .A1( u0_u11_u6_n122 ) , .ZN( u0_u11_u6_n131 ) );
  AND3_X1 u0_u11_u6_U27 (.ZN( u0_u11_u6_n120 ) , .A2( u0_u11_u6_n127 ) , .A1( u0_u11_u6_n132 ) , .A3( u0_u11_u6_n145 ) );
  INV_X1 u0_u11_u6_U28 (.A( u0_u11_u6_n146 ) , .ZN( u0_u11_u6_n163 ) );
  AOI222_X1 u0_u11_u6_U29 (.ZN( u0_u11_u6_n114 ) , .A1( u0_u11_u6_n118 ) , .A2( u0_u11_u6_n126 ) , .B2( u0_u11_u6_n151 ) , .C2( u0_u11_u6_n159 ) , .C1( u0_u11_u6_n168 ) , .B1( u0_u11_u6_n169 ) );
  INV_X1 u0_u11_u6_U3 (.A( u0_u11_u6_n110 ) , .ZN( u0_u11_u6_n166 ) );
  NOR2_X1 u0_u11_u6_U30 (.A1( u0_u11_u6_n162 ) , .A2( u0_u11_u6_n165 ) , .ZN( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U31 (.A1( u0_u11_u6_n144 ) , .ZN( u0_u11_u6_n151 ) , .A2( u0_u11_u6_n158 ) );
  NAND2_X1 u0_u11_u6_U32 (.ZN( u0_u11_u6_n132 ) , .A1( u0_u11_u6_n91 ) , .A2( u0_u11_u6_n97 ) );
  AOI22_X1 u0_u11_u6_U33 (.B2( u0_u11_u6_n110 ) , .B1( u0_u11_u6_n111 ) , .A1( u0_u11_u6_n112 ) , .ZN( u0_u11_u6_n115 ) , .A2( u0_u11_u6_n161 ) );
  NAND4_X1 u0_u11_u6_U34 (.A3( u0_u11_u6_n109 ) , .ZN( u0_u11_u6_n112 ) , .A4( u0_u11_u6_n132 ) , .A2( u0_u11_u6_n147 ) , .A1( u0_u11_u6_n166 ) );
  NOR2_X1 u0_u11_u6_U35 (.ZN( u0_u11_u6_n109 ) , .A1( u0_u11_u6_n170 ) , .A2( u0_u11_u6_n173 ) );
  NOR2_X1 u0_u11_u6_U36 (.A2( u0_u11_u6_n126 ) , .ZN( u0_u11_u6_n155 ) , .A1( u0_u11_u6_n160 ) );
  NAND2_X1 u0_u11_u6_U37 (.ZN( u0_u11_u6_n146 ) , .A2( u0_u11_u6_n94 ) , .A1( u0_u11_u6_n99 ) );
  AOI21_X1 u0_u11_u6_U38 (.A( u0_u11_u6_n144 ) , .B2( u0_u11_u6_n145 ) , .B1( u0_u11_u6_n146 ) , .ZN( u0_u11_u6_n150 ) );
  AOI211_X1 u0_u11_u6_U39 (.B( u0_u11_u6_n134 ) , .A( u0_u11_u6_n135 ) , .C1( u0_u11_u6_n136 ) , .ZN( u0_u11_u6_n137 ) , .C2( u0_u11_u6_n151 ) );
  INV_X1 u0_u11_u6_U4 (.A( u0_u11_u6_n142 ) , .ZN( u0_u11_u6_n174 ) );
  NAND4_X1 u0_u11_u6_U40 (.A4( u0_u11_u6_n127 ) , .A3( u0_u11_u6_n128 ) , .A2( u0_u11_u6_n129 ) , .A1( u0_u11_u6_n130 ) , .ZN( u0_u11_u6_n136 ) );
  AOI21_X1 u0_u11_u6_U41 (.B2( u0_u11_u6_n132 ) , .B1( u0_u11_u6_n133 ) , .ZN( u0_u11_u6_n134 ) , .A( u0_u11_u6_n158 ) );
  AOI21_X1 u0_u11_u6_U42 (.B1( u0_u11_u6_n131 ) , .ZN( u0_u11_u6_n135 ) , .A( u0_u11_u6_n144 ) , .B2( u0_u11_u6_n146 ) );
  INV_X1 u0_u11_u6_U43 (.A( u0_u11_u6_n111 ) , .ZN( u0_u11_u6_n158 ) );
  NAND2_X1 u0_u11_u6_U44 (.ZN( u0_u11_u6_n127 ) , .A1( u0_u11_u6_n91 ) , .A2( u0_u11_u6_n92 ) );
  NAND2_X1 u0_u11_u6_U45 (.ZN( u0_u11_u6_n129 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n96 ) );
  INV_X1 u0_u11_u6_U46 (.A( u0_u11_u6_n144 ) , .ZN( u0_u11_u6_n159 ) );
  NAND2_X1 u0_u11_u6_U47 (.ZN( u0_u11_u6_n145 ) , .A2( u0_u11_u6_n97 ) , .A1( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U48 (.ZN( u0_u11_u6_n148 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n94 ) );
  NAND2_X1 u0_u11_u6_U49 (.ZN( u0_u11_u6_n108 ) , .A2( u0_u11_u6_n139 ) , .A1( u0_u11_u6_n144 ) );
  NAND2_X1 u0_u11_u6_U5 (.A2( u0_u11_u6_n143 ) , .ZN( u0_u11_u6_n152 ) , .A1( u0_u11_u6_n166 ) );
  NAND2_X1 u0_u11_u6_U50 (.ZN( u0_u11_u6_n121 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n97 ) );
  NAND2_X1 u0_u11_u6_U51 (.ZN( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n95 ) );
  AND2_X1 u0_u11_u6_U52 (.ZN( u0_u11_u6_n118 ) , .A2( u0_u11_u6_n91 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U53 (.ZN( u0_u11_u6_n147 ) , .A2( u0_u11_u6_n98 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U54 (.ZN( u0_u11_u6_n128 ) , .A1( u0_u11_u6_n94 ) , .A2( u0_u11_u6_n96 ) );
  NAND2_X1 u0_u11_u6_U55 (.ZN( u0_u11_u6_n119 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U56 (.ZN( u0_u11_u6_n123 ) , .A2( u0_u11_u6_n91 ) , .A1( u0_u11_u6_n96 ) );
  NAND2_X1 u0_u11_u6_U57 (.ZN( u0_u11_u6_n100 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U58 (.ZN( u0_u11_u6_n122 ) , .A1( u0_u11_u6_n94 ) , .A2( u0_u11_u6_n97 ) );
  INV_X1 u0_u11_u6_U59 (.A( u0_u11_u6_n139 ) , .ZN( u0_u11_u6_n160 ) );
  AOI22_X1 u0_u11_u6_U6 (.B2( u0_u11_u6_n101 ) , .A1( u0_u11_u6_n102 ) , .ZN( u0_u11_u6_n103 ) , .B1( u0_u11_u6_n160 ) , .A2( u0_u11_u6_n161 ) );
  NAND2_X1 u0_u11_u6_U60 (.ZN( u0_u11_u6_n113 ) , .A1( u0_u11_u6_n96 ) , .A2( u0_u11_u6_n98 ) );
  NOR2_X1 u0_u11_u6_U61 (.A2( u0_u11_X_40 ) , .A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n126 ) );
  NOR2_X1 u0_u11_u6_U62 (.A2( u0_u11_X_39 ) , .A1( u0_u11_X_42 ) , .ZN( u0_u11_u6_n92 ) );
  NOR2_X1 u0_u11_u6_U63 (.A2( u0_u11_X_39 ) , .A1( u0_u11_u6_n156 ) , .ZN( u0_u11_u6_n97 ) );
  NOR2_X1 u0_u11_u6_U64 (.A2( u0_u11_X_38 ) , .A1( u0_u11_u6_n165 ) , .ZN( u0_u11_u6_n95 ) );
  NOR2_X1 u0_u11_u6_U65 (.A2( u0_u11_X_41 ) , .ZN( u0_u11_u6_n111 ) , .A1( u0_u11_u6_n157 ) );
  NOR2_X1 u0_u11_u6_U66 (.A2( u0_u11_X_37 ) , .A1( u0_u11_u6_n162 ) , .ZN( u0_u11_u6_n94 ) );
  NOR2_X1 u0_u11_u6_U67 (.A2( u0_u11_X_37 ) , .A1( u0_u11_X_38 ) , .ZN( u0_u11_u6_n91 ) );
  NAND2_X1 u0_u11_u6_U68 (.A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n144 ) , .A2( u0_u11_u6_n157 ) );
  NAND2_X1 u0_u11_u6_U69 (.A2( u0_u11_X_40 ) , .A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n139 ) );
  NOR2_X1 u0_u11_u6_U7 (.A1( u0_u11_u6_n118 ) , .ZN( u0_u11_u6_n143 ) , .A2( u0_u11_u6_n168 ) );
  AND2_X1 u0_u11_u6_U70 (.A1( u0_u11_X_39 ) , .A2( u0_u11_u6_n156 ) , .ZN( u0_u11_u6_n96 ) );
  AND2_X1 u0_u11_u6_U71 (.A1( u0_u11_X_39 ) , .A2( u0_u11_X_42 ) , .ZN( u0_u11_u6_n99 ) );
  INV_X1 u0_u11_u6_U72 (.A( u0_u11_X_40 ) , .ZN( u0_u11_u6_n157 ) );
  INV_X1 u0_u11_u6_U73 (.A( u0_u11_X_37 ) , .ZN( u0_u11_u6_n165 ) );
  INV_X1 u0_u11_u6_U74 (.A( u0_u11_X_38 ) , .ZN( u0_u11_u6_n162 ) );
  INV_X1 u0_u11_u6_U75 (.A( u0_u11_X_42 ) , .ZN( u0_u11_u6_n156 ) );
  NAND4_X1 u0_u11_u6_U76 (.ZN( u0_out11_32 ) , .A4( u0_u11_u6_n103 ) , .A3( u0_u11_u6_n104 ) , .A2( u0_u11_u6_n105 ) , .A1( u0_u11_u6_n106 ) );
  AOI22_X1 u0_u11_u6_U77 (.ZN( u0_u11_u6_n105 ) , .A2( u0_u11_u6_n108 ) , .A1( u0_u11_u6_n118 ) , .B2( u0_u11_u6_n126 ) , .B1( u0_u11_u6_n171 ) );
  AOI22_X1 u0_u11_u6_U78 (.ZN( u0_u11_u6_n104 ) , .A1( u0_u11_u6_n111 ) , .B1( u0_u11_u6_n124 ) , .B2( u0_u11_u6_n151 ) , .A2( u0_u11_u6_n93 ) );
  NAND4_X1 u0_u11_u6_U79 (.ZN( u0_out11_12 ) , .A4( u0_u11_u6_n114 ) , .A3( u0_u11_u6_n115 ) , .A2( u0_u11_u6_n116 ) , .A1( u0_u11_u6_n117 ) );
  AOI21_X1 u0_u11_u6_U8 (.B1( u0_u11_u6_n107 ) , .B2( u0_u11_u6_n132 ) , .A( u0_u11_u6_n158 ) , .ZN( u0_u11_u6_n88 ) );
  OAI22_X1 u0_u11_u6_U80 (.B2( u0_u11_u6_n111 ) , .ZN( u0_u11_u6_n116 ) , .B1( u0_u11_u6_n126 ) , .A2( u0_u11_u6_n164 ) , .A1( u0_u11_u6_n167 ) );
  OAI21_X1 u0_u11_u6_U81 (.A( u0_u11_u6_n108 ) , .ZN( u0_u11_u6_n117 ) , .B2( u0_u11_u6_n141 ) , .B1( u0_u11_u6_n163 ) );
  OAI211_X1 u0_u11_u6_U82 (.ZN( u0_out11_7 ) , .B( u0_u11_u6_n153 ) , .C2( u0_u11_u6_n154 ) , .C1( u0_u11_u6_n155 ) , .A( u0_u11_u6_n174 ) );
  NOR3_X1 u0_u11_u6_U83 (.A1( u0_u11_u6_n141 ) , .ZN( u0_u11_u6_n154 ) , .A3( u0_u11_u6_n164 ) , .A2( u0_u11_u6_n171 ) );
  AOI211_X1 u0_u11_u6_U84 (.B( u0_u11_u6_n149 ) , .A( u0_u11_u6_n150 ) , .C2( u0_u11_u6_n151 ) , .C1( u0_u11_u6_n152 ) , .ZN( u0_u11_u6_n153 ) );
  OAI211_X1 u0_u11_u6_U85 (.ZN( u0_out11_22 ) , .B( u0_u11_u6_n137 ) , .A( u0_u11_u6_n138 ) , .C2( u0_u11_u6_n139 ) , .C1( u0_u11_u6_n140 ) );
  AOI22_X1 u0_u11_u6_U86 (.B1( u0_u11_u6_n124 ) , .A2( u0_u11_u6_n125 ) , .A1( u0_u11_u6_n126 ) , .ZN( u0_u11_u6_n138 ) , .B2( u0_u11_u6_n161 ) );
  AND4_X1 u0_u11_u6_U87 (.A3( u0_u11_u6_n119 ) , .A1( u0_u11_u6_n120 ) , .A4( u0_u11_u6_n129 ) , .ZN( u0_u11_u6_n140 ) , .A2( u0_u11_u6_n143 ) );
  NAND3_X1 u0_u11_u6_U88 (.A2( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n125 ) , .A1( u0_u11_u6_n130 ) , .A3( u0_u11_u6_n131 ) );
  NAND3_X1 u0_u11_u6_U89 (.A3( u0_u11_u6_n133 ) , .ZN( u0_u11_u6_n141 ) , .A1( u0_u11_u6_n145 ) , .A2( u0_u11_u6_n148 ) );
  AOI21_X1 u0_u11_u6_U9 (.B2( u0_u11_u6_n147 ) , .B1( u0_u11_u6_n148 ) , .ZN( u0_u11_u6_n149 ) , .A( u0_u11_u6_n158 ) );
  NAND3_X1 u0_u11_u6_U90 (.ZN( u0_u11_u6_n101 ) , .A3( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n121 ) , .A1( u0_u11_u6_n127 ) );
  NAND3_X1 u0_u11_u6_U91 (.ZN( u0_u11_u6_n102 ) , .A3( u0_u11_u6_n130 ) , .A2( u0_u11_u6_n145 ) , .A1( u0_u11_u6_n166 ) );
  NAND3_X1 u0_u11_u6_U92 (.A3( u0_u11_u6_n113 ) , .A1( u0_u11_u6_n119 ) , .A2( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n93 ) );
  NAND3_X1 u0_u11_u6_U93 (.ZN( u0_u11_u6_n142 ) , .A2( u0_u11_u6_n172 ) , .A3( u0_u11_u6_n89 ) , .A1( u0_u11_u6_n90 ) );
  XOR2_X1 u0_u12_U1 (.B( u0_K13_9 ) , .A( u0_R11_6 ) , .Z( u0_u12_X_9 ) );
  XOR2_X1 u0_u12_U12 (.B( u0_K13_43 ) , .A( u0_R11_28 ) , .Z( u0_u12_X_43 ) );
  XOR2_X1 u0_u12_U14 (.B( u0_K13_41 ) , .A( u0_R11_28 ) , .Z( u0_u12_X_41 ) );
  XOR2_X1 u0_u12_U16 (.B( u0_K13_3 ) , .A( u0_R11_2 ) , .Z( u0_u12_X_3 ) );
  XOR2_X1 u0_u12_U2 (.B( u0_K13_8 ) , .A( u0_R11_5 ) , .Z( u0_u12_X_8 ) );
  XOR2_X1 u0_u12_U34 (.B( u0_K13_23 ) , .A( u0_R11_16 ) , .Z( u0_u12_X_23 ) );
  XOR2_X1 u0_u12_U35 (.B( u0_K13_22 ) , .A( u0_R11_15 ) , .Z( u0_u12_X_22 ) );
  XOR2_X1 u0_u12_U36 (.B( u0_K13_21 ) , .A( u0_R11_14 ) , .Z( u0_u12_X_21 ) );
  XOR2_X1 u0_u12_U37 (.B( u0_K13_20 ) , .A( u0_R11_13 ) , .Z( u0_u12_X_20 ) );
  XOR2_X1 u0_u12_U38 (.B( u0_K13_1 ) , .A( u0_R11_32 ) , .Z( u0_u12_X_1 ) );
  XOR2_X1 u0_u12_U39 (.B( u0_K13_19 ) , .A( u0_R11_12 ) , .Z( u0_u12_X_19 ) );
  XOR2_X1 u0_u12_U4 (.B( u0_K13_6 ) , .A( u0_R11_5 ) , .Z( u0_u12_X_6 ) );
  XOR2_X1 u0_u12_U40 (.B( u0_K13_18 ) , .A( u0_R11_13 ) , .Z( u0_u12_X_18 ) );
  XOR2_X1 u0_u12_U41 (.B( u0_K13_17 ) , .A( u0_R11_12 ) , .Z( u0_u12_X_17 ) );
  XOR2_X1 u0_u12_U42 (.B( u0_K13_16 ) , .A( u0_R11_11 ) , .Z( u0_u12_X_16 ) );
  XOR2_X1 u0_u12_U43 (.B( u0_K13_15 ) , .A( u0_R11_10 ) , .Z( u0_u12_X_15 ) );
  XOR2_X1 u0_u12_U6 (.B( u0_K13_4 ) , .A( u0_R11_3 ) , .Z( u0_u12_X_4 ) );
  XOR2_X1 u0_u12_U8 (.B( u0_K13_47 ) , .A( u0_R11_32 ) , .Z( u0_u12_X_47 ) );
  NAND2_X1 u0_u12_u0_U10 (.ZN( u0_u12_u0_n113 ) , .A1( u0_u12_u0_n139 ) , .A2( u0_u12_u0_n149 ) );
  AND3_X1 u0_u12_u0_U11 (.A2( u0_u12_u0_n112 ) , .ZN( u0_u12_u0_n127 ) , .A3( u0_u12_u0_n130 ) , .A1( u0_u12_u0_n148 ) );
  AND2_X1 u0_u12_u0_U12 (.ZN( u0_u12_u0_n107 ) , .A1( u0_u12_u0_n130 ) , .A2( u0_u12_u0_n140 ) );
  AND2_X1 u0_u12_u0_U13 (.A2( u0_u12_u0_n129 ) , .A1( u0_u12_u0_n130 ) , .ZN( u0_u12_u0_n151 ) );
  AND2_X1 u0_u12_u0_U14 (.A1( u0_u12_u0_n108 ) , .A2( u0_u12_u0_n125 ) , .ZN( u0_u12_u0_n145 ) );
  INV_X1 u0_u12_u0_U15 (.A( u0_u12_u0_n143 ) , .ZN( u0_u12_u0_n173 ) );
  NOR2_X1 u0_u12_u0_U16 (.A2( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n147 ) , .A1( u0_u12_u0_n160 ) );
  AOI21_X1 u0_u12_u0_U17 (.B1( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n132 ) , .A( u0_u12_u0_n165 ) , .B2( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U18 (.A( u0_u12_u0_n142 ) , .ZN( u0_u12_u0_n165 ) );
  OAI22_X1 u0_u12_u0_U19 (.B1( u0_u12_u0_n131 ) , .A1( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n147 ) , .A2( u0_u12_u0_n90 ) , .ZN( u0_u12_u0_n91 ) );
  AND3_X1 u0_u12_u0_U20 (.A3( u0_u12_u0_n121 ) , .A2( u0_u12_u0_n125 ) , .A1( u0_u12_u0_n148 ) , .ZN( u0_u12_u0_n90 ) );
  OAI22_X1 u0_u12_u0_U21 (.B1( u0_u12_u0_n125 ) , .ZN( u0_u12_u0_n126 ) , .A1( u0_u12_u0_n138 ) , .A2( u0_u12_u0_n146 ) , .B2( u0_u12_u0_n147 ) );
  INV_X1 u0_u12_u0_U22 (.A( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n161 ) );
  AOI22_X1 u0_u12_u0_U23 (.B2( u0_u12_u0_n109 ) , .A2( u0_u12_u0_n110 ) , .ZN( u0_u12_u0_n111 ) , .B1( u0_u12_u0_n118 ) , .A1( u0_u12_u0_n160 ) );
  NAND2_X1 u0_u12_u0_U24 (.A2( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n140 ) , .A1( u0_u12_u0_n94 ) );
  NAND2_X1 u0_u12_u0_U25 (.A2( u0_u12_u0_n102 ) , .A1( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n149 ) );
  INV_X1 u0_u12_u0_U26 (.A( u0_u12_u0_n118 ) , .ZN( u0_u12_u0_n158 ) );
  NAND2_X1 u0_u12_u0_U27 (.A2( u0_u12_u0_n100 ) , .ZN( u0_u12_u0_n131 ) , .A1( u0_u12_u0_n92 ) );
  NAND2_X1 u0_u12_u0_U28 (.ZN( u0_u12_u0_n108 ) , .A1( u0_u12_u0_n92 ) , .A2( u0_u12_u0_n94 ) );
  AOI21_X1 u0_u12_u0_U29 (.ZN( u0_u12_u0_n104 ) , .B1( u0_u12_u0_n107 ) , .B2( u0_u12_u0_n141 ) , .A( u0_u12_u0_n144 ) );
  INV_X1 u0_u12_u0_U3 (.A( u0_u12_u0_n113 ) , .ZN( u0_u12_u0_n166 ) );
  AOI21_X1 u0_u12_u0_U30 (.ZN( u0_u12_u0_n116 ) , .B2( u0_u12_u0_n142 ) , .A( u0_u12_u0_n144 ) , .B1( u0_u12_u0_n166 ) );
  AOI21_X1 u0_u12_u0_U31 (.B1( u0_u12_u0_n127 ) , .B2( u0_u12_u0_n129 ) , .A( u0_u12_u0_n138 ) , .ZN( u0_u12_u0_n96 ) );
  NAND2_X1 u0_u12_u0_U32 (.A2( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n114 ) , .A1( u0_u12_u0_n92 ) );
  NOR2_X1 u0_u12_u0_U33 (.A1( u0_u12_u0_n120 ) , .ZN( u0_u12_u0_n143 ) , .A2( u0_u12_u0_n167 ) );
  OAI221_X1 u0_u12_u0_U34 (.C1( u0_u12_u0_n112 ) , .ZN( u0_u12_u0_n120 ) , .B1( u0_u12_u0_n138 ) , .B2( u0_u12_u0_n141 ) , .C2( u0_u12_u0_n147 ) , .A( u0_u12_u0_n172 ) );
  AOI211_X1 u0_u12_u0_U35 (.B( u0_u12_u0_n115 ) , .A( u0_u12_u0_n116 ) , .C2( u0_u12_u0_n117 ) , .C1( u0_u12_u0_n118 ) , .ZN( u0_u12_u0_n119 ) );
  NAND2_X1 u0_u12_u0_U36 (.A1( u0_u12_u0_n100 ) , .A2( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n125 ) );
  NAND2_X1 u0_u12_u0_U37 (.A1( u0_u12_u0_n101 ) , .A2( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n150 ) );
  INV_X1 u0_u12_u0_U38 (.A( u0_u12_u0_n138 ) , .ZN( u0_u12_u0_n160 ) );
  NAND2_X1 u0_u12_u0_U39 (.A2( u0_u12_u0_n100 ) , .A1( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n139 ) );
  AOI21_X1 u0_u12_u0_U4 (.B1( u0_u12_u0_n114 ) , .ZN( u0_u12_u0_n115 ) , .B2( u0_u12_u0_n129 ) , .A( u0_u12_u0_n161 ) );
  NAND2_X1 u0_u12_u0_U40 (.A1( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n130 ) , .A2( u0_u12_u0_n94 ) );
  NAND2_X1 u0_u12_u0_U41 (.ZN( u0_u12_u0_n112 ) , .A2( u0_u12_u0_n92 ) , .A1( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U42 (.ZN( u0_u12_u0_n172 ) , .A( u0_u12_u0_n88 ) );
  OAI222_X1 u0_u12_u0_U43 (.C1( u0_u12_u0_n108 ) , .A1( u0_u12_u0_n125 ) , .B2( u0_u12_u0_n128 ) , .B1( u0_u12_u0_n144 ) , .A2( u0_u12_u0_n158 ) , .C2( u0_u12_u0_n161 ) , .ZN( u0_u12_u0_n88 ) );
  NAND2_X1 u0_u12_u0_U44 (.A2( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n121 ) , .A1( u0_u12_u0_n93 ) );
  OR3_X1 u0_u12_u0_U45 (.A3( u0_u12_u0_n152 ) , .A2( u0_u12_u0_n153 ) , .A1( u0_u12_u0_n154 ) , .ZN( u0_u12_u0_n155 ) );
  AOI21_X1 u0_u12_u0_U46 (.A( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n145 ) , .B1( u0_u12_u0_n146 ) , .ZN( u0_u12_u0_n154 ) );
  AOI21_X1 u0_u12_u0_U47 (.B2( u0_u12_u0_n150 ) , .B1( u0_u12_u0_n151 ) , .ZN( u0_u12_u0_n152 ) , .A( u0_u12_u0_n158 ) );
  AOI21_X1 u0_u12_u0_U48 (.A( u0_u12_u0_n147 ) , .B2( u0_u12_u0_n148 ) , .B1( u0_u12_u0_n149 ) , .ZN( u0_u12_u0_n153 ) );
  INV_X1 u0_u12_u0_U49 (.ZN( u0_u12_u0_n171 ) , .A( u0_u12_u0_n99 ) );
  AOI21_X1 u0_u12_u0_U5 (.B2( u0_u12_u0_n131 ) , .ZN( u0_u12_u0_n134 ) , .B1( u0_u12_u0_n151 ) , .A( u0_u12_u0_n158 ) );
  OAI211_X1 u0_u12_u0_U50 (.C2( u0_u12_u0_n140 ) , .C1( u0_u12_u0_n161 ) , .A( u0_u12_u0_n169 ) , .B( u0_u12_u0_n98 ) , .ZN( u0_u12_u0_n99 ) );
  INV_X1 u0_u12_u0_U51 (.ZN( u0_u12_u0_n169 ) , .A( u0_u12_u0_n91 ) );
  AOI211_X1 u0_u12_u0_U52 (.C1( u0_u12_u0_n118 ) , .A( u0_u12_u0_n123 ) , .B( u0_u12_u0_n96 ) , .C2( u0_u12_u0_n97 ) , .ZN( u0_u12_u0_n98 ) );
  NOR2_X1 u0_u12_u0_U53 (.A2( u0_u12_X_4 ) , .A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n118 ) );
  NOR2_X1 u0_u12_u0_U54 (.A2( u0_u12_X_1 ) , .ZN( u0_u12_u0_n101 ) , .A1( u0_u12_u0_n163 ) );
  NOR2_X1 u0_u12_u0_U55 (.A2( u0_u12_X_6 ) , .ZN( u0_u12_u0_n100 ) , .A1( u0_u12_u0_n162 ) );
  NAND2_X1 u0_u12_u0_U56 (.A2( u0_u12_X_4 ) , .A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n144 ) );
  NOR2_X1 u0_u12_u0_U57 (.A2( u0_u12_X_5 ) , .ZN( u0_u12_u0_n136 ) , .A1( u0_u12_u0_n159 ) );
  NAND2_X1 u0_u12_u0_U58 (.A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n138 ) , .A2( u0_u12_u0_n159 ) );
  AND2_X1 u0_u12_u0_U59 (.A2( u0_u12_X_3 ) , .A1( u0_u12_X_6 ) , .ZN( u0_u12_u0_n102 ) );
  NOR2_X1 u0_u12_u0_U6 (.A1( u0_u12_u0_n108 ) , .ZN( u0_u12_u0_n123 ) , .A2( u0_u12_u0_n158 ) );
  AND2_X1 u0_u12_u0_U60 (.A1( u0_u12_X_6 ) , .A2( u0_u12_u0_n162 ) , .ZN( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U61 (.A( u0_u12_X_4 ) , .ZN( u0_u12_u0_n159 ) );
  INV_X1 u0_u12_u0_U62 (.A( u0_u12_X_3 ) , .ZN( u0_u12_u0_n162 ) );
  INV_X1 u0_u12_u0_U63 (.A( u0_u12_u0_n126 ) , .ZN( u0_u12_u0_n168 ) );
  AOI211_X1 u0_u12_u0_U64 (.B( u0_u12_u0_n133 ) , .A( u0_u12_u0_n134 ) , .C2( u0_u12_u0_n135 ) , .C1( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n137 ) );
  OR4_X1 u0_u12_u0_U65 (.ZN( u0_out12_17 ) , .A4( u0_u12_u0_n122 ) , .A2( u0_u12_u0_n123 ) , .A1( u0_u12_u0_n124 ) , .A3( u0_u12_u0_n170 ) );
  AOI21_X1 u0_u12_u0_U66 (.B2( u0_u12_u0_n107 ) , .ZN( u0_u12_u0_n124 ) , .B1( u0_u12_u0_n128 ) , .A( u0_u12_u0_n161 ) );
  INV_X1 u0_u12_u0_U67 (.A( u0_u12_u0_n111 ) , .ZN( u0_u12_u0_n170 ) );
  OR4_X1 u0_u12_u0_U68 (.ZN( u0_out12_31 ) , .A4( u0_u12_u0_n155 ) , .A2( u0_u12_u0_n156 ) , .A1( u0_u12_u0_n157 ) , .A3( u0_u12_u0_n173 ) );
  AOI21_X1 u0_u12_u0_U69 (.A( u0_u12_u0_n138 ) , .B2( u0_u12_u0_n139 ) , .B1( u0_u12_u0_n140 ) , .ZN( u0_u12_u0_n157 ) );
  OAI21_X1 u0_u12_u0_U7 (.B1( u0_u12_u0_n150 ) , .B2( u0_u12_u0_n158 ) , .A( u0_u12_u0_n172 ) , .ZN( u0_u12_u0_n89 ) );
  AOI21_X1 u0_u12_u0_U70 (.B2( u0_u12_u0_n141 ) , .B1( u0_u12_u0_n142 ) , .ZN( u0_u12_u0_n156 ) , .A( u0_u12_u0_n161 ) );
  INV_X1 u0_u12_u0_U71 (.ZN( u0_u12_u0_n174 ) , .A( u0_u12_u0_n89 ) );
  AOI211_X1 u0_u12_u0_U72 (.B( u0_u12_u0_n104 ) , .A( u0_u12_u0_n105 ) , .ZN( u0_u12_u0_n106 ) , .C2( u0_u12_u0_n113 ) , .C1( u0_u12_u0_n160 ) );
  AND2_X1 u0_u12_u0_U73 (.A2( u0_u12_X_1 ) , .A1( u0_u12_X_2 ) , .ZN( u0_u12_u0_n95 ) );
  INV_X1 u0_u12_u0_U74 (.A( u0_u12_X_1 ) , .ZN( u0_u12_u0_n164 ) );
  NOR2_X1 u0_u12_u0_U75 (.A2( u0_u12_X_3 ) , .A1( u0_u12_X_6 ) , .ZN( u0_u12_u0_n94 ) );
  OAI221_X1 u0_u12_u0_U76 (.C1( u0_u12_u0_n121 ) , .ZN( u0_u12_u0_n122 ) , .B2( u0_u12_u0_n127 ) , .A( u0_u12_u0_n143 ) , .B1( u0_u12_u0_n144 ) , .C2( u0_u12_u0_n147 ) );
  AOI21_X1 u0_u12_u0_U77 (.B1( u0_u12_u0_n132 ) , .ZN( u0_u12_u0_n133 ) , .A( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n166 ) );
  OAI22_X1 u0_u12_u0_U78 (.ZN( u0_u12_u0_n105 ) , .A2( u0_u12_u0_n132 ) , .B1( u0_u12_u0_n146 ) , .A1( u0_u12_u0_n147 ) , .B2( u0_u12_u0_n161 ) );
  NAND2_X1 u0_u12_u0_U79 (.ZN( u0_u12_u0_n110 ) , .A2( u0_u12_u0_n132 ) , .A1( u0_u12_u0_n145 ) );
  AND2_X1 u0_u12_u0_U8 (.A1( u0_u12_u0_n114 ) , .A2( u0_u12_u0_n121 ) , .ZN( u0_u12_u0_n146 ) );
  INV_X1 u0_u12_u0_U80 (.A( u0_u12_u0_n119 ) , .ZN( u0_u12_u0_n167 ) );
  NAND2_X1 u0_u12_u0_U81 (.ZN( u0_u12_u0_n148 ) , .A1( u0_u12_u0_n93 ) , .A2( u0_u12_u0_n95 ) );
  NAND2_X1 u0_u12_u0_U82 (.A1( u0_u12_u0_n100 ) , .ZN( u0_u12_u0_n129 ) , .A2( u0_u12_u0_n95 ) );
  NAND2_X1 u0_u12_u0_U83 (.A1( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n128 ) , .A2( u0_u12_u0_n95 ) );
  NOR2_X1 u0_u12_u0_U84 (.A2( u0_u12_X_1 ) , .A1( u0_u12_X_2 ) , .ZN( u0_u12_u0_n92 ) );
  NAND2_X1 u0_u12_u0_U85 (.ZN( u0_u12_u0_n142 ) , .A1( u0_u12_u0_n94 ) , .A2( u0_u12_u0_n95 ) );
  NOR2_X1 u0_u12_u0_U86 (.A2( u0_u12_X_2 ) , .ZN( u0_u12_u0_n103 ) , .A1( u0_u12_u0_n164 ) );
  INV_X1 u0_u12_u0_U87 (.A( u0_u12_X_2 ) , .ZN( u0_u12_u0_n163 ) );
  NAND3_X1 u0_u12_u0_U88 (.ZN( u0_out12_23 ) , .A3( u0_u12_u0_n137 ) , .A1( u0_u12_u0_n168 ) , .A2( u0_u12_u0_n171 ) );
  NAND3_X1 u0_u12_u0_U89 (.A3( u0_u12_u0_n127 ) , .A2( u0_u12_u0_n128 ) , .ZN( u0_u12_u0_n135 ) , .A1( u0_u12_u0_n150 ) );
  AND2_X1 u0_u12_u0_U9 (.A1( u0_u12_u0_n131 ) , .ZN( u0_u12_u0_n141 ) , .A2( u0_u12_u0_n150 ) );
  NAND3_X1 u0_u12_u0_U90 (.ZN( u0_u12_u0_n117 ) , .A3( u0_u12_u0_n132 ) , .A2( u0_u12_u0_n139 ) , .A1( u0_u12_u0_n148 ) );
  NAND3_X1 u0_u12_u0_U91 (.ZN( u0_u12_u0_n109 ) , .A2( u0_u12_u0_n114 ) , .A3( u0_u12_u0_n140 ) , .A1( u0_u12_u0_n149 ) );
  NAND3_X1 u0_u12_u0_U92 (.ZN( u0_out12_9 ) , .A3( u0_u12_u0_n106 ) , .A2( u0_u12_u0_n171 ) , .A1( u0_u12_u0_n174 ) );
  NAND3_X1 u0_u12_u0_U93 (.A2( u0_u12_u0_n128 ) , .A1( u0_u12_u0_n132 ) , .A3( u0_u12_u0_n146 ) , .ZN( u0_u12_u0_n97 ) );
  NOR2_X1 u0_u12_u1_U10 (.A1( u0_u12_u1_n112 ) , .A2( u0_u12_u1_n116 ) , .ZN( u0_u12_u1_n118 ) );
  NAND3_X1 u0_u12_u1_U100 (.ZN( u0_u12_u1_n113 ) , .A1( u0_u12_u1_n120 ) , .A3( u0_u12_u1_n133 ) , .A2( u0_u12_u1_n155 ) );
  OAI21_X1 u0_u12_u1_U11 (.ZN( u0_u12_u1_n101 ) , .B1( u0_u12_u1_n141 ) , .A( u0_u12_u1_n146 ) , .B2( u0_u12_u1_n183 ) );
  AOI21_X1 u0_u12_u1_U12 (.B2( u0_u12_u1_n155 ) , .B1( u0_u12_u1_n156 ) , .ZN( u0_u12_u1_n157 ) , .A( u0_u12_u1_n174 ) );
  OR4_X1 u0_u12_u1_U13 (.A4( u0_u12_u1_n106 ) , .A3( u0_u12_u1_n107 ) , .ZN( u0_u12_u1_n108 ) , .A1( u0_u12_u1_n117 ) , .A2( u0_u12_u1_n184 ) );
  AOI21_X1 u0_u12_u1_U14 (.ZN( u0_u12_u1_n106 ) , .A( u0_u12_u1_n112 ) , .B1( u0_u12_u1_n154 ) , .B2( u0_u12_u1_n156 ) );
  INV_X1 u0_u12_u1_U15 (.A( u0_u12_u1_n101 ) , .ZN( u0_u12_u1_n184 ) );
  AOI21_X1 u0_u12_u1_U16 (.ZN( u0_u12_u1_n107 ) , .B1( u0_u12_u1_n134 ) , .B2( u0_u12_u1_n149 ) , .A( u0_u12_u1_n174 ) );
  NAND2_X1 u0_u12_u1_U17 (.ZN( u0_u12_u1_n140 ) , .A2( u0_u12_u1_n150 ) , .A1( u0_u12_u1_n155 ) );
  NAND2_X1 u0_u12_u1_U18 (.A1( u0_u12_u1_n131 ) , .ZN( u0_u12_u1_n147 ) , .A2( u0_u12_u1_n153 ) );
  INV_X1 u0_u12_u1_U19 (.A( u0_u12_u1_n139 ) , .ZN( u0_u12_u1_n174 ) );
  INV_X1 u0_u12_u1_U20 (.A( u0_u12_u1_n112 ) , .ZN( u0_u12_u1_n171 ) );
  NAND2_X1 u0_u12_u1_U21 (.ZN( u0_u12_u1_n141 ) , .A1( u0_u12_u1_n153 ) , .A2( u0_u12_u1_n156 ) );
  AND2_X1 u0_u12_u1_U22 (.A1( u0_u12_u1_n123 ) , .ZN( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n161 ) );
  NAND2_X1 u0_u12_u1_U23 (.A2( u0_u12_u1_n115 ) , .A1( u0_u12_u1_n116 ) , .ZN( u0_u12_u1_n148 ) );
  NAND2_X1 u0_u12_u1_U24 (.A2( u0_u12_u1_n133 ) , .A1( u0_u12_u1_n135 ) , .ZN( u0_u12_u1_n159 ) );
  NAND2_X1 u0_u12_u1_U25 (.A2( u0_u12_u1_n115 ) , .A1( u0_u12_u1_n120 ) , .ZN( u0_u12_u1_n132 ) );
  INV_X1 u0_u12_u1_U26 (.A( u0_u12_u1_n154 ) , .ZN( u0_u12_u1_n178 ) );
  INV_X1 u0_u12_u1_U27 (.A( u0_u12_u1_n151 ) , .ZN( u0_u12_u1_n183 ) );
  AND2_X1 u0_u12_u1_U28 (.A1( u0_u12_u1_n129 ) , .A2( u0_u12_u1_n133 ) , .ZN( u0_u12_u1_n149 ) );
  INV_X1 u0_u12_u1_U29 (.A( u0_u12_u1_n131 ) , .ZN( u0_u12_u1_n180 ) );
  INV_X1 u0_u12_u1_U3 (.A( u0_u12_u1_n159 ) , .ZN( u0_u12_u1_n182 ) );
  AOI221_X1 u0_u12_u1_U30 (.B1( u0_u12_u1_n140 ) , .ZN( u0_u12_u1_n167 ) , .B2( u0_u12_u1_n172 ) , .C2( u0_u12_u1_n175 ) , .C1( u0_u12_u1_n178 ) , .A( u0_u12_u1_n188 ) );
  INV_X1 u0_u12_u1_U31 (.ZN( u0_u12_u1_n188 ) , .A( u0_u12_u1_n97 ) );
  AOI211_X1 u0_u12_u1_U32 (.A( u0_u12_u1_n118 ) , .C1( u0_u12_u1_n132 ) , .C2( u0_u12_u1_n139 ) , .B( u0_u12_u1_n96 ) , .ZN( u0_u12_u1_n97 ) );
  AOI21_X1 u0_u12_u1_U33 (.B2( u0_u12_u1_n121 ) , .B1( u0_u12_u1_n135 ) , .A( u0_u12_u1_n152 ) , .ZN( u0_u12_u1_n96 ) );
  OAI221_X1 u0_u12_u1_U34 (.A( u0_u12_u1_n119 ) , .C2( u0_u12_u1_n129 ) , .ZN( u0_u12_u1_n138 ) , .B2( u0_u12_u1_n152 ) , .C1( u0_u12_u1_n174 ) , .B1( u0_u12_u1_n187 ) );
  INV_X1 u0_u12_u1_U35 (.A( u0_u12_u1_n148 ) , .ZN( u0_u12_u1_n187 ) );
  AOI211_X1 u0_u12_u1_U36 (.B( u0_u12_u1_n117 ) , .A( u0_u12_u1_n118 ) , .ZN( u0_u12_u1_n119 ) , .C2( u0_u12_u1_n146 ) , .C1( u0_u12_u1_n159 ) );
  NOR2_X1 u0_u12_u1_U37 (.A1( u0_u12_u1_n168 ) , .A2( u0_u12_u1_n176 ) , .ZN( u0_u12_u1_n98 ) );
  AOI211_X1 u0_u12_u1_U38 (.B( u0_u12_u1_n162 ) , .A( u0_u12_u1_n163 ) , .C2( u0_u12_u1_n164 ) , .ZN( u0_u12_u1_n165 ) , .C1( u0_u12_u1_n171 ) );
  AOI21_X1 u0_u12_u1_U39 (.A( u0_u12_u1_n160 ) , .B2( u0_u12_u1_n161 ) , .ZN( u0_u12_u1_n162 ) , .B1( u0_u12_u1_n182 ) );
  AOI221_X1 u0_u12_u1_U4 (.A( u0_u12_u1_n138 ) , .C2( u0_u12_u1_n139 ) , .C1( u0_u12_u1_n140 ) , .B2( u0_u12_u1_n141 ) , .ZN( u0_u12_u1_n142 ) , .B1( u0_u12_u1_n175 ) );
  OR2_X1 u0_u12_u1_U40 (.A2( u0_u12_u1_n157 ) , .A1( u0_u12_u1_n158 ) , .ZN( u0_u12_u1_n163 ) );
  NAND2_X1 u0_u12_u1_U41 (.A1( u0_u12_u1_n128 ) , .ZN( u0_u12_u1_n146 ) , .A2( u0_u12_u1_n160 ) );
  NAND2_X1 u0_u12_u1_U42 (.A2( u0_u12_u1_n112 ) , .ZN( u0_u12_u1_n139 ) , .A1( u0_u12_u1_n152 ) );
  NAND2_X1 u0_u12_u1_U43 (.A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n156 ) , .A2( u0_u12_u1_n99 ) );
  NOR2_X1 u0_u12_u1_U44 (.ZN( u0_u12_u1_n117 ) , .A1( u0_u12_u1_n121 ) , .A2( u0_u12_u1_n160 ) );
  OAI21_X1 u0_u12_u1_U45 (.B2( u0_u12_u1_n123 ) , .ZN( u0_u12_u1_n145 ) , .B1( u0_u12_u1_n160 ) , .A( u0_u12_u1_n185 ) );
  INV_X1 u0_u12_u1_U46 (.A( u0_u12_u1_n122 ) , .ZN( u0_u12_u1_n185 ) );
  AOI21_X1 u0_u12_u1_U47 (.B2( u0_u12_u1_n120 ) , .B1( u0_u12_u1_n121 ) , .ZN( u0_u12_u1_n122 ) , .A( u0_u12_u1_n128 ) );
  AOI21_X1 u0_u12_u1_U48 (.A( u0_u12_u1_n128 ) , .B2( u0_u12_u1_n129 ) , .ZN( u0_u12_u1_n130 ) , .B1( u0_u12_u1_n150 ) );
  NAND2_X1 u0_u12_u1_U49 (.ZN( u0_u12_u1_n112 ) , .A1( u0_u12_u1_n169 ) , .A2( u0_u12_u1_n170 ) );
  AOI211_X1 u0_u12_u1_U5 (.ZN( u0_u12_u1_n124 ) , .A( u0_u12_u1_n138 ) , .C2( u0_u12_u1_n139 ) , .B( u0_u12_u1_n145 ) , .C1( u0_u12_u1_n147 ) );
  NAND2_X1 u0_u12_u1_U50 (.ZN( u0_u12_u1_n129 ) , .A2( u0_u12_u1_n95 ) , .A1( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U51 (.A1( u0_u12_u1_n102 ) , .ZN( u0_u12_u1_n154 ) , .A2( u0_u12_u1_n99 ) );
  NAND2_X1 u0_u12_u1_U52 (.A2( u0_u12_u1_n100 ) , .ZN( u0_u12_u1_n135 ) , .A1( u0_u12_u1_n99 ) );
  AOI21_X1 u0_u12_u1_U53 (.A( u0_u12_u1_n152 ) , .B2( u0_u12_u1_n153 ) , .B1( u0_u12_u1_n154 ) , .ZN( u0_u12_u1_n158 ) );
  INV_X1 u0_u12_u1_U54 (.A( u0_u12_u1_n160 ) , .ZN( u0_u12_u1_n175 ) );
  NAND2_X1 u0_u12_u1_U55 (.A1( u0_u12_u1_n100 ) , .ZN( u0_u12_u1_n116 ) , .A2( u0_u12_u1_n95 ) );
  NAND2_X1 u0_u12_u1_U56 (.A1( u0_u12_u1_n102 ) , .ZN( u0_u12_u1_n131 ) , .A2( u0_u12_u1_n95 ) );
  NAND2_X1 u0_u12_u1_U57 (.A2( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n121 ) , .A1( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U58 (.A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n153 ) , .A2( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U59 (.A2( u0_u12_u1_n104 ) , .A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n133 ) );
  AOI22_X1 u0_u12_u1_U6 (.B2( u0_u12_u1_n113 ) , .A2( u0_u12_u1_n114 ) , .ZN( u0_u12_u1_n125 ) , .A1( u0_u12_u1_n171 ) , .B1( u0_u12_u1_n173 ) );
  NAND2_X1 u0_u12_u1_U60 (.ZN( u0_u12_u1_n150 ) , .A2( u0_u12_u1_n98 ) , .A1( u0_u12_u1_n99 ) );
  NAND2_X1 u0_u12_u1_U61 (.A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n155 ) , .A2( u0_u12_u1_n95 ) );
  OAI21_X1 u0_u12_u1_U62 (.ZN( u0_u12_u1_n109 ) , .B1( u0_u12_u1_n129 ) , .B2( u0_u12_u1_n160 ) , .A( u0_u12_u1_n167 ) );
  NAND2_X1 u0_u12_u1_U63 (.A2( u0_u12_u1_n100 ) , .A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n120 ) );
  NAND2_X1 u0_u12_u1_U64 (.A1( u0_u12_u1_n102 ) , .A2( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n115 ) );
  NAND2_X1 u0_u12_u1_U65 (.A2( u0_u12_u1_n100 ) , .A1( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n151 ) );
  NAND2_X1 u0_u12_u1_U66 (.A2( u0_u12_u1_n103 ) , .A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n161 ) );
  INV_X1 u0_u12_u1_U67 (.A( u0_u12_u1_n152 ) , .ZN( u0_u12_u1_n173 ) );
  INV_X1 u0_u12_u1_U68 (.A( u0_u12_u1_n128 ) , .ZN( u0_u12_u1_n172 ) );
  NAND2_X1 u0_u12_u1_U69 (.A2( u0_u12_u1_n102 ) , .A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n123 ) );
  NAND2_X1 u0_u12_u1_U7 (.ZN( u0_u12_u1_n114 ) , .A1( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n156 ) );
  NOR2_X1 u0_u12_u1_U70 (.A2( u0_u12_X_7 ) , .A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n95 ) );
  NOR2_X1 u0_u12_u1_U71 (.A1( u0_u12_X_12 ) , .A2( u0_u12_X_9 ) , .ZN( u0_u12_u1_n100 ) );
  NOR2_X1 u0_u12_u1_U72 (.A2( u0_u12_X_8 ) , .A1( u0_u12_u1_n177 ) , .ZN( u0_u12_u1_n99 ) );
  NOR2_X1 u0_u12_u1_U73 (.A2( u0_u12_X_12 ) , .ZN( u0_u12_u1_n102 ) , .A1( u0_u12_u1_n176 ) );
  NOR2_X1 u0_u12_u1_U74 (.A2( u0_u12_X_9 ) , .ZN( u0_u12_u1_n105 ) , .A1( u0_u12_u1_n168 ) );
  NAND2_X1 u0_u12_u1_U75 (.A1( u0_u12_X_10 ) , .ZN( u0_u12_u1_n160 ) , .A2( u0_u12_u1_n169 ) );
  NAND2_X1 u0_u12_u1_U76 (.A2( u0_u12_X_10 ) , .A1( u0_u12_X_11 ) , .ZN( u0_u12_u1_n152 ) );
  NAND2_X1 u0_u12_u1_U77 (.A1( u0_u12_X_11 ) , .ZN( u0_u12_u1_n128 ) , .A2( u0_u12_u1_n170 ) );
  AND2_X1 u0_u12_u1_U78 (.A2( u0_u12_X_7 ) , .A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n104 ) );
  AND2_X1 u0_u12_u1_U79 (.A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n103 ) , .A2( u0_u12_u1_n177 ) );
  AOI22_X1 u0_u12_u1_U8 (.B2( u0_u12_u1_n136 ) , .A2( u0_u12_u1_n137 ) , .ZN( u0_u12_u1_n143 ) , .A1( u0_u12_u1_n171 ) , .B1( u0_u12_u1_n173 ) );
  INV_X1 u0_u12_u1_U80 (.A( u0_u12_X_10 ) , .ZN( u0_u12_u1_n170 ) );
  INV_X1 u0_u12_u1_U81 (.A( u0_u12_X_9 ) , .ZN( u0_u12_u1_n176 ) );
  INV_X1 u0_u12_u1_U82 (.A( u0_u12_X_11 ) , .ZN( u0_u12_u1_n169 ) );
  INV_X1 u0_u12_u1_U83 (.A( u0_u12_X_12 ) , .ZN( u0_u12_u1_n168 ) );
  INV_X1 u0_u12_u1_U84 (.A( u0_u12_X_7 ) , .ZN( u0_u12_u1_n177 ) );
  NAND4_X1 u0_u12_u1_U85 (.ZN( u0_out12_28 ) , .A4( u0_u12_u1_n124 ) , .A3( u0_u12_u1_n125 ) , .A2( u0_u12_u1_n126 ) , .A1( u0_u12_u1_n127 ) );
  OAI21_X1 u0_u12_u1_U86 (.ZN( u0_u12_u1_n127 ) , .B2( u0_u12_u1_n139 ) , .B1( u0_u12_u1_n175 ) , .A( u0_u12_u1_n183 ) );
  OAI21_X1 u0_u12_u1_U87 (.ZN( u0_u12_u1_n126 ) , .B2( u0_u12_u1_n140 ) , .A( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n178 ) );
  NAND4_X1 u0_u12_u1_U88 (.ZN( u0_out12_18 ) , .A4( u0_u12_u1_n165 ) , .A3( u0_u12_u1_n166 ) , .A1( u0_u12_u1_n167 ) , .A2( u0_u12_u1_n186 ) );
  AOI22_X1 u0_u12_u1_U89 (.B2( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n147 ) , .A2( u0_u12_u1_n148 ) , .ZN( u0_u12_u1_n166 ) , .A1( u0_u12_u1_n172 ) );
  INV_X1 u0_u12_u1_U9 (.A( u0_u12_u1_n147 ) , .ZN( u0_u12_u1_n181 ) );
  INV_X1 u0_u12_u1_U90 (.A( u0_u12_u1_n145 ) , .ZN( u0_u12_u1_n186 ) );
  NAND4_X1 u0_u12_u1_U91 (.ZN( u0_out12_2 ) , .A4( u0_u12_u1_n142 ) , .A3( u0_u12_u1_n143 ) , .A2( u0_u12_u1_n144 ) , .A1( u0_u12_u1_n179 ) );
  OAI21_X1 u0_u12_u1_U92 (.B2( u0_u12_u1_n132 ) , .ZN( u0_u12_u1_n144 ) , .A( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n180 ) );
  INV_X1 u0_u12_u1_U93 (.A( u0_u12_u1_n130 ) , .ZN( u0_u12_u1_n179 ) );
  OR4_X1 u0_u12_u1_U94 (.ZN( u0_out12_13 ) , .A4( u0_u12_u1_n108 ) , .A3( u0_u12_u1_n109 ) , .A2( u0_u12_u1_n110 ) , .A1( u0_u12_u1_n111 ) );
  AOI21_X1 u0_u12_u1_U95 (.ZN( u0_u12_u1_n111 ) , .A( u0_u12_u1_n128 ) , .B2( u0_u12_u1_n131 ) , .B1( u0_u12_u1_n135 ) );
  AOI21_X1 u0_u12_u1_U96 (.ZN( u0_u12_u1_n110 ) , .A( u0_u12_u1_n116 ) , .B1( u0_u12_u1_n152 ) , .B2( u0_u12_u1_n160 ) );
  NAND3_X1 u0_u12_u1_U97 (.A3( u0_u12_u1_n149 ) , .A2( u0_u12_u1_n150 ) , .A1( u0_u12_u1_n151 ) , .ZN( u0_u12_u1_n164 ) );
  NAND3_X1 u0_u12_u1_U98 (.A3( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n135 ) , .ZN( u0_u12_u1_n136 ) , .A1( u0_u12_u1_n151 ) );
  NAND3_X1 u0_u12_u1_U99 (.A1( u0_u12_u1_n133 ) , .ZN( u0_u12_u1_n137 ) , .A2( u0_u12_u1_n154 ) , .A3( u0_u12_u1_n181 ) );
  OAI22_X1 u0_u12_u2_U10 (.B1( u0_u12_u2_n151 ) , .A2( u0_u12_u2_n152 ) , .A1( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n160 ) , .B2( u0_u12_u2_n168 ) );
  NAND3_X1 u0_u12_u2_U100 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n104 ) , .A3( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n98 ) );
  NOR3_X1 u0_u12_u2_U11 (.A1( u0_u12_u2_n150 ) , .ZN( u0_u12_u2_n151 ) , .A3( u0_u12_u2_n175 ) , .A2( u0_u12_u2_n188 ) );
  AOI21_X1 u0_u12_u2_U12 (.B2( u0_u12_u2_n123 ) , .ZN( u0_u12_u2_n125 ) , .A( u0_u12_u2_n171 ) , .B1( u0_u12_u2_n184 ) );
  INV_X1 u0_u12_u2_U13 (.A( u0_u12_u2_n150 ) , .ZN( u0_u12_u2_n184 ) );
  AOI21_X1 u0_u12_u2_U14 (.ZN( u0_u12_u2_n144 ) , .B2( u0_u12_u2_n155 ) , .A( u0_u12_u2_n172 ) , .B1( u0_u12_u2_n185 ) );
  AOI21_X1 u0_u12_u2_U15 (.B2( u0_u12_u2_n143 ) , .ZN( u0_u12_u2_n145 ) , .B1( u0_u12_u2_n152 ) , .A( u0_u12_u2_n171 ) );
  INV_X1 u0_u12_u2_U16 (.A( u0_u12_u2_n156 ) , .ZN( u0_u12_u2_n171 ) );
  INV_X1 u0_u12_u2_U17 (.A( u0_u12_u2_n120 ) , .ZN( u0_u12_u2_n188 ) );
  NAND2_X1 u0_u12_u2_U18 (.A2( u0_u12_u2_n122 ) , .ZN( u0_u12_u2_n150 ) , .A1( u0_u12_u2_n152 ) );
  INV_X1 u0_u12_u2_U19 (.A( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n170 ) );
  INV_X1 u0_u12_u2_U20 (.A( u0_u12_u2_n137 ) , .ZN( u0_u12_u2_n173 ) );
  NAND2_X1 u0_u12_u2_U21 (.A1( u0_u12_u2_n132 ) , .A2( u0_u12_u2_n139 ) , .ZN( u0_u12_u2_n157 ) );
  INV_X1 u0_u12_u2_U22 (.A( u0_u12_u2_n113 ) , .ZN( u0_u12_u2_n178 ) );
  INV_X1 u0_u12_u2_U23 (.A( u0_u12_u2_n139 ) , .ZN( u0_u12_u2_n175 ) );
  INV_X1 u0_u12_u2_U24 (.A( u0_u12_u2_n155 ) , .ZN( u0_u12_u2_n181 ) );
  INV_X1 u0_u12_u2_U25 (.A( u0_u12_u2_n119 ) , .ZN( u0_u12_u2_n177 ) );
  INV_X1 u0_u12_u2_U26 (.A( u0_u12_u2_n116 ) , .ZN( u0_u12_u2_n180 ) );
  INV_X1 u0_u12_u2_U27 (.A( u0_u12_u2_n131 ) , .ZN( u0_u12_u2_n179 ) );
  INV_X1 u0_u12_u2_U28 (.A( u0_u12_u2_n154 ) , .ZN( u0_u12_u2_n176 ) );
  NAND2_X1 u0_u12_u2_U29 (.A2( u0_u12_u2_n116 ) , .A1( u0_u12_u2_n117 ) , .ZN( u0_u12_u2_n118 ) );
  NOR2_X1 u0_u12_u2_U3 (.ZN( u0_u12_u2_n121 ) , .A2( u0_u12_u2_n177 ) , .A1( u0_u12_u2_n180 ) );
  INV_X1 u0_u12_u2_U30 (.A( u0_u12_u2_n132 ) , .ZN( u0_u12_u2_n182 ) );
  INV_X1 u0_u12_u2_U31 (.A( u0_u12_u2_n158 ) , .ZN( u0_u12_u2_n183 ) );
  OAI21_X1 u0_u12_u2_U32 (.A( u0_u12_u2_n156 ) , .B1( u0_u12_u2_n157 ) , .ZN( u0_u12_u2_n158 ) , .B2( u0_u12_u2_n179 ) );
  NOR2_X1 u0_u12_u2_U33 (.ZN( u0_u12_u2_n156 ) , .A1( u0_u12_u2_n166 ) , .A2( u0_u12_u2_n169 ) );
  NOR2_X1 u0_u12_u2_U34 (.A2( u0_u12_u2_n114 ) , .ZN( u0_u12_u2_n137 ) , .A1( u0_u12_u2_n140 ) );
  NOR2_X1 u0_u12_u2_U35 (.A2( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n153 ) , .A1( u0_u12_u2_n156 ) );
  AOI211_X1 u0_u12_u2_U36 (.ZN( u0_u12_u2_n130 ) , .C1( u0_u12_u2_n138 ) , .C2( u0_u12_u2_n179 ) , .B( u0_u12_u2_n96 ) , .A( u0_u12_u2_n97 ) );
  OAI22_X1 u0_u12_u2_U37 (.B1( u0_u12_u2_n133 ) , .A2( u0_u12_u2_n137 ) , .A1( u0_u12_u2_n152 ) , .B2( u0_u12_u2_n168 ) , .ZN( u0_u12_u2_n97 ) );
  OAI221_X1 u0_u12_u2_U38 (.B1( u0_u12_u2_n113 ) , .C1( u0_u12_u2_n132 ) , .A( u0_u12_u2_n149 ) , .B2( u0_u12_u2_n171 ) , .C2( u0_u12_u2_n172 ) , .ZN( u0_u12_u2_n96 ) );
  OAI221_X1 u0_u12_u2_U39 (.A( u0_u12_u2_n115 ) , .C2( u0_u12_u2_n123 ) , .B2( u0_u12_u2_n143 ) , .B1( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n163 ) , .C1( u0_u12_u2_n168 ) );
  INV_X1 u0_u12_u2_U4 (.A( u0_u12_u2_n134 ) , .ZN( u0_u12_u2_n185 ) );
  OAI21_X1 u0_u12_u2_U40 (.A( u0_u12_u2_n114 ) , .ZN( u0_u12_u2_n115 ) , .B1( u0_u12_u2_n176 ) , .B2( u0_u12_u2_n178 ) );
  OAI221_X1 u0_u12_u2_U41 (.A( u0_u12_u2_n135 ) , .B2( u0_u12_u2_n136 ) , .B1( u0_u12_u2_n137 ) , .ZN( u0_u12_u2_n162 ) , .C2( u0_u12_u2_n167 ) , .C1( u0_u12_u2_n185 ) );
  AND3_X1 u0_u12_u2_U42 (.A3( u0_u12_u2_n131 ) , .A2( u0_u12_u2_n132 ) , .A1( u0_u12_u2_n133 ) , .ZN( u0_u12_u2_n136 ) );
  AOI22_X1 u0_u12_u2_U43 (.ZN( u0_u12_u2_n135 ) , .B1( u0_u12_u2_n140 ) , .A1( u0_u12_u2_n156 ) , .B2( u0_u12_u2_n180 ) , .A2( u0_u12_u2_n188 ) );
  AOI21_X1 u0_u12_u2_U44 (.ZN( u0_u12_u2_n149 ) , .B1( u0_u12_u2_n173 ) , .B2( u0_u12_u2_n188 ) , .A( u0_u12_u2_n95 ) );
  AND3_X1 u0_u12_u2_U45 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n104 ) , .A3( u0_u12_u2_n156 ) , .ZN( u0_u12_u2_n95 ) );
  OAI21_X1 u0_u12_u2_U46 (.A( u0_u12_u2_n101 ) , .B2( u0_u12_u2_n121 ) , .B1( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n164 ) );
  NAND2_X1 u0_u12_u2_U47 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n107 ) , .ZN( u0_u12_u2_n155 ) );
  NAND2_X1 u0_u12_u2_U48 (.A2( u0_u12_u2_n105 ) , .A1( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n143 ) );
  NAND2_X1 u0_u12_u2_U49 (.A1( u0_u12_u2_n104 ) , .A2( u0_u12_u2_n106 ) , .ZN( u0_u12_u2_n152 ) );
  NOR4_X1 u0_u12_u2_U5 (.A4( u0_u12_u2_n124 ) , .A3( u0_u12_u2_n125 ) , .A2( u0_u12_u2_n126 ) , .A1( u0_u12_u2_n127 ) , .ZN( u0_u12_u2_n128 ) );
  NAND2_X1 u0_u12_u2_U50 (.A1( u0_u12_u2_n100 ) , .A2( u0_u12_u2_n105 ) , .ZN( u0_u12_u2_n132 ) );
  INV_X1 u0_u12_u2_U51 (.A( u0_u12_u2_n140 ) , .ZN( u0_u12_u2_n168 ) );
  INV_X1 u0_u12_u2_U52 (.A( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n167 ) );
  OAI21_X1 u0_u12_u2_U53 (.A( u0_u12_u2_n141 ) , .B2( u0_u12_u2_n142 ) , .ZN( u0_u12_u2_n146 ) , .B1( u0_u12_u2_n153 ) );
  OAI21_X1 u0_u12_u2_U54 (.A( u0_u12_u2_n140 ) , .ZN( u0_u12_u2_n141 ) , .B1( u0_u12_u2_n176 ) , .B2( u0_u12_u2_n177 ) );
  NOR3_X1 u0_u12_u2_U55 (.ZN( u0_u12_u2_n142 ) , .A3( u0_u12_u2_n175 ) , .A2( u0_u12_u2_n178 ) , .A1( u0_u12_u2_n181 ) );
  NAND2_X1 u0_u12_u2_U56 (.A1( u0_u12_u2_n102 ) , .A2( u0_u12_u2_n106 ) , .ZN( u0_u12_u2_n113 ) );
  NAND2_X1 u0_u12_u2_U57 (.A1( u0_u12_u2_n106 ) , .A2( u0_u12_u2_n107 ) , .ZN( u0_u12_u2_n131 ) );
  NAND2_X1 u0_u12_u2_U58 (.A1( u0_u12_u2_n103 ) , .A2( u0_u12_u2_n107 ) , .ZN( u0_u12_u2_n139 ) );
  NAND2_X1 u0_u12_u2_U59 (.A1( u0_u12_u2_n103 ) , .A2( u0_u12_u2_n105 ) , .ZN( u0_u12_u2_n133 ) );
  AOI21_X1 u0_u12_u2_U6 (.B2( u0_u12_u2_n119 ) , .ZN( u0_u12_u2_n127 ) , .A( u0_u12_u2_n137 ) , .B1( u0_u12_u2_n155 ) );
  NAND2_X1 u0_u12_u2_U60 (.A1( u0_u12_u2_n102 ) , .A2( u0_u12_u2_n103 ) , .ZN( u0_u12_u2_n154 ) );
  NAND2_X1 u0_u12_u2_U61 (.A2( u0_u12_u2_n103 ) , .A1( u0_u12_u2_n104 ) , .ZN( u0_u12_u2_n119 ) );
  NAND2_X1 u0_u12_u2_U62 (.A2( u0_u12_u2_n107 ) , .A1( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n123 ) );
  NAND2_X1 u0_u12_u2_U63 (.A1( u0_u12_u2_n104 ) , .A2( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n122 ) );
  INV_X1 u0_u12_u2_U64 (.A( u0_u12_u2_n114 ) , .ZN( u0_u12_u2_n172 ) );
  NAND2_X1 u0_u12_u2_U65 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n102 ) , .ZN( u0_u12_u2_n116 ) );
  NAND2_X1 u0_u12_u2_U66 (.A1( u0_u12_u2_n102 ) , .A2( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n120 ) );
  NAND2_X1 u0_u12_u2_U67 (.A2( u0_u12_u2_n105 ) , .A1( u0_u12_u2_n106 ) , .ZN( u0_u12_u2_n117 ) );
  INV_X1 u0_u12_u2_U68 (.ZN( u0_u12_u2_n187 ) , .A( u0_u12_u2_n99 ) );
  OAI21_X1 u0_u12_u2_U69 (.B1( u0_u12_u2_n137 ) , .B2( u0_u12_u2_n143 ) , .A( u0_u12_u2_n98 ) , .ZN( u0_u12_u2_n99 ) );
  AOI21_X1 u0_u12_u2_U7 (.ZN( u0_u12_u2_n124 ) , .B1( u0_u12_u2_n131 ) , .B2( u0_u12_u2_n143 ) , .A( u0_u12_u2_n172 ) );
  NOR2_X1 u0_u12_u2_U70 (.A2( u0_u12_X_16 ) , .ZN( u0_u12_u2_n140 ) , .A1( u0_u12_u2_n166 ) );
  NOR2_X1 u0_u12_u2_U71 (.A2( u0_u12_X_13 ) , .A1( u0_u12_X_14 ) , .ZN( u0_u12_u2_n100 ) );
  NOR2_X1 u0_u12_u2_U72 (.A2( u0_u12_X_16 ) , .A1( u0_u12_X_17 ) , .ZN( u0_u12_u2_n138 ) );
  NOR2_X1 u0_u12_u2_U73 (.A2( u0_u12_X_15 ) , .A1( u0_u12_X_18 ) , .ZN( u0_u12_u2_n104 ) );
  NOR2_X1 u0_u12_u2_U74 (.A2( u0_u12_X_14 ) , .ZN( u0_u12_u2_n103 ) , .A1( u0_u12_u2_n174 ) );
  NOR2_X1 u0_u12_u2_U75 (.A2( u0_u12_X_15 ) , .ZN( u0_u12_u2_n102 ) , .A1( u0_u12_u2_n165 ) );
  NOR2_X1 u0_u12_u2_U76 (.A2( u0_u12_X_17 ) , .ZN( u0_u12_u2_n114 ) , .A1( u0_u12_u2_n169 ) );
  AND2_X1 u0_u12_u2_U77 (.A1( u0_u12_X_15 ) , .ZN( u0_u12_u2_n105 ) , .A2( u0_u12_u2_n165 ) );
  AND2_X1 u0_u12_u2_U78 (.A2( u0_u12_X_15 ) , .A1( u0_u12_X_18 ) , .ZN( u0_u12_u2_n107 ) );
  AND2_X1 u0_u12_u2_U79 (.A1( u0_u12_X_14 ) , .ZN( u0_u12_u2_n106 ) , .A2( u0_u12_u2_n174 ) );
  AOI21_X1 u0_u12_u2_U8 (.B2( u0_u12_u2_n120 ) , .B1( u0_u12_u2_n121 ) , .ZN( u0_u12_u2_n126 ) , .A( u0_u12_u2_n167 ) );
  AND2_X1 u0_u12_u2_U80 (.A1( u0_u12_X_13 ) , .A2( u0_u12_X_14 ) , .ZN( u0_u12_u2_n108 ) );
  INV_X1 u0_u12_u2_U81 (.A( u0_u12_X_16 ) , .ZN( u0_u12_u2_n169 ) );
  INV_X1 u0_u12_u2_U82 (.A( u0_u12_X_17 ) , .ZN( u0_u12_u2_n166 ) );
  INV_X1 u0_u12_u2_U83 (.A( u0_u12_X_13 ) , .ZN( u0_u12_u2_n174 ) );
  INV_X1 u0_u12_u2_U84 (.A( u0_u12_X_18 ) , .ZN( u0_u12_u2_n165 ) );
  NAND4_X1 u0_u12_u2_U85 (.ZN( u0_out12_30 ) , .A4( u0_u12_u2_n147 ) , .A3( u0_u12_u2_n148 ) , .A2( u0_u12_u2_n149 ) , .A1( u0_u12_u2_n187 ) );
  AOI21_X1 u0_u12_u2_U86 (.B2( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n148 ) , .A( u0_u12_u2_n162 ) , .B1( u0_u12_u2_n182 ) );
  NOR3_X1 u0_u12_u2_U87 (.A3( u0_u12_u2_n144 ) , .A2( u0_u12_u2_n145 ) , .A1( u0_u12_u2_n146 ) , .ZN( u0_u12_u2_n147 ) );
  NAND4_X1 u0_u12_u2_U88 (.ZN( u0_out12_24 ) , .A4( u0_u12_u2_n111 ) , .A3( u0_u12_u2_n112 ) , .A1( u0_u12_u2_n130 ) , .A2( u0_u12_u2_n187 ) );
  AOI221_X1 u0_u12_u2_U89 (.A( u0_u12_u2_n109 ) , .B1( u0_u12_u2_n110 ) , .ZN( u0_u12_u2_n111 ) , .C1( u0_u12_u2_n134 ) , .C2( u0_u12_u2_n170 ) , .B2( u0_u12_u2_n173 ) );
  OAI22_X1 u0_u12_u2_U9 (.ZN( u0_u12_u2_n109 ) , .A2( u0_u12_u2_n113 ) , .B2( u0_u12_u2_n133 ) , .B1( u0_u12_u2_n167 ) , .A1( u0_u12_u2_n168 ) );
  AOI21_X1 u0_u12_u2_U90 (.ZN( u0_u12_u2_n112 ) , .B2( u0_u12_u2_n156 ) , .A( u0_u12_u2_n164 ) , .B1( u0_u12_u2_n181 ) );
  NAND4_X1 u0_u12_u2_U91 (.ZN( u0_out12_16 ) , .A4( u0_u12_u2_n128 ) , .A3( u0_u12_u2_n129 ) , .A1( u0_u12_u2_n130 ) , .A2( u0_u12_u2_n186 ) );
  AOI22_X1 u0_u12_u2_U92 (.A2( u0_u12_u2_n118 ) , .ZN( u0_u12_u2_n129 ) , .A1( u0_u12_u2_n140 ) , .B1( u0_u12_u2_n157 ) , .B2( u0_u12_u2_n170 ) );
  INV_X1 u0_u12_u2_U93 (.A( u0_u12_u2_n163 ) , .ZN( u0_u12_u2_n186 ) );
  OR4_X1 u0_u12_u2_U94 (.ZN( u0_out12_6 ) , .A4( u0_u12_u2_n161 ) , .A3( u0_u12_u2_n162 ) , .A2( u0_u12_u2_n163 ) , .A1( u0_u12_u2_n164 ) );
  OR3_X1 u0_u12_u2_U95 (.A2( u0_u12_u2_n159 ) , .A1( u0_u12_u2_n160 ) , .ZN( u0_u12_u2_n161 ) , .A3( u0_u12_u2_n183 ) );
  AOI21_X1 u0_u12_u2_U96 (.B2( u0_u12_u2_n154 ) , .B1( u0_u12_u2_n155 ) , .ZN( u0_u12_u2_n159 ) , .A( u0_u12_u2_n167 ) );
  NAND3_X1 u0_u12_u2_U97 (.A2( u0_u12_u2_n117 ) , .A1( u0_u12_u2_n122 ) , .A3( u0_u12_u2_n123 ) , .ZN( u0_u12_u2_n134 ) );
  NAND3_X1 u0_u12_u2_U98 (.ZN( u0_u12_u2_n110 ) , .A2( u0_u12_u2_n131 ) , .A3( u0_u12_u2_n139 ) , .A1( u0_u12_u2_n154 ) );
  NAND3_X1 u0_u12_u2_U99 (.A2( u0_u12_u2_n100 ) , .ZN( u0_u12_u2_n101 ) , .A1( u0_u12_u2_n104 ) , .A3( u0_u12_u2_n114 ) );
  OAI22_X1 u0_u12_u3_U10 (.B1( u0_u12_u3_n113 ) , .A2( u0_u12_u3_n135 ) , .A1( u0_u12_u3_n150 ) , .B2( u0_u12_u3_n164 ) , .ZN( u0_u12_u3_n98 ) );
  OAI211_X1 u0_u12_u3_U11 (.B( u0_u12_u3_n106 ) , .ZN( u0_u12_u3_n119 ) , .C2( u0_u12_u3_n128 ) , .C1( u0_u12_u3_n167 ) , .A( u0_u12_u3_n181 ) );
  AOI221_X1 u0_u12_u3_U12 (.C1( u0_u12_u3_n105 ) , .ZN( u0_u12_u3_n106 ) , .A( u0_u12_u3_n131 ) , .B2( u0_u12_u3_n132 ) , .C2( u0_u12_u3_n133 ) , .B1( u0_u12_u3_n169 ) );
  INV_X1 u0_u12_u3_U13 (.ZN( u0_u12_u3_n181 ) , .A( u0_u12_u3_n98 ) );
  NAND2_X1 u0_u12_u3_U14 (.ZN( u0_u12_u3_n105 ) , .A2( u0_u12_u3_n130 ) , .A1( u0_u12_u3_n155 ) );
  AOI22_X1 u0_u12_u3_U15 (.B1( u0_u12_u3_n115 ) , .A2( u0_u12_u3_n116 ) , .ZN( u0_u12_u3_n123 ) , .B2( u0_u12_u3_n133 ) , .A1( u0_u12_u3_n169 ) );
  NAND2_X1 u0_u12_u3_U16 (.ZN( u0_u12_u3_n116 ) , .A2( u0_u12_u3_n151 ) , .A1( u0_u12_u3_n182 ) );
  NOR2_X1 u0_u12_u3_U17 (.ZN( u0_u12_u3_n126 ) , .A2( u0_u12_u3_n150 ) , .A1( u0_u12_u3_n164 ) );
  AOI21_X1 u0_u12_u3_U18 (.ZN( u0_u12_u3_n112 ) , .B2( u0_u12_u3_n146 ) , .B1( u0_u12_u3_n155 ) , .A( u0_u12_u3_n167 ) );
  NAND2_X1 u0_u12_u3_U19 (.A1( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n142 ) , .A2( u0_u12_u3_n164 ) );
  NAND2_X1 u0_u12_u3_U20 (.ZN( u0_u12_u3_n132 ) , .A2( u0_u12_u3_n152 ) , .A1( u0_u12_u3_n156 ) );
  AND2_X1 u0_u12_u3_U21 (.A2( u0_u12_u3_n113 ) , .A1( u0_u12_u3_n114 ) , .ZN( u0_u12_u3_n151 ) );
  INV_X1 u0_u12_u3_U22 (.A( u0_u12_u3_n133 ) , .ZN( u0_u12_u3_n165 ) );
  INV_X1 u0_u12_u3_U23 (.A( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n170 ) );
  NAND2_X1 u0_u12_u3_U24 (.A1( u0_u12_u3_n107 ) , .A2( u0_u12_u3_n108 ) , .ZN( u0_u12_u3_n140 ) );
  NAND2_X1 u0_u12_u3_U25 (.ZN( u0_u12_u3_n117 ) , .A1( u0_u12_u3_n124 ) , .A2( u0_u12_u3_n148 ) );
  NAND2_X1 u0_u12_u3_U26 (.ZN( u0_u12_u3_n143 ) , .A1( u0_u12_u3_n165 ) , .A2( u0_u12_u3_n167 ) );
  INV_X1 u0_u12_u3_U27 (.A( u0_u12_u3_n130 ) , .ZN( u0_u12_u3_n177 ) );
  INV_X1 u0_u12_u3_U28 (.A( u0_u12_u3_n128 ) , .ZN( u0_u12_u3_n176 ) );
  INV_X1 u0_u12_u3_U29 (.A( u0_u12_u3_n155 ) , .ZN( u0_u12_u3_n174 ) );
  INV_X1 u0_u12_u3_U3 (.A( u0_u12_u3_n129 ) , .ZN( u0_u12_u3_n183 ) );
  INV_X1 u0_u12_u3_U30 (.A( u0_u12_u3_n139 ) , .ZN( u0_u12_u3_n185 ) );
  NOR2_X1 u0_u12_u3_U31 (.ZN( u0_u12_u3_n135 ) , .A2( u0_u12_u3_n141 ) , .A1( u0_u12_u3_n169 ) );
  OAI222_X1 u0_u12_u3_U32 (.C2( u0_u12_u3_n107 ) , .A2( u0_u12_u3_n108 ) , .B1( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n138 ) , .B2( u0_u12_u3_n146 ) , .C1( u0_u12_u3_n154 ) , .A1( u0_u12_u3_n164 ) );
  NOR4_X1 u0_u12_u3_U33 (.A4( u0_u12_u3_n157 ) , .A3( u0_u12_u3_n158 ) , .A2( u0_u12_u3_n159 ) , .A1( u0_u12_u3_n160 ) , .ZN( u0_u12_u3_n161 ) );
  AOI21_X1 u0_u12_u3_U34 (.B2( u0_u12_u3_n152 ) , .B1( u0_u12_u3_n153 ) , .ZN( u0_u12_u3_n158 ) , .A( u0_u12_u3_n164 ) );
  AOI21_X1 u0_u12_u3_U35 (.A( u0_u12_u3_n154 ) , .B2( u0_u12_u3_n155 ) , .B1( u0_u12_u3_n156 ) , .ZN( u0_u12_u3_n157 ) );
  AOI21_X1 u0_u12_u3_U36 (.A( u0_u12_u3_n149 ) , .B2( u0_u12_u3_n150 ) , .B1( u0_u12_u3_n151 ) , .ZN( u0_u12_u3_n159 ) );
  AOI211_X1 u0_u12_u3_U37 (.ZN( u0_u12_u3_n109 ) , .A( u0_u12_u3_n119 ) , .C2( u0_u12_u3_n129 ) , .B( u0_u12_u3_n138 ) , .C1( u0_u12_u3_n141 ) );
  AOI211_X1 u0_u12_u3_U38 (.B( u0_u12_u3_n119 ) , .A( u0_u12_u3_n120 ) , .C2( u0_u12_u3_n121 ) , .ZN( u0_u12_u3_n122 ) , .C1( u0_u12_u3_n179 ) );
  INV_X1 u0_u12_u3_U39 (.A( u0_u12_u3_n156 ) , .ZN( u0_u12_u3_n179 ) );
  INV_X1 u0_u12_u3_U4 (.A( u0_u12_u3_n140 ) , .ZN( u0_u12_u3_n182 ) );
  OAI22_X1 u0_u12_u3_U40 (.B1( u0_u12_u3_n118 ) , .ZN( u0_u12_u3_n120 ) , .A1( u0_u12_u3_n135 ) , .B2( u0_u12_u3_n154 ) , .A2( u0_u12_u3_n178 ) );
  AND3_X1 u0_u12_u3_U41 (.ZN( u0_u12_u3_n118 ) , .A2( u0_u12_u3_n124 ) , .A1( u0_u12_u3_n144 ) , .A3( u0_u12_u3_n152 ) );
  INV_X1 u0_u12_u3_U42 (.A( u0_u12_u3_n121 ) , .ZN( u0_u12_u3_n164 ) );
  NAND2_X1 u0_u12_u3_U43 (.ZN( u0_u12_u3_n133 ) , .A1( u0_u12_u3_n154 ) , .A2( u0_u12_u3_n164 ) );
  OAI211_X1 u0_u12_u3_U44 (.B( u0_u12_u3_n127 ) , .ZN( u0_u12_u3_n139 ) , .C1( u0_u12_u3_n150 ) , .C2( u0_u12_u3_n154 ) , .A( u0_u12_u3_n184 ) );
  INV_X1 u0_u12_u3_U45 (.A( u0_u12_u3_n125 ) , .ZN( u0_u12_u3_n184 ) );
  AOI221_X1 u0_u12_u3_U46 (.A( u0_u12_u3_n126 ) , .ZN( u0_u12_u3_n127 ) , .C2( u0_u12_u3_n132 ) , .C1( u0_u12_u3_n169 ) , .B2( u0_u12_u3_n170 ) , .B1( u0_u12_u3_n174 ) );
  OAI22_X1 u0_u12_u3_U47 (.A1( u0_u12_u3_n124 ) , .ZN( u0_u12_u3_n125 ) , .B2( u0_u12_u3_n145 ) , .A2( u0_u12_u3_n165 ) , .B1( u0_u12_u3_n167 ) );
  NOR2_X1 u0_u12_u3_U48 (.A1( u0_u12_u3_n113 ) , .ZN( u0_u12_u3_n131 ) , .A2( u0_u12_u3_n154 ) );
  NAND2_X1 u0_u12_u3_U49 (.A1( u0_u12_u3_n103 ) , .ZN( u0_u12_u3_n150 ) , .A2( u0_u12_u3_n99 ) );
  INV_X1 u0_u12_u3_U5 (.A( u0_u12_u3_n117 ) , .ZN( u0_u12_u3_n178 ) );
  NAND2_X1 u0_u12_u3_U50 (.A2( u0_u12_u3_n102 ) , .ZN( u0_u12_u3_n155 ) , .A1( u0_u12_u3_n97 ) );
  INV_X1 u0_u12_u3_U51 (.A( u0_u12_u3_n141 ) , .ZN( u0_u12_u3_n167 ) );
  AOI21_X1 u0_u12_u3_U52 (.B2( u0_u12_u3_n114 ) , .B1( u0_u12_u3_n146 ) , .A( u0_u12_u3_n154 ) , .ZN( u0_u12_u3_n94 ) );
  AOI21_X1 u0_u12_u3_U53 (.ZN( u0_u12_u3_n110 ) , .B2( u0_u12_u3_n142 ) , .B1( u0_u12_u3_n186 ) , .A( u0_u12_u3_n95 ) );
  INV_X1 u0_u12_u3_U54 (.A( u0_u12_u3_n145 ) , .ZN( u0_u12_u3_n186 ) );
  AOI21_X1 u0_u12_u3_U55 (.B1( u0_u12_u3_n124 ) , .A( u0_u12_u3_n149 ) , .B2( u0_u12_u3_n155 ) , .ZN( u0_u12_u3_n95 ) );
  INV_X1 u0_u12_u3_U56 (.A( u0_u12_u3_n149 ) , .ZN( u0_u12_u3_n169 ) );
  NAND2_X1 u0_u12_u3_U57 (.ZN( u0_u12_u3_n124 ) , .A1( u0_u12_u3_n96 ) , .A2( u0_u12_u3_n97 ) );
  NAND2_X1 u0_u12_u3_U58 (.A2( u0_u12_u3_n100 ) , .ZN( u0_u12_u3_n146 ) , .A1( u0_u12_u3_n96 ) );
  NAND2_X1 u0_u12_u3_U59 (.A1( u0_u12_u3_n101 ) , .ZN( u0_u12_u3_n145 ) , .A2( u0_u12_u3_n99 ) );
  AOI221_X1 u0_u12_u3_U6 (.A( u0_u12_u3_n131 ) , .C2( u0_u12_u3_n132 ) , .C1( u0_u12_u3_n133 ) , .ZN( u0_u12_u3_n134 ) , .B1( u0_u12_u3_n143 ) , .B2( u0_u12_u3_n177 ) );
  NAND2_X1 u0_u12_u3_U60 (.A1( u0_u12_u3_n100 ) , .ZN( u0_u12_u3_n156 ) , .A2( u0_u12_u3_n99 ) );
  NAND2_X1 u0_u12_u3_U61 (.A2( u0_u12_u3_n101 ) , .A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n148 ) );
  NAND2_X1 u0_u12_u3_U62 (.A1( u0_u12_u3_n100 ) , .A2( u0_u12_u3_n102 ) , .ZN( u0_u12_u3_n128 ) );
  NAND2_X1 u0_u12_u3_U63 (.A2( u0_u12_u3_n101 ) , .A1( u0_u12_u3_n102 ) , .ZN( u0_u12_u3_n152 ) );
  NAND2_X1 u0_u12_u3_U64 (.A2( u0_u12_u3_n101 ) , .ZN( u0_u12_u3_n114 ) , .A1( u0_u12_u3_n96 ) );
  NAND2_X1 u0_u12_u3_U65 (.ZN( u0_u12_u3_n107 ) , .A1( u0_u12_u3_n97 ) , .A2( u0_u12_u3_n99 ) );
  NAND2_X1 u0_u12_u3_U66 (.A2( u0_u12_u3_n100 ) , .A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n113 ) );
  NAND2_X1 u0_u12_u3_U67 (.A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n153 ) , .A2( u0_u12_u3_n97 ) );
  NAND2_X1 u0_u12_u3_U68 (.A2( u0_u12_u3_n103 ) , .A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n130 ) );
  NAND2_X1 u0_u12_u3_U69 (.A2( u0_u12_u3_n103 ) , .ZN( u0_u12_u3_n144 ) , .A1( u0_u12_u3_n96 ) );
  OAI22_X1 u0_u12_u3_U7 (.B2( u0_u12_u3_n147 ) , .A2( u0_u12_u3_n148 ) , .ZN( u0_u12_u3_n160 ) , .B1( u0_u12_u3_n165 ) , .A1( u0_u12_u3_n168 ) );
  NAND2_X1 u0_u12_u3_U70 (.A1( u0_u12_u3_n102 ) , .A2( u0_u12_u3_n103 ) , .ZN( u0_u12_u3_n108 ) );
  NOR2_X1 u0_u12_u3_U71 (.A2( u0_u12_X_19 ) , .A1( u0_u12_X_20 ) , .ZN( u0_u12_u3_n99 ) );
  NOR2_X1 u0_u12_u3_U72 (.A2( u0_u12_X_21 ) , .A1( u0_u12_X_24 ) , .ZN( u0_u12_u3_n103 ) );
  NOR2_X1 u0_u12_u3_U73 (.A2( u0_u12_X_24 ) , .A1( u0_u12_u3_n171 ) , .ZN( u0_u12_u3_n97 ) );
  NOR2_X1 u0_u12_u3_U74 (.A2( u0_u12_X_23 ) , .ZN( u0_u12_u3_n141 ) , .A1( u0_u12_u3_n166 ) );
  NOR2_X1 u0_u12_u3_U75 (.A2( u0_u12_X_19 ) , .A1( u0_u12_u3_n172 ) , .ZN( u0_u12_u3_n96 ) );
  NAND2_X1 u0_u12_u3_U76 (.A1( u0_u12_X_22 ) , .A2( u0_u12_X_23 ) , .ZN( u0_u12_u3_n154 ) );
  NAND2_X1 u0_u12_u3_U77 (.A1( u0_u12_X_23 ) , .ZN( u0_u12_u3_n149 ) , .A2( u0_u12_u3_n166 ) );
  NOR2_X1 u0_u12_u3_U78 (.A2( u0_u12_X_22 ) , .A1( u0_u12_X_23 ) , .ZN( u0_u12_u3_n121 ) );
  AND2_X1 u0_u12_u3_U79 (.A1( u0_u12_X_24 ) , .ZN( u0_u12_u3_n101 ) , .A2( u0_u12_u3_n171 ) );
  AND3_X1 u0_u12_u3_U8 (.A3( u0_u12_u3_n144 ) , .A2( u0_u12_u3_n145 ) , .A1( u0_u12_u3_n146 ) , .ZN( u0_u12_u3_n147 ) );
  AND2_X1 u0_u12_u3_U80 (.A1( u0_u12_X_19 ) , .ZN( u0_u12_u3_n102 ) , .A2( u0_u12_u3_n172 ) );
  AND2_X1 u0_u12_u3_U81 (.A1( u0_u12_X_21 ) , .A2( u0_u12_X_24 ) , .ZN( u0_u12_u3_n100 ) );
  AND2_X1 u0_u12_u3_U82 (.A2( u0_u12_X_19 ) , .A1( u0_u12_X_20 ) , .ZN( u0_u12_u3_n104 ) );
  INV_X1 u0_u12_u3_U83 (.A( u0_u12_X_22 ) , .ZN( u0_u12_u3_n166 ) );
  INV_X1 u0_u12_u3_U84 (.A( u0_u12_X_21 ) , .ZN( u0_u12_u3_n171 ) );
  INV_X1 u0_u12_u3_U85 (.A( u0_u12_X_20 ) , .ZN( u0_u12_u3_n172 ) );
  OR4_X1 u0_u12_u3_U86 (.ZN( u0_out12_10 ) , .A4( u0_u12_u3_n136 ) , .A3( u0_u12_u3_n137 ) , .A1( u0_u12_u3_n138 ) , .A2( u0_u12_u3_n139 ) );
  OAI222_X1 u0_u12_u3_U87 (.C1( u0_u12_u3_n128 ) , .ZN( u0_u12_u3_n137 ) , .B1( u0_u12_u3_n148 ) , .A2( u0_u12_u3_n150 ) , .B2( u0_u12_u3_n154 ) , .C2( u0_u12_u3_n164 ) , .A1( u0_u12_u3_n167 ) );
  OAI221_X1 u0_u12_u3_U88 (.A( u0_u12_u3_n134 ) , .B2( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n136 ) , .C1( u0_u12_u3_n149 ) , .B1( u0_u12_u3_n151 ) , .C2( u0_u12_u3_n183 ) );
  NAND4_X1 u0_u12_u3_U89 (.ZN( u0_out12_26 ) , .A4( u0_u12_u3_n109 ) , .A3( u0_u12_u3_n110 ) , .A2( u0_u12_u3_n111 ) , .A1( u0_u12_u3_n173 ) );
  INV_X1 u0_u12_u3_U9 (.A( u0_u12_u3_n143 ) , .ZN( u0_u12_u3_n168 ) );
  INV_X1 u0_u12_u3_U90 (.ZN( u0_u12_u3_n173 ) , .A( u0_u12_u3_n94 ) );
  OAI21_X1 u0_u12_u3_U91 (.ZN( u0_u12_u3_n111 ) , .B2( u0_u12_u3_n117 ) , .A( u0_u12_u3_n133 ) , .B1( u0_u12_u3_n176 ) );
  NAND4_X1 u0_u12_u3_U92 (.ZN( u0_out12_20 ) , .A4( u0_u12_u3_n122 ) , .A3( u0_u12_u3_n123 ) , .A1( u0_u12_u3_n175 ) , .A2( u0_u12_u3_n180 ) );
  INV_X1 u0_u12_u3_U93 (.A( u0_u12_u3_n126 ) , .ZN( u0_u12_u3_n180 ) );
  INV_X1 u0_u12_u3_U94 (.A( u0_u12_u3_n112 ) , .ZN( u0_u12_u3_n175 ) );
  NAND4_X1 u0_u12_u3_U95 (.ZN( u0_out12_1 ) , .A4( u0_u12_u3_n161 ) , .A3( u0_u12_u3_n162 ) , .A2( u0_u12_u3_n163 ) , .A1( u0_u12_u3_n185 ) );
  NAND2_X1 u0_u12_u3_U96 (.ZN( u0_u12_u3_n163 ) , .A2( u0_u12_u3_n170 ) , .A1( u0_u12_u3_n176 ) );
  AOI22_X1 u0_u12_u3_U97 (.B2( u0_u12_u3_n140 ) , .B1( u0_u12_u3_n141 ) , .A2( u0_u12_u3_n142 ) , .ZN( u0_u12_u3_n162 ) , .A1( u0_u12_u3_n177 ) );
  NAND3_X1 u0_u12_u3_U98 (.A1( u0_u12_u3_n114 ) , .ZN( u0_u12_u3_n115 ) , .A2( u0_u12_u3_n145 ) , .A3( u0_u12_u3_n153 ) );
  NAND3_X1 u0_u12_u3_U99 (.ZN( u0_u12_u3_n129 ) , .A2( u0_u12_u3_n144 ) , .A1( u0_u12_u3_n153 ) , .A3( u0_u12_u3_n182 ) );
  AOI22_X1 u0_u12_u6_U10 (.A2( u0_u12_u6_n151 ) , .B2( u0_u12_u6_n161 ) , .A1( u0_u12_u6_n167 ) , .B1( u0_u12_u6_n170 ) , .ZN( u0_u12_u6_n89 ) );
  AOI21_X1 u0_u12_u6_U11 (.B1( u0_u12_u6_n107 ) , .B2( u0_u12_u6_n132 ) , .A( u0_u12_u6_n158 ) , .ZN( u0_u12_u6_n88 ) );
  AOI21_X1 u0_u12_u6_U12 (.B2( u0_u12_u6_n147 ) , .B1( u0_u12_u6_n148 ) , .ZN( u0_u12_u6_n149 ) , .A( u0_u12_u6_n158 ) );
  AOI21_X1 u0_u12_u6_U13 (.ZN( u0_u12_u6_n106 ) , .A( u0_u12_u6_n142 ) , .B2( u0_u12_u6_n159 ) , .B1( u0_u12_u6_n164 ) );
  INV_X1 u0_u12_u6_U14 (.A( u0_u12_u6_n155 ) , .ZN( u0_u12_u6_n161 ) );
  INV_X1 u0_u12_u6_U15 (.A( u0_u12_u6_n128 ) , .ZN( u0_u12_u6_n164 ) );
  NAND2_X1 u0_u12_u6_U16 (.ZN( u0_u12_u6_n110 ) , .A1( u0_u12_u6_n122 ) , .A2( u0_u12_u6_n129 ) );
  NAND2_X1 u0_u12_u6_U17 (.ZN( u0_u12_u6_n124 ) , .A2( u0_u12_u6_n146 ) , .A1( u0_u12_u6_n148 ) );
  INV_X1 u0_u12_u6_U18 (.A( u0_u12_u6_n132 ) , .ZN( u0_u12_u6_n171 ) );
  AND2_X1 u0_u12_u6_U19 (.A1( u0_u12_u6_n100 ) , .ZN( u0_u12_u6_n130 ) , .A2( u0_u12_u6_n147 ) );
  INV_X1 u0_u12_u6_U20 (.A( u0_u12_u6_n127 ) , .ZN( u0_u12_u6_n173 ) );
  INV_X1 u0_u12_u6_U21 (.A( u0_u12_u6_n121 ) , .ZN( u0_u12_u6_n167 ) );
  INV_X1 u0_u12_u6_U22 (.A( u0_u12_u6_n100 ) , .ZN( u0_u12_u6_n169 ) );
  INV_X1 u0_u12_u6_U23 (.A( u0_u12_u6_n123 ) , .ZN( u0_u12_u6_n170 ) );
  INV_X1 u0_u12_u6_U24 (.A( u0_u12_u6_n113 ) , .ZN( u0_u12_u6_n168 ) );
  AND2_X1 u0_u12_u6_U25 (.A1( u0_u12_u6_n107 ) , .A2( u0_u12_u6_n119 ) , .ZN( u0_u12_u6_n133 ) );
  AND2_X1 u0_u12_u6_U26 (.A2( u0_u12_u6_n121 ) , .A1( u0_u12_u6_n122 ) , .ZN( u0_u12_u6_n131 ) );
  AND3_X1 u0_u12_u6_U27 (.ZN( u0_u12_u6_n120 ) , .A2( u0_u12_u6_n127 ) , .A1( u0_u12_u6_n132 ) , .A3( u0_u12_u6_n145 ) );
  INV_X1 u0_u12_u6_U28 (.A( u0_u12_u6_n146 ) , .ZN( u0_u12_u6_n163 ) );
  AOI222_X1 u0_u12_u6_U29 (.ZN( u0_u12_u6_n114 ) , .A1( u0_u12_u6_n118 ) , .A2( u0_u12_u6_n126 ) , .B2( u0_u12_u6_n151 ) , .C2( u0_u12_u6_n159 ) , .C1( u0_u12_u6_n168 ) , .B1( u0_u12_u6_n169 ) );
  INV_X1 u0_u12_u6_U3 (.A( u0_u12_u6_n110 ) , .ZN( u0_u12_u6_n166 ) );
  NOR2_X1 u0_u12_u6_U30 (.A1( u0_u12_u6_n162 ) , .A2( u0_u12_u6_n165 ) , .ZN( u0_u12_u6_n98 ) );
  AOI211_X1 u0_u12_u6_U31 (.B( u0_u12_u6_n134 ) , .A( u0_u12_u6_n135 ) , .C1( u0_u12_u6_n136 ) , .ZN( u0_u12_u6_n137 ) , .C2( u0_u12_u6_n151 ) );
  AOI21_X1 u0_u12_u6_U32 (.B2( u0_u12_u6_n132 ) , .B1( u0_u12_u6_n133 ) , .ZN( u0_u12_u6_n134 ) , .A( u0_u12_u6_n158 ) );
  AOI21_X1 u0_u12_u6_U33 (.B1( u0_u12_u6_n131 ) , .ZN( u0_u12_u6_n135 ) , .A( u0_u12_u6_n144 ) , .B2( u0_u12_u6_n146 ) );
  NAND4_X1 u0_u12_u6_U34 (.A4( u0_u12_u6_n127 ) , .A3( u0_u12_u6_n128 ) , .A2( u0_u12_u6_n129 ) , .A1( u0_u12_u6_n130 ) , .ZN( u0_u12_u6_n136 ) );
  NAND2_X1 u0_u12_u6_U35 (.A1( u0_u12_u6_n144 ) , .ZN( u0_u12_u6_n151 ) , .A2( u0_u12_u6_n158 ) );
  NAND2_X1 u0_u12_u6_U36 (.ZN( u0_u12_u6_n132 ) , .A1( u0_u12_u6_n91 ) , .A2( u0_u12_u6_n97 ) );
  AOI22_X1 u0_u12_u6_U37 (.B2( u0_u12_u6_n110 ) , .B1( u0_u12_u6_n111 ) , .A1( u0_u12_u6_n112 ) , .ZN( u0_u12_u6_n115 ) , .A2( u0_u12_u6_n161 ) );
  NAND4_X1 u0_u12_u6_U38 (.A3( u0_u12_u6_n109 ) , .ZN( u0_u12_u6_n112 ) , .A4( u0_u12_u6_n132 ) , .A2( u0_u12_u6_n147 ) , .A1( u0_u12_u6_n166 ) );
  NOR2_X1 u0_u12_u6_U39 (.ZN( u0_u12_u6_n109 ) , .A1( u0_u12_u6_n170 ) , .A2( u0_u12_u6_n173 ) );
  INV_X1 u0_u12_u6_U4 (.A( u0_u12_u6_n142 ) , .ZN( u0_u12_u6_n174 ) );
  NOR2_X1 u0_u12_u6_U40 (.A2( u0_u12_u6_n126 ) , .ZN( u0_u12_u6_n155 ) , .A1( u0_u12_u6_n160 ) );
  NAND2_X1 u0_u12_u6_U41 (.ZN( u0_u12_u6_n146 ) , .A2( u0_u12_u6_n94 ) , .A1( u0_u12_u6_n99 ) );
  AOI21_X1 u0_u12_u6_U42 (.A( u0_u12_u6_n144 ) , .B2( u0_u12_u6_n145 ) , .B1( u0_u12_u6_n146 ) , .ZN( u0_u12_u6_n150 ) );
  INV_X1 u0_u12_u6_U43 (.A( u0_u12_u6_n111 ) , .ZN( u0_u12_u6_n158 ) );
  NAND2_X1 u0_u12_u6_U44 (.ZN( u0_u12_u6_n127 ) , .A1( u0_u12_u6_n91 ) , .A2( u0_u12_u6_n92 ) );
  NAND2_X1 u0_u12_u6_U45 (.ZN( u0_u12_u6_n129 ) , .A2( u0_u12_u6_n95 ) , .A1( u0_u12_u6_n96 ) );
  INV_X1 u0_u12_u6_U46 (.A( u0_u12_u6_n144 ) , .ZN( u0_u12_u6_n159 ) );
  NAND2_X1 u0_u12_u6_U47 (.ZN( u0_u12_u6_n145 ) , .A2( u0_u12_u6_n97 ) , .A1( u0_u12_u6_n98 ) );
  NAND2_X1 u0_u12_u6_U48 (.ZN( u0_u12_u6_n148 ) , .A2( u0_u12_u6_n92 ) , .A1( u0_u12_u6_n94 ) );
  NAND2_X1 u0_u12_u6_U49 (.ZN( u0_u12_u6_n108 ) , .A2( u0_u12_u6_n139 ) , .A1( u0_u12_u6_n144 ) );
  NAND2_X1 u0_u12_u6_U5 (.A2( u0_u12_u6_n143 ) , .ZN( u0_u12_u6_n152 ) , .A1( u0_u12_u6_n166 ) );
  NAND2_X1 u0_u12_u6_U50 (.ZN( u0_u12_u6_n121 ) , .A2( u0_u12_u6_n95 ) , .A1( u0_u12_u6_n97 ) );
  NAND2_X1 u0_u12_u6_U51 (.ZN( u0_u12_u6_n107 ) , .A2( u0_u12_u6_n92 ) , .A1( u0_u12_u6_n95 ) );
  AND2_X1 u0_u12_u6_U52 (.ZN( u0_u12_u6_n118 ) , .A2( u0_u12_u6_n91 ) , .A1( u0_u12_u6_n99 ) );
  NAND2_X1 u0_u12_u6_U53 (.ZN( u0_u12_u6_n147 ) , .A2( u0_u12_u6_n98 ) , .A1( u0_u12_u6_n99 ) );
  NAND2_X1 u0_u12_u6_U54 (.ZN( u0_u12_u6_n128 ) , .A1( u0_u12_u6_n94 ) , .A2( u0_u12_u6_n96 ) );
  NAND2_X1 u0_u12_u6_U55 (.ZN( u0_u12_u6_n119 ) , .A2( u0_u12_u6_n95 ) , .A1( u0_u12_u6_n99 ) );
  NAND2_X1 u0_u12_u6_U56 (.ZN( u0_u12_u6_n123 ) , .A2( u0_u12_u6_n91 ) , .A1( u0_u12_u6_n96 ) );
  NAND2_X1 u0_u12_u6_U57 (.ZN( u0_u12_u6_n100 ) , .A2( u0_u12_u6_n92 ) , .A1( u0_u12_u6_n98 ) );
  NAND2_X1 u0_u12_u6_U58 (.ZN( u0_u12_u6_n122 ) , .A1( u0_u12_u6_n94 ) , .A2( u0_u12_u6_n97 ) );
  INV_X1 u0_u12_u6_U59 (.A( u0_u12_u6_n139 ) , .ZN( u0_u12_u6_n160 ) );
  AOI22_X1 u0_u12_u6_U6 (.B2( u0_u12_u6_n101 ) , .A1( u0_u12_u6_n102 ) , .ZN( u0_u12_u6_n103 ) , .B1( u0_u12_u6_n160 ) , .A2( u0_u12_u6_n161 ) );
  NAND2_X1 u0_u12_u6_U60 (.ZN( u0_u12_u6_n113 ) , .A1( u0_u12_u6_n96 ) , .A2( u0_u12_u6_n98 ) );
  NOR2_X1 u0_u12_u6_U61 (.A2( u0_u12_X_40 ) , .A1( u0_u12_X_41 ) , .ZN( u0_u12_u6_n126 ) );
  NOR2_X1 u0_u12_u6_U62 (.A2( u0_u12_X_39 ) , .A1( u0_u12_X_42 ) , .ZN( u0_u12_u6_n92 ) );
  NOR2_X1 u0_u12_u6_U63 (.A2( u0_u12_X_39 ) , .A1( u0_u12_u6_n156 ) , .ZN( u0_u12_u6_n97 ) );
  NOR2_X1 u0_u12_u6_U64 (.A2( u0_u12_X_38 ) , .A1( u0_u12_u6_n165 ) , .ZN( u0_u12_u6_n95 ) );
  NOR2_X1 u0_u12_u6_U65 (.A2( u0_u12_X_41 ) , .ZN( u0_u12_u6_n111 ) , .A1( u0_u12_u6_n157 ) );
  NOR2_X1 u0_u12_u6_U66 (.A2( u0_u12_X_37 ) , .A1( u0_u12_u6_n162 ) , .ZN( u0_u12_u6_n94 ) );
  NOR2_X1 u0_u12_u6_U67 (.A2( u0_u12_X_37 ) , .A1( u0_u12_X_38 ) , .ZN( u0_u12_u6_n91 ) );
  NAND2_X1 u0_u12_u6_U68 (.A1( u0_u12_X_41 ) , .ZN( u0_u12_u6_n144 ) , .A2( u0_u12_u6_n157 ) );
  NAND2_X1 u0_u12_u6_U69 (.A2( u0_u12_X_40 ) , .A1( u0_u12_X_41 ) , .ZN( u0_u12_u6_n139 ) );
  NOR2_X1 u0_u12_u6_U7 (.A1( u0_u12_u6_n118 ) , .ZN( u0_u12_u6_n143 ) , .A2( u0_u12_u6_n168 ) );
  AND2_X1 u0_u12_u6_U70 (.A1( u0_u12_X_39 ) , .A2( u0_u12_u6_n156 ) , .ZN( u0_u12_u6_n96 ) );
  AND2_X1 u0_u12_u6_U71 (.A1( u0_u12_X_39 ) , .A2( u0_u12_X_42 ) , .ZN( u0_u12_u6_n99 ) );
  INV_X1 u0_u12_u6_U72 (.A( u0_u12_X_40 ) , .ZN( u0_u12_u6_n157 ) );
  INV_X1 u0_u12_u6_U73 (.A( u0_u12_X_37 ) , .ZN( u0_u12_u6_n165 ) );
  INV_X1 u0_u12_u6_U74 (.A( u0_u12_X_38 ) , .ZN( u0_u12_u6_n162 ) );
  INV_X1 u0_u12_u6_U75 (.A( u0_u12_X_42 ) , .ZN( u0_u12_u6_n156 ) );
  NAND4_X1 u0_u12_u6_U76 (.ZN( u0_out12_32 ) , .A4( u0_u12_u6_n103 ) , .A3( u0_u12_u6_n104 ) , .A2( u0_u12_u6_n105 ) , .A1( u0_u12_u6_n106 ) );
  AOI22_X1 u0_u12_u6_U77 (.ZN( u0_u12_u6_n105 ) , .A2( u0_u12_u6_n108 ) , .A1( u0_u12_u6_n118 ) , .B2( u0_u12_u6_n126 ) , .B1( u0_u12_u6_n171 ) );
  AOI22_X1 u0_u12_u6_U78 (.ZN( u0_u12_u6_n104 ) , .A1( u0_u12_u6_n111 ) , .B1( u0_u12_u6_n124 ) , .B2( u0_u12_u6_n151 ) , .A2( u0_u12_u6_n93 ) );
  NAND4_X1 u0_u12_u6_U79 (.ZN( u0_out12_12 ) , .A4( u0_u12_u6_n114 ) , .A3( u0_u12_u6_n115 ) , .A2( u0_u12_u6_n116 ) , .A1( u0_u12_u6_n117 ) );
  INV_X1 u0_u12_u6_U8 (.ZN( u0_u12_u6_n172 ) , .A( u0_u12_u6_n88 ) );
  OAI22_X1 u0_u12_u6_U80 (.B2( u0_u12_u6_n111 ) , .ZN( u0_u12_u6_n116 ) , .B1( u0_u12_u6_n126 ) , .A2( u0_u12_u6_n164 ) , .A1( u0_u12_u6_n167 ) );
  OAI21_X1 u0_u12_u6_U81 (.A( u0_u12_u6_n108 ) , .ZN( u0_u12_u6_n117 ) , .B2( u0_u12_u6_n141 ) , .B1( u0_u12_u6_n163 ) );
  OAI211_X1 u0_u12_u6_U82 (.ZN( u0_out12_22 ) , .B( u0_u12_u6_n137 ) , .A( u0_u12_u6_n138 ) , .C2( u0_u12_u6_n139 ) , .C1( u0_u12_u6_n140 ) );
  AOI22_X1 u0_u12_u6_U83 (.B1( u0_u12_u6_n124 ) , .A2( u0_u12_u6_n125 ) , .A1( u0_u12_u6_n126 ) , .ZN( u0_u12_u6_n138 ) , .B2( u0_u12_u6_n161 ) );
  AND4_X1 u0_u12_u6_U84 (.A3( u0_u12_u6_n119 ) , .A1( u0_u12_u6_n120 ) , .A4( u0_u12_u6_n129 ) , .ZN( u0_u12_u6_n140 ) , .A2( u0_u12_u6_n143 ) );
  OAI211_X1 u0_u12_u6_U85 (.ZN( u0_out12_7 ) , .B( u0_u12_u6_n153 ) , .C2( u0_u12_u6_n154 ) , .C1( u0_u12_u6_n155 ) , .A( u0_u12_u6_n174 ) );
  NOR3_X1 u0_u12_u6_U86 (.A1( u0_u12_u6_n141 ) , .ZN( u0_u12_u6_n154 ) , .A3( u0_u12_u6_n164 ) , .A2( u0_u12_u6_n171 ) );
  AOI211_X1 u0_u12_u6_U87 (.B( u0_u12_u6_n149 ) , .A( u0_u12_u6_n150 ) , .C2( u0_u12_u6_n151 ) , .C1( u0_u12_u6_n152 ) , .ZN( u0_u12_u6_n153 ) );
  NAND3_X1 u0_u12_u6_U88 (.A2( u0_u12_u6_n123 ) , .ZN( u0_u12_u6_n125 ) , .A1( u0_u12_u6_n130 ) , .A3( u0_u12_u6_n131 ) );
  NAND3_X1 u0_u12_u6_U89 (.A3( u0_u12_u6_n133 ) , .ZN( u0_u12_u6_n141 ) , .A1( u0_u12_u6_n145 ) , .A2( u0_u12_u6_n148 ) );
  OAI21_X1 u0_u12_u6_U9 (.A( u0_u12_u6_n159 ) , .B1( u0_u12_u6_n169 ) , .B2( u0_u12_u6_n173 ) , .ZN( u0_u12_u6_n90 ) );
  NAND3_X1 u0_u12_u6_U90 (.ZN( u0_u12_u6_n101 ) , .A3( u0_u12_u6_n107 ) , .A2( u0_u12_u6_n121 ) , .A1( u0_u12_u6_n127 ) );
  NAND3_X1 u0_u12_u6_U91 (.ZN( u0_u12_u6_n102 ) , .A3( u0_u12_u6_n130 ) , .A2( u0_u12_u6_n145 ) , .A1( u0_u12_u6_n166 ) );
  NAND3_X1 u0_u12_u6_U92 (.A3( u0_u12_u6_n113 ) , .A1( u0_u12_u6_n119 ) , .A2( u0_u12_u6_n123 ) , .ZN( u0_u12_u6_n93 ) );
  NAND3_X1 u0_u12_u6_U93 (.ZN( u0_u12_u6_n142 ) , .A2( u0_u12_u6_n172 ) , .A3( u0_u12_u6_n89 ) , .A1( u0_u12_u6_n90 ) );
  AND3_X1 u0_u12_u7_U10 (.A3( u0_u12_u7_n110 ) , .A2( u0_u12_u7_n127 ) , .A1( u0_u12_u7_n132 ) , .ZN( u0_u12_u7_n92 ) );
  OAI21_X1 u0_u12_u7_U11 (.A( u0_u12_u7_n161 ) , .B1( u0_u12_u7_n168 ) , .B2( u0_u12_u7_n173 ) , .ZN( u0_u12_u7_n91 ) );
  AOI211_X1 u0_u12_u7_U12 (.A( u0_u12_u7_n117 ) , .ZN( u0_u12_u7_n118 ) , .C2( u0_u12_u7_n126 ) , .C1( u0_u12_u7_n177 ) , .B( u0_u12_u7_n180 ) );
  OAI22_X1 u0_u12_u7_U13 (.B1( u0_u12_u7_n115 ) , .ZN( u0_u12_u7_n117 ) , .A2( u0_u12_u7_n133 ) , .A1( u0_u12_u7_n137 ) , .B2( u0_u12_u7_n162 ) );
  INV_X1 u0_u12_u7_U14 (.A( u0_u12_u7_n116 ) , .ZN( u0_u12_u7_n180 ) );
  NOR3_X1 u0_u12_u7_U15 (.ZN( u0_u12_u7_n115 ) , .A3( u0_u12_u7_n145 ) , .A2( u0_u12_u7_n168 ) , .A1( u0_u12_u7_n169 ) );
  OAI211_X1 u0_u12_u7_U16 (.B( u0_u12_u7_n122 ) , .A( u0_u12_u7_n123 ) , .C2( u0_u12_u7_n124 ) , .ZN( u0_u12_u7_n154 ) , .C1( u0_u12_u7_n162 ) );
  AOI222_X1 u0_u12_u7_U17 (.ZN( u0_u12_u7_n122 ) , .C2( u0_u12_u7_n126 ) , .C1( u0_u12_u7_n145 ) , .B1( u0_u12_u7_n161 ) , .A2( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n170 ) , .A1( u0_u12_u7_n176 ) );
  INV_X1 u0_u12_u7_U18 (.A( u0_u12_u7_n133 ) , .ZN( u0_u12_u7_n176 ) );
  NOR3_X1 u0_u12_u7_U19 (.A2( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n135 ) , .ZN( u0_u12_u7_n136 ) , .A3( u0_u12_u7_n171 ) );
  NOR2_X1 u0_u12_u7_U20 (.A1( u0_u12_u7_n130 ) , .A2( u0_u12_u7_n134 ) , .ZN( u0_u12_u7_n153 ) );
  INV_X1 u0_u12_u7_U21 (.A( u0_u12_u7_n101 ) , .ZN( u0_u12_u7_n165 ) );
  NOR2_X1 u0_u12_u7_U22 (.ZN( u0_u12_u7_n111 ) , .A2( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n169 ) );
  AOI21_X1 u0_u12_u7_U23 (.ZN( u0_u12_u7_n104 ) , .B2( u0_u12_u7_n112 ) , .B1( u0_u12_u7_n127 ) , .A( u0_u12_u7_n164 ) );
  AOI21_X1 u0_u12_u7_U24 (.ZN( u0_u12_u7_n106 ) , .B1( u0_u12_u7_n133 ) , .B2( u0_u12_u7_n146 ) , .A( u0_u12_u7_n162 ) );
  AOI21_X1 u0_u12_u7_U25 (.A( u0_u12_u7_n101 ) , .ZN( u0_u12_u7_n107 ) , .B2( u0_u12_u7_n128 ) , .B1( u0_u12_u7_n175 ) );
  INV_X1 u0_u12_u7_U26 (.A( u0_u12_u7_n138 ) , .ZN( u0_u12_u7_n171 ) );
  INV_X1 u0_u12_u7_U27 (.A( u0_u12_u7_n131 ) , .ZN( u0_u12_u7_n177 ) );
  INV_X1 u0_u12_u7_U28 (.A( u0_u12_u7_n110 ) , .ZN( u0_u12_u7_n174 ) );
  NAND2_X1 u0_u12_u7_U29 (.A1( u0_u12_u7_n129 ) , .A2( u0_u12_u7_n132 ) , .ZN( u0_u12_u7_n149 ) );
  OAI21_X1 u0_u12_u7_U3 (.ZN( u0_u12_u7_n159 ) , .A( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n171 ) , .B1( u0_u12_u7_n174 ) );
  NAND2_X1 u0_u12_u7_U30 (.A1( u0_u12_u7_n113 ) , .A2( u0_u12_u7_n124 ) , .ZN( u0_u12_u7_n130 ) );
  INV_X1 u0_u12_u7_U31 (.A( u0_u12_u7_n112 ) , .ZN( u0_u12_u7_n173 ) );
  INV_X1 u0_u12_u7_U32 (.A( u0_u12_u7_n128 ) , .ZN( u0_u12_u7_n168 ) );
  INV_X1 u0_u12_u7_U33 (.A( u0_u12_u7_n148 ) , .ZN( u0_u12_u7_n169 ) );
  INV_X1 u0_u12_u7_U34 (.A( u0_u12_u7_n127 ) , .ZN( u0_u12_u7_n179 ) );
  NOR2_X1 u0_u12_u7_U35 (.ZN( u0_u12_u7_n101 ) , .A2( u0_u12_u7_n150 ) , .A1( u0_u12_u7_n156 ) );
  AOI211_X1 u0_u12_u7_U36 (.B( u0_u12_u7_n154 ) , .A( u0_u12_u7_n155 ) , .C1( u0_u12_u7_n156 ) , .ZN( u0_u12_u7_n157 ) , .C2( u0_u12_u7_n172 ) );
  INV_X1 u0_u12_u7_U37 (.A( u0_u12_u7_n153 ) , .ZN( u0_u12_u7_n172 ) );
  AOI211_X1 u0_u12_u7_U38 (.B( u0_u12_u7_n139 ) , .A( u0_u12_u7_n140 ) , .C2( u0_u12_u7_n141 ) , .ZN( u0_u12_u7_n142 ) , .C1( u0_u12_u7_n156 ) );
  NAND4_X1 u0_u12_u7_U39 (.A3( u0_u12_u7_n127 ) , .A2( u0_u12_u7_n128 ) , .A1( u0_u12_u7_n129 ) , .ZN( u0_u12_u7_n141 ) , .A4( u0_u12_u7_n147 ) );
  INV_X1 u0_u12_u7_U4 (.A( u0_u12_u7_n111 ) , .ZN( u0_u12_u7_n170 ) );
  AOI21_X1 u0_u12_u7_U40 (.A( u0_u12_u7_n137 ) , .B1( u0_u12_u7_n138 ) , .ZN( u0_u12_u7_n139 ) , .B2( u0_u12_u7_n146 ) );
  OAI22_X1 u0_u12_u7_U41 (.B1( u0_u12_u7_n136 ) , .ZN( u0_u12_u7_n140 ) , .A1( u0_u12_u7_n153 ) , .B2( u0_u12_u7_n162 ) , .A2( u0_u12_u7_n164 ) );
  AOI21_X1 u0_u12_u7_U42 (.ZN( u0_u12_u7_n123 ) , .B1( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n177 ) , .A( u0_u12_u7_n97 ) );
  AOI21_X1 u0_u12_u7_U43 (.B2( u0_u12_u7_n113 ) , .B1( u0_u12_u7_n124 ) , .A( u0_u12_u7_n125 ) , .ZN( u0_u12_u7_n97 ) );
  INV_X1 u0_u12_u7_U44 (.A( u0_u12_u7_n125 ) , .ZN( u0_u12_u7_n161 ) );
  INV_X1 u0_u12_u7_U45 (.A( u0_u12_u7_n152 ) , .ZN( u0_u12_u7_n162 ) );
  AOI22_X1 u0_u12_u7_U46 (.A2( u0_u12_u7_n114 ) , .ZN( u0_u12_u7_n119 ) , .B1( u0_u12_u7_n130 ) , .A1( u0_u12_u7_n156 ) , .B2( u0_u12_u7_n165 ) );
  NAND2_X1 u0_u12_u7_U47 (.A2( u0_u12_u7_n112 ) , .ZN( u0_u12_u7_n114 ) , .A1( u0_u12_u7_n175 ) );
  AND2_X1 u0_u12_u7_U48 (.ZN( u0_u12_u7_n145 ) , .A2( u0_u12_u7_n98 ) , .A1( u0_u12_u7_n99 ) );
  NOR2_X1 u0_u12_u7_U49 (.ZN( u0_u12_u7_n137 ) , .A1( u0_u12_u7_n150 ) , .A2( u0_u12_u7_n161 ) );
  INV_X1 u0_u12_u7_U5 (.A( u0_u12_u7_n149 ) , .ZN( u0_u12_u7_n175 ) );
  AOI21_X1 u0_u12_u7_U50 (.ZN( u0_u12_u7_n105 ) , .B2( u0_u12_u7_n110 ) , .A( u0_u12_u7_n125 ) , .B1( u0_u12_u7_n147 ) );
  NAND2_X1 u0_u12_u7_U51 (.ZN( u0_u12_u7_n146 ) , .A1( u0_u12_u7_n95 ) , .A2( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U52 (.A2( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n147 ) , .A1( u0_u12_u7_n93 ) );
  NAND2_X1 u0_u12_u7_U53 (.A1( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n127 ) , .A2( u0_u12_u7_n99 ) );
  OR2_X1 u0_u12_u7_U54 (.ZN( u0_u12_u7_n126 ) , .A2( u0_u12_u7_n152 ) , .A1( u0_u12_u7_n156 ) );
  NAND2_X1 u0_u12_u7_U55 (.A2( u0_u12_u7_n102 ) , .A1( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n133 ) );
  NAND2_X1 u0_u12_u7_U56 (.ZN( u0_u12_u7_n112 ) , .A2( u0_u12_u7_n96 ) , .A1( u0_u12_u7_n99 ) );
  NAND2_X1 u0_u12_u7_U57 (.A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n128 ) , .A1( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U58 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n113 ) , .A2( u0_u12_u7_n93 ) );
  NAND2_X1 u0_u12_u7_U59 (.A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n124 ) , .A1( u0_u12_u7_n96 ) );
  INV_X1 u0_u12_u7_U6 (.A( u0_u12_u7_n154 ) , .ZN( u0_u12_u7_n178 ) );
  NAND2_X1 u0_u12_u7_U60 (.ZN( u0_u12_u7_n110 ) , .A1( u0_u12_u7_n95 ) , .A2( u0_u12_u7_n96 ) );
  INV_X1 u0_u12_u7_U61 (.A( u0_u12_u7_n150 ) , .ZN( u0_u12_u7_n164 ) );
  AND2_X1 u0_u12_u7_U62 (.ZN( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n93 ) , .A2( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U63 (.A1( u0_u12_u7_n100 ) , .A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n129 ) );
  NAND2_X1 u0_u12_u7_U64 (.A2( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n131 ) , .A1( u0_u12_u7_n95 ) );
  NAND2_X1 u0_u12_u7_U65 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n138 ) , .A2( u0_u12_u7_n99 ) );
  NAND2_X1 u0_u12_u7_U66 (.ZN( u0_u12_u7_n132 ) , .A1( u0_u12_u7_n93 ) , .A2( u0_u12_u7_n96 ) );
  NAND2_X1 u0_u12_u7_U67 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n148 ) , .A2( u0_u12_u7_n95 ) );
  NOR2_X1 u0_u12_u7_U68 (.A2( u0_u12_X_47 ) , .ZN( u0_u12_u7_n150 ) , .A1( u0_u12_u7_n163 ) );
  NOR2_X1 u0_u12_u7_U69 (.A2( u0_u12_X_43 ) , .A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n103 ) );
  AOI211_X1 u0_u12_u7_U7 (.ZN( u0_u12_u7_n116 ) , .A( u0_u12_u7_n155 ) , .C1( u0_u12_u7_n161 ) , .C2( u0_u12_u7_n171 ) , .B( u0_u12_u7_n94 ) );
  NOR2_X1 u0_u12_u7_U70 (.A2( u0_u12_X_48 ) , .A1( u0_u12_u7_n166 ) , .ZN( u0_u12_u7_n95 ) );
  NOR2_X1 u0_u12_u7_U71 (.A2( u0_u12_X_45 ) , .A1( u0_u12_X_48 ) , .ZN( u0_u12_u7_n99 ) );
  NOR2_X1 u0_u12_u7_U72 (.A2( u0_u12_X_44 ) , .A1( u0_u12_u7_n167 ) , .ZN( u0_u12_u7_n98 ) );
  NOR2_X1 u0_u12_u7_U73 (.A2( u0_u12_X_46 ) , .A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n152 ) );
  AND2_X1 u0_u12_u7_U74 (.A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n156 ) , .A2( u0_u12_u7_n163 ) );
  NAND2_X1 u0_u12_u7_U75 (.A2( u0_u12_X_46 ) , .A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n125 ) );
  AND2_X1 u0_u12_u7_U76 (.A2( u0_u12_X_45 ) , .A1( u0_u12_X_48 ) , .ZN( u0_u12_u7_n102 ) );
  AND2_X1 u0_u12_u7_U77 (.A2( u0_u12_X_43 ) , .A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n96 ) );
  AND2_X1 u0_u12_u7_U78 (.A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n100 ) , .A2( u0_u12_u7_n167 ) );
  AND2_X1 u0_u12_u7_U79 (.A1( u0_u12_X_48 ) , .A2( u0_u12_u7_n166 ) , .ZN( u0_u12_u7_n93 ) );
  OAI222_X1 u0_u12_u7_U8 (.C2( u0_u12_u7_n101 ) , .B2( u0_u12_u7_n111 ) , .A1( u0_u12_u7_n113 ) , .C1( u0_u12_u7_n146 ) , .A2( u0_u12_u7_n162 ) , .B1( u0_u12_u7_n164 ) , .ZN( u0_u12_u7_n94 ) );
  INV_X1 u0_u12_u7_U80 (.A( u0_u12_X_46 ) , .ZN( u0_u12_u7_n163 ) );
  INV_X1 u0_u12_u7_U81 (.A( u0_u12_X_43 ) , .ZN( u0_u12_u7_n167 ) );
  INV_X1 u0_u12_u7_U82 (.A( u0_u12_X_45 ) , .ZN( u0_u12_u7_n166 ) );
  NAND4_X1 u0_u12_u7_U83 (.ZN( u0_out12_27 ) , .A4( u0_u12_u7_n118 ) , .A3( u0_u12_u7_n119 ) , .A2( u0_u12_u7_n120 ) , .A1( u0_u12_u7_n121 ) );
  OAI21_X1 u0_u12_u7_U84 (.ZN( u0_u12_u7_n121 ) , .B2( u0_u12_u7_n145 ) , .A( u0_u12_u7_n150 ) , .B1( u0_u12_u7_n174 ) );
  OAI21_X1 u0_u12_u7_U85 (.ZN( u0_u12_u7_n120 ) , .A( u0_u12_u7_n161 ) , .B2( u0_u12_u7_n170 ) , .B1( u0_u12_u7_n179 ) );
  NAND4_X1 u0_u12_u7_U86 (.ZN( u0_out12_21 ) , .A4( u0_u12_u7_n157 ) , .A3( u0_u12_u7_n158 ) , .A2( u0_u12_u7_n159 ) , .A1( u0_u12_u7_n160 ) );
  OAI21_X1 u0_u12_u7_U87 (.B1( u0_u12_u7_n145 ) , .ZN( u0_u12_u7_n160 ) , .A( u0_u12_u7_n161 ) , .B2( u0_u12_u7_n177 ) );
  AOI22_X1 u0_u12_u7_U88 (.B2( u0_u12_u7_n149 ) , .B1( u0_u12_u7_n150 ) , .A2( u0_u12_u7_n151 ) , .A1( u0_u12_u7_n152 ) , .ZN( u0_u12_u7_n158 ) );
  NAND4_X1 u0_u12_u7_U89 (.ZN( u0_out12_15 ) , .A4( u0_u12_u7_n142 ) , .A3( u0_u12_u7_n143 ) , .A2( u0_u12_u7_n144 ) , .A1( u0_u12_u7_n178 ) );
  OAI221_X1 u0_u12_u7_U9 (.C1( u0_u12_u7_n101 ) , .C2( u0_u12_u7_n147 ) , .ZN( u0_u12_u7_n155 ) , .B2( u0_u12_u7_n162 ) , .A( u0_u12_u7_n91 ) , .B1( u0_u12_u7_n92 ) );
  OR2_X1 u0_u12_u7_U90 (.A2( u0_u12_u7_n125 ) , .A1( u0_u12_u7_n129 ) , .ZN( u0_u12_u7_n144 ) );
  AOI22_X1 u0_u12_u7_U91 (.A2( u0_u12_u7_n126 ) , .ZN( u0_u12_u7_n143 ) , .B2( u0_u12_u7_n165 ) , .B1( u0_u12_u7_n173 ) , .A1( u0_u12_u7_n174 ) );
  NAND4_X1 u0_u12_u7_U92 (.ZN( u0_out12_5 ) , .A4( u0_u12_u7_n108 ) , .A3( u0_u12_u7_n109 ) , .A1( u0_u12_u7_n116 ) , .A2( u0_u12_u7_n123 ) );
  AOI22_X1 u0_u12_u7_U93 (.ZN( u0_u12_u7_n109 ) , .A2( u0_u12_u7_n126 ) , .B2( u0_u12_u7_n145 ) , .B1( u0_u12_u7_n156 ) , .A1( u0_u12_u7_n171 ) );
  NOR4_X1 u0_u12_u7_U94 (.A4( u0_u12_u7_n104 ) , .A3( u0_u12_u7_n105 ) , .A2( u0_u12_u7_n106 ) , .A1( u0_u12_u7_n107 ) , .ZN( u0_u12_u7_n108 ) );
  NAND3_X1 u0_u12_u7_U95 (.A3( u0_u12_u7_n146 ) , .A2( u0_u12_u7_n147 ) , .A1( u0_u12_u7_n148 ) , .ZN( u0_u12_u7_n151 ) );
  NAND3_X1 u0_u12_u7_U96 (.A3( u0_u12_u7_n131 ) , .A2( u0_u12_u7_n132 ) , .A1( u0_u12_u7_n133 ) , .ZN( u0_u12_u7_n135 ) );
  XOR2_X1 u0_u13_U10 (.B( u0_K14_45 ) , .A( u0_R12_30 ) , .Z( u0_u13_X_45 ) );
  AND3_X1 u0_u13_u7_U10 (.A3( u0_u13_u7_n110 ) , .A2( u0_u13_u7_n127 ) , .A1( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n92 ) );
  OAI21_X1 u0_u13_u7_U11 (.A( u0_u13_u7_n161 ) , .B1( u0_u13_u7_n168 ) , .B2( u0_u13_u7_n173 ) , .ZN( u0_u13_u7_n91 ) );
  AOI211_X1 u0_u13_u7_U12 (.A( u0_u13_u7_n117 ) , .ZN( u0_u13_u7_n118 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n177 ) , .B( u0_u13_u7_n180 ) );
  OAI22_X1 u0_u13_u7_U13 (.B1( u0_u13_u7_n115 ) , .ZN( u0_u13_u7_n117 ) , .A2( u0_u13_u7_n133 ) , .A1( u0_u13_u7_n137 ) , .B2( u0_u13_u7_n162 ) );
  INV_X1 u0_u13_u7_U14 (.A( u0_u13_u7_n116 ) , .ZN( u0_u13_u7_n180 ) );
  NOR3_X1 u0_u13_u7_U15 (.ZN( u0_u13_u7_n115 ) , .A3( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n168 ) , .A1( u0_u13_u7_n169 ) );
  OAI211_X1 u0_u13_u7_U16 (.B( u0_u13_u7_n122 ) , .A( u0_u13_u7_n123 ) , .C2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n154 ) , .C1( u0_u13_u7_n162 ) );
  AOI222_X1 u0_u13_u7_U17 (.ZN( u0_u13_u7_n122 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n161 ) , .A2( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n170 ) , .A1( u0_u13_u7_n176 ) );
  INV_X1 u0_u13_u7_U18 (.A( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n176 ) );
  NOR3_X1 u0_u13_u7_U19 (.A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n135 ) , .ZN( u0_u13_u7_n136 ) , .A3( u0_u13_u7_n171 ) );
  NOR2_X1 u0_u13_u7_U20 (.A1( u0_u13_u7_n130 ) , .A2( u0_u13_u7_n134 ) , .ZN( u0_u13_u7_n153 ) );
  INV_X1 u0_u13_u7_U21 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n165 ) );
  NOR2_X1 u0_u13_u7_U22 (.ZN( u0_u13_u7_n111 ) , .A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n169 ) );
  AOI21_X1 u0_u13_u7_U23 (.ZN( u0_u13_u7_n104 ) , .B2( u0_u13_u7_n112 ) , .B1( u0_u13_u7_n127 ) , .A( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U24 (.ZN( u0_u13_u7_n106 ) , .B1( u0_u13_u7_n133 ) , .B2( u0_u13_u7_n146 ) , .A( u0_u13_u7_n162 ) );
  AOI21_X1 u0_u13_u7_U25 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n107 ) , .B2( u0_u13_u7_n128 ) , .B1( u0_u13_u7_n175 ) );
  INV_X1 u0_u13_u7_U26 (.A( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n171 ) );
  INV_X1 u0_u13_u7_U27 (.A( u0_u13_u7_n131 ) , .ZN( u0_u13_u7_n177 ) );
  INV_X1 u0_u13_u7_U28 (.A( u0_u13_u7_n110 ) , .ZN( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U29 (.A1( u0_u13_u7_n129 ) , .A2( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n149 ) );
  OAI21_X1 u0_u13_u7_U3 (.ZN( u0_u13_u7_n159 ) , .A( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n171 ) , .B1( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U30 (.A1( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n130 ) );
  INV_X1 u0_u13_u7_U31 (.A( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n173 ) );
  INV_X1 u0_u13_u7_U32 (.A( u0_u13_u7_n128 ) , .ZN( u0_u13_u7_n168 ) );
  INV_X1 u0_u13_u7_U33 (.A( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n169 ) );
  INV_X1 u0_u13_u7_U34 (.A( u0_u13_u7_n127 ) , .ZN( u0_u13_u7_n179 ) );
  NOR2_X1 u0_u13_u7_U35 (.ZN( u0_u13_u7_n101 ) , .A2( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n156 ) );
  AOI211_X1 u0_u13_u7_U36 (.B( u0_u13_u7_n154 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n156 ) , .ZN( u0_u13_u7_n157 ) , .C2( u0_u13_u7_n172 ) );
  INV_X1 u0_u13_u7_U37 (.A( u0_u13_u7_n153 ) , .ZN( u0_u13_u7_n172 ) );
  AOI211_X1 u0_u13_u7_U38 (.B( u0_u13_u7_n139 ) , .A( u0_u13_u7_n140 ) , .C2( u0_u13_u7_n141 ) , .ZN( u0_u13_u7_n142 ) , .C1( u0_u13_u7_n156 ) );
  NAND4_X1 u0_u13_u7_U39 (.A3( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n141 ) , .A4( u0_u13_u7_n147 ) );
  INV_X1 u0_u13_u7_U4 (.A( u0_u13_u7_n111 ) , .ZN( u0_u13_u7_n170 ) );
  AOI21_X1 u0_u13_u7_U40 (.A( u0_u13_u7_n137 ) , .B1( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n139 ) , .B2( u0_u13_u7_n146 ) );
  OAI22_X1 u0_u13_u7_U41 (.B1( u0_u13_u7_n136 ) , .ZN( u0_u13_u7_n140 ) , .A1( u0_u13_u7_n153 ) , .B2( u0_u13_u7_n162 ) , .A2( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U42 (.ZN( u0_u13_u7_n123 ) , .B1( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n177 ) , .A( u0_u13_u7_n97 ) );
  AOI21_X1 u0_u13_u7_U43 (.B2( u0_u13_u7_n113 ) , .B1( u0_u13_u7_n124 ) , .A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n97 ) );
  INV_X1 u0_u13_u7_U44 (.A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U45 (.A( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n162 ) );
  AOI22_X1 u0_u13_u7_U46 (.A2( u0_u13_u7_n114 ) , .ZN( u0_u13_u7_n119 ) , .B1( u0_u13_u7_n130 ) , .A1( u0_u13_u7_n156 ) , .B2( u0_u13_u7_n165 ) );
  NAND2_X1 u0_u13_u7_U47 (.A2( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n114 ) , .A1( u0_u13_u7_n175 ) );
  AND2_X1 u0_u13_u7_U48 (.ZN( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n98 ) , .A1( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U49 (.ZN( u0_u13_u7_n137 ) , .A1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U5 (.A( u0_u13_u7_n149 ) , .ZN( u0_u13_u7_n175 ) );
  AOI21_X1 u0_u13_u7_U50 (.ZN( u0_u13_u7_n105 ) , .B2( u0_u13_u7_n110 ) , .A( u0_u13_u7_n125 ) , .B1( u0_u13_u7_n147 ) );
  NAND2_X1 u0_u13_u7_U51 (.ZN( u0_u13_u7_n146 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U52 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U53 (.A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n99 ) );
  OR2_X1 u0_u13_u7_U54 (.ZN( u0_u13_u7_n126 ) , .A2( u0_u13_u7_n152 ) , .A1( u0_u13_u7_n156 ) );
  NAND2_X1 u0_u13_u7_U55 (.A2( u0_u13_u7_n102 ) , .A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n133 ) );
  NAND2_X1 u0_u13_u7_U56 (.ZN( u0_u13_u7_n112 ) , .A2( u0_u13_u7_n96 ) , .A1( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U57 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U58 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U59 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n124 ) , .A1( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U6 (.A( u0_u13_u7_n154 ) , .ZN( u0_u13_u7_n178 ) );
  NAND2_X1 u0_u13_u7_U60 (.ZN( u0_u13_u7_n110 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U61 (.A( u0_u13_u7_n150 ) , .ZN( u0_u13_u7_n164 ) );
  AND2_X1 u0_u13_u7_U62 (.ZN( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U63 (.A1( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n129 ) );
  NAND2_X1 u0_u13_u7_U64 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n131 ) , .A1( u0_u13_u7_n95 ) );
  NAND2_X1 u0_u13_u7_U65 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n138 ) , .A2( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U66 (.ZN( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n96 ) );
  NAND2_X1 u0_u13_u7_U67 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n148 ) , .A2( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U68 (.A2( u0_u13_X_47 ) , .ZN( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n163 ) );
  NOR2_X1 u0_u13_u7_U69 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n103 ) );
  AOI211_X1 u0_u13_u7_U7 (.ZN( u0_u13_u7_n116 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n161 ) , .C2( u0_u13_u7_n171 ) , .B( u0_u13_u7_n94 ) );
  NOR2_X1 u0_u13_u7_U70 (.A2( u0_u13_X_48 ) , .A1( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U71 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U72 (.A2( u0_u13_X_44 ) , .A1( u0_u13_u7_n167 ) , .ZN( u0_u13_u7_n98 ) );
  NOR2_X1 u0_u13_u7_U73 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n152 ) );
  AND2_X1 u0_u13_u7_U74 (.A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n156 ) , .A2( u0_u13_u7_n163 ) );
  NAND2_X1 u0_u13_u7_U75 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n125 ) );
  AND2_X1 u0_u13_u7_U76 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n102 ) );
  AND2_X1 u0_u13_u7_U77 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n96 ) );
  AND2_X1 u0_u13_u7_U78 (.A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n167 ) );
  AND2_X1 u0_u13_u7_U79 (.A1( u0_u13_X_48 ) , .A2( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n93 ) );
  OAI222_X1 u0_u13_u7_U8 (.C2( u0_u13_u7_n101 ) , .B2( u0_u13_u7_n111 ) , .A1( u0_u13_u7_n113 ) , .C1( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n162 ) , .B1( u0_u13_u7_n164 ) , .ZN( u0_u13_u7_n94 ) );
  INV_X1 u0_u13_u7_U80 (.A( u0_u13_X_46 ) , .ZN( u0_u13_u7_n163 ) );
  INV_X1 u0_u13_u7_U81 (.A( u0_u13_X_43 ) , .ZN( u0_u13_u7_n167 ) );
  INV_X1 u0_u13_u7_U82 (.A( u0_u13_X_45 ) , .ZN( u0_u13_u7_n166 ) );
  NAND4_X1 u0_u13_u7_U83 (.ZN( u0_out13_27 ) , .A4( u0_u13_u7_n118 ) , .A3( u0_u13_u7_n119 ) , .A2( u0_u13_u7_n120 ) , .A1( u0_u13_u7_n121 ) );
  OAI21_X1 u0_u13_u7_U84 (.ZN( u0_u13_u7_n121 ) , .B2( u0_u13_u7_n145 ) , .A( u0_u13_u7_n150 ) , .B1( u0_u13_u7_n174 ) );
  OAI21_X1 u0_u13_u7_U85 (.ZN( u0_u13_u7_n120 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n170 ) , .B1( u0_u13_u7_n179 ) );
  NAND4_X1 u0_u13_u7_U86 (.ZN( u0_out13_21 ) , .A4( u0_u13_u7_n157 ) , .A3( u0_u13_u7_n158 ) , .A2( u0_u13_u7_n159 ) , .A1( u0_u13_u7_n160 ) );
  OAI21_X1 u0_u13_u7_U87 (.B1( u0_u13_u7_n145 ) , .ZN( u0_u13_u7_n160 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n177 ) );
  AOI22_X1 u0_u13_u7_U88 (.B2( u0_u13_u7_n149 ) , .B1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n151 ) , .A1( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n158 ) );
  NAND4_X1 u0_u13_u7_U89 (.ZN( u0_out13_15 ) , .A4( u0_u13_u7_n142 ) , .A3( u0_u13_u7_n143 ) , .A2( u0_u13_u7_n144 ) , .A1( u0_u13_u7_n178 ) );
  OAI221_X1 u0_u13_u7_U9 (.C1( u0_u13_u7_n101 ) , .C2( u0_u13_u7_n147 ) , .ZN( u0_u13_u7_n155 ) , .B2( u0_u13_u7_n162 ) , .A( u0_u13_u7_n91 ) , .B1( u0_u13_u7_n92 ) );
  OR2_X1 u0_u13_u7_U90 (.A2( u0_u13_u7_n125 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n144 ) );
  AOI22_X1 u0_u13_u7_U91 (.A2( u0_u13_u7_n126 ) , .ZN( u0_u13_u7_n143 ) , .B2( u0_u13_u7_n165 ) , .B1( u0_u13_u7_n173 ) , .A1( u0_u13_u7_n174 ) );
  NAND4_X1 u0_u13_u7_U92 (.ZN( u0_out13_5 ) , .A4( u0_u13_u7_n108 ) , .A3( u0_u13_u7_n109 ) , .A1( u0_u13_u7_n116 ) , .A2( u0_u13_u7_n123 ) );
  AOI22_X1 u0_u13_u7_U93 (.ZN( u0_u13_u7_n109 ) , .A2( u0_u13_u7_n126 ) , .B2( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n156 ) , .A1( u0_u13_u7_n171 ) );
  NOR4_X1 u0_u13_u7_U94 (.A4( u0_u13_u7_n104 ) , .A3( u0_u13_u7_n105 ) , .A2( u0_u13_u7_n106 ) , .A1( u0_u13_u7_n107 ) , .ZN( u0_u13_u7_n108 ) );
  NAND3_X1 u0_u13_u7_U95 (.A3( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n151 ) );
  NAND3_X1 u0_u13_u7_U96 (.A3( u0_u13_u7_n131 ) , .A2( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n135 ) );
  XOR2_X1 u0_u14_U45 (.B( u0_K15_13 ) , .A( u0_R13_8 ) , .Z( u0_u14_X_13 ) );
  XOR2_X1 u0_u14_U47 (.B( u0_K15_11 ) , .A( u0_R13_8 ) , .Z( u0_u14_X_11 ) );
  AOI21_X1 u0_u14_u1_U10 (.ZN( u0_u14_u1_n106 ) , .A( u0_u14_u1_n112 ) , .B1( u0_u14_u1_n154 ) , .B2( u0_u14_u1_n156 ) );
  NAND3_X1 u0_u14_u1_U100 (.ZN( u0_u14_u1_n113 ) , .A1( u0_u14_u1_n120 ) , .A3( u0_u14_u1_n133 ) , .A2( u0_u14_u1_n155 ) );
  INV_X1 u0_u14_u1_U11 (.A( u0_u14_u1_n101 ) , .ZN( u0_u14_u1_n184 ) );
  AOI21_X1 u0_u14_u1_U12 (.ZN( u0_u14_u1_n107 ) , .B1( u0_u14_u1_n134 ) , .B2( u0_u14_u1_n149 ) , .A( u0_u14_u1_n174 ) );
  NAND2_X1 u0_u14_u1_U13 (.ZN( u0_u14_u1_n140 ) , .A2( u0_u14_u1_n150 ) , .A1( u0_u14_u1_n155 ) );
  NAND2_X1 u0_u14_u1_U14 (.A1( u0_u14_u1_n131 ) , .ZN( u0_u14_u1_n147 ) , .A2( u0_u14_u1_n153 ) );
  AOI22_X1 u0_u14_u1_U15 (.B2( u0_u14_u1_n136 ) , .A2( u0_u14_u1_n137 ) , .ZN( u0_u14_u1_n143 ) , .A1( u0_u14_u1_n171 ) , .B1( u0_u14_u1_n173 ) );
  INV_X1 u0_u14_u1_U16 (.A( u0_u14_u1_n147 ) , .ZN( u0_u14_u1_n181 ) );
  INV_X1 u0_u14_u1_U17 (.A( u0_u14_u1_n139 ) , .ZN( u0_u14_u1_n174 ) );
  INV_X1 u0_u14_u1_U18 (.A( u0_u14_u1_n112 ) , .ZN( u0_u14_u1_n171 ) );
  NAND2_X1 u0_u14_u1_U19 (.ZN( u0_u14_u1_n141 ) , .A1( u0_u14_u1_n153 ) , .A2( u0_u14_u1_n156 ) );
  AND2_X1 u0_u14_u1_U20 (.A1( u0_u14_u1_n123 ) , .ZN( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n161 ) );
  NAND2_X1 u0_u14_u1_U21 (.A2( u0_u14_u1_n115 ) , .A1( u0_u14_u1_n116 ) , .ZN( u0_u14_u1_n148 ) );
  NAND2_X1 u0_u14_u1_U22 (.A2( u0_u14_u1_n133 ) , .A1( u0_u14_u1_n135 ) , .ZN( u0_u14_u1_n159 ) );
  NAND2_X1 u0_u14_u1_U23 (.A2( u0_u14_u1_n115 ) , .A1( u0_u14_u1_n120 ) , .ZN( u0_u14_u1_n132 ) );
  INV_X1 u0_u14_u1_U24 (.A( u0_u14_u1_n154 ) , .ZN( u0_u14_u1_n178 ) );
  AOI22_X1 u0_u14_u1_U25 (.B2( u0_u14_u1_n113 ) , .A2( u0_u14_u1_n114 ) , .ZN( u0_u14_u1_n125 ) , .A1( u0_u14_u1_n171 ) , .B1( u0_u14_u1_n173 ) );
  NAND2_X1 u0_u14_u1_U26 (.ZN( u0_u14_u1_n114 ) , .A1( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n156 ) );
  INV_X1 u0_u14_u1_U27 (.A( u0_u14_u1_n151 ) , .ZN( u0_u14_u1_n183 ) );
  AND2_X1 u0_u14_u1_U28 (.A1( u0_u14_u1_n129 ) , .A2( u0_u14_u1_n133 ) , .ZN( u0_u14_u1_n149 ) );
  INV_X1 u0_u14_u1_U29 (.A( u0_u14_u1_n131 ) , .ZN( u0_u14_u1_n180 ) );
  INV_X1 u0_u14_u1_U3 (.A( u0_u14_u1_n159 ) , .ZN( u0_u14_u1_n182 ) );
  AOI221_X1 u0_u14_u1_U30 (.B1( u0_u14_u1_n140 ) , .ZN( u0_u14_u1_n167 ) , .B2( u0_u14_u1_n172 ) , .C2( u0_u14_u1_n175 ) , .C1( u0_u14_u1_n178 ) , .A( u0_u14_u1_n188 ) );
  INV_X1 u0_u14_u1_U31 (.ZN( u0_u14_u1_n188 ) , .A( u0_u14_u1_n97 ) );
  AOI211_X1 u0_u14_u1_U32 (.A( u0_u14_u1_n118 ) , .C1( u0_u14_u1_n132 ) , .C2( u0_u14_u1_n139 ) , .B( u0_u14_u1_n96 ) , .ZN( u0_u14_u1_n97 ) );
  AOI21_X1 u0_u14_u1_U33 (.B2( u0_u14_u1_n121 ) , .B1( u0_u14_u1_n135 ) , .A( u0_u14_u1_n152 ) , .ZN( u0_u14_u1_n96 ) );
  OAI221_X1 u0_u14_u1_U34 (.A( u0_u14_u1_n119 ) , .C2( u0_u14_u1_n129 ) , .ZN( u0_u14_u1_n138 ) , .B2( u0_u14_u1_n152 ) , .C1( u0_u14_u1_n174 ) , .B1( u0_u14_u1_n187 ) );
  INV_X1 u0_u14_u1_U35 (.A( u0_u14_u1_n148 ) , .ZN( u0_u14_u1_n187 ) );
  AOI211_X1 u0_u14_u1_U36 (.B( u0_u14_u1_n117 ) , .A( u0_u14_u1_n118 ) , .ZN( u0_u14_u1_n119 ) , .C2( u0_u14_u1_n146 ) , .C1( u0_u14_u1_n159 ) );
  NOR2_X1 u0_u14_u1_U37 (.A1( u0_u14_u1_n168 ) , .A2( u0_u14_u1_n176 ) , .ZN( u0_u14_u1_n98 ) );
  AOI211_X1 u0_u14_u1_U38 (.B( u0_u14_u1_n162 ) , .A( u0_u14_u1_n163 ) , .C2( u0_u14_u1_n164 ) , .ZN( u0_u14_u1_n165 ) , .C1( u0_u14_u1_n171 ) );
  AOI21_X1 u0_u14_u1_U39 (.A( u0_u14_u1_n160 ) , .B2( u0_u14_u1_n161 ) , .ZN( u0_u14_u1_n162 ) , .B1( u0_u14_u1_n182 ) );
  AOI221_X1 u0_u14_u1_U4 (.A( u0_u14_u1_n138 ) , .C2( u0_u14_u1_n139 ) , .C1( u0_u14_u1_n140 ) , .B2( u0_u14_u1_n141 ) , .ZN( u0_u14_u1_n142 ) , .B1( u0_u14_u1_n175 ) );
  OR2_X1 u0_u14_u1_U40 (.A2( u0_u14_u1_n157 ) , .A1( u0_u14_u1_n158 ) , .ZN( u0_u14_u1_n163 ) );
  OAI21_X1 u0_u14_u1_U41 (.B2( u0_u14_u1_n123 ) , .ZN( u0_u14_u1_n145 ) , .B1( u0_u14_u1_n160 ) , .A( u0_u14_u1_n185 ) );
  INV_X1 u0_u14_u1_U42 (.A( u0_u14_u1_n122 ) , .ZN( u0_u14_u1_n185 ) );
  AOI21_X1 u0_u14_u1_U43 (.B2( u0_u14_u1_n120 ) , .B1( u0_u14_u1_n121 ) , .ZN( u0_u14_u1_n122 ) , .A( u0_u14_u1_n128 ) );
  NAND2_X1 u0_u14_u1_U44 (.A1( u0_u14_u1_n128 ) , .ZN( u0_u14_u1_n146 ) , .A2( u0_u14_u1_n160 ) );
  NAND2_X1 u0_u14_u1_U45 (.A2( u0_u14_u1_n112 ) , .ZN( u0_u14_u1_n139 ) , .A1( u0_u14_u1_n152 ) );
  NAND2_X1 u0_u14_u1_U46 (.A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n156 ) , .A2( u0_u14_u1_n99 ) );
  NOR2_X1 u0_u14_u1_U47 (.ZN( u0_u14_u1_n117 ) , .A1( u0_u14_u1_n121 ) , .A2( u0_u14_u1_n160 ) );
  AOI21_X1 u0_u14_u1_U48 (.A( u0_u14_u1_n128 ) , .B2( u0_u14_u1_n129 ) , .ZN( u0_u14_u1_n130 ) , .B1( u0_u14_u1_n150 ) );
  NAND2_X1 u0_u14_u1_U49 (.ZN( u0_u14_u1_n112 ) , .A1( u0_u14_u1_n169 ) , .A2( u0_u14_u1_n170 ) );
  AOI211_X1 u0_u14_u1_U5 (.ZN( u0_u14_u1_n124 ) , .A( u0_u14_u1_n138 ) , .C2( u0_u14_u1_n139 ) , .B( u0_u14_u1_n145 ) , .C1( u0_u14_u1_n147 ) );
  NAND2_X1 u0_u14_u1_U50 (.ZN( u0_u14_u1_n129 ) , .A2( u0_u14_u1_n95 ) , .A1( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U51 (.A1( u0_u14_u1_n102 ) , .ZN( u0_u14_u1_n154 ) , .A2( u0_u14_u1_n99 ) );
  NAND2_X1 u0_u14_u1_U52 (.A2( u0_u14_u1_n100 ) , .ZN( u0_u14_u1_n135 ) , .A1( u0_u14_u1_n99 ) );
  AOI21_X1 u0_u14_u1_U53 (.A( u0_u14_u1_n152 ) , .B2( u0_u14_u1_n153 ) , .B1( u0_u14_u1_n154 ) , .ZN( u0_u14_u1_n158 ) );
  INV_X1 u0_u14_u1_U54 (.A( u0_u14_u1_n160 ) , .ZN( u0_u14_u1_n175 ) );
  NAND2_X1 u0_u14_u1_U55 (.A1( u0_u14_u1_n100 ) , .ZN( u0_u14_u1_n116 ) , .A2( u0_u14_u1_n95 ) );
  NAND2_X1 u0_u14_u1_U56 (.A1( u0_u14_u1_n102 ) , .ZN( u0_u14_u1_n131 ) , .A2( u0_u14_u1_n95 ) );
  NAND2_X1 u0_u14_u1_U57 (.A2( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n121 ) , .A1( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U58 (.A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n153 ) , .A2( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U59 (.A2( u0_u14_u1_n104 ) , .A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n133 ) );
  NOR2_X1 u0_u14_u1_U6 (.A1( u0_u14_u1_n112 ) , .A2( u0_u14_u1_n116 ) , .ZN( u0_u14_u1_n118 ) );
  NAND2_X1 u0_u14_u1_U60 (.ZN( u0_u14_u1_n150 ) , .A2( u0_u14_u1_n98 ) , .A1( u0_u14_u1_n99 ) );
  NAND2_X1 u0_u14_u1_U61 (.A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n155 ) , .A2( u0_u14_u1_n95 ) );
  OAI21_X1 u0_u14_u1_U62 (.ZN( u0_u14_u1_n109 ) , .B1( u0_u14_u1_n129 ) , .B2( u0_u14_u1_n160 ) , .A( u0_u14_u1_n167 ) );
  NAND2_X1 u0_u14_u1_U63 (.A2( u0_u14_u1_n100 ) , .A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n120 ) );
  NAND2_X1 u0_u14_u1_U64 (.A1( u0_u14_u1_n102 ) , .A2( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n115 ) );
  NAND2_X1 u0_u14_u1_U65 (.A2( u0_u14_u1_n100 ) , .A1( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n151 ) );
  NAND2_X1 u0_u14_u1_U66 (.A2( u0_u14_u1_n103 ) , .A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n161 ) );
  INV_X1 u0_u14_u1_U67 (.A( u0_u14_u1_n152 ) , .ZN( u0_u14_u1_n173 ) );
  INV_X1 u0_u14_u1_U68 (.A( u0_u14_u1_n128 ) , .ZN( u0_u14_u1_n172 ) );
  NAND2_X1 u0_u14_u1_U69 (.A2( u0_u14_u1_n102 ) , .A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n123 ) );
  OAI21_X1 u0_u14_u1_U7 (.ZN( u0_u14_u1_n101 ) , .B1( u0_u14_u1_n141 ) , .A( u0_u14_u1_n146 ) , .B2( u0_u14_u1_n183 ) );
  NOR2_X1 u0_u14_u1_U70 (.A2( u0_u14_X_7 ) , .A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n95 ) );
  NOR2_X1 u0_u14_u1_U71 (.A1( u0_u14_X_12 ) , .A2( u0_u14_X_9 ) , .ZN( u0_u14_u1_n100 ) );
  NOR2_X1 u0_u14_u1_U72 (.A2( u0_u14_X_8 ) , .A1( u0_u14_u1_n177 ) , .ZN( u0_u14_u1_n99 ) );
  NOR2_X1 u0_u14_u1_U73 (.A2( u0_u14_X_12 ) , .ZN( u0_u14_u1_n102 ) , .A1( u0_u14_u1_n176 ) );
  NOR2_X1 u0_u14_u1_U74 (.A2( u0_u14_X_9 ) , .ZN( u0_u14_u1_n105 ) , .A1( u0_u14_u1_n168 ) );
  NAND2_X1 u0_u14_u1_U75 (.A1( u0_u14_X_10 ) , .ZN( u0_u14_u1_n160 ) , .A2( u0_u14_u1_n169 ) );
  NAND2_X1 u0_u14_u1_U76 (.A2( u0_u14_X_10 ) , .A1( u0_u14_X_11 ) , .ZN( u0_u14_u1_n152 ) );
  NAND2_X1 u0_u14_u1_U77 (.A1( u0_u14_X_11 ) , .ZN( u0_u14_u1_n128 ) , .A2( u0_u14_u1_n170 ) );
  AND2_X1 u0_u14_u1_U78 (.A2( u0_u14_X_7 ) , .A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n104 ) );
  AND2_X1 u0_u14_u1_U79 (.A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n103 ) , .A2( u0_u14_u1_n177 ) );
  AOI21_X1 u0_u14_u1_U8 (.B2( u0_u14_u1_n155 ) , .B1( u0_u14_u1_n156 ) , .ZN( u0_u14_u1_n157 ) , .A( u0_u14_u1_n174 ) );
  INV_X1 u0_u14_u1_U80 (.A( u0_u14_X_10 ) , .ZN( u0_u14_u1_n170 ) );
  INV_X1 u0_u14_u1_U81 (.A( u0_u14_X_9 ) , .ZN( u0_u14_u1_n176 ) );
  INV_X1 u0_u14_u1_U82 (.A( u0_u14_X_11 ) , .ZN( u0_u14_u1_n169 ) );
  INV_X1 u0_u14_u1_U83 (.A( u0_u14_X_12 ) , .ZN( u0_u14_u1_n168 ) );
  INV_X1 u0_u14_u1_U84 (.A( u0_u14_X_7 ) , .ZN( u0_u14_u1_n177 ) );
  NAND4_X1 u0_u14_u1_U85 (.ZN( u0_out14_28 ) , .A4( u0_u14_u1_n124 ) , .A3( u0_u14_u1_n125 ) , .A2( u0_u14_u1_n126 ) , .A1( u0_u14_u1_n127 ) );
  OAI21_X1 u0_u14_u1_U86 (.ZN( u0_u14_u1_n127 ) , .B2( u0_u14_u1_n139 ) , .B1( u0_u14_u1_n175 ) , .A( u0_u14_u1_n183 ) );
  OAI21_X1 u0_u14_u1_U87 (.ZN( u0_u14_u1_n126 ) , .B2( u0_u14_u1_n140 ) , .A( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n178 ) );
  NAND4_X1 u0_u14_u1_U88 (.ZN( u0_out14_18 ) , .A4( u0_u14_u1_n165 ) , .A3( u0_u14_u1_n166 ) , .A1( u0_u14_u1_n167 ) , .A2( u0_u14_u1_n186 ) );
  AOI22_X1 u0_u14_u1_U89 (.B2( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n147 ) , .A2( u0_u14_u1_n148 ) , .ZN( u0_u14_u1_n166 ) , .A1( u0_u14_u1_n172 ) );
  OR4_X1 u0_u14_u1_U9 (.A4( u0_u14_u1_n106 ) , .A3( u0_u14_u1_n107 ) , .ZN( u0_u14_u1_n108 ) , .A1( u0_u14_u1_n117 ) , .A2( u0_u14_u1_n184 ) );
  INV_X1 u0_u14_u1_U90 (.A( u0_u14_u1_n145 ) , .ZN( u0_u14_u1_n186 ) );
  NAND4_X1 u0_u14_u1_U91 (.ZN( u0_out14_2 ) , .A4( u0_u14_u1_n142 ) , .A3( u0_u14_u1_n143 ) , .A2( u0_u14_u1_n144 ) , .A1( u0_u14_u1_n179 ) );
  OAI21_X1 u0_u14_u1_U92 (.B2( u0_u14_u1_n132 ) , .ZN( u0_u14_u1_n144 ) , .A( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n180 ) );
  INV_X1 u0_u14_u1_U93 (.A( u0_u14_u1_n130 ) , .ZN( u0_u14_u1_n179 ) );
  OR4_X1 u0_u14_u1_U94 (.ZN( u0_out14_13 ) , .A4( u0_u14_u1_n108 ) , .A3( u0_u14_u1_n109 ) , .A2( u0_u14_u1_n110 ) , .A1( u0_u14_u1_n111 ) );
  AOI21_X1 u0_u14_u1_U95 (.ZN( u0_u14_u1_n111 ) , .A( u0_u14_u1_n128 ) , .B2( u0_u14_u1_n131 ) , .B1( u0_u14_u1_n135 ) );
  AOI21_X1 u0_u14_u1_U96 (.ZN( u0_u14_u1_n110 ) , .A( u0_u14_u1_n116 ) , .B1( u0_u14_u1_n152 ) , .B2( u0_u14_u1_n160 ) );
  NAND3_X1 u0_u14_u1_U97 (.A3( u0_u14_u1_n149 ) , .A2( u0_u14_u1_n150 ) , .A1( u0_u14_u1_n151 ) , .ZN( u0_u14_u1_n164 ) );
  NAND3_X1 u0_u14_u1_U98 (.A3( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n135 ) , .ZN( u0_u14_u1_n136 ) , .A1( u0_u14_u1_n151 ) );
  NAND3_X1 u0_u14_u1_U99 (.A1( u0_u14_u1_n133 ) , .ZN( u0_u14_u1_n137 ) , .A2( u0_u14_u1_n154 ) , .A3( u0_u14_u1_n181 ) );
  OAI22_X1 u0_u14_u2_U10 (.ZN( u0_u14_u2_n109 ) , .A2( u0_u14_u2_n113 ) , .B2( u0_u14_u2_n133 ) , .B1( u0_u14_u2_n167 ) , .A1( u0_u14_u2_n168 ) );
  NAND3_X1 u0_u14_u2_U100 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n98 ) );
  OAI22_X1 u0_u14_u2_U11 (.B1( u0_u14_u2_n151 ) , .A2( u0_u14_u2_n152 ) , .A1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n160 ) , .B2( u0_u14_u2_n168 ) );
  NOR3_X1 u0_u14_u2_U12 (.A1( u0_u14_u2_n150 ) , .ZN( u0_u14_u2_n151 ) , .A3( u0_u14_u2_n175 ) , .A2( u0_u14_u2_n188 ) );
  AOI21_X1 u0_u14_u2_U13 (.ZN( u0_u14_u2_n144 ) , .B2( u0_u14_u2_n155 ) , .A( u0_u14_u2_n172 ) , .B1( u0_u14_u2_n185 ) );
  AOI21_X1 u0_u14_u2_U14 (.B2( u0_u14_u2_n143 ) , .ZN( u0_u14_u2_n145 ) , .B1( u0_u14_u2_n152 ) , .A( u0_u14_u2_n171 ) );
  AOI21_X1 u0_u14_u2_U15 (.B2( u0_u14_u2_n120 ) , .B1( u0_u14_u2_n121 ) , .ZN( u0_u14_u2_n126 ) , .A( u0_u14_u2_n167 ) );
  INV_X1 u0_u14_u2_U16 (.A( u0_u14_u2_n156 ) , .ZN( u0_u14_u2_n171 ) );
  INV_X1 u0_u14_u2_U17 (.A( u0_u14_u2_n120 ) , .ZN( u0_u14_u2_n188 ) );
  NAND2_X1 u0_u14_u2_U18 (.A2( u0_u14_u2_n122 ) , .ZN( u0_u14_u2_n150 ) , .A1( u0_u14_u2_n152 ) );
  INV_X1 u0_u14_u2_U19 (.A( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n170 ) );
  INV_X1 u0_u14_u2_U20 (.A( u0_u14_u2_n137 ) , .ZN( u0_u14_u2_n173 ) );
  NAND2_X1 u0_u14_u2_U21 (.A1( u0_u14_u2_n132 ) , .A2( u0_u14_u2_n139 ) , .ZN( u0_u14_u2_n157 ) );
  INV_X1 u0_u14_u2_U22 (.A( u0_u14_u2_n113 ) , .ZN( u0_u14_u2_n178 ) );
  INV_X1 u0_u14_u2_U23 (.A( u0_u14_u2_n139 ) , .ZN( u0_u14_u2_n175 ) );
  INV_X1 u0_u14_u2_U24 (.A( u0_u14_u2_n155 ) , .ZN( u0_u14_u2_n181 ) );
  INV_X1 u0_u14_u2_U25 (.A( u0_u14_u2_n119 ) , .ZN( u0_u14_u2_n177 ) );
  INV_X1 u0_u14_u2_U26 (.A( u0_u14_u2_n116 ) , .ZN( u0_u14_u2_n180 ) );
  INV_X1 u0_u14_u2_U27 (.A( u0_u14_u2_n131 ) , .ZN( u0_u14_u2_n179 ) );
  INV_X1 u0_u14_u2_U28 (.A( u0_u14_u2_n154 ) , .ZN( u0_u14_u2_n176 ) );
  NAND2_X1 u0_u14_u2_U29 (.A2( u0_u14_u2_n116 ) , .A1( u0_u14_u2_n117 ) , .ZN( u0_u14_u2_n118 ) );
  NOR2_X1 u0_u14_u2_U3 (.ZN( u0_u14_u2_n121 ) , .A2( u0_u14_u2_n177 ) , .A1( u0_u14_u2_n180 ) );
  INV_X1 u0_u14_u2_U30 (.A( u0_u14_u2_n132 ) , .ZN( u0_u14_u2_n182 ) );
  INV_X1 u0_u14_u2_U31 (.A( u0_u14_u2_n158 ) , .ZN( u0_u14_u2_n183 ) );
  OAI21_X1 u0_u14_u2_U32 (.A( u0_u14_u2_n156 ) , .B1( u0_u14_u2_n157 ) , .ZN( u0_u14_u2_n158 ) , .B2( u0_u14_u2_n179 ) );
  NOR2_X1 u0_u14_u2_U33 (.ZN( u0_u14_u2_n156 ) , .A1( u0_u14_u2_n166 ) , .A2( u0_u14_u2_n169 ) );
  NOR2_X1 u0_u14_u2_U34 (.A2( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n137 ) , .A1( u0_u14_u2_n140 ) );
  NOR2_X1 u0_u14_u2_U35 (.A2( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n153 ) , .A1( u0_u14_u2_n156 ) );
  AOI211_X1 u0_u14_u2_U36 (.ZN( u0_u14_u2_n130 ) , .C1( u0_u14_u2_n138 ) , .C2( u0_u14_u2_n179 ) , .B( u0_u14_u2_n96 ) , .A( u0_u14_u2_n97 ) );
  OAI22_X1 u0_u14_u2_U37 (.B1( u0_u14_u2_n133 ) , .A2( u0_u14_u2_n137 ) , .A1( u0_u14_u2_n152 ) , .B2( u0_u14_u2_n168 ) , .ZN( u0_u14_u2_n97 ) );
  OAI221_X1 u0_u14_u2_U38 (.B1( u0_u14_u2_n113 ) , .C1( u0_u14_u2_n132 ) , .A( u0_u14_u2_n149 ) , .B2( u0_u14_u2_n171 ) , .C2( u0_u14_u2_n172 ) , .ZN( u0_u14_u2_n96 ) );
  OAI221_X1 u0_u14_u2_U39 (.A( u0_u14_u2_n115 ) , .C2( u0_u14_u2_n123 ) , .B2( u0_u14_u2_n143 ) , .B1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n163 ) , .C1( u0_u14_u2_n168 ) );
  INV_X1 u0_u14_u2_U4 (.A( u0_u14_u2_n134 ) , .ZN( u0_u14_u2_n185 ) );
  OAI21_X1 u0_u14_u2_U40 (.A( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n115 ) , .B1( u0_u14_u2_n176 ) , .B2( u0_u14_u2_n178 ) );
  OAI221_X1 u0_u14_u2_U41 (.A( u0_u14_u2_n135 ) , .B2( u0_u14_u2_n136 ) , .B1( u0_u14_u2_n137 ) , .ZN( u0_u14_u2_n162 ) , .C2( u0_u14_u2_n167 ) , .C1( u0_u14_u2_n185 ) );
  AND3_X1 u0_u14_u2_U42 (.A3( u0_u14_u2_n131 ) , .A2( u0_u14_u2_n132 ) , .A1( u0_u14_u2_n133 ) , .ZN( u0_u14_u2_n136 ) );
  AOI22_X1 u0_u14_u2_U43 (.ZN( u0_u14_u2_n135 ) , .B1( u0_u14_u2_n140 ) , .A1( u0_u14_u2_n156 ) , .B2( u0_u14_u2_n180 ) , .A2( u0_u14_u2_n188 ) );
  AOI21_X1 u0_u14_u2_U44 (.ZN( u0_u14_u2_n149 ) , .B1( u0_u14_u2_n173 ) , .B2( u0_u14_u2_n188 ) , .A( u0_u14_u2_n95 ) );
  AND3_X1 u0_u14_u2_U45 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n156 ) , .ZN( u0_u14_u2_n95 ) );
  OAI21_X1 u0_u14_u2_U46 (.A( u0_u14_u2_n141 ) , .B2( u0_u14_u2_n142 ) , .ZN( u0_u14_u2_n146 ) , .B1( u0_u14_u2_n153 ) );
  OAI21_X1 u0_u14_u2_U47 (.A( u0_u14_u2_n140 ) , .ZN( u0_u14_u2_n141 ) , .B1( u0_u14_u2_n176 ) , .B2( u0_u14_u2_n177 ) );
  NOR3_X1 u0_u14_u2_U48 (.ZN( u0_u14_u2_n142 ) , .A3( u0_u14_u2_n175 ) , .A2( u0_u14_u2_n178 ) , .A1( u0_u14_u2_n181 ) );
  OAI21_X1 u0_u14_u2_U49 (.A( u0_u14_u2_n101 ) , .B2( u0_u14_u2_n121 ) , .B1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n164 ) );
  INV_X1 u0_u14_u2_U5 (.A( u0_u14_u2_n150 ) , .ZN( u0_u14_u2_n184 ) );
  NAND2_X1 u0_u14_u2_U50 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n155 ) );
  NAND2_X1 u0_u14_u2_U51 (.A2( u0_u14_u2_n105 ) , .A1( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n143 ) );
  NAND2_X1 u0_u14_u2_U52 (.A1( u0_u14_u2_n104 ) , .A2( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n152 ) );
  NAND2_X1 u0_u14_u2_U53 (.A1( u0_u14_u2_n100 ) , .A2( u0_u14_u2_n105 ) , .ZN( u0_u14_u2_n132 ) );
  INV_X1 u0_u14_u2_U54 (.A( u0_u14_u2_n140 ) , .ZN( u0_u14_u2_n168 ) );
  INV_X1 u0_u14_u2_U55 (.A( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n167 ) );
  INV_X1 u0_u14_u2_U56 (.ZN( u0_u14_u2_n187 ) , .A( u0_u14_u2_n99 ) );
  OAI21_X1 u0_u14_u2_U57 (.B1( u0_u14_u2_n137 ) , .B2( u0_u14_u2_n143 ) , .A( u0_u14_u2_n98 ) , .ZN( u0_u14_u2_n99 ) );
  NAND2_X1 u0_u14_u2_U58 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n113 ) );
  NAND2_X1 u0_u14_u2_U59 (.A1( u0_u14_u2_n106 ) , .A2( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n131 ) );
  NOR4_X1 u0_u14_u2_U6 (.A4( u0_u14_u2_n124 ) , .A3( u0_u14_u2_n125 ) , .A2( u0_u14_u2_n126 ) , .A1( u0_u14_u2_n127 ) , .ZN( u0_u14_u2_n128 ) );
  NAND2_X1 u0_u14_u2_U60 (.A1( u0_u14_u2_n103 ) , .A2( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n139 ) );
  NAND2_X1 u0_u14_u2_U61 (.A1( u0_u14_u2_n103 ) , .A2( u0_u14_u2_n105 ) , .ZN( u0_u14_u2_n133 ) );
  NAND2_X1 u0_u14_u2_U62 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n103 ) , .ZN( u0_u14_u2_n154 ) );
  NAND2_X1 u0_u14_u2_U63 (.A2( u0_u14_u2_n103 ) , .A1( u0_u14_u2_n104 ) , .ZN( u0_u14_u2_n119 ) );
  NAND2_X1 u0_u14_u2_U64 (.A2( u0_u14_u2_n107 ) , .A1( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n123 ) );
  NAND2_X1 u0_u14_u2_U65 (.A1( u0_u14_u2_n104 ) , .A2( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n122 ) );
  INV_X1 u0_u14_u2_U66 (.A( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n172 ) );
  NAND2_X1 u0_u14_u2_U67 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n102 ) , .ZN( u0_u14_u2_n116 ) );
  NAND2_X1 u0_u14_u2_U68 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n120 ) );
  NAND2_X1 u0_u14_u2_U69 (.A2( u0_u14_u2_n105 ) , .A1( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n117 ) );
  AOI21_X1 u0_u14_u2_U7 (.B2( u0_u14_u2_n119 ) , .ZN( u0_u14_u2_n127 ) , .A( u0_u14_u2_n137 ) , .B1( u0_u14_u2_n155 ) );
  NOR2_X1 u0_u14_u2_U70 (.A2( u0_u14_X_16 ) , .ZN( u0_u14_u2_n140 ) , .A1( u0_u14_u2_n166 ) );
  NOR2_X1 u0_u14_u2_U71 (.A2( u0_u14_X_13 ) , .A1( u0_u14_X_14 ) , .ZN( u0_u14_u2_n100 ) );
  NOR2_X1 u0_u14_u2_U72 (.A2( u0_u14_X_16 ) , .A1( u0_u14_X_17 ) , .ZN( u0_u14_u2_n138 ) );
  NOR2_X1 u0_u14_u2_U73 (.A2( u0_u14_X_15 ) , .A1( u0_u14_X_18 ) , .ZN( u0_u14_u2_n104 ) );
  NOR2_X1 u0_u14_u2_U74 (.A2( u0_u14_X_14 ) , .ZN( u0_u14_u2_n103 ) , .A1( u0_u14_u2_n174 ) );
  NOR2_X1 u0_u14_u2_U75 (.A2( u0_u14_X_15 ) , .ZN( u0_u14_u2_n102 ) , .A1( u0_u14_u2_n165 ) );
  NOR2_X1 u0_u14_u2_U76 (.A2( u0_u14_X_17 ) , .ZN( u0_u14_u2_n114 ) , .A1( u0_u14_u2_n169 ) );
  AND2_X1 u0_u14_u2_U77 (.A1( u0_u14_X_15 ) , .ZN( u0_u14_u2_n105 ) , .A2( u0_u14_u2_n165 ) );
  AND2_X1 u0_u14_u2_U78 (.A2( u0_u14_X_15 ) , .A1( u0_u14_X_18 ) , .ZN( u0_u14_u2_n107 ) );
  AND2_X1 u0_u14_u2_U79 (.A1( u0_u14_X_14 ) , .ZN( u0_u14_u2_n106 ) , .A2( u0_u14_u2_n174 ) );
  AOI21_X1 u0_u14_u2_U8 (.ZN( u0_u14_u2_n124 ) , .B1( u0_u14_u2_n131 ) , .B2( u0_u14_u2_n143 ) , .A( u0_u14_u2_n172 ) );
  AND2_X1 u0_u14_u2_U80 (.A1( u0_u14_X_13 ) , .A2( u0_u14_X_14 ) , .ZN( u0_u14_u2_n108 ) );
  INV_X1 u0_u14_u2_U81 (.A( u0_u14_X_16 ) , .ZN( u0_u14_u2_n169 ) );
  INV_X1 u0_u14_u2_U82 (.A( u0_u14_X_17 ) , .ZN( u0_u14_u2_n166 ) );
  INV_X1 u0_u14_u2_U83 (.A( u0_u14_X_13 ) , .ZN( u0_u14_u2_n174 ) );
  INV_X1 u0_u14_u2_U84 (.A( u0_u14_X_18 ) , .ZN( u0_u14_u2_n165 ) );
  NAND4_X1 u0_u14_u2_U85 (.ZN( u0_out14_30 ) , .A4( u0_u14_u2_n147 ) , .A3( u0_u14_u2_n148 ) , .A2( u0_u14_u2_n149 ) , .A1( u0_u14_u2_n187 ) );
  NOR3_X1 u0_u14_u2_U86 (.A3( u0_u14_u2_n144 ) , .A2( u0_u14_u2_n145 ) , .A1( u0_u14_u2_n146 ) , .ZN( u0_u14_u2_n147 ) );
  AOI21_X1 u0_u14_u2_U87 (.B2( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n148 ) , .A( u0_u14_u2_n162 ) , .B1( u0_u14_u2_n182 ) );
  NAND4_X1 u0_u14_u2_U88 (.ZN( u0_out14_24 ) , .A4( u0_u14_u2_n111 ) , .A3( u0_u14_u2_n112 ) , .A1( u0_u14_u2_n130 ) , .A2( u0_u14_u2_n187 ) );
  AOI221_X1 u0_u14_u2_U89 (.A( u0_u14_u2_n109 ) , .B1( u0_u14_u2_n110 ) , .ZN( u0_u14_u2_n111 ) , .C1( u0_u14_u2_n134 ) , .C2( u0_u14_u2_n170 ) , .B2( u0_u14_u2_n173 ) );
  AOI21_X1 u0_u14_u2_U9 (.B2( u0_u14_u2_n123 ) , .ZN( u0_u14_u2_n125 ) , .A( u0_u14_u2_n171 ) , .B1( u0_u14_u2_n184 ) );
  AOI21_X1 u0_u14_u2_U90 (.ZN( u0_u14_u2_n112 ) , .B2( u0_u14_u2_n156 ) , .A( u0_u14_u2_n164 ) , .B1( u0_u14_u2_n181 ) );
  NAND4_X1 u0_u14_u2_U91 (.ZN( u0_out14_16 ) , .A4( u0_u14_u2_n128 ) , .A3( u0_u14_u2_n129 ) , .A1( u0_u14_u2_n130 ) , .A2( u0_u14_u2_n186 ) );
  AOI22_X1 u0_u14_u2_U92 (.A2( u0_u14_u2_n118 ) , .ZN( u0_u14_u2_n129 ) , .A1( u0_u14_u2_n140 ) , .B1( u0_u14_u2_n157 ) , .B2( u0_u14_u2_n170 ) );
  INV_X1 u0_u14_u2_U93 (.A( u0_u14_u2_n163 ) , .ZN( u0_u14_u2_n186 ) );
  OR4_X1 u0_u14_u2_U94 (.ZN( u0_out14_6 ) , .A4( u0_u14_u2_n161 ) , .A3( u0_u14_u2_n162 ) , .A2( u0_u14_u2_n163 ) , .A1( u0_u14_u2_n164 ) );
  OR3_X1 u0_u14_u2_U95 (.A2( u0_u14_u2_n159 ) , .A1( u0_u14_u2_n160 ) , .ZN( u0_u14_u2_n161 ) , .A3( u0_u14_u2_n183 ) );
  AOI21_X1 u0_u14_u2_U96 (.B2( u0_u14_u2_n154 ) , .B1( u0_u14_u2_n155 ) , .ZN( u0_u14_u2_n159 ) , .A( u0_u14_u2_n167 ) );
  NAND3_X1 u0_u14_u2_U97 (.A2( u0_u14_u2_n117 ) , .A1( u0_u14_u2_n122 ) , .A3( u0_u14_u2_n123 ) , .ZN( u0_u14_u2_n134 ) );
  NAND3_X1 u0_u14_u2_U98 (.ZN( u0_u14_u2_n110 ) , .A2( u0_u14_u2_n131 ) , .A3( u0_u14_u2_n139 ) , .A1( u0_u14_u2_n154 ) );
  NAND3_X1 u0_u14_u2_U99 (.A2( u0_u14_u2_n100 ) , .ZN( u0_u14_u2_n101 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n114 ) );
  OAI22_X1 u0_u14_u3_U10 (.B1( u0_u14_u3_n113 ) , .A2( u0_u14_u3_n135 ) , .A1( u0_u14_u3_n150 ) , .B2( u0_u14_u3_n164 ) , .ZN( u0_u14_u3_n98 ) );
  OAI211_X1 u0_u14_u3_U11 (.B( u0_u14_u3_n106 ) , .ZN( u0_u14_u3_n119 ) , .C2( u0_u14_u3_n128 ) , .C1( u0_u14_u3_n167 ) , .A( u0_u14_u3_n181 ) );
  AOI221_X1 u0_u14_u3_U12 (.C1( u0_u14_u3_n105 ) , .ZN( u0_u14_u3_n106 ) , .A( u0_u14_u3_n131 ) , .B2( u0_u14_u3_n132 ) , .C2( u0_u14_u3_n133 ) , .B1( u0_u14_u3_n169 ) );
  INV_X1 u0_u14_u3_U13 (.ZN( u0_u14_u3_n181 ) , .A( u0_u14_u3_n98 ) );
  NAND2_X1 u0_u14_u3_U14 (.ZN( u0_u14_u3_n105 ) , .A2( u0_u14_u3_n130 ) , .A1( u0_u14_u3_n155 ) );
  AOI22_X1 u0_u14_u3_U15 (.B1( u0_u14_u3_n115 ) , .A2( u0_u14_u3_n116 ) , .ZN( u0_u14_u3_n123 ) , .B2( u0_u14_u3_n133 ) , .A1( u0_u14_u3_n169 ) );
  NAND2_X1 u0_u14_u3_U16 (.ZN( u0_u14_u3_n116 ) , .A2( u0_u14_u3_n151 ) , .A1( u0_u14_u3_n182 ) );
  NOR2_X1 u0_u14_u3_U17 (.ZN( u0_u14_u3_n126 ) , .A2( u0_u14_u3_n150 ) , .A1( u0_u14_u3_n164 ) );
  AOI21_X1 u0_u14_u3_U18 (.ZN( u0_u14_u3_n112 ) , .B2( u0_u14_u3_n146 ) , .B1( u0_u14_u3_n155 ) , .A( u0_u14_u3_n167 ) );
  NAND2_X1 u0_u14_u3_U19 (.A1( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n142 ) , .A2( u0_u14_u3_n164 ) );
  NAND2_X1 u0_u14_u3_U20 (.ZN( u0_u14_u3_n132 ) , .A2( u0_u14_u3_n152 ) , .A1( u0_u14_u3_n156 ) );
  AND2_X1 u0_u14_u3_U21 (.A2( u0_u14_u3_n113 ) , .A1( u0_u14_u3_n114 ) , .ZN( u0_u14_u3_n151 ) );
  INV_X1 u0_u14_u3_U22 (.A( u0_u14_u3_n133 ) , .ZN( u0_u14_u3_n165 ) );
  INV_X1 u0_u14_u3_U23 (.A( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n170 ) );
  NAND2_X1 u0_u14_u3_U24 (.A1( u0_u14_u3_n107 ) , .A2( u0_u14_u3_n108 ) , .ZN( u0_u14_u3_n140 ) );
  NAND2_X1 u0_u14_u3_U25 (.ZN( u0_u14_u3_n117 ) , .A1( u0_u14_u3_n124 ) , .A2( u0_u14_u3_n148 ) );
  NAND2_X1 u0_u14_u3_U26 (.ZN( u0_u14_u3_n143 ) , .A1( u0_u14_u3_n165 ) , .A2( u0_u14_u3_n167 ) );
  INV_X1 u0_u14_u3_U27 (.A( u0_u14_u3_n130 ) , .ZN( u0_u14_u3_n177 ) );
  INV_X1 u0_u14_u3_U28 (.A( u0_u14_u3_n128 ) , .ZN( u0_u14_u3_n176 ) );
  INV_X1 u0_u14_u3_U29 (.A( u0_u14_u3_n155 ) , .ZN( u0_u14_u3_n174 ) );
  INV_X1 u0_u14_u3_U3 (.A( u0_u14_u3_n129 ) , .ZN( u0_u14_u3_n183 ) );
  INV_X1 u0_u14_u3_U30 (.A( u0_u14_u3_n139 ) , .ZN( u0_u14_u3_n185 ) );
  NOR2_X1 u0_u14_u3_U31 (.ZN( u0_u14_u3_n135 ) , .A2( u0_u14_u3_n141 ) , .A1( u0_u14_u3_n169 ) );
  OAI222_X1 u0_u14_u3_U32 (.C2( u0_u14_u3_n107 ) , .A2( u0_u14_u3_n108 ) , .B1( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n138 ) , .B2( u0_u14_u3_n146 ) , .C1( u0_u14_u3_n154 ) , .A1( u0_u14_u3_n164 ) );
  NOR4_X1 u0_u14_u3_U33 (.A4( u0_u14_u3_n157 ) , .A3( u0_u14_u3_n158 ) , .A2( u0_u14_u3_n159 ) , .A1( u0_u14_u3_n160 ) , .ZN( u0_u14_u3_n161 ) );
  AOI21_X1 u0_u14_u3_U34 (.B2( u0_u14_u3_n152 ) , .B1( u0_u14_u3_n153 ) , .ZN( u0_u14_u3_n158 ) , .A( u0_u14_u3_n164 ) );
  AOI21_X1 u0_u14_u3_U35 (.A( u0_u14_u3_n154 ) , .B2( u0_u14_u3_n155 ) , .B1( u0_u14_u3_n156 ) , .ZN( u0_u14_u3_n157 ) );
  AOI21_X1 u0_u14_u3_U36 (.A( u0_u14_u3_n149 ) , .B2( u0_u14_u3_n150 ) , .B1( u0_u14_u3_n151 ) , .ZN( u0_u14_u3_n159 ) );
  AOI211_X1 u0_u14_u3_U37 (.ZN( u0_u14_u3_n109 ) , .A( u0_u14_u3_n119 ) , .C2( u0_u14_u3_n129 ) , .B( u0_u14_u3_n138 ) , .C1( u0_u14_u3_n141 ) );
  AOI211_X1 u0_u14_u3_U38 (.B( u0_u14_u3_n119 ) , .A( u0_u14_u3_n120 ) , .C2( u0_u14_u3_n121 ) , .ZN( u0_u14_u3_n122 ) , .C1( u0_u14_u3_n179 ) );
  INV_X1 u0_u14_u3_U39 (.A( u0_u14_u3_n156 ) , .ZN( u0_u14_u3_n179 ) );
  INV_X1 u0_u14_u3_U4 (.A( u0_u14_u3_n140 ) , .ZN( u0_u14_u3_n182 ) );
  OAI22_X1 u0_u14_u3_U40 (.B1( u0_u14_u3_n118 ) , .ZN( u0_u14_u3_n120 ) , .A1( u0_u14_u3_n135 ) , .B2( u0_u14_u3_n154 ) , .A2( u0_u14_u3_n178 ) );
  AND3_X1 u0_u14_u3_U41 (.ZN( u0_u14_u3_n118 ) , .A2( u0_u14_u3_n124 ) , .A1( u0_u14_u3_n144 ) , .A3( u0_u14_u3_n152 ) );
  INV_X1 u0_u14_u3_U42 (.A( u0_u14_u3_n121 ) , .ZN( u0_u14_u3_n164 ) );
  NAND2_X1 u0_u14_u3_U43 (.ZN( u0_u14_u3_n133 ) , .A1( u0_u14_u3_n154 ) , .A2( u0_u14_u3_n164 ) );
  OAI211_X1 u0_u14_u3_U44 (.B( u0_u14_u3_n127 ) , .ZN( u0_u14_u3_n139 ) , .C1( u0_u14_u3_n150 ) , .C2( u0_u14_u3_n154 ) , .A( u0_u14_u3_n184 ) );
  INV_X1 u0_u14_u3_U45 (.A( u0_u14_u3_n125 ) , .ZN( u0_u14_u3_n184 ) );
  AOI221_X1 u0_u14_u3_U46 (.A( u0_u14_u3_n126 ) , .ZN( u0_u14_u3_n127 ) , .C2( u0_u14_u3_n132 ) , .C1( u0_u14_u3_n169 ) , .B2( u0_u14_u3_n170 ) , .B1( u0_u14_u3_n174 ) );
  OAI22_X1 u0_u14_u3_U47 (.A1( u0_u14_u3_n124 ) , .ZN( u0_u14_u3_n125 ) , .B2( u0_u14_u3_n145 ) , .A2( u0_u14_u3_n165 ) , .B1( u0_u14_u3_n167 ) );
  NOR2_X1 u0_u14_u3_U48 (.A1( u0_u14_u3_n113 ) , .ZN( u0_u14_u3_n131 ) , .A2( u0_u14_u3_n154 ) );
  NAND2_X1 u0_u14_u3_U49 (.A1( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n150 ) , .A2( u0_u14_u3_n99 ) );
  INV_X1 u0_u14_u3_U5 (.A( u0_u14_u3_n117 ) , .ZN( u0_u14_u3_n178 ) );
  NAND2_X1 u0_u14_u3_U50 (.A2( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n155 ) , .A1( u0_u14_u3_n97 ) );
  INV_X1 u0_u14_u3_U51 (.A( u0_u14_u3_n141 ) , .ZN( u0_u14_u3_n167 ) );
  AOI21_X1 u0_u14_u3_U52 (.B2( u0_u14_u3_n114 ) , .B1( u0_u14_u3_n146 ) , .A( u0_u14_u3_n154 ) , .ZN( u0_u14_u3_n94 ) );
  AOI21_X1 u0_u14_u3_U53 (.ZN( u0_u14_u3_n110 ) , .B2( u0_u14_u3_n142 ) , .B1( u0_u14_u3_n186 ) , .A( u0_u14_u3_n95 ) );
  INV_X1 u0_u14_u3_U54 (.A( u0_u14_u3_n145 ) , .ZN( u0_u14_u3_n186 ) );
  AOI21_X1 u0_u14_u3_U55 (.B1( u0_u14_u3_n124 ) , .A( u0_u14_u3_n149 ) , .B2( u0_u14_u3_n155 ) , .ZN( u0_u14_u3_n95 ) );
  INV_X1 u0_u14_u3_U56 (.A( u0_u14_u3_n149 ) , .ZN( u0_u14_u3_n169 ) );
  NAND2_X1 u0_u14_u3_U57 (.ZN( u0_u14_u3_n124 ) , .A1( u0_u14_u3_n96 ) , .A2( u0_u14_u3_n97 ) );
  NAND2_X1 u0_u14_u3_U58 (.A2( u0_u14_u3_n100 ) , .ZN( u0_u14_u3_n146 ) , .A1( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U59 (.A1( u0_u14_u3_n101 ) , .ZN( u0_u14_u3_n145 ) , .A2( u0_u14_u3_n99 ) );
  AOI221_X1 u0_u14_u3_U6 (.A( u0_u14_u3_n131 ) , .C2( u0_u14_u3_n132 ) , .C1( u0_u14_u3_n133 ) , .ZN( u0_u14_u3_n134 ) , .B1( u0_u14_u3_n143 ) , .B2( u0_u14_u3_n177 ) );
  NAND2_X1 u0_u14_u3_U60 (.A1( u0_u14_u3_n100 ) , .ZN( u0_u14_u3_n156 ) , .A2( u0_u14_u3_n99 ) );
  NAND2_X1 u0_u14_u3_U61 (.A2( u0_u14_u3_n101 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n148 ) );
  NAND2_X1 u0_u14_u3_U62 (.A1( u0_u14_u3_n100 ) , .A2( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n128 ) );
  NAND2_X1 u0_u14_u3_U63 (.A2( u0_u14_u3_n101 ) , .A1( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n152 ) );
  NAND2_X1 u0_u14_u3_U64 (.A2( u0_u14_u3_n101 ) , .ZN( u0_u14_u3_n114 ) , .A1( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U65 (.ZN( u0_u14_u3_n107 ) , .A1( u0_u14_u3_n97 ) , .A2( u0_u14_u3_n99 ) );
  NAND2_X1 u0_u14_u3_U66 (.A2( u0_u14_u3_n100 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n113 ) );
  NAND2_X1 u0_u14_u3_U67 (.A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n153 ) , .A2( u0_u14_u3_n97 ) );
  NAND2_X1 u0_u14_u3_U68 (.A2( u0_u14_u3_n103 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n130 ) );
  NAND2_X1 u0_u14_u3_U69 (.A2( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n144 ) , .A1( u0_u14_u3_n96 ) );
  OAI22_X1 u0_u14_u3_U7 (.B2( u0_u14_u3_n147 ) , .A2( u0_u14_u3_n148 ) , .ZN( u0_u14_u3_n160 ) , .B1( u0_u14_u3_n165 ) , .A1( u0_u14_u3_n168 ) );
  NAND2_X1 u0_u14_u3_U70 (.A1( u0_u14_u3_n102 ) , .A2( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n108 ) );
  NOR2_X1 u0_u14_u3_U71 (.A2( u0_u14_X_19 ) , .A1( u0_u14_X_20 ) , .ZN( u0_u14_u3_n99 ) );
  NOR2_X1 u0_u14_u3_U72 (.A2( u0_u14_X_21 ) , .A1( u0_u14_X_24 ) , .ZN( u0_u14_u3_n103 ) );
  NOR2_X1 u0_u14_u3_U73 (.A2( u0_u14_X_24 ) , .A1( u0_u14_u3_n171 ) , .ZN( u0_u14_u3_n97 ) );
  NOR2_X1 u0_u14_u3_U74 (.A2( u0_u14_X_23 ) , .ZN( u0_u14_u3_n141 ) , .A1( u0_u14_u3_n166 ) );
  NOR2_X1 u0_u14_u3_U75 (.A2( u0_u14_X_19 ) , .A1( u0_u14_u3_n172 ) , .ZN( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U76 (.A1( u0_u14_X_22 ) , .A2( u0_u14_X_23 ) , .ZN( u0_u14_u3_n154 ) );
  NAND2_X1 u0_u14_u3_U77 (.A1( u0_u14_X_23 ) , .ZN( u0_u14_u3_n149 ) , .A2( u0_u14_u3_n166 ) );
  NOR2_X1 u0_u14_u3_U78 (.A2( u0_u14_X_22 ) , .A1( u0_u14_X_23 ) , .ZN( u0_u14_u3_n121 ) );
  AND2_X1 u0_u14_u3_U79 (.A1( u0_u14_X_24 ) , .ZN( u0_u14_u3_n101 ) , .A2( u0_u14_u3_n171 ) );
  AND3_X1 u0_u14_u3_U8 (.A3( u0_u14_u3_n144 ) , .A2( u0_u14_u3_n145 ) , .A1( u0_u14_u3_n146 ) , .ZN( u0_u14_u3_n147 ) );
  AND2_X1 u0_u14_u3_U80 (.A1( u0_u14_X_19 ) , .ZN( u0_u14_u3_n102 ) , .A2( u0_u14_u3_n172 ) );
  AND2_X1 u0_u14_u3_U81 (.A1( u0_u14_X_21 ) , .A2( u0_u14_X_24 ) , .ZN( u0_u14_u3_n100 ) );
  AND2_X1 u0_u14_u3_U82 (.A2( u0_u14_X_19 ) , .A1( u0_u14_X_20 ) , .ZN( u0_u14_u3_n104 ) );
  INV_X1 u0_u14_u3_U83 (.A( u0_u14_X_22 ) , .ZN( u0_u14_u3_n166 ) );
  INV_X1 u0_u14_u3_U84 (.A( u0_u14_X_21 ) , .ZN( u0_u14_u3_n171 ) );
  INV_X1 u0_u14_u3_U85 (.A( u0_u14_X_20 ) , .ZN( u0_u14_u3_n172 ) );
  NAND4_X1 u0_u14_u3_U86 (.ZN( u0_out14_26 ) , .A4( u0_u14_u3_n109 ) , .A3( u0_u14_u3_n110 ) , .A2( u0_u14_u3_n111 ) , .A1( u0_u14_u3_n173 ) );
  INV_X1 u0_u14_u3_U87 (.ZN( u0_u14_u3_n173 ) , .A( u0_u14_u3_n94 ) );
  OAI21_X1 u0_u14_u3_U88 (.ZN( u0_u14_u3_n111 ) , .B2( u0_u14_u3_n117 ) , .A( u0_u14_u3_n133 ) , .B1( u0_u14_u3_n176 ) );
  NAND4_X1 u0_u14_u3_U89 (.ZN( u0_out14_20 ) , .A4( u0_u14_u3_n122 ) , .A3( u0_u14_u3_n123 ) , .A1( u0_u14_u3_n175 ) , .A2( u0_u14_u3_n180 ) );
  INV_X1 u0_u14_u3_U9 (.A( u0_u14_u3_n143 ) , .ZN( u0_u14_u3_n168 ) );
  INV_X1 u0_u14_u3_U90 (.A( u0_u14_u3_n126 ) , .ZN( u0_u14_u3_n180 ) );
  INV_X1 u0_u14_u3_U91 (.A( u0_u14_u3_n112 ) , .ZN( u0_u14_u3_n175 ) );
  NAND4_X1 u0_u14_u3_U92 (.ZN( u0_out14_1 ) , .A4( u0_u14_u3_n161 ) , .A3( u0_u14_u3_n162 ) , .A2( u0_u14_u3_n163 ) , .A1( u0_u14_u3_n185 ) );
  NAND2_X1 u0_u14_u3_U93 (.ZN( u0_u14_u3_n163 ) , .A2( u0_u14_u3_n170 ) , .A1( u0_u14_u3_n176 ) );
  AOI22_X1 u0_u14_u3_U94 (.B2( u0_u14_u3_n140 ) , .B1( u0_u14_u3_n141 ) , .A2( u0_u14_u3_n142 ) , .ZN( u0_u14_u3_n162 ) , .A1( u0_u14_u3_n177 ) );
  OR4_X1 u0_u14_u3_U95 (.ZN( u0_out14_10 ) , .A4( u0_u14_u3_n136 ) , .A3( u0_u14_u3_n137 ) , .A1( u0_u14_u3_n138 ) , .A2( u0_u14_u3_n139 ) );
  OAI222_X1 u0_u14_u3_U96 (.C1( u0_u14_u3_n128 ) , .ZN( u0_u14_u3_n137 ) , .B1( u0_u14_u3_n148 ) , .A2( u0_u14_u3_n150 ) , .B2( u0_u14_u3_n154 ) , .C2( u0_u14_u3_n164 ) , .A1( u0_u14_u3_n167 ) );
  OAI221_X1 u0_u14_u3_U97 (.A( u0_u14_u3_n134 ) , .B2( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n136 ) , .C1( u0_u14_u3_n149 ) , .B1( u0_u14_u3_n151 ) , .C2( u0_u14_u3_n183 ) );
  NAND3_X1 u0_u14_u3_U98 (.A1( u0_u14_u3_n114 ) , .ZN( u0_u14_u3_n115 ) , .A2( u0_u14_u3_n145 ) , .A3( u0_u14_u3_n153 ) );
  NAND3_X1 u0_u14_u3_U99 (.ZN( u0_u14_u3_n129 ) , .A2( u0_u14_u3_n144 ) , .A1( u0_u14_u3_n153 ) , .A3( u0_u14_u3_n182 ) );
  XOR2_X1 u0_u15_U14 (.A( u0_FP_60 ) , .B( u0_K16_41 ) , .Z( u0_u15_X_41 ) );
  XOR2_X1 u0_u15_U15 (.A( u0_FP_59 ) , .B( u0_K16_40 ) , .Z( u0_u15_X_40 ) );
  XOR2_X1 u0_u15_U17 (.A( u0_FP_58 ) , .B( u0_K16_39 ) , .Z( u0_u15_X_39 ) );
  XOR2_X1 u0_u15_U18 (.A( u0_FP_57 ) , .B( u0_K16_38 ) , .Z( u0_u15_X_38 ) );
  XOR2_X1 u0_u15_U19 (.A( u0_FP_56 ) , .B( u0_K16_37 ) , .Z( u0_u15_X_37 ) );
  INV_X1 u0_u15_u6_U10 (.ZN( u0_u15_u6_n172 ) , .A( u0_u15_u6_n88 ) );
  OAI21_X1 u0_u15_u6_U11 (.A( u0_u15_u6_n159 ) , .B1( u0_u15_u6_n169 ) , .B2( u0_u15_u6_n173 ) , .ZN( u0_u15_u6_n90 ) );
  AOI22_X1 u0_u15_u6_U12 (.A2( u0_u15_u6_n151 ) , .B2( u0_u15_u6_n161 ) , .A1( u0_u15_u6_n167 ) , .B1( u0_u15_u6_n170 ) , .ZN( u0_u15_u6_n89 ) );
  AOI21_X1 u0_u15_u6_U13 (.ZN( u0_u15_u6_n106 ) , .A( u0_u15_u6_n142 ) , .B2( u0_u15_u6_n159 ) , .B1( u0_u15_u6_n164 ) );
  INV_X1 u0_u15_u6_U14 (.A( u0_u15_u6_n155 ) , .ZN( u0_u15_u6_n161 ) );
  INV_X1 u0_u15_u6_U15 (.A( u0_u15_u6_n128 ) , .ZN( u0_u15_u6_n164 ) );
  NAND2_X1 u0_u15_u6_U16 (.ZN( u0_u15_u6_n110 ) , .A1( u0_u15_u6_n122 ) , .A2( u0_u15_u6_n129 ) );
  NAND2_X1 u0_u15_u6_U17 (.ZN( u0_u15_u6_n124 ) , .A2( u0_u15_u6_n146 ) , .A1( u0_u15_u6_n148 ) );
  INV_X1 u0_u15_u6_U18 (.A( u0_u15_u6_n132 ) , .ZN( u0_u15_u6_n171 ) );
  AND2_X1 u0_u15_u6_U19 (.A1( u0_u15_u6_n100 ) , .ZN( u0_u15_u6_n130 ) , .A2( u0_u15_u6_n147 ) );
  INV_X1 u0_u15_u6_U20 (.A( u0_u15_u6_n127 ) , .ZN( u0_u15_u6_n173 ) );
  INV_X1 u0_u15_u6_U21 (.A( u0_u15_u6_n121 ) , .ZN( u0_u15_u6_n167 ) );
  INV_X1 u0_u15_u6_U22 (.A( u0_u15_u6_n100 ) , .ZN( u0_u15_u6_n169 ) );
  INV_X1 u0_u15_u6_U23 (.A( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n170 ) );
  INV_X1 u0_u15_u6_U24 (.A( u0_u15_u6_n113 ) , .ZN( u0_u15_u6_n168 ) );
  AND2_X1 u0_u15_u6_U25 (.A1( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n119 ) , .ZN( u0_u15_u6_n133 ) );
  AND2_X1 u0_u15_u6_U26 (.A2( u0_u15_u6_n121 ) , .A1( u0_u15_u6_n122 ) , .ZN( u0_u15_u6_n131 ) );
  AND3_X1 u0_u15_u6_U27 (.ZN( u0_u15_u6_n120 ) , .A2( u0_u15_u6_n127 ) , .A1( u0_u15_u6_n132 ) , .A3( u0_u15_u6_n145 ) );
  INV_X1 u0_u15_u6_U28 (.A( u0_u15_u6_n146 ) , .ZN( u0_u15_u6_n163 ) );
  AOI222_X1 u0_u15_u6_U29 (.ZN( u0_u15_u6_n114 ) , .A1( u0_u15_u6_n118 ) , .A2( u0_u15_u6_n126 ) , .B2( u0_u15_u6_n151 ) , .C2( u0_u15_u6_n159 ) , .C1( u0_u15_u6_n168 ) , .B1( u0_u15_u6_n169 ) );
  INV_X1 u0_u15_u6_U3 (.A( u0_u15_u6_n110 ) , .ZN( u0_u15_u6_n166 ) );
  NOR2_X1 u0_u15_u6_U30 (.A1( u0_u15_u6_n162 ) , .A2( u0_u15_u6_n165 ) , .ZN( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U31 (.A1( u0_u15_u6_n144 ) , .ZN( u0_u15_u6_n151 ) , .A2( u0_u15_u6_n158 ) );
  NAND2_X1 u0_u15_u6_U32 (.ZN( u0_u15_u6_n132 ) , .A1( u0_u15_u6_n91 ) , .A2( u0_u15_u6_n97 ) );
  AOI22_X1 u0_u15_u6_U33 (.B2( u0_u15_u6_n110 ) , .B1( u0_u15_u6_n111 ) , .A1( u0_u15_u6_n112 ) , .ZN( u0_u15_u6_n115 ) , .A2( u0_u15_u6_n161 ) );
  NAND4_X1 u0_u15_u6_U34 (.A3( u0_u15_u6_n109 ) , .ZN( u0_u15_u6_n112 ) , .A4( u0_u15_u6_n132 ) , .A2( u0_u15_u6_n147 ) , .A1( u0_u15_u6_n166 ) );
  NOR2_X1 u0_u15_u6_U35 (.ZN( u0_u15_u6_n109 ) , .A1( u0_u15_u6_n170 ) , .A2( u0_u15_u6_n173 ) );
  NOR2_X1 u0_u15_u6_U36 (.A2( u0_u15_u6_n126 ) , .ZN( u0_u15_u6_n155 ) , .A1( u0_u15_u6_n160 ) );
  NAND2_X1 u0_u15_u6_U37 (.ZN( u0_u15_u6_n146 ) , .A2( u0_u15_u6_n94 ) , .A1( u0_u15_u6_n99 ) );
  AOI21_X1 u0_u15_u6_U38 (.A( u0_u15_u6_n144 ) , .B2( u0_u15_u6_n145 ) , .B1( u0_u15_u6_n146 ) , .ZN( u0_u15_u6_n150 ) );
  AOI211_X1 u0_u15_u6_U39 (.B( u0_u15_u6_n134 ) , .A( u0_u15_u6_n135 ) , .C1( u0_u15_u6_n136 ) , .ZN( u0_u15_u6_n137 ) , .C2( u0_u15_u6_n151 ) );
  INV_X1 u0_u15_u6_U4 (.A( u0_u15_u6_n142 ) , .ZN( u0_u15_u6_n174 ) );
  NAND4_X1 u0_u15_u6_U40 (.A4( u0_u15_u6_n127 ) , .A3( u0_u15_u6_n128 ) , .A2( u0_u15_u6_n129 ) , .A1( u0_u15_u6_n130 ) , .ZN( u0_u15_u6_n136 ) );
  AOI21_X1 u0_u15_u6_U41 (.B2( u0_u15_u6_n132 ) , .B1( u0_u15_u6_n133 ) , .ZN( u0_u15_u6_n134 ) , .A( u0_u15_u6_n158 ) );
  AOI21_X1 u0_u15_u6_U42 (.B1( u0_u15_u6_n131 ) , .ZN( u0_u15_u6_n135 ) , .A( u0_u15_u6_n144 ) , .B2( u0_u15_u6_n146 ) );
  INV_X1 u0_u15_u6_U43 (.A( u0_u15_u6_n111 ) , .ZN( u0_u15_u6_n158 ) );
  NAND2_X1 u0_u15_u6_U44 (.ZN( u0_u15_u6_n127 ) , .A1( u0_u15_u6_n91 ) , .A2( u0_u15_u6_n92 ) );
  NAND2_X1 u0_u15_u6_U45 (.ZN( u0_u15_u6_n129 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n96 ) );
  INV_X1 u0_u15_u6_U46 (.A( u0_u15_u6_n144 ) , .ZN( u0_u15_u6_n159 ) );
  NAND2_X1 u0_u15_u6_U47 (.ZN( u0_u15_u6_n145 ) , .A2( u0_u15_u6_n97 ) , .A1( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U48 (.ZN( u0_u15_u6_n148 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n94 ) );
  NAND2_X1 u0_u15_u6_U49 (.ZN( u0_u15_u6_n108 ) , .A2( u0_u15_u6_n139 ) , .A1( u0_u15_u6_n144 ) );
  NAND2_X1 u0_u15_u6_U5 (.A2( u0_u15_u6_n143 ) , .ZN( u0_u15_u6_n152 ) , .A1( u0_u15_u6_n166 ) );
  NAND2_X1 u0_u15_u6_U50 (.ZN( u0_u15_u6_n121 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n97 ) );
  NAND2_X1 u0_u15_u6_U51 (.ZN( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n95 ) );
  AND2_X1 u0_u15_u6_U52 (.ZN( u0_u15_u6_n118 ) , .A2( u0_u15_u6_n91 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U53 (.ZN( u0_u15_u6_n147 ) , .A2( u0_u15_u6_n98 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U54 (.ZN( u0_u15_u6_n128 ) , .A1( u0_u15_u6_n94 ) , .A2( u0_u15_u6_n96 ) );
  NAND2_X1 u0_u15_u6_U55 (.ZN( u0_u15_u6_n119 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U56 (.ZN( u0_u15_u6_n123 ) , .A2( u0_u15_u6_n91 ) , .A1( u0_u15_u6_n96 ) );
  NAND2_X1 u0_u15_u6_U57 (.ZN( u0_u15_u6_n100 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U58 (.ZN( u0_u15_u6_n122 ) , .A1( u0_u15_u6_n94 ) , .A2( u0_u15_u6_n97 ) );
  INV_X1 u0_u15_u6_U59 (.A( u0_u15_u6_n139 ) , .ZN( u0_u15_u6_n160 ) );
  AOI22_X1 u0_u15_u6_U6 (.B2( u0_u15_u6_n101 ) , .A1( u0_u15_u6_n102 ) , .ZN( u0_u15_u6_n103 ) , .B1( u0_u15_u6_n160 ) , .A2( u0_u15_u6_n161 ) );
  NAND2_X1 u0_u15_u6_U60 (.ZN( u0_u15_u6_n113 ) , .A1( u0_u15_u6_n96 ) , .A2( u0_u15_u6_n98 ) );
  NOR2_X1 u0_u15_u6_U61 (.A2( u0_u15_X_40 ) , .A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n126 ) );
  NOR2_X1 u0_u15_u6_U62 (.A2( u0_u15_X_39 ) , .A1( u0_u15_X_42 ) , .ZN( u0_u15_u6_n92 ) );
  NOR2_X1 u0_u15_u6_U63 (.A2( u0_u15_X_39 ) , .A1( u0_u15_u6_n156 ) , .ZN( u0_u15_u6_n97 ) );
  NOR2_X1 u0_u15_u6_U64 (.A2( u0_u15_X_38 ) , .A1( u0_u15_u6_n165 ) , .ZN( u0_u15_u6_n95 ) );
  NOR2_X1 u0_u15_u6_U65 (.A2( u0_u15_X_41 ) , .ZN( u0_u15_u6_n111 ) , .A1( u0_u15_u6_n157 ) );
  NOR2_X1 u0_u15_u6_U66 (.A2( u0_u15_X_37 ) , .A1( u0_u15_u6_n162 ) , .ZN( u0_u15_u6_n94 ) );
  NOR2_X1 u0_u15_u6_U67 (.A2( u0_u15_X_37 ) , .A1( u0_u15_X_38 ) , .ZN( u0_u15_u6_n91 ) );
  NAND2_X1 u0_u15_u6_U68 (.A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n144 ) , .A2( u0_u15_u6_n157 ) );
  NAND2_X1 u0_u15_u6_U69 (.A2( u0_u15_X_40 ) , .A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n139 ) );
  NOR2_X1 u0_u15_u6_U7 (.A1( u0_u15_u6_n118 ) , .ZN( u0_u15_u6_n143 ) , .A2( u0_u15_u6_n168 ) );
  AND2_X1 u0_u15_u6_U70 (.A1( u0_u15_X_39 ) , .A2( u0_u15_u6_n156 ) , .ZN( u0_u15_u6_n96 ) );
  AND2_X1 u0_u15_u6_U71 (.A1( u0_u15_X_39 ) , .A2( u0_u15_X_42 ) , .ZN( u0_u15_u6_n99 ) );
  INV_X1 u0_u15_u6_U72 (.A( u0_u15_X_40 ) , .ZN( u0_u15_u6_n157 ) );
  INV_X1 u0_u15_u6_U73 (.A( u0_u15_X_37 ) , .ZN( u0_u15_u6_n165 ) );
  INV_X1 u0_u15_u6_U74 (.A( u0_u15_X_38 ) , .ZN( u0_u15_u6_n162 ) );
  INV_X1 u0_u15_u6_U75 (.A( u0_u15_X_42 ) , .ZN( u0_u15_u6_n156 ) );
  NAND4_X1 u0_u15_u6_U76 (.ZN( u0_out15_12 ) , .A4( u0_u15_u6_n114 ) , .A3( u0_u15_u6_n115 ) , .A2( u0_u15_u6_n116 ) , .A1( u0_u15_u6_n117 ) );
  OAI22_X1 u0_u15_u6_U77 (.B2( u0_u15_u6_n111 ) , .ZN( u0_u15_u6_n116 ) , .B1( u0_u15_u6_n126 ) , .A2( u0_u15_u6_n164 ) , .A1( u0_u15_u6_n167 ) );
  OAI21_X1 u0_u15_u6_U78 (.A( u0_u15_u6_n108 ) , .ZN( u0_u15_u6_n117 ) , .B2( u0_u15_u6_n141 ) , .B1( u0_u15_u6_n163 ) );
  NAND4_X1 u0_u15_u6_U79 (.ZN( u0_out15_32 ) , .A4( u0_u15_u6_n103 ) , .A3( u0_u15_u6_n104 ) , .A2( u0_u15_u6_n105 ) , .A1( u0_u15_u6_n106 ) );
  AOI21_X1 u0_u15_u6_U8 (.B1( u0_u15_u6_n107 ) , .B2( u0_u15_u6_n132 ) , .A( u0_u15_u6_n158 ) , .ZN( u0_u15_u6_n88 ) );
  AOI22_X1 u0_u15_u6_U80 (.ZN( u0_u15_u6_n105 ) , .A2( u0_u15_u6_n108 ) , .A1( u0_u15_u6_n118 ) , .B2( u0_u15_u6_n126 ) , .B1( u0_u15_u6_n171 ) );
  AOI22_X1 u0_u15_u6_U81 (.ZN( u0_u15_u6_n104 ) , .A1( u0_u15_u6_n111 ) , .B1( u0_u15_u6_n124 ) , .B2( u0_u15_u6_n151 ) , .A2( u0_u15_u6_n93 ) );
  OAI211_X1 u0_u15_u6_U82 (.ZN( u0_out15_22 ) , .B( u0_u15_u6_n137 ) , .A( u0_u15_u6_n138 ) , .C2( u0_u15_u6_n139 ) , .C1( u0_u15_u6_n140 ) );
  AOI22_X1 u0_u15_u6_U83 (.B1( u0_u15_u6_n124 ) , .A2( u0_u15_u6_n125 ) , .A1( u0_u15_u6_n126 ) , .ZN( u0_u15_u6_n138 ) , .B2( u0_u15_u6_n161 ) );
  AND4_X1 u0_u15_u6_U84 (.A3( u0_u15_u6_n119 ) , .A1( u0_u15_u6_n120 ) , .A4( u0_u15_u6_n129 ) , .ZN( u0_u15_u6_n140 ) , .A2( u0_u15_u6_n143 ) );
  OAI211_X1 u0_u15_u6_U85 (.ZN( u0_out15_7 ) , .B( u0_u15_u6_n153 ) , .C2( u0_u15_u6_n154 ) , .C1( u0_u15_u6_n155 ) , .A( u0_u15_u6_n174 ) );
  NOR3_X1 u0_u15_u6_U86 (.A1( u0_u15_u6_n141 ) , .ZN( u0_u15_u6_n154 ) , .A3( u0_u15_u6_n164 ) , .A2( u0_u15_u6_n171 ) );
  AOI211_X1 u0_u15_u6_U87 (.B( u0_u15_u6_n149 ) , .A( u0_u15_u6_n150 ) , .C2( u0_u15_u6_n151 ) , .C1( u0_u15_u6_n152 ) , .ZN( u0_u15_u6_n153 ) );
  NAND3_X1 u0_u15_u6_U88 (.A2( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n125 ) , .A1( u0_u15_u6_n130 ) , .A3( u0_u15_u6_n131 ) );
  NAND3_X1 u0_u15_u6_U89 (.A3( u0_u15_u6_n133 ) , .ZN( u0_u15_u6_n141 ) , .A1( u0_u15_u6_n145 ) , .A2( u0_u15_u6_n148 ) );
  AOI21_X1 u0_u15_u6_U9 (.B2( u0_u15_u6_n147 ) , .B1( u0_u15_u6_n148 ) , .ZN( u0_u15_u6_n149 ) , .A( u0_u15_u6_n158 ) );
  NAND3_X1 u0_u15_u6_U90 (.ZN( u0_u15_u6_n101 ) , .A3( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n121 ) , .A1( u0_u15_u6_n127 ) );
  NAND3_X1 u0_u15_u6_U91 (.ZN( u0_u15_u6_n102 ) , .A3( u0_u15_u6_n130 ) , .A2( u0_u15_u6_n145 ) , .A1( u0_u15_u6_n166 ) );
  NAND3_X1 u0_u15_u6_U92 (.A3( u0_u15_u6_n113 ) , .A1( u0_u15_u6_n119 ) , .A2( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n93 ) );
  NAND3_X1 u0_u15_u6_U93 (.ZN( u0_u15_u6_n142 ) , .A2( u0_u15_u6_n172 ) , .A3( u0_u15_u6_n89 ) , .A1( u0_u15_u6_n90 ) );
  XOR2_X1 u0_u1_U14 (.B( u0_K2_41 ) , .A( u0_R0_28 ) , .Z( u0_u1_X_41 ) );
  XOR2_X1 u0_u1_U24 (.B( u0_K2_32 ) , .A( u0_R0_21 ) , .Z( u0_u1_X_32 ) );
  XOR2_X1 u0_u1_U25 (.B( u0_K2_31 ) , .A( u0_R0_20 ) , .Z( u0_u1_X_31 ) );
  XOR2_X1 u0_u1_U26 (.B( u0_K2_30 ) , .A( u0_R0_21 ) , .Z( u0_u1_X_30 ) );
  XOR2_X1 u0_u1_U28 (.B( u0_K2_29 ) , .A( u0_R0_20 ) , .Z( u0_u1_X_29 ) );
  XOR2_X1 u0_u1_U29 (.B( u0_K2_28 ) , .A( u0_R0_19 ) , .Z( u0_u1_X_28 ) );
  XOR2_X1 u0_u1_U30 (.B( u0_K2_27 ) , .A( u0_R0_18 ) , .Z( u0_u1_X_27 ) );
  OAI22_X1 u0_u1_u4_U10 (.B2( u0_u1_u4_n135 ) , .ZN( u0_u1_u4_n137 ) , .B1( u0_u1_u4_n153 ) , .A1( u0_u1_u4_n155 ) , .A2( u0_u1_u4_n171 ) );
  AND3_X1 u0_u1_u4_U11 (.A2( u0_u1_u4_n134 ) , .ZN( u0_u1_u4_n135 ) , .A3( u0_u1_u4_n145 ) , .A1( u0_u1_u4_n157 ) );
  NAND2_X1 u0_u1_u4_U12 (.ZN( u0_u1_u4_n132 ) , .A2( u0_u1_u4_n170 ) , .A1( u0_u1_u4_n173 ) );
  AOI21_X1 u0_u1_u4_U13 (.B2( u0_u1_u4_n160 ) , .B1( u0_u1_u4_n161 ) , .ZN( u0_u1_u4_n162 ) , .A( u0_u1_u4_n170 ) );
  AOI21_X1 u0_u1_u4_U14 (.ZN( u0_u1_u4_n107 ) , .B2( u0_u1_u4_n143 ) , .A( u0_u1_u4_n174 ) , .B1( u0_u1_u4_n184 ) );
  AOI21_X1 u0_u1_u4_U15 (.B2( u0_u1_u4_n158 ) , .B1( u0_u1_u4_n159 ) , .ZN( u0_u1_u4_n163 ) , .A( u0_u1_u4_n174 ) );
  AOI21_X1 u0_u1_u4_U16 (.A( u0_u1_u4_n153 ) , .B2( u0_u1_u4_n154 ) , .B1( u0_u1_u4_n155 ) , .ZN( u0_u1_u4_n165 ) );
  AOI21_X1 u0_u1_u4_U17 (.A( u0_u1_u4_n156 ) , .B2( u0_u1_u4_n157 ) , .ZN( u0_u1_u4_n164 ) , .B1( u0_u1_u4_n184 ) );
  INV_X1 u0_u1_u4_U18 (.A( u0_u1_u4_n138 ) , .ZN( u0_u1_u4_n170 ) );
  AND2_X1 u0_u1_u4_U19 (.A2( u0_u1_u4_n120 ) , .ZN( u0_u1_u4_n155 ) , .A1( u0_u1_u4_n160 ) );
  INV_X1 u0_u1_u4_U20 (.A( u0_u1_u4_n156 ) , .ZN( u0_u1_u4_n175 ) );
  NAND2_X1 u0_u1_u4_U21 (.A2( u0_u1_u4_n118 ) , .ZN( u0_u1_u4_n131 ) , .A1( u0_u1_u4_n147 ) );
  NAND2_X1 u0_u1_u4_U22 (.A1( u0_u1_u4_n119 ) , .A2( u0_u1_u4_n120 ) , .ZN( u0_u1_u4_n130 ) );
  NAND2_X1 u0_u1_u4_U23 (.ZN( u0_u1_u4_n117 ) , .A2( u0_u1_u4_n118 ) , .A1( u0_u1_u4_n148 ) );
  NAND2_X1 u0_u1_u4_U24 (.ZN( u0_u1_u4_n129 ) , .A1( u0_u1_u4_n134 ) , .A2( u0_u1_u4_n148 ) );
  AND3_X1 u0_u1_u4_U25 (.A1( u0_u1_u4_n119 ) , .A2( u0_u1_u4_n143 ) , .A3( u0_u1_u4_n154 ) , .ZN( u0_u1_u4_n161 ) );
  AND2_X1 u0_u1_u4_U26 (.A1( u0_u1_u4_n145 ) , .A2( u0_u1_u4_n147 ) , .ZN( u0_u1_u4_n159 ) );
  OR3_X1 u0_u1_u4_U27 (.A3( u0_u1_u4_n114 ) , .A2( u0_u1_u4_n115 ) , .A1( u0_u1_u4_n116 ) , .ZN( u0_u1_u4_n136 ) );
  AOI21_X1 u0_u1_u4_U28 (.A( u0_u1_u4_n113 ) , .ZN( u0_u1_u4_n116 ) , .B2( u0_u1_u4_n173 ) , .B1( u0_u1_u4_n174 ) );
  AOI21_X1 u0_u1_u4_U29 (.ZN( u0_u1_u4_n115 ) , .B2( u0_u1_u4_n145 ) , .B1( u0_u1_u4_n146 ) , .A( u0_u1_u4_n156 ) );
  NOR2_X1 u0_u1_u4_U3 (.ZN( u0_u1_u4_n121 ) , .A1( u0_u1_u4_n181 ) , .A2( u0_u1_u4_n182 ) );
  OAI22_X1 u0_u1_u4_U30 (.ZN( u0_u1_u4_n114 ) , .A2( u0_u1_u4_n121 ) , .B1( u0_u1_u4_n160 ) , .B2( u0_u1_u4_n170 ) , .A1( u0_u1_u4_n171 ) );
  INV_X1 u0_u1_u4_U31 (.A( u0_u1_u4_n158 ) , .ZN( u0_u1_u4_n182 ) );
  INV_X1 u0_u1_u4_U32 (.ZN( u0_u1_u4_n181 ) , .A( u0_u1_u4_n96 ) );
  INV_X1 u0_u1_u4_U33 (.A( u0_u1_u4_n144 ) , .ZN( u0_u1_u4_n179 ) );
  INV_X1 u0_u1_u4_U34 (.A( u0_u1_u4_n157 ) , .ZN( u0_u1_u4_n178 ) );
  NAND2_X1 u0_u1_u4_U35 (.A2( u0_u1_u4_n154 ) , .A1( u0_u1_u4_n96 ) , .ZN( u0_u1_u4_n97 ) );
  INV_X1 u0_u1_u4_U36 (.ZN( u0_u1_u4_n186 ) , .A( u0_u1_u4_n95 ) );
  OAI221_X1 u0_u1_u4_U37 (.C1( u0_u1_u4_n134 ) , .B1( u0_u1_u4_n158 ) , .B2( u0_u1_u4_n171 ) , .C2( u0_u1_u4_n173 ) , .A( u0_u1_u4_n94 ) , .ZN( u0_u1_u4_n95 ) );
  AOI222_X1 u0_u1_u4_U38 (.B2( u0_u1_u4_n132 ) , .A1( u0_u1_u4_n138 ) , .C2( u0_u1_u4_n175 ) , .A2( u0_u1_u4_n179 ) , .C1( u0_u1_u4_n181 ) , .B1( u0_u1_u4_n185 ) , .ZN( u0_u1_u4_n94 ) );
  INV_X1 u0_u1_u4_U39 (.A( u0_u1_u4_n113 ) , .ZN( u0_u1_u4_n185 ) );
  INV_X1 u0_u1_u4_U4 (.A( u0_u1_u4_n117 ) , .ZN( u0_u1_u4_n184 ) );
  INV_X1 u0_u1_u4_U40 (.A( u0_u1_u4_n143 ) , .ZN( u0_u1_u4_n183 ) );
  NOR2_X1 u0_u1_u4_U41 (.ZN( u0_u1_u4_n138 ) , .A1( u0_u1_u4_n168 ) , .A2( u0_u1_u4_n169 ) );
  NOR2_X1 u0_u1_u4_U42 (.A1( u0_u1_u4_n150 ) , .A2( u0_u1_u4_n152 ) , .ZN( u0_u1_u4_n153 ) );
  NOR2_X1 u0_u1_u4_U43 (.A2( u0_u1_u4_n128 ) , .A1( u0_u1_u4_n138 ) , .ZN( u0_u1_u4_n156 ) );
  AOI22_X1 u0_u1_u4_U44 (.B2( u0_u1_u4_n122 ) , .A1( u0_u1_u4_n123 ) , .ZN( u0_u1_u4_n124 ) , .B1( u0_u1_u4_n128 ) , .A2( u0_u1_u4_n172 ) );
  NAND2_X1 u0_u1_u4_U45 (.A2( u0_u1_u4_n120 ) , .ZN( u0_u1_u4_n123 ) , .A1( u0_u1_u4_n161 ) );
  INV_X1 u0_u1_u4_U46 (.A( u0_u1_u4_n153 ) , .ZN( u0_u1_u4_n172 ) );
  AOI22_X1 u0_u1_u4_U47 (.B2( u0_u1_u4_n132 ) , .A2( u0_u1_u4_n133 ) , .ZN( u0_u1_u4_n140 ) , .A1( u0_u1_u4_n150 ) , .B1( u0_u1_u4_n179 ) );
  NAND2_X1 u0_u1_u4_U48 (.ZN( u0_u1_u4_n133 ) , .A2( u0_u1_u4_n146 ) , .A1( u0_u1_u4_n154 ) );
  NAND2_X1 u0_u1_u4_U49 (.A1( u0_u1_u4_n103 ) , .ZN( u0_u1_u4_n154 ) , .A2( u0_u1_u4_n98 ) );
  NOR4_X1 u0_u1_u4_U5 (.A4( u0_u1_u4_n106 ) , .A3( u0_u1_u4_n107 ) , .A2( u0_u1_u4_n108 ) , .A1( u0_u1_u4_n109 ) , .ZN( u0_u1_u4_n110 ) );
  NAND2_X1 u0_u1_u4_U50 (.A1( u0_u1_u4_n101 ) , .ZN( u0_u1_u4_n158 ) , .A2( u0_u1_u4_n99 ) );
  AOI21_X1 u0_u1_u4_U51 (.ZN( u0_u1_u4_n127 ) , .A( u0_u1_u4_n136 ) , .B2( u0_u1_u4_n150 ) , .B1( u0_u1_u4_n180 ) );
  INV_X1 u0_u1_u4_U52 (.A( u0_u1_u4_n160 ) , .ZN( u0_u1_u4_n180 ) );
  NAND2_X1 u0_u1_u4_U53 (.A2( u0_u1_u4_n104 ) , .A1( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n146 ) );
  NAND2_X1 u0_u1_u4_U54 (.A2( u0_u1_u4_n101 ) , .A1( u0_u1_u4_n102 ) , .ZN( u0_u1_u4_n160 ) );
  NAND2_X1 u0_u1_u4_U55 (.ZN( u0_u1_u4_n134 ) , .A1( u0_u1_u4_n98 ) , .A2( u0_u1_u4_n99 ) );
  NAND2_X1 u0_u1_u4_U56 (.A1( u0_u1_u4_n103 ) , .A2( u0_u1_u4_n104 ) , .ZN( u0_u1_u4_n143 ) );
  NAND2_X1 u0_u1_u4_U57 (.A2( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n145 ) , .A1( u0_u1_u4_n98 ) );
  NAND2_X1 u0_u1_u4_U58 (.A1( u0_u1_u4_n100 ) , .A2( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n120 ) );
  NAND2_X1 u0_u1_u4_U59 (.A1( u0_u1_u4_n102 ) , .A2( u0_u1_u4_n104 ) , .ZN( u0_u1_u4_n148 ) );
  AOI21_X1 u0_u1_u4_U6 (.ZN( u0_u1_u4_n106 ) , .B2( u0_u1_u4_n146 ) , .B1( u0_u1_u4_n158 ) , .A( u0_u1_u4_n170 ) );
  NAND2_X1 u0_u1_u4_U60 (.A2( u0_u1_u4_n100 ) , .A1( u0_u1_u4_n103 ) , .ZN( u0_u1_u4_n157 ) );
  INV_X1 u0_u1_u4_U61 (.A( u0_u1_u4_n150 ) , .ZN( u0_u1_u4_n173 ) );
  INV_X1 u0_u1_u4_U62 (.A( u0_u1_u4_n152 ) , .ZN( u0_u1_u4_n171 ) );
  NAND2_X1 u0_u1_u4_U63 (.A1( u0_u1_u4_n100 ) , .ZN( u0_u1_u4_n118 ) , .A2( u0_u1_u4_n99 ) );
  NAND2_X1 u0_u1_u4_U64 (.A2( u0_u1_u4_n100 ) , .A1( u0_u1_u4_n102 ) , .ZN( u0_u1_u4_n144 ) );
  NAND2_X1 u0_u1_u4_U65 (.A2( u0_u1_u4_n101 ) , .A1( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n96 ) );
  INV_X1 u0_u1_u4_U66 (.A( u0_u1_u4_n128 ) , .ZN( u0_u1_u4_n174 ) );
  NAND2_X1 u0_u1_u4_U67 (.A2( u0_u1_u4_n102 ) , .ZN( u0_u1_u4_n119 ) , .A1( u0_u1_u4_n98 ) );
  NAND2_X1 u0_u1_u4_U68 (.A2( u0_u1_u4_n101 ) , .A1( u0_u1_u4_n103 ) , .ZN( u0_u1_u4_n147 ) );
  NAND2_X1 u0_u1_u4_U69 (.A2( u0_u1_u4_n104 ) , .ZN( u0_u1_u4_n113 ) , .A1( u0_u1_u4_n99 ) );
  AOI21_X1 u0_u1_u4_U7 (.ZN( u0_u1_u4_n108 ) , .B2( u0_u1_u4_n134 ) , .B1( u0_u1_u4_n155 ) , .A( u0_u1_u4_n156 ) );
  NOR2_X1 u0_u1_u4_U70 (.A2( u0_u1_X_28 ) , .ZN( u0_u1_u4_n150 ) , .A1( u0_u1_u4_n168 ) );
  NOR2_X1 u0_u1_u4_U71 (.A2( u0_u1_X_29 ) , .ZN( u0_u1_u4_n152 ) , .A1( u0_u1_u4_n169 ) );
  NOR2_X1 u0_u1_u4_U72 (.A2( u0_u1_X_30 ) , .ZN( u0_u1_u4_n105 ) , .A1( u0_u1_u4_n176 ) );
  NOR2_X1 u0_u1_u4_U73 (.A2( u0_u1_X_26 ) , .ZN( u0_u1_u4_n100 ) , .A1( u0_u1_u4_n177 ) );
  NOR2_X1 u0_u1_u4_U74 (.A2( u0_u1_X_28 ) , .A1( u0_u1_X_29 ) , .ZN( u0_u1_u4_n128 ) );
  NOR2_X1 u0_u1_u4_U75 (.A2( u0_u1_X_27 ) , .A1( u0_u1_X_30 ) , .ZN( u0_u1_u4_n102 ) );
  NOR2_X1 u0_u1_u4_U76 (.A2( u0_u1_X_25 ) , .A1( u0_u1_X_26 ) , .ZN( u0_u1_u4_n98 ) );
  AND2_X1 u0_u1_u4_U77 (.A2( u0_u1_X_25 ) , .A1( u0_u1_X_26 ) , .ZN( u0_u1_u4_n104 ) );
  AND2_X1 u0_u1_u4_U78 (.A1( u0_u1_X_30 ) , .A2( u0_u1_u4_n176 ) , .ZN( u0_u1_u4_n99 ) );
  AND2_X1 u0_u1_u4_U79 (.A1( u0_u1_X_26 ) , .ZN( u0_u1_u4_n101 ) , .A2( u0_u1_u4_n177 ) );
  AOI21_X1 u0_u1_u4_U8 (.ZN( u0_u1_u4_n109 ) , .A( u0_u1_u4_n153 ) , .B1( u0_u1_u4_n159 ) , .B2( u0_u1_u4_n184 ) );
  AND2_X1 u0_u1_u4_U80 (.A1( u0_u1_X_27 ) , .A2( u0_u1_X_30 ) , .ZN( u0_u1_u4_n103 ) );
  INV_X1 u0_u1_u4_U81 (.A( u0_u1_X_28 ) , .ZN( u0_u1_u4_n169 ) );
  INV_X1 u0_u1_u4_U82 (.A( u0_u1_X_29 ) , .ZN( u0_u1_u4_n168 ) );
  INV_X1 u0_u1_u4_U83 (.A( u0_u1_X_25 ) , .ZN( u0_u1_u4_n177 ) );
  INV_X1 u0_u1_u4_U84 (.A( u0_u1_X_27 ) , .ZN( u0_u1_u4_n176 ) );
  NAND4_X1 u0_u1_u4_U85 (.ZN( u0_out1_25 ) , .A4( u0_u1_u4_n139 ) , .A3( u0_u1_u4_n140 ) , .A2( u0_u1_u4_n141 ) , .A1( u0_u1_u4_n142 ) );
  OAI21_X1 u0_u1_u4_U86 (.A( u0_u1_u4_n128 ) , .B2( u0_u1_u4_n129 ) , .B1( u0_u1_u4_n130 ) , .ZN( u0_u1_u4_n142 ) );
  OAI21_X1 u0_u1_u4_U87 (.B2( u0_u1_u4_n131 ) , .ZN( u0_u1_u4_n141 ) , .A( u0_u1_u4_n175 ) , .B1( u0_u1_u4_n183 ) );
  NAND4_X1 u0_u1_u4_U88 (.ZN( u0_out1_14 ) , .A4( u0_u1_u4_n124 ) , .A3( u0_u1_u4_n125 ) , .A2( u0_u1_u4_n126 ) , .A1( u0_u1_u4_n127 ) );
  AOI22_X1 u0_u1_u4_U89 (.B2( u0_u1_u4_n117 ) , .ZN( u0_u1_u4_n126 ) , .A1( u0_u1_u4_n129 ) , .B1( u0_u1_u4_n152 ) , .A2( u0_u1_u4_n175 ) );
  AOI211_X1 u0_u1_u4_U9 (.B( u0_u1_u4_n136 ) , .A( u0_u1_u4_n137 ) , .C2( u0_u1_u4_n138 ) , .ZN( u0_u1_u4_n139 ) , .C1( u0_u1_u4_n182 ) );
  AOI22_X1 u0_u1_u4_U90 (.ZN( u0_u1_u4_n125 ) , .B2( u0_u1_u4_n131 ) , .A2( u0_u1_u4_n132 ) , .B1( u0_u1_u4_n138 ) , .A1( u0_u1_u4_n178 ) );
  NAND4_X1 u0_u1_u4_U91 (.ZN( u0_out1_8 ) , .A4( u0_u1_u4_n110 ) , .A3( u0_u1_u4_n111 ) , .A2( u0_u1_u4_n112 ) , .A1( u0_u1_u4_n186 ) );
  NAND2_X1 u0_u1_u4_U92 (.ZN( u0_u1_u4_n112 ) , .A2( u0_u1_u4_n130 ) , .A1( u0_u1_u4_n150 ) );
  AOI22_X1 u0_u1_u4_U93 (.ZN( u0_u1_u4_n111 ) , .B2( u0_u1_u4_n132 ) , .A1( u0_u1_u4_n152 ) , .B1( u0_u1_u4_n178 ) , .A2( u0_u1_u4_n97 ) );
  AOI22_X1 u0_u1_u4_U94 (.B2( u0_u1_u4_n149 ) , .B1( u0_u1_u4_n150 ) , .A2( u0_u1_u4_n151 ) , .A1( u0_u1_u4_n152 ) , .ZN( u0_u1_u4_n167 ) );
  NOR4_X1 u0_u1_u4_U95 (.A4( u0_u1_u4_n162 ) , .A3( u0_u1_u4_n163 ) , .A2( u0_u1_u4_n164 ) , .A1( u0_u1_u4_n165 ) , .ZN( u0_u1_u4_n166 ) );
  NAND3_X1 u0_u1_u4_U96 (.ZN( u0_out1_3 ) , .A3( u0_u1_u4_n166 ) , .A1( u0_u1_u4_n167 ) , .A2( u0_u1_u4_n186 ) );
  NAND3_X1 u0_u1_u4_U97 (.A3( u0_u1_u4_n146 ) , .A2( u0_u1_u4_n147 ) , .A1( u0_u1_u4_n148 ) , .ZN( u0_u1_u4_n149 ) );
  NAND3_X1 u0_u1_u4_U98 (.A3( u0_u1_u4_n143 ) , .A2( u0_u1_u4_n144 ) , .A1( u0_u1_u4_n145 ) , .ZN( u0_u1_u4_n151 ) );
  NAND3_X1 u0_u1_u4_U99 (.A3( u0_u1_u4_n121 ) , .ZN( u0_u1_u4_n122 ) , .A2( u0_u1_u4_n144 ) , .A1( u0_u1_u4_n154 ) );
  INV_X1 u0_u1_u5_U10 (.A( u0_u1_u5_n121 ) , .ZN( u0_u1_u5_n177 ) );
  NOR3_X1 u0_u1_u5_U100 (.A3( u0_u1_u5_n141 ) , .A1( u0_u1_u5_n142 ) , .ZN( u0_u1_u5_n143 ) , .A2( u0_u1_u5_n191 ) );
  NAND4_X1 u0_u1_u5_U101 (.ZN( u0_out1_4 ) , .A4( u0_u1_u5_n112 ) , .A2( u0_u1_u5_n113 ) , .A1( u0_u1_u5_n114 ) , .A3( u0_u1_u5_n195 ) );
  AOI211_X1 u0_u1_u5_U102 (.A( u0_u1_u5_n110 ) , .C1( u0_u1_u5_n111 ) , .ZN( u0_u1_u5_n112 ) , .B( u0_u1_u5_n118 ) , .C2( u0_u1_u5_n177 ) );
  AOI222_X1 u0_u1_u5_U103 (.ZN( u0_u1_u5_n113 ) , .A1( u0_u1_u5_n131 ) , .C1( u0_u1_u5_n148 ) , .B2( u0_u1_u5_n174 ) , .C2( u0_u1_u5_n178 ) , .A2( u0_u1_u5_n179 ) , .B1( u0_u1_u5_n99 ) );
  NAND3_X1 u0_u1_u5_U104 (.A2( u0_u1_u5_n154 ) , .A3( u0_u1_u5_n158 ) , .A1( u0_u1_u5_n161 ) , .ZN( u0_u1_u5_n99 ) );
  NOR2_X1 u0_u1_u5_U11 (.ZN( u0_u1_u5_n160 ) , .A2( u0_u1_u5_n173 ) , .A1( u0_u1_u5_n177 ) );
  INV_X1 u0_u1_u5_U12 (.A( u0_u1_u5_n150 ) , .ZN( u0_u1_u5_n174 ) );
  AOI21_X1 u0_u1_u5_U13 (.A( u0_u1_u5_n160 ) , .B2( u0_u1_u5_n161 ) , .ZN( u0_u1_u5_n162 ) , .B1( u0_u1_u5_n192 ) );
  INV_X1 u0_u1_u5_U14 (.A( u0_u1_u5_n159 ) , .ZN( u0_u1_u5_n192 ) );
  AOI21_X1 u0_u1_u5_U15 (.A( u0_u1_u5_n156 ) , .B2( u0_u1_u5_n157 ) , .B1( u0_u1_u5_n158 ) , .ZN( u0_u1_u5_n163 ) );
  AOI21_X1 u0_u1_u5_U16 (.B2( u0_u1_u5_n139 ) , .B1( u0_u1_u5_n140 ) , .ZN( u0_u1_u5_n141 ) , .A( u0_u1_u5_n150 ) );
  OAI21_X1 u0_u1_u5_U17 (.A( u0_u1_u5_n133 ) , .B2( u0_u1_u5_n134 ) , .B1( u0_u1_u5_n135 ) , .ZN( u0_u1_u5_n142 ) );
  OAI21_X1 u0_u1_u5_U18 (.ZN( u0_u1_u5_n133 ) , .B2( u0_u1_u5_n147 ) , .A( u0_u1_u5_n173 ) , .B1( u0_u1_u5_n188 ) );
  NAND2_X1 u0_u1_u5_U19 (.A2( u0_u1_u5_n119 ) , .A1( u0_u1_u5_n123 ) , .ZN( u0_u1_u5_n137 ) );
  INV_X1 u0_u1_u5_U20 (.A( u0_u1_u5_n155 ) , .ZN( u0_u1_u5_n194 ) );
  NAND2_X1 u0_u1_u5_U21 (.A1( u0_u1_u5_n121 ) , .ZN( u0_u1_u5_n132 ) , .A2( u0_u1_u5_n172 ) );
  NAND2_X1 u0_u1_u5_U22 (.A2( u0_u1_u5_n122 ) , .ZN( u0_u1_u5_n136 ) , .A1( u0_u1_u5_n154 ) );
  NAND2_X1 u0_u1_u5_U23 (.A2( u0_u1_u5_n119 ) , .A1( u0_u1_u5_n120 ) , .ZN( u0_u1_u5_n159 ) );
  INV_X1 u0_u1_u5_U24 (.A( u0_u1_u5_n156 ) , .ZN( u0_u1_u5_n175 ) );
  INV_X1 u0_u1_u5_U25 (.A( u0_u1_u5_n158 ) , .ZN( u0_u1_u5_n188 ) );
  INV_X1 u0_u1_u5_U26 (.A( u0_u1_u5_n152 ) , .ZN( u0_u1_u5_n179 ) );
  INV_X1 u0_u1_u5_U27 (.A( u0_u1_u5_n140 ) , .ZN( u0_u1_u5_n182 ) );
  INV_X1 u0_u1_u5_U28 (.A( u0_u1_u5_n151 ) , .ZN( u0_u1_u5_n183 ) );
  INV_X1 u0_u1_u5_U29 (.A( u0_u1_u5_n123 ) , .ZN( u0_u1_u5_n185 ) );
  NOR2_X1 u0_u1_u5_U3 (.ZN( u0_u1_u5_n134 ) , .A1( u0_u1_u5_n183 ) , .A2( u0_u1_u5_n190 ) );
  INV_X1 u0_u1_u5_U30 (.A( u0_u1_u5_n161 ) , .ZN( u0_u1_u5_n184 ) );
  INV_X1 u0_u1_u5_U31 (.A( u0_u1_u5_n139 ) , .ZN( u0_u1_u5_n189 ) );
  INV_X1 u0_u1_u5_U32 (.A( u0_u1_u5_n157 ) , .ZN( u0_u1_u5_n190 ) );
  INV_X1 u0_u1_u5_U33 (.A( u0_u1_u5_n120 ) , .ZN( u0_u1_u5_n193 ) );
  NAND2_X1 u0_u1_u5_U34 (.ZN( u0_u1_u5_n111 ) , .A1( u0_u1_u5_n140 ) , .A2( u0_u1_u5_n155 ) );
  INV_X1 u0_u1_u5_U35 (.A( u0_u1_u5_n117 ) , .ZN( u0_u1_u5_n196 ) );
  OAI221_X1 u0_u1_u5_U36 (.A( u0_u1_u5_n116 ) , .ZN( u0_u1_u5_n117 ) , .B2( u0_u1_u5_n119 ) , .C1( u0_u1_u5_n153 ) , .C2( u0_u1_u5_n158 ) , .B1( u0_u1_u5_n172 ) );
  AOI222_X1 u0_u1_u5_U37 (.ZN( u0_u1_u5_n116 ) , .B2( u0_u1_u5_n145 ) , .C1( u0_u1_u5_n148 ) , .A2( u0_u1_u5_n174 ) , .C2( u0_u1_u5_n177 ) , .B1( u0_u1_u5_n187 ) , .A1( u0_u1_u5_n193 ) );
  INV_X1 u0_u1_u5_U38 (.A( u0_u1_u5_n115 ) , .ZN( u0_u1_u5_n187 ) );
  NOR2_X1 u0_u1_u5_U39 (.ZN( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n170 ) , .A2( u0_u1_u5_n180 ) );
  INV_X1 u0_u1_u5_U4 (.A( u0_u1_u5_n138 ) , .ZN( u0_u1_u5_n191 ) );
  AOI22_X1 u0_u1_u5_U40 (.B2( u0_u1_u5_n131 ) , .A2( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n169 ) , .B1( u0_u1_u5_n174 ) , .A1( u0_u1_u5_n185 ) );
  NOR2_X1 u0_u1_u5_U41 (.A1( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n150 ) , .A2( u0_u1_u5_n173 ) );
  AOI21_X1 u0_u1_u5_U42 (.A( u0_u1_u5_n118 ) , .B2( u0_u1_u5_n145 ) , .ZN( u0_u1_u5_n168 ) , .B1( u0_u1_u5_n186 ) );
  INV_X1 u0_u1_u5_U43 (.A( u0_u1_u5_n122 ) , .ZN( u0_u1_u5_n186 ) );
  NOR2_X1 u0_u1_u5_U44 (.A1( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n152 ) , .A2( u0_u1_u5_n176 ) );
  NOR2_X1 u0_u1_u5_U45 (.A1( u0_u1_u5_n115 ) , .ZN( u0_u1_u5_n118 ) , .A2( u0_u1_u5_n153 ) );
  NOR2_X1 u0_u1_u5_U46 (.A2( u0_u1_u5_n145 ) , .ZN( u0_u1_u5_n156 ) , .A1( u0_u1_u5_n174 ) );
  NOR2_X1 u0_u1_u5_U47 (.ZN( u0_u1_u5_n121 ) , .A2( u0_u1_u5_n145 ) , .A1( u0_u1_u5_n176 ) );
  AOI22_X1 u0_u1_u5_U48 (.ZN( u0_u1_u5_n114 ) , .A2( u0_u1_u5_n137 ) , .A1( u0_u1_u5_n145 ) , .B2( u0_u1_u5_n175 ) , .B1( u0_u1_u5_n193 ) );
  OAI211_X1 u0_u1_u5_U49 (.B( u0_u1_u5_n124 ) , .A( u0_u1_u5_n125 ) , .C2( u0_u1_u5_n126 ) , .C1( u0_u1_u5_n127 ) , .ZN( u0_u1_u5_n128 ) );
  OAI21_X1 u0_u1_u5_U5 (.B2( u0_u1_u5_n136 ) , .B1( u0_u1_u5_n137 ) , .ZN( u0_u1_u5_n138 ) , .A( u0_u1_u5_n177 ) );
  OAI21_X1 u0_u1_u5_U50 (.ZN( u0_u1_u5_n124 ) , .A( u0_u1_u5_n177 ) , .B2( u0_u1_u5_n183 ) , .B1( u0_u1_u5_n189 ) );
  NOR3_X1 u0_u1_u5_U51 (.ZN( u0_u1_u5_n127 ) , .A1( u0_u1_u5_n136 ) , .A3( u0_u1_u5_n148 ) , .A2( u0_u1_u5_n182 ) );
  OAI21_X1 u0_u1_u5_U52 (.ZN( u0_u1_u5_n125 ) , .A( u0_u1_u5_n174 ) , .B2( u0_u1_u5_n185 ) , .B1( u0_u1_u5_n190 ) );
  AOI21_X1 u0_u1_u5_U53 (.A( u0_u1_u5_n153 ) , .B2( u0_u1_u5_n154 ) , .B1( u0_u1_u5_n155 ) , .ZN( u0_u1_u5_n164 ) );
  AOI21_X1 u0_u1_u5_U54 (.ZN( u0_u1_u5_n110 ) , .B1( u0_u1_u5_n122 ) , .B2( u0_u1_u5_n139 ) , .A( u0_u1_u5_n153 ) );
  INV_X1 u0_u1_u5_U55 (.A( u0_u1_u5_n153 ) , .ZN( u0_u1_u5_n176 ) );
  INV_X1 u0_u1_u5_U56 (.A( u0_u1_u5_n126 ) , .ZN( u0_u1_u5_n173 ) );
  AND2_X1 u0_u1_u5_U57 (.A2( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n107 ) , .ZN( u0_u1_u5_n147 ) );
  AND2_X1 u0_u1_u5_U58 (.A2( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n108 ) , .ZN( u0_u1_u5_n148 ) );
  NAND2_X1 u0_u1_u5_U59 (.A1( u0_u1_u5_n105 ) , .A2( u0_u1_u5_n106 ) , .ZN( u0_u1_u5_n158 ) );
  INV_X1 u0_u1_u5_U6 (.A( u0_u1_u5_n135 ) , .ZN( u0_u1_u5_n178 ) );
  NAND2_X1 u0_u1_u5_U60 (.A2( u0_u1_u5_n108 ) , .A1( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n139 ) );
  NAND2_X1 u0_u1_u5_U61 (.A1( u0_u1_u5_n106 ) , .A2( u0_u1_u5_n108 ) , .ZN( u0_u1_u5_n119 ) );
  NAND2_X1 u0_u1_u5_U62 (.A2( u0_u1_u5_n103 ) , .A1( u0_u1_u5_n105 ) , .ZN( u0_u1_u5_n140 ) );
  NAND2_X1 u0_u1_u5_U63 (.A2( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n105 ) , .ZN( u0_u1_u5_n155 ) );
  NAND2_X1 u0_u1_u5_U64 (.A2( u0_u1_u5_n106 ) , .A1( u0_u1_u5_n107 ) , .ZN( u0_u1_u5_n122 ) );
  NAND2_X1 u0_u1_u5_U65 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n106 ) , .ZN( u0_u1_u5_n115 ) );
  NAND2_X1 u0_u1_u5_U66 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n103 ) , .ZN( u0_u1_u5_n161 ) );
  NAND2_X1 u0_u1_u5_U67 (.A1( u0_u1_u5_n105 ) , .A2( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n154 ) );
  INV_X1 u0_u1_u5_U68 (.A( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n172 ) );
  NAND2_X1 u0_u1_u5_U69 (.A1( u0_u1_u5_n103 ) , .A2( u0_u1_u5_n108 ) , .ZN( u0_u1_u5_n123 ) );
  OAI22_X1 u0_u1_u5_U7 (.B2( u0_u1_u5_n149 ) , .B1( u0_u1_u5_n150 ) , .A2( u0_u1_u5_n151 ) , .A1( u0_u1_u5_n152 ) , .ZN( u0_u1_u5_n165 ) );
  NAND2_X1 u0_u1_u5_U70 (.A2( u0_u1_u5_n103 ) , .A1( u0_u1_u5_n107 ) , .ZN( u0_u1_u5_n151 ) );
  NAND2_X1 u0_u1_u5_U71 (.A2( u0_u1_u5_n107 ) , .A1( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n120 ) );
  NAND2_X1 u0_u1_u5_U72 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n157 ) );
  AND2_X1 u0_u1_u5_U73 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n104 ) , .ZN( u0_u1_u5_n131 ) );
  INV_X1 u0_u1_u5_U74 (.A( u0_u1_u5_n102 ) , .ZN( u0_u1_u5_n195 ) );
  OAI221_X1 u0_u1_u5_U75 (.A( u0_u1_u5_n101 ) , .ZN( u0_u1_u5_n102 ) , .C2( u0_u1_u5_n115 ) , .C1( u0_u1_u5_n126 ) , .B1( u0_u1_u5_n134 ) , .B2( u0_u1_u5_n160 ) );
  OAI21_X1 u0_u1_u5_U76 (.ZN( u0_u1_u5_n101 ) , .B1( u0_u1_u5_n137 ) , .A( u0_u1_u5_n146 ) , .B2( u0_u1_u5_n147 ) );
  NOR2_X1 u0_u1_u5_U77 (.A2( u0_u1_X_34 ) , .A1( u0_u1_X_35 ) , .ZN( u0_u1_u5_n145 ) );
  NOR2_X1 u0_u1_u5_U78 (.A2( u0_u1_X_34 ) , .ZN( u0_u1_u5_n146 ) , .A1( u0_u1_u5_n171 ) );
  NOR2_X1 u0_u1_u5_U79 (.A2( u0_u1_X_31 ) , .A1( u0_u1_X_32 ) , .ZN( u0_u1_u5_n103 ) );
  NOR3_X1 u0_u1_u5_U8 (.A2( u0_u1_u5_n147 ) , .A1( u0_u1_u5_n148 ) , .ZN( u0_u1_u5_n149 ) , .A3( u0_u1_u5_n194 ) );
  NOR2_X1 u0_u1_u5_U80 (.A2( u0_u1_X_36 ) , .ZN( u0_u1_u5_n105 ) , .A1( u0_u1_u5_n180 ) );
  NOR2_X1 u0_u1_u5_U81 (.A2( u0_u1_X_33 ) , .ZN( u0_u1_u5_n108 ) , .A1( u0_u1_u5_n170 ) );
  NOR2_X1 u0_u1_u5_U82 (.A2( u0_u1_X_33 ) , .A1( u0_u1_X_36 ) , .ZN( u0_u1_u5_n107 ) );
  NOR2_X1 u0_u1_u5_U83 (.A2( u0_u1_X_31 ) , .ZN( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n181 ) );
  NAND2_X1 u0_u1_u5_U84 (.A2( u0_u1_X_34 ) , .A1( u0_u1_X_35 ) , .ZN( u0_u1_u5_n153 ) );
  NAND2_X1 u0_u1_u5_U85 (.A1( u0_u1_X_34 ) , .ZN( u0_u1_u5_n126 ) , .A2( u0_u1_u5_n171 ) );
  AND2_X1 u0_u1_u5_U86 (.A1( u0_u1_X_31 ) , .A2( u0_u1_X_32 ) , .ZN( u0_u1_u5_n106 ) );
  AND2_X1 u0_u1_u5_U87 (.A1( u0_u1_X_31 ) , .ZN( u0_u1_u5_n109 ) , .A2( u0_u1_u5_n181 ) );
  INV_X1 u0_u1_u5_U88 (.A( u0_u1_X_33 ) , .ZN( u0_u1_u5_n180 ) );
  INV_X1 u0_u1_u5_U89 (.A( u0_u1_X_35 ) , .ZN( u0_u1_u5_n171 ) );
  NOR2_X1 u0_u1_u5_U9 (.ZN( u0_u1_u5_n135 ) , .A1( u0_u1_u5_n173 ) , .A2( u0_u1_u5_n176 ) );
  INV_X1 u0_u1_u5_U90 (.A( u0_u1_X_36 ) , .ZN( u0_u1_u5_n170 ) );
  INV_X1 u0_u1_u5_U91 (.A( u0_u1_X_32 ) , .ZN( u0_u1_u5_n181 ) );
  NAND4_X1 u0_u1_u5_U92 (.ZN( u0_out1_29 ) , .A4( u0_u1_u5_n129 ) , .A3( u0_u1_u5_n130 ) , .A2( u0_u1_u5_n168 ) , .A1( u0_u1_u5_n196 ) );
  AOI221_X1 u0_u1_u5_U93 (.A( u0_u1_u5_n128 ) , .ZN( u0_u1_u5_n129 ) , .C2( u0_u1_u5_n132 ) , .B2( u0_u1_u5_n159 ) , .B1( u0_u1_u5_n176 ) , .C1( u0_u1_u5_n184 ) );
  AOI222_X1 u0_u1_u5_U94 (.ZN( u0_u1_u5_n130 ) , .A2( u0_u1_u5_n146 ) , .B1( u0_u1_u5_n147 ) , .C2( u0_u1_u5_n175 ) , .B2( u0_u1_u5_n179 ) , .A1( u0_u1_u5_n188 ) , .C1( u0_u1_u5_n194 ) );
  NAND4_X1 u0_u1_u5_U95 (.ZN( u0_out1_19 ) , .A4( u0_u1_u5_n166 ) , .A3( u0_u1_u5_n167 ) , .A2( u0_u1_u5_n168 ) , .A1( u0_u1_u5_n169 ) );
  AOI22_X1 u0_u1_u5_U96 (.B2( u0_u1_u5_n145 ) , .A2( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n167 ) , .B1( u0_u1_u5_n182 ) , .A1( u0_u1_u5_n189 ) );
  NOR4_X1 u0_u1_u5_U97 (.A4( u0_u1_u5_n162 ) , .A3( u0_u1_u5_n163 ) , .A2( u0_u1_u5_n164 ) , .A1( u0_u1_u5_n165 ) , .ZN( u0_u1_u5_n166 ) );
  NAND4_X1 u0_u1_u5_U98 (.ZN( u0_out1_11 ) , .A4( u0_u1_u5_n143 ) , .A3( u0_u1_u5_n144 ) , .A2( u0_u1_u5_n169 ) , .A1( u0_u1_u5_n196 ) );
  AOI22_X1 u0_u1_u5_U99 (.A2( u0_u1_u5_n132 ) , .ZN( u0_u1_u5_n144 ) , .B2( u0_u1_u5_n145 ) , .B1( u0_u1_u5_n184 ) , .A1( u0_u1_u5_n194 ) );
  AOI22_X1 u0_u1_u6_U10 (.A2( u0_u1_u6_n151 ) , .B2( u0_u1_u6_n161 ) , .A1( u0_u1_u6_n167 ) , .B1( u0_u1_u6_n170 ) , .ZN( u0_u1_u6_n89 ) );
  AOI21_X1 u0_u1_u6_U11 (.B1( u0_u1_u6_n107 ) , .B2( u0_u1_u6_n132 ) , .A( u0_u1_u6_n158 ) , .ZN( u0_u1_u6_n88 ) );
  AOI21_X1 u0_u1_u6_U12 (.B2( u0_u1_u6_n147 ) , .B1( u0_u1_u6_n148 ) , .ZN( u0_u1_u6_n149 ) , .A( u0_u1_u6_n158 ) );
  AOI21_X1 u0_u1_u6_U13 (.ZN( u0_u1_u6_n106 ) , .A( u0_u1_u6_n142 ) , .B2( u0_u1_u6_n159 ) , .B1( u0_u1_u6_n164 ) );
  INV_X1 u0_u1_u6_U14 (.A( u0_u1_u6_n155 ) , .ZN( u0_u1_u6_n161 ) );
  INV_X1 u0_u1_u6_U15 (.A( u0_u1_u6_n128 ) , .ZN( u0_u1_u6_n164 ) );
  NAND2_X1 u0_u1_u6_U16 (.ZN( u0_u1_u6_n110 ) , .A1( u0_u1_u6_n122 ) , .A2( u0_u1_u6_n129 ) );
  NAND2_X1 u0_u1_u6_U17 (.ZN( u0_u1_u6_n124 ) , .A2( u0_u1_u6_n146 ) , .A1( u0_u1_u6_n148 ) );
  INV_X1 u0_u1_u6_U18 (.A( u0_u1_u6_n132 ) , .ZN( u0_u1_u6_n171 ) );
  AND2_X1 u0_u1_u6_U19 (.A1( u0_u1_u6_n100 ) , .ZN( u0_u1_u6_n130 ) , .A2( u0_u1_u6_n147 ) );
  INV_X1 u0_u1_u6_U20 (.A( u0_u1_u6_n127 ) , .ZN( u0_u1_u6_n173 ) );
  INV_X1 u0_u1_u6_U21 (.A( u0_u1_u6_n121 ) , .ZN( u0_u1_u6_n167 ) );
  INV_X1 u0_u1_u6_U22 (.A( u0_u1_u6_n100 ) , .ZN( u0_u1_u6_n169 ) );
  INV_X1 u0_u1_u6_U23 (.A( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n170 ) );
  INV_X1 u0_u1_u6_U24 (.A( u0_u1_u6_n113 ) , .ZN( u0_u1_u6_n168 ) );
  AND2_X1 u0_u1_u6_U25 (.A1( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n119 ) , .ZN( u0_u1_u6_n133 ) );
  AND2_X1 u0_u1_u6_U26 (.A2( u0_u1_u6_n121 ) , .A1( u0_u1_u6_n122 ) , .ZN( u0_u1_u6_n131 ) );
  AND3_X1 u0_u1_u6_U27 (.ZN( u0_u1_u6_n120 ) , .A2( u0_u1_u6_n127 ) , .A1( u0_u1_u6_n132 ) , .A3( u0_u1_u6_n145 ) );
  INV_X1 u0_u1_u6_U28 (.A( u0_u1_u6_n146 ) , .ZN( u0_u1_u6_n163 ) );
  AOI222_X1 u0_u1_u6_U29 (.ZN( u0_u1_u6_n114 ) , .A1( u0_u1_u6_n118 ) , .A2( u0_u1_u6_n126 ) , .B2( u0_u1_u6_n151 ) , .C2( u0_u1_u6_n159 ) , .C1( u0_u1_u6_n168 ) , .B1( u0_u1_u6_n169 ) );
  INV_X1 u0_u1_u6_U3 (.A( u0_u1_u6_n110 ) , .ZN( u0_u1_u6_n166 ) );
  NOR2_X1 u0_u1_u6_U30 (.A1( u0_u1_u6_n162 ) , .A2( u0_u1_u6_n165 ) , .ZN( u0_u1_u6_n98 ) );
  AOI211_X1 u0_u1_u6_U31 (.B( u0_u1_u6_n134 ) , .A( u0_u1_u6_n135 ) , .C1( u0_u1_u6_n136 ) , .ZN( u0_u1_u6_n137 ) , .C2( u0_u1_u6_n151 ) );
  AOI21_X1 u0_u1_u6_U32 (.B1( u0_u1_u6_n131 ) , .ZN( u0_u1_u6_n135 ) , .A( u0_u1_u6_n144 ) , .B2( u0_u1_u6_n146 ) );
  NAND4_X1 u0_u1_u6_U33 (.A4( u0_u1_u6_n127 ) , .A3( u0_u1_u6_n128 ) , .A2( u0_u1_u6_n129 ) , .A1( u0_u1_u6_n130 ) , .ZN( u0_u1_u6_n136 ) );
  AOI21_X1 u0_u1_u6_U34 (.B2( u0_u1_u6_n132 ) , .B1( u0_u1_u6_n133 ) , .ZN( u0_u1_u6_n134 ) , .A( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U35 (.A1( u0_u1_u6_n144 ) , .ZN( u0_u1_u6_n151 ) , .A2( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U36 (.ZN( u0_u1_u6_n132 ) , .A1( u0_u1_u6_n91 ) , .A2( u0_u1_u6_n97 ) );
  AOI22_X1 u0_u1_u6_U37 (.B2( u0_u1_u6_n110 ) , .B1( u0_u1_u6_n111 ) , .A1( u0_u1_u6_n112 ) , .ZN( u0_u1_u6_n115 ) , .A2( u0_u1_u6_n161 ) );
  NAND4_X1 u0_u1_u6_U38 (.A3( u0_u1_u6_n109 ) , .ZN( u0_u1_u6_n112 ) , .A4( u0_u1_u6_n132 ) , .A2( u0_u1_u6_n147 ) , .A1( u0_u1_u6_n166 ) );
  NOR2_X1 u0_u1_u6_U39 (.ZN( u0_u1_u6_n109 ) , .A1( u0_u1_u6_n170 ) , .A2( u0_u1_u6_n173 ) );
  INV_X1 u0_u1_u6_U4 (.A( u0_u1_u6_n142 ) , .ZN( u0_u1_u6_n174 ) );
  NOR2_X1 u0_u1_u6_U40 (.A2( u0_u1_u6_n126 ) , .ZN( u0_u1_u6_n155 ) , .A1( u0_u1_u6_n160 ) );
  NAND2_X1 u0_u1_u6_U41 (.ZN( u0_u1_u6_n146 ) , .A2( u0_u1_u6_n94 ) , .A1( u0_u1_u6_n99 ) );
  AOI21_X1 u0_u1_u6_U42 (.A( u0_u1_u6_n144 ) , .B2( u0_u1_u6_n145 ) , .B1( u0_u1_u6_n146 ) , .ZN( u0_u1_u6_n150 ) );
  INV_X1 u0_u1_u6_U43 (.A( u0_u1_u6_n111 ) , .ZN( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U44 (.ZN( u0_u1_u6_n127 ) , .A1( u0_u1_u6_n91 ) , .A2( u0_u1_u6_n92 ) );
  NAND2_X1 u0_u1_u6_U45 (.ZN( u0_u1_u6_n129 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n96 ) );
  INV_X1 u0_u1_u6_U46 (.A( u0_u1_u6_n144 ) , .ZN( u0_u1_u6_n159 ) );
  NAND2_X1 u0_u1_u6_U47 (.ZN( u0_u1_u6_n145 ) , .A2( u0_u1_u6_n97 ) , .A1( u0_u1_u6_n98 ) );
  NAND2_X1 u0_u1_u6_U48 (.ZN( u0_u1_u6_n148 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n94 ) );
  NAND2_X1 u0_u1_u6_U49 (.ZN( u0_u1_u6_n108 ) , .A2( u0_u1_u6_n139 ) , .A1( u0_u1_u6_n144 ) );
  NAND2_X1 u0_u1_u6_U5 (.A2( u0_u1_u6_n143 ) , .ZN( u0_u1_u6_n152 ) , .A1( u0_u1_u6_n166 ) );
  NAND2_X1 u0_u1_u6_U50 (.ZN( u0_u1_u6_n121 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n97 ) );
  NAND2_X1 u0_u1_u6_U51 (.ZN( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n95 ) );
  AND2_X1 u0_u1_u6_U52 (.ZN( u0_u1_u6_n118 ) , .A2( u0_u1_u6_n91 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U53 (.ZN( u0_u1_u6_n147 ) , .A2( u0_u1_u6_n98 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U54 (.ZN( u0_u1_u6_n128 ) , .A1( u0_u1_u6_n94 ) , .A2( u0_u1_u6_n96 ) );
  NAND2_X1 u0_u1_u6_U55 (.ZN( u0_u1_u6_n119 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U56 (.ZN( u0_u1_u6_n123 ) , .A2( u0_u1_u6_n91 ) , .A1( u0_u1_u6_n96 ) );
  NAND2_X1 u0_u1_u6_U57 (.ZN( u0_u1_u6_n100 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n98 ) );
  NAND2_X1 u0_u1_u6_U58 (.ZN( u0_u1_u6_n122 ) , .A1( u0_u1_u6_n94 ) , .A2( u0_u1_u6_n97 ) );
  INV_X1 u0_u1_u6_U59 (.A( u0_u1_u6_n139 ) , .ZN( u0_u1_u6_n160 ) );
  AOI22_X1 u0_u1_u6_U6 (.B2( u0_u1_u6_n101 ) , .A1( u0_u1_u6_n102 ) , .ZN( u0_u1_u6_n103 ) , .B1( u0_u1_u6_n160 ) , .A2( u0_u1_u6_n161 ) );
  NAND2_X1 u0_u1_u6_U60 (.ZN( u0_u1_u6_n113 ) , .A1( u0_u1_u6_n96 ) , .A2( u0_u1_u6_n98 ) );
  NOR2_X1 u0_u1_u6_U61 (.A2( u0_u1_X_40 ) , .A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n126 ) );
  NOR2_X1 u0_u1_u6_U62 (.A2( u0_u1_X_39 ) , .A1( u0_u1_X_42 ) , .ZN( u0_u1_u6_n92 ) );
  NOR2_X1 u0_u1_u6_U63 (.A2( u0_u1_X_39 ) , .A1( u0_u1_u6_n156 ) , .ZN( u0_u1_u6_n97 ) );
  NOR2_X1 u0_u1_u6_U64 (.A2( u0_u1_X_38 ) , .A1( u0_u1_u6_n165 ) , .ZN( u0_u1_u6_n95 ) );
  NOR2_X1 u0_u1_u6_U65 (.A2( u0_u1_X_41 ) , .ZN( u0_u1_u6_n111 ) , .A1( u0_u1_u6_n157 ) );
  NOR2_X1 u0_u1_u6_U66 (.A2( u0_u1_X_37 ) , .A1( u0_u1_u6_n162 ) , .ZN( u0_u1_u6_n94 ) );
  NOR2_X1 u0_u1_u6_U67 (.A2( u0_u1_X_37 ) , .A1( u0_u1_X_38 ) , .ZN( u0_u1_u6_n91 ) );
  NAND2_X1 u0_u1_u6_U68 (.A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n144 ) , .A2( u0_u1_u6_n157 ) );
  NAND2_X1 u0_u1_u6_U69 (.A2( u0_u1_X_40 ) , .A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n139 ) );
  NOR2_X1 u0_u1_u6_U7 (.A1( u0_u1_u6_n118 ) , .ZN( u0_u1_u6_n143 ) , .A2( u0_u1_u6_n168 ) );
  AND2_X1 u0_u1_u6_U70 (.A1( u0_u1_X_39 ) , .A2( u0_u1_u6_n156 ) , .ZN( u0_u1_u6_n96 ) );
  AND2_X1 u0_u1_u6_U71 (.A1( u0_u1_X_39 ) , .A2( u0_u1_X_42 ) , .ZN( u0_u1_u6_n99 ) );
  INV_X1 u0_u1_u6_U72 (.A( u0_u1_X_40 ) , .ZN( u0_u1_u6_n157 ) );
  INV_X1 u0_u1_u6_U73 (.A( u0_u1_X_37 ) , .ZN( u0_u1_u6_n165 ) );
  INV_X1 u0_u1_u6_U74 (.A( u0_u1_X_38 ) , .ZN( u0_u1_u6_n162 ) );
  INV_X1 u0_u1_u6_U75 (.A( u0_u1_X_42 ) , .ZN( u0_u1_u6_n156 ) );
  NAND4_X1 u0_u1_u6_U76 (.ZN( u0_out1_12 ) , .A4( u0_u1_u6_n114 ) , .A3( u0_u1_u6_n115 ) , .A2( u0_u1_u6_n116 ) , .A1( u0_u1_u6_n117 ) );
  OAI22_X1 u0_u1_u6_U77 (.B2( u0_u1_u6_n111 ) , .ZN( u0_u1_u6_n116 ) , .B1( u0_u1_u6_n126 ) , .A2( u0_u1_u6_n164 ) , .A1( u0_u1_u6_n167 ) );
  OAI21_X1 u0_u1_u6_U78 (.A( u0_u1_u6_n108 ) , .ZN( u0_u1_u6_n117 ) , .B2( u0_u1_u6_n141 ) , .B1( u0_u1_u6_n163 ) );
  NAND4_X1 u0_u1_u6_U79 (.ZN( u0_out1_32 ) , .A4( u0_u1_u6_n103 ) , .A3( u0_u1_u6_n104 ) , .A2( u0_u1_u6_n105 ) , .A1( u0_u1_u6_n106 ) );
  OAI21_X1 u0_u1_u6_U8 (.A( u0_u1_u6_n159 ) , .B1( u0_u1_u6_n169 ) , .B2( u0_u1_u6_n173 ) , .ZN( u0_u1_u6_n90 ) );
  AOI22_X1 u0_u1_u6_U80 (.ZN( u0_u1_u6_n105 ) , .A2( u0_u1_u6_n108 ) , .A1( u0_u1_u6_n118 ) , .B2( u0_u1_u6_n126 ) , .B1( u0_u1_u6_n171 ) );
  AOI22_X1 u0_u1_u6_U81 (.ZN( u0_u1_u6_n104 ) , .A1( u0_u1_u6_n111 ) , .B1( u0_u1_u6_n124 ) , .B2( u0_u1_u6_n151 ) , .A2( u0_u1_u6_n93 ) );
  OAI211_X1 u0_u1_u6_U82 (.ZN( u0_out1_22 ) , .B( u0_u1_u6_n137 ) , .A( u0_u1_u6_n138 ) , .C2( u0_u1_u6_n139 ) , .C1( u0_u1_u6_n140 ) );
  AND4_X1 u0_u1_u6_U83 (.A3( u0_u1_u6_n119 ) , .A1( u0_u1_u6_n120 ) , .A4( u0_u1_u6_n129 ) , .ZN( u0_u1_u6_n140 ) , .A2( u0_u1_u6_n143 ) );
  AOI22_X1 u0_u1_u6_U84 (.B1( u0_u1_u6_n124 ) , .A2( u0_u1_u6_n125 ) , .A1( u0_u1_u6_n126 ) , .ZN( u0_u1_u6_n138 ) , .B2( u0_u1_u6_n161 ) );
  OAI211_X1 u0_u1_u6_U85 (.ZN( u0_out1_7 ) , .B( u0_u1_u6_n153 ) , .C2( u0_u1_u6_n154 ) , .C1( u0_u1_u6_n155 ) , .A( u0_u1_u6_n174 ) );
  NOR3_X1 u0_u1_u6_U86 (.A1( u0_u1_u6_n141 ) , .ZN( u0_u1_u6_n154 ) , .A3( u0_u1_u6_n164 ) , .A2( u0_u1_u6_n171 ) );
  AOI211_X1 u0_u1_u6_U87 (.B( u0_u1_u6_n149 ) , .A( u0_u1_u6_n150 ) , .C2( u0_u1_u6_n151 ) , .C1( u0_u1_u6_n152 ) , .ZN( u0_u1_u6_n153 ) );
  NAND3_X1 u0_u1_u6_U88 (.A2( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n125 ) , .A1( u0_u1_u6_n130 ) , .A3( u0_u1_u6_n131 ) );
  NAND3_X1 u0_u1_u6_U89 (.A3( u0_u1_u6_n133 ) , .ZN( u0_u1_u6_n141 ) , .A1( u0_u1_u6_n145 ) , .A2( u0_u1_u6_n148 ) );
  INV_X1 u0_u1_u6_U9 (.ZN( u0_u1_u6_n172 ) , .A( u0_u1_u6_n88 ) );
  NAND3_X1 u0_u1_u6_U90 (.ZN( u0_u1_u6_n101 ) , .A3( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n121 ) , .A1( u0_u1_u6_n127 ) );
  NAND3_X1 u0_u1_u6_U91 (.ZN( u0_u1_u6_n102 ) , .A3( u0_u1_u6_n130 ) , .A2( u0_u1_u6_n145 ) , .A1( u0_u1_u6_n166 ) );
  NAND3_X1 u0_u1_u6_U92 (.A3( u0_u1_u6_n113 ) , .A1( u0_u1_u6_n119 ) , .A2( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n93 ) );
  NAND3_X1 u0_u1_u6_U93 (.ZN( u0_u1_u6_n142 ) , .A2( u0_u1_u6_n172 ) , .A3( u0_u1_u6_n89 ) , .A1( u0_u1_u6_n90 ) );
  XOR2_X1 u0_u2_U2 (.B( u0_K3_8 ) , .A( u0_R1_5 ) , .Z( u0_u2_X_8 ) );
  XOR2_X1 u0_u2_U27 (.B( u0_K3_2 ) , .A( u0_R1_1 ) , .Z( u0_u2_X_2 ) );
  XOR2_X1 u0_u2_U3 (.B( u0_K3_7 ) , .A( u0_R1_4 ) , .Z( u0_u2_X_7 ) );
  XOR2_X1 u0_u2_U38 (.B( u0_K3_1 ) , .A( u0_R1_32 ) , .Z( u0_u2_X_1 ) );
  XOR2_X1 u0_u2_U4 (.B( u0_K3_6 ) , .A( u0_R1_5 ) , .Z( u0_u2_X_6 ) );
  XOR2_X1 u0_u2_U40 (.B( u0_K3_18 ) , .A( u0_R1_13 ) , .Z( u0_u2_X_18 ) );
  XOR2_X1 u0_u2_U41 (.B( u0_K3_17 ) , .A( u0_R1_12 ) , .Z( u0_u2_X_17 ) );
  XOR2_X1 u0_u2_U44 (.B( u0_K3_14 ) , .A( u0_R1_9 ) , .Z( u0_u2_X_14 ) );
  XOR2_X1 u0_u2_U45 (.B( u0_K3_13 ) , .A( u0_R1_8 ) , .Z( u0_u2_X_13 ) );
  XOR2_X1 u0_u2_U46 (.B( u0_K3_12 ) , .A( u0_R1_9 ) , .Z( u0_u2_X_12 ) );
  XOR2_X1 u0_u2_U47 (.B( u0_K3_11 ) , .A( u0_R1_8 ) , .Z( u0_u2_X_11 ) );
  XOR2_X1 u0_u2_U5 (.B( u0_K3_5 ) , .A( u0_R1_4 ) , .Z( u0_u2_X_5 ) );
  XOR2_X1 u0_u2_U6 (.B( u0_K3_4 ) , .A( u0_R1_3 ) , .Z( u0_u2_X_4 ) );
  AND3_X1 u0_u2_u0_U10 (.A2( u0_u2_u0_n112 ) , .ZN( u0_u2_u0_n127 ) , .A3( u0_u2_u0_n130 ) , .A1( u0_u2_u0_n148 ) );
  NAND2_X1 u0_u2_u0_U11 (.ZN( u0_u2_u0_n113 ) , .A1( u0_u2_u0_n139 ) , .A2( u0_u2_u0_n149 ) );
  AND2_X1 u0_u2_u0_U12 (.ZN( u0_u2_u0_n107 ) , .A1( u0_u2_u0_n130 ) , .A2( u0_u2_u0_n140 ) );
  AND2_X1 u0_u2_u0_U13 (.A2( u0_u2_u0_n129 ) , .A1( u0_u2_u0_n130 ) , .ZN( u0_u2_u0_n151 ) );
  AND2_X1 u0_u2_u0_U14 (.A1( u0_u2_u0_n108 ) , .A2( u0_u2_u0_n125 ) , .ZN( u0_u2_u0_n145 ) );
  INV_X1 u0_u2_u0_U15 (.A( u0_u2_u0_n143 ) , .ZN( u0_u2_u0_n173 ) );
  NOR2_X1 u0_u2_u0_U16 (.A2( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n147 ) , .A1( u0_u2_u0_n160 ) );
  INV_X1 u0_u2_u0_U17 (.ZN( u0_u2_u0_n172 ) , .A( u0_u2_u0_n88 ) );
  OAI222_X1 u0_u2_u0_U18 (.C1( u0_u2_u0_n108 ) , .A1( u0_u2_u0_n125 ) , .B2( u0_u2_u0_n128 ) , .B1( u0_u2_u0_n144 ) , .A2( u0_u2_u0_n158 ) , .C2( u0_u2_u0_n161 ) , .ZN( u0_u2_u0_n88 ) );
  NOR2_X1 u0_u2_u0_U19 (.A1( u0_u2_u0_n163 ) , .A2( u0_u2_u0_n164 ) , .ZN( u0_u2_u0_n95 ) );
  AOI21_X1 u0_u2_u0_U20 (.B1( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n132 ) , .A( u0_u2_u0_n165 ) , .B2( u0_u2_u0_n93 ) );
  INV_X1 u0_u2_u0_U21 (.A( u0_u2_u0_n142 ) , .ZN( u0_u2_u0_n165 ) );
  OAI221_X1 u0_u2_u0_U22 (.C1( u0_u2_u0_n121 ) , .ZN( u0_u2_u0_n122 ) , .B2( u0_u2_u0_n127 ) , .A( u0_u2_u0_n143 ) , .B1( u0_u2_u0_n144 ) , .C2( u0_u2_u0_n147 ) );
  OAI22_X1 u0_u2_u0_U23 (.B1( u0_u2_u0_n125 ) , .ZN( u0_u2_u0_n126 ) , .A1( u0_u2_u0_n138 ) , .A2( u0_u2_u0_n146 ) , .B2( u0_u2_u0_n147 ) );
  OAI22_X1 u0_u2_u0_U24 (.B1( u0_u2_u0_n131 ) , .A1( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n147 ) , .A2( u0_u2_u0_n90 ) , .ZN( u0_u2_u0_n91 ) );
  AND3_X1 u0_u2_u0_U25 (.A3( u0_u2_u0_n121 ) , .A2( u0_u2_u0_n125 ) , .A1( u0_u2_u0_n148 ) , .ZN( u0_u2_u0_n90 ) );
  INV_X1 u0_u2_u0_U26 (.A( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n161 ) );
  NOR2_X1 u0_u2_u0_U27 (.A1( u0_u2_u0_n120 ) , .ZN( u0_u2_u0_n143 ) , .A2( u0_u2_u0_n167 ) );
  OAI221_X1 u0_u2_u0_U28 (.C1( u0_u2_u0_n112 ) , .ZN( u0_u2_u0_n120 ) , .B1( u0_u2_u0_n138 ) , .B2( u0_u2_u0_n141 ) , .C2( u0_u2_u0_n147 ) , .A( u0_u2_u0_n172 ) );
  AOI211_X1 u0_u2_u0_U29 (.B( u0_u2_u0_n115 ) , .A( u0_u2_u0_n116 ) , .C2( u0_u2_u0_n117 ) , .C1( u0_u2_u0_n118 ) , .ZN( u0_u2_u0_n119 ) );
  INV_X1 u0_u2_u0_U3 (.A( u0_u2_u0_n113 ) , .ZN( u0_u2_u0_n166 ) );
  AOI22_X1 u0_u2_u0_U30 (.B2( u0_u2_u0_n109 ) , .A2( u0_u2_u0_n110 ) , .ZN( u0_u2_u0_n111 ) , .B1( u0_u2_u0_n118 ) , .A1( u0_u2_u0_n160 ) );
  INV_X1 u0_u2_u0_U31 (.A( u0_u2_u0_n118 ) , .ZN( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U32 (.ZN( u0_u2_u0_n104 ) , .B1( u0_u2_u0_n107 ) , .B2( u0_u2_u0_n141 ) , .A( u0_u2_u0_n144 ) );
  AOI21_X1 u0_u2_u0_U33 (.B1( u0_u2_u0_n127 ) , .B2( u0_u2_u0_n129 ) , .A( u0_u2_u0_n138 ) , .ZN( u0_u2_u0_n96 ) );
  AOI21_X1 u0_u2_u0_U34 (.ZN( u0_u2_u0_n116 ) , .B2( u0_u2_u0_n142 ) , .A( u0_u2_u0_n144 ) , .B1( u0_u2_u0_n166 ) );
  NAND2_X1 u0_u2_u0_U35 (.A1( u0_u2_u0_n100 ) , .A2( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n125 ) );
  NAND2_X1 u0_u2_u0_U36 (.A1( u0_u2_u0_n101 ) , .A2( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n150 ) );
  INV_X1 u0_u2_u0_U37 (.A( u0_u2_u0_n138 ) , .ZN( u0_u2_u0_n160 ) );
  NAND2_X1 u0_u2_u0_U38 (.A1( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n128 ) , .A2( u0_u2_u0_n95 ) );
  NAND2_X1 u0_u2_u0_U39 (.A1( u0_u2_u0_n100 ) , .ZN( u0_u2_u0_n129 ) , .A2( u0_u2_u0_n95 ) );
  AOI21_X1 u0_u2_u0_U4 (.B1( u0_u2_u0_n114 ) , .ZN( u0_u2_u0_n115 ) , .B2( u0_u2_u0_n129 ) , .A( u0_u2_u0_n161 ) );
  NAND2_X1 u0_u2_u0_U40 (.A2( u0_u2_u0_n100 ) , .ZN( u0_u2_u0_n131 ) , .A1( u0_u2_u0_n92 ) );
  NAND2_X1 u0_u2_u0_U41 (.A2( u0_u2_u0_n100 ) , .A1( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n139 ) );
  NAND2_X1 u0_u2_u0_U42 (.ZN( u0_u2_u0_n148 ) , .A1( u0_u2_u0_n93 ) , .A2( u0_u2_u0_n95 ) );
  NAND2_X1 u0_u2_u0_U43 (.A2( u0_u2_u0_n102 ) , .A1( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n149 ) );
  NAND2_X1 u0_u2_u0_U44 (.A2( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n114 ) , .A1( u0_u2_u0_n92 ) );
  NAND2_X1 u0_u2_u0_U45 (.A2( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n121 ) , .A1( u0_u2_u0_n93 ) );
  NAND2_X1 u0_u2_u0_U46 (.ZN( u0_u2_u0_n112 ) , .A2( u0_u2_u0_n92 ) , .A1( u0_u2_u0_n93 ) );
  OR3_X1 u0_u2_u0_U47 (.A3( u0_u2_u0_n152 ) , .A2( u0_u2_u0_n153 ) , .A1( u0_u2_u0_n154 ) , .ZN( u0_u2_u0_n155 ) );
  AOI21_X1 u0_u2_u0_U48 (.B2( u0_u2_u0_n150 ) , .B1( u0_u2_u0_n151 ) , .ZN( u0_u2_u0_n152 ) , .A( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U49 (.A( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n145 ) , .B1( u0_u2_u0_n146 ) , .ZN( u0_u2_u0_n154 ) );
  AOI21_X1 u0_u2_u0_U5 (.B2( u0_u2_u0_n131 ) , .ZN( u0_u2_u0_n134 ) , .B1( u0_u2_u0_n151 ) , .A( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U50 (.A( u0_u2_u0_n147 ) , .B2( u0_u2_u0_n148 ) , .B1( u0_u2_u0_n149 ) , .ZN( u0_u2_u0_n153 ) );
  INV_X1 u0_u2_u0_U51 (.ZN( u0_u2_u0_n171 ) , .A( u0_u2_u0_n99 ) );
  OAI211_X1 u0_u2_u0_U52 (.C2( u0_u2_u0_n140 ) , .C1( u0_u2_u0_n161 ) , .A( u0_u2_u0_n169 ) , .B( u0_u2_u0_n98 ) , .ZN( u0_u2_u0_n99 ) );
  AOI211_X1 u0_u2_u0_U53 (.C1( u0_u2_u0_n118 ) , .A( u0_u2_u0_n123 ) , .B( u0_u2_u0_n96 ) , .C2( u0_u2_u0_n97 ) , .ZN( u0_u2_u0_n98 ) );
  INV_X1 u0_u2_u0_U54 (.ZN( u0_u2_u0_n169 ) , .A( u0_u2_u0_n91 ) );
  NOR2_X1 u0_u2_u0_U55 (.A2( u0_u2_X_6 ) , .ZN( u0_u2_u0_n100 ) , .A1( u0_u2_u0_n162 ) );
  NOR2_X1 u0_u2_u0_U56 (.A2( u0_u2_X_4 ) , .A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n118 ) );
  NOR2_X1 u0_u2_u0_U57 (.A2( u0_u2_X_2 ) , .ZN( u0_u2_u0_n103 ) , .A1( u0_u2_u0_n164 ) );
  NOR2_X1 u0_u2_u0_U58 (.A2( u0_u2_X_1 ) , .A1( u0_u2_X_2 ) , .ZN( u0_u2_u0_n92 ) );
  NOR2_X1 u0_u2_u0_U59 (.A2( u0_u2_X_1 ) , .ZN( u0_u2_u0_n101 ) , .A1( u0_u2_u0_n163 ) );
  NOR2_X1 u0_u2_u0_U6 (.A1( u0_u2_u0_n108 ) , .ZN( u0_u2_u0_n123 ) , .A2( u0_u2_u0_n158 ) );
  NAND2_X1 u0_u2_u0_U60 (.A2( u0_u2_X_4 ) , .A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n144 ) );
  NOR2_X1 u0_u2_u0_U61 (.A2( u0_u2_X_5 ) , .ZN( u0_u2_u0_n136 ) , .A1( u0_u2_u0_n159 ) );
  NAND2_X1 u0_u2_u0_U62 (.A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n138 ) , .A2( u0_u2_u0_n159 ) );
  AND2_X1 u0_u2_u0_U63 (.A2( u0_u2_X_3 ) , .A1( u0_u2_X_6 ) , .ZN( u0_u2_u0_n102 ) );
  AND2_X1 u0_u2_u0_U64 (.A1( u0_u2_X_6 ) , .A2( u0_u2_u0_n162 ) , .ZN( u0_u2_u0_n93 ) );
  INV_X1 u0_u2_u0_U65 (.A( u0_u2_X_4 ) , .ZN( u0_u2_u0_n159 ) );
  INV_X1 u0_u2_u0_U66 (.A( u0_u2_X_1 ) , .ZN( u0_u2_u0_n164 ) );
  INV_X1 u0_u2_u0_U67 (.A( u0_u2_X_2 ) , .ZN( u0_u2_u0_n163 ) );
  INV_X1 u0_u2_u0_U68 (.ZN( u0_u2_u0_n174 ) , .A( u0_u2_u0_n89 ) );
  AOI211_X1 u0_u2_u0_U69 (.B( u0_u2_u0_n104 ) , .A( u0_u2_u0_n105 ) , .ZN( u0_u2_u0_n106 ) , .C2( u0_u2_u0_n113 ) , .C1( u0_u2_u0_n160 ) );
  OAI21_X1 u0_u2_u0_U7 (.B1( u0_u2_u0_n150 ) , .B2( u0_u2_u0_n158 ) , .A( u0_u2_u0_n172 ) , .ZN( u0_u2_u0_n89 ) );
  INV_X1 u0_u2_u0_U70 (.A( u0_u2_u0_n126 ) , .ZN( u0_u2_u0_n168 ) );
  AOI211_X1 u0_u2_u0_U71 (.B( u0_u2_u0_n133 ) , .A( u0_u2_u0_n134 ) , .C2( u0_u2_u0_n135 ) , .C1( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n137 ) );
  OR4_X1 u0_u2_u0_U72 (.ZN( u0_out2_31 ) , .A4( u0_u2_u0_n155 ) , .A2( u0_u2_u0_n156 ) , .A1( u0_u2_u0_n157 ) , .A3( u0_u2_u0_n173 ) );
  AOI21_X1 u0_u2_u0_U73 (.A( u0_u2_u0_n138 ) , .B2( u0_u2_u0_n139 ) , .B1( u0_u2_u0_n140 ) , .ZN( u0_u2_u0_n157 ) );
  AOI21_X1 u0_u2_u0_U74 (.B2( u0_u2_u0_n141 ) , .B1( u0_u2_u0_n142 ) , .ZN( u0_u2_u0_n156 ) , .A( u0_u2_u0_n161 ) );
  OR4_X1 u0_u2_u0_U75 (.ZN( u0_out2_17 ) , .A4( u0_u2_u0_n122 ) , .A2( u0_u2_u0_n123 ) , .A1( u0_u2_u0_n124 ) , .A3( u0_u2_u0_n170 ) );
  AOI21_X1 u0_u2_u0_U76 (.B2( u0_u2_u0_n107 ) , .ZN( u0_u2_u0_n124 ) , .B1( u0_u2_u0_n128 ) , .A( u0_u2_u0_n161 ) );
  INV_X1 u0_u2_u0_U77 (.A( u0_u2_u0_n111 ) , .ZN( u0_u2_u0_n170 ) );
  AOI21_X1 u0_u2_u0_U78 (.B1( u0_u2_u0_n132 ) , .ZN( u0_u2_u0_n133 ) , .A( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n166 ) );
  OAI22_X1 u0_u2_u0_U79 (.ZN( u0_u2_u0_n105 ) , .A2( u0_u2_u0_n132 ) , .B1( u0_u2_u0_n146 ) , .A1( u0_u2_u0_n147 ) , .B2( u0_u2_u0_n161 ) );
  AND2_X1 u0_u2_u0_U8 (.A1( u0_u2_u0_n114 ) , .A2( u0_u2_u0_n121 ) , .ZN( u0_u2_u0_n146 ) );
  NAND2_X1 u0_u2_u0_U80 (.ZN( u0_u2_u0_n110 ) , .A2( u0_u2_u0_n132 ) , .A1( u0_u2_u0_n145 ) );
  INV_X1 u0_u2_u0_U81 (.A( u0_u2_u0_n119 ) , .ZN( u0_u2_u0_n167 ) );
  NAND2_X1 u0_u2_u0_U82 (.A2( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n140 ) , .A1( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U83 (.A1( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n130 ) , .A2( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U84 (.ZN( u0_u2_u0_n108 ) , .A1( u0_u2_u0_n92 ) , .A2( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U85 (.ZN( u0_u2_u0_n142 ) , .A1( u0_u2_u0_n94 ) , .A2( u0_u2_u0_n95 ) );
  INV_X1 u0_u2_u0_U86 (.A( u0_u2_X_3 ) , .ZN( u0_u2_u0_n162 ) );
  NOR2_X1 u0_u2_u0_U87 (.A2( u0_u2_X_3 ) , .A1( u0_u2_X_6 ) , .ZN( u0_u2_u0_n94 ) );
  NAND3_X1 u0_u2_u0_U88 (.ZN( u0_out2_23 ) , .A3( u0_u2_u0_n137 ) , .A1( u0_u2_u0_n168 ) , .A2( u0_u2_u0_n171 ) );
  NAND3_X1 u0_u2_u0_U89 (.A3( u0_u2_u0_n127 ) , .A2( u0_u2_u0_n128 ) , .ZN( u0_u2_u0_n135 ) , .A1( u0_u2_u0_n150 ) );
  AND2_X1 u0_u2_u0_U9 (.A1( u0_u2_u0_n131 ) , .ZN( u0_u2_u0_n141 ) , .A2( u0_u2_u0_n150 ) );
  NAND3_X1 u0_u2_u0_U90 (.ZN( u0_u2_u0_n117 ) , .A3( u0_u2_u0_n132 ) , .A2( u0_u2_u0_n139 ) , .A1( u0_u2_u0_n148 ) );
  NAND3_X1 u0_u2_u0_U91 (.ZN( u0_u2_u0_n109 ) , .A2( u0_u2_u0_n114 ) , .A3( u0_u2_u0_n140 ) , .A1( u0_u2_u0_n149 ) );
  NAND3_X1 u0_u2_u0_U92 (.ZN( u0_out2_9 ) , .A3( u0_u2_u0_n106 ) , .A2( u0_u2_u0_n171 ) , .A1( u0_u2_u0_n174 ) );
  NAND3_X1 u0_u2_u0_U93 (.A2( u0_u2_u0_n128 ) , .A1( u0_u2_u0_n132 ) , .A3( u0_u2_u0_n146 ) , .ZN( u0_u2_u0_n97 ) );
  NOR2_X1 u0_u2_u1_U10 (.A1( u0_u2_u1_n112 ) , .A2( u0_u2_u1_n116 ) , .ZN( u0_u2_u1_n118 ) );
  NAND3_X1 u0_u2_u1_U100 (.ZN( u0_u2_u1_n113 ) , .A1( u0_u2_u1_n120 ) , .A3( u0_u2_u1_n133 ) , .A2( u0_u2_u1_n155 ) );
  OAI21_X1 u0_u2_u1_U11 (.ZN( u0_u2_u1_n101 ) , .B1( u0_u2_u1_n141 ) , .A( u0_u2_u1_n146 ) , .B2( u0_u2_u1_n183 ) );
  AOI21_X1 u0_u2_u1_U12 (.B2( u0_u2_u1_n155 ) , .B1( u0_u2_u1_n156 ) , .ZN( u0_u2_u1_n157 ) , .A( u0_u2_u1_n174 ) );
  OR4_X1 u0_u2_u1_U13 (.A4( u0_u2_u1_n106 ) , .A3( u0_u2_u1_n107 ) , .ZN( u0_u2_u1_n108 ) , .A1( u0_u2_u1_n117 ) , .A2( u0_u2_u1_n184 ) );
  AOI21_X1 u0_u2_u1_U14 (.ZN( u0_u2_u1_n106 ) , .A( u0_u2_u1_n112 ) , .B1( u0_u2_u1_n154 ) , .B2( u0_u2_u1_n156 ) );
  INV_X1 u0_u2_u1_U15 (.A( u0_u2_u1_n101 ) , .ZN( u0_u2_u1_n184 ) );
  AOI21_X1 u0_u2_u1_U16 (.ZN( u0_u2_u1_n107 ) , .B1( u0_u2_u1_n134 ) , .B2( u0_u2_u1_n149 ) , .A( u0_u2_u1_n174 ) );
  NAND2_X1 u0_u2_u1_U17 (.ZN( u0_u2_u1_n140 ) , .A2( u0_u2_u1_n150 ) , .A1( u0_u2_u1_n155 ) );
  NAND2_X1 u0_u2_u1_U18 (.A1( u0_u2_u1_n131 ) , .ZN( u0_u2_u1_n147 ) , .A2( u0_u2_u1_n153 ) );
  INV_X1 u0_u2_u1_U19 (.A( u0_u2_u1_n139 ) , .ZN( u0_u2_u1_n174 ) );
  INV_X1 u0_u2_u1_U20 (.A( u0_u2_u1_n112 ) , .ZN( u0_u2_u1_n171 ) );
  NAND2_X1 u0_u2_u1_U21 (.ZN( u0_u2_u1_n141 ) , .A1( u0_u2_u1_n153 ) , .A2( u0_u2_u1_n156 ) );
  AND2_X1 u0_u2_u1_U22 (.A1( u0_u2_u1_n123 ) , .ZN( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n161 ) );
  NAND2_X1 u0_u2_u1_U23 (.A2( u0_u2_u1_n115 ) , .A1( u0_u2_u1_n116 ) , .ZN( u0_u2_u1_n148 ) );
  NAND2_X1 u0_u2_u1_U24 (.A2( u0_u2_u1_n133 ) , .A1( u0_u2_u1_n135 ) , .ZN( u0_u2_u1_n159 ) );
  NAND2_X1 u0_u2_u1_U25 (.A2( u0_u2_u1_n115 ) , .A1( u0_u2_u1_n120 ) , .ZN( u0_u2_u1_n132 ) );
  INV_X1 u0_u2_u1_U26 (.A( u0_u2_u1_n154 ) , .ZN( u0_u2_u1_n178 ) );
  INV_X1 u0_u2_u1_U27 (.A( u0_u2_u1_n151 ) , .ZN( u0_u2_u1_n183 ) );
  AND2_X1 u0_u2_u1_U28 (.A1( u0_u2_u1_n129 ) , .A2( u0_u2_u1_n133 ) , .ZN( u0_u2_u1_n149 ) );
  INV_X1 u0_u2_u1_U29 (.A( u0_u2_u1_n131 ) , .ZN( u0_u2_u1_n180 ) );
  INV_X1 u0_u2_u1_U3 (.A( u0_u2_u1_n159 ) , .ZN( u0_u2_u1_n182 ) );
  OAI221_X1 u0_u2_u1_U30 (.A( u0_u2_u1_n119 ) , .C2( u0_u2_u1_n129 ) , .ZN( u0_u2_u1_n138 ) , .B2( u0_u2_u1_n152 ) , .C1( u0_u2_u1_n174 ) , .B1( u0_u2_u1_n187 ) );
  INV_X1 u0_u2_u1_U31 (.A( u0_u2_u1_n148 ) , .ZN( u0_u2_u1_n187 ) );
  AOI211_X1 u0_u2_u1_U32 (.B( u0_u2_u1_n117 ) , .A( u0_u2_u1_n118 ) , .ZN( u0_u2_u1_n119 ) , .C2( u0_u2_u1_n146 ) , .C1( u0_u2_u1_n159 ) );
  NOR2_X1 u0_u2_u1_U33 (.A1( u0_u2_u1_n168 ) , .A2( u0_u2_u1_n176 ) , .ZN( u0_u2_u1_n98 ) );
  AOI211_X1 u0_u2_u1_U34 (.B( u0_u2_u1_n162 ) , .A( u0_u2_u1_n163 ) , .C2( u0_u2_u1_n164 ) , .ZN( u0_u2_u1_n165 ) , .C1( u0_u2_u1_n171 ) );
  AOI21_X1 u0_u2_u1_U35 (.A( u0_u2_u1_n160 ) , .B2( u0_u2_u1_n161 ) , .ZN( u0_u2_u1_n162 ) , .B1( u0_u2_u1_n182 ) );
  OR2_X1 u0_u2_u1_U36 (.A2( u0_u2_u1_n157 ) , .A1( u0_u2_u1_n158 ) , .ZN( u0_u2_u1_n163 ) );
  OAI21_X1 u0_u2_u1_U37 (.B2( u0_u2_u1_n123 ) , .ZN( u0_u2_u1_n145 ) , .B1( u0_u2_u1_n160 ) , .A( u0_u2_u1_n185 ) );
  INV_X1 u0_u2_u1_U38 (.A( u0_u2_u1_n122 ) , .ZN( u0_u2_u1_n185 ) );
  AOI21_X1 u0_u2_u1_U39 (.B2( u0_u2_u1_n120 ) , .B1( u0_u2_u1_n121 ) , .ZN( u0_u2_u1_n122 ) , .A( u0_u2_u1_n128 ) );
  AOI221_X1 u0_u2_u1_U4 (.A( u0_u2_u1_n138 ) , .C2( u0_u2_u1_n139 ) , .C1( u0_u2_u1_n140 ) , .B2( u0_u2_u1_n141 ) , .ZN( u0_u2_u1_n142 ) , .B1( u0_u2_u1_n175 ) );
  NAND2_X1 u0_u2_u1_U40 (.A1( u0_u2_u1_n128 ) , .ZN( u0_u2_u1_n146 ) , .A2( u0_u2_u1_n160 ) );
  NAND2_X1 u0_u2_u1_U41 (.A2( u0_u2_u1_n112 ) , .ZN( u0_u2_u1_n139 ) , .A1( u0_u2_u1_n152 ) );
  NAND2_X1 u0_u2_u1_U42 (.A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n156 ) , .A2( u0_u2_u1_n99 ) );
  AOI221_X1 u0_u2_u1_U43 (.B1( u0_u2_u1_n140 ) , .ZN( u0_u2_u1_n167 ) , .B2( u0_u2_u1_n172 ) , .C2( u0_u2_u1_n175 ) , .C1( u0_u2_u1_n178 ) , .A( u0_u2_u1_n188 ) );
  INV_X1 u0_u2_u1_U44 (.ZN( u0_u2_u1_n188 ) , .A( u0_u2_u1_n97 ) );
  AOI211_X1 u0_u2_u1_U45 (.A( u0_u2_u1_n118 ) , .C1( u0_u2_u1_n132 ) , .C2( u0_u2_u1_n139 ) , .B( u0_u2_u1_n96 ) , .ZN( u0_u2_u1_n97 ) );
  AOI21_X1 u0_u2_u1_U46 (.B2( u0_u2_u1_n121 ) , .B1( u0_u2_u1_n135 ) , .A( u0_u2_u1_n152 ) , .ZN( u0_u2_u1_n96 ) );
  NOR2_X1 u0_u2_u1_U47 (.ZN( u0_u2_u1_n117 ) , .A1( u0_u2_u1_n121 ) , .A2( u0_u2_u1_n160 ) );
  AOI21_X1 u0_u2_u1_U48 (.A( u0_u2_u1_n128 ) , .B2( u0_u2_u1_n129 ) , .ZN( u0_u2_u1_n130 ) , .B1( u0_u2_u1_n150 ) );
  NAND2_X1 u0_u2_u1_U49 (.ZN( u0_u2_u1_n112 ) , .A1( u0_u2_u1_n169 ) , .A2( u0_u2_u1_n170 ) );
  AOI211_X1 u0_u2_u1_U5 (.ZN( u0_u2_u1_n124 ) , .A( u0_u2_u1_n138 ) , .C2( u0_u2_u1_n139 ) , .B( u0_u2_u1_n145 ) , .C1( u0_u2_u1_n147 ) );
  NAND2_X1 u0_u2_u1_U50 (.ZN( u0_u2_u1_n129 ) , .A2( u0_u2_u1_n95 ) , .A1( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U51 (.A1( u0_u2_u1_n102 ) , .ZN( u0_u2_u1_n154 ) , .A2( u0_u2_u1_n99 ) );
  NAND2_X1 u0_u2_u1_U52 (.A2( u0_u2_u1_n100 ) , .ZN( u0_u2_u1_n135 ) , .A1( u0_u2_u1_n99 ) );
  AOI21_X1 u0_u2_u1_U53 (.A( u0_u2_u1_n152 ) , .B2( u0_u2_u1_n153 ) , .B1( u0_u2_u1_n154 ) , .ZN( u0_u2_u1_n158 ) );
  INV_X1 u0_u2_u1_U54 (.A( u0_u2_u1_n160 ) , .ZN( u0_u2_u1_n175 ) );
  NAND2_X1 u0_u2_u1_U55 (.A1( u0_u2_u1_n100 ) , .ZN( u0_u2_u1_n116 ) , .A2( u0_u2_u1_n95 ) );
  NAND2_X1 u0_u2_u1_U56 (.A1( u0_u2_u1_n102 ) , .ZN( u0_u2_u1_n131 ) , .A2( u0_u2_u1_n95 ) );
  NAND2_X1 u0_u2_u1_U57 (.A2( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n121 ) , .A1( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U58 (.A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n153 ) , .A2( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U59 (.A2( u0_u2_u1_n104 ) , .A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n133 ) );
  AOI22_X1 u0_u2_u1_U6 (.B2( u0_u2_u1_n113 ) , .A2( u0_u2_u1_n114 ) , .ZN( u0_u2_u1_n125 ) , .A1( u0_u2_u1_n171 ) , .B1( u0_u2_u1_n173 ) );
  NAND2_X1 u0_u2_u1_U60 (.ZN( u0_u2_u1_n150 ) , .A2( u0_u2_u1_n98 ) , .A1( u0_u2_u1_n99 ) );
  NAND2_X1 u0_u2_u1_U61 (.A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n155 ) , .A2( u0_u2_u1_n95 ) );
  OAI21_X1 u0_u2_u1_U62 (.ZN( u0_u2_u1_n109 ) , .B1( u0_u2_u1_n129 ) , .B2( u0_u2_u1_n160 ) , .A( u0_u2_u1_n167 ) );
  NAND2_X1 u0_u2_u1_U63 (.A2( u0_u2_u1_n100 ) , .A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n120 ) );
  NAND2_X1 u0_u2_u1_U64 (.A1( u0_u2_u1_n102 ) , .A2( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n115 ) );
  NAND2_X1 u0_u2_u1_U65 (.A2( u0_u2_u1_n100 ) , .A1( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n151 ) );
  NAND2_X1 u0_u2_u1_U66 (.A2( u0_u2_u1_n103 ) , .A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n161 ) );
  INV_X1 u0_u2_u1_U67 (.A( u0_u2_u1_n152 ) , .ZN( u0_u2_u1_n173 ) );
  INV_X1 u0_u2_u1_U68 (.A( u0_u2_u1_n128 ) , .ZN( u0_u2_u1_n172 ) );
  NAND2_X1 u0_u2_u1_U69 (.A2( u0_u2_u1_n102 ) , .A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n123 ) );
  NAND2_X1 u0_u2_u1_U7 (.ZN( u0_u2_u1_n114 ) , .A1( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n156 ) );
  NOR2_X1 u0_u2_u1_U70 (.A2( u0_u2_X_7 ) , .A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n95 ) );
  NOR2_X1 u0_u2_u1_U71 (.A1( u0_u2_X_12 ) , .A2( u0_u2_X_9 ) , .ZN( u0_u2_u1_n100 ) );
  NOR2_X1 u0_u2_u1_U72 (.A2( u0_u2_X_8 ) , .A1( u0_u2_u1_n177 ) , .ZN( u0_u2_u1_n99 ) );
  NOR2_X1 u0_u2_u1_U73 (.A2( u0_u2_X_12 ) , .ZN( u0_u2_u1_n102 ) , .A1( u0_u2_u1_n176 ) );
  NOR2_X1 u0_u2_u1_U74 (.A2( u0_u2_X_9 ) , .ZN( u0_u2_u1_n105 ) , .A1( u0_u2_u1_n168 ) );
  NAND2_X1 u0_u2_u1_U75 (.A1( u0_u2_X_10 ) , .ZN( u0_u2_u1_n160 ) , .A2( u0_u2_u1_n169 ) );
  NAND2_X1 u0_u2_u1_U76 (.A2( u0_u2_X_10 ) , .A1( u0_u2_X_11 ) , .ZN( u0_u2_u1_n152 ) );
  NAND2_X1 u0_u2_u1_U77 (.A1( u0_u2_X_11 ) , .ZN( u0_u2_u1_n128 ) , .A2( u0_u2_u1_n170 ) );
  AND2_X1 u0_u2_u1_U78 (.A2( u0_u2_X_7 ) , .A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n104 ) );
  AND2_X1 u0_u2_u1_U79 (.A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n103 ) , .A2( u0_u2_u1_n177 ) );
  AOI22_X1 u0_u2_u1_U8 (.B2( u0_u2_u1_n136 ) , .A2( u0_u2_u1_n137 ) , .ZN( u0_u2_u1_n143 ) , .A1( u0_u2_u1_n171 ) , .B1( u0_u2_u1_n173 ) );
  INV_X1 u0_u2_u1_U80 (.A( u0_u2_X_10 ) , .ZN( u0_u2_u1_n170 ) );
  INV_X1 u0_u2_u1_U81 (.A( u0_u2_X_9 ) , .ZN( u0_u2_u1_n176 ) );
  INV_X1 u0_u2_u1_U82 (.A( u0_u2_X_11 ) , .ZN( u0_u2_u1_n169 ) );
  INV_X1 u0_u2_u1_U83 (.A( u0_u2_X_12 ) , .ZN( u0_u2_u1_n168 ) );
  INV_X1 u0_u2_u1_U84 (.A( u0_u2_X_7 ) , .ZN( u0_u2_u1_n177 ) );
  NAND4_X1 u0_u2_u1_U85 (.ZN( u0_out2_28 ) , .A4( u0_u2_u1_n124 ) , .A3( u0_u2_u1_n125 ) , .A2( u0_u2_u1_n126 ) , .A1( u0_u2_u1_n127 ) );
  OAI21_X1 u0_u2_u1_U86 (.ZN( u0_u2_u1_n127 ) , .B2( u0_u2_u1_n139 ) , .B1( u0_u2_u1_n175 ) , .A( u0_u2_u1_n183 ) );
  OAI21_X1 u0_u2_u1_U87 (.ZN( u0_u2_u1_n126 ) , .B2( u0_u2_u1_n140 ) , .A( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n178 ) );
  NAND4_X1 u0_u2_u1_U88 (.ZN( u0_out2_18 ) , .A4( u0_u2_u1_n165 ) , .A3( u0_u2_u1_n166 ) , .A1( u0_u2_u1_n167 ) , .A2( u0_u2_u1_n186 ) );
  AOI22_X1 u0_u2_u1_U89 (.B2( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n147 ) , .A2( u0_u2_u1_n148 ) , .ZN( u0_u2_u1_n166 ) , .A1( u0_u2_u1_n172 ) );
  INV_X1 u0_u2_u1_U9 (.A( u0_u2_u1_n147 ) , .ZN( u0_u2_u1_n181 ) );
  INV_X1 u0_u2_u1_U90 (.A( u0_u2_u1_n145 ) , .ZN( u0_u2_u1_n186 ) );
  NAND4_X1 u0_u2_u1_U91 (.ZN( u0_out2_2 ) , .A4( u0_u2_u1_n142 ) , .A3( u0_u2_u1_n143 ) , .A2( u0_u2_u1_n144 ) , .A1( u0_u2_u1_n179 ) );
  OAI21_X1 u0_u2_u1_U92 (.B2( u0_u2_u1_n132 ) , .ZN( u0_u2_u1_n144 ) , .A( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n180 ) );
  INV_X1 u0_u2_u1_U93 (.A( u0_u2_u1_n130 ) , .ZN( u0_u2_u1_n179 ) );
  OR4_X1 u0_u2_u1_U94 (.ZN( u0_out2_13 ) , .A4( u0_u2_u1_n108 ) , .A3( u0_u2_u1_n109 ) , .A2( u0_u2_u1_n110 ) , .A1( u0_u2_u1_n111 ) );
  AOI21_X1 u0_u2_u1_U95 (.ZN( u0_u2_u1_n111 ) , .A( u0_u2_u1_n128 ) , .B2( u0_u2_u1_n131 ) , .B1( u0_u2_u1_n135 ) );
  AOI21_X1 u0_u2_u1_U96 (.ZN( u0_u2_u1_n110 ) , .A( u0_u2_u1_n116 ) , .B1( u0_u2_u1_n152 ) , .B2( u0_u2_u1_n160 ) );
  NAND3_X1 u0_u2_u1_U97 (.A3( u0_u2_u1_n149 ) , .A2( u0_u2_u1_n150 ) , .A1( u0_u2_u1_n151 ) , .ZN( u0_u2_u1_n164 ) );
  NAND3_X1 u0_u2_u1_U98 (.A3( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n135 ) , .ZN( u0_u2_u1_n136 ) , .A1( u0_u2_u1_n151 ) );
  NAND3_X1 u0_u2_u1_U99 (.A1( u0_u2_u1_n133 ) , .ZN( u0_u2_u1_n137 ) , .A2( u0_u2_u1_n154 ) , .A3( u0_u2_u1_n181 ) );
  OAI22_X1 u0_u2_u2_U10 (.B1( u0_u2_u2_n151 ) , .A2( u0_u2_u2_n152 ) , .A1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n160 ) , .B2( u0_u2_u2_n168 ) );
  NAND3_X1 u0_u2_u2_U100 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n98 ) );
  NOR3_X1 u0_u2_u2_U11 (.A1( u0_u2_u2_n150 ) , .ZN( u0_u2_u2_n151 ) , .A3( u0_u2_u2_n175 ) , .A2( u0_u2_u2_n188 ) );
  AOI21_X1 u0_u2_u2_U12 (.B2( u0_u2_u2_n123 ) , .ZN( u0_u2_u2_n125 ) , .A( u0_u2_u2_n171 ) , .B1( u0_u2_u2_n184 ) );
  INV_X1 u0_u2_u2_U13 (.A( u0_u2_u2_n150 ) , .ZN( u0_u2_u2_n184 ) );
  AOI21_X1 u0_u2_u2_U14 (.ZN( u0_u2_u2_n144 ) , .B2( u0_u2_u2_n155 ) , .A( u0_u2_u2_n172 ) , .B1( u0_u2_u2_n185 ) );
  AOI21_X1 u0_u2_u2_U15 (.B2( u0_u2_u2_n143 ) , .ZN( u0_u2_u2_n145 ) , .B1( u0_u2_u2_n152 ) , .A( u0_u2_u2_n171 ) );
  INV_X1 u0_u2_u2_U16 (.A( u0_u2_u2_n156 ) , .ZN( u0_u2_u2_n171 ) );
  INV_X1 u0_u2_u2_U17 (.A( u0_u2_u2_n120 ) , .ZN( u0_u2_u2_n188 ) );
  NAND2_X1 u0_u2_u2_U18 (.A2( u0_u2_u2_n122 ) , .ZN( u0_u2_u2_n150 ) , .A1( u0_u2_u2_n152 ) );
  INV_X1 u0_u2_u2_U19 (.A( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n170 ) );
  INV_X1 u0_u2_u2_U20 (.A( u0_u2_u2_n137 ) , .ZN( u0_u2_u2_n173 ) );
  NAND2_X1 u0_u2_u2_U21 (.A1( u0_u2_u2_n132 ) , .A2( u0_u2_u2_n139 ) , .ZN( u0_u2_u2_n157 ) );
  INV_X1 u0_u2_u2_U22 (.A( u0_u2_u2_n113 ) , .ZN( u0_u2_u2_n178 ) );
  INV_X1 u0_u2_u2_U23 (.A( u0_u2_u2_n139 ) , .ZN( u0_u2_u2_n175 ) );
  INV_X1 u0_u2_u2_U24 (.A( u0_u2_u2_n155 ) , .ZN( u0_u2_u2_n181 ) );
  INV_X1 u0_u2_u2_U25 (.A( u0_u2_u2_n119 ) , .ZN( u0_u2_u2_n177 ) );
  INV_X1 u0_u2_u2_U26 (.A( u0_u2_u2_n116 ) , .ZN( u0_u2_u2_n180 ) );
  INV_X1 u0_u2_u2_U27 (.A( u0_u2_u2_n131 ) , .ZN( u0_u2_u2_n179 ) );
  INV_X1 u0_u2_u2_U28 (.A( u0_u2_u2_n154 ) , .ZN( u0_u2_u2_n176 ) );
  NAND2_X1 u0_u2_u2_U29 (.A2( u0_u2_u2_n116 ) , .A1( u0_u2_u2_n117 ) , .ZN( u0_u2_u2_n118 ) );
  NOR2_X1 u0_u2_u2_U3 (.ZN( u0_u2_u2_n121 ) , .A2( u0_u2_u2_n177 ) , .A1( u0_u2_u2_n180 ) );
  INV_X1 u0_u2_u2_U30 (.A( u0_u2_u2_n132 ) , .ZN( u0_u2_u2_n182 ) );
  INV_X1 u0_u2_u2_U31 (.A( u0_u2_u2_n158 ) , .ZN( u0_u2_u2_n183 ) );
  OAI21_X1 u0_u2_u2_U32 (.A( u0_u2_u2_n156 ) , .B1( u0_u2_u2_n157 ) , .ZN( u0_u2_u2_n158 ) , .B2( u0_u2_u2_n179 ) );
  NOR2_X1 u0_u2_u2_U33 (.ZN( u0_u2_u2_n156 ) , .A1( u0_u2_u2_n166 ) , .A2( u0_u2_u2_n169 ) );
  NOR2_X1 u0_u2_u2_U34 (.A2( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n137 ) , .A1( u0_u2_u2_n140 ) );
  NOR2_X1 u0_u2_u2_U35 (.A2( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n153 ) , .A1( u0_u2_u2_n156 ) );
  AOI211_X1 u0_u2_u2_U36 (.ZN( u0_u2_u2_n130 ) , .C1( u0_u2_u2_n138 ) , .C2( u0_u2_u2_n179 ) , .B( u0_u2_u2_n96 ) , .A( u0_u2_u2_n97 ) );
  OAI22_X1 u0_u2_u2_U37 (.B1( u0_u2_u2_n133 ) , .A2( u0_u2_u2_n137 ) , .A1( u0_u2_u2_n152 ) , .B2( u0_u2_u2_n168 ) , .ZN( u0_u2_u2_n97 ) );
  OAI221_X1 u0_u2_u2_U38 (.B1( u0_u2_u2_n113 ) , .C1( u0_u2_u2_n132 ) , .A( u0_u2_u2_n149 ) , .B2( u0_u2_u2_n171 ) , .C2( u0_u2_u2_n172 ) , .ZN( u0_u2_u2_n96 ) );
  OAI221_X1 u0_u2_u2_U39 (.A( u0_u2_u2_n115 ) , .C2( u0_u2_u2_n123 ) , .B2( u0_u2_u2_n143 ) , .B1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n163 ) , .C1( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U4 (.A( u0_u2_u2_n134 ) , .ZN( u0_u2_u2_n185 ) );
  OAI21_X1 u0_u2_u2_U40 (.A( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n115 ) , .B1( u0_u2_u2_n176 ) , .B2( u0_u2_u2_n178 ) );
  OAI221_X1 u0_u2_u2_U41 (.A( u0_u2_u2_n135 ) , .B2( u0_u2_u2_n136 ) , .B1( u0_u2_u2_n137 ) , .ZN( u0_u2_u2_n162 ) , .C2( u0_u2_u2_n167 ) , .C1( u0_u2_u2_n185 ) );
  AND3_X1 u0_u2_u2_U42 (.A3( u0_u2_u2_n131 ) , .A2( u0_u2_u2_n132 ) , .A1( u0_u2_u2_n133 ) , .ZN( u0_u2_u2_n136 ) );
  AOI22_X1 u0_u2_u2_U43 (.ZN( u0_u2_u2_n135 ) , .B1( u0_u2_u2_n140 ) , .A1( u0_u2_u2_n156 ) , .B2( u0_u2_u2_n180 ) , .A2( u0_u2_u2_n188 ) );
  AOI21_X1 u0_u2_u2_U44 (.ZN( u0_u2_u2_n149 ) , .B1( u0_u2_u2_n173 ) , .B2( u0_u2_u2_n188 ) , .A( u0_u2_u2_n95 ) );
  AND3_X1 u0_u2_u2_U45 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n156 ) , .ZN( u0_u2_u2_n95 ) );
  OAI21_X1 u0_u2_u2_U46 (.A( u0_u2_u2_n141 ) , .B2( u0_u2_u2_n142 ) , .ZN( u0_u2_u2_n146 ) , .B1( u0_u2_u2_n153 ) );
  OAI21_X1 u0_u2_u2_U47 (.A( u0_u2_u2_n140 ) , .ZN( u0_u2_u2_n141 ) , .B1( u0_u2_u2_n176 ) , .B2( u0_u2_u2_n177 ) );
  NOR3_X1 u0_u2_u2_U48 (.ZN( u0_u2_u2_n142 ) , .A3( u0_u2_u2_n175 ) , .A2( u0_u2_u2_n178 ) , .A1( u0_u2_u2_n181 ) );
  OAI21_X1 u0_u2_u2_U49 (.A( u0_u2_u2_n101 ) , .B2( u0_u2_u2_n121 ) , .B1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n164 ) );
  NOR4_X1 u0_u2_u2_U5 (.A4( u0_u2_u2_n124 ) , .A3( u0_u2_u2_n125 ) , .A2( u0_u2_u2_n126 ) , .A1( u0_u2_u2_n127 ) , .ZN( u0_u2_u2_n128 ) );
  NAND2_X1 u0_u2_u2_U50 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n155 ) );
  NAND2_X1 u0_u2_u2_U51 (.A2( u0_u2_u2_n105 ) , .A1( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n143 ) );
  NAND2_X1 u0_u2_u2_U52 (.A1( u0_u2_u2_n104 ) , .A2( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n152 ) );
  NAND2_X1 u0_u2_u2_U53 (.A1( u0_u2_u2_n100 ) , .A2( u0_u2_u2_n105 ) , .ZN( u0_u2_u2_n132 ) );
  INV_X1 u0_u2_u2_U54 (.A( u0_u2_u2_n140 ) , .ZN( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U55 (.A( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n167 ) );
  INV_X1 u0_u2_u2_U56 (.ZN( u0_u2_u2_n187 ) , .A( u0_u2_u2_n99 ) );
  OAI21_X1 u0_u2_u2_U57 (.B1( u0_u2_u2_n137 ) , .B2( u0_u2_u2_n143 ) , .A( u0_u2_u2_n98 ) , .ZN( u0_u2_u2_n99 ) );
  NAND2_X1 u0_u2_u2_U58 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n113 ) );
  NAND2_X1 u0_u2_u2_U59 (.A1( u0_u2_u2_n106 ) , .A2( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n131 ) );
  AOI21_X1 u0_u2_u2_U6 (.B2( u0_u2_u2_n119 ) , .ZN( u0_u2_u2_n127 ) , .A( u0_u2_u2_n137 ) , .B1( u0_u2_u2_n155 ) );
  NAND2_X1 u0_u2_u2_U60 (.A1( u0_u2_u2_n103 ) , .A2( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n139 ) );
  NAND2_X1 u0_u2_u2_U61 (.A1( u0_u2_u2_n103 ) , .A2( u0_u2_u2_n105 ) , .ZN( u0_u2_u2_n133 ) );
  NAND2_X1 u0_u2_u2_U62 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n103 ) , .ZN( u0_u2_u2_n154 ) );
  NAND2_X1 u0_u2_u2_U63 (.A2( u0_u2_u2_n103 ) , .A1( u0_u2_u2_n104 ) , .ZN( u0_u2_u2_n119 ) );
  NAND2_X1 u0_u2_u2_U64 (.A2( u0_u2_u2_n107 ) , .A1( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n123 ) );
  NAND2_X1 u0_u2_u2_U65 (.A1( u0_u2_u2_n104 ) , .A2( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n122 ) );
  INV_X1 u0_u2_u2_U66 (.A( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n172 ) );
  NAND2_X1 u0_u2_u2_U67 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n102 ) , .ZN( u0_u2_u2_n116 ) );
  NAND2_X1 u0_u2_u2_U68 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n120 ) );
  NAND2_X1 u0_u2_u2_U69 (.A2( u0_u2_u2_n105 ) , .A1( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n117 ) );
  AOI21_X1 u0_u2_u2_U7 (.ZN( u0_u2_u2_n124 ) , .B1( u0_u2_u2_n131 ) , .B2( u0_u2_u2_n143 ) , .A( u0_u2_u2_n172 ) );
  NOR2_X1 u0_u2_u2_U70 (.A2( u0_u2_X_16 ) , .ZN( u0_u2_u2_n140 ) , .A1( u0_u2_u2_n166 ) );
  NOR2_X1 u0_u2_u2_U71 (.A2( u0_u2_X_13 ) , .A1( u0_u2_X_14 ) , .ZN( u0_u2_u2_n100 ) );
  NOR2_X1 u0_u2_u2_U72 (.A2( u0_u2_X_16 ) , .A1( u0_u2_X_17 ) , .ZN( u0_u2_u2_n138 ) );
  NOR2_X1 u0_u2_u2_U73 (.A2( u0_u2_X_15 ) , .A1( u0_u2_X_18 ) , .ZN( u0_u2_u2_n104 ) );
  NOR2_X1 u0_u2_u2_U74 (.A2( u0_u2_X_14 ) , .ZN( u0_u2_u2_n103 ) , .A1( u0_u2_u2_n174 ) );
  NOR2_X1 u0_u2_u2_U75 (.A2( u0_u2_X_15 ) , .ZN( u0_u2_u2_n102 ) , .A1( u0_u2_u2_n165 ) );
  NOR2_X1 u0_u2_u2_U76 (.A2( u0_u2_X_17 ) , .ZN( u0_u2_u2_n114 ) , .A1( u0_u2_u2_n169 ) );
  AND2_X1 u0_u2_u2_U77 (.A1( u0_u2_X_15 ) , .ZN( u0_u2_u2_n105 ) , .A2( u0_u2_u2_n165 ) );
  AND2_X1 u0_u2_u2_U78 (.A2( u0_u2_X_15 ) , .A1( u0_u2_X_18 ) , .ZN( u0_u2_u2_n107 ) );
  AND2_X1 u0_u2_u2_U79 (.A1( u0_u2_X_14 ) , .ZN( u0_u2_u2_n106 ) , .A2( u0_u2_u2_n174 ) );
  AOI21_X1 u0_u2_u2_U8 (.B2( u0_u2_u2_n120 ) , .B1( u0_u2_u2_n121 ) , .ZN( u0_u2_u2_n126 ) , .A( u0_u2_u2_n167 ) );
  AND2_X1 u0_u2_u2_U80 (.A1( u0_u2_X_13 ) , .A2( u0_u2_X_14 ) , .ZN( u0_u2_u2_n108 ) );
  INV_X1 u0_u2_u2_U81 (.A( u0_u2_X_16 ) , .ZN( u0_u2_u2_n169 ) );
  INV_X1 u0_u2_u2_U82 (.A( u0_u2_X_17 ) , .ZN( u0_u2_u2_n166 ) );
  INV_X1 u0_u2_u2_U83 (.A( u0_u2_X_13 ) , .ZN( u0_u2_u2_n174 ) );
  INV_X1 u0_u2_u2_U84 (.A( u0_u2_X_18 ) , .ZN( u0_u2_u2_n165 ) );
  NAND4_X1 u0_u2_u2_U85 (.ZN( u0_out2_24 ) , .A4( u0_u2_u2_n111 ) , .A3( u0_u2_u2_n112 ) , .A1( u0_u2_u2_n130 ) , .A2( u0_u2_u2_n187 ) );
  AOI21_X1 u0_u2_u2_U86 (.ZN( u0_u2_u2_n112 ) , .B2( u0_u2_u2_n156 ) , .A( u0_u2_u2_n164 ) , .B1( u0_u2_u2_n181 ) );
  AOI221_X1 u0_u2_u2_U87 (.A( u0_u2_u2_n109 ) , .B1( u0_u2_u2_n110 ) , .ZN( u0_u2_u2_n111 ) , .C1( u0_u2_u2_n134 ) , .C2( u0_u2_u2_n170 ) , .B2( u0_u2_u2_n173 ) );
  NAND4_X1 u0_u2_u2_U88 (.ZN( u0_out2_16 ) , .A4( u0_u2_u2_n128 ) , .A3( u0_u2_u2_n129 ) , .A1( u0_u2_u2_n130 ) , .A2( u0_u2_u2_n186 ) );
  AOI22_X1 u0_u2_u2_U89 (.A2( u0_u2_u2_n118 ) , .ZN( u0_u2_u2_n129 ) , .A1( u0_u2_u2_n140 ) , .B1( u0_u2_u2_n157 ) , .B2( u0_u2_u2_n170 ) );
  OAI22_X1 u0_u2_u2_U9 (.ZN( u0_u2_u2_n109 ) , .A2( u0_u2_u2_n113 ) , .B2( u0_u2_u2_n133 ) , .B1( u0_u2_u2_n167 ) , .A1( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U90 (.A( u0_u2_u2_n163 ) , .ZN( u0_u2_u2_n186 ) );
  NAND4_X1 u0_u2_u2_U91 (.ZN( u0_out2_30 ) , .A4( u0_u2_u2_n147 ) , .A3( u0_u2_u2_n148 ) , .A2( u0_u2_u2_n149 ) , .A1( u0_u2_u2_n187 ) );
  NOR3_X1 u0_u2_u2_U92 (.A3( u0_u2_u2_n144 ) , .A2( u0_u2_u2_n145 ) , .A1( u0_u2_u2_n146 ) , .ZN( u0_u2_u2_n147 ) );
  AOI21_X1 u0_u2_u2_U93 (.B2( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n148 ) , .A( u0_u2_u2_n162 ) , .B1( u0_u2_u2_n182 ) );
  OR4_X1 u0_u2_u2_U94 (.ZN( u0_out2_6 ) , .A4( u0_u2_u2_n161 ) , .A3( u0_u2_u2_n162 ) , .A2( u0_u2_u2_n163 ) , .A1( u0_u2_u2_n164 ) );
  OR3_X1 u0_u2_u2_U95 (.A2( u0_u2_u2_n159 ) , .A1( u0_u2_u2_n160 ) , .ZN( u0_u2_u2_n161 ) , .A3( u0_u2_u2_n183 ) );
  AOI21_X1 u0_u2_u2_U96 (.B2( u0_u2_u2_n154 ) , .B1( u0_u2_u2_n155 ) , .ZN( u0_u2_u2_n159 ) , .A( u0_u2_u2_n167 ) );
  NAND3_X1 u0_u2_u2_U97 (.A2( u0_u2_u2_n117 ) , .A1( u0_u2_u2_n122 ) , .A3( u0_u2_u2_n123 ) , .ZN( u0_u2_u2_n134 ) );
  NAND3_X1 u0_u2_u2_U98 (.ZN( u0_u2_u2_n110 ) , .A2( u0_u2_u2_n131 ) , .A3( u0_u2_u2_n139 ) , .A1( u0_u2_u2_n154 ) );
  NAND3_X1 u0_u2_u2_U99 (.A2( u0_u2_u2_n100 ) , .ZN( u0_u2_u2_n101 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n114 ) );
  XOR2_X1 u0_u5_U10 (.B( u0_K6_45 ) , .A( u0_R4_30 ) , .Z( u0_u5_X_45 ) );
  XOR2_X1 u0_u5_U11 (.B( u0_K6_44 ) , .A( u0_R4_29 ) , .Z( u0_u5_X_44 ) );
  XOR2_X1 u0_u5_U12 (.B( u0_K6_43 ) , .A( u0_R4_28 ) , .Z( u0_u5_X_43 ) );
  XOR2_X1 u0_u5_U13 (.B( u0_K6_42 ) , .A( u0_R4_29 ) , .Z( u0_u5_X_42 ) );
  XOR2_X1 u0_u5_U14 (.B( u0_K6_41 ) , .A( u0_R4_28 ) , .Z( u0_u5_X_41 ) );
  XOR2_X1 u0_u5_U15 (.B( u0_K6_40 ) , .A( u0_R4_27 ) , .Z( u0_u5_X_40 ) );
  XOR2_X1 u0_u5_U17 (.B( u0_K6_39 ) , .A( u0_R4_26 ) , .Z( u0_u5_X_39 ) );
  XOR2_X1 u0_u5_U18 (.B( u0_K6_38 ) , .A( u0_R4_25 ) , .Z( u0_u5_X_38 ) );
  XOR2_X1 u0_u5_U19 (.B( u0_K6_37 ) , .A( u0_R4_24 ) , .Z( u0_u5_X_37 ) );
  XOR2_X1 u0_u5_U2 (.B( u0_K6_8 ) , .A( u0_R4_5 ) , .Z( u0_u5_X_8 ) );
  XOR2_X1 u0_u5_U20 (.B( u0_K6_36 ) , .A( u0_R4_25 ) , .Z( u0_u5_X_36 ) );
  XOR2_X1 u0_u5_U21 (.B( u0_K6_35 ) , .A( u0_R4_24 ) , .Z( u0_u5_X_35 ) );
  XOR2_X1 u0_u5_U23 (.B( u0_K6_33 ) , .A( u0_R4_22 ) , .Z( u0_u5_X_33 ) );
  XOR2_X1 u0_u5_U24 (.B( u0_K6_32 ) , .A( u0_R4_21 ) , .Z( u0_u5_X_32 ) );
  XOR2_X1 u0_u5_U25 (.B( u0_K6_31 ) , .A( u0_R4_20 ) , .Z( u0_u5_X_31 ) );
  XOR2_X1 u0_u5_U26 (.B( u0_K6_30 ) , .A( u0_R4_21 ) , .Z( u0_u5_X_30 ) );
  XOR2_X1 u0_u5_U27 (.B( u0_K6_2 ) , .A( u0_R4_1 ) , .Z( u0_u5_X_2 ) );
  XOR2_X1 u0_u5_U28 (.B( u0_K6_29 ) , .A( u0_R4_20 ) , .Z( u0_u5_X_29 ) );
  XOR2_X1 u0_u5_U29 (.B( u0_K6_28 ) , .A( u0_R4_19 ) , .Z( u0_u5_X_28 ) );
  XOR2_X1 u0_u5_U3 (.B( u0_K6_7 ) , .A( u0_R4_4 ) , .Z( u0_u5_X_7 ) );
  XOR2_X1 u0_u5_U31 (.B( u0_K6_26 ) , .A( u0_R4_17 ) , .Z( u0_u5_X_26 ) );
  XOR2_X1 u0_u5_U32 (.B( u0_K6_25 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_25 ) );
  XOR2_X1 u0_u5_U33 (.B( u0_K6_24 ) , .A( u0_R4_17 ) , .Z( u0_u5_X_24 ) );
  XOR2_X1 u0_u5_U34 (.B( u0_K6_23 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_23 ) );
  XOR2_X1 u0_u5_U37 (.B( u0_K6_20 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_20 ) );
  XOR2_X1 u0_u5_U38 (.B( u0_K6_1 ) , .A( u0_R4_32 ) , .Z( u0_u5_X_1 ) );
  XOR2_X1 u0_u5_U39 (.B( u0_K6_19 ) , .A( u0_R4_12 ) , .Z( u0_u5_X_19 ) );
  XOR2_X1 u0_u5_U4 (.B( u0_K6_6 ) , .A( u0_R4_5 ) , .Z( u0_u5_X_6 ) );
  XOR2_X1 u0_u5_U40 (.B( u0_K6_18 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_18 ) );
  XOR2_X1 u0_u5_U41 (.B( u0_K6_17 ) , .A( u0_R4_12 ) , .Z( u0_u5_X_17 ) );
  XOR2_X1 u0_u5_U44 (.B( u0_K6_14 ) , .A( u0_R4_9 ) , .Z( u0_u5_X_14 ) );
  XOR2_X1 u0_u5_U45 (.B( u0_K6_13 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_13 ) );
  XOR2_X1 u0_u5_U46 (.B( u0_K6_12 ) , .A( u0_R4_9 ) , .Z( u0_u5_X_12 ) );
  XOR2_X1 u0_u5_U47 (.B( u0_K6_11 ) , .A( u0_R4_8 ) , .Z( u0_u5_X_11 ) );
  XOR2_X1 u0_u5_U5 (.B( u0_K6_5 ) , .A( u0_R4_4 ) , .Z( u0_u5_X_5 ) );
  XOR2_X1 u0_u5_U6 (.B( u0_K6_4 ) , .A( u0_R4_3 ) , .Z( u0_u5_X_4 ) );
  XOR2_X1 u0_u5_U7 (.B( u0_K6_48 ) , .A( u0_R4_1 ) , .Z( u0_u5_X_48 ) );
  XOR2_X1 u0_u5_U8 (.B( u0_K6_47 ) , .A( u0_R4_32 ) , .Z( u0_u5_X_47 ) );
  AND2_X1 u0_u5_u0_U10 (.A1( u0_u5_u0_n131 ) , .ZN( u0_u5_u0_n141 ) , .A2( u0_u5_u0_n150 ) );
  AND3_X1 u0_u5_u0_U11 (.A2( u0_u5_u0_n112 ) , .ZN( u0_u5_u0_n127 ) , .A3( u0_u5_u0_n130 ) , .A1( u0_u5_u0_n148 ) );
  AND2_X1 u0_u5_u0_U12 (.ZN( u0_u5_u0_n107 ) , .A1( u0_u5_u0_n130 ) , .A2( u0_u5_u0_n140 ) );
  AND2_X1 u0_u5_u0_U13 (.A2( u0_u5_u0_n129 ) , .A1( u0_u5_u0_n130 ) , .ZN( u0_u5_u0_n151 ) );
  AND2_X1 u0_u5_u0_U14 (.A1( u0_u5_u0_n108 ) , .A2( u0_u5_u0_n125 ) , .ZN( u0_u5_u0_n145 ) );
  INV_X1 u0_u5_u0_U15 (.A( u0_u5_u0_n143 ) , .ZN( u0_u5_u0_n173 ) );
  NOR2_X1 u0_u5_u0_U16 (.A2( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n147 ) , .A1( u0_u5_u0_n160 ) );
  AOI21_X1 u0_u5_u0_U17 (.B1( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n132 ) , .A( u0_u5_u0_n165 ) , .B2( u0_u5_u0_n93 ) );
  OAI22_X1 u0_u5_u0_U18 (.B1( u0_u5_u0_n131 ) , .A1( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n147 ) , .A2( u0_u5_u0_n90 ) , .ZN( u0_u5_u0_n91 ) );
  AND3_X1 u0_u5_u0_U19 (.A3( u0_u5_u0_n121 ) , .A2( u0_u5_u0_n125 ) , .A1( u0_u5_u0_n148 ) , .ZN( u0_u5_u0_n90 ) );
  OAI22_X1 u0_u5_u0_U20 (.B1( u0_u5_u0_n125 ) , .ZN( u0_u5_u0_n126 ) , .A1( u0_u5_u0_n138 ) , .A2( u0_u5_u0_n146 ) , .B2( u0_u5_u0_n147 ) );
  NOR2_X1 u0_u5_u0_U21 (.A1( u0_u5_u0_n163 ) , .A2( u0_u5_u0_n164 ) , .ZN( u0_u5_u0_n95 ) );
  AOI22_X1 u0_u5_u0_U22 (.B2( u0_u5_u0_n109 ) , .A2( u0_u5_u0_n110 ) , .ZN( u0_u5_u0_n111 ) , .B1( u0_u5_u0_n118 ) , .A1( u0_u5_u0_n160 ) );
  NAND2_X1 u0_u5_u0_U23 (.A2( u0_u5_u0_n102 ) , .A1( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n149 ) );
  INV_X1 u0_u5_u0_U24 (.A( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n161 ) );
  INV_X1 u0_u5_u0_U25 (.A( u0_u5_u0_n118 ) , .ZN( u0_u5_u0_n158 ) );
  NAND2_X1 u0_u5_u0_U26 (.A2( u0_u5_u0_n100 ) , .ZN( u0_u5_u0_n131 ) , .A1( u0_u5_u0_n92 ) );
  NAND2_X1 u0_u5_u0_U27 (.ZN( u0_u5_u0_n108 ) , .A1( u0_u5_u0_n92 ) , .A2( u0_u5_u0_n94 ) );
  AOI21_X1 u0_u5_u0_U28 (.ZN( u0_u5_u0_n104 ) , .B1( u0_u5_u0_n107 ) , .B2( u0_u5_u0_n141 ) , .A( u0_u5_u0_n144 ) );
  AOI21_X1 u0_u5_u0_U29 (.B1( u0_u5_u0_n127 ) , .B2( u0_u5_u0_n129 ) , .A( u0_u5_u0_n138 ) , .ZN( u0_u5_u0_n96 ) );
  INV_X1 u0_u5_u0_U3 (.A( u0_u5_u0_n113 ) , .ZN( u0_u5_u0_n166 ) );
  NAND2_X1 u0_u5_u0_U30 (.A2( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n114 ) , .A1( u0_u5_u0_n92 ) );
  NOR2_X1 u0_u5_u0_U31 (.A1( u0_u5_u0_n120 ) , .ZN( u0_u5_u0_n143 ) , .A2( u0_u5_u0_n167 ) );
  OAI221_X1 u0_u5_u0_U32 (.C1( u0_u5_u0_n112 ) , .ZN( u0_u5_u0_n120 ) , .B1( u0_u5_u0_n138 ) , .B2( u0_u5_u0_n141 ) , .C2( u0_u5_u0_n147 ) , .A( u0_u5_u0_n172 ) );
  AOI211_X1 u0_u5_u0_U33 (.B( u0_u5_u0_n115 ) , .A( u0_u5_u0_n116 ) , .C2( u0_u5_u0_n117 ) , .C1( u0_u5_u0_n118 ) , .ZN( u0_u5_u0_n119 ) );
  NAND2_X1 u0_u5_u0_U34 (.A2( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n140 ) , .A1( u0_u5_u0_n94 ) );
  NAND2_X1 u0_u5_u0_U35 (.A1( u0_u5_u0_n100 ) , .A2( u0_u5_u0_n103 ) , .ZN( u0_u5_u0_n125 ) );
  NAND2_X1 u0_u5_u0_U36 (.A1( u0_u5_u0_n101 ) , .A2( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n150 ) );
  INV_X1 u0_u5_u0_U37 (.A( u0_u5_u0_n138 ) , .ZN( u0_u5_u0_n160 ) );
  NAND2_X1 u0_u5_u0_U38 (.A2( u0_u5_u0_n100 ) , .A1( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n139 ) );
  NAND2_X1 u0_u5_u0_U39 (.ZN( u0_u5_u0_n112 ) , .A2( u0_u5_u0_n92 ) , .A1( u0_u5_u0_n93 ) );
  AOI21_X1 u0_u5_u0_U4 (.B1( u0_u5_u0_n114 ) , .ZN( u0_u5_u0_n115 ) , .B2( u0_u5_u0_n129 ) , .A( u0_u5_u0_n161 ) );
  NAND2_X1 u0_u5_u0_U40 (.A1( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n130 ) , .A2( u0_u5_u0_n94 ) );
  INV_X1 u0_u5_u0_U41 (.ZN( u0_u5_u0_n172 ) , .A( u0_u5_u0_n88 ) );
  OAI222_X1 u0_u5_u0_U42 (.C1( u0_u5_u0_n108 ) , .A1( u0_u5_u0_n125 ) , .B2( u0_u5_u0_n128 ) , .B1( u0_u5_u0_n144 ) , .A2( u0_u5_u0_n158 ) , .C2( u0_u5_u0_n161 ) , .ZN( u0_u5_u0_n88 ) );
  NAND2_X1 u0_u5_u0_U43 (.A2( u0_u5_u0_n101 ) , .ZN( u0_u5_u0_n121 ) , .A1( u0_u5_u0_n93 ) );
  OR3_X1 u0_u5_u0_U44 (.A3( u0_u5_u0_n152 ) , .A2( u0_u5_u0_n153 ) , .A1( u0_u5_u0_n154 ) , .ZN( u0_u5_u0_n155 ) );
  AOI21_X1 u0_u5_u0_U45 (.A( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n145 ) , .B1( u0_u5_u0_n146 ) , .ZN( u0_u5_u0_n154 ) );
  AOI21_X1 u0_u5_u0_U46 (.B2( u0_u5_u0_n150 ) , .B1( u0_u5_u0_n151 ) , .ZN( u0_u5_u0_n152 ) , .A( u0_u5_u0_n158 ) );
  AOI21_X1 u0_u5_u0_U47 (.A( u0_u5_u0_n147 ) , .B2( u0_u5_u0_n148 ) , .B1( u0_u5_u0_n149 ) , .ZN( u0_u5_u0_n153 ) );
  INV_X1 u0_u5_u0_U48 (.ZN( u0_u5_u0_n171 ) , .A( u0_u5_u0_n99 ) );
  OAI211_X1 u0_u5_u0_U49 (.C2( u0_u5_u0_n140 ) , .C1( u0_u5_u0_n161 ) , .A( u0_u5_u0_n169 ) , .B( u0_u5_u0_n98 ) , .ZN( u0_u5_u0_n99 ) );
  AOI21_X1 u0_u5_u0_U5 (.B2( u0_u5_u0_n131 ) , .ZN( u0_u5_u0_n134 ) , .B1( u0_u5_u0_n151 ) , .A( u0_u5_u0_n158 ) );
  AOI211_X1 u0_u5_u0_U50 (.C1( u0_u5_u0_n118 ) , .A( u0_u5_u0_n123 ) , .B( u0_u5_u0_n96 ) , .C2( u0_u5_u0_n97 ) , .ZN( u0_u5_u0_n98 ) );
  INV_X1 u0_u5_u0_U51 (.ZN( u0_u5_u0_n169 ) , .A( u0_u5_u0_n91 ) );
  NOR2_X1 u0_u5_u0_U52 (.A2( u0_u5_X_4 ) , .A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n118 ) );
  NOR2_X1 u0_u5_u0_U53 (.A2( u0_u5_X_1 ) , .ZN( u0_u5_u0_n101 ) , .A1( u0_u5_u0_n163 ) );
  NOR2_X1 u0_u5_u0_U54 (.A2( u0_u5_X_3 ) , .A1( u0_u5_X_6 ) , .ZN( u0_u5_u0_n94 ) );
  NOR2_X1 u0_u5_u0_U55 (.A2( u0_u5_X_6 ) , .ZN( u0_u5_u0_n100 ) , .A1( u0_u5_u0_n162 ) );
  NAND2_X1 u0_u5_u0_U56 (.A2( u0_u5_X_4 ) , .A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n144 ) );
  NOR2_X1 u0_u5_u0_U57 (.A2( u0_u5_X_5 ) , .ZN( u0_u5_u0_n136 ) , .A1( u0_u5_u0_n159 ) );
  NAND2_X1 u0_u5_u0_U58 (.A1( u0_u5_X_5 ) , .ZN( u0_u5_u0_n138 ) , .A2( u0_u5_u0_n159 ) );
  AND2_X1 u0_u5_u0_U59 (.A2( u0_u5_X_3 ) , .A1( u0_u5_X_6 ) , .ZN( u0_u5_u0_n102 ) );
  NOR2_X1 u0_u5_u0_U6 (.A1( u0_u5_u0_n108 ) , .ZN( u0_u5_u0_n123 ) , .A2( u0_u5_u0_n158 ) );
  AND2_X1 u0_u5_u0_U60 (.A1( u0_u5_X_6 ) , .A2( u0_u5_u0_n162 ) , .ZN( u0_u5_u0_n93 ) );
  INV_X1 u0_u5_u0_U61 (.A( u0_u5_X_4 ) , .ZN( u0_u5_u0_n159 ) );
  INV_X1 u0_u5_u0_U62 (.A( u0_u5_X_1 ) , .ZN( u0_u5_u0_n164 ) );
  INV_X1 u0_u5_u0_U63 (.A( u0_u5_X_3 ) , .ZN( u0_u5_u0_n162 ) );
  AOI211_X1 u0_u5_u0_U64 (.B( u0_u5_u0_n133 ) , .A( u0_u5_u0_n134 ) , .C2( u0_u5_u0_n135 ) , .C1( u0_u5_u0_n136 ) , .ZN( u0_u5_u0_n137 ) );
  INV_X1 u0_u5_u0_U65 (.A( u0_u5_u0_n126 ) , .ZN( u0_u5_u0_n168 ) );
  OR4_X1 u0_u5_u0_U66 (.ZN( u0_out5_17 ) , .A4( u0_u5_u0_n122 ) , .A2( u0_u5_u0_n123 ) , .A1( u0_u5_u0_n124 ) , .A3( u0_u5_u0_n170 ) );
  AOI21_X1 u0_u5_u0_U67 (.B2( u0_u5_u0_n107 ) , .ZN( u0_u5_u0_n124 ) , .B1( u0_u5_u0_n128 ) , .A( u0_u5_u0_n161 ) );
  INV_X1 u0_u5_u0_U68 (.A( u0_u5_u0_n111 ) , .ZN( u0_u5_u0_n170 ) );
  OR4_X1 u0_u5_u0_U69 (.ZN( u0_out5_31 ) , .A4( u0_u5_u0_n155 ) , .A2( u0_u5_u0_n156 ) , .A1( u0_u5_u0_n157 ) , .A3( u0_u5_u0_n173 ) );
  OAI21_X1 u0_u5_u0_U7 (.B1( u0_u5_u0_n150 ) , .B2( u0_u5_u0_n158 ) , .A( u0_u5_u0_n172 ) , .ZN( u0_u5_u0_n89 ) );
  AOI21_X1 u0_u5_u0_U70 (.A( u0_u5_u0_n138 ) , .B2( u0_u5_u0_n139 ) , .B1( u0_u5_u0_n140 ) , .ZN( u0_u5_u0_n157 ) );
  INV_X1 u0_u5_u0_U71 (.ZN( u0_u5_u0_n174 ) , .A( u0_u5_u0_n89 ) );
  AOI211_X1 u0_u5_u0_U72 (.B( u0_u5_u0_n104 ) , .A( u0_u5_u0_n105 ) , .ZN( u0_u5_u0_n106 ) , .C2( u0_u5_u0_n113 ) , .C1( u0_u5_u0_n160 ) );
  INV_X1 u0_u5_u0_U73 (.A( u0_u5_u0_n142 ) , .ZN( u0_u5_u0_n165 ) );
  AOI21_X1 u0_u5_u0_U74 (.ZN( u0_u5_u0_n116 ) , .B2( u0_u5_u0_n142 ) , .A( u0_u5_u0_n144 ) , .B1( u0_u5_u0_n166 ) );
  AOI21_X1 u0_u5_u0_U75 (.B2( u0_u5_u0_n141 ) , .B1( u0_u5_u0_n142 ) , .ZN( u0_u5_u0_n156 ) , .A( u0_u5_u0_n161 ) );
  OAI221_X1 u0_u5_u0_U76 (.C1( u0_u5_u0_n121 ) , .ZN( u0_u5_u0_n122 ) , .B2( u0_u5_u0_n127 ) , .A( u0_u5_u0_n143 ) , .B1( u0_u5_u0_n144 ) , .C2( u0_u5_u0_n147 ) );
  AOI21_X1 u0_u5_u0_U77 (.B1( u0_u5_u0_n132 ) , .ZN( u0_u5_u0_n133 ) , .A( u0_u5_u0_n144 ) , .B2( u0_u5_u0_n166 ) );
  OAI22_X1 u0_u5_u0_U78 (.ZN( u0_u5_u0_n105 ) , .A2( u0_u5_u0_n132 ) , .B1( u0_u5_u0_n146 ) , .A1( u0_u5_u0_n147 ) , .B2( u0_u5_u0_n161 ) );
  NAND2_X1 u0_u5_u0_U79 (.ZN( u0_u5_u0_n110 ) , .A2( u0_u5_u0_n132 ) , .A1( u0_u5_u0_n145 ) );
  AND2_X1 u0_u5_u0_U8 (.A1( u0_u5_u0_n114 ) , .A2( u0_u5_u0_n121 ) , .ZN( u0_u5_u0_n146 ) );
  INV_X1 u0_u5_u0_U80 (.A( u0_u5_u0_n119 ) , .ZN( u0_u5_u0_n167 ) );
  NAND2_X1 u0_u5_u0_U81 (.ZN( u0_u5_u0_n148 ) , .A1( u0_u5_u0_n93 ) , .A2( u0_u5_u0_n95 ) );
  NAND2_X1 u0_u5_u0_U82 (.A1( u0_u5_u0_n100 ) , .ZN( u0_u5_u0_n129 ) , .A2( u0_u5_u0_n95 ) );
  NAND2_X1 u0_u5_u0_U83 (.A1( u0_u5_u0_n102 ) , .ZN( u0_u5_u0_n128 ) , .A2( u0_u5_u0_n95 ) );
  NOR2_X1 u0_u5_u0_U84 (.A2( u0_u5_X_1 ) , .A1( u0_u5_X_2 ) , .ZN( u0_u5_u0_n92 ) );
  NAND2_X1 u0_u5_u0_U85 (.ZN( u0_u5_u0_n142 ) , .A1( u0_u5_u0_n94 ) , .A2( u0_u5_u0_n95 ) );
  NOR2_X1 u0_u5_u0_U86 (.A2( u0_u5_X_2 ) , .ZN( u0_u5_u0_n103 ) , .A1( u0_u5_u0_n164 ) );
  INV_X1 u0_u5_u0_U87 (.A( u0_u5_X_2 ) , .ZN( u0_u5_u0_n163 ) );
  NAND3_X1 u0_u5_u0_U88 (.ZN( u0_out5_23 ) , .A3( u0_u5_u0_n137 ) , .A1( u0_u5_u0_n168 ) , .A2( u0_u5_u0_n171 ) );
  NAND3_X1 u0_u5_u0_U89 (.A3( u0_u5_u0_n127 ) , .A2( u0_u5_u0_n128 ) , .ZN( u0_u5_u0_n135 ) , .A1( u0_u5_u0_n150 ) );
  NAND2_X1 u0_u5_u0_U9 (.ZN( u0_u5_u0_n113 ) , .A1( u0_u5_u0_n139 ) , .A2( u0_u5_u0_n149 ) );
  NAND3_X1 u0_u5_u0_U90 (.ZN( u0_u5_u0_n117 ) , .A3( u0_u5_u0_n132 ) , .A2( u0_u5_u0_n139 ) , .A1( u0_u5_u0_n148 ) );
  NAND3_X1 u0_u5_u0_U91 (.ZN( u0_u5_u0_n109 ) , .A2( u0_u5_u0_n114 ) , .A3( u0_u5_u0_n140 ) , .A1( u0_u5_u0_n149 ) );
  NAND3_X1 u0_u5_u0_U92 (.ZN( u0_out5_9 ) , .A3( u0_u5_u0_n106 ) , .A2( u0_u5_u0_n171 ) , .A1( u0_u5_u0_n174 ) );
  NAND3_X1 u0_u5_u0_U93 (.A2( u0_u5_u0_n128 ) , .A1( u0_u5_u0_n132 ) , .A3( u0_u5_u0_n146 ) , .ZN( u0_u5_u0_n97 ) );
  NOR2_X1 u0_u5_u1_U10 (.A1( u0_u5_u1_n112 ) , .A2( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n118 ) );
  NAND3_X1 u0_u5_u1_U100 (.ZN( u0_u5_u1_n113 ) , .A1( u0_u5_u1_n120 ) , .A3( u0_u5_u1_n133 ) , .A2( u0_u5_u1_n155 ) );
  OAI21_X1 u0_u5_u1_U11 (.ZN( u0_u5_u1_n101 ) , .B1( u0_u5_u1_n141 ) , .A( u0_u5_u1_n146 ) , .B2( u0_u5_u1_n183 ) );
  AOI21_X1 u0_u5_u1_U12 (.B2( u0_u5_u1_n155 ) , .B1( u0_u5_u1_n156 ) , .ZN( u0_u5_u1_n157 ) , .A( u0_u5_u1_n174 ) );
  NAND2_X1 u0_u5_u1_U13 (.ZN( u0_u5_u1_n140 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n155 ) );
  NAND2_X1 u0_u5_u1_U14 (.A1( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n153 ) );
  INV_X1 u0_u5_u1_U15 (.A( u0_u5_u1_n139 ) , .ZN( u0_u5_u1_n174 ) );
  OR4_X1 u0_u5_u1_U16 (.A4( u0_u5_u1_n106 ) , .A3( u0_u5_u1_n107 ) , .ZN( u0_u5_u1_n108 ) , .A1( u0_u5_u1_n117 ) , .A2( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U17 (.ZN( u0_u5_u1_n106 ) , .A( u0_u5_u1_n112 ) , .B1( u0_u5_u1_n154 ) , .B2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U18 (.A( u0_u5_u1_n101 ) , .ZN( u0_u5_u1_n184 ) );
  AOI21_X1 u0_u5_u1_U19 (.ZN( u0_u5_u1_n107 ) , .B1( u0_u5_u1_n134 ) , .B2( u0_u5_u1_n149 ) , .A( u0_u5_u1_n174 ) );
  INV_X1 u0_u5_u1_U20 (.A( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n171 ) );
  NAND2_X1 u0_u5_u1_U21 (.ZN( u0_u5_u1_n141 ) , .A1( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n156 ) );
  AND2_X1 u0_u5_u1_U22 (.A1( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n161 ) );
  NAND2_X1 u0_u5_u1_U23 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n116 ) , .ZN( u0_u5_u1_n148 ) );
  NAND2_X1 u0_u5_u1_U24 (.A2( u0_u5_u1_n133 ) , .A1( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n159 ) );
  NAND2_X1 u0_u5_u1_U25 (.A2( u0_u5_u1_n115 ) , .A1( u0_u5_u1_n120 ) , .ZN( u0_u5_u1_n132 ) );
  INV_X1 u0_u5_u1_U26 (.A( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n178 ) );
  INV_X1 u0_u5_u1_U27 (.A( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n183 ) );
  AND2_X1 u0_u5_u1_U28 (.A1( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n149 ) );
  INV_X1 u0_u5_u1_U29 (.A( u0_u5_u1_n131 ) , .ZN( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U3 (.A( u0_u5_u1_n159 ) , .ZN( u0_u5_u1_n182 ) );
  OAI221_X1 u0_u5_u1_U30 (.A( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n138 ) , .B2( u0_u5_u1_n152 ) , .C1( u0_u5_u1_n174 ) , .B1( u0_u5_u1_n187 ) );
  INV_X1 u0_u5_u1_U31 (.A( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n187 ) );
  AOI211_X1 u0_u5_u1_U32 (.B( u0_u5_u1_n117 ) , .A( u0_u5_u1_n118 ) , .ZN( u0_u5_u1_n119 ) , .C2( u0_u5_u1_n146 ) , .C1( u0_u5_u1_n159 ) );
  NOR2_X1 u0_u5_u1_U33 (.A1( u0_u5_u1_n168 ) , .A2( u0_u5_u1_n176 ) , .ZN( u0_u5_u1_n98 ) );
  OAI21_X1 u0_u5_u1_U34 (.B2( u0_u5_u1_n123 ) , .ZN( u0_u5_u1_n145 ) , .B1( u0_u5_u1_n160 ) , .A( u0_u5_u1_n185 ) );
  INV_X1 u0_u5_u1_U35 (.A( u0_u5_u1_n122 ) , .ZN( u0_u5_u1_n185 ) );
  AOI21_X1 u0_u5_u1_U36 (.B2( u0_u5_u1_n120 ) , .B1( u0_u5_u1_n121 ) , .ZN( u0_u5_u1_n122 ) , .A( u0_u5_u1_n128 ) );
  NAND2_X1 u0_u5_u1_U37 (.A1( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n146 ) , .A2( u0_u5_u1_n160 ) );
  NAND2_X1 u0_u5_u1_U38 (.A2( u0_u5_u1_n112 ) , .ZN( u0_u5_u1_n139 ) , .A1( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U39 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n156 ) , .A2( u0_u5_u1_n99 ) );
  AOI221_X1 u0_u5_u1_U4 (.A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .C1( u0_u5_u1_n140 ) , .B2( u0_u5_u1_n141 ) , .ZN( u0_u5_u1_n142 ) , .B1( u0_u5_u1_n175 ) );
  AOI221_X1 u0_u5_u1_U40 (.B1( u0_u5_u1_n140 ) , .ZN( u0_u5_u1_n167 ) , .B2( u0_u5_u1_n172 ) , .C2( u0_u5_u1_n175 ) , .C1( u0_u5_u1_n178 ) , .A( u0_u5_u1_n188 ) );
  INV_X1 u0_u5_u1_U41 (.ZN( u0_u5_u1_n188 ) , .A( u0_u5_u1_n97 ) );
  AOI211_X1 u0_u5_u1_U42 (.A( u0_u5_u1_n118 ) , .C1( u0_u5_u1_n132 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n96 ) , .ZN( u0_u5_u1_n97 ) );
  AOI21_X1 u0_u5_u1_U43 (.B2( u0_u5_u1_n121 ) , .B1( u0_u5_u1_n135 ) , .A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n96 ) );
  NOR2_X1 u0_u5_u1_U44 (.ZN( u0_u5_u1_n117 ) , .A1( u0_u5_u1_n121 ) , .A2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U45 (.A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n129 ) , .ZN( u0_u5_u1_n130 ) , .B1( u0_u5_u1_n150 ) );
  NAND2_X1 u0_u5_u1_U46 (.ZN( u0_u5_u1_n112 ) , .A1( u0_u5_u1_n169 ) , .A2( u0_u5_u1_n170 ) );
  NAND2_X1 u0_u5_u1_U47 (.ZN( u0_u5_u1_n129 ) , .A2( u0_u5_u1_n95 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U48 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n154 ) , .A2( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U49 (.A2( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n135 ) , .A1( u0_u5_u1_n99 ) );
  AOI211_X1 u0_u5_u1_U5 (.ZN( u0_u5_u1_n124 ) , .A( u0_u5_u1_n138 ) , .C2( u0_u5_u1_n139 ) , .B( u0_u5_u1_n145 ) , .C1( u0_u5_u1_n147 ) );
  AOI21_X1 u0_u5_u1_U50 (.A( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n153 ) , .B1( u0_u5_u1_n154 ) , .ZN( u0_u5_u1_n158 ) );
  INV_X1 u0_u5_u1_U51 (.A( u0_u5_u1_n160 ) , .ZN( u0_u5_u1_n175 ) );
  NAND2_X1 u0_u5_u1_U52 (.A1( u0_u5_u1_n100 ) , .ZN( u0_u5_u1_n116 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U53 (.A1( u0_u5_u1_n102 ) , .ZN( u0_u5_u1_n131 ) , .A2( u0_u5_u1_n95 ) );
  NAND2_X1 u0_u5_u1_U54 (.A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n121 ) , .A1( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U55 (.A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n153 ) , .A2( u0_u5_u1_n98 ) );
  NAND2_X1 u0_u5_u1_U56 (.A2( u0_u5_u1_n104 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n133 ) );
  NAND2_X1 u0_u5_u1_U57 (.ZN( u0_u5_u1_n150 ) , .A2( u0_u5_u1_n98 ) , .A1( u0_u5_u1_n99 ) );
  NAND2_X1 u0_u5_u1_U58 (.A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n155 ) , .A2( u0_u5_u1_n95 ) );
  OAI21_X1 u0_u5_u1_U59 (.ZN( u0_u5_u1_n109 ) , .B1( u0_u5_u1_n129 ) , .B2( u0_u5_u1_n160 ) , .A( u0_u5_u1_n167 ) );
  AOI22_X1 u0_u5_u1_U6 (.B2( u0_u5_u1_n136 ) , .A2( u0_u5_u1_n137 ) , .ZN( u0_u5_u1_n143 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  NAND2_X1 u0_u5_u1_U60 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n120 ) );
  NAND2_X1 u0_u5_u1_U61 (.A1( u0_u5_u1_n102 ) , .A2( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n115 ) );
  NAND2_X1 u0_u5_u1_U62 (.A2( u0_u5_u1_n100 ) , .A1( u0_u5_u1_n104 ) , .ZN( u0_u5_u1_n151 ) );
  NAND2_X1 u0_u5_u1_U63 (.A2( u0_u5_u1_n103 ) , .A1( u0_u5_u1_n105 ) , .ZN( u0_u5_u1_n161 ) );
  INV_X1 u0_u5_u1_U64 (.A( u0_u5_u1_n152 ) , .ZN( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U65 (.A( u0_u5_u1_n128 ) , .ZN( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U66 (.A2( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n103 ) , .ZN( u0_u5_u1_n123 ) );
  AOI211_X1 u0_u5_u1_U67 (.B( u0_u5_u1_n162 ) , .A( u0_u5_u1_n163 ) , .C2( u0_u5_u1_n164 ) , .ZN( u0_u5_u1_n165 ) , .C1( u0_u5_u1_n171 ) );
  AOI21_X1 u0_u5_u1_U68 (.A( u0_u5_u1_n160 ) , .B2( u0_u5_u1_n161 ) , .ZN( u0_u5_u1_n162 ) , .B1( u0_u5_u1_n182 ) );
  OR2_X1 u0_u5_u1_U69 (.A2( u0_u5_u1_n157 ) , .A1( u0_u5_u1_n158 ) , .ZN( u0_u5_u1_n163 ) );
  INV_X1 u0_u5_u1_U7 (.A( u0_u5_u1_n147 ) , .ZN( u0_u5_u1_n181 ) );
  NOR2_X1 u0_u5_u1_U70 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n95 ) );
  NOR2_X1 u0_u5_u1_U71 (.A1( u0_u5_X_12 ) , .A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n100 ) );
  NOR2_X1 u0_u5_u1_U72 (.A2( u0_u5_X_8 ) , .A1( u0_u5_u1_n177 ) , .ZN( u0_u5_u1_n99 ) );
  NOR2_X1 u0_u5_u1_U73 (.A2( u0_u5_X_12 ) , .ZN( u0_u5_u1_n102 ) , .A1( u0_u5_u1_n176 ) );
  NOR2_X1 u0_u5_u1_U74 (.A2( u0_u5_X_9 ) , .ZN( u0_u5_u1_n105 ) , .A1( u0_u5_u1_n168 ) );
  NAND2_X1 u0_u5_u1_U75 (.A1( u0_u5_X_10 ) , .ZN( u0_u5_u1_n160 ) , .A2( u0_u5_u1_n169 ) );
  NAND2_X1 u0_u5_u1_U76 (.A2( u0_u5_X_10 ) , .A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n152 ) );
  NAND2_X1 u0_u5_u1_U77 (.A1( u0_u5_X_11 ) , .ZN( u0_u5_u1_n128 ) , .A2( u0_u5_u1_n170 ) );
  AND2_X1 u0_u5_u1_U78 (.A2( u0_u5_X_7 ) , .A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n104 ) );
  AND2_X1 u0_u5_u1_U79 (.A1( u0_u5_X_8 ) , .ZN( u0_u5_u1_n103 ) , .A2( u0_u5_u1_n177 ) );
  AOI22_X1 u0_u5_u1_U8 (.B2( u0_u5_u1_n113 ) , .A2( u0_u5_u1_n114 ) , .ZN( u0_u5_u1_n125 ) , .A1( u0_u5_u1_n171 ) , .B1( u0_u5_u1_n173 ) );
  INV_X1 u0_u5_u1_U80 (.A( u0_u5_X_10 ) , .ZN( u0_u5_u1_n170 ) );
  INV_X1 u0_u5_u1_U81 (.A( u0_u5_X_9 ) , .ZN( u0_u5_u1_n176 ) );
  INV_X1 u0_u5_u1_U82 (.A( u0_u5_X_11 ) , .ZN( u0_u5_u1_n169 ) );
  INV_X1 u0_u5_u1_U83 (.A( u0_u5_X_12 ) , .ZN( u0_u5_u1_n168 ) );
  INV_X1 u0_u5_u1_U84 (.A( u0_u5_X_7 ) , .ZN( u0_u5_u1_n177 ) );
  NAND4_X1 u0_u5_u1_U85 (.ZN( u0_out5_28 ) , .A4( u0_u5_u1_n124 ) , .A3( u0_u5_u1_n125 ) , .A2( u0_u5_u1_n126 ) , .A1( u0_u5_u1_n127 ) );
  OAI21_X1 u0_u5_u1_U86 (.ZN( u0_u5_u1_n127 ) , .B2( u0_u5_u1_n139 ) , .B1( u0_u5_u1_n175 ) , .A( u0_u5_u1_n183 ) );
  OAI21_X1 u0_u5_u1_U87 (.ZN( u0_u5_u1_n126 ) , .B2( u0_u5_u1_n140 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n178 ) );
  NAND4_X1 u0_u5_u1_U88 (.ZN( u0_out5_18 ) , .A4( u0_u5_u1_n165 ) , .A3( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n167 ) , .A2( u0_u5_u1_n186 ) );
  AOI22_X1 u0_u5_u1_U89 (.B2( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n147 ) , .A2( u0_u5_u1_n148 ) , .ZN( u0_u5_u1_n166 ) , .A1( u0_u5_u1_n172 ) );
  NAND2_X1 u0_u5_u1_U9 (.ZN( u0_u5_u1_n114 ) , .A1( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n156 ) );
  INV_X1 u0_u5_u1_U90 (.A( u0_u5_u1_n145 ) , .ZN( u0_u5_u1_n186 ) );
  NAND4_X1 u0_u5_u1_U91 (.ZN( u0_out5_2 ) , .A4( u0_u5_u1_n142 ) , .A3( u0_u5_u1_n143 ) , .A2( u0_u5_u1_n144 ) , .A1( u0_u5_u1_n179 ) );
  OAI21_X1 u0_u5_u1_U92 (.B2( u0_u5_u1_n132 ) , .ZN( u0_u5_u1_n144 ) , .A( u0_u5_u1_n146 ) , .B1( u0_u5_u1_n180 ) );
  INV_X1 u0_u5_u1_U93 (.A( u0_u5_u1_n130 ) , .ZN( u0_u5_u1_n179 ) );
  OR4_X1 u0_u5_u1_U94 (.ZN( u0_out5_13 ) , .A4( u0_u5_u1_n108 ) , .A3( u0_u5_u1_n109 ) , .A2( u0_u5_u1_n110 ) , .A1( u0_u5_u1_n111 ) );
  AOI21_X1 u0_u5_u1_U95 (.ZN( u0_u5_u1_n110 ) , .A( u0_u5_u1_n116 ) , .B1( u0_u5_u1_n152 ) , .B2( u0_u5_u1_n160 ) );
  AOI21_X1 u0_u5_u1_U96 (.ZN( u0_u5_u1_n111 ) , .A( u0_u5_u1_n128 ) , .B2( u0_u5_u1_n131 ) , .B1( u0_u5_u1_n135 ) );
  NAND3_X1 u0_u5_u1_U97 (.A3( u0_u5_u1_n149 ) , .A2( u0_u5_u1_n150 ) , .A1( u0_u5_u1_n151 ) , .ZN( u0_u5_u1_n164 ) );
  NAND3_X1 u0_u5_u1_U98 (.A3( u0_u5_u1_n134 ) , .A2( u0_u5_u1_n135 ) , .ZN( u0_u5_u1_n136 ) , .A1( u0_u5_u1_n151 ) );
  NAND3_X1 u0_u5_u1_U99 (.A1( u0_u5_u1_n133 ) , .ZN( u0_u5_u1_n137 ) , .A2( u0_u5_u1_n154 ) , .A3( u0_u5_u1_n181 ) );
  OAI22_X1 u0_u5_u2_U10 (.ZN( u0_u5_u2_n109 ) , .A2( u0_u5_u2_n113 ) , .B2( u0_u5_u2_n133 ) , .B1( u0_u5_u2_n167 ) , .A1( u0_u5_u2_n168 ) );
  NAND3_X1 u0_u5_u2_U100 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n98 ) );
  OAI22_X1 u0_u5_u2_U11 (.B1( u0_u5_u2_n151 ) , .A2( u0_u5_u2_n152 ) , .A1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n160 ) , .B2( u0_u5_u2_n168 ) );
  NOR3_X1 u0_u5_u2_U12 (.A1( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n151 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U13 (.ZN( u0_u5_u2_n144 ) , .B2( u0_u5_u2_n155 ) , .A( u0_u5_u2_n172 ) , .B1( u0_u5_u2_n185 ) );
  AOI21_X1 u0_u5_u2_U14 (.B2( u0_u5_u2_n143 ) , .ZN( u0_u5_u2_n145 ) , .B1( u0_u5_u2_n152 ) , .A( u0_u5_u2_n171 ) );
  AOI21_X1 u0_u5_u2_U15 (.B2( u0_u5_u2_n120 ) , .B1( u0_u5_u2_n121 ) , .ZN( u0_u5_u2_n126 ) , .A( u0_u5_u2_n167 ) );
  INV_X1 u0_u5_u2_U16 (.A( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n171 ) );
  INV_X1 u0_u5_u2_U17 (.A( u0_u5_u2_n120 ) , .ZN( u0_u5_u2_n188 ) );
  NAND2_X1 u0_u5_u2_U18 (.A2( u0_u5_u2_n122 ) , .ZN( u0_u5_u2_n150 ) , .A1( u0_u5_u2_n152 ) );
  INV_X1 u0_u5_u2_U19 (.A( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U20 (.A( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n173 ) );
  NAND2_X1 u0_u5_u2_U21 (.A1( u0_u5_u2_n132 ) , .A2( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n157 ) );
  INV_X1 u0_u5_u2_U22 (.A( u0_u5_u2_n113 ) , .ZN( u0_u5_u2_n178 ) );
  INV_X1 u0_u5_u2_U23 (.A( u0_u5_u2_n139 ) , .ZN( u0_u5_u2_n175 ) );
  INV_X1 u0_u5_u2_U24 (.A( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n181 ) );
  INV_X1 u0_u5_u2_U25 (.A( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n177 ) );
  INV_X1 u0_u5_u2_U26 (.A( u0_u5_u2_n116 ) , .ZN( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U27 (.A( u0_u5_u2_n131 ) , .ZN( u0_u5_u2_n179 ) );
  INV_X1 u0_u5_u2_U28 (.A( u0_u5_u2_n154 ) , .ZN( u0_u5_u2_n176 ) );
  NAND2_X1 u0_u5_u2_U29 (.A2( u0_u5_u2_n116 ) , .A1( u0_u5_u2_n117 ) , .ZN( u0_u5_u2_n118 ) );
  NOR2_X1 u0_u5_u2_U3 (.ZN( u0_u5_u2_n121 ) , .A2( u0_u5_u2_n177 ) , .A1( u0_u5_u2_n180 ) );
  INV_X1 u0_u5_u2_U30 (.A( u0_u5_u2_n132 ) , .ZN( u0_u5_u2_n182 ) );
  INV_X1 u0_u5_u2_U31 (.A( u0_u5_u2_n158 ) , .ZN( u0_u5_u2_n183 ) );
  OAI21_X1 u0_u5_u2_U32 (.A( u0_u5_u2_n156 ) , .B1( u0_u5_u2_n157 ) , .ZN( u0_u5_u2_n158 ) , .B2( u0_u5_u2_n179 ) );
  NOR2_X1 u0_u5_u2_U33 (.ZN( u0_u5_u2_n156 ) , .A1( u0_u5_u2_n166 ) , .A2( u0_u5_u2_n169 ) );
  NOR2_X1 u0_u5_u2_U34 (.A2( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n140 ) );
  NOR2_X1 u0_u5_u2_U35 (.A2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n153 ) , .A1( u0_u5_u2_n156 ) );
  AOI211_X1 u0_u5_u2_U36 (.ZN( u0_u5_u2_n130 ) , .C1( u0_u5_u2_n138 ) , .C2( u0_u5_u2_n179 ) , .B( u0_u5_u2_n96 ) , .A( u0_u5_u2_n97 ) );
  OAI22_X1 u0_u5_u2_U37 (.B1( u0_u5_u2_n133 ) , .A2( u0_u5_u2_n137 ) , .A1( u0_u5_u2_n152 ) , .B2( u0_u5_u2_n168 ) , .ZN( u0_u5_u2_n97 ) );
  OAI221_X1 u0_u5_u2_U38 (.B1( u0_u5_u2_n113 ) , .C1( u0_u5_u2_n132 ) , .A( u0_u5_u2_n149 ) , .B2( u0_u5_u2_n171 ) , .C2( u0_u5_u2_n172 ) , .ZN( u0_u5_u2_n96 ) );
  OAI221_X1 u0_u5_u2_U39 (.A( u0_u5_u2_n115 ) , .C2( u0_u5_u2_n123 ) , .B2( u0_u5_u2_n143 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n163 ) , .C1( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U4 (.A( u0_u5_u2_n134 ) , .ZN( u0_u5_u2_n185 ) );
  OAI21_X1 u0_u5_u2_U40 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n115 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n178 ) );
  OAI221_X1 u0_u5_u2_U41 (.A( u0_u5_u2_n135 ) , .B2( u0_u5_u2_n136 ) , .B1( u0_u5_u2_n137 ) , .ZN( u0_u5_u2_n162 ) , .C2( u0_u5_u2_n167 ) , .C1( u0_u5_u2_n185 ) );
  AND3_X1 u0_u5_u2_U42 (.A3( u0_u5_u2_n131 ) , .A2( u0_u5_u2_n132 ) , .A1( u0_u5_u2_n133 ) , .ZN( u0_u5_u2_n136 ) );
  AOI22_X1 u0_u5_u2_U43 (.ZN( u0_u5_u2_n135 ) , .B1( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n156 ) , .B2( u0_u5_u2_n180 ) , .A2( u0_u5_u2_n188 ) );
  AOI21_X1 u0_u5_u2_U44 (.ZN( u0_u5_u2_n149 ) , .B1( u0_u5_u2_n173 ) , .B2( u0_u5_u2_n188 ) , .A( u0_u5_u2_n95 ) );
  AND3_X1 u0_u5_u2_U45 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n156 ) , .ZN( u0_u5_u2_n95 ) );
  OAI21_X1 u0_u5_u2_U46 (.A( u0_u5_u2_n141 ) , .B2( u0_u5_u2_n142 ) , .ZN( u0_u5_u2_n146 ) , .B1( u0_u5_u2_n153 ) );
  OAI21_X1 u0_u5_u2_U47 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n141 ) , .B1( u0_u5_u2_n176 ) , .B2( u0_u5_u2_n177 ) );
  NOR3_X1 u0_u5_u2_U48 (.ZN( u0_u5_u2_n142 ) , .A3( u0_u5_u2_n175 ) , .A2( u0_u5_u2_n178 ) , .A1( u0_u5_u2_n181 ) );
  OAI21_X1 u0_u5_u2_U49 (.A( u0_u5_u2_n101 ) , .B2( u0_u5_u2_n121 ) , .B1( u0_u5_u2_n153 ) , .ZN( u0_u5_u2_n164 ) );
  INV_X1 u0_u5_u2_U5 (.A( u0_u5_u2_n150 ) , .ZN( u0_u5_u2_n184 ) );
  NAND2_X1 u0_u5_u2_U50 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n155 ) );
  NAND2_X1 u0_u5_u2_U51 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n143 ) );
  NAND2_X1 u0_u5_u2_U52 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n152 ) );
  NAND2_X1 u0_u5_u2_U53 (.A1( u0_u5_u2_n100 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n132 ) );
  INV_X1 u0_u5_u2_U54 (.A( u0_u5_u2_n140 ) , .ZN( u0_u5_u2_n168 ) );
  INV_X1 u0_u5_u2_U55 (.A( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n167 ) );
  NAND2_X1 u0_u5_u2_U56 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n113 ) );
  NAND2_X1 u0_u5_u2_U57 (.A1( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n131 ) );
  NAND2_X1 u0_u5_u2_U58 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n107 ) , .ZN( u0_u5_u2_n139 ) );
  NAND2_X1 u0_u5_u2_U59 (.A1( u0_u5_u2_n103 ) , .A2( u0_u5_u2_n105 ) , .ZN( u0_u5_u2_n133 ) );
  NOR4_X1 u0_u5_u2_U6 (.A4( u0_u5_u2_n124 ) , .A3( u0_u5_u2_n125 ) , .A2( u0_u5_u2_n126 ) , .A1( u0_u5_u2_n127 ) , .ZN( u0_u5_u2_n128 ) );
  NAND2_X1 u0_u5_u2_U60 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n103 ) , .ZN( u0_u5_u2_n154 ) );
  NAND2_X1 u0_u5_u2_U61 (.A2( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n104 ) , .ZN( u0_u5_u2_n119 ) );
  NAND2_X1 u0_u5_u2_U62 (.A2( u0_u5_u2_n107 ) , .A1( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n123 ) );
  NAND2_X1 u0_u5_u2_U63 (.A1( u0_u5_u2_n104 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n122 ) );
  INV_X1 u0_u5_u2_U64 (.A( u0_u5_u2_n114 ) , .ZN( u0_u5_u2_n172 ) );
  NAND2_X1 u0_u5_u2_U65 (.A2( u0_u5_u2_n100 ) , .A1( u0_u5_u2_n102 ) , .ZN( u0_u5_u2_n116 ) );
  NAND2_X1 u0_u5_u2_U66 (.A1( u0_u5_u2_n102 ) , .A2( u0_u5_u2_n108 ) , .ZN( u0_u5_u2_n120 ) );
  NAND2_X1 u0_u5_u2_U67 (.A2( u0_u5_u2_n105 ) , .A1( u0_u5_u2_n106 ) , .ZN( u0_u5_u2_n117 ) );
  INV_X1 u0_u5_u2_U68 (.ZN( u0_u5_u2_n187 ) , .A( u0_u5_u2_n99 ) );
  OAI21_X1 u0_u5_u2_U69 (.B1( u0_u5_u2_n137 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n98 ) , .ZN( u0_u5_u2_n99 ) );
  AOI21_X1 u0_u5_u2_U7 (.B2( u0_u5_u2_n119 ) , .ZN( u0_u5_u2_n127 ) , .A( u0_u5_u2_n137 ) , .B1( u0_u5_u2_n155 ) );
  NOR2_X1 u0_u5_u2_U70 (.A2( u0_u5_X_16 ) , .ZN( u0_u5_u2_n140 ) , .A1( u0_u5_u2_n166 ) );
  NOR2_X1 u0_u5_u2_U71 (.A2( u0_u5_X_13 ) , .A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n100 ) );
  NOR2_X1 u0_u5_u2_U72 (.A2( u0_u5_X_16 ) , .A1( u0_u5_X_17 ) , .ZN( u0_u5_u2_n138 ) );
  NOR2_X1 u0_u5_u2_U73 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n104 ) );
  NOR2_X1 u0_u5_u2_U74 (.A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n103 ) , .A1( u0_u5_u2_n174 ) );
  NOR2_X1 u0_u5_u2_U75 (.A2( u0_u5_X_15 ) , .ZN( u0_u5_u2_n102 ) , .A1( u0_u5_u2_n165 ) );
  NOR2_X1 u0_u5_u2_U76 (.A2( u0_u5_X_17 ) , .ZN( u0_u5_u2_n114 ) , .A1( u0_u5_u2_n169 ) );
  AND2_X1 u0_u5_u2_U77 (.A1( u0_u5_X_15 ) , .ZN( u0_u5_u2_n105 ) , .A2( u0_u5_u2_n165 ) );
  AND2_X1 u0_u5_u2_U78 (.A2( u0_u5_X_15 ) , .A1( u0_u5_X_18 ) , .ZN( u0_u5_u2_n107 ) );
  AND2_X1 u0_u5_u2_U79 (.A1( u0_u5_X_14 ) , .ZN( u0_u5_u2_n106 ) , .A2( u0_u5_u2_n174 ) );
  AOI21_X1 u0_u5_u2_U8 (.ZN( u0_u5_u2_n124 ) , .B1( u0_u5_u2_n131 ) , .B2( u0_u5_u2_n143 ) , .A( u0_u5_u2_n172 ) );
  AND2_X1 u0_u5_u2_U80 (.A1( u0_u5_X_13 ) , .A2( u0_u5_X_14 ) , .ZN( u0_u5_u2_n108 ) );
  INV_X1 u0_u5_u2_U81 (.A( u0_u5_X_16 ) , .ZN( u0_u5_u2_n169 ) );
  INV_X1 u0_u5_u2_U82 (.A( u0_u5_X_17 ) , .ZN( u0_u5_u2_n166 ) );
  INV_X1 u0_u5_u2_U83 (.A( u0_u5_X_13 ) , .ZN( u0_u5_u2_n174 ) );
  INV_X1 u0_u5_u2_U84 (.A( u0_u5_X_18 ) , .ZN( u0_u5_u2_n165 ) );
  NAND4_X1 u0_u5_u2_U85 (.ZN( u0_out5_30 ) , .A4( u0_u5_u2_n147 ) , .A3( u0_u5_u2_n148 ) , .A2( u0_u5_u2_n149 ) , .A1( u0_u5_u2_n187 ) );
  NOR3_X1 u0_u5_u2_U86 (.A3( u0_u5_u2_n144 ) , .A2( u0_u5_u2_n145 ) , .A1( u0_u5_u2_n146 ) , .ZN( u0_u5_u2_n147 ) );
  AOI21_X1 u0_u5_u2_U87 (.B2( u0_u5_u2_n138 ) , .ZN( u0_u5_u2_n148 ) , .A( u0_u5_u2_n162 ) , .B1( u0_u5_u2_n182 ) );
  NAND4_X1 u0_u5_u2_U88 (.ZN( u0_out5_24 ) , .A4( u0_u5_u2_n111 ) , .A3( u0_u5_u2_n112 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n187 ) );
  AOI221_X1 u0_u5_u2_U89 (.A( u0_u5_u2_n109 ) , .B1( u0_u5_u2_n110 ) , .ZN( u0_u5_u2_n111 ) , .C1( u0_u5_u2_n134 ) , .C2( u0_u5_u2_n170 ) , .B2( u0_u5_u2_n173 ) );
  AOI21_X1 u0_u5_u2_U9 (.B2( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n125 ) , .A( u0_u5_u2_n171 ) , .B1( u0_u5_u2_n184 ) );
  AOI21_X1 u0_u5_u2_U90 (.ZN( u0_u5_u2_n112 ) , .B2( u0_u5_u2_n156 ) , .A( u0_u5_u2_n164 ) , .B1( u0_u5_u2_n181 ) );
  NAND4_X1 u0_u5_u2_U91 (.ZN( u0_out5_16 ) , .A4( u0_u5_u2_n128 ) , .A3( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n130 ) , .A2( u0_u5_u2_n186 ) );
  AOI22_X1 u0_u5_u2_U92 (.A2( u0_u5_u2_n118 ) , .ZN( u0_u5_u2_n129 ) , .A1( u0_u5_u2_n140 ) , .B1( u0_u5_u2_n157 ) , .B2( u0_u5_u2_n170 ) );
  INV_X1 u0_u5_u2_U93 (.A( u0_u5_u2_n163 ) , .ZN( u0_u5_u2_n186 ) );
  OR4_X1 u0_u5_u2_U94 (.ZN( u0_out5_6 ) , .A4( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n162 ) , .A2( u0_u5_u2_n163 ) , .A1( u0_u5_u2_n164 ) );
  OR3_X1 u0_u5_u2_U95 (.A2( u0_u5_u2_n159 ) , .A1( u0_u5_u2_n160 ) , .ZN( u0_u5_u2_n161 ) , .A3( u0_u5_u2_n183 ) );
  AOI21_X1 u0_u5_u2_U96 (.B2( u0_u5_u2_n154 ) , .B1( u0_u5_u2_n155 ) , .ZN( u0_u5_u2_n159 ) , .A( u0_u5_u2_n167 ) );
  NAND3_X1 u0_u5_u2_U97 (.A2( u0_u5_u2_n117 ) , .A1( u0_u5_u2_n122 ) , .A3( u0_u5_u2_n123 ) , .ZN( u0_u5_u2_n134 ) );
  NAND3_X1 u0_u5_u2_U98 (.ZN( u0_u5_u2_n110 ) , .A2( u0_u5_u2_n131 ) , .A3( u0_u5_u2_n139 ) , .A1( u0_u5_u2_n154 ) );
  NAND3_X1 u0_u5_u2_U99 (.A2( u0_u5_u2_n100 ) , .ZN( u0_u5_u2_n101 ) , .A1( u0_u5_u2_n104 ) , .A3( u0_u5_u2_n114 ) );
  OAI22_X1 u0_u5_u3_U10 (.B1( u0_u5_u3_n113 ) , .A2( u0_u5_u3_n135 ) , .A1( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n164 ) , .ZN( u0_u5_u3_n98 ) );
  OAI211_X1 u0_u5_u3_U11 (.B( u0_u5_u3_n106 ) , .ZN( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n128 ) , .C1( u0_u5_u3_n167 ) , .A( u0_u5_u3_n181 ) );
  AOI221_X1 u0_u5_u3_U12 (.C1( u0_u5_u3_n105 ) , .ZN( u0_u5_u3_n106 ) , .A( u0_u5_u3_n131 ) , .B2( u0_u5_u3_n132 ) , .C2( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n169 ) );
  INV_X1 u0_u5_u3_U13 (.ZN( u0_u5_u3_n181 ) , .A( u0_u5_u3_n98 ) );
  NAND2_X1 u0_u5_u3_U14 (.ZN( u0_u5_u3_n105 ) , .A2( u0_u5_u3_n130 ) , .A1( u0_u5_u3_n155 ) );
  AOI22_X1 u0_u5_u3_U15 (.B1( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n116 ) , .ZN( u0_u5_u3_n123 ) , .B2( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U16 (.ZN( u0_u5_u3_n116 ) , .A2( u0_u5_u3_n151 ) , .A1( u0_u5_u3_n182 ) );
  NOR2_X1 u0_u5_u3_U17 (.ZN( u0_u5_u3_n126 ) , .A2( u0_u5_u3_n150 ) , .A1( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U18 (.ZN( u0_u5_u3_n112 ) , .B2( u0_u5_u3_n146 ) , .B1( u0_u5_u3_n155 ) , .A( u0_u5_u3_n167 ) );
  NAND2_X1 u0_u5_u3_U19 (.A1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n142 ) , .A2( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U20 (.ZN( u0_u5_u3_n132 ) , .A2( u0_u5_u3_n152 ) , .A1( u0_u5_u3_n156 ) );
  AND2_X1 u0_u5_u3_U21 (.A2( u0_u5_u3_n113 ) , .A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n151 ) );
  INV_X1 u0_u5_u3_U22 (.A( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n165 ) );
  INV_X1 u0_u5_u3_U23 (.A( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n170 ) );
  NAND2_X1 u0_u5_u3_U24 (.A1( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .ZN( u0_u5_u3_n140 ) );
  NAND2_X1 u0_u5_u3_U25 (.ZN( u0_u5_u3_n117 ) , .A1( u0_u5_u3_n124 ) , .A2( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U26 (.ZN( u0_u5_u3_n143 ) , .A1( u0_u5_u3_n165 ) , .A2( u0_u5_u3_n167 ) );
  INV_X1 u0_u5_u3_U27 (.A( u0_u5_u3_n130 ) , .ZN( u0_u5_u3_n177 ) );
  INV_X1 u0_u5_u3_U28 (.A( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n176 ) );
  INV_X1 u0_u5_u3_U29 (.A( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n174 ) );
  INV_X1 u0_u5_u3_U3 (.A( u0_u5_u3_n129 ) , .ZN( u0_u5_u3_n183 ) );
  INV_X1 u0_u5_u3_U30 (.A( u0_u5_u3_n139 ) , .ZN( u0_u5_u3_n185 ) );
  NOR2_X1 u0_u5_u3_U31 (.ZN( u0_u5_u3_n135 ) , .A2( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n169 ) );
  OAI222_X1 u0_u5_u3_U32 (.C2( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .B1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n138 ) , .B2( u0_u5_u3_n146 ) , .C1( u0_u5_u3_n154 ) , .A1( u0_u5_u3_n164 ) );
  NOR4_X1 u0_u5_u3_U33 (.A4( u0_u5_u3_n157 ) , .A3( u0_u5_u3_n158 ) , .A2( u0_u5_u3_n159 ) , .A1( u0_u5_u3_n160 ) , .ZN( u0_u5_u3_n161 ) );
  AOI21_X1 u0_u5_u3_U34 (.B2( u0_u5_u3_n152 ) , .B1( u0_u5_u3_n153 ) , .ZN( u0_u5_u3_n158 ) , .A( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U35 (.A( u0_u5_u3_n154 ) , .B2( u0_u5_u3_n155 ) , .B1( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n157 ) );
  AOI21_X1 u0_u5_u3_U36 (.A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n150 ) , .B1( u0_u5_u3_n151 ) , .ZN( u0_u5_u3_n159 ) );
  AOI211_X1 u0_u5_u3_U37 (.ZN( u0_u5_u3_n109 ) , .A( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n129 ) , .B( u0_u5_u3_n138 ) , .C1( u0_u5_u3_n141 ) );
  AOI211_X1 u0_u5_u3_U38 (.B( u0_u5_u3_n119 ) , .A( u0_u5_u3_n120 ) , .C2( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n122 ) , .C1( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U39 (.A( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U4 (.A( u0_u5_u3_n140 ) , .ZN( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u3_U40 (.B1( u0_u5_u3_n118 ) , .ZN( u0_u5_u3_n120 ) , .A1( u0_u5_u3_n135 ) , .B2( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n178 ) );
  AND3_X1 u0_u5_u3_U41 (.ZN( u0_u5_u3_n118 ) , .A2( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n144 ) , .A3( u0_u5_u3_n152 ) );
  INV_X1 u0_u5_u3_U42 (.A( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U43 (.ZN( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n164 ) );
  OAI211_X1 u0_u5_u3_U44 (.B( u0_u5_u3_n127 ) , .ZN( u0_u5_u3_n139 ) , .C1( u0_u5_u3_n150 ) , .C2( u0_u5_u3_n154 ) , .A( u0_u5_u3_n184 ) );
  INV_X1 u0_u5_u3_U45 (.A( u0_u5_u3_n125 ) , .ZN( u0_u5_u3_n184 ) );
  AOI221_X1 u0_u5_u3_U46 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n127 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n169 ) , .B2( u0_u5_u3_n170 ) , .B1( u0_u5_u3_n174 ) );
  OAI22_X1 u0_u5_u3_U47 (.A1( u0_u5_u3_n124 ) , .ZN( u0_u5_u3_n125 ) , .B2( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n165 ) , .B1( u0_u5_u3_n167 ) );
  NOR2_X1 u0_u5_u3_U48 (.A1( u0_u5_u3_n113 ) , .ZN( u0_u5_u3_n131 ) , .A2( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U49 (.A1( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n150 ) , .A2( u0_u5_u3_n99 ) );
  INV_X1 u0_u5_u3_U5 (.A( u0_u5_u3_n117 ) , .ZN( u0_u5_u3_n178 ) );
  NAND2_X1 u0_u5_u3_U50 (.A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n155 ) , .A1( u0_u5_u3_n97 ) );
  INV_X1 u0_u5_u3_U51 (.A( u0_u5_u3_n141 ) , .ZN( u0_u5_u3_n167 ) );
  AOI21_X1 u0_u5_u3_U52 (.B2( u0_u5_u3_n114 ) , .B1( u0_u5_u3_n146 ) , .A( u0_u5_u3_n154 ) , .ZN( u0_u5_u3_n94 ) );
  AOI21_X1 u0_u5_u3_U53 (.ZN( u0_u5_u3_n110 ) , .B2( u0_u5_u3_n142 ) , .B1( u0_u5_u3_n186 ) , .A( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U54 (.A( u0_u5_u3_n145 ) , .ZN( u0_u5_u3_n186 ) );
  AOI21_X1 u0_u5_u3_U55 (.B1( u0_u5_u3_n124 ) , .A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U56 (.A( u0_u5_u3_n149 ) , .ZN( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U57 (.ZN( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n96 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U58 (.A2( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n146 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U59 (.A1( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n99 ) );
  AOI221_X1 u0_u5_u3_U6 (.A( u0_u5_u3_n131 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n134 ) , .B1( u0_u5_u3_n143 ) , .B2( u0_u5_u3_n177 ) );
  NAND2_X1 u0_u5_u3_U60 (.A1( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n156 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U61 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U62 (.A1( u0_u5_u3_n100 ) , .A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n128 ) );
  NAND2_X1 u0_u5_u3_U63 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n152 ) );
  NAND2_X1 u0_u5_u3_U64 (.A2( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n114 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U65 (.ZN( u0_u5_u3_n107 ) , .A1( u0_u5_u3_n97 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U66 (.A2( u0_u5_u3_n100 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n113 ) );
  NAND2_X1 u0_u5_u3_U67 (.A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n153 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U68 (.A2( u0_u5_u3_n103 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n130 ) );
  NAND2_X1 u0_u5_u3_U69 (.A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n96 ) );
  OAI22_X1 u0_u5_u3_U7 (.B2( u0_u5_u3_n147 ) , .A2( u0_u5_u3_n148 ) , .ZN( u0_u5_u3_n160 ) , .B1( u0_u5_u3_n165 ) , .A1( u0_u5_u3_n168 ) );
  NAND2_X1 u0_u5_u3_U70 (.A1( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n108 ) );
  NOR2_X1 u0_u5_u3_U71 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n99 ) );
  NOR2_X1 u0_u5_u3_U72 (.A2( u0_u5_X_21 ) , .A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n103 ) );
  NOR2_X1 u0_u5_u3_U73 (.A2( u0_u5_X_24 ) , .A1( u0_u5_u3_n171 ) , .ZN( u0_u5_u3_n97 ) );
  NOR2_X1 u0_u5_u3_U74 (.A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U75 (.A2( u0_u5_X_19 ) , .A1( u0_u5_u3_n172 ) , .ZN( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U76 (.A1( u0_u5_X_22 ) , .A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U77 (.A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n149 ) , .A2( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U78 (.A2( u0_u5_X_22 ) , .A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n121 ) );
  AND2_X1 u0_u5_u3_U79 (.A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n101 ) , .A2( u0_u5_u3_n171 ) );
  AND3_X1 u0_u5_u3_U8 (.A3( u0_u5_u3_n144 ) , .A2( u0_u5_u3_n145 ) , .A1( u0_u5_u3_n146 ) , .ZN( u0_u5_u3_n147 ) );
  AND2_X1 u0_u5_u3_U80 (.A1( u0_u5_X_19 ) , .ZN( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n172 ) );
  AND2_X1 u0_u5_u3_U81 (.A1( u0_u5_X_21 ) , .A2( u0_u5_X_24 ) , .ZN( u0_u5_u3_n100 ) );
  AND2_X1 u0_u5_u3_U82 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n104 ) );
  INV_X1 u0_u5_u3_U83 (.A( u0_u5_X_22 ) , .ZN( u0_u5_u3_n166 ) );
  INV_X1 u0_u5_u3_U84 (.A( u0_u5_X_21 ) , .ZN( u0_u5_u3_n171 ) );
  INV_X1 u0_u5_u3_U85 (.A( u0_u5_X_20 ) , .ZN( u0_u5_u3_n172 ) );
  NAND4_X1 u0_u5_u3_U86 (.ZN( u0_out5_26 ) , .A4( u0_u5_u3_n109 ) , .A3( u0_u5_u3_n110 ) , .A2( u0_u5_u3_n111 ) , .A1( u0_u5_u3_n173 ) );
  INV_X1 u0_u5_u3_U87 (.ZN( u0_u5_u3_n173 ) , .A( u0_u5_u3_n94 ) );
  OAI21_X1 u0_u5_u3_U88 (.ZN( u0_u5_u3_n111 ) , .B2( u0_u5_u3_n117 ) , .A( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n176 ) );
  NAND4_X1 u0_u5_u3_U89 (.ZN( u0_out5_20 ) , .A4( u0_u5_u3_n122 ) , .A3( u0_u5_u3_n123 ) , .A1( u0_u5_u3_n175 ) , .A2( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U9 (.A( u0_u5_u3_n143 ) , .ZN( u0_u5_u3_n168 ) );
  INV_X1 u0_u5_u3_U90 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U91 (.A( u0_u5_u3_n112 ) , .ZN( u0_u5_u3_n175 ) );
  NAND4_X1 u0_u5_u3_U92 (.ZN( u0_out5_1 ) , .A4( u0_u5_u3_n161 ) , .A3( u0_u5_u3_n162 ) , .A2( u0_u5_u3_n163 ) , .A1( u0_u5_u3_n185 ) );
  NAND2_X1 u0_u5_u3_U93 (.ZN( u0_u5_u3_n163 ) , .A2( u0_u5_u3_n170 ) , .A1( u0_u5_u3_n176 ) );
  AOI22_X1 u0_u5_u3_U94 (.B2( u0_u5_u3_n140 ) , .B1( u0_u5_u3_n141 ) , .A2( u0_u5_u3_n142 ) , .ZN( u0_u5_u3_n162 ) , .A1( u0_u5_u3_n177 ) );
  OR4_X1 u0_u5_u3_U95 (.ZN( u0_out5_10 ) , .A4( u0_u5_u3_n136 ) , .A3( u0_u5_u3_n137 ) , .A1( u0_u5_u3_n138 ) , .A2( u0_u5_u3_n139 ) );
  OAI222_X1 u0_u5_u3_U96 (.C1( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n137 ) , .B1( u0_u5_u3_n148 ) , .A2( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n154 ) , .C2( u0_u5_u3_n164 ) , .A1( u0_u5_u3_n167 ) );
  OAI221_X1 u0_u5_u3_U97 (.A( u0_u5_u3_n134 ) , .B2( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n136 ) , .C1( u0_u5_u3_n149 ) , .B1( u0_u5_u3_n151 ) , .C2( u0_u5_u3_n183 ) );
  NAND3_X1 u0_u5_u3_U98 (.A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n145 ) , .A3( u0_u5_u3_n153 ) );
  NAND3_X1 u0_u5_u3_U99 (.ZN( u0_u5_u3_n129 ) , .A2( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n153 ) , .A3( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u4_U10 (.B2( u0_u5_u4_n135 ) , .ZN( u0_u5_u4_n137 ) , .B1( u0_u5_u4_n153 ) , .A1( u0_u5_u4_n155 ) , .A2( u0_u5_u4_n171 ) );
  AND3_X1 u0_u5_u4_U11 (.A2( u0_u5_u4_n134 ) , .ZN( u0_u5_u4_n135 ) , .A3( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n157 ) );
  NAND2_X1 u0_u5_u4_U12 (.ZN( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n173 ) );
  AOI21_X1 u0_u5_u4_U13 (.B2( u0_u5_u4_n160 ) , .B1( u0_u5_u4_n161 ) , .ZN( u0_u5_u4_n162 ) , .A( u0_u5_u4_n170 ) );
  AOI21_X1 u0_u5_u4_U14 (.ZN( u0_u5_u4_n107 ) , .B2( u0_u5_u4_n143 ) , .A( u0_u5_u4_n174 ) , .B1( u0_u5_u4_n184 ) );
  AOI21_X1 u0_u5_u4_U15 (.B2( u0_u5_u4_n158 ) , .B1( u0_u5_u4_n159 ) , .ZN( u0_u5_u4_n163 ) , .A( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U16 (.A( u0_u5_u4_n153 ) , .B2( u0_u5_u4_n154 ) , .B1( u0_u5_u4_n155 ) , .ZN( u0_u5_u4_n165 ) );
  AOI21_X1 u0_u5_u4_U17 (.A( u0_u5_u4_n156 ) , .B2( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n164 ) , .B1( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U18 (.A( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n170 ) );
  AND2_X1 u0_u5_u4_U19 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n155 ) , .A1( u0_u5_u4_n160 ) );
  INV_X1 u0_u5_u4_U20 (.A( u0_u5_u4_n156 ) , .ZN( u0_u5_u4_n175 ) );
  NAND2_X1 u0_u5_u4_U21 (.A2( u0_u5_u4_n118 ) , .ZN( u0_u5_u4_n131 ) , .A1( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U22 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n130 ) );
  NAND2_X1 u0_u5_u4_U23 (.ZN( u0_u5_u4_n117 ) , .A2( u0_u5_u4_n118 ) , .A1( u0_u5_u4_n148 ) );
  NAND2_X1 u0_u5_u4_U24 (.ZN( u0_u5_u4_n129 ) , .A1( u0_u5_u4_n134 ) , .A2( u0_u5_u4_n148 ) );
  AND3_X1 u0_u5_u4_U25 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n143 ) , .A3( u0_u5_u4_n154 ) , .ZN( u0_u5_u4_n161 ) );
  AND2_X1 u0_u5_u4_U26 (.A1( u0_u5_u4_n145 ) , .A2( u0_u5_u4_n147 ) , .ZN( u0_u5_u4_n159 ) );
  OR3_X1 u0_u5_u4_U27 (.A3( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n115 ) , .A1( u0_u5_u4_n116 ) , .ZN( u0_u5_u4_n136 ) );
  AOI21_X1 u0_u5_u4_U28 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n116 ) , .B2( u0_u5_u4_n173 ) , .B1( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U29 (.ZN( u0_u5_u4_n115 ) , .B2( u0_u5_u4_n145 ) , .B1( u0_u5_u4_n146 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U3 (.ZN( u0_u5_u4_n121 ) , .A1( u0_u5_u4_n181 ) , .A2( u0_u5_u4_n182 ) );
  OAI22_X1 u0_u5_u4_U30 (.ZN( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n121 ) , .B1( u0_u5_u4_n160 ) , .B2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n171 ) );
  INV_X1 u0_u5_u4_U31 (.A( u0_u5_u4_n158 ) , .ZN( u0_u5_u4_n182 ) );
  INV_X1 u0_u5_u4_U32 (.ZN( u0_u5_u4_n181 ) , .A( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U33 (.A( u0_u5_u4_n144 ) , .ZN( u0_u5_u4_n179 ) );
  INV_X1 u0_u5_u4_U34 (.A( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n178 ) );
  NAND2_X1 u0_u5_u4_U35 (.A2( u0_u5_u4_n154 ) , .A1( u0_u5_u4_n96 ) , .ZN( u0_u5_u4_n97 ) );
  INV_X1 u0_u5_u4_U36 (.ZN( u0_u5_u4_n186 ) , .A( u0_u5_u4_n95 ) );
  OAI221_X1 u0_u5_u4_U37 (.C1( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n158 ) , .B2( u0_u5_u4_n171 ) , .C2( u0_u5_u4_n173 ) , .A( u0_u5_u4_n94 ) , .ZN( u0_u5_u4_n95 ) );
  AOI222_X1 u0_u5_u4_U38 (.B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n138 ) , .C2( u0_u5_u4_n175 ) , .A2( u0_u5_u4_n179 ) , .C1( u0_u5_u4_n181 ) , .B1( u0_u5_u4_n185 ) , .ZN( u0_u5_u4_n94 ) );
  INV_X1 u0_u5_u4_U39 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n185 ) );
  INV_X1 u0_u5_u4_U4 (.A( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U40 (.A( u0_u5_u4_n143 ) , .ZN( u0_u5_u4_n183 ) );
  NOR2_X1 u0_u5_u4_U41 (.ZN( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n168 ) , .A2( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U42 (.A1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n153 ) );
  NOR2_X1 u0_u5_u4_U43 (.A2( u0_u5_u4_n128 ) , .A1( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n156 ) );
  AOI22_X1 u0_u5_u4_U44 (.B2( u0_u5_u4_n122 ) , .A1( u0_u5_u4_n123 ) , .ZN( u0_u5_u4_n124 ) , .B1( u0_u5_u4_n128 ) , .A2( u0_u5_u4_n172 ) );
  INV_X1 u0_u5_u4_U45 (.A( u0_u5_u4_n153 ) , .ZN( u0_u5_u4_n172 ) );
  NAND2_X1 u0_u5_u4_U46 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n123 ) , .A1( u0_u5_u4_n161 ) );
  AOI22_X1 u0_u5_u4_U47 (.B2( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n133 ) , .ZN( u0_u5_u4_n140 ) , .A1( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n179 ) );
  NAND2_X1 u0_u5_u4_U48 (.ZN( u0_u5_u4_n133 ) , .A2( u0_u5_u4_n146 ) , .A1( u0_u5_u4_n154 ) );
  NAND2_X1 u0_u5_u4_U49 (.A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n154 ) , .A2( u0_u5_u4_n98 ) );
  NOR4_X1 u0_u5_u4_U5 (.A4( u0_u5_u4_n106 ) , .A3( u0_u5_u4_n107 ) , .A2( u0_u5_u4_n108 ) , .A1( u0_u5_u4_n109 ) , .ZN( u0_u5_u4_n110 ) );
  NAND2_X1 u0_u5_u4_U50 (.A1( u0_u5_u4_n101 ) , .ZN( u0_u5_u4_n158 ) , .A2( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U51 (.ZN( u0_u5_u4_n127 ) , .A( u0_u5_u4_n136 ) , .B2( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n180 ) );
  INV_X1 u0_u5_u4_U52 (.A( u0_u5_u4_n160 ) , .ZN( u0_u5_u4_n180 ) );
  NAND2_X1 u0_u5_u4_U53 (.A2( u0_u5_u4_n104 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n146 ) );
  NAND2_X1 u0_u5_u4_U54 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n160 ) );
  NAND2_X1 u0_u5_u4_U55 (.ZN( u0_u5_u4_n134 ) , .A1( u0_u5_u4_n98 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U56 (.A1( u0_u5_u4_n103 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n143 ) );
  NAND2_X1 u0_u5_u4_U57 (.A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U58 (.A1( u0_u5_u4_n100 ) , .A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n120 ) );
  NAND2_X1 u0_u5_u4_U59 (.A1( u0_u5_u4_n102 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n148 ) );
  AOI21_X1 u0_u5_u4_U6 (.ZN( u0_u5_u4_n106 ) , .B2( u0_u5_u4_n146 ) , .B1( u0_u5_u4_n158 ) , .A( u0_u5_u4_n170 ) );
  NAND2_X1 u0_u5_u4_U60 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n157 ) );
  INV_X1 u0_u5_u4_U61 (.A( u0_u5_u4_n150 ) , .ZN( u0_u5_u4_n173 ) );
  INV_X1 u0_u5_u4_U62 (.A( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n171 ) );
  NAND2_X1 u0_u5_u4_U63 (.A1( u0_u5_u4_n100 ) , .ZN( u0_u5_u4_n118 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U64 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n144 ) );
  NAND2_X1 u0_u5_u4_U65 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U66 (.A( u0_u5_u4_n128 ) , .ZN( u0_u5_u4_n174 ) );
  NAND2_X1 u0_u5_u4_U67 (.A2( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n119 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U68 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U69 (.A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n113 ) , .A1( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U7 (.ZN( u0_u5_u4_n108 ) , .B2( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n155 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U70 (.A2( u0_u5_X_28 ) , .ZN( u0_u5_u4_n150 ) , .A1( u0_u5_u4_n168 ) );
  NOR2_X1 u0_u5_u4_U71 (.A2( u0_u5_X_29 ) , .ZN( u0_u5_u4_n152 ) , .A1( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U72 (.A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n105 ) , .A1( u0_u5_u4_n176 ) );
  NOR2_X1 u0_u5_u4_U73 (.A2( u0_u5_X_26 ) , .ZN( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n177 ) );
  NOR2_X1 u0_u5_u4_U74 (.A2( u0_u5_X_28 ) , .A1( u0_u5_X_29 ) , .ZN( u0_u5_u4_n128 ) );
  NOR2_X1 u0_u5_u4_U75 (.A2( u0_u5_X_27 ) , .A1( u0_u5_X_30 ) , .ZN( u0_u5_u4_n102 ) );
  NOR2_X1 u0_u5_u4_U76 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n98 ) );
  AND2_X1 u0_u5_u4_U77 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n104 ) );
  AND2_X1 u0_u5_u4_U78 (.A1( u0_u5_X_30 ) , .A2( u0_u5_u4_n176 ) , .ZN( u0_u5_u4_n99 ) );
  AND2_X1 u0_u5_u4_U79 (.A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n101 ) , .A2( u0_u5_u4_n177 ) );
  AOI21_X1 u0_u5_u4_U8 (.ZN( u0_u5_u4_n109 ) , .A( u0_u5_u4_n153 ) , .B1( u0_u5_u4_n159 ) , .B2( u0_u5_u4_n184 ) );
  AND2_X1 u0_u5_u4_U80 (.A1( u0_u5_X_27 ) , .A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n103 ) );
  INV_X1 u0_u5_u4_U81 (.A( u0_u5_X_28 ) , .ZN( u0_u5_u4_n169 ) );
  INV_X1 u0_u5_u4_U82 (.A( u0_u5_X_29 ) , .ZN( u0_u5_u4_n168 ) );
  INV_X1 u0_u5_u4_U83 (.A( u0_u5_X_25 ) , .ZN( u0_u5_u4_n177 ) );
  INV_X1 u0_u5_u4_U84 (.A( u0_u5_X_27 ) , .ZN( u0_u5_u4_n176 ) );
  NAND4_X1 u0_u5_u4_U85 (.ZN( u0_out5_25 ) , .A4( u0_u5_u4_n139 ) , .A3( u0_u5_u4_n140 ) , .A2( u0_u5_u4_n141 ) , .A1( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U86 (.A( u0_u5_u4_n128 ) , .B2( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n130 ) , .ZN( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U87 (.B2( u0_u5_u4_n131 ) , .ZN( u0_u5_u4_n141 ) , .A( u0_u5_u4_n175 ) , .B1( u0_u5_u4_n183 ) );
  NAND4_X1 u0_u5_u4_U88 (.ZN( u0_out5_14 ) , .A4( u0_u5_u4_n124 ) , .A3( u0_u5_u4_n125 ) , .A2( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n127 ) );
  AOI22_X1 u0_u5_u4_U89 (.B2( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n152 ) , .A2( u0_u5_u4_n175 ) );
  AOI211_X1 u0_u5_u4_U9 (.B( u0_u5_u4_n136 ) , .A( u0_u5_u4_n137 ) , .C2( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n139 ) , .C1( u0_u5_u4_n182 ) );
  AOI22_X1 u0_u5_u4_U90 (.ZN( u0_u5_u4_n125 ) , .B2( u0_u5_u4_n131 ) , .A2( u0_u5_u4_n132 ) , .B1( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n178 ) );
  NAND4_X1 u0_u5_u4_U91 (.ZN( u0_out5_8 ) , .A4( u0_u5_u4_n110 ) , .A3( u0_u5_u4_n111 ) , .A2( u0_u5_u4_n112 ) , .A1( u0_u5_u4_n186 ) );
  NAND2_X1 u0_u5_u4_U92 (.ZN( u0_u5_u4_n112 ) , .A2( u0_u5_u4_n130 ) , .A1( u0_u5_u4_n150 ) );
  AOI22_X1 u0_u5_u4_U93 (.ZN( u0_u5_u4_n111 ) , .B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n152 ) , .B1( u0_u5_u4_n178 ) , .A2( u0_u5_u4_n97 ) );
  AOI22_X1 u0_u5_u4_U94 (.B2( u0_u5_u4_n149 ) , .B1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n151 ) , .A1( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n167 ) );
  NOR4_X1 u0_u5_u4_U95 (.A4( u0_u5_u4_n162 ) , .A3( u0_u5_u4_n163 ) , .A2( u0_u5_u4_n164 ) , .A1( u0_u5_u4_n165 ) , .ZN( u0_u5_u4_n166 ) );
  NAND3_X1 u0_u5_u4_U96 (.ZN( u0_out5_3 ) , .A3( u0_u5_u4_n166 ) , .A1( u0_u5_u4_n167 ) , .A2( u0_u5_u4_n186 ) );
  NAND3_X1 u0_u5_u4_U97 (.A3( u0_u5_u4_n146 ) , .A2( u0_u5_u4_n147 ) , .A1( u0_u5_u4_n148 ) , .ZN( u0_u5_u4_n149 ) );
  NAND3_X1 u0_u5_u4_U98 (.A3( u0_u5_u4_n143 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n145 ) , .ZN( u0_u5_u4_n151 ) );
  NAND3_X1 u0_u5_u4_U99 (.A3( u0_u5_u4_n121 ) , .ZN( u0_u5_u4_n122 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n154 ) );
  INV_X1 u0_u5_u5_U10 (.A( u0_u5_u5_n121 ) , .ZN( u0_u5_u5_n177 ) );
  NOR3_X1 u0_u5_u5_U100 (.A3( u0_u5_u5_n141 ) , .A1( u0_u5_u5_n142 ) , .ZN( u0_u5_u5_n143 ) , .A2( u0_u5_u5_n191 ) );
  NAND4_X1 u0_u5_u5_U101 (.ZN( u0_out5_4 ) , .A4( u0_u5_u5_n112 ) , .A2( u0_u5_u5_n113 ) , .A1( u0_u5_u5_n114 ) , .A3( u0_u5_u5_n195 ) );
  AOI211_X1 u0_u5_u5_U102 (.A( u0_u5_u5_n110 ) , .C1( u0_u5_u5_n111 ) , .ZN( u0_u5_u5_n112 ) , .B( u0_u5_u5_n118 ) , .C2( u0_u5_u5_n177 ) );
  AOI222_X1 u0_u5_u5_U103 (.ZN( u0_u5_u5_n113 ) , .A1( u0_u5_u5_n131 ) , .C1( u0_u5_u5_n148 ) , .B2( u0_u5_u5_n174 ) , .C2( u0_u5_u5_n178 ) , .A2( u0_u5_u5_n179 ) , .B1( u0_u5_u5_n99 ) );
  NAND3_X1 u0_u5_u5_U104 (.A2( u0_u5_u5_n154 ) , .A3( u0_u5_u5_n158 ) , .A1( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n99 ) );
  NOR2_X1 u0_u5_u5_U11 (.ZN( u0_u5_u5_n160 ) , .A2( u0_u5_u5_n173 ) , .A1( u0_u5_u5_n177 ) );
  INV_X1 u0_u5_u5_U12 (.A( u0_u5_u5_n150 ) , .ZN( u0_u5_u5_n174 ) );
  AOI21_X1 u0_u5_u5_U13 (.A( u0_u5_u5_n160 ) , .B2( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n162 ) , .B1( u0_u5_u5_n192 ) );
  INV_X1 u0_u5_u5_U14 (.A( u0_u5_u5_n159 ) , .ZN( u0_u5_u5_n192 ) );
  AOI21_X1 u0_u5_u5_U15 (.A( u0_u5_u5_n156 ) , .B2( u0_u5_u5_n157 ) , .B1( u0_u5_u5_n158 ) , .ZN( u0_u5_u5_n163 ) );
  AOI21_X1 u0_u5_u5_U16 (.B2( u0_u5_u5_n139 ) , .B1( u0_u5_u5_n140 ) , .ZN( u0_u5_u5_n141 ) , .A( u0_u5_u5_n150 ) );
  OAI21_X1 u0_u5_u5_U17 (.A( u0_u5_u5_n133 ) , .B2( u0_u5_u5_n134 ) , .B1( u0_u5_u5_n135 ) , .ZN( u0_u5_u5_n142 ) );
  OAI21_X1 u0_u5_u5_U18 (.ZN( u0_u5_u5_n133 ) , .B2( u0_u5_u5_n147 ) , .A( u0_u5_u5_n173 ) , .B1( u0_u5_u5_n188 ) );
  NAND2_X1 u0_u5_u5_U19 (.A2( u0_u5_u5_n119 ) , .A1( u0_u5_u5_n123 ) , .ZN( u0_u5_u5_n137 ) );
  INV_X1 u0_u5_u5_U20 (.A( u0_u5_u5_n155 ) , .ZN( u0_u5_u5_n194 ) );
  NAND2_X1 u0_u5_u5_U21 (.A1( u0_u5_u5_n121 ) , .ZN( u0_u5_u5_n132 ) , .A2( u0_u5_u5_n172 ) );
  NAND2_X1 u0_u5_u5_U22 (.A2( u0_u5_u5_n122 ) , .ZN( u0_u5_u5_n136 ) , .A1( u0_u5_u5_n154 ) );
  NAND2_X1 u0_u5_u5_U23 (.A2( u0_u5_u5_n119 ) , .A1( u0_u5_u5_n120 ) , .ZN( u0_u5_u5_n159 ) );
  INV_X1 u0_u5_u5_U24 (.A( u0_u5_u5_n156 ) , .ZN( u0_u5_u5_n175 ) );
  INV_X1 u0_u5_u5_U25 (.A( u0_u5_u5_n158 ) , .ZN( u0_u5_u5_n188 ) );
  INV_X1 u0_u5_u5_U26 (.A( u0_u5_u5_n152 ) , .ZN( u0_u5_u5_n179 ) );
  INV_X1 u0_u5_u5_U27 (.A( u0_u5_u5_n140 ) , .ZN( u0_u5_u5_n182 ) );
  INV_X1 u0_u5_u5_U28 (.A( u0_u5_u5_n151 ) , .ZN( u0_u5_u5_n183 ) );
  INV_X1 u0_u5_u5_U29 (.A( u0_u5_u5_n123 ) , .ZN( u0_u5_u5_n185 ) );
  NOR2_X1 u0_u5_u5_U3 (.ZN( u0_u5_u5_n134 ) , .A1( u0_u5_u5_n183 ) , .A2( u0_u5_u5_n190 ) );
  INV_X1 u0_u5_u5_U30 (.A( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n184 ) );
  INV_X1 u0_u5_u5_U31 (.A( u0_u5_u5_n139 ) , .ZN( u0_u5_u5_n189 ) );
  INV_X1 u0_u5_u5_U32 (.A( u0_u5_u5_n157 ) , .ZN( u0_u5_u5_n190 ) );
  INV_X1 u0_u5_u5_U33 (.A( u0_u5_u5_n120 ) , .ZN( u0_u5_u5_n193 ) );
  NAND2_X1 u0_u5_u5_U34 (.ZN( u0_u5_u5_n111 ) , .A1( u0_u5_u5_n140 ) , .A2( u0_u5_u5_n155 ) );
  NOR2_X1 u0_u5_u5_U35 (.ZN( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n170 ) , .A2( u0_u5_u5_n180 ) );
  INV_X1 u0_u5_u5_U36 (.A( u0_u5_u5_n117 ) , .ZN( u0_u5_u5_n196 ) );
  OAI221_X1 u0_u5_u5_U37 (.A( u0_u5_u5_n116 ) , .ZN( u0_u5_u5_n117 ) , .B2( u0_u5_u5_n119 ) , .C1( u0_u5_u5_n153 ) , .C2( u0_u5_u5_n158 ) , .B1( u0_u5_u5_n172 ) );
  AOI222_X1 u0_u5_u5_U38 (.ZN( u0_u5_u5_n116 ) , .B2( u0_u5_u5_n145 ) , .C1( u0_u5_u5_n148 ) , .A2( u0_u5_u5_n174 ) , .C2( u0_u5_u5_n177 ) , .B1( u0_u5_u5_n187 ) , .A1( u0_u5_u5_n193 ) );
  INV_X1 u0_u5_u5_U39 (.A( u0_u5_u5_n115 ) , .ZN( u0_u5_u5_n187 ) );
  INV_X1 u0_u5_u5_U4 (.A( u0_u5_u5_n138 ) , .ZN( u0_u5_u5_n191 ) );
  AOI22_X1 u0_u5_u5_U40 (.B2( u0_u5_u5_n131 ) , .A2( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n169 ) , .B1( u0_u5_u5_n174 ) , .A1( u0_u5_u5_n185 ) );
  NOR2_X1 u0_u5_u5_U41 (.A1( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n150 ) , .A2( u0_u5_u5_n173 ) );
  AOI21_X1 u0_u5_u5_U42 (.A( u0_u5_u5_n118 ) , .B2( u0_u5_u5_n145 ) , .ZN( u0_u5_u5_n168 ) , .B1( u0_u5_u5_n186 ) );
  INV_X1 u0_u5_u5_U43 (.A( u0_u5_u5_n122 ) , .ZN( u0_u5_u5_n186 ) );
  NOR2_X1 u0_u5_u5_U44 (.A1( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n152 ) , .A2( u0_u5_u5_n176 ) );
  NOR2_X1 u0_u5_u5_U45 (.A1( u0_u5_u5_n115 ) , .ZN( u0_u5_u5_n118 ) , .A2( u0_u5_u5_n153 ) );
  NOR2_X1 u0_u5_u5_U46 (.A2( u0_u5_u5_n145 ) , .ZN( u0_u5_u5_n156 ) , .A1( u0_u5_u5_n174 ) );
  NOR2_X1 u0_u5_u5_U47 (.ZN( u0_u5_u5_n121 ) , .A2( u0_u5_u5_n145 ) , .A1( u0_u5_u5_n176 ) );
  AOI22_X1 u0_u5_u5_U48 (.ZN( u0_u5_u5_n114 ) , .A2( u0_u5_u5_n137 ) , .A1( u0_u5_u5_n145 ) , .B2( u0_u5_u5_n175 ) , .B1( u0_u5_u5_n193 ) );
  OAI211_X1 u0_u5_u5_U49 (.B( u0_u5_u5_n124 ) , .A( u0_u5_u5_n125 ) , .C2( u0_u5_u5_n126 ) , .C1( u0_u5_u5_n127 ) , .ZN( u0_u5_u5_n128 ) );
  OAI21_X1 u0_u5_u5_U5 (.B2( u0_u5_u5_n136 ) , .B1( u0_u5_u5_n137 ) , .ZN( u0_u5_u5_n138 ) , .A( u0_u5_u5_n177 ) );
  NOR3_X1 u0_u5_u5_U50 (.ZN( u0_u5_u5_n127 ) , .A1( u0_u5_u5_n136 ) , .A3( u0_u5_u5_n148 ) , .A2( u0_u5_u5_n182 ) );
  OAI21_X1 u0_u5_u5_U51 (.ZN( u0_u5_u5_n124 ) , .A( u0_u5_u5_n177 ) , .B2( u0_u5_u5_n183 ) , .B1( u0_u5_u5_n189 ) );
  OAI21_X1 u0_u5_u5_U52 (.ZN( u0_u5_u5_n125 ) , .A( u0_u5_u5_n174 ) , .B2( u0_u5_u5_n185 ) , .B1( u0_u5_u5_n190 ) );
  AOI21_X1 u0_u5_u5_U53 (.A( u0_u5_u5_n153 ) , .B2( u0_u5_u5_n154 ) , .B1( u0_u5_u5_n155 ) , .ZN( u0_u5_u5_n164 ) );
  AOI21_X1 u0_u5_u5_U54 (.ZN( u0_u5_u5_n110 ) , .B1( u0_u5_u5_n122 ) , .B2( u0_u5_u5_n139 ) , .A( u0_u5_u5_n153 ) );
  INV_X1 u0_u5_u5_U55 (.A( u0_u5_u5_n153 ) , .ZN( u0_u5_u5_n176 ) );
  INV_X1 u0_u5_u5_U56 (.A( u0_u5_u5_n126 ) , .ZN( u0_u5_u5_n173 ) );
  AND2_X1 u0_u5_u5_U57 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n147 ) );
  AND2_X1 u0_u5_u5_U58 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n148 ) );
  NAND2_X1 u0_u5_u5_U59 (.A1( u0_u5_u5_n105 ) , .A2( u0_u5_u5_n106 ) , .ZN( u0_u5_u5_n158 ) );
  INV_X1 u0_u5_u5_U6 (.A( u0_u5_u5_n135 ) , .ZN( u0_u5_u5_n178 ) );
  NAND2_X1 u0_u5_u5_U60 (.A2( u0_u5_u5_n108 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n139 ) );
  NAND2_X1 u0_u5_u5_U61 (.A1( u0_u5_u5_n106 ) , .A2( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n119 ) );
  NAND2_X1 u0_u5_u5_U62 (.A2( u0_u5_u5_n103 ) , .A1( u0_u5_u5_n105 ) , .ZN( u0_u5_u5_n140 ) );
  NAND2_X1 u0_u5_u5_U63 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n105 ) , .ZN( u0_u5_u5_n155 ) );
  NAND2_X1 u0_u5_u5_U64 (.A2( u0_u5_u5_n106 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n122 ) );
  NAND2_X1 u0_u5_u5_U65 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n106 ) , .ZN( u0_u5_u5_n115 ) );
  NAND2_X1 u0_u5_u5_U66 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n103 ) , .ZN( u0_u5_u5_n161 ) );
  NAND2_X1 u0_u5_u5_U67 (.A1( u0_u5_u5_n105 ) , .A2( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n154 ) );
  INV_X1 u0_u5_u5_U68 (.A( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n172 ) );
  NAND2_X1 u0_u5_u5_U69 (.A1( u0_u5_u5_n103 ) , .A2( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n123 ) );
  OAI22_X1 u0_u5_u5_U7 (.B2( u0_u5_u5_n149 ) , .B1( u0_u5_u5_n150 ) , .A2( u0_u5_u5_n151 ) , .A1( u0_u5_u5_n152 ) , .ZN( u0_u5_u5_n165 ) );
  NAND2_X1 u0_u5_u5_U70 (.A2( u0_u5_u5_n103 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n151 ) );
  NAND2_X1 u0_u5_u5_U71 (.A2( u0_u5_u5_n107 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n120 ) );
  NAND2_X1 u0_u5_u5_U72 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n157 ) );
  AND2_X1 u0_u5_u5_U73 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n104 ) , .ZN( u0_u5_u5_n131 ) );
  INV_X1 u0_u5_u5_U74 (.A( u0_u5_u5_n102 ) , .ZN( u0_u5_u5_n195 ) );
  OAI221_X1 u0_u5_u5_U75 (.A( u0_u5_u5_n101 ) , .ZN( u0_u5_u5_n102 ) , .C2( u0_u5_u5_n115 ) , .C1( u0_u5_u5_n126 ) , .B1( u0_u5_u5_n134 ) , .B2( u0_u5_u5_n160 ) );
  OAI21_X1 u0_u5_u5_U76 (.ZN( u0_u5_u5_n101 ) , .B1( u0_u5_u5_n137 ) , .A( u0_u5_u5_n146 ) , .B2( u0_u5_u5_n147 ) );
  NOR2_X1 u0_u5_u5_U77 (.A2( u0_u5_X_34 ) , .A1( u0_u5_X_35 ) , .ZN( u0_u5_u5_n145 ) );
  NOR2_X1 u0_u5_u5_U78 (.A2( u0_u5_X_34 ) , .ZN( u0_u5_u5_n146 ) , .A1( u0_u5_u5_n171 ) );
  NOR2_X1 u0_u5_u5_U79 (.A2( u0_u5_X_31 ) , .A1( u0_u5_X_32 ) , .ZN( u0_u5_u5_n103 ) );
  NOR3_X1 u0_u5_u5_U8 (.A2( u0_u5_u5_n147 ) , .A1( u0_u5_u5_n148 ) , .ZN( u0_u5_u5_n149 ) , .A3( u0_u5_u5_n194 ) );
  NOR2_X1 u0_u5_u5_U80 (.A2( u0_u5_X_36 ) , .ZN( u0_u5_u5_n105 ) , .A1( u0_u5_u5_n180 ) );
  NOR2_X1 u0_u5_u5_U81 (.A2( u0_u5_X_33 ) , .ZN( u0_u5_u5_n108 ) , .A1( u0_u5_u5_n170 ) );
  NOR2_X1 u0_u5_u5_U82 (.A2( u0_u5_X_33 ) , .A1( u0_u5_X_36 ) , .ZN( u0_u5_u5_n107 ) );
  NOR2_X1 u0_u5_u5_U83 (.A2( u0_u5_X_31 ) , .ZN( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n181 ) );
  NAND2_X1 u0_u5_u5_U84 (.A2( u0_u5_X_34 ) , .A1( u0_u5_X_35 ) , .ZN( u0_u5_u5_n153 ) );
  NAND2_X1 u0_u5_u5_U85 (.A1( u0_u5_X_34 ) , .ZN( u0_u5_u5_n126 ) , .A2( u0_u5_u5_n171 ) );
  AND2_X1 u0_u5_u5_U86 (.A1( u0_u5_X_31 ) , .A2( u0_u5_X_32 ) , .ZN( u0_u5_u5_n106 ) );
  AND2_X1 u0_u5_u5_U87 (.A1( u0_u5_X_31 ) , .ZN( u0_u5_u5_n109 ) , .A2( u0_u5_u5_n181 ) );
  INV_X1 u0_u5_u5_U88 (.A( u0_u5_X_33 ) , .ZN( u0_u5_u5_n180 ) );
  INV_X1 u0_u5_u5_U89 (.A( u0_u5_X_35 ) , .ZN( u0_u5_u5_n171 ) );
  NOR2_X1 u0_u5_u5_U9 (.ZN( u0_u5_u5_n135 ) , .A1( u0_u5_u5_n173 ) , .A2( u0_u5_u5_n176 ) );
  INV_X1 u0_u5_u5_U90 (.A( u0_u5_X_36 ) , .ZN( u0_u5_u5_n170 ) );
  INV_X1 u0_u5_u5_U91 (.A( u0_u5_X_32 ) , .ZN( u0_u5_u5_n181 ) );
  NAND4_X1 u0_u5_u5_U92 (.ZN( u0_out5_29 ) , .A4( u0_u5_u5_n129 ) , .A3( u0_u5_u5_n130 ) , .A2( u0_u5_u5_n168 ) , .A1( u0_u5_u5_n196 ) );
  AOI221_X1 u0_u5_u5_U93 (.A( u0_u5_u5_n128 ) , .ZN( u0_u5_u5_n129 ) , .C2( u0_u5_u5_n132 ) , .B2( u0_u5_u5_n159 ) , .B1( u0_u5_u5_n176 ) , .C1( u0_u5_u5_n184 ) );
  AOI222_X1 u0_u5_u5_U94 (.ZN( u0_u5_u5_n130 ) , .A2( u0_u5_u5_n146 ) , .B1( u0_u5_u5_n147 ) , .C2( u0_u5_u5_n175 ) , .B2( u0_u5_u5_n179 ) , .A1( u0_u5_u5_n188 ) , .C1( u0_u5_u5_n194 ) );
  NAND4_X1 u0_u5_u5_U95 (.ZN( u0_out5_19 ) , .A4( u0_u5_u5_n166 ) , .A3( u0_u5_u5_n167 ) , .A2( u0_u5_u5_n168 ) , .A1( u0_u5_u5_n169 ) );
  AOI22_X1 u0_u5_u5_U96 (.B2( u0_u5_u5_n145 ) , .A2( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n167 ) , .B1( u0_u5_u5_n182 ) , .A1( u0_u5_u5_n189 ) );
  NOR4_X1 u0_u5_u5_U97 (.A4( u0_u5_u5_n162 ) , .A3( u0_u5_u5_n163 ) , .A2( u0_u5_u5_n164 ) , .A1( u0_u5_u5_n165 ) , .ZN( u0_u5_u5_n166 ) );
  NAND4_X1 u0_u5_u5_U98 (.ZN( u0_out5_11 ) , .A4( u0_u5_u5_n143 ) , .A3( u0_u5_u5_n144 ) , .A2( u0_u5_u5_n169 ) , .A1( u0_u5_u5_n196 ) );
  AOI22_X1 u0_u5_u5_U99 (.A2( u0_u5_u5_n132 ) , .ZN( u0_u5_u5_n144 ) , .B2( u0_u5_u5_n145 ) , .B1( u0_u5_u5_n184 ) , .A1( u0_u5_u5_n194 ) );
  OAI21_X1 u0_u5_u6_U10 (.A( u0_u5_u6_n159 ) , .B1( u0_u5_u6_n169 ) , .B2( u0_u5_u6_n173 ) , .ZN( u0_u5_u6_n90 ) );
  INV_X1 u0_u5_u6_U11 (.ZN( u0_u5_u6_n172 ) , .A( u0_u5_u6_n88 ) );
  AOI22_X1 u0_u5_u6_U12 (.A2( u0_u5_u6_n151 ) , .B2( u0_u5_u6_n161 ) , .A1( u0_u5_u6_n167 ) , .B1( u0_u5_u6_n170 ) , .ZN( u0_u5_u6_n89 ) );
  AOI21_X1 u0_u5_u6_U13 (.ZN( u0_u5_u6_n106 ) , .A( u0_u5_u6_n142 ) , .B2( u0_u5_u6_n159 ) , .B1( u0_u5_u6_n164 ) );
  INV_X1 u0_u5_u6_U14 (.A( u0_u5_u6_n155 ) , .ZN( u0_u5_u6_n161 ) );
  INV_X1 u0_u5_u6_U15 (.A( u0_u5_u6_n128 ) , .ZN( u0_u5_u6_n164 ) );
  NAND2_X1 u0_u5_u6_U16 (.ZN( u0_u5_u6_n110 ) , .A1( u0_u5_u6_n122 ) , .A2( u0_u5_u6_n129 ) );
  NAND2_X1 u0_u5_u6_U17 (.ZN( u0_u5_u6_n124 ) , .A2( u0_u5_u6_n146 ) , .A1( u0_u5_u6_n148 ) );
  INV_X1 u0_u5_u6_U18 (.A( u0_u5_u6_n132 ) , .ZN( u0_u5_u6_n171 ) );
  AND2_X1 u0_u5_u6_U19 (.A1( u0_u5_u6_n100 ) , .ZN( u0_u5_u6_n130 ) , .A2( u0_u5_u6_n147 ) );
  INV_X1 u0_u5_u6_U20 (.A( u0_u5_u6_n127 ) , .ZN( u0_u5_u6_n173 ) );
  INV_X1 u0_u5_u6_U21 (.A( u0_u5_u6_n121 ) , .ZN( u0_u5_u6_n167 ) );
  INV_X1 u0_u5_u6_U22 (.A( u0_u5_u6_n100 ) , .ZN( u0_u5_u6_n169 ) );
  INV_X1 u0_u5_u6_U23 (.A( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n170 ) );
  INV_X1 u0_u5_u6_U24 (.A( u0_u5_u6_n113 ) , .ZN( u0_u5_u6_n168 ) );
  AND2_X1 u0_u5_u6_U25 (.A1( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n119 ) , .ZN( u0_u5_u6_n133 ) );
  AND2_X1 u0_u5_u6_U26 (.A2( u0_u5_u6_n121 ) , .A1( u0_u5_u6_n122 ) , .ZN( u0_u5_u6_n131 ) );
  AND3_X1 u0_u5_u6_U27 (.ZN( u0_u5_u6_n120 ) , .A2( u0_u5_u6_n127 ) , .A1( u0_u5_u6_n132 ) , .A3( u0_u5_u6_n145 ) );
  INV_X1 u0_u5_u6_U28 (.A( u0_u5_u6_n146 ) , .ZN( u0_u5_u6_n163 ) );
  AOI222_X1 u0_u5_u6_U29 (.ZN( u0_u5_u6_n114 ) , .A1( u0_u5_u6_n118 ) , .A2( u0_u5_u6_n126 ) , .B2( u0_u5_u6_n151 ) , .C2( u0_u5_u6_n159 ) , .C1( u0_u5_u6_n168 ) , .B1( u0_u5_u6_n169 ) );
  INV_X1 u0_u5_u6_U3 (.A( u0_u5_u6_n110 ) , .ZN( u0_u5_u6_n166 ) );
  NOR2_X1 u0_u5_u6_U30 (.A1( u0_u5_u6_n162 ) , .A2( u0_u5_u6_n165 ) , .ZN( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U31 (.A1( u0_u5_u6_n144 ) , .ZN( u0_u5_u6_n151 ) , .A2( u0_u5_u6_n158 ) );
  NAND2_X1 u0_u5_u6_U32 (.ZN( u0_u5_u6_n132 ) , .A1( u0_u5_u6_n91 ) , .A2( u0_u5_u6_n97 ) );
  NOR2_X1 u0_u5_u6_U33 (.A2( u0_u5_u6_n126 ) , .ZN( u0_u5_u6_n155 ) , .A1( u0_u5_u6_n160 ) );
  NAND2_X1 u0_u5_u6_U34 (.ZN( u0_u5_u6_n146 ) , .A2( u0_u5_u6_n94 ) , .A1( u0_u5_u6_n99 ) );
  AOI21_X1 u0_u5_u6_U35 (.A( u0_u5_u6_n144 ) , .B2( u0_u5_u6_n145 ) , .B1( u0_u5_u6_n146 ) , .ZN( u0_u5_u6_n150 ) );
  INV_X1 u0_u5_u6_U36 (.A( u0_u5_u6_n111 ) , .ZN( u0_u5_u6_n158 ) );
  NAND2_X1 u0_u5_u6_U37 (.ZN( u0_u5_u6_n127 ) , .A1( u0_u5_u6_n91 ) , .A2( u0_u5_u6_n92 ) );
  NAND2_X1 u0_u5_u6_U38 (.ZN( u0_u5_u6_n129 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n96 ) );
  INV_X1 u0_u5_u6_U39 (.A( u0_u5_u6_n144 ) , .ZN( u0_u5_u6_n159 ) );
  INV_X1 u0_u5_u6_U4 (.A( u0_u5_u6_n142 ) , .ZN( u0_u5_u6_n174 ) );
  NAND2_X1 u0_u5_u6_U40 (.ZN( u0_u5_u6_n145 ) , .A2( u0_u5_u6_n97 ) , .A1( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U41 (.ZN( u0_u5_u6_n148 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n94 ) );
  NAND2_X1 u0_u5_u6_U42 (.ZN( u0_u5_u6_n108 ) , .A2( u0_u5_u6_n139 ) , .A1( u0_u5_u6_n144 ) );
  NAND2_X1 u0_u5_u6_U43 (.ZN( u0_u5_u6_n121 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n97 ) );
  NAND2_X1 u0_u5_u6_U44 (.ZN( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n95 ) );
  AND2_X1 u0_u5_u6_U45 (.ZN( u0_u5_u6_n118 ) , .A2( u0_u5_u6_n91 ) , .A1( u0_u5_u6_n99 ) );
  AOI22_X1 u0_u5_u6_U46 (.B2( u0_u5_u6_n110 ) , .B1( u0_u5_u6_n111 ) , .A1( u0_u5_u6_n112 ) , .ZN( u0_u5_u6_n115 ) , .A2( u0_u5_u6_n161 ) );
  NAND4_X1 u0_u5_u6_U47 (.A3( u0_u5_u6_n109 ) , .ZN( u0_u5_u6_n112 ) , .A4( u0_u5_u6_n132 ) , .A2( u0_u5_u6_n147 ) , .A1( u0_u5_u6_n166 ) );
  NOR2_X1 u0_u5_u6_U48 (.ZN( u0_u5_u6_n109 ) , .A1( u0_u5_u6_n170 ) , .A2( u0_u5_u6_n173 ) );
  NAND2_X1 u0_u5_u6_U49 (.ZN( u0_u5_u6_n147 ) , .A2( u0_u5_u6_n98 ) , .A1( u0_u5_u6_n99 ) );
  NAND2_X1 u0_u5_u6_U5 (.A2( u0_u5_u6_n143 ) , .ZN( u0_u5_u6_n152 ) , .A1( u0_u5_u6_n166 ) );
  NAND2_X1 u0_u5_u6_U50 (.ZN( u0_u5_u6_n128 ) , .A1( u0_u5_u6_n94 ) , .A2( u0_u5_u6_n96 ) );
  AOI211_X1 u0_u5_u6_U51 (.B( u0_u5_u6_n134 ) , .A( u0_u5_u6_n135 ) , .C1( u0_u5_u6_n136 ) , .ZN( u0_u5_u6_n137 ) , .C2( u0_u5_u6_n151 ) );
  AOI21_X1 u0_u5_u6_U52 (.B2( u0_u5_u6_n132 ) , .B1( u0_u5_u6_n133 ) , .ZN( u0_u5_u6_n134 ) , .A( u0_u5_u6_n158 ) );
  AOI21_X1 u0_u5_u6_U53 (.B1( u0_u5_u6_n131 ) , .ZN( u0_u5_u6_n135 ) , .A( u0_u5_u6_n144 ) , .B2( u0_u5_u6_n146 ) );
  NAND4_X1 u0_u5_u6_U54 (.A4( u0_u5_u6_n127 ) , .A3( u0_u5_u6_n128 ) , .A2( u0_u5_u6_n129 ) , .A1( u0_u5_u6_n130 ) , .ZN( u0_u5_u6_n136 ) );
  NAND2_X1 u0_u5_u6_U55 (.ZN( u0_u5_u6_n119 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n99 ) );
  NAND2_X1 u0_u5_u6_U56 (.ZN( u0_u5_u6_n123 ) , .A2( u0_u5_u6_n91 ) , .A1( u0_u5_u6_n96 ) );
  NAND2_X1 u0_u5_u6_U57 (.ZN( u0_u5_u6_n100 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U58 (.ZN( u0_u5_u6_n122 ) , .A1( u0_u5_u6_n94 ) , .A2( u0_u5_u6_n97 ) );
  INV_X1 u0_u5_u6_U59 (.A( u0_u5_u6_n139 ) , .ZN( u0_u5_u6_n160 ) );
  AOI22_X1 u0_u5_u6_U6 (.B2( u0_u5_u6_n101 ) , .A1( u0_u5_u6_n102 ) , .ZN( u0_u5_u6_n103 ) , .B1( u0_u5_u6_n160 ) , .A2( u0_u5_u6_n161 ) );
  NAND2_X1 u0_u5_u6_U60 (.ZN( u0_u5_u6_n113 ) , .A1( u0_u5_u6_n96 ) , .A2( u0_u5_u6_n98 ) );
  NOR2_X1 u0_u5_u6_U61 (.A2( u0_u5_X_40 ) , .A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n126 ) );
  NOR2_X1 u0_u5_u6_U62 (.A2( u0_u5_X_39 ) , .A1( u0_u5_X_42 ) , .ZN( u0_u5_u6_n92 ) );
  NOR2_X1 u0_u5_u6_U63 (.A2( u0_u5_X_39 ) , .A1( u0_u5_u6_n156 ) , .ZN( u0_u5_u6_n97 ) );
  NOR2_X1 u0_u5_u6_U64 (.A2( u0_u5_X_38 ) , .A1( u0_u5_u6_n165 ) , .ZN( u0_u5_u6_n95 ) );
  NOR2_X1 u0_u5_u6_U65 (.A2( u0_u5_X_41 ) , .ZN( u0_u5_u6_n111 ) , .A1( u0_u5_u6_n157 ) );
  NOR2_X1 u0_u5_u6_U66 (.A2( u0_u5_X_37 ) , .A1( u0_u5_u6_n162 ) , .ZN( u0_u5_u6_n94 ) );
  NOR2_X1 u0_u5_u6_U67 (.A2( u0_u5_X_37 ) , .A1( u0_u5_X_38 ) , .ZN( u0_u5_u6_n91 ) );
  NAND2_X1 u0_u5_u6_U68 (.A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n144 ) , .A2( u0_u5_u6_n157 ) );
  NAND2_X1 u0_u5_u6_U69 (.A2( u0_u5_X_40 ) , .A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n139 ) );
  NOR2_X1 u0_u5_u6_U7 (.A1( u0_u5_u6_n118 ) , .ZN( u0_u5_u6_n143 ) , .A2( u0_u5_u6_n168 ) );
  AND2_X1 u0_u5_u6_U70 (.A1( u0_u5_X_39 ) , .A2( u0_u5_u6_n156 ) , .ZN( u0_u5_u6_n96 ) );
  AND2_X1 u0_u5_u6_U71 (.A1( u0_u5_X_39 ) , .A2( u0_u5_X_42 ) , .ZN( u0_u5_u6_n99 ) );
  INV_X1 u0_u5_u6_U72 (.A( u0_u5_X_40 ) , .ZN( u0_u5_u6_n157 ) );
  INV_X1 u0_u5_u6_U73 (.A( u0_u5_X_37 ) , .ZN( u0_u5_u6_n165 ) );
  INV_X1 u0_u5_u6_U74 (.A( u0_u5_X_38 ) , .ZN( u0_u5_u6_n162 ) );
  INV_X1 u0_u5_u6_U75 (.A( u0_u5_X_42 ) , .ZN( u0_u5_u6_n156 ) );
  NAND4_X1 u0_u5_u6_U76 (.ZN( u0_out5_32 ) , .A4( u0_u5_u6_n103 ) , .A3( u0_u5_u6_n104 ) , .A2( u0_u5_u6_n105 ) , .A1( u0_u5_u6_n106 ) );
  AOI22_X1 u0_u5_u6_U77 (.ZN( u0_u5_u6_n105 ) , .A2( u0_u5_u6_n108 ) , .A1( u0_u5_u6_n118 ) , .B2( u0_u5_u6_n126 ) , .B1( u0_u5_u6_n171 ) );
  AOI22_X1 u0_u5_u6_U78 (.ZN( u0_u5_u6_n104 ) , .A1( u0_u5_u6_n111 ) , .B1( u0_u5_u6_n124 ) , .B2( u0_u5_u6_n151 ) , .A2( u0_u5_u6_n93 ) );
  NAND4_X1 u0_u5_u6_U79 (.ZN( u0_out5_12 ) , .A4( u0_u5_u6_n114 ) , .A3( u0_u5_u6_n115 ) , .A2( u0_u5_u6_n116 ) , .A1( u0_u5_u6_n117 ) );
  AOI21_X1 u0_u5_u6_U8 (.B1( u0_u5_u6_n107 ) , .B2( u0_u5_u6_n132 ) , .A( u0_u5_u6_n158 ) , .ZN( u0_u5_u6_n88 ) );
  OAI22_X1 u0_u5_u6_U80 (.B2( u0_u5_u6_n111 ) , .ZN( u0_u5_u6_n116 ) , .B1( u0_u5_u6_n126 ) , .A2( u0_u5_u6_n164 ) , .A1( u0_u5_u6_n167 ) );
  OAI21_X1 u0_u5_u6_U81 (.A( u0_u5_u6_n108 ) , .ZN( u0_u5_u6_n117 ) , .B2( u0_u5_u6_n141 ) , .B1( u0_u5_u6_n163 ) );
  OAI211_X1 u0_u5_u6_U82 (.ZN( u0_out5_22 ) , .B( u0_u5_u6_n137 ) , .A( u0_u5_u6_n138 ) , .C2( u0_u5_u6_n139 ) , .C1( u0_u5_u6_n140 ) );
  AOI22_X1 u0_u5_u6_U83 (.B1( u0_u5_u6_n124 ) , .A2( u0_u5_u6_n125 ) , .A1( u0_u5_u6_n126 ) , .ZN( u0_u5_u6_n138 ) , .B2( u0_u5_u6_n161 ) );
  AND4_X1 u0_u5_u6_U84 (.A3( u0_u5_u6_n119 ) , .A1( u0_u5_u6_n120 ) , .A4( u0_u5_u6_n129 ) , .ZN( u0_u5_u6_n140 ) , .A2( u0_u5_u6_n143 ) );
  OAI211_X1 u0_u5_u6_U85 (.ZN( u0_out5_7 ) , .B( u0_u5_u6_n153 ) , .C2( u0_u5_u6_n154 ) , .C1( u0_u5_u6_n155 ) , .A( u0_u5_u6_n174 ) );
  NOR3_X1 u0_u5_u6_U86 (.A1( u0_u5_u6_n141 ) , .ZN( u0_u5_u6_n154 ) , .A3( u0_u5_u6_n164 ) , .A2( u0_u5_u6_n171 ) );
  AOI211_X1 u0_u5_u6_U87 (.B( u0_u5_u6_n149 ) , .A( u0_u5_u6_n150 ) , .C2( u0_u5_u6_n151 ) , .C1( u0_u5_u6_n152 ) , .ZN( u0_u5_u6_n153 ) );
  NAND3_X1 u0_u5_u6_U88 (.A2( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n125 ) , .A1( u0_u5_u6_n130 ) , .A3( u0_u5_u6_n131 ) );
  NAND3_X1 u0_u5_u6_U89 (.A3( u0_u5_u6_n133 ) , .ZN( u0_u5_u6_n141 ) , .A1( u0_u5_u6_n145 ) , .A2( u0_u5_u6_n148 ) );
  AOI21_X1 u0_u5_u6_U9 (.B2( u0_u5_u6_n147 ) , .B1( u0_u5_u6_n148 ) , .ZN( u0_u5_u6_n149 ) , .A( u0_u5_u6_n158 ) );
  NAND3_X1 u0_u5_u6_U90 (.ZN( u0_u5_u6_n101 ) , .A3( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n121 ) , .A1( u0_u5_u6_n127 ) );
  NAND3_X1 u0_u5_u6_U91 (.ZN( u0_u5_u6_n102 ) , .A3( u0_u5_u6_n130 ) , .A2( u0_u5_u6_n145 ) , .A1( u0_u5_u6_n166 ) );
  NAND3_X1 u0_u5_u6_U92 (.A3( u0_u5_u6_n113 ) , .A1( u0_u5_u6_n119 ) , .A2( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n93 ) );
  NAND3_X1 u0_u5_u6_U93 (.ZN( u0_u5_u6_n142 ) , .A2( u0_u5_u6_n172 ) , .A3( u0_u5_u6_n89 ) , .A1( u0_u5_u6_n90 ) );
  AND3_X1 u0_u5_u7_U10 (.A3( u0_u5_u7_n110 ) , .A2( u0_u5_u7_n127 ) , .A1( u0_u5_u7_n132 ) , .ZN( u0_u5_u7_n92 ) );
  OAI21_X1 u0_u5_u7_U11 (.A( u0_u5_u7_n161 ) , .B1( u0_u5_u7_n168 ) , .B2( u0_u5_u7_n173 ) , .ZN( u0_u5_u7_n91 ) );
  AOI211_X1 u0_u5_u7_U12 (.A( u0_u5_u7_n117 ) , .ZN( u0_u5_u7_n118 ) , .C2( u0_u5_u7_n126 ) , .C1( u0_u5_u7_n177 ) , .B( u0_u5_u7_n180 ) );
  OAI22_X1 u0_u5_u7_U13 (.B1( u0_u5_u7_n115 ) , .ZN( u0_u5_u7_n117 ) , .A2( u0_u5_u7_n133 ) , .A1( u0_u5_u7_n137 ) , .B2( u0_u5_u7_n162 ) );
  INV_X1 u0_u5_u7_U14 (.A( u0_u5_u7_n116 ) , .ZN( u0_u5_u7_n180 ) );
  NOR3_X1 u0_u5_u7_U15 (.ZN( u0_u5_u7_n115 ) , .A3( u0_u5_u7_n145 ) , .A2( u0_u5_u7_n168 ) , .A1( u0_u5_u7_n169 ) );
  OAI211_X1 u0_u5_u7_U16 (.B( u0_u5_u7_n122 ) , .A( u0_u5_u7_n123 ) , .C2( u0_u5_u7_n124 ) , .ZN( u0_u5_u7_n154 ) , .C1( u0_u5_u7_n162 ) );
  AOI222_X1 u0_u5_u7_U17 (.ZN( u0_u5_u7_n122 ) , .C2( u0_u5_u7_n126 ) , .C1( u0_u5_u7_n145 ) , .B1( u0_u5_u7_n161 ) , .A2( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n170 ) , .A1( u0_u5_u7_n176 ) );
  INV_X1 u0_u5_u7_U18 (.A( u0_u5_u7_n133 ) , .ZN( u0_u5_u7_n176 ) );
  NOR3_X1 u0_u5_u7_U19 (.A2( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n135 ) , .ZN( u0_u5_u7_n136 ) , .A3( u0_u5_u7_n171 ) );
  NOR2_X1 u0_u5_u7_U20 (.A1( u0_u5_u7_n130 ) , .A2( u0_u5_u7_n134 ) , .ZN( u0_u5_u7_n153 ) );
  INV_X1 u0_u5_u7_U21 (.A( u0_u5_u7_n101 ) , .ZN( u0_u5_u7_n165 ) );
  NOR2_X1 u0_u5_u7_U22 (.ZN( u0_u5_u7_n111 ) , .A2( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n169 ) );
  AOI21_X1 u0_u5_u7_U23 (.ZN( u0_u5_u7_n104 ) , .B2( u0_u5_u7_n112 ) , .B1( u0_u5_u7_n127 ) , .A( u0_u5_u7_n164 ) );
  AOI21_X1 u0_u5_u7_U24 (.ZN( u0_u5_u7_n106 ) , .B1( u0_u5_u7_n133 ) , .B2( u0_u5_u7_n146 ) , .A( u0_u5_u7_n162 ) );
  AOI21_X1 u0_u5_u7_U25 (.A( u0_u5_u7_n101 ) , .ZN( u0_u5_u7_n107 ) , .B2( u0_u5_u7_n128 ) , .B1( u0_u5_u7_n175 ) );
  INV_X1 u0_u5_u7_U26 (.A( u0_u5_u7_n138 ) , .ZN( u0_u5_u7_n171 ) );
  INV_X1 u0_u5_u7_U27 (.A( u0_u5_u7_n131 ) , .ZN( u0_u5_u7_n177 ) );
  INV_X1 u0_u5_u7_U28 (.A( u0_u5_u7_n110 ) , .ZN( u0_u5_u7_n174 ) );
  NAND2_X1 u0_u5_u7_U29 (.A1( u0_u5_u7_n129 ) , .A2( u0_u5_u7_n132 ) , .ZN( u0_u5_u7_n149 ) );
  OAI21_X1 u0_u5_u7_U3 (.ZN( u0_u5_u7_n159 ) , .A( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n171 ) , .B1( u0_u5_u7_n174 ) );
  NAND2_X1 u0_u5_u7_U30 (.A1( u0_u5_u7_n113 ) , .A2( u0_u5_u7_n124 ) , .ZN( u0_u5_u7_n130 ) );
  INV_X1 u0_u5_u7_U31 (.A( u0_u5_u7_n112 ) , .ZN( u0_u5_u7_n173 ) );
  INV_X1 u0_u5_u7_U32 (.A( u0_u5_u7_n128 ) , .ZN( u0_u5_u7_n168 ) );
  INV_X1 u0_u5_u7_U33 (.A( u0_u5_u7_n148 ) , .ZN( u0_u5_u7_n169 ) );
  INV_X1 u0_u5_u7_U34 (.A( u0_u5_u7_n127 ) , .ZN( u0_u5_u7_n179 ) );
  NOR2_X1 u0_u5_u7_U35 (.ZN( u0_u5_u7_n101 ) , .A2( u0_u5_u7_n150 ) , .A1( u0_u5_u7_n156 ) );
  AOI211_X1 u0_u5_u7_U36 (.B( u0_u5_u7_n154 ) , .A( u0_u5_u7_n155 ) , .C1( u0_u5_u7_n156 ) , .ZN( u0_u5_u7_n157 ) , .C2( u0_u5_u7_n172 ) );
  INV_X1 u0_u5_u7_U37 (.A( u0_u5_u7_n153 ) , .ZN( u0_u5_u7_n172 ) );
  AOI211_X1 u0_u5_u7_U38 (.B( u0_u5_u7_n139 ) , .A( u0_u5_u7_n140 ) , .C2( u0_u5_u7_n141 ) , .ZN( u0_u5_u7_n142 ) , .C1( u0_u5_u7_n156 ) );
  NAND4_X1 u0_u5_u7_U39 (.A3( u0_u5_u7_n127 ) , .A2( u0_u5_u7_n128 ) , .A1( u0_u5_u7_n129 ) , .ZN( u0_u5_u7_n141 ) , .A4( u0_u5_u7_n147 ) );
  INV_X1 u0_u5_u7_U4 (.A( u0_u5_u7_n111 ) , .ZN( u0_u5_u7_n170 ) );
  AOI21_X1 u0_u5_u7_U40 (.A( u0_u5_u7_n137 ) , .B1( u0_u5_u7_n138 ) , .ZN( u0_u5_u7_n139 ) , .B2( u0_u5_u7_n146 ) );
  OAI22_X1 u0_u5_u7_U41 (.B1( u0_u5_u7_n136 ) , .ZN( u0_u5_u7_n140 ) , .A1( u0_u5_u7_n153 ) , .B2( u0_u5_u7_n162 ) , .A2( u0_u5_u7_n164 ) );
  AOI21_X1 u0_u5_u7_U42 (.ZN( u0_u5_u7_n123 ) , .B1( u0_u5_u7_n165 ) , .B2( u0_u5_u7_n177 ) , .A( u0_u5_u7_n97 ) );
  AOI21_X1 u0_u5_u7_U43 (.B2( u0_u5_u7_n113 ) , .B1( u0_u5_u7_n124 ) , .A( u0_u5_u7_n125 ) , .ZN( u0_u5_u7_n97 ) );
  INV_X1 u0_u5_u7_U44 (.A( u0_u5_u7_n125 ) , .ZN( u0_u5_u7_n161 ) );
  INV_X1 u0_u5_u7_U45 (.A( u0_u5_u7_n152 ) , .ZN( u0_u5_u7_n162 ) );
  AOI22_X1 u0_u5_u7_U46 (.A2( u0_u5_u7_n114 ) , .ZN( u0_u5_u7_n119 ) , .B1( u0_u5_u7_n130 ) , .A1( u0_u5_u7_n156 ) , .B2( u0_u5_u7_n165 ) );
  NAND2_X1 u0_u5_u7_U47 (.A2( u0_u5_u7_n112 ) , .ZN( u0_u5_u7_n114 ) , .A1( u0_u5_u7_n175 ) );
  AND2_X1 u0_u5_u7_U48 (.ZN( u0_u5_u7_n145 ) , .A2( u0_u5_u7_n98 ) , .A1( u0_u5_u7_n99 ) );
  NOR2_X1 u0_u5_u7_U49 (.ZN( u0_u5_u7_n137 ) , .A1( u0_u5_u7_n150 ) , .A2( u0_u5_u7_n161 ) );
  INV_X1 u0_u5_u7_U5 (.A( u0_u5_u7_n149 ) , .ZN( u0_u5_u7_n175 ) );
  AOI21_X1 u0_u5_u7_U50 (.ZN( u0_u5_u7_n105 ) , .B2( u0_u5_u7_n110 ) , .A( u0_u5_u7_n125 ) , .B1( u0_u5_u7_n147 ) );
  NAND2_X1 u0_u5_u7_U51 (.ZN( u0_u5_u7_n146 ) , .A1( u0_u5_u7_n95 ) , .A2( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U52 (.A2( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n147 ) , .A1( u0_u5_u7_n93 ) );
  NAND2_X1 u0_u5_u7_U53 (.A1( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n127 ) , .A2( u0_u5_u7_n99 ) );
  OR2_X1 u0_u5_u7_U54 (.ZN( u0_u5_u7_n126 ) , .A2( u0_u5_u7_n152 ) , .A1( u0_u5_u7_n156 ) );
  NAND2_X1 u0_u5_u7_U55 (.A2( u0_u5_u7_n102 ) , .A1( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n133 ) );
  NAND2_X1 u0_u5_u7_U56 (.ZN( u0_u5_u7_n112 ) , .A2( u0_u5_u7_n96 ) , .A1( u0_u5_u7_n99 ) );
  NAND2_X1 u0_u5_u7_U57 (.A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n128 ) , .A1( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U58 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n113 ) , .A2( u0_u5_u7_n93 ) );
  NAND2_X1 u0_u5_u7_U59 (.A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n124 ) , .A1( u0_u5_u7_n96 ) );
  INV_X1 u0_u5_u7_U6 (.A( u0_u5_u7_n154 ) , .ZN( u0_u5_u7_n178 ) );
  NAND2_X1 u0_u5_u7_U60 (.ZN( u0_u5_u7_n110 ) , .A1( u0_u5_u7_n95 ) , .A2( u0_u5_u7_n96 ) );
  INV_X1 u0_u5_u7_U61 (.A( u0_u5_u7_n150 ) , .ZN( u0_u5_u7_n164 ) );
  AND2_X1 u0_u5_u7_U62 (.ZN( u0_u5_u7_n134 ) , .A1( u0_u5_u7_n93 ) , .A2( u0_u5_u7_n98 ) );
  NAND2_X1 u0_u5_u7_U63 (.A1( u0_u5_u7_n100 ) , .A2( u0_u5_u7_n102 ) , .ZN( u0_u5_u7_n129 ) );
  NAND2_X1 u0_u5_u7_U64 (.A2( u0_u5_u7_n103 ) , .ZN( u0_u5_u7_n131 ) , .A1( u0_u5_u7_n95 ) );
  NAND2_X1 u0_u5_u7_U65 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n138 ) , .A2( u0_u5_u7_n99 ) );
  NAND2_X1 u0_u5_u7_U66 (.ZN( u0_u5_u7_n132 ) , .A1( u0_u5_u7_n93 ) , .A2( u0_u5_u7_n96 ) );
  NAND2_X1 u0_u5_u7_U67 (.A1( u0_u5_u7_n100 ) , .ZN( u0_u5_u7_n148 ) , .A2( u0_u5_u7_n95 ) );
  NOR2_X1 u0_u5_u7_U68 (.A2( u0_u5_X_47 ) , .ZN( u0_u5_u7_n150 ) , .A1( u0_u5_u7_n163 ) );
  NOR2_X1 u0_u5_u7_U69 (.A2( u0_u5_X_43 ) , .A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n103 ) );
  AOI211_X1 u0_u5_u7_U7 (.ZN( u0_u5_u7_n116 ) , .A( u0_u5_u7_n155 ) , .C1( u0_u5_u7_n161 ) , .C2( u0_u5_u7_n171 ) , .B( u0_u5_u7_n94 ) );
  NOR2_X1 u0_u5_u7_U70 (.A2( u0_u5_X_48 ) , .A1( u0_u5_u7_n166 ) , .ZN( u0_u5_u7_n95 ) );
  NOR2_X1 u0_u5_u7_U71 (.A2( u0_u5_X_45 ) , .A1( u0_u5_X_48 ) , .ZN( u0_u5_u7_n99 ) );
  NOR2_X1 u0_u5_u7_U72 (.A2( u0_u5_X_44 ) , .A1( u0_u5_u7_n167 ) , .ZN( u0_u5_u7_n98 ) );
  NOR2_X1 u0_u5_u7_U73 (.A2( u0_u5_X_46 ) , .A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n152 ) );
  AND2_X1 u0_u5_u7_U74 (.A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n156 ) , .A2( u0_u5_u7_n163 ) );
  NAND2_X1 u0_u5_u7_U75 (.A2( u0_u5_X_46 ) , .A1( u0_u5_X_47 ) , .ZN( u0_u5_u7_n125 ) );
  AND2_X1 u0_u5_u7_U76 (.A2( u0_u5_X_45 ) , .A1( u0_u5_X_48 ) , .ZN( u0_u5_u7_n102 ) );
  AND2_X1 u0_u5_u7_U77 (.A2( u0_u5_X_43 ) , .A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n96 ) );
  AND2_X1 u0_u5_u7_U78 (.A1( u0_u5_X_44 ) , .ZN( u0_u5_u7_n100 ) , .A2( u0_u5_u7_n167 ) );
  AND2_X1 u0_u5_u7_U79 (.A1( u0_u5_X_48 ) , .A2( u0_u5_u7_n166 ) , .ZN( u0_u5_u7_n93 ) );
  OAI222_X1 u0_u5_u7_U8 (.C2( u0_u5_u7_n101 ) , .B2( u0_u5_u7_n111 ) , .A1( u0_u5_u7_n113 ) , .C1( u0_u5_u7_n146 ) , .A2( u0_u5_u7_n162 ) , .B1( u0_u5_u7_n164 ) , .ZN( u0_u5_u7_n94 ) );
  INV_X1 u0_u5_u7_U80 (.A( u0_u5_X_46 ) , .ZN( u0_u5_u7_n163 ) );
  INV_X1 u0_u5_u7_U81 (.A( u0_u5_X_43 ) , .ZN( u0_u5_u7_n167 ) );
  INV_X1 u0_u5_u7_U82 (.A( u0_u5_X_45 ) , .ZN( u0_u5_u7_n166 ) );
  NAND4_X1 u0_u5_u7_U83 (.ZN( u0_out5_27 ) , .A4( u0_u5_u7_n118 ) , .A3( u0_u5_u7_n119 ) , .A2( u0_u5_u7_n120 ) , .A1( u0_u5_u7_n121 ) );
  OAI21_X1 u0_u5_u7_U84 (.ZN( u0_u5_u7_n121 ) , .B2( u0_u5_u7_n145 ) , .A( u0_u5_u7_n150 ) , .B1( u0_u5_u7_n174 ) );
  OAI21_X1 u0_u5_u7_U85 (.ZN( u0_u5_u7_n120 ) , .A( u0_u5_u7_n161 ) , .B2( u0_u5_u7_n170 ) , .B1( u0_u5_u7_n179 ) );
  NAND4_X1 u0_u5_u7_U86 (.ZN( u0_out5_21 ) , .A4( u0_u5_u7_n157 ) , .A3( u0_u5_u7_n158 ) , .A2( u0_u5_u7_n159 ) , .A1( u0_u5_u7_n160 ) );
  OAI21_X1 u0_u5_u7_U87 (.B1( u0_u5_u7_n145 ) , .ZN( u0_u5_u7_n160 ) , .A( u0_u5_u7_n161 ) , .B2( u0_u5_u7_n177 ) );
  AOI22_X1 u0_u5_u7_U88 (.B2( u0_u5_u7_n149 ) , .B1( u0_u5_u7_n150 ) , .A2( u0_u5_u7_n151 ) , .A1( u0_u5_u7_n152 ) , .ZN( u0_u5_u7_n158 ) );
  NAND4_X1 u0_u5_u7_U89 (.ZN( u0_out5_15 ) , .A4( u0_u5_u7_n142 ) , .A3( u0_u5_u7_n143 ) , .A2( u0_u5_u7_n144 ) , .A1( u0_u5_u7_n178 ) );
  OAI221_X1 u0_u5_u7_U9 (.C1( u0_u5_u7_n101 ) , .C2( u0_u5_u7_n147 ) , .ZN( u0_u5_u7_n155 ) , .B2( u0_u5_u7_n162 ) , .A( u0_u5_u7_n91 ) , .B1( u0_u5_u7_n92 ) );
  OR2_X1 u0_u5_u7_U90 (.A2( u0_u5_u7_n125 ) , .A1( u0_u5_u7_n129 ) , .ZN( u0_u5_u7_n144 ) );
  AOI22_X1 u0_u5_u7_U91 (.A2( u0_u5_u7_n126 ) , .ZN( u0_u5_u7_n143 ) , .B2( u0_u5_u7_n165 ) , .B1( u0_u5_u7_n173 ) , .A1( u0_u5_u7_n174 ) );
  NAND4_X1 u0_u5_u7_U92 (.ZN( u0_out5_5 ) , .A4( u0_u5_u7_n108 ) , .A3( u0_u5_u7_n109 ) , .A1( u0_u5_u7_n116 ) , .A2( u0_u5_u7_n123 ) );
  AOI22_X1 u0_u5_u7_U93 (.ZN( u0_u5_u7_n109 ) , .A2( u0_u5_u7_n126 ) , .B2( u0_u5_u7_n145 ) , .B1( u0_u5_u7_n156 ) , .A1( u0_u5_u7_n171 ) );
  NOR4_X1 u0_u5_u7_U94 (.A4( u0_u5_u7_n104 ) , .A3( u0_u5_u7_n105 ) , .A2( u0_u5_u7_n106 ) , .A1( u0_u5_u7_n107 ) , .ZN( u0_u5_u7_n108 ) );
  NAND3_X1 u0_u5_u7_U95 (.A3( u0_u5_u7_n146 ) , .A2( u0_u5_u7_n147 ) , .A1( u0_u5_u7_n148 ) , .ZN( u0_u5_u7_n151 ) );
  NAND3_X1 u0_u5_u7_U96 (.A3( u0_u5_u7_n131 ) , .A2( u0_u5_u7_n132 ) , .A1( u0_u5_u7_n133 ) , .ZN( u0_u5_u7_n135 ) );
  INV_X1 u0_uk_U10 (.A( u0_uk_n252 ) , .ZN( u0_uk_n31 ) );
  OAI21_X1 u0_uk_U1030 (.ZN( u0_K16_41 ) , .B1( u0_uk_n142 ) , .B2( u0_uk_n643 ) , .A( u0_uk_n898 ) );
  INV_X1 u0_uk_U1064 (.A( u0_key_r_6 ) , .ZN( u0_uk_n712 ) );
  INV_X1 u0_uk_U1065 (.A( u0_key_r_54 ) , .ZN( u0_uk_n673 ) );
  OAI22_X1 u0_uk_U107 (.ZN( u0_K1_5 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n708 ) , .A2( u0_uk_n712 ) , .B1( u0_uk_n99 ) );
  INV_X1 u0_uk_U1073 (.A( u0_key_r_20 ) , .ZN( u0_uk_n703 ) );
  INV_X1 u0_uk_U1078 (.A( u0_key_r_13 ) , .ZN( u0_uk_n708 ) );
  INV_X1 u0_uk_U1081 (.A( u0_key_r_19 ) , .ZN( u0_uk_n704 ) );
  INV_X1 u0_uk_U1082 (.A( u0_key_r_4 ) , .ZN( u0_uk_n713 ) );
  OAI21_X1 u0_uk_U1093 (.ZN( u0_K16_39 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n657 ) , .A( u0_uk_n899 ) );
  NAND2_X1 u0_uk_U1094 (.A1( u0_uk_K_r14_15 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n899 ) );
  OAI22_X1 u0_uk_U110 (.ZN( u0_K12_41 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n144 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n153 ) );
  INV_X1 u0_uk_U1100 (.A( u0_key_r_47 ) , .ZN( u0_uk_n679 ) );
  INV_X1 u0_uk_U1103 (.ZN( u0_K1_11 ) , .A( u0_uk_n892 ) );
  INV_X1 u0_uk_U1105 (.ZN( u0_K1_18 ) , .A( u0_uk_n887 ) );
  AOI22_X1 u0_uk_U1106 (.A2( u0_key_r_5 ) , .B2( u0_key_r_55 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n887 ) );
  INV_X1 u0_uk_U1109 (.ZN( u0_K11_8 ) , .A( u0_uk_n982 ) );
  INV_X1 u0_uk_U1111 (.ZN( u0_K11_12 ) , .A( u0_uk_n1003 ) );
  AOI22_X1 u0_uk_U1112 (.B2( u0_uk_K_r9_25 ) , .A2( u0_uk_K_r9_6 ) , .ZN( u0_uk_n1003 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n207 ) );
  INV_X1 u0_uk_U1115 (.ZN( u0_K1_20 ) , .A( u0_uk_n886 ) );
  AOI22_X1 u0_uk_U1116 (.B2( u0_key_r_48 ) , .A2( u0_key_r_55 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n886 ) );
  OAI22_X1 u0_uk_U113 (.ZN( u0_K13_47 ) , .B2( u0_uk_n106 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n96 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U1131 (.ZN( u0_K12_42 ) , .A( u0_uk_n966 ) );
  AOI22_X1 u0_uk_U1132 (.B2( u0_uk_K_r10_28 ) , .A2( u0_uk_K_r10_9 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n966 ) );
  INV_X1 u0_uk_U1156 (.ZN( u0_K6_2 ) , .A( u0_uk_n793 ) );
  OAI22_X1 u0_uk_U1157 (.ZN( u0_K1_1 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n679 ) , .B2( u0_uk_n684 ) );
  INV_X1 u0_uk_U1159 (.ZN( u0_K13_6 ) , .A( u0_uk_n940 ) );
  OAI21_X1 u0_uk_U120 (.ZN( u0_K6_47 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n439 ) , .A( u0_uk_n789 ) );
  NAND2_X1 u0_uk_U121 (.A1( u0_uk_K_r4_23 ) , .ZN( u0_uk_n789 ) , .A2( u0_uk_n93 ) );
  INV_X1 u0_uk_U13 (.A( u0_uk_n252 ) , .ZN( u0_uk_n60 ) );
  INV_X1 u0_uk_U130 (.ZN( u0_K13_15 ) , .A( u0_uk_n956 ) );
  INV_X1 u0_uk_U136 (.ZN( u0_K13_19 ) , .A( u0_uk_n953 ) );
  AOI22_X1 u0_uk_U137 (.B2( u0_uk_K_r11_19 ) , .A2( u0_uk_K_r11_39 ) , .B1( u0_uk_n207 ) , .A1( u0_uk_n94 ) , .ZN( u0_uk_n953 ) );
  OAI22_X1 u0_uk_U139 (.ZN( u0_K11_15 ) , .A1( u0_uk_n147 ) , .A2( u0_uk_n197 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U144 (.ZN( u0_K1_19 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n673 ) , .B2( u0_uk_n713 ) );
  INV_X1 u0_uk_U151 (.ZN( u0_K11_19 ) , .A( u0_uk_n1000 ) );
  INV_X1 u0_uk_U16 (.ZN( u0_uk_n110 ) , .A( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U179 (.ZN( u0_K12_24 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n143 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n172 ) );
  INV_X1 u0_uk_U18 (.ZN( u0_uk_n117 ) , .A( u0_uk_n182 ) );
  INV_X1 u0_uk_U180 (.ZN( u0_K11_14 ) , .A( u0_uk_n1002 ) );
  OAI22_X1 u0_uk_U186 (.ZN( u0_K6_14 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n442 ) , .A2( u0_uk_n448 ) );
  OAI22_X1 u0_uk_U189 (.ZN( u0_K1_24 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n703 ) , .B2( u0_uk_n708 ) );
  INV_X1 u0_uk_U21 (.ZN( u0_uk_n102 ) , .A( u0_uk_n162 ) );
  OAI21_X1 u0_uk_U216 (.ZN( u0_K12_31 ) , .B2( u0_uk_n173 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n973 ) );
  NAND2_X1 u0_uk_U217 (.A1( u0_uk_K_r10_44 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n973 ) );
  OAI22_X1 u0_uk_U228 (.ZN( u0_K6_31 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n428 ) , .B2( u0_uk_n433 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U23 (.ZN( u0_uk_n10 ) , .A( u0_uk_n148 ) );
  INV_X1 u0_uk_U24 (.ZN( u0_uk_n11 ) , .A( u0_uk_n242 ) );
  INV_X1 u0_uk_U26 (.ZN( u0_uk_n129 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U268 (.ZN( u0_K6_44 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n412 ) , .B2( u0_uk_n430 ) );
  OAI22_X1 u0_uk_U269 (.ZN( u0_K6_48 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n425 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U27 (.Z( u0_uk_n163 ) , .A( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U279 (.ZN( u0_K6_6 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n410 ) , .B2( u0_uk_n414 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U28 (.Z( u0_uk_n147 ) , .A( u0_uk_n250 ) );
  OAI21_X1 u0_uk_U280 (.ZN( u0_K6_8 ) , .B2( u0_uk_n442 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n786 ) );
  OAI22_X1 u0_uk_U283 (.ZN( u0_K1_8 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n699 ) , .A2( u0_uk_n712 ) );
  BUF_X1 u0_uk_U29 (.Z( u0_uk_n162 ) , .A( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U293 (.ZN( u0_K3_8 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n562 ) , .A2( u0_uk_n578 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U3 (.ZN( u0_uk_n142 ) , .A( u0_uk_n191 ) );
  OAI21_X1 u0_uk_U306 (.ZN( u0_K6_26 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n419 ) , .A( u0_uk_n795 ) );
  NAND2_X1 u0_uk_U307 (.A1( u0_uk_K_r4_35 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n795 ) );
  INV_X1 u0_uk_U341 (.ZN( u0_K6_4 ) , .A( u0_uk_n788 ) );
  AOI22_X1 u0_uk_U342 (.B2( u0_uk_K_r4_41 ) , .A2( u0_uk_K_r4_47 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n788 ) );
  OAI22_X1 u0_uk_U347 (.ZN( u0_K3_4 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n557 ) , .B2( u0_uk_n565 ) , .B1( u0_uk_n63 ) );
  OAI21_X1 u0_uk_U349 (.ZN( u0_K1_4 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n674 ) , .A( u0_uk_n869 ) );
  OAI22_X1 u0_uk_U351 (.ZN( u0_K16_40 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n632 ) , .B2( u0_uk_n670 ) );
  OAI22_X1 u0_uk_U352 (.ZN( u0_K6_40 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n438 ) , .A2( u0_uk_n446 ) );
  BUF_X1 u0_uk_U37 (.Z( u0_uk_n182 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U375 (.ZN( u0_K6_28 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n411 ) , .B2( u0_uk_n438 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U38 (.Z( u0_uk_n203 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U389 (.ZN( u0_K3_1 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n568 ) , .B2( u0_uk_n573 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U39 (.Z( u0_uk_n202 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U391 (.ZN( u0_K1_9 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n673 ) , .B2( u0_uk_n679 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U392 (.ZN( u0_K13_16 ) , .A1( u0_uk_n118 ) , .A2( u0_uk_n122 ) , .B2( u0_uk_n127 ) , .B1( u0_uk_n242 ) );
  INV_X1 u0_uk_U4 (.ZN( u0_uk_n145 ) , .A( u0_uk_n242 ) );
  OAI22_X1 u0_uk_U406 (.ZN( u0_K13_9 ) , .A2( u0_uk_n115 ) , .B2( u0_uk_n127 ) , .A1( u0_uk_n230 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U408 (.ZN( u0_K11_9 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n195 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n225 ) );
  INV_X1 u0_uk_U410 (.ZN( u0_K2_28 ) , .A( u0_uk_n861 ) );
  AOI22_X1 u0_uk_U411 (.B2( u0_uk_K_r0_15 ) , .A2( u0_uk_K_r0_49 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n861 ) );
  BUF_X1 u0_uk_U42 (.Z( u0_uk_n238 ) , .A( u0_uk_n252 ) );
  BUF_X1 u0_uk_U43 (.Z( u0_uk_n220 ) , .A( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U448 (.ZN( u0_K6_33 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n425 ) , .B2( u0_uk_n430 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U452 (.ZN( u0_K16_37 ) , .A( u0_uk_n900 ) );
  AOI22_X1 u0_uk_U453 (.B2( u0_uk_K_r14_2 ) , .A2( u0_uk_K_r14_50 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n900 ) );
  OAI22_X1 u0_uk_U456 (.ZN( u0_K12_37 ) , .A2( u0_uk_n139 ) , .B2( u0_uk_n179 ) , .A1( u0_uk_n238 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U461 (.ZN( u0_K6_37 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n420 ) , .A( u0_uk_n791 ) );
  NAND2_X1 u0_uk_U462 (.A1( u0_uk_K_r4_38 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n791 ) );
  BUF_X1 u0_uk_U47 (.Z( u0_uk_n217 ) , .A( u0_uk_n240 ) );
  OAI21_X1 u0_uk_U477 (.ZN( u0_K6_29 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n446 ) , .A( u0_uk_n794 ) );
  NAND2_X1 u0_uk_U478 (.A1( u0_uk_K_r4_0 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n794 ) );
  BUF_X1 u0_uk_U48 (.Z( u0_uk_n222 ) , .A( u0_uk_n250 ) );
  BUF_X1 u0_uk_U49 (.Z( u0_uk_n231 ) , .A( u0_uk_n250 ) );
  OAI22_X1 u0_uk_U491 (.ZN( u0_K3_2 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n552 ) , .B2( u0_uk_n557 ) , .B1( u0_uk_n63 ) );
  OAI21_X1 u0_uk_U495 (.ZN( u0_K1_2 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n713 ) , .A( u0_uk_n881 ) );
  NAND2_X1 u0_uk_U496 (.A1( u0_key_r_11 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n881 ) );
  OAI21_X1 u0_uk_U499 (.ZN( u0_K1_12 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n704 ) , .A( u0_uk_n891 ) );
  INV_X1 u0_uk_U5 (.ZN( u0_uk_n141 ) , .A( u0_uk_n191 ) );
  NAND2_X1 u0_uk_U500 (.A1( u0_key_r_12 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n891 ) );
  OAI21_X1 u0_uk_U501 (.ZN( u0_K13_17 ) , .B2( u0_uk_n115 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n955 ) );
  NAND2_X1 u0_uk_U502 (.A1( u0_uk_K_r11_27 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n955 ) );
  INV_X1 u0_uk_U508 (.ZN( u0_K11_17 ) , .A( u0_uk_n1001 ) );
  BUF_X1 u0_uk_U51 (.A( u0_uk_n161 ) , .Z( u0_uk_n242 ) );
  BUF_X1 u0_uk_U52 (.Z( u0_uk_n207 ) , .A( u0_uk_n217 ) );
  BUF_X1 u0_uk_U53 (.A( u0_uk_n163 ) , .Z( u0_uk_n208 ) );
  BUF_X1 u0_uk_U54 (.Z( u0_uk_n251 ) , .A( u0_uk_n257 ) );
  INV_X1 u0_uk_U540 (.ZN( u0_K12_17 ) , .A( u0_uk_n979 ) );
  AOI22_X1 u0_uk_U541 (.B2( u0_uk_K_r10_18 ) , .A2( u0_uk_K_r10_41 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n979 ) );
  INV_X1 u0_uk_U542 (.ZN( u0_K6_17 ) , .A( u0_uk_n800 ) );
  BUF_X1 u0_uk_U55 (.A( u0_uk_n250 ) , .Z( u0_uk_n252 ) );
  OAI22_X1 u0_uk_U555 (.ZN( u0_K12_38 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n153 ) , .B2( u0_uk_n180 ) );
  BUF_X1 u0_uk_U56 (.Z( u0_uk_n250 ) , .A( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U567 (.ZN( u0_K6_38 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n433 ) , .B2( u0_uk_n440 ) , .B1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U575 (.ZN( u0_K11_10 ) , .A( u0_uk_n1004 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n225 ) );
  INV_X1 u0_uk_U586 (.ZN( u0_K1_10 ) , .A( u0_uk_n893 ) );
  AOI22_X1 u0_uk_U587 (.B2( u0_key_r_41 ) , .A2( u0_key_r_48 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n893 ) );
  INV_X1 u0_uk_U590 (.ZN( u0_K13_22 ) , .A( u0_uk_n949 ) );
  OAI22_X1 u0_uk_U618 (.ZN( u0_K6_35 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n412 ) , .B2( u0_uk_n419 ) , .B1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U624 (.ZN( u0_K15_11 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n8 ) , .A( u0_uk_n924 ) );
  NAND2_X1 u0_uk_U625 (.A1( u0_uk_K_r13_25 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n924 ) );
  OAI22_X1 u0_uk_U627 (.ZN( u0_K11_11 ) , .A1( u0_uk_n145 ) , .A2( u0_uk_n206 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U634 (.ZN( u0_K3_11 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n573 ) , .A2( u0_uk_n578 ) );
  INV_X1 u0_uk_U641 (.ZN( u0_K12_23 ) , .A( u0_uk_n975 ) );
  AOI22_X1 u0_uk_U642 (.B2( u0_uk_K_r10_32 ) , .A2( u0_uk_K_r10_41 ) , .A1( u0_uk_n220 ) , .B1( u0_uk_n83 ) , .ZN( u0_uk_n975 ) );
  OAI22_X1 u0_uk_U656 (.ZN( u0_K1_7 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n696 ) , .B2( u0_uk_n703 ) );
  OAI21_X1 u0_uk_U662 (.ZN( u0_K14_45 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n58 ) , .A( u0_uk_n929 ) );
  NAND2_X1 u0_uk_U663 (.A1( u0_uk_K_r12_16 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n929 ) );
  OAI21_X1 u0_uk_U664 (.ZN( u0_K13_43 ) , .B1( u0_uk_n252 ) , .A( u0_uk_n943 ) , .B2( u0_uk_n96 ) );
  NAND2_X1 u0_uk_U665 (.A1( u0_uk_K_r11_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n943 ) );
  OAI21_X1 u0_uk_U682 (.ZN( u0_K11_7 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n197 ) , .A( u0_uk_n983 ) );
  NAND2_X1 u0_uk_U683 (.A1( u0_uk_K_r9_33 ) , .A2( u0_uk_n146 ) , .ZN( u0_uk_n983 ) );
  OAI21_X1 u0_uk_U699 (.ZN( u0_K6_7 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n423 ) , .A( u0_uk_n787 ) );
  NAND2_X1 u0_uk_U700 (.A1( u0_uk_K_r4_33 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n787 ) );
  OAI22_X1 u0_uk_U721 (.ZN( u0_K6_32 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n424 ) , .B2( u0_uk_n440 ) );
  INV_X1 u0_uk_U738 (.ZN( u0_K12_32 ) , .A( u0_uk_n972 ) );
  AOI22_X1 u0_uk_U739 (.B2( u0_uk_K_r10_23 ) , .A2( u0_uk_K_r10_28 ) , .A1( u0_uk_n251 ) , .B1( u0_uk_n60 ) , .ZN( u0_uk_n972 ) );
  INV_X1 u0_uk_U740 (.ZN( u0_K2_32 ) , .A( u0_uk_n860 ) );
  AOI22_X1 u0_uk_U741 (.B2( u0_uk_K_r0_15 ) , .A2( u0_uk_K_r0_36 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n231 ) , .ZN( u0_uk_n860 ) );
  OAI21_X1 u0_uk_U75 (.ZN( u0_K11_23 ) , .B2( u0_uk_n190 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n996 ) );
  OAI22_X1 u0_uk_U752 (.ZN( u0_K11_13 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n196 ) , .B2( u0_uk_n200 ) );
  NAND2_X1 u0_uk_U76 (.A1( u0_uk_K_r9_27 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n996 ) );
  INV_X1 u0_uk_U776 (.ZN( u0_K2_27 ) , .A( u0_uk_n862 ) );
  AOI22_X1 u0_uk_U777 (.B2( u0_uk_K_r0_28 ) , .A2( u0_uk_K_r0_7 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n862 ) );
  INV_X1 u0_uk_U782 (.ZN( u0_K13_21 ) , .A( u0_uk_n950 ) );
  INV_X1 u0_uk_U784 (.ZN( u0_K12_21 ) , .A( u0_uk_n976 ) );
  OAI22_X1 u0_uk_U799 (.ZN( u0_K6_1 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n410 ) , .B2( u0_uk_n426 ) );
  OAI21_X1 u0_uk_U808 (.ZN( u0_K13_20 ) , .B2( u0_uk_n126 ) , .B1( u0_uk_n92 ) , .A( u0_uk_n951 ) );
  NAND2_X1 u0_uk_U809 (.A1( u0_uk_K_r11_33 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n951 ) );
  OAI21_X1 u0_uk_U819 (.ZN( u0_K13_18 ) , .B2( u0_uk_n108 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n954 ) );
  NAND2_X1 u0_uk_U820 (.A1( u0_uk_K_r11_20 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n954 ) );
  INV_X1 u0_uk_U827 (.ZN( u0_K6_18 ) , .A( u0_uk_n799 ) );
  INV_X1 u0_uk_U829 (.ZN( u0_K11_20 ) , .A( u0_uk_n999 ) );
  OAI21_X1 u0_uk_U835 (.ZN( u0_K13_1 ) , .B2( u0_uk_n131 ) , .B1( u0_uk_n31 ) , .A( u0_uk_n952 ) );
  NAND2_X1 u0_uk_U836 (.A1( u0_uk_K_r11_25 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n952 ) );
  OAI22_X1 u0_uk_U840 (.ZN( u0_K1_6 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n683 ) , .B2( u0_uk_n690 ) );
  INV_X1 u0_uk_U841 (.A( u0_key_r_41 ) , .ZN( u0_uk_n683 ) );
  OAI21_X1 u0_uk_U847 (.ZN( u0_K13_3 ) , .B2( u0_uk_n107 ) , .B1( u0_uk_n31 ) , .A( u0_uk_n944 ) );
  NAND2_X1 u0_uk_U848 (.A1( u0_uk_K_r11_4 ) , .A2( u0_uk_n129 ) , .ZN( u0_uk_n944 ) );
  INV_X1 u0_uk_U86 (.ZN( u0_K2_41 ) , .A( u0_uk_n858 ) );
  AOI22_X1 u0_uk_U866 (.B2( u0_uk_K_r11_19 ) , .A2( u0_uk_K_r11_24 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n940 ) );
  AOI22_X1 u0_uk_U87 (.B2( u0_uk_K_r0_28 ) , .A2( u0_uk_K_r0_49 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n858 ) );
  OAI22_X1 u0_uk_U880 (.ZN( u0_K6_5 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n432 ) , .B2( u0_uk_n436 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U889 (.ZN( u0_K6_45 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n429 ) , .B2( u0_uk_n434 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U897 (.ZN( u0_K6_12 ) , .A1( u0_uk_n257 ) , .B2( u0_uk_n432 ) , .A2( u0_uk_n448 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U918 (.ZN( u0_K6_30 ) , .A1( u0_uk_n203 ) , .A2( u0_uk_n445 ) , .B2( u0_uk_n450 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U923 (.ZN( u0_K6_42 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n413 ) , .B2( u0_uk_n420 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U924 (.ZN( u0_K6_39 ) , .A1( u0_uk_n162 ) , .B2( u0_uk_n428 ) , .A2( u0_uk_n447 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U929 (.ZN( u0_K13_23 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n121 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n91 ) );
  OAI22_X1 u0_uk_U933 (.ZN( u0_K11_16 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n190 ) , .B2( u0_uk_n196 ) );
  OAI22_X1 u0_uk_U942 (.ZN( u0_K11_24 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n201 ) , .B2( u0_uk_n206 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U952 (.ZN( u0_K13_4 ) , .A1( u0_uk_n117 ) , .A2( u0_uk_n121 ) , .B2( u0_uk_n126 ) , .B1( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U957 (.ZN( u0_K13_8 ) , .A2( u0_uk_n101 ) , .B2( u0_uk_n107 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n147 ) );
  OAI22_X1 u0_uk_U959 (.ZN( u0_K11_18 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n215 ) , .B2( u0_uk_n221 ) );
  OAI22_X1 u0_uk_U965 (.ZN( u0_K6_36 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n439 ) , .A2( u0_uk_n447 ) );
  OAI22_X1 u0_uk_U977 (.ZN( u0_K6_43 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n411 ) , .B2( u0_uk_n450 ) );
  OAI22_X1 u0_uk_U985 (.ZN( u0_K3_7 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n547 ) , .B2( u0_uk_n565 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U988 (.ZN( u0_K6_25 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n434 ) );
  OAI22_X1 u0_uk_U993 (.ZN( u0_K1_3 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n697 ) , .B2( u0_uk_n704 ) );
  XOR2_X1 u1_u0_U12 (.B( u1_K1_43 ) , .A( u1_desIn_r_25 ) , .Z( u1_u0_X_43 ) );
  XOR2_X1 u1_u0_U14 (.B( u1_K1_41 ) , .A( u1_desIn_r_25 ) , .Z( u1_u0_X_41 ) );
  XOR2_X1 u1_u0_U2 (.B( u1_K1_8 ) , .A( u1_desIn_r_39 ) , .Z( u1_u0_X_8 ) );
  XOR2_X1 u1_u0_U38 (.B( u1_K1_1 ) , .A( u1_desIn_r_57 ) , .Z( u1_u0_X_1 ) );
  XOR2_X1 u1_u0_U4 (.B( u1_K1_6 ) , .A( u1_desIn_r_39 ) , .Z( u1_u0_X_6 ) );
  XOR2_X1 u1_u0_U8 (.B( u1_K1_47 ) , .A( u1_desIn_r_57 ) , .Z( u1_u0_X_47 ) );
  NAND2_X1 u1_u0_u0_U10 (.ZN( u1_u0_u0_n113 ) , .A1( u1_u0_u0_n139 ) , .A2( u1_u0_u0_n149 ) );
  AND3_X1 u1_u0_u0_U11 (.A2( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n127 ) , .A3( u1_u0_u0_n130 ) , .A1( u1_u0_u0_n148 ) );
  AND2_X1 u1_u0_u0_U12 (.ZN( u1_u0_u0_n107 ) , .A1( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n140 ) );
  AND2_X1 u1_u0_u0_U13 (.A2( u1_u0_u0_n129 ) , .A1( u1_u0_u0_n130 ) , .ZN( u1_u0_u0_n151 ) );
  AND2_X1 u1_u0_u0_U14 (.A1( u1_u0_u0_n108 ) , .A2( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U15 (.A( u1_u0_u0_n143 ) , .ZN( u1_u0_u0_n173 ) );
  NOR2_X1 u1_u0_u0_U16 (.A2( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n147 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U17 (.ZN( u1_u0_u0_n172 ) , .A( u1_u0_u0_n88 ) );
  OAI222_X1 u1_u0_u0_U18 (.C1( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n125 ) , .B2( u1_u0_u0_n128 ) , .B1( u1_u0_u0_n144 ) , .A2( u1_u0_u0_n158 ) , .C2( u1_u0_u0_n161 ) , .ZN( u1_u0_u0_n88 ) );
  AOI21_X1 u1_u0_u0_U19 (.B1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n132 ) , .A( u1_u0_u0_n165 ) , .B2( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U20 (.A( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n165 ) );
  OAI22_X1 u1_u0_u0_U21 (.B1( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n126 ) , .A1( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n146 ) , .B2( u1_u0_u0_n147 ) );
  OAI22_X1 u1_u0_u0_U22 (.B1( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n147 ) , .A2( u1_u0_u0_n90 ) , .ZN( u1_u0_u0_n91 ) );
  AND3_X1 u1_u0_u0_U23 (.A3( u1_u0_u0_n121 ) , .A2( u1_u0_u0_n125 ) , .A1( u1_u0_u0_n148 ) , .ZN( u1_u0_u0_n90 ) );
  INV_X1 u1_u0_u0_U24 (.A( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n161 ) );
  AOI22_X1 u1_u0_u0_U25 (.B2( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n110 ) , .ZN( u1_u0_u0_n111 ) , .B1( u1_u0_u0_n118 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U26 (.A( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U27 (.B1( u1_u0_u0_n127 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n96 ) );
  AOI21_X1 u1_u0_u0_U28 (.ZN( u1_u0_u0_n104 ) , .B1( u1_u0_u0_n107 ) , .B2( u1_u0_u0_n141 ) , .A( u1_u0_u0_n144 ) );
  NAND2_X1 u1_u0_u0_U29 (.A1( u1_u0_u0_n100 ) , .A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n125 ) );
  INV_X1 u1_u0_u0_U3 (.A( u1_u0_u0_n113 ) , .ZN( u1_u0_u0_n166 ) );
  NAND2_X1 u1_u0_u0_U30 (.A2( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n92 ) );
  NAND2_X1 u1_u0_u0_U31 (.A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n114 ) , .A1( u1_u0_u0_n92 ) );
  NOR2_X1 u1_u0_u0_U32 (.A1( u1_u0_u0_n120 ) , .ZN( u1_u0_u0_n143 ) , .A2( u1_u0_u0_n167 ) );
  OAI221_X1 u1_u0_u0_U33 (.C1( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n120 ) , .B1( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n141 ) , .C2( u1_u0_u0_n147 ) , .A( u1_u0_u0_n172 ) );
  AOI21_X1 u1_u0_u0_U34 (.ZN( u1_u0_u0_n116 ) , .B2( u1_u0_u0_n142 ) , .A( u1_u0_u0_n144 ) , .B1( u1_u0_u0_n166 ) );
  INV_X1 u1_u0_u0_U35 (.A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n160 ) );
  NAND2_X1 u1_u0_u0_U36 (.A2( u1_u0_u0_n102 ) , .A1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n149 ) );
  NAND2_X1 u1_u0_u0_U37 (.ZN( u1_u0_u0_n112 ) , .A2( u1_u0_u0_n92 ) , .A1( u1_u0_u0_n93 ) );
  OR3_X1 u1_u0_u0_U38 (.A3( u1_u0_u0_n152 ) , .A2( u1_u0_u0_n153 ) , .A1( u1_u0_u0_n154 ) , .ZN( u1_u0_u0_n155 ) );
  AOI21_X1 u1_u0_u0_U39 (.B2( u1_u0_u0_n150 ) , .B1( u1_u0_u0_n151 ) , .ZN( u1_u0_u0_n152 ) , .A( u1_u0_u0_n158 ) );
  NOR2_X1 u1_u0_u0_U4 (.A1( u1_u0_u0_n108 ) , .ZN( u1_u0_u0_n123 ) , .A2( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U40 (.A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n145 ) , .B1( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n154 ) );
  AOI21_X1 u1_u0_u0_U41 (.A( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n148 ) , .B1( u1_u0_u0_n149 ) , .ZN( u1_u0_u0_n153 ) );
  INV_X1 u1_u0_u0_U42 (.ZN( u1_u0_u0_n171 ) , .A( u1_u0_u0_n99 ) );
  OAI211_X1 u1_u0_u0_U43 (.C2( u1_u0_u0_n140 ) , .C1( u1_u0_u0_n161 ) , .A( u1_u0_u0_n169 ) , .B( u1_u0_u0_n98 ) , .ZN( u1_u0_u0_n99 ) );
  AOI211_X1 u1_u0_u0_U44 (.C1( u1_u0_u0_n118 ) , .A( u1_u0_u0_n123 ) , .B( u1_u0_u0_n96 ) , .C2( u1_u0_u0_n97 ) , .ZN( u1_u0_u0_n98 ) );
  INV_X1 u1_u0_u0_U45 (.ZN( u1_u0_u0_n169 ) , .A( u1_u0_u0_n91 ) );
  NOR2_X1 u1_u0_u0_U46 (.A2( u1_u0_X_2 ) , .ZN( u1_u0_u0_n103 ) , .A1( u1_u0_u0_n164 ) );
  NOR2_X1 u1_u0_u0_U47 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n118 ) );
  NAND2_X1 u1_u0_u0_U48 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n144 ) );
  NOR2_X1 u1_u0_u0_U49 (.A2( u1_u0_X_5 ) , .ZN( u1_u0_u0_n136 ) , .A1( u1_u0_u0_n159 ) );
  AOI21_X1 u1_u0_u0_U5 (.B2( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n134 ) , .B1( u1_u0_u0_n151 ) , .A( u1_u0_u0_n158 ) );
  NAND2_X1 u1_u0_u0_U50 (.A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n159 ) );
  AND2_X1 u1_u0_u0_U51 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n102 ) );
  AND2_X1 u1_u0_u0_U52 (.A1( u1_u0_X_6 ) , .A2( u1_u0_u0_n162 ) , .ZN( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U53 (.A( u1_u0_X_4 ) , .ZN( u1_u0_u0_n159 ) );
  INV_X1 u1_u0_u0_U54 (.A( u1_u0_X_2 ) , .ZN( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U55 (.A( u1_u0_X_3 ) , .ZN( u1_u0_u0_n162 ) );
  INV_X1 u1_u0_u0_U56 (.A( u1_u0_u0_n126 ) , .ZN( u1_u0_u0_n168 ) );
  AOI211_X1 u1_u0_u0_U57 (.B( u1_u0_u0_n133 ) , .A( u1_u0_u0_n134 ) , .C2( u1_u0_u0_n135 ) , .C1( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n137 ) );
  OR4_X1 u1_u0_u0_U58 (.ZN( u1_out0_17 ) , .A4( u1_u0_u0_n122 ) , .A2( u1_u0_u0_n123 ) , .A1( u1_u0_u0_n124 ) , .A3( u1_u0_u0_n170 ) );
  AOI21_X1 u1_u0_u0_U59 (.B2( u1_u0_u0_n107 ) , .ZN( u1_u0_u0_n124 ) , .B1( u1_u0_u0_n128 ) , .A( u1_u0_u0_n161 ) );
  OAI21_X1 u1_u0_u0_U6 (.B1( u1_u0_u0_n150 ) , .B2( u1_u0_u0_n158 ) , .A( u1_u0_u0_n172 ) , .ZN( u1_u0_u0_n89 ) );
  INV_X1 u1_u0_u0_U60 (.A( u1_u0_u0_n111 ) , .ZN( u1_u0_u0_n170 ) );
  OR4_X1 u1_u0_u0_U61 (.ZN( u1_out0_31 ) , .A4( u1_u0_u0_n155 ) , .A2( u1_u0_u0_n156 ) , .A1( u1_u0_u0_n157 ) , .A3( u1_u0_u0_n173 ) );
  AOI21_X1 u1_u0_u0_U62 (.A( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n139 ) , .B1( u1_u0_u0_n140 ) , .ZN( u1_u0_u0_n157 ) );
  AOI21_X1 u1_u0_u0_U63 (.B2( u1_u0_u0_n141 ) , .B1( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n156 ) , .A( u1_u0_u0_n161 ) );
  INV_X1 u1_u0_u0_U64 (.ZN( u1_u0_u0_n174 ) , .A( u1_u0_u0_n89 ) );
  AOI211_X1 u1_u0_u0_U65 (.B( u1_u0_u0_n104 ) , .A( u1_u0_u0_n105 ) , .ZN( u1_u0_u0_n106 ) , .C2( u1_u0_u0_n113 ) , .C1( u1_u0_u0_n160 ) );
  AOI211_X1 u1_u0_u0_U66 (.B( u1_u0_u0_n115 ) , .A( u1_u0_u0_n116 ) , .C2( u1_u0_u0_n117 ) , .C1( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n119 ) );
  NAND2_X1 u1_u0_u0_U67 (.A2( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n121 ) , .A1( u1_u0_u0_n93 ) );
  NAND2_X1 u1_u0_u0_U68 (.A1( u1_u0_u0_n101 ) , .A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n150 ) );
  NOR2_X1 u1_u0_u0_U69 (.A2( u1_u0_X_1 ) , .A1( u1_u0_X_2 ) , .ZN( u1_u0_u0_n92 ) );
  AOI21_X1 u1_u0_u0_U7 (.B1( u1_u0_u0_n114 ) , .ZN( u1_u0_u0_n115 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n161 ) );
  NAND2_X1 u1_u0_u0_U70 (.A2( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n139 ) );
  NOR2_X1 u1_u0_u0_U71 (.A2( u1_u0_X_1 ) , .ZN( u1_u0_u0_n101 ) , .A1( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U72 (.A( u1_u0_X_1 ) , .ZN( u1_u0_u0_n164 ) );
  NAND2_X1 u1_u0_u0_U73 (.A1( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n128 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U74 (.A1( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n129 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U75 (.ZN( u1_u0_u0_n148 ) , .A1( u1_u0_u0_n93 ) , .A2( u1_u0_u0_n95 ) );
  OAI221_X1 u1_u0_u0_U76 (.C1( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n122 ) , .B2( u1_u0_u0_n127 ) , .A( u1_u0_u0_n143 ) , .B1( u1_u0_u0_n144 ) , .C2( u1_u0_u0_n147 ) );
  NOR2_X1 u1_u0_u0_U77 (.A1( u1_u0_u0_n163 ) , .A2( u1_u0_u0_n164 ) , .ZN( u1_u0_u0_n95 ) );
  AOI21_X1 u1_u0_u0_U78 (.B1( u1_u0_u0_n132 ) , .ZN( u1_u0_u0_n133 ) , .A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n166 ) );
  OAI22_X1 u1_u0_u0_U79 (.ZN( u1_u0_u0_n105 ) , .A2( u1_u0_u0_n132 ) , .B1( u1_u0_u0_n146 ) , .A1( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n161 ) );
  AND2_X1 u1_u0_u0_U8 (.A1( u1_u0_u0_n114 ) , .A2( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n146 ) );
  NAND2_X1 u1_u0_u0_U80 (.ZN( u1_u0_u0_n110 ) , .A2( u1_u0_u0_n132 ) , .A1( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U81 (.A( u1_u0_u0_n119 ) , .ZN( u1_u0_u0_n167 ) );
  NAND2_X1 u1_u0_u0_U82 (.A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U83 (.A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U84 (.ZN( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n92 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U85 (.ZN( u1_u0_u0_n142 ) , .A1( u1_u0_u0_n94 ) , .A2( u1_u0_u0_n95 ) );
  NOR2_X1 u1_u0_u0_U86 (.A2( u1_u0_X_6 ) , .ZN( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n162 ) );
  NOR2_X1 u1_u0_u0_U87 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n94 ) );
  NAND3_X1 u1_u0_u0_U88 (.ZN( u1_out0_23 ) , .A3( u1_u0_u0_n137 ) , .A1( u1_u0_u0_n168 ) , .A2( u1_u0_u0_n171 ) );
  NAND3_X1 u1_u0_u0_U89 (.A3( u1_u0_u0_n127 ) , .A2( u1_u0_u0_n128 ) , .ZN( u1_u0_u0_n135 ) , .A1( u1_u0_u0_n150 ) );
  AND2_X1 u1_u0_u0_U9 (.A1( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n141 ) , .A2( u1_u0_u0_n150 ) );
  NAND3_X1 u1_u0_u0_U90 (.ZN( u1_u0_u0_n117 ) , .A3( u1_u0_u0_n132 ) , .A2( u1_u0_u0_n139 ) , .A1( u1_u0_u0_n148 ) );
  NAND3_X1 u1_u0_u0_U91 (.ZN( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n114 ) , .A3( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n149 ) );
  NAND3_X1 u1_u0_u0_U92 (.ZN( u1_out0_9 ) , .A3( u1_u0_u0_n106 ) , .A2( u1_u0_u0_n171 ) , .A1( u1_u0_u0_n174 ) );
  NAND3_X1 u1_u0_u0_U93 (.A2( u1_u0_u0_n128 ) , .A1( u1_u0_u0_n132 ) , .A3( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n97 ) );
  AOI21_X1 u1_u0_u1_U10 (.B2( u1_u0_u1_n155 ) , .B1( u1_u0_u1_n156 ) , .ZN( u1_u0_u1_n157 ) , .A( u1_u0_u1_n174 ) );
  NAND3_X1 u1_u0_u1_U100 (.ZN( u1_u0_u1_n113 ) , .A1( u1_u0_u1_n120 ) , .A3( u1_u0_u1_n133 ) , .A2( u1_u0_u1_n155 ) );
  NAND2_X1 u1_u0_u1_U11 (.ZN( u1_u0_u1_n140 ) , .A2( u1_u0_u1_n150 ) , .A1( u1_u0_u1_n155 ) );
  NAND2_X1 u1_u0_u1_U12 (.A1( u1_u0_u1_n131 ) , .ZN( u1_u0_u1_n147 ) , .A2( u1_u0_u1_n153 ) );
  AOI22_X1 u1_u0_u1_U13 (.B2( u1_u0_u1_n136 ) , .A2( u1_u0_u1_n137 ) , .ZN( u1_u0_u1_n143 ) , .A1( u1_u0_u1_n171 ) , .B1( u1_u0_u1_n173 ) );
  INV_X1 u1_u0_u1_U14 (.A( u1_u0_u1_n147 ) , .ZN( u1_u0_u1_n181 ) );
  INV_X1 u1_u0_u1_U15 (.A( u1_u0_u1_n139 ) , .ZN( u1_u0_u1_n174 ) );
  OR4_X1 u1_u0_u1_U16 (.A4( u1_u0_u1_n106 ) , .A3( u1_u0_u1_n107 ) , .ZN( u1_u0_u1_n108 ) , .A1( u1_u0_u1_n117 ) , .A2( u1_u0_u1_n184 ) );
  AOI21_X1 u1_u0_u1_U17 (.ZN( u1_u0_u1_n106 ) , .A( u1_u0_u1_n112 ) , .B1( u1_u0_u1_n154 ) , .B2( u1_u0_u1_n156 ) );
  AOI21_X1 u1_u0_u1_U18 (.ZN( u1_u0_u1_n107 ) , .B1( u1_u0_u1_n134 ) , .B2( u1_u0_u1_n149 ) , .A( u1_u0_u1_n174 ) );
  INV_X1 u1_u0_u1_U19 (.A( u1_u0_u1_n101 ) , .ZN( u1_u0_u1_n184 ) );
  INV_X1 u1_u0_u1_U20 (.A( u1_u0_u1_n112 ) , .ZN( u1_u0_u1_n171 ) );
  NAND2_X1 u1_u0_u1_U21 (.ZN( u1_u0_u1_n141 ) , .A1( u1_u0_u1_n153 ) , .A2( u1_u0_u1_n156 ) );
  AND2_X1 u1_u0_u1_U22 (.A1( u1_u0_u1_n123 ) , .ZN( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n161 ) );
  NAND2_X1 u1_u0_u1_U23 (.A2( u1_u0_u1_n115 ) , .A1( u1_u0_u1_n116 ) , .ZN( u1_u0_u1_n148 ) );
  NAND2_X1 u1_u0_u1_U24 (.A2( u1_u0_u1_n133 ) , .A1( u1_u0_u1_n135 ) , .ZN( u1_u0_u1_n159 ) );
  NAND2_X1 u1_u0_u1_U25 (.A2( u1_u0_u1_n115 ) , .A1( u1_u0_u1_n120 ) , .ZN( u1_u0_u1_n132 ) );
  INV_X1 u1_u0_u1_U26 (.A( u1_u0_u1_n154 ) , .ZN( u1_u0_u1_n178 ) );
  INV_X1 u1_u0_u1_U27 (.A( u1_u0_u1_n151 ) , .ZN( u1_u0_u1_n183 ) );
  AND2_X1 u1_u0_u1_U28 (.A1( u1_u0_u1_n129 ) , .A2( u1_u0_u1_n133 ) , .ZN( u1_u0_u1_n149 ) );
  INV_X1 u1_u0_u1_U29 (.A( u1_u0_u1_n131 ) , .ZN( u1_u0_u1_n180 ) );
  INV_X1 u1_u0_u1_U3 (.A( u1_u0_u1_n159 ) , .ZN( u1_u0_u1_n182 ) );
  AOI221_X1 u1_u0_u1_U30 (.B1( u1_u0_u1_n140 ) , .ZN( u1_u0_u1_n167 ) , .B2( u1_u0_u1_n172 ) , .C2( u1_u0_u1_n175 ) , .C1( u1_u0_u1_n178 ) , .A( u1_u0_u1_n188 ) );
  INV_X1 u1_u0_u1_U31 (.ZN( u1_u0_u1_n188 ) , .A( u1_u0_u1_n97 ) );
  AOI211_X1 u1_u0_u1_U32 (.A( u1_u0_u1_n118 ) , .C1( u1_u0_u1_n132 ) , .C2( u1_u0_u1_n139 ) , .B( u1_u0_u1_n96 ) , .ZN( u1_u0_u1_n97 ) );
  AOI21_X1 u1_u0_u1_U33 (.B2( u1_u0_u1_n121 ) , .B1( u1_u0_u1_n135 ) , .A( u1_u0_u1_n152 ) , .ZN( u1_u0_u1_n96 ) );
  OAI221_X1 u1_u0_u1_U34 (.A( u1_u0_u1_n119 ) , .C2( u1_u0_u1_n129 ) , .ZN( u1_u0_u1_n138 ) , .B2( u1_u0_u1_n152 ) , .C1( u1_u0_u1_n174 ) , .B1( u1_u0_u1_n187 ) );
  INV_X1 u1_u0_u1_U35 (.A( u1_u0_u1_n148 ) , .ZN( u1_u0_u1_n187 ) );
  AOI211_X1 u1_u0_u1_U36 (.B( u1_u0_u1_n117 ) , .A( u1_u0_u1_n118 ) , .ZN( u1_u0_u1_n119 ) , .C2( u1_u0_u1_n146 ) , .C1( u1_u0_u1_n159 ) );
  NOR2_X1 u1_u0_u1_U37 (.A1( u1_u0_u1_n168 ) , .A2( u1_u0_u1_n176 ) , .ZN( u1_u0_u1_n98 ) );
  AOI211_X1 u1_u0_u1_U38 (.B( u1_u0_u1_n162 ) , .A( u1_u0_u1_n163 ) , .C2( u1_u0_u1_n164 ) , .ZN( u1_u0_u1_n165 ) , .C1( u1_u0_u1_n171 ) );
  AOI21_X1 u1_u0_u1_U39 (.A( u1_u0_u1_n160 ) , .B2( u1_u0_u1_n161 ) , .ZN( u1_u0_u1_n162 ) , .B1( u1_u0_u1_n182 ) );
  AOI221_X1 u1_u0_u1_U4 (.A( u1_u0_u1_n138 ) , .C2( u1_u0_u1_n139 ) , .C1( u1_u0_u1_n140 ) , .B2( u1_u0_u1_n141 ) , .ZN( u1_u0_u1_n142 ) , .B1( u1_u0_u1_n175 ) );
  OR2_X1 u1_u0_u1_U40 (.A2( u1_u0_u1_n157 ) , .A1( u1_u0_u1_n158 ) , .ZN( u1_u0_u1_n163 ) );
  OAI21_X1 u1_u0_u1_U41 (.B2( u1_u0_u1_n123 ) , .ZN( u1_u0_u1_n145 ) , .B1( u1_u0_u1_n160 ) , .A( u1_u0_u1_n185 ) );
  INV_X1 u1_u0_u1_U42 (.A( u1_u0_u1_n122 ) , .ZN( u1_u0_u1_n185 ) );
  AOI21_X1 u1_u0_u1_U43 (.B2( u1_u0_u1_n120 ) , .B1( u1_u0_u1_n121 ) , .ZN( u1_u0_u1_n122 ) , .A( u1_u0_u1_n128 ) );
  NAND2_X1 u1_u0_u1_U44 (.A1( u1_u0_u1_n128 ) , .ZN( u1_u0_u1_n146 ) , .A2( u1_u0_u1_n160 ) );
  NAND2_X1 u1_u0_u1_U45 (.A2( u1_u0_u1_n112 ) , .ZN( u1_u0_u1_n139 ) , .A1( u1_u0_u1_n152 ) );
  NAND2_X1 u1_u0_u1_U46 (.A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n156 ) , .A2( u1_u0_u1_n99 ) );
  NOR2_X1 u1_u0_u1_U47 (.ZN( u1_u0_u1_n117 ) , .A1( u1_u0_u1_n121 ) , .A2( u1_u0_u1_n160 ) );
  AOI21_X1 u1_u0_u1_U48 (.A( u1_u0_u1_n128 ) , .B2( u1_u0_u1_n129 ) , .ZN( u1_u0_u1_n130 ) , .B1( u1_u0_u1_n150 ) );
  NAND2_X1 u1_u0_u1_U49 (.ZN( u1_u0_u1_n112 ) , .A1( u1_u0_u1_n169 ) , .A2( u1_u0_u1_n170 ) );
  AOI211_X1 u1_u0_u1_U5 (.ZN( u1_u0_u1_n124 ) , .A( u1_u0_u1_n138 ) , .C2( u1_u0_u1_n139 ) , .B( u1_u0_u1_n145 ) , .C1( u1_u0_u1_n147 ) );
  NAND2_X1 u1_u0_u1_U50 (.ZN( u1_u0_u1_n129 ) , .A2( u1_u0_u1_n95 ) , .A1( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U51 (.A1( u1_u0_u1_n102 ) , .ZN( u1_u0_u1_n154 ) , .A2( u1_u0_u1_n99 ) );
  NAND2_X1 u1_u0_u1_U52 (.A2( u1_u0_u1_n100 ) , .ZN( u1_u0_u1_n135 ) , .A1( u1_u0_u1_n99 ) );
  AOI21_X1 u1_u0_u1_U53 (.A( u1_u0_u1_n152 ) , .B2( u1_u0_u1_n153 ) , .B1( u1_u0_u1_n154 ) , .ZN( u1_u0_u1_n158 ) );
  INV_X1 u1_u0_u1_U54 (.A( u1_u0_u1_n160 ) , .ZN( u1_u0_u1_n175 ) );
  NAND2_X1 u1_u0_u1_U55 (.A1( u1_u0_u1_n100 ) , .ZN( u1_u0_u1_n116 ) , .A2( u1_u0_u1_n95 ) );
  NAND2_X1 u1_u0_u1_U56 (.A1( u1_u0_u1_n102 ) , .ZN( u1_u0_u1_n131 ) , .A2( u1_u0_u1_n95 ) );
  NAND2_X1 u1_u0_u1_U57 (.A2( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n121 ) , .A1( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U58 (.A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n153 ) , .A2( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U59 (.A2( u1_u0_u1_n104 ) , .A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n133 ) );
  AOI22_X1 u1_u0_u1_U6 (.B2( u1_u0_u1_n113 ) , .A2( u1_u0_u1_n114 ) , .ZN( u1_u0_u1_n125 ) , .A1( u1_u0_u1_n171 ) , .B1( u1_u0_u1_n173 ) );
  NAND2_X1 u1_u0_u1_U60 (.ZN( u1_u0_u1_n150 ) , .A2( u1_u0_u1_n98 ) , .A1( u1_u0_u1_n99 ) );
  NAND2_X1 u1_u0_u1_U61 (.A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n155 ) , .A2( u1_u0_u1_n95 ) );
  OAI21_X1 u1_u0_u1_U62 (.ZN( u1_u0_u1_n109 ) , .B1( u1_u0_u1_n129 ) , .B2( u1_u0_u1_n160 ) , .A( u1_u0_u1_n167 ) );
  NAND2_X1 u1_u0_u1_U63 (.A2( u1_u0_u1_n100 ) , .A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n120 ) );
  NAND2_X1 u1_u0_u1_U64 (.A1( u1_u0_u1_n102 ) , .A2( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n115 ) );
  NAND2_X1 u1_u0_u1_U65 (.A2( u1_u0_u1_n100 ) , .A1( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n151 ) );
  NAND2_X1 u1_u0_u1_U66 (.A2( u1_u0_u1_n103 ) , .A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n161 ) );
  INV_X1 u1_u0_u1_U67 (.A( u1_u0_u1_n152 ) , .ZN( u1_u0_u1_n173 ) );
  INV_X1 u1_u0_u1_U68 (.A( u1_u0_u1_n128 ) , .ZN( u1_u0_u1_n172 ) );
  NAND2_X1 u1_u0_u1_U69 (.A2( u1_u0_u1_n102 ) , .A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n123 ) );
  NAND2_X1 u1_u0_u1_U7 (.ZN( u1_u0_u1_n114 ) , .A1( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n156 ) );
  NOR2_X1 u1_u0_u1_U70 (.A2( u1_u0_X_7 ) , .A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n95 ) );
  NOR2_X1 u1_u0_u1_U71 (.A1( u1_u0_X_12 ) , .A2( u1_u0_X_9 ) , .ZN( u1_u0_u1_n100 ) );
  NOR2_X1 u1_u0_u1_U72 (.A2( u1_u0_X_8 ) , .A1( u1_u0_u1_n177 ) , .ZN( u1_u0_u1_n99 ) );
  NOR2_X1 u1_u0_u1_U73 (.A2( u1_u0_X_12 ) , .ZN( u1_u0_u1_n102 ) , .A1( u1_u0_u1_n176 ) );
  NOR2_X1 u1_u0_u1_U74 (.A2( u1_u0_X_9 ) , .ZN( u1_u0_u1_n105 ) , .A1( u1_u0_u1_n168 ) );
  NAND2_X1 u1_u0_u1_U75 (.A1( u1_u0_X_10 ) , .ZN( u1_u0_u1_n160 ) , .A2( u1_u0_u1_n169 ) );
  NAND2_X1 u1_u0_u1_U76 (.A2( u1_u0_X_10 ) , .A1( u1_u0_X_11 ) , .ZN( u1_u0_u1_n152 ) );
  NAND2_X1 u1_u0_u1_U77 (.A1( u1_u0_X_11 ) , .ZN( u1_u0_u1_n128 ) , .A2( u1_u0_u1_n170 ) );
  AND2_X1 u1_u0_u1_U78 (.A2( u1_u0_X_7 ) , .A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n104 ) );
  AND2_X1 u1_u0_u1_U79 (.A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n103 ) , .A2( u1_u0_u1_n177 ) );
  NOR2_X1 u1_u0_u1_U8 (.A1( u1_u0_u1_n112 ) , .A2( u1_u0_u1_n116 ) , .ZN( u1_u0_u1_n118 ) );
  INV_X1 u1_u0_u1_U80 (.A( u1_u0_X_10 ) , .ZN( u1_u0_u1_n170 ) );
  INV_X1 u1_u0_u1_U81 (.A( u1_u0_X_9 ) , .ZN( u1_u0_u1_n176 ) );
  INV_X1 u1_u0_u1_U82 (.A( u1_u0_X_11 ) , .ZN( u1_u0_u1_n169 ) );
  INV_X1 u1_u0_u1_U83 (.A( u1_u0_X_12 ) , .ZN( u1_u0_u1_n168 ) );
  INV_X1 u1_u0_u1_U84 (.A( u1_u0_X_7 ) , .ZN( u1_u0_u1_n177 ) );
  NAND4_X1 u1_u0_u1_U85 (.ZN( u1_out0_28 ) , .A4( u1_u0_u1_n124 ) , .A3( u1_u0_u1_n125 ) , .A2( u1_u0_u1_n126 ) , .A1( u1_u0_u1_n127 ) );
  OAI21_X1 u1_u0_u1_U86 (.ZN( u1_u0_u1_n127 ) , .B2( u1_u0_u1_n139 ) , .B1( u1_u0_u1_n175 ) , .A( u1_u0_u1_n183 ) );
  OAI21_X1 u1_u0_u1_U87 (.ZN( u1_u0_u1_n126 ) , .B2( u1_u0_u1_n140 ) , .A( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n178 ) );
  NAND4_X1 u1_u0_u1_U88 (.ZN( u1_out0_18 ) , .A4( u1_u0_u1_n165 ) , .A3( u1_u0_u1_n166 ) , .A1( u1_u0_u1_n167 ) , .A2( u1_u0_u1_n186 ) );
  AOI22_X1 u1_u0_u1_U89 (.B2( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n147 ) , .A2( u1_u0_u1_n148 ) , .ZN( u1_u0_u1_n166 ) , .A1( u1_u0_u1_n172 ) );
  OAI21_X1 u1_u0_u1_U9 (.ZN( u1_u0_u1_n101 ) , .B1( u1_u0_u1_n141 ) , .A( u1_u0_u1_n146 ) , .B2( u1_u0_u1_n183 ) );
  INV_X1 u1_u0_u1_U90 (.A( u1_u0_u1_n145 ) , .ZN( u1_u0_u1_n186 ) );
  NAND4_X1 u1_u0_u1_U91 (.ZN( u1_out0_2 ) , .A4( u1_u0_u1_n142 ) , .A3( u1_u0_u1_n143 ) , .A2( u1_u0_u1_n144 ) , .A1( u1_u0_u1_n179 ) );
  OAI21_X1 u1_u0_u1_U92 (.B2( u1_u0_u1_n132 ) , .ZN( u1_u0_u1_n144 ) , .A( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n180 ) );
  INV_X1 u1_u0_u1_U93 (.A( u1_u0_u1_n130 ) , .ZN( u1_u0_u1_n179 ) );
  OR4_X1 u1_u0_u1_U94 (.ZN( u1_out0_13 ) , .A4( u1_u0_u1_n108 ) , .A3( u1_u0_u1_n109 ) , .A2( u1_u0_u1_n110 ) , .A1( u1_u0_u1_n111 ) );
  AOI21_X1 u1_u0_u1_U95 (.ZN( u1_u0_u1_n111 ) , .A( u1_u0_u1_n128 ) , .B2( u1_u0_u1_n131 ) , .B1( u1_u0_u1_n135 ) );
  AOI21_X1 u1_u0_u1_U96 (.ZN( u1_u0_u1_n110 ) , .A( u1_u0_u1_n116 ) , .B1( u1_u0_u1_n152 ) , .B2( u1_u0_u1_n160 ) );
  NAND3_X1 u1_u0_u1_U97 (.A3( u1_u0_u1_n149 ) , .A2( u1_u0_u1_n150 ) , .A1( u1_u0_u1_n151 ) , .ZN( u1_u0_u1_n164 ) );
  NAND3_X1 u1_u0_u1_U98 (.A3( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n135 ) , .ZN( u1_u0_u1_n136 ) , .A1( u1_u0_u1_n151 ) );
  NAND3_X1 u1_u0_u1_U99 (.A1( u1_u0_u1_n133 ) , .ZN( u1_u0_u1_n137 ) , .A2( u1_u0_u1_n154 ) , .A3( u1_u0_u1_n181 ) );
  INV_X1 u1_u0_u5_U10 (.A( u1_u0_u5_n121 ) , .ZN( u1_u0_u5_n177 ) );
  NOR3_X1 u1_u0_u5_U100 (.A3( u1_u0_u5_n141 ) , .A1( u1_u0_u5_n142 ) , .ZN( u1_u0_u5_n143 ) , .A2( u1_u0_u5_n191 ) );
  NAND4_X1 u1_u0_u5_U101 (.ZN( u1_out0_4 ) , .A4( u1_u0_u5_n112 ) , .A2( u1_u0_u5_n113 ) , .A1( u1_u0_u5_n114 ) , .A3( u1_u0_u5_n195 ) );
  AOI211_X1 u1_u0_u5_U102 (.A( u1_u0_u5_n110 ) , .C1( u1_u0_u5_n111 ) , .ZN( u1_u0_u5_n112 ) , .B( u1_u0_u5_n118 ) , .C2( u1_u0_u5_n177 ) );
  AOI222_X1 u1_u0_u5_U103 (.ZN( u1_u0_u5_n113 ) , .A1( u1_u0_u5_n131 ) , .C1( u1_u0_u5_n148 ) , .B2( u1_u0_u5_n174 ) , .C2( u1_u0_u5_n178 ) , .A2( u1_u0_u5_n179 ) , .B1( u1_u0_u5_n99 ) );
  NAND3_X1 u1_u0_u5_U104 (.A2( u1_u0_u5_n154 ) , .A3( u1_u0_u5_n158 ) , .A1( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n99 ) );
  NOR2_X1 u1_u0_u5_U11 (.ZN( u1_u0_u5_n160 ) , .A2( u1_u0_u5_n173 ) , .A1( u1_u0_u5_n177 ) );
  INV_X1 u1_u0_u5_U12 (.A( u1_u0_u5_n150 ) , .ZN( u1_u0_u5_n174 ) );
  AOI21_X1 u1_u0_u5_U13 (.A( u1_u0_u5_n160 ) , .B2( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n162 ) , .B1( u1_u0_u5_n192 ) );
  INV_X1 u1_u0_u5_U14 (.A( u1_u0_u5_n159 ) , .ZN( u1_u0_u5_n192 ) );
  AOI21_X1 u1_u0_u5_U15 (.A( u1_u0_u5_n156 ) , .B2( u1_u0_u5_n157 ) , .B1( u1_u0_u5_n158 ) , .ZN( u1_u0_u5_n163 ) );
  AOI21_X1 u1_u0_u5_U16 (.B2( u1_u0_u5_n139 ) , .B1( u1_u0_u5_n140 ) , .ZN( u1_u0_u5_n141 ) , .A( u1_u0_u5_n150 ) );
  OAI21_X1 u1_u0_u5_U17 (.A( u1_u0_u5_n133 ) , .B2( u1_u0_u5_n134 ) , .B1( u1_u0_u5_n135 ) , .ZN( u1_u0_u5_n142 ) );
  OAI21_X1 u1_u0_u5_U18 (.ZN( u1_u0_u5_n133 ) , .B2( u1_u0_u5_n147 ) , .A( u1_u0_u5_n173 ) , .B1( u1_u0_u5_n188 ) );
  NAND2_X1 u1_u0_u5_U19 (.A2( u1_u0_u5_n119 ) , .A1( u1_u0_u5_n123 ) , .ZN( u1_u0_u5_n137 ) );
  INV_X1 u1_u0_u5_U20 (.A( u1_u0_u5_n155 ) , .ZN( u1_u0_u5_n194 ) );
  NAND2_X1 u1_u0_u5_U21 (.A1( u1_u0_u5_n121 ) , .ZN( u1_u0_u5_n132 ) , .A2( u1_u0_u5_n172 ) );
  NAND2_X1 u1_u0_u5_U22 (.A2( u1_u0_u5_n122 ) , .ZN( u1_u0_u5_n136 ) , .A1( u1_u0_u5_n154 ) );
  NAND2_X1 u1_u0_u5_U23 (.A2( u1_u0_u5_n119 ) , .A1( u1_u0_u5_n120 ) , .ZN( u1_u0_u5_n159 ) );
  INV_X1 u1_u0_u5_U24 (.A( u1_u0_u5_n156 ) , .ZN( u1_u0_u5_n175 ) );
  INV_X1 u1_u0_u5_U25 (.A( u1_u0_u5_n158 ) , .ZN( u1_u0_u5_n188 ) );
  INV_X1 u1_u0_u5_U26 (.A( u1_u0_u5_n152 ) , .ZN( u1_u0_u5_n179 ) );
  INV_X1 u1_u0_u5_U27 (.A( u1_u0_u5_n140 ) , .ZN( u1_u0_u5_n182 ) );
  INV_X1 u1_u0_u5_U28 (.A( u1_u0_u5_n151 ) , .ZN( u1_u0_u5_n183 ) );
  INV_X1 u1_u0_u5_U29 (.A( u1_u0_u5_n123 ) , .ZN( u1_u0_u5_n185 ) );
  NOR2_X1 u1_u0_u5_U3 (.ZN( u1_u0_u5_n134 ) , .A1( u1_u0_u5_n183 ) , .A2( u1_u0_u5_n190 ) );
  INV_X1 u1_u0_u5_U30 (.A( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n184 ) );
  INV_X1 u1_u0_u5_U31 (.A( u1_u0_u5_n139 ) , .ZN( u1_u0_u5_n189 ) );
  INV_X1 u1_u0_u5_U32 (.A( u1_u0_u5_n157 ) , .ZN( u1_u0_u5_n190 ) );
  INV_X1 u1_u0_u5_U33 (.A( u1_u0_u5_n120 ) , .ZN( u1_u0_u5_n193 ) );
  NAND2_X1 u1_u0_u5_U34 (.ZN( u1_u0_u5_n111 ) , .A1( u1_u0_u5_n140 ) , .A2( u1_u0_u5_n155 ) );
  INV_X1 u1_u0_u5_U35 (.A( u1_u0_u5_n117 ) , .ZN( u1_u0_u5_n196 ) );
  OAI221_X1 u1_u0_u5_U36 (.A( u1_u0_u5_n116 ) , .ZN( u1_u0_u5_n117 ) , .B2( u1_u0_u5_n119 ) , .C1( u1_u0_u5_n153 ) , .C2( u1_u0_u5_n158 ) , .B1( u1_u0_u5_n172 ) );
  AOI222_X1 u1_u0_u5_U37 (.ZN( u1_u0_u5_n116 ) , .B2( u1_u0_u5_n145 ) , .C1( u1_u0_u5_n148 ) , .A2( u1_u0_u5_n174 ) , .C2( u1_u0_u5_n177 ) , .B1( u1_u0_u5_n187 ) , .A1( u1_u0_u5_n193 ) );
  INV_X1 u1_u0_u5_U38 (.A( u1_u0_u5_n115 ) , .ZN( u1_u0_u5_n187 ) );
  NOR2_X1 u1_u0_u5_U39 (.ZN( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n170 ) , .A2( u1_u0_u5_n180 ) );
  INV_X1 u1_u0_u5_U4 (.A( u1_u0_u5_n138 ) , .ZN( u1_u0_u5_n191 ) );
  AOI22_X1 u1_u0_u5_U40 (.B2( u1_u0_u5_n131 ) , .A2( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n169 ) , .B1( u1_u0_u5_n174 ) , .A1( u1_u0_u5_n185 ) );
  NOR2_X1 u1_u0_u5_U41 (.A1( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n150 ) , .A2( u1_u0_u5_n173 ) );
  AOI21_X1 u1_u0_u5_U42 (.A( u1_u0_u5_n118 ) , .B2( u1_u0_u5_n145 ) , .ZN( u1_u0_u5_n168 ) , .B1( u1_u0_u5_n186 ) );
  INV_X1 u1_u0_u5_U43 (.A( u1_u0_u5_n122 ) , .ZN( u1_u0_u5_n186 ) );
  NOR2_X1 u1_u0_u5_U44 (.A1( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n152 ) , .A2( u1_u0_u5_n176 ) );
  NOR2_X1 u1_u0_u5_U45 (.A1( u1_u0_u5_n115 ) , .ZN( u1_u0_u5_n118 ) , .A2( u1_u0_u5_n153 ) );
  NOR2_X1 u1_u0_u5_U46 (.A2( u1_u0_u5_n145 ) , .ZN( u1_u0_u5_n156 ) , .A1( u1_u0_u5_n174 ) );
  NOR2_X1 u1_u0_u5_U47 (.ZN( u1_u0_u5_n121 ) , .A2( u1_u0_u5_n145 ) , .A1( u1_u0_u5_n176 ) );
  AOI22_X1 u1_u0_u5_U48 (.ZN( u1_u0_u5_n114 ) , .A2( u1_u0_u5_n137 ) , .A1( u1_u0_u5_n145 ) , .B2( u1_u0_u5_n175 ) , .B1( u1_u0_u5_n193 ) );
  OAI211_X1 u1_u0_u5_U49 (.B( u1_u0_u5_n124 ) , .A( u1_u0_u5_n125 ) , .C2( u1_u0_u5_n126 ) , .C1( u1_u0_u5_n127 ) , .ZN( u1_u0_u5_n128 ) );
  OAI21_X1 u1_u0_u5_U5 (.B2( u1_u0_u5_n136 ) , .B1( u1_u0_u5_n137 ) , .ZN( u1_u0_u5_n138 ) , .A( u1_u0_u5_n177 ) );
  NOR3_X1 u1_u0_u5_U50 (.ZN( u1_u0_u5_n127 ) , .A1( u1_u0_u5_n136 ) , .A3( u1_u0_u5_n148 ) , .A2( u1_u0_u5_n182 ) );
  OAI21_X1 u1_u0_u5_U51 (.ZN( u1_u0_u5_n124 ) , .A( u1_u0_u5_n177 ) , .B2( u1_u0_u5_n183 ) , .B1( u1_u0_u5_n189 ) );
  OAI21_X1 u1_u0_u5_U52 (.ZN( u1_u0_u5_n125 ) , .A( u1_u0_u5_n174 ) , .B2( u1_u0_u5_n185 ) , .B1( u1_u0_u5_n190 ) );
  AOI21_X1 u1_u0_u5_U53 (.A( u1_u0_u5_n153 ) , .B2( u1_u0_u5_n154 ) , .B1( u1_u0_u5_n155 ) , .ZN( u1_u0_u5_n164 ) );
  AOI21_X1 u1_u0_u5_U54 (.ZN( u1_u0_u5_n110 ) , .B1( u1_u0_u5_n122 ) , .B2( u1_u0_u5_n139 ) , .A( u1_u0_u5_n153 ) );
  INV_X1 u1_u0_u5_U55 (.A( u1_u0_u5_n153 ) , .ZN( u1_u0_u5_n176 ) );
  INV_X1 u1_u0_u5_U56 (.A( u1_u0_u5_n126 ) , .ZN( u1_u0_u5_n173 ) );
  AND2_X1 u1_u0_u5_U57 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n147 ) );
  AND2_X1 u1_u0_u5_U58 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n148 ) );
  NAND2_X1 u1_u0_u5_U59 (.A1( u1_u0_u5_n105 ) , .A2( u1_u0_u5_n106 ) , .ZN( u1_u0_u5_n158 ) );
  INV_X1 u1_u0_u5_U6 (.A( u1_u0_u5_n135 ) , .ZN( u1_u0_u5_n178 ) );
  NAND2_X1 u1_u0_u5_U60 (.A2( u1_u0_u5_n108 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n139 ) );
  NAND2_X1 u1_u0_u5_U61 (.A1( u1_u0_u5_n106 ) , .A2( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n119 ) );
  NAND2_X1 u1_u0_u5_U62 (.A2( u1_u0_u5_n103 ) , .A1( u1_u0_u5_n105 ) , .ZN( u1_u0_u5_n140 ) );
  NAND2_X1 u1_u0_u5_U63 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n105 ) , .ZN( u1_u0_u5_n155 ) );
  NAND2_X1 u1_u0_u5_U64 (.A2( u1_u0_u5_n106 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n122 ) );
  NAND2_X1 u1_u0_u5_U65 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n106 ) , .ZN( u1_u0_u5_n115 ) );
  NAND2_X1 u1_u0_u5_U66 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n103 ) , .ZN( u1_u0_u5_n161 ) );
  NAND2_X1 u1_u0_u5_U67 (.A1( u1_u0_u5_n105 ) , .A2( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n154 ) );
  INV_X1 u1_u0_u5_U68 (.A( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n172 ) );
  NAND2_X1 u1_u0_u5_U69 (.A1( u1_u0_u5_n103 ) , .A2( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n123 ) );
  OAI22_X1 u1_u0_u5_U7 (.B2( u1_u0_u5_n149 ) , .B1( u1_u0_u5_n150 ) , .A2( u1_u0_u5_n151 ) , .A1( u1_u0_u5_n152 ) , .ZN( u1_u0_u5_n165 ) );
  NAND2_X1 u1_u0_u5_U70 (.A2( u1_u0_u5_n103 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n151 ) );
  NAND2_X1 u1_u0_u5_U71 (.A2( u1_u0_u5_n107 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n120 ) );
  NAND2_X1 u1_u0_u5_U72 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n157 ) );
  AND2_X1 u1_u0_u5_U73 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n104 ) , .ZN( u1_u0_u5_n131 ) );
  INV_X1 u1_u0_u5_U74 (.A( u1_u0_u5_n102 ) , .ZN( u1_u0_u5_n195 ) );
  OAI221_X1 u1_u0_u5_U75 (.A( u1_u0_u5_n101 ) , .ZN( u1_u0_u5_n102 ) , .C2( u1_u0_u5_n115 ) , .C1( u1_u0_u5_n126 ) , .B1( u1_u0_u5_n134 ) , .B2( u1_u0_u5_n160 ) );
  OAI21_X1 u1_u0_u5_U76 (.ZN( u1_u0_u5_n101 ) , .B1( u1_u0_u5_n137 ) , .A( u1_u0_u5_n146 ) , .B2( u1_u0_u5_n147 ) );
  NOR2_X1 u1_u0_u5_U77 (.A2( u1_u0_X_34 ) , .A1( u1_u0_X_35 ) , .ZN( u1_u0_u5_n145 ) );
  NOR2_X1 u1_u0_u5_U78 (.A2( u1_u0_X_34 ) , .ZN( u1_u0_u5_n146 ) , .A1( u1_u0_u5_n171 ) );
  NOR2_X1 u1_u0_u5_U79 (.A2( u1_u0_X_31 ) , .A1( u1_u0_X_32 ) , .ZN( u1_u0_u5_n103 ) );
  NOR3_X1 u1_u0_u5_U8 (.A2( u1_u0_u5_n147 ) , .A1( u1_u0_u5_n148 ) , .ZN( u1_u0_u5_n149 ) , .A3( u1_u0_u5_n194 ) );
  NOR2_X1 u1_u0_u5_U80 (.A2( u1_u0_X_36 ) , .ZN( u1_u0_u5_n105 ) , .A1( u1_u0_u5_n180 ) );
  NOR2_X1 u1_u0_u5_U81 (.A2( u1_u0_X_33 ) , .ZN( u1_u0_u5_n108 ) , .A1( u1_u0_u5_n170 ) );
  NOR2_X1 u1_u0_u5_U82 (.A2( u1_u0_X_33 ) , .A1( u1_u0_X_36 ) , .ZN( u1_u0_u5_n107 ) );
  NOR2_X1 u1_u0_u5_U83 (.A2( u1_u0_X_31 ) , .ZN( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n181 ) );
  NAND2_X1 u1_u0_u5_U84 (.A2( u1_u0_X_34 ) , .A1( u1_u0_X_35 ) , .ZN( u1_u0_u5_n153 ) );
  NAND2_X1 u1_u0_u5_U85 (.A1( u1_u0_X_34 ) , .ZN( u1_u0_u5_n126 ) , .A2( u1_u0_u5_n171 ) );
  AND2_X1 u1_u0_u5_U86 (.A1( u1_u0_X_31 ) , .A2( u1_u0_X_32 ) , .ZN( u1_u0_u5_n106 ) );
  AND2_X1 u1_u0_u5_U87 (.A1( u1_u0_X_31 ) , .ZN( u1_u0_u5_n109 ) , .A2( u1_u0_u5_n181 ) );
  INV_X1 u1_u0_u5_U88 (.A( u1_u0_X_33 ) , .ZN( u1_u0_u5_n180 ) );
  INV_X1 u1_u0_u5_U89 (.A( u1_u0_X_35 ) , .ZN( u1_u0_u5_n171 ) );
  NOR2_X1 u1_u0_u5_U9 (.ZN( u1_u0_u5_n135 ) , .A1( u1_u0_u5_n173 ) , .A2( u1_u0_u5_n176 ) );
  INV_X1 u1_u0_u5_U90 (.A( u1_u0_X_36 ) , .ZN( u1_u0_u5_n170 ) );
  INV_X1 u1_u0_u5_U91 (.A( u1_u0_X_32 ) , .ZN( u1_u0_u5_n181 ) );
  NAND4_X1 u1_u0_u5_U92 (.ZN( u1_out0_29 ) , .A4( u1_u0_u5_n129 ) , .A3( u1_u0_u5_n130 ) , .A2( u1_u0_u5_n168 ) , .A1( u1_u0_u5_n196 ) );
  AOI221_X1 u1_u0_u5_U93 (.A( u1_u0_u5_n128 ) , .ZN( u1_u0_u5_n129 ) , .C2( u1_u0_u5_n132 ) , .B2( u1_u0_u5_n159 ) , .B1( u1_u0_u5_n176 ) , .C1( u1_u0_u5_n184 ) );
  AOI222_X1 u1_u0_u5_U94 (.ZN( u1_u0_u5_n130 ) , .A2( u1_u0_u5_n146 ) , .B1( u1_u0_u5_n147 ) , .C2( u1_u0_u5_n175 ) , .B2( u1_u0_u5_n179 ) , .A1( u1_u0_u5_n188 ) , .C1( u1_u0_u5_n194 ) );
  NAND4_X1 u1_u0_u5_U95 (.ZN( u1_out0_19 ) , .A4( u1_u0_u5_n166 ) , .A3( u1_u0_u5_n167 ) , .A2( u1_u0_u5_n168 ) , .A1( u1_u0_u5_n169 ) );
  AOI22_X1 u1_u0_u5_U96 (.B2( u1_u0_u5_n145 ) , .A2( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n167 ) , .B1( u1_u0_u5_n182 ) , .A1( u1_u0_u5_n189 ) );
  NOR4_X1 u1_u0_u5_U97 (.A4( u1_u0_u5_n162 ) , .A3( u1_u0_u5_n163 ) , .A2( u1_u0_u5_n164 ) , .A1( u1_u0_u5_n165 ) , .ZN( u1_u0_u5_n166 ) );
  NAND4_X1 u1_u0_u5_U98 (.ZN( u1_out0_11 ) , .A4( u1_u0_u5_n143 ) , .A3( u1_u0_u5_n144 ) , .A2( u1_u0_u5_n169 ) , .A1( u1_u0_u5_n196 ) );
  AOI22_X1 u1_u0_u5_U99 (.A2( u1_u0_u5_n132 ) , .ZN( u1_u0_u5_n144 ) , .B2( u1_u0_u5_n145 ) , .B1( u1_u0_u5_n184 ) , .A1( u1_u0_u5_n194 ) );
  AOI22_X1 u1_u0_u6_U10 (.A2( u1_u0_u6_n151 ) , .B2( u1_u0_u6_n161 ) , .A1( u1_u0_u6_n167 ) , .B1( u1_u0_u6_n170 ) , .ZN( u1_u0_u6_n89 ) );
  AOI21_X1 u1_u0_u6_U11 (.B1( u1_u0_u6_n107 ) , .B2( u1_u0_u6_n132 ) , .A( u1_u0_u6_n158 ) , .ZN( u1_u0_u6_n88 ) );
  AOI21_X1 u1_u0_u6_U12 (.B2( u1_u0_u6_n147 ) , .B1( u1_u0_u6_n148 ) , .ZN( u1_u0_u6_n149 ) , .A( u1_u0_u6_n158 ) );
  AOI21_X1 u1_u0_u6_U13 (.ZN( u1_u0_u6_n106 ) , .A( u1_u0_u6_n142 ) , .B2( u1_u0_u6_n159 ) , .B1( u1_u0_u6_n164 ) );
  INV_X1 u1_u0_u6_U14 (.A( u1_u0_u6_n155 ) , .ZN( u1_u0_u6_n161 ) );
  INV_X1 u1_u0_u6_U15 (.A( u1_u0_u6_n128 ) , .ZN( u1_u0_u6_n164 ) );
  NAND2_X1 u1_u0_u6_U16 (.ZN( u1_u0_u6_n110 ) , .A1( u1_u0_u6_n122 ) , .A2( u1_u0_u6_n129 ) );
  NAND2_X1 u1_u0_u6_U17 (.ZN( u1_u0_u6_n124 ) , .A2( u1_u0_u6_n146 ) , .A1( u1_u0_u6_n148 ) );
  INV_X1 u1_u0_u6_U18 (.A( u1_u0_u6_n132 ) , .ZN( u1_u0_u6_n171 ) );
  AND2_X1 u1_u0_u6_U19 (.A1( u1_u0_u6_n100 ) , .ZN( u1_u0_u6_n130 ) , .A2( u1_u0_u6_n147 ) );
  INV_X1 u1_u0_u6_U20 (.A( u1_u0_u6_n127 ) , .ZN( u1_u0_u6_n173 ) );
  INV_X1 u1_u0_u6_U21 (.A( u1_u0_u6_n121 ) , .ZN( u1_u0_u6_n167 ) );
  INV_X1 u1_u0_u6_U22 (.A( u1_u0_u6_n100 ) , .ZN( u1_u0_u6_n169 ) );
  INV_X1 u1_u0_u6_U23 (.A( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n170 ) );
  INV_X1 u1_u0_u6_U24 (.A( u1_u0_u6_n113 ) , .ZN( u1_u0_u6_n168 ) );
  AND2_X1 u1_u0_u6_U25 (.A1( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n119 ) , .ZN( u1_u0_u6_n133 ) );
  AND2_X1 u1_u0_u6_U26 (.A2( u1_u0_u6_n121 ) , .A1( u1_u0_u6_n122 ) , .ZN( u1_u0_u6_n131 ) );
  AND3_X1 u1_u0_u6_U27 (.ZN( u1_u0_u6_n120 ) , .A2( u1_u0_u6_n127 ) , .A1( u1_u0_u6_n132 ) , .A3( u1_u0_u6_n145 ) );
  INV_X1 u1_u0_u6_U28 (.A( u1_u0_u6_n146 ) , .ZN( u1_u0_u6_n163 ) );
  AOI222_X1 u1_u0_u6_U29 (.ZN( u1_u0_u6_n114 ) , .A1( u1_u0_u6_n118 ) , .A2( u1_u0_u6_n126 ) , .B2( u1_u0_u6_n151 ) , .C2( u1_u0_u6_n159 ) , .C1( u1_u0_u6_n168 ) , .B1( u1_u0_u6_n169 ) );
  INV_X1 u1_u0_u6_U3 (.A( u1_u0_u6_n110 ) , .ZN( u1_u0_u6_n166 ) );
  NOR2_X1 u1_u0_u6_U30 (.A1( u1_u0_u6_n162 ) , .A2( u1_u0_u6_n165 ) , .ZN( u1_u0_u6_n98 ) );
  AOI211_X1 u1_u0_u6_U31 (.B( u1_u0_u6_n134 ) , .A( u1_u0_u6_n135 ) , .C1( u1_u0_u6_n136 ) , .ZN( u1_u0_u6_n137 ) , .C2( u1_u0_u6_n151 ) );
  AOI21_X1 u1_u0_u6_U32 (.B2( u1_u0_u6_n132 ) , .B1( u1_u0_u6_n133 ) , .ZN( u1_u0_u6_n134 ) , .A( u1_u0_u6_n158 ) );
  NAND4_X1 u1_u0_u6_U33 (.A4( u1_u0_u6_n127 ) , .A3( u1_u0_u6_n128 ) , .A2( u1_u0_u6_n129 ) , .A1( u1_u0_u6_n130 ) , .ZN( u1_u0_u6_n136 ) );
  AOI21_X1 u1_u0_u6_U34 (.B1( u1_u0_u6_n131 ) , .ZN( u1_u0_u6_n135 ) , .A( u1_u0_u6_n144 ) , .B2( u1_u0_u6_n146 ) );
  NAND2_X1 u1_u0_u6_U35 (.A1( u1_u0_u6_n144 ) , .ZN( u1_u0_u6_n151 ) , .A2( u1_u0_u6_n158 ) );
  NAND2_X1 u1_u0_u6_U36 (.ZN( u1_u0_u6_n132 ) , .A1( u1_u0_u6_n91 ) , .A2( u1_u0_u6_n97 ) );
  AOI22_X1 u1_u0_u6_U37 (.B2( u1_u0_u6_n110 ) , .B1( u1_u0_u6_n111 ) , .A1( u1_u0_u6_n112 ) , .ZN( u1_u0_u6_n115 ) , .A2( u1_u0_u6_n161 ) );
  NAND4_X1 u1_u0_u6_U38 (.A3( u1_u0_u6_n109 ) , .ZN( u1_u0_u6_n112 ) , .A4( u1_u0_u6_n132 ) , .A2( u1_u0_u6_n147 ) , .A1( u1_u0_u6_n166 ) );
  NOR2_X1 u1_u0_u6_U39 (.ZN( u1_u0_u6_n109 ) , .A1( u1_u0_u6_n170 ) , .A2( u1_u0_u6_n173 ) );
  INV_X1 u1_u0_u6_U4 (.A( u1_u0_u6_n142 ) , .ZN( u1_u0_u6_n174 ) );
  NOR2_X1 u1_u0_u6_U40 (.A2( u1_u0_u6_n126 ) , .ZN( u1_u0_u6_n155 ) , .A1( u1_u0_u6_n160 ) );
  NAND2_X1 u1_u0_u6_U41 (.ZN( u1_u0_u6_n146 ) , .A2( u1_u0_u6_n94 ) , .A1( u1_u0_u6_n99 ) );
  AOI21_X1 u1_u0_u6_U42 (.A( u1_u0_u6_n144 ) , .B2( u1_u0_u6_n145 ) , .B1( u1_u0_u6_n146 ) , .ZN( u1_u0_u6_n150 ) );
  INV_X1 u1_u0_u6_U43 (.A( u1_u0_u6_n111 ) , .ZN( u1_u0_u6_n158 ) );
  NAND2_X1 u1_u0_u6_U44 (.ZN( u1_u0_u6_n127 ) , .A1( u1_u0_u6_n91 ) , .A2( u1_u0_u6_n92 ) );
  NAND2_X1 u1_u0_u6_U45 (.ZN( u1_u0_u6_n129 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n96 ) );
  INV_X1 u1_u0_u6_U46 (.A( u1_u0_u6_n144 ) , .ZN( u1_u0_u6_n159 ) );
  NAND2_X1 u1_u0_u6_U47 (.ZN( u1_u0_u6_n145 ) , .A2( u1_u0_u6_n97 ) , .A1( u1_u0_u6_n98 ) );
  NAND2_X1 u1_u0_u6_U48 (.ZN( u1_u0_u6_n148 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n94 ) );
  NAND2_X1 u1_u0_u6_U49 (.ZN( u1_u0_u6_n108 ) , .A2( u1_u0_u6_n139 ) , .A1( u1_u0_u6_n144 ) );
  NAND2_X1 u1_u0_u6_U5 (.A2( u1_u0_u6_n143 ) , .ZN( u1_u0_u6_n152 ) , .A1( u1_u0_u6_n166 ) );
  NAND2_X1 u1_u0_u6_U50 (.ZN( u1_u0_u6_n121 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n97 ) );
  NAND2_X1 u1_u0_u6_U51 (.ZN( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n95 ) );
  AND2_X1 u1_u0_u6_U52 (.ZN( u1_u0_u6_n118 ) , .A2( u1_u0_u6_n91 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U53 (.ZN( u1_u0_u6_n147 ) , .A2( u1_u0_u6_n98 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U54 (.ZN( u1_u0_u6_n128 ) , .A1( u1_u0_u6_n94 ) , .A2( u1_u0_u6_n96 ) );
  NAND2_X1 u1_u0_u6_U55 (.ZN( u1_u0_u6_n119 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U56 (.ZN( u1_u0_u6_n123 ) , .A2( u1_u0_u6_n91 ) , .A1( u1_u0_u6_n96 ) );
  NAND2_X1 u1_u0_u6_U57 (.ZN( u1_u0_u6_n100 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n98 ) );
  NAND2_X1 u1_u0_u6_U58 (.ZN( u1_u0_u6_n122 ) , .A1( u1_u0_u6_n94 ) , .A2( u1_u0_u6_n97 ) );
  INV_X1 u1_u0_u6_U59 (.A( u1_u0_u6_n139 ) , .ZN( u1_u0_u6_n160 ) );
  AOI22_X1 u1_u0_u6_U6 (.B2( u1_u0_u6_n101 ) , .A1( u1_u0_u6_n102 ) , .ZN( u1_u0_u6_n103 ) , .B1( u1_u0_u6_n160 ) , .A2( u1_u0_u6_n161 ) );
  NAND2_X1 u1_u0_u6_U60 (.ZN( u1_u0_u6_n113 ) , .A1( u1_u0_u6_n96 ) , .A2( u1_u0_u6_n98 ) );
  NOR2_X1 u1_u0_u6_U61 (.A2( u1_u0_X_40 ) , .A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n126 ) );
  NOR2_X1 u1_u0_u6_U62 (.A2( u1_u0_X_39 ) , .A1( u1_u0_X_42 ) , .ZN( u1_u0_u6_n92 ) );
  NOR2_X1 u1_u0_u6_U63 (.A2( u1_u0_X_39 ) , .A1( u1_u0_u6_n156 ) , .ZN( u1_u0_u6_n97 ) );
  NOR2_X1 u1_u0_u6_U64 (.A2( u1_u0_X_38 ) , .A1( u1_u0_u6_n165 ) , .ZN( u1_u0_u6_n95 ) );
  NOR2_X1 u1_u0_u6_U65 (.A2( u1_u0_X_41 ) , .ZN( u1_u0_u6_n111 ) , .A1( u1_u0_u6_n157 ) );
  NOR2_X1 u1_u0_u6_U66 (.A2( u1_u0_X_37 ) , .A1( u1_u0_u6_n162 ) , .ZN( u1_u0_u6_n94 ) );
  NOR2_X1 u1_u0_u6_U67 (.A2( u1_u0_X_37 ) , .A1( u1_u0_X_38 ) , .ZN( u1_u0_u6_n91 ) );
  NAND2_X1 u1_u0_u6_U68 (.A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n144 ) , .A2( u1_u0_u6_n157 ) );
  NAND2_X1 u1_u0_u6_U69 (.A2( u1_u0_X_40 ) , .A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n139 ) );
  NOR2_X1 u1_u0_u6_U7 (.A1( u1_u0_u6_n118 ) , .ZN( u1_u0_u6_n143 ) , .A2( u1_u0_u6_n168 ) );
  AND2_X1 u1_u0_u6_U70 (.A1( u1_u0_X_39 ) , .A2( u1_u0_u6_n156 ) , .ZN( u1_u0_u6_n96 ) );
  AND2_X1 u1_u0_u6_U71 (.A1( u1_u0_X_39 ) , .A2( u1_u0_X_42 ) , .ZN( u1_u0_u6_n99 ) );
  INV_X1 u1_u0_u6_U72 (.A( u1_u0_X_40 ) , .ZN( u1_u0_u6_n157 ) );
  INV_X1 u1_u0_u6_U73 (.A( u1_u0_X_37 ) , .ZN( u1_u0_u6_n165 ) );
  INV_X1 u1_u0_u6_U74 (.A( u1_u0_X_38 ) , .ZN( u1_u0_u6_n162 ) );
  INV_X1 u1_u0_u6_U75 (.A( u1_u0_X_42 ) , .ZN( u1_u0_u6_n156 ) );
  NAND4_X1 u1_u0_u6_U76 (.ZN( u1_out0_32 ) , .A4( u1_u0_u6_n103 ) , .A3( u1_u0_u6_n104 ) , .A2( u1_u0_u6_n105 ) , .A1( u1_u0_u6_n106 ) );
  AOI22_X1 u1_u0_u6_U77 (.ZN( u1_u0_u6_n105 ) , .A2( u1_u0_u6_n108 ) , .A1( u1_u0_u6_n118 ) , .B2( u1_u0_u6_n126 ) , .B1( u1_u0_u6_n171 ) );
  AOI22_X1 u1_u0_u6_U78 (.ZN( u1_u0_u6_n104 ) , .A1( u1_u0_u6_n111 ) , .B1( u1_u0_u6_n124 ) , .B2( u1_u0_u6_n151 ) , .A2( u1_u0_u6_n93 ) );
  NAND4_X1 u1_u0_u6_U79 (.ZN( u1_out0_12 ) , .A4( u1_u0_u6_n114 ) , .A3( u1_u0_u6_n115 ) , .A2( u1_u0_u6_n116 ) , .A1( u1_u0_u6_n117 ) );
  OAI21_X1 u1_u0_u6_U8 (.A( u1_u0_u6_n159 ) , .B1( u1_u0_u6_n169 ) , .B2( u1_u0_u6_n173 ) , .ZN( u1_u0_u6_n90 ) );
  OAI22_X1 u1_u0_u6_U80 (.B2( u1_u0_u6_n111 ) , .ZN( u1_u0_u6_n116 ) , .B1( u1_u0_u6_n126 ) , .A2( u1_u0_u6_n164 ) , .A1( u1_u0_u6_n167 ) );
  OAI21_X1 u1_u0_u6_U81 (.A( u1_u0_u6_n108 ) , .ZN( u1_u0_u6_n117 ) , .B2( u1_u0_u6_n141 ) , .B1( u1_u0_u6_n163 ) );
  OAI211_X1 u1_u0_u6_U82 (.ZN( u1_out0_7 ) , .B( u1_u0_u6_n153 ) , .C2( u1_u0_u6_n154 ) , .C1( u1_u0_u6_n155 ) , .A( u1_u0_u6_n174 ) );
  NOR3_X1 u1_u0_u6_U83 (.A1( u1_u0_u6_n141 ) , .ZN( u1_u0_u6_n154 ) , .A3( u1_u0_u6_n164 ) , .A2( u1_u0_u6_n171 ) );
  AOI211_X1 u1_u0_u6_U84 (.B( u1_u0_u6_n149 ) , .A( u1_u0_u6_n150 ) , .C2( u1_u0_u6_n151 ) , .C1( u1_u0_u6_n152 ) , .ZN( u1_u0_u6_n153 ) );
  OAI211_X1 u1_u0_u6_U85 (.ZN( u1_out0_22 ) , .B( u1_u0_u6_n137 ) , .A( u1_u0_u6_n138 ) , .C2( u1_u0_u6_n139 ) , .C1( u1_u0_u6_n140 ) );
  AOI22_X1 u1_u0_u6_U86 (.B1( u1_u0_u6_n124 ) , .A2( u1_u0_u6_n125 ) , .A1( u1_u0_u6_n126 ) , .ZN( u1_u0_u6_n138 ) , .B2( u1_u0_u6_n161 ) );
  AND4_X1 u1_u0_u6_U87 (.A3( u1_u0_u6_n119 ) , .A1( u1_u0_u6_n120 ) , .A4( u1_u0_u6_n129 ) , .ZN( u1_u0_u6_n140 ) , .A2( u1_u0_u6_n143 ) );
  NAND3_X1 u1_u0_u6_U88 (.A2( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n125 ) , .A1( u1_u0_u6_n130 ) , .A3( u1_u0_u6_n131 ) );
  NAND3_X1 u1_u0_u6_U89 (.A3( u1_u0_u6_n133 ) , .ZN( u1_u0_u6_n141 ) , .A1( u1_u0_u6_n145 ) , .A2( u1_u0_u6_n148 ) );
  INV_X1 u1_u0_u6_U9 (.ZN( u1_u0_u6_n172 ) , .A( u1_u0_u6_n88 ) );
  NAND3_X1 u1_u0_u6_U90 (.ZN( u1_u0_u6_n101 ) , .A3( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n121 ) , .A1( u1_u0_u6_n127 ) );
  NAND3_X1 u1_u0_u6_U91 (.ZN( u1_u0_u6_n102 ) , .A3( u1_u0_u6_n130 ) , .A2( u1_u0_u6_n145 ) , .A1( u1_u0_u6_n166 ) );
  NAND3_X1 u1_u0_u6_U92 (.A3( u1_u0_u6_n113 ) , .A1( u1_u0_u6_n119 ) , .A2( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n93 ) );
  NAND3_X1 u1_u0_u6_U93 (.ZN( u1_u0_u6_n142 ) , .A2( u1_u0_u6_n172 ) , .A3( u1_u0_u6_n89 ) , .A1( u1_u0_u6_n90 ) );
  OAI21_X1 u1_u0_u7_U10 (.A( u1_u0_u7_n161 ) , .B1( u1_u0_u7_n168 ) , .B2( u1_u0_u7_n173 ) , .ZN( u1_u0_u7_n91 ) );
  AOI211_X1 u1_u0_u7_U11 (.A( u1_u0_u7_n117 ) , .ZN( u1_u0_u7_n118 ) , .C2( u1_u0_u7_n126 ) , .C1( u1_u0_u7_n177 ) , .B( u1_u0_u7_n180 ) );
  OAI22_X1 u1_u0_u7_U12 (.B1( u1_u0_u7_n115 ) , .ZN( u1_u0_u7_n117 ) , .A2( u1_u0_u7_n133 ) , .A1( u1_u0_u7_n137 ) , .B2( u1_u0_u7_n162 ) );
  INV_X1 u1_u0_u7_U13 (.A( u1_u0_u7_n116 ) , .ZN( u1_u0_u7_n180 ) );
  NOR3_X1 u1_u0_u7_U14 (.ZN( u1_u0_u7_n115 ) , .A3( u1_u0_u7_n145 ) , .A2( u1_u0_u7_n168 ) , .A1( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U15 (.A( u1_u0_u7_n133 ) , .ZN( u1_u0_u7_n176 ) );
  NOR3_X1 u1_u0_u7_U16 (.A2( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n135 ) , .ZN( u1_u0_u7_n136 ) , .A3( u1_u0_u7_n171 ) );
  NOR2_X1 u1_u0_u7_U17 (.A1( u1_u0_u7_n130 ) , .A2( u1_u0_u7_n134 ) , .ZN( u1_u0_u7_n153 ) );
  AOI21_X1 u1_u0_u7_U18 (.ZN( u1_u0_u7_n104 ) , .B2( u1_u0_u7_n112 ) , .B1( u1_u0_u7_n127 ) , .A( u1_u0_u7_n164 ) );
  AOI21_X1 u1_u0_u7_U19 (.ZN( u1_u0_u7_n106 ) , .B1( u1_u0_u7_n133 ) , .B2( u1_u0_u7_n146 ) , .A( u1_u0_u7_n162 ) );
  AOI21_X1 u1_u0_u7_U20 (.A( u1_u0_u7_n101 ) , .ZN( u1_u0_u7_n107 ) , .B2( u1_u0_u7_n128 ) , .B1( u1_u0_u7_n175 ) );
  INV_X1 u1_u0_u7_U21 (.A( u1_u0_u7_n101 ) , .ZN( u1_u0_u7_n165 ) );
  NOR2_X1 u1_u0_u7_U22 (.ZN( u1_u0_u7_n111 ) , .A2( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U23 (.A( u1_u0_u7_n138 ) , .ZN( u1_u0_u7_n171 ) );
  INV_X1 u1_u0_u7_U24 (.A( u1_u0_u7_n131 ) , .ZN( u1_u0_u7_n177 ) );
  INV_X1 u1_u0_u7_U25 (.A( u1_u0_u7_n110 ) , .ZN( u1_u0_u7_n174 ) );
  NAND2_X1 u1_u0_u7_U26 (.A1( u1_u0_u7_n129 ) , .A2( u1_u0_u7_n132 ) , .ZN( u1_u0_u7_n149 ) );
  NAND2_X1 u1_u0_u7_U27 (.A1( u1_u0_u7_n113 ) , .A2( u1_u0_u7_n124 ) , .ZN( u1_u0_u7_n130 ) );
  INV_X1 u1_u0_u7_U28 (.A( u1_u0_u7_n112 ) , .ZN( u1_u0_u7_n173 ) );
  INV_X1 u1_u0_u7_U29 (.A( u1_u0_u7_n128 ) , .ZN( u1_u0_u7_n168 ) );
  OAI21_X1 u1_u0_u7_U3 (.ZN( u1_u0_u7_n159 ) , .A( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n171 ) , .B1( u1_u0_u7_n174 ) );
  INV_X1 u1_u0_u7_U30 (.A( u1_u0_u7_n148 ) , .ZN( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U31 (.A( u1_u0_u7_n127 ) , .ZN( u1_u0_u7_n179 ) );
  INV_X1 u1_u0_u7_U32 (.A( u1_u0_u7_n153 ) , .ZN( u1_u0_u7_n172 ) );
  NOR2_X1 u1_u0_u7_U33 (.ZN( u1_u0_u7_n101 ) , .A2( u1_u0_u7_n150 ) , .A1( u1_u0_u7_n156 ) );
  AOI211_X1 u1_u0_u7_U34 (.B( u1_u0_u7_n139 ) , .A( u1_u0_u7_n140 ) , .C2( u1_u0_u7_n141 ) , .ZN( u1_u0_u7_n142 ) , .C1( u1_u0_u7_n156 ) );
  NAND4_X1 u1_u0_u7_U35 (.A3( u1_u0_u7_n127 ) , .A2( u1_u0_u7_n128 ) , .A1( u1_u0_u7_n129 ) , .ZN( u1_u0_u7_n141 ) , .A4( u1_u0_u7_n147 ) );
  AOI21_X1 u1_u0_u7_U36 (.A( u1_u0_u7_n137 ) , .B1( u1_u0_u7_n138 ) , .ZN( u1_u0_u7_n139 ) , .B2( u1_u0_u7_n146 ) );
  OAI22_X1 u1_u0_u7_U37 (.B1( u1_u0_u7_n136 ) , .ZN( u1_u0_u7_n140 ) , .A1( u1_u0_u7_n153 ) , .B2( u1_u0_u7_n162 ) , .A2( u1_u0_u7_n164 ) );
  INV_X1 u1_u0_u7_U38 (.A( u1_u0_u7_n125 ) , .ZN( u1_u0_u7_n161 ) );
  AOI21_X1 u1_u0_u7_U39 (.ZN( u1_u0_u7_n123 ) , .B1( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n177 ) , .A( u1_u0_u7_n97 ) );
  INV_X1 u1_u0_u7_U4 (.A( u1_u0_u7_n149 ) , .ZN( u1_u0_u7_n175 ) );
  AOI21_X1 u1_u0_u7_U40 (.B2( u1_u0_u7_n113 ) , .B1( u1_u0_u7_n124 ) , .A( u1_u0_u7_n125 ) , .ZN( u1_u0_u7_n97 ) );
  INV_X1 u1_u0_u7_U41 (.A( u1_u0_u7_n152 ) , .ZN( u1_u0_u7_n162 ) );
  AOI22_X1 u1_u0_u7_U42 (.A2( u1_u0_u7_n114 ) , .ZN( u1_u0_u7_n119 ) , .B1( u1_u0_u7_n130 ) , .A1( u1_u0_u7_n156 ) , .B2( u1_u0_u7_n165 ) );
  NAND2_X1 u1_u0_u7_U43 (.A2( u1_u0_u7_n112 ) , .ZN( u1_u0_u7_n114 ) , .A1( u1_u0_u7_n175 ) );
  NOR2_X1 u1_u0_u7_U44 (.ZN( u1_u0_u7_n137 ) , .A1( u1_u0_u7_n150 ) , .A2( u1_u0_u7_n161 ) );
  AND2_X1 u1_u0_u7_U45 (.ZN( u1_u0_u7_n145 ) , .A2( u1_u0_u7_n98 ) , .A1( u1_u0_u7_n99 ) );
  AOI21_X1 u1_u0_u7_U46 (.ZN( u1_u0_u7_n105 ) , .B2( u1_u0_u7_n110 ) , .A( u1_u0_u7_n125 ) , .B1( u1_u0_u7_n147 ) );
  NAND2_X1 u1_u0_u7_U47 (.ZN( u1_u0_u7_n146 ) , .A1( u1_u0_u7_n95 ) , .A2( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U48 (.A2( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n147 ) , .A1( u1_u0_u7_n93 ) );
  NAND2_X1 u1_u0_u7_U49 (.A1( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n127 ) , .A2( u1_u0_u7_n99 ) );
  INV_X1 u1_u0_u7_U5 (.A( u1_u0_u7_n154 ) , .ZN( u1_u0_u7_n178 ) );
  NAND2_X1 u1_u0_u7_U50 (.A2( u1_u0_u7_n102 ) , .A1( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n133 ) );
  OR2_X1 u1_u0_u7_U51 (.ZN( u1_u0_u7_n126 ) , .A2( u1_u0_u7_n152 ) , .A1( u1_u0_u7_n156 ) );
  NAND2_X1 u1_u0_u7_U52 (.ZN( u1_u0_u7_n112 ) , .A2( u1_u0_u7_n96 ) , .A1( u1_u0_u7_n99 ) );
  NAND2_X1 u1_u0_u7_U53 (.A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n128 ) , .A1( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U54 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n113 ) , .A2( u1_u0_u7_n93 ) );
  NAND2_X1 u1_u0_u7_U55 (.ZN( u1_u0_u7_n110 ) , .A1( u1_u0_u7_n95 ) , .A2( u1_u0_u7_n96 ) );
  INV_X1 u1_u0_u7_U56 (.A( u1_u0_u7_n150 ) , .ZN( u1_u0_u7_n164 ) );
  AND2_X1 u1_u0_u7_U57 (.ZN( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n93 ) , .A2( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U58 (.A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n124 ) , .A1( u1_u0_u7_n96 ) );
  NAND2_X1 u1_u0_u7_U59 (.A1( u1_u0_u7_n100 ) , .A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n129 ) );
  AOI211_X1 u1_u0_u7_U6 (.ZN( u1_u0_u7_n116 ) , .A( u1_u0_u7_n155 ) , .C1( u1_u0_u7_n161 ) , .C2( u1_u0_u7_n171 ) , .B( u1_u0_u7_n94 ) );
  NAND2_X1 u1_u0_u7_U60 (.A2( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n131 ) , .A1( u1_u0_u7_n95 ) );
  NAND2_X1 u1_u0_u7_U61 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n138 ) , .A2( u1_u0_u7_n99 ) );
  NAND2_X1 u1_u0_u7_U62 (.ZN( u1_u0_u7_n132 ) , .A1( u1_u0_u7_n93 ) , .A2( u1_u0_u7_n96 ) );
  NAND2_X1 u1_u0_u7_U63 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n148 ) , .A2( u1_u0_u7_n95 ) );
  NOR2_X1 u1_u0_u7_U64 (.A2( u1_u0_X_47 ) , .ZN( u1_u0_u7_n150 ) , .A1( u1_u0_u7_n163 ) );
  NOR2_X1 u1_u0_u7_U65 (.A2( u1_u0_X_43 ) , .A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n103 ) );
  NOR2_X1 u1_u0_u7_U66 (.A2( u1_u0_X_48 ) , .A1( u1_u0_u7_n166 ) , .ZN( u1_u0_u7_n95 ) );
  NOR2_X1 u1_u0_u7_U67 (.A2( u1_u0_X_45 ) , .A1( u1_u0_X_48 ) , .ZN( u1_u0_u7_n99 ) );
  NOR2_X1 u1_u0_u7_U68 (.A2( u1_u0_X_44 ) , .A1( u1_u0_u7_n167 ) , .ZN( u1_u0_u7_n98 ) );
  NOR2_X1 u1_u0_u7_U69 (.A2( u1_u0_X_46 ) , .A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n152 ) );
  OAI222_X1 u1_u0_u7_U7 (.C2( u1_u0_u7_n101 ) , .B2( u1_u0_u7_n111 ) , .A1( u1_u0_u7_n113 ) , .C1( u1_u0_u7_n146 ) , .A2( u1_u0_u7_n162 ) , .B1( u1_u0_u7_n164 ) , .ZN( u1_u0_u7_n94 ) );
  NAND2_X1 u1_u0_u7_U70 (.A2( u1_u0_X_46 ) , .A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n125 ) );
  AND2_X1 u1_u0_u7_U71 (.A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n156 ) , .A2( u1_u0_u7_n163 ) );
  AND2_X1 u1_u0_u7_U72 (.A2( u1_u0_X_45 ) , .A1( u1_u0_X_48 ) , .ZN( u1_u0_u7_n102 ) );
  AND2_X1 u1_u0_u7_U73 (.A2( u1_u0_X_43 ) , .A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n96 ) );
  AND2_X1 u1_u0_u7_U74 (.A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n100 ) , .A2( u1_u0_u7_n167 ) );
  AND2_X1 u1_u0_u7_U75 (.A1( u1_u0_X_48 ) , .A2( u1_u0_u7_n166 ) , .ZN( u1_u0_u7_n93 ) );
  INV_X1 u1_u0_u7_U76 (.A( u1_u0_X_46 ) , .ZN( u1_u0_u7_n163 ) );
  INV_X1 u1_u0_u7_U77 (.A( u1_u0_X_45 ) , .ZN( u1_u0_u7_n166 ) );
  NAND4_X1 u1_u0_u7_U78 (.ZN( u1_out0_5 ) , .A4( u1_u0_u7_n108 ) , .A3( u1_u0_u7_n109 ) , .A1( u1_u0_u7_n116 ) , .A2( u1_u0_u7_n123 ) );
  AOI22_X1 u1_u0_u7_U79 (.ZN( u1_u0_u7_n109 ) , .A2( u1_u0_u7_n126 ) , .B2( u1_u0_u7_n145 ) , .B1( u1_u0_u7_n156 ) , .A1( u1_u0_u7_n171 ) );
  OAI221_X1 u1_u0_u7_U8 (.C1( u1_u0_u7_n101 ) , .C2( u1_u0_u7_n147 ) , .ZN( u1_u0_u7_n155 ) , .B2( u1_u0_u7_n162 ) , .A( u1_u0_u7_n91 ) , .B1( u1_u0_u7_n92 ) );
  NOR4_X1 u1_u0_u7_U80 (.A4( u1_u0_u7_n104 ) , .A3( u1_u0_u7_n105 ) , .A2( u1_u0_u7_n106 ) , .A1( u1_u0_u7_n107 ) , .ZN( u1_u0_u7_n108 ) );
  NAND4_X1 u1_u0_u7_U81 (.ZN( u1_out0_27 ) , .A4( u1_u0_u7_n118 ) , .A3( u1_u0_u7_n119 ) , .A2( u1_u0_u7_n120 ) , .A1( u1_u0_u7_n121 ) );
  OAI21_X1 u1_u0_u7_U82 (.ZN( u1_u0_u7_n121 ) , .B2( u1_u0_u7_n145 ) , .A( u1_u0_u7_n150 ) , .B1( u1_u0_u7_n174 ) );
  OAI21_X1 u1_u0_u7_U83 (.ZN( u1_u0_u7_n120 ) , .A( u1_u0_u7_n161 ) , .B2( u1_u0_u7_n170 ) , .B1( u1_u0_u7_n179 ) );
  NAND4_X1 u1_u0_u7_U84 (.ZN( u1_out0_21 ) , .A4( u1_u0_u7_n157 ) , .A3( u1_u0_u7_n158 ) , .A2( u1_u0_u7_n159 ) , .A1( u1_u0_u7_n160 ) );
  OAI21_X1 u1_u0_u7_U85 (.B1( u1_u0_u7_n145 ) , .ZN( u1_u0_u7_n160 ) , .A( u1_u0_u7_n161 ) , .B2( u1_u0_u7_n177 ) );
  AOI22_X1 u1_u0_u7_U86 (.B2( u1_u0_u7_n149 ) , .B1( u1_u0_u7_n150 ) , .A2( u1_u0_u7_n151 ) , .A1( u1_u0_u7_n152 ) , .ZN( u1_u0_u7_n158 ) );
  NAND4_X1 u1_u0_u7_U87 (.ZN( u1_out0_15 ) , .A4( u1_u0_u7_n142 ) , .A3( u1_u0_u7_n143 ) , .A2( u1_u0_u7_n144 ) , .A1( u1_u0_u7_n178 ) );
  OR2_X1 u1_u0_u7_U88 (.A2( u1_u0_u7_n125 ) , .A1( u1_u0_u7_n129 ) , .ZN( u1_u0_u7_n144 ) );
  AOI22_X1 u1_u0_u7_U89 (.A2( u1_u0_u7_n126 ) , .ZN( u1_u0_u7_n143 ) , .B2( u1_u0_u7_n165 ) , .B1( u1_u0_u7_n173 ) , .A1( u1_u0_u7_n174 ) );
  AND3_X1 u1_u0_u7_U9 (.A3( u1_u0_u7_n110 ) , .A2( u1_u0_u7_n127 ) , .A1( u1_u0_u7_n132 ) , .ZN( u1_u0_u7_n92 ) );
  INV_X1 u1_u0_u7_U90 (.A( u1_u0_X_43 ) , .ZN( u1_u0_u7_n167 ) );
  AOI211_X1 u1_u0_u7_U91 (.B( u1_u0_u7_n154 ) , .A( u1_u0_u7_n155 ) , .C1( u1_u0_u7_n156 ) , .ZN( u1_u0_u7_n157 ) , .C2( u1_u0_u7_n172 ) );
  OAI211_X1 u1_u0_u7_U92 (.B( u1_u0_u7_n122 ) , .A( u1_u0_u7_n123 ) , .C2( u1_u0_u7_n124 ) , .ZN( u1_u0_u7_n154 ) , .C1( u1_u0_u7_n162 ) );
  AOI222_X1 u1_u0_u7_U93 (.ZN( u1_u0_u7_n122 ) , .C2( u1_u0_u7_n126 ) , .C1( u1_u0_u7_n145 ) , .B1( u1_u0_u7_n161 ) , .A2( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n170 ) , .A1( u1_u0_u7_n176 ) );
  INV_X1 u1_u0_u7_U94 (.A( u1_u0_u7_n111 ) , .ZN( u1_u0_u7_n170 ) );
  NAND3_X1 u1_u0_u7_U95 (.A3( u1_u0_u7_n146 ) , .A2( u1_u0_u7_n147 ) , .A1( u1_u0_u7_n148 ) , .ZN( u1_u0_u7_n151 ) );
  NAND3_X1 u1_u0_u7_U96 (.A3( u1_u0_u7_n131 ) , .A2( u1_u0_u7_n132 ) , .A1( u1_u0_u7_n133 ) , .ZN( u1_u0_u7_n135 ) );
  XOR2_X1 u1_u10_U18 (.B( u1_K11_38 ) , .A( u1_R9_25 ) , .Z( u1_u10_X_38 ) );
  XOR2_X1 u1_u10_U19 (.B( u1_K11_37 ) , .A( u1_R9_24 ) , .Z( u1_u10_X_37 ) );
  XOR2_X1 u1_u10_U20 (.B( u1_K11_36 ) , .A( u1_R9_25 ) , .Z( u1_u10_X_36 ) );
  XOR2_X1 u1_u10_U21 (.B( u1_K11_35 ) , .A( u1_R9_24 ) , .Z( u1_u10_X_35 ) );
  XOR2_X1 u1_u10_U22 (.B( u1_K11_34 ) , .A( u1_R9_23 ) , .Z( u1_u10_X_34 ) );
  XOR2_X1 u1_u10_U24 (.B( u1_K11_32 ) , .A( u1_R9_21 ) , .Z( u1_u10_X_32 ) );
  XOR2_X1 u1_u10_U25 (.B( u1_K11_31 ) , .A( u1_R9_20 ) , .Z( u1_u10_X_31 ) );
  XOR2_X1 u1_u10_U27 (.B( u1_K11_2 ) , .A( u1_R9_1 ) , .Z( u1_u10_X_2 ) );
  XOR2_X1 u1_u10_U3 (.B( u1_K11_7 ) , .A( u1_R9_4 ) , .Z( u1_u10_X_7 ) );
  XOR2_X1 u1_u10_U41 (.B( u1_K11_17 ) , .A( u1_R9_12 ) , .Z( u1_u10_X_17 ) );
  XOR2_X1 u1_u10_U44 (.B( u1_K11_14 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_14 ) );
  XOR2_X1 u1_u10_U45 (.B( u1_K11_13 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_13 ) );
  XOR2_X1 u1_u10_U46 (.B( u1_K11_12 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_12 ) );
  XOR2_X1 u1_u10_U47 (.B( u1_K11_11 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_11 ) );
  XOR2_X1 u1_u10_U5 (.B( u1_K11_5 ) , .A( u1_R9_4 ) , .Z( u1_u10_X_5 ) );
  XOR2_X1 u1_u10_U7 (.B( u1_K11_48 ) , .A( u1_R9_1 ) , .Z( u1_u10_X_48 ) );
  AND3_X1 u1_u10_u0_U10 (.A2( u1_u10_u0_n112 ) , .ZN( u1_u10_u0_n127 ) , .A3( u1_u10_u0_n130 ) , .A1( u1_u10_u0_n148 ) );
  NAND2_X1 u1_u10_u0_U11 (.ZN( u1_u10_u0_n113 ) , .A1( u1_u10_u0_n139 ) , .A2( u1_u10_u0_n149 ) );
  AND2_X1 u1_u10_u0_U12 (.ZN( u1_u10_u0_n107 ) , .A1( u1_u10_u0_n130 ) , .A2( u1_u10_u0_n140 ) );
  AND2_X1 u1_u10_u0_U13 (.A2( u1_u10_u0_n129 ) , .A1( u1_u10_u0_n130 ) , .ZN( u1_u10_u0_n151 ) );
  AND2_X1 u1_u10_u0_U14 (.A1( u1_u10_u0_n108 ) , .A2( u1_u10_u0_n125 ) , .ZN( u1_u10_u0_n145 ) );
  INV_X1 u1_u10_u0_U15 (.A( u1_u10_u0_n143 ) , .ZN( u1_u10_u0_n173 ) );
  NOR2_X1 u1_u10_u0_U16 (.A2( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n147 ) , .A1( u1_u10_u0_n160 ) );
  NOR2_X1 u1_u10_u0_U17 (.A1( u1_u10_u0_n163 ) , .A2( u1_u10_u0_n164 ) , .ZN( u1_u10_u0_n95 ) );
  AOI21_X1 u1_u10_u0_U18 (.B1( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n132 ) , .A( u1_u10_u0_n165 ) , .B2( u1_u10_u0_n93 ) );
  INV_X1 u1_u10_u0_U19 (.A( u1_u10_u0_n142 ) , .ZN( u1_u10_u0_n165 ) );
  OAI221_X1 u1_u10_u0_U20 (.C1( u1_u10_u0_n121 ) , .ZN( u1_u10_u0_n122 ) , .B2( u1_u10_u0_n127 ) , .A( u1_u10_u0_n143 ) , .B1( u1_u10_u0_n144 ) , .C2( u1_u10_u0_n147 ) );
  OAI22_X1 u1_u10_u0_U21 (.B1( u1_u10_u0_n125 ) , .ZN( u1_u10_u0_n126 ) , .A1( u1_u10_u0_n138 ) , .A2( u1_u10_u0_n146 ) , .B2( u1_u10_u0_n147 ) );
  OAI22_X1 u1_u10_u0_U22 (.B1( u1_u10_u0_n131 ) , .A1( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n147 ) , .A2( u1_u10_u0_n90 ) , .ZN( u1_u10_u0_n91 ) );
  AND3_X1 u1_u10_u0_U23 (.A3( u1_u10_u0_n121 ) , .A2( u1_u10_u0_n125 ) , .A1( u1_u10_u0_n148 ) , .ZN( u1_u10_u0_n90 ) );
  INV_X1 u1_u10_u0_U24 (.A( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n161 ) );
  NOR2_X1 u1_u10_u0_U25 (.A1( u1_u10_u0_n120 ) , .ZN( u1_u10_u0_n143 ) , .A2( u1_u10_u0_n167 ) );
  OAI221_X1 u1_u10_u0_U26 (.C1( u1_u10_u0_n112 ) , .ZN( u1_u10_u0_n120 ) , .B1( u1_u10_u0_n138 ) , .B2( u1_u10_u0_n141 ) , .C2( u1_u10_u0_n147 ) , .A( u1_u10_u0_n172 ) );
  AOI22_X1 u1_u10_u0_U27 (.B2( u1_u10_u0_n109 ) , .A2( u1_u10_u0_n110 ) , .ZN( u1_u10_u0_n111 ) , .B1( u1_u10_u0_n118 ) , .A1( u1_u10_u0_n160 ) );
  INV_X1 u1_u10_u0_U28 (.A( u1_u10_u0_n118 ) , .ZN( u1_u10_u0_n158 ) );
  AOI21_X1 u1_u10_u0_U29 (.B1( u1_u10_u0_n132 ) , .ZN( u1_u10_u0_n133 ) , .A( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n166 ) );
  INV_X1 u1_u10_u0_U3 (.A( u1_u10_u0_n113 ) , .ZN( u1_u10_u0_n166 ) );
  AOI21_X1 u1_u10_u0_U30 (.ZN( u1_u10_u0_n104 ) , .B1( u1_u10_u0_n107 ) , .B2( u1_u10_u0_n141 ) , .A( u1_u10_u0_n144 ) );
  AOI21_X1 u1_u10_u0_U31 (.B1( u1_u10_u0_n127 ) , .B2( u1_u10_u0_n129 ) , .A( u1_u10_u0_n138 ) , .ZN( u1_u10_u0_n96 ) );
  AOI21_X1 u1_u10_u0_U32 (.ZN( u1_u10_u0_n116 ) , .B2( u1_u10_u0_n142 ) , .A( u1_u10_u0_n144 ) , .B1( u1_u10_u0_n166 ) );
  NAND2_X1 u1_u10_u0_U33 (.A1( u1_u10_u0_n100 ) , .A2( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n125 ) );
  NAND2_X1 u1_u10_u0_U34 (.A2( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n140 ) , .A1( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U35 (.A1( u1_u10_u0_n101 ) , .A2( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n150 ) );
  INV_X1 u1_u10_u0_U36 (.A( u1_u10_u0_n138 ) , .ZN( u1_u10_u0_n160 ) );
  NAND2_X1 u1_u10_u0_U37 (.ZN( u1_u10_u0_n142 ) , .A1( u1_u10_u0_n94 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U38 (.A1( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n128 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U39 (.A2( u1_u10_u0_n102 ) , .A1( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n149 ) );
  AOI21_X1 u1_u10_u0_U4 (.B2( u1_u10_u0_n131 ) , .ZN( u1_u10_u0_n134 ) , .B1( u1_u10_u0_n151 ) , .A( u1_u10_u0_n158 ) );
  NAND2_X1 u1_u10_u0_U40 (.A1( u1_u10_u0_n100 ) , .ZN( u1_u10_u0_n129 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U41 (.A2( u1_u10_u0_n100 ) , .A1( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n139 ) );
  NAND2_X1 u1_u10_u0_U42 (.A2( u1_u10_u0_n100 ) , .ZN( u1_u10_u0_n131 ) , .A1( u1_u10_u0_n92 ) );
  NAND2_X1 u1_u10_u0_U43 (.ZN( u1_u10_u0_n108 ) , .A1( u1_u10_u0_n92 ) , .A2( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U44 (.ZN( u1_u10_u0_n148 ) , .A1( u1_u10_u0_n93 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U45 (.A2( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n114 ) , .A1( u1_u10_u0_n92 ) );
  NAND2_X1 u1_u10_u0_U46 (.A1( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n130 ) , .A2( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U47 (.A2( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n121 ) , .A1( u1_u10_u0_n93 ) );
  INV_X1 u1_u10_u0_U48 (.ZN( u1_u10_u0_n172 ) , .A( u1_u10_u0_n88 ) );
  OAI222_X1 u1_u10_u0_U49 (.C1( u1_u10_u0_n108 ) , .A1( u1_u10_u0_n125 ) , .B2( u1_u10_u0_n128 ) , .B1( u1_u10_u0_n144 ) , .A2( u1_u10_u0_n158 ) , .C2( u1_u10_u0_n161 ) , .ZN( u1_u10_u0_n88 ) );
  NOR2_X1 u1_u10_u0_U5 (.A1( u1_u10_u0_n108 ) , .ZN( u1_u10_u0_n123 ) , .A2( u1_u10_u0_n158 ) );
  NAND2_X1 u1_u10_u0_U50 (.ZN( u1_u10_u0_n112 ) , .A2( u1_u10_u0_n92 ) , .A1( u1_u10_u0_n93 ) );
  OR3_X1 u1_u10_u0_U51 (.A3( u1_u10_u0_n152 ) , .A2( u1_u10_u0_n153 ) , .A1( u1_u10_u0_n154 ) , .ZN( u1_u10_u0_n155 ) );
  AOI21_X1 u1_u10_u0_U52 (.A( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n145 ) , .B1( u1_u10_u0_n146 ) , .ZN( u1_u10_u0_n154 ) );
  AOI21_X1 u1_u10_u0_U53 (.B2( u1_u10_u0_n150 ) , .B1( u1_u10_u0_n151 ) , .ZN( u1_u10_u0_n152 ) , .A( u1_u10_u0_n158 ) );
  AOI21_X1 u1_u10_u0_U54 (.A( u1_u10_u0_n147 ) , .B2( u1_u10_u0_n148 ) , .B1( u1_u10_u0_n149 ) , .ZN( u1_u10_u0_n153 ) );
  INV_X1 u1_u10_u0_U55 (.ZN( u1_u10_u0_n171 ) , .A( u1_u10_u0_n99 ) );
  OAI211_X1 u1_u10_u0_U56 (.C2( u1_u10_u0_n140 ) , .C1( u1_u10_u0_n161 ) , .A( u1_u10_u0_n169 ) , .B( u1_u10_u0_n98 ) , .ZN( u1_u10_u0_n99 ) );
  INV_X1 u1_u10_u0_U57 (.ZN( u1_u10_u0_n169 ) , .A( u1_u10_u0_n91 ) );
  AOI211_X1 u1_u10_u0_U58 (.C1( u1_u10_u0_n118 ) , .A( u1_u10_u0_n123 ) , .B( u1_u10_u0_n96 ) , .C2( u1_u10_u0_n97 ) , .ZN( u1_u10_u0_n98 ) );
  NOR2_X1 u1_u10_u0_U59 (.A2( u1_u10_X_2 ) , .ZN( u1_u10_u0_n103 ) , .A1( u1_u10_u0_n164 ) );
  OAI21_X1 u1_u10_u0_U6 (.B1( u1_u10_u0_n150 ) , .B2( u1_u10_u0_n158 ) , .A( u1_u10_u0_n172 ) , .ZN( u1_u10_u0_n89 ) );
  NOR2_X1 u1_u10_u0_U60 (.A2( u1_u10_X_3 ) , .A1( u1_u10_X_6 ) , .ZN( u1_u10_u0_n94 ) );
  NOR2_X1 u1_u10_u0_U61 (.A2( u1_u10_X_6 ) , .ZN( u1_u10_u0_n100 ) , .A1( u1_u10_u0_n162 ) );
  NOR2_X1 u1_u10_u0_U62 (.A2( u1_u10_X_1 ) , .A1( u1_u10_X_2 ) , .ZN( u1_u10_u0_n92 ) );
  NOR2_X1 u1_u10_u0_U63 (.A2( u1_u10_X_1 ) , .ZN( u1_u10_u0_n101 ) , .A1( u1_u10_u0_n163 ) );
  NOR2_X1 u1_u10_u0_U64 (.A2( u1_u10_X_4 ) , .A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n118 ) );
  NAND2_X1 u1_u10_u0_U65 (.A2( u1_u10_X_4 ) , .A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n144 ) );
  NOR2_X1 u1_u10_u0_U66 (.A2( u1_u10_X_5 ) , .ZN( u1_u10_u0_n136 ) , .A1( u1_u10_u0_n159 ) );
  NAND2_X1 u1_u10_u0_U67 (.A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n138 ) , .A2( u1_u10_u0_n159 ) );
  AND2_X1 u1_u10_u0_U68 (.A2( u1_u10_X_3 ) , .A1( u1_u10_X_6 ) , .ZN( u1_u10_u0_n102 ) );
  AND2_X1 u1_u10_u0_U69 (.A1( u1_u10_X_6 ) , .A2( u1_u10_u0_n162 ) , .ZN( u1_u10_u0_n93 ) );
  AOI21_X1 u1_u10_u0_U7 (.B1( u1_u10_u0_n114 ) , .ZN( u1_u10_u0_n115 ) , .B2( u1_u10_u0_n129 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U70 (.A( u1_u10_X_4 ) , .ZN( u1_u10_u0_n159 ) );
  INV_X1 u1_u10_u0_U71 (.A( u1_u10_X_1 ) , .ZN( u1_u10_u0_n164 ) );
  INV_X1 u1_u10_u0_U72 (.A( u1_u10_X_2 ) , .ZN( u1_u10_u0_n163 ) );
  INV_X1 u1_u10_u0_U73 (.A( u1_u10_X_3 ) , .ZN( u1_u10_u0_n162 ) );
  INV_X1 u1_u10_u0_U74 (.ZN( u1_u10_u0_n174 ) , .A( u1_u10_u0_n89 ) );
  AOI211_X1 u1_u10_u0_U75 (.B( u1_u10_u0_n104 ) , .A( u1_u10_u0_n105 ) , .ZN( u1_u10_u0_n106 ) , .C2( u1_u10_u0_n113 ) , .C1( u1_u10_u0_n160 ) );
  OR4_X1 u1_u10_u0_U76 (.ZN( u1_out10_17 ) , .A4( u1_u10_u0_n122 ) , .A2( u1_u10_u0_n123 ) , .A1( u1_u10_u0_n124 ) , .A3( u1_u10_u0_n170 ) );
  AOI21_X1 u1_u10_u0_U77 (.B2( u1_u10_u0_n107 ) , .ZN( u1_u10_u0_n124 ) , .B1( u1_u10_u0_n128 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U78 (.A( u1_u10_u0_n111 ) , .ZN( u1_u10_u0_n170 ) );
  OR4_X1 u1_u10_u0_U79 (.ZN( u1_out10_31 ) , .A4( u1_u10_u0_n155 ) , .A2( u1_u10_u0_n156 ) , .A1( u1_u10_u0_n157 ) , .A3( u1_u10_u0_n173 ) );
  AND2_X1 u1_u10_u0_U8 (.A1( u1_u10_u0_n114 ) , .A2( u1_u10_u0_n121 ) , .ZN( u1_u10_u0_n146 ) );
  AOI21_X1 u1_u10_u0_U80 (.A( u1_u10_u0_n138 ) , .B2( u1_u10_u0_n139 ) , .B1( u1_u10_u0_n140 ) , .ZN( u1_u10_u0_n157 ) );
  AOI21_X1 u1_u10_u0_U81 (.B2( u1_u10_u0_n141 ) , .B1( u1_u10_u0_n142 ) , .ZN( u1_u10_u0_n156 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U82 (.A( u1_u10_u0_n126 ) , .ZN( u1_u10_u0_n168 ) );
  AOI211_X1 u1_u10_u0_U83 (.B( u1_u10_u0_n133 ) , .A( u1_u10_u0_n134 ) , .C2( u1_u10_u0_n135 ) , .C1( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n137 ) );
  AOI211_X1 u1_u10_u0_U84 (.B( u1_u10_u0_n115 ) , .A( u1_u10_u0_n116 ) , .C2( u1_u10_u0_n117 ) , .C1( u1_u10_u0_n118 ) , .ZN( u1_u10_u0_n119 ) );
  INV_X1 u1_u10_u0_U85 (.A( u1_u10_u0_n119 ) , .ZN( u1_u10_u0_n167 ) );
  NAND2_X1 u1_u10_u0_U86 (.ZN( u1_u10_u0_n110 ) , .A2( u1_u10_u0_n132 ) , .A1( u1_u10_u0_n145 ) );
  OAI22_X1 u1_u10_u0_U87 (.ZN( u1_u10_u0_n105 ) , .A2( u1_u10_u0_n132 ) , .B1( u1_u10_u0_n146 ) , .A1( u1_u10_u0_n147 ) , .B2( u1_u10_u0_n161 ) );
  NAND3_X1 u1_u10_u0_U88 (.ZN( u1_out10_23 ) , .A3( u1_u10_u0_n137 ) , .A1( u1_u10_u0_n168 ) , .A2( u1_u10_u0_n171 ) );
  NAND3_X1 u1_u10_u0_U89 (.A3( u1_u10_u0_n127 ) , .A2( u1_u10_u0_n128 ) , .ZN( u1_u10_u0_n135 ) , .A1( u1_u10_u0_n150 ) );
  AND2_X1 u1_u10_u0_U9 (.A1( u1_u10_u0_n131 ) , .ZN( u1_u10_u0_n141 ) , .A2( u1_u10_u0_n150 ) );
  NAND3_X1 u1_u10_u0_U90 (.ZN( u1_u10_u0_n117 ) , .A3( u1_u10_u0_n132 ) , .A2( u1_u10_u0_n139 ) , .A1( u1_u10_u0_n148 ) );
  NAND3_X1 u1_u10_u0_U91 (.ZN( u1_u10_u0_n109 ) , .A2( u1_u10_u0_n114 ) , .A3( u1_u10_u0_n140 ) , .A1( u1_u10_u0_n149 ) );
  NAND3_X1 u1_u10_u0_U92 (.ZN( u1_out10_9 ) , .A3( u1_u10_u0_n106 ) , .A2( u1_u10_u0_n171 ) , .A1( u1_u10_u0_n174 ) );
  NAND3_X1 u1_u10_u0_U93 (.A2( u1_u10_u0_n128 ) , .A1( u1_u10_u0_n132 ) , .A3( u1_u10_u0_n146 ) , .ZN( u1_u10_u0_n97 ) );
  AOI21_X1 u1_u10_u1_U10 (.B2( u1_u10_u1_n155 ) , .B1( u1_u10_u1_n156 ) , .ZN( u1_u10_u1_n157 ) , .A( u1_u10_u1_n174 ) );
  NAND3_X1 u1_u10_u1_U100 (.ZN( u1_u10_u1_n113 ) , .A1( u1_u10_u1_n120 ) , .A3( u1_u10_u1_n133 ) , .A2( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U11 (.ZN( u1_u10_u1_n140 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U12 (.A1( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n153 ) );
  AOI22_X1 u1_u10_u1_U13 (.B2( u1_u10_u1_n136 ) , .A2( u1_u10_u1_n137 ) , .ZN( u1_u10_u1_n143 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U14 (.A( u1_u10_u1_n147 ) , .ZN( u1_u10_u1_n181 ) );
  INV_X1 u1_u10_u1_U15 (.A( u1_u10_u1_n139 ) , .ZN( u1_u10_u1_n174 ) );
  OR4_X1 u1_u10_u1_U16 (.A4( u1_u10_u1_n106 ) , .A3( u1_u10_u1_n107 ) , .ZN( u1_u10_u1_n108 ) , .A1( u1_u10_u1_n117 ) , .A2( u1_u10_u1_n184 ) );
  AOI21_X1 u1_u10_u1_U17 (.ZN( u1_u10_u1_n106 ) , .A( u1_u10_u1_n112 ) , .B1( u1_u10_u1_n154 ) , .B2( u1_u10_u1_n156 ) );
  AOI21_X1 u1_u10_u1_U18 (.ZN( u1_u10_u1_n107 ) , .B1( u1_u10_u1_n134 ) , .B2( u1_u10_u1_n149 ) , .A( u1_u10_u1_n174 ) );
  INV_X1 u1_u10_u1_U19 (.A( u1_u10_u1_n101 ) , .ZN( u1_u10_u1_n184 ) );
  INV_X1 u1_u10_u1_U20 (.A( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n171 ) );
  NAND2_X1 u1_u10_u1_U21 (.ZN( u1_u10_u1_n141 ) , .A1( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n156 ) );
  AND2_X1 u1_u10_u1_U22 (.A1( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n161 ) );
  NAND2_X1 u1_u10_u1_U23 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n148 ) );
  NAND2_X1 u1_u10_u1_U24 (.A2( u1_u10_u1_n133 ) , .A1( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n159 ) );
  NAND2_X1 u1_u10_u1_U25 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n120 ) , .ZN( u1_u10_u1_n132 ) );
  INV_X1 u1_u10_u1_U26 (.A( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n178 ) );
  INV_X1 u1_u10_u1_U27 (.A( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n183 ) );
  AND2_X1 u1_u10_u1_U28 (.A1( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n149 ) );
  INV_X1 u1_u10_u1_U29 (.A( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n180 ) );
  INV_X1 u1_u10_u1_U3 (.A( u1_u10_u1_n159 ) , .ZN( u1_u10_u1_n182 ) );
  OAI221_X1 u1_u10_u1_U30 (.A( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n138 ) , .B2( u1_u10_u1_n152 ) , .C1( u1_u10_u1_n174 ) , .B1( u1_u10_u1_n187 ) );
  INV_X1 u1_u10_u1_U31 (.A( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n187 ) );
  AOI211_X1 u1_u10_u1_U32 (.B( u1_u10_u1_n117 ) , .A( u1_u10_u1_n118 ) , .ZN( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n146 ) , .C1( u1_u10_u1_n159 ) );
  NOR2_X1 u1_u10_u1_U33 (.A1( u1_u10_u1_n168 ) , .A2( u1_u10_u1_n176 ) , .ZN( u1_u10_u1_n98 ) );
  AOI211_X1 u1_u10_u1_U34 (.B( u1_u10_u1_n162 ) , .A( u1_u10_u1_n163 ) , .C2( u1_u10_u1_n164 ) , .ZN( u1_u10_u1_n165 ) , .C1( u1_u10_u1_n171 ) );
  AOI21_X1 u1_u10_u1_U35 (.A( u1_u10_u1_n160 ) , .B2( u1_u10_u1_n161 ) , .ZN( u1_u10_u1_n162 ) , .B1( u1_u10_u1_n182 ) );
  OR2_X1 u1_u10_u1_U36 (.A2( u1_u10_u1_n157 ) , .A1( u1_u10_u1_n158 ) , .ZN( u1_u10_u1_n163 ) );
  OAI21_X1 u1_u10_u1_U37 (.B2( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n145 ) , .B1( u1_u10_u1_n160 ) , .A( u1_u10_u1_n185 ) );
  INV_X1 u1_u10_u1_U38 (.A( u1_u10_u1_n122 ) , .ZN( u1_u10_u1_n185 ) );
  AOI21_X1 u1_u10_u1_U39 (.B2( u1_u10_u1_n120 ) , .B1( u1_u10_u1_n121 ) , .ZN( u1_u10_u1_n122 ) , .A( u1_u10_u1_n128 ) );
  AOI221_X1 u1_u10_u1_U4 (.A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .C1( u1_u10_u1_n140 ) , .B2( u1_u10_u1_n141 ) , .ZN( u1_u10_u1_n142 ) , .B1( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U40 (.A1( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n146 ) , .A2( u1_u10_u1_n160 ) );
  NAND2_X1 u1_u10_u1_U41 (.A2( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n139 ) , .A1( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U42 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n156 ) , .A2( u1_u10_u1_n99 ) );
  AOI221_X1 u1_u10_u1_U43 (.B1( u1_u10_u1_n140 ) , .ZN( u1_u10_u1_n167 ) , .B2( u1_u10_u1_n172 ) , .C2( u1_u10_u1_n175 ) , .C1( u1_u10_u1_n178 ) , .A( u1_u10_u1_n188 ) );
  INV_X1 u1_u10_u1_U44 (.ZN( u1_u10_u1_n188 ) , .A( u1_u10_u1_n97 ) );
  AOI211_X1 u1_u10_u1_U45 (.A( u1_u10_u1_n118 ) , .C1( u1_u10_u1_n132 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n96 ) , .ZN( u1_u10_u1_n97 ) );
  AOI21_X1 u1_u10_u1_U46 (.B2( u1_u10_u1_n121 ) , .B1( u1_u10_u1_n135 ) , .A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n96 ) );
  NOR2_X1 u1_u10_u1_U47 (.ZN( u1_u10_u1_n117 ) , .A1( u1_u10_u1_n121 ) , .A2( u1_u10_u1_n160 ) );
  AOI21_X1 u1_u10_u1_U48 (.A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n130 ) , .B1( u1_u10_u1_n150 ) );
  NAND2_X1 u1_u10_u1_U49 (.ZN( u1_u10_u1_n112 ) , .A1( u1_u10_u1_n169 ) , .A2( u1_u10_u1_n170 ) );
  AOI211_X1 u1_u10_u1_U5 (.ZN( u1_u10_u1_n124 ) , .A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n145 ) , .C1( u1_u10_u1_n147 ) );
  NAND2_X1 u1_u10_u1_U50 (.ZN( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n95 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U51 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n154 ) , .A2( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U52 (.A2( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n135 ) , .A1( u1_u10_u1_n99 ) );
  AOI21_X1 u1_u10_u1_U53 (.A( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n153 ) , .B1( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n158 ) );
  INV_X1 u1_u10_u1_U54 (.A( u1_u10_u1_n160 ) , .ZN( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U55 (.A1( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n116 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U56 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n131 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U57 (.A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n121 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U58 (.A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U59 (.A2( u1_u10_u1_n104 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n133 ) );
  AOI22_X1 u1_u10_u1_U6 (.B2( u1_u10_u1_n113 ) , .A2( u1_u10_u1_n114 ) , .ZN( u1_u10_u1_n125 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  NAND2_X1 u1_u10_u1_U60 (.ZN( u1_u10_u1_n150 ) , .A2( u1_u10_u1_n98 ) , .A1( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U61 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n155 ) , .A2( u1_u10_u1_n95 ) );
  OAI21_X1 u1_u10_u1_U62 (.ZN( u1_u10_u1_n109 ) , .B1( u1_u10_u1_n129 ) , .B2( u1_u10_u1_n160 ) , .A( u1_u10_u1_n167 ) );
  NAND2_X1 u1_u10_u1_U63 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n120 ) );
  NAND2_X1 u1_u10_u1_U64 (.A1( u1_u10_u1_n102 ) , .A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n115 ) );
  NAND2_X1 u1_u10_u1_U65 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n151 ) );
  NAND2_X1 u1_u10_u1_U66 (.A2( u1_u10_u1_n103 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n161 ) );
  INV_X1 u1_u10_u1_U67 (.A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U68 (.A( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n172 ) );
  NAND2_X1 u1_u10_u1_U69 (.A2( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n123 ) );
  NAND2_X1 u1_u10_u1_U7 (.ZN( u1_u10_u1_n114 ) , .A1( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n156 ) );
  NOR2_X1 u1_u10_u1_U70 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n95 ) );
  NOR2_X1 u1_u10_u1_U71 (.A1( u1_u10_X_12 ) , .A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n100 ) );
  NOR2_X1 u1_u10_u1_U72 (.A2( u1_u10_X_8 ) , .A1( u1_u10_u1_n177 ) , .ZN( u1_u10_u1_n99 ) );
  NOR2_X1 u1_u10_u1_U73 (.A2( u1_u10_X_12 ) , .ZN( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n176 ) );
  NOR2_X1 u1_u10_u1_U74 (.A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n105 ) , .A1( u1_u10_u1_n168 ) );
  NAND2_X1 u1_u10_u1_U75 (.A1( u1_u10_X_10 ) , .ZN( u1_u10_u1_n160 ) , .A2( u1_u10_u1_n169 ) );
  NAND2_X1 u1_u10_u1_U76 (.A2( u1_u10_X_10 ) , .A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U77 (.A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n128 ) , .A2( u1_u10_u1_n170 ) );
  AND2_X1 u1_u10_u1_U78 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n104 ) );
  AND2_X1 u1_u10_u1_U79 (.A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n103 ) , .A2( u1_u10_u1_n177 ) );
  NOR2_X1 u1_u10_u1_U8 (.A1( u1_u10_u1_n112 ) , .A2( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n118 ) );
  INV_X1 u1_u10_u1_U80 (.A( u1_u10_X_10 ) , .ZN( u1_u10_u1_n170 ) );
  INV_X1 u1_u10_u1_U81 (.A( u1_u10_X_9 ) , .ZN( u1_u10_u1_n176 ) );
  INV_X1 u1_u10_u1_U82 (.A( u1_u10_X_11 ) , .ZN( u1_u10_u1_n169 ) );
  INV_X1 u1_u10_u1_U83 (.A( u1_u10_X_12 ) , .ZN( u1_u10_u1_n168 ) );
  INV_X1 u1_u10_u1_U84 (.A( u1_u10_X_7 ) , .ZN( u1_u10_u1_n177 ) );
  NAND4_X1 u1_u10_u1_U85 (.ZN( u1_out10_18 ) , .A4( u1_u10_u1_n165 ) , .A3( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n167 ) , .A2( u1_u10_u1_n186 ) );
  AOI22_X1 u1_u10_u1_U86 (.B2( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n172 ) );
  INV_X1 u1_u10_u1_U87 (.A( u1_u10_u1_n145 ) , .ZN( u1_u10_u1_n186 ) );
  NAND4_X1 u1_u10_u1_U88 (.ZN( u1_out10_2 ) , .A4( u1_u10_u1_n142 ) , .A3( u1_u10_u1_n143 ) , .A2( u1_u10_u1_n144 ) , .A1( u1_u10_u1_n179 ) );
  OAI21_X1 u1_u10_u1_U89 (.B2( u1_u10_u1_n132 ) , .ZN( u1_u10_u1_n144 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n180 ) );
  OAI21_X1 u1_u10_u1_U9 (.ZN( u1_u10_u1_n101 ) , .B1( u1_u10_u1_n141 ) , .A( u1_u10_u1_n146 ) , .B2( u1_u10_u1_n183 ) );
  INV_X1 u1_u10_u1_U90 (.A( u1_u10_u1_n130 ) , .ZN( u1_u10_u1_n179 ) );
  OR4_X1 u1_u10_u1_U91 (.ZN( u1_out10_13 ) , .A4( u1_u10_u1_n108 ) , .A3( u1_u10_u1_n109 ) , .A2( u1_u10_u1_n110 ) , .A1( u1_u10_u1_n111 ) );
  AOI21_X1 u1_u10_u1_U92 (.ZN( u1_u10_u1_n111 ) , .A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n131 ) , .B1( u1_u10_u1_n135 ) );
  AOI21_X1 u1_u10_u1_U93 (.ZN( u1_u10_u1_n110 ) , .A( u1_u10_u1_n116 ) , .B1( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n160 ) );
  NAND4_X1 u1_u10_u1_U94 (.ZN( u1_out10_28 ) , .A4( u1_u10_u1_n124 ) , .A3( u1_u10_u1_n125 ) , .A2( u1_u10_u1_n126 ) , .A1( u1_u10_u1_n127 ) );
  OAI21_X1 u1_u10_u1_U95 (.ZN( u1_u10_u1_n127 ) , .B2( u1_u10_u1_n139 ) , .B1( u1_u10_u1_n175 ) , .A( u1_u10_u1_n183 ) );
  OAI21_X1 u1_u10_u1_U96 (.ZN( u1_u10_u1_n126 ) , .B2( u1_u10_u1_n140 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n178 ) );
  NAND3_X1 u1_u10_u1_U97 (.A3( u1_u10_u1_n149 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n164 ) );
  NAND3_X1 u1_u10_u1_U98 (.A3( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n136 ) , .A1( u1_u10_u1_n151 ) );
  NAND3_X1 u1_u10_u1_U99 (.A1( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n137 ) , .A2( u1_u10_u1_n154 ) , .A3( u1_u10_u1_n181 ) );
  OAI22_X1 u1_u10_u2_U10 (.ZN( u1_u10_u2_n109 ) , .A2( u1_u10_u2_n113 ) , .B2( u1_u10_u2_n133 ) , .B1( u1_u10_u2_n167 ) , .A1( u1_u10_u2_n168 ) );
  NAND3_X1 u1_u10_u2_U100 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n98 ) );
  OAI22_X1 u1_u10_u2_U11 (.B1( u1_u10_u2_n151 ) , .A2( u1_u10_u2_n152 ) , .A1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n160 ) , .B2( u1_u10_u2_n168 ) );
  NOR3_X1 u1_u10_u2_U12 (.A1( u1_u10_u2_n150 ) , .ZN( u1_u10_u2_n151 ) , .A3( u1_u10_u2_n175 ) , .A2( u1_u10_u2_n188 ) );
  AOI21_X1 u1_u10_u2_U13 (.ZN( u1_u10_u2_n144 ) , .B2( u1_u10_u2_n155 ) , .A( u1_u10_u2_n172 ) , .B1( u1_u10_u2_n185 ) );
  AOI21_X1 u1_u10_u2_U14 (.B2( u1_u10_u2_n143 ) , .ZN( u1_u10_u2_n145 ) , .B1( u1_u10_u2_n152 ) , .A( u1_u10_u2_n171 ) );
  AOI21_X1 u1_u10_u2_U15 (.B2( u1_u10_u2_n120 ) , .B1( u1_u10_u2_n121 ) , .ZN( u1_u10_u2_n126 ) , .A( u1_u10_u2_n167 ) );
  INV_X1 u1_u10_u2_U16 (.A( u1_u10_u2_n156 ) , .ZN( u1_u10_u2_n171 ) );
  INV_X1 u1_u10_u2_U17 (.A( u1_u10_u2_n120 ) , .ZN( u1_u10_u2_n188 ) );
  NAND2_X1 u1_u10_u2_U18 (.A2( u1_u10_u2_n122 ) , .ZN( u1_u10_u2_n150 ) , .A1( u1_u10_u2_n152 ) );
  INV_X1 u1_u10_u2_U19 (.A( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n170 ) );
  INV_X1 u1_u10_u2_U20 (.A( u1_u10_u2_n137 ) , .ZN( u1_u10_u2_n173 ) );
  NAND2_X1 u1_u10_u2_U21 (.A1( u1_u10_u2_n132 ) , .A2( u1_u10_u2_n139 ) , .ZN( u1_u10_u2_n157 ) );
  INV_X1 u1_u10_u2_U22 (.A( u1_u10_u2_n113 ) , .ZN( u1_u10_u2_n178 ) );
  INV_X1 u1_u10_u2_U23 (.A( u1_u10_u2_n139 ) , .ZN( u1_u10_u2_n175 ) );
  INV_X1 u1_u10_u2_U24 (.A( u1_u10_u2_n155 ) , .ZN( u1_u10_u2_n181 ) );
  INV_X1 u1_u10_u2_U25 (.A( u1_u10_u2_n119 ) , .ZN( u1_u10_u2_n177 ) );
  INV_X1 u1_u10_u2_U26 (.A( u1_u10_u2_n116 ) , .ZN( u1_u10_u2_n180 ) );
  INV_X1 u1_u10_u2_U27 (.A( u1_u10_u2_n131 ) , .ZN( u1_u10_u2_n179 ) );
  INV_X1 u1_u10_u2_U28 (.A( u1_u10_u2_n154 ) , .ZN( u1_u10_u2_n176 ) );
  NAND2_X1 u1_u10_u2_U29 (.A2( u1_u10_u2_n116 ) , .A1( u1_u10_u2_n117 ) , .ZN( u1_u10_u2_n118 ) );
  NOR2_X1 u1_u10_u2_U3 (.ZN( u1_u10_u2_n121 ) , .A2( u1_u10_u2_n177 ) , .A1( u1_u10_u2_n180 ) );
  INV_X1 u1_u10_u2_U30 (.A( u1_u10_u2_n132 ) , .ZN( u1_u10_u2_n182 ) );
  INV_X1 u1_u10_u2_U31 (.A( u1_u10_u2_n158 ) , .ZN( u1_u10_u2_n183 ) );
  OAI21_X1 u1_u10_u2_U32 (.A( u1_u10_u2_n156 ) , .B1( u1_u10_u2_n157 ) , .ZN( u1_u10_u2_n158 ) , .B2( u1_u10_u2_n179 ) );
  NOR2_X1 u1_u10_u2_U33 (.ZN( u1_u10_u2_n156 ) , .A1( u1_u10_u2_n166 ) , .A2( u1_u10_u2_n169 ) );
  NOR2_X1 u1_u10_u2_U34 (.A2( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n137 ) , .A1( u1_u10_u2_n140 ) );
  NOR2_X1 u1_u10_u2_U35 (.A2( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n153 ) , .A1( u1_u10_u2_n156 ) );
  AOI211_X1 u1_u10_u2_U36 (.ZN( u1_u10_u2_n130 ) , .C1( u1_u10_u2_n138 ) , .C2( u1_u10_u2_n179 ) , .B( u1_u10_u2_n96 ) , .A( u1_u10_u2_n97 ) );
  OAI22_X1 u1_u10_u2_U37 (.B1( u1_u10_u2_n133 ) , .A2( u1_u10_u2_n137 ) , .A1( u1_u10_u2_n152 ) , .B2( u1_u10_u2_n168 ) , .ZN( u1_u10_u2_n97 ) );
  OAI221_X1 u1_u10_u2_U38 (.B1( u1_u10_u2_n113 ) , .C1( u1_u10_u2_n132 ) , .A( u1_u10_u2_n149 ) , .B2( u1_u10_u2_n171 ) , .C2( u1_u10_u2_n172 ) , .ZN( u1_u10_u2_n96 ) );
  OAI221_X1 u1_u10_u2_U39 (.A( u1_u10_u2_n115 ) , .C2( u1_u10_u2_n123 ) , .B2( u1_u10_u2_n143 ) , .B1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n163 ) , .C1( u1_u10_u2_n168 ) );
  INV_X1 u1_u10_u2_U4 (.A( u1_u10_u2_n134 ) , .ZN( u1_u10_u2_n185 ) );
  OAI21_X1 u1_u10_u2_U40 (.A( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n115 ) , .B1( u1_u10_u2_n176 ) , .B2( u1_u10_u2_n178 ) );
  OAI221_X1 u1_u10_u2_U41 (.A( u1_u10_u2_n135 ) , .B2( u1_u10_u2_n136 ) , .B1( u1_u10_u2_n137 ) , .ZN( u1_u10_u2_n162 ) , .C2( u1_u10_u2_n167 ) , .C1( u1_u10_u2_n185 ) );
  AND3_X1 u1_u10_u2_U42 (.A3( u1_u10_u2_n131 ) , .A2( u1_u10_u2_n132 ) , .A1( u1_u10_u2_n133 ) , .ZN( u1_u10_u2_n136 ) );
  AOI22_X1 u1_u10_u2_U43 (.ZN( u1_u10_u2_n135 ) , .B1( u1_u10_u2_n140 ) , .A1( u1_u10_u2_n156 ) , .B2( u1_u10_u2_n180 ) , .A2( u1_u10_u2_n188 ) );
  AOI21_X1 u1_u10_u2_U44 (.ZN( u1_u10_u2_n149 ) , .B1( u1_u10_u2_n173 ) , .B2( u1_u10_u2_n188 ) , .A( u1_u10_u2_n95 ) );
  AND3_X1 u1_u10_u2_U45 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n156 ) , .ZN( u1_u10_u2_n95 ) );
  OAI21_X1 u1_u10_u2_U46 (.A( u1_u10_u2_n101 ) , .B2( u1_u10_u2_n121 ) , .B1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n164 ) );
  NAND2_X1 u1_u10_u2_U47 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n155 ) );
  NAND2_X1 u1_u10_u2_U48 (.A2( u1_u10_u2_n105 ) , .A1( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n143 ) );
  NAND2_X1 u1_u10_u2_U49 (.A1( u1_u10_u2_n104 ) , .A2( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n152 ) );
  INV_X1 u1_u10_u2_U5 (.A( u1_u10_u2_n150 ) , .ZN( u1_u10_u2_n184 ) );
  NAND2_X1 u1_u10_u2_U50 (.A1( u1_u10_u2_n100 ) , .A2( u1_u10_u2_n105 ) , .ZN( u1_u10_u2_n132 ) );
  INV_X1 u1_u10_u2_U51 (.A( u1_u10_u2_n140 ) , .ZN( u1_u10_u2_n168 ) );
  INV_X1 u1_u10_u2_U52 (.A( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n167 ) );
  OAI21_X1 u1_u10_u2_U53 (.A( u1_u10_u2_n141 ) , .B2( u1_u10_u2_n142 ) , .ZN( u1_u10_u2_n146 ) , .B1( u1_u10_u2_n153 ) );
  OAI21_X1 u1_u10_u2_U54 (.A( u1_u10_u2_n140 ) , .ZN( u1_u10_u2_n141 ) , .B1( u1_u10_u2_n176 ) , .B2( u1_u10_u2_n177 ) );
  NOR3_X1 u1_u10_u2_U55 (.ZN( u1_u10_u2_n142 ) , .A3( u1_u10_u2_n175 ) , .A2( u1_u10_u2_n178 ) , .A1( u1_u10_u2_n181 ) );
  NAND2_X1 u1_u10_u2_U56 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n113 ) );
  NAND2_X1 u1_u10_u2_U57 (.A1( u1_u10_u2_n106 ) , .A2( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n131 ) );
  NAND2_X1 u1_u10_u2_U58 (.A1( u1_u10_u2_n103 ) , .A2( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n139 ) );
  NAND2_X1 u1_u10_u2_U59 (.A1( u1_u10_u2_n103 ) , .A2( u1_u10_u2_n105 ) , .ZN( u1_u10_u2_n133 ) );
  NOR4_X1 u1_u10_u2_U6 (.A4( u1_u10_u2_n124 ) , .A3( u1_u10_u2_n125 ) , .A2( u1_u10_u2_n126 ) , .A1( u1_u10_u2_n127 ) , .ZN( u1_u10_u2_n128 ) );
  NAND2_X1 u1_u10_u2_U60 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n103 ) , .ZN( u1_u10_u2_n154 ) );
  NAND2_X1 u1_u10_u2_U61 (.A2( u1_u10_u2_n103 ) , .A1( u1_u10_u2_n104 ) , .ZN( u1_u10_u2_n119 ) );
  NAND2_X1 u1_u10_u2_U62 (.A2( u1_u10_u2_n107 ) , .A1( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n123 ) );
  NAND2_X1 u1_u10_u2_U63 (.A1( u1_u10_u2_n104 ) , .A2( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n122 ) );
  INV_X1 u1_u10_u2_U64 (.A( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n172 ) );
  NAND2_X1 u1_u10_u2_U65 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n102 ) , .ZN( u1_u10_u2_n116 ) );
  NAND2_X1 u1_u10_u2_U66 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n120 ) );
  NAND2_X1 u1_u10_u2_U67 (.A2( u1_u10_u2_n105 ) , .A1( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n117 ) );
  INV_X1 u1_u10_u2_U68 (.ZN( u1_u10_u2_n187 ) , .A( u1_u10_u2_n99 ) );
  OAI21_X1 u1_u10_u2_U69 (.B1( u1_u10_u2_n137 ) , .B2( u1_u10_u2_n143 ) , .A( u1_u10_u2_n98 ) , .ZN( u1_u10_u2_n99 ) );
  AOI21_X1 u1_u10_u2_U7 (.ZN( u1_u10_u2_n124 ) , .B1( u1_u10_u2_n131 ) , .B2( u1_u10_u2_n143 ) , .A( u1_u10_u2_n172 ) );
  NOR2_X1 u1_u10_u2_U70 (.A2( u1_u10_X_16 ) , .ZN( u1_u10_u2_n140 ) , .A1( u1_u10_u2_n166 ) );
  NOR2_X1 u1_u10_u2_U71 (.A2( u1_u10_X_13 ) , .A1( u1_u10_X_14 ) , .ZN( u1_u10_u2_n100 ) );
  NOR2_X1 u1_u10_u2_U72 (.A2( u1_u10_X_16 ) , .A1( u1_u10_X_17 ) , .ZN( u1_u10_u2_n138 ) );
  NOR2_X1 u1_u10_u2_U73 (.A2( u1_u10_X_15 ) , .A1( u1_u10_X_18 ) , .ZN( u1_u10_u2_n104 ) );
  NOR2_X1 u1_u10_u2_U74 (.A2( u1_u10_X_14 ) , .ZN( u1_u10_u2_n103 ) , .A1( u1_u10_u2_n174 ) );
  NOR2_X1 u1_u10_u2_U75 (.A2( u1_u10_X_15 ) , .ZN( u1_u10_u2_n102 ) , .A1( u1_u10_u2_n165 ) );
  NOR2_X1 u1_u10_u2_U76 (.A2( u1_u10_X_17 ) , .ZN( u1_u10_u2_n114 ) , .A1( u1_u10_u2_n169 ) );
  AND2_X1 u1_u10_u2_U77 (.A1( u1_u10_X_15 ) , .ZN( u1_u10_u2_n105 ) , .A2( u1_u10_u2_n165 ) );
  AND2_X1 u1_u10_u2_U78 (.A2( u1_u10_X_15 ) , .A1( u1_u10_X_18 ) , .ZN( u1_u10_u2_n107 ) );
  AND2_X1 u1_u10_u2_U79 (.A1( u1_u10_X_14 ) , .ZN( u1_u10_u2_n106 ) , .A2( u1_u10_u2_n174 ) );
  AOI21_X1 u1_u10_u2_U8 (.B2( u1_u10_u2_n119 ) , .ZN( u1_u10_u2_n127 ) , .A( u1_u10_u2_n137 ) , .B1( u1_u10_u2_n155 ) );
  AND2_X1 u1_u10_u2_U80 (.A1( u1_u10_X_13 ) , .A2( u1_u10_X_14 ) , .ZN( u1_u10_u2_n108 ) );
  INV_X1 u1_u10_u2_U81 (.A( u1_u10_X_16 ) , .ZN( u1_u10_u2_n169 ) );
  INV_X1 u1_u10_u2_U82 (.A( u1_u10_X_17 ) , .ZN( u1_u10_u2_n166 ) );
  INV_X1 u1_u10_u2_U83 (.A( u1_u10_X_13 ) , .ZN( u1_u10_u2_n174 ) );
  INV_X1 u1_u10_u2_U84 (.A( u1_u10_X_18 ) , .ZN( u1_u10_u2_n165 ) );
  NAND4_X1 u1_u10_u2_U85 (.ZN( u1_out10_30 ) , .A4( u1_u10_u2_n147 ) , .A3( u1_u10_u2_n148 ) , .A2( u1_u10_u2_n149 ) , .A1( u1_u10_u2_n187 ) );
  NOR3_X1 u1_u10_u2_U86 (.A3( u1_u10_u2_n144 ) , .A2( u1_u10_u2_n145 ) , .A1( u1_u10_u2_n146 ) , .ZN( u1_u10_u2_n147 ) );
  AOI21_X1 u1_u10_u2_U87 (.B2( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n148 ) , .A( u1_u10_u2_n162 ) , .B1( u1_u10_u2_n182 ) );
  NAND4_X1 u1_u10_u2_U88 (.ZN( u1_out10_24 ) , .A4( u1_u10_u2_n111 ) , .A3( u1_u10_u2_n112 ) , .A1( u1_u10_u2_n130 ) , .A2( u1_u10_u2_n187 ) );
  AOI221_X1 u1_u10_u2_U89 (.A( u1_u10_u2_n109 ) , .B1( u1_u10_u2_n110 ) , .ZN( u1_u10_u2_n111 ) , .C1( u1_u10_u2_n134 ) , .C2( u1_u10_u2_n170 ) , .B2( u1_u10_u2_n173 ) );
  AOI21_X1 u1_u10_u2_U9 (.B2( u1_u10_u2_n123 ) , .ZN( u1_u10_u2_n125 ) , .A( u1_u10_u2_n171 ) , .B1( u1_u10_u2_n184 ) );
  AOI21_X1 u1_u10_u2_U90 (.ZN( u1_u10_u2_n112 ) , .B2( u1_u10_u2_n156 ) , .A( u1_u10_u2_n164 ) , .B1( u1_u10_u2_n181 ) );
  NAND4_X1 u1_u10_u2_U91 (.ZN( u1_out10_16 ) , .A4( u1_u10_u2_n128 ) , .A3( u1_u10_u2_n129 ) , .A1( u1_u10_u2_n130 ) , .A2( u1_u10_u2_n186 ) );
  AOI22_X1 u1_u10_u2_U92 (.A2( u1_u10_u2_n118 ) , .ZN( u1_u10_u2_n129 ) , .A1( u1_u10_u2_n140 ) , .B1( u1_u10_u2_n157 ) , .B2( u1_u10_u2_n170 ) );
  INV_X1 u1_u10_u2_U93 (.A( u1_u10_u2_n163 ) , .ZN( u1_u10_u2_n186 ) );
  OR4_X1 u1_u10_u2_U94 (.ZN( u1_out10_6 ) , .A4( u1_u10_u2_n161 ) , .A3( u1_u10_u2_n162 ) , .A2( u1_u10_u2_n163 ) , .A1( u1_u10_u2_n164 ) );
  OR3_X1 u1_u10_u2_U95 (.A2( u1_u10_u2_n159 ) , .A1( u1_u10_u2_n160 ) , .ZN( u1_u10_u2_n161 ) , .A3( u1_u10_u2_n183 ) );
  AOI21_X1 u1_u10_u2_U96 (.B2( u1_u10_u2_n154 ) , .B1( u1_u10_u2_n155 ) , .ZN( u1_u10_u2_n159 ) , .A( u1_u10_u2_n167 ) );
  NAND3_X1 u1_u10_u2_U97 (.A2( u1_u10_u2_n117 ) , .A1( u1_u10_u2_n122 ) , .A3( u1_u10_u2_n123 ) , .ZN( u1_u10_u2_n134 ) );
  NAND3_X1 u1_u10_u2_U98 (.ZN( u1_u10_u2_n110 ) , .A2( u1_u10_u2_n131 ) , .A3( u1_u10_u2_n139 ) , .A1( u1_u10_u2_n154 ) );
  NAND3_X1 u1_u10_u2_U99 (.A2( u1_u10_u2_n100 ) , .ZN( u1_u10_u2_n101 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n114 ) );
  INV_X1 u1_u10_u5_U10 (.A( u1_u10_u5_n121 ) , .ZN( u1_u10_u5_n177 ) );
  NOR3_X1 u1_u10_u5_U100 (.A3( u1_u10_u5_n141 ) , .A1( u1_u10_u5_n142 ) , .ZN( u1_u10_u5_n143 ) , .A2( u1_u10_u5_n191 ) );
  NAND4_X1 u1_u10_u5_U101 (.ZN( u1_out10_4 ) , .A4( u1_u10_u5_n112 ) , .A2( u1_u10_u5_n113 ) , .A1( u1_u10_u5_n114 ) , .A3( u1_u10_u5_n195 ) );
  AOI211_X1 u1_u10_u5_U102 (.A( u1_u10_u5_n110 ) , .C1( u1_u10_u5_n111 ) , .ZN( u1_u10_u5_n112 ) , .B( u1_u10_u5_n118 ) , .C2( u1_u10_u5_n177 ) );
  AOI222_X1 u1_u10_u5_U103 (.ZN( u1_u10_u5_n113 ) , .A1( u1_u10_u5_n131 ) , .C1( u1_u10_u5_n148 ) , .B2( u1_u10_u5_n174 ) , .C2( u1_u10_u5_n178 ) , .A2( u1_u10_u5_n179 ) , .B1( u1_u10_u5_n99 ) );
  NAND3_X1 u1_u10_u5_U104 (.A2( u1_u10_u5_n154 ) , .A3( u1_u10_u5_n158 ) , .A1( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n99 ) );
  NOR2_X1 u1_u10_u5_U11 (.ZN( u1_u10_u5_n160 ) , .A2( u1_u10_u5_n173 ) , .A1( u1_u10_u5_n177 ) );
  INV_X1 u1_u10_u5_U12 (.A( u1_u10_u5_n150 ) , .ZN( u1_u10_u5_n174 ) );
  AOI21_X1 u1_u10_u5_U13 (.A( u1_u10_u5_n160 ) , .B2( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n162 ) , .B1( u1_u10_u5_n192 ) );
  INV_X1 u1_u10_u5_U14 (.A( u1_u10_u5_n159 ) , .ZN( u1_u10_u5_n192 ) );
  AOI21_X1 u1_u10_u5_U15 (.A( u1_u10_u5_n156 ) , .B2( u1_u10_u5_n157 ) , .B1( u1_u10_u5_n158 ) , .ZN( u1_u10_u5_n163 ) );
  AOI21_X1 u1_u10_u5_U16 (.B2( u1_u10_u5_n139 ) , .B1( u1_u10_u5_n140 ) , .ZN( u1_u10_u5_n141 ) , .A( u1_u10_u5_n150 ) );
  OAI21_X1 u1_u10_u5_U17 (.A( u1_u10_u5_n133 ) , .B2( u1_u10_u5_n134 ) , .B1( u1_u10_u5_n135 ) , .ZN( u1_u10_u5_n142 ) );
  OAI21_X1 u1_u10_u5_U18 (.ZN( u1_u10_u5_n133 ) , .B2( u1_u10_u5_n147 ) , .A( u1_u10_u5_n173 ) , .B1( u1_u10_u5_n188 ) );
  NAND2_X1 u1_u10_u5_U19 (.A2( u1_u10_u5_n119 ) , .A1( u1_u10_u5_n123 ) , .ZN( u1_u10_u5_n137 ) );
  INV_X1 u1_u10_u5_U20 (.A( u1_u10_u5_n155 ) , .ZN( u1_u10_u5_n194 ) );
  NAND2_X1 u1_u10_u5_U21 (.A1( u1_u10_u5_n121 ) , .ZN( u1_u10_u5_n132 ) , .A2( u1_u10_u5_n172 ) );
  NAND2_X1 u1_u10_u5_U22 (.A2( u1_u10_u5_n122 ) , .ZN( u1_u10_u5_n136 ) , .A1( u1_u10_u5_n154 ) );
  NAND2_X1 u1_u10_u5_U23 (.A2( u1_u10_u5_n119 ) , .A1( u1_u10_u5_n120 ) , .ZN( u1_u10_u5_n159 ) );
  INV_X1 u1_u10_u5_U24 (.A( u1_u10_u5_n156 ) , .ZN( u1_u10_u5_n175 ) );
  INV_X1 u1_u10_u5_U25 (.A( u1_u10_u5_n158 ) , .ZN( u1_u10_u5_n188 ) );
  INV_X1 u1_u10_u5_U26 (.A( u1_u10_u5_n152 ) , .ZN( u1_u10_u5_n179 ) );
  INV_X1 u1_u10_u5_U27 (.A( u1_u10_u5_n140 ) , .ZN( u1_u10_u5_n182 ) );
  INV_X1 u1_u10_u5_U28 (.A( u1_u10_u5_n151 ) , .ZN( u1_u10_u5_n183 ) );
  INV_X1 u1_u10_u5_U29 (.A( u1_u10_u5_n123 ) , .ZN( u1_u10_u5_n185 ) );
  NOR2_X1 u1_u10_u5_U3 (.ZN( u1_u10_u5_n134 ) , .A1( u1_u10_u5_n183 ) , .A2( u1_u10_u5_n190 ) );
  INV_X1 u1_u10_u5_U30 (.A( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n184 ) );
  INV_X1 u1_u10_u5_U31 (.A( u1_u10_u5_n139 ) , .ZN( u1_u10_u5_n189 ) );
  INV_X1 u1_u10_u5_U32 (.A( u1_u10_u5_n157 ) , .ZN( u1_u10_u5_n190 ) );
  INV_X1 u1_u10_u5_U33 (.A( u1_u10_u5_n120 ) , .ZN( u1_u10_u5_n193 ) );
  NAND2_X1 u1_u10_u5_U34 (.ZN( u1_u10_u5_n111 ) , .A1( u1_u10_u5_n140 ) , .A2( u1_u10_u5_n155 ) );
  INV_X1 u1_u10_u5_U35 (.A( u1_u10_u5_n117 ) , .ZN( u1_u10_u5_n196 ) );
  OAI221_X1 u1_u10_u5_U36 (.A( u1_u10_u5_n116 ) , .ZN( u1_u10_u5_n117 ) , .B2( u1_u10_u5_n119 ) , .C1( u1_u10_u5_n153 ) , .C2( u1_u10_u5_n158 ) , .B1( u1_u10_u5_n172 ) );
  AOI222_X1 u1_u10_u5_U37 (.ZN( u1_u10_u5_n116 ) , .B2( u1_u10_u5_n145 ) , .C1( u1_u10_u5_n148 ) , .A2( u1_u10_u5_n174 ) , .C2( u1_u10_u5_n177 ) , .B1( u1_u10_u5_n187 ) , .A1( u1_u10_u5_n193 ) );
  INV_X1 u1_u10_u5_U38 (.A( u1_u10_u5_n115 ) , .ZN( u1_u10_u5_n187 ) );
  NOR2_X1 u1_u10_u5_U39 (.ZN( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n170 ) , .A2( u1_u10_u5_n180 ) );
  INV_X1 u1_u10_u5_U4 (.A( u1_u10_u5_n138 ) , .ZN( u1_u10_u5_n191 ) );
  AOI22_X1 u1_u10_u5_U40 (.B2( u1_u10_u5_n131 ) , .A2( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n169 ) , .B1( u1_u10_u5_n174 ) , .A1( u1_u10_u5_n185 ) );
  NOR2_X1 u1_u10_u5_U41 (.A1( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n150 ) , .A2( u1_u10_u5_n173 ) );
  AOI21_X1 u1_u10_u5_U42 (.A( u1_u10_u5_n118 ) , .B2( u1_u10_u5_n145 ) , .ZN( u1_u10_u5_n168 ) , .B1( u1_u10_u5_n186 ) );
  INV_X1 u1_u10_u5_U43 (.A( u1_u10_u5_n122 ) , .ZN( u1_u10_u5_n186 ) );
  NOR2_X1 u1_u10_u5_U44 (.A1( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n152 ) , .A2( u1_u10_u5_n176 ) );
  NOR2_X1 u1_u10_u5_U45 (.A1( u1_u10_u5_n115 ) , .ZN( u1_u10_u5_n118 ) , .A2( u1_u10_u5_n153 ) );
  NOR2_X1 u1_u10_u5_U46 (.A2( u1_u10_u5_n145 ) , .ZN( u1_u10_u5_n156 ) , .A1( u1_u10_u5_n174 ) );
  NOR2_X1 u1_u10_u5_U47 (.ZN( u1_u10_u5_n121 ) , .A2( u1_u10_u5_n145 ) , .A1( u1_u10_u5_n176 ) );
  AOI22_X1 u1_u10_u5_U48 (.ZN( u1_u10_u5_n114 ) , .A2( u1_u10_u5_n137 ) , .A1( u1_u10_u5_n145 ) , .B2( u1_u10_u5_n175 ) , .B1( u1_u10_u5_n193 ) );
  OAI211_X1 u1_u10_u5_U49 (.B( u1_u10_u5_n124 ) , .A( u1_u10_u5_n125 ) , .C2( u1_u10_u5_n126 ) , .C1( u1_u10_u5_n127 ) , .ZN( u1_u10_u5_n128 ) );
  OAI21_X1 u1_u10_u5_U5 (.B2( u1_u10_u5_n136 ) , .B1( u1_u10_u5_n137 ) , .ZN( u1_u10_u5_n138 ) , .A( u1_u10_u5_n177 ) );
  NOR3_X1 u1_u10_u5_U50 (.ZN( u1_u10_u5_n127 ) , .A1( u1_u10_u5_n136 ) , .A3( u1_u10_u5_n148 ) , .A2( u1_u10_u5_n182 ) );
  OAI21_X1 u1_u10_u5_U51 (.ZN( u1_u10_u5_n124 ) , .A( u1_u10_u5_n177 ) , .B2( u1_u10_u5_n183 ) , .B1( u1_u10_u5_n189 ) );
  OAI21_X1 u1_u10_u5_U52 (.ZN( u1_u10_u5_n125 ) , .A( u1_u10_u5_n174 ) , .B2( u1_u10_u5_n185 ) , .B1( u1_u10_u5_n190 ) );
  AOI21_X1 u1_u10_u5_U53 (.A( u1_u10_u5_n153 ) , .B2( u1_u10_u5_n154 ) , .B1( u1_u10_u5_n155 ) , .ZN( u1_u10_u5_n164 ) );
  AOI21_X1 u1_u10_u5_U54 (.ZN( u1_u10_u5_n110 ) , .B1( u1_u10_u5_n122 ) , .B2( u1_u10_u5_n139 ) , .A( u1_u10_u5_n153 ) );
  INV_X1 u1_u10_u5_U55 (.A( u1_u10_u5_n153 ) , .ZN( u1_u10_u5_n176 ) );
  INV_X1 u1_u10_u5_U56 (.A( u1_u10_u5_n126 ) , .ZN( u1_u10_u5_n173 ) );
  AND2_X1 u1_u10_u5_U57 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n147 ) );
  AND2_X1 u1_u10_u5_U58 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n148 ) );
  NAND2_X1 u1_u10_u5_U59 (.A1( u1_u10_u5_n105 ) , .A2( u1_u10_u5_n106 ) , .ZN( u1_u10_u5_n158 ) );
  INV_X1 u1_u10_u5_U6 (.A( u1_u10_u5_n135 ) , .ZN( u1_u10_u5_n178 ) );
  NAND2_X1 u1_u10_u5_U60 (.A2( u1_u10_u5_n108 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n139 ) );
  NAND2_X1 u1_u10_u5_U61 (.A1( u1_u10_u5_n106 ) , .A2( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n119 ) );
  NAND2_X1 u1_u10_u5_U62 (.A2( u1_u10_u5_n103 ) , .A1( u1_u10_u5_n105 ) , .ZN( u1_u10_u5_n140 ) );
  NAND2_X1 u1_u10_u5_U63 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n105 ) , .ZN( u1_u10_u5_n155 ) );
  NAND2_X1 u1_u10_u5_U64 (.A2( u1_u10_u5_n106 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n122 ) );
  NAND2_X1 u1_u10_u5_U65 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n106 ) , .ZN( u1_u10_u5_n115 ) );
  NAND2_X1 u1_u10_u5_U66 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n103 ) , .ZN( u1_u10_u5_n161 ) );
  NAND2_X1 u1_u10_u5_U67 (.A1( u1_u10_u5_n105 ) , .A2( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n154 ) );
  INV_X1 u1_u10_u5_U68 (.A( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n172 ) );
  NAND2_X1 u1_u10_u5_U69 (.A1( u1_u10_u5_n103 ) , .A2( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n123 ) );
  OAI22_X1 u1_u10_u5_U7 (.B2( u1_u10_u5_n149 ) , .B1( u1_u10_u5_n150 ) , .A2( u1_u10_u5_n151 ) , .A1( u1_u10_u5_n152 ) , .ZN( u1_u10_u5_n165 ) );
  NAND2_X1 u1_u10_u5_U70 (.A2( u1_u10_u5_n103 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n151 ) );
  NAND2_X1 u1_u10_u5_U71 (.A2( u1_u10_u5_n107 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n120 ) );
  NAND2_X1 u1_u10_u5_U72 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n157 ) );
  AND2_X1 u1_u10_u5_U73 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n104 ) , .ZN( u1_u10_u5_n131 ) );
  INV_X1 u1_u10_u5_U74 (.A( u1_u10_u5_n102 ) , .ZN( u1_u10_u5_n195 ) );
  OAI221_X1 u1_u10_u5_U75 (.A( u1_u10_u5_n101 ) , .ZN( u1_u10_u5_n102 ) , .C2( u1_u10_u5_n115 ) , .C1( u1_u10_u5_n126 ) , .B1( u1_u10_u5_n134 ) , .B2( u1_u10_u5_n160 ) );
  OAI21_X1 u1_u10_u5_U76 (.ZN( u1_u10_u5_n101 ) , .B1( u1_u10_u5_n137 ) , .A( u1_u10_u5_n146 ) , .B2( u1_u10_u5_n147 ) );
  NOR2_X1 u1_u10_u5_U77 (.A2( u1_u10_X_34 ) , .A1( u1_u10_X_35 ) , .ZN( u1_u10_u5_n145 ) );
  NOR2_X1 u1_u10_u5_U78 (.A2( u1_u10_X_34 ) , .ZN( u1_u10_u5_n146 ) , .A1( u1_u10_u5_n171 ) );
  NOR2_X1 u1_u10_u5_U79 (.A2( u1_u10_X_31 ) , .A1( u1_u10_X_32 ) , .ZN( u1_u10_u5_n103 ) );
  NOR3_X1 u1_u10_u5_U8 (.A2( u1_u10_u5_n147 ) , .A1( u1_u10_u5_n148 ) , .ZN( u1_u10_u5_n149 ) , .A3( u1_u10_u5_n194 ) );
  NOR2_X1 u1_u10_u5_U80 (.A2( u1_u10_X_36 ) , .ZN( u1_u10_u5_n105 ) , .A1( u1_u10_u5_n180 ) );
  NOR2_X1 u1_u10_u5_U81 (.A2( u1_u10_X_33 ) , .ZN( u1_u10_u5_n108 ) , .A1( u1_u10_u5_n170 ) );
  NOR2_X1 u1_u10_u5_U82 (.A2( u1_u10_X_33 ) , .A1( u1_u10_X_36 ) , .ZN( u1_u10_u5_n107 ) );
  NOR2_X1 u1_u10_u5_U83 (.A2( u1_u10_X_31 ) , .ZN( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n181 ) );
  NAND2_X1 u1_u10_u5_U84 (.A2( u1_u10_X_34 ) , .A1( u1_u10_X_35 ) , .ZN( u1_u10_u5_n153 ) );
  NAND2_X1 u1_u10_u5_U85 (.A1( u1_u10_X_34 ) , .ZN( u1_u10_u5_n126 ) , .A2( u1_u10_u5_n171 ) );
  AND2_X1 u1_u10_u5_U86 (.A1( u1_u10_X_31 ) , .A2( u1_u10_X_32 ) , .ZN( u1_u10_u5_n106 ) );
  AND2_X1 u1_u10_u5_U87 (.A1( u1_u10_X_31 ) , .ZN( u1_u10_u5_n109 ) , .A2( u1_u10_u5_n181 ) );
  INV_X1 u1_u10_u5_U88 (.A( u1_u10_X_33 ) , .ZN( u1_u10_u5_n180 ) );
  INV_X1 u1_u10_u5_U89 (.A( u1_u10_X_35 ) , .ZN( u1_u10_u5_n171 ) );
  NOR2_X1 u1_u10_u5_U9 (.ZN( u1_u10_u5_n135 ) , .A1( u1_u10_u5_n173 ) , .A2( u1_u10_u5_n176 ) );
  INV_X1 u1_u10_u5_U90 (.A( u1_u10_X_36 ) , .ZN( u1_u10_u5_n170 ) );
  INV_X1 u1_u10_u5_U91 (.A( u1_u10_X_32 ) , .ZN( u1_u10_u5_n181 ) );
  NAND4_X1 u1_u10_u5_U92 (.ZN( u1_out10_29 ) , .A4( u1_u10_u5_n129 ) , .A3( u1_u10_u5_n130 ) , .A2( u1_u10_u5_n168 ) , .A1( u1_u10_u5_n196 ) );
  AOI221_X1 u1_u10_u5_U93 (.A( u1_u10_u5_n128 ) , .ZN( u1_u10_u5_n129 ) , .C2( u1_u10_u5_n132 ) , .B2( u1_u10_u5_n159 ) , .B1( u1_u10_u5_n176 ) , .C1( u1_u10_u5_n184 ) );
  AOI222_X1 u1_u10_u5_U94 (.ZN( u1_u10_u5_n130 ) , .A2( u1_u10_u5_n146 ) , .B1( u1_u10_u5_n147 ) , .C2( u1_u10_u5_n175 ) , .B2( u1_u10_u5_n179 ) , .A1( u1_u10_u5_n188 ) , .C1( u1_u10_u5_n194 ) );
  NAND4_X1 u1_u10_u5_U95 (.ZN( u1_out10_19 ) , .A4( u1_u10_u5_n166 ) , .A3( u1_u10_u5_n167 ) , .A2( u1_u10_u5_n168 ) , .A1( u1_u10_u5_n169 ) );
  AOI22_X1 u1_u10_u5_U96 (.B2( u1_u10_u5_n145 ) , .A2( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n167 ) , .B1( u1_u10_u5_n182 ) , .A1( u1_u10_u5_n189 ) );
  NOR4_X1 u1_u10_u5_U97 (.A4( u1_u10_u5_n162 ) , .A3( u1_u10_u5_n163 ) , .A2( u1_u10_u5_n164 ) , .A1( u1_u10_u5_n165 ) , .ZN( u1_u10_u5_n166 ) );
  NAND4_X1 u1_u10_u5_U98 (.ZN( u1_out10_11 ) , .A4( u1_u10_u5_n143 ) , .A3( u1_u10_u5_n144 ) , .A2( u1_u10_u5_n169 ) , .A1( u1_u10_u5_n196 ) );
  AOI22_X1 u1_u10_u5_U99 (.A2( u1_u10_u5_n132 ) , .ZN( u1_u10_u5_n144 ) , .B2( u1_u10_u5_n145 ) , .B1( u1_u10_u5_n184 ) , .A1( u1_u10_u5_n194 ) );
  AOI22_X1 u1_u10_u6_U10 (.A2( u1_u10_u6_n151 ) , .B2( u1_u10_u6_n161 ) , .A1( u1_u10_u6_n167 ) , .B1( u1_u10_u6_n170 ) , .ZN( u1_u10_u6_n89 ) );
  AOI21_X1 u1_u10_u6_U11 (.B1( u1_u10_u6_n107 ) , .B2( u1_u10_u6_n132 ) , .A( u1_u10_u6_n158 ) , .ZN( u1_u10_u6_n88 ) );
  AOI21_X1 u1_u10_u6_U12 (.B2( u1_u10_u6_n147 ) , .B1( u1_u10_u6_n148 ) , .ZN( u1_u10_u6_n149 ) , .A( u1_u10_u6_n158 ) );
  AOI21_X1 u1_u10_u6_U13 (.ZN( u1_u10_u6_n106 ) , .A( u1_u10_u6_n142 ) , .B2( u1_u10_u6_n159 ) , .B1( u1_u10_u6_n164 ) );
  INV_X1 u1_u10_u6_U14 (.A( u1_u10_u6_n155 ) , .ZN( u1_u10_u6_n161 ) );
  INV_X1 u1_u10_u6_U15 (.A( u1_u10_u6_n128 ) , .ZN( u1_u10_u6_n164 ) );
  NAND2_X1 u1_u10_u6_U16 (.ZN( u1_u10_u6_n110 ) , .A1( u1_u10_u6_n122 ) , .A2( u1_u10_u6_n129 ) );
  NAND2_X1 u1_u10_u6_U17 (.ZN( u1_u10_u6_n124 ) , .A2( u1_u10_u6_n146 ) , .A1( u1_u10_u6_n148 ) );
  INV_X1 u1_u10_u6_U18 (.A( u1_u10_u6_n132 ) , .ZN( u1_u10_u6_n171 ) );
  AND2_X1 u1_u10_u6_U19 (.A1( u1_u10_u6_n100 ) , .ZN( u1_u10_u6_n130 ) , .A2( u1_u10_u6_n147 ) );
  INV_X1 u1_u10_u6_U20 (.A( u1_u10_u6_n127 ) , .ZN( u1_u10_u6_n173 ) );
  INV_X1 u1_u10_u6_U21 (.A( u1_u10_u6_n121 ) , .ZN( u1_u10_u6_n167 ) );
  INV_X1 u1_u10_u6_U22 (.A( u1_u10_u6_n100 ) , .ZN( u1_u10_u6_n169 ) );
  INV_X1 u1_u10_u6_U23 (.A( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n170 ) );
  INV_X1 u1_u10_u6_U24 (.A( u1_u10_u6_n113 ) , .ZN( u1_u10_u6_n168 ) );
  AND2_X1 u1_u10_u6_U25 (.A1( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n119 ) , .ZN( u1_u10_u6_n133 ) );
  AND2_X1 u1_u10_u6_U26 (.A2( u1_u10_u6_n121 ) , .A1( u1_u10_u6_n122 ) , .ZN( u1_u10_u6_n131 ) );
  AND3_X1 u1_u10_u6_U27 (.ZN( u1_u10_u6_n120 ) , .A2( u1_u10_u6_n127 ) , .A1( u1_u10_u6_n132 ) , .A3( u1_u10_u6_n145 ) );
  INV_X1 u1_u10_u6_U28 (.A( u1_u10_u6_n146 ) , .ZN( u1_u10_u6_n163 ) );
  AOI222_X1 u1_u10_u6_U29 (.ZN( u1_u10_u6_n114 ) , .A1( u1_u10_u6_n118 ) , .A2( u1_u10_u6_n126 ) , .B2( u1_u10_u6_n151 ) , .C2( u1_u10_u6_n159 ) , .C1( u1_u10_u6_n168 ) , .B1( u1_u10_u6_n169 ) );
  INV_X1 u1_u10_u6_U3 (.A( u1_u10_u6_n110 ) , .ZN( u1_u10_u6_n166 ) );
  NOR2_X1 u1_u10_u6_U30 (.A1( u1_u10_u6_n162 ) , .A2( u1_u10_u6_n165 ) , .ZN( u1_u10_u6_n98 ) );
  AOI211_X1 u1_u10_u6_U31 (.B( u1_u10_u6_n134 ) , .A( u1_u10_u6_n135 ) , .C1( u1_u10_u6_n136 ) , .ZN( u1_u10_u6_n137 ) , .C2( u1_u10_u6_n151 ) );
  NAND4_X1 u1_u10_u6_U32 (.A4( u1_u10_u6_n127 ) , .A3( u1_u10_u6_n128 ) , .A2( u1_u10_u6_n129 ) , .A1( u1_u10_u6_n130 ) , .ZN( u1_u10_u6_n136 ) );
  AOI21_X1 u1_u10_u6_U33 (.B2( u1_u10_u6_n132 ) , .B1( u1_u10_u6_n133 ) , .ZN( u1_u10_u6_n134 ) , .A( u1_u10_u6_n158 ) );
  AOI21_X1 u1_u10_u6_U34 (.B1( u1_u10_u6_n131 ) , .ZN( u1_u10_u6_n135 ) , .A( u1_u10_u6_n144 ) , .B2( u1_u10_u6_n146 ) );
  NAND2_X1 u1_u10_u6_U35 (.A1( u1_u10_u6_n144 ) , .ZN( u1_u10_u6_n151 ) , .A2( u1_u10_u6_n158 ) );
  NAND2_X1 u1_u10_u6_U36 (.ZN( u1_u10_u6_n132 ) , .A1( u1_u10_u6_n91 ) , .A2( u1_u10_u6_n97 ) );
  AOI22_X1 u1_u10_u6_U37 (.B2( u1_u10_u6_n110 ) , .B1( u1_u10_u6_n111 ) , .A1( u1_u10_u6_n112 ) , .ZN( u1_u10_u6_n115 ) , .A2( u1_u10_u6_n161 ) );
  NAND4_X1 u1_u10_u6_U38 (.A3( u1_u10_u6_n109 ) , .ZN( u1_u10_u6_n112 ) , .A4( u1_u10_u6_n132 ) , .A2( u1_u10_u6_n147 ) , .A1( u1_u10_u6_n166 ) );
  NOR2_X1 u1_u10_u6_U39 (.ZN( u1_u10_u6_n109 ) , .A1( u1_u10_u6_n170 ) , .A2( u1_u10_u6_n173 ) );
  INV_X1 u1_u10_u6_U4 (.A( u1_u10_u6_n142 ) , .ZN( u1_u10_u6_n174 ) );
  NOR2_X1 u1_u10_u6_U40 (.A2( u1_u10_u6_n126 ) , .ZN( u1_u10_u6_n155 ) , .A1( u1_u10_u6_n160 ) );
  NAND2_X1 u1_u10_u6_U41 (.ZN( u1_u10_u6_n146 ) , .A2( u1_u10_u6_n94 ) , .A1( u1_u10_u6_n99 ) );
  AOI21_X1 u1_u10_u6_U42 (.A( u1_u10_u6_n144 ) , .B2( u1_u10_u6_n145 ) , .B1( u1_u10_u6_n146 ) , .ZN( u1_u10_u6_n150 ) );
  INV_X1 u1_u10_u6_U43 (.A( u1_u10_u6_n111 ) , .ZN( u1_u10_u6_n158 ) );
  NAND2_X1 u1_u10_u6_U44 (.ZN( u1_u10_u6_n127 ) , .A1( u1_u10_u6_n91 ) , .A2( u1_u10_u6_n92 ) );
  NAND2_X1 u1_u10_u6_U45 (.ZN( u1_u10_u6_n129 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n96 ) );
  INV_X1 u1_u10_u6_U46 (.A( u1_u10_u6_n144 ) , .ZN( u1_u10_u6_n159 ) );
  NAND2_X1 u1_u10_u6_U47 (.ZN( u1_u10_u6_n145 ) , .A2( u1_u10_u6_n97 ) , .A1( u1_u10_u6_n98 ) );
  NAND2_X1 u1_u10_u6_U48 (.ZN( u1_u10_u6_n148 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n94 ) );
  NAND2_X1 u1_u10_u6_U49 (.ZN( u1_u10_u6_n108 ) , .A2( u1_u10_u6_n139 ) , .A1( u1_u10_u6_n144 ) );
  NAND2_X1 u1_u10_u6_U5 (.A2( u1_u10_u6_n143 ) , .ZN( u1_u10_u6_n152 ) , .A1( u1_u10_u6_n166 ) );
  NAND2_X1 u1_u10_u6_U50 (.ZN( u1_u10_u6_n121 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n97 ) );
  NAND2_X1 u1_u10_u6_U51 (.ZN( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n95 ) );
  AND2_X1 u1_u10_u6_U52 (.ZN( u1_u10_u6_n118 ) , .A2( u1_u10_u6_n91 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U53 (.ZN( u1_u10_u6_n147 ) , .A2( u1_u10_u6_n98 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U54 (.ZN( u1_u10_u6_n128 ) , .A1( u1_u10_u6_n94 ) , .A2( u1_u10_u6_n96 ) );
  NAND2_X1 u1_u10_u6_U55 (.ZN( u1_u10_u6_n119 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U56 (.ZN( u1_u10_u6_n123 ) , .A2( u1_u10_u6_n91 ) , .A1( u1_u10_u6_n96 ) );
  NAND2_X1 u1_u10_u6_U57 (.ZN( u1_u10_u6_n100 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n98 ) );
  NAND2_X1 u1_u10_u6_U58 (.ZN( u1_u10_u6_n122 ) , .A1( u1_u10_u6_n94 ) , .A2( u1_u10_u6_n97 ) );
  INV_X1 u1_u10_u6_U59 (.A( u1_u10_u6_n139 ) , .ZN( u1_u10_u6_n160 ) );
  AOI22_X1 u1_u10_u6_U6 (.B2( u1_u10_u6_n101 ) , .A1( u1_u10_u6_n102 ) , .ZN( u1_u10_u6_n103 ) , .B1( u1_u10_u6_n160 ) , .A2( u1_u10_u6_n161 ) );
  NAND2_X1 u1_u10_u6_U60 (.ZN( u1_u10_u6_n113 ) , .A1( u1_u10_u6_n96 ) , .A2( u1_u10_u6_n98 ) );
  NOR2_X1 u1_u10_u6_U61 (.A2( u1_u10_X_40 ) , .A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n126 ) );
  NOR2_X1 u1_u10_u6_U62 (.A2( u1_u10_X_39 ) , .A1( u1_u10_X_42 ) , .ZN( u1_u10_u6_n92 ) );
  NOR2_X1 u1_u10_u6_U63 (.A2( u1_u10_X_39 ) , .A1( u1_u10_u6_n156 ) , .ZN( u1_u10_u6_n97 ) );
  NOR2_X1 u1_u10_u6_U64 (.A2( u1_u10_X_38 ) , .A1( u1_u10_u6_n165 ) , .ZN( u1_u10_u6_n95 ) );
  NOR2_X1 u1_u10_u6_U65 (.A2( u1_u10_X_41 ) , .ZN( u1_u10_u6_n111 ) , .A1( u1_u10_u6_n157 ) );
  NOR2_X1 u1_u10_u6_U66 (.A2( u1_u10_X_37 ) , .A1( u1_u10_u6_n162 ) , .ZN( u1_u10_u6_n94 ) );
  NOR2_X1 u1_u10_u6_U67 (.A2( u1_u10_X_37 ) , .A1( u1_u10_X_38 ) , .ZN( u1_u10_u6_n91 ) );
  NAND2_X1 u1_u10_u6_U68 (.A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n144 ) , .A2( u1_u10_u6_n157 ) );
  NAND2_X1 u1_u10_u6_U69 (.A2( u1_u10_X_40 ) , .A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n139 ) );
  NOR2_X1 u1_u10_u6_U7 (.A1( u1_u10_u6_n118 ) , .ZN( u1_u10_u6_n143 ) , .A2( u1_u10_u6_n168 ) );
  AND2_X1 u1_u10_u6_U70 (.A1( u1_u10_X_39 ) , .A2( u1_u10_u6_n156 ) , .ZN( u1_u10_u6_n96 ) );
  AND2_X1 u1_u10_u6_U71 (.A1( u1_u10_X_39 ) , .A2( u1_u10_X_42 ) , .ZN( u1_u10_u6_n99 ) );
  INV_X1 u1_u10_u6_U72 (.A( u1_u10_X_40 ) , .ZN( u1_u10_u6_n157 ) );
  INV_X1 u1_u10_u6_U73 (.A( u1_u10_X_37 ) , .ZN( u1_u10_u6_n165 ) );
  INV_X1 u1_u10_u6_U74 (.A( u1_u10_X_38 ) , .ZN( u1_u10_u6_n162 ) );
  INV_X1 u1_u10_u6_U75 (.A( u1_u10_X_42 ) , .ZN( u1_u10_u6_n156 ) );
  NAND4_X1 u1_u10_u6_U76 (.ZN( u1_out10_32 ) , .A4( u1_u10_u6_n103 ) , .A3( u1_u10_u6_n104 ) , .A2( u1_u10_u6_n105 ) , .A1( u1_u10_u6_n106 ) );
  AOI22_X1 u1_u10_u6_U77 (.ZN( u1_u10_u6_n105 ) , .A2( u1_u10_u6_n108 ) , .A1( u1_u10_u6_n118 ) , .B2( u1_u10_u6_n126 ) , .B1( u1_u10_u6_n171 ) );
  AOI22_X1 u1_u10_u6_U78 (.ZN( u1_u10_u6_n104 ) , .A1( u1_u10_u6_n111 ) , .B1( u1_u10_u6_n124 ) , .B2( u1_u10_u6_n151 ) , .A2( u1_u10_u6_n93 ) );
  NAND4_X1 u1_u10_u6_U79 (.ZN( u1_out10_12 ) , .A4( u1_u10_u6_n114 ) , .A3( u1_u10_u6_n115 ) , .A2( u1_u10_u6_n116 ) , .A1( u1_u10_u6_n117 ) );
  INV_X1 u1_u10_u6_U8 (.ZN( u1_u10_u6_n172 ) , .A( u1_u10_u6_n88 ) );
  OAI22_X1 u1_u10_u6_U80 (.B2( u1_u10_u6_n111 ) , .ZN( u1_u10_u6_n116 ) , .B1( u1_u10_u6_n126 ) , .A2( u1_u10_u6_n164 ) , .A1( u1_u10_u6_n167 ) );
  OAI21_X1 u1_u10_u6_U81 (.A( u1_u10_u6_n108 ) , .ZN( u1_u10_u6_n117 ) , .B2( u1_u10_u6_n141 ) , .B1( u1_u10_u6_n163 ) );
  OAI211_X1 u1_u10_u6_U82 (.ZN( u1_out10_7 ) , .B( u1_u10_u6_n153 ) , .C2( u1_u10_u6_n154 ) , .C1( u1_u10_u6_n155 ) , .A( u1_u10_u6_n174 ) );
  NOR3_X1 u1_u10_u6_U83 (.A1( u1_u10_u6_n141 ) , .ZN( u1_u10_u6_n154 ) , .A3( u1_u10_u6_n164 ) , .A2( u1_u10_u6_n171 ) );
  AOI211_X1 u1_u10_u6_U84 (.B( u1_u10_u6_n149 ) , .A( u1_u10_u6_n150 ) , .C2( u1_u10_u6_n151 ) , .C1( u1_u10_u6_n152 ) , .ZN( u1_u10_u6_n153 ) );
  OAI211_X1 u1_u10_u6_U85 (.ZN( u1_out10_22 ) , .B( u1_u10_u6_n137 ) , .A( u1_u10_u6_n138 ) , .C2( u1_u10_u6_n139 ) , .C1( u1_u10_u6_n140 ) );
  AOI22_X1 u1_u10_u6_U86 (.B1( u1_u10_u6_n124 ) , .A2( u1_u10_u6_n125 ) , .A1( u1_u10_u6_n126 ) , .ZN( u1_u10_u6_n138 ) , .B2( u1_u10_u6_n161 ) );
  AND4_X1 u1_u10_u6_U87 (.A3( u1_u10_u6_n119 ) , .A1( u1_u10_u6_n120 ) , .A4( u1_u10_u6_n129 ) , .ZN( u1_u10_u6_n140 ) , .A2( u1_u10_u6_n143 ) );
  NAND3_X1 u1_u10_u6_U88 (.A2( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n125 ) , .A1( u1_u10_u6_n130 ) , .A3( u1_u10_u6_n131 ) );
  NAND3_X1 u1_u10_u6_U89 (.A3( u1_u10_u6_n133 ) , .ZN( u1_u10_u6_n141 ) , .A1( u1_u10_u6_n145 ) , .A2( u1_u10_u6_n148 ) );
  OAI21_X1 u1_u10_u6_U9 (.A( u1_u10_u6_n159 ) , .B1( u1_u10_u6_n169 ) , .B2( u1_u10_u6_n173 ) , .ZN( u1_u10_u6_n90 ) );
  NAND3_X1 u1_u10_u6_U90 (.ZN( u1_u10_u6_n101 ) , .A3( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n121 ) , .A1( u1_u10_u6_n127 ) );
  NAND3_X1 u1_u10_u6_U91 (.ZN( u1_u10_u6_n102 ) , .A3( u1_u10_u6_n130 ) , .A2( u1_u10_u6_n145 ) , .A1( u1_u10_u6_n166 ) );
  NAND3_X1 u1_u10_u6_U92 (.A3( u1_u10_u6_n113 ) , .A1( u1_u10_u6_n119 ) , .A2( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n93 ) );
  NAND3_X1 u1_u10_u6_U93 (.ZN( u1_u10_u6_n142 ) , .A2( u1_u10_u6_n172 ) , .A3( u1_u10_u6_n89 ) , .A1( u1_u10_u6_n90 ) );
  AND3_X1 u1_u10_u7_U10 (.A3( u1_u10_u7_n110 ) , .A2( u1_u10_u7_n127 ) , .A1( u1_u10_u7_n132 ) , .ZN( u1_u10_u7_n92 ) );
  OAI21_X1 u1_u10_u7_U11 (.A( u1_u10_u7_n161 ) , .B1( u1_u10_u7_n168 ) , .B2( u1_u10_u7_n173 ) , .ZN( u1_u10_u7_n91 ) );
  AOI211_X1 u1_u10_u7_U12 (.A( u1_u10_u7_n117 ) , .ZN( u1_u10_u7_n118 ) , .C2( u1_u10_u7_n126 ) , .C1( u1_u10_u7_n177 ) , .B( u1_u10_u7_n180 ) );
  OAI22_X1 u1_u10_u7_U13 (.B1( u1_u10_u7_n115 ) , .ZN( u1_u10_u7_n117 ) , .A2( u1_u10_u7_n133 ) , .A1( u1_u10_u7_n137 ) , .B2( u1_u10_u7_n162 ) );
  INV_X1 u1_u10_u7_U14 (.A( u1_u10_u7_n116 ) , .ZN( u1_u10_u7_n180 ) );
  NOR3_X1 u1_u10_u7_U15 (.ZN( u1_u10_u7_n115 ) , .A3( u1_u10_u7_n145 ) , .A2( u1_u10_u7_n168 ) , .A1( u1_u10_u7_n169 ) );
  OAI211_X1 u1_u10_u7_U16 (.B( u1_u10_u7_n122 ) , .A( u1_u10_u7_n123 ) , .C2( u1_u10_u7_n124 ) , .ZN( u1_u10_u7_n154 ) , .C1( u1_u10_u7_n162 ) );
  AOI222_X1 u1_u10_u7_U17 (.ZN( u1_u10_u7_n122 ) , .C2( u1_u10_u7_n126 ) , .C1( u1_u10_u7_n145 ) , .B1( u1_u10_u7_n161 ) , .A2( u1_u10_u7_n165 ) , .B2( u1_u10_u7_n170 ) , .A1( u1_u10_u7_n176 ) );
  INV_X1 u1_u10_u7_U18 (.A( u1_u10_u7_n133 ) , .ZN( u1_u10_u7_n176 ) );
  NOR3_X1 u1_u10_u7_U19 (.A2( u1_u10_u7_n134 ) , .A1( u1_u10_u7_n135 ) , .ZN( u1_u10_u7_n136 ) , .A3( u1_u10_u7_n171 ) );
  NOR2_X1 u1_u10_u7_U20 (.A1( u1_u10_u7_n130 ) , .A2( u1_u10_u7_n134 ) , .ZN( u1_u10_u7_n153 ) );
  INV_X1 u1_u10_u7_U21 (.A( u1_u10_u7_n101 ) , .ZN( u1_u10_u7_n165 ) );
  NOR2_X1 u1_u10_u7_U22 (.ZN( u1_u10_u7_n111 ) , .A2( u1_u10_u7_n134 ) , .A1( u1_u10_u7_n169 ) );
  AOI21_X1 u1_u10_u7_U23 (.ZN( u1_u10_u7_n104 ) , .B2( u1_u10_u7_n112 ) , .B1( u1_u10_u7_n127 ) , .A( u1_u10_u7_n164 ) );
  AOI21_X1 u1_u10_u7_U24 (.ZN( u1_u10_u7_n106 ) , .B1( u1_u10_u7_n133 ) , .B2( u1_u10_u7_n146 ) , .A( u1_u10_u7_n162 ) );
  AOI21_X1 u1_u10_u7_U25 (.A( u1_u10_u7_n101 ) , .ZN( u1_u10_u7_n107 ) , .B2( u1_u10_u7_n128 ) , .B1( u1_u10_u7_n175 ) );
  INV_X1 u1_u10_u7_U26 (.A( u1_u10_u7_n138 ) , .ZN( u1_u10_u7_n171 ) );
  INV_X1 u1_u10_u7_U27 (.A( u1_u10_u7_n131 ) , .ZN( u1_u10_u7_n177 ) );
  INV_X1 u1_u10_u7_U28 (.A( u1_u10_u7_n110 ) , .ZN( u1_u10_u7_n174 ) );
  NAND2_X1 u1_u10_u7_U29 (.A1( u1_u10_u7_n129 ) , .A2( u1_u10_u7_n132 ) , .ZN( u1_u10_u7_n149 ) );
  OAI21_X1 u1_u10_u7_U3 (.ZN( u1_u10_u7_n159 ) , .A( u1_u10_u7_n165 ) , .B2( u1_u10_u7_n171 ) , .B1( u1_u10_u7_n174 ) );
  NAND2_X1 u1_u10_u7_U30 (.A1( u1_u10_u7_n113 ) , .A2( u1_u10_u7_n124 ) , .ZN( u1_u10_u7_n130 ) );
  INV_X1 u1_u10_u7_U31 (.A( u1_u10_u7_n112 ) , .ZN( u1_u10_u7_n173 ) );
  INV_X1 u1_u10_u7_U32 (.A( u1_u10_u7_n128 ) , .ZN( u1_u10_u7_n168 ) );
  INV_X1 u1_u10_u7_U33 (.A( u1_u10_u7_n148 ) , .ZN( u1_u10_u7_n169 ) );
  INV_X1 u1_u10_u7_U34 (.A( u1_u10_u7_n127 ) , .ZN( u1_u10_u7_n179 ) );
  NOR2_X1 u1_u10_u7_U35 (.ZN( u1_u10_u7_n101 ) , .A2( u1_u10_u7_n150 ) , .A1( u1_u10_u7_n156 ) );
  AOI211_X1 u1_u10_u7_U36 (.B( u1_u10_u7_n154 ) , .A( u1_u10_u7_n155 ) , .C1( u1_u10_u7_n156 ) , .ZN( u1_u10_u7_n157 ) , .C2( u1_u10_u7_n172 ) );
  INV_X1 u1_u10_u7_U37 (.A( u1_u10_u7_n153 ) , .ZN( u1_u10_u7_n172 ) );
  AOI211_X1 u1_u10_u7_U38 (.B( u1_u10_u7_n139 ) , .A( u1_u10_u7_n140 ) , .C2( u1_u10_u7_n141 ) , .ZN( u1_u10_u7_n142 ) , .C1( u1_u10_u7_n156 ) );
  NAND4_X1 u1_u10_u7_U39 (.A3( u1_u10_u7_n127 ) , .A2( u1_u10_u7_n128 ) , .A1( u1_u10_u7_n129 ) , .ZN( u1_u10_u7_n141 ) , .A4( u1_u10_u7_n147 ) );
  INV_X1 u1_u10_u7_U4 (.A( u1_u10_u7_n111 ) , .ZN( u1_u10_u7_n170 ) );
  AOI21_X1 u1_u10_u7_U40 (.A( u1_u10_u7_n137 ) , .B1( u1_u10_u7_n138 ) , .ZN( u1_u10_u7_n139 ) , .B2( u1_u10_u7_n146 ) );
  OAI22_X1 u1_u10_u7_U41 (.B1( u1_u10_u7_n136 ) , .ZN( u1_u10_u7_n140 ) , .A1( u1_u10_u7_n153 ) , .B2( u1_u10_u7_n162 ) , .A2( u1_u10_u7_n164 ) );
  AOI21_X1 u1_u10_u7_U42 (.ZN( u1_u10_u7_n123 ) , .B1( u1_u10_u7_n165 ) , .B2( u1_u10_u7_n177 ) , .A( u1_u10_u7_n97 ) );
  AOI21_X1 u1_u10_u7_U43 (.B2( u1_u10_u7_n113 ) , .B1( u1_u10_u7_n124 ) , .A( u1_u10_u7_n125 ) , .ZN( u1_u10_u7_n97 ) );
  INV_X1 u1_u10_u7_U44 (.A( u1_u10_u7_n125 ) , .ZN( u1_u10_u7_n161 ) );
  INV_X1 u1_u10_u7_U45 (.A( u1_u10_u7_n152 ) , .ZN( u1_u10_u7_n162 ) );
  AOI22_X1 u1_u10_u7_U46 (.A2( u1_u10_u7_n114 ) , .ZN( u1_u10_u7_n119 ) , .B1( u1_u10_u7_n130 ) , .A1( u1_u10_u7_n156 ) , .B2( u1_u10_u7_n165 ) );
  NAND2_X1 u1_u10_u7_U47 (.A2( u1_u10_u7_n112 ) , .ZN( u1_u10_u7_n114 ) , .A1( u1_u10_u7_n175 ) );
  AND2_X1 u1_u10_u7_U48 (.ZN( u1_u10_u7_n145 ) , .A2( u1_u10_u7_n98 ) , .A1( u1_u10_u7_n99 ) );
  NOR2_X1 u1_u10_u7_U49 (.ZN( u1_u10_u7_n137 ) , .A1( u1_u10_u7_n150 ) , .A2( u1_u10_u7_n161 ) );
  INV_X1 u1_u10_u7_U5 (.A( u1_u10_u7_n149 ) , .ZN( u1_u10_u7_n175 ) );
  AOI21_X1 u1_u10_u7_U50 (.ZN( u1_u10_u7_n105 ) , .B2( u1_u10_u7_n110 ) , .A( u1_u10_u7_n125 ) , .B1( u1_u10_u7_n147 ) );
  NAND2_X1 u1_u10_u7_U51 (.ZN( u1_u10_u7_n146 ) , .A1( u1_u10_u7_n95 ) , .A2( u1_u10_u7_n98 ) );
  NAND2_X1 u1_u10_u7_U52 (.A2( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n147 ) , .A1( u1_u10_u7_n93 ) );
  NAND2_X1 u1_u10_u7_U53 (.A1( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n127 ) , .A2( u1_u10_u7_n99 ) );
  OR2_X1 u1_u10_u7_U54 (.ZN( u1_u10_u7_n126 ) , .A2( u1_u10_u7_n152 ) , .A1( u1_u10_u7_n156 ) );
  NAND2_X1 u1_u10_u7_U55 (.A2( u1_u10_u7_n102 ) , .A1( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n133 ) );
  NAND2_X1 u1_u10_u7_U56 (.ZN( u1_u10_u7_n112 ) , .A2( u1_u10_u7_n96 ) , .A1( u1_u10_u7_n99 ) );
  NAND2_X1 u1_u10_u7_U57 (.A2( u1_u10_u7_n102 ) , .ZN( u1_u10_u7_n128 ) , .A1( u1_u10_u7_n98 ) );
  NAND2_X1 u1_u10_u7_U58 (.A1( u1_u10_u7_n100 ) , .ZN( u1_u10_u7_n113 ) , .A2( u1_u10_u7_n93 ) );
  NAND2_X1 u1_u10_u7_U59 (.A2( u1_u10_u7_n102 ) , .ZN( u1_u10_u7_n124 ) , .A1( u1_u10_u7_n96 ) );
  INV_X1 u1_u10_u7_U6 (.A( u1_u10_u7_n154 ) , .ZN( u1_u10_u7_n178 ) );
  NAND2_X1 u1_u10_u7_U60 (.ZN( u1_u10_u7_n110 ) , .A1( u1_u10_u7_n95 ) , .A2( u1_u10_u7_n96 ) );
  INV_X1 u1_u10_u7_U61 (.A( u1_u10_u7_n150 ) , .ZN( u1_u10_u7_n164 ) );
  AND2_X1 u1_u10_u7_U62 (.ZN( u1_u10_u7_n134 ) , .A1( u1_u10_u7_n93 ) , .A2( u1_u10_u7_n98 ) );
  NAND2_X1 u1_u10_u7_U63 (.A1( u1_u10_u7_n100 ) , .A2( u1_u10_u7_n102 ) , .ZN( u1_u10_u7_n129 ) );
  NAND2_X1 u1_u10_u7_U64 (.A2( u1_u10_u7_n103 ) , .ZN( u1_u10_u7_n131 ) , .A1( u1_u10_u7_n95 ) );
  NAND2_X1 u1_u10_u7_U65 (.A1( u1_u10_u7_n100 ) , .ZN( u1_u10_u7_n138 ) , .A2( u1_u10_u7_n99 ) );
  NAND2_X1 u1_u10_u7_U66 (.ZN( u1_u10_u7_n132 ) , .A1( u1_u10_u7_n93 ) , .A2( u1_u10_u7_n96 ) );
  NAND2_X1 u1_u10_u7_U67 (.A1( u1_u10_u7_n100 ) , .ZN( u1_u10_u7_n148 ) , .A2( u1_u10_u7_n95 ) );
  NOR2_X1 u1_u10_u7_U68 (.A2( u1_u10_X_47 ) , .ZN( u1_u10_u7_n150 ) , .A1( u1_u10_u7_n163 ) );
  NOR2_X1 u1_u10_u7_U69 (.A2( u1_u10_X_43 ) , .A1( u1_u10_X_44 ) , .ZN( u1_u10_u7_n103 ) );
  AOI211_X1 u1_u10_u7_U7 (.ZN( u1_u10_u7_n116 ) , .A( u1_u10_u7_n155 ) , .C1( u1_u10_u7_n161 ) , .C2( u1_u10_u7_n171 ) , .B( u1_u10_u7_n94 ) );
  NOR2_X1 u1_u10_u7_U70 (.A2( u1_u10_X_48 ) , .A1( u1_u10_u7_n166 ) , .ZN( u1_u10_u7_n95 ) );
  NOR2_X1 u1_u10_u7_U71 (.A2( u1_u10_X_45 ) , .A1( u1_u10_X_48 ) , .ZN( u1_u10_u7_n99 ) );
  NOR2_X1 u1_u10_u7_U72 (.A2( u1_u10_X_44 ) , .A1( u1_u10_u7_n167 ) , .ZN( u1_u10_u7_n98 ) );
  NOR2_X1 u1_u10_u7_U73 (.A2( u1_u10_X_46 ) , .A1( u1_u10_X_47 ) , .ZN( u1_u10_u7_n152 ) );
  AND2_X1 u1_u10_u7_U74 (.A1( u1_u10_X_47 ) , .ZN( u1_u10_u7_n156 ) , .A2( u1_u10_u7_n163 ) );
  NAND2_X1 u1_u10_u7_U75 (.A2( u1_u10_X_46 ) , .A1( u1_u10_X_47 ) , .ZN( u1_u10_u7_n125 ) );
  AND2_X1 u1_u10_u7_U76 (.A2( u1_u10_X_45 ) , .A1( u1_u10_X_48 ) , .ZN( u1_u10_u7_n102 ) );
  AND2_X1 u1_u10_u7_U77 (.A2( u1_u10_X_43 ) , .A1( u1_u10_X_44 ) , .ZN( u1_u10_u7_n96 ) );
  AND2_X1 u1_u10_u7_U78 (.A1( u1_u10_X_44 ) , .ZN( u1_u10_u7_n100 ) , .A2( u1_u10_u7_n167 ) );
  AND2_X1 u1_u10_u7_U79 (.A1( u1_u10_X_48 ) , .A2( u1_u10_u7_n166 ) , .ZN( u1_u10_u7_n93 ) );
  OAI222_X1 u1_u10_u7_U8 (.C2( u1_u10_u7_n101 ) , .B2( u1_u10_u7_n111 ) , .A1( u1_u10_u7_n113 ) , .C1( u1_u10_u7_n146 ) , .A2( u1_u10_u7_n162 ) , .B1( u1_u10_u7_n164 ) , .ZN( u1_u10_u7_n94 ) );
  INV_X1 u1_u10_u7_U80 (.A( u1_u10_X_46 ) , .ZN( u1_u10_u7_n163 ) );
  INV_X1 u1_u10_u7_U81 (.A( u1_u10_X_43 ) , .ZN( u1_u10_u7_n167 ) );
  INV_X1 u1_u10_u7_U82 (.A( u1_u10_X_45 ) , .ZN( u1_u10_u7_n166 ) );
  NAND4_X1 u1_u10_u7_U83 (.ZN( u1_out10_27 ) , .A4( u1_u10_u7_n118 ) , .A3( u1_u10_u7_n119 ) , .A2( u1_u10_u7_n120 ) , .A1( u1_u10_u7_n121 ) );
  OAI21_X1 u1_u10_u7_U84 (.ZN( u1_u10_u7_n121 ) , .B2( u1_u10_u7_n145 ) , .A( u1_u10_u7_n150 ) , .B1( u1_u10_u7_n174 ) );
  OAI21_X1 u1_u10_u7_U85 (.ZN( u1_u10_u7_n120 ) , .A( u1_u10_u7_n161 ) , .B2( u1_u10_u7_n170 ) , .B1( u1_u10_u7_n179 ) );
  NAND4_X1 u1_u10_u7_U86 (.ZN( u1_out10_21 ) , .A4( u1_u10_u7_n157 ) , .A3( u1_u10_u7_n158 ) , .A2( u1_u10_u7_n159 ) , .A1( u1_u10_u7_n160 ) );
  OAI21_X1 u1_u10_u7_U87 (.B1( u1_u10_u7_n145 ) , .ZN( u1_u10_u7_n160 ) , .A( u1_u10_u7_n161 ) , .B2( u1_u10_u7_n177 ) );
  AOI22_X1 u1_u10_u7_U88 (.B2( u1_u10_u7_n149 ) , .B1( u1_u10_u7_n150 ) , .A2( u1_u10_u7_n151 ) , .A1( u1_u10_u7_n152 ) , .ZN( u1_u10_u7_n158 ) );
  NAND4_X1 u1_u10_u7_U89 (.ZN( u1_out10_15 ) , .A4( u1_u10_u7_n142 ) , .A3( u1_u10_u7_n143 ) , .A2( u1_u10_u7_n144 ) , .A1( u1_u10_u7_n178 ) );
  OAI221_X1 u1_u10_u7_U9 (.C1( u1_u10_u7_n101 ) , .C2( u1_u10_u7_n147 ) , .ZN( u1_u10_u7_n155 ) , .B2( u1_u10_u7_n162 ) , .A( u1_u10_u7_n91 ) , .B1( u1_u10_u7_n92 ) );
  OR2_X1 u1_u10_u7_U90 (.A2( u1_u10_u7_n125 ) , .A1( u1_u10_u7_n129 ) , .ZN( u1_u10_u7_n144 ) );
  AOI22_X1 u1_u10_u7_U91 (.A2( u1_u10_u7_n126 ) , .ZN( u1_u10_u7_n143 ) , .B2( u1_u10_u7_n165 ) , .B1( u1_u10_u7_n173 ) , .A1( u1_u10_u7_n174 ) );
  NAND4_X1 u1_u10_u7_U92 (.ZN( u1_out10_5 ) , .A4( u1_u10_u7_n108 ) , .A3( u1_u10_u7_n109 ) , .A1( u1_u10_u7_n116 ) , .A2( u1_u10_u7_n123 ) );
  AOI22_X1 u1_u10_u7_U93 (.ZN( u1_u10_u7_n109 ) , .A2( u1_u10_u7_n126 ) , .B2( u1_u10_u7_n145 ) , .B1( u1_u10_u7_n156 ) , .A1( u1_u10_u7_n171 ) );
  NOR4_X1 u1_u10_u7_U94 (.A4( u1_u10_u7_n104 ) , .A3( u1_u10_u7_n105 ) , .A2( u1_u10_u7_n106 ) , .A1( u1_u10_u7_n107 ) , .ZN( u1_u10_u7_n108 ) );
  NAND3_X1 u1_u10_u7_U95 (.A3( u1_u10_u7_n146 ) , .A2( u1_u10_u7_n147 ) , .A1( u1_u10_u7_n148 ) , .ZN( u1_u10_u7_n151 ) );
  NAND3_X1 u1_u10_u7_U96 (.A3( u1_u10_u7_n131 ) , .A2( u1_u10_u7_n132 ) , .A1( u1_u10_u7_n133 ) , .ZN( u1_u10_u7_n135 ) );
  XOR2_X1 u1_u12_U2 (.B( u1_K13_8 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_8 ) );
  XOR2_X1 u1_u12_U27 (.B( u1_K13_2 ) , .A( u1_R11_1 ) , .Z( u1_u12_X_2 ) );
  XOR2_X1 u1_u12_U3 (.B( u1_K13_7 ) , .A( u1_R11_4 ) , .Z( u1_u12_X_7 ) );
  XOR2_X1 u1_u12_U37 (.B( u1_K13_20 ) , .A( u1_R11_13 ) , .Z( u1_u12_X_20 ) );
  XOR2_X1 u1_u12_U39 (.B( u1_K13_19 ) , .A( u1_R11_12 ) , .Z( u1_u12_X_19 ) );
  XOR2_X1 u1_u12_U4 (.B( u1_K13_6 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_6 ) );
  XOR2_X1 u1_u12_U40 (.B( u1_K13_18 ) , .A( u1_R11_13 ) , .Z( u1_u12_X_18 ) );
  XOR2_X1 u1_u12_U41 (.B( u1_K13_17 ) , .A( u1_R11_12 ) , .Z( u1_u12_X_17 ) );
  XOR2_X1 u1_u12_U43 (.B( u1_K13_15 ) , .A( u1_R11_10 ) , .Z( u1_u12_X_15 ) );
  XOR2_X1 u1_u12_U44 (.B( u1_K13_14 ) , .A( u1_R11_9 ) , .Z( u1_u12_X_14 ) );
  XOR2_X1 u1_u12_U45 (.B( u1_K13_13 ) , .A( u1_R11_8 ) , .Z( u1_u12_X_13 ) );
  XOR2_X1 u1_u12_U46 (.B( u1_K13_12 ) , .A( u1_R11_9 ) , .Z( u1_u12_X_12 ) );
  XOR2_X1 u1_u12_U47 (.B( u1_K13_11 ) , .A( u1_R11_8 ) , .Z( u1_u12_X_11 ) );
  XOR2_X1 u1_u12_U5 (.B( u1_K13_5 ) , .A( u1_R11_4 ) , .Z( u1_u12_X_5 ) );
  XOR2_X1 u1_u12_U7 (.B( u1_K13_48 ) , .A( u1_R11_1 ) , .Z( u1_u12_X_48 ) );
  NAND2_X1 u1_u12_u0_U10 (.ZN( u1_u12_u0_n113 ) , .A1( u1_u12_u0_n139 ) , .A2( u1_u12_u0_n149 ) );
  AND3_X1 u1_u12_u0_U11 (.A2( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n127 ) , .A3( u1_u12_u0_n130 ) , .A1( u1_u12_u0_n148 ) );
  AND2_X1 u1_u12_u0_U12 (.ZN( u1_u12_u0_n107 ) , .A1( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n140 ) );
  AND2_X1 u1_u12_u0_U13 (.A2( u1_u12_u0_n129 ) , .A1( u1_u12_u0_n130 ) , .ZN( u1_u12_u0_n151 ) );
  AND2_X1 u1_u12_u0_U14 (.A1( u1_u12_u0_n108 ) , .A2( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n145 ) );
  INV_X1 u1_u12_u0_U15 (.A( u1_u12_u0_n143 ) , .ZN( u1_u12_u0_n173 ) );
  NOR2_X1 u1_u12_u0_U16 (.A2( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n147 ) , .A1( u1_u12_u0_n160 ) );
  AOI21_X1 u1_u12_u0_U17 (.B1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n132 ) , .A( u1_u12_u0_n165 ) , .B2( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U18 (.A( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n165 ) );
  OAI22_X1 u1_u12_u0_U19 (.B1( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n147 ) , .A2( u1_u12_u0_n90 ) , .ZN( u1_u12_u0_n91 ) );
  AND3_X1 u1_u12_u0_U20 (.A3( u1_u12_u0_n121 ) , .A2( u1_u12_u0_n125 ) , .A1( u1_u12_u0_n148 ) , .ZN( u1_u12_u0_n90 ) );
  OAI22_X1 u1_u12_u0_U21 (.B1( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n126 ) , .A1( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n146 ) , .B2( u1_u12_u0_n147 ) );
  INV_X1 u1_u12_u0_U22 (.A( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n161 ) );
  AOI22_X1 u1_u12_u0_U23 (.B2( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n110 ) , .ZN( u1_u12_u0_n111 ) , .B1( u1_u12_u0_n118 ) , .A1( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U24 (.A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U25 (.A2( u1_u12_u0_n102 ) , .A1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n149 ) );
  INV_X1 u1_u12_u0_U26 (.A( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n158 ) );
  NAND2_X1 u1_u12_u0_U27 (.A2( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U28 (.ZN( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n92 ) , .A2( u1_u12_u0_n94 ) );
  AOI21_X1 u1_u12_u0_U29 (.ZN( u1_u12_u0_n104 ) , .B1( u1_u12_u0_n107 ) , .B2( u1_u12_u0_n141 ) , .A( u1_u12_u0_n144 ) );
  INV_X1 u1_u12_u0_U3 (.A( u1_u12_u0_n113 ) , .ZN( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U30 (.ZN( u1_u12_u0_n116 ) , .B2( u1_u12_u0_n142 ) , .A( u1_u12_u0_n144 ) , .B1( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U31 (.B1( u1_u12_u0_n127 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n96 ) );
  NAND2_X1 u1_u12_u0_U32 (.A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n114 ) , .A1( u1_u12_u0_n92 ) );
  NOR2_X1 u1_u12_u0_U33 (.A1( u1_u12_u0_n120 ) , .ZN( u1_u12_u0_n143 ) , .A2( u1_u12_u0_n167 ) );
  OAI221_X1 u1_u12_u0_U34 (.C1( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n120 ) , .B1( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n141 ) , .C2( u1_u12_u0_n147 ) , .A( u1_u12_u0_n172 ) );
  AOI211_X1 u1_u12_u0_U35 (.B( u1_u12_u0_n115 ) , .A( u1_u12_u0_n116 ) , .C2( u1_u12_u0_n117 ) , .C1( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n119 ) );
  NAND2_X1 u1_u12_u0_U36 (.A1( u1_u12_u0_n100 ) , .A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n125 ) );
  NAND2_X1 u1_u12_u0_U37 (.A1( u1_u12_u0_n101 ) , .A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n150 ) );
  INV_X1 u1_u12_u0_U38 (.A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U39 (.A2( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n139 ) );
  AOI21_X1 u1_u12_u0_U4 (.B1( u1_u12_u0_n114 ) , .ZN( u1_u12_u0_n115 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U40 (.A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U41 (.ZN( u1_u12_u0_n112 ) , .A2( u1_u12_u0_n92 ) , .A1( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U42 (.ZN( u1_u12_u0_n172 ) , .A( u1_u12_u0_n88 ) );
  OAI222_X1 u1_u12_u0_U43 (.C1( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n125 ) , .B2( u1_u12_u0_n128 ) , .B1( u1_u12_u0_n144 ) , .A2( u1_u12_u0_n158 ) , .C2( u1_u12_u0_n161 ) , .ZN( u1_u12_u0_n88 ) );
  NAND2_X1 u1_u12_u0_U44 (.A2( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n121 ) , .A1( u1_u12_u0_n93 ) );
  OR3_X1 u1_u12_u0_U45 (.A3( u1_u12_u0_n152 ) , .A2( u1_u12_u0_n153 ) , .A1( u1_u12_u0_n154 ) , .ZN( u1_u12_u0_n155 ) );
  AOI21_X1 u1_u12_u0_U46 (.B2( u1_u12_u0_n150 ) , .B1( u1_u12_u0_n151 ) , .ZN( u1_u12_u0_n152 ) , .A( u1_u12_u0_n158 ) );
  AOI21_X1 u1_u12_u0_U47 (.A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n145 ) , .B1( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n154 ) );
  AOI21_X1 u1_u12_u0_U48 (.A( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n148 ) , .B1( u1_u12_u0_n149 ) , .ZN( u1_u12_u0_n153 ) );
  INV_X1 u1_u12_u0_U49 (.ZN( u1_u12_u0_n171 ) , .A( u1_u12_u0_n99 ) );
  AOI21_X1 u1_u12_u0_U5 (.B2( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n134 ) , .B1( u1_u12_u0_n151 ) , .A( u1_u12_u0_n158 ) );
  OAI211_X1 u1_u12_u0_U50 (.C2( u1_u12_u0_n140 ) , .C1( u1_u12_u0_n161 ) , .A( u1_u12_u0_n169 ) , .B( u1_u12_u0_n98 ) , .ZN( u1_u12_u0_n99 ) );
  INV_X1 u1_u12_u0_U51 (.ZN( u1_u12_u0_n169 ) , .A( u1_u12_u0_n91 ) );
  AOI211_X1 u1_u12_u0_U52 (.C1( u1_u12_u0_n118 ) , .A( u1_u12_u0_n123 ) , .B( u1_u12_u0_n96 ) , .C2( u1_u12_u0_n97 ) , .ZN( u1_u12_u0_n98 ) );
  NOR2_X1 u1_u12_u0_U53 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n118 ) );
  NOR2_X1 u1_u12_u0_U54 (.A2( u1_u12_X_1 ) , .ZN( u1_u12_u0_n101 ) , .A1( u1_u12_u0_n163 ) );
  NOR2_X1 u1_u12_u0_U55 (.A2( u1_u12_X_6 ) , .ZN( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n162 ) );
  NAND2_X1 u1_u12_u0_U56 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n144 ) );
  NOR2_X1 u1_u12_u0_U57 (.A2( u1_u12_X_5 ) , .ZN( u1_u12_u0_n136 ) , .A1( u1_u12_u0_n159 ) );
  NAND2_X1 u1_u12_u0_U58 (.A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n159 ) );
  AND2_X1 u1_u12_u0_U59 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n102 ) );
  NOR2_X1 u1_u12_u0_U6 (.A1( u1_u12_u0_n108 ) , .ZN( u1_u12_u0_n123 ) , .A2( u1_u12_u0_n158 ) );
  AND2_X1 u1_u12_u0_U60 (.A1( u1_u12_X_6 ) , .A2( u1_u12_u0_n162 ) , .ZN( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U61 (.A( u1_u12_X_4 ) , .ZN( u1_u12_u0_n159 ) );
  INV_X1 u1_u12_u0_U62 (.A( u1_u12_X_1 ) , .ZN( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U63 (.A( u1_u12_X_3 ) , .ZN( u1_u12_u0_n162 ) );
  OR4_X1 u1_u12_u0_U64 (.ZN( u1_out12_17 ) , .A4( u1_u12_u0_n122 ) , .A2( u1_u12_u0_n123 ) , .A1( u1_u12_u0_n124 ) , .A3( u1_u12_u0_n170 ) );
  AOI21_X1 u1_u12_u0_U65 (.B2( u1_u12_u0_n107 ) , .ZN( u1_u12_u0_n124 ) , .B1( u1_u12_u0_n128 ) , .A( u1_u12_u0_n161 ) );
  INV_X1 u1_u12_u0_U66 (.A( u1_u12_u0_n111 ) , .ZN( u1_u12_u0_n170 ) );
  OR4_X1 u1_u12_u0_U67 (.ZN( u1_out12_31 ) , .A4( u1_u12_u0_n155 ) , .A2( u1_u12_u0_n156 ) , .A1( u1_u12_u0_n157 ) , .A3( u1_u12_u0_n173 ) );
  AOI21_X1 u1_u12_u0_U68 (.A( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n139 ) , .B1( u1_u12_u0_n140 ) , .ZN( u1_u12_u0_n157 ) );
  AOI21_X1 u1_u12_u0_U69 (.B2( u1_u12_u0_n141 ) , .B1( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n156 ) , .A( u1_u12_u0_n161 ) );
  OAI21_X1 u1_u12_u0_U7 (.B1( u1_u12_u0_n150 ) , .B2( u1_u12_u0_n158 ) , .A( u1_u12_u0_n172 ) , .ZN( u1_u12_u0_n89 ) );
  INV_X1 u1_u12_u0_U70 (.ZN( u1_u12_u0_n174 ) , .A( u1_u12_u0_n89 ) );
  AOI211_X1 u1_u12_u0_U71 (.B( u1_u12_u0_n104 ) , .A( u1_u12_u0_n105 ) , .ZN( u1_u12_u0_n106 ) , .C2( u1_u12_u0_n113 ) , .C1( u1_u12_u0_n160 ) );
  INV_X1 u1_u12_u0_U72 (.A( u1_u12_u0_n126 ) , .ZN( u1_u12_u0_n168 ) );
  AOI211_X1 u1_u12_u0_U73 (.B( u1_u12_u0_n133 ) , .A( u1_u12_u0_n134 ) , .C2( u1_u12_u0_n135 ) , .C1( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n137 ) );
  NOR2_X1 u1_u12_u0_U74 (.A1( u1_u12_u0_n163 ) , .A2( u1_u12_u0_n164 ) , .ZN( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U75 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n94 ) );
  OAI221_X1 u1_u12_u0_U76 (.C1( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n122 ) , .B2( u1_u12_u0_n127 ) , .A( u1_u12_u0_n143 ) , .B1( u1_u12_u0_n144 ) , .C2( u1_u12_u0_n147 ) );
  AOI21_X1 u1_u12_u0_U77 (.B1( u1_u12_u0_n132 ) , .ZN( u1_u12_u0_n133 ) , .A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n166 ) );
  OAI22_X1 u1_u12_u0_U78 (.ZN( u1_u12_u0_n105 ) , .A2( u1_u12_u0_n132 ) , .B1( u1_u12_u0_n146 ) , .A1( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U79 (.ZN( u1_u12_u0_n110 ) , .A2( u1_u12_u0_n132 ) , .A1( u1_u12_u0_n145 ) );
  AND2_X1 u1_u12_u0_U8 (.A1( u1_u12_u0_n114 ) , .A2( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n146 ) );
  INV_X1 u1_u12_u0_U80 (.A( u1_u12_u0_n119 ) , .ZN( u1_u12_u0_n167 ) );
  NAND2_X1 u1_u12_u0_U81 (.ZN( u1_u12_u0_n148 ) , .A1( u1_u12_u0_n93 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U82 (.A1( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n129 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U83 (.A1( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n128 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U84 (.A2( u1_u12_X_1 ) , .A1( u1_u12_X_2 ) , .ZN( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U85 (.ZN( u1_u12_u0_n142 ) , .A1( u1_u12_u0_n94 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U86 (.A2( u1_u12_X_2 ) , .ZN( u1_u12_u0_n103 ) , .A1( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U87 (.A( u1_u12_X_2 ) , .ZN( u1_u12_u0_n163 ) );
  NAND3_X1 u1_u12_u0_U88 (.ZN( u1_out12_23 ) , .A3( u1_u12_u0_n137 ) , .A1( u1_u12_u0_n168 ) , .A2( u1_u12_u0_n171 ) );
  NAND3_X1 u1_u12_u0_U89 (.A3( u1_u12_u0_n127 ) , .A2( u1_u12_u0_n128 ) , .ZN( u1_u12_u0_n135 ) , .A1( u1_u12_u0_n150 ) );
  AND2_X1 u1_u12_u0_U9 (.A1( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n141 ) , .A2( u1_u12_u0_n150 ) );
  NAND3_X1 u1_u12_u0_U90 (.ZN( u1_u12_u0_n117 ) , .A3( u1_u12_u0_n132 ) , .A2( u1_u12_u0_n139 ) , .A1( u1_u12_u0_n148 ) );
  NAND3_X1 u1_u12_u0_U91 (.ZN( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n114 ) , .A3( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n149 ) );
  NAND3_X1 u1_u12_u0_U92 (.ZN( u1_out12_9 ) , .A3( u1_u12_u0_n106 ) , .A2( u1_u12_u0_n171 ) , .A1( u1_u12_u0_n174 ) );
  NAND3_X1 u1_u12_u0_U93 (.A2( u1_u12_u0_n128 ) , .A1( u1_u12_u0_n132 ) , .A3( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n97 ) );
  NOR2_X1 u1_u12_u1_U10 (.A1( u1_u12_u1_n112 ) , .A2( u1_u12_u1_n116 ) , .ZN( u1_u12_u1_n118 ) );
  NAND3_X1 u1_u12_u1_U100 (.ZN( u1_u12_u1_n113 ) , .A1( u1_u12_u1_n120 ) , .A3( u1_u12_u1_n133 ) , .A2( u1_u12_u1_n155 ) );
  OAI21_X1 u1_u12_u1_U11 (.ZN( u1_u12_u1_n101 ) , .B1( u1_u12_u1_n141 ) , .A( u1_u12_u1_n146 ) , .B2( u1_u12_u1_n183 ) );
  AOI21_X1 u1_u12_u1_U12 (.B2( u1_u12_u1_n155 ) , .B1( u1_u12_u1_n156 ) , .ZN( u1_u12_u1_n157 ) , .A( u1_u12_u1_n174 ) );
  NAND2_X1 u1_u12_u1_U13 (.ZN( u1_u12_u1_n140 ) , .A2( u1_u12_u1_n150 ) , .A1( u1_u12_u1_n155 ) );
  NAND2_X1 u1_u12_u1_U14 (.A1( u1_u12_u1_n131 ) , .ZN( u1_u12_u1_n147 ) , .A2( u1_u12_u1_n153 ) );
  INV_X1 u1_u12_u1_U15 (.A( u1_u12_u1_n139 ) , .ZN( u1_u12_u1_n174 ) );
  OR4_X1 u1_u12_u1_U16 (.A4( u1_u12_u1_n106 ) , .A3( u1_u12_u1_n107 ) , .ZN( u1_u12_u1_n108 ) , .A1( u1_u12_u1_n117 ) , .A2( u1_u12_u1_n184 ) );
  AOI21_X1 u1_u12_u1_U17 (.ZN( u1_u12_u1_n106 ) , .A( u1_u12_u1_n112 ) , .B1( u1_u12_u1_n154 ) , .B2( u1_u12_u1_n156 ) );
  INV_X1 u1_u12_u1_U18 (.A( u1_u12_u1_n101 ) , .ZN( u1_u12_u1_n184 ) );
  AOI21_X1 u1_u12_u1_U19 (.ZN( u1_u12_u1_n107 ) , .B1( u1_u12_u1_n134 ) , .B2( u1_u12_u1_n149 ) , .A( u1_u12_u1_n174 ) );
  INV_X1 u1_u12_u1_U20 (.A( u1_u12_u1_n112 ) , .ZN( u1_u12_u1_n171 ) );
  NAND2_X1 u1_u12_u1_U21 (.ZN( u1_u12_u1_n141 ) , .A1( u1_u12_u1_n153 ) , .A2( u1_u12_u1_n156 ) );
  AND2_X1 u1_u12_u1_U22 (.A1( u1_u12_u1_n123 ) , .ZN( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n161 ) );
  NAND2_X1 u1_u12_u1_U23 (.A2( u1_u12_u1_n115 ) , .A1( u1_u12_u1_n116 ) , .ZN( u1_u12_u1_n148 ) );
  NAND2_X1 u1_u12_u1_U24 (.A2( u1_u12_u1_n133 ) , .A1( u1_u12_u1_n135 ) , .ZN( u1_u12_u1_n159 ) );
  NAND2_X1 u1_u12_u1_U25 (.A2( u1_u12_u1_n115 ) , .A1( u1_u12_u1_n120 ) , .ZN( u1_u12_u1_n132 ) );
  INV_X1 u1_u12_u1_U26 (.A( u1_u12_u1_n154 ) , .ZN( u1_u12_u1_n178 ) );
  INV_X1 u1_u12_u1_U27 (.A( u1_u12_u1_n151 ) , .ZN( u1_u12_u1_n183 ) );
  AND2_X1 u1_u12_u1_U28 (.A1( u1_u12_u1_n129 ) , .A2( u1_u12_u1_n133 ) , .ZN( u1_u12_u1_n149 ) );
  INV_X1 u1_u12_u1_U29 (.A( u1_u12_u1_n131 ) , .ZN( u1_u12_u1_n180 ) );
  INV_X1 u1_u12_u1_U3 (.A( u1_u12_u1_n159 ) , .ZN( u1_u12_u1_n182 ) );
  AOI221_X1 u1_u12_u1_U30 (.B1( u1_u12_u1_n140 ) , .ZN( u1_u12_u1_n167 ) , .B2( u1_u12_u1_n172 ) , .C2( u1_u12_u1_n175 ) , .C1( u1_u12_u1_n178 ) , .A( u1_u12_u1_n188 ) );
  INV_X1 u1_u12_u1_U31 (.ZN( u1_u12_u1_n188 ) , .A( u1_u12_u1_n97 ) );
  AOI211_X1 u1_u12_u1_U32 (.A( u1_u12_u1_n118 ) , .C1( u1_u12_u1_n132 ) , .C2( u1_u12_u1_n139 ) , .B( u1_u12_u1_n96 ) , .ZN( u1_u12_u1_n97 ) );
  AOI21_X1 u1_u12_u1_U33 (.B2( u1_u12_u1_n121 ) , .B1( u1_u12_u1_n135 ) , .A( u1_u12_u1_n152 ) , .ZN( u1_u12_u1_n96 ) );
  OAI221_X1 u1_u12_u1_U34 (.A( u1_u12_u1_n119 ) , .C2( u1_u12_u1_n129 ) , .ZN( u1_u12_u1_n138 ) , .B2( u1_u12_u1_n152 ) , .C1( u1_u12_u1_n174 ) , .B1( u1_u12_u1_n187 ) );
  INV_X1 u1_u12_u1_U35 (.A( u1_u12_u1_n148 ) , .ZN( u1_u12_u1_n187 ) );
  AOI211_X1 u1_u12_u1_U36 (.B( u1_u12_u1_n117 ) , .A( u1_u12_u1_n118 ) , .ZN( u1_u12_u1_n119 ) , .C2( u1_u12_u1_n146 ) , .C1( u1_u12_u1_n159 ) );
  NOR2_X1 u1_u12_u1_U37 (.A1( u1_u12_u1_n168 ) , .A2( u1_u12_u1_n176 ) , .ZN( u1_u12_u1_n98 ) );
  AOI211_X1 u1_u12_u1_U38 (.B( u1_u12_u1_n162 ) , .A( u1_u12_u1_n163 ) , .C2( u1_u12_u1_n164 ) , .ZN( u1_u12_u1_n165 ) , .C1( u1_u12_u1_n171 ) );
  AOI21_X1 u1_u12_u1_U39 (.A( u1_u12_u1_n160 ) , .B2( u1_u12_u1_n161 ) , .ZN( u1_u12_u1_n162 ) , .B1( u1_u12_u1_n182 ) );
  AOI221_X1 u1_u12_u1_U4 (.A( u1_u12_u1_n138 ) , .C2( u1_u12_u1_n139 ) , .C1( u1_u12_u1_n140 ) , .B2( u1_u12_u1_n141 ) , .ZN( u1_u12_u1_n142 ) , .B1( u1_u12_u1_n175 ) );
  OR2_X1 u1_u12_u1_U40 (.A2( u1_u12_u1_n157 ) , .A1( u1_u12_u1_n158 ) , .ZN( u1_u12_u1_n163 ) );
  NAND2_X1 u1_u12_u1_U41 (.A1( u1_u12_u1_n128 ) , .ZN( u1_u12_u1_n146 ) , .A2( u1_u12_u1_n160 ) );
  NAND2_X1 u1_u12_u1_U42 (.A2( u1_u12_u1_n112 ) , .ZN( u1_u12_u1_n139 ) , .A1( u1_u12_u1_n152 ) );
  NAND2_X1 u1_u12_u1_U43 (.A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n156 ) , .A2( u1_u12_u1_n99 ) );
  NOR2_X1 u1_u12_u1_U44 (.ZN( u1_u12_u1_n117 ) , .A1( u1_u12_u1_n121 ) , .A2( u1_u12_u1_n160 ) );
  OAI21_X1 u1_u12_u1_U45 (.B2( u1_u12_u1_n123 ) , .ZN( u1_u12_u1_n145 ) , .B1( u1_u12_u1_n160 ) , .A( u1_u12_u1_n185 ) );
  INV_X1 u1_u12_u1_U46 (.A( u1_u12_u1_n122 ) , .ZN( u1_u12_u1_n185 ) );
  AOI21_X1 u1_u12_u1_U47 (.B2( u1_u12_u1_n120 ) , .B1( u1_u12_u1_n121 ) , .ZN( u1_u12_u1_n122 ) , .A( u1_u12_u1_n128 ) );
  AOI21_X1 u1_u12_u1_U48 (.A( u1_u12_u1_n128 ) , .B2( u1_u12_u1_n129 ) , .ZN( u1_u12_u1_n130 ) , .B1( u1_u12_u1_n150 ) );
  NAND2_X1 u1_u12_u1_U49 (.ZN( u1_u12_u1_n112 ) , .A1( u1_u12_u1_n169 ) , .A2( u1_u12_u1_n170 ) );
  AOI211_X1 u1_u12_u1_U5 (.ZN( u1_u12_u1_n124 ) , .A( u1_u12_u1_n138 ) , .C2( u1_u12_u1_n139 ) , .B( u1_u12_u1_n145 ) , .C1( u1_u12_u1_n147 ) );
  NAND2_X1 u1_u12_u1_U50 (.ZN( u1_u12_u1_n129 ) , .A2( u1_u12_u1_n95 ) , .A1( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U51 (.A1( u1_u12_u1_n102 ) , .ZN( u1_u12_u1_n154 ) , .A2( u1_u12_u1_n99 ) );
  NAND2_X1 u1_u12_u1_U52 (.A2( u1_u12_u1_n100 ) , .ZN( u1_u12_u1_n135 ) , .A1( u1_u12_u1_n99 ) );
  AOI21_X1 u1_u12_u1_U53 (.A( u1_u12_u1_n152 ) , .B2( u1_u12_u1_n153 ) , .B1( u1_u12_u1_n154 ) , .ZN( u1_u12_u1_n158 ) );
  INV_X1 u1_u12_u1_U54 (.A( u1_u12_u1_n160 ) , .ZN( u1_u12_u1_n175 ) );
  NAND2_X1 u1_u12_u1_U55 (.A1( u1_u12_u1_n100 ) , .ZN( u1_u12_u1_n116 ) , .A2( u1_u12_u1_n95 ) );
  NAND2_X1 u1_u12_u1_U56 (.A1( u1_u12_u1_n102 ) , .ZN( u1_u12_u1_n131 ) , .A2( u1_u12_u1_n95 ) );
  NAND2_X1 u1_u12_u1_U57 (.A2( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n121 ) , .A1( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U58 (.A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n153 ) , .A2( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U59 (.A2( u1_u12_u1_n104 ) , .A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n133 ) );
  AOI22_X1 u1_u12_u1_U6 (.B2( u1_u12_u1_n113 ) , .A2( u1_u12_u1_n114 ) , .ZN( u1_u12_u1_n125 ) , .A1( u1_u12_u1_n171 ) , .B1( u1_u12_u1_n173 ) );
  NAND2_X1 u1_u12_u1_U60 (.ZN( u1_u12_u1_n150 ) , .A2( u1_u12_u1_n98 ) , .A1( u1_u12_u1_n99 ) );
  NAND2_X1 u1_u12_u1_U61 (.A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n155 ) , .A2( u1_u12_u1_n95 ) );
  OAI21_X1 u1_u12_u1_U62 (.ZN( u1_u12_u1_n109 ) , .B1( u1_u12_u1_n129 ) , .B2( u1_u12_u1_n160 ) , .A( u1_u12_u1_n167 ) );
  NAND2_X1 u1_u12_u1_U63 (.A2( u1_u12_u1_n100 ) , .A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n120 ) );
  NAND2_X1 u1_u12_u1_U64 (.A1( u1_u12_u1_n102 ) , .A2( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n115 ) );
  NAND2_X1 u1_u12_u1_U65 (.A2( u1_u12_u1_n100 ) , .A1( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n151 ) );
  NAND2_X1 u1_u12_u1_U66 (.A2( u1_u12_u1_n103 ) , .A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n161 ) );
  INV_X1 u1_u12_u1_U67 (.A( u1_u12_u1_n152 ) , .ZN( u1_u12_u1_n173 ) );
  INV_X1 u1_u12_u1_U68 (.A( u1_u12_u1_n128 ) , .ZN( u1_u12_u1_n172 ) );
  NAND2_X1 u1_u12_u1_U69 (.A2( u1_u12_u1_n102 ) , .A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n123 ) );
  NAND2_X1 u1_u12_u1_U7 (.ZN( u1_u12_u1_n114 ) , .A1( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n156 ) );
  NOR2_X1 u1_u12_u1_U70 (.A2( u1_u12_X_7 ) , .A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n95 ) );
  NOR2_X1 u1_u12_u1_U71 (.A1( u1_u12_X_12 ) , .A2( u1_u12_X_9 ) , .ZN( u1_u12_u1_n100 ) );
  NOR2_X1 u1_u12_u1_U72 (.A2( u1_u12_X_8 ) , .A1( u1_u12_u1_n177 ) , .ZN( u1_u12_u1_n99 ) );
  NOR2_X1 u1_u12_u1_U73 (.A2( u1_u12_X_12 ) , .ZN( u1_u12_u1_n102 ) , .A1( u1_u12_u1_n176 ) );
  NOR2_X1 u1_u12_u1_U74 (.A2( u1_u12_X_9 ) , .ZN( u1_u12_u1_n105 ) , .A1( u1_u12_u1_n168 ) );
  NAND2_X1 u1_u12_u1_U75 (.A1( u1_u12_X_10 ) , .ZN( u1_u12_u1_n160 ) , .A2( u1_u12_u1_n169 ) );
  NAND2_X1 u1_u12_u1_U76 (.A2( u1_u12_X_10 ) , .A1( u1_u12_X_11 ) , .ZN( u1_u12_u1_n152 ) );
  NAND2_X1 u1_u12_u1_U77 (.A1( u1_u12_X_11 ) , .ZN( u1_u12_u1_n128 ) , .A2( u1_u12_u1_n170 ) );
  AND2_X1 u1_u12_u1_U78 (.A2( u1_u12_X_7 ) , .A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n104 ) );
  AND2_X1 u1_u12_u1_U79 (.A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n103 ) , .A2( u1_u12_u1_n177 ) );
  AOI22_X1 u1_u12_u1_U8 (.B2( u1_u12_u1_n136 ) , .A2( u1_u12_u1_n137 ) , .ZN( u1_u12_u1_n143 ) , .A1( u1_u12_u1_n171 ) , .B1( u1_u12_u1_n173 ) );
  INV_X1 u1_u12_u1_U80 (.A( u1_u12_X_10 ) , .ZN( u1_u12_u1_n170 ) );
  INV_X1 u1_u12_u1_U81 (.A( u1_u12_X_9 ) , .ZN( u1_u12_u1_n176 ) );
  INV_X1 u1_u12_u1_U82 (.A( u1_u12_X_11 ) , .ZN( u1_u12_u1_n169 ) );
  INV_X1 u1_u12_u1_U83 (.A( u1_u12_X_12 ) , .ZN( u1_u12_u1_n168 ) );
  INV_X1 u1_u12_u1_U84 (.A( u1_u12_X_7 ) , .ZN( u1_u12_u1_n177 ) );
  NAND4_X1 u1_u12_u1_U85 (.ZN( u1_out12_28 ) , .A4( u1_u12_u1_n124 ) , .A3( u1_u12_u1_n125 ) , .A2( u1_u12_u1_n126 ) , .A1( u1_u12_u1_n127 ) );
  OAI21_X1 u1_u12_u1_U86 (.ZN( u1_u12_u1_n127 ) , .B2( u1_u12_u1_n139 ) , .B1( u1_u12_u1_n175 ) , .A( u1_u12_u1_n183 ) );
  OAI21_X1 u1_u12_u1_U87 (.ZN( u1_u12_u1_n126 ) , .B2( u1_u12_u1_n140 ) , .A( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n178 ) );
  NAND4_X1 u1_u12_u1_U88 (.ZN( u1_out12_18 ) , .A4( u1_u12_u1_n165 ) , .A3( u1_u12_u1_n166 ) , .A1( u1_u12_u1_n167 ) , .A2( u1_u12_u1_n186 ) );
  AOI22_X1 u1_u12_u1_U89 (.B2( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n147 ) , .A2( u1_u12_u1_n148 ) , .ZN( u1_u12_u1_n166 ) , .A1( u1_u12_u1_n172 ) );
  INV_X1 u1_u12_u1_U9 (.A( u1_u12_u1_n147 ) , .ZN( u1_u12_u1_n181 ) );
  INV_X1 u1_u12_u1_U90 (.A( u1_u12_u1_n145 ) , .ZN( u1_u12_u1_n186 ) );
  NAND4_X1 u1_u12_u1_U91 (.ZN( u1_out12_2 ) , .A4( u1_u12_u1_n142 ) , .A3( u1_u12_u1_n143 ) , .A2( u1_u12_u1_n144 ) , .A1( u1_u12_u1_n179 ) );
  OAI21_X1 u1_u12_u1_U92 (.B2( u1_u12_u1_n132 ) , .ZN( u1_u12_u1_n144 ) , .A( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n180 ) );
  INV_X1 u1_u12_u1_U93 (.A( u1_u12_u1_n130 ) , .ZN( u1_u12_u1_n179 ) );
  OR4_X1 u1_u12_u1_U94 (.ZN( u1_out12_13 ) , .A4( u1_u12_u1_n108 ) , .A3( u1_u12_u1_n109 ) , .A2( u1_u12_u1_n110 ) , .A1( u1_u12_u1_n111 ) );
  AOI21_X1 u1_u12_u1_U95 (.ZN( u1_u12_u1_n111 ) , .A( u1_u12_u1_n128 ) , .B2( u1_u12_u1_n131 ) , .B1( u1_u12_u1_n135 ) );
  AOI21_X1 u1_u12_u1_U96 (.ZN( u1_u12_u1_n110 ) , .A( u1_u12_u1_n116 ) , .B1( u1_u12_u1_n152 ) , .B2( u1_u12_u1_n160 ) );
  NAND3_X1 u1_u12_u1_U97 (.A3( u1_u12_u1_n149 ) , .A2( u1_u12_u1_n150 ) , .A1( u1_u12_u1_n151 ) , .ZN( u1_u12_u1_n164 ) );
  NAND3_X1 u1_u12_u1_U98 (.A3( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n135 ) , .ZN( u1_u12_u1_n136 ) , .A1( u1_u12_u1_n151 ) );
  NAND3_X1 u1_u12_u1_U99 (.A1( u1_u12_u1_n133 ) , .ZN( u1_u12_u1_n137 ) , .A2( u1_u12_u1_n154 ) , .A3( u1_u12_u1_n181 ) );
  OAI22_X1 u1_u12_u2_U10 (.B1( u1_u12_u2_n151 ) , .A2( u1_u12_u2_n152 ) , .A1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n160 ) , .B2( u1_u12_u2_n168 ) );
  NAND3_X1 u1_u12_u2_U100 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n98 ) );
  NOR3_X1 u1_u12_u2_U11 (.A1( u1_u12_u2_n150 ) , .ZN( u1_u12_u2_n151 ) , .A3( u1_u12_u2_n175 ) , .A2( u1_u12_u2_n188 ) );
  AOI21_X1 u1_u12_u2_U12 (.B2( u1_u12_u2_n123 ) , .ZN( u1_u12_u2_n125 ) , .A( u1_u12_u2_n171 ) , .B1( u1_u12_u2_n184 ) );
  INV_X1 u1_u12_u2_U13 (.A( u1_u12_u2_n150 ) , .ZN( u1_u12_u2_n184 ) );
  AOI21_X1 u1_u12_u2_U14 (.ZN( u1_u12_u2_n144 ) , .B2( u1_u12_u2_n155 ) , .A( u1_u12_u2_n172 ) , .B1( u1_u12_u2_n185 ) );
  AOI21_X1 u1_u12_u2_U15 (.B2( u1_u12_u2_n143 ) , .ZN( u1_u12_u2_n145 ) , .B1( u1_u12_u2_n152 ) , .A( u1_u12_u2_n171 ) );
  INV_X1 u1_u12_u2_U16 (.A( u1_u12_u2_n156 ) , .ZN( u1_u12_u2_n171 ) );
  INV_X1 u1_u12_u2_U17 (.A( u1_u12_u2_n120 ) , .ZN( u1_u12_u2_n188 ) );
  NAND2_X1 u1_u12_u2_U18 (.A2( u1_u12_u2_n122 ) , .ZN( u1_u12_u2_n150 ) , .A1( u1_u12_u2_n152 ) );
  INV_X1 u1_u12_u2_U19 (.A( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n170 ) );
  INV_X1 u1_u12_u2_U20 (.A( u1_u12_u2_n137 ) , .ZN( u1_u12_u2_n173 ) );
  NAND2_X1 u1_u12_u2_U21 (.A1( u1_u12_u2_n132 ) , .A2( u1_u12_u2_n139 ) , .ZN( u1_u12_u2_n157 ) );
  INV_X1 u1_u12_u2_U22 (.A( u1_u12_u2_n113 ) , .ZN( u1_u12_u2_n178 ) );
  INV_X1 u1_u12_u2_U23 (.A( u1_u12_u2_n139 ) , .ZN( u1_u12_u2_n175 ) );
  INV_X1 u1_u12_u2_U24 (.A( u1_u12_u2_n155 ) , .ZN( u1_u12_u2_n181 ) );
  INV_X1 u1_u12_u2_U25 (.A( u1_u12_u2_n119 ) , .ZN( u1_u12_u2_n177 ) );
  INV_X1 u1_u12_u2_U26 (.A( u1_u12_u2_n116 ) , .ZN( u1_u12_u2_n180 ) );
  INV_X1 u1_u12_u2_U27 (.A( u1_u12_u2_n131 ) , .ZN( u1_u12_u2_n179 ) );
  INV_X1 u1_u12_u2_U28 (.A( u1_u12_u2_n154 ) , .ZN( u1_u12_u2_n176 ) );
  NAND2_X1 u1_u12_u2_U29 (.A2( u1_u12_u2_n116 ) , .A1( u1_u12_u2_n117 ) , .ZN( u1_u12_u2_n118 ) );
  NOR2_X1 u1_u12_u2_U3 (.ZN( u1_u12_u2_n121 ) , .A2( u1_u12_u2_n177 ) , .A1( u1_u12_u2_n180 ) );
  INV_X1 u1_u12_u2_U30 (.A( u1_u12_u2_n132 ) , .ZN( u1_u12_u2_n182 ) );
  INV_X1 u1_u12_u2_U31 (.A( u1_u12_u2_n158 ) , .ZN( u1_u12_u2_n183 ) );
  OAI21_X1 u1_u12_u2_U32 (.A( u1_u12_u2_n156 ) , .B1( u1_u12_u2_n157 ) , .ZN( u1_u12_u2_n158 ) , .B2( u1_u12_u2_n179 ) );
  NOR2_X1 u1_u12_u2_U33 (.ZN( u1_u12_u2_n156 ) , .A1( u1_u12_u2_n166 ) , .A2( u1_u12_u2_n169 ) );
  NOR2_X1 u1_u12_u2_U34 (.A2( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n137 ) , .A1( u1_u12_u2_n140 ) );
  NOR2_X1 u1_u12_u2_U35 (.A2( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n153 ) , .A1( u1_u12_u2_n156 ) );
  AOI211_X1 u1_u12_u2_U36 (.ZN( u1_u12_u2_n130 ) , .C1( u1_u12_u2_n138 ) , .C2( u1_u12_u2_n179 ) , .B( u1_u12_u2_n96 ) , .A( u1_u12_u2_n97 ) );
  OAI22_X1 u1_u12_u2_U37 (.B1( u1_u12_u2_n133 ) , .A2( u1_u12_u2_n137 ) , .A1( u1_u12_u2_n152 ) , .B2( u1_u12_u2_n168 ) , .ZN( u1_u12_u2_n97 ) );
  OAI221_X1 u1_u12_u2_U38 (.B1( u1_u12_u2_n113 ) , .C1( u1_u12_u2_n132 ) , .A( u1_u12_u2_n149 ) , .B2( u1_u12_u2_n171 ) , .C2( u1_u12_u2_n172 ) , .ZN( u1_u12_u2_n96 ) );
  OAI221_X1 u1_u12_u2_U39 (.A( u1_u12_u2_n115 ) , .C2( u1_u12_u2_n123 ) , .B2( u1_u12_u2_n143 ) , .B1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n163 ) , .C1( u1_u12_u2_n168 ) );
  INV_X1 u1_u12_u2_U4 (.A( u1_u12_u2_n134 ) , .ZN( u1_u12_u2_n185 ) );
  OAI21_X1 u1_u12_u2_U40 (.A( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n115 ) , .B1( u1_u12_u2_n176 ) , .B2( u1_u12_u2_n178 ) );
  OAI221_X1 u1_u12_u2_U41 (.A( u1_u12_u2_n135 ) , .B2( u1_u12_u2_n136 ) , .B1( u1_u12_u2_n137 ) , .ZN( u1_u12_u2_n162 ) , .C2( u1_u12_u2_n167 ) , .C1( u1_u12_u2_n185 ) );
  AND3_X1 u1_u12_u2_U42 (.A3( u1_u12_u2_n131 ) , .A2( u1_u12_u2_n132 ) , .A1( u1_u12_u2_n133 ) , .ZN( u1_u12_u2_n136 ) );
  AOI22_X1 u1_u12_u2_U43 (.ZN( u1_u12_u2_n135 ) , .B1( u1_u12_u2_n140 ) , .A1( u1_u12_u2_n156 ) , .B2( u1_u12_u2_n180 ) , .A2( u1_u12_u2_n188 ) );
  AOI21_X1 u1_u12_u2_U44 (.ZN( u1_u12_u2_n149 ) , .B1( u1_u12_u2_n173 ) , .B2( u1_u12_u2_n188 ) , .A( u1_u12_u2_n95 ) );
  AND3_X1 u1_u12_u2_U45 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n156 ) , .ZN( u1_u12_u2_n95 ) );
  OAI21_X1 u1_u12_u2_U46 (.A( u1_u12_u2_n101 ) , .B2( u1_u12_u2_n121 ) , .B1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n164 ) );
  NAND2_X1 u1_u12_u2_U47 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n155 ) );
  NAND2_X1 u1_u12_u2_U48 (.A2( u1_u12_u2_n105 ) , .A1( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n143 ) );
  NAND2_X1 u1_u12_u2_U49 (.A1( u1_u12_u2_n104 ) , .A2( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n152 ) );
  NOR4_X1 u1_u12_u2_U5 (.A4( u1_u12_u2_n124 ) , .A3( u1_u12_u2_n125 ) , .A2( u1_u12_u2_n126 ) , .A1( u1_u12_u2_n127 ) , .ZN( u1_u12_u2_n128 ) );
  NAND2_X1 u1_u12_u2_U50 (.A1( u1_u12_u2_n100 ) , .A2( u1_u12_u2_n105 ) , .ZN( u1_u12_u2_n132 ) );
  INV_X1 u1_u12_u2_U51 (.A( u1_u12_u2_n140 ) , .ZN( u1_u12_u2_n168 ) );
  INV_X1 u1_u12_u2_U52 (.A( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n167 ) );
  OAI21_X1 u1_u12_u2_U53 (.A( u1_u12_u2_n141 ) , .B2( u1_u12_u2_n142 ) , .ZN( u1_u12_u2_n146 ) , .B1( u1_u12_u2_n153 ) );
  OAI21_X1 u1_u12_u2_U54 (.A( u1_u12_u2_n140 ) , .ZN( u1_u12_u2_n141 ) , .B1( u1_u12_u2_n176 ) , .B2( u1_u12_u2_n177 ) );
  NOR3_X1 u1_u12_u2_U55 (.ZN( u1_u12_u2_n142 ) , .A3( u1_u12_u2_n175 ) , .A2( u1_u12_u2_n178 ) , .A1( u1_u12_u2_n181 ) );
  NAND2_X1 u1_u12_u2_U56 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n113 ) );
  NAND2_X1 u1_u12_u2_U57 (.A1( u1_u12_u2_n106 ) , .A2( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n131 ) );
  NAND2_X1 u1_u12_u2_U58 (.A1( u1_u12_u2_n103 ) , .A2( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n139 ) );
  NAND2_X1 u1_u12_u2_U59 (.A1( u1_u12_u2_n103 ) , .A2( u1_u12_u2_n105 ) , .ZN( u1_u12_u2_n133 ) );
  AOI21_X1 u1_u12_u2_U6 (.B2( u1_u12_u2_n119 ) , .ZN( u1_u12_u2_n127 ) , .A( u1_u12_u2_n137 ) , .B1( u1_u12_u2_n155 ) );
  NAND2_X1 u1_u12_u2_U60 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n103 ) , .ZN( u1_u12_u2_n154 ) );
  NAND2_X1 u1_u12_u2_U61 (.A2( u1_u12_u2_n103 ) , .A1( u1_u12_u2_n104 ) , .ZN( u1_u12_u2_n119 ) );
  NAND2_X1 u1_u12_u2_U62 (.A2( u1_u12_u2_n107 ) , .A1( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n123 ) );
  NAND2_X1 u1_u12_u2_U63 (.A1( u1_u12_u2_n104 ) , .A2( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n122 ) );
  INV_X1 u1_u12_u2_U64 (.A( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n172 ) );
  NAND2_X1 u1_u12_u2_U65 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n102 ) , .ZN( u1_u12_u2_n116 ) );
  NAND2_X1 u1_u12_u2_U66 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n120 ) );
  NAND2_X1 u1_u12_u2_U67 (.A2( u1_u12_u2_n105 ) , .A1( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n117 ) );
  INV_X1 u1_u12_u2_U68 (.ZN( u1_u12_u2_n187 ) , .A( u1_u12_u2_n99 ) );
  OAI21_X1 u1_u12_u2_U69 (.B1( u1_u12_u2_n137 ) , .B2( u1_u12_u2_n143 ) , .A( u1_u12_u2_n98 ) , .ZN( u1_u12_u2_n99 ) );
  AOI21_X1 u1_u12_u2_U7 (.ZN( u1_u12_u2_n124 ) , .B1( u1_u12_u2_n131 ) , .B2( u1_u12_u2_n143 ) , .A( u1_u12_u2_n172 ) );
  NOR2_X1 u1_u12_u2_U70 (.A2( u1_u12_X_16 ) , .ZN( u1_u12_u2_n140 ) , .A1( u1_u12_u2_n166 ) );
  NOR2_X1 u1_u12_u2_U71 (.A2( u1_u12_X_13 ) , .A1( u1_u12_X_14 ) , .ZN( u1_u12_u2_n100 ) );
  NOR2_X1 u1_u12_u2_U72 (.A2( u1_u12_X_16 ) , .A1( u1_u12_X_17 ) , .ZN( u1_u12_u2_n138 ) );
  NOR2_X1 u1_u12_u2_U73 (.A2( u1_u12_X_15 ) , .A1( u1_u12_X_18 ) , .ZN( u1_u12_u2_n104 ) );
  NOR2_X1 u1_u12_u2_U74 (.A2( u1_u12_X_14 ) , .ZN( u1_u12_u2_n103 ) , .A1( u1_u12_u2_n174 ) );
  NOR2_X1 u1_u12_u2_U75 (.A2( u1_u12_X_15 ) , .ZN( u1_u12_u2_n102 ) , .A1( u1_u12_u2_n165 ) );
  NOR2_X1 u1_u12_u2_U76 (.A2( u1_u12_X_17 ) , .ZN( u1_u12_u2_n114 ) , .A1( u1_u12_u2_n169 ) );
  AND2_X1 u1_u12_u2_U77 (.A1( u1_u12_X_15 ) , .ZN( u1_u12_u2_n105 ) , .A2( u1_u12_u2_n165 ) );
  AND2_X1 u1_u12_u2_U78 (.A2( u1_u12_X_15 ) , .A1( u1_u12_X_18 ) , .ZN( u1_u12_u2_n107 ) );
  AND2_X1 u1_u12_u2_U79 (.A1( u1_u12_X_14 ) , .ZN( u1_u12_u2_n106 ) , .A2( u1_u12_u2_n174 ) );
  AOI21_X1 u1_u12_u2_U8 (.B2( u1_u12_u2_n120 ) , .B1( u1_u12_u2_n121 ) , .ZN( u1_u12_u2_n126 ) , .A( u1_u12_u2_n167 ) );
  AND2_X1 u1_u12_u2_U80 (.A1( u1_u12_X_13 ) , .A2( u1_u12_X_14 ) , .ZN( u1_u12_u2_n108 ) );
  INV_X1 u1_u12_u2_U81 (.A( u1_u12_X_16 ) , .ZN( u1_u12_u2_n169 ) );
  INV_X1 u1_u12_u2_U82 (.A( u1_u12_X_17 ) , .ZN( u1_u12_u2_n166 ) );
  INV_X1 u1_u12_u2_U83 (.A( u1_u12_X_13 ) , .ZN( u1_u12_u2_n174 ) );
  INV_X1 u1_u12_u2_U84 (.A( u1_u12_X_18 ) , .ZN( u1_u12_u2_n165 ) );
  NAND4_X1 u1_u12_u2_U85 (.ZN( u1_out12_30 ) , .A4( u1_u12_u2_n147 ) , .A3( u1_u12_u2_n148 ) , .A2( u1_u12_u2_n149 ) , .A1( u1_u12_u2_n187 ) );
  AOI21_X1 u1_u12_u2_U86 (.B2( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n148 ) , .A( u1_u12_u2_n162 ) , .B1( u1_u12_u2_n182 ) );
  NOR3_X1 u1_u12_u2_U87 (.A3( u1_u12_u2_n144 ) , .A2( u1_u12_u2_n145 ) , .A1( u1_u12_u2_n146 ) , .ZN( u1_u12_u2_n147 ) );
  NAND4_X1 u1_u12_u2_U88 (.ZN( u1_out12_24 ) , .A4( u1_u12_u2_n111 ) , .A3( u1_u12_u2_n112 ) , .A1( u1_u12_u2_n130 ) , .A2( u1_u12_u2_n187 ) );
  AOI221_X1 u1_u12_u2_U89 (.A( u1_u12_u2_n109 ) , .B1( u1_u12_u2_n110 ) , .ZN( u1_u12_u2_n111 ) , .C1( u1_u12_u2_n134 ) , .C2( u1_u12_u2_n170 ) , .B2( u1_u12_u2_n173 ) );
  OAI22_X1 u1_u12_u2_U9 (.ZN( u1_u12_u2_n109 ) , .A2( u1_u12_u2_n113 ) , .B2( u1_u12_u2_n133 ) , .B1( u1_u12_u2_n167 ) , .A1( u1_u12_u2_n168 ) );
  AOI21_X1 u1_u12_u2_U90 (.ZN( u1_u12_u2_n112 ) , .B2( u1_u12_u2_n156 ) , .A( u1_u12_u2_n164 ) , .B1( u1_u12_u2_n181 ) );
  NAND4_X1 u1_u12_u2_U91 (.ZN( u1_out12_16 ) , .A4( u1_u12_u2_n128 ) , .A3( u1_u12_u2_n129 ) , .A1( u1_u12_u2_n130 ) , .A2( u1_u12_u2_n186 ) );
  AOI22_X1 u1_u12_u2_U92 (.A2( u1_u12_u2_n118 ) , .ZN( u1_u12_u2_n129 ) , .A1( u1_u12_u2_n140 ) , .B1( u1_u12_u2_n157 ) , .B2( u1_u12_u2_n170 ) );
  INV_X1 u1_u12_u2_U93 (.A( u1_u12_u2_n163 ) , .ZN( u1_u12_u2_n186 ) );
  OR4_X1 u1_u12_u2_U94 (.ZN( u1_out12_6 ) , .A4( u1_u12_u2_n161 ) , .A3( u1_u12_u2_n162 ) , .A2( u1_u12_u2_n163 ) , .A1( u1_u12_u2_n164 ) );
  OR3_X1 u1_u12_u2_U95 (.A2( u1_u12_u2_n159 ) , .A1( u1_u12_u2_n160 ) , .ZN( u1_u12_u2_n161 ) , .A3( u1_u12_u2_n183 ) );
  AOI21_X1 u1_u12_u2_U96 (.B2( u1_u12_u2_n154 ) , .B1( u1_u12_u2_n155 ) , .ZN( u1_u12_u2_n159 ) , .A( u1_u12_u2_n167 ) );
  NAND3_X1 u1_u12_u2_U97 (.A2( u1_u12_u2_n117 ) , .A1( u1_u12_u2_n122 ) , .A3( u1_u12_u2_n123 ) , .ZN( u1_u12_u2_n134 ) );
  NAND3_X1 u1_u12_u2_U98 (.ZN( u1_u12_u2_n110 ) , .A2( u1_u12_u2_n131 ) , .A3( u1_u12_u2_n139 ) , .A1( u1_u12_u2_n154 ) );
  NAND3_X1 u1_u12_u2_U99 (.A2( u1_u12_u2_n100 ) , .ZN( u1_u12_u2_n101 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n114 ) );
  OAI22_X1 u1_u12_u3_U10 (.B1( u1_u12_u3_n113 ) , .A2( u1_u12_u3_n135 ) , .A1( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n164 ) , .ZN( u1_u12_u3_n98 ) );
  OAI211_X1 u1_u12_u3_U11 (.B( u1_u12_u3_n106 ) , .ZN( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n128 ) , .C1( u1_u12_u3_n167 ) , .A( u1_u12_u3_n181 ) );
  AOI221_X1 u1_u12_u3_U12 (.C1( u1_u12_u3_n105 ) , .ZN( u1_u12_u3_n106 ) , .A( u1_u12_u3_n131 ) , .B2( u1_u12_u3_n132 ) , .C2( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n169 ) );
  INV_X1 u1_u12_u3_U13 (.ZN( u1_u12_u3_n181 ) , .A( u1_u12_u3_n98 ) );
  NAND2_X1 u1_u12_u3_U14 (.ZN( u1_u12_u3_n105 ) , .A2( u1_u12_u3_n130 ) , .A1( u1_u12_u3_n155 ) );
  AOI22_X1 u1_u12_u3_U15 (.B1( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n116 ) , .ZN( u1_u12_u3_n123 ) , .B2( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U16 (.ZN( u1_u12_u3_n116 ) , .A2( u1_u12_u3_n151 ) , .A1( u1_u12_u3_n182 ) );
  NOR2_X1 u1_u12_u3_U17 (.ZN( u1_u12_u3_n126 ) , .A2( u1_u12_u3_n150 ) , .A1( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U18 (.ZN( u1_u12_u3_n112 ) , .B2( u1_u12_u3_n146 ) , .B1( u1_u12_u3_n155 ) , .A( u1_u12_u3_n167 ) );
  NAND2_X1 u1_u12_u3_U19 (.A1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n142 ) , .A2( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U20 (.ZN( u1_u12_u3_n132 ) , .A2( u1_u12_u3_n152 ) , .A1( u1_u12_u3_n156 ) );
  AND2_X1 u1_u12_u3_U21 (.A2( u1_u12_u3_n113 ) , .A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n151 ) );
  INV_X1 u1_u12_u3_U22 (.A( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n165 ) );
  INV_X1 u1_u12_u3_U23 (.A( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n170 ) );
  NAND2_X1 u1_u12_u3_U24 (.A1( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .ZN( u1_u12_u3_n140 ) );
  NAND2_X1 u1_u12_u3_U25 (.ZN( u1_u12_u3_n117 ) , .A1( u1_u12_u3_n124 ) , .A2( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U26 (.ZN( u1_u12_u3_n143 ) , .A1( u1_u12_u3_n165 ) , .A2( u1_u12_u3_n167 ) );
  INV_X1 u1_u12_u3_U27 (.A( u1_u12_u3_n130 ) , .ZN( u1_u12_u3_n177 ) );
  INV_X1 u1_u12_u3_U28 (.A( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n176 ) );
  INV_X1 u1_u12_u3_U29 (.A( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n174 ) );
  INV_X1 u1_u12_u3_U3 (.A( u1_u12_u3_n129 ) , .ZN( u1_u12_u3_n183 ) );
  INV_X1 u1_u12_u3_U30 (.A( u1_u12_u3_n139 ) , .ZN( u1_u12_u3_n185 ) );
  NOR2_X1 u1_u12_u3_U31 (.ZN( u1_u12_u3_n135 ) , .A2( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n169 ) );
  OAI222_X1 u1_u12_u3_U32 (.C2( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .B1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n138 ) , .B2( u1_u12_u3_n146 ) , .C1( u1_u12_u3_n154 ) , .A1( u1_u12_u3_n164 ) );
  NOR4_X1 u1_u12_u3_U33 (.A4( u1_u12_u3_n157 ) , .A3( u1_u12_u3_n158 ) , .A2( u1_u12_u3_n159 ) , .A1( u1_u12_u3_n160 ) , .ZN( u1_u12_u3_n161 ) );
  AOI21_X1 u1_u12_u3_U34 (.B2( u1_u12_u3_n152 ) , .B1( u1_u12_u3_n153 ) , .ZN( u1_u12_u3_n158 ) , .A( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U35 (.A( u1_u12_u3_n154 ) , .B2( u1_u12_u3_n155 ) , .B1( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n157 ) );
  AOI21_X1 u1_u12_u3_U36 (.A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n150 ) , .B1( u1_u12_u3_n151 ) , .ZN( u1_u12_u3_n159 ) );
  AOI211_X1 u1_u12_u3_U37 (.ZN( u1_u12_u3_n109 ) , .A( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n129 ) , .B( u1_u12_u3_n138 ) , .C1( u1_u12_u3_n141 ) );
  AOI211_X1 u1_u12_u3_U38 (.B( u1_u12_u3_n119 ) , .A( u1_u12_u3_n120 ) , .C2( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n122 ) , .C1( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U39 (.A( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U4 (.A( u1_u12_u3_n140 ) , .ZN( u1_u12_u3_n182 ) );
  OAI22_X1 u1_u12_u3_U40 (.B1( u1_u12_u3_n118 ) , .ZN( u1_u12_u3_n120 ) , .A1( u1_u12_u3_n135 ) , .B2( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n178 ) );
  AND3_X1 u1_u12_u3_U41 (.ZN( u1_u12_u3_n118 ) , .A2( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n144 ) , .A3( u1_u12_u3_n152 ) );
  INV_X1 u1_u12_u3_U42 (.A( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U43 (.ZN( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n164 ) );
  OAI211_X1 u1_u12_u3_U44 (.B( u1_u12_u3_n127 ) , .ZN( u1_u12_u3_n139 ) , .C1( u1_u12_u3_n150 ) , .C2( u1_u12_u3_n154 ) , .A( u1_u12_u3_n184 ) );
  INV_X1 u1_u12_u3_U45 (.A( u1_u12_u3_n125 ) , .ZN( u1_u12_u3_n184 ) );
  AOI221_X1 u1_u12_u3_U46 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n127 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n169 ) , .B2( u1_u12_u3_n170 ) , .B1( u1_u12_u3_n174 ) );
  OAI22_X1 u1_u12_u3_U47 (.A1( u1_u12_u3_n124 ) , .ZN( u1_u12_u3_n125 ) , .B2( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n165 ) , .B1( u1_u12_u3_n167 ) );
  NOR2_X1 u1_u12_u3_U48 (.A1( u1_u12_u3_n113 ) , .ZN( u1_u12_u3_n131 ) , .A2( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U49 (.A1( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n150 ) , .A2( u1_u12_u3_n99 ) );
  INV_X1 u1_u12_u3_U5 (.A( u1_u12_u3_n117 ) , .ZN( u1_u12_u3_n178 ) );
  NAND2_X1 u1_u12_u3_U50 (.A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n155 ) , .A1( u1_u12_u3_n97 ) );
  INV_X1 u1_u12_u3_U51 (.A( u1_u12_u3_n141 ) , .ZN( u1_u12_u3_n167 ) );
  AOI21_X1 u1_u12_u3_U52 (.B2( u1_u12_u3_n114 ) , .B1( u1_u12_u3_n146 ) , .A( u1_u12_u3_n154 ) , .ZN( u1_u12_u3_n94 ) );
  AOI21_X1 u1_u12_u3_U53 (.ZN( u1_u12_u3_n110 ) , .B2( u1_u12_u3_n142 ) , .B1( u1_u12_u3_n186 ) , .A( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U54 (.A( u1_u12_u3_n145 ) , .ZN( u1_u12_u3_n186 ) );
  AOI21_X1 u1_u12_u3_U55 (.B1( u1_u12_u3_n124 ) , .A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U56 (.A( u1_u12_u3_n149 ) , .ZN( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U57 (.ZN( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n96 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U58 (.A2( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n146 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U59 (.A1( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n99 ) );
  AOI221_X1 u1_u12_u3_U6 (.A( u1_u12_u3_n131 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n134 ) , .B1( u1_u12_u3_n143 ) , .B2( u1_u12_u3_n177 ) );
  NAND2_X1 u1_u12_u3_U60 (.A1( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n156 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U61 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U62 (.A1( u1_u12_u3_n100 ) , .A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n128 ) );
  NAND2_X1 u1_u12_u3_U63 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n152 ) );
  NAND2_X1 u1_u12_u3_U64 (.A2( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n114 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U65 (.ZN( u1_u12_u3_n107 ) , .A1( u1_u12_u3_n97 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U66 (.A2( u1_u12_u3_n100 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n113 ) );
  NAND2_X1 u1_u12_u3_U67 (.A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n153 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U68 (.A2( u1_u12_u3_n103 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n130 ) );
  NAND2_X1 u1_u12_u3_U69 (.A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n96 ) );
  OAI22_X1 u1_u12_u3_U7 (.B2( u1_u12_u3_n147 ) , .A2( u1_u12_u3_n148 ) , .ZN( u1_u12_u3_n160 ) , .B1( u1_u12_u3_n165 ) , .A1( u1_u12_u3_n168 ) );
  NAND2_X1 u1_u12_u3_U70 (.A1( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n108 ) );
  NOR2_X1 u1_u12_u3_U71 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n99 ) );
  NOR2_X1 u1_u12_u3_U72 (.A2( u1_u12_X_21 ) , .A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n103 ) );
  NOR2_X1 u1_u12_u3_U73 (.A2( u1_u12_X_24 ) , .A1( u1_u12_u3_n171 ) , .ZN( u1_u12_u3_n97 ) );
  NOR2_X1 u1_u12_u3_U74 (.A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U75 (.A2( u1_u12_X_19 ) , .A1( u1_u12_u3_n172 ) , .ZN( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U76 (.A1( u1_u12_X_22 ) , .A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U77 (.A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n149 ) , .A2( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U78 (.A2( u1_u12_X_22 ) , .A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n121 ) );
  AND2_X1 u1_u12_u3_U79 (.A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n101 ) , .A2( u1_u12_u3_n171 ) );
  AND3_X1 u1_u12_u3_U8 (.A3( u1_u12_u3_n144 ) , .A2( u1_u12_u3_n145 ) , .A1( u1_u12_u3_n146 ) , .ZN( u1_u12_u3_n147 ) );
  AND2_X1 u1_u12_u3_U80 (.A1( u1_u12_X_19 ) , .ZN( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n172 ) );
  AND2_X1 u1_u12_u3_U81 (.A1( u1_u12_X_21 ) , .A2( u1_u12_X_24 ) , .ZN( u1_u12_u3_n100 ) );
  AND2_X1 u1_u12_u3_U82 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n104 ) );
  INV_X1 u1_u12_u3_U83 (.A( u1_u12_X_22 ) , .ZN( u1_u12_u3_n166 ) );
  INV_X1 u1_u12_u3_U84 (.A( u1_u12_X_21 ) , .ZN( u1_u12_u3_n171 ) );
  INV_X1 u1_u12_u3_U85 (.A( u1_u12_X_20 ) , .ZN( u1_u12_u3_n172 ) );
  NAND4_X1 u1_u12_u3_U86 (.ZN( u1_out12_26 ) , .A4( u1_u12_u3_n109 ) , .A3( u1_u12_u3_n110 ) , .A2( u1_u12_u3_n111 ) , .A1( u1_u12_u3_n173 ) );
  INV_X1 u1_u12_u3_U87 (.ZN( u1_u12_u3_n173 ) , .A( u1_u12_u3_n94 ) );
  OAI21_X1 u1_u12_u3_U88 (.ZN( u1_u12_u3_n111 ) , .B2( u1_u12_u3_n117 ) , .A( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n176 ) );
  NAND4_X1 u1_u12_u3_U89 (.ZN( u1_out12_20 ) , .A4( u1_u12_u3_n122 ) , .A3( u1_u12_u3_n123 ) , .A1( u1_u12_u3_n175 ) , .A2( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U9 (.A( u1_u12_u3_n143 ) , .ZN( u1_u12_u3_n168 ) );
  INV_X1 u1_u12_u3_U90 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U91 (.A( u1_u12_u3_n112 ) , .ZN( u1_u12_u3_n175 ) );
  NAND4_X1 u1_u12_u3_U92 (.ZN( u1_out12_1 ) , .A4( u1_u12_u3_n161 ) , .A3( u1_u12_u3_n162 ) , .A2( u1_u12_u3_n163 ) , .A1( u1_u12_u3_n185 ) );
  NAND2_X1 u1_u12_u3_U93 (.ZN( u1_u12_u3_n163 ) , .A2( u1_u12_u3_n170 ) , .A1( u1_u12_u3_n176 ) );
  AOI22_X1 u1_u12_u3_U94 (.B2( u1_u12_u3_n140 ) , .B1( u1_u12_u3_n141 ) , .A2( u1_u12_u3_n142 ) , .ZN( u1_u12_u3_n162 ) , .A1( u1_u12_u3_n177 ) );
  OR4_X1 u1_u12_u3_U95 (.ZN( u1_out12_10 ) , .A4( u1_u12_u3_n136 ) , .A3( u1_u12_u3_n137 ) , .A1( u1_u12_u3_n138 ) , .A2( u1_u12_u3_n139 ) );
  OAI222_X1 u1_u12_u3_U96 (.C1( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n137 ) , .B1( u1_u12_u3_n148 ) , .A2( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n154 ) , .C2( u1_u12_u3_n164 ) , .A1( u1_u12_u3_n167 ) );
  OAI221_X1 u1_u12_u3_U97 (.A( u1_u12_u3_n134 ) , .B2( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n136 ) , .C1( u1_u12_u3_n149 ) , .B1( u1_u12_u3_n151 ) , .C2( u1_u12_u3_n183 ) );
  NAND3_X1 u1_u12_u3_U98 (.A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n145 ) , .A3( u1_u12_u3_n153 ) );
  NAND3_X1 u1_u12_u3_U99 (.ZN( u1_u12_u3_n129 ) , .A2( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n153 ) , .A3( u1_u12_u3_n182 ) );
  AND3_X1 u1_u12_u7_U10 (.A3( u1_u12_u7_n110 ) , .A2( u1_u12_u7_n127 ) , .A1( u1_u12_u7_n132 ) , .ZN( u1_u12_u7_n92 ) );
  OAI21_X1 u1_u12_u7_U11 (.A( u1_u12_u7_n161 ) , .B1( u1_u12_u7_n168 ) , .B2( u1_u12_u7_n173 ) , .ZN( u1_u12_u7_n91 ) );
  AOI211_X1 u1_u12_u7_U12 (.A( u1_u12_u7_n117 ) , .ZN( u1_u12_u7_n118 ) , .C2( u1_u12_u7_n126 ) , .C1( u1_u12_u7_n177 ) , .B( u1_u12_u7_n180 ) );
  OAI22_X1 u1_u12_u7_U13 (.B1( u1_u12_u7_n115 ) , .ZN( u1_u12_u7_n117 ) , .A2( u1_u12_u7_n133 ) , .A1( u1_u12_u7_n137 ) , .B2( u1_u12_u7_n162 ) );
  INV_X1 u1_u12_u7_U14 (.A( u1_u12_u7_n116 ) , .ZN( u1_u12_u7_n180 ) );
  NOR3_X1 u1_u12_u7_U15 (.ZN( u1_u12_u7_n115 ) , .A3( u1_u12_u7_n145 ) , .A2( u1_u12_u7_n168 ) , .A1( u1_u12_u7_n169 ) );
  OAI211_X1 u1_u12_u7_U16 (.B( u1_u12_u7_n122 ) , .A( u1_u12_u7_n123 ) , .C2( u1_u12_u7_n124 ) , .ZN( u1_u12_u7_n154 ) , .C1( u1_u12_u7_n162 ) );
  AOI222_X1 u1_u12_u7_U17 (.ZN( u1_u12_u7_n122 ) , .C2( u1_u12_u7_n126 ) , .C1( u1_u12_u7_n145 ) , .B1( u1_u12_u7_n161 ) , .A2( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n170 ) , .A1( u1_u12_u7_n176 ) );
  INV_X1 u1_u12_u7_U18 (.A( u1_u12_u7_n133 ) , .ZN( u1_u12_u7_n176 ) );
  NOR3_X1 u1_u12_u7_U19 (.A2( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n135 ) , .ZN( u1_u12_u7_n136 ) , .A3( u1_u12_u7_n171 ) );
  NOR2_X1 u1_u12_u7_U20 (.A1( u1_u12_u7_n130 ) , .A2( u1_u12_u7_n134 ) , .ZN( u1_u12_u7_n153 ) );
  INV_X1 u1_u12_u7_U21 (.A( u1_u12_u7_n101 ) , .ZN( u1_u12_u7_n165 ) );
  NOR2_X1 u1_u12_u7_U22 (.ZN( u1_u12_u7_n111 ) , .A2( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n169 ) );
  AOI21_X1 u1_u12_u7_U23 (.ZN( u1_u12_u7_n104 ) , .B2( u1_u12_u7_n112 ) , .B1( u1_u12_u7_n127 ) , .A( u1_u12_u7_n164 ) );
  AOI21_X1 u1_u12_u7_U24 (.ZN( u1_u12_u7_n106 ) , .B1( u1_u12_u7_n133 ) , .B2( u1_u12_u7_n146 ) , .A( u1_u12_u7_n162 ) );
  AOI21_X1 u1_u12_u7_U25 (.A( u1_u12_u7_n101 ) , .ZN( u1_u12_u7_n107 ) , .B2( u1_u12_u7_n128 ) , .B1( u1_u12_u7_n175 ) );
  INV_X1 u1_u12_u7_U26 (.A( u1_u12_u7_n138 ) , .ZN( u1_u12_u7_n171 ) );
  INV_X1 u1_u12_u7_U27 (.A( u1_u12_u7_n131 ) , .ZN( u1_u12_u7_n177 ) );
  INV_X1 u1_u12_u7_U28 (.A( u1_u12_u7_n110 ) , .ZN( u1_u12_u7_n174 ) );
  NAND2_X1 u1_u12_u7_U29 (.A1( u1_u12_u7_n129 ) , .A2( u1_u12_u7_n132 ) , .ZN( u1_u12_u7_n149 ) );
  OAI21_X1 u1_u12_u7_U3 (.ZN( u1_u12_u7_n159 ) , .A( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n171 ) , .B1( u1_u12_u7_n174 ) );
  NAND2_X1 u1_u12_u7_U30 (.A1( u1_u12_u7_n113 ) , .A2( u1_u12_u7_n124 ) , .ZN( u1_u12_u7_n130 ) );
  INV_X1 u1_u12_u7_U31 (.A( u1_u12_u7_n112 ) , .ZN( u1_u12_u7_n173 ) );
  INV_X1 u1_u12_u7_U32 (.A( u1_u12_u7_n128 ) , .ZN( u1_u12_u7_n168 ) );
  INV_X1 u1_u12_u7_U33 (.A( u1_u12_u7_n148 ) , .ZN( u1_u12_u7_n169 ) );
  INV_X1 u1_u12_u7_U34 (.A( u1_u12_u7_n127 ) , .ZN( u1_u12_u7_n179 ) );
  NOR2_X1 u1_u12_u7_U35 (.ZN( u1_u12_u7_n101 ) , .A2( u1_u12_u7_n150 ) , .A1( u1_u12_u7_n156 ) );
  AOI211_X1 u1_u12_u7_U36 (.B( u1_u12_u7_n154 ) , .A( u1_u12_u7_n155 ) , .C1( u1_u12_u7_n156 ) , .ZN( u1_u12_u7_n157 ) , .C2( u1_u12_u7_n172 ) );
  INV_X1 u1_u12_u7_U37 (.A( u1_u12_u7_n153 ) , .ZN( u1_u12_u7_n172 ) );
  AOI211_X1 u1_u12_u7_U38 (.B( u1_u12_u7_n139 ) , .A( u1_u12_u7_n140 ) , .C2( u1_u12_u7_n141 ) , .ZN( u1_u12_u7_n142 ) , .C1( u1_u12_u7_n156 ) );
  NAND4_X1 u1_u12_u7_U39 (.A3( u1_u12_u7_n127 ) , .A2( u1_u12_u7_n128 ) , .A1( u1_u12_u7_n129 ) , .ZN( u1_u12_u7_n141 ) , .A4( u1_u12_u7_n147 ) );
  INV_X1 u1_u12_u7_U4 (.A( u1_u12_u7_n111 ) , .ZN( u1_u12_u7_n170 ) );
  AOI21_X1 u1_u12_u7_U40 (.A( u1_u12_u7_n137 ) , .B1( u1_u12_u7_n138 ) , .ZN( u1_u12_u7_n139 ) , .B2( u1_u12_u7_n146 ) );
  OAI22_X1 u1_u12_u7_U41 (.B1( u1_u12_u7_n136 ) , .ZN( u1_u12_u7_n140 ) , .A1( u1_u12_u7_n153 ) , .B2( u1_u12_u7_n162 ) , .A2( u1_u12_u7_n164 ) );
  AOI21_X1 u1_u12_u7_U42 (.ZN( u1_u12_u7_n123 ) , .B1( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n177 ) , .A( u1_u12_u7_n97 ) );
  AOI21_X1 u1_u12_u7_U43 (.B2( u1_u12_u7_n113 ) , .B1( u1_u12_u7_n124 ) , .A( u1_u12_u7_n125 ) , .ZN( u1_u12_u7_n97 ) );
  INV_X1 u1_u12_u7_U44 (.A( u1_u12_u7_n125 ) , .ZN( u1_u12_u7_n161 ) );
  INV_X1 u1_u12_u7_U45 (.A( u1_u12_u7_n152 ) , .ZN( u1_u12_u7_n162 ) );
  AOI22_X1 u1_u12_u7_U46 (.A2( u1_u12_u7_n114 ) , .ZN( u1_u12_u7_n119 ) , .B1( u1_u12_u7_n130 ) , .A1( u1_u12_u7_n156 ) , .B2( u1_u12_u7_n165 ) );
  NAND2_X1 u1_u12_u7_U47 (.A2( u1_u12_u7_n112 ) , .ZN( u1_u12_u7_n114 ) , .A1( u1_u12_u7_n175 ) );
  AND2_X1 u1_u12_u7_U48 (.ZN( u1_u12_u7_n145 ) , .A2( u1_u12_u7_n98 ) , .A1( u1_u12_u7_n99 ) );
  NOR2_X1 u1_u12_u7_U49 (.ZN( u1_u12_u7_n137 ) , .A1( u1_u12_u7_n150 ) , .A2( u1_u12_u7_n161 ) );
  INV_X1 u1_u12_u7_U5 (.A( u1_u12_u7_n149 ) , .ZN( u1_u12_u7_n175 ) );
  AOI21_X1 u1_u12_u7_U50 (.ZN( u1_u12_u7_n105 ) , .B2( u1_u12_u7_n110 ) , .A( u1_u12_u7_n125 ) , .B1( u1_u12_u7_n147 ) );
  NAND2_X1 u1_u12_u7_U51 (.ZN( u1_u12_u7_n146 ) , .A1( u1_u12_u7_n95 ) , .A2( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U52 (.A2( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n147 ) , .A1( u1_u12_u7_n93 ) );
  NAND2_X1 u1_u12_u7_U53 (.A1( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n127 ) , .A2( u1_u12_u7_n99 ) );
  OR2_X1 u1_u12_u7_U54 (.ZN( u1_u12_u7_n126 ) , .A2( u1_u12_u7_n152 ) , .A1( u1_u12_u7_n156 ) );
  NAND2_X1 u1_u12_u7_U55 (.A2( u1_u12_u7_n102 ) , .A1( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n133 ) );
  NAND2_X1 u1_u12_u7_U56 (.ZN( u1_u12_u7_n112 ) , .A2( u1_u12_u7_n96 ) , .A1( u1_u12_u7_n99 ) );
  NAND2_X1 u1_u12_u7_U57 (.A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n128 ) , .A1( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U58 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n113 ) , .A2( u1_u12_u7_n93 ) );
  NAND2_X1 u1_u12_u7_U59 (.A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n124 ) , .A1( u1_u12_u7_n96 ) );
  INV_X1 u1_u12_u7_U6 (.A( u1_u12_u7_n154 ) , .ZN( u1_u12_u7_n178 ) );
  NAND2_X1 u1_u12_u7_U60 (.ZN( u1_u12_u7_n110 ) , .A1( u1_u12_u7_n95 ) , .A2( u1_u12_u7_n96 ) );
  INV_X1 u1_u12_u7_U61 (.A( u1_u12_u7_n150 ) , .ZN( u1_u12_u7_n164 ) );
  AND2_X1 u1_u12_u7_U62 (.ZN( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n93 ) , .A2( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U63 (.A1( u1_u12_u7_n100 ) , .A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n129 ) );
  NAND2_X1 u1_u12_u7_U64 (.A2( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n131 ) , .A1( u1_u12_u7_n95 ) );
  NAND2_X1 u1_u12_u7_U65 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n138 ) , .A2( u1_u12_u7_n99 ) );
  NAND2_X1 u1_u12_u7_U66 (.ZN( u1_u12_u7_n132 ) , .A1( u1_u12_u7_n93 ) , .A2( u1_u12_u7_n96 ) );
  NAND2_X1 u1_u12_u7_U67 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n148 ) , .A2( u1_u12_u7_n95 ) );
  NOR2_X1 u1_u12_u7_U68 (.A2( u1_u12_X_47 ) , .ZN( u1_u12_u7_n150 ) , .A1( u1_u12_u7_n163 ) );
  NOR2_X1 u1_u12_u7_U69 (.A2( u1_u12_X_43 ) , .A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n103 ) );
  AOI211_X1 u1_u12_u7_U7 (.ZN( u1_u12_u7_n116 ) , .A( u1_u12_u7_n155 ) , .C1( u1_u12_u7_n161 ) , .C2( u1_u12_u7_n171 ) , .B( u1_u12_u7_n94 ) );
  NOR2_X1 u1_u12_u7_U70 (.A2( u1_u12_X_48 ) , .A1( u1_u12_u7_n166 ) , .ZN( u1_u12_u7_n95 ) );
  NOR2_X1 u1_u12_u7_U71 (.A2( u1_u12_X_45 ) , .A1( u1_u12_X_48 ) , .ZN( u1_u12_u7_n99 ) );
  NOR2_X1 u1_u12_u7_U72 (.A2( u1_u12_X_44 ) , .A1( u1_u12_u7_n167 ) , .ZN( u1_u12_u7_n98 ) );
  NOR2_X1 u1_u12_u7_U73 (.A2( u1_u12_X_46 ) , .A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n152 ) );
  AND2_X1 u1_u12_u7_U74 (.A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n156 ) , .A2( u1_u12_u7_n163 ) );
  NAND2_X1 u1_u12_u7_U75 (.A2( u1_u12_X_46 ) , .A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n125 ) );
  AND2_X1 u1_u12_u7_U76 (.A2( u1_u12_X_45 ) , .A1( u1_u12_X_48 ) , .ZN( u1_u12_u7_n102 ) );
  AND2_X1 u1_u12_u7_U77 (.A2( u1_u12_X_43 ) , .A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n96 ) );
  AND2_X1 u1_u12_u7_U78 (.A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n100 ) , .A2( u1_u12_u7_n167 ) );
  AND2_X1 u1_u12_u7_U79 (.A1( u1_u12_X_48 ) , .A2( u1_u12_u7_n166 ) , .ZN( u1_u12_u7_n93 ) );
  OAI222_X1 u1_u12_u7_U8 (.C2( u1_u12_u7_n101 ) , .B2( u1_u12_u7_n111 ) , .A1( u1_u12_u7_n113 ) , .C1( u1_u12_u7_n146 ) , .A2( u1_u12_u7_n162 ) , .B1( u1_u12_u7_n164 ) , .ZN( u1_u12_u7_n94 ) );
  INV_X1 u1_u12_u7_U80 (.A( u1_u12_X_46 ) , .ZN( u1_u12_u7_n163 ) );
  INV_X1 u1_u12_u7_U81 (.A( u1_u12_X_43 ) , .ZN( u1_u12_u7_n167 ) );
  INV_X1 u1_u12_u7_U82 (.A( u1_u12_X_45 ) , .ZN( u1_u12_u7_n166 ) );
  NAND4_X1 u1_u12_u7_U83 (.ZN( u1_out12_5 ) , .A4( u1_u12_u7_n108 ) , .A3( u1_u12_u7_n109 ) , .A1( u1_u12_u7_n116 ) , .A2( u1_u12_u7_n123 ) );
  AOI22_X1 u1_u12_u7_U84 (.ZN( u1_u12_u7_n109 ) , .A2( u1_u12_u7_n126 ) , .B2( u1_u12_u7_n145 ) , .B1( u1_u12_u7_n156 ) , .A1( u1_u12_u7_n171 ) );
  NOR4_X1 u1_u12_u7_U85 (.A4( u1_u12_u7_n104 ) , .A3( u1_u12_u7_n105 ) , .A2( u1_u12_u7_n106 ) , .A1( u1_u12_u7_n107 ) , .ZN( u1_u12_u7_n108 ) );
  NAND4_X1 u1_u12_u7_U86 (.ZN( u1_out12_27 ) , .A4( u1_u12_u7_n118 ) , .A3( u1_u12_u7_n119 ) , .A2( u1_u12_u7_n120 ) , .A1( u1_u12_u7_n121 ) );
  OAI21_X1 u1_u12_u7_U87 (.ZN( u1_u12_u7_n121 ) , .B2( u1_u12_u7_n145 ) , .A( u1_u12_u7_n150 ) , .B1( u1_u12_u7_n174 ) );
  OAI21_X1 u1_u12_u7_U88 (.ZN( u1_u12_u7_n120 ) , .A( u1_u12_u7_n161 ) , .B2( u1_u12_u7_n170 ) , .B1( u1_u12_u7_n179 ) );
  NAND4_X1 u1_u12_u7_U89 (.ZN( u1_out12_21 ) , .A4( u1_u12_u7_n157 ) , .A3( u1_u12_u7_n158 ) , .A2( u1_u12_u7_n159 ) , .A1( u1_u12_u7_n160 ) );
  OAI221_X1 u1_u12_u7_U9 (.C1( u1_u12_u7_n101 ) , .C2( u1_u12_u7_n147 ) , .ZN( u1_u12_u7_n155 ) , .B2( u1_u12_u7_n162 ) , .A( u1_u12_u7_n91 ) , .B1( u1_u12_u7_n92 ) );
  OAI21_X1 u1_u12_u7_U90 (.B1( u1_u12_u7_n145 ) , .ZN( u1_u12_u7_n160 ) , .A( u1_u12_u7_n161 ) , .B2( u1_u12_u7_n177 ) );
  AOI22_X1 u1_u12_u7_U91 (.B2( u1_u12_u7_n149 ) , .B1( u1_u12_u7_n150 ) , .A2( u1_u12_u7_n151 ) , .A1( u1_u12_u7_n152 ) , .ZN( u1_u12_u7_n158 ) );
  NAND4_X1 u1_u12_u7_U92 (.ZN( u1_out12_15 ) , .A4( u1_u12_u7_n142 ) , .A3( u1_u12_u7_n143 ) , .A2( u1_u12_u7_n144 ) , .A1( u1_u12_u7_n178 ) );
  OR2_X1 u1_u12_u7_U93 (.A2( u1_u12_u7_n125 ) , .A1( u1_u12_u7_n129 ) , .ZN( u1_u12_u7_n144 ) );
  AOI22_X1 u1_u12_u7_U94 (.A2( u1_u12_u7_n126 ) , .ZN( u1_u12_u7_n143 ) , .B2( u1_u12_u7_n165 ) , .B1( u1_u12_u7_n173 ) , .A1( u1_u12_u7_n174 ) );
  NAND3_X1 u1_u12_u7_U95 (.A3( u1_u12_u7_n146 ) , .A2( u1_u12_u7_n147 ) , .A1( u1_u12_u7_n148 ) , .ZN( u1_u12_u7_n151 ) );
  NAND3_X1 u1_u12_u7_U96 (.A3( u1_u12_u7_n131 ) , .A2( u1_u12_u7_n132 ) , .A1( u1_u12_u7_n133 ) , .ZN( u1_u12_u7_n135 ) );
  XOR2_X1 u1_u13_U11 (.B( u1_K14_44 ) , .A( u1_R12_29 ) , .Z( u1_u13_X_44 ) );
  XOR2_X1 u1_u13_U13 (.B( u1_K14_42 ) , .A( u1_R12_29 ) , .Z( u1_u13_X_42 ) );
  XOR2_X1 u1_u13_U27 (.B( u1_K14_2 ) , .A( u1_R12_1 ) , .Z( u1_u13_X_2 ) );
  XOR2_X1 u1_u13_U38 (.B( u1_K14_1 ) , .A( u1_R12_32 ) , .Z( u1_u13_X_1 ) );
  XOR2_X1 u1_u13_U7 (.B( u1_K14_48 ) , .A( u1_R12_1 ) , .Z( u1_u13_X_48 ) );
  XOR2_X1 u1_u13_U8 (.B( u1_K14_47 ) , .A( u1_R12_32 ) , .Z( u1_u13_X_47 ) );
  AND3_X1 u1_u13_u0_U10 (.A2( u1_u13_u0_n112 ) , .ZN( u1_u13_u0_n127 ) , .A3( u1_u13_u0_n130 ) , .A1( u1_u13_u0_n148 ) );
  NAND2_X1 u1_u13_u0_U11 (.ZN( u1_u13_u0_n113 ) , .A1( u1_u13_u0_n139 ) , .A2( u1_u13_u0_n149 ) );
  AND2_X1 u1_u13_u0_U12 (.ZN( u1_u13_u0_n107 ) , .A1( u1_u13_u0_n130 ) , .A2( u1_u13_u0_n140 ) );
  AND2_X1 u1_u13_u0_U13 (.A2( u1_u13_u0_n129 ) , .A1( u1_u13_u0_n130 ) , .ZN( u1_u13_u0_n151 ) );
  AND2_X1 u1_u13_u0_U14 (.A1( u1_u13_u0_n108 ) , .A2( u1_u13_u0_n125 ) , .ZN( u1_u13_u0_n145 ) );
  INV_X1 u1_u13_u0_U15 (.A( u1_u13_u0_n143 ) , .ZN( u1_u13_u0_n173 ) );
  NOR2_X1 u1_u13_u0_U16 (.A2( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n147 ) , .A1( u1_u13_u0_n160 ) );
  INV_X1 u1_u13_u0_U17 (.ZN( u1_u13_u0_n172 ) , .A( u1_u13_u0_n88 ) );
  OAI222_X1 u1_u13_u0_U18 (.C1( u1_u13_u0_n108 ) , .A1( u1_u13_u0_n125 ) , .B2( u1_u13_u0_n128 ) , .B1( u1_u13_u0_n144 ) , .A2( u1_u13_u0_n158 ) , .C2( u1_u13_u0_n161 ) , .ZN( u1_u13_u0_n88 ) );
  NOR2_X1 u1_u13_u0_U19 (.A1( u1_u13_u0_n163 ) , .A2( u1_u13_u0_n164 ) , .ZN( u1_u13_u0_n95 ) );
  AOI21_X1 u1_u13_u0_U20 (.B1( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n132 ) , .A( u1_u13_u0_n165 ) , .B2( u1_u13_u0_n93 ) );
  INV_X1 u1_u13_u0_U21 (.A( u1_u13_u0_n142 ) , .ZN( u1_u13_u0_n165 ) );
  OAI221_X1 u1_u13_u0_U22 (.C1( u1_u13_u0_n121 ) , .ZN( u1_u13_u0_n122 ) , .B2( u1_u13_u0_n127 ) , .A( u1_u13_u0_n143 ) , .B1( u1_u13_u0_n144 ) , .C2( u1_u13_u0_n147 ) );
  OAI22_X1 u1_u13_u0_U23 (.B1( u1_u13_u0_n125 ) , .ZN( u1_u13_u0_n126 ) , .A1( u1_u13_u0_n138 ) , .A2( u1_u13_u0_n146 ) , .B2( u1_u13_u0_n147 ) );
  OAI22_X1 u1_u13_u0_U24 (.B1( u1_u13_u0_n131 ) , .A1( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n147 ) , .A2( u1_u13_u0_n90 ) , .ZN( u1_u13_u0_n91 ) );
  AND3_X1 u1_u13_u0_U25 (.A3( u1_u13_u0_n121 ) , .A2( u1_u13_u0_n125 ) , .A1( u1_u13_u0_n148 ) , .ZN( u1_u13_u0_n90 ) );
  INV_X1 u1_u13_u0_U26 (.A( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n161 ) );
  NOR2_X1 u1_u13_u0_U27 (.A1( u1_u13_u0_n120 ) , .ZN( u1_u13_u0_n143 ) , .A2( u1_u13_u0_n167 ) );
  OAI221_X1 u1_u13_u0_U28 (.C1( u1_u13_u0_n112 ) , .ZN( u1_u13_u0_n120 ) , .B1( u1_u13_u0_n138 ) , .B2( u1_u13_u0_n141 ) , .C2( u1_u13_u0_n147 ) , .A( u1_u13_u0_n172 ) );
  AOI211_X1 u1_u13_u0_U29 (.B( u1_u13_u0_n115 ) , .A( u1_u13_u0_n116 ) , .C2( u1_u13_u0_n117 ) , .C1( u1_u13_u0_n118 ) , .ZN( u1_u13_u0_n119 ) );
  INV_X1 u1_u13_u0_U3 (.A( u1_u13_u0_n113 ) , .ZN( u1_u13_u0_n166 ) );
  AOI22_X1 u1_u13_u0_U30 (.B2( u1_u13_u0_n109 ) , .A2( u1_u13_u0_n110 ) , .ZN( u1_u13_u0_n111 ) , .B1( u1_u13_u0_n118 ) , .A1( u1_u13_u0_n160 ) );
  INV_X1 u1_u13_u0_U31 (.A( u1_u13_u0_n118 ) , .ZN( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U32 (.ZN( u1_u13_u0_n104 ) , .B1( u1_u13_u0_n107 ) , .B2( u1_u13_u0_n141 ) , .A( u1_u13_u0_n144 ) );
  AOI21_X1 u1_u13_u0_U33 (.B1( u1_u13_u0_n127 ) , .B2( u1_u13_u0_n129 ) , .A( u1_u13_u0_n138 ) , .ZN( u1_u13_u0_n96 ) );
  AOI21_X1 u1_u13_u0_U34 (.ZN( u1_u13_u0_n116 ) , .B2( u1_u13_u0_n142 ) , .A( u1_u13_u0_n144 ) , .B1( u1_u13_u0_n166 ) );
  NAND2_X1 u1_u13_u0_U35 (.A1( u1_u13_u0_n100 ) , .A2( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n125 ) );
  NAND2_X1 u1_u13_u0_U36 (.A1( u1_u13_u0_n101 ) , .A2( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n150 ) );
  INV_X1 u1_u13_u0_U37 (.A( u1_u13_u0_n138 ) , .ZN( u1_u13_u0_n160 ) );
  NAND2_X1 u1_u13_u0_U38 (.A1( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n128 ) , .A2( u1_u13_u0_n95 ) );
  NAND2_X1 u1_u13_u0_U39 (.A1( u1_u13_u0_n100 ) , .ZN( u1_u13_u0_n129 ) , .A2( u1_u13_u0_n95 ) );
  AOI21_X1 u1_u13_u0_U4 (.B1( u1_u13_u0_n114 ) , .ZN( u1_u13_u0_n115 ) , .B2( u1_u13_u0_n129 ) , .A( u1_u13_u0_n161 ) );
  NAND2_X1 u1_u13_u0_U40 (.A2( u1_u13_u0_n100 ) , .ZN( u1_u13_u0_n131 ) , .A1( u1_u13_u0_n92 ) );
  NAND2_X1 u1_u13_u0_U41 (.A2( u1_u13_u0_n100 ) , .A1( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n139 ) );
  NAND2_X1 u1_u13_u0_U42 (.ZN( u1_u13_u0_n148 ) , .A1( u1_u13_u0_n93 ) , .A2( u1_u13_u0_n95 ) );
  NAND2_X1 u1_u13_u0_U43 (.A2( u1_u13_u0_n102 ) , .A1( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n149 ) );
  NAND2_X1 u1_u13_u0_U44 (.A2( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n114 ) , .A1( u1_u13_u0_n92 ) );
  NAND2_X1 u1_u13_u0_U45 (.A2( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n121 ) , .A1( u1_u13_u0_n93 ) );
  NAND2_X1 u1_u13_u0_U46 (.ZN( u1_u13_u0_n112 ) , .A2( u1_u13_u0_n92 ) , .A1( u1_u13_u0_n93 ) );
  OR3_X1 u1_u13_u0_U47 (.A3( u1_u13_u0_n152 ) , .A2( u1_u13_u0_n153 ) , .A1( u1_u13_u0_n154 ) , .ZN( u1_u13_u0_n155 ) );
  AOI21_X1 u1_u13_u0_U48 (.B2( u1_u13_u0_n150 ) , .B1( u1_u13_u0_n151 ) , .ZN( u1_u13_u0_n152 ) , .A( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U49 (.A( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n145 ) , .B1( u1_u13_u0_n146 ) , .ZN( u1_u13_u0_n154 ) );
  AOI21_X1 u1_u13_u0_U5 (.B2( u1_u13_u0_n131 ) , .ZN( u1_u13_u0_n134 ) , .B1( u1_u13_u0_n151 ) , .A( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U50 (.A( u1_u13_u0_n147 ) , .B2( u1_u13_u0_n148 ) , .B1( u1_u13_u0_n149 ) , .ZN( u1_u13_u0_n153 ) );
  INV_X1 u1_u13_u0_U51 (.ZN( u1_u13_u0_n171 ) , .A( u1_u13_u0_n99 ) );
  OAI211_X1 u1_u13_u0_U52 (.C2( u1_u13_u0_n140 ) , .C1( u1_u13_u0_n161 ) , .A( u1_u13_u0_n169 ) , .B( u1_u13_u0_n98 ) , .ZN( u1_u13_u0_n99 ) );
  AOI211_X1 u1_u13_u0_U53 (.C1( u1_u13_u0_n118 ) , .A( u1_u13_u0_n123 ) , .B( u1_u13_u0_n96 ) , .C2( u1_u13_u0_n97 ) , .ZN( u1_u13_u0_n98 ) );
  INV_X1 u1_u13_u0_U54 (.ZN( u1_u13_u0_n169 ) , .A( u1_u13_u0_n91 ) );
  NOR2_X1 u1_u13_u0_U55 (.A2( u1_u13_X_6 ) , .ZN( u1_u13_u0_n100 ) , .A1( u1_u13_u0_n162 ) );
  NOR2_X1 u1_u13_u0_U56 (.A2( u1_u13_X_4 ) , .A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n118 ) );
  NOR2_X1 u1_u13_u0_U57 (.A2( u1_u13_X_2 ) , .ZN( u1_u13_u0_n103 ) , .A1( u1_u13_u0_n164 ) );
  NOR2_X1 u1_u13_u0_U58 (.A2( u1_u13_X_1 ) , .A1( u1_u13_X_2 ) , .ZN( u1_u13_u0_n92 ) );
  NOR2_X1 u1_u13_u0_U59 (.A2( u1_u13_X_1 ) , .ZN( u1_u13_u0_n101 ) , .A1( u1_u13_u0_n163 ) );
  NOR2_X1 u1_u13_u0_U6 (.A1( u1_u13_u0_n108 ) , .ZN( u1_u13_u0_n123 ) , .A2( u1_u13_u0_n158 ) );
  NAND2_X1 u1_u13_u0_U60 (.A2( u1_u13_X_4 ) , .A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n144 ) );
  NOR2_X1 u1_u13_u0_U61 (.A2( u1_u13_X_5 ) , .ZN( u1_u13_u0_n136 ) , .A1( u1_u13_u0_n159 ) );
  NAND2_X1 u1_u13_u0_U62 (.A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n138 ) , .A2( u1_u13_u0_n159 ) );
  AND2_X1 u1_u13_u0_U63 (.A2( u1_u13_X_3 ) , .A1( u1_u13_X_6 ) , .ZN( u1_u13_u0_n102 ) );
  AND2_X1 u1_u13_u0_U64 (.A1( u1_u13_X_6 ) , .A2( u1_u13_u0_n162 ) , .ZN( u1_u13_u0_n93 ) );
  INV_X1 u1_u13_u0_U65 (.A( u1_u13_X_4 ) , .ZN( u1_u13_u0_n159 ) );
  INV_X1 u1_u13_u0_U66 (.A( u1_u13_X_1 ) , .ZN( u1_u13_u0_n164 ) );
  INV_X1 u1_u13_u0_U67 (.A( u1_u13_X_2 ) , .ZN( u1_u13_u0_n163 ) );
  INV_X1 u1_u13_u0_U68 (.A( u1_u13_u0_n126 ) , .ZN( u1_u13_u0_n168 ) );
  AOI211_X1 u1_u13_u0_U69 (.B( u1_u13_u0_n133 ) , .A( u1_u13_u0_n134 ) , .C2( u1_u13_u0_n135 ) , .C1( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n137 ) );
  OAI21_X1 u1_u13_u0_U7 (.B1( u1_u13_u0_n150 ) , .B2( u1_u13_u0_n158 ) , .A( u1_u13_u0_n172 ) , .ZN( u1_u13_u0_n89 ) );
  INV_X1 u1_u13_u0_U70 (.ZN( u1_u13_u0_n174 ) , .A( u1_u13_u0_n89 ) );
  AOI211_X1 u1_u13_u0_U71 (.B( u1_u13_u0_n104 ) , .A( u1_u13_u0_n105 ) , .ZN( u1_u13_u0_n106 ) , .C2( u1_u13_u0_n113 ) , .C1( u1_u13_u0_n160 ) );
  OR4_X1 u1_u13_u0_U72 (.ZN( u1_out13_17 ) , .A4( u1_u13_u0_n122 ) , .A2( u1_u13_u0_n123 ) , .A1( u1_u13_u0_n124 ) , .A3( u1_u13_u0_n170 ) );
  AOI21_X1 u1_u13_u0_U73 (.B2( u1_u13_u0_n107 ) , .ZN( u1_u13_u0_n124 ) , .B1( u1_u13_u0_n128 ) , .A( u1_u13_u0_n161 ) );
  INV_X1 u1_u13_u0_U74 (.A( u1_u13_u0_n111 ) , .ZN( u1_u13_u0_n170 ) );
  OR4_X1 u1_u13_u0_U75 (.ZN( u1_out13_31 ) , .A4( u1_u13_u0_n155 ) , .A2( u1_u13_u0_n156 ) , .A1( u1_u13_u0_n157 ) , .A3( u1_u13_u0_n173 ) );
  AOI21_X1 u1_u13_u0_U76 (.A( u1_u13_u0_n138 ) , .B2( u1_u13_u0_n139 ) , .B1( u1_u13_u0_n140 ) , .ZN( u1_u13_u0_n157 ) );
  AOI21_X1 u1_u13_u0_U77 (.B2( u1_u13_u0_n141 ) , .B1( u1_u13_u0_n142 ) , .ZN( u1_u13_u0_n156 ) , .A( u1_u13_u0_n161 ) );
  AOI21_X1 u1_u13_u0_U78 (.B1( u1_u13_u0_n132 ) , .ZN( u1_u13_u0_n133 ) , .A( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n166 ) );
  OAI22_X1 u1_u13_u0_U79 (.ZN( u1_u13_u0_n105 ) , .A2( u1_u13_u0_n132 ) , .B1( u1_u13_u0_n146 ) , .A1( u1_u13_u0_n147 ) , .B2( u1_u13_u0_n161 ) );
  AND2_X1 u1_u13_u0_U8 (.A1( u1_u13_u0_n114 ) , .A2( u1_u13_u0_n121 ) , .ZN( u1_u13_u0_n146 ) );
  NAND2_X1 u1_u13_u0_U80 (.ZN( u1_u13_u0_n110 ) , .A2( u1_u13_u0_n132 ) , .A1( u1_u13_u0_n145 ) );
  INV_X1 u1_u13_u0_U81 (.A( u1_u13_u0_n119 ) , .ZN( u1_u13_u0_n167 ) );
  NAND2_X1 u1_u13_u0_U82 (.A2( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n140 ) , .A1( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U83 (.A1( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n130 ) , .A2( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U84 (.ZN( u1_u13_u0_n108 ) , .A1( u1_u13_u0_n92 ) , .A2( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U85 (.ZN( u1_u13_u0_n142 ) , .A1( u1_u13_u0_n94 ) , .A2( u1_u13_u0_n95 ) );
  INV_X1 u1_u13_u0_U86 (.A( u1_u13_X_3 ) , .ZN( u1_u13_u0_n162 ) );
  NOR2_X1 u1_u13_u0_U87 (.A2( u1_u13_X_3 ) , .A1( u1_u13_X_6 ) , .ZN( u1_u13_u0_n94 ) );
  NAND3_X1 u1_u13_u0_U88 (.ZN( u1_out13_23 ) , .A3( u1_u13_u0_n137 ) , .A1( u1_u13_u0_n168 ) , .A2( u1_u13_u0_n171 ) );
  NAND3_X1 u1_u13_u0_U89 (.A3( u1_u13_u0_n127 ) , .A2( u1_u13_u0_n128 ) , .ZN( u1_u13_u0_n135 ) , .A1( u1_u13_u0_n150 ) );
  AND2_X1 u1_u13_u0_U9 (.A1( u1_u13_u0_n131 ) , .ZN( u1_u13_u0_n141 ) , .A2( u1_u13_u0_n150 ) );
  NAND3_X1 u1_u13_u0_U90 (.ZN( u1_u13_u0_n117 ) , .A3( u1_u13_u0_n132 ) , .A2( u1_u13_u0_n139 ) , .A1( u1_u13_u0_n148 ) );
  NAND3_X1 u1_u13_u0_U91 (.ZN( u1_u13_u0_n109 ) , .A2( u1_u13_u0_n114 ) , .A3( u1_u13_u0_n140 ) , .A1( u1_u13_u0_n149 ) );
  NAND3_X1 u1_u13_u0_U92 (.ZN( u1_out13_9 ) , .A3( u1_u13_u0_n106 ) , .A2( u1_u13_u0_n171 ) , .A1( u1_u13_u0_n174 ) );
  NAND3_X1 u1_u13_u0_U93 (.A2( u1_u13_u0_n128 ) , .A1( u1_u13_u0_n132 ) , .A3( u1_u13_u0_n146 ) , .ZN( u1_u13_u0_n97 ) );
  NAND2_X1 u1_u13_u1_U10 (.A1( u1_u13_u1_n131 ) , .ZN( u1_u13_u1_n147 ) , .A2( u1_u13_u1_n153 ) );
  NAND3_X1 u1_u13_u1_U100 (.ZN( u1_u13_u1_n113 ) , .A1( u1_u13_u1_n120 ) , .A3( u1_u13_u1_n133 ) , .A2( u1_u13_u1_n155 ) );
  AOI22_X1 u1_u13_u1_U11 (.B2( u1_u13_u1_n136 ) , .A2( u1_u13_u1_n137 ) , .ZN( u1_u13_u1_n143 ) , .A1( u1_u13_u1_n171 ) , .B1( u1_u13_u1_n173 ) );
  INV_X1 u1_u13_u1_U12 (.A( u1_u13_u1_n147 ) , .ZN( u1_u13_u1_n181 ) );
  INV_X1 u1_u13_u1_U13 (.A( u1_u13_u1_n139 ) , .ZN( u1_u13_u1_n174 ) );
  OR4_X1 u1_u13_u1_U14 (.A4( u1_u13_u1_n106 ) , .A3( u1_u13_u1_n107 ) , .ZN( u1_u13_u1_n108 ) , .A1( u1_u13_u1_n117 ) , .A2( u1_u13_u1_n184 ) );
  AOI21_X1 u1_u13_u1_U15 (.ZN( u1_u13_u1_n106 ) , .A( u1_u13_u1_n112 ) , .B1( u1_u13_u1_n154 ) , .B2( u1_u13_u1_n156 ) );
  AOI21_X1 u1_u13_u1_U16 (.ZN( u1_u13_u1_n107 ) , .B1( u1_u13_u1_n134 ) , .B2( u1_u13_u1_n149 ) , .A( u1_u13_u1_n174 ) );
  INV_X1 u1_u13_u1_U17 (.A( u1_u13_u1_n101 ) , .ZN( u1_u13_u1_n184 ) );
  INV_X1 u1_u13_u1_U18 (.A( u1_u13_u1_n112 ) , .ZN( u1_u13_u1_n171 ) );
  NAND2_X1 u1_u13_u1_U19 (.ZN( u1_u13_u1_n141 ) , .A1( u1_u13_u1_n153 ) , .A2( u1_u13_u1_n156 ) );
  AND2_X1 u1_u13_u1_U20 (.A1( u1_u13_u1_n123 ) , .ZN( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n161 ) );
  NAND2_X1 u1_u13_u1_U21 (.A2( u1_u13_u1_n115 ) , .A1( u1_u13_u1_n116 ) , .ZN( u1_u13_u1_n148 ) );
  NAND2_X1 u1_u13_u1_U22 (.A2( u1_u13_u1_n133 ) , .A1( u1_u13_u1_n135 ) , .ZN( u1_u13_u1_n159 ) );
  NAND2_X1 u1_u13_u1_U23 (.A2( u1_u13_u1_n115 ) , .A1( u1_u13_u1_n120 ) , .ZN( u1_u13_u1_n132 ) );
  INV_X1 u1_u13_u1_U24 (.A( u1_u13_u1_n154 ) , .ZN( u1_u13_u1_n178 ) );
  AOI22_X1 u1_u13_u1_U25 (.B2( u1_u13_u1_n113 ) , .A2( u1_u13_u1_n114 ) , .ZN( u1_u13_u1_n125 ) , .A1( u1_u13_u1_n171 ) , .B1( u1_u13_u1_n173 ) );
  NAND2_X1 u1_u13_u1_U26 (.ZN( u1_u13_u1_n114 ) , .A1( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n156 ) );
  INV_X1 u1_u13_u1_U27 (.A( u1_u13_u1_n151 ) , .ZN( u1_u13_u1_n183 ) );
  AND2_X1 u1_u13_u1_U28 (.A1( u1_u13_u1_n129 ) , .A2( u1_u13_u1_n133 ) , .ZN( u1_u13_u1_n149 ) );
  INV_X1 u1_u13_u1_U29 (.A( u1_u13_u1_n131 ) , .ZN( u1_u13_u1_n180 ) );
  INV_X1 u1_u13_u1_U3 (.A( u1_u13_u1_n159 ) , .ZN( u1_u13_u1_n182 ) );
  OAI221_X1 u1_u13_u1_U30 (.A( u1_u13_u1_n119 ) , .C2( u1_u13_u1_n129 ) , .ZN( u1_u13_u1_n138 ) , .B2( u1_u13_u1_n152 ) , .C1( u1_u13_u1_n174 ) , .B1( u1_u13_u1_n187 ) );
  INV_X1 u1_u13_u1_U31 (.A( u1_u13_u1_n148 ) , .ZN( u1_u13_u1_n187 ) );
  AOI211_X1 u1_u13_u1_U32 (.B( u1_u13_u1_n117 ) , .A( u1_u13_u1_n118 ) , .ZN( u1_u13_u1_n119 ) , .C2( u1_u13_u1_n146 ) , .C1( u1_u13_u1_n159 ) );
  NOR2_X1 u1_u13_u1_U33 (.A1( u1_u13_u1_n168 ) , .A2( u1_u13_u1_n176 ) , .ZN( u1_u13_u1_n98 ) );
  AOI211_X1 u1_u13_u1_U34 (.B( u1_u13_u1_n162 ) , .A( u1_u13_u1_n163 ) , .C2( u1_u13_u1_n164 ) , .ZN( u1_u13_u1_n165 ) , .C1( u1_u13_u1_n171 ) );
  AOI21_X1 u1_u13_u1_U35 (.A( u1_u13_u1_n160 ) , .B2( u1_u13_u1_n161 ) , .ZN( u1_u13_u1_n162 ) , .B1( u1_u13_u1_n182 ) );
  OR2_X1 u1_u13_u1_U36 (.A2( u1_u13_u1_n157 ) , .A1( u1_u13_u1_n158 ) , .ZN( u1_u13_u1_n163 ) );
  OAI21_X1 u1_u13_u1_U37 (.B2( u1_u13_u1_n123 ) , .ZN( u1_u13_u1_n145 ) , .B1( u1_u13_u1_n160 ) , .A( u1_u13_u1_n185 ) );
  INV_X1 u1_u13_u1_U38 (.A( u1_u13_u1_n122 ) , .ZN( u1_u13_u1_n185 ) );
  AOI21_X1 u1_u13_u1_U39 (.B2( u1_u13_u1_n120 ) , .B1( u1_u13_u1_n121 ) , .ZN( u1_u13_u1_n122 ) , .A( u1_u13_u1_n128 ) );
  AOI221_X1 u1_u13_u1_U4 (.A( u1_u13_u1_n138 ) , .C2( u1_u13_u1_n139 ) , .C1( u1_u13_u1_n140 ) , .B2( u1_u13_u1_n141 ) , .ZN( u1_u13_u1_n142 ) , .B1( u1_u13_u1_n175 ) );
  NAND2_X1 u1_u13_u1_U40 (.A1( u1_u13_u1_n128 ) , .ZN( u1_u13_u1_n146 ) , .A2( u1_u13_u1_n160 ) );
  NAND2_X1 u1_u13_u1_U41 (.A2( u1_u13_u1_n112 ) , .ZN( u1_u13_u1_n139 ) , .A1( u1_u13_u1_n152 ) );
  NAND2_X1 u1_u13_u1_U42 (.A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n156 ) , .A2( u1_u13_u1_n99 ) );
  AOI221_X1 u1_u13_u1_U43 (.B1( u1_u13_u1_n140 ) , .ZN( u1_u13_u1_n167 ) , .B2( u1_u13_u1_n172 ) , .C2( u1_u13_u1_n175 ) , .C1( u1_u13_u1_n178 ) , .A( u1_u13_u1_n188 ) );
  INV_X1 u1_u13_u1_U44 (.ZN( u1_u13_u1_n188 ) , .A( u1_u13_u1_n97 ) );
  AOI211_X1 u1_u13_u1_U45 (.A( u1_u13_u1_n118 ) , .C1( u1_u13_u1_n132 ) , .C2( u1_u13_u1_n139 ) , .B( u1_u13_u1_n96 ) , .ZN( u1_u13_u1_n97 ) );
  AOI21_X1 u1_u13_u1_U46 (.B2( u1_u13_u1_n121 ) , .B1( u1_u13_u1_n135 ) , .A( u1_u13_u1_n152 ) , .ZN( u1_u13_u1_n96 ) );
  NOR2_X1 u1_u13_u1_U47 (.ZN( u1_u13_u1_n117 ) , .A1( u1_u13_u1_n121 ) , .A2( u1_u13_u1_n160 ) );
  AOI21_X1 u1_u13_u1_U48 (.A( u1_u13_u1_n128 ) , .B2( u1_u13_u1_n129 ) , .ZN( u1_u13_u1_n130 ) , .B1( u1_u13_u1_n150 ) );
  NAND2_X1 u1_u13_u1_U49 (.ZN( u1_u13_u1_n112 ) , .A1( u1_u13_u1_n169 ) , .A2( u1_u13_u1_n170 ) );
  AOI211_X1 u1_u13_u1_U5 (.ZN( u1_u13_u1_n124 ) , .A( u1_u13_u1_n138 ) , .C2( u1_u13_u1_n139 ) , .B( u1_u13_u1_n145 ) , .C1( u1_u13_u1_n147 ) );
  NAND2_X1 u1_u13_u1_U50 (.ZN( u1_u13_u1_n129 ) , .A2( u1_u13_u1_n95 ) , .A1( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U51 (.A1( u1_u13_u1_n102 ) , .ZN( u1_u13_u1_n154 ) , .A2( u1_u13_u1_n99 ) );
  NAND2_X1 u1_u13_u1_U52 (.A2( u1_u13_u1_n100 ) , .ZN( u1_u13_u1_n135 ) , .A1( u1_u13_u1_n99 ) );
  AOI21_X1 u1_u13_u1_U53 (.A( u1_u13_u1_n152 ) , .B2( u1_u13_u1_n153 ) , .B1( u1_u13_u1_n154 ) , .ZN( u1_u13_u1_n158 ) );
  INV_X1 u1_u13_u1_U54 (.A( u1_u13_u1_n160 ) , .ZN( u1_u13_u1_n175 ) );
  NAND2_X1 u1_u13_u1_U55 (.A1( u1_u13_u1_n100 ) , .ZN( u1_u13_u1_n116 ) , .A2( u1_u13_u1_n95 ) );
  NAND2_X1 u1_u13_u1_U56 (.A1( u1_u13_u1_n102 ) , .ZN( u1_u13_u1_n131 ) , .A2( u1_u13_u1_n95 ) );
  NAND2_X1 u1_u13_u1_U57 (.A2( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n121 ) , .A1( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U58 (.A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n153 ) , .A2( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U59 (.A2( u1_u13_u1_n104 ) , .A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n133 ) );
  NOR2_X1 u1_u13_u1_U6 (.A1( u1_u13_u1_n112 ) , .A2( u1_u13_u1_n116 ) , .ZN( u1_u13_u1_n118 ) );
  NAND2_X1 u1_u13_u1_U60 (.ZN( u1_u13_u1_n150 ) , .A2( u1_u13_u1_n98 ) , .A1( u1_u13_u1_n99 ) );
  NAND2_X1 u1_u13_u1_U61 (.A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n155 ) , .A2( u1_u13_u1_n95 ) );
  OAI21_X1 u1_u13_u1_U62 (.ZN( u1_u13_u1_n109 ) , .B1( u1_u13_u1_n129 ) , .B2( u1_u13_u1_n160 ) , .A( u1_u13_u1_n167 ) );
  NAND2_X1 u1_u13_u1_U63 (.A2( u1_u13_u1_n100 ) , .A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n120 ) );
  NAND2_X1 u1_u13_u1_U64 (.A1( u1_u13_u1_n102 ) , .A2( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n115 ) );
  NAND2_X1 u1_u13_u1_U65 (.A2( u1_u13_u1_n100 ) , .A1( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n151 ) );
  NAND2_X1 u1_u13_u1_U66 (.A2( u1_u13_u1_n103 ) , .A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n161 ) );
  INV_X1 u1_u13_u1_U67 (.A( u1_u13_u1_n152 ) , .ZN( u1_u13_u1_n173 ) );
  INV_X1 u1_u13_u1_U68 (.A( u1_u13_u1_n128 ) , .ZN( u1_u13_u1_n172 ) );
  NAND2_X1 u1_u13_u1_U69 (.A2( u1_u13_u1_n102 ) , .A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n123 ) );
  OAI21_X1 u1_u13_u1_U7 (.ZN( u1_u13_u1_n101 ) , .B1( u1_u13_u1_n141 ) , .A( u1_u13_u1_n146 ) , .B2( u1_u13_u1_n183 ) );
  NOR2_X1 u1_u13_u1_U70 (.A2( u1_u13_X_7 ) , .A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n95 ) );
  NOR2_X1 u1_u13_u1_U71 (.A1( u1_u13_X_12 ) , .A2( u1_u13_X_9 ) , .ZN( u1_u13_u1_n100 ) );
  NOR2_X1 u1_u13_u1_U72 (.A2( u1_u13_X_8 ) , .A1( u1_u13_u1_n177 ) , .ZN( u1_u13_u1_n99 ) );
  NOR2_X1 u1_u13_u1_U73 (.A2( u1_u13_X_12 ) , .ZN( u1_u13_u1_n102 ) , .A1( u1_u13_u1_n176 ) );
  NOR2_X1 u1_u13_u1_U74 (.A2( u1_u13_X_9 ) , .ZN( u1_u13_u1_n105 ) , .A1( u1_u13_u1_n168 ) );
  NAND2_X1 u1_u13_u1_U75 (.A1( u1_u13_X_10 ) , .ZN( u1_u13_u1_n160 ) , .A2( u1_u13_u1_n169 ) );
  NAND2_X1 u1_u13_u1_U76 (.A2( u1_u13_X_10 ) , .A1( u1_u13_X_11 ) , .ZN( u1_u13_u1_n152 ) );
  NAND2_X1 u1_u13_u1_U77 (.A1( u1_u13_X_11 ) , .ZN( u1_u13_u1_n128 ) , .A2( u1_u13_u1_n170 ) );
  AND2_X1 u1_u13_u1_U78 (.A2( u1_u13_X_7 ) , .A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n104 ) );
  AND2_X1 u1_u13_u1_U79 (.A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n103 ) , .A2( u1_u13_u1_n177 ) );
  AOI21_X1 u1_u13_u1_U8 (.B2( u1_u13_u1_n155 ) , .B1( u1_u13_u1_n156 ) , .ZN( u1_u13_u1_n157 ) , .A( u1_u13_u1_n174 ) );
  INV_X1 u1_u13_u1_U80 (.A( u1_u13_X_10 ) , .ZN( u1_u13_u1_n170 ) );
  INV_X1 u1_u13_u1_U81 (.A( u1_u13_X_9 ) , .ZN( u1_u13_u1_n176 ) );
  INV_X1 u1_u13_u1_U82 (.A( u1_u13_X_11 ) , .ZN( u1_u13_u1_n169 ) );
  INV_X1 u1_u13_u1_U83 (.A( u1_u13_X_12 ) , .ZN( u1_u13_u1_n168 ) );
  INV_X1 u1_u13_u1_U84 (.A( u1_u13_X_7 ) , .ZN( u1_u13_u1_n177 ) );
  NAND4_X1 u1_u13_u1_U85 (.ZN( u1_out13_18 ) , .A4( u1_u13_u1_n165 ) , .A3( u1_u13_u1_n166 ) , .A1( u1_u13_u1_n167 ) , .A2( u1_u13_u1_n186 ) );
  AOI22_X1 u1_u13_u1_U86 (.B2( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n147 ) , .A2( u1_u13_u1_n148 ) , .ZN( u1_u13_u1_n166 ) , .A1( u1_u13_u1_n172 ) );
  INV_X1 u1_u13_u1_U87 (.A( u1_u13_u1_n145 ) , .ZN( u1_u13_u1_n186 ) );
  NAND4_X1 u1_u13_u1_U88 (.ZN( u1_out13_2 ) , .A4( u1_u13_u1_n142 ) , .A3( u1_u13_u1_n143 ) , .A2( u1_u13_u1_n144 ) , .A1( u1_u13_u1_n179 ) );
  OAI21_X1 u1_u13_u1_U89 (.B2( u1_u13_u1_n132 ) , .ZN( u1_u13_u1_n144 ) , .A( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n180 ) );
  NAND2_X1 u1_u13_u1_U9 (.ZN( u1_u13_u1_n140 ) , .A2( u1_u13_u1_n150 ) , .A1( u1_u13_u1_n155 ) );
  INV_X1 u1_u13_u1_U90 (.A( u1_u13_u1_n130 ) , .ZN( u1_u13_u1_n179 ) );
  NAND4_X1 u1_u13_u1_U91 (.ZN( u1_out13_28 ) , .A4( u1_u13_u1_n124 ) , .A3( u1_u13_u1_n125 ) , .A2( u1_u13_u1_n126 ) , .A1( u1_u13_u1_n127 ) );
  OAI21_X1 u1_u13_u1_U92 (.ZN( u1_u13_u1_n127 ) , .B2( u1_u13_u1_n139 ) , .B1( u1_u13_u1_n175 ) , .A( u1_u13_u1_n183 ) );
  OAI21_X1 u1_u13_u1_U93 (.ZN( u1_u13_u1_n126 ) , .B2( u1_u13_u1_n140 ) , .A( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n178 ) );
  OR4_X1 u1_u13_u1_U94 (.ZN( u1_out13_13 ) , .A4( u1_u13_u1_n108 ) , .A3( u1_u13_u1_n109 ) , .A2( u1_u13_u1_n110 ) , .A1( u1_u13_u1_n111 ) );
  AOI21_X1 u1_u13_u1_U95 (.ZN( u1_u13_u1_n111 ) , .A( u1_u13_u1_n128 ) , .B2( u1_u13_u1_n131 ) , .B1( u1_u13_u1_n135 ) );
  AOI21_X1 u1_u13_u1_U96 (.ZN( u1_u13_u1_n110 ) , .A( u1_u13_u1_n116 ) , .B1( u1_u13_u1_n152 ) , .B2( u1_u13_u1_n160 ) );
  NAND3_X1 u1_u13_u1_U97 (.A3( u1_u13_u1_n149 ) , .A2( u1_u13_u1_n150 ) , .A1( u1_u13_u1_n151 ) , .ZN( u1_u13_u1_n164 ) );
  NAND3_X1 u1_u13_u1_U98 (.A3( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n135 ) , .ZN( u1_u13_u1_n136 ) , .A1( u1_u13_u1_n151 ) );
  NAND3_X1 u1_u13_u1_U99 (.A1( u1_u13_u1_n133 ) , .ZN( u1_u13_u1_n137 ) , .A2( u1_u13_u1_n154 ) , .A3( u1_u13_u1_n181 ) );
  AOI22_X1 u1_u13_u6_U10 (.A2( u1_u13_u6_n151 ) , .B2( u1_u13_u6_n161 ) , .A1( u1_u13_u6_n167 ) , .B1( u1_u13_u6_n170 ) , .ZN( u1_u13_u6_n89 ) );
  AOI21_X1 u1_u13_u6_U11 (.B1( u1_u13_u6_n107 ) , .B2( u1_u13_u6_n132 ) , .A( u1_u13_u6_n158 ) , .ZN( u1_u13_u6_n88 ) );
  AOI21_X1 u1_u13_u6_U12 (.B2( u1_u13_u6_n147 ) , .B1( u1_u13_u6_n148 ) , .ZN( u1_u13_u6_n149 ) , .A( u1_u13_u6_n158 ) );
  AOI21_X1 u1_u13_u6_U13 (.ZN( u1_u13_u6_n106 ) , .A( u1_u13_u6_n142 ) , .B2( u1_u13_u6_n159 ) , .B1( u1_u13_u6_n164 ) );
  INV_X1 u1_u13_u6_U14 (.A( u1_u13_u6_n155 ) , .ZN( u1_u13_u6_n161 ) );
  INV_X1 u1_u13_u6_U15 (.A( u1_u13_u6_n128 ) , .ZN( u1_u13_u6_n164 ) );
  NAND2_X1 u1_u13_u6_U16 (.ZN( u1_u13_u6_n110 ) , .A1( u1_u13_u6_n122 ) , .A2( u1_u13_u6_n129 ) );
  NAND2_X1 u1_u13_u6_U17 (.ZN( u1_u13_u6_n124 ) , .A2( u1_u13_u6_n146 ) , .A1( u1_u13_u6_n148 ) );
  INV_X1 u1_u13_u6_U18 (.A( u1_u13_u6_n132 ) , .ZN( u1_u13_u6_n171 ) );
  AND2_X1 u1_u13_u6_U19 (.A1( u1_u13_u6_n100 ) , .ZN( u1_u13_u6_n130 ) , .A2( u1_u13_u6_n147 ) );
  INV_X1 u1_u13_u6_U20 (.A( u1_u13_u6_n127 ) , .ZN( u1_u13_u6_n173 ) );
  INV_X1 u1_u13_u6_U21 (.A( u1_u13_u6_n121 ) , .ZN( u1_u13_u6_n167 ) );
  INV_X1 u1_u13_u6_U22 (.A( u1_u13_u6_n100 ) , .ZN( u1_u13_u6_n169 ) );
  INV_X1 u1_u13_u6_U23 (.A( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n170 ) );
  INV_X1 u1_u13_u6_U24 (.A( u1_u13_u6_n113 ) , .ZN( u1_u13_u6_n168 ) );
  AND2_X1 u1_u13_u6_U25 (.A1( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n119 ) , .ZN( u1_u13_u6_n133 ) );
  AND2_X1 u1_u13_u6_U26 (.A2( u1_u13_u6_n121 ) , .A1( u1_u13_u6_n122 ) , .ZN( u1_u13_u6_n131 ) );
  AND3_X1 u1_u13_u6_U27 (.ZN( u1_u13_u6_n120 ) , .A2( u1_u13_u6_n127 ) , .A1( u1_u13_u6_n132 ) , .A3( u1_u13_u6_n145 ) );
  INV_X1 u1_u13_u6_U28 (.A( u1_u13_u6_n146 ) , .ZN( u1_u13_u6_n163 ) );
  AOI222_X1 u1_u13_u6_U29 (.ZN( u1_u13_u6_n114 ) , .A1( u1_u13_u6_n118 ) , .A2( u1_u13_u6_n126 ) , .B2( u1_u13_u6_n151 ) , .C2( u1_u13_u6_n159 ) , .C1( u1_u13_u6_n168 ) , .B1( u1_u13_u6_n169 ) );
  INV_X1 u1_u13_u6_U3 (.A( u1_u13_u6_n110 ) , .ZN( u1_u13_u6_n166 ) );
  NOR2_X1 u1_u13_u6_U30 (.A1( u1_u13_u6_n162 ) , .A2( u1_u13_u6_n165 ) , .ZN( u1_u13_u6_n98 ) );
  AOI211_X1 u1_u13_u6_U31 (.B( u1_u13_u6_n134 ) , .A( u1_u13_u6_n135 ) , .C1( u1_u13_u6_n136 ) , .ZN( u1_u13_u6_n137 ) , .C2( u1_u13_u6_n151 ) );
  AOI21_X1 u1_u13_u6_U32 (.B2( u1_u13_u6_n132 ) , .B1( u1_u13_u6_n133 ) , .ZN( u1_u13_u6_n134 ) , .A( u1_u13_u6_n158 ) );
  AOI21_X1 u1_u13_u6_U33 (.B1( u1_u13_u6_n131 ) , .ZN( u1_u13_u6_n135 ) , .A( u1_u13_u6_n144 ) , .B2( u1_u13_u6_n146 ) );
  NAND4_X1 u1_u13_u6_U34 (.A4( u1_u13_u6_n127 ) , .A3( u1_u13_u6_n128 ) , .A2( u1_u13_u6_n129 ) , .A1( u1_u13_u6_n130 ) , .ZN( u1_u13_u6_n136 ) );
  NAND2_X1 u1_u13_u6_U35 (.A1( u1_u13_u6_n144 ) , .ZN( u1_u13_u6_n151 ) , .A2( u1_u13_u6_n158 ) );
  NAND2_X1 u1_u13_u6_U36 (.ZN( u1_u13_u6_n132 ) , .A1( u1_u13_u6_n91 ) , .A2( u1_u13_u6_n97 ) );
  AOI22_X1 u1_u13_u6_U37 (.B2( u1_u13_u6_n110 ) , .B1( u1_u13_u6_n111 ) , .A1( u1_u13_u6_n112 ) , .ZN( u1_u13_u6_n115 ) , .A2( u1_u13_u6_n161 ) );
  NAND4_X1 u1_u13_u6_U38 (.A3( u1_u13_u6_n109 ) , .ZN( u1_u13_u6_n112 ) , .A4( u1_u13_u6_n132 ) , .A2( u1_u13_u6_n147 ) , .A1( u1_u13_u6_n166 ) );
  NOR2_X1 u1_u13_u6_U39 (.ZN( u1_u13_u6_n109 ) , .A1( u1_u13_u6_n170 ) , .A2( u1_u13_u6_n173 ) );
  INV_X1 u1_u13_u6_U4 (.A( u1_u13_u6_n142 ) , .ZN( u1_u13_u6_n174 ) );
  NOR2_X1 u1_u13_u6_U40 (.A2( u1_u13_u6_n126 ) , .ZN( u1_u13_u6_n155 ) , .A1( u1_u13_u6_n160 ) );
  NAND2_X1 u1_u13_u6_U41 (.ZN( u1_u13_u6_n146 ) , .A2( u1_u13_u6_n94 ) , .A1( u1_u13_u6_n99 ) );
  AOI21_X1 u1_u13_u6_U42 (.A( u1_u13_u6_n144 ) , .B2( u1_u13_u6_n145 ) , .B1( u1_u13_u6_n146 ) , .ZN( u1_u13_u6_n150 ) );
  INV_X1 u1_u13_u6_U43 (.A( u1_u13_u6_n111 ) , .ZN( u1_u13_u6_n158 ) );
  NAND2_X1 u1_u13_u6_U44 (.ZN( u1_u13_u6_n127 ) , .A1( u1_u13_u6_n91 ) , .A2( u1_u13_u6_n92 ) );
  NAND2_X1 u1_u13_u6_U45 (.ZN( u1_u13_u6_n129 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n96 ) );
  INV_X1 u1_u13_u6_U46 (.A( u1_u13_u6_n144 ) , .ZN( u1_u13_u6_n159 ) );
  NAND2_X1 u1_u13_u6_U47 (.ZN( u1_u13_u6_n145 ) , .A2( u1_u13_u6_n97 ) , .A1( u1_u13_u6_n98 ) );
  NAND2_X1 u1_u13_u6_U48 (.ZN( u1_u13_u6_n148 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n94 ) );
  NAND2_X1 u1_u13_u6_U49 (.ZN( u1_u13_u6_n108 ) , .A2( u1_u13_u6_n139 ) , .A1( u1_u13_u6_n144 ) );
  NAND2_X1 u1_u13_u6_U5 (.A2( u1_u13_u6_n143 ) , .ZN( u1_u13_u6_n152 ) , .A1( u1_u13_u6_n166 ) );
  NAND2_X1 u1_u13_u6_U50 (.ZN( u1_u13_u6_n121 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n97 ) );
  NAND2_X1 u1_u13_u6_U51 (.ZN( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n95 ) );
  AND2_X1 u1_u13_u6_U52 (.ZN( u1_u13_u6_n118 ) , .A2( u1_u13_u6_n91 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U53 (.ZN( u1_u13_u6_n147 ) , .A2( u1_u13_u6_n98 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U54 (.ZN( u1_u13_u6_n128 ) , .A1( u1_u13_u6_n94 ) , .A2( u1_u13_u6_n96 ) );
  NAND2_X1 u1_u13_u6_U55 (.ZN( u1_u13_u6_n119 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U56 (.ZN( u1_u13_u6_n123 ) , .A2( u1_u13_u6_n91 ) , .A1( u1_u13_u6_n96 ) );
  NAND2_X1 u1_u13_u6_U57 (.ZN( u1_u13_u6_n100 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n98 ) );
  NAND2_X1 u1_u13_u6_U58 (.ZN( u1_u13_u6_n122 ) , .A1( u1_u13_u6_n94 ) , .A2( u1_u13_u6_n97 ) );
  INV_X1 u1_u13_u6_U59 (.A( u1_u13_u6_n139 ) , .ZN( u1_u13_u6_n160 ) );
  AOI22_X1 u1_u13_u6_U6 (.B2( u1_u13_u6_n101 ) , .A1( u1_u13_u6_n102 ) , .ZN( u1_u13_u6_n103 ) , .B1( u1_u13_u6_n160 ) , .A2( u1_u13_u6_n161 ) );
  NAND2_X1 u1_u13_u6_U60 (.ZN( u1_u13_u6_n113 ) , .A1( u1_u13_u6_n96 ) , .A2( u1_u13_u6_n98 ) );
  NOR2_X1 u1_u13_u6_U61 (.A2( u1_u13_X_40 ) , .A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n126 ) );
  NOR2_X1 u1_u13_u6_U62 (.A2( u1_u13_X_39 ) , .A1( u1_u13_X_42 ) , .ZN( u1_u13_u6_n92 ) );
  NOR2_X1 u1_u13_u6_U63 (.A2( u1_u13_X_39 ) , .A1( u1_u13_u6_n156 ) , .ZN( u1_u13_u6_n97 ) );
  NOR2_X1 u1_u13_u6_U64 (.A2( u1_u13_X_38 ) , .A1( u1_u13_u6_n165 ) , .ZN( u1_u13_u6_n95 ) );
  NOR2_X1 u1_u13_u6_U65 (.A2( u1_u13_X_41 ) , .ZN( u1_u13_u6_n111 ) , .A1( u1_u13_u6_n157 ) );
  NOR2_X1 u1_u13_u6_U66 (.A2( u1_u13_X_37 ) , .A1( u1_u13_u6_n162 ) , .ZN( u1_u13_u6_n94 ) );
  NOR2_X1 u1_u13_u6_U67 (.A2( u1_u13_X_37 ) , .A1( u1_u13_X_38 ) , .ZN( u1_u13_u6_n91 ) );
  NAND2_X1 u1_u13_u6_U68 (.A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n144 ) , .A2( u1_u13_u6_n157 ) );
  NAND2_X1 u1_u13_u6_U69 (.A2( u1_u13_X_40 ) , .A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n139 ) );
  NOR2_X1 u1_u13_u6_U7 (.A1( u1_u13_u6_n118 ) , .ZN( u1_u13_u6_n143 ) , .A2( u1_u13_u6_n168 ) );
  AND2_X1 u1_u13_u6_U70 (.A1( u1_u13_X_39 ) , .A2( u1_u13_u6_n156 ) , .ZN( u1_u13_u6_n96 ) );
  AND2_X1 u1_u13_u6_U71 (.A1( u1_u13_X_39 ) , .A2( u1_u13_X_42 ) , .ZN( u1_u13_u6_n99 ) );
  INV_X1 u1_u13_u6_U72 (.A( u1_u13_X_40 ) , .ZN( u1_u13_u6_n157 ) );
  INV_X1 u1_u13_u6_U73 (.A( u1_u13_X_37 ) , .ZN( u1_u13_u6_n165 ) );
  INV_X1 u1_u13_u6_U74 (.A( u1_u13_X_38 ) , .ZN( u1_u13_u6_n162 ) );
  INV_X1 u1_u13_u6_U75 (.A( u1_u13_X_42 ) , .ZN( u1_u13_u6_n156 ) );
  NAND4_X1 u1_u13_u6_U76 (.ZN( u1_out13_32 ) , .A4( u1_u13_u6_n103 ) , .A3( u1_u13_u6_n104 ) , .A2( u1_u13_u6_n105 ) , .A1( u1_u13_u6_n106 ) );
  AOI22_X1 u1_u13_u6_U77 (.ZN( u1_u13_u6_n105 ) , .A2( u1_u13_u6_n108 ) , .A1( u1_u13_u6_n118 ) , .B2( u1_u13_u6_n126 ) , .B1( u1_u13_u6_n171 ) );
  AOI22_X1 u1_u13_u6_U78 (.ZN( u1_u13_u6_n104 ) , .A1( u1_u13_u6_n111 ) , .B1( u1_u13_u6_n124 ) , .B2( u1_u13_u6_n151 ) , .A2( u1_u13_u6_n93 ) );
  NAND4_X1 u1_u13_u6_U79 (.ZN( u1_out13_12 ) , .A4( u1_u13_u6_n114 ) , .A3( u1_u13_u6_n115 ) , .A2( u1_u13_u6_n116 ) , .A1( u1_u13_u6_n117 ) );
  OAI21_X1 u1_u13_u6_U8 (.A( u1_u13_u6_n159 ) , .B1( u1_u13_u6_n169 ) , .B2( u1_u13_u6_n173 ) , .ZN( u1_u13_u6_n90 ) );
  OAI22_X1 u1_u13_u6_U80 (.B2( u1_u13_u6_n111 ) , .ZN( u1_u13_u6_n116 ) , .B1( u1_u13_u6_n126 ) , .A2( u1_u13_u6_n164 ) , .A1( u1_u13_u6_n167 ) );
  OAI21_X1 u1_u13_u6_U81 (.A( u1_u13_u6_n108 ) , .ZN( u1_u13_u6_n117 ) , .B2( u1_u13_u6_n141 ) , .B1( u1_u13_u6_n163 ) );
  OAI211_X1 u1_u13_u6_U82 (.ZN( u1_out13_7 ) , .B( u1_u13_u6_n153 ) , .C2( u1_u13_u6_n154 ) , .C1( u1_u13_u6_n155 ) , .A( u1_u13_u6_n174 ) );
  NOR3_X1 u1_u13_u6_U83 (.A1( u1_u13_u6_n141 ) , .ZN( u1_u13_u6_n154 ) , .A3( u1_u13_u6_n164 ) , .A2( u1_u13_u6_n171 ) );
  AOI211_X1 u1_u13_u6_U84 (.B( u1_u13_u6_n149 ) , .A( u1_u13_u6_n150 ) , .C2( u1_u13_u6_n151 ) , .C1( u1_u13_u6_n152 ) , .ZN( u1_u13_u6_n153 ) );
  OAI211_X1 u1_u13_u6_U85 (.ZN( u1_out13_22 ) , .B( u1_u13_u6_n137 ) , .A( u1_u13_u6_n138 ) , .C2( u1_u13_u6_n139 ) , .C1( u1_u13_u6_n140 ) );
  AOI22_X1 u1_u13_u6_U86 (.B1( u1_u13_u6_n124 ) , .A2( u1_u13_u6_n125 ) , .A1( u1_u13_u6_n126 ) , .ZN( u1_u13_u6_n138 ) , .B2( u1_u13_u6_n161 ) );
  AND4_X1 u1_u13_u6_U87 (.A3( u1_u13_u6_n119 ) , .A1( u1_u13_u6_n120 ) , .A4( u1_u13_u6_n129 ) , .ZN( u1_u13_u6_n140 ) , .A2( u1_u13_u6_n143 ) );
  NAND3_X1 u1_u13_u6_U88 (.A2( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n125 ) , .A1( u1_u13_u6_n130 ) , .A3( u1_u13_u6_n131 ) );
  NAND3_X1 u1_u13_u6_U89 (.A3( u1_u13_u6_n133 ) , .ZN( u1_u13_u6_n141 ) , .A1( u1_u13_u6_n145 ) , .A2( u1_u13_u6_n148 ) );
  INV_X1 u1_u13_u6_U9 (.ZN( u1_u13_u6_n172 ) , .A( u1_u13_u6_n88 ) );
  NAND3_X1 u1_u13_u6_U90 (.ZN( u1_u13_u6_n101 ) , .A3( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n121 ) , .A1( u1_u13_u6_n127 ) );
  NAND3_X1 u1_u13_u6_U91 (.ZN( u1_u13_u6_n102 ) , .A3( u1_u13_u6_n130 ) , .A2( u1_u13_u6_n145 ) , .A1( u1_u13_u6_n166 ) );
  NAND3_X1 u1_u13_u6_U92 (.A3( u1_u13_u6_n113 ) , .A1( u1_u13_u6_n119 ) , .A2( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n93 ) );
  NAND3_X1 u1_u13_u6_U93 (.ZN( u1_u13_u6_n142 ) , .A2( u1_u13_u6_n172 ) , .A3( u1_u13_u6_n89 ) , .A1( u1_u13_u6_n90 ) );
  AND3_X1 u1_u13_u7_U10 (.A3( u1_u13_u7_n110 ) , .A2( u1_u13_u7_n127 ) , .A1( u1_u13_u7_n132 ) , .ZN( u1_u13_u7_n92 ) );
  OAI21_X1 u1_u13_u7_U11 (.A( u1_u13_u7_n161 ) , .B1( u1_u13_u7_n168 ) , .B2( u1_u13_u7_n173 ) , .ZN( u1_u13_u7_n91 ) );
  AOI211_X1 u1_u13_u7_U12 (.A( u1_u13_u7_n117 ) , .ZN( u1_u13_u7_n118 ) , .C2( u1_u13_u7_n126 ) , .C1( u1_u13_u7_n177 ) , .B( u1_u13_u7_n180 ) );
  OAI22_X1 u1_u13_u7_U13 (.B1( u1_u13_u7_n115 ) , .ZN( u1_u13_u7_n117 ) , .A2( u1_u13_u7_n133 ) , .A1( u1_u13_u7_n137 ) , .B2( u1_u13_u7_n162 ) );
  INV_X1 u1_u13_u7_U14 (.A( u1_u13_u7_n116 ) , .ZN( u1_u13_u7_n180 ) );
  NOR3_X1 u1_u13_u7_U15 (.ZN( u1_u13_u7_n115 ) , .A3( u1_u13_u7_n145 ) , .A2( u1_u13_u7_n168 ) , .A1( u1_u13_u7_n169 ) );
  OAI211_X1 u1_u13_u7_U16 (.B( u1_u13_u7_n122 ) , .A( u1_u13_u7_n123 ) , .C2( u1_u13_u7_n124 ) , .ZN( u1_u13_u7_n154 ) , .C1( u1_u13_u7_n162 ) );
  AOI222_X1 u1_u13_u7_U17 (.ZN( u1_u13_u7_n122 ) , .C2( u1_u13_u7_n126 ) , .C1( u1_u13_u7_n145 ) , .B1( u1_u13_u7_n161 ) , .A2( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n170 ) , .A1( u1_u13_u7_n176 ) );
  INV_X1 u1_u13_u7_U18 (.A( u1_u13_u7_n133 ) , .ZN( u1_u13_u7_n176 ) );
  NOR3_X1 u1_u13_u7_U19 (.A2( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n135 ) , .ZN( u1_u13_u7_n136 ) , .A3( u1_u13_u7_n171 ) );
  NOR2_X1 u1_u13_u7_U20 (.A1( u1_u13_u7_n130 ) , .A2( u1_u13_u7_n134 ) , .ZN( u1_u13_u7_n153 ) );
  INV_X1 u1_u13_u7_U21 (.A( u1_u13_u7_n101 ) , .ZN( u1_u13_u7_n165 ) );
  NOR2_X1 u1_u13_u7_U22 (.ZN( u1_u13_u7_n111 ) , .A2( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n169 ) );
  AOI21_X1 u1_u13_u7_U23 (.ZN( u1_u13_u7_n104 ) , .B2( u1_u13_u7_n112 ) , .B1( u1_u13_u7_n127 ) , .A( u1_u13_u7_n164 ) );
  AOI21_X1 u1_u13_u7_U24 (.ZN( u1_u13_u7_n106 ) , .B1( u1_u13_u7_n133 ) , .B2( u1_u13_u7_n146 ) , .A( u1_u13_u7_n162 ) );
  AOI21_X1 u1_u13_u7_U25 (.A( u1_u13_u7_n101 ) , .ZN( u1_u13_u7_n107 ) , .B2( u1_u13_u7_n128 ) , .B1( u1_u13_u7_n175 ) );
  INV_X1 u1_u13_u7_U26 (.A( u1_u13_u7_n138 ) , .ZN( u1_u13_u7_n171 ) );
  INV_X1 u1_u13_u7_U27 (.A( u1_u13_u7_n131 ) , .ZN( u1_u13_u7_n177 ) );
  INV_X1 u1_u13_u7_U28 (.A( u1_u13_u7_n110 ) , .ZN( u1_u13_u7_n174 ) );
  NAND2_X1 u1_u13_u7_U29 (.A1( u1_u13_u7_n129 ) , .A2( u1_u13_u7_n132 ) , .ZN( u1_u13_u7_n149 ) );
  OAI21_X1 u1_u13_u7_U3 (.ZN( u1_u13_u7_n159 ) , .A( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n171 ) , .B1( u1_u13_u7_n174 ) );
  NAND2_X1 u1_u13_u7_U30 (.A1( u1_u13_u7_n113 ) , .A2( u1_u13_u7_n124 ) , .ZN( u1_u13_u7_n130 ) );
  INV_X1 u1_u13_u7_U31 (.A( u1_u13_u7_n112 ) , .ZN( u1_u13_u7_n173 ) );
  INV_X1 u1_u13_u7_U32 (.A( u1_u13_u7_n128 ) , .ZN( u1_u13_u7_n168 ) );
  INV_X1 u1_u13_u7_U33 (.A( u1_u13_u7_n148 ) , .ZN( u1_u13_u7_n169 ) );
  INV_X1 u1_u13_u7_U34 (.A( u1_u13_u7_n127 ) , .ZN( u1_u13_u7_n179 ) );
  NOR2_X1 u1_u13_u7_U35 (.ZN( u1_u13_u7_n101 ) , .A2( u1_u13_u7_n150 ) , .A1( u1_u13_u7_n156 ) );
  AOI211_X1 u1_u13_u7_U36 (.B( u1_u13_u7_n154 ) , .A( u1_u13_u7_n155 ) , .C1( u1_u13_u7_n156 ) , .ZN( u1_u13_u7_n157 ) , .C2( u1_u13_u7_n172 ) );
  INV_X1 u1_u13_u7_U37 (.A( u1_u13_u7_n153 ) , .ZN( u1_u13_u7_n172 ) );
  AOI211_X1 u1_u13_u7_U38 (.B( u1_u13_u7_n139 ) , .A( u1_u13_u7_n140 ) , .C2( u1_u13_u7_n141 ) , .ZN( u1_u13_u7_n142 ) , .C1( u1_u13_u7_n156 ) );
  NAND4_X1 u1_u13_u7_U39 (.A3( u1_u13_u7_n127 ) , .A2( u1_u13_u7_n128 ) , .A1( u1_u13_u7_n129 ) , .ZN( u1_u13_u7_n141 ) , .A4( u1_u13_u7_n147 ) );
  INV_X1 u1_u13_u7_U4 (.A( u1_u13_u7_n111 ) , .ZN( u1_u13_u7_n170 ) );
  AOI21_X1 u1_u13_u7_U40 (.A( u1_u13_u7_n137 ) , .B1( u1_u13_u7_n138 ) , .ZN( u1_u13_u7_n139 ) , .B2( u1_u13_u7_n146 ) );
  OAI22_X1 u1_u13_u7_U41 (.B1( u1_u13_u7_n136 ) , .ZN( u1_u13_u7_n140 ) , .A1( u1_u13_u7_n153 ) , .B2( u1_u13_u7_n162 ) , .A2( u1_u13_u7_n164 ) );
  AOI21_X1 u1_u13_u7_U42 (.ZN( u1_u13_u7_n123 ) , .B1( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n177 ) , .A( u1_u13_u7_n97 ) );
  AOI21_X1 u1_u13_u7_U43 (.B2( u1_u13_u7_n113 ) , .B1( u1_u13_u7_n124 ) , .A( u1_u13_u7_n125 ) , .ZN( u1_u13_u7_n97 ) );
  INV_X1 u1_u13_u7_U44 (.A( u1_u13_u7_n125 ) , .ZN( u1_u13_u7_n161 ) );
  INV_X1 u1_u13_u7_U45 (.A( u1_u13_u7_n152 ) , .ZN( u1_u13_u7_n162 ) );
  AOI22_X1 u1_u13_u7_U46 (.A2( u1_u13_u7_n114 ) , .ZN( u1_u13_u7_n119 ) , .B1( u1_u13_u7_n130 ) , .A1( u1_u13_u7_n156 ) , .B2( u1_u13_u7_n165 ) );
  NAND2_X1 u1_u13_u7_U47 (.A2( u1_u13_u7_n112 ) , .ZN( u1_u13_u7_n114 ) , .A1( u1_u13_u7_n175 ) );
  AND2_X1 u1_u13_u7_U48 (.ZN( u1_u13_u7_n145 ) , .A2( u1_u13_u7_n98 ) , .A1( u1_u13_u7_n99 ) );
  NOR2_X1 u1_u13_u7_U49 (.ZN( u1_u13_u7_n137 ) , .A1( u1_u13_u7_n150 ) , .A2( u1_u13_u7_n161 ) );
  INV_X1 u1_u13_u7_U5 (.A( u1_u13_u7_n149 ) , .ZN( u1_u13_u7_n175 ) );
  AOI21_X1 u1_u13_u7_U50 (.ZN( u1_u13_u7_n105 ) , .B2( u1_u13_u7_n110 ) , .A( u1_u13_u7_n125 ) , .B1( u1_u13_u7_n147 ) );
  NAND2_X1 u1_u13_u7_U51 (.ZN( u1_u13_u7_n146 ) , .A1( u1_u13_u7_n95 ) , .A2( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U52 (.A2( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n147 ) , .A1( u1_u13_u7_n93 ) );
  NAND2_X1 u1_u13_u7_U53 (.A1( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n127 ) , .A2( u1_u13_u7_n99 ) );
  OR2_X1 u1_u13_u7_U54 (.ZN( u1_u13_u7_n126 ) , .A2( u1_u13_u7_n152 ) , .A1( u1_u13_u7_n156 ) );
  NAND2_X1 u1_u13_u7_U55 (.A2( u1_u13_u7_n102 ) , .A1( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n133 ) );
  NAND2_X1 u1_u13_u7_U56 (.ZN( u1_u13_u7_n112 ) , .A2( u1_u13_u7_n96 ) , .A1( u1_u13_u7_n99 ) );
  NAND2_X1 u1_u13_u7_U57 (.A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n128 ) , .A1( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U58 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n113 ) , .A2( u1_u13_u7_n93 ) );
  NAND2_X1 u1_u13_u7_U59 (.A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n124 ) , .A1( u1_u13_u7_n96 ) );
  INV_X1 u1_u13_u7_U6 (.A( u1_u13_u7_n154 ) , .ZN( u1_u13_u7_n178 ) );
  NAND2_X1 u1_u13_u7_U60 (.ZN( u1_u13_u7_n110 ) , .A1( u1_u13_u7_n95 ) , .A2( u1_u13_u7_n96 ) );
  INV_X1 u1_u13_u7_U61 (.A( u1_u13_u7_n150 ) , .ZN( u1_u13_u7_n164 ) );
  AND2_X1 u1_u13_u7_U62 (.ZN( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n93 ) , .A2( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U63 (.A1( u1_u13_u7_n100 ) , .A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n129 ) );
  NAND2_X1 u1_u13_u7_U64 (.A2( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n131 ) , .A1( u1_u13_u7_n95 ) );
  NAND2_X1 u1_u13_u7_U65 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n138 ) , .A2( u1_u13_u7_n99 ) );
  NAND2_X1 u1_u13_u7_U66 (.ZN( u1_u13_u7_n132 ) , .A1( u1_u13_u7_n93 ) , .A2( u1_u13_u7_n96 ) );
  NAND2_X1 u1_u13_u7_U67 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n148 ) , .A2( u1_u13_u7_n95 ) );
  NOR2_X1 u1_u13_u7_U68 (.A2( u1_u13_X_47 ) , .ZN( u1_u13_u7_n150 ) , .A1( u1_u13_u7_n163 ) );
  NOR2_X1 u1_u13_u7_U69 (.A2( u1_u13_X_43 ) , .A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n103 ) );
  AOI211_X1 u1_u13_u7_U7 (.ZN( u1_u13_u7_n116 ) , .A( u1_u13_u7_n155 ) , .C1( u1_u13_u7_n161 ) , .C2( u1_u13_u7_n171 ) , .B( u1_u13_u7_n94 ) );
  NOR2_X1 u1_u13_u7_U70 (.A2( u1_u13_X_48 ) , .A1( u1_u13_u7_n166 ) , .ZN( u1_u13_u7_n95 ) );
  NOR2_X1 u1_u13_u7_U71 (.A2( u1_u13_X_45 ) , .A1( u1_u13_X_48 ) , .ZN( u1_u13_u7_n99 ) );
  NOR2_X1 u1_u13_u7_U72 (.A2( u1_u13_X_44 ) , .A1( u1_u13_u7_n167 ) , .ZN( u1_u13_u7_n98 ) );
  NOR2_X1 u1_u13_u7_U73 (.A2( u1_u13_X_46 ) , .A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n152 ) );
  AND2_X1 u1_u13_u7_U74 (.A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n156 ) , .A2( u1_u13_u7_n163 ) );
  NAND2_X1 u1_u13_u7_U75 (.A2( u1_u13_X_46 ) , .A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n125 ) );
  AND2_X1 u1_u13_u7_U76 (.A2( u1_u13_X_45 ) , .A1( u1_u13_X_48 ) , .ZN( u1_u13_u7_n102 ) );
  AND2_X1 u1_u13_u7_U77 (.A2( u1_u13_X_43 ) , .A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n96 ) );
  AND2_X1 u1_u13_u7_U78 (.A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n100 ) , .A2( u1_u13_u7_n167 ) );
  AND2_X1 u1_u13_u7_U79 (.A1( u1_u13_X_48 ) , .A2( u1_u13_u7_n166 ) , .ZN( u1_u13_u7_n93 ) );
  OAI222_X1 u1_u13_u7_U8 (.C2( u1_u13_u7_n101 ) , .B2( u1_u13_u7_n111 ) , .A1( u1_u13_u7_n113 ) , .C1( u1_u13_u7_n146 ) , .A2( u1_u13_u7_n162 ) , .B1( u1_u13_u7_n164 ) , .ZN( u1_u13_u7_n94 ) );
  INV_X1 u1_u13_u7_U80 (.A( u1_u13_X_46 ) , .ZN( u1_u13_u7_n163 ) );
  INV_X1 u1_u13_u7_U81 (.A( u1_u13_X_43 ) , .ZN( u1_u13_u7_n167 ) );
  INV_X1 u1_u13_u7_U82 (.A( u1_u13_X_45 ) , .ZN( u1_u13_u7_n166 ) );
  NAND4_X1 u1_u13_u7_U83 (.ZN( u1_out13_5 ) , .A4( u1_u13_u7_n108 ) , .A3( u1_u13_u7_n109 ) , .A1( u1_u13_u7_n116 ) , .A2( u1_u13_u7_n123 ) );
  AOI22_X1 u1_u13_u7_U84 (.ZN( u1_u13_u7_n109 ) , .A2( u1_u13_u7_n126 ) , .B2( u1_u13_u7_n145 ) , .B1( u1_u13_u7_n156 ) , .A1( u1_u13_u7_n171 ) );
  NOR4_X1 u1_u13_u7_U85 (.A4( u1_u13_u7_n104 ) , .A3( u1_u13_u7_n105 ) , .A2( u1_u13_u7_n106 ) , .A1( u1_u13_u7_n107 ) , .ZN( u1_u13_u7_n108 ) );
  NAND4_X1 u1_u13_u7_U86 (.ZN( u1_out13_27 ) , .A4( u1_u13_u7_n118 ) , .A3( u1_u13_u7_n119 ) , .A2( u1_u13_u7_n120 ) , .A1( u1_u13_u7_n121 ) );
  OAI21_X1 u1_u13_u7_U87 (.ZN( u1_u13_u7_n121 ) , .B2( u1_u13_u7_n145 ) , .A( u1_u13_u7_n150 ) , .B1( u1_u13_u7_n174 ) );
  OAI21_X1 u1_u13_u7_U88 (.ZN( u1_u13_u7_n120 ) , .A( u1_u13_u7_n161 ) , .B2( u1_u13_u7_n170 ) , .B1( u1_u13_u7_n179 ) );
  NAND4_X1 u1_u13_u7_U89 (.ZN( u1_out13_21 ) , .A4( u1_u13_u7_n157 ) , .A3( u1_u13_u7_n158 ) , .A2( u1_u13_u7_n159 ) , .A1( u1_u13_u7_n160 ) );
  OAI221_X1 u1_u13_u7_U9 (.C1( u1_u13_u7_n101 ) , .C2( u1_u13_u7_n147 ) , .ZN( u1_u13_u7_n155 ) , .B2( u1_u13_u7_n162 ) , .A( u1_u13_u7_n91 ) , .B1( u1_u13_u7_n92 ) );
  OAI21_X1 u1_u13_u7_U90 (.B1( u1_u13_u7_n145 ) , .ZN( u1_u13_u7_n160 ) , .A( u1_u13_u7_n161 ) , .B2( u1_u13_u7_n177 ) );
  AOI22_X1 u1_u13_u7_U91 (.B2( u1_u13_u7_n149 ) , .B1( u1_u13_u7_n150 ) , .A2( u1_u13_u7_n151 ) , .A1( u1_u13_u7_n152 ) , .ZN( u1_u13_u7_n158 ) );
  NAND4_X1 u1_u13_u7_U92 (.ZN( u1_out13_15 ) , .A4( u1_u13_u7_n142 ) , .A3( u1_u13_u7_n143 ) , .A2( u1_u13_u7_n144 ) , .A1( u1_u13_u7_n178 ) );
  OR2_X1 u1_u13_u7_U93 (.A2( u1_u13_u7_n125 ) , .A1( u1_u13_u7_n129 ) , .ZN( u1_u13_u7_n144 ) );
  AOI22_X1 u1_u13_u7_U94 (.A2( u1_u13_u7_n126 ) , .ZN( u1_u13_u7_n143 ) , .B2( u1_u13_u7_n165 ) , .B1( u1_u13_u7_n173 ) , .A1( u1_u13_u7_n174 ) );
  NAND3_X1 u1_u13_u7_U95 (.A3( u1_u13_u7_n146 ) , .A2( u1_u13_u7_n147 ) , .A1( u1_u13_u7_n148 ) , .ZN( u1_u13_u7_n151 ) );
  NAND3_X1 u1_u13_u7_U96 (.A3( u1_u13_u7_n131 ) , .A2( u1_u13_u7_n132 ) , .A1( u1_u13_u7_n133 ) , .ZN( u1_u13_u7_n135 ) );
  XOR2_X1 u1_u14_U11 (.B( u1_K15_44 ) , .A( u1_R13_29 ) , .Z( u1_u14_X_44 ) );
  XOR2_X1 u1_u14_U12 (.B( u1_K15_43 ) , .A( u1_R13_28 ) , .Z( u1_u14_X_43 ) );
  XOR2_X1 u1_u14_U13 (.B( u1_K15_42 ) , .A( u1_R13_29 ) , .Z( u1_u14_X_42 ) );
  XOR2_X1 u1_u14_U14 (.B( u1_K15_41 ) , .A( u1_R13_28 ) , .Z( u1_u14_X_41 ) );
  XOR2_X1 u1_u14_U18 (.B( u1_K15_38 ) , .A( u1_R13_25 ) , .Z( u1_u14_X_38 ) );
  XOR2_X1 u1_u14_U19 (.B( u1_K15_37 ) , .A( u1_R13_24 ) , .Z( u1_u14_X_37 ) );
  XOR2_X1 u1_u14_U2 (.B( u1_K15_8 ) , .A( u1_R13_5 ) , .Z( u1_u14_X_8 ) );
  XOR2_X1 u1_u14_U20 (.B( u1_K15_36 ) , .A( u1_R13_25 ) , .Z( u1_u14_X_36 ) );
  XOR2_X1 u1_u14_U21 (.B( u1_K15_35 ) , .A( u1_R13_24 ) , .Z( u1_u14_X_35 ) );
  XOR2_X1 u1_u14_U24 (.B( u1_K15_32 ) , .A( u1_R13_21 ) , .Z( u1_u14_X_32 ) );
  XOR2_X1 u1_u14_U25 (.B( u1_K15_31 ) , .A( u1_R13_20 ) , .Z( u1_u14_X_31 ) );
  XOR2_X1 u1_u14_U26 (.B( u1_K15_30 ) , .A( u1_R13_21 ) , .Z( u1_u14_X_30 ) );
  XOR2_X1 u1_u14_U27 (.B( u1_K15_2 ) , .A( u1_R13_1 ) , .Z( u1_u14_X_2 ) );
  XOR2_X1 u1_u14_U28 (.B( u1_K15_29 ) , .A( u1_R13_20 ) , .Z( u1_u14_X_29 ) );
  XOR2_X1 u1_u14_U3 (.B( u1_K15_7 ) , .A( u1_R13_4 ) , .Z( u1_u14_X_7 ) );
  XOR2_X1 u1_u14_U31 (.B( u1_K15_26 ) , .A( u1_R13_17 ) , .Z( u1_u14_X_26 ) );
  XOR2_X1 u1_u14_U32 (.B( u1_K15_25 ) , .A( u1_R13_16 ) , .Z( u1_u14_X_25 ) );
  XOR2_X1 u1_u14_U33 (.B( u1_K15_24 ) , .A( u1_R13_17 ) , .Z( u1_u14_X_24 ) );
  XOR2_X1 u1_u14_U34 (.B( u1_K15_23 ) , .A( u1_R13_16 ) , .Z( u1_u14_X_23 ) );
  XOR2_X1 u1_u14_U37 (.B( u1_K15_20 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_20 ) );
  XOR2_X1 u1_u14_U4 (.B( u1_K15_6 ) , .A( u1_R13_5 ) , .Z( u1_u14_X_6 ) );
  XOR2_X1 u1_u14_U40 (.B( u1_K15_18 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_18 ) );
  XOR2_X1 u1_u14_U44 (.B( u1_K15_14 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_14 ) );
  XOR2_X1 u1_u14_U45 (.B( u1_K15_13 ) , .A( u1_R13_8 ) , .Z( u1_u14_X_13 ) );
  XOR2_X1 u1_u14_U46 (.B( u1_K15_12 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_12 ) );
  XOR2_X1 u1_u14_U47 (.B( u1_K15_11 ) , .A( u1_R13_8 ) , .Z( u1_u14_X_11 ) );
  XOR2_X1 u1_u14_U5 (.B( u1_K15_5 ) , .A( u1_R13_4 ) , .Z( u1_u14_X_5 ) );
  XOR2_X1 u1_u14_U7 (.B( u1_K15_48 ) , .A( u1_R13_1 ) , .Z( u1_u14_X_48 ) );
  AND3_X1 u1_u14_u0_U10 (.A2( u1_u14_u0_n112 ) , .ZN( u1_u14_u0_n127 ) , .A3( u1_u14_u0_n130 ) , .A1( u1_u14_u0_n148 ) );
  NAND2_X1 u1_u14_u0_U11 (.ZN( u1_u14_u0_n113 ) , .A1( u1_u14_u0_n139 ) , .A2( u1_u14_u0_n149 ) );
  AND2_X1 u1_u14_u0_U12 (.ZN( u1_u14_u0_n107 ) , .A1( u1_u14_u0_n130 ) , .A2( u1_u14_u0_n140 ) );
  AND2_X1 u1_u14_u0_U13 (.A2( u1_u14_u0_n129 ) , .A1( u1_u14_u0_n130 ) , .ZN( u1_u14_u0_n151 ) );
  AND2_X1 u1_u14_u0_U14 (.A1( u1_u14_u0_n108 ) , .A2( u1_u14_u0_n125 ) , .ZN( u1_u14_u0_n145 ) );
  INV_X1 u1_u14_u0_U15 (.A( u1_u14_u0_n143 ) , .ZN( u1_u14_u0_n173 ) );
  NOR2_X1 u1_u14_u0_U16 (.A2( u1_u14_u0_n136 ) , .ZN( u1_u14_u0_n147 ) , .A1( u1_u14_u0_n160 ) );
  NOR2_X1 u1_u14_u0_U17 (.A1( u1_u14_u0_n163 ) , .A2( u1_u14_u0_n164 ) , .ZN( u1_u14_u0_n95 ) );
  AOI21_X1 u1_u14_u0_U18 (.B1( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n132 ) , .A( u1_u14_u0_n165 ) , .B2( u1_u14_u0_n93 ) );
  INV_X1 u1_u14_u0_U19 (.A( u1_u14_u0_n142 ) , .ZN( u1_u14_u0_n165 ) );
  OAI221_X1 u1_u14_u0_U20 (.C1( u1_u14_u0_n121 ) , .ZN( u1_u14_u0_n122 ) , .B2( u1_u14_u0_n127 ) , .A( u1_u14_u0_n143 ) , .B1( u1_u14_u0_n144 ) , .C2( u1_u14_u0_n147 ) );
  OAI22_X1 u1_u14_u0_U21 (.B1( u1_u14_u0_n125 ) , .ZN( u1_u14_u0_n126 ) , .A1( u1_u14_u0_n138 ) , .A2( u1_u14_u0_n146 ) , .B2( u1_u14_u0_n147 ) );
  OAI22_X1 u1_u14_u0_U22 (.B1( u1_u14_u0_n131 ) , .A1( u1_u14_u0_n144 ) , .B2( u1_u14_u0_n147 ) , .A2( u1_u14_u0_n90 ) , .ZN( u1_u14_u0_n91 ) );
  AND3_X1 u1_u14_u0_U23 (.A3( u1_u14_u0_n121 ) , .A2( u1_u14_u0_n125 ) , .A1( u1_u14_u0_n148 ) , .ZN( u1_u14_u0_n90 ) );
  NAND2_X1 u1_u14_u0_U24 (.A1( u1_u14_u0_n100 ) , .A2( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n125 ) );
  INV_X1 u1_u14_u0_U25 (.A( u1_u14_u0_n136 ) , .ZN( u1_u14_u0_n161 ) );
  NOR2_X1 u1_u14_u0_U26 (.A1( u1_u14_u0_n120 ) , .ZN( u1_u14_u0_n143 ) , .A2( u1_u14_u0_n167 ) );
  OAI221_X1 u1_u14_u0_U27 (.C1( u1_u14_u0_n112 ) , .ZN( u1_u14_u0_n120 ) , .B1( u1_u14_u0_n138 ) , .B2( u1_u14_u0_n141 ) , .C2( u1_u14_u0_n147 ) , .A( u1_u14_u0_n172 ) );
  AOI211_X1 u1_u14_u0_U28 (.B( u1_u14_u0_n115 ) , .A( u1_u14_u0_n116 ) , .C2( u1_u14_u0_n117 ) , .C1( u1_u14_u0_n118 ) , .ZN( u1_u14_u0_n119 ) );
  AOI22_X1 u1_u14_u0_U29 (.B2( u1_u14_u0_n109 ) , .A2( u1_u14_u0_n110 ) , .ZN( u1_u14_u0_n111 ) , .B1( u1_u14_u0_n118 ) , .A1( u1_u14_u0_n160 ) );
  INV_X1 u1_u14_u0_U3 (.A( u1_u14_u0_n113 ) , .ZN( u1_u14_u0_n166 ) );
  NAND2_X1 u1_u14_u0_U30 (.A1( u1_u14_u0_n100 ) , .ZN( u1_u14_u0_n129 ) , .A2( u1_u14_u0_n95 ) );
  INV_X1 u1_u14_u0_U31 (.A( u1_u14_u0_n118 ) , .ZN( u1_u14_u0_n158 ) );
  AOI21_X1 u1_u14_u0_U32 (.ZN( u1_u14_u0_n104 ) , .B1( u1_u14_u0_n107 ) , .B2( u1_u14_u0_n141 ) , .A( u1_u14_u0_n144 ) );
  AOI21_X1 u1_u14_u0_U33 (.B1( u1_u14_u0_n127 ) , .B2( u1_u14_u0_n129 ) , .A( u1_u14_u0_n138 ) , .ZN( u1_u14_u0_n96 ) );
  AOI21_X1 u1_u14_u0_U34 (.ZN( u1_u14_u0_n116 ) , .B2( u1_u14_u0_n142 ) , .A( u1_u14_u0_n144 ) , .B1( u1_u14_u0_n166 ) );
  NAND2_X1 u1_u14_u0_U35 (.A2( u1_u14_u0_n100 ) , .A1( u1_u14_u0_n101 ) , .ZN( u1_u14_u0_n139 ) );
  NAND2_X1 u1_u14_u0_U36 (.A2( u1_u14_u0_n100 ) , .ZN( u1_u14_u0_n131 ) , .A1( u1_u14_u0_n92 ) );
  NAND2_X1 u1_u14_u0_U37 (.A1( u1_u14_u0_n101 ) , .A2( u1_u14_u0_n102 ) , .ZN( u1_u14_u0_n150 ) );
  INV_X1 u1_u14_u0_U38 (.A( u1_u14_u0_n138 ) , .ZN( u1_u14_u0_n160 ) );
  NAND2_X1 u1_u14_u0_U39 (.A1( u1_u14_u0_n102 ) , .ZN( u1_u14_u0_n128 ) , .A2( u1_u14_u0_n95 ) );
  AOI21_X1 u1_u14_u0_U4 (.B1( u1_u14_u0_n114 ) , .ZN( u1_u14_u0_n115 ) , .B2( u1_u14_u0_n129 ) , .A( u1_u14_u0_n161 ) );
  NAND2_X1 u1_u14_u0_U40 (.ZN( u1_u14_u0_n148 ) , .A1( u1_u14_u0_n93 ) , .A2( u1_u14_u0_n95 ) );
  NAND2_X1 u1_u14_u0_U41 (.A2( u1_u14_u0_n102 ) , .A1( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n149 ) );
  NAND2_X1 u1_u14_u0_U42 (.A2( u1_u14_u0_n102 ) , .ZN( u1_u14_u0_n114 ) , .A1( u1_u14_u0_n92 ) );
  NAND2_X1 u1_u14_u0_U43 (.A2( u1_u14_u0_n101 ) , .ZN( u1_u14_u0_n121 ) , .A1( u1_u14_u0_n93 ) );
  INV_X1 u1_u14_u0_U44 (.ZN( u1_u14_u0_n172 ) , .A( u1_u14_u0_n88 ) );
  OAI222_X1 u1_u14_u0_U45 (.C1( u1_u14_u0_n108 ) , .A1( u1_u14_u0_n125 ) , .B2( u1_u14_u0_n128 ) , .B1( u1_u14_u0_n144 ) , .A2( u1_u14_u0_n158 ) , .C2( u1_u14_u0_n161 ) , .ZN( u1_u14_u0_n88 ) );
  NAND2_X1 u1_u14_u0_U46 (.ZN( u1_u14_u0_n112 ) , .A2( u1_u14_u0_n92 ) , .A1( u1_u14_u0_n93 ) );
  OR3_X1 u1_u14_u0_U47 (.A3( u1_u14_u0_n152 ) , .A2( u1_u14_u0_n153 ) , .A1( u1_u14_u0_n154 ) , .ZN( u1_u14_u0_n155 ) );
  AOI21_X1 u1_u14_u0_U48 (.B2( u1_u14_u0_n150 ) , .B1( u1_u14_u0_n151 ) , .ZN( u1_u14_u0_n152 ) , .A( u1_u14_u0_n158 ) );
  AOI21_X1 u1_u14_u0_U49 (.A( u1_u14_u0_n144 ) , .B2( u1_u14_u0_n145 ) , .B1( u1_u14_u0_n146 ) , .ZN( u1_u14_u0_n154 ) );
  AOI21_X1 u1_u14_u0_U5 (.B2( u1_u14_u0_n131 ) , .ZN( u1_u14_u0_n134 ) , .B1( u1_u14_u0_n151 ) , .A( u1_u14_u0_n158 ) );
  AOI21_X1 u1_u14_u0_U50 (.A( u1_u14_u0_n147 ) , .B2( u1_u14_u0_n148 ) , .B1( u1_u14_u0_n149 ) , .ZN( u1_u14_u0_n153 ) );
  INV_X1 u1_u14_u0_U51 (.ZN( u1_u14_u0_n171 ) , .A( u1_u14_u0_n99 ) );
  OAI211_X1 u1_u14_u0_U52 (.C2( u1_u14_u0_n140 ) , .C1( u1_u14_u0_n161 ) , .A( u1_u14_u0_n169 ) , .B( u1_u14_u0_n98 ) , .ZN( u1_u14_u0_n99 ) );
  AOI211_X1 u1_u14_u0_U53 (.C1( u1_u14_u0_n118 ) , .A( u1_u14_u0_n123 ) , .B( u1_u14_u0_n96 ) , .C2( u1_u14_u0_n97 ) , .ZN( u1_u14_u0_n98 ) );
  INV_X1 u1_u14_u0_U54 (.ZN( u1_u14_u0_n169 ) , .A( u1_u14_u0_n91 ) );
  NOR2_X1 u1_u14_u0_U55 (.A2( u1_u14_X_4 ) , .A1( u1_u14_X_5 ) , .ZN( u1_u14_u0_n118 ) );
  NOR2_X1 u1_u14_u0_U56 (.A2( u1_u14_X_2 ) , .ZN( u1_u14_u0_n103 ) , .A1( u1_u14_u0_n164 ) );
  NOR2_X1 u1_u14_u0_U57 (.A2( u1_u14_X_1 ) , .A1( u1_u14_X_2 ) , .ZN( u1_u14_u0_n92 ) );
  NOR2_X1 u1_u14_u0_U58 (.A2( u1_u14_X_1 ) , .ZN( u1_u14_u0_n101 ) , .A1( u1_u14_u0_n163 ) );
  NAND2_X1 u1_u14_u0_U59 (.A2( u1_u14_X_4 ) , .A1( u1_u14_X_5 ) , .ZN( u1_u14_u0_n144 ) );
  NOR2_X1 u1_u14_u0_U6 (.A1( u1_u14_u0_n108 ) , .ZN( u1_u14_u0_n123 ) , .A2( u1_u14_u0_n158 ) );
  NOR2_X1 u1_u14_u0_U60 (.A2( u1_u14_X_5 ) , .ZN( u1_u14_u0_n136 ) , .A1( u1_u14_u0_n159 ) );
  NAND2_X1 u1_u14_u0_U61 (.A1( u1_u14_X_5 ) , .ZN( u1_u14_u0_n138 ) , .A2( u1_u14_u0_n159 ) );
  AND2_X1 u1_u14_u0_U62 (.A2( u1_u14_X_3 ) , .A1( u1_u14_X_6 ) , .ZN( u1_u14_u0_n102 ) );
  AND2_X1 u1_u14_u0_U63 (.A1( u1_u14_X_6 ) , .A2( u1_u14_u0_n162 ) , .ZN( u1_u14_u0_n93 ) );
  INV_X1 u1_u14_u0_U64 (.A( u1_u14_X_4 ) , .ZN( u1_u14_u0_n159 ) );
  INV_X1 u1_u14_u0_U65 (.A( u1_u14_X_1 ) , .ZN( u1_u14_u0_n164 ) );
  INV_X1 u1_u14_u0_U66 (.A( u1_u14_X_2 ) , .ZN( u1_u14_u0_n163 ) );
  INV_X1 u1_u14_u0_U67 (.A( u1_u14_X_3 ) , .ZN( u1_u14_u0_n162 ) );
  INV_X1 u1_u14_u0_U68 (.A( u1_u14_u0_n126 ) , .ZN( u1_u14_u0_n168 ) );
  AOI211_X1 u1_u14_u0_U69 (.B( u1_u14_u0_n133 ) , .A( u1_u14_u0_n134 ) , .C2( u1_u14_u0_n135 ) , .C1( u1_u14_u0_n136 ) , .ZN( u1_u14_u0_n137 ) );
  OAI21_X1 u1_u14_u0_U7 (.B1( u1_u14_u0_n150 ) , .B2( u1_u14_u0_n158 ) , .A( u1_u14_u0_n172 ) , .ZN( u1_u14_u0_n89 ) );
  INV_X1 u1_u14_u0_U70 (.ZN( u1_u14_u0_n174 ) , .A( u1_u14_u0_n89 ) );
  AOI211_X1 u1_u14_u0_U71 (.B( u1_u14_u0_n104 ) , .A( u1_u14_u0_n105 ) , .ZN( u1_u14_u0_n106 ) , .C2( u1_u14_u0_n113 ) , .C1( u1_u14_u0_n160 ) );
  OR4_X1 u1_u14_u0_U72 (.ZN( u1_out14_17 ) , .A4( u1_u14_u0_n122 ) , .A2( u1_u14_u0_n123 ) , .A1( u1_u14_u0_n124 ) , .A3( u1_u14_u0_n170 ) );
  AOI21_X1 u1_u14_u0_U73 (.B2( u1_u14_u0_n107 ) , .ZN( u1_u14_u0_n124 ) , .B1( u1_u14_u0_n128 ) , .A( u1_u14_u0_n161 ) );
  INV_X1 u1_u14_u0_U74 (.A( u1_u14_u0_n111 ) , .ZN( u1_u14_u0_n170 ) );
  OR4_X1 u1_u14_u0_U75 (.ZN( u1_out14_31 ) , .A4( u1_u14_u0_n155 ) , .A2( u1_u14_u0_n156 ) , .A1( u1_u14_u0_n157 ) , .A3( u1_u14_u0_n173 ) );
  AOI21_X1 u1_u14_u0_U76 (.A( u1_u14_u0_n138 ) , .B2( u1_u14_u0_n139 ) , .B1( u1_u14_u0_n140 ) , .ZN( u1_u14_u0_n157 ) );
  AOI21_X1 u1_u14_u0_U77 (.B2( u1_u14_u0_n141 ) , .B1( u1_u14_u0_n142 ) , .ZN( u1_u14_u0_n156 ) , .A( u1_u14_u0_n161 ) );
  AOI21_X1 u1_u14_u0_U78 (.B1( u1_u14_u0_n132 ) , .ZN( u1_u14_u0_n133 ) , .A( u1_u14_u0_n144 ) , .B2( u1_u14_u0_n166 ) );
  OAI22_X1 u1_u14_u0_U79 (.ZN( u1_u14_u0_n105 ) , .A2( u1_u14_u0_n132 ) , .B1( u1_u14_u0_n146 ) , .A1( u1_u14_u0_n147 ) , .B2( u1_u14_u0_n161 ) );
  AND2_X1 u1_u14_u0_U8 (.A1( u1_u14_u0_n114 ) , .A2( u1_u14_u0_n121 ) , .ZN( u1_u14_u0_n146 ) );
  NAND2_X1 u1_u14_u0_U80 (.ZN( u1_u14_u0_n110 ) , .A2( u1_u14_u0_n132 ) , .A1( u1_u14_u0_n145 ) );
  INV_X1 u1_u14_u0_U81 (.A( u1_u14_u0_n119 ) , .ZN( u1_u14_u0_n167 ) );
  NAND2_X1 u1_u14_u0_U82 (.A2( u1_u14_u0_n103 ) , .ZN( u1_u14_u0_n140 ) , .A1( u1_u14_u0_n94 ) );
  NAND2_X1 u1_u14_u0_U83 (.A1( u1_u14_u0_n101 ) , .ZN( u1_u14_u0_n130 ) , .A2( u1_u14_u0_n94 ) );
  NAND2_X1 u1_u14_u0_U84 (.ZN( u1_u14_u0_n108 ) , .A1( u1_u14_u0_n92 ) , .A2( u1_u14_u0_n94 ) );
  NAND2_X1 u1_u14_u0_U85 (.ZN( u1_u14_u0_n142 ) , .A1( u1_u14_u0_n94 ) , .A2( u1_u14_u0_n95 ) );
  NOR2_X1 u1_u14_u0_U86 (.A2( u1_u14_X_6 ) , .ZN( u1_u14_u0_n100 ) , .A1( u1_u14_u0_n162 ) );
  NOR2_X1 u1_u14_u0_U87 (.A2( u1_u14_X_3 ) , .A1( u1_u14_X_6 ) , .ZN( u1_u14_u0_n94 ) );
  NAND3_X1 u1_u14_u0_U88 (.ZN( u1_out14_23 ) , .A3( u1_u14_u0_n137 ) , .A1( u1_u14_u0_n168 ) , .A2( u1_u14_u0_n171 ) );
  NAND3_X1 u1_u14_u0_U89 (.A3( u1_u14_u0_n127 ) , .A2( u1_u14_u0_n128 ) , .ZN( u1_u14_u0_n135 ) , .A1( u1_u14_u0_n150 ) );
  AND2_X1 u1_u14_u0_U9 (.A1( u1_u14_u0_n131 ) , .ZN( u1_u14_u0_n141 ) , .A2( u1_u14_u0_n150 ) );
  NAND3_X1 u1_u14_u0_U90 (.ZN( u1_u14_u0_n117 ) , .A3( u1_u14_u0_n132 ) , .A2( u1_u14_u0_n139 ) , .A1( u1_u14_u0_n148 ) );
  NAND3_X1 u1_u14_u0_U91 (.ZN( u1_u14_u0_n109 ) , .A2( u1_u14_u0_n114 ) , .A3( u1_u14_u0_n140 ) , .A1( u1_u14_u0_n149 ) );
  NAND3_X1 u1_u14_u0_U92 (.ZN( u1_out14_9 ) , .A3( u1_u14_u0_n106 ) , .A2( u1_u14_u0_n171 ) , .A1( u1_u14_u0_n174 ) );
  NAND3_X1 u1_u14_u0_U93 (.A2( u1_u14_u0_n128 ) , .A1( u1_u14_u0_n132 ) , .A3( u1_u14_u0_n146 ) , .ZN( u1_u14_u0_n97 ) );
  AOI21_X1 u1_u14_u1_U10 (.ZN( u1_u14_u1_n106 ) , .A( u1_u14_u1_n112 ) , .B1( u1_u14_u1_n154 ) , .B2( u1_u14_u1_n156 ) );
  NAND3_X1 u1_u14_u1_U100 (.ZN( u1_u14_u1_n113 ) , .A1( u1_u14_u1_n120 ) , .A3( u1_u14_u1_n133 ) , .A2( u1_u14_u1_n155 ) );
  INV_X1 u1_u14_u1_U11 (.A( u1_u14_u1_n101 ) , .ZN( u1_u14_u1_n184 ) );
  AOI21_X1 u1_u14_u1_U12 (.ZN( u1_u14_u1_n107 ) , .B1( u1_u14_u1_n134 ) , .B2( u1_u14_u1_n149 ) , .A( u1_u14_u1_n174 ) );
  NAND2_X1 u1_u14_u1_U13 (.ZN( u1_u14_u1_n140 ) , .A2( u1_u14_u1_n150 ) , .A1( u1_u14_u1_n155 ) );
  NAND2_X1 u1_u14_u1_U14 (.A1( u1_u14_u1_n131 ) , .ZN( u1_u14_u1_n147 ) , .A2( u1_u14_u1_n153 ) );
  AOI22_X1 u1_u14_u1_U15 (.B2( u1_u14_u1_n136 ) , .A2( u1_u14_u1_n137 ) , .ZN( u1_u14_u1_n143 ) , .A1( u1_u14_u1_n171 ) , .B1( u1_u14_u1_n173 ) );
  INV_X1 u1_u14_u1_U16 (.A( u1_u14_u1_n147 ) , .ZN( u1_u14_u1_n181 ) );
  INV_X1 u1_u14_u1_U17 (.A( u1_u14_u1_n139 ) , .ZN( u1_u14_u1_n174 ) );
  INV_X1 u1_u14_u1_U18 (.A( u1_u14_u1_n112 ) , .ZN( u1_u14_u1_n171 ) );
  NAND2_X1 u1_u14_u1_U19 (.ZN( u1_u14_u1_n141 ) , .A1( u1_u14_u1_n153 ) , .A2( u1_u14_u1_n156 ) );
  AND2_X1 u1_u14_u1_U20 (.A1( u1_u14_u1_n123 ) , .ZN( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n161 ) );
  NAND2_X1 u1_u14_u1_U21 (.A2( u1_u14_u1_n115 ) , .A1( u1_u14_u1_n116 ) , .ZN( u1_u14_u1_n148 ) );
  NAND2_X1 u1_u14_u1_U22 (.A2( u1_u14_u1_n133 ) , .A1( u1_u14_u1_n135 ) , .ZN( u1_u14_u1_n159 ) );
  NAND2_X1 u1_u14_u1_U23 (.A2( u1_u14_u1_n115 ) , .A1( u1_u14_u1_n120 ) , .ZN( u1_u14_u1_n132 ) );
  INV_X1 u1_u14_u1_U24 (.A( u1_u14_u1_n154 ) , .ZN( u1_u14_u1_n178 ) );
  AOI22_X1 u1_u14_u1_U25 (.B2( u1_u14_u1_n113 ) , .A2( u1_u14_u1_n114 ) , .ZN( u1_u14_u1_n125 ) , .A1( u1_u14_u1_n171 ) , .B1( u1_u14_u1_n173 ) );
  NAND2_X1 u1_u14_u1_U26 (.ZN( u1_u14_u1_n114 ) , .A1( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n156 ) );
  INV_X1 u1_u14_u1_U27 (.A( u1_u14_u1_n151 ) , .ZN( u1_u14_u1_n183 ) );
  AND2_X1 u1_u14_u1_U28 (.A1( u1_u14_u1_n129 ) , .A2( u1_u14_u1_n133 ) , .ZN( u1_u14_u1_n149 ) );
  INV_X1 u1_u14_u1_U29 (.A( u1_u14_u1_n131 ) , .ZN( u1_u14_u1_n180 ) );
  INV_X1 u1_u14_u1_U3 (.A( u1_u14_u1_n159 ) , .ZN( u1_u14_u1_n182 ) );
  AOI221_X1 u1_u14_u1_U30 (.B1( u1_u14_u1_n140 ) , .ZN( u1_u14_u1_n167 ) , .B2( u1_u14_u1_n172 ) , .C2( u1_u14_u1_n175 ) , .C1( u1_u14_u1_n178 ) , .A( u1_u14_u1_n188 ) );
  INV_X1 u1_u14_u1_U31 (.ZN( u1_u14_u1_n188 ) , .A( u1_u14_u1_n97 ) );
  AOI211_X1 u1_u14_u1_U32 (.A( u1_u14_u1_n118 ) , .C1( u1_u14_u1_n132 ) , .C2( u1_u14_u1_n139 ) , .B( u1_u14_u1_n96 ) , .ZN( u1_u14_u1_n97 ) );
  AOI21_X1 u1_u14_u1_U33 (.B2( u1_u14_u1_n121 ) , .B1( u1_u14_u1_n135 ) , .A( u1_u14_u1_n152 ) , .ZN( u1_u14_u1_n96 ) );
  OAI221_X1 u1_u14_u1_U34 (.A( u1_u14_u1_n119 ) , .C2( u1_u14_u1_n129 ) , .ZN( u1_u14_u1_n138 ) , .B2( u1_u14_u1_n152 ) , .C1( u1_u14_u1_n174 ) , .B1( u1_u14_u1_n187 ) );
  INV_X1 u1_u14_u1_U35 (.A( u1_u14_u1_n148 ) , .ZN( u1_u14_u1_n187 ) );
  AOI211_X1 u1_u14_u1_U36 (.B( u1_u14_u1_n117 ) , .A( u1_u14_u1_n118 ) , .ZN( u1_u14_u1_n119 ) , .C2( u1_u14_u1_n146 ) , .C1( u1_u14_u1_n159 ) );
  NOR2_X1 u1_u14_u1_U37 (.A1( u1_u14_u1_n168 ) , .A2( u1_u14_u1_n176 ) , .ZN( u1_u14_u1_n98 ) );
  AOI211_X1 u1_u14_u1_U38 (.B( u1_u14_u1_n162 ) , .A( u1_u14_u1_n163 ) , .C2( u1_u14_u1_n164 ) , .ZN( u1_u14_u1_n165 ) , .C1( u1_u14_u1_n171 ) );
  AOI21_X1 u1_u14_u1_U39 (.A( u1_u14_u1_n160 ) , .B2( u1_u14_u1_n161 ) , .ZN( u1_u14_u1_n162 ) , .B1( u1_u14_u1_n182 ) );
  AOI221_X1 u1_u14_u1_U4 (.A( u1_u14_u1_n138 ) , .C2( u1_u14_u1_n139 ) , .C1( u1_u14_u1_n140 ) , .B2( u1_u14_u1_n141 ) , .ZN( u1_u14_u1_n142 ) , .B1( u1_u14_u1_n175 ) );
  OR2_X1 u1_u14_u1_U40 (.A2( u1_u14_u1_n157 ) , .A1( u1_u14_u1_n158 ) , .ZN( u1_u14_u1_n163 ) );
  OAI21_X1 u1_u14_u1_U41 (.B2( u1_u14_u1_n123 ) , .ZN( u1_u14_u1_n145 ) , .B1( u1_u14_u1_n160 ) , .A( u1_u14_u1_n185 ) );
  INV_X1 u1_u14_u1_U42 (.A( u1_u14_u1_n122 ) , .ZN( u1_u14_u1_n185 ) );
  AOI21_X1 u1_u14_u1_U43 (.B2( u1_u14_u1_n120 ) , .B1( u1_u14_u1_n121 ) , .ZN( u1_u14_u1_n122 ) , .A( u1_u14_u1_n128 ) );
  NAND2_X1 u1_u14_u1_U44 (.A1( u1_u14_u1_n128 ) , .ZN( u1_u14_u1_n146 ) , .A2( u1_u14_u1_n160 ) );
  NAND2_X1 u1_u14_u1_U45 (.A2( u1_u14_u1_n112 ) , .ZN( u1_u14_u1_n139 ) , .A1( u1_u14_u1_n152 ) );
  NAND2_X1 u1_u14_u1_U46 (.A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n156 ) , .A2( u1_u14_u1_n99 ) );
  NOR2_X1 u1_u14_u1_U47 (.ZN( u1_u14_u1_n117 ) , .A1( u1_u14_u1_n121 ) , .A2( u1_u14_u1_n160 ) );
  AOI21_X1 u1_u14_u1_U48 (.A( u1_u14_u1_n128 ) , .B2( u1_u14_u1_n129 ) , .ZN( u1_u14_u1_n130 ) , .B1( u1_u14_u1_n150 ) );
  NAND2_X1 u1_u14_u1_U49 (.ZN( u1_u14_u1_n112 ) , .A1( u1_u14_u1_n169 ) , .A2( u1_u14_u1_n170 ) );
  AOI211_X1 u1_u14_u1_U5 (.ZN( u1_u14_u1_n124 ) , .A( u1_u14_u1_n138 ) , .C2( u1_u14_u1_n139 ) , .B( u1_u14_u1_n145 ) , .C1( u1_u14_u1_n147 ) );
  NAND2_X1 u1_u14_u1_U50 (.ZN( u1_u14_u1_n129 ) , .A2( u1_u14_u1_n95 ) , .A1( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U51 (.A1( u1_u14_u1_n102 ) , .ZN( u1_u14_u1_n154 ) , .A2( u1_u14_u1_n99 ) );
  NAND2_X1 u1_u14_u1_U52 (.A2( u1_u14_u1_n100 ) , .ZN( u1_u14_u1_n135 ) , .A1( u1_u14_u1_n99 ) );
  AOI21_X1 u1_u14_u1_U53 (.A( u1_u14_u1_n152 ) , .B2( u1_u14_u1_n153 ) , .B1( u1_u14_u1_n154 ) , .ZN( u1_u14_u1_n158 ) );
  INV_X1 u1_u14_u1_U54 (.A( u1_u14_u1_n160 ) , .ZN( u1_u14_u1_n175 ) );
  NAND2_X1 u1_u14_u1_U55 (.A1( u1_u14_u1_n100 ) , .ZN( u1_u14_u1_n116 ) , .A2( u1_u14_u1_n95 ) );
  NAND2_X1 u1_u14_u1_U56 (.A1( u1_u14_u1_n102 ) , .ZN( u1_u14_u1_n131 ) , .A2( u1_u14_u1_n95 ) );
  NAND2_X1 u1_u14_u1_U57 (.A2( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n121 ) , .A1( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U58 (.A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n153 ) , .A2( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U59 (.A2( u1_u14_u1_n104 ) , .A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n133 ) );
  NOR2_X1 u1_u14_u1_U6 (.A1( u1_u14_u1_n112 ) , .A2( u1_u14_u1_n116 ) , .ZN( u1_u14_u1_n118 ) );
  NAND2_X1 u1_u14_u1_U60 (.ZN( u1_u14_u1_n150 ) , .A2( u1_u14_u1_n98 ) , .A1( u1_u14_u1_n99 ) );
  NAND2_X1 u1_u14_u1_U61 (.A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n155 ) , .A2( u1_u14_u1_n95 ) );
  OAI21_X1 u1_u14_u1_U62 (.ZN( u1_u14_u1_n109 ) , .B1( u1_u14_u1_n129 ) , .B2( u1_u14_u1_n160 ) , .A( u1_u14_u1_n167 ) );
  NAND2_X1 u1_u14_u1_U63 (.A2( u1_u14_u1_n100 ) , .A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n120 ) );
  NAND2_X1 u1_u14_u1_U64 (.A1( u1_u14_u1_n102 ) , .A2( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n115 ) );
  NAND2_X1 u1_u14_u1_U65 (.A2( u1_u14_u1_n100 ) , .A1( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n151 ) );
  NAND2_X1 u1_u14_u1_U66 (.A2( u1_u14_u1_n103 ) , .A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n161 ) );
  INV_X1 u1_u14_u1_U67 (.A( u1_u14_u1_n152 ) , .ZN( u1_u14_u1_n173 ) );
  INV_X1 u1_u14_u1_U68 (.A( u1_u14_u1_n128 ) , .ZN( u1_u14_u1_n172 ) );
  NAND2_X1 u1_u14_u1_U69 (.A2( u1_u14_u1_n102 ) , .A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n123 ) );
  OAI21_X1 u1_u14_u1_U7 (.ZN( u1_u14_u1_n101 ) , .B1( u1_u14_u1_n141 ) , .A( u1_u14_u1_n146 ) , .B2( u1_u14_u1_n183 ) );
  NOR2_X1 u1_u14_u1_U70 (.A2( u1_u14_X_7 ) , .A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n95 ) );
  NOR2_X1 u1_u14_u1_U71 (.A1( u1_u14_X_12 ) , .A2( u1_u14_X_9 ) , .ZN( u1_u14_u1_n100 ) );
  NOR2_X1 u1_u14_u1_U72 (.A2( u1_u14_X_8 ) , .A1( u1_u14_u1_n177 ) , .ZN( u1_u14_u1_n99 ) );
  NOR2_X1 u1_u14_u1_U73 (.A2( u1_u14_X_12 ) , .ZN( u1_u14_u1_n102 ) , .A1( u1_u14_u1_n176 ) );
  NOR2_X1 u1_u14_u1_U74 (.A2( u1_u14_X_9 ) , .ZN( u1_u14_u1_n105 ) , .A1( u1_u14_u1_n168 ) );
  NAND2_X1 u1_u14_u1_U75 (.A1( u1_u14_X_10 ) , .ZN( u1_u14_u1_n160 ) , .A2( u1_u14_u1_n169 ) );
  NAND2_X1 u1_u14_u1_U76 (.A2( u1_u14_X_10 ) , .A1( u1_u14_X_11 ) , .ZN( u1_u14_u1_n152 ) );
  NAND2_X1 u1_u14_u1_U77 (.A1( u1_u14_X_11 ) , .ZN( u1_u14_u1_n128 ) , .A2( u1_u14_u1_n170 ) );
  AND2_X1 u1_u14_u1_U78 (.A2( u1_u14_X_7 ) , .A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n104 ) );
  AND2_X1 u1_u14_u1_U79 (.A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n103 ) , .A2( u1_u14_u1_n177 ) );
  AOI21_X1 u1_u14_u1_U8 (.B2( u1_u14_u1_n155 ) , .B1( u1_u14_u1_n156 ) , .ZN( u1_u14_u1_n157 ) , .A( u1_u14_u1_n174 ) );
  INV_X1 u1_u14_u1_U80 (.A( u1_u14_X_10 ) , .ZN( u1_u14_u1_n170 ) );
  INV_X1 u1_u14_u1_U81 (.A( u1_u14_X_9 ) , .ZN( u1_u14_u1_n176 ) );
  INV_X1 u1_u14_u1_U82 (.A( u1_u14_X_11 ) , .ZN( u1_u14_u1_n169 ) );
  INV_X1 u1_u14_u1_U83 (.A( u1_u14_X_12 ) , .ZN( u1_u14_u1_n168 ) );
  INV_X1 u1_u14_u1_U84 (.A( u1_u14_X_7 ) , .ZN( u1_u14_u1_n177 ) );
  NAND4_X1 u1_u14_u1_U85 (.ZN( u1_out14_18 ) , .A4( u1_u14_u1_n165 ) , .A3( u1_u14_u1_n166 ) , .A1( u1_u14_u1_n167 ) , .A2( u1_u14_u1_n186 ) );
  AOI22_X1 u1_u14_u1_U86 (.B2( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n147 ) , .A2( u1_u14_u1_n148 ) , .ZN( u1_u14_u1_n166 ) , .A1( u1_u14_u1_n172 ) );
  INV_X1 u1_u14_u1_U87 (.A( u1_u14_u1_n145 ) , .ZN( u1_u14_u1_n186 ) );
  OR4_X1 u1_u14_u1_U88 (.ZN( u1_out14_13 ) , .A4( u1_u14_u1_n108 ) , .A3( u1_u14_u1_n109 ) , .A2( u1_u14_u1_n110 ) , .A1( u1_u14_u1_n111 ) );
  AOI21_X1 u1_u14_u1_U89 (.ZN( u1_u14_u1_n111 ) , .A( u1_u14_u1_n128 ) , .B2( u1_u14_u1_n131 ) , .B1( u1_u14_u1_n135 ) );
  OR4_X1 u1_u14_u1_U9 (.A4( u1_u14_u1_n106 ) , .A3( u1_u14_u1_n107 ) , .ZN( u1_u14_u1_n108 ) , .A1( u1_u14_u1_n117 ) , .A2( u1_u14_u1_n184 ) );
  AOI21_X1 u1_u14_u1_U90 (.ZN( u1_u14_u1_n110 ) , .A( u1_u14_u1_n116 ) , .B1( u1_u14_u1_n152 ) , .B2( u1_u14_u1_n160 ) );
  NAND4_X1 u1_u14_u1_U91 (.ZN( u1_out14_2 ) , .A4( u1_u14_u1_n142 ) , .A3( u1_u14_u1_n143 ) , .A2( u1_u14_u1_n144 ) , .A1( u1_u14_u1_n179 ) );
  OAI21_X1 u1_u14_u1_U92 (.B2( u1_u14_u1_n132 ) , .ZN( u1_u14_u1_n144 ) , .A( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n180 ) );
  INV_X1 u1_u14_u1_U93 (.A( u1_u14_u1_n130 ) , .ZN( u1_u14_u1_n179 ) );
  NAND4_X1 u1_u14_u1_U94 (.ZN( u1_out14_28 ) , .A4( u1_u14_u1_n124 ) , .A3( u1_u14_u1_n125 ) , .A2( u1_u14_u1_n126 ) , .A1( u1_u14_u1_n127 ) );
  OAI21_X1 u1_u14_u1_U95 (.ZN( u1_u14_u1_n127 ) , .B2( u1_u14_u1_n139 ) , .B1( u1_u14_u1_n175 ) , .A( u1_u14_u1_n183 ) );
  OAI21_X1 u1_u14_u1_U96 (.ZN( u1_u14_u1_n126 ) , .B2( u1_u14_u1_n140 ) , .A( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n178 ) );
  NAND3_X1 u1_u14_u1_U97 (.A3( u1_u14_u1_n149 ) , .A2( u1_u14_u1_n150 ) , .A1( u1_u14_u1_n151 ) , .ZN( u1_u14_u1_n164 ) );
  NAND3_X1 u1_u14_u1_U98 (.A3( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n135 ) , .ZN( u1_u14_u1_n136 ) , .A1( u1_u14_u1_n151 ) );
  NAND3_X1 u1_u14_u1_U99 (.A1( u1_u14_u1_n133 ) , .ZN( u1_u14_u1_n137 ) , .A2( u1_u14_u1_n154 ) , .A3( u1_u14_u1_n181 ) );
  OAI22_X1 u1_u14_u2_U10 (.ZN( u1_u14_u2_n109 ) , .A2( u1_u14_u2_n113 ) , .B2( u1_u14_u2_n133 ) , .B1( u1_u14_u2_n167 ) , .A1( u1_u14_u2_n168 ) );
  NAND3_X1 u1_u14_u2_U100 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n98 ) );
  OAI22_X1 u1_u14_u2_U11 (.B1( u1_u14_u2_n151 ) , .A2( u1_u14_u2_n152 ) , .A1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n160 ) , .B2( u1_u14_u2_n168 ) );
  NOR3_X1 u1_u14_u2_U12 (.A1( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n151 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U13 (.ZN( u1_u14_u2_n144 ) , .B2( u1_u14_u2_n155 ) , .A( u1_u14_u2_n172 ) , .B1( u1_u14_u2_n185 ) );
  AOI21_X1 u1_u14_u2_U14 (.B2( u1_u14_u2_n143 ) , .ZN( u1_u14_u2_n145 ) , .B1( u1_u14_u2_n152 ) , .A( u1_u14_u2_n171 ) );
  AOI21_X1 u1_u14_u2_U15 (.B2( u1_u14_u2_n120 ) , .B1( u1_u14_u2_n121 ) , .ZN( u1_u14_u2_n126 ) , .A( u1_u14_u2_n167 ) );
  INV_X1 u1_u14_u2_U16 (.A( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n171 ) );
  INV_X1 u1_u14_u2_U17 (.A( u1_u14_u2_n120 ) , .ZN( u1_u14_u2_n188 ) );
  NAND2_X1 u1_u14_u2_U18 (.A2( u1_u14_u2_n122 ) , .ZN( u1_u14_u2_n150 ) , .A1( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U19 (.A( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U20 (.A( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n173 ) );
  NAND2_X1 u1_u14_u2_U21 (.A1( u1_u14_u2_n132 ) , .A2( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n157 ) );
  INV_X1 u1_u14_u2_U22 (.A( u1_u14_u2_n113 ) , .ZN( u1_u14_u2_n178 ) );
  INV_X1 u1_u14_u2_U23 (.A( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n175 ) );
  INV_X1 u1_u14_u2_U24 (.A( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U25 (.A( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n177 ) );
  INV_X1 u1_u14_u2_U26 (.A( u1_u14_u2_n116 ) , .ZN( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U27 (.A( u1_u14_u2_n131 ) , .ZN( u1_u14_u2_n179 ) );
  INV_X1 u1_u14_u2_U28 (.A( u1_u14_u2_n154 ) , .ZN( u1_u14_u2_n176 ) );
  NAND2_X1 u1_u14_u2_U29 (.A2( u1_u14_u2_n116 ) , .A1( u1_u14_u2_n117 ) , .ZN( u1_u14_u2_n118 ) );
  NOR2_X1 u1_u14_u2_U3 (.ZN( u1_u14_u2_n121 ) , .A2( u1_u14_u2_n177 ) , .A1( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U30 (.A( u1_u14_u2_n132 ) , .ZN( u1_u14_u2_n182 ) );
  INV_X1 u1_u14_u2_U31 (.A( u1_u14_u2_n158 ) , .ZN( u1_u14_u2_n183 ) );
  OAI21_X1 u1_u14_u2_U32 (.A( u1_u14_u2_n156 ) , .B1( u1_u14_u2_n157 ) , .ZN( u1_u14_u2_n158 ) , .B2( u1_u14_u2_n179 ) );
  NOR2_X1 u1_u14_u2_U33 (.ZN( u1_u14_u2_n156 ) , .A1( u1_u14_u2_n166 ) , .A2( u1_u14_u2_n169 ) );
  NOR2_X1 u1_u14_u2_U34 (.A2( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n140 ) );
  NOR2_X1 u1_u14_u2_U35 (.A2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n153 ) , .A1( u1_u14_u2_n156 ) );
  AOI211_X1 u1_u14_u2_U36 (.ZN( u1_u14_u2_n130 ) , .C1( u1_u14_u2_n138 ) , .C2( u1_u14_u2_n179 ) , .B( u1_u14_u2_n96 ) , .A( u1_u14_u2_n97 ) );
  OAI22_X1 u1_u14_u2_U37 (.B1( u1_u14_u2_n133 ) , .A2( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n152 ) , .B2( u1_u14_u2_n168 ) , .ZN( u1_u14_u2_n97 ) );
  OAI221_X1 u1_u14_u2_U38 (.B1( u1_u14_u2_n113 ) , .C1( u1_u14_u2_n132 ) , .A( u1_u14_u2_n149 ) , .B2( u1_u14_u2_n171 ) , .C2( u1_u14_u2_n172 ) , .ZN( u1_u14_u2_n96 ) );
  OAI221_X1 u1_u14_u2_U39 (.A( u1_u14_u2_n115 ) , .C2( u1_u14_u2_n123 ) , .B2( u1_u14_u2_n143 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n163 ) , .C1( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U4 (.A( u1_u14_u2_n134 ) , .ZN( u1_u14_u2_n185 ) );
  OAI21_X1 u1_u14_u2_U40 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n115 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n178 ) );
  OAI221_X1 u1_u14_u2_U41 (.A( u1_u14_u2_n135 ) , .B2( u1_u14_u2_n136 ) , .B1( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n162 ) , .C2( u1_u14_u2_n167 ) , .C1( u1_u14_u2_n185 ) );
  AND3_X1 u1_u14_u2_U42 (.A3( u1_u14_u2_n131 ) , .A2( u1_u14_u2_n132 ) , .A1( u1_u14_u2_n133 ) , .ZN( u1_u14_u2_n136 ) );
  AOI22_X1 u1_u14_u2_U43 (.ZN( u1_u14_u2_n135 ) , .B1( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n156 ) , .B2( u1_u14_u2_n180 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U44 (.ZN( u1_u14_u2_n149 ) , .B1( u1_u14_u2_n173 ) , .B2( u1_u14_u2_n188 ) , .A( u1_u14_u2_n95 ) );
  AND3_X1 u1_u14_u2_U45 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n95 ) );
  OAI21_X1 u1_u14_u2_U46 (.A( u1_u14_u2_n101 ) , .B2( u1_u14_u2_n121 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n164 ) );
  NAND2_X1 u1_u14_u2_U47 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n155 ) );
  NAND2_X1 u1_u14_u2_U48 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n143 ) );
  NAND2_X1 u1_u14_u2_U49 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U5 (.A( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n184 ) );
  NAND2_X1 u1_u14_u2_U50 (.A1( u1_u14_u2_n100 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n132 ) );
  INV_X1 u1_u14_u2_U51 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U52 (.A( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n167 ) );
  OAI21_X1 u1_u14_u2_U53 (.A( u1_u14_u2_n141 ) , .B2( u1_u14_u2_n142 ) , .ZN( u1_u14_u2_n146 ) , .B1( u1_u14_u2_n153 ) );
  OAI21_X1 u1_u14_u2_U54 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n141 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n177 ) );
  NOR3_X1 u1_u14_u2_U55 (.ZN( u1_u14_u2_n142 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n178 ) , .A1( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U56 (.ZN( u1_u14_u2_n187 ) , .A( u1_u14_u2_n99 ) );
  OAI21_X1 u1_u14_u2_U57 (.B1( u1_u14_u2_n137 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n98 ) , .ZN( u1_u14_u2_n99 ) );
  NAND2_X1 u1_u14_u2_U58 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n113 ) );
  NAND2_X1 u1_u14_u2_U59 (.A1( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n131 ) );
  NOR4_X1 u1_u14_u2_U6 (.A4( u1_u14_u2_n124 ) , .A3( u1_u14_u2_n125 ) , .A2( u1_u14_u2_n126 ) , .A1( u1_u14_u2_n127 ) , .ZN( u1_u14_u2_n128 ) );
  NAND2_X1 u1_u14_u2_U60 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n139 ) );
  NAND2_X1 u1_u14_u2_U61 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n133 ) );
  NAND2_X1 u1_u14_u2_U62 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n103 ) , .ZN( u1_u14_u2_n154 ) );
  NAND2_X1 u1_u14_u2_U63 (.A2( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n104 ) , .ZN( u1_u14_u2_n119 ) );
  NAND2_X1 u1_u14_u2_U64 (.A2( u1_u14_u2_n107 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n123 ) );
  NAND2_X1 u1_u14_u2_U65 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n122 ) );
  INV_X1 u1_u14_u2_U66 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n172 ) );
  NAND2_X1 u1_u14_u2_U67 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n102 ) , .ZN( u1_u14_u2_n116 ) );
  NAND2_X1 u1_u14_u2_U68 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n120 ) );
  NAND2_X1 u1_u14_u2_U69 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n117 ) );
  AOI21_X1 u1_u14_u2_U7 (.B2( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n127 ) , .A( u1_u14_u2_n137 ) , .B1( u1_u14_u2_n155 ) );
  NOR2_X1 u1_u14_u2_U70 (.A2( u1_u14_X_16 ) , .ZN( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n166 ) );
  NOR2_X1 u1_u14_u2_U71 (.A2( u1_u14_X_13 ) , .A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n100 ) );
  NOR2_X1 u1_u14_u2_U72 (.A2( u1_u14_X_16 ) , .A1( u1_u14_X_17 ) , .ZN( u1_u14_u2_n138 ) );
  NOR2_X1 u1_u14_u2_U73 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n104 ) );
  NOR2_X1 u1_u14_u2_U74 (.A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n174 ) );
  NOR2_X1 u1_u14_u2_U75 (.A2( u1_u14_X_15 ) , .ZN( u1_u14_u2_n102 ) , .A1( u1_u14_u2_n165 ) );
  NOR2_X1 u1_u14_u2_U76 (.A2( u1_u14_X_17 ) , .ZN( u1_u14_u2_n114 ) , .A1( u1_u14_u2_n169 ) );
  AND2_X1 u1_u14_u2_U77 (.A1( u1_u14_X_15 ) , .ZN( u1_u14_u2_n105 ) , .A2( u1_u14_u2_n165 ) );
  AND2_X1 u1_u14_u2_U78 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n107 ) );
  AND2_X1 u1_u14_u2_U79 (.A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n174 ) );
  AOI21_X1 u1_u14_u2_U8 (.ZN( u1_u14_u2_n124 ) , .B1( u1_u14_u2_n131 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n172 ) );
  AND2_X1 u1_u14_u2_U80 (.A1( u1_u14_X_13 ) , .A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n108 ) );
  INV_X1 u1_u14_u2_U81 (.A( u1_u14_X_16 ) , .ZN( u1_u14_u2_n169 ) );
  INV_X1 u1_u14_u2_U82 (.A( u1_u14_X_17 ) , .ZN( u1_u14_u2_n166 ) );
  INV_X1 u1_u14_u2_U83 (.A( u1_u14_X_13 ) , .ZN( u1_u14_u2_n174 ) );
  INV_X1 u1_u14_u2_U84 (.A( u1_u14_X_18 ) , .ZN( u1_u14_u2_n165 ) );
  NAND4_X1 u1_u14_u2_U85 (.ZN( u1_out14_30 ) , .A4( u1_u14_u2_n147 ) , .A3( u1_u14_u2_n148 ) , .A2( u1_u14_u2_n149 ) , .A1( u1_u14_u2_n187 ) );
  NOR3_X1 u1_u14_u2_U86 (.A3( u1_u14_u2_n144 ) , .A2( u1_u14_u2_n145 ) , .A1( u1_u14_u2_n146 ) , .ZN( u1_u14_u2_n147 ) );
  AOI21_X1 u1_u14_u2_U87 (.B2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n148 ) , .A( u1_u14_u2_n162 ) , .B1( u1_u14_u2_n182 ) );
  NAND4_X1 u1_u14_u2_U88 (.ZN( u1_out14_24 ) , .A4( u1_u14_u2_n111 ) , .A3( u1_u14_u2_n112 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n187 ) );
  AOI221_X1 u1_u14_u2_U89 (.A( u1_u14_u2_n109 ) , .B1( u1_u14_u2_n110 ) , .ZN( u1_u14_u2_n111 ) , .C1( u1_u14_u2_n134 ) , .C2( u1_u14_u2_n170 ) , .B2( u1_u14_u2_n173 ) );
  AOI21_X1 u1_u14_u2_U9 (.B2( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n125 ) , .A( u1_u14_u2_n171 ) , .B1( u1_u14_u2_n184 ) );
  AOI21_X1 u1_u14_u2_U90 (.ZN( u1_u14_u2_n112 ) , .B2( u1_u14_u2_n156 ) , .A( u1_u14_u2_n164 ) , .B1( u1_u14_u2_n181 ) );
  NAND4_X1 u1_u14_u2_U91 (.ZN( u1_out14_16 ) , .A4( u1_u14_u2_n128 ) , .A3( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n186 ) );
  AOI22_X1 u1_u14_u2_U92 (.A2( u1_u14_u2_n118 ) , .ZN( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n140 ) , .B1( u1_u14_u2_n157 ) , .B2( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U93 (.A( u1_u14_u2_n163 ) , .ZN( u1_u14_u2_n186 ) );
  OR4_X1 u1_u14_u2_U94 (.ZN( u1_out14_6 ) , .A4( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n162 ) , .A2( u1_u14_u2_n163 ) , .A1( u1_u14_u2_n164 ) );
  OR3_X1 u1_u14_u2_U95 (.A2( u1_u14_u2_n159 ) , .A1( u1_u14_u2_n160 ) , .ZN( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n183 ) );
  AOI21_X1 u1_u14_u2_U96 (.B2( u1_u14_u2_n154 ) , .B1( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n159 ) , .A( u1_u14_u2_n167 ) );
  NAND3_X1 u1_u14_u2_U97 (.A2( u1_u14_u2_n117 ) , .A1( u1_u14_u2_n122 ) , .A3( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n134 ) );
  NAND3_X1 u1_u14_u2_U98 (.ZN( u1_u14_u2_n110 ) , .A2( u1_u14_u2_n131 ) , .A3( u1_u14_u2_n139 ) , .A1( u1_u14_u2_n154 ) );
  NAND3_X1 u1_u14_u2_U99 (.A2( u1_u14_u2_n100 ) , .ZN( u1_u14_u2_n101 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n114 ) );
  OAI22_X1 u1_u14_u3_U10 (.B1( u1_u14_u3_n113 ) , .A2( u1_u14_u3_n135 ) , .A1( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n164 ) , .ZN( u1_u14_u3_n98 ) );
  OAI211_X1 u1_u14_u3_U11 (.B( u1_u14_u3_n106 ) , .ZN( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n128 ) , .C1( u1_u14_u3_n167 ) , .A( u1_u14_u3_n181 ) );
  AOI221_X1 u1_u14_u3_U12 (.C1( u1_u14_u3_n105 ) , .ZN( u1_u14_u3_n106 ) , .A( u1_u14_u3_n131 ) , .B2( u1_u14_u3_n132 ) , .C2( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n169 ) );
  INV_X1 u1_u14_u3_U13 (.ZN( u1_u14_u3_n181 ) , .A( u1_u14_u3_n98 ) );
  NAND2_X1 u1_u14_u3_U14 (.ZN( u1_u14_u3_n105 ) , .A2( u1_u14_u3_n130 ) , .A1( u1_u14_u3_n155 ) );
  AOI22_X1 u1_u14_u3_U15 (.B1( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n116 ) , .ZN( u1_u14_u3_n123 ) , .B2( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U16 (.ZN( u1_u14_u3_n116 ) , .A2( u1_u14_u3_n151 ) , .A1( u1_u14_u3_n182 ) );
  NOR2_X1 u1_u14_u3_U17 (.ZN( u1_u14_u3_n126 ) , .A2( u1_u14_u3_n150 ) , .A1( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U18 (.ZN( u1_u14_u3_n112 ) , .B2( u1_u14_u3_n146 ) , .B1( u1_u14_u3_n155 ) , .A( u1_u14_u3_n167 ) );
  NAND2_X1 u1_u14_u3_U19 (.A1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n142 ) , .A2( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U20 (.ZN( u1_u14_u3_n132 ) , .A2( u1_u14_u3_n152 ) , .A1( u1_u14_u3_n156 ) );
  AND2_X1 u1_u14_u3_U21 (.A2( u1_u14_u3_n113 ) , .A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n151 ) );
  INV_X1 u1_u14_u3_U22 (.A( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n165 ) );
  INV_X1 u1_u14_u3_U23 (.A( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n170 ) );
  NAND2_X1 u1_u14_u3_U24 (.A1( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .ZN( u1_u14_u3_n140 ) );
  NAND2_X1 u1_u14_u3_U25 (.ZN( u1_u14_u3_n117 ) , .A1( u1_u14_u3_n124 ) , .A2( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U26 (.ZN( u1_u14_u3_n143 ) , .A1( u1_u14_u3_n165 ) , .A2( u1_u14_u3_n167 ) );
  INV_X1 u1_u14_u3_U27 (.A( u1_u14_u3_n130 ) , .ZN( u1_u14_u3_n177 ) );
  INV_X1 u1_u14_u3_U28 (.A( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n176 ) );
  INV_X1 u1_u14_u3_U29 (.A( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n174 ) );
  INV_X1 u1_u14_u3_U3 (.A( u1_u14_u3_n129 ) , .ZN( u1_u14_u3_n183 ) );
  INV_X1 u1_u14_u3_U30 (.A( u1_u14_u3_n139 ) , .ZN( u1_u14_u3_n185 ) );
  NOR2_X1 u1_u14_u3_U31 (.ZN( u1_u14_u3_n135 ) , .A2( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n169 ) );
  OAI222_X1 u1_u14_u3_U32 (.C2( u1_u14_u3_n107 ) , .A2( u1_u14_u3_n108 ) , .B1( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n138 ) , .B2( u1_u14_u3_n146 ) , .C1( u1_u14_u3_n154 ) , .A1( u1_u14_u3_n164 ) );
  NOR4_X1 u1_u14_u3_U33 (.A4( u1_u14_u3_n157 ) , .A3( u1_u14_u3_n158 ) , .A2( u1_u14_u3_n159 ) , .A1( u1_u14_u3_n160 ) , .ZN( u1_u14_u3_n161 ) );
  AOI21_X1 u1_u14_u3_U34 (.B2( u1_u14_u3_n152 ) , .B1( u1_u14_u3_n153 ) , .ZN( u1_u14_u3_n158 ) , .A( u1_u14_u3_n164 ) );
  AOI21_X1 u1_u14_u3_U35 (.A( u1_u14_u3_n154 ) , .B2( u1_u14_u3_n155 ) , .B1( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n157 ) );
  AOI21_X1 u1_u14_u3_U36 (.A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n150 ) , .B1( u1_u14_u3_n151 ) , .ZN( u1_u14_u3_n159 ) );
  AOI211_X1 u1_u14_u3_U37 (.ZN( u1_u14_u3_n109 ) , .A( u1_u14_u3_n119 ) , .C2( u1_u14_u3_n129 ) , .B( u1_u14_u3_n138 ) , .C1( u1_u14_u3_n141 ) );
  AOI211_X1 u1_u14_u3_U38 (.B( u1_u14_u3_n119 ) , .A( u1_u14_u3_n120 ) , .C2( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n122 ) , .C1( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U39 (.A( u1_u14_u3_n156 ) , .ZN( u1_u14_u3_n179 ) );
  INV_X1 u1_u14_u3_U4 (.A( u1_u14_u3_n140 ) , .ZN( u1_u14_u3_n182 ) );
  OAI22_X1 u1_u14_u3_U40 (.B1( u1_u14_u3_n118 ) , .ZN( u1_u14_u3_n120 ) , .A1( u1_u14_u3_n135 ) , .B2( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n178 ) );
  AND3_X1 u1_u14_u3_U41 (.ZN( u1_u14_u3_n118 ) , .A2( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n144 ) , .A3( u1_u14_u3_n152 ) );
  INV_X1 u1_u14_u3_U42 (.A( u1_u14_u3_n121 ) , .ZN( u1_u14_u3_n164 ) );
  NAND2_X1 u1_u14_u3_U43 (.ZN( u1_u14_u3_n133 ) , .A1( u1_u14_u3_n154 ) , .A2( u1_u14_u3_n164 ) );
  OAI211_X1 u1_u14_u3_U44 (.B( u1_u14_u3_n127 ) , .ZN( u1_u14_u3_n139 ) , .C1( u1_u14_u3_n150 ) , .C2( u1_u14_u3_n154 ) , .A( u1_u14_u3_n184 ) );
  INV_X1 u1_u14_u3_U45 (.A( u1_u14_u3_n125 ) , .ZN( u1_u14_u3_n184 ) );
  AOI221_X1 u1_u14_u3_U46 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n127 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n169 ) , .B2( u1_u14_u3_n170 ) , .B1( u1_u14_u3_n174 ) );
  OAI22_X1 u1_u14_u3_U47 (.A1( u1_u14_u3_n124 ) , .ZN( u1_u14_u3_n125 ) , .B2( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n165 ) , .B1( u1_u14_u3_n167 ) );
  NOR2_X1 u1_u14_u3_U48 (.A1( u1_u14_u3_n113 ) , .ZN( u1_u14_u3_n131 ) , .A2( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U49 (.A1( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n150 ) , .A2( u1_u14_u3_n99 ) );
  INV_X1 u1_u14_u3_U5 (.A( u1_u14_u3_n117 ) , .ZN( u1_u14_u3_n178 ) );
  NAND2_X1 u1_u14_u3_U50 (.A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n155 ) , .A1( u1_u14_u3_n97 ) );
  INV_X1 u1_u14_u3_U51 (.A( u1_u14_u3_n141 ) , .ZN( u1_u14_u3_n167 ) );
  AOI21_X1 u1_u14_u3_U52 (.B2( u1_u14_u3_n114 ) , .B1( u1_u14_u3_n146 ) , .A( u1_u14_u3_n154 ) , .ZN( u1_u14_u3_n94 ) );
  AOI21_X1 u1_u14_u3_U53 (.ZN( u1_u14_u3_n110 ) , .B2( u1_u14_u3_n142 ) , .B1( u1_u14_u3_n186 ) , .A( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U54 (.A( u1_u14_u3_n145 ) , .ZN( u1_u14_u3_n186 ) );
  AOI21_X1 u1_u14_u3_U55 (.B1( u1_u14_u3_n124 ) , .A( u1_u14_u3_n149 ) , .B2( u1_u14_u3_n155 ) , .ZN( u1_u14_u3_n95 ) );
  INV_X1 u1_u14_u3_U56 (.A( u1_u14_u3_n149 ) , .ZN( u1_u14_u3_n169 ) );
  NAND2_X1 u1_u14_u3_U57 (.ZN( u1_u14_u3_n124 ) , .A1( u1_u14_u3_n96 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U58 (.A2( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n146 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U59 (.A1( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n145 ) , .A2( u1_u14_u3_n99 ) );
  AOI221_X1 u1_u14_u3_U6 (.A( u1_u14_u3_n131 ) , .C2( u1_u14_u3_n132 ) , .C1( u1_u14_u3_n133 ) , .ZN( u1_u14_u3_n134 ) , .B1( u1_u14_u3_n143 ) , .B2( u1_u14_u3_n177 ) );
  NAND2_X1 u1_u14_u3_U60 (.A1( u1_u14_u3_n100 ) , .ZN( u1_u14_u3_n156 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U61 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n148 ) );
  NAND2_X1 u1_u14_u3_U62 (.A1( u1_u14_u3_n100 ) , .A2( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n128 ) );
  NAND2_X1 u1_u14_u3_U63 (.A2( u1_u14_u3_n101 ) , .A1( u1_u14_u3_n102 ) , .ZN( u1_u14_u3_n152 ) );
  NAND2_X1 u1_u14_u3_U64 (.A2( u1_u14_u3_n101 ) , .ZN( u1_u14_u3_n114 ) , .A1( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U65 (.ZN( u1_u14_u3_n107 ) , .A1( u1_u14_u3_n97 ) , .A2( u1_u14_u3_n99 ) );
  NAND2_X1 u1_u14_u3_U66 (.A2( u1_u14_u3_n100 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n113 ) );
  NAND2_X1 u1_u14_u3_U67 (.A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n153 ) , .A2( u1_u14_u3_n97 ) );
  NAND2_X1 u1_u14_u3_U68 (.A2( u1_u14_u3_n103 ) , .A1( u1_u14_u3_n104 ) , .ZN( u1_u14_u3_n130 ) );
  NAND2_X1 u1_u14_u3_U69 (.A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n96 ) );
  OAI22_X1 u1_u14_u3_U7 (.B2( u1_u14_u3_n147 ) , .A2( u1_u14_u3_n148 ) , .ZN( u1_u14_u3_n160 ) , .B1( u1_u14_u3_n165 ) , .A1( u1_u14_u3_n168 ) );
  NAND2_X1 u1_u14_u3_U70 (.A1( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n103 ) , .ZN( u1_u14_u3_n108 ) );
  NOR2_X1 u1_u14_u3_U71 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n99 ) );
  NOR2_X1 u1_u14_u3_U72 (.A2( u1_u14_X_21 ) , .A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n103 ) );
  NOR2_X1 u1_u14_u3_U73 (.A2( u1_u14_X_24 ) , .A1( u1_u14_u3_n171 ) , .ZN( u1_u14_u3_n97 ) );
  NOR2_X1 u1_u14_u3_U74 (.A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n141 ) , .A1( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U75 (.A2( u1_u14_X_19 ) , .A1( u1_u14_u3_n172 ) , .ZN( u1_u14_u3_n96 ) );
  NAND2_X1 u1_u14_u3_U76 (.A1( u1_u14_X_22 ) , .A2( u1_u14_X_23 ) , .ZN( u1_u14_u3_n154 ) );
  NAND2_X1 u1_u14_u3_U77 (.A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n149 ) , .A2( u1_u14_u3_n166 ) );
  NOR2_X1 u1_u14_u3_U78 (.A2( u1_u14_X_22 ) , .A1( u1_u14_X_23 ) , .ZN( u1_u14_u3_n121 ) );
  AND2_X1 u1_u14_u3_U79 (.A1( u1_u14_X_24 ) , .ZN( u1_u14_u3_n101 ) , .A2( u1_u14_u3_n171 ) );
  AND3_X1 u1_u14_u3_U8 (.A3( u1_u14_u3_n144 ) , .A2( u1_u14_u3_n145 ) , .A1( u1_u14_u3_n146 ) , .ZN( u1_u14_u3_n147 ) );
  AND2_X1 u1_u14_u3_U80 (.A1( u1_u14_X_19 ) , .ZN( u1_u14_u3_n102 ) , .A2( u1_u14_u3_n172 ) );
  AND2_X1 u1_u14_u3_U81 (.A1( u1_u14_X_21 ) , .A2( u1_u14_X_24 ) , .ZN( u1_u14_u3_n100 ) );
  AND2_X1 u1_u14_u3_U82 (.A2( u1_u14_X_19 ) , .A1( u1_u14_X_20 ) , .ZN( u1_u14_u3_n104 ) );
  INV_X1 u1_u14_u3_U83 (.A( u1_u14_X_22 ) , .ZN( u1_u14_u3_n166 ) );
  INV_X1 u1_u14_u3_U84 (.A( u1_u14_X_21 ) , .ZN( u1_u14_u3_n171 ) );
  INV_X1 u1_u14_u3_U85 (.A( u1_u14_X_20 ) , .ZN( u1_u14_u3_n172 ) );
  NAND4_X1 u1_u14_u3_U86 (.ZN( u1_out14_26 ) , .A4( u1_u14_u3_n109 ) , .A3( u1_u14_u3_n110 ) , .A2( u1_u14_u3_n111 ) , .A1( u1_u14_u3_n173 ) );
  INV_X1 u1_u14_u3_U87 (.ZN( u1_u14_u3_n173 ) , .A( u1_u14_u3_n94 ) );
  OAI21_X1 u1_u14_u3_U88 (.ZN( u1_u14_u3_n111 ) , .B2( u1_u14_u3_n117 ) , .A( u1_u14_u3_n133 ) , .B1( u1_u14_u3_n176 ) );
  NAND4_X1 u1_u14_u3_U89 (.ZN( u1_out14_20 ) , .A4( u1_u14_u3_n122 ) , .A3( u1_u14_u3_n123 ) , .A1( u1_u14_u3_n175 ) , .A2( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U9 (.A( u1_u14_u3_n143 ) , .ZN( u1_u14_u3_n168 ) );
  INV_X1 u1_u14_u3_U90 (.A( u1_u14_u3_n126 ) , .ZN( u1_u14_u3_n180 ) );
  INV_X1 u1_u14_u3_U91 (.A( u1_u14_u3_n112 ) , .ZN( u1_u14_u3_n175 ) );
  NAND4_X1 u1_u14_u3_U92 (.ZN( u1_out14_1 ) , .A4( u1_u14_u3_n161 ) , .A3( u1_u14_u3_n162 ) , .A2( u1_u14_u3_n163 ) , .A1( u1_u14_u3_n185 ) );
  NAND2_X1 u1_u14_u3_U93 (.ZN( u1_u14_u3_n163 ) , .A2( u1_u14_u3_n170 ) , .A1( u1_u14_u3_n176 ) );
  AOI22_X1 u1_u14_u3_U94 (.B2( u1_u14_u3_n140 ) , .B1( u1_u14_u3_n141 ) , .A2( u1_u14_u3_n142 ) , .ZN( u1_u14_u3_n162 ) , .A1( u1_u14_u3_n177 ) );
  OR4_X1 u1_u14_u3_U95 (.ZN( u1_out14_10 ) , .A4( u1_u14_u3_n136 ) , .A3( u1_u14_u3_n137 ) , .A1( u1_u14_u3_n138 ) , .A2( u1_u14_u3_n139 ) );
  OAI222_X1 u1_u14_u3_U96 (.C1( u1_u14_u3_n128 ) , .ZN( u1_u14_u3_n137 ) , .B1( u1_u14_u3_n148 ) , .A2( u1_u14_u3_n150 ) , .B2( u1_u14_u3_n154 ) , .C2( u1_u14_u3_n164 ) , .A1( u1_u14_u3_n167 ) );
  OAI221_X1 u1_u14_u3_U97 (.A( u1_u14_u3_n134 ) , .B2( u1_u14_u3_n135 ) , .ZN( u1_u14_u3_n136 ) , .C1( u1_u14_u3_n149 ) , .B1( u1_u14_u3_n151 ) , .C2( u1_u14_u3_n183 ) );
  NAND3_X1 u1_u14_u3_U98 (.A1( u1_u14_u3_n114 ) , .ZN( u1_u14_u3_n115 ) , .A2( u1_u14_u3_n145 ) , .A3( u1_u14_u3_n153 ) );
  NAND3_X1 u1_u14_u3_U99 (.ZN( u1_u14_u3_n129 ) , .A2( u1_u14_u3_n144 ) , .A1( u1_u14_u3_n153 ) , .A3( u1_u14_u3_n182 ) );
  OAI22_X1 u1_u14_u4_U10 (.B2( u1_u14_u4_n135 ) , .ZN( u1_u14_u4_n137 ) , .B1( u1_u14_u4_n153 ) , .A1( u1_u14_u4_n155 ) , .A2( u1_u14_u4_n171 ) );
  AND3_X1 u1_u14_u4_U11 (.A2( u1_u14_u4_n134 ) , .ZN( u1_u14_u4_n135 ) , .A3( u1_u14_u4_n145 ) , .A1( u1_u14_u4_n157 ) );
  NAND2_X1 u1_u14_u4_U12 (.ZN( u1_u14_u4_n132 ) , .A2( u1_u14_u4_n170 ) , .A1( u1_u14_u4_n173 ) );
  AOI21_X1 u1_u14_u4_U13 (.B2( u1_u14_u4_n160 ) , .B1( u1_u14_u4_n161 ) , .ZN( u1_u14_u4_n162 ) , .A( u1_u14_u4_n170 ) );
  AOI21_X1 u1_u14_u4_U14 (.ZN( u1_u14_u4_n107 ) , .B2( u1_u14_u4_n143 ) , .A( u1_u14_u4_n174 ) , .B1( u1_u14_u4_n184 ) );
  AOI21_X1 u1_u14_u4_U15 (.B2( u1_u14_u4_n158 ) , .B1( u1_u14_u4_n159 ) , .ZN( u1_u14_u4_n163 ) , .A( u1_u14_u4_n174 ) );
  AOI21_X1 u1_u14_u4_U16 (.A( u1_u14_u4_n153 ) , .B2( u1_u14_u4_n154 ) , .B1( u1_u14_u4_n155 ) , .ZN( u1_u14_u4_n165 ) );
  AOI21_X1 u1_u14_u4_U17 (.A( u1_u14_u4_n156 ) , .B2( u1_u14_u4_n157 ) , .ZN( u1_u14_u4_n164 ) , .B1( u1_u14_u4_n184 ) );
  INV_X1 u1_u14_u4_U18 (.A( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n170 ) );
  AND2_X1 u1_u14_u4_U19 (.A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n155 ) , .A1( u1_u14_u4_n160 ) );
  INV_X1 u1_u14_u4_U20 (.A( u1_u14_u4_n156 ) , .ZN( u1_u14_u4_n175 ) );
  NAND2_X1 u1_u14_u4_U21 (.A2( u1_u14_u4_n118 ) , .ZN( u1_u14_u4_n131 ) , .A1( u1_u14_u4_n147 ) );
  NAND2_X1 u1_u14_u4_U22 (.A1( u1_u14_u4_n119 ) , .A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n130 ) );
  NAND2_X1 u1_u14_u4_U23 (.ZN( u1_u14_u4_n117 ) , .A2( u1_u14_u4_n118 ) , .A1( u1_u14_u4_n148 ) );
  NAND2_X1 u1_u14_u4_U24 (.ZN( u1_u14_u4_n129 ) , .A1( u1_u14_u4_n134 ) , .A2( u1_u14_u4_n148 ) );
  AND3_X1 u1_u14_u4_U25 (.A1( u1_u14_u4_n119 ) , .A2( u1_u14_u4_n143 ) , .A3( u1_u14_u4_n154 ) , .ZN( u1_u14_u4_n161 ) );
  AND2_X1 u1_u14_u4_U26 (.A1( u1_u14_u4_n145 ) , .A2( u1_u14_u4_n147 ) , .ZN( u1_u14_u4_n159 ) );
  OR3_X1 u1_u14_u4_U27 (.A3( u1_u14_u4_n114 ) , .A2( u1_u14_u4_n115 ) , .A1( u1_u14_u4_n116 ) , .ZN( u1_u14_u4_n136 ) );
  AOI21_X1 u1_u14_u4_U28 (.A( u1_u14_u4_n113 ) , .ZN( u1_u14_u4_n116 ) , .B2( u1_u14_u4_n173 ) , .B1( u1_u14_u4_n174 ) );
  AOI21_X1 u1_u14_u4_U29 (.ZN( u1_u14_u4_n115 ) , .B2( u1_u14_u4_n145 ) , .B1( u1_u14_u4_n146 ) , .A( u1_u14_u4_n156 ) );
  NOR2_X1 u1_u14_u4_U3 (.ZN( u1_u14_u4_n121 ) , .A1( u1_u14_u4_n181 ) , .A2( u1_u14_u4_n182 ) );
  OAI22_X1 u1_u14_u4_U30 (.ZN( u1_u14_u4_n114 ) , .A2( u1_u14_u4_n121 ) , .B1( u1_u14_u4_n160 ) , .B2( u1_u14_u4_n170 ) , .A1( u1_u14_u4_n171 ) );
  INV_X1 u1_u14_u4_U31 (.A( u1_u14_u4_n158 ) , .ZN( u1_u14_u4_n182 ) );
  INV_X1 u1_u14_u4_U32 (.ZN( u1_u14_u4_n181 ) , .A( u1_u14_u4_n96 ) );
  INV_X1 u1_u14_u4_U33 (.A( u1_u14_u4_n144 ) , .ZN( u1_u14_u4_n179 ) );
  INV_X1 u1_u14_u4_U34 (.A( u1_u14_u4_n157 ) , .ZN( u1_u14_u4_n178 ) );
  NAND2_X1 u1_u14_u4_U35 (.A2( u1_u14_u4_n154 ) , .A1( u1_u14_u4_n96 ) , .ZN( u1_u14_u4_n97 ) );
  INV_X1 u1_u14_u4_U36 (.ZN( u1_u14_u4_n186 ) , .A( u1_u14_u4_n95 ) );
  OAI221_X1 u1_u14_u4_U37 (.C1( u1_u14_u4_n134 ) , .B1( u1_u14_u4_n158 ) , .B2( u1_u14_u4_n171 ) , .C2( u1_u14_u4_n173 ) , .A( u1_u14_u4_n94 ) , .ZN( u1_u14_u4_n95 ) );
  AOI222_X1 u1_u14_u4_U38 (.B2( u1_u14_u4_n132 ) , .A1( u1_u14_u4_n138 ) , .C2( u1_u14_u4_n175 ) , .A2( u1_u14_u4_n179 ) , .C1( u1_u14_u4_n181 ) , .B1( u1_u14_u4_n185 ) , .ZN( u1_u14_u4_n94 ) );
  INV_X1 u1_u14_u4_U39 (.A( u1_u14_u4_n113 ) , .ZN( u1_u14_u4_n185 ) );
  INV_X1 u1_u14_u4_U4 (.A( u1_u14_u4_n117 ) , .ZN( u1_u14_u4_n184 ) );
  INV_X1 u1_u14_u4_U40 (.A( u1_u14_u4_n143 ) , .ZN( u1_u14_u4_n183 ) );
  NOR2_X1 u1_u14_u4_U41 (.ZN( u1_u14_u4_n138 ) , .A1( u1_u14_u4_n168 ) , .A2( u1_u14_u4_n169 ) );
  NOR2_X1 u1_u14_u4_U42 (.A1( u1_u14_u4_n150 ) , .A2( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n153 ) );
  NOR2_X1 u1_u14_u4_U43 (.A2( u1_u14_u4_n128 ) , .A1( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n156 ) );
  AOI22_X1 u1_u14_u4_U44 (.B2( u1_u14_u4_n122 ) , .A1( u1_u14_u4_n123 ) , .ZN( u1_u14_u4_n124 ) , .B1( u1_u14_u4_n128 ) , .A2( u1_u14_u4_n172 ) );
  INV_X1 u1_u14_u4_U45 (.A( u1_u14_u4_n153 ) , .ZN( u1_u14_u4_n172 ) );
  NAND2_X1 u1_u14_u4_U46 (.A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n123 ) , .A1( u1_u14_u4_n161 ) );
  AOI22_X1 u1_u14_u4_U47 (.B2( u1_u14_u4_n132 ) , .A2( u1_u14_u4_n133 ) , .ZN( u1_u14_u4_n140 ) , .A1( u1_u14_u4_n150 ) , .B1( u1_u14_u4_n179 ) );
  NAND2_X1 u1_u14_u4_U48 (.ZN( u1_u14_u4_n133 ) , .A2( u1_u14_u4_n146 ) , .A1( u1_u14_u4_n154 ) );
  NAND2_X1 u1_u14_u4_U49 (.A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n154 ) , .A2( u1_u14_u4_n98 ) );
  NOR4_X1 u1_u14_u4_U5 (.A4( u1_u14_u4_n106 ) , .A3( u1_u14_u4_n107 ) , .A2( u1_u14_u4_n108 ) , .A1( u1_u14_u4_n109 ) , .ZN( u1_u14_u4_n110 ) );
  NAND2_X1 u1_u14_u4_U50 (.A1( u1_u14_u4_n101 ) , .ZN( u1_u14_u4_n158 ) , .A2( u1_u14_u4_n99 ) );
  AOI21_X1 u1_u14_u4_U51 (.ZN( u1_u14_u4_n127 ) , .A( u1_u14_u4_n136 ) , .B2( u1_u14_u4_n150 ) , .B1( u1_u14_u4_n180 ) );
  INV_X1 u1_u14_u4_U52 (.A( u1_u14_u4_n160 ) , .ZN( u1_u14_u4_n180 ) );
  NAND2_X1 u1_u14_u4_U53 (.A2( u1_u14_u4_n104 ) , .A1( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n146 ) );
  NAND2_X1 u1_u14_u4_U54 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n160 ) );
  NAND2_X1 u1_u14_u4_U55 (.ZN( u1_u14_u4_n134 ) , .A1( u1_u14_u4_n98 ) , .A2( u1_u14_u4_n99 ) );
  NAND2_X1 u1_u14_u4_U56 (.A1( u1_u14_u4_n103 ) , .A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n143 ) );
  NAND2_X1 u1_u14_u4_U57 (.A2( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n145 ) , .A1( u1_u14_u4_n98 ) );
  NAND2_X1 u1_u14_u4_U58 (.A1( u1_u14_u4_n100 ) , .A2( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n120 ) );
  NAND2_X1 u1_u14_u4_U59 (.A1( u1_u14_u4_n102 ) , .A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n148 ) );
  AOI21_X1 u1_u14_u4_U6 (.ZN( u1_u14_u4_n106 ) , .B2( u1_u14_u4_n146 ) , .B1( u1_u14_u4_n158 ) , .A( u1_u14_u4_n170 ) );
  NAND2_X1 u1_u14_u4_U60 (.A2( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n157 ) );
  INV_X1 u1_u14_u4_U61 (.A( u1_u14_u4_n150 ) , .ZN( u1_u14_u4_n173 ) );
  INV_X1 u1_u14_u4_U62 (.A( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n171 ) );
  NAND2_X1 u1_u14_u4_U63 (.A1( u1_u14_u4_n100 ) , .ZN( u1_u14_u4_n118 ) , .A2( u1_u14_u4_n99 ) );
  NAND2_X1 u1_u14_u4_U64 (.A2( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n144 ) );
  NAND2_X1 u1_u14_u4_U65 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n96 ) );
  INV_X1 u1_u14_u4_U66 (.A( u1_u14_u4_n128 ) , .ZN( u1_u14_u4_n174 ) );
  NAND2_X1 u1_u14_u4_U67 (.A2( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n119 ) , .A1( u1_u14_u4_n98 ) );
  NAND2_X1 u1_u14_u4_U68 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n147 ) );
  NAND2_X1 u1_u14_u4_U69 (.A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n113 ) , .A1( u1_u14_u4_n99 ) );
  AOI21_X1 u1_u14_u4_U7 (.ZN( u1_u14_u4_n108 ) , .B2( u1_u14_u4_n134 ) , .B1( u1_u14_u4_n155 ) , .A( u1_u14_u4_n156 ) );
  NOR2_X1 u1_u14_u4_U70 (.A2( u1_u14_X_28 ) , .ZN( u1_u14_u4_n150 ) , .A1( u1_u14_u4_n168 ) );
  NOR2_X1 u1_u14_u4_U71 (.A2( u1_u14_X_29 ) , .ZN( u1_u14_u4_n152 ) , .A1( u1_u14_u4_n169 ) );
  NOR2_X1 u1_u14_u4_U72 (.A2( u1_u14_X_30 ) , .ZN( u1_u14_u4_n105 ) , .A1( u1_u14_u4_n176 ) );
  NOR2_X1 u1_u14_u4_U73 (.A2( u1_u14_X_26 ) , .ZN( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n177 ) );
  NOR2_X1 u1_u14_u4_U74 (.A2( u1_u14_X_28 ) , .A1( u1_u14_X_29 ) , .ZN( u1_u14_u4_n128 ) );
  NOR2_X1 u1_u14_u4_U75 (.A2( u1_u14_X_27 ) , .A1( u1_u14_X_30 ) , .ZN( u1_u14_u4_n102 ) );
  NOR2_X1 u1_u14_u4_U76 (.A2( u1_u14_X_25 ) , .A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n98 ) );
  AND2_X1 u1_u14_u4_U77 (.A2( u1_u14_X_25 ) , .A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n104 ) );
  AND2_X1 u1_u14_u4_U78 (.A1( u1_u14_X_30 ) , .A2( u1_u14_u4_n176 ) , .ZN( u1_u14_u4_n99 ) );
  AND2_X1 u1_u14_u4_U79 (.A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n101 ) , .A2( u1_u14_u4_n177 ) );
  AOI21_X1 u1_u14_u4_U8 (.ZN( u1_u14_u4_n109 ) , .A( u1_u14_u4_n153 ) , .B1( u1_u14_u4_n159 ) , .B2( u1_u14_u4_n184 ) );
  AND2_X1 u1_u14_u4_U80 (.A1( u1_u14_X_27 ) , .A2( u1_u14_X_30 ) , .ZN( u1_u14_u4_n103 ) );
  INV_X1 u1_u14_u4_U81 (.A( u1_u14_X_28 ) , .ZN( u1_u14_u4_n169 ) );
  INV_X1 u1_u14_u4_U82 (.A( u1_u14_X_29 ) , .ZN( u1_u14_u4_n168 ) );
  INV_X1 u1_u14_u4_U83 (.A( u1_u14_X_25 ) , .ZN( u1_u14_u4_n177 ) );
  INV_X1 u1_u14_u4_U84 (.A( u1_u14_X_27 ) , .ZN( u1_u14_u4_n176 ) );
  NAND4_X1 u1_u14_u4_U85 (.ZN( u1_out14_25 ) , .A4( u1_u14_u4_n139 ) , .A3( u1_u14_u4_n140 ) , .A2( u1_u14_u4_n141 ) , .A1( u1_u14_u4_n142 ) );
  OAI21_X1 u1_u14_u4_U86 (.A( u1_u14_u4_n128 ) , .B2( u1_u14_u4_n129 ) , .B1( u1_u14_u4_n130 ) , .ZN( u1_u14_u4_n142 ) );
  OAI21_X1 u1_u14_u4_U87 (.B2( u1_u14_u4_n131 ) , .ZN( u1_u14_u4_n141 ) , .A( u1_u14_u4_n175 ) , .B1( u1_u14_u4_n183 ) );
  NAND4_X1 u1_u14_u4_U88 (.ZN( u1_out14_14 ) , .A4( u1_u14_u4_n124 ) , .A3( u1_u14_u4_n125 ) , .A2( u1_u14_u4_n126 ) , .A1( u1_u14_u4_n127 ) );
  AOI22_X1 u1_u14_u4_U89 (.B2( u1_u14_u4_n117 ) , .ZN( u1_u14_u4_n126 ) , .A1( u1_u14_u4_n129 ) , .B1( u1_u14_u4_n152 ) , .A2( u1_u14_u4_n175 ) );
  AOI211_X1 u1_u14_u4_U9 (.B( u1_u14_u4_n136 ) , .A( u1_u14_u4_n137 ) , .C2( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n139 ) , .C1( u1_u14_u4_n182 ) );
  AOI22_X1 u1_u14_u4_U90 (.ZN( u1_u14_u4_n125 ) , .B2( u1_u14_u4_n131 ) , .A2( u1_u14_u4_n132 ) , .B1( u1_u14_u4_n138 ) , .A1( u1_u14_u4_n178 ) );
  NAND4_X1 u1_u14_u4_U91 (.ZN( u1_out14_8 ) , .A4( u1_u14_u4_n110 ) , .A3( u1_u14_u4_n111 ) , .A2( u1_u14_u4_n112 ) , .A1( u1_u14_u4_n186 ) );
  NAND2_X1 u1_u14_u4_U92 (.ZN( u1_u14_u4_n112 ) , .A2( u1_u14_u4_n130 ) , .A1( u1_u14_u4_n150 ) );
  AOI22_X1 u1_u14_u4_U93 (.ZN( u1_u14_u4_n111 ) , .B2( u1_u14_u4_n132 ) , .A1( u1_u14_u4_n152 ) , .B1( u1_u14_u4_n178 ) , .A2( u1_u14_u4_n97 ) );
  AOI22_X1 u1_u14_u4_U94 (.B2( u1_u14_u4_n149 ) , .B1( u1_u14_u4_n150 ) , .A2( u1_u14_u4_n151 ) , .A1( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n167 ) );
  NOR4_X1 u1_u14_u4_U95 (.A4( u1_u14_u4_n162 ) , .A3( u1_u14_u4_n163 ) , .A2( u1_u14_u4_n164 ) , .A1( u1_u14_u4_n165 ) , .ZN( u1_u14_u4_n166 ) );
  NAND3_X1 u1_u14_u4_U96 (.ZN( u1_out14_3 ) , .A3( u1_u14_u4_n166 ) , .A1( u1_u14_u4_n167 ) , .A2( u1_u14_u4_n186 ) );
  NAND3_X1 u1_u14_u4_U97 (.A3( u1_u14_u4_n146 ) , .A2( u1_u14_u4_n147 ) , .A1( u1_u14_u4_n148 ) , .ZN( u1_u14_u4_n149 ) );
  NAND3_X1 u1_u14_u4_U98 (.A3( u1_u14_u4_n143 ) , .A2( u1_u14_u4_n144 ) , .A1( u1_u14_u4_n145 ) , .ZN( u1_u14_u4_n151 ) );
  NAND3_X1 u1_u14_u4_U99 (.A3( u1_u14_u4_n121 ) , .ZN( u1_u14_u4_n122 ) , .A2( u1_u14_u4_n144 ) , .A1( u1_u14_u4_n154 ) );
  INV_X1 u1_u14_u5_U10 (.A( u1_u14_u5_n121 ) , .ZN( u1_u14_u5_n177 ) );
  NOR3_X1 u1_u14_u5_U100 (.A3( u1_u14_u5_n141 ) , .A1( u1_u14_u5_n142 ) , .ZN( u1_u14_u5_n143 ) , .A2( u1_u14_u5_n191 ) );
  NAND4_X1 u1_u14_u5_U101 (.ZN( u1_out14_4 ) , .A4( u1_u14_u5_n112 ) , .A2( u1_u14_u5_n113 ) , .A1( u1_u14_u5_n114 ) , .A3( u1_u14_u5_n195 ) );
  AOI211_X1 u1_u14_u5_U102 (.A( u1_u14_u5_n110 ) , .C1( u1_u14_u5_n111 ) , .ZN( u1_u14_u5_n112 ) , .B( u1_u14_u5_n118 ) , .C2( u1_u14_u5_n177 ) );
  AOI222_X1 u1_u14_u5_U103 (.ZN( u1_u14_u5_n113 ) , .A1( u1_u14_u5_n131 ) , .C1( u1_u14_u5_n148 ) , .B2( u1_u14_u5_n174 ) , .C2( u1_u14_u5_n178 ) , .A2( u1_u14_u5_n179 ) , .B1( u1_u14_u5_n99 ) );
  NAND3_X1 u1_u14_u5_U104 (.A2( u1_u14_u5_n154 ) , .A3( u1_u14_u5_n158 ) , .A1( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n99 ) );
  NOR2_X1 u1_u14_u5_U11 (.ZN( u1_u14_u5_n160 ) , .A2( u1_u14_u5_n173 ) , .A1( u1_u14_u5_n177 ) );
  INV_X1 u1_u14_u5_U12 (.A( u1_u14_u5_n150 ) , .ZN( u1_u14_u5_n174 ) );
  AOI21_X1 u1_u14_u5_U13 (.A( u1_u14_u5_n160 ) , .B2( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n162 ) , .B1( u1_u14_u5_n192 ) );
  INV_X1 u1_u14_u5_U14 (.A( u1_u14_u5_n159 ) , .ZN( u1_u14_u5_n192 ) );
  AOI21_X1 u1_u14_u5_U15 (.A( u1_u14_u5_n156 ) , .B2( u1_u14_u5_n157 ) , .B1( u1_u14_u5_n158 ) , .ZN( u1_u14_u5_n163 ) );
  AOI21_X1 u1_u14_u5_U16 (.B2( u1_u14_u5_n139 ) , .B1( u1_u14_u5_n140 ) , .ZN( u1_u14_u5_n141 ) , .A( u1_u14_u5_n150 ) );
  OAI21_X1 u1_u14_u5_U17 (.A( u1_u14_u5_n133 ) , .B2( u1_u14_u5_n134 ) , .B1( u1_u14_u5_n135 ) , .ZN( u1_u14_u5_n142 ) );
  OAI21_X1 u1_u14_u5_U18 (.ZN( u1_u14_u5_n133 ) , .B2( u1_u14_u5_n147 ) , .A( u1_u14_u5_n173 ) , .B1( u1_u14_u5_n188 ) );
  NAND2_X1 u1_u14_u5_U19 (.A2( u1_u14_u5_n119 ) , .A1( u1_u14_u5_n123 ) , .ZN( u1_u14_u5_n137 ) );
  INV_X1 u1_u14_u5_U20 (.A( u1_u14_u5_n155 ) , .ZN( u1_u14_u5_n194 ) );
  NAND2_X1 u1_u14_u5_U21 (.A1( u1_u14_u5_n121 ) , .ZN( u1_u14_u5_n132 ) , .A2( u1_u14_u5_n172 ) );
  NAND2_X1 u1_u14_u5_U22 (.A2( u1_u14_u5_n122 ) , .ZN( u1_u14_u5_n136 ) , .A1( u1_u14_u5_n154 ) );
  NAND2_X1 u1_u14_u5_U23 (.A2( u1_u14_u5_n119 ) , .A1( u1_u14_u5_n120 ) , .ZN( u1_u14_u5_n159 ) );
  INV_X1 u1_u14_u5_U24 (.A( u1_u14_u5_n156 ) , .ZN( u1_u14_u5_n175 ) );
  INV_X1 u1_u14_u5_U25 (.A( u1_u14_u5_n158 ) , .ZN( u1_u14_u5_n188 ) );
  INV_X1 u1_u14_u5_U26 (.A( u1_u14_u5_n152 ) , .ZN( u1_u14_u5_n179 ) );
  INV_X1 u1_u14_u5_U27 (.A( u1_u14_u5_n140 ) , .ZN( u1_u14_u5_n182 ) );
  INV_X1 u1_u14_u5_U28 (.A( u1_u14_u5_n151 ) , .ZN( u1_u14_u5_n183 ) );
  INV_X1 u1_u14_u5_U29 (.A( u1_u14_u5_n123 ) , .ZN( u1_u14_u5_n185 ) );
  NOR2_X1 u1_u14_u5_U3 (.ZN( u1_u14_u5_n134 ) , .A1( u1_u14_u5_n183 ) , .A2( u1_u14_u5_n190 ) );
  INV_X1 u1_u14_u5_U30 (.A( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n184 ) );
  INV_X1 u1_u14_u5_U31 (.A( u1_u14_u5_n139 ) , .ZN( u1_u14_u5_n189 ) );
  INV_X1 u1_u14_u5_U32 (.A( u1_u14_u5_n157 ) , .ZN( u1_u14_u5_n190 ) );
  INV_X1 u1_u14_u5_U33 (.A( u1_u14_u5_n120 ) , .ZN( u1_u14_u5_n193 ) );
  NAND2_X1 u1_u14_u5_U34 (.ZN( u1_u14_u5_n111 ) , .A1( u1_u14_u5_n140 ) , .A2( u1_u14_u5_n155 ) );
  INV_X1 u1_u14_u5_U35 (.A( u1_u14_u5_n117 ) , .ZN( u1_u14_u5_n196 ) );
  OAI221_X1 u1_u14_u5_U36 (.A( u1_u14_u5_n116 ) , .ZN( u1_u14_u5_n117 ) , .B2( u1_u14_u5_n119 ) , .C1( u1_u14_u5_n153 ) , .C2( u1_u14_u5_n158 ) , .B1( u1_u14_u5_n172 ) );
  AOI222_X1 u1_u14_u5_U37 (.ZN( u1_u14_u5_n116 ) , .B2( u1_u14_u5_n145 ) , .C1( u1_u14_u5_n148 ) , .A2( u1_u14_u5_n174 ) , .C2( u1_u14_u5_n177 ) , .B1( u1_u14_u5_n187 ) , .A1( u1_u14_u5_n193 ) );
  INV_X1 u1_u14_u5_U38 (.A( u1_u14_u5_n115 ) , .ZN( u1_u14_u5_n187 ) );
  NOR2_X1 u1_u14_u5_U39 (.ZN( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n170 ) , .A2( u1_u14_u5_n180 ) );
  INV_X1 u1_u14_u5_U4 (.A( u1_u14_u5_n138 ) , .ZN( u1_u14_u5_n191 ) );
  AOI22_X1 u1_u14_u5_U40 (.B2( u1_u14_u5_n131 ) , .A2( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n169 ) , .B1( u1_u14_u5_n174 ) , .A1( u1_u14_u5_n185 ) );
  NOR2_X1 u1_u14_u5_U41 (.A1( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n150 ) , .A2( u1_u14_u5_n173 ) );
  AOI21_X1 u1_u14_u5_U42 (.A( u1_u14_u5_n118 ) , .B2( u1_u14_u5_n145 ) , .ZN( u1_u14_u5_n168 ) , .B1( u1_u14_u5_n186 ) );
  INV_X1 u1_u14_u5_U43 (.A( u1_u14_u5_n122 ) , .ZN( u1_u14_u5_n186 ) );
  NOR2_X1 u1_u14_u5_U44 (.A1( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n152 ) , .A2( u1_u14_u5_n176 ) );
  NOR2_X1 u1_u14_u5_U45 (.A1( u1_u14_u5_n115 ) , .ZN( u1_u14_u5_n118 ) , .A2( u1_u14_u5_n153 ) );
  NOR2_X1 u1_u14_u5_U46 (.A2( u1_u14_u5_n145 ) , .ZN( u1_u14_u5_n156 ) , .A1( u1_u14_u5_n174 ) );
  NOR2_X1 u1_u14_u5_U47 (.ZN( u1_u14_u5_n121 ) , .A2( u1_u14_u5_n145 ) , .A1( u1_u14_u5_n176 ) );
  AOI22_X1 u1_u14_u5_U48 (.ZN( u1_u14_u5_n114 ) , .A2( u1_u14_u5_n137 ) , .A1( u1_u14_u5_n145 ) , .B2( u1_u14_u5_n175 ) , .B1( u1_u14_u5_n193 ) );
  OAI211_X1 u1_u14_u5_U49 (.B( u1_u14_u5_n124 ) , .A( u1_u14_u5_n125 ) , .C2( u1_u14_u5_n126 ) , .C1( u1_u14_u5_n127 ) , .ZN( u1_u14_u5_n128 ) );
  OAI21_X1 u1_u14_u5_U5 (.B2( u1_u14_u5_n136 ) , .B1( u1_u14_u5_n137 ) , .ZN( u1_u14_u5_n138 ) , .A( u1_u14_u5_n177 ) );
  NOR3_X1 u1_u14_u5_U50 (.ZN( u1_u14_u5_n127 ) , .A1( u1_u14_u5_n136 ) , .A3( u1_u14_u5_n148 ) , .A2( u1_u14_u5_n182 ) );
  OAI21_X1 u1_u14_u5_U51 (.ZN( u1_u14_u5_n124 ) , .A( u1_u14_u5_n177 ) , .B2( u1_u14_u5_n183 ) , .B1( u1_u14_u5_n189 ) );
  OAI21_X1 u1_u14_u5_U52 (.ZN( u1_u14_u5_n125 ) , .A( u1_u14_u5_n174 ) , .B2( u1_u14_u5_n185 ) , .B1( u1_u14_u5_n190 ) );
  AOI21_X1 u1_u14_u5_U53 (.A( u1_u14_u5_n153 ) , .B2( u1_u14_u5_n154 ) , .B1( u1_u14_u5_n155 ) , .ZN( u1_u14_u5_n164 ) );
  AOI21_X1 u1_u14_u5_U54 (.ZN( u1_u14_u5_n110 ) , .B1( u1_u14_u5_n122 ) , .B2( u1_u14_u5_n139 ) , .A( u1_u14_u5_n153 ) );
  INV_X1 u1_u14_u5_U55 (.A( u1_u14_u5_n153 ) , .ZN( u1_u14_u5_n176 ) );
  INV_X1 u1_u14_u5_U56 (.A( u1_u14_u5_n126 ) , .ZN( u1_u14_u5_n173 ) );
  AND2_X1 u1_u14_u5_U57 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n147 ) );
  AND2_X1 u1_u14_u5_U58 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n148 ) );
  NAND2_X1 u1_u14_u5_U59 (.A1( u1_u14_u5_n105 ) , .A2( u1_u14_u5_n106 ) , .ZN( u1_u14_u5_n158 ) );
  INV_X1 u1_u14_u5_U6 (.A( u1_u14_u5_n135 ) , .ZN( u1_u14_u5_n178 ) );
  NAND2_X1 u1_u14_u5_U60 (.A2( u1_u14_u5_n108 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n139 ) );
  NAND2_X1 u1_u14_u5_U61 (.A1( u1_u14_u5_n106 ) , .A2( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n119 ) );
  NAND2_X1 u1_u14_u5_U62 (.A2( u1_u14_u5_n103 ) , .A1( u1_u14_u5_n105 ) , .ZN( u1_u14_u5_n140 ) );
  NAND2_X1 u1_u14_u5_U63 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n105 ) , .ZN( u1_u14_u5_n155 ) );
  NAND2_X1 u1_u14_u5_U64 (.A2( u1_u14_u5_n106 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n122 ) );
  NAND2_X1 u1_u14_u5_U65 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n106 ) , .ZN( u1_u14_u5_n115 ) );
  NAND2_X1 u1_u14_u5_U66 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n103 ) , .ZN( u1_u14_u5_n161 ) );
  NAND2_X1 u1_u14_u5_U67 (.A1( u1_u14_u5_n105 ) , .A2( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n154 ) );
  INV_X1 u1_u14_u5_U68 (.A( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n172 ) );
  NAND2_X1 u1_u14_u5_U69 (.A1( u1_u14_u5_n103 ) , .A2( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n123 ) );
  OAI22_X1 u1_u14_u5_U7 (.B2( u1_u14_u5_n149 ) , .B1( u1_u14_u5_n150 ) , .A2( u1_u14_u5_n151 ) , .A1( u1_u14_u5_n152 ) , .ZN( u1_u14_u5_n165 ) );
  NAND2_X1 u1_u14_u5_U70 (.A2( u1_u14_u5_n103 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n151 ) );
  NAND2_X1 u1_u14_u5_U71 (.A2( u1_u14_u5_n107 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n120 ) );
  NAND2_X1 u1_u14_u5_U72 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n157 ) );
  AND2_X1 u1_u14_u5_U73 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n104 ) , .ZN( u1_u14_u5_n131 ) );
  INV_X1 u1_u14_u5_U74 (.A( u1_u14_u5_n102 ) , .ZN( u1_u14_u5_n195 ) );
  OAI221_X1 u1_u14_u5_U75 (.A( u1_u14_u5_n101 ) , .ZN( u1_u14_u5_n102 ) , .C2( u1_u14_u5_n115 ) , .C1( u1_u14_u5_n126 ) , .B1( u1_u14_u5_n134 ) , .B2( u1_u14_u5_n160 ) );
  OAI21_X1 u1_u14_u5_U76 (.ZN( u1_u14_u5_n101 ) , .B1( u1_u14_u5_n137 ) , .A( u1_u14_u5_n146 ) , .B2( u1_u14_u5_n147 ) );
  NOR2_X1 u1_u14_u5_U77 (.A2( u1_u14_X_34 ) , .A1( u1_u14_X_35 ) , .ZN( u1_u14_u5_n145 ) );
  NOR2_X1 u1_u14_u5_U78 (.A2( u1_u14_X_34 ) , .ZN( u1_u14_u5_n146 ) , .A1( u1_u14_u5_n171 ) );
  NOR2_X1 u1_u14_u5_U79 (.A2( u1_u14_X_31 ) , .A1( u1_u14_X_32 ) , .ZN( u1_u14_u5_n103 ) );
  NOR3_X1 u1_u14_u5_U8 (.A2( u1_u14_u5_n147 ) , .A1( u1_u14_u5_n148 ) , .ZN( u1_u14_u5_n149 ) , .A3( u1_u14_u5_n194 ) );
  NOR2_X1 u1_u14_u5_U80 (.A2( u1_u14_X_36 ) , .ZN( u1_u14_u5_n105 ) , .A1( u1_u14_u5_n180 ) );
  NOR2_X1 u1_u14_u5_U81 (.A2( u1_u14_X_33 ) , .ZN( u1_u14_u5_n108 ) , .A1( u1_u14_u5_n170 ) );
  NOR2_X1 u1_u14_u5_U82 (.A2( u1_u14_X_33 ) , .A1( u1_u14_X_36 ) , .ZN( u1_u14_u5_n107 ) );
  NOR2_X1 u1_u14_u5_U83 (.A2( u1_u14_X_31 ) , .ZN( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n181 ) );
  NAND2_X1 u1_u14_u5_U84 (.A2( u1_u14_X_34 ) , .A1( u1_u14_X_35 ) , .ZN( u1_u14_u5_n153 ) );
  NAND2_X1 u1_u14_u5_U85 (.A1( u1_u14_X_34 ) , .ZN( u1_u14_u5_n126 ) , .A2( u1_u14_u5_n171 ) );
  AND2_X1 u1_u14_u5_U86 (.A1( u1_u14_X_31 ) , .A2( u1_u14_X_32 ) , .ZN( u1_u14_u5_n106 ) );
  AND2_X1 u1_u14_u5_U87 (.A1( u1_u14_X_31 ) , .ZN( u1_u14_u5_n109 ) , .A2( u1_u14_u5_n181 ) );
  INV_X1 u1_u14_u5_U88 (.A( u1_u14_X_33 ) , .ZN( u1_u14_u5_n180 ) );
  INV_X1 u1_u14_u5_U89 (.A( u1_u14_X_35 ) , .ZN( u1_u14_u5_n171 ) );
  NOR2_X1 u1_u14_u5_U9 (.ZN( u1_u14_u5_n135 ) , .A1( u1_u14_u5_n173 ) , .A2( u1_u14_u5_n176 ) );
  INV_X1 u1_u14_u5_U90 (.A( u1_u14_X_36 ) , .ZN( u1_u14_u5_n170 ) );
  INV_X1 u1_u14_u5_U91 (.A( u1_u14_X_32 ) , .ZN( u1_u14_u5_n181 ) );
  NAND4_X1 u1_u14_u5_U92 (.ZN( u1_out14_29 ) , .A4( u1_u14_u5_n129 ) , .A3( u1_u14_u5_n130 ) , .A2( u1_u14_u5_n168 ) , .A1( u1_u14_u5_n196 ) );
  AOI221_X1 u1_u14_u5_U93 (.A( u1_u14_u5_n128 ) , .ZN( u1_u14_u5_n129 ) , .C2( u1_u14_u5_n132 ) , .B2( u1_u14_u5_n159 ) , .B1( u1_u14_u5_n176 ) , .C1( u1_u14_u5_n184 ) );
  AOI222_X1 u1_u14_u5_U94 (.ZN( u1_u14_u5_n130 ) , .A2( u1_u14_u5_n146 ) , .B1( u1_u14_u5_n147 ) , .C2( u1_u14_u5_n175 ) , .B2( u1_u14_u5_n179 ) , .A1( u1_u14_u5_n188 ) , .C1( u1_u14_u5_n194 ) );
  NAND4_X1 u1_u14_u5_U95 (.ZN( u1_out14_19 ) , .A4( u1_u14_u5_n166 ) , .A3( u1_u14_u5_n167 ) , .A2( u1_u14_u5_n168 ) , .A1( u1_u14_u5_n169 ) );
  AOI22_X1 u1_u14_u5_U96 (.B2( u1_u14_u5_n145 ) , .A2( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n167 ) , .B1( u1_u14_u5_n182 ) , .A1( u1_u14_u5_n189 ) );
  NOR4_X1 u1_u14_u5_U97 (.A4( u1_u14_u5_n162 ) , .A3( u1_u14_u5_n163 ) , .A2( u1_u14_u5_n164 ) , .A1( u1_u14_u5_n165 ) , .ZN( u1_u14_u5_n166 ) );
  NAND4_X1 u1_u14_u5_U98 (.ZN( u1_out14_11 ) , .A4( u1_u14_u5_n143 ) , .A3( u1_u14_u5_n144 ) , .A2( u1_u14_u5_n169 ) , .A1( u1_u14_u5_n196 ) );
  AOI22_X1 u1_u14_u5_U99 (.A2( u1_u14_u5_n132 ) , .ZN( u1_u14_u5_n144 ) , .B2( u1_u14_u5_n145 ) , .B1( u1_u14_u5_n184 ) , .A1( u1_u14_u5_n194 ) );
  AOI22_X1 u1_u14_u6_U10 (.A2( u1_u14_u6_n151 ) , .B2( u1_u14_u6_n161 ) , .A1( u1_u14_u6_n167 ) , .B1( u1_u14_u6_n170 ) , .ZN( u1_u14_u6_n89 ) );
  AOI21_X1 u1_u14_u6_U11 (.B1( u1_u14_u6_n107 ) , .B2( u1_u14_u6_n132 ) , .A( u1_u14_u6_n158 ) , .ZN( u1_u14_u6_n88 ) );
  AOI21_X1 u1_u14_u6_U12 (.B2( u1_u14_u6_n147 ) , .B1( u1_u14_u6_n148 ) , .ZN( u1_u14_u6_n149 ) , .A( u1_u14_u6_n158 ) );
  AOI21_X1 u1_u14_u6_U13 (.ZN( u1_u14_u6_n106 ) , .A( u1_u14_u6_n142 ) , .B2( u1_u14_u6_n159 ) , .B1( u1_u14_u6_n164 ) );
  INV_X1 u1_u14_u6_U14 (.A( u1_u14_u6_n155 ) , .ZN( u1_u14_u6_n161 ) );
  INV_X1 u1_u14_u6_U15 (.A( u1_u14_u6_n128 ) , .ZN( u1_u14_u6_n164 ) );
  NAND2_X1 u1_u14_u6_U16 (.ZN( u1_u14_u6_n110 ) , .A1( u1_u14_u6_n122 ) , .A2( u1_u14_u6_n129 ) );
  NAND2_X1 u1_u14_u6_U17 (.ZN( u1_u14_u6_n124 ) , .A2( u1_u14_u6_n146 ) , .A1( u1_u14_u6_n148 ) );
  INV_X1 u1_u14_u6_U18 (.A( u1_u14_u6_n132 ) , .ZN( u1_u14_u6_n171 ) );
  AND2_X1 u1_u14_u6_U19 (.A1( u1_u14_u6_n100 ) , .ZN( u1_u14_u6_n130 ) , .A2( u1_u14_u6_n147 ) );
  INV_X1 u1_u14_u6_U20 (.A( u1_u14_u6_n127 ) , .ZN( u1_u14_u6_n173 ) );
  INV_X1 u1_u14_u6_U21 (.A( u1_u14_u6_n121 ) , .ZN( u1_u14_u6_n167 ) );
  INV_X1 u1_u14_u6_U22 (.A( u1_u14_u6_n100 ) , .ZN( u1_u14_u6_n169 ) );
  INV_X1 u1_u14_u6_U23 (.A( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n170 ) );
  INV_X1 u1_u14_u6_U24 (.A( u1_u14_u6_n113 ) , .ZN( u1_u14_u6_n168 ) );
  AND2_X1 u1_u14_u6_U25 (.A1( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n119 ) , .ZN( u1_u14_u6_n133 ) );
  AND2_X1 u1_u14_u6_U26 (.A2( u1_u14_u6_n121 ) , .A1( u1_u14_u6_n122 ) , .ZN( u1_u14_u6_n131 ) );
  AND3_X1 u1_u14_u6_U27 (.ZN( u1_u14_u6_n120 ) , .A2( u1_u14_u6_n127 ) , .A1( u1_u14_u6_n132 ) , .A3( u1_u14_u6_n145 ) );
  INV_X1 u1_u14_u6_U28 (.A( u1_u14_u6_n146 ) , .ZN( u1_u14_u6_n163 ) );
  AOI222_X1 u1_u14_u6_U29 (.ZN( u1_u14_u6_n114 ) , .A1( u1_u14_u6_n118 ) , .A2( u1_u14_u6_n126 ) , .B2( u1_u14_u6_n151 ) , .C2( u1_u14_u6_n159 ) , .C1( u1_u14_u6_n168 ) , .B1( u1_u14_u6_n169 ) );
  INV_X1 u1_u14_u6_U3 (.A( u1_u14_u6_n110 ) , .ZN( u1_u14_u6_n166 ) );
  NOR2_X1 u1_u14_u6_U30 (.A1( u1_u14_u6_n162 ) , .A2( u1_u14_u6_n165 ) , .ZN( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U31 (.A1( u1_u14_u6_n144 ) , .ZN( u1_u14_u6_n151 ) , .A2( u1_u14_u6_n158 ) );
  NAND2_X1 u1_u14_u6_U32 (.ZN( u1_u14_u6_n132 ) , .A1( u1_u14_u6_n91 ) , .A2( u1_u14_u6_n97 ) );
  AOI22_X1 u1_u14_u6_U33 (.B2( u1_u14_u6_n110 ) , .B1( u1_u14_u6_n111 ) , .A1( u1_u14_u6_n112 ) , .ZN( u1_u14_u6_n115 ) , .A2( u1_u14_u6_n161 ) );
  NAND4_X1 u1_u14_u6_U34 (.A3( u1_u14_u6_n109 ) , .ZN( u1_u14_u6_n112 ) , .A4( u1_u14_u6_n132 ) , .A2( u1_u14_u6_n147 ) , .A1( u1_u14_u6_n166 ) );
  NOR2_X1 u1_u14_u6_U35 (.ZN( u1_u14_u6_n109 ) , .A1( u1_u14_u6_n170 ) , .A2( u1_u14_u6_n173 ) );
  NOR2_X1 u1_u14_u6_U36 (.A2( u1_u14_u6_n126 ) , .ZN( u1_u14_u6_n155 ) , .A1( u1_u14_u6_n160 ) );
  NAND2_X1 u1_u14_u6_U37 (.ZN( u1_u14_u6_n146 ) , .A2( u1_u14_u6_n94 ) , .A1( u1_u14_u6_n99 ) );
  AOI21_X1 u1_u14_u6_U38 (.A( u1_u14_u6_n144 ) , .B2( u1_u14_u6_n145 ) , .B1( u1_u14_u6_n146 ) , .ZN( u1_u14_u6_n150 ) );
  AOI211_X1 u1_u14_u6_U39 (.B( u1_u14_u6_n134 ) , .A( u1_u14_u6_n135 ) , .C1( u1_u14_u6_n136 ) , .ZN( u1_u14_u6_n137 ) , .C2( u1_u14_u6_n151 ) );
  INV_X1 u1_u14_u6_U4 (.A( u1_u14_u6_n142 ) , .ZN( u1_u14_u6_n174 ) );
  AOI21_X1 u1_u14_u6_U40 (.B2( u1_u14_u6_n132 ) , .B1( u1_u14_u6_n133 ) , .ZN( u1_u14_u6_n134 ) , .A( u1_u14_u6_n158 ) );
  NAND4_X1 u1_u14_u6_U41 (.A4( u1_u14_u6_n127 ) , .A3( u1_u14_u6_n128 ) , .A2( u1_u14_u6_n129 ) , .A1( u1_u14_u6_n130 ) , .ZN( u1_u14_u6_n136 ) );
  AOI21_X1 u1_u14_u6_U42 (.B1( u1_u14_u6_n131 ) , .ZN( u1_u14_u6_n135 ) , .A( u1_u14_u6_n144 ) , .B2( u1_u14_u6_n146 ) );
  INV_X1 u1_u14_u6_U43 (.A( u1_u14_u6_n111 ) , .ZN( u1_u14_u6_n158 ) );
  NAND2_X1 u1_u14_u6_U44 (.ZN( u1_u14_u6_n127 ) , .A1( u1_u14_u6_n91 ) , .A2( u1_u14_u6_n92 ) );
  NAND2_X1 u1_u14_u6_U45 (.ZN( u1_u14_u6_n129 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n96 ) );
  INV_X1 u1_u14_u6_U46 (.A( u1_u14_u6_n144 ) , .ZN( u1_u14_u6_n159 ) );
  NAND2_X1 u1_u14_u6_U47 (.ZN( u1_u14_u6_n145 ) , .A2( u1_u14_u6_n97 ) , .A1( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U48 (.ZN( u1_u14_u6_n148 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n94 ) );
  NAND2_X1 u1_u14_u6_U49 (.ZN( u1_u14_u6_n108 ) , .A2( u1_u14_u6_n139 ) , .A1( u1_u14_u6_n144 ) );
  NAND2_X1 u1_u14_u6_U5 (.A2( u1_u14_u6_n143 ) , .ZN( u1_u14_u6_n152 ) , .A1( u1_u14_u6_n166 ) );
  NAND2_X1 u1_u14_u6_U50 (.ZN( u1_u14_u6_n121 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n97 ) );
  NAND2_X1 u1_u14_u6_U51 (.ZN( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n95 ) );
  AND2_X1 u1_u14_u6_U52 (.ZN( u1_u14_u6_n118 ) , .A2( u1_u14_u6_n91 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U53 (.ZN( u1_u14_u6_n147 ) , .A2( u1_u14_u6_n98 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U54 (.ZN( u1_u14_u6_n128 ) , .A1( u1_u14_u6_n94 ) , .A2( u1_u14_u6_n96 ) );
  NAND2_X1 u1_u14_u6_U55 (.ZN( u1_u14_u6_n119 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U56 (.ZN( u1_u14_u6_n123 ) , .A2( u1_u14_u6_n91 ) , .A1( u1_u14_u6_n96 ) );
  NAND2_X1 u1_u14_u6_U57 (.ZN( u1_u14_u6_n100 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U58 (.ZN( u1_u14_u6_n122 ) , .A1( u1_u14_u6_n94 ) , .A2( u1_u14_u6_n97 ) );
  INV_X1 u1_u14_u6_U59 (.A( u1_u14_u6_n139 ) , .ZN( u1_u14_u6_n160 ) );
  AOI22_X1 u1_u14_u6_U6 (.B2( u1_u14_u6_n101 ) , .A1( u1_u14_u6_n102 ) , .ZN( u1_u14_u6_n103 ) , .B1( u1_u14_u6_n160 ) , .A2( u1_u14_u6_n161 ) );
  NAND2_X1 u1_u14_u6_U60 (.ZN( u1_u14_u6_n113 ) , .A1( u1_u14_u6_n96 ) , .A2( u1_u14_u6_n98 ) );
  NOR2_X1 u1_u14_u6_U61 (.A2( u1_u14_X_40 ) , .A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n126 ) );
  NOR2_X1 u1_u14_u6_U62 (.A2( u1_u14_X_39 ) , .A1( u1_u14_X_42 ) , .ZN( u1_u14_u6_n92 ) );
  NOR2_X1 u1_u14_u6_U63 (.A2( u1_u14_X_39 ) , .A1( u1_u14_u6_n156 ) , .ZN( u1_u14_u6_n97 ) );
  NOR2_X1 u1_u14_u6_U64 (.A2( u1_u14_X_38 ) , .A1( u1_u14_u6_n165 ) , .ZN( u1_u14_u6_n95 ) );
  NOR2_X1 u1_u14_u6_U65 (.A2( u1_u14_X_41 ) , .ZN( u1_u14_u6_n111 ) , .A1( u1_u14_u6_n157 ) );
  NOR2_X1 u1_u14_u6_U66 (.A2( u1_u14_X_37 ) , .A1( u1_u14_u6_n162 ) , .ZN( u1_u14_u6_n94 ) );
  NOR2_X1 u1_u14_u6_U67 (.A2( u1_u14_X_37 ) , .A1( u1_u14_X_38 ) , .ZN( u1_u14_u6_n91 ) );
  NAND2_X1 u1_u14_u6_U68 (.A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n144 ) , .A2( u1_u14_u6_n157 ) );
  NAND2_X1 u1_u14_u6_U69 (.A2( u1_u14_X_40 ) , .A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n139 ) );
  NOR2_X1 u1_u14_u6_U7 (.A1( u1_u14_u6_n118 ) , .ZN( u1_u14_u6_n143 ) , .A2( u1_u14_u6_n168 ) );
  AND2_X1 u1_u14_u6_U70 (.A1( u1_u14_X_39 ) , .A2( u1_u14_u6_n156 ) , .ZN( u1_u14_u6_n96 ) );
  AND2_X1 u1_u14_u6_U71 (.A1( u1_u14_X_39 ) , .A2( u1_u14_X_42 ) , .ZN( u1_u14_u6_n99 ) );
  INV_X1 u1_u14_u6_U72 (.A( u1_u14_X_40 ) , .ZN( u1_u14_u6_n157 ) );
  INV_X1 u1_u14_u6_U73 (.A( u1_u14_X_37 ) , .ZN( u1_u14_u6_n165 ) );
  INV_X1 u1_u14_u6_U74 (.A( u1_u14_X_38 ) , .ZN( u1_u14_u6_n162 ) );
  INV_X1 u1_u14_u6_U75 (.A( u1_u14_X_42 ) , .ZN( u1_u14_u6_n156 ) );
  NAND4_X1 u1_u14_u6_U76 (.ZN( u1_out14_32 ) , .A4( u1_u14_u6_n103 ) , .A3( u1_u14_u6_n104 ) , .A2( u1_u14_u6_n105 ) , .A1( u1_u14_u6_n106 ) );
  AOI22_X1 u1_u14_u6_U77 (.ZN( u1_u14_u6_n105 ) , .A2( u1_u14_u6_n108 ) , .A1( u1_u14_u6_n118 ) , .B2( u1_u14_u6_n126 ) , .B1( u1_u14_u6_n171 ) );
  AOI22_X1 u1_u14_u6_U78 (.ZN( u1_u14_u6_n104 ) , .A1( u1_u14_u6_n111 ) , .B1( u1_u14_u6_n124 ) , .B2( u1_u14_u6_n151 ) , .A2( u1_u14_u6_n93 ) );
  NAND4_X1 u1_u14_u6_U79 (.ZN( u1_out14_12 ) , .A4( u1_u14_u6_n114 ) , .A3( u1_u14_u6_n115 ) , .A2( u1_u14_u6_n116 ) , .A1( u1_u14_u6_n117 ) );
  INV_X1 u1_u14_u6_U8 (.ZN( u1_u14_u6_n172 ) , .A( u1_u14_u6_n88 ) );
  OAI22_X1 u1_u14_u6_U80 (.B2( u1_u14_u6_n111 ) , .ZN( u1_u14_u6_n116 ) , .B1( u1_u14_u6_n126 ) , .A2( u1_u14_u6_n164 ) , .A1( u1_u14_u6_n167 ) );
  OAI21_X1 u1_u14_u6_U81 (.A( u1_u14_u6_n108 ) , .ZN( u1_u14_u6_n117 ) , .B2( u1_u14_u6_n141 ) , .B1( u1_u14_u6_n163 ) );
  OAI211_X1 u1_u14_u6_U82 (.ZN( u1_out14_22 ) , .B( u1_u14_u6_n137 ) , .A( u1_u14_u6_n138 ) , .C2( u1_u14_u6_n139 ) , .C1( u1_u14_u6_n140 ) );
  AOI22_X1 u1_u14_u6_U83 (.B1( u1_u14_u6_n124 ) , .A2( u1_u14_u6_n125 ) , .A1( u1_u14_u6_n126 ) , .ZN( u1_u14_u6_n138 ) , .B2( u1_u14_u6_n161 ) );
  AND4_X1 u1_u14_u6_U84 (.A3( u1_u14_u6_n119 ) , .A1( u1_u14_u6_n120 ) , .A4( u1_u14_u6_n129 ) , .ZN( u1_u14_u6_n140 ) , .A2( u1_u14_u6_n143 ) );
  OAI211_X1 u1_u14_u6_U85 (.ZN( u1_out14_7 ) , .B( u1_u14_u6_n153 ) , .C2( u1_u14_u6_n154 ) , .C1( u1_u14_u6_n155 ) , .A( u1_u14_u6_n174 ) );
  NOR3_X1 u1_u14_u6_U86 (.A1( u1_u14_u6_n141 ) , .ZN( u1_u14_u6_n154 ) , .A3( u1_u14_u6_n164 ) , .A2( u1_u14_u6_n171 ) );
  AOI211_X1 u1_u14_u6_U87 (.B( u1_u14_u6_n149 ) , .A( u1_u14_u6_n150 ) , .C2( u1_u14_u6_n151 ) , .C1( u1_u14_u6_n152 ) , .ZN( u1_u14_u6_n153 ) );
  NAND3_X1 u1_u14_u6_U88 (.A2( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n125 ) , .A1( u1_u14_u6_n130 ) , .A3( u1_u14_u6_n131 ) );
  NAND3_X1 u1_u14_u6_U89 (.A3( u1_u14_u6_n133 ) , .ZN( u1_u14_u6_n141 ) , .A1( u1_u14_u6_n145 ) , .A2( u1_u14_u6_n148 ) );
  OAI21_X1 u1_u14_u6_U9 (.A( u1_u14_u6_n159 ) , .B1( u1_u14_u6_n169 ) , .B2( u1_u14_u6_n173 ) , .ZN( u1_u14_u6_n90 ) );
  NAND3_X1 u1_u14_u6_U90 (.ZN( u1_u14_u6_n101 ) , .A3( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n121 ) , .A1( u1_u14_u6_n127 ) );
  NAND3_X1 u1_u14_u6_U91 (.ZN( u1_u14_u6_n102 ) , .A3( u1_u14_u6_n130 ) , .A2( u1_u14_u6_n145 ) , .A1( u1_u14_u6_n166 ) );
  NAND3_X1 u1_u14_u6_U92 (.A3( u1_u14_u6_n113 ) , .A1( u1_u14_u6_n119 ) , .A2( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n93 ) );
  NAND3_X1 u1_u14_u6_U93 (.ZN( u1_u14_u6_n142 ) , .A2( u1_u14_u6_n172 ) , .A3( u1_u14_u6_n89 ) , .A1( u1_u14_u6_n90 ) );
  OAI21_X1 u1_u14_u7_U10 (.A( u1_u14_u7_n161 ) , .B1( u1_u14_u7_n168 ) , .B2( u1_u14_u7_n173 ) , .ZN( u1_u14_u7_n91 ) );
  AOI211_X1 u1_u14_u7_U11 (.A( u1_u14_u7_n117 ) , .ZN( u1_u14_u7_n118 ) , .C2( u1_u14_u7_n126 ) , .C1( u1_u14_u7_n177 ) , .B( u1_u14_u7_n180 ) );
  OAI22_X1 u1_u14_u7_U12 (.B1( u1_u14_u7_n115 ) , .ZN( u1_u14_u7_n117 ) , .A2( u1_u14_u7_n133 ) , .A1( u1_u14_u7_n137 ) , .B2( u1_u14_u7_n162 ) );
  INV_X1 u1_u14_u7_U13 (.A( u1_u14_u7_n116 ) , .ZN( u1_u14_u7_n180 ) );
  NOR3_X1 u1_u14_u7_U14 (.ZN( u1_u14_u7_n115 ) , .A3( u1_u14_u7_n145 ) , .A2( u1_u14_u7_n168 ) , .A1( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U15 (.A( u1_u14_u7_n133 ) , .ZN( u1_u14_u7_n176 ) );
  NOR3_X1 u1_u14_u7_U16 (.A2( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n135 ) , .ZN( u1_u14_u7_n136 ) , .A3( u1_u14_u7_n171 ) );
  NOR2_X1 u1_u14_u7_U17 (.A1( u1_u14_u7_n130 ) , .A2( u1_u14_u7_n134 ) , .ZN( u1_u14_u7_n153 ) );
  AOI21_X1 u1_u14_u7_U18 (.ZN( u1_u14_u7_n104 ) , .B2( u1_u14_u7_n112 ) , .B1( u1_u14_u7_n127 ) , .A( u1_u14_u7_n164 ) );
  AOI21_X1 u1_u14_u7_U19 (.ZN( u1_u14_u7_n106 ) , .B1( u1_u14_u7_n133 ) , .B2( u1_u14_u7_n146 ) , .A( u1_u14_u7_n162 ) );
  AOI21_X1 u1_u14_u7_U20 (.A( u1_u14_u7_n101 ) , .ZN( u1_u14_u7_n107 ) , .B2( u1_u14_u7_n128 ) , .B1( u1_u14_u7_n175 ) );
  INV_X1 u1_u14_u7_U21 (.A( u1_u14_u7_n101 ) , .ZN( u1_u14_u7_n165 ) );
  NOR2_X1 u1_u14_u7_U22 (.ZN( u1_u14_u7_n111 ) , .A2( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U23 (.A( u1_u14_u7_n138 ) , .ZN( u1_u14_u7_n171 ) );
  INV_X1 u1_u14_u7_U24 (.A( u1_u14_u7_n131 ) , .ZN( u1_u14_u7_n177 ) );
  INV_X1 u1_u14_u7_U25 (.A( u1_u14_u7_n110 ) , .ZN( u1_u14_u7_n174 ) );
  NAND2_X1 u1_u14_u7_U26 (.A1( u1_u14_u7_n129 ) , .A2( u1_u14_u7_n132 ) , .ZN( u1_u14_u7_n149 ) );
  NAND2_X1 u1_u14_u7_U27 (.A1( u1_u14_u7_n113 ) , .A2( u1_u14_u7_n124 ) , .ZN( u1_u14_u7_n130 ) );
  INV_X1 u1_u14_u7_U28 (.A( u1_u14_u7_n112 ) , .ZN( u1_u14_u7_n173 ) );
  INV_X1 u1_u14_u7_U29 (.A( u1_u14_u7_n128 ) , .ZN( u1_u14_u7_n168 ) );
  OAI21_X1 u1_u14_u7_U3 (.ZN( u1_u14_u7_n159 ) , .A( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n171 ) , .B1( u1_u14_u7_n174 ) );
  INV_X1 u1_u14_u7_U30 (.A( u1_u14_u7_n148 ) , .ZN( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U31 (.A( u1_u14_u7_n127 ) , .ZN( u1_u14_u7_n179 ) );
  NOR2_X1 u1_u14_u7_U32 (.ZN( u1_u14_u7_n101 ) , .A2( u1_u14_u7_n150 ) , .A1( u1_u14_u7_n156 ) );
  AOI211_X1 u1_u14_u7_U33 (.B( u1_u14_u7_n139 ) , .A( u1_u14_u7_n140 ) , .C2( u1_u14_u7_n141 ) , .ZN( u1_u14_u7_n142 ) , .C1( u1_u14_u7_n156 ) );
  NAND4_X1 u1_u14_u7_U34 (.A3( u1_u14_u7_n127 ) , .A2( u1_u14_u7_n128 ) , .A1( u1_u14_u7_n129 ) , .ZN( u1_u14_u7_n141 ) , .A4( u1_u14_u7_n147 ) );
  AOI21_X1 u1_u14_u7_U35 (.A( u1_u14_u7_n137 ) , .B1( u1_u14_u7_n138 ) , .ZN( u1_u14_u7_n139 ) , .B2( u1_u14_u7_n146 ) );
  OAI22_X1 u1_u14_u7_U36 (.B1( u1_u14_u7_n136 ) , .ZN( u1_u14_u7_n140 ) , .A1( u1_u14_u7_n153 ) , .B2( u1_u14_u7_n162 ) , .A2( u1_u14_u7_n164 ) );
  INV_X1 u1_u14_u7_U37 (.A( u1_u14_u7_n125 ) , .ZN( u1_u14_u7_n161 ) );
  AOI21_X1 u1_u14_u7_U38 (.ZN( u1_u14_u7_n123 ) , .B1( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n177 ) , .A( u1_u14_u7_n97 ) );
  AOI21_X1 u1_u14_u7_U39 (.B2( u1_u14_u7_n113 ) , .B1( u1_u14_u7_n124 ) , .A( u1_u14_u7_n125 ) , .ZN( u1_u14_u7_n97 ) );
  INV_X1 u1_u14_u7_U4 (.A( u1_u14_u7_n149 ) , .ZN( u1_u14_u7_n175 ) );
  INV_X1 u1_u14_u7_U40 (.A( u1_u14_u7_n152 ) , .ZN( u1_u14_u7_n162 ) );
  AOI22_X1 u1_u14_u7_U41 (.A2( u1_u14_u7_n114 ) , .ZN( u1_u14_u7_n119 ) , .B1( u1_u14_u7_n130 ) , .A1( u1_u14_u7_n156 ) , .B2( u1_u14_u7_n165 ) );
  NAND2_X1 u1_u14_u7_U42 (.A2( u1_u14_u7_n112 ) , .ZN( u1_u14_u7_n114 ) , .A1( u1_u14_u7_n175 ) );
  NOR2_X1 u1_u14_u7_U43 (.ZN( u1_u14_u7_n137 ) , .A1( u1_u14_u7_n150 ) , .A2( u1_u14_u7_n161 ) );
  AND2_X1 u1_u14_u7_U44 (.ZN( u1_u14_u7_n145 ) , .A2( u1_u14_u7_n98 ) , .A1( u1_u14_u7_n99 ) );
  AOI21_X1 u1_u14_u7_U45 (.ZN( u1_u14_u7_n105 ) , .B2( u1_u14_u7_n110 ) , .A( u1_u14_u7_n125 ) , .B1( u1_u14_u7_n147 ) );
  NAND2_X1 u1_u14_u7_U46 (.ZN( u1_u14_u7_n146 ) , .A1( u1_u14_u7_n95 ) , .A2( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U47 (.A2( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n147 ) , .A1( u1_u14_u7_n93 ) );
  NAND2_X1 u1_u14_u7_U48 (.A1( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n127 ) , .A2( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U49 (.A2( u1_u14_u7_n102 ) , .A1( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n133 ) );
  INV_X1 u1_u14_u7_U5 (.A( u1_u14_u7_n154 ) , .ZN( u1_u14_u7_n178 ) );
  OR2_X1 u1_u14_u7_U50 (.ZN( u1_u14_u7_n126 ) , .A2( u1_u14_u7_n152 ) , .A1( u1_u14_u7_n156 ) );
  NAND2_X1 u1_u14_u7_U51 (.ZN( u1_u14_u7_n112 ) , .A2( u1_u14_u7_n96 ) , .A1( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U52 (.A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n128 ) , .A1( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U53 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n113 ) , .A2( u1_u14_u7_n93 ) );
  NAND2_X1 u1_u14_u7_U54 (.ZN( u1_u14_u7_n110 ) , .A1( u1_u14_u7_n95 ) , .A2( u1_u14_u7_n96 ) );
  INV_X1 u1_u14_u7_U55 (.A( u1_u14_u7_n150 ) , .ZN( u1_u14_u7_n164 ) );
  AND2_X1 u1_u14_u7_U56 (.ZN( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n93 ) , .A2( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U57 (.A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n124 ) , .A1( u1_u14_u7_n96 ) );
  NAND2_X1 u1_u14_u7_U58 (.A1( u1_u14_u7_n100 ) , .A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n129 ) );
  NAND2_X1 u1_u14_u7_U59 (.A2( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n131 ) , .A1( u1_u14_u7_n95 ) );
  AOI211_X1 u1_u14_u7_U6 (.ZN( u1_u14_u7_n116 ) , .A( u1_u14_u7_n155 ) , .C1( u1_u14_u7_n161 ) , .C2( u1_u14_u7_n171 ) , .B( u1_u14_u7_n94 ) );
  NAND2_X1 u1_u14_u7_U60 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n138 ) , .A2( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U61 (.ZN( u1_u14_u7_n132 ) , .A1( u1_u14_u7_n93 ) , .A2( u1_u14_u7_n96 ) );
  NAND2_X1 u1_u14_u7_U62 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n148 ) , .A2( u1_u14_u7_n95 ) );
  AOI211_X1 u1_u14_u7_U63 (.B( u1_u14_u7_n154 ) , .A( u1_u14_u7_n155 ) , .C1( u1_u14_u7_n156 ) , .ZN( u1_u14_u7_n157 ) , .C2( u1_u14_u7_n172 ) );
  INV_X1 u1_u14_u7_U64 (.A( u1_u14_u7_n153 ) , .ZN( u1_u14_u7_n172 ) );
  NOR2_X1 u1_u14_u7_U65 (.A2( u1_u14_X_47 ) , .ZN( u1_u14_u7_n150 ) , .A1( u1_u14_u7_n163 ) );
  NOR2_X1 u1_u14_u7_U66 (.A2( u1_u14_X_43 ) , .A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n103 ) );
  NOR2_X1 u1_u14_u7_U67 (.A2( u1_u14_X_48 ) , .A1( u1_u14_u7_n166 ) , .ZN( u1_u14_u7_n95 ) );
  NOR2_X1 u1_u14_u7_U68 (.A2( u1_u14_X_45 ) , .A1( u1_u14_X_48 ) , .ZN( u1_u14_u7_n99 ) );
  NOR2_X1 u1_u14_u7_U69 (.A2( u1_u14_X_44 ) , .A1( u1_u14_u7_n167 ) , .ZN( u1_u14_u7_n98 ) );
  OAI222_X1 u1_u14_u7_U7 (.C2( u1_u14_u7_n101 ) , .B2( u1_u14_u7_n111 ) , .A1( u1_u14_u7_n113 ) , .C1( u1_u14_u7_n146 ) , .A2( u1_u14_u7_n162 ) , .B1( u1_u14_u7_n164 ) , .ZN( u1_u14_u7_n94 ) );
  NOR2_X1 u1_u14_u7_U70 (.A2( u1_u14_X_46 ) , .A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n152 ) );
  NAND2_X1 u1_u14_u7_U71 (.A2( u1_u14_X_46 ) , .A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n125 ) );
  AND2_X1 u1_u14_u7_U72 (.A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n156 ) , .A2( u1_u14_u7_n163 ) );
  AND2_X1 u1_u14_u7_U73 (.A2( u1_u14_X_45 ) , .A1( u1_u14_X_48 ) , .ZN( u1_u14_u7_n102 ) );
  AND2_X1 u1_u14_u7_U74 (.A2( u1_u14_X_43 ) , .A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n96 ) );
  AND2_X1 u1_u14_u7_U75 (.A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n100 ) , .A2( u1_u14_u7_n167 ) );
  AND2_X1 u1_u14_u7_U76 (.A1( u1_u14_X_48 ) , .A2( u1_u14_u7_n166 ) , .ZN( u1_u14_u7_n93 ) );
  INV_X1 u1_u14_u7_U77 (.A( u1_u14_X_46 ) , .ZN( u1_u14_u7_n163 ) );
  INV_X1 u1_u14_u7_U78 (.A( u1_u14_X_43 ) , .ZN( u1_u14_u7_n167 ) );
  INV_X1 u1_u14_u7_U79 (.A( u1_u14_X_45 ) , .ZN( u1_u14_u7_n166 ) );
  OAI221_X1 u1_u14_u7_U8 (.C1( u1_u14_u7_n101 ) , .C2( u1_u14_u7_n147 ) , .ZN( u1_u14_u7_n155 ) , .B2( u1_u14_u7_n162 ) , .A( u1_u14_u7_n91 ) , .B1( u1_u14_u7_n92 ) );
  NAND4_X1 u1_u14_u7_U80 (.ZN( u1_out14_5 ) , .A4( u1_u14_u7_n108 ) , .A3( u1_u14_u7_n109 ) , .A1( u1_u14_u7_n116 ) , .A2( u1_u14_u7_n123 ) );
  AOI22_X1 u1_u14_u7_U81 (.ZN( u1_u14_u7_n109 ) , .A2( u1_u14_u7_n126 ) , .B2( u1_u14_u7_n145 ) , .B1( u1_u14_u7_n156 ) , .A1( u1_u14_u7_n171 ) );
  NOR4_X1 u1_u14_u7_U82 (.A4( u1_u14_u7_n104 ) , .A3( u1_u14_u7_n105 ) , .A2( u1_u14_u7_n106 ) , .A1( u1_u14_u7_n107 ) , .ZN( u1_u14_u7_n108 ) );
  NAND4_X1 u1_u14_u7_U83 (.ZN( u1_out14_27 ) , .A4( u1_u14_u7_n118 ) , .A3( u1_u14_u7_n119 ) , .A2( u1_u14_u7_n120 ) , .A1( u1_u14_u7_n121 ) );
  OAI21_X1 u1_u14_u7_U84 (.ZN( u1_u14_u7_n121 ) , .B2( u1_u14_u7_n145 ) , .A( u1_u14_u7_n150 ) , .B1( u1_u14_u7_n174 ) );
  OAI21_X1 u1_u14_u7_U85 (.ZN( u1_u14_u7_n120 ) , .A( u1_u14_u7_n161 ) , .B2( u1_u14_u7_n170 ) , .B1( u1_u14_u7_n179 ) );
  NAND4_X1 u1_u14_u7_U86 (.ZN( u1_out14_21 ) , .A4( u1_u14_u7_n157 ) , .A3( u1_u14_u7_n158 ) , .A2( u1_u14_u7_n159 ) , .A1( u1_u14_u7_n160 ) );
  OAI21_X1 u1_u14_u7_U87 (.B1( u1_u14_u7_n145 ) , .ZN( u1_u14_u7_n160 ) , .A( u1_u14_u7_n161 ) , .B2( u1_u14_u7_n177 ) );
  AOI22_X1 u1_u14_u7_U88 (.B2( u1_u14_u7_n149 ) , .B1( u1_u14_u7_n150 ) , .A2( u1_u14_u7_n151 ) , .A1( u1_u14_u7_n152 ) , .ZN( u1_u14_u7_n158 ) );
  NAND4_X1 u1_u14_u7_U89 (.ZN( u1_out14_15 ) , .A4( u1_u14_u7_n142 ) , .A3( u1_u14_u7_n143 ) , .A2( u1_u14_u7_n144 ) , .A1( u1_u14_u7_n178 ) );
  AND3_X1 u1_u14_u7_U9 (.A3( u1_u14_u7_n110 ) , .A2( u1_u14_u7_n127 ) , .A1( u1_u14_u7_n132 ) , .ZN( u1_u14_u7_n92 ) );
  OR2_X1 u1_u14_u7_U90 (.A2( u1_u14_u7_n125 ) , .A1( u1_u14_u7_n129 ) , .ZN( u1_u14_u7_n144 ) );
  AOI22_X1 u1_u14_u7_U91 (.A2( u1_u14_u7_n126 ) , .ZN( u1_u14_u7_n143 ) , .B2( u1_u14_u7_n165 ) , .B1( u1_u14_u7_n173 ) , .A1( u1_u14_u7_n174 ) );
  OAI211_X1 u1_u14_u7_U92 (.B( u1_u14_u7_n122 ) , .A( u1_u14_u7_n123 ) , .C2( u1_u14_u7_n124 ) , .ZN( u1_u14_u7_n154 ) , .C1( u1_u14_u7_n162 ) );
  AOI222_X1 u1_u14_u7_U93 (.ZN( u1_u14_u7_n122 ) , .C2( u1_u14_u7_n126 ) , .C1( u1_u14_u7_n145 ) , .B1( u1_u14_u7_n161 ) , .A2( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n170 ) , .A1( u1_u14_u7_n176 ) );
  INV_X1 u1_u14_u7_U94 (.A( u1_u14_u7_n111 ) , .ZN( u1_u14_u7_n170 ) );
  NAND3_X1 u1_u14_u7_U95 (.A3( u1_u14_u7_n146 ) , .A2( u1_u14_u7_n147 ) , .A1( u1_u14_u7_n148 ) , .ZN( u1_u14_u7_n151 ) );
  NAND3_X1 u1_u14_u7_U96 (.A3( u1_u14_u7_n131 ) , .A2( u1_u14_u7_n132 ) , .A1( u1_u14_u7_n133 ) , .ZN( u1_u14_u7_n135 ) );
  XOR2_X1 u1_u15_U21 (.A( u1_FP_56 ) , .B( u1_K16_35 ) , .Z( u1_u15_X_35 ) );
  XOR2_X1 u1_u15_U22 (.A( u1_FP_55 ) , .B( u1_K16_34 ) , .Z( u1_u15_X_34 ) );
  XOR2_X1 u1_u15_U24 (.A( u1_FP_53 ) , .B( u1_K16_32 ) , .Z( u1_u15_X_32 ) );
  XOR2_X1 u1_u15_U25 (.A( u1_FP_52 ) , .B( u1_K16_31 ) , .Z( u1_u15_X_31 ) );
  XOR2_X1 u1_u15_U26 (.A( u1_FP_53 ) , .B( u1_K16_30 ) , .Z( u1_u15_X_30 ) );
  XOR2_X1 u1_u15_U28 (.A( u1_FP_52 ) , .B( u1_K16_29 ) , .Z( u1_u15_X_29 ) );
  XOR2_X1 u1_u15_U37 (.A( u1_FP_45 ) , .B( u1_K16_20 ) , .Z( u1_u15_X_20 ) );
  XOR2_X1 u1_u15_U39 (.A( u1_FP_44 ) , .B( u1_K16_19 ) , .Z( u1_u15_X_19 ) );
  XOR2_X1 u1_u15_U40 (.A( u1_FP_45 ) , .B( u1_K16_18 ) , .Z( u1_u15_X_18 ) );
  XOR2_X1 u1_u15_U41 (.A( u1_FP_44 ) , .B( u1_K16_17 ) , .Z( u1_u15_X_17 ) );
  XOR2_X1 u1_u15_U44 (.A( u1_FP_41 ) , .B( u1_K16_14 ) , .Z( u1_u15_X_14 ) );
  XOR2_X1 u1_u15_U45 (.A( u1_FP_40 ) , .B( u1_K16_13 ) , .Z( u1_u15_X_13 ) );
  OAI22_X1 u1_u15_u2_U10 (.B1( u1_u15_u2_n151 ) , .A2( u1_u15_u2_n152 ) , .A1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n160 ) , .B2( u1_u15_u2_n168 ) );
  NAND3_X1 u1_u15_u2_U100 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n98 ) );
  NOR3_X1 u1_u15_u2_U11 (.A1( u1_u15_u2_n150 ) , .ZN( u1_u15_u2_n151 ) , .A3( u1_u15_u2_n175 ) , .A2( u1_u15_u2_n188 ) );
  AOI21_X1 u1_u15_u2_U12 (.B2( u1_u15_u2_n123 ) , .ZN( u1_u15_u2_n125 ) , .A( u1_u15_u2_n171 ) , .B1( u1_u15_u2_n184 ) );
  INV_X1 u1_u15_u2_U13 (.A( u1_u15_u2_n150 ) , .ZN( u1_u15_u2_n184 ) );
  AOI21_X1 u1_u15_u2_U14 (.ZN( u1_u15_u2_n144 ) , .B2( u1_u15_u2_n155 ) , .A( u1_u15_u2_n172 ) , .B1( u1_u15_u2_n185 ) );
  AOI21_X1 u1_u15_u2_U15 (.B2( u1_u15_u2_n143 ) , .ZN( u1_u15_u2_n145 ) , .B1( u1_u15_u2_n152 ) , .A( u1_u15_u2_n171 ) );
  INV_X1 u1_u15_u2_U16 (.A( u1_u15_u2_n156 ) , .ZN( u1_u15_u2_n171 ) );
  INV_X1 u1_u15_u2_U17 (.A( u1_u15_u2_n120 ) , .ZN( u1_u15_u2_n188 ) );
  NAND2_X1 u1_u15_u2_U18 (.A2( u1_u15_u2_n122 ) , .ZN( u1_u15_u2_n150 ) , .A1( u1_u15_u2_n152 ) );
  INV_X1 u1_u15_u2_U19 (.A( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n170 ) );
  INV_X1 u1_u15_u2_U20 (.A( u1_u15_u2_n137 ) , .ZN( u1_u15_u2_n173 ) );
  NAND2_X1 u1_u15_u2_U21 (.A1( u1_u15_u2_n132 ) , .A2( u1_u15_u2_n139 ) , .ZN( u1_u15_u2_n157 ) );
  INV_X1 u1_u15_u2_U22 (.A( u1_u15_u2_n113 ) , .ZN( u1_u15_u2_n178 ) );
  INV_X1 u1_u15_u2_U23 (.A( u1_u15_u2_n139 ) , .ZN( u1_u15_u2_n175 ) );
  INV_X1 u1_u15_u2_U24 (.A( u1_u15_u2_n155 ) , .ZN( u1_u15_u2_n181 ) );
  INV_X1 u1_u15_u2_U25 (.A( u1_u15_u2_n119 ) , .ZN( u1_u15_u2_n177 ) );
  INV_X1 u1_u15_u2_U26 (.A( u1_u15_u2_n116 ) , .ZN( u1_u15_u2_n180 ) );
  INV_X1 u1_u15_u2_U27 (.A( u1_u15_u2_n131 ) , .ZN( u1_u15_u2_n179 ) );
  INV_X1 u1_u15_u2_U28 (.A( u1_u15_u2_n154 ) , .ZN( u1_u15_u2_n176 ) );
  NAND2_X1 u1_u15_u2_U29 (.A2( u1_u15_u2_n116 ) , .A1( u1_u15_u2_n117 ) , .ZN( u1_u15_u2_n118 ) );
  NOR2_X1 u1_u15_u2_U3 (.ZN( u1_u15_u2_n121 ) , .A2( u1_u15_u2_n177 ) , .A1( u1_u15_u2_n180 ) );
  INV_X1 u1_u15_u2_U30 (.A( u1_u15_u2_n132 ) , .ZN( u1_u15_u2_n182 ) );
  INV_X1 u1_u15_u2_U31 (.A( u1_u15_u2_n158 ) , .ZN( u1_u15_u2_n183 ) );
  OAI21_X1 u1_u15_u2_U32 (.A( u1_u15_u2_n156 ) , .B1( u1_u15_u2_n157 ) , .ZN( u1_u15_u2_n158 ) , .B2( u1_u15_u2_n179 ) );
  NOR2_X1 u1_u15_u2_U33 (.ZN( u1_u15_u2_n156 ) , .A1( u1_u15_u2_n166 ) , .A2( u1_u15_u2_n169 ) );
  NOR2_X1 u1_u15_u2_U34 (.A2( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n137 ) , .A1( u1_u15_u2_n140 ) );
  NOR2_X1 u1_u15_u2_U35 (.A2( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n153 ) , .A1( u1_u15_u2_n156 ) );
  AOI211_X1 u1_u15_u2_U36 (.ZN( u1_u15_u2_n130 ) , .C1( u1_u15_u2_n138 ) , .C2( u1_u15_u2_n179 ) , .B( u1_u15_u2_n96 ) , .A( u1_u15_u2_n97 ) );
  OAI22_X1 u1_u15_u2_U37 (.B1( u1_u15_u2_n133 ) , .A2( u1_u15_u2_n137 ) , .A1( u1_u15_u2_n152 ) , .B2( u1_u15_u2_n168 ) , .ZN( u1_u15_u2_n97 ) );
  OAI221_X1 u1_u15_u2_U38 (.B1( u1_u15_u2_n113 ) , .C1( u1_u15_u2_n132 ) , .A( u1_u15_u2_n149 ) , .B2( u1_u15_u2_n171 ) , .C2( u1_u15_u2_n172 ) , .ZN( u1_u15_u2_n96 ) );
  OAI221_X1 u1_u15_u2_U39 (.A( u1_u15_u2_n115 ) , .C2( u1_u15_u2_n123 ) , .B2( u1_u15_u2_n143 ) , .B1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n163 ) , .C1( u1_u15_u2_n168 ) );
  INV_X1 u1_u15_u2_U4 (.A( u1_u15_u2_n134 ) , .ZN( u1_u15_u2_n185 ) );
  OAI21_X1 u1_u15_u2_U40 (.A( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n115 ) , .B1( u1_u15_u2_n176 ) , .B2( u1_u15_u2_n178 ) );
  OAI221_X1 u1_u15_u2_U41 (.A( u1_u15_u2_n135 ) , .B2( u1_u15_u2_n136 ) , .B1( u1_u15_u2_n137 ) , .ZN( u1_u15_u2_n162 ) , .C2( u1_u15_u2_n167 ) , .C1( u1_u15_u2_n185 ) );
  AND3_X1 u1_u15_u2_U42 (.A3( u1_u15_u2_n131 ) , .A2( u1_u15_u2_n132 ) , .A1( u1_u15_u2_n133 ) , .ZN( u1_u15_u2_n136 ) );
  AOI22_X1 u1_u15_u2_U43 (.ZN( u1_u15_u2_n135 ) , .B1( u1_u15_u2_n140 ) , .A1( u1_u15_u2_n156 ) , .B2( u1_u15_u2_n180 ) , .A2( u1_u15_u2_n188 ) );
  AOI21_X1 u1_u15_u2_U44 (.ZN( u1_u15_u2_n149 ) , .B1( u1_u15_u2_n173 ) , .B2( u1_u15_u2_n188 ) , .A( u1_u15_u2_n95 ) );
  AND3_X1 u1_u15_u2_U45 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n156 ) , .ZN( u1_u15_u2_n95 ) );
  OAI21_X1 u1_u15_u2_U46 (.A( u1_u15_u2_n101 ) , .B2( u1_u15_u2_n121 ) , .B1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n164 ) );
  NAND2_X1 u1_u15_u2_U47 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n155 ) );
  NAND2_X1 u1_u15_u2_U48 (.A2( u1_u15_u2_n105 ) , .A1( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n143 ) );
  NAND2_X1 u1_u15_u2_U49 (.A1( u1_u15_u2_n104 ) , .A2( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n152 ) );
  NOR4_X1 u1_u15_u2_U5 (.A4( u1_u15_u2_n124 ) , .A3( u1_u15_u2_n125 ) , .A2( u1_u15_u2_n126 ) , .A1( u1_u15_u2_n127 ) , .ZN( u1_u15_u2_n128 ) );
  NAND2_X1 u1_u15_u2_U50 (.A1( u1_u15_u2_n100 ) , .A2( u1_u15_u2_n105 ) , .ZN( u1_u15_u2_n132 ) );
  INV_X1 u1_u15_u2_U51 (.A( u1_u15_u2_n140 ) , .ZN( u1_u15_u2_n168 ) );
  INV_X1 u1_u15_u2_U52 (.A( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n167 ) );
  OAI21_X1 u1_u15_u2_U53 (.A( u1_u15_u2_n141 ) , .B2( u1_u15_u2_n142 ) , .ZN( u1_u15_u2_n146 ) , .B1( u1_u15_u2_n153 ) );
  OAI21_X1 u1_u15_u2_U54 (.A( u1_u15_u2_n140 ) , .ZN( u1_u15_u2_n141 ) , .B1( u1_u15_u2_n176 ) , .B2( u1_u15_u2_n177 ) );
  NOR3_X1 u1_u15_u2_U55 (.ZN( u1_u15_u2_n142 ) , .A3( u1_u15_u2_n175 ) , .A2( u1_u15_u2_n178 ) , .A1( u1_u15_u2_n181 ) );
  INV_X1 u1_u15_u2_U56 (.ZN( u1_u15_u2_n187 ) , .A( u1_u15_u2_n99 ) );
  OAI21_X1 u1_u15_u2_U57 (.B1( u1_u15_u2_n137 ) , .B2( u1_u15_u2_n143 ) , .A( u1_u15_u2_n98 ) , .ZN( u1_u15_u2_n99 ) );
  NAND2_X1 u1_u15_u2_U58 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n113 ) );
  NAND2_X1 u1_u15_u2_U59 (.A1( u1_u15_u2_n106 ) , .A2( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n131 ) );
  AOI21_X1 u1_u15_u2_U6 (.B2( u1_u15_u2_n119 ) , .ZN( u1_u15_u2_n127 ) , .A( u1_u15_u2_n137 ) , .B1( u1_u15_u2_n155 ) );
  NAND2_X1 u1_u15_u2_U60 (.A1( u1_u15_u2_n103 ) , .A2( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n139 ) );
  NAND2_X1 u1_u15_u2_U61 (.A1( u1_u15_u2_n103 ) , .A2( u1_u15_u2_n105 ) , .ZN( u1_u15_u2_n133 ) );
  NAND2_X1 u1_u15_u2_U62 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n103 ) , .ZN( u1_u15_u2_n154 ) );
  NAND2_X1 u1_u15_u2_U63 (.A2( u1_u15_u2_n103 ) , .A1( u1_u15_u2_n104 ) , .ZN( u1_u15_u2_n119 ) );
  NAND2_X1 u1_u15_u2_U64 (.A2( u1_u15_u2_n107 ) , .A1( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n123 ) );
  NAND2_X1 u1_u15_u2_U65 (.A1( u1_u15_u2_n104 ) , .A2( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n122 ) );
  INV_X1 u1_u15_u2_U66 (.A( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n172 ) );
  NAND2_X1 u1_u15_u2_U67 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n102 ) , .ZN( u1_u15_u2_n116 ) );
  NAND2_X1 u1_u15_u2_U68 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n120 ) );
  NAND2_X1 u1_u15_u2_U69 (.A2( u1_u15_u2_n105 ) , .A1( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n117 ) );
  AOI21_X1 u1_u15_u2_U7 (.ZN( u1_u15_u2_n124 ) , .B1( u1_u15_u2_n131 ) , .B2( u1_u15_u2_n143 ) , .A( u1_u15_u2_n172 ) );
  NOR2_X1 u1_u15_u2_U70 (.A2( u1_u15_X_16 ) , .ZN( u1_u15_u2_n140 ) , .A1( u1_u15_u2_n166 ) );
  NOR2_X1 u1_u15_u2_U71 (.A2( u1_u15_X_13 ) , .A1( u1_u15_X_14 ) , .ZN( u1_u15_u2_n100 ) );
  NOR2_X1 u1_u15_u2_U72 (.A2( u1_u15_X_16 ) , .A1( u1_u15_X_17 ) , .ZN( u1_u15_u2_n138 ) );
  NOR2_X1 u1_u15_u2_U73 (.A2( u1_u15_X_15 ) , .A1( u1_u15_X_18 ) , .ZN( u1_u15_u2_n104 ) );
  NOR2_X1 u1_u15_u2_U74 (.A2( u1_u15_X_14 ) , .ZN( u1_u15_u2_n103 ) , .A1( u1_u15_u2_n174 ) );
  NOR2_X1 u1_u15_u2_U75 (.A2( u1_u15_X_15 ) , .ZN( u1_u15_u2_n102 ) , .A1( u1_u15_u2_n165 ) );
  NOR2_X1 u1_u15_u2_U76 (.A2( u1_u15_X_17 ) , .ZN( u1_u15_u2_n114 ) , .A1( u1_u15_u2_n169 ) );
  AND2_X1 u1_u15_u2_U77 (.A1( u1_u15_X_15 ) , .ZN( u1_u15_u2_n105 ) , .A2( u1_u15_u2_n165 ) );
  AND2_X1 u1_u15_u2_U78 (.A2( u1_u15_X_15 ) , .A1( u1_u15_X_18 ) , .ZN( u1_u15_u2_n107 ) );
  AND2_X1 u1_u15_u2_U79 (.A1( u1_u15_X_14 ) , .ZN( u1_u15_u2_n106 ) , .A2( u1_u15_u2_n174 ) );
  AOI21_X1 u1_u15_u2_U8 (.B2( u1_u15_u2_n120 ) , .B1( u1_u15_u2_n121 ) , .ZN( u1_u15_u2_n126 ) , .A( u1_u15_u2_n167 ) );
  AND2_X1 u1_u15_u2_U80 (.A1( u1_u15_X_13 ) , .A2( u1_u15_X_14 ) , .ZN( u1_u15_u2_n108 ) );
  INV_X1 u1_u15_u2_U81 (.A( u1_u15_X_16 ) , .ZN( u1_u15_u2_n169 ) );
  INV_X1 u1_u15_u2_U82 (.A( u1_u15_X_17 ) , .ZN( u1_u15_u2_n166 ) );
  INV_X1 u1_u15_u2_U83 (.A( u1_u15_X_13 ) , .ZN( u1_u15_u2_n174 ) );
  INV_X1 u1_u15_u2_U84 (.A( u1_u15_X_18 ) , .ZN( u1_u15_u2_n165 ) );
  NAND4_X1 u1_u15_u2_U85 (.ZN( u1_out15_30 ) , .A4( u1_u15_u2_n147 ) , .A3( u1_u15_u2_n148 ) , .A2( u1_u15_u2_n149 ) , .A1( u1_u15_u2_n187 ) );
  NOR3_X1 u1_u15_u2_U86 (.A3( u1_u15_u2_n144 ) , .A2( u1_u15_u2_n145 ) , .A1( u1_u15_u2_n146 ) , .ZN( u1_u15_u2_n147 ) );
  AOI21_X1 u1_u15_u2_U87 (.B2( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n148 ) , .A( u1_u15_u2_n162 ) , .B1( u1_u15_u2_n182 ) );
  NAND4_X1 u1_u15_u2_U88 (.ZN( u1_out15_24 ) , .A4( u1_u15_u2_n111 ) , .A3( u1_u15_u2_n112 ) , .A1( u1_u15_u2_n130 ) , .A2( u1_u15_u2_n187 ) );
  AOI221_X1 u1_u15_u2_U89 (.A( u1_u15_u2_n109 ) , .B1( u1_u15_u2_n110 ) , .ZN( u1_u15_u2_n111 ) , .C1( u1_u15_u2_n134 ) , .C2( u1_u15_u2_n170 ) , .B2( u1_u15_u2_n173 ) );
  OAI22_X1 u1_u15_u2_U9 (.ZN( u1_u15_u2_n109 ) , .A2( u1_u15_u2_n113 ) , .B2( u1_u15_u2_n133 ) , .B1( u1_u15_u2_n167 ) , .A1( u1_u15_u2_n168 ) );
  AOI21_X1 u1_u15_u2_U90 (.ZN( u1_u15_u2_n112 ) , .B2( u1_u15_u2_n156 ) , .A( u1_u15_u2_n164 ) , .B1( u1_u15_u2_n181 ) );
  NAND4_X1 u1_u15_u2_U91 (.ZN( u1_out15_16 ) , .A4( u1_u15_u2_n128 ) , .A3( u1_u15_u2_n129 ) , .A1( u1_u15_u2_n130 ) , .A2( u1_u15_u2_n186 ) );
  AOI22_X1 u1_u15_u2_U92 (.A2( u1_u15_u2_n118 ) , .ZN( u1_u15_u2_n129 ) , .A1( u1_u15_u2_n140 ) , .B1( u1_u15_u2_n157 ) , .B2( u1_u15_u2_n170 ) );
  INV_X1 u1_u15_u2_U93 (.A( u1_u15_u2_n163 ) , .ZN( u1_u15_u2_n186 ) );
  OR4_X1 u1_u15_u2_U94 (.ZN( u1_out15_6 ) , .A4( u1_u15_u2_n161 ) , .A3( u1_u15_u2_n162 ) , .A2( u1_u15_u2_n163 ) , .A1( u1_u15_u2_n164 ) );
  OR3_X1 u1_u15_u2_U95 (.A2( u1_u15_u2_n159 ) , .A1( u1_u15_u2_n160 ) , .ZN( u1_u15_u2_n161 ) , .A3( u1_u15_u2_n183 ) );
  AOI21_X1 u1_u15_u2_U96 (.B2( u1_u15_u2_n154 ) , .B1( u1_u15_u2_n155 ) , .ZN( u1_u15_u2_n159 ) , .A( u1_u15_u2_n167 ) );
  NAND3_X1 u1_u15_u2_U97 (.A2( u1_u15_u2_n117 ) , .A1( u1_u15_u2_n122 ) , .A3( u1_u15_u2_n123 ) , .ZN( u1_u15_u2_n134 ) );
  NAND3_X1 u1_u15_u2_U98 (.ZN( u1_u15_u2_n110 ) , .A2( u1_u15_u2_n131 ) , .A3( u1_u15_u2_n139 ) , .A1( u1_u15_u2_n154 ) );
  NAND3_X1 u1_u15_u2_U99 (.A2( u1_u15_u2_n100 ) , .ZN( u1_u15_u2_n101 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n114 ) );
  OAI22_X1 u1_u15_u3_U10 (.B1( u1_u15_u3_n113 ) , .A2( u1_u15_u3_n135 ) , .A1( u1_u15_u3_n150 ) , .B2( u1_u15_u3_n164 ) , .ZN( u1_u15_u3_n98 ) );
  OAI211_X1 u1_u15_u3_U11 (.B( u1_u15_u3_n106 ) , .ZN( u1_u15_u3_n119 ) , .C2( u1_u15_u3_n128 ) , .C1( u1_u15_u3_n167 ) , .A( u1_u15_u3_n181 ) );
  AOI221_X1 u1_u15_u3_U12 (.C1( u1_u15_u3_n105 ) , .ZN( u1_u15_u3_n106 ) , .A( u1_u15_u3_n131 ) , .B2( u1_u15_u3_n132 ) , .C2( u1_u15_u3_n133 ) , .B1( u1_u15_u3_n169 ) );
  INV_X1 u1_u15_u3_U13 (.ZN( u1_u15_u3_n181 ) , .A( u1_u15_u3_n98 ) );
  NAND2_X1 u1_u15_u3_U14 (.ZN( u1_u15_u3_n105 ) , .A2( u1_u15_u3_n130 ) , .A1( u1_u15_u3_n155 ) );
  AOI22_X1 u1_u15_u3_U15 (.B1( u1_u15_u3_n115 ) , .A2( u1_u15_u3_n116 ) , .ZN( u1_u15_u3_n123 ) , .B2( u1_u15_u3_n133 ) , .A1( u1_u15_u3_n169 ) );
  NAND2_X1 u1_u15_u3_U16 (.ZN( u1_u15_u3_n116 ) , .A2( u1_u15_u3_n151 ) , .A1( u1_u15_u3_n182 ) );
  NOR2_X1 u1_u15_u3_U17 (.ZN( u1_u15_u3_n126 ) , .A2( u1_u15_u3_n150 ) , .A1( u1_u15_u3_n164 ) );
  AOI21_X1 u1_u15_u3_U18 (.ZN( u1_u15_u3_n112 ) , .B2( u1_u15_u3_n146 ) , .B1( u1_u15_u3_n155 ) , .A( u1_u15_u3_n167 ) );
  NAND2_X1 u1_u15_u3_U19 (.A1( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n142 ) , .A2( u1_u15_u3_n164 ) );
  NAND2_X1 u1_u15_u3_U20 (.ZN( u1_u15_u3_n132 ) , .A2( u1_u15_u3_n152 ) , .A1( u1_u15_u3_n156 ) );
  AND2_X1 u1_u15_u3_U21 (.A2( u1_u15_u3_n113 ) , .A1( u1_u15_u3_n114 ) , .ZN( u1_u15_u3_n151 ) );
  INV_X1 u1_u15_u3_U22 (.A( u1_u15_u3_n133 ) , .ZN( u1_u15_u3_n165 ) );
  INV_X1 u1_u15_u3_U23 (.A( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n170 ) );
  NAND2_X1 u1_u15_u3_U24 (.A1( u1_u15_u3_n107 ) , .A2( u1_u15_u3_n108 ) , .ZN( u1_u15_u3_n140 ) );
  NAND2_X1 u1_u15_u3_U25 (.ZN( u1_u15_u3_n117 ) , .A1( u1_u15_u3_n124 ) , .A2( u1_u15_u3_n148 ) );
  NAND2_X1 u1_u15_u3_U26 (.ZN( u1_u15_u3_n143 ) , .A1( u1_u15_u3_n165 ) , .A2( u1_u15_u3_n167 ) );
  INV_X1 u1_u15_u3_U27 (.A( u1_u15_u3_n130 ) , .ZN( u1_u15_u3_n177 ) );
  INV_X1 u1_u15_u3_U28 (.A( u1_u15_u3_n128 ) , .ZN( u1_u15_u3_n176 ) );
  INV_X1 u1_u15_u3_U29 (.A( u1_u15_u3_n155 ) , .ZN( u1_u15_u3_n174 ) );
  INV_X1 u1_u15_u3_U3 (.A( u1_u15_u3_n129 ) , .ZN( u1_u15_u3_n183 ) );
  INV_X1 u1_u15_u3_U30 (.A( u1_u15_u3_n139 ) , .ZN( u1_u15_u3_n185 ) );
  NOR2_X1 u1_u15_u3_U31 (.ZN( u1_u15_u3_n135 ) , .A2( u1_u15_u3_n141 ) , .A1( u1_u15_u3_n169 ) );
  OAI222_X1 u1_u15_u3_U32 (.C2( u1_u15_u3_n107 ) , .A2( u1_u15_u3_n108 ) , .B1( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n138 ) , .B2( u1_u15_u3_n146 ) , .C1( u1_u15_u3_n154 ) , .A1( u1_u15_u3_n164 ) );
  NOR4_X1 u1_u15_u3_U33 (.A4( u1_u15_u3_n157 ) , .A3( u1_u15_u3_n158 ) , .A2( u1_u15_u3_n159 ) , .A1( u1_u15_u3_n160 ) , .ZN( u1_u15_u3_n161 ) );
  AOI21_X1 u1_u15_u3_U34 (.B2( u1_u15_u3_n152 ) , .B1( u1_u15_u3_n153 ) , .ZN( u1_u15_u3_n158 ) , .A( u1_u15_u3_n164 ) );
  AOI21_X1 u1_u15_u3_U35 (.A( u1_u15_u3_n154 ) , .B2( u1_u15_u3_n155 ) , .B1( u1_u15_u3_n156 ) , .ZN( u1_u15_u3_n157 ) );
  AOI21_X1 u1_u15_u3_U36 (.A( u1_u15_u3_n149 ) , .B2( u1_u15_u3_n150 ) , .B1( u1_u15_u3_n151 ) , .ZN( u1_u15_u3_n159 ) );
  AOI211_X1 u1_u15_u3_U37 (.ZN( u1_u15_u3_n109 ) , .A( u1_u15_u3_n119 ) , .C2( u1_u15_u3_n129 ) , .B( u1_u15_u3_n138 ) , .C1( u1_u15_u3_n141 ) );
  AOI211_X1 u1_u15_u3_U38 (.B( u1_u15_u3_n119 ) , .A( u1_u15_u3_n120 ) , .C2( u1_u15_u3_n121 ) , .ZN( u1_u15_u3_n122 ) , .C1( u1_u15_u3_n179 ) );
  INV_X1 u1_u15_u3_U39 (.A( u1_u15_u3_n156 ) , .ZN( u1_u15_u3_n179 ) );
  INV_X1 u1_u15_u3_U4 (.A( u1_u15_u3_n140 ) , .ZN( u1_u15_u3_n182 ) );
  OAI22_X1 u1_u15_u3_U40 (.B1( u1_u15_u3_n118 ) , .ZN( u1_u15_u3_n120 ) , .A1( u1_u15_u3_n135 ) , .B2( u1_u15_u3_n154 ) , .A2( u1_u15_u3_n178 ) );
  AND3_X1 u1_u15_u3_U41 (.ZN( u1_u15_u3_n118 ) , .A2( u1_u15_u3_n124 ) , .A1( u1_u15_u3_n144 ) , .A3( u1_u15_u3_n152 ) );
  INV_X1 u1_u15_u3_U42 (.A( u1_u15_u3_n121 ) , .ZN( u1_u15_u3_n164 ) );
  NAND2_X1 u1_u15_u3_U43 (.ZN( u1_u15_u3_n133 ) , .A1( u1_u15_u3_n154 ) , .A2( u1_u15_u3_n164 ) );
  OAI211_X1 u1_u15_u3_U44 (.B( u1_u15_u3_n127 ) , .ZN( u1_u15_u3_n139 ) , .C1( u1_u15_u3_n150 ) , .C2( u1_u15_u3_n154 ) , .A( u1_u15_u3_n184 ) );
  INV_X1 u1_u15_u3_U45 (.A( u1_u15_u3_n125 ) , .ZN( u1_u15_u3_n184 ) );
  AOI221_X1 u1_u15_u3_U46 (.A( u1_u15_u3_n126 ) , .ZN( u1_u15_u3_n127 ) , .C2( u1_u15_u3_n132 ) , .C1( u1_u15_u3_n169 ) , .B2( u1_u15_u3_n170 ) , .B1( u1_u15_u3_n174 ) );
  OAI22_X1 u1_u15_u3_U47 (.A1( u1_u15_u3_n124 ) , .ZN( u1_u15_u3_n125 ) , .B2( u1_u15_u3_n145 ) , .A2( u1_u15_u3_n165 ) , .B1( u1_u15_u3_n167 ) );
  NOR2_X1 u1_u15_u3_U48 (.A1( u1_u15_u3_n113 ) , .ZN( u1_u15_u3_n131 ) , .A2( u1_u15_u3_n154 ) );
  NAND2_X1 u1_u15_u3_U49 (.A1( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n150 ) , .A2( u1_u15_u3_n99 ) );
  INV_X1 u1_u15_u3_U5 (.A( u1_u15_u3_n117 ) , .ZN( u1_u15_u3_n178 ) );
  NAND2_X1 u1_u15_u3_U50 (.A2( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n155 ) , .A1( u1_u15_u3_n97 ) );
  INV_X1 u1_u15_u3_U51 (.A( u1_u15_u3_n141 ) , .ZN( u1_u15_u3_n167 ) );
  AOI21_X1 u1_u15_u3_U52 (.B2( u1_u15_u3_n114 ) , .B1( u1_u15_u3_n146 ) , .A( u1_u15_u3_n154 ) , .ZN( u1_u15_u3_n94 ) );
  AOI21_X1 u1_u15_u3_U53 (.ZN( u1_u15_u3_n110 ) , .B2( u1_u15_u3_n142 ) , .B1( u1_u15_u3_n186 ) , .A( u1_u15_u3_n95 ) );
  INV_X1 u1_u15_u3_U54 (.A( u1_u15_u3_n145 ) , .ZN( u1_u15_u3_n186 ) );
  AOI21_X1 u1_u15_u3_U55 (.B1( u1_u15_u3_n124 ) , .A( u1_u15_u3_n149 ) , .B2( u1_u15_u3_n155 ) , .ZN( u1_u15_u3_n95 ) );
  INV_X1 u1_u15_u3_U56 (.A( u1_u15_u3_n149 ) , .ZN( u1_u15_u3_n169 ) );
  NAND2_X1 u1_u15_u3_U57 (.ZN( u1_u15_u3_n124 ) , .A1( u1_u15_u3_n96 ) , .A2( u1_u15_u3_n97 ) );
  NAND2_X1 u1_u15_u3_U58 (.A2( u1_u15_u3_n100 ) , .ZN( u1_u15_u3_n146 ) , .A1( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U59 (.A1( u1_u15_u3_n101 ) , .ZN( u1_u15_u3_n145 ) , .A2( u1_u15_u3_n99 ) );
  AOI221_X1 u1_u15_u3_U6 (.A( u1_u15_u3_n131 ) , .C2( u1_u15_u3_n132 ) , .C1( u1_u15_u3_n133 ) , .ZN( u1_u15_u3_n134 ) , .B1( u1_u15_u3_n143 ) , .B2( u1_u15_u3_n177 ) );
  NAND2_X1 u1_u15_u3_U60 (.A1( u1_u15_u3_n100 ) , .ZN( u1_u15_u3_n156 ) , .A2( u1_u15_u3_n99 ) );
  NAND2_X1 u1_u15_u3_U61 (.A2( u1_u15_u3_n101 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n148 ) );
  NAND2_X1 u1_u15_u3_U62 (.A1( u1_u15_u3_n100 ) , .A2( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n128 ) );
  NAND2_X1 u1_u15_u3_U63 (.A2( u1_u15_u3_n101 ) , .A1( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n152 ) );
  NAND2_X1 u1_u15_u3_U64 (.A2( u1_u15_u3_n101 ) , .ZN( u1_u15_u3_n114 ) , .A1( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U65 (.ZN( u1_u15_u3_n107 ) , .A1( u1_u15_u3_n97 ) , .A2( u1_u15_u3_n99 ) );
  NAND2_X1 u1_u15_u3_U66 (.A2( u1_u15_u3_n100 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n113 ) );
  NAND2_X1 u1_u15_u3_U67 (.A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n153 ) , .A2( u1_u15_u3_n97 ) );
  NAND2_X1 u1_u15_u3_U68 (.A2( u1_u15_u3_n103 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n130 ) );
  NAND2_X1 u1_u15_u3_U69 (.A2( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n144 ) , .A1( u1_u15_u3_n96 ) );
  OAI22_X1 u1_u15_u3_U7 (.B2( u1_u15_u3_n147 ) , .A2( u1_u15_u3_n148 ) , .ZN( u1_u15_u3_n160 ) , .B1( u1_u15_u3_n165 ) , .A1( u1_u15_u3_n168 ) );
  NAND2_X1 u1_u15_u3_U70 (.A1( u1_u15_u3_n102 ) , .A2( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n108 ) );
  NOR2_X1 u1_u15_u3_U71 (.A2( u1_u15_X_19 ) , .A1( u1_u15_X_20 ) , .ZN( u1_u15_u3_n99 ) );
  NOR2_X1 u1_u15_u3_U72 (.A2( u1_u15_X_21 ) , .A1( u1_u15_X_24 ) , .ZN( u1_u15_u3_n103 ) );
  NOR2_X1 u1_u15_u3_U73 (.A2( u1_u15_X_24 ) , .A1( u1_u15_u3_n171 ) , .ZN( u1_u15_u3_n97 ) );
  NOR2_X1 u1_u15_u3_U74 (.A2( u1_u15_X_23 ) , .ZN( u1_u15_u3_n141 ) , .A1( u1_u15_u3_n166 ) );
  NOR2_X1 u1_u15_u3_U75 (.A2( u1_u15_X_19 ) , .A1( u1_u15_u3_n172 ) , .ZN( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U76 (.A1( u1_u15_X_22 ) , .A2( u1_u15_X_23 ) , .ZN( u1_u15_u3_n154 ) );
  NAND2_X1 u1_u15_u3_U77 (.A1( u1_u15_X_23 ) , .ZN( u1_u15_u3_n149 ) , .A2( u1_u15_u3_n166 ) );
  NOR2_X1 u1_u15_u3_U78 (.A2( u1_u15_X_22 ) , .A1( u1_u15_X_23 ) , .ZN( u1_u15_u3_n121 ) );
  AND2_X1 u1_u15_u3_U79 (.A1( u1_u15_X_24 ) , .ZN( u1_u15_u3_n101 ) , .A2( u1_u15_u3_n171 ) );
  AND3_X1 u1_u15_u3_U8 (.A3( u1_u15_u3_n144 ) , .A2( u1_u15_u3_n145 ) , .A1( u1_u15_u3_n146 ) , .ZN( u1_u15_u3_n147 ) );
  AND2_X1 u1_u15_u3_U80 (.A1( u1_u15_X_19 ) , .ZN( u1_u15_u3_n102 ) , .A2( u1_u15_u3_n172 ) );
  AND2_X1 u1_u15_u3_U81 (.A1( u1_u15_X_21 ) , .A2( u1_u15_X_24 ) , .ZN( u1_u15_u3_n100 ) );
  AND2_X1 u1_u15_u3_U82 (.A2( u1_u15_X_19 ) , .A1( u1_u15_X_20 ) , .ZN( u1_u15_u3_n104 ) );
  INV_X1 u1_u15_u3_U83 (.A( u1_u15_X_22 ) , .ZN( u1_u15_u3_n166 ) );
  INV_X1 u1_u15_u3_U84 (.A( u1_u15_X_21 ) , .ZN( u1_u15_u3_n171 ) );
  INV_X1 u1_u15_u3_U85 (.A( u1_u15_X_20 ) , .ZN( u1_u15_u3_n172 ) );
  OR4_X1 u1_u15_u3_U86 (.ZN( u1_out15_10 ) , .A4( u1_u15_u3_n136 ) , .A3( u1_u15_u3_n137 ) , .A1( u1_u15_u3_n138 ) , .A2( u1_u15_u3_n139 ) );
  OAI222_X1 u1_u15_u3_U87 (.C1( u1_u15_u3_n128 ) , .ZN( u1_u15_u3_n137 ) , .B1( u1_u15_u3_n148 ) , .A2( u1_u15_u3_n150 ) , .B2( u1_u15_u3_n154 ) , .C2( u1_u15_u3_n164 ) , .A1( u1_u15_u3_n167 ) );
  OAI221_X1 u1_u15_u3_U88 (.A( u1_u15_u3_n134 ) , .B2( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n136 ) , .C1( u1_u15_u3_n149 ) , .B1( u1_u15_u3_n151 ) , .C2( u1_u15_u3_n183 ) );
  NAND4_X1 u1_u15_u3_U89 (.ZN( u1_out15_1 ) , .A4( u1_u15_u3_n161 ) , .A3( u1_u15_u3_n162 ) , .A2( u1_u15_u3_n163 ) , .A1( u1_u15_u3_n185 ) );
  INV_X1 u1_u15_u3_U9 (.A( u1_u15_u3_n143 ) , .ZN( u1_u15_u3_n168 ) );
  NAND2_X1 u1_u15_u3_U90 (.ZN( u1_u15_u3_n163 ) , .A2( u1_u15_u3_n170 ) , .A1( u1_u15_u3_n176 ) );
  AOI22_X1 u1_u15_u3_U91 (.B2( u1_u15_u3_n140 ) , .B1( u1_u15_u3_n141 ) , .A2( u1_u15_u3_n142 ) , .ZN( u1_u15_u3_n162 ) , .A1( u1_u15_u3_n177 ) );
  NAND4_X1 u1_u15_u3_U92 (.ZN( u1_out15_26 ) , .A4( u1_u15_u3_n109 ) , .A3( u1_u15_u3_n110 ) , .A2( u1_u15_u3_n111 ) , .A1( u1_u15_u3_n173 ) );
  INV_X1 u1_u15_u3_U93 (.ZN( u1_u15_u3_n173 ) , .A( u1_u15_u3_n94 ) );
  OAI21_X1 u1_u15_u3_U94 (.ZN( u1_u15_u3_n111 ) , .B2( u1_u15_u3_n117 ) , .A( u1_u15_u3_n133 ) , .B1( u1_u15_u3_n176 ) );
  NAND4_X1 u1_u15_u3_U95 (.ZN( u1_out15_20 ) , .A4( u1_u15_u3_n122 ) , .A3( u1_u15_u3_n123 ) , .A1( u1_u15_u3_n175 ) , .A2( u1_u15_u3_n180 ) );
  INV_X1 u1_u15_u3_U96 (.A( u1_u15_u3_n126 ) , .ZN( u1_u15_u3_n180 ) );
  INV_X1 u1_u15_u3_U97 (.A( u1_u15_u3_n112 ) , .ZN( u1_u15_u3_n175 ) );
  NAND3_X1 u1_u15_u3_U98 (.A1( u1_u15_u3_n114 ) , .ZN( u1_u15_u3_n115 ) , .A2( u1_u15_u3_n145 ) , .A3( u1_u15_u3_n153 ) );
  NAND3_X1 u1_u15_u3_U99 (.ZN( u1_u15_u3_n129 ) , .A2( u1_u15_u3_n144 ) , .A1( u1_u15_u3_n153 ) , .A3( u1_u15_u3_n182 ) );
  OAI22_X1 u1_u15_u4_U10 (.B2( u1_u15_u4_n135 ) , .ZN( u1_u15_u4_n137 ) , .B1( u1_u15_u4_n153 ) , .A1( u1_u15_u4_n155 ) , .A2( u1_u15_u4_n171 ) );
  AND3_X1 u1_u15_u4_U11 (.A2( u1_u15_u4_n134 ) , .ZN( u1_u15_u4_n135 ) , .A3( u1_u15_u4_n145 ) , .A1( u1_u15_u4_n157 ) );
  NAND2_X1 u1_u15_u4_U12 (.ZN( u1_u15_u4_n132 ) , .A2( u1_u15_u4_n170 ) , .A1( u1_u15_u4_n173 ) );
  AOI21_X1 u1_u15_u4_U13 (.B2( u1_u15_u4_n160 ) , .B1( u1_u15_u4_n161 ) , .ZN( u1_u15_u4_n162 ) , .A( u1_u15_u4_n170 ) );
  AOI21_X1 u1_u15_u4_U14 (.ZN( u1_u15_u4_n107 ) , .B2( u1_u15_u4_n143 ) , .A( u1_u15_u4_n174 ) , .B1( u1_u15_u4_n184 ) );
  AOI21_X1 u1_u15_u4_U15 (.B2( u1_u15_u4_n158 ) , .B1( u1_u15_u4_n159 ) , .ZN( u1_u15_u4_n163 ) , .A( u1_u15_u4_n174 ) );
  AOI21_X1 u1_u15_u4_U16 (.A( u1_u15_u4_n153 ) , .B2( u1_u15_u4_n154 ) , .B1( u1_u15_u4_n155 ) , .ZN( u1_u15_u4_n165 ) );
  AOI21_X1 u1_u15_u4_U17 (.A( u1_u15_u4_n156 ) , .B2( u1_u15_u4_n157 ) , .ZN( u1_u15_u4_n164 ) , .B1( u1_u15_u4_n184 ) );
  INV_X1 u1_u15_u4_U18 (.A( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n170 ) );
  AND2_X1 u1_u15_u4_U19 (.A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n155 ) , .A1( u1_u15_u4_n160 ) );
  INV_X1 u1_u15_u4_U20 (.A( u1_u15_u4_n156 ) , .ZN( u1_u15_u4_n175 ) );
  NAND2_X1 u1_u15_u4_U21 (.A2( u1_u15_u4_n118 ) , .ZN( u1_u15_u4_n131 ) , .A1( u1_u15_u4_n147 ) );
  NAND2_X1 u1_u15_u4_U22 (.A1( u1_u15_u4_n119 ) , .A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n130 ) );
  NAND2_X1 u1_u15_u4_U23 (.ZN( u1_u15_u4_n117 ) , .A2( u1_u15_u4_n118 ) , .A1( u1_u15_u4_n148 ) );
  NAND2_X1 u1_u15_u4_U24 (.ZN( u1_u15_u4_n129 ) , .A1( u1_u15_u4_n134 ) , .A2( u1_u15_u4_n148 ) );
  AND3_X1 u1_u15_u4_U25 (.A1( u1_u15_u4_n119 ) , .A2( u1_u15_u4_n143 ) , .A3( u1_u15_u4_n154 ) , .ZN( u1_u15_u4_n161 ) );
  AND2_X1 u1_u15_u4_U26 (.A1( u1_u15_u4_n145 ) , .A2( u1_u15_u4_n147 ) , .ZN( u1_u15_u4_n159 ) );
  OR3_X1 u1_u15_u4_U27 (.A3( u1_u15_u4_n114 ) , .A2( u1_u15_u4_n115 ) , .A1( u1_u15_u4_n116 ) , .ZN( u1_u15_u4_n136 ) );
  AOI21_X1 u1_u15_u4_U28 (.A( u1_u15_u4_n113 ) , .ZN( u1_u15_u4_n116 ) , .B2( u1_u15_u4_n173 ) , .B1( u1_u15_u4_n174 ) );
  AOI21_X1 u1_u15_u4_U29 (.ZN( u1_u15_u4_n115 ) , .B2( u1_u15_u4_n145 ) , .B1( u1_u15_u4_n146 ) , .A( u1_u15_u4_n156 ) );
  NOR2_X1 u1_u15_u4_U3 (.ZN( u1_u15_u4_n121 ) , .A1( u1_u15_u4_n181 ) , .A2( u1_u15_u4_n182 ) );
  OAI22_X1 u1_u15_u4_U30 (.ZN( u1_u15_u4_n114 ) , .A2( u1_u15_u4_n121 ) , .B1( u1_u15_u4_n160 ) , .B2( u1_u15_u4_n170 ) , .A1( u1_u15_u4_n171 ) );
  INV_X1 u1_u15_u4_U31 (.A( u1_u15_u4_n158 ) , .ZN( u1_u15_u4_n182 ) );
  INV_X1 u1_u15_u4_U32 (.ZN( u1_u15_u4_n181 ) , .A( u1_u15_u4_n96 ) );
  INV_X1 u1_u15_u4_U33 (.A( u1_u15_u4_n144 ) , .ZN( u1_u15_u4_n179 ) );
  INV_X1 u1_u15_u4_U34 (.A( u1_u15_u4_n157 ) , .ZN( u1_u15_u4_n178 ) );
  NAND2_X1 u1_u15_u4_U35 (.A2( u1_u15_u4_n154 ) , .A1( u1_u15_u4_n96 ) , .ZN( u1_u15_u4_n97 ) );
  INV_X1 u1_u15_u4_U36 (.ZN( u1_u15_u4_n186 ) , .A( u1_u15_u4_n95 ) );
  OAI221_X1 u1_u15_u4_U37 (.C1( u1_u15_u4_n134 ) , .B1( u1_u15_u4_n158 ) , .B2( u1_u15_u4_n171 ) , .C2( u1_u15_u4_n173 ) , .A( u1_u15_u4_n94 ) , .ZN( u1_u15_u4_n95 ) );
  AOI222_X1 u1_u15_u4_U38 (.B2( u1_u15_u4_n132 ) , .A1( u1_u15_u4_n138 ) , .C2( u1_u15_u4_n175 ) , .A2( u1_u15_u4_n179 ) , .C1( u1_u15_u4_n181 ) , .B1( u1_u15_u4_n185 ) , .ZN( u1_u15_u4_n94 ) );
  INV_X1 u1_u15_u4_U39 (.A( u1_u15_u4_n113 ) , .ZN( u1_u15_u4_n185 ) );
  INV_X1 u1_u15_u4_U4 (.A( u1_u15_u4_n117 ) , .ZN( u1_u15_u4_n184 ) );
  INV_X1 u1_u15_u4_U40 (.A( u1_u15_u4_n143 ) , .ZN( u1_u15_u4_n183 ) );
  NOR2_X1 u1_u15_u4_U41 (.ZN( u1_u15_u4_n138 ) , .A1( u1_u15_u4_n168 ) , .A2( u1_u15_u4_n169 ) );
  NOR2_X1 u1_u15_u4_U42 (.A1( u1_u15_u4_n150 ) , .A2( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n153 ) );
  NOR2_X1 u1_u15_u4_U43 (.A2( u1_u15_u4_n128 ) , .A1( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n156 ) );
  AOI22_X1 u1_u15_u4_U44 (.B2( u1_u15_u4_n122 ) , .A1( u1_u15_u4_n123 ) , .ZN( u1_u15_u4_n124 ) , .B1( u1_u15_u4_n128 ) , .A2( u1_u15_u4_n172 ) );
  NAND2_X1 u1_u15_u4_U45 (.A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n123 ) , .A1( u1_u15_u4_n161 ) );
  INV_X1 u1_u15_u4_U46 (.A( u1_u15_u4_n153 ) , .ZN( u1_u15_u4_n172 ) );
  AOI22_X1 u1_u15_u4_U47 (.B2( u1_u15_u4_n132 ) , .A2( u1_u15_u4_n133 ) , .ZN( u1_u15_u4_n140 ) , .A1( u1_u15_u4_n150 ) , .B1( u1_u15_u4_n179 ) );
  NAND2_X1 u1_u15_u4_U48 (.ZN( u1_u15_u4_n133 ) , .A2( u1_u15_u4_n146 ) , .A1( u1_u15_u4_n154 ) );
  NAND2_X1 u1_u15_u4_U49 (.A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n154 ) , .A2( u1_u15_u4_n98 ) );
  NOR4_X1 u1_u15_u4_U5 (.A4( u1_u15_u4_n106 ) , .A3( u1_u15_u4_n107 ) , .A2( u1_u15_u4_n108 ) , .A1( u1_u15_u4_n109 ) , .ZN( u1_u15_u4_n110 ) );
  NAND2_X1 u1_u15_u4_U50 (.A1( u1_u15_u4_n101 ) , .ZN( u1_u15_u4_n158 ) , .A2( u1_u15_u4_n99 ) );
  AOI21_X1 u1_u15_u4_U51 (.ZN( u1_u15_u4_n127 ) , .A( u1_u15_u4_n136 ) , .B2( u1_u15_u4_n150 ) , .B1( u1_u15_u4_n180 ) );
  INV_X1 u1_u15_u4_U52 (.A( u1_u15_u4_n160 ) , .ZN( u1_u15_u4_n180 ) );
  NAND2_X1 u1_u15_u4_U53 (.A2( u1_u15_u4_n104 ) , .A1( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n146 ) );
  NAND2_X1 u1_u15_u4_U54 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n160 ) );
  NAND2_X1 u1_u15_u4_U55 (.ZN( u1_u15_u4_n134 ) , .A1( u1_u15_u4_n98 ) , .A2( u1_u15_u4_n99 ) );
  NAND2_X1 u1_u15_u4_U56 (.A1( u1_u15_u4_n103 ) , .A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n143 ) );
  NAND2_X1 u1_u15_u4_U57 (.A2( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n145 ) , .A1( u1_u15_u4_n98 ) );
  NAND2_X1 u1_u15_u4_U58 (.A1( u1_u15_u4_n100 ) , .A2( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n120 ) );
  NAND2_X1 u1_u15_u4_U59 (.A1( u1_u15_u4_n102 ) , .A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n148 ) );
  AOI21_X1 u1_u15_u4_U6 (.ZN( u1_u15_u4_n106 ) , .B2( u1_u15_u4_n146 ) , .B1( u1_u15_u4_n158 ) , .A( u1_u15_u4_n170 ) );
  NAND2_X1 u1_u15_u4_U60 (.A2( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n157 ) );
  INV_X1 u1_u15_u4_U61 (.A( u1_u15_u4_n150 ) , .ZN( u1_u15_u4_n173 ) );
  INV_X1 u1_u15_u4_U62 (.A( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n171 ) );
  NAND2_X1 u1_u15_u4_U63 (.A1( u1_u15_u4_n100 ) , .ZN( u1_u15_u4_n118 ) , .A2( u1_u15_u4_n99 ) );
  NAND2_X1 u1_u15_u4_U64 (.A2( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n144 ) );
  NAND2_X1 u1_u15_u4_U65 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n96 ) );
  INV_X1 u1_u15_u4_U66 (.A( u1_u15_u4_n128 ) , .ZN( u1_u15_u4_n174 ) );
  NAND2_X1 u1_u15_u4_U67 (.A2( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n119 ) , .A1( u1_u15_u4_n98 ) );
  NAND2_X1 u1_u15_u4_U68 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n147 ) );
  NAND2_X1 u1_u15_u4_U69 (.A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n113 ) , .A1( u1_u15_u4_n99 ) );
  AOI21_X1 u1_u15_u4_U7 (.ZN( u1_u15_u4_n108 ) , .B2( u1_u15_u4_n134 ) , .B1( u1_u15_u4_n155 ) , .A( u1_u15_u4_n156 ) );
  NOR2_X1 u1_u15_u4_U70 (.A2( u1_u15_X_28 ) , .ZN( u1_u15_u4_n150 ) , .A1( u1_u15_u4_n168 ) );
  NOR2_X1 u1_u15_u4_U71 (.A2( u1_u15_X_29 ) , .ZN( u1_u15_u4_n152 ) , .A1( u1_u15_u4_n169 ) );
  NOR2_X1 u1_u15_u4_U72 (.A2( u1_u15_X_26 ) , .ZN( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n177 ) );
  NOR2_X1 u1_u15_u4_U73 (.A2( u1_u15_X_30 ) , .ZN( u1_u15_u4_n105 ) , .A1( u1_u15_u4_n176 ) );
  NOR2_X1 u1_u15_u4_U74 (.A2( u1_u15_X_28 ) , .A1( u1_u15_X_29 ) , .ZN( u1_u15_u4_n128 ) );
  NOR2_X1 u1_u15_u4_U75 (.A2( u1_u15_X_25 ) , .A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n98 ) );
  NOR2_X1 u1_u15_u4_U76 (.A2( u1_u15_X_27 ) , .A1( u1_u15_X_30 ) , .ZN( u1_u15_u4_n102 ) );
  AND2_X1 u1_u15_u4_U77 (.A2( u1_u15_X_25 ) , .A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n104 ) );
  AND2_X1 u1_u15_u4_U78 (.A1( u1_u15_X_30 ) , .A2( u1_u15_u4_n176 ) , .ZN( u1_u15_u4_n99 ) );
  AND2_X1 u1_u15_u4_U79 (.A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n101 ) , .A2( u1_u15_u4_n177 ) );
  AOI21_X1 u1_u15_u4_U8 (.ZN( u1_u15_u4_n109 ) , .A( u1_u15_u4_n153 ) , .B1( u1_u15_u4_n159 ) , .B2( u1_u15_u4_n184 ) );
  AND2_X1 u1_u15_u4_U80 (.A1( u1_u15_X_27 ) , .A2( u1_u15_X_30 ) , .ZN( u1_u15_u4_n103 ) );
  INV_X1 u1_u15_u4_U81 (.A( u1_u15_X_28 ) , .ZN( u1_u15_u4_n169 ) );
  INV_X1 u1_u15_u4_U82 (.A( u1_u15_X_29 ) , .ZN( u1_u15_u4_n168 ) );
  INV_X1 u1_u15_u4_U83 (.A( u1_u15_X_25 ) , .ZN( u1_u15_u4_n177 ) );
  INV_X1 u1_u15_u4_U84 (.A( u1_u15_X_27 ) , .ZN( u1_u15_u4_n176 ) );
  NAND4_X1 u1_u15_u4_U85 (.ZN( u1_out15_25 ) , .A4( u1_u15_u4_n139 ) , .A3( u1_u15_u4_n140 ) , .A2( u1_u15_u4_n141 ) , .A1( u1_u15_u4_n142 ) );
  OAI21_X1 u1_u15_u4_U86 (.A( u1_u15_u4_n128 ) , .B2( u1_u15_u4_n129 ) , .B1( u1_u15_u4_n130 ) , .ZN( u1_u15_u4_n142 ) );
  OAI21_X1 u1_u15_u4_U87 (.B2( u1_u15_u4_n131 ) , .ZN( u1_u15_u4_n141 ) , .A( u1_u15_u4_n175 ) , .B1( u1_u15_u4_n183 ) );
  NAND4_X1 u1_u15_u4_U88 (.ZN( u1_out15_14 ) , .A4( u1_u15_u4_n124 ) , .A3( u1_u15_u4_n125 ) , .A2( u1_u15_u4_n126 ) , .A1( u1_u15_u4_n127 ) );
  AOI22_X1 u1_u15_u4_U89 (.B2( u1_u15_u4_n117 ) , .ZN( u1_u15_u4_n126 ) , .A1( u1_u15_u4_n129 ) , .B1( u1_u15_u4_n152 ) , .A2( u1_u15_u4_n175 ) );
  AOI211_X1 u1_u15_u4_U9 (.B( u1_u15_u4_n136 ) , .A( u1_u15_u4_n137 ) , .C2( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n139 ) , .C1( u1_u15_u4_n182 ) );
  AOI22_X1 u1_u15_u4_U90 (.ZN( u1_u15_u4_n125 ) , .B2( u1_u15_u4_n131 ) , .A2( u1_u15_u4_n132 ) , .B1( u1_u15_u4_n138 ) , .A1( u1_u15_u4_n178 ) );
  AOI22_X1 u1_u15_u4_U91 (.B2( u1_u15_u4_n149 ) , .B1( u1_u15_u4_n150 ) , .A2( u1_u15_u4_n151 ) , .A1( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n167 ) );
  NOR4_X1 u1_u15_u4_U92 (.A4( u1_u15_u4_n162 ) , .A3( u1_u15_u4_n163 ) , .A2( u1_u15_u4_n164 ) , .A1( u1_u15_u4_n165 ) , .ZN( u1_u15_u4_n166 ) );
  NAND4_X1 u1_u15_u4_U93 (.ZN( u1_out15_8 ) , .A4( u1_u15_u4_n110 ) , .A3( u1_u15_u4_n111 ) , .A2( u1_u15_u4_n112 ) , .A1( u1_u15_u4_n186 ) );
  NAND2_X1 u1_u15_u4_U94 (.ZN( u1_u15_u4_n112 ) , .A2( u1_u15_u4_n130 ) , .A1( u1_u15_u4_n150 ) );
  AOI22_X1 u1_u15_u4_U95 (.ZN( u1_u15_u4_n111 ) , .B2( u1_u15_u4_n132 ) , .A1( u1_u15_u4_n152 ) , .B1( u1_u15_u4_n178 ) , .A2( u1_u15_u4_n97 ) );
  NAND3_X1 u1_u15_u4_U96 (.ZN( u1_out15_3 ) , .A3( u1_u15_u4_n166 ) , .A1( u1_u15_u4_n167 ) , .A2( u1_u15_u4_n186 ) );
  NAND3_X1 u1_u15_u4_U97 (.A3( u1_u15_u4_n146 ) , .A2( u1_u15_u4_n147 ) , .A1( u1_u15_u4_n148 ) , .ZN( u1_u15_u4_n149 ) );
  NAND3_X1 u1_u15_u4_U98 (.A3( u1_u15_u4_n143 ) , .A2( u1_u15_u4_n144 ) , .A1( u1_u15_u4_n145 ) , .ZN( u1_u15_u4_n151 ) );
  NAND3_X1 u1_u15_u4_U99 (.A3( u1_u15_u4_n121 ) , .ZN( u1_u15_u4_n122 ) , .A2( u1_u15_u4_n144 ) , .A1( u1_u15_u4_n154 ) );
  INV_X1 u1_u15_u5_U10 (.A( u1_u15_u5_n121 ) , .ZN( u1_u15_u5_n177 ) );
  AOI222_X1 u1_u15_u5_U100 (.ZN( u1_u15_u5_n113 ) , .A1( u1_u15_u5_n131 ) , .C1( u1_u15_u5_n148 ) , .B2( u1_u15_u5_n174 ) , .C2( u1_u15_u5_n178 ) , .A2( u1_u15_u5_n179 ) , .B1( u1_u15_u5_n99 ) );
  NAND4_X1 u1_u15_u5_U101 (.ZN( u1_out15_29 ) , .A4( u1_u15_u5_n129 ) , .A3( u1_u15_u5_n130 ) , .A2( u1_u15_u5_n168 ) , .A1( u1_u15_u5_n196 ) );
  AOI221_X1 u1_u15_u5_U102 (.A( u1_u15_u5_n128 ) , .ZN( u1_u15_u5_n129 ) , .C2( u1_u15_u5_n132 ) , .B2( u1_u15_u5_n159 ) , .B1( u1_u15_u5_n176 ) , .C1( u1_u15_u5_n184 ) );
  AOI222_X1 u1_u15_u5_U103 (.ZN( u1_u15_u5_n130 ) , .A2( u1_u15_u5_n146 ) , .B1( u1_u15_u5_n147 ) , .C2( u1_u15_u5_n175 ) , .B2( u1_u15_u5_n179 ) , .A1( u1_u15_u5_n188 ) , .C1( u1_u15_u5_n194 ) );
  NAND3_X1 u1_u15_u5_U104 (.A2( u1_u15_u5_n154 ) , .A3( u1_u15_u5_n158 ) , .A1( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n99 ) );
  NOR2_X1 u1_u15_u5_U11 (.ZN( u1_u15_u5_n160 ) , .A2( u1_u15_u5_n173 ) , .A1( u1_u15_u5_n177 ) );
  INV_X1 u1_u15_u5_U12 (.A( u1_u15_u5_n150 ) , .ZN( u1_u15_u5_n174 ) );
  AOI21_X1 u1_u15_u5_U13 (.A( u1_u15_u5_n160 ) , .B2( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n162 ) , .B1( u1_u15_u5_n192 ) );
  INV_X1 u1_u15_u5_U14 (.A( u1_u15_u5_n159 ) , .ZN( u1_u15_u5_n192 ) );
  AOI21_X1 u1_u15_u5_U15 (.A( u1_u15_u5_n156 ) , .B2( u1_u15_u5_n157 ) , .B1( u1_u15_u5_n158 ) , .ZN( u1_u15_u5_n163 ) );
  AOI21_X1 u1_u15_u5_U16 (.B2( u1_u15_u5_n139 ) , .B1( u1_u15_u5_n140 ) , .ZN( u1_u15_u5_n141 ) , .A( u1_u15_u5_n150 ) );
  OAI21_X1 u1_u15_u5_U17 (.A( u1_u15_u5_n133 ) , .B2( u1_u15_u5_n134 ) , .B1( u1_u15_u5_n135 ) , .ZN( u1_u15_u5_n142 ) );
  OAI21_X1 u1_u15_u5_U18 (.ZN( u1_u15_u5_n133 ) , .B2( u1_u15_u5_n147 ) , .A( u1_u15_u5_n173 ) , .B1( u1_u15_u5_n188 ) );
  NAND2_X1 u1_u15_u5_U19 (.A2( u1_u15_u5_n119 ) , .A1( u1_u15_u5_n123 ) , .ZN( u1_u15_u5_n137 ) );
  INV_X1 u1_u15_u5_U20 (.A( u1_u15_u5_n155 ) , .ZN( u1_u15_u5_n194 ) );
  NAND2_X1 u1_u15_u5_U21 (.A1( u1_u15_u5_n121 ) , .ZN( u1_u15_u5_n132 ) , .A2( u1_u15_u5_n172 ) );
  NAND2_X1 u1_u15_u5_U22 (.A2( u1_u15_u5_n122 ) , .ZN( u1_u15_u5_n136 ) , .A1( u1_u15_u5_n154 ) );
  NAND2_X1 u1_u15_u5_U23 (.A2( u1_u15_u5_n119 ) , .A1( u1_u15_u5_n120 ) , .ZN( u1_u15_u5_n159 ) );
  INV_X1 u1_u15_u5_U24 (.A( u1_u15_u5_n156 ) , .ZN( u1_u15_u5_n175 ) );
  INV_X1 u1_u15_u5_U25 (.A( u1_u15_u5_n158 ) , .ZN( u1_u15_u5_n188 ) );
  INV_X1 u1_u15_u5_U26 (.A( u1_u15_u5_n152 ) , .ZN( u1_u15_u5_n179 ) );
  INV_X1 u1_u15_u5_U27 (.A( u1_u15_u5_n140 ) , .ZN( u1_u15_u5_n182 ) );
  INV_X1 u1_u15_u5_U28 (.A( u1_u15_u5_n151 ) , .ZN( u1_u15_u5_n183 ) );
  INV_X1 u1_u15_u5_U29 (.A( u1_u15_u5_n123 ) , .ZN( u1_u15_u5_n185 ) );
  NOR2_X1 u1_u15_u5_U3 (.ZN( u1_u15_u5_n134 ) , .A1( u1_u15_u5_n183 ) , .A2( u1_u15_u5_n190 ) );
  INV_X1 u1_u15_u5_U30 (.A( u1_u15_u5_n161 ) , .ZN( u1_u15_u5_n184 ) );
  INV_X1 u1_u15_u5_U31 (.A( u1_u15_u5_n139 ) , .ZN( u1_u15_u5_n189 ) );
  INV_X1 u1_u15_u5_U32 (.A( u1_u15_u5_n157 ) , .ZN( u1_u15_u5_n190 ) );
  INV_X1 u1_u15_u5_U33 (.A( u1_u15_u5_n120 ) , .ZN( u1_u15_u5_n193 ) );
  NAND2_X1 u1_u15_u5_U34 (.ZN( u1_u15_u5_n111 ) , .A1( u1_u15_u5_n140 ) , .A2( u1_u15_u5_n155 ) );
  NOR2_X1 u1_u15_u5_U35 (.ZN( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n170 ) , .A2( u1_u15_u5_n180 ) );
  INV_X1 u1_u15_u5_U36 (.A( u1_u15_u5_n117 ) , .ZN( u1_u15_u5_n196 ) );
  OAI221_X1 u1_u15_u5_U37 (.A( u1_u15_u5_n116 ) , .ZN( u1_u15_u5_n117 ) , .B2( u1_u15_u5_n119 ) , .C1( u1_u15_u5_n153 ) , .C2( u1_u15_u5_n158 ) , .B1( u1_u15_u5_n172 ) );
  AOI222_X1 u1_u15_u5_U38 (.ZN( u1_u15_u5_n116 ) , .B2( u1_u15_u5_n145 ) , .C1( u1_u15_u5_n148 ) , .A2( u1_u15_u5_n174 ) , .C2( u1_u15_u5_n177 ) , .B1( u1_u15_u5_n187 ) , .A1( u1_u15_u5_n193 ) );
  INV_X1 u1_u15_u5_U39 (.A( u1_u15_u5_n115 ) , .ZN( u1_u15_u5_n187 ) );
  INV_X1 u1_u15_u5_U4 (.A( u1_u15_u5_n138 ) , .ZN( u1_u15_u5_n191 ) );
  AOI22_X1 u1_u15_u5_U40 (.B2( u1_u15_u5_n131 ) , .A2( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n169 ) , .B1( u1_u15_u5_n174 ) , .A1( u1_u15_u5_n185 ) );
  NOR2_X1 u1_u15_u5_U41 (.A1( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n150 ) , .A2( u1_u15_u5_n173 ) );
  AOI21_X1 u1_u15_u5_U42 (.A( u1_u15_u5_n118 ) , .B2( u1_u15_u5_n145 ) , .ZN( u1_u15_u5_n168 ) , .B1( u1_u15_u5_n186 ) );
  INV_X1 u1_u15_u5_U43 (.A( u1_u15_u5_n122 ) , .ZN( u1_u15_u5_n186 ) );
  NOR2_X1 u1_u15_u5_U44 (.A1( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n152 ) , .A2( u1_u15_u5_n176 ) );
  NOR2_X1 u1_u15_u5_U45 (.A1( u1_u15_u5_n115 ) , .ZN( u1_u15_u5_n118 ) , .A2( u1_u15_u5_n153 ) );
  NOR2_X1 u1_u15_u5_U46 (.A2( u1_u15_u5_n145 ) , .ZN( u1_u15_u5_n156 ) , .A1( u1_u15_u5_n174 ) );
  NOR2_X1 u1_u15_u5_U47 (.ZN( u1_u15_u5_n121 ) , .A2( u1_u15_u5_n145 ) , .A1( u1_u15_u5_n176 ) );
  AOI22_X1 u1_u15_u5_U48 (.ZN( u1_u15_u5_n114 ) , .A2( u1_u15_u5_n137 ) , .A1( u1_u15_u5_n145 ) , .B2( u1_u15_u5_n175 ) , .B1( u1_u15_u5_n193 ) );
  OAI211_X1 u1_u15_u5_U49 (.B( u1_u15_u5_n124 ) , .A( u1_u15_u5_n125 ) , .C2( u1_u15_u5_n126 ) , .C1( u1_u15_u5_n127 ) , .ZN( u1_u15_u5_n128 ) );
  OAI21_X1 u1_u15_u5_U5 (.B2( u1_u15_u5_n136 ) , .B1( u1_u15_u5_n137 ) , .ZN( u1_u15_u5_n138 ) , .A( u1_u15_u5_n177 ) );
  NOR3_X1 u1_u15_u5_U50 (.ZN( u1_u15_u5_n127 ) , .A1( u1_u15_u5_n136 ) , .A3( u1_u15_u5_n148 ) , .A2( u1_u15_u5_n182 ) );
  OAI21_X1 u1_u15_u5_U51 (.ZN( u1_u15_u5_n124 ) , .A( u1_u15_u5_n177 ) , .B2( u1_u15_u5_n183 ) , .B1( u1_u15_u5_n189 ) );
  OAI21_X1 u1_u15_u5_U52 (.ZN( u1_u15_u5_n125 ) , .A( u1_u15_u5_n174 ) , .B2( u1_u15_u5_n185 ) , .B1( u1_u15_u5_n190 ) );
  AOI21_X1 u1_u15_u5_U53 (.A( u1_u15_u5_n153 ) , .B2( u1_u15_u5_n154 ) , .B1( u1_u15_u5_n155 ) , .ZN( u1_u15_u5_n164 ) );
  AOI21_X1 u1_u15_u5_U54 (.ZN( u1_u15_u5_n110 ) , .B1( u1_u15_u5_n122 ) , .B2( u1_u15_u5_n139 ) , .A( u1_u15_u5_n153 ) );
  INV_X1 u1_u15_u5_U55 (.A( u1_u15_u5_n153 ) , .ZN( u1_u15_u5_n176 ) );
  INV_X1 u1_u15_u5_U56 (.A( u1_u15_u5_n126 ) , .ZN( u1_u15_u5_n173 ) );
  AND2_X1 u1_u15_u5_U57 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n147 ) );
  AND2_X1 u1_u15_u5_U58 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n148 ) );
  NAND2_X1 u1_u15_u5_U59 (.A1( u1_u15_u5_n105 ) , .A2( u1_u15_u5_n106 ) , .ZN( u1_u15_u5_n158 ) );
  INV_X1 u1_u15_u5_U6 (.A( u1_u15_u5_n135 ) , .ZN( u1_u15_u5_n178 ) );
  NAND2_X1 u1_u15_u5_U60 (.A2( u1_u15_u5_n108 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n139 ) );
  NAND2_X1 u1_u15_u5_U61 (.A1( u1_u15_u5_n106 ) , .A2( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n119 ) );
  NAND2_X1 u1_u15_u5_U62 (.A2( u1_u15_u5_n103 ) , .A1( u1_u15_u5_n105 ) , .ZN( u1_u15_u5_n140 ) );
  NAND2_X1 u1_u15_u5_U63 (.A2( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n105 ) , .ZN( u1_u15_u5_n155 ) );
  NAND2_X1 u1_u15_u5_U64 (.A2( u1_u15_u5_n106 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n122 ) );
  NAND2_X1 u1_u15_u5_U65 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n106 ) , .ZN( u1_u15_u5_n115 ) );
  NAND2_X1 u1_u15_u5_U66 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n103 ) , .ZN( u1_u15_u5_n161 ) );
  NAND2_X1 u1_u15_u5_U67 (.A1( u1_u15_u5_n105 ) , .A2( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n154 ) );
  INV_X1 u1_u15_u5_U68 (.A( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n172 ) );
  NAND2_X1 u1_u15_u5_U69 (.A1( u1_u15_u5_n103 ) , .A2( u1_u15_u5_n108 ) , .ZN( u1_u15_u5_n123 ) );
  OAI22_X1 u1_u15_u5_U7 (.B2( u1_u15_u5_n149 ) , .B1( u1_u15_u5_n150 ) , .A2( u1_u15_u5_n151 ) , .A1( u1_u15_u5_n152 ) , .ZN( u1_u15_u5_n165 ) );
  NAND2_X1 u1_u15_u5_U70 (.A2( u1_u15_u5_n103 ) , .A1( u1_u15_u5_n107 ) , .ZN( u1_u15_u5_n151 ) );
  NAND2_X1 u1_u15_u5_U71 (.A2( u1_u15_u5_n107 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n120 ) );
  NAND2_X1 u1_u15_u5_U72 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n109 ) , .ZN( u1_u15_u5_n157 ) );
  AND2_X1 u1_u15_u5_U73 (.A2( u1_u15_u5_n100 ) , .A1( u1_u15_u5_n104 ) , .ZN( u1_u15_u5_n131 ) );
  INV_X1 u1_u15_u5_U74 (.A( u1_u15_u5_n102 ) , .ZN( u1_u15_u5_n195 ) );
  OAI221_X1 u1_u15_u5_U75 (.A( u1_u15_u5_n101 ) , .ZN( u1_u15_u5_n102 ) , .C2( u1_u15_u5_n115 ) , .C1( u1_u15_u5_n126 ) , .B1( u1_u15_u5_n134 ) , .B2( u1_u15_u5_n160 ) );
  OAI21_X1 u1_u15_u5_U76 (.ZN( u1_u15_u5_n101 ) , .B1( u1_u15_u5_n137 ) , .A( u1_u15_u5_n146 ) , .B2( u1_u15_u5_n147 ) );
  NOR2_X1 u1_u15_u5_U77 (.A2( u1_u15_X_34 ) , .A1( u1_u15_X_35 ) , .ZN( u1_u15_u5_n145 ) );
  NOR2_X1 u1_u15_u5_U78 (.A2( u1_u15_X_34 ) , .ZN( u1_u15_u5_n146 ) , .A1( u1_u15_u5_n171 ) );
  NOR2_X1 u1_u15_u5_U79 (.A2( u1_u15_X_31 ) , .A1( u1_u15_X_32 ) , .ZN( u1_u15_u5_n103 ) );
  NOR3_X1 u1_u15_u5_U8 (.A2( u1_u15_u5_n147 ) , .A1( u1_u15_u5_n148 ) , .ZN( u1_u15_u5_n149 ) , .A3( u1_u15_u5_n194 ) );
  NOR2_X1 u1_u15_u5_U80 (.A2( u1_u15_X_36 ) , .ZN( u1_u15_u5_n105 ) , .A1( u1_u15_u5_n180 ) );
  NOR2_X1 u1_u15_u5_U81 (.A2( u1_u15_X_33 ) , .ZN( u1_u15_u5_n108 ) , .A1( u1_u15_u5_n170 ) );
  NOR2_X1 u1_u15_u5_U82 (.A2( u1_u15_X_33 ) , .A1( u1_u15_X_36 ) , .ZN( u1_u15_u5_n107 ) );
  NOR2_X1 u1_u15_u5_U83 (.A2( u1_u15_X_31 ) , .ZN( u1_u15_u5_n104 ) , .A1( u1_u15_u5_n181 ) );
  NAND2_X1 u1_u15_u5_U84 (.A2( u1_u15_X_34 ) , .A1( u1_u15_X_35 ) , .ZN( u1_u15_u5_n153 ) );
  NAND2_X1 u1_u15_u5_U85 (.A1( u1_u15_X_34 ) , .ZN( u1_u15_u5_n126 ) , .A2( u1_u15_u5_n171 ) );
  AND2_X1 u1_u15_u5_U86 (.A1( u1_u15_X_31 ) , .A2( u1_u15_X_32 ) , .ZN( u1_u15_u5_n106 ) );
  AND2_X1 u1_u15_u5_U87 (.A1( u1_u15_X_31 ) , .ZN( u1_u15_u5_n109 ) , .A2( u1_u15_u5_n181 ) );
  INV_X1 u1_u15_u5_U88 (.A( u1_u15_X_33 ) , .ZN( u1_u15_u5_n180 ) );
  INV_X1 u1_u15_u5_U89 (.A( u1_u15_X_35 ) , .ZN( u1_u15_u5_n171 ) );
  NOR2_X1 u1_u15_u5_U9 (.ZN( u1_u15_u5_n135 ) , .A1( u1_u15_u5_n173 ) , .A2( u1_u15_u5_n176 ) );
  INV_X1 u1_u15_u5_U90 (.A( u1_u15_X_36 ) , .ZN( u1_u15_u5_n170 ) );
  INV_X1 u1_u15_u5_U91 (.A( u1_u15_X_32 ) , .ZN( u1_u15_u5_n181 ) );
  NAND4_X1 u1_u15_u5_U92 (.ZN( u1_out15_19 ) , .A4( u1_u15_u5_n166 ) , .A3( u1_u15_u5_n167 ) , .A2( u1_u15_u5_n168 ) , .A1( u1_u15_u5_n169 ) );
  AOI22_X1 u1_u15_u5_U93 (.B2( u1_u15_u5_n145 ) , .A2( u1_u15_u5_n146 ) , .ZN( u1_u15_u5_n167 ) , .B1( u1_u15_u5_n182 ) , .A1( u1_u15_u5_n189 ) );
  NOR4_X1 u1_u15_u5_U94 (.A4( u1_u15_u5_n162 ) , .A3( u1_u15_u5_n163 ) , .A2( u1_u15_u5_n164 ) , .A1( u1_u15_u5_n165 ) , .ZN( u1_u15_u5_n166 ) );
  NAND4_X1 u1_u15_u5_U95 (.ZN( u1_out15_11 ) , .A4( u1_u15_u5_n143 ) , .A3( u1_u15_u5_n144 ) , .A2( u1_u15_u5_n169 ) , .A1( u1_u15_u5_n196 ) );
  AOI22_X1 u1_u15_u5_U96 (.A2( u1_u15_u5_n132 ) , .ZN( u1_u15_u5_n144 ) , .B2( u1_u15_u5_n145 ) , .B1( u1_u15_u5_n184 ) , .A1( u1_u15_u5_n194 ) );
  NOR3_X1 u1_u15_u5_U97 (.A3( u1_u15_u5_n141 ) , .A1( u1_u15_u5_n142 ) , .ZN( u1_u15_u5_n143 ) , .A2( u1_u15_u5_n191 ) );
  NAND4_X1 u1_u15_u5_U98 (.ZN( u1_out15_4 ) , .A4( u1_u15_u5_n112 ) , .A2( u1_u15_u5_n113 ) , .A1( u1_u15_u5_n114 ) , .A3( u1_u15_u5_n195 ) );
  AOI211_X1 u1_u15_u5_U99 (.A( u1_u15_u5_n110 ) , .C1( u1_u15_u5_n111 ) , .ZN( u1_u15_u5_n112 ) , .B( u1_u15_u5_n118 ) , .C2( u1_u15_u5_n177 ) );
  XOR2_X1 u1_u1_U11 (.B( u1_K2_44 ) , .A( u1_R0_29 ) , .Z( u1_u1_X_44 ) );
  XOR2_X1 u1_u1_U12 (.B( u1_K2_43 ) , .A( u1_R0_28 ) , .Z( u1_u1_X_43 ) );
  XOR2_X1 u1_u1_U13 (.B( u1_K2_42 ) , .A( u1_R0_29 ) , .Z( u1_u1_X_42 ) );
  XOR2_X1 u1_u1_U14 (.B( u1_K2_41 ) , .A( u1_R0_28 ) , .Z( u1_u1_X_41 ) );
  XOR2_X1 u1_u1_U26 (.B( u1_K2_30 ) , .A( u1_R0_21 ) , .Z( u1_u1_X_30 ) );
  XOR2_X1 u1_u1_U28 (.B( u1_K2_29 ) , .A( u1_R0_20 ) , .Z( u1_u1_X_29 ) );
  XOR2_X1 u1_u1_U31 (.B( u1_K2_26 ) , .A( u1_R0_17 ) , .Z( u1_u1_X_26 ) );
  XOR2_X1 u1_u1_U32 (.B( u1_K2_25 ) , .A( u1_R0_16 ) , .Z( u1_u1_X_25 ) );
  XOR2_X1 u1_u1_U33 (.B( u1_K2_24 ) , .A( u1_R0_17 ) , .Z( u1_u1_X_24 ) );
  XOR2_X1 u1_u1_U34 (.B( u1_K2_23 ) , .A( u1_R0_16 ) , .Z( u1_u1_X_23 ) );
  XOR2_X1 u1_u1_U37 (.B( u1_K2_20 ) , .A( u1_R0_13 ) , .Z( u1_u1_X_20 ) );
  XOR2_X1 u1_u1_U39 (.B( u1_K2_19 ) , .A( u1_R0_12 ) , .Z( u1_u1_X_19 ) );
  XOR2_X1 u1_u1_U7 (.B( u1_K2_48 ) , .A( u1_R0_1 ) , .Z( u1_u1_X_48 ) );
  XOR2_X1 u1_u1_U8 (.B( u1_K2_47 ) , .A( u1_R0_32 ) , .Z( u1_u1_X_47 ) );
  OAI22_X1 u1_u1_u3_U10 (.B1( u1_u1_u3_n113 ) , .A2( u1_u1_u3_n135 ) , .A1( u1_u1_u3_n150 ) , .B2( u1_u1_u3_n164 ) , .ZN( u1_u1_u3_n98 ) );
  OAI211_X1 u1_u1_u3_U11 (.B( u1_u1_u3_n106 ) , .ZN( u1_u1_u3_n119 ) , .C2( u1_u1_u3_n128 ) , .C1( u1_u1_u3_n167 ) , .A( u1_u1_u3_n181 ) );
  AOI221_X1 u1_u1_u3_U12 (.C1( u1_u1_u3_n105 ) , .ZN( u1_u1_u3_n106 ) , .A( u1_u1_u3_n131 ) , .B2( u1_u1_u3_n132 ) , .C2( u1_u1_u3_n133 ) , .B1( u1_u1_u3_n169 ) );
  INV_X1 u1_u1_u3_U13 (.ZN( u1_u1_u3_n181 ) , .A( u1_u1_u3_n98 ) );
  NAND2_X1 u1_u1_u3_U14 (.ZN( u1_u1_u3_n105 ) , .A2( u1_u1_u3_n130 ) , .A1( u1_u1_u3_n155 ) );
  AOI22_X1 u1_u1_u3_U15 (.B1( u1_u1_u3_n115 ) , .A2( u1_u1_u3_n116 ) , .ZN( u1_u1_u3_n123 ) , .B2( u1_u1_u3_n133 ) , .A1( u1_u1_u3_n169 ) );
  NAND2_X1 u1_u1_u3_U16 (.ZN( u1_u1_u3_n116 ) , .A2( u1_u1_u3_n151 ) , .A1( u1_u1_u3_n182 ) );
  NOR2_X1 u1_u1_u3_U17 (.ZN( u1_u1_u3_n126 ) , .A2( u1_u1_u3_n150 ) , .A1( u1_u1_u3_n164 ) );
  AOI21_X1 u1_u1_u3_U18 (.ZN( u1_u1_u3_n112 ) , .B2( u1_u1_u3_n146 ) , .B1( u1_u1_u3_n155 ) , .A( u1_u1_u3_n167 ) );
  NAND2_X1 u1_u1_u3_U19 (.A1( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n142 ) , .A2( u1_u1_u3_n164 ) );
  NAND2_X1 u1_u1_u3_U20 (.ZN( u1_u1_u3_n132 ) , .A2( u1_u1_u3_n152 ) , .A1( u1_u1_u3_n156 ) );
  AND2_X1 u1_u1_u3_U21 (.A2( u1_u1_u3_n113 ) , .A1( u1_u1_u3_n114 ) , .ZN( u1_u1_u3_n151 ) );
  INV_X1 u1_u1_u3_U22 (.A( u1_u1_u3_n133 ) , .ZN( u1_u1_u3_n165 ) );
  INV_X1 u1_u1_u3_U23 (.A( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n170 ) );
  NAND2_X1 u1_u1_u3_U24 (.A1( u1_u1_u3_n107 ) , .A2( u1_u1_u3_n108 ) , .ZN( u1_u1_u3_n140 ) );
  NAND2_X1 u1_u1_u3_U25 (.ZN( u1_u1_u3_n117 ) , .A1( u1_u1_u3_n124 ) , .A2( u1_u1_u3_n148 ) );
  NAND2_X1 u1_u1_u3_U26 (.ZN( u1_u1_u3_n143 ) , .A1( u1_u1_u3_n165 ) , .A2( u1_u1_u3_n167 ) );
  INV_X1 u1_u1_u3_U27 (.A( u1_u1_u3_n130 ) , .ZN( u1_u1_u3_n177 ) );
  INV_X1 u1_u1_u3_U28 (.A( u1_u1_u3_n128 ) , .ZN( u1_u1_u3_n176 ) );
  INV_X1 u1_u1_u3_U29 (.A( u1_u1_u3_n155 ) , .ZN( u1_u1_u3_n174 ) );
  INV_X1 u1_u1_u3_U3 (.A( u1_u1_u3_n129 ) , .ZN( u1_u1_u3_n183 ) );
  INV_X1 u1_u1_u3_U30 (.A( u1_u1_u3_n139 ) , .ZN( u1_u1_u3_n185 ) );
  NOR2_X1 u1_u1_u3_U31 (.ZN( u1_u1_u3_n135 ) , .A2( u1_u1_u3_n141 ) , .A1( u1_u1_u3_n169 ) );
  OAI222_X1 u1_u1_u3_U32 (.C2( u1_u1_u3_n107 ) , .A2( u1_u1_u3_n108 ) , .B1( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n138 ) , .B2( u1_u1_u3_n146 ) , .C1( u1_u1_u3_n154 ) , .A1( u1_u1_u3_n164 ) );
  NOR4_X1 u1_u1_u3_U33 (.A4( u1_u1_u3_n157 ) , .A3( u1_u1_u3_n158 ) , .A2( u1_u1_u3_n159 ) , .A1( u1_u1_u3_n160 ) , .ZN( u1_u1_u3_n161 ) );
  AOI21_X1 u1_u1_u3_U34 (.B2( u1_u1_u3_n152 ) , .B1( u1_u1_u3_n153 ) , .ZN( u1_u1_u3_n158 ) , .A( u1_u1_u3_n164 ) );
  AOI21_X1 u1_u1_u3_U35 (.A( u1_u1_u3_n154 ) , .B2( u1_u1_u3_n155 ) , .B1( u1_u1_u3_n156 ) , .ZN( u1_u1_u3_n157 ) );
  AOI21_X1 u1_u1_u3_U36 (.A( u1_u1_u3_n149 ) , .B2( u1_u1_u3_n150 ) , .B1( u1_u1_u3_n151 ) , .ZN( u1_u1_u3_n159 ) );
  AOI211_X1 u1_u1_u3_U37 (.ZN( u1_u1_u3_n109 ) , .A( u1_u1_u3_n119 ) , .C2( u1_u1_u3_n129 ) , .B( u1_u1_u3_n138 ) , .C1( u1_u1_u3_n141 ) );
  AOI211_X1 u1_u1_u3_U38 (.B( u1_u1_u3_n119 ) , .A( u1_u1_u3_n120 ) , .C2( u1_u1_u3_n121 ) , .ZN( u1_u1_u3_n122 ) , .C1( u1_u1_u3_n179 ) );
  INV_X1 u1_u1_u3_U39 (.A( u1_u1_u3_n156 ) , .ZN( u1_u1_u3_n179 ) );
  INV_X1 u1_u1_u3_U4 (.A( u1_u1_u3_n140 ) , .ZN( u1_u1_u3_n182 ) );
  OAI22_X1 u1_u1_u3_U40 (.B1( u1_u1_u3_n118 ) , .ZN( u1_u1_u3_n120 ) , .A1( u1_u1_u3_n135 ) , .B2( u1_u1_u3_n154 ) , .A2( u1_u1_u3_n178 ) );
  AND3_X1 u1_u1_u3_U41 (.ZN( u1_u1_u3_n118 ) , .A2( u1_u1_u3_n124 ) , .A1( u1_u1_u3_n144 ) , .A3( u1_u1_u3_n152 ) );
  INV_X1 u1_u1_u3_U42 (.A( u1_u1_u3_n121 ) , .ZN( u1_u1_u3_n164 ) );
  NAND2_X1 u1_u1_u3_U43 (.ZN( u1_u1_u3_n133 ) , .A1( u1_u1_u3_n154 ) , .A2( u1_u1_u3_n164 ) );
  OAI211_X1 u1_u1_u3_U44 (.B( u1_u1_u3_n127 ) , .ZN( u1_u1_u3_n139 ) , .C1( u1_u1_u3_n150 ) , .C2( u1_u1_u3_n154 ) , .A( u1_u1_u3_n184 ) );
  INV_X1 u1_u1_u3_U45 (.A( u1_u1_u3_n125 ) , .ZN( u1_u1_u3_n184 ) );
  AOI221_X1 u1_u1_u3_U46 (.A( u1_u1_u3_n126 ) , .ZN( u1_u1_u3_n127 ) , .C2( u1_u1_u3_n132 ) , .C1( u1_u1_u3_n169 ) , .B2( u1_u1_u3_n170 ) , .B1( u1_u1_u3_n174 ) );
  OAI22_X1 u1_u1_u3_U47 (.A1( u1_u1_u3_n124 ) , .ZN( u1_u1_u3_n125 ) , .B2( u1_u1_u3_n145 ) , .A2( u1_u1_u3_n165 ) , .B1( u1_u1_u3_n167 ) );
  NOR2_X1 u1_u1_u3_U48 (.A1( u1_u1_u3_n113 ) , .ZN( u1_u1_u3_n131 ) , .A2( u1_u1_u3_n154 ) );
  NAND2_X1 u1_u1_u3_U49 (.A1( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n150 ) , .A2( u1_u1_u3_n99 ) );
  INV_X1 u1_u1_u3_U5 (.A( u1_u1_u3_n117 ) , .ZN( u1_u1_u3_n178 ) );
  NAND2_X1 u1_u1_u3_U50 (.A2( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n155 ) , .A1( u1_u1_u3_n97 ) );
  INV_X1 u1_u1_u3_U51 (.A( u1_u1_u3_n141 ) , .ZN( u1_u1_u3_n167 ) );
  AOI21_X1 u1_u1_u3_U52 (.B2( u1_u1_u3_n114 ) , .B1( u1_u1_u3_n146 ) , .A( u1_u1_u3_n154 ) , .ZN( u1_u1_u3_n94 ) );
  AOI21_X1 u1_u1_u3_U53 (.ZN( u1_u1_u3_n110 ) , .B2( u1_u1_u3_n142 ) , .B1( u1_u1_u3_n186 ) , .A( u1_u1_u3_n95 ) );
  INV_X1 u1_u1_u3_U54 (.A( u1_u1_u3_n145 ) , .ZN( u1_u1_u3_n186 ) );
  AOI21_X1 u1_u1_u3_U55 (.B1( u1_u1_u3_n124 ) , .A( u1_u1_u3_n149 ) , .B2( u1_u1_u3_n155 ) , .ZN( u1_u1_u3_n95 ) );
  INV_X1 u1_u1_u3_U56 (.A( u1_u1_u3_n149 ) , .ZN( u1_u1_u3_n169 ) );
  NAND2_X1 u1_u1_u3_U57 (.ZN( u1_u1_u3_n124 ) , .A1( u1_u1_u3_n96 ) , .A2( u1_u1_u3_n97 ) );
  NAND2_X1 u1_u1_u3_U58 (.A2( u1_u1_u3_n100 ) , .ZN( u1_u1_u3_n146 ) , .A1( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U59 (.A1( u1_u1_u3_n101 ) , .ZN( u1_u1_u3_n145 ) , .A2( u1_u1_u3_n99 ) );
  AOI221_X1 u1_u1_u3_U6 (.A( u1_u1_u3_n131 ) , .C2( u1_u1_u3_n132 ) , .C1( u1_u1_u3_n133 ) , .ZN( u1_u1_u3_n134 ) , .B1( u1_u1_u3_n143 ) , .B2( u1_u1_u3_n177 ) );
  NAND2_X1 u1_u1_u3_U60 (.A1( u1_u1_u3_n100 ) , .ZN( u1_u1_u3_n156 ) , .A2( u1_u1_u3_n99 ) );
  NAND2_X1 u1_u1_u3_U61 (.A2( u1_u1_u3_n101 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n148 ) );
  NAND2_X1 u1_u1_u3_U62 (.A1( u1_u1_u3_n100 ) , .A2( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n128 ) );
  NAND2_X1 u1_u1_u3_U63 (.A2( u1_u1_u3_n101 ) , .A1( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n152 ) );
  NAND2_X1 u1_u1_u3_U64 (.A2( u1_u1_u3_n101 ) , .ZN( u1_u1_u3_n114 ) , .A1( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U65 (.ZN( u1_u1_u3_n107 ) , .A1( u1_u1_u3_n97 ) , .A2( u1_u1_u3_n99 ) );
  NAND2_X1 u1_u1_u3_U66 (.A2( u1_u1_u3_n100 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n113 ) );
  NAND2_X1 u1_u1_u3_U67 (.A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n153 ) , .A2( u1_u1_u3_n97 ) );
  NAND2_X1 u1_u1_u3_U68 (.A2( u1_u1_u3_n103 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n130 ) );
  NAND2_X1 u1_u1_u3_U69 (.A2( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n144 ) , .A1( u1_u1_u3_n96 ) );
  OAI22_X1 u1_u1_u3_U7 (.B2( u1_u1_u3_n147 ) , .A2( u1_u1_u3_n148 ) , .ZN( u1_u1_u3_n160 ) , .B1( u1_u1_u3_n165 ) , .A1( u1_u1_u3_n168 ) );
  NAND2_X1 u1_u1_u3_U70 (.A1( u1_u1_u3_n102 ) , .A2( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n108 ) );
  NOR2_X1 u1_u1_u3_U71 (.A2( u1_u1_X_19 ) , .A1( u1_u1_X_20 ) , .ZN( u1_u1_u3_n99 ) );
  NOR2_X1 u1_u1_u3_U72 (.A2( u1_u1_X_21 ) , .A1( u1_u1_X_24 ) , .ZN( u1_u1_u3_n103 ) );
  NOR2_X1 u1_u1_u3_U73 (.A2( u1_u1_X_24 ) , .A1( u1_u1_u3_n171 ) , .ZN( u1_u1_u3_n97 ) );
  NOR2_X1 u1_u1_u3_U74 (.A2( u1_u1_X_23 ) , .ZN( u1_u1_u3_n141 ) , .A1( u1_u1_u3_n166 ) );
  NOR2_X1 u1_u1_u3_U75 (.A2( u1_u1_X_19 ) , .A1( u1_u1_u3_n172 ) , .ZN( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U76 (.A1( u1_u1_X_22 ) , .A2( u1_u1_X_23 ) , .ZN( u1_u1_u3_n154 ) );
  NAND2_X1 u1_u1_u3_U77 (.A1( u1_u1_X_23 ) , .ZN( u1_u1_u3_n149 ) , .A2( u1_u1_u3_n166 ) );
  NOR2_X1 u1_u1_u3_U78 (.A2( u1_u1_X_22 ) , .A1( u1_u1_X_23 ) , .ZN( u1_u1_u3_n121 ) );
  AND2_X1 u1_u1_u3_U79 (.A1( u1_u1_X_24 ) , .ZN( u1_u1_u3_n101 ) , .A2( u1_u1_u3_n171 ) );
  AND3_X1 u1_u1_u3_U8 (.A3( u1_u1_u3_n144 ) , .A2( u1_u1_u3_n145 ) , .A1( u1_u1_u3_n146 ) , .ZN( u1_u1_u3_n147 ) );
  AND2_X1 u1_u1_u3_U80 (.A1( u1_u1_X_19 ) , .ZN( u1_u1_u3_n102 ) , .A2( u1_u1_u3_n172 ) );
  AND2_X1 u1_u1_u3_U81 (.A1( u1_u1_X_21 ) , .A2( u1_u1_X_24 ) , .ZN( u1_u1_u3_n100 ) );
  AND2_X1 u1_u1_u3_U82 (.A2( u1_u1_X_19 ) , .A1( u1_u1_X_20 ) , .ZN( u1_u1_u3_n104 ) );
  INV_X1 u1_u1_u3_U83 (.A( u1_u1_X_22 ) , .ZN( u1_u1_u3_n166 ) );
  INV_X1 u1_u1_u3_U84 (.A( u1_u1_X_21 ) , .ZN( u1_u1_u3_n171 ) );
  INV_X1 u1_u1_u3_U85 (.A( u1_u1_X_20 ) , .ZN( u1_u1_u3_n172 ) );
  OR4_X1 u1_u1_u3_U86 (.ZN( u1_out1_10 ) , .A4( u1_u1_u3_n136 ) , .A3( u1_u1_u3_n137 ) , .A1( u1_u1_u3_n138 ) , .A2( u1_u1_u3_n139 ) );
  OAI222_X1 u1_u1_u3_U87 (.C1( u1_u1_u3_n128 ) , .ZN( u1_u1_u3_n137 ) , .B1( u1_u1_u3_n148 ) , .A2( u1_u1_u3_n150 ) , .B2( u1_u1_u3_n154 ) , .C2( u1_u1_u3_n164 ) , .A1( u1_u1_u3_n167 ) );
  OAI221_X1 u1_u1_u3_U88 (.A( u1_u1_u3_n134 ) , .B2( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n136 ) , .C1( u1_u1_u3_n149 ) , .B1( u1_u1_u3_n151 ) , .C2( u1_u1_u3_n183 ) );
  NAND4_X1 u1_u1_u3_U89 (.ZN( u1_out1_26 ) , .A4( u1_u1_u3_n109 ) , .A3( u1_u1_u3_n110 ) , .A2( u1_u1_u3_n111 ) , .A1( u1_u1_u3_n173 ) );
  INV_X1 u1_u1_u3_U9 (.A( u1_u1_u3_n143 ) , .ZN( u1_u1_u3_n168 ) );
  INV_X1 u1_u1_u3_U90 (.ZN( u1_u1_u3_n173 ) , .A( u1_u1_u3_n94 ) );
  OAI21_X1 u1_u1_u3_U91 (.ZN( u1_u1_u3_n111 ) , .B2( u1_u1_u3_n117 ) , .A( u1_u1_u3_n133 ) , .B1( u1_u1_u3_n176 ) );
  NAND4_X1 u1_u1_u3_U92 (.ZN( u1_out1_20 ) , .A4( u1_u1_u3_n122 ) , .A3( u1_u1_u3_n123 ) , .A1( u1_u1_u3_n175 ) , .A2( u1_u1_u3_n180 ) );
  INV_X1 u1_u1_u3_U93 (.A( u1_u1_u3_n112 ) , .ZN( u1_u1_u3_n175 ) );
  INV_X1 u1_u1_u3_U94 (.A( u1_u1_u3_n126 ) , .ZN( u1_u1_u3_n180 ) );
  NAND4_X1 u1_u1_u3_U95 (.ZN( u1_out1_1 ) , .A4( u1_u1_u3_n161 ) , .A3( u1_u1_u3_n162 ) , .A2( u1_u1_u3_n163 ) , .A1( u1_u1_u3_n185 ) );
  NAND2_X1 u1_u1_u3_U96 (.ZN( u1_u1_u3_n163 ) , .A2( u1_u1_u3_n170 ) , .A1( u1_u1_u3_n176 ) );
  AOI22_X1 u1_u1_u3_U97 (.B2( u1_u1_u3_n140 ) , .B1( u1_u1_u3_n141 ) , .A2( u1_u1_u3_n142 ) , .ZN( u1_u1_u3_n162 ) , .A1( u1_u1_u3_n177 ) );
  NAND3_X1 u1_u1_u3_U98 (.A1( u1_u1_u3_n114 ) , .ZN( u1_u1_u3_n115 ) , .A2( u1_u1_u3_n145 ) , .A3( u1_u1_u3_n153 ) );
  NAND3_X1 u1_u1_u3_U99 (.ZN( u1_u1_u3_n129 ) , .A2( u1_u1_u3_n144 ) , .A1( u1_u1_u3_n153 ) , .A3( u1_u1_u3_n182 ) );
  OAI22_X1 u1_u1_u4_U10 (.B2( u1_u1_u4_n135 ) , .ZN( u1_u1_u4_n137 ) , .B1( u1_u1_u4_n153 ) , .A1( u1_u1_u4_n155 ) , .A2( u1_u1_u4_n171 ) );
  AND3_X1 u1_u1_u4_U11 (.A2( u1_u1_u4_n134 ) , .ZN( u1_u1_u4_n135 ) , .A3( u1_u1_u4_n145 ) , .A1( u1_u1_u4_n157 ) );
  NAND2_X1 u1_u1_u4_U12 (.ZN( u1_u1_u4_n132 ) , .A2( u1_u1_u4_n170 ) , .A1( u1_u1_u4_n173 ) );
  AOI21_X1 u1_u1_u4_U13 (.B2( u1_u1_u4_n160 ) , .B1( u1_u1_u4_n161 ) , .ZN( u1_u1_u4_n162 ) , .A( u1_u1_u4_n170 ) );
  AOI21_X1 u1_u1_u4_U14 (.ZN( u1_u1_u4_n107 ) , .B2( u1_u1_u4_n143 ) , .A( u1_u1_u4_n174 ) , .B1( u1_u1_u4_n184 ) );
  AOI21_X1 u1_u1_u4_U15 (.B2( u1_u1_u4_n158 ) , .B1( u1_u1_u4_n159 ) , .ZN( u1_u1_u4_n163 ) , .A( u1_u1_u4_n174 ) );
  AOI21_X1 u1_u1_u4_U16 (.A( u1_u1_u4_n153 ) , .B2( u1_u1_u4_n154 ) , .B1( u1_u1_u4_n155 ) , .ZN( u1_u1_u4_n165 ) );
  AOI21_X1 u1_u1_u4_U17 (.A( u1_u1_u4_n156 ) , .B2( u1_u1_u4_n157 ) , .ZN( u1_u1_u4_n164 ) , .B1( u1_u1_u4_n184 ) );
  INV_X1 u1_u1_u4_U18 (.A( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n170 ) );
  AND2_X1 u1_u1_u4_U19 (.A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n155 ) , .A1( u1_u1_u4_n160 ) );
  INV_X1 u1_u1_u4_U20 (.A( u1_u1_u4_n156 ) , .ZN( u1_u1_u4_n175 ) );
  NAND2_X1 u1_u1_u4_U21 (.A2( u1_u1_u4_n118 ) , .ZN( u1_u1_u4_n131 ) , .A1( u1_u1_u4_n147 ) );
  NAND2_X1 u1_u1_u4_U22 (.A1( u1_u1_u4_n119 ) , .A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n130 ) );
  NAND2_X1 u1_u1_u4_U23 (.ZN( u1_u1_u4_n117 ) , .A2( u1_u1_u4_n118 ) , .A1( u1_u1_u4_n148 ) );
  NAND2_X1 u1_u1_u4_U24 (.ZN( u1_u1_u4_n129 ) , .A1( u1_u1_u4_n134 ) , .A2( u1_u1_u4_n148 ) );
  AND3_X1 u1_u1_u4_U25 (.A1( u1_u1_u4_n119 ) , .A2( u1_u1_u4_n143 ) , .A3( u1_u1_u4_n154 ) , .ZN( u1_u1_u4_n161 ) );
  AND2_X1 u1_u1_u4_U26 (.A1( u1_u1_u4_n145 ) , .A2( u1_u1_u4_n147 ) , .ZN( u1_u1_u4_n159 ) );
  OR3_X1 u1_u1_u4_U27 (.A3( u1_u1_u4_n114 ) , .A2( u1_u1_u4_n115 ) , .A1( u1_u1_u4_n116 ) , .ZN( u1_u1_u4_n136 ) );
  AOI21_X1 u1_u1_u4_U28 (.A( u1_u1_u4_n113 ) , .ZN( u1_u1_u4_n116 ) , .B2( u1_u1_u4_n173 ) , .B1( u1_u1_u4_n174 ) );
  AOI21_X1 u1_u1_u4_U29 (.ZN( u1_u1_u4_n115 ) , .B2( u1_u1_u4_n145 ) , .B1( u1_u1_u4_n146 ) , .A( u1_u1_u4_n156 ) );
  NOR2_X1 u1_u1_u4_U3 (.ZN( u1_u1_u4_n121 ) , .A1( u1_u1_u4_n181 ) , .A2( u1_u1_u4_n182 ) );
  OAI22_X1 u1_u1_u4_U30 (.ZN( u1_u1_u4_n114 ) , .A2( u1_u1_u4_n121 ) , .B1( u1_u1_u4_n160 ) , .B2( u1_u1_u4_n170 ) , .A1( u1_u1_u4_n171 ) );
  INV_X1 u1_u1_u4_U31 (.A( u1_u1_u4_n158 ) , .ZN( u1_u1_u4_n182 ) );
  INV_X1 u1_u1_u4_U32 (.ZN( u1_u1_u4_n181 ) , .A( u1_u1_u4_n96 ) );
  INV_X1 u1_u1_u4_U33 (.A( u1_u1_u4_n144 ) , .ZN( u1_u1_u4_n179 ) );
  INV_X1 u1_u1_u4_U34 (.A( u1_u1_u4_n157 ) , .ZN( u1_u1_u4_n178 ) );
  NAND2_X1 u1_u1_u4_U35 (.A2( u1_u1_u4_n154 ) , .A1( u1_u1_u4_n96 ) , .ZN( u1_u1_u4_n97 ) );
  INV_X1 u1_u1_u4_U36 (.ZN( u1_u1_u4_n186 ) , .A( u1_u1_u4_n95 ) );
  OAI221_X1 u1_u1_u4_U37 (.C1( u1_u1_u4_n134 ) , .B1( u1_u1_u4_n158 ) , .B2( u1_u1_u4_n171 ) , .C2( u1_u1_u4_n173 ) , .A( u1_u1_u4_n94 ) , .ZN( u1_u1_u4_n95 ) );
  AOI222_X1 u1_u1_u4_U38 (.B2( u1_u1_u4_n132 ) , .A1( u1_u1_u4_n138 ) , .C2( u1_u1_u4_n175 ) , .A2( u1_u1_u4_n179 ) , .C1( u1_u1_u4_n181 ) , .B1( u1_u1_u4_n185 ) , .ZN( u1_u1_u4_n94 ) );
  INV_X1 u1_u1_u4_U39 (.A( u1_u1_u4_n113 ) , .ZN( u1_u1_u4_n185 ) );
  INV_X1 u1_u1_u4_U4 (.A( u1_u1_u4_n117 ) , .ZN( u1_u1_u4_n184 ) );
  INV_X1 u1_u1_u4_U40 (.A( u1_u1_u4_n143 ) , .ZN( u1_u1_u4_n183 ) );
  NOR2_X1 u1_u1_u4_U41 (.ZN( u1_u1_u4_n138 ) , .A1( u1_u1_u4_n168 ) , .A2( u1_u1_u4_n169 ) );
  NOR2_X1 u1_u1_u4_U42 (.A1( u1_u1_u4_n150 ) , .A2( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n153 ) );
  NOR2_X1 u1_u1_u4_U43 (.A2( u1_u1_u4_n128 ) , .A1( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n156 ) );
  AOI22_X1 u1_u1_u4_U44 (.B2( u1_u1_u4_n122 ) , .A1( u1_u1_u4_n123 ) , .ZN( u1_u1_u4_n124 ) , .B1( u1_u1_u4_n128 ) , .A2( u1_u1_u4_n172 ) );
  NAND2_X1 u1_u1_u4_U45 (.A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n123 ) , .A1( u1_u1_u4_n161 ) );
  INV_X1 u1_u1_u4_U46 (.A( u1_u1_u4_n153 ) , .ZN( u1_u1_u4_n172 ) );
  AOI22_X1 u1_u1_u4_U47 (.B2( u1_u1_u4_n132 ) , .A2( u1_u1_u4_n133 ) , .ZN( u1_u1_u4_n140 ) , .A1( u1_u1_u4_n150 ) , .B1( u1_u1_u4_n179 ) );
  NAND2_X1 u1_u1_u4_U48 (.ZN( u1_u1_u4_n133 ) , .A2( u1_u1_u4_n146 ) , .A1( u1_u1_u4_n154 ) );
  NAND2_X1 u1_u1_u4_U49 (.A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n154 ) , .A2( u1_u1_u4_n98 ) );
  NOR4_X1 u1_u1_u4_U5 (.A4( u1_u1_u4_n106 ) , .A3( u1_u1_u4_n107 ) , .A2( u1_u1_u4_n108 ) , .A1( u1_u1_u4_n109 ) , .ZN( u1_u1_u4_n110 ) );
  NAND2_X1 u1_u1_u4_U50 (.A1( u1_u1_u4_n101 ) , .ZN( u1_u1_u4_n158 ) , .A2( u1_u1_u4_n99 ) );
  AOI21_X1 u1_u1_u4_U51 (.ZN( u1_u1_u4_n127 ) , .A( u1_u1_u4_n136 ) , .B2( u1_u1_u4_n150 ) , .B1( u1_u1_u4_n180 ) );
  INV_X1 u1_u1_u4_U52 (.A( u1_u1_u4_n160 ) , .ZN( u1_u1_u4_n180 ) );
  NAND2_X1 u1_u1_u4_U53 (.A2( u1_u1_u4_n104 ) , .A1( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n146 ) );
  NAND2_X1 u1_u1_u4_U54 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n160 ) );
  NAND2_X1 u1_u1_u4_U55 (.ZN( u1_u1_u4_n134 ) , .A1( u1_u1_u4_n98 ) , .A2( u1_u1_u4_n99 ) );
  NAND2_X1 u1_u1_u4_U56 (.A1( u1_u1_u4_n103 ) , .A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n143 ) );
  NAND2_X1 u1_u1_u4_U57 (.A2( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n145 ) , .A1( u1_u1_u4_n98 ) );
  NAND2_X1 u1_u1_u4_U58 (.A1( u1_u1_u4_n100 ) , .A2( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n120 ) );
  NAND2_X1 u1_u1_u4_U59 (.A1( u1_u1_u4_n102 ) , .A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n148 ) );
  AOI21_X1 u1_u1_u4_U6 (.ZN( u1_u1_u4_n106 ) , .B2( u1_u1_u4_n146 ) , .B1( u1_u1_u4_n158 ) , .A( u1_u1_u4_n170 ) );
  NAND2_X1 u1_u1_u4_U60 (.A2( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n157 ) );
  INV_X1 u1_u1_u4_U61 (.A( u1_u1_u4_n150 ) , .ZN( u1_u1_u4_n173 ) );
  INV_X1 u1_u1_u4_U62 (.A( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n171 ) );
  NAND2_X1 u1_u1_u4_U63 (.A1( u1_u1_u4_n100 ) , .ZN( u1_u1_u4_n118 ) , .A2( u1_u1_u4_n99 ) );
  NAND2_X1 u1_u1_u4_U64 (.A2( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n144 ) );
  NAND2_X1 u1_u1_u4_U65 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n96 ) );
  INV_X1 u1_u1_u4_U66 (.A( u1_u1_u4_n128 ) , .ZN( u1_u1_u4_n174 ) );
  NAND2_X1 u1_u1_u4_U67 (.A2( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n119 ) , .A1( u1_u1_u4_n98 ) );
  NAND2_X1 u1_u1_u4_U68 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n147 ) );
  NAND2_X1 u1_u1_u4_U69 (.A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n113 ) , .A1( u1_u1_u4_n99 ) );
  AOI21_X1 u1_u1_u4_U7 (.ZN( u1_u1_u4_n108 ) , .B2( u1_u1_u4_n134 ) , .B1( u1_u1_u4_n155 ) , .A( u1_u1_u4_n156 ) );
  NOR2_X1 u1_u1_u4_U70 (.A2( u1_u1_X_28 ) , .ZN( u1_u1_u4_n150 ) , .A1( u1_u1_u4_n168 ) );
  NOR2_X1 u1_u1_u4_U71 (.A2( u1_u1_X_29 ) , .ZN( u1_u1_u4_n152 ) , .A1( u1_u1_u4_n169 ) );
  NOR2_X1 u1_u1_u4_U72 (.A2( u1_u1_X_30 ) , .ZN( u1_u1_u4_n105 ) , .A1( u1_u1_u4_n176 ) );
  NOR2_X1 u1_u1_u4_U73 (.A2( u1_u1_X_26 ) , .ZN( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n177 ) );
  NOR2_X1 u1_u1_u4_U74 (.A2( u1_u1_X_28 ) , .A1( u1_u1_X_29 ) , .ZN( u1_u1_u4_n128 ) );
  NOR2_X1 u1_u1_u4_U75 (.A2( u1_u1_X_27 ) , .A1( u1_u1_X_30 ) , .ZN( u1_u1_u4_n102 ) );
  NOR2_X1 u1_u1_u4_U76 (.A2( u1_u1_X_25 ) , .A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n98 ) );
  AND2_X1 u1_u1_u4_U77 (.A2( u1_u1_X_25 ) , .A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n104 ) );
  AND2_X1 u1_u1_u4_U78 (.A1( u1_u1_X_30 ) , .A2( u1_u1_u4_n176 ) , .ZN( u1_u1_u4_n99 ) );
  AND2_X1 u1_u1_u4_U79 (.A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n101 ) , .A2( u1_u1_u4_n177 ) );
  AOI21_X1 u1_u1_u4_U8 (.ZN( u1_u1_u4_n109 ) , .A( u1_u1_u4_n153 ) , .B1( u1_u1_u4_n159 ) , .B2( u1_u1_u4_n184 ) );
  AND2_X1 u1_u1_u4_U80 (.A1( u1_u1_X_27 ) , .A2( u1_u1_X_30 ) , .ZN( u1_u1_u4_n103 ) );
  INV_X1 u1_u1_u4_U81 (.A( u1_u1_X_28 ) , .ZN( u1_u1_u4_n169 ) );
  INV_X1 u1_u1_u4_U82 (.A( u1_u1_X_29 ) , .ZN( u1_u1_u4_n168 ) );
  INV_X1 u1_u1_u4_U83 (.A( u1_u1_X_25 ) , .ZN( u1_u1_u4_n177 ) );
  INV_X1 u1_u1_u4_U84 (.A( u1_u1_X_27 ) , .ZN( u1_u1_u4_n176 ) );
  NAND4_X1 u1_u1_u4_U85 (.ZN( u1_out1_25 ) , .A4( u1_u1_u4_n139 ) , .A3( u1_u1_u4_n140 ) , .A2( u1_u1_u4_n141 ) , .A1( u1_u1_u4_n142 ) );
  OAI21_X1 u1_u1_u4_U86 (.A( u1_u1_u4_n128 ) , .B2( u1_u1_u4_n129 ) , .B1( u1_u1_u4_n130 ) , .ZN( u1_u1_u4_n142 ) );
  OAI21_X1 u1_u1_u4_U87 (.B2( u1_u1_u4_n131 ) , .ZN( u1_u1_u4_n141 ) , .A( u1_u1_u4_n175 ) , .B1( u1_u1_u4_n183 ) );
  NAND4_X1 u1_u1_u4_U88 (.ZN( u1_out1_14 ) , .A4( u1_u1_u4_n124 ) , .A3( u1_u1_u4_n125 ) , .A2( u1_u1_u4_n126 ) , .A1( u1_u1_u4_n127 ) );
  AOI22_X1 u1_u1_u4_U89 (.B2( u1_u1_u4_n117 ) , .ZN( u1_u1_u4_n126 ) , .A1( u1_u1_u4_n129 ) , .B1( u1_u1_u4_n152 ) , .A2( u1_u1_u4_n175 ) );
  AOI211_X1 u1_u1_u4_U9 (.B( u1_u1_u4_n136 ) , .A( u1_u1_u4_n137 ) , .C2( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n139 ) , .C1( u1_u1_u4_n182 ) );
  AOI22_X1 u1_u1_u4_U90 (.ZN( u1_u1_u4_n125 ) , .B2( u1_u1_u4_n131 ) , .A2( u1_u1_u4_n132 ) , .B1( u1_u1_u4_n138 ) , .A1( u1_u1_u4_n178 ) );
  NAND4_X1 u1_u1_u4_U91 (.ZN( u1_out1_8 ) , .A4( u1_u1_u4_n110 ) , .A3( u1_u1_u4_n111 ) , .A2( u1_u1_u4_n112 ) , .A1( u1_u1_u4_n186 ) );
  NAND2_X1 u1_u1_u4_U92 (.ZN( u1_u1_u4_n112 ) , .A2( u1_u1_u4_n130 ) , .A1( u1_u1_u4_n150 ) );
  AOI22_X1 u1_u1_u4_U93 (.ZN( u1_u1_u4_n111 ) , .B2( u1_u1_u4_n132 ) , .A1( u1_u1_u4_n152 ) , .B1( u1_u1_u4_n178 ) , .A2( u1_u1_u4_n97 ) );
  AOI22_X1 u1_u1_u4_U94 (.B2( u1_u1_u4_n149 ) , .B1( u1_u1_u4_n150 ) , .A2( u1_u1_u4_n151 ) , .A1( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n167 ) );
  NOR4_X1 u1_u1_u4_U95 (.A4( u1_u1_u4_n162 ) , .A3( u1_u1_u4_n163 ) , .A2( u1_u1_u4_n164 ) , .A1( u1_u1_u4_n165 ) , .ZN( u1_u1_u4_n166 ) );
  NAND3_X1 u1_u1_u4_U96 (.ZN( u1_out1_3 ) , .A3( u1_u1_u4_n166 ) , .A1( u1_u1_u4_n167 ) , .A2( u1_u1_u4_n186 ) );
  NAND3_X1 u1_u1_u4_U97 (.A3( u1_u1_u4_n146 ) , .A2( u1_u1_u4_n147 ) , .A1( u1_u1_u4_n148 ) , .ZN( u1_u1_u4_n149 ) );
  NAND3_X1 u1_u1_u4_U98 (.A3( u1_u1_u4_n143 ) , .A2( u1_u1_u4_n144 ) , .A1( u1_u1_u4_n145 ) , .ZN( u1_u1_u4_n151 ) );
  NAND3_X1 u1_u1_u4_U99 (.A3( u1_u1_u4_n121 ) , .ZN( u1_u1_u4_n122 ) , .A2( u1_u1_u4_n144 ) , .A1( u1_u1_u4_n154 ) );
  AOI22_X1 u1_u1_u6_U10 (.A2( u1_u1_u6_n151 ) , .B2( u1_u1_u6_n161 ) , .A1( u1_u1_u6_n167 ) , .B1( u1_u1_u6_n170 ) , .ZN( u1_u1_u6_n89 ) );
  AOI21_X1 u1_u1_u6_U11 (.B1( u1_u1_u6_n107 ) , .B2( u1_u1_u6_n132 ) , .A( u1_u1_u6_n158 ) , .ZN( u1_u1_u6_n88 ) );
  AOI21_X1 u1_u1_u6_U12 (.B2( u1_u1_u6_n147 ) , .B1( u1_u1_u6_n148 ) , .ZN( u1_u1_u6_n149 ) , .A( u1_u1_u6_n158 ) );
  AOI21_X1 u1_u1_u6_U13 (.ZN( u1_u1_u6_n106 ) , .A( u1_u1_u6_n142 ) , .B2( u1_u1_u6_n159 ) , .B1( u1_u1_u6_n164 ) );
  INV_X1 u1_u1_u6_U14 (.A( u1_u1_u6_n155 ) , .ZN( u1_u1_u6_n161 ) );
  INV_X1 u1_u1_u6_U15 (.A( u1_u1_u6_n128 ) , .ZN( u1_u1_u6_n164 ) );
  NAND2_X1 u1_u1_u6_U16 (.ZN( u1_u1_u6_n110 ) , .A1( u1_u1_u6_n122 ) , .A2( u1_u1_u6_n129 ) );
  NAND2_X1 u1_u1_u6_U17 (.ZN( u1_u1_u6_n124 ) , .A2( u1_u1_u6_n146 ) , .A1( u1_u1_u6_n148 ) );
  INV_X1 u1_u1_u6_U18 (.A( u1_u1_u6_n132 ) , .ZN( u1_u1_u6_n171 ) );
  AND2_X1 u1_u1_u6_U19 (.A1( u1_u1_u6_n100 ) , .ZN( u1_u1_u6_n130 ) , .A2( u1_u1_u6_n147 ) );
  INV_X1 u1_u1_u6_U20 (.A( u1_u1_u6_n127 ) , .ZN( u1_u1_u6_n173 ) );
  INV_X1 u1_u1_u6_U21 (.A( u1_u1_u6_n121 ) , .ZN( u1_u1_u6_n167 ) );
  INV_X1 u1_u1_u6_U22 (.A( u1_u1_u6_n100 ) , .ZN( u1_u1_u6_n169 ) );
  INV_X1 u1_u1_u6_U23 (.A( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n170 ) );
  INV_X1 u1_u1_u6_U24 (.A( u1_u1_u6_n113 ) , .ZN( u1_u1_u6_n168 ) );
  AND2_X1 u1_u1_u6_U25 (.A1( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n119 ) , .ZN( u1_u1_u6_n133 ) );
  AND2_X1 u1_u1_u6_U26 (.A2( u1_u1_u6_n121 ) , .A1( u1_u1_u6_n122 ) , .ZN( u1_u1_u6_n131 ) );
  AND3_X1 u1_u1_u6_U27 (.ZN( u1_u1_u6_n120 ) , .A2( u1_u1_u6_n127 ) , .A1( u1_u1_u6_n132 ) , .A3( u1_u1_u6_n145 ) );
  INV_X1 u1_u1_u6_U28 (.A( u1_u1_u6_n146 ) , .ZN( u1_u1_u6_n163 ) );
  AOI222_X1 u1_u1_u6_U29 (.ZN( u1_u1_u6_n114 ) , .A1( u1_u1_u6_n118 ) , .A2( u1_u1_u6_n126 ) , .B2( u1_u1_u6_n151 ) , .C2( u1_u1_u6_n159 ) , .C1( u1_u1_u6_n168 ) , .B1( u1_u1_u6_n169 ) );
  INV_X1 u1_u1_u6_U3 (.A( u1_u1_u6_n110 ) , .ZN( u1_u1_u6_n166 ) );
  NOR2_X1 u1_u1_u6_U30 (.A1( u1_u1_u6_n162 ) , .A2( u1_u1_u6_n165 ) , .ZN( u1_u1_u6_n98 ) );
  AOI211_X1 u1_u1_u6_U31 (.B( u1_u1_u6_n134 ) , .A( u1_u1_u6_n135 ) , .C1( u1_u1_u6_n136 ) , .ZN( u1_u1_u6_n137 ) , .C2( u1_u1_u6_n151 ) );
  AOI21_X1 u1_u1_u6_U32 (.B1( u1_u1_u6_n131 ) , .ZN( u1_u1_u6_n135 ) , .A( u1_u1_u6_n144 ) , .B2( u1_u1_u6_n146 ) );
  NAND4_X1 u1_u1_u6_U33 (.A4( u1_u1_u6_n127 ) , .A3( u1_u1_u6_n128 ) , .A2( u1_u1_u6_n129 ) , .A1( u1_u1_u6_n130 ) , .ZN( u1_u1_u6_n136 ) );
  AOI21_X1 u1_u1_u6_U34 (.B2( u1_u1_u6_n132 ) , .B1( u1_u1_u6_n133 ) , .ZN( u1_u1_u6_n134 ) , .A( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U35 (.A1( u1_u1_u6_n144 ) , .ZN( u1_u1_u6_n151 ) , .A2( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U36 (.ZN( u1_u1_u6_n132 ) , .A1( u1_u1_u6_n91 ) , .A2( u1_u1_u6_n97 ) );
  AOI22_X1 u1_u1_u6_U37 (.B2( u1_u1_u6_n110 ) , .B1( u1_u1_u6_n111 ) , .A1( u1_u1_u6_n112 ) , .ZN( u1_u1_u6_n115 ) , .A2( u1_u1_u6_n161 ) );
  NAND4_X1 u1_u1_u6_U38 (.A3( u1_u1_u6_n109 ) , .ZN( u1_u1_u6_n112 ) , .A4( u1_u1_u6_n132 ) , .A2( u1_u1_u6_n147 ) , .A1( u1_u1_u6_n166 ) );
  NOR2_X1 u1_u1_u6_U39 (.ZN( u1_u1_u6_n109 ) , .A1( u1_u1_u6_n170 ) , .A2( u1_u1_u6_n173 ) );
  INV_X1 u1_u1_u6_U4 (.A( u1_u1_u6_n142 ) , .ZN( u1_u1_u6_n174 ) );
  NOR2_X1 u1_u1_u6_U40 (.A2( u1_u1_u6_n126 ) , .ZN( u1_u1_u6_n155 ) , .A1( u1_u1_u6_n160 ) );
  NAND2_X1 u1_u1_u6_U41 (.ZN( u1_u1_u6_n146 ) , .A2( u1_u1_u6_n94 ) , .A1( u1_u1_u6_n99 ) );
  AOI21_X1 u1_u1_u6_U42 (.A( u1_u1_u6_n144 ) , .B2( u1_u1_u6_n145 ) , .B1( u1_u1_u6_n146 ) , .ZN( u1_u1_u6_n150 ) );
  INV_X1 u1_u1_u6_U43 (.A( u1_u1_u6_n111 ) , .ZN( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U44 (.ZN( u1_u1_u6_n127 ) , .A1( u1_u1_u6_n91 ) , .A2( u1_u1_u6_n92 ) );
  NAND2_X1 u1_u1_u6_U45 (.ZN( u1_u1_u6_n129 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n96 ) );
  INV_X1 u1_u1_u6_U46 (.A( u1_u1_u6_n144 ) , .ZN( u1_u1_u6_n159 ) );
  NAND2_X1 u1_u1_u6_U47 (.ZN( u1_u1_u6_n145 ) , .A2( u1_u1_u6_n97 ) , .A1( u1_u1_u6_n98 ) );
  NAND2_X1 u1_u1_u6_U48 (.ZN( u1_u1_u6_n148 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n94 ) );
  NAND2_X1 u1_u1_u6_U49 (.ZN( u1_u1_u6_n108 ) , .A2( u1_u1_u6_n139 ) , .A1( u1_u1_u6_n144 ) );
  NAND2_X1 u1_u1_u6_U5 (.A2( u1_u1_u6_n143 ) , .ZN( u1_u1_u6_n152 ) , .A1( u1_u1_u6_n166 ) );
  NAND2_X1 u1_u1_u6_U50 (.ZN( u1_u1_u6_n121 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n97 ) );
  NAND2_X1 u1_u1_u6_U51 (.ZN( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n95 ) );
  AND2_X1 u1_u1_u6_U52 (.ZN( u1_u1_u6_n118 ) , .A2( u1_u1_u6_n91 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U53 (.ZN( u1_u1_u6_n147 ) , .A2( u1_u1_u6_n98 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U54 (.ZN( u1_u1_u6_n128 ) , .A1( u1_u1_u6_n94 ) , .A2( u1_u1_u6_n96 ) );
  NAND2_X1 u1_u1_u6_U55 (.ZN( u1_u1_u6_n119 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U56 (.ZN( u1_u1_u6_n123 ) , .A2( u1_u1_u6_n91 ) , .A1( u1_u1_u6_n96 ) );
  NAND2_X1 u1_u1_u6_U57 (.ZN( u1_u1_u6_n100 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n98 ) );
  NAND2_X1 u1_u1_u6_U58 (.ZN( u1_u1_u6_n122 ) , .A1( u1_u1_u6_n94 ) , .A2( u1_u1_u6_n97 ) );
  INV_X1 u1_u1_u6_U59 (.A( u1_u1_u6_n139 ) , .ZN( u1_u1_u6_n160 ) );
  AOI22_X1 u1_u1_u6_U6 (.B2( u1_u1_u6_n101 ) , .A1( u1_u1_u6_n102 ) , .ZN( u1_u1_u6_n103 ) , .B1( u1_u1_u6_n160 ) , .A2( u1_u1_u6_n161 ) );
  NAND2_X1 u1_u1_u6_U60 (.ZN( u1_u1_u6_n113 ) , .A1( u1_u1_u6_n96 ) , .A2( u1_u1_u6_n98 ) );
  NOR2_X1 u1_u1_u6_U61 (.A2( u1_u1_X_40 ) , .A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n126 ) );
  NOR2_X1 u1_u1_u6_U62 (.A2( u1_u1_X_39 ) , .A1( u1_u1_X_42 ) , .ZN( u1_u1_u6_n92 ) );
  NOR2_X1 u1_u1_u6_U63 (.A2( u1_u1_X_39 ) , .A1( u1_u1_u6_n156 ) , .ZN( u1_u1_u6_n97 ) );
  NOR2_X1 u1_u1_u6_U64 (.A2( u1_u1_X_38 ) , .A1( u1_u1_u6_n165 ) , .ZN( u1_u1_u6_n95 ) );
  NOR2_X1 u1_u1_u6_U65 (.A2( u1_u1_X_41 ) , .ZN( u1_u1_u6_n111 ) , .A1( u1_u1_u6_n157 ) );
  NOR2_X1 u1_u1_u6_U66 (.A2( u1_u1_X_37 ) , .A1( u1_u1_u6_n162 ) , .ZN( u1_u1_u6_n94 ) );
  NOR2_X1 u1_u1_u6_U67 (.A2( u1_u1_X_37 ) , .A1( u1_u1_X_38 ) , .ZN( u1_u1_u6_n91 ) );
  NAND2_X1 u1_u1_u6_U68 (.A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n144 ) , .A2( u1_u1_u6_n157 ) );
  NAND2_X1 u1_u1_u6_U69 (.A2( u1_u1_X_40 ) , .A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n139 ) );
  NOR2_X1 u1_u1_u6_U7 (.A1( u1_u1_u6_n118 ) , .ZN( u1_u1_u6_n143 ) , .A2( u1_u1_u6_n168 ) );
  AND2_X1 u1_u1_u6_U70 (.A1( u1_u1_X_39 ) , .A2( u1_u1_u6_n156 ) , .ZN( u1_u1_u6_n96 ) );
  AND2_X1 u1_u1_u6_U71 (.A1( u1_u1_X_39 ) , .A2( u1_u1_X_42 ) , .ZN( u1_u1_u6_n99 ) );
  INV_X1 u1_u1_u6_U72 (.A( u1_u1_X_40 ) , .ZN( u1_u1_u6_n157 ) );
  INV_X1 u1_u1_u6_U73 (.A( u1_u1_X_37 ) , .ZN( u1_u1_u6_n165 ) );
  INV_X1 u1_u1_u6_U74 (.A( u1_u1_X_38 ) , .ZN( u1_u1_u6_n162 ) );
  INV_X1 u1_u1_u6_U75 (.A( u1_u1_X_42 ) , .ZN( u1_u1_u6_n156 ) );
  NAND4_X1 u1_u1_u6_U76 (.ZN( u1_out1_32 ) , .A4( u1_u1_u6_n103 ) , .A3( u1_u1_u6_n104 ) , .A2( u1_u1_u6_n105 ) , .A1( u1_u1_u6_n106 ) );
  AOI22_X1 u1_u1_u6_U77 (.ZN( u1_u1_u6_n105 ) , .A2( u1_u1_u6_n108 ) , .A1( u1_u1_u6_n118 ) , .B2( u1_u1_u6_n126 ) , .B1( u1_u1_u6_n171 ) );
  AOI22_X1 u1_u1_u6_U78 (.ZN( u1_u1_u6_n104 ) , .A1( u1_u1_u6_n111 ) , .B1( u1_u1_u6_n124 ) , .B2( u1_u1_u6_n151 ) , .A2( u1_u1_u6_n93 ) );
  NAND4_X1 u1_u1_u6_U79 (.ZN( u1_out1_12 ) , .A4( u1_u1_u6_n114 ) , .A3( u1_u1_u6_n115 ) , .A2( u1_u1_u6_n116 ) , .A1( u1_u1_u6_n117 ) );
  OAI21_X1 u1_u1_u6_U8 (.A( u1_u1_u6_n159 ) , .B1( u1_u1_u6_n169 ) , .B2( u1_u1_u6_n173 ) , .ZN( u1_u1_u6_n90 ) );
  OAI22_X1 u1_u1_u6_U80 (.B2( u1_u1_u6_n111 ) , .ZN( u1_u1_u6_n116 ) , .B1( u1_u1_u6_n126 ) , .A2( u1_u1_u6_n164 ) , .A1( u1_u1_u6_n167 ) );
  OAI21_X1 u1_u1_u6_U81 (.A( u1_u1_u6_n108 ) , .ZN( u1_u1_u6_n117 ) , .B2( u1_u1_u6_n141 ) , .B1( u1_u1_u6_n163 ) );
  OAI211_X1 u1_u1_u6_U82 (.ZN( u1_out1_7 ) , .B( u1_u1_u6_n153 ) , .C2( u1_u1_u6_n154 ) , .C1( u1_u1_u6_n155 ) , .A( u1_u1_u6_n174 ) );
  NOR3_X1 u1_u1_u6_U83 (.A1( u1_u1_u6_n141 ) , .ZN( u1_u1_u6_n154 ) , .A3( u1_u1_u6_n164 ) , .A2( u1_u1_u6_n171 ) );
  AOI211_X1 u1_u1_u6_U84 (.B( u1_u1_u6_n149 ) , .A( u1_u1_u6_n150 ) , .C2( u1_u1_u6_n151 ) , .C1( u1_u1_u6_n152 ) , .ZN( u1_u1_u6_n153 ) );
  OAI211_X1 u1_u1_u6_U85 (.ZN( u1_out1_22 ) , .B( u1_u1_u6_n137 ) , .A( u1_u1_u6_n138 ) , .C2( u1_u1_u6_n139 ) , .C1( u1_u1_u6_n140 ) );
  AND4_X1 u1_u1_u6_U86 (.A3( u1_u1_u6_n119 ) , .A1( u1_u1_u6_n120 ) , .A4( u1_u1_u6_n129 ) , .ZN( u1_u1_u6_n140 ) , .A2( u1_u1_u6_n143 ) );
  AOI22_X1 u1_u1_u6_U87 (.B1( u1_u1_u6_n124 ) , .A2( u1_u1_u6_n125 ) , .A1( u1_u1_u6_n126 ) , .ZN( u1_u1_u6_n138 ) , .B2( u1_u1_u6_n161 ) );
  NAND3_X1 u1_u1_u6_U88 (.A2( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n125 ) , .A1( u1_u1_u6_n130 ) , .A3( u1_u1_u6_n131 ) );
  NAND3_X1 u1_u1_u6_U89 (.A3( u1_u1_u6_n133 ) , .ZN( u1_u1_u6_n141 ) , .A1( u1_u1_u6_n145 ) , .A2( u1_u1_u6_n148 ) );
  INV_X1 u1_u1_u6_U9 (.ZN( u1_u1_u6_n172 ) , .A( u1_u1_u6_n88 ) );
  NAND3_X1 u1_u1_u6_U90 (.ZN( u1_u1_u6_n101 ) , .A3( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n121 ) , .A1( u1_u1_u6_n127 ) );
  NAND3_X1 u1_u1_u6_U91 (.ZN( u1_u1_u6_n102 ) , .A3( u1_u1_u6_n130 ) , .A2( u1_u1_u6_n145 ) , .A1( u1_u1_u6_n166 ) );
  NAND3_X1 u1_u1_u6_U92 (.A3( u1_u1_u6_n113 ) , .A1( u1_u1_u6_n119 ) , .A2( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n93 ) );
  NAND3_X1 u1_u1_u6_U93 (.ZN( u1_u1_u6_n142 ) , .A2( u1_u1_u6_n172 ) , .A3( u1_u1_u6_n89 ) , .A1( u1_u1_u6_n90 ) );
  AND3_X1 u1_u1_u7_U10 (.A3( u1_u1_u7_n110 ) , .A2( u1_u1_u7_n127 ) , .A1( u1_u1_u7_n132 ) , .ZN( u1_u1_u7_n92 ) );
  OAI21_X1 u1_u1_u7_U11 (.A( u1_u1_u7_n161 ) , .B1( u1_u1_u7_n168 ) , .B2( u1_u1_u7_n173 ) , .ZN( u1_u1_u7_n91 ) );
  AOI211_X1 u1_u1_u7_U12 (.A( u1_u1_u7_n117 ) , .ZN( u1_u1_u7_n118 ) , .C2( u1_u1_u7_n126 ) , .C1( u1_u1_u7_n177 ) , .B( u1_u1_u7_n180 ) );
  OAI22_X1 u1_u1_u7_U13 (.B1( u1_u1_u7_n115 ) , .ZN( u1_u1_u7_n117 ) , .A2( u1_u1_u7_n133 ) , .A1( u1_u1_u7_n137 ) , .B2( u1_u1_u7_n162 ) );
  INV_X1 u1_u1_u7_U14 (.A( u1_u1_u7_n116 ) , .ZN( u1_u1_u7_n180 ) );
  NOR3_X1 u1_u1_u7_U15 (.ZN( u1_u1_u7_n115 ) , .A3( u1_u1_u7_n145 ) , .A2( u1_u1_u7_n168 ) , .A1( u1_u1_u7_n169 ) );
  OAI211_X1 u1_u1_u7_U16 (.B( u1_u1_u7_n122 ) , .A( u1_u1_u7_n123 ) , .C2( u1_u1_u7_n124 ) , .ZN( u1_u1_u7_n154 ) , .C1( u1_u1_u7_n162 ) );
  AOI222_X1 u1_u1_u7_U17 (.ZN( u1_u1_u7_n122 ) , .C2( u1_u1_u7_n126 ) , .C1( u1_u1_u7_n145 ) , .B1( u1_u1_u7_n161 ) , .A2( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n170 ) , .A1( u1_u1_u7_n176 ) );
  INV_X1 u1_u1_u7_U18 (.A( u1_u1_u7_n133 ) , .ZN( u1_u1_u7_n176 ) );
  NOR3_X1 u1_u1_u7_U19 (.A2( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n135 ) , .ZN( u1_u1_u7_n136 ) , .A3( u1_u1_u7_n171 ) );
  NOR2_X1 u1_u1_u7_U20 (.A1( u1_u1_u7_n130 ) , .A2( u1_u1_u7_n134 ) , .ZN( u1_u1_u7_n153 ) );
  INV_X1 u1_u1_u7_U21 (.A( u1_u1_u7_n101 ) , .ZN( u1_u1_u7_n165 ) );
  NOR2_X1 u1_u1_u7_U22 (.ZN( u1_u1_u7_n111 ) , .A2( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n169 ) );
  AOI21_X1 u1_u1_u7_U23 (.ZN( u1_u1_u7_n104 ) , .B2( u1_u1_u7_n112 ) , .B1( u1_u1_u7_n127 ) , .A( u1_u1_u7_n164 ) );
  AOI21_X1 u1_u1_u7_U24 (.ZN( u1_u1_u7_n106 ) , .B1( u1_u1_u7_n133 ) , .B2( u1_u1_u7_n146 ) , .A( u1_u1_u7_n162 ) );
  AOI21_X1 u1_u1_u7_U25 (.A( u1_u1_u7_n101 ) , .ZN( u1_u1_u7_n107 ) , .B2( u1_u1_u7_n128 ) , .B1( u1_u1_u7_n175 ) );
  INV_X1 u1_u1_u7_U26 (.A( u1_u1_u7_n138 ) , .ZN( u1_u1_u7_n171 ) );
  INV_X1 u1_u1_u7_U27 (.A( u1_u1_u7_n131 ) , .ZN( u1_u1_u7_n177 ) );
  INV_X1 u1_u1_u7_U28 (.A( u1_u1_u7_n110 ) , .ZN( u1_u1_u7_n174 ) );
  NAND2_X1 u1_u1_u7_U29 (.A1( u1_u1_u7_n129 ) , .A2( u1_u1_u7_n132 ) , .ZN( u1_u1_u7_n149 ) );
  OAI21_X1 u1_u1_u7_U3 (.ZN( u1_u1_u7_n159 ) , .A( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n171 ) , .B1( u1_u1_u7_n174 ) );
  NAND2_X1 u1_u1_u7_U30 (.A1( u1_u1_u7_n113 ) , .A2( u1_u1_u7_n124 ) , .ZN( u1_u1_u7_n130 ) );
  INV_X1 u1_u1_u7_U31 (.A( u1_u1_u7_n112 ) , .ZN( u1_u1_u7_n173 ) );
  INV_X1 u1_u1_u7_U32 (.A( u1_u1_u7_n128 ) , .ZN( u1_u1_u7_n168 ) );
  INV_X1 u1_u1_u7_U33 (.A( u1_u1_u7_n148 ) , .ZN( u1_u1_u7_n169 ) );
  INV_X1 u1_u1_u7_U34 (.A( u1_u1_u7_n127 ) , .ZN( u1_u1_u7_n179 ) );
  NOR2_X1 u1_u1_u7_U35 (.ZN( u1_u1_u7_n101 ) , .A2( u1_u1_u7_n150 ) , .A1( u1_u1_u7_n156 ) );
  AOI211_X1 u1_u1_u7_U36 (.B( u1_u1_u7_n154 ) , .A( u1_u1_u7_n155 ) , .C1( u1_u1_u7_n156 ) , .ZN( u1_u1_u7_n157 ) , .C2( u1_u1_u7_n172 ) );
  INV_X1 u1_u1_u7_U37 (.A( u1_u1_u7_n153 ) , .ZN( u1_u1_u7_n172 ) );
  AOI211_X1 u1_u1_u7_U38 (.B( u1_u1_u7_n139 ) , .A( u1_u1_u7_n140 ) , .C2( u1_u1_u7_n141 ) , .ZN( u1_u1_u7_n142 ) , .C1( u1_u1_u7_n156 ) );
  NAND4_X1 u1_u1_u7_U39 (.A3( u1_u1_u7_n127 ) , .A2( u1_u1_u7_n128 ) , .A1( u1_u1_u7_n129 ) , .ZN( u1_u1_u7_n141 ) , .A4( u1_u1_u7_n147 ) );
  INV_X1 u1_u1_u7_U4 (.A( u1_u1_u7_n111 ) , .ZN( u1_u1_u7_n170 ) );
  AOI21_X1 u1_u1_u7_U40 (.A( u1_u1_u7_n137 ) , .B1( u1_u1_u7_n138 ) , .ZN( u1_u1_u7_n139 ) , .B2( u1_u1_u7_n146 ) );
  OAI22_X1 u1_u1_u7_U41 (.B1( u1_u1_u7_n136 ) , .ZN( u1_u1_u7_n140 ) , .A1( u1_u1_u7_n153 ) , .B2( u1_u1_u7_n162 ) , .A2( u1_u1_u7_n164 ) );
  AOI21_X1 u1_u1_u7_U42 (.ZN( u1_u1_u7_n123 ) , .B1( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n177 ) , .A( u1_u1_u7_n97 ) );
  AOI21_X1 u1_u1_u7_U43 (.B2( u1_u1_u7_n113 ) , .B1( u1_u1_u7_n124 ) , .A( u1_u1_u7_n125 ) , .ZN( u1_u1_u7_n97 ) );
  INV_X1 u1_u1_u7_U44 (.A( u1_u1_u7_n125 ) , .ZN( u1_u1_u7_n161 ) );
  INV_X1 u1_u1_u7_U45 (.A( u1_u1_u7_n152 ) , .ZN( u1_u1_u7_n162 ) );
  AOI22_X1 u1_u1_u7_U46 (.A2( u1_u1_u7_n114 ) , .ZN( u1_u1_u7_n119 ) , .B1( u1_u1_u7_n130 ) , .A1( u1_u1_u7_n156 ) , .B2( u1_u1_u7_n165 ) );
  NAND2_X1 u1_u1_u7_U47 (.A2( u1_u1_u7_n112 ) , .ZN( u1_u1_u7_n114 ) , .A1( u1_u1_u7_n175 ) );
  AND2_X1 u1_u1_u7_U48 (.ZN( u1_u1_u7_n145 ) , .A2( u1_u1_u7_n98 ) , .A1( u1_u1_u7_n99 ) );
  NOR2_X1 u1_u1_u7_U49 (.ZN( u1_u1_u7_n137 ) , .A1( u1_u1_u7_n150 ) , .A2( u1_u1_u7_n161 ) );
  INV_X1 u1_u1_u7_U5 (.A( u1_u1_u7_n149 ) , .ZN( u1_u1_u7_n175 ) );
  AOI21_X1 u1_u1_u7_U50 (.ZN( u1_u1_u7_n105 ) , .B2( u1_u1_u7_n110 ) , .A( u1_u1_u7_n125 ) , .B1( u1_u1_u7_n147 ) );
  NAND2_X1 u1_u1_u7_U51 (.ZN( u1_u1_u7_n146 ) , .A1( u1_u1_u7_n95 ) , .A2( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U52 (.A2( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n147 ) , .A1( u1_u1_u7_n93 ) );
  NAND2_X1 u1_u1_u7_U53 (.A1( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n127 ) , .A2( u1_u1_u7_n99 ) );
  OR2_X1 u1_u1_u7_U54 (.ZN( u1_u1_u7_n126 ) , .A2( u1_u1_u7_n152 ) , .A1( u1_u1_u7_n156 ) );
  NAND2_X1 u1_u1_u7_U55 (.A2( u1_u1_u7_n102 ) , .A1( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n133 ) );
  NAND2_X1 u1_u1_u7_U56 (.ZN( u1_u1_u7_n112 ) , .A2( u1_u1_u7_n96 ) , .A1( u1_u1_u7_n99 ) );
  NAND2_X1 u1_u1_u7_U57 (.A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n128 ) , .A1( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U58 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n113 ) , .A2( u1_u1_u7_n93 ) );
  NAND2_X1 u1_u1_u7_U59 (.A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n124 ) , .A1( u1_u1_u7_n96 ) );
  INV_X1 u1_u1_u7_U6 (.A( u1_u1_u7_n154 ) , .ZN( u1_u1_u7_n178 ) );
  NAND2_X1 u1_u1_u7_U60 (.ZN( u1_u1_u7_n110 ) , .A1( u1_u1_u7_n95 ) , .A2( u1_u1_u7_n96 ) );
  INV_X1 u1_u1_u7_U61 (.A( u1_u1_u7_n150 ) , .ZN( u1_u1_u7_n164 ) );
  AND2_X1 u1_u1_u7_U62 (.ZN( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n93 ) , .A2( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U63 (.A1( u1_u1_u7_n100 ) , .A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n129 ) );
  NAND2_X1 u1_u1_u7_U64 (.A2( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n131 ) , .A1( u1_u1_u7_n95 ) );
  NAND2_X1 u1_u1_u7_U65 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n138 ) , .A2( u1_u1_u7_n99 ) );
  NAND2_X1 u1_u1_u7_U66 (.ZN( u1_u1_u7_n132 ) , .A1( u1_u1_u7_n93 ) , .A2( u1_u1_u7_n96 ) );
  NAND2_X1 u1_u1_u7_U67 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n148 ) , .A2( u1_u1_u7_n95 ) );
  NOR2_X1 u1_u1_u7_U68 (.A2( u1_u1_X_47 ) , .ZN( u1_u1_u7_n150 ) , .A1( u1_u1_u7_n163 ) );
  NOR2_X1 u1_u1_u7_U69 (.A2( u1_u1_X_43 ) , .A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n103 ) );
  AOI211_X1 u1_u1_u7_U7 (.ZN( u1_u1_u7_n116 ) , .A( u1_u1_u7_n155 ) , .C1( u1_u1_u7_n161 ) , .C2( u1_u1_u7_n171 ) , .B( u1_u1_u7_n94 ) );
  NOR2_X1 u1_u1_u7_U70 (.A2( u1_u1_X_48 ) , .A1( u1_u1_u7_n166 ) , .ZN( u1_u1_u7_n95 ) );
  NOR2_X1 u1_u1_u7_U71 (.A2( u1_u1_X_45 ) , .A1( u1_u1_X_48 ) , .ZN( u1_u1_u7_n99 ) );
  NOR2_X1 u1_u1_u7_U72 (.A2( u1_u1_X_44 ) , .A1( u1_u1_u7_n167 ) , .ZN( u1_u1_u7_n98 ) );
  NOR2_X1 u1_u1_u7_U73 (.A2( u1_u1_X_46 ) , .A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n152 ) );
  AND2_X1 u1_u1_u7_U74 (.A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n156 ) , .A2( u1_u1_u7_n163 ) );
  NAND2_X1 u1_u1_u7_U75 (.A2( u1_u1_X_46 ) , .A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n125 ) );
  AND2_X1 u1_u1_u7_U76 (.A2( u1_u1_X_45 ) , .A1( u1_u1_X_48 ) , .ZN( u1_u1_u7_n102 ) );
  AND2_X1 u1_u1_u7_U77 (.A2( u1_u1_X_43 ) , .A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n96 ) );
  AND2_X1 u1_u1_u7_U78 (.A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n100 ) , .A2( u1_u1_u7_n167 ) );
  AND2_X1 u1_u1_u7_U79 (.A1( u1_u1_X_48 ) , .A2( u1_u1_u7_n166 ) , .ZN( u1_u1_u7_n93 ) );
  OAI222_X1 u1_u1_u7_U8 (.C2( u1_u1_u7_n101 ) , .B2( u1_u1_u7_n111 ) , .A1( u1_u1_u7_n113 ) , .C1( u1_u1_u7_n146 ) , .A2( u1_u1_u7_n162 ) , .B1( u1_u1_u7_n164 ) , .ZN( u1_u1_u7_n94 ) );
  INV_X1 u1_u1_u7_U80 (.A( u1_u1_X_46 ) , .ZN( u1_u1_u7_n163 ) );
  INV_X1 u1_u1_u7_U81 (.A( u1_u1_X_43 ) , .ZN( u1_u1_u7_n167 ) );
  INV_X1 u1_u1_u7_U82 (.A( u1_u1_X_45 ) , .ZN( u1_u1_u7_n166 ) );
  NAND4_X1 u1_u1_u7_U83 (.ZN( u1_out1_5 ) , .A4( u1_u1_u7_n108 ) , .A3( u1_u1_u7_n109 ) , .A1( u1_u1_u7_n116 ) , .A2( u1_u1_u7_n123 ) );
  AOI22_X1 u1_u1_u7_U84 (.ZN( u1_u1_u7_n109 ) , .A2( u1_u1_u7_n126 ) , .B2( u1_u1_u7_n145 ) , .B1( u1_u1_u7_n156 ) , .A1( u1_u1_u7_n171 ) );
  NOR4_X1 u1_u1_u7_U85 (.A4( u1_u1_u7_n104 ) , .A3( u1_u1_u7_n105 ) , .A2( u1_u1_u7_n106 ) , .A1( u1_u1_u7_n107 ) , .ZN( u1_u1_u7_n108 ) );
  NAND4_X1 u1_u1_u7_U86 (.ZN( u1_out1_27 ) , .A4( u1_u1_u7_n118 ) , .A3( u1_u1_u7_n119 ) , .A2( u1_u1_u7_n120 ) , .A1( u1_u1_u7_n121 ) );
  OAI21_X1 u1_u1_u7_U87 (.ZN( u1_u1_u7_n121 ) , .B2( u1_u1_u7_n145 ) , .A( u1_u1_u7_n150 ) , .B1( u1_u1_u7_n174 ) );
  OAI21_X1 u1_u1_u7_U88 (.ZN( u1_u1_u7_n120 ) , .A( u1_u1_u7_n161 ) , .B2( u1_u1_u7_n170 ) , .B1( u1_u1_u7_n179 ) );
  NAND4_X1 u1_u1_u7_U89 (.ZN( u1_out1_21 ) , .A4( u1_u1_u7_n157 ) , .A3( u1_u1_u7_n158 ) , .A2( u1_u1_u7_n159 ) , .A1( u1_u1_u7_n160 ) );
  OAI221_X1 u1_u1_u7_U9 (.C1( u1_u1_u7_n101 ) , .C2( u1_u1_u7_n147 ) , .ZN( u1_u1_u7_n155 ) , .B2( u1_u1_u7_n162 ) , .A( u1_u1_u7_n91 ) , .B1( u1_u1_u7_n92 ) );
  OAI21_X1 u1_u1_u7_U90 (.B1( u1_u1_u7_n145 ) , .ZN( u1_u1_u7_n160 ) , .A( u1_u1_u7_n161 ) , .B2( u1_u1_u7_n177 ) );
  AOI22_X1 u1_u1_u7_U91 (.B2( u1_u1_u7_n149 ) , .B1( u1_u1_u7_n150 ) , .A2( u1_u1_u7_n151 ) , .A1( u1_u1_u7_n152 ) , .ZN( u1_u1_u7_n158 ) );
  NAND4_X1 u1_u1_u7_U92 (.ZN( u1_out1_15 ) , .A4( u1_u1_u7_n142 ) , .A3( u1_u1_u7_n143 ) , .A2( u1_u1_u7_n144 ) , .A1( u1_u1_u7_n178 ) );
  OR2_X1 u1_u1_u7_U93 (.A2( u1_u1_u7_n125 ) , .A1( u1_u1_u7_n129 ) , .ZN( u1_u1_u7_n144 ) );
  AOI22_X1 u1_u1_u7_U94 (.A2( u1_u1_u7_n126 ) , .ZN( u1_u1_u7_n143 ) , .B2( u1_u1_u7_n165 ) , .B1( u1_u1_u7_n173 ) , .A1( u1_u1_u7_n174 ) );
  NAND3_X1 u1_u1_u7_U95 (.A3( u1_u1_u7_n146 ) , .A2( u1_u1_u7_n147 ) , .A1( u1_u1_u7_n148 ) , .ZN( u1_u1_u7_n151 ) );
  NAND3_X1 u1_u1_u7_U96 (.A3( u1_u1_u7_n131 ) , .A2( u1_u1_u7_n132 ) , .A1( u1_u1_u7_n133 ) , .ZN( u1_u1_u7_n135 ) );
  XOR2_X1 u1_u2_U11 (.B( u1_K3_44 ) , .A( u1_R1_29 ) , .Z( u1_u2_X_44 ) );
  XOR2_X1 u1_u2_U12 (.B( u1_K3_43 ) , .A( u1_R1_28 ) , .Z( u1_u2_X_43 ) );
  XOR2_X1 u1_u2_U13 (.B( u1_K3_42 ) , .A( u1_R1_29 ) , .Z( u1_u2_X_42 ) );
  XOR2_X1 u1_u2_U14 (.B( u1_K3_41 ) , .A( u1_R1_28 ) , .Z( u1_u2_X_41 ) );
  XOR2_X1 u1_u2_U18 (.B( u1_K3_38 ) , .A( u1_R1_25 ) , .Z( u1_u2_X_38 ) );
  XOR2_X1 u1_u2_U19 (.B( u1_K3_37 ) , .A( u1_R1_24 ) , .Z( u1_u2_X_37 ) );
  XOR2_X1 u1_u2_U27 (.B( u1_K3_2 ) , .A( u1_R1_1 ) , .Z( u1_u2_X_2 ) );
  XOR2_X1 u1_u2_U38 (.B( u1_K3_1 ) , .A( u1_R1_32 ) , .Z( u1_u2_X_1 ) );
  XOR2_X1 u1_u2_U4 (.B( u1_K3_6 ) , .A( u1_R1_5 ) , .Z( u1_u2_X_6 ) );
  XOR2_X1 u1_u2_U5 (.B( u1_K3_5 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_5 ) );
  XOR2_X1 u1_u2_U7 (.B( u1_K3_48 ) , .A( u1_R1_1 ) , .Z( u1_u2_X_48 ) );
  XOR2_X1 u1_u2_U8 (.B( u1_K3_47 ) , .A( u1_R1_32 ) , .Z( u1_u2_X_47 ) );
  AND3_X1 u1_u2_u0_U10 (.A2( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n127 ) , .A3( u1_u2_u0_n130 ) , .A1( u1_u2_u0_n148 ) );
  NAND2_X1 u1_u2_u0_U11 (.ZN( u1_u2_u0_n113 ) , .A1( u1_u2_u0_n139 ) , .A2( u1_u2_u0_n149 ) );
  AND2_X1 u1_u2_u0_U12 (.ZN( u1_u2_u0_n107 ) , .A1( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n140 ) );
  AND2_X1 u1_u2_u0_U13 (.A2( u1_u2_u0_n129 ) , .A1( u1_u2_u0_n130 ) , .ZN( u1_u2_u0_n151 ) );
  AND2_X1 u1_u2_u0_U14 (.A1( u1_u2_u0_n108 ) , .A2( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U15 (.A( u1_u2_u0_n143 ) , .ZN( u1_u2_u0_n173 ) );
  NOR2_X1 u1_u2_u0_U16 (.A2( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n147 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U17 (.ZN( u1_u2_u0_n172 ) , .A( u1_u2_u0_n88 ) );
  OAI222_X1 u1_u2_u0_U18 (.C1( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n125 ) , .B2( u1_u2_u0_n128 ) , .B1( u1_u2_u0_n144 ) , .A2( u1_u2_u0_n158 ) , .C2( u1_u2_u0_n161 ) , .ZN( u1_u2_u0_n88 ) );
  NOR2_X1 u1_u2_u0_U19 (.A1( u1_u2_u0_n163 ) , .A2( u1_u2_u0_n164 ) , .ZN( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U20 (.B1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n132 ) , .A( u1_u2_u0_n165 ) , .B2( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U21 (.A( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n165 ) );
  OAI221_X1 u1_u2_u0_U22 (.C1( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n122 ) , .B2( u1_u2_u0_n127 ) , .A( u1_u2_u0_n143 ) , .B1( u1_u2_u0_n144 ) , .C2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U23 (.B1( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n126 ) , .A1( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n146 ) , .B2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U24 (.B1( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n147 ) , .A2( u1_u2_u0_n90 ) , .ZN( u1_u2_u0_n91 ) );
  AND3_X1 u1_u2_u0_U25 (.A3( u1_u2_u0_n121 ) , .A2( u1_u2_u0_n125 ) , .A1( u1_u2_u0_n148 ) , .ZN( u1_u2_u0_n90 ) );
  INV_X1 u1_u2_u0_U26 (.A( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n161 ) );
  NOR2_X1 u1_u2_u0_U27 (.A1( u1_u2_u0_n120 ) , .ZN( u1_u2_u0_n143 ) , .A2( u1_u2_u0_n167 ) );
  OAI221_X1 u1_u2_u0_U28 (.C1( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n120 ) , .B1( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n141 ) , .C2( u1_u2_u0_n147 ) , .A( u1_u2_u0_n172 ) );
  AOI211_X1 u1_u2_u0_U29 (.B( u1_u2_u0_n115 ) , .A( u1_u2_u0_n116 ) , .C2( u1_u2_u0_n117 ) , .C1( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n119 ) );
  INV_X1 u1_u2_u0_U3 (.A( u1_u2_u0_n113 ) , .ZN( u1_u2_u0_n166 ) );
  AOI22_X1 u1_u2_u0_U30 (.B2( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n110 ) , .ZN( u1_u2_u0_n111 ) , .B1( u1_u2_u0_n118 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U31 (.A( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U32 (.ZN( u1_u2_u0_n104 ) , .B1( u1_u2_u0_n107 ) , .B2( u1_u2_u0_n141 ) , .A( u1_u2_u0_n144 ) );
  AOI21_X1 u1_u2_u0_U33 (.B1( u1_u2_u0_n127 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n96 ) );
  AOI21_X1 u1_u2_u0_U34 (.ZN( u1_u2_u0_n116 ) , .B2( u1_u2_u0_n142 ) , .A( u1_u2_u0_n144 ) , .B1( u1_u2_u0_n166 ) );
  NAND2_X1 u1_u2_u0_U35 (.A1( u1_u2_u0_n100 ) , .A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n125 ) );
  NAND2_X1 u1_u2_u0_U36 (.A1( u1_u2_u0_n101 ) , .A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n150 ) );
  INV_X1 u1_u2_u0_U37 (.A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n160 ) );
  NAND2_X1 u1_u2_u0_U38 (.A1( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n128 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U39 (.A1( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n129 ) , .A2( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U4 (.B1( u1_u2_u0_n114 ) , .ZN( u1_u2_u0_n115 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n161 ) );
  NAND2_X1 u1_u2_u0_U40 (.A2( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U41 (.A2( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n139 ) );
  NAND2_X1 u1_u2_u0_U42 (.ZN( u1_u2_u0_n148 ) , .A1( u1_u2_u0_n93 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U43 (.A2( u1_u2_u0_n102 ) , .A1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n149 ) );
  NAND2_X1 u1_u2_u0_U44 (.A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n114 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U45 (.A2( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n121 ) , .A1( u1_u2_u0_n93 ) );
  NAND2_X1 u1_u2_u0_U46 (.ZN( u1_u2_u0_n112 ) , .A2( u1_u2_u0_n92 ) , .A1( u1_u2_u0_n93 ) );
  OR3_X1 u1_u2_u0_U47 (.A3( u1_u2_u0_n152 ) , .A2( u1_u2_u0_n153 ) , .A1( u1_u2_u0_n154 ) , .ZN( u1_u2_u0_n155 ) );
  AOI21_X1 u1_u2_u0_U48 (.B2( u1_u2_u0_n150 ) , .B1( u1_u2_u0_n151 ) , .ZN( u1_u2_u0_n152 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U49 (.A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n145 ) , .B1( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n154 ) );
  AOI21_X1 u1_u2_u0_U5 (.B2( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n134 ) , .B1( u1_u2_u0_n151 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U50 (.A( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n148 ) , .B1( u1_u2_u0_n149 ) , .ZN( u1_u2_u0_n153 ) );
  INV_X1 u1_u2_u0_U51 (.ZN( u1_u2_u0_n171 ) , .A( u1_u2_u0_n99 ) );
  OAI211_X1 u1_u2_u0_U52 (.C2( u1_u2_u0_n140 ) , .C1( u1_u2_u0_n161 ) , .A( u1_u2_u0_n169 ) , .B( u1_u2_u0_n98 ) , .ZN( u1_u2_u0_n99 ) );
  AOI211_X1 u1_u2_u0_U53 (.C1( u1_u2_u0_n118 ) , .A( u1_u2_u0_n123 ) , .B( u1_u2_u0_n96 ) , .C2( u1_u2_u0_n97 ) , .ZN( u1_u2_u0_n98 ) );
  INV_X1 u1_u2_u0_U54 (.ZN( u1_u2_u0_n169 ) , .A( u1_u2_u0_n91 ) );
  NOR2_X1 u1_u2_u0_U55 (.A2( u1_u2_X_6 ) , .ZN( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U56 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n118 ) );
  NOR2_X1 u1_u2_u0_U57 (.A2( u1_u2_X_2 ) , .ZN( u1_u2_u0_n103 ) , .A1( u1_u2_u0_n164 ) );
  NOR2_X1 u1_u2_u0_U58 (.A2( u1_u2_X_1 ) , .A1( u1_u2_X_2 ) , .ZN( u1_u2_u0_n92 ) );
  NOR2_X1 u1_u2_u0_U59 (.A2( u1_u2_X_1 ) , .ZN( u1_u2_u0_n101 ) , .A1( u1_u2_u0_n163 ) );
  NOR2_X1 u1_u2_u0_U6 (.A1( u1_u2_u0_n108 ) , .ZN( u1_u2_u0_n123 ) , .A2( u1_u2_u0_n158 ) );
  NAND2_X1 u1_u2_u0_U60 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n144 ) );
  NOR2_X1 u1_u2_u0_U61 (.A2( u1_u2_X_5 ) , .ZN( u1_u2_u0_n136 ) , .A1( u1_u2_u0_n159 ) );
  NAND2_X1 u1_u2_u0_U62 (.A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n159 ) );
  AND2_X1 u1_u2_u0_U63 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n102 ) );
  AND2_X1 u1_u2_u0_U64 (.A1( u1_u2_X_6 ) , .A2( u1_u2_u0_n162 ) , .ZN( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U65 (.A( u1_u2_X_4 ) , .ZN( u1_u2_u0_n159 ) );
  INV_X1 u1_u2_u0_U66 (.A( u1_u2_X_1 ) , .ZN( u1_u2_u0_n164 ) );
  INV_X1 u1_u2_u0_U67 (.A( u1_u2_X_2 ) , .ZN( u1_u2_u0_n163 ) );
  INV_X1 u1_u2_u0_U68 (.ZN( u1_u2_u0_n174 ) , .A( u1_u2_u0_n89 ) );
  AOI211_X1 u1_u2_u0_U69 (.B( u1_u2_u0_n104 ) , .A( u1_u2_u0_n105 ) , .ZN( u1_u2_u0_n106 ) , .C2( u1_u2_u0_n113 ) , .C1( u1_u2_u0_n160 ) );
  OAI21_X1 u1_u2_u0_U7 (.B1( u1_u2_u0_n150 ) , .B2( u1_u2_u0_n158 ) , .A( u1_u2_u0_n172 ) , .ZN( u1_u2_u0_n89 ) );
  OR4_X1 u1_u2_u0_U70 (.ZN( u1_out2_17 ) , .A4( u1_u2_u0_n122 ) , .A2( u1_u2_u0_n123 ) , .A1( u1_u2_u0_n124 ) , .A3( u1_u2_u0_n170 ) );
  AOI21_X1 u1_u2_u0_U71 (.B2( u1_u2_u0_n107 ) , .ZN( u1_u2_u0_n124 ) , .B1( u1_u2_u0_n128 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U72 (.A( u1_u2_u0_n111 ) , .ZN( u1_u2_u0_n170 ) );
  OR4_X1 u1_u2_u0_U73 (.ZN( u1_out2_31 ) , .A4( u1_u2_u0_n155 ) , .A2( u1_u2_u0_n156 ) , .A1( u1_u2_u0_n157 ) , .A3( u1_u2_u0_n173 ) );
  AOI21_X1 u1_u2_u0_U74 (.A( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n139 ) , .B1( u1_u2_u0_n140 ) , .ZN( u1_u2_u0_n157 ) );
  AOI21_X1 u1_u2_u0_U75 (.B2( u1_u2_u0_n141 ) , .B1( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n156 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U76 (.A( u1_u2_u0_n126 ) , .ZN( u1_u2_u0_n168 ) );
  AOI211_X1 u1_u2_u0_U77 (.B( u1_u2_u0_n133 ) , .A( u1_u2_u0_n134 ) , .C2( u1_u2_u0_n135 ) , .C1( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n137 ) );
  AOI21_X1 u1_u2_u0_U78 (.B1( u1_u2_u0_n132 ) , .ZN( u1_u2_u0_n133 ) , .A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n166 ) );
  OAI22_X1 u1_u2_u0_U79 (.ZN( u1_u2_u0_n105 ) , .A2( u1_u2_u0_n132 ) , .B1( u1_u2_u0_n146 ) , .A1( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n161 ) );
  AND2_X1 u1_u2_u0_U8 (.A1( u1_u2_u0_n114 ) , .A2( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n146 ) );
  NAND2_X1 u1_u2_u0_U80 (.ZN( u1_u2_u0_n110 ) , .A2( u1_u2_u0_n132 ) , .A1( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U81 (.A( u1_u2_u0_n119 ) , .ZN( u1_u2_u0_n167 ) );
  NAND2_X1 u1_u2_u0_U82 (.A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U83 (.A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U84 (.ZN( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n92 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U85 (.ZN( u1_u2_u0_n142 ) , .A1( u1_u2_u0_n94 ) , .A2( u1_u2_u0_n95 ) );
  INV_X1 u1_u2_u0_U86 (.A( u1_u2_X_3 ) , .ZN( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U87 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n94 ) );
  NAND3_X1 u1_u2_u0_U88 (.ZN( u1_out2_23 ) , .A3( u1_u2_u0_n137 ) , .A1( u1_u2_u0_n168 ) , .A2( u1_u2_u0_n171 ) );
  NAND3_X1 u1_u2_u0_U89 (.A3( u1_u2_u0_n127 ) , .A2( u1_u2_u0_n128 ) , .ZN( u1_u2_u0_n135 ) , .A1( u1_u2_u0_n150 ) );
  AND2_X1 u1_u2_u0_U9 (.A1( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n141 ) , .A2( u1_u2_u0_n150 ) );
  NAND3_X1 u1_u2_u0_U90 (.ZN( u1_u2_u0_n117 ) , .A3( u1_u2_u0_n132 ) , .A2( u1_u2_u0_n139 ) , .A1( u1_u2_u0_n148 ) );
  NAND3_X1 u1_u2_u0_U91 (.ZN( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n114 ) , .A3( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n149 ) );
  NAND3_X1 u1_u2_u0_U92 (.ZN( u1_out2_9 ) , .A3( u1_u2_u0_n106 ) , .A2( u1_u2_u0_n171 ) , .A1( u1_u2_u0_n174 ) );
  NAND3_X1 u1_u2_u0_U93 (.A2( u1_u2_u0_n128 ) , .A1( u1_u2_u0_n132 ) , .A3( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n97 ) );
  OAI21_X1 u1_u2_u6_U10 (.A( u1_u2_u6_n159 ) , .B1( u1_u2_u6_n169 ) , .B2( u1_u2_u6_n173 ) , .ZN( u1_u2_u6_n90 ) );
  INV_X1 u1_u2_u6_U11 (.ZN( u1_u2_u6_n172 ) , .A( u1_u2_u6_n88 ) );
  AOI22_X1 u1_u2_u6_U12 (.A2( u1_u2_u6_n151 ) , .B2( u1_u2_u6_n161 ) , .A1( u1_u2_u6_n167 ) , .B1( u1_u2_u6_n170 ) , .ZN( u1_u2_u6_n89 ) );
  AOI21_X1 u1_u2_u6_U13 (.ZN( u1_u2_u6_n106 ) , .A( u1_u2_u6_n142 ) , .B2( u1_u2_u6_n159 ) , .B1( u1_u2_u6_n164 ) );
  INV_X1 u1_u2_u6_U14 (.A( u1_u2_u6_n155 ) , .ZN( u1_u2_u6_n161 ) );
  INV_X1 u1_u2_u6_U15 (.A( u1_u2_u6_n128 ) , .ZN( u1_u2_u6_n164 ) );
  NAND2_X1 u1_u2_u6_U16 (.ZN( u1_u2_u6_n110 ) , .A1( u1_u2_u6_n122 ) , .A2( u1_u2_u6_n129 ) );
  NAND2_X1 u1_u2_u6_U17 (.ZN( u1_u2_u6_n124 ) , .A2( u1_u2_u6_n146 ) , .A1( u1_u2_u6_n148 ) );
  INV_X1 u1_u2_u6_U18 (.A( u1_u2_u6_n132 ) , .ZN( u1_u2_u6_n171 ) );
  AND2_X1 u1_u2_u6_U19 (.A1( u1_u2_u6_n100 ) , .ZN( u1_u2_u6_n130 ) , .A2( u1_u2_u6_n147 ) );
  INV_X1 u1_u2_u6_U20 (.A( u1_u2_u6_n127 ) , .ZN( u1_u2_u6_n173 ) );
  INV_X1 u1_u2_u6_U21 (.A( u1_u2_u6_n121 ) , .ZN( u1_u2_u6_n167 ) );
  INV_X1 u1_u2_u6_U22 (.A( u1_u2_u6_n100 ) , .ZN( u1_u2_u6_n169 ) );
  INV_X1 u1_u2_u6_U23 (.A( u1_u2_u6_n123 ) , .ZN( u1_u2_u6_n170 ) );
  INV_X1 u1_u2_u6_U24 (.A( u1_u2_u6_n113 ) , .ZN( u1_u2_u6_n168 ) );
  AND2_X1 u1_u2_u6_U25 (.A1( u1_u2_u6_n107 ) , .A2( u1_u2_u6_n119 ) , .ZN( u1_u2_u6_n133 ) );
  AND2_X1 u1_u2_u6_U26 (.A2( u1_u2_u6_n121 ) , .A1( u1_u2_u6_n122 ) , .ZN( u1_u2_u6_n131 ) );
  AND3_X1 u1_u2_u6_U27 (.ZN( u1_u2_u6_n120 ) , .A2( u1_u2_u6_n127 ) , .A1( u1_u2_u6_n132 ) , .A3( u1_u2_u6_n145 ) );
  INV_X1 u1_u2_u6_U28 (.A( u1_u2_u6_n146 ) , .ZN( u1_u2_u6_n163 ) );
  AOI222_X1 u1_u2_u6_U29 (.ZN( u1_u2_u6_n114 ) , .A1( u1_u2_u6_n118 ) , .A2( u1_u2_u6_n126 ) , .B2( u1_u2_u6_n151 ) , .C2( u1_u2_u6_n159 ) , .C1( u1_u2_u6_n168 ) , .B1( u1_u2_u6_n169 ) );
  INV_X1 u1_u2_u6_U3 (.A( u1_u2_u6_n110 ) , .ZN( u1_u2_u6_n166 ) );
  NOR2_X1 u1_u2_u6_U30 (.A1( u1_u2_u6_n162 ) , .A2( u1_u2_u6_n165 ) , .ZN( u1_u2_u6_n98 ) );
  NAND2_X1 u1_u2_u6_U31 (.A1( u1_u2_u6_n144 ) , .ZN( u1_u2_u6_n151 ) , .A2( u1_u2_u6_n158 ) );
  NAND2_X1 u1_u2_u6_U32 (.ZN( u1_u2_u6_n132 ) , .A1( u1_u2_u6_n91 ) , .A2( u1_u2_u6_n97 ) );
  AOI22_X1 u1_u2_u6_U33 (.B2( u1_u2_u6_n110 ) , .B1( u1_u2_u6_n111 ) , .A1( u1_u2_u6_n112 ) , .ZN( u1_u2_u6_n115 ) , .A2( u1_u2_u6_n161 ) );
  NAND4_X1 u1_u2_u6_U34 (.A3( u1_u2_u6_n109 ) , .ZN( u1_u2_u6_n112 ) , .A4( u1_u2_u6_n132 ) , .A2( u1_u2_u6_n147 ) , .A1( u1_u2_u6_n166 ) );
  NOR2_X1 u1_u2_u6_U35 (.ZN( u1_u2_u6_n109 ) , .A1( u1_u2_u6_n170 ) , .A2( u1_u2_u6_n173 ) );
  NOR2_X1 u1_u2_u6_U36 (.A2( u1_u2_u6_n126 ) , .ZN( u1_u2_u6_n155 ) , .A1( u1_u2_u6_n160 ) );
  NAND2_X1 u1_u2_u6_U37 (.ZN( u1_u2_u6_n146 ) , .A2( u1_u2_u6_n94 ) , .A1( u1_u2_u6_n99 ) );
  AOI21_X1 u1_u2_u6_U38 (.A( u1_u2_u6_n144 ) , .B2( u1_u2_u6_n145 ) , .B1( u1_u2_u6_n146 ) , .ZN( u1_u2_u6_n150 ) );
  INV_X1 u1_u2_u6_U39 (.A( u1_u2_u6_n111 ) , .ZN( u1_u2_u6_n158 ) );
  INV_X1 u1_u2_u6_U4 (.A( u1_u2_u6_n142 ) , .ZN( u1_u2_u6_n174 ) );
  NAND2_X1 u1_u2_u6_U40 (.ZN( u1_u2_u6_n127 ) , .A1( u1_u2_u6_n91 ) , .A2( u1_u2_u6_n92 ) );
  NAND2_X1 u1_u2_u6_U41 (.ZN( u1_u2_u6_n129 ) , .A2( u1_u2_u6_n95 ) , .A1( u1_u2_u6_n96 ) );
  INV_X1 u1_u2_u6_U42 (.A( u1_u2_u6_n144 ) , .ZN( u1_u2_u6_n159 ) );
  NAND2_X1 u1_u2_u6_U43 (.ZN( u1_u2_u6_n145 ) , .A2( u1_u2_u6_n97 ) , .A1( u1_u2_u6_n98 ) );
  NAND2_X1 u1_u2_u6_U44 (.ZN( u1_u2_u6_n148 ) , .A2( u1_u2_u6_n92 ) , .A1( u1_u2_u6_n94 ) );
  NAND2_X1 u1_u2_u6_U45 (.ZN( u1_u2_u6_n108 ) , .A2( u1_u2_u6_n139 ) , .A1( u1_u2_u6_n144 ) );
  NAND2_X1 u1_u2_u6_U46 (.ZN( u1_u2_u6_n121 ) , .A2( u1_u2_u6_n95 ) , .A1( u1_u2_u6_n97 ) );
  NAND2_X1 u1_u2_u6_U47 (.ZN( u1_u2_u6_n107 ) , .A2( u1_u2_u6_n92 ) , .A1( u1_u2_u6_n95 ) );
  AND2_X1 u1_u2_u6_U48 (.ZN( u1_u2_u6_n118 ) , .A2( u1_u2_u6_n91 ) , .A1( u1_u2_u6_n99 ) );
  NAND2_X1 u1_u2_u6_U49 (.ZN( u1_u2_u6_n147 ) , .A2( u1_u2_u6_n98 ) , .A1( u1_u2_u6_n99 ) );
  NAND2_X1 u1_u2_u6_U5 (.A2( u1_u2_u6_n143 ) , .ZN( u1_u2_u6_n152 ) , .A1( u1_u2_u6_n166 ) );
  NAND2_X1 u1_u2_u6_U50 (.ZN( u1_u2_u6_n128 ) , .A1( u1_u2_u6_n94 ) , .A2( u1_u2_u6_n96 ) );
  AOI211_X1 u1_u2_u6_U51 (.B( u1_u2_u6_n134 ) , .A( u1_u2_u6_n135 ) , .C1( u1_u2_u6_n136 ) , .ZN( u1_u2_u6_n137 ) , .C2( u1_u2_u6_n151 ) );
  AOI21_X1 u1_u2_u6_U52 (.B2( u1_u2_u6_n132 ) , .B1( u1_u2_u6_n133 ) , .ZN( u1_u2_u6_n134 ) , .A( u1_u2_u6_n158 ) );
  AOI21_X1 u1_u2_u6_U53 (.B1( u1_u2_u6_n131 ) , .ZN( u1_u2_u6_n135 ) , .A( u1_u2_u6_n144 ) , .B2( u1_u2_u6_n146 ) );
  NAND4_X1 u1_u2_u6_U54 (.A4( u1_u2_u6_n127 ) , .A3( u1_u2_u6_n128 ) , .A2( u1_u2_u6_n129 ) , .A1( u1_u2_u6_n130 ) , .ZN( u1_u2_u6_n136 ) );
  NAND2_X1 u1_u2_u6_U55 (.ZN( u1_u2_u6_n119 ) , .A2( u1_u2_u6_n95 ) , .A1( u1_u2_u6_n99 ) );
  NAND2_X1 u1_u2_u6_U56 (.ZN( u1_u2_u6_n123 ) , .A2( u1_u2_u6_n91 ) , .A1( u1_u2_u6_n96 ) );
  NAND2_X1 u1_u2_u6_U57 (.ZN( u1_u2_u6_n100 ) , .A2( u1_u2_u6_n92 ) , .A1( u1_u2_u6_n98 ) );
  NAND2_X1 u1_u2_u6_U58 (.ZN( u1_u2_u6_n122 ) , .A1( u1_u2_u6_n94 ) , .A2( u1_u2_u6_n97 ) );
  INV_X1 u1_u2_u6_U59 (.A( u1_u2_u6_n139 ) , .ZN( u1_u2_u6_n160 ) );
  AOI22_X1 u1_u2_u6_U6 (.B2( u1_u2_u6_n101 ) , .A1( u1_u2_u6_n102 ) , .ZN( u1_u2_u6_n103 ) , .B1( u1_u2_u6_n160 ) , .A2( u1_u2_u6_n161 ) );
  NAND2_X1 u1_u2_u6_U60 (.ZN( u1_u2_u6_n113 ) , .A1( u1_u2_u6_n96 ) , .A2( u1_u2_u6_n98 ) );
  NOR2_X1 u1_u2_u6_U61 (.A2( u1_u2_X_40 ) , .A1( u1_u2_X_41 ) , .ZN( u1_u2_u6_n126 ) );
  NOR2_X1 u1_u2_u6_U62 (.A2( u1_u2_X_39 ) , .A1( u1_u2_X_42 ) , .ZN( u1_u2_u6_n92 ) );
  NOR2_X1 u1_u2_u6_U63 (.A2( u1_u2_X_39 ) , .A1( u1_u2_u6_n156 ) , .ZN( u1_u2_u6_n97 ) );
  NOR2_X1 u1_u2_u6_U64 (.A2( u1_u2_X_38 ) , .A1( u1_u2_u6_n165 ) , .ZN( u1_u2_u6_n95 ) );
  NOR2_X1 u1_u2_u6_U65 (.A2( u1_u2_X_41 ) , .ZN( u1_u2_u6_n111 ) , .A1( u1_u2_u6_n157 ) );
  NOR2_X1 u1_u2_u6_U66 (.A2( u1_u2_X_37 ) , .A1( u1_u2_u6_n162 ) , .ZN( u1_u2_u6_n94 ) );
  NOR2_X1 u1_u2_u6_U67 (.A2( u1_u2_X_37 ) , .A1( u1_u2_X_38 ) , .ZN( u1_u2_u6_n91 ) );
  NAND2_X1 u1_u2_u6_U68 (.A1( u1_u2_X_41 ) , .ZN( u1_u2_u6_n144 ) , .A2( u1_u2_u6_n157 ) );
  NAND2_X1 u1_u2_u6_U69 (.A2( u1_u2_X_40 ) , .A1( u1_u2_X_41 ) , .ZN( u1_u2_u6_n139 ) );
  NOR2_X1 u1_u2_u6_U7 (.A1( u1_u2_u6_n118 ) , .ZN( u1_u2_u6_n143 ) , .A2( u1_u2_u6_n168 ) );
  AND2_X1 u1_u2_u6_U70 (.A1( u1_u2_X_39 ) , .A2( u1_u2_u6_n156 ) , .ZN( u1_u2_u6_n96 ) );
  AND2_X1 u1_u2_u6_U71 (.A1( u1_u2_X_39 ) , .A2( u1_u2_X_42 ) , .ZN( u1_u2_u6_n99 ) );
  INV_X1 u1_u2_u6_U72 (.A( u1_u2_X_40 ) , .ZN( u1_u2_u6_n157 ) );
  INV_X1 u1_u2_u6_U73 (.A( u1_u2_X_37 ) , .ZN( u1_u2_u6_n165 ) );
  INV_X1 u1_u2_u6_U74 (.A( u1_u2_X_38 ) , .ZN( u1_u2_u6_n162 ) );
  INV_X1 u1_u2_u6_U75 (.A( u1_u2_X_42 ) , .ZN( u1_u2_u6_n156 ) );
  NAND4_X1 u1_u2_u6_U76 (.ZN( u1_out2_32 ) , .A4( u1_u2_u6_n103 ) , .A3( u1_u2_u6_n104 ) , .A2( u1_u2_u6_n105 ) , .A1( u1_u2_u6_n106 ) );
  AOI22_X1 u1_u2_u6_U77 (.ZN( u1_u2_u6_n105 ) , .A2( u1_u2_u6_n108 ) , .A1( u1_u2_u6_n118 ) , .B2( u1_u2_u6_n126 ) , .B1( u1_u2_u6_n171 ) );
  AOI22_X1 u1_u2_u6_U78 (.ZN( u1_u2_u6_n104 ) , .A1( u1_u2_u6_n111 ) , .B1( u1_u2_u6_n124 ) , .B2( u1_u2_u6_n151 ) , .A2( u1_u2_u6_n93 ) );
  NAND4_X1 u1_u2_u6_U79 (.ZN( u1_out2_12 ) , .A4( u1_u2_u6_n114 ) , .A3( u1_u2_u6_n115 ) , .A2( u1_u2_u6_n116 ) , .A1( u1_u2_u6_n117 ) );
  AOI21_X1 u1_u2_u6_U8 (.B1( u1_u2_u6_n107 ) , .B2( u1_u2_u6_n132 ) , .A( u1_u2_u6_n158 ) , .ZN( u1_u2_u6_n88 ) );
  OAI22_X1 u1_u2_u6_U80 (.B2( u1_u2_u6_n111 ) , .ZN( u1_u2_u6_n116 ) , .B1( u1_u2_u6_n126 ) , .A2( u1_u2_u6_n164 ) , .A1( u1_u2_u6_n167 ) );
  OAI21_X1 u1_u2_u6_U81 (.A( u1_u2_u6_n108 ) , .ZN( u1_u2_u6_n117 ) , .B2( u1_u2_u6_n141 ) , .B1( u1_u2_u6_n163 ) );
  OAI211_X1 u1_u2_u6_U82 (.ZN( u1_out2_7 ) , .B( u1_u2_u6_n153 ) , .C2( u1_u2_u6_n154 ) , .C1( u1_u2_u6_n155 ) , .A( u1_u2_u6_n174 ) );
  NOR3_X1 u1_u2_u6_U83 (.A1( u1_u2_u6_n141 ) , .ZN( u1_u2_u6_n154 ) , .A3( u1_u2_u6_n164 ) , .A2( u1_u2_u6_n171 ) );
  AOI211_X1 u1_u2_u6_U84 (.B( u1_u2_u6_n149 ) , .A( u1_u2_u6_n150 ) , .C2( u1_u2_u6_n151 ) , .C1( u1_u2_u6_n152 ) , .ZN( u1_u2_u6_n153 ) );
  OAI211_X1 u1_u2_u6_U85 (.ZN( u1_out2_22 ) , .B( u1_u2_u6_n137 ) , .A( u1_u2_u6_n138 ) , .C2( u1_u2_u6_n139 ) , .C1( u1_u2_u6_n140 ) );
  AOI22_X1 u1_u2_u6_U86 (.B1( u1_u2_u6_n124 ) , .A2( u1_u2_u6_n125 ) , .A1( u1_u2_u6_n126 ) , .ZN( u1_u2_u6_n138 ) , .B2( u1_u2_u6_n161 ) );
  AND4_X1 u1_u2_u6_U87 (.A3( u1_u2_u6_n119 ) , .A1( u1_u2_u6_n120 ) , .A4( u1_u2_u6_n129 ) , .ZN( u1_u2_u6_n140 ) , .A2( u1_u2_u6_n143 ) );
  NAND3_X1 u1_u2_u6_U88 (.A2( u1_u2_u6_n123 ) , .ZN( u1_u2_u6_n125 ) , .A1( u1_u2_u6_n130 ) , .A3( u1_u2_u6_n131 ) );
  NAND3_X1 u1_u2_u6_U89 (.A3( u1_u2_u6_n133 ) , .ZN( u1_u2_u6_n141 ) , .A1( u1_u2_u6_n145 ) , .A2( u1_u2_u6_n148 ) );
  AOI21_X1 u1_u2_u6_U9 (.B2( u1_u2_u6_n147 ) , .B1( u1_u2_u6_n148 ) , .ZN( u1_u2_u6_n149 ) , .A( u1_u2_u6_n158 ) );
  NAND3_X1 u1_u2_u6_U90 (.ZN( u1_u2_u6_n101 ) , .A3( u1_u2_u6_n107 ) , .A2( u1_u2_u6_n121 ) , .A1( u1_u2_u6_n127 ) );
  NAND3_X1 u1_u2_u6_U91 (.ZN( u1_u2_u6_n102 ) , .A3( u1_u2_u6_n130 ) , .A2( u1_u2_u6_n145 ) , .A1( u1_u2_u6_n166 ) );
  NAND3_X1 u1_u2_u6_U92 (.A3( u1_u2_u6_n113 ) , .A1( u1_u2_u6_n119 ) , .A2( u1_u2_u6_n123 ) , .ZN( u1_u2_u6_n93 ) );
  NAND3_X1 u1_u2_u6_U93 (.ZN( u1_u2_u6_n142 ) , .A2( u1_u2_u6_n172 ) , .A3( u1_u2_u6_n89 ) , .A1( u1_u2_u6_n90 ) );
  AND3_X1 u1_u2_u7_U10 (.A3( u1_u2_u7_n110 ) , .A2( u1_u2_u7_n127 ) , .A1( u1_u2_u7_n132 ) , .ZN( u1_u2_u7_n92 ) );
  OAI21_X1 u1_u2_u7_U11 (.A( u1_u2_u7_n161 ) , .B1( u1_u2_u7_n168 ) , .B2( u1_u2_u7_n173 ) , .ZN( u1_u2_u7_n91 ) );
  AOI211_X1 u1_u2_u7_U12 (.A( u1_u2_u7_n117 ) , .ZN( u1_u2_u7_n118 ) , .C2( u1_u2_u7_n126 ) , .C1( u1_u2_u7_n177 ) , .B( u1_u2_u7_n180 ) );
  OAI22_X1 u1_u2_u7_U13 (.B1( u1_u2_u7_n115 ) , .ZN( u1_u2_u7_n117 ) , .A2( u1_u2_u7_n133 ) , .A1( u1_u2_u7_n137 ) , .B2( u1_u2_u7_n162 ) );
  INV_X1 u1_u2_u7_U14 (.A( u1_u2_u7_n116 ) , .ZN( u1_u2_u7_n180 ) );
  NOR3_X1 u1_u2_u7_U15 (.ZN( u1_u2_u7_n115 ) , .A3( u1_u2_u7_n145 ) , .A2( u1_u2_u7_n168 ) , .A1( u1_u2_u7_n169 ) );
  OAI211_X1 u1_u2_u7_U16 (.B( u1_u2_u7_n122 ) , .A( u1_u2_u7_n123 ) , .C2( u1_u2_u7_n124 ) , .ZN( u1_u2_u7_n154 ) , .C1( u1_u2_u7_n162 ) );
  AOI222_X1 u1_u2_u7_U17 (.ZN( u1_u2_u7_n122 ) , .C2( u1_u2_u7_n126 ) , .C1( u1_u2_u7_n145 ) , .B1( u1_u2_u7_n161 ) , .A2( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n170 ) , .A1( u1_u2_u7_n176 ) );
  INV_X1 u1_u2_u7_U18 (.A( u1_u2_u7_n133 ) , .ZN( u1_u2_u7_n176 ) );
  NOR3_X1 u1_u2_u7_U19 (.A2( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n135 ) , .ZN( u1_u2_u7_n136 ) , .A3( u1_u2_u7_n171 ) );
  NOR2_X1 u1_u2_u7_U20 (.A1( u1_u2_u7_n130 ) , .A2( u1_u2_u7_n134 ) , .ZN( u1_u2_u7_n153 ) );
  INV_X1 u1_u2_u7_U21 (.A( u1_u2_u7_n101 ) , .ZN( u1_u2_u7_n165 ) );
  NOR2_X1 u1_u2_u7_U22 (.ZN( u1_u2_u7_n111 ) , .A2( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n169 ) );
  AOI21_X1 u1_u2_u7_U23 (.ZN( u1_u2_u7_n104 ) , .B2( u1_u2_u7_n112 ) , .B1( u1_u2_u7_n127 ) , .A( u1_u2_u7_n164 ) );
  AOI21_X1 u1_u2_u7_U24 (.ZN( u1_u2_u7_n106 ) , .B1( u1_u2_u7_n133 ) , .B2( u1_u2_u7_n146 ) , .A( u1_u2_u7_n162 ) );
  AOI21_X1 u1_u2_u7_U25 (.A( u1_u2_u7_n101 ) , .ZN( u1_u2_u7_n107 ) , .B2( u1_u2_u7_n128 ) , .B1( u1_u2_u7_n175 ) );
  INV_X1 u1_u2_u7_U26 (.A( u1_u2_u7_n138 ) , .ZN( u1_u2_u7_n171 ) );
  INV_X1 u1_u2_u7_U27 (.A( u1_u2_u7_n131 ) , .ZN( u1_u2_u7_n177 ) );
  INV_X1 u1_u2_u7_U28 (.A( u1_u2_u7_n110 ) , .ZN( u1_u2_u7_n174 ) );
  NAND2_X1 u1_u2_u7_U29 (.A1( u1_u2_u7_n129 ) , .A2( u1_u2_u7_n132 ) , .ZN( u1_u2_u7_n149 ) );
  OAI21_X1 u1_u2_u7_U3 (.ZN( u1_u2_u7_n159 ) , .A( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n171 ) , .B1( u1_u2_u7_n174 ) );
  NAND2_X1 u1_u2_u7_U30 (.A1( u1_u2_u7_n113 ) , .A2( u1_u2_u7_n124 ) , .ZN( u1_u2_u7_n130 ) );
  INV_X1 u1_u2_u7_U31 (.A( u1_u2_u7_n112 ) , .ZN( u1_u2_u7_n173 ) );
  INV_X1 u1_u2_u7_U32 (.A( u1_u2_u7_n128 ) , .ZN( u1_u2_u7_n168 ) );
  INV_X1 u1_u2_u7_U33 (.A( u1_u2_u7_n148 ) , .ZN( u1_u2_u7_n169 ) );
  INV_X1 u1_u2_u7_U34 (.A( u1_u2_u7_n127 ) , .ZN( u1_u2_u7_n179 ) );
  NOR2_X1 u1_u2_u7_U35 (.ZN( u1_u2_u7_n101 ) , .A2( u1_u2_u7_n150 ) , .A1( u1_u2_u7_n156 ) );
  AOI211_X1 u1_u2_u7_U36 (.B( u1_u2_u7_n154 ) , .A( u1_u2_u7_n155 ) , .C1( u1_u2_u7_n156 ) , .ZN( u1_u2_u7_n157 ) , .C2( u1_u2_u7_n172 ) );
  INV_X1 u1_u2_u7_U37 (.A( u1_u2_u7_n153 ) , .ZN( u1_u2_u7_n172 ) );
  AOI211_X1 u1_u2_u7_U38 (.B( u1_u2_u7_n139 ) , .A( u1_u2_u7_n140 ) , .C2( u1_u2_u7_n141 ) , .ZN( u1_u2_u7_n142 ) , .C1( u1_u2_u7_n156 ) );
  NAND4_X1 u1_u2_u7_U39 (.A3( u1_u2_u7_n127 ) , .A2( u1_u2_u7_n128 ) , .A1( u1_u2_u7_n129 ) , .ZN( u1_u2_u7_n141 ) , .A4( u1_u2_u7_n147 ) );
  INV_X1 u1_u2_u7_U4 (.A( u1_u2_u7_n111 ) , .ZN( u1_u2_u7_n170 ) );
  AOI21_X1 u1_u2_u7_U40 (.A( u1_u2_u7_n137 ) , .B1( u1_u2_u7_n138 ) , .ZN( u1_u2_u7_n139 ) , .B2( u1_u2_u7_n146 ) );
  OAI22_X1 u1_u2_u7_U41 (.B1( u1_u2_u7_n136 ) , .ZN( u1_u2_u7_n140 ) , .A1( u1_u2_u7_n153 ) , .B2( u1_u2_u7_n162 ) , .A2( u1_u2_u7_n164 ) );
  AOI21_X1 u1_u2_u7_U42 (.ZN( u1_u2_u7_n123 ) , .B1( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n177 ) , .A( u1_u2_u7_n97 ) );
  AOI21_X1 u1_u2_u7_U43 (.B2( u1_u2_u7_n113 ) , .B1( u1_u2_u7_n124 ) , .A( u1_u2_u7_n125 ) , .ZN( u1_u2_u7_n97 ) );
  INV_X1 u1_u2_u7_U44 (.A( u1_u2_u7_n125 ) , .ZN( u1_u2_u7_n161 ) );
  INV_X1 u1_u2_u7_U45 (.A( u1_u2_u7_n152 ) , .ZN( u1_u2_u7_n162 ) );
  AOI22_X1 u1_u2_u7_U46 (.A2( u1_u2_u7_n114 ) , .ZN( u1_u2_u7_n119 ) , .B1( u1_u2_u7_n130 ) , .A1( u1_u2_u7_n156 ) , .B2( u1_u2_u7_n165 ) );
  NAND2_X1 u1_u2_u7_U47 (.A2( u1_u2_u7_n112 ) , .ZN( u1_u2_u7_n114 ) , .A1( u1_u2_u7_n175 ) );
  AND2_X1 u1_u2_u7_U48 (.ZN( u1_u2_u7_n145 ) , .A2( u1_u2_u7_n98 ) , .A1( u1_u2_u7_n99 ) );
  NOR2_X1 u1_u2_u7_U49 (.ZN( u1_u2_u7_n137 ) , .A1( u1_u2_u7_n150 ) , .A2( u1_u2_u7_n161 ) );
  INV_X1 u1_u2_u7_U5 (.A( u1_u2_u7_n149 ) , .ZN( u1_u2_u7_n175 ) );
  AOI21_X1 u1_u2_u7_U50 (.ZN( u1_u2_u7_n105 ) , .B2( u1_u2_u7_n110 ) , .A( u1_u2_u7_n125 ) , .B1( u1_u2_u7_n147 ) );
  NAND2_X1 u1_u2_u7_U51 (.ZN( u1_u2_u7_n146 ) , .A1( u1_u2_u7_n95 ) , .A2( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U52 (.A2( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n147 ) , .A1( u1_u2_u7_n93 ) );
  NAND2_X1 u1_u2_u7_U53 (.A1( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n127 ) , .A2( u1_u2_u7_n99 ) );
  OR2_X1 u1_u2_u7_U54 (.ZN( u1_u2_u7_n126 ) , .A2( u1_u2_u7_n152 ) , .A1( u1_u2_u7_n156 ) );
  NAND2_X1 u1_u2_u7_U55 (.A2( u1_u2_u7_n102 ) , .A1( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n133 ) );
  NAND2_X1 u1_u2_u7_U56 (.ZN( u1_u2_u7_n112 ) , .A2( u1_u2_u7_n96 ) , .A1( u1_u2_u7_n99 ) );
  NAND2_X1 u1_u2_u7_U57 (.A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n128 ) , .A1( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U58 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n113 ) , .A2( u1_u2_u7_n93 ) );
  NAND2_X1 u1_u2_u7_U59 (.A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n124 ) , .A1( u1_u2_u7_n96 ) );
  INV_X1 u1_u2_u7_U6 (.A( u1_u2_u7_n154 ) , .ZN( u1_u2_u7_n178 ) );
  NAND2_X1 u1_u2_u7_U60 (.ZN( u1_u2_u7_n110 ) , .A1( u1_u2_u7_n95 ) , .A2( u1_u2_u7_n96 ) );
  INV_X1 u1_u2_u7_U61 (.A( u1_u2_u7_n150 ) , .ZN( u1_u2_u7_n164 ) );
  AND2_X1 u1_u2_u7_U62 (.ZN( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n93 ) , .A2( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U63 (.A1( u1_u2_u7_n100 ) , .A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n129 ) );
  NAND2_X1 u1_u2_u7_U64 (.A2( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n131 ) , .A1( u1_u2_u7_n95 ) );
  NAND2_X1 u1_u2_u7_U65 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n138 ) , .A2( u1_u2_u7_n99 ) );
  NAND2_X1 u1_u2_u7_U66 (.ZN( u1_u2_u7_n132 ) , .A1( u1_u2_u7_n93 ) , .A2( u1_u2_u7_n96 ) );
  NAND2_X1 u1_u2_u7_U67 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n148 ) , .A2( u1_u2_u7_n95 ) );
  NOR2_X1 u1_u2_u7_U68 (.A2( u1_u2_X_47 ) , .ZN( u1_u2_u7_n150 ) , .A1( u1_u2_u7_n163 ) );
  NOR2_X1 u1_u2_u7_U69 (.A2( u1_u2_X_43 ) , .A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n103 ) );
  AOI211_X1 u1_u2_u7_U7 (.ZN( u1_u2_u7_n116 ) , .A( u1_u2_u7_n155 ) , .C1( u1_u2_u7_n161 ) , .C2( u1_u2_u7_n171 ) , .B( u1_u2_u7_n94 ) );
  NOR2_X1 u1_u2_u7_U70 (.A2( u1_u2_X_48 ) , .A1( u1_u2_u7_n166 ) , .ZN( u1_u2_u7_n95 ) );
  NOR2_X1 u1_u2_u7_U71 (.A2( u1_u2_X_45 ) , .A1( u1_u2_X_48 ) , .ZN( u1_u2_u7_n99 ) );
  NOR2_X1 u1_u2_u7_U72 (.A2( u1_u2_X_44 ) , .A1( u1_u2_u7_n167 ) , .ZN( u1_u2_u7_n98 ) );
  NOR2_X1 u1_u2_u7_U73 (.A2( u1_u2_X_46 ) , .A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n152 ) );
  AND2_X1 u1_u2_u7_U74 (.A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n156 ) , .A2( u1_u2_u7_n163 ) );
  NAND2_X1 u1_u2_u7_U75 (.A2( u1_u2_X_46 ) , .A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n125 ) );
  AND2_X1 u1_u2_u7_U76 (.A2( u1_u2_X_45 ) , .A1( u1_u2_X_48 ) , .ZN( u1_u2_u7_n102 ) );
  AND2_X1 u1_u2_u7_U77 (.A2( u1_u2_X_43 ) , .A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n96 ) );
  AND2_X1 u1_u2_u7_U78 (.A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n100 ) , .A2( u1_u2_u7_n167 ) );
  AND2_X1 u1_u2_u7_U79 (.A1( u1_u2_X_48 ) , .A2( u1_u2_u7_n166 ) , .ZN( u1_u2_u7_n93 ) );
  OAI222_X1 u1_u2_u7_U8 (.C2( u1_u2_u7_n101 ) , .B2( u1_u2_u7_n111 ) , .A1( u1_u2_u7_n113 ) , .C1( u1_u2_u7_n146 ) , .A2( u1_u2_u7_n162 ) , .B1( u1_u2_u7_n164 ) , .ZN( u1_u2_u7_n94 ) );
  INV_X1 u1_u2_u7_U80 (.A( u1_u2_X_46 ) , .ZN( u1_u2_u7_n163 ) );
  INV_X1 u1_u2_u7_U81 (.A( u1_u2_X_43 ) , .ZN( u1_u2_u7_n167 ) );
  INV_X1 u1_u2_u7_U82 (.A( u1_u2_X_45 ) , .ZN( u1_u2_u7_n166 ) );
  NAND4_X1 u1_u2_u7_U83 (.ZN( u1_out2_5 ) , .A4( u1_u2_u7_n108 ) , .A3( u1_u2_u7_n109 ) , .A1( u1_u2_u7_n116 ) , .A2( u1_u2_u7_n123 ) );
  AOI22_X1 u1_u2_u7_U84 (.ZN( u1_u2_u7_n109 ) , .A2( u1_u2_u7_n126 ) , .B2( u1_u2_u7_n145 ) , .B1( u1_u2_u7_n156 ) , .A1( u1_u2_u7_n171 ) );
  NOR4_X1 u1_u2_u7_U85 (.A4( u1_u2_u7_n104 ) , .A3( u1_u2_u7_n105 ) , .A2( u1_u2_u7_n106 ) , .A1( u1_u2_u7_n107 ) , .ZN( u1_u2_u7_n108 ) );
  NAND4_X1 u1_u2_u7_U86 (.ZN( u1_out2_27 ) , .A4( u1_u2_u7_n118 ) , .A3( u1_u2_u7_n119 ) , .A2( u1_u2_u7_n120 ) , .A1( u1_u2_u7_n121 ) );
  OAI21_X1 u1_u2_u7_U87 (.ZN( u1_u2_u7_n121 ) , .B2( u1_u2_u7_n145 ) , .A( u1_u2_u7_n150 ) , .B1( u1_u2_u7_n174 ) );
  OAI21_X1 u1_u2_u7_U88 (.ZN( u1_u2_u7_n120 ) , .A( u1_u2_u7_n161 ) , .B2( u1_u2_u7_n170 ) , .B1( u1_u2_u7_n179 ) );
  NAND4_X1 u1_u2_u7_U89 (.ZN( u1_out2_21 ) , .A4( u1_u2_u7_n157 ) , .A3( u1_u2_u7_n158 ) , .A2( u1_u2_u7_n159 ) , .A1( u1_u2_u7_n160 ) );
  OAI221_X1 u1_u2_u7_U9 (.C1( u1_u2_u7_n101 ) , .C2( u1_u2_u7_n147 ) , .ZN( u1_u2_u7_n155 ) , .B2( u1_u2_u7_n162 ) , .A( u1_u2_u7_n91 ) , .B1( u1_u2_u7_n92 ) );
  OAI21_X1 u1_u2_u7_U90 (.B1( u1_u2_u7_n145 ) , .ZN( u1_u2_u7_n160 ) , .A( u1_u2_u7_n161 ) , .B2( u1_u2_u7_n177 ) );
  AOI22_X1 u1_u2_u7_U91 (.B2( u1_u2_u7_n149 ) , .B1( u1_u2_u7_n150 ) , .A2( u1_u2_u7_n151 ) , .A1( u1_u2_u7_n152 ) , .ZN( u1_u2_u7_n158 ) );
  NAND4_X1 u1_u2_u7_U92 (.ZN( u1_out2_15 ) , .A4( u1_u2_u7_n142 ) , .A3( u1_u2_u7_n143 ) , .A2( u1_u2_u7_n144 ) , .A1( u1_u2_u7_n178 ) );
  OR2_X1 u1_u2_u7_U93 (.A2( u1_u2_u7_n125 ) , .A1( u1_u2_u7_n129 ) , .ZN( u1_u2_u7_n144 ) );
  AOI22_X1 u1_u2_u7_U94 (.A2( u1_u2_u7_n126 ) , .ZN( u1_u2_u7_n143 ) , .B2( u1_u2_u7_n165 ) , .B1( u1_u2_u7_n173 ) , .A1( u1_u2_u7_n174 ) );
  NAND3_X1 u1_u2_u7_U95 (.A3( u1_u2_u7_n146 ) , .A2( u1_u2_u7_n147 ) , .A1( u1_u2_u7_n148 ) , .ZN( u1_u2_u7_n151 ) );
  NAND3_X1 u1_u2_u7_U96 (.A3( u1_u2_u7_n131 ) , .A2( u1_u2_u7_n132 ) , .A1( u1_u2_u7_n133 ) , .ZN( u1_u2_u7_n135 ) );
  XOR2_X1 u1_u3_U16 (.B( u1_K4_3 ) , .A( u1_R2_2 ) , .Z( u1_u3_X_3 ) );
  XOR2_X1 u1_u3_U2 (.B( u1_K4_8 ) , .A( u1_R2_5 ) , .Z( u1_u3_X_8 ) );
  XOR2_X1 u1_u3_U27 (.B( u1_K4_2 ) , .A( u1_R2_1 ) , .Z( u1_u3_X_2 ) );
  XOR2_X1 u1_u3_U38 (.B( u1_K4_1 ) , .A( u1_R2_32 ) , .Z( u1_u3_X_1 ) );
  XOR2_X1 u1_u3_U4 (.B( u1_K4_6 ) , .A( u1_R2_5 ) , .Z( u1_u3_X_6 ) );
  XOR2_X1 u1_u3_U46 (.B( u1_K4_12 ) , .A( u1_R2_9 ) , .Z( u1_u3_X_12 ) );
  XOR2_X1 u1_u3_U47 (.B( u1_K4_11 ) , .A( u1_R2_8 ) , .Z( u1_u3_X_11 ) );
  XOR2_X1 u1_u3_U48 (.B( u1_K4_10 ) , .A( u1_R2_7 ) , .Z( u1_u3_X_10 ) );
  AND2_X1 u1_u3_u0_U10 (.A1( u1_u3_u0_n131 ) , .ZN( u1_u3_u0_n141 ) , .A2( u1_u3_u0_n150 ) );
  AND3_X1 u1_u3_u0_U11 (.A2( u1_u3_u0_n112 ) , .ZN( u1_u3_u0_n127 ) , .A3( u1_u3_u0_n130 ) , .A1( u1_u3_u0_n148 ) );
  AND2_X1 u1_u3_u0_U12 (.ZN( u1_u3_u0_n107 ) , .A1( u1_u3_u0_n130 ) , .A2( u1_u3_u0_n140 ) );
  AND2_X1 u1_u3_u0_U13 (.A2( u1_u3_u0_n129 ) , .A1( u1_u3_u0_n130 ) , .ZN( u1_u3_u0_n151 ) );
  AND2_X1 u1_u3_u0_U14 (.A1( u1_u3_u0_n108 ) , .A2( u1_u3_u0_n125 ) , .ZN( u1_u3_u0_n145 ) );
  INV_X1 u1_u3_u0_U15 (.A( u1_u3_u0_n143 ) , .ZN( u1_u3_u0_n173 ) );
  NOR2_X1 u1_u3_u0_U16 (.A2( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n147 ) , .A1( u1_u3_u0_n160 ) );
  AOI21_X1 u1_u3_u0_U17 (.B1( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n132 ) , .A( u1_u3_u0_n165 ) , .B2( u1_u3_u0_n93 ) );
  OAI22_X1 u1_u3_u0_U18 (.B1( u1_u3_u0_n131 ) , .A1( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n147 ) , .A2( u1_u3_u0_n90 ) , .ZN( u1_u3_u0_n91 ) );
  AND3_X1 u1_u3_u0_U19 (.A3( u1_u3_u0_n121 ) , .A2( u1_u3_u0_n125 ) , .A1( u1_u3_u0_n148 ) , .ZN( u1_u3_u0_n90 ) );
  OAI22_X1 u1_u3_u0_U20 (.B1( u1_u3_u0_n125 ) , .ZN( u1_u3_u0_n126 ) , .A1( u1_u3_u0_n138 ) , .A2( u1_u3_u0_n146 ) , .B2( u1_u3_u0_n147 ) );
  NOR2_X1 u1_u3_u0_U21 (.A1( u1_u3_u0_n163 ) , .A2( u1_u3_u0_n164 ) , .ZN( u1_u3_u0_n95 ) );
  AOI22_X1 u1_u3_u0_U22 (.B2( u1_u3_u0_n109 ) , .A2( u1_u3_u0_n110 ) , .ZN( u1_u3_u0_n111 ) , .B1( u1_u3_u0_n118 ) , .A1( u1_u3_u0_n160 ) );
  NAND2_X1 u1_u3_u0_U23 (.A2( u1_u3_u0_n102 ) , .A1( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n149 ) );
  INV_X1 u1_u3_u0_U24 (.A( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n161 ) );
  INV_X1 u1_u3_u0_U25 (.A( u1_u3_u0_n118 ) , .ZN( u1_u3_u0_n158 ) );
  NAND2_X1 u1_u3_u0_U26 (.A2( u1_u3_u0_n100 ) , .ZN( u1_u3_u0_n131 ) , .A1( u1_u3_u0_n92 ) );
  NAND2_X1 u1_u3_u0_U27 (.ZN( u1_u3_u0_n108 ) , .A1( u1_u3_u0_n92 ) , .A2( u1_u3_u0_n94 ) );
  AOI21_X1 u1_u3_u0_U28 (.ZN( u1_u3_u0_n104 ) , .B1( u1_u3_u0_n107 ) , .B2( u1_u3_u0_n141 ) , .A( u1_u3_u0_n144 ) );
  AOI21_X1 u1_u3_u0_U29 (.B1( u1_u3_u0_n127 ) , .B2( u1_u3_u0_n129 ) , .A( u1_u3_u0_n138 ) , .ZN( u1_u3_u0_n96 ) );
  INV_X1 u1_u3_u0_U3 (.A( u1_u3_u0_n113 ) , .ZN( u1_u3_u0_n166 ) );
  NAND2_X1 u1_u3_u0_U30 (.A2( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n114 ) , .A1( u1_u3_u0_n92 ) );
  NOR2_X1 u1_u3_u0_U31 (.A1( u1_u3_u0_n120 ) , .ZN( u1_u3_u0_n143 ) , .A2( u1_u3_u0_n167 ) );
  OAI221_X1 u1_u3_u0_U32 (.C1( u1_u3_u0_n112 ) , .ZN( u1_u3_u0_n120 ) , .B1( u1_u3_u0_n138 ) , .B2( u1_u3_u0_n141 ) , .C2( u1_u3_u0_n147 ) , .A( u1_u3_u0_n172 ) );
  AOI211_X1 u1_u3_u0_U33 (.B( u1_u3_u0_n115 ) , .A( u1_u3_u0_n116 ) , .C2( u1_u3_u0_n117 ) , .C1( u1_u3_u0_n118 ) , .ZN( u1_u3_u0_n119 ) );
  NAND2_X1 u1_u3_u0_U34 (.A2( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n140 ) , .A1( u1_u3_u0_n94 ) );
  NAND2_X1 u1_u3_u0_U35 (.A1( u1_u3_u0_n100 ) , .A2( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n125 ) );
  NAND2_X1 u1_u3_u0_U36 (.A1( u1_u3_u0_n101 ) , .A2( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n150 ) );
  INV_X1 u1_u3_u0_U37 (.A( u1_u3_u0_n138 ) , .ZN( u1_u3_u0_n160 ) );
  NAND2_X1 u1_u3_u0_U38 (.A2( u1_u3_u0_n100 ) , .A1( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n139 ) );
  NAND2_X1 u1_u3_u0_U39 (.ZN( u1_u3_u0_n112 ) , .A2( u1_u3_u0_n92 ) , .A1( u1_u3_u0_n93 ) );
  AOI21_X1 u1_u3_u0_U4 (.B1( u1_u3_u0_n114 ) , .ZN( u1_u3_u0_n115 ) , .B2( u1_u3_u0_n129 ) , .A( u1_u3_u0_n161 ) );
  NAND2_X1 u1_u3_u0_U40 (.A1( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n130 ) , .A2( u1_u3_u0_n94 ) );
  INV_X1 u1_u3_u0_U41 (.ZN( u1_u3_u0_n172 ) , .A( u1_u3_u0_n88 ) );
  OAI222_X1 u1_u3_u0_U42 (.C1( u1_u3_u0_n108 ) , .A1( u1_u3_u0_n125 ) , .B2( u1_u3_u0_n128 ) , .B1( u1_u3_u0_n144 ) , .A2( u1_u3_u0_n158 ) , .C2( u1_u3_u0_n161 ) , .ZN( u1_u3_u0_n88 ) );
  NAND2_X1 u1_u3_u0_U43 (.A2( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n121 ) , .A1( u1_u3_u0_n93 ) );
  OR3_X1 u1_u3_u0_U44 (.A3( u1_u3_u0_n152 ) , .A2( u1_u3_u0_n153 ) , .A1( u1_u3_u0_n154 ) , .ZN( u1_u3_u0_n155 ) );
  AOI21_X1 u1_u3_u0_U45 (.A( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n145 ) , .B1( u1_u3_u0_n146 ) , .ZN( u1_u3_u0_n154 ) );
  AOI21_X1 u1_u3_u0_U46 (.B2( u1_u3_u0_n150 ) , .B1( u1_u3_u0_n151 ) , .ZN( u1_u3_u0_n152 ) , .A( u1_u3_u0_n158 ) );
  AOI21_X1 u1_u3_u0_U47 (.A( u1_u3_u0_n147 ) , .B2( u1_u3_u0_n148 ) , .B1( u1_u3_u0_n149 ) , .ZN( u1_u3_u0_n153 ) );
  INV_X1 u1_u3_u0_U48 (.ZN( u1_u3_u0_n171 ) , .A( u1_u3_u0_n99 ) );
  OAI211_X1 u1_u3_u0_U49 (.C2( u1_u3_u0_n140 ) , .C1( u1_u3_u0_n161 ) , .A( u1_u3_u0_n169 ) , .B( u1_u3_u0_n98 ) , .ZN( u1_u3_u0_n99 ) );
  AOI21_X1 u1_u3_u0_U5 (.B2( u1_u3_u0_n131 ) , .ZN( u1_u3_u0_n134 ) , .B1( u1_u3_u0_n151 ) , .A( u1_u3_u0_n158 ) );
  AOI211_X1 u1_u3_u0_U50 (.C1( u1_u3_u0_n118 ) , .A( u1_u3_u0_n123 ) , .B( u1_u3_u0_n96 ) , .C2( u1_u3_u0_n97 ) , .ZN( u1_u3_u0_n98 ) );
  INV_X1 u1_u3_u0_U51 (.ZN( u1_u3_u0_n169 ) , .A( u1_u3_u0_n91 ) );
  NOR2_X1 u1_u3_u0_U52 (.A2( u1_u3_X_4 ) , .A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n118 ) );
  NOR2_X1 u1_u3_u0_U53 (.A2( u1_u3_X_1 ) , .ZN( u1_u3_u0_n101 ) , .A1( u1_u3_u0_n163 ) );
  NOR2_X1 u1_u3_u0_U54 (.A2( u1_u3_X_3 ) , .A1( u1_u3_X_6 ) , .ZN( u1_u3_u0_n94 ) );
  NOR2_X1 u1_u3_u0_U55 (.A2( u1_u3_X_6 ) , .ZN( u1_u3_u0_n100 ) , .A1( u1_u3_u0_n162 ) );
  NAND2_X1 u1_u3_u0_U56 (.A2( u1_u3_X_4 ) , .A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n144 ) );
  NOR2_X1 u1_u3_u0_U57 (.A2( u1_u3_X_5 ) , .ZN( u1_u3_u0_n136 ) , .A1( u1_u3_u0_n159 ) );
  NAND2_X1 u1_u3_u0_U58 (.A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n138 ) , .A2( u1_u3_u0_n159 ) );
  AND2_X1 u1_u3_u0_U59 (.A2( u1_u3_X_3 ) , .A1( u1_u3_X_6 ) , .ZN( u1_u3_u0_n102 ) );
  NOR2_X1 u1_u3_u0_U6 (.A1( u1_u3_u0_n108 ) , .ZN( u1_u3_u0_n123 ) , .A2( u1_u3_u0_n158 ) );
  AND2_X1 u1_u3_u0_U60 (.A1( u1_u3_X_6 ) , .A2( u1_u3_u0_n162 ) , .ZN( u1_u3_u0_n93 ) );
  INV_X1 u1_u3_u0_U61 (.A( u1_u3_X_4 ) , .ZN( u1_u3_u0_n159 ) );
  INV_X1 u1_u3_u0_U62 (.A( u1_u3_X_1 ) , .ZN( u1_u3_u0_n164 ) );
  INV_X1 u1_u3_u0_U63 (.A( u1_u3_X_3 ) , .ZN( u1_u3_u0_n162 ) );
  INV_X1 u1_u3_u0_U64 (.A( u1_u3_u0_n126 ) , .ZN( u1_u3_u0_n168 ) );
  AOI211_X1 u1_u3_u0_U65 (.B( u1_u3_u0_n133 ) , .A( u1_u3_u0_n134 ) , .C2( u1_u3_u0_n135 ) , .C1( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n137 ) );
  OR4_X1 u1_u3_u0_U66 (.ZN( u1_out3_17 ) , .A4( u1_u3_u0_n122 ) , .A2( u1_u3_u0_n123 ) , .A1( u1_u3_u0_n124 ) , .A3( u1_u3_u0_n170 ) );
  AOI21_X1 u1_u3_u0_U67 (.B2( u1_u3_u0_n107 ) , .ZN( u1_u3_u0_n124 ) , .B1( u1_u3_u0_n128 ) , .A( u1_u3_u0_n161 ) );
  INV_X1 u1_u3_u0_U68 (.A( u1_u3_u0_n111 ) , .ZN( u1_u3_u0_n170 ) );
  OR4_X1 u1_u3_u0_U69 (.ZN( u1_out3_31 ) , .A4( u1_u3_u0_n155 ) , .A2( u1_u3_u0_n156 ) , .A1( u1_u3_u0_n157 ) , .A3( u1_u3_u0_n173 ) );
  OAI21_X1 u1_u3_u0_U7 (.B1( u1_u3_u0_n150 ) , .B2( u1_u3_u0_n158 ) , .A( u1_u3_u0_n172 ) , .ZN( u1_u3_u0_n89 ) );
  AOI21_X1 u1_u3_u0_U70 (.A( u1_u3_u0_n138 ) , .B2( u1_u3_u0_n139 ) , .B1( u1_u3_u0_n140 ) , .ZN( u1_u3_u0_n157 ) );
  INV_X1 u1_u3_u0_U71 (.ZN( u1_u3_u0_n174 ) , .A( u1_u3_u0_n89 ) );
  AOI211_X1 u1_u3_u0_U72 (.B( u1_u3_u0_n104 ) , .A( u1_u3_u0_n105 ) , .ZN( u1_u3_u0_n106 ) , .C2( u1_u3_u0_n113 ) , .C1( u1_u3_u0_n160 ) );
  AOI21_X1 u1_u3_u0_U73 (.B2( u1_u3_u0_n141 ) , .B1( u1_u3_u0_n142 ) , .ZN( u1_u3_u0_n156 ) , .A( u1_u3_u0_n161 ) );
  AOI21_X1 u1_u3_u0_U74 (.ZN( u1_u3_u0_n116 ) , .B2( u1_u3_u0_n142 ) , .A( u1_u3_u0_n144 ) , .B1( u1_u3_u0_n166 ) );
  INV_X1 u1_u3_u0_U75 (.A( u1_u3_u0_n142 ) , .ZN( u1_u3_u0_n165 ) );
  NOR2_X1 u1_u3_u0_U76 (.A2( u1_u3_X_1 ) , .A1( u1_u3_X_2 ) , .ZN( u1_u3_u0_n92 ) );
  NOR2_X1 u1_u3_u0_U77 (.A2( u1_u3_X_2 ) , .ZN( u1_u3_u0_n103 ) , .A1( u1_u3_u0_n164 ) );
  INV_X1 u1_u3_u0_U78 (.A( u1_u3_X_2 ) , .ZN( u1_u3_u0_n163 ) );
  OAI221_X1 u1_u3_u0_U79 (.C1( u1_u3_u0_n121 ) , .ZN( u1_u3_u0_n122 ) , .B2( u1_u3_u0_n127 ) , .A( u1_u3_u0_n143 ) , .B1( u1_u3_u0_n144 ) , .C2( u1_u3_u0_n147 ) );
  AND2_X1 u1_u3_u0_U8 (.A1( u1_u3_u0_n114 ) , .A2( u1_u3_u0_n121 ) , .ZN( u1_u3_u0_n146 ) );
  AOI21_X1 u1_u3_u0_U80 (.B1( u1_u3_u0_n132 ) , .ZN( u1_u3_u0_n133 ) , .A( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n166 ) );
  OAI22_X1 u1_u3_u0_U81 (.ZN( u1_u3_u0_n105 ) , .A2( u1_u3_u0_n132 ) , .B1( u1_u3_u0_n146 ) , .A1( u1_u3_u0_n147 ) , .B2( u1_u3_u0_n161 ) );
  NAND2_X1 u1_u3_u0_U82 (.ZN( u1_u3_u0_n110 ) , .A2( u1_u3_u0_n132 ) , .A1( u1_u3_u0_n145 ) );
  INV_X1 u1_u3_u0_U83 (.A( u1_u3_u0_n119 ) , .ZN( u1_u3_u0_n167 ) );
  NAND2_X1 u1_u3_u0_U84 (.ZN( u1_u3_u0_n148 ) , .A1( u1_u3_u0_n93 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U85 (.A1( u1_u3_u0_n100 ) , .ZN( u1_u3_u0_n129 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U86 (.A1( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n128 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U87 (.ZN( u1_u3_u0_n142 ) , .A1( u1_u3_u0_n94 ) , .A2( u1_u3_u0_n95 ) );
  NAND3_X1 u1_u3_u0_U88 (.ZN( u1_out3_23 ) , .A3( u1_u3_u0_n137 ) , .A1( u1_u3_u0_n168 ) , .A2( u1_u3_u0_n171 ) );
  NAND3_X1 u1_u3_u0_U89 (.A3( u1_u3_u0_n127 ) , .A2( u1_u3_u0_n128 ) , .ZN( u1_u3_u0_n135 ) , .A1( u1_u3_u0_n150 ) );
  NAND2_X1 u1_u3_u0_U9 (.ZN( u1_u3_u0_n113 ) , .A1( u1_u3_u0_n139 ) , .A2( u1_u3_u0_n149 ) );
  NAND3_X1 u1_u3_u0_U90 (.ZN( u1_u3_u0_n117 ) , .A3( u1_u3_u0_n132 ) , .A2( u1_u3_u0_n139 ) , .A1( u1_u3_u0_n148 ) );
  NAND3_X1 u1_u3_u0_U91 (.ZN( u1_u3_u0_n109 ) , .A2( u1_u3_u0_n114 ) , .A3( u1_u3_u0_n140 ) , .A1( u1_u3_u0_n149 ) );
  NAND3_X1 u1_u3_u0_U92 (.ZN( u1_out3_9 ) , .A3( u1_u3_u0_n106 ) , .A2( u1_u3_u0_n171 ) , .A1( u1_u3_u0_n174 ) );
  NAND3_X1 u1_u3_u0_U93 (.A2( u1_u3_u0_n128 ) , .A1( u1_u3_u0_n132 ) , .A3( u1_u3_u0_n146 ) , .ZN( u1_u3_u0_n97 ) );
  AOI21_X1 u1_u3_u1_U10 (.B2( u1_u3_u1_n155 ) , .B1( u1_u3_u1_n156 ) , .ZN( u1_u3_u1_n157 ) , .A( u1_u3_u1_n174 ) );
  NAND3_X1 u1_u3_u1_U100 (.ZN( u1_u3_u1_n113 ) , .A1( u1_u3_u1_n120 ) , .A3( u1_u3_u1_n133 ) , .A2( u1_u3_u1_n155 ) );
  NAND2_X1 u1_u3_u1_U11 (.ZN( u1_u3_u1_n140 ) , .A2( u1_u3_u1_n150 ) , .A1( u1_u3_u1_n155 ) );
  NAND2_X1 u1_u3_u1_U12 (.A1( u1_u3_u1_n131 ) , .ZN( u1_u3_u1_n147 ) , .A2( u1_u3_u1_n153 ) );
  INV_X1 u1_u3_u1_U13 (.A( u1_u3_u1_n139 ) , .ZN( u1_u3_u1_n174 ) );
  OR4_X1 u1_u3_u1_U14 (.A4( u1_u3_u1_n106 ) , .A3( u1_u3_u1_n107 ) , .ZN( u1_u3_u1_n108 ) , .A1( u1_u3_u1_n117 ) , .A2( u1_u3_u1_n184 ) );
  AOI21_X1 u1_u3_u1_U15 (.ZN( u1_u3_u1_n106 ) , .A( u1_u3_u1_n112 ) , .B1( u1_u3_u1_n154 ) , .B2( u1_u3_u1_n156 ) );
  INV_X1 u1_u3_u1_U16 (.A( u1_u3_u1_n101 ) , .ZN( u1_u3_u1_n184 ) );
  AOI21_X1 u1_u3_u1_U17 (.ZN( u1_u3_u1_n107 ) , .B1( u1_u3_u1_n134 ) , .B2( u1_u3_u1_n149 ) , .A( u1_u3_u1_n174 ) );
  INV_X1 u1_u3_u1_U18 (.A( u1_u3_u1_n112 ) , .ZN( u1_u3_u1_n171 ) );
  NAND2_X1 u1_u3_u1_U19 (.ZN( u1_u3_u1_n141 ) , .A1( u1_u3_u1_n153 ) , .A2( u1_u3_u1_n156 ) );
  AND2_X1 u1_u3_u1_U20 (.A1( u1_u3_u1_n123 ) , .ZN( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n161 ) );
  NAND2_X1 u1_u3_u1_U21 (.A2( u1_u3_u1_n115 ) , .A1( u1_u3_u1_n116 ) , .ZN( u1_u3_u1_n148 ) );
  NAND2_X1 u1_u3_u1_U22 (.A2( u1_u3_u1_n133 ) , .A1( u1_u3_u1_n135 ) , .ZN( u1_u3_u1_n159 ) );
  NAND2_X1 u1_u3_u1_U23 (.A2( u1_u3_u1_n115 ) , .A1( u1_u3_u1_n120 ) , .ZN( u1_u3_u1_n132 ) );
  INV_X1 u1_u3_u1_U24 (.A( u1_u3_u1_n154 ) , .ZN( u1_u3_u1_n178 ) );
  AOI22_X1 u1_u3_u1_U25 (.B2( u1_u3_u1_n113 ) , .A2( u1_u3_u1_n114 ) , .ZN( u1_u3_u1_n125 ) , .A1( u1_u3_u1_n171 ) , .B1( u1_u3_u1_n173 ) );
  NAND2_X1 u1_u3_u1_U26 (.ZN( u1_u3_u1_n114 ) , .A1( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n156 ) );
  INV_X1 u1_u3_u1_U27 (.A( u1_u3_u1_n151 ) , .ZN( u1_u3_u1_n183 ) );
  AND2_X1 u1_u3_u1_U28 (.A1( u1_u3_u1_n129 ) , .A2( u1_u3_u1_n133 ) , .ZN( u1_u3_u1_n149 ) );
  INV_X1 u1_u3_u1_U29 (.A( u1_u3_u1_n131 ) , .ZN( u1_u3_u1_n180 ) );
  INV_X1 u1_u3_u1_U3 (.A( u1_u3_u1_n159 ) , .ZN( u1_u3_u1_n182 ) );
  AOI221_X1 u1_u3_u1_U30 (.B1( u1_u3_u1_n140 ) , .ZN( u1_u3_u1_n167 ) , .B2( u1_u3_u1_n172 ) , .C2( u1_u3_u1_n175 ) , .C1( u1_u3_u1_n178 ) , .A( u1_u3_u1_n188 ) );
  INV_X1 u1_u3_u1_U31 (.ZN( u1_u3_u1_n188 ) , .A( u1_u3_u1_n97 ) );
  AOI211_X1 u1_u3_u1_U32 (.A( u1_u3_u1_n118 ) , .C1( u1_u3_u1_n132 ) , .C2( u1_u3_u1_n139 ) , .B( u1_u3_u1_n96 ) , .ZN( u1_u3_u1_n97 ) );
  AOI21_X1 u1_u3_u1_U33 (.B2( u1_u3_u1_n121 ) , .B1( u1_u3_u1_n135 ) , .A( u1_u3_u1_n152 ) , .ZN( u1_u3_u1_n96 ) );
  OAI221_X1 u1_u3_u1_U34 (.A( u1_u3_u1_n119 ) , .C2( u1_u3_u1_n129 ) , .ZN( u1_u3_u1_n138 ) , .B2( u1_u3_u1_n152 ) , .C1( u1_u3_u1_n174 ) , .B1( u1_u3_u1_n187 ) );
  INV_X1 u1_u3_u1_U35 (.A( u1_u3_u1_n148 ) , .ZN( u1_u3_u1_n187 ) );
  AOI211_X1 u1_u3_u1_U36 (.B( u1_u3_u1_n117 ) , .A( u1_u3_u1_n118 ) , .ZN( u1_u3_u1_n119 ) , .C2( u1_u3_u1_n146 ) , .C1( u1_u3_u1_n159 ) );
  NOR2_X1 u1_u3_u1_U37 (.A1( u1_u3_u1_n168 ) , .A2( u1_u3_u1_n176 ) , .ZN( u1_u3_u1_n98 ) );
  AOI211_X1 u1_u3_u1_U38 (.B( u1_u3_u1_n162 ) , .A( u1_u3_u1_n163 ) , .C2( u1_u3_u1_n164 ) , .ZN( u1_u3_u1_n165 ) , .C1( u1_u3_u1_n171 ) );
  AOI21_X1 u1_u3_u1_U39 (.A( u1_u3_u1_n160 ) , .B2( u1_u3_u1_n161 ) , .ZN( u1_u3_u1_n162 ) , .B1( u1_u3_u1_n182 ) );
  AOI221_X1 u1_u3_u1_U4 (.A( u1_u3_u1_n138 ) , .C2( u1_u3_u1_n139 ) , .C1( u1_u3_u1_n140 ) , .B2( u1_u3_u1_n141 ) , .ZN( u1_u3_u1_n142 ) , .B1( u1_u3_u1_n175 ) );
  OR2_X1 u1_u3_u1_U40 (.A2( u1_u3_u1_n157 ) , .A1( u1_u3_u1_n158 ) , .ZN( u1_u3_u1_n163 ) );
  NAND2_X1 u1_u3_u1_U41 (.A1( u1_u3_u1_n128 ) , .ZN( u1_u3_u1_n146 ) , .A2( u1_u3_u1_n160 ) );
  NAND2_X1 u1_u3_u1_U42 (.A2( u1_u3_u1_n112 ) , .ZN( u1_u3_u1_n139 ) , .A1( u1_u3_u1_n152 ) );
  NAND2_X1 u1_u3_u1_U43 (.A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n156 ) , .A2( u1_u3_u1_n99 ) );
  NOR2_X1 u1_u3_u1_U44 (.ZN( u1_u3_u1_n117 ) , .A1( u1_u3_u1_n121 ) , .A2( u1_u3_u1_n160 ) );
  OAI21_X1 u1_u3_u1_U45 (.B2( u1_u3_u1_n123 ) , .ZN( u1_u3_u1_n145 ) , .B1( u1_u3_u1_n160 ) , .A( u1_u3_u1_n185 ) );
  INV_X1 u1_u3_u1_U46 (.A( u1_u3_u1_n122 ) , .ZN( u1_u3_u1_n185 ) );
  AOI21_X1 u1_u3_u1_U47 (.B2( u1_u3_u1_n120 ) , .B1( u1_u3_u1_n121 ) , .ZN( u1_u3_u1_n122 ) , .A( u1_u3_u1_n128 ) );
  AOI21_X1 u1_u3_u1_U48 (.A( u1_u3_u1_n128 ) , .B2( u1_u3_u1_n129 ) , .ZN( u1_u3_u1_n130 ) , .B1( u1_u3_u1_n150 ) );
  NAND2_X1 u1_u3_u1_U49 (.ZN( u1_u3_u1_n112 ) , .A1( u1_u3_u1_n169 ) , .A2( u1_u3_u1_n170 ) );
  AOI211_X1 u1_u3_u1_U5 (.ZN( u1_u3_u1_n124 ) , .A( u1_u3_u1_n138 ) , .C2( u1_u3_u1_n139 ) , .B( u1_u3_u1_n145 ) , .C1( u1_u3_u1_n147 ) );
  NAND2_X1 u1_u3_u1_U50 (.ZN( u1_u3_u1_n129 ) , .A2( u1_u3_u1_n95 ) , .A1( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U51 (.A1( u1_u3_u1_n102 ) , .ZN( u1_u3_u1_n154 ) , .A2( u1_u3_u1_n99 ) );
  NAND2_X1 u1_u3_u1_U52 (.A2( u1_u3_u1_n100 ) , .ZN( u1_u3_u1_n135 ) , .A1( u1_u3_u1_n99 ) );
  AOI21_X1 u1_u3_u1_U53 (.A( u1_u3_u1_n152 ) , .B2( u1_u3_u1_n153 ) , .B1( u1_u3_u1_n154 ) , .ZN( u1_u3_u1_n158 ) );
  INV_X1 u1_u3_u1_U54 (.A( u1_u3_u1_n160 ) , .ZN( u1_u3_u1_n175 ) );
  NAND2_X1 u1_u3_u1_U55 (.A1( u1_u3_u1_n100 ) , .ZN( u1_u3_u1_n116 ) , .A2( u1_u3_u1_n95 ) );
  NAND2_X1 u1_u3_u1_U56 (.A1( u1_u3_u1_n102 ) , .ZN( u1_u3_u1_n131 ) , .A2( u1_u3_u1_n95 ) );
  NAND2_X1 u1_u3_u1_U57 (.A2( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n121 ) , .A1( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U58 (.A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n153 ) , .A2( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U59 (.A2( u1_u3_u1_n104 ) , .A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n133 ) );
  AOI22_X1 u1_u3_u1_U6 (.B2( u1_u3_u1_n136 ) , .A2( u1_u3_u1_n137 ) , .ZN( u1_u3_u1_n143 ) , .A1( u1_u3_u1_n171 ) , .B1( u1_u3_u1_n173 ) );
  NAND2_X1 u1_u3_u1_U60 (.ZN( u1_u3_u1_n150 ) , .A2( u1_u3_u1_n98 ) , .A1( u1_u3_u1_n99 ) );
  NAND2_X1 u1_u3_u1_U61 (.A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n155 ) , .A2( u1_u3_u1_n95 ) );
  OAI21_X1 u1_u3_u1_U62 (.ZN( u1_u3_u1_n109 ) , .B1( u1_u3_u1_n129 ) , .B2( u1_u3_u1_n160 ) , .A( u1_u3_u1_n167 ) );
  NAND2_X1 u1_u3_u1_U63 (.A2( u1_u3_u1_n100 ) , .A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n120 ) );
  NAND2_X1 u1_u3_u1_U64 (.A1( u1_u3_u1_n102 ) , .A2( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n115 ) );
  NAND2_X1 u1_u3_u1_U65 (.A2( u1_u3_u1_n100 ) , .A1( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n151 ) );
  NAND2_X1 u1_u3_u1_U66 (.A2( u1_u3_u1_n103 ) , .A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n161 ) );
  INV_X1 u1_u3_u1_U67 (.A( u1_u3_u1_n152 ) , .ZN( u1_u3_u1_n173 ) );
  INV_X1 u1_u3_u1_U68 (.A( u1_u3_u1_n128 ) , .ZN( u1_u3_u1_n172 ) );
  NAND2_X1 u1_u3_u1_U69 (.A2( u1_u3_u1_n102 ) , .A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n123 ) );
  INV_X1 u1_u3_u1_U7 (.A( u1_u3_u1_n147 ) , .ZN( u1_u3_u1_n181 ) );
  NOR2_X1 u1_u3_u1_U70 (.A2( u1_u3_X_7 ) , .A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n95 ) );
  NOR2_X1 u1_u3_u1_U71 (.A1( u1_u3_X_12 ) , .A2( u1_u3_X_9 ) , .ZN( u1_u3_u1_n100 ) );
  NOR2_X1 u1_u3_u1_U72 (.A2( u1_u3_X_8 ) , .A1( u1_u3_u1_n177 ) , .ZN( u1_u3_u1_n99 ) );
  NOR2_X1 u1_u3_u1_U73 (.A2( u1_u3_X_12 ) , .ZN( u1_u3_u1_n102 ) , .A1( u1_u3_u1_n176 ) );
  NOR2_X1 u1_u3_u1_U74 (.A2( u1_u3_X_9 ) , .ZN( u1_u3_u1_n105 ) , .A1( u1_u3_u1_n168 ) );
  NAND2_X1 u1_u3_u1_U75 (.A1( u1_u3_X_10 ) , .ZN( u1_u3_u1_n160 ) , .A2( u1_u3_u1_n169 ) );
  NAND2_X1 u1_u3_u1_U76 (.A2( u1_u3_X_10 ) , .A1( u1_u3_X_11 ) , .ZN( u1_u3_u1_n152 ) );
  NAND2_X1 u1_u3_u1_U77 (.A1( u1_u3_X_11 ) , .ZN( u1_u3_u1_n128 ) , .A2( u1_u3_u1_n170 ) );
  AND2_X1 u1_u3_u1_U78 (.A2( u1_u3_X_7 ) , .A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n104 ) );
  AND2_X1 u1_u3_u1_U79 (.A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n103 ) , .A2( u1_u3_u1_n177 ) );
  NOR2_X1 u1_u3_u1_U8 (.A1( u1_u3_u1_n112 ) , .A2( u1_u3_u1_n116 ) , .ZN( u1_u3_u1_n118 ) );
  INV_X1 u1_u3_u1_U80 (.A( u1_u3_X_10 ) , .ZN( u1_u3_u1_n170 ) );
  INV_X1 u1_u3_u1_U81 (.A( u1_u3_X_9 ) , .ZN( u1_u3_u1_n176 ) );
  INV_X1 u1_u3_u1_U82 (.A( u1_u3_X_11 ) , .ZN( u1_u3_u1_n169 ) );
  INV_X1 u1_u3_u1_U83 (.A( u1_u3_X_12 ) , .ZN( u1_u3_u1_n168 ) );
  INV_X1 u1_u3_u1_U84 (.A( u1_u3_X_7 ) , .ZN( u1_u3_u1_n177 ) );
  NAND4_X1 u1_u3_u1_U85 (.ZN( u1_out3_18 ) , .A4( u1_u3_u1_n165 ) , .A3( u1_u3_u1_n166 ) , .A1( u1_u3_u1_n167 ) , .A2( u1_u3_u1_n186 ) );
  AOI22_X1 u1_u3_u1_U86 (.B2( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n147 ) , .A2( u1_u3_u1_n148 ) , .ZN( u1_u3_u1_n166 ) , .A1( u1_u3_u1_n172 ) );
  INV_X1 u1_u3_u1_U87 (.A( u1_u3_u1_n145 ) , .ZN( u1_u3_u1_n186 ) );
  OR4_X1 u1_u3_u1_U88 (.ZN( u1_out3_13 ) , .A4( u1_u3_u1_n108 ) , .A3( u1_u3_u1_n109 ) , .A2( u1_u3_u1_n110 ) , .A1( u1_u3_u1_n111 ) );
  AOI21_X1 u1_u3_u1_U89 (.ZN( u1_u3_u1_n111 ) , .A( u1_u3_u1_n128 ) , .B2( u1_u3_u1_n131 ) , .B1( u1_u3_u1_n135 ) );
  OAI21_X1 u1_u3_u1_U9 (.ZN( u1_u3_u1_n101 ) , .B1( u1_u3_u1_n141 ) , .A( u1_u3_u1_n146 ) , .B2( u1_u3_u1_n183 ) );
  AOI21_X1 u1_u3_u1_U90 (.ZN( u1_u3_u1_n110 ) , .A( u1_u3_u1_n116 ) , .B1( u1_u3_u1_n152 ) , .B2( u1_u3_u1_n160 ) );
  NAND4_X1 u1_u3_u1_U91 (.ZN( u1_out3_2 ) , .A4( u1_u3_u1_n142 ) , .A3( u1_u3_u1_n143 ) , .A2( u1_u3_u1_n144 ) , .A1( u1_u3_u1_n179 ) );
  INV_X1 u1_u3_u1_U92 (.A( u1_u3_u1_n130 ) , .ZN( u1_u3_u1_n179 ) );
  OAI21_X1 u1_u3_u1_U93 (.B2( u1_u3_u1_n132 ) , .ZN( u1_u3_u1_n144 ) , .A( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n180 ) );
  NAND4_X1 u1_u3_u1_U94 (.ZN( u1_out3_28 ) , .A4( u1_u3_u1_n124 ) , .A3( u1_u3_u1_n125 ) , .A2( u1_u3_u1_n126 ) , .A1( u1_u3_u1_n127 ) );
  OAI21_X1 u1_u3_u1_U95 (.ZN( u1_u3_u1_n127 ) , .B2( u1_u3_u1_n139 ) , .B1( u1_u3_u1_n175 ) , .A( u1_u3_u1_n183 ) );
  OAI21_X1 u1_u3_u1_U96 (.ZN( u1_u3_u1_n126 ) , .B2( u1_u3_u1_n140 ) , .A( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n178 ) );
  NAND3_X1 u1_u3_u1_U97 (.A3( u1_u3_u1_n149 ) , .A2( u1_u3_u1_n150 ) , .A1( u1_u3_u1_n151 ) , .ZN( u1_u3_u1_n164 ) );
  NAND3_X1 u1_u3_u1_U98 (.A3( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n135 ) , .ZN( u1_u3_u1_n136 ) , .A1( u1_u3_u1_n151 ) );
  NAND3_X1 u1_u3_u1_U99 (.A1( u1_u3_u1_n133 ) , .ZN( u1_u3_u1_n137 ) , .A2( u1_u3_u1_n154 ) , .A3( u1_u3_u1_n181 ) );
  XOR2_X1 u1_u4_U33 (.B( u1_K5_24 ) , .A( u1_R3_17 ) , .Z( u1_u4_X_24 ) );
  XOR2_X1 u1_u4_U34 (.B( u1_K5_23 ) , .A( u1_R3_16 ) , .Z( u1_u4_X_23 ) );
  XOR2_X1 u1_u4_U35 (.B( u1_K5_22 ) , .A( u1_R3_15 ) , .Z( u1_u4_X_22 ) );
  XOR2_X1 u1_u4_U37 (.B( u1_K5_20 ) , .A( u1_R3_13 ) , .Z( u1_u4_X_20 ) );
  XOR2_X1 u1_u4_U39 (.B( u1_K5_19 ) , .A( u1_R3_12 ) , .Z( u1_u4_X_19 ) );
  OAI22_X1 u1_u4_u3_U10 (.B1( u1_u4_u3_n113 ) , .A2( u1_u4_u3_n135 ) , .A1( u1_u4_u3_n150 ) , .B2( u1_u4_u3_n164 ) , .ZN( u1_u4_u3_n98 ) );
  OAI211_X1 u1_u4_u3_U11 (.B( u1_u4_u3_n106 ) , .ZN( u1_u4_u3_n119 ) , .C2( u1_u4_u3_n128 ) , .C1( u1_u4_u3_n167 ) , .A( u1_u4_u3_n181 ) );
  AOI221_X1 u1_u4_u3_U12 (.C1( u1_u4_u3_n105 ) , .ZN( u1_u4_u3_n106 ) , .A( u1_u4_u3_n131 ) , .B2( u1_u4_u3_n132 ) , .C2( u1_u4_u3_n133 ) , .B1( u1_u4_u3_n169 ) );
  INV_X1 u1_u4_u3_U13 (.ZN( u1_u4_u3_n181 ) , .A( u1_u4_u3_n98 ) );
  NAND2_X1 u1_u4_u3_U14 (.ZN( u1_u4_u3_n105 ) , .A2( u1_u4_u3_n130 ) , .A1( u1_u4_u3_n155 ) );
  AOI22_X1 u1_u4_u3_U15 (.B1( u1_u4_u3_n115 ) , .A2( u1_u4_u3_n116 ) , .ZN( u1_u4_u3_n123 ) , .B2( u1_u4_u3_n133 ) , .A1( u1_u4_u3_n169 ) );
  NAND2_X1 u1_u4_u3_U16 (.ZN( u1_u4_u3_n116 ) , .A2( u1_u4_u3_n151 ) , .A1( u1_u4_u3_n182 ) );
  NOR2_X1 u1_u4_u3_U17 (.ZN( u1_u4_u3_n126 ) , .A2( u1_u4_u3_n150 ) , .A1( u1_u4_u3_n164 ) );
  AOI21_X1 u1_u4_u3_U18 (.ZN( u1_u4_u3_n112 ) , .B2( u1_u4_u3_n146 ) , .B1( u1_u4_u3_n155 ) , .A( u1_u4_u3_n167 ) );
  NAND2_X1 u1_u4_u3_U19 (.A1( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n142 ) , .A2( u1_u4_u3_n164 ) );
  NAND2_X1 u1_u4_u3_U20 (.ZN( u1_u4_u3_n132 ) , .A2( u1_u4_u3_n152 ) , .A1( u1_u4_u3_n156 ) );
  AND2_X1 u1_u4_u3_U21 (.A2( u1_u4_u3_n113 ) , .A1( u1_u4_u3_n114 ) , .ZN( u1_u4_u3_n151 ) );
  INV_X1 u1_u4_u3_U22 (.A( u1_u4_u3_n133 ) , .ZN( u1_u4_u3_n165 ) );
  INV_X1 u1_u4_u3_U23 (.A( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n170 ) );
  NAND2_X1 u1_u4_u3_U24 (.A1( u1_u4_u3_n107 ) , .A2( u1_u4_u3_n108 ) , .ZN( u1_u4_u3_n140 ) );
  NAND2_X1 u1_u4_u3_U25 (.ZN( u1_u4_u3_n117 ) , .A1( u1_u4_u3_n124 ) , .A2( u1_u4_u3_n148 ) );
  NAND2_X1 u1_u4_u3_U26 (.ZN( u1_u4_u3_n143 ) , .A1( u1_u4_u3_n165 ) , .A2( u1_u4_u3_n167 ) );
  INV_X1 u1_u4_u3_U27 (.A( u1_u4_u3_n130 ) , .ZN( u1_u4_u3_n177 ) );
  INV_X1 u1_u4_u3_U28 (.A( u1_u4_u3_n128 ) , .ZN( u1_u4_u3_n176 ) );
  INV_X1 u1_u4_u3_U29 (.A( u1_u4_u3_n155 ) , .ZN( u1_u4_u3_n174 ) );
  INV_X1 u1_u4_u3_U3 (.A( u1_u4_u3_n129 ) , .ZN( u1_u4_u3_n183 ) );
  INV_X1 u1_u4_u3_U30 (.A( u1_u4_u3_n139 ) , .ZN( u1_u4_u3_n185 ) );
  NOR2_X1 u1_u4_u3_U31 (.ZN( u1_u4_u3_n135 ) , .A2( u1_u4_u3_n141 ) , .A1( u1_u4_u3_n169 ) );
  OAI222_X1 u1_u4_u3_U32 (.C2( u1_u4_u3_n107 ) , .A2( u1_u4_u3_n108 ) , .B1( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n138 ) , .B2( u1_u4_u3_n146 ) , .C1( u1_u4_u3_n154 ) , .A1( u1_u4_u3_n164 ) );
  NOR4_X1 u1_u4_u3_U33 (.A4( u1_u4_u3_n157 ) , .A3( u1_u4_u3_n158 ) , .A2( u1_u4_u3_n159 ) , .A1( u1_u4_u3_n160 ) , .ZN( u1_u4_u3_n161 ) );
  AOI21_X1 u1_u4_u3_U34 (.B2( u1_u4_u3_n152 ) , .B1( u1_u4_u3_n153 ) , .ZN( u1_u4_u3_n158 ) , .A( u1_u4_u3_n164 ) );
  AOI21_X1 u1_u4_u3_U35 (.A( u1_u4_u3_n149 ) , .B2( u1_u4_u3_n150 ) , .B1( u1_u4_u3_n151 ) , .ZN( u1_u4_u3_n159 ) );
  AOI21_X1 u1_u4_u3_U36 (.A( u1_u4_u3_n154 ) , .B2( u1_u4_u3_n155 ) , .B1( u1_u4_u3_n156 ) , .ZN( u1_u4_u3_n157 ) );
  AOI211_X1 u1_u4_u3_U37 (.ZN( u1_u4_u3_n109 ) , .A( u1_u4_u3_n119 ) , .C2( u1_u4_u3_n129 ) , .B( u1_u4_u3_n138 ) , .C1( u1_u4_u3_n141 ) );
  AOI211_X1 u1_u4_u3_U38 (.B( u1_u4_u3_n119 ) , .A( u1_u4_u3_n120 ) , .C2( u1_u4_u3_n121 ) , .ZN( u1_u4_u3_n122 ) , .C1( u1_u4_u3_n179 ) );
  INV_X1 u1_u4_u3_U39 (.A( u1_u4_u3_n156 ) , .ZN( u1_u4_u3_n179 ) );
  INV_X1 u1_u4_u3_U4 (.A( u1_u4_u3_n140 ) , .ZN( u1_u4_u3_n182 ) );
  OAI22_X1 u1_u4_u3_U40 (.B1( u1_u4_u3_n118 ) , .ZN( u1_u4_u3_n120 ) , .A1( u1_u4_u3_n135 ) , .B2( u1_u4_u3_n154 ) , .A2( u1_u4_u3_n178 ) );
  AND3_X1 u1_u4_u3_U41 (.ZN( u1_u4_u3_n118 ) , .A2( u1_u4_u3_n124 ) , .A1( u1_u4_u3_n144 ) , .A3( u1_u4_u3_n152 ) );
  INV_X1 u1_u4_u3_U42 (.A( u1_u4_u3_n121 ) , .ZN( u1_u4_u3_n164 ) );
  NAND2_X1 u1_u4_u3_U43 (.ZN( u1_u4_u3_n133 ) , .A1( u1_u4_u3_n154 ) , .A2( u1_u4_u3_n164 ) );
  OAI211_X1 u1_u4_u3_U44 (.B( u1_u4_u3_n127 ) , .ZN( u1_u4_u3_n139 ) , .C1( u1_u4_u3_n150 ) , .C2( u1_u4_u3_n154 ) , .A( u1_u4_u3_n184 ) );
  INV_X1 u1_u4_u3_U45 (.A( u1_u4_u3_n125 ) , .ZN( u1_u4_u3_n184 ) );
  AOI221_X1 u1_u4_u3_U46 (.A( u1_u4_u3_n126 ) , .ZN( u1_u4_u3_n127 ) , .C2( u1_u4_u3_n132 ) , .C1( u1_u4_u3_n169 ) , .B2( u1_u4_u3_n170 ) , .B1( u1_u4_u3_n174 ) );
  OAI22_X1 u1_u4_u3_U47 (.A1( u1_u4_u3_n124 ) , .ZN( u1_u4_u3_n125 ) , .B2( u1_u4_u3_n145 ) , .A2( u1_u4_u3_n165 ) , .B1( u1_u4_u3_n167 ) );
  NOR2_X1 u1_u4_u3_U48 (.A1( u1_u4_u3_n113 ) , .ZN( u1_u4_u3_n131 ) , .A2( u1_u4_u3_n154 ) );
  NAND2_X1 u1_u4_u3_U49 (.A1( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n150 ) , .A2( u1_u4_u3_n99 ) );
  INV_X1 u1_u4_u3_U5 (.A( u1_u4_u3_n117 ) , .ZN( u1_u4_u3_n178 ) );
  NAND2_X1 u1_u4_u3_U50 (.A2( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n155 ) , .A1( u1_u4_u3_n97 ) );
  INV_X1 u1_u4_u3_U51 (.A( u1_u4_u3_n141 ) , .ZN( u1_u4_u3_n167 ) );
  AOI21_X1 u1_u4_u3_U52 (.B2( u1_u4_u3_n114 ) , .B1( u1_u4_u3_n146 ) , .A( u1_u4_u3_n154 ) , .ZN( u1_u4_u3_n94 ) );
  AOI21_X1 u1_u4_u3_U53 (.ZN( u1_u4_u3_n110 ) , .B2( u1_u4_u3_n142 ) , .B1( u1_u4_u3_n186 ) , .A( u1_u4_u3_n95 ) );
  INV_X1 u1_u4_u3_U54 (.A( u1_u4_u3_n145 ) , .ZN( u1_u4_u3_n186 ) );
  AOI21_X1 u1_u4_u3_U55 (.B1( u1_u4_u3_n124 ) , .A( u1_u4_u3_n149 ) , .B2( u1_u4_u3_n155 ) , .ZN( u1_u4_u3_n95 ) );
  INV_X1 u1_u4_u3_U56 (.A( u1_u4_u3_n149 ) , .ZN( u1_u4_u3_n169 ) );
  NAND2_X1 u1_u4_u3_U57 (.ZN( u1_u4_u3_n124 ) , .A1( u1_u4_u3_n96 ) , .A2( u1_u4_u3_n97 ) );
  NAND2_X1 u1_u4_u3_U58 (.A2( u1_u4_u3_n100 ) , .ZN( u1_u4_u3_n146 ) , .A1( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U59 (.A1( u1_u4_u3_n101 ) , .ZN( u1_u4_u3_n145 ) , .A2( u1_u4_u3_n99 ) );
  AOI221_X1 u1_u4_u3_U6 (.A( u1_u4_u3_n131 ) , .C2( u1_u4_u3_n132 ) , .C1( u1_u4_u3_n133 ) , .ZN( u1_u4_u3_n134 ) , .B1( u1_u4_u3_n143 ) , .B2( u1_u4_u3_n177 ) );
  NAND2_X1 u1_u4_u3_U60 (.A1( u1_u4_u3_n100 ) , .ZN( u1_u4_u3_n156 ) , .A2( u1_u4_u3_n99 ) );
  NAND2_X1 u1_u4_u3_U61 (.A2( u1_u4_u3_n101 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n148 ) );
  NAND2_X1 u1_u4_u3_U62 (.A1( u1_u4_u3_n100 ) , .A2( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n128 ) );
  NAND2_X1 u1_u4_u3_U63 (.A2( u1_u4_u3_n101 ) , .A1( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n152 ) );
  NAND2_X1 u1_u4_u3_U64 (.A2( u1_u4_u3_n101 ) , .ZN( u1_u4_u3_n114 ) , .A1( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U65 (.ZN( u1_u4_u3_n107 ) , .A1( u1_u4_u3_n97 ) , .A2( u1_u4_u3_n99 ) );
  NAND2_X1 u1_u4_u3_U66 (.A2( u1_u4_u3_n100 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n113 ) );
  NAND2_X1 u1_u4_u3_U67 (.A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n153 ) , .A2( u1_u4_u3_n97 ) );
  NAND2_X1 u1_u4_u3_U68 (.A2( u1_u4_u3_n103 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n130 ) );
  NAND2_X1 u1_u4_u3_U69 (.A2( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n144 ) , .A1( u1_u4_u3_n96 ) );
  OAI22_X1 u1_u4_u3_U7 (.B2( u1_u4_u3_n147 ) , .A2( u1_u4_u3_n148 ) , .ZN( u1_u4_u3_n160 ) , .B1( u1_u4_u3_n165 ) , .A1( u1_u4_u3_n168 ) );
  NAND2_X1 u1_u4_u3_U70 (.A1( u1_u4_u3_n102 ) , .A2( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n108 ) );
  NOR2_X1 u1_u4_u3_U71 (.A2( u1_u4_X_19 ) , .A1( u1_u4_X_20 ) , .ZN( u1_u4_u3_n99 ) );
  NOR2_X1 u1_u4_u3_U72 (.A2( u1_u4_X_21 ) , .A1( u1_u4_X_24 ) , .ZN( u1_u4_u3_n103 ) );
  NOR2_X1 u1_u4_u3_U73 (.A2( u1_u4_X_24 ) , .A1( u1_u4_u3_n171 ) , .ZN( u1_u4_u3_n97 ) );
  NOR2_X1 u1_u4_u3_U74 (.A2( u1_u4_X_23 ) , .ZN( u1_u4_u3_n141 ) , .A1( u1_u4_u3_n166 ) );
  NOR2_X1 u1_u4_u3_U75 (.A2( u1_u4_X_19 ) , .A1( u1_u4_u3_n172 ) , .ZN( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U76 (.A1( u1_u4_X_22 ) , .A2( u1_u4_X_23 ) , .ZN( u1_u4_u3_n154 ) );
  NAND2_X1 u1_u4_u3_U77 (.A1( u1_u4_X_23 ) , .ZN( u1_u4_u3_n149 ) , .A2( u1_u4_u3_n166 ) );
  NOR2_X1 u1_u4_u3_U78 (.A2( u1_u4_X_22 ) , .A1( u1_u4_X_23 ) , .ZN( u1_u4_u3_n121 ) );
  AND2_X1 u1_u4_u3_U79 (.A1( u1_u4_X_24 ) , .ZN( u1_u4_u3_n101 ) , .A2( u1_u4_u3_n171 ) );
  AND3_X1 u1_u4_u3_U8 (.A3( u1_u4_u3_n144 ) , .A2( u1_u4_u3_n145 ) , .A1( u1_u4_u3_n146 ) , .ZN( u1_u4_u3_n147 ) );
  AND2_X1 u1_u4_u3_U80 (.A1( u1_u4_X_19 ) , .ZN( u1_u4_u3_n102 ) , .A2( u1_u4_u3_n172 ) );
  AND2_X1 u1_u4_u3_U81 (.A1( u1_u4_X_21 ) , .A2( u1_u4_X_24 ) , .ZN( u1_u4_u3_n100 ) );
  AND2_X1 u1_u4_u3_U82 (.A2( u1_u4_X_19 ) , .A1( u1_u4_X_20 ) , .ZN( u1_u4_u3_n104 ) );
  INV_X1 u1_u4_u3_U83 (.A( u1_u4_X_22 ) , .ZN( u1_u4_u3_n166 ) );
  INV_X1 u1_u4_u3_U84 (.A( u1_u4_X_21 ) , .ZN( u1_u4_u3_n171 ) );
  INV_X1 u1_u4_u3_U85 (.A( u1_u4_X_20 ) , .ZN( u1_u4_u3_n172 ) );
  NAND4_X1 u1_u4_u3_U86 (.ZN( u1_out4_26 ) , .A4( u1_u4_u3_n109 ) , .A3( u1_u4_u3_n110 ) , .A2( u1_u4_u3_n111 ) , .A1( u1_u4_u3_n173 ) );
  INV_X1 u1_u4_u3_U87 (.ZN( u1_u4_u3_n173 ) , .A( u1_u4_u3_n94 ) );
  OAI21_X1 u1_u4_u3_U88 (.ZN( u1_u4_u3_n111 ) , .B2( u1_u4_u3_n117 ) , .A( u1_u4_u3_n133 ) , .B1( u1_u4_u3_n176 ) );
  NAND4_X1 u1_u4_u3_U89 (.ZN( u1_out4_20 ) , .A4( u1_u4_u3_n122 ) , .A3( u1_u4_u3_n123 ) , .A1( u1_u4_u3_n175 ) , .A2( u1_u4_u3_n180 ) );
  INV_X1 u1_u4_u3_U9 (.A( u1_u4_u3_n143 ) , .ZN( u1_u4_u3_n168 ) );
  INV_X1 u1_u4_u3_U90 (.A( u1_u4_u3_n126 ) , .ZN( u1_u4_u3_n180 ) );
  INV_X1 u1_u4_u3_U91 (.A( u1_u4_u3_n112 ) , .ZN( u1_u4_u3_n175 ) );
  NAND4_X1 u1_u4_u3_U92 (.ZN( u1_out4_1 ) , .A4( u1_u4_u3_n161 ) , .A3( u1_u4_u3_n162 ) , .A2( u1_u4_u3_n163 ) , .A1( u1_u4_u3_n185 ) );
  NAND2_X1 u1_u4_u3_U93 (.ZN( u1_u4_u3_n163 ) , .A2( u1_u4_u3_n170 ) , .A1( u1_u4_u3_n176 ) );
  AOI22_X1 u1_u4_u3_U94 (.B2( u1_u4_u3_n140 ) , .B1( u1_u4_u3_n141 ) , .A2( u1_u4_u3_n142 ) , .ZN( u1_u4_u3_n162 ) , .A1( u1_u4_u3_n177 ) );
  OR4_X1 u1_u4_u3_U95 (.ZN( u1_out4_10 ) , .A4( u1_u4_u3_n136 ) , .A3( u1_u4_u3_n137 ) , .A1( u1_u4_u3_n138 ) , .A2( u1_u4_u3_n139 ) );
  OAI222_X1 u1_u4_u3_U96 (.C1( u1_u4_u3_n128 ) , .ZN( u1_u4_u3_n137 ) , .B1( u1_u4_u3_n148 ) , .A2( u1_u4_u3_n150 ) , .B2( u1_u4_u3_n154 ) , .C2( u1_u4_u3_n164 ) , .A1( u1_u4_u3_n167 ) );
  OAI221_X1 u1_u4_u3_U97 (.A( u1_u4_u3_n134 ) , .B2( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n136 ) , .C1( u1_u4_u3_n149 ) , .B1( u1_u4_u3_n151 ) , .C2( u1_u4_u3_n183 ) );
  NAND3_X1 u1_u4_u3_U98 (.A1( u1_u4_u3_n114 ) , .ZN( u1_u4_u3_n115 ) , .A2( u1_u4_u3_n145 ) , .A3( u1_u4_u3_n153 ) );
  NAND3_X1 u1_u4_u3_U99 (.ZN( u1_u4_u3_n129 ) , .A2( u1_u4_u3_n144 ) , .A1( u1_u4_u3_n153 ) , .A3( u1_u4_u3_n182 ) );
  XOR2_X1 u1_u5_U20 (.B( u1_K6_36 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_36 ) );
  XOR2_X1 u1_u5_U21 (.B( u1_K6_35 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_35 ) );
  XOR2_X1 u1_u5_U24 (.B( u1_K6_32 ) , .A( u1_R4_21 ) , .Z( u1_u5_X_32 ) );
  XOR2_X1 u1_u5_U25 (.B( u1_K6_31 ) , .A( u1_R4_20 ) , .Z( u1_u5_X_31 ) );
  XOR2_X1 u1_u5_U26 (.B( u1_K6_30 ) , .A( u1_R4_21 ) , .Z( u1_u5_X_30 ) );
  XOR2_X1 u1_u5_U28 (.B( u1_K6_29 ) , .A( u1_R4_20 ) , .Z( u1_u5_X_29 ) );
  XOR2_X1 u1_u5_U31 (.B( u1_K6_26 ) , .A( u1_R4_17 ) , .Z( u1_u5_X_26 ) );
  XOR2_X1 u1_u5_U32 (.B( u1_K6_25 ) , .A( u1_R4_16 ) , .Z( u1_u5_X_25 ) );
  OAI22_X1 u1_u5_u4_U10 (.B2( u1_u5_u4_n135 ) , .ZN( u1_u5_u4_n137 ) , .B1( u1_u5_u4_n153 ) , .A1( u1_u5_u4_n155 ) , .A2( u1_u5_u4_n171 ) );
  AND3_X1 u1_u5_u4_U11 (.A2( u1_u5_u4_n134 ) , .ZN( u1_u5_u4_n135 ) , .A3( u1_u5_u4_n145 ) , .A1( u1_u5_u4_n157 ) );
  NAND2_X1 u1_u5_u4_U12 (.ZN( u1_u5_u4_n132 ) , .A2( u1_u5_u4_n170 ) , .A1( u1_u5_u4_n173 ) );
  AOI21_X1 u1_u5_u4_U13 (.B2( u1_u5_u4_n160 ) , .B1( u1_u5_u4_n161 ) , .ZN( u1_u5_u4_n162 ) , .A( u1_u5_u4_n170 ) );
  AOI21_X1 u1_u5_u4_U14 (.ZN( u1_u5_u4_n107 ) , .B2( u1_u5_u4_n143 ) , .A( u1_u5_u4_n174 ) , .B1( u1_u5_u4_n184 ) );
  AOI21_X1 u1_u5_u4_U15 (.B2( u1_u5_u4_n158 ) , .B1( u1_u5_u4_n159 ) , .ZN( u1_u5_u4_n163 ) , .A( u1_u5_u4_n174 ) );
  AOI21_X1 u1_u5_u4_U16 (.A( u1_u5_u4_n153 ) , .B2( u1_u5_u4_n154 ) , .B1( u1_u5_u4_n155 ) , .ZN( u1_u5_u4_n165 ) );
  AOI21_X1 u1_u5_u4_U17 (.A( u1_u5_u4_n156 ) , .B2( u1_u5_u4_n157 ) , .ZN( u1_u5_u4_n164 ) , .B1( u1_u5_u4_n184 ) );
  INV_X1 u1_u5_u4_U18 (.A( u1_u5_u4_n138 ) , .ZN( u1_u5_u4_n170 ) );
  AND2_X1 u1_u5_u4_U19 (.A2( u1_u5_u4_n120 ) , .ZN( u1_u5_u4_n155 ) , .A1( u1_u5_u4_n160 ) );
  INV_X1 u1_u5_u4_U20 (.A( u1_u5_u4_n156 ) , .ZN( u1_u5_u4_n175 ) );
  NAND2_X1 u1_u5_u4_U21 (.A2( u1_u5_u4_n118 ) , .ZN( u1_u5_u4_n131 ) , .A1( u1_u5_u4_n147 ) );
  NAND2_X1 u1_u5_u4_U22 (.A1( u1_u5_u4_n119 ) , .A2( u1_u5_u4_n120 ) , .ZN( u1_u5_u4_n130 ) );
  NAND2_X1 u1_u5_u4_U23 (.ZN( u1_u5_u4_n117 ) , .A2( u1_u5_u4_n118 ) , .A1( u1_u5_u4_n148 ) );
  NAND2_X1 u1_u5_u4_U24 (.ZN( u1_u5_u4_n129 ) , .A1( u1_u5_u4_n134 ) , .A2( u1_u5_u4_n148 ) );
  AND3_X1 u1_u5_u4_U25 (.A1( u1_u5_u4_n119 ) , .A2( u1_u5_u4_n143 ) , .A3( u1_u5_u4_n154 ) , .ZN( u1_u5_u4_n161 ) );
  AND2_X1 u1_u5_u4_U26 (.A1( u1_u5_u4_n145 ) , .A2( u1_u5_u4_n147 ) , .ZN( u1_u5_u4_n159 ) );
  OR3_X1 u1_u5_u4_U27 (.A3( u1_u5_u4_n114 ) , .A2( u1_u5_u4_n115 ) , .A1( u1_u5_u4_n116 ) , .ZN( u1_u5_u4_n136 ) );
  AOI21_X1 u1_u5_u4_U28 (.A( u1_u5_u4_n113 ) , .ZN( u1_u5_u4_n116 ) , .B2( u1_u5_u4_n173 ) , .B1( u1_u5_u4_n174 ) );
  AOI21_X1 u1_u5_u4_U29 (.ZN( u1_u5_u4_n115 ) , .B2( u1_u5_u4_n145 ) , .B1( u1_u5_u4_n146 ) , .A( u1_u5_u4_n156 ) );
  NOR2_X1 u1_u5_u4_U3 (.ZN( u1_u5_u4_n121 ) , .A1( u1_u5_u4_n181 ) , .A2( u1_u5_u4_n182 ) );
  OAI22_X1 u1_u5_u4_U30 (.ZN( u1_u5_u4_n114 ) , .A2( u1_u5_u4_n121 ) , .B1( u1_u5_u4_n160 ) , .B2( u1_u5_u4_n170 ) , .A1( u1_u5_u4_n171 ) );
  INV_X1 u1_u5_u4_U31 (.A( u1_u5_u4_n158 ) , .ZN( u1_u5_u4_n182 ) );
  INV_X1 u1_u5_u4_U32 (.ZN( u1_u5_u4_n181 ) , .A( u1_u5_u4_n96 ) );
  INV_X1 u1_u5_u4_U33 (.A( u1_u5_u4_n144 ) , .ZN( u1_u5_u4_n179 ) );
  INV_X1 u1_u5_u4_U34 (.A( u1_u5_u4_n157 ) , .ZN( u1_u5_u4_n178 ) );
  NAND2_X1 u1_u5_u4_U35 (.A2( u1_u5_u4_n154 ) , .A1( u1_u5_u4_n96 ) , .ZN( u1_u5_u4_n97 ) );
  INV_X1 u1_u5_u4_U36 (.ZN( u1_u5_u4_n186 ) , .A( u1_u5_u4_n95 ) );
  OAI221_X1 u1_u5_u4_U37 (.C1( u1_u5_u4_n134 ) , .B1( u1_u5_u4_n158 ) , .B2( u1_u5_u4_n171 ) , .C2( u1_u5_u4_n173 ) , .A( u1_u5_u4_n94 ) , .ZN( u1_u5_u4_n95 ) );
  AOI222_X1 u1_u5_u4_U38 (.B2( u1_u5_u4_n132 ) , .A1( u1_u5_u4_n138 ) , .C2( u1_u5_u4_n175 ) , .A2( u1_u5_u4_n179 ) , .C1( u1_u5_u4_n181 ) , .B1( u1_u5_u4_n185 ) , .ZN( u1_u5_u4_n94 ) );
  INV_X1 u1_u5_u4_U39 (.A( u1_u5_u4_n113 ) , .ZN( u1_u5_u4_n185 ) );
  INV_X1 u1_u5_u4_U4 (.A( u1_u5_u4_n117 ) , .ZN( u1_u5_u4_n184 ) );
  INV_X1 u1_u5_u4_U40 (.A( u1_u5_u4_n143 ) , .ZN( u1_u5_u4_n183 ) );
  NOR2_X1 u1_u5_u4_U41 (.ZN( u1_u5_u4_n138 ) , .A1( u1_u5_u4_n168 ) , .A2( u1_u5_u4_n169 ) );
  NOR2_X1 u1_u5_u4_U42 (.A1( u1_u5_u4_n150 ) , .A2( u1_u5_u4_n152 ) , .ZN( u1_u5_u4_n153 ) );
  NOR2_X1 u1_u5_u4_U43 (.A2( u1_u5_u4_n128 ) , .A1( u1_u5_u4_n138 ) , .ZN( u1_u5_u4_n156 ) );
  AOI22_X1 u1_u5_u4_U44 (.B2( u1_u5_u4_n122 ) , .A1( u1_u5_u4_n123 ) , .ZN( u1_u5_u4_n124 ) , .B1( u1_u5_u4_n128 ) , .A2( u1_u5_u4_n172 ) );
  INV_X1 u1_u5_u4_U45 (.A( u1_u5_u4_n153 ) , .ZN( u1_u5_u4_n172 ) );
  NAND2_X1 u1_u5_u4_U46 (.A2( u1_u5_u4_n120 ) , .ZN( u1_u5_u4_n123 ) , .A1( u1_u5_u4_n161 ) );
  AOI22_X1 u1_u5_u4_U47 (.B2( u1_u5_u4_n132 ) , .A2( u1_u5_u4_n133 ) , .ZN( u1_u5_u4_n140 ) , .A1( u1_u5_u4_n150 ) , .B1( u1_u5_u4_n179 ) );
  NAND2_X1 u1_u5_u4_U48 (.ZN( u1_u5_u4_n133 ) , .A2( u1_u5_u4_n146 ) , .A1( u1_u5_u4_n154 ) );
  NAND2_X1 u1_u5_u4_U49 (.A1( u1_u5_u4_n103 ) , .ZN( u1_u5_u4_n154 ) , .A2( u1_u5_u4_n98 ) );
  NOR4_X1 u1_u5_u4_U5 (.A4( u1_u5_u4_n106 ) , .A3( u1_u5_u4_n107 ) , .A2( u1_u5_u4_n108 ) , .A1( u1_u5_u4_n109 ) , .ZN( u1_u5_u4_n110 ) );
  NAND2_X1 u1_u5_u4_U50 (.A1( u1_u5_u4_n101 ) , .ZN( u1_u5_u4_n158 ) , .A2( u1_u5_u4_n99 ) );
  AOI21_X1 u1_u5_u4_U51 (.ZN( u1_u5_u4_n127 ) , .A( u1_u5_u4_n136 ) , .B2( u1_u5_u4_n150 ) , .B1( u1_u5_u4_n180 ) );
  INV_X1 u1_u5_u4_U52 (.A( u1_u5_u4_n160 ) , .ZN( u1_u5_u4_n180 ) );
  NAND2_X1 u1_u5_u4_U53 (.A2( u1_u5_u4_n104 ) , .A1( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n146 ) );
  NAND2_X1 u1_u5_u4_U54 (.A2( u1_u5_u4_n101 ) , .A1( u1_u5_u4_n102 ) , .ZN( u1_u5_u4_n160 ) );
  NAND2_X1 u1_u5_u4_U55 (.ZN( u1_u5_u4_n134 ) , .A1( u1_u5_u4_n98 ) , .A2( u1_u5_u4_n99 ) );
  NAND2_X1 u1_u5_u4_U56 (.A1( u1_u5_u4_n103 ) , .A2( u1_u5_u4_n104 ) , .ZN( u1_u5_u4_n143 ) );
  NAND2_X1 u1_u5_u4_U57 (.A2( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n145 ) , .A1( u1_u5_u4_n98 ) );
  NAND2_X1 u1_u5_u4_U58 (.A1( u1_u5_u4_n100 ) , .A2( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n120 ) );
  NAND2_X1 u1_u5_u4_U59 (.A1( u1_u5_u4_n102 ) , .A2( u1_u5_u4_n104 ) , .ZN( u1_u5_u4_n148 ) );
  AOI21_X1 u1_u5_u4_U6 (.ZN( u1_u5_u4_n106 ) , .B2( u1_u5_u4_n146 ) , .B1( u1_u5_u4_n158 ) , .A( u1_u5_u4_n170 ) );
  NAND2_X1 u1_u5_u4_U60 (.A2( u1_u5_u4_n100 ) , .A1( u1_u5_u4_n103 ) , .ZN( u1_u5_u4_n157 ) );
  INV_X1 u1_u5_u4_U61 (.A( u1_u5_u4_n150 ) , .ZN( u1_u5_u4_n173 ) );
  INV_X1 u1_u5_u4_U62 (.A( u1_u5_u4_n152 ) , .ZN( u1_u5_u4_n171 ) );
  NAND2_X1 u1_u5_u4_U63 (.A1( u1_u5_u4_n100 ) , .ZN( u1_u5_u4_n118 ) , .A2( u1_u5_u4_n99 ) );
  NAND2_X1 u1_u5_u4_U64 (.A2( u1_u5_u4_n100 ) , .A1( u1_u5_u4_n102 ) , .ZN( u1_u5_u4_n144 ) );
  NAND2_X1 u1_u5_u4_U65 (.A2( u1_u5_u4_n101 ) , .A1( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n96 ) );
  INV_X1 u1_u5_u4_U66 (.A( u1_u5_u4_n128 ) , .ZN( u1_u5_u4_n174 ) );
  NAND2_X1 u1_u5_u4_U67 (.A2( u1_u5_u4_n102 ) , .ZN( u1_u5_u4_n119 ) , .A1( u1_u5_u4_n98 ) );
  NAND2_X1 u1_u5_u4_U68 (.A2( u1_u5_u4_n101 ) , .A1( u1_u5_u4_n103 ) , .ZN( u1_u5_u4_n147 ) );
  NAND2_X1 u1_u5_u4_U69 (.A2( u1_u5_u4_n104 ) , .ZN( u1_u5_u4_n113 ) , .A1( u1_u5_u4_n99 ) );
  AOI21_X1 u1_u5_u4_U7 (.ZN( u1_u5_u4_n108 ) , .B2( u1_u5_u4_n134 ) , .B1( u1_u5_u4_n155 ) , .A( u1_u5_u4_n156 ) );
  NOR2_X1 u1_u5_u4_U70 (.A2( u1_u5_X_28 ) , .ZN( u1_u5_u4_n150 ) , .A1( u1_u5_u4_n168 ) );
  NOR2_X1 u1_u5_u4_U71 (.A2( u1_u5_X_29 ) , .ZN( u1_u5_u4_n152 ) , .A1( u1_u5_u4_n169 ) );
  NOR2_X1 u1_u5_u4_U72 (.A2( u1_u5_X_30 ) , .ZN( u1_u5_u4_n105 ) , .A1( u1_u5_u4_n176 ) );
  NOR2_X1 u1_u5_u4_U73 (.A2( u1_u5_X_26 ) , .ZN( u1_u5_u4_n100 ) , .A1( u1_u5_u4_n177 ) );
  NOR2_X1 u1_u5_u4_U74 (.A2( u1_u5_X_28 ) , .A1( u1_u5_X_29 ) , .ZN( u1_u5_u4_n128 ) );
  NOR2_X1 u1_u5_u4_U75 (.A2( u1_u5_X_27 ) , .A1( u1_u5_X_30 ) , .ZN( u1_u5_u4_n102 ) );
  NOR2_X1 u1_u5_u4_U76 (.A2( u1_u5_X_25 ) , .A1( u1_u5_X_26 ) , .ZN( u1_u5_u4_n98 ) );
  AND2_X1 u1_u5_u4_U77 (.A2( u1_u5_X_25 ) , .A1( u1_u5_X_26 ) , .ZN( u1_u5_u4_n104 ) );
  AND2_X1 u1_u5_u4_U78 (.A1( u1_u5_X_30 ) , .A2( u1_u5_u4_n176 ) , .ZN( u1_u5_u4_n99 ) );
  AND2_X1 u1_u5_u4_U79 (.A1( u1_u5_X_26 ) , .ZN( u1_u5_u4_n101 ) , .A2( u1_u5_u4_n177 ) );
  AOI21_X1 u1_u5_u4_U8 (.ZN( u1_u5_u4_n109 ) , .A( u1_u5_u4_n153 ) , .B1( u1_u5_u4_n159 ) , .B2( u1_u5_u4_n184 ) );
  AND2_X1 u1_u5_u4_U80 (.A1( u1_u5_X_27 ) , .A2( u1_u5_X_30 ) , .ZN( u1_u5_u4_n103 ) );
  INV_X1 u1_u5_u4_U81 (.A( u1_u5_X_28 ) , .ZN( u1_u5_u4_n169 ) );
  INV_X1 u1_u5_u4_U82 (.A( u1_u5_X_29 ) , .ZN( u1_u5_u4_n168 ) );
  INV_X1 u1_u5_u4_U83 (.A( u1_u5_X_25 ) , .ZN( u1_u5_u4_n177 ) );
  INV_X1 u1_u5_u4_U84 (.A( u1_u5_X_27 ) , .ZN( u1_u5_u4_n176 ) );
  NAND4_X1 u1_u5_u4_U85 (.ZN( u1_out5_25 ) , .A4( u1_u5_u4_n139 ) , .A3( u1_u5_u4_n140 ) , .A2( u1_u5_u4_n141 ) , .A1( u1_u5_u4_n142 ) );
  OAI21_X1 u1_u5_u4_U86 (.A( u1_u5_u4_n128 ) , .B2( u1_u5_u4_n129 ) , .B1( u1_u5_u4_n130 ) , .ZN( u1_u5_u4_n142 ) );
  OAI21_X1 u1_u5_u4_U87 (.B2( u1_u5_u4_n131 ) , .ZN( u1_u5_u4_n141 ) , .A( u1_u5_u4_n175 ) , .B1( u1_u5_u4_n183 ) );
  NAND4_X1 u1_u5_u4_U88 (.ZN( u1_out5_14 ) , .A4( u1_u5_u4_n124 ) , .A3( u1_u5_u4_n125 ) , .A2( u1_u5_u4_n126 ) , .A1( u1_u5_u4_n127 ) );
  AOI22_X1 u1_u5_u4_U89 (.B2( u1_u5_u4_n117 ) , .ZN( u1_u5_u4_n126 ) , .A1( u1_u5_u4_n129 ) , .B1( u1_u5_u4_n152 ) , .A2( u1_u5_u4_n175 ) );
  AOI211_X1 u1_u5_u4_U9 (.B( u1_u5_u4_n136 ) , .A( u1_u5_u4_n137 ) , .C2( u1_u5_u4_n138 ) , .ZN( u1_u5_u4_n139 ) , .C1( u1_u5_u4_n182 ) );
  AOI22_X1 u1_u5_u4_U90 (.ZN( u1_u5_u4_n125 ) , .B2( u1_u5_u4_n131 ) , .A2( u1_u5_u4_n132 ) , .B1( u1_u5_u4_n138 ) , .A1( u1_u5_u4_n178 ) );
  NAND4_X1 u1_u5_u4_U91 (.ZN( u1_out5_8 ) , .A4( u1_u5_u4_n110 ) , .A3( u1_u5_u4_n111 ) , .A2( u1_u5_u4_n112 ) , .A1( u1_u5_u4_n186 ) );
  NAND2_X1 u1_u5_u4_U92 (.ZN( u1_u5_u4_n112 ) , .A2( u1_u5_u4_n130 ) , .A1( u1_u5_u4_n150 ) );
  AOI22_X1 u1_u5_u4_U93 (.ZN( u1_u5_u4_n111 ) , .B2( u1_u5_u4_n132 ) , .A1( u1_u5_u4_n152 ) , .B1( u1_u5_u4_n178 ) , .A2( u1_u5_u4_n97 ) );
  AOI22_X1 u1_u5_u4_U94 (.B2( u1_u5_u4_n149 ) , .B1( u1_u5_u4_n150 ) , .A2( u1_u5_u4_n151 ) , .A1( u1_u5_u4_n152 ) , .ZN( u1_u5_u4_n167 ) );
  NOR4_X1 u1_u5_u4_U95 (.A4( u1_u5_u4_n162 ) , .A3( u1_u5_u4_n163 ) , .A2( u1_u5_u4_n164 ) , .A1( u1_u5_u4_n165 ) , .ZN( u1_u5_u4_n166 ) );
  NAND3_X1 u1_u5_u4_U96 (.ZN( u1_out5_3 ) , .A3( u1_u5_u4_n166 ) , .A1( u1_u5_u4_n167 ) , .A2( u1_u5_u4_n186 ) );
  NAND3_X1 u1_u5_u4_U97 (.A3( u1_u5_u4_n146 ) , .A2( u1_u5_u4_n147 ) , .A1( u1_u5_u4_n148 ) , .ZN( u1_u5_u4_n149 ) );
  NAND3_X1 u1_u5_u4_U98 (.A3( u1_u5_u4_n143 ) , .A2( u1_u5_u4_n144 ) , .A1( u1_u5_u4_n145 ) , .ZN( u1_u5_u4_n151 ) );
  NAND3_X1 u1_u5_u4_U99 (.A3( u1_u5_u4_n121 ) , .ZN( u1_u5_u4_n122 ) , .A2( u1_u5_u4_n144 ) , .A1( u1_u5_u4_n154 ) );
  INV_X1 u1_u5_u5_U10 (.A( u1_u5_u5_n121 ) , .ZN( u1_u5_u5_n177 ) );
  NOR3_X1 u1_u5_u5_U100 (.A3( u1_u5_u5_n141 ) , .A1( u1_u5_u5_n142 ) , .ZN( u1_u5_u5_n143 ) , .A2( u1_u5_u5_n191 ) );
  NAND4_X1 u1_u5_u5_U101 (.ZN( u1_out5_4 ) , .A4( u1_u5_u5_n112 ) , .A2( u1_u5_u5_n113 ) , .A1( u1_u5_u5_n114 ) , .A3( u1_u5_u5_n195 ) );
  AOI211_X1 u1_u5_u5_U102 (.A( u1_u5_u5_n110 ) , .C1( u1_u5_u5_n111 ) , .ZN( u1_u5_u5_n112 ) , .B( u1_u5_u5_n118 ) , .C2( u1_u5_u5_n177 ) );
  AOI222_X1 u1_u5_u5_U103 (.ZN( u1_u5_u5_n113 ) , .A1( u1_u5_u5_n131 ) , .C1( u1_u5_u5_n148 ) , .B2( u1_u5_u5_n174 ) , .C2( u1_u5_u5_n178 ) , .A2( u1_u5_u5_n179 ) , .B1( u1_u5_u5_n99 ) );
  NAND3_X1 u1_u5_u5_U104 (.A2( u1_u5_u5_n154 ) , .A3( u1_u5_u5_n158 ) , .A1( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n99 ) );
  NOR2_X1 u1_u5_u5_U11 (.ZN( u1_u5_u5_n160 ) , .A2( u1_u5_u5_n173 ) , .A1( u1_u5_u5_n177 ) );
  INV_X1 u1_u5_u5_U12 (.A( u1_u5_u5_n150 ) , .ZN( u1_u5_u5_n174 ) );
  AOI21_X1 u1_u5_u5_U13 (.A( u1_u5_u5_n160 ) , .B2( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n162 ) , .B1( u1_u5_u5_n192 ) );
  INV_X1 u1_u5_u5_U14 (.A( u1_u5_u5_n159 ) , .ZN( u1_u5_u5_n192 ) );
  AOI21_X1 u1_u5_u5_U15 (.A( u1_u5_u5_n156 ) , .B2( u1_u5_u5_n157 ) , .B1( u1_u5_u5_n158 ) , .ZN( u1_u5_u5_n163 ) );
  AOI21_X1 u1_u5_u5_U16 (.B2( u1_u5_u5_n139 ) , .B1( u1_u5_u5_n140 ) , .ZN( u1_u5_u5_n141 ) , .A( u1_u5_u5_n150 ) );
  OAI21_X1 u1_u5_u5_U17 (.A( u1_u5_u5_n133 ) , .B2( u1_u5_u5_n134 ) , .B1( u1_u5_u5_n135 ) , .ZN( u1_u5_u5_n142 ) );
  OAI21_X1 u1_u5_u5_U18 (.ZN( u1_u5_u5_n133 ) , .B2( u1_u5_u5_n147 ) , .A( u1_u5_u5_n173 ) , .B1( u1_u5_u5_n188 ) );
  NAND2_X1 u1_u5_u5_U19 (.A2( u1_u5_u5_n119 ) , .A1( u1_u5_u5_n123 ) , .ZN( u1_u5_u5_n137 ) );
  INV_X1 u1_u5_u5_U20 (.A( u1_u5_u5_n155 ) , .ZN( u1_u5_u5_n194 ) );
  NAND2_X1 u1_u5_u5_U21 (.A1( u1_u5_u5_n121 ) , .ZN( u1_u5_u5_n132 ) , .A2( u1_u5_u5_n172 ) );
  NAND2_X1 u1_u5_u5_U22 (.A2( u1_u5_u5_n122 ) , .ZN( u1_u5_u5_n136 ) , .A1( u1_u5_u5_n154 ) );
  NAND2_X1 u1_u5_u5_U23 (.A2( u1_u5_u5_n119 ) , .A1( u1_u5_u5_n120 ) , .ZN( u1_u5_u5_n159 ) );
  INV_X1 u1_u5_u5_U24 (.A( u1_u5_u5_n156 ) , .ZN( u1_u5_u5_n175 ) );
  INV_X1 u1_u5_u5_U25 (.A( u1_u5_u5_n158 ) , .ZN( u1_u5_u5_n188 ) );
  INV_X1 u1_u5_u5_U26 (.A( u1_u5_u5_n152 ) , .ZN( u1_u5_u5_n179 ) );
  INV_X1 u1_u5_u5_U27 (.A( u1_u5_u5_n140 ) , .ZN( u1_u5_u5_n182 ) );
  INV_X1 u1_u5_u5_U28 (.A( u1_u5_u5_n151 ) , .ZN( u1_u5_u5_n183 ) );
  INV_X1 u1_u5_u5_U29 (.A( u1_u5_u5_n123 ) , .ZN( u1_u5_u5_n185 ) );
  NOR2_X1 u1_u5_u5_U3 (.ZN( u1_u5_u5_n134 ) , .A1( u1_u5_u5_n183 ) , .A2( u1_u5_u5_n190 ) );
  INV_X1 u1_u5_u5_U30 (.A( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n184 ) );
  INV_X1 u1_u5_u5_U31 (.A( u1_u5_u5_n139 ) , .ZN( u1_u5_u5_n189 ) );
  INV_X1 u1_u5_u5_U32 (.A( u1_u5_u5_n157 ) , .ZN( u1_u5_u5_n190 ) );
  INV_X1 u1_u5_u5_U33 (.A( u1_u5_u5_n120 ) , .ZN( u1_u5_u5_n193 ) );
  NAND2_X1 u1_u5_u5_U34 (.ZN( u1_u5_u5_n111 ) , .A1( u1_u5_u5_n140 ) , .A2( u1_u5_u5_n155 ) );
  NOR2_X1 u1_u5_u5_U35 (.ZN( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n170 ) , .A2( u1_u5_u5_n180 ) );
  INV_X1 u1_u5_u5_U36 (.A( u1_u5_u5_n117 ) , .ZN( u1_u5_u5_n196 ) );
  OAI221_X1 u1_u5_u5_U37 (.A( u1_u5_u5_n116 ) , .ZN( u1_u5_u5_n117 ) , .B2( u1_u5_u5_n119 ) , .C1( u1_u5_u5_n153 ) , .C2( u1_u5_u5_n158 ) , .B1( u1_u5_u5_n172 ) );
  AOI222_X1 u1_u5_u5_U38 (.ZN( u1_u5_u5_n116 ) , .B2( u1_u5_u5_n145 ) , .C1( u1_u5_u5_n148 ) , .A2( u1_u5_u5_n174 ) , .C2( u1_u5_u5_n177 ) , .B1( u1_u5_u5_n187 ) , .A1( u1_u5_u5_n193 ) );
  INV_X1 u1_u5_u5_U39 (.A( u1_u5_u5_n115 ) , .ZN( u1_u5_u5_n187 ) );
  INV_X1 u1_u5_u5_U4 (.A( u1_u5_u5_n138 ) , .ZN( u1_u5_u5_n191 ) );
  AOI22_X1 u1_u5_u5_U40 (.B2( u1_u5_u5_n131 ) , .A2( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n169 ) , .B1( u1_u5_u5_n174 ) , .A1( u1_u5_u5_n185 ) );
  NOR2_X1 u1_u5_u5_U41 (.A1( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n150 ) , .A2( u1_u5_u5_n173 ) );
  AOI21_X1 u1_u5_u5_U42 (.A( u1_u5_u5_n118 ) , .B2( u1_u5_u5_n145 ) , .ZN( u1_u5_u5_n168 ) , .B1( u1_u5_u5_n186 ) );
  INV_X1 u1_u5_u5_U43 (.A( u1_u5_u5_n122 ) , .ZN( u1_u5_u5_n186 ) );
  NOR2_X1 u1_u5_u5_U44 (.A1( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n152 ) , .A2( u1_u5_u5_n176 ) );
  NOR2_X1 u1_u5_u5_U45 (.A1( u1_u5_u5_n115 ) , .ZN( u1_u5_u5_n118 ) , .A2( u1_u5_u5_n153 ) );
  NOR2_X1 u1_u5_u5_U46 (.A2( u1_u5_u5_n145 ) , .ZN( u1_u5_u5_n156 ) , .A1( u1_u5_u5_n174 ) );
  NOR2_X1 u1_u5_u5_U47 (.ZN( u1_u5_u5_n121 ) , .A2( u1_u5_u5_n145 ) , .A1( u1_u5_u5_n176 ) );
  AOI22_X1 u1_u5_u5_U48 (.ZN( u1_u5_u5_n114 ) , .A2( u1_u5_u5_n137 ) , .A1( u1_u5_u5_n145 ) , .B2( u1_u5_u5_n175 ) , .B1( u1_u5_u5_n193 ) );
  OAI211_X1 u1_u5_u5_U49 (.B( u1_u5_u5_n124 ) , .A( u1_u5_u5_n125 ) , .C2( u1_u5_u5_n126 ) , .C1( u1_u5_u5_n127 ) , .ZN( u1_u5_u5_n128 ) );
  OAI21_X1 u1_u5_u5_U5 (.B2( u1_u5_u5_n136 ) , .B1( u1_u5_u5_n137 ) , .ZN( u1_u5_u5_n138 ) , .A( u1_u5_u5_n177 ) );
  NOR3_X1 u1_u5_u5_U50 (.ZN( u1_u5_u5_n127 ) , .A1( u1_u5_u5_n136 ) , .A3( u1_u5_u5_n148 ) , .A2( u1_u5_u5_n182 ) );
  OAI21_X1 u1_u5_u5_U51 (.ZN( u1_u5_u5_n124 ) , .A( u1_u5_u5_n177 ) , .B2( u1_u5_u5_n183 ) , .B1( u1_u5_u5_n189 ) );
  OAI21_X1 u1_u5_u5_U52 (.ZN( u1_u5_u5_n125 ) , .A( u1_u5_u5_n174 ) , .B2( u1_u5_u5_n185 ) , .B1( u1_u5_u5_n190 ) );
  AOI21_X1 u1_u5_u5_U53 (.A( u1_u5_u5_n153 ) , .B2( u1_u5_u5_n154 ) , .B1( u1_u5_u5_n155 ) , .ZN( u1_u5_u5_n164 ) );
  AOI21_X1 u1_u5_u5_U54 (.ZN( u1_u5_u5_n110 ) , .B1( u1_u5_u5_n122 ) , .B2( u1_u5_u5_n139 ) , .A( u1_u5_u5_n153 ) );
  INV_X1 u1_u5_u5_U55 (.A( u1_u5_u5_n153 ) , .ZN( u1_u5_u5_n176 ) );
  INV_X1 u1_u5_u5_U56 (.A( u1_u5_u5_n126 ) , .ZN( u1_u5_u5_n173 ) );
  AND2_X1 u1_u5_u5_U57 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n147 ) );
  AND2_X1 u1_u5_u5_U58 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n148 ) );
  NAND2_X1 u1_u5_u5_U59 (.A1( u1_u5_u5_n105 ) , .A2( u1_u5_u5_n106 ) , .ZN( u1_u5_u5_n158 ) );
  INV_X1 u1_u5_u5_U6 (.A( u1_u5_u5_n135 ) , .ZN( u1_u5_u5_n178 ) );
  NAND2_X1 u1_u5_u5_U60 (.A2( u1_u5_u5_n108 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n139 ) );
  NAND2_X1 u1_u5_u5_U61 (.A1( u1_u5_u5_n106 ) , .A2( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n119 ) );
  NAND2_X1 u1_u5_u5_U62 (.A2( u1_u5_u5_n103 ) , .A1( u1_u5_u5_n105 ) , .ZN( u1_u5_u5_n140 ) );
  NAND2_X1 u1_u5_u5_U63 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n105 ) , .ZN( u1_u5_u5_n155 ) );
  NAND2_X1 u1_u5_u5_U64 (.A2( u1_u5_u5_n106 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n122 ) );
  NAND2_X1 u1_u5_u5_U65 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n106 ) , .ZN( u1_u5_u5_n115 ) );
  NAND2_X1 u1_u5_u5_U66 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n103 ) , .ZN( u1_u5_u5_n161 ) );
  NAND2_X1 u1_u5_u5_U67 (.A1( u1_u5_u5_n105 ) , .A2( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n154 ) );
  INV_X1 u1_u5_u5_U68 (.A( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n172 ) );
  NAND2_X1 u1_u5_u5_U69 (.A1( u1_u5_u5_n103 ) , .A2( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n123 ) );
  OAI22_X1 u1_u5_u5_U7 (.B2( u1_u5_u5_n149 ) , .B1( u1_u5_u5_n150 ) , .A2( u1_u5_u5_n151 ) , .A1( u1_u5_u5_n152 ) , .ZN( u1_u5_u5_n165 ) );
  NAND2_X1 u1_u5_u5_U70 (.A2( u1_u5_u5_n103 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n151 ) );
  NAND2_X1 u1_u5_u5_U71 (.A2( u1_u5_u5_n107 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n120 ) );
  NAND2_X1 u1_u5_u5_U72 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n157 ) );
  AND2_X1 u1_u5_u5_U73 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n104 ) , .ZN( u1_u5_u5_n131 ) );
  INV_X1 u1_u5_u5_U74 (.A( u1_u5_u5_n102 ) , .ZN( u1_u5_u5_n195 ) );
  OAI221_X1 u1_u5_u5_U75 (.A( u1_u5_u5_n101 ) , .ZN( u1_u5_u5_n102 ) , .C2( u1_u5_u5_n115 ) , .C1( u1_u5_u5_n126 ) , .B1( u1_u5_u5_n134 ) , .B2( u1_u5_u5_n160 ) );
  OAI21_X1 u1_u5_u5_U76 (.ZN( u1_u5_u5_n101 ) , .B1( u1_u5_u5_n137 ) , .A( u1_u5_u5_n146 ) , .B2( u1_u5_u5_n147 ) );
  NOR2_X1 u1_u5_u5_U77 (.A2( u1_u5_X_34 ) , .A1( u1_u5_X_35 ) , .ZN( u1_u5_u5_n145 ) );
  NOR2_X1 u1_u5_u5_U78 (.A2( u1_u5_X_34 ) , .ZN( u1_u5_u5_n146 ) , .A1( u1_u5_u5_n171 ) );
  NOR2_X1 u1_u5_u5_U79 (.A2( u1_u5_X_31 ) , .A1( u1_u5_X_32 ) , .ZN( u1_u5_u5_n103 ) );
  NOR3_X1 u1_u5_u5_U8 (.A2( u1_u5_u5_n147 ) , .A1( u1_u5_u5_n148 ) , .ZN( u1_u5_u5_n149 ) , .A3( u1_u5_u5_n194 ) );
  NOR2_X1 u1_u5_u5_U80 (.A2( u1_u5_X_36 ) , .ZN( u1_u5_u5_n105 ) , .A1( u1_u5_u5_n180 ) );
  NOR2_X1 u1_u5_u5_U81 (.A2( u1_u5_X_33 ) , .ZN( u1_u5_u5_n108 ) , .A1( u1_u5_u5_n170 ) );
  NOR2_X1 u1_u5_u5_U82 (.A2( u1_u5_X_33 ) , .A1( u1_u5_X_36 ) , .ZN( u1_u5_u5_n107 ) );
  NOR2_X1 u1_u5_u5_U83 (.A2( u1_u5_X_31 ) , .ZN( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n181 ) );
  NAND2_X1 u1_u5_u5_U84 (.A2( u1_u5_X_34 ) , .A1( u1_u5_X_35 ) , .ZN( u1_u5_u5_n153 ) );
  NAND2_X1 u1_u5_u5_U85 (.A1( u1_u5_X_34 ) , .ZN( u1_u5_u5_n126 ) , .A2( u1_u5_u5_n171 ) );
  AND2_X1 u1_u5_u5_U86 (.A1( u1_u5_X_31 ) , .A2( u1_u5_X_32 ) , .ZN( u1_u5_u5_n106 ) );
  AND2_X1 u1_u5_u5_U87 (.A1( u1_u5_X_31 ) , .ZN( u1_u5_u5_n109 ) , .A2( u1_u5_u5_n181 ) );
  INV_X1 u1_u5_u5_U88 (.A( u1_u5_X_33 ) , .ZN( u1_u5_u5_n180 ) );
  INV_X1 u1_u5_u5_U89 (.A( u1_u5_X_35 ) , .ZN( u1_u5_u5_n171 ) );
  NOR2_X1 u1_u5_u5_U9 (.ZN( u1_u5_u5_n135 ) , .A1( u1_u5_u5_n173 ) , .A2( u1_u5_u5_n176 ) );
  INV_X1 u1_u5_u5_U90 (.A( u1_u5_X_36 ) , .ZN( u1_u5_u5_n170 ) );
  INV_X1 u1_u5_u5_U91 (.A( u1_u5_X_32 ) , .ZN( u1_u5_u5_n181 ) );
  NAND4_X1 u1_u5_u5_U92 (.ZN( u1_out5_29 ) , .A4( u1_u5_u5_n129 ) , .A3( u1_u5_u5_n130 ) , .A2( u1_u5_u5_n168 ) , .A1( u1_u5_u5_n196 ) );
  AOI221_X1 u1_u5_u5_U93 (.A( u1_u5_u5_n128 ) , .ZN( u1_u5_u5_n129 ) , .C2( u1_u5_u5_n132 ) , .B2( u1_u5_u5_n159 ) , .B1( u1_u5_u5_n176 ) , .C1( u1_u5_u5_n184 ) );
  AOI222_X1 u1_u5_u5_U94 (.ZN( u1_u5_u5_n130 ) , .A2( u1_u5_u5_n146 ) , .B1( u1_u5_u5_n147 ) , .C2( u1_u5_u5_n175 ) , .B2( u1_u5_u5_n179 ) , .A1( u1_u5_u5_n188 ) , .C1( u1_u5_u5_n194 ) );
  NAND4_X1 u1_u5_u5_U95 (.ZN( u1_out5_19 ) , .A4( u1_u5_u5_n166 ) , .A3( u1_u5_u5_n167 ) , .A2( u1_u5_u5_n168 ) , .A1( u1_u5_u5_n169 ) );
  AOI22_X1 u1_u5_u5_U96 (.B2( u1_u5_u5_n145 ) , .A2( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n167 ) , .B1( u1_u5_u5_n182 ) , .A1( u1_u5_u5_n189 ) );
  NOR4_X1 u1_u5_u5_U97 (.A4( u1_u5_u5_n162 ) , .A3( u1_u5_u5_n163 ) , .A2( u1_u5_u5_n164 ) , .A1( u1_u5_u5_n165 ) , .ZN( u1_u5_u5_n166 ) );
  NAND4_X1 u1_u5_u5_U98 (.ZN( u1_out5_11 ) , .A4( u1_u5_u5_n143 ) , .A3( u1_u5_u5_n144 ) , .A2( u1_u5_u5_n169 ) , .A1( u1_u5_u5_n196 ) );
  AOI22_X1 u1_u5_u5_U99 (.A2( u1_u5_u5_n132 ) , .ZN( u1_u5_u5_n144 ) , .B2( u1_u5_u5_n145 ) , .B1( u1_u5_u5_n184 ) , .A1( u1_u5_u5_n194 ) );
  XOR2_X1 u1_u6_U11 (.B( u1_K7_44 ) , .A( u1_R5_29 ) , .Z( u1_u6_X_44 ) );
  XOR2_X1 u1_u6_U12 (.B( u1_K7_43 ) , .A( u1_R5_28 ) , .Z( u1_u6_X_43 ) );
  XOR2_X1 u1_u6_U13 (.B( u1_K7_42 ) , .A( u1_R5_29 ) , .Z( u1_u6_X_42 ) );
  XOR2_X1 u1_u6_U14 (.B( u1_K7_41 ) , .A( u1_R5_28 ) , .Z( u1_u6_X_41 ) );
  XOR2_X1 u1_u6_U18 (.B( u1_K7_38 ) , .A( u1_R5_25 ) , .Z( u1_u6_X_38 ) );
  XOR2_X1 u1_u6_U19 (.B( u1_K7_37 ) , .A( u1_R5_24 ) , .Z( u1_u6_X_37 ) );
  XOR2_X1 u1_u6_U2 (.B( u1_K7_8 ) , .A( u1_R5_5 ) , .Z( u1_u6_X_8 ) );
  XOR2_X1 u1_u6_U27 (.B( u1_K7_2 ) , .A( u1_R5_1 ) , .Z( u1_u6_X_2 ) );
  XOR2_X1 u1_u6_U3 (.B( u1_K7_7 ) , .A( u1_R5_4 ) , .Z( u1_u6_X_7 ) );
  XOR2_X1 u1_u6_U38 (.B( u1_K7_1 ) , .A( u1_R5_32 ) , .Z( u1_u6_X_1 ) );
  XOR2_X1 u1_u6_U4 (.B( u1_K7_6 ) , .A( u1_R5_5 ) , .Z( u1_u6_X_6 ) );
  XOR2_X1 u1_u6_U40 (.B( u1_K7_18 ) , .A( u1_R5_13 ) , .Z( u1_u6_X_18 ) );
  XOR2_X1 u1_u6_U41 (.B( u1_K7_17 ) , .A( u1_R5_12 ) , .Z( u1_u6_X_17 ) );
  XOR2_X1 u1_u6_U44 (.B( u1_K7_14 ) , .A( u1_R5_9 ) , .Z( u1_u6_X_14 ) );
  XOR2_X1 u1_u6_U45 (.B( u1_K7_13 ) , .A( u1_R5_8 ) , .Z( u1_u6_X_13 ) );
  XOR2_X1 u1_u6_U46 (.B( u1_K7_12 ) , .A( u1_R5_9 ) , .Z( u1_u6_X_12 ) );
  XOR2_X1 u1_u6_U47 (.B( u1_K7_11 ) , .A( u1_R5_8 ) , .Z( u1_u6_X_11 ) );
  XOR2_X1 u1_u6_U5 (.B( u1_K7_5 ) , .A( u1_R5_4 ) , .Z( u1_u6_X_5 ) );
  XOR2_X1 u1_u6_U7 (.B( u1_K7_48 ) , .A( u1_R5_1 ) , .Z( u1_u6_X_48 ) );
  XOR2_X1 u1_u6_U8 (.B( u1_K7_47 ) , .A( u1_R5_32 ) , .Z( u1_u6_X_47 ) );
  XOR2_X1 u1_u6_U9 (.B( u1_K7_46 ) , .A( u1_R5_31 ) , .Z( u1_u6_X_46 ) );
  AND3_X1 u1_u6_u0_U10 (.A2( u1_u6_u0_n112 ) , .ZN( u1_u6_u0_n127 ) , .A3( u1_u6_u0_n130 ) , .A1( u1_u6_u0_n148 ) );
  NAND2_X1 u1_u6_u0_U11 (.ZN( u1_u6_u0_n113 ) , .A1( u1_u6_u0_n139 ) , .A2( u1_u6_u0_n149 ) );
  AND2_X1 u1_u6_u0_U12 (.ZN( u1_u6_u0_n107 ) , .A1( u1_u6_u0_n130 ) , .A2( u1_u6_u0_n140 ) );
  AND2_X1 u1_u6_u0_U13 (.A2( u1_u6_u0_n129 ) , .A1( u1_u6_u0_n130 ) , .ZN( u1_u6_u0_n151 ) );
  AND2_X1 u1_u6_u0_U14 (.A1( u1_u6_u0_n108 ) , .A2( u1_u6_u0_n125 ) , .ZN( u1_u6_u0_n145 ) );
  INV_X1 u1_u6_u0_U15 (.A( u1_u6_u0_n143 ) , .ZN( u1_u6_u0_n173 ) );
  NOR2_X1 u1_u6_u0_U16 (.A2( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n147 ) , .A1( u1_u6_u0_n160 ) );
  NOR2_X1 u1_u6_u0_U17 (.A1( u1_u6_u0_n163 ) , .A2( u1_u6_u0_n164 ) , .ZN( u1_u6_u0_n95 ) );
  AOI21_X1 u1_u6_u0_U18 (.B1( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n132 ) , .A( u1_u6_u0_n165 ) , .B2( u1_u6_u0_n93 ) );
  INV_X1 u1_u6_u0_U19 (.A( u1_u6_u0_n142 ) , .ZN( u1_u6_u0_n165 ) );
  OAI221_X1 u1_u6_u0_U20 (.C1( u1_u6_u0_n112 ) , .ZN( u1_u6_u0_n120 ) , .B1( u1_u6_u0_n138 ) , .B2( u1_u6_u0_n141 ) , .C2( u1_u6_u0_n147 ) , .A( u1_u6_u0_n172 ) );
  AOI211_X1 u1_u6_u0_U21 (.B( u1_u6_u0_n115 ) , .A( u1_u6_u0_n116 ) , .C2( u1_u6_u0_n117 ) , .C1( u1_u6_u0_n118 ) , .ZN( u1_u6_u0_n119 ) );
  OAI22_X1 u1_u6_u0_U22 (.B1( u1_u6_u0_n125 ) , .ZN( u1_u6_u0_n126 ) , .A1( u1_u6_u0_n138 ) , .A2( u1_u6_u0_n146 ) , .B2( u1_u6_u0_n147 ) );
  OAI22_X1 u1_u6_u0_U23 (.B1( u1_u6_u0_n131 ) , .A1( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n147 ) , .A2( u1_u6_u0_n90 ) , .ZN( u1_u6_u0_n91 ) );
  AND3_X1 u1_u6_u0_U24 (.A3( u1_u6_u0_n121 ) , .A2( u1_u6_u0_n125 ) , .A1( u1_u6_u0_n148 ) , .ZN( u1_u6_u0_n90 ) );
  NAND2_X1 u1_u6_u0_U25 (.A1( u1_u6_u0_n100 ) , .A2( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n125 ) );
  INV_X1 u1_u6_u0_U26 (.A( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n161 ) );
  AOI22_X1 u1_u6_u0_U27 (.B2( u1_u6_u0_n109 ) , .A2( u1_u6_u0_n110 ) , .ZN( u1_u6_u0_n111 ) , .B1( u1_u6_u0_n118 ) , .A1( u1_u6_u0_n160 ) );
  NAND2_X1 u1_u6_u0_U28 (.A1( u1_u6_u0_n100 ) , .ZN( u1_u6_u0_n129 ) , .A2( u1_u6_u0_n95 ) );
  INV_X1 u1_u6_u0_U29 (.A( u1_u6_u0_n118 ) , .ZN( u1_u6_u0_n158 ) );
  INV_X1 u1_u6_u0_U3 (.A( u1_u6_u0_n113 ) , .ZN( u1_u6_u0_n166 ) );
  AOI21_X1 u1_u6_u0_U30 (.ZN( u1_u6_u0_n104 ) , .B1( u1_u6_u0_n107 ) , .B2( u1_u6_u0_n141 ) , .A( u1_u6_u0_n144 ) );
  AOI21_X1 u1_u6_u0_U31 (.B1( u1_u6_u0_n127 ) , .B2( u1_u6_u0_n129 ) , .A( u1_u6_u0_n138 ) , .ZN( u1_u6_u0_n96 ) );
  AOI21_X1 u1_u6_u0_U32 (.ZN( u1_u6_u0_n116 ) , .B2( u1_u6_u0_n142 ) , .A( u1_u6_u0_n144 ) , .B1( u1_u6_u0_n166 ) );
  NAND2_X1 u1_u6_u0_U33 (.A2( u1_u6_u0_n100 ) , .A1( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n139 ) );
  NAND2_X1 u1_u6_u0_U34 (.A2( u1_u6_u0_n100 ) , .ZN( u1_u6_u0_n131 ) , .A1( u1_u6_u0_n92 ) );
  NAND2_X1 u1_u6_u0_U35 (.A1( u1_u6_u0_n101 ) , .A2( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n150 ) );
  INV_X1 u1_u6_u0_U36 (.A( u1_u6_u0_n138 ) , .ZN( u1_u6_u0_n160 ) );
  NAND2_X1 u1_u6_u0_U37 (.A1( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n128 ) , .A2( u1_u6_u0_n95 ) );
  NAND2_X1 u1_u6_u0_U38 (.ZN( u1_u6_u0_n148 ) , .A1( u1_u6_u0_n93 ) , .A2( u1_u6_u0_n95 ) );
  NAND2_X1 u1_u6_u0_U39 (.A2( u1_u6_u0_n102 ) , .A1( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n149 ) );
  AOI21_X1 u1_u6_u0_U4 (.B1( u1_u6_u0_n114 ) , .ZN( u1_u6_u0_n115 ) , .B2( u1_u6_u0_n129 ) , .A( u1_u6_u0_n161 ) );
  NAND2_X1 u1_u6_u0_U40 (.A2( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n114 ) , .A1( u1_u6_u0_n92 ) );
  NAND2_X1 u1_u6_u0_U41 (.A2( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n121 ) , .A1( u1_u6_u0_n93 ) );
  NAND2_X1 u1_u6_u0_U42 (.ZN( u1_u6_u0_n112 ) , .A2( u1_u6_u0_n92 ) , .A1( u1_u6_u0_n93 ) );
  INV_X1 u1_u6_u0_U43 (.ZN( u1_u6_u0_n172 ) , .A( u1_u6_u0_n88 ) );
  OAI222_X1 u1_u6_u0_U44 (.C1( u1_u6_u0_n108 ) , .A1( u1_u6_u0_n125 ) , .B2( u1_u6_u0_n128 ) , .B1( u1_u6_u0_n144 ) , .A2( u1_u6_u0_n158 ) , .C2( u1_u6_u0_n161 ) , .ZN( u1_u6_u0_n88 ) );
  OR3_X1 u1_u6_u0_U45 (.A3( u1_u6_u0_n152 ) , .A2( u1_u6_u0_n153 ) , .A1( u1_u6_u0_n154 ) , .ZN( u1_u6_u0_n155 ) );
  AOI21_X1 u1_u6_u0_U46 (.A( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n145 ) , .B1( u1_u6_u0_n146 ) , .ZN( u1_u6_u0_n154 ) );
  AOI21_X1 u1_u6_u0_U47 (.B2( u1_u6_u0_n150 ) , .B1( u1_u6_u0_n151 ) , .ZN( u1_u6_u0_n152 ) , .A( u1_u6_u0_n158 ) );
  AOI21_X1 u1_u6_u0_U48 (.A( u1_u6_u0_n147 ) , .B2( u1_u6_u0_n148 ) , .B1( u1_u6_u0_n149 ) , .ZN( u1_u6_u0_n153 ) );
  INV_X1 u1_u6_u0_U49 (.ZN( u1_u6_u0_n171 ) , .A( u1_u6_u0_n99 ) );
  AOI21_X1 u1_u6_u0_U5 (.B2( u1_u6_u0_n131 ) , .ZN( u1_u6_u0_n134 ) , .B1( u1_u6_u0_n151 ) , .A( u1_u6_u0_n158 ) );
  OAI211_X1 u1_u6_u0_U50 (.C2( u1_u6_u0_n140 ) , .C1( u1_u6_u0_n161 ) , .A( u1_u6_u0_n169 ) , .B( u1_u6_u0_n98 ) , .ZN( u1_u6_u0_n99 ) );
  INV_X1 u1_u6_u0_U51 (.ZN( u1_u6_u0_n169 ) , .A( u1_u6_u0_n91 ) );
  AOI211_X1 u1_u6_u0_U52 (.C1( u1_u6_u0_n118 ) , .A( u1_u6_u0_n123 ) , .B( u1_u6_u0_n96 ) , .C2( u1_u6_u0_n97 ) , .ZN( u1_u6_u0_n98 ) );
  NOR2_X1 u1_u6_u0_U53 (.A2( u1_u6_X_4 ) , .A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n118 ) );
  NOR2_X1 u1_u6_u0_U54 (.A2( u1_u6_X_2 ) , .ZN( u1_u6_u0_n103 ) , .A1( u1_u6_u0_n164 ) );
  NOR2_X1 u1_u6_u0_U55 (.A2( u1_u6_X_1 ) , .A1( u1_u6_X_2 ) , .ZN( u1_u6_u0_n92 ) );
  NOR2_X1 u1_u6_u0_U56 (.A2( u1_u6_X_1 ) , .ZN( u1_u6_u0_n101 ) , .A1( u1_u6_u0_n163 ) );
  NAND2_X1 u1_u6_u0_U57 (.A2( u1_u6_X_4 ) , .A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n144 ) );
  NOR2_X1 u1_u6_u0_U58 (.A2( u1_u6_X_5 ) , .ZN( u1_u6_u0_n136 ) , .A1( u1_u6_u0_n159 ) );
  NAND2_X1 u1_u6_u0_U59 (.A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n138 ) , .A2( u1_u6_u0_n159 ) );
  NOR2_X1 u1_u6_u0_U6 (.A1( u1_u6_u0_n108 ) , .ZN( u1_u6_u0_n123 ) , .A2( u1_u6_u0_n158 ) );
  AND2_X1 u1_u6_u0_U60 (.A2( u1_u6_X_3 ) , .A1( u1_u6_X_6 ) , .ZN( u1_u6_u0_n102 ) );
  INV_X1 u1_u6_u0_U61 (.A( u1_u6_X_4 ) , .ZN( u1_u6_u0_n159 ) );
  INV_X1 u1_u6_u0_U62 (.A( u1_u6_X_1 ) , .ZN( u1_u6_u0_n164 ) );
  INV_X1 u1_u6_u0_U63 (.A( u1_u6_X_2 ) , .ZN( u1_u6_u0_n163 ) );
  INV_X1 u1_u6_u0_U64 (.A( u1_u6_X_3 ) , .ZN( u1_u6_u0_n162 ) );
  INV_X1 u1_u6_u0_U65 (.A( u1_u6_u0_n126 ) , .ZN( u1_u6_u0_n168 ) );
  AOI211_X1 u1_u6_u0_U66 (.B( u1_u6_u0_n133 ) , .A( u1_u6_u0_n134 ) , .C2( u1_u6_u0_n135 ) , .C1( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n137 ) );
  OR4_X1 u1_u6_u0_U67 (.ZN( u1_out6_17 ) , .A4( u1_u6_u0_n122 ) , .A2( u1_u6_u0_n123 ) , .A1( u1_u6_u0_n124 ) , .A3( u1_u6_u0_n170 ) );
  AOI21_X1 u1_u6_u0_U68 (.B2( u1_u6_u0_n107 ) , .ZN( u1_u6_u0_n124 ) , .B1( u1_u6_u0_n128 ) , .A( u1_u6_u0_n161 ) );
  INV_X1 u1_u6_u0_U69 (.A( u1_u6_u0_n111 ) , .ZN( u1_u6_u0_n170 ) );
  OAI21_X1 u1_u6_u0_U7 (.B1( u1_u6_u0_n150 ) , .B2( u1_u6_u0_n158 ) , .A( u1_u6_u0_n172 ) , .ZN( u1_u6_u0_n89 ) );
  OR4_X1 u1_u6_u0_U70 (.ZN( u1_out6_31 ) , .A4( u1_u6_u0_n155 ) , .A2( u1_u6_u0_n156 ) , .A1( u1_u6_u0_n157 ) , .A3( u1_u6_u0_n173 ) );
  AOI21_X1 u1_u6_u0_U71 (.A( u1_u6_u0_n138 ) , .B2( u1_u6_u0_n139 ) , .B1( u1_u6_u0_n140 ) , .ZN( u1_u6_u0_n157 ) );
  AOI21_X1 u1_u6_u0_U72 (.B2( u1_u6_u0_n141 ) , .B1( u1_u6_u0_n142 ) , .ZN( u1_u6_u0_n156 ) , .A( u1_u6_u0_n161 ) );
  INV_X1 u1_u6_u0_U73 (.ZN( u1_u6_u0_n174 ) , .A( u1_u6_u0_n89 ) );
  AOI211_X1 u1_u6_u0_U74 (.B( u1_u6_u0_n104 ) , .A( u1_u6_u0_n105 ) , .ZN( u1_u6_u0_n106 ) , .C2( u1_u6_u0_n113 ) , .C1( u1_u6_u0_n160 ) );
  OAI221_X1 u1_u6_u0_U75 (.C1( u1_u6_u0_n121 ) , .ZN( u1_u6_u0_n122 ) , .B2( u1_u6_u0_n127 ) , .A( u1_u6_u0_n143 ) , .B1( u1_u6_u0_n144 ) , .C2( u1_u6_u0_n147 ) );
  NOR2_X1 u1_u6_u0_U76 (.A1( u1_u6_u0_n120 ) , .ZN( u1_u6_u0_n143 ) , .A2( u1_u6_u0_n167 ) );
  AOI21_X1 u1_u6_u0_U77 (.B1( u1_u6_u0_n132 ) , .ZN( u1_u6_u0_n133 ) , .A( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n166 ) );
  OAI22_X1 u1_u6_u0_U78 (.ZN( u1_u6_u0_n105 ) , .A2( u1_u6_u0_n132 ) , .B1( u1_u6_u0_n146 ) , .A1( u1_u6_u0_n147 ) , .B2( u1_u6_u0_n161 ) );
  NAND2_X1 u1_u6_u0_U79 (.ZN( u1_u6_u0_n110 ) , .A2( u1_u6_u0_n132 ) , .A1( u1_u6_u0_n145 ) );
  AND2_X1 u1_u6_u0_U8 (.A1( u1_u6_u0_n114 ) , .A2( u1_u6_u0_n121 ) , .ZN( u1_u6_u0_n146 ) );
  INV_X1 u1_u6_u0_U80 (.A( u1_u6_u0_n119 ) , .ZN( u1_u6_u0_n167 ) );
  NAND2_X1 u1_u6_u0_U81 (.A2( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n140 ) , .A1( u1_u6_u0_n94 ) );
  NAND2_X1 u1_u6_u0_U82 (.A1( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n130 ) , .A2( u1_u6_u0_n94 ) );
  NAND2_X1 u1_u6_u0_U83 (.ZN( u1_u6_u0_n108 ) , .A1( u1_u6_u0_n92 ) , .A2( u1_u6_u0_n94 ) );
  AND2_X1 u1_u6_u0_U84 (.A1( u1_u6_X_6 ) , .A2( u1_u6_u0_n162 ) , .ZN( u1_u6_u0_n93 ) );
  NAND2_X1 u1_u6_u0_U85 (.ZN( u1_u6_u0_n142 ) , .A1( u1_u6_u0_n94 ) , .A2( u1_u6_u0_n95 ) );
  NOR2_X1 u1_u6_u0_U86 (.A2( u1_u6_X_6 ) , .ZN( u1_u6_u0_n100 ) , .A1( u1_u6_u0_n162 ) );
  NOR2_X1 u1_u6_u0_U87 (.A2( u1_u6_X_3 ) , .A1( u1_u6_X_6 ) , .ZN( u1_u6_u0_n94 ) );
  NAND3_X1 u1_u6_u0_U88 (.ZN( u1_out6_23 ) , .A3( u1_u6_u0_n137 ) , .A1( u1_u6_u0_n168 ) , .A2( u1_u6_u0_n171 ) );
  NAND3_X1 u1_u6_u0_U89 (.A3( u1_u6_u0_n127 ) , .A2( u1_u6_u0_n128 ) , .ZN( u1_u6_u0_n135 ) , .A1( u1_u6_u0_n150 ) );
  AND2_X1 u1_u6_u0_U9 (.A1( u1_u6_u0_n131 ) , .ZN( u1_u6_u0_n141 ) , .A2( u1_u6_u0_n150 ) );
  NAND3_X1 u1_u6_u0_U90 (.ZN( u1_u6_u0_n117 ) , .A3( u1_u6_u0_n132 ) , .A2( u1_u6_u0_n139 ) , .A1( u1_u6_u0_n148 ) );
  NAND3_X1 u1_u6_u0_U91 (.ZN( u1_u6_u0_n109 ) , .A2( u1_u6_u0_n114 ) , .A3( u1_u6_u0_n140 ) , .A1( u1_u6_u0_n149 ) );
  NAND3_X1 u1_u6_u0_U92 (.ZN( u1_out6_9 ) , .A3( u1_u6_u0_n106 ) , .A2( u1_u6_u0_n171 ) , .A1( u1_u6_u0_n174 ) );
  NAND3_X1 u1_u6_u0_U93 (.A2( u1_u6_u0_n128 ) , .A1( u1_u6_u0_n132 ) , .A3( u1_u6_u0_n146 ) , .ZN( u1_u6_u0_n97 ) );
  NOR2_X1 u1_u6_u1_U10 (.A1( u1_u6_u1_n112 ) , .A2( u1_u6_u1_n116 ) , .ZN( u1_u6_u1_n118 ) );
  NAND3_X1 u1_u6_u1_U100 (.ZN( u1_u6_u1_n113 ) , .A1( u1_u6_u1_n120 ) , .A3( u1_u6_u1_n133 ) , .A2( u1_u6_u1_n155 ) );
  OAI21_X1 u1_u6_u1_U11 (.ZN( u1_u6_u1_n101 ) , .B1( u1_u6_u1_n141 ) , .A( u1_u6_u1_n146 ) , .B2( u1_u6_u1_n183 ) );
  AOI21_X1 u1_u6_u1_U12 (.B2( u1_u6_u1_n155 ) , .B1( u1_u6_u1_n156 ) , .ZN( u1_u6_u1_n157 ) , .A( u1_u6_u1_n174 ) );
  NAND2_X1 u1_u6_u1_U13 (.ZN( u1_u6_u1_n140 ) , .A2( u1_u6_u1_n150 ) , .A1( u1_u6_u1_n155 ) );
  NAND2_X1 u1_u6_u1_U14 (.A1( u1_u6_u1_n131 ) , .ZN( u1_u6_u1_n147 ) , .A2( u1_u6_u1_n153 ) );
  INV_X1 u1_u6_u1_U15 (.A( u1_u6_u1_n139 ) , .ZN( u1_u6_u1_n174 ) );
  OR4_X1 u1_u6_u1_U16 (.A4( u1_u6_u1_n106 ) , .A3( u1_u6_u1_n107 ) , .ZN( u1_u6_u1_n108 ) , .A1( u1_u6_u1_n117 ) , .A2( u1_u6_u1_n184 ) );
  AOI21_X1 u1_u6_u1_U17 (.ZN( u1_u6_u1_n106 ) , .A( u1_u6_u1_n112 ) , .B1( u1_u6_u1_n154 ) , .B2( u1_u6_u1_n156 ) );
  AOI21_X1 u1_u6_u1_U18 (.ZN( u1_u6_u1_n107 ) , .B1( u1_u6_u1_n134 ) , .B2( u1_u6_u1_n149 ) , .A( u1_u6_u1_n174 ) );
  INV_X1 u1_u6_u1_U19 (.A( u1_u6_u1_n101 ) , .ZN( u1_u6_u1_n184 ) );
  INV_X1 u1_u6_u1_U20 (.A( u1_u6_u1_n112 ) , .ZN( u1_u6_u1_n171 ) );
  NAND2_X1 u1_u6_u1_U21 (.ZN( u1_u6_u1_n141 ) , .A1( u1_u6_u1_n153 ) , .A2( u1_u6_u1_n156 ) );
  AND2_X1 u1_u6_u1_U22 (.A1( u1_u6_u1_n123 ) , .ZN( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n161 ) );
  NAND2_X1 u1_u6_u1_U23 (.A2( u1_u6_u1_n115 ) , .A1( u1_u6_u1_n116 ) , .ZN( u1_u6_u1_n148 ) );
  NAND2_X1 u1_u6_u1_U24 (.A2( u1_u6_u1_n133 ) , .A1( u1_u6_u1_n135 ) , .ZN( u1_u6_u1_n159 ) );
  NAND2_X1 u1_u6_u1_U25 (.A2( u1_u6_u1_n115 ) , .A1( u1_u6_u1_n120 ) , .ZN( u1_u6_u1_n132 ) );
  INV_X1 u1_u6_u1_U26 (.A( u1_u6_u1_n154 ) , .ZN( u1_u6_u1_n178 ) );
  INV_X1 u1_u6_u1_U27 (.A( u1_u6_u1_n151 ) , .ZN( u1_u6_u1_n183 ) );
  AND2_X1 u1_u6_u1_U28 (.A1( u1_u6_u1_n129 ) , .A2( u1_u6_u1_n133 ) , .ZN( u1_u6_u1_n149 ) );
  INV_X1 u1_u6_u1_U29 (.A( u1_u6_u1_n131 ) , .ZN( u1_u6_u1_n180 ) );
  INV_X1 u1_u6_u1_U3 (.A( u1_u6_u1_n159 ) , .ZN( u1_u6_u1_n182 ) );
  AOI221_X1 u1_u6_u1_U30 (.B1( u1_u6_u1_n140 ) , .ZN( u1_u6_u1_n167 ) , .B2( u1_u6_u1_n172 ) , .C2( u1_u6_u1_n175 ) , .C1( u1_u6_u1_n178 ) , .A( u1_u6_u1_n188 ) );
  INV_X1 u1_u6_u1_U31 (.ZN( u1_u6_u1_n188 ) , .A( u1_u6_u1_n97 ) );
  AOI211_X1 u1_u6_u1_U32 (.A( u1_u6_u1_n118 ) , .C1( u1_u6_u1_n132 ) , .C2( u1_u6_u1_n139 ) , .B( u1_u6_u1_n96 ) , .ZN( u1_u6_u1_n97 ) );
  AOI21_X1 u1_u6_u1_U33 (.B2( u1_u6_u1_n121 ) , .B1( u1_u6_u1_n135 ) , .A( u1_u6_u1_n152 ) , .ZN( u1_u6_u1_n96 ) );
  OAI221_X1 u1_u6_u1_U34 (.A( u1_u6_u1_n119 ) , .C2( u1_u6_u1_n129 ) , .ZN( u1_u6_u1_n138 ) , .B2( u1_u6_u1_n152 ) , .C1( u1_u6_u1_n174 ) , .B1( u1_u6_u1_n187 ) );
  INV_X1 u1_u6_u1_U35 (.A( u1_u6_u1_n148 ) , .ZN( u1_u6_u1_n187 ) );
  AOI211_X1 u1_u6_u1_U36 (.B( u1_u6_u1_n117 ) , .A( u1_u6_u1_n118 ) , .ZN( u1_u6_u1_n119 ) , .C2( u1_u6_u1_n146 ) , .C1( u1_u6_u1_n159 ) );
  NOR2_X1 u1_u6_u1_U37 (.A1( u1_u6_u1_n168 ) , .A2( u1_u6_u1_n176 ) , .ZN( u1_u6_u1_n98 ) );
  AOI211_X1 u1_u6_u1_U38 (.B( u1_u6_u1_n162 ) , .A( u1_u6_u1_n163 ) , .C2( u1_u6_u1_n164 ) , .ZN( u1_u6_u1_n165 ) , .C1( u1_u6_u1_n171 ) );
  AOI21_X1 u1_u6_u1_U39 (.A( u1_u6_u1_n160 ) , .B2( u1_u6_u1_n161 ) , .ZN( u1_u6_u1_n162 ) , .B1( u1_u6_u1_n182 ) );
  AOI221_X1 u1_u6_u1_U4 (.A( u1_u6_u1_n138 ) , .C2( u1_u6_u1_n139 ) , .C1( u1_u6_u1_n140 ) , .B2( u1_u6_u1_n141 ) , .ZN( u1_u6_u1_n142 ) , .B1( u1_u6_u1_n175 ) );
  OR2_X1 u1_u6_u1_U40 (.A2( u1_u6_u1_n157 ) , .A1( u1_u6_u1_n158 ) , .ZN( u1_u6_u1_n163 ) );
  NAND2_X1 u1_u6_u1_U41 (.A1( u1_u6_u1_n128 ) , .ZN( u1_u6_u1_n146 ) , .A2( u1_u6_u1_n160 ) );
  NAND2_X1 u1_u6_u1_U42 (.A2( u1_u6_u1_n112 ) , .ZN( u1_u6_u1_n139 ) , .A1( u1_u6_u1_n152 ) );
  NAND2_X1 u1_u6_u1_U43 (.A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n156 ) , .A2( u1_u6_u1_n99 ) );
  NOR2_X1 u1_u6_u1_U44 (.ZN( u1_u6_u1_n117 ) , .A1( u1_u6_u1_n121 ) , .A2( u1_u6_u1_n160 ) );
  OAI21_X1 u1_u6_u1_U45 (.B2( u1_u6_u1_n123 ) , .ZN( u1_u6_u1_n145 ) , .B1( u1_u6_u1_n160 ) , .A( u1_u6_u1_n185 ) );
  INV_X1 u1_u6_u1_U46 (.A( u1_u6_u1_n122 ) , .ZN( u1_u6_u1_n185 ) );
  AOI21_X1 u1_u6_u1_U47 (.B2( u1_u6_u1_n120 ) , .B1( u1_u6_u1_n121 ) , .ZN( u1_u6_u1_n122 ) , .A( u1_u6_u1_n128 ) );
  AOI21_X1 u1_u6_u1_U48 (.A( u1_u6_u1_n128 ) , .B2( u1_u6_u1_n129 ) , .ZN( u1_u6_u1_n130 ) , .B1( u1_u6_u1_n150 ) );
  NAND2_X1 u1_u6_u1_U49 (.ZN( u1_u6_u1_n112 ) , .A1( u1_u6_u1_n169 ) , .A2( u1_u6_u1_n170 ) );
  AOI211_X1 u1_u6_u1_U5 (.ZN( u1_u6_u1_n124 ) , .A( u1_u6_u1_n138 ) , .C2( u1_u6_u1_n139 ) , .B( u1_u6_u1_n145 ) , .C1( u1_u6_u1_n147 ) );
  NAND2_X1 u1_u6_u1_U50 (.ZN( u1_u6_u1_n129 ) , .A2( u1_u6_u1_n95 ) , .A1( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U51 (.A1( u1_u6_u1_n102 ) , .ZN( u1_u6_u1_n154 ) , .A2( u1_u6_u1_n99 ) );
  NAND2_X1 u1_u6_u1_U52 (.A2( u1_u6_u1_n100 ) , .ZN( u1_u6_u1_n135 ) , .A1( u1_u6_u1_n99 ) );
  AOI21_X1 u1_u6_u1_U53 (.A( u1_u6_u1_n152 ) , .B2( u1_u6_u1_n153 ) , .B1( u1_u6_u1_n154 ) , .ZN( u1_u6_u1_n158 ) );
  INV_X1 u1_u6_u1_U54 (.A( u1_u6_u1_n160 ) , .ZN( u1_u6_u1_n175 ) );
  NAND2_X1 u1_u6_u1_U55 (.A1( u1_u6_u1_n100 ) , .ZN( u1_u6_u1_n116 ) , .A2( u1_u6_u1_n95 ) );
  NAND2_X1 u1_u6_u1_U56 (.A1( u1_u6_u1_n102 ) , .ZN( u1_u6_u1_n131 ) , .A2( u1_u6_u1_n95 ) );
  NAND2_X1 u1_u6_u1_U57 (.A2( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n121 ) , .A1( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U58 (.A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n153 ) , .A2( u1_u6_u1_n98 ) );
  NAND2_X1 u1_u6_u1_U59 (.A2( u1_u6_u1_n104 ) , .A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n133 ) );
  AOI22_X1 u1_u6_u1_U6 (.B2( u1_u6_u1_n113 ) , .A2( u1_u6_u1_n114 ) , .ZN( u1_u6_u1_n125 ) , .A1( u1_u6_u1_n171 ) , .B1( u1_u6_u1_n173 ) );
  NAND2_X1 u1_u6_u1_U60 (.ZN( u1_u6_u1_n150 ) , .A2( u1_u6_u1_n98 ) , .A1( u1_u6_u1_n99 ) );
  NAND2_X1 u1_u6_u1_U61 (.A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n155 ) , .A2( u1_u6_u1_n95 ) );
  OAI21_X1 u1_u6_u1_U62 (.ZN( u1_u6_u1_n109 ) , .B1( u1_u6_u1_n129 ) , .B2( u1_u6_u1_n160 ) , .A( u1_u6_u1_n167 ) );
  NAND2_X1 u1_u6_u1_U63 (.A2( u1_u6_u1_n100 ) , .A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n120 ) );
  NAND2_X1 u1_u6_u1_U64 (.A1( u1_u6_u1_n102 ) , .A2( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n115 ) );
  NAND2_X1 u1_u6_u1_U65 (.A2( u1_u6_u1_n100 ) , .A1( u1_u6_u1_n104 ) , .ZN( u1_u6_u1_n151 ) );
  NAND2_X1 u1_u6_u1_U66 (.A2( u1_u6_u1_n103 ) , .A1( u1_u6_u1_n105 ) , .ZN( u1_u6_u1_n161 ) );
  INV_X1 u1_u6_u1_U67 (.A( u1_u6_u1_n152 ) , .ZN( u1_u6_u1_n173 ) );
  INV_X1 u1_u6_u1_U68 (.A( u1_u6_u1_n128 ) , .ZN( u1_u6_u1_n172 ) );
  NAND2_X1 u1_u6_u1_U69 (.A2( u1_u6_u1_n102 ) , .A1( u1_u6_u1_n103 ) , .ZN( u1_u6_u1_n123 ) );
  NAND2_X1 u1_u6_u1_U7 (.ZN( u1_u6_u1_n114 ) , .A1( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n156 ) );
  NOR2_X1 u1_u6_u1_U70 (.A2( u1_u6_X_7 ) , .A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n95 ) );
  NOR2_X1 u1_u6_u1_U71 (.A1( u1_u6_X_12 ) , .A2( u1_u6_X_9 ) , .ZN( u1_u6_u1_n100 ) );
  NOR2_X1 u1_u6_u1_U72 (.A2( u1_u6_X_8 ) , .A1( u1_u6_u1_n177 ) , .ZN( u1_u6_u1_n99 ) );
  NOR2_X1 u1_u6_u1_U73 (.A2( u1_u6_X_12 ) , .ZN( u1_u6_u1_n102 ) , .A1( u1_u6_u1_n176 ) );
  NOR2_X1 u1_u6_u1_U74 (.A2( u1_u6_X_9 ) , .ZN( u1_u6_u1_n105 ) , .A1( u1_u6_u1_n168 ) );
  NAND2_X1 u1_u6_u1_U75 (.A1( u1_u6_X_10 ) , .ZN( u1_u6_u1_n160 ) , .A2( u1_u6_u1_n169 ) );
  NAND2_X1 u1_u6_u1_U76 (.A2( u1_u6_X_10 ) , .A1( u1_u6_X_11 ) , .ZN( u1_u6_u1_n152 ) );
  NAND2_X1 u1_u6_u1_U77 (.A1( u1_u6_X_11 ) , .ZN( u1_u6_u1_n128 ) , .A2( u1_u6_u1_n170 ) );
  AND2_X1 u1_u6_u1_U78 (.A2( u1_u6_X_7 ) , .A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n104 ) );
  AND2_X1 u1_u6_u1_U79 (.A1( u1_u6_X_8 ) , .ZN( u1_u6_u1_n103 ) , .A2( u1_u6_u1_n177 ) );
  AOI22_X1 u1_u6_u1_U8 (.B2( u1_u6_u1_n136 ) , .A2( u1_u6_u1_n137 ) , .ZN( u1_u6_u1_n143 ) , .A1( u1_u6_u1_n171 ) , .B1( u1_u6_u1_n173 ) );
  INV_X1 u1_u6_u1_U80 (.A( u1_u6_X_10 ) , .ZN( u1_u6_u1_n170 ) );
  INV_X1 u1_u6_u1_U81 (.A( u1_u6_X_9 ) , .ZN( u1_u6_u1_n176 ) );
  INV_X1 u1_u6_u1_U82 (.A( u1_u6_X_11 ) , .ZN( u1_u6_u1_n169 ) );
  INV_X1 u1_u6_u1_U83 (.A( u1_u6_X_12 ) , .ZN( u1_u6_u1_n168 ) );
  INV_X1 u1_u6_u1_U84 (.A( u1_u6_X_7 ) , .ZN( u1_u6_u1_n177 ) );
  NAND4_X1 u1_u6_u1_U85 (.ZN( u1_out6_18 ) , .A4( u1_u6_u1_n165 ) , .A3( u1_u6_u1_n166 ) , .A1( u1_u6_u1_n167 ) , .A2( u1_u6_u1_n186 ) );
  AOI22_X1 u1_u6_u1_U86 (.B2( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n147 ) , .A2( u1_u6_u1_n148 ) , .ZN( u1_u6_u1_n166 ) , .A1( u1_u6_u1_n172 ) );
  INV_X1 u1_u6_u1_U87 (.A( u1_u6_u1_n145 ) , .ZN( u1_u6_u1_n186 ) );
  NAND4_X1 u1_u6_u1_U88 (.ZN( u1_out6_2 ) , .A4( u1_u6_u1_n142 ) , .A3( u1_u6_u1_n143 ) , .A2( u1_u6_u1_n144 ) , .A1( u1_u6_u1_n179 ) );
  OAI21_X1 u1_u6_u1_U89 (.B2( u1_u6_u1_n132 ) , .ZN( u1_u6_u1_n144 ) , .A( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n180 ) );
  INV_X1 u1_u6_u1_U9 (.A( u1_u6_u1_n147 ) , .ZN( u1_u6_u1_n181 ) );
  INV_X1 u1_u6_u1_U90 (.A( u1_u6_u1_n130 ) , .ZN( u1_u6_u1_n179 ) );
  NAND4_X1 u1_u6_u1_U91 (.ZN( u1_out6_28 ) , .A4( u1_u6_u1_n124 ) , .A3( u1_u6_u1_n125 ) , .A2( u1_u6_u1_n126 ) , .A1( u1_u6_u1_n127 ) );
  OAI21_X1 u1_u6_u1_U92 (.ZN( u1_u6_u1_n127 ) , .B2( u1_u6_u1_n139 ) , .B1( u1_u6_u1_n175 ) , .A( u1_u6_u1_n183 ) );
  OAI21_X1 u1_u6_u1_U93 (.ZN( u1_u6_u1_n126 ) , .B2( u1_u6_u1_n140 ) , .A( u1_u6_u1_n146 ) , .B1( u1_u6_u1_n178 ) );
  OR4_X1 u1_u6_u1_U94 (.ZN( u1_out6_13 ) , .A4( u1_u6_u1_n108 ) , .A3( u1_u6_u1_n109 ) , .A2( u1_u6_u1_n110 ) , .A1( u1_u6_u1_n111 ) );
  AOI21_X1 u1_u6_u1_U95 (.ZN( u1_u6_u1_n111 ) , .A( u1_u6_u1_n128 ) , .B2( u1_u6_u1_n131 ) , .B1( u1_u6_u1_n135 ) );
  AOI21_X1 u1_u6_u1_U96 (.ZN( u1_u6_u1_n110 ) , .A( u1_u6_u1_n116 ) , .B1( u1_u6_u1_n152 ) , .B2( u1_u6_u1_n160 ) );
  NAND3_X1 u1_u6_u1_U97 (.A3( u1_u6_u1_n149 ) , .A2( u1_u6_u1_n150 ) , .A1( u1_u6_u1_n151 ) , .ZN( u1_u6_u1_n164 ) );
  NAND3_X1 u1_u6_u1_U98 (.A3( u1_u6_u1_n134 ) , .A2( u1_u6_u1_n135 ) , .ZN( u1_u6_u1_n136 ) , .A1( u1_u6_u1_n151 ) );
  NAND3_X1 u1_u6_u1_U99 (.A1( u1_u6_u1_n133 ) , .ZN( u1_u6_u1_n137 ) , .A2( u1_u6_u1_n154 ) , .A3( u1_u6_u1_n181 ) );
  OAI22_X1 u1_u6_u2_U10 (.B1( u1_u6_u2_n151 ) , .A2( u1_u6_u2_n152 ) , .A1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n160 ) , .B2( u1_u6_u2_n168 ) );
  NAND3_X1 u1_u6_u2_U100 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n98 ) );
  NOR3_X1 u1_u6_u2_U11 (.A1( u1_u6_u2_n150 ) , .ZN( u1_u6_u2_n151 ) , .A3( u1_u6_u2_n175 ) , .A2( u1_u6_u2_n188 ) );
  AOI21_X1 u1_u6_u2_U12 (.B2( u1_u6_u2_n123 ) , .ZN( u1_u6_u2_n125 ) , .A( u1_u6_u2_n171 ) , .B1( u1_u6_u2_n184 ) );
  INV_X1 u1_u6_u2_U13 (.A( u1_u6_u2_n150 ) , .ZN( u1_u6_u2_n184 ) );
  AOI21_X1 u1_u6_u2_U14 (.ZN( u1_u6_u2_n144 ) , .B2( u1_u6_u2_n155 ) , .A( u1_u6_u2_n172 ) , .B1( u1_u6_u2_n185 ) );
  AOI21_X1 u1_u6_u2_U15 (.B2( u1_u6_u2_n143 ) , .ZN( u1_u6_u2_n145 ) , .B1( u1_u6_u2_n152 ) , .A( u1_u6_u2_n171 ) );
  INV_X1 u1_u6_u2_U16 (.A( u1_u6_u2_n156 ) , .ZN( u1_u6_u2_n171 ) );
  INV_X1 u1_u6_u2_U17 (.A( u1_u6_u2_n120 ) , .ZN( u1_u6_u2_n188 ) );
  NAND2_X1 u1_u6_u2_U18 (.A2( u1_u6_u2_n122 ) , .ZN( u1_u6_u2_n150 ) , .A1( u1_u6_u2_n152 ) );
  INV_X1 u1_u6_u2_U19 (.A( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n170 ) );
  INV_X1 u1_u6_u2_U20 (.A( u1_u6_u2_n137 ) , .ZN( u1_u6_u2_n173 ) );
  NAND2_X1 u1_u6_u2_U21 (.A1( u1_u6_u2_n132 ) , .A2( u1_u6_u2_n139 ) , .ZN( u1_u6_u2_n157 ) );
  INV_X1 u1_u6_u2_U22 (.A( u1_u6_u2_n113 ) , .ZN( u1_u6_u2_n178 ) );
  INV_X1 u1_u6_u2_U23 (.A( u1_u6_u2_n139 ) , .ZN( u1_u6_u2_n175 ) );
  INV_X1 u1_u6_u2_U24 (.A( u1_u6_u2_n155 ) , .ZN( u1_u6_u2_n181 ) );
  INV_X1 u1_u6_u2_U25 (.A( u1_u6_u2_n119 ) , .ZN( u1_u6_u2_n177 ) );
  INV_X1 u1_u6_u2_U26 (.A( u1_u6_u2_n116 ) , .ZN( u1_u6_u2_n180 ) );
  INV_X1 u1_u6_u2_U27 (.A( u1_u6_u2_n131 ) , .ZN( u1_u6_u2_n179 ) );
  INV_X1 u1_u6_u2_U28 (.A( u1_u6_u2_n154 ) , .ZN( u1_u6_u2_n176 ) );
  NAND2_X1 u1_u6_u2_U29 (.A2( u1_u6_u2_n116 ) , .A1( u1_u6_u2_n117 ) , .ZN( u1_u6_u2_n118 ) );
  NOR2_X1 u1_u6_u2_U3 (.ZN( u1_u6_u2_n121 ) , .A2( u1_u6_u2_n177 ) , .A1( u1_u6_u2_n180 ) );
  INV_X1 u1_u6_u2_U30 (.A( u1_u6_u2_n132 ) , .ZN( u1_u6_u2_n182 ) );
  INV_X1 u1_u6_u2_U31 (.A( u1_u6_u2_n158 ) , .ZN( u1_u6_u2_n183 ) );
  OAI21_X1 u1_u6_u2_U32 (.A( u1_u6_u2_n156 ) , .B1( u1_u6_u2_n157 ) , .ZN( u1_u6_u2_n158 ) , .B2( u1_u6_u2_n179 ) );
  NOR2_X1 u1_u6_u2_U33 (.ZN( u1_u6_u2_n156 ) , .A1( u1_u6_u2_n166 ) , .A2( u1_u6_u2_n169 ) );
  NOR2_X1 u1_u6_u2_U34 (.A2( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n137 ) , .A1( u1_u6_u2_n140 ) );
  NOR2_X1 u1_u6_u2_U35 (.A2( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n153 ) , .A1( u1_u6_u2_n156 ) );
  AOI211_X1 u1_u6_u2_U36 (.ZN( u1_u6_u2_n130 ) , .C1( u1_u6_u2_n138 ) , .C2( u1_u6_u2_n179 ) , .B( u1_u6_u2_n96 ) , .A( u1_u6_u2_n97 ) );
  OAI22_X1 u1_u6_u2_U37 (.B1( u1_u6_u2_n133 ) , .A2( u1_u6_u2_n137 ) , .A1( u1_u6_u2_n152 ) , .B2( u1_u6_u2_n168 ) , .ZN( u1_u6_u2_n97 ) );
  OAI221_X1 u1_u6_u2_U38 (.B1( u1_u6_u2_n113 ) , .C1( u1_u6_u2_n132 ) , .A( u1_u6_u2_n149 ) , .B2( u1_u6_u2_n171 ) , .C2( u1_u6_u2_n172 ) , .ZN( u1_u6_u2_n96 ) );
  OAI221_X1 u1_u6_u2_U39 (.A( u1_u6_u2_n115 ) , .C2( u1_u6_u2_n123 ) , .B2( u1_u6_u2_n143 ) , .B1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n163 ) , .C1( u1_u6_u2_n168 ) );
  INV_X1 u1_u6_u2_U4 (.A( u1_u6_u2_n134 ) , .ZN( u1_u6_u2_n185 ) );
  OAI21_X1 u1_u6_u2_U40 (.A( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n115 ) , .B1( u1_u6_u2_n176 ) , .B2( u1_u6_u2_n178 ) );
  OAI221_X1 u1_u6_u2_U41 (.A( u1_u6_u2_n135 ) , .B2( u1_u6_u2_n136 ) , .B1( u1_u6_u2_n137 ) , .ZN( u1_u6_u2_n162 ) , .C2( u1_u6_u2_n167 ) , .C1( u1_u6_u2_n185 ) );
  AND3_X1 u1_u6_u2_U42 (.A3( u1_u6_u2_n131 ) , .A2( u1_u6_u2_n132 ) , .A1( u1_u6_u2_n133 ) , .ZN( u1_u6_u2_n136 ) );
  AOI22_X1 u1_u6_u2_U43 (.ZN( u1_u6_u2_n135 ) , .B1( u1_u6_u2_n140 ) , .A1( u1_u6_u2_n156 ) , .B2( u1_u6_u2_n180 ) , .A2( u1_u6_u2_n188 ) );
  AOI21_X1 u1_u6_u2_U44 (.ZN( u1_u6_u2_n149 ) , .B1( u1_u6_u2_n173 ) , .B2( u1_u6_u2_n188 ) , .A( u1_u6_u2_n95 ) );
  AND3_X1 u1_u6_u2_U45 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n156 ) , .ZN( u1_u6_u2_n95 ) );
  OAI21_X1 u1_u6_u2_U46 (.A( u1_u6_u2_n101 ) , .B2( u1_u6_u2_n121 ) , .B1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n164 ) );
  NAND2_X1 u1_u6_u2_U47 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n155 ) );
  NAND2_X1 u1_u6_u2_U48 (.A2( u1_u6_u2_n105 ) , .A1( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n143 ) );
  NAND2_X1 u1_u6_u2_U49 (.A1( u1_u6_u2_n104 ) , .A2( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n152 ) );
  NOR4_X1 u1_u6_u2_U5 (.A4( u1_u6_u2_n124 ) , .A3( u1_u6_u2_n125 ) , .A2( u1_u6_u2_n126 ) , .A1( u1_u6_u2_n127 ) , .ZN( u1_u6_u2_n128 ) );
  NAND2_X1 u1_u6_u2_U50 (.A1( u1_u6_u2_n100 ) , .A2( u1_u6_u2_n105 ) , .ZN( u1_u6_u2_n132 ) );
  INV_X1 u1_u6_u2_U51 (.A( u1_u6_u2_n140 ) , .ZN( u1_u6_u2_n168 ) );
  INV_X1 u1_u6_u2_U52 (.A( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n167 ) );
  OAI21_X1 u1_u6_u2_U53 (.A( u1_u6_u2_n141 ) , .B2( u1_u6_u2_n142 ) , .ZN( u1_u6_u2_n146 ) , .B1( u1_u6_u2_n153 ) );
  OAI21_X1 u1_u6_u2_U54 (.A( u1_u6_u2_n140 ) , .ZN( u1_u6_u2_n141 ) , .B1( u1_u6_u2_n176 ) , .B2( u1_u6_u2_n177 ) );
  NOR3_X1 u1_u6_u2_U55 (.ZN( u1_u6_u2_n142 ) , .A3( u1_u6_u2_n175 ) , .A2( u1_u6_u2_n178 ) , .A1( u1_u6_u2_n181 ) );
  NAND2_X1 u1_u6_u2_U56 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n113 ) );
  NAND2_X1 u1_u6_u2_U57 (.A1( u1_u6_u2_n106 ) , .A2( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n131 ) );
  NAND2_X1 u1_u6_u2_U58 (.A1( u1_u6_u2_n103 ) , .A2( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n139 ) );
  NAND2_X1 u1_u6_u2_U59 (.A1( u1_u6_u2_n103 ) , .A2( u1_u6_u2_n105 ) , .ZN( u1_u6_u2_n133 ) );
  AOI21_X1 u1_u6_u2_U6 (.B2( u1_u6_u2_n119 ) , .ZN( u1_u6_u2_n127 ) , .A( u1_u6_u2_n137 ) , .B1( u1_u6_u2_n155 ) );
  NAND2_X1 u1_u6_u2_U60 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n103 ) , .ZN( u1_u6_u2_n154 ) );
  NAND2_X1 u1_u6_u2_U61 (.A2( u1_u6_u2_n103 ) , .A1( u1_u6_u2_n104 ) , .ZN( u1_u6_u2_n119 ) );
  NAND2_X1 u1_u6_u2_U62 (.A2( u1_u6_u2_n107 ) , .A1( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n123 ) );
  NAND2_X1 u1_u6_u2_U63 (.A1( u1_u6_u2_n104 ) , .A2( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n122 ) );
  INV_X1 u1_u6_u2_U64 (.A( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n172 ) );
  NAND2_X1 u1_u6_u2_U65 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n102 ) , .ZN( u1_u6_u2_n116 ) );
  NAND2_X1 u1_u6_u2_U66 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n120 ) );
  NAND2_X1 u1_u6_u2_U67 (.A2( u1_u6_u2_n105 ) , .A1( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n117 ) );
  INV_X1 u1_u6_u2_U68 (.ZN( u1_u6_u2_n187 ) , .A( u1_u6_u2_n99 ) );
  OAI21_X1 u1_u6_u2_U69 (.B1( u1_u6_u2_n137 ) , .B2( u1_u6_u2_n143 ) , .A( u1_u6_u2_n98 ) , .ZN( u1_u6_u2_n99 ) );
  AOI21_X1 u1_u6_u2_U7 (.ZN( u1_u6_u2_n124 ) , .B1( u1_u6_u2_n131 ) , .B2( u1_u6_u2_n143 ) , .A( u1_u6_u2_n172 ) );
  NOR2_X1 u1_u6_u2_U70 (.A2( u1_u6_X_16 ) , .ZN( u1_u6_u2_n140 ) , .A1( u1_u6_u2_n166 ) );
  NOR2_X1 u1_u6_u2_U71 (.A2( u1_u6_X_13 ) , .A1( u1_u6_X_14 ) , .ZN( u1_u6_u2_n100 ) );
  NOR2_X1 u1_u6_u2_U72 (.A2( u1_u6_X_16 ) , .A1( u1_u6_X_17 ) , .ZN( u1_u6_u2_n138 ) );
  NOR2_X1 u1_u6_u2_U73 (.A2( u1_u6_X_15 ) , .A1( u1_u6_X_18 ) , .ZN( u1_u6_u2_n104 ) );
  NOR2_X1 u1_u6_u2_U74 (.A2( u1_u6_X_14 ) , .ZN( u1_u6_u2_n103 ) , .A1( u1_u6_u2_n174 ) );
  NOR2_X1 u1_u6_u2_U75 (.A2( u1_u6_X_15 ) , .ZN( u1_u6_u2_n102 ) , .A1( u1_u6_u2_n165 ) );
  NOR2_X1 u1_u6_u2_U76 (.A2( u1_u6_X_17 ) , .ZN( u1_u6_u2_n114 ) , .A1( u1_u6_u2_n169 ) );
  AND2_X1 u1_u6_u2_U77 (.A1( u1_u6_X_15 ) , .ZN( u1_u6_u2_n105 ) , .A2( u1_u6_u2_n165 ) );
  AND2_X1 u1_u6_u2_U78 (.A2( u1_u6_X_15 ) , .A1( u1_u6_X_18 ) , .ZN( u1_u6_u2_n107 ) );
  AND2_X1 u1_u6_u2_U79 (.A1( u1_u6_X_14 ) , .ZN( u1_u6_u2_n106 ) , .A2( u1_u6_u2_n174 ) );
  AOI21_X1 u1_u6_u2_U8 (.B2( u1_u6_u2_n120 ) , .B1( u1_u6_u2_n121 ) , .ZN( u1_u6_u2_n126 ) , .A( u1_u6_u2_n167 ) );
  AND2_X1 u1_u6_u2_U80 (.A1( u1_u6_X_13 ) , .A2( u1_u6_X_14 ) , .ZN( u1_u6_u2_n108 ) );
  INV_X1 u1_u6_u2_U81 (.A( u1_u6_X_16 ) , .ZN( u1_u6_u2_n169 ) );
  INV_X1 u1_u6_u2_U82 (.A( u1_u6_X_17 ) , .ZN( u1_u6_u2_n166 ) );
  INV_X1 u1_u6_u2_U83 (.A( u1_u6_X_13 ) , .ZN( u1_u6_u2_n174 ) );
  INV_X1 u1_u6_u2_U84 (.A( u1_u6_X_18 ) , .ZN( u1_u6_u2_n165 ) );
  NAND4_X1 u1_u6_u2_U85 (.ZN( u1_out6_16 ) , .A4( u1_u6_u2_n128 ) , .A3( u1_u6_u2_n129 ) , .A1( u1_u6_u2_n130 ) , .A2( u1_u6_u2_n186 ) );
  AOI22_X1 u1_u6_u2_U86 (.A2( u1_u6_u2_n118 ) , .ZN( u1_u6_u2_n129 ) , .A1( u1_u6_u2_n140 ) , .B1( u1_u6_u2_n157 ) , .B2( u1_u6_u2_n170 ) );
  INV_X1 u1_u6_u2_U87 (.A( u1_u6_u2_n163 ) , .ZN( u1_u6_u2_n186 ) );
  NAND4_X1 u1_u6_u2_U88 (.ZN( u1_out6_24 ) , .A4( u1_u6_u2_n111 ) , .A3( u1_u6_u2_n112 ) , .A1( u1_u6_u2_n130 ) , .A2( u1_u6_u2_n187 ) );
  AOI221_X1 u1_u6_u2_U89 (.A( u1_u6_u2_n109 ) , .B1( u1_u6_u2_n110 ) , .ZN( u1_u6_u2_n111 ) , .C1( u1_u6_u2_n134 ) , .C2( u1_u6_u2_n170 ) , .B2( u1_u6_u2_n173 ) );
  OAI22_X1 u1_u6_u2_U9 (.ZN( u1_u6_u2_n109 ) , .A2( u1_u6_u2_n113 ) , .B2( u1_u6_u2_n133 ) , .B1( u1_u6_u2_n167 ) , .A1( u1_u6_u2_n168 ) );
  AOI21_X1 u1_u6_u2_U90 (.ZN( u1_u6_u2_n112 ) , .B2( u1_u6_u2_n156 ) , .A( u1_u6_u2_n164 ) , .B1( u1_u6_u2_n181 ) );
  NAND4_X1 u1_u6_u2_U91 (.ZN( u1_out6_30 ) , .A4( u1_u6_u2_n147 ) , .A3( u1_u6_u2_n148 ) , .A2( u1_u6_u2_n149 ) , .A1( u1_u6_u2_n187 ) );
  AOI21_X1 u1_u6_u2_U92 (.B2( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n148 ) , .A( u1_u6_u2_n162 ) , .B1( u1_u6_u2_n182 ) );
  NOR3_X1 u1_u6_u2_U93 (.A3( u1_u6_u2_n144 ) , .A2( u1_u6_u2_n145 ) , .A1( u1_u6_u2_n146 ) , .ZN( u1_u6_u2_n147 ) );
  OR4_X1 u1_u6_u2_U94 (.ZN( u1_out6_6 ) , .A4( u1_u6_u2_n161 ) , .A3( u1_u6_u2_n162 ) , .A2( u1_u6_u2_n163 ) , .A1( u1_u6_u2_n164 ) );
  OR3_X1 u1_u6_u2_U95 (.A2( u1_u6_u2_n159 ) , .A1( u1_u6_u2_n160 ) , .ZN( u1_u6_u2_n161 ) , .A3( u1_u6_u2_n183 ) );
  AOI21_X1 u1_u6_u2_U96 (.B2( u1_u6_u2_n154 ) , .B1( u1_u6_u2_n155 ) , .ZN( u1_u6_u2_n159 ) , .A( u1_u6_u2_n167 ) );
  NAND3_X1 u1_u6_u2_U97 (.A2( u1_u6_u2_n117 ) , .A1( u1_u6_u2_n122 ) , .A3( u1_u6_u2_n123 ) , .ZN( u1_u6_u2_n134 ) );
  NAND3_X1 u1_u6_u2_U98 (.ZN( u1_u6_u2_n110 ) , .A2( u1_u6_u2_n131 ) , .A3( u1_u6_u2_n139 ) , .A1( u1_u6_u2_n154 ) );
  NAND3_X1 u1_u6_u2_U99 (.A2( u1_u6_u2_n100 ) , .ZN( u1_u6_u2_n101 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n114 ) );
  AOI21_X1 u1_u6_u6_U10 (.ZN( u1_u6_u6_n106 ) , .A( u1_u6_u6_n142 ) , .B2( u1_u6_u6_n159 ) , .B1( u1_u6_u6_n164 ) );
  INV_X1 u1_u6_u6_U11 (.A( u1_u6_u6_n155 ) , .ZN( u1_u6_u6_n161 ) );
  INV_X1 u1_u6_u6_U12 (.A( u1_u6_u6_n128 ) , .ZN( u1_u6_u6_n164 ) );
  NAND2_X1 u1_u6_u6_U13 (.ZN( u1_u6_u6_n110 ) , .A1( u1_u6_u6_n122 ) , .A2( u1_u6_u6_n129 ) );
  NAND2_X1 u1_u6_u6_U14 (.ZN( u1_u6_u6_n124 ) , .A2( u1_u6_u6_n146 ) , .A1( u1_u6_u6_n148 ) );
  INV_X1 u1_u6_u6_U15 (.A( u1_u6_u6_n132 ) , .ZN( u1_u6_u6_n171 ) );
  AND2_X1 u1_u6_u6_U16 (.A1( u1_u6_u6_n100 ) , .ZN( u1_u6_u6_n130 ) , .A2( u1_u6_u6_n147 ) );
  INV_X1 u1_u6_u6_U17 (.A( u1_u6_u6_n127 ) , .ZN( u1_u6_u6_n173 ) );
  INV_X1 u1_u6_u6_U18 (.A( u1_u6_u6_n121 ) , .ZN( u1_u6_u6_n167 ) );
  INV_X1 u1_u6_u6_U19 (.A( u1_u6_u6_n100 ) , .ZN( u1_u6_u6_n169 ) );
  INV_X1 u1_u6_u6_U20 (.A( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n170 ) );
  INV_X1 u1_u6_u6_U21 (.A( u1_u6_u6_n113 ) , .ZN( u1_u6_u6_n168 ) );
  AND2_X1 u1_u6_u6_U22 (.A1( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n119 ) , .ZN( u1_u6_u6_n133 ) );
  AND2_X1 u1_u6_u6_U23 (.A2( u1_u6_u6_n121 ) , .A1( u1_u6_u6_n122 ) , .ZN( u1_u6_u6_n131 ) );
  AND3_X1 u1_u6_u6_U24 (.ZN( u1_u6_u6_n120 ) , .A2( u1_u6_u6_n127 ) , .A1( u1_u6_u6_n132 ) , .A3( u1_u6_u6_n145 ) );
  INV_X1 u1_u6_u6_U25 (.A( u1_u6_u6_n146 ) , .ZN( u1_u6_u6_n163 ) );
  AOI222_X1 u1_u6_u6_U26 (.ZN( u1_u6_u6_n114 ) , .A1( u1_u6_u6_n118 ) , .A2( u1_u6_u6_n126 ) , .B2( u1_u6_u6_n151 ) , .C2( u1_u6_u6_n159 ) , .C1( u1_u6_u6_n168 ) , .B1( u1_u6_u6_n169 ) );
  NOR2_X1 u1_u6_u6_U27 (.A1( u1_u6_u6_n162 ) , .A2( u1_u6_u6_n165 ) , .ZN( u1_u6_u6_n98 ) );
  AOI211_X1 u1_u6_u6_U28 (.B( u1_u6_u6_n149 ) , .A( u1_u6_u6_n150 ) , .C2( u1_u6_u6_n151 ) , .C1( u1_u6_u6_n152 ) , .ZN( u1_u6_u6_n153 ) );
  AOI21_X1 u1_u6_u6_U29 (.B2( u1_u6_u6_n147 ) , .B1( u1_u6_u6_n148 ) , .ZN( u1_u6_u6_n149 ) , .A( u1_u6_u6_n158 ) );
  INV_X1 u1_u6_u6_U3 (.A( u1_u6_u6_n110 ) , .ZN( u1_u6_u6_n166 ) );
  AOI21_X1 u1_u6_u6_U30 (.A( u1_u6_u6_n144 ) , .B2( u1_u6_u6_n145 ) , .B1( u1_u6_u6_n146 ) , .ZN( u1_u6_u6_n150 ) );
  NAND2_X1 u1_u6_u6_U31 (.A2( u1_u6_u6_n143 ) , .ZN( u1_u6_u6_n152 ) , .A1( u1_u6_u6_n166 ) );
  NAND2_X1 u1_u6_u6_U32 (.A1( u1_u6_u6_n144 ) , .ZN( u1_u6_u6_n151 ) , .A2( u1_u6_u6_n158 ) );
  NAND2_X1 u1_u6_u6_U33 (.ZN( u1_u6_u6_n132 ) , .A1( u1_u6_u6_n91 ) , .A2( u1_u6_u6_n97 ) );
  AOI22_X1 u1_u6_u6_U34 (.B2( u1_u6_u6_n110 ) , .B1( u1_u6_u6_n111 ) , .A1( u1_u6_u6_n112 ) , .ZN( u1_u6_u6_n115 ) , .A2( u1_u6_u6_n161 ) );
  NAND4_X1 u1_u6_u6_U35 (.A3( u1_u6_u6_n109 ) , .ZN( u1_u6_u6_n112 ) , .A4( u1_u6_u6_n132 ) , .A2( u1_u6_u6_n147 ) , .A1( u1_u6_u6_n166 ) );
  NOR2_X1 u1_u6_u6_U36 (.ZN( u1_u6_u6_n109 ) , .A1( u1_u6_u6_n170 ) , .A2( u1_u6_u6_n173 ) );
  NOR2_X1 u1_u6_u6_U37 (.A2( u1_u6_u6_n126 ) , .ZN( u1_u6_u6_n155 ) , .A1( u1_u6_u6_n160 ) );
  NAND2_X1 u1_u6_u6_U38 (.ZN( u1_u6_u6_n146 ) , .A2( u1_u6_u6_n94 ) , .A1( u1_u6_u6_n99 ) );
  AOI211_X1 u1_u6_u6_U39 (.B( u1_u6_u6_n134 ) , .A( u1_u6_u6_n135 ) , .C1( u1_u6_u6_n136 ) , .ZN( u1_u6_u6_n137 ) , .C2( u1_u6_u6_n151 ) );
  AOI22_X1 u1_u6_u6_U4 (.B2( u1_u6_u6_n101 ) , .A1( u1_u6_u6_n102 ) , .ZN( u1_u6_u6_n103 ) , .B1( u1_u6_u6_n160 ) , .A2( u1_u6_u6_n161 ) );
  NAND4_X1 u1_u6_u6_U40 (.A4( u1_u6_u6_n127 ) , .A3( u1_u6_u6_n128 ) , .A2( u1_u6_u6_n129 ) , .A1( u1_u6_u6_n130 ) , .ZN( u1_u6_u6_n136 ) );
  AOI21_X1 u1_u6_u6_U41 (.B2( u1_u6_u6_n132 ) , .B1( u1_u6_u6_n133 ) , .ZN( u1_u6_u6_n134 ) , .A( u1_u6_u6_n158 ) );
  AOI21_X1 u1_u6_u6_U42 (.B1( u1_u6_u6_n131 ) , .ZN( u1_u6_u6_n135 ) , .A( u1_u6_u6_n144 ) , .B2( u1_u6_u6_n146 ) );
  INV_X1 u1_u6_u6_U43 (.A( u1_u6_u6_n111 ) , .ZN( u1_u6_u6_n158 ) );
  NAND2_X1 u1_u6_u6_U44 (.ZN( u1_u6_u6_n127 ) , .A1( u1_u6_u6_n91 ) , .A2( u1_u6_u6_n92 ) );
  NAND2_X1 u1_u6_u6_U45 (.ZN( u1_u6_u6_n129 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n96 ) );
  INV_X1 u1_u6_u6_U46 (.A( u1_u6_u6_n144 ) , .ZN( u1_u6_u6_n159 ) );
  NAND2_X1 u1_u6_u6_U47 (.ZN( u1_u6_u6_n145 ) , .A2( u1_u6_u6_n97 ) , .A1( u1_u6_u6_n98 ) );
  NAND2_X1 u1_u6_u6_U48 (.ZN( u1_u6_u6_n148 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n94 ) );
  NAND2_X1 u1_u6_u6_U49 (.ZN( u1_u6_u6_n108 ) , .A2( u1_u6_u6_n139 ) , .A1( u1_u6_u6_n144 ) );
  NOR2_X1 u1_u6_u6_U5 (.A1( u1_u6_u6_n118 ) , .ZN( u1_u6_u6_n143 ) , .A2( u1_u6_u6_n168 ) );
  NAND2_X1 u1_u6_u6_U50 (.ZN( u1_u6_u6_n121 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n97 ) );
  NAND2_X1 u1_u6_u6_U51 (.ZN( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n95 ) );
  AND2_X1 u1_u6_u6_U52 (.ZN( u1_u6_u6_n118 ) , .A2( u1_u6_u6_n91 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U53 (.ZN( u1_u6_u6_n147 ) , .A2( u1_u6_u6_n98 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U54 (.ZN( u1_u6_u6_n128 ) , .A1( u1_u6_u6_n94 ) , .A2( u1_u6_u6_n96 ) );
  NAND2_X1 u1_u6_u6_U55 (.ZN( u1_u6_u6_n119 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U56 (.ZN( u1_u6_u6_n123 ) , .A2( u1_u6_u6_n91 ) , .A1( u1_u6_u6_n96 ) );
  NAND2_X1 u1_u6_u6_U57 (.ZN( u1_u6_u6_n100 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n98 ) );
  NAND2_X1 u1_u6_u6_U58 (.ZN( u1_u6_u6_n122 ) , .A1( u1_u6_u6_n94 ) , .A2( u1_u6_u6_n97 ) );
  INV_X1 u1_u6_u6_U59 (.A( u1_u6_u6_n139 ) , .ZN( u1_u6_u6_n160 ) );
  AOI21_X1 u1_u6_u6_U6 (.B1( u1_u6_u6_n107 ) , .B2( u1_u6_u6_n132 ) , .A( u1_u6_u6_n158 ) , .ZN( u1_u6_u6_n88 ) );
  NAND2_X1 u1_u6_u6_U60 (.ZN( u1_u6_u6_n113 ) , .A1( u1_u6_u6_n96 ) , .A2( u1_u6_u6_n98 ) );
  NOR2_X1 u1_u6_u6_U61 (.A2( u1_u6_X_40 ) , .A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n126 ) );
  NOR2_X1 u1_u6_u6_U62 (.A2( u1_u6_X_39 ) , .A1( u1_u6_X_42 ) , .ZN( u1_u6_u6_n92 ) );
  NOR2_X1 u1_u6_u6_U63 (.A2( u1_u6_X_39 ) , .A1( u1_u6_u6_n156 ) , .ZN( u1_u6_u6_n97 ) );
  NOR2_X1 u1_u6_u6_U64 (.A2( u1_u6_X_38 ) , .A1( u1_u6_u6_n165 ) , .ZN( u1_u6_u6_n95 ) );
  NOR2_X1 u1_u6_u6_U65 (.A2( u1_u6_X_41 ) , .ZN( u1_u6_u6_n111 ) , .A1( u1_u6_u6_n157 ) );
  NOR2_X1 u1_u6_u6_U66 (.A2( u1_u6_X_37 ) , .A1( u1_u6_u6_n162 ) , .ZN( u1_u6_u6_n94 ) );
  NOR2_X1 u1_u6_u6_U67 (.A2( u1_u6_X_37 ) , .A1( u1_u6_X_38 ) , .ZN( u1_u6_u6_n91 ) );
  NAND2_X1 u1_u6_u6_U68 (.A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n144 ) , .A2( u1_u6_u6_n157 ) );
  NAND2_X1 u1_u6_u6_U69 (.A2( u1_u6_X_40 ) , .A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n139 ) );
  OAI21_X1 u1_u6_u6_U7 (.A( u1_u6_u6_n159 ) , .B1( u1_u6_u6_n169 ) , .B2( u1_u6_u6_n173 ) , .ZN( u1_u6_u6_n90 ) );
  AND2_X1 u1_u6_u6_U70 (.A1( u1_u6_X_39 ) , .A2( u1_u6_u6_n156 ) , .ZN( u1_u6_u6_n96 ) );
  AND2_X1 u1_u6_u6_U71 (.A1( u1_u6_X_39 ) , .A2( u1_u6_X_42 ) , .ZN( u1_u6_u6_n99 ) );
  INV_X1 u1_u6_u6_U72 (.A( u1_u6_X_40 ) , .ZN( u1_u6_u6_n157 ) );
  INV_X1 u1_u6_u6_U73 (.A( u1_u6_X_37 ) , .ZN( u1_u6_u6_n165 ) );
  INV_X1 u1_u6_u6_U74 (.A( u1_u6_X_38 ) , .ZN( u1_u6_u6_n162 ) );
  INV_X1 u1_u6_u6_U75 (.A( u1_u6_X_42 ) , .ZN( u1_u6_u6_n156 ) );
  NAND4_X1 u1_u6_u6_U76 (.ZN( u1_out6_12 ) , .A4( u1_u6_u6_n114 ) , .A3( u1_u6_u6_n115 ) , .A2( u1_u6_u6_n116 ) , .A1( u1_u6_u6_n117 ) );
  OAI22_X1 u1_u6_u6_U77 (.B2( u1_u6_u6_n111 ) , .ZN( u1_u6_u6_n116 ) , .B1( u1_u6_u6_n126 ) , .A2( u1_u6_u6_n164 ) , .A1( u1_u6_u6_n167 ) );
  OAI21_X1 u1_u6_u6_U78 (.A( u1_u6_u6_n108 ) , .ZN( u1_u6_u6_n117 ) , .B2( u1_u6_u6_n141 ) , .B1( u1_u6_u6_n163 ) );
  NAND4_X1 u1_u6_u6_U79 (.ZN( u1_out6_32 ) , .A4( u1_u6_u6_n103 ) , .A3( u1_u6_u6_n104 ) , .A2( u1_u6_u6_n105 ) , .A1( u1_u6_u6_n106 ) );
  INV_X1 u1_u6_u6_U8 (.ZN( u1_u6_u6_n172 ) , .A( u1_u6_u6_n88 ) );
  AOI22_X1 u1_u6_u6_U80 (.ZN( u1_u6_u6_n104 ) , .A1( u1_u6_u6_n111 ) , .B1( u1_u6_u6_n124 ) , .B2( u1_u6_u6_n151 ) , .A2( u1_u6_u6_n93 ) );
  AOI22_X1 u1_u6_u6_U81 (.ZN( u1_u6_u6_n105 ) , .A2( u1_u6_u6_n108 ) , .A1( u1_u6_u6_n118 ) , .B2( u1_u6_u6_n126 ) , .B1( u1_u6_u6_n171 ) );
  OAI211_X1 u1_u6_u6_U82 (.ZN( u1_out6_22 ) , .B( u1_u6_u6_n137 ) , .A( u1_u6_u6_n138 ) , .C2( u1_u6_u6_n139 ) , .C1( u1_u6_u6_n140 ) );
  AOI22_X1 u1_u6_u6_U83 (.B1( u1_u6_u6_n124 ) , .A2( u1_u6_u6_n125 ) , .A1( u1_u6_u6_n126 ) , .ZN( u1_u6_u6_n138 ) , .B2( u1_u6_u6_n161 ) );
  AND4_X1 u1_u6_u6_U84 (.A3( u1_u6_u6_n119 ) , .A1( u1_u6_u6_n120 ) , .A4( u1_u6_u6_n129 ) , .ZN( u1_u6_u6_n140 ) , .A2( u1_u6_u6_n143 ) );
  OAI211_X1 u1_u6_u6_U85 (.ZN( u1_out6_7 ) , .B( u1_u6_u6_n153 ) , .C2( u1_u6_u6_n154 ) , .C1( u1_u6_u6_n155 ) , .A( u1_u6_u6_n174 ) );
  NOR3_X1 u1_u6_u6_U86 (.A1( u1_u6_u6_n141 ) , .ZN( u1_u6_u6_n154 ) , .A3( u1_u6_u6_n164 ) , .A2( u1_u6_u6_n171 ) );
  INV_X1 u1_u6_u6_U87 (.A( u1_u6_u6_n142 ) , .ZN( u1_u6_u6_n174 ) );
  NAND3_X1 u1_u6_u6_U88 (.A2( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n125 ) , .A1( u1_u6_u6_n130 ) , .A3( u1_u6_u6_n131 ) );
  NAND3_X1 u1_u6_u6_U89 (.A3( u1_u6_u6_n133 ) , .ZN( u1_u6_u6_n141 ) , .A1( u1_u6_u6_n145 ) , .A2( u1_u6_u6_n148 ) );
  AOI22_X1 u1_u6_u6_U9 (.A2( u1_u6_u6_n151 ) , .B2( u1_u6_u6_n161 ) , .A1( u1_u6_u6_n167 ) , .B1( u1_u6_u6_n170 ) , .ZN( u1_u6_u6_n89 ) );
  NAND3_X1 u1_u6_u6_U90 (.ZN( u1_u6_u6_n101 ) , .A3( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n121 ) , .A1( u1_u6_u6_n127 ) );
  NAND3_X1 u1_u6_u6_U91 (.ZN( u1_u6_u6_n102 ) , .A3( u1_u6_u6_n130 ) , .A2( u1_u6_u6_n145 ) , .A1( u1_u6_u6_n166 ) );
  NAND3_X1 u1_u6_u6_U92 (.A3( u1_u6_u6_n113 ) , .A1( u1_u6_u6_n119 ) , .A2( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n93 ) );
  NAND3_X1 u1_u6_u6_U93 (.ZN( u1_u6_u6_n142 ) , .A2( u1_u6_u6_n172 ) , .A3( u1_u6_u6_n89 ) , .A1( u1_u6_u6_n90 ) );
  AND3_X1 u1_u6_u7_U10 (.A3( u1_u6_u7_n110 ) , .A2( u1_u6_u7_n127 ) , .A1( u1_u6_u7_n132 ) , .ZN( u1_u6_u7_n92 ) );
  OAI21_X1 u1_u6_u7_U11 (.A( u1_u6_u7_n161 ) , .B1( u1_u6_u7_n168 ) , .B2( u1_u6_u7_n173 ) , .ZN( u1_u6_u7_n91 ) );
  AOI211_X1 u1_u6_u7_U12 (.A( u1_u6_u7_n117 ) , .ZN( u1_u6_u7_n118 ) , .C2( u1_u6_u7_n126 ) , .C1( u1_u6_u7_n177 ) , .B( u1_u6_u7_n180 ) );
  OAI22_X1 u1_u6_u7_U13 (.B1( u1_u6_u7_n115 ) , .ZN( u1_u6_u7_n117 ) , .A2( u1_u6_u7_n133 ) , .A1( u1_u6_u7_n137 ) , .B2( u1_u6_u7_n162 ) );
  INV_X1 u1_u6_u7_U14 (.A( u1_u6_u7_n116 ) , .ZN( u1_u6_u7_n180 ) );
  NOR3_X1 u1_u6_u7_U15 (.ZN( u1_u6_u7_n115 ) , .A3( u1_u6_u7_n145 ) , .A2( u1_u6_u7_n168 ) , .A1( u1_u6_u7_n169 ) );
  OAI211_X1 u1_u6_u7_U16 (.B( u1_u6_u7_n122 ) , .A( u1_u6_u7_n123 ) , .C2( u1_u6_u7_n124 ) , .ZN( u1_u6_u7_n154 ) , .C1( u1_u6_u7_n162 ) );
  AOI222_X1 u1_u6_u7_U17 (.ZN( u1_u6_u7_n122 ) , .C2( u1_u6_u7_n126 ) , .C1( u1_u6_u7_n145 ) , .B1( u1_u6_u7_n161 ) , .A2( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n170 ) , .A1( u1_u6_u7_n176 ) );
  INV_X1 u1_u6_u7_U18 (.A( u1_u6_u7_n133 ) , .ZN( u1_u6_u7_n176 ) );
  NOR3_X1 u1_u6_u7_U19 (.A2( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n135 ) , .ZN( u1_u6_u7_n136 ) , .A3( u1_u6_u7_n171 ) );
  NOR2_X1 u1_u6_u7_U20 (.A1( u1_u6_u7_n130 ) , .A2( u1_u6_u7_n134 ) , .ZN( u1_u6_u7_n153 ) );
  INV_X1 u1_u6_u7_U21 (.A( u1_u6_u7_n101 ) , .ZN( u1_u6_u7_n165 ) );
  NOR2_X1 u1_u6_u7_U22 (.ZN( u1_u6_u7_n111 ) , .A2( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n169 ) );
  AOI21_X1 u1_u6_u7_U23 (.ZN( u1_u6_u7_n104 ) , .B2( u1_u6_u7_n112 ) , .B1( u1_u6_u7_n127 ) , .A( u1_u6_u7_n164 ) );
  AOI21_X1 u1_u6_u7_U24 (.ZN( u1_u6_u7_n106 ) , .B1( u1_u6_u7_n133 ) , .B2( u1_u6_u7_n146 ) , .A( u1_u6_u7_n162 ) );
  AOI21_X1 u1_u6_u7_U25 (.A( u1_u6_u7_n101 ) , .ZN( u1_u6_u7_n107 ) , .B2( u1_u6_u7_n128 ) , .B1( u1_u6_u7_n175 ) );
  INV_X1 u1_u6_u7_U26 (.A( u1_u6_u7_n138 ) , .ZN( u1_u6_u7_n171 ) );
  INV_X1 u1_u6_u7_U27 (.A( u1_u6_u7_n131 ) , .ZN( u1_u6_u7_n177 ) );
  INV_X1 u1_u6_u7_U28 (.A( u1_u6_u7_n110 ) , .ZN( u1_u6_u7_n174 ) );
  NAND2_X1 u1_u6_u7_U29 (.A1( u1_u6_u7_n129 ) , .A2( u1_u6_u7_n132 ) , .ZN( u1_u6_u7_n149 ) );
  OAI21_X1 u1_u6_u7_U3 (.ZN( u1_u6_u7_n159 ) , .A( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n171 ) , .B1( u1_u6_u7_n174 ) );
  NAND2_X1 u1_u6_u7_U30 (.A1( u1_u6_u7_n113 ) , .A2( u1_u6_u7_n124 ) , .ZN( u1_u6_u7_n130 ) );
  INV_X1 u1_u6_u7_U31 (.A( u1_u6_u7_n112 ) , .ZN( u1_u6_u7_n173 ) );
  INV_X1 u1_u6_u7_U32 (.A( u1_u6_u7_n128 ) , .ZN( u1_u6_u7_n168 ) );
  INV_X1 u1_u6_u7_U33 (.A( u1_u6_u7_n148 ) , .ZN( u1_u6_u7_n169 ) );
  INV_X1 u1_u6_u7_U34 (.A( u1_u6_u7_n127 ) , .ZN( u1_u6_u7_n179 ) );
  NOR2_X1 u1_u6_u7_U35 (.ZN( u1_u6_u7_n101 ) , .A2( u1_u6_u7_n150 ) , .A1( u1_u6_u7_n156 ) );
  AOI211_X1 u1_u6_u7_U36 (.B( u1_u6_u7_n154 ) , .A( u1_u6_u7_n155 ) , .C1( u1_u6_u7_n156 ) , .ZN( u1_u6_u7_n157 ) , .C2( u1_u6_u7_n172 ) );
  INV_X1 u1_u6_u7_U37 (.A( u1_u6_u7_n153 ) , .ZN( u1_u6_u7_n172 ) );
  AOI211_X1 u1_u6_u7_U38 (.B( u1_u6_u7_n139 ) , .A( u1_u6_u7_n140 ) , .C2( u1_u6_u7_n141 ) , .ZN( u1_u6_u7_n142 ) , .C1( u1_u6_u7_n156 ) );
  NAND4_X1 u1_u6_u7_U39 (.A3( u1_u6_u7_n127 ) , .A2( u1_u6_u7_n128 ) , .A1( u1_u6_u7_n129 ) , .ZN( u1_u6_u7_n141 ) , .A4( u1_u6_u7_n147 ) );
  INV_X1 u1_u6_u7_U4 (.A( u1_u6_u7_n111 ) , .ZN( u1_u6_u7_n170 ) );
  AOI21_X1 u1_u6_u7_U40 (.A( u1_u6_u7_n137 ) , .B1( u1_u6_u7_n138 ) , .ZN( u1_u6_u7_n139 ) , .B2( u1_u6_u7_n146 ) );
  OAI22_X1 u1_u6_u7_U41 (.B1( u1_u6_u7_n136 ) , .ZN( u1_u6_u7_n140 ) , .A1( u1_u6_u7_n153 ) , .B2( u1_u6_u7_n162 ) , .A2( u1_u6_u7_n164 ) );
  AOI21_X1 u1_u6_u7_U42 (.ZN( u1_u6_u7_n123 ) , .B1( u1_u6_u7_n165 ) , .B2( u1_u6_u7_n177 ) , .A( u1_u6_u7_n97 ) );
  AOI21_X1 u1_u6_u7_U43 (.B2( u1_u6_u7_n113 ) , .B1( u1_u6_u7_n124 ) , .A( u1_u6_u7_n125 ) , .ZN( u1_u6_u7_n97 ) );
  INV_X1 u1_u6_u7_U44 (.A( u1_u6_u7_n125 ) , .ZN( u1_u6_u7_n161 ) );
  INV_X1 u1_u6_u7_U45 (.A( u1_u6_u7_n152 ) , .ZN( u1_u6_u7_n162 ) );
  AOI22_X1 u1_u6_u7_U46 (.A2( u1_u6_u7_n114 ) , .ZN( u1_u6_u7_n119 ) , .B1( u1_u6_u7_n130 ) , .A1( u1_u6_u7_n156 ) , .B2( u1_u6_u7_n165 ) );
  NAND2_X1 u1_u6_u7_U47 (.A2( u1_u6_u7_n112 ) , .ZN( u1_u6_u7_n114 ) , .A1( u1_u6_u7_n175 ) );
  AND2_X1 u1_u6_u7_U48 (.ZN( u1_u6_u7_n145 ) , .A2( u1_u6_u7_n98 ) , .A1( u1_u6_u7_n99 ) );
  NOR2_X1 u1_u6_u7_U49 (.ZN( u1_u6_u7_n137 ) , .A1( u1_u6_u7_n150 ) , .A2( u1_u6_u7_n161 ) );
  INV_X1 u1_u6_u7_U5 (.A( u1_u6_u7_n149 ) , .ZN( u1_u6_u7_n175 ) );
  AOI21_X1 u1_u6_u7_U50 (.ZN( u1_u6_u7_n105 ) , .B2( u1_u6_u7_n110 ) , .A( u1_u6_u7_n125 ) , .B1( u1_u6_u7_n147 ) );
  NAND2_X1 u1_u6_u7_U51 (.ZN( u1_u6_u7_n146 ) , .A1( u1_u6_u7_n95 ) , .A2( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U52 (.A2( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n147 ) , .A1( u1_u6_u7_n93 ) );
  NAND2_X1 u1_u6_u7_U53 (.A1( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n127 ) , .A2( u1_u6_u7_n99 ) );
  OR2_X1 u1_u6_u7_U54 (.ZN( u1_u6_u7_n126 ) , .A2( u1_u6_u7_n152 ) , .A1( u1_u6_u7_n156 ) );
  NAND2_X1 u1_u6_u7_U55 (.A2( u1_u6_u7_n102 ) , .A1( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n133 ) );
  NAND2_X1 u1_u6_u7_U56 (.ZN( u1_u6_u7_n112 ) , .A2( u1_u6_u7_n96 ) , .A1( u1_u6_u7_n99 ) );
  NAND2_X1 u1_u6_u7_U57 (.A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n128 ) , .A1( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U58 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n113 ) , .A2( u1_u6_u7_n93 ) );
  NAND2_X1 u1_u6_u7_U59 (.A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n124 ) , .A1( u1_u6_u7_n96 ) );
  INV_X1 u1_u6_u7_U6 (.A( u1_u6_u7_n154 ) , .ZN( u1_u6_u7_n178 ) );
  NAND2_X1 u1_u6_u7_U60 (.ZN( u1_u6_u7_n110 ) , .A1( u1_u6_u7_n95 ) , .A2( u1_u6_u7_n96 ) );
  INV_X1 u1_u6_u7_U61 (.A( u1_u6_u7_n150 ) , .ZN( u1_u6_u7_n164 ) );
  AND2_X1 u1_u6_u7_U62 (.ZN( u1_u6_u7_n134 ) , .A1( u1_u6_u7_n93 ) , .A2( u1_u6_u7_n98 ) );
  NAND2_X1 u1_u6_u7_U63 (.A1( u1_u6_u7_n100 ) , .A2( u1_u6_u7_n102 ) , .ZN( u1_u6_u7_n129 ) );
  NAND2_X1 u1_u6_u7_U64 (.A2( u1_u6_u7_n103 ) , .ZN( u1_u6_u7_n131 ) , .A1( u1_u6_u7_n95 ) );
  NAND2_X1 u1_u6_u7_U65 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n138 ) , .A2( u1_u6_u7_n99 ) );
  NAND2_X1 u1_u6_u7_U66 (.ZN( u1_u6_u7_n132 ) , .A1( u1_u6_u7_n93 ) , .A2( u1_u6_u7_n96 ) );
  NAND2_X1 u1_u6_u7_U67 (.A1( u1_u6_u7_n100 ) , .ZN( u1_u6_u7_n148 ) , .A2( u1_u6_u7_n95 ) );
  NOR2_X1 u1_u6_u7_U68 (.A2( u1_u6_X_47 ) , .ZN( u1_u6_u7_n150 ) , .A1( u1_u6_u7_n163 ) );
  NOR2_X1 u1_u6_u7_U69 (.A2( u1_u6_X_43 ) , .A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n103 ) );
  AOI211_X1 u1_u6_u7_U7 (.ZN( u1_u6_u7_n116 ) , .A( u1_u6_u7_n155 ) , .C1( u1_u6_u7_n161 ) , .C2( u1_u6_u7_n171 ) , .B( u1_u6_u7_n94 ) );
  NOR2_X1 u1_u6_u7_U70 (.A2( u1_u6_X_48 ) , .A1( u1_u6_u7_n166 ) , .ZN( u1_u6_u7_n95 ) );
  NOR2_X1 u1_u6_u7_U71 (.A2( u1_u6_X_45 ) , .A1( u1_u6_X_48 ) , .ZN( u1_u6_u7_n99 ) );
  NOR2_X1 u1_u6_u7_U72 (.A2( u1_u6_X_44 ) , .A1( u1_u6_u7_n167 ) , .ZN( u1_u6_u7_n98 ) );
  NOR2_X1 u1_u6_u7_U73 (.A2( u1_u6_X_46 ) , .A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n152 ) );
  AND2_X1 u1_u6_u7_U74 (.A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n156 ) , .A2( u1_u6_u7_n163 ) );
  NAND2_X1 u1_u6_u7_U75 (.A2( u1_u6_X_46 ) , .A1( u1_u6_X_47 ) , .ZN( u1_u6_u7_n125 ) );
  AND2_X1 u1_u6_u7_U76 (.A2( u1_u6_X_45 ) , .A1( u1_u6_X_48 ) , .ZN( u1_u6_u7_n102 ) );
  AND2_X1 u1_u6_u7_U77 (.A2( u1_u6_X_43 ) , .A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n96 ) );
  AND2_X1 u1_u6_u7_U78 (.A1( u1_u6_X_44 ) , .ZN( u1_u6_u7_n100 ) , .A2( u1_u6_u7_n167 ) );
  AND2_X1 u1_u6_u7_U79 (.A1( u1_u6_X_48 ) , .A2( u1_u6_u7_n166 ) , .ZN( u1_u6_u7_n93 ) );
  OAI222_X1 u1_u6_u7_U8 (.C2( u1_u6_u7_n101 ) , .B2( u1_u6_u7_n111 ) , .A1( u1_u6_u7_n113 ) , .C1( u1_u6_u7_n146 ) , .A2( u1_u6_u7_n162 ) , .B1( u1_u6_u7_n164 ) , .ZN( u1_u6_u7_n94 ) );
  INV_X1 u1_u6_u7_U80 (.A( u1_u6_X_46 ) , .ZN( u1_u6_u7_n163 ) );
  INV_X1 u1_u6_u7_U81 (.A( u1_u6_X_43 ) , .ZN( u1_u6_u7_n167 ) );
  INV_X1 u1_u6_u7_U82 (.A( u1_u6_X_45 ) , .ZN( u1_u6_u7_n166 ) );
  NAND4_X1 u1_u6_u7_U83 (.ZN( u1_out6_5 ) , .A4( u1_u6_u7_n108 ) , .A3( u1_u6_u7_n109 ) , .A1( u1_u6_u7_n116 ) , .A2( u1_u6_u7_n123 ) );
  AOI22_X1 u1_u6_u7_U84 (.ZN( u1_u6_u7_n109 ) , .A2( u1_u6_u7_n126 ) , .B2( u1_u6_u7_n145 ) , .B1( u1_u6_u7_n156 ) , .A1( u1_u6_u7_n171 ) );
  NOR4_X1 u1_u6_u7_U85 (.A4( u1_u6_u7_n104 ) , .A3( u1_u6_u7_n105 ) , .A2( u1_u6_u7_n106 ) , .A1( u1_u6_u7_n107 ) , .ZN( u1_u6_u7_n108 ) );
  NAND4_X1 u1_u6_u7_U86 (.ZN( u1_out6_21 ) , .A4( u1_u6_u7_n157 ) , .A3( u1_u6_u7_n158 ) , .A2( u1_u6_u7_n159 ) , .A1( u1_u6_u7_n160 ) );
  OAI21_X1 u1_u6_u7_U87 (.B1( u1_u6_u7_n145 ) , .ZN( u1_u6_u7_n160 ) , .A( u1_u6_u7_n161 ) , .B2( u1_u6_u7_n177 ) );
  AOI22_X1 u1_u6_u7_U88 (.B2( u1_u6_u7_n149 ) , .B1( u1_u6_u7_n150 ) , .A2( u1_u6_u7_n151 ) , .A1( u1_u6_u7_n152 ) , .ZN( u1_u6_u7_n158 ) );
  NAND4_X1 u1_u6_u7_U89 (.ZN( u1_out6_15 ) , .A4( u1_u6_u7_n142 ) , .A3( u1_u6_u7_n143 ) , .A2( u1_u6_u7_n144 ) , .A1( u1_u6_u7_n178 ) );
  OAI221_X1 u1_u6_u7_U9 (.C1( u1_u6_u7_n101 ) , .C2( u1_u6_u7_n147 ) , .ZN( u1_u6_u7_n155 ) , .B2( u1_u6_u7_n162 ) , .A( u1_u6_u7_n91 ) , .B1( u1_u6_u7_n92 ) );
  OR2_X1 u1_u6_u7_U90 (.A2( u1_u6_u7_n125 ) , .A1( u1_u6_u7_n129 ) , .ZN( u1_u6_u7_n144 ) );
  AOI22_X1 u1_u6_u7_U91 (.A2( u1_u6_u7_n126 ) , .ZN( u1_u6_u7_n143 ) , .B2( u1_u6_u7_n165 ) , .B1( u1_u6_u7_n173 ) , .A1( u1_u6_u7_n174 ) );
  NAND4_X1 u1_u6_u7_U92 (.ZN( u1_out6_27 ) , .A4( u1_u6_u7_n118 ) , .A3( u1_u6_u7_n119 ) , .A2( u1_u6_u7_n120 ) , .A1( u1_u6_u7_n121 ) );
  OAI21_X1 u1_u6_u7_U93 (.ZN( u1_u6_u7_n121 ) , .B2( u1_u6_u7_n145 ) , .A( u1_u6_u7_n150 ) , .B1( u1_u6_u7_n174 ) );
  OAI21_X1 u1_u6_u7_U94 (.ZN( u1_u6_u7_n120 ) , .A( u1_u6_u7_n161 ) , .B2( u1_u6_u7_n170 ) , .B1( u1_u6_u7_n179 ) );
  NAND3_X1 u1_u6_u7_U95 (.A3( u1_u6_u7_n146 ) , .A2( u1_u6_u7_n147 ) , .A1( u1_u6_u7_n148 ) , .ZN( u1_u6_u7_n151 ) );
  NAND3_X1 u1_u6_u7_U96 (.A3( u1_u6_u7_n131 ) , .A2( u1_u6_u7_n132 ) , .A1( u1_u6_u7_n133 ) , .ZN( u1_u6_u7_n135 ) );
  XOR2_X1 u1_u8_U11 (.B( u1_K9_44 ) , .A( u1_R7_29 ) , .Z( u1_u8_X_44 ) );
  XOR2_X1 u1_u8_U12 (.B( u1_K9_43 ) , .A( u1_R7_28 ) , .Z( u1_u8_X_43 ) );
  XOR2_X1 u1_u8_U13 (.B( u1_K9_42 ) , .A( u1_R7_29 ) , .Z( u1_u8_X_42 ) );
  XOR2_X1 u1_u8_U14 (.B( u1_K9_41 ) , .A( u1_R7_28 ) , .Z( u1_u8_X_41 ) );
  XOR2_X1 u1_u8_U18 (.B( u1_K9_38 ) , .A( u1_R7_25 ) , .Z( u1_u8_X_38 ) );
  XOR2_X1 u1_u8_U19 (.B( u1_K9_37 ) , .A( u1_R7_24 ) , .Z( u1_u8_X_37 ) );
  XOR2_X1 u1_u8_U20 (.B( u1_K9_36 ) , .A( u1_R7_25 ) , .Z( u1_u8_X_36 ) );
  XOR2_X1 u1_u8_U21 (.B( u1_K9_35 ) , .A( u1_R7_24 ) , .Z( u1_u8_X_35 ) );
  XOR2_X1 u1_u8_U25 (.B( u1_K9_31 ) , .A( u1_R7_20 ) , .Z( u1_u8_X_31 ) );
  XOR2_X1 u1_u8_U27 (.B( u1_K9_2 ) , .A( u1_R7_1 ) , .Z( u1_u8_X_2 ) );
  XOR2_X1 u1_u8_U28 (.B( u1_K9_29 ) , .A( u1_R7_20 ) , .Z( u1_u8_X_29 ) );
  XOR2_X1 u1_u8_U30 (.B( u1_K9_27 ) , .A( u1_R7_18 ) , .Z( u1_u8_X_27 ) );
  XOR2_X1 u1_u8_U31 (.B( u1_K9_26 ) , .A( u1_R7_17 ) , .Z( u1_u8_X_26 ) );
  XOR2_X1 u1_u8_U32 (.B( u1_K9_25 ) , .A( u1_R7_16 ) , .Z( u1_u8_X_25 ) );
  XOR2_X1 u1_u8_U33 (.B( u1_K9_24 ) , .A( u1_R7_17 ) , .Z( u1_u8_X_24 ) );
  XOR2_X1 u1_u8_U34 (.B( u1_K9_23 ) , .A( u1_R7_16 ) , .Z( u1_u8_X_23 ) );
  XOR2_X1 u1_u8_U35 (.B( u1_K9_22 ) , .A( u1_R7_15 ) , .Z( u1_u8_X_22 ) );
  XOR2_X1 u1_u8_U37 (.B( u1_K9_20 ) , .A( u1_R7_13 ) , .Z( u1_u8_X_20 ) );
  XOR2_X1 u1_u8_U38 (.B( u1_K9_1 ) , .A( u1_R7_32 ) , .Z( u1_u8_X_1 ) );
  XOR2_X1 u1_u8_U39 (.B( u1_K9_19 ) , .A( u1_R7_12 ) , .Z( u1_u8_X_19 ) );
  XOR2_X1 u1_u8_U4 (.B( u1_K9_6 ) , .A( u1_R7_5 ) , .Z( u1_u8_X_6 ) );
  XOR2_X1 u1_u8_U5 (.B( u1_K9_5 ) , .A( u1_R7_4 ) , .Z( u1_u8_X_5 ) );
  XOR2_X1 u1_u8_U7 (.B( u1_K9_48 ) , .A( u1_R7_1 ) , .Z( u1_u8_X_48 ) );
  XOR2_X1 u1_u8_U8 (.B( u1_K9_47 ) , .A( u1_R7_32 ) , .Z( u1_u8_X_47 ) );
  AND2_X1 u1_u8_u0_U10 (.A1( u1_u8_u0_n131 ) , .ZN( u1_u8_u0_n141 ) , .A2( u1_u8_u0_n150 ) );
  AND3_X1 u1_u8_u0_U11 (.A2( u1_u8_u0_n112 ) , .ZN( u1_u8_u0_n127 ) , .A3( u1_u8_u0_n130 ) , .A1( u1_u8_u0_n148 ) );
  AND2_X1 u1_u8_u0_U12 (.ZN( u1_u8_u0_n107 ) , .A1( u1_u8_u0_n130 ) , .A2( u1_u8_u0_n140 ) );
  AND2_X1 u1_u8_u0_U13 (.A2( u1_u8_u0_n129 ) , .A1( u1_u8_u0_n130 ) , .ZN( u1_u8_u0_n151 ) );
  AND2_X1 u1_u8_u0_U14 (.A1( u1_u8_u0_n108 ) , .A2( u1_u8_u0_n125 ) , .ZN( u1_u8_u0_n145 ) );
  INV_X1 u1_u8_u0_U15 (.A( u1_u8_u0_n143 ) , .ZN( u1_u8_u0_n173 ) );
  NOR2_X1 u1_u8_u0_U16 (.A2( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n147 ) , .A1( u1_u8_u0_n160 ) );
  AOI21_X1 u1_u8_u0_U17 (.B1( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n132 ) , .A( u1_u8_u0_n165 ) , .B2( u1_u8_u0_n93 ) );
  OAI22_X1 u1_u8_u0_U18 (.B1( u1_u8_u0_n131 ) , .A1( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n147 ) , .A2( u1_u8_u0_n90 ) , .ZN( u1_u8_u0_n91 ) );
  AND3_X1 u1_u8_u0_U19 (.A3( u1_u8_u0_n121 ) , .A2( u1_u8_u0_n125 ) , .A1( u1_u8_u0_n148 ) , .ZN( u1_u8_u0_n90 ) );
  OAI22_X1 u1_u8_u0_U20 (.B1( u1_u8_u0_n125 ) , .ZN( u1_u8_u0_n126 ) , .A1( u1_u8_u0_n138 ) , .A2( u1_u8_u0_n146 ) , .B2( u1_u8_u0_n147 ) );
  NOR2_X1 u1_u8_u0_U21 (.A1( u1_u8_u0_n163 ) , .A2( u1_u8_u0_n164 ) , .ZN( u1_u8_u0_n95 ) );
  AOI22_X1 u1_u8_u0_U22 (.B2( u1_u8_u0_n109 ) , .A2( u1_u8_u0_n110 ) , .ZN( u1_u8_u0_n111 ) , .B1( u1_u8_u0_n118 ) , .A1( u1_u8_u0_n160 ) );
  NAND2_X1 u1_u8_u0_U23 (.A2( u1_u8_u0_n102 ) , .A1( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n149 ) );
  INV_X1 u1_u8_u0_U24 (.A( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n161 ) );
  INV_X1 u1_u8_u0_U25 (.A( u1_u8_u0_n118 ) , .ZN( u1_u8_u0_n158 ) );
  NAND2_X1 u1_u8_u0_U26 (.A2( u1_u8_u0_n100 ) , .ZN( u1_u8_u0_n131 ) , .A1( u1_u8_u0_n92 ) );
  NAND2_X1 u1_u8_u0_U27 (.ZN( u1_u8_u0_n108 ) , .A1( u1_u8_u0_n92 ) , .A2( u1_u8_u0_n94 ) );
  AOI21_X1 u1_u8_u0_U28 (.ZN( u1_u8_u0_n104 ) , .B1( u1_u8_u0_n107 ) , .B2( u1_u8_u0_n141 ) , .A( u1_u8_u0_n144 ) );
  AOI21_X1 u1_u8_u0_U29 (.B1( u1_u8_u0_n127 ) , .B2( u1_u8_u0_n129 ) , .A( u1_u8_u0_n138 ) , .ZN( u1_u8_u0_n96 ) );
  INV_X1 u1_u8_u0_U3 (.A( u1_u8_u0_n113 ) , .ZN( u1_u8_u0_n166 ) );
  NAND2_X1 u1_u8_u0_U30 (.A2( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n114 ) , .A1( u1_u8_u0_n92 ) );
  NOR2_X1 u1_u8_u0_U31 (.A1( u1_u8_u0_n120 ) , .ZN( u1_u8_u0_n143 ) , .A2( u1_u8_u0_n167 ) );
  OAI221_X1 u1_u8_u0_U32 (.C1( u1_u8_u0_n112 ) , .ZN( u1_u8_u0_n120 ) , .B1( u1_u8_u0_n138 ) , .B2( u1_u8_u0_n141 ) , .C2( u1_u8_u0_n147 ) , .A( u1_u8_u0_n172 ) );
  AOI211_X1 u1_u8_u0_U33 (.B( u1_u8_u0_n115 ) , .A( u1_u8_u0_n116 ) , .C2( u1_u8_u0_n117 ) , .C1( u1_u8_u0_n118 ) , .ZN( u1_u8_u0_n119 ) );
  NAND2_X1 u1_u8_u0_U34 (.A2( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n140 ) , .A1( u1_u8_u0_n94 ) );
  NAND2_X1 u1_u8_u0_U35 (.A1( u1_u8_u0_n100 ) , .A2( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n125 ) );
  NAND2_X1 u1_u8_u0_U36 (.A1( u1_u8_u0_n101 ) , .A2( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n150 ) );
  INV_X1 u1_u8_u0_U37 (.A( u1_u8_u0_n138 ) , .ZN( u1_u8_u0_n160 ) );
  NAND2_X1 u1_u8_u0_U38 (.A2( u1_u8_u0_n100 ) , .A1( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n139 ) );
  NAND2_X1 u1_u8_u0_U39 (.ZN( u1_u8_u0_n112 ) , .A2( u1_u8_u0_n92 ) , .A1( u1_u8_u0_n93 ) );
  AOI21_X1 u1_u8_u0_U4 (.B1( u1_u8_u0_n114 ) , .ZN( u1_u8_u0_n115 ) , .B2( u1_u8_u0_n129 ) , .A( u1_u8_u0_n161 ) );
  NAND2_X1 u1_u8_u0_U40 (.A1( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n130 ) , .A2( u1_u8_u0_n94 ) );
  INV_X1 u1_u8_u0_U41 (.ZN( u1_u8_u0_n172 ) , .A( u1_u8_u0_n88 ) );
  OAI222_X1 u1_u8_u0_U42 (.C1( u1_u8_u0_n108 ) , .A1( u1_u8_u0_n125 ) , .B2( u1_u8_u0_n128 ) , .B1( u1_u8_u0_n144 ) , .A2( u1_u8_u0_n158 ) , .C2( u1_u8_u0_n161 ) , .ZN( u1_u8_u0_n88 ) );
  NAND2_X1 u1_u8_u0_U43 (.A2( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n121 ) , .A1( u1_u8_u0_n93 ) );
  OR3_X1 u1_u8_u0_U44 (.A3( u1_u8_u0_n152 ) , .A2( u1_u8_u0_n153 ) , .A1( u1_u8_u0_n154 ) , .ZN( u1_u8_u0_n155 ) );
  AOI21_X1 u1_u8_u0_U45 (.A( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n145 ) , .B1( u1_u8_u0_n146 ) , .ZN( u1_u8_u0_n154 ) );
  AOI21_X1 u1_u8_u0_U46 (.B2( u1_u8_u0_n150 ) , .B1( u1_u8_u0_n151 ) , .ZN( u1_u8_u0_n152 ) , .A( u1_u8_u0_n158 ) );
  AOI21_X1 u1_u8_u0_U47 (.A( u1_u8_u0_n147 ) , .B2( u1_u8_u0_n148 ) , .B1( u1_u8_u0_n149 ) , .ZN( u1_u8_u0_n153 ) );
  INV_X1 u1_u8_u0_U48 (.ZN( u1_u8_u0_n171 ) , .A( u1_u8_u0_n99 ) );
  OAI211_X1 u1_u8_u0_U49 (.C2( u1_u8_u0_n140 ) , .C1( u1_u8_u0_n161 ) , .A( u1_u8_u0_n169 ) , .B( u1_u8_u0_n98 ) , .ZN( u1_u8_u0_n99 ) );
  AOI21_X1 u1_u8_u0_U5 (.B2( u1_u8_u0_n131 ) , .ZN( u1_u8_u0_n134 ) , .B1( u1_u8_u0_n151 ) , .A( u1_u8_u0_n158 ) );
  INV_X1 u1_u8_u0_U50 (.ZN( u1_u8_u0_n169 ) , .A( u1_u8_u0_n91 ) );
  AOI211_X1 u1_u8_u0_U51 (.C1( u1_u8_u0_n118 ) , .A( u1_u8_u0_n123 ) , .B( u1_u8_u0_n96 ) , .C2( u1_u8_u0_n97 ) , .ZN( u1_u8_u0_n98 ) );
  NOR2_X1 u1_u8_u0_U52 (.A2( u1_u8_X_4 ) , .A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n118 ) );
  NOR2_X1 u1_u8_u0_U53 (.A2( u1_u8_X_1 ) , .ZN( u1_u8_u0_n101 ) , .A1( u1_u8_u0_n163 ) );
  NOR2_X1 u1_u8_u0_U54 (.A2( u1_u8_X_3 ) , .A1( u1_u8_X_6 ) , .ZN( u1_u8_u0_n94 ) );
  NOR2_X1 u1_u8_u0_U55 (.A2( u1_u8_X_6 ) , .ZN( u1_u8_u0_n100 ) , .A1( u1_u8_u0_n162 ) );
  NAND2_X1 u1_u8_u0_U56 (.A2( u1_u8_X_4 ) , .A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n144 ) );
  NOR2_X1 u1_u8_u0_U57 (.A2( u1_u8_X_5 ) , .ZN( u1_u8_u0_n136 ) , .A1( u1_u8_u0_n159 ) );
  NAND2_X1 u1_u8_u0_U58 (.A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n138 ) , .A2( u1_u8_u0_n159 ) );
  AND2_X1 u1_u8_u0_U59 (.A2( u1_u8_X_3 ) , .A1( u1_u8_X_6 ) , .ZN( u1_u8_u0_n102 ) );
  NOR2_X1 u1_u8_u0_U6 (.A1( u1_u8_u0_n108 ) , .ZN( u1_u8_u0_n123 ) , .A2( u1_u8_u0_n158 ) );
  AND2_X1 u1_u8_u0_U60 (.A1( u1_u8_X_6 ) , .A2( u1_u8_u0_n162 ) , .ZN( u1_u8_u0_n93 ) );
  INV_X1 u1_u8_u0_U61 (.A( u1_u8_X_4 ) , .ZN( u1_u8_u0_n159 ) );
  INV_X1 u1_u8_u0_U62 (.A( u1_u8_X_1 ) , .ZN( u1_u8_u0_n164 ) );
  INV_X1 u1_u8_u0_U63 (.A( u1_u8_X_3 ) , .ZN( u1_u8_u0_n162 ) );
  INV_X1 u1_u8_u0_U64 (.A( u1_u8_u0_n126 ) , .ZN( u1_u8_u0_n168 ) );
  AOI211_X1 u1_u8_u0_U65 (.B( u1_u8_u0_n133 ) , .A( u1_u8_u0_n134 ) , .C2( u1_u8_u0_n135 ) , .C1( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n137 ) );
  OR4_X1 u1_u8_u0_U66 (.ZN( u1_out8_17 ) , .A4( u1_u8_u0_n122 ) , .A2( u1_u8_u0_n123 ) , .A1( u1_u8_u0_n124 ) , .A3( u1_u8_u0_n170 ) );
  AOI21_X1 u1_u8_u0_U67 (.B2( u1_u8_u0_n107 ) , .ZN( u1_u8_u0_n124 ) , .B1( u1_u8_u0_n128 ) , .A( u1_u8_u0_n161 ) );
  INV_X1 u1_u8_u0_U68 (.A( u1_u8_u0_n111 ) , .ZN( u1_u8_u0_n170 ) );
  OR4_X1 u1_u8_u0_U69 (.ZN( u1_out8_31 ) , .A4( u1_u8_u0_n155 ) , .A2( u1_u8_u0_n156 ) , .A1( u1_u8_u0_n157 ) , .A3( u1_u8_u0_n173 ) );
  OAI21_X1 u1_u8_u0_U7 (.B1( u1_u8_u0_n150 ) , .B2( u1_u8_u0_n158 ) , .A( u1_u8_u0_n172 ) , .ZN( u1_u8_u0_n89 ) );
  AOI21_X1 u1_u8_u0_U70 (.A( u1_u8_u0_n138 ) , .B2( u1_u8_u0_n139 ) , .B1( u1_u8_u0_n140 ) , .ZN( u1_u8_u0_n157 ) );
  AOI211_X1 u1_u8_u0_U71 (.B( u1_u8_u0_n104 ) , .A( u1_u8_u0_n105 ) , .ZN( u1_u8_u0_n106 ) , .C2( u1_u8_u0_n113 ) , .C1( u1_u8_u0_n160 ) );
  INV_X1 u1_u8_u0_U72 (.ZN( u1_u8_u0_n174 ) , .A( u1_u8_u0_n89 ) );
  AOI21_X1 u1_u8_u0_U73 (.B2( u1_u8_u0_n141 ) , .B1( u1_u8_u0_n142 ) , .ZN( u1_u8_u0_n156 ) , .A( u1_u8_u0_n161 ) );
  AOI21_X1 u1_u8_u0_U74 (.ZN( u1_u8_u0_n116 ) , .B2( u1_u8_u0_n142 ) , .A( u1_u8_u0_n144 ) , .B1( u1_u8_u0_n166 ) );
  INV_X1 u1_u8_u0_U75 (.A( u1_u8_u0_n142 ) , .ZN( u1_u8_u0_n165 ) );
  NOR2_X1 u1_u8_u0_U76 (.A2( u1_u8_X_1 ) , .A1( u1_u8_X_2 ) , .ZN( u1_u8_u0_n92 ) );
  NOR2_X1 u1_u8_u0_U77 (.A2( u1_u8_X_2 ) , .ZN( u1_u8_u0_n103 ) , .A1( u1_u8_u0_n164 ) );
  INV_X1 u1_u8_u0_U78 (.A( u1_u8_X_2 ) , .ZN( u1_u8_u0_n163 ) );
  OAI221_X1 u1_u8_u0_U79 (.C1( u1_u8_u0_n121 ) , .ZN( u1_u8_u0_n122 ) , .B2( u1_u8_u0_n127 ) , .A( u1_u8_u0_n143 ) , .B1( u1_u8_u0_n144 ) , .C2( u1_u8_u0_n147 ) );
  AND2_X1 u1_u8_u0_U8 (.A1( u1_u8_u0_n114 ) , .A2( u1_u8_u0_n121 ) , .ZN( u1_u8_u0_n146 ) );
  AOI21_X1 u1_u8_u0_U80 (.B1( u1_u8_u0_n132 ) , .ZN( u1_u8_u0_n133 ) , .A( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n166 ) );
  OAI22_X1 u1_u8_u0_U81 (.ZN( u1_u8_u0_n105 ) , .A2( u1_u8_u0_n132 ) , .B1( u1_u8_u0_n146 ) , .A1( u1_u8_u0_n147 ) , .B2( u1_u8_u0_n161 ) );
  NAND2_X1 u1_u8_u0_U82 (.ZN( u1_u8_u0_n110 ) , .A2( u1_u8_u0_n132 ) , .A1( u1_u8_u0_n145 ) );
  INV_X1 u1_u8_u0_U83 (.A( u1_u8_u0_n119 ) , .ZN( u1_u8_u0_n167 ) );
  NAND2_X1 u1_u8_u0_U84 (.ZN( u1_u8_u0_n148 ) , .A1( u1_u8_u0_n93 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U85 (.A1( u1_u8_u0_n100 ) , .ZN( u1_u8_u0_n129 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U86 (.A1( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n128 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U87 (.ZN( u1_u8_u0_n142 ) , .A1( u1_u8_u0_n94 ) , .A2( u1_u8_u0_n95 ) );
  NAND3_X1 u1_u8_u0_U88 (.ZN( u1_out8_23 ) , .A3( u1_u8_u0_n137 ) , .A1( u1_u8_u0_n168 ) , .A2( u1_u8_u0_n171 ) );
  NAND3_X1 u1_u8_u0_U89 (.A3( u1_u8_u0_n127 ) , .A2( u1_u8_u0_n128 ) , .ZN( u1_u8_u0_n135 ) , .A1( u1_u8_u0_n150 ) );
  NAND2_X1 u1_u8_u0_U9 (.ZN( u1_u8_u0_n113 ) , .A1( u1_u8_u0_n139 ) , .A2( u1_u8_u0_n149 ) );
  NAND3_X1 u1_u8_u0_U90 (.ZN( u1_u8_u0_n117 ) , .A3( u1_u8_u0_n132 ) , .A2( u1_u8_u0_n139 ) , .A1( u1_u8_u0_n148 ) );
  NAND3_X1 u1_u8_u0_U91 (.ZN( u1_u8_u0_n109 ) , .A2( u1_u8_u0_n114 ) , .A3( u1_u8_u0_n140 ) , .A1( u1_u8_u0_n149 ) );
  NAND3_X1 u1_u8_u0_U92 (.ZN( u1_out8_9 ) , .A3( u1_u8_u0_n106 ) , .A2( u1_u8_u0_n171 ) , .A1( u1_u8_u0_n174 ) );
  NAND3_X1 u1_u8_u0_U93 (.A2( u1_u8_u0_n128 ) , .A1( u1_u8_u0_n132 ) , .A3( u1_u8_u0_n146 ) , .ZN( u1_u8_u0_n97 ) );
  OAI22_X1 u1_u8_u3_U10 (.B1( u1_u8_u3_n113 ) , .A2( u1_u8_u3_n135 ) , .A1( u1_u8_u3_n150 ) , .B2( u1_u8_u3_n164 ) , .ZN( u1_u8_u3_n98 ) );
  OAI211_X1 u1_u8_u3_U11 (.B( u1_u8_u3_n106 ) , .ZN( u1_u8_u3_n119 ) , .C2( u1_u8_u3_n128 ) , .C1( u1_u8_u3_n167 ) , .A( u1_u8_u3_n181 ) );
  AOI221_X1 u1_u8_u3_U12 (.C1( u1_u8_u3_n105 ) , .ZN( u1_u8_u3_n106 ) , .A( u1_u8_u3_n131 ) , .B2( u1_u8_u3_n132 ) , .C2( u1_u8_u3_n133 ) , .B1( u1_u8_u3_n169 ) );
  INV_X1 u1_u8_u3_U13 (.ZN( u1_u8_u3_n181 ) , .A( u1_u8_u3_n98 ) );
  NAND2_X1 u1_u8_u3_U14 (.ZN( u1_u8_u3_n105 ) , .A2( u1_u8_u3_n130 ) , .A1( u1_u8_u3_n155 ) );
  AOI22_X1 u1_u8_u3_U15 (.B1( u1_u8_u3_n115 ) , .A2( u1_u8_u3_n116 ) , .ZN( u1_u8_u3_n123 ) , .B2( u1_u8_u3_n133 ) , .A1( u1_u8_u3_n169 ) );
  NAND2_X1 u1_u8_u3_U16 (.ZN( u1_u8_u3_n116 ) , .A2( u1_u8_u3_n151 ) , .A1( u1_u8_u3_n182 ) );
  NOR2_X1 u1_u8_u3_U17 (.ZN( u1_u8_u3_n126 ) , .A2( u1_u8_u3_n150 ) , .A1( u1_u8_u3_n164 ) );
  AOI21_X1 u1_u8_u3_U18 (.ZN( u1_u8_u3_n112 ) , .B2( u1_u8_u3_n146 ) , .B1( u1_u8_u3_n155 ) , .A( u1_u8_u3_n167 ) );
  NAND2_X1 u1_u8_u3_U19 (.A1( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n142 ) , .A2( u1_u8_u3_n164 ) );
  NAND2_X1 u1_u8_u3_U20 (.ZN( u1_u8_u3_n132 ) , .A2( u1_u8_u3_n152 ) , .A1( u1_u8_u3_n156 ) );
  AND2_X1 u1_u8_u3_U21 (.A2( u1_u8_u3_n113 ) , .A1( u1_u8_u3_n114 ) , .ZN( u1_u8_u3_n151 ) );
  INV_X1 u1_u8_u3_U22 (.A( u1_u8_u3_n133 ) , .ZN( u1_u8_u3_n165 ) );
  INV_X1 u1_u8_u3_U23 (.A( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n170 ) );
  NAND2_X1 u1_u8_u3_U24 (.A1( u1_u8_u3_n107 ) , .A2( u1_u8_u3_n108 ) , .ZN( u1_u8_u3_n140 ) );
  NAND2_X1 u1_u8_u3_U25 (.ZN( u1_u8_u3_n117 ) , .A1( u1_u8_u3_n124 ) , .A2( u1_u8_u3_n148 ) );
  NAND2_X1 u1_u8_u3_U26 (.ZN( u1_u8_u3_n143 ) , .A1( u1_u8_u3_n165 ) , .A2( u1_u8_u3_n167 ) );
  INV_X1 u1_u8_u3_U27 (.A( u1_u8_u3_n130 ) , .ZN( u1_u8_u3_n177 ) );
  INV_X1 u1_u8_u3_U28 (.A( u1_u8_u3_n128 ) , .ZN( u1_u8_u3_n176 ) );
  INV_X1 u1_u8_u3_U29 (.A( u1_u8_u3_n155 ) , .ZN( u1_u8_u3_n174 ) );
  INV_X1 u1_u8_u3_U3 (.A( u1_u8_u3_n129 ) , .ZN( u1_u8_u3_n183 ) );
  INV_X1 u1_u8_u3_U30 (.A( u1_u8_u3_n139 ) , .ZN( u1_u8_u3_n185 ) );
  NOR2_X1 u1_u8_u3_U31 (.ZN( u1_u8_u3_n135 ) , .A2( u1_u8_u3_n141 ) , .A1( u1_u8_u3_n169 ) );
  OAI222_X1 u1_u8_u3_U32 (.C2( u1_u8_u3_n107 ) , .A2( u1_u8_u3_n108 ) , .B1( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n138 ) , .B2( u1_u8_u3_n146 ) , .C1( u1_u8_u3_n154 ) , .A1( u1_u8_u3_n164 ) );
  NOR4_X1 u1_u8_u3_U33 (.A4( u1_u8_u3_n157 ) , .A3( u1_u8_u3_n158 ) , .A2( u1_u8_u3_n159 ) , .A1( u1_u8_u3_n160 ) , .ZN( u1_u8_u3_n161 ) );
  AOI21_X1 u1_u8_u3_U34 (.B2( u1_u8_u3_n152 ) , .B1( u1_u8_u3_n153 ) , .ZN( u1_u8_u3_n158 ) , .A( u1_u8_u3_n164 ) );
  AOI21_X1 u1_u8_u3_U35 (.A( u1_u8_u3_n149 ) , .B2( u1_u8_u3_n150 ) , .B1( u1_u8_u3_n151 ) , .ZN( u1_u8_u3_n159 ) );
  AOI21_X1 u1_u8_u3_U36 (.A( u1_u8_u3_n154 ) , .B2( u1_u8_u3_n155 ) , .B1( u1_u8_u3_n156 ) , .ZN( u1_u8_u3_n157 ) );
  AOI211_X1 u1_u8_u3_U37 (.ZN( u1_u8_u3_n109 ) , .A( u1_u8_u3_n119 ) , .C2( u1_u8_u3_n129 ) , .B( u1_u8_u3_n138 ) , .C1( u1_u8_u3_n141 ) );
  AOI211_X1 u1_u8_u3_U38 (.B( u1_u8_u3_n119 ) , .A( u1_u8_u3_n120 ) , .C2( u1_u8_u3_n121 ) , .ZN( u1_u8_u3_n122 ) , .C1( u1_u8_u3_n179 ) );
  INV_X1 u1_u8_u3_U39 (.A( u1_u8_u3_n156 ) , .ZN( u1_u8_u3_n179 ) );
  INV_X1 u1_u8_u3_U4 (.A( u1_u8_u3_n140 ) , .ZN( u1_u8_u3_n182 ) );
  OAI22_X1 u1_u8_u3_U40 (.B1( u1_u8_u3_n118 ) , .ZN( u1_u8_u3_n120 ) , .A1( u1_u8_u3_n135 ) , .B2( u1_u8_u3_n154 ) , .A2( u1_u8_u3_n178 ) );
  AND3_X1 u1_u8_u3_U41 (.ZN( u1_u8_u3_n118 ) , .A2( u1_u8_u3_n124 ) , .A1( u1_u8_u3_n144 ) , .A3( u1_u8_u3_n152 ) );
  INV_X1 u1_u8_u3_U42 (.A( u1_u8_u3_n121 ) , .ZN( u1_u8_u3_n164 ) );
  NAND2_X1 u1_u8_u3_U43 (.ZN( u1_u8_u3_n133 ) , .A1( u1_u8_u3_n154 ) , .A2( u1_u8_u3_n164 ) );
  OAI211_X1 u1_u8_u3_U44 (.B( u1_u8_u3_n127 ) , .ZN( u1_u8_u3_n139 ) , .C1( u1_u8_u3_n150 ) , .C2( u1_u8_u3_n154 ) , .A( u1_u8_u3_n184 ) );
  INV_X1 u1_u8_u3_U45 (.A( u1_u8_u3_n125 ) , .ZN( u1_u8_u3_n184 ) );
  AOI221_X1 u1_u8_u3_U46 (.A( u1_u8_u3_n126 ) , .ZN( u1_u8_u3_n127 ) , .C2( u1_u8_u3_n132 ) , .C1( u1_u8_u3_n169 ) , .B2( u1_u8_u3_n170 ) , .B1( u1_u8_u3_n174 ) );
  OAI22_X1 u1_u8_u3_U47 (.A1( u1_u8_u3_n124 ) , .ZN( u1_u8_u3_n125 ) , .B2( u1_u8_u3_n145 ) , .A2( u1_u8_u3_n165 ) , .B1( u1_u8_u3_n167 ) );
  NOR2_X1 u1_u8_u3_U48 (.A1( u1_u8_u3_n113 ) , .ZN( u1_u8_u3_n131 ) , .A2( u1_u8_u3_n154 ) );
  NAND2_X1 u1_u8_u3_U49 (.A1( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n150 ) , .A2( u1_u8_u3_n99 ) );
  INV_X1 u1_u8_u3_U5 (.A( u1_u8_u3_n117 ) , .ZN( u1_u8_u3_n178 ) );
  NAND2_X1 u1_u8_u3_U50 (.A2( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n155 ) , .A1( u1_u8_u3_n97 ) );
  INV_X1 u1_u8_u3_U51 (.A( u1_u8_u3_n141 ) , .ZN( u1_u8_u3_n167 ) );
  AOI21_X1 u1_u8_u3_U52 (.B2( u1_u8_u3_n114 ) , .B1( u1_u8_u3_n146 ) , .A( u1_u8_u3_n154 ) , .ZN( u1_u8_u3_n94 ) );
  AOI21_X1 u1_u8_u3_U53 (.ZN( u1_u8_u3_n110 ) , .B2( u1_u8_u3_n142 ) , .B1( u1_u8_u3_n186 ) , .A( u1_u8_u3_n95 ) );
  INV_X1 u1_u8_u3_U54 (.A( u1_u8_u3_n145 ) , .ZN( u1_u8_u3_n186 ) );
  AOI21_X1 u1_u8_u3_U55 (.B1( u1_u8_u3_n124 ) , .A( u1_u8_u3_n149 ) , .B2( u1_u8_u3_n155 ) , .ZN( u1_u8_u3_n95 ) );
  INV_X1 u1_u8_u3_U56 (.A( u1_u8_u3_n149 ) , .ZN( u1_u8_u3_n169 ) );
  NAND2_X1 u1_u8_u3_U57 (.ZN( u1_u8_u3_n124 ) , .A1( u1_u8_u3_n96 ) , .A2( u1_u8_u3_n97 ) );
  NAND2_X1 u1_u8_u3_U58 (.A2( u1_u8_u3_n100 ) , .ZN( u1_u8_u3_n146 ) , .A1( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U59 (.A1( u1_u8_u3_n101 ) , .ZN( u1_u8_u3_n145 ) , .A2( u1_u8_u3_n99 ) );
  AOI221_X1 u1_u8_u3_U6 (.A( u1_u8_u3_n131 ) , .C2( u1_u8_u3_n132 ) , .C1( u1_u8_u3_n133 ) , .ZN( u1_u8_u3_n134 ) , .B1( u1_u8_u3_n143 ) , .B2( u1_u8_u3_n177 ) );
  NAND2_X1 u1_u8_u3_U60 (.A1( u1_u8_u3_n100 ) , .ZN( u1_u8_u3_n156 ) , .A2( u1_u8_u3_n99 ) );
  NAND2_X1 u1_u8_u3_U61 (.A2( u1_u8_u3_n101 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n148 ) );
  NAND2_X1 u1_u8_u3_U62 (.A1( u1_u8_u3_n100 ) , .A2( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n128 ) );
  NAND2_X1 u1_u8_u3_U63 (.A2( u1_u8_u3_n101 ) , .A1( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n152 ) );
  NAND2_X1 u1_u8_u3_U64 (.A2( u1_u8_u3_n101 ) , .ZN( u1_u8_u3_n114 ) , .A1( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U65 (.ZN( u1_u8_u3_n107 ) , .A1( u1_u8_u3_n97 ) , .A2( u1_u8_u3_n99 ) );
  NAND2_X1 u1_u8_u3_U66 (.A2( u1_u8_u3_n100 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n113 ) );
  NAND2_X1 u1_u8_u3_U67 (.A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n153 ) , .A2( u1_u8_u3_n97 ) );
  NAND2_X1 u1_u8_u3_U68 (.A2( u1_u8_u3_n103 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n130 ) );
  NAND2_X1 u1_u8_u3_U69 (.A2( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n144 ) , .A1( u1_u8_u3_n96 ) );
  OAI22_X1 u1_u8_u3_U7 (.B2( u1_u8_u3_n147 ) , .A2( u1_u8_u3_n148 ) , .ZN( u1_u8_u3_n160 ) , .B1( u1_u8_u3_n165 ) , .A1( u1_u8_u3_n168 ) );
  NAND2_X1 u1_u8_u3_U70 (.A1( u1_u8_u3_n102 ) , .A2( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n108 ) );
  NOR2_X1 u1_u8_u3_U71 (.A2( u1_u8_X_19 ) , .A1( u1_u8_X_20 ) , .ZN( u1_u8_u3_n99 ) );
  NOR2_X1 u1_u8_u3_U72 (.A2( u1_u8_X_21 ) , .A1( u1_u8_X_24 ) , .ZN( u1_u8_u3_n103 ) );
  NOR2_X1 u1_u8_u3_U73 (.A2( u1_u8_X_24 ) , .A1( u1_u8_u3_n171 ) , .ZN( u1_u8_u3_n97 ) );
  NOR2_X1 u1_u8_u3_U74 (.A2( u1_u8_X_23 ) , .ZN( u1_u8_u3_n141 ) , .A1( u1_u8_u3_n166 ) );
  NOR2_X1 u1_u8_u3_U75 (.A2( u1_u8_X_19 ) , .A1( u1_u8_u3_n172 ) , .ZN( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U76 (.A1( u1_u8_X_22 ) , .A2( u1_u8_X_23 ) , .ZN( u1_u8_u3_n154 ) );
  NAND2_X1 u1_u8_u3_U77 (.A1( u1_u8_X_23 ) , .ZN( u1_u8_u3_n149 ) , .A2( u1_u8_u3_n166 ) );
  NOR2_X1 u1_u8_u3_U78 (.A2( u1_u8_X_22 ) , .A1( u1_u8_X_23 ) , .ZN( u1_u8_u3_n121 ) );
  AND2_X1 u1_u8_u3_U79 (.A1( u1_u8_X_24 ) , .ZN( u1_u8_u3_n101 ) , .A2( u1_u8_u3_n171 ) );
  AND3_X1 u1_u8_u3_U8 (.A3( u1_u8_u3_n144 ) , .A2( u1_u8_u3_n145 ) , .A1( u1_u8_u3_n146 ) , .ZN( u1_u8_u3_n147 ) );
  AND2_X1 u1_u8_u3_U80 (.A1( u1_u8_X_19 ) , .ZN( u1_u8_u3_n102 ) , .A2( u1_u8_u3_n172 ) );
  AND2_X1 u1_u8_u3_U81 (.A1( u1_u8_X_21 ) , .A2( u1_u8_X_24 ) , .ZN( u1_u8_u3_n100 ) );
  AND2_X1 u1_u8_u3_U82 (.A2( u1_u8_X_19 ) , .A1( u1_u8_X_20 ) , .ZN( u1_u8_u3_n104 ) );
  INV_X1 u1_u8_u3_U83 (.A( u1_u8_X_22 ) , .ZN( u1_u8_u3_n166 ) );
  INV_X1 u1_u8_u3_U84 (.A( u1_u8_X_21 ) , .ZN( u1_u8_u3_n171 ) );
  INV_X1 u1_u8_u3_U85 (.A( u1_u8_X_20 ) , .ZN( u1_u8_u3_n172 ) );
  OR4_X1 u1_u8_u3_U86 (.ZN( u1_out8_10 ) , .A4( u1_u8_u3_n136 ) , .A3( u1_u8_u3_n137 ) , .A1( u1_u8_u3_n138 ) , .A2( u1_u8_u3_n139 ) );
  OAI222_X1 u1_u8_u3_U87 (.C1( u1_u8_u3_n128 ) , .ZN( u1_u8_u3_n137 ) , .B1( u1_u8_u3_n148 ) , .A2( u1_u8_u3_n150 ) , .B2( u1_u8_u3_n154 ) , .C2( u1_u8_u3_n164 ) , .A1( u1_u8_u3_n167 ) );
  OAI221_X1 u1_u8_u3_U88 (.A( u1_u8_u3_n134 ) , .B2( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n136 ) , .C1( u1_u8_u3_n149 ) , .B1( u1_u8_u3_n151 ) , .C2( u1_u8_u3_n183 ) );
  NAND4_X1 u1_u8_u3_U89 (.ZN( u1_out8_26 ) , .A4( u1_u8_u3_n109 ) , .A3( u1_u8_u3_n110 ) , .A2( u1_u8_u3_n111 ) , .A1( u1_u8_u3_n173 ) );
  INV_X1 u1_u8_u3_U9 (.A( u1_u8_u3_n143 ) , .ZN( u1_u8_u3_n168 ) );
  INV_X1 u1_u8_u3_U90 (.ZN( u1_u8_u3_n173 ) , .A( u1_u8_u3_n94 ) );
  OAI21_X1 u1_u8_u3_U91 (.ZN( u1_u8_u3_n111 ) , .B2( u1_u8_u3_n117 ) , .A( u1_u8_u3_n133 ) , .B1( u1_u8_u3_n176 ) );
  NAND4_X1 u1_u8_u3_U92 (.ZN( u1_out8_20 ) , .A4( u1_u8_u3_n122 ) , .A3( u1_u8_u3_n123 ) , .A1( u1_u8_u3_n175 ) , .A2( u1_u8_u3_n180 ) );
  INV_X1 u1_u8_u3_U93 (.A( u1_u8_u3_n126 ) , .ZN( u1_u8_u3_n180 ) );
  INV_X1 u1_u8_u3_U94 (.A( u1_u8_u3_n112 ) , .ZN( u1_u8_u3_n175 ) );
  NAND4_X1 u1_u8_u3_U95 (.ZN( u1_out8_1 ) , .A4( u1_u8_u3_n161 ) , .A3( u1_u8_u3_n162 ) , .A2( u1_u8_u3_n163 ) , .A1( u1_u8_u3_n185 ) );
  NAND2_X1 u1_u8_u3_U96 (.ZN( u1_u8_u3_n163 ) , .A2( u1_u8_u3_n170 ) , .A1( u1_u8_u3_n176 ) );
  AOI22_X1 u1_u8_u3_U97 (.B2( u1_u8_u3_n140 ) , .B1( u1_u8_u3_n141 ) , .A2( u1_u8_u3_n142 ) , .ZN( u1_u8_u3_n162 ) , .A1( u1_u8_u3_n177 ) );
  NAND3_X1 u1_u8_u3_U98 (.A1( u1_u8_u3_n114 ) , .ZN( u1_u8_u3_n115 ) , .A2( u1_u8_u3_n145 ) , .A3( u1_u8_u3_n153 ) );
  NAND3_X1 u1_u8_u3_U99 (.ZN( u1_u8_u3_n129 ) , .A2( u1_u8_u3_n144 ) , .A1( u1_u8_u3_n153 ) , .A3( u1_u8_u3_n182 ) );
  OAI22_X1 u1_u8_u4_U10 (.B2( u1_u8_u4_n135 ) , .ZN( u1_u8_u4_n137 ) , .B1( u1_u8_u4_n153 ) , .A1( u1_u8_u4_n155 ) , .A2( u1_u8_u4_n171 ) );
  AND3_X1 u1_u8_u4_U11 (.A2( u1_u8_u4_n134 ) , .ZN( u1_u8_u4_n135 ) , .A3( u1_u8_u4_n145 ) , .A1( u1_u8_u4_n157 ) );
  NAND2_X1 u1_u8_u4_U12 (.ZN( u1_u8_u4_n132 ) , .A2( u1_u8_u4_n170 ) , .A1( u1_u8_u4_n173 ) );
  AOI21_X1 u1_u8_u4_U13 (.B2( u1_u8_u4_n160 ) , .B1( u1_u8_u4_n161 ) , .ZN( u1_u8_u4_n162 ) , .A( u1_u8_u4_n170 ) );
  AOI21_X1 u1_u8_u4_U14 (.ZN( u1_u8_u4_n107 ) , .B2( u1_u8_u4_n143 ) , .A( u1_u8_u4_n174 ) , .B1( u1_u8_u4_n184 ) );
  AOI21_X1 u1_u8_u4_U15 (.B2( u1_u8_u4_n158 ) , .B1( u1_u8_u4_n159 ) , .ZN( u1_u8_u4_n163 ) , .A( u1_u8_u4_n174 ) );
  AOI21_X1 u1_u8_u4_U16 (.A( u1_u8_u4_n153 ) , .B2( u1_u8_u4_n154 ) , .B1( u1_u8_u4_n155 ) , .ZN( u1_u8_u4_n165 ) );
  AOI21_X1 u1_u8_u4_U17 (.A( u1_u8_u4_n156 ) , .B2( u1_u8_u4_n157 ) , .ZN( u1_u8_u4_n164 ) , .B1( u1_u8_u4_n184 ) );
  INV_X1 u1_u8_u4_U18 (.A( u1_u8_u4_n138 ) , .ZN( u1_u8_u4_n170 ) );
  AND2_X1 u1_u8_u4_U19 (.A2( u1_u8_u4_n120 ) , .ZN( u1_u8_u4_n155 ) , .A1( u1_u8_u4_n160 ) );
  INV_X1 u1_u8_u4_U20 (.A( u1_u8_u4_n156 ) , .ZN( u1_u8_u4_n175 ) );
  NAND2_X1 u1_u8_u4_U21 (.A2( u1_u8_u4_n118 ) , .ZN( u1_u8_u4_n131 ) , .A1( u1_u8_u4_n147 ) );
  NAND2_X1 u1_u8_u4_U22 (.A1( u1_u8_u4_n119 ) , .A2( u1_u8_u4_n120 ) , .ZN( u1_u8_u4_n130 ) );
  NAND2_X1 u1_u8_u4_U23 (.ZN( u1_u8_u4_n117 ) , .A2( u1_u8_u4_n118 ) , .A1( u1_u8_u4_n148 ) );
  NAND2_X1 u1_u8_u4_U24 (.ZN( u1_u8_u4_n129 ) , .A1( u1_u8_u4_n134 ) , .A2( u1_u8_u4_n148 ) );
  AND3_X1 u1_u8_u4_U25 (.A1( u1_u8_u4_n119 ) , .A2( u1_u8_u4_n143 ) , .A3( u1_u8_u4_n154 ) , .ZN( u1_u8_u4_n161 ) );
  AND2_X1 u1_u8_u4_U26 (.A1( u1_u8_u4_n145 ) , .A2( u1_u8_u4_n147 ) , .ZN( u1_u8_u4_n159 ) );
  OR3_X1 u1_u8_u4_U27 (.A3( u1_u8_u4_n114 ) , .A2( u1_u8_u4_n115 ) , .A1( u1_u8_u4_n116 ) , .ZN( u1_u8_u4_n136 ) );
  AOI21_X1 u1_u8_u4_U28 (.A( u1_u8_u4_n113 ) , .ZN( u1_u8_u4_n116 ) , .B2( u1_u8_u4_n173 ) , .B1( u1_u8_u4_n174 ) );
  AOI21_X1 u1_u8_u4_U29 (.ZN( u1_u8_u4_n115 ) , .B2( u1_u8_u4_n145 ) , .B1( u1_u8_u4_n146 ) , .A( u1_u8_u4_n156 ) );
  NOR2_X1 u1_u8_u4_U3 (.ZN( u1_u8_u4_n121 ) , .A1( u1_u8_u4_n181 ) , .A2( u1_u8_u4_n182 ) );
  OAI22_X1 u1_u8_u4_U30 (.ZN( u1_u8_u4_n114 ) , .A2( u1_u8_u4_n121 ) , .B1( u1_u8_u4_n160 ) , .B2( u1_u8_u4_n170 ) , .A1( u1_u8_u4_n171 ) );
  INV_X1 u1_u8_u4_U31 (.A( u1_u8_u4_n158 ) , .ZN( u1_u8_u4_n182 ) );
  INV_X1 u1_u8_u4_U32 (.ZN( u1_u8_u4_n181 ) , .A( u1_u8_u4_n96 ) );
  INV_X1 u1_u8_u4_U33 (.A( u1_u8_u4_n144 ) , .ZN( u1_u8_u4_n179 ) );
  INV_X1 u1_u8_u4_U34 (.A( u1_u8_u4_n157 ) , .ZN( u1_u8_u4_n178 ) );
  NAND2_X1 u1_u8_u4_U35 (.A2( u1_u8_u4_n154 ) , .A1( u1_u8_u4_n96 ) , .ZN( u1_u8_u4_n97 ) );
  INV_X1 u1_u8_u4_U36 (.ZN( u1_u8_u4_n186 ) , .A( u1_u8_u4_n95 ) );
  OAI221_X1 u1_u8_u4_U37 (.C1( u1_u8_u4_n134 ) , .B1( u1_u8_u4_n158 ) , .B2( u1_u8_u4_n171 ) , .C2( u1_u8_u4_n173 ) , .A( u1_u8_u4_n94 ) , .ZN( u1_u8_u4_n95 ) );
  AOI222_X1 u1_u8_u4_U38 (.B2( u1_u8_u4_n132 ) , .A1( u1_u8_u4_n138 ) , .C2( u1_u8_u4_n175 ) , .A2( u1_u8_u4_n179 ) , .C1( u1_u8_u4_n181 ) , .B1( u1_u8_u4_n185 ) , .ZN( u1_u8_u4_n94 ) );
  INV_X1 u1_u8_u4_U39 (.A( u1_u8_u4_n113 ) , .ZN( u1_u8_u4_n185 ) );
  INV_X1 u1_u8_u4_U4 (.A( u1_u8_u4_n117 ) , .ZN( u1_u8_u4_n184 ) );
  INV_X1 u1_u8_u4_U40 (.A( u1_u8_u4_n143 ) , .ZN( u1_u8_u4_n183 ) );
  NOR2_X1 u1_u8_u4_U41 (.ZN( u1_u8_u4_n138 ) , .A1( u1_u8_u4_n168 ) , .A2( u1_u8_u4_n169 ) );
  NOR2_X1 u1_u8_u4_U42 (.A1( u1_u8_u4_n150 ) , .A2( u1_u8_u4_n152 ) , .ZN( u1_u8_u4_n153 ) );
  NOR2_X1 u1_u8_u4_U43 (.A2( u1_u8_u4_n128 ) , .A1( u1_u8_u4_n138 ) , .ZN( u1_u8_u4_n156 ) );
  AOI22_X1 u1_u8_u4_U44 (.B2( u1_u8_u4_n122 ) , .A1( u1_u8_u4_n123 ) , .ZN( u1_u8_u4_n124 ) , .B1( u1_u8_u4_n128 ) , .A2( u1_u8_u4_n172 ) );
  INV_X1 u1_u8_u4_U45 (.A( u1_u8_u4_n153 ) , .ZN( u1_u8_u4_n172 ) );
  NAND2_X1 u1_u8_u4_U46 (.A2( u1_u8_u4_n120 ) , .ZN( u1_u8_u4_n123 ) , .A1( u1_u8_u4_n161 ) );
  AOI22_X1 u1_u8_u4_U47 (.B2( u1_u8_u4_n132 ) , .A2( u1_u8_u4_n133 ) , .ZN( u1_u8_u4_n140 ) , .A1( u1_u8_u4_n150 ) , .B1( u1_u8_u4_n179 ) );
  NAND2_X1 u1_u8_u4_U48 (.ZN( u1_u8_u4_n133 ) , .A2( u1_u8_u4_n146 ) , .A1( u1_u8_u4_n154 ) );
  NAND2_X1 u1_u8_u4_U49 (.A1( u1_u8_u4_n103 ) , .ZN( u1_u8_u4_n154 ) , .A2( u1_u8_u4_n98 ) );
  NOR4_X1 u1_u8_u4_U5 (.A4( u1_u8_u4_n106 ) , .A3( u1_u8_u4_n107 ) , .A2( u1_u8_u4_n108 ) , .A1( u1_u8_u4_n109 ) , .ZN( u1_u8_u4_n110 ) );
  NAND2_X1 u1_u8_u4_U50 (.A1( u1_u8_u4_n101 ) , .ZN( u1_u8_u4_n158 ) , .A2( u1_u8_u4_n99 ) );
  AOI21_X1 u1_u8_u4_U51 (.ZN( u1_u8_u4_n127 ) , .A( u1_u8_u4_n136 ) , .B2( u1_u8_u4_n150 ) , .B1( u1_u8_u4_n180 ) );
  INV_X1 u1_u8_u4_U52 (.A( u1_u8_u4_n160 ) , .ZN( u1_u8_u4_n180 ) );
  NAND2_X1 u1_u8_u4_U53 (.A2( u1_u8_u4_n104 ) , .A1( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n146 ) );
  NAND2_X1 u1_u8_u4_U54 (.A2( u1_u8_u4_n101 ) , .A1( u1_u8_u4_n102 ) , .ZN( u1_u8_u4_n160 ) );
  NAND2_X1 u1_u8_u4_U55 (.ZN( u1_u8_u4_n134 ) , .A1( u1_u8_u4_n98 ) , .A2( u1_u8_u4_n99 ) );
  NAND2_X1 u1_u8_u4_U56 (.A1( u1_u8_u4_n103 ) , .A2( u1_u8_u4_n104 ) , .ZN( u1_u8_u4_n143 ) );
  NAND2_X1 u1_u8_u4_U57 (.A2( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n145 ) , .A1( u1_u8_u4_n98 ) );
  NAND2_X1 u1_u8_u4_U58 (.A1( u1_u8_u4_n100 ) , .A2( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n120 ) );
  NAND2_X1 u1_u8_u4_U59 (.A1( u1_u8_u4_n102 ) , .A2( u1_u8_u4_n104 ) , .ZN( u1_u8_u4_n148 ) );
  AOI21_X1 u1_u8_u4_U6 (.ZN( u1_u8_u4_n106 ) , .B2( u1_u8_u4_n146 ) , .B1( u1_u8_u4_n158 ) , .A( u1_u8_u4_n170 ) );
  NAND2_X1 u1_u8_u4_U60 (.A2( u1_u8_u4_n100 ) , .A1( u1_u8_u4_n103 ) , .ZN( u1_u8_u4_n157 ) );
  INV_X1 u1_u8_u4_U61 (.A( u1_u8_u4_n150 ) , .ZN( u1_u8_u4_n173 ) );
  INV_X1 u1_u8_u4_U62 (.A( u1_u8_u4_n152 ) , .ZN( u1_u8_u4_n171 ) );
  NAND2_X1 u1_u8_u4_U63 (.A1( u1_u8_u4_n100 ) , .ZN( u1_u8_u4_n118 ) , .A2( u1_u8_u4_n99 ) );
  NAND2_X1 u1_u8_u4_U64 (.A2( u1_u8_u4_n100 ) , .A1( u1_u8_u4_n102 ) , .ZN( u1_u8_u4_n144 ) );
  NAND2_X1 u1_u8_u4_U65 (.A2( u1_u8_u4_n101 ) , .A1( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n96 ) );
  INV_X1 u1_u8_u4_U66 (.A( u1_u8_u4_n128 ) , .ZN( u1_u8_u4_n174 ) );
  NAND2_X1 u1_u8_u4_U67 (.A2( u1_u8_u4_n102 ) , .ZN( u1_u8_u4_n119 ) , .A1( u1_u8_u4_n98 ) );
  NAND2_X1 u1_u8_u4_U68 (.A2( u1_u8_u4_n101 ) , .A1( u1_u8_u4_n103 ) , .ZN( u1_u8_u4_n147 ) );
  NAND2_X1 u1_u8_u4_U69 (.A2( u1_u8_u4_n104 ) , .ZN( u1_u8_u4_n113 ) , .A1( u1_u8_u4_n99 ) );
  AOI21_X1 u1_u8_u4_U7 (.ZN( u1_u8_u4_n108 ) , .B2( u1_u8_u4_n134 ) , .B1( u1_u8_u4_n155 ) , .A( u1_u8_u4_n156 ) );
  NOR2_X1 u1_u8_u4_U70 (.A2( u1_u8_X_28 ) , .ZN( u1_u8_u4_n150 ) , .A1( u1_u8_u4_n168 ) );
  NOR2_X1 u1_u8_u4_U71 (.A2( u1_u8_X_29 ) , .ZN( u1_u8_u4_n152 ) , .A1( u1_u8_u4_n169 ) );
  NOR2_X1 u1_u8_u4_U72 (.A2( u1_u8_X_30 ) , .ZN( u1_u8_u4_n105 ) , .A1( u1_u8_u4_n176 ) );
  NOR2_X1 u1_u8_u4_U73 (.A2( u1_u8_X_26 ) , .ZN( u1_u8_u4_n100 ) , .A1( u1_u8_u4_n177 ) );
  NOR2_X1 u1_u8_u4_U74 (.A2( u1_u8_X_28 ) , .A1( u1_u8_X_29 ) , .ZN( u1_u8_u4_n128 ) );
  NOR2_X1 u1_u8_u4_U75 (.A2( u1_u8_X_27 ) , .A1( u1_u8_X_30 ) , .ZN( u1_u8_u4_n102 ) );
  NOR2_X1 u1_u8_u4_U76 (.A2( u1_u8_X_25 ) , .A1( u1_u8_X_26 ) , .ZN( u1_u8_u4_n98 ) );
  AND2_X1 u1_u8_u4_U77 (.A2( u1_u8_X_25 ) , .A1( u1_u8_X_26 ) , .ZN( u1_u8_u4_n104 ) );
  AND2_X1 u1_u8_u4_U78 (.A1( u1_u8_X_30 ) , .A2( u1_u8_u4_n176 ) , .ZN( u1_u8_u4_n99 ) );
  AND2_X1 u1_u8_u4_U79 (.A1( u1_u8_X_26 ) , .ZN( u1_u8_u4_n101 ) , .A2( u1_u8_u4_n177 ) );
  AOI21_X1 u1_u8_u4_U8 (.ZN( u1_u8_u4_n109 ) , .A( u1_u8_u4_n153 ) , .B1( u1_u8_u4_n159 ) , .B2( u1_u8_u4_n184 ) );
  AND2_X1 u1_u8_u4_U80 (.A1( u1_u8_X_27 ) , .A2( u1_u8_X_30 ) , .ZN( u1_u8_u4_n103 ) );
  INV_X1 u1_u8_u4_U81 (.A( u1_u8_X_28 ) , .ZN( u1_u8_u4_n169 ) );
  INV_X1 u1_u8_u4_U82 (.A( u1_u8_X_29 ) , .ZN( u1_u8_u4_n168 ) );
  INV_X1 u1_u8_u4_U83 (.A( u1_u8_X_25 ) , .ZN( u1_u8_u4_n177 ) );
  INV_X1 u1_u8_u4_U84 (.A( u1_u8_X_27 ) , .ZN( u1_u8_u4_n176 ) );
  NAND4_X1 u1_u8_u4_U85 (.ZN( u1_out8_25 ) , .A4( u1_u8_u4_n139 ) , .A3( u1_u8_u4_n140 ) , .A2( u1_u8_u4_n141 ) , .A1( u1_u8_u4_n142 ) );
  OAI21_X1 u1_u8_u4_U86 (.B2( u1_u8_u4_n131 ) , .ZN( u1_u8_u4_n141 ) , .A( u1_u8_u4_n175 ) , .B1( u1_u8_u4_n183 ) );
  OAI21_X1 u1_u8_u4_U87 (.A( u1_u8_u4_n128 ) , .B2( u1_u8_u4_n129 ) , .B1( u1_u8_u4_n130 ) , .ZN( u1_u8_u4_n142 ) );
  NAND4_X1 u1_u8_u4_U88 (.ZN( u1_out8_14 ) , .A4( u1_u8_u4_n124 ) , .A3( u1_u8_u4_n125 ) , .A2( u1_u8_u4_n126 ) , .A1( u1_u8_u4_n127 ) );
  AOI22_X1 u1_u8_u4_U89 (.B2( u1_u8_u4_n117 ) , .ZN( u1_u8_u4_n126 ) , .A1( u1_u8_u4_n129 ) , .B1( u1_u8_u4_n152 ) , .A2( u1_u8_u4_n175 ) );
  AOI211_X1 u1_u8_u4_U9 (.B( u1_u8_u4_n136 ) , .A( u1_u8_u4_n137 ) , .C2( u1_u8_u4_n138 ) , .ZN( u1_u8_u4_n139 ) , .C1( u1_u8_u4_n182 ) );
  AOI22_X1 u1_u8_u4_U90 (.ZN( u1_u8_u4_n125 ) , .B2( u1_u8_u4_n131 ) , .A2( u1_u8_u4_n132 ) , .B1( u1_u8_u4_n138 ) , .A1( u1_u8_u4_n178 ) );
  NAND4_X1 u1_u8_u4_U91 (.ZN( u1_out8_8 ) , .A4( u1_u8_u4_n110 ) , .A3( u1_u8_u4_n111 ) , .A2( u1_u8_u4_n112 ) , .A1( u1_u8_u4_n186 ) );
  NAND2_X1 u1_u8_u4_U92 (.ZN( u1_u8_u4_n112 ) , .A2( u1_u8_u4_n130 ) , .A1( u1_u8_u4_n150 ) );
  AOI22_X1 u1_u8_u4_U93 (.ZN( u1_u8_u4_n111 ) , .B2( u1_u8_u4_n132 ) , .A1( u1_u8_u4_n152 ) , .B1( u1_u8_u4_n178 ) , .A2( u1_u8_u4_n97 ) );
  AOI22_X1 u1_u8_u4_U94 (.B2( u1_u8_u4_n149 ) , .B1( u1_u8_u4_n150 ) , .A2( u1_u8_u4_n151 ) , .A1( u1_u8_u4_n152 ) , .ZN( u1_u8_u4_n167 ) );
  NOR4_X1 u1_u8_u4_U95 (.A4( u1_u8_u4_n162 ) , .A3( u1_u8_u4_n163 ) , .A2( u1_u8_u4_n164 ) , .A1( u1_u8_u4_n165 ) , .ZN( u1_u8_u4_n166 ) );
  NAND3_X1 u1_u8_u4_U96 (.ZN( u1_out8_3 ) , .A3( u1_u8_u4_n166 ) , .A1( u1_u8_u4_n167 ) , .A2( u1_u8_u4_n186 ) );
  NAND3_X1 u1_u8_u4_U97 (.A3( u1_u8_u4_n146 ) , .A2( u1_u8_u4_n147 ) , .A1( u1_u8_u4_n148 ) , .ZN( u1_u8_u4_n149 ) );
  NAND3_X1 u1_u8_u4_U98 (.A3( u1_u8_u4_n143 ) , .A2( u1_u8_u4_n144 ) , .A1( u1_u8_u4_n145 ) , .ZN( u1_u8_u4_n151 ) );
  NAND3_X1 u1_u8_u4_U99 (.A3( u1_u8_u4_n121 ) , .ZN( u1_u8_u4_n122 ) , .A2( u1_u8_u4_n144 ) , .A1( u1_u8_u4_n154 ) );
  NOR2_X1 u1_u8_u5_U10 (.ZN( u1_u8_u5_n135 ) , .A1( u1_u8_u5_n173 ) , .A2( u1_u8_u5_n176 ) );
  NOR3_X1 u1_u8_u5_U100 (.A3( u1_u8_u5_n141 ) , .A1( u1_u8_u5_n142 ) , .ZN( u1_u8_u5_n143 ) , .A2( u1_u8_u5_n191 ) );
  NAND4_X1 u1_u8_u5_U101 (.ZN( u1_out8_4 ) , .A4( u1_u8_u5_n112 ) , .A2( u1_u8_u5_n113 ) , .A1( u1_u8_u5_n114 ) , .A3( u1_u8_u5_n195 ) );
  AOI211_X1 u1_u8_u5_U102 (.A( u1_u8_u5_n110 ) , .C1( u1_u8_u5_n111 ) , .ZN( u1_u8_u5_n112 ) , .B( u1_u8_u5_n118 ) , .C2( u1_u8_u5_n177 ) );
  INV_X1 u1_u8_u5_U103 (.A( u1_u8_u5_n102 ) , .ZN( u1_u8_u5_n195 ) );
  NAND3_X1 u1_u8_u5_U104 (.A2( u1_u8_u5_n154 ) , .A3( u1_u8_u5_n158 ) , .A1( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n99 ) );
  INV_X1 u1_u8_u5_U11 (.A( u1_u8_u5_n121 ) , .ZN( u1_u8_u5_n177 ) );
  NOR2_X1 u1_u8_u5_U12 (.ZN( u1_u8_u5_n160 ) , .A2( u1_u8_u5_n173 ) , .A1( u1_u8_u5_n177 ) );
  INV_X1 u1_u8_u5_U13 (.A( u1_u8_u5_n150 ) , .ZN( u1_u8_u5_n174 ) );
  AOI21_X1 u1_u8_u5_U14 (.A( u1_u8_u5_n160 ) , .B2( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n162 ) , .B1( u1_u8_u5_n192 ) );
  INV_X1 u1_u8_u5_U15 (.A( u1_u8_u5_n159 ) , .ZN( u1_u8_u5_n192 ) );
  AOI21_X1 u1_u8_u5_U16 (.A( u1_u8_u5_n156 ) , .B2( u1_u8_u5_n157 ) , .B1( u1_u8_u5_n158 ) , .ZN( u1_u8_u5_n163 ) );
  AOI21_X1 u1_u8_u5_U17 (.B2( u1_u8_u5_n139 ) , .B1( u1_u8_u5_n140 ) , .ZN( u1_u8_u5_n141 ) , .A( u1_u8_u5_n150 ) );
  OAI21_X1 u1_u8_u5_U18 (.A( u1_u8_u5_n133 ) , .B2( u1_u8_u5_n134 ) , .B1( u1_u8_u5_n135 ) , .ZN( u1_u8_u5_n142 ) );
  OAI21_X1 u1_u8_u5_U19 (.ZN( u1_u8_u5_n133 ) , .B2( u1_u8_u5_n147 ) , .A( u1_u8_u5_n173 ) , .B1( u1_u8_u5_n188 ) );
  NAND2_X1 u1_u8_u5_U20 (.A2( u1_u8_u5_n119 ) , .A1( u1_u8_u5_n123 ) , .ZN( u1_u8_u5_n137 ) );
  INV_X1 u1_u8_u5_U21 (.A( u1_u8_u5_n155 ) , .ZN( u1_u8_u5_n194 ) );
  NAND2_X1 u1_u8_u5_U22 (.A1( u1_u8_u5_n121 ) , .ZN( u1_u8_u5_n132 ) , .A2( u1_u8_u5_n172 ) );
  NAND2_X1 u1_u8_u5_U23 (.A2( u1_u8_u5_n122 ) , .ZN( u1_u8_u5_n136 ) , .A1( u1_u8_u5_n154 ) );
  NAND2_X1 u1_u8_u5_U24 (.A2( u1_u8_u5_n119 ) , .A1( u1_u8_u5_n120 ) , .ZN( u1_u8_u5_n159 ) );
  INV_X1 u1_u8_u5_U25 (.A( u1_u8_u5_n156 ) , .ZN( u1_u8_u5_n175 ) );
  INV_X1 u1_u8_u5_U26 (.A( u1_u8_u5_n158 ) , .ZN( u1_u8_u5_n188 ) );
  INV_X1 u1_u8_u5_U27 (.A( u1_u8_u5_n152 ) , .ZN( u1_u8_u5_n179 ) );
  INV_X1 u1_u8_u5_U28 (.A( u1_u8_u5_n140 ) , .ZN( u1_u8_u5_n182 ) );
  INV_X1 u1_u8_u5_U29 (.A( u1_u8_u5_n151 ) , .ZN( u1_u8_u5_n183 ) );
  NOR2_X1 u1_u8_u5_U3 (.ZN( u1_u8_u5_n134 ) , .A1( u1_u8_u5_n183 ) , .A2( u1_u8_u5_n190 ) );
  INV_X1 u1_u8_u5_U30 (.A( u1_u8_u5_n123 ) , .ZN( u1_u8_u5_n185 ) );
  INV_X1 u1_u8_u5_U31 (.A( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n184 ) );
  INV_X1 u1_u8_u5_U32 (.A( u1_u8_u5_n139 ) , .ZN( u1_u8_u5_n189 ) );
  INV_X1 u1_u8_u5_U33 (.A( u1_u8_u5_n157 ) , .ZN( u1_u8_u5_n190 ) );
  INV_X1 u1_u8_u5_U34 (.A( u1_u8_u5_n120 ) , .ZN( u1_u8_u5_n193 ) );
  NAND2_X1 u1_u8_u5_U35 (.ZN( u1_u8_u5_n111 ) , .A1( u1_u8_u5_n140 ) , .A2( u1_u8_u5_n155 ) );
  INV_X1 u1_u8_u5_U36 (.A( u1_u8_u5_n117 ) , .ZN( u1_u8_u5_n196 ) );
  OAI221_X1 u1_u8_u5_U37 (.A( u1_u8_u5_n116 ) , .ZN( u1_u8_u5_n117 ) , .B2( u1_u8_u5_n119 ) , .C1( u1_u8_u5_n153 ) , .C2( u1_u8_u5_n158 ) , .B1( u1_u8_u5_n172 ) );
  AOI222_X1 u1_u8_u5_U38 (.ZN( u1_u8_u5_n116 ) , .B2( u1_u8_u5_n145 ) , .C1( u1_u8_u5_n148 ) , .A2( u1_u8_u5_n174 ) , .C2( u1_u8_u5_n177 ) , .B1( u1_u8_u5_n187 ) , .A1( u1_u8_u5_n193 ) );
  INV_X1 u1_u8_u5_U39 (.A( u1_u8_u5_n115 ) , .ZN( u1_u8_u5_n187 ) );
  INV_X1 u1_u8_u5_U4 (.A( u1_u8_u5_n138 ) , .ZN( u1_u8_u5_n191 ) );
  NOR2_X1 u1_u8_u5_U40 (.ZN( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n170 ) , .A2( u1_u8_u5_n180 ) );
  OAI221_X1 u1_u8_u5_U41 (.A( u1_u8_u5_n101 ) , .ZN( u1_u8_u5_n102 ) , .C2( u1_u8_u5_n115 ) , .C1( u1_u8_u5_n126 ) , .B1( u1_u8_u5_n134 ) , .B2( u1_u8_u5_n160 ) );
  OAI21_X1 u1_u8_u5_U42 (.ZN( u1_u8_u5_n101 ) , .B1( u1_u8_u5_n137 ) , .A( u1_u8_u5_n146 ) , .B2( u1_u8_u5_n147 ) );
  AOI22_X1 u1_u8_u5_U43 (.B2( u1_u8_u5_n131 ) , .A2( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n169 ) , .B1( u1_u8_u5_n174 ) , .A1( u1_u8_u5_n185 ) );
  NOR2_X1 u1_u8_u5_U44 (.A1( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n150 ) , .A2( u1_u8_u5_n173 ) );
  AOI21_X1 u1_u8_u5_U45 (.A( u1_u8_u5_n118 ) , .B2( u1_u8_u5_n145 ) , .ZN( u1_u8_u5_n168 ) , .B1( u1_u8_u5_n186 ) );
  INV_X1 u1_u8_u5_U46 (.A( u1_u8_u5_n122 ) , .ZN( u1_u8_u5_n186 ) );
  NOR2_X1 u1_u8_u5_U47 (.A1( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n152 ) , .A2( u1_u8_u5_n176 ) );
  NOR2_X1 u1_u8_u5_U48 (.A1( u1_u8_u5_n115 ) , .ZN( u1_u8_u5_n118 ) , .A2( u1_u8_u5_n153 ) );
  NOR2_X1 u1_u8_u5_U49 (.A2( u1_u8_u5_n145 ) , .ZN( u1_u8_u5_n156 ) , .A1( u1_u8_u5_n174 ) );
  OAI21_X1 u1_u8_u5_U5 (.B2( u1_u8_u5_n136 ) , .B1( u1_u8_u5_n137 ) , .ZN( u1_u8_u5_n138 ) , .A( u1_u8_u5_n177 ) );
  NOR2_X1 u1_u8_u5_U50 (.ZN( u1_u8_u5_n121 ) , .A2( u1_u8_u5_n145 ) , .A1( u1_u8_u5_n176 ) );
  AOI22_X1 u1_u8_u5_U51 (.ZN( u1_u8_u5_n114 ) , .A2( u1_u8_u5_n137 ) , .A1( u1_u8_u5_n145 ) , .B2( u1_u8_u5_n175 ) , .B1( u1_u8_u5_n193 ) );
  OAI211_X1 u1_u8_u5_U52 (.B( u1_u8_u5_n124 ) , .A( u1_u8_u5_n125 ) , .C2( u1_u8_u5_n126 ) , .C1( u1_u8_u5_n127 ) , .ZN( u1_u8_u5_n128 ) );
  NOR3_X1 u1_u8_u5_U53 (.ZN( u1_u8_u5_n127 ) , .A1( u1_u8_u5_n136 ) , .A3( u1_u8_u5_n148 ) , .A2( u1_u8_u5_n182 ) );
  OAI21_X1 u1_u8_u5_U54 (.ZN( u1_u8_u5_n124 ) , .A( u1_u8_u5_n177 ) , .B2( u1_u8_u5_n183 ) , .B1( u1_u8_u5_n189 ) );
  OAI21_X1 u1_u8_u5_U55 (.ZN( u1_u8_u5_n125 ) , .A( u1_u8_u5_n174 ) , .B2( u1_u8_u5_n185 ) , .B1( u1_u8_u5_n190 ) );
  AOI21_X1 u1_u8_u5_U56 (.A( u1_u8_u5_n153 ) , .B2( u1_u8_u5_n154 ) , .B1( u1_u8_u5_n155 ) , .ZN( u1_u8_u5_n164 ) );
  AOI21_X1 u1_u8_u5_U57 (.ZN( u1_u8_u5_n110 ) , .B1( u1_u8_u5_n122 ) , .B2( u1_u8_u5_n139 ) , .A( u1_u8_u5_n153 ) );
  INV_X1 u1_u8_u5_U58 (.A( u1_u8_u5_n153 ) , .ZN( u1_u8_u5_n176 ) );
  INV_X1 u1_u8_u5_U59 (.A( u1_u8_u5_n126 ) , .ZN( u1_u8_u5_n173 ) );
  AOI222_X1 u1_u8_u5_U6 (.ZN( u1_u8_u5_n113 ) , .A1( u1_u8_u5_n131 ) , .C1( u1_u8_u5_n148 ) , .B2( u1_u8_u5_n174 ) , .C2( u1_u8_u5_n178 ) , .A2( u1_u8_u5_n179 ) , .B1( u1_u8_u5_n99 ) );
  AND2_X1 u1_u8_u5_U60 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n147 ) );
  AND2_X1 u1_u8_u5_U61 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n148 ) );
  NAND2_X1 u1_u8_u5_U62 (.A1( u1_u8_u5_n105 ) , .A2( u1_u8_u5_n106 ) , .ZN( u1_u8_u5_n158 ) );
  NAND2_X1 u1_u8_u5_U63 (.A2( u1_u8_u5_n108 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n139 ) );
  NAND2_X1 u1_u8_u5_U64 (.A1( u1_u8_u5_n106 ) , .A2( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n119 ) );
  NAND2_X1 u1_u8_u5_U65 (.A2( u1_u8_u5_n103 ) , .A1( u1_u8_u5_n105 ) , .ZN( u1_u8_u5_n140 ) );
  NAND2_X1 u1_u8_u5_U66 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n105 ) , .ZN( u1_u8_u5_n155 ) );
  NAND2_X1 u1_u8_u5_U67 (.A2( u1_u8_u5_n106 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n122 ) );
  NAND2_X1 u1_u8_u5_U68 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n106 ) , .ZN( u1_u8_u5_n115 ) );
  NAND2_X1 u1_u8_u5_U69 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n103 ) , .ZN( u1_u8_u5_n161 ) );
  INV_X1 u1_u8_u5_U7 (.A( u1_u8_u5_n135 ) , .ZN( u1_u8_u5_n178 ) );
  NAND2_X1 u1_u8_u5_U70 (.A1( u1_u8_u5_n105 ) , .A2( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n154 ) );
  INV_X1 u1_u8_u5_U71 (.A( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n172 ) );
  NAND2_X1 u1_u8_u5_U72 (.A1( u1_u8_u5_n103 ) , .A2( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n123 ) );
  NAND2_X1 u1_u8_u5_U73 (.A2( u1_u8_u5_n103 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n151 ) );
  NAND2_X1 u1_u8_u5_U74 (.A2( u1_u8_u5_n107 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n120 ) );
  NAND2_X1 u1_u8_u5_U75 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n157 ) );
  AND2_X1 u1_u8_u5_U76 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n104 ) , .ZN( u1_u8_u5_n131 ) );
  NOR2_X1 u1_u8_u5_U77 (.A2( u1_u8_X_34 ) , .A1( u1_u8_X_35 ) , .ZN( u1_u8_u5_n145 ) );
  NOR2_X1 u1_u8_u5_U78 (.A2( u1_u8_X_34 ) , .ZN( u1_u8_u5_n146 ) , .A1( u1_u8_u5_n171 ) );
  NOR2_X1 u1_u8_u5_U79 (.A2( u1_u8_X_31 ) , .A1( u1_u8_X_32 ) , .ZN( u1_u8_u5_n103 ) );
  OAI22_X1 u1_u8_u5_U8 (.B2( u1_u8_u5_n149 ) , .B1( u1_u8_u5_n150 ) , .A2( u1_u8_u5_n151 ) , .A1( u1_u8_u5_n152 ) , .ZN( u1_u8_u5_n165 ) );
  NOR2_X1 u1_u8_u5_U80 (.A2( u1_u8_X_36 ) , .ZN( u1_u8_u5_n105 ) , .A1( u1_u8_u5_n180 ) );
  NOR2_X1 u1_u8_u5_U81 (.A2( u1_u8_X_33 ) , .ZN( u1_u8_u5_n108 ) , .A1( u1_u8_u5_n170 ) );
  NOR2_X1 u1_u8_u5_U82 (.A2( u1_u8_X_33 ) , .A1( u1_u8_X_36 ) , .ZN( u1_u8_u5_n107 ) );
  NOR2_X1 u1_u8_u5_U83 (.A2( u1_u8_X_31 ) , .ZN( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n181 ) );
  NAND2_X1 u1_u8_u5_U84 (.A2( u1_u8_X_34 ) , .A1( u1_u8_X_35 ) , .ZN( u1_u8_u5_n153 ) );
  NAND2_X1 u1_u8_u5_U85 (.A1( u1_u8_X_34 ) , .ZN( u1_u8_u5_n126 ) , .A2( u1_u8_u5_n171 ) );
  AND2_X1 u1_u8_u5_U86 (.A1( u1_u8_X_31 ) , .A2( u1_u8_X_32 ) , .ZN( u1_u8_u5_n106 ) );
  AND2_X1 u1_u8_u5_U87 (.A1( u1_u8_X_31 ) , .ZN( u1_u8_u5_n109 ) , .A2( u1_u8_u5_n181 ) );
  INV_X1 u1_u8_u5_U88 (.A( u1_u8_X_33 ) , .ZN( u1_u8_u5_n180 ) );
  INV_X1 u1_u8_u5_U89 (.A( u1_u8_X_35 ) , .ZN( u1_u8_u5_n171 ) );
  NOR3_X1 u1_u8_u5_U9 (.A2( u1_u8_u5_n147 ) , .A1( u1_u8_u5_n148 ) , .ZN( u1_u8_u5_n149 ) , .A3( u1_u8_u5_n194 ) );
  INV_X1 u1_u8_u5_U90 (.A( u1_u8_X_36 ) , .ZN( u1_u8_u5_n170 ) );
  INV_X1 u1_u8_u5_U91 (.A( u1_u8_X_32 ) , .ZN( u1_u8_u5_n181 ) );
  NAND4_X1 u1_u8_u5_U92 (.ZN( u1_out8_29 ) , .A4( u1_u8_u5_n129 ) , .A3( u1_u8_u5_n130 ) , .A2( u1_u8_u5_n168 ) , .A1( u1_u8_u5_n196 ) );
  AOI221_X1 u1_u8_u5_U93 (.A( u1_u8_u5_n128 ) , .ZN( u1_u8_u5_n129 ) , .C2( u1_u8_u5_n132 ) , .B2( u1_u8_u5_n159 ) , .B1( u1_u8_u5_n176 ) , .C1( u1_u8_u5_n184 ) );
  AOI222_X1 u1_u8_u5_U94 (.ZN( u1_u8_u5_n130 ) , .A2( u1_u8_u5_n146 ) , .B1( u1_u8_u5_n147 ) , .C2( u1_u8_u5_n175 ) , .B2( u1_u8_u5_n179 ) , .A1( u1_u8_u5_n188 ) , .C1( u1_u8_u5_n194 ) );
  NAND4_X1 u1_u8_u5_U95 (.ZN( u1_out8_19 ) , .A4( u1_u8_u5_n166 ) , .A3( u1_u8_u5_n167 ) , .A2( u1_u8_u5_n168 ) , .A1( u1_u8_u5_n169 ) );
  AOI22_X1 u1_u8_u5_U96 (.B2( u1_u8_u5_n145 ) , .A2( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n167 ) , .B1( u1_u8_u5_n182 ) , .A1( u1_u8_u5_n189 ) );
  NOR4_X1 u1_u8_u5_U97 (.A4( u1_u8_u5_n162 ) , .A3( u1_u8_u5_n163 ) , .A2( u1_u8_u5_n164 ) , .A1( u1_u8_u5_n165 ) , .ZN( u1_u8_u5_n166 ) );
  NAND4_X1 u1_u8_u5_U98 (.ZN( u1_out8_11 ) , .A4( u1_u8_u5_n143 ) , .A3( u1_u8_u5_n144 ) , .A2( u1_u8_u5_n169 ) , .A1( u1_u8_u5_n196 ) );
  AOI22_X1 u1_u8_u5_U99 (.A2( u1_u8_u5_n132 ) , .ZN( u1_u8_u5_n144 ) , .B2( u1_u8_u5_n145 ) , .B1( u1_u8_u5_n184 ) , .A1( u1_u8_u5_n194 ) );
  AOI22_X1 u1_u8_u6_U10 (.A2( u1_u8_u6_n151 ) , .B2( u1_u8_u6_n161 ) , .A1( u1_u8_u6_n167 ) , .B1( u1_u8_u6_n170 ) , .ZN( u1_u8_u6_n89 ) );
  AOI21_X1 u1_u8_u6_U11 (.B1( u1_u8_u6_n107 ) , .B2( u1_u8_u6_n132 ) , .A( u1_u8_u6_n158 ) , .ZN( u1_u8_u6_n88 ) );
  AOI21_X1 u1_u8_u6_U12 (.B2( u1_u8_u6_n147 ) , .B1( u1_u8_u6_n148 ) , .ZN( u1_u8_u6_n149 ) , .A( u1_u8_u6_n158 ) );
  AOI21_X1 u1_u8_u6_U13 (.ZN( u1_u8_u6_n106 ) , .A( u1_u8_u6_n142 ) , .B2( u1_u8_u6_n159 ) , .B1( u1_u8_u6_n164 ) );
  INV_X1 u1_u8_u6_U14 (.A( u1_u8_u6_n155 ) , .ZN( u1_u8_u6_n161 ) );
  INV_X1 u1_u8_u6_U15 (.A( u1_u8_u6_n128 ) , .ZN( u1_u8_u6_n164 ) );
  NAND2_X1 u1_u8_u6_U16 (.ZN( u1_u8_u6_n110 ) , .A1( u1_u8_u6_n122 ) , .A2( u1_u8_u6_n129 ) );
  NAND2_X1 u1_u8_u6_U17 (.ZN( u1_u8_u6_n124 ) , .A2( u1_u8_u6_n146 ) , .A1( u1_u8_u6_n148 ) );
  INV_X1 u1_u8_u6_U18 (.A( u1_u8_u6_n132 ) , .ZN( u1_u8_u6_n171 ) );
  AND2_X1 u1_u8_u6_U19 (.A1( u1_u8_u6_n100 ) , .ZN( u1_u8_u6_n130 ) , .A2( u1_u8_u6_n147 ) );
  INV_X1 u1_u8_u6_U20 (.A( u1_u8_u6_n127 ) , .ZN( u1_u8_u6_n173 ) );
  INV_X1 u1_u8_u6_U21 (.A( u1_u8_u6_n121 ) , .ZN( u1_u8_u6_n167 ) );
  INV_X1 u1_u8_u6_U22 (.A( u1_u8_u6_n100 ) , .ZN( u1_u8_u6_n169 ) );
  INV_X1 u1_u8_u6_U23 (.A( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n170 ) );
  INV_X1 u1_u8_u6_U24 (.A( u1_u8_u6_n113 ) , .ZN( u1_u8_u6_n168 ) );
  AND2_X1 u1_u8_u6_U25 (.A1( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n119 ) , .ZN( u1_u8_u6_n133 ) );
  AND2_X1 u1_u8_u6_U26 (.A2( u1_u8_u6_n121 ) , .A1( u1_u8_u6_n122 ) , .ZN( u1_u8_u6_n131 ) );
  AND3_X1 u1_u8_u6_U27 (.ZN( u1_u8_u6_n120 ) , .A2( u1_u8_u6_n127 ) , .A1( u1_u8_u6_n132 ) , .A3( u1_u8_u6_n145 ) );
  INV_X1 u1_u8_u6_U28 (.A( u1_u8_u6_n146 ) , .ZN( u1_u8_u6_n163 ) );
  AOI222_X1 u1_u8_u6_U29 (.ZN( u1_u8_u6_n114 ) , .A1( u1_u8_u6_n118 ) , .A2( u1_u8_u6_n126 ) , .B2( u1_u8_u6_n151 ) , .C2( u1_u8_u6_n159 ) , .C1( u1_u8_u6_n168 ) , .B1( u1_u8_u6_n169 ) );
  INV_X1 u1_u8_u6_U3 (.A( u1_u8_u6_n110 ) , .ZN( u1_u8_u6_n166 ) );
  NOR2_X1 u1_u8_u6_U30 (.A1( u1_u8_u6_n162 ) , .A2( u1_u8_u6_n165 ) , .ZN( u1_u8_u6_n98 ) );
  AOI211_X1 u1_u8_u6_U31 (.B( u1_u8_u6_n134 ) , .A( u1_u8_u6_n135 ) , .C1( u1_u8_u6_n136 ) , .ZN( u1_u8_u6_n137 ) , .C2( u1_u8_u6_n151 ) );
  AOI21_X1 u1_u8_u6_U32 (.B2( u1_u8_u6_n132 ) , .B1( u1_u8_u6_n133 ) , .ZN( u1_u8_u6_n134 ) , .A( u1_u8_u6_n158 ) );
  NAND4_X1 u1_u8_u6_U33 (.A4( u1_u8_u6_n127 ) , .A3( u1_u8_u6_n128 ) , .A2( u1_u8_u6_n129 ) , .A1( u1_u8_u6_n130 ) , .ZN( u1_u8_u6_n136 ) );
  AOI21_X1 u1_u8_u6_U34 (.B1( u1_u8_u6_n131 ) , .ZN( u1_u8_u6_n135 ) , .A( u1_u8_u6_n144 ) , .B2( u1_u8_u6_n146 ) );
  NAND2_X1 u1_u8_u6_U35 (.A1( u1_u8_u6_n144 ) , .ZN( u1_u8_u6_n151 ) , .A2( u1_u8_u6_n158 ) );
  NAND2_X1 u1_u8_u6_U36 (.ZN( u1_u8_u6_n132 ) , .A1( u1_u8_u6_n91 ) , .A2( u1_u8_u6_n97 ) );
  AOI22_X1 u1_u8_u6_U37 (.B2( u1_u8_u6_n110 ) , .B1( u1_u8_u6_n111 ) , .A1( u1_u8_u6_n112 ) , .ZN( u1_u8_u6_n115 ) , .A2( u1_u8_u6_n161 ) );
  NAND4_X1 u1_u8_u6_U38 (.A3( u1_u8_u6_n109 ) , .ZN( u1_u8_u6_n112 ) , .A4( u1_u8_u6_n132 ) , .A2( u1_u8_u6_n147 ) , .A1( u1_u8_u6_n166 ) );
  NOR2_X1 u1_u8_u6_U39 (.ZN( u1_u8_u6_n109 ) , .A1( u1_u8_u6_n170 ) , .A2( u1_u8_u6_n173 ) );
  INV_X1 u1_u8_u6_U4 (.A( u1_u8_u6_n142 ) , .ZN( u1_u8_u6_n174 ) );
  NOR2_X1 u1_u8_u6_U40 (.A2( u1_u8_u6_n126 ) , .ZN( u1_u8_u6_n155 ) , .A1( u1_u8_u6_n160 ) );
  NAND2_X1 u1_u8_u6_U41 (.ZN( u1_u8_u6_n146 ) , .A2( u1_u8_u6_n94 ) , .A1( u1_u8_u6_n99 ) );
  AOI21_X1 u1_u8_u6_U42 (.A( u1_u8_u6_n144 ) , .B2( u1_u8_u6_n145 ) , .B1( u1_u8_u6_n146 ) , .ZN( u1_u8_u6_n150 ) );
  INV_X1 u1_u8_u6_U43 (.A( u1_u8_u6_n111 ) , .ZN( u1_u8_u6_n158 ) );
  NAND2_X1 u1_u8_u6_U44 (.ZN( u1_u8_u6_n127 ) , .A1( u1_u8_u6_n91 ) , .A2( u1_u8_u6_n92 ) );
  NAND2_X1 u1_u8_u6_U45 (.ZN( u1_u8_u6_n129 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n96 ) );
  INV_X1 u1_u8_u6_U46 (.A( u1_u8_u6_n144 ) , .ZN( u1_u8_u6_n159 ) );
  NAND2_X1 u1_u8_u6_U47 (.ZN( u1_u8_u6_n145 ) , .A2( u1_u8_u6_n97 ) , .A1( u1_u8_u6_n98 ) );
  NAND2_X1 u1_u8_u6_U48 (.ZN( u1_u8_u6_n148 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n94 ) );
  NAND2_X1 u1_u8_u6_U49 (.ZN( u1_u8_u6_n108 ) , .A2( u1_u8_u6_n139 ) , .A1( u1_u8_u6_n144 ) );
  NAND2_X1 u1_u8_u6_U5 (.A2( u1_u8_u6_n143 ) , .ZN( u1_u8_u6_n152 ) , .A1( u1_u8_u6_n166 ) );
  NAND2_X1 u1_u8_u6_U50 (.ZN( u1_u8_u6_n121 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n97 ) );
  NAND2_X1 u1_u8_u6_U51 (.ZN( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n95 ) );
  AND2_X1 u1_u8_u6_U52 (.ZN( u1_u8_u6_n118 ) , .A2( u1_u8_u6_n91 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U53 (.ZN( u1_u8_u6_n147 ) , .A2( u1_u8_u6_n98 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U54 (.ZN( u1_u8_u6_n128 ) , .A1( u1_u8_u6_n94 ) , .A2( u1_u8_u6_n96 ) );
  NAND2_X1 u1_u8_u6_U55 (.ZN( u1_u8_u6_n119 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U56 (.ZN( u1_u8_u6_n123 ) , .A2( u1_u8_u6_n91 ) , .A1( u1_u8_u6_n96 ) );
  NAND2_X1 u1_u8_u6_U57 (.ZN( u1_u8_u6_n100 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n98 ) );
  NAND2_X1 u1_u8_u6_U58 (.ZN( u1_u8_u6_n122 ) , .A1( u1_u8_u6_n94 ) , .A2( u1_u8_u6_n97 ) );
  INV_X1 u1_u8_u6_U59 (.A( u1_u8_u6_n139 ) , .ZN( u1_u8_u6_n160 ) );
  AOI22_X1 u1_u8_u6_U6 (.B2( u1_u8_u6_n101 ) , .A1( u1_u8_u6_n102 ) , .ZN( u1_u8_u6_n103 ) , .B1( u1_u8_u6_n160 ) , .A2( u1_u8_u6_n161 ) );
  NAND2_X1 u1_u8_u6_U60 (.ZN( u1_u8_u6_n113 ) , .A1( u1_u8_u6_n96 ) , .A2( u1_u8_u6_n98 ) );
  NOR2_X1 u1_u8_u6_U61 (.A2( u1_u8_X_40 ) , .A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n126 ) );
  NOR2_X1 u1_u8_u6_U62 (.A2( u1_u8_X_39 ) , .A1( u1_u8_X_42 ) , .ZN( u1_u8_u6_n92 ) );
  NOR2_X1 u1_u8_u6_U63 (.A2( u1_u8_X_39 ) , .A1( u1_u8_u6_n156 ) , .ZN( u1_u8_u6_n97 ) );
  NOR2_X1 u1_u8_u6_U64 (.A2( u1_u8_X_38 ) , .A1( u1_u8_u6_n165 ) , .ZN( u1_u8_u6_n95 ) );
  NOR2_X1 u1_u8_u6_U65 (.A2( u1_u8_X_41 ) , .ZN( u1_u8_u6_n111 ) , .A1( u1_u8_u6_n157 ) );
  NOR2_X1 u1_u8_u6_U66 (.A2( u1_u8_X_37 ) , .A1( u1_u8_u6_n162 ) , .ZN( u1_u8_u6_n94 ) );
  NOR2_X1 u1_u8_u6_U67 (.A2( u1_u8_X_37 ) , .A1( u1_u8_X_38 ) , .ZN( u1_u8_u6_n91 ) );
  NAND2_X1 u1_u8_u6_U68 (.A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n144 ) , .A2( u1_u8_u6_n157 ) );
  NAND2_X1 u1_u8_u6_U69 (.A2( u1_u8_X_40 ) , .A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n139 ) );
  NOR2_X1 u1_u8_u6_U7 (.A1( u1_u8_u6_n118 ) , .ZN( u1_u8_u6_n143 ) , .A2( u1_u8_u6_n168 ) );
  AND2_X1 u1_u8_u6_U70 (.A1( u1_u8_X_39 ) , .A2( u1_u8_u6_n156 ) , .ZN( u1_u8_u6_n96 ) );
  AND2_X1 u1_u8_u6_U71 (.A1( u1_u8_X_39 ) , .A2( u1_u8_X_42 ) , .ZN( u1_u8_u6_n99 ) );
  INV_X1 u1_u8_u6_U72 (.A( u1_u8_X_40 ) , .ZN( u1_u8_u6_n157 ) );
  INV_X1 u1_u8_u6_U73 (.A( u1_u8_X_37 ) , .ZN( u1_u8_u6_n165 ) );
  INV_X1 u1_u8_u6_U74 (.A( u1_u8_X_38 ) , .ZN( u1_u8_u6_n162 ) );
  INV_X1 u1_u8_u6_U75 (.A( u1_u8_X_42 ) , .ZN( u1_u8_u6_n156 ) );
  NAND4_X1 u1_u8_u6_U76 (.ZN( u1_out8_12 ) , .A4( u1_u8_u6_n114 ) , .A3( u1_u8_u6_n115 ) , .A2( u1_u8_u6_n116 ) , .A1( u1_u8_u6_n117 ) );
  OAI22_X1 u1_u8_u6_U77 (.B2( u1_u8_u6_n111 ) , .ZN( u1_u8_u6_n116 ) , .B1( u1_u8_u6_n126 ) , .A2( u1_u8_u6_n164 ) , .A1( u1_u8_u6_n167 ) );
  OAI21_X1 u1_u8_u6_U78 (.A( u1_u8_u6_n108 ) , .ZN( u1_u8_u6_n117 ) , .B2( u1_u8_u6_n141 ) , .B1( u1_u8_u6_n163 ) );
  NAND4_X1 u1_u8_u6_U79 (.ZN( u1_out8_32 ) , .A4( u1_u8_u6_n103 ) , .A3( u1_u8_u6_n104 ) , .A2( u1_u8_u6_n105 ) , .A1( u1_u8_u6_n106 ) );
  OAI21_X1 u1_u8_u6_U8 (.A( u1_u8_u6_n159 ) , .B1( u1_u8_u6_n169 ) , .B2( u1_u8_u6_n173 ) , .ZN( u1_u8_u6_n90 ) );
  AOI22_X1 u1_u8_u6_U80 (.ZN( u1_u8_u6_n105 ) , .A2( u1_u8_u6_n108 ) , .A1( u1_u8_u6_n118 ) , .B2( u1_u8_u6_n126 ) , .B1( u1_u8_u6_n171 ) );
  AOI22_X1 u1_u8_u6_U81 (.ZN( u1_u8_u6_n104 ) , .A1( u1_u8_u6_n111 ) , .B1( u1_u8_u6_n124 ) , .B2( u1_u8_u6_n151 ) , .A2( u1_u8_u6_n93 ) );
  OAI211_X1 u1_u8_u6_U82 (.ZN( u1_out8_7 ) , .B( u1_u8_u6_n153 ) , .C2( u1_u8_u6_n154 ) , .C1( u1_u8_u6_n155 ) , .A( u1_u8_u6_n174 ) );
  NOR3_X1 u1_u8_u6_U83 (.A1( u1_u8_u6_n141 ) , .ZN( u1_u8_u6_n154 ) , .A3( u1_u8_u6_n164 ) , .A2( u1_u8_u6_n171 ) );
  AOI211_X1 u1_u8_u6_U84 (.B( u1_u8_u6_n149 ) , .A( u1_u8_u6_n150 ) , .C2( u1_u8_u6_n151 ) , .C1( u1_u8_u6_n152 ) , .ZN( u1_u8_u6_n153 ) );
  OAI211_X1 u1_u8_u6_U85 (.ZN( u1_out8_22 ) , .B( u1_u8_u6_n137 ) , .A( u1_u8_u6_n138 ) , .C2( u1_u8_u6_n139 ) , .C1( u1_u8_u6_n140 ) );
  AOI22_X1 u1_u8_u6_U86 (.B1( u1_u8_u6_n124 ) , .A2( u1_u8_u6_n125 ) , .A1( u1_u8_u6_n126 ) , .ZN( u1_u8_u6_n138 ) , .B2( u1_u8_u6_n161 ) );
  AND4_X1 u1_u8_u6_U87 (.A3( u1_u8_u6_n119 ) , .A1( u1_u8_u6_n120 ) , .A4( u1_u8_u6_n129 ) , .ZN( u1_u8_u6_n140 ) , .A2( u1_u8_u6_n143 ) );
  NAND3_X1 u1_u8_u6_U88 (.A2( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n125 ) , .A1( u1_u8_u6_n130 ) , .A3( u1_u8_u6_n131 ) );
  NAND3_X1 u1_u8_u6_U89 (.A3( u1_u8_u6_n133 ) , .ZN( u1_u8_u6_n141 ) , .A1( u1_u8_u6_n145 ) , .A2( u1_u8_u6_n148 ) );
  INV_X1 u1_u8_u6_U9 (.ZN( u1_u8_u6_n172 ) , .A( u1_u8_u6_n88 ) );
  NAND3_X1 u1_u8_u6_U90 (.ZN( u1_u8_u6_n101 ) , .A3( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n121 ) , .A1( u1_u8_u6_n127 ) );
  NAND3_X1 u1_u8_u6_U91 (.ZN( u1_u8_u6_n102 ) , .A3( u1_u8_u6_n130 ) , .A2( u1_u8_u6_n145 ) , .A1( u1_u8_u6_n166 ) );
  NAND3_X1 u1_u8_u6_U92 (.A3( u1_u8_u6_n113 ) , .A1( u1_u8_u6_n119 ) , .A2( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n93 ) );
  NAND3_X1 u1_u8_u6_U93 (.ZN( u1_u8_u6_n142 ) , .A2( u1_u8_u6_n172 ) , .A3( u1_u8_u6_n89 ) , .A1( u1_u8_u6_n90 ) );
  AND3_X1 u1_u8_u7_U10 (.A3( u1_u8_u7_n110 ) , .A2( u1_u8_u7_n127 ) , .A1( u1_u8_u7_n132 ) , .ZN( u1_u8_u7_n92 ) );
  OAI21_X1 u1_u8_u7_U11 (.A( u1_u8_u7_n161 ) , .B1( u1_u8_u7_n168 ) , .B2( u1_u8_u7_n173 ) , .ZN( u1_u8_u7_n91 ) );
  AOI211_X1 u1_u8_u7_U12 (.A( u1_u8_u7_n117 ) , .ZN( u1_u8_u7_n118 ) , .C2( u1_u8_u7_n126 ) , .C1( u1_u8_u7_n177 ) , .B( u1_u8_u7_n180 ) );
  OAI22_X1 u1_u8_u7_U13 (.B1( u1_u8_u7_n115 ) , .ZN( u1_u8_u7_n117 ) , .A2( u1_u8_u7_n133 ) , .A1( u1_u8_u7_n137 ) , .B2( u1_u8_u7_n162 ) );
  INV_X1 u1_u8_u7_U14 (.A( u1_u8_u7_n116 ) , .ZN( u1_u8_u7_n180 ) );
  NOR3_X1 u1_u8_u7_U15 (.ZN( u1_u8_u7_n115 ) , .A3( u1_u8_u7_n145 ) , .A2( u1_u8_u7_n168 ) , .A1( u1_u8_u7_n169 ) );
  OAI211_X1 u1_u8_u7_U16 (.B( u1_u8_u7_n122 ) , .A( u1_u8_u7_n123 ) , .C2( u1_u8_u7_n124 ) , .ZN( u1_u8_u7_n154 ) , .C1( u1_u8_u7_n162 ) );
  AOI222_X1 u1_u8_u7_U17 (.ZN( u1_u8_u7_n122 ) , .C2( u1_u8_u7_n126 ) , .C1( u1_u8_u7_n145 ) , .B1( u1_u8_u7_n161 ) , .A2( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n170 ) , .A1( u1_u8_u7_n176 ) );
  INV_X1 u1_u8_u7_U18 (.A( u1_u8_u7_n133 ) , .ZN( u1_u8_u7_n176 ) );
  NOR3_X1 u1_u8_u7_U19 (.A2( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n135 ) , .ZN( u1_u8_u7_n136 ) , .A3( u1_u8_u7_n171 ) );
  NOR2_X1 u1_u8_u7_U20 (.A1( u1_u8_u7_n130 ) , .A2( u1_u8_u7_n134 ) , .ZN( u1_u8_u7_n153 ) );
  INV_X1 u1_u8_u7_U21 (.A( u1_u8_u7_n101 ) , .ZN( u1_u8_u7_n165 ) );
  NOR2_X1 u1_u8_u7_U22 (.ZN( u1_u8_u7_n111 ) , .A2( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n169 ) );
  AOI21_X1 u1_u8_u7_U23 (.ZN( u1_u8_u7_n104 ) , .B2( u1_u8_u7_n112 ) , .B1( u1_u8_u7_n127 ) , .A( u1_u8_u7_n164 ) );
  AOI21_X1 u1_u8_u7_U24 (.ZN( u1_u8_u7_n106 ) , .B1( u1_u8_u7_n133 ) , .B2( u1_u8_u7_n146 ) , .A( u1_u8_u7_n162 ) );
  AOI21_X1 u1_u8_u7_U25 (.A( u1_u8_u7_n101 ) , .ZN( u1_u8_u7_n107 ) , .B2( u1_u8_u7_n128 ) , .B1( u1_u8_u7_n175 ) );
  INV_X1 u1_u8_u7_U26 (.A( u1_u8_u7_n138 ) , .ZN( u1_u8_u7_n171 ) );
  INV_X1 u1_u8_u7_U27 (.A( u1_u8_u7_n131 ) , .ZN( u1_u8_u7_n177 ) );
  INV_X1 u1_u8_u7_U28 (.A( u1_u8_u7_n110 ) , .ZN( u1_u8_u7_n174 ) );
  NAND2_X1 u1_u8_u7_U29 (.A1( u1_u8_u7_n129 ) , .A2( u1_u8_u7_n132 ) , .ZN( u1_u8_u7_n149 ) );
  OAI21_X1 u1_u8_u7_U3 (.ZN( u1_u8_u7_n159 ) , .A( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n171 ) , .B1( u1_u8_u7_n174 ) );
  NAND2_X1 u1_u8_u7_U30 (.A1( u1_u8_u7_n113 ) , .A2( u1_u8_u7_n124 ) , .ZN( u1_u8_u7_n130 ) );
  INV_X1 u1_u8_u7_U31 (.A( u1_u8_u7_n112 ) , .ZN( u1_u8_u7_n173 ) );
  INV_X1 u1_u8_u7_U32 (.A( u1_u8_u7_n128 ) , .ZN( u1_u8_u7_n168 ) );
  INV_X1 u1_u8_u7_U33 (.A( u1_u8_u7_n148 ) , .ZN( u1_u8_u7_n169 ) );
  INV_X1 u1_u8_u7_U34 (.A( u1_u8_u7_n127 ) , .ZN( u1_u8_u7_n179 ) );
  NOR2_X1 u1_u8_u7_U35 (.ZN( u1_u8_u7_n101 ) , .A2( u1_u8_u7_n150 ) , .A1( u1_u8_u7_n156 ) );
  AOI211_X1 u1_u8_u7_U36 (.B( u1_u8_u7_n154 ) , .A( u1_u8_u7_n155 ) , .C1( u1_u8_u7_n156 ) , .ZN( u1_u8_u7_n157 ) , .C2( u1_u8_u7_n172 ) );
  INV_X1 u1_u8_u7_U37 (.A( u1_u8_u7_n153 ) , .ZN( u1_u8_u7_n172 ) );
  AOI211_X1 u1_u8_u7_U38 (.B( u1_u8_u7_n139 ) , .A( u1_u8_u7_n140 ) , .C2( u1_u8_u7_n141 ) , .ZN( u1_u8_u7_n142 ) , .C1( u1_u8_u7_n156 ) );
  NAND4_X1 u1_u8_u7_U39 (.A3( u1_u8_u7_n127 ) , .A2( u1_u8_u7_n128 ) , .A1( u1_u8_u7_n129 ) , .ZN( u1_u8_u7_n141 ) , .A4( u1_u8_u7_n147 ) );
  INV_X1 u1_u8_u7_U4 (.A( u1_u8_u7_n111 ) , .ZN( u1_u8_u7_n170 ) );
  AOI21_X1 u1_u8_u7_U40 (.A( u1_u8_u7_n137 ) , .B1( u1_u8_u7_n138 ) , .ZN( u1_u8_u7_n139 ) , .B2( u1_u8_u7_n146 ) );
  OAI22_X1 u1_u8_u7_U41 (.B1( u1_u8_u7_n136 ) , .ZN( u1_u8_u7_n140 ) , .A1( u1_u8_u7_n153 ) , .B2( u1_u8_u7_n162 ) , .A2( u1_u8_u7_n164 ) );
  AOI21_X1 u1_u8_u7_U42 (.ZN( u1_u8_u7_n123 ) , .B1( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n177 ) , .A( u1_u8_u7_n97 ) );
  AOI21_X1 u1_u8_u7_U43 (.B2( u1_u8_u7_n113 ) , .B1( u1_u8_u7_n124 ) , .A( u1_u8_u7_n125 ) , .ZN( u1_u8_u7_n97 ) );
  INV_X1 u1_u8_u7_U44 (.A( u1_u8_u7_n125 ) , .ZN( u1_u8_u7_n161 ) );
  INV_X1 u1_u8_u7_U45 (.A( u1_u8_u7_n152 ) , .ZN( u1_u8_u7_n162 ) );
  AOI22_X1 u1_u8_u7_U46 (.A2( u1_u8_u7_n114 ) , .ZN( u1_u8_u7_n119 ) , .B1( u1_u8_u7_n130 ) , .A1( u1_u8_u7_n156 ) , .B2( u1_u8_u7_n165 ) );
  NAND2_X1 u1_u8_u7_U47 (.A2( u1_u8_u7_n112 ) , .ZN( u1_u8_u7_n114 ) , .A1( u1_u8_u7_n175 ) );
  AND2_X1 u1_u8_u7_U48 (.ZN( u1_u8_u7_n145 ) , .A2( u1_u8_u7_n98 ) , .A1( u1_u8_u7_n99 ) );
  NOR2_X1 u1_u8_u7_U49 (.ZN( u1_u8_u7_n137 ) , .A1( u1_u8_u7_n150 ) , .A2( u1_u8_u7_n161 ) );
  INV_X1 u1_u8_u7_U5 (.A( u1_u8_u7_n149 ) , .ZN( u1_u8_u7_n175 ) );
  AOI21_X1 u1_u8_u7_U50 (.ZN( u1_u8_u7_n105 ) , .B2( u1_u8_u7_n110 ) , .A( u1_u8_u7_n125 ) , .B1( u1_u8_u7_n147 ) );
  NAND2_X1 u1_u8_u7_U51 (.ZN( u1_u8_u7_n146 ) , .A1( u1_u8_u7_n95 ) , .A2( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U52 (.A2( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n147 ) , .A1( u1_u8_u7_n93 ) );
  NAND2_X1 u1_u8_u7_U53 (.A1( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n127 ) , .A2( u1_u8_u7_n99 ) );
  OR2_X1 u1_u8_u7_U54 (.ZN( u1_u8_u7_n126 ) , .A2( u1_u8_u7_n152 ) , .A1( u1_u8_u7_n156 ) );
  NAND2_X1 u1_u8_u7_U55 (.A2( u1_u8_u7_n102 ) , .A1( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n133 ) );
  NAND2_X1 u1_u8_u7_U56 (.ZN( u1_u8_u7_n112 ) , .A2( u1_u8_u7_n96 ) , .A1( u1_u8_u7_n99 ) );
  NAND2_X1 u1_u8_u7_U57 (.A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n128 ) , .A1( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U58 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n113 ) , .A2( u1_u8_u7_n93 ) );
  NAND2_X1 u1_u8_u7_U59 (.A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n124 ) , .A1( u1_u8_u7_n96 ) );
  INV_X1 u1_u8_u7_U6 (.A( u1_u8_u7_n154 ) , .ZN( u1_u8_u7_n178 ) );
  NAND2_X1 u1_u8_u7_U60 (.ZN( u1_u8_u7_n110 ) , .A1( u1_u8_u7_n95 ) , .A2( u1_u8_u7_n96 ) );
  INV_X1 u1_u8_u7_U61 (.A( u1_u8_u7_n150 ) , .ZN( u1_u8_u7_n164 ) );
  AND2_X1 u1_u8_u7_U62 (.ZN( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n93 ) , .A2( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U63 (.A1( u1_u8_u7_n100 ) , .A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n129 ) );
  NAND2_X1 u1_u8_u7_U64 (.A2( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n131 ) , .A1( u1_u8_u7_n95 ) );
  NAND2_X1 u1_u8_u7_U65 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n138 ) , .A2( u1_u8_u7_n99 ) );
  NAND2_X1 u1_u8_u7_U66 (.ZN( u1_u8_u7_n132 ) , .A1( u1_u8_u7_n93 ) , .A2( u1_u8_u7_n96 ) );
  NAND2_X1 u1_u8_u7_U67 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n148 ) , .A2( u1_u8_u7_n95 ) );
  NOR2_X1 u1_u8_u7_U68 (.A2( u1_u8_X_47 ) , .ZN( u1_u8_u7_n150 ) , .A1( u1_u8_u7_n163 ) );
  NOR2_X1 u1_u8_u7_U69 (.A2( u1_u8_X_43 ) , .A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n103 ) );
  AOI211_X1 u1_u8_u7_U7 (.ZN( u1_u8_u7_n116 ) , .A( u1_u8_u7_n155 ) , .C1( u1_u8_u7_n161 ) , .C2( u1_u8_u7_n171 ) , .B( u1_u8_u7_n94 ) );
  NOR2_X1 u1_u8_u7_U70 (.A2( u1_u8_X_48 ) , .A1( u1_u8_u7_n166 ) , .ZN( u1_u8_u7_n95 ) );
  NOR2_X1 u1_u8_u7_U71 (.A2( u1_u8_X_45 ) , .A1( u1_u8_X_48 ) , .ZN( u1_u8_u7_n99 ) );
  NOR2_X1 u1_u8_u7_U72 (.A2( u1_u8_X_44 ) , .A1( u1_u8_u7_n167 ) , .ZN( u1_u8_u7_n98 ) );
  NOR2_X1 u1_u8_u7_U73 (.A2( u1_u8_X_46 ) , .A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n152 ) );
  AND2_X1 u1_u8_u7_U74 (.A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n156 ) , .A2( u1_u8_u7_n163 ) );
  NAND2_X1 u1_u8_u7_U75 (.A2( u1_u8_X_46 ) , .A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n125 ) );
  AND2_X1 u1_u8_u7_U76 (.A2( u1_u8_X_45 ) , .A1( u1_u8_X_48 ) , .ZN( u1_u8_u7_n102 ) );
  AND2_X1 u1_u8_u7_U77 (.A2( u1_u8_X_43 ) , .A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n96 ) );
  AND2_X1 u1_u8_u7_U78 (.A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n100 ) , .A2( u1_u8_u7_n167 ) );
  AND2_X1 u1_u8_u7_U79 (.A1( u1_u8_X_48 ) , .A2( u1_u8_u7_n166 ) , .ZN( u1_u8_u7_n93 ) );
  OAI222_X1 u1_u8_u7_U8 (.C2( u1_u8_u7_n101 ) , .B2( u1_u8_u7_n111 ) , .A1( u1_u8_u7_n113 ) , .C1( u1_u8_u7_n146 ) , .A2( u1_u8_u7_n162 ) , .B1( u1_u8_u7_n164 ) , .ZN( u1_u8_u7_n94 ) );
  INV_X1 u1_u8_u7_U80 (.A( u1_u8_X_46 ) , .ZN( u1_u8_u7_n163 ) );
  INV_X1 u1_u8_u7_U81 (.A( u1_u8_X_43 ) , .ZN( u1_u8_u7_n167 ) );
  INV_X1 u1_u8_u7_U82 (.A( u1_u8_X_45 ) , .ZN( u1_u8_u7_n166 ) );
  NAND4_X1 u1_u8_u7_U83 (.ZN( u1_out8_5 ) , .A4( u1_u8_u7_n108 ) , .A3( u1_u8_u7_n109 ) , .A1( u1_u8_u7_n116 ) , .A2( u1_u8_u7_n123 ) );
  AOI22_X1 u1_u8_u7_U84 (.ZN( u1_u8_u7_n109 ) , .A2( u1_u8_u7_n126 ) , .B2( u1_u8_u7_n145 ) , .B1( u1_u8_u7_n156 ) , .A1( u1_u8_u7_n171 ) );
  NOR4_X1 u1_u8_u7_U85 (.A4( u1_u8_u7_n104 ) , .A3( u1_u8_u7_n105 ) , .A2( u1_u8_u7_n106 ) , .A1( u1_u8_u7_n107 ) , .ZN( u1_u8_u7_n108 ) );
  NAND4_X1 u1_u8_u7_U86 (.ZN( u1_out8_27 ) , .A4( u1_u8_u7_n118 ) , .A3( u1_u8_u7_n119 ) , .A2( u1_u8_u7_n120 ) , .A1( u1_u8_u7_n121 ) );
  OAI21_X1 u1_u8_u7_U87 (.ZN( u1_u8_u7_n121 ) , .B2( u1_u8_u7_n145 ) , .A( u1_u8_u7_n150 ) , .B1( u1_u8_u7_n174 ) );
  OAI21_X1 u1_u8_u7_U88 (.ZN( u1_u8_u7_n120 ) , .A( u1_u8_u7_n161 ) , .B2( u1_u8_u7_n170 ) , .B1( u1_u8_u7_n179 ) );
  NAND4_X1 u1_u8_u7_U89 (.ZN( u1_out8_21 ) , .A4( u1_u8_u7_n157 ) , .A3( u1_u8_u7_n158 ) , .A2( u1_u8_u7_n159 ) , .A1( u1_u8_u7_n160 ) );
  OAI221_X1 u1_u8_u7_U9 (.C1( u1_u8_u7_n101 ) , .C2( u1_u8_u7_n147 ) , .ZN( u1_u8_u7_n155 ) , .B2( u1_u8_u7_n162 ) , .A( u1_u8_u7_n91 ) , .B1( u1_u8_u7_n92 ) );
  OAI21_X1 u1_u8_u7_U90 (.B1( u1_u8_u7_n145 ) , .ZN( u1_u8_u7_n160 ) , .A( u1_u8_u7_n161 ) , .B2( u1_u8_u7_n177 ) );
  AOI22_X1 u1_u8_u7_U91 (.B2( u1_u8_u7_n149 ) , .B1( u1_u8_u7_n150 ) , .A2( u1_u8_u7_n151 ) , .A1( u1_u8_u7_n152 ) , .ZN( u1_u8_u7_n158 ) );
  NAND4_X1 u1_u8_u7_U92 (.ZN( u1_out8_15 ) , .A4( u1_u8_u7_n142 ) , .A3( u1_u8_u7_n143 ) , .A2( u1_u8_u7_n144 ) , .A1( u1_u8_u7_n178 ) );
  OR2_X1 u1_u8_u7_U93 (.A2( u1_u8_u7_n125 ) , .A1( u1_u8_u7_n129 ) , .ZN( u1_u8_u7_n144 ) );
  AOI22_X1 u1_u8_u7_U94 (.A2( u1_u8_u7_n126 ) , .ZN( u1_u8_u7_n143 ) , .B2( u1_u8_u7_n165 ) , .B1( u1_u8_u7_n173 ) , .A1( u1_u8_u7_n174 ) );
  NAND3_X1 u1_u8_u7_U95 (.A3( u1_u8_u7_n146 ) , .A2( u1_u8_u7_n147 ) , .A1( u1_u8_u7_n148 ) , .ZN( u1_u8_u7_n151 ) );
  NAND3_X1 u1_u8_u7_U96 (.A3( u1_u8_u7_n131 ) , .A2( u1_u8_u7_n132 ) , .A1( u1_u8_u7_n133 ) , .ZN( u1_u8_u7_n135 ) );
  XOR2_X1 u1_u9_U11 (.B( u1_K10_44 ) , .A( u1_R8_29 ) , .Z( u1_u9_X_44 ) );
  XOR2_X1 u1_u9_U12 (.B( u1_K10_43 ) , .A( u1_R8_28 ) , .Z( u1_u9_X_43 ) );
  XOR2_X1 u1_u9_U13 (.B( u1_K10_42 ) , .A( u1_R8_29 ) , .Z( u1_u9_X_42 ) );
  XOR2_X1 u1_u9_U14 (.B( u1_K10_41 ) , .A( u1_R8_28 ) , .Z( u1_u9_X_41 ) );
  XOR2_X1 u1_u9_U18 (.B( u1_K10_38 ) , .A( u1_R8_25 ) , .Z( u1_u9_X_38 ) );
  XOR2_X1 u1_u9_U19 (.B( u1_K10_37 ) , .A( u1_R8_24 ) , .Z( u1_u9_X_37 ) );
  XOR2_X1 u1_u9_U20 (.B( u1_K10_36 ) , .A( u1_R8_25 ) , .Z( u1_u9_X_36 ) );
  XOR2_X1 u1_u9_U21 (.B( u1_K10_35 ) , .A( u1_R8_24 ) , .Z( u1_u9_X_35 ) );
  XOR2_X1 u1_u9_U23 (.B( u1_K10_33 ) , .A( u1_R8_22 ) , .Z( u1_u9_X_33 ) );
  XOR2_X1 u1_u9_U24 (.B( u1_K10_32 ) , .A( u1_R8_21 ) , .Z( u1_u9_X_32 ) );
  XOR2_X1 u1_u9_U25 (.B( u1_K10_31 ) , .A( u1_R8_20 ) , .Z( u1_u9_X_31 ) );
  XOR2_X1 u1_u9_U7 (.B( u1_K10_48 ) , .A( u1_R8_1 ) , .Z( u1_u9_X_48 ) );
  XOR2_X1 u1_u9_U8 (.B( u1_K10_47 ) , .A( u1_R8_32 ) , .Z( u1_u9_X_47 ) );
  NOR2_X1 u1_u9_u5_U10 (.ZN( u1_u9_u5_n135 ) , .A1( u1_u9_u5_n173 ) , .A2( u1_u9_u5_n176 ) );
  NOR3_X1 u1_u9_u5_U100 (.A3( u1_u9_u5_n141 ) , .A1( u1_u9_u5_n142 ) , .ZN( u1_u9_u5_n143 ) , .A2( u1_u9_u5_n191 ) );
  NAND4_X1 u1_u9_u5_U101 (.ZN( u1_out9_4 ) , .A4( u1_u9_u5_n112 ) , .A2( u1_u9_u5_n113 ) , .A1( u1_u9_u5_n114 ) , .A3( u1_u9_u5_n195 ) );
  AOI211_X1 u1_u9_u5_U102 (.A( u1_u9_u5_n110 ) , .C1( u1_u9_u5_n111 ) , .ZN( u1_u9_u5_n112 ) , .B( u1_u9_u5_n118 ) , .C2( u1_u9_u5_n177 ) );
  INV_X1 u1_u9_u5_U103 (.A( u1_u9_u5_n102 ) , .ZN( u1_u9_u5_n195 ) );
  NAND3_X1 u1_u9_u5_U104 (.A2( u1_u9_u5_n154 ) , .A3( u1_u9_u5_n158 ) , .A1( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n99 ) );
  INV_X1 u1_u9_u5_U11 (.A( u1_u9_u5_n121 ) , .ZN( u1_u9_u5_n177 ) );
  NOR2_X1 u1_u9_u5_U12 (.ZN( u1_u9_u5_n160 ) , .A2( u1_u9_u5_n173 ) , .A1( u1_u9_u5_n177 ) );
  INV_X1 u1_u9_u5_U13 (.A( u1_u9_u5_n150 ) , .ZN( u1_u9_u5_n174 ) );
  AOI21_X1 u1_u9_u5_U14 (.A( u1_u9_u5_n160 ) , .B2( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n162 ) , .B1( u1_u9_u5_n192 ) );
  INV_X1 u1_u9_u5_U15 (.A( u1_u9_u5_n159 ) , .ZN( u1_u9_u5_n192 ) );
  AOI21_X1 u1_u9_u5_U16 (.A( u1_u9_u5_n156 ) , .B2( u1_u9_u5_n157 ) , .B1( u1_u9_u5_n158 ) , .ZN( u1_u9_u5_n163 ) );
  AOI21_X1 u1_u9_u5_U17 (.B2( u1_u9_u5_n139 ) , .B1( u1_u9_u5_n140 ) , .ZN( u1_u9_u5_n141 ) , .A( u1_u9_u5_n150 ) );
  OAI21_X1 u1_u9_u5_U18 (.A( u1_u9_u5_n133 ) , .B2( u1_u9_u5_n134 ) , .B1( u1_u9_u5_n135 ) , .ZN( u1_u9_u5_n142 ) );
  OAI21_X1 u1_u9_u5_U19 (.ZN( u1_u9_u5_n133 ) , .B2( u1_u9_u5_n147 ) , .A( u1_u9_u5_n173 ) , .B1( u1_u9_u5_n188 ) );
  NAND2_X1 u1_u9_u5_U20 (.A2( u1_u9_u5_n119 ) , .A1( u1_u9_u5_n123 ) , .ZN( u1_u9_u5_n137 ) );
  INV_X1 u1_u9_u5_U21 (.A( u1_u9_u5_n155 ) , .ZN( u1_u9_u5_n194 ) );
  NAND2_X1 u1_u9_u5_U22 (.A1( u1_u9_u5_n121 ) , .ZN( u1_u9_u5_n132 ) , .A2( u1_u9_u5_n172 ) );
  NAND2_X1 u1_u9_u5_U23 (.A2( u1_u9_u5_n122 ) , .ZN( u1_u9_u5_n136 ) , .A1( u1_u9_u5_n154 ) );
  NAND2_X1 u1_u9_u5_U24 (.A2( u1_u9_u5_n119 ) , .A1( u1_u9_u5_n120 ) , .ZN( u1_u9_u5_n159 ) );
  INV_X1 u1_u9_u5_U25 (.A( u1_u9_u5_n156 ) , .ZN( u1_u9_u5_n175 ) );
  INV_X1 u1_u9_u5_U26 (.A( u1_u9_u5_n158 ) , .ZN( u1_u9_u5_n188 ) );
  INV_X1 u1_u9_u5_U27 (.A( u1_u9_u5_n152 ) , .ZN( u1_u9_u5_n179 ) );
  INV_X1 u1_u9_u5_U28 (.A( u1_u9_u5_n140 ) , .ZN( u1_u9_u5_n182 ) );
  INV_X1 u1_u9_u5_U29 (.A( u1_u9_u5_n151 ) , .ZN( u1_u9_u5_n183 ) );
  NOR2_X1 u1_u9_u5_U3 (.ZN( u1_u9_u5_n134 ) , .A1( u1_u9_u5_n183 ) , .A2( u1_u9_u5_n190 ) );
  INV_X1 u1_u9_u5_U30 (.A( u1_u9_u5_n123 ) , .ZN( u1_u9_u5_n185 ) );
  INV_X1 u1_u9_u5_U31 (.A( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n184 ) );
  INV_X1 u1_u9_u5_U32 (.A( u1_u9_u5_n139 ) , .ZN( u1_u9_u5_n189 ) );
  INV_X1 u1_u9_u5_U33 (.A( u1_u9_u5_n157 ) , .ZN( u1_u9_u5_n190 ) );
  INV_X1 u1_u9_u5_U34 (.A( u1_u9_u5_n120 ) , .ZN( u1_u9_u5_n193 ) );
  NAND2_X1 u1_u9_u5_U35 (.ZN( u1_u9_u5_n111 ) , .A1( u1_u9_u5_n140 ) , .A2( u1_u9_u5_n155 ) );
  NOR2_X1 u1_u9_u5_U36 (.ZN( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n170 ) , .A2( u1_u9_u5_n180 ) );
  INV_X1 u1_u9_u5_U37 (.A( u1_u9_u5_n117 ) , .ZN( u1_u9_u5_n196 ) );
  OAI221_X1 u1_u9_u5_U38 (.A( u1_u9_u5_n116 ) , .ZN( u1_u9_u5_n117 ) , .B2( u1_u9_u5_n119 ) , .C1( u1_u9_u5_n153 ) , .C2( u1_u9_u5_n158 ) , .B1( u1_u9_u5_n172 ) );
  AOI222_X1 u1_u9_u5_U39 (.ZN( u1_u9_u5_n116 ) , .B2( u1_u9_u5_n145 ) , .C1( u1_u9_u5_n148 ) , .A2( u1_u9_u5_n174 ) , .C2( u1_u9_u5_n177 ) , .B1( u1_u9_u5_n187 ) , .A1( u1_u9_u5_n193 ) );
  INV_X1 u1_u9_u5_U4 (.A( u1_u9_u5_n138 ) , .ZN( u1_u9_u5_n191 ) );
  INV_X1 u1_u9_u5_U40 (.A( u1_u9_u5_n115 ) , .ZN( u1_u9_u5_n187 ) );
  OAI221_X1 u1_u9_u5_U41 (.A( u1_u9_u5_n101 ) , .ZN( u1_u9_u5_n102 ) , .C2( u1_u9_u5_n115 ) , .C1( u1_u9_u5_n126 ) , .B1( u1_u9_u5_n134 ) , .B2( u1_u9_u5_n160 ) );
  OAI21_X1 u1_u9_u5_U42 (.ZN( u1_u9_u5_n101 ) , .B1( u1_u9_u5_n137 ) , .A( u1_u9_u5_n146 ) , .B2( u1_u9_u5_n147 ) );
  AOI22_X1 u1_u9_u5_U43 (.B2( u1_u9_u5_n131 ) , .A2( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n169 ) , .B1( u1_u9_u5_n174 ) , .A1( u1_u9_u5_n185 ) );
  NOR2_X1 u1_u9_u5_U44 (.A1( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n150 ) , .A2( u1_u9_u5_n173 ) );
  AOI21_X1 u1_u9_u5_U45 (.A( u1_u9_u5_n118 ) , .B2( u1_u9_u5_n145 ) , .ZN( u1_u9_u5_n168 ) , .B1( u1_u9_u5_n186 ) );
  INV_X1 u1_u9_u5_U46 (.A( u1_u9_u5_n122 ) , .ZN( u1_u9_u5_n186 ) );
  NOR2_X1 u1_u9_u5_U47 (.A1( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n152 ) , .A2( u1_u9_u5_n176 ) );
  NOR2_X1 u1_u9_u5_U48 (.A1( u1_u9_u5_n115 ) , .ZN( u1_u9_u5_n118 ) , .A2( u1_u9_u5_n153 ) );
  NOR2_X1 u1_u9_u5_U49 (.A2( u1_u9_u5_n145 ) , .ZN( u1_u9_u5_n156 ) , .A1( u1_u9_u5_n174 ) );
  OAI21_X1 u1_u9_u5_U5 (.B2( u1_u9_u5_n136 ) , .B1( u1_u9_u5_n137 ) , .ZN( u1_u9_u5_n138 ) , .A( u1_u9_u5_n177 ) );
  NOR2_X1 u1_u9_u5_U50 (.ZN( u1_u9_u5_n121 ) , .A2( u1_u9_u5_n145 ) , .A1( u1_u9_u5_n176 ) );
  AOI22_X1 u1_u9_u5_U51 (.ZN( u1_u9_u5_n114 ) , .A2( u1_u9_u5_n137 ) , .A1( u1_u9_u5_n145 ) , .B2( u1_u9_u5_n175 ) , .B1( u1_u9_u5_n193 ) );
  OAI211_X1 u1_u9_u5_U52 (.B( u1_u9_u5_n124 ) , .A( u1_u9_u5_n125 ) , .C2( u1_u9_u5_n126 ) , .C1( u1_u9_u5_n127 ) , .ZN( u1_u9_u5_n128 ) );
  NOR3_X1 u1_u9_u5_U53 (.ZN( u1_u9_u5_n127 ) , .A1( u1_u9_u5_n136 ) , .A3( u1_u9_u5_n148 ) , .A2( u1_u9_u5_n182 ) );
  OAI21_X1 u1_u9_u5_U54 (.ZN( u1_u9_u5_n124 ) , .A( u1_u9_u5_n177 ) , .B2( u1_u9_u5_n183 ) , .B1( u1_u9_u5_n189 ) );
  OAI21_X1 u1_u9_u5_U55 (.ZN( u1_u9_u5_n125 ) , .A( u1_u9_u5_n174 ) , .B2( u1_u9_u5_n185 ) , .B1( u1_u9_u5_n190 ) );
  AOI21_X1 u1_u9_u5_U56 (.A( u1_u9_u5_n153 ) , .B2( u1_u9_u5_n154 ) , .B1( u1_u9_u5_n155 ) , .ZN( u1_u9_u5_n164 ) );
  AOI21_X1 u1_u9_u5_U57 (.ZN( u1_u9_u5_n110 ) , .B1( u1_u9_u5_n122 ) , .B2( u1_u9_u5_n139 ) , .A( u1_u9_u5_n153 ) );
  INV_X1 u1_u9_u5_U58 (.A( u1_u9_u5_n153 ) , .ZN( u1_u9_u5_n176 ) );
  INV_X1 u1_u9_u5_U59 (.A( u1_u9_u5_n126 ) , .ZN( u1_u9_u5_n173 ) );
  AOI222_X1 u1_u9_u5_U6 (.ZN( u1_u9_u5_n113 ) , .A1( u1_u9_u5_n131 ) , .C1( u1_u9_u5_n148 ) , .B2( u1_u9_u5_n174 ) , .C2( u1_u9_u5_n178 ) , .A2( u1_u9_u5_n179 ) , .B1( u1_u9_u5_n99 ) );
  AND2_X1 u1_u9_u5_U60 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n147 ) );
  AND2_X1 u1_u9_u5_U61 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n148 ) );
  NAND2_X1 u1_u9_u5_U62 (.A1( u1_u9_u5_n105 ) , .A2( u1_u9_u5_n106 ) , .ZN( u1_u9_u5_n158 ) );
  NAND2_X1 u1_u9_u5_U63 (.A2( u1_u9_u5_n108 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n139 ) );
  NAND2_X1 u1_u9_u5_U64 (.A1( u1_u9_u5_n106 ) , .A2( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n119 ) );
  NAND2_X1 u1_u9_u5_U65 (.A2( u1_u9_u5_n103 ) , .A1( u1_u9_u5_n105 ) , .ZN( u1_u9_u5_n140 ) );
  NAND2_X1 u1_u9_u5_U66 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n105 ) , .ZN( u1_u9_u5_n155 ) );
  NAND2_X1 u1_u9_u5_U67 (.A2( u1_u9_u5_n106 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n122 ) );
  NAND2_X1 u1_u9_u5_U68 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n106 ) , .ZN( u1_u9_u5_n115 ) );
  NAND2_X1 u1_u9_u5_U69 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n103 ) , .ZN( u1_u9_u5_n161 ) );
  INV_X1 u1_u9_u5_U7 (.A( u1_u9_u5_n135 ) , .ZN( u1_u9_u5_n178 ) );
  NAND2_X1 u1_u9_u5_U70 (.A1( u1_u9_u5_n105 ) , .A2( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n154 ) );
  INV_X1 u1_u9_u5_U71 (.A( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n172 ) );
  NAND2_X1 u1_u9_u5_U72 (.A1( u1_u9_u5_n103 ) , .A2( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n123 ) );
  NAND2_X1 u1_u9_u5_U73 (.A2( u1_u9_u5_n103 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n151 ) );
  NAND2_X1 u1_u9_u5_U74 (.A2( u1_u9_u5_n107 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n120 ) );
  NAND2_X1 u1_u9_u5_U75 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n157 ) );
  AND2_X1 u1_u9_u5_U76 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n104 ) , .ZN( u1_u9_u5_n131 ) );
  NOR2_X1 u1_u9_u5_U77 (.A2( u1_u9_X_34 ) , .A1( u1_u9_X_35 ) , .ZN( u1_u9_u5_n145 ) );
  NOR2_X1 u1_u9_u5_U78 (.A2( u1_u9_X_34 ) , .ZN( u1_u9_u5_n146 ) , .A1( u1_u9_u5_n171 ) );
  NOR2_X1 u1_u9_u5_U79 (.A2( u1_u9_X_31 ) , .A1( u1_u9_X_32 ) , .ZN( u1_u9_u5_n103 ) );
  OAI22_X1 u1_u9_u5_U8 (.B2( u1_u9_u5_n149 ) , .B1( u1_u9_u5_n150 ) , .A2( u1_u9_u5_n151 ) , .A1( u1_u9_u5_n152 ) , .ZN( u1_u9_u5_n165 ) );
  NOR2_X1 u1_u9_u5_U80 (.A2( u1_u9_X_36 ) , .ZN( u1_u9_u5_n105 ) , .A1( u1_u9_u5_n180 ) );
  NOR2_X1 u1_u9_u5_U81 (.A2( u1_u9_X_33 ) , .ZN( u1_u9_u5_n108 ) , .A1( u1_u9_u5_n170 ) );
  NOR2_X1 u1_u9_u5_U82 (.A2( u1_u9_X_33 ) , .A1( u1_u9_X_36 ) , .ZN( u1_u9_u5_n107 ) );
  NOR2_X1 u1_u9_u5_U83 (.A2( u1_u9_X_31 ) , .ZN( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n181 ) );
  NAND2_X1 u1_u9_u5_U84 (.A2( u1_u9_X_34 ) , .A1( u1_u9_X_35 ) , .ZN( u1_u9_u5_n153 ) );
  NAND2_X1 u1_u9_u5_U85 (.A1( u1_u9_X_34 ) , .ZN( u1_u9_u5_n126 ) , .A2( u1_u9_u5_n171 ) );
  AND2_X1 u1_u9_u5_U86 (.A1( u1_u9_X_31 ) , .A2( u1_u9_X_32 ) , .ZN( u1_u9_u5_n106 ) );
  AND2_X1 u1_u9_u5_U87 (.A1( u1_u9_X_31 ) , .ZN( u1_u9_u5_n109 ) , .A2( u1_u9_u5_n181 ) );
  INV_X1 u1_u9_u5_U88 (.A( u1_u9_X_33 ) , .ZN( u1_u9_u5_n180 ) );
  INV_X1 u1_u9_u5_U89 (.A( u1_u9_X_35 ) , .ZN( u1_u9_u5_n171 ) );
  NOR3_X1 u1_u9_u5_U9 (.A2( u1_u9_u5_n147 ) , .A1( u1_u9_u5_n148 ) , .ZN( u1_u9_u5_n149 ) , .A3( u1_u9_u5_n194 ) );
  INV_X1 u1_u9_u5_U90 (.A( u1_u9_X_36 ) , .ZN( u1_u9_u5_n170 ) );
  INV_X1 u1_u9_u5_U91 (.A( u1_u9_X_32 ) , .ZN( u1_u9_u5_n181 ) );
  NAND4_X1 u1_u9_u5_U92 (.ZN( u1_out9_29 ) , .A4( u1_u9_u5_n129 ) , .A3( u1_u9_u5_n130 ) , .A2( u1_u9_u5_n168 ) , .A1( u1_u9_u5_n196 ) );
  AOI221_X1 u1_u9_u5_U93 (.A( u1_u9_u5_n128 ) , .ZN( u1_u9_u5_n129 ) , .C2( u1_u9_u5_n132 ) , .B2( u1_u9_u5_n159 ) , .B1( u1_u9_u5_n176 ) , .C1( u1_u9_u5_n184 ) );
  AOI222_X1 u1_u9_u5_U94 (.ZN( u1_u9_u5_n130 ) , .A2( u1_u9_u5_n146 ) , .B1( u1_u9_u5_n147 ) , .C2( u1_u9_u5_n175 ) , .B2( u1_u9_u5_n179 ) , .A1( u1_u9_u5_n188 ) , .C1( u1_u9_u5_n194 ) );
  NAND4_X1 u1_u9_u5_U95 (.ZN( u1_out9_19 ) , .A4( u1_u9_u5_n166 ) , .A3( u1_u9_u5_n167 ) , .A2( u1_u9_u5_n168 ) , .A1( u1_u9_u5_n169 ) );
  AOI22_X1 u1_u9_u5_U96 (.B2( u1_u9_u5_n145 ) , .A2( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n167 ) , .B1( u1_u9_u5_n182 ) , .A1( u1_u9_u5_n189 ) );
  NOR4_X1 u1_u9_u5_U97 (.A4( u1_u9_u5_n162 ) , .A3( u1_u9_u5_n163 ) , .A2( u1_u9_u5_n164 ) , .A1( u1_u9_u5_n165 ) , .ZN( u1_u9_u5_n166 ) );
  NAND4_X1 u1_u9_u5_U98 (.ZN( u1_out9_11 ) , .A4( u1_u9_u5_n143 ) , .A3( u1_u9_u5_n144 ) , .A2( u1_u9_u5_n169 ) , .A1( u1_u9_u5_n196 ) );
  AOI22_X1 u1_u9_u5_U99 (.A2( u1_u9_u5_n132 ) , .ZN( u1_u9_u5_n144 ) , .B2( u1_u9_u5_n145 ) , .B1( u1_u9_u5_n184 ) , .A1( u1_u9_u5_n194 ) );
  AOI22_X1 u1_u9_u6_U10 (.A2( u1_u9_u6_n151 ) , .B2( u1_u9_u6_n161 ) , .A1( u1_u9_u6_n167 ) , .B1( u1_u9_u6_n170 ) , .ZN( u1_u9_u6_n89 ) );
  AOI21_X1 u1_u9_u6_U11 (.B1( u1_u9_u6_n107 ) , .B2( u1_u9_u6_n132 ) , .A( u1_u9_u6_n158 ) , .ZN( u1_u9_u6_n88 ) );
  AOI21_X1 u1_u9_u6_U12 (.B2( u1_u9_u6_n147 ) , .B1( u1_u9_u6_n148 ) , .ZN( u1_u9_u6_n149 ) , .A( u1_u9_u6_n158 ) );
  AOI21_X1 u1_u9_u6_U13 (.ZN( u1_u9_u6_n106 ) , .A( u1_u9_u6_n142 ) , .B2( u1_u9_u6_n159 ) , .B1( u1_u9_u6_n164 ) );
  INV_X1 u1_u9_u6_U14 (.A( u1_u9_u6_n155 ) , .ZN( u1_u9_u6_n161 ) );
  INV_X1 u1_u9_u6_U15 (.A( u1_u9_u6_n128 ) , .ZN( u1_u9_u6_n164 ) );
  NAND2_X1 u1_u9_u6_U16 (.ZN( u1_u9_u6_n110 ) , .A1( u1_u9_u6_n122 ) , .A2( u1_u9_u6_n129 ) );
  NAND2_X1 u1_u9_u6_U17 (.ZN( u1_u9_u6_n124 ) , .A2( u1_u9_u6_n146 ) , .A1( u1_u9_u6_n148 ) );
  INV_X1 u1_u9_u6_U18 (.A( u1_u9_u6_n132 ) , .ZN( u1_u9_u6_n171 ) );
  AND2_X1 u1_u9_u6_U19 (.A1( u1_u9_u6_n100 ) , .ZN( u1_u9_u6_n130 ) , .A2( u1_u9_u6_n147 ) );
  INV_X1 u1_u9_u6_U20 (.A( u1_u9_u6_n127 ) , .ZN( u1_u9_u6_n173 ) );
  INV_X1 u1_u9_u6_U21 (.A( u1_u9_u6_n121 ) , .ZN( u1_u9_u6_n167 ) );
  INV_X1 u1_u9_u6_U22 (.A( u1_u9_u6_n100 ) , .ZN( u1_u9_u6_n169 ) );
  INV_X1 u1_u9_u6_U23 (.A( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n170 ) );
  INV_X1 u1_u9_u6_U24 (.A( u1_u9_u6_n113 ) , .ZN( u1_u9_u6_n168 ) );
  AND2_X1 u1_u9_u6_U25 (.A1( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n119 ) , .ZN( u1_u9_u6_n133 ) );
  AND2_X1 u1_u9_u6_U26 (.A2( u1_u9_u6_n121 ) , .A1( u1_u9_u6_n122 ) , .ZN( u1_u9_u6_n131 ) );
  AND3_X1 u1_u9_u6_U27 (.ZN( u1_u9_u6_n120 ) , .A2( u1_u9_u6_n127 ) , .A1( u1_u9_u6_n132 ) , .A3( u1_u9_u6_n145 ) );
  INV_X1 u1_u9_u6_U28 (.A( u1_u9_u6_n146 ) , .ZN( u1_u9_u6_n163 ) );
  AOI222_X1 u1_u9_u6_U29 (.ZN( u1_u9_u6_n114 ) , .A1( u1_u9_u6_n118 ) , .A2( u1_u9_u6_n126 ) , .B2( u1_u9_u6_n151 ) , .C2( u1_u9_u6_n159 ) , .C1( u1_u9_u6_n168 ) , .B1( u1_u9_u6_n169 ) );
  INV_X1 u1_u9_u6_U3 (.A( u1_u9_u6_n110 ) , .ZN( u1_u9_u6_n166 ) );
  NOR2_X1 u1_u9_u6_U30 (.A1( u1_u9_u6_n162 ) , .A2( u1_u9_u6_n165 ) , .ZN( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U31 (.A1( u1_u9_u6_n144 ) , .ZN( u1_u9_u6_n151 ) , .A2( u1_u9_u6_n158 ) );
  NAND2_X1 u1_u9_u6_U32 (.ZN( u1_u9_u6_n132 ) , .A1( u1_u9_u6_n91 ) , .A2( u1_u9_u6_n97 ) );
  AOI22_X1 u1_u9_u6_U33 (.B2( u1_u9_u6_n110 ) , .B1( u1_u9_u6_n111 ) , .A1( u1_u9_u6_n112 ) , .ZN( u1_u9_u6_n115 ) , .A2( u1_u9_u6_n161 ) );
  NAND4_X1 u1_u9_u6_U34 (.A3( u1_u9_u6_n109 ) , .ZN( u1_u9_u6_n112 ) , .A4( u1_u9_u6_n132 ) , .A2( u1_u9_u6_n147 ) , .A1( u1_u9_u6_n166 ) );
  NOR2_X1 u1_u9_u6_U35 (.ZN( u1_u9_u6_n109 ) , .A1( u1_u9_u6_n170 ) , .A2( u1_u9_u6_n173 ) );
  NOR2_X1 u1_u9_u6_U36 (.A2( u1_u9_u6_n126 ) , .ZN( u1_u9_u6_n155 ) , .A1( u1_u9_u6_n160 ) );
  NAND2_X1 u1_u9_u6_U37 (.ZN( u1_u9_u6_n146 ) , .A2( u1_u9_u6_n94 ) , .A1( u1_u9_u6_n99 ) );
  AOI21_X1 u1_u9_u6_U38 (.A( u1_u9_u6_n144 ) , .B2( u1_u9_u6_n145 ) , .B1( u1_u9_u6_n146 ) , .ZN( u1_u9_u6_n150 ) );
  AOI211_X1 u1_u9_u6_U39 (.B( u1_u9_u6_n134 ) , .A( u1_u9_u6_n135 ) , .C1( u1_u9_u6_n136 ) , .ZN( u1_u9_u6_n137 ) , .C2( u1_u9_u6_n151 ) );
  INV_X1 u1_u9_u6_U4 (.A( u1_u9_u6_n142 ) , .ZN( u1_u9_u6_n174 ) );
  NAND4_X1 u1_u9_u6_U40 (.A4( u1_u9_u6_n127 ) , .A3( u1_u9_u6_n128 ) , .A2( u1_u9_u6_n129 ) , .A1( u1_u9_u6_n130 ) , .ZN( u1_u9_u6_n136 ) );
  AOI21_X1 u1_u9_u6_U41 (.B2( u1_u9_u6_n132 ) , .B1( u1_u9_u6_n133 ) , .ZN( u1_u9_u6_n134 ) , .A( u1_u9_u6_n158 ) );
  AOI21_X1 u1_u9_u6_U42 (.B1( u1_u9_u6_n131 ) , .ZN( u1_u9_u6_n135 ) , .A( u1_u9_u6_n144 ) , .B2( u1_u9_u6_n146 ) );
  INV_X1 u1_u9_u6_U43 (.A( u1_u9_u6_n111 ) , .ZN( u1_u9_u6_n158 ) );
  NAND2_X1 u1_u9_u6_U44 (.ZN( u1_u9_u6_n127 ) , .A1( u1_u9_u6_n91 ) , .A2( u1_u9_u6_n92 ) );
  NAND2_X1 u1_u9_u6_U45 (.ZN( u1_u9_u6_n129 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n96 ) );
  INV_X1 u1_u9_u6_U46 (.A( u1_u9_u6_n144 ) , .ZN( u1_u9_u6_n159 ) );
  NAND2_X1 u1_u9_u6_U47 (.ZN( u1_u9_u6_n145 ) , .A2( u1_u9_u6_n97 ) , .A1( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U48 (.ZN( u1_u9_u6_n148 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n94 ) );
  NAND2_X1 u1_u9_u6_U49 (.ZN( u1_u9_u6_n108 ) , .A2( u1_u9_u6_n139 ) , .A1( u1_u9_u6_n144 ) );
  NAND2_X1 u1_u9_u6_U5 (.A2( u1_u9_u6_n143 ) , .ZN( u1_u9_u6_n152 ) , .A1( u1_u9_u6_n166 ) );
  NAND2_X1 u1_u9_u6_U50 (.ZN( u1_u9_u6_n121 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n97 ) );
  NAND2_X1 u1_u9_u6_U51 (.ZN( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n95 ) );
  AND2_X1 u1_u9_u6_U52 (.ZN( u1_u9_u6_n118 ) , .A2( u1_u9_u6_n91 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U53 (.ZN( u1_u9_u6_n147 ) , .A2( u1_u9_u6_n98 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U54 (.ZN( u1_u9_u6_n128 ) , .A1( u1_u9_u6_n94 ) , .A2( u1_u9_u6_n96 ) );
  NAND2_X1 u1_u9_u6_U55 (.ZN( u1_u9_u6_n119 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U56 (.ZN( u1_u9_u6_n123 ) , .A2( u1_u9_u6_n91 ) , .A1( u1_u9_u6_n96 ) );
  NAND2_X1 u1_u9_u6_U57 (.ZN( u1_u9_u6_n100 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U58 (.ZN( u1_u9_u6_n122 ) , .A1( u1_u9_u6_n94 ) , .A2( u1_u9_u6_n97 ) );
  INV_X1 u1_u9_u6_U59 (.A( u1_u9_u6_n139 ) , .ZN( u1_u9_u6_n160 ) );
  AOI22_X1 u1_u9_u6_U6 (.B2( u1_u9_u6_n101 ) , .A1( u1_u9_u6_n102 ) , .ZN( u1_u9_u6_n103 ) , .B1( u1_u9_u6_n160 ) , .A2( u1_u9_u6_n161 ) );
  NAND2_X1 u1_u9_u6_U60 (.ZN( u1_u9_u6_n113 ) , .A1( u1_u9_u6_n96 ) , .A2( u1_u9_u6_n98 ) );
  NOR2_X1 u1_u9_u6_U61 (.A2( u1_u9_X_40 ) , .A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n126 ) );
  NOR2_X1 u1_u9_u6_U62 (.A2( u1_u9_X_39 ) , .A1( u1_u9_X_42 ) , .ZN( u1_u9_u6_n92 ) );
  NOR2_X1 u1_u9_u6_U63 (.A2( u1_u9_X_39 ) , .A1( u1_u9_u6_n156 ) , .ZN( u1_u9_u6_n97 ) );
  NOR2_X1 u1_u9_u6_U64 (.A2( u1_u9_X_38 ) , .A1( u1_u9_u6_n165 ) , .ZN( u1_u9_u6_n95 ) );
  NOR2_X1 u1_u9_u6_U65 (.A2( u1_u9_X_41 ) , .ZN( u1_u9_u6_n111 ) , .A1( u1_u9_u6_n157 ) );
  NOR2_X1 u1_u9_u6_U66 (.A2( u1_u9_X_37 ) , .A1( u1_u9_u6_n162 ) , .ZN( u1_u9_u6_n94 ) );
  NOR2_X1 u1_u9_u6_U67 (.A2( u1_u9_X_37 ) , .A1( u1_u9_X_38 ) , .ZN( u1_u9_u6_n91 ) );
  NAND2_X1 u1_u9_u6_U68 (.A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n144 ) , .A2( u1_u9_u6_n157 ) );
  NAND2_X1 u1_u9_u6_U69 (.A2( u1_u9_X_40 ) , .A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n139 ) );
  NOR2_X1 u1_u9_u6_U7 (.A1( u1_u9_u6_n118 ) , .ZN( u1_u9_u6_n143 ) , .A2( u1_u9_u6_n168 ) );
  AND2_X1 u1_u9_u6_U70 (.A1( u1_u9_X_39 ) , .A2( u1_u9_u6_n156 ) , .ZN( u1_u9_u6_n96 ) );
  AND2_X1 u1_u9_u6_U71 (.A1( u1_u9_X_39 ) , .A2( u1_u9_X_42 ) , .ZN( u1_u9_u6_n99 ) );
  INV_X1 u1_u9_u6_U72 (.A( u1_u9_X_40 ) , .ZN( u1_u9_u6_n157 ) );
  INV_X1 u1_u9_u6_U73 (.A( u1_u9_X_37 ) , .ZN( u1_u9_u6_n165 ) );
  INV_X1 u1_u9_u6_U74 (.A( u1_u9_X_38 ) , .ZN( u1_u9_u6_n162 ) );
  INV_X1 u1_u9_u6_U75 (.A( u1_u9_X_42 ) , .ZN( u1_u9_u6_n156 ) );
  NAND4_X1 u1_u9_u6_U76 (.ZN( u1_out9_12 ) , .A4( u1_u9_u6_n114 ) , .A3( u1_u9_u6_n115 ) , .A2( u1_u9_u6_n116 ) , .A1( u1_u9_u6_n117 ) );
  OAI22_X1 u1_u9_u6_U77 (.B2( u1_u9_u6_n111 ) , .ZN( u1_u9_u6_n116 ) , .B1( u1_u9_u6_n126 ) , .A2( u1_u9_u6_n164 ) , .A1( u1_u9_u6_n167 ) );
  OAI21_X1 u1_u9_u6_U78 (.A( u1_u9_u6_n108 ) , .ZN( u1_u9_u6_n117 ) , .B2( u1_u9_u6_n141 ) , .B1( u1_u9_u6_n163 ) );
  NAND4_X1 u1_u9_u6_U79 (.ZN( u1_out9_32 ) , .A4( u1_u9_u6_n103 ) , .A3( u1_u9_u6_n104 ) , .A2( u1_u9_u6_n105 ) , .A1( u1_u9_u6_n106 ) );
  OAI21_X1 u1_u9_u6_U8 (.A( u1_u9_u6_n159 ) , .B1( u1_u9_u6_n169 ) , .B2( u1_u9_u6_n173 ) , .ZN( u1_u9_u6_n90 ) );
  AOI22_X1 u1_u9_u6_U80 (.ZN( u1_u9_u6_n105 ) , .A2( u1_u9_u6_n108 ) , .A1( u1_u9_u6_n118 ) , .B2( u1_u9_u6_n126 ) , .B1( u1_u9_u6_n171 ) );
  AOI22_X1 u1_u9_u6_U81 (.ZN( u1_u9_u6_n104 ) , .A1( u1_u9_u6_n111 ) , .B1( u1_u9_u6_n124 ) , .B2( u1_u9_u6_n151 ) , .A2( u1_u9_u6_n93 ) );
  OAI211_X1 u1_u9_u6_U82 (.ZN( u1_out9_7 ) , .B( u1_u9_u6_n153 ) , .C2( u1_u9_u6_n154 ) , .C1( u1_u9_u6_n155 ) , .A( u1_u9_u6_n174 ) );
  NOR3_X1 u1_u9_u6_U83 (.A1( u1_u9_u6_n141 ) , .ZN( u1_u9_u6_n154 ) , .A3( u1_u9_u6_n164 ) , .A2( u1_u9_u6_n171 ) );
  AOI211_X1 u1_u9_u6_U84 (.B( u1_u9_u6_n149 ) , .A( u1_u9_u6_n150 ) , .C2( u1_u9_u6_n151 ) , .C1( u1_u9_u6_n152 ) , .ZN( u1_u9_u6_n153 ) );
  OAI211_X1 u1_u9_u6_U85 (.ZN( u1_out9_22 ) , .B( u1_u9_u6_n137 ) , .A( u1_u9_u6_n138 ) , .C2( u1_u9_u6_n139 ) , .C1( u1_u9_u6_n140 ) );
  AOI22_X1 u1_u9_u6_U86 (.B1( u1_u9_u6_n124 ) , .A2( u1_u9_u6_n125 ) , .A1( u1_u9_u6_n126 ) , .ZN( u1_u9_u6_n138 ) , .B2( u1_u9_u6_n161 ) );
  AND4_X1 u1_u9_u6_U87 (.A3( u1_u9_u6_n119 ) , .A1( u1_u9_u6_n120 ) , .A4( u1_u9_u6_n129 ) , .ZN( u1_u9_u6_n140 ) , .A2( u1_u9_u6_n143 ) );
  NAND3_X1 u1_u9_u6_U88 (.A2( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n125 ) , .A1( u1_u9_u6_n130 ) , .A3( u1_u9_u6_n131 ) );
  NAND3_X1 u1_u9_u6_U89 (.A3( u1_u9_u6_n133 ) , .ZN( u1_u9_u6_n141 ) , .A1( u1_u9_u6_n145 ) , .A2( u1_u9_u6_n148 ) );
  INV_X1 u1_u9_u6_U9 (.ZN( u1_u9_u6_n172 ) , .A( u1_u9_u6_n88 ) );
  NAND3_X1 u1_u9_u6_U90 (.ZN( u1_u9_u6_n101 ) , .A3( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n121 ) , .A1( u1_u9_u6_n127 ) );
  NAND3_X1 u1_u9_u6_U91 (.ZN( u1_u9_u6_n102 ) , .A3( u1_u9_u6_n130 ) , .A2( u1_u9_u6_n145 ) , .A1( u1_u9_u6_n166 ) );
  NAND3_X1 u1_u9_u6_U92 (.A3( u1_u9_u6_n113 ) , .A1( u1_u9_u6_n119 ) , .A2( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n93 ) );
  NAND3_X1 u1_u9_u6_U93 (.ZN( u1_u9_u6_n142 ) , .A2( u1_u9_u6_n172 ) , .A3( u1_u9_u6_n89 ) , .A1( u1_u9_u6_n90 ) );
  AND3_X1 u1_u9_u7_U10 (.A3( u1_u9_u7_n110 ) , .A2( u1_u9_u7_n127 ) , .A1( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U11 (.A( u1_u9_u7_n161 ) , .B1( u1_u9_u7_n168 ) , .B2( u1_u9_u7_n173 ) , .ZN( u1_u9_u7_n91 ) );
  AOI211_X1 u1_u9_u7_U12 (.A( u1_u9_u7_n117 ) , .ZN( u1_u9_u7_n118 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n177 ) , .B( u1_u9_u7_n180 ) );
  OAI22_X1 u1_u9_u7_U13 (.B1( u1_u9_u7_n115 ) , .ZN( u1_u9_u7_n117 ) , .A2( u1_u9_u7_n133 ) , .A1( u1_u9_u7_n137 ) , .B2( u1_u9_u7_n162 ) );
  INV_X1 u1_u9_u7_U14 (.A( u1_u9_u7_n116 ) , .ZN( u1_u9_u7_n180 ) );
  NOR3_X1 u1_u9_u7_U15 (.ZN( u1_u9_u7_n115 ) , .A3( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n168 ) , .A1( u1_u9_u7_n169 ) );
  OAI211_X1 u1_u9_u7_U16 (.B( u1_u9_u7_n122 ) , .A( u1_u9_u7_n123 ) , .C2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n154 ) , .C1( u1_u9_u7_n162 ) );
  AOI222_X1 u1_u9_u7_U17 (.ZN( u1_u9_u7_n122 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n161 ) , .A2( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n170 ) , .A1( u1_u9_u7_n176 ) );
  INV_X1 u1_u9_u7_U18 (.A( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n176 ) );
  NOR3_X1 u1_u9_u7_U19 (.A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n135 ) , .ZN( u1_u9_u7_n136 ) , .A3( u1_u9_u7_n171 ) );
  NOR2_X1 u1_u9_u7_U20 (.A1( u1_u9_u7_n130 ) , .A2( u1_u9_u7_n134 ) , .ZN( u1_u9_u7_n153 ) );
  INV_X1 u1_u9_u7_U21 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n165 ) );
  NOR2_X1 u1_u9_u7_U22 (.ZN( u1_u9_u7_n111 ) , .A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n169 ) );
  AOI21_X1 u1_u9_u7_U23 (.ZN( u1_u9_u7_n104 ) , .B2( u1_u9_u7_n112 ) , .B1( u1_u9_u7_n127 ) , .A( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U24 (.ZN( u1_u9_u7_n106 ) , .B1( u1_u9_u7_n133 ) , .B2( u1_u9_u7_n146 ) , .A( u1_u9_u7_n162 ) );
  AOI21_X1 u1_u9_u7_U25 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n107 ) , .B2( u1_u9_u7_n128 ) , .B1( u1_u9_u7_n175 ) );
  INV_X1 u1_u9_u7_U26 (.A( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n171 ) );
  INV_X1 u1_u9_u7_U27 (.A( u1_u9_u7_n131 ) , .ZN( u1_u9_u7_n177 ) );
  INV_X1 u1_u9_u7_U28 (.A( u1_u9_u7_n110 ) , .ZN( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U29 (.A1( u1_u9_u7_n129 ) , .A2( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n149 ) );
  OAI21_X1 u1_u9_u7_U3 (.ZN( u1_u9_u7_n159 ) , .A( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n171 ) , .B1( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U30 (.A1( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n130 ) );
  INV_X1 u1_u9_u7_U31 (.A( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n173 ) );
  INV_X1 u1_u9_u7_U32 (.A( u1_u9_u7_n128 ) , .ZN( u1_u9_u7_n168 ) );
  INV_X1 u1_u9_u7_U33 (.A( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n169 ) );
  INV_X1 u1_u9_u7_U34 (.A( u1_u9_u7_n127 ) , .ZN( u1_u9_u7_n179 ) );
  NOR2_X1 u1_u9_u7_U35 (.ZN( u1_u9_u7_n101 ) , .A2( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n156 ) );
  AOI211_X1 u1_u9_u7_U36 (.B( u1_u9_u7_n154 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n156 ) , .ZN( u1_u9_u7_n157 ) , .C2( u1_u9_u7_n172 ) );
  INV_X1 u1_u9_u7_U37 (.A( u1_u9_u7_n153 ) , .ZN( u1_u9_u7_n172 ) );
  AOI211_X1 u1_u9_u7_U38 (.B( u1_u9_u7_n139 ) , .A( u1_u9_u7_n140 ) , .C2( u1_u9_u7_n141 ) , .ZN( u1_u9_u7_n142 ) , .C1( u1_u9_u7_n156 ) );
  NAND4_X1 u1_u9_u7_U39 (.A3( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n141 ) , .A4( u1_u9_u7_n147 ) );
  INV_X1 u1_u9_u7_U4 (.A( u1_u9_u7_n111 ) , .ZN( u1_u9_u7_n170 ) );
  AOI21_X1 u1_u9_u7_U40 (.A( u1_u9_u7_n137 ) , .B1( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n139 ) , .B2( u1_u9_u7_n146 ) );
  OAI22_X1 u1_u9_u7_U41 (.B1( u1_u9_u7_n136 ) , .ZN( u1_u9_u7_n140 ) , .A1( u1_u9_u7_n153 ) , .B2( u1_u9_u7_n162 ) , .A2( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U42 (.ZN( u1_u9_u7_n123 ) , .B1( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n177 ) , .A( u1_u9_u7_n97 ) );
  AOI21_X1 u1_u9_u7_U43 (.B2( u1_u9_u7_n113 ) , .B1( u1_u9_u7_n124 ) , .A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n97 ) );
  INV_X1 u1_u9_u7_U44 (.A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U45 (.A( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n162 ) );
  AOI22_X1 u1_u9_u7_U46 (.A2( u1_u9_u7_n114 ) , .ZN( u1_u9_u7_n119 ) , .B1( u1_u9_u7_n130 ) , .A1( u1_u9_u7_n156 ) , .B2( u1_u9_u7_n165 ) );
  NAND2_X1 u1_u9_u7_U47 (.A2( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n114 ) , .A1( u1_u9_u7_n175 ) );
  AND2_X1 u1_u9_u7_U48 (.ZN( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n98 ) , .A1( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U49 (.ZN( u1_u9_u7_n137 ) , .A1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U5 (.A( u1_u9_u7_n149 ) , .ZN( u1_u9_u7_n175 ) );
  AOI21_X1 u1_u9_u7_U50 (.ZN( u1_u9_u7_n105 ) , .B2( u1_u9_u7_n110 ) , .A( u1_u9_u7_n125 ) , .B1( u1_u9_u7_n147 ) );
  NAND2_X1 u1_u9_u7_U51 (.ZN( u1_u9_u7_n146 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U52 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U53 (.A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n99 ) );
  OR2_X1 u1_u9_u7_U54 (.ZN( u1_u9_u7_n126 ) , .A2( u1_u9_u7_n152 ) , .A1( u1_u9_u7_n156 ) );
  NAND2_X1 u1_u9_u7_U55 (.A2( u1_u9_u7_n102 ) , .A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n133 ) );
  NAND2_X1 u1_u9_u7_U56 (.ZN( u1_u9_u7_n112 ) , .A2( u1_u9_u7_n96 ) , .A1( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U57 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U58 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U59 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n124 ) , .A1( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U6 (.A( u1_u9_u7_n154 ) , .ZN( u1_u9_u7_n178 ) );
  NAND2_X1 u1_u9_u7_U60 (.ZN( u1_u9_u7_n110 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U61 (.A( u1_u9_u7_n150 ) , .ZN( u1_u9_u7_n164 ) );
  AND2_X1 u1_u9_u7_U62 (.ZN( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U63 (.A1( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n129 ) );
  NAND2_X1 u1_u9_u7_U64 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n131 ) , .A1( u1_u9_u7_n95 ) );
  NAND2_X1 u1_u9_u7_U65 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n138 ) , .A2( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U66 (.ZN( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n96 ) );
  NAND2_X1 u1_u9_u7_U67 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n148 ) , .A2( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U68 (.A2( u1_u9_X_47 ) , .ZN( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n163 ) );
  NOR2_X1 u1_u9_u7_U69 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n103 ) );
  AOI211_X1 u1_u9_u7_U7 (.ZN( u1_u9_u7_n116 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n161 ) , .C2( u1_u9_u7_n171 ) , .B( u1_u9_u7_n94 ) );
  NOR2_X1 u1_u9_u7_U70 (.A2( u1_u9_X_48 ) , .A1( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U71 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U72 (.A2( u1_u9_X_44 ) , .A1( u1_u9_u7_n167 ) , .ZN( u1_u9_u7_n98 ) );
  NOR2_X1 u1_u9_u7_U73 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n152 ) );
  AND2_X1 u1_u9_u7_U74 (.A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n156 ) , .A2( u1_u9_u7_n163 ) );
  NAND2_X1 u1_u9_u7_U75 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n125 ) );
  AND2_X1 u1_u9_u7_U76 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n102 ) );
  AND2_X1 u1_u9_u7_U77 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n96 ) );
  AND2_X1 u1_u9_u7_U78 (.A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n167 ) );
  AND2_X1 u1_u9_u7_U79 (.A1( u1_u9_X_48 ) , .A2( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n93 ) );
  OAI222_X1 u1_u9_u7_U8 (.C2( u1_u9_u7_n101 ) , .B2( u1_u9_u7_n111 ) , .A1( u1_u9_u7_n113 ) , .C1( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n162 ) , .B1( u1_u9_u7_n164 ) , .ZN( u1_u9_u7_n94 ) );
  INV_X1 u1_u9_u7_U80 (.A( u1_u9_X_46 ) , .ZN( u1_u9_u7_n163 ) );
  INV_X1 u1_u9_u7_U81 (.A( u1_u9_X_43 ) , .ZN( u1_u9_u7_n167 ) );
  INV_X1 u1_u9_u7_U82 (.A( u1_u9_X_45 ) , .ZN( u1_u9_u7_n166 ) );
  NAND4_X1 u1_u9_u7_U83 (.ZN( u1_out9_5 ) , .A4( u1_u9_u7_n108 ) , .A3( u1_u9_u7_n109 ) , .A1( u1_u9_u7_n116 ) , .A2( u1_u9_u7_n123 ) );
  AOI22_X1 u1_u9_u7_U84 (.ZN( u1_u9_u7_n109 ) , .A2( u1_u9_u7_n126 ) , .B2( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n156 ) , .A1( u1_u9_u7_n171 ) );
  NOR4_X1 u1_u9_u7_U85 (.A4( u1_u9_u7_n104 ) , .A3( u1_u9_u7_n105 ) , .A2( u1_u9_u7_n106 ) , .A1( u1_u9_u7_n107 ) , .ZN( u1_u9_u7_n108 ) );
  NAND4_X1 u1_u9_u7_U86 (.ZN( u1_out9_27 ) , .A4( u1_u9_u7_n118 ) , .A3( u1_u9_u7_n119 ) , .A2( u1_u9_u7_n120 ) , .A1( u1_u9_u7_n121 ) );
  OAI21_X1 u1_u9_u7_U87 (.ZN( u1_u9_u7_n121 ) , .B2( u1_u9_u7_n145 ) , .A( u1_u9_u7_n150 ) , .B1( u1_u9_u7_n174 ) );
  OAI21_X1 u1_u9_u7_U88 (.ZN( u1_u9_u7_n120 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n170 ) , .B1( u1_u9_u7_n179 ) );
  NAND4_X1 u1_u9_u7_U89 (.ZN( u1_out9_21 ) , .A4( u1_u9_u7_n157 ) , .A3( u1_u9_u7_n158 ) , .A2( u1_u9_u7_n159 ) , .A1( u1_u9_u7_n160 ) );
  OAI221_X1 u1_u9_u7_U9 (.C1( u1_u9_u7_n101 ) , .C2( u1_u9_u7_n147 ) , .ZN( u1_u9_u7_n155 ) , .B2( u1_u9_u7_n162 ) , .A( u1_u9_u7_n91 ) , .B1( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U90 (.B1( u1_u9_u7_n145 ) , .ZN( u1_u9_u7_n160 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n177 ) );
  AOI22_X1 u1_u9_u7_U91 (.B2( u1_u9_u7_n149 ) , .B1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n151 ) , .A1( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n158 ) );
  NAND4_X1 u1_u9_u7_U92 (.ZN( u1_out9_15 ) , .A4( u1_u9_u7_n142 ) , .A3( u1_u9_u7_n143 ) , .A2( u1_u9_u7_n144 ) , .A1( u1_u9_u7_n178 ) );
  OR2_X1 u1_u9_u7_U93 (.A2( u1_u9_u7_n125 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n144 ) );
  AOI22_X1 u1_u9_u7_U94 (.A2( u1_u9_u7_n126 ) , .ZN( u1_u9_u7_n143 ) , .B2( u1_u9_u7_n165 ) , .B1( u1_u9_u7_n173 ) , .A1( u1_u9_u7_n174 ) );
  NAND3_X1 u1_u9_u7_U95 (.A3( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n151 ) );
  NAND3_X1 u1_u9_u7_U96 (.A3( u1_u9_u7_n131 ) , .A2( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n135 ) );
  INV_X1 u1_uk_U105 (.ZN( u1_K11_5 ) , .A( u1_uk_n496 ) );
  INV_X1 u1_uk_U112 (.ZN( u1_K13_5 ) , .A( u1_uk_n948 ) );
  INV_X1 u1_uk_U1127 (.ZN( u1_K1_41 ) , .A( u1_uk_n1015 ) );
  INV_X1 u1_uk_U1131 (.ZN( u1_K11_12 ) , .A( u1_uk_n379 ) );
  INV_X1 u1_uk_U1145 (.ZN( u1_K9_20 ) , .A( u1_uk_n1156 ) );
  INV_X1 u1_uk_U1149 (.ZN( u1_K7_13 ) , .A( u1_uk_n1106 ) );
  INV_X1 u1_uk_U1163 (.ZN( u1_K13_12 ) , .A( u1_uk_n676 ) );
  INV_X1 u1_uk_U1166 (.ZN( u1_K15_43 ) , .A( u1_uk_n974 ) );
  INV_X1 u1_uk_U1168 (.ZN( u1_K13_2 ) , .A( u1_uk_n702 ) );
  INV_X1 u1_uk_U1170 (.ZN( u1_K9_2 ) , .A( u1_uk_n1160 ) );
  INV_X1 u1_uk_U1171 (.ZN( u1_K4_2 ) , .A( u1_uk_n1061 ) );
  INV_X1 u1_uk_U1172 (.ZN( u1_K13_6 ) , .A( u1_uk_n949 ) );
  INV_X1 u1_uk_U141 (.ZN( u1_K13_15 ) , .A( u1_uk_n678 ) );
  INV_X1 u1_uk_U147 (.ZN( u1_K13_19 ) , .A( u1_uk_n685 ) );
  INV_X1 u1_uk_U163 (.ZN( u1_K9_19 ) , .A( u1_uk_n1154 ) );
  INV_X1 u1_uk_U169 (.ZN( u1_K2_19 ) , .A( u1_uk_n1025 ) );
  INV_X1 u1_uk_U190 (.ZN( u1_K11_14 ) , .A( u1_uk_n382 ) );
  INV_X1 u1_uk_U215 (.ZN( u1_K15_30 ) , .A( u1_uk_n970 ) );
  INV_X1 u1_uk_U226 (.ZN( u1_K11_31 ) , .A( u1_uk_n437 ) );
  INV_X1 u1_uk_U276 (.ZN( u1_K9_48 ) , .A( u1_uk_n1170 ) );
  INV_X1 u1_uk_U299 (.ZN( u1_K15_8 ) , .A( u1_uk_n976 ) );
  INV_X1 u1_uk_U303 (.ZN( u1_K7_8 ) , .A( u1_uk_n1126 ) );
  INV_X1 u1_uk_U306 (.ZN( u1_K4_8 ) , .A( u1_uk_n1070 ) );
  INV_X1 u1_uk_U315 (.ZN( u1_K9_26 ) , .A( u1_uk_n1158 ) );
  INV_X1 u1_uk_U319 (.ZN( u1_K15_26 ) , .A( u1_uk_n969 ) );
  INV_X1 u1_uk_U369 (.ZN( u1_K7_46 ) , .A( u1_uk_n1124 ) );
  INV_X1 u1_uk_U441 (.ZN( u1_K10_37 ) , .A( u1_uk_n366 ) );
  INV_X1 u1_uk_U463 (.ZN( u1_K10_33 ) , .A( u1_uk_n349 ) );
  INV_X1 u1_uk_U495 (.ZN( u1_K16_29 ) , .A( u1_uk_n985 ) );
  INV_X1 u1_uk_U536 (.ZN( u1_K11_17 ) , .A( u1_uk_n385 ) );
  INV_X1 u1_uk_U538 (.ZN( u1_K7_12 ) , .A( u1_uk_n1105 ) );
  INV_X1 u1_uk_U568 (.ZN( u1_K11_36 ) , .A( u1_uk_n454 ) );
  INV_X1 u1_uk_U572 (.ZN( u1_K15_38 ) , .A( u1_uk_n973 ) );
  INV_X1 u1_uk_U574 (.ZN( u1_K10_38 ) , .A( u1_uk_n369 ) );
  INV_X1 u1_uk_U592 (.ZN( u1_K4_10 ) , .A( u1_uk_n1050 ) );
  INV_X1 u1_uk_U605 (.ZN( u1_K9_22 ) , .A( u1_uk_n1157 ) );
  INV_X1 u1_uk_U608 (.ZN( u1_K5_22 ) , .A( u1_uk_n1074 ) );
  INV_X1 u1_uk_U622 (.ZN( u1_K10_35 ) , .A( u1_uk_n353 ) );
  INV_X1 u1_uk_U624 (.ZN( u1_K9_35 ) , .A( u1_uk_n1163 ) );
  INV_X1 u1_uk_U642 (.ZN( u1_K13_11 ) , .A( u1_uk_n672 ) );
  INV_X1 u1_uk_U67 (.ZN( u1_K16_34 ) , .A( u1_uk_n988 ) );
  INV_X1 u1_uk_U69 (.ZN( u1_K11_34 ) , .A( u1_uk_n443 ) );
  INV_X1 u1_uk_U707 (.ZN( u1_K4_3 ) , .A( u1_uk_n1065 ) );
  INV_X1 u1_uk_U709 (.ZN( u1_K13_7 ) , .A( u1_uk_n950 ) );
  INV_X1 u1_uk_U742 (.ZN( u1_K9_42 ) , .A( u1_uk_n1167 ) );
  INV_X1 u1_uk_U744 (.ZN( u1_K7_42 ) , .A( u1_uk_n1123 ) );
  INV_X1 u1_uk_U781 (.ZN( u1_K13_13 ) , .A( u1_uk_n677 ) );
  INV_X1 u1_uk_U800 (.ZN( u1_K9_27 ) , .A( u1_uk_n1159 ) );
  INV_X1 u1_uk_U806 (.ZN( u1_K9_1 ) , .A( u1_uk_n1155 ) );
  INV_X1 u1_uk_U839 (.ZN( u1_K5_20 ) , .A( u1_uk_n1073 ) );
  INV_X1 u1_uk_U851 (.ZN( u1_K7_6 ) , .A( u1_uk_n1125 ) );
  INV_X1 u1_uk_U97 (.ZN( u1_K9_41 ) , .A( u1_uk_n1166 ) );
  INV_X1 u1_uk_U99 (.ZN( u1_K2_41 ) , .A( u1_uk_n1031 ) );
  XOR2_X1 u2_u10_U41 (.B( u2_K11_17 ) , .A( u2_R9_12 ) , .Z( u2_u10_X_17 ) );
  XOR2_X1 u2_u10_U44 (.B( u2_K11_14 ) , .A( u2_R9_9 ) , .Z( u2_u10_X_14 ) );
  XOR2_X1 u2_u10_U45 (.B( u2_K11_13 ) , .A( u2_R9_8 ) , .Z( u2_u10_X_13 ) );
  XOR2_X1 u2_u10_U46 (.B( u2_K11_12 ) , .A( u2_R9_9 ) , .Z( u2_u10_X_12 ) );
  XOR2_X1 u2_u10_U47 (.B( u2_K11_11 ) , .A( u2_R9_8 ) , .Z( u2_u10_X_11 ) );
  AOI21_X1 u2_u10_u1_U10 (.B2( u2_u10_u1_n155 ) , .B1( u2_u10_u1_n156 ) , .ZN( u2_u10_u1_n157 ) , .A( u2_u10_u1_n174 ) );
  NAND3_X1 u2_u10_u1_U100 (.ZN( u2_u10_u1_n113 ) , .A1( u2_u10_u1_n120 ) , .A3( u2_u10_u1_n133 ) , .A2( u2_u10_u1_n155 ) );
  NAND2_X1 u2_u10_u1_U11 (.ZN( u2_u10_u1_n140 ) , .A2( u2_u10_u1_n150 ) , .A1( u2_u10_u1_n155 ) );
  NAND2_X1 u2_u10_u1_U12 (.A1( u2_u10_u1_n131 ) , .ZN( u2_u10_u1_n147 ) , .A2( u2_u10_u1_n153 ) );
  AOI22_X1 u2_u10_u1_U13 (.B2( u2_u10_u1_n136 ) , .A2( u2_u10_u1_n137 ) , .ZN( u2_u10_u1_n143 ) , .A1( u2_u10_u1_n171 ) , .B1( u2_u10_u1_n173 ) );
  INV_X1 u2_u10_u1_U14 (.A( u2_u10_u1_n147 ) , .ZN( u2_u10_u1_n181 ) );
  INV_X1 u2_u10_u1_U15 (.A( u2_u10_u1_n139 ) , .ZN( u2_u10_u1_n174 ) );
  OR4_X1 u2_u10_u1_U16 (.A4( u2_u10_u1_n106 ) , .A3( u2_u10_u1_n107 ) , .ZN( u2_u10_u1_n108 ) , .A1( u2_u10_u1_n117 ) , .A2( u2_u10_u1_n184 ) );
  AOI21_X1 u2_u10_u1_U17 (.ZN( u2_u10_u1_n106 ) , .A( u2_u10_u1_n112 ) , .B1( u2_u10_u1_n154 ) , .B2( u2_u10_u1_n156 ) );
  AOI21_X1 u2_u10_u1_U18 (.ZN( u2_u10_u1_n107 ) , .B1( u2_u10_u1_n134 ) , .B2( u2_u10_u1_n149 ) , .A( u2_u10_u1_n174 ) );
  INV_X1 u2_u10_u1_U19 (.A( u2_u10_u1_n101 ) , .ZN( u2_u10_u1_n184 ) );
  INV_X1 u2_u10_u1_U20 (.A( u2_u10_u1_n112 ) , .ZN( u2_u10_u1_n171 ) );
  NAND2_X1 u2_u10_u1_U21 (.ZN( u2_u10_u1_n141 ) , .A1( u2_u10_u1_n153 ) , .A2( u2_u10_u1_n156 ) );
  AND2_X1 u2_u10_u1_U22 (.A1( u2_u10_u1_n123 ) , .ZN( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n161 ) );
  NAND2_X1 u2_u10_u1_U23 (.A2( u2_u10_u1_n115 ) , .A1( u2_u10_u1_n116 ) , .ZN( u2_u10_u1_n148 ) );
  NAND2_X1 u2_u10_u1_U24 (.A2( u2_u10_u1_n133 ) , .A1( u2_u10_u1_n135 ) , .ZN( u2_u10_u1_n159 ) );
  NAND2_X1 u2_u10_u1_U25 (.A2( u2_u10_u1_n115 ) , .A1( u2_u10_u1_n120 ) , .ZN( u2_u10_u1_n132 ) );
  INV_X1 u2_u10_u1_U26 (.A( u2_u10_u1_n154 ) , .ZN( u2_u10_u1_n178 ) );
  INV_X1 u2_u10_u1_U27 (.A( u2_u10_u1_n151 ) , .ZN( u2_u10_u1_n183 ) );
  AND2_X1 u2_u10_u1_U28 (.A1( u2_u10_u1_n129 ) , .A2( u2_u10_u1_n133 ) , .ZN( u2_u10_u1_n149 ) );
  INV_X1 u2_u10_u1_U29 (.A( u2_u10_u1_n131 ) , .ZN( u2_u10_u1_n180 ) );
  INV_X1 u2_u10_u1_U3 (.A( u2_u10_u1_n159 ) , .ZN( u2_u10_u1_n182 ) );
  OAI221_X1 u2_u10_u1_U30 (.A( u2_u10_u1_n119 ) , .C2( u2_u10_u1_n129 ) , .ZN( u2_u10_u1_n138 ) , .B2( u2_u10_u1_n152 ) , .C1( u2_u10_u1_n174 ) , .B1( u2_u10_u1_n187 ) );
  INV_X1 u2_u10_u1_U31 (.A( u2_u10_u1_n148 ) , .ZN( u2_u10_u1_n187 ) );
  AOI211_X1 u2_u10_u1_U32 (.B( u2_u10_u1_n117 ) , .A( u2_u10_u1_n118 ) , .ZN( u2_u10_u1_n119 ) , .C2( u2_u10_u1_n146 ) , .C1( u2_u10_u1_n159 ) );
  NOR2_X1 u2_u10_u1_U33 (.A1( u2_u10_u1_n168 ) , .A2( u2_u10_u1_n176 ) , .ZN( u2_u10_u1_n98 ) );
  OAI21_X1 u2_u10_u1_U34 (.B2( u2_u10_u1_n123 ) , .ZN( u2_u10_u1_n145 ) , .B1( u2_u10_u1_n160 ) , .A( u2_u10_u1_n185 ) );
  INV_X1 u2_u10_u1_U35 (.A( u2_u10_u1_n122 ) , .ZN( u2_u10_u1_n185 ) );
  AOI21_X1 u2_u10_u1_U36 (.B2( u2_u10_u1_n120 ) , .B1( u2_u10_u1_n121 ) , .ZN( u2_u10_u1_n122 ) , .A( u2_u10_u1_n128 ) );
  NAND2_X1 u2_u10_u1_U37 (.A1( u2_u10_u1_n128 ) , .ZN( u2_u10_u1_n146 ) , .A2( u2_u10_u1_n160 ) );
  NAND2_X1 u2_u10_u1_U38 (.A2( u2_u10_u1_n112 ) , .ZN( u2_u10_u1_n139 ) , .A1( u2_u10_u1_n152 ) );
  NAND2_X1 u2_u10_u1_U39 (.A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n156 ) , .A2( u2_u10_u1_n99 ) );
  AOI221_X1 u2_u10_u1_U4 (.A( u2_u10_u1_n138 ) , .C2( u2_u10_u1_n139 ) , .C1( u2_u10_u1_n140 ) , .B2( u2_u10_u1_n141 ) , .ZN( u2_u10_u1_n142 ) , .B1( u2_u10_u1_n175 ) );
  AOI221_X1 u2_u10_u1_U40 (.B1( u2_u10_u1_n140 ) , .ZN( u2_u10_u1_n167 ) , .B2( u2_u10_u1_n172 ) , .C2( u2_u10_u1_n175 ) , .C1( u2_u10_u1_n178 ) , .A( u2_u10_u1_n188 ) );
  INV_X1 u2_u10_u1_U41 (.ZN( u2_u10_u1_n188 ) , .A( u2_u10_u1_n97 ) );
  AOI211_X1 u2_u10_u1_U42 (.A( u2_u10_u1_n118 ) , .C1( u2_u10_u1_n132 ) , .C2( u2_u10_u1_n139 ) , .B( u2_u10_u1_n96 ) , .ZN( u2_u10_u1_n97 ) );
  AOI21_X1 u2_u10_u1_U43 (.B2( u2_u10_u1_n121 ) , .B1( u2_u10_u1_n135 ) , .A( u2_u10_u1_n152 ) , .ZN( u2_u10_u1_n96 ) );
  NOR2_X1 u2_u10_u1_U44 (.ZN( u2_u10_u1_n117 ) , .A1( u2_u10_u1_n121 ) , .A2( u2_u10_u1_n160 ) );
  AOI21_X1 u2_u10_u1_U45 (.A( u2_u10_u1_n128 ) , .B2( u2_u10_u1_n129 ) , .ZN( u2_u10_u1_n130 ) , .B1( u2_u10_u1_n150 ) );
  NAND2_X1 u2_u10_u1_U46 (.ZN( u2_u10_u1_n112 ) , .A1( u2_u10_u1_n169 ) , .A2( u2_u10_u1_n170 ) );
  NAND2_X1 u2_u10_u1_U47 (.ZN( u2_u10_u1_n129 ) , .A2( u2_u10_u1_n95 ) , .A1( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U48 (.A1( u2_u10_u1_n102 ) , .ZN( u2_u10_u1_n154 ) , .A2( u2_u10_u1_n99 ) );
  NAND2_X1 u2_u10_u1_U49 (.A2( u2_u10_u1_n100 ) , .ZN( u2_u10_u1_n135 ) , .A1( u2_u10_u1_n99 ) );
  AOI211_X1 u2_u10_u1_U5 (.ZN( u2_u10_u1_n124 ) , .A( u2_u10_u1_n138 ) , .C2( u2_u10_u1_n139 ) , .B( u2_u10_u1_n145 ) , .C1( u2_u10_u1_n147 ) );
  AOI21_X1 u2_u10_u1_U50 (.A( u2_u10_u1_n152 ) , .B2( u2_u10_u1_n153 ) , .B1( u2_u10_u1_n154 ) , .ZN( u2_u10_u1_n158 ) );
  INV_X1 u2_u10_u1_U51 (.A( u2_u10_u1_n160 ) , .ZN( u2_u10_u1_n175 ) );
  NAND2_X1 u2_u10_u1_U52 (.A1( u2_u10_u1_n100 ) , .ZN( u2_u10_u1_n116 ) , .A2( u2_u10_u1_n95 ) );
  NAND2_X1 u2_u10_u1_U53 (.A1( u2_u10_u1_n102 ) , .ZN( u2_u10_u1_n131 ) , .A2( u2_u10_u1_n95 ) );
  NAND2_X1 u2_u10_u1_U54 (.A2( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n121 ) , .A1( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U55 (.A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n153 ) , .A2( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U56 (.A2( u2_u10_u1_n104 ) , .A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n133 ) );
  NAND2_X1 u2_u10_u1_U57 (.ZN( u2_u10_u1_n150 ) , .A2( u2_u10_u1_n98 ) , .A1( u2_u10_u1_n99 ) );
  NAND2_X1 u2_u10_u1_U58 (.A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n155 ) , .A2( u2_u10_u1_n95 ) );
  OAI21_X1 u2_u10_u1_U59 (.ZN( u2_u10_u1_n109 ) , .B1( u2_u10_u1_n129 ) , .B2( u2_u10_u1_n160 ) , .A( u2_u10_u1_n167 ) );
  AOI22_X1 u2_u10_u1_U6 (.B2( u2_u10_u1_n113 ) , .A2( u2_u10_u1_n114 ) , .ZN( u2_u10_u1_n125 ) , .A1( u2_u10_u1_n171 ) , .B1( u2_u10_u1_n173 ) );
  NAND2_X1 u2_u10_u1_U60 (.A2( u2_u10_u1_n100 ) , .A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n120 ) );
  NAND2_X1 u2_u10_u1_U61 (.A1( u2_u10_u1_n102 ) , .A2( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n115 ) );
  NAND2_X1 u2_u10_u1_U62 (.A2( u2_u10_u1_n100 ) , .A1( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n151 ) );
  NAND2_X1 u2_u10_u1_U63 (.A2( u2_u10_u1_n103 ) , .A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n161 ) );
  INV_X1 u2_u10_u1_U64 (.A( u2_u10_u1_n152 ) , .ZN( u2_u10_u1_n173 ) );
  INV_X1 u2_u10_u1_U65 (.A( u2_u10_u1_n128 ) , .ZN( u2_u10_u1_n172 ) );
  NAND2_X1 u2_u10_u1_U66 (.A2( u2_u10_u1_n102 ) , .A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n123 ) );
  AOI211_X1 u2_u10_u1_U67 (.B( u2_u10_u1_n162 ) , .A( u2_u10_u1_n163 ) , .C2( u2_u10_u1_n164 ) , .ZN( u2_u10_u1_n165 ) , .C1( u2_u10_u1_n171 ) );
  AOI21_X1 u2_u10_u1_U68 (.A( u2_u10_u1_n160 ) , .B2( u2_u10_u1_n161 ) , .ZN( u2_u10_u1_n162 ) , .B1( u2_u10_u1_n182 ) );
  OR2_X1 u2_u10_u1_U69 (.A2( u2_u10_u1_n157 ) , .A1( u2_u10_u1_n158 ) , .ZN( u2_u10_u1_n163 ) );
  NAND2_X1 u2_u10_u1_U7 (.ZN( u2_u10_u1_n114 ) , .A1( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n156 ) );
  NOR2_X1 u2_u10_u1_U70 (.A2( u2_u10_X_7 ) , .A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n95 ) );
  NOR2_X1 u2_u10_u1_U71 (.A1( u2_u10_X_12 ) , .A2( u2_u10_X_9 ) , .ZN( u2_u10_u1_n100 ) );
  NOR2_X1 u2_u10_u1_U72 (.A2( u2_u10_X_8 ) , .A1( u2_u10_u1_n177 ) , .ZN( u2_u10_u1_n99 ) );
  NOR2_X1 u2_u10_u1_U73 (.A2( u2_u10_X_12 ) , .ZN( u2_u10_u1_n102 ) , .A1( u2_u10_u1_n176 ) );
  NOR2_X1 u2_u10_u1_U74 (.A2( u2_u10_X_9 ) , .ZN( u2_u10_u1_n105 ) , .A1( u2_u10_u1_n168 ) );
  NAND2_X1 u2_u10_u1_U75 (.A1( u2_u10_X_10 ) , .ZN( u2_u10_u1_n160 ) , .A2( u2_u10_u1_n169 ) );
  NAND2_X1 u2_u10_u1_U76 (.A2( u2_u10_X_10 ) , .A1( u2_u10_X_11 ) , .ZN( u2_u10_u1_n152 ) );
  NAND2_X1 u2_u10_u1_U77 (.A1( u2_u10_X_11 ) , .ZN( u2_u10_u1_n128 ) , .A2( u2_u10_u1_n170 ) );
  AND2_X1 u2_u10_u1_U78 (.A2( u2_u10_X_7 ) , .A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n104 ) );
  AND2_X1 u2_u10_u1_U79 (.A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n103 ) , .A2( u2_u10_u1_n177 ) );
  NOR2_X1 u2_u10_u1_U8 (.A1( u2_u10_u1_n112 ) , .A2( u2_u10_u1_n116 ) , .ZN( u2_u10_u1_n118 ) );
  INV_X1 u2_u10_u1_U80 (.A( u2_u10_X_10 ) , .ZN( u2_u10_u1_n170 ) );
  INV_X1 u2_u10_u1_U81 (.A( u2_u10_X_9 ) , .ZN( u2_u10_u1_n176 ) );
  INV_X1 u2_u10_u1_U82 (.A( u2_u10_X_11 ) , .ZN( u2_u10_u1_n169 ) );
  INV_X1 u2_u10_u1_U83 (.A( u2_u10_X_12 ) , .ZN( u2_u10_u1_n168 ) );
  INV_X1 u2_u10_u1_U84 (.A( u2_u10_X_7 ) , .ZN( u2_u10_u1_n177 ) );
  NAND4_X1 u2_u10_u1_U85 (.ZN( u2_out10_28 ) , .A4( u2_u10_u1_n124 ) , .A3( u2_u10_u1_n125 ) , .A2( u2_u10_u1_n126 ) , .A1( u2_u10_u1_n127 ) );
  OAI21_X1 u2_u10_u1_U86 (.ZN( u2_u10_u1_n127 ) , .B2( u2_u10_u1_n139 ) , .B1( u2_u10_u1_n175 ) , .A( u2_u10_u1_n183 ) );
  OAI21_X1 u2_u10_u1_U87 (.ZN( u2_u10_u1_n126 ) , .B2( u2_u10_u1_n140 ) , .A( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n178 ) );
  NAND4_X1 u2_u10_u1_U88 (.ZN( u2_out10_18 ) , .A4( u2_u10_u1_n165 ) , .A3( u2_u10_u1_n166 ) , .A1( u2_u10_u1_n167 ) , .A2( u2_u10_u1_n186 ) );
  AOI22_X1 u2_u10_u1_U89 (.B2( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n147 ) , .A2( u2_u10_u1_n148 ) , .ZN( u2_u10_u1_n166 ) , .A1( u2_u10_u1_n172 ) );
  OAI21_X1 u2_u10_u1_U9 (.ZN( u2_u10_u1_n101 ) , .B1( u2_u10_u1_n141 ) , .A( u2_u10_u1_n146 ) , .B2( u2_u10_u1_n183 ) );
  INV_X1 u2_u10_u1_U90 (.A( u2_u10_u1_n145 ) , .ZN( u2_u10_u1_n186 ) );
  NAND4_X1 u2_u10_u1_U91 (.ZN( u2_out10_2 ) , .A4( u2_u10_u1_n142 ) , .A3( u2_u10_u1_n143 ) , .A2( u2_u10_u1_n144 ) , .A1( u2_u10_u1_n179 ) );
  OAI21_X1 u2_u10_u1_U92 (.B2( u2_u10_u1_n132 ) , .ZN( u2_u10_u1_n144 ) , .A( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n180 ) );
  INV_X1 u2_u10_u1_U93 (.A( u2_u10_u1_n130 ) , .ZN( u2_u10_u1_n179 ) );
  OR4_X1 u2_u10_u1_U94 (.ZN( u2_out10_13 ) , .A4( u2_u10_u1_n108 ) , .A3( u2_u10_u1_n109 ) , .A2( u2_u10_u1_n110 ) , .A1( u2_u10_u1_n111 ) );
  AOI21_X1 u2_u10_u1_U95 (.ZN( u2_u10_u1_n111 ) , .A( u2_u10_u1_n128 ) , .B2( u2_u10_u1_n131 ) , .B1( u2_u10_u1_n135 ) );
  AOI21_X1 u2_u10_u1_U96 (.ZN( u2_u10_u1_n110 ) , .A( u2_u10_u1_n116 ) , .B1( u2_u10_u1_n152 ) , .B2( u2_u10_u1_n160 ) );
  NAND3_X1 u2_u10_u1_U97 (.A3( u2_u10_u1_n149 ) , .A2( u2_u10_u1_n150 ) , .A1( u2_u10_u1_n151 ) , .ZN( u2_u10_u1_n164 ) );
  NAND3_X1 u2_u10_u1_U98 (.A3( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n135 ) , .ZN( u2_u10_u1_n136 ) , .A1( u2_u10_u1_n151 ) );
  NAND3_X1 u2_u10_u1_U99 (.A1( u2_u10_u1_n133 ) , .ZN( u2_u10_u1_n137 ) , .A2( u2_u10_u1_n154 ) , .A3( u2_u10_u1_n181 ) );
  OAI22_X1 u2_u10_u2_U10 (.ZN( u2_u10_u2_n109 ) , .A2( u2_u10_u2_n113 ) , .B2( u2_u10_u2_n133 ) , .B1( u2_u10_u2_n167 ) , .A1( u2_u10_u2_n168 ) );
  NAND3_X1 u2_u10_u2_U100 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n98 ) );
  OAI22_X1 u2_u10_u2_U11 (.B1( u2_u10_u2_n151 ) , .A2( u2_u10_u2_n152 ) , .A1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n160 ) , .B2( u2_u10_u2_n168 ) );
  NOR3_X1 u2_u10_u2_U12 (.A1( u2_u10_u2_n150 ) , .ZN( u2_u10_u2_n151 ) , .A3( u2_u10_u2_n175 ) , .A2( u2_u10_u2_n188 ) );
  AOI21_X1 u2_u10_u2_U13 (.ZN( u2_u10_u2_n144 ) , .B2( u2_u10_u2_n155 ) , .A( u2_u10_u2_n172 ) , .B1( u2_u10_u2_n185 ) );
  AOI21_X1 u2_u10_u2_U14 (.B2( u2_u10_u2_n143 ) , .ZN( u2_u10_u2_n145 ) , .B1( u2_u10_u2_n152 ) , .A( u2_u10_u2_n171 ) );
  AOI21_X1 u2_u10_u2_U15 (.B2( u2_u10_u2_n120 ) , .B1( u2_u10_u2_n121 ) , .ZN( u2_u10_u2_n126 ) , .A( u2_u10_u2_n167 ) );
  INV_X1 u2_u10_u2_U16 (.A( u2_u10_u2_n156 ) , .ZN( u2_u10_u2_n171 ) );
  INV_X1 u2_u10_u2_U17 (.A( u2_u10_u2_n120 ) , .ZN( u2_u10_u2_n188 ) );
  NAND2_X1 u2_u10_u2_U18 (.A2( u2_u10_u2_n122 ) , .ZN( u2_u10_u2_n150 ) , .A1( u2_u10_u2_n152 ) );
  INV_X1 u2_u10_u2_U19 (.A( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n170 ) );
  INV_X1 u2_u10_u2_U20 (.A( u2_u10_u2_n137 ) , .ZN( u2_u10_u2_n173 ) );
  NAND2_X1 u2_u10_u2_U21 (.A1( u2_u10_u2_n132 ) , .A2( u2_u10_u2_n139 ) , .ZN( u2_u10_u2_n157 ) );
  INV_X1 u2_u10_u2_U22 (.A( u2_u10_u2_n113 ) , .ZN( u2_u10_u2_n178 ) );
  INV_X1 u2_u10_u2_U23 (.A( u2_u10_u2_n139 ) , .ZN( u2_u10_u2_n175 ) );
  INV_X1 u2_u10_u2_U24 (.A( u2_u10_u2_n155 ) , .ZN( u2_u10_u2_n181 ) );
  INV_X1 u2_u10_u2_U25 (.A( u2_u10_u2_n119 ) , .ZN( u2_u10_u2_n177 ) );
  INV_X1 u2_u10_u2_U26 (.A( u2_u10_u2_n116 ) , .ZN( u2_u10_u2_n180 ) );
  INV_X1 u2_u10_u2_U27 (.A( u2_u10_u2_n131 ) , .ZN( u2_u10_u2_n179 ) );
  INV_X1 u2_u10_u2_U28 (.A( u2_u10_u2_n154 ) , .ZN( u2_u10_u2_n176 ) );
  NAND2_X1 u2_u10_u2_U29 (.A2( u2_u10_u2_n116 ) , .A1( u2_u10_u2_n117 ) , .ZN( u2_u10_u2_n118 ) );
  NOR2_X1 u2_u10_u2_U3 (.ZN( u2_u10_u2_n121 ) , .A2( u2_u10_u2_n177 ) , .A1( u2_u10_u2_n180 ) );
  INV_X1 u2_u10_u2_U30 (.A( u2_u10_u2_n132 ) , .ZN( u2_u10_u2_n182 ) );
  INV_X1 u2_u10_u2_U31 (.A( u2_u10_u2_n158 ) , .ZN( u2_u10_u2_n183 ) );
  OAI21_X1 u2_u10_u2_U32 (.A( u2_u10_u2_n156 ) , .B1( u2_u10_u2_n157 ) , .ZN( u2_u10_u2_n158 ) , .B2( u2_u10_u2_n179 ) );
  NOR2_X1 u2_u10_u2_U33 (.ZN( u2_u10_u2_n156 ) , .A1( u2_u10_u2_n166 ) , .A2( u2_u10_u2_n169 ) );
  NOR2_X1 u2_u10_u2_U34 (.A2( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n137 ) , .A1( u2_u10_u2_n140 ) );
  NOR2_X1 u2_u10_u2_U35 (.A2( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n153 ) , .A1( u2_u10_u2_n156 ) );
  AOI211_X1 u2_u10_u2_U36 (.ZN( u2_u10_u2_n130 ) , .C1( u2_u10_u2_n138 ) , .C2( u2_u10_u2_n179 ) , .B( u2_u10_u2_n96 ) , .A( u2_u10_u2_n97 ) );
  OAI22_X1 u2_u10_u2_U37 (.B1( u2_u10_u2_n133 ) , .A2( u2_u10_u2_n137 ) , .A1( u2_u10_u2_n152 ) , .B2( u2_u10_u2_n168 ) , .ZN( u2_u10_u2_n97 ) );
  OAI221_X1 u2_u10_u2_U38 (.B1( u2_u10_u2_n113 ) , .C1( u2_u10_u2_n132 ) , .A( u2_u10_u2_n149 ) , .B2( u2_u10_u2_n171 ) , .C2( u2_u10_u2_n172 ) , .ZN( u2_u10_u2_n96 ) );
  OAI221_X1 u2_u10_u2_U39 (.A( u2_u10_u2_n115 ) , .C2( u2_u10_u2_n123 ) , .B2( u2_u10_u2_n143 ) , .B1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n163 ) , .C1( u2_u10_u2_n168 ) );
  INV_X1 u2_u10_u2_U4 (.A( u2_u10_u2_n134 ) , .ZN( u2_u10_u2_n185 ) );
  OAI21_X1 u2_u10_u2_U40 (.A( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n115 ) , .B1( u2_u10_u2_n176 ) , .B2( u2_u10_u2_n178 ) );
  OAI221_X1 u2_u10_u2_U41 (.A( u2_u10_u2_n135 ) , .B2( u2_u10_u2_n136 ) , .B1( u2_u10_u2_n137 ) , .ZN( u2_u10_u2_n162 ) , .C2( u2_u10_u2_n167 ) , .C1( u2_u10_u2_n185 ) );
  AND3_X1 u2_u10_u2_U42 (.A3( u2_u10_u2_n131 ) , .A2( u2_u10_u2_n132 ) , .A1( u2_u10_u2_n133 ) , .ZN( u2_u10_u2_n136 ) );
  AOI22_X1 u2_u10_u2_U43 (.ZN( u2_u10_u2_n135 ) , .B1( u2_u10_u2_n140 ) , .A1( u2_u10_u2_n156 ) , .B2( u2_u10_u2_n180 ) , .A2( u2_u10_u2_n188 ) );
  AOI21_X1 u2_u10_u2_U44 (.ZN( u2_u10_u2_n149 ) , .B1( u2_u10_u2_n173 ) , .B2( u2_u10_u2_n188 ) , .A( u2_u10_u2_n95 ) );
  AND3_X1 u2_u10_u2_U45 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n156 ) , .ZN( u2_u10_u2_n95 ) );
  OAI21_X1 u2_u10_u2_U46 (.A( u2_u10_u2_n141 ) , .B2( u2_u10_u2_n142 ) , .ZN( u2_u10_u2_n146 ) , .B1( u2_u10_u2_n153 ) );
  OAI21_X1 u2_u10_u2_U47 (.A( u2_u10_u2_n140 ) , .ZN( u2_u10_u2_n141 ) , .B1( u2_u10_u2_n176 ) , .B2( u2_u10_u2_n177 ) );
  NOR3_X1 u2_u10_u2_U48 (.ZN( u2_u10_u2_n142 ) , .A3( u2_u10_u2_n175 ) , .A2( u2_u10_u2_n178 ) , .A1( u2_u10_u2_n181 ) );
  OAI21_X1 u2_u10_u2_U49 (.A( u2_u10_u2_n101 ) , .B2( u2_u10_u2_n121 ) , .B1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n164 ) );
  INV_X1 u2_u10_u2_U5 (.A( u2_u10_u2_n150 ) , .ZN( u2_u10_u2_n184 ) );
  NAND2_X1 u2_u10_u2_U50 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n155 ) );
  NAND2_X1 u2_u10_u2_U51 (.A2( u2_u10_u2_n105 ) , .A1( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n143 ) );
  NAND2_X1 u2_u10_u2_U52 (.A1( u2_u10_u2_n104 ) , .A2( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n152 ) );
  NAND2_X1 u2_u10_u2_U53 (.A1( u2_u10_u2_n100 ) , .A2( u2_u10_u2_n105 ) , .ZN( u2_u10_u2_n132 ) );
  INV_X1 u2_u10_u2_U54 (.A( u2_u10_u2_n140 ) , .ZN( u2_u10_u2_n168 ) );
  INV_X1 u2_u10_u2_U55 (.A( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n167 ) );
  NAND2_X1 u2_u10_u2_U56 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n113 ) );
  NAND2_X1 u2_u10_u2_U57 (.A1( u2_u10_u2_n106 ) , .A2( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n131 ) );
  NAND2_X1 u2_u10_u2_U58 (.A1( u2_u10_u2_n103 ) , .A2( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n139 ) );
  NAND2_X1 u2_u10_u2_U59 (.A1( u2_u10_u2_n103 ) , .A2( u2_u10_u2_n105 ) , .ZN( u2_u10_u2_n133 ) );
  NOR4_X1 u2_u10_u2_U6 (.A4( u2_u10_u2_n124 ) , .A3( u2_u10_u2_n125 ) , .A2( u2_u10_u2_n126 ) , .A1( u2_u10_u2_n127 ) , .ZN( u2_u10_u2_n128 ) );
  NAND2_X1 u2_u10_u2_U60 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n103 ) , .ZN( u2_u10_u2_n154 ) );
  NAND2_X1 u2_u10_u2_U61 (.A2( u2_u10_u2_n103 ) , .A1( u2_u10_u2_n104 ) , .ZN( u2_u10_u2_n119 ) );
  NAND2_X1 u2_u10_u2_U62 (.A2( u2_u10_u2_n107 ) , .A1( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n123 ) );
  NAND2_X1 u2_u10_u2_U63 (.A1( u2_u10_u2_n104 ) , .A2( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n122 ) );
  INV_X1 u2_u10_u2_U64 (.A( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n172 ) );
  NAND2_X1 u2_u10_u2_U65 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n102 ) , .ZN( u2_u10_u2_n116 ) );
  NAND2_X1 u2_u10_u2_U66 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n120 ) );
  NAND2_X1 u2_u10_u2_U67 (.A2( u2_u10_u2_n105 ) , .A1( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n117 ) );
  INV_X1 u2_u10_u2_U68 (.ZN( u2_u10_u2_n187 ) , .A( u2_u10_u2_n99 ) );
  OAI21_X1 u2_u10_u2_U69 (.B1( u2_u10_u2_n137 ) , .B2( u2_u10_u2_n143 ) , .A( u2_u10_u2_n98 ) , .ZN( u2_u10_u2_n99 ) );
  AOI21_X1 u2_u10_u2_U7 (.ZN( u2_u10_u2_n124 ) , .B1( u2_u10_u2_n131 ) , .B2( u2_u10_u2_n143 ) , .A( u2_u10_u2_n172 ) );
  NOR2_X1 u2_u10_u2_U70 (.A2( u2_u10_X_16 ) , .ZN( u2_u10_u2_n140 ) , .A1( u2_u10_u2_n166 ) );
  NOR2_X1 u2_u10_u2_U71 (.A2( u2_u10_X_13 ) , .A1( u2_u10_X_14 ) , .ZN( u2_u10_u2_n100 ) );
  NOR2_X1 u2_u10_u2_U72 (.A2( u2_u10_X_16 ) , .A1( u2_u10_X_17 ) , .ZN( u2_u10_u2_n138 ) );
  NOR2_X1 u2_u10_u2_U73 (.A2( u2_u10_X_15 ) , .A1( u2_u10_X_18 ) , .ZN( u2_u10_u2_n104 ) );
  NOR2_X1 u2_u10_u2_U74 (.A2( u2_u10_X_14 ) , .ZN( u2_u10_u2_n103 ) , .A1( u2_u10_u2_n174 ) );
  NOR2_X1 u2_u10_u2_U75 (.A2( u2_u10_X_15 ) , .ZN( u2_u10_u2_n102 ) , .A1( u2_u10_u2_n165 ) );
  NOR2_X1 u2_u10_u2_U76 (.A2( u2_u10_X_17 ) , .ZN( u2_u10_u2_n114 ) , .A1( u2_u10_u2_n169 ) );
  AND2_X1 u2_u10_u2_U77 (.A1( u2_u10_X_15 ) , .ZN( u2_u10_u2_n105 ) , .A2( u2_u10_u2_n165 ) );
  AND2_X1 u2_u10_u2_U78 (.A2( u2_u10_X_15 ) , .A1( u2_u10_X_18 ) , .ZN( u2_u10_u2_n107 ) );
  AND2_X1 u2_u10_u2_U79 (.A1( u2_u10_X_14 ) , .ZN( u2_u10_u2_n106 ) , .A2( u2_u10_u2_n174 ) );
  AOI21_X1 u2_u10_u2_U8 (.B2( u2_u10_u2_n119 ) , .ZN( u2_u10_u2_n127 ) , .A( u2_u10_u2_n137 ) , .B1( u2_u10_u2_n155 ) );
  AND2_X1 u2_u10_u2_U80 (.A1( u2_u10_X_13 ) , .A2( u2_u10_X_14 ) , .ZN( u2_u10_u2_n108 ) );
  INV_X1 u2_u10_u2_U81 (.A( u2_u10_X_16 ) , .ZN( u2_u10_u2_n169 ) );
  INV_X1 u2_u10_u2_U82 (.A( u2_u10_X_17 ) , .ZN( u2_u10_u2_n166 ) );
  INV_X1 u2_u10_u2_U83 (.A( u2_u10_X_13 ) , .ZN( u2_u10_u2_n174 ) );
  INV_X1 u2_u10_u2_U84 (.A( u2_u10_X_18 ) , .ZN( u2_u10_u2_n165 ) );
  NAND4_X1 u2_u10_u2_U85 (.ZN( u2_out10_24 ) , .A4( u2_u10_u2_n111 ) , .A3( u2_u10_u2_n112 ) , .A1( u2_u10_u2_n130 ) , .A2( u2_u10_u2_n187 ) );
  AOI221_X1 u2_u10_u2_U86 (.A( u2_u10_u2_n109 ) , .B1( u2_u10_u2_n110 ) , .ZN( u2_u10_u2_n111 ) , .C1( u2_u10_u2_n134 ) , .C2( u2_u10_u2_n170 ) , .B2( u2_u10_u2_n173 ) );
  AOI21_X1 u2_u10_u2_U87 (.ZN( u2_u10_u2_n112 ) , .B2( u2_u10_u2_n156 ) , .A( u2_u10_u2_n164 ) , .B1( u2_u10_u2_n181 ) );
  NAND4_X1 u2_u10_u2_U88 (.ZN( u2_out10_16 ) , .A4( u2_u10_u2_n128 ) , .A3( u2_u10_u2_n129 ) , .A1( u2_u10_u2_n130 ) , .A2( u2_u10_u2_n186 ) );
  AOI22_X1 u2_u10_u2_U89 (.A2( u2_u10_u2_n118 ) , .ZN( u2_u10_u2_n129 ) , .A1( u2_u10_u2_n140 ) , .B1( u2_u10_u2_n157 ) , .B2( u2_u10_u2_n170 ) );
  AOI21_X1 u2_u10_u2_U9 (.B2( u2_u10_u2_n123 ) , .ZN( u2_u10_u2_n125 ) , .A( u2_u10_u2_n171 ) , .B1( u2_u10_u2_n184 ) );
  INV_X1 u2_u10_u2_U90 (.A( u2_u10_u2_n163 ) , .ZN( u2_u10_u2_n186 ) );
  NAND4_X1 u2_u10_u2_U91 (.ZN( u2_out10_30 ) , .A4( u2_u10_u2_n147 ) , .A3( u2_u10_u2_n148 ) , .A2( u2_u10_u2_n149 ) , .A1( u2_u10_u2_n187 ) );
  NOR3_X1 u2_u10_u2_U92 (.A3( u2_u10_u2_n144 ) , .A2( u2_u10_u2_n145 ) , .A1( u2_u10_u2_n146 ) , .ZN( u2_u10_u2_n147 ) );
  AOI21_X1 u2_u10_u2_U93 (.B2( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n148 ) , .A( u2_u10_u2_n162 ) , .B1( u2_u10_u2_n182 ) );
  OR4_X1 u2_u10_u2_U94 (.ZN( u2_out10_6 ) , .A4( u2_u10_u2_n161 ) , .A3( u2_u10_u2_n162 ) , .A2( u2_u10_u2_n163 ) , .A1( u2_u10_u2_n164 ) );
  OR3_X1 u2_u10_u2_U95 (.A2( u2_u10_u2_n159 ) , .A1( u2_u10_u2_n160 ) , .ZN( u2_u10_u2_n161 ) , .A3( u2_u10_u2_n183 ) );
  AOI21_X1 u2_u10_u2_U96 (.B2( u2_u10_u2_n154 ) , .B1( u2_u10_u2_n155 ) , .ZN( u2_u10_u2_n159 ) , .A( u2_u10_u2_n167 ) );
  NAND3_X1 u2_u10_u2_U97 (.A2( u2_u10_u2_n117 ) , .A1( u2_u10_u2_n122 ) , .A3( u2_u10_u2_n123 ) , .ZN( u2_u10_u2_n134 ) );
  NAND3_X1 u2_u10_u2_U98 (.ZN( u2_u10_u2_n110 ) , .A2( u2_u10_u2_n131 ) , .A3( u2_u10_u2_n139 ) , .A1( u2_u10_u2_n154 ) );
  NAND3_X1 u2_u10_u2_U99 (.A2( u2_u10_u2_n100 ) , .ZN( u2_u10_u2_n101 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n114 ) );
  XOR2_X1 u2_u15_U11 (.A( u2_FP_61 ) , .B( u2_K16_44 ) , .Z( u2_u15_X_44 ) );
  XOR2_X1 u2_u15_U12 (.A( u2_FP_60 ) , .B( u2_K16_43 ) , .Z( u2_u15_X_43 ) );
  XOR2_X1 u2_u15_U13 (.A( u2_FP_61 ) , .B( u2_K16_42 ) , .Z( u2_u15_X_42 ) );
  XOR2_X1 u2_u15_U14 (.A( u2_FP_60 ) , .B( u2_K16_41 ) , .Z( u2_u15_X_41 ) );
  XOR2_X1 u2_u15_U18 (.A( u2_FP_57 ) , .B( u2_K16_38 ) , .Z( u2_u15_X_38 ) );
  XOR2_X1 u2_u15_U19 (.A( u2_FP_56 ) , .B( u2_K16_37 ) , .Z( u2_u15_X_37 ) );
  XOR2_X1 u2_u15_U2 (.A( u2_FP_37 ) , .B( u2_K16_8 ) , .Z( u2_u15_X_8 ) );
  XOR2_X1 u2_u15_U20 (.A( u2_FP_57 ) , .B( u2_K16_36 ) , .Z( u2_u15_X_36 ) );
  XOR2_X1 u2_u15_U21 (.A( u2_FP_56 ) , .B( u2_K16_35 ) , .Z( u2_u15_X_35 ) );
  XOR2_X1 u2_u15_U22 (.A( u2_FP_55 ) , .B( u2_K16_34 ) , .Z( u2_u15_X_34 ) );
  XOR2_X1 u2_u15_U24 (.A( u2_FP_53 ) , .B( u2_K16_32 ) , .Z( u2_u15_X_32 ) );
  XOR2_X1 u2_u15_U25 (.A( u2_FP_52 ) , .B( u2_K16_31 ) , .Z( u2_u15_X_31 ) );
  XOR2_X1 u2_u15_U26 (.A( u2_FP_53 ) , .B( u2_K16_30 ) , .Z( u2_u15_X_30 ) );
  XOR2_X1 u2_u15_U27 (.A( u2_FP_33 ) , .B( u2_K16_2 ) , .Z( u2_u15_X_2 ) );
  XOR2_X1 u2_u15_U28 (.A( u2_FP_52 ) , .B( u2_K16_29 ) , .Z( u2_u15_X_29 ) );
  XOR2_X1 u2_u15_U3 (.A( u2_FP_36 ) , .B( u2_K16_7 ) , .Z( u2_u15_X_7 ) );
  XOR2_X1 u2_u15_U31 (.A( u2_FP_49 ) , .B( u2_K16_26 ) , .Z( u2_u15_X_26 ) );
  XOR2_X1 u2_u15_U32 (.A( u2_FP_48 ) , .B( u2_K16_25 ) , .Z( u2_u15_X_25 ) );
  XOR2_X1 u2_u15_U33 (.A( u2_FP_49 ) , .B( u2_K16_24 ) , .Z( u2_u15_X_24 ) );
  XOR2_X1 u2_u15_U34 (.A( u2_FP_48 ) , .B( u2_K16_23 ) , .Z( u2_u15_X_23 ) );
  XOR2_X1 u2_u15_U37 (.A( u2_FP_45 ) , .B( u2_K16_20 ) , .Z( u2_u15_X_20 ) );
  XOR2_X1 u2_u15_U38 (.A( u2_FP_64 ) , .B( u2_K16_1 ) , .Z( u2_u15_X_1 ) );
  XOR2_X1 u2_u15_U39 (.A( u2_FP_44 ) , .B( u2_K16_19 ) , .Z( u2_u15_X_19 ) );
  XOR2_X1 u2_u15_U4 (.A( u2_FP_37 ) , .B( u2_K16_6 ) , .Z( u2_u15_X_6 ) );
  XOR2_X1 u2_u15_U40 (.A( u2_FP_45 ) , .B( u2_K16_18 ) , .Z( u2_u15_X_18 ) );
  XOR2_X1 u2_u15_U41 (.A( u2_FP_44 ) , .B( u2_K16_17 ) , .Z( u2_u15_X_17 ) );
  XOR2_X1 u2_u15_U44 (.A( u2_FP_41 ) , .B( u2_K16_14 ) , .Z( u2_u15_X_14 ) );
  XOR2_X1 u2_u15_U45 (.A( u2_FP_40 ) , .B( u2_K16_13 ) , .Z( u2_u15_X_13 ) );
  XOR2_X1 u2_u15_U46 (.A( u2_FP_41 ) , .B( u2_K16_12 ) , .Z( u2_u15_X_12 ) );
  XOR2_X1 u2_u15_U47 (.A( u2_FP_40 ) , .B( u2_K16_11 ) , .Z( u2_u15_X_11 ) );
  XOR2_X1 u2_u15_U5 (.A( u2_FP_36 ) , .B( u2_K16_5 ) , .Z( u2_u15_X_5 ) );
  XOR2_X1 u2_u15_U7 (.A( u2_FP_33 ) , .B( u2_K16_48 ) , .Z( u2_u15_X_48 ) );
  XOR2_X1 u2_u15_U8 (.A( u2_FP_64 ) , .B( u2_K16_47 ) , .Z( u2_u15_X_47 ) );
  AND3_X1 u2_u15_u0_U10 (.A2( u2_u15_u0_n112 ) , .ZN( u2_u15_u0_n127 ) , .A3( u2_u15_u0_n130 ) , .A1( u2_u15_u0_n148 ) );
  NAND2_X1 u2_u15_u0_U11 (.ZN( u2_u15_u0_n113 ) , .A1( u2_u15_u0_n139 ) , .A2( u2_u15_u0_n149 ) );
  AND2_X1 u2_u15_u0_U12 (.ZN( u2_u15_u0_n107 ) , .A1( u2_u15_u0_n130 ) , .A2( u2_u15_u0_n140 ) );
  AND2_X1 u2_u15_u0_U13 (.A2( u2_u15_u0_n129 ) , .A1( u2_u15_u0_n130 ) , .ZN( u2_u15_u0_n151 ) );
  AND2_X1 u2_u15_u0_U14 (.A1( u2_u15_u0_n108 ) , .A2( u2_u15_u0_n125 ) , .ZN( u2_u15_u0_n145 ) );
  INV_X1 u2_u15_u0_U15 (.A( u2_u15_u0_n143 ) , .ZN( u2_u15_u0_n173 ) );
  NOR2_X1 u2_u15_u0_U16 (.A2( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n147 ) , .A1( u2_u15_u0_n160 ) );
  AOI21_X1 u2_u15_u0_U17 (.B1( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n132 ) , .A( u2_u15_u0_n165 ) , .B2( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U18 (.A( u2_u15_u0_n142 ) , .ZN( u2_u15_u0_n165 ) );
  OAI221_X1 u2_u15_u0_U19 (.C1( u2_u15_u0_n112 ) , .ZN( u2_u15_u0_n120 ) , .B1( u2_u15_u0_n138 ) , .B2( u2_u15_u0_n141 ) , .C2( u2_u15_u0_n147 ) , .A( u2_u15_u0_n172 ) );
  AOI211_X1 u2_u15_u0_U20 (.B( u2_u15_u0_n115 ) , .A( u2_u15_u0_n116 ) , .C2( u2_u15_u0_n117 ) , .C1( u2_u15_u0_n118 ) , .ZN( u2_u15_u0_n119 ) );
  OAI22_X1 u2_u15_u0_U21 (.B1( u2_u15_u0_n125 ) , .ZN( u2_u15_u0_n126 ) , .A1( u2_u15_u0_n138 ) , .A2( u2_u15_u0_n146 ) , .B2( u2_u15_u0_n147 ) );
  OAI22_X1 u2_u15_u0_U22 (.B1( u2_u15_u0_n131 ) , .A1( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n147 ) , .A2( u2_u15_u0_n90 ) , .ZN( u2_u15_u0_n91 ) );
  AND3_X1 u2_u15_u0_U23 (.A3( u2_u15_u0_n121 ) , .A2( u2_u15_u0_n125 ) , .A1( u2_u15_u0_n148 ) , .ZN( u2_u15_u0_n90 ) );
  INV_X1 u2_u15_u0_U24 (.A( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n161 ) );
  AOI22_X1 u2_u15_u0_U25 (.B2( u2_u15_u0_n109 ) , .A2( u2_u15_u0_n110 ) , .ZN( u2_u15_u0_n111 ) , .B1( u2_u15_u0_n118 ) , .A1( u2_u15_u0_n160 ) );
  INV_X1 u2_u15_u0_U26 (.A( u2_u15_u0_n118 ) , .ZN( u2_u15_u0_n158 ) );
  AOI21_X1 u2_u15_u0_U27 (.ZN( u2_u15_u0_n104 ) , .B1( u2_u15_u0_n107 ) , .B2( u2_u15_u0_n141 ) , .A( u2_u15_u0_n144 ) );
  AOI21_X1 u2_u15_u0_U28 (.B1( u2_u15_u0_n127 ) , .B2( u2_u15_u0_n129 ) , .A( u2_u15_u0_n138 ) , .ZN( u2_u15_u0_n96 ) );
  AOI21_X1 u2_u15_u0_U29 (.ZN( u2_u15_u0_n116 ) , .B2( u2_u15_u0_n142 ) , .A( u2_u15_u0_n144 ) , .B1( u2_u15_u0_n166 ) );
  INV_X1 u2_u15_u0_U3 (.A( u2_u15_u0_n113 ) , .ZN( u2_u15_u0_n166 ) );
  NAND2_X1 u2_u15_u0_U30 (.A1( u2_u15_u0_n100 ) , .A2( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n125 ) );
  NAND2_X1 u2_u15_u0_U31 (.A2( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n140 ) , .A1( u2_u15_u0_n94 ) );
  NAND2_X1 u2_u15_u0_U32 (.A1( u2_u15_u0_n101 ) , .A2( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n150 ) );
  INV_X1 u2_u15_u0_U33 (.A( u2_u15_u0_n138 ) , .ZN( u2_u15_u0_n160 ) );
  NAND2_X1 u2_u15_u0_U34 (.A2( u2_u15_u0_n102 ) , .A1( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n149 ) );
  NAND2_X1 u2_u15_u0_U35 (.A2( u2_u15_u0_n100 ) , .A1( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n139 ) );
  NAND2_X1 u2_u15_u0_U36 (.A2( u2_u15_u0_n100 ) , .ZN( u2_u15_u0_n131 ) , .A1( u2_u15_u0_n92 ) );
  NAND2_X1 u2_u15_u0_U37 (.ZN( u2_u15_u0_n108 ) , .A1( u2_u15_u0_n92 ) , .A2( u2_u15_u0_n94 ) );
  NAND2_X1 u2_u15_u0_U38 (.A2( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n114 ) , .A1( u2_u15_u0_n92 ) );
  NAND2_X1 u2_u15_u0_U39 (.A1( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n130 ) , .A2( u2_u15_u0_n94 ) );
  AOI21_X1 u2_u15_u0_U4 (.B1( u2_u15_u0_n114 ) , .ZN( u2_u15_u0_n115 ) , .B2( u2_u15_u0_n129 ) , .A( u2_u15_u0_n161 ) );
  NAND2_X1 u2_u15_u0_U40 (.A2( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n121 ) , .A1( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U41 (.ZN( u2_u15_u0_n172 ) , .A( u2_u15_u0_n88 ) );
  OAI222_X1 u2_u15_u0_U42 (.C1( u2_u15_u0_n108 ) , .A1( u2_u15_u0_n125 ) , .B2( u2_u15_u0_n128 ) , .B1( u2_u15_u0_n144 ) , .A2( u2_u15_u0_n158 ) , .C2( u2_u15_u0_n161 ) , .ZN( u2_u15_u0_n88 ) );
  NAND2_X1 u2_u15_u0_U43 (.ZN( u2_u15_u0_n112 ) , .A2( u2_u15_u0_n92 ) , .A1( u2_u15_u0_n93 ) );
  OR3_X1 u2_u15_u0_U44 (.A3( u2_u15_u0_n152 ) , .A2( u2_u15_u0_n153 ) , .A1( u2_u15_u0_n154 ) , .ZN( u2_u15_u0_n155 ) );
  AOI21_X1 u2_u15_u0_U45 (.B2( u2_u15_u0_n150 ) , .B1( u2_u15_u0_n151 ) , .ZN( u2_u15_u0_n152 ) , .A( u2_u15_u0_n158 ) );
  AOI21_X1 u2_u15_u0_U46 (.A( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n145 ) , .B1( u2_u15_u0_n146 ) , .ZN( u2_u15_u0_n154 ) );
  AOI21_X1 u2_u15_u0_U47 (.A( u2_u15_u0_n147 ) , .B2( u2_u15_u0_n148 ) , .B1( u2_u15_u0_n149 ) , .ZN( u2_u15_u0_n153 ) );
  INV_X1 u2_u15_u0_U48 (.ZN( u2_u15_u0_n171 ) , .A( u2_u15_u0_n99 ) );
  OAI211_X1 u2_u15_u0_U49 (.C2( u2_u15_u0_n140 ) , .C1( u2_u15_u0_n161 ) , .A( u2_u15_u0_n169 ) , .B( u2_u15_u0_n98 ) , .ZN( u2_u15_u0_n99 ) );
  AOI21_X1 u2_u15_u0_U5 (.B2( u2_u15_u0_n131 ) , .ZN( u2_u15_u0_n134 ) , .B1( u2_u15_u0_n151 ) , .A( u2_u15_u0_n158 ) );
  AOI211_X1 u2_u15_u0_U50 (.C1( u2_u15_u0_n118 ) , .A( u2_u15_u0_n123 ) , .B( u2_u15_u0_n96 ) , .C2( u2_u15_u0_n97 ) , .ZN( u2_u15_u0_n98 ) );
  INV_X1 u2_u15_u0_U51 (.ZN( u2_u15_u0_n169 ) , .A( u2_u15_u0_n91 ) );
  NOR2_X1 u2_u15_u0_U52 (.A2( u2_u15_X_2 ) , .ZN( u2_u15_u0_n103 ) , .A1( u2_u15_u0_n164 ) );
  NOR2_X1 u2_u15_u0_U53 (.A2( u2_u15_X_4 ) , .A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n118 ) );
  NOR2_X1 u2_u15_u0_U54 (.A2( u2_u15_X_1 ) , .A1( u2_u15_X_2 ) , .ZN( u2_u15_u0_n92 ) );
  NOR2_X1 u2_u15_u0_U55 (.A2( u2_u15_X_1 ) , .ZN( u2_u15_u0_n101 ) , .A1( u2_u15_u0_n163 ) );
  NOR2_X1 u2_u15_u0_U56 (.A2( u2_u15_X_3 ) , .A1( u2_u15_X_6 ) , .ZN( u2_u15_u0_n94 ) );
  NOR2_X1 u2_u15_u0_U57 (.A2( u2_u15_X_6 ) , .ZN( u2_u15_u0_n100 ) , .A1( u2_u15_u0_n162 ) );
  NAND2_X1 u2_u15_u0_U58 (.A2( u2_u15_X_4 ) , .A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n144 ) );
  NOR2_X1 u2_u15_u0_U59 (.A2( u2_u15_X_5 ) , .ZN( u2_u15_u0_n136 ) , .A1( u2_u15_u0_n159 ) );
  NOR2_X1 u2_u15_u0_U6 (.A1( u2_u15_u0_n108 ) , .ZN( u2_u15_u0_n123 ) , .A2( u2_u15_u0_n158 ) );
  NAND2_X1 u2_u15_u0_U60 (.A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n138 ) , .A2( u2_u15_u0_n159 ) );
  AND2_X1 u2_u15_u0_U61 (.A2( u2_u15_X_3 ) , .A1( u2_u15_X_6 ) , .ZN( u2_u15_u0_n102 ) );
  AND2_X1 u2_u15_u0_U62 (.A1( u2_u15_X_6 ) , .A2( u2_u15_u0_n162 ) , .ZN( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U63 (.A( u2_u15_X_4 ) , .ZN( u2_u15_u0_n159 ) );
  INV_X1 u2_u15_u0_U64 (.A( u2_u15_X_1 ) , .ZN( u2_u15_u0_n164 ) );
  INV_X1 u2_u15_u0_U65 (.A( u2_u15_X_2 ) , .ZN( u2_u15_u0_n163 ) );
  INV_X1 u2_u15_u0_U66 (.A( u2_u15_X_3 ) , .ZN( u2_u15_u0_n162 ) );
  INV_X1 u2_u15_u0_U67 (.A( u2_u15_u0_n126 ) , .ZN( u2_u15_u0_n168 ) );
  AOI211_X1 u2_u15_u0_U68 (.B( u2_u15_u0_n133 ) , .A( u2_u15_u0_n134 ) , .C2( u2_u15_u0_n135 ) , .C1( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n137 ) );
  OR4_X1 u2_u15_u0_U69 (.ZN( u2_out15_17 ) , .A4( u2_u15_u0_n122 ) , .A2( u2_u15_u0_n123 ) , .A1( u2_u15_u0_n124 ) , .A3( u2_u15_u0_n170 ) );
  OAI21_X1 u2_u15_u0_U7 (.B1( u2_u15_u0_n150 ) , .B2( u2_u15_u0_n158 ) , .A( u2_u15_u0_n172 ) , .ZN( u2_u15_u0_n89 ) );
  AOI21_X1 u2_u15_u0_U70 (.B2( u2_u15_u0_n107 ) , .ZN( u2_u15_u0_n124 ) , .B1( u2_u15_u0_n128 ) , .A( u2_u15_u0_n161 ) );
  INV_X1 u2_u15_u0_U71 (.A( u2_u15_u0_n111 ) , .ZN( u2_u15_u0_n170 ) );
  OR4_X1 u2_u15_u0_U72 (.ZN( u2_out15_31 ) , .A4( u2_u15_u0_n155 ) , .A2( u2_u15_u0_n156 ) , .A1( u2_u15_u0_n157 ) , .A3( u2_u15_u0_n173 ) );
  AOI21_X1 u2_u15_u0_U73 (.A( u2_u15_u0_n138 ) , .B2( u2_u15_u0_n139 ) , .B1( u2_u15_u0_n140 ) , .ZN( u2_u15_u0_n157 ) );
  AOI21_X1 u2_u15_u0_U74 (.B2( u2_u15_u0_n141 ) , .B1( u2_u15_u0_n142 ) , .ZN( u2_u15_u0_n156 ) , .A( u2_u15_u0_n161 ) );
  INV_X1 u2_u15_u0_U75 (.ZN( u2_u15_u0_n174 ) , .A( u2_u15_u0_n89 ) );
  AOI211_X1 u2_u15_u0_U76 (.B( u2_u15_u0_n104 ) , .A( u2_u15_u0_n105 ) , .ZN( u2_u15_u0_n106 ) , .C2( u2_u15_u0_n113 ) , .C1( u2_u15_u0_n160 ) );
  NOR2_X1 u2_u15_u0_U77 (.A1( u2_u15_u0_n163 ) , .A2( u2_u15_u0_n164 ) , .ZN( u2_u15_u0_n95 ) );
  OAI221_X1 u2_u15_u0_U78 (.C1( u2_u15_u0_n121 ) , .ZN( u2_u15_u0_n122 ) , .B2( u2_u15_u0_n127 ) , .A( u2_u15_u0_n143 ) , .B1( u2_u15_u0_n144 ) , .C2( u2_u15_u0_n147 ) );
  NOR2_X1 u2_u15_u0_U79 (.A1( u2_u15_u0_n120 ) , .ZN( u2_u15_u0_n143 ) , .A2( u2_u15_u0_n167 ) );
  AND2_X1 u2_u15_u0_U8 (.A1( u2_u15_u0_n114 ) , .A2( u2_u15_u0_n121 ) , .ZN( u2_u15_u0_n146 ) );
  AOI21_X1 u2_u15_u0_U80 (.B1( u2_u15_u0_n132 ) , .ZN( u2_u15_u0_n133 ) , .A( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n166 ) );
  OAI22_X1 u2_u15_u0_U81 (.ZN( u2_u15_u0_n105 ) , .A2( u2_u15_u0_n132 ) , .B1( u2_u15_u0_n146 ) , .A1( u2_u15_u0_n147 ) , .B2( u2_u15_u0_n161 ) );
  NAND2_X1 u2_u15_u0_U82 (.ZN( u2_u15_u0_n110 ) , .A2( u2_u15_u0_n132 ) , .A1( u2_u15_u0_n145 ) );
  INV_X1 u2_u15_u0_U83 (.A( u2_u15_u0_n119 ) , .ZN( u2_u15_u0_n167 ) );
  NAND2_X1 u2_u15_u0_U84 (.ZN( u2_u15_u0_n148 ) , .A1( u2_u15_u0_n93 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U85 (.A1( u2_u15_u0_n100 ) , .ZN( u2_u15_u0_n129 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U86 (.A1( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n128 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U87 (.ZN( u2_u15_u0_n142 ) , .A1( u2_u15_u0_n94 ) , .A2( u2_u15_u0_n95 ) );
  NAND3_X1 u2_u15_u0_U88 (.ZN( u2_out15_23 ) , .A3( u2_u15_u0_n137 ) , .A1( u2_u15_u0_n168 ) , .A2( u2_u15_u0_n171 ) );
  NAND3_X1 u2_u15_u0_U89 (.A3( u2_u15_u0_n127 ) , .A2( u2_u15_u0_n128 ) , .ZN( u2_u15_u0_n135 ) , .A1( u2_u15_u0_n150 ) );
  AND2_X1 u2_u15_u0_U9 (.A1( u2_u15_u0_n131 ) , .ZN( u2_u15_u0_n141 ) , .A2( u2_u15_u0_n150 ) );
  NAND3_X1 u2_u15_u0_U90 (.ZN( u2_u15_u0_n117 ) , .A3( u2_u15_u0_n132 ) , .A2( u2_u15_u0_n139 ) , .A1( u2_u15_u0_n148 ) );
  NAND3_X1 u2_u15_u0_U91 (.ZN( u2_u15_u0_n109 ) , .A2( u2_u15_u0_n114 ) , .A3( u2_u15_u0_n140 ) , .A1( u2_u15_u0_n149 ) );
  NAND3_X1 u2_u15_u0_U92 (.ZN( u2_out15_9 ) , .A3( u2_u15_u0_n106 ) , .A2( u2_u15_u0_n171 ) , .A1( u2_u15_u0_n174 ) );
  NAND3_X1 u2_u15_u0_U93 (.A2( u2_u15_u0_n128 ) , .A1( u2_u15_u0_n132 ) , .A3( u2_u15_u0_n146 ) , .ZN( u2_u15_u0_n97 ) );
  NOR2_X1 u2_u15_u1_U10 (.A1( u2_u15_u1_n112 ) , .A2( u2_u15_u1_n116 ) , .ZN( u2_u15_u1_n118 ) );
  NAND3_X1 u2_u15_u1_U100 (.ZN( u2_u15_u1_n113 ) , .A1( u2_u15_u1_n120 ) , .A3( u2_u15_u1_n133 ) , .A2( u2_u15_u1_n155 ) );
  OAI21_X1 u2_u15_u1_U11 (.ZN( u2_u15_u1_n101 ) , .B1( u2_u15_u1_n141 ) , .A( u2_u15_u1_n146 ) , .B2( u2_u15_u1_n183 ) );
  AOI21_X1 u2_u15_u1_U12 (.B2( u2_u15_u1_n155 ) , .B1( u2_u15_u1_n156 ) , .ZN( u2_u15_u1_n157 ) , .A( u2_u15_u1_n174 ) );
  NAND2_X1 u2_u15_u1_U13 (.ZN( u2_u15_u1_n140 ) , .A2( u2_u15_u1_n150 ) , .A1( u2_u15_u1_n155 ) );
  NAND2_X1 u2_u15_u1_U14 (.A1( u2_u15_u1_n131 ) , .ZN( u2_u15_u1_n147 ) , .A2( u2_u15_u1_n153 ) );
  INV_X1 u2_u15_u1_U15 (.A( u2_u15_u1_n139 ) , .ZN( u2_u15_u1_n174 ) );
  OR4_X1 u2_u15_u1_U16 (.A4( u2_u15_u1_n106 ) , .A3( u2_u15_u1_n107 ) , .ZN( u2_u15_u1_n108 ) , .A1( u2_u15_u1_n117 ) , .A2( u2_u15_u1_n184 ) );
  AOI21_X1 u2_u15_u1_U17 (.ZN( u2_u15_u1_n106 ) , .A( u2_u15_u1_n112 ) , .B1( u2_u15_u1_n154 ) , .B2( u2_u15_u1_n156 ) );
  AOI21_X1 u2_u15_u1_U18 (.ZN( u2_u15_u1_n107 ) , .B1( u2_u15_u1_n134 ) , .B2( u2_u15_u1_n149 ) , .A( u2_u15_u1_n174 ) );
  INV_X1 u2_u15_u1_U19 (.A( u2_u15_u1_n101 ) , .ZN( u2_u15_u1_n184 ) );
  INV_X1 u2_u15_u1_U20 (.A( u2_u15_u1_n112 ) , .ZN( u2_u15_u1_n171 ) );
  NAND2_X1 u2_u15_u1_U21 (.ZN( u2_u15_u1_n141 ) , .A1( u2_u15_u1_n153 ) , .A2( u2_u15_u1_n156 ) );
  AND2_X1 u2_u15_u1_U22 (.A1( u2_u15_u1_n123 ) , .ZN( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n161 ) );
  NAND2_X1 u2_u15_u1_U23 (.A2( u2_u15_u1_n115 ) , .A1( u2_u15_u1_n116 ) , .ZN( u2_u15_u1_n148 ) );
  NAND2_X1 u2_u15_u1_U24 (.A2( u2_u15_u1_n133 ) , .A1( u2_u15_u1_n135 ) , .ZN( u2_u15_u1_n159 ) );
  NAND2_X1 u2_u15_u1_U25 (.A2( u2_u15_u1_n115 ) , .A1( u2_u15_u1_n120 ) , .ZN( u2_u15_u1_n132 ) );
  INV_X1 u2_u15_u1_U26 (.A( u2_u15_u1_n154 ) , .ZN( u2_u15_u1_n178 ) );
  INV_X1 u2_u15_u1_U27 (.A( u2_u15_u1_n151 ) , .ZN( u2_u15_u1_n183 ) );
  AND2_X1 u2_u15_u1_U28 (.A1( u2_u15_u1_n129 ) , .A2( u2_u15_u1_n133 ) , .ZN( u2_u15_u1_n149 ) );
  INV_X1 u2_u15_u1_U29 (.A( u2_u15_u1_n131 ) , .ZN( u2_u15_u1_n180 ) );
  INV_X1 u2_u15_u1_U3 (.A( u2_u15_u1_n159 ) , .ZN( u2_u15_u1_n182 ) );
  OAI221_X1 u2_u15_u1_U30 (.A( u2_u15_u1_n119 ) , .C2( u2_u15_u1_n129 ) , .ZN( u2_u15_u1_n138 ) , .B2( u2_u15_u1_n152 ) , .C1( u2_u15_u1_n174 ) , .B1( u2_u15_u1_n187 ) );
  INV_X1 u2_u15_u1_U31 (.A( u2_u15_u1_n148 ) , .ZN( u2_u15_u1_n187 ) );
  AOI211_X1 u2_u15_u1_U32 (.B( u2_u15_u1_n117 ) , .A( u2_u15_u1_n118 ) , .ZN( u2_u15_u1_n119 ) , .C2( u2_u15_u1_n146 ) , .C1( u2_u15_u1_n159 ) );
  NOR2_X1 u2_u15_u1_U33 (.A1( u2_u15_u1_n168 ) , .A2( u2_u15_u1_n176 ) , .ZN( u2_u15_u1_n98 ) );
  AOI211_X1 u2_u15_u1_U34 (.B( u2_u15_u1_n162 ) , .A( u2_u15_u1_n163 ) , .C2( u2_u15_u1_n164 ) , .ZN( u2_u15_u1_n165 ) , .C1( u2_u15_u1_n171 ) );
  AOI21_X1 u2_u15_u1_U35 (.A( u2_u15_u1_n160 ) , .B2( u2_u15_u1_n161 ) , .ZN( u2_u15_u1_n162 ) , .B1( u2_u15_u1_n182 ) );
  OR2_X1 u2_u15_u1_U36 (.A2( u2_u15_u1_n157 ) , .A1( u2_u15_u1_n158 ) , .ZN( u2_u15_u1_n163 ) );
  NAND2_X1 u2_u15_u1_U37 (.A1( u2_u15_u1_n128 ) , .ZN( u2_u15_u1_n146 ) , .A2( u2_u15_u1_n160 ) );
  NAND2_X1 u2_u15_u1_U38 (.A2( u2_u15_u1_n112 ) , .ZN( u2_u15_u1_n139 ) , .A1( u2_u15_u1_n152 ) );
  NAND2_X1 u2_u15_u1_U39 (.A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n156 ) , .A2( u2_u15_u1_n99 ) );
  AOI221_X1 u2_u15_u1_U4 (.A( u2_u15_u1_n138 ) , .C2( u2_u15_u1_n139 ) , .C1( u2_u15_u1_n140 ) , .B2( u2_u15_u1_n141 ) , .ZN( u2_u15_u1_n142 ) , .B1( u2_u15_u1_n175 ) );
  AOI221_X1 u2_u15_u1_U40 (.B1( u2_u15_u1_n140 ) , .ZN( u2_u15_u1_n167 ) , .B2( u2_u15_u1_n172 ) , .C2( u2_u15_u1_n175 ) , .C1( u2_u15_u1_n178 ) , .A( u2_u15_u1_n188 ) );
  INV_X1 u2_u15_u1_U41 (.ZN( u2_u15_u1_n188 ) , .A( u2_u15_u1_n97 ) );
  AOI211_X1 u2_u15_u1_U42 (.A( u2_u15_u1_n118 ) , .C1( u2_u15_u1_n132 ) , .C2( u2_u15_u1_n139 ) , .B( u2_u15_u1_n96 ) , .ZN( u2_u15_u1_n97 ) );
  AOI21_X1 u2_u15_u1_U43 (.B2( u2_u15_u1_n121 ) , .B1( u2_u15_u1_n135 ) , .A( u2_u15_u1_n152 ) , .ZN( u2_u15_u1_n96 ) );
  NOR2_X1 u2_u15_u1_U44 (.ZN( u2_u15_u1_n117 ) , .A1( u2_u15_u1_n121 ) , .A2( u2_u15_u1_n160 ) );
  AOI21_X1 u2_u15_u1_U45 (.A( u2_u15_u1_n128 ) , .B2( u2_u15_u1_n129 ) , .ZN( u2_u15_u1_n130 ) , .B1( u2_u15_u1_n150 ) );
  OAI21_X1 u2_u15_u1_U46 (.B2( u2_u15_u1_n123 ) , .ZN( u2_u15_u1_n145 ) , .B1( u2_u15_u1_n160 ) , .A( u2_u15_u1_n185 ) );
  INV_X1 u2_u15_u1_U47 (.A( u2_u15_u1_n122 ) , .ZN( u2_u15_u1_n185 ) );
  AOI21_X1 u2_u15_u1_U48 (.B2( u2_u15_u1_n120 ) , .B1( u2_u15_u1_n121 ) , .ZN( u2_u15_u1_n122 ) , .A( u2_u15_u1_n128 ) );
  NAND2_X1 u2_u15_u1_U49 (.ZN( u2_u15_u1_n112 ) , .A1( u2_u15_u1_n169 ) , .A2( u2_u15_u1_n170 ) );
  AOI211_X1 u2_u15_u1_U5 (.ZN( u2_u15_u1_n124 ) , .A( u2_u15_u1_n138 ) , .C2( u2_u15_u1_n139 ) , .B( u2_u15_u1_n145 ) , .C1( u2_u15_u1_n147 ) );
  NAND2_X1 u2_u15_u1_U50 (.ZN( u2_u15_u1_n129 ) , .A2( u2_u15_u1_n95 ) , .A1( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U51 (.A1( u2_u15_u1_n102 ) , .ZN( u2_u15_u1_n154 ) , .A2( u2_u15_u1_n99 ) );
  NAND2_X1 u2_u15_u1_U52 (.A2( u2_u15_u1_n100 ) , .ZN( u2_u15_u1_n135 ) , .A1( u2_u15_u1_n99 ) );
  AOI21_X1 u2_u15_u1_U53 (.A( u2_u15_u1_n152 ) , .B2( u2_u15_u1_n153 ) , .B1( u2_u15_u1_n154 ) , .ZN( u2_u15_u1_n158 ) );
  INV_X1 u2_u15_u1_U54 (.A( u2_u15_u1_n160 ) , .ZN( u2_u15_u1_n175 ) );
  NAND2_X1 u2_u15_u1_U55 (.A1( u2_u15_u1_n100 ) , .ZN( u2_u15_u1_n116 ) , .A2( u2_u15_u1_n95 ) );
  NAND2_X1 u2_u15_u1_U56 (.A1( u2_u15_u1_n102 ) , .ZN( u2_u15_u1_n131 ) , .A2( u2_u15_u1_n95 ) );
  NAND2_X1 u2_u15_u1_U57 (.A2( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n121 ) , .A1( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U58 (.A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n153 ) , .A2( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U59 (.A2( u2_u15_u1_n104 ) , .A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n133 ) );
  AOI22_X1 u2_u15_u1_U6 (.B2( u2_u15_u1_n136 ) , .A2( u2_u15_u1_n137 ) , .ZN( u2_u15_u1_n143 ) , .A1( u2_u15_u1_n171 ) , .B1( u2_u15_u1_n173 ) );
  NAND2_X1 u2_u15_u1_U60 (.ZN( u2_u15_u1_n150 ) , .A2( u2_u15_u1_n98 ) , .A1( u2_u15_u1_n99 ) );
  NAND2_X1 u2_u15_u1_U61 (.A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n155 ) , .A2( u2_u15_u1_n95 ) );
  OAI21_X1 u2_u15_u1_U62 (.ZN( u2_u15_u1_n109 ) , .B1( u2_u15_u1_n129 ) , .B2( u2_u15_u1_n160 ) , .A( u2_u15_u1_n167 ) );
  NAND2_X1 u2_u15_u1_U63 (.A2( u2_u15_u1_n100 ) , .A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n120 ) );
  NAND2_X1 u2_u15_u1_U64 (.A1( u2_u15_u1_n102 ) , .A2( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n115 ) );
  NAND2_X1 u2_u15_u1_U65 (.A2( u2_u15_u1_n100 ) , .A1( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n151 ) );
  NAND2_X1 u2_u15_u1_U66 (.A2( u2_u15_u1_n103 ) , .A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n161 ) );
  INV_X1 u2_u15_u1_U67 (.A( u2_u15_u1_n152 ) , .ZN( u2_u15_u1_n173 ) );
  INV_X1 u2_u15_u1_U68 (.A( u2_u15_u1_n128 ) , .ZN( u2_u15_u1_n172 ) );
  NAND2_X1 u2_u15_u1_U69 (.A2( u2_u15_u1_n102 ) , .A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n123 ) );
  INV_X1 u2_u15_u1_U7 (.A( u2_u15_u1_n147 ) , .ZN( u2_u15_u1_n181 ) );
  NOR2_X1 u2_u15_u1_U70 (.A2( u2_u15_X_7 ) , .A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n95 ) );
  NOR2_X1 u2_u15_u1_U71 (.A1( u2_u15_X_12 ) , .A2( u2_u15_X_9 ) , .ZN( u2_u15_u1_n100 ) );
  NOR2_X1 u2_u15_u1_U72 (.A2( u2_u15_X_8 ) , .A1( u2_u15_u1_n177 ) , .ZN( u2_u15_u1_n99 ) );
  NOR2_X1 u2_u15_u1_U73 (.A2( u2_u15_X_12 ) , .ZN( u2_u15_u1_n102 ) , .A1( u2_u15_u1_n176 ) );
  NOR2_X1 u2_u15_u1_U74 (.A2( u2_u15_X_9 ) , .ZN( u2_u15_u1_n105 ) , .A1( u2_u15_u1_n168 ) );
  NAND2_X1 u2_u15_u1_U75 (.A1( u2_u15_X_10 ) , .ZN( u2_u15_u1_n160 ) , .A2( u2_u15_u1_n169 ) );
  NAND2_X1 u2_u15_u1_U76 (.A2( u2_u15_X_10 ) , .A1( u2_u15_X_11 ) , .ZN( u2_u15_u1_n152 ) );
  NAND2_X1 u2_u15_u1_U77 (.A1( u2_u15_X_11 ) , .ZN( u2_u15_u1_n128 ) , .A2( u2_u15_u1_n170 ) );
  AND2_X1 u2_u15_u1_U78 (.A2( u2_u15_X_7 ) , .A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n104 ) );
  AND2_X1 u2_u15_u1_U79 (.A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n103 ) , .A2( u2_u15_u1_n177 ) );
  AOI22_X1 u2_u15_u1_U8 (.B2( u2_u15_u1_n113 ) , .A2( u2_u15_u1_n114 ) , .ZN( u2_u15_u1_n125 ) , .A1( u2_u15_u1_n171 ) , .B1( u2_u15_u1_n173 ) );
  INV_X1 u2_u15_u1_U80 (.A( u2_u15_X_10 ) , .ZN( u2_u15_u1_n170 ) );
  INV_X1 u2_u15_u1_U81 (.A( u2_u15_X_9 ) , .ZN( u2_u15_u1_n176 ) );
  INV_X1 u2_u15_u1_U82 (.A( u2_u15_X_11 ) , .ZN( u2_u15_u1_n169 ) );
  INV_X1 u2_u15_u1_U83 (.A( u2_u15_X_12 ) , .ZN( u2_u15_u1_n168 ) );
  INV_X1 u2_u15_u1_U84 (.A( u2_u15_X_7 ) , .ZN( u2_u15_u1_n177 ) );
  NAND4_X1 u2_u15_u1_U85 (.ZN( u2_out15_18 ) , .A4( u2_u15_u1_n165 ) , .A3( u2_u15_u1_n166 ) , .A1( u2_u15_u1_n167 ) , .A2( u2_u15_u1_n186 ) );
  AOI22_X1 u2_u15_u1_U86 (.B2( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n147 ) , .A2( u2_u15_u1_n148 ) , .ZN( u2_u15_u1_n166 ) , .A1( u2_u15_u1_n172 ) );
  INV_X1 u2_u15_u1_U87 (.A( u2_u15_u1_n145 ) , .ZN( u2_u15_u1_n186 ) );
  NAND4_X1 u2_u15_u1_U88 (.ZN( u2_out15_2 ) , .A4( u2_u15_u1_n142 ) , .A3( u2_u15_u1_n143 ) , .A2( u2_u15_u1_n144 ) , .A1( u2_u15_u1_n179 ) );
  OAI21_X1 u2_u15_u1_U89 (.B2( u2_u15_u1_n132 ) , .ZN( u2_u15_u1_n144 ) , .A( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n180 ) );
  NAND2_X1 u2_u15_u1_U9 (.ZN( u2_u15_u1_n114 ) , .A1( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n156 ) );
  INV_X1 u2_u15_u1_U90 (.A( u2_u15_u1_n130 ) , .ZN( u2_u15_u1_n179 ) );
  NAND4_X1 u2_u15_u1_U91 (.ZN( u2_out15_28 ) , .A4( u2_u15_u1_n124 ) , .A3( u2_u15_u1_n125 ) , .A2( u2_u15_u1_n126 ) , .A1( u2_u15_u1_n127 ) );
  OAI21_X1 u2_u15_u1_U92 (.ZN( u2_u15_u1_n127 ) , .B2( u2_u15_u1_n139 ) , .B1( u2_u15_u1_n175 ) , .A( u2_u15_u1_n183 ) );
  OAI21_X1 u2_u15_u1_U93 (.ZN( u2_u15_u1_n126 ) , .B2( u2_u15_u1_n140 ) , .A( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n178 ) );
  OR4_X1 u2_u15_u1_U94 (.ZN( u2_out15_13 ) , .A4( u2_u15_u1_n108 ) , .A3( u2_u15_u1_n109 ) , .A2( u2_u15_u1_n110 ) , .A1( u2_u15_u1_n111 ) );
  AOI21_X1 u2_u15_u1_U95 (.ZN( u2_u15_u1_n111 ) , .A( u2_u15_u1_n128 ) , .B2( u2_u15_u1_n131 ) , .B1( u2_u15_u1_n135 ) );
  AOI21_X1 u2_u15_u1_U96 (.ZN( u2_u15_u1_n110 ) , .A( u2_u15_u1_n116 ) , .B1( u2_u15_u1_n152 ) , .B2( u2_u15_u1_n160 ) );
  NAND3_X1 u2_u15_u1_U97 (.A3( u2_u15_u1_n149 ) , .A2( u2_u15_u1_n150 ) , .A1( u2_u15_u1_n151 ) , .ZN( u2_u15_u1_n164 ) );
  NAND3_X1 u2_u15_u1_U98 (.A3( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n135 ) , .ZN( u2_u15_u1_n136 ) , .A1( u2_u15_u1_n151 ) );
  NAND3_X1 u2_u15_u1_U99 (.A1( u2_u15_u1_n133 ) , .ZN( u2_u15_u1_n137 ) , .A2( u2_u15_u1_n154 ) , .A3( u2_u15_u1_n181 ) );
  OAI22_X1 u2_u15_u2_U10 (.B1( u2_u15_u2_n151 ) , .A2( u2_u15_u2_n152 ) , .A1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n160 ) , .B2( u2_u15_u2_n168 ) );
  NAND3_X1 u2_u15_u2_U100 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n98 ) );
  NOR3_X1 u2_u15_u2_U11 (.A1( u2_u15_u2_n150 ) , .ZN( u2_u15_u2_n151 ) , .A3( u2_u15_u2_n175 ) , .A2( u2_u15_u2_n188 ) );
  AOI21_X1 u2_u15_u2_U12 (.B2( u2_u15_u2_n123 ) , .ZN( u2_u15_u2_n125 ) , .A( u2_u15_u2_n171 ) , .B1( u2_u15_u2_n184 ) );
  INV_X1 u2_u15_u2_U13 (.A( u2_u15_u2_n150 ) , .ZN( u2_u15_u2_n184 ) );
  AOI21_X1 u2_u15_u2_U14 (.ZN( u2_u15_u2_n144 ) , .B2( u2_u15_u2_n155 ) , .A( u2_u15_u2_n172 ) , .B1( u2_u15_u2_n185 ) );
  AOI21_X1 u2_u15_u2_U15 (.B2( u2_u15_u2_n143 ) , .ZN( u2_u15_u2_n145 ) , .B1( u2_u15_u2_n152 ) , .A( u2_u15_u2_n171 ) );
  INV_X1 u2_u15_u2_U16 (.A( u2_u15_u2_n156 ) , .ZN( u2_u15_u2_n171 ) );
  INV_X1 u2_u15_u2_U17 (.A( u2_u15_u2_n120 ) , .ZN( u2_u15_u2_n188 ) );
  NAND2_X1 u2_u15_u2_U18 (.A2( u2_u15_u2_n122 ) , .ZN( u2_u15_u2_n150 ) , .A1( u2_u15_u2_n152 ) );
  INV_X1 u2_u15_u2_U19 (.A( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n170 ) );
  INV_X1 u2_u15_u2_U20 (.A( u2_u15_u2_n137 ) , .ZN( u2_u15_u2_n173 ) );
  NAND2_X1 u2_u15_u2_U21 (.A1( u2_u15_u2_n132 ) , .A2( u2_u15_u2_n139 ) , .ZN( u2_u15_u2_n157 ) );
  INV_X1 u2_u15_u2_U22 (.A( u2_u15_u2_n113 ) , .ZN( u2_u15_u2_n178 ) );
  INV_X1 u2_u15_u2_U23 (.A( u2_u15_u2_n139 ) , .ZN( u2_u15_u2_n175 ) );
  INV_X1 u2_u15_u2_U24 (.A( u2_u15_u2_n155 ) , .ZN( u2_u15_u2_n181 ) );
  INV_X1 u2_u15_u2_U25 (.A( u2_u15_u2_n119 ) , .ZN( u2_u15_u2_n177 ) );
  INV_X1 u2_u15_u2_U26 (.A( u2_u15_u2_n116 ) , .ZN( u2_u15_u2_n180 ) );
  INV_X1 u2_u15_u2_U27 (.A( u2_u15_u2_n131 ) , .ZN( u2_u15_u2_n179 ) );
  INV_X1 u2_u15_u2_U28 (.A( u2_u15_u2_n154 ) , .ZN( u2_u15_u2_n176 ) );
  NAND2_X1 u2_u15_u2_U29 (.A2( u2_u15_u2_n116 ) , .A1( u2_u15_u2_n117 ) , .ZN( u2_u15_u2_n118 ) );
  NOR2_X1 u2_u15_u2_U3 (.ZN( u2_u15_u2_n121 ) , .A2( u2_u15_u2_n177 ) , .A1( u2_u15_u2_n180 ) );
  INV_X1 u2_u15_u2_U30 (.A( u2_u15_u2_n132 ) , .ZN( u2_u15_u2_n182 ) );
  INV_X1 u2_u15_u2_U31 (.A( u2_u15_u2_n158 ) , .ZN( u2_u15_u2_n183 ) );
  OAI21_X1 u2_u15_u2_U32 (.A( u2_u15_u2_n156 ) , .B1( u2_u15_u2_n157 ) , .ZN( u2_u15_u2_n158 ) , .B2( u2_u15_u2_n179 ) );
  NOR2_X1 u2_u15_u2_U33 (.ZN( u2_u15_u2_n156 ) , .A1( u2_u15_u2_n166 ) , .A2( u2_u15_u2_n169 ) );
  NOR2_X1 u2_u15_u2_U34 (.A2( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n137 ) , .A1( u2_u15_u2_n140 ) );
  NOR2_X1 u2_u15_u2_U35 (.A2( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n153 ) , .A1( u2_u15_u2_n156 ) );
  AOI211_X1 u2_u15_u2_U36 (.ZN( u2_u15_u2_n130 ) , .C1( u2_u15_u2_n138 ) , .C2( u2_u15_u2_n179 ) , .B( u2_u15_u2_n96 ) , .A( u2_u15_u2_n97 ) );
  OAI22_X1 u2_u15_u2_U37 (.B1( u2_u15_u2_n133 ) , .A2( u2_u15_u2_n137 ) , .A1( u2_u15_u2_n152 ) , .B2( u2_u15_u2_n168 ) , .ZN( u2_u15_u2_n97 ) );
  OAI221_X1 u2_u15_u2_U38 (.B1( u2_u15_u2_n113 ) , .C1( u2_u15_u2_n132 ) , .A( u2_u15_u2_n149 ) , .B2( u2_u15_u2_n171 ) , .C2( u2_u15_u2_n172 ) , .ZN( u2_u15_u2_n96 ) );
  OAI221_X1 u2_u15_u2_U39 (.A( u2_u15_u2_n115 ) , .C2( u2_u15_u2_n123 ) , .B2( u2_u15_u2_n143 ) , .B1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n163 ) , .C1( u2_u15_u2_n168 ) );
  INV_X1 u2_u15_u2_U4 (.A( u2_u15_u2_n134 ) , .ZN( u2_u15_u2_n185 ) );
  OAI21_X1 u2_u15_u2_U40 (.A( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n115 ) , .B1( u2_u15_u2_n176 ) , .B2( u2_u15_u2_n178 ) );
  OAI221_X1 u2_u15_u2_U41 (.A( u2_u15_u2_n135 ) , .B2( u2_u15_u2_n136 ) , .B1( u2_u15_u2_n137 ) , .ZN( u2_u15_u2_n162 ) , .C2( u2_u15_u2_n167 ) , .C1( u2_u15_u2_n185 ) );
  AND3_X1 u2_u15_u2_U42 (.A3( u2_u15_u2_n131 ) , .A2( u2_u15_u2_n132 ) , .A1( u2_u15_u2_n133 ) , .ZN( u2_u15_u2_n136 ) );
  AOI22_X1 u2_u15_u2_U43 (.ZN( u2_u15_u2_n135 ) , .B1( u2_u15_u2_n140 ) , .A1( u2_u15_u2_n156 ) , .B2( u2_u15_u2_n180 ) , .A2( u2_u15_u2_n188 ) );
  AOI21_X1 u2_u15_u2_U44 (.ZN( u2_u15_u2_n149 ) , .B1( u2_u15_u2_n173 ) , .B2( u2_u15_u2_n188 ) , .A( u2_u15_u2_n95 ) );
  AND3_X1 u2_u15_u2_U45 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n156 ) , .ZN( u2_u15_u2_n95 ) );
  OAI21_X1 u2_u15_u2_U46 (.A( u2_u15_u2_n141 ) , .B2( u2_u15_u2_n142 ) , .ZN( u2_u15_u2_n146 ) , .B1( u2_u15_u2_n153 ) );
  OAI21_X1 u2_u15_u2_U47 (.A( u2_u15_u2_n140 ) , .ZN( u2_u15_u2_n141 ) , .B1( u2_u15_u2_n176 ) , .B2( u2_u15_u2_n177 ) );
  NOR3_X1 u2_u15_u2_U48 (.ZN( u2_u15_u2_n142 ) , .A3( u2_u15_u2_n175 ) , .A2( u2_u15_u2_n178 ) , .A1( u2_u15_u2_n181 ) );
  OAI21_X1 u2_u15_u2_U49 (.A( u2_u15_u2_n101 ) , .B2( u2_u15_u2_n121 ) , .B1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n164 ) );
  NOR4_X1 u2_u15_u2_U5 (.A4( u2_u15_u2_n124 ) , .A3( u2_u15_u2_n125 ) , .A2( u2_u15_u2_n126 ) , .A1( u2_u15_u2_n127 ) , .ZN( u2_u15_u2_n128 ) );
  NAND2_X1 u2_u15_u2_U50 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n155 ) );
  NAND2_X1 u2_u15_u2_U51 (.A2( u2_u15_u2_n105 ) , .A1( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n143 ) );
  NAND2_X1 u2_u15_u2_U52 (.A1( u2_u15_u2_n104 ) , .A2( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n152 ) );
  NAND2_X1 u2_u15_u2_U53 (.A1( u2_u15_u2_n100 ) , .A2( u2_u15_u2_n105 ) , .ZN( u2_u15_u2_n132 ) );
  INV_X1 u2_u15_u2_U54 (.A( u2_u15_u2_n140 ) , .ZN( u2_u15_u2_n168 ) );
  INV_X1 u2_u15_u2_U55 (.A( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n167 ) );
  INV_X1 u2_u15_u2_U56 (.ZN( u2_u15_u2_n187 ) , .A( u2_u15_u2_n99 ) );
  OAI21_X1 u2_u15_u2_U57 (.B1( u2_u15_u2_n137 ) , .B2( u2_u15_u2_n143 ) , .A( u2_u15_u2_n98 ) , .ZN( u2_u15_u2_n99 ) );
  NAND2_X1 u2_u15_u2_U58 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n113 ) );
  NAND2_X1 u2_u15_u2_U59 (.A1( u2_u15_u2_n106 ) , .A2( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n131 ) );
  AOI21_X1 u2_u15_u2_U6 (.B2( u2_u15_u2_n119 ) , .ZN( u2_u15_u2_n127 ) , .A( u2_u15_u2_n137 ) , .B1( u2_u15_u2_n155 ) );
  NAND2_X1 u2_u15_u2_U60 (.A1( u2_u15_u2_n103 ) , .A2( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n139 ) );
  NAND2_X1 u2_u15_u2_U61 (.A1( u2_u15_u2_n103 ) , .A2( u2_u15_u2_n105 ) , .ZN( u2_u15_u2_n133 ) );
  NAND2_X1 u2_u15_u2_U62 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n103 ) , .ZN( u2_u15_u2_n154 ) );
  NAND2_X1 u2_u15_u2_U63 (.A2( u2_u15_u2_n103 ) , .A1( u2_u15_u2_n104 ) , .ZN( u2_u15_u2_n119 ) );
  NAND2_X1 u2_u15_u2_U64 (.A2( u2_u15_u2_n107 ) , .A1( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n123 ) );
  NAND2_X1 u2_u15_u2_U65 (.A1( u2_u15_u2_n104 ) , .A2( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n122 ) );
  INV_X1 u2_u15_u2_U66 (.A( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n172 ) );
  NAND2_X1 u2_u15_u2_U67 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n102 ) , .ZN( u2_u15_u2_n116 ) );
  NAND2_X1 u2_u15_u2_U68 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n120 ) );
  NAND2_X1 u2_u15_u2_U69 (.A2( u2_u15_u2_n105 ) , .A1( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n117 ) );
  AOI21_X1 u2_u15_u2_U7 (.ZN( u2_u15_u2_n124 ) , .B1( u2_u15_u2_n131 ) , .B2( u2_u15_u2_n143 ) , .A( u2_u15_u2_n172 ) );
  NOR2_X1 u2_u15_u2_U70 (.A2( u2_u15_X_16 ) , .ZN( u2_u15_u2_n140 ) , .A1( u2_u15_u2_n166 ) );
  NOR2_X1 u2_u15_u2_U71 (.A2( u2_u15_X_13 ) , .A1( u2_u15_X_14 ) , .ZN( u2_u15_u2_n100 ) );
  NOR2_X1 u2_u15_u2_U72 (.A2( u2_u15_X_16 ) , .A1( u2_u15_X_17 ) , .ZN( u2_u15_u2_n138 ) );
  NOR2_X1 u2_u15_u2_U73 (.A2( u2_u15_X_15 ) , .A1( u2_u15_X_18 ) , .ZN( u2_u15_u2_n104 ) );
  NOR2_X1 u2_u15_u2_U74 (.A2( u2_u15_X_14 ) , .ZN( u2_u15_u2_n103 ) , .A1( u2_u15_u2_n174 ) );
  NOR2_X1 u2_u15_u2_U75 (.A2( u2_u15_X_15 ) , .ZN( u2_u15_u2_n102 ) , .A1( u2_u15_u2_n165 ) );
  NOR2_X1 u2_u15_u2_U76 (.A2( u2_u15_X_17 ) , .ZN( u2_u15_u2_n114 ) , .A1( u2_u15_u2_n169 ) );
  AND2_X1 u2_u15_u2_U77 (.A1( u2_u15_X_15 ) , .ZN( u2_u15_u2_n105 ) , .A2( u2_u15_u2_n165 ) );
  AND2_X1 u2_u15_u2_U78 (.A2( u2_u15_X_15 ) , .A1( u2_u15_X_18 ) , .ZN( u2_u15_u2_n107 ) );
  AND2_X1 u2_u15_u2_U79 (.A1( u2_u15_X_14 ) , .ZN( u2_u15_u2_n106 ) , .A2( u2_u15_u2_n174 ) );
  AOI21_X1 u2_u15_u2_U8 (.B2( u2_u15_u2_n120 ) , .B1( u2_u15_u2_n121 ) , .ZN( u2_u15_u2_n126 ) , .A( u2_u15_u2_n167 ) );
  AND2_X1 u2_u15_u2_U80 (.A1( u2_u15_X_13 ) , .A2( u2_u15_X_14 ) , .ZN( u2_u15_u2_n108 ) );
  INV_X1 u2_u15_u2_U81 (.A( u2_u15_X_16 ) , .ZN( u2_u15_u2_n169 ) );
  INV_X1 u2_u15_u2_U82 (.A( u2_u15_X_17 ) , .ZN( u2_u15_u2_n166 ) );
  INV_X1 u2_u15_u2_U83 (.A( u2_u15_X_13 ) , .ZN( u2_u15_u2_n174 ) );
  INV_X1 u2_u15_u2_U84 (.A( u2_u15_X_18 ) , .ZN( u2_u15_u2_n165 ) );
  NAND4_X1 u2_u15_u2_U85 (.ZN( u2_out15_30 ) , .A4( u2_u15_u2_n147 ) , .A3( u2_u15_u2_n148 ) , .A2( u2_u15_u2_n149 ) , .A1( u2_u15_u2_n187 ) );
  NOR3_X1 u2_u15_u2_U86 (.A3( u2_u15_u2_n144 ) , .A2( u2_u15_u2_n145 ) , .A1( u2_u15_u2_n146 ) , .ZN( u2_u15_u2_n147 ) );
  AOI21_X1 u2_u15_u2_U87 (.B2( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n148 ) , .A( u2_u15_u2_n162 ) , .B1( u2_u15_u2_n182 ) );
  NAND4_X1 u2_u15_u2_U88 (.ZN( u2_out15_24 ) , .A4( u2_u15_u2_n111 ) , .A3( u2_u15_u2_n112 ) , .A1( u2_u15_u2_n130 ) , .A2( u2_u15_u2_n187 ) );
  AOI221_X1 u2_u15_u2_U89 (.A( u2_u15_u2_n109 ) , .B1( u2_u15_u2_n110 ) , .ZN( u2_u15_u2_n111 ) , .C1( u2_u15_u2_n134 ) , .C2( u2_u15_u2_n170 ) , .B2( u2_u15_u2_n173 ) );
  OAI22_X1 u2_u15_u2_U9 (.ZN( u2_u15_u2_n109 ) , .A2( u2_u15_u2_n113 ) , .B2( u2_u15_u2_n133 ) , .B1( u2_u15_u2_n167 ) , .A1( u2_u15_u2_n168 ) );
  AOI21_X1 u2_u15_u2_U90 (.ZN( u2_u15_u2_n112 ) , .B2( u2_u15_u2_n156 ) , .A( u2_u15_u2_n164 ) , .B1( u2_u15_u2_n181 ) );
  NAND4_X1 u2_u15_u2_U91 (.ZN( u2_out15_16 ) , .A4( u2_u15_u2_n128 ) , .A3( u2_u15_u2_n129 ) , .A1( u2_u15_u2_n130 ) , .A2( u2_u15_u2_n186 ) );
  AOI22_X1 u2_u15_u2_U92 (.A2( u2_u15_u2_n118 ) , .ZN( u2_u15_u2_n129 ) , .A1( u2_u15_u2_n140 ) , .B1( u2_u15_u2_n157 ) , .B2( u2_u15_u2_n170 ) );
  INV_X1 u2_u15_u2_U93 (.A( u2_u15_u2_n163 ) , .ZN( u2_u15_u2_n186 ) );
  OR4_X1 u2_u15_u2_U94 (.ZN( u2_out15_6 ) , .A4( u2_u15_u2_n161 ) , .A3( u2_u15_u2_n162 ) , .A2( u2_u15_u2_n163 ) , .A1( u2_u15_u2_n164 ) );
  OR3_X1 u2_u15_u2_U95 (.A2( u2_u15_u2_n159 ) , .A1( u2_u15_u2_n160 ) , .ZN( u2_u15_u2_n161 ) , .A3( u2_u15_u2_n183 ) );
  AOI21_X1 u2_u15_u2_U96 (.B2( u2_u15_u2_n154 ) , .B1( u2_u15_u2_n155 ) , .ZN( u2_u15_u2_n159 ) , .A( u2_u15_u2_n167 ) );
  NAND3_X1 u2_u15_u2_U97 (.A2( u2_u15_u2_n117 ) , .A1( u2_u15_u2_n122 ) , .A3( u2_u15_u2_n123 ) , .ZN( u2_u15_u2_n134 ) );
  NAND3_X1 u2_u15_u2_U98 (.ZN( u2_u15_u2_n110 ) , .A2( u2_u15_u2_n131 ) , .A3( u2_u15_u2_n139 ) , .A1( u2_u15_u2_n154 ) );
  NAND3_X1 u2_u15_u2_U99 (.A2( u2_u15_u2_n100 ) , .ZN( u2_u15_u2_n101 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n114 ) );
  OAI22_X1 u2_u15_u3_U10 (.B1( u2_u15_u3_n113 ) , .A2( u2_u15_u3_n135 ) , .A1( u2_u15_u3_n150 ) , .B2( u2_u15_u3_n164 ) , .ZN( u2_u15_u3_n98 ) );
  OAI211_X1 u2_u15_u3_U11 (.B( u2_u15_u3_n106 ) , .ZN( u2_u15_u3_n119 ) , .C2( u2_u15_u3_n128 ) , .C1( u2_u15_u3_n167 ) , .A( u2_u15_u3_n181 ) );
  AOI221_X1 u2_u15_u3_U12 (.C1( u2_u15_u3_n105 ) , .ZN( u2_u15_u3_n106 ) , .A( u2_u15_u3_n131 ) , .B2( u2_u15_u3_n132 ) , .C2( u2_u15_u3_n133 ) , .B1( u2_u15_u3_n169 ) );
  INV_X1 u2_u15_u3_U13 (.ZN( u2_u15_u3_n181 ) , .A( u2_u15_u3_n98 ) );
  NAND2_X1 u2_u15_u3_U14 (.ZN( u2_u15_u3_n105 ) , .A2( u2_u15_u3_n130 ) , .A1( u2_u15_u3_n155 ) );
  AOI22_X1 u2_u15_u3_U15 (.B1( u2_u15_u3_n115 ) , .A2( u2_u15_u3_n116 ) , .ZN( u2_u15_u3_n123 ) , .B2( u2_u15_u3_n133 ) , .A1( u2_u15_u3_n169 ) );
  NAND2_X1 u2_u15_u3_U16 (.ZN( u2_u15_u3_n116 ) , .A2( u2_u15_u3_n151 ) , .A1( u2_u15_u3_n182 ) );
  NOR2_X1 u2_u15_u3_U17 (.ZN( u2_u15_u3_n126 ) , .A2( u2_u15_u3_n150 ) , .A1( u2_u15_u3_n164 ) );
  AOI21_X1 u2_u15_u3_U18 (.ZN( u2_u15_u3_n112 ) , .B2( u2_u15_u3_n146 ) , .B1( u2_u15_u3_n155 ) , .A( u2_u15_u3_n167 ) );
  NAND2_X1 u2_u15_u3_U19 (.A1( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n142 ) , .A2( u2_u15_u3_n164 ) );
  NAND2_X1 u2_u15_u3_U20 (.ZN( u2_u15_u3_n132 ) , .A2( u2_u15_u3_n152 ) , .A1( u2_u15_u3_n156 ) );
  AND2_X1 u2_u15_u3_U21 (.A2( u2_u15_u3_n113 ) , .A1( u2_u15_u3_n114 ) , .ZN( u2_u15_u3_n151 ) );
  INV_X1 u2_u15_u3_U22 (.A( u2_u15_u3_n133 ) , .ZN( u2_u15_u3_n165 ) );
  INV_X1 u2_u15_u3_U23 (.A( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n170 ) );
  NAND2_X1 u2_u15_u3_U24 (.A1( u2_u15_u3_n107 ) , .A2( u2_u15_u3_n108 ) , .ZN( u2_u15_u3_n140 ) );
  NAND2_X1 u2_u15_u3_U25 (.ZN( u2_u15_u3_n117 ) , .A1( u2_u15_u3_n124 ) , .A2( u2_u15_u3_n148 ) );
  NAND2_X1 u2_u15_u3_U26 (.ZN( u2_u15_u3_n143 ) , .A1( u2_u15_u3_n165 ) , .A2( u2_u15_u3_n167 ) );
  INV_X1 u2_u15_u3_U27 (.A( u2_u15_u3_n130 ) , .ZN( u2_u15_u3_n177 ) );
  INV_X1 u2_u15_u3_U28 (.A( u2_u15_u3_n128 ) , .ZN( u2_u15_u3_n176 ) );
  INV_X1 u2_u15_u3_U29 (.A( u2_u15_u3_n155 ) , .ZN( u2_u15_u3_n174 ) );
  INV_X1 u2_u15_u3_U3 (.A( u2_u15_u3_n129 ) , .ZN( u2_u15_u3_n183 ) );
  INV_X1 u2_u15_u3_U30 (.A( u2_u15_u3_n139 ) , .ZN( u2_u15_u3_n185 ) );
  NOR2_X1 u2_u15_u3_U31 (.ZN( u2_u15_u3_n135 ) , .A2( u2_u15_u3_n141 ) , .A1( u2_u15_u3_n169 ) );
  OAI222_X1 u2_u15_u3_U32 (.C2( u2_u15_u3_n107 ) , .A2( u2_u15_u3_n108 ) , .B1( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n138 ) , .B2( u2_u15_u3_n146 ) , .C1( u2_u15_u3_n154 ) , .A1( u2_u15_u3_n164 ) );
  NOR4_X1 u2_u15_u3_U33 (.A4( u2_u15_u3_n157 ) , .A3( u2_u15_u3_n158 ) , .A2( u2_u15_u3_n159 ) , .A1( u2_u15_u3_n160 ) , .ZN( u2_u15_u3_n161 ) );
  AOI21_X1 u2_u15_u3_U34 (.B2( u2_u15_u3_n152 ) , .B1( u2_u15_u3_n153 ) , .ZN( u2_u15_u3_n158 ) , .A( u2_u15_u3_n164 ) );
  AOI21_X1 u2_u15_u3_U35 (.A( u2_u15_u3_n154 ) , .B2( u2_u15_u3_n155 ) , .B1( u2_u15_u3_n156 ) , .ZN( u2_u15_u3_n157 ) );
  AOI21_X1 u2_u15_u3_U36 (.A( u2_u15_u3_n149 ) , .B2( u2_u15_u3_n150 ) , .B1( u2_u15_u3_n151 ) , .ZN( u2_u15_u3_n159 ) );
  AOI211_X1 u2_u15_u3_U37 (.ZN( u2_u15_u3_n109 ) , .A( u2_u15_u3_n119 ) , .C2( u2_u15_u3_n129 ) , .B( u2_u15_u3_n138 ) , .C1( u2_u15_u3_n141 ) );
  AOI211_X1 u2_u15_u3_U38 (.B( u2_u15_u3_n119 ) , .A( u2_u15_u3_n120 ) , .C2( u2_u15_u3_n121 ) , .ZN( u2_u15_u3_n122 ) , .C1( u2_u15_u3_n179 ) );
  INV_X1 u2_u15_u3_U39 (.A( u2_u15_u3_n156 ) , .ZN( u2_u15_u3_n179 ) );
  INV_X1 u2_u15_u3_U4 (.A( u2_u15_u3_n140 ) , .ZN( u2_u15_u3_n182 ) );
  OAI22_X1 u2_u15_u3_U40 (.B1( u2_u15_u3_n118 ) , .ZN( u2_u15_u3_n120 ) , .A1( u2_u15_u3_n135 ) , .B2( u2_u15_u3_n154 ) , .A2( u2_u15_u3_n178 ) );
  AND3_X1 u2_u15_u3_U41 (.ZN( u2_u15_u3_n118 ) , .A2( u2_u15_u3_n124 ) , .A1( u2_u15_u3_n144 ) , .A3( u2_u15_u3_n152 ) );
  INV_X1 u2_u15_u3_U42 (.A( u2_u15_u3_n121 ) , .ZN( u2_u15_u3_n164 ) );
  NAND2_X1 u2_u15_u3_U43 (.ZN( u2_u15_u3_n133 ) , .A1( u2_u15_u3_n154 ) , .A2( u2_u15_u3_n164 ) );
  OAI211_X1 u2_u15_u3_U44 (.B( u2_u15_u3_n127 ) , .ZN( u2_u15_u3_n139 ) , .C1( u2_u15_u3_n150 ) , .C2( u2_u15_u3_n154 ) , .A( u2_u15_u3_n184 ) );
  INV_X1 u2_u15_u3_U45 (.A( u2_u15_u3_n125 ) , .ZN( u2_u15_u3_n184 ) );
  AOI221_X1 u2_u15_u3_U46 (.A( u2_u15_u3_n126 ) , .ZN( u2_u15_u3_n127 ) , .C2( u2_u15_u3_n132 ) , .C1( u2_u15_u3_n169 ) , .B2( u2_u15_u3_n170 ) , .B1( u2_u15_u3_n174 ) );
  OAI22_X1 u2_u15_u3_U47 (.A1( u2_u15_u3_n124 ) , .ZN( u2_u15_u3_n125 ) , .B2( u2_u15_u3_n145 ) , .A2( u2_u15_u3_n165 ) , .B1( u2_u15_u3_n167 ) );
  NOR2_X1 u2_u15_u3_U48 (.A1( u2_u15_u3_n113 ) , .ZN( u2_u15_u3_n131 ) , .A2( u2_u15_u3_n154 ) );
  NAND2_X1 u2_u15_u3_U49 (.A1( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n150 ) , .A2( u2_u15_u3_n99 ) );
  INV_X1 u2_u15_u3_U5 (.A( u2_u15_u3_n117 ) , .ZN( u2_u15_u3_n178 ) );
  NAND2_X1 u2_u15_u3_U50 (.A2( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n155 ) , .A1( u2_u15_u3_n97 ) );
  INV_X1 u2_u15_u3_U51 (.A( u2_u15_u3_n141 ) , .ZN( u2_u15_u3_n167 ) );
  AOI21_X1 u2_u15_u3_U52 (.B2( u2_u15_u3_n114 ) , .B1( u2_u15_u3_n146 ) , .A( u2_u15_u3_n154 ) , .ZN( u2_u15_u3_n94 ) );
  AOI21_X1 u2_u15_u3_U53 (.ZN( u2_u15_u3_n110 ) , .B2( u2_u15_u3_n142 ) , .B1( u2_u15_u3_n186 ) , .A( u2_u15_u3_n95 ) );
  INV_X1 u2_u15_u3_U54 (.A( u2_u15_u3_n145 ) , .ZN( u2_u15_u3_n186 ) );
  AOI21_X1 u2_u15_u3_U55 (.B1( u2_u15_u3_n124 ) , .A( u2_u15_u3_n149 ) , .B2( u2_u15_u3_n155 ) , .ZN( u2_u15_u3_n95 ) );
  INV_X1 u2_u15_u3_U56 (.A( u2_u15_u3_n149 ) , .ZN( u2_u15_u3_n169 ) );
  NAND2_X1 u2_u15_u3_U57 (.ZN( u2_u15_u3_n124 ) , .A1( u2_u15_u3_n96 ) , .A2( u2_u15_u3_n97 ) );
  NAND2_X1 u2_u15_u3_U58 (.A2( u2_u15_u3_n100 ) , .ZN( u2_u15_u3_n146 ) , .A1( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U59 (.A1( u2_u15_u3_n101 ) , .ZN( u2_u15_u3_n145 ) , .A2( u2_u15_u3_n99 ) );
  AOI221_X1 u2_u15_u3_U6 (.A( u2_u15_u3_n131 ) , .C2( u2_u15_u3_n132 ) , .C1( u2_u15_u3_n133 ) , .ZN( u2_u15_u3_n134 ) , .B1( u2_u15_u3_n143 ) , .B2( u2_u15_u3_n177 ) );
  NAND2_X1 u2_u15_u3_U60 (.A1( u2_u15_u3_n100 ) , .ZN( u2_u15_u3_n156 ) , .A2( u2_u15_u3_n99 ) );
  NAND2_X1 u2_u15_u3_U61 (.A2( u2_u15_u3_n101 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n148 ) );
  NAND2_X1 u2_u15_u3_U62 (.A1( u2_u15_u3_n100 ) , .A2( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n128 ) );
  NAND2_X1 u2_u15_u3_U63 (.A2( u2_u15_u3_n101 ) , .A1( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n152 ) );
  NAND2_X1 u2_u15_u3_U64 (.A2( u2_u15_u3_n101 ) , .ZN( u2_u15_u3_n114 ) , .A1( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U65 (.ZN( u2_u15_u3_n107 ) , .A1( u2_u15_u3_n97 ) , .A2( u2_u15_u3_n99 ) );
  NAND2_X1 u2_u15_u3_U66 (.A2( u2_u15_u3_n100 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n113 ) );
  NAND2_X1 u2_u15_u3_U67 (.A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n153 ) , .A2( u2_u15_u3_n97 ) );
  NAND2_X1 u2_u15_u3_U68 (.A2( u2_u15_u3_n103 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n130 ) );
  NAND2_X1 u2_u15_u3_U69 (.A2( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n144 ) , .A1( u2_u15_u3_n96 ) );
  OAI22_X1 u2_u15_u3_U7 (.B2( u2_u15_u3_n147 ) , .A2( u2_u15_u3_n148 ) , .ZN( u2_u15_u3_n160 ) , .B1( u2_u15_u3_n165 ) , .A1( u2_u15_u3_n168 ) );
  NAND2_X1 u2_u15_u3_U70 (.A1( u2_u15_u3_n102 ) , .A2( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n108 ) );
  NOR2_X1 u2_u15_u3_U71 (.A2( u2_u15_X_19 ) , .A1( u2_u15_X_20 ) , .ZN( u2_u15_u3_n99 ) );
  NOR2_X1 u2_u15_u3_U72 (.A2( u2_u15_X_21 ) , .A1( u2_u15_X_24 ) , .ZN( u2_u15_u3_n103 ) );
  NOR2_X1 u2_u15_u3_U73 (.A2( u2_u15_X_24 ) , .A1( u2_u15_u3_n171 ) , .ZN( u2_u15_u3_n97 ) );
  NOR2_X1 u2_u15_u3_U74 (.A2( u2_u15_X_23 ) , .ZN( u2_u15_u3_n141 ) , .A1( u2_u15_u3_n166 ) );
  NOR2_X1 u2_u15_u3_U75 (.A2( u2_u15_X_19 ) , .A1( u2_u15_u3_n172 ) , .ZN( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U76 (.A1( u2_u15_X_22 ) , .A2( u2_u15_X_23 ) , .ZN( u2_u15_u3_n154 ) );
  NAND2_X1 u2_u15_u3_U77 (.A1( u2_u15_X_23 ) , .ZN( u2_u15_u3_n149 ) , .A2( u2_u15_u3_n166 ) );
  NOR2_X1 u2_u15_u3_U78 (.A2( u2_u15_X_22 ) , .A1( u2_u15_X_23 ) , .ZN( u2_u15_u3_n121 ) );
  AND2_X1 u2_u15_u3_U79 (.A1( u2_u15_X_24 ) , .ZN( u2_u15_u3_n101 ) , .A2( u2_u15_u3_n171 ) );
  AND3_X1 u2_u15_u3_U8 (.A3( u2_u15_u3_n144 ) , .A2( u2_u15_u3_n145 ) , .A1( u2_u15_u3_n146 ) , .ZN( u2_u15_u3_n147 ) );
  AND2_X1 u2_u15_u3_U80 (.A1( u2_u15_X_19 ) , .ZN( u2_u15_u3_n102 ) , .A2( u2_u15_u3_n172 ) );
  AND2_X1 u2_u15_u3_U81 (.A1( u2_u15_X_21 ) , .A2( u2_u15_X_24 ) , .ZN( u2_u15_u3_n100 ) );
  AND2_X1 u2_u15_u3_U82 (.A2( u2_u15_X_19 ) , .A1( u2_u15_X_20 ) , .ZN( u2_u15_u3_n104 ) );
  INV_X1 u2_u15_u3_U83 (.A( u2_u15_X_22 ) , .ZN( u2_u15_u3_n166 ) );
  INV_X1 u2_u15_u3_U84 (.A( u2_u15_X_21 ) , .ZN( u2_u15_u3_n171 ) );
  INV_X1 u2_u15_u3_U85 (.A( u2_u15_X_20 ) , .ZN( u2_u15_u3_n172 ) );
  OR4_X1 u2_u15_u3_U86 (.ZN( u2_out15_10 ) , .A4( u2_u15_u3_n136 ) , .A3( u2_u15_u3_n137 ) , .A1( u2_u15_u3_n138 ) , .A2( u2_u15_u3_n139 ) );
  OAI222_X1 u2_u15_u3_U87 (.C1( u2_u15_u3_n128 ) , .ZN( u2_u15_u3_n137 ) , .B1( u2_u15_u3_n148 ) , .A2( u2_u15_u3_n150 ) , .B2( u2_u15_u3_n154 ) , .C2( u2_u15_u3_n164 ) , .A1( u2_u15_u3_n167 ) );
  OAI221_X1 u2_u15_u3_U88 (.A( u2_u15_u3_n134 ) , .B2( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n136 ) , .C1( u2_u15_u3_n149 ) , .B1( u2_u15_u3_n151 ) , .C2( u2_u15_u3_n183 ) );
  NAND4_X1 u2_u15_u3_U89 (.ZN( u2_out15_1 ) , .A4( u2_u15_u3_n161 ) , .A3( u2_u15_u3_n162 ) , .A2( u2_u15_u3_n163 ) , .A1( u2_u15_u3_n185 ) );
  INV_X1 u2_u15_u3_U9 (.A( u2_u15_u3_n143 ) , .ZN( u2_u15_u3_n168 ) );
  NAND2_X1 u2_u15_u3_U90 (.ZN( u2_u15_u3_n163 ) , .A2( u2_u15_u3_n170 ) , .A1( u2_u15_u3_n176 ) );
  AOI22_X1 u2_u15_u3_U91 (.B2( u2_u15_u3_n140 ) , .B1( u2_u15_u3_n141 ) , .A2( u2_u15_u3_n142 ) , .ZN( u2_u15_u3_n162 ) , .A1( u2_u15_u3_n177 ) );
  NAND4_X1 u2_u15_u3_U92 (.ZN( u2_out15_26 ) , .A4( u2_u15_u3_n109 ) , .A3( u2_u15_u3_n110 ) , .A2( u2_u15_u3_n111 ) , .A1( u2_u15_u3_n173 ) );
  INV_X1 u2_u15_u3_U93 (.ZN( u2_u15_u3_n173 ) , .A( u2_u15_u3_n94 ) );
  OAI21_X1 u2_u15_u3_U94 (.ZN( u2_u15_u3_n111 ) , .B2( u2_u15_u3_n117 ) , .A( u2_u15_u3_n133 ) , .B1( u2_u15_u3_n176 ) );
  NAND4_X1 u2_u15_u3_U95 (.ZN( u2_out15_20 ) , .A4( u2_u15_u3_n122 ) , .A3( u2_u15_u3_n123 ) , .A1( u2_u15_u3_n175 ) , .A2( u2_u15_u3_n180 ) );
  INV_X1 u2_u15_u3_U96 (.A( u2_u15_u3_n126 ) , .ZN( u2_u15_u3_n180 ) );
  INV_X1 u2_u15_u3_U97 (.A( u2_u15_u3_n112 ) , .ZN( u2_u15_u3_n175 ) );
  NAND3_X1 u2_u15_u3_U98 (.A1( u2_u15_u3_n114 ) , .ZN( u2_u15_u3_n115 ) , .A2( u2_u15_u3_n145 ) , .A3( u2_u15_u3_n153 ) );
  NAND3_X1 u2_u15_u3_U99 (.ZN( u2_u15_u3_n129 ) , .A2( u2_u15_u3_n144 ) , .A1( u2_u15_u3_n153 ) , .A3( u2_u15_u3_n182 ) );
  OAI22_X1 u2_u15_u4_U10 (.B2( u2_u15_u4_n135 ) , .ZN( u2_u15_u4_n137 ) , .B1( u2_u15_u4_n153 ) , .A1( u2_u15_u4_n155 ) , .A2( u2_u15_u4_n171 ) );
  AND3_X1 u2_u15_u4_U11 (.A2( u2_u15_u4_n134 ) , .ZN( u2_u15_u4_n135 ) , .A3( u2_u15_u4_n145 ) , .A1( u2_u15_u4_n157 ) );
  OR3_X1 u2_u15_u4_U12 (.A3( u2_u15_u4_n114 ) , .A2( u2_u15_u4_n115 ) , .A1( u2_u15_u4_n116 ) , .ZN( u2_u15_u4_n136 ) );
  AOI21_X1 u2_u15_u4_U13 (.A( u2_u15_u4_n113 ) , .ZN( u2_u15_u4_n116 ) , .B2( u2_u15_u4_n173 ) , .B1( u2_u15_u4_n174 ) );
  AOI21_X1 u2_u15_u4_U14 (.ZN( u2_u15_u4_n115 ) , .B2( u2_u15_u4_n145 ) , .B1( u2_u15_u4_n146 ) , .A( u2_u15_u4_n156 ) );
  OAI22_X1 u2_u15_u4_U15 (.ZN( u2_u15_u4_n114 ) , .A2( u2_u15_u4_n121 ) , .B1( u2_u15_u4_n160 ) , .B2( u2_u15_u4_n170 ) , .A1( u2_u15_u4_n171 ) );
  NAND2_X1 u2_u15_u4_U16 (.ZN( u2_u15_u4_n132 ) , .A2( u2_u15_u4_n170 ) , .A1( u2_u15_u4_n173 ) );
  AOI21_X1 u2_u15_u4_U17 (.B2( u2_u15_u4_n160 ) , .B1( u2_u15_u4_n161 ) , .ZN( u2_u15_u4_n162 ) , .A( u2_u15_u4_n170 ) );
  AOI21_X1 u2_u15_u4_U18 (.ZN( u2_u15_u4_n107 ) , .B2( u2_u15_u4_n143 ) , .A( u2_u15_u4_n174 ) , .B1( u2_u15_u4_n184 ) );
  AOI21_X1 u2_u15_u4_U19 (.B2( u2_u15_u4_n158 ) , .B1( u2_u15_u4_n159 ) , .ZN( u2_u15_u4_n163 ) , .A( u2_u15_u4_n174 ) );
  AOI21_X1 u2_u15_u4_U20 (.A( u2_u15_u4_n153 ) , .B2( u2_u15_u4_n154 ) , .B1( u2_u15_u4_n155 ) , .ZN( u2_u15_u4_n165 ) );
  AOI21_X1 u2_u15_u4_U21 (.A( u2_u15_u4_n156 ) , .B2( u2_u15_u4_n157 ) , .ZN( u2_u15_u4_n164 ) , .B1( u2_u15_u4_n184 ) );
  INV_X1 u2_u15_u4_U22 (.A( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n170 ) );
  AND2_X1 u2_u15_u4_U23 (.A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n155 ) , .A1( u2_u15_u4_n160 ) );
  INV_X1 u2_u15_u4_U24 (.A( u2_u15_u4_n156 ) , .ZN( u2_u15_u4_n175 ) );
  NAND2_X1 u2_u15_u4_U25 (.A2( u2_u15_u4_n118 ) , .ZN( u2_u15_u4_n131 ) , .A1( u2_u15_u4_n147 ) );
  NAND2_X1 u2_u15_u4_U26 (.A1( u2_u15_u4_n119 ) , .A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n130 ) );
  NAND2_X1 u2_u15_u4_U27 (.ZN( u2_u15_u4_n117 ) , .A2( u2_u15_u4_n118 ) , .A1( u2_u15_u4_n148 ) );
  NAND2_X1 u2_u15_u4_U28 (.ZN( u2_u15_u4_n129 ) , .A1( u2_u15_u4_n134 ) , .A2( u2_u15_u4_n148 ) );
  AND3_X1 u2_u15_u4_U29 (.A1( u2_u15_u4_n119 ) , .A2( u2_u15_u4_n143 ) , .A3( u2_u15_u4_n154 ) , .ZN( u2_u15_u4_n161 ) );
  NOR2_X1 u2_u15_u4_U3 (.ZN( u2_u15_u4_n121 ) , .A1( u2_u15_u4_n181 ) , .A2( u2_u15_u4_n182 ) );
  AND2_X1 u2_u15_u4_U30 (.A1( u2_u15_u4_n145 ) , .A2( u2_u15_u4_n147 ) , .ZN( u2_u15_u4_n159 ) );
  INV_X1 u2_u15_u4_U31 (.A( u2_u15_u4_n158 ) , .ZN( u2_u15_u4_n182 ) );
  INV_X1 u2_u15_u4_U32 (.ZN( u2_u15_u4_n181 ) , .A( u2_u15_u4_n96 ) );
  INV_X1 u2_u15_u4_U33 (.A( u2_u15_u4_n144 ) , .ZN( u2_u15_u4_n179 ) );
  INV_X1 u2_u15_u4_U34 (.A( u2_u15_u4_n157 ) , .ZN( u2_u15_u4_n178 ) );
  NAND2_X1 u2_u15_u4_U35 (.A2( u2_u15_u4_n154 ) , .A1( u2_u15_u4_n96 ) , .ZN( u2_u15_u4_n97 ) );
  INV_X1 u2_u15_u4_U36 (.ZN( u2_u15_u4_n186 ) , .A( u2_u15_u4_n95 ) );
  OAI221_X1 u2_u15_u4_U37 (.C1( u2_u15_u4_n134 ) , .B1( u2_u15_u4_n158 ) , .B2( u2_u15_u4_n171 ) , .C2( u2_u15_u4_n173 ) , .A( u2_u15_u4_n94 ) , .ZN( u2_u15_u4_n95 ) );
  AOI222_X1 u2_u15_u4_U38 (.B2( u2_u15_u4_n132 ) , .A1( u2_u15_u4_n138 ) , .C2( u2_u15_u4_n175 ) , .A2( u2_u15_u4_n179 ) , .C1( u2_u15_u4_n181 ) , .B1( u2_u15_u4_n185 ) , .ZN( u2_u15_u4_n94 ) );
  INV_X1 u2_u15_u4_U39 (.A( u2_u15_u4_n113 ) , .ZN( u2_u15_u4_n185 ) );
  INV_X1 u2_u15_u4_U4 (.A( u2_u15_u4_n117 ) , .ZN( u2_u15_u4_n184 ) );
  INV_X1 u2_u15_u4_U40 (.A( u2_u15_u4_n143 ) , .ZN( u2_u15_u4_n183 ) );
  NOR2_X1 u2_u15_u4_U41 (.ZN( u2_u15_u4_n138 ) , .A1( u2_u15_u4_n168 ) , .A2( u2_u15_u4_n169 ) );
  NOR2_X1 u2_u15_u4_U42 (.A1( u2_u15_u4_n150 ) , .A2( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n153 ) );
  NOR2_X1 u2_u15_u4_U43 (.A2( u2_u15_u4_n128 ) , .A1( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n156 ) );
  AOI22_X1 u2_u15_u4_U44 (.B2( u2_u15_u4_n122 ) , .A1( u2_u15_u4_n123 ) , .ZN( u2_u15_u4_n124 ) , .B1( u2_u15_u4_n128 ) , .A2( u2_u15_u4_n172 ) );
  NAND2_X1 u2_u15_u4_U45 (.A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n123 ) , .A1( u2_u15_u4_n161 ) );
  INV_X1 u2_u15_u4_U46 (.A( u2_u15_u4_n153 ) , .ZN( u2_u15_u4_n172 ) );
  AOI22_X1 u2_u15_u4_U47 (.B2( u2_u15_u4_n132 ) , .A2( u2_u15_u4_n133 ) , .ZN( u2_u15_u4_n140 ) , .A1( u2_u15_u4_n150 ) , .B1( u2_u15_u4_n179 ) );
  NAND2_X1 u2_u15_u4_U48 (.ZN( u2_u15_u4_n133 ) , .A2( u2_u15_u4_n146 ) , .A1( u2_u15_u4_n154 ) );
  NAND2_X1 u2_u15_u4_U49 (.A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n154 ) , .A2( u2_u15_u4_n98 ) );
  NOR4_X1 u2_u15_u4_U5 (.A4( u2_u15_u4_n106 ) , .A3( u2_u15_u4_n107 ) , .A2( u2_u15_u4_n108 ) , .A1( u2_u15_u4_n109 ) , .ZN( u2_u15_u4_n110 ) );
  NAND2_X1 u2_u15_u4_U50 (.A1( u2_u15_u4_n101 ) , .ZN( u2_u15_u4_n158 ) , .A2( u2_u15_u4_n99 ) );
  AOI21_X1 u2_u15_u4_U51 (.ZN( u2_u15_u4_n127 ) , .A( u2_u15_u4_n136 ) , .B2( u2_u15_u4_n150 ) , .B1( u2_u15_u4_n180 ) );
  INV_X1 u2_u15_u4_U52 (.A( u2_u15_u4_n160 ) , .ZN( u2_u15_u4_n180 ) );
  NAND2_X1 u2_u15_u4_U53 (.A2( u2_u15_u4_n104 ) , .A1( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n146 ) );
  NAND2_X1 u2_u15_u4_U54 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n160 ) );
  NAND2_X1 u2_u15_u4_U55 (.ZN( u2_u15_u4_n134 ) , .A1( u2_u15_u4_n98 ) , .A2( u2_u15_u4_n99 ) );
  NAND2_X1 u2_u15_u4_U56 (.A1( u2_u15_u4_n103 ) , .A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n143 ) );
  NAND2_X1 u2_u15_u4_U57 (.A2( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n145 ) , .A1( u2_u15_u4_n98 ) );
  NAND2_X1 u2_u15_u4_U58 (.A1( u2_u15_u4_n100 ) , .A2( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n120 ) );
  NAND2_X1 u2_u15_u4_U59 (.A1( u2_u15_u4_n102 ) , .A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n148 ) );
  AOI21_X1 u2_u15_u4_U6 (.ZN( u2_u15_u4_n106 ) , .B2( u2_u15_u4_n146 ) , .B1( u2_u15_u4_n158 ) , .A( u2_u15_u4_n170 ) );
  NAND2_X1 u2_u15_u4_U60 (.A2( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n157 ) );
  INV_X1 u2_u15_u4_U61 (.A( u2_u15_u4_n150 ) , .ZN( u2_u15_u4_n173 ) );
  INV_X1 u2_u15_u4_U62 (.A( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n171 ) );
  NAND2_X1 u2_u15_u4_U63 (.A1( u2_u15_u4_n100 ) , .ZN( u2_u15_u4_n118 ) , .A2( u2_u15_u4_n99 ) );
  NAND2_X1 u2_u15_u4_U64 (.A2( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n144 ) );
  NAND2_X1 u2_u15_u4_U65 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n96 ) );
  INV_X1 u2_u15_u4_U66 (.A( u2_u15_u4_n128 ) , .ZN( u2_u15_u4_n174 ) );
  NAND2_X1 u2_u15_u4_U67 (.A2( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n119 ) , .A1( u2_u15_u4_n98 ) );
  NAND2_X1 u2_u15_u4_U68 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n147 ) );
  NAND2_X1 u2_u15_u4_U69 (.A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n113 ) , .A1( u2_u15_u4_n99 ) );
  AOI21_X1 u2_u15_u4_U7 (.ZN( u2_u15_u4_n108 ) , .B2( u2_u15_u4_n134 ) , .B1( u2_u15_u4_n155 ) , .A( u2_u15_u4_n156 ) );
  NOR2_X1 u2_u15_u4_U70 (.A2( u2_u15_X_28 ) , .ZN( u2_u15_u4_n150 ) , .A1( u2_u15_u4_n168 ) );
  NOR2_X1 u2_u15_u4_U71 (.A2( u2_u15_X_29 ) , .ZN( u2_u15_u4_n152 ) , .A1( u2_u15_u4_n169 ) );
  NOR2_X1 u2_u15_u4_U72 (.A2( u2_u15_X_26 ) , .ZN( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n177 ) );
  NOR2_X1 u2_u15_u4_U73 (.A2( u2_u15_X_30 ) , .ZN( u2_u15_u4_n105 ) , .A1( u2_u15_u4_n176 ) );
  NOR2_X1 u2_u15_u4_U74 (.A2( u2_u15_X_28 ) , .A1( u2_u15_X_29 ) , .ZN( u2_u15_u4_n128 ) );
  NOR2_X1 u2_u15_u4_U75 (.A2( u2_u15_X_25 ) , .A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n98 ) );
  NOR2_X1 u2_u15_u4_U76 (.A2( u2_u15_X_27 ) , .A1( u2_u15_X_30 ) , .ZN( u2_u15_u4_n102 ) );
  AND2_X1 u2_u15_u4_U77 (.A2( u2_u15_X_25 ) , .A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n104 ) );
  AND2_X1 u2_u15_u4_U78 (.A1( u2_u15_X_30 ) , .A2( u2_u15_u4_n176 ) , .ZN( u2_u15_u4_n99 ) );
  AND2_X1 u2_u15_u4_U79 (.A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n101 ) , .A2( u2_u15_u4_n177 ) );
  AOI21_X1 u2_u15_u4_U8 (.ZN( u2_u15_u4_n109 ) , .A( u2_u15_u4_n153 ) , .B1( u2_u15_u4_n159 ) , .B2( u2_u15_u4_n184 ) );
  AND2_X1 u2_u15_u4_U80 (.A1( u2_u15_X_27 ) , .A2( u2_u15_X_30 ) , .ZN( u2_u15_u4_n103 ) );
  INV_X1 u2_u15_u4_U81 (.A( u2_u15_X_28 ) , .ZN( u2_u15_u4_n169 ) );
  INV_X1 u2_u15_u4_U82 (.A( u2_u15_X_29 ) , .ZN( u2_u15_u4_n168 ) );
  INV_X1 u2_u15_u4_U83 (.A( u2_u15_X_25 ) , .ZN( u2_u15_u4_n177 ) );
  INV_X1 u2_u15_u4_U84 (.A( u2_u15_X_27 ) , .ZN( u2_u15_u4_n176 ) );
  NAND4_X1 u2_u15_u4_U85 (.ZN( u2_out15_14 ) , .A4( u2_u15_u4_n124 ) , .A3( u2_u15_u4_n125 ) , .A2( u2_u15_u4_n126 ) , .A1( u2_u15_u4_n127 ) );
  AOI22_X1 u2_u15_u4_U86 (.B2( u2_u15_u4_n117 ) , .ZN( u2_u15_u4_n126 ) , .A1( u2_u15_u4_n129 ) , .B1( u2_u15_u4_n152 ) , .A2( u2_u15_u4_n175 ) );
  AOI22_X1 u2_u15_u4_U87 (.ZN( u2_u15_u4_n125 ) , .B2( u2_u15_u4_n131 ) , .A2( u2_u15_u4_n132 ) , .B1( u2_u15_u4_n138 ) , .A1( u2_u15_u4_n178 ) );
  AOI22_X1 u2_u15_u4_U88 (.B2( u2_u15_u4_n149 ) , .B1( u2_u15_u4_n150 ) , .A2( u2_u15_u4_n151 ) , .A1( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n167 ) );
  NOR4_X1 u2_u15_u4_U89 (.A4( u2_u15_u4_n162 ) , .A3( u2_u15_u4_n163 ) , .A2( u2_u15_u4_n164 ) , .A1( u2_u15_u4_n165 ) , .ZN( u2_u15_u4_n166 ) );
  AOI211_X1 u2_u15_u4_U9 (.B( u2_u15_u4_n136 ) , .A( u2_u15_u4_n137 ) , .C2( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n139 ) , .C1( u2_u15_u4_n182 ) );
  NAND4_X1 u2_u15_u4_U90 (.ZN( u2_out15_8 ) , .A4( u2_u15_u4_n110 ) , .A3( u2_u15_u4_n111 ) , .A2( u2_u15_u4_n112 ) , .A1( u2_u15_u4_n186 ) );
  NAND2_X1 u2_u15_u4_U91 (.ZN( u2_u15_u4_n112 ) , .A2( u2_u15_u4_n130 ) , .A1( u2_u15_u4_n150 ) );
  AOI22_X1 u2_u15_u4_U92 (.ZN( u2_u15_u4_n111 ) , .B2( u2_u15_u4_n132 ) , .A1( u2_u15_u4_n152 ) , .B1( u2_u15_u4_n178 ) , .A2( u2_u15_u4_n97 ) );
  NAND4_X1 u2_u15_u4_U93 (.ZN( u2_out15_25 ) , .A4( u2_u15_u4_n139 ) , .A3( u2_u15_u4_n140 ) , .A2( u2_u15_u4_n141 ) , .A1( u2_u15_u4_n142 ) );
  OAI21_X1 u2_u15_u4_U94 (.A( u2_u15_u4_n128 ) , .B2( u2_u15_u4_n129 ) , .B1( u2_u15_u4_n130 ) , .ZN( u2_u15_u4_n142 ) );
  OAI21_X1 u2_u15_u4_U95 (.B2( u2_u15_u4_n131 ) , .ZN( u2_u15_u4_n141 ) , .A( u2_u15_u4_n175 ) , .B1( u2_u15_u4_n183 ) );
  NAND3_X1 u2_u15_u4_U96 (.ZN( u2_out15_3 ) , .A3( u2_u15_u4_n166 ) , .A1( u2_u15_u4_n167 ) , .A2( u2_u15_u4_n186 ) );
  NAND3_X1 u2_u15_u4_U97 (.A3( u2_u15_u4_n146 ) , .A2( u2_u15_u4_n147 ) , .A1( u2_u15_u4_n148 ) , .ZN( u2_u15_u4_n149 ) );
  NAND3_X1 u2_u15_u4_U98 (.A3( u2_u15_u4_n143 ) , .A2( u2_u15_u4_n144 ) , .A1( u2_u15_u4_n145 ) , .ZN( u2_u15_u4_n151 ) );
  NAND3_X1 u2_u15_u4_U99 (.A3( u2_u15_u4_n121 ) , .ZN( u2_u15_u4_n122 ) , .A2( u2_u15_u4_n144 ) , .A1( u2_u15_u4_n154 ) );
  INV_X1 u2_u15_u5_U10 (.A( u2_u15_u5_n121 ) , .ZN( u2_u15_u5_n177 ) );
  AOI222_X1 u2_u15_u5_U100 (.ZN( u2_u15_u5_n113 ) , .A1( u2_u15_u5_n131 ) , .C1( u2_u15_u5_n148 ) , .B2( u2_u15_u5_n174 ) , .C2( u2_u15_u5_n178 ) , .A2( u2_u15_u5_n179 ) , .B1( u2_u15_u5_n99 ) );
  NAND4_X1 u2_u15_u5_U101 (.ZN( u2_out15_29 ) , .A4( u2_u15_u5_n129 ) , .A3( u2_u15_u5_n130 ) , .A2( u2_u15_u5_n168 ) , .A1( u2_u15_u5_n196 ) );
  AOI221_X1 u2_u15_u5_U102 (.A( u2_u15_u5_n128 ) , .ZN( u2_u15_u5_n129 ) , .C2( u2_u15_u5_n132 ) , .B2( u2_u15_u5_n159 ) , .B1( u2_u15_u5_n176 ) , .C1( u2_u15_u5_n184 ) );
  AOI222_X1 u2_u15_u5_U103 (.ZN( u2_u15_u5_n130 ) , .A2( u2_u15_u5_n146 ) , .B1( u2_u15_u5_n147 ) , .C2( u2_u15_u5_n175 ) , .B2( u2_u15_u5_n179 ) , .A1( u2_u15_u5_n188 ) , .C1( u2_u15_u5_n194 ) );
  NAND3_X1 u2_u15_u5_U104 (.A2( u2_u15_u5_n154 ) , .A3( u2_u15_u5_n158 ) , .A1( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n99 ) );
  NOR2_X1 u2_u15_u5_U11 (.ZN( u2_u15_u5_n160 ) , .A2( u2_u15_u5_n173 ) , .A1( u2_u15_u5_n177 ) );
  INV_X1 u2_u15_u5_U12 (.A( u2_u15_u5_n150 ) , .ZN( u2_u15_u5_n174 ) );
  AOI21_X1 u2_u15_u5_U13 (.A( u2_u15_u5_n160 ) , .B2( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n162 ) , .B1( u2_u15_u5_n192 ) );
  INV_X1 u2_u15_u5_U14 (.A( u2_u15_u5_n159 ) , .ZN( u2_u15_u5_n192 ) );
  AOI21_X1 u2_u15_u5_U15 (.A( u2_u15_u5_n156 ) , .B2( u2_u15_u5_n157 ) , .B1( u2_u15_u5_n158 ) , .ZN( u2_u15_u5_n163 ) );
  AOI21_X1 u2_u15_u5_U16 (.B2( u2_u15_u5_n139 ) , .B1( u2_u15_u5_n140 ) , .ZN( u2_u15_u5_n141 ) , .A( u2_u15_u5_n150 ) );
  OAI21_X1 u2_u15_u5_U17 (.A( u2_u15_u5_n133 ) , .B2( u2_u15_u5_n134 ) , .B1( u2_u15_u5_n135 ) , .ZN( u2_u15_u5_n142 ) );
  OAI21_X1 u2_u15_u5_U18 (.ZN( u2_u15_u5_n133 ) , .B2( u2_u15_u5_n147 ) , .A( u2_u15_u5_n173 ) , .B1( u2_u15_u5_n188 ) );
  NAND2_X1 u2_u15_u5_U19 (.A2( u2_u15_u5_n119 ) , .A1( u2_u15_u5_n123 ) , .ZN( u2_u15_u5_n137 ) );
  INV_X1 u2_u15_u5_U20 (.A( u2_u15_u5_n155 ) , .ZN( u2_u15_u5_n194 ) );
  NAND2_X1 u2_u15_u5_U21 (.A1( u2_u15_u5_n121 ) , .ZN( u2_u15_u5_n132 ) , .A2( u2_u15_u5_n172 ) );
  NAND2_X1 u2_u15_u5_U22 (.A2( u2_u15_u5_n122 ) , .ZN( u2_u15_u5_n136 ) , .A1( u2_u15_u5_n154 ) );
  NAND2_X1 u2_u15_u5_U23 (.A2( u2_u15_u5_n119 ) , .A1( u2_u15_u5_n120 ) , .ZN( u2_u15_u5_n159 ) );
  INV_X1 u2_u15_u5_U24 (.A( u2_u15_u5_n156 ) , .ZN( u2_u15_u5_n175 ) );
  INV_X1 u2_u15_u5_U25 (.A( u2_u15_u5_n158 ) , .ZN( u2_u15_u5_n188 ) );
  INV_X1 u2_u15_u5_U26 (.A( u2_u15_u5_n152 ) , .ZN( u2_u15_u5_n179 ) );
  INV_X1 u2_u15_u5_U27 (.A( u2_u15_u5_n140 ) , .ZN( u2_u15_u5_n182 ) );
  INV_X1 u2_u15_u5_U28 (.A( u2_u15_u5_n151 ) , .ZN( u2_u15_u5_n183 ) );
  INV_X1 u2_u15_u5_U29 (.A( u2_u15_u5_n123 ) , .ZN( u2_u15_u5_n185 ) );
  NOR2_X1 u2_u15_u5_U3 (.ZN( u2_u15_u5_n134 ) , .A1( u2_u15_u5_n183 ) , .A2( u2_u15_u5_n190 ) );
  INV_X1 u2_u15_u5_U30 (.A( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n184 ) );
  INV_X1 u2_u15_u5_U31 (.A( u2_u15_u5_n139 ) , .ZN( u2_u15_u5_n189 ) );
  INV_X1 u2_u15_u5_U32 (.A( u2_u15_u5_n157 ) , .ZN( u2_u15_u5_n190 ) );
  INV_X1 u2_u15_u5_U33 (.A( u2_u15_u5_n120 ) , .ZN( u2_u15_u5_n193 ) );
  NAND2_X1 u2_u15_u5_U34 (.ZN( u2_u15_u5_n111 ) , .A1( u2_u15_u5_n140 ) , .A2( u2_u15_u5_n155 ) );
  NOR2_X1 u2_u15_u5_U35 (.ZN( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n170 ) , .A2( u2_u15_u5_n180 ) );
  INV_X1 u2_u15_u5_U36 (.A( u2_u15_u5_n117 ) , .ZN( u2_u15_u5_n196 ) );
  OAI221_X1 u2_u15_u5_U37 (.A( u2_u15_u5_n116 ) , .ZN( u2_u15_u5_n117 ) , .B2( u2_u15_u5_n119 ) , .C1( u2_u15_u5_n153 ) , .C2( u2_u15_u5_n158 ) , .B1( u2_u15_u5_n172 ) );
  AOI222_X1 u2_u15_u5_U38 (.ZN( u2_u15_u5_n116 ) , .B2( u2_u15_u5_n145 ) , .C1( u2_u15_u5_n148 ) , .A2( u2_u15_u5_n174 ) , .C2( u2_u15_u5_n177 ) , .B1( u2_u15_u5_n187 ) , .A1( u2_u15_u5_n193 ) );
  INV_X1 u2_u15_u5_U39 (.A( u2_u15_u5_n115 ) , .ZN( u2_u15_u5_n187 ) );
  INV_X1 u2_u15_u5_U4 (.A( u2_u15_u5_n138 ) , .ZN( u2_u15_u5_n191 ) );
  AOI22_X1 u2_u15_u5_U40 (.B2( u2_u15_u5_n131 ) , .A2( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n169 ) , .B1( u2_u15_u5_n174 ) , .A1( u2_u15_u5_n185 ) );
  NOR2_X1 u2_u15_u5_U41 (.A1( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n150 ) , .A2( u2_u15_u5_n173 ) );
  AOI21_X1 u2_u15_u5_U42 (.A( u2_u15_u5_n118 ) , .B2( u2_u15_u5_n145 ) , .ZN( u2_u15_u5_n168 ) , .B1( u2_u15_u5_n186 ) );
  INV_X1 u2_u15_u5_U43 (.A( u2_u15_u5_n122 ) , .ZN( u2_u15_u5_n186 ) );
  NOR2_X1 u2_u15_u5_U44 (.A1( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n152 ) , .A2( u2_u15_u5_n176 ) );
  NOR2_X1 u2_u15_u5_U45 (.A1( u2_u15_u5_n115 ) , .ZN( u2_u15_u5_n118 ) , .A2( u2_u15_u5_n153 ) );
  NOR2_X1 u2_u15_u5_U46 (.A2( u2_u15_u5_n145 ) , .ZN( u2_u15_u5_n156 ) , .A1( u2_u15_u5_n174 ) );
  NOR2_X1 u2_u15_u5_U47 (.ZN( u2_u15_u5_n121 ) , .A2( u2_u15_u5_n145 ) , .A1( u2_u15_u5_n176 ) );
  AOI22_X1 u2_u15_u5_U48 (.ZN( u2_u15_u5_n114 ) , .A2( u2_u15_u5_n137 ) , .A1( u2_u15_u5_n145 ) , .B2( u2_u15_u5_n175 ) , .B1( u2_u15_u5_n193 ) );
  OAI211_X1 u2_u15_u5_U49 (.B( u2_u15_u5_n124 ) , .A( u2_u15_u5_n125 ) , .C2( u2_u15_u5_n126 ) , .C1( u2_u15_u5_n127 ) , .ZN( u2_u15_u5_n128 ) );
  OAI21_X1 u2_u15_u5_U5 (.B2( u2_u15_u5_n136 ) , .B1( u2_u15_u5_n137 ) , .ZN( u2_u15_u5_n138 ) , .A( u2_u15_u5_n177 ) );
  NOR3_X1 u2_u15_u5_U50 (.ZN( u2_u15_u5_n127 ) , .A1( u2_u15_u5_n136 ) , .A3( u2_u15_u5_n148 ) , .A2( u2_u15_u5_n182 ) );
  OAI21_X1 u2_u15_u5_U51 (.ZN( u2_u15_u5_n124 ) , .A( u2_u15_u5_n177 ) , .B2( u2_u15_u5_n183 ) , .B1( u2_u15_u5_n189 ) );
  OAI21_X1 u2_u15_u5_U52 (.ZN( u2_u15_u5_n125 ) , .A( u2_u15_u5_n174 ) , .B2( u2_u15_u5_n185 ) , .B1( u2_u15_u5_n190 ) );
  AOI21_X1 u2_u15_u5_U53 (.A( u2_u15_u5_n153 ) , .B2( u2_u15_u5_n154 ) , .B1( u2_u15_u5_n155 ) , .ZN( u2_u15_u5_n164 ) );
  AOI21_X1 u2_u15_u5_U54 (.ZN( u2_u15_u5_n110 ) , .B1( u2_u15_u5_n122 ) , .B2( u2_u15_u5_n139 ) , .A( u2_u15_u5_n153 ) );
  INV_X1 u2_u15_u5_U55 (.A( u2_u15_u5_n153 ) , .ZN( u2_u15_u5_n176 ) );
  INV_X1 u2_u15_u5_U56 (.A( u2_u15_u5_n126 ) , .ZN( u2_u15_u5_n173 ) );
  AND2_X1 u2_u15_u5_U57 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n147 ) );
  AND2_X1 u2_u15_u5_U58 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n148 ) );
  NAND2_X1 u2_u15_u5_U59 (.A1( u2_u15_u5_n105 ) , .A2( u2_u15_u5_n106 ) , .ZN( u2_u15_u5_n158 ) );
  INV_X1 u2_u15_u5_U6 (.A( u2_u15_u5_n135 ) , .ZN( u2_u15_u5_n178 ) );
  NAND2_X1 u2_u15_u5_U60 (.A2( u2_u15_u5_n108 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n139 ) );
  NAND2_X1 u2_u15_u5_U61 (.A1( u2_u15_u5_n106 ) , .A2( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n119 ) );
  NAND2_X1 u2_u15_u5_U62 (.A2( u2_u15_u5_n103 ) , .A1( u2_u15_u5_n105 ) , .ZN( u2_u15_u5_n140 ) );
  NAND2_X1 u2_u15_u5_U63 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n105 ) , .ZN( u2_u15_u5_n155 ) );
  NAND2_X1 u2_u15_u5_U64 (.A2( u2_u15_u5_n106 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n122 ) );
  NAND2_X1 u2_u15_u5_U65 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n106 ) , .ZN( u2_u15_u5_n115 ) );
  NAND2_X1 u2_u15_u5_U66 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n103 ) , .ZN( u2_u15_u5_n161 ) );
  NAND2_X1 u2_u15_u5_U67 (.A1( u2_u15_u5_n105 ) , .A2( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n154 ) );
  INV_X1 u2_u15_u5_U68 (.A( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n172 ) );
  NAND2_X1 u2_u15_u5_U69 (.A1( u2_u15_u5_n103 ) , .A2( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n123 ) );
  OAI22_X1 u2_u15_u5_U7 (.B2( u2_u15_u5_n149 ) , .B1( u2_u15_u5_n150 ) , .A2( u2_u15_u5_n151 ) , .A1( u2_u15_u5_n152 ) , .ZN( u2_u15_u5_n165 ) );
  NAND2_X1 u2_u15_u5_U70 (.A2( u2_u15_u5_n103 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n151 ) );
  NAND2_X1 u2_u15_u5_U71 (.A2( u2_u15_u5_n107 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n120 ) );
  NAND2_X1 u2_u15_u5_U72 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n157 ) );
  AND2_X1 u2_u15_u5_U73 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n104 ) , .ZN( u2_u15_u5_n131 ) );
  INV_X1 u2_u15_u5_U74 (.A( u2_u15_u5_n102 ) , .ZN( u2_u15_u5_n195 ) );
  OAI221_X1 u2_u15_u5_U75 (.A( u2_u15_u5_n101 ) , .ZN( u2_u15_u5_n102 ) , .C2( u2_u15_u5_n115 ) , .C1( u2_u15_u5_n126 ) , .B1( u2_u15_u5_n134 ) , .B2( u2_u15_u5_n160 ) );
  OAI21_X1 u2_u15_u5_U76 (.ZN( u2_u15_u5_n101 ) , .B1( u2_u15_u5_n137 ) , .A( u2_u15_u5_n146 ) , .B2( u2_u15_u5_n147 ) );
  NOR2_X1 u2_u15_u5_U77 (.A2( u2_u15_X_34 ) , .A1( u2_u15_X_35 ) , .ZN( u2_u15_u5_n145 ) );
  NOR2_X1 u2_u15_u5_U78 (.A2( u2_u15_X_34 ) , .ZN( u2_u15_u5_n146 ) , .A1( u2_u15_u5_n171 ) );
  NOR2_X1 u2_u15_u5_U79 (.A2( u2_u15_X_31 ) , .A1( u2_u15_X_32 ) , .ZN( u2_u15_u5_n103 ) );
  NOR3_X1 u2_u15_u5_U8 (.A2( u2_u15_u5_n147 ) , .A1( u2_u15_u5_n148 ) , .ZN( u2_u15_u5_n149 ) , .A3( u2_u15_u5_n194 ) );
  NOR2_X1 u2_u15_u5_U80 (.A2( u2_u15_X_36 ) , .ZN( u2_u15_u5_n105 ) , .A1( u2_u15_u5_n180 ) );
  NOR2_X1 u2_u15_u5_U81 (.A2( u2_u15_X_33 ) , .ZN( u2_u15_u5_n108 ) , .A1( u2_u15_u5_n170 ) );
  NOR2_X1 u2_u15_u5_U82 (.A2( u2_u15_X_33 ) , .A1( u2_u15_X_36 ) , .ZN( u2_u15_u5_n107 ) );
  NOR2_X1 u2_u15_u5_U83 (.A2( u2_u15_X_31 ) , .ZN( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n181 ) );
  NAND2_X1 u2_u15_u5_U84 (.A2( u2_u15_X_34 ) , .A1( u2_u15_X_35 ) , .ZN( u2_u15_u5_n153 ) );
  NAND2_X1 u2_u15_u5_U85 (.A1( u2_u15_X_34 ) , .ZN( u2_u15_u5_n126 ) , .A2( u2_u15_u5_n171 ) );
  AND2_X1 u2_u15_u5_U86 (.A1( u2_u15_X_31 ) , .A2( u2_u15_X_32 ) , .ZN( u2_u15_u5_n106 ) );
  AND2_X1 u2_u15_u5_U87 (.A1( u2_u15_X_31 ) , .ZN( u2_u15_u5_n109 ) , .A2( u2_u15_u5_n181 ) );
  INV_X1 u2_u15_u5_U88 (.A( u2_u15_X_33 ) , .ZN( u2_u15_u5_n180 ) );
  INV_X1 u2_u15_u5_U89 (.A( u2_u15_X_35 ) , .ZN( u2_u15_u5_n171 ) );
  NOR2_X1 u2_u15_u5_U9 (.ZN( u2_u15_u5_n135 ) , .A1( u2_u15_u5_n173 ) , .A2( u2_u15_u5_n176 ) );
  INV_X1 u2_u15_u5_U90 (.A( u2_u15_X_36 ) , .ZN( u2_u15_u5_n170 ) );
  INV_X1 u2_u15_u5_U91 (.A( u2_u15_X_32 ) , .ZN( u2_u15_u5_n181 ) );
  NAND4_X1 u2_u15_u5_U92 (.ZN( u2_out15_19 ) , .A4( u2_u15_u5_n166 ) , .A3( u2_u15_u5_n167 ) , .A2( u2_u15_u5_n168 ) , .A1( u2_u15_u5_n169 ) );
  AOI22_X1 u2_u15_u5_U93 (.B2( u2_u15_u5_n145 ) , .A2( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n167 ) , .B1( u2_u15_u5_n182 ) , .A1( u2_u15_u5_n189 ) );
  NOR4_X1 u2_u15_u5_U94 (.A4( u2_u15_u5_n162 ) , .A3( u2_u15_u5_n163 ) , .A2( u2_u15_u5_n164 ) , .A1( u2_u15_u5_n165 ) , .ZN( u2_u15_u5_n166 ) );
  NAND4_X1 u2_u15_u5_U95 (.ZN( u2_out15_11 ) , .A4( u2_u15_u5_n143 ) , .A3( u2_u15_u5_n144 ) , .A2( u2_u15_u5_n169 ) , .A1( u2_u15_u5_n196 ) );
  AOI22_X1 u2_u15_u5_U96 (.A2( u2_u15_u5_n132 ) , .ZN( u2_u15_u5_n144 ) , .B2( u2_u15_u5_n145 ) , .B1( u2_u15_u5_n184 ) , .A1( u2_u15_u5_n194 ) );
  NOR3_X1 u2_u15_u5_U97 (.A3( u2_u15_u5_n141 ) , .A1( u2_u15_u5_n142 ) , .ZN( u2_u15_u5_n143 ) , .A2( u2_u15_u5_n191 ) );
  NAND4_X1 u2_u15_u5_U98 (.ZN( u2_out15_4 ) , .A4( u2_u15_u5_n112 ) , .A2( u2_u15_u5_n113 ) , .A1( u2_u15_u5_n114 ) , .A3( u2_u15_u5_n195 ) );
  AOI211_X1 u2_u15_u5_U99 (.A( u2_u15_u5_n110 ) , .C1( u2_u15_u5_n111 ) , .ZN( u2_u15_u5_n112 ) , .B( u2_u15_u5_n118 ) , .C2( u2_u15_u5_n177 ) );
  INV_X1 u2_u15_u6_U10 (.ZN( u2_u15_u6_n172 ) , .A( u2_u15_u6_n88 ) );
  OAI21_X1 u2_u15_u6_U11 (.A( u2_u15_u6_n159 ) , .B1( u2_u15_u6_n169 ) , .B2( u2_u15_u6_n173 ) , .ZN( u2_u15_u6_n90 ) );
  AOI22_X1 u2_u15_u6_U12 (.A2( u2_u15_u6_n151 ) , .B2( u2_u15_u6_n161 ) , .A1( u2_u15_u6_n167 ) , .B1( u2_u15_u6_n170 ) , .ZN( u2_u15_u6_n89 ) );
  AOI21_X1 u2_u15_u6_U13 (.ZN( u2_u15_u6_n106 ) , .A( u2_u15_u6_n142 ) , .B2( u2_u15_u6_n159 ) , .B1( u2_u15_u6_n164 ) );
  INV_X1 u2_u15_u6_U14 (.A( u2_u15_u6_n155 ) , .ZN( u2_u15_u6_n161 ) );
  INV_X1 u2_u15_u6_U15 (.A( u2_u15_u6_n128 ) , .ZN( u2_u15_u6_n164 ) );
  NAND2_X1 u2_u15_u6_U16 (.ZN( u2_u15_u6_n110 ) , .A1( u2_u15_u6_n122 ) , .A2( u2_u15_u6_n129 ) );
  NAND2_X1 u2_u15_u6_U17 (.ZN( u2_u15_u6_n124 ) , .A2( u2_u15_u6_n146 ) , .A1( u2_u15_u6_n148 ) );
  INV_X1 u2_u15_u6_U18 (.A( u2_u15_u6_n132 ) , .ZN( u2_u15_u6_n171 ) );
  AND2_X1 u2_u15_u6_U19 (.A1( u2_u15_u6_n100 ) , .ZN( u2_u15_u6_n130 ) , .A2( u2_u15_u6_n147 ) );
  INV_X1 u2_u15_u6_U20 (.A( u2_u15_u6_n127 ) , .ZN( u2_u15_u6_n173 ) );
  INV_X1 u2_u15_u6_U21 (.A( u2_u15_u6_n121 ) , .ZN( u2_u15_u6_n167 ) );
  INV_X1 u2_u15_u6_U22 (.A( u2_u15_u6_n100 ) , .ZN( u2_u15_u6_n169 ) );
  INV_X1 u2_u15_u6_U23 (.A( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n170 ) );
  INV_X1 u2_u15_u6_U24 (.A( u2_u15_u6_n113 ) , .ZN( u2_u15_u6_n168 ) );
  AND2_X1 u2_u15_u6_U25 (.A1( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n119 ) , .ZN( u2_u15_u6_n133 ) );
  AND2_X1 u2_u15_u6_U26 (.A2( u2_u15_u6_n121 ) , .A1( u2_u15_u6_n122 ) , .ZN( u2_u15_u6_n131 ) );
  AND3_X1 u2_u15_u6_U27 (.ZN( u2_u15_u6_n120 ) , .A2( u2_u15_u6_n127 ) , .A1( u2_u15_u6_n132 ) , .A3( u2_u15_u6_n145 ) );
  INV_X1 u2_u15_u6_U28 (.A( u2_u15_u6_n146 ) , .ZN( u2_u15_u6_n163 ) );
  AOI222_X1 u2_u15_u6_U29 (.ZN( u2_u15_u6_n114 ) , .A1( u2_u15_u6_n118 ) , .A2( u2_u15_u6_n126 ) , .B2( u2_u15_u6_n151 ) , .C2( u2_u15_u6_n159 ) , .C1( u2_u15_u6_n168 ) , .B1( u2_u15_u6_n169 ) );
  INV_X1 u2_u15_u6_U3 (.A( u2_u15_u6_n110 ) , .ZN( u2_u15_u6_n166 ) );
  NOR2_X1 u2_u15_u6_U30 (.A1( u2_u15_u6_n162 ) , .A2( u2_u15_u6_n165 ) , .ZN( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U31 (.A1( u2_u15_u6_n144 ) , .ZN( u2_u15_u6_n151 ) , .A2( u2_u15_u6_n158 ) );
  NAND2_X1 u2_u15_u6_U32 (.ZN( u2_u15_u6_n132 ) , .A1( u2_u15_u6_n91 ) , .A2( u2_u15_u6_n97 ) );
  AOI22_X1 u2_u15_u6_U33 (.B2( u2_u15_u6_n110 ) , .B1( u2_u15_u6_n111 ) , .A1( u2_u15_u6_n112 ) , .ZN( u2_u15_u6_n115 ) , .A2( u2_u15_u6_n161 ) );
  NAND4_X1 u2_u15_u6_U34 (.A3( u2_u15_u6_n109 ) , .ZN( u2_u15_u6_n112 ) , .A4( u2_u15_u6_n132 ) , .A2( u2_u15_u6_n147 ) , .A1( u2_u15_u6_n166 ) );
  NOR2_X1 u2_u15_u6_U35 (.ZN( u2_u15_u6_n109 ) , .A1( u2_u15_u6_n170 ) , .A2( u2_u15_u6_n173 ) );
  NOR2_X1 u2_u15_u6_U36 (.A2( u2_u15_u6_n126 ) , .ZN( u2_u15_u6_n155 ) , .A1( u2_u15_u6_n160 ) );
  NAND2_X1 u2_u15_u6_U37 (.ZN( u2_u15_u6_n146 ) , .A2( u2_u15_u6_n94 ) , .A1( u2_u15_u6_n99 ) );
  AOI21_X1 u2_u15_u6_U38 (.A( u2_u15_u6_n144 ) , .B2( u2_u15_u6_n145 ) , .B1( u2_u15_u6_n146 ) , .ZN( u2_u15_u6_n150 ) );
  AOI211_X1 u2_u15_u6_U39 (.B( u2_u15_u6_n134 ) , .A( u2_u15_u6_n135 ) , .C1( u2_u15_u6_n136 ) , .ZN( u2_u15_u6_n137 ) , .C2( u2_u15_u6_n151 ) );
  INV_X1 u2_u15_u6_U4 (.A( u2_u15_u6_n142 ) , .ZN( u2_u15_u6_n174 ) );
  NAND4_X1 u2_u15_u6_U40 (.A4( u2_u15_u6_n127 ) , .A3( u2_u15_u6_n128 ) , .A2( u2_u15_u6_n129 ) , .A1( u2_u15_u6_n130 ) , .ZN( u2_u15_u6_n136 ) );
  AOI21_X1 u2_u15_u6_U41 (.B2( u2_u15_u6_n132 ) , .B1( u2_u15_u6_n133 ) , .ZN( u2_u15_u6_n134 ) , .A( u2_u15_u6_n158 ) );
  AOI21_X1 u2_u15_u6_U42 (.B1( u2_u15_u6_n131 ) , .ZN( u2_u15_u6_n135 ) , .A( u2_u15_u6_n144 ) , .B2( u2_u15_u6_n146 ) );
  INV_X1 u2_u15_u6_U43 (.A( u2_u15_u6_n111 ) , .ZN( u2_u15_u6_n158 ) );
  NAND2_X1 u2_u15_u6_U44 (.ZN( u2_u15_u6_n127 ) , .A1( u2_u15_u6_n91 ) , .A2( u2_u15_u6_n92 ) );
  NAND2_X1 u2_u15_u6_U45 (.ZN( u2_u15_u6_n129 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n96 ) );
  INV_X1 u2_u15_u6_U46 (.A( u2_u15_u6_n144 ) , .ZN( u2_u15_u6_n159 ) );
  NAND2_X1 u2_u15_u6_U47 (.ZN( u2_u15_u6_n145 ) , .A2( u2_u15_u6_n97 ) , .A1( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U48 (.ZN( u2_u15_u6_n148 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n94 ) );
  NAND2_X1 u2_u15_u6_U49 (.ZN( u2_u15_u6_n108 ) , .A2( u2_u15_u6_n139 ) , .A1( u2_u15_u6_n144 ) );
  NAND2_X1 u2_u15_u6_U5 (.A2( u2_u15_u6_n143 ) , .ZN( u2_u15_u6_n152 ) , .A1( u2_u15_u6_n166 ) );
  NAND2_X1 u2_u15_u6_U50 (.ZN( u2_u15_u6_n121 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n97 ) );
  NAND2_X1 u2_u15_u6_U51 (.ZN( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n95 ) );
  AND2_X1 u2_u15_u6_U52 (.ZN( u2_u15_u6_n118 ) , .A2( u2_u15_u6_n91 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U53 (.ZN( u2_u15_u6_n147 ) , .A2( u2_u15_u6_n98 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U54 (.ZN( u2_u15_u6_n128 ) , .A1( u2_u15_u6_n94 ) , .A2( u2_u15_u6_n96 ) );
  NAND2_X1 u2_u15_u6_U55 (.ZN( u2_u15_u6_n119 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U56 (.ZN( u2_u15_u6_n123 ) , .A2( u2_u15_u6_n91 ) , .A1( u2_u15_u6_n96 ) );
  NAND2_X1 u2_u15_u6_U57 (.ZN( u2_u15_u6_n100 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U58 (.ZN( u2_u15_u6_n122 ) , .A1( u2_u15_u6_n94 ) , .A2( u2_u15_u6_n97 ) );
  INV_X1 u2_u15_u6_U59 (.A( u2_u15_u6_n139 ) , .ZN( u2_u15_u6_n160 ) );
  AOI22_X1 u2_u15_u6_U6 (.B2( u2_u15_u6_n101 ) , .A1( u2_u15_u6_n102 ) , .ZN( u2_u15_u6_n103 ) , .B1( u2_u15_u6_n160 ) , .A2( u2_u15_u6_n161 ) );
  NAND2_X1 u2_u15_u6_U60 (.ZN( u2_u15_u6_n113 ) , .A1( u2_u15_u6_n96 ) , .A2( u2_u15_u6_n98 ) );
  NOR2_X1 u2_u15_u6_U61 (.A2( u2_u15_X_40 ) , .A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n126 ) );
  NOR2_X1 u2_u15_u6_U62 (.A2( u2_u15_X_39 ) , .A1( u2_u15_X_42 ) , .ZN( u2_u15_u6_n92 ) );
  NOR2_X1 u2_u15_u6_U63 (.A2( u2_u15_X_39 ) , .A1( u2_u15_u6_n156 ) , .ZN( u2_u15_u6_n97 ) );
  NOR2_X1 u2_u15_u6_U64 (.A2( u2_u15_X_38 ) , .A1( u2_u15_u6_n165 ) , .ZN( u2_u15_u6_n95 ) );
  NOR2_X1 u2_u15_u6_U65 (.A2( u2_u15_X_41 ) , .ZN( u2_u15_u6_n111 ) , .A1( u2_u15_u6_n157 ) );
  NOR2_X1 u2_u15_u6_U66 (.A2( u2_u15_X_37 ) , .A1( u2_u15_u6_n162 ) , .ZN( u2_u15_u6_n94 ) );
  NOR2_X1 u2_u15_u6_U67 (.A2( u2_u15_X_37 ) , .A1( u2_u15_X_38 ) , .ZN( u2_u15_u6_n91 ) );
  NAND2_X1 u2_u15_u6_U68 (.A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n144 ) , .A2( u2_u15_u6_n157 ) );
  NAND2_X1 u2_u15_u6_U69 (.A2( u2_u15_X_40 ) , .A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n139 ) );
  NOR2_X1 u2_u15_u6_U7 (.A1( u2_u15_u6_n118 ) , .ZN( u2_u15_u6_n143 ) , .A2( u2_u15_u6_n168 ) );
  AND2_X1 u2_u15_u6_U70 (.A1( u2_u15_X_39 ) , .A2( u2_u15_u6_n156 ) , .ZN( u2_u15_u6_n96 ) );
  AND2_X1 u2_u15_u6_U71 (.A1( u2_u15_X_39 ) , .A2( u2_u15_X_42 ) , .ZN( u2_u15_u6_n99 ) );
  INV_X1 u2_u15_u6_U72 (.A( u2_u15_X_40 ) , .ZN( u2_u15_u6_n157 ) );
  INV_X1 u2_u15_u6_U73 (.A( u2_u15_X_37 ) , .ZN( u2_u15_u6_n165 ) );
  INV_X1 u2_u15_u6_U74 (.A( u2_u15_X_38 ) , .ZN( u2_u15_u6_n162 ) );
  INV_X1 u2_u15_u6_U75 (.A( u2_u15_X_42 ) , .ZN( u2_u15_u6_n156 ) );
  NAND4_X1 u2_u15_u6_U76 (.ZN( u2_out15_12 ) , .A4( u2_u15_u6_n114 ) , .A3( u2_u15_u6_n115 ) , .A2( u2_u15_u6_n116 ) , .A1( u2_u15_u6_n117 ) );
  OAI22_X1 u2_u15_u6_U77 (.B2( u2_u15_u6_n111 ) , .ZN( u2_u15_u6_n116 ) , .B1( u2_u15_u6_n126 ) , .A2( u2_u15_u6_n164 ) , .A1( u2_u15_u6_n167 ) );
  OAI21_X1 u2_u15_u6_U78 (.A( u2_u15_u6_n108 ) , .ZN( u2_u15_u6_n117 ) , .B2( u2_u15_u6_n141 ) , .B1( u2_u15_u6_n163 ) );
  NAND4_X1 u2_u15_u6_U79 (.ZN( u2_out15_32 ) , .A4( u2_u15_u6_n103 ) , .A3( u2_u15_u6_n104 ) , .A2( u2_u15_u6_n105 ) , .A1( u2_u15_u6_n106 ) );
  AOI21_X1 u2_u15_u6_U8 (.B1( u2_u15_u6_n107 ) , .B2( u2_u15_u6_n132 ) , .A( u2_u15_u6_n158 ) , .ZN( u2_u15_u6_n88 ) );
  AOI22_X1 u2_u15_u6_U80 (.ZN( u2_u15_u6_n105 ) , .A2( u2_u15_u6_n108 ) , .A1( u2_u15_u6_n118 ) , .B2( u2_u15_u6_n126 ) , .B1( u2_u15_u6_n171 ) );
  AOI22_X1 u2_u15_u6_U81 (.ZN( u2_u15_u6_n104 ) , .A1( u2_u15_u6_n111 ) , .B1( u2_u15_u6_n124 ) , .B2( u2_u15_u6_n151 ) , .A2( u2_u15_u6_n93 ) );
  OAI211_X1 u2_u15_u6_U82 (.ZN( u2_out15_22 ) , .B( u2_u15_u6_n137 ) , .A( u2_u15_u6_n138 ) , .C2( u2_u15_u6_n139 ) , .C1( u2_u15_u6_n140 ) );
  AOI22_X1 u2_u15_u6_U83 (.B1( u2_u15_u6_n124 ) , .A2( u2_u15_u6_n125 ) , .A1( u2_u15_u6_n126 ) , .ZN( u2_u15_u6_n138 ) , .B2( u2_u15_u6_n161 ) );
  AND4_X1 u2_u15_u6_U84 (.A3( u2_u15_u6_n119 ) , .A1( u2_u15_u6_n120 ) , .A4( u2_u15_u6_n129 ) , .ZN( u2_u15_u6_n140 ) , .A2( u2_u15_u6_n143 ) );
  OAI211_X1 u2_u15_u6_U85 (.ZN( u2_out15_7 ) , .B( u2_u15_u6_n153 ) , .C2( u2_u15_u6_n154 ) , .C1( u2_u15_u6_n155 ) , .A( u2_u15_u6_n174 ) );
  NOR3_X1 u2_u15_u6_U86 (.A1( u2_u15_u6_n141 ) , .ZN( u2_u15_u6_n154 ) , .A3( u2_u15_u6_n164 ) , .A2( u2_u15_u6_n171 ) );
  AOI211_X1 u2_u15_u6_U87 (.B( u2_u15_u6_n149 ) , .A( u2_u15_u6_n150 ) , .C2( u2_u15_u6_n151 ) , .C1( u2_u15_u6_n152 ) , .ZN( u2_u15_u6_n153 ) );
  NAND3_X1 u2_u15_u6_U88 (.A2( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n125 ) , .A1( u2_u15_u6_n130 ) , .A3( u2_u15_u6_n131 ) );
  NAND3_X1 u2_u15_u6_U89 (.A3( u2_u15_u6_n133 ) , .ZN( u2_u15_u6_n141 ) , .A1( u2_u15_u6_n145 ) , .A2( u2_u15_u6_n148 ) );
  AOI21_X1 u2_u15_u6_U9 (.B2( u2_u15_u6_n147 ) , .B1( u2_u15_u6_n148 ) , .ZN( u2_u15_u6_n149 ) , .A( u2_u15_u6_n158 ) );
  NAND3_X1 u2_u15_u6_U90 (.ZN( u2_u15_u6_n101 ) , .A3( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n121 ) , .A1( u2_u15_u6_n127 ) );
  NAND3_X1 u2_u15_u6_U91 (.ZN( u2_u15_u6_n102 ) , .A3( u2_u15_u6_n130 ) , .A2( u2_u15_u6_n145 ) , .A1( u2_u15_u6_n166 ) );
  NAND3_X1 u2_u15_u6_U92 (.A3( u2_u15_u6_n113 ) , .A1( u2_u15_u6_n119 ) , .A2( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n93 ) );
  NAND3_X1 u2_u15_u6_U93 (.ZN( u2_u15_u6_n142 ) , .A2( u2_u15_u6_n172 ) , .A3( u2_u15_u6_n89 ) , .A1( u2_u15_u6_n90 ) );
  OAI21_X1 u2_u15_u7_U10 (.A( u2_u15_u7_n161 ) , .B1( u2_u15_u7_n168 ) , .B2( u2_u15_u7_n173 ) , .ZN( u2_u15_u7_n91 ) );
  AOI211_X1 u2_u15_u7_U11 (.A( u2_u15_u7_n117 ) , .ZN( u2_u15_u7_n118 ) , .C2( u2_u15_u7_n126 ) , .C1( u2_u15_u7_n177 ) , .B( u2_u15_u7_n180 ) );
  OAI22_X1 u2_u15_u7_U12 (.B1( u2_u15_u7_n115 ) , .ZN( u2_u15_u7_n117 ) , .A2( u2_u15_u7_n133 ) , .A1( u2_u15_u7_n137 ) , .B2( u2_u15_u7_n162 ) );
  INV_X1 u2_u15_u7_U13 (.A( u2_u15_u7_n116 ) , .ZN( u2_u15_u7_n180 ) );
  NOR3_X1 u2_u15_u7_U14 (.ZN( u2_u15_u7_n115 ) , .A3( u2_u15_u7_n145 ) , .A2( u2_u15_u7_n168 ) , .A1( u2_u15_u7_n169 ) );
  OAI211_X1 u2_u15_u7_U15 (.B( u2_u15_u7_n122 ) , .A( u2_u15_u7_n123 ) , .C2( u2_u15_u7_n124 ) , .ZN( u2_u15_u7_n154 ) , .C1( u2_u15_u7_n162 ) );
  AOI222_X1 u2_u15_u7_U16 (.ZN( u2_u15_u7_n122 ) , .C2( u2_u15_u7_n126 ) , .C1( u2_u15_u7_n145 ) , .B1( u2_u15_u7_n161 ) , .A2( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n170 ) , .A1( u2_u15_u7_n176 ) );
  INV_X1 u2_u15_u7_U17 (.A( u2_u15_u7_n133 ) , .ZN( u2_u15_u7_n176 ) );
  NOR3_X1 u2_u15_u7_U18 (.A2( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n135 ) , .ZN( u2_u15_u7_n136 ) , .A3( u2_u15_u7_n171 ) );
  NOR2_X1 u2_u15_u7_U19 (.A1( u2_u15_u7_n130 ) , .A2( u2_u15_u7_n134 ) , .ZN( u2_u15_u7_n153 ) );
  INV_X1 u2_u15_u7_U20 (.A( u2_u15_u7_n101 ) , .ZN( u2_u15_u7_n165 ) );
  NOR2_X1 u2_u15_u7_U21 (.ZN( u2_u15_u7_n111 ) , .A2( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n169 ) );
  AOI21_X1 u2_u15_u7_U22 (.ZN( u2_u15_u7_n104 ) , .B2( u2_u15_u7_n112 ) , .B1( u2_u15_u7_n127 ) , .A( u2_u15_u7_n164 ) );
  AOI21_X1 u2_u15_u7_U23 (.ZN( u2_u15_u7_n106 ) , .B1( u2_u15_u7_n133 ) , .B2( u2_u15_u7_n146 ) , .A( u2_u15_u7_n162 ) );
  AOI21_X1 u2_u15_u7_U24 (.A( u2_u15_u7_n101 ) , .ZN( u2_u15_u7_n107 ) , .B2( u2_u15_u7_n128 ) , .B1( u2_u15_u7_n175 ) );
  INV_X1 u2_u15_u7_U25 (.A( u2_u15_u7_n138 ) , .ZN( u2_u15_u7_n171 ) );
  INV_X1 u2_u15_u7_U26 (.A( u2_u15_u7_n131 ) , .ZN( u2_u15_u7_n177 ) );
  INV_X1 u2_u15_u7_U27 (.A( u2_u15_u7_n110 ) , .ZN( u2_u15_u7_n174 ) );
  NAND2_X1 u2_u15_u7_U28 (.A1( u2_u15_u7_n129 ) , .A2( u2_u15_u7_n132 ) , .ZN( u2_u15_u7_n149 ) );
  NAND2_X1 u2_u15_u7_U29 (.A1( u2_u15_u7_n113 ) , .A2( u2_u15_u7_n124 ) , .ZN( u2_u15_u7_n130 ) );
  INV_X1 u2_u15_u7_U3 (.A( u2_u15_u7_n111 ) , .ZN( u2_u15_u7_n170 ) );
  INV_X1 u2_u15_u7_U30 (.A( u2_u15_u7_n112 ) , .ZN( u2_u15_u7_n173 ) );
  INV_X1 u2_u15_u7_U31 (.A( u2_u15_u7_n128 ) , .ZN( u2_u15_u7_n168 ) );
  INV_X1 u2_u15_u7_U32 (.A( u2_u15_u7_n148 ) , .ZN( u2_u15_u7_n169 ) );
  INV_X1 u2_u15_u7_U33 (.A( u2_u15_u7_n127 ) , .ZN( u2_u15_u7_n179 ) );
  NOR2_X1 u2_u15_u7_U34 (.ZN( u2_u15_u7_n101 ) , .A2( u2_u15_u7_n150 ) , .A1( u2_u15_u7_n156 ) );
  AOI211_X1 u2_u15_u7_U35 (.B( u2_u15_u7_n154 ) , .A( u2_u15_u7_n155 ) , .C1( u2_u15_u7_n156 ) , .ZN( u2_u15_u7_n157 ) , .C2( u2_u15_u7_n172 ) );
  INV_X1 u2_u15_u7_U36 (.A( u2_u15_u7_n153 ) , .ZN( u2_u15_u7_n172 ) );
  AOI211_X1 u2_u15_u7_U37 (.B( u2_u15_u7_n139 ) , .A( u2_u15_u7_n140 ) , .C2( u2_u15_u7_n141 ) , .ZN( u2_u15_u7_n142 ) , .C1( u2_u15_u7_n156 ) );
  NAND4_X1 u2_u15_u7_U38 (.A3( u2_u15_u7_n127 ) , .A2( u2_u15_u7_n128 ) , .A1( u2_u15_u7_n129 ) , .ZN( u2_u15_u7_n141 ) , .A4( u2_u15_u7_n147 ) );
  AOI21_X1 u2_u15_u7_U39 (.A( u2_u15_u7_n137 ) , .B1( u2_u15_u7_n138 ) , .ZN( u2_u15_u7_n139 ) , .B2( u2_u15_u7_n146 ) );
  INV_X1 u2_u15_u7_U4 (.A( u2_u15_u7_n149 ) , .ZN( u2_u15_u7_n175 ) );
  OAI22_X1 u2_u15_u7_U40 (.B1( u2_u15_u7_n136 ) , .ZN( u2_u15_u7_n140 ) , .A1( u2_u15_u7_n153 ) , .B2( u2_u15_u7_n162 ) , .A2( u2_u15_u7_n164 ) );
  AOI21_X1 u2_u15_u7_U41 (.ZN( u2_u15_u7_n123 ) , .B1( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n177 ) , .A( u2_u15_u7_n97 ) );
  AOI21_X1 u2_u15_u7_U42 (.B2( u2_u15_u7_n113 ) , .B1( u2_u15_u7_n124 ) , .A( u2_u15_u7_n125 ) , .ZN( u2_u15_u7_n97 ) );
  INV_X1 u2_u15_u7_U43 (.A( u2_u15_u7_n125 ) , .ZN( u2_u15_u7_n161 ) );
  INV_X1 u2_u15_u7_U44 (.A( u2_u15_u7_n152 ) , .ZN( u2_u15_u7_n162 ) );
  AOI22_X1 u2_u15_u7_U45 (.A2( u2_u15_u7_n114 ) , .ZN( u2_u15_u7_n119 ) , .B1( u2_u15_u7_n130 ) , .A1( u2_u15_u7_n156 ) , .B2( u2_u15_u7_n165 ) );
  NAND2_X1 u2_u15_u7_U46 (.A2( u2_u15_u7_n112 ) , .ZN( u2_u15_u7_n114 ) , .A1( u2_u15_u7_n175 ) );
  AOI22_X1 u2_u15_u7_U47 (.B2( u2_u15_u7_n149 ) , .B1( u2_u15_u7_n150 ) , .A2( u2_u15_u7_n151 ) , .A1( u2_u15_u7_n152 ) , .ZN( u2_u15_u7_n158 ) );
  AND2_X1 u2_u15_u7_U48 (.ZN( u2_u15_u7_n145 ) , .A2( u2_u15_u7_n98 ) , .A1( u2_u15_u7_n99 ) );
  NOR2_X1 u2_u15_u7_U49 (.ZN( u2_u15_u7_n137 ) , .A1( u2_u15_u7_n150 ) , .A2( u2_u15_u7_n161 ) );
  INV_X1 u2_u15_u7_U5 (.A( u2_u15_u7_n154 ) , .ZN( u2_u15_u7_n178 ) );
  AOI21_X1 u2_u15_u7_U50 (.ZN( u2_u15_u7_n105 ) , .B2( u2_u15_u7_n110 ) , .A( u2_u15_u7_n125 ) , .B1( u2_u15_u7_n147 ) );
  NAND2_X1 u2_u15_u7_U51 (.ZN( u2_u15_u7_n146 ) , .A1( u2_u15_u7_n95 ) , .A2( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U52 (.A2( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n147 ) , .A1( u2_u15_u7_n93 ) );
  NAND2_X1 u2_u15_u7_U53 (.A1( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n127 ) , .A2( u2_u15_u7_n99 ) );
  OR2_X1 u2_u15_u7_U54 (.ZN( u2_u15_u7_n126 ) , .A2( u2_u15_u7_n152 ) , .A1( u2_u15_u7_n156 ) );
  NAND2_X1 u2_u15_u7_U55 (.A2( u2_u15_u7_n102 ) , .A1( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n133 ) );
  NAND2_X1 u2_u15_u7_U56 (.ZN( u2_u15_u7_n112 ) , .A2( u2_u15_u7_n96 ) , .A1( u2_u15_u7_n99 ) );
  NAND2_X1 u2_u15_u7_U57 (.A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n128 ) , .A1( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U58 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n113 ) , .A2( u2_u15_u7_n93 ) );
  NAND2_X1 u2_u15_u7_U59 (.A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n124 ) , .A1( u2_u15_u7_n96 ) );
  AOI211_X1 u2_u15_u7_U6 (.ZN( u2_u15_u7_n116 ) , .A( u2_u15_u7_n155 ) , .C1( u2_u15_u7_n161 ) , .C2( u2_u15_u7_n171 ) , .B( u2_u15_u7_n94 ) );
  NAND2_X1 u2_u15_u7_U60 (.ZN( u2_u15_u7_n110 ) , .A1( u2_u15_u7_n95 ) , .A2( u2_u15_u7_n96 ) );
  INV_X1 u2_u15_u7_U61 (.A( u2_u15_u7_n150 ) , .ZN( u2_u15_u7_n164 ) );
  AND2_X1 u2_u15_u7_U62 (.ZN( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n93 ) , .A2( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U63 (.A1( u2_u15_u7_n100 ) , .A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n129 ) );
  NAND2_X1 u2_u15_u7_U64 (.A2( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n131 ) , .A1( u2_u15_u7_n95 ) );
  NAND2_X1 u2_u15_u7_U65 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n138 ) , .A2( u2_u15_u7_n99 ) );
  NAND2_X1 u2_u15_u7_U66 (.ZN( u2_u15_u7_n132 ) , .A1( u2_u15_u7_n93 ) , .A2( u2_u15_u7_n96 ) );
  NAND2_X1 u2_u15_u7_U67 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n148 ) , .A2( u2_u15_u7_n95 ) );
  NOR2_X1 u2_u15_u7_U68 (.A2( u2_u15_X_47 ) , .ZN( u2_u15_u7_n150 ) , .A1( u2_u15_u7_n163 ) );
  NOR2_X1 u2_u15_u7_U69 (.A2( u2_u15_X_43 ) , .A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n103 ) );
  OAI222_X1 u2_u15_u7_U7 (.C2( u2_u15_u7_n101 ) , .B2( u2_u15_u7_n111 ) , .A1( u2_u15_u7_n113 ) , .C1( u2_u15_u7_n146 ) , .A2( u2_u15_u7_n162 ) , .B1( u2_u15_u7_n164 ) , .ZN( u2_u15_u7_n94 ) );
  NOR2_X1 u2_u15_u7_U70 (.A2( u2_u15_X_48 ) , .A1( u2_u15_u7_n166 ) , .ZN( u2_u15_u7_n95 ) );
  NOR2_X1 u2_u15_u7_U71 (.A2( u2_u15_X_45 ) , .A1( u2_u15_X_48 ) , .ZN( u2_u15_u7_n99 ) );
  NOR2_X1 u2_u15_u7_U72 (.A2( u2_u15_X_44 ) , .A1( u2_u15_u7_n167 ) , .ZN( u2_u15_u7_n98 ) );
  NOR2_X1 u2_u15_u7_U73 (.A2( u2_u15_X_46 ) , .A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n152 ) );
  AND2_X1 u2_u15_u7_U74 (.A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n156 ) , .A2( u2_u15_u7_n163 ) );
  NAND2_X1 u2_u15_u7_U75 (.A2( u2_u15_X_46 ) , .A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n125 ) );
  AND2_X1 u2_u15_u7_U76 (.A2( u2_u15_X_45 ) , .A1( u2_u15_X_48 ) , .ZN( u2_u15_u7_n102 ) );
  AND2_X1 u2_u15_u7_U77 (.A2( u2_u15_X_43 ) , .A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n96 ) );
  AND2_X1 u2_u15_u7_U78 (.A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n100 ) , .A2( u2_u15_u7_n167 ) );
  AND2_X1 u2_u15_u7_U79 (.A1( u2_u15_X_48 ) , .A2( u2_u15_u7_n166 ) , .ZN( u2_u15_u7_n93 ) );
  OAI221_X1 u2_u15_u7_U8 (.C1( u2_u15_u7_n101 ) , .C2( u2_u15_u7_n147 ) , .ZN( u2_u15_u7_n155 ) , .B2( u2_u15_u7_n162 ) , .A( u2_u15_u7_n91 ) , .B1( u2_u15_u7_n92 ) );
  INV_X1 u2_u15_u7_U80 (.A( u2_u15_X_46 ) , .ZN( u2_u15_u7_n163 ) );
  INV_X1 u2_u15_u7_U81 (.A( u2_u15_X_45 ) , .ZN( u2_u15_u7_n166 ) );
  INV_X1 u2_u15_u7_U82 (.A( u2_u15_X_43 ) , .ZN( u2_u15_u7_n167 ) );
  NAND4_X1 u2_u15_u7_U83 (.ZN( u2_out15_5 ) , .A4( u2_u15_u7_n108 ) , .A3( u2_u15_u7_n109 ) , .A1( u2_u15_u7_n116 ) , .A2( u2_u15_u7_n123 ) );
  AOI22_X1 u2_u15_u7_U84 (.ZN( u2_u15_u7_n109 ) , .A2( u2_u15_u7_n126 ) , .B2( u2_u15_u7_n145 ) , .B1( u2_u15_u7_n156 ) , .A1( u2_u15_u7_n171 ) );
  NOR4_X1 u2_u15_u7_U85 (.A4( u2_u15_u7_n104 ) , .A3( u2_u15_u7_n105 ) , .A2( u2_u15_u7_n106 ) , .A1( u2_u15_u7_n107 ) , .ZN( u2_u15_u7_n108 ) );
  NAND4_X1 u2_u15_u7_U86 (.ZN( u2_out15_27 ) , .A4( u2_u15_u7_n118 ) , .A3( u2_u15_u7_n119 ) , .A2( u2_u15_u7_n120 ) , .A1( u2_u15_u7_n121 ) );
  OAI21_X1 u2_u15_u7_U87 (.ZN( u2_u15_u7_n121 ) , .B2( u2_u15_u7_n145 ) , .A( u2_u15_u7_n150 ) , .B1( u2_u15_u7_n174 ) );
  OAI21_X1 u2_u15_u7_U88 (.ZN( u2_u15_u7_n120 ) , .A( u2_u15_u7_n161 ) , .B2( u2_u15_u7_n170 ) , .B1( u2_u15_u7_n179 ) );
  NAND4_X1 u2_u15_u7_U89 (.ZN( u2_out15_21 ) , .A4( u2_u15_u7_n157 ) , .A3( u2_u15_u7_n158 ) , .A2( u2_u15_u7_n159 ) , .A1( u2_u15_u7_n160 ) );
  AND3_X1 u2_u15_u7_U9 (.A3( u2_u15_u7_n110 ) , .A2( u2_u15_u7_n127 ) , .A1( u2_u15_u7_n132 ) , .ZN( u2_u15_u7_n92 ) );
  OAI21_X1 u2_u15_u7_U90 (.B1( u2_u15_u7_n145 ) , .ZN( u2_u15_u7_n160 ) , .A( u2_u15_u7_n161 ) , .B2( u2_u15_u7_n177 ) );
  OAI21_X1 u2_u15_u7_U91 (.ZN( u2_u15_u7_n159 ) , .A( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n171 ) , .B1( u2_u15_u7_n174 ) );
  NAND4_X1 u2_u15_u7_U92 (.ZN( u2_out15_15 ) , .A4( u2_u15_u7_n142 ) , .A3( u2_u15_u7_n143 ) , .A2( u2_u15_u7_n144 ) , .A1( u2_u15_u7_n178 ) );
  OR2_X1 u2_u15_u7_U93 (.A2( u2_u15_u7_n125 ) , .A1( u2_u15_u7_n129 ) , .ZN( u2_u15_u7_n144 ) );
  AOI22_X1 u2_u15_u7_U94 (.A2( u2_u15_u7_n126 ) , .ZN( u2_u15_u7_n143 ) , .B2( u2_u15_u7_n165 ) , .B1( u2_u15_u7_n173 ) , .A1( u2_u15_u7_n174 ) );
  NAND3_X1 u2_u15_u7_U95 (.A3( u2_u15_u7_n146 ) , .A2( u2_u15_u7_n147 ) , .A1( u2_u15_u7_n148 ) , .ZN( u2_u15_u7_n151 ) );
  NAND3_X1 u2_u15_u7_U96 (.A3( u2_u15_u7_n131 ) , .A2( u2_u15_u7_n132 ) , .A1( u2_u15_u7_n133 ) , .ZN( u2_u15_u7_n135 ) );
  XOR2_X1 u2_u7_U12 (.B( u2_K8_43 ) , .A( u2_R6_28 ) , .Z( u2_u7_X_43 ) );
  XOR2_X1 u2_u7_U16 (.B( u2_K8_3 ) , .A( u2_R6_2 ) , .Z( u2_u7_X_3 ) );
  XOR2_X1 u2_u7_U2 (.B( u2_K8_8 ) , .A( u2_R6_5 ) , .Z( u2_u7_X_8 ) );
  XOR2_X1 u2_u7_U27 (.B( u2_K8_2 ) , .A( u2_R6_1 ) , .Z( u2_u7_X_2 ) );
  XOR2_X1 u2_u7_U3 (.B( u2_K8_7 ) , .A( u2_R6_4 ) , .Z( u2_u7_X_7 ) );
  XOR2_X1 u2_u7_U37 (.B( u2_K8_20 ) , .A( u2_R6_13 ) , .Z( u2_u7_X_20 ) );
  XOR2_X1 u2_u7_U38 (.B( u2_K8_1 ) , .A( u2_R6_32 ) , .Z( u2_u7_X_1 ) );
  XOR2_X1 u2_u7_U39 (.B( u2_K8_19 ) , .A( u2_R6_12 ) , .Z( u2_u7_X_19 ) );
  XOR2_X1 u2_u7_U4 (.B( u2_K8_6 ) , .A( u2_R6_5 ) , .Z( u2_u7_X_6 ) );
  XOR2_X1 u2_u7_U40 (.B( u2_K8_18 ) , .A( u2_R6_13 ) , .Z( u2_u7_X_18 ) );
  XOR2_X1 u2_u7_U41 (.B( u2_K8_17 ) , .A( u2_R6_12 ) , .Z( u2_u7_X_17 ) );
  XOR2_X1 u2_u7_U44 (.B( u2_K8_14 ) , .A( u2_R6_9 ) , .Z( u2_u7_X_14 ) );
  XOR2_X1 u2_u7_U45 (.B( u2_K8_13 ) , .A( u2_R6_8 ) , .Z( u2_u7_X_13 ) );
  XOR2_X1 u2_u7_U46 (.B( u2_K8_12 ) , .A( u2_R6_9 ) , .Z( u2_u7_X_12 ) );
  XOR2_X1 u2_u7_U47 (.B( u2_K8_11 ) , .A( u2_R6_8 ) , .Z( u2_u7_X_11 ) );
  XOR2_X1 u2_u7_U5 (.B( u2_K8_5 ) , .A( u2_R6_4 ) , .Z( u2_u7_X_5 ) );
  XOR2_X1 u2_u7_U7 (.B( u2_K8_48 ) , .A( u2_R6_1 ) , .Z( u2_u7_X_48 ) );
  XOR2_X1 u2_u7_U8 (.B( u2_K8_47 ) , .A( u2_R6_32 ) , .Z( u2_u7_X_47 ) );
  AND3_X1 u2_u7_u0_U10 (.A2( u2_u7_u0_n112 ) , .ZN( u2_u7_u0_n127 ) , .A3( u2_u7_u0_n130 ) , .A1( u2_u7_u0_n148 ) );
  NAND2_X1 u2_u7_u0_U11 (.ZN( u2_u7_u0_n113 ) , .A1( u2_u7_u0_n139 ) , .A2( u2_u7_u0_n149 ) );
  AND2_X1 u2_u7_u0_U12 (.ZN( u2_u7_u0_n107 ) , .A1( u2_u7_u0_n130 ) , .A2( u2_u7_u0_n140 ) );
  AND2_X1 u2_u7_u0_U13 (.A2( u2_u7_u0_n129 ) , .A1( u2_u7_u0_n130 ) , .ZN( u2_u7_u0_n151 ) );
  AND2_X1 u2_u7_u0_U14 (.A1( u2_u7_u0_n108 ) , .A2( u2_u7_u0_n125 ) , .ZN( u2_u7_u0_n145 ) );
  INV_X1 u2_u7_u0_U15 (.A( u2_u7_u0_n143 ) , .ZN( u2_u7_u0_n173 ) );
  NOR2_X1 u2_u7_u0_U16 (.A2( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n147 ) , .A1( u2_u7_u0_n160 ) );
  INV_X1 u2_u7_u0_U17 (.ZN( u2_u7_u0_n172 ) , .A( u2_u7_u0_n88 ) );
  OAI222_X1 u2_u7_u0_U18 (.C1( u2_u7_u0_n108 ) , .A1( u2_u7_u0_n125 ) , .B2( u2_u7_u0_n128 ) , .B1( u2_u7_u0_n144 ) , .A2( u2_u7_u0_n158 ) , .C2( u2_u7_u0_n161 ) , .ZN( u2_u7_u0_n88 ) );
  NOR2_X1 u2_u7_u0_U19 (.A1( u2_u7_u0_n163 ) , .A2( u2_u7_u0_n164 ) , .ZN( u2_u7_u0_n95 ) );
  OAI22_X1 u2_u7_u0_U20 (.B1( u2_u7_u0_n125 ) , .ZN( u2_u7_u0_n126 ) , .A1( u2_u7_u0_n138 ) , .A2( u2_u7_u0_n146 ) , .B2( u2_u7_u0_n147 ) );
  OAI22_X1 u2_u7_u0_U21 (.B1( u2_u7_u0_n131 ) , .A1( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n147 ) , .A2( u2_u7_u0_n90 ) , .ZN( u2_u7_u0_n91 ) );
  AND3_X1 u2_u7_u0_U22 (.A3( u2_u7_u0_n121 ) , .A2( u2_u7_u0_n125 ) , .A1( u2_u7_u0_n148 ) , .ZN( u2_u7_u0_n90 ) );
  INV_X1 u2_u7_u0_U23 (.A( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n161 ) );
  AOI22_X1 u2_u7_u0_U24 (.B2( u2_u7_u0_n109 ) , .A2( u2_u7_u0_n110 ) , .ZN( u2_u7_u0_n111 ) , .B1( u2_u7_u0_n118 ) , .A1( u2_u7_u0_n160 ) );
  INV_X1 u2_u7_u0_U25 (.A( u2_u7_u0_n118 ) , .ZN( u2_u7_u0_n158 ) );
  AOI21_X1 u2_u7_u0_U26 (.ZN( u2_u7_u0_n104 ) , .B1( u2_u7_u0_n107 ) , .B2( u2_u7_u0_n141 ) , .A( u2_u7_u0_n144 ) );
  AOI21_X1 u2_u7_u0_U27 (.B1( u2_u7_u0_n127 ) , .B2( u2_u7_u0_n129 ) , .A( u2_u7_u0_n138 ) , .ZN( u2_u7_u0_n96 ) );
  AOI21_X1 u2_u7_u0_U28 (.ZN( u2_u7_u0_n116 ) , .B2( u2_u7_u0_n142 ) , .A( u2_u7_u0_n144 ) , .B1( u2_u7_u0_n166 ) );
  INV_X1 u2_u7_u0_U29 (.ZN( u2_u7_u0_n171 ) , .A( u2_u7_u0_n99 ) );
  INV_X1 u2_u7_u0_U3 (.A( u2_u7_u0_n113 ) , .ZN( u2_u7_u0_n166 ) );
  OAI211_X1 u2_u7_u0_U30 (.C2( u2_u7_u0_n140 ) , .C1( u2_u7_u0_n161 ) , .A( u2_u7_u0_n169 ) , .B( u2_u7_u0_n98 ) , .ZN( u2_u7_u0_n99 ) );
  INV_X1 u2_u7_u0_U31 (.ZN( u2_u7_u0_n169 ) , .A( u2_u7_u0_n91 ) );
  AOI211_X1 u2_u7_u0_U32 (.C1( u2_u7_u0_n118 ) , .A( u2_u7_u0_n123 ) , .B( u2_u7_u0_n96 ) , .C2( u2_u7_u0_n97 ) , .ZN( u2_u7_u0_n98 ) );
  NOR2_X1 u2_u7_u0_U33 (.A1( u2_u7_u0_n120 ) , .ZN( u2_u7_u0_n143 ) , .A2( u2_u7_u0_n167 ) );
  OAI221_X1 u2_u7_u0_U34 (.C1( u2_u7_u0_n112 ) , .ZN( u2_u7_u0_n120 ) , .B1( u2_u7_u0_n138 ) , .B2( u2_u7_u0_n141 ) , .C2( u2_u7_u0_n147 ) , .A( u2_u7_u0_n172 ) );
  AOI211_X1 u2_u7_u0_U35 (.B( u2_u7_u0_n115 ) , .A( u2_u7_u0_n116 ) , .C2( u2_u7_u0_n117 ) , .C1( u2_u7_u0_n118 ) , .ZN( u2_u7_u0_n119 ) );
  NAND2_X1 u2_u7_u0_U36 (.A1( u2_u7_u0_n101 ) , .A2( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n150 ) );
  INV_X1 u2_u7_u0_U37 (.A( u2_u7_u0_n138 ) , .ZN( u2_u7_u0_n160 ) );
  NAND2_X1 u2_u7_u0_U38 (.A1( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n128 ) , .A2( u2_u7_u0_n95 ) );
  NAND2_X1 u2_u7_u0_U39 (.ZN( u2_u7_u0_n148 ) , .A1( u2_u7_u0_n93 ) , .A2( u2_u7_u0_n95 ) );
  AOI21_X1 u2_u7_u0_U4 (.B1( u2_u7_u0_n114 ) , .ZN( u2_u7_u0_n115 ) , .B2( u2_u7_u0_n129 ) , .A( u2_u7_u0_n161 ) );
  NAND2_X1 u2_u7_u0_U40 (.A2( u2_u7_u0_n102 ) , .A1( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n149 ) );
  NAND2_X1 u2_u7_u0_U41 (.A2( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n114 ) , .A1( u2_u7_u0_n92 ) );
  NAND2_X1 u2_u7_u0_U42 (.A2( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n121 ) , .A1( u2_u7_u0_n93 ) );
  NAND2_X1 u2_u7_u0_U43 (.ZN( u2_u7_u0_n112 ) , .A2( u2_u7_u0_n92 ) , .A1( u2_u7_u0_n93 ) );
  AOI21_X1 u2_u7_u0_U44 (.B1( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n132 ) , .A( u2_u7_u0_n165 ) , .B2( u2_u7_u0_n93 ) );
  INV_X1 u2_u7_u0_U45 (.A( u2_u7_u0_n142 ) , .ZN( u2_u7_u0_n165 ) );
  OR3_X1 u2_u7_u0_U46 (.A3( u2_u7_u0_n152 ) , .A2( u2_u7_u0_n153 ) , .A1( u2_u7_u0_n154 ) , .ZN( u2_u7_u0_n155 ) );
  AOI21_X1 u2_u7_u0_U47 (.A( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n145 ) , .B1( u2_u7_u0_n146 ) , .ZN( u2_u7_u0_n154 ) );
  AOI21_X1 u2_u7_u0_U48 (.B2( u2_u7_u0_n150 ) , .B1( u2_u7_u0_n151 ) , .ZN( u2_u7_u0_n152 ) , .A( u2_u7_u0_n158 ) );
  AOI21_X1 u2_u7_u0_U49 (.A( u2_u7_u0_n147 ) , .B2( u2_u7_u0_n148 ) , .B1( u2_u7_u0_n149 ) , .ZN( u2_u7_u0_n153 ) );
  AOI21_X1 u2_u7_u0_U5 (.B2( u2_u7_u0_n131 ) , .ZN( u2_u7_u0_n134 ) , .B1( u2_u7_u0_n151 ) , .A( u2_u7_u0_n158 ) );
  NOR2_X1 u2_u7_u0_U50 (.A2( u2_u7_X_4 ) , .A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n118 ) );
  NAND2_X1 u2_u7_u0_U51 (.A2( u2_u7_X_4 ) , .A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n144 ) );
  NOR2_X1 u2_u7_u0_U52 (.A2( u2_u7_X_1 ) , .A1( u2_u7_X_2 ) , .ZN( u2_u7_u0_n92 ) );
  NOR2_X1 u2_u7_u0_U53 (.A2( u2_u7_X_1 ) , .ZN( u2_u7_u0_n101 ) , .A1( u2_u7_u0_n163 ) );
  NOR2_X1 u2_u7_u0_U54 (.A2( u2_u7_X_2 ) , .ZN( u2_u7_u0_n103 ) , .A1( u2_u7_u0_n164 ) );
  NOR2_X1 u2_u7_u0_U55 (.A2( u2_u7_X_5 ) , .ZN( u2_u7_u0_n136 ) , .A1( u2_u7_u0_n159 ) );
  NAND2_X1 u2_u7_u0_U56 (.A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n138 ) , .A2( u2_u7_u0_n159 ) );
  AND2_X1 u2_u7_u0_U57 (.A2( u2_u7_X_3 ) , .A1( u2_u7_X_6 ) , .ZN( u2_u7_u0_n102 ) );
  AND2_X1 u2_u7_u0_U58 (.A1( u2_u7_X_6 ) , .A2( u2_u7_u0_n162 ) , .ZN( u2_u7_u0_n93 ) );
  INV_X1 u2_u7_u0_U59 (.A( u2_u7_X_4 ) , .ZN( u2_u7_u0_n159 ) );
  NOR2_X1 u2_u7_u0_U6 (.A1( u2_u7_u0_n108 ) , .ZN( u2_u7_u0_n123 ) , .A2( u2_u7_u0_n158 ) );
  INV_X1 u2_u7_u0_U60 (.A( u2_u7_X_1 ) , .ZN( u2_u7_u0_n164 ) );
  INV_X1 u2_u7_u0_U61 (.A( u2_u7_X_2 ) , .ZN( u2_u7_u0_n163 ) );
  INV_X1 u2_u7_u0_U62 (.A( u2_u7_u0_n126 ) , .ZN( u2_u7_u0_n168 ) );
  AOI211_X1 u2_u7_u0_U63 (.B( u2_u7_u0_n133 ) , .A( u2_u7_u0_n134 ) , .C2( u2_u7_u0_n135 ) , .C1( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n137 ) );
  OR4_X1 u2_u7_u0_U64 (.ZN( u2_out7_17 ) , .A4( u2_u7_u0_n122 ) , .A2( u2_u7_u0_n123 ) , .A1( u2_u7_u0_n124 ) , .A3( u2_u7_u0_n170 ) );
  AOI21_X1 u2_u7_u0_U65 (.B2( u2_u7_u0_n107 ) , .ZN( u2_u7_u0_n124 ) , .B1( u2_u7_u0_n128 ) , .A( u2_u7_u0_n161 ) );
  INV_X1 u2_u7_u0_U66 (.A( u2_u7_u0_n111 ) , .ZN( u2_u7_u0_n170 ) );
  OR4_X1 u2_u7_u0_U67 (.ZN( u2_out7_31 ) , .A4( u2_u7_u0_n155 ) , .A2( u2_u7_u0_n156 ) , .A1( u2_u7_u0_n157 ) , .A3( u2_u7_u0_n173 ) );
  AOI21_X1 u2_u7_u0_U68 (.A( u2_u7_u0_n138 ) , .B2( u2_u7_u0_n139 ) , .B1( u2_u7_u0_n140 ) , .ZN( u2_u7_u0_n157 ) );
  AOI21_X1 u2_u7_u0_U69 (.B2( u2_u7_u0_n141 ) , .B1( u2_u7_u0_n142 ) , .ZN( u2_u7_u0_n156 ) , .A( u2_u7_u0_n161 ) );
  OAI21_X1 u2_u7_u0_U7 (.B1( u2_u7_u0_n150 ) , .B2( u2_u7_u0_n158 ) , .A( u2_u7_u0_n172 ) , .ZN( u2_u7_u0_n89 ) );
  INV_X1 u2_u7_u0_U70 (.ZN( u2_u7_u0_n174 ) , .A( u2_u7_u0_n89 ) );
  AOI211_X1 u2_u7_u0_U71 (.B( u2_u7_u0_n104 ) , .A( u2_u7_u0_n105 ) , .ZN( u2_u7_u0_n106 ) , .C2( u2_u7_u0_n113 ) , .C1( u2_u7_u0_n160 ) );
  NAND2_X1 u2_u7_u0_U72 (.A2( u2_u7_u0_n100 ) , .A1( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n139 ) );
  NAND2_X1 u2_u7_u0_U73 (.A1( u2_u7_u0_n100 ) , .A2( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n125 ) );
  NAND2_X1 u2_u7_u0_U74 (.A1( u2_u7_u0_n100 ) , .ZN( u2_u7_u0_n129 ) , .A2( u2_u7_u0_n95 ) );
  NAND2_X1 u2_u7_u0_U75 (.A2( u2_u7_u0_n100 ) , .ZN( u2_u7_u0_n131 ) , .A1( u2_u7_u0_n92 ) );
  OAI221_X1 u2_u7_u0_U76 (.C1( u2_u7_u0_n121 ) , .ZN( u2_u7_u0_n122 ) , .B2( u2_u7_u0_n127 ) , .A( u2_u7_u0_n143 ) , .B1( u2_u7_u0_n144 ) , .C2( u2_u7_u0_n147 ) );
  NOR2_X1 u2_u7_u0_U77 (.A2( u2_u7_X_6 ) , .ZN( u2_u7_u0_n100 ) , .A1( u2_u7_u0_n162 ) );
  AOI21_X1 u2_u7_u0_U78 (.B1( u2_u7_u0_n132 ) , .ZN( u2_u7_u0_n133 ) , .A( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n166 ) );
  OAI22_X1 u2_u7_u0_U79 (.ZN( u2_u7_u0_n105 ) , .A2( u2_u7_u0_n132 ) , .B1( u2_u7_u0_n146 ) , .A1( u2_u7_u0_n147 ) , .B2( u2_u7_u0_n161 ) );
  AND2_X1 u2_u7_u0_U8 (.A1( u2_u7_u0_n114 ) , .A2( u2_u7_u0_n121 ) , .ZN( u2_u7_u0_n146 ) );
  NAND2_X1 u2_u7_u0_U80 (.ZN( u2_u7_u0_n110 ) , .A2( u2_u7_u0_n132 ) , .A1( u2_u7_u0_n145 ) );
  INV_X1 u2_u7_u0_U81 (.A( u2_u7_u0_n119 ) , .ZN( u2_u7_u0_n167 ) );
  NAND2_X1 u2_u7_u0_U82 (.A2( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n140 ) , .A1( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U83 (.A1( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n130 ) , .A2( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U84 (.ZN( u2_u7_u0_n108 ) , .A1( u2_u7_u0_n92 ) , .A2( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U85 (.ZN( u2_u7_u0_n142 ) , .A1( u2_u7_u0_n94 ) , .A2( u2_u7_u0_n95 ) );
  INV_X1 u2_u7_u0_U86 (.A( u2_u7_X_3 ) , .ZN( u2_u7_u0_n162 ) );
  NOR2_X1 u2_u7_u0_U87 (.A2( u2_u7_X_3 ) , .A1( u2_u7_X_6 ) , .ZN( u2_u7_u0_n94 ) );
  NAND3_X1 u2_u7_u0_U88 (.ZN( u2_out7_23 ) , .A3( u2_u7_u0_n137 ) , .A1( u2_u7_u0_n168 ) , .A2( u2_u7_u0_n171 ) );
  NAND3_X1 u2_u7_u0_U89 (.A3( u2_u7_u0_n127 ) , .A2( u2_u7_u0_n128 ) , .ZN( u2_u7_u0_n135 ) , .A1( u2_u7_u0_n150 ) );
  AND2_X1 u2_u7_u0_U9 (.A1( u2_u7_u0_n131 ) , .ZN( u2_u7_u0_n141 ) , .A2( u2_u7_u0_n150 ) );
  NAND3_X1 u2_u7_u0_U90 (.ZN( u2_u7_u0_n117 ) , .A3( u2_u7_u0_n132 ) , .A2( u2_u7_u0_n139 ) , .A1( u2_u7_u0_n148 ) );
  NAND3_X1 u2_u7_u0_U91 (.ZN( u2_u7_u0_n109 ) , .A2( u2_u7_u0_n114 ) , .A3( u2_u7_u0_n140 ) , .A1( u2_u7_u0_n149 ) );
  NAND3_X1 u2_u7_u0_U92 (.ZN( u2_out7_9 ) , .A3( u2_u7_u0_n106 ) , .A2( u2_u7_u0_n171 ) , .A1( u2_u7_u0_n174 ) );
  NAND3_X1 u2_u7_u0_U93 (.A2( u2_u7_u0_n128 ) , .A1( u2_u7_u0_n132 ) , .A3( u2_u7_u0_n146 ) , .ZN( u2_u7_u0_n97 ) );
  AOI21_X1 u2_u7_u1_U10 (.B2( u2_u7_u1_n155 ) , .B1( u2_u7_u1_n156 ) , .ZN( u2_u7_u1_n157 ) , .A( u2_u7_u1_n174 ) );
  NAND3_X1 u2_u7_u1_U100 (.ZN( u2_u7_u1_n113 ) , .A1( u2_u7_u1_n120 ) , .A3( u2_u7_u1_n133 ) , .A2( u2_u7_u1_n155 ) );
  NAND2_X1 u2_u7_u1_U11 (.ZN( u2_u7_u1_n140 ) , .A2( u2_u7_u1_n150 ) , .A1( u2_u7_u1_n155 ) );
  NAND2_X1 u2_u7_u1_U12 (.A1( u2_u7_u1_n131 ) , .ZN( u2_u7_u1_n147 ) , .A2( u2_u7_u1_n153 ) );
  AOI22_X1 u2_u7_u1_U13 (.B2( u2_u7_u1_n136 ) , .A2( u2_u7_u1_n137 ) , .ZN( u2_u7_u1_n143 ) , .A1( u2_u7_u1_n171 ) , .B1( u2_u7_u1_n173 ) );
  INV_X1 u2_u7_u1_U14 (.A( u2_u7_u1_n147 ) , .ZN( u2_u7_u1_n181 ) );
  INV_X1 u2_u7_u1_U15 (.A( u2_u7_u1_n139 ) , .ZN( u2_u7_u1_n174 ) );
  OR4_X1 u2_u7_u1_U16 (.A4( u2_u7_u1_n106 ) , .A3( u2_u7_u1_n107 ) , .ZN( u2_u7_u1_n108 ) , .A1( u2_u7_u1_n117 ) , .A2( u2_u7_u1_n184 ) );
  AOI21_X1 u2_u7_u1_U17 (.ZN( u2_u7_u1_n106 ) , .A( u2_u7_u1_n112 ) , .B1( u2_u7_u1_n154 ) , .B2( u2_u7_u1_n156 ) );
  AOI21_X1 u2_u7_u1_U18 (.ZN( u2_u7_u1_n107 ) , .B1( u2_u7_u1_n134 ) , .B2( u2_u7_u1_n149 ) , .A( u2_u7_u1_n174 ) );
  INV_X1 u2_u7_u1_U19 (.A( u2_u7_u1_n101 ) , .ZN( u2_u7_u1_n184 ) );
  INV_X1 u2_u7_u1_U20 (.A( u2_u7_u1_n112 ) , .ZN( u2_u7_u1_n171 ) );
  NAND2_X1 u2_u7_u1_U21 (.ZN( u2_u7_u1_n141 ) , .A1( u2_u7_u1_n153 ) , .A2( u2_u7_u1_n156 ) );
  AND2_X1 u2_u7_u1_U22 (.A1( u2_u7_u1_n123 ) , .ZN( u2_u7_u1_n134 ) , .A2( u2_u7_u1_n161 ) );
  NAND2_X1 u2_u7_u1_U23 (.A2( u2_u7_u1_n115 ) , .A1( u2_u7_u1_n116 ) , .ZN( u2_u7_u1_n148 ) );
  NAND2_X1 u2_u7_u1_U24 (.A2( u2_u7_u1_n133 ) , .A1( u2_u7_u1_n135 ) , .ZN( u2_u7_u1_n159 ) );
  NAND2_X1 u2_u7_u1_U25 (.A2( u2_u7_u1_n115 ) , .A1( u2_u7_u1_n120 ) , .ZN( u2_u7_u1_n132 ) );
  INV_X1 u2_u7_u1_U26 (.A( u2_u7_u1_n154 ) , .ZN( u2_u7_u1_n178 ) );
  INV_X1 u2_u7_u1_U27 (.A( u2_u7_u1_n151 ) , .ZN( u2_u7_u1_n183 ) );
  AND2_X1 u2_u7_u1_U28 (.A1( u2_u7_u1_n129 ) , .A2( u2_u7_u1_n133 ) , .ZN( u2_u7_u1_n149 ) );
  INV_X1 u2_u7_u1_U29 (.A( u2_u7_u1_n131 ) , .ZN( u2_u7_u1_n180 ) );
  INV_X1 u2_u7_u1_U3 (.A( u2_u7_u1_n159 ) , .ZN( u2_u7_u1_n182 ) );
  OAI221_X1 u2_u7_u1_U30 (.A( u2_u7_u1_n119 ) , .C2( u2_u7_u1_n129 ) , .ZN( u2_u7_u1_n138 ) , .B2( u2_u7_u1_n152 ) , .C1( u2_u7_u1_n174 ) , .B1( u2_u7_u1_n187 ) );
  INV_X1 u2_u7_u1_U31 (.A( u2_u7_u1_n148 ) , .ZN( u2_u7_u1_n187 ) );
  AOI211_X1 u2_u7_u1_U32 (.B( u2_u7_u1_n117 ) , .A( u2_u7_u1_n118 ) , .ZN( u2_u7_u1_n119 ) , .C2( u2_u7_u1_n146 ) , .C1( u2_u7_u1_n159 ) );
  NOR2_X1 u2_u7_u1_U33 (.A1( u2_u7_u1_n168 ) , .A2( u2_u7_u1_n176 ) , .ZN( u2_u7_u1_n98 ) );
  AOI211_X1 u2_u7_u1_U34 (.B( u2_u7_u1_n162 ) , .A( u2_u7_u1_n163 ) , .C2( u2_u7_u1_n164 ) , .ZN( u2_u7_u1_n165 ) , .C1( u2_u7_u1_n171 ) );
  AOI21_X1 u2_u7_u1_U35 (.A( u2_u7_u1_n160 ) , .B2( u2_u7_u1_n161 ) , .ZN( u2_u7_u1_n162 ) , .B1( u2_u7_u1_n182 ) );
  OR2_X1 u2_u7_u1_U36 (.A2( u2_u7_u1_n157 ) , .A1( u2_u7_u1_n158 ) , .ZN( u2_u7_u1_n163 ) );
  NAND2_X1 u2_u7_u1_U37 (.A1( u2_u7_u1_n128 ) , .ZN( u2_u7_u1_n146 ) , .A2( u2_u7_u1_n160 ) );
  NAND2_X1 u2_u7_u1_U38 (.A2( u2_u7_u1_n112 ) , .ZN( u2_u7_u1_n139 ) , .A1( u2_u7_u1_n152 ) );
  NAND2_X1 u2_u7_u1_U39 (.A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n156 ) , .A2( u2_u7_u1_n99 ) );
  AOI221_X1 u2_u7_u1_U4 (.A( u2_u7_u1_n138 ) , .C2( u2_u7_u1_n139 ) , .C1( u2_u7_u1_n140 ) , .B2( u2_u7_u1_n141 ) , .ZN( u2_u7_u1_n142 ) , .B1( u2_u7_u1_n175 ) );
  AOI221_X1 u2_u7_u1_U40 (.B1( u2_u7_u1_n140 ) , .ZN( u2_u7_u1_n167 ) , .B2( u2_u7_u1_n172 ) , .C2( u2_u7_u1_n175 ) , .C1( u2_u7_u1_n178 ) , .A( u2_u7_u1_n188 ) );
  INV_X1 u2_u7_u1_U41 (.ZN( u2_u7_u1_n188 ) , .A( u2_u7_u1_n97 ) );
  AOI211_X1 u2_u7_u1_U42 (.A( u2_u7_u1_n118 ) , .C1( u2_u7_u1_n132 ) , .C2( u2_u7_u1_n139 ) , .B( u2_u7_u1_n96 ) , .ZN( u2_u7_u1_n97 ) );
  AOI21_X1 u2_u7_u1_U43 (.B2( u2_u7_u1_n121 ) , .B1( u2_u7_u1_n135 ) , .A( u2_u7_u1_n152 ) , .ZN( u2_u7_u1_n96 ) );
  NOR2_X1 u2_u7_u1_U44 (.ZN( u2_u7_u1_n117 ) , .A1( u2_u7_u1_n121 ) , .A2( u2_u7_u1_n160 ) );
  OAI21_X1 u2_u7_u1_U45 (.B2( u2_u7_u1_n123 ) , .ZN( u2_u7_u1_n145 ) , .B1( u2_u7_u1_n160 ) , .A( u2_u7_u1_n185 ) );
  INV_X1 u2_u7_u1_U46 (.A( u2_u7_u1_n122 ) , .ZN( u2_u7_u1_n185 ) );
  AOI21_X1 u2_u7_u1_U47 (.B2( u2_u7_u1_n120 ) , .B1( u2_u7_u1_n121 ) , .ZN( u2_u7_u1_n122 ) , .A( u2_u7_u1_n128 ) );
  AOI21_X1 u2_u7_u1_U48 (.A( u2_u7_u1_n128 ) , .B2( u2_u7_u1_n129 ) , .ZN( u2_u7_u1_n130 ) , .B1( u2_u7_u1_n150 ) );
  NAND2_X1 u2_u7_u1_U49 (.ZN( u2_u7_u1_n112 ) , .A1( u2_u7_u1_n169 ) , .A2( u2_u7_u1_n170 ) );
  AOI211_X1 u2_u7_u1_U5 (.ZN( u2_u7_u1_n124 ) , .A( u2_u7_u1_n138 ) , .C2( u2_u7_u1_n139 ) , .B( u2_u7_u1_n145 ) , .C1( u2_u7_u1_n147 ) );
  NAND2_X1 u2_u7_u1_U50 (.ZN( u2_u7_u1_n129 ) , .A2( u2_u7_u1_n95 ) , .A1( u2_u7_u1_n98 ) );
  NAND2_X1 u2_u7_u1_U51 (.A1( u2_u7_u1_n102 ) , .ZN( u2_u7_u1_n154 ) , .A2( u2_u7_u1_n99 ) );
  NAND2_X1 u2_u7_u1_U52 (.A2( u2_u7_u1_n100 ) , .ZN( u2_u7_u1_n135 ) , .A1( u2_u7_u1_n99 ) );
  AOI21_X1 u2_u7_u1_U53 (.A( u2_u7_u1_n152 ) , .B2( u2_u7_u1_n153 ) , .B1( u2_u7_u1_n154 ) , .ZN( u2_u7_u1_n158 ) );
  INV_X1 u2_u7_u1_U54 (.A( u2_u7_u1_n160 ) , .ZN( u2_u7_u1_n175 ) );
  NAND2_X1 u2_u7_u1_U55 (.A1( u2_u7_u1_n100 ) , .ZN( u2_u7_u1_n116 ) , .A2( u2_u7_u1_n95 ) );
  NAND2_X1 u2_u7_u1_U56 (.A1( u2_u7_u1_n102 ) , .ZN( u2_u7_u1_n131 ) , .A2( u2_u7_u1_n95 ) );
  NAND2_X1 u2_u7_u1_U57 (.A2( u2_u7_u1_n104 ) , .ZN( u2_u7_u1_n121 ) , .A1( u2_u7_u1_n98 ) );
  NAND2_X1 u2_u7_u1_U58 (.A1( u2_u7_u1_n103 ) , .ZN( u2_u7_u1_n153 ) , .A2( u2_u7_u1_n98 ) );
  NAND2_X1 u2_u7_u1_U59 (.A2( u2_u7_u1_n104 ) , .A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n133 ) );
  AOI22_X1 u2_u7_u1_U6 (.B2( u2_u7_u1_n113 ) , .A2( u2_u7_u1_n114 ) , .ZN( u2_u7_u1_n125 ) , .A1( u2_u7_u1_n171 ) , .B1( u2_u7_u1_n173 ) );
  NAND2_X1 u2_u7_u1_U60 (.ZN( u2_u7_u1_n150 ) , .A2( u2_u7_u1_n98 ) , .A1( u2_u7_u1_n99 ) );
  NAND2_X1 u2_u7_u1_U61 (.A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n155 ) , .A2( u2_u7_u1_n95 ) );
  OAI21_X1 u2_u7_u1_U62 (.ZN( u2_u7_u1_n109 ) , .B1( u2_u7_u1_n129 ) , .B2( u2_u7_u1_n160 ) , .A( u2_u7_u1_n167 ) );
  NAND2_X1 u2_u7_u1_U63 (.A2( u2_u7_u1_n100 ) , .A1( u2_u7_u1_n103 ) , .ZN( u2_u7_u1_n120 ) );
  NAND2_X1 u2_u7_u1_U64 (.A1( u2_u7_u1_n102 ) , .A2( u2_u7_u1_n104 ) , .ZN( u2_u7_u1_n115 ) );
  NAND2_X1 u2_u7_u1_U65 (.A2( u2_u7_u1_n100 ) , .A1( u2_u7_u1_n104 ) , .ZN( u2_u7_u1_n151 ) );
  NAND2_X1 u2_u7_u1_U66 (.A2( u2_u7_u1_n103 ) , .A1( u2_u7_u1_n105 ) , .ZN( u2_u7_u1_n161 ) );
  INV_X1 u2_u7_u1_U67 (.A( u2_u7_u1_n152 ) , .ZN( u2_u7_u1_n173 ) );
  INV_X1 u2_u7_u1_U68 (.A( u2_u7_u1_n128 ) , .ZN( u2_u7_u1_n172 ) );
  NAND2_X1 u2_u7_u1_U69 (.A2( u2_u7_u1_n102 ) , .A1( u2_u7_u1_n103 ) , .ZN( u2_u7_u1_n123 ) );
  NAND2_X1 u2_u7_u1_U7 (.ZN( u2_u7_u1_n114 ) , .A1( u2_u7_u1_n134 ) , .A2( u2_u7_u1_n156 ) );
  NOR2_X1 u2_u7_u1_U70 (.A2( u2_u7_X_7 ) , .A1( u2_u7_X_8 ) , .ZN( u2_u7_u1_n95 ) );
  NOR2_X1 u2_u7_u1_U71 (.A1( u2_u7_X_12 ) , .A2( u2_u7_X_9 ) , .ZN( u2_u7_u1_n100 ) );
  NOR2_X1 u2_u7_u1_U72 (.A2( u2_u7_X_8 ) , .A1( u2_u7_u1_n177 ) , .ZN( u2_u7_u1_n99 ) );
  NOR2_X1 u2_u7_u1_U73 (.A2( u2_u7_X_12 ) , .ZN( u2_u7_u1_n102 ) , .A1( u2_u7_u1_n176 ) );
  NOR2_X1 u2_u7_u1_U74 (.A2( u2_u7_X_9 ) , .ZN( u2_u7_u1_n105 ) , .A1( u2_u7_u1_n168 ) );
  NAND2_X1 u2_u7_u1_U75 (.A1( u2_u7_X_10 ) , .ZN( u2_u7_u1_n160 ) , .A2( u2_u7_u1_n169 ) );
  NAND2_X1 u2_u7_u1_U76 (.A2( u2_u7_X_10 ) , .A1( u2_u7_X_11 ) , .ZN( u2_u7_u1_n152 ) );
  NAND2_X1 u2_u7_u1_U77 (.A1( u2_u7_X_11 ) , .ZN( u2_u7_u1_n128 ) , .A2( u2_u7_u1_n170 ) );
  AND2_X1 u2_u7_u1_U78 (.A2( u2_u7_X_7 ) , .A1( u2_u7_X_8 ) , .ZN( u2_u7_u1_n104 ) );
  AND2_X1 u2_u7_u1_U79 (.A1( u2_u7_X_8 ) , .ZN( u2_u7_u1_n103 ) , .A2( u2_u7_u1_n177 ) );
  NOR2_X1 u2_u7_u1_U8 (.A1( u2_u7_u1_n112 ) , .A2( u2_u7_u1_n116 ) , .ZN( u2_u7_u1_n118 ) );
  INV_X1 u2_u7_u1_U80 (.A( u2_u7_X_10 ) , .ZN( u2_u7_u1_n170 ) );
  INV_X1 u2_u7_u1_U81 (.A( u2_u7_X_9 ) , .ZN( u2_u7_u1_n176 ) );
  INV_X1 u2_u7_u1_U82 (.A( u2_u7_X_11 ) , .ZN( u2_u7_u1_n169 ) );
  INV_X1 u2_u7_u1_U83 (.A( u2_u7_X_12 ) , .ZN( u2_u7_u1_n168 ) );
  INV_X1 u2_u7_u1_U84 (.A( u2_u7_X_7 ) , .ZN( u2_u7_u1_n177 ) );
  NAND4_X1 u2_u7_u1_U85 (.ZN( u2_out7_28 ) , .A4( u2_u7_u1_n124 ) , .A3( u2_u7_u1_n125 ) , .A2( u2_u7_u1_n126 ) , .A1( u2_u7_u1_n127 ) );
  OAI21_X1 u2_u7_u1_U86 (.ZN( u2_u7_u1_n127 ) , .B2( u2_u7_u1_n139 ) , .B1( u2_u7_u1_n175 ) , .A( u2_u7_u1_n183 ) );
  OAI21_X1 u2_u7_u1_U87 (.ZN( u2_u7_u1_n126 ) , .B2( u2_u7_u1_n140 ) , .A( u2_u7_u1_n146 ) , .B1( u2_u7_u1_n178 ) );
  NAND4_X1 u2_u7_u1_U88 (.ZN( u2_out7_18 ) , .A4( u2_u7_u1_n165 ) , .A3( u2_u7_u1_n166 ) , .A1( u2_u7_u1_n167 ) , .A2( u2_u7_u1_n186 ) );
  AOI22_X1 u2_u7_u1_U89 (.B2( u2_u7_u1_n146 ) , .B1( u2_u7_u1_n147 ) , .A2( u2_u7_u1_n148 ) , .ZN( u2_u7_u1_n166 ) , .A1( u2_u7_u1_n172 ) );
  OAI21_X1 u2_u7_u1_U9 (.ZN( u2_u7_u1_n101 ) , .B1( u2_u7_u1_n141 ) , .A( u2_u7_u1_n146 ) , .B2( u2_u7_u1_n183 ) );
  INV_X1 u2_u7_u1_U90 (.A( u2_u7_u1_n145 ) , .ZN( u2_u7_u1_n186 ) );
  NAND4_X1 u2_u7_u1_U91 (.ZN( u2_out7_2 ) , .A4( u2_u7_u1_n142 ) , .A3( u2_u7_u1_n143 ) , .A2( u2_u7_u1_n144 ) , .A1( u2_u7_u1_n179 ) );
  OAI21_X1 u2_u7_u1_U92 (.B2( u2_u7_u1_n132 ) , .ZN( u2_u7_u1_n144 ) , .A( u2_u7_u1_n146 ) , .B1( u2_u7_u1_n180 ) );
  INV_X1 u2_u7_u1_U93 (.A( u2_u7_u1_n130 ) , .ZN( u2_u7_u1_n179 ) );
  OR4_X1 u2_u7_u1_U94 (.ZN( u2_out7_13 ) , .A4( u2_u7_u1_n108 ) , .A3( u2_u7_u1_n109 ) , .A2( u2_u7_u1_n110 ) , .A1( u2_u7_u1_n111 ) );
  AOI21_X1 u2_u7_u1_U95 (.ZN( u2_u7_u1_n111 ) , .A( u2_u7_u1_n128 ) , .B2( u2_u7_u1_n131 ) , .B1( u2_u7_u1_n135 ) );
  AOI21_X1 u2_u7_u1_U96 (.ZN( u2_u7_u1_n110 ) , .A( u2_u7_u1_n116 ) , .B1( u2_u7_u1_n152 ) , .B2( u2_u7_u1_n160 ) );
  NAND3_X1 u2_u7_u1_U97 (.A3( u2_u7_u1_n149 ) , .A2( u2_u7_u1_n150 ) , .A1( u2_u7_u1_n151 ) , .ZN( u2_u7_u1_n164 ) );
  NAND3_X1 u2_u7_u1_U98 (.A3( u2_u7_u1_n134 ) , .A2( u2_u7_u1_n135 ) , .ZN( u2_u7_u1_n136 ) , .A1( u2_u7_u1_n151 ) );
  NAND3_X1 u2_u7_u1_U99 (.A1( u2_u7_u1_n133 ) , .ZN( u2_u7_u1_n137 ) , .A2( u2_u7_u1_n154 ) , .A3( u2_u7_u1_n181 ) );
  OAI22_X1 u2_u7_u2_U10 (.ZN( u2_u7_u2_n109 ) , .A2( u2_u7_u2_n113 ) , .B2( u2_u7_u2_n133 ) , .B1( u2_u7_u2_n167 ) , .A1( u2_u7_u2_n168 ) );
  NAND3_X1 u2_u7_u2_U100 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n104 ) , .A3( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n98 ) );
  OAI22_X1 u2_u7_u2_U11 (.B1( u2_u7_u2_n151 ) , .A2( u2_u7_u2_n152 ) , .A1( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n160 ) , .B2( u2_u7_u2_n168 ) );
  NOR3_X1 u2_u7_u2_U12 (.A1( u2_u7_u2_n150 ) , .ZN( u2_u7_u2_n151 ) , .A3( u2_u7_u2_n175 ) , .A2( u2_u7_u2_n188 ) );
  AOI21_X1 u2_u7_u2_U13 (.ZN( u2_u7_u2_n144 ) , .B2( u2_u7_u2_n155 ) , .A( u2_u7_u2_n172 ) , .B1( u2_u7_u2_n185 ) );
  AOI21_X1 u2_u7_u2_U14 (.B2( u2_u7_u2_n143 ) , .ZN( u2_u7_u2_n145 ) , .B1( u2_u7_u2_n152 ) , .A( u2_u7_u2_n171 ) );
  AOI21_X1 u2_u7_u2_U15 (.B2( u2_u7_u2_n120 ) , .B1( u2_u7_u2_n121 ) , .ZN( u2_u7_u2_n126 ) , .A( u2_u7_u2_n167 ) );
  INV_X1 u2_u7_u2_U16 (.A( u2_u7_u2_n156 ) , .ZN( u2_u7_u2_n171 ) );
  INV_X1 u2_u7_u2_U17 (.A( u2_u7_u2_n120 ) , .ZN( u2_u7_u2_n188 ) );
  NAND2_X1 u2_u7_u2_U18 (.A2( u2_u7_u2_n122 ) , .ZN( u2_u7_u2_n150 ) , .A1( u2_u7_u2_n152 ) );
  INV_X1 u2_u7_u2_U19 (.A( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n170 ) );
  INV_X1 u2_u7_u2_U20 (.A( u2_u7_u2_n137 ) , .ZN( u2_u7_u2_n173 ) );
  NAND2_X1 u2_u7_u2_U21 (.A1( u2_u7_u2_n132 ) , .A2( u2_u7_u2_n139 ) , .ZN( u2_u7_u2_n157 ) );
  INV_X1 u2_u7_u2_U22 (.A( u2_u7_u2_n113 ) , .ZN( u2_u7_u2_n178 ) );
  INV_X1 u2_u7_u2_U23 (.A( u2_u7_u2_n139 ) , .ZN( u2_u7_u2_n175 ) );
  INV_X1 u2_u7_u2_U24 (.A( u2_u7_u2_n155 ) , .ZN( u2_u7_u2_n181 ) );
  INV_X1 u2_u7_u2_U25 (.A( u2_u7_u2_n119 ) , .ZN( u2_u7_u2_n177 ) );
  INV_X1 u2_u7_u2_U26 (.A( u2_u7_u2_n116 ) , .ZN( u2_u7_u2_n180 ) );
  INV_X1 u2_u7_u2_U27 (.A( u2_u7_u2_n131 ) , .ZN( u2_u7_u2_n179 ) );
  INV_X1 u2_u7_u2_U28 (.A( u2_u7_u2_n154 ) , .ZN( u2_u7_u2_n176 ) );
  NAND2_X1 u2_u7_u2_U29 (.A2( u2_u7_u2_n116 ) , .A1( u2_u7_u2_n117 ) , .ZN( u2_u7_u2_n118 ) );
  NOR2_X1 u2_u7_u2_U3 (.ZN( u2_u7_u2_n121 ) , .A2( u2_u7_u2_n177 ) , .A1( u2_u7_u2_n180 ) );
  INV_X1 u2_u7_u2_U30 (.A( u2_u7_u2_n132 ) , .ZN( u2_u7_u2_n182 ) );
  INV_X1 u2_u7_u2_U31 (.A( u2_u7_u2_n158 ) , .ZN( u2_u7_u2_n183 ) );
  OAI21_X1 u2_u7_u2_U32 (.A( u2_u7_u2_n156 ) , .B1( u2_u7_u2_n157 ) , .ZN( u2_u7_u2_n158 ) , .B2( u2_u7_u2_n179 ) );
  NOR2_X1 u2_u7_u2_U33 (.ZN( u2_u7_u2_n156 ) , .A1( u2_u7_u2_n166 ) , .A2( u2_u7_u2_n169 ) );
  NOR2_X1 u2_u7_u2_U34 (.A2( u2_u7_u2_n114 ) , .ZN( u2_u7_u2_n137 ) , .A1( u2_u7_u2_n140 ) );
  NOR2_X1 u2_u7_u2_U35 (.A2( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n153 ) , .A1( u2_u7_u2_n156 ) );
  AOI211_X1 u2_u7_u2_U36 (.ZN( u2_u7_u2_n130 ) , .C1( u2_u7_u2_n138 ) , .C2( u2_u7_u2_n179 ) , .B( u2_u7_u2_n96 ) , .A( u2_u7_u2_n97 ) );
  OAI22_X1 u2_u7_u2_U37 (.B1( u2_u7_u2_n133 ) , .A2( u2_u7_u2_n137 ) , .A1( u2_u7_u2_n152 ) , .B2( u2_u7_u2_n168 ) , .ZN( u2_u7_u2_n97 ) );
  OAI221_X1 u2_u7_u2_U38 (.B1( u2_u7_u2_n113 ) , .C1( u2_u7_u2_n132 ) , .A( u2_u7_u2_n149 ) , .B2( u2_u7_u2_n171 ) , .C2( u2_u7_u2_n172 ) , .ZN( u2_u7_u2_n96 ) );
  OAI221_X1 u2_u7_u2_U39 (.A( u2_u7_u2_n115 ) , .C2( u2_u7_u2_n123 ) , .B2( u2_u7_u2_n143 ) , .B1( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n163 ) , .C1( u2_u7_u2_n168 ) );
  INV_X1 u2_u7_u2_U4 (.A( u2_u7_u2_n134 ) , .ZN( u2_u7_u2_n185 ) );
  OAI21_X1 u2_u7_u2_U40 (.A( u2_u7_u2_n114 ) , .ZN( u2_u7_u2_n115 ) , .B1( u2_u7_u2_n176 ) , .B2( u2_u7_u2_n178 ) );
  OAI221_X1 u2_u7_u2_U41 (.A( u2_u7_u2_n135 ) , .B2( u2_u7_u2_n136 ) , .B1( u2_u7_u2_n137 ) , .ZN( u2_u7_u2_n162 ) , .C2( u2_u7_u2_n167 ) , .C1( u2_u7_u2_n185 ) );
  AND3_X1 u2_u7_u2_U42 (.A3( u2_u7_u2_n131 ) , .A2( u2_u7_u2_n132 ) , .A1( u2_u7_u2_n133 ) , .ZN( u2_u7_u2_n136 ) );
  AOI22_X1 u2_u7_u2_U43 (.ZN( u2_u7_u2_n135 ) , .B1( u2_u7_u2_n140 ) , .A1( u2_u7_u2_n156 ) , .B2( u2_u7_u2_n180 ) , .A2( u2_u7_u2_n188 ) );
  AOI21_X1 u2_u7_u2_U44 (.ZN( u2_u7_u2_n149 ) , .B1( u2_u7_u2_n173 ) , .B2( u2_u7_u2_n188 ) , .A( u2_u7_u2_n95 ) );
  AND3_X1 u2_u7_u2_U45 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n104 ) , .A3( u2_u7_u2_n156 ) , .ZN( u2_u7_u2_n95 ) );
  OAI21_X1 u2_u7_u2_U46 (.A( u2_u7_u2_n101 ) , .B2( u2_u7_u2_n121 ) , .B1( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n164 ) );
  NAND2_X1 u2_u7_u2_U47 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n107 ) , .ZN( u2_u7_u2_n155 ) );
  NAND2_X1 u2_u7_u2_U48 (.A2( u2_u7_u2_n105 ) , .A1( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n143 ) );
  NAND2_X1 u2_u7_u2_U49 (.A1( u2_u7_u2_n104 ) , .A2( u2_u7_u2_n106 ) , .ZN( u2_u7_u2_n152 ) );
  INV_X1 u2_u7_u2_U5 (.A( u2_u7_u2_n150 ) , .ZN( u2_u7_u2_n184 ) );
  NAND2_X1 u2_u7_u2_U50 (.A1( u2_u7_u2_n100 ) , .A2( u2_u7_u2_n105 ) , .ZN( u2_u7_u2_n132 ) );
  INV_X1 u2_u7_u2_U51 (.A( u2_u7_u2_n140 ) , .ZN( u2_u7_u2_n168 ) );
  INV_X1 u2_u7_u2_U52 (.A( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n167 ) );
  OAI21_X1 u2_u7_u2_U53 (.A( u2_u7_u2_n141 ) , .B2( u2_u7_u2_n142 ) , .ZN( u2_u7_u2_n146 ) , .B1( u2_u7_u2_n153 ) );
  OAI21_X1 u2_u7_u2_U54 (.A( u2_u7_u2_n140 ) , .ZN( u2_u7_u2_n141 ) , .B1( u2_u7_u2_n176 ) , .B2( u2_u7_u2_n177 ) );
  NOR3_X1 u2_u7_u2_U55 (.ZN( u2_u7_u2_n142 ) , .A3( u2_u7_u2_n175 ) , .A2( u2_u7_u2_n178 ) , .A1( u2_u7_u2_n181 ) );
  INV_X1 u2_u7_u2_U56 (.ZN( u2_u7_u2_n187 ) , .A( u2_u7_u2_n99 ) );
  OAI21_X1 u2_u7_u2_U57 (.B1( u2_u7_u2_n137 ) , .B2( u2_u7_u2_n143 ) , .A( u2_u7_u2_n98 ) , .ZN( u2_u7_u2_n99 ) );
  NAND2_X1 u2_u7_u2_U58 (.A1( u2_u7_u2_n102 ) , .A2( u2_u7_u2_n106 ) , .ZN( u2_u7_u2_n113 ) );
  NAND2_X1 u2_u7_u2_U59 (.A1( u2_u7_u2_n106 ) , .A2( u2_u7_u2_n107 ) , .ZN( u2_u7_u2_n131 ) );
  NOR4_X1 u2_u7_u2_U6 (.A4( u2_u7_u2_n124 ) , .A3( u2_u7_u2_n125 ) , .A2( u2_u7_u2_n126 ) , .A1( u2_u7_u2_n127 ) , .ZN( u2_u7_u2_n128 ) );
  NAND2_X1 u2_u7_u2_U60 (.A1( u2_u7_u2_n103 ) , .A2( u2_u7_u2_n107 ) , .ZN( u2_u7_u2_n139 ) );
  NAND2_X1 u2_u7_u2_U61 (.A1( u2_u7_u2_n103 ) , .A2( u2_u7_u2_n105 ) , .ZN( u2_u7_u2_n133 ) );
  NAND2_X1 u2_u7_u2_U62 (.A1( u2_u7_u2_n102 ) , .A2( u2_u7_u2_n103 ) , .ZN( u2_u7_u2_n154 ) );
  NAND2_X1 u2_u7_u2_U63 (.A2( u2_u7_u2_n103 ) , .A1( u2_u7_u2_n104 ) , .ZN( u2_u7_u2_n119 ) );
  NAND2_X1 u2_u7_u2_U64 (.A2( u2_u7_u2_n107 ) , .A1( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n123 ) );
  NAND2_X1 u2_u7_u2_U65 (.A1( u2_u7_u2_n104 ) , .A2( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n122 ) );
  INV_X1 u2_u7_u2_U66 (.A( u2_u7_u2_n114 ) , .ZN( u2_u7_u2_n172 ) );
  NAND2_X1 u2_u7_u2_U67 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n102 ) , .ZN( u2_u7_u2_n116 ) );
  NAND2_X1 u2_u7_u2_U68 (.A1( u2_u7_u2_n102 ) , .A2( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n120 ) );
  NAND2_X1 u2_u7_u2_U69 (.A2( u2_u7_u2_n105 ) , .A1( u2_u7_u2_n106 ) , .ZN( u2_u7_u2_n117 ) );
  AOI21_X1 u2_u7_u2_U7 (.B2( u2_u7_u2_n119 ) , .ZN( u2_u7_u2_n127 ) , .A( u2_u7_u2_n137 ) , .B1( u2_u7_u2_n155 ) );
  NOR2_X1 u2_u7_u2_U70 (.A2( u2_u7_X_16 ) , .ZN( u2_u7_u2_n140 ) , .A1( u2_u7_u2_n166 ) );
  NOR2_X1 u2_u7_u2_U71 (.A2( u2_u7_X_13 ) , .A1( u2_u7_X_14 ) , .ZN( u2_u7_u2_n100 ) );
  NOR2_X1 u2_u7_u2_U72 (.A2( u2_u7_X_16 ) , .A1( u2_u7_X_17 ) , .ZN( u2_u7_u2_n138 ) );
  NOR2_X1 u2_u7_u2_U73 (.A2( u2_u7_X_15 ) , .A1( u2_u7_X_18 ) , .ZN( u2_u7_u2_n104 ) );
  NOR2_X1 u2_u7_u2_U74 (.A2( u2_u7_X_14 ) , .ZN( u2_u7_u2_n103 ) , .A1( u2_u7_u2_n174 ) );
  NOR2_X1 u2_u7_u2_U75 (.A2( u2_u7_X_15 ) , .ZN( u2_u7_u2_n102 ) , .A1( u2_u7_u2_n165 ) );
  NOR2_X1 u2_u7_u2_U76 (.A2( u2_u7_X_17 ) , .ZN( u2_u7_u2_n114 ) , .A1( u2_u7_u2_n169 ) );
  AND2_X1 u2_u7_u2_U77 (.A1( u2_u7_X_15 ) , .ZN( u2_u7_u2_n105 ) , .A2( u2_u7_u2_n165 ) );
  AND2_X1 u2_u7_u2_U78 (.A2( u2_u7_X_15 ) , .A1( u2_u7_X_18 ) , .ZN( u2_u7_u2_n107 ) );
  AND2_X1 u2_u7_u2_U79 (.A1( u2_u7_X_14 ) , .ZN( u2_u7_u2_n106 ) , .A2( u2_u7_u2_n174 ) );
  AOI21_X1 u2_u7_u2_U8 (.ZN( u2_u7_u2_n124 ) , .B1( u2_u7_u2_n131 ) , .B2( u2_u7_u2_n143 ) , .A( u2_u7_u2_n172 ) );
  AND2_X1 u2_u7_u2_U80 (.A1( u2_u7_X_13 ) , .A2( u2_u7_X_14 ) , .ZN( u2_u7_u2_n108 ) );
  INV_X1 u2_u7_u2_U81 (.A( u2_u7_X_16 ) , .ZN( u2_u7_u2_n169 ) );
  INV_X1 u2_u7_u2_U82 (.A( u2_u7_X_17 ) , .ZN( u2_u7_u2_n166 ) );
  INV_X1 u2_u7_u2_U83 (.A( u2_u7_X_13 ) , .ZN( u2_u7_u2_n174 ) );
  INV_X1 u2_u7_u2_U84 (.A( u2_u7_X_18 ) , .ZN( u2_u7_u2_n165 ) );
  NAND4_X1 u2_u7_u2_U85 (.ZN( u2_out7_24 ) , .A4( u2_u7_u2_n111 ) , .A3( u2_u7_u2_n112 ) , .A1( u2_u7_u2_n130 ) , .A2( u2_u7_u2_n187 ) );
  AOI221_X1 u2_u7_u2_U86 (.A( u2_u7_u2_n109 ) , .B1( u2_u7_u2_n110 ) , .ZN( u2_u7_u2_n111 ) , .C1( u2_u7_u2_n134 ) , .C2( u2_u7_u2_n170 ) , .B2( u2_u7_u2_n173 ) );
  AOI21_X1 u2_u7_u2_U87 (.ZN( u2_u7_u2_n112 ) , .B2( u2_u7_u2_n156 ) , .A( u2_u7_u2_n164 ) , .B1( u2_u7_u2_n181 ) );
  NAND4_X1 u2_u7_u2_U88 (.ZN( u2_out7_16 ) , .A4( u2_u7_u2_n128 ) , .A3( u2_u7_u2_n129 ) , .A1( u2_u7_u2_n130 ) , .A2( u2_u7_u2_n186 ) );
  AOI22_X1 u2_u7_u2_U89 (.A2( u2_u7_u2_n118 ) , .ZN( u2_u7_u2_n129 ) , .A1( u2_u7_u2_n140 ) , .B1( u2_u7_u2_n157 ) , .B2( u2_u7_u2_n170 ) );
  AOI21_X1 u2_u7_u2_U9 (.B2( u2_u7_u2_n123 ) , .ZN( u2_u7_u2_n125 ) , .A( u2_u7_u2_n171 ) , .B1( u2_u7_u2_n184 ) );
  INV_X1 u2_u7_u2_U90 (.A( u2_u7_u2_n163 ) , .ZN( u2_u7_u2_n186 ) );
  NAND4_X1 u2_u7_u2_U91 (.ZN( u2_out7_30 ) , .A4( u2_u7_u2_n147 ) , .A3( u2_u7_u2_n148 ) , .A2( u2_u7_u2_n149 ) , .A1( u2_u7_u2_n187 ) );
  NOR3_X1 u2_u7_u2_U92 (.A3( u2_u7_u2_n144 ) , .A2( u2_u7_u2_n145 ) , .A1( u2_u7_u2_n146 ) , .ZN( u2_u7_u2_n147 ) );
  AOI21_X1 u2_u7_u2_U93 (.B2( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n148 ) , .A( u2_u7_u2_n162 ) , .B1( u2_u7_u2_n182 ) );
  OR4_X1 u2_u7_u2_U94 (.ZN( u2_out7_6 ) , .A4( u2_u7_u2_n161 ) , .A3( u2_u7_u2_n162 ) , .A2( u2_u7_u2_n163 ) , .A1( u2_u7_u2_n164 ) );
  OR3_X1 u2_u7_u2_U95 (.A2( u2_u7_u2_n159 ) , .A1( u2_u7_u2_n160 ) , .ZN( u2_u7_u2_n161 ) , .A3( u2_u7_u2_n183 ) );
  AOI21_X1 u2_u7_u2_U96 (.B2( u2_u7_u2_n154 ) , .B1( u2_u7_u2_n155 ) , .ZN( u2_u7_u2_n159 ) , .A( u2_u7_u2_n167 ) );
  NAND3_X1 u2_u7_u2_U97 (.A2( u2_u7_u2_n117 ) , .A1( u2_u7_u2_n122 ) , .A3( u2_u7_u2_n123 ) , .ZN( u2_u7_u2_n134 ) );
  NAND3_X1 u2_u7_u2_U98 (.ZN( u2_u7_u2_n110 ) , .A2( u2_u7_u2_n131 ) , .A3( u2_u7_u2_n139 ) , .A1( u2_u7_u2_n154 ) );
  NAND3_X1 u2_u7_u2_U99 (.A2( u2_u7_u2_n100 ) , .ZN( u2_u7_u2_n101 ) , .A1( u2_u7_u2_n104 ) , .A3( u2_u7_u2_n114 ) );
  OAI22_X1 u2_u7_u3_U10 (.B1( u2_u7_u3_n113 ) , .A2( u2_u7_u3_n135 ) , .A1( u2_u7_u3_n150 ) , .B2( u2_u7_u3_n164 ) , .ZN( u2_u7_u3_n98 ) );
  OAI211_X1 u2_u7_u3_U11 (.B( u2_u7_u3_n106 ) , .ZN( u2_u7_u3_n119 ) , .C2( u2_u7_u3_n128 ) , .C1( u2_u7_u3_n167 ) , .A( u2_u7_u3_n181 ) );
  AOI221_X1 u2_u7_u3_U12 (.C1( u2_u7_u3_n105 ) , .ZN( u2_u7_u3_n106 ) , .A( u2_u7_u3_n131 ) , .B2( u2_u7_u3_n132 ) , .C2( u2_u7_u3_n133 ) , .B1( u2_u7_u3_n169 ) );
  INV_X1 u2_u7_u3_U13 (.ZN( u2_u7_u3_n181 ) , .A( u2_u7_u3_n98 ) );
  NAND2_X1 u2_u7_u3_U14 (.ZN( u2_u7_u3_n105 ) , .A2( u2_u7_u3_n130 ) , .A1( u2_u7_u3_n155 ) );
  AOI22_X1 u2_u7_u3_U15 (.B1( u2_u7_u3_n115 ) , .A2( u2_u7_u3_n116 ) , .ZN( u2_u7_u3_n123 ) , .B2( u2_u7_u3_n133 ) , .A1( u2_u7_u3_n169 ) );
  NAND2_X1 u2_u7_u3_U16 (.ZN( u2_u7_u3_n116 ) , .A2( u2_u7_u3_n151 ) , .A1( u2_u7_u3_n182 ) );
  NOR2_X1 u2_u7_u3_U17 (.ZN( u2_u7_u3_n126 ) , .A2( u2_u7_u3_n150 ) , .A1( u2_u7_u3_n164 ) );
  AOI21_X1 u2_u7_u3_U18 (.ZN( u2_u7_u3_n112 ) , .B2( u2_u7_u3_n146 ) , .B1( u2_u7_u3_n155 ) , .A( u2_u7_u3_n167 ) );
  NAND2_X1 u2_u7_u3_U19 (.A1( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n142 ) , .A2( u2_u7_u3_n164 ) );
  NAND2_X1 u2_u7_u3_U20 (.ZN( u2_u7_u3_n132 ) , .A2( u2_u7_u3_n152 ) , .A1( u2_u7_u3_n156 ) );
  AND2_X1 u2_u7_u3_U21 (.A2( u2_u7_u3_n113 ) , .A1( u2_u7_u3_n114 ) , .ZN( u2_u7_u3_n151 ) );
  INV_X1 u2_u7_u3_U22 (.A( u2_u7_u3_n133 ) , .ZN( u2_u7_u3_n165 ) );
  INV_X1 u2_u7_u3_U23 (.A( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n170 ) );
  NAND2_X1 u2_u7_u3_U24 (.A1( u2_u7_u3_n107 ) , .A2( u2_u7_u3_n108 ) , .ZN( u2_u7_u3_n140 ) );
  NAND2_X1 u2_u7_u3_U25 (.ZN( u2_u7_u3_n117 ) , .A1( u2_u7_u3_n124 ) , .A2( u2_u7_u3_n148 ) );
  NAND2_X1 u2_u7_u3_U26 (.ZN( u2_u7_u3_n143 ) , .A1( u2_u7_u3_n165 ) , .A2( u2_u7_u3_n167 ) );
  INV_X1 u2_u7_u3_U27 (.A( u2_u7_u3_n130 ) , .ZN( u2_u7_u3_n177 ) );
  INV_X1 u2_u7_u3_U28 (.A( u2_u7_u3_n128 ) , .ZN( u2_u7_u3_n176 ) );
  INV_X1 u2_u7_u3_U29 (.A( u2_u7_u3_n155 ) , .ZN( u2_u7_u3_n174 ) );
  INV_X1 u2_u7_u3_U3 (.A( u2_u7_u3_n129 ) , .ZN( u2_u7_u3_n183 ) );
  INV_X1 u2_u7_u3_U30 (.A( u2_u7_u3_n139 ) , .ZN( u2_u7_u3_n185 ) );
  NOR2_X1 u2_u7_u3_U31 (.ZN( u2_u7_u3_n135 ) , .A2( u2_u7_u3_n141 ) , .A1( u2_u7_u3_n169 ) );
  OAI222_X1 u2_u7_u3_U32 (.C2( u2_u7_u3_n107 ) , .A2( u2_u7_u3_n108 ) , .B1( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n138 ) , .B2( u2_u7_u3_n146 ) , .C1( u2_u7_u3_n154 ) , .A1( u2_u7_u3_n164 ) );
  NOR4_X1 u2_u7_u3_U33 (.A4( u2_u7_u3_n157 ) , .A3( u2_u7_u3_n158 ) , .A2( u2_u7_u3_n159 ) , .A1( u2_u7_u3_n160 ) , .ZN( u2_u7_u3_n161 ) );
  AOI21_X1 u2_u7_u3_U34 (.B2( u2_u7_u3_n152 ) , .B1( u2_u7_u3_n153 ) , .ZN( u2_u7_u3_n158 ) , .A( u2_u7_u3_n164 ) );
  AOI21_X1 u2_u7_u3_U35 (.A( u2_u7_u3_n154 ) , .B2( u2_u7_u3_n155 ) , .B1( u2_u7_u3_n156 ) , .ZN( u2_u7_u3_n157 ) );
  AOI21_X1 u2_u7_u3_U36 (.A( u2_u7_u3_n149 ) , .B2( u2_u7_u3_n150 ) , .B1( u2_u7_u3_n151 ) , .ZN( u2_u7_u3_n159 ) );
  AOI211_X1 u2_u7_u3_U37 (.ZN( u2_u7_u3_n109 ) , .A( u2_u7_u3_n119 ) , .C2( u2_u7_u3_n129 ) , .B( u2_u7_u3_n138 ) , .C1( u2_u7_u3_n141 ) );
  AOI211_X1 u2_u7_u3_U38 (.B( u2_u7_u3_n119 ) , .A( u2_u7_u3_n120 ) , .C2( u2_u7_u3_n121 ) , .ZN( u2_u7_u3_n122 ) , .C1( u2_u7_u3_n179 ) );
  INV_X1 u2_u7_u3_U39 (.A( u2_u7_u3_n156 ) , .ZN( u2_u7_u3_n179 ) );
  INV_X1 u2_u7_u3_U4 (.A( u2_u7_u3_n140 ) , .ZN( u2_u7_u3_n182 ) );
  OAI22_X1 u2_u7_u3_U40 (.B1( u2_u7_u3_n118 ) , .ZN( u2_u7_u3_n120 ) , .A1( u2_u7_u3_n135 ) , .B2( u2_u7_u3_n154 ) , .A2( u2_u7_u3_n178 ) );
  AND3_X1 u2_u7_u3_U41 (.ZN( u2_u7_u3_n118 ) , .A2( u2_u7_u3_n124 ) , .A1( u2_u7_u3_n144 ) , .A3( u2_u7_u3_n152 ) );
  INV_X1 u2_u7_u3_U42 (.A( u2_u7_u3_n121 ) , .ZN( u2_u7_u3_n164 ) );
  NAND2_X1 u2_u7_u3_U43 (.ZN( u2_u7_u3_n133 ) , .A1( u2_u7_u3_n154 ) , .A2( u2_u7_u3_n164 ) );
  OAI211_X1 u2_u7_u3_U44 (.B( u2_u7_u3_n127 ) , .ZN( u2_u7_u3_n139 ) , .C1( u2_u7_u3_n150 ) , .C2( u2_u7_u3_n154 ) , .A( u2_u7_u3_n184 ) );
  INV_X1 u2_u7_u3_U45 (.A( u2_u7_u3_n125 ) , .ZN( u2_u7_u3_n184 ) );
  AOI221_X1 u2_u7_u3_U46 (.A( u2_u7_u3_n126 ) , .ZN( u2_u7_u3_n127 ) , .C2( u2_u7_u3_n132 ) , .C1( u2_u7_u3_n169 ) , .B2( u2_u7_u3_n170 ) , .B1( u2_u7_u3_n174 ) );
  OAI22_X1 u2_u7_u3_U47 (.A1( u2_u7_u3_n124 ) , .ZN( u2_u7_u3_n125 ) , .B2( u2_u7_u3_n145 ) , .A2( u2_u7_u3_n165 ) , .B1( u2_u7_u3_n167 ) );
  NOR2_X1 u2_u7_u3_U48 (.A1( u2_u7_u3_n113 ) , .ZN( u2_u7_u3_n131 ) , .A2( u2_u7_u3_n154 ) );
  NAND2_X1 u2_u7_u3_U49 (.A1( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n150 ) , .A2( u2_u7_u3_n99 ) );
  INV_X1 u2_u7_u3_U5 (.A( u2_u7_u3_n117 ) , .ZN( u2_u7_u3_n178 ) );
  NAND2_X1 u2_u7_u3_U50 (.A2( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n155 ) , .A1( u2_u7_u3_n97 ) );
  INV_X1 u2_u7_u3_U51 (.A( u2_u7_u3_n141 ) , .ZN( u2_u7_u3_n167 ) );
  AOI21_X1 u2_u7_u3_U52 (.B2( u2_u7_u3_n114 ) , .B1( u2_u7_u3_n146 ) , .A( u2_u7_u3_n154 ) , .ZN( u2_u7_u3_n94 ) );
  AOI21_X1 u2_u7_u3_U53 (.ZN( u2_u7_u3_n110 ) , .B2( u2_u7_u3_n142 ) , .B1( u2_u7_u3_n186 ) , .A( u2_u7_u3_n95 ) );
  INV_X1 u2_u7_u3_U54 (.A( u2_u7_u3_n145 ) , .ZN( u2_u7_u3_n186 ) );
  AOI21_X1 u2_u7_u3_U55 (.B1( u2_u7_u3_n124 ) , .A( u2_u7_u3_n149 ) , .B2( u2_u7_u3_n155 ) , .ZN( u2_u7_u3_n95 ) );
  INV_X1 u2_u7_u3_U56 (.A( u2_u7_u3_n149 ) , .ZN( u2_u7_u3_n169 ) );
  NAND2_X1 u2_u7_u3_U57 (.ZN( u2_u7_u3_n124 ) , .A1( u2_u7_u3_n96 ) , .A2( u2_u7_u3_n97 ) );
  NAND2_X1 u2_u7_u3_U58 (.A2( u2_u7_u3_n100 ) , .ZN( u2_u7_u3_n146 ) , .A1( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U59 (.A1( u2_u7_u3_n101 ) , .ZN( u2_u7_u3_n145 ) , .A2( u2_u7_u3_n99 ) );
  AOI221_X1 u2_u7_u3_U6 (.A( u2_u7_u3_n131 ) , .C2( u2_u7_u3_n132 ) , .C1( u2_u7_u3_n133 ) , .ZN( u2_u7_u3_n134 ) , .B1( u2_u7_u3_n143 ) , .B2( u2_u7_u3_n177 ) );
  NAND2_X1 u2_u7_u3_U60 (.A1( u2_u7_u3_n100 ) , .ZN( u2_u7_u3_n156 ) , .A2( u2_u7_u3_n99 ) );
  NAND2_X1 u2_u7_u3_U61 (.A2( u2_u7_u3_n101 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n148 ) );
  NAND2_X1 u2_u7_u3_U62 (.A1( u2_u7_u3_n100 ) , .A2( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n128 ) );
  NAND2_X1 u2_u7_u3_U63 (.A2( u2_u7_u3_n101 ) , .A1( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n152 ) );
  NAND2_X1 u2_u7_u3_U64 (.A2( u2_u7_u3_n101 ) , .ZN( u2_u7_u3_n114 ) , .A1( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U65 (.ZN( u2_u7_u3_n107 ) , .A1( u2_u7_u3_n97 ) , .A2( u2_u7_u3_n99 ) );
  NAND2_X1 u2_u7_u3_U66 (.A2( u2_u7_u3_n100 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n113 ) );
  NAND2_X1 u2_u7_u3_U67 (.A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n153 ) , .A2( u2_u7_u3_n97 ) );
  NAND2_X1 u2_u7_u3_U68 (.A2( u2_u7_u3_n103 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n130 ) );
  NAND2_X1 u2_u7_u3_U69 (.A2( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n144 ) , .A1( u2_u7_u3_n96 ) );
  OAI22_X1 u2_u7_u3_U7 (.B2( u2_u7_u3_n147 ) , .A2( u2_u7_u3_n148 ) , .ZN( u2_u7_u3_n160 ) , .B1( u2_u7_u3_n165 ) , .A1( u2_u7_u3_n168 ) );
  NAND2_X1 u2_u7_u3_U70 (.A1( u2_u7_u3_n102 ) , .A2( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n108 ) );
  NOR2_X1 u2_u7_u3_U71 (.A2( u2_u7_X_19 ) , .A1( u2_u7_X_20 ) , .ZN( u2_u7_u3_n99 ) );
  NOR2_X1 u2_u7_u3_U72 (.A2( u2_u7_X_21 ) , .A1( u2_u7_X_24 ) , .ZN( u2_u7_u3_n103 ) );
  NOR2_X1 u2_u7_u3_U73 (.A2( u2_u7_X_24 ) , .A1( u2_u7_u3_n171 ) , .ZN( u2_u7_u3_n97 ) );
  NOR2_X1 u2_u7_u3_U74 (.A2( u2_u7_X_23 ) , .ZN( u2_u7_u3_n141 ) , .A1( u2_u7_u3_n166 ) );
  NOR2_X1 u2_u7_u3_U75 (.A2( u2_u7_X_19 ) , .A1( u2_u7_u3_n172 ) , .ZN( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U76 (.A1( u2_u7_X_22 ) , .A2( u2_u7_X_23 ) , .ZN( u2_u7_u3_n154 ) );
  NAND2_X1 u2_u7_u3_U77 (.A1( u2_u7_X_23 ) , .ZN( u2_u7_u3_n149 ) , .A2( u2_u7_u3_n166 ) );
  NOR2_X1 u2_u7_u3_U78 (.A2( u2_u7_X_22 ) , .A1( u2_u7_X_23 ) , .ZN( u2_u7_u3_n121 ) );
  AND2_X1 u2_u7_u3_U79 (.A1( u2_u7_X_24 ) , .ZN( u2_u7_u3_n101 ) , .A2( u2_u7_u3_n171 ) );
  AND3_X1 u2_u7_u3_U8 (.A3( u2_u7_u3_n144 ) , .A2( u2_u7_u3_n145 ) , .A1( u2_u7_u3_n146 ) , .ZN( u2_u7_u3_n147 ) );
  AND2_X1 u2_u7_u3_U80 (.A1( u2_u7_X_19 ) , .ZN( u2_u7_u3_n102 ) , .A2( u2_u7_u3_n172 ) );
  AND2_X1 u2_u7_u3_U81 (.A1( u2_u7_X_21 ) , .A2( u2_u7_X_24 ) , .ZN( u2_u7_u3_n100 ) );
  AND2_X1 u2_u7_u3_U82 (.A2( u2_u7_X_19 ) , .A1( u2_u7_X_20 ) , .ZN( u2_u7_u3_n104 ) );
  INV_X1 u2_u7_u3_U83 (.A( u2_u7_X_22 ) , .ZN( u2_u7_u3_n166 ) );
  INV_X1 u2_u7_u3_U84 (.A( u2_u7_X_21 ) , .ZN( u2_u7_u3_n171 ) );
  INV_X1 u2_u7_u3_U85 (.A( u2_u7_X_20 ) , .ZN( u2_u7_u3_n172 ) );
  OR4_X1 u2_u7_u3_U86 (.ZN( u2_out7_10 ) , .A4( u2_u7_u3_n136 ) , .A3( u2_u7_u3_n137 ) , .A1( u2_u7_u3_n138 ) , .A2( u2_u7_u3_n139 ) );
  OAI222_X1 u2_u7_u3_U87 (.C1( u2_u7_u3_n128 ) , .ZN( u2_u7_u3_n137 ) , .B1( u2_u7_u3_n148 ) , .A2( u2_u7_u3_n150 ) , .B2( u2_u7_u3_n154 ) , .C2( u2_u7_u3_n164 ) , .A1( u2_u7_u3_n167 ) );
  OAI221_X1 u2_u7_u3_U88 (.A( u2_u7_u3_n134 ) , .B2( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n136 ) , .C1( u2_u7_u3_n149 ) , .B1( u2_u7_u3_n151 ) , .C2( u2_u7_u3_n183 ) );
  NAND4_X1 u2_u7_u3_U89 (.ZN( u2_out7_26 ) , .A4( u2_u7_u3_n109 ) , .A3( u2_u7_u3_n110 ) , .A2( u2_u7_u3_n111 ) , .A1( u2_u7_u3_n173 ) );
  INV_X1 u2_u7_u3_U9 (.A( u2_u7_u3_n143 ) , .ZN( u2_u7_u3_n168 ) );
  INV_X1 u2_u7_u3_U90 (.ZN( u2_u7_u3_n173 ) , .A( u2_u7_u3_n94 ) );
  OAI21_X1 u2_u7_u3_U91 (.ZN( u2_u7_u3_n111 ) , .B2( u2_u7_u3_n117 ) , .A( u2_u7_u3_n133 ) , .B1( u2_u7_u3_n176 ) );
  NAND4_X1 u2_u7_u3_U92 (.ZN( u2_out7_20 ) , .A4( u2_u7_u3_n122 ) , .A3( u2_u7_u3_n123 ) , .A1( u2_u7_u3_n175 ) , .A2( u2_u7_u3_n180 ) );
  INV_X1 u2_u7_u3_U93 (.A( u2_u7_u3_n126 ) , .ZN( u2_u7_u3_n180 ) );
  INV_X1 u2_u7_u3_U94 (.A( u2_u7_u3_n112 ) , .ZN( u2_u7_u3_n175 ) );
  NAND4_X1 u2_u7_u3_U95 (.ZN( u2_out7_1 ) , .A4( u2_u7_u3_n161 ) , .A3( u2_u7_u3_n162 ) , .A2( u2_u7_u3_n163 ) , .A1( u2_u7_u3_n185 ) );
  NAND2_X1 u2_u7_u3_U96 (.ZN( u2_u7_u3_n163 ) , .A2( u2_u7_u3_n170 ) , .A1( u2_u7_u3_n176 ) );
  AOI22_X1 u2_u7_u3_U97 (.B2( u2_u7_u3_n140 ) , .B1( u2_u7_u3_n141 ) , .A2( u2_u7_u3_n142 ) , .ZN( u2_u7_u3_n162 ) , .A1( u2_u7_u3_n177 ) );
  NAND3_X1 u2_u7_u3_U98 (.A1( u2_u7_u3_n114 ) , .ZN( u2_u7_u3_n115 ) , .A2( u2_u7_u3_n145 ) , .A3( u2_u7_u3_n153 ) );
  NAND3_X1 u2_u7_u3_U99 (.ZN( u2_u7_u3_n129 ) , .A2( u2_u7_u3_n144 ) , .A1( u2_u7_u3_n153 ) , .A3( u2_u7_u3_n182 ) );
  OAI21_X1 u2_u7_u7_U10 (.A( u2_u7_u7_n161 ) , .B1( u2_u7_u7_n168 ) , .B2( u2_u7_u7_n173 ) , .ZN( u2_u7_u7_n91 ) );
  AOI211_X1 u2_u7_u7_U11 (.A( u2_u7_u7_n117 ) , .ZN( u2_u7_u7_n118 ) , .C2( u2_u7_u7_n126 ) , .C1( u2_u7_u7_n177 ) , .B( u2_u7_u7_n180 ) );
  OAI22_X1 u2_u7_u7_U12 (.B1( u2_u7_u7_n115 ) , .ZN( u2_u7_u7_n117 ) , .A2( u2_u7_u7_n133 ) , .A1( u2_u7_u7_n137 ) , .B2( u2_u7_u7_n162 ) );
  INV_X1 u2_u7_u7_U13 (.A( u2_u7_u7_n116 ) , .ZN( u2_u7_u7_n180 ) );
  NOR3_X1 u2_u7_u7_U14 (.ZN( u2_u7_u7_n115 ) , .A3( u2_u7_u7_n145 ) , .A2( u2_u7_u7_n168 ) , .A1( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U15 (.A( u2_u7_u7_n133 ) , .ZN( u2_u7_u7_n176 ) );
  NOR3_X1 u2_u7_u7_U16 (.A2( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n135 ) , .ZN( u2_u7_u7_n136 ) , .A3( u2_u7_u7_n171 ) );
  NOR2_X1 u2_u7_u7_U17 (.A1( u2_u7_u7_n130 ) , .A2( u2_u7_u7_n134 ) , .ZN( u2_u7_u7_n153 ) );
  AOI21_X1 u2_u7_u7_U18 (.ZN( u2_u7_u7_n104 ) , .B2( u2_u7_u7_n112 ) , .B1( u2_u7_u7_n127 ) , .A( u2_u7_u7_n164 ) );
  AOI21_X1 u2_u7_u7_U19 (.ZN( u2_u7_u7_n106 ) , .B1( u2_u7_u7_n133 ) , .B2( u2_u7_u7_n146 ) , .A( u2_u7_u7_n162 ) );
  AOI21_X1 u2_u7_u7_U20 (.A( u2_u7_u7_n101 ) , .ZN( u2_u7_u7_n107 ) , .B2( u2_u7_u7_n128 ) , .B1( u2_u7_u7_n175 ) );
  INV_X1 u2_u7_u7_U21 (.A( u2_u7_u7_n101 ) , .ZN( u2_u7_u7_n165 ) );
  NOR2_X1 u2_u7_u7_U22 (.ZN( u2_u7_u7_n111 ) , .A2( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U23 (.A( u2_u7_u7_n138 ) , .ZN( u2_u7_u7_n171 ) );
  INV_X1 u2_u7_u7_U24 (.A( u2_u7_u7_n131 ) , .ZN( u2_u7_u7_n177 ) );
  INV_X1 u2_u7_u7_U25 (.A( u2_u7_u7_n110 ) , .ZN( u2_u7_u7_n174 ) );
  NAND2_X1 u2_u7_u7_U26 (.A1( u2_u7_u7_n129 ) , .A2( u2_u7_u7_n132 ) , .ZN( u2_u7_u7_n149 ) );
  NAND2_X1 u2_u7_u7_U27 (.A1( u2_u7_u7_n113 ) , .A2( u2_u7_u7_n124 ) , .ZN( u2_u7_u7_n130 ) );
  INV_X1 u2_u7_u7_U28 (.A( u2_u7_u7_n112 ) , .ZN( u2_u7_u7_n173 ) );
  INV_X1 u2_u7_u7_U29 (.A( u2_u7_u7_n128 ) , .ZN( u2_u7_u7_n168 ) );
  OAI21_X1 u2_u7_u7_U3 (.ZN( u2_u7_u7_n159 ) , .A( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n171 ) , .B1( u2_u7_u7_n174 ) );
  INV_X1 u2_u7_u7_U30 (.A( u2_u7_u7_n148 ) , .ZN( u2_u7_u7_n169 ) );
  INV_X1 u2_u7_u7_U31 (.A( u2_u7_u7_n127 ) , .ZN( u2_u7_u7_n179 ) );
  NOR2_X1 u2_u7_u7_U32 (.ZN( u2_u7_u7_n101 ) , .A2( u2_u7_u7_n150 ) , .A1( u2_u7_u7_n156 ) );
  AOI211_X1 u2_u7_u7_U33 (.B( u2_u7_u7_n139 ) , .A( u2_u7_u7_n140 ) , .C2( u2_u7_u7_n141 ) , .ZN( u2_u7_u7_n142 ) , .C1( u2_u7_u7_n156 ) );
  NAND4_X1 u2_u7_u7_U34 (.A3( u2_u7_u7_n127 ) , .A2( u2_u7_u7_n128 ) , .A1( u2_u7_u7_n129 ) , .ZN( u2_u7_u7_n141 ) , .A4( u2_u7_u7_n147 ) );
  AOI21_X1 u2_u7_u7_U35 (.A( u2_u7_u7_n137 ) , .B1( u2_u7_u7_n138 ) , .ZN( u2_u7_u7_n139 ) , .B2( u2_u7_u7_n146 ) );
  OAI22_X1 u2_u7_u7_U36 (.B1( u2_u7_u7_n136 ) , .ZN( u2_u7_u7_n140 ) , .A1( u2_u7_u7_n153 ) , .B2( u2_u7_u7_n162 ) , .A2( u2_u7_u7_n164 ) );
  INV_X1 u2_u7_u7_U37 (.A( u2_u7_u7_n125 ) , .ZN( u2_u7_u7_n161 ) );
  AOI21_X1 u2_u7_u7_U38 (.ZN( u2_u7_u7_n123 ) , .B1( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n177 ) , .A( u2_u7_u7_n97 ) );
  AOI21_X1 u2_u7_u7_U39 (.B2( u2_u7_u7_n113 ) , .B1( u2_u7_u7_n124 ) , .A( u2_u7_u7_n125 ) , .ZN( u2_u7_u7_n97 ) );
  INV_X1 u2_u7_u7_U4 (.A( u2_u7_u7_n149 ) , .ZN( u2_u7_u7_n175 ) );
  INV_X1 u2_u7_u7_U40 (.A( u2_u7_u7_n152 ) , .ZN( u2_u7_u7_n162 ) );
  AOI22_X1 u2_u7_u7_U41 (.A2( u2_u7_u7_n114 ) , .ZN( u2_u7_u7_n119 ) , .B1( u2_u7_u7_n130 ) , .A1( u2_u7_u7_n156 ) , .B2( u2_u7_u7_n165 ) );
  NAND2_X1 u2_u7_u7_U42 (.A2( u2_u7_u7_n112 ) , .ZN( u2_u7_u7_n114 ) , .A1( u2_u7_u7_n175 ) );
  NOR2_X1 u2_u7_u7_U43 (.ZN( u2_u7_u7_n137 ) , .A1( u2_u7_u7_n150 ) , .A2( u2_u7_u7_n161 ) );
  AND2_X1 u2_u7_u7_U44 (.ZN( u2_u7_u7_n145 ) , .A2( u2_u7_u7_n98 ) , .A1( u2_u7_u7_n99 ) );
  AOI21_X1 u2_u7_u7_U45 (.ZN( u2_u7_u7_n105 ) , .B2( u2_u7_u7_n110 ) , .A( u2_u7_u7_n125 ) , .B1( u2_u7_u7_n147 ) );
  NAND2_X1 u2_u7_u7_U46 (.ZN( u2_u7_u7_n146 ) , .A1( u2_u7_u7_n95 ) , .A2( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U47 (.A2( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n147 ) , .A1( u2_u7_u7_n93 ) );
  NAND2_X1 u2_u7_u7_U48 (.A1( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n127 ) , .A2( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U49 (.A2( u2_u7_u7_n102 ) , .A1( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n133 ) );
  INV_X1 u2_u7_u7_U5 (.A( u2_u7_u7_n154 ) , .ZN( u2_u7_u7_n178 ) );
  OR2_X1 u2_u7_u7_U50 (.ZN( u2_u7_u7_n126 ) , .A2( u2_u7_u7_n152 ) , .A1( u2_u7_u7_n156 ) );
  NAND2_X1 u2_u7_u7_U51 (.ZN( u2_u7_u7_n112 ) , .A2( u2_u7_u7_n96 ) , .A1( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U52 (.A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n128 ) , .A1( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U53 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n113 ) , .A2( u2_u7_u7_n93 ) );
  NAND2_X1 u2_u7_u7_U54 (.ZN( u2_u7_u7_n110 ) , .A1( u2_u7_u7_n95 ) , .A2( u2_u7_u7_n96 ) );
  INV_X1 u2_u7_u7_U55 (.A( u2_u7_u7_n150 ) , .ZN( u2_u7_u7_n164 ) );
  AND2_X1 u2_u7_u7_U56 (.ZN( u2_u7_u7_n134 ) , .A1( u2_u7_u7_n93 ) , .A2( u2_u7_u7_n98 ) );
  NAND2_X1 u2_u7_u7_U57 (.A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n124 ) , .A1( u2_u7_u7_n96 ) );
  NAND2_X1 u2_u7_u7_U58 (.A1( u2_u7_u7_n100 ) , .A2( u2_u7_u7_n102 ) , .ZN( u2_u7_u7_n129 ) );
  NAND2_X1 u2_u7_u7_U59 (.A2( u2_u7_u7_n103 ) , .ZN( u2_u7_u7_n131 ) , .A1( u2_u7_u7_n95 ) );
  AOI211_X1 u2_u7_u7_U6 (.ZN( u2_u7_u7_n116 ) , .A( u2_u7_u7_n155 ) , .C1( u2_u7_u7_n161 ) , .C2( u2_u7_u7_n171 ) , .B( u2_u7_u7_n94 ) );
  NAND2_X1 u2_u7_u7_U60 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n138 ) , .A2( u2_u7_u7_n99 ) );
  NAND2_X1 u2_u7_u7_U61 (.ZN( u2_u7_u7_n132 ) , .A1( u2_u7_u7_n93 ) , .A2( u2_u7_u7_n96 ) );
  NAND2_X1 u2_u7_u7_U62 (.A1( u2_u7_u7_n100 ) , .ZN( u2_u7_u7_n148 ) , .A2( u2_u7_u7_n95 ) );
  AOI211_X1 u2_u7_u7_U63 (.B( u2_u7_u7_n154 ) , .A( u2_u7_u7_n155 ) , .C1( u2_u7_u7_n156 ) , .ZN( u2_u7_u7_n157 ) , .C2( u2_u7_u7_n172 ) );
  INV_X1 u2_u7_u7_U64 (.A( u2_u7_u7_n153 ) , .ZN( u2_u7_u7_n172 ) );
  NOR2_X1 u2_u7_u7_U65 (.A2( u2_u7_X_47 ) , .ZN( u2_u7_u7_n150 ) , .A1( u2_u7_u7_n163 ) );
  NOR2_X1 u2_u7_u7_U66 (.A2( u2_u7_X_43 ) , .A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n103 ) );
  NOR2_X1 u2_u7_u7_U67 (.A2( u2_u7_X_48 ) , .A1( u2_u7_u7_n166 ) , .ZN( u2_u7_u7_n95 ) );
  NOR2_X1 u2_u7_u7_U68 (.A2( u2_u7_X_45 ) , .A1( u2_u7_X_48 ) , .ZN( u2_u7_u7_n99 ) );
  NOR2_X1 u2_u7_u7_U69 (.A2( u2_u7_X_44 ) , .A1( u2_u7_u7_n167 ) , .ZN( u2_u7_u7_n98 ) );
  OAI222_X1 u2_u7_u7_U7 (.C2( u2_u7_u7_n101 ) , .B2( u2_u7_u7_n111 ) , .A1( u2_u7_u7_n113 ) , .C1( u2_u7_u7_n146 ) , .A2( u2_u7_u7_n162 ) , .B1( u2_u7_u7_n164 ) , .ZN( u2_u7_u7_n94 ) );
  NOR2_X1 u2_u7_u7_U70 (.A2( u2_u7_X_46 ) , .A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n152 ) );
  NAND2_X1 u2_u7_u7_U71 (.A2( u2_u7_X_46 ) , .A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n125 ) );
  AND2_X1 u2_u7_u7_U72 (.A1( u2_u7_X_47 ) , .ZN( u2_u7_u7_n156 ) , .A2( u2_u7_u7_n163 ) );
  AND2_X1 u2_u7_u7_U73 (.A2( u2_u7_X_45 ) , .A1( u2_u7_X_48 ) , .ZN( u2_u7_u7_n102 ) );
  AND2_X1 u2_u7_u7_U74 (.A2( u2_u7_X_43 ) , .A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n96 ) );
  AND2_X1 u2_u7_u7_U75 (.A1( u2_u7_X_44 ) , .ZN( u2_u7_u7_n100 ) , .A2( u2_u7_u7_n167 ) );
  AND2_X1 u2_u7_u7_U76 (.A1( u2_u7_X_48 ) , .A2( u2_u7_u7_n166 ) , .ZN( u2_u7_u7_n93 ) );
  INV_X1 u2_u7_u7_U77 (.A( u2_u7_X_46 ) , .ZN( u2_u7_u7_n163 ) );
  INV_X1 u2_u7_u7_U78 (.A( u2_u7_X_43 ) , .ZN( u2_u7_u7_n167 ) );
  INV_X1 u2_u7_u7_U79 (.A( u2_u7_X_45 ) , .ZN( u2_u7_u7_n166 ) );
  OAI221_X1 u2_u7_u7_U8 (.C1( u2_u7_u7_n101 ) , .C2( u2_u7_u7_n147 ) , .ZN( u2_u7_u7_n155 ) , .B2( u2_u7_u7_n162 ) , .A( u2_u7_u7_n91 ) , .B1( u2_u7_u7_n92 ) );
  NAND4_X1 u2_u7_u7_U80 (.ZN( u2_out7_5 ) , .A4( u2_u7_u7_n108 ) , .A3( u2_u7_u7_n109 ) , .A1( u2_u7_u7_n116 ) , .A2( u2_u7_u7_n123 ) );
  AOI22_X1 u2_u7_u7_U81 (.ZN( u2_u7_u7_n109 ) , .A2( u2_u7_u7_n126 ) , .B2( u2_u7_u7_n145 ) , .B1( u2_u7_u7_n156 ) , .A1( u2_u7_u7_n171 ) );
  NOR4_X1 u2_u7_u7_U82 (.A4( u2_u7_u7_n104 ) , .A3( u2_u7_u7_n105 ) , .A2( u2_u7_u7_n106 ) , .A1( u2_u7_u7_n107 ) , .ZN( u2_u7_u7_n108 ) );
  NAND4_X1 u2_u7_u7_U83 (.ZN( u2_out7_27 ) , .A4( u2_u7_u7_n118 ) , .A3( u2_u7_u7_n119 ) , .A2( u2_u7_u7_n120 ) , .A1( u2_u7_u7_n121 ) );
  OAI21_X1 u2_u7_u7_U84 (.ZN( u2_u7_u7_n121 ) , .B2( u2_u7_u7_n145 ) , .A( u2_u7_u7_n150 ) , .B1( u2_u7_u7_n174 ) );
  OAI21_X1 u2_u7_u7_U85 (.ZN( u2_u7_u7_n120 ) , .A( u2_u7_u7_n161 ) , .B2( u2_u7_u7_n170 ) , .B1( u2_u7_u7_n179 ) );
  NAND4_X1 u2_u7_u7_U86 (.ZN( u2_out7_21 ) , .A4( u2_u7_u7_n157 ) , .A3( u2_u7_u7_n158 ) , .A2( u2_u7_u7_n159 ) , .A1( u2_u7_u7_n160 ) );
  OAI21_X1 u2_u7_u7_U87 (.B1( u2_u7_u7_n145 ) , .ZN( u2_u7_u7_n160 ) , .A( u2_u7_u7_n161 ) , .B2( u2_u7_u7_n177 ) );
  AOI22_X1 u2_u7_u7_U88 (.B2( u2_u7_u7_n149 ) , .B1( u2_u7_u7_n150 ) , .A2( u2_u7_u7_n151 ) , .A1( u2_u7_u7_n152 ) , .ZN( u2_u7_u7_n158 ) );
  NAND4_X1 u2_u7_u7_U89 (.ZN( u2_out7_15 ) , .A4( u2_u7_u7_n142 ) , .A3( u2_u7_u7_n143 ) , .A2( u2_u7_u7_n144 ) , .A1( u2_u7_u7_n178 ) );
  AND3_X1 u2_u7_u7_U9 (.A3( u2_u7_u7_n110 ) , .A2( u2_u7_u7_n127 ) , .A1( u2_u7_u7_n132 ) , .ZN( u2_u7_u7_n92 ) );
  OR2_X1 u2_u7_u7_U90 (.A2( u2_u7_u7_n125 ) , .A1( u2_u7_u7_n129 ) , .ZN( u2_u7_u7_n144 ) );
  AOI22_X1 u2_u7_u7_U91 (.A2( u2_u7_u7_n126 ) , .ZN( u2_u7_u7_n143 ) , .B2( u2_u7_u7_n165 ) , .B1( u2_u7_u7_n173 ) , .A1( u2_u7_u7_n174 ) );
  OAI211_X1 u2_u7_u7_U92 (.B( u2_u7_u7_n122 ) , .A( u2_u7_u7_n123 ) , .C2( u2_u7_u7_n124 ) , .ZN( u2_u7_u7_n154 ) , .C1( u2_u7_u7_n162 ) );
  AOI222_X1 u2_u7_u7_U93 (.ZN( u2_u7_u7_n122 ) , .C2( u2_u7_u7_n126 ) , .C1( u2_u7_u7_n145 ) , .B1( u2_u7_u7_n161 ) , .A2( u2_u7_u7_n165 ) , .B2( u2_u7_u7_n170 ) , .A1( u2_u7_u7_n176 ) );
  INV_X1 u2_u7_u7_U94 (.A( u2_u7_u7_n111 ) , .ZN( u2_u7_u7_n170 ) );
  NAND3_X1 u2_u7_u7_U95 (.A3( u2_u7_u7_n146 ) , .A2( u2_u7_u7_n147 ) , .A1( u2_u7_u7_n148 ) , .ZN( u2_u7_u7_n151 ) );
  NAND3_X1 u2_u7_u7_U96 (.A3( u2_u7_u7_n131 ) , .A2( u2_u7_u7_n132 ) , .A1( u2_u7_u7_n133 ) , .ZN( u2_u7_u7_n135 ) );
  XOR2_X1 u2_u8_U11 (.B( u2_K9_44 ) , .A( u2_R7_29 ) , .Z( u2_u8_X_44 ) );
  XOR2_X1 u2_u8_U12 (.B( u2_K9_43 ) , .A( u2_R7_28 ) , .Z( u2_u8_X_43 ) );
  XOR2_X1 u2_u8_U13 (.B( u2_K9_42 ) , .A( u2_R7_29 ) , .Z( u2_u8_X_42 ) );
  XOR2_X1 u2_u8_U14 (.B( u2_K9_41 ) , .A( u2_R7_28 ) , .Z( u2_u8_X_41 ) );
  XOR2_X1 u2_u8_U18 (.B( u2_K9_38 ) , .A( u2_R7_25 ) , .Z( u2_u8_X_38 ) );
  XOR2_X1 u2_u8_U19 (.B( u2_K9_37 ) , .A( u2_R7_24 ) , .Z( u2_u8_X_37 ) );
  XOR2_X1 u2_u8_U20 (.B( u2_K9_36 ) , .A( u2_R7_25 ) , .Z( u2_u8_X_36 ) );
  XOR2_X1 u2_u8_U21 (.B( u2_K9_35 ) , .A( u2_R7_24 ) , .Z( u2_u8_X_35 ) );
  XOR2_X1 u2_u8_U23 (.B( u2_K9_33 ) , .A( u2_R7_22 ) , .Z( u2_u8_X_33 ) );
  XOR2_X1 u2_u8_U7 (.B( u2_K9_48 ) , .A( u2_R7_1 ) , .Z( u2_u8_X_48 ) );
  NOR2_X1 u2_u8_u5_U10 (.ZN( u2_u8_u5_n135 ) , .A1( u2_u8_u5_n173 ) , .A2( u2_u8_u5_n176 ) );
  NOR3_X1 u2_u8_u5_U100 (.A3( u2_u8_u5_n141 ) , .A1( u2_u8_u5_n142 ) , .ZN( u2_u8_u5_n143 ) , .A2( u2_u8_u5_n191 ) );
  NAND4_X1 u2_u8_u5_U101 (.ZN( u2_out8_4 ) , .A4( u2_u8_u5_n112 ) , .A2( u2_u8_u5_n113 ) , .A1( u2_u8_u5_n114 ) , .A3( u2_u8_u5_n195 ) );
  AOI211_X1 u2_u8_u5_U102 (.A( u2_u8_u5_n110 ) , .C1( u2_u8_u5_n111 ) , .ZN( u2_u8_u5_n112 ) , .B( u2_u8_u5_n118 ) , .C2( u2_u8_u5_n177 ) );
  INV_X1 u2_u8_u5_U103 (.A( u2_u8_u5_n102 ) , .ZN( u2_u8_u5_n195 ) );
  NAND3_X1 u2_u8_u5_U104 (.A2( u2_u8_u5_n154 ) , .A3( u2_u8_u5_n158 ) , .A1( u2_u8_u5_n161 ) , .ZN( u2_u8_u5_n99 ) );
  INV_X1 u2_u8_u5_U11 (.A( u2_u8_u5_n121 ) , .ZN( u2_u8_u5_n177 ) );
  NOR2_X1 u2_u8_u5_U12 (.ZN( u2_u8_u5_n160 ) , .A2( u2_u8_u5_n173 ) , .A1( u2_u8_u5_n177 ) );
  INV_X1 u2_u8_u5_U13 (.A( u2_u8_u5_n150 ) , .ZN( u2_u8_u5_n174 ) );
  AOI21_X1 u2_u8_u5_U14 (.A( u2_u8_u5_n160 ) , .B2( u2_u8_u5_n161 ) , .ZN( u2_u8_u5_n162 ) , .B1( u2_u8_u5_n192 ) );
  INV_X1 u2_u8_u5_U15 (.A( u2_u8_u5_n159 ) , .ZN( u2_u8_u5_n192 ) );
  AOI21_X1 u2_u8_u5_U16 (.A( u2_u8_u5_n156 ) , .B2( u2_u8_u5_n157 ) , .B1( u2_u8_u5_n158 ) , .ZN( u2_u8_u5_n163 ) );
  AOI21_X1 u2_u8_u5_U17 (.B2( u2_u8_u5_n139 ) , .B1( u2_u8_u5_n140 ) , .ZN( u2_u8_u5_n141 ) , .A( u2_u8_u5_n150 ) );
  OAI21_X1 u2_u8_u5_U18 (.A( u2_u8_u5_n133 ) , .B2( u2_u8_u5_n134 ) , .B1( u2_u8_u5_n135 ) , .ZN( u2_u8_u5_n142 ) );
  OAI21_X1 u2_u8_u5_U19 (.ZN( u2_u8_u5_n133 ) , .B2( u2_u8_u5_n147 ) , .A( u2_u8_u5_n173 ) , .B1( u2_u8_u5_n188 ) );
  NAND2_X1 u2_u8_u5_U20 (.A2( u2_u8_u5_n119 ) , .A1( u2_u8_u5_n123 ) , .ZN( u2_u8_u5_n137 ) );
  INV_X1 u2_u8_u5_U21 (.A( u2_u8_u5_n155 ) , .ZN( u2_u8_u5_n194 ) );
  NAND2_X1 u2_u8_u5_U22 (.A1( u2_u8_u5_n121 ) , .ZN( u2_u8_u5_n132 ) , .A2( u2_u8_u5_n172 ) );
  NAND2_X1 u2_u8_u5_U23 (.A2( u2_u8_u5_n122 ) , .ZN( u2_u8_u5_n136 ) , .A1( u2_u8_u5_n154 ) );
  NAND2_X1 u2_u8_u5_U24 (.A2( u2_u8_u5_n119 ) , .A1( u2_u8_u5_n120 ) , .ZN( u2_u8_u5_n159 ) );
  INV_X1 u2_u8_u5_U25 (.A( u2_u8_u5_n156 ) , .ZN( u2_u8_u5_n175 ) );
  INV_X1 u2_u8_u5_U26 (.A( u2_u8_u5_n158 ) , .ZN( u2_u8_u5_n188 ) );
  INV_X1 u2_u8_u5_U27 (.A( u2_u8_u5_n152 ) , .ZN( u2_u8_u5_n179 ) );
  INV_X1 u2_u8_u5_U28 (.A( u2_u8_u5_n140 ) , .ZN( u2_u8_u5_n182 ) );
  INV_X1 u2_u8_u5_U29 (.A( u2_u8_u5_n151 ) , .ZN( u2_u8_u5_n183 ) );
  NOR2_X1 u2_u8_u5_U3 (.ZN( u2_u8_u5_n134 ) , .A1( u2_u8_u5_n183 ) , .A2( u2_u8_u5_n190 ) );
  INV_X1 u2_u8_u5_U30 (.A( u2_u8_u5_n123 ) , .ZN( u2_u8_u5_n185 ) );
  INV_X1 u2_u8_u5_U31 (.A( u2_u8_u5_n161 ) , .ZN( u2_u8_u5_n184 ) );
  INV_X1 u2_u8_u5_U32 (.A( u2_u8_u5_n139 ) , .ZN( u2_u8_u5_n189 ) );
  INV_X1 u2_u8_u5_U33 (.A( u2_u8_u5_n157 ) , .ZN( u2_u8_u5_n190 ) );
  INV_X1 u2_u8_u5_U34 (.A( u2_u8_u5_n120 ) , .ZN( u2_u8_u5_n193 ) );
  NAND2_X1 u2_u8_u5_U35 (.ZN( u2_u8_u5_n111 ) , .A1( u2_u8_u5_n140 ) , .A2( u2_u8_u5_n155 ) );
  NOR2_X1 u2_u8_u5_U36 (.ZN( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n170 ) , .A2( u2_u8_u5_n180 ) );
  INV_X1 u2_u8_u5_U37 (.A( u2_u8_u5_n117 ) , .ZN( u2_u8_u5_n196 ) );
  OAI221_X1 u2_u8_u5_U38 (.A( u2_u8_u5_n116 ) , .ZN( u2_u8_u5_n117 ) , .B2( u2_u8_u5_n119 ) , .C1( u2_u8_u5_n153 ) , .C2( u2_u8_u5_n158 ) , .B1( u2_u8_u5_n172 ) );
  AOI222_X1 u2_u8_u5_U39 (.ZN( u2_u8_u5_n116 ) , .B2( u2_u8_u5_n145 ) , .C1( u2_u8_u5_n148 ) , .A2( u2_u8_u5_n174 ) , .C2( u2_u8_u5_n177 ) , .B1( u2_u8_u5_n187 ) , .A1( u2_u8_u5_n193 ) );
  INV_X1 u2_u8_u5_U4 (.A( u2_u8_u5_n138 ) , .ZN( u2_u8_u5_n191 ) );
  INV_X1 u2_u8_u5_U40 (.A( u2_u8_u5_n115 ) , .ZN( u2_u8_u5_n187 ) );
  OAI221_X1 u2_u8_u5_U41 (.A( u2_u8_u5_n101 ) , .ZN( u2_u8_u5_n102 ) , .C2( u2_u8_u5_n115 ) , .C1( u2_u8_u5_n126 ) , .B1( u2_u8_u5_n134 ) , .B2( u2_u8_u5_n160 ) );
  OAI21_X1 u2_u8_u5_U42 (.ZN( u2_u8_u5_n101 ) , .B1( u2_u8_u5_n137 ) , .A( u2_u8_u5_n146 ) , .B2( u2_u8_u5_n147 ) );
  AOI22_X1 u2_u8_u5_U43 (.B2( u2_u8_u5_n131 ) , .A2( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n169 ) , .B1( u2_u8_u5_n174 ) , .A1( u2_u8_u5_n185 ) );
  NOR2_X1 u2_u8_u5_U44 (.A1( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n150 ) , .A2( u2_u8_u5_n173 ) );
  AOI21_X1 u2_u8_u5_U45 (.A( u2_u8_u5_n118 ) , .B2( u2_u8_u5_n145 ) , .ZN( u2_u8_u5_n168 ) , .B1( u2_u8_u5_n186 ) );
  INV_X1 u2_u8_u5_U46 (.A( u2_u8_u5_n122 ) , .ZN( u2_u8_u5_n186 ) );
  NOR2_X1 u2_u8_u5_U47 (.A1( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n152 ) , .A2( u2_u8_u5_n176 ) );
  NOR2_X1 u2_u8_u5_U48 (.A1( u2_u8_u5_n115 ) , .ZN( u2_u8_u5_n118 ) , .A2( u2_u8_u5_n153 ) );
  NOR2_X1 u2_u8_u5_U49 (.A2( u2_u8_u5_n145 ) , .ZN( u2_u8_u5_n156 ) , .A1( u2_u8_u5_n174 ) );
  OAI21_X1 u2_u8_u5_U5 (.B2( u2_u8_u5_n136 ) , .B1( u2_u8_u5_n137 ) , .ZN( u2_u8_u5_n138 ) , .A( u2_u8_u5_n177 ) );
  NOR2_X1 u2_u8_u5_U50 (.ZN( u2_u8_u5_n121 ) , .A2( u2_u8_u5_n145 ) , .A1( u2_u8_u5_n176 ) );
  AOI22_X1 u2_u8_u5_U51 (.ZN( u2_u8_u5_n114 ) , .A2( u2_u8_u5_n137 ) , .A1( u2_u8_u5_n145 ) , .B2( u2_u8_u5_n175 ) , .B1( u2_u8_u5_n193 ) );
  OAI211_X1 u2_u8_u5_U52 (.B( u2_u8_u5_n124 ) , .A( u2_u8_u5_n125 ) , .C2( u2_u8_u5_n126 ) , .C1( u2_u8_u5_n127 ) , .ZN( u2_u8_u5_n128 ) );
  NOR3_X1 u2_u8_u5_U53 (.ZN( u2_u8_u5_n127 ) , .A1( u2_u8_u5_n136 ) , .A3( u2_u8_u5_n148 ) , .A2( u2_u8_u5_n182 ) );
  OAI21_X1 u2_u8_u5_U54 (.ZN( u2_u8_u5_n124 ) , .A( u2_u8_u5_n177 ) , .B2( u2_u8_u5_n183 ) , .B1( u2_u8_u5_n189 ) );
  OAI21_X1 u2_u8_u5_U55 (.ZN( u2_u8_u5_n125 ) , .A( u2_u8_u5_n174 ) , .B2( u2_u8_u5_n185 ) , .B1( u2_u8_u5_n190 ) );
  AOI21_X1 u2_u8_u5_U56 (.A( u2_u8_u5_n153 ) , .B2( u2_u8_u5_n154 ) , .B1( u2_u8_u5_n155 ) , .ZN( u2_u8_u5_n164 ) );
  AOI21_X1 u2_u8_u5_U57 (.ZN( u2_u8_u5_n110 ) , .B1( u2_u8_u5_n122 ) , .B2( u2_u8_u5_n139 ) , .A( u2_u8_u5_n153 ) );
  INV_X1 u2_u8_u5_U58 (.A( u2_u8_u5_n153 ) , .ZN( u2_u8_u5_n176 ) );
  INV_X1 u2_u8_u5_U59 (.A( u2_u8_u5_n126 ) , .ZN( u2_u8_u5_n173 ) );
  AOI222_X1 u2_u8_u5_U6 (.ZN( u2_u8_u5_n113 ) , .A1( u2_u8_u5_n131 ) , .C1( u2_u8_u5_n148 ) , .B2( u2_u8_u5_n174 ) , .C2( u2_u8_u5_n178 ) , .A2( u2_u8_u5_n179 ) , .B1( u2_u8_u5_n99 ) );
  AND2_X1 u2_u8_u5_U60 (.A2( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n107 ) , .ZN( u2_u8_u5_n147 ) );
  AND2_X1 u2_u8_u5_U61 (.A2( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n108 ) , .ZN( u2_u8_u5_n148 ) );
  NAND2_X1 u2_u8_u5_U62 (.A1( u2_u8_u5_n105 ) , .A2( u2_u8_u5_n106 ) , .ZN( u2_u8_u5_n158 ) );
  NAND2_X1 u2_u8_u5_U63 (.A2( u2_u8_u5_n108 ) , .A1( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n139 ) );
  NAND2_X1 u2_u8_u5_U64 (.A1( u2_u8_u5_n106 ) , .A2( u2_u8_u5_n108 ) , .ZN( u2_u8_u5_n119 ) );
  NAND2_X1 u2_u8_u5_U65 (.A2( u2_u8_u5_n103 ) , .A1( u2_u8_u5_n105 ) , .ZN( u2_u8_u5_n140 ) );
  NAND2_X1 u2_u8_u5_U66 (.A2( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n105 ) , .ZN( u2_u8_u5_n155 ) );
  NAND2_X1 u2_u8_u5_U67 (.A2( u2_u8_u5_n106 ) , .A1( u2_u8_u5_n107 ) , .ZN( u2_u8_u5_n122 ) );
  NAND2_X1 u2_u8_u5_U68 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n106 ) , .ZN( u2_u8_u5_n115 ) );
  NAND2_X1 u2_u8_u5_U69 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n103 ) , .ZN( u2_u8_u5_n161 ) );
  INV_X1 u2_u8_u5_U7 (.A( u2_u8_u5_n135 ) , .ZN( u2_u8_u5_n178 ) );
  NAND2_X1 u2_u8_u5_U70 (.A1( u2_u8_u5_n105 ) , .A2( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n154 ) );
  INV_X1 u2_u8_u5_U71 (.A( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n172 ) );
  NAND2_X1 u2_u8_u5_U72 (.A1( u2_u8_u5_n103 ) , .A2( u2_u8_u5_n108 ) , .ZN( u2_u8_u5_n123 ) );
  NAND2_X1 u2_u8_u5_U73 (.A2( u2_u8_u5_n103 ) , .A1( u2_u8_u5_n107 ) , .ZN( u2_u8_u5_n151 ) );
  NAND2_X1 u2_u8_u5_U74 (.A2( u2_u8_u5_n107 ) , .A1( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n120 ) );
  NAND2_X1 u2_u8_u5_U75 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n157 ) );
  AND2_X1 u2_u8_u5_U76 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n104 ) , .ZN( u2_u8_u5_n131 ) );
  NOR2_X1 u2_u8_u5_U77 (.A2( u2_u8_X_34 ) , .A1( u2_u8_X_35 ) , .ZN( u2_u8_u5_n145 ) );
  NOR2_X1 u2_u8_u5_U78 (.A2( u2_u8_X_34 ) , .ZN( u2_u8_u5_n146 ) , .A1( u2_u8_u5_n171 ) );
  NOR2_X1 u2_u8_u5_U79 (.A2( u2_u8_X_31 ) , .A1( u2_u8_X_32 ) , .ZN( u2_u8_u5_n103 ) );
  OAI22_X1 u2_u8_u5_U8 (.B2( u2_u8_u5_n149 ) , .B1( u2_u8_u5_n150 ) , .A2( u2_u8_u5_n151 ) , .A1( u2_u8_u5_n152 ) , .ZN( u2_u8_u5_n165 ) );
  NOR2_X1 u2_u8_u5_U80 (.A2( u2_u8_X_36 ) , .ZN( u2_u8_u5_n105 ) , .A1( u2_u8_u5_n180 ) );
  NOR2_X1 u2_u8_u5_U81 (.A2( u2_u8_X_33 ) , .ZN( u2_u8_u5_n108 ) , .A1( u2_u8_u5_n170 ) );
  NOR2_X1 u2_u8_u5_U82 (.A2( u2_u8_X_33 ) , .A1( u2_u8_X_36 ) , .ZN( u2_u8_u5_n107 ) );
  NOR2_X1 u2_u8_u5_U83 (.A2( u2_u8_X_31 ) , .ZN( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n181 ) );
  NAND2_X1 u2_u8_u5_U84 (.A2( u2_u8_X_34 ) , .A1( u2_u8_X_35 ) , .ZN( u2_u8_u5_n153 ) );
  NAND2_X1 u2_u8_u5_U85 (.A1( u2_u8_X_34 ) , .ZN( u2_u8_u5_n126 ) , .A2( u2_u8_u5_n171 ) );
  AND2_X1 u2_u8_u5_U86 (.A1( u2_u8_X_31 ) , .A2( u2_u8_X_32 ) , .ZN( u2_u8_u5_n106 ) );
  AND2_X1 u2_u8_u5_U87 (.A1( u2_u8_X_31 ) , .ZN( u2_u8_u5_n109 ) , .A2( u2_u8_u5_n181 ) );
  INV_X1 u2_u8_u5_U88 (.A( u2_u8_X_33 ) , .ZN( u2_u8_u5_n180 ) );
  INV_X1 u2_u8_u5_U89 (.A( u2_u8_X_35 ) , .ZN( u2_u8_u5_n171 ) );
  NOR3_X1 u2_u8_u5_U9 (.A2( u2_u8_u5_n147 ) , .A1( u2_u8_u5_n148 ) , .ZN( u2_u8_u5_n149 ) , .A3( u2_u8_u5_n194 ) );
  INV_X1 u2_u8_u5_U90 (.A( u2_u8_X_36 ) , .ZN( u2_u8_u5_n170 ) );
  INV_X1 u2_u8_u5_U91 (.A( u2_u8_X_32 ) , .ZN( u2_u8_u5_n181 ) );
  NAND4_X1 u2_u8_u5_U92 (.ZN( u2_out8_29 ) , .A4( u2_u8_u5_n129 ) , .A3( u2_u8_u5_n130 ) , .A2( u2_u8_u5_n168 ) , .A1( u2_u8_u5_n196 ) );
  AOI221_X1 u2_u8_u5_U93 (.A( u2_u8_u5_n128 ) , .ZN( u2_u8_u5_n129 ) , .C2( u2_u8_u5_n132 ) , .B2( u2_u8_u5_n159 ) , .B1( u2_u8_u5_n176 ) , .C1( u2_u8_u5_n184 ) );
  AOI222_X1 u2_u8_u5_U94 (.ZN( u2_u8_u5_n130 ) , .A2( u2_u8_u5_n146 ) , .B1( u2_u8_u5_n147 ) , .C2( u2_u8_u5_n175 ) , .B2( u2_u8_u5_n179 ) , .A1( u2_u8_u5_n188 ) , .C1( u2_u8_u5_n194 ) );
  NAND4_X1 u2_u8_u5_U95 (.ZN( u2_out8_19 ) , .A4( u2_u8_u5_n166 ) , .A3( u2_u8_u5_n167 ) , .A2( u2_u8_u5_n168 ) , .A1( u2_u8_u5_n169 ) );
  AOI22_X1 u2_u8_u5_U96 (.B2( u2_u8_u5_n145 ) , .A2( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n167 ) , .B1( u2_u8_u5_n182 ) , .A1( u2_u8_u5_n189 ) );
  NOR4_X1 u2_u8_u5_U97 (.A4( u2_u8_u5_n162 ) , .A3( u2_u8_u5_n163 ) , .A2( u2_u8_u5_n164 ) , .A1( u2_u8_u5_n165 ) , .ZN( u2_u8_u5_n166 ) );
  NAND4_X1 u2_u8_u5_U98 (.ZN( u2_out8_11 ) , .A4( u2_u8_u5_n143 ) , .A3( u2_u8_u5_n144 ) , .A2( u2_u8_u5_n169 ) , .A1( u2_u8_u5_n196 ) );
  AOI22_X1 u2_u8_u5_U99 (.A2( u2_u8_u5_n132 ) , .ZN( u2_u8_u5_n144 ) , .B2( u2_u8_u5_n145 ) , .B1( u2_u8_u5_n184 ) , .A1( u2_u8_u5_n194 ) );
  AOI22_X1 u2_u8_u6_U10 (.A2( u2_u8_u6_n151 ) , .B2( u2_u8_u6_n161 ) , .A1( u2_u8_u6_n167 ) , .B1( u2_u8_u6_n170 ) , .ZN( u2_u8_u6_n89 ) );
  AOI21_X1 u2_u8_u6_U11 (.B1( u2_u8_u6_n107 ) , .B2( u2_u8_u6_n132 ) , .A( u2_u8_u6_n158 ) , .ZN( u2_u8_u6_n88 ) );
  AOI21_X1 u2_u8_u6_U12 (.B2( u2_u8_u6_n147 ) , .B1( u2_u8_u6_n148 ) , .ZN( u2_u8_u6_n149 ) , .A( u2_u8_u6_n158 ) );
  AOI21_X1 u2_u8_u6_U13 (.ZN( u2_u8_u6_n106 ) , .A( u2_u8_u6_n142 ) , .B2( u2_u8_u6_n159 ) , .B1( u2_u8_u6_n164 ) );
  INV_X1 u2_u8_u6_U14 (.A( u2_u8_u6_n155 ) , .ZN( u2_u8_u6_n161 ) );
  INV_X1 u2_u8_u6_U15 (.A( u2_u8_u6_n128 ) , .ZN( u2_u8_u6_n164 ) );
  NAND2_X1 u2_u8_u6_U16 (.ZN( u2_u8_u6_n110 ) , .A1( u2_u8_u6_n122 ) , .A2( u2_u8_u6_n129 ) );
  NAND2_X1 u2_u8_u6_U17 (.ZN( u2_u8_u6_n124 ) , .A2( u2_u8_u6_n146 ) , .A1( u2_u8_u6_n148 ) );
  INV_X1 u2_u8_u6_U18 (.A( u2_u8_u6_n132 ) , .ZN( u2_u8_u6_n171 ) );
  AND2_X1 u2_u8_u6_U19 (.A1( u2_u8_u6_n100 ) , .ZN( u2_u8_u6_n130 ) , .A2( u2_u8_u6_n147 ) );
  INV_X1 u2_u8_u6_U20 (.A( u2_u8_u6_n127 ) , .ZN( u2_u8_u6_n173 ) );
  INV_X1 u2_u8_u6_U21 (.A( u2_u8_u6_n121 ) , .ZN( u2_u8_u6_n167 ) );
  INV_X1 u2_u8_u6_U22 (.A( u2_u8_u6_n100 ) , .ZN( u2_u8_u6_n169 ) );
  INV_X1 u2_u8_u6_U23 (.A( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n170 ) );
  INV_X1 u2_u8_u6_U24 (.A( u2_u8_u6_n113 ) , .ZN( u2_u8_u6_n168 ) );
  AND2_X1 u2_u8_u6_U25 (.A1( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n119 ) , .ZN( u2_u8_u6_n133 ) );
  AND2_X1 u2_u8_u6_U26 (.A2( u2_u8_u6_n121 ) , .A1( u2_u8_u6_n122 ) , .ZN( u2_u8_u6_n131 ) );
  AND3_X1 u2_u8_u6_U27 (.ZN( u2_u8_u6_n120 ) , .A2( u2_u8_u6_n127 ) , .A1( u2_u8_u6_n132 ) , .A3( u2_u8_u6_n145 ) );
  INV_X1 u2_u8_u6_U28 (.A( u2_u8_u6_n146 ) , .ZN( u2_u8_u6_n163 ) );
  AOI222_X1 u2_u8_u6_U29 (.ZN( u2_u8_u6_n114 ) , .A1( u2_u8_u6_n118 ) , .A2( u2_u8_u6_n126 ) , .B2( u2_u8_u6_n151 ) , .C2( u2_u8_u6_n159 ) , .C1( u2_u8_u6_n168 ) , .B1( u2_u8_u6_n169 ) );
  INV_X1 u2_u8_u6_U3 (.A( u2_u8_u6_n110 ) , .ZN( u2_u8_u6_n166 ) );
  NOR2_X1 u2_u8_u6_U30 (.A1( u2_u8_u6_n162 ) , .A2( u2_u8_u6_n165 ) , .ZN( u2_u8_u6_n98 ) );
  AOI211_X1 u2_u8_u6_U31 (.B( u2_u8_u6_n134 ) , .A( u2_u8_u6_n135 ) , .C1( u2_u8_u6_n136 ) , .ZN( u2_u8_u6_n137 ) , .C2( u2_u8_u6_n151 ) );
  AOI21_X1 u2_u8_u6_U32 (.B2( u2_u8_u6_n132 ) , .B1( u2_u8_u6_n133 ) , .ZN( u2_u8_u6_n134 ) , .A( u2_u8_u6_n158 ) );
  NAND4_X1 u2_u8_u6_U33 (.A4( u2_u8_u6_n127 ) , .A3( u2_u8_u6_n128 ) , .A2( u2_u8_u6_n129 ) , .A1( u2_u8_u6_n130 ) , .ZN( u2_u8_u6_n136 ) );
  AOI21_X1 u2_u8_u6_U34 (.B1( u2_u8_u6_n131 ) , .ZN( u2_u8_u6_n135 ) , .A( u2_u8_u6_n144 ) , .B2( u2_u8_u6_n146 ) );
  NAND2_X1 u2_u8_u6_U35 (.A1( u2_u8_u6_n144 ) , .ZN( u2_u8_u6_n151 ) , .A2( u2_u8_u6_n158 ) );
  NAND2_X1 u2_u8_u6_U36 (.ZN( u2_u8_u6_n132 ) , .A1( u2_u8_u6_n91 ) , .A2( u2_u8_u6_n97 ) );
  AOI22_X1 u2_u8_u6_U37 (.B2( u2_u8_u6_n110 ) , .B1( u2_u8_u6_n111 ) , .A1( u2_u8_u6_n112 ) , .ZN( u2_u8_u6_n115 ) , .A2( u2_u8_u6_n161 ) );
  NAND4_X1 u2_u8_u6_U38 (.A3( u2_u8_u6_n109 ) , .ZN( u2_u8_u6_n112 ) , .A4( u2_u8_u6_n132 ) , .A2( u2_u8_u6_n147 ) , .A1( u2_u8_u6_n166 ) );
  NOR2_X1 u2_u8_u6_U39 (.ZN( u2_u8_u6_n109 ) , .A1( u2_u8_u6_n170 ) , .A2( u2_u8_u6_n173 ) );
  INV_X1 u2_u8_u6_U4 (.A( u2_u8_u6_n142 ) , .ZN( u2_u8_u6_n174 ) );
  NOR2_X1 u2_u8_u6_U40 (.A2( u2_u8_u6_n126 ) , .ZN( u2_u8_u6_n155 ) , .A1( u2_u8_u6_n160 ) );
  NAND2_X1 u2_u8_u6_U41 (.ZN( u2_u8_u6_n146 ) , .A2( u2_u8_u6_n94 ) , .A1( u2_u8_u6_n99 ) );
  AOI21_X1 u2_u8_u6_U42 (.A( u2_u8_u6_n144 ) , .B2( u2_u8_u6_n145 ) , .B1( u2_u8_u6_n146 ) , .ZN( u2_u8_u6_n150 ) );
  INV_X1 u2_u8_u6_U43 (.A( u2_u8_u6_n111 ) , .ZN( u2_u8_u6_n158 ) );
  NAND2_X1 u2_u8_u6_U44 (.ZN( u2_u8_u6_n127 ) , .A1( u2_u8_u6_n91 ) , .A2( u2_u8_u6_n92 ) );
  NAND2_X1 u2_u8_u6_U45 (.ZN( u2_u8_u6_n129 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n96 ) );
  INV_X1 u2_u8_u6_U46 (.A( u2_u8_u6_n144 ) , .ZN( u2_u8_u6_n159 ) );
  NAND2_X1 u2_u8_u6_U47 (.ZN( u2_u8_u6_n145 ) , .A2( u2_u8_u6_n97 ) , .A1( u2_u8_u6_n98 ) );
  NAND2_X1 u2_u8_u6_U48 (.ZN( u2_u8_u6_n148 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n94 ) );
  NAND2_X1 u2_u8_u6_U49 (.ZN( u2_u8_u6_n108 ) , .A2( u2_u8_u6_n139 ) , .A1( u2_u8_u6_n144 ) );
  NAND2_X1 u2_u8_u6_U5 (.A2( u2_u8_u6_n143 ) , .ZN( u2_u8_u6_n152 ) , .A1( u2_u8_u6_n166 ) );
  NAND2_X1 u2_u8_u6_U50 (.ZN( u2_u8_u6_n121 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n97 ) );
  NAND2_X1 u2_u8_u6_U51 (.ZN( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n95 ) );
  AND2_X1 u2_u8_u6_U52 (.ZN( u2_u8_u6_n118 ) , .A2( u2_u8_u6_n91 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U53 (.ZN( u2_u8_u6_n147 ) , .A2( u2_u8_u6_n98 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U54 (.ZN( u2_u8_u6_n128 ) , .A1( u2_u8_u6_n94 ) , .A2( u2_u8_u6_n96 ) );
  NAND2_X1 u2_u8_u6_U55 (.ZN( u2_u8_u6_n119 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U56 (.ZN( u2_u8_u6_n123 ) , .A2( u2_u8_u6_n91 ) , .A1( u2_u8_u6_n96 ) );
  NAND2_X1 u2_u8_u6_U57 (.ZN( u2_u8_u6_n100 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n98 ) );
  NAND2_X1 u2_u8_u6_U58 (.ZN( u2_u8_u6_n122 ) , .A1( u2_u8_u6_n94 ) , .A2( u2_u8_u6_n97 ) );
  INV_X1 u2_u8_u6_U59 (.A( u2_u8_u6_n139 ) , .ZN( u2_u8_u6_n160 ) );
  AOI22_X1 u2_u8_u6_U6 (.B2( u2_u8_u6_n101 ) , .A1( u2_u8_u6_n102 ) , .ZN( u2_u8_u6_n103 ) , .B1( u2_u8_u6_n160 ) , .A2( u2_u8_u6_n161 ) );
  NAND2_X1 u2_u8_u6_U60 (.ZN( u2_u8_u6_n113 ) , .A1( u2_u8_u6_n96 ) , .A2( u2_u8_u6_n98 ) );
  NOR2_X1 u2_u8_u6_U61 (.A2( u2_u8_X_40 ) , .A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n126 ) );
  NOR2_X1 u2_u8_u6_U62 (.A2( u2_u8_X_39 ) , .A1( u2_u8_X_42 ) , .ZN( u2_u8_u6_n92 ) );
  NOR2_X1 u2_u8_u6_U63 (.A2( u2_u8_X_39 ) , .A1( u2_u8_u6_n156 ) , .ZN( u2_u8_u6_n97 ) );
  NOR2_X1 u2_u8_u6_U64 (.A2( u2_u8_X_38 ) , .A1( u2_u8_u6_n165 ) , .ZN( u2_u8_u6_n95 ) );
  NOR2_X1 u2_u8_u6_U65 (.A2( u2_u8_X_41 ) , .ZN( u2_u8_u6_n111 ) , .A1( u2_u8_u6_n157 ) );
  NOR2_X1 u2_u8_u6_U66 (.A2( u2_u8_X_37 ) , .A1( u2_u8_u6_n162 ) , .ZN( u2_u8_u6_n94 ) );
  NOR2_X1 u2_u8_u6_U67 (.A2( u2_u8_X_37 ) , .A1( u2_u8_X_38 ) , .ZN( u2_u8_u6_n91 ) );
  NAND2_X1 u2_u8_u6_U68 (.A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n144 ) , .A2( u2_u8_u6_n157 ) );
  NAND2_X1 u2_u8_u6_U69 (.A2( u2_u8_X_40 ) , .A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n139 ) );
  NOR2_X1 u2_u8_u6_U7 (.A1( u2_u8_u6_n118 ) , .ZN( u2_u8_u6_n143 ) , .A2( u2_u8_u6_n168 ) );
  AND2_X1 u2_u8_u6_U70 (.A1( u2_u8_X_39 ) , .A2( u2_u8_u6_n156 ) , .ZN( u2_u8_u6_n96 ) );
  AND2_X1 u2_u8_u6_U71 (.A1( u2_u8_X_39 ) , .A2( u2_u8_X_42 ) , .ZN( u2_u8_u6_n99 ) );
  INV_X1 u2_u8_u6_U72 (.A( u2_u8_X_40 ) , .ZN( u2_u8_u6_n157 ) );
  INV_X1 u2_u8_u6_U73 (.A( u2_u8_X_37 ) , .ZN( u2_u8_u6_n165 ) );
  INV_X1 u2_u8_u6_U74 (.A( u2_u8_X_38 ) , .ZN( u2_u8_u6_n162 ) );
  INV_X1 u2_u8_u6_U75 (.A( u2_u8_X_42 ) , .ZN( u2_u8_u6_n156 ) );
  NAND4_X1 u2_u8_u6_U76 (.ZN( u2_out8_32 ) , .A4( u2_u8_u6_n103 ) , .A3( u2_u8_u6_n104 ) , .A2( u2_u8_u6_n105 ) , .A1( u2_u8_u6_n106 ) );
  AOI22_X1 u2_u8_u6_U77 (.ZN( u2_u8_u6_n105 ) , .A2( u2_u8_u6_n108 ) , .A1( u2_u8_u6_n118 ) , .B2( u2_u8_u6_n126 ) , .B1( u2_u8_u6_n171 ) );
  AOI22_X1 u2_u8_u6_U78 (.ZN( u2_u8_u6_n104 ) , .A1( u2_u8_u6_n111 ) , .B1( u2_u8_u6_n124 ) , .B2( u2_u8_u6_n151 ) , .A2( u2_u8_u6_n93 ) );
  NAND4_X1 u2_u8_u6_U79 (.ZN( u2_out8_12 ) , .A4( u2_u8_u6_n114 ) , .A3( u2_u8_u6_n115 ) , .A2( u2_u8_u6_n116 ) , .A1( u2_u8_u6_n117 ) );
  OAI21_X1 u2_u8_u6_U8 (.A( u2_u8_u6_n159 ) , .B1( u2_u8_u6_n169 ) , .B2( u2_u8_u6_n173 ) , .ZN( u2_u8_u6_n90 ) );
  OAI22_X1 u2_u8_u6_U80 (.B2( u2_u8_u6_n111 ) , .ZN( u2_u8_u6_n116 ) , .B1( u2_u8_u6_n126 ) , .A2( u2_u8_u6_n164 ) , .A1( u2_u8_u6_n167 ) );
  OAI21_X1 u2_u8_u6_U81 (.A( u2_u8_u6_n108 ) , .ZN( u2_u8_u6_n117 ) , .B2( u2_u8_u6_n141 ) , .B1( u2_u8_u6_n163 ) );
  OAI211_X1 u2_u8_u6_U82 (.ZN( u2_out8_7 ) , .B( u2_u8_u6_n153 ) , .C2( u2_u8_u6_n154 ) , .C1( u2_u8_u6_n155 ) , .A( u2_u8_u6_n174 ) );
  NOR3_X1 u2_u8_u6_U83 (.A1( u2_u8_u6_n141 ) , .ZN( u2_u8_u6_n154 ) , .A3( u2_u8_u6_n164 ) , .A2( u2_u8_u6_n171 ) );
  AOI211_X1 u2_u8_u6_U84 (.B( u2_u8_u6_n149 ) , .A( u2_u8_u6_n150 ) , .C2( u2_u8_u6_n151 ) , .C1( u2_u8_u6_n152 ) , .ZN( u2_u8_u6_n153 ) );
  OAI211_X1 u2_u8_u6_U85 (.ZN( u2_out8_22 ) , .B( u2_u8_u6_n137 ) , .A( u2_u8_u6_n138 ) , .C2( u2_u8_u6_n139 ) , .C1( u2_u8_u6_n140 ) );
  AOI22_X1 u2_u8_u6_U86 (.B1( u2_u8_u6_n124 ) , .A2( u2_u8_u6_n125 ) , .A1( u2_u8_u6_n126 ) , .ZN( u2_u8_u6_n138 ) , .B2( u2_u8_u6_n161 ) );
  AND4_X1 u2_u8_u6_U87 (.A3( u2_u8_u6_n119 ) , .A1( u2_u8_u6_n120 ) , .A4( u2_u8_u6_n129 ) , .ZN( u2_u8_u6_n140 ) , .A2( u2_u8_u6_n143 ) );
  NAND3_X1 u2_u8_u6_U88 (.A2( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n125 ) , .A1( u2_u8_u6_n130 ) , .A3( u2_u8_u6_n131 ) );
  NAND3_X1 u2_u8_u6_U89 (.A3( u2_u8_u6_n133 ) , .ZN( u2_u8_u6_n141 ) , .A1( u2_u8_u6_n145 ) , .A2( u2_u8_u6_n148 ) );
  INV_X1 u2_u8_u6_U9 (.ZN( u2_u8_u6_n172 ) , .A( u2_u8_u6_n88 ) );
  NAND3_X1 u2_u8_u6_U90 (.ZN( u2_u8_u6_n101 ) , .A3( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n121 ) , .A1( u2_u8_u6_n127 ) );
  NAND3_X1 u2_u8_u6_U91 (.ZN( u2_u8_u6_n102 ) , .A3( u2_u8_u6_n130 ) , .A2( u2_u8_u6_n145 ) , .A1( u2_u8_u6_n166 ) );
  NAND3_X1 u2_u8_u6_U92 (.A3( u2_u8_u6_n113 ) , .A1( u2_u8_u6_n119 ) , .A2( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n93 ) );
  NAND3_X1 u2_u8_u6_U93 (.ZN( u2_u8_u6_n142 ) , .A2( u2_u8_u6_n172 ) , .A3( u2_u8_u6_n89 ) , .A1( u2_u8_u6_n90 ) );
  AND3_X1 u2_u8_u7_U10 (.A3( u2_u8_u7_n110 ) , .A2( u2_u8_u7_n127 ) , .A1( u2_u8_u7_n132 ) , .ZN( u2_u8_u7_n92 ) );
  OAI21_X1 u2_u8_u7_U11 (.A( u2_u8_u7_n161 ) , .B1( u2_u8_u7_n168 ) , .B2( u2_u8_u7_n173 ) , .ZN( u2_u8_u7_n91 ) );
  AOI211_X1 u2_u8_u7_U12 (.A( u2_u8_u7_n117 ) , .ZN( u2_u8_u7_n118 ) , .C2( u2_u8_u7_n126 ) , .C1( u2_u8_u7_n177 ) , .B( u2_u8_u7_n180 ) );
  OAI22_X1 u2_u8_u7_U13 (.B1( u2_u8_u7_n115 ) , .ZN( u2_u8_u7_n117 ) , .A2( u2_u8_u7_n133 ) , .A1( u2_u8_u7_n137 ) , .B2( u2_u8_u7_n162 ) );
  INV_X1 u2_u8_u7_U14 (.A( u2_u8_u7_n116 ) , .ZN( u2_u8_u7_n180 ) );
  NOR3_X1 u2_u8_u7_U15 (.ZN( u2_u8_u7_n115 ) , .A3( u2_u8_u7_n145 ) , .A2( u2_u8_u7_n168 ) , .A1( u2_u8_u7_n169 ) );
  OAI211_X1 u2_u8_u7_U16 (.B( u2_u8_u7_n122 ) , .A( u2_u8_u7_n123 ) , .C2( u2_u8_u7_n124 ) , .ZN( u2_u8_u7_n154 ) , .C1( u2_u8_u7_n162 ) );
  AOI222_X1 u2_u8_u7_U17 (.ZN( u2_u8_u7_n122 ) , .C2( u2_u8_u7_n126 ) , .C1( u2_u8_u7_n145 ) , .B1( u2_u8_u7_n161 ) , .A2( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n170 ) , .A1( u2_u8_u7_n176 ) );
  INV_X1 u2_u8_u7_U18 (.A( u2_u8_u7_n133 ) , .ZN( u2_u8_u7_n176 ) );
  NOR3_X1 u2_u8_u7_U19 (.A2( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n135 ) , .ZN( u2_u8_u7_n136 ) , .A3( u2_u8_u7_n171 ) );
  NOR2_X1 u2_u8_u7_U20 (.A1( u2_u8_u7_n130 ) , .A2( u2_u8_u7_n134 ) , .ZN( u2_u8_u7_n153 ) );
  INV_X1 u2_u8_u7_U21 (.A( u2_u8_u7_n101 ) , .ZN( u2_u8_u7_n165 ) );
  NOR2_X1 u2_u8_u7_U22 (.ZN( u2_u8_u7_n111 ) , .A2( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n169 ) );
  AOI21_X1 u2_u8_u7_U23 (.ZN( u2_u8_u7_n104 ) , .B2( u2_u8_u7_n112 ) , .B1( u2_u8_u7_n127 ) , .A( u2_u8_u7_n164 ) );
  AOI21_X1 u2_u8_u7_U24 (.ZN( u2_u8_u7_n106 ) , .B1( u2_u8_u7_n133 ) , .B2( u2_u8_u7_n146 ) , .A( u2_u8_u7_n162 ) );
  AOI21_X1 u2_u8_u7_U25 (.A( u2_u8_u7_n101 ) , .ZN( u2_u8_u7_n107 ) , .B2( u2_u8_u7_n128 ) , .B1( u2_u8_u7_n175 ) );
  INV_X1 u2_u8_u7_U26 (.A( u2_u8_u7_n138 ) , .ZN( u2_u8_u7_n171 ) );
  INV_X1 u2_u8_u7_U27 (.A( u2_u8_u7_n131 ) , .ZN( u2_u8_u7_n177 ) );
  INV_X1 u2_u8_u7_U28 (.A( u2_u8_u7_n110 ) , .ZN( u2_u8_u7_n174 ) );
  NAND2_X1 u2_u8_u7_U29 (.A1( u2_u8_u7_n129 ) , .A2( u2_u8_u7_n132 ) , .ZN( u2_u8_u7_n149 ) );
  OAI21_X1 u2_u8_u7_U3 (.ZN( u2_u8_u7_n159 ) , .A( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n171 ) , .B1( u2_u8_u7_n174 ) );
  NAND2_X1 u2_u8_u7_U30 (.A1( u2_u8_u7_n113 ) , .A2( u2_u8_u7_n124 ) , .ZN( u2_u8_u7_n130 ) );
  INV_X1 u2_u8_u7_U31 (.A( u2_u8_u7_n112 ) , .ZN( u2_u8_u7_n173 ) );
  INV_X1 u2_u8_u7_U32 (.A( u2_u8_u7_n128 ) , .ZN( u2_u8_u7_n168 ) );
  INV_X1 u2_u8_u7_U33 (.A( u2_u8_u7_n148 ) , .ZN( u2_u8_u7_n169 ) );
  INV_X1 u2_u8_u7_U34 (.A( u2_u8_u7_n127 ) , .ZN( u2_u8_u7_n179 ) );
  NOR2_X1 u2_u8_u7_U35 (.ZN( u2_u8_u7_n101 ) , .A2( u2_u8_u7_n150 ) , .A1( u2_u8_u7_n156 ) );
  AOI211_X1 u2_u8_u7_U36 (.B( u2_u8_u7_n154 ) , .A( u2_u8_u7_n155 ) , .C1( u2_u8_u7_n156 ) , .ZN( u2_u8_u7_n157 ) , .C2( u2_u8_u7_n172 ) );
  INV_X1 u2_u8_u7_U37 (.A( u2_u8_u7_n153 ) , .ZN( u2_u8_u7_n172 ) );
  AOI211_X1 u2_u8_u7_U38 (.B( u2_u8_u7_n139 ) , .A( u2_u8_u7_n140 ) , .C2( u2_u8_u7_n141 ) , .ZN( u2_u8_u7_n142 ) , .C1( u2_u8_u7_n156 ) );
  NAND4_X1 u2_u8_u7_U39 (.A3( u2_u8_u7_n127 ) , .A2( u2_u8_u7_n128 ) , .A1( u2_u8_u7_n129 ) , .ZN( u2_u8_u7_n141 ) , .A4( u2_u8_u7_n147 ) );
  INV_X1 u2_u8_u7_U4 (.A( u2_u8_u7_n111 ) , .ZN( u2_u8_u7_n170 ) );
  AOI21_X1 u2_u8_u7_U40 (.A( u2_u8_u7_n137 ) , .B1( u2_u8_u7_n138 ) , .ZN( u2_u8_u7_n139 ) , .B2( u2_u8_u7_n146 ) );
  OAI22_X1 u2_u8_u7_U41 (.B1( u2_u8_u7_n136 ) , .ZN( u2_u8_u7_n140 ) , .A1( u2_u8_u7_n153 ) , .B2( u2_u8_u7_n162 ) , .A2( u2_u8_u7_n164 ) );
  AOI21_X1 u2_u8_u7_U42 (.ZN( u2_u8_u7_n123 ) , .B1( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n177 ) , .A( u2_u8_u7_n97 ) );
  AOI21_X1 u2_u8_u7_U43 (.B2( u2_u8_u7_n113 ) , .B1( u2_u8_u7_n124 ) , .A( u2_u8_u7_n125 ) , .ZN( u2_u8_u7_n97 ) );
  INV_X1 u2_u8_u7_U44 (.A( u2_u8_u7_n125 ) , .ZN( u2_u8_u7_n161 ) );
  INV_X1 u2_u8_u7_U45 (.A( u2_u8_u7_n152 ) , .ZN( u2_u8_u7_n162 ) );
  AOI22_X1 u2_u8_u7_U46 (.A2( u2_u8_u7_n114 ) , .ZN( u2_u8_u7_n119 ) , .B1( u2_u8_u7_n130 ) , .A1( u2_u8_u7_n156 ) , .B2( u2_u8_u7_n165 ) );
  NAND2_X1 u2_u8_u7_U47 (.A2( u2_u8_u7_n112 ) , .ZN( u2_u8_u7_n114 ) , .A1( u2_u8_u7_n175 ) );
  AND2_X1 u2_u8_u7_U48 (.ZN( u2_u8_u7_n145 ) , .A2( u2_u8_u7_n98 ) , .A1( u2_u8_u7_n99 ) );
  NOR2_X1 u2_u8_u7_U49 (.ZN( u2_u8_u7_n137 ) , .A1( u2_u8_u7_n150 ) , .A2( u2_u8_u7_n161 ) );
  INV_X1 u2_u8_u7_U5 (.A( u2_u8_u7_n149 ) , .ZN( u2_u8_u7_n175 ) );
  AOI21_X1 u2_u8_u7_U50 (.ZN( u2_u8_u7_n105 ) , .B2( u2_u8_u7_n110 ) , .A( u2_u8_u7_n125 ) , .B1( u2_u8_u7_n147 ) );
  NAND2_X1 u2_u8_u7_U51 (.ZN( u2_u8_u7_n146 ) , .A1( u2_u8_u7_n95 ) , .A2( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U52 (.A2( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n147 ) , .A1( u2_u8_u7_n93 ) );
  NAND2_X1 u2_u8_u7_U53 (.A1( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n127 ) , .A2( u2_u8_u7_n99 ) );
  OR2_X1 u2_u8_u7_U54 (.ZN( u2_u8_u7_n126 ) , .A2( u2_u8_u7_n152 ) , .A1( u2_u8_u7_n156 ) );
  NAND2_X1 u2_u8_u7_U55 (.A2( u2_u8_u7_n102 ) , .A1( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n133 ) );
  NAND2_X1 u2_u8_u7_U56 (.ZN( u2_u8_u7_n112 ) , .A2( u2_u8_u7_n96 ) , .A1( u2_u8_u7_n99 ) );
  NAND2_X1 u2_u8_u7_U57 (.A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n128 ) , .A1( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U58 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n113 ) , .A2( u2_u8_u7_n93 ) );
  NAND2_X1 u2_u8_u7_U59 (.A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n124 ) , .A1( u2_u8_u7_n96 ) );
  INV_X1 u2_u8_u7_U6 (.A( u2_u8_u7_n154 ) , .ZN( u2_u8_u7_n178 ) );
  NAND2_X1 u2_u8_u7_U60 (.ZN( u2_u8_u7_n110 ) , .A1( u2_u8_u7_n95 ) , .A2( u2_u8_u7_n96 ) );
  INV_X1 u2_u8_u7_U61 (.A( u2_u8_u7_n150 ) , .ZN( u2_u8_u7_n164 ) );
  AND2_X1 u2_u8_u7_U62 (.ZN( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n93 ) , .A2( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U63 (.A1( u2_u8_u7_n100 ) , .A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n129 ) );
  NAND2_X1 u2_u8_u7_U64 (.A2( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n131 ) , .A1( u2_u8_u7_n95 ) );
  NAND2_X1 u2_u8_u7_U65 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n138 ) , .A2( u2_u8_u7_n99 ) );
  NAND2_X1 u2_u8_u7_U66 (.ZN( u2_u8_u7_n132 ) , .A1( u2_u8_u7_n93 ) , .A2( u2_u8_u7_n96 ) );
  NAND2_X1 u2_u8_u7_U67 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n148 ) , .A2( u2_u8_u7_n95 ) );
  NOR2_X1 u2_u8_u7_U68 (.A2( u2_u8_X_47 ) , .ZN( u2_u8_u7_n150 ) , .A1( u2_u8_u7_n163 ) );
  NOR2_X1 u2_u8_u7_U69 (.A2( u2_u8_X_43 ) , .A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n103 ) );
  AOI211_X1 u2_u8_u7_U7 (.ZN( u2_u8_u7_n116 ) , .A( u2_u8_u7_n155 ) , .C1( u2_u8_u7_n161 ) , .C2( u2_u8_u7_n171 ) , .B( u2_u8_u7_n94 ) );
  NOR2_X1 u2_u8_u7_U70 (.A2( u2_u8_X_48 ) , .A1( u2_u8_u7_n166 ) , .ZN( u2_u8_u7_n95 ) );
  NOR2_X1 u2_u8_u7_U71 (.A2( u2_u8_X_45 ) , .A1( u2_u8_X_48 ) , .ZN( u2_u8_u7_n99 ) );
  NOR2_X1 u2_u8_u7_U72 (.A2( u2_u8_X_44 ) , .A1( u2_u8_u7_n167 ) , .ZN( u2_u8_u7_n98 ) );
  NOR2_X1 u2_u8_u7_U73 (.A2( u2_u8_X_46 ) , .A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n152 ) );
  AND2_X1 u2_u8_u7_U74 (.A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n156 ) , .A2( u2_u8_u7_n163 ) );
  NAND2_X1 u2_u8_u7_U75 (.A2( u2_u8_X_46 ) , .A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n125 ) );
  AND2_X1 u2_u8_u7_U76 (.A2( u2_u8_X_45 ) , .A1( u2_u8_X_48 ) , .ZN( u2_u8_u7_n102 ) );
  AND2_X1 u2_u8_u7_U77 (.A2( u2_u8_X_43 ) , .A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n96 ) );
  AND2_X1 u2_u8_u7_U78 (.A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n100 ) , .A2( u2_u8_u7_n167 ) );
  AND2_X1 u2_u8_u7_U79 (.A1( u2_u8_X_48 ) , .A2( u2_u8_u7_n166 ) , .ZN( u2_u8_u7_n93 ) );
  OAI222_X1 u2_u8_u7_U8 (.C2( u2_u8_u7_n101 ) , .B2( u2_u8_u7_n111 ) , .A1( u2_u8_u7_n113 ) , .C1( u2_u8_u7_n146 ) , .A2( u2_u8_u7_n162 ) , .B1( u2_u8_u7_n164 ) , .ZN( u2_u8_u7_n94 ) );
  INV_X1 u2_u8_u7_U80 (.A( u2_u8_X_46 ) , .ZN( u2_u8_u7_n163 ) );
  INV_X1 u2_u8_u7_U81 (.A( u2_u8_X_43 ) , .ZN( u2_u8_u7_n167 ) );
  INV_X1 u2_u8_u7_U82 (.A( u2_u8_X_45 ) , .ZN( u2_u8_u7_n166 ) );
  NAND4_X1 u2_u8_u7_U83 (.ZN( u2_out8_27 ) , .A4( u2_u8_u7_n118 ) , .A3( u2_u8_u7_n119 ) , .A2( u2_u8_u7_n120 ) , .A1( u2_u8_u7_n121 ) );
  OAI21_X1 u2_u8_u7_U84 (.ZN( u2_u8_u7_n121 ) , .B2( u2_u8_u7_n145 ) , .A( u2_u8_u7_n150 ) , .B1( u2_u8_u7_n174 ) );
  OAI21_X1 u2_u8_u7_U85 (.ZN( u2_u8_u7_n120 ) , .A( u2_u8_u7_n161 ) , .B2( u2_u8_u7_n170 ) , .B1( u2_u8_u7_n179 ) );
  NAND4_X1 u2_u8_u7_U86 (.ZN( u2_out8_21 ) , .A4( u2_u8_u7_n157 ) , .A3( u2_u8_u7_n158 ) , .A2( u2_u8_u7_n159 ) , .A1( u2_u8_u7_n160 ) );
  OAI21_X1 u2_u8_u7_U87 (.B1( u2_u8_u7_n145 ) , .ZN( u2_u8_u7_n160 ) , .A( u2_u8_u7_n161 ) , .B2( u2_u8_u7_n177 ) );
  AOI22_X1 u2_u8_u7_U88 (.B2( u2_u8_u7_n149 ) , .B1( u2_u8_u7_n150 ) , .A2( u2_u8_u7_n151 ) , .A1( u2_u8_u7_n152 ) , .ZN( u2_u8_u7_n158 ) );
  NAND4_X1 u2_u8_u7_U89 (.ZN( u2_out8_15 ) , .A4( u2_u8_u7_n142 ) , .A3( u2_u8_u7_n143 ) , .A2( u2_u8_u7_n144 ) , .A1( u2_u8_u7_n178 ) );
  OAI221_X1 u2_u8_u7_U9 (.C1( u2_u8_u7_n101 ) , .C2( u2_u8_u7_n147 ) , .ZN( u2_u8_u7_n155 ) , .B2( u2_u8_u7_n162 ) , .A( u2_u8_u7_n91 ) , .B1( u2_u8_u7_n92 ) );
  OR2_X1 u2_u8_u7_U90 (.A2( u2_u8_u7_n125 ) , .A1( u2_u8_u7_n129 ) , .ZN( u2_u8_u7_n144 ) );
  AOI22_X1 u2_u8_u7_U91 (.A2( u2_u8_u7_n126 ) , .ZN( u2_u8_u7_n143 ) , .B2( u2_u8_u7_n165 ) , .B1( u2_u8_u7_n173 ) , .A1( u2_u8_u7_n174 ) );
  NAND4_X1 u2_u8_u7_U92 (.ZN( u2_out8_5 ) , .A4( u2_u8_u7_n108 ) , .A3( u2_u8_u7_n109 ) , .A1( u2_u8_u7_n116 ) , .A2( u2_u8_u7_n123 ) );
  AOI22_X1 u2_u8_u7_U93 (.ZN( u2_u8_u7_n109 ) , .A2( u2_u8_u7_n126 ) , .B2( u2_u8_u7_n145 ) , .B1( u2_u8_u7_n156 ) , .A1( u2_u8_u7_n171 ) );
  NOR4_X1 u2_u8_u7_U94 (.A4( u2_u8_u7_n104 ) , .A3( u2_u8_u7_n105 ) , .A2( u2_u8_u7_n106 ) , .A1( u2_u8_u7_n107 ) , .ZN( u2_u8_u7_n108 ) );
  NAND3_X1 u2_u8_u7_U95 (.A3( u2_u8_u7_n146 ) , .A2( u2_u8_u7_n147 ) , .A1( u2_u8_u7_n148 ) , .ZN( u2_u8_u7_n151 ) );
  NAND3_X1 u2_u8_u7_U96 (.A3( u2_u8_u7_n131 ) , .A2( u2_u8_u7_n132 ) , .A1( u2_u8_u7_n133 ) , .ZN( u2_u8_u7_n135 ) );
  OAI21_X1 u2_uk_U1013 (.ZN( u2_K9_44 ) , .A( u2_uk_n1138 ) , .B2( u2_uk_n1585 ) , .B1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U1014 (.A1( u2_uk_K_r7_0 ) , .ZN( u2_uk_n1138 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1088 (.ZN( u2_K8_3 ) , .A( u2_uk_n1110 ) );
  INV_X1 u2_uk_U1096 (.ZN( u2_K11_12 ) , .A( u2_uk_n313 ) );
  INV_X1 u2_uk_U1098 (.ZN( u2_K8_12 ) , .A( u2_uk_n1098 ) );
  INV_X1 u2_uk_U1139 (.ZN( u2_K8_43 ) , .A( u2_uk_n1113 ) );
  INV_X1 u2_uk_U177 (.ZN( u2_K11_14 ) , .A( u2_uk_n319 ) );
  INV_X1 u2_uk_U262 (.ZN( u2_K9_48 ) , .A( u2_uk_n1140 ) );
  INV_X1 u2_uk_U441 (.ZN( u2_K16_37 ) , .A( u2_uk_n959 ) );
  INV_X1 u2_uk_U444 (.ZN( u2_K9_33 ) , .A( u2_uk_n1132 ) );
  INV_X1 u2_uk_U481 (.ZN( u2_K16_29 ) , .A( u2_uk_n955 ) );
  INV_X1 u2_uk_U52 (.ZN( u2_K16_34 ) , .A( u2_uk_n958 ) );
  INV_X1 u2_uk_U544 (.ZN( u2_K11_17 ) , .A( u2_uk_n335 ) );
  INV_X1 u2_uk_U616 (.ZN( u2_K9_35 ) , .A( u2_uk_n1133 ) );
  INV_X1 u2_uk_U661 (.ZN( u2_K16_43 ) , .A( u2_uk_n963 ) );
  INV_X1 u2_uk_U968 (.ZN( u2_K9_41 ) , .A( u2_uk_n1136 ) );
  INV_X1 u2_uk_U972 (.ZN( u2_K9_42 ) , .A( u2_uk_n1137 ) );
endmodule

