module des_des_die_8 ( n116, u0_K10_25, u0_K10_27, u0_K10_32, u0_K10_34, u0_K10_36, u0_K14_10, u0_K14_12, u0_K14_13, 
       u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_21, u0_K14_24, u0_K14_27, u0_K14_9, u0_L12_1, u0_L12_10, 
       u0_L12_13, u0_L12_14, u0_L12_16, u0_L12_18, u0_L12_2, u0_L12_20, u0_L12_24, u0_L12_25, u0_L12_26, 
       u0_L12_28, u0_L12_3, u0_L12_30, u0_L12_6, u0_L12_8, u0_L8_11, u0_L8_14, u0_L8_15, u0_L8_19, 
       u0_L8_21, u0_L8_25, u0_L8_27, u0_L8_29, u0_L8_3, u0_L8_4, u0_L8_5, u0_L8_8, u0_R12_10, 
       u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, u0_R12_16, u0_R12_17, u0_R12_18, u0_R12_19, 
       u0_R12_20, u0_R12_21, u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R8_1, 
       u0_R8_16, u0_R8_17, u0_R8_18, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_23, u0_R8_24, 
       u0_R8_25, u0_R8_28, u0_R8_29, u0_R8_30, u0_R8_31, u0_R8_32, u0_uk_K_r12_25, u0_uk_K_r12_33, u0_uk_K_r12_44, 
       u0_uk_K_r8_16, u0_uk_K_r8_2, u0_uk_K_r8_37, u0_uk_n100, u0_uk_n1012, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, 
       u0_uk_n117, u0_uk_n118, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n162, u0_uk_n164, 
       u0_uk_n17, u0_uk_n182, u0_uk_n188, u0_uk_n203, u0_uk_n207, u0_uk_n213, u0_uk_n214, u0_uk_n222, u0_uk_n223, 
       u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n237, u0_uk_n240, u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n247, 
       u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n256, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n265, u0_uk_n46, 
       u0_uk_n48, u0_uk_n49, u0_uk_n50, u0_uk_n51, u0_uk_n53, u0_uk_n54, u0_uk_n61, u0_uk_n66, u0_uk_n67, 
       u0_uk_n69, u0_uk_n72, u0_uk_n75, u0_uk_n77, u0_uk_n78, u0_uk_n79, u0_uk_n80, u0_uk_n82, u0_uk_n83, 
       u0_uk_n84, u0_uk_n86, u0_uk_n87, u0_uk_n88, u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_L13_11, u1_L13_12, 
       u1_L13_15, u1_L13_19, u1_L13_21, u1_L13_22, u1_L13_27, u1_L13_29, u1_L13_32, u1_L13_4, u1_L13_5, 
       u1_L13_7, u1_L2_13, u1_L2_18, u1_L2_2, u1_L2_28, u1_L3_11, u1_L3_19, u1_L3_29, u1_L3_4, 
       u1_L4_1, u1_L4_10, u1_L4_11, u1_L4_12, u1_L4_14, u1_L4_16, u1_L4_17, u1_L4_19, u1_L4_20, 
       u1_L4_22, u1_L4_23, u1_L4_24, u1_L4_25, u1_L4_26, u1_L4_29, u1_L4_3, u1_L4_30, u1_L4_31, 
       u1_L4_32, u1_L4_4, u1_L4_6, u1_L4_7, u1_L4_8, u1_L4_9, u1_L7_1, u1_L7_10, u1_L7_13, 
       u1_L7_16, u1_L7_17, u1_L7_18, u1_L7_2, u1_L7_20, u1_L7_23, u1_L7_24, u1_L7_26, u1_L7_28, 
       u1_L7_30, u1_L7_31, u1_L7_6, u1_L7_9, u1_L8_15, u1_L8_21, u1_L8_27, u1_L8_5, u1_R13_1, 
       u1_R13_20, u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, u1_R13_28, 
       u1_R13_29, u1_R13_30, u1_R13_31, u1_R13_32, u1_R2_4, u1_R2_5, u1_R2_6, u1_R2_7, u1_R2_8, 
       u1_R2_9, u1_R3_20, u1_R3_21, u1_R3_22, u1_R3_23, u1_R3_24, u1_R3_25, u1_R4_1, u1_R4_10, 
       u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, u1_R4_16, u1_R4_17, u1_R4_18, u1_R4_19, 
       u1_R4_2, u1_R4_20, u1_R4_21, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, u1_R4_27, 
       u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_8, u1_R4_9, u1_R7_1, 
       u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_2, 
       u1_R7_3, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, 
       u1_R8_28, u1_R8_29, u1_R8_30, u1_R8_31, u1_R8_32, u1_desIn_r_0, u1_desIn_r_1, u1_desIn_r_11, u1_desIn_r_16, 
       u1_desIn_r_17, u1_desIn_r_18, u1_desIn_r_19, u1_desIn_r_20, u1_desIn_r_22, u1_desIn_r_25, u1_desIn_r_27, u1_desIn_r_28, u1_desIn_r_3, 
       u1_desIn_r_30, u1_desIn_r_32, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_38, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_43, 
       u1_desIn_r_44, u1_desIn_r_49, u1_desIn_r_51, u1_desIn_r_52, u1_desIn_r_54, u1_desIn_r_56, u1_desIn_r_57, u1_desIn_r_59, u1_desIn_r_61, 
       u1_desIn_r_62, u1_desIn_r_7, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_2, 
       u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_28, u1_key_r_29, u1_key_r_30, u1_key_r_31, u1_key_r_35, u1_key_r_36, 
       u1_key_r_37, u1_key_r_38, u1_key_r_42, u1_key_r_43, u1_key_r_44, u1_key_r_45, u1_key_r_49, u1_key_r_50, u1_key_r_51, 
       u1_key_r_52, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r13_2, u1_uk_K_r13_23, u1_uk_K_r13_31, u1_uk_K_r13_35, u1_uk_K_r13_36, 
       u1_uk_K_r13_44, u1_uk_K_r2_26, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_6, u1_uk_K_r3_14, u1_uk_K_r3_29, u1_uk_K_r3_38, u1_uk_K_r3_44, 
       u1_uk_K_r3_52, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_27, u1_uk_K_r4_31, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, 
       u1_uk_K_r4_41, u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_55, u1_uk_K_r7_13, u1_uk_K_r7_20, u1_uk_K_r7_24, 
       u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_32, u1_uk_K_r7_34, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, 
       u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, 
       u1_uk_n110, u1_uk_n117, u1_uk_n118, u1_uk_n128, u1_uk_n129, u1_uk_n1353, u1_uk_n1357, u1_uk_n1359, u1_uk_n1363, 
       u1_uk_n1369, u1_uk_n1371, u1_uk_n1391, u1_uk_n1401, u1_uk_n1408, u1_uk_n1412, u1_uk_n1414, u1_uk_n142, u1_uk_n1431, 
       u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, 
       u1_uk_n1448, u1_uk_n1449, u1_uk_n145, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, 
       u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n146, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, 
       u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, u1_uk_n147, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, 
       u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n148, u1_uk_n155, u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, 
       u1_uk_n1578, u1_uk_n1579, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1592, u1_uk_n1593, u1_uk_n1598, u1_uk_n1603, 
       u1_uk_n1604, u1_uk_n161, u1_uk_n1610, u1_uk_n1616, u1_uk_n162, u1_uk_n1623, u1_uk_n1624, u1_uk_n1627, u1_uk_n1628, 
       u1_uk_n163, u1_uk_n1632, u1_uk_n1639, u1_uk_n164, u1_uk_n1640, u1_uk_n1641, u1_uk_n1644, u1_uk_n1647, u1_uk_n1651, 
       u1_uk_n1656, u1_uk_n17, u1_uk_n182, u1_uk_n1843, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1854, u1_uk_n1855, 
       u1_uk_n1856, u1_uk_n1860, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, u1_uk_n187, u1_uk_n1870, u1_uk_n1875, u1_uk_n1876, 
       u1_uk_n1879, u1_uk_n188, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n191, u1_uk_n202, u1_uk_n203, 
       u1_uk_n207, u1_uk_n208, u1_uk_n209, u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n230, 
       u1_uk_n231, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, 
       u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, 
       u1_uk_n31, u1_uk_n83, u1_uk_n92, u1_uk_n93, u1_uk_n94, u1_uk_n99, u2_K2_16, u2_K2_18, u2_K9_32, 
       u2_K9_36, u2_K9_38, u2_K9_40, u2_L0_16, u2_L0_24, u2_L0_30, u2_L0_6, u2_L7_11, u2_L7_12, 
       u2_L7_19, u2_L7_22, u2_L7_29, u2_L7_32, u2_L7_4, u2_L7_7, u2_R0_10, u2_R0_11, u2_R0_12, 
       u2_R0_13, u2_R0_8, u2_R0_9, u2_R7_20, u2_R7_21, u2_R7_22, u2_R7_23, u2_R7_24, u2_R7_25, 
       u2_R7_26, u2_R7_27, u2_R7_28, u2_R7_29, u2_uk_K_r0_11, u2_uk_K_r0_32, u2_uk_K_r7_16, u2_uk_K_r7_23, u2_uk_K_r7_31, 
       u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n1132, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n118, 
       u2_uk_n1231, u2_uk_n1247, u2_uk_n1260, u2_uk_n1261, u2_uk_n142, u2_uk_n145, u2_uk_n148, u2_uk_n1542, u2_uk_n1551, 
       u2_uk_n1558, u2_uk_n1571, u2_uk_n1583, u2_uk_n161, u2_uk_n162, u2_uk_n230, u2_uk_n94, u2_uk_n99, u2_uk_n994, u0_N290, u0_N291, u0_N292, u0_N295, u0_N298, u0_N301, u0_N302, u0_N306, u0_N308, 
        u0_N312, u0_N314, u0_N316, u0_N416, u0_N417, u0_N418, u0_N421, u0_N423, u0_N425, 
        u0_N428, u0_N429, u0_N431, u0_N433, u0_N435, u0_N439, u0_N440, u0_N441, u0_N443, 
        u0_N445, u1_N10, u1_N108, u1_N11, u1_N113, u1_N123, u1_N13, u1_N131, u1_N138, 
        u1_N14, u1_N146, u1_N156, u1_N160, u1_N162, u1_N163, u1_N165, u1_N166, u1_N167, 
        u1_N168, u1_N169, u1_N170, u1_N171, u1_N173, u1_N175, u1_N176, u1_N178, u1_N179, 
        u1_N18, u1_N181, u1_N182, u1_N183, u1_N184, u1_N185, u1_N188, u1_N189, u1_N190, 
        u1_N191, u1_N2, u1_N20, u1_N21, u1_N24, u1_N256, u1_N257, u1_N26, u1_N261, 
        u1_N264, u1_N265, u1_N268, u1_N271, u1_N272, u1_N273, u1_N275, u1_N278, u1_N279, 
        u1_N28, u1_N281, u1_N283, u1_N285, u1_N286, u1_N292, u1_N3, u1_N302, u1_N308, 
        u1_N31, u1_N314, u1_N4, u1_N451, u1_N452, u1_N454, u1_N458, u1_N459, u1_N462, 
        u1_N466, u1_N468, u1_N469, u1_N474, u1_N476, u1_N479, u1_N6, u1_N7, u1_N97, 
        u1_uk_n213, u1_uk_n60, u2_N259, u2_N262, u2_N266, u2_N267, u2_N274, u2_N277, u2_N284, 
        u2_N287, u2_N37, u2_N47, u2_N55, u2_N61 );
  input n116, u0_K10_25, u0_K10_27, u0_K10_32, u0_K10_34, u0_K10_36, u0_K14_10, u0_K14_12, u0_K14_13, 
        u0_K14_14, u0_K14_15, u0_K14_18, u0_K14_21, u0_K14_24, u0_K14_27, u0_K14_9, u0_L12_1, u0_L12_10, 
        u0_L12_13, u0_L12_14, u0_L12_16, u0_L12_18, u0_L12_2, u0_L12_20, u0_L12_24, u0_L12_25, u0_L12_26, 
        u0_L12_28, u0_L12_3, u0_L12_30, u0_L12_6, u0_L12_8, u0_L8_11, u0_L8_14, u0_L8_15, u0_L8_19, 
        u0_L8_21, u0_L8_25, u0_L8_27, u0_L8_29, u0_L8_3, u0_L8_4, u0_L8_5, u0_L8_8, u0_R12_10, 
        u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, u0_R12_16, u0_R12_17, u0_R12_18, u0_R12_19, 
        u0_R12_20, u0_R12_21, u0_R12_4, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R8_1, 
        u0_R8_16, u0_R8_17, u0_R8_18, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, u0_R8_23, u0_R8_24, 
        u0_R8_25, u0_R8_28, u0_R8_29, u0_R8_30, u0_R8_31, u0_R8_32, u0_uk_K_r12_25, u0_uk_K_r12_33, u0_uk_K_r12_44, 
        u0_uk_K_r8_16, u0_uk_K_r8_2, u0_uk_K_r8_37, u0_uk_n100, u0_uk_n1012, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, 
        u0_uk_n117, u0_uk_n118, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n162, u0_uk_n164, 
        u0_uk_n17, u0_uk_n182, u0_uk_n188, u0_uk_n203, u0_uk_n207, u0_uk_n213, u0_uk_n214, u0_uk_n222, u0_uk_n223, 
        u0_uk_n231, u0_uk_n232, u0_uk_n233, u0_uk_n237, u0_uk_n240, u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n247, 
        u0_uk_n248, u0_uk_n249, u0_uk_n250, u0_uk_n256, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n265, u0_uk_n46, 
        u0_uk_n48, u0_uk_n49, u0_uk_n50, u0_uk_n51, u0_uk_n53, u0_uk_n54, u0_uk_n61, u0_uk_n66, u0_uk_n67, 
        u0_uk_n69, u0_uk_n72, u0_uk_n75, u0_uk_n77, u0_uk_n78, u0_uk_n79, u0_uk_n80, u0_uk_n82, u0_uk_n83, 
        u0_uk_n84, u0_uk_n86, u0_uk_n87, u0_uk_n88, u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_L13_11, u1_L13_12, 
        u1_L13_15, u1_L13_19, u1_L13_21, u1_L13_22, u1_L13_27, u1_L13_29, u1_L13_32, u1_L13_4, u1_L13_5, 
        u1_L13_7, u1_L2_13, u1_L2_18, u1_L2_2, u1_L2_28, u1_L3_11, u1_L3_19, u1_L3_29, u1_L3_4, 
        u1_L4_1, u1_L4_10, u1_L4_11, u1_L4_12, u1_L4_14, u1_L4_16, u1_L4_17, u1_L4_19, u1_L4_20, 
        u1_L4_22, u1_L4_23, u1_L4_24, u1_L4_25, u1_L4_26, u1_L4_29, u1_L4_3, u1_L4_30, u1_L4_31, 
        u1_L4_32, u1_L4_4, u1_L4_6, u1_L4_7, u1_L4_8, u1_L4_9, u1_L7_1, u1_L7_10, u1_L7_13, 
        u1_L7_16, u1_L7_17, u1_L7_18, u1_L7_2, u1_L7_20, u1_L7_23, u1_L7_24, u1_L7_26, u1_L7_28, 
        u1_L7_30, u1_L7_31, u1_L7_6, u1_L7_9, u1_L8_15, u1_L8_21, u1_L8_27, u1_L8_5, u1_R13_1, 
        u1_R13_20, u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, u1_R13_27, u1_R13_28, 
        u1_R13_29, u1_R13_30, u1_R13_31, u1_R13_32, u1_R2_4, u1_R2_5, u1_R2_6, u1_R2_7, u1_R2_8, 
        u1_R2_9, u1_R3_20, u1_R3_21, u1_R3_22, u1_R3_23, u1_R3_24, u1_R3_25, u1_R4_1, u1_R4_10, 
        u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, u1_R4_16, u1_R4_17, u1_R4_18, u1_R4_19, 
        u1_R4_2, u1_R4_20, u1_R4_21, u1_R4_22, u1_R4_23, u1_R4_24, u1_R4_25, u1_R4_26, u1_R4_27, 
        u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_8, u1_R4_9, u1_R7_1, 
        u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_2, 
        u1_R7_3, u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, 
        u1_R8_28, u1_R8_29, u1_R8_30, u1_R8_31, u1_R8_32, u1_desIn_r_0, u1_desIn_r_1, u1_desIn_r_11, u1_desIn_r_16, 
        u1_desIn_r_17, u1_desIn_r_18, u1_desIn_r_19, u1_desIn_r_20, u1_desIn_r_22, u1_desIn_r_25, u1_desIn_r_27, u1_desIn_r_28, u1_desIn_r_3, 
        u1_desIn_r_30, u1_desIn_r_32, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_38, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_43, 
        u1_desIn_r_44, u1_desIn_r_49, u1_desIn_r_51, u1_desIn_r_52, u1_desIn_r_54, u1_desIn_r_56, u1_desIn_r_57, u1_desIn_r_59, u1_desIn_r_61, 
        u1_desIn_r_62, u1_desIn_r_7, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_2, 
        u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_28, u1_key_r_29, u1_key_r_30, u1_key_r_31, u1_key_r_35, u1_key_r_36, 
        u1_key_r_37, u1_key_r_38, u1_key_r_42, u1_key_r_43, u1_key_r_44, u1_key_r_45, u1_key_r_49, u1_key_r_50, u1_key_r_51, 
        u1_key_r_52, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r13_2, u1_uk_K_r13_23, u1_uk_K_r13_31, u1_uk_K_r13_35, u1_uk_K_r13_36, 
        u1_uk_K_r13_44, u1_uk_K_r2_26, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_6, u1_uk_K_r3_14, u1_uk_K_r3_29, u1_uk_K_r3_38, u1_uk_K_r3_44, 
        u1_uk_K_r3_52, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_27, u1_uk_K_r4_31, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, 
        u1_uk_K_r4_41, u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_55, u1_uk_K_r7_13, u1_uk_K_r7_20, u1_uk_K_r7_24, 
        u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_32, u1_uk_K_r7_34, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, 
        u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, 
        u1_uk_n110, u1_uk_n117, u1_uk_n118, u1_uk_n128, u1_uk_n129, u1_uk_n1353, u1_uk_n1357, u1_uk_n1359, u1_uk_n1363, 
        u1_uk_n1369, u1_uk_n1371, u1_uk_n1391, u1_uk_n1401, u1_uk_n1408, u1_uk_n1412, u1_uk_n1414, u1_uk_n142, u1_uk_n1431, 
        u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, 
        u1_uk_n1448, u1_uk_n1449, u1_uk_n145, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, 
        u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n146, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, 
        u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, u1_uk_n147, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, 
        u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n148, u1_uk_n155, u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, 
        u1_uk_n1578, u1_uk_n1579, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1592, u1_uk_n1593, u1_uk_n1598, u1_uk_n1603, 
        u1_uk_n1604, u1_uk_n161, u1_uk_n1610, u1_uk_n1616, u1_uk_n162, u1_uk_n1623, u1_uk_n1624, u1_uk_n1627, u1_uk_n1628, 
        u1_uk_n163, u1_uk_n1632, u1_uk_n1639, u1_uk_n164, u1_uk_n1640, u1_uk_n1641, u1_uk_n1644, u1_uk_n1647, u1_uk_n1651, 
        u1_uk_n1656, u1_uk_n17, u1_uk_n182, u1_uk_n1843, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1854, u1_uk_n1855, 
        u1_uk_n1856, u1_uk_n1860, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, u1_uk_n187, u1_uk_n1870, u1_uk_n1875, u1_uk_n1876, 
        u1_uk_n1879, u1_uk_n188, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n191, u1_uk_n202, u1_uk_n203, 
        u1_uk_n207, u1_uk_n208, u1_uk_n209, u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n230, 
        u1_uk_n231, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, 
        u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, 
        u1_uk_n31, u1_uk_n83, u1_uk_n92, u1_uk_n93, u1_uk_n94, u1_uk_n99, u2_K2_16, u2_K2_18, u2_K9_32, 
        u2_K9_36, u2_K9_38, u2_K9_40, u2_L0_16, u2_L0_24, u2_L0_30, u2_L0_6, u2_L7_11, u2_L7_12, 
        u2_L7_19, u2_L7_22, u2_L7_29, u2_L7_32, u2_L7_4, u2_L7_7, u2_R0_10, u2_R0_11, u2_R0_12, 
        u2_R0_13, u2_R0_8, u2_R0_9, u2_R7_20, u2_R7_21, u2_R7_22, u2_R7_23, u2_R7_24, u2_R7_25, 
        u2_R7_26, u2_R7_27, u2_R7_28, u2_R7_29, u2_uk_K_r0_11, u2_uk_K_r0_32, u2_uk_K_r7_16, u2_uk_K_r7_23, u2_uk_K_r7_31, 
        u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n1132, u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n118, 
        u2_uk_n1231, u2_uk_n1247, u2_uk_n1260, u2_uk_n1261, u2_uk_n142, u2_uk_n145, u2_uk_n148, u2_uk_n1542, u2_uk_n1551, 
        u2_uk_n1558, u2_uk_n1571, u2_uk_n1583, u2_uk_n161, u2_uk_n162, u2_uk_n230, u2_uk_n94, u2_uk_n99, u2_uk_n994;
  output u0_N290, u0_N291, u0_N292, u0_N295, u0_N298, u0_N301, u0_N302, u0_N306, u0_N308, 
        u0_N312, u0_N314, u0_N316, u0_N416, u0_N417, u0_N418, u0_N421, u0_N423, u0_N425, 
        u0_N428, u0_N429, u0_N431, u0_N433, u0_N435, u0_N439, u0_N440, u0_N441, u0_N443, 
        u0_N445, u1_N10, u1_N108, u1_N11, u1_N113, u1_N123, u1_N13, u1_N131, u1_N138, 
        u1_N14, u1_N146, u1_N156, u1_N160, u1_N162, u1_N163, u1_N165, u1_N166, u1_N167, 
        u1_N168, u1_N169, u1_N170, u1_N171, u1_N173, u1_N175, u1_N176, u1_N178, u1_N179, 
        u1_N18, u1_N181, u1_N182, u1_N183, u1_N184, u1_N185, u1_N188, u1_N189, u1_N190, 
        u1_N191, u1_N2, u1_N20, u1_N21, u1_N24, u1_N256, u1_N257, u1_N26, u1_N261, 
        u1_N264, u1_N265, u1_N268, u1_N271, u1_N272, u1_N273, u1_N275, u1_N278, u1_N279, 
        u1_N28, u1_N281, u1_N283, u1_N285, u1_N286, u1_N292, u1_N3, u1_N302, u1_N308, 
        u1_N31, u1_N314, u1_N4, u1_N451, u1_N452, u1_N454, u1_N458, u1_N459, u1_N462, 
        u1_N466, u1_N468, u1_N469, u1_N474, u1_N476, u1_N479, u1_N6, u1_N7, u1_N97, 
        u1_uk_n213, u1_uk_n60, u2_N259, u2_N262, u2_N266, u2_N267, u2_N274, u2_N277, u2_N284, 
        u2_N287, u2_N37, u2_N47, u2_N55, u2_N61;
  wire u0_K10_26, u0_K10_28, u0_K10_29, u0_K10_30, u0_K10_31, u0_K10_33, u0_K10_35, u0_K10_43, u0_K10_44, 
       u0_K10_45, u0_K10_46, u0_K10_47, u0_K10_48, u0_K14_11, u0_K14_16, u0_K14_17, u0_K14_19, u0_K14_20, 
       u0_K14_22, u0_K14_23, u0_K14_25, u0_K14_26, u0_K14_28, u0_K14_29, u0_K14_30, u0_K14_7, u0_K14_8, 
       u0_out13_1, u0_out13_10, u0_out13_13, u0_out13_14, u0_out13_16, u0_out13_18, u0_out13_2, u0_out13_20, u0_out13_24, 
       u0_out13_25, u0_out13_26, u0_out13_28, u0_out13_3, u0_out13_30, u0_out13_6, u0_out13_8, u0_out9_11, u0_out9_14, 
       u0_out9_15, u0_out9_19, u0_out9_21, u0_out9_25, u0_out9_27, u0_out9_29, u0_out9_3, u0_out9_4, u0_out9_5, 
       u0_out9_8, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_13, u0_u13_X_14, u0_u13_X_15, u0_u13_X_16, u0_u13_X_17, 
       u0_u13_X_18, u0_u13_X_19, u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_23, u0_u13_X_24, u0_u13_X_25, u0_u13_X_26, 
       u0_u13_X_27, u0_u13_X_28, u0_u13_X_29, u0_u13_X_30, u0_u13_X_7, u0_u13_X_8, u0_u13_X_9, u0_u13_u1_n100, u0_u13_u1_n101, 
       u0_u13_u1_n102, u0_u13_u1_n103, u0_u13_u1_n104, u0_u13_u1_n105, u0_u13_u1_n106, u0_u13_u1_n107, u0_u13_u1_n108, u0_u13_u1_n109, u0_u13_u1_n110, 
       u0_u13_u1_n111, u0_u13_u1_n112, u0_u13_u1_n113, u0_u13_u1_n114, u0_u13_u1_n115, u0_u13_u1_n116, u0_u13_u1_n117, u0_u13_u1_n118, u0_u13_u1_n119, 
       u0_u13_u1_n120, u0_u13_u1_n121, u0_u13_u1_n122, u0_u13_u1_n123, u0_u13_u1_n124, u0_u13_u1_n125, u0_u13_u1_n126, u0_u13_u1_n127, u0_u13_u1_n128, 
       u0_u13_u1_n129, u0_u13_u1_n130, u0_u13_u1_n131, u0_u13_u1_n132, u0_u13_u1_n133, u0_u13_u1_n134, u0_u13_u1_n135, u0_u13_u1_n136, u0_u13_u1_n137, 
       u0_u13_u1_n138, u0_u13_u1_n139, u0_u13_u1_n140, u0_u13_u1_n141, u0_u13_u1_n142, u0_u13_u1_n143, u0_u13_u1_n144, u0_u13_u1_n145, u0_u13_u1_n146, 
       u0_u13_u1_n147, u0_u13_u1_n148, u0_u13_u1_n149, u0_u13_u1_n150, u0_u13_u1_n151, u0_u13_u1_n152, u0_u13_u1_n153, u0_u13_u1_n154, u0_u13_u1_n155, 
       u0_u13_u1_n156, u0_u13_u1_n157, u0_u13_u1_n158, u0_u13_u1_n159, u0_u13_u1_n160, u0_u13_u1_n161, u0_u13_u1_n162, u0_u13_u1_n163, u0_u13_u1_n164, 
       u0_u13_u1_n165, u0_u13_u1_n166, u0_u13_u1_n167, u0_u13_u1_n168, u0_u13_u1_n169, u0_u13_u1_n170, u0_u13_u1_n171, u0_u13_u1_n172, u0_u13_u1_n173, 
       u0_u13_u1_n174, u0_u13_u1_n175, u0_u13_u1_n176, u0_u13_u1_n177, u0_u13_u1_n178, u0_u13_u1_n179, u0_u13_u1_n180, u0_u13_u1_n181, u0_u13_u1_n182, 
       u0_u13_u1_n183, u0_u13_u1_n184, u0_u13_u1_n185, u0_u13_u1_n186, u0_u13_u1_n187, u0_u13_u1_n188, u0_u13_u1_n95, u0_u13_u1_n96, u0_u13_u1_n97, 
       u0_u13_u1_n98, u0_u13_u1_n99, u0_u13_u2_n100, u0_u13_u2_n101, u0_u13_u2_n102, u0_u13_u2_n103, u0_u13_u2_n104, u0_u13_u2_n105, u0_u13_u2_n106, 
       u0_u13_u2_n107, u0_u13_u2_n108, u0_u13_u2_n109, u0_u13_u2_n110, u0_u13_u2_n111, u0_u13_u2_n112, u0_u13_u2_n113, u0_u13_u2_n114, u0_u13_u2_n115, 
       u0_u13_u2_n116, u0_u13_u2_n117, u0_u13_u2_n118, u0_u13_u2_n119, u0_u13_u2_n120, u0_u13_u2_n121, u0_u13_u2_n122, u0_u13_u2_n123, u0_u13_u2_n124, 
       u0_u13_u2_n125, u0_u13_u2_n126, u0_u13_u2_n127, u0_u13_u2_n128, u0_u13_u2_n129, u0_u13_u2_n130, u0_u13_u2_n131, u0_u13_u2_n132, u0_u13_u2_n133, 
       u0_u13_u2_n134, u0_u13_u2_n135, u0_u13_u2_n136, u0_u13_u2_n137, u0_u13_u2_n138, u0_u13_u2_n139, u0_u13_u2_n140, u0_u13_u2_n141, u0_u13_u2_n142, 
       u0_u13_u2_n143, u0_u13_u2_n144, u0_u13_u2_n145, u0_u13_u2_n146, u0_u13_u2_n147, u0_u13_u2_n148, u0_u13_u2_n149, u0_u13_u2_n150, u0_u13_u2_n151, 
       u0_u13_u2_n152, u0_u13_u2_n153, u0_u13_u2_n154, u0_u13_u2_n155, u0_u13_u2_n156, u0_u13_u2_n157, u0_u13_u2_n158, u0_u13_u2_n159, u0_u13_u2_n160, 
       u0_u13_u2_n161, u0_u13_u2_n162, u0_u13_u2_n163, u0_u13_u2_n164, u0_u13_u2_n165, u0_u13_u2_n166, u0_u13_u2_n167, u0_u13_u2_n168, u0_u13_u2_n169, 
       u0_u13_u2_n170, u0_u13_u2_n171, u0_u13_u2_n172, u0_u13_u2_n173, u0_u13_u2_n174, u0_u13_u2_n175, u0_u13_u2_n176, u0_u13_u2_n177, u0_u13_u2_n178, 
       u0_u13_u2_n179, u0_u13_u2_n180, u0_u13_u2_n181, u0_u13_u2_n182, u0_u13_u2_n183, u0_u13_u2_n184, u0_u13_u2_n185, u0_u13_u2_n186, u0_u13_u2_n187, 
       u0_u13_u2_n188, u0_u13_u2_n95, u0_u13_u2_n96, u0_u13_u2_n97, u0_u13_u2_n98, u0_u13_u2_n99, u0_u13_u3_n100, u0_u13_u3_n101, u0_u13_u3_n102, 
       u0_u13_u3_n103, u0_u13_u3_n104, u0_u13_u3_n105, u0_u13_u3_n106, u0_u13_u3_n107, u0_u13_u3_n108, u0_u13_u3_n109, u0_u13_u3_n110, u0_u13_u3_n111, 
       u0_u13_u3_n112, u0_u13_u3_n113, u0_u13_u3_n114, u0_u13_u3_n115, u0_u13_u3_n116, u0_u13_u3_n117, u0_u13_u3_n118, u0_u13_u3_n119, u0_u13_u3_n120, 
       u0_u13_u3_n121, u0_u13_u3_n122, u0_u13_u3_n123, u0_u13_u3_n124, u0_u13_u3_n125, u0_u13_u3_n126, u0_u13_u3_n127, u0_u13_u3_n128, u0_u13_u3_n129, 
       u0_u13_u3_n130, u0_u13_u3_n131, u0_u13_u3_n132, u0_u13_u3_n133, u0_u13_u3_n134, u0_u13_u3_n135, u0_u13_u3_n136, u0_u13_u3_n137, u0_u13_u3_n138, 
       u0_u13_u3_n139, u0_u13_u3_n140, u0_u13_u3_n141, u0_u13_u3_n142, u0_u13_u3_n143, u0_u13_u3_n144, u0_u13_u3_n145, u0_u13_u3_n146, u0_u13_u3_n147, 
       u0_u13_u3_n148, u0_u13_u3_n149, u0_u13_u3_n150, u0_u13_u3_n151, u0_u13_u3_n152, u0_u13_u3_n153, u0_u13_u3_n154, u0_u13_u3_n155, u0_u13_u3_n156, 
       u0_u13_u3_n157, u0_u13_u3_n158, u0_u13_u3_n159, u0_u13_u3_n160, u0_u13_u3_n161, u0_u13_u3_n162, u0_u13_u3_n163, u0_u13_u3_n164, u0_u13_u3_n165, 
       u0_u13_u3_n166, u0_u13_u3_n167, u0_u13_u3_n168, u0_u13_u3_n169, u0_u13_u3_n170, u0_u13_u3_n171, u0_u13_u3_n172, u0_u13_u3_n173, u0_u13_u3_n174, 
       u0_u13_u3_n175, u0_u13_u3_n176, u0_u13_u3_n177, u0_u13_u3_n178, u0_u13_u3_n179, u0_u13_u3_n180, u0_u13_u3_n181, u0_u13_u3_n182, u0_u13_u3_n183, 
       u0_u13_u3_n184, u0_u13_u3_n185, u0_u13_u3_n186, u0_u13_u3_n94, u0_u13_u3_n95, u0_u13_u3_n96, u0_u13_u3_n97, u0_u13_u3_n98, u0_u13_u3_n99, 
       u0_u13_u4_n100, u0_u13_u4_n101, u0_u13_u4_n102, u0_u13_u4_n103, u0_u13_u4_n104, u0_u13_u4_n105, u0_u13_u4_n106, u0_u13_u4_n107, u0_u13_u4_n108, 
       u0_u13_u4_n109, u0_u13_u4_n110, u0_u13_u4_n111, u0_u13_u4_n112, u0_u13_u4_n113, u0_u13_u4_n114, u0_u13_u4_n115, u0_u13_u4_n116, u0_u13_u4_n117, 
       u0_u13_u4_n118, u0_u13_u4_n119, u0_u13_u4_n120, u0_u13_u4_n121, u0_u13_u4_n122, u0_u13_u4_n123, u0_u13_u4_n124, u0_u13_u4_n125, u0_u13_u4_n126, 
       u0_u13_u4_n127, u0_u13_u4_n128, u0_u13_u4_n129, u0_u13_u4_n130, u0_u13_u4_n131, u0_u13_u4_n132, u0_u13_u4_n133, u0_u13_u4_n134, u0_u13_u4_n135, 
       u0_u13_u4_n136, u0_u13_u4_n137, u0_u13_u4_n138, u0_u13_u4_n139, u0_u13_u4_n140, u0_u13_u4_n141, u0_u13_u4_n142, u0_u13_u4_n143, u0_u13_u4_n144, 
       u0_u13_u4_n145, u0_u13_u4_n146, u0_u13_u4_n147, u0_u13_u4_n148, u0_u13_u4_n149, u0_u13_u4_n150, u0_u13_u4_n151, u0_u13_u4_n152, u0_u13_u4_n153, 
       u0_u13_u4_n154, u0_u13_u4_n155, u0_u13_u4_n156, u0_u13_u4_n157, u0_u13_u4_n158, u0_u13_u4_n159, u0_u13_u4_n160, u0_u13_u4_n161, u0_u13_u4_n162, 
       u0_u13_u4_n163, u0_u13_u4_n164, u0_u13_u4_n165, u0_u13_u4_n166, u0_u13_u4_n167, u0_u13_u4_n168, u0_u13_u4_n169, u0_u13_u4_n170, u0_u13_u4_n171, 
       u0_u13_u4_n172, u0_u13_u4_n173, u0_u13_u4_n174, u0_u13_u4_n175, u0_u13_u4_n176, u0_u13_u4_n177, u0_u13_u4_n178, u0_u13_u4_n179, u0_u13_u4_n180, 
       u0_u13_u4_n181, u0_u13_u4_n182, u0_u13_u4_n183, u0_u13_u4_n184, u0_u13_u4_n185, u0_u13_u4_n186, u0_u13_u4_n94, u0_u13_u4_n95, u0_u13_u4_n96, 
       u0_u13_u4_n97, u0_u13_u4_n98, u0_u13_u4_n99, u0_u9_X_25, u0_u9_X_26, u0_u9_X_27, u0_u9_X_28, u0_u9_X_29, u0_u9_X_30, 
       u0_u9_X_31, u0_u9_X_32, u0_u9_X_33, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_43, u0_u9_X_44, u0_u9_X_45, 
       u0_u9_X_46, u0_u9_X_47, u0_u9_X_48, u0_u9_u4_n100, u0_u9_u4_n101, u0_u9_u4_n102, u0_u9_u4_n103, u0_u9_u4_n104, u0_u9_u4_n105, 
       u0_u9_u4_n106, u0_u9_u4_n107, u0_u9_u4_n108, u0_u9_u4_n109, u0_u9_u4_n110, u0_u9_u4_n111, u0_u9_u4_n112, u0_u9_u4_n113, u0_u9_u4_n114, 
       u0_u9_u4_n115, u0_u9_u4_n116, u0_u9_u4_n117, u0_u9_u4_n118, u0_u9_u4_n119, u0_u9_u4_n120, u0_u9_u4_n121, u0_u9_u4_n122, u0_u9_u4_n123, 
       u0_u9_u4_n124, u0_u9_u4_n125, u0_u9_u4_n126, u0_u9_u4_n127, u0_u9_u4_n128, u0_u9_u4_n129, u0_u9_u4_n130, u0_u9_u4_n131, u0_u9_u4_n132, 
       u0_u9_u4_n133, u0_u9_u4_n134, u0_u9_u4_n135, u0_u9_u4_n136, u0_u9_u4_n137, u0_u9_u4_n138, u0_u9_u4_n139, u0_u9_u4_n140, u0_u9_u4_n141, 
       u0_u9_u4_n142, u0_u9_u4_n143, u0_u9_u4_n144, u0_u9_u4_n145, u0_u9_u4_n146, u0_u9_u4_n147, u0_u9_u4_n148, u0_u9_u4_n149, u0_u9_u4_n150, 
       u0_u9_u4_n151, u0_u9_u4_n152, u0_u9_u4_n153, u0_u9_u4_n154, u0_u9_u4_n155, u0_u9_u4_n156, u0_u9_u4_n157, u0_u9_u4_n158, u0_u9_u4_n159, 
       u0_u9_u4_n160, u0_u9_u4_n161, u0_u9_u4_n162, u0_u9_u4_n163, u0_u9_u4_n164, u0_u9_u4_n165, u0_u9_u4_n166, u0_u9_u4_n167, u0_u9_u4_n168, 
       u0_u9_u4_n169, u0_u9_u4_n170, u0_u9_u4_n171, u0_u9_u4_n172, u0_u9_u4_n173, u0_u9_u4_n174, u0_u9_u4_n175, u0_u9_u4_n176, u0_u9_u4_n177, 
       u0_u9_u4_n178, u0_u9_u4_n179, u0_u9_u4_n180, u0_u9_u4_n181, u0_u9_u4_n182, u0_u9_u4_n183, u0_u9_u4_n184, u0_u9_u4_n185, u0_u9_u4_n186, 
       u0_u9_u4_n94, u0_u9_u4_n95, u0_u9_u4_n96, u0_u9_u4_n97, u0_u9_u4_n98, u0_u9_u4_n99, u0_u9_u5_n100, u0_u9_u5_n101, u0_u9_u5_n102, 
       u0_u9_u5_n103, u0_u9_u5_n104, u0_u9_u5_n105, u0_u9_u5_n106, u0_u9_u5_n107, u0_u9_u5_n108, u0_u9_u5_n109, u0_u9_u5_n110, u0_u9_u5_n111, 
       u0_u9_u5_n112, u0_u9_u5_n113, u0_u9_u5_n114, u0_u9_u5_n115, u0_u9_u5_n116, u0_u9_u5_n117, u0_u9_u5_n118, u0_u9_u5_n119, u0_u9_u5_n120, 
       u0_u9_u5_n121, u0_u9_u5_n122, u0_u9_u5_n123, u0_u9_u5_n124, u0_u9_u5_n125, u0_u9_u5_n126, u0_u9_u5_n127, u0_u9_u5_n128, u0_u9_u5_n129, 
       u0_u9_u5_n130, u0_u9_u5_n131, u0_u9_u5_n132, u0_u9_u5_n133, u0_u9_u5_n134, u0_u9_u5_n135, u0_u9_u5_n136, u0_u9_u5_n137, u0_u9_u5_n138, 
       u0_u9_u5_n139, u0_u9_u5_n140, u0_u9_u5_n141, u0_u9_u5_n142, u0_u9_u5_n143, u0_u9_u5_n144, u0_u9_u5_n145, u0_u9_u5_n146, u0_u9_u5_n147, 
       u0_u9_u5_n148, u0_u9_u5_n149, u0_u9_u5_n150, u0_u9_u5_n151, u0_u9_u5_n152, u0_u9_u5_n153, u0_u9_u5_n154, u0_u9_u5_n155, u0_u9_u5_n156, 
       u0_u9_u5_n157, u0_u9_u5_n158, u0_u9_u5_n159, u0_u9_u5_n160, u0_u9_u5_n161, u0_u9_u5_n162, u0_u9_u5_n163, u0_u9_u5_n164, u0_u9_u5_n165, 
       u0_u9_u5_n166, u0_u9_u5_n167, u0_u9_u5_n168, u0_u9_u5_n169, u0_u9_u5_n170, u0_u9_u5_n171, u0_u9_u5_n172, u0_u9_u5_n173, u0_u9_u5_n174, 
       u0_u9_u5_n175, u0_u9_u5_n176, u0_u9_u5_n177, u0_u9_u5_n178, u0_u9_u5_n179, u0_u9_u5_n180, u0_u9_u5_n181, u0_u9_u5_n182, u0_u9_u5_n183, 
       u0_u9_u5_n184, u0_u9_u5_n185, u0_u9_u5_n186, u0_u9_u5_n187, u0_u9_u5_n188, u0_u9_u5_n189, u0_u9_u5_n190, u0_u9_u5_n191, u0_u9_u5_n192, 
       u0_u9_u5_n193, u0_u9_u5_n194, u0_u9_u5_n195, u0_u9_u5_n196, u0_u9_u5_n99, u0_u9_u7_n100, u0_u9_u7_n101, u0_u9_u7_n102, u0_u9_u7_n103, 
       u0_u9_u7_n104, u0_u9_u7_n105, u0_u9_u7_n106, u0_u9_u7_n107, u0_u9_u7_n108, u0_u9_u7_n109, u0_u9_u7_n110, u0_u9_u7_n111, u0_u9_u7_n112, 
       u0_u9_u7_n113, u0_u9_u7_n114, u0_u9_u7_n115, u0_u9_u7_n116, u0_u9_u7_n117, u0_u9_u7_n118, u0_u9_u7_n119, u0_u9_u7_n120, u0_u9_u7_n121, 
       u0_u9_u7_n122, u0_u9_u7_n123, u0_u9_u7_n124, u0_u9_u7_n125, u0_u9_u7_n126, u0_u9_u7_n127, u0_u9_u7_n128, u0_u9_u7_n129, u0_u9_u7_n130, 
       u0_u9_u7_n131, u0_u9_u7_n132, u0_u9_u7_n133, u0_u9_u7_n134, u0_u9_u7_n135, u0_u9_u7_n136, u0_u9_u7_n137, u0_u9_u7_n138, u0_u9_u7_n139, 
       u0_u9_u7_n140, u0_u9_u7_n141, u0_u9_u7_n142, u0_u9_u7_n143, u0_u9_u7_n144, u0_u9_u7_n145, u0_u9_u7_n146, u0_u9_u7_n147, u0_u9_u7_n148, 
       u0_u9_u7_n149, u0_u9_u7_n150, u0_u9_u7_n151, u0_u9_u7_n152, u0_u9_u7_n153, u0_u9_u7_n154, u0_u9_u7_n155, u0_u9_u7_n156, u0_u9_u7_n157, 
       u0_u9_u7_n158, u0_u9_u7_n159, u0_u9_u7_n160, u0_u9_u7_n161, u0_u9_u7_n162, u0_u9_u7_n163, u0_u9_u7_n164, u0_u9_u7_n165, u0_u9_u7_n166, 
       u0_u9_u7_n167, u0_u9_u7_n168, u0_u9_u7_n169, u0_u9_u7_n170, u0_u9_u7_n171, u0_u9_u7_n172, u0_u9_u7_n173, u0_u9_u7_n174, u0_u9_u7_n175, 
       u0_u9_u7_n176, u0_u9_u7_n177, u0_u9_u7_n178, u0_u9_u7_n179, u0_u9_u7_n180, u0_u9_u7_n91, u0_u9_u7_n92, u0_u9_u7_n93, u0_u9_u7_n94, 
       u0_u9_u7_n95, u0_u9_u7_n96, u0_u9_u7_n97, u0_u9_u7_n98, u0_u9_u7_n99, u0_uk_n1011, u0_uk_n1014, u0_uk_n935, u0_uk_n938, 
       u1_K10_43, u1_K10_44, u1_K10_45, u1_K10_46, u1_K10_47, u1_K10_48, u1_K15_31, u1_K15_32, u1_K15_33, 
       u1_K15_34, u1_K15_35, u1_K15_36, u1_K15_37, u1_K15_38, u1_K15_39, u1_K15_40, u1_K15_41, u1_K15_42, 
       u1_K15_43, u1_K15_44, u1_K15_45, u1_K15_46, u1_K15_47, u1_K15_48, u1_K1_25, u1_K1_26, u1_K1_27, 
       u1_K1_28, u1_K1_29, u1_K1_30, u1_K1_31, u1_K1_32, u1_K1_33, u1_K1_34, u1_K1_35, u1_K1_36, 
       u1_K1_37, u1_K1_38, u1_K1_39, u1_K1_40, u1_K1_41, u1_K1_42, u1_K1_43, u1_K1_44, u1_K1_45, 
       u1_K1_46, u1_K1_47, u1_K1_48, u1_K4_10, u1_K4_11, u1_K4_12, u1_K4_7, u1_K4_8, u1_K4_9, 
       u1_K5_31, u1_K5_32, u1_K5_33, u1_K5_34, u1_K5_35, u1_K5_36, u1_K6_1, u1_K6_13, u1_K6_14, 
       u1_K6_15, u1_K6_16, u1_K6_17, u1_K6_18, u1_K6_19, u1_K6_2, u1_K6_20, u1_K6_21, u1_K6_22, 
       u1_K6_23, u1_K6_24, u1_K6_25, u1_K6_26, u1_K6_27, u1_K6_28, u1_K6_29, u1_K6_3, u1_K6_30, 
       u1_K6_31, u1_K6_32, u1_K6_33, u1_K6_34, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, u1_K6_39, 
       u1_K6_4, u1_K6_40, u1_K6_41, u1_K6_42, u1_K6_5, u1_K6_6, u1_K9_1, u1_K9_10, u1_K9_11, 
       u1_K9_12, u1_K9_13, u1_K9_14, u1_K9_15, u1_K9_16, u1_K9_17, u1_K9_18, u1_K9_19, u1_K9_2, 
       u1_K9_20, u1_K9_21, u1_K9_22, u1_K9_23, u1_K9_24, u1_K9_3, u1_K9_4, u1_K9_5, u1_K9_6, 
       u1_K9_7, u1_K9_8, u1_K9_9, u1_out0_11, u1_out0_12, u1_out0_14, u1_out0_15, u1_out0_19, u1_out0_21, 
       u1_out0_22, u1_out0_25, u1_out0_27, u1_out0_29, u1_out0_3, u1_out0_32, u1_out0_4, u1_out0_5, u1_out0_7, 
       u1_out0_8, u1_out14_11, u1_out14_12, u1_out14_15, u1_out14_19, u1_out14_21, u1_out14_22, u1_out14_27, u1_out14_29, 
       u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_7, u1_out3_13, u1_out3_18, u1_out3_2, u1_out3_28, u1_out4_11, 
       u1_out4_19, u1_out4_29, u1_out4_4, u1_out5_1, u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_14, u1_out5_16, 
       u1_out5_17, u1_out5_19, u1_out5_20, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_25, u1_out5_26, u1_out5_29, 
       u1_out5_3, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_6, u1_out5_7, u1_out5_8, u1_out5_9, 
       u1_out8_1, u1_out8_10, u1_out8_13, u1_out8_16, u1_out8_17, u1_out8_18, u1_out8_2, u1_out8_20, u1_out8_23, 
       u1_out8_24, u1_out8_26, u1_out8_28, u1_out8_30, u1_out8_31, u1_out8_6, u1_out8_9, u1_out9_15, u1_out9_21, 
       u1_out9_27, u1_out9_5, u1_u0_X_25, u1_u0_X_26, u1_u0_X_27, u1_u0_X_28, u1_u0_X_29, u1_u0_X_30, u1_u0_X_31, 
       u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_39, u1_u0_X_40, 
       u1_u0_X_41, u1_u0_X_42, u1_u0_X_43, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, u1_u0_X_47, u1_u0_X_48, u1_u0_u4_n100, 
       u1_u0_u4_n101, u1_u0_u4_n102, u1_u0_u4_n103, u1_u0_u4_n104, u1_u0_u4_n105, u1_u0_u4_n106, u1_u0_u4_n107, u1_u0_u4_n108, u1_u0_u4_n109, 
       u1_u0_u4_n110, u1_u0_u4_n111, u1_u0_u4_n112, u1_u0_u4_n113, u1_u0_u4_n114, u1_u0_u4_n115, u1_u0_u4_n116, u1_u0_u4_n117, u1_u0_u4_n118, 
       u1_u0_u4_n119, u1_u0_u4_n120, u1_u0_u4_n121, u1_u0_u4_n122, u1_u0_u4_n123, u1_u0_u4_n124, u1_u0_u4_n125, u1_u0_u4_n126, u1_u0_u4_n127, 
       u1_u0_u4_n128, u1_u0_u4_n129, u1_u0_u4_n130, u1_u0_u4_n131, u1_u0_u4_n132, u1_u0_u4_n133, u1_u0_u4_n134, u1_u0_u4_n135, u1_u0_u4_n136, 
       u1_u0_u4_n137, u1_u0_u4_n138, u1_u0_u4_n139, u1_u0_u4_n140, u1_u0_u4_n141, u1_u0_u4_n142, u1_u0_u4_n143, u1_u0_u4_n144, u1_u0_u4_n145, 
       u1_u0_u4_n146, u1_u0_u4_n147, u1_u0_u4_n148, u1_u0_u4_n149, u1_u0_u4_n150, u1_u0_u4_n151, u1_u0_u4_n152, u1_u0_u4_n153, u1_u0_u4_n154, 
       u1_u0_u4_n155, u1_u0_u4_n156, u1_u0_u4_n157, u1_u0_u4_n158, u1_u0_u4_n159, u1_u0_u4_n160, u1_u0_u4_n161, u1_u0_u4_n162, u1_u0_u4_n163, 
       u1_u0_u4_n164, u1_u0_u4_n165, u1_u0_u4_n166, u1_u0_u4_n167, u1_u0_u4_n168, u1_u0_u4_n169, u1_u0_u4_n170, u1_u0_u4_n171, u1_u0_u4_n172, 
       u1_u0_u4_n173, u1_u0_u4_n174, u1_u0_u4_n175, u1_u0_u4_n176, u1_u0_u4_n177, u1_u0_u4_n178, u1_u0_u4_n179, u1_u0_u4_n180, u1_u0_u4_n181, 
       u1_u0_u4_n182, u1_u0_u4_n183, u1_u0_u4_n184, u1_u0_u4_n185, u1_u0_u4_n186, u1_u0_u4_n94, u1_u0_u4_n95, u1_u0_u4_n96, u1_u0_u4_n97, 
       u1_u0_u4_n98, u1_u0_u4_n99, u1_u0_u5_n100, u1_u0_u5_n101, u1_u0_u5_n102, u1_u0_u5_n103, u1_u0_u5_n104, u1_u0_u5_n105, u1_u0_u5_n106, 
       u1_u0_u5_n107, u1_u0_u5_n108, u1_u0_u5_n109, u1_u0_u5_n110, u1_u0_u5_n111, u1_u0_u5_n112, u1_u0_u5_n113, u1_u0_u5_n114, u1_u0_u5_n115, 
       u1_u0_u5_n116, u1_u0_u5_n117, u1_u0_u5_n118, u1_u0_u5_n119, u1_u0_u5_n120, u1_u0_u5_n121, u1_u0_u5_n122, u1_u0_u5_n123, u1_u0_u5_n124, 
       u1_u0_u5_n125, u1_u0_u5_n126, u1_u0_u5_n127, u1_u0_u5_n128, u1_u0_u5_n129, u1_u0_u5_n130, u1_u0_u5_n131, u1_u0_u5_n132, u1_u0_u5_n133, 
       u1_u0_u5_n134, u1_u0_u5_n135, u1_u0_u5_n136, u1_u0_u5_n137, u1_u0_u5_n138, u1_u0_u5_n139, u1_u0_u5_n140, u1_u0_u5_n141, u1_u0_u5_n142, 
       u1_u0_u5_n143, u1_u0_u5_n144, u1_u0_u5_n145, u1_u0_u5_n146, u1_u0_u5_n147, u1_u0_u5_n148, u1_u0_u5_n149, u1_u0_u5_n150, u1_u0_u5_n151, 
       u1_u0_u5_n152, u1_u0_u5_n153, u1_u0_u5_n154, u1_u0_u5_n155, u1_u0_u5_n156, u1_u0_u5_n157, u1_u0_u5_n158, u1_u0_u5_n159, u1_u0_u5_n160, 
       u1_u0_u5_n161, u1_u0_u5_n162, u1_u0_u5_n163, u1_u0_u5_n164, u1_u0_u5_n165, u1_u0_u5_n166, u1_u0_u5_n167, u1_u0_u5_n168, u1_u0_u5_n169, 
       u1_u0_u5_n170, u1_u0_u5_n171, u1_u0_u5_n172, u1_u0_u5_n173, u1_u0_u5_n174, u1_u0_u5_n175, u1_u0_u5_n176, u1_u0_u5_n177, u1_u0_u5_n178, 
       u1_u0_u5_n179, u1_u0_u5_n180, u1_u0_u5_n181, u1_u0_u5_n182, u1_u0_u5_n183, u1_u0_u5_n184, u1_u0_u5_n185, u1_u0_u5_n186, u1_u0_u5_n187, 
       u1_u0_u5_n188, u1_u0_u5_n189, u1_u0_u5_n190, u1_u0_u5_n191, u1_u0_u5_n192, u1_u0_u5_n193, u1_u0_u5_n194, u1_u0_u5_n195, u1_u0_u5_n196, 
       u1_u0_u5_n99, u1_u0_u6_n100, u1_u0_u6_n101, u1_u0_u6_n102, u1_u0_u6_n103, u1_u0_u6_n104, u1_u0_u6_n105, u1_u0_u6_n106, u1_u0_u6_n107, 
       u1_u0_u6_n108, u1_u0_u6_n109, u1_u0_u6_n110, u1_u0_u6_n111, u1_u0_u6_n112, u1_u0_u6_n113, u1_u0_u6_n114, u1_u0_u6_n115, u1_u0_u6_n116, 
       u1_u0_u6_n117, u1_u0_u6_n118, u1_u0_u6_n119, u1_u0_u6_n120, u1_u0_u6_n121, u1_u0_u6_n122, u1_u0_u6_n123, u1_u0_u6_n124, u1_u0_u6_n125, 
       u1_u0_u6_n126, u1_u0_u6_n127, u1_u0_u6_n128, u1_u0_u6_n129, u1_u0_u6_n130, u1_u0_u6_n131, u1_u0_u6_n132, u1_u0_u6_n133, u1_u0_u6_n134, 
       u1_u0_u6_n135, u1_u0_u6_n136, u1_u0_u6_n137, u1_u0_u6_n138, u1_u0_u6_n139, u1_u0_u6_n140, u1_u0_u6_n141, u1_u0_u6_n142, u1_u0_u6_n143, 
       u1_u0_u6_n144, u1_u0_u6_n145, u1_u0_u6_n146, u1_u0_u6_n147, u1_u0_u6_n148, u1_u0_u6_n149, u1_u0_u6_n150, u1_u0_u6_n151, u1_u0_u6_n152, 
       u1_u0_u6_n153, u1_u0_u6_n154, u1_u0_u6_n155, u1_u0_u6_n156, u1_u0_u6_n157, u1_u0_u6_n158, u1_u0_u6_n159, u1_u0_u6_n160, u1_u0_u6_n161, 
       u1_u0_u6_n162, u1_u0_u6_n163, u1_u0_u6_n164, u1_u0_u6_n165, u1_u0_u6_n166, u1_u0_u6_n167, u1_u0_u6_n168, u1_u0_u6_n169, u1_u0_u6_n170, 
       u1_u0_u6_n171, u1_u0_u6_n172, u1_u0_u6_n173, u1_u0_u6_n174, u1_u0_u6_n88, u1_u0_u6_n89, u1_u0_u6_n90, u1_u0_u6_n91, u1_u0_u6_n92, 
       u1_u0_u6_n93, u1_u0_u6_n94, u1_u0_u6_n95, u1_u0_u6_n96, u1_u0_u6_n97, u1_u0_u6_n98, u1_u0_u6_n99, u1_u0_u7_n100, u1_u0_u7_n101, 
       u1_u0_u7_n102, u1_u0_u7_n103, u1_u0_u7_n104, u1_u0_u7_n105, u1_u0_u7_n106, u1_u0_u7_n107, u1_u0_u7_n108, u1_u0_u7_n109, u1_u0_u7_n110, 
       u1_u0_u7_n111, u1_u0_u7_n112, u1_u0_u7_n113, u1_u0_u7_n114, u1_u0_u7_n115, u1_u0_u7_n116, u1_u0_u7_n117, u1_u0_u7_n118, u1_u0_u7_n119, 
       u1_u0_u7_n120, u1_u0_u7_n121, u1_u0_u7_n122, u1_u0_u7_n123, u1_u0_u7_n124, u1_u0_u7_n125, u1_u0_u7_n126, u1_u0_u7_n127, u1_u0_u7_n128, 
       u1_u0_u7_n129, u1_u0_u7_n130, u1_u0_u7_n131, u1_u0_u7_n132, u1_u0_u7_n133, u1_u0_u7_n134, u1_u0_u7_n135, u1_u0_u7_n136, u1_u0_u7_n137, 
       u1_u0_u7_n138, u1_u0_u7_n139, u1_u0_u7_n140, u1_u0_u7_n141, u1_u0_u7_n142, u1_u0_u7_n143, u1_u0_u7_n144, u1_u0_u7_n145, u1_u0_u7_n146, 
       u1_u0_u7_n147, u1_u0_u7_n148, u1_u0_u7_n149, u1_u0_u7_n150, u1_u0_u7_n151, u1_u0_u7_n152, u1_u0_u7_n153, u1_u0_u7_n154, u1_u0_u7_n155, 
       u1_u0_u7_n156, u1_u0_u7_n157, u1_u0_u7_n158, u1_u0_u7_n159, u1_u0_u7_n160, u1_u0_u7_n161, u1_u0_u7_n162, u1_u0_u7_n163, u1_u0_u7_n164, 
       u1_u0_u7_n165, u1_u0_u7_n166, u1_u0_u7_n167, u1_u0_u7_n168, u1_u0_u7_n169, u1_u0_u7_n170, u1_u0_u7_n171, u1_u0_u7_n172, u1_u0_u7_n173, 
       u1_u0_u7_n174, u1_u0_u7_n175, u1_u0_u7_n176, u1_u0_u7_n177, u1_u0_u7_n178, u1_u0_u7_n179, u1_u0_u7_n180, u1_u0_u7_n91, u1_u0_u7_n92, 
       u1_u0_u7_n93, u1_u0_u7_n94, u1_u0_u7_n95, u1_u0_u7_n96, u1_u0_u7_n97, u1_u0_u7_n98, u1_u0_u7_n99, u1_u14_X_31, u1_u14_X_32, 
       u1_u14_X_33, u1_u14_X_34, u1_u14_X_35, u1_u14_X_36, u1_u14_X_37, u1_u14_X_38, u1_u14_X_39, u1_u14_X_40, u1_u14_X_41, 
       u1_u14_X_42, u1_u14_X_43, u1_u14_X_44, u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, u1_u14_X_48, u1_u14_u5_n100, u1_u14_u5_n101, 
       u1_u14_u5_n102, u1_u14_u5_n103, u1_u14_u5_n104, u1_u14_u5_n105, u1_u14_u5_n106, u1_u14_u5_n107, u1_u14_u5_n108, u1_u14_u5_n109, u1_u14_u5_n110, 
       u1_u14_u5_n111, u1_u14_u5_n112, u1_u14_u5_n113, u1_u14_u5_n114, u1_u14_u5_n115, u1_u14_u5_n116, u1_u14_u5_n117, u1_u14_u5_n118, u1_u14_u5_n119, 
       u1_u14_u5_n120, u1_u14_u5_n121, u1_u14_u5_n122, u1_u14_u5_n123, u1_u14_u5_n124, u1_u14_u5_n125, u1_u14_u5_n126, u1_u14_u5_n127, u1_u14_u5_n128, 
       u1_u14_u5_n129, u1_u14_u5_n130, u1_u14_u5_n131, u1_u14_u5_n132, u1_u14_u5_n133, u1_u14_u5_n134, u1_u14_u5_n135, u1_u14_u5_n136, u1_u14_u5_n137, 
       u1_u14_u5_n138, u1_u14_u5_n139, u1_u14_u5_n140, u1_u14_u5_n141, u1_u14_u5_n142, u1_u14_u5_n143, u1_u14_u5_n144, u1_u14_u5_n145, u1_u14_u5_n146, 
       u1_u14_u5_n147, u1_u14_u5_n148, u1_u14_u5_n149, u1_u14_u5_n150, u1_u14_u5_n151, u1_u14_u5_n152, u1_u14_u5_n153, u1_u14_u5_n154, u1_u14_u5_n155, 
       u1_u14_u5_n156, u1_u14_u5_n157, u1_u14_u5_n158, u1_u14_u5_n159, u1_u14_u5_n160, u1_u14_u5_n161, u1_u14_u5_n162, u1_u14_u5_n163, u1_u14_u5_n164, 
       u1_u14_u5_n165, u1_u14_u5_n166, u1_u14_u5_n167, u1_u14_u5_n168, u1_u14_u5_n169, u1_u14_u5_n170, u1_u14_u5_n171, u1_u14_u5_n172, u1_u14_u5_n173, 
       u1_u14_u5_n174, u1_u14_u5_n175, u1_u14_u5_n176, u1_u14_u5_n177, u1_u14_u5_n178, u1_u14_u5_n179, u1_u14_u5_n180, u1_u14_u5_n181, u1_u14_u5_n182, 
       u1_u14_u5_n183, u1_u14_u5_n184, u1_u14_u5_n185, u1_u14_u5_n186, u1_u14_u5_n187, u1_u14_u5_n188, u1_u14_u5_n189, u1_u14_u5_n190, u1_u14_u5_n191, 
       u1_u14_u5_n192, u1_u14_u5_n193, u1_u14_u5_n194, u1_u14_u5_n195, u1_u14_u5_n196, u1_u14_u5_n99, u1_u14_u6_n100, u1_u14_u6_n101, u1_u14_u6_n102, 
       u1_u14_u6_n103, u1_u14_u6_n104, u1_u14_u6_n105, u1_u14_u6_n106, u1_u14_u6_n107, u1_u14_u6_n108, u1_u14_u6_n109, u1_u14_u6_n110, u1_u14_u6_n111, 
       u1_u14_u6_n112, u1_u14_u6_n113, u1_u14_u6_n114, u1_u14_u6_n115, u1_u14_u6_n116, u1_u14_u6_n117, u1_u14_u6_n118, u1_u14_u6_n119, u1_u14_u6_n120, 
       u1_u14_u6_n121, u1_u14_u6_n122, u1_u14_u6_n123, u1_u14_u6_n124, u1_u14_u6_n125, u1_u14_u6_n126, u1_u14_u6_n127, u1_u14_u6_n128, u1_u14_u6_n129, 
       u1_u14_u6_n130, u1_u14_u6_n131, u1_u14_u6_n132, u1_u14_u6_n133, u1_u14_u6_n134, u1_u14_u6_n135, u1_u14_u6_n136, u1_u14_u6_n137, u1_u14_u6_n138, 
       u1_u14_u6_n139, u1_u14_u6_n140, u1_u14_u6_n141, u1_u14_u6_n142, u1_u14_u6_n143, u1_u14_u6_n144, u1_u14_u6_n145, u1_u14_u6_n146, u1_u14_u6_n147, 
       u1_u14_u6_n148, u1_u14_u6_n149, u1_u14_u6_n150, u1_u14_u6_n151, u1_u14_u6_n152, u1_u14_u6_n153, u1_u14_u6_n154, u1_u14_u6_n155, u1_u14_u6_n156, 
       u1_u14_u6_n157, u1_u14_u6_n158, u1_u14_u6_n159, u1_u14_u6_n160, u1_u14_u6_n161, u1_u14_u6_n162, u1_u14_u6_n163, u1_u14_u6_n164, u1_u14_u6_n165, 
       u1_u14_u6_n166, u1_u14_u6_n167, u1_u14_u6_n168, u1_u14_u6_n169, u1_u14_u6_n170, u1_u14_u6_n171, u1_u14_u6_n172, u1_u14_u6_n173, u1_u14_u6_n174, 
       u1_u14_u6_n88, u1_u14_u6_n89, u1_u14_u6_n90, u1_u14_u6_n91, u1_u14_u6_n92, u1_u14_u6_n93, u1_u14_u6_n94, u1_u14_u6_n95, u1_u14_u6_n96, 
       u1_u14_u6_n97, u1_u14_u6_n98, u1_u14_u6_n99, u1_u14_u7_n100, u1_u14_u7_n101, u1_u14_u7_n102, u1_u14_u7_n103, u1_u14_u7_n104, u1_u14_u7_n105, 
       u1_u14_u7_n106, u1_u14_u7_n107, u1_u14_u7_n108, u1_u14_u7_n109, u1_u14_u7_n110, u1_u14_u7_n111, u1_u14_u7_n112, u1_u14_u7_n113, u1_u14_u7_n114, 
       u1_u14_u7_n115, u1_u14_u7_n116, u1_u14_u7_n117, u1_u14_u7_n118, u1_u14_u7_n119, u1_u14_u7_n120, u1_u14_u7_n121, u1_u14_u7_n122, u1_u14_u7_n123, 
       u1_u14_u7_n124, u1_u14_u7_n125, u1_u14_u7_n126, u1_u14_u7_n127, u1_u14_u7_n128, u1_u14_u7_n129, u1_u14_u7_n130, u1_u14_u7_n131, u1_u14_u7_n132, 
       u1_u14_u7_n133, u1_u14_u7_n134, u1_u14_u7_n135, u1_u14_u7_n136, u1_u14_u7_n137, u1_u14_u7_n138, u1_u14_u7_n139, u1_u14_u7_n140, u1_u14_u7_n141, 
       u1_u14_u7_n142, u1_u14_u7_n143, u1_u14_u7_n144, u1_u14_u7_n145, u1_u14_u7_n146, u1_u14_u7_n147, u1_u14_u7_n148, u1_u14_u7_n149, u1_u14_u7_n150, 
       u1_u14_u7_n151, u1_u14_u7_n152, u1_u14_u7_n153, u1_u14_u7_n154, u1_u14_u7_n155, u1_u14_u7_n156, u1_u14_u7_n157, u1_u14_u7_n158, u1_u14_u7_n159, 
       u1_u14_u7_n160, u1_u14_u7_n161, u1_u14_u7_n162, u1_u14_u7_n163, u1_u14_u7_n164, u1_u14_u7_n165, u1_u14_u7_n166, u1_u14_u7_n167, u1_u14_u7_n168, 
       u1_u14_u7_n169, u1_u14_u7_n170, u1_u14_u7_n171, u1_u14_u7_n172, u1_u14_u7_n173, u1_u14_u7_n174, u1_u14_u7_n175, u1_u14_u7_n176, u1_u14_u7_n177, 
       u1_u14_u7_n178, u1_u14_u7_n179, u1_u14_u7_n180, u1_u14_u7_n91, u1_u14_u7_n92, u1_u14_u7_n93, u1_u14_u7_n94, u1_u14_u7_n95, u1_u14_u7_n96, 
       u1_u14_u7_n97, u1_u14_u7_n98, u1_u14_u7_n99, u1_u3_X_10, u1_u3_X_11, u1_u3_X_12, u1_u3_X_7, u1_u3_X_8, u1_u3_X_9, 
       u1_u3_u1_n100, u1_u3_u1_n101, u1_u3_u1_n102, u1_u3_u1_n103, u1_u3_u1_n104, u1_u3_u1_n105, u1_u3_u1_n106, u1_u3_u1_n107, u1_u3_u1_n108, 
       u1_u3_u1_n109, u1_u3_u1_n110, u1_u3_u1_n111, u1_u3_u1_n112, u1_u3_u1_n113, u1_u3_u1_n114, u1_u3_u1_n115, u1_u3_u1_n116, u1_u3_u1_n117, 
       u1_u3_u1_n118, u1_u3_u1_n119, u1_u3_u1_n120, u1_u3_u1_n121, u1_u3_u1_n122, u1_u3_u1_n123, u1_u3_u1_n124, u1_u3_u1_n125, u1_u3_u1_n126, 
       u1_u3_u1_n127, u1_u3_u1_n128, u1_u3_u1_n129, u1_u3_u1_n130, u1_u3_u1_n131, u1_u3_u1_n132, u1_u3_u1_n133, u1_u3_u1_n134, u1_u3_u1_n135, 
       u1_u3_u1_n136, u1_u3_u1_n137, u1_u3_u1_n138, u1_u3_u1_n139, u1_u3_u1_n140, u1_u3_u1_n141, u1_u3_u1_n142, u1_u3_u1_n143, u1_u3_u1_n144, 
       u1_u3_u1_n145, u1_u3_u1_n146, u1_u3_u1_n147, u1_u3_u1_n148, u1_u3_u1_n149, u1_u3_u1_n150, u1_u3_u1_n151, u1_u3_u1_n152, u1_u3_u1_n153, 
       u1_u3_u1_n154, u1_u3_u1_n155, u1_u3_u1_n156, u1_u3_u1_n157, u1_u3_u1_n158, u1_u3_u1_n159, u1_u3_u1_n160, u1_u3_u1_n161, u1_u3_u1_n162, 
       u1_u3_u1_n163, u1_u3_u1_n164, u1_u3_u1_n165, u1_u3_u1_n166, u1_u3_u1_n167, u1_u3_u1_n168, u1_u3_u1_n169, u1_u3_u1_n170, u1_u3_u1_n171, 
       u1_u3_u1_n172, u1_u3_u1_n173, u1_u3_u1_n174, u1_u3_u1_n175, u1_u3_u1_n176, u1_u3_u1_n177, u1_u3_u1_n178, u1_u3_u1_n179, u1_u3_u1_n180, 
       u1_u3_u1_n181, u1_u3_u1_n182, u1_u3_u1_n183, u1_u3_u1_n184, u1_u3_u1_n185, u1_u3_u1_n186, u1_u3_u1_n187, u1_u3_u1_n188, u1_u3_u1_n95, 
       u1_u3_u1_n96, u1_u3_u1_n97, u1_u3_u1_n98, u1_u3_u1_n99, u1_u4_X_31, u1_u4_X_32, u1_u4_X_33, u1_u4_X_34, u1_u4_X_35, 
       u1_u4_X_36, u1_u4_u5_n100, u1_u4_u5_n101, u1_u4_u5_n102, u1_u4_u5_n103, u1_u4_u5_n104, u1_u4_u5_n105, u1_u4_u5_n106, u1_u4_u5_n107, 
       u1_u4_u5_n108, u1_u4_u5_n109, u1_u4_u5_n110, u1_u4_u5_n111, u1_u4_u5_n112, u1_u4_u5_n113, u1_u4_u5_n114, u1_u4_u5_n115, u1_u4_u5_n116, 
       u1_u4_u5_n117, u1_u4_u5_n118, u1_u4_u5_n119, u1_u4_u5_n120, u1_u4_u5_n121, u1_u4_u5_n122, u1_u4_u5_n123, u1_u4_u5_n124, u1_u4_u5_n125, 
       u1_u4_u5_n126, u1_u4_u5_n127, u1_u4_u5_n128, u1_u4_u5_n129, u1_u4_u5_n130, u1_u4_u5_n131, u1_u4_u5_n132, u1_u4_u5_n133, u1_u4_u5_n134, 
       u1_u4_u5_n135, u1_u4_u5_n136, u1_u4_u5_n137, u1_u4_u5_n138, u1_u4_u5_n139, u1_u4_u5_n140, u1_u4_u5_n141, u1_u4_u5_n142, u1_u4_u5_n143, 
       u1_u4_u5_n144, u1_u4_u5_n145, u1_u4_u5_n146, u1_u4_u5_n147, u1_u4_u5_n148, u1_u4_u5_n149, u1_u4_u5_n150, u1_u4_u5_n151, u1_u4_u5_n152, 
       u1_u4_u5_n153, u1_u4_u5_n154, u1_u4_u5_n155, u1_u4_u5_n156, u1_u4_u5_n157, u1_u4_u5_n158, u1_u4_u5_n159, u1_u4_u5_n160, u1_u4_u5_n161, 
       u1_u4_u5_n162, u1_u4_u5_n163, u1_u4_u5_n164, u1_u4_u5_n165, u1_u4_u5_n166, u1_u4_u5_n167, u1_u4_u5_n168, u1_u4_u5_n169, u1_u4_u5_n170, 
       u1_u4_u5_n171, u1_u4_u5_n172, u1_u4_u5_n173, u1_u4_u5_n174, u1_u4_u5_n175, u1_u4_u5_n176, u1_u4_u5_n177, u1_u4_u5_n178, u1_u4_u5_n179, 
       u1_u4_u5_n180, u1_u4_u5_n181, u1_u4_u5_n182, u1_u4_u5_n183, u1_u4_u5_n184, u1_u4_u5_n185, u1_u4_u5_n186, u1_u4_u5_n187, u1_u4_u5_n188, 
       u1_u4_u5_n189, u1_u4_u5_n190, u1_u4_u5_n191, u1_u4_u5_n192, u1_u4_u5_n193, u1_u4_u5_n194, u1_u4_u5_n195, u1_u4_u5_n196, u1_u4_u5_n99, 
       u1_u5_X_1, u1_u5_X_13, u1_u5_X_14, u1_u5_X_15, u1_u5_X_16, u1_u5_X_17, u1_u5_X_18, u1_u5_X_19, u1_u5_X_2, 
       u1_u5_X_20, u1_u5_X_21, u1_u5_X_22, u1_u5_X_23, u1_u5_X_24, u1_u5_X_25, u1_u5_X_26, u1_u5_X_27, u1_u5_X_28, 
       u1_u5_X_29, u1_u5_X_3, u1_u5_X_30, u1_u5_X_31, u1_u5_X_32, u1_u5_X_33, u1_u5_X_34, u1_u5_X_35, u1_u5_X_36, 
       u1_u5_X_37, u1_u5_X_38, u1_u5_X_39, u1_u5_X_4, u1_u5_X_40, u1_u5_X_41, u1_u5_X_42, u1_u5_X_5, u1_u5_X_6, 
       u1_u5_u0_n100, u1_u5_u0_n101, u1_u5_u0_n102, u1_u5_u0_n103, u1_u5_u0_n104, u1_u5_u0_n105, u1_u5_u0_n106, u1_u5_u0_n107, u1_u5_u0_n108, 
       u1_u5_u0_n109, u1_u5_u0_n110, u1_u5_u0_n111, u1_u5_u0_n112, u1_u5_u0_n113, u1_u5_u0_n114, u1_u5_u0_n115, u1_u5_u0_n116, u1_u5_u0_n117, 
       u1_u5_u0_n118, u1_u5_u0_n119, u1_u5_u0_n120, u1_u5_u0_n121, u1_u5_u0_n122, u1_u5_u0_n123, u1_u5_u0_n124, u1_u5_u0_n125, u1_u5_u0_n126, 
       u1_u5_u0_n127, u1_u5_u0_n128, u1_u5_u0_n129, u1_u5_u0_n130, u1_u5_u0_n131, u1_u5_u0_n132, u1_u5_u0_n133, u1_u5_u0_n134, u1_u5_u0_n135, 
       u1_u5_u0_n136, u1_u5_u0_n137, u1_u5_u0_n138, u1_u5_u0_n139, u1_u5_u0_n140, u1_u5_u0_n141, u1_u5_u0_n142, u1_u5_u0_n143, u1_u5_u0_n144, 
       u1_u5_u0_n145, u1_u5_u0_n146, u1_u5_u0_n147, u1_u5_u0_n148, u1_u5_u0_n149, u1_u5_u0_n150, u1_u5_u0_n151, u1_u5_u0_n152, u1_u5_u0_n153, 
       u1_u5_u0_n154, u1_u5_u0_n155, u1_u5_u0_n156, u1_u5_u0_n157, u1_u5_u0_n158, u1_u5_u0_n159, u1_u5_u0_n160, u1_u5_u0_n161, u1_u5_u0_n162, 
       u1_u5_u0_n163, u1_u5_u0_n164, u1_u5_u0_n165, u1_u5_u0_n166, u1_u5_u0_n167, u1_u5_u0_n168, u1_u5_u0_n169, u1_u5_u0_n170, u1_u5_u0_n171, 
       u1_u5_u0_n172, u1_u5_u0_n173, u1_u5_u0_n174, u1_u5_u0_n88, u1_u5_u0_n89, u1_u5_u0_n90, u1_u5_u0_n91, u1_u5_u0_n92, u1_u5_u0_n93, 
       u1_u5_u0_n94, u1_u5_u0_n95, u1_u5_u0_n96, u1_u5_u0_n97, u1_u5_u0_n98, u1_u5_u0_n99, u1_u5_u2_n100, u1_u5_u2_n101, u1_u5_u2_n102, 
       u1_u5_u2_n103, u1_u5_u2_n104, u1_u5_u2_n105, u1_u5_u2_n106, u1_u5_u2_n107, u1_u5_u2_n108, u1_u5_u2_n109, u1_u5_u2_n110, u1_u5_u2_n111, 
       u1_u5_u2_n112, u1_u5_u2_n113, u1_u5_u2_n114, u1_u5_u2_n115, u1_u5_u2_n116, u1_u5_u2_n117, u1_u5_u2_n118, u1_u5_u2_n119, u1_u5_u2_n120, 
       u1_u5_u2_n121, u1_u5_u2_n122, u1_u5_u2_n123, u1_u5_u2_n124, u1_u5_u2_n125, u1_u5_u2_n126, u1_u5_u2_n127, u1_u5_u2_n128, u1_u5_u2_n129, 
       u1_u5_u2_n130, u1_u5_u2_n131, u1_u5_u2_n132, u1_u5_u2_n133, u1_u5_u2_n134, u1_u5_u2_n135, u1_u5_u2_n136, u1_u5_u2_n137, u1_u5_u2_n138, 
       u1_u5_u2_n139, u1_u5_u2_n140, u1_u5_u2_n141, u1_u5_u2_n142, u1_u5_u2_n143, u1_u5_u2_n144, u1_u5_u2_n145, u1_u5_u2_n146, u1_u5_u2_n147, 
       u1_u5_u2_n148, u1_u5_u2_n149, u1_u5_u2_n150, u1_u5_u2_n151, u1_u5_u2_n152, u1_u5_u2_n153, u1_u5_u2_n154, u1_u5_u2_n155, u1_u5_u2_n156, 
       u1_u5_u2_n157, u1_u5_u2_n158, u1_u5_u2_n159, u1_u5_u2_n160, u1_u5_u2_n161, u1_u5_u2_n162, u1_u5_u2_n163, u1_u5_u2_n164, u1_u5_u2_n165, 
       u1_u5_u2_n166, u1_u5_u2_n167, u1_u5_u2_n168, u1_u5_u2_n169, u1_u5_u2_n170, u1_u5_u2_n171, u1_u5_u2_n172, u1_u5_u2_n173, u1_u5_u2_n174, 
       u1_u5_u2_n175, u1_u5_u2_n176, u1_u5_u2_n177, u1_u5_u2_n178, u1_u5_u2_n179, u1_u5_u2_n180, u1_u5_u2_n181, u1_u5_u2_n182, u1_u5_u2_n183, 
       u1_u5_u2_n184, u1_u5_u2_n185, u1_u5_u2_n186, u1_u5_u2_n187, u1_u5_u2_n188, u1_u5_u2_n95, u1_u5_u2_n96, u1_u5_u2_n97, u1_u5_u2_n98, 
       u1_u5_u2_n99, u1_u5_u3_n100, u1_u5_u3_n101, u1_u5_u3_n102, u1_u5_u3_n103, u1_u5_u3_n104, u1_u5_u3_n105, u1_u5_u3_n106, u1_u5_u3_n107, 
       u1_u5_u3_n108, u1_u5_u3_n109, u1_u5_u3_n110, u1_u5_u3_n111, u1_u5_u3_n112, u1_u5_u3_n113, u1_u5_u3_n114, u1_u5_u3_n115, u1_u5_u3_n116, 
       u1_u5_u3_n117, u1_u5_u3_n118, u1_u5_u3_n119, u1_u5_u3_n120, u1_u5_u3_n121, u1_u5_u3_n122, u1_u5_u3_n123, u1_u5_u3_n124, u1_u5_u3_n125, 
       u1_u5_u3_n126, u1_u5_u3_n127, u1_u5_u3_n128, u1_u5_u3_n129, u1_u5_u3_n130, u1_u5_u3_n131, u1_u5_u3_n132, u1_u5_u3_n133, u1_u5_u3_n134, 
       u1_u5_u3_n135, u1_u5_u3_n136, u1_u5_u3_n137, u1_u5_u3_n138, u1_u5_u3_n139, u1_u5_u3_n140, u1_u5_u3_n141, u1_u5_u3_n142, u1_u5_u3_n143, 
       u1_u5_u3_n144, u1_u5_u3_n145, u1_u5_u3_n146, u1_u5_u3_n147, u1_u5_u3_n148, u1_u5_u3_n149, u1_u5_u3_n150, u1_u5_u3_n151, u1_u5_u3_n152, 
       u1_u5_u3_n153, u1_u5_u3_n154, u1_u5_u3_n155, u1_u5_u3_n156, u1_u5_u3_n157, u1_u5_u3_n158, u1_u5_u3_n159, u1_u5_u3_n160, u1_u5_u3_n161, 
       u1_u5_u3_n162, u1_u5_u3_n163, u1_u5_u3_n164, u1_u5_u3_n165, u1_u5_u3_n166, u1_u5_u3_n167, u1_u5_u3_n168, u1_u5_u3_n169, u1_u5_u3_n170, 
       u1_u5_u3_n171, u1_u5_u3_n172, u1_u5_u3_n173, u1_u5_u3_n174, u1_u5_u3_n175, u1_u5_u3_n176, u1_u5_u3_n177, u1_u5_u3_n178, u1_u5_u3_n179, 
       u1_u5_u3_n180, u1_u5_u3_n181, u1_u5_u3_n182, u1_u5_u3_n183, u1_u5_u3_n184, u1_u5_u3_n185, u1_u5_u3_n186, u1_u5_u3_n94, u1_u5_u3_n95, 
       u1_u5_u3_n96, u1_u5_u3_n97, u1_u5_u3_n98, u1_u5_u3_n99, u1_u5_u4_n100, u1_u5_u4_n101, u1_u5_u4_n102, u1_u5_u4_n103, u1_u5_u4_n104, 
       u1_u5_u4_n105, u1_u5_u4_n106, u1_u5_u4_n107, u1_u5_u4_n108, u1_u5_u4_n109, u1_u5_u4_n110, u1_u5_u4_n111, u1_u5_u4_n112, u1_u5_u4_n113, 
       u1_u5_u4_n114, u1_u5_u4_n115, u1_u5_u4_n116, u1_u5_u4_n117, u1_u5_u4_n118, u1_u5_u4_n119, u1_u5_u4_n120, u1_u5_u4_n121, u1_u5_u4_n122, 
       u1_u5_u4_n123, u1_u5_u4_n124, u1_u5_u4_n125, u1_u5_u4_n126, u1_u5_u4_n127, u1_u5_u4_n128, u1_u5_u4_n129, u1_u5_u4_n130, u1_u5_u4_n131, 
       u1_u5_u4_n132, u1_u5_u4_n133, u1_u5_u4_n134, u1_u5_u4_n135, u1_u5_u4_n136, u1_u5_u4_n137, u1_u5_u4_n138, u1_u5_u4_n139, u1_u5_u4_n140, 
       u1_u5_u4_n141, u1_u5_u4_n142, u1_u5_u4_n143, u1_u5_u4_n144, u1_u5_u4_n145, u1_u5_u4_n146, u1_u5_u4_n147, u1_u5_u4_n148, u1_u5_u4_n149, 
       u1_u5_u4_n150, u1_u5_u4_n151, u1_u5_u4_n152, u1_u5_u4_n153, u1_u5_u4_n154, u1_u5_u4_n155, u1_u5_u4_n156, u1_u5_u4_n157, u1_u5_u4_n158, 
       u1_u5_u4_n159, u1_u5_u4_n160, u1_u5_u4_n161, u1_u5_u4_n162, u1_u5_u4_n163, u1_u5_u4_n164, u1_u5_u4_n165, u1_u5_u4_n166, u1_u5_u4_n167, 
       u1_u5_u4_n168, u1_u5_u4_n169, u1_u5_u4_n170, u1_u5_u4_n171, u1_u5_u4_n172, u1_u5_u4_n173, u1_u5_u4_n174, u1_u5_u4_n175, u1_u5_u4_n176, 
       u1_u5_u4_n177, u1_u5_u4_n178, u1_u5_u4_n179, u1_u5_u4_n180, u1_u5_u4_n181, u1_u5_u4_n182, u1_u5_u4_n183, u1_u5_u4_n184, u1_u5_u4_n185, 
       u1_u5_u4_n186, u1_u5_u4_n94, u1_u5_u4_n95, u1_u5_u4_n96, u1_u5_u4_n97, u1_u5_u4_n98, u1_u5_u4_n99, u1_u5_u5_n100, u1_u5_u5_n101, 
       u1_u5_u5_n102, u1_u5_u5_n103, u1_u5_u5_n104, u1_u5_u5_n105, u1_u5_u5_n106, u1_u5_u5_n107, u1_u5_u5_n108, u1_u5_u5_n109, u1_u5_u5_n110, 
       u1_u5_u5_n111, u1_u5_u5_n112, u1_u5_u5_n113, u1_u5_u5_n114, u1_u5_u5_n115, u1_u5_u5_n116, u1_u5_u5_n117, u1_u5_u5_n118, u1_u5_u5_n119, 
       u1_u5_u5_n120, u1_u5_u5_n121, u1_u5_u5_n122, u1_u5_u5_n123, u1_u5_u5_n124, u1_u5_u5_n125, u1_u5_u5_n126, u1_u5_u5_n127, u1_u5_u5_n128, 
       u1_u5_u5_n129, u1_u5_u5_n130, u1_u5_u5_n131, u1_u5_u5_n132, u1_u5_u5_n133, u1_u5_u5_n134, u1_u5_u5_n135, u1_u5_u5_n136, u1_u5_u5_n137, 
       u1_u5_u5_n138, u1_u5_u5_n139, u1_u5_u5_n140, u1_u5_u5_n141, u1_u5_u5_n142, u1_u5_u5_n143, u1_u5_u5_n144, u1_u5_u5_n145, u1_u5_u5_n146, 
       u1_u5_u5_n147, u1_u5_u5_n148, u1_u5_u5_n149, u1_u5_u5_n150, u1_u5_u5_n151, u1_u5_u5_n152, u1_u5_u5_n153, u1_u5_u5_n154, u1_u5_u5_n155, 
       u1_u5_u5_n156, u1_u5_u5_n157, u1_u5_u5_n158, u1_u5_u5_n159, u1_u5_u5_n160, u1_u5_u5_n161, u1_u5_u5_n162, u1_u5_u5_n163, u1_u5_u5_n164, 
       u1_u5_u5_n165, u1_u5_u5_n166, u1_u5_u5_n167, u1_u5_u5_n168, u1_u5_u5_n169, u1_u5_u5_n170, u1_u5_u5_n171, u1_u5_u5_n172, u1_u5_u5_n173, 
       u1_u5_u5_n174, u1_u5_u5_n175, u1_u5_u5_n176, u1_u5_u5_n177, u1_u5_u5_n178, u1_u5_u5_n179, u1_u5_u5_n180, u1_u5_u5_n181, u1_u5_u5_n182, 
       u1_u5_u5_n183, u1_u5_u5_n184, u1_u5_u5_n185, u1_u5_u5_n186, u1_u5_u5_n187, u1_u5_u5_n188, u1_u5_u5_n189, u1_u5_u5_n190, u1_u5_u5_n191, 
       u1_u5_u5_n192, u1_u5_u5_n193, u1_u5_u5_n194, u1_u5_u5_n195, u1_u5_u5_n196, u1_u5_u5_n99, u1_u5_u6_n100, u1_u5_u6_n101, u1_u5_u6_n102, 
       u1_u5_u6_n103, u1_u5_u6_n104, u1_u5_u6_n105, u1_u5_u6_n106, u1_u5_u6_n107, u1_u5_u6_n108, u1_u5_u6_n109, u1_u5_u6_n110, u1_u5_u6_n111, 
       u1_u5_u6_n112, u1_u5_u6_n113, u1_u5_u6_n114, u1_u5_u6_n115, u1_u5_u6_n116, u1_u5_u6_n117, u1_u5_u6_n118, u1_u5_u6_n119, u1_u5_u6_n120, 
       u1_u5_u6_n121, u1_u5_u6_n122, u1_u5_u6_n123, u1_u5_u6_n124, u1_u5_u6_n125, u1_u5_u6_n126, u1_u5_u6_n127, u1_u5_u6_n128, u1_u5_u6_n129, 
       u1_u5_u6_n130, u1_u5_u6_n131, u1_u5_u6_n132, u1_u5_u6_n133, u1_u5_u6_n134, u1_u5_u6_n135, u1_u5_u6_n136, u1_u5_u6_n137, u1_u5_u6_n138, 
       u1_u5_u6_n139, u1_u5_u6_n140, u1_u5_u6_n141, u1_u5_u6_n142, u1_u5_u6_n143, u1_u5_u6_n144, u1_u5_u6_n145, u1_u5_u6_n146, u1_u5_u6_n147, 
       u1_u5_u6_n148, u1_u5_u6_n149, u1_u5_u6_n150, u1_u5_u6_n151, u1_u5_u6_n152, u1_u5_u6_n153, u1_u5_u6_n154, u1_u5_u6_n155, u1_u5_u6_n156, 
       u1_u5_u6_n157, u1_u5_u6_n158, u1_u5_u6_n159, u1_u5_u6_n160, u1_u5_u6_n161, u1_u5_u6_n162, u1_u5_u6_n163, u1_u5_u6_n164, u1_u5_u6_n165, 
       u1_u5_u6_n166, u1_u5_u6_n167, u1_u5_u6_n168, u1_u5_u6_n169, u1_u5_u6_n170, u1_u5_u6_n171, u1_u5_u6_n172, u1_u5_u6_n173, u1_u5_u6_n174, 
       u1_u5_u6_n88, u1_u5_u6_n89, u1_u5_u6_n90, u1_u5_u6_n91, u1_u5_u6_n92, u1_u5_u6_n93, u1_u5_u6_n94, u1_u5_u6_n95, u1_u5_u6_n96, 
       u1_u5_u6_n97, u1_u5_u6_n98, u1_u5_u6_n99, u1_u8_X_1, u1_u8_X_10, u1_u8_X_11, u1_u8_X_12, u1_u8_X_13, u1_u8_X_14, 
       u1_u8_X_15, u1_u8_X_16, u1_u8_X_17, u1_u8_X_18, u1_u8_X_19, u1_u8_X_2, u1_u8_X_20, u1_u8_X_21, u1_u8_X_22, 
       u1_u8_X_23, u1_u8_X_24, u1_u8_X_3, u1_u8_X_4, u1_u8_X_5, u1_u8_X_6, u1_u8_X_7, u1_u8_X_8, u1_u8_X_9, 
       u1_u8_u0_n100, u1_u8_u0_n101, u1_u8_u0_n102, u1_u8_u0_n103, u1_u8_u0_n104, u1_u8_u0_n105, u1_u8_u0_n106, u1_u8_u0_n107, u1_u8_u0_n108, 
       u1_u8_u0_n109, u1_u8_u0_n110, u1_u8_u0_n111, u1_u8_u0_n112, u1_u8_u0_n113, u1_u8_u0_n114, u1_u8_u0_n115, u1_u8_u0_n116, u1_u8_u0_n117, 
       u1_u8_u0_n118, u1_u8_u0_n119, u1_u8_u0_n120, u1_u8_u0_n121, u1_u8_u0_n122, u1_u8_u0_n123, u1_u8_u0_n124, u1_u8_u0_n125, u1_u8_u0_n126, 
       u1_u8_u0_n127, u1_u8_u0_n128, u1_u8_u0_n129, u1_u8_u0_n130, u1_u8_u0_n131, u1_u8_u0_n132, u1_u8_u0_n133, u1_u8_u0_n134, u1_u8_u0_n135, 
       u1_u8_u0_n136, u1_u8_u0_n137, u1_u8_u0_n138, u1_u8_u0_n139, u1_u8_u0_n140, u1_u8_u0_n141, u1_u8_u0_n142, u1_u8_u0_n143, u1_u8_u0_n144, 
       u1_u8_u0_n145, u1_u8_u0_n146, u1_u8_u0_n147, u1_u8_u0_n148, u1_u8_u0_n149, u1_u8_u0_n150, u1_u8_u0_n151, u1_u8_u0_n152, u1_u8_u0_n153, 
       u1_u8_u0_n154, u1_u8_u0_n155, u1_u8_u0_n156, u1_u8_u0_n157, u1_u8_u0_n158, u1_u8_u0_n159, u1_u8_u0_n160, u1_u8_u0_n161, u1_u8_u0_n162, 
       u1_u8_u0_n163, u1_u8_u0_n164, u1_u8_u0_n165, u1_u8_u0_n166, u1_u8_u0_n167, u1_u8_u0_n168, u1_u8_u0_n169, u1_u8_u0_n170, u1_u8_u0_n171, 
       u1_u8_u0_n172, u1_u8_u0_n173, u1_u8_u0_n174, u1_u8_u0_n88, u1_u8_u0_n89, u1_u8_u0_n90, u1_u8_u0_n91, u1_u8_u0_n92, u1_u8_u0_n93, 
       u1_u8_u0_n94, u1_u8_u0_n95, u1_u8_u0_n96, u1_u8_u0_n97, u1_u8_u0_n98, u1_u8_u0_n99, u1_u8_u1_n100, u1_u8_u1_n101, u1_u8_u1_n102, 
       u1_u8_u1_n103, u1_u8_u1_n104, u1_u8_u1_n105, u1_u8_u1_n106, u1_u8_u1_n107, u1_u8_u1_n108, u1_u8_u1_n109, u1_u8_u1_n110, u1_u8_u1_n111, 
       u1_u8_u1_n112, u1_u8_u1_n113, u1_u8_u1_n114, u1_u8_u1_n115, u1_u8_u1_n116, u1_u8_u1_n117, u1_u8_u1_n118, u1_u8_u1_n119, u1_u8_u1_n120, 
       u1_u8_u1_n121, u1_u8_u1_n122, u1_u8_u1_n123, u1_u8_u1_n124, u1_u8_u1_n125, u1_u8_u1_n126, u1_u8_u1_n127, u1_u8_u1_n128, u1_u8_u1_n129, 
       u1_u8_u1_n130, u1_u8_u1_n131, u1_u8_u1_n132, u1_u8_u1_n133, u1_u8_u1_n134, u1_u8_u1_n135, u1_u8_u1_n136, u1_u8_u1_n137, u1_u8_u1_n138, 
       u1_u8_u1_n139, u1_u8_u1_n140, u1_u8_u1_n141, u1_u8_u1_n142, u1_u8_u1_n143, u1_u8_u1_n144, u1_u8_u1_n145, u1_u8_u1_n146, u1_u8_u1_n147, 
       u1_u8_u1_n148, u1_u8_u1_n149, u1_u8_u1_n150, u1_u8_u1_n151, u1_u8_u1_n152, u1_u8_u1_n153, u1_u8_u1_n154, u1_u8_u1_n155, u1_u8_u1_n156, 
       u1_u8_u1_n157, u1_u8_u1_n158, u1_u8_u1_n159, u1_u8_u1_n160, u1_u8_u1_n161, u1_u8_u1_n162, u1_u8_u1_n163, u1_u8_u1_n164, u1_u8_u1_n165, 
       u1_u8_u1_n166, u1_u8_u1_n167, u1_u8_u1_n168, u1_u8_u1_n169, u1_u8_u1_n170, u1_u8_u1_n171, u1_u8_u1_n172, u1_u8_u1_n173, u1_u8_u1_n174, 
       u1_u8_u1_n175, u1_u8_u1_n176, u1_u8_u1_n177, u1_u8_u1_n178, u1_u8_u1_n179, u1_u8_u1_n180, u1_u8_u1_n181, u1_u8_u1_n182, u1_u8_u1_n183, 
       u1_u8_u1_n184, u1_u8_u1_n185, u1_u8_u1_n186, u1_u8_u1_n187, u1_u8_u1_n188, u1_u8_u1_n95, u1_u8_u1_n96, u1_u8_u1_n97, u1_u8_u1_n98, 
       u1_u8_u1_n99, u1_u8_u2_n100, u1_u8_u2_n101, u1_u8_u2_n102, u1_u8_u2_n103, u1_u8_u2_n104, u1_u8_u2_n105, u1_u8_u2_n106, u1_u8_u2_n107, 
       u1_u8_u2_n108, u1_u8_u2_n109, u1_u8_u2_n110, u1_u8_u2_n111, u1_u8_u2_n112, u1_u8_u2_n113, u1_u8_u2_n114, u1_u8_u2_n115, u1_u8_u2_n116, 
       u1_u8_u2_n117, u1_u8_u2_n118, u1_u8_u2_n119, u1_u8_u2_n120, u1_u8_u2_n121, u1_u8_u2_n122, u1_u8_u2_n123, u1_u8_u2_n124, u1_u8_u2_n125, 
       u1_u8_u2_n126, u1_u8_u2_n127, u1_u8_u2_n128, u1_u8_u2_n129, u1_u8_u2_n130, u1_u8_u2_n131, u1_u8_u2_n132, u1_u8_u2_n133, u1_u8_u2_n134, 
       u1_u8_u2_n135, u1_u8_u2_n136, u1_u8_u2_n137, u1_u8_u2_n138, u1_u8_u2_n139, u1_u8_u2_n140, u1_u8_u2_n141, u1_u8_u2_n142, u1_u8_u2_n143, 
       u1_u8_u2_n144, u1_u8_u2_n145, u1_u8_u2_n146, u1_u8_u2_n147, u1_u8_u2_n148, u1_u8_u2_n149, u1_u8_u2_n150, u1_u8_u2_n151, u1_u8_u2_n152, 
       u1_u8_u2_n153, u1_u8_u2_n154, u1_u8_u2_n155, u1_u8_u2_n156, u1_u8_u2_n157, u1_u8_u2_n158, u1_u8_u2_n159, u1_u8_u2_n160, u1_u8_u2_n161, 
       u1_u8_u2_n162, u1_u8_u2_n163, u1_u8_u2_n164, u1_u8_u2_n165, u1_u8_u2_n166, u1_u8_u2_n167, u1_u8_u2_n168, u1_u8_u2_n169, u1_u8_u2_n170, 
       u1_u8_u2_n171, u1_u8_u2_n172, u1_u8_u2_n173, u1_u8_u2_n174, u1_u8_u2_n175, u1_u8_u2_n176, u1_u8_u2_n177, u1_u8_u2_n178, u1_u8_u2_n179, 
       u1_u8_u2_n180, u1_u8_u2_n181, u1_u8_u2_n182, u1_u8_u2_n183, u1_u8_u2_n184, u1_u8_u2_n185, u1_u8_u2_n186, u1_u8_u2_n187, u1_u8_u2_n188, 
       u1_u8_u2_n95, u1_u8_u2_n96, u1_u8_u2_n97, u1_u8_u2_n98, u1_u8_u2_n99, u1_u8_u3_n100, u1_u8_u3_n101, u1_u8_u3_n102, u1_u8_u3_n103, 
       u1_u8_u3_n104, u1_u8_u3_n105, u1_u8_u3_n106, u1_u8_u3_n107, u1_u8_u3_n108, u1_u8_u3_n109, u1_u8_u3_n110, u1_u8_u3_n111, u1_u8_u3_n112, 
       u1_u8_u3_n113, u1_u8_u3_n114, u1_u8_u3_n115, u1_u8_u3_n116, u1_u8_u3_n117, u1_u8_u3_n118, u1_u8_u3_n119, u1_u8_u3_n120, u1_u8_u3_n121, 
       u1_u8_u3_n122, u1_u8_u3_n123, u1_u8_u3_n124, u1_u8_u3_n125, u1_u8_u3_n126, u1_u8_u3_n127, u1_u8_u3_n128, u1_u8_u3_n129, u1_u8_u3_n130, 
       u1_u8_u3_n131, u1_u8_u3_n132, u1_u8_u3_n133, u1_u8_u3_n134, u1_u8_u3_n135, u1_u8_u3_n136, u1_u8_u3_n137, u1_u8_u3_n138, u1_u8_u3_n139, 
       u1_u8_u3_n140, u1_u8_u3_n141, u1_u8_u3_n142, u1_u8_u3_n143, u1_u8_u3_n144, u1_u8_u3_n145, u1_u8_u3_n146, u1_u8_u3_n147, u1_u8_u3_n148, 
       u1_u8_u3_n149, u1_u8_u3_n150, u1_u8_u3_n151, u1_u8_u3_n152, u1_u8_u3_n153, u1_u8_u3_n154, u1_u8_u3_n155, u1_u8_u3_n156, u1_u8_u3_n157, 
       u1_u8_u3_n158, u1_u8_u3_n159, u1_u8_u3_n160, u1_u8_u3_n161, u1_u8_u3_n162, u1_u8_u3_n163, u1_u8_u3_n164, u1_u8_u3_n165, u1_u8_u3_n166, 
       u1_u8_u3_n167, u1_u8_u3_n168, u1_u8_u3_n169, u1_u8_u3_n170, u1_u8_u3_n171, u1_u8_u3_n172, u1_u8_u3_n173, u1_u8_u3_n174, u1_u8_u3_n175, 
       u1_u8_u3_n176, u1_u8_u3_n177, u1_u8_u3_n178, u1_u8_u3_n179, u1_u8_u3_n180, u1_u8_u3_n181, u1_u8_u3_n182, u1_u8_u3_n183, u1_u8_u3_n184, 
       u1_u8_u3_n185, u1_u8_u3_n186, u1_u8_u3_n94, u1_u8_u3_n95, u1_u8_u3_n96, u1_u8_u3_n97, u1_u8_u3_n98, u1_u8_u3_n99, u1_u9_X_43, 
       u1_u9_X_44, u1_u9_X_45, u1_u9_X_46, u1_u9_X_47, u1_u9_X_48, u1_u9_u7_n100, u1_u9_u7_n101, u1_u9_u7_n102, u1_u9_u7_n103, 
       u1_u9_u7_n104, u1_u9_u7_n105, u1_u9_u7_n106, u1_u9_u7_n107, u1_u9_u7_n108, u1_u9_u7_n109, u1_u9_u7_n110, u1_u9_u7_n111, u1_u9_u7_n112, 
       u1_u9_u7_n113, u1_u9_u7_n114, u1_u9_u7_n115, u1_u9_u7_n116, u1_u9_u7_n117, u1_u9_u7_n118, u1_u9_u7_n119, u1_u9_u7_n120, u1_u9_u7_n121, 
       u1_u9_u7_n122, u1_u9_u7_n123, u1_u9_u7_n124, u1_u9_u7_n125, u1_u9_u7_n126, u1_u9_u7_n127, u1_u9_u7_n128, u1_u9_u7_n129, u1_u9_u7_n130, 
       u1_u9_u7_n131, u1_u9_u7_n132, u1_u9_u7_n133, u1_u9_u7_n134, u1_u9_u7_n135, u1_u9_u7_n136, u1_u9_u7_n137, u1_u9_u7_n138, u1_u9_u7_n139, 
       u1_u9_u7_n140, u1_u9_u7_n141, u1_u9_u7_n142, u1_u9_u7_n143, u1_u9_u7_n144, u1_u9_u7_n145, u1_u9_u7_n146, u1_u9_u7_n147, u1_u9_u7_n148, 
       u1_u9_u7_n149, u1_u9_u7_n150, u1_u9_u7_n151, u1_u9_u7_n152, u1_u9_u7_n153, u1_u9_u7_n154, u1_u9_u7_n155, u1_u9_u7_n156, u1_u9_u7_n157, 
       u1_u9_u7_n158, u1_u9_u7_n159, u1_u9_u7_n160, u1_u9_u7_n161, u1_u9_u7_n162, u1_u9_u7_n163, u1_u9_u7_n164, u1_u9_u7_n165, u1_u9_u7_n166, 
       u1_u9_u7_n167, u1_u9_u7_n168, u1_u9_u7_n169, u1_u9_u7_n170, u1_u9_u7_n171, u1_u9_u7_n172, u1_u9_u7_n173, u1_u9_u7_n174, u1_u9_u7_n175, 
       u1_u9_u7_n176, u1_u9_u7_n177, u1_u9_u7_n178, u1_u9_u7_n179, u1_u9_u7_n180, u1_u9_u7_n91, u1_u9_u7_n92, u1_u9_u7_n93, u1_u9_u7_n94, 
       u1_u9_u7_n95, u1_u9_u7_n96, u1_u9_u7_n97, u1_u9_u7_n98, u1_u9_u7_n99, u1_uk_n1005, u1_uk_n1006, u1_uk_n1007, u1_uk_n1009, 
       u1_uk_n1010, u1_uk_n1011, u1_uk_n1012, u1_uk_n1013, u1_uk_n1014, u1_uk_n1015, u1_uk_n1016, u1_uk_n1017, u1_uk_n1018, 
       u1_uk_n1019, u1_uk_n1050, u1_uk_n1070, u1_uk_n1077, u1_uk_n1078, u1_uk_n1079, u1_uk_n1080, u1_uk_n1089, u1_uk_n1090, 
       u1_uk_n1091, u1_uk_n1092, u1_uk_n1093, u1_uk_n1094, u1_uk_n1095, u1_uk_n1096, u1_uk_n1097, u1_uk_n1098, u1_uk_n1099, 
       u1_uk_n1101, u1_uk_n1147, u1_uk_n1148, u1_uk_n1149, u1_uk_n1150, u1_uk_n1151, u1_uk_n1152, u1_uk_n1153, u1_uk_n1154, 
       u1_uk_n1155, u1_uk_n1156, u1_uk_n1157, u1_uk_n1160, u1_uk_n1171, u1_uk_n1172, u1_uk_n1173, u1_uk_n1174, u1_uk_n1177, 
       u1_uk_n1178, u1_uk_n1179, u1_uk_n1181, u1_uk_n1182, u1_uk_n1187, u1_uk_n1188, u1_uk_n1195, u1_uk_n1201, u1_uk_n1208, 
       u1_uk_n1213, u1_uk_n971, u1_uk_n972, u1_uk_n973, u1_uk_n974, u1_uk_n975, u2_K2_13, u2_K2_14, u2_K2_15, 
       u2_K2_17, u2_K9_31, u2_K9_33, u2_K9_34, u2_K9_35, u2_K9_37, u2_K9_39, u2_K9_41, u2_K9_42, 
       u2_out1_16, u2_out1_24, u2_out1_30, u2_out1_6, u2_out8_11, u2_out8_12, u2_out8_19, u2_out8_22, u2_out8_29, 
       u2_out8_32, u2_out8_4, u2_out8_7, u2_u1_X_13, u2_u1_X_14, u2_u1_X_15, u2_u1_X_16, u2_u1_X_17, u2_u1_X_18, 
       u2_u1_u2_n100, u2_u1_u2_n101, u2_u1_u2_n102, u2_u1_u2_n103, u2_u1_u2_n104, u2_u1_u2_n105, u2_u1_u2_n106, u2_u1_u2_n107, u2_u1_u2_n108, 
       u2_u1_u2_n109, u2_u1_u2_n110, u2_u1_u2_n111, u2_u1_u2_n112, u2_u1_u2_n113, u2_u1_u2_n114, u2_u1_u2_n115, u2_u1_u2_n116, u2_u1_u2_n117, 
       u2_u1_u2_n118, u2_u1_u2_n119, u2_u1_u2_n120, u2_u1_u2_n121, u2_u1_u2_n122, u2_u1_u2_n123, u2_u1_u2_n124, u2_u1_u2_n125, u2_u1_u2_n126, 
       u2_u1_u2_n127, u2_u1_u2_n128, u2_u1_u2_n129, u2_u1_u2_n130, u2_u1_u2_n131, u2_u1_u2_n132, u2_u1_u2_n133, u2_u1_u2_n134, u2_u1_u2_n135, 
       u2_u1_u2_n136, u2_u1_u2_n137, u2_u1_u2_n138, u2_u1_u2_n139, u2_u1_u2_n140, u2_u1_u2_n141, u2_u1_u2_n142, u2_u1_u2_n143, u2_u1_u2_n144, 
       u2_u1_u2_n145, u2_u1_u2_n146, u2_u1_u2_n147, u2_u1_u2_n148, u2_u1_u2_n149, u2_u1_u2_n150, u2_u1_u2_n151, u2_u1_u2_n152, u2_u1_u2_n153, 
       u2_u1_u2_n154, u2_u1_u2_n155, u2_u1_u2_n156, u2_u1_u2_n157, u2_u1_u2_n158, u2_u1_u2_n159, u2_u1_u2_n160, u2_u1_u2_n161, u2_u1_u2_n162, 
       u2_u1_u2_n163, u2_u1_u2_n164, u2_u1_u2_n165, u2_u1_u2_n166, u2_u1_u2_n167, u2_u1_u2_n168, u2_u1_u2_n169, u2_u1_u2_n170, u2_u1_u2_n171, 
       u2_u1_u2_n172, u2_u1_u2_n173, u2_u1_u2_n174, u2_u1_u2_n175, u2_u1_u2_n176, u2_u1_u2_n177, u2_u1_u2_n178, u2_u1_u2_n179, u2_u1_u2_n180, 
       u2_u1_u2_n181, u2_u1_u2_n182, u2_u1_u2_n183, u2_u1_u2_n184, u2_u1_u2_n185, u2_u1_u2_n186, u2_u1_u2_n187, u2_u1_u2_n188, u2_u1_u2_n95, 
       u2_u1_u2_n96, u2_u1_u2_n97, u2_u1_u2_n98, u2_u1_u2_n99, u2_u8_X_31, u2_u8_X_32, u2_u8_X_33, u2_u8_X_34, u2_u8_X_35, 
       u2_u8_X_36, u2_u8_X_37, u2_u8_X_38, u2_u8_X_39, u2_u8_X_40, u2_u8_X_41, u2_u8_X_42, u2_u8_u5_n100, u2_u8_u5_n101, 
       u2_u8_u5_n102, u2_u8_u5_n103, u2_u8_u5_n104, u2_u8_u5_n105, u2_u8_u5_n106, u2_u8_u5_n107, u2_u8_u5_n108, u2_u8_u5_n109, u2_u8_u5_n110, 
       u2_u8_u5_n111, u2_u8_u5_n112, u2_u8_u5_n113, u2_u8_u5_n114, u2_u8_u5_n115, u2_u8_u5_n116, u2_u8_u5_n117, u2_u8_u5_n118, u2_u8_u5_n119, 
       u2_u8_u5_n120, u2_u8_u5_n121, u2_u8_u5_n122, u2_u8_u5_n123, u2_u8_u5_n124, u2_u8_u5_n125, u2_u8_u5_n126, u2_u8_u5_n127, u2_u8_u5_n128, 
       u2_u8_u5_n129, u2_u8_u5_n130, u2_u8_u5_n131, u2_u8_u5_n132, u2_u8_u5_n133, u2_u8_u5_n134, u2_u8_u5_n135, u2_u8_u5_n136, u2_u8_u5_n137, 
       u2_u8_u5_n138, u2_u8_u5_n139, u2_u8_u5_n140, u2_u8_u5_n141, u2_u8_u5_n142, u2_u8_u5_n143, u2_u8_u5_n144, u2_u8_u5_n145, u2_u8_u5_n146, 
       u2_u8_u5_n147, u2_u8_u5_n148, u2_u8_u5_n149, u2_u8_u5_n150, u2_u8_u5_n151, u2_u8_u5_n152, u2_u8_u5_n153, u2_u8_u5_n154, u2_u8_u5_n155, 
       u2_u8_u5_n156, u2_u8_u5_n157, u2_u8_u5_n158, u2_u8_u5_n159, u2_u8_u5_n160, u2_u8_u5_n161, u2_u8_u5_n162, u2_u8_u5_n163, u2_u8_u5_n164, 
       u2_u8_u5_n165, u2_u8_u5_n166, u2_u8_u5_n167, u2_u8_u5_n168, u2_u8_u5_n169, u2_u8_u5_n170, u2_u8_u5_n171, u2_u8_u5_n172, u2_u8_u5_n173, 
       u2_u8_u5_n174, u2_u8_u5_n175, u2_u8_u5_n176, u2_u8_u5_n177, u2_u8_u5_n178, u2_u8_u5_n179, u2_u8_u5_n180, u2_u8_u5_n181, u2_u8_u5_n182, 
       u2_u8_u5_n183, u2_u8_u5_n184, u2_u8_u5_n185, u2_u8_u5_n186, u2_u8_u5_n187, u2_u8_u5_n188, u2_u8_u5_n189, u2_u8_u5_n190, u2_u8_u5_n191, 
       u2_u8_u5_n192, u2_u8_u5_n193, u2_u8_u5_n194, u2_u8_u5_n195, u2_u8_u5_n196, u2_u8_u5_n99, u2_u8_u6_n100, u2_u8_u6_n101, u2_u8_u6_n102, 
       u2_u8_u6_n103, u2_u8_u6_n104, u2_u8_u6_n105, u2_u8_u6_n106, u2_u8_u6_n107, u2_u8_u6_n108, u2_u8_u6_n109, u2_u8_u6_n110, u2_u8_u6_n111, 
       u2_u8_u6_n112, u2_u8_u6_n113, u2_u8_u6_n114, u2_u8_u6_n115, u2_u8_u6_n116, u2_u8_u6_n117, u2_u8_u6_n118, u2_u8_u6_n119, u2_u8_u6_n120, 
       u2_u8_u6_n121, u2_u8_u6_n122, u2_u8_u6_n123, u2_u8_u6_n124, u2_u8_u6_n125, u2_u8_u6_n126, u2_u8_u6_n127, u2_u8_u6_n128, u2_u8_u6_n129, 
       u2_u8_u6_n130, u2_u8_u6_n131, u2_u8_u6_n132, u2_u8_u6_n133, u2_u8_u6_n134, u2_u8_u6_n135, u2_u8_u6_n136, u2_u8_u6_n137, u2_u8_u6_n138, 
       u2_u8_u6_n139, u2_u8_u6_n140, u2_u8_u6_n141, u2_u8_u6_n142, u2_u8_u6_n143, u2_u8_u6_n144, u2_u8_u6_n145, u2_u8_u6_n146, u2_u8_u6_n147, 
       u2_u8_u6_n148, u2_u8_u6_n149, u2_u8_u6_n150, u2_u8_u6_n151, u2_u8_u6_n152, u2_u8_u6_n153, u2_u8_u6_n154, u2_u8_u6_n155, u2_u8_u6_n156, 
       u2_u8_u6_n157, u2_u8_u6_n158, u2_u8_u6_n159, u2_u8_u6_n160, u2_u8_u6_n161, u2_u8_u6_n162, u2_u8_u6_n163, u2_u8_u6_n164, u2_u8_u6_n165, 
       u2_u8_u6_n166, u2_u8_u6_n167, u2_u8_u6_n168, u2_u8_u6_n169, u2_u8_u6_n170, u2_u8_u6_n171, u2_u8_u6_n172, u2_u8_u6_n173, u2_u8_u6_n174, 
       u2_u8_u6_n88, u2_u8_u6_n89, u2_u8_u6_n90, u2_u8_u6_n91, u2_u8_u6_n92, u2_u8_u6_n93, u2_u8_u6_n94, u2_u8_u6_n95, u2_u8_u6_n96, 
       u2_u8_u6_n97, u2_u8_u6_n98, u2_u8_u6_n99, u2_uk_n1133, u2_uk_n1135,  u2_uk_n993;
  XOR2_X1 u0_U101 (.B( u0_L12_26 ) , .Z( u0_N441 ) , .A( u0_out13_26 ) );
  XOR2_X1 u0_U102 (.B( u0_L12_25 ) , .Z( u0_N440 ) , .A( u0_out13_25 ) );
  XOR2_X1 u0_U104 (.B( u0_L12_24 ) , .Z( u0_N439 ) , .A( u0_out13_24 ) );
  XOR2_X1 u0_U108 (.B( u0_L12_20 ) , .Z( u0_N435 ) , .A( u0_out13_20 ) );
  XOR2_X1 u0_U110 (.B( u0_L12_18 ) , .Z( u0_N433 ) , .A( u0_out13_18 ) );
  XOR2_X1 u0_U112 (.B( u0_L12_16 ) , .Z( u0_N431 ) , .A( u0_out13_16 ) );
  XOR2_X1 u0_U115 (.B( u0_L12_14 ) , .Z( u0_N429 ) , .A( u0_out13_14 ) );
  XOR2_X1 u0_U116 (.B( u0_L12_13 ) , .Z( u0_N428 ) , .A( u0_out13_13 ) );
  XOR2_X1 u0_U119 (.B( u0_L12_10 ) , .Z( u0_N425 ) , .A( u0_out13_10 ) );
  XOR2_X1 u0_U121 (.B( u0_L12_8 ) , .Z( u0_N423 ) , .A( u0_out13_8 ) );
  XOR2_X1 u0_U123 (.B( u0_L12_6 ) , .Z( u0_N421 ) , .A( u0_out13_6 ) );
  XOR2_X1 u0_U127 (.B( u0_L12_3 ) , .Z( u0_N418 ) , .A( u0_out13_3 ) );
  XOR2_X1 u0_U128 (.B( u0_L12_2 ) , .Z( u0_N417 ) , .A( u0_out13_2 ) );
  XOR2_X1 u0_U129 (.B( u0_L12_1 ) , .Z( u0_N416 ) , .A( u0_out13_1 ) );
  XOR2_X1 u0_U240 (.B( u0_L8_29 ) , .Z( u0_N316 ) , .A( u0_out9_29 ) );
  XOR2_X1 u0_U242 (.B( u0_L8_27 ) , .Z( u0_N314 ) , .A( u0_out9_27 ) );
  XOR2_X1 u0_U244 (.B( u0_L8_25 ) , .Z( u0_N312 ) , .A( u0_out9_25 ) );
  XOR2_X1 u0_U249 (.B( u0_L8_21 ) , .Z( u0_N308 ) , .A( u0_out9_21 ) );
  XOR2_X1 u0_U251 (.B( u0_L8_19 ) , .Z( u0_N306 ) , .A( u0_out9_19 ) );
  XOR2_X1 u0_U255 (.B( u0_L8_15 ) , .Z( u0_N302 ) , .A( u0_out9_15 ) );
  XOR2_X1 u0_U256 (.B( u0_L8_14 ) , .Z( u0_N301 ) , .A( u0_out9_14 ) );
  XOR2_X1 u0_U261 (.B( u0_L8_11 ) , .Z( u0_N298 ) , .A( u0_out9_11 ) );
  XOR2_X1 u0_U264 (.B( u0_L8_8 ) , .Z( u0_N295 ) , .A( u0_out9_8 ) );
  XOR2_X1 u0_U267 (.B( u0_L8_5 ) , .Z( u0_N292 ) , .A( u0_out9_5 ) );
  XOR2_X1 u0_U268 (.B( u0_L8_4 ) , .Z( u0_N291 ) , .A( u0_out9_4 ) );
  XOR2_X1 u0_U269 (.B( u0_L8_3 ) , .Z( u0_N290 ) , .A( u0_out9_3 ) );
  XOR2_X1 u0_U97 (.B( u0_L12_30 ) , .Z( u0_N445 ) , .A( u0_out13_30 ) );
  XOR2_X1 u0_U99 (.B( u0_L12_28 ) , .Z( u0_N443 ) , .A( u0_out13_28 ) );
  XOR2_X1 u0_u13_U1 (.B( u0_K14_9 ) , .A( u0_R12_6 ) , .Z( u0_u13_X_9 ) );
  XOR2_X1 u0_u13_U2 (.B( u0_K14_8 ) , .A( u0_R12_5 ) , .Z( u0_u13_X_8 ) );
  XOR2_X1 u0_u13_U26 (.B( u0_K14_30 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_30 ) );
  XOR2_X1 u0_u13_U28 (.B( u0_K14_29 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_29 ) );
  XOR2_X1 u0_u13_U29 (.B( u0_K14_28 ) , .A( u0_R12_19 ) , .Z( u0_u13_X_28 ) );
  XOR2_X1 u0_u13_U3 (.B( u0_K14_7 ) , .A( u0_R12_4 ) , .Z( u0_u13_X_7 ) );
  XOR2_X1 u0_u13_U30 (.B( u0_K14_27 ) , .A( u0_R12_18 ) , .Z( u0_u13_X_27 ) );
  XOR2_X1 u0_u13_U31 (.B( u0_K14_26 ) , .A( u0_R12_17 ) , .Z( u0_u13_X_26 ) );
  XOR2_X1 u0_u13_U32 (.B( u0_K14_25 ) , .A( u0_R12_16 ) , .Z( u0_u13_X_25 ) );
  XOR2_X1 u0_u13_U33 (.B( u0_K14_24 ) , .A( u0_R12_17 ) , .Z( u0_u13_X_24 ) );
  XOR2_X1 u0_u13_U34 (.B( u0_K14_23 ) , .A( u0_R12_16 ) , .Z( u0_u13_X_23 ) );
  XOR2_X1 u0_u13_U35 (.B( u0_K14_22 ) , .A( u0_R12_15 ) , .Z( u0_u13_X_22 ) );
  XOR2_X1 u0_u13_U36 (.B( u0_K14_21 ) , .A( u0_R12_14 ) , .Z( u0_u13_X_21 ) );
  XOR2_X1 u0_u13_U37 (.B( u0_K14_20 ) , .A( u0_R12_13 ) , .Z( u0_u13_X_20 ) );
  XOR2_X1 u0_u13_U39 (.B( u0_K14_19 ) , .A( u0_R12_12 ) , .Z( u0_u13_X_19 ) );
  XOR2_X1 u0_u13_U40 (.B( u0_K14_18 ) , .A( u0_R12_13 ) , .Z( u0_u13_X_18 ) );
  XOR2_X1 u0_u13_U41 (.B( u0_K14_17 ) , .A( u0_R12_12 ) , .Z( u0_u13_X_17 ) );
  XOR2_X1 u0_u13_U42 (.B( u0_K14_16 ) , .A( u0_R12_11 ) , .Z( u0_u13_X_16 ) );
  XOR2_X1 u0_u13_U43 (.B( u0_K14_15 ) , .A( u0_R12_10 ) , .Z( u0_u13_X_15 ) );
  XOR2_X1 u0_u13_U44 (.B( u0_K14_14 ) , .A( u0_R12_9 ) , .Z( u0_u13_X_14 ) );
  XOR2_X1 u0_u13_U45 (.B( u0_K14_13 ) , .A( u0_R12_8 ) , .Z( u0_u13_X_13 ) );
  XOR2_X1 u0_u13_U46 (.B( u0_K14_12 ) , .A( u0_R12_9 ) , .Z( u0_u13_X_12 ) );
  XOR2_X1 u0_u13_U47 (.B( u0_K14_11 ) , .A( u0_R12_8 ) , .Z( u0_u13_X_11 ) );
  XOR2_X1 u0_u13_U48 (.B( u0_K14_10 ) , .A( u0_R12_7 ) , .Z( u0_u13_X_10 ) );
  AOI21_X1 u0_u13_u1_U10 (.B2( u0_u13_u1_n155 ) , .B1( u0_u13_u1_n156 ) , .ZN( u0_u13_u1_n157 ) , .A( u0_u13_u1_n174 ) );
  NAND3_X1 u0_u13_u1_U100 (.ZN( u0_u13_u1_n113 ) , .A1( u0_u13_u1_n120 ) , .A3( u0_u13_u1_n133 ) , .A2( u0_u13_u1_n155 ) );
  NAND2_X1 u0_u13_u1_U11 (.ZN( u0_u13_u1_n140 ) , .A2( u0_u13_u1_n150 ) , .A1( u0_u13_u1_n155 ) );
  NAND2_X1 u0_u13_u1_U12 (.A1( u0_u13_u1_n131 ) , .ZN( u0_u13_u1_n147 ) , .A2( u0_u13_u1_n153 ) );
  INV_X1 u0_u13_u1_U13 (.A( u0_u13_u1_n139 ) , .ZN( u0_u13_u1_n174 ) );
  OR4_X1 u0_u13_u1_U14 (.A4( u0_u13_u1_n106 ) , .A3( u0_u13_u1_n107 ) , .ZN( u0_u13_u1_n108 ) , .A1( u0_u13_u1_n117 ) , .A2( u0_u13_u1_n184 ) );
  AOI21_X1 u0_u13_u1_U15 (.ZN( u0_u13_u1_n106 ) , .A( u0_u13_u1_n112 ) , .B1( u0_u13_u1_n154 ) , .B2( u0_u13_u1_n156 ) );
  AOI21_X1 u0_u13_u1_U16 (.ZN( u0_u13_u1_n107 ) , .B1( u0_u13_u1_n134 ) , .B2( u0_u13_u1_n149 ) , .A( u0_u13_u1_n174 ) );
  INV_X1 u0_u13_u1_U17 (.A( u0_u13_u1_n101 ) , .ZN( u0_u13_u1_n184 ) );
  INV_X1 u0_u13_u1_U18 (.A( u0_u13_u1_n112 ) , .ZN( u0_u13_u1_n171 ) );
  NAND2_X1 u0_u13_u1_U19 (.ZN( u0_u13_u1_n141 ) , .A1( u0_u13_u1_n153 ) , .A2( u0_u13_u1_n156 ) );
  AND2_X1 u0_u13_u1_U20 (.A1( u0_u13_u1_n123 ) , .ZN( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n161 ) );
  NAND2_X1 u0_u13_u1_U21 (.A2( u0_u13_u1_n115 ) , .A1( u0_u13_u1_n116 ) , .ZN( u0_u13_u1_n148 ) );
  NAND2_X1 u0_u13_u1_U22 (.A2( u0_u13_u1_n133 ) , .A1( u0_u13_u1_n135 ) , .ZN( u0_u13_u1_n159 ) );
  NAND2_X1 u0_u13_u1_U23 (.A2( u0_u13_u1_n115 ) , .A1( u0_u13_u1_n120 ) , .ZN( u0_u13_u1_n132 ) );
  INV_X1 u0_u13_u1_U24 (.A( u0_u13_u1_n154 ) , .ZN( u0_u13_u1_n178 ) );
  AOI22_X1 u0_u13_u1_U25 (.B2( u0_u13_u1_n113 ) , .A2( u0_u13_u1_n114 ) , .ZN( u0_u13_u1_n125 ) , .A1( u0_u13_u1_n171 ) , .B1( u0_u13_u1_n173 ) );
  NAND2_X1 u0_u13_u1_U26 (.ZN( u0_u13_u1_n114 ) , .A1( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n156 ) );
  INV_X1 u0_u13_u1_U27 (.A( u0_u13_u1_n151 ) , .ZN( u0_u13_u1_n183 ) );
  AND2_X1 u0_u13_u1_U28 (.A1( u0_u13_u1_n129 ) , .A2( u0_u13_u1_n133 ) , .ZN( u0_u13_u1_n149 ) );
  INV_X1 u0_u13_u1_U29 (.A( u0_u13_u1_n131 ) , .ZN( u0_u13_u1_n180 ) );
  INV_X1 u0_u13_u1_U3 (.A( u0_u13_u1_n159 ) , .ZN( u0_u13_u1_n182 ) );
  OAI221_X1 u0_u13_u1_U30 (.A( u0_u13_u1_n119 ) , .C2( u0_u13_u1_n129 ) , .ZN( u0_u13_u1_n138 ) , .B2( u0_u13_u1_n152 ) , .C1( u0_u13_u1_n174 ) , .B1( u0_u13_u1_n187 ) );
  INV_X1 u0_u13_u1_U31 (.A( u0_u13_u1_n148 ) , .ZN( u0_u13_u1_n187 ) );
  AOI211_X1 u0_u13_u1_U32 (.B( u0_u13_u1_n117 ) , .A( u0_u13_u1_n118 ) , .ZN( u0_u13_u1_n119 ) , .C2( u0_u13_u1_n146 ) , .C1( u0_u13_u1_n159 ) );
  NOR2_X1 u0_u13_u1_U33 (.A1( u0_u13_u1_n168 ) , .A2( u0_u13_u1_n176 ) , .ZN( u0_u13_u1_n98 ) );
  AOI211_X1 u0_u13_u1_U34 (.B( u0_u13_u1_n162 ) , .A( u0_u13_u1_n163 ) , .C2( u0_u13_u1_n164 ) , .ZN( u0_u13_u1_n165 ) , .C1( u0_u13_u1_n171 ) );
  AOI21_X1 u0_u13_u1_U35 (.A( u0_u13_u1_n160 ) , .B2( u0_u13_u1_n161 ) , .ZN( u0_u13_u1_n162 ) , .B1( u0_u13_u1_n182 ) );
  OR2_X1 u0_u13_u1_U36 (.A2( u0_u13_u1_n157 ) , .A1( u0_u13_u1_n158 ) , .ZN( u0_u13_u1_n163 ) );
  OAI21_X1 u0_u13_u1_U37 (.B2( u0_u13_u1_n123 ) , .ZN( u0_u13_u1_n145 ) , .B1( u0_u13_u1_n160 ) , .A( u0_u13_u1_n185 ) );
  INV_X1 u0_u13_u1_U38 (.A( u0_u13_u1_n122 ) , .ZN( u0_u13_u1_n185 ) );
  AOI21_X1 u0_u13_u1_U39 (.B2( u0_u13_u1_n120 ) , .B1( u0_u13_u1_n121 ) , .ZN( u0_u13_u1_n122 ) , .A( u0_u13_u1_n128 ) );
  AOI221_X1 u0_u13_u1_U4 (.A( u0_u13_u1_n138 ) , .C2( u0_u13_u1_n139 ) , .C1( u0_u13_u1_n140 ) , .B2( u0_u13_u1_n141 ) , .ZN( u0_u13_u1_n142 ) , .B1( u0_u13_u1_n175 ) );
  NAND2_X1 u0_u13_u1_U40 (.A1( u0_u13_u1_n128 ) , .ZN( u0_u13_u1_n146 ) , .A2( u0_u13_u1_n160 ) );
  NAND2_X1 u0_u13_u1_U41 (.A2( u0_u13_u1_n112 ) , .ZN( u0_u13_u1_n139 ) , .A1( u0_u13_u1_n152 ) );
  NAND2_X1 u0_u13_u1_U42 (.A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n156 ) , .A2( u0_u13_u1_n99 ) );
  AOI221_X1 u0_u13_u1_U43 (.B1( u0_u13_u1_n140 ) , .ZN( u0_u13_u1_n167 ) , .B2( u0_u13_u1_n172 ) , .C2( u0_u13_u1_n175 ) , .C1( u0_u13_u1_n178 ) , .A( u0_u13_u1_n188 ) );
  INV_X1 u0_u13_u1_U44 (.ZN( u0_u13_u1_n188 ) , .A( u0_u13_u1_n97 ) );
  AOI211_X1 u0_u13_u1_U45 (.A( u0_u13_u1_n118 ) , .C1( u0_u13_u1_n132 ) , .C2( u0_u13_u1_n139 ) , .B( u0_u13_u1_n96 ) , .ZN( u0_u13_u1_n97 ) );
  AOI21_X1 u0_u13_u1_U46 (.B2( u0_u13_u1_n121 ) , .B1( u0_u13_u1_n135 ) , .A( u0_u13_u1_n152 ) , .ZN( u0_u13_u1_n96 ) );
  NOR2_X1 u0_u13_u1_U47 (.ZN( u0_u13_u1_n117 ) , .A1( u0_u13_u1_n121 ) , .A2( u0_u13_u1_n160 ) );
  AOI21_X1 u0_u13_u1_U48 (.A( u0_u13_u1_n128 ) , .B2( u0_u13_u1_n129 ) , .ZN( u0_u13_u1_n130 ) , .B1( u0_u13_u1_n150 ) );
  NAND2_X1 u0_u13_u1_U49 (.ZN( u0_u13_u1_n112 ) , .A1( u0_u13_u1_n169 ) , .A2( u0_u13_u1_n170 ) );
  AOI211_X1 u0_u13_u1_U5 (.ZN( u0_u13_u1_n124 ) , .A( u0_u13_u1_n138 ) , .C2( u0_u13_u1_n139 ) , .B( u0_u13_u1_n145 ) , .C1( u0_u13_u1_n147 ) );
  NAND2_X1 u0_u13_u1_U50 (.ZN( u0_u13_u1_n129 ) , .A2( u0_u13_u1_n95 ) , .A1( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U51 (.A1( u0_u13_u1_n102 ) , .ZN( u0_u13_u1_n154 ) , .A2( u0_u13_u1_n99 ) );
  NAND2_X1 u0_u13_u1_U52 (.A2( u0_u13_u1_n100 ) , .ZN( u0_u13_u1_n135 ) , .A1( u0_u13_u1_n99 ) );
  AOI21_X1 u0_u13_u1_U53 (.A( u0_u13_u1_n152 ) , .B2( u0_u13_u1_n153 ) , .B1( u0_u13_u1_n154 ) , .ZN( u0_u13_u1_n158 ) );
  INV_X1 u0_u13_u1_U54 (.A( u0_u13_u1_n160 ) , .ZN( u0_u13_u1_n175 ) );
  NAND2_X1 u0_u13_u1_U55 (.A1( u0_u13_u1_n100 ) , .ZN( u0_u13_u1_n116 ) , .A2( u0_u13_u1_n95 ) );
  NAND2_X1 u0_u13_u1_U56 (.A1( u0_u13_u1_n102 ) , .ZN( u0_u13_u1_n131 ) , .A2( u0_u13_u1_n95 ) );
  NAND2_X1 u0_u13_u1_U57 (.A2( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n121 ) , .A1( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U58 (.A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n153 ) , .A2( u0_u13_u1_n98 ) );
  NAND2_X1 u0_u13_u1_U59 (.A2( u0_u13_u1_n104 ) , .A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n133 ) );
  AOI22_X1 u0_u13_u1_U6 (.B2( u0_u13_u1_n136 ) , .A2( u0_u13_u1_n137 ) , .ZN( u0_u13_u1_n143 ) , .A1( u0_u13_u1_n171 ) , .B1( u0_u13_u1_n173 ) );
  NAND2_X1 u0_u13_u1_U60 (.ZN( u0_u13_u1_n150 ) , .A2( u0_u13_u1_n98 ) , .A1( u0_u13_u1_n99 ) );
  NAND2_X1 u0_u13_u1_U61 (.A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n155 ) , .A2( u0_u13_u1_n95 ) );
  OAI21_X1 u0_u13_u1_U62 (.ZN( u0_u13_u1_n109 ) , .B1( u0_u13_u1_n129 ) , .B2( u0_u13_u1_n160 ) , .A( u0_u13_u1_n167 ) );
  NAND2_X1 u0_u13_u1_U63 (.A2( u0_u13_u1_n100 ) , .A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n120 ) );
  NAND2_X1 u0_u13_u1_U64 (.A1( u0_u13_u1_n102 ) , .A2( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n115 ) );
  NAND2_X1 u0_u13_u1_U65 (.A2( u0_u13_u1_n100 ) , .A1( u0_u13_u1_n104 ) , .ZN( u0_u13_u1_n151 ) );
  NAND2_X1 u0_u13_u1_U66 (.A2( u0_u13_u1_n103 ) , .A1( u0_u13_u1_n105 ) , .ZN( u0_u13_u1_n161 ) );
  INV_X1 u0_u13_u1_U67 (.A( u0_u13_u1_n152 ) , .ZN( u0_u13_u1_n173 ) );
  INV_X1 u0_u13_u1_U68 (.A( u0_u13_u1_n128 ) , .ZN( u0_u13_u1_n172 ) );
  NAND2_X1 u0_u13_u1_U69 (.A2( u0_u13_u1_n102 ) , .A1( u0_u13_u1_n103 ) , .ZN( u0_u13_u1_n123 ) );
  INV_X1 u0_u13_u1_U7 (.A( u0_u13_u1_n147 ) , .ZN( u0_u13_u1_n181 ) );
  NOR2_X1 u0_u13_u1_U70 (.A2( u0_u13_X_7 ) , .A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n95 ) );
  NOR2_X1 u0_u13_u1_U71 (.A1( u0_u13_X_12 ) , .A2( u0_u13_X_9 ) , .ZN( u0_u13_u1_n100 ) );
  NOR2_X1 u0_u13_u1_U72 (.A2( u0_u13_X_8 ) , .A1( u0_u13_u1_n177 ) , .ZN( u0_u13_u1_n99 ) );
  NOR2_X1 u0_u13_u1_U73 (.A2( u0_u13_X_12 ) , .ZN( u0_u13_u1_n102 ) , .A1( u0_u13_u1_n176 ) );
  NOR2_X1 u0_u13_u1_U74 (.A2( u0_u13_X_9 ) , .ZN( u0_u13_u1_n105 ) , .A1( u0_u13_u1_n168 ) );
  NAND2_X1 u0_u13_u1_U75 (.A1( u0_u13_X_10 ) , .ZN( u0_u13_u1_n160 ) , .A2( u0_u13_u1_n169 ) );
  NAND2_X1 u0_u13_u1_U76 (.A2( u0_u13_X_10 ) , .A1( u0_u13_X_11 ) , .ZN( u0_u13_u1_n152 ) );
  NAND2_X1 u0_u13_u1_U77 (.A1( u0_u13_X_11 ) , .ZN( u0_u13_u1_n128 ) , .A2( u0_u13_u1_n170 ) );
  AND2_X1 u0_u13_u1_U78 (.A2( u0_u13_X_7 ) , .A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n104 ) );
  AND2_X1 u0_u13_u1_U79 (.A1( u0_u13_X_8 ) , .ZN( u0_u13_u1_n103 ) , .A2( u0_u13_u1_n177 ) );
  NOR2_X1 u0_u13_u1_U8 (.A1( u0_u13_u1_n112 ) , .A2( u0_u13_u1_n116 ) , .ZN( u0_u13_u1_n118 ) );
  INV_X1 u0_u13_u1_U80 (.A( u0_u13_X_10 ) , .ZN( u0_u13_u1_n170 ) );
  INV_X1 u0_u13_u1_U81 (.A( u0_u13_X_9 ) , .ZN( u0_u13_u1_n176 ) );
  INV_X1 u0_u13_u1_U82 (.A( u0_u13_X_11 ) , .ZN( u0_u13_u1_n169 ) );
  INV_X1 u0_u13_u1_U83 (.A( u0_u13_X_12 ) , .ZN( u0_u13_u1_n168 ) );
  INV_X1 u0_u13_u1_U84 (.A( u0_u13_X_7 ) , .ZN( u0_u13_u1_n177 ) );
  NAND4_X1 u0_u13_u1_U85 (.ZN( u0_out13_28 ) , .A4( u0_u13_u1_n124 ) , .A3( u0_u13_u1_n125 ) , .A2( u0_u13_u1_n126 ) , .A1( u0_u13_u1_n127 ) );
  OAI21_X1 u0_u13_u1_U86 (.ZN( u0_u13_u1_n127 ) , .B2( u0_u13_u1_n139 ) , .B1( u0_u13_u1_n175 ) , .A( u0_u13_u1_n183 ) );
  OAI21_X1 u0_u13_u1_U87 (.ZN( u0_u13_u1_n126 ) , .B2( u0_u13_u1_n140 ) , .A( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n178 ) );
  NAND4_X1 u0_u13_u1_U88 (.ZN( u0_out13_18 ) , .A4( u0_u13_u1_n165 ) , .A3( u0_u13_u1_n166 ) , .A1( u0_u13_u1_n167 ) , .A2( u0_u13_u1_n186 ) );
  AOI22_X1 u0_u13_u1_U89 (.B2( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n147 ) , .A2( u0_u13_u1_n148 ) , .ZN( u0_u13_u1_n166 ) , .A1( u0_u13_u1_n172 ) );
  OAI21_X1 u0_u13_u1_U9 (.ZN( u0_u13_u1_n101 ) , .B1( u0_u13_u1_n141 ) , .A( u0_u13_u1_n146 ) , .B2( u0_u13_u1_n183 ) );
  INV_X1 u0_u13_u1_U90 (.A( u0_u13_u1_n145 ) , .ZN( u0_u13_u1_n186 ) );
  NAND4_X1 u0_u13_u1_U91 (.ZN( u0_out13_2 ) , .A4( u0_u13_u1_n142 ) , .A3( u0_u13_u1_n143 ) , .A2( u0_u13_u1_n144 ) , .A1( u0_u13_u1_n179 ) );
  OAI21_X1 u0_u13_u1_U92 (.B2( u0_u13_u1_n132 ) , .ZN( u0_u13_u1_n144 ) , .A( u0_u13_u1_n146 ) , .B1( u0_u13_u1_n180 ) );
  INV_X1 u0_u13_u1_U93 (.A( u0_u13_u1_n130 ) , .ZN( u0_u13_u1_n179 ) );
  OR4_X1 u0_u13_u1_U94 (.ZN( u0_out13_13 ) , .A4( u0_u13_u1_n108 ) , .A3( u0_u13_u1_n109 ) , .A2( u0_u13_u1_n110 ) , .A1( u0_u13_u1_n111 ) );
  AOI21_X1 u0_u13_u1_U95 (.ZN( u0_u13_u1_n111 ) , .A( u0_u13_u1_n128 ) , .B2( u0_u13_u1_n131 ) , .B1( u0_u13_u1_n135 ) );
  AOI21_X1 u0_u13_u1_U96 (.ZN( u0_u13_u1_n110 ) , .A( u0_u13_u1_n116 ) , .B1( u0_u13_u1_n152 ) , .B2( u0_u13_u1_n160 ) );
  NAND3_X1 u0_u13_u1_U97 (.A3( u0_u13_u1_n149 ) , .A2( u0_u13_u1_n150 ) , .A1( u0_u13_u1_n151 ) , .ZN( u0_u13_u1_n164 ) );
  NAND3_X1 u0_u13_u1_U98 (.A3( u0_u13_u1_n134 ) , .A2( u0_u13_u1_n135 ) , .ZN( u0_u13_u1_n136 ) , .A1( u0_u13_u1_n151 ) );
  NAND3_X1 u0_u13_u1_U99 (.A1( u0_u13_u1_n133 ) , .ZN( u0_u13_u1_n137 ) , .A2( u0_u13_u1_n154 ) , .A3( u0_u13_u1_n181 ) );
  OAI22_X1 u0_u13_u2_U10 (.B1( u0_u13_u2_n151 ) , .A2( u0_u13_u2_n152 ) , .A1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n160 ) , .B2( u0_u13_u2_n168 ) );
  NAND3_X1 u0_u13_u2_U100 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n98 ) );
  NOR3_X1 u0_u13_u2_U11 (.A1( u0_u13_u2_n150 ) , .ZN( u0_u13_u2_n151 ) , .A3( u0_u13_u2_n175 ) , .A2( u0_u13_u2_n188 ) );
  AOI21_X1 u0_u13_u2_U12 (.B2( u0_u13_u2_n123 ) , .ZN( u0_u13_u2_n125 ) , .A( u0_u13_u2_n171 ) , .B1( u0_u13_u2_n184 ) );
  INV_X1 u0_u13_u2_U13 (.A( u0_u13_u2_n150 ) , .ZN( u0_u13_u2_n184 ) );
  AOI21_X1 u0_u13_u2_U14 (.ZN( u0_u13_u2_n144 ) , .B2( u0_u13_u2_n155 ) , .A( u0_u13_u2_n172 ) , .B1( u0_u13_u2_n185 ) );
  AOI21_X1 u0_u13_u2_U15 (.B2( u0_u13_u2_n143 ) , .ZN( u0_u13_u2_n145 ) , .B1( u0_u13_u2_n152 ) , .A( u0_u13_u2_n171 ) );
  INV_X1 u0_u13_u2_U16 (.A( u0_u13_u2_n156 ) , .ZN( u0_u13_u2_n171 ) );
  INV_X1 u0_u13_u2_U17 (.A( u0_u13_u2_n120 ) , .ZN( u0_u13_u2_n188 ) );
  NAND2_X1 u0_u13_u2_U18 (.A2( u0_u13_u2_n122 ) , .ZN( u0_u13_u2_n150 ) , .A1( u0_u13_u2_n152 ) );
  INV_X1 u0_u13_u2_U19 (.A( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n170 ) );
  INV_X1 u0_u13_u2_U20 (.A( u0_u13_u2_n137 ) , .ZN( u0_u13_u2_n173 ) );
  NAND2_X1 u0_u13_u2_U21 (.A1( u0_u13_u2_n132 ) , .A2( u0_u13_u2_n139 ) , .ZN( u0_u13_u2_n157 ) );
  INV_X1 u0_u13_u2_U22 (.A( u0_u13_u2_n113 ) , .ZN( u0_u13_u2_n178 ) );
  INV_X1 u0_u13_u2_U23 (.A( u0_u13_u2_n139 ) , .ZN( u0_u13_u2_n175 ) );
  INV_X1 u0_u13_u2_U24 (.A( u0_u13_u2_n155 ) , .ZN( u0_u13_u2_n181 ) );
  INV_X1 u0_u13_u2_U25 (.A( u0_u13_u2_n119 ) , .ZN( u0_u13_u2_n177 ) );
  INV_X1 u0_u13_u2_U26 (.A( u0_u13_u2_n116 ) , .ZN( u0_u13_u2_n180 ) );
  INV_X1 u0_u13_u2_U27 (.A( u0_u13_u2_n131 ) , .ZN( u0_u13_u2_n179 ) );
  INV_X1 u0_u13_u2_U28 (.A( u0_u13_u2_n154 ) , .ZN( u0_u13_u2_n176 ) );
  NAND2_X1 u0_u13_u2_U29 (.A2( u0_u13_u2_n116 ) , .A1( u0_u13_u2_n117 ) , .ZN( u0_u13_u2_n118 ) );
  NOR2_X1 u0_u13_u2_U3 (.ZN( u0_u13_u2_n121 ) , .A2( u0_u13_u2_n177 ) , .A1( u0_u13_u2_n180 ) );
  INV_X1 u0_u13_u2_U30 (.A( u0_u13_u2_n132 ) , .ZN( u0_u13_u2_n182 ) );
  INV_X1 u0_u13_u2_U31 (.A( u0_u13_u2_n158 ) , .ZN( u0_u13_u2_n183 ) );
  OAI21_X1 u0_u13_u2_U32 (.A( u0_u13_u2_n156 ) , .B1( u0_u13_u2_n157 ) , .ZN( u0_u13_u2_n158 ) , .B2( u0_u13_u2_n179 ) );
  NOR2_X1 u0_u13_u2_U33 (.ZN( u0_u13_u2_n156 ) , .A1( u0_u13_u2_n166 ) , .A2( u0_u13_u2_n169 ) );
  NOR2_X1 u0_u13_u2_U34 (.A2( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n137 ) , .A1( u0_u13_u2_n140 ) );
  NOR2_X1 u0_u13_u2_U35 (.A2( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n153 ) , .A1( u0_u13_u2_n156 ) );
  AOI211_X1 u0_u13_u2_U36 (.ZN( u0_u13_u2_n130 ) , .C1( u0_u13_u2_n138 ) , .C2( u0_u13_u2_n179 ) , .B( u0_u13_u2_n96 ) , .A( u0_u13_u2_n97 ) );
  OAI22_X1 u0_u13_u2_U37 (.B1( u0_u13_u2_n133 ) , .A2( u0_u13_u2_n137 ) , .A1( u0_u13_u2_n152 ) , .B2( u0_u13_u2_n168 ) , .ZN( u0_u13_u2_n97 ) );
  OAI221_X1 u0_u13_u2_U38 (.B1( u0_u13_u2_n113 ) , .C1( u0_u13_u2_n132 ) , .A( u0_u13_u2_n149 ) , .B2( u0_u13_u2_n171 ) , .C2( u0_u13_u2_n172 ) , .ZN( u0_u13_u2_n96 ) );
  OAI221_X1 u0_u13_u2_U39 (.A( u0_u13_u2_n115 ) , .C2( u0_u13_u2_n123 ) , .B2( u0_u13_u2_n143 ) , .B1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n163 ) , .C1( u0_u13_u2_n168 ) );
  INV_X1 u0_u13_u2_U4 (.A( u0_u13_u2_n134 ) , .ZN( u0_u13_u2_n185 ) );
  OAI21_X1 u0_u13_u2_U40 (.A( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n115 ) , .B1( u0_u13_u2_n176 ) , .B2( u0_u13_u2_n178 ) );
  OAI221_X1 u0_u13_u2_U41 (.A( u0_u13_u2_n135 ) , .B2( u0_u13_u2_n136 ) , .B1( u0_u13_u2_n137 ) , .ZN( u0_u13_u2_n162 ) , .C2( u0_u13_u2_n167 ) , .C1( u0_u13_u2_n185 ) );
  AND3_X1 u0_u13_u2_U42 (.A3( u0_u13_u2_n131 ) , .A2( u0_u13_u2_n132 ) , .A1( u0_u13_u2_n133 ) , .ZN( u0_u13_u2_n136 ) );
  AOI22_X1 u0_u13_u2_U43 (.ZN( u0_u13_u2_n135 ) , .B1( u0_u13_u2_n140 ) , .A1( u0_u13_u2_n156 ) , .B2( u0_u13_u2_n180 ) , .A2( u0_u13_u2_n188 ) );
  AOI21_X1 u0_u13_u2_U44 (.ZN( u0_u13_u2_n149 ) , .B1( u0_u13_u2_n173 ) , .B2( u0_u13_u2_n188 ) , .A( u0_u13_u2_n95 ) );
  AND3_X1 u0_u13_u2_U45 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n156 ) , .ZN( u0_u13_u2_n95 ) );
  OAI21_X1 u0_u13_u2_U46 (.A( u0_u13_u2_n141 ) , .B2( u0_u13_u2_n142 ) , .ZN( u0_u13_u2_n146 ) , .B1( u0_u13_u2_n153 ) );
  OAI21_X1 u0_u13_u2_U47 (.A( u0_u13_u2_n140 ) , .ZN( u0_u13_u2_n141 ) , .B1( u0_u13_u2_n176 ) , .B2( u0_u13_u2_n177 ) );
  NOR3_X1 u0_u13_u2_U48 (.ZN( u0_u13_u2_n142 ) , .A3( u0_u13_u2_n175 ) , .A2( u0_u13_u2_n178 ) , .A1( u0_u13_u2_n181 ) );
  OAI21_X1 u0_u13_u2_U49 (.A( u0_u13_u2_n101 ) , .B2( u0_u13_u2_n121 ) , .B1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n164 ) );
  NOR4_X1 u0_u13_u2_U5 (.A4( u0_u13_u2_n124 ) , .A3( u0_u13_u2_n125 ) , .A2( u0_u13_u2_n126 ) , .A1( u0_u13_u2_n127 ) , .ZN( u0_u13_u2_n128 ) );
  NAND2_X1 u0_u13_u2_U50 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n155 ) );
  NAND2_X1 u0_u13_u2_U51 (.A2( u0_u13_u2_n105 ) , .A1( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n143 ) );
  NAND2_X1 u0_u13_u2_U52 (.A1( u0_u13_u2_n104 ) , .A2( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n152 ) );
  NAND2_X1 u0_u13_u2_U53 (.A1( u0_u13_u2_n100 ) , .A2( u0_u13_u2_n105 ) , .ZN( u0_u13_u2_n132 ) );
  INV_X1 u0_u13_u2_U54 (.A( u0_u13_u2_n140 ) , .ZN( u0_u13_u2_n168 ) );
  INV_X1 u0_u13_u2_U55 (.A( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n167 ) );
  NAND2_X1 u0_u13_u2_U56 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n113 ) );
  NAND2_X1 u0_u13_u2_U57 (.A1( u0_u13_u2_n106 ) , .A2( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n131 ) );
  NAND2_X1 u0_u13_u2_U58 (.A1( u0_u13_u2_n103 ) , .A2( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n139 ) );
  NAND2_X1 u0_u13_u2_U59 (.A1( u0_u13_u2_n103 ) , .A2( u0_u13_u2_n105 ) , .ZN( u0_u13_u2_n133 ) );
  AOI21_X1 u0_u13_u2_U6 (.B2( u0_u13_u2_n119 ) , .ZN( u0_u13_u2_n127 ) , .A( u0_u13_u2_n137 ) , .B1( u0_u13_u2_n155 ) );
  NAND2_X1 u0_u13_u2_U60 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n103 ) , .ZN( u0_u13_u2_n154 ) );
  NAND2_X1 u0_u13_u2_U61 (.A2( u0_u13_u2_n103 ) , .A1( u0_u13_u2_n104 ) , .ZN( u0_u13_u2_n119 ) );
  NAND2_X1 u0_u13_u2_U62 (.A2( u0_u13_u2_n107 ) , .A1( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n123 ) );
  NAND2_X1 u0_u13_u2_U63 (.A1( u0_u13_u2_n104 ) , .A2( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n122 ) );
  INV_X1 u0_u13_u2_U64 (.A( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n172 ) );
  NAND2_X1 u0_u13_u2_U65 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n102 ) , .ZN( u0_u13_u2_n116 ) );
  NAND2_X1 u0_u13_u2_U66 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n120 ) );
  NAND2_X1 u0_u13_u2_U67 (.A2( u0_u13_u2_n105 ) , .A1( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n117 ) );
  INV_X1 u0_u13_u2_U68 (.ZN( u0_u13_u2_n187 ) , .A( u0_u13_u2_n99 ) );
  OAI21_X1 u0_u13_u2_U69 (.B1( u0_u13_u2_n137 ) , .B2( u0_u13_u2_n143 ) , .A( u0_u13_u2_n98 ) , .ZN( u0_u13_u2_n99 ) );
  AOI21_X1 u0_u13_u2_U7 (.ZN( u0_u13_u2_n124 ) , .B1( u0_u13_u2_n131 ) , .B2( u0_u13_u2_n143 ) , .A( u0_u13_u2_n172 ) );
  NOR2_X1 u0_u13_u2_U70 (.A2( u0_u13_X_16 ) , .ZN( u0_u13_u2_n140 ) , .A1( u0_u13_u2_n166 ) );
  NOR2_X1 u0_u13_u2_U71 (.A2( u0_u13_X_13 ) , .A1( u0_u13_X_14 ) , .ZN( u0_u13_u2_n100 ) );
  NOR2_X1 u0_u13_u2_U72 (.A2( u0_u13_X_16 ) , .A1( u0_u13_X_17 ) , .ZN( u0_u13_u2_n138 ) );
  NOR2_X1 u0_u13_u2_U73 (.A2( u0_u13_X_15 ) , .A1( u0_u13_X_18 ) , .ZN( u0_u13_u2_n104 ) );
  NOR2_X1 u0_u13_u2_U74 (.A2( u0_u13_X_14 ) , .ZN( u0_u13_u2_n103 ) , .A1( u0_u13_u2_n174 ) );
  NOR2_X1 u0_u13_u2_U75 (.A2( u0_u13_X_15 ) , .ZN( u0_u13_u2_n102 ) , .A1( u0_u13_u2_n165 ) );
  NOR2_X1 u0_u13_u2_U76 (.A2( u0_u13_X_17 ) , .ZN( u0_u13_u2_n114 ) , .A1( u0_u13_u2_n169 ) );
  AND2_X1 u0_u13_u2_U77 (.A1( u0_u13_X_15 ) , .ZN( u0_u13_u2_n105 ) , .A2( u0_u13_u2_n165 ) );
  AND2_X1 u0_u13_u2_U78 (.A2( u0_u13_X_15 ) , .A1( u0_u13_X_18 ) , .ZN( u0_u13_u2_n107 ) );
  AND2_X1 u0_u13_u2_U79 (.A1( u0_u13_X_14 ) , .ZN( u0_u13_u2_n106 ) , .A2( u0_u13_u2_n174 ) );
  AOI21_X1 u0_u13_u2_U8 (.B2( u0_u13_u2_n120 ) , .B1( u0_u13_u2_n121 ) , .ZN( u0_u13_u2_n126 ) , .A( u0_u13_u2_n167 ) );
  AND2_X1 u0_u13_u2_U80 (.A1( u0_u13_X_13 ) , .A2( u0_u13_X_14 ) , .ZN( u0_u13_u2_n108 ) );
  INV_X1 u0_u13_u2_U81 (.A( u0_u13_X_16 ) , .ZN( u0_u13_u2_n169 ) );
  INV_X1 u0_u13_u2_U82 (.A( u0_u13_X_17 ) , .ZN( u0_u13_u2_n166 ) );
  INV_X1 u0_u13_u2_U83 (.A( u0_u13_X_13 ) , .ZN( u0_u13_u2_n174 ) );
  INV_X1 u0_u13_u2_U84 (.A( u0_u13_X_18 ) , .ZN( u0_u13_u2_n165 ) );
  NAND4_X1 u0_u13_u2_U85 (.ZN( u0_out13_30 ) , .A4( u0_u13_u2_n147 ) , .A3( u0_u13_u2_n148 ) , .A2( u0_u13_u2_n149 ) , .A1( u0_u13_u2_n187 ) );
  NOR3_X1 u0_u13_u2_U86 (.A3( u0_u13_u2_n144 ) , .A2( u0_u13_u2_n145 ) , .A1( u0_u13_u2_n146 ) , .ZN( u0_u13_u2_n147 ) );
  AOI21_X1 u0_u13_u2_U87 (.B2( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n148 ) , .A( u0_u13_u2_n162 ) , .B1( u0_u13_u2_n182 ) );
  NAND4_X1 u0_u13_u2_U88 (.ZN( u0_out13_24 ) , .A4( u0_u13_u2_n111 ) , .A3( u0_u13_u2_n112 ) , .A1( u0_u13_u2_n130 ) , .A2( u0_u13_u2_n187 ) );
  AOI221_X1 u0_u13_u2_U89 (.A( u0_u13_u2_n109 ) , .B1( u0_u13_u2_n110 ) , .ZN( u0_u13_u2_n111 ) , .C1( u0_u13_u2_n134 ) , .C2( u0_u13_u2_n170 ) , .B2( u0_u13_u2_n173 ) );
  OAI22_X1 u0_u13_u2_U9 (.ZN( u0_u13_u2_n109 ) , .A2( u0_u13_u2_n113 ) , .B2( u0_u13_u2_n133 ) , .B1( u0_u13_u2_n167 ) , .A1( u0_u13_u2_n168 ) );
  AOI21_X1 u0_u13_u2_U90 (.ZN( u0_u13_u2_n112 ) , .B2( u0_u13_u2_n156 ) , .A( u0_u13_u2_n164 ) , .B1( u0_u13_u2_n181 ) );
  NAND4_X1 u0_u13_u2_U91 (.ZN( u0_out13_16 ) , .A4( u0_u13_u2_n128 ) , .A3( u0_u13_u2_n129 ) , .A1( u0_u13_u2_n130 ) , .A2( u0_u13_u2_n186 ) );
  AOI22_X1 u0_u13_u2_U92 (.A2( u0_u13_u2_n118 ) , .ZN( u0_u13_u2_n129 ) , .A1( u0_u13_u2_n140 ) , .B1( u0_u13_u2_n157 ) , .B2( u0_u13_u2_n170 ) );
  INV_X1 u0_u13_u2_U93 (.A( u0_u13_u2_n163 ) , .ZN( u0_u13_u2_n186 ) );
  OR4_X1 u0_u13_u2_U94 (.ZN( u0_out13_6 ) , .A4( u0_u13_u2_n161 ) , .A3( u0_u13_u2_n162 ) , .A2( u0_u13_u2_n163 ) , .A1( u0_u13_u2_n164 ) );
  OR3_X1 u0_u13_u2_U95 (.A2( u0_u13_u2_n159 ) , .A1( u0_u13_u2_n160 ) , .ZN( u0_u13_u2_n161 ) , .A3( u0_u13_u2_n183 ) );
  AOI21_X1 u0_u13_u2_U96 (.B2( u0_u13_u2_n154 ) , .B1( u0_u13_u2_n155 ) , .ZN( u0_u13_u2_n159 ) , .A( u0_u13_u2_n167 ) );
  NAND3_X1 u0_u13_u2_U97 (.A2( u0_u13_u2_n117 ) , .A1( u0_u13_u2_n122 ) , .A3( u0_u13_u2_n123 ) , .ZN( u0_u13_u2_n134 ) );
  NAND3_X1 u0_u13_u2_U98 (.ZN( u0_u13_u2_n110 ) , .A2( u0_u13_u2_n131 ) , .A3( u0_u13_u2_n139 ) , .A1( u0_u13_u2_n154 ) );
  NAND3_X1 u0_u13_u2_U99 (.A2( u0_u13_u2_n100 ) , .ZN( u0_u13_u2_n101 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n114 ) );
  OAI22_X1 u0_u13_u3_U10 (.B1( u0_u13_u3_n113 ) , .A2( u0_u13_u3_n135 ) , .A1( u0_u13_u3_n150 ) , .B2( u0_u13_u3_n164 ) , .ZN( u0_u13_u3_n98 ) );
  OAI211_X1 u0_u13_u3_U11 (.B( u0_u13_u3_n106 ) , .ZN( u0_u13_u3_n119 ) , .C2( u0_u13_u3_n128 ) , .C1( u0_u13_u3_n167 ) , .A( u0_u13_u3_n181 ) );
  AOI221_X1 u0_u13_u3_U12 (.C1( u0_u13_u3_n105 ) , .ZN( u0_u13_u3_n106 ) , .A( u0_u13_u3_n131 ) , .B2( u0_u13_u3_n132 ) , .C2( u0_u13_u3_n133 ) , .B1( u0_u13_u3_n169 ) );
  INV_X1 u0_u13_u3_U13 (.ZN( u0_u13_u3_n181 ) , .A( u0_u13_u3_n98 ) );
  NAND2_X1 u0_u13_u3_U14 (.ZN( u0_u13_u3_n105 ) , .A2( u0_u13_u3_n130 ) , .A1( u0_u13_u3_n155 ) );
  AOI22_X1 u0_u13_u3_U15 (.B1( u0_u13_u3_n115 ) , .A2( u0_u13_u3_n116 ) , .ZN( u0_u13_u3_n123 ) , .B2( u0_u13_u3_n133 ) , .A1( u0_u13_u3_n169 ) );
  NAND2_X1 u0_u13_u3_U16 (.ZN( u0_u13_u3_n116 ) , .A2( u0_u13_u3_n151 ) , .A1( u0_u13_u3_n182 ) );
  NOR2_X1 u0_u13_u3_U17 (.ZN( u0_u13_u3_n126 ) , .A2( u0_u13_u3_n150 ) , .A1( u0_u13_u3_n164 ) );
  AOI21_X1 u0_u13_u3_U18 (.ZN( u0_u13_u3_n112 ) , .B2( u0_u13_u3_n146 ) , .B1( u0_u13_u3_n155 ) , .A( u0_u13_u3_n167 ) );
  NAND2_X1 u0_u13_u3_U19 (.A1( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n142 ) , .A2( u0_u13_u3_n164 ) );
  NAND2_X1 u0_u13_u3_U20 (.ZN( u0_u13_u3_n132 ) , .A2( u0_u13_u3_n152 ) , .A1( u0_u13_u3_n156 ) );
  AND2_X1 u0_u13_u3_U21 (.A2( u0_u13_u3_n113 ) , .A1( u0_u13_u3_n114 ) , .ZN( u0_u13_u3_n151 ) );
  INV_X1 u0_u13_u3_U22 (.A( u0_u13_u3_n133 ) , .ZN( u0_u13_u3_n165 ) );
  INV_X1 u0_u13_u3_U23 (.A( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n170 ) );
  NAND2_X1 u0_u13_u3_U24 (.A1( u0_u13_u3_n107 ) , .A2( u0_u13_u3_n108 ) , .ZN( u0_u13_u3_n140 ) );
  NAND2_X1 u0_u13_u3_U25 (.ZN( u0_u13_u3_n117 ) , .A1( u0_u13_u3_n124 ) , .A2( u0_u13_u3_n148 ) );
  NAND2_X1 u0_u13_u3_U26 (.ZN( u0_u13_u3_n143 ) , .A1( u0_u13_u3_n165 ) , .A2( u0_u13_u3_n167 ) );
  INV_X1 u0_u13_u3_U27 (.A( u0_u13_u3_n130 ) , .ZN( u0_u13_u3_n177 ) );
  INV_X1 u0_u13_u3_U28 (.A( u0_u13_u3_n128 ) , .ZN( u0_u13_u3_n176 ) );
  INV_X1 u0_u13_u3_U29 (.A( u0_u13_u3_n155 ) , .ZN( u0_u13_u3_n174 ) );
  INV_X1 u0_u13_u3_U3 (.A( u0_u13_u3_n129 ) , .ZN( u0_u13_u3_n183 ) );
  INV_X1 u0_u13_u3_U30 (.A( u0_u13_u3_n139 ) , .ZN( u0_u13_u3_n185 ) );
  NOR2_X1 u0_u13_u3_U31 (.ZN( u0_u13_u3_n135 ) , .A2( u0_u13_u3_n141 ) , .A1( u0_u13_u3_n169 ) );
  OAI222_X1 u0_u13_u3_U32 (.C2( u0_u13_u3_n107 ) , .A2( u0_u13_u3_n108 ) , .B1( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n138 ) , .B2( u0_u13_u3_n146 ) , .C1( u0_u13_u3_n154 ) , .A1( u0_u13_u3_n164 ) );
  NOR4_X1 u0_u13_u3_U33 (.A4( u0_u13_u3_n157 ) , .A3( u0_u13_u3_n158 ) , .A2( u0_u13_u3_n159 ) , .A1( u0_u13_u3_n160 ) , .ZN( u0_u13_u3_n161 ) );
  AOI21_X1 u0_u13_u3_U34 (.B2( u0_u13_u3_n152 ) , .B1( u0_u13_u3_n153 ) , .ZN( u0_u13_u3_n158 ) , .A( u0_u13_u3_n164 ) );
  AOI21_X1 u0_u13_u3_U35 (.A( u0_u13_u3_n154 ) , .B2( u0_u13_u3_n155 ) , .B1( u0_u13_u3_n156 ) , .ZN( u0_u13_u3_n157 ) );
  AOI21_X1 u0_u13_u3_U36 (.A( u0_u13_u3_n149 ) , .B2( u0_u13_u3_n150 ) , .B1( u0_u13_u3_n151 ) , .ZN( u0_u13_u3_n159 ) );
  AOI211_X1 u0_u13_u3_U37 (.ZN( u0_u13_u3_n109 ) , .A( u0_u13_u3_n119 ) , .C2( u0_u13_u3_n129 ) , .B( u0_u13_u3_n138 ) , .C1( u0_u13_u3_n141 ) );
  AOI211_X1 u0_u13_u3_U38 (.B( u0_u13_u3_n119 ) , .A( u0_u13_u3_n120 ) , .C2( u0_u13_u3_n121 ) , .ZN( u0_u13_u3_n122 ) , .C1( u0_u13_u3_n179 ) );
  INV_X1 u0_u13_u3_U39 (.A( u0_u13_u3_n156 ) , .ZN( u0_u13_u3_n179 ) );
  INV_X1 u0_u13_u3_U4 (.A( u0_u13_u3_n140 ) , .ZN( u0_u13_u3_n182 ) );
  OAI22_X1 u0_u13_u3_U40 (.B1( u0_u13_u3_n118 ) , .ZN( u0_u13_u3_n120 ) , .A1( u0_u13_u3_n135 ) , .B2( u0_u13_u3_n154 ) , .A2( u0_u13_u3_n178 ) );
  AND3_X1 u0_u13_u3_U41 (.ZN( u0_u13_u3_n118 ) , .A2( u0_u13_u3_n124 ) , .A1( u0_u13_u3_n144 ) , .A3( u0_u13_u3_n152 ) );
  INV_X1 u0_u13_u3_U42 (.A( u0_u13_u3_n121 ) , .ZN( u0_u13_u3_n164 ) );
  NAND2_X1 u0_u13_u3_U43 (.ZN( u0_u13_u3_n133 ) , .A1( u0_u13_u3_n154 ) , .A2( u0_u13_u3_n164 ) );
  OAI211_X1 u0_u13_u3_U44 (.B( u0_u13_u3_n127 ) , .ZN( u0_u13_u3_n139 ) , .C1( u0_u13_u3_n150 ) , .C2( u0_u13_u3_n154 ) , .A( u0_u13_u3_n184 ) );
  INV_X1 u0_u13_u3_U45 (.A( u0_u13_u3_n125 ) , .ZN( u0_u13_u3_n184 ) );
  AOI221_X1 u0_u13_u3_U46 (.A( u0_u13_u3_n126 ) , .ZN( u0_u13_u3_n127 ) , .C2( u0_u13_u3_n132 ) , .C1( u0_u13_u3_n169 ) , .B2( u0_u13_u3_n170 ) , .B1( u0_u13_u3_n174 ) );
  OAI22_X1 u0_u13_u3_U47 (.A1( u0_u13_u3_n124 ) , .ZN( u0_u13_u3_n125 ) , .B2( u0_u13_u3_n145 ) , .A2( u0_u13_u3_n165 ) , .B1( u0_u13_u3_n167 ) );
  NOR2_X1 u0_u13_u3_U48 (.A1( u0_u13_u3_n113 ) , .ZN( u0_u13_u3_n131 ) , .A2( u0_u13_u3_n154 ) );
  NAND2_X1 u0_u13_u3_U49 (.A1( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n150 ) , .A2( u0_u13_u3_n99 ) );
  INV_X1 u0_u13_u3_U5 (.A( u0_u13_u3_n117 ) , .ZN( u0_u13_u3_n178 ) );
  NAND2_X1 u0_u13_u3_U50 (.A2( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n155 ) , .A1( u0_u13_u3_n97 ) );
  INV_X1 u0_u13_u3_U51 (.A( u0_u13_u3_n141 ) , .ZN( u0_u13_u3_n167 ) );
  AOI21_X1 u0_u13_u3_U52 (.B2( u0_u13_u3_n114 ) , .B1( u0_u13_u3_n146 ) , .A( u0_u13_u3_n154 ) , .ZN( u0_u13_u3_n94 ) );
  AOI21_X1 u0_u13_u3_U53 (.ZN( u0_u13_u3_n110 ) , .B2( u0_u13_u3_n142 ) , .B1( u0_u13_u3_n186 ) , .A( u0_u13_u3_n95 ) );
  INV_X1 u0_u13_u3_U54 (.A( u0_u13_u3_n145 ) , .ZN( u0_u13_u3_n186 ) );
  AOI21_X1 u0_u13_u3_U55 (.B1( u0_u13_u3_n124 ) , .A( u0_u13_u3_n149 ) , .B2( u0_u13_u3_n155 ) , .ZN( u0_u13_u3_n95 ) );
  INV_X1 u0_u13_u3_U56 (.A( u0_u13_u3_n149 ) , .ZN( u0_u13_u3_n169 ) );
  NAND2_X1 u0_u13_u3_U57 (.ZN( u0_u13_u3_n124 ) , .A1( u0_u13_u3_n96 ) , .A2( u0_u13_u3_n97 ) );
  NAND2_X1 u0_u13_u3_U58 (.A2( u0_u13_u3_n100 ) , .ZN( u0_u13_u3_n146 ) , .A1( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U59 (.A1( u0_u13_u3_n101 ) , .ZN( u0_u13_u3_n145 ) , .A2( u0_u13_u3_n99 ) );
  AOI221_X1 u0_u13_u3_U6 (.A( u0_u13_u3_n131 ) , .C2( u0_u13_u3_n132 ) , .C1( u0_u13_u3_n133 ) , .ZN( u0_u13_u3_n134 ) , .B1( u0_u13_u3_n143 ) , .B2( u0_u13_u3_n177 ) );
  NAND2_X1 u0_u13_u3_U60 (.A1( u0_u13_u3_n100 ) , .ZN( u0_u13_u3_n156 ) , .A2( u0_u13_u3_n99 ) );
  NAND2_X1 u0_u13_u3_U61 (.A2( u0_u13_u3_n101 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n148 ) );
  NAND2_X1 u0_u13_u3_U62 (.A1( u0_u13_u3_n100 ) , .A2( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n128 ) );
  NAND2_X1 u0_u13_u3_U63 (.A2( u0_u13_u3_n101 ) , .A1( u0_u13_u3_n102 ) , .ZN( u0_u13_u3_n152 ) );
  NAND2_X1 u0_u13_u3_U64 (.A2( u0_u13_u3_n101 ) , .ZN( u0_u13_u3_n114 ) , .A1( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U65 (.ZN( u0_u13_u3_n107 ) , .A1( u0_u13_u3_n97 ) , .A2( u0_u13_u3_n99 ) );
  NAND2_X1 u0_u13_u3_U66 (.A2( u0_u13_u3_n100 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n113 ) );
  NAND2_X1 u0_u13_u3_U67 (.A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n153 ) , .A2( u0_u13_u3_n97 ) );
  NAND2_X1 u0_u13_u3_U68 (.A2( u0_u13_u3_n103 ) , .A1( u0_u13_u3_n104 ) , .ZN( u0_u13_u3_n130 ) );
  NAND2_X1 u0_u13_u3_U69 (.A2( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n144 ) , .A1( u0_u13_u3_n96 ) );
  OAI22_X1 u0_u13_u3_U7 (.B2( u0_u13_u3_n147 ) , .A2( u0_u13_u3_n148 ) , .ZN( u0_u13_u3_n160 ) , .B1( u0_u13_u3_n165 ) , .A1( u0_u13_u3_n168 ) );
  NAND2_X1 u0_u13_u3_U70 (.A1( u0_u13_u3_n102 ) , .A2( u0_u13_u3_n103 ) , .ZN( u0_u13_u3_n108 ) );
  NOR2_X1 u0_u13_u3_U71 (.A2( u0_u13_X_19 ) , .A1( u0_u13_X_20 ) , .ZN( u0_u13_u3_n99 ) );
  NOR2_X1 u0_u13_u3_U72 (.A2( u0_u13_X_21 ) , .A1( u0_u13_X_24 ) , .ZN( u0_u13_u3_n103 ) );
  NOR2_X1 u0_u13_u3_U73 (.A2( u0_u13_X_24 ) , .A1( u0_u13_u3_n171 ) , .ZN( u0_u13_u3_n97 ) );
  NOR2_X1 u0_u13_u3_U74 (.A2( u0_u13_X_23 ) , .ZN( u0_u13_u3_n141 ) , .A1( u0_u13_u3_n166 ) );
  NOR2_X1 u0_u13_u3_U75 (.A2( u0_u13_X_19 ) , .A1( u0_u13_u3_n172 ) , .ZN( u0_u13_u3_n96 ) );
  NAND2_X1 u0_u13_u3_U76 (.A1( u0_u13_X_22 ) , .A2( u0_u13_X_23 ) , .ZN( u0_u13_u3_n154 ) );
  NAND2_X1 u0_u13_u3_U77 (.A1( u0_u13_X_23 ) , .ZN( u0_u13_u3_n149 ) , .A2( u0_u13_u3_n166 ) );
  NOR2_X1 u0_u13_u3_U78 (.A2( u0_u13_X_22 ) , .A1( u0_u13_X_23 ) , .ZN( u0_u13_u3_n121 ) );
  AND2_X1 u0_u13_u3_U79 (.A1( u0_u13_X_24 ) , .ZN( u0_u13_u3_n101 ) , .A2( u0_u13_u3_n171 ) );
  AND3_X1 u0_u13_u3_U8 (.A3( u0_u13_u3_n144 ) , .A2( u0_u13_u3_n145 ) , .A1( u0_u13_u3_n146 ) , .ZN( u0_u13_u3_n147 ) );
  AND2_X1 u0_u13_u3_U80 (.A1( u0_u13_X_19 ) , .ZN( u0_u13_u3_n102 ) , .A2( u0_u13_u3_n172 ) );
  AND2_X1 u0_u13_u3_U81 (.A1( u0_u13_X_21 ) , .A2( u0_u13_X_24 ) , .ZN( u0_u13_u3_n100 ) );
  AND2_X1 u0_u13_u3_U82 (.A2( u0_u13_X_19 ) , .A1( u0_u13_X_20 ) , .ZN( u0_u13_u3_n104 ) );
  INV_X1 u0_u13_u3_U83 (.A( u0_u13_X_22 ) , .ZN( u0_u13_u3_n166 ) );
  INV_X1 u0_u13_u3_U84 (.A( u0_u13_X_21 ) , .ZN( u0_u13_u3_n171 ) );
  INV_X1 u0_u13_u3_U85 (.A( u0_u13_X_20 ) , .ZN( u0_u13_u3_n172 ) );
  NAND4_X1 u0_u13_u3_U86 (.ZN( u0_out13_26 ) , .A4( u0_u13_u3_n109 ) , .A3( u0_u13_u3_n110 ) , .A2( u0_u13_u3_n111 ) , .A1( u0_u13_u3_n173 ) );
  INV_X1 u0_u13_u3_U87 (.ZN( u0_u13_u3_n173 ) , .A( u0_u13_u3_n94 ) );
  OAI21_X1 u0_u13_u3_U88 (.ZN( u0_u13_u3_n111 ) , .B2( u0_u13_u3_n117 ) , .A( u0_u13_u3_n133 ) , .B1( u0_u13_u3_n176 ) );
  NAND4_X1 u0_u13_u3_U89 (.ZN( u0_out13_20 ) , .A4( u0_u13_u3_n122 ) , .A3( u0_u13_u3_n123 ) , .A1( u0_u13_u3_n175 ) , .A2( u0_u13_u3_n180 ) );
  INV_X1 u0_u13_u3_U9 (.A( u0_u13_u3_n143 ) , .ZN( u0_u13_u3_n168 ) );
  INV_X1 u0_u13_u3_U90 (.A( u0_u13_u3_n112 ) , .ZN( u0_u13_u3_n175 ) );
  INV_X1 u0_u13_u3_U91 (.A( u0_u13_u3_n126 ) , .ZN( u0_u13_u3_n180 ) );
  NAND4_X1 u0_u13_u3_U92 (.ZN( u0_out13_1 ) , .A4( u0_u13_u3_n161 ) , .A3( u0_u13_u3_n162 ) , .A2( u0_u13_u3_n163 ) , .A1( u0_u13_u3_n185 ) );
  NAND2_X1 u0_u13_u3_U93 (.ZN( u0_u13_u3_n163 ) , .A2( u0_u13_u3_n170 ) , .A1( u0_u13_u3_n176 ) );
  AOI22_X1 u0_u13_u3_U94 (.B2( u0_u13_u3_n140 ) , .B1( u0_u13_u3_n141 ) , .A2( u0_u13_u3_n142 ) , .ZN( u0_u13_u3_n162 ) , .A1( u0_u13_u3_n177 ) );
  OR4_X1 u0_u13_u3_U95 (.ZN( u0_out13_10 ) , .A4( u0_u13_u3_n136 ) , .A3( u0_u13_u3_n137 ) , .A1( u0_u13_u3_n138 ) , .A2( u0_u13_u3_n139 ) );
  OAI222_X1 u0_u13_u3_U96 (.C1( u0_u13_u3_n128 ) , .ZN( u0_u13_u3_n137 ) , .B1( u0_u13_u3_n148 ) , .A2( u0_u13_u3_n150 ) , .B2( u0_u13_u3_n154 ) , .C2( u0_u13_u3_n164 ) , .A1( u0_u13_u3_n167 ) );
  OAI221_X1 u0_u13_u3_U97 (.A( u0_u13_u3_n134 ) , .B2( u0_u13_u3_n135 ) , .ZN( u0_u13_u3_n136 ) , .C1( u0_u13_u3_n149 ) , .B1( u0_u13_u3_n151 ) , .C2( u0_u13_u3_n183 ) );
  NAND3_X1 u0_u13_u3_U98 (.A1( u0_u13_u3_n114 ) , .ZN( u0_u13_u3_n115 ) , .A2( u0_u13_u3_n145 ) , .A3( u0_u13_u3_n153 ) );
  NAND3_X1 u0_u13_u3_U99 (.ZN( u0_u13_u3_n129 ) , .A2( u0_u13_u3_n144 ) , .A1( u0_u13_u3_n153 ) , .A3( u0_u13_u3_n182 ) );
  AOI21_X1 u0_u13_u4_U10 (.ZN( u0_u13_u4_n106 ) , .B2( u0_u13_u4_n146 ) , .B1( u0_u13_u4_n158 ) , .A( u0_u13_u4_n170 ) );
  AOI21_X1 u0_u13_u4_U11 (.ZN( u0_u13_u4_n108 ) , .B2( u0_u13_u4_n134 ) , .B1( u0_u13_u4_n155 ) , .A( u0_u13_u4_n156 ) );
  AOI21_X1 u0_u13_u4_U12 (.ZN( u0_u13_u4_n109 ) , .A( u0_u13_u4_n153 ) , .B1( u0_u13_u4_n159 ) , .B2( u0_u13_u4_n184 ) );
  AOI211_X1 u0_u13_u4_U13 (.B( u0_u13_u4_n136 ) , .A( u0_u13_u4_n137 ) , .C2( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n139 ) , .C1( u0_u13_u4_n182 ) );
  OAI22_X1 u0_u13_u4_U14 (.B2( u0_u13_u4_n135 ) , .ZN( u0_u13_u4_n137 ) , .B1( u0_u13_u4_n153 ) , .A1( u0_u13_u4_n155 ) , .A2( u0_u13_u4_n171 ) );
  AND3_X1 u0_u13_u4_U15 (.A2( u0_u13_u4_n134 ) , .ZN( u0_u13_u4_n135 ) , .A3( u0_u13_u4_n145 ) , .A1( u0_u13_u4_n157 ) );
  NAND2_X1 u0_u13_u4_U16 (.ZN( u0_u13_u4_n132 ) , .A2( u0_u13_u4_n170 ) , .A1( u0_u13_u4_n173 ) );
  AOI21_X1 u0_u13_u4_U17 (.B2( u0_u13_u4_n160 ) , .B1( u0_u13_u4_n161 ) , .ZN( u0_u13_u4_n162 ) , .A( u0_u13_u4_n170 ) );
  AOI21_X1 u0_u13_u4_U18 (.ZN( u0_u13_u4_n107 ) , .B2( u0_u13_u4_n143 ) , .A( u0_u13_u4_n174 ) , .B1( u0_u13_u4_n184 ) );
  AOI21_X1 u0_u13_u4_U19 (.B2( u0_u13_u4_n158 ) , .B1( u0_u13_u4_n159 ) , .ZN( u0_u13_u4_n163 ) , .A( u0_u13_u4_n174 ) );
  AOI21_X1 u0_u13_u4_U20 (.A( u0_u13_u4_n153 ) , .B2( u0_u13_u4_n154 ) , .B1( u0_u13_u4_n155 ) , .ZN( u0_u13_u4_n165 ) );
  AOI21_X1 u0_u13_u4_U21 (.A( u0_u13_u4_n156 ) , .B2( u0_u13_u4_n157 ) , .ZN( u0_u13_u4_n164 ) , .B1( u0_u13_u4_n184 ) );
  INV_X1 u0_u13_u4_U22 (.A( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n170 ) );
  AND2_X1 u0_u13_u4_U23 (.A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n155 ) , .A1( u0_u13_u4_n160 ) );
  INV_X1 u0_u13_u4_U24 (.A( u0_u13_u4_n156 ) , .ZN( u0_u13_u4_n175 ) );
  NAND2_X1 u0_u13_u4_U25 (.A2( u0_u13_u4_n118 ) , .ZN( u0_u13_u4_n131 ) , .A1( u0_u13_u4_n147 ) );
  NAND2_X1 u0_u13_u4_U26 (.A1( u0_u13_u4_n119 ) , .A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n130 ) );
  NAND2_X1 u0_u13_u4_U27 (.ZN( u0_u13_u4_n117 ) , .A2( u0_u13_u4_n118 ) , .A1( u0_u13_u4_n148 ) );
  NAND2_X1 u0_u13_u4_U28 (.ZN( u0_u13_u4_n129 ) , .A1( u0_u13_u4_n134 ) , .A2( u0_u13_u4_n148 ) );
  AND3_X1 u0_u13_u4_U29 (.A1( u0_u13_u4_n119 ) , .A2( u0_u13_u4_n143 ) , .A3( u0_u13_u4_n154 ) , .ZN( u0_u13_u4_n161 ) );
  NOR2_X1 u0_u13_u4_U3 (.ZN( u0_u13_u4_n121 ) , .A1( u0_u13_u4_n181 ) , .A2( u0_u13_u4_n182 ) );
  AND2_X1 u0_u13_u4_U30 (.A1( u0_u13_u4_n145 ) , .A2( u0_u13_u4_n147 ) , .ZN( u0_u13_u4_n159 ) );
  OR3_X1 u0_u13_u4_U31 (.A3( u0_u13_u4_n114 ) , .A2( u0_u13_u4_n115 ) , .A1( u0_u13_u4_n116 ) , .ZN( u0_u13_u4_n136 ) );
  AOI21_X1 u0_u13_u4_U32 (.A( u0_u13_u4_n113 ) , .ZN( u0_u13_u4_n116 ) , .B2( u0_u13_u4_n173 ) , .B1( u0_u13_u4_n174 ) );
  AOI21_X1 u0_u13_u4_U33 (.ZN( u0_u13_u4_n115 ) , .B2( u0_u13_u4_n145 ) , .B1( u0_u13_u4_n146 ) , .A( u0_u13_u4_n156 ) );
  OAI22_X1 u0_u13_u4_U34 (.ZN( u0_u13_u4_n114 ) , .A2( u0_u13_u4_n121 ) , .B1( u0_u13_u4_n160 ) , .B2( u0_u13_u4_n170 ) , .A1( u0_u13_u4_n171 ) );
  INV_X1 u0_u13_u4_U35 (.A( u0_u13_u4_n158 ) , .ZN( u0_u13_u4_n182 ) );
  INV_X1 u0_u13_u4_U36 (.ZN( u0_u13_u4_n181 ) , .A( u0_u13_u4_n96 ) );
  INV_X1 u0_u13_u4_U37 (.A( u0_u13_u4_n144 ) , .ZN( u0_u13_u4_n179 ) );
  INV_X1 u0_u13_u4_U38 (.A( u0_u13_u4_n157 ) , .ZN( u0_u13_u4_n178 ) );
  NAND2_X1 u0_u13_u4_U39 (.A2( u0_u13_u4_n154 ) , .A1( u0_u13_u4_n96 ) , .ZN( u0_u13_u4_n97 ) );
  INV_X1 u0_u13_u4_U4 (.A( u0_u13_u4_n117 ) , .ZN( u0_u13_u4_n184 ) );
  INV_X1 u0_u13_u4_U40 (.A( u0_u13_u4_n143 ) , .ZN( u0_u13_u4_n183 ) );
  NOR2_X1 u0_u13_u4_U41 (.ZN( u0_u13_u4_n138 ) , .A1( u0_u13_u4_n168 ) , .A2( u0_u13_u4_n169 ) );
  NOR2_X1 u0_u13_u4_U42 (.A1( u0_u13_u4_n150 ) , .A2( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n153 ) );
  NOR2_X1 u0_u13_u4_U43 (.A2( u0_u13_u4_n128 ) , .A1( u0_u13_u4_n138 ) , .ZN( u0_u13_u4_n156 ) );
  AOI22_X1 u0_u13_u4_U44 (.B2( u0_u13_u4_n122 ) , .A1( u0_u13_u4_n123 ) , .ZN( u0_u13_u4_n124 ) , .B1( u0_u13_u4_n128 ) , .A2( u0_u13_u4_n172 ) );
  NAND2_X1 u0_u13_u4_U45 (.A2( u0_u13_u4_n120 ) , .ZN( u0_u13_u4_n123 ) , .A1( u0_u13_u4_n161 ) );
  INV_X1 u0_u13_u4_U46 (.A( u0_u13_u4_n153 ) , .ZN( u0_u13_u4_n172 ) );
  AOI22_X1 u0_u13_u4_U47 (.B2( u0_u13_u4_n132 ) , .A2( u0_u13_u4_n133 ) , .ZN( u0_u13_u4_n140 ) , .A1( u0_u13_u4_n150 ) , .B1( u0_u13_u4_n179 ) );
  NAND2_X1 u0_u13_u4_U48 (.ZN( u0_u13_u4_n133 ) , .A2( u0_u13_u4_n146 ) , .A1( u0_u13_u4_n154 ) );
  NAND2_X1 u0_u13_u4_U49 (.A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n154 ) , .A2( u0_u13_u4_n98 ) );
  INV_X1 u0_u13_u4_U5 (.ZN( u0_u13_u4_n186 ) , .A( u0_u13_u4_n95 ) );
  NAND2_X1 u0_u13_u4_U50 (.A1( u0_u13_u4_n101 ) , .ZN( u0_u13_u4_n158 ) , .A2( u0_u13_u4_n99 ) );
  AOI21_X1 u0_u13_u4_U51 (.ZN( u0_u13_u4_n127 ) , .A( u0_u13_u4_n136 ) , .B2( u0_u13_u4_n150 ) , .B1( u0_u13_u4_n180 ) );
  INV_X1 u0_u13_u4_U52 (.A( u0_u13_u4_n160 ) , .ZN( u0_u13_u4_n180 ) );
  NAND2_X1 u0_u13_u4_U53 (.A2( u0_u13_u4_n104 ) , .A1( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n146 ) );
  NAND2_X1 u0_u13_u4_U54 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n160 ) );
  NAND2_X1 u0_u13_u4_U55 (.ZN( u0_u13_u4_n134 ) , .A1( u0_u13_u4_n98 ) , .A2( u0_u13_u4_n99 ) );
  NAND2_X1 u0_u13_u4_U56 (.A1( u0_u13_u4_n103 ) , .A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n143 ) );
  NAND2_X1 u0_u13_u4_U57 (.A2( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n145 ) , .A1( u0_u13_u4_n98 ) );
  NAND2_X1 u0_u13_u4_U58 (.A1( u0_u13_u4_n100 ) , .A2( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n120 ) );
  NAND2_X1 u0_u13_u4_U59 (.A1( u0_u13_u4_n102 ) , .A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n148 ) );
  OAI221_X1 u0_u13_u4_U6 (.C1( u0_u13_u4_n134 ) , .B1( u0_u13_u4_n158 ) , .B2( u0_u13_u4_n171 ) , .C2( u0_u13_u4_n173 ) , .A( u0_u13_u4_n94 ) , .ZN( u0_u13_u4_n95 ) );
  NAND2_X1 u0_u13_u4_U60 (.A2( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n157 ) );
  INV_X1 u0_u13_u4_U61 (.A( u0_u13_u4_n150 ) , .ZN( u0_u13_u4_n173 ) );
  INV_X1 u0_u13_u4_U62 (.A( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n171 ) );
  NAND2_X1 u0_u13_u4_U63 (.A1( u0_u13_u4_n100 ) , .ZN( u0_u13_u4_n118 ) , .A2( u0_u13_u4_n99 ) );
  NAND2_X1 u0_u13_u4_U64 (.A2( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n144 ) );
  NAND2_X1 u0_u13_u4_U65 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n105 ) , .ZN( u0_u13_u4_n96 ) );
  INV_X1 u0_u13_u4_U66 (.A( u0_u13_u4_n128 ) , .ZN( u0_u13_u4_n174 ) );
  NAND2_X1 u0_u13_u4_U67 (.A2( u0_u13_u4_n102 ) , .ZN( u0_u13_u4_n119 ) , .A1( u0_u13_u4_n98 ) );
  NAND2_X1 u0_u13_u4_U68 (.A2( u0_u13_u4_n101 ) , .A1( u0_u13_u4_n103 ) , .ZN( u0_u13_u4_n147 ) );
  NAND2_X1 u0_u13_u4_U69 (.A2( u0_u13_u4_n104 ) , .ZN( u0_u13_u4_n113 ) , .A1( u0_u13_u4_n99 ) );
  AOI222_X1 u0_u13_u4_U7 (.B2( u0_u13_u4_n132 ) , .A1( u0_u13_u4_n138 ) , .C2( u0_u13_u4_n175 ) , .A2( u0_u13_u4_n179 ) , .C1( u0_u13_u4_n181 ) , .B1( u0_u13_u4_n185 ) , .ZN( u0_u13_u4_n94 ) );
  NOR2_X1 u0_u13_u4_U70 (.A2( u0_u13_X_28 ) , .ZN( u0_u13_u4_n150 ) , .A1( u0_u13_u4_n168 ) );
  NOR2_X1 u0_u13_u4_U71 (.A2( u0_u13_X_29 ) , .ZN( u0_u13_u4_n152 ) , .A1( u0_u13_u4_n169 ) );
  NOR2_X1 u0_u13_u4_U72 (.A2( u0_u13_X_30 ) , .ZN( u0_u13_u4_n105 ) , .A1( u0_u13_u4_n176 ) );
  NOR2_X1 u0_u13_u4_U73 (.A2( u0_u13_X_26 ) , .ZN( u0_u13_u4_n100 ) , .A1( u0_u13_u4_n177 ) );
  NOR2_X1 u0_u13_u4_U74 (.A2( u0_u13_X_28 ) , .A1( u0_u13_X_29 ) , .ZN( u0_u13_u4_n128 ) );
  NOR2_X1 u0_u13_u4_U75 (.A2( u0_u13_X_27 ) , .A1( u0_u13_X_30 ) , .ZN( u0_u13_u4_n102 ) );
  NOR2_X1 u0_u13_u4_U76 (.A2( u0_u13_X_25 ) , .A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n98 ) );
  AND2_X1 u0_u13_u4_U77 (.A2( u0_u13_X_25 ) , .A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n104 ) );
  AND2_X1 u0_u13_u4_U78 (.A1( u0_u13_X_30 ) , .A2( u0_u13_u4_n176 ) , .ZN( u0_u13_u4_n99 ) );
  AND2_X1 u0_u13_u4_U79 (.A1( u0_u13_X_26 ) , .ZN( u0_u13_u4_n101 ) , .A2( u0_u13_u4_n177 ) );
  INV_X1 u0_u13_u4_U8 (.A( u0_u13_u4_n113 ) , .ZN( u0_u13_u4_n185 ) );
  AND2_X1 u0_u13_u4_U80 (.A1( u0_u13_X_27 ) , .A2( u0_u13_X_30 ) , .ZN( u0_u13_u4_n103 ) );
  INV_X1 u0_u13_u4_U81 (.A( u0_u13_X_28 ) , .ZN( u0_u13_u4_n169 ) );
  INV_X1 u0_u13_u4_U82 (.A( u0_u13_X_29 ) , .ZN( u0_u13_u4_n168 ) );
  INV_X1 u0_u13_u4_U83 (.A( u0_u13_X_25 ) , .ZN( u0_u13_u4_n177 ) );
  INV_X1 u0_u13_u4_U84 (.A( u0_u13_X_27 ) , .ZN( u0_u13_u4_n176 ) );
  NAND4_X1 u0_u13_u4_U85 (.ZN( u0_out13_25 ) , .A4( u0_u13_u4_n139 ) , .A3( u0_u13_u4_n140 ) , .A2( u0_u13_u4_n141 ) , .A1( u0_u13_u4_n142 ) );
  OAI21_X1 u0_u13_u4_U86 (.A( u0_u13_u4_n128 ) , .B2( u0_u13_u4_n129 ) , .B1( u0_u13_u4_n130 ) , .ZN( u0_u13_u4_n142 ) );
  OAI21_X1 u0_u13_u4_U87 (.B2( u0_u13_u4_n131 ) , .ZN( u0_u13_u4_n141 ) , .A( u0_u13_u4_n175 ) , .B1( u0_u13_u4_n183 ) );
  NAND4_X1 u0_u13_u4_U88 (.ZN( u0_out13_14 ) , .A4( u0_u13_u4_n124 ) , .A3( u0_u13_u4_n125 ) , .A2( u0_u13_u4_n126 ) , .A1( u0_u13_u4_n127 ) );
  AOI22_X1 u0_u13_u4_U89 (.B2( u0_u13_u4_n117 ) , .ZN( u0_u13_u4_n126 ) , .A1( u0_u13_u4_n129 ) , .B1( u0_u13_u4_n152 ) , .A2( u0_u13_u4_n175 ) );
  NOR4_X1 u0_u13_u4_U9 (.A4( u0_u13_u4_n106 ) , .A3( u0_u13_u4_n107 ) , .A2( u0_u13_u4_n108 ) , .A1( u0_u13_u4_n109 ) , .ZN( u0_u13_u4_n110 ) );
  AOI22_X1 u0_u13_u4_U90 (.ZN( u0_u13_u4_n125 ) , .B2( u0_u13_u4_n131 ) , .A2( u0_u13_u4_n132 ) , .B1( u0_u13_u4_n138 ) , .A1( u0_u13_u4_n178 ) );
  NAND4_X1 u0_u13_u4_U91 (.ZN( u0_out13_8 ) , .A4( u0_u13_u4_n110 ) , .A3( u0_u13_u4_n111 ) , .A2( u0_u13_u4_n112 ) , .A1( u0_u13_u4_n186 ) );
  NAND2_X1 u0_u13_u4_U92 (.ZN( u0_u13_u4_n112 ) , .A2( u0_u13_u4_n130 ) , .A1( u0_u13_u4_n150 ) );
  AOI22_X1 u0_u13_u4_U93 (.ZN( u0_u13_u4_n111 ) , .B2( u0_u13_u4_n132 ) , .A1( u0_u13_u4_n152 ) , .B1( u0_u13_u4_n178 ) , .A2( u0_u13_u4_n97 ) );
  AOI22_X1 u0_u13_u4_U94 (.B2( u0_u13_u4_n149 ) , .B1( u0_u13_u4_n150 ) , .A2( u0_u13_u4_n151 ) , .A1( u0_u13_u4_n152 ) , .ZN( u0_u13_u4_n167 ) );
  NOR4_X1 u0_u13_u4_U95 (.A4( u0_u13_u4_n162 ) , .A3( u0_u13_u4_n163 ) , .A2( u0_u13_u4_n164 ) , .A1( u0_u13_u4_n165 ) , .ZN( u0_u13_u4_n166 ) );
  NAND3_X1 u0_u13_u4_U96 (.ZN( u0_out13_3 ) , .A3( u0_u13_u4_n166 ) , .A1( u0_u13_u4_n167 ) , .A2( u0_u13_u4_n186 ) );
  NAND3_X1 u0_u13_u4_U97 (.A3( u0_u13_u4_n146 ) , .A2( u0_u13_u4_n147 ) , .A1( u0_u13_u4_n148 ) , .ZN( u0_u13_u4_n149 ) );
  NAND3_X1 u0_u13_u4_U98 (.A3( u0_u13_u4_n143 ) , .A2( u0_u13_u4_n144 ) , .A1( u0_u13_u4_n145 ) , .ZN( u0_u13_u4_n151 ) );
  NAND3_X1 u0_u13_u4_U99 (.A3( u0_u13_u4_n121 ) , .ZN( u0_u13_u4_n122 ) , .A2( u0_u13_u4_n144 ) , .A1( u0_u13_u4_n154 ) );
  XOR2_X1 u0_u9_U10 (.B( u0_K10_45 ) , .A( u0_R8_30 ) , .Z( u0_u9_X_45 ) );
  XOR2_X1 u0_u9_U11 (.B( u0_K10_44 ) , .A( u0_R8_29 ) , .Z( u0_u9_X_44 ) );
  XOR2_X1 u0_u9_U12 (.B( u0_K10_43 ) , .A( u0_R8_28 ) , .Z( u0_u9_X_43 ) );
  XOR2_X1 u0_u9_U20 (.B( u0_K10_36 ) , .A( u0_R8_25 ) , .Z( u0_u9_X_36 ) );
  XOR2_X1 u0_u9_U21 (.B( u0_K10_35 ) , .A( u0_R8_24 ) , .Z( u0_u9_X_35 ) );
  XOR2_X1 u0_u9_U22 (.B( u0_K10_34 ) , .A( u0_R8_23 ) , .Z( u0_u9_X_34 ) );
  XOR2_X1 u0_u9_U23 (.B( u0_K10_33 ) , .A( u0_R8_22 ) , .Z( u0_u9_X_33 ) );
  XOR2_X1 u0_u9_U24 (.B( u0_K10_32 ) , .A( u0_R8_21 ) , .Z( u0_u9_X_32 ) );
  XOR2_X1 u0_u9_U25 (.B( u0_K10_31 ) , .A( u0_R8_20 ) , .Z( u0_u9_X_31 ) );
  XOR2_X1 u0_u9_U26 (.B( u0_K10_30 ) , .A( u0_R8_21 ) , .Z( u0_u9_X_30 ) );
  XOR2_X1 u0_u9_U28 (.B( u0_K10_29 ) , .A( u0_R8_20 ) , .Z( u0_u9_X_29 ) );
  XOR2_X1 u0_u9_U29 (.B( u0_K10_28 ) , .A( u0_R8_19 ) , .Z( u0_u9_X_28 ) );
  XOR2_X1 u0_u9_U30 (.B( u0_K10_27 ) , .A( u0_R8_18 ) , .Z( u0_u9_X_27 ) );
  XOR2_X1 u0_u9_U31 (.B( u0_K10_26 ) , .A( u0_R8_17 ) , .Z( u0_u9_X_26 ) );
  XOR2_X1 u0_u9_U32 (.B( u0_K10_25 ) , .A( u0_R8_16 ) , .Z( u0_u9_X_25 ) );
  XOR2_X1 u0_u9_U7 (.B( u0_K10_48 ) , .A( u0_R8_1 ) , .Z( u0_u9_X_48 ) );
  XOR2_X1 u0_u9_U8 (.B( u0_K10_47 ) , .A( u0_R8_32 ) , .Z( u0_u9_X_47 ) );
  XOR2_X1 u0_u9_U9 (.B( u0_K10_46 ) , .A( u0_R8_31 ) , .Z( u0_u9_X_46 ) );
  OAI22_X1 u0_u9_u4_U10 (.B2( u0_u9_u4_n135 ) , .ZN( u0_u9_u4_n137 ) , .B1( u0_u9_u4_n153 ) , .A1( u0_u9_u4_n155 ) , .A2( u0_u9_u4_n171 ) );
  AND3_X1 u0_u9_u4_U11 (.A2( u0_u9_u4_n134 ) , .ZN( u0_u9_u4_n135 ) , .A3( u0_u9_u4_n145 ) , .A1( u0_u9_u4_n157 ) );
  NAND2_X1 u0_u9_u4_U12 (.ZN( u0_u9_u4_n132 ) , .A2( u0_u9_u4_n170 ) , .A1( u0_u9_u4_n173 ) );
  AOI21_X1 u0_u9_u4_U13 (.B2( u0_u9_u4_n160 ) , .B1( u0_u9_u4_n161 ) , .ZN( u0_u9_u4_n162 ) , .A( u0_u9_u4_n170 ) );
  AOI21_X1 u0_u9_u4_U14 (.ZN( u0_u9_u4_n107 ) , .B2( u0_u9_u4_n143 ) , .A( u0_u9_u4_n174 ) , .B1( u0_u9_u4_n184 ) );
  AOI21_X1 u0_u9_u4_U15 (.B2( u0_u9_u4_n158 ) , .B1( u0_u9_u4_n159 ) , .ZN( u0_u9_u4_n163 ) , .A( u0_u9_u4_n174 ) );
  AOI21_X1 u0_u9_u4_U16 (.A( u0_u9_u4_n153 ) , .B2( u0_u9_u4_n154 ) , .B1( u0_u9_u4_n155 ) , .ZN( u0_u9_u4_n165 ) );
  AOI21_X1 u0_u9_u4_U17 (.A( u0_u9_u4_n156 ) , .B2( u0_u9_u4_n157 ) , .ZN( u0_u9_u4_n164 ) , .B1( u0_u9_u4_n184 ) );
  INV_X1 u0_u9_u4_U18 (.A( u0_u9_u4_n138 ) , .ZN( u0_u9_u4_n170 ) );
  AND2_X1 u0_u9_u4_U19 (.A2( u0_u9_u4_n120 ) , .ZN( u0_u9_u4_n155 ) , .A1( u0_u9_u4_n160 ) );
  INV_X1 u0_u9_u4_U20 (.A( u0_u9_u4_n156 ) , .ZN( u0_u9_u4_n175 ) );
  NAND2_X1 u0_u9_u4_U21 (.A2( u0_u9_u4_n118 ) , .ZN( u0_u9_u4_n131 ) , .A1( u0_u9_u4_n147 ) );
  NAND2_X1 u0_u9_u4_U22 (.A1( u0_u9_u4_n119 ) , .A2( u0_u9_u4_n120 ) , .ZN( u0_u9_u4_n130 ) );
  NAND2_X1 u0_u9_u4_U23 (.ZN( u0_u9_u4_n117 ) , .A2( u0_u9_u4_n118 ) , .A1( u0_u9_u4_n148 ) );
  NAND2_X1 u0_u9_u4_U24 (.ZN( u0_u9_u4_n129 ) , .A1( u0_u9_u4_n134 ) , .A2( u0_u9_u4_n148 ) );
  AND3_X1 u0_u9_u4_U25 (.A1( u0_u9_u4_n119 ) , .A2( u0_u9_u4_n143 ) , .A3( u0_u9_u4_n154 ) , .ZN( u0_u9_u4_n161 ) );
  AND2_X1 u0_u9_u4_U26 (.A1( u0_u9_u4_n145 ) , .A2( u0_u9_u4_n147 ) , .ZN( u0_u9_u4_n159 ) );
  OR3_X1 u0_u9_u4_U27 (.A3( u0_u9_u4_n114 ) , .A2( u0_u9_u4_n115 ) , .A1( u0_u9_u4_n116 ) , .ZN( u0_u9_u4_n136 ) );
  AOI21_X1 u0_u9_u4_U28 (.A( u0_u9_u4_n113 ) , .ZN( u0_u9_u4_n116 ) , .B2( u0_u9_u4_n173 ) , .B1( u0_u9_u4_n174 ) );
  AOI21_X1 u0_u9_u4_U29 (.ZN( u0_u9_u4_n115 ) , .B2( u0_u9_u4_n145 ) , .B1( u0_u9_u4_n146 ) , .A( u0_u9_u4_n156 ) );
  NOR2_X1 u0_u9_u4_U3 (.ZN( u0_u9_u4_n121 ) , .A1( u0_u9_u4_n181 ) , .A2( u0_u9_u4_n182 ) );
  OAI22_X1 u0_u9_u4_U30 (.ZN( u0_u9_u4_n114 ) , .A2( u0_u9_u4_n121 ) , .B1( u0_u9_u4_n160 ) , .B2( u0_u9_u4_n170 ) , .A1( u0_u9_u4_n171 ) );
  INV_X1 u0_u9_u4_U31 (.A( u0_u9_u4_n158 ) , .ZN( u0_u9_u4_n182 ) );
  INV_X1 u0_u9_u4_U32 (.ZN( u0_u9_u4_n181 ) , .A( u0_u9_u4_n96 ) );
  INV_X1 u0_u9_u4_U33 (.A( u0_u9_u4_n144 ) , .ZN( u0_u9_u4_n179 ) );
  INV_X1 u0_u9_u4_U34 (.A( u0_u9_u4_n157 ) , .ZN( u0_u9_u4_n178 ) );
  NAND2_X1 u0_u9_u4_U35 (.A2( u0_u9_u4_n154 ) , .A1( u0_u9_u4_n96 ) , .ZN( u0_u9_u4_n97 ) );
  INV_X1 u0_u9_u4_U36 (.ZN( u0_u9_u4_n186 ) , .A( u0_u9_u4_n95 ) );
  OAI221_X1 u0_u9_u4_U37 (.C1( u0_u9_u4_n134 ) , .B1( u0_u9_u4_n158 ) , .B2( u0_u9_u4_n171 ) , .C2( u0_u9_u4_n173 ) , .A( u0_u9_u4_n94 ) , .ZN( u0_u9_u4_n95 ) );
  AOI222_X1 u0_u9_u4_U38 (.B2( u0_u9_u4_n132 ) , .A1( u0_u9_u4_n138 ) , .C2( u0_u9_u4_n175 ) , .A2( u0_u9_u4_n179 ) , .C1( u0_u9_u4_n181 ) , .B1( u0_u9_u4_n185 ) , .ZN( u0_u9_u4_n94 ) );
  INV_X1 u0_u9_u4_U39 (.A( u0_u9_u4_n113 ) , .ZN( u0_u9_u4_n185 ) );
  INV_X1 u0_u9_u4_U4 (.A( u0_u9_u4_n117 ) , .ZN( u0_u9_u4_n184 ) );
  INV_X1 u0_u9_u4_U40 (.A( u0_u9_u4_n143 ) , .ZN( u0_u9_u4_n183 ) );
  NOR2_X1 u0_u9_u4_U41 (.ZN( u0_u9_u4_n138 ) , .A1( u0_u9_u4_n168 ) , .A2( u0_u9_u4_n169 ) );
  NOR2_X1 u0_u9_u4_U42 (.A1( u0_u9_u4_n150 ) , .A2( u0_u9_u4_n152 ) , .ZN( u0_u9_u4_n153 ) );
  NOR2_X1 u0_u9_u4_U43 (.A2( u0_u9_u4_n128 ) , .A1( u0_u9_u4_n138 ) , .ZN( u0_u9_u4_n156 ) );
  AOI22_X1 u0_u9_u4_U44 (.B2( u0_u9_u4_n122 ) , .A1( u0_u9_u4_n123 ) , .ZN( u0_u9_u4_n124 ) , .B1( u0_u9_u4_n128 ) , .A2( u0_u9_u4_n172 ) );
  INV_X1 u0_u9_u4_U45 (.A( u0_u9_u4_n153 ) , .ZN( u0_u9_u4_n172 ) );
  NAND2_X1 u0_u9_u4_U46 (.A2( u0_u9_u4_n120 ) , .ZN( u0_u9_u4_n123 ) , .A1( u0_u9_u4_n161 ) );
  AOI22_X1 u0_u9_u4_U47 (.B2( u0_u9_u4_n132 ) , .A2( u0_u9_u4_n133 ) , .ZN( u0_u9_u4_n140 ) , .A1( u0_u9_u4_n150 ) , .B1( u0_u9_u4_n179 ) );
  NAND2_X1 u0_u9_u4_U48 (.ZN( u0_u9_u4_n133 ) , .A2( u0_u9_u4_n146 ) , .A1( u0_u9_u4_n154 ) );
  NAND2_X1 u0_u9_u4_U49 (.A1( u0_u9_u4_n103 ) , .ZN( u0_u9_u4_n154 ) , .A2( u0_u9_u4_n98 ) );
  NOR4_X1 u0_u9_u4_U5 (.A4( u0_u9_u4_n106 ) , .A3( u0_u9_u4_n107 ) , .A2( u0_u9_u4_n108 ) , .A1( u0_u9_u4_n109 ) , .ZN( u0_u9_u4_n110 ) );
  NAND2_X1 u0_u9_u4_U50 (.A1( u0_u9_u4_n101 ) , .ZN( u0_u9_u4_n158 ) , .A2( u0_u9_u4_n99 ) );
  AOI21_X1 u0_u9_u4_U51 (.ZN( u0_u9_u4_n127 ) , .A( u0_u9_u4_n136 ) , .B2( u0_u9_u4_n150 ) , .B1( u0_u9_u4_n180 ) );
  INV_X1 u0_u9_u4_U52 (.A( u0_u9_u4_n160 ) , .ZN( u0_u9_u4_n180 ) );
  NAND2_X1 u0_u9_u4_U53 (.A2( u0_u9_u4_n104 ) , .A1( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n146 ) );
  NAND2_X1 u0_u9_u4_U54 (.A2( u0_u9_u4_n101 ) , .A1( u0_u9_u4_n102 ) , .ZN( u0_u9_u4_n160 ) );
  NAND2_X1 u0_u9_u4_U55 (.ZN( u0_u9_u4_n134 ) , .A1( u0_u9_u4_n98 ) , .A2( u0_u9_u4_n99 ) );
  NAND2_X1 u0_u9_u4_U56 (.A1( u0_u9_u4_n103 ) , .A2( u0_u9_u4_n104 ) , .ZN( u0_u9_u4_n143 ) );
  NAND2_X1 u0_u9_u4_U57 (.A2( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n145 ) , .A1( u0_u9_u4_n98 ) );
  NAND2_X1 u0_u9_u4_U58 (.A1( u0_u9_u4_n100 ) , .A2( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n120 ) );
  NAND2_X1 u0_u9_u4_U59 (.A1( u0_u9_u4_n102 ) , .A2( u0_u9_u4_n104 ) , .ZN( u0_u9_u4_n148 ) );
  AOI21_X1 u0_u9_u4_U6 (.ZN( u0_u9_u4_n106 ) , .B2( u0_u9_u4_n146 ) , .B1( u0_u9_u4_n158 ) , .A( u0_u9_u4_n170 ) );
  NAND2_X1 u0_u9_u4_U60 (.A2( u0_u9_u4_n100 ) , .A1( u0_u9_u4_n103 ) , .ZN( u0_u9_u4_n157 ) );
  INV_X1 u0_u9_u4_U61 (.A( u0_u9_u4_n150 ) , .ZN( u0_u9_u4_n173 ) );
  INV_X1 u0_u9_u4_U62 (.A( u0_u9_u4_n152 ) , .ZN( u0_u9_u4_n171 ) );
  NAND2_X1 u0_u9_u4_U63 (.A1( u0_u9_u4_n100 ) , .ZN( u0_u9_u4_n118 ) , .A2( u0_u9_u4_n99 ) );
  NAND2_X1 u0_u9_u4_U64 (.A2( u0_u9_u4_n100 ) , .A1( u0_u9_u4_n102 ) , .ZN( u0_u9_u4_n144 ) );
  NAND2_X1 u0_u9_u4_U65 (.A2( u0_u9_u4_n101 ) , .A1( u0_u9_u4_n105 ) , .ZN( u0_u9_u4_n96 ) );
  INV_X1 u0_u9_u4_U66 (.A( u0_u9_u4_n128 ) , .ZN( u0_u9_u4_n174 ) );
  NAND2_X1 u0_u9_u4_U67 (.A2( u0_u9_u4_n102 ) , .ZN( u0_u9_u4_n119 ) , .A1( u0_u9_u4_n98 ) );
  NAND2_X1 u0_u9_u4_U68 (.A2( u0_u9_u4_n101 ) , .A1( u0_u9_u4_n103 ) , .ZN( u0_u9_u4_n147 ) );
  NAND2_X1 u0_u9_u4_U69 (.A2( u0_u9_u4_n104 ) , .ZN( u0_u9_u4_n113 ) , .A1( u0_u9_u4_n99 ) );
  AOI21_X1 u0_u9_u4_U7 (.ZN( u0_u9_u4_n108 ) , .B2( u0_u9_u4_n134 ) , .B1( u0_u9_u4_n155 ) , .A( u0_u9_u4_n156 ) );
  NOR2_X1 u0_u9_u4_U70 (.A2( u0_u9_X_28 ) , .ZN( u0_u9_u4_n150 ) , .A1( u0_u9_u4_n168 ) );
  NOR2_X1 u0_u9_u4_U71 (.A2( u0_u9_X_29 ) , .ZN( u0_u9_u4_n152 ) , .A1( u0_u9_u4_n169 ) );
  NOR2_X1 u0_u9_u4_U72 (.A2( u0_u9_X_30 ) , .ZN( u0_u9_u4_n105 ) , .A1( u0_u9_u4_n176 ) );
  NOR2_X1 u0_u9_u4_U73 (.A2( u0_u9_X_26 ) , .ZN( u0_u9_u4_n100 ) , .A1( u0_u9_u4_n177 ) );
  NOR2_X1 u0_u9_u4_U74 (.A2( u0_u9_X_28 ) , .A1( u0_u9_X_29 ) , .ZN( u0_u9_u4_n128 ) );
  NOR2_X1 u0_u9_u4_U75 (.A2( u0_u9_X_27 ) , .A1( u0_u9_X_30 ) , .ZN( u0_u9_u4_n102 ) );
  NOR2_X1 u0_u9_u4_U76 (.A2( u0_u9_X_25 ) , .A1( u0_u9_X_26 ) , .ZN( u0_u9_u4_n98 ) );
  AND2_X1 u0_u9_u4_U77 (.A2( u0_u9_X_25 ) , .A1( u0_u9_X_26 ) , .ZN( u0_u9_u4_n104 ) );
  AND2_X1 u0_u9_u4_U78 (.A1( u0_u9_X_30 ) , .A2( u0_u9_u4_n176 ) , .ZN( u0_u9_u4_n99 ) );
  AND2_X1 u0_u9_u4_U79 (.A1( u0_u9_X_26 ) , .ZN( u0_u9_u4_n101 ) , .A2( u0_u9_u4_n177 ) );
  AOI21_X1 u0_u9_u4_U8 (.ZN( u0_u9_u4_n109 ) , .A( u0_u9_u4_n153 ) , .B1( u0_u9_u4_n159 ) , .B2( u0_u9_u4_n184 ) );
  AND2_X1 u0_u9_u4_U80 (.A1( u0_u9_X_27 ) , .A2( u0_u9_X_30 ) , .ZN( u0_u9_u4_n103 ) );
  INV_X1 u0_u9_u4_U81 (.A( u0_u9_X_28 ) , .ZN( u0_u9_u4_n169 ) );
  INV_X1 u0_u9_u4_U82 (.A( u0_u9_X_29 ) , .ZN( u0_u9_u4_n168 ) );
  INV_X1 u0_u9_u4_U83 (.A( u0_u9_X_25 ) , .ZN( u0_u9_u4_n177 ) );
  INV_X1 u0_u9_u4_U84 (.A( u0_u9_X_27 ) , .ZN( u0_u9_u4_n176 ) );
  NAND4_X1 u0_u9_u4_U85 (.ZN( u0_out9_25 ) , .A4( u0_u9_u4_n139 ) , .A3( u0_u9_u4_n140 ) , .A2( u0_u9_u4_n141 ) , .A1( u0_u9_u4_n142 ) );
  OAI21_X1 u0_u9_u4_U86 (.A( u0_u9_u4_n128 ) , .B2( u0_u9_u4_n129 ) , .B1( u0_u9_u4_n130 ) , .ZN( u0_u9_u4_n142 ) );
  OAI21_X1 u0_u9_u4_U87 (.B2( u0_u9_u4_n131 ) , .ZN( u0_u9_u4_n141 ) , .A( u0_u9_u4_n175 ) , .B1( u0_u9_u4_n183 ) );
  NAND4_X1 u0_u9_u4_U88 (.ZN( u0_out9_14 ) , .A4( u0_u9_u4_n124 ) , .A3( u0_u9_u4_n125 ) , .A2( u0_u9_u4_n126 ) , .A1( u0_u9_u4_n127 ) );
  AOI22_X1 u0_u9_u4_U89 (.B2( u0_u9_u4_n117 ) , .ZN( u0_u9_u4_n126 ) , .A1( u0_u9_u4_n129 ) , .B1( u0_u9_u4_n152 ) , .A2( u0_u9_u4_n175 ) );
  AOI211_X1 u0_u9_u4_U9 (.B( u0_u9_u4_n136 ) , .A( u0_u9_u4_n137 ) , .C2( u0_u9_u4_n138 ) , .ZN( u0_u9_u4_n139 ) , .C1( u0_u9_u4_n182 ) );
  AOI22_X1 u0_u9_u4_U90 (.ZN( u0_u9_u4_n125 ) , .B2( u0_u9_u4_n131 ) , .A2( u0_u9_u4_n132 ) , .B1( u0_u9_u4_n138 ) , .A1( u0_u9_u4_n178 ) );
  NAND4_X1 u0_u9_u4_U91 (.ZN( u0_out9_8 ) , .A4( u0_u9_u4_n110 ) , .A3( u0_u9_u4_n111 ) , .A2( u0_u9_u4_n112 ) , .A1( u0_u9_u4_n186 ) );
  NAND2_X1 u0_u9_u4_U92 (.ZN( u0_u9_u4_n112 ) , .A2( u0_u9_u4_n130 ) , .A1( u0_u9_u4_n150 ) );
  AOI22_X1 u0_u9_u4_U93 (.ZN( u0_u9_u4_n111 ) , .B2( u0_u9_u4_n132 ) , .A1( u0_u9_u4_n152 ) , .B1( u0_u9_u4_n178 ) , .A2( u0_u9_u4_n97 ) );
  AOI22_X1 u0_u9_u4_U94 (.B2( u0_u9_u4_n149 ) , .B1( u0_u9_u4_n150 ) , .A2( u0_u9_u4_n151 ) , .A1( u0_u9_u4_n152 ) , .ZN( u0_u9_u4_n167 ) );
  NOR4_X1 u0_u9_u4_U95 (.A4( u0_u9_u4_n162 ) , .A3( u0_u9_u4_n163 ) , .A2( u0_u9_u4_n164 ) , .A1( u0_u9_u4_n165 ) , .ZN( u0_u9_u4_n166 ) );
  NAND3_X1 u0_u9_u4_U96 (.ZN( u0_out9_3 ) , .A3( u0_u9_u4_n166 ) , .A1( u0_u9_u4_n167 ) , .A2( u0_u9_u4_n186 ) );
  NAND3_X1 u0_u9_u4_U97 (.A3( u0_u9_u4_n146 ) , .A2( u0_u9_u4_n147 ) , .A1( u0_u9_u4_n148 ) , .ZN( u0_u9_u4_n149 ) );
  NAND3_X1 u0_u9_u4_U98 (.A3( u0_u9_u4_n143 ) , .A2( u0_u9_u4_n144 ) , .A1( u0_u9_u4_n145 ) , .ZN( u0_u9_u4_n151 ) );
  NAND3_X1 u0_u9_u4_U99 (.A3( u0_u9_u4_n121 ) , .ZN( u0_u9_u4_n122 ) , .A2( u0_u9_u4_n144 ) , .A1( u0_u9_u4_n154 ) );
  NOR2_X1 u0_u9_u5_U10 (.ZN( u0_u9_u5_n135 ) , .A1( u0_u9_u5_n173 ) , .A2( u0_u9_u5_n176 ) );
  NOR3_X1 u0_u9_u5_U100 (.A3( u0_u9_u5_n141 ) , .A1( u0_u9_u5_n142 ) , .ZN( u0_u9_u5_n143 ) , .A2( u0_u9_u5_n191 ) );
  NAND4_X1 u0_u9_u5_U101 (.ZN( u0_out9_4 ) , .A4( u0_u9_u5_n112 ) , .A2( u0_u9_u5_n113 ) , .A1( u0_u9_u5_n114 ) , .A3( u0_u9_u5_n195 ) );
  AOI211_X1 u0_u9_u5_U102 (.A( u0_u9_u5_n110 ) , .C1( u0_u9_u5_n111 ) , .ZN( u0_u9_u5_n112 ) , .B( u0_u9_u5_n118 ) , .C2( u0_u9_u5_n177 ) );
  INV_X1 u0_u9_u5_U103 (.A( u0_u9_u5_n102 ) , .ZN( u0_u9_u5_n195 ) );
  NAND3_X1 u0_u9_u5_U104 (.A2( u0_u9_u5_n154 ) , .A3( u0_u9_u5_n158 ) , .A1( u0_u9_u5_n161 ) , .ZN( u0_u9_u5_n99 ) );
  INV_X1 u0_u9_u5_U11 (.A( u0_u9_u5_n121 ) , .ZN( u0_u9_u5_n177 ) );
  NOR2_X1 u0_u9_u5_U12 (.ZN( u0_u9_u5_n160 ) , .A2( u0_u9_u5_n173 ) , .A1( u0_u9_u5_n177 ) );
  INV_X1 u0_u9_u5_U13 (.A( u0_u9_u5_n150 ) , .ZN( u0_u9_u5_n174 ) );
  AOI21_X1 u0_u9_u5_U14 (.A( u0_u9_u5_n160 ) , .B2( u0_u9_u5_n161 ) , .ZN( u0_u9_u5_n162 ) , .B1( u0_u9_u5_n192 ) );
  INV_X1 u0_u9_u5_U15 (.A( u0_u9_u5_n159 ) , .ZN( u0_u9_u5_n192 ) );
  AOI21_X1 u0_u9_u5_U16 (.A( u0_u9_u5_n156 ) , .B2( u0_u9_u5_n157 ) , .B1( u0_u9_u5_n158 ) , .ZN( u0_u9_u5_n163 ) );
  AOI21_X1 u0_u9_u5_U17 (.B2( u0_u9_u5_n139 ) , .B1( u0_u9_u5_n140 ) , .ZN( u0_u9_u5_n141 ) , .A( u0_u9_u5_n150 ) );
  OAI21_X1 u0_u9_u5_U18 (.A( u0_u9_u5_n133 ) , .B2( u0_u9_u5_n134 ) , .B1( u0_u9_u5_n135 ) , .ZN( u0_u9_u5_n142 ) );
  OAI21_X1 u0_u9_u5_U19 (.ZN( u0_u9_u5_n133 ) , .B2( u0_u9_u5_n147 ) , .A( u0_u9_u5_n173 ) , .B1( u0_u9_u5_n188 ) );
  NAND2_X1 u0_u9_u5_U20 (.A2( u0_u9_u5_n119 ) , .A1( u0_u9_u5_n123 ) , .ZN( u0_u9_u5_n137 ) );
  INV_X1 u0_u9_u5_U21 (.A( u0_u9_u5_n155 ) , .ZN( u0_u9_u5_n194 ) );
  NAND2_X1 u0_u9_u5_U22 (.A1( u0_u9_u5_n121 ) , .ZN( u0_u9_u5_n132 ) , .A2( u0_u9_u5_n172 ) );
  NAND2_X1 u0_u9_u5_U23 (.A2( u0_u9_u5_n122 ) , .ZN( u0_u9_u5_n136 ) , .A1( u0_u9_u5_n154 ) );
  NAND2_X1 u0_u9_u5_U24 (.A2( u0_u9_u5_n119 ) , .A1( u0_u9_u5_n120 ) , .ZN( u0_u9_u5_n159 ) );
  INV_X1 u0_u9_u5_U25 (.A( u0_u9_u5_n156 ) , .ZN( u0_u9_u5_n175 ) );
  INV_X1 u0_u9_u5_U26 (.A( u0_u9_u5_n158 ) , .ZN( u0_u9_u5_n188 ) );
  INV_X1 u0_u9_u5_U27 (.A( u0_u9_u5_n152 ) , .ZN( u0_u9_u5_n179 ) );
  INV_X1 u0_u9_u5_U28 (.A( u0_u9_u5_n140 ) , .ZN( u0_u9_u5_n182 ) );
  INV_X1 u0_u9_u5_U29 (.A( u0_u9_u5_n151 ) , .ZN( u0_u9_u5_n183 ) );
  NOR2_X1 u0_u9_u5_U3 (.ZN( u0_u9_u5_n134 ) , .A1( u0_u9_u5_n183 ) , .A2( u0_u9_u5_n190 ) );
  INV_X1 u0_u9_u5_U30 (.A( u0_u9_u5_n123 ) , .ZN( u0_u9_u5_n185 ) );
  INV_X1 u0_u9_u5_U31 (.A( u0_u9_u5_n161 ) , .ZN( u0_u9_u5_n184 ) );
  INV_X1 u0_u9_u5_U32 (.A( u0_u9_u5_n139 ) , .ZN( u0_u9_u5_n189 ) );
  INV_X1 u0_u9_u5_U33 (.A( u0_u9_u5_n157 ) , .ZN( u0_u9_u5_n190 ) );
  INV_X1 u0_u9_u5_U34 (.A( u0_u9_u5_n120 ) , .ZN( u0_u9_u5_n193 ) );
  NAND2_X1 u0_u9_u5_U35 (.ZN( u0_u9_u5_n111 ) , .A1( u0_u9_u5_n140 ) , .A2( u0_u9_u5_n155 ) );
  NOR2_X1 u0_u9_u5_U36 (.ZN( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n170 ) , .A2( u0_u9_u5_n180 ) );
  INV_X1 u0_u9_u5_U37 (.A( u0_u9_u5_n117 ) , .ZN( u0_u9_u5_n196 ) );
  OAI221_X1 u0_u9_u5_U38 (.A( u0_u9_u5_n116 ) , .ZN( u0_u9_u5_n117 ) , .B2( u0_u9_u5_n119 ) , .C1( u0_u9_u5_n153 ) , .C2( u0_u9_u5_n158 ) , .B1( u0_u9_u5_n172 ) );
  AOI222_X1 u0_u9_u5_U39 (.ZN( u0_u9_u5_n116 ) , .B2( u0_u9_u5_n145 ) , .C1( u0_u9_u5_n148 ) , .A2( u0_u9_u5_n174 ) , .C2( u0_u9_u5_n177 ) , .B1( u0_u9_u5_n187 ) , .A1( u0_u9_u5_n193 ) );
  INV_X1 u0_u9_u5_U4 (.A( u0_u9_u5_n138 ) , .ZN( u0_u9_u5_n191 ) );
  INV_X1 u0_u9_u5_U40 (.A( u0_u9_u5_n115 ) , .ZN( u0_u9_u5_n187 ) );
  OAI221_X1 u0_u9_u5_U41 (.A( u0_u9_u5_n101 ) , .ZN( u0_u9_u5_n102 ) , .C2( u0_u9_u5_n115 ) , .C1( u0_u9_u5_n126 ) , .B1( u0_u9_u5_n134 ) , .B2( u0_u9_u5_n160 ) );
  OAI21_X1 u0_u9_u5_U42 (.ZN( u0_u9_u5_n101 ) , .B1( u0_u9_u5_n137 ) , .A( u0_u9_u5_n146 ) , .B2( u0_u9_u5_n147 ) );
  AOI22_X1 u0_u9_u5_U43 (.B2( u0_u9_u5_n131 ) , .A2( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n169 ) , .B1( u0_u9_u5_n174 ) , .A1( u0_u9_u5_n185 ) );
  NOR2_X1 u0_u9_u5_U44 (.A1( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n150 ) , .A2( u0_u9_u5_n173 ) );
  AOI21_X1 u0_u9_u5_U45 (.A( u0_u9_u5_n118 ) , .B2( u0_u9_u5_n145 ) , .ZN( u0_u9_u5_n168 ) , .B1( u0_u9_u5_n186 ) );
  INV_X1 u0_u9_u5_U46 (.A( u0_u9_u5_n122 ) , .ZN( u0_u9_u5_n186 ) );
  NOR2_X1 u0_u9_u5_U47 (.A1( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n152 ) , .A2( u0_u9_u5_n176 ) );
  NOR2_X1 u0_u9_u5_U48 (.A1( u0_u9_u5_n115 ) , .ZN( u0_u9_u5_n118 ) , .A2( u0_u9_u5_n153 ) );
  NOR2_X1 u0_u9_u5_U49 (.A2( u0_u9_u5_n145 ) , .ZN( u0_u9_u5_n156 ) , .A1( u0_u9_u5_n174 ) );
  OAI21_X1 u0_u9_u5_U5 (.B2( u0_u9_u5_n136 ) , .B1( u0_u9_u5_n137 ) , .ZN( u0_u9_u5_n138 ) , .A( u0_u9_u5_n177 ) );
  NOR2_X1 u0_u9_u5_U50 (.ZN( u0_u9_u5_n121 ) , .A2( u0_u9_u5_n145 ) , .A1( u0_u9_u5_n176 ) );
  AOI22_X1 u0_u9_u5_U51 (.ZN( u0_u9_u5_n114 ) , .A2( u0_u9_u5_n137 ) , .A1( u0_u9_u5_n145 ) , .B2( u0_u9_u5_n175 ) , .B1( u0_u9_u5_n193 ) );
  OAI211_X1 u0_u9_u5_U52 (.B( u0_u9_u5_n124 ) , .A( u0_u9_u5_n125 ) , .C2( u0_u9_u5_n126 ) , .C1( u0_u9_u5_n127 ) , .ZN( u0_u9_u5_n128 ) );
  NOR3_X1 u0_u9_u5_U53 (.ZN( u0_u9_u5_n127 ) , .A1( u0_u9_u5_n136 ) , .A3( u0_u9_u5_n148 ) , .A2( u0_u9_u5_n182 ) );
  OAI21_X1 u0_u9_u5_U54 (.ZN( u0_u9_u5_n124 ) , .A( u0_u9_u5_n177 ) , .B2( u0_u9_u5_n183 ) , .B1( u0_u9_u5_n189 ) );
  OAI21_X1 u0_u9_u5_U55 (.ZN( u0_u9_u5_n125 ) , .A( u0_u9_u5_n174 ) , .B2( u0_u9_u5_n185 ) , .B1( u0_u9_u5_n190 ) );
  AOI21_X1 u0_u9_u5_U56 (.A( u0_u9_u5_n153 ) , .B2( u0_u9_u5_n154 ) , .B1( u0_u9_u5_n155 ) , .ZN( u0_u9_u5_n164 ) );
  AOI21_X1 u0_u9_u5_U57 (.ZN( u0_u9_u5_n110 ) , .B1( u0_u9_u5_n122 ) , .B2( u0_u9_u5_n139 ) , .A( u0_u9_u5_n153 ) );
  INV_X1 u0_u9_u5_U58 (.A( u0_u9_u5_n153 ) , .ZN( u0_u9_u5_n176 ) );
  INV_X1 u0_u9_u5_U59 (.A( u0_u9_u5_n126 ) , .ZN( u0_u9_u5_n173 ) );
  AOI222_X1 u0_u9_u5_U6 (.ZN( u0_u9_u5_n113 ) , .A1( u0_u9_u5_n131 ) , .C1( u0_u9_u5_n148 ) , .B2( u0_u9_u5_n174 ) , .C2( u0_u9_u5_n178 ) , .A2( u0_u9_u5_n179 ) , .B1( u0_u9_u5_n99 ) );
  AND2_X1 u0_u9_u5_U60 (.A2( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n107 ) , .ZN( u0_u9_u5_n147 ) );
  AND2_X1 u0_u9_u5_U61 (.A2( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n108 ) , .ZN( u0_u9_u5_n148 ) );
  NAND2_X1 u0_u9_u5_U62 (.A1( u0_u9_u5_n105 ) , .A2( u0_u9_u5_n106 ) , .ZN( u0_u9_u5_n158 ) );
  NAND2_X1 u0_u9_u5_U63 (.A2( u0_u9_u5_n108 ) , .A1( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n139 ) );
  NAND2_X1 u0_u9_u5_U64 (.A1( u0_u9_u5_n106 ) , .A2( u0_u9_u5_n108 ) , .ZN( u0_u9_u5_n119 ) );
  NAND2_X1 u0_u9_u5_U65 (.A2( u0_u9_u5_n103 ) , .A1( u0_u9_u5_n105 ) , .ZN( u0_u9_u5_n140 ) );
  NAND2_X1 u0_u9_u5_U66 (.A2( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n105 ) , .ZN( u0_u9_u5_n155 ) );
  NAND2_X1 u0_u9_u5_U67 (.A2( u0_u9_u5_n106 ) , .A1( u0_u9_u5_n107 ) , .ZN( u0_u9_u5_n122 ) );
  NAND2_X1 u0_u9_u5_U68 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n106 ) , .ZN( u0_u9_u5_n115 ) );
  NAND2_X1 u0_u9_u5_U69 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n103 ) , .ZN( u0_u9_u5_n161 ) );
  INV_X1 u0_u9_u5_U7 (.A( u0_u9_u5_n135 ) , .ZN( u0_u9_u5_n178 ) );
  NAND2_X1 u0_u9_u5_U70 (.A1( u0_u9_u5_n105 ) , .A2( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n154 ) );
  INV_X1 u0_u9_u5_U71 (.A( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n172 ) );
  NAND2_X1 u0_u9_u5_U72 (.A1( u0_u9_u5_n103 ) , .A2( u0_u9_u5_n108 ) , .ZN( u0_u9_u5_n123 ) );
  NAND2_X1 u0_u9_u5_U73 (.A2( u0_u9_u5_n103 ) , .A1( u0_u9_u5_n107 ) , .ZN( u0_u9_u5_n151 ) );
  NAND2_X1 u0_u9_u5_U74 (.A2( u0_u9_u5_n107 ) , .A1( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n120 ) );
  NAND2_X1 u0_u9_u5_U75 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n109 ) , .ZN( u0_u9_u5_n157 ) );
  AND2_X1 u0_u9_u5_U76 (.A2( u0_u9_u5_n100 ) , .A1( u0_u9_u5_n104 ) , .ZN( u0_u9_u5_n131 ) );
  NOR2_X1 u0_u9_u5_U77 (.A2( u0_u9_X_34 ) , .A1( u0_u9_X_35 ) , .ZN( u0_u9_u5_n145 ) );
  NOR2_X1 u0_u9_u5_U78 (.A2( u0_u9_X_34 ) , .ZN( u0_u9_u5_n146 ) , .A1( u0_u9_u5_n171 ) );
  NOR2_X1 u0_u9_u5_U79 (.A2( u0_u9_X_31 ) , .A1( u0_u9_X_32 ) , .ZN( u0_u9_u5_n103 ) );
  OAI22_X1 u0_u9_u5_U8 (.B2( u0_u9_u5_n149 ) , .B1( u0_u9_u5_n150 ) , .A2( u0_u9_u5_n151 ) , .A1( u0_u9_u5_n152 ) , .ZN( u0_u9_u5_n165 ) );
  NOR2_X1 u0_u9_u5_U80 (.A2( u0_u9_X_36 ) , .ZN( u0_u9_u5_n105 ) , .A1( u0_u9_u5_n180 ) );
  NOR2_X1 u0_u9_u5_U81 (.A2( u0_u9_X_33 ) , .ZN( u0_u9_u5_n108 ) , .A1( u0_u9_u5_n170 ) );
  NOR2_X1 u0_u9_u5_U82 (.A2( u0_u9_X_33 ) , .A1( u0_u9_X_36 ) , .ZN( u0_u9_u5_n107 ) );
  NOR2_X1 u0_u9_u5_U83 (.A2( u0_u9_X_31 ) , .ZN( u0_u9_u5_n104 ) , .A1( u0_u9_u5_n181 ) );
  NAND2_X1 u0_u9_u5_U84 (.A2( u0_u9_X_34 ) , .A1( u0_u9_X_35 ) , .ZN( u0_u9_u5_n153 ) );
  NAND2_X1 u0_u9_u5_U85 (.A1( u0_u9_X_34 ) , .ZN( u0_u9_u5_n126 ) , .A2( u0_u9_u5_n171 ) );
  AND2_X1 u0_u9_u5_U86 (.A1( u0_u9_X_31 ) , .A2( u0_u9_X_32 ) , .ZN( u0_u9_u5_n106 ) );
  AND2_X1 u0_u9_u5_U87 (.A1( u0_u9_X_31 ) , .ZN( u0_u9_u5_n109 ) , .A2( u0_u9_u5_n181 ) );
  INV_X1 u0_u9_u5_U88 (.A( u0_u9_X_33 ) , .ZN( u0_u9_u5_n180 ) );
  INV_X1 u0_u9_u5_U89 (.A( u0_u9_X_35 ) , .ZN( u0_u9_u5_n171 ) );
  NOR3_X1 u0_u9_u5_U9 (.A2( u0_u9_u5_n147 ) , .A1( u0_u9_u5_n148 ) , .ZN( u0_u9_u5_n149 ) , .A3( u0_u9_u5_n194 ) );
  INV_X1 u0_u9_u5_U90 (.A( u0_u9_X_36 ) , .ZN( u0_u9_u5_n170 ) );
  INV_X1 u0_u9_u5_U91 (.A( u0_u9_X_32 ) , .ZN( u0_u9_u5_n181 ) );
  NAND4_X1 u0_u9_u5_U92 (.ZN( u0_out9_29 ) , .A4( u0_u9_u5_n129 ) , .A3( u0_u9_u5_n130 ) , .A2( u0_u9_u5_n168 ) , .A1( u0_u9_u5_n196 ) );
  AOI221_X1 u0_u9_u5_U93 (.A( u0_u9_u5_n128 ) , .ZN( u0_u9_u5_n129 ) , .C2( u0_u9_u5_n132 ) , .B2( u0_u9_u5_n159 ) , .B1( u0_u9_u5_n176 ) , .C1( u0_u9_u5_n184 ) );
  AOI222_X1 u0_u9_u5_U94 (.ZN( u0_u9_u5_n130 ) , .A2( u0_u9_u5_n146 ) , .B1( u0_u9_u5_n147 ) , .C2( u0_u9_u5_n175 ) , .B2( u0_u9_u5_n179 ) , .A1( u0_u9_u5_n188 ) , .C1( u0_u9_u5_n194 ) );
  NAND4_X1 u0_u9_u5_U95 (.ZN( u0_out9_19 ) , .A4( u0_u9_u5_n166 ) , .A3( u0_u9_u5_n167 ) , .A2( u0_u9_u5_n168 ) , .A1( u0_u9_u5_n169 ) );
  AOI22_X1 u0_u9_u5_U96 (.B2( u0_u9_u5_n145 ) , .A2( u0_u9_u5_n146 ) , .ZN( u0_u9_u5_n167 ) , .B1( u0_u9_u5_n182 ) , .A1( u0_u9_u5_n189 ) );
  NOR4_X1 u0_u9_u5_U97 (.A4( u0_u9_u5_n162 ) , .A3( u0_u9_u5_n163 ) , .A2( u0_u9_u5_n164 ) , .A1( u0_u9_u5_n165 ) , .ZN( u0_u9_u5_n166 ) );
  NAND4_X1 u0_u9_u5_U98 (.ZN( u0_out9_11 ) , .A4( u0_u9_u5_n143 ) , .A3( u0_u9_u5_n144 ) , .A2( u0_u9_u5_n169 ) , .A1( u0_u9_u5_n196 ) );
  AOI22_X1 u0_u9_u5_U99 (.A2( u0_u9_u5_n132 ) , .ZN( u0_u9_u5_n144 ) , .B2( u0_u9_u5_n145 ) , .B1( u0_u9_u5_n184 ) , .A1( u0_u9_u5_n194 ) );
  AND3_X1 u0_u9_u7_U10 (.A3( u0_u9_u7_n110 ) , .A2( u0_u9_u7_n127 ) , .A1( u0_u9_u7_n132 ) , .ZN( u0_u9_u7_n92 ) );
  OAI21_X1 u0_u9_u7_U11 (.A( u0_u9_u7_n161 ) , .B1( u0_u9_u7_n168 ) , .B2( u0_u9_u7_n173 ) , .ZN( u0_u9_u7_n91 ) );
  AOI211_X1 u0_u9_u7_U12 (.A( u0_u9_u7_n117 ) , .ZN( u0_u9_u7_n118 ) , .C2( u0_u9_u7_n126 ) , .C1( u0_u9_u7_n177 ) , .B( u0_u9_u7_n180 ) );
  OAI22_X1 u0_u9_u7_U13 (.B1( u0_u9_u7_n115 ) , .ZN( u0_u9_u7_n117 ) , .A2( u0_u9_u7_n133 ) , .A1( u0_u9_u7_n137 ) , .B2( u0_u9_u7_n162 ) );
  INV_X1 u0_u9_u7_U14 (.A( u0_u9_u7_n116 ) , .ZN( u0_u9_u7_n180 ) );
  NOR3_X1 u0_u9_u7_U15 (.ZN( u0_u9_u7_n115 ) , .A3( u0_u9_u7_n145 ) , .A2( u0_u9_u7_n168 ) , .A1( u0_u9_u7_n169 ) );
  OAI211_X1 u0_u9_u7_U16 (.B( u0_u9_u7_n122 ) , .A( u0_u9_u7_n123 ) , .C2( u0_u9_u7_n124 ) , .ZN( u0_u9_u7_n154 ) , .C1( u0_u9_u7_n162 ) );
  AOI222_X1 u0_u9_u7_U17 (.ZN( u0_u9_u7_n122 ) , .C2( u0_u9_u7_n126 ) , .C1( u0_u9_u7_n145 ) , .B1( u0_u9_u7_n161 ) , .A2( u0_u9_u7_n165 ) , .B2( u0_u9_u7_n170 ) , .A1( u0_u9_u7_n176 ) );
  INV_X1 u0_u9_u7_U18 (.A( u0_u9_u7_n133 ) , .ZN( u0_u9_u7_n176 ) );
  NOR3_X1 u0_u9_u7_U19 (.A2( u0_u9_u7_n134 ) , .A1( u0_u9_u7_n135 ) , .ZN( u0_u9_u7_n136 ) , .A3( u0_u9_u7_n171 ) );
  NOR2_X1 u0_u9_u7_U20 (.A1( u0_u9_u7_n130 ) , .A2( u0_u9_u7_n134 ) , .ZN( u0_u9_u7_n153 ) );
  INV_X1 u0_u9_u7_U21 (.A( u0_u9_u7_n101 ) , .ZN( u0_u9_u7_n165 ) );
  NOR2_X1 u0_u9_u7_U22 (.ZN( u0_u9_u7_n111 ) , .A2( u0_u9_u7_n134 ) , .A1( u0_u9_u7_n169 ) );
  AOI21_X1 u0_u9_u7_U23 (.ZN( u0_u9_u7_n104 ) , .B2( u0_u9_u7_n112 ) , .B1( u0_u9_u7_n127 ) , .A( u0_u9_u7_n164 ) );
  AOI21_X1 u0_u9_u7_U24 (.ZN( u0_u9_u7_n106 ) , .B1( u0_u9_u7_n133 ) , .B2( u0_u9_u7_n146 ) , .A( u0_u9_u7_n162 ) );
  AOI21_X1 u0_u9_u7_U25 (.A( u0_u9_u7_n101 ) , .ZN( u0_u9_u7_n107 ) , .B2( u0_u9_u7_n128 ) , .B1( u0_u9_u7_n175 ) );
  INV_X1 u0_u9_u7_U26 (.A( u0_u9_u7_n138 ) , .ZN( u0_u9_u7_n171 ) );
  INV_X1 u0_u9_u7_U27 (.A( u0_u9_u7_n131 ) , .ZN( u0_u9_u7_n177 ) );
  INV_X1 u0_u9_u7_U28 (.A( u0_u9_u7_n110 ) , .ZN( u0_u9_u7_n174 ) );
  NAND2_X1 u0_u9_u7_U29 (.A1( u0_u9_u7_n129 ) , .A2( u0_u9_u7_n132 ) , .ZN( u0_u9_u7_n149 ) );
  OAI21_X1 u0_u9_u7_U3 (.ZN( u0_u9_u7_n159 ) , .A( u0_u9_u7_n165 ) , .B2( u0_u9_u7_n171 ) , .B1( u0_u9_u7_n174 ) );
  NAND2_X1 u0_u9_u7_U30 (.A1( u0_u9_u7_n113 ) , .A2( u0_u9_u7_n124 ) , .ZN( u0_u9_u7_n130 ) );
  INV_X1 u0_u9_u7_U31 (.A( u0_u9_u7_n112 ) , .ZN( u0_u9_u7_n173 ) );
  INV_X1 u0_u9_u7_U32 (.A( u0_u9_u7_n128 ) , .ZN( u0_u9_u7_n168 ) );
  INV_X1 u0_u9_u7_U33 (.A( u0_u9_u7_n148 ) , .ZN( u0_u9_u7_n169 ) );
  INV_X1 u0_u9_u7_U34 (.A( u0_u9_u7_n127 ) , .ZN( u0_u9_u7_n179 ) );
  NOR2_X1 u0_u9_u7_U35 (.ZN( u0_u9_u7_n101 ) , .A2( u0_u9_u7_n150 ) , .A1( u0_u9_u7_n156 ) );
  AOI211_X1 u0_u9_u7_U36 (.B( u0_u9_u7_n154 ) , .A( u0_u9_u7_n155 ) , .C1( u0_u9_u7_n156 ) , .ZN( u0_u9_u7_n157 ) , .C2( u0_u9_u7_n172 ) );
  INV_X1 u0_u9_u7_U37 (.A( u0_u9_u7_n153 ) , .ZN( u0_u9_u7_n172 ) );
  AOI211_X1 u0_u9_u7_U38 (.B( u0_u9_u7_n139 ) , .A( u0_u9_u7_n140 ) , .C2( u0_u9_u7_n141 ) , .ZN( u0_u9_u7_n142 ) , .C1( u0_u9_u7_n156 ) );
  NAND4_X1 u0_u9_u7_U39 (.A3( u0_u9_u7_n127 ) , .A2( u0_u9_u7_n128 ) , .A1( u0_u9_u7_n129 ) , .ZN( u0_u9_u7_n141 ) , .A4( u0_u9_u7_n147 ) );
  INV_X1 u0_u9_u7_U4 (.A( u0_u9_u7_n111 ) , .ZN( u0_u9_u7_n170 ) );
  AOI21_X1 u0_u9_u7_U40 (.A( u0_u9_u7_n137 ) , .B1( u0_u9_u7_n138 ) , .ZN( u0_u9_u7_n139 ) , .B2( u0_u9_u7_n146 ) );
  OAI22_X1 u0_u9_u7_U41 (.B1( u0_u9_u7_n136 ) , .ZN( u0_u9_u7_n140 ) , .A1( u0_u9_u7_n153 ) , .B2( u0_u9_u7_n162 ) , .A2( u0_u9_u7_n164 ) );
  AOI21_X1 u0_u9_u7_U42 (.ZN( u0_u9_u7_n123 ) , .B1( u0_u9_u7_n165 ) , .B2( u0_u9_u7_n177 ) , .A( u0_u9_u7_n97 ) );
  AOI21_X1 u0_u9_u7_U43 (.B2( u0_u9_u7_n113 ) , .B1( u0_u9_u7_n124 ) , .A( u0_u9_u7_n125 ) , .ZN( u0_u9_u7_n97 ) );
  INV_X1 u0_u9_u7_U44 (.A( u0_u9_u7_n125 ) , .ZN( u0_u9_u7_n161 ) );
  INV_X1 u0_u9_u7_U45 (.A( u0_u9_u7_n152 ) , .ZN( u0_u9_u7_n162 ) );
  AOI22_X1 u0_u9_u7_U46 (.A2( u0_u9_u7_n114 ) , .ZN( u0_u9_u7_n119 ) , .B1( u0_u9_u7_n130 ) , .A1( u0_u9_u7_n156 ) , .B2( u0_u9_u7_n165 ) );
  NAND2_X1 u0_u9_u7_U47 (.A2( u0_u9_u7_n112 ) , .ZN( u0_u9_u7_n114 ) , .A1( u0_u9_u7_n175 ) );
  AND2_X1 u0_u9_u7_U48 (.ZN( u0_u9_u7_n145 ) , .A2( u0_u9_u7_n98 ) , .A1( u0_u9_u7_n99 ) );
  NOR2_X1 u0_u9_u7_U49 (.ZN( u0_u9_u7_n137 ) , .A1( u0_u9_u7_n150 ) , .A2( u0_u9_u7_n161 ) );
  INV_X1 u0_u9_u7_U5 (.A( u0_u9_u7_n149 ) , .ZN( u0_u9_u7_n175 ) );
  AOI21_X1 u0_u9_u7_U50 (.ZN( u0_u9_u7_n105 ) , .B2( u0_u9_u7_n110 ) , .A( u0_u9_u7_n125 ) , .B1( u0_u9_u7_n147 ) );
  NAND2_X1 u0_u9_u7_U51 (.ZN( u0_u9_u7_n146 ) , .A1( u0_u9_u7_n95 ) , .A2( u0_u9_u7_n98 ) );
  NAND2_X1 u0_u9_u7_U52 (.A2( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n147 ) , .A1( u0_u9_u7_n93 ) );
  NAND2_X1 u0_u9_u7_U53 (.A1( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n127 ) , .A2( u0_u9_u7_n99 ) );
  OR2_X1 u0_u9_u7_U54 (.ZN( u0_u9_u7_n126 ) , .A2( u0_u9_u7_n152 ) , .A1( u0_u9_u7_n156 ) );
  NAND2_X1 u0_u9_u7_U55 (.A2( u0_u9_u7_n102 ) , .A1( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n133 ) );
  NAND2_X1 u0_u9_u7_U56 (.ZN( u0_u9_u7_n112 ) , .A2( u0_u9_u7_n96 ) , .A1( u0_u9_u7_n99 ) );
  NAND2_X1 u0_u9_u7_U57 (.A2( u0_u9_u7_n102 ) , .ZN( u0_u9_u7_n128 ) , .A1( u0_u9_u7_n98 ) );
  NAND2_X1 u0_u9_u7_U58 (.A1( u0_u9_u7_n100 ) , .ZN( u0_u9_u7_n113 ) , .A2( u0_u9_u7_n93 ) );
  NAND2_X1 u0_u9_u7_U59 (.A2( u0_u9_u7_n102 ) , .ZN( u0_u9_u7_n124 ) , .A1( u0_u9_u7_n96 ) );
  INV_X1 u0_u9_u7_U6 (.A( u0_u9_u7_n154 ) , .ZN( u0_u9_u7_n178 ) );
  NAND2_X1 u0_u9_u7_U60 (.ZN( u0_u9_u7_n110 ) , .A1( u0_u9_u7_n95 ) , .A2( u0_u9_u7_n96 ) );
  INV_X1 u0_u9_u7_U61 (.A( u0_u9_u7_n150 ) , .ZN( u0_u9_u7_n164 ) );
  AND2_X1 u0_u9_u7_U62 (.ZN( u0_u9_u7_n134 ) , .A1( u0_u9_u7_n93 ) , .A2( u0_u9_u7_n98 ) );
  NAND2_X1 u0_u9_u7_U63 (.A1( u0_u9_u7_n100 ) , .A2( u0_u9_u7_n102 ) , .ZN( u0_u9_u7_n129 ) );
  NAND2_X1 u0_u9_u7_U64 (.A2( u0_u9_u7_n103 ) , .ZN( u0_u9_u7_n131 ) , .A1( u0_u9_u7_n95 ) );
  NAND2_X1 u0_u9_u7_U65 (.A1( u0_u9_u7_n100 ) , .ZN( u0_u9_u7_n138 ) , .A2( u0_u9_u7_n99 ) );
  NAND2_X1 u0_u9_u7_U66 (.ZN( u0_u9_u7_n132 ) , .A1( u0_u9_u7_n93 ) , .A2( u0_u9_u7_n96 ) );
  NAND2_X1 u0_u9_u7_U67 (.A1( u0_u9_u7_n100 ) , .ZN( u0_u9_u7_n148 ) , .A2( u0_u9_u7_n95 ) );
  NOR2_X1 u0_u9_u7_U68 (.A2( u0_u9_X_47 ) , .ZN( u0_u9_u7_n150 ) , .A1( u0_u9_u7_n163 ) );
  NOR2_X1 u0_u9_u7_U69 (.A2( u0_u9_X_43 ) , .A1( u0_u9_X_44 ) , .ZN( u0_u9_u7_n103 ) );
  AOI211_X1 u0_u9_u7_U7 (.ZN( u0_u9_u7_n116 ) , .A( u0_u9_u7_n155 ) , .C1( u0_u9_u7_n161 ) , .C2( u0_u9_u7_n171 ) , .B( u0_u9_u7_n94 ) );
  NOR2_X1 u0_u9_u7_U70 (.A2( u0_u9_X_48 ) , .A1( u0_u9_u7_n166 ) , .ZN( u0_u9_u7_n95 ) );
  NOR2_X1 u0_u9_u7_U71 (.A2( u0_u9_X_45 ) , .A1( u0_u9_X_48 ) , .ZN( u0_u9_u7_n99 ) );
  NOR2_X1 u0_u9_u7_U72 (.A2( u0_u9_X_44 ) , .A1( u0_u9_u7_n167 ) , .ZN( u0_u9_u7_n98 ) );
  NOR2_X1 u0_u9_u7_U73 (.A2( u0_u9_X_46 ) , .A1( u0_u9_X_47 ) , .ZN( u0_u9_u7_n152 ) );
  AND2_X1 u0_u9_u7_U74 (.A1( u0_u9_X_47 ) , .ZN( u0_u9_u7_n156 ) , .A2( u0_u9_u7_n163 ) );
  NAND2_X1 u0_u9_u7_U75 (.A2( u0_u9_X_46 ) , .A1( u0_u9_X_47 ) , .ZN( u0_u9_u7_n125 ) );
  AND2_X1 u0_u9_u7_U76 (.A2( u0_u9_X_45 ) , .A1( u0_u9_X_48 ) , .ZN( u0_u9_u7_n102 ) );
  AND2_X1 u0_u9_u7_U77 (.A2( u0_u9_X_43 ) , .A1( u0_u9_X_44 ) , .ZN( u0_u9_u7_n96 ) );
  AND2_X1 u0_u9_u7_U78 (.A1( u0_u9_X_44 ) , .ZN( u0_u9_u7_n100 ) , .A2( u0_u9_u7_n167 ) );
  AND2_X1 u0_u9_u7_U79 (.A1( u0_u9_X_48 ) , .A2( u0_u9_u7_n166 ) , .ZN( u0_u9_u7_n93 ) );
  OAI222_X1 u0_u9_u7_U8 (.C2( u0_u9_u7_n101 ) , .B2( u0_u9_u7_n111 ) , .A1( u0_u9_u7_n113 ) , .C1( u0_u9_u7_n146 ) , .A2( u0_u9_u7_n162 ) , .B1( u0_u9_u7_n164 ) , .ZN( u0_u9_u7_n94 ) );
  INV_X1 u0_u9_u7_U80 (.A( u0_u9_X_46 ) , .ZN( u0_u9_u7_n163 ) );
  INV_X1 u0_u9_u7_U81 (.A( u0_u9_X_45 ) , .ZN( u0_u9_u7_n166 ) );
  INV_X1 u0_u9_u7_U82 (.A( u0_u9_X_43 ) , .ZN( u0_u9_u7_n167 ) );
  NAND4_X1 u0_u9_u7_U83 (.ZN( u0_out9_27 ) , .A4( u0_u9_u7_n118 ) , .A3( u0_u9_u7_n119 ) , .A2( u0_u9_u7_n120 ) , .A1( u0_u9_u7_n121 ) );
  OAI21_X1 u0_u9_u7_U84 (.ZN( u0_u9_u7_n121 ) , .B2( u0_u9_u7_n145 ) , .A( u0_u9_u7_n150 ) , .B1( u0_u9_u7_n174 ) );
  OAI21_X1 u0_u9_u7_U85 (.ZN( u0_u9_u7_n120 ) , .A( u0_u9_u7_n161 ) , .B2( u0_u9_u7_n170 ) , .B1( u0_u9_u7_n179 ) );
  NAND4_X1 u0_u9_u7_U86 (.ZN( u0_out9_21 ) , .A4( u0_u9_u7_n157 ) , .A3( u0_u9_u7_n158 ) , .A2( u0_u9_u7_n159 ) , .A1( u0_u9_u7_n160 ) );
  OAI21_X1 u0_u9_u7_U87 (.B1( u0_u9_u7_n145 ) , .ZN( u0_u9_u7_n160 ) , .A( u0_u9_u7_n161 ) , .B2( u0_u9_u7_n177 ) );
  AOI22_X1 u0_u9_u7_U88 (.B2( u0_u9_u7_n149 ) , .B1( u0_u9_u7_n150 ) , .A2( u0_u9_u7_n151 ) , .A1( u0_u9_u7_n152 ) , .ZN( u0_u9_u7_n158 ) );
  NAND4_X1 u0_u9_u7_U89 (.ZN( u0_out9_15 ) , .A4( u0_u9_u7_n142 ) , .A3( u0_u9_u7_n143 ) , .A2( u0_u9_u7_n144 ) , .A1( u0_u9_u7_n178 ) );
  OAI221_X1 u0_u9_u7_U9 (.C1( u0_u9_u7_n101 ) , .C2( u0_u9_u7_n147 ) , .ZN( u0_u9_u7_n155 ) , .B2( u0_u9_u7_n162 ) , .A( u0_u9_u7_n91 ) , .B1( u0_u9_u7_n92 ) );
  OR2_X1 u0_u9_u7_U90 (.A2( u0_u9_u7_n125 ) , .A1( u0_u9_u7_n129 ) , .ZN( u0_u9_u7_n144 ) );
  AOI22_X1 u0_u9_u7_U91 (.A2( u0_u9_u7_n126 ) , .ZN( u0_u9_u7_n143 ) , .B2( u0_u9_u7_n165 ) , .B1( u0_u9_u7_n173 ) , .A1( u0_u9_u7_n174 ) );
  NAND4_X1 u0_u9_u7_U92 (.ZN( u0_out9_5 ) , .A4( u0_u9_u7_n108 ) , .A3( u0_u9_u7_n109 ) , .A1( u0_u9_u7_n116 ) , .A2( u0_u9_u7_n123 ) );
  AOI22_X1 u0_u9_u7_U93 (.ZN( u0_u9_u7_n109 ) , .A2( u0_u9_u7_n126 ) , .B2( u0_u9_u7_n145 ) , .B1( u0_u9_u7_n156 ) , .A1( u0_u9_u7_n171 ) );
  NOR4_X1 u0_u9_u7_U94 (.A4( u0_u9_u7_n104 ) , .A3( u0_u9_u7_n105 ) , .A2( u0_u9_u7_n106 ) , .A1( u0_u9_u7_n107 ) , .ZN( u0_u9_u7_n108 ) );
  NAND3_X1 u0_u9_u7_U95 (.A3( u0_u9_u7_n146 ) , .A2( u0_u9_u7_n147 ) , .A1( u0_u9_u7_n148 ) , .ZN( u0_u9_u7_n151 ) );
  NAND3_X1 u0_u9_u7_U96 (.A3( u0_u9_u7_n131 ) , .A2( u0_u9_u7_n132 ) , .A1( u0_u9_u7_n133 ) , .ZN( u0_u9_u7_n135 ) );
  OAI22_X1 u0_uk_U117 (.ZN( u0_K10_47 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n249 ) , .A2( u0_uk_n264 ) );
  INV_X1 u0_uk_U149 (.ZN( u0_K14_19 ) , .A( u0_uk_n938 ) );
  AOI22_X1 u0_uk_U150 (.B2( u0_uk_K_r12_25 ) , .A2( u0_uk_K_r12_33 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n207 ) , .ZN( u0_uk_n938 ) );
  OAI22_X1 u0_uk_U166 (.ZN( u0_K14_30 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n250 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n77 ) );
  OAI22_X1 u0_uk_U169 (.ZN( u0_K10_30 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n232 ) , .B2( u0_uk_n260 ) );
  OAI21_X1 u0_uk_U226 (.ZN( u0_K10_31 ) , .A( u0_uk_n1014 ) , .B2( u0_uk_n243 ) , .B1( u0_uk_n250 ) );
  NAND2_X1 u0_uk_U227 (.A1( u0_uk_K_r8_16 ) , .ZN( u0_uk_n1014 ) , .A2( u0_uk_n207 ) );
  OAI22_X1 u0_uk_U262 (.ZN( u0_K10_44 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n241 ) , .B2( u0_uk_n261 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U263 (.ZN( u0_K10_48 ) , .A2( u0_uk_n232 ) , .A1( u0_uk_n240 ) , .B2( u0_uk_n248 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U315 (.ZN( u0_K14_26 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n49 ) , .B2( u0_uk_n66 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U317 (.ZN( u0_K10_26 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n233 ) , .B2( u0_uk_n249 ) );
  OAI22_X1 u0_uk_U373 (.ZN( u0_K14_28 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n61 ) , .B2( u0_uk_n67 ) );
  OAI22_X1 u0_uk_U383 (.ZN( u0_K10_28 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n241 ) , .B2( u0_uk_n248 ) );
  INV_X1 u0_uk_U439 (.ZN( u0_K10_33 ) , .A( u0_uk_n1012 ) );
  OAI21_X1 u0_uk_U472 (.ZN( u0_K14_29 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n51 ) , .A( u0_uk_n935 ) );
  NAND2_X1 u0_uk_U473 (.A1( u0_uk_K_r12_44 ) , .A2( u0_uk_n145 ) , .ZN( u0_uk_n935 ) );
  OAI22_X1 u0_uk_U483 (.ZN( u0_K10_29 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n233 ) , .B2( u0_uk_n261 ) );
  OAI22_X1 u0_uk_U538 (.ZN( u0_K14_17 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n54 ) , .B2( u0_uk_n78 ) );
  INV_X1 u0_uk_U614 (.ZN( u0_K10_35 ) , .A( u0_uk_n1011 ) );
  AOI22_X1 u0_uk_U615 (.B2( u0_uk_K_r8_2 ) , .A2( u0_uk_K_r8_37 ) , .ZN( u0_uk_n1011 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U626 (.ZN( u0_K14_11 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n80 ) , .B1( u0_uk_n83 ) , .A2( u0_uk_n87 ) );
  OAI22_X1 u0_uk_U669 (.ZN( u0_K10_43 ) , .A1( u0_uk_n214 ) , .B2( u0_uk_n237 ) , .A2( u0_uk_n265 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U670 (.ZN( u0_K10_45 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n244 ) , .B2( u0_uk_n260 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U868 (.ZN( u0_K14_22 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n48 ) , .B2( u0_uk_n86 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U874 (.ZN( u0_K14_23 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n79 ) , .A2( u0_uk_n86 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U899 (.ZN( u0_K14_7 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n53 ) , .B2( u0_uk_n72 ) );
  OAI22_X1 u0_uk_U938 (.ZN( u0_K14_8 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n69 ) , .A2( u0_uk_n87 ) );
  OAI22_X1 u0_uk_U940 (.ZN( u0_K14_20 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n69 ) , .B2( u0_uk_n75 ) , .A1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U948 (.ZN( u0_K10_46 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n247 ) , .B2( u0_uk_n256 ) );
  OAI22_X1 u0_uk_U964 (.ZN( u0_K14_16 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n46 ) , .A2( u0_uk_n84 ) );
  OAI22_X1 u0_uk_U989 (.ZN( u0_K14_25 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n82 ) , .B2( u0_uk_n88 ) );
  XOR2_X1 u1_U148 (.Z( u1_N4 ) , .B( u1_desIn_r_38 ) , .A( u1_out0_5 ) );
  XOR2_X1 u1_U242 (.B( u1_L8_27 ) , .Z( u1_N314 ) , .A( u1_out9_27 ) );
  XOR2_X1 u1_U247 (.Z( u1_N31 ) , .B( u1_desIn_r_56 ) , .A( u1_out0_32 ) );
  XOR2_X1 u1_U249 (.B( u1_L8_21 ) , .Z( u1_N308 ) , .A( u1_out9_21 ) );
  XOR2_X1 u1_U255 (.B( u1_L8_15 ) , .Z( u1_N302 ) , .A( u1_out9_15 ) );
  XOR2_X1 u1_U259 (.Z( u1_N3 ) , .B( u1_desIn_r_30 ) , .A( u1_out0_4 ) );
  XOR2_X1 u1_U267 (.B( u1_L8_5 ) , .Z( u1_N292 ) , .A( u1_out9_5 ) );
  XOR2_X1 u1_U274 (.B( u1_L7_31 ) , .Z( u1_N286 ) , .A( u1_out8_31 ) );
  XOR2_X1 u1_U275 (.B( u1_L7_30 ) , .Z( u1_N285 ) , .A( u1_out8_30 ) );
  XOR2_X1 u1_U277 (.B( u1_L7_28 ) , .Z( u1_N283 ) , .A( u1_out8_28 ) );
  XOR2_X1 u1_U279 (.B( u1_L7_26 ) , .Z( u1_N281 ) , .A( u1_out8_26 ) );
  XOR2_X1 u1_U281 (.Z( u1_N28 ) , .B( u1_desIn_r_32 ) , .A( u1_out0_29 ) );
  XOR2_X1 u1_U282 (.B( u1_L7_24 ) , .Z( u1_N279 ) , .A( u1_out8_24 ) );
  XOR2_X1 u1_U283 (.B( u1_L7_23 ) , .Z( u1_N278 ) , .A( u1_out8_23 ) );
  XOR2_X1 u1_U286 (.B( u1_L7_20 ) , .Z( u1_N275 ) , .A( u1_out8_20 ) );
  XOR2_X1 u1_U288 (.B( u1_L7_18 ) , .Z( u1_N273 ) , .A( u1_out8_18 ) );
  XOR2_X1 u1_U289 (.B( u1_L7_17 ) , .Z( u1_N272 ) , .A( u1_out8_17 ) );
  XOR2_X1 u1_U290 (.B( u1_L7_16 ) , .Z( u1_N271 ) , .A( u1_out8_16 ) );
  XOR2_X1 u1_U294 (.B( u1_L7_13 ) , .Z( u1_N268 ) , .A( u1_out8_13 ) );
  XOR2_X1 u1_U297 (.B( u1_L7_10 ) , .Z( u1_N265 ) , .A( u1_out8_10 ) );
  XOR2_X1 u1_U298 (.B( u1_L7_9 ) , .Z( u1_N264 ) , .A( u1_out8_9 ) );
  XOR2_X1 u1_U301 (.B( u1_L7_6 ) , .Z( u1_N261 ) , .A( u1_out8_6 ) );
  XOR2_X1 u1_U303 (.Z( u1_N26 ) , .B( u1_desIn_r_16 ) , .A( u1_out0_27 ) );
  XOR2_X1 u1_U306 (.B( u1_L7_2 ) , .Z( u1_N257 ) , .A( u1_out8_2 ) );
  XOR2_X1 u1_U307 (.B( u1_L7_1 ) , .Z( u1_N256 ) , .A( u1_out8_1 ) );
  XOR2_X1 u1_U325 (.Z( u1_N24 ) , .B( u1_desIn_r_0 ) , .A( u1_out0_25 ) );
  XOR2_X1 u1_U35 (.Z( u1_N7 ) , .B( u1_desIn_r_62 ) , .A( u1_out0_8 ) );
  XOR2_X1 u1_U358 (.Z( u1_N21 ) , .B( u1_desIn_r_42 ) , .A( u1_out0_22 ) );
  XOR2_X1 u1_U369 (.Z( u1_N20 ) , .B( u1_desIn_r_34 ) , .A( u1_out0_21 ) );
  XOR2_X1 u1_U370 (.Z( u1_N2 ) , .B( u1_desIn_r_22 ) , .A( u1_out0_3 ) );
  XOR2_X1 u1_U379 (.B( u1_L4_32 ) , .Z( u1_N191 ) , .A( u1_out5_32 ) );
  XOR2_X1 u1_U380 (.B( u1_L4_31 ) , .Z( u1_N190 ) , .A( u1_out5_31 ) );
  XOR2_X1 u1_U382 (.B( u1_L4_30 ) , .Z( u1_N189 ) , .A( u1_out5_30 ) );
  XOR2_X1 u1_U383 (.B( u1_L4_29 ) , .Z( u1_N188 ) , .A( u1_out5_29 ) );
  XOR2_X1 u1_U386 (.B( u1_L4_26 ) , .Z( u1_N185 ) , .A( u1_out5_26 ) );
  XOR2_X1 u1_U387 (.B( u1_L4_25 ) , .Z( u1_N184 ) , .A( u1_out5_25 ) );
  XOR2_X1 u1_U388 (.B( u1_L4_24 ) , .Z( u1_N183 ) , .A( u1_out5_24 ) );
  XOR2_X1 u1_U389 (.B( u1_L4_23 ) , .Z( u1_N182 ) , .A( u1_out5_23 ) );
  XOR2_X1 u1_U390 (.B( u1_L4_22 ) , .Z( u1_N181 ) , .A( u1_out5_22 ) );
  XOR2_X1 u1_U392 (.Z( u1_N18 ) , .B( u1_desIn_r_18 ) , .A( u1_out0_19 ) );
  XOR2_X1 u1_U393 (.B( u1_L4_20 ) , .Z( u1_N179 ) , .A( u1_out5_20 ) );
  XOR2_X1 u1_U394 (.B( u1_L4_19 ) , .Z( u1_N178 ) , .A( u1_out5_19 ) );
  XOR2_X1 u1_U396 (.B( u1_L4_17 ) , .Z( u1_N176 ) , .A( u1_out5_17 ) );
  XOR2_X1 u1_U397 (.B( u1_L4_16 ) , .Z( u1_N175 ) , .A( u1_out5_16 ) );
  XOR2_X1 u1_U399 (.B( u1_L4_14 ) , .Z( u1_N173 ) , .A( u1_out5_14 ) );
  XOR2_X1 u1_U401 (.B( u1_L4_12 ) , .Z( u1_N171 ) , .A( u1_out5_12 ) );
  XOR2_X1 u1_U402 (.B( u1_L4_11 ) , .Z( u1_N170 ) , .A( u1_out5_11 ) );
  XOR2_X1 u1_U404 (.B( u1_L4_10 ) , .Z( u1_N169 ) , .A( u1_out5_10 ) );
  XOR2_X1 u1_U405 (.B( u1_L4_9 ) , .Z( u1_N168 ) , .A( u1_out5_9 ) );
  XOR2_X1 u1_U406 (.B( u1_L4_8 ) , .Z( u1_N167 ) , .A( u1_out5_8 ) );
  XOR2_X1 u1_U407 (.B( u1_L4_7 ) , .Z( u1_N166 ) , .A( u1_out5_7 ) );
  XOR2_X1 u1_U408 (.B( u1_L4_6 ) , .Z( u1_N165 ) , .A( u1_out5_6 ) );
  XOR2_X1 u1_U410 (.B( u1_L4_4 ) , .Z( u1_N163 ) , .A( u1_out5_4 ) );
  XOR2_X1 u1_U411 (.B( u1_L4_3 ) , .Z( u1_N162 ) , .A( u1_out5_3 ) );
  XOR2_X1 u1_U413 (.B( u1_L4_1 ) , .Z( u1_N160 ) , .A( u1_out5_1 ) );
  XOR2_X1 u1_U418 (.B( u1_L3_29 ) , .Z( u1_N156 ) , .A( u1_out4_29 ) );
  XOR2_X1 u1_U429 (.B( u1_L3_19 ) , .Z( u1_N146 ) , .A( u1_out4_19 ) );
  XOR2_X1 u1_U436 (.Z( u1_N14 ) , .B( u1_desIn_r_52 ) , .A( u1_out0_15 ) );
  XOR2_X1 u1_U438 (.B( u1_L3_11 ) , .Z( u1_N138 ) , .A( u1_out4_11 ) );
  XOR2_X1 u1_U445 (.B( u1_L3_4 ) , .Z( u1_N131 ) , .A( u1_out4_4 ) );
  XOR2_X1 u1_U447 (.Z( u1_N13 ) , .B( u1_desIn_r_44 ) , .A( u1_out0_14 ) );
  XOR2_X1 u1_U454 (.B( u1_L2_28 ) , .Z( u1_N123 ) , .A( u1_out3_28 ) );
  XOR2_X1 u1_U46 (.Z( u1_N6 ) , .B( u1_desIn_r_54 ) , .A( u1_out0_7 ) );
  XOR2_X1 u1_U465 (.B( u1_L2_18 ) , .Z( u1_N113 ) , .A( u1_out3_18 ) );
  XOR2_X1 u1_U469 (.Z( u1_N11 ) , .B( u1_desIn_r_28 ) , .A( u1_out0_12 ) );
  XOR2_X1 u1_U471 (.B( u1_L2_13 ) , .Z( u1_N108 ) , .A( u1_out3_13 ) );
  XOR2_X1 u1_U480 (.Z( u1_N10 ) , .B( u1_desIn_r_20 ) , .A( u1_out0_11 ) );
  XOR2_X1 u1_U5 (.B( u1_L2_2 ) , .Z( u1_N97 ) , .A( u1_out3_2 ) );
  XOR2_X1 u1_U60 (.B( u1_L13_32 ) , .Z( u1_N479 ) , .A( u1_out14_32 ) );
  XOR2_X1 u1_U63 (.B( u1_L13_29 ) , .Z( u1_N476 ) , .A( u1_out14_29 ) );
  XOR2_X1 u1_U65 (.B( u1_L13_27 ) , .Z( u1_N474 ) , .A( u1_out14_27 ) );
  XOR2_X1 u1_U71 (.B( u1_L13_22 ) , .Z( u1_N469 ) , .A( u1_out14_22 ) );
  XOR2_X1 u1_U72 (.B( u1_L13_21 ) , .Z( u1_N468 ) , .A( u1_out14_21 ) );
  XOR2_X1 u1_U74 (.B( u1_L13_19 ) , .Z( u1_N466 ) , .A( u1_out14_19 ) );
  XOR2_X1 u1_U78 (.B( u1_L13_15 ) , .Z( u1_N462 ) , .A( u1_out14_15 ) );
  XOR2_X1 u1_U82 (.B( u1_L13_12 ) , .Z( u1_N459 ) , .A( u1_out14_12 ) );
  XOR2_X1 u1_U83 (.B( u1_L13_11 ) , .Z( u1_N458 ) , .A( u1_out14_11 ) );
  XOR2_X1 u1_U87 (.B( u1_L13_7 ) , .Z( u1_N454 ) , .A( u1_out14_7 ) );
  XOR2_X1 u1_U89 (.B( u1_L13_5 ) , .Z( u1_N452 ) , .A( u1_out14_5 ) );
  XOR2_X1 u1_U90 (.B( u1_L13_4 ) , .Z( u1_N451 ) , .A( u1_out14_4 ) );
  XOR2_X1 u1_u0_U10 (.B( u1_K1_45 ) , .A( u1_desIn_r_41 ) , .Z( u1_u0_X_45 ) );
  XOR2_X1 u1_u0_U11 (.B( u1_K1_44 ) , .A( u1_desIn_r_33 ) , .Z( u1_u0_X_44 ) );
  XOR2_X1 u1_u0_U12 (.B( u1_K1_43 ) , .A( u1_desIn_r_25 ) , .Z( u1_u0_X_43 ) );
  XOR2_X1 u1_u0_U13 (.B( u1_K1_42 ) , .A( u1_desIn_r_33 ) , .Z( u1_u0_X_42 ) );
  XOR2_X1 u1_u0_U14 (.B( u1_K1_41 ) , .A( u1_desIn_r_25 ) , .Z( u1_u0_X_41 ) );
  XOR2_X1 u1_u0_U15 (.B( u1_K1_40 ) , .A( u1_desIn_r_17 ) , .Z( u1_u0_X_40 ) );
  XOR2_X1 u1_u0_U17 (.B( u1_K1_39 ) , .A( u1_desIn_r_9 ) , .Z( u1_u0_X_39 ) );
  XOR2_X1 u1_u0_U18 (.B( u1_K1_38 ) , .A( u1_desIn_r_1 ) , .Z( u1_u0_X_38 ) );
  XOR2_X1 u1_u0_U19 (.B( u1_K1_37 ) , .A( u1_desIn_r_59 ) , .Z( u1_u0_X_37 ) );
  XOR2_X1 u1_u0_U20 (.B( u1_K1_36 ) , .A( u1_desIn_r_1 ) , .Z( u1_u0_X_36 ) );
  XOR2_X1 u1_u0_U21 (.B( u1_K1_35 ) , .A( u1_desIn_r_59 ) , .Z( u1_u0_X_35 ) );
  XOR2_X1 u1_u0_U22 (.B( u1_K1_34 ) , .A( u1_desIn_r_51 ) , .Z( u1_u0_X_34 ) );
  XOR2_X1 u1_u0_U23 (.B( u1_K1_33 ) , .A( u1_desIn_r_43 ) , .Z( u1_u0_X_33 ) );
  XOR2_X1 u1_u0_U24 (.B( u1_K1_32 ) , .A( u1_desIn_r_35 ) , .Z( u1_u0_X_32 ) );
  XOR2_X1 u1_u0_U25 (.B( u1_K1_31 ) , .A( u1_desIn_r_27 ) , .Z( u1_u0_X_31 ) );
  XOR2_X1 u1_u0_U26 (.B( u1_K1_30 ) , .A( u1_desIn_r_35 ) , .Z( u1_u0_X_30 ) );
  XOR2_X1 u1_u0_U28 (.B( u1_K1_29 ) , .A( u1_desIn_r_27 ) , .Z( u1_u0_X_29 ) );
  XOR2_X1 u1_u0_U29 (.B( u1_K1_28 ) , .A( u1_desIn_r_19 ) , .Z( u1_u0_X_28 ) );
  XOR2_X1 u1_u0_U30 (.B( u1_K1_27 ) , .A( u1_desIn_r_11 ) , .Z( u1_u0_X_27 ) );
  XOR2_X1 u1_u0_U31 (.B( u1_K1_26 ) , .A( u1_desIn_r_3 ) , .Z( u1_u0_X_26 ) );
  XOR2_X1 u1_u0_U32 (.B( u1_K1_25 ) , .A( u1_desIn_r_61 ) , .Z( u1_u0_X_25 ) );
  XOR2_X1 u1_u0_U7 (.B( u1_K1_48 ) , .A( u1_desIn_r_7 ) , .Z( u1_u0_X_48 ) );
  XOR2_X1 u1_u0_U8 (.B( u1_K1_47 ) , .A( u1_desIn_r_57 ) , .Z( u1_u0_X_47 ) );
  XOR2_X1 u1_u0_U9 (.B( u1_K1_46 ) , .A( u1_desIn_r_49 ) , .Z( u1_u0_X_46 ) );
  OAI22_X1 u1_u0_u4_U10 (.B2( u1_u0_u4_n135 ) , .ZN( u1_u0_u4_n137 ) , .B1( u1_u0_u4_n153 ) , .A1( u1_u0_u4_n155 ) , .A2( u1_u0_u4_n171 ) );
  AND3_X1 u1_u0_u4_U11 (.A2( u1_u0_u4_n134 ) , .ZN( u1_u0_u4_n135 ) , .A3( u1_u0_u4_n145 ) , .A1( u1_u0_u4_n157 ) );
  NAND2_X1 u1_u0_u4_U12 (.ZN( u1_u0_u4_n132 ) , .A2( u1_u0_u4_n170 ) , .A1( u1_u0_u4_n173 ) );
  AOI21_X1 u1_u0_u4_U13 (.B2( u1_u0_u4_n160 ) , .B1( u1_u0_u4_n161 ) , .ZN( u1_u0_u4_n162 ) , .A( u1_u0_u4_n170 ) );
  AOI21_X1 u1_u0_u4_U14 (.ZN( u1_u0_u4_n107 ) , .B2( u1_u0_u4_n143 ) , .A( u1_u0_u4_n174 ) , .B1( u1_u0_u4_n184 ) );
  AOI21_X1 u1_u0_u4_U15 (.B2( u1_u0_u4_n158 ) , .B1( u1_u0_u4_n159 ) , .ZN( u1_u0_u4_n163 ) , .A( u1_u0_u4_n174 ) );
  AOI21_X1 u1_u0_u4_U16 (.A( u1_u0_u4_n153 ) , .B2( u1_u0_u4_n154 ) , .B1( u1_u0_u4_n155 ) , .ZN( u1_u0_u4_n165 ) );
  AOI21_X1 u1_u0_u4_U17 (.A( u1_u0_u4_n156 ) , .B2( u1_u0_u4_n157 ) , .ZN( u1_u0_u4_n164 ) , .B1( u1_u0_u4_n184 ) );
  INV_X1 u1_u0_u4_U18 (.A( u1_u0_u4_n138 ) , .ZN( u1_u0_u4_n170 ) );
  AND2_X1 u1_u0_u4_U19 (.A2( u1_u0_u4_n120 ) , .ZN( u1_u0_u4_n155 ) , .A1( u1_u0_u4_n160 ) );
  INV_X1 u1_u0_u4_U20 (.A( u1_u0_u4_n156 ) , .ZN( u1_u0_u4_n175 ) );
  NAND2_X1 u1_u0_u4_U21 (.A2( u1_u0_u4_n118 ) , .ZN( u1_u0_u4_n131 ) , .A1( u1_u0_u4_n147 ) );
  NAND2_X1 u1_u0_u4_U22 (.A1( u1_u0_u4_n119 ) , .A2( u1_u0_u4_n120 ) , .ZN( u1_u0_u4_n130 ) );
  NAND2_X1 u1_u0_u4_U23 (.ZN( u1_u0_u4_n117 ) , .A2( u1_u0_u4_n118 ) , .A1( u1_u0_u4_n148 ) );
  NAND2_X1 u1_u0_u4_U24 (.ZN( u1_u0_u4_n129 ) , .A1( u1_u0_u4_n134 ) , .A2( u1_u0_u4_n148 ) );
  AND3_X1 u1_u0_u4_U25 (.A1( u1_u0_u4_n119 ) , .A2( u1_u0_u4_n143 ) , .A3( u1_u0_u4_n154 ) , .ZN( u1_u0_u4_n161 ) );
  AND2_X1 u1_u0_u4_U26 (.A1( u1_u0_u4_n145 ) , .A2( u1_u0_u4_n147 ) , .ZN( u1_u0_u4_n159 ) );
  OR3_X1 u1_u0_u4_U27 (.A3( u1_u0_u4_n114 ) , .A2( u1_u0_u4_n115 ) , .A1( u1_u0_u4_n116 ) , .ZN( u1_u0_u4_n136 ) );
  AOI21_X1 u1_u0_u4_U28 (.A( u1_u0_u4_n113 ) , .ZN( u1_u0_u4_n116 ) , .B2( u1_u0_u4_n173 ) , .B1( u1_u0_u4_n174 ) );
  AOI21_X1 u1_u0_u4_U29 (.ZN( u1_u0_u4_n115 ) , .B2( u1_u0_u4_n145 ) , .B1( u1_u0_u4_n146 ) , .A( u1_u0_u4_n156 ) );
  NOR2_X1 u1_u0_u4_U3 (.ZN( u1_u0_u4_n121 ) , .A1( u1_u0_u4_n181 ) , .A2( u1_u0_u4_n182 ) );
  OAI22_X1 u1_u0_u4_U30 (.ZN( u1_u0_u4_n114 ) , .A2( u1_u0_u4_n121 ) , .B1( u1_u0_u4_n160 ) , .B2( u1_u0_u4_n170 ) , .A1( u1_u0_u4_n171 ) );
  INV_X1 u1_u0_u4_U31 (.A( u1_u0_u4_n158 ) , .ZN( u1_u0_u4_n182 ) );
  INV_X1 u1_u0_u4_U32 (.ZN( u1_u0_u4_n181 ) , .A( u1_u0_u4_n96 ) );
  INV_X1 u1_u0_u4_U33 (.A( u1_u0_u4_n144 ) , .ZN( u1_u0_u4_n179 ) );
  INV_X1 u1_u0_u4_U34 (.A( u1_u0_u4_n157 ) , .ZN( u1_u0_u4_n178 ) );
  NAND2_X1 u1_u0_u4_U35 (.A2( u1_u0_u4_n154 ) , .A1( u1_u0_u4_n96 ) , .ZN( u1_u0_u4_n97 ) );
  INV_X1 u1_u0_u4_U36 (.ZN( u1_u0_u4_n186 ) , .A( u1_u0_u4_n95 ) );
  OAI221_X1 u1_u0_u4_U37 (.C1( u1_u0_u4_n134 ) , .B1( u1_u0_u4_n158 ) , .B2( u1_u0_u4_n171 ) , .C2( u1_u0_u4_n173 ) , .A( u1_u0_u4_n94 ) , .ZN( u1_u0_u4_n95 ) );
  AOI222_X1 u1_u0_u4_U38 (.B2( u1_u0_u4_n132 ) , .A1( u1_u0_u4_n138 ) , .C2( u1_u0_u4_n175 ) , .A2( u1_u0_u4_n179 ) , .C1( u1_u0_u4_n181 ) , .B1( u1_u0_u4_n185 ) , .ZN( u1_u0_u4_n94 ) );
  INV_X1 u1_u0_u4_U39 (.A( u1_u0_u4_n113 ) , .ZN( u1_u0_u4_n185 ) );
  INV_X1 u1_u0_u4_U4 (.A( u1_u0_u4_n117 ) , .ZN( u1_u0_u4_n184 ) );
  INV_X1 u1_u0_u4_U40 (.A( u1_u0_u4_n143 ) , .ZN( u1_u0_u4_n183 ) );
  NOR2_X1 u1_u0_u4_U41 (.ZN( u1_u0_u4_n138 ) , .A1( u1_u0_u4_n168 ) , .A2( u1_u0_u4_n169 ) );
  NOR2_X1 u1_u0_u4_U42 (.A1( u1_u0_u4_n150 ) , .A2( u1_u0_u4_n152 ) , .ZN( u1_u0_u4_n153 ) );
  NOR2_X1 u1_u0_u4_U43 (.A2( u1_u0_u4_n128 ) , .A1( u1_u0_u4_n138 ) , .ZN( u1_u0_u4_n156 ) );
  AOI22_X1 u1_u0_u4_U44 (.B2( u1_u0_u4_n122 ) , .A1( u1_u0_u4_n123 ) , .ZN( u1_u0_u4_n124 ) , .B1( u1_u0_u4_n128 ) , .A2( u1_u0_u4_n172 ) );
  INV_X1 u1_u0_u4_U45 (.A( u1_u0_u4_n153 ) , .ZN( u1_u0_u4_n172 ) );
  NAND2_X1 u1_u0_u4_U46 (.A2( u1_u0_u4_n120 ) , .ZN( u1_u0_u4_n123 ) , .A1( u1_u0_u4_n161 ) );
  AOI22_X1 u1_u0_u4_U47 (.B2( u1_u0_u4_n132 ) , .A2( u1_u0_u4_n133 ) , .ZN( u1_u0_u4_n140 ) , .A1( u1_u0_u4_n150 ) , .B1( u1_u0_u4_n179 ) );
  NAND2_X1 u1_u0_u4_U48 (.ZN( u1_u0_u4_n133 ) , .A2( u1_u0_u4_n146 ) , .A1( u1_u0_u4_n154 ) );
  NAND2_X1 u1_u0_u4_U49 (.A1( u1_u0_u4_n103 ) , .ZN( u1_u0_u4_n154 ) , .A2( u1_u0_u4_n98 ) );
  NOR4_X1 u1_u0_u4_U5 (.A4( u1_u0_u4_n106 ) , .A3( u1_u0_u4_n107 ) , .A2( u1_u0_u4_n108 ) , .A1( u1_u0_u4_n109 ) , .ZN( u1_u0_u4_n110 ) );
  NAND2_X1 u1_u0_u4_U50 (.A1( u1_u0_u4_n101 ) , .ZN( u1_u0_u4_n158 ) , .A2( u1_u0_u4_n99 ) );
  AOI21_X1 u1_u0_u4_U51 (.ZN( u1_u0_u4_n127 ) , .A( u1_u0_u4_n136 ) , .B2( u1_u0_u4_n150 ) , .B1( u1_u0_u4_n180 ) );
  INV_X1 u1_u0_u4_U52 (.A( u1_u0_u4_n160 ) , .ZN( u1_u0_u4_n180 ) );
  NAND2_X1 u1_u0_u4_U53 (.A2( u1_u0_u4_n104 ) , .A1( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n146 ) );
  NAND2_X1 u1_u0_u4_U54 (.A2( u1_u0_u4_n101 ) , .A1( u1_u0_u4_n102 ) , .ZN( u1_u0_u4_n160 ) );
  NAND2_X1 u1_u0_u4_U55 (.ZN( u1_u0_u4_n134 ) , .A1( u1_u0_u4_n98 ) , .A2( u1_u0_u4_n99 ) );
  NAND2_X1 u1_u0_u4_U56 (.A1( u1_u0_u4_n103 ) , .A2( u1_u0_u4_n104 ) , .ZN( u1_u0_u4_n143 ) );
  NAND2_X1 u1_u0_u4_U57 (.A2( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n145 ) , .A1( u1_u0_u4_n98 ) );
  NAND2_X1 u1_u0_u4_U58 (.A1( u1_u0_u4_n100 ) , .A2( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n120 ) );
  NAND2_X1 u1_u0_u4_U59 (.A1( u1_u0_u4_n102 ) , .A2( u1_u0_u4_n104 ) , .ZN( u1_u0_u4_n148 ) );
  AOI21_X1 u1_u0_u4_U6 (.ZN( u1_u0_u4_n106 ) , .B2( u1_u0_u4_n146 ) , .B1( u1_u0_u4_n158 ) , .A( u1_u0_u4_n170 ) );
  NAND2_X1 u1_u0_u4_U60 (.A2( u1_u0_u4_n100 ) , .A1( u1_u0_u4_n103 ) , .ZN( u1_u0_u4_n157 ) );
  INV_X1 u1_u0_u4_U61 (.A( u1_u0_u4_n150 ) , .ZN( u1_u0_u4_n173 ) );
  INV_X1 u1_u0_u4_U62 (.A( u1_u0_u4_n152 ) , .ZN( u1_u0_u4_n171 ) );
  NAND2_X1 u1_u0_u4_U63 (.A1( u1_u0_u4_n100 ) , .ZN( u1_u0_u4_n118 ) , .A2( u1_u0_u4_n99 ) );
  NAND2_X1 u1_u0_u4_U64 (.A2( u1_u0_u4_n100 ) , .A1( u1_u0_u4_n102 ) , .ZN( u1_u0_u4_n144 ) );
  NAND2_X1 u1_u0_u4_U65 (.A2( u1_u0_u4_n101 ) , .A1( u1_u0_u4_n105 ) , .ZN( u1_u0_u4_n96 ) );
  INV_X1 u1_u0_u4_U66 (.A( u1_u0_u4_n128 ) , .ZN( u1_u0_u4_n174 ) );
  NAND2_X1 u1_u0_u4_U67 (.A2( u1_u0_u4_n102 ) , .ZN( u1_u0_u4_n119 ) , .A1( u1_u0_u4_n98 ) );
  NAND2_X1 u1_u0_u4_U68 (.A2( u1_u0_u4_n101 ) , .A1( u1_u0_u4_n103 ) , .ZN( u1_u0_u4_n147 ) );
  NAND2_X1 u1_u0_u4_U69 (.A2( u1_u0_u4_n104 ) , .ZN( u1_u0_u4_n113 ) , .A1( u1_u0_u4_n99 ) );
  AOI21_X1 u1_u0_u4_U7 (.ZN( u1_u0_u4_n108 ) , .B2( u1_u0_u4_n134 ) , .B1( u1_u0_u4_n155 ) , .A( u1_u0_u4_n156 ) );
  NOR2_X1 u1_u0_u4_U70 (.A2( u1_u0_X_28 ) , .ZN( u1_u0_u4_n150 ) , .A1( u1_u0_u4_n168 ) );
  NOR2_X1 u1_u0_u4_U71 (.A2( u1_u0_X_29 ) , .ZN( u1_u0_u4_n152 ) , .A1( u1_u0_u4_n169 ) );
  NOR2_X1 u1_u0_u4_U72 (.A2( u1_u0_X_30 ) , .ZN( u1_u0_u4_n105 ) , .A1( u1_u0_u4_n176 ) );
  NOR2_X1 u1_u0_u4_U73 (.A2( u1_u0_X_26 ) , .ZN( u1_u0_u4_n100 ) , .A1( u1_u0_u4_n177 ) );
  NOR2_X1 u1_u0_u4_U74 (.A2( u1_u0_X_28 ) , .A1( u1_u0_X_29 ) , .ZN( u1_u0_u4_n128 ) );
  NOR2_X1 u1_u0_u4_U75 (.A2( u1_u0_X_27 ) , .A1( u1_u0_X_30 ) , .ZN( u1_u0_u4_n102 ) );
  NOR2_X1 u1_u0_u4_U76 (.A2( u1_u0_X_25 ) , .A1( u1_u0_X_26 ) , .ZN( u1_u0_u4_n98 ) );
  AND2_X1 u1_u0_u4_U77 (.A2( u1_u0_X_25 ) , .A1( u1_u0_X_26 ) , .ZN( u1_u0_u4_n104 ) );
  AND2_X1 u1_u0_u4_U78 (.A1( u1_u0_X_30 ) , .A2( u1_u0_u4_n176 ) , .ZN( u1_u0_u4_n99 ) );
  AND2_X1 u1_u0_u4_U79 (.A1( u1_u0_X_26 ) , .ZN( u1_u0_u4_n101 ) , .A2( u1_u0_u4_n177 ) );
  AOI21_X1 u1_u0_u4_U8 (.ZN( u1_u0_u4_n109 ) , .A( u1_u0_u4_n153 ) , .B1( u1_u0_u4_n159 ) , .B2( u1_u0_u4_n184 ) );
  AND2_X1 u1_u0_u4_U80 (.A1( u1_u0_X_27 ) , .A2( u1_u0_X_30 ) , .ZN( u1_u0_u4_n103 ) );
  INV_X1 u1_u0_u4_U81 (.A( u1_u0_X_28 ) , .ZN( u1_u0_u4_n169 ) );
  INV_X1 u1_u0_u4_U82 (.A( u1_u0_X_29 ) , .ZN( u1_u0_u4_n168 ) );
  INV_X1 u1_u0_u4_U83 (.A( u1_u0_X_25 ) , .ZN( u1_u0_u4_n177 ) );
  INV_X1 u1_u0_u4_U84 (.A( u1_u0_X_27 ) , .ZN( u1_u0_u4_n176 ) );
  NAND4_X1 u1_u0_u4_U85 (.ZN( u1_out0_25 ) , .A4( u1_u0_u4_n139 ) , .A3( u1_u0_u4_n140 ) , .A2( u1_u0_u4_n141 ) , .A1( u1_u0_u4_n142 ) );
  OAI21_X1 u1_u0_u4_U86 (.A( u1_u0_u4_n128 ) , .B2( u1_u0_u4_n129 ) , .B1( u1_u0_u4_n130 ) , .ZN( u1_u0_u4_n142 ) );
  OAI21_X1 u1_u0_u4_U87 (.B2( u1_u0_u4_n131 ) , .ZN( u1_u0_u4_n141 ) , .A( u1_u0_u4_n175 ) , .B1( u1_u0_u4_n183 ) );
  NAND4_X1 u1_u0_u4_U88 (.ZN( u1_out0_14 ) , .A4( u1_u0_u4_n124 ) , .A3( u1_u0_u4_n125 ) , .A2( u1_u0_u4_n126 ) , .A1( u1_u0_u4_n127 ) );
  AOI22_X1 u1_u0_u4_U89 (.B2( u1_u0_u4_n117 ) , .ZN( u1_u0_u4_n126 ) , .A1( u1_u0_u4_n129 ) , .B1( u1_u0_u4_n152 ) , .A2( u1_u0_u4_n175 ) );
  AOI211_X1 u1_u0_u4_U9 (.B( u1_u0_u4_n136 ) , .A( u1_u0_u4_n137 ) , .C2( u1_u0_u4_n138 ) , .ZN( u1_u0_u4_n139 ) , .C1( u1_u0_u4_n182 ) );
  AOI22_X1 u1_u0_u4_U90 (.ZN( u1_u0_u4_n125 ) , .B2( u1_u0_u4_n131 ) , .A2( u1_u0_u4_n132 ) , .B1( u1_u0_u4_n138 ) , .A1( u1_u0_u4_n178 ) );
  NAND4_X1 u1_u0_u4_U91 (.ZN( u1_out0_8 ) , .A4( u1_u0_u4_n110 ) , .A3( u1_u0_u4_n111 ) , .A2( u1_u0_u4_n112 ) , .A1( u1_u0_u4_n186 ) );
  NAND2_X1 u1_u0_u4_U92 (.ZN( u1_u0_u4_n112 ) , .A2( u1_u0_u4_n130 ) , .A1( u1_u0_u4_n150 ) );
  AOI22_X1 u1_u0_u4_U93 (.ZN( u1_u0_u4_n111 ) , .B2( u1_u0_u4_n132 ) , .A1( u1_u0_u4_n152 ) , .B1( u1_u0_u4_n178 ) , .A2( u1_u0_u4_n97 ) );
  AOI22_X1 u1_u0_u4_U94 (.B2( u1_u0_u4_n149 ) , .B1( u1_u0_u4_n150 ) , .A2( u1_u0_u4_n151 ) , .A1( u1_u0_u4_n152 ) , .ZN( u1_u0_u4_n167 ) );
  NOR4_X1 u1_u0_u4_U95 (.A4( u1_u0_u4_n162 ) , .A3( u1_u0_u4_n163 ) , .A2( u1_u0_u4_n164 ) , .A1( u1_u0_u4_n165 ) , .ZN( u1_u0_u4_n166 ) );
  NAND3_X1 u1_u0_u4_U96 (.ZN( u1_out0_3 ) , .A3( u1_u0_u4_n166 ) , .A1( u1_u0_u4_n167 ) , .A2( u1_u0_u4_n186 ) );
  NAND3_X1 u1_u0_u4_U97 (.A3( u1_u0_u4_n146 ) , .A2( u1_u0_u4_n147 ) , .A1( u1_u0_u4_n148 ) , .ZN( u1_u0_u4_n149 ) );
  NAND3_X1 u1_u0_u4_U98 (.A3( u1_u0_u4_n143 ) , .A2( u1_u0_u4_n144 ) , .A1( u1_u0_u4_n145 ) , .ZN( u1_u0_u4_n151 ) );
  NAND3_X1 u1_u0_u4_U99 (.A3( u1_u0_u4_n121 ) , .ZN( u1_u0_u4_n122 ) , .A2( u1_u0_u4_n144 ) , .A1( u1_u0_u4_n154 ) );
  INV_X1 u1_u0_u5_U10 (.A( u1_u0_u5_n121 ) , .ZN( u1_u0_u5_n177 ) );
  NOR3_X1 u1_u0_u5_U100 (.A3( u1_u0_u5_n141 ) , .A1( u1_u0_u5_n142 ) , .ZN( u1_u0_u5_n143 ) , .A2( u1_u0_u5_n191 ) );
  NAND4_X1 u1_u0_u5_U101 (.ZN( u1_out0_4 ) , .A4( u1_u0_u5_n112 ) , .A2( u1_u0_u5_n113 ) , .A1( u1_u0_u5_n114 ) , .A3( u1_u0_u5_n195 ) );
  AOI211_X1 u1_u0_u5_U102 (.A( u1_u0_u5_n110 ) , .C1( u1_u0_u5_n111 ) , .ZN( u1_u0_u5_n112 ) , .B( u1_u0_u5_n118 ) , .C2( u1_u0_u5_n177 ) );
  AOI222_X1 u1_u0_u5_U103 (.ZN( u1_u0_u5_n113 ) , .A1( u1_u0_u5_n131 ) , .C1( u1_u0_u5_n148 ) , .B2( u1_u0_u5_n174 ) , .C2( u1_u0_u5_n178 ) , .A2( u1_u0_u5_n179 ) , .B1( u1_u0_u5_n99 ) );
  NAND3_X1 u1_u0_u5_U104 (.A2( u1_u0_u5_n154 ) , .A3( u1_u0_u5_n158 ) , .A1( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n99 ) );
  NOR2_X1 u1_u0_u5_U11 (.ZN( u1_u0_u5_n160 ) , .A2( u1_u0_u5_n173 ) , .A1( u1_u0_u5_n177 ) );
  INV_X1 u1_u0_u5_U12 (.A( u1_u0_u5_n150 ) , .ZN( u1_u0_u5_n174 ) );
  AOI21_X1 u1_u0_u5_U13 (.A( u1_u0_u5_n160 ) , .B2( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n162 ) , .B1( u1_u0_u5_n192 ) );
  INV_X1 u1_u0_u5_U14 (.A( u1_u0_u5_n159 ) , .ZN( u1_u0_u5_n192 ) );
  AOI21_X1 u1_u0_u5_U15 (.A( u1_u0_u5_n156 ) , .B2( u1_u0_u5_n157 ) , .B1( u1_u0_u5_n158 ) , .ZN( u1_u0_u5_n163 ) );
  AOI21_X1 u1_u0_u5_U16 (.B2( u1_u0_u5_n139 ) , .B1( u1_u0_u5_n140 ) , .ZN( u1_u0_u5_n141 ) , .A( u1_u0_u5_n150 ) );
  OAI21_X1 u1_u0_u5_U17 (.A( u1_u0_u5_n133 ) , .B2( u1_u0_u5_n134 ) , .B1( u1_u0_u5_n135 ) , .ZN( u1_u0_u5_n142 ) );
  OAI21_X1 u1_u0_u5_U18 (.ZN( u1_u0_u5_n133 ) , .B2( u1_u0_u5_n147 ) , .A( u1_u0_u5_n173 ) , .B1( u1_u0_u5_n188 ) );
  NAND2_X1 u1_u0_u5_U19 (.A2( u1_u0_u5_n119 ) , .A1( u1_u0_u5_n123 ) , .ZN( u1_u0_u5_n137 ) );
  INV_X1 u1_u0_u5_U20 (.A( u1_u0_u5_n155 ) , .ZN( u1_u0_u5_n194 ) );
  NAND2_X1 u1_u0_u5_U21 (.A1( u1_u0_u5_n121 ) , .ZN( u1_u0_u5_n132 ) , .A2( u1_u0_u5_n172 ) );
  NAND2_X1 u1_u0_u5_U22 (.A2( u1_u0_u5_n122 ) , .ZN( u1_u0_u5_n136 ) , .A1( u1_u0_u5_n154 ) );
  NAND2_X1 u1_u0_u5_U23 (.A2( u1_u0_u5_n119 ) , .A1( u1_u0_u5_n120 ) , .ZN( u1_u0_u5_n159 ) );
  INV_X1 u1_u0_u5_U24 (.A( u1_u0_u5_n156 ) , .ZN( u1_u0_u5_n175 ) );
  INV_X1 u1_u0_u5_U25 (.A( u1_u0_u5_n158 ) , .ZN( u1_u0_u5_n188 ) );
  INV_X1 u1_u0_u5_U26 (.A( u1_u0_u5_n152 ) , .ZN( u1_u0_u5_n179 ) );
  INV_X1 u1_u0_u5_U27 (.A( u1_u0_u5_n140 ) , .ZN( u1_u0_u5_n182 ) );
  INV_X1 u1_u0_u5_U28 (.A( u1_u0_u5_n151 ) , .ZN( u1_u0_u5_n183 ) );
  INV_X1 u1_u0_u5_U29 (.A( u1_u0_u5_n123 ) , .ZN( u1_u0_u5_n185 ) );
  NOR2_X1 u1_u0_u5_U3 (.ZN( u1_u0_u5_n134 ) , .A1( u1_u0_u5_n183 ) , .A2( u1_u0_u5_n190 ) );
  INV_X1 u1_u0_u5_U30 (.A( u1_u0_u5_n161 ) , .ZN( u1_u0_u5_n184 ) );
  INV_X1 u1_u0_u5_U31 (.A( u1_u0_u5_n139 ) , .ZN( u1_u0_u5_n189 ) );
  INV_X1 u1_u0_u5_U32 (.A( u1_u0_u5_n157 ) , .ZN( u1_u0_u5_n190 ) );
  INV_X1 u1_u0_u5_U33 (.A( u1_u0_u5_n120 ) , .ZN( u1_u0_u5_n193 ) );
  NAND2_X1 u1_u0_u5_U34 (.ZN( u1_u0_u5_n111 ) , .A1( u1_u0_u5_n140 ) , .A2( u1_u0_u5_n155 ) );
  INV_X1 u1_u0_u5_U35 (.A( u1_u0_u5_n117 ) , .ZN( u1_u0_u5_n196 ) );
  OAI221_X1 u1_u0_u5_U36 (.A( u1_u0_u5_n116 ) , .ZN( u1_u0_u5_n117 ) , .B2( u1_u0_u5_n119 ) , .C1( u1_u0_u5_n153 ) , .C2( u1_u0_u5_n158 ) , .B1( u1_u0_u5_n172 ) );
  AOI222_X1 u1_u0_u5_U37 (.ZN( u1_u0_u5_n116 ) , .B2( u1_u0_u5_n145 ) , .C1( u1_u0_u5_n148 ) , .A2( u1_u0_u5_n174 ) , .C2( u1_u0_u5_n177 ) , .B1( u1_u0_u5_n187 ) , .A1( u1_u0_u5_n193 ) );
  INV_X1 u1_u0_u5_U38 (.A( u1_u0_u5_n115 ) , .ZN( u1_u0_u5_n187 ) );
  NOR2_X1 u1_u0_u5_U39 (.ZN( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n170 ) , .A2( u1_u0_u5_n180 ) );
  INV_X1 u1_u0_u5_U4 (.A( u1_u0_u5_n138 ) , .ZN( u1_u0_u5_n191 ) );
  AOI22_X1 u1_u0_u5_U40 (.B2( u1_u0_u5_n131 ) , .A2( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n169 ) , .B1( u1_u0_u5_n174 ) , .A1( u1_u0_u5_n185 ) );
  NOR2_X1 u1_u0_u5_U41 (.A1( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n150 ) , .A2( u1_u0_u5_n173 ) );
  AOI21_X1 u1_u0_u5_U42 (.A( u1_u0_u5_n118 ) , .B2( u1_u0_u5_n145 ) , .ZN( u1_u0_u5_n168 ) , .B1( u1_u0_u5_n186 ) );
  INV_X1 u1_u0_u5_U43 (.A( u1_u0_u5_n122 ) , .ZN( u1_u0_u5_n186 ) );
  NOR2_X1 u1_u0_u5_U44 (.A1( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n152 ) , .A2( u1_u0_u5_n176 ) );
  NOR2_X1 u1_u0_u5_U45 (.A1( u1_u0_u5_n115 ) , .ZN( u1_u0_u5_n118 ) , .A2( u1_u0_u5_n153 ) );
  NOR2_X1 u1_u0_u5_U46 (.A2( u1_u0_u5_n145 ) , .ZN( u1_u0_u5_n156 ) , .A1( u1_u0_u5_n174 ) );
  NOR2_X1 u1_u0_u5_U47 (.ZN( u1_u0_u5_n121 ) , .A2( u1_u0_u5_n145 ) , .A1( u1_u0_u5_n176 ) );
  AOI22_X1 u1_u0_u5_U48 (.ZN( u1_u0_u5_n114 ) , .A2( u1_u0_u5_n137 ) , .A1( u1_u0_u5_n145 ) , .B2( u1_u0_u5_n175 ) , .B1( u1_u0_u5_n193 ) );
  OAI211_X1 u1_u0_u5_U49 (.B( u1_u0_u5_n124 ) , .A( u1_u0_u5_n125 ) , .C2( u1_u0_u5_n126 ) , .C1( u1_u0_u5_n127 ) , .ZN( u1_u0_u5_n128 ) );
  OAI21_X1 u1_u0_u5_U5 (.B2( u1_u0_u5_n136 ) , .B1( u1_u0_u5_n137 ) , .ZN( u1_u0_u5_n138 ) , .A( u1_u0_u5_n177 ) );
  NOR3_X1 u1_u0_u5_U50 (.ZN( u1_u0_u5_n127 ) , .A1( u1_u0_u5_n136 ) , .A3( u1_u0_u5_n148 ) , .A2( u1_u0_u5_n182 ) );
  OAI21_X1 u1_u0_u5_U51 (.ZN( u1_u0_u5_n124 ) , .A( u1_u0_u5_n177 ) , .B2( u1_u0_u5_n183 ) , .B1( u1_u0_u5_n189 ) );
  OAI21_X1 u1_u0_u5_U52 (.ZN( u1_u0_u5_n125 ) , .A( u1_u0_u5_n174 ) , .B2( u1_u0_u5_n185 ) , .B1( u1_u0_u5_n190 ) );
  AOI21_X1 u1_u0_u5_U53 (.A( u1_u0_u5_n153 ) , .B2( u1_u0_u5_n154 ) , .B1( u1_u0_u5_n155 ) , .ZN( u1_u0_u5_n164 ) );
  AOI21_X1 u1_u0_u5_U54 (.ZN( u1_u0_u5_n110 ) , .B1( u1_u0_u5_n122 ) , .B2( u1_u0_u5_n139 ) , .A( u1_u0_u5_n153 ) );
  INV_X1 u1_u0_u5_U55 (.A( u1_u0_u5_n153 ) , .ZN( u1_u0_u5_n176 ) );
  INV_X1 u1_u0_u5_U56 (.A( u1_u0_u5_n126 ) , .ZN( u1_u0_u5_n173 ) );
  AND2_X1 u1_u0_u5_U57 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n147 ) );
  AND2_X1 u1_u0_u5_U58 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n148 ) );
  NAND2_X1 u1_u0_u5_U59 (.A1( u1_u0_u5_n105 ) , .A2( u1_u0_u5_n106 ) , .ZN( u1_u0_u5_n158 ) );
  INV_X1 u1_u0_u5_U6 (.A( u1_u0_u5_n135 ) , .ZN( u1_u0_u5_n178 ) );
  NAND2_X1 u1_u0_u5_U60 (.A2( u1_u0_u5_n108 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n139 ) );
  NAND2_X1 u1_u0_u5_U61 (.A1( u1_u0_u5_n106 ) , .A2( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n119 ) );
  NAND2_X1 u1_u0_u5_U62 (.A2( u1_u0_u5_n103 ) , .A1( u1_u0_u5_n105 ) , .ZN( u1_u0_u5_n140 ) );
  NAND2_X1 u1_u0_u5_U63 (.A2( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n105 ) , .ZN( u1_u0_u5_n155 ) );
  NAND2_X1 u1_u0_u5_U64 (.A2( u1_u0_u5_n106 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n122 ) );
  NAND2_X1 u1_u0_u5_U65 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n106 ) , .ZN( u1_u0_u5_n115 ) );
  NAND2_X1 u1_u0_u5_U66 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n103 ) , .ZN( u1_u0_u5_n161 ) );
  NAND2_X1 u1_u0_u5_U67 (.A1( u1_u0_u5_n105 ) , .A2( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n154 ) );
  INV_X1 u1_u0_u5_U68 (.A( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n172 ) );
  NAND2_X1 u1_u0_u5_U69 (.A1( u1_u0_u5_n103 ) , .A2( u1_u0_u5_n108 ) , .ZN( u1_u0_u5_n123 ) );
  OAI22_X1 u1_u0_u5_U7 (.B2( u1_u0_u5_n149 ) , .B1( u1_u0_u5_n150 ) , .A2( u1_u0_u5_n151 ) , .A1( u1_u0_u5_n152 ) , .ZN( u1_u0_u5_n165 ) );
  NAND2_X1 u1_u0_u5_U70 (.A2( u1_u0_u5_n103 ) , .A1( u1_u0_u5_n107 ) , .ZN( u1_u0_u5_n151 ) );
  NAND2_X1 u1_u0_u5_U71 (.A2( u1_u0_u5_n107 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n120 ) );
  NAND2_X1 u1_u0_u5_U72 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n109 ) , .ZN( u1_u0_u5_n157 ) );
  AND2_X1 u1_u0_u5_U73 (.A2( u1_u0_u5_n100 ) , .A1( u1_u0_u5_n104 ) , .ZN( u1_u0_u5_n131 ) );
  INV_X1 u1_u0_u5_U74 (.A( u1_u0_u5_n102 ) , .ZN( u1_u0_u5_n195 ) );
  OAI221_X1 u1_u0_u5_U75 (.A( u1_u0_u5_n101 ) , .ZN( u1_u0_u5_n102 ) , .C2( u1_u0_u5_n115 ) , .C1( u1_u0_u5_n126 ) , .B1( u1_u0_u5_n134 ) , .B2( u1_u0_u5_n160 ) );
  OAI21_X1 u1_u0_u5_U76 (.ZN( u1_u0_u5_n101 ) , .B1( u1_u0_u5_n137 ) , .A( u1_u0_u5_n146 ) , .B2( u1_u0_u5_n147 ) );
  NOR2_X1 u1_u0_u5_U77 (.A2( u1_u0_X_34 ) , .A1( u1_u0_X_35 ) , .ZN( u1_u0_u5_n145 ) );
  NOR2_X1 u1_u0_u5_U78 (.A2( u1_u0_X_34 ) , .ZN( u1_u0_u5_n146 ) , .A1( u1_u0_u5_n171 ) );
  NOR2_X1 u1_u0_u5_U79 (.A2( u1_u0_X_31 ) , .A1( u1_u0_X_32 ) , .ZN( u1_u0_u5_n103 ) );
  NOR3_X1 u1_u0_u5_U8 (.A2( u1_u0_u5_n147 ) , .A1( u1_u0_u5_n148 ) , .ZN( u1_u0_u5_n149 ) , .A3( u1_u0_u5_n194 ) );
  NOR2_X1 u1_u0_u5_U80 (.A2( u1_u0_X_36 ) , .ZN( u1_u0_u5_n105 ) , .A1( u1_u0_u5_n180 ) );
  NOR2_X1 u1_u0_u5_U81 (.A2( u1_u0_X_33 ) , .ZN( u1_u0_u5_n108 ) , .A1( u1_u0_u5_n170 ) );
  NOR2_X1 u1_u0_u5_U82 (.A2( u1_u0_X_33 ) , .A1( u1_u0_X_36 ) , .ZN( u1_u0_u5_n107 ) );
  NOR2_X1 u1_u0_u5_U83 (.A2( u1_u0_X_31 ) , .ZN( u1_u0_u5_n104 ) , .A1( u1_u0_u5_n181 ) );
  NAND2_X1 u1_u0_u5_U84 (.A2( u1_u0_X_34 ) , .A1( u1_u0_X_35 ) , .ZN( u1_u0_u5_n153 ) );
  NAND2_X1 u1_u0_u5_U85 (.A1( u1_u0_X_34 ) , .ZN( u1_u0_u5_n126 ) , .A2( u1_u0_u5_n171 ) );
  AND2_X1 u1_u0_u5_U86 (.A1( u1_u0_X_31 ) , .A2( u1_u0_X_32 ) , .ZN( u1_u0_u5_n106 ) );
  AND2_X1 u1_u0_u5_U87 (.A1( u1_u0_X_31 ) , .ZN( u1_u0_u5_n109 ) , .A2( u1_u0_u5_n181 ) );
  INV_X1 u1_u0_u5_U88 (.A( u1_u0_X_33 ) , .ZN( u1_u0_u5_n180 ) );
  INV_X1 u1_u0_u5_U89 (.A( u1_u0_X_35 ) , .ZN( u1_u0_u5_n171 ) );
  NOR2_X1 u1_u0_u5_U9 (.ZN( u1_u0_u5_n135 ) , .A1( u1_u0_u5_n173 ) , .A2( u1_u0_u5_n176 ) );
  INV_X1 u1_u0_u5_U90 (.A( u1_u0_X_36 ) , .ZN( u1_u0_u5_n170 ) );
  INV_X1 u1_u0_u5_U91 (.A( u1_u0_X_32 ) , .ZN( u1_u0_u5_n181 ) );
  NAND4_X1 u1_u0_u5_U92 (.ZN( u1_out0_29 ) , .A4( u1_u0_u5_n129 ) , .A3( u1_u0_u5_n130 ) , .A2( u1_u0_u5_n168 ) , .A1( u1_u0_u5_n196 ) );
  AOI221_X1 u1_u0_u5_U93 (.A( u1_u0_u5_n128 ) , .ZN( u1_u0_u5_n129 ) , .C2( u1_u0_u5_n132 ) , .B2( u1_u0_u5_n159 ) , .B1( u1_u0_u5_n176 ) , .C1( u1_u0_u5_n184 ) );
  AOI222_X1 u1_u0_u5_U94 (.ZN( u1_u0_u5_n130 ) , .A2( u1_u0_u5_n146 ) , .B1( u1_u0_u5_n147 ) , .C2( u1_u0_u5_n175 ) , .B2( u1_u0_u5_n179 ) , .A1( u1_u0_u5_n188 ) , .C1( u1_u0_u5_n194 ) );
  NAND4_X1 u1_u0_u5_U95 (.ZN( u1_out0_19 ) , .A4( u1_u0_u5_n166 ) , .A3( u1_u0_u5_n167 ) , .A2( u1_u0_u5_n168 ) , .A1( u1_u0_u5_n169 ) );
  AOI22_X1 u1_u0_u5_U96 (.B2( u1_u0_u5_n145 ) , .A2( u1_u0_u5_n146 ) , .ZN( u1_u0_u5_n167 ) , .B1( u1_u0_u5_n182 ) , .A1( u1_u0_u5_n189 ) );
  NOR4_X1 u1_u0_u5_U97 (.A4( u1_u0_u5_n162 ) , .A3( u1_u0_u5_n163 ) , .A2( u1_u0_u5_n164 ) , .A1( u1_u0_u5_n165 ) , .ZN( u1_u0_u5_n166 ) );
  NAND4_X1 u1_u0_u5_U98 (.ZN( u1_out0_11 ) , .A4( u1_u0_u5_n143 ) , .A3( u1_u0_u5_n144 ) , .A2( u1_u0_u5_n169 ) , .A1( u1_u0_u5_n196 ) );
  AOI22_X1 u1_u0_u5_U99 (.A2( u1_u0_u5_n132 ) , .ZN( u1_u0_u5_n144 ) , .B2( u1_u0_u5_n145 ) , .B1( u1_u0_u5_n184 ) , .A1( u1_u0_u5_n194 ) );
  AOI22_X1 u1_u0_u6_U10 (.A2( u1_u0_u6_n151 ) , .B2( u1_u0_u6_n161 ) , .A1( u1_u0_u6_n167 ) , .B1( u1_u0_u6_n170 ) , .ZN( u1_u0_u6_n89 ) );
  AOI21_X1 u1_u0_u6_U11 (.B1( u1_u0_u6_n107 ) , .B2( u1_u0_u6_n132 ) , .A( u1_u0_u6_n158 ) , .ZN( u1_u0_u6_n88 ) );
  AOI21_X1 u1_u0_u6_U12 (.B2( u1_u0_u6_n147 ) , .B1( u1_u0_u6_n148 ) , .ZN( u1_u0_u6_n149 ) , .A( u1_u0_u6_n158 ) );
  AOI21_X1 u1_u0_u6_U13 (.ZN( u1_u0_u6_n106 ) , .A( u1_u0_u6_n142 ) , .B2( u1_u0_u6_n159 ) , .B1( u1_u0_u6_n164 ) );
  INV_X1 u1_u0_u6_U14 (.A( u1_u0_u6_n155 ) , .ZN( u1_u0_u6_n161 ) );
  INV_X1 u1_u0_u6_U15 (.A( u1_u0_u6_n128 ) , .ZN( u1_u0_u6_n164 ) );
  NAND2_X1 u1_u0_u6_U16 (.ZN( u1_u0_u6_n110 ) , .A1( u1_u0_u6_n122 ) , .A2( u1_u0_u6_n129 ) );
  NAND2_X1 u1_u0_u6_U17 (.ZN( u1_u0_u6_n124 ) , .A2( u1_u0_u6_n146 ) , .A1( u1_u0_u6_n148 ) );
  INV_X1 u1_u0_u6_U18 (.A( u1_u0_u6_n132 ) , .ZN( u1_u0_u6_n171 ) );
  AND2_X1 u1_u0_u6_U19 (.A1( u1_u0_u6_n100 ) , .ZN( u1_u0_u6_n130 ) , .A2( u1_u0_u6_n147 ) );
  INV_X1 u1_u0_u6_U20 (.A( u1_u0_u6_n127 ) , .ZN( u1_u0_u6_n173 ) );
  INV_X1 u1_u0_u6_U21 (.A( u1_u0_u6_n121 ) , .ZN( u1_u0_u6_n167 ) );
  INV_X1 u1_u0_u6_U22 (.A( u1_u0_u6_n100 ) , .ZN( u1_u0_u6_n169 ) );
  INV_X1 u1_u0_u6_U23 (.A( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n170 ) );
  INV_X1 u1_u0_u6_U24 (.A( u1_u0_u6_n113 ) , .ZN( u1_u0_u6_n168 ) );
  AND2_X1 u1_u0_u6_U25 (.A1( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n119 ) , .ZN( u1_u0_u6_n133 ) );
  AND2_X1 u1_u0_u6_U26 (.A2( u1_u0_u6_n121 ) , .A1( u1_u0_u6_n122 ) , .ZN( u1_u0_u6_n131 ) );
  AND3_X1 u1_u0_u6_U27 (.ZN( u1_u0_u6_n120 ) , .A2( u1_u0_u6_n127 ) , .A1( u1_u0_u6_n132 ) , .A3( u1_u0_u6_n145 ) );
  INV_X1 u1_u0_u6_U28 (.A( u1_u0_u6_n146 ) , .ZN( u1_u0_u6_n163 ) );
  AOI222_X1 u1_u0_u6_U29 (.ZN( u1_u0_u6_n114 ) , .A1( u1_u0_u6_n118 ) , .A2( u1_u0_u6_n126 ) , .B2( u1_u0_u6_n151 ) , .C2( u1_u0_u6_n159 ) , .C1( u1_u0_u6_n168 ) , .B1( u1_u0_u6_n169 ) );
  INV_X1 u1_u0_u6_U3 (.A( u1_u0_u6_n110 ) , .ZN( u1_u0_u6_n166 ) );
  NOR2_X1 u1_u0_u6_U30 (.A1( u1_u0_u6_n162 ) , .A2( u1_u0_u6_n165 ) , .ZN( u1_u0_u6_n98 ) );
  AOI211_X1 u1_u0_u6_U31 (.B( u1_u0_u6_n134 ) , .A( u1_u0_u6_n135 ) , .C1( u1_u0_u6_n136 ) , .ZN( u1_u0_u6_n137 ) , .C2( u1_u0_u6_n151 ) );
  AOI21_X1 u1_u0_u6_U32 (.B2( u1_u0_u6_n132 ) , .B1( u1_u0_u6_n133 ) , .ZN( u1_u0_u6_n134 ) , .A( u1_u0_u6_n158 ) );
  NAND4_X1 u1_u0_u6_U33 (.A4( u1_u0_u6_n127 ) , .A3( u1_u0_u6_n128 ) , .A2( u1_u0_u6_n129 ) , .A1( u1_u0_u6_n130 ) , .ZN( u1_u0_u6_n136 ) );
  AOI21_X1 u1_u0_u6_U34 (.B1( u1_u0_u6_n131 ) , .ZN( u1_u0_u6_n135 ) , .A( u1_u0_u6_n144 ) , .B2( u1_u0_u6_n146 ) );
  NAND2_X1 u1_u0_u6_U35 (.A1( u1_u0_u6_n144 ) , .ZN( u1_u0_u6_n151 ) , .A2( u1_u0_u6_n158 ) );
  NAND2_X1 u1_u0_u6_U36 (.ZN( u1_u0_u6_n132 ) , .A1( u1_u0_u6_n91 ) , .A2( u1_u0_u6_n97 ) );
  AOI22_X1 u1_u0_u6_U37 (.B2( u1_u0_u6_n110 ) , .B1( u1_u0_u6_n111 ) , .A1( u1_u0_u6_n112 ) , .ZN( u1_u0_u6_n115 ) , .A2( u1_u0_u6_n161 ) );
  NAND4_X1 u1_u0_u6_U38 (.A3( u1_u0_u6_n109 ) , .ZN( u1_u0_u6_n112 ) , .A4( u1_u0_u6_n132 ) , .A2( u1_u0_u6_n147 ) , .A1( u1_u0_u6_n166 ) );
  NOR2_X1 u1_u0_u6_U39 (.ZN( u1_u0_u6_n109 ) , .A1( u1_u0_u6_n170 ) , .A2( u1_u0_u6_n173 ) );
  INV_X1 u1_u0_u6_U4 (.A( u1_u0_u6_n142 ) , .ZN( u1_u0_u6_n174 ) );
  NOR2_X1 u1_u0_u6_U40 (.A2( u1_u0_u6_n126 ) , .ZN( u1_u0_u6_n155 ) , .A1( u1_u0_u6_n160 ) );
  NAND2_X1 u1_u0_u6_U41 (.ZN( u1_u0_u6_n146 ) , .A2( u1_u0_u6_n94 ) , .A1( u1_u0_u6_n99 ) );
  AOI21_X1 u1_u0_u6_U42 (.A( u1_u0_u6_n144 ) , .B2( u1_u0_u6_n145 ) , .B1( u1_u0_u6_n146 ) , .ZN( u1_u0_u6_n150 ) );
  INV_X1 u1_u0_u6_U43 (.A( u1_u0_u6_n111 ) , .ZN( u1_u0_u6_n158 ) );
  NAND2_X1 u1_u0_u6_U44 (.ZN( u1_u0_u6_n127 ) , .A1( u1_u0_u6_n91 ) , .A2( u1_u0_u6_n92 ) );
  NAND2_X1 u1_u0_u6_U45 (.ZN( u1_u0_u6_n129 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n96 ) );
  INV_X1 u1_u0_u6_U46 (.A( u1_u0_u6_n144 ) , .ZN( u1_u0_u6_n159 ) );
  NAND2_X1 u1_u0_u6_U47 (.ZN( u1_u0_u6_n145 ) , .A2( u1_u0_u6_n97 ) , .A1( u1_u0_u6_n98 ) );
  NAND2_X1 u1_u0_u6_U48 (.ZN( u1_u0_u6_n148 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n94 ) );
  NAND2_X1 u1_u0_u6_U49 (.ZN( u1_u0_u6_n108 ) , .A2( u1_u0_u6_n139 ) , .A1( u1_u0_u6_n144 ) );
  NAND2_X1 u1_u0_u6_U5 (.A2( u1_u0_u6_n143 ) , .ZN( u1_u0_u6_n152 ) , .A1( u1_u0_u6_n166 ) );
  NAND2_X1 u1_u0_u6_U50 (.ZN( u1_u0_u6_n121 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n97 ) );
  NAND2_X1 u1_u0_u6_U51 (.ZN( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n95 ) );
  AND2_X1 u1_u0_u6_U52 (.ZN( u1_u0_u6_n118 ) , .A2( u1_u0_u6_n91 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U53 (.ZN( u1_u0_u6_n147 ) , .A2( u1_u0_u6_n98 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U54 (.ZN( u1_u0_u6_n128 ) , .A1( u1_u0_u6_n94 ) , .A2( u1_u0_u6_n96 ) );
  NAND2_X1 u1_u0_u6_U55 (.ZN( u1_u0_u6_n119 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U56 (.ZN( u1_u0_u6_n123 ) , .A2( u1_u0_u6_n91 ) , .A1( u1_u0_u6_n96 ) );
  NAND2_X1 u1_u0_u6_U57 (.ZN( u1_u0_u6_n100 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n98 ) );
  NAND2_X1 u1_u0_u6_U58 (.ZN( u1_u0_u6_n122 ) , .A1( u1_u0_u6_n94 ) , .A2( u1_u0_u6_n97 ) );
  INV_X1 u1_u0_u6_U59 (.A( u1_u0_u6_n139 ) , .ZN( u1_u0_u6_n160 ) );
  AOI22_X1 u1_u0_u6_U6 (.B2( u1_u0_u6_n101 ) , .A1( u1_u0_u6_n102 ) , .ZN( u1_u0_u6_n103 ) , .B1( u1_u0_u6_n160 ) , .A2( u1_u0_u6_n161 ) );
  NAND2_X1 u1_u0_u6_U60 (.ZN( u1_u0_u6_n113 ) , .A1( u1_u0_u6_n96 ) , .A2( u1_u0_u6_n98 ) );
  NOR2_X1 u1_u0_u6_U61 (.A2( u1_u0_X_40 ) , .A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n126 ) );
  NOR2_X1 u1_u0_u6_U62 (.A2( u1_u0_X_39 ) , .A1( u1_u0_X_42 ) , .ZN( u1_u0_u6_n92 ) );
  NOR2_X1 u1_u0_u6_U63 (.A2( u1_u0_X_39 ) , .A1( u1_u0_u6_n156 ) , .ZN( u1_u0_u6_n97 ) );
  NOR2_X1 u1_u0_u6_U64 (.A2( u1_u0_X_38 ) , .A1( u1_u0_u6_n165 ) , .ZN( u1_u0_u6_n95 ) );
  NOR2_X1 u1_u0_u6_U65 (.A2( u1_u0_X_41 ) , .ZN( u1_u0_u6_n111 ) , .A1( u1_u0_u6_n157 ) );
  NOR2_X1 u1_u0_u6_U66 (.A2( u1_u0_X_37 ) , .A1( u1_u0_u6_n162 ) , .ZN( u1_u0_u6_n94 ) );
  NOR2_X1 u1_u0_u6_U67 (.A2( u1_u0_X_37 ) , .A1( u1_u0_X_38 ) , .ZN( u1_u0_u6_n91 ) );
  NAND2_X1 u1_u0_u6_U68 (.A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n144 ) , .A2( u1_u0_u6_n157 ) );
  NAND2_X1 u1_u0_u6_U69 (.A2( u1_u0_X_40 ) , .A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n139 ) );
  NOR2_X1 u1_u0_u6_U7 (.A1( u1_u0_u6_n118 ) , .ZN( u1_u0_u6_n143 ) , .A2( u1_u0_u6_n168 ) );
  AND2_X1 u1_u0_u6_U70 (.A1( u1_u0_X_39 ) , .A2( u1_u0_u6_n156 ) , .ZN( u1_u0_u6_n96 ) );
  AND2_X1 u1_u0_u6_U71 (.A1( u1_u0_X_39 ) , .A2( u1_u0_X_42 ) , .ZN( u1_u0_u6_n99 ) );
  INV_X1 u1_u0_u6_U72 (.A( u1_u0_X_40 ) , .ZN( u1_u0_u6_n157 ) );
  INV_X1 u1_u0_u6_U73 (.A( u1_u0_X_37 ) , .ZN( u1_u0_u6_n165 ) );
  INV_X1 u1_u0_u6_U74 (.A( u1_u0_X_38 ) , .ZN( u1_u0_u6_n162 ) );
  INV_X1 u1_u0_u6_U75 (.A( u1_u0_X_42 ) , .ZN( u1_u0_u6_n156 ) );
  NAND4_X1 u1_u0_u6_U76 (.ZN( u1_out0_32 ) , .A4( u1_u0_u6_n103 ) , .A3( u1_u0_u6_n104 ) , .A2( u1_u0_u6_n105 ) , .A1( u1_u0_u6_n106 ) );
  AOI22_X1 u1_u0_u6_U77 (.ZN( u1_u0_u6_n105 ) , .A2( u1_u0_u6_n108 ) , .A1( u1_u0_u6_n118 ) , .B2( u1_u0_u6_n126 ) , .B1( u1_u0_u6_n171 ) );
  AOI22_X1 u1_u0_u6_U78 (.ZN( u1_u0_u6_n104 ) , .A1( u1_u0_u6_n111 ) , .B1( u1_u0_u6_n124 ) , .B2( u1_u0_u6_n151 ) , .A2( u1_u0_u6_n93 ) );
  NAND4_X1 u1_u0_u6_U79 (.ZN( u1_out0_12 ) , .A4( u1_u0_u6_n114 ) , .A3( u1_u0_u6_n115 ) , .A2( u1_u0_u6_n116 ) , .A1( u1_u0_u6_n117 ) );
  OAI21_X1 u1_u0_u6_U8 (.A( u1_u0_u6_n159 ) , .B1( u1_u0_u6_n169 ) , .B2( u1_u0_u6_n173 ) , .ZN( u1_u0_u6_n90 ) );
  OAI22_X1 u1_u0_u6_U80 (.B2( u1_u0_u6_n111 ) , .ZN( u1_u0_u6_n116 ) , .B1( u1_u0_u6_n126 ) , .A2( u1_u0_u6_n164 ) , .A1( u1_u0_u6_n167 ) );
  OAI21_X1 u1_u0_u6_U81 (.A( u1_u0_u6_n108 ) , .ZN( u1_u0_u6_n117 ) , .B2( u1_u0_u6_n141 ) , .B1( u1_u0_u6_n163 ) );
  OAI211_X1 u1_u0_u6_U82 (.ZN( u1_out0_7 ) , .B( u1_u0_u6_n153 ) , .C2( u1_u0_u6_n154 ) , .C1( u1_u0_u6_n155 ) , .A( u1_u0_u6_n174 ) );
  NOR3_X1 u1_u0_u6_U83 (.A1( u1_u0_u6_n141 ) , .ZN( u1_u0_u6_n154 ) , .A3( u1_u0_u6_n164 ) , .A2( u1_u0_u6_n171 ) );
  AOI211_X1 u1_u0_u6_U84 (.B( u1_u0_u6_n149 ) , .A( u1_u0_u6_n150 ) , .C2( u1_u0_u6_n151 ) , .C1( u1_u0_u6_n152 ) , .ZN( u1_u0_u6_n153 ) );
  OAI211_X1 u1_u0_u6_U85 (.ZN( u1_out0_22 ) , .B( u1_u0_u6_n137 ) , .A( u1_u0_u6_n138 ) , .C2( u1_u0_u6_n139 ) , .C1( u1_u0_u6_n140 ) );
  AOI22_X1 u1_u0_u6_U86 (.B1( u1_u0_u6_n124 ) , .A2( u1_u0_u6_n125 ) , .A1( u1_u0_u6_n126 ) , .ZN( u1_u0_u6_n138 ) , .B2( u1_u0_u6_n161 ) );
  AND4_X1 u1_u0_u6_U87 (.A3( u1_u0_u6_n119 ) , .A1( u1_u0_u6_n120 ) , .A4( u1_u0_u6_n129 ) , .ZN( u1_u0_u6_n140 ) , .A2( u1_u0_u6_n143 ) );
  NAND3_X1 u1_u0_u6_U88 (.A2( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n125 ) , .A1( u1_u0_u6_n130 ) , .A3( u1_u0_u6_n131 ) );
  NAND3_X1 u1_u0_u6_U89 (.A3( u1_u0_u6_n133 ) , .ZN( u1_u0_u6_n141 ) , .A1( u1_u0_u6_n145 ) , .A2( u1_u0_u6_n148 ) );
  INV_X1 u1_u0_u6_U9 (.ZN( u1_u0_u6_n172 ) , .A( u1_u0_u6_n88 ) );
  NAND3_X1 u1_u0_u6_U90 (.ZN( u1_u0_u6_n101 ) , .A3( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n121 ) , .A1( u1_u0_u6_n127 ) );
  NAND3_X1 u1_u0_u6_U91 (.ZN( u1_u0_u6_n102 ) , .A3( u1_u0_u6_n130 ) , .A2( u1_u0_u6_n145 ) , .A1( u1_u0_u6_n166 ) );
  NAND3_X1 u1_u0_u6_U92 (.A3( u1_u0_u6_n113 ) , .A1( u1_u0_u6_n119 ) , .A2( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n93 ) );
  NAND3_X1 u1_u0_u6_U93 (.ZN( u1_u0_u6_n142 ) , .A2( u1_u0_u6_n172 ) , .A3( u1_u0_u6_n89 ) , .A1( u1_u0_u6_n90 ) );
  OAI21_X1 u1_u0_u7_U10 (.A( u1_u0_u7_n161 ) , .B1( u1_u0_u7_n168 ) , .B2( u1_u0_u7_n173 ) , .ZN( u1_u0_u7_n91 ) );
  AOI211_X1 u1_u0_u7_U11 (.A( u1_u0_u7_n117 ) , .ZN( u1_u0_u7_n118 ) , .C2( u1_u0_u7_n126 ) , .C1( u1_u0_u7_n177 ) , .B( u1_u0_u7_n180 ) );
  OAI22_X1 u1_u0_u7_U12 (.B1( u1_u0_u7_n115 ) , .ZN( u1_u0_u7_n117 ) , .A2( u1_u0_u7_n133 ) , .A1( u1_u0_u7_n137 ) , .B2( u1_u0_u7_n162 ) );
  INV_X1 u1_u0_u7_U13 (.A( u1_u0_u7_n116 ) , .ZN( u1_u0_u7_n180 ) );
  NOR3_X1 u1_u0_u7_U14 (.ZN( u1_u0_u7_n115 ) , .A3( u1_u0_u7_n145 ) , .A2( u1_u0_u7_n168 ) , .A1( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U15 (.A( u1_u0_u7_n133 ) , .ZN( u1_u0_u7_n176 ) );
  NOR3_X1 u1_u0_u7_U16 (.A2( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n135 ) , .ZN( u1_u0_u7_n136 ) , .A3( u1_u0_u7_n171 ) );
  NOR2_X1 u1_u0_u7_U17 (.A1( u1_u0_u7_n130 ) , .A2( u1_u0_u7_n134 ) , .ZN( u1_u0_u7_n153 ) );
  AOI21_X1 u1_u0_u7_U18 (.ZN( u1_u0_u7_n104 ) , .B2( u1_u0_u7_n112 ) , .B1( u1_u0_u7_n127 ) , .A( u1_u0_u7_n164 ) );
  AOI21_X1 u1_u0_u7_U19 (.ZN( u1_u0_u7_n106 ) , .B1( u1_u0_u7_n133 ) , .B2( u1_u0_u7_n146 ) , .A( u1_u0_u7_n162 ) );
  AOI21_X1 u1_u0_u7_U20 (.A( u1_u0_u7_n101 ) , .ZN( u1_u0_u7_n107 ) , .B2( u1_u0_u7_n128 ) , .B1( u1_u0_u7_n175 ) );
  INV_X1 u1_u0_u7_U21 (.A( u1_u0_u7_n101 ) , .ZN( u1_u0_u7_n165 ) );
  NOR2_X1 u1_u0_u7_U22 (.ZN( u1_u0_u7_n111 ) , .A2( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U23 (.A( u1_u0_u7_n138 ) , .ZN( u1_u0_u7_n171 ) );
  INV_X1 u1_u0_u7_U24 (.A( u1_u0_u7_n131 ) , .ZN( u1_u0_u7_n177 ) );
  INV_X1 u1_u0_u7_U25 (.A( u1_u0_u7_n110 ) , .ZN( u1_u0_u7_n174 ) );
  NAND2_X1 u1_u0_u7_U26 (.A1( u1_u0_u7_n129 ) , .A2( u1_u0_u7_n132 ) , .ZN( u1_u0_u7_n149 ) );
  NAND2_X1 u1_u0_u7_U27 (.A1( u1_u0_u7_n113 ) , .A2( u1_u0_u7_n124 ) , .ZN( u1_u0_u7_n130 ) );
  INV_X1 u1_u0_u7_U28 (.A( u1_u0_u7_n112 ) , .ZN( u1_u0_u7_n173 ) );
  INV_X1 u1_u0_u7_U29 (.A( u1_u0_u7_n128 ) , .ZN( u1_u0_u7_n168 ) );
  OAI21_X1 u1_u0_u7_U3 (.ZN( u1_u0_u7_n159 ) , .A( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n171 ) , .B1( u1_u0_u7_n174 ) );
  INV_X1 u1_u0_u7_U30 (.A( u1_u0_u7_n148 ) , .ZN( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U31 (.A( u1_u0_u7_n127 ) , .ZN( u1_u0_u7_n179 ) );
  INV_X1 u1_u0_u7_U32 (.A( u1_u0_u7_n153 ) , .ZN( u1_u0_u7_n172 ) );
  NOR2_X1 u1_u0_u7_U33 (.ZN( u1_u0_u7_n101 ) , .A2( u1_u0_u7_n150 ) , .A1( u1_u0_u7_n156 ) );
  AOI211_X1 u1_u0_u7_U34 (.B( u1_u0_u7_n139 ) , .A( u1_u0_u7_n140 ) , .C2( u1_u0_u7_n141 ) , .ZN( u1_u0_u7_n142 ) , .C1( u1_u0_u7_n156 ) );
  NAND4_X1 u1_u0_u7_U35 (.A3( u1_u0_u7_n127 ) , .A2( u1_u0_u7_n128 ) , .A1( u1_u0_u7_n129 ) , .ZN( u1_u0_u7_n141 ) , .A4( u1_u0_u7_n147 ) );
  AOI21_X1 u1_u0_u7_U36 (.A( u1_u0_u7_n137 ) , .B1( u1_u0_u7_n138 ) , .ZN( u1_u0_u7_n139 ) , .B2( u1_u0_u7_n146 ) );
  OAI22_X1 u1_u0_u7_U37 (.B1( u1_u0_u7_n136 ) , .ZN( u1_u0_u7_n140 ) , .A1( u1_u0_u7_n153 ) , .B2( u1_u0_u7_n162 ) , .A2( u1_u0_u7_n164 ) );
  INV_X1 u1_u0_u7_U38 (.A( u1_u0_u7_n125 ) , .ZN( u1_u0_u7_n161 ) );
  AOI21_X1 u1_u0_u7_U39 (.ZN( u1_u0_u7_n123 ) , .B1( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n177 ) , .A( u1_u0_u7_n97 ) );
  INV_X1 u1_u0_u7_U4 (.A( u1_u0_u7_n149 ) , .ZN( u1_u0_u7_n175 ) );
  AOI21_X1 u1_u0_u7_U40 (.B2( u1_u0_u7_n113 ) , .B1( u1_u0_u7_n124 ) , .A( u1_u0_u7_n125 ) , .ZN( u1_u0_u7_n97 ) );
  INV_X1 u1_u0_u7_U41 (.A( u1_u0_u7_n152 ) , .ZN( u1_u0_u7_n162 ) );
  AOI22_X1 u1_u0_u7_U42 (.A2( u1_u0_u7_n114 ) , .ZN( u1_u0_u7_n119 ) , .B1( u1_u0_u7_n130 ) , .A1( u1_u0_u7_n156 ) , .B2( u1_u0_u7_n165 ) );
  NAND2_X1 u1_u0_u7_U43 (.A2( u1_u0_u7_n112 ) , .ZN( u1_u0_u7_n114 ) , .A1( u1_u0_u7_n175 ) );
  NOR2_X1 u1_u0_u7_U44 (.ZN( u1_u0_u7_n137 ) , .A1( u1_u0_u7_n150 ) , .A2( u1_u0_u7_n161 ) );
  AND2_X1 u1_u0_u7_U45 (.ZN( u1_u0_u7_n145 ) , .A2( u1_u0_u7_n98 ) , .A1( u1_u0_u7_n99 ) );
  AOI21_X1 u1_u0_u7_U46 (.ZN( u1_u0_u7_n105 ) , .B2( u1_u0_u7_n110 ) , .A( u1_u0_u7_n125 ) , .B1( u1_u0_u7_n147 ) );
  NAND2_X1 u1_u0_u7_U47 (.ZN( u1_u0_u7_n146 ) , .A1( u1_u0_u7_n95 ) , .A2( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U48 (.A2( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n147 ) , .A1( u1_u0_u7_n93 ) );
  NAND2_X1 u1_u0_u7_U49 (.A1( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n127 ) , .A2( u1_u0_u7_n99 ) );
  INV_X1 u1_u0_u7_U5 (.A( u1_u0_u7_n154 ) , .ZN( u1_u0_u7_n178 ) );
  NAND2_X1 u1_u0_u7_U50 (.A2( u1_u0_u7_n102 ) , .A1( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n133 ) );
  OR2_X1 u1_u0_u7_U51 (.ZN( u1_u0_u7_n126 ) , .A2( u1_u0_u7_n152 ) , .A1( u1_u0_u7_n156 ) );
  NAND2_X1 u1_u0_u7_U52 (.ZN( u1_u0_u7_n112 ) , .A2( u1_u0_u7_n96 ) , .A1( u1_u0_u7_n99 ) );
  NAND2_X1 u1_u0_u7_U53 (.A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n128 ) , .A1( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U54 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n113 ) , .A2( u1_u0_u7_n93 ) );
  NAND2_X1 u1_u0_u7_U55 (.ZN( u1_u0_u7_n110 ) , .A1( u1_u0_u7_n95 ) , .A2( u1_u0_u7_n96 ) );
  INV_X1 u1_u0_u7_U56 (.A( u1_u0_u7_n150 ) , .ZN( u1_u0_u7_n164 ) );
  AND2_X1 u1_u0_u7_U57 (.ZN( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n93 ) , .A2( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U58 (.A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n124 ) , .A1( u1_u0_u7_n96 ) );
  NAND2_X1 u1_u0_u7_U59 (.A1( u1_u0_u7_n100 ) , .A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n129 ) );
  AOI211_X1 u1_u0_u7_U6 (.ZN( u1_u0_u7_n116 ) , .A( u1_u0_u7_n155 ) , .C1( u1_u0_u7_n161 ) , .C2( u1_u0_u7_n171 ) , .B( u1_u0_u7_n94 ) );
  NAND2_X1 u1_u0_u7_U60 (.A2( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n131 ) , .A1( u1_u0_u7_n95 ) );
  NAND2_X1 u1_u0_u7_U61 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n138 ) , .A2( u1_u0_u7_n99 ) );
  NAND2_X1 u1_u0_u7_U62 (.ZN( u1_u0_u7_n132 ) , .A1( u1_u0_u7_n93 ) , .A2( u1_u0_u7_n96 ) );
  NAND2_X1 u1_u0_u7_U63 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n148 ) , .A2( u1_u0_u7_n95 ) );
  NOR2_X1 u1_u0_u7_U64 (.A2( u1_u0_X_47 ) , .ZN( u1_u0_u7_n150 ) , .A1( u1_u0_u7_n163 ) );
  NOR2_X1 u1_u0_u7_U65 (.A2( u1_u0_X_43 ) , .A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n103 ) );
  NOR2_X1 u1_u0_u7_U66 (.A2( u1_u0_X_48 ) , .A1( u1_u0_u7_n166 ) , .ZN( u1_u0_u7_n95 ) );
  NOR2_X1 u1_u0_u7_U67 (.A2( u1_u0_X_45 ) , .A1( u1_u0_X_48 ) , .ZN( u1_u0_u7_n99 ) );
  NOR2_X1 u1_u0_u7_U68 (.A2( u1_u0_X_44 ) , .A1( u1_u0_u7_n167 ) , .ZN( u1_u0_u7_n98 ) );
  NOR2_X1 u1_u0_u7_U69 (.A2( u1_u0_X_46 ) , .A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n152 ) );
  OAI222_X1 u1_u0_u7_U7 (.C2( u1_u0_u7_n101 ) , .B2( u1_u0_u7_n111 ) , .A1( u1_u0_u7_n113 ) , .C1( u1_u0_u7_n146 ) , .A2( u1_u0_u7_n162 ) , .B1( u1_u0_u7_n164 ) , .ZN( u1_u0_u7_n94 ) );
  NAND2_X1 u1_u0_u7_U70 (.A2( u1_u0_X_46 ) , .A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n125 ) );
  AND2_X1 u1_u0_u7_U71 (.A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n156 ) , .A2( u1_u0_u7_n163 ) );
  AND2_X1 u1_u0_u7_U72 (.A2( u1_u0_X_45 ) , .A1( u1_u0_X_48 ) , .ZN( u1_u0_u7_n102 ) );
  AND2_X1 u1_u0_u7_U73 (.A2( u1_u0_X_43 ) , .A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n96 ) );
  AND2_X1 u1_u0_u7_U74 (.A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n100 ) , .A2( u1_u0_u7_n167 ) );
  AND2_X1 u1_u0_u7_U75 (.A1( u1_u0_X_48 ) , .A2( u1_u0_u7_n166 ) , .ZN( u1_u0_u7_n93 ) );
  INV_X1 u1_u0_u7_U76 (.A( u1_u0_X_46 ) , .ZN( u1_u0_u7_n163 ) );
  INV_X1 u1_u0_u7_U77 (.A( u1_u0_X_45 ) , .ZN( u1_u0_u7_n166 ) );
  NAND4_X1 u1_u0_u7_U78 (.ZN( u1_out0_5 ) , .A4( u1_u0_u7_n108 ) , .A3( u1_u0_u7_n109 ) , .A1( u1_u0_u7_n116 ) , .A2( u1_u0_u7_n123 ) );
  AOI22_X1 u1_u0_u7_U79 (.ZN( u1_u0_u7_n109 ) , .A2( u1_u0_u7_n126 ) , .B2( u1_u0_u7_n145 ) , .B1( u1_u0_u7_n156 ) , .A1( u1_u0_u7_n171 ) );
  OAI221_X1 u1_u0_u7_U8 (.C1( u1_u0_u7_n101 ) , .C2( u1_u0_u7_n147 ) , .ZN( u1_u0_u7_n155 ) , .B2( u1_u0_u7_n162 ) , .A( u1_u0_u7_n91 ) , .B1( u1_u0_u7_n92 ) );
  NOR4_X1 u1_u0_u7_U80 (.A4( u1_u0_u7_n104 ) , .A3( u1_u0_u7_n105 ) , .A2( u1_u0_u7_n106 ) , .A1( u1_u0_u7_n107 ) , .ZN( u1_u0_u7_n108 ) );
  NAND4_X1 u1_u0_u7_U81 (.ZN( u1_out0_27 ) , .A4( u1_u0_u7_n118 ) , .A3( u1_u0_u7_n119 ) , .A2( u1_u0_u7_n120 ) , .A1( u1_u0_u7_n121 ) );
  OAI21_X1 u1_u0_u7_U82 (.ZN( u1_u0_u7_n121 ) , .B2( u1_u0_u7_n145 ) , .A( u1_u0_u7_n150 ) , .B1( u1_u0_u7_n174 ) );
  OAI21_X1 u1_u0_u7_U83 (.ZN( u1_u0_u7_n120 ) , .A( u1_u0_u7_n161 ) , .B2( u1_u0_u7_n170 ) , .B1( u1_u0_u7_n179 ) );
  NAND4_X1 u1_u0_u7_U84 (.ZN( u1_out0_21 ) , .A4( u1_u0_u7_n157 ) , .A3( u1_u0_u7_n158 ) , .A2( u1_u0_u7_n159 ) , .A1( u1_u0_u7_n160 ) );
  OAI21_X1 u1_u0_u7_U85 (.B1( u1_u0_u7_n145 ) , .ZN( u1_u0_u7_n160 ) , .A( u1_u0_u7_n161 ) , .B2( u1_u0_u7_n177 ) );
  AOI22_X1 u1_u0_u7_U86 (.B2( u1_u0_u7_n149 ) , .B1( u1_u0_u7_n150 ) , .A2( u1_u0_u7_n151 ) , .A1( u1_u0_u7_n152 ) , .ZN( u1_u0_u7_n158 ) );
  NAND4_X1 u1_u0_u7_U87 (.ZN( u1_out0_15 ) , .A4( u1_u0_u7_n142 ) , .A3( u1_u0_u7_n143 ) , .A2( u1_u0_u7_n144 ) , .A1( u1_u0_u7_n178 ) );
  OR2_X1 u1_u0_u7_U88 (.A2( u1_u0_u7_n125 ) , .A1( u1_u0_u7_n129 ) , .ZN( u1_u0_u7_n144 ) );
  AOI22_X1 u1_u0_u7_U89 (.A2( u1_u0_u7_n126 ) , .ZN( u1_u0_u7_n143 ) , .B2( u1_u0_u7_n165 ) , .B1( u1_u0_u7_n173 ) , .A1( u1_u0_u7_n174 ) );
  AND3_X1 u1_u0_u7_U9 (.A3( u1_u0_u7_n110 ) , .A2( u1_u0_u7_n127 ) , .A1( u1_u0_u7_n132 ) , .ZN( u1_u0_u7_n92 ) );
  INV_X1 u1_u0_u7_U90 (.A( u1_u0_X_43 ) , .ZN( u1_u0_u7_n167 ) );
  AOI211_X1 u1_u0_u7_U91 (.B( u1_u0_u7_n154 ) , .A( u1_u0_u7_n155 ) , .C1( u1_u0_u7_n156 ) , .ZN( u1_u0_u7_n157 ) , .C2( u1_u0_u7_n172 ) );
  OAI211_X1 u1_u0_u7_U92 (.B( u1_u0_u7_n122 ) , .A( u1_u0_u7_n123 ) , .C2( u1_u0_u7_n124 ) , .ZN( u1_u0_u7_n154 ) , .C1( u1_u0_u7_n162 ) );
  AOI222_X1 u1_u0_u7_U93 (.ZN( u1_u0_u7_n122 ) , .C2( u1_u0_u7_n126 ) , .C1( u1_u0_u7_n145 ) , .B1( u1_u0_u7_n161 ) , .A2( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n170 ) , .A1( u1_u0_u7_n176 ) );
  INV_X1 u1_u0_u7_U94 (.A( u1_u0_u7_n111 ) , .ZN( u1_u0_u7_n170 ) );
  NAND3_X1 u1_u0_u7_U95 (.A3( u1_u0_u7_n146 ) , .A2( u1_u0_u7_n147 ) , .A1( u1_u0_u7_n148 ) , .ZN( u1_u0_u7_n151 ) );
  NAND3_X1 u1_u0_u7_U96 (.A3( u1_u0_u7_n131 ) , .A2( u1_u0_u7_n132 ) , .A1( u1_u0_u7_n133 ) , .ZN( u1_u0_u7_n135 ) );
  XOR2_X1 u1_u14_U10 (.B( u1_K15_45 ) , .A( u1_R13_30 ) , .Z( u1_u14_X_45 ) );
  XOR2_X1 u1_u14_U11 (.B( u1_K15_44 ) , .A( u1_R13_29 ) , .Z( u1_u14_X_44 ) );
  XOR2_X1 u1_u14_U12 (.B( u1_K15_43 ) , .A( u1_R13_28 ) , .Z( u1_u14_X_43 ) );
  XOR2_X1 u1_u14_U13 (.B( u1_K15_42 ) , .A( u1_R13_29 ) , .Z( u1_u14_X_42 ) );
  XOR2_X1 u1_u14_U14 (.B( u1_K15_41 ) , .A( u1_R13_28 ) , .Z( u1_u14_X_41 ) );
  XOR2_X1 u1_u14_U15 (.B( u1_K15_40 ) , .A( u1_R13_27 ) , .Z( u1_u14_X_40 ) );
  XOR2_X1 u1_u14_U17 (.B( u1_K15_39 ) , .A( u1_R13_26 ) , .Z( u1_u14_X_39 ) );
  XOR2_X1 u1_u14_U18 (.B( u1_K15_38 ) , .A( u1_R13_25 ) , .Z( u1_u14_X_38 ) );
  XOR2_X1 u1_u14_U19 (.B( u1_K15_37 ) , .A( u1_R13_24 ) , .Z( u1_u14_X_37 ) );
  XOR2_X1 u1_u14_U20 (.B( u1_K15_36 ) , .A( u1_R13_25 ) , .Z( u1_u14_X_36 ) );
  XOR2_X1 u1_u14_U21 (.B( u1_K15_35 ) , .A( u1_R13_24 ) , .Z( u1_u14_X_35 ) );
  XOR2_X1 u1_u14_U22 (.B( u1_K15_34 ) , .A( u1_R13_23 ) , .Z( u1_u14_X_34 ) );
  XOR2_X1 u1_u14_U23 (.B( u1_K15_33 ) , .A( u1_R13_22 ) , .Z( u1_u14_X_33 ) );
  XOR2_X1 u1_u14_U24 (.B( u1_K15_32 ) , .A( u1_R13_21 ) , .Z( u1_u14_X_32 ) );
  XOR2_X1 u1_u14_U25 (.B( u1_K15_31 ) , .A( u1_R13_20 ) , .Z( u1_u14_X_31 ) );
  XOR2_X1 u1_u14_U7 (.B( u1_K15_48 ) , .A( u1_R13_1 ) , .Z( u1_u14_X_48 ) );
  XOR2_X1 u1_u14_U8 (.B( u1_K15_47 ) , .A( u1_R13_32 ) , .Z( u1_u14_X_47 ) );
  XOR2_X1 u1_u14_U9 (.B( u1_K15_46 ) , .A( u1_R13_31 ) , .Z( u1_u14_X_46 ) );
  INV_X1 u1_u14_u5_U10 (.A( u1_u14_u5_n121 ) , .ZN( u1_u14_u5_n177 ) );
  NOR3_X1 u1_u14_u5_U100 (.A3( u1_u14_u5_n141 ) , .A1( u1_u14_u5_n142 ) , .ZN( u1_u14_u5_n143 ) , .A2( u1_u14_u5_n191 ) );
  NAND4_X1 u1_u14_u5_U101 (.ZN( u1_out14_4 ) , .A4( u1_u14_u5_n112 ) , .A2( u1_u14_u5_n113 ) , .A1( u1_u14_u5_n114 ) , .A3( u1_u14_u5_n195 ) );
  AOI211_X1 u1_u14_u5_U102 (.A( u1_u14_u5_n110 ) , .C1( u1_u14_u5_n111 ) , .ZN( u1_u14_u5_n112 ) , .B( u1_u14_u5_n118 ) , .C2( u1_u14_u5_n177 ) );
  AOI222_X1 u1_u14_u5_U103 (.ZN( u1_u14_u5_n113 ) , .A1( u1_u14_u5_n131 ) , .C1( u1_u14_u5_n148 ) , .B2( u1_u14_u5_n174 ) , .C2( u1_u14_u5_n178 ) , .A2( u1_u14_u5_n179 ) , .B1( u1_u14_u5_n99 ) );
  NAND3_X1 u1_u14_u5_U104 (.A2( u1_u14_u5_n154 ) , .A3( u1_u14_u5_n158 ) , .A1( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n99 ) );
  NOR2_X1 u1_u14_u5_U11 (.ZN( u1_u14_u5_n160 ) , .A2( u1_u14_u5_n173 ) , .A1( u1_u14_u5_n177 ) );
  INV_X1 u1_u14_u5_U12 (.A( u1_u14_u5_n150 ) , .ZN( u1_u14_u5_n174 ) );
  AOI21_X1 u1_u14_u5_U13 (.A( u1_u14_u5_n160 ) , .B2( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n162 ) , .B1( u1_u14_u5_n192 ) );
  INV_X1 u1_u14_u5_U14 (.A( u1_u14_u5_n159 ) , .ZN( u1_u14_u5_n192 ) );
  AOI21_X1 u1_u14_u5_U15 (.A( u1_u14_u5_n156 ) , .B2( u1_u14_u5_n157 ) , .B1( u1_u14_u5_n158 ) , .ZN( u1_u14_u5_n163 ) );
  AOI21_X1 u1_u14_u5_U16 (.B2( u1_u14_u5_n139 ) , .B1( u1_u14_u5_n140 ) , .ZN( u1_u14_u5_n141 ) , .A( u1_u14_u5_n150 ) );
  OAI21_X1 u1_u14_u5_U17 (.A( u1_u14_u5_n133 ) , .B2( u1_u14_u5_n134 ) , .B1( u1_u14_u5_n135 ) , .ZN( u1_u14_u5_n142 ) );
  OAI21_X1 u1_u14_u5_U18 (.ZN( u1_u14_u5_n133 ) , .B2( u1_u14_u5_n147 ) , .A( u1_u14_u5_n173 ) , .B1( u1_u14_u5_n188 ) );
  NAND2_X1 u1_u14_u5_U19 (.A2( u1_u14_u5_n119 ) , .A1( u1_u14_u5_n123 ) , .ZN( u1_u14_u5_n137 ) );
  INV_X1 u1_u14_u5_U20 (.A( u1_u14_u5_n155 ) , .ZN( u1_u14_u5_n194 ) );
  NAND2_X1 u1_u14_u5_U21 (.A1( u1_u14_u5_n121 ) , .ZN( u1_u14_u5_n132 ) , .A2( u1_u14_u5_n172 ) );
  NAND2_X1 u1_u14_u5_U22 (.A2( u1_u14_u5_n122 ) , .ZN( u1_u14_u5_n136 ) , .A1( u1_u14_u5_n154 ) );
  NAND2_X1 u1_u14_u5_U23 (.A2( u1_u14_u5_n119 ) , .A1( u1_u14_u5_n120 ) , .ZN( u1_u14_u5_n159 ) );
  INV_X1 u1_u14_u5_U24 (.A( u1_u14_u5_n156 ) , .ZN( u1_u14_u5_n175 ) );
  INV_X1 u1_u14_u5_U25 (.A( u1_u14_u5_n158 ) , .ZN( u1_u14_u5_n188 ) );
  INV_X1 u1_u14_u5_U26 (.A( u1_u14_u5_n152 ) , .ZN( u1_u14_u5_n179 ) );
  INV_X1 u1_u14_u5_U27 (.A( u1_u14_u5_n140 ) , .ZN( u1_u14_u5_n182 ) );
  INV_X1 u1_u14_u5_U28 (.A( u1_u14_u5_n151 ) , .ZN( u1_u14_u5_n183 ) );
  INV_X1 u1_u14_u5_U29 (.A( u1_u14_u5_n123 ) , .ZN( u1_u14_u5_n185 ) );
  NOR2_X1 u1_u14_u5_U3 (.ZN( u1_u14_u5_n134 ) , .A1( u1_u14_u5_n183 ) , .A2( u1_u14_u5_n190 ) );
  INV_X1 u1_u14_u5_U30 (.A( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n184 ) );
  INV_X1 u1_u14_u5_U31 (.A( u1_u14_u5_n139 ) , .ZN( u1_u14_u5_n189 ) );
  INV_X1 u1_u14_u5_U32 (.A( u1_u14_u5_n157 ) , .ZN( u1_u14_u5_n190 ) );
  INV_X1 u1_u14_u5_U33 (.A( u1_u14_u5_n120 ) , .ZN( u1_u14_u5_n193 ) );
  NAND2_X1 u1_u14_u5_U34 (.ZN( u1_u14_u5_n111 ) , .A1( u1_u14_u5_n140 ) , .A2( u1_u14_u5_n155 ) );
  INV_X1 u1_u14_u5_U35 (.A( u1_u14_u5_n117 ) , .ZN( u1_u14_u5_n196 ) );
  OAI221_X1 u1_u14_u5_U36 (.A( u1_u14_u5_n116 ) , .ZN( u1_u14_u5_n117 ) , .B2( u1_u14_u5_n119 ) , .C1( u1_u14_u5_n153 ) , .C2( u1_u14_u5_n158 ) , .B1( u1_u14_u5_n172 ) );
  AOI222_X1 u1_u14_u5_U37 (.ZN( u1_u14_u5_n116 ) , .B2( u1_u14_u5_n145 ) , .C1( u1_u14_u5_n148 ) , .A2( u1_u14_u5_n174 ) , .C2( u1_u14_u5_n177 ) , .B1( u1_u14_u5_n187 ) , .A1( u1_u14_u5_n193 ) );
  INV_X1 u1_u14_u5_U38 (.A( u1_u14_u5_n115 ) , .ZN( u1_u14_u5_n187 ) );
  NOR2_X1 u1_u14_u5_U39 (.ZN( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n170 ) , .A2( u1_u14_u5_n180 ) );
  INV_X1 u1_u14_u5_U4 (.A( u1_u14_u5_n138 ) , .ZN( u1_u14_u5_n191 ) );
  AOI22_X1 u1_u14_u5_U40 (.B2( u1_u14_u5_n131 ) , .A2( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n169 ) , .B1( u1_u14_u5_n174 ) , .A1( u1_u14_u5_n185 ) );
  NOR2_X1 u1_u14_u5_U41 (.A1( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n150 ) , .A2( u1_u14_u5_n173 ) );
  AOI21_X1 u1_u14_u5_U42 (.A( u1_u14_u5_n118 ) , .B2( u1_u14_u5_n145 ) , .ZN( u1_u14_u5_n168 ) , .B1( u1_u14_u5_n186 ) );
  INV_X1 u1_u14_u5_U43 (.A( u1_u14_u5_n122 ) , .ZN( u1_u14_u5_n186 ) );
  NOR2_X1 u1_u14_u5_U44 (.A1( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n152 ) , .A2( u1_u14_u5_n176 ) );
  NOR2_X1 u1_u14_u5_U45 (.A1( u1_u14_u5_n115 ) , .ZN( u1_u14_u5_n118 ) , .A2( u1_u14_u5_n153 ) );
  NOR2_X1 u1_u14_u5_U46 (.A2( u1_u14_u5_n145 ) , .ZN( u1_u14_u5_n156 ) , .A1( u1_u14_u5_n174 ) );
  NOR2_X1 u1_u14_u5_U47 (.ZN( u1_u14_u5_n121 ) , .A2( u1_u14_u5_n145 ) , .A1( u1_u14_u5_n176 ) );
  AOI22_X1 u1_u14_u5_U48 (.ZN( u1_u14_u5_n114 ) , .A2( u1_u14_u5_n137 ) , .A1( u1_u14_u5_n145 ) , .B2( u1_u14_u5_n175 ) , .B1( u1_u14_u5_n193 ) );
  OAI211_X1 u1_u14_u5_U49 (.B( u1_u14_u5_n124 ) , .A( u1_u14_u5_n125 ) , .C2( u1_u14_u5_n126 ) , .C1( u1_u14_u5_n127 ) , .ZN( u1_u14_u5_n128 ) );
  OAI21_X1 u1_u14_u5_U5 (.B2( u1_u14_u5_n136 ) , .B1( u1_u14_u5_n137 ) , .ZN( u1_u14_u5_n138 ) , .A( u1_u14_u5_n177 ) );
  NOR3_X1 u1_u14_u5_U50 (.ZN( u1_u14_u5_n127 ) , .A1( u1_u14_u5_n136 ) , .A3( u1_u14_u5_n148 ) , .A2( u1_u14_u5_n182 ) );
  OAI21_X1 u1_u14_u5_U51 (.ZN( u1_u14_u5_n124 ) , .A( u1_u14_u5_n177 ) , .B2( u1_u14_u5_n183 ) , .B1( u1_u14_u5_n189 ) );
  OAI21_X1 u1_u14_u5_U52 (.ZN( u1_u14_u5_n125 ) , .A( u1_u14_u5_n174 ) , .B2( u1_u14_u5_n185 ) , .B1( u1_u14_u5_n190 ) );
  AOI21_X1 u1_u14_u5_U53 (.A( u1_u14_u5_n153 ) , .B2( u1_u14_u5_n154 ) , .B1( u1_u14_u5_n155 ) , .ZN( u1_u14_u5_n164 ) );
  AOI21_X1 u1_u14_u5_U54 (.ZN( u1_u14_u5_n110 ) , .B1( u1_u14_u5_n122 ) , .B2( u1_u14_u5_n139 ) , .A( u1_u14_u5_n153 ) );
  INV_X1 u1_u14_u5_U55 (.A( u1_u14_u5_n153 ) , .ZN( u1_u14_u5_n176 ) );
  INV_X1 u1_u14_u5_U56 (.A( u1_u14_u5_n126 ) , .ZN( u1_u14_u5_n173 ) );
  AND2_X1 u1_u14_u5_U57 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n147 ) );
  AND2_X1 u1_u14_u5_U58 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n148 ) );
  NAND2_X1 u1_u14_u5_U59 (.A1( u1_u14_u5_n105 ) , .A2( u1_u14_u5_n106 ) , .ZN( u1_u14_u5_n158 ) );
  INV_X1 u1_u14_u5_U6 (.A( u1_u14_u5_n135 ) , .ZN( u1_u14_u5_n178 ) );
  NAND2_X1 u1_u14_u5_U60 (.A2( u1_u14_u5_n108 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n139 ) );
  NAND2_X1 u1_u14_u5_U61 (.A1( u1_u14_u5_n106 ) , .A2( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n119 ) );
  NAND2_X1 u1_u14_u5_U62 (.A2( u1_u14_u5_n103 ) , .A1( u1_u14_u5_n105 ) , .ZN( u1_u14_u5_n140 ) );
  NAND2_X1 u1_u14_u5_U63 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n105 ) , .ZN( u1_u14_u5_n155 ) );
  NAND2_X1 u1_u14_u5_U64 (.A2( u1_u14_u5_n106 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n122 ) );
  NAND2_X1 u1_u14_u5_U65 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n106 ) , .ZN( u1_u14_u5_n115 ) );
  NAND2_X1 u1_u14_u5_U66 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n103 ) , .ZN( u1_u14_u5_n161 ) );
  NAND2_X1 u1_u14_u5_U67 (.A1( u1_u14_u5_n105 ) , .A2( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n154 ) );
  INV_X1 u1_u14_u5_U68 (.A( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n172 ) );
  NAND2_X1 u1_u14_u5_U69 (.A1( u1_u14_u5_n103 ) , .A2( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n123 ) );
  OAI22_X1 u1_u14_u5_U7 (.B2( u1_u14_u5_n149 ) , .B1( u1_u14_u5_n150 ) , .A2( u1_u14_u5_n151 ) , .A1( u1_u14_u5_n152 ) , .ZN( u1_u14_u5_n165 ) );
  NAND2_X1 u1_u14_u5_U70 (.A2( u1_u14_u5_n103 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n151 ) );
  NAND2_X1 u1_u14_u5_U71 (.A2( u1_u14_u5_n107 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n120 ) );
  NAND2_X1 u1_u14_u5_U72 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n157 ) );
  AND2_X1 u1_u14_u5_U73 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n104 ) , .ZN( u1_u14_u5_n131 ) );
  INV_X1 u1_u14_u5_U74 (.A( u1_u14_u5_n102 ) , .ZN( u1_u14_u5_n195 ) );
  OAI221_X1 u1_u14_u5_U75 (.A( u1_u14_u5_n101 ) , .ZN( u1_u14_u5_n102 ) , .C2( u1_u14_u5_n115 ) , .C1( u1_u14_u5_n126 ) , .B1( u1_u14_u5_n134 ) , .B2( u1_u14_u5_n160 ) );
  OAI21_X1 u1_u14_u5_U76 (.ZN( u1_u14_u5_n101 ) , .B1( u1_u14_u5_n137 ) , .A( u1_u14_u5_n146 ) , .B2( u1_u14_u5_n147 ) );
  NOR2_X1 u1_u14_u5_U77 (.A2( u1_u14_X_34 ) , .A1( u1_u14_X_35 ) , .ZN( u1_u14_u5_n145 ) );
  NOR2_X1 u1_u14_u5_U78 (.A2( u1_u14_X_34 ) , .ZN( u1_u14_u5_n146 ) , .A1( u1_u14_u5_n171 ) );
  NOR2_X1 u1_u14_u5_U79 (.A2( u1_u14_X_31 ) , .A1( u1_u14_X_32 ) , .ZN( u1_u14_u5_n103 ) );
  NOR3_X1 u1_u14_u5_U8 (.A2( u1_u14_u5_n147 ) , .A1( u1_u14_u5_n148 ) , .ZN( u1_u14_u5_n149 ) , .A3( u1_u14_u5_n194 ) );
  NOR2_X1 u1_u14_u5_U80 (.A2( u1_u14_X_36 ) , .ZN( u1_u14_u5_n105 ) , .A1( u1_u14_u5_n180 ) );
  NOR2_X1 u1_u14_u5_U81 (.A2( u1_u14_X_33 ) , .ZN( u1_u14_u5_n108 ) , .A1( u1_u14_u5_n170 ) );
  NOR2_X1 u1_u14_u5_U82 (.A2( u1_u14_X_33 ) , .A1( u1_u14_X_36 ) , .ZN( u1_u14_u5_n107 ) );
  NOR2_X1 u1_u14_u5_U83 (.A2( u1_u14_X_31 ) , .ZN( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n181 ) );
  NAND2_X1 u1_u14_u5_U84 (.A2( u1_u14_X_34 ) , .A1( u1_u14_X_35 ) , .ZN( u1_u14_u5_n153 ) );
  NAND2_X1 u1_u14_u5_U85 (.A1( u1_u14_X_34 ) , .ZN( u1_u14_u5_n126 ) , .A2( u1_u14_u5_n171 ) );
  AND2_X1 u1_u14_u5_U86 (.A1( u1_u14_X_31 ) , .A2( u1_u14_X_32 ) , .ZN( u1_u14_u5_n106 ) );
  AND2_X1 u1_u14_u5_U87 (.A1( u1_u14_X_31 ) , .ZN( u1_u14_u5_n109 ) , .A2( u1_u14_u5_n181 ) );
  INV_X1 u1_u14_u5_U88 (.A( u1_u14_X_33 ) , .ZN( u1_u14_u5_n180 ) );
  INV_X1 u1_u14_u5_U89 (.A( u1_u14_X_35 ) , .ZN( u1_u14_u5_n171 ) );
  NOR2_X1 u1_u14_u5_U9 (.ZN( u1_u14_u5_n135 ) , .A1( u1_u14_u5_n173 ) , .A2( u1_u14_u5_n176 ) );
  INV_X1 u1_u14_u5_U90 (.A( u1_u14_X_36 ) , .ZN( u1_u14_u5_n170 ) );
  INV_X1 u1_u14_u5_U91 (.A( u1_u14_X_32 ) , .ZN( u1_u14_u5_n181 ) );
  NAND4_X1 u1_u14_u5_U92 (.ZN( u1_out14_29 ) , .A4( u1_u14_u5_n129 ) , .A3( u1_u14_u5_n130 ) , .A2( u1_u14_u5_n168 ) , .A1( u1_u14_u5_n196 ) );
  AOI221_X1 u1_u14_u5_U93 (.A( u1_u14_u5_n128 ) , .ZN( u1_u14_u5_n129 ) , .C2( u1_u14_u5_n132 ) , .B2( u1_u14_u5_n159 ) , .B1( u1_u14_u5_n176 ) , .C1( u1_u14_u5_n184 ) );
  AOI222_X1 u1_u14_u5_U94 (.ZN( u1_u14_u5_n130 ) , .A2( u1_u14_u5_n146 ) , .B1( u1_u14_u5_n147 ) , .C2( u1_u14_u5_n175 ) , .B2( u1_u14_u5_n179 ) , .A1( u1_u14_u5_n188 ) , .C1( u1_u14_u5_n194 ) );
  NAND4_X1 u1_u14_u5_U95 (.ZN( u1_out14_19 ) , .A4( u1_u14_u5_n166 ) , .A3( u1_u14_u5_n167 ) , .A2( u1_u14_u5_n168 ) , .A1( u1_u14_u5_n169 ) );
  AOI22_X1 u1_u14_u5_U96 (.B2( u1_u14_u5_n145 ) , .A2( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n167 ) , .B1( u1_u14_u5_n182 ) , .A1( u1_u14_u5_n189 ) );
  NOR4_X1 u1_u14_u5_U97 (.A4( u1_u14_u5_n162 ) , .A3( u1_u14_u5_n163 ) , .A2( u1_u14_u5_n164 ) , .A1( u1_u14_u5_n165 ) , .ZN( u1_u14_u5_n166 ) );
  NAND4_X1 u1_u14_u5_U98 (.ZN( u1_out14_11 ) , .A4( u1_u14_u5_n143 ) , .A3( u1_u14_u5_n144 ) , .A2( u1_u14_u5_n169 ) , .A1( u1_u14_u5_n196 ) );
  AOI22_X1 u1_u14_u5_U99 (.A2( u1_u14_u5_n132 ) , .ZN( u1_u14_u5_n144 ) , .B2( u1_u14_u5_n145 ) , .B1( u1_u14_u5_n184 ) , .A1( u1_u14_u5_n194 ) );
  AOI22_X1 u1_u14_u6_U10 (.A2( u1_u14_u6_n151 ) , .B2( u1_u14_u6_n161 ) , .A1( u1_u14_u6_n167 ) , .B1( u1_u14_u6_n170 ) , .ZN( u1_u14_u6_n89 ) );
  AOI21_X1 u1_u14_u6_U11 (.B1( u1_u14_u6_n107 ) , .B2( u1_u14_u6_n132 ) , .A( u1_u14_u6_n158 ) , .ZN( u1_u14_u6_n88 ) );
  AOI21_X1 u1_u14_u6_U12 (.B2( u1_u14_u6_n147 ) , .B1( u1_u14_u6_n148 ) , .ZN( u1_u14_u6_n149 ) , .A( u1_u14_u6_n158 ) );
  AOI21_X1 u1_u14_u6_U13 (.ZN( u1_u14_u6_n106 ) , .A( u1_u14_u6_n142 ) , .B2( u1_u14_u6_n159 ) , .B1( u1_u14_u6_n164 ) );
  INV_X1 u1_u14_u6_U14 (.A( u1_u14_u6_n155 ) , .ZN( u1_u14_u6_n161 ) );
  INV_X1 u1_u14_u6_U15 (.A( u1_u14_u6_n128 ) , .ZN( u1_u14_u6_n164 ) );
  NAND2_X1 u1_u14_u6_U16 (.ZN( u1_u14_u6_n110 ) , .A1( u1_u14_u6_n122 ) , .A2( u1_u14_u6_n129 ) );
  NAND2_X1 u1_u14_u6_U17 (.ZN( u1_u14_u6_n124 ) , .A2( u1_u14_u6_n146 ) , .A1( u1_u14_u6_n148 ) );
  INV_X1 u1_u14_u6_U18 (.A( u1_u14_u6_n132 ) , .ZN( u1_u14_u6_n171 ) );
  AND2_X1 u1_u14_u6_U19 (.A1( u1_u14_u6_n100 ) , .ZN( u1_u14_u6_n130 ) , .A2( u1_u14_u6_n147 ) );
  INV_X1 u1_u14_u6_U20 (.A( u1_u14_u6_n127 ) , .ZN( u1_u14_u6_n173 ) );
  INV_X1 u1_u14_u6_U21 (.A( u1_u14_u6_n121 ) , .ZN( u1_u14_u6_n167 ) );
  INV_X1 u1_u14_u6_U22 (.A( u1_u14_u6_n100 ) , .ZN( u1_u14_u6_n169 ) );
  INV_X1 u1_u14_u6_U23 (.A( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n170 ) );
  INV_X1 u1_u14_u6_U24 (.A( u1_u14_u6_n113 ) , .ZN( u1_u14_u6_n168 ) );
  AND2_X1 u1_u14_u6_U25 (.A1( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n119 ) , .ZN( u1_u14_u6_n133 ) );
  AND2_X1 u1_u14_u6_U26 (.A2( u1_u14_u6_n121 ) , .A1( u1_u14_u6_n122 ) , .ZN( u1_u14_u6_n131 ) );
  AND3_X1 u1_u14_u6_U27 (.ZN( u1_u14_u6_n120 ) , .A2( u1_u14_u6_n127 ) , .A1( u1_u14_u6_n132 ) , .A3( u1_u14_u6_n145 ) );
  INV_X1 u1_u14_u6_U28 (.A( u1_u14_u6_n146 ) , .ZN( u1_u14_u6_n163 ) );
  AOI222_X1 u1_u14_u6_U29 (.ZN( u1_u14_u6_n114 ) , .A1( u1_u14_u6_n118 ) , .A2( u1_u14_u6_n126 ) , .B2( u1_u14_u6_n151 ) , .C2( u1_u14_u6_n159 ) , .C1( u1_u14_u6_n168 ) , .B1( u1_u14_u6_n169 ) );
  INV_X1 u1_u14_u6_U3 (.A( u1_u14_u6_n110 ) , .ZN( u1_u14_u6_n166 ) );
  NOR2_X1 u1_u14_u6_U30 (.A1( u1_u14_u6_n162 ) , .A2( u1_u14_u6_n165 ) , .ZN( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U31 (.A1( u1_u14_u6_n144 ) , .ZN( u1_u14_u6_n151 ) , .A2( u1_u14_u6_n158 ) );
  NAND2_X1 u1_u14_u6_U32 (.ZN( u1_u14_u6_n132 ) , .A1( u1_u14_u6_n91 ) , .A2( u1_u14_u6_n97 ) );
  AOI22_X1 u1_u14_u6_U33 (.B2( u1_u14_u6_n110 ) , .B1( u1_u14_u6_n111 ) , .A1( u1_u14_u6_n112 ) , .ZN( u1_u14_u6_n115 ) , .A2( u1_u14_u6_n161 ) );
  NAND4_X1 u1_u14_u6_U34 (.A3( u1_u14_u6_n109 ) , .ZN( u1_u14_u6_n112 ) , .A4( u1_u14_u6_n132 ) , .A2( u1_u14_u6_n147 ) , .A1( u1_u14_u6_n166 ) );
  NOR2_X1 u1_u14_u6_U35 (.ZN( u1_u14_u6_n109 ) , .A1( u1_u14_u6_n170 ) , .A2( u1_u14_u6_n173 ) );
  NOR2_X1 u1_u14_u6_U36 (.A2( u1_u14_u6_n126 ) , .ZN( u1_u14_u6_n155 ) , .A1( u1_u14_u6_n160 ) );
  NAND2_X1 u1_u14_u6_U37 (.ZN( u1_u14_u6_n146 ) , .A2( u1_u14_u6_n94 ) , .A1( u1_u14_u6_n99 ) );
  AOI21_X1 u1_u14_u6_U38 (.A( u1_u14_u6_n144 ) , .B2( u1_u14_u6_n145 ) , .B1( u1_u14_u6_n146 ) , .ZN( u1_u14_u6_n150 ) );
  AOI211_X1 u1_u14_u6_U39 (.B( u1_u14_u6_n134 ) , .A( u1_u14_u6_n135 ) , .C1( u1_u14_u6_n136 ) , .ZN( u1_u14_u6_n137 ) , .C2( u1_u14_u6_n151 ) );
  INV_X1 u1_u14_u6_U4 (.A( u1_u14_u6_n142 ) , .ZN( u1_u14_u6_n174 ) );
  AOI21_X1 u1_u14_u6_U40 (.B2( u1_u14_u6_n132 ) , .B1( u1_u14_u6_n133 ) , .ZN( u1_u14_u6_n134 ) , .A( u1_u14_u6_n158 ) );
  NAND4_X1 u1_u14_u6_U41 (.A4( u1_u14_u6_n127 ) , .A3( u1_u14_u6_n128 ) , .A2( u1_u14_u6_n129 ) , .A1( u1_u14_u6_n130 ) , .ZN( u1_u14_u6_n136 ) );
  AOI21_X1 u1_u14_u6_U42 (.B1( u1_u14_u6_n131 ) , .ZN( u1_u14_u6_n135 ) , .A( u1_u14_u6_n144 ) , .B2( u1_u14_u6_n146 ) );
  INV_X1 u1_u14_u6_U43 (.A( u1_u14_u6_n111 ) , .ZN( u1_u14_u6_n158 ) );
  NAND2_X1 u1_u14_u6_U44 (.ZN( u1_u14_u6_n127 ) , .A1( u1_u14_u6_n91 ) , .A2( u1_u14_u6_n92 ) );
  NAND2_X1 u1_u14_u6_U45 (.ZN( u1_u14_u6_n129 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n96 ) );
  INV_X1 u1_u14_u6_U46 (.A( u1_u14_u6_n144 ) , .ZN( u1_u14_u6_n159 ) );
  NAND2_X1 u1_u14_u6_U47 (.ZN( u1_u14_u6_n145 ) , .A2( u1_u14_u6_n97 ) , .A1( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U48 (.ZN( u1_u14_u6_n148 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n94 ) );
  NAND2_X1 u1_u14_u6_U49 (.ZN( u1_u14_u6_n108 ) , .A2( u1_u14_u6_n139 ) , .A1( u1_u14_u6_n144 ) );
  NAND2_X1 u1_u14_u6_U5 (.A2( u1_u14_u6_n143 ) , .ZN( u1_u14_u6_n152 ) , .A1( u1_u14_u6_n166 ) );
  NAND2_X1 u1_u14_u6_U50 (.ZN( u1_u14_u6_n121 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n97 ) );
  NAND2_X1 u1_u14_u6_U51 (.ZN( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n95 ) );
  AND2_X1 u1_u14_u6_U52 (.ZN( u1_u14_u6_n118 ) , .A2( u1_u14_u6_n91 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U53 (.ZN( u1_u14_u6_n147 ) , .A2( u1_u14_u6_n98 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U54 (.ZN( u1_u14_u6_n128 ) , .A1( u1_u14_u6_n94 ) , .A2( u1_u14_u6_n96 ) );
  NAND2_X1 u1_u14_u6_U55 (.ZN( u1_u14_u6_n119 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U56 (.ZN( u1_u14_u6_n123 ) , .A2( u1_u14_u6_n91 ) , .A1( u1_u14_u6_n96 ) );
  NAND2_X1 u1_u14_u6_U57 (.ZN( u1_u14_u6_n100 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U58 (.ZN( u1_u14_u6_n122 ) , .A1( u1_u14_u6_n94 ) , .A2( u1_u14_u6_n97 ) );
  INV_X1 u1_u14_u6_U59 (.A( u1_u14_u6_n139 ) , .ZN( u1_u14_u6_n160 ) );
  AOI22_X1 u1_u14_u6_U6 (.B2( u1_u14_u6_n101 ) , .A1( u1_u14_u6_n102 ) , .ZN( u1_u14_u6_n103 ) , .B1( u1_u14_u6_n160 ) , .A2( u1_u14_u6_n161 ) );
  NAND2_X1 u1_u14_u6_U60 (.ZN( u1_u14_u6_n113 ) , .A1( u1_u14_u6_n96 ) , .A2( u1_u14_u6_n98 ) );
  NOR2_X1 u1_u14_u6_U61 (.A2( u1_u14_X_40 ) , .A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n126 ) );
  NOR2_X1 u1_u14_u6_U62 (.A2( u1_u14_X_39 ) , .A1( u1_u14_X_42 ) , .ZN( u1_u14_u6_n92 ) );
  NOR2_X1 u1_u14_u6_U63 (.A2( u1_u14_X_39 ) , .A1( u1_u14_u6_n156 ) , .ZN( u1_u14_u6_n97 ) );
  NOR2_X1 u1_u14_u6_U64 (.A2( u1_u14_X_38 ) , .A1( u1_u14_u6_n165 ) , .ZN( u1_u14_u6_n95 ) );
  NOR2_X1 u1_u14_u6_U65 (.A2( u1_u14_X_41 ) , .ZN( u1_u14_u6_n111 ) , .A1( u1_u14_u6_n157 ) );
  NOR2_X1 u1_u14_u6_U66 (.A2( u1_u14_X_37 ) , .A1( u1_u14_u6_n162 ) , .ZN( u1_u14_u6_n94 ) );
  NOR2_X1 u1_u14_u6_U67 (.A2( u1_u14_X_37 ) , .A1( u1_u14_X_38 ) , .ZN( u1_u14_u6_n91 ) );
  NAND2_X1 u1_u14_u6_U68 (.A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n144 ) , .A2( u1_u14_u6_n157 ) );
  NAND2_X1 u1_u14_u6_U69 (.A2( u1_u14_X_40 ) , .A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n139 ) );
  NOR2_X1 u1_u14_u6_U7 (.A1( u1_u14_u6_n118 ) , .ZN( u1_u14_u6_n143 ) , .A2( u1_u14_u6_n168 ) );
  AND2_X1 u1_u14_u6_U70 (.A1( u1_u14_X_39 ) , .A2( u1_u14_u6_n156 ) , .ZN( u1_u14_u6_n96 ) );
  AND2_X1 u1_u14_u6_U71 (.A1( u1_u14_X_39 ) , .A2( u1_u14_X_42 ) , .ZN( u1_u14_u6_n99 ) );
  INV_X1 u1_u14_u6_U72 (.A( u1_u14_X_40 ) , .ZN( u1_u14_u6_n157 ) );
  INV_X1 u1_u14_u6_U73 (.A( u1_u14_X_37 ) , .ZN( u1_u14_u6_n165 ) );
  INV_X1 u1_u14_u6_U74 (.A( u1_u14_X_38 ) , .ZN( u1_u14_u6_n162 ) );
  INV_X1 u1_u14_u6_U75 (.A( u1_u14_X_42 ) , .ZN( u1_u14_u6_n156 ) );
  NAND4_X1 u1_u14_u6_U76 (.ZN( u1_out14_32 ) , .A4( u1_u14_u6_n103 ) , .A3( u1_u14_u6_n104 ) , .A2( u1_u14_u6_n105 ) , .A1( u1_u14_u6_n106 ) );
  AOI22_X1 u1_u14_u6_U77 (.ZN( u1_u14_u6_n105 ) , .A2( u1_u14_u6_n108 ) , .A1( u1_u14_u6_n118 ) , .B2( u1_u14_u6_n126 ) , .B1( u1_u14_u6_n171 ) );
  AOI22_X1 u1_u14_u6_U78 (.ZN( u1_u14_u6_n104 ) , .A1( u1_u14_u6_n111 ) , .B1( u1_u14_u6_n124 ) , .B2( u1_u14_u6_n151 ) , .A2( u1_u14_u6_n93 ) );
  NAND4_X1 u1_u14_u6_U79 (.ZN( u1_out14_12 ) , .A4( u1_u14_u6_n114 ) , .A3( u1_u14_u6_n115 ) , .A2( u1_u14_u6_n116 ) , .A1( u1_u14_u6_n117 ) );
  INV_X1 u1_u14_u6_U8 (.ZN( u1_u14_u6_n172 ) , .A( u1_u14_u6_n88 ) );
  OAI22_X1 u1_u14_u6_U80 (.B2( u1_u14_u6_n111 ) , .ZN( u1_u14_u6_n116 ) , .B1( u1_u14_u6_n126 ) , .A2( u1_u14_u6_n164 ) , .A1( u1_u14_u6_n167 ) );
  OAI21_X1 u1_u14_u6_U81 (.A( u1_u14_u6_n108 ) , .ZN( u1_u14_u6_n117 ) , .B2( u1_u14_u6_n141 ) , .B1( u1_u14_u6_n163 ) );
  OAI211_X1 u1_u14_u6_U82 (.ZN( u1_out14_22 ) , .B( u1_u14_u6_n137 ) , .A( u1_u14_u6_n138 ) , .C2( u1_u14_u6_n139 ) , .C1( u1_u14_u6_n140 ) );
  AOI22_X1 u1_u14_u6_U83 (.B1( u1_u14_u6_n124 ) , .A2( u1_u14_u6_n125 ) , .A1( u1_u14_u6_n126 ) , .ZN( u1_u14_u6_n138 ) , .B2( u1_u14_u6_n161 ) );
  AND4_X1 u1_u14_u6_U84 (.A3( u1_u14_u6_n119 ) , .A1( u1_u14_u6_n120 ) , .A4( u1_u14_u6_n129 ) , .ZN( u1_u14_u6_n140 ) , .A2( u1_u14_u6_n143 ) );
  OAI211_X1 u1_u14_u6_U85 (.ZN( u1_out14_7 ) , .B( u1_u14_u6_n153 ) , .C2( u1_u14_u6_n154 ) , .C1( u1_u14_u6_n155 ) , .A( u1_u14_u6_n174 ) );
  NOR3_X1 u1_u14_u6_U86 (.A1( u1_u14_u6_n141 ) , .ZN( u1_u14_u6_n154 ) , .A3( u1_u14_u6_n164 ) , .A2( u1_u14_u6_n171 ) );
  AOI211_X1 u1_u14_u6_U87 (.B( u1_u14_u6_n149 ) , .A( u1_u14_u6_n150 ) , .C2( u1_u14_u6_n151 ) , .C1( u1_u14_u6_n152 ) , .ZN( u1_u14_u6_n153 ) );
  NAND3_X1 u1_u14_u6_U88 (.A2( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n125 ) , .A1( u1_u14_u6_n130 ) , .A3( u1_u14_u6_n131 ) );
  NAND3_X1 u1_u14_u6_U89 (.A3( u1_u14_u6_n133 ) , .ZN( u1_u14_u6_n141 ) , .A1( u1_u14_u6_n145 ) , .A2( u1_u14_u6_n148 ) );
  OAI21_X1 u1_u14_u6_U9 (.A( u1_u14_u6_n159 ) , .B1( u1_u14_u6_n169 ) , .B2( u1_u14_u6_n173 ) , .ZN( u1_u14_u6_n90 ) );
  NAND3_X1 u1_u14_u6_U90 (.ZN( u1_u14_u6_n101 ) , .A3( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n121 ) , .A1( u1_u14_u6_n127 ) );
  NAND3_X1 u1_u14_u6_U91 (.ZN( u1_u14_u6_n102 ) , .A3( u1_u14_u6_n130 ) , .A2( u1_u14_u6_n145 ) , .A1( u1_u14_u6_n166 ) );
  NAND3_X1 u1_u14_u6_U92 (.A3( u1_u14_u6_n113 ) , .A1( u1_u14_u6_n119 ) , .A2( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n93 ) );
  NAND3_X1 u1_u14_u6_U93 (.ZN( u1_u14_u6_n142 ) , .A2( u1_u14_u6_n172 ) , .A3( u1_u14_u6_n89 ) , .A1( u1_u14_u6_n90 ) );
  OAI21_X1 u1_u14_u7_U10 (.A( u1_u14_u7_n161 ) , .B1( u1_u14_u7_n168 ) , .B2( u1_u14_u7_n173 ) , .ZN( u1_u14_u7_n91 ) );
  AOI211_X1 u1_u14_u7_U11 (.A( u1_u14_u7_n117 ) , .ZN( u1_u14_u7_n118 ) , .C2( u1_u14_u7_n126 ) , .C1( u1_u14_u7_n177 ) , .B( u1_u14_u7_n180 ) );
  OAI22_X1 u1_u14_u7_U12 (.B1( u1_u14_u7_n115 ) , .ZN( u1_u14_u7_n117 ) , .A2( u1_u14_u7_n133 ) , .A1( u1_u14_u7_n137 ) , .B2( u1_u14_u7_n162 ) );
  INV_X1 u1_u14_u7_U13 (.A( u1_u14_u7_n116 ) , .ZN( u1_u14_u7_n180 ) );
  NOR3_X1 u1_u14_u7_U14 (.ZN( u1_u14_u7_n115 ) , .A3( u1_u14_u7_n145 ) , .A2( u1_u14_u7_n168 ) , .A1( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U15 (.A( u1_u14_u7_n133 ) , .ZN( u1_u14_u7_n176 ) );
  NOR3_X1 u1_u14_u7_U16 (.A2( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n135 ) , .ZN( u1_u14_u7_n136 ) , .A3( u1_u14_u7_n171 ) );
  NOR2_X1 u1_u14_u7_U17 (.A1( u1_u14_u7_n130 ) , .A2( u1_u14_u7_n134 ) , .ZN( u1_u14_u7_n153 ) );
  AOI21_X1 u1_u14_u7_U18 (.ZN( u1_u14_u7_n104 ) , .B2( u1_u14_u7_n112 ) , .B1( u1_u14_u7_n127 ) , .A( u1_u14_u7_n164 ) );
  AOI21_X1 u1_u14_u7_U19 (.ZN( u1_u14_u7_n106 ) , .B1( u1_u14_u7_n133 ) , .B2( u1_u14_u7_n146 ) , .A( u1_u14_u7_n162 ) );
  AOI21_X1 u1_u14_u7_U20 (.A( u1_u14_u7_n101 ) , .ZN( u1_u14_u7_n107 ) , .B2( u1_u14_u7_n128 ) , .B1( u1_u14_u7_n175 ) );
  INV_X1 u1_u14_u7_U21 (.A( u1_u14_u7_n101 ) , .ZN( u1_u14_u7_n165 ) );
  NOR2_X1 u1_u14_u7_U22 (.ZN( u1_u14_u7_n111 ) , .A2( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U23 (.A( u1_u14_u7_n138 ) , .ZN( u1_u14_u7_n171 ) );
  INV_X1 u1_u14_u7_U24 (.A( u1_u14_u7_n131 ) , .ZN( u1_u14_u7_n177 ) );
  INV_X1 u1_u14_u7_U25 (.A( u1_u14_u7_n110 ) , .ZN( u1_u14_u7_n174 ) );
  NAND2_X1 u1_u14_u7_U26 (.A1( u1_u14_u7_n129 ) , .A2( u1_u14_u7_n132 ) , .ZN( u1_u14_u7_n149 ) );
  NAND2_X1 u1_u14_u7_U27 (.A1( u1_u14_u7_n113 ) , .A2( u1_u14_u7_n124 ) , .ZN( u1_u14_u7_n130 ) );
  INV_X1 u1_u14_u7_U28 (.A( u1_u14_u7_n112 ) , .ZN( u1_u14_u7_n173 ) );
  INV_X1 u1_u14_u7_U29 (.A( u1_u14_u7_n128 ) , .ZN( u1_u14_u7_n168 ) );
  OAI21_X1 u1_u14_u7_U3 (.ZN( u1_u14_u7_n159 ) , .A( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n171 ) , .B1( u1_u14_u7_n174 ) );
  INV_X1 u1_u14_u7_U30 (.A( u1_u14_u7_n148 ) , .ZN( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U31 (.A( u1_u14_u7_n127 ) , .ZN( u1_u14_u7_n179 ) );
  NOR2_X1 u1_u14_u7_U32 (.ZN( u1_u14_u7_n101 ) , .A2( u1_u14_u7_n150 ) , .A1( u1_u14_u7_n156 ) );
  AOI211_X1 u1_u14_u7_U33 (.B( u1_u14_u7_n139 ) , .A( u1_u14_u7_n140 ) , .C2( u1_u14_u7_n141 ) , .ZN( u1_u14_u7_n142 ) , .C1( u1_u14_u7_n156 ) );
  NAND4_X1 u1_u14_u7_U34 (.A3( u1_u14_u7_n127 ) , .A2( u1_u14_u7_n128 ) , .A1( u1_u14_u7_n129 ) , .ZN( u1_u14_u7_n141 ) , .A4( u1_u14_u7_n147 ) );
  AOI21_X1 u1_u14_u7_U35 (.A( u1_u14_u7_n137 ) , .B1( u1_u14_u7_n138 ) , .ZN( u1_u14_u7_n139 ) , .B2( u1_u14_u7_n146 ) );
  OAI22_X1 u1_u14_u7_U36 (.B1( u1_u14_u7_n136 ) , .ZN( u1_u14_u7_n140 ) , .A1( u1_u14_u7_n153 ) , .B2( u1_u14_u7_n162 ) , .A2( u1_u14_u7_n164 ) );
  INV_X1 u1_u14_u7_U37 (.A( u1_u14_u7_n125 ) , .ZN( u1_u14_u7_n161 ) );
  AOI21_X1 u1_u14_u7_U38 (.ZN( u1_u14_u7_n123 ) , .B1( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n177 ) , .A( u1_u14_u7_n97 ) );
  AOI21_X1 u1_u14_u7_U39 (.B2( u1_u14_u7_n113 ) , .B1( u1_u14_u7_n124 ) , .A( u1_u14_u7_n125 ) , .ZN( u1_u14_u7_n97 ) );
  INV_X1 u1_u14_u7_U4 (.A( u1_u14_u7_n149 ) , .ZN( u1_u14_u7_n175 ) );
  INV_X1 u1_u14_u7_U40 (.A( u1_u14_u7_n152 ) , .ZN( u1_u14_u7_n162 ) );
  AOI22_X1 u1_u14_u7_U41 (.A2( u1_u14_u7_n114 ) , .ZN( u1_u14_u7_n119 ) , .B1( u1_u14_u7_n130 ) , .A1( u1_u14_u7_n156 ) , .B2( u1_u14_u7_n165 ) );
  NAND2_X1 u1_u14_u7_U42 (.A2( u1_u14_u7_n112 ) , .ZN( u1_u14_u7_n114 ) , .A1( u1_u14_u7_n175 ) );
  NOR2_X1 u1_u14_u7_U43 (.ZN( u1_u14_u7_n137 ) , .A1( u1_u14_u7_n150 ) , .A2( u1_u14_u7_n161 ) );
  AND2_X1 u1_u14_u7_U44 (.ZN( u1_u14_u7_n145 ) , .A2( u1_u14_u7_n98 ) , .A1( u1_u14_u7_n99 ) );
  AOI21_X1 u1_u14_u7_U45 (.ZN( u1_u14_u7_n105 ) , .B2( u1_u14_u7_n110 ) , .A( u1_u14_u7_n125 ) , .B1( u1_u14_u7_n147 ) );
  NAND2_X1 u1_u14_u7_U46 (.ZN( u1_u14_u7_n146 ) , .A1( u1_u14_u7_n95 ) , .A2( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U47 (.A2( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n147 ) , .A1( u1_u14_u7_n93 ) );
  NAND2_X1 u1_u14_u7_U48 (.A1( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n127 ) , .A2( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U49 (.A2( u1_u14_u7_n102 ) , .A1( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n133 ) );
  INV_X1 u1_u14_u7_U5 (.A( u1_u14_u7_n154 ) , .ZN( u1_u14_u7_n178 ) );
  OR2_X1 u1_u14_u7_U50 (.ZN( u1_u14_u7_n126 ) , .A2( u1_u14_u7_n152 ) , .A1( u1_u14_u7_n156 ) );
  NAND2_X1 u1_u14_u7_U51 (.ZN( u1_u14_u7_n112 ) , .A2( u1_u14_u7_n96 ) , .A1( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U52 (.A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n128 ) , .A1( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U53 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n113 ) , .A2( u1_u14_u7_n93 ) );
  NAND2_X1 u1_u14_u7_U54 (.ZN( u1_u14_u7_n110 ) , .A1( u1_u14_u7_n95 ) , .A2( u1_u14_u7_n96 ) );
  INV_X1 u1_u14_u7_U55 (.A( u1_u14_u7_n150 ) , .ZN( u1_u14_u7_n164 ) );
  AND2_X1 u1_u14_u7_U56 (.ZN( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n93 ) , .A2( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U57 (.A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n124 ) , .A1( u1_u14_u7_n96 ) );
  NAND2_X1 u1_u14_u7_U58 (.A1( u1_u14_u7_n100 ) , .A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n129 ) );
  NAND2_X1 u1_u14_u7_U59 (.A2( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n131 ) , .A1( u1_u14_u7_n95 ) );
  AOI211_X1 u1_u14_u7_U6 (.ZN( u1_u14_u7_n116 ) , .A( u1_u14_u7_n155 ) , .C1( u1_u14_u7_n161 ) , .C2( u1_u14_u7_n171 ) , .B( u1_u14_u7_n94 ) );
  NAND2_X1 u1_u14_u7_U60 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n138 ) , .A2( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U61 (.ZN( u1_u14_u7_n132 ) , .A1( u1_u14_u7_n93 ) , .A2( u1_u14_u7_n96 ) );
  NAND2_X1 u1_u14_u7_U62 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n148 ) , .A2( u1_u14_u7_n95 ) );
  AOI211_X1 u1_u14_u7_U63 (.B( u1_u14_u7_n154 ) , .A( u1_u14_u7_n155 ) , .C1( u1_u14_u7_n156 ) , .ZN( u1_u14_u7_n157 ) , .C2( u1_u14_u7_n172 ) );
  INV_X1 u1_u14_u7_U64 (.A( u1_u14_u7_n153 ) , .ZN( u1_u14_u7_n172 ) );
  NOR2_X1 u1_u14_u7_U65 (.A2( u1_u14_X_47 ) , .ZN( u1_u14_u7_n150 ) , .A1( u1_u14_u7_n163 ) );
  NOR2_X1 u1_u14_u7_U66 (.A2( u1_u14_X_43 ) , .A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n103 ) );
  NOR2_X1 u1_u14_u7_U67 (.A2( u1_u14_X_48 ) , .A1( u1_u14_u7_n166 ) , .ZN( u1_u14_u7_n95 ) );
  NOR2_X1 u1_u14_u7_U68 (.A2( u1_u14_X_45 ) , .A1( u1_u14_X_48 ) , .ZN( u1_u14_u7_n99 ) );
  NOR2_X1 u1_u14_u7_U69 (.A2( u1_u14_X_44 ) , .A1( u1_u14_u7_n167 ) , .ZN( u1_u14_u7_n98 ) );
  OAI222_X1 u1_u14_u7_U7 (.C2( u1_u14_u7_n101 ) , .B2( u1_u14_u7_n111 ) , .A1( u1_u14_u7_n113 ) , .C1( u1_u14_u7_n146 ) , .A2( u1_u14_u7_n162 ) , .B1( u1_u14_u7_n164 ) , .ZN( u1_u14_u7_n94 ) );
  NOR2_X1 u1_u14_u7_U70 (.A2( u1_u14_X_46 ) , .A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n152 ) );
  NAND2_X1 u1_u14_u7_U71 (.A2( u1_u14_X_46 ) , .A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n125 ) );
  AND2_X1 u1_u14_u7_U72 (.A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n156 ) , .A2( u1_u14_u7_n163 ) );
  AND2_X1 u1_u14_u7_U73 (.A2( u1_u14_X_45 ) , .A1( u1_u14_X_48 ) , .ZN( u1_u14_u7_n102 ) );
  AND2_X1 u1_u14_u7_U74 (.A2( u1_u14_X_43 ) , .A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n96 ) );
  AND2_X1 u1_u14_u7_U75 (.A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n100 ) , .A2( u1_u14_u7_n167 ) );
  AND2_X1 u1_u14_u7_U76 (.A1( u1_u14_X_48 ) , .A2( u1_u14_u7_n166 ) , .ZN( u1_u14_u7_n93 ) );
  INV_X1 u1_u14_u7_U77 (.A( u1_u14_X_46 ) , .ZN( u1_u14_u7_n163 ) );
  INV_X1 u1_u14_u7_U78 (.A( u1_u14_X_43 ) , .ZN( u1_u14_u7_n167 ) );
  INV_X1 u1_u14_u7_U79 (.A( u1_u14_X_45 ) , .ZN( u1_u14_u7_n166 ) );
  OAI221_X1 u1_u14_u7_U8 (.C1( u1_u14_u7_n101 ) , .C2( u1_u14_u7_n147 ) , .ZN( u1_u14_u7_n155 ) , .B2( u1_u14_u7_n162 ) , .A( u1_u14_u7_n91 ) , .B1( u1_u14_u7_n92 ) );
  NAND4_X1 u1_u14_u7_U80 (.ZN( u1_out14_5 ) , .A4( u1_u14_u7_n108 ) , .A3( u1_u14_u7_n109 ) , .A1( u1_u14_u7_n116 ) , .A2( u1_u14_u7_n123 ) );
  AOI22_X1 u1_u14_u7_U81 (.ZN( u1_u14_u7_n109 ) , .A2( u1_u14_u7_n126 ) , .B2( u1_u14_u7_n145 ) , .B1( u1_u14_u7_n156 ) , .A1( u1_u14_u7_n171 ) );
  NOR4_X1 u1_u14_u7_U82 (.A4( u1_u14_u7_n104 ) , .A3( u1_u14_u7_n105 ) , .A2( u1_u14_u7_n106 ) , .A1( u1_u14_u7_n107 ) , .ZN( u1_u14_u7_n108 ) );
  NAND4_X1 u1_u14_u7_U83 (.ZN( u1_out14_27 ) , .A4( u1_u14_u7_n118 ) , .A3( u1_u14_u7_n119 ) , .A2( u1_u14_u7_n120 ) , .A1( u1_u14_u7_n121 ) );
  OAI21_X1 u1_u14_u7_U84 (.ZN( u1_u14_u7_n121 ) , .B2( u1_u14_u7_n145 ) , .A( u1_u14_u7_n150 ) , .B1( u1_u14_u7_n174 ) );
  OAI21_X1 u1_u14_u7_U85 (.ZN( u1_u14_u7_n120 ) , .A( u1_u14_u7_n161 ) , .B2( u1_u14_u7_n170 ) , .B1( u1_u14_u7_n179 ) );
  NAND4_X1 u1_u14_u7_U86 (.ZN( u1_out14_21 ) , .A4( u1_u14_u7_n157 ) , .A3( u1_u14_u7_n158 ) , .A2( u1_u14_u7_n159 ) , .A1( u1_u14_u7_n160 ) );
  OAI21_X1 u1_u14_u7_U87 (.B1( u1_u14_u7_n145 ) , .ZN( u1_u14_u7_n160 ) , .A( u1_u14_u7_n161 ) , .B2( u1_u14_u7_n177 ) );
  AOI22_X1 u1_u14_u7_U88 (.B2( u1_u14_u7_n149 ) , .B1( u1_u14_u7_n150 ) , .A2( u1_u14_u7_n151 ) , .A1( u1_u14_u7_n152 ) , .ZN( u1_u14_u7_n158 ) );
  NAND4_X1 u1_u14_u7_U89 (.ZN( u1_out14_15 ) , .A4( u1_u14_u7_n142 ) , .A3( u1_u14_u7_n143 ) , .A2( u1_u14_u7_n144 ) , .A1( u1_u14_u7_n178 ) );
  AND3_X1 u1_u14_u7_U9 (.A3( u1_u14_u7_n110 ) , .A2( u1_u14_u7_n127 ) , .A1( u1_u14_u7_n132 ) , .ZN( u1_u14_u7_n92 ) );
  OR2_X1 u1_u14_u7_U90 (.A2( u1_u14_u7_n125 ) , .A1( u1_u14_u7_n129 ) , .ZN( u1_u14_u7_n144 ) );
  AOI22_X1 u1_u14_u7_U91 (.A2( u1_u14_u7_n126 ) , .ZN( u1_u14_u7_n143 ) , .B2( u1_u14_u7_n165 ) , .B1( u1_u14_u7_n173 ) , .A1( u1_u14_u7_n174 ) );
  OAI211_X1 u1_u14_u7_U92 (.B( u1_u14_u7_n122 ) , .A( u1_u14_u7_n123 ) , .C2( u1_u14_u7_n124 ) , .ZN( u1_u14_u7_n154 ) , .C1( u1_u14_u7_n162 ) );
  AOI222_X1 u1_u14_u7_U93 (.ZN( u1_u14_u7_n122 ) , .C2( u1_u14_u7_n126 ) , .C1( u1_u14_u7_n145 ) , .B1( u1_u14_u7_n161 ) , .A2( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n170 ) , .A1( u1_u14_u7_n176 ) );
  INV_X1 u1_u14_u7_U94 (.A( u1_u14_u7_n111 ) , .ZN( u1_u14_u7_n170 ) );
  NAND3_X1 u1_u14_u7_U95 (.A3( u1_u14_u7_n146 ) , .A2( u1_u14_u7_n147 ) , .A1( u1_u14_u7_n148 ) , .ZN( u1_u14_u7_n151 ) );
  NAND3_X1 u1_u14_u7_U96 (.A3( u1_u14_u7_n131 ) , .A2( u1_u14_u7_n132 ) , .A1( u1_u14_u7_n133 ) , .ZN( u1_u14_u7_n135 ) );
  XOR2_X1 u1_u3_U1 (.B( u1_K4_9 ) , .A( u1_R2_6 ) , .Z( u1_u3_X_9 ) );
  XOR2_X1 u1_u3_U2 (.B( u1_K4_8 ) , .A( u1_R2_5 ) , .Z( u1_u3_X_8 ) );
  XOR2_X1 u1_u3_U3 (.B( u1_K4_7 ) , .A( u1_R2_4 ) , .Z( u1_u3_X_7 ) );
  XOR2_X1 u1_u3_U46 (.B( u1_K4_12 ) , .A( u1_R2_9 ) , .Z( u1_u3_X_12 ) );
  XOR2_X1 u1_u3_U47 (.B( u1_K4_11 ) , .A( u1_R2_8 ) , .Z( u1_u3_X_11 ) );
  XOR2_X1 u1_u3_U48 (.B( u1_K4_10 ) , .A( u1_R2_7 ) , .Z( u1_u3_X_10 ) );
  AOI21_X1 u1_u3_u1_U10 (.B2( u1_u3_u1_n155 ) , .B1( u1_u3_u1_n156 ) , .ZN( u1_u3_u1_n157 ) , .A( u1_u3_u1_n174 ) );
  NAND3_X1 u1_u3_u1_U100 (.ZN( u1_u3_u1_n113 ) , .A1( u1_u3_u1_n120 ) , .A3( u1_u3_u1_n133 ) , .A2( u1_u3_u1_n155 ) );
  NAND2_X1 u1_u3_u1_U11 (.ZN( u1_u3_u1_n140 ) , .A2( u1_u3_u1_n150 ) , .A1( u1_u3_u1_n155 ) );
  NAND2_X1 u1_u3_u1_U12 (.A1( u1_u3_u1_n131 ) , .ZN( u1_u3_u1_n147 ) , .A2( u1_u3_u1_n153 ) );
  INV_X1 u1_u3_u1_U13 (.A( u1_u3_u1_n139 ) , .ZN( u1_u3_u1_n174 ) );
  OR4_X1 u1_u3_u1_U14 (.A4( u1_u3_u1_n106 ) , .A3( u1_u3_u1_n107 ) , .ZN( u1_u3_u1_n108 ) , .A1( u1_u3_u1_n117 ) , .A2( u1_u3_u1_n184 ) );
  AOI21_X1 u1_u3_u1_U15 (.ZN( u1_u3_u1_n106 ) , .A( u1_u3_u1_n112 ) , .B1( u1_u3_u1_n154 ) , .B2( u1_u3_u1_n156 ) );
  INV_X1 u1_u3_u1_U16 (.A( u1_u3_u1_n101 ) , .ZN( u1_u3_u1_n184 ) );
  AOI21_X1 u1_u3_u1_U17 (.ZN( u1_u3_u1_n107 ) , .B1( u1_u3_u1_n134 ) , .B2( u1_u3_u1_n149 ) , .A( u1_u3_u1_n174 ) );
  INV_X1 u1_u3_u1_U18 (.A( u1_u3_u1_n112 ) , .ZN( u1_u3_u1_n171 ) );
  NAND2_X1 u1_u3_u1_U19 (.ZN( u1_u3_u1_n141 ) , .A1( u1_u3_u1_n153 ) , .A2( u1_u3_u1_n156 ) );
  AND2_X1 u1_u3_u1_U20 (.A1( u1_u3_u1_n123 ) , .ZN( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n161 ) );
  NAND2_X1 u1_u3_u1_U21 (.A2( u1_u3_u1_n115 ) , .A1( u1_u3_u1_n116 ) , .ZN( u1_u3_u1_n148 ) );
  NAND2_X1 u1_u3_u1_U22 (.A2( u1_u3_u1_n133 ) , .A1( u1_u3_u1_n135 ) , .ZN( u1_u3_u1_n159 ) );
  NAND2_X1 u1_u3_u1_U23 (.A2( u1_u3_u1_n115 ) , .A1( u1_u3_u1_n120 ) , .ZN( u1_u3_u1_n132 ) );
  INV_X1 u1_u3_u1_U24 (.A( u1_u3_u1_n154 ) , .ZN( u1_u3_u1_n178 ) );
  AOI22_X1 u1_u3_u1_U25 (.B2( u1_u3_u1_n113 ) , .A2( u1_u3_u1_n114 ) , .ZN( u1_u3_u1_n125 ) , .A1( u1_u3_u1_n171 ) , .B1( u1_u3_u1_n173 ) );
  NAND2_X1 u1_u3_u1_U26 (.ZN( u1_u3_u1_n114 ) , .A1( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n156 ) );
  INV_X1 u1_u3_u1_U27 (.A( u1_u3_u1_n151 ) , .ZN( u1_u3_u1_n183 ) );
  AND2_X1 u1_u3_u1_U28 (.A1( u1_u3_u1_n129 ) , .A2( u1_u3_u1_n133 ) , .ZN( u1_u3_u1_n149 ) );
  INV_X1 u1_u3_u1_U29 (.A( u1_u3_u1_n131 ) , .ZN( u1_u3_u1_n180 ) );
  INV_X1 u1_u3_u1_U3 (.A( u1_u3_u1_n159 ) , .ZN( u1_u3_u1_n182 ) );
  AOI221_X1 u1_u3_u1_U30 (.B1( u1_u3_u1_n140 ) , .ZN( u1_u3_u1_n167 ) , .B2( u1_u3_u1_n172 ) , .C2( u1_u3_u1_n175 ) , .C1( u1_u3_u1_n178 ) , .A( u1_u3_u1_n188 ) );
  INV_X1 u1_u3_u1_U31 (.ZN( u1_u3_u1_n188 ) , .A( u1_u3_u1_n97 ) );
  AOI211_X1 u1_u3_u1_U32 (.A( u1_u3_u1_n118 ) , .C1( u1_u3_u1_n132 ) , .C2( u1_u3_u1_n139 ) , .B( u1_u3_u1_n96 ) , .ZN( u1_u3_u1_n97 ) );
  AOI21_X1 u1_u3_u1_U33 (.B2( u1_u3_u1_n121 ) , .B1( u1_u3_u1_n135 ) , .A( u1_u3_u1_n152 ) , .ZN( u1_u3_u1_n96 ) );
  OAI221_X1 u1_u3_u1_U34 (.A( u1_u3_u1_n119 ) , .C2( u1_u3_u1_n129 ) , .ZN( u1_u3_u1_n138 ) , .B2( u1_u3_u1_n152 ) , .C1( u1_u3_u1_n174 ) , .B1( u1_u3_u1_n187 ) );
  INV_X1 u1_u3_u1_U35 (.A( u1_u3_u1_n148 ) , .ZN( u1_u3_u1_n187 ) );
  AOI211_X1 u1_u3_u1_U36 (.B( u1_u3_u1_n117 ) , .A( u1_u3_u1_n118 ) , .ZN( u1_u3_u1_n119 ) , .C2( u1_u3_u1_n146 ) , .C1( u1_u3_u1_n159 ) );
  NOR2_X1 u1_u3_u1_U37 (.A1( u1_u3_u1_n168 ) , .A2( u1_u3_u1_n176 ) , .ZN( u1_u3_u1_n98 ) );
  AOI211_X1 u1_u3_u1_U38 (.B( u1_u3_u1_n162 ) , .A( u1_u3_u1_n163 ) , .C2( u1_u3_u1_n164 ) , .ZN( u1_u3_u1_n165 ) , .C1( u1_u3_u1_n171 ) );
  AOI21_X1 u1_u3_u1_U39 (.A( u1_u3_u1_n160 ) , .B2( u1_u3_u1_n161 ) , .ZN( u1_u3_u1_n162 ) , .B1( u1_u3_u1_n182 ) );
  AOI221_X1 u1_u3_u1_U4 (.A( u1_u3_u1_n138 ) , .C2( u1_u3_u1_n139 ) , .C1( u1_u3_u1_n140 ) , .B2( u1_u3_u1_n141 ) , .ZN( u1_u3_u1_n142 ) , .B1( u1_u3_u1_n175 ) );
  OR2_X1 u1_u3_u1_U40 (.A2( u1_u3_u1_n157 ) , .A1( u1_u3_u1_n158 ) , .ZN( u1_u3_u1_n163 ) );
  NAND2_X1 u1_u3_u1_U41 (.A1( u1_u3_u1_n128 ) , .ZN( u1_u3_u1_n146 ) , .A2( u1_u3_u1_n160 ) );
  NAND2_X1 u1_u3_u1_U42 (.A2( u1_u3_u1_n112 ) , .ZN( u1_u3_u1_n139 ) , .A1( u1_u3_u1_n152 ) );
  NAND2_X1 u1_u3_u1_U43 (.A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n156 ) , .A2( u1_u3_u1_n99 ) );
  NOR2_X1 u1_u3_u1_U44 (.ZN( u1_u3_u1_n117 ) , .A1( u1_u3_u1_n121 ) , .A2( u1_u3_u1_n160 ) );
  OAI21_X1 u1_u3_u1_U45 (.B2( u1_u3_u1_n123 ) , .ZN( u1_u3_u1_n145 ) , .B1( u1_u3_u1_n160 ) , .A( u1_u3_u1_n185 ) );
  INV_X1 u1_u3_u1_U46 (.A( u1_u3_u1_n122 ) , .ZN( u1_u3_u1_n185 ) );
  AOI21_X1 u1_u3_u1_U47 (.B2( u1_u3_u1_n120 ) , .B1( u1_u3_u1_n121 ) , .ZN( u1_u3_u1_n122 ) , .A( u1_u3_u1_n128 ) );
  AOI21_X1 u1_u3_u1_U48 (.A( u1_u3_u1_n128 ) , .B2( u1_u3_u1_n129 ) , .ZN( u1_u3_u1_n130 ) , .B1( u1_u3_u1_n150 ) );
  NAND2_X1 u1_u3_u1_U49 (.ZN( u1_u3_u1_n112 ) , .A1( u1_u3_u1_n169 ) , .A2( u1_u3_u1_n170 ) );
  AOI211_X1 u1_u3_u1_U5 (.ZN( u1_u3_u1_n124 ) , .A( u1_u3_u1_n138 ) , .C2( u1_u3_u1_n139 ) , .B( u1_u3_u1_n145 ) , .C1( u1_u3_u1_n147 ) );
  NAND2_X1 u1_u3_u1_U50 (.ZN( u1_u3_u1_n129 ) , .A2( u1_u3_u1_n95 ) , .A1( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U51 (.A1( u1_u3_u1_n102 ) , .ZN( u1_u3_u1_n154 ) , .A2( u1_u3_u1_n99 ) );
  NAND2_X1 u1_u3_u1_U52 (.A2( u1_u3_u1_n100 ) , .ZN( u1_u3_u1_n135 ) , .A1( u1_u3_u1_n99 ) );
  AOI21_X1 u1_u3_u1_U53 (.A( u1_u3_u1_n152 ) , .B2( u1_u3_u1_n153 ) , .B1( u1_u3_u1_n154 ) , .ZN( u1_u3_u1_n158 ) );
  INV_X1 u1_u3_u1_U54 (.A( u1_u3_u1_n160 ) , .ZN( u1_u3_u1_n175 ) );
  NAND2_X1 u1_u3_u1_U55 (.A1( u1_u3_u1_n100 ) , .ZN( u1_u3_u1_n116 ) , .A2( u1_u3_u1_n95 ) );
  NAND2_X1 u1_u3_u1_U56 (.A1( u1_u3_u1_n102 ) , .ZN( u1_u3_u1_n131 ) , .A2( u1_u3_u1_n95 ) );
  NAND2_X1 u1_u3_u1_U57 (.A2( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n121 ) , .A1( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U58 (.A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n153 ) , .A2( u1_u3_u1_n98 ) );
  NAND2_X1 u1_u3_u1_U59 (.A2( u1_u3_u1_n104 ) , .A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n133 ) );
  AOI22_X1 u1_u3_u1_U6 (.B2( u1_u3_u1_n136 ) , .A2( u1_u3_u1_n137 ) , .ZN( u1_u3_u1_n143 ) , .A1( u1_u3_u1_n171 ) , .B1( u1_u3_u1_n173 ) );
  NAND2_X1 u1_u3_u1_U60 (.ZN( u1_u3_u1_n150 ) , .A2( u1_u3_u1_n98 ) , .A1( u1_u3_u1_n99 ) );
  NAND2_X1 u1_u3_u1_U61 (.A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n155 ) , .A2( u1_u3_u1_n95 ) );
  OAI21_X1 u1_u3_u1_U62 (.ZN( u1_u3_u1_n109 ) , .B1( u1_u3_u1_n129 ) , .B2( u1_u3_u1_n160 ) , .A( u1_u3_u1_n167 ) );
  NAND2_X1 u1_u3_u1_U63 (.A2( u1_u3_u1_n100 ) , .A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n120 ) );
  NAND2_X1 u1_u3_u1_U64 (.A1( u1_u3_u1_n102 ) , .A2( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n115 ) );
  NAND2_X1 u1_u3_u1_U65 (.A2( u1_u3_u1_n100 ) , .A1( u1_u3_u1_n104 ) , .ZN( u1_u3_u1_n151 ) );
  NAND2_X1 u1_u3_u1_U66 (.A2( u1_u3_u1_n103 ) , .A1( u1_u3_u1_n105 ) , .ZN( u1_u3_u1_n161 ) );
  INV_X1 u1_u3_u1_U67 (.A( u1_u3_u1_n152 ) , .ZN( u1_u3_u1_n173 ) );
  INV_X1 u1_u3_u1_U68 (.A( u1_u3_u1_n128 ) , .ZN( u1_u3_u1_n172 ) );
  NAND2_X1 u1_u3_u1_U69 (.A2( u1_u3_u1_n102 ) , .A1( u1_u3_u1_n103 ) , .ZN( u1_u3_u1_n123 ) );
  INV_X1 u1_u3_u1_U7 (.A( u1_u3_u1_n147 ) , .ZN( u1_u3_u1_n181 ) );
  NOR2_X1 u1_u3_u1_U70 (.A2( u1_u3_X_7 ) , .A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n95 ) );
  NOR2_X1 u1_u3_u1_U71 (.A1( u1_u3_X_12 ) , .A2( u1_u3_X_9 ) , .ZN( u1_u3_u1_n100 ) );
  NOR2_X1 u1_u3_u1_U72 (.A2( u1_u3_X_8 ) , .A1( u1_u3_u1_n177 ) , .ZN( u1_u3_u1_n99 ) );
  NOR2_X1 u1_u3_u1_U73 (.A2( u1_u3_X_12 ) , .ZN( u1_u3_u1_n102 ) , .A1( u1_u3_u1_n176 ) );
  NOR2_X1 u1_u3_u1_U74 (.A2( u1_u3_X_9 ) , .ZN( u1_u3_u1_n105 ) , .A1( u1_u3_u1_n168 ) );
  NAND2_X1 u1_u3_u1_U75 (.A1( u1_u3_X_10 ) , .ZN( u1_u3_u1_n160 ) , .A2( u1_u3_u1_n169 ) );
  NAND2_X1 u1_u3_u1_U76 (.A2( u1_u3_X_10 ) , .A1( u1_u3_X_11 ) , .ZN( u1_u3_u1_n152 ) );
  NAND2_X1 u1_u3_u1_U77 (.A1( u1_u3_X_11 ) , .ZN( u1_u3_u1_n128 ) , .A2( u1_u3_u1_n170 ) );
  AND2_X1 u1_u3_u1_U78 (.A2( u1_u3_X_7 ) , .A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n104 ) );
  AND2_X1 u1_u3_u1_U79 (.A1( u1_u3_X_8 ) , .ZN( u1_u3_u1_n103 ) , .A2( u1_u3_u1_n177 ) );
  NOR2_X1 u1_u3_u1_U8 (.A1( u1_u3_u1_n112 ) , .A2( u1_u3_u1_n116 ) , .ZN( u1_u3_u1_n118 ) );
  INV_X1 u1_u3_u1_U80 (.A( u1_u3_X_10 ) , .ZN( u1_u3_u1_n170 ) );
  INV_X1 u1_u3_u1_U81 (.A( u1_u3_X_9 ) , .ZN( u1_u3_u1_n176 ) );
  INV_X1 u1_u3_u1_U82 (.A( u1_u3_X_11 ) , .ZN( u1_u3_u1_n169 ) );
  INV_X1 u1_u3_u1_U83 (.A( u1_u3_X_12 ) , .ZN( u1_u3_u1_n168 ) );
  INV_X1 u1_u3_u1_U84 (.A( u1_u3_X_7 ) , .ZN( u1_u3_u1_n177 ) );
  NAND4_X1 u1_u3_u1_U85 (.ZN( u1_out3_18 ) , .A4( u1_u3_u1_n165 ) , .A3( u1_u3_u1_n166 ) , .A1( u1_u3_u1_n167 ) , .A2( u1_u3_u1_n186 ) );
  AOI22_X1 u1_u3_u1_U86 (.B2( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n147 ) , .A2( u1_u3_u1_n148 ) , .ZN( u1_u3_u1_n166 ) , .A1( u1_u3_u1_n172 ) );
  INV_X1 u1_u3_u1_U87 (.A( u1_u3_u1_n145 ) , .ZN( u1_u3_u1_n186 ) );
  OR4_X1 u1_u3_u1_U88 (.ZN( u1_out3_13 ) , .A4( u1_u3_u1_n108 ) , .A3( u1_u3_u1_n109 ) , .A2( u1_u3_u1_n110 ) , .A1( u1_u3_u1_n111 ) );
  AOI21_X1 u1_u3_u1_U89 (.ZN( u1_u3_u1_n111 ) , .A( u1_u3_u1_n128 ) , .B2( u1_u3_u1_n131 ) , .B1( u1_u3_u1_n135 ) );
  OAI21_X1 u1_u3_u1_U9 (.ZN( u1_u3_u1_n101 ) , .B1( u1_u3_u1_n141 ) , .A( u1_u3_u1_n146 ) , .B2( u1_u3_u1_n183 ) );
  AOI21_X1 u1_u3_u1_U90 (.ZN( u1_u3_u1_n110 ) , .A( u1_u3_u1_n116 ) , .B1( u1_u3_u1_n152 ) , .B2( u1_u3_u1_n160 ) );
  NAND4_X1 u1_u3_u1_U91 (.ZN( u1_out3_2 ) , .A4( u1_u3_u1_n142 ) , .A3( u1_u3_u1_n143 ) , .A2( u1_u3_u1_n144 ) , .A1( u1_u3_u1_n179 ) );
  INV_X1 u1_u3_u1_U92 (.A( u1_u3_u1_n130 ) , .ZN( u1_u3_u1_n179 ) );
  OAI21_X1 u1_u3_u1_U93 (.B2( u1_u3_u1_n132 ) , .ZN( u1_u3_u1_n144 ) , .A( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n180 ) );
  NAND4_X1 u1_u3_u1_U94 (.ZN( u1_out3_28 ) , .A4( u1_u3_u1_n124 ) , .A3( u1_u3_u1_n125 ) , .A2( u1_u3_u1_n126 ) , .A1( u1_u3_u1_n127 ) );
  OAI21_X1 u1_u3_u1_U95 (.ZN( u1_u3_u1_n127 ) , .B2( u1_u3_u1_n139 ) , .B1( u1_u3_u1_n175 ) , .A( u1_u3_u1_n183 ) );
  OAI21_X1 u1_u3_u1_U96 (.ZN( u1_u3_u1_n126 ) , .B2( u1_u3_u1_n140 ) , .A( u1_u3_u1_n146 ) , .B1( u1_u3_u1_n178 ) );
  NAND3_X1 u1_u3_u1_U97 (.A3( u1_u3_u1_n149 ) , .A2( u1_u3_u1_n150 ) , .A1( u1_u3_u1_n151 ) , .ZN( u1_u3_u1_n164 ) );
  NAND3_X1 u1_u3_u1_U98 (.A3( u1_u3_u1_n134 ) , .A2( u1_u3_u1_n135 ) , .ZN( u1_u3_u1_n136 ) , .A1( u1_u3_u1_n151 ) );
  NAND3_X1 u1_u3_u1_U99 (.A1( u1_u3_u1_n133 ) , .ZN( u1_u3_u1_n137 ) , .A2( u1_u3_u1_n154 ) , .A3( u1_u3_u1_n181 ) );
  XOR2_X1 u1_u4_U20 (.B( u1_K5_36 ) , .A( u1_R3_25 ) , .Z( u1_u4_X_36 ) );
  XOR2_X1 u1_u4_U21 (.B( u1_K5_35 ) , .A( u1_R3_24 ) , .Z( u1_u4_X_35 ) );
  XOR2_X1 u1_u4_U22 (.B( u1_K5_34 ) , .A( u1_R3_23 ) , .Z( u1_u4_X_34 ) );
  XOR2_X1 u1_u4_U23 (.B( u1_K5_33 ) , .A( u1_R3_22 ) , .Z( u1_u4_X_33 ) );
  XOR2_X1 u1_u4_U24 (.B( u1_K5_32 ) , .A( u1_R3_21 ) , .Z( u1_u4_X_32 ) );
  XOR2_X1 u1_u4_U25 (.B( u1_K5_31 ) , .A( u1_R3_20 ) , .Z( u1_u4_X_31 ) );
  NOR2_X1 u1_u4_u5_U10 (.ZN( u1_u4_u5_n135 ) , .A1( u1_u4_u5_n173 ) , .A2( u1_u4_u5_n176 ) );
  NOR3_X1 u1_u4_u5_U100 (.A3( u1_u4_u5_n141 ) , .A1( u1_u4_u5_n142 ) , .ZN( u1_u4_u5_n143 ) , .A2( u1_u4_u5_n191 ) );
  NAND4_X1 u1_u4_u5_U101 (.ZN( u1_out4_4 ) , .A4( u1_u4_u5_n112 ) , .A2( u1_u4_u5_n113 ) , .A1( u1_u4_u5_n114 ) , .A3( u1_u4_u5_n195 ) );
  AOI211_X1 u1_u4_u5_U102 (.A( u1_u4_u5_n110 ) , .C1( u1_u4_u5_n111 ) , .ZN( u1_u4_u5_n112 ) , .B( u1_u4_u5_n118 ) , .C2( u1_u4_u5_n177 ) );
  INV_X1 u1_u4_u5_U103 (.A( u1_u4_u5_n102 ) , .ZN( u1_u4_u5_n195 ) );
  NAND3_X1 u1_u4_u5_U104 (.A2( u1_u4_u5_n154 ) , .A3( u1_u4_u5_n158 ) , .A1( u1_u4_u5_n161 ) , .ZN( u1_u4_u5_n99 ) );
  INV_X1 u1_u4_u5_U11 (.A( u1_u4_u5_n121 ) , .ZN( u1_u4_u5_n177 ) );
  NOR2_X1 u1_u4_u5_U12 (.ZN( u1_u4_u5_n160 ) , .A2( u1_u4_u5_n173 ) , .A1( u1_u4_u5_n177 ) );
  INV_X1 u1_u4_u5_U13 (.A( u1_u4_u5_n150 ) , .ZN( u1_u4_u5_n174 ) );
  AOI21_X1 u1_u4_u5_U14 (.A( u1_u4_u5_n160 ) , .B2( u1_u4_u5_n161 ) , .ZN( u1_u4_u5_n162 ) , .B1( u1_u4_u5_n192 ) );
  INV_X1 u1_u4_u5_U15 (.A( u1_u4_u5_n159 ) , .ZN( u1_u4_u5_n192 ) );
  AOI21_X1 u1_u4_u5_U16 (.A( u1_u4_u5_n156 ) , .B2( u1_u4_u5_n157 ) , .B1( u1_u4_u5_n158 ) , .ZN( u1_u4_u5_n163 ) );
  AOI21_X1 u1_u4_u5_U17 (.B2( u1_u4_u5_n139 ) , .B1( u1_u4_u5_n140 ) , .ZN( u1_u4_u5_n141 ) , .A( u1_u4_u5_n150 ) );
  OAI21_X1 u1_u4_u5_U18 (.A( u1_u4_u5_n133 ) , .B2( u1_u4_u5_n134 ) , .B1( u1_u4_u5_n135 ) , .ZN( u1_u4_u5_n142 ) );
  OAI21_X1 u1_u4_u5_U19 (.ZN( u1_u4_u5_n133 ) , .B2( u1_u4_u5_n147 ) , .A( u1_u4_u5_n173 ) , .B1( u1_u4_u5_n188 ) );
  NAND2_X1 u1_u4_u5_U20 (.A2( u1_u4_u5_n119 ) , .A1( u1_u4_u5_n123 ) , .ZN( u1_u4_u5_n137 ) );
  INV_X1 u1_u4_u5_U21 (.A( u1_u4_u5_n155 ) , .ZN( u1_u4_u5_n194 ) );
  NAND2_X1 u1_u4_u5_U22 (.A1( u1_u4_u5_n121 ) , .ZN( u1_u4_u5_n132 ) , .A2( u1_u4_u5_n172 ) );
  NAND2_X1 u1_u4_u5_U23 (.A2( u1_u4_u5_n122 ) , .ZN( u1_u4_u5_n136 ) , .A1( u1_u4_u5_n154 ) );
  NAND2_X1 u1_u4_u5_U24 (.A2( u1_u4_u5_n119 ) , .A1( u1_u4_u5_n120 ) , .ZN( u1_u4_u5_n159 ) );
  INV_X1 u1_u4_u5_U25 (.A( u1_u4_u5_n156 ) , .ZN( u1_u4_u5_n175 ) );
  INV_X1 u1_u4_u5_U26 (.A( u1_u4_u5_n158 ) , .ZN( u1_u4_u5_n188 ) );
  INV_X1 u1_u4_u5_U27 (.A( u1_u4_u5_n152 ) , .ZN( u1_u4_u5_n179 ) );
  INV_X1 u1_u4_u5_U28 (.A( u1_u4_u5_n140 ) , .ZN( u1_u4_u5_n182 ) );
  INV_X1 u1_u4_u5_U29 (.A( u1_u4_u5_n151 ) , .ZN( u1_u4_u5_n183 ) );
  NOR2_X1 u1_u4_u5_U3 (.ZN( u1_u4_u5_n134 ) , .A1( u1_u4_u5_n183 ) , .A2( u1_u4_u5_n190 ) );
  INV_X1 u1_u4_u5_U30 (.A( u1_u4_u5_n123 ) , .ZN( u1_u4_u5_n185 ) );
  INV_X1 u1_u4_u5_U31 (.A( u1_u4_u5_n161 ) , .ZN( u1_u4_u5_n184 ) );
  INV_X1 u1_u4_u5_U32 (.A( u1_u4_u5_n139 ) , .ZN( u1_u4_u5_n189 ) );
  INV_X1 u1_u4_u5_U33 (.A( u1_u4_u5_n157 ) , .ZN( u1_u4_u5_n190 ) );
  INV_X1 u1_u4_u5_U34 (.A( u1_u4_u5_n120 ) , .ZN( u1_u4_u5_n193 ) );
  NAND2_X1 u1_u4_u5_U35 (.ZN( u1_u4_u5_n111 ) , .A1( u1_u4_u5_n140 ) , .A2( u1_u4_u5_n155 ) );
  INV_X1 u1_u4_u5_U36 (.A( u1_u4_u5_n117 ) , .ZN( u1_u4_u5_n196 ) );
  OAI221_X1 u1_u4_u5_U37 (.A( u1_u4_u5_n116 ) , .ZN( u1_u4_u5_n117 ) , .B2( u1_u4_u5_n119 ) , .C1( u1_u4_u5_n153 ) , .C2( u1_u4_u5_n158 ) , .B1( u1_u4_u5_n172 ) );
  AOI222_X1 u1_u4_u5_U38 (.ZN( u1_u4_u5_n116 ) , .B2( u1_u4_u5_n145 ) , .C1( u1_u4_u5_n148 ) , .A2( u1_u4_u5_n174 ) , .C2( u1_u4_u5_n177 ) , .B1( u1_u4_u5_n187 ) , .A1( u1_u4_u5_n193 ) );
  INV_X1 u1_u4_u5_U39 (.A( u1_u4_u5_n115 ) , .ZN( u1_u4_u5_n187 ) );
  INV_X1 u1_u4_u5_U4 (.A( u1_u4_u5_n138 ) , .ZN( u1_u4_u5_n191 ) );
  NOR2_X1 u1_u4_u5_U40 (.ZN( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n170 ) , .A2( u1_u4_u5_n180 ) );
  OAI221_X1 u1_u4_u5_U41 (.A( u1_u4_u5_n101 ) , .ZN( u1_u4_u5_n102 ) , .C2( u1_u4_u5_n115 ) , .C1( u1_u4_u5_n126 ) , .B1( u1_u4_u5_n134 ) , .B2( u1_u4_u5_n160 ) );
  OAI21_X1 u1_u4_u5_U42 (.ZN( u1_u4_u5_n101 ) , .B1( u1_u4_u5_n137 ) , .A( u1_u4_u5_n146 ) , .B2( u1_u4_u5_n147 ) );
  AOI22_X1 u1_u4_u5_U43 (.B2( u1_u4_u5_n131 ) , .A2( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n169 ) , .B1( u1_u4_u5_n174 ) , .A1( u1_u4_u5_n185 ) );
  NOR2_X1 u1_u4_u5_U44 (.A1( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n150 ) , .A2( u1_u4_u5_n173 ) );
  AOI21_X1 u1_u4_u5_U45 (.A( u1_u4_u5_n118 ) , .B2( u1_u4_u5_n145 ) , .ZN( u1_u4_u5_n168 ) , .B1( u1_u4_u5_n186 ) );
  INV_X1 u1_u4_u5_U46 (.A( u1_u4_u5_n122 ) , .ZN( u1_u4_u5_n186 ) );
  NOR2_X1 u1_u4_u5_U47 (.A1( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n152 ) , .A2( u1_u4_u5_n176 ) );
  NOR2_X1 u1_u4_u5_U48 (.A1( u1_u4_u5_n115 ) , .ZN( u1_u4_u5_n118 ) , .A2( u1_u4_u5_n153 ) );
  NOR2_X1 u1_u4_u5_U49 (.A2( u1_u4_u5_n145 ) , .ZN( u1_u4_u5_n156 ) , .A1( u1_u4_u5_n174 ) );
  OAI21_X1 u1_u4_u5_U5 (.B2( u1_u4_u5_n136 ) , .B1( u1_u4_u5_n137 ) , .ZN( u1_u4_u5_n138 ) , .A( u1_u4_u5_n177 ) );
  NOR2_X1 u1_u4_u5_U50 (.ZN( u1_u4_u5_n121 ) , .A2( u1_u4_u5_n145 ) , .A1( u1_u4_u5_n176 ) );
  AOI22_X1 u1_u4_u5_U51 (.ZN( u1_u4_u5_n114 ) , .A2( u1_u4_u5_n137 ) , .A1( u1_u4_u5_n145 ) , .B2( u1_u4_u5_n175 ) , .B1( u1_u4_u5_n193 ) );
  OAI211_X1 u1_u4_u5_U52 (.B( u1_u4_u5_n124 ) , .A( u1_u4_u5_n125 ) , .C2( u1_u4_u5_n126 ) , .C1( u1_u4_u5_n127 ) , .ZN( u1_u4_u5_n128 ) );
  NOR3_X1 u1_u4_u5_U53 (.ZN( u1_u4_u5_n127 ) , .A1( u1_u4_u5_n136 ) , .A3( u1_u4_u5_n148 ) , .A2( u1_u4_u5_n182 ) );
  OAI21_X1 u1_u4_u5_U54 (.ZN( u1_u4_u5_n124 ) , .A( u1_u4_u5_n177 ) , .B2( u1_u4_u5_n183 ) , .B1( u1_u4_u5_n189 ) );
  OAI21_X1 u1_u4_u5_U55 (.ZN( u1_u4_u5_n125 ) , .A( u1_u4_u5_n174 ) , .B2( u1_u4_u5_n185 ) , .B1( u1_u4_u5_n190 ) );
  AOI21_X1 u1_u4_u5_U56 (.A( u1_u4_u5_n153 ) , .B2( u1_u4_u5_n154 ) , .B1( u1_u4_u5_n155 ) , .ZN( u1_u4_u5_n164 ) );
  AOI21_X1 u1_u4_u5_U57 (.ZN( u1_u4_u5_n110 ) , .B1( u1_u4_u5_n122 ) , .B2( u1_u4_u5_n139 ) , .A( u1_u4_u5_n153 ) );
  INV_X1 u1_u4_u5_U58 (.A( u1_u4_u5_n153 ) , .ZN( u1_u4_u5_n176 ) );
  INV_X1 u1_u4_u5_U59 (.A( u1_u4_u5_n126 ) , .ZN( u1_u4_u5_n173 ) );
  AOI222_X1 u1_u4_u5_U6 (.ZN( u1_u4_u5_n113 ) , .A1( u1_u4_u5_n131 ) , .C1( u1_u4_u5_n148 ) , .B2( u1_u4_u5_n174 ) , .C2( u1_u4_u5_n178 ) , .A2( u1_u4_u5_n179 ) , .B1( u1_u4_u5_n99 ) );
  AND2_X1 u1_u4_u5_U60 (.A2( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n107 ) , .ZN( u1_u4_u5_n147 ) );
  AND2_X1 u1_u4_u5_U61 (.A2( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n108 ) , .ZN( u1_u4_u5_n148 ) );
  NAND2_X1 u1_u4_u5_U62 (.A1( u1_u4_u5_n105 ) , .A2( u1_u4_u5_n106 ) , .ZN( u1_u4_u5_n158 ) );
  NAND2_X1 u1_u4_u5_U63 (.A2( u1_u4_u5_n108 ) , .A1( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n139 ) );
  NAND2_X1 u1_u4_u5_U64 (.A1( u1_u4_u5_n106 ) , .A2( u1_u4_u5_n108 ) , .ZN( u1_u4_u5_n119 ) );
  NAND2_X1 u1_u4_u5_U65 (.A2( u1_u4_u5_n103 ) , .A1( u1_u4_u5_n105 ) , .ZN( u1_u4_u5_n140 ) );
  NAND2_X1 u1_u4_u5_U66 (.A2( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n105 ) , .ZN( u1_u4_u5_n155 ) );
  NAND2_X1 u1_u4_u5_U67 (.A2( u1_u4_u5_n106 ) , .A1( u1_u4_u5_n107 ) , .ZN( u1_u4_u5_n122 ) );
  NAND2_X1 u1_u4_u5_U68 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n106 ) , .ZN( u1_u4_u5_n115 ) );
  NAND2_X1 u1_u4_u5_U69 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n103 ) , .ZN( u1_u4_u5_n161 ) );
  INV_X1 u1_u4_u5_U7 (.A( u1_u4_u5_n135 ) , .ZN( u1_u4_u5_n178 ) );
  NAND2_X1 u1_u4_u5_U70 (.A1( u1_u4_u5_n105 ) , .A2( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n154 ) );
  INV_X1 u1_u4_u5_U71 (.A( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n172 ) );
  NAND2_X1 u1_u4_u5_U72 (.A1( u1_u4_u5_n103 ) , .A2( u1_u4_u5_n108 ) , .ZN( u1_u4_u5_n123 ) );
  NAND2_X1 u1_u4_u5_U73 (.A2( u1_u4_u5_n103 ) , .A1( u1_u4_u5_n107 ) , .ZN( u1_u4_u5_n151 ) );
  NAND2_X1 u1_u4_u5_U74 (.A2( u1_u4_u5_n107 ) , .A1( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n120 ) );
  NAND2_X1 u1_u4_u5_U75 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n157 ) );
  AND2_X1 u1_u4_u5_U76 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n104 ) , .ZN( u1_u4_u5_n131 ) );
  NOR2_X1 u1_u4_u5_U77 (.A2( u1_u4_X_34 ) , .A1( u1_u4_X_35 ) , .ZN( u1_u4_u5_n145 ) );
  NOR2_X1 u1_u4_u5_U78 (.A2( u1_u4_X_34 ) , .ZN( u1_u4_u5_n146 ) , .A1( u1_u4_u5_n171 ) );
  NOR2_X1 u1_u4_u5_U79 (.A2( u1_u4_X_31 ) , .A1( u1_u4_X_32 ) , .ZN( u1_u4_u5_n103 ) );
  OAI22_X1 u1_u4_u5_U8 (.B2( u1_u4_u5_n149 ) , .B1( u1_u4_u5_n150 ) , .A2( u1_u4_u5_n151 ) , .A1( u1_u4_u5_n152 ) , .ZN( u1_u4_u5_n165 ) );
  NOR2_X1 u1_u4_u5_U80 (.A2( u1_u4_X_36 ) , .ZN( u1_u4_u5_n105 ) , .A1( u1_u4_u5_n180 ) );
  NOR2_X1 u1_u4_u5_U81 (.A2( u1_u4_X_33 ) , .ZN( u1_u4_u5_n108 ) , .A1( u1_u4_u5_n170 ) );
  NOR2_X1 u1_u4_u5_U82 (.A2( u1_u4_X_33 ) , .A1( u1_u4_X_36 ) , .ZN( u1_u4_u5_n107 ) );
  NOR2_X1 u1_u4_u5_U83 (.A2( u1_u4_X_31 ) , .ZN( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n181 ) );
  NAND2_X1 u1_u4_u5_U84 (.A2( u1_u4_X_34 ) , .A1( u1_u4_X_35 ) , .ZN( u1_u4_u5_n153 ) );
  NAND2_X1 u1_u4_u5_U85 (.A1( u1_u4_X_34 ) , .ZN( u1_u4_u5_n126 ) , .A2( u1_u4_u5_n171 ) );
  AND2_X1 u1_u4_u5_U86 (.A1( u1_u4_X_31 ) , .A2( u1_u4_X_32 ) , .ZN( u1_u4_u5_n106 ) );
  AND2_X1 u1_u4_u5_U87 (.A1( u1_u4_X_31 ) , .ZN( u1_u4_u5_n109 ) , .A2( u1_u4_u5_n181 ) );
  INV_X1 u1_u4_u5_U88 (.A( u1_u4_X_33 ) , .ZN( u1_u4_u5_n180 ) );
  INV_X1 u1_u4_u5_U89 (.A( u1_u4_X_35 ) , .ZN( u1_u4_u5_n171 ) );
  NOR3_X1 u1_u4_u5_U9 (.A2( u1_u4_u5_n147 ) , .A1( u1_u4_u5_n148 ) , .ZN( u1_u4_u5_n149 ) , .A3( u1_u4_u5_n194 ) );
  INV_X1 u1_u4_u5_U90 (.A( u1_u4_X_36 ) , .ZN( u1_u4_u5_n170 ) );
  INV_X1 u1_u4_u5_U91 (.A( u1_u4_X_32 ) , .ZN( u1_u4_u5_n181 ) );
  NAND4_X1 u1_u4_u5_U92 (.ZN( u1_out4_29 ) , .A4( u1_u4_u5_n129 ) , .A3( u1_u4_u5_n130 ) , .A2( u1_u4_u5_n168 ) , .A1( u1_u4_u5_n196 ) );
  AOI221_X1 u1_u4_u5_U93 (.A( u1_u4_u5_n128 ) , .ZN( u1_u4_u5_n129 ) , .C2( u1_u4_u5_n132 ) , .B2( u1_u4_u5_n159 ) , .B1( u1_u4_u5_n176 ) , .C1( u1_u4_u5_n184 ) );
  AOI222_X1 u1_u4_u5_U94 (.ZN( u1_u4_u5_n130 ) , .A2( u1_u4_u5_n146 ) , .B1( u1_u4_u5_n147 ) , .C2( u1_u4_u5_n175 ) , .B2( u1_u4_u5_n179 ) , .A1( u1_u4_u5_n188 ) , .C1( u1_u4_u5_n194 ) );
  NAND4_X1 u1_u4_u5_U95 (.ZN( u1_out4_19 ) , .A4( u1_u4_u5_n166 ) , .A3( u1_u4_u5_n167 ) , .A2( u1_u4_u5_n168 ) , .A1( u1_u4_u5_n169 ) );
  AOI22_X1 u1_u4_u5_U96 (.B2( u1_u4_u5_n145 ) , .A2( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n167 ) , .B1( u1_u4_u5_n182 ) , .A1( u1_u4_u5_n189 ) );
  NOR4_X1 u1_u4_u5_U97 (.A4( u1_u4_u5_n162 ) , .A3( u1_u4_u5_n163 ) , .A2( u1_u4_u5_n164 ) , .A1( u1_u4_u5_n165 ) , .ZN( u1_u4_u5_n166 ) );
  NAND4_X1 u1_u4_u5_U98 (.ZN( u1_out4_11 ) , .A4( u1_u4_u5_n143 ) , .A3( u1_u4_u5_n144 ) , .A2( u1_u4_u5_n169 ) , .A1( u1_u4_u5_n196 ) );
  AOI22_X1 u1_u4_u5_U99 (.A2( u1_u4_u5_n132 ) , .ZN( u1_u4_u5_n144 ) , .B2( u1_u4_u5_n145 ) , .B1( u1_u4_u5_n184 ) , .A1( u1_u4_u5_n194 ) );
  XOR2_X1 u1_u5_U13 (.B( u1_K6_42 ) , .A( u1_R4_29 ) , .Z( u1_u5_X_42 ) );
  XOR2_X1 u1_u5_U14 (.B( u1_K6_41 ) , .A( u1_R4_28 ) , .Z( u1_u5_X_41 ) );
  XOR2_X1 u1_u5_U15 (.B( u1_K6_40 ) , .A( u1_R4_27 ) , .Z( u1_u5_X_40 ) );
  XOR2_X1 u1_u5_U16 (.B( u1_K6_3 ) , .A( u1_R4_2 ) , .Z( u1_u5_X_3 ) );
  XOR2_X1 u1_u5_U17 (.B( u1_K6_39 ) , .A( u1_R4_26 ) , .Z( u1_u5_X_39 ) );
  XOR2_X1 u1_u5_U18 (.B( u1_K6_38 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_38 ) );
  XOR2_X1 u1_u5_U19 (.B( u1_K6_37 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_37 ) );
  XOR2_X1 u1_u5_U20 (.B( u1_K6_36 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_36 ) );
  XOR2_X1 u1_u5_U21 (.B( u1_K6_35 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_35 ) );
  XOR2_X1 u1_u5_U22 (.B( u1_K6_34 ) , .A( u1_R4_23 ) , .Z( u1_u5_X_34 ) );
  XOR2_X1 u1_u5_U23 (.B( u1_K6_33 ) , .A( u1_R4_22 ) , .Z( u1_u5_X_33 ) );
  XOR2_X1 u1_u5_U24 (.B( u1_K6_32 ) , .A( u1_R4_21 ) , .Z( u1_u5_X_32 ) );
  XOR2_X1 u1_u5_U25 (.B( u1_K6_31 ) , .A( u1_R4_20 ) , .Z( u1_u5_X_31 ) );
  XOR2_X1 u1_u5_U26 (.B( u1_K6_30 ) , .A( u1_R4_21 ) , .Z( u1_u5_X_30 ) );
  XOR2_X1 u1_u5_U27 (.B( u1_K6_2 ) , .A( u1_R4_1 ) , .Z( u1_u5_X_2 ) );
  XOR2_X1 u1_u5_U28 (.B( u1_K6_29 ) , .A( u1_R4_20 ) , .Z( u1_u5_X_29 ) );
  XOR2_X1 u1_u5_U29 (.B( u1_K6_28 ) , .A( u1_R4_19 ) , .Z( u1_u5_X_28 ) );
  XOR2_X1 u1_u5_U30 (.B( u1_K6_27 ) , .A( u1_R4_18 ) , .Z( u1_u5_X_27 ) );
  XOR2_X1 u1_u5_U31 (.B( u1_K6_26 ) , .A( u1_R4_17 ) , .Z( u1_u5_X_26 ) );
  XOR2_X1 u1_u5_U32 (.B( u1_K6_25 ) , .A( u1_R4_16 ) , .Z( u1_u5_X_25 ) );
  XOR2_X1 u1_u5_U33 (.B( u1_K6_24 ) , .A( u1_R4_17 ) , .Z( u1_u5_X_24 ) );
  XOR2_X1 u1_u5_U34 (.B( u1_K6_23 ) , .A( u1_R4_16 ) , .Z( u1_u5_X_23 ) );
  XOR2_X1 u1_u5_U35 (.B( u1_K6_22 ) , .A( u1_R4_15 ) , .Z( u1_u5_X_22 ) );
  XOR2_X1 u1_u5_U36 (.B( u1_K6_21 ) , .A( u1_R4_14 ) , .Z( u1_u5_X_21 ) );
  XOR2_X1 u1_u5_U37 (.B( u1_K6_20 ) , .A( u1_R4_13 ) , .Z( u1_u5_X_20 ) );
  XOR2_X1 u1_u5_U38 (.B( u1_K6_1 ) , .A( u1_R4_32 ) , .Z( u1_u5_X_1 ) );
  XOR2_X1 u1_u5_U39 (.B( u1_K6_19 ) , .A( u1_R4_12 ) , .Z( u1_u5_X_19 ) );
  XOR2_X1 u1_u5_U4 (.B( u1_K6_6 ) , .A( u1_R4_5 ) , .Z( u1_u5_X_6 ) );
  XOR2_X1 u1_u5_U40 (.B( u1_K6_18 ) , .A( u1_R4_13 ) , .Z( u1_u5_X_18 ) );
  XOR2_X1 u1_u5_U41 (.B( u1_K6_17 ) , .A( u1_R4_12 ) , .Z( u1_u5_X_17 ) );
  XOR2_X1 u1_u5_U42 (.B( u1_K6_16 ) , .A( u1_R4_11 ) , .Z( u1_u5_X_16 ) );
  XOR2_X1 u1_u5_U43 (.B( u1_K6_15 ) , .A( u1_R4_10 ) , .Z( u1_u5_X_15 ) );
  XOR2_X1 u1_u5_U44 (.B( u1_K6_14 ) , .A( u1_R4_9 ) , .Z( u1_u5_X_14 ) );
  XOR2_X1 u1_u5_U45 (.B( u1_K6_13 ) , .A( u1_R4_8 ) , .Z( u1_u5_X_13 ) );
  XOR2_X1 u1_u5_U5 (.B( u1_K6_5 ) , .A( u1_R4_4 ) , .Z( u1_u5_X_5 ) );
  XOR2_X1 u1_u5_U6 (.B( u1_K6_4 ) , .A( u1_R4_3 ) , .Z( u1_u5_X_4 ) );
  NAND2_X1 u1_u5_u0_U10 (.ZN( u1_u5_u0_n113 ) , .A1( u1_u5_u0_n139 ) , .A2( u1_u5_u0_n149 ) );
  AND3_X1 u1_u5_u0_U11 (.A2( u1_u5_u0_n112 ) , .ZN( u1_u5_u0_n127 ) , .A3( u1_u5_u0_n130 ) , .A1( u1_u5_u0_n148 ) );
  AND2_X1 u1_u5_u0_U12 (.ZN( u1_u5_u0_n107 ) , .A1( u1_u5_u0_n130 ) , .A2( u1_u5_u0_n140 ) );
  AND2_X1 u1_u5_u0_U13 (.A2( u1_u5_u0_n129 ) , .A1( u1_u5_u0_n130 ) , .ZN( u1_u5_u0_n151 ) );
  AND2_X1 u1_u5_u0_U14 (.A1( u1_u5_u0_n108 ) , .A2( u1_u5_u0_n125 ) , .ZN( u1_u5_u0_n145 ) );
  INV_X1 u1_u5_u0_U15 (.A( u1_u5_u0_n143 ) , .ZN( u1_u5_u0_n173 ) );
  NOR2_X1 u1_u5_u0_U16 (.A2( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n147 ) , .A1( u1_u5_u0_n160 ) );
  AOI21_X1 u1_u5_u0_U17 (.B1( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n132 ) , .A( u1_u5_u0_n165 ) , .B2( u1_u5_u0_n93 ) );
  INV_X1 u1_u5_u0_U18 (.A( u1_u5_u0_n142 ) , .ZN( u1_u5_u0_n165 ) );
  OAI22_X1 u1_u5_u0_U19 (.B1( u1_u5_u0_n131 ) , .A1( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n147 ) , .A2( u1_u5_u0_n90 ) , .ZN( u1_u5_u0_n91 ) );
  AND3_X1 u1_u5_u0_U20 (.A3( u1_u5_u0_n121 ) , .A2( u1_u5_u0_n125 ) , .A1( u1_u5_u0_n148 ) , .ZN( u1_u5_u0_n90 ) );
  OAI22_X1 u1_u5_u0_U21 (.B1( u1_u5_u0_n125 ) , .ZN( u1_u5_u0_n126 ) , .A1( u1_u5_u0_n138 ) , .A2( u1_u5_u0_n146 ) , .B2( u1_u5_u0_n147 ) );
  NOR2_X1 u1_u5_u0_U22 (.A1( u1_u5_u0_n163 ) , .A2( u1_u5_u0_n164 ) , .ZN( u1_u5_u0_n95 ) );
  INV_X1 u1_u5_u0_U23 (.A( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n161 ) );
  AOI22_X1 u1_u5_u0_U24 (.B2( u1_u5_u0_n109 ) , .A2( u1_u5_u0_n110 ) , .ZN( u1_u5_u0_n111 ) , .B1( u1_u5_u0_n118 ) , .A1( u1_u5_u0_n160 ) );
  NAND2_X1 u1_u5_u0_U25 (.A2( u1_u5_u0_n102 ) , .A1( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n149 ) );
  INV_X1 u1_u5_u0_U26 (.A( u1_u5_u0_n118 ) , .ZN( u1_u5_u0_n158 ) );
  NAND2_X1 u1_u5_u0_U27 (.A2( u1_u5_u0_n100 ) , .ZN( u1_u5_u0_n131 ) , .A1( u1_u5_u0_n92 ) );
  NAND2_X1 u1_u5_u0_U28 (.ZN( u1_u5_u0_n108 ) , .A1( u1_u5_u0_n92 ) , .A2( u1_u5_u0_n94 ) );
  AOI21_X1 u1_u5_u0_U29 (.ZN( u1_u5_u0_n104 ) , .B1( u1_u5_u0_n107 ) , .B2( u1_u5_u0_n141 ) , .A( u1_u5_u0_n144 ) );
  INV_X1 u1_u5_u0_U3 (.A( u1_u5_u0_n113 ) , .ZN( u1_u5_u0_n166 ) );
  AOI21_X1 u1_u5_u0_U30 (.B1( u1_u5_u0_n127 ) , .B2( u1_u5_u0_n129 ) , .A( u1_u5_u0_n138 ) , .ZN( u1_u5_u0_n96 ) );
  NAND2_X1 u1_u5_u0_U31 (.A2( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n114 ) , .A1( u1_u5_u0_n92 ) );
  AOI21_X1 u1_u5_u0_U32 (.ZN( u1_u5_u0_n116 ) , .B2( u1_u5_u0_n142 ) , .A( u1_u5_u0_n144 ) , .B1( u1_u5_u0_n166 ) );
  NOR2_X1 u1_u5_u0_U33 (.A1( u1_u5_u0_n120 ) , .ZN( u1_u5_u0_n143 ) , .A2( u1_u5_u0_n167 ) );
  OAI221_X1 u1_u5_u0_U34 (.C1( u1_u5_u0_n112 ) , .ZN( u1_u5_u0_n120 ) , .B1( u1_u5_u0_n138 ) , .B2( u1_u5_u0_n141 ) , .C2( u1_u5_u0_n147 ) , .A( u1_u5_u0_n172 ) );
  AOI211_X1 u1_u5_u0_U35 (.B( u1_u5_u0_n115 ) , .A( u1_u5_u0_n116 ) , .C2( u1_u5_u0_n117 ) , .C1( u1_u5_u0_n118 ) , .ZN( u1_u5_u0_n119 ) );
  NAND2_X1 u1_u5_u0_U36 (.A2( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n140 ) , .A1( u1_u5_u0_n94 ) );
  NAND2_X1 u1_u5_u0_U37 (.A1( u1_u5_u0_n100 ) , .A2( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n125 ) );
  NAND2_X1 u1_u5_u0_U38 (.A1( u1_u5_u0_n101 ) , .A2( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n150 ) );
  INV_X1 u1_u5_u0_U39 (.A( u1_u5_u0_n138 ) , .ZN( u1_u5_u0_n160 ) );
  AOI21_X1 u1_u5_u0_U4 (.B1( u1_u5_u0_n114 ) , .ZN( u1_u5_u0_n115 ) , .B2( u1_u5_u0_n129 ) , .A( u1_u5_u0_n161 ) );
  NAND2_X1 u1_u5_u0_U40 (.A2( u1_u5_u0_n100 ) , .A1( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n139 ) );
  NAND2_X1 u1_u5_u0_U41 (.ZN( u1_u5_u0_n112 ) , .A2( u1_u5_u0_n92 ) , .A1( u1_u5_u0_n93 ) );
  NAND2_X1 u1_u5_u0_U42 (.A1( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n130 ) , .A2( u1_u5_u0_n94 ) );
  INV_X1 u1_u5_u0_U43 (.ZN( u1_u5_u0_n172 ) , .A( u1_u5_u0_n88 ) );
  OAI222_X1 u1_u5_u0_U44 (.C1( u1_u5_u0_n108 ) , .A1( u1_u5_u0_n125 ) , .B2( u1_u5_u0_n128 ) , .B1( u1_u5_u0_n144 ) , .A2( u1_u5_u0_n158 ) , .C2( u1_u5_u0_n161 ) , .ZN( u1_u5_u0_n88 ) );
  NAND2_X1 u1_u5_u0_U45 (.A2( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n121 ) , .A1( u1_u5_u0_n93 ) );
  OR3_X1 u1_u5_u0_U46 (.A3( u1_u5_u0_n152 ) , .A2( u1_u5_u0_n153 ) , .A1( u1_u5_u0_n154 ) , .ZN( u1_u5_u0_n155 ) );
  AOI21_X1 u1_u5_u0_U47 (.A( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n145 ) , .B1( u1_u5_u0_n146 ) , .ZN( u1_u5_u0_n154 ) );
  AOI21_X1 u1_u5_u0_U48 (.B2( u1_u5_u0_n150 ) , .B1( u1_u5_u0_n151 ) , .ZN( u1_u5_u0_n152 ) , .A( u1_u5_u0_n158 ) );
  AOI21_X1 u1_u5_u0_U49 (.A( u1_u5_u0_n147 ) , .B2( u1_u5_u0_n148 ) , .B1( u1_u5_u0_n149 ) , .ZN( u1_u5_u0_n153 ) );
  AOI21_X1 u1_u5_u0_U5 (.B2( u1_u5_u0_n131 ) , .ZN( u1_u5_u0_n134 ) , .B1( u1_u5_u0_n151 ) , .A( u1_u5_u0_n158 ) );
  INV_X1 u1_u5_u0_U50 (.ZN( u1_u5_u0_n171 ) , .A( u1_u5_u0_n99 ) );
  OAI211_X1 u1_u5_u0_U51 (.C2( u1_u5_u0_n140 ) , .C1( u1_u5_u0_n161 ) , .A( u1_u5_u0_n169 ) , .B( u1_u5_u0_n98 ) , .ZN( u1_u5_u0_n99 ) );
  INV_X1 u1_u5_u0_U52 (.ZN( u1_u5_u0_n169 ) , .A( u1_u5_u0_n91 ) );
  AOI211_X1 u1_u5_u0_U53 (.C1( u1_u5_u0_n118 ) , .A( u1_u5_u0_n123 ) , .B( u1_u5_u0_n96 ) , .C2( u1_u5_u0_n97 ) , .ZN( u1_u5_u0_n98 ) );
  NOR2_X1 u1_u5_u0_U54 (.A2( u1_u5_X_4 ) , .A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n118 ) );
  NOR2_X1 u1_u5_u0_U55 (.A2( u1_u5_X_1 ) , .ZN( u1_u5_u0_n101 ) , .A1( u1_u5_u0_n163 ) );
  NOR2_X1 u1_u5_u0_U56 (.A2( u1_u5_X_3 ) , .A1( u1_u5_X_6 ) , .ZN( u1_u5_u0_n94 ) );
  NOR2_X1 u1_u5_u0_U57 (.A2( u1_u5_X_6 ) , .ZN( u1_u5_u0_n100 ) , .A1( u1_u5_u0_n162 ) );
  NAND2_X1 u1_u5_u0_U58 (.A2( u1_u5_X_4 ) , .A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n144 ) );
  NOR2_X1 u1_u5_u0_U59 (.A2( u1_u5_X_5 ) , .ZN( u1_u5_u0_n136 ) , .A1( u1_u5_u0_n159 ) );
  NOR2_X1 u1_u5_u0_U6 (.A1( u1_u5_u0_n108 ) , .ZN( u1_u5_u0_n123 ) , .A2( u1_u5_u0_n158 ) );
  NAND2_X1 u1_u5_u0_U60 (.A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n138 ) , .A2( u1_u5_u0_n159 ) );
  AND2_X1 u1_u5_u0_U61 (.A2( u1_u5_X_3 ) , .A1( u1_u5_X_6 ) , .ZN( u1_u5_u0_n102 ) );
  AND2_X1 u1_u5_u0_U62 (.A1( u1_u5_X_6 ) , .A2( u1_u5_u0_n162 ) , .ZN( u1_u5_u0_n93 ) );
  INV_X1 u1_u5_u0_U63 (.A( u1_u5_X_4 ) , .ZN( u1_u5_u0_n159 ) );
  INV_X1 u1_u5_u0_U64 (.A( u1_u5_X_1 ) , .ZN( u1_u5_u0_n164 ) );
  INV_X1 u1_u5_u0_U65 (.A( u1_u5_X_3 ) , .ZN( u1_u5_u0_n162 ) );
  INV_X1 u1_u5_u0_U66 (.A( u1_u5_u0_n126 ) , .ZN( u1_u5_u0_n168 ) );
  AOI211_X1 u1_u5_u0_U67 (.B( u1_u5_u0_n133 ) , .A( u1_u5_u0_n134 ) , .C2( u1_u5_u0_n135 ) , .C1( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n137 ) );
  OR4_X1 u1_u5_u0_U68 (.ZN( u1_out5_17 ) , .A1( u1_u5_u0_n122 ) , .A2( u1_u5_u0_n123 ) , .A4( u1_u5_u0_n124 ) , .A3( u1_u5_u0_n170 ) );
  AOI21_X1 u1_u5_u0_U69 (.B2( u1_u5_u0_n107 ) , .ZN( u1_u5_u0_n124 ) , .B1( u1_u5_u0_n128 ) , .A( u1_u5_u0_n161 ) );
  OAI21_X1 u1_u5_u0_U7 (.B1( u1_u5_u0_n150 ) , .B2( u1_u5_u0_n158 ) , .A( u1_u5_u0_n172 ) , .ZN( u1_u5_u0_n89 ) );
  INV_X1 u1_u5_u0_U70 (.A( u1_u5_u0_n111 ) , .ZN( u1_u5_u0_n170 ) );
  OR4_X1 u1_u5_u0_U71 (.ZN( u1_out5_31 ) , .A4( u1_u5_u0_n155 ) , .A2( u1_u5_u0_n156 ) , .A1( u1_u5_u0_n157 ) , .A3( u1_u5_u0_n173 ) );
  AOI21_X1 u1_u5_u0_U72 (.A( u1_u5_u0_n138 ) , .B2( u1_u5_u0_n139 ) , .B1( u1_u5_u0_n140 ) , .ZN( u1_u5_u0_n157 ) );
  AOI21_X1 u1_u5_u0_U73 (.B2( u1_u5_u0_n141 ) , .B1( u1_u5_u0_n142 ) , .ZN( u1_u5_u0_n156 ) , .A( u1_u5_u0_n161 ) );
  INV_X1 u1_u5_u0_U74 (.ZN( u1_u5_u0_n174 ) , .A( u1_u5_u0_n89 ) );
  AOI211_X1 u1_u5_u0_U75 (.B( u1_u5_u0_n104 ) , .A( u1_u5_u0_n105 ) , .ZN( u1_u5_u0_n106 ) , .C2( u1_u5_u0_n113 ) , .C1( u1_u5_u0_n160 ) );
  OAI221_X1 u1_u5_u0_U76 (.C1( u1_u5_u0_n121 ) , .ZN( u1_u5_u0_n122 ) , .B2( u1_u5_u0_n127 ) , .A( u1_u5_u0_n143 ) , .B1( u1_u5_u0_n144 ) , .C2( u1_u5_u0_n147 ) );
  AOI21_X1 u1_u5_u0_U77 (.B1( u1_u5_u0_n132 ) , .ZN( u1_u5_u0_n133 ) , .A( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n166 ) );
  OAI22_X1 u1_u5_u0_U78 (.ZN( u1_u5_u0_n105 ) , .A2( u1_u5_u0_n132 ) , .B1( u1_u5_u0_n146 ) , .A1( u1_u5_u0_n147 ) , .B2( u1_u5_u0_n161 ) );
  NAND2_X1 u1_u5_u0_U79 (.ZN( u1_u5_u0_n110 ) , .A2( u1_u5_u0_n132 ) , .A1( u1_u5_u0_n145 ) );
  AND2_X1 u1_u5_u0_U8 (.A1( u1_u5_u0_n114 ) , .A2( u1_u5_u0_n121 ) , .ZN( u1_u5_u0_n146 ) );
  INV_X1 u1_u5_u0_U80 (.A( u1_u5_u0_n119 ) , .ZN( u1_u5_u0_n167 ) );
  NAND2_X1 u1_u5_u0_U81 (.ZN( u1_u5_u0_n148 ) , .A1( u1_u5_u0_n93 ) , .A2( u1_u5_u0_n95 ) );
  NAND2_X1 u1_u5_u0_U82 (.A1( u1_u5_u0_n100 ) , .ZN( u1_u5_u0_n129 ) , .A2( u1_u5_u0_n95 ) );
  NAND2_X1 u1_u5_u0_U83 (.A1( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n128 ) , .A2( u1_u5_u0_n95 ) );
  NOR2_X1 u1_u5_u0_U84 (.A2( u1_u5_X_1 ) , .A1( u1_u5_X_2 ) , .ZN( u1_u5_u0_n92 ) );
  NAND2_X1 u1_u5_u0_U85 (.ZN( u1_u5_u0_n142 ) , .A1( u1_u5_u0_n94 ) , .A2( u1_u5_u0_n95 ) );
  NOR2_X1 u1_u5_u0_U86 (.A2( u1_u5_X_2 ) , .ZN( u1_u5_u0_n103 ) , .A1( u1_u5_u0_n164 ) );
  INV_X1 u1_u5_u0_U87 (.A( u1_u5_X_2 ) , .ZN( u1_u5_u0_n163 ) );
  NAND3_X1 u1_u5_u0_U88 (.ZN( u1_out5_23 ) , .A3( u1_u5_u0_n137 ) , .A1( u1_u5_u0_n168 ) , .A2( u1_u5_u0_n171 ) );
  NAND3_X1 u1_u5_u0_U89 (.A3( u1_u5_u0_n127 ) , .A2( u1_u5_u0_n128 ) , .ZN( u1_u5_u0_n135 ) , .A1( u1_u5_u0_n150 ) );
  AND2_X1 u1_u5_u0_U9 (.A1( u1_u5_u0_n131 ) , .ZN( u1_u5_u0_n141 ) , .A2( u1_u5_u0_n150 ) );
  NAND3_X1 u1_u5_u0_U90 (.ZN( u1_u5_u0_n117 ) , .A3( u1_u5_u0_n132 ) , .A2( u1_u5_u0_n139 ) , .A1( u1_u5_u0_n148 ) );
  NAND3_X1 u1_u5_u0_U91 (.ZN( u1_u5_u0_n109 ) , .A2( u1_u5_u0_n114 ) , .A3( u1_u5_u0_n140 ) , .A1( u1_u5_u0_n149 ) );
  NAND3_X1 u1_u5_u0_U92 (.ZN( u1_out5_9 ) , .A3( u1_u5_u0_n106 ) , .A2( u1_u5_u0_n171 ) , .A1( u1_u5_u0_n174 ) );
  NAND3_X1 u1_u5_u0_U93 (.A2( u1_u5_u0_n128 ) , .A1( u1_u5_u0_n132 ) , .A3( u1_u5_u0_n146 ) , .ZN( u1_u5_u0_n97 ) );
  OAI22_X1 u1_u5_u2_U10 (.ZN( u1_u5_u2_n109 ) , .A2( u1_u5_u2_n113 ) , .B2( u1_u5_u2_n133 ) , .B1( u1_u5_u2_n167 ) , .A1( u1_u5_u2_n168 ) );
  NAND3_X1 u1_u5_u2_U100 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n104 ) , .A3( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n98 ) );
  OAI22_X1 u1_u5_u2_U11 (.B1( u1_u5_u2_n151 ) , .A2( u1_u5_u2_n152 ) , .A1( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n160 ) , .B2( u1_u5_u2_n168 ) );
  NOR3_X1 u1_u5_u2_U12 (.A1( u1_u5_u2_n150 ) , .ZN( u1_u5_u2_n151 ) , .A3( u1_u5_u2_n175 ) , .A2( u1_u5_u2_n188 ) );
  AOI21_X1 u1_u5_u2_U13 (.ZN( u1_u5_u2_n144 ) , .B2( u1_u5_u2_n155 ) , .A( u1_u5_u2_n172 ) , .B1( u1_u5_u2_n185 ) );
  AOI21_X1 u1_u5_u2_U14 (.B2( u1_u5_u2_n143 ) , .ZN( u1_u5_u2_n145 ) , .B1( u1_u5_u2_n152 ) , .A( u1_u5_u2_n171 ) );
  AOI21_X1 u1_u5_u2_U15 (.B2( u1_u5_u2_n120 ) , .B1( u1_u5_u2_n121 ) , .ZN( u1_u5_u2_n126 ) , .A( u1_u5_u2_n167 ) );
  INV_X1 u1_u5_u2_U16 (.A( u1_u5_u2_n156 ) , .ZN( u1_u5_u2_n171 ) );
  INV_X1 u1_u5_u2_U17 (.A( u1_u5_u2_n120 ) , .ZN( u1_u5_u2_n188 ) );
  NAND2_X1 u1_u5_u2_U18 (.A2( u1_u5_u2_n122 ) , .ZN( u1_u5_u2_n150 ) , .A1( u1_u5_u2_n152 ) );
  INV_X1 u1_u5_u2_U19 (.A( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n170 ) );
  INV_X1 u1_u5_u2_U20 (.A( u1_u5_u2_n137 ) , .ZN( u1_u5_u2_n173 ) );
  NAND2_X1 u1_u5_u2_U21 (.A1( u1_u5_u2_n132 ) , .A2( u1_u5_u2_n139 ) , .ZN( u1_u5_u2_n157 ) );
  INV_X1 u1_u5_u2_U22 (.A( u1_u5_u2_n113 ) , .ZN( u1_u5_u2_n178 ) );
  INV_X1 u1_u5_u2_U23 (.A( u1_u5_u2_n139 ) , .ZN( u1_u5_u2_n175 ) );
  INV_X1 u1_u5_u2_U24 (.A( u1_u5_u2_n155 ) , .ZN( u1_u5_u2_n181 ) );
  INV_X1 u1_u5_u2_U25 (.A( u1_u5_u2_n119 ) , .ZN( u1_u5_u2_n177 ) );
  INV_X1 u1_u5_u2_U26 (.A( u1_u5_u2_n116 ) , .ZN( u1_u5_u2_n180 ) );
  INV_X1 u1_u5_u2_U27 (.A( u1_u5_u2_n131 ) , .ZN( u1_u5_u2_n179 ) );
  INV_X1 u1_u5_u2_U28 (.A( u1_u5_u2_n154 ) , .ZN( u1_u5_u2_n176 ) );
  NAND2_X1 u1_u5_u2_U29 (.A2( u1_u5_u2_n116 ) , .A1( u1_u5_u2_n117 ) , .ZN( u1_u5_u2_n118 ) );
  NOR2_X1 u1_u5_u2_U3 (.ZN( u1_u5_u2_n121 ) , .A2( u1_u5_u2_n177 ) , .A1( u1_u5_u2_n180 ) );
  INV_X1 u1_u5_u2_U30 (.A( u1_u5_u2_n132 ) , .ZN( u1_u5_u2_n182 ) );
  INV_X1 u1_u5_u2_U31 (.A( u1_u5_u2_n158 ) , .ZN( u1_u5_u2_n183 ) );
  OAI21_X1 u1_u5_u2_U32 (.A( u1_u5_u2_n156 ) , .B1( u1_u5_u2_n157 ) , .ZN( u1_u5_u2_n158 ) , .B2( u1_u5_u2_n179 ) );
  NOR2_X1 u1_u5_u2_U33 (.ZN( u1_u5_u2_n156 ) , .A1( u1_u5_u2_n166 ) , .A2( u1_u5_u2_n169 ) );
  NOR2_X1 u1_u5_u2_U34 (.A2( u1_u5_u2_n114 ) , .ZN( u1_u5_u2_n137 ) , .A1( u1_u5_u2_n140 ) );
  NOR2_X1 u1_u5_u2_U35 (.A2( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n153 ) , .A1( u1_u5_u2_n156 ) );
  AOI211_X1 u1_u5_u2_U36 (.ZN( u1_u5_u2_n130 ) , .C1( u1_u5_u2_n138 ) , .C2( u1_u5_u2_n179 ) , .B( u1_u5_u2_n96 ) , .A( u1_u5_u2_n97 ) );
  OAI22_X1 u1_u5_u2_U37 (.B1( u1_u5_u2_n133 ) , .A2( u1_u5_u2_n137 ) , .A1( u1_u5_u2_n152 ) , .B2( u1_u5_u2_n168 ) , .ZN( u1_u5_u2_n97 ) );
  OAI221_X1 u1_u5_u2_U38 (.B1( u1_u5_u2_n113 ) , .C1( u1_u5_u2_n132 ) , .A( u1_u5_u2_n149 ) , .B2( u1_u5_u2_n171 ) , .C2( u1_u5_u2_n172 ) , .ZN( u1_u5_u2_n96 ) );
  OAI221_X1 u1_u5_u2_U39 (.A( u1_u5_u2_n115 ) , .C2( u1_u5_u2_n123 ) , .B2( u1_u5_u2_n143 ) , .B1( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n163 ) , .C1( u1_u5_u2_n168 ) );
  INV_X1 u1_u5_u2_U4 (.A( u1_u5_u2_n134 ) , .ZN( u1_u5_u2_n185 ) );
  OAI21_X1 u1_u5_u2_U40 (.A( u1_u5_u2_n114 ) , .ZN( u1_u5_u2_n115 ) , .B1( u1_u5_u2_n176 ) , .B2( u1_u5_u2_n178 ) );
  OAI221_X1 u1_u5_u2_U41 (.A( u1_u5_u2_n135 ) , .B2( u1_u5_u2_n136 ) , .B1( u1_u5_u2_n137 ) , .ZN( u1_u5_u2_n162 ) , .C2( u1_u5_u2_n167 ) , .C1( u1_u5_u2_n185 ) );
  AND3_X1 u1_u5_u2_U42 (.A3( u1_u5_u2_n131 ) , .A2( u1_u5_u2_n132 ) , .A1( u1_u5_u2_n133 ) , .ZN( u1_u5_u2_n136 ) );
  AOI22_X1 u1_u5_u2_U43 (.ZN( u1_u5_u2_n135 ) , .B1( u1_u5_u2_n140 ) , .A1( u1_u5_u2_n156 ) , .B2( u1_u5_u2_n180 ) , .A2( u1_u5_u2_n188 ) );
  AOI21_X1 u1_u5_u2_U44 (.ZN( u1_u5_u2_n149 ) , .B1( u1_u5_u2_n173 ) , .B2( u1_u5_u2_n188 ) , .A( u1_u5_u2_n95 ) );
  AND3_X1 u1_u5_u2_U45 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n104 ) , .A3( u1_u5_u2_n156 ) , .ZN( u1_u5_u2_n95 ) );
  OAI21_X1 u1_u5_u2_U46 (.A( u1_u5_u2_n101 ) , .B2( u1_u5_u2_n121 ) , .B1( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n164 ) );
  NAND2_X1 u1_u5_u2_U47 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n107 ) , .ZN( u1_u5_u2_n155 ) );
  NAND2_X1 u1_u5_u2_U48 (.A2( u1_u5_u2_n105 ) , .A1( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n143 ) );
  NAND2_X1 u1_u5_u2_U49 (.A1( u1_u5_u2_n104 ) , .A2( u1_u5_u2_n106 ) , .ZN( u1_u5_u2_n152 ) );
  INV_X1 u1_u5_u2_U5 (.A( u1_u5_u2_n150 ) , .ZN( u1_u5_u2_n184 ) );
  NAND2_X1 u1_u5_u2_U50 (.A1( u1_u5_u2_n100 ) , .A2( u1_u5_u2_n105 ) , .ZN( u1_u5_u2_n132 ) );
  INV_X1 u1_u5_u2_U51 (.A( u1_u5_u2_n140 ) , .ZN( u1_u5_u2_n168 ) );
  INV_X1 u1_u5_u2_U52 (.A( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n167 ) );
  OAI21_X1 u1_u5_u2_U53 (.A( u1_u5_u2_n141 ) , .B2( u1_u5_u2_n142 ) , .ZN( u1_u5_u2_n146 ) , .B1( u1_u5_u2_n153 ) );
  OAI21_X1 u1_u5_u2_U54 (.A( u1_u5_u2_n140 ) , .ZN( u1_u5_u2_n141 ) , .B1( u1_u5_u2_n176 ) , .B2( u1_u5_u2_n177 ) );
  NOR3_X1 u1_u5_u2_U55 (.ZN( u1_u5_u2_n142 ) , .A3( u1_u5_u2_n175 ) , .A2( u1_u5_u2_n178 ) , .A1( u1_u5_u2_n181 ) );
  INV_X1 u1_u5_u2_U56 (.ZN( u1_u5_u2_n187 ) , .A( u1_u5_u2_n99 ) );
  OAI21_X1 u1_u5_u2_U57 (.B1( u1_u5_u2_n137 ) , .B2( u1_u5_u2_n143 ) , .A( u1_u5_u2_n98 ) , .ZN( u1_u5_u2_n99 ) );
  NAND2_X1 u1_u5_u2_U58 (.A1( u1_u5_u2_n102 ) , .A2( u1_u5_u2_n106 ) , .ZN( u1_u5_u2_n113 ) );
  NAND2_X1 u1_u5_u2_U59 (.A1( u1_u5_u2_n106 ) , .A2( u1_u5_u2_n107 ) , .ZN( u1_u5_u2_n131 ) );
  NOR4_X1 u1_u5_u2_U6 (.A4( u1_u5_u2_n124 ) , .A3( u1_u5_u2_n125 ) , .A2( u1_u5_u2_n126 ) , .A1( u1_u5_u2_n127 ) , .ZN( u1_u5_u2_n128 ) );
  NAND2_X1 u1_u5_u2_U60 (.A1( u1_u5_u2_n103 ) , .A2( u1_u5_u2_n107 ) , .ZN( u1_u5_u2_n139 ) );
  NAND2_X1 u1_u5_u2_U61 (.A1( u1_u5_u2_n103 ) , .A2( u1_u5_u2_n105 ) , .ZN( u1_u5_u2_n133 ) );
  NAND2_X1 u1_u5_u2_U62 (.A1( u1_u5_u2_n102 ) , .A2( u1_u5_u2_n103 ) , .ZN( u1_u5_u2_n154 ) );
  NAND2_X1 u1_u5_u2_U63 (.A2( u1_u5_u2_n103 ) , .A1( u1_u5_u2_n104 ) , .ZN( u1_u5_u2_n119 ) );
  NAND2_X1 u1_u5_u2_U64 (.A2( u1_u5_u2_n107 ) , .A1( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n123 ) );
  NAND2_X1 u1_u5_u2_U65 (.A1( u1_u5_u2_n104 ) , .A2( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n122 ) );
  INV_X1 u1_u5_u2_U66 (.A( u1_u5_u2_n114 ) , .ZN( u1_u5_u2_n172 ) );
  NAND2_X1 u1_u5_u2_U67 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n102 ) , .ZN( u1_u5_u2_n116 ) );
  NAND2_X1 u1_u5_u2_U68 (.A1( u1_u5_u2_n102 ) , .A2( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n120 ) );
  NAND2_X1 u1_u5_u2_U69 (.A2( u1_u5_u2_n105 ) , .A1( u1_u5_u2_n106 ) , .ZN( u1_u5_u2_n117 ) );
  AOI21_X1 u1_u5_u2_U7 (.B2( u1_u5_u2_n119 ) , .ZN( u1_u5_u2_n127 ) , .A( u1_u5_u2_n137 ) , .B1( u1_u5_u2_n155 ) );
  NOR2_X1 u1_u5_u2_U70 (.A2( u1_u5_X_16 ) , .ZN( u1_u5_u2_n140 ) , .A1( u1_u5_u2_n166 ) );
  NOR2_X1 u1_u5_u2_U71 (.A2( u1_u5_X_13 ) , .A1( u1_u5_X_14 ) , .ZN( u1_u5_u2_n100 ) );
  NOR2_X1 u1_u5_u2_U72 (.A2( u1_u5_X_16 ) , .A1( u1_u5_X_17 ) , .ZN( u1_u5_u2_n138 ) );
  NOR2_X1 u1_u5_u2_U73 (.A2( u1_u5_X_15 ) , .A1( u1_u5_X_18 ) , .ZN( u1_u5_u2_n104 ) );
  NOR2_X1 u1_u5_u2_U74 (.A2( u1_u5_X_14 ) , .ZN( u1_u5_u2_n103 ) , .A1( u1_u5_u2_n174 ) );
  NOR2_X1 u1_u5_u2_U75 (.A2( u1_u5_X_15 ) , .ZN( u1_u5_u2_n102 ) , .A1( u1_u5_u2_n165 ) );
  NOR2_X1 u1_u5_u2_U76 (.A2( u1_u5_X_17 ) , .ZN( u1_u5_u2_n114 ) , .A1( u1_u5_u2_n169 ) );
  AND2_X1 u1_u5_u2_U77 (.A1( u1_u5_X_15 ) , .ZN( u1_u5_u2_n105 ) , .A2( u1_u5_u2_n165 ) );
  AND2_X1 u1_u5_u2_U78 (.A2( u1_u5_X_15 ) , .A1( u1_u5_X_18 ) , .ZN( u1_u5_u2_n107 ) );
  AND2_X1 u1_u5_u2_U79 (.A1( u1_u5_X_14 ) , .ZN( u1_u5_u2_n106 ) , .A2( u1_u5_u2_n174 ) );
  AOI21_X1 u1_u5_u2_U8 (.ZN( u1_u5_u2_n124 ) , .B1( u1_u5_u2_n131 ) , .B2( u1_u5_u2_n143 ) , .A( u1_u5_u2_n172 ) );
  AND2_X1 u1_u5_u2_U80 (.A1( u1_u5_X_13 ) , .A2( u1_u5_X_14 ) , .ZN( u1_u5_u2_n108 ) );
  INV_X1 u1_u5_u2_U81 (.A( u1_u5_X_16 ) , .ZN( u1_u5_u2_n169 ) );
  INV_X1 u1_u5_u2_U82 (.A( u1_u5_X_17 ) , .ZN( u1_u5_u2_n166 ) );
  INV_X1 u1_u5_u2_U83 (.A( u1_u5_X_13 ) , .ZN( u1_u5_u2_n174 ) );
  INV_X1 u1_u5_u2_U84 (.A( u1_u5_X_18 ) , .ZN( u1_u5_u2_n165 ) );
  NAND4_X1 u1_u5_u2_U85 (.ZN( u1_out5_30 ) , .A4( u1_u5_u2_n147 ) , .A3( u1_u5_u2_n148 ) , .A2( u1_u5_u2_n149 ) , .A1( u1_u5_u2_n187 ) );
  NOR3_X1 u1_u5_u2_U86 (.A3( u1_u5_u2_n144 ) , .A2( u1_u5_u2_n145 ) , .A1( u1_u5_u2_n146 ) , .ZN( u1_u5_u2_n147 ) );
  AOI21_X1 u1_u5_u2_U87 (.B2( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n148 ) , .A( u1_u5_u2_n162 ) , .B1( u1_u5_u2_n182 ) );
  NAND4_X1 u1_u5_u2_U88 (.ZN( u1_out5_24 ) , .A4( u1_u5_u2_n111 ) , .A3( u1_u5_u2_n112 ) , .A1( u1_u5_u2_n130 ) , .A2( u1_u5_u2_n187 ) );
  AOI221_X1 u1_u5_u2_U89 (.A( u1_u5_u2_n109 ) , .B1( u1_u5_u2_n110 ) , .ZN( u1_u5_u2_n111 ) , .C1( u1_u5_u2_n134 ) , .C2( u1_u5_u2_n170 ) , .B2( u1_u5_u2_n173 ) );
  AOI21_X1 u1_u5_u2_U9 (.B2( u1_u5_u2_n123 ) , .ZN( u1_u5_u2_n125 ) , .A( u1_u5_u2_n171 ) , .B1( u1_u5_u2_n184 ) );
  AOI21_X1 u1_u5_u2_U90 (.ZN( u1_u5_u2_n112 ) , .B2( u1_u5_u2_n156 ) , .A( u1_u5_u2_n164 ) , .B1( u1_u5_u2_n181 ) );
  NAND4_X1 u1_u5_u2_U91 (.ZN( u1_out5_16 ) , .A4( u1_u5_u2_n128 ) , .A3( u1_u5_u2_n129 ) , .A1( u1_u5_u2_n130 ) , .A2( u1_u5_u2_n186 ) );
  AOI22_X1 u1_u5_u2_U92 (.A2( u1_u5_u2_n118 ) , .ZN( u1_u5_u2_n129 ) , .A1( u1_u5_u2_n140 ) , .B1( u1_u5_u2_n157 ) , .B2( u1_u5_u2_n170 ) );
  INV_X1 u1_u5_u2_U93 (.A( u1_u5_u2_n163 ) , .ZN( u1_u5_u2_n186 ) );
  OR4_X1 u1_u5_u2_U94 (.ZN( u1_out5_6 ) , .A4( u1_u5_u2_n161 ) , .A3( u1_u5_u2_n162 ) , .A2( u1_u5_u2_n163 ) , .A1( u1_u5_u2_n164 ) );
  OR3_X1 u1_u5_u2_U95 (.A2( u1_u5_u2_n159 ) , .A1( u1_u5_u2_n160 ) , .ZN( u1_u5_u2_n161 ) , .A3( u1_u5_u2_n183 ) );
  AOI21_X1 u1_u5_u2_U96 (.B2( u1_u5_u2_n154 ) , .B1( u1_u5_u2_n155 ) , .ZN( u1_u5_u2_n159 ) , .A( u1_u5_u2_n167 ) );
  NAND3_X1 u1_u5_u2_U97 (.A2( u1_u5_u2_n117 ) , .A1( u1_u5_u2_n122 ) , .A3( u1_u5_u2_n123 ) , .ZN( u1_u5_u2_n134 ) );
  NAND3_X1 u1_u5_u2_U98 (.ZN( u1_u5_u2_n110 ) , .A2( u1_u5_u2_n131 ) , .A3( u1_u5_u2_n139 ) , .A1( u1_u5_u2_n154 ) );
  NAND3_X1 u1_u5_u2_U99 (.A2( u1_u5_u2_n100 ) , .ZN( u1_u5_u2_n101 ) , .A1( u1_u5_u2_n104 ) , .A3( u1_u5_u2_n114 ) );
  OAI22_X1 u1_u5_u3_U10 (.B1( u1_u5_u3_n113 ) , .A2( u1_u5_u3_n135 ) , .A1( u1_u5_u3_n150 ) , .B2( u1_u5_u3_n164 ) , .ZN( u1_u5_u3_n98 ) );
  OAI211_X1 u1_u5_u3_U11 (.B( u1_u5_u3_n106 ) , .ZN( u1_u5_u3_n119 ) , .C2( u1_u5_u3_n128 ) , .C1( u1_u5_u3_n167 ) , .A( u1_u5_u3_n181 ) );
  AOI221_X1 u1_u5_u3_U12 (.C1( u1_u5_u3_n105 ) , .ZN( u1_u5_u3_n106 ) , .A( u1_u5_u3_n131 ) , .B2( u1_u5_u3_n132 ) , .C2( u1_u5_u3_n133 ) , .B1( u1_u5_u3_n169 ) );
  INV_X1 u1_u5_u3_U13 (.ZN( u1_u5_u3_n181 ) , .A( u1_u5_u3_n98 ) );
  NAND2_X1 u1_u5_u3_U14 (.ZN( u1_u5_u3_n105 ) , .A2( u1_u5_u3_n130 ) , .A1( u1_u5_u3_n155 ) );
  AOI22_X1 u1_u5_u3_U15 (.B1( u1_u5_u3_n115 ) , .A2( u1_u5_u3_n116 ) , .ZN( u1_u5_u3_n123 ) , .B2( u1_u5_u3_n133 ) , .A1( u1_u5_u3_n169 ) );
  NAND2_X1 u1_u5_u3_U16 (.ZN( u1_u5_u3_n116 ) , .A2( u1_u5_u3_n151 ) , .A1( u1_u5_u3_n182 ) );
  NOR2_X1 u1_u5_u3_U17 (.ZN( u1_u5_u3_n126 ) , .A2( u1_u5_u3_n150 ) , .A1( u1_u5_u3_n164 ) );
  AOI21_X1 u1_u5_u3_U18 (.ZN( u1_u5_u3_n112 ) , .B2( u1_u5_u3_n146 ) , .B1( u1_u5_u3_n155 ) , .A( u1_u5_u3_n167 ) );
  NAND2_X1 u1_u5_u3_U19 (.A1( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n142 ) , .A2( u1_u5_u3_n164 ) );
  NAND2_X1 u1_u5_u3_U20 (.ZN( u1_u5_u3_n132 ) , .A2( u1_u5_u3_n152 ) , .A1( u1_u5_u3_n156 ) );
  AND2_X1 u1_u5_u3_U21 (.A2( u1_u5_u3_n113 ) , .A1( u1_u5_u3_n114 ) , .ZN( u1_u5_u3_n151 ) );
  INV_X1 u1_u5_u3_U22 (.A( u1_u5_u3_n133 ) , .ZN( u1_u5_u3_n165 ) );
  INV_X1 u1_u5_u3_U23 (.A( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n170 ) );
  NAND2_X1 u1_u5_u3_U24 (.A1( u1_u5_u3_n107 ) , .A2( u1_u5_u3_n108 ) , .ZN( u1_u5_u3_n140 ) );
  NAND2_X1 u1_u5_u3_U25 (.ZN( u1_u5_u3_n117 ) , .A1( u1_u5_u3_n124 ) , .A2( u1_u5_u3_n148 ) );
  NAND2_X1 u1_u5_u3_U26 (.ZN( u1_u5_u3_n143 ) , .A1( u1_u5_u3_n165 ) , .A2( u1_u5_u3_n167 ) );
  INV_X1 u1_u5_u3_U27 (.A( u1_u5_u3_n130 ) , .ZN( u1_u5_u3_n177 ) );
  INV_X1 u1_u5_u3_U28 (.A( u1_u5_u3_n128 ) , .ZN( u1_u5_u3_n176 ) );
  INV_X1 u1_u5_u3_U29 (.A( u1_u5_u3_n155 ) , .ZN( u1_u5_u3_n174 ) );
  INV_X1 u1_u5_u3_U3 (.A( u1_u5_u3_n129 ) , .ZN( u1_u5_u3_n183 ) );
  INV_X1 u1_u5_u3_U30 (.A( u1_u5_u3_n139 ) , .ZN( u1_u5_u3_n185 ) );
  NOR2_X1 u1_u5_u3_U31 (.ZN( u1_u5_u3_n135 ) , .A2( u1_u5_u3_n141 ) , .A1( u1_u5_u3_n169 ) );
  OAI222_X1 u1_u5_u3_U32 (.C2( u1_u5_u3_n107 ) , .A2( u1_u5_u3_n108 ) , .B1( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n138 ) , .B2( u1_u5_u3_n146 ) , .C1( u1_u5_u3_n154 ) , .A1( u1_u5_u3_n164 ) );
  NOR4_X1 u1_u5_u3_U33 (.A4( u1_u5_u3_n157 ) , .A3( u1_u5_u3_n158 ) , .A2( u1_u5_u3_n159 ) , .A1( u1_u5_u3_n160 ) , .ZN( u1_u5_u3_n161 ) );
  AOI21_X1 u1_u5_u3_U34 (.B2( u1_u5_u3_n152 ) , .B1( u1_u5_u3_n153 ) , .ZN( u1_u5_u3_n158 ) , .A( u1_u5_u3_n164 ) );
  AOI21_X1 u1_u5_u3_U35 (.A( u1_u5_u3_n154 ) , .B2( u1_u5_u3_n155 ) , .B1( u1_u5_u3_n156 ) , .ZN( u1_u5_u3_n157 ) );
  AOI21_X1 u1_u5_u3_U36 (.A( u1_u5_u3_n149 ) , .B2( u1_u5_u3_n150 ) , .B1( u1_u5_u3_n151 ) , .ZN( u1_u5_u3_n159 ) );
  AOI211_X1 u1_u5_u3_U37 (.ZN( u1_u5_u3_n109 ) , .A( u1_u5_u3_n119 ) , .C2( u1_u5_u3_n129 ) , .B( u1_u5_u3_n138 ) , .C1( u1_u5_u3_n141 ) );
  AOI211_X1 u1_u5_u3_U38 (.B( u1_u5_u3_n119 ) , .A( u1_u5_u3_n120 ) , .C2( u1_u5_u3_n121 ) , .ZN( u1_u5_u3_n122 ) , .C1( u1_u5_u3_n179 ) );
  INV_X1 u1_u5_u3_U39 (.A( u1_u5_u3_n156 ) , .ZN( u1_u5_u3_n179 ) );
  INV_X1 u1_u5_u3_U4 (.A( u1_u5_u3_n140 ) , .ZN( u1_u5_u3_n182 ) );
  OAI22_X1 u1_u5_u3_U40 (.B1( u1_u5_u3_n118 ) , .ZN( u1_u5_u3_n120 ) , .A1( u1_u5_u3_n135 ) , .B2( u1_u5_u3_n154 ) , .A2( u1_u5_u3_n178 ) );
  AND3_X1 u1_u5_u3_U41 (.ZN( u1_u5_u3_n118 ) , .A2( u1_u5_u3_n124 ) , .A1( u1_u5_u3_n144 ) , .A3( u1_u5_u3_n152 ) );
  INV_X1 u1_u5_u3_U42 (.A( u1_u5_u3_n121 ) , .ZN( u1_u5_u3_n164 ) );
  NAND2_X1 u1_u5_u3_U43 (.ZN( u1_u5_u3_n133 ) , .A1( u1_u5_u3_n154 ) , .A2( u1_u5_u3_n164 ) );
  OAI211_X1 u1_u5_u3_U44 (.B( u1_u5_u3_n127 ) , .ZN( u1_u5_u3_n139 ) , .C1( u1_u5_u3_n150 ) , .C2( u1_u5_u3_n154 ) , .A( u1_u5_u3_n184 ) );
  INV_X1 u1_u5_u3_U45 (.A( u1_u5_u3_n125 ) , .ZN( u1_u5_u3_n184 ) );
  AOI221_X1 u1_u5_u3_U46 (.A( u1_u5_u3_n126 ) , .ZN( u1_u5_u3_n127 ) , .C2( u1_u5_u3_n132 ) , .C1( u1_u5_u3_n169 ) , .B2( u1_u5_u3_n170 ) , .B1( u1_u5_u3_n174 ) );
  OAI22_X1 u1_u5_u3_U47 (.A1( u1_u5_u3_n124 ) , .ZN( u1_u5_u3_n125 ) , .B2( u1_u5_u3_n145 ) , .A2( u1_u5_u3_n165 ) , .B1( u1_u5_u3_n167 ) );
  NOR2_X1 u1_u5_u3_U48 (.A1( u1_u5_u3_n113 ) , .ZN( u1_u5_u3_n131 ) , .A2( u1_u5_u3_n154 ) );
  NAND2_X1 u1_u5_u3_U49 (.A1( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n150 ) , .A2( u1_u5_u3_n99 ) );
  INV_X1 u1_u5_u3_U5 (.A( u1_u5_u3_n117 ) , .ZN( u1_u5_u3_n178 ) );
  NAND2_X1 u1_u5_u3_U50 (.A2( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n155 ) , .A1( u1_u5_u3_n97 ) );
  INV_X1 u1_u5_u3_U51 (.A( u1_u5_u3_n141 ) , .ZN( u1_u5_u3_n167 ) );
  AOI21_X1 u1_u5_u3_U52 (.B2( u1_u5_u3_n114 ) , .B1( u1_u5_u3_n146 ) , .A( u1_u5_u3_n154 ) , .ZN( u1_u5_u3_n94 ) );
  AOI21_X1 u1_u5_u3_U53 (.ZN( u1_u5_u3_n110 ) , .B2( u1_u5_u3_n142 ) , .B1( u1_u5_u3_n186 ) , .A( u1_u5_u3_n95 ) );
  INV_X1 u1_u5_u3_U54 (.A( u1_u5_u3_n145 ) , .ZN( u1_u5_u3_n186 ) );
  AOI21_X1 u1_u5_u3_U55 (.B1( u1_u5_u3_n124 ) , .A( u1_u5_u3_n149 ) , .B2( u1_u5_u3_n155 ) , .ZN( u1_u5_u3_n95 ) );
  INV_X1 u1_u5_u3_U56 (.A( u1_u5_u3_n149 ) , .ZN( u1_u5_u3_n169 ) );
  NAND2_X1 u1_u5_u3_U57 (.ZN( u1_u5_u3_n124 ) , .A1( u1_u5_u3_n96 ) , .A2( u1_u5_u3_n97 ) );
  NAND2_X1 u1_u5_u3_U58 (.A2( u1_u5_u3_n100 ) , .ZN( u1_u5_u3_n146 ) , .A1( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U59 (.A1( u1_u5_u3_n101 ) , .ZN( u1_u5_u3_n145 ) , .A2( u1_u5_u3_n99 ) );
  AOI221_X1 u1_u5_u3_U6 (.A( u1_u5_u3_n131 ) , .C2( u1_u5_u3_n132 ) , .C1( u1_u5_u3_n133 ) , .ZN( u1_u5_u3_n134 ) , .B1( u1_u5_u3_n143 ) , .B2( u1_u5_u3_n177 ) );
  NAND2_X1 u1_u5_u3_U60 (.A1( u1_u5_u3_n100 ) , .ZN( u1_u5_u3_n156 ) , .A2( u1_u5_u3_n99 ) );
  NAND2_X1 u1_u5_u3_U61 (.A2( u1_u5_u3_n101 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n148 ) );
  NAND2_X1 u1_u5_u3_U62 (.A1( u1_u5_u3_n100 ) , .A2( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n128 ) );
  NAND2_X1 u1_u5_u3_U63 (.A2( u1_u5_u3_n101 ) , .A1( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n152 ) );
  NAND2_X1 u1_u5_u3_U64 (.A2( u1_u5_u3_n101 ) , .ZN( u1_u5_u3_n114 ) , .A1( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U65 (.ZN( u1_u5_u3_n107 ) , .A1( u1_u5_u3_n97 ) , .A2( u1_u5_u3_n99 ) );
  NAND2_X1 u1_u5_u3_U66 (.A2( u1_u5_u3_n100 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n113 ) );
  NAND2_X1 u1_u5_u3_U67 (.A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n153 ) , .A2( u1_u5_u3_n97 ) );
  NAND2_X1 u1_u5_u3_U68 (.A2( u1_u5_u3_n103 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n130 ) );
  NAND2_X1 u1_u5_u3_U69 (.A2( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n144 ) , .A1( u1_u5_u3_n96 ) );
  OAI22_X1 u1_u5_u3_U7 (.B2( u1_u5_u3_n147 ) , .A2( u1_u5_u3_n148 ) , .ZN( u1_u5_u3_n160 ) , .B1( u1_u5_u3_n165 ) , .A1( u1_u5_u3_n168 ) );
  NAND2_X1 u1_u5_u3_U70 (.A1( u1_u5_u3_n102 ) , .A2( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n108 ) );
  NOR2_X1 u1_u5_u3_U71 (.A2( u1_u5_X_19 ) , .A1( u1_u5_X_20 ) , .ZN( u1_u5_u3_n99 ) );
  NOR2_X1 u1_u5_u3_U72 (.A2( u1_u5_X_21 ) , .A1( u1_u5_X_24 ) , .ZN( u1_u5_u3_n103 ) );
  NOR2_X1 u1_u5_u3_U73 (.A2( u1_u5_X_24 ) , .A1( u1_u5_u3_n171 ) , .ZN( u1_u5_u3_n97 ) );
  NOR2_X1 u1_u5_u3_U74 (.A2( u1_u5_X_23 ) , .ZN( u1_u5_u3_n141 ) , .A1( u1_u5_u3_n166 ) );
  NOR2_X1 u1_u5_u3_U75 (.A2( u1_u5_X_19 ) , .A1( u1_u5_u3_n172 ) , .ZN( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U76 (.A1( u1_u5_X_22 ) , .A2( u1_u5_X_23 ) , .ZN( u1_u5_u3_n154 ) );
  NAND2_X1 u1_u5_u3_U77 (.A1( u1_u5_X_23 ) , .ZN( u1_u5_u3_n149 ) , .A2( u1_u5_u3_n166 ) );
  NOR2_X1 u1_u5_u3_U78 (.A2( u1_u5_X_22 ) , .A1( u1_u5_X_23 ) , .ZN( u1_u5_u3_n121 ) );
  AND2_X1 u1_u5_u3_U79 (.A1( u1_u5_X_24 ) , .ZN( u1_u5_u3_n101 ) , .A2( u1_u5_u3_n171 ) );
  AND3_X1 u1_u5_u3_U8 (.A3( u1_u5_u3_n144 ) , .A2( u1_u5_u3_n145 ) , .A1( u1_u5_u3_n146 ) , .ZN( u1_u5_u3_n147 ) );
  AND2_X1 u1_u5_u3_U80 (.A1( u1_u5_X_19 ) , .ZN( u1_u5_u3_n102 ) , .A2( u1_u5_u3_n172 ) );
  AND2_X1 u1_u5_u3_U81 (.A1( u1_u5_X_21 ) , .A2( u1_u5_X_24 ) , .ZN( u1_u5_u3_n100 ) );
  AND2_X1 u1_u5_u3_U82 (.A2( u1_u5_X_19 ) , .A1( u1_u5_X_20 ) , .ZN( u1_u5_u3_n104 ) );
  INV_X1 u1_u5_u3_U83 (.A( u1_u5_X_22 ) , .ZN( u1_u5_u3_n166 ) );
  INV_X1 u1_u5_u3_U84 (.A( u1_u5_X_21 ) , .ZN( u1_u5_u3_n171 ) );
  INV_X1 u1_u5_u3_U85 (.A( u1_u5_X_20 ) , .ZN( u1_u5_u3_n172 ) );
  NAND4_X1 u1_u5_u3_U86 (.ZN( u1_out5_26 ) , .A4( u1_u5_u3_n109 ) , .A3( u1_u5_u3_n110 ) , .A2( u1_u5_u3_n111 ) , .A1( u1_u5_u3_n173 ) );
  INV_X1 u1_u5_u3_U87 (.ZN( u1_u5_u3_n173 ) , .A( u1_u5_u3_n94 ) );
  OAI21_X1 u1_u5_u3_U88 (.ZN( u1_u5_u3_n111 ) , .B2( u1_u5_u3_n117 ) , .A( u1_u5_u3_n133 ) , .B1( u1_u5_u3_n176 ) );
  NAND4_X1 u1_u5_u3_U89 (.ZN( u1_out5_20 ) , .A4( u1_u5_u3_n122 ) , .A3( u1_u5_u3_n123 ) , .A1( u1_u5_u3_n175 ) , .A2( u1_u5_u3_n180 ) );
  INV_X1 u1_u5_u3_U9 (.A( u1_u5_u3_n143 ) , .ZN( u1_u5_u3_n168 ) );
  INV_X1 u1_u5_u3_U90 (.A( u1_u5_u3_n126 ) , .ZN( u1_u5_u3_n180 ) );
  INV_X1 u1_u5_u3_U91 (.A( u1_u5_u3_n112 ) , .ZN( u1_u5_u3_n175 ) );
  OR4_X1 u1_u5_u3_U92 (.ZN( u1_out5_10 ) , .A4( u1_u5_u3_n136 ) , .A3( u1_u5_u3_n137 ) , .A1( u1_u5_u3_n138 ) , .A2( u1_u5_u3_n139 ) );
  OAI222_X1 u1_u5_u3_U93 (.C1( u1_u5_u3_n128 ) , .ZN( u1_u5_u3_n137 ) , .B1( u1_u5_u3_n148 ) , .A2( u1_u5_u3_n150 ) , .B2( u1_u5_u3_n154 ) , .C2( u1_u5_u3_n164 ) , .A1( u1_u5_u3_n167 ) );
  OAI221_X1 u1_u5_u3_U94 (.A( u1_u5_u3_n134 ) , .B2( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n136 ) , .C1( u1_u5_u3_n149 ) , .B1( u1_u5_u3_n151 ) , .C2( u1_u5_u3_n183 ) );
  NAND4_X1 u1_u5_u3_U95 (.ZN( u1_out5_1 ) , .A4( u1_u5_u3_n161 ) , .A3( u1_u5_u3_n162 ) , .A2( u1_u5_u3_n163 ) , .A1( u1_u5_u3_n185 ) );
  NAND2_X1 u1_u5_u3_U96 (.ZN( u1_u5_u3_n163 ) , .A2( u1_u5_u3_n170 ) , .A1( u1_u5_u3_n176 ) );
  AOI22_X1 u1_u5_u3_U97 (.B2( u1_u5_u3_n140 ) , .B1( u1_u5_u3_n141 ) , .A2( u1_u5_u3_n142 ) , .ZN( u1_u5_u3_n162 ) , .A1( u1_u5_u3_n177 ) );
  NAND3_X1 u1_u5_u3_U98 (.A1( u1_u5_u3_n114 ) , .ZN( u1_u5_u3_n115 ) , .A2( u1_u5_u3_n145 ) , .A3( u1_u5_u3_n153 ) );
  NAND3_X1 u1_u5_u3_U99 (.ZN( u1_u5_u3_n129 ) , .A2( u1_u5_u3_n144 ) , .A1( u1_u5_u3_n153 ) , .A3( u1_u5_u3_n182 ) );
  OAI22_X1 u1_u5_u4_U10 (.B2( u1_u5_u4_n135 ) , .ZN( u1_u5_u4_n137 ) , .B1( u1_u5_u4_n153 ) , .A1( u1_u5_u4_n155 ) , .A2( u1_u5_u4_n171 ) );
  AND3_X1 u1_u5_u4_U11 (.A2( u1_u5_u4_n134 ) , .ZN( u1_u5_u4_n135 ) , .A3( u1_u5_u4_n145 ) , .A1( u1_u5_u4_n157 ) );
  NAND2_X1 u1_u5_u4_U12 (.ZN( u1_u5_u4_n132 ) , .A2( u1_u5_u4_n170 ) , .A1( u1_u5_u4_n173 ) );
  AOI21_X1 u1_u5_u4_U13 (.B2( u1_u5_u4_n160 ) , .B1( u1_u5_u4_n161 ) , .ZN( u1_u5_u4_n162 ) , .A( u1_u5_u4_n170 ) );
  AOI21_X1 u1_u5_u4_U14 (.ZN( u1_u5_u4_n107 ) , .B2( u1_u5_u4_n143 ) , .A( u1_u5_u4_n174 ) , .B1( u1_u5_u4_n184 ) );
  AOI21_X1 u1_u5_u4_U15 (.B2( u1_u5_u4_n158 ) , .B1( u1_u5_u4_n159 ) , .ZN( u1_u5_u4_n163 ) , .A( u1_u5_u4_n174 ) );
  AOI21_X1 u1_u5_u4_U16 (.A( u1_u5_u4_n153 ) , .B2( u1_u5_u4_n154 ) , .B1( u1_u5_u4_n155 ) , .ZN( u1_u5_u4_n165 ) );
  AOI21_X1 u1_u5_u4_U17 (.A( u1_u5_u4_n156 ) , .B2( u1_u5_u4_n157 ) , .ZN( u1_u5_u4_n164 ) , .B1( u1_u5_u4_n184 ) );
  INV_X1 u1_u5_u4_U18 (.A( u1_u5_u4_n138 ) , .ZN( u1_u5_u4_n170 ) );
  AND2_X1 u1_u5_u4_U19 (.A2( u1_u5_u4_n120 ) , .ZN( u1_u5_u4_n155 ) , .A1( u1_u5_u4_n160 ) );
  INV_X1 u1_u5_u4_U20 (.A( u1_u5_u4_n156 ) , .ZN( u1_u5_u4_n175 ) );
  NAND2_X1 u1_u5_u4_U21 (.A2( u1_u5_u4_n118 ) , .ZN( u1_u5_u4_n131 ) , .A1( u1_u5_u4_n147 ) );
  NAND2_X1 u1_u5_u4_U22 (.A1( u1_u5_u4_n119 ) , .A2( u1_u5_u4_n120 ) , .ZN( u1_u5_u4_n130 ) );
  NAND2_X1 u1_u5_u4_U23 (.ZN( u1_u5_u4_n117 ) , .A2( u1_u5_u4_n118 ) , .A1( u1_u5_u4_n148 ) );
  NAND2_X1 u1_u5_u4_U24 (.ZN( u1_u5_u4_n129 ) , .A1( u1_u5_u4_n134 ) , .A2( u1_u5_u4_n148 ) );
  AND3_X1 u1_u5_u4_U25 (.A1( u1_u5_u4_n119 ) , .A2( u1_u5_u4_n143 ) , .A3( u1_u5_u4_n154 ) , .ZN( u1_u5_u4_n161 ) );
  AND2_X1 u1_u5_u4_U26 (.A1( u1_u5_u4_n145 ) , .A2( u1_u5_u4_n147 ) , .ZN( u1_u5_u4_n159 ) );
  OR3_X1 u1_u5_u4_U27 (.A3( u1_u5_u4_n114 ) , .A2( u1_u5_u4_n115 ) , .A1( u1_u5_u4_n116 ) , .ZN( u1_u5_u4_n136 ) );
  AOI21_X1 u1_u5_u4_U28 (.A( u1_u5_u4_n113 ) , .ZN( u1_u5_u4_n116 ) , .B2( u1_u5_u4_n173 ) , .B1( u1_u5_u4_n174 ) );
  AOI21_X1 u1_u5_u4_U29 (.ZN( u1_u5_u4_n115 ) , .B2( u1_u5_u4_n145 ) , .B1( u1_u5_u4_n146 ) , .A( u1_u5_u4_n156 ) );
  NOR2_X1 u1_u5_u4_U3 (.ZN( u1_u5_u4_n121 ) , .A1( u1_u5_u4_n181 ) , .A2( u1_u5_u4_n182 ) );
  OAI22_X1 u1_u5_u4_U30 (.ZN( u1_u5_u4_n114 ) , .A2( u1_u5_u4_n121 ) , .B1( u1_u5_u4_n160 ) , .B2( u1_u5_u4_n170 ) , .A1( u1_u5_u4_n171 ) );
  INV_X1 u1_u5_u4_U31 (.A( u1_u5_u4_n158 ) , .ZN( u1_u5_u4_n182 ) );
  INV_X1 u1_u5_u4_U32 (.ZN( u1_u5_u4_n181 ) , .A( u1_u5_u4_n96 ) );
  INV_X1 u1_u5_u4_U33 (.A( u1_u5_u4_n144 ) , .ZN( u1_u5_u4_n179 ) );
  INV_X1 u1_u5_u4_U34 (.A( u1_u5_u4_n157 ) , .ZN( u1_u5_u4_n178 ) );
  NAND2_X1 u1_u5_u4_U35 (.A2( u1_u5_u4_n154 ) , .A1( u1_u5_u4_n96 ) , .ZN( u1_u5_u4_n97 ) );
  INV_X1 u1_u5_u4_U36 (.ZN( u1_u5_u4_n186 ) , .A( u1_u5_u4_n95 ) );
  OAI221_X1 u1_u5_u4_U37 (.C1( u1_u5_u4_n134 ) , .B1( u1_u5_u4_n158 ) , .B2( u1_u5_u4_n171 ) , .C2( u1_u5_u4_n173 ) , .A( u1_u5_u4_n94 ) , .ZN( u1_u5_u4_n95 ) );
  AOI222_X1 u1_u5_u4_U38 (.B2( u1_u5_u4_n132 ) , .A1( u1_u5_u4_n138 ) , .C2( u1_u5_u4_n175 ) , .A2( u1_u5_u4_n179 ) , .C1( u1_u5_u4_n181 ) , .B1( u1_u5_u4_n185 ) , .ZN( u1_u5_u4_n94 ) );
  INV_X1 u1_u5_u4_U39 (.A( u1_u5_u4_n113 ) , .ZN( u1_u5_u4_n185 ) );
  INV_X1 u1_u5_u4_U4 (.A( u1_u5_u4_n117 ) , .ZN( u1_u5_u4_n184 ) );
  INV_X1 u1_u5_u4_U40 (.A( u1_u5_u4_n143 ) , .ZN( u1_u5_u4_n183 ) );
  NOR2_X1 u1_u5_u4_U41 (.ZN( u1_u5_u4_n138 ) , .A1( u1_u5_u4_n168 ) , .A2( u1_u5_u4_n169 ) );
  NOR2_X1 u1_u5_u4_U42 (.A1( u1_u5_u4_n150 ) , .A2( u1_u5_u4_n152 ) , .ZN( u1_u5_u4_n153 ) );
  NOR2_X1 u1_u5_u4_U43 (.A2( u1_u5_u4_n128 ) , .A1( u1_u5_u4_n138 ) , .ZN( u1_u5_u4_n156 ) );
  AOI22_X1 u1_u5_u4_U44 (.B2( u1_u5_u4_n122 ) , .A1( u1_u5_u4_n123 ) , .ZN( u1_u5_u4_n124 ) , .B1( u1_u5_u4_n128 ) , .A2( u1_u5_u4_n172 ) );
  INV_X1 u1_u5_u4_U45 (.A( u1_u5_u4_n153 ) , .ZN( u1_u5_u4_n172 ) );
  NAND2_X1 u1_u5_u4_U46 (.A2( u1_u5_u4_n120 ) , .ZN( u1_u5_u4_n123 ) , .A1( u1_u5_u4_n161 ) );
  AOI22_X1 u1_u5_u4_U47 (.B2( u1_u5_u4_n132 ) , .A2( u1_u5_u4_n133 ) , .ZN( u1_u5_u4_n140 ) , .A1( u1_u5_u4_n150 ) , .B1( u1_u5_u4_n179 ) );
  NAND2_X1 u1_u5_u4_U48 (.ZN( u1_u5_u4_n133 ) , .A2( u1_u5_u4_n146 ) , .A1( u1_u5_u4_n154 ) );
  NAND2_X1 u1_u5_u4_U49 (.A1( u1_u5_u4_n103 ) , .ZN( u1_u5_u4_n154 ) , .A2( u1_u5_u4_n98 ) );
  NOR4_X1 u1_u5_u4_U5 (.A4( u1_u5_u4_n106 ) , .A3( u1_u5_u4_n107 ) , .A2( u1_u5_u4_n108 ) , .A1( u1_u5_u4_n109 ) , .ZN( u1_u5_u4_n110 ) );
  NAND2_X1 u1_u5_u4_U50 (.A1( u1_u5_u4_n101 ) , .ZN( u1_u5_u4_n158 ) , .A2( u1_u5_u4_n99 ) );
  AOI21_X1 u1_u5_u4_U51 (.ZN( u1_u5_u4_n127 ) , .A( u1_u5_u4_n136 ) , .B2( u1_u5_u4_n150 ) , .B1( u1_u5_u4_n180 ) );
  INV_X1 u1_u5_u4_U52 (.A( u1_u5_u4_n160 ) , .ZN( u1_u5_u4_n180 ) );
  NAND2_X1 u1_u5_u4_U53 (.A2( u1_u5_u4_n104 ) , .A1( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n146 ) );
  NAND2_X1 u1_u5_u4_U54 (.A2( u1_u5_u4_n101 ) , .A1( u1_u5_u4_n102 ) , .ZN( u1_u5_u4_n160 ) );
  NAND2_X1 u1_u5_u4_U55 (.ZN( u1_u5_u4_n134 ) , .A1( u1_u5_u4_n98 ) , .A2( u1_u5_u4_n99 ) );
  NAND2_X1 u1_u5_u4_U56 (.A1( u1_u5_u4_n103 ) , .A2( u1_u5_u4_n104 ) , .ZN( u1_u5_u4_n143 ) );
  NAND2_X1 u1_u5_u4_U57 (.A2( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n145 ) , .A1( u1_u5_u4_n98 ) );
  NAND2_X1 u1_u5_u4_U58 (.A1( u1_u5_u4_n100 ) , .A2( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n120 ) );
  NAND2_X1 u1_u5_u4_U59 (.A1( u1_u5_u4_n102 ) , .A2( u1_u5_u4_n104 ) , .ZN( u1_u5_u4_n148 ) );
  AOI21_X1 u1_u5_u4_U6 (.ZN( u1_u5_u4_n106 ) , .B2( u1_u5_u4_n146 ) , .B1( u1_u5_u4_n158 ) , .A( u1_u5_u4_n170 ) );
  NAND2_X1 u1_u5_u4_U60 (.A2( u1_u5_u4_n100 ) , .A1( u1_u5_u4_n103 ) , .ZN( u1_u5_u4_n157 ) );
  INV_X1 u1_u5_u4_U61 (.A( u1_u5_u4_n150 ) , .ZN( u1_u5_u4_n173 ) );
  INV_X1 u1_u5_u4_U62 (.A( u1_u5_u4_n152 ) , .ZN( u1_u5_u4_n171 ) );
  NAND2_X1 u1_u5_u4_U63 (.A1( u1_u5_u4_n100 ) , .ZN( u1_u5_u4_n118 ) , .A2( u1_u5_u4_n99 ) );
  NAND2_X1 u1_u5_u4_U64 (.A2( u1_u5_u4_n100 ) , .A1( u1_u5_u4_n102 ) , .ZN( u1_u5_u4_n144 ) );
  NAND2_X1 u1_u5_u4_U65 (.A2( u1_u5_u4_n101 ) , .A1( u1_u5_u4_n105 ) , .ZN( u1_u5_u4_n96 ) );
  INV_X1 u1_u5_u4_U66 (.A( u1_u5_u4_n128 ) , .ZN( u1_u5_u4_n174 ) );
  NAND2_X1 u1_u5_u4_U67 (.A2( u1_u5_u4_n102 ) , .ZN( u1_u5_u4_n119 ) , .A1( u1_u5_u4_n98 ) );
  NAND2_X1 u1_u5_u4_U68 (.A2( u1_u5_u4_n101 ) , .A1( u1_u5_u4_n103 ) , .ZN( u1_u5_u4_n147 ) );
  NAND2_X1 u1_u5_u4_U69 (.A2( u1_u5_u4_n104 ) , .ZN( u1_u5_u4_n113 ) , .A1( u1_u5_u4_n99 ) );
  AOI21_X1 u1_u5_u4_U7 (.ZN( u1_u5_u4_n108 ) , .B2( u1_u5_u4_n134 ) , .B1( u1_u5_u4_n155 ) , .A( u1_u5_u4_n156 ) );
  NOR2_X1 u1_u5_u4_U70 (.A2( u1_u5_X_28 ) , .ZN( u1_u5_u4_n150 ) , .A1( u1_u5_u4_n168 ) );
  NOR2_X1 u1_u5_u4_U71 (.A2( u1_u5_X_29 ) , .ZN( u1_u5_u4_n152 ) , .A1( u1_u5_u4_n169 ) );
  NOR2_X1 u1_u5_u4_U72 (.A2( u1_u5_X_30 ) , .ZN( u1_u5_u4_n105 ) , .A1( u1_u5_u4_n176 ) );
  NOR2_X1 u1_u5_u4_U73 (.A2( u1_u5_X_26 ) , .ZN( u1_u5_u4_n100 ) , .A1( u1_u5_u4_n177 ) );
  NOR2_X1 u1_u5_u4_U74 (.A2( u1_u5_X_28 ) , .A1( u1_u5_X_29 ) , .ZN( u1_u5_u4_n128 ) );
  NOR2_X1 u1_u5_u4_U75 (.A2( u1_u5_X_27 ) , .A1( u1_u5_X_30 ) , .ZN( u1_u5_u4_n102 ) );
  NOR2_X1 u1_u5_u4_U76 (.A2( u1_u5_X_25 ) , .A1( u1_u5_X_26 ) , .ZN( u1_u5_u4_n98 ) );
  AND2_X1 u1_u5_u4_U77 (.A2( u1_u5_X_25 ) , .A1( u1_u5_X_26 ) , .ZN( u1_u5_u4_n104 ) );
  AND2_X1 u1_u5_u4_U78 (.A1( u1_u5_X_30 ) , .A2( u1_u5_u4_n176 ) , .ZN( u1_u5_u4_n99 ) );
  AND2_X1 u1_u5_u4_U79 (.A1( u1_u5_X_26 ) , .ZN( u1_u5_u4_n101 ) , .A2( u1_u5_u4_n177 ) );
  AOI21_X1 u1_u5_u4_U8 (.ZN( u1_u5_u4_n109 ) , .A( u1_u5_u4_n153 ) , .B1( u1_u5_u4_n159 ) , .B2( u1_u5_u4_n184 ) );
  AND2_X1 u1_u5_u4_U80 (.A1( u1_u5_X_27 ) , .A2( u1_u5_X_30 ) , .ZN( u1_u5_u4_n103 ) );
  INV_X1 u1_u5_u4_U81 (.A( u1_u5_X_28 ) , .ZN( u1_u5_u4_n169 ) );
  INV_X1 u1_u5_u4_U82 (.A( u1_u5_X_29 ) , .ZN( u1_u5_u4_n168 ) );
  INV_X1 u1_u5_u4_U83 (.A( u1_u5_X_25 ) , .ZN( u1_u5_u4_n177 ) );
  INV_X1 u1_u5_u4_U84 (.A( u1_u5_X_27 ) , .ZN( u1_u5_u4_n176 ) );
  NAND4_X1 u1_u5_u4_U85 (.ZN( u1_out5_25 ) , .A4( u1_u5_u4_n139 ) , .A3( u1_u5_u4_n140 ) , .A2( u1_u5_u4_n141 ) , .A1( u1_u5_u4_n142 ) );
  OAI21_X1 u1_u5_u4_U86 (.A( u1_u5_u4_n128 ) , .B2( u1_u5_u4_n129 ) , .B1( u1_u5_u4_n130 ) , .ZN( u1_u5_u4_n142 ) );
  OAI21_X1 u1_u5_u4_U87 (.B2( u1_u5_u4_n131 ) , .ZN( u1_u5_u4_n141 ) , .A( u1_u5_u4_n175 ) , .B1( u1_u5_u4_n183 ) );
  NAND4_X1 u1_u5_u4_U88 (.ZN( u1_out5_14 ) , .A4( u1_u5_u4_n124 ) , .A3( u1_u5_u4_n125 ) , .A2( u1_u5_u4_n126 ) , .A1( u1_u5_u4_n127 ) );
  AOI22_X1 u1_u5_u4_U89 (.B2( u1_u5_u4_n117 ) , .ZN( u1_u5_u4_n126 ) , .A1( u1_u5_u4_n129 ) , .B1( u1_u5_u4_n152 ) , .A2( u1_u5_u4_n175 ) );
  AOI211_X1 u1_u5_u4_U9 (.B( u1_u5_u4_n136 ) , .A( u1_u5_u4_n137 ) , .C2( u1_u5_u4_n138 ) , .ZN( u1_u5_u4_n139 ) , .C1( u1_u5_u4_n182 ) );
  AOI22_X1 u1_u5_u4_U90 (.ZN( u1_u5_u4_n125 ) , .B2( u1_u5_u4_n131 ) , .A2( u1_u5_u4_n132 ) , .B1( u1_u5_u4_n138 ) , .A1( u1_u5_u4_n178 ) );
  NAND4_X1 u1_u5_u4_U91 (.ZN( u1_out5_8 ) , .A4( u1_u5_u4_n110 ) , .A3( u1_u5_u4_n111 ) , .A2( u1_u5_u4_n112 ) , .A1( u1_u5_u4_n186 ) );
  NAND2_X1 u1_u5_u4_U92 (.ZN( u1_u5_u4_n112 ) , .A2( u1_u5_u4_n130 ) , .A1( u1_u5_u4_n150 ) );
  AOI22_X1 u1_u5_u4_U93 (.ZN( u1_u5_u4_n111 ) , .B2( u1_u5_u4_n132 ) , .A1( u1_u5_u4_n152 ) , .B1( u1_u5_u4_n178 ) , .A2( u1_u5_u4_n97 ) );
  AOI22_X1 u1_u5_u4_U94 (.B2( u1_u5_u4_n149 ) , .B1( u1_u5_u4_n150 ) , .A2( u1_u5_u4_n151 ) , .A1( u1_u5_u4_n152 ) , .ZN( u1_u5_u4_n167 ) );
  NOR4_X1 u1_u5_u4_U95 (.A4( u1_u5_u4_n162 ) , .A3( u1_u5_u4_n163 ) , .A2( u1_u5_u4_n164 ) , .A1( u1_u5_u4_n165 ) , .ZN( u1_u5_u4_n166 ) );
  NAND3_X1 u1_u5_u4_U96 (.ZN( u1_out5_3 ) , .A3( u1_u5_u4_n166 ) , .A1( u1_u5_u4_n167 ) , .A2( u1_u5_u4_n186 ) );
  NAND3_X1 u1_u5_u4_U97 (.A3( u1_u5_u4_n146 ) , .A2( u1_u5_u4_n147 ) , .A1( u1_u5_u4_n148 ) , .ZN( u1_u5_u4_n149 ) );
  NAND3_X1 u1_u5_u4_U98 (.A3( u1_u5_u4_n143 ) , .A2( u1_u5_u4_n144 ) , .A1( u1_u5_u4_n145 ) , .ZN( u1_u5_u4_n151 ) );
  NAND3_X1 u1_u5_u4_U99 (.A3( u1_u5_u4_n121 ) , .ZN( u1_u5_u4_n122 ) , .A2( u1_u5_u4_n144 ) , .A1( u1_u5_u4_n154 ) );
  INV_X1 u1_u5_u5_U10 (.A( u1_u5_u5_n121 ) , .ZN( u1_u5_u5_n177 ) );
  NOR3_X1 u1_u5_u5_U100 (.A3( u1_u5_u5_n141 ) , .A1( u1_u5_u5_n142 ) , .ZN( u1_u5_u5_n143 ) , .A2( u1_u5_u5_n191 ) );
  NAND4_X1 u1_u5_u5_U101 (.ZN( u1_out5_4 ) , .A4( u1_u5_u5_n112 ) , .A2( u1_u5_u5_n113 ) , .A1( u1_u5_u5_n114 ) , .A3( u1_u5_u5_n195 ) );
  AOI211_X1 u1_u5_u5_U102 (.A( u1_u5_u5_n110 ) , .C1( u1_u5_u5_n111 ) , .ZN( u1_u5_u5_n112 ) , .B( u1_u5_u5_n118 ) , .C2( u1_u5_u5_n177 ) );
  AOI222_X1 u1_u5_u5_U103 (.ZN( u1_u5_u5_n113 ) , .A1( u1_u5_u5_n131 ) , .C1( u1_u5_u5_n148 ) , .B2( u1_u5_u5_n174 ) , .C2( u1_u5_u5_n178 ) , .A2( u1_u5_u5_n179 ) , .B1( u1_u5_u5_n99 ) );
  NAND3_X1 u1_u5_u5_U104 (.A2( u1_u5_u5_n154 ) , .A3( u1_u5_u5_n158 ) , .A1( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n99 ) );
  NOR2_X1 u1_u5_u5_U11 (.ZN( u1_u5_u5_n160 ) , .A2( u1_u5_u5_n173 ) , .A1( u1_u5_u5_n177 ) );
  INV_X1 u1_u5_u5_U12 (.A( u1_u5_u5_n150 ) , .ZN( u1_u5_u5_n174 ) );
  AOI21_X1 u1_u5_u5_U13 (.A( u1_u5_u5_n160 ) , .B2( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n162 ) , .B1( u1_u5_u5_n192 ) );
  INV_X1 u1_u5_u5_U14 (.A( u1_u5_u5_n159 ) , .ZN( u1_u5_u5_n192 ) );
  AOI21_X1 u1_u5_u5_U15 (.A( u1_u5_u5_n156 ) , .B2( u1_u5_u5_n157 ) , .B1( u1_u5_u5_n158 ) , .ZN( u1_u5_u5_n163 ) );
  AOI21_X1 u1_u5_u5_U16 (.B2( u1_u5_u5_n139 ) , .B1( u1_u5_u5_n140 ) , .ZN( u1_u5_u5_n141 ) , .A( u1_u5_u5_n150 ) );
  OAI21_X1 u1_u5_u5_U17 (.A( u1_u5_u5_n133 ) , .B2( u1_u5_u5_n134 ) , .B1( u1_u5_u5_n135 ) , .ZN( u1_u5_u5_n142 ) );
  OAI21_X1 u1_u5_u5_U18 (.ZN( u1_u5_u5_n133 ) , .B2( u1_u5_u5_n147 ) , .A( u1_u5_u5_n173 ) , .B1( u1_u5_u5_n188 ) );
  NAND2_X1 u1_u5_u5_U19 (.A2( u1_u5_u5_n119 ) , .A1( u1_u5_u5_n123 ) , .ZN( u1_u5_u5_n137 ) );
  INV_X1 u1_u5_u5_U20 (.A( u1_u5_u5_n155 ) , .ZN( u1_u5_u5_n194 ) );
  NAND2_X1 u1_u5_u5_U21 (.A1( u1_u5_u5_n121 ) , .ZN( u1_u5_u5_n132 ) , .A2( u1_u5_u5_n172 ) );
  NAND2_X1 u1_u5_u5_U22 (.A2( u1_u5_u5_n122 ) , .ZN( u1_u5_u5_n136 ) , .A1( u1_u5_u5_n154 ) );
  NAND2_X1 u1_u5_u5_U23 (.A2( u1_u5_u5_n119 ) , .A1( u1_u5_u5_n120 ) , .ZN( u1_u5_u5_n159 ) );
  INV_X1 u1_u5_u5_U24 (.A( u1_u5_u5_n156 ) , .ZN( u1_u5_u5_n175 ) );
  INV_X1 u1_u5_u5_U25 (.A( u1_u5_u5_n158 ) , .ZN( u1_u5_u5_n188 ) );
  INV_X1 u1_u5_u5_U26 (.A( u1_u5_u5_n152 ) , .ZN( u1_u5_u5_n179 ) );
  INV_X1 u1_u5_u5_U27 (.A( u1_u5_u5_n140 ) , .ZN( u1_u5_u5_n182 ) );
  INV_X1 u1_u5_u5_U28 (.A( u1_u5_u5_n151 ) , .ZN( u1_u5_u5_n183 ) );
  INV_X1 u1_u5_u5_U29 (.A( u1_u5_u5_n123 ) , .ZN( u1_u5_u5_n185 ) );
  NOR2_X1 u1_u5_u5_U3 (.ZN( u1_u5_u5_n134 ) , .A1( u1_u5_u5_n183 ) , .A2( u1_u5_u5_n190 ) );
  INV_X1 u1_u5_u5_U30 (.A( u1_u5_u5_n161 ) , .ZN( u1_u5_u5_n184 ) );
  INV_X1 u1_u5_u5_U31 (.A( u1_u5_u5_n139 ) , .ZN( u1_u5_u5_n189 ) );
  INV_X1 u1_u5_u5_U32 (.A( u1_u5_u5_n157 ) , .ZN( u1_u5_u5_n190 ) );
  INV_X1 u1_u5_u5_U33 (.A( u1_u5_u5_n120 ) , .ZN( u1_u5_u5_n193 ) );
  NAND2_X1 u1_u5_u5_U34 (.ZN( u1_u5_u5_n111 ) , .A1( u1_u5_u5_n140 ) , .A2( u1_u5_u5_n155 ) );
  NOR2_X1 u1_u5_u5_U35 (.ZN( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n170 ) , .A2( u1_u5_u5_n180 ) );
  INV_X1 u1_u5_u5_U36 (.A( u1_u5_u5_n117 ) , .ZN( u1_u5_u5_n196 ) );
  OAI221_X1 u1_u5_u5_U37 (.A( u1_u5_u5_n116 ) , .ZN( u1_u5_u5_n117 ) , .B2( u1_u5_u5_n119 ) , .C1( u1_u5_u5_n153 ) , .C2( u1_u5_u5_n158 ) , .B1( u1_u5_u5_n172 ) );
  AOI222_X1 u1_u5_u5_U38 (.ZN( u1_u5_u5_n116 ) , .B2( u1_u5_u5_n145 ) , .C1( u1_u5_u5_n148 ) , .A2( u1_u5_u5_n174 ) , .C2( u1_u5_u5_n177 ) , .B1( u1_u5_u5_n187 ) , .A1( u1_u5_u5_n193 ) );
  INV_X1 u1_u5_u5_U39 (.A( u1_u5_u5_n115 ) , .ZN( u1_u5_u5_n187 ) );
  INV_X1 u1_u5_u5_U4 (.A( u1_u5_u5_n138 ) , .ZN( u1_u5_u5_n191 ) );
  AOI22_X1 u1_u5_u5_U40 (.B2( u1_u5_u5_n131 ) , .A2( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n169 ) , .B1( u1_u5_u5_n174 ) , .A1( u1_u5_u5_n185 ) );
  NOR2_X1 u1_u5_u5_U41 (.A1( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n150 ) , .A2( u1_u5_u5_n173 ) );
  AOI21_X1 u1_u5_u5_U42 (.A( u1_u5_u5_n118 ) , .B2( u1_u5_u5_n145 ) , .ZN( u1_u5_u5_n168 ) , .B1( u1_u5_u5_n186 ) );
  INV_X1 u1_u5_u5_U43 (.A( u1_u5_u5_n122 ) , .ZN( u1_u5_u5_n186 ) );
  NOR2_X1 u1_u5_u5_U44 (.A1( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n152 ) , .A2( u1_u5_u5_n176 ) );
  NOR2_X1 u1_u5_u5_U45 (.A1( u1_u5_u5_n115 ) , .ZN( u1_u5_u5_n118 ) , .A2( u1_u5_u5_n153 ) );
  NOR2_X1 u1_u5_u5_U46 (.A2( u1_u5_u5_n145 ) , .ZN( u1_u5_u5_n156 ) , .A1( u1_u5_u5_n174 ) );
  NOR2_X1 u1_u5_u5_U47 (.ZN( u1_u5_u5_n121 ) , .A2( u1_u5_u5_n145 ) , .A1( u1_u5_u5_n176 ) );
  AOI22_X1 u1_u5_u5_U48 (.ZN( u1_u5_u5_n114 ) , .A2( u1_u5_u5_n137 ) , .A1( u1_u5_u5_n145 ) , .B2( u1_u5_u5_n175 ) , .B1( u1_u5_u5_n193 ) );
  OAI211_X1 u1_u5_u5_U49 (.B( u1_u5_u5_n124 ) , .A( u1_u5_u5_n125 ) , .C2( u1_u5_u5_n126 ) , .C1( u1_u5_u5_n127 ) , .ZN( u1_u5_u5_n128 ) );
  OAI21_X1 u1_u5_u5_U5 (.B2( u1_u5_u5_n136 ) , .B1( u1_u5_u5_n137 ) , .ZN( u1_u5_u5_n138 ) , .A( u1_u5_u5_n177 ) );
  NOR3_X1 u1_u5_u5_U50 (.ZN( u1_u5_u5_n127 ) , .A1( u1_u5_u5_n136 ) , .A3( u1_u5_u5_n148 ) , .A2( u1_u5_u5_n182 ) );
  OAI21_X1 u1_u5_u5_U51 (.ZN( u1_u5_u5_n124 ) , .A( u1_u5_u5_n177 ) , .B2( u1_u5_u5_n183 ) , .B1( u1_u5_u5_n189 ) );
  OAI21_X1 u1_u5_u5_U52 (.ZN( u1_u5_u5_n125 ) , .A( u1_u5_u5_n174 ) , .B2( u1_u5_u5_n185 ) , .B1( u1_u5_u5_n190 ) );
  AOI21_X1 u1_u5_u5_U53 (.A( u1_u5_u5_n153 ) , .B2( u1_u5_u5_n154 ) , .B1( u1_u5_u5_n155 ) , .ZN( u1_u5_u5_n164 ) );
  AOI21_X1 u1_u5_u5_U54 (.ZN( u1_u5_u5_n110 ) , .B1( u1_u5_u5_n122 ) , .B2( u1_u5_u5_n139 ) , .A( u1_u5_u5_n153 ) );
  INV_X1 u1_u5_u5_U55 (.A( u1_u5_u5_n153 ) , .ZN( u1_u5_u5_n176 ) );
  INV_X1 u1_u5_u5_U56 (.A( u1_u5_u5_n126 ) , .ZN( u1_u5_u5_n173 ) );
  AND2_X1 u1_u5_u5_U57 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n147 ) );
  AND2_X1 u1_u5_u5_U58 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n148 ) );
  NAND2_X1 u1_u5_u5_U59 (.A1( u1_u5_u5_n105 ) , .A2( u1_u5_u5_n106 ) , .ZN( u1_u5_u5_n158 ) );
  INV_X1 u1_u5_u5_U6 (.A( u1_u5_u5_n135 ) , .ZN( u1_u5_u5_n178 ) );
  NAND2_X1 u1_u5_u5_U60 (.A2( u1_u5_u5_n108 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n139 ) );
  NAND2_X1 u1_u5_u5_U61 (.A1( u1_u5_u5_n106 ) , .A2( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n119 ) );
  NAND2_X1 u1_u5_u5_U62 (.A2( u1_u5_u5_n103 ) , .A1( u1_u5_u5_n105 ) , .ZN( u1_u5_u5_n140 ) );
  NAND2_X1 u1_u5_u5_U63 (.A2( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n105 ) , .ZN( u1_u5_u5_n155 ) );
  NAND2_X1 u1_u5_u5_U64 (.A2( u1_u5_u5_n106 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n122 ) );
  NAND2_X1 u1_u5_u5_U65 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n106 ) , .ZN( u1_u5_u5_n115 ) );
  NAND2_X1 u1_u5_u5_U66 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n103 ) , .ZN( u1_u5_u5_n161 ) );
  NAND2_X1 u1_u5_u5_U67 (.A1( u1_u5_u5_n105 ) , .A2( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n154 ) );
  INV_X1 u1_u5_u5_U68 (.A( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n172 ) );
  NAND2_X1 u1_u5_u5_U69 (.A1( u1_u5_u5_n103 ) , .A2( u1_u5_u5_n108 ) , .ZN( u1_u5_u5_n123 ) );
  OAI22_X1 u1_u5_u5_U7 (.B2( u1_u5_u5_n149 ) , .B1( u1_u5_u5_n150 ) , .A2( u1_u5_u5_n151 ) , .A1( u1_u5_u5_n152 ) , .ZN( u1_u5_u5_n165 ) );
  NAND2_X1 u1_u5_u5_U70 (.A2( u1_u5_u5_n103 ) , .A1( u1_u5_u5_n107 ) , .ZN( u1_u5_u5_n151 ) );
  NAND2_X1 u1_u5_u5_U71 (.A2( u1_u5_u5_n107 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n120 ) );
  NAND2_X1 u1_u5_u5_U72 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n109 ) , .ZN( u1_u5_u5_n157 ) );
  AND2_X1 u1_u5_u5_U73 (.A2( u1_u5_u5_n100 ) , .A1( u1_u5_u5_n104 ) , .ZN( u1_u5_u5_n131 ) );
  INV_X1 u1_u5_u5_U74 (.A( u1_u5_u5_n102 ) , .ZN( u1_u5_u5_n195 ) );
  OAI221_X1 u1_u5_u5_U75 (.A( u1_u5_u5_n101 ) , .ZN( u1_u5_u5_n102 ) , .C2( u1_u5_u5_n115 ) , .C1( u1_u5_u5_n126 ) , .B1( u1_u5_u5_n134 ) , .B2( u1_u5_u5_n160 ) );
  OAI21_X1 u1_u5_u5_U76 (.ZN( u1_u5_u5_n101 ) , .B1( u1_u5_u5_n137 ) , .A( u1_u5_u5_n146 ) , .B2( u1_u5_u5_n147 ) );
  NOR2_X1 u1_u5_u5_U77 (.A2( u1_u5_X_34 ) , .A1( u1_u5_X_35 ) , .ZN( u1_u5_u5_n145 ) );
  NOR2_X1 u1_u5_u5_U78 (.A2( u1_u5_X_34 ) , .ZN( u1_u5_u5_n146 ) , .A1( u1_u5_u5_n171 ) );
  NOR2_X1 u1_u5_u5_U79 (.A2( u1_u5_X_31 ) , .A1( u1_u5_X_32 ) , .ZN( u1_u5_u5_n103 ) );
  NOR3_X1 u1_u5_u5_U8 (.A2( u1_u5_u5_n147 ) , .A1( u1_u5_u5_n148 ) , .ZN( u1_u5_u5_n149 ) , .A3( u1_u5_u5_n194 ) );
  NOR2_X1 u1_u5_u5_U80 (.A2( u1_u5_X_36 ) , .ZN( u1_u5_u5_n105 ) , .A1( u1_u5_u5_n180 ) );
  NOR2_X1 u1_u5_u5_U81 (.A2( u1_u5_X_33 ) , .ZN( u1_u5_u5_n108 ) , .A1( u1_u5_u5_n170 ) );
  NOR2_X1 u1_u5_u5_U82 (.A2( u1_u5_X_33 ) , .A1( u1_u5_X_36 ) , .ZN( u1_u5_u5_n107 ) );
  NOR2_X1 u1_u5_u5_U83 (.A2( u1_u5_X_31 ) , .ZN( u1_u5_u5_n104 ) , .A1( u1_u5_u5_n181 ) );
  NAND2_X1 u1_u5_u5_U84 (.A2( u1_u5_X_34 ) , .A1( u1_u5_X_35 ) , .ZN( u1_u5_u5_n153 ) );
  NAND2_X1 u1_u5_u5_U85 (.A1( u1_u5_X_34 ) , .ZN( u1_u5_u5_n126 ) , .A2( u1_u5_u5_n171 ) );
  AND2_X1 u1_u5_u5_U86 (.A1( u1_u5_X_31 ) , .A2( u1_u5_X_32 ) , .ZN( u1_u5_u5_n106 ) );
  AND2_X1 u1_u5_u5_U87 (.A1( u1_u5_X_31 ) , .ZN( u1_u5_u5_n109 ) , .A2( u1_u5_u5_n181 ) );
  INV_X1 u1_u5_u5_U88 (.A( u1_u5_X_33 ) , .ZN( u1_u5_u5_n180 ) );
  INV_X1 u1_u5_u5_U89 (.A( u1_u5_X_35 ) , .ZN( u1_u5_u5_n171 ) );
  NOR2_X1 u1_u5_u5_U9 (.ZN( u1_u5_u5_n135 ) , .A1( u1_u5_u5_n173 ) , .A2( u1_u5_u5_n176 ) );
  INV_X1 u1_u5_u5_U90 (.A( u1_u5_X_36 ) , .ZN( u1_u5_u5_n170 ) );
  INV_X1 u1_u5_u5_U91 (.A( u1_u5_X_32 ) , .ZN( u1_u5_u5_n181 ) );
  NAND4_X1 u1_u5_u5_U92 (.ZN( u1_out5_29 ) , .A4( u1_u5_u5_n129 ) , .A3( u1_u5_u5_n130 ) , .A2( u1_u5_u5_n168 ) , .A1( u1_u5_u5_n196 ) );
  AOI221_X1 u1_u5_u5_U93 (.A( u1_u5_u5_n128 ) , .ZN( u1_u5_u5_n129 ) , .C2( u1_u5_u5_n132 ) , .B2( u1_u5_u5_n159 ) , .B1( u1_u5_u5_n176 ) , .C1( u1_u5_u5_n184 ) );
  AOI222_X1 u1_u5_u5_U94 (.ZN( u1_u5_u5_n130 ) , .A2( u1_u5_u5_n146 ) , .B1( u1_u5_u5_n147 ) , .C2( u1_u5_u5_n175 ) , .B2( u1_u5_u5_n179 ) , .A1( u1_u5_u5_n188 ) , .C1( u1_u5_u5_n194 ) );
  NAND4_X1 u1_u5_u5_U95 (.ZN( u1_out5_19 ) , .A4( u1_u5_u5_n166 ) , .A3( u1_u5_u5_n167 ) , .A2( u1_u5_u5_n168 ) , .A1( u1_u5_u5_n169 ) );
  AOI22_X1 u1_u5_u5_U96 (.B2( u1_u5_u5_n145 ) , .A2( u1_u5_u5_n146 ) , .ZN( u1_u5_u5_n167 ) , .B1( u1_u5_u5_n182 ) , .A1( u1_u5_u5_n189 ) );
  NOR4_X1 u1_u5_u5_U97 (.A4( u1_u5_u5_n162 ) , .A3( u1_u5_u5_n163 ) , .A2( u1_u5_u5_n164 ) , .A1( u1_u5_u5_n165 ) , .ZN( u1_u5_u5_n166 ) );
  NAND4_X1 u1_u5_u5_U98 (.ZN( u1_out5_11 ) , .A4( u1_u5_u5_n143 ) , .A3( u1_u5_u5_n144 ) , .A2( u1_u5_u5_n169 ) , .A1( u1_u5_u5_n196 ) );
  AOI22_X1 u1_u5_u5_U99 (.A2( u1_u5_u5_n132 ) , .ZN( u1_u5_u5_n144 ) , .B2( u1_u5_u5_n145 ) , .B1( u1_u5_u5_n184 ) , .A1( u1_u5_u5_n194 ) );
  OAI21_X1 u1_u5_u6_U10 (.A( u1_u5_u6_n159 ) , .B1( u1_u5_u6_n169 ) , .B2( u1_u5_u6_n173 ) , .ZN( u1_u5_u6_n90 ) );
  INV_X1 u1_u5_u6_U11 (.ZN( u1_u5_u6_n172 ) , .A( u1_u5_u6_n88 ) );
  AOI22_X1 u1_u5_u6_U12 (.A2( u1_u5_u6_n151 ) , .B2( u1_u5_u6_n161 ) , .A1( u1_u5_u6_n167 ) , .B1( u1_u5_u6_n170 ) , .ZN( u1_u5_u6_n89 ) );
  AOI21_X1 u1_u5_u6_U13 (.ZN( u1_u5_u6_n106 ) , .A( u1_u5_u6_n142 ) , .B2( u1_u5_u6_n159 ) , .B1( u1_u5_u6_n164 ) );
  INV_X1 u1_u5_u6_U14 (.A( u1_u5_u6_n155 ) , .ZN( u1_u5_u6_n161 ) );
  INV_X1 u1_u5_u6_U15 (.A( u1_u5_u6_n128 ) , .ZN( u1_u5_u6_n164 ) );
  NAND2_X1 u1_u5_u6_U16 (.ZN( u1_u5_u6_n110 ) , .A1( u1_u5_u6_n122 ) , .A2( u1_u5_u6_n129 ) );
  NAND2_X1 u1_u5_u6_U17 (.ZN( u1_u5_u6_n124 ) , .A2( u1_u5_u6_n146 ) , .A1( u1_u5_u6_n148 ) );
  INV_X1 u1_u5_u6_U18 (.A( u1_u5_u6_n132 ) , .ZN( u1_u5_u6_n171 ) );
  AND2_X1 u1_u5_u6_U19 (.A1( u1_u5_u6_n100 ) , .ZN( u1_u5_u6_n130 ) , .A2( u1_u5_u6_n147 ) );
  INV_X1 u1_u5_u6_U20 (.A( u1_u5_u6_n127 ) , .ZN( u1_u5_u6_n173 ) );
  INV_X1 u1_u5_u6_U21 (.A( u1_u5_u6_n121 ) , .ZN( u1_u5_u6_n167 ) );
  INV_X1 u1_u5_u6_U22 (.A( u1_u5_u6_n100 ) , .ZN( u1_u5_u6_n169 ) );
  INV_X1 u1_u5_u6_U23 (.A( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n170 ) );
  INV_X1 u1_u5_u6_U24 (.A( u1_u5_u6_n113 ) , .ZN( u1_u5_u6_n168 ) );
  AND2_X1 u1_u5_u6_U25 (.A1( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n119 ) , .ZN( u1_u5_u6_n133 ) );
  AND2_X1 u1_u5_u6_U26 (.A2( u1_u5_u6_n121 ) , .A1( u1_u5_u6_n122 ) , .ZN( u1_u5_u6_n131 ) );
  AND3_X1 u1_u5_u6_U27 (.ZN( u1_u5_u6_n120 ) , .A2( u1_u5_u6_n127 ) , .A1( u1_u5_u6_n132 ) , .A3( u1_u5_u6_n145 ) );
  INV_X1 u1_u5_u6_U28 (.A( u1_u5_u6_n146 ) , .ZN( u1_u5_u6_n163 ) );
  AOI222_X1 u1_u5_u6_U29 (.ZN( u1_u5_u6_n114 ) , .A1( u1_u5_u6_n118 ) , .A2( u1_u5_u6_n126 ) , .B2( u1_u5_u6_n151 ) , .C2( u1_u5_u6_n159 ) , .C1( u1_u5_u6_n168 ) , .B1( u1_u5_u6_n169 ) );
  INV_X1 u1_u5_u6_U3 (.A( u1_u5_u6_n110 ) , .ZN( u1_u5_u6_n166 ) );
  NOR2_X1 u1_u5_u6_U30 (.A1( u1_u5_u6_n162 ) , .A2( u1_u5_u6_n165 ) , .ZN( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U31 (.A1( u1_u5_u6_n144 ) , .ZN( u1_u5_u6_n151 ) , .A2( u1_u5_u6_n158 ) );
  NAND2_X1 u1_u5_u6_U32 (.ZN( u1_u5_u6_n132 ) , .A1( u1_u5_u6_n91 ) , .A2( u1_u5_u6_n97 ) );
  NOR2_X1 u1_u5_u6_U33 (.A2( u1_u5_u6_n126 ) , .ZN( u1_u5_u6_n155 ) , .A1( u1_u5_u6_n160 ) );
  NAND2_X1 u1_u5_u6_U34 (.ZN( u1_u5_u6_n146 ) , .A2( u1_u5_u6_n94 ) , .A1( u1_u5_u6_n99 ) );
  AOI21_X1 u1_u5_u6_U35 (.A( u1_u5_u6_n144 ) , .B2( u1_u5_u6_n145 ) , .B1( u1_u5_u6_n146 ) , .ZN( u1_u5_u6_n150 ) );
  INV_X1 u1_u5_u6_U36 (.A( u1_u5_u6_n111 ) , .ZN( u1_u5_u6_n158 ) );
  NAND2_X1 u1_u5_u6_U37 (.ZN( u1_u5_u6_n127 ) , .A1( u1_u5_u6_n91 ) , .A2( u1_u5_u6_n92 ) );
  NAND2_X1 u1_u5_u6_U38 (.ZN( u1_u5_u6_n129 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n96 ) );
  INV_X1 u1_u5_u6_U39 (.A( u1_u5_u6_n144 ) , .ZN( u1_u5_u6_n159 ) );
  INV_X1 u1_u5_u6_U4 (.A( u1_u5_u6_n142 ) , .ZN( u1_u5_u6_n174 ) );
  NAND2_X1 u1_u5_u6_U40 (.ZN( u1_u5_u6_n145 ) , .A2( u1_u5_u6_n97 ) , .A1( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U41 (.ZN( u1_u5_u6_n148 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n94 ) );
  NAND2_X1 u1_u5_u6_U42 (.ZN( u1_u5_u6_n108 ) , .A2( u1_u5_u6_n139 ) , .A1( u1_u5_u6_n144 ) );
  NAND2_X1 u1_u5_u6_U43 (.ZN( u1_u5_u6_n121 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n97 ) );
  NAND2_X1 u1_u5_u6_U44 (.ZN( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n95 ) );
  AND2_X1 u1_u5_u6_U45 (.ZN( u1_u5_u6_n118 ) , .A2( u1_u5_u6_n91 ) , .A1( u1_u5_u6_n99 ) );
  AOI22_X1 u1_u5_u6_U46 (.B2( u1_u5_u6_n110 ) , .B1( u1_u5_u6_n111 ) , .A1( u1_u5_u6_n112 ) , .ZN( u1_u5_u6_n115 ) , .A2( u1_u5_u6_n161 ) );
  NAND4_X1 u1_u5_u6_U47 (.A3( u1_u5_u6_n109 ) , .ZN( u1_u5_u6_n112 ) , .A4( u1_u5_u6_n132 ) , .A2( u1_u5_u6_n147 ) , .A1( u1_u5_u6_n166 ) );
  NOR2_X1 u1_u5_u6_U48 (.ZN( u1_u5_u6_n109 ) , .A1( u1_u5_u6_n170 ) , .A2( u1_u5_u6_n173 ) );
  NAND2_X1 u1_u5_u6_U49 (.ZN( u1_u5_u6_n147 ) , .A2( u1_u5_u6_n98 ) , .A1( u1_u5_u6_n99 ) );
  NAND2_X1 u1_u5_u6_U5 (.A2( u1_u5_u6_n143 ) , .ZN( u1_u5_u6_n152 ) , .A1( u1_u5_u6_n166 ) );
  NAND2_X1 u1_u5_u6_U50 (.ZN( u1_u5_u6_n128 ) , .A1( u1_u5_u6_n94 ) , .A2( u1_u5_u6_n96 ) );
  AOI211_X1 u1_u5_u6_U51 (.B( u1_u5_u6_n134 ) , .A( u1_u5_u6_n135 ) , .C1( u1_u5_u6_n136 ) , .ZN( u1_u5_u6_n137 ) , .C2( u1_u5_u6_n151 ) );
  AOI21_X1 u1_u5_u6_U52 (.B2( u1_u5_u6_n132 ) , .B1( u1_u5_u6_n133 ) , .ZN( u1_u5_u6_n134 ) , .A( u1_u5_u6_n158 ) );
  AOI21_X1 u1_u5_u6_U53 (.B1( u1_u5_u6_n131 ) , .ZN( u1_u5_u6_n135 ) , .A( u1_u5_u6_n144 ) , .B2( u1_u5_u6_n146 ) );
  NAND4_X1 u1_u5_u6_U54 (.A4( u1_u5_u6_n127 ) , .A3( u1_u5_u6_n128 ) , .A2( u1_u5_u6_n129 ) , .A1( u1_u5_u6_n130 ) , .ZN( u1_u5_u6_n136 ) );
  NAND2_X1 u1_u5_u6_U55 (.ZN( u1_u5_u6_n119 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n99 ) );
  NAND2_X1 u1_u5_u6_U56 (.ZN( u1_u5_u6_n123 ) , .A2( u1_u5_u6_n91 ) , .A1( u1_u5_u6_n96 ) );
  NAND2_X1 u1_u5_u6_U57 (.ZN( u1_u5_u6_n100 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U58 (.ZN( u1_u5_u6_n122 ) , .A1( u1_u5_u6_n94 ) , .A2( u1_u5_u6_n97 ) );
  INV_X1 u1_u5_u6_U59 (.A( u1_u5_u6_n139 ) , .ZN( u1_u5_u6_n160 ) );
  AOI22_X1 u1_u5_u6_U6 (.B2( u1_u5_u6_n101 ) , .A1( u1_u5_u6_n102 ) , .ZN( u1_u5_u6_n103 ) , .B1( u1_u5_u6_n160 ) , .A2( u1_u5_u6_n161 ) );
  NAND2_X1 u1_u5_u6_U60 (.ZN( u1_u5_u6_n113 ) , .A1( u1_u5_u6_n96 ) , .A2( u1_u5_u6_n98 ) );
  NOR2_X1 u1_u5_u6_U61 (.A2( u1_u5_X_40 ) , .A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n126 ) );
  NOR2_X1 u1_u5_u6_U62 (.A2( u1_u5_X_39 ) , .A1( u1_u5_X_42 ) , .ZN( u1_u5_u6_n92 ) );
  NOR2_X1 u1_u5_u6_U63 (.A2( u1_u5_X_39 ) , .A1( u1_u5_u6_n156 ) , .ZN( u1_u5_u6_n97 ) );
  NOR2_X1 u1_u5_u6_U64 (.A2( u1_u5_X_38 ) , .A1( u1_u5_u6_n165 ) , .ZN( u1_u5_u6_n95 ) );
  NOR2_X1 u1_u5_u6_U65 (.A2( u1_u5_X_41 ) , .ZN( u1_u5_u6_n111 ) , .A1( u1_u5_u6_n157 ) );
  NOR2_X1 u1_u5_u6_U66 (.A2( u1_u5_X_37 ) , .A1( u1_u5_u6_n162 ) , .ZN( u1_u5_u6_n94 ) );
  NOR2_X1 u1_u5_u6_U67 (.A2( u1_u5_X_37 ) , .A1( u1_u5_X_38 ) , .ZN( u1_u5_u6_n91 ) );
  NAND2_X1 u1_u5_u6_U68 (.A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n144 ) , .A2( u1_u5_u6_n157 ) );
  NAND2_X1 u1_u5_u6_U69 (.A2( u1_u5_X_40 ) , .A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n139 ) );
  NOR2_X1 u1_u5_u6_U7 (.A1( u1_u5_u6_n118 ) , .ZN( u1_u5_u6_n143 ) , .A2( u1_u5_u6_n168 ) );
  AND2_X1 u1_u5_u6_U70 (.A1( u1_u5_X_39 ) , .A2( u1_u5_u6_n156 ) , .ZN( u1_u5_u6_n96 ) );
  AND2_X1 u1_u5_u6_U71 (.A1( u1_u5_X_39 ) , .A2( u1_u5_X_42 ) , .ZN( u1_u5_u6_n99 ) );
  INV_X1 u1_u5_u6_U72 (.A( u1_u5_X_40 ) , .ZN( u1_u5_u6_n157 ) );
  INV_X1 u1_u5_u6_U73 (.A( u1_u5_X_37 ) , .ZN( u1_u5_u6_n165 ) );
  INV_X1 u1_u5_u6_U74 (.A( u1_u5_X_38 ) , .ZN( u1_u5_u6_n162 ) );
  INV_X1 u1_u5_u6_U75 (.A( u1_u5_X_42 ) , .ZN( u1_u5_u6_n156 ) );
  NAND4_X1 u1_u5_u6_U76 (.ZN( u1_out5_32 ) , .A4( u1_u5_u6_n103 ) , .A3( u1_u5_u6_n104 ) , .A2( u1_u5_u6_n105 ) , .A1( u1_u5_u6_n106 ) );
  AOI22_X1 u1_u5_u6_U77 (.ZN( u1_u5_u6_n105 ) , .A2( u1_u5_u6_n108 ) , .A1( u1_u5_u6_n118 ) , .B2( u1_u5_u6_n126 ) , .B1( u1_u5_u6_n171 ) );
  AOI22_X1 u1_u5_u6_U78 (.ZN( u1_u5_u6_n104 ) , .A1( u1_u5_u6_n111 ) , .B1( u1_u5_u6_n124 ) , .B2( u1_u5_u6_n151 ) , .A2( u1_u5_u6_n93 ) );
  NAND4_X1 u1_u5_u6_U79 (.ZN( u1_out5_12 ) , .A4( u1_u5_u6_n114 ) , .A3( u1_u5_u6_n115 ) , .A2( u1_u5_u6_n116 ) , .A1( u1_u5_u6_n117 ) );
  AOI21_X1 u1_u5_u6_U8 (.B1( u1_u5_u6_n107 ) , .B2( u1_u5_u6_n132 ) , .A( u1_u5_u6_n158 ) , .ZN( u1_u5_u6_n88 ) );
  OAI22_X1 u1_u5_u6_U80 (.B2( u1_u5_u6_n111 ) , .ZN( u1_u5_u6_n116 ) , .B1( u1_u5_u6_n126 ) , .A2( u1_u5_u6_n164 ) , .A1( u1_u5_u6_n167 ) );
  OAI21_X1 u1_u5_u6_U81 (.A( u1_u5_u6_n108 ) , .ZN( u1_u5_u6_n117 ) , .B2( u1_u5_u6_n141 ) , .B1( u1_u5_u6_n163 ) );
  OAI211_X1 u1_u5_u6_U82 (.ZN( u1_out5_7 ) , .B( u1_u5_u6_n153 ) , .C2( u1_u5_u6_n154 ) , .C1( u1_u5_u6_n155 ) , .A( u1_u5_u6_n174 ) );
  NOR3_X1 u1_u5_u6_U83 (.A1( u1_u5_u6_n141 ) , .ZN( u1_u5_u6_n154 ) , .A3( u1_u5_u6_n164 ) , .A2( u1_u5_u6_n171 ) );
  AOI211_X1 u1_u5_u6_U84 (.B( u1_u5_u6_n149 ) , .A( u1_u5_u6_n150 ) , .C2( u1_u5_u6_n151 ) , .C1( u1_u5_u6_n152 ) , .ZN( u1_u5_u6_n153 ) );
  OAI211_X1 u1_u5_u6_U85 (.ZN( u1_out5_22 ) , .B( u1_u5_u6_n137 ) , .A( u1_u5_u6_n138 ) , .C2( u1_u5_u6_n139 ) , .C1( u1_u5_u6_n140 ) );
  AOI22_X1 u1_u5_u6_U86 (.B1( u1_u5_u6_n124 ) , .A2( u1_u5_u6_n125 ) , .A1( u1_u5_u6_n126 ) , .ZN( u1_u5_u6_n138 ) , .B2( u1_u5_u6_n161 ) );
  AND4_X1 u1_u5_u6_U87 (.A3( u1_u5_u6_n119 ) , .A1( u1_u5_u6_n120 ) , .A4( u1_u5_u6_n129 ) , .ZN( u1_u5_u6_n140 ) , .A2( u1_u5_u6_n143 ) );
  NAND3_X1 u1_u5_u6_U88 (.A2( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n125 ) , .A1( u1_u5_u6_n130 ) , .A3( u1_u5_u6_n131 ) );
  NAND3_X1 u1_u5_u6_U89 (.A3( u1_u5_u6_n133 ) , .ZN( u1_u5_u6_n141 ) , .A1( u1_u5_u6_n145 ) , .A2( u1_u5_u6_n148 ) );
  AOI21_X1 u1_u5_u6_U9 (.B2( u1_u5_u6_n147 ) , .B1( u1_u5_u6_n148 ) , .ZN( u1_u5_u6_n149 ) , .A( u1_u5_u6_n158 ) );
  NAND3_X1 u1_u5_u6_U90 (.ZN( u1_u5_u6_n101 ) , .A3( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n121 ) , .A1( u1_u5_u6_n127 ) );
  NAND3_X1 u1_u5_u6_U91 (.ZN( u1_u5_u6_n102 ) , .A3( u1_u5_u6_n130 ) , .A2( u1_u5_u6_n145 ) , .A1( u1_u5_u6_n166 ) );
  NAND3_X1 u1_u5_u6_U92 (.A3( u1_u5_u6_n113 ) , .A1( u1_u5_u6_n119 ) , .A2( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n93 ) );
  NAND3_X1 u1_u5_u6_U93 (.ZN( u1_u5_u6_n142 ) , .A2( u1_u5_u6_n172 ) , .A3( u1_u5_u6_n89 ) , .A1( u1_u5_u6_n90 ) );
  XOR2_X1 u1_u8_U1 (.B( u1_K9_9 ) , .A( u1_R7_6 ) , .Z( u1_u8_X_9 ) );
  XOR2_X1 u1_u8_U16 (.B( u1_K9_3 ) , .A( u1_R7_2 ) , .Z( u1_u8_X_3 ) );
  XOR2_X1 u1_u8_U2 (.B( u1_K9_8 ) , .A( u1_R7_5 ) , .Z( u1_u8_X_8 ) );
  XOR2_X1 u1_u8_U27 (.B( u1_K9_2 ) , .A( u1_R7_1 ) , .Z( u1_u8_X_2 ) );
  XOR2_X1 u1_u8_U3 (.B( u1_K9_7 ) , .A( u1_R7_4 ) , .Z( u1_u8_X_7 ) );
  XOR2_X1 u1_u8_U33 (.B( u1_K9_24 ) , .A( u1_R7_17 ) , .Z( u1_u8_X_24 ) );
  XOR2_X1 u1_u8_U34 (.B( u1_K9_23 ) , .A( u1_R7_16 ) , .Z( u1_u8_X_23 ) );
  XOR2_X1 u1_u8_U35 (.B( u1_K9_22 ) , .A( u1_R7_15 ) , .Z( u1_u8_X_22 ) );
  XOR2_X1 u1_u8_U36 (.B( u1_K9_21 ) , .A( u1_R7_14 ) , .Z( u1_u8_X_21 ) );
  XOR2_X1 u1_u8_U37 (.B( u1_K9_20 ) , .A( u1_R7_13 ) , .Z( u1_u8_X_20 ) );
  XOR2_X1 u1_u8_U38 (.B( u1_K9_1 ) , .A( u1_R7_32 ) , .Z( u1_u8_X_1 ) );
  XOR2_X1 u1_u8_U39 (.B( u1_K9_19 ) , .A( u1_R7_12 ) , .Z( u1_u8_X_19 ) );
  XOR2_X1 u1_u8_U4 (.B( u1_K9_6 ) , .A( u1_R7_5 ) , .Z( u1_u8_X_6 ) );
  XOR2_X1 u1_u8_U40 (.B( u1_K9_18 ) , .A( u1_R7_13 ) , .Z( u1_u8_X_18 ) );
  XOR2_X1 u1_u8_U41 (.B( u1_K9_17 ) , .A( u1_R7_12 ) , .Z( u1_u8_X_17 ) );
  XOR2_X1 u1_u8_U42 (.B( u1_K9_16 ) , .A( u1_R7_11 ) , .Z( u1_u8_X_16 ) );
  XOR2_X1 u1_u8_U43 (.B( u1_K9_15 ) , .A( u1_R7_10 ) , .Z( u1_u8_X_15 ) );
  XOR2_X1 u1_u8_U44 (.B( u1_K9_14 ) , .A( u1_R7_9 ) , .Z( u1_u8_X_14 ) );
  XOR2_X1 u1_u8_U45 (.B( u1_K9_13 ) , .A( u1_R7_8 ) , .Z( u1_u8_X_13 ) );
  XOR2_X1 u1_u8_U46 (.B( u1_K9_12 ) , .A( u1_R7_9 ) , .Z( u1_u8_X_12 ) );
  XOR2_X1 u1_u8_U47 (.B( u1_K9_11 ) , .A( u1_R7_8 ) , .Z( u1_u8_X_11 ) );
  XOR2_X1 u1_u8_U48 (.B( u1_K9_10 ) , .A( u1_R7_7 ) , .Z( u1_u8_X_10 ) );
  XOR2_X1 u1_u8_U5 (.B( u1_K9_5 ) , .A( u1_R7_4 ) , .Z( u1_u8_X_5 ) );
  XOR2_X1 u1_u8_U6 (.B( u1_K9_4 ) , .A( u1_R7_3 ) , .Z( u1_u8_X_4 ) );
  AND2_X1 u1_u8_u0_U10 (.A1( u1_u8_u0_n131 ) , .ZN( u1_u8_u0_n141 ) , .A2( u1_u8_u0_n150 ) );
  AND3_X1 u1_u8_u0_U11 (.A2( u1_u8_u0_n112 ) , .ZN( u1_u8_u0_n127 ) , .A3( u1_u8_u0_n130 ) , .A1( u1_u8_u0_n148 ) );
  AND2_X1 u1_u8_u0_U12 (.ZN( u1_u8_u0_n107 ) , .A1( u1_u8_u0_n130 ) , .A2( u1_u8_u0_n140 ) );
  AND2_X1 u1_u8_u0_U13 (.A2( u1_u8_u0_n129 ) , .A1( u1_u8_u0_n130 ) , .ZN( u1_u8_u0_n151 ) );
  AND2_X1 u1_u8_u0_U14 (.A1( u1_u8_u0_n108 ) , .A2( u1_u8_u0_n125 ) , .ZN( u1_u8_u0_n145 ) );
  INV_X1 u1_u8_u0_U15 (.A( u1_u8_u0_n143 ) , .ZN( u1_u8_u0_n173 ) );
  NOR2_X1 u1_u8_u0_U16 (.A2( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n147 ) , .A1( u1_u8_u0_n160 ) );
  AOI21_X1 u1_u8_u0_U17 (.B1( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n132 ) , .A( u1_u8_u0_n165 ) , .B2( u1_u8_u0_n93 ) );
  OAI22_X1 u1_u8_u0_U18 (.B1( u1_u8_u0_n131 ) , .A1( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n147 ) , .A2( u1_u8_u0_n90 ) , .ZN( u1_u8_u0_n91 ) );
  AND3_X1 u1_u8_u0_U19 (.A3( u1_u8_u0_n121 ) , .A2( u1_u8_u0_n125 ) , .A1( u1_u8_u0_n148 ) , .ZN( u1_u8_u0_n90 ) );
  OAI22_X1 u1_u8_u0_U20 (.B1( u1_u8_u0_n125 ) , .ZN( u1_u8_u0_n126 ) , .A1( u1_u8_u0_n138 ) , .A2( u1_u8_u0_n146 ) , .B2( u1_u8_u0_n147 ) );
  NOR2_X1 u1_u8_u0_U21 (.A1( u1_u8_u0_n163 ) , .A2( u1_u8_u0_n164 ) , .ZN( u1_u8_u0_n95 ) );
  AOI22_X1 u1_u8_u0_U22 (.B2( u1_u8_u0_n109 ) , .A2( u1_u8_u0_n110 ) , .ZN( u1_u8_u0_n111 ) , .B1( u1_u8_u0_n118 ) , .A1( u1_u8_u0_n160 ) );
  NAND2_X1 u1_u8_u0_U23 (.A2( u1_u8_u0_n102 ) , .A1( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n149 ) );
  INV_X1 u1_u8_u0_U24 (.A( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n161 ) );
  INV_X1 u1_u8_u0_U25 (.A( u1_u8_u0_n118 ) , .ZN( u1_u8_u0_n158 ) );
  NAND2_X1 u1_u8_u0_U26 (.A2( u1_u8_u0_n100 ) , .ZN( u1_u8_u0_n131 ) , .A1( u1_u8_u0_n92 ) );
  NAND2_X1 u1_u8_u0_U27 (.ZN( u1_u8_u0_n108 ) , .A1( u1_u8_u0_n92 ) , .A2( u1_u8_u0_n94 ) );
  AOI21_X1 u1_u8_u0_U28 (.ZN( u1_u8_u0_n104 ) , .B1( u1_u8_u0_n107 ) , .B2( u1_u8_u0_n141 ) , .A( u1_u8_u0_n144 ) );
  AOI21_X1 u1_u8_u0_U29 (.B1( u1_u8_u0_n127 ) , .B2( u1_u8_u0_n129 ) , .A( u1_u8_u0_n138 ) , .ZN( u1_u8_u0_n96 ) );
  INV_X1 u1_u8_u0_U3 (.A( u1_u8_u0_n113 ) , .ZN( u1_u8_u0_n166 ) );
  NAND2_X1 u1_u8_u0_U30 (.A2( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n114 ) , .A1( u1_u8_u0_n92 ) );
  NOR2_X1 u1_u8_u0_U31 (.A1( u1_u8_u0_n120 ) , .ZN( u1_u8_u0_n143 ) , .A2( u1_u8_u0_n167 ) );
  OAI221_X1 u1_u8_u0_U32 (.C1( u1_u8_u0_n112 ) , .ZN( u1_u8_u0_n120 ) , .B1( u1_u8_u0_n138 ) , .B2( u1_u8_u0_n141 ) , .C2( u1_u8_u0_n147 ) , .A( u1_u8_u0_n172 ) );
  AOI211_X1 u1_u8_u0_U33 (.B( u1_u8_u0_n115 ) , .A( u1_u8_u0_n116 ) , .C2( u1_u8_u0_n117 ) , .C1( u1_u8_u0_n118 ) , .ZN( u1_u8_u0_n119 ) );
  NAND2_X1 u1_u8_u0_U34 (.A2( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n140 ) , .A1( u1_u8_u0_n94 ) );
  NAND2_X1 u1_u8_u0_U35 (.A1( u1_u8_u0_n100 ) , .A2( u1_u8_u0_n103 ) , .ZN( u1_u8_u0_n125 ) );
  NAND2_X1 u1_u8_u0_U36 (.A1( u1_u8_u0_n101 ) , .A2( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n150 ) );
  INV_X1 u1_u8_u0_U37 (.A( u1_u8_u0_n138 ) , .ZN( u1_u8_u0_n160 ) );
  NAND2_X1 u1_u8_u0_U38 (.A2( u1_u8_u0_n100 ) , .A1( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n139 ) );
  NAND2_X1 u1_u8_u0_U39 (.ZN( u1_u8_u0_n112 ) , .A2( u1_u8_u0_n92 ) , .A1( u1_u8_u0_n93 ) );
  AOI21_X1 u1_u8_u0_U4 (.B1( u1_u8_u0_n114 ) , .ZN( u1_u8_u0_n115 ) , .B2( u1_u8_u0_n129 ) , .A( u1_u8_u0_n161 ) );
  NAND2_X1 u1_u8_u0_U40 (.A1( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n130 ) , .A2( u1_u8_u0_n94 ) );
  INV_X1 u1_u8_u0_U41 (.ZN( u1_u8_u0_n172 ) , .A( u1_u8_u0_n88 ) );
  OAI222_X1 u1_u8_u0_U42 (.C1( u1_u8_u0_n108 ) , .A1( u1_u8_u0_n125 ) , .B2( u1_u8_u0_n128 ) , .B1( u1_u8_u0_n144 ) , .A2( u1_u8_u0_n158 ) , .C2( u1_u8_u0_n161 ) , .ZN( u1_u8_u0_n88 ) );
  NAND2_X1 u1_u8_u0_U43 (.A2( u1_u8_u0_n101 ) , .ZN( u1_u8_u0_n121 ) , .A1( u1_u8_u0_n93 ) );
  OR3_X1 u1_u8_u0_U44 (.A3( u1_u8_u0_n152 ) , .A2( u1_u8_u0_n153 ) , .A1( u1_u8_u0_n154 ) , .ZN( u1_u8_u0_n155 ) );
  AOI21_X1 u1_u8_u0_U45 (.A( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n145 ) , .B1( u1_u8_u0_n146 ) , .ZN( u1_u8_u0_n154 ) );
  AOI21_X1 u1_u8_u0_U46 (.B2( u1_u8_u0_n150 ) , .B1( u1_u8_u0_n151 ) , .ZN( u1_u8_u0_n152 ) , .A( u1_u8_u0_n158 ) );
  AOI21_X1 u1_u8_u0_U47 (.A( u1_u8_u0_n147 ) , .B2( u1_u8_u0_n148 ) , .B1( u1_u8_u0_n149 ) , .ZN( u1_u8_u0_n153 ) );
  INV_X1 u1_u8_u0_U48 (.ZN( u1_u8_u0_n171 ) , .A( u1_u8_u0_n99 ) );
  OAI211_X1 u1_u8_u0_U49 (.C2( u1_u8_u0_n140 ) , .C1( u1_u8_u0_n161 ) , .A( u1_u8_u0_n169 ) , .B( u1_u8_u0_n98 ) , .ZN( u1_u8_u0_n99 ) );
  AOI21_X1 u1_u8_u0_U5 (.B2( u1_u8_u0_n131 ) , .ZN( u1_u8_u0_n134 ) , .B1( u1_u8_u0_n151 ) , .A( u1_u8_u0_n158 ) );
  INV_X1 u1_u8_u0_U50 (.ZN( u1_u8_u0_n169 ) , .A( u1_u8_u0_n91 ) );
  AOI211_X1 u1_u8_u0_U51 (.C1( u1_u8_u0_n118 ) , .A( u1_u8_u0_n123 ) , .B( u1_u8_u0_n96 ) , .C2( u1_u8_u0_n97 ) , .ZN( u1_u8_u0_n98 ) );
  NOR2_X1 u1_u8_u0_U52 (.A2( u1_u8_X_4 ) , .A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n118 ) );
  NOR2_X1 u1_u8_u0_U53 (.A2( u1_u8_X_1 ) , .ZN( u1_u8_u0_n101 ) , .A1( u1_u8_u0_n163 ) );
  NOR2_X1 u1_u8_u0_U54 (.A2( u1_u8_X_3 ) , .A1( u1_u8_X_6 ) , .ZN( u1_u8_u0_n94 ) );
  NOR2_X1 u1_u8_u0_U55 (.A2( u1_u8_X_6 ) , .ZN( u1_u8_u0_n100 ) , .A1( u1_u8_u0_n162 ) );
  NAND2_X1 u1_u8_u0_U56 (.A2( u1_u8_X_4 ) , .A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n144 ) );
  NOR2_X1 u1_u8_u0_U57 (.A2( u1_u8_X_5 ) , .ZN( u1_u8_u0_n136 ) , .A1( u1_u8_u0_n159 ) );
  NAND2_X1 u1_u8_u0_U58 (.A1( u1_u8_X_5 ) , .ZN( u1_u8_u0_n138 ) , .A2( u1_u8_u0_n159 ) );
  AND2_X1 u1_u8_u0_U59 (.A2( u1_u8_X_3 ) , .A1( u1_u8_X_6 ) , .ZN( u1_u8_u0_n102 ) );
  NOR2_X1 u1_u8_u0_U6 (.A1( u1_u8_u0_n108 ) , .ZN( u1_u8_u0_n123 ) , .A2( u1_u8_u0_n158 ) );
  AND2_X1 u1_u8_u0_U60 (.A1( u1_u8_X_6 ) , .A2( u1_u8_u0_n162 ) , .ZN( u1_u8_u0_n93 ) );
  INV_X1 u1_u8_u0_U61 (.A( u1_u8_X_4 ) , .ZN( u1_u8_u0_n159 ) );
  INV_X1 u1_u8_u0_U62 (.A( u1_u8_X_1 ) , .ZN( u1_u8_u0_n164 ) );
  INV_X1 u1_u8_u0_U63 (.A( u1_u8_X_3 ) , .ZN( u1_u8_u0_n162 ) );
  INV_X1 u1_u8_u0_U64 (.A( u1_u8_u0_n126 ) , .ZN( u1_u8_u0_n168 ) );
  AOI211_X1 u1_u8_u0_U65 (.B( u1_u8_u0_n133 ) , .A( u1_u8_u0_n134 ) , .C2( u1_u8_u0_n135 ) , .C1( u1_u8_u0_n136 ) , .ZN( u1_u8_u0_n137 ) );
  OR4_X1 u1_u8_u0_U66 (.ZN( u1_out8_17 ) , .A4( u1_u8_u0_n122 ) , .A2( u1_u8_u0_n123 ) , .A1( u1_u8_u0_n124 ) , .A3( u1_u8_u0_n170 ) );
  AOI21_X1 u1_u8_u0_U67 (.B2( u1_u8_u0_n107 ) , .ZN( u1_u8_u0_n124 ) , .B1( u1_u8_u0_n128 ) , .A( u1_u8_u0_n161 ) );
  INV_X1 u1_u8_u0_U68 (.A( u1_u8_u0_n111 ) , .ZN( u1_u8_u0_n170 ) );
  OR4_X1 u1_u8_u0_U69 (.ZN( u1_out8_31 ) , .A4( u1_u8_u0_n155 ) , .A2( u1_u8_u0_n156 ) , .A1( u1_u8_u0_n157 ) , .A3( u1_u8_u0_n173 ) );
  OAI21_X1 u1_u8_u0_U7 (.B1( u1_u8_u0_n150 ) , .B2( u1_u8_u0_n158 ) , .A( u1_u8_u0_n172 ) , .ZN( u1_u8_u0_n89 ) );
  AOI21_X1 u1_u8_u0_U70 (.A( u1_u8_u0_n138 ) , .B2( u1_u8_u0_n139 ) , .B1( u1_u8_u0_n140 ) , .ZN( u1_u8_u0_n157 ) );
  AOI211_X1 u1_u8_u0_U71 (.B( u1_u8_u0_n104 ) , .A( u1_u8_u0_n105 ) , .ZN( u1_u8_u0_n106 ) , .C2( u1_u8_u0_n113 ) , .C1( u1_u8_u0_n160 ) );
  INV_X1 u1_u8_u0_U72 (.ZN( u1_u8_u0_n174 ) , .A( u1_u8_u0_n89 ) );
  AOI21_X1 u1_u8_u0_U73 (.B2( u1_u8_u0_n141 ) , .B1( u1_u8_u0_n142 ) , .ZN( u1_u8_u0_n156 ) , .A( u1_u8_u0_n161 ) );
  AOI21_X1 u1_u8_u0_U74 (.ZN( u1_u8_u0_n116 ) , .B2( u1_u8_u0_n142 ) , .A( u1_u8_u0_n144 ) , .B1( u1_u8_u0_n166 ) );
  INV_X1 u1_u8_u0_U75 (.A( u1_u8_u0_n142 ) , .ZN( u1_u8_u0_n165 ) );
  NOR2_X1 u1_u8_u0_U76 (.A2( u1_u8_X_1 ) , .A1( u1_u8_X_2 ) , .ZN( u1_u8_u0_n92 ) );
  NOR2_X1 u1_u8_u0_U77 (.A2( u1_u8_X_2 ) , .ZN( u1_u8_u0_n103 ) , .A1( u1_u8_u0_n164 ) );
  INV_X1 u1_u8_u0_U78 (.A( u1_u8_X_2 ) , .ZN( u1_u8_u0_n163 ) );
  OAI221_X1 u1_u8_u0_U79 (.C1( u1_u8_u0_n121 ) , .ZN( u1_u8_u0_n122 ) , .B2( u1_u8_u0_n127 ) , .A( u1_u8_u0_n143 ) , .B1( u1_u8_u0_n144 ) , .C2( u1_u8_u0_n147 ) );
  AND2_X1 u1_u8_u0_U8 (.A1( u1_u8_u0_n114 ) , .A2( u1_u8_u0_n121 ) , .ZN( u1_u8_u0_n146 ) );
  AOI21_X1 u1_u8_u0_U80 (.B1( u1_u8_u0_n132 ) , .ZN( u1_u8_u0_n133 ) , .A( u1_u8_u0_n144 ) , .B2( u1_u8_u0_n166 ) );
  OAI22_X1 u1_u8_u0_U81 (.ZN( u1_u8_u0_n105 ) , .A2( u1_u8_u0_n132 ) , .B1( u1_u8_u0_n146 ) , .A1( u1_u8_u0_n147 ) , .B2( u1_u8_u0_n161 ) );
  NAND2_X1 u1_u8_u0_U82 (.ZN( u1_u8_u0_n110 ) , .A2( u1_u8_u0_n132 ) , .A1( u1_u8_u0_n145 ) );
  INV_X1 u1_u8_u0_U83 (.A( u1_u8_u0_n119 ) , .ZN( u1_u8_u0_n167 ) );
  NAND2_X1 u1_u8_u0_U84 (.ZN( u1_u8_u0_n148 ) , .A1( u1_u8_u0_n93 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U85 (.A1( u1_u8_u0_n100 ) , .ZN( u1_u8_u0_n129 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U86 (.A1( u1_u8_u0_n102 ) , .ZN( u1_u8_u0_n128 ) , .A2( u1_u8_u0_n95 ) );
  NAND2_X1 u1_u8_u0_U87 (.ZN( u1_u8_u0_n142 ) , .A1( u1_u8_u0_n94 ) , .A2( u1_u8_u0_n95 ) );
  NAND3_X1 u1_u8_u0_U88 (.ZN( u1_out8_23 ) , .A3( u1_u8_u0_n137 ) , .A1( u1_u8_u0_n168 ) , .A2( u1_u8_u0_n171 ) );
  NAND3_X1 u1_u8_u0_U89 (.A3( u1_u8_u0_n127 ) , .A2( u1_u8_u0_n128 ) , .ZN( u1_u8_u0_n135 ) , .A1( u1_u8_u0_n150 ) );
  NAND2_X1 u1_u8_u0_U9 (.ZN( u1_u8_u0_n113 ) , .A1( u1_u8_u0_n139 ) , .A2( u1_u8_u0_n149 ) );
  NAND3_X1 u1_u8_u0_U90 (.ZN( u1_u8_u0_n117 ) , .A3( u1_u8_u0_n132 ) , .A2( u1_u8_u0_n139 ) , .A1( u1_u8_u0_n148 ) );
  NAND3_X1 u1_u8_u0_U91 (.ZN( u1_u8_u0_n109 ) , .A2( u1_u8_u0_n114 ) , .A3( u1_u8_u0_n140 ) , .A1( u1_u8_u0_n149 ) );
  NAND3_X1 u1_u8_u0_U92 (.ZN( u1_out8_9 ) , .A3( u1_u8_u0_n106 ) , .A2( u1_u8_u0_n171 ) , .A1( u1_u8_u0_n174 ) );
  NAND3_X1 u1_u8_u0_U93 (.A2( u1_u8_u0_n128 ) , .A1( u1_u8_u0_n132 ) , .A3( u1_u8_u0_n146 ) , .ZN( u1_u8_u0_n97 ) );
  AOI21_X1 u1_u8_u1_U10 (.B2( u1_u8_u1_n155 ) , .B1( u1_u8_u1_n156 ) , .ZN( u1_u8_u1_n157 ) , .A( u1_u8_u1_n174 ) );
  NAND3_X1 u1_u8_u1_U100 (.ZN( u1_u8_u1_n113 ) , .A1( u1_u8_u1_n120 ) , .A3( u1_u8_u1_n133 ) , .A2( u1_u8_u1_n155 ) );
  NAND2_X1 u1_u8_u1_U11 (.ZN( u1_u8_u1_n140 ) , .A2( u1_u8_u1_n150 ) , .A1( u1_u8_u1_n155 ) );
  NAND2_X1 u1_u8_u1_U12 (.A1( u1_u8_u1_n131 ) , .ZN( u1_u8_u1_n147 ) , .A2( u1_u8_u1_n153 ) );
  AOI22_X1 u1_u8_u1_U13 (.B2( u1_u8_u1_n136 ) , .A2( u1_u8_u1_n137 ) , .ZN( u1_u8_u1_n143 ) , .A1( u1_u8_u1_n171 ) , .B1( u1_u8_u1_n173 ) );
  INV_X1 u1_u8_u1_U14 (.A( u1_u8_u1_n147 ) , .ZN( u1_u8_u1_n181 ) );
  INV_X1 u1_u8_u1_U15 (.A( u1_u8_u1_n139 ) , .ZN( u1_u8_u1_n174 ) );
  INV_X1 u1_u8_u1_U16 (.A( u1_u8_u1_n112 ) , .ZN( u1_u8_u1_n171 ) );
  NAND2_X1 u1_u8_u1_U17 (.ZN( u1_u8_u1_n141 ) , .A1( u1_u8_u1_n153 ) , .A2( u1_u8_u1_n156 ) );
  AND2_X1 u1_u8_u1_U18 (.A1( u1_u8_u1_n123 ) , .ZN( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n161 ) );
  NAND2_X1 u1_u8_u1_U19 (.A2( u1_u8_u1_n115 ) , .A1( u1_u8_u1_n116 ) , .ZN( u1_u8_u1_n148 ) );
  NAND2_X1 u1_u8_u1_U20 (.A2( u1_u8_u1_n133 ) , .A1( u1_u8_u1_n135 ) , .ZN( u1_u8_u1_n159 ) );
  NAND2_X1 u1_u8_u1_U21 (.A2( u1_u8_u1_n115 ) , .A1( u1_u8_u1_n120 ) , .ZN( u1_u8_u1_n132 ) );
  INV_X1 u1_u8_u1_U22 (.A( u1_u8_u1_n154 ) , .ZN( u1_u8_u1_n178 ) );
  INV_X1 u1_u8_u1_U23 (.A( u1_u8_u1_n151 ) , .ZN( u1_u8_u1_n183 ) );
  AND2_X1 u1_u8_u1_U24 (.A1( u1_u8_u1_n129 ) , .A2( u1_u8_u1_n133 ) , .ZN( u1_u8_u1_n149 ) );
  INV_X1 u1_u8_u1_U25 (.A( u1_u8_u1_n131 ) , .ZN( u1_u8_u1_n180 ) );
  OR4_X1 u1_u8_u1_U26 (.A4( u1_u8_u1_n106 ) , .A3( u1_u8_u1_n107 ) , .ZN( u1_u8_u1_n108 ) , .A1( u1_u8_u1_n117 ) , .A2( u1_u8_u1_n184 ) );
  AOI21_X1 u1_u8_u1_U27 (.ZN( u1_u8_u1_n106 ) , .A( u1_u8_u1_n112 ) , .B1( u1_u8_u1_n154 ) , .B2( u1_u8_u1_n156 ) );
  AOI21_X1 u1_u8_u1_U28 (.ZN( u1_u8_u1_n107 ) , .B1( u1_u8_u1_n134 ) , .B2( u1_u8_u1_n149 ) , .A( u1_u8_u1_n174 ) );
  INV_X1 u1_u8_u1_U29 (.A( u1_u8_u1_n101 ) , .ZN( u1_u8_u1_n184 ) );
  INV_X1 u1_u8_u1_U3 (.A( u1_u8_u1_n159 ) , .ZN( u1_u8_u1_n182 ) );
  AOI221_X1 u1_u8_u1_U30 (.B1( u1_u8_u1_n140 ) , .ZN( u1_u8_u1_n167 ) , .B2( u1_u8_u1_n172 ) , .C2( u1_u8_u1_n175 ) , .C1( u1_u8_u1_n178 ) , .A( u1_u8_u1_n188 ) );
  INV_X1 u1_u8_u1_U31 (.ZN( u1_u8_u1_n188 ) , .A( u1_u8_u1_n97 ) );
  AOI211_X1 u1_u8_u1_U32 (.A( u1_u8_u1_n118 ) , .C1( u1_u8_u1_n132 ) , .C2( u1_u8_u1_n139 ) , .B( u1_u8_u1_n96 ) , .ZN( u1_u8_u1_n97 ) );
  AOI21_X1 u1_u8_u1_U33 (.B2( u1_u8_u1_n121 ) , .B1( u1_u8_u1_n135 ) , .A( u1_u8_u1_n152 ) , .ZN( u1_u8_u1_n96 ) );
  OAI221_X1 u1_u8_u1_U34 (.A( u1_u8_u1_n119 ) , .C2( u1_u8_u1_n129 ) , .ZN( u1_u8_u1_n138 ) , .B2( u1_u8_u1_n152 ) , .C1( u1_u8_u1_n174 ) , .B1( u1_u8_u1_n187 ) );
  INV_X1 u1_u8_u1_U35 (.A( u1_u8_u1_n148 ) , .ZN( u1_u8_u1_n187 ) );
  AOI211_X1 u1_u8_u1_U36 (.B( u1_u8_u1_n117 ) , .A( u1_u8_u1_n118 ) , .ZN( u1_u8_u1_n119 ) , .C2( u1_u8_u1_n146 ) , .C1( u1_u8_u1_n159 ) );
  NOR2_X1 u1_u8_u1_U37 (.A1( u1_u8_u1_n168 ) , .A2( u1_u8_u1_n176 ) , .ZN( u1_u8_u1_n98 ) );
  AOI211_X1 u1_u8_u1_U38 (.B( u1_u8_u1_n162 ) , .A( u1_u8_u1_n163 ) , .C2( u1_u8_u1_n164 ) , .ZN( u1_u8_u1_n165 ) , .C1( u1_u8_u1_n171 ) );
  AOI21_X1 u1_u8_u1_U39 (.A( u1_u8_u1_n160 ) , .B2( u1_u8_u1_n161 ) , .ZN( u1_u8_u1_n162 ) , .B1( u1_u8_u1_n182 ) );
  AOI221_X1 u1_u8_u1_U4 (.A( u1_u8_u1_n138 ) , .C2( u1_u8_u1_n139 ) , .C1( u1_u8_u1_n140 ) , .B2( u1_u8_u1_n141 ) , .ZN( u1_u8_u1_n142 ) , .B1( u1_u8_u1_n175 ) );
  OR2_X1 u1_u8_u1_U40 (.A2( u1_u8_u1_n157 ) , .A1( u1_u8_u1_n158 ) , .ZN( u1_u8_u1_n163 ) );
  NAND2_X1 u1_u8_u1_U41 (.A1( u1_u8_u1_n128 ) , .ZN( u1_u8_u1_n146 ) , .A2( u1_u8_u1_n160 ) );
  NAND2_X1 u1_u8_u1_U42 (.A2( u1_u8_u1_n112 ) , .ZN( u1_u8_u1_n139 ) , .A1( u1_u8_u1_n152 ) );
  NAND2_X1 u1_u8_u1_U43 (.A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n156 ) , .A2( u1_u8_u1_n99 ) );
  NOR2_X1 u1_u8_u1_U44 (.ZN( u1_u8_u1_n117 ) , .A1( u1_u8_u1_n121 ) , .A2( u1_u8_u1_n160 ) );
  OAI21_X1 u1_u8_u1_U45 (.B2( u1_u8_u1_n123 ) , .ZN( u1_u8_u1_n145 ) , .B1( u1_u8_u1_n160 ) , .A( u1_u8_u1_n185 ) );
  INV_X1 u1_u8_u1_U46 (.A( u1_u8_u1_n122 ) , .ZN( u1_u8_u1_n185 ) );
  AOI21_X1 u1_u8_u1_U47 (.B2( u1_u8_u1_n120 ) , .B1( u1_u8_u1_n121 ) , .ZN( u1_u8_u1_n122 ) , .A( u1_u8_u1_n128 ) );
  AOI21_X1 u1_u8_u1_U48 (.A( u1_u8_u1_n128 ) , .B2( u1_u8_u1_n129 ) , .ZN( u1_u8_u1_n130 ) , .B1( u1_u8_u1_n150 ) );
  NAND2_X1 u1_u8_u1_U49 (.ZN( u1_u8_u1_n112 ) , .A1( u1_u8_u1_n169 ) , .A2( u1_u8_u1_n170 ) );
  AOI211_X1 u1_u8_u1_U5 (.ZN( u1_u8_u1_n124 ) , .A( u1_u8_u1_n138 ) , .C2( u1_u8_u1_n139 ) , .B( u1_u8_u1_n145 ) , .C1( u1_u8_u1_n147 ) );
  NAND2_X1 u1_u8_u1_U50 (.ZN( u1_u8_u1_n129 ) , .A2( u1_u8_u1_n95 ) , .A1( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U51 (.A1( u1_u8_u1_n102 ) , .ZN( u1_u8_u1_n154 ) , .A2( u1_u8_u1_n99 ) );
  NAND2_X1 u1_u8_u1_U52 (.A2( u1_u8_u1_n100 ) , .ZN( u1_u8_u1_n135 ) , .A1( u1_u8_u1_n99 ) );
  AOI21_X1 u1_u8_u1_U53 (.A( u1_u8_u1_n152 ) , .B2( u1_u8_u1_n153 ) , .B1( u1_u8_u1_n154 ) , .ZN( u1_u8_u1_n158 ) );
  INV_X1 u1_u8_u1_U54 (.A( u1_u8_u1_n160 ) , .ZN( u1_u8_u1_n175 ) );
  NAND2_X1 u1_u8_u1_U55 (.A1( u1_u8_u1_n100 ) , .ZN( u1_u8_u1_n116 ) , .A2( u1_u8_u1_n95 ) );
  NAND2_X1 u1_u8_u1_U56 (.A1( u1_u8_u1_n102 ) , .ZN( u1_u8_u1_n131 ) , .A2( u1_u8_u1_n95 ) );
  NAND2_X1 u1_u8_u1_U57 (.A2( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n121 ) , .A1( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U58 (.A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n153 ) , .A2( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U59 (.A2( u1_u8_u1_n104 ) , .A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n133 ) );
  AOI22_X1 u1_u8_u1_U6 (.B2( u1_u8_u1_n113 ) , .A2( u1_u8_u1_n114 ) , .ZN( u1_u8_u1_n125 ) , .A1( u1_u8_u1_n171 ) , .B1( u1_u8_u1_n173 ) );
  NAND2_X1 u1_u8_u1_U60 (.ZN( u1_u8_u1_n150 ) , .A2( u1_u8_u1_n98 ) , .A1( u1_u8_u1_n99 ) );
  NAND2_X1 u1_u8_u1_U61 (.A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n155 ) , .A2( u1_u8_u1_n95 ) );
  OAI21_X1 u1_u8_u1_U62 (.ZN( u1_u8_u1_n109 ) , .B1( u1_u8_u1_n129 ) , .B2( u1_u8_u1_n160 ) , .A( u1_u8_u1_n167 ) );
  NAND2_X1 u1_u8_u1_U63 (.A2( u1_u8_u1_n100 ) , .A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n120 ) );
  NAND2_X1 u1_u8_u1_U64 (.A1( u1_u8_u1_n102 ) , .A2( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n115 ) );
  NAND2_X1 u1_u8_u1_U65 (.A2( u1_u8_u1_n100 ) , .A1( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n151 ) );
  NAND2_X1 u1_u8_u1_U66 (.A2( u1_u8_u1_n103 ) , .A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n161 ) );
  INV_X1 u1_u8_u1_U67 (.A( u1_u8_u1_n152 ) , .ZN( u1_u8_u1_n173 ) );
  INV_X1 u1_u8_u1_U68 (.A( u1_u8_u1_n128 ) , .ZN( u1_u8_u1_n172 ) );
  NAND2_X1 u1_u8_u1_U69 (.A2( u1_u8_u1_n102 ) , .A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n123 ) );
  NAND2_X1 u1_u8_u1_U7 (.ZN( u1_u8_u1_n114 ) , .A1( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n156 ) );
  NOR2_X1 u1_u8_u1_U70 (.A2( u1_u8_X_7 ) , .A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n95 ) );
  NOR2_X1 u1_u8_u1_U71 (.A1( u1_u8_X_12 ) , .A2( u1_u8_X_9 ) , .ZN( u1_u8_u1_n100 ) );
  NOR2_X1 u1_u8_u1_U72 (.A2( u1_u8_X_8 ) , .A1( u1_u8_u1_n177 ) , .ZN( u1_u8_u1_n99 ) );
  NOR2_X1 u1_u8_u1_U73 (.A2( u1_u8_X_12 ) , .ZN( u1_u8_u1_n102 ) , .A1( u1_u8_u1_n176 ) );
  NOR2_X1 u1_u8_u1_U74 (.A2( u1_u8_X_9 ) , .ZN( u1_u8_u1_n105 ) , .A1( u1_u8_u1_n168 ) );
  NAND2_X1 u1_u8_u1_U75 (.A1( u1_u8_X_10 ) , .ZN( u1_u8_u1_n160 ) , .A2( u1_u8_u1_n169 ) );
  NAND2_X1 u1_u8_u1_U76 (.A2( u1_u8_X_10 ) , .A1( u1_u8_X_11 ) , .ZN( u1_u8_u1_n152 ) );
  NAND2_X1 u1_u8_u1_U77 (.A1( u1_u8_X_11 ) , .ZN( u1_u8_u1_n128 ) , .A2( u1_u8_u1_n170 ) );
  AND2_X1 u1_u8_u1_U78 (.A2( u1_u8_X_7 ) , .A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n104 ) );
  AND2_X1 u1_u8_u1_U79 (.A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n103 ) , .A2( u1_u8_u1_n177 ) );
  NOR2_X1 u1_u8_u1_U8 (.A1( u1_u8_u1_n112 ) , .A2( u1_u8_u1_n116 ) , .ZN( u1_u8_u1_n118 ) );
  INV_X1 u1_u8_u1_U80 (.A( u1_u8_X_10 ) , .ZN( u1_u8_u1_n170 ) );
  INV_X1 u1_u8_u1_U81 (.A( u1_u8_X_9 ) , .ZN( u1_u8_u1_n176 ) );
  INV_X1 u1_u8_u1_U82 (.A( u1_u8_X_11 ) , .ZN( u1_u8_u1_n169 ) );
  INV_X1 u1_u8_u1_U83 (.A( u1_u8_X_12 ) , .ZN( u1_u8_u1_n168 ) );
  INV_X1 u1_u8_u1_U84 (.A( u1_u8_X_7 ) , .ZN( u1_u8_u1_n177 ) );
  NAND4_X1 u1_u8_u1_U85 (.ZN( u1_out8_28 ) , .A4( u1_u8_u1_n124 ) , .A3( u1_u8_u1_n125 ) , .A2( u1_u8_u1_n126 ) , .A1( u1_u8_u1_n127 ) );
  OAI21_X1 u1_u8_u1_U86 (.ZN( u1_u8_u1_n127 ) , .B2( u1_u8_u1_n139 ) , .B1( u1_u8_u1_n175 ) , .A( u1_u8_u1_n183 ) );
  OAI21_X1 u1_u8_u1_U87 (.ZN( u1_u8_u1_n126 ) , .B2( u1_u8_u1_n140 ) , .A( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n178 ) );
  NAND4_X1 u1_u8_u1_U88 (.ZN( u1_out8_18 ) , .A4( u1_u8_u1_n165 ) , .A3( u1_u8_u1_n166 ) , .A1( u1_u8_u1_n167 ) , .A2( u1_u8_u1_n186 ) );
  AOI22_X1 u1_u8_u1_U89 (.B2( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n147 ) , .A2( u1_u8_u1_n148 ) , .ZN( u1_u8_u1_n166 ) , .A1( u1_u8_u1_n172 ) );
  OAI21_X1 u1_u8_u1_U9 (.ZN( u1_u8_u1_n101 ) , .B1( u1_u8_u1_n141 ) , .A( u1_u8_u1_n146 ) , .B2( u1_u8_u1_n183 ) );
  INV_X1 u1_u8_u1_U90 (.A( u1_u8_u1_n145 ) , .ZN( u1_u8_u1_n186 ) );
  NAND4_X1 u1_u8_u1_U91 (.ZN( u1_out8_2 ) , .A4( u1_u8_u1_n142 ) , .A3( u1_u8_u1_n143 ) , .A2( u1_u8_u1_n144 ) , .A1( u1_u8_u1_n179 ) );
  OAI21_X1 u1_u8_u1_U92 (.B2( u1_u8_u1_n132 ) , .ZN( u1_u8_u1_n144 ) , .A( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n180 ) );
  INV_X1 u1_u8_u1_U93 (.A( u1_u8_u1_n130 ) , .ZN( u1_u8_u1_n179 ) );
  OR4_X1 u1_u8_u1_U94 (.ZN( u1_out8_13 ) , .A4( u1_u8_u1_n108 ) , .A3( u1_u8_u1_n109 ) , .A2( u1_u8_u1_n110 ) , .A1( u1_u8_u1_n111 ) );
  AOI21_X1 u1_u8_u1_U95 (.ZN( u1_u8_u1_n111 ) , .A( u1_u8_u1_n128 ) , .B2( u1_u8_u1_n131 ) , .B1( u1_u8_u1_n135 ) );
  AOI21_X1 u1_u8_u1_U96 (.ZN( u1_u8_u1_n110 ) , .A( u1_u8_u1_n116 ) , .B1( u1_u8_u1_n152 ) , .B2( u1_u8_u1_n160 ) );
  NAND3_X1 u1_u8_u1_U97 (.A3( u1_u8_u1_n149 ) , .A2( u1_u8_u1_n150 ) , .A1( u1_u8_u1_n151 ) , .ZN( u1_u8_u1_n164 ) );
  NAND3_X1 u1_u8_u1_U98 (.A3( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n135 ) , .ZN( u1_u8_u1_n136 ) , .A1( u1_u8_u1_n151 ) );
  NAND3_X1 u1_u8_u1_U99 (.A1( u1_u8_u1_n133 ) , .ZN( u1_u8_u1_n137 ) , .A2( u1_u8_u1_n154 ) , .A3( u1_u8_u1_n181 ) );
  OAI22_X1 u1_u8_u2_U10 (.B1( u1_u8_u2_n151 ) , .A2( u1_u8_u2_n152 ) , .A1( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n160 ) , .B2( u1_u8_u2_n168 ) );
  NAND3_X1 u1_u8_u2_U100 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n104 ) , .A3( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n98 ) );
  NOR3_X1 u1_u8_u2_U11 (.A1( u1_u8_u2_n150 ) , .ZN( u1_u8_u2_n151 ) , .A3( u1_u8_u2_n175 ) , .A2( u1_u8_u2_n188 ) );
  AOI21_X1 u1_u8_u2_U12 (.B2( u1_u8_u2_n123 ) , .ZN( u1_u8_u2_n125 ) , .A( u1_u8_u2_n171 ) , .B1( u1_u8_u2_n184 ) );
  INV_X1 u1_u8_u2_U13 (.A( u1_u8_u2_n150 ) , .ZN( u1_u8_u2_n184 ) );
  AOI21_X1 u1_u8_u2_U14 (.ZN( u1_u8_u2_n144 ) , .B2( u1_u8_u2_n155 ) , .A( u1_u8_u2_n172 ) , .B1( u1_u8_u2_n185 ) );
  AOI21_X1 u1_u8_u2_U15 (.B2( u1_u8_u2_n143 ) , .ZN( u1_u8_u2_n145 ) , .B1( u1_u8_u2_n152 ) , .A( u1_u8_u2_n171 ) );
  INV_X1 u1_u8_u2_U16 (.A( u1_u8_u2_n156 ) , .ZN( u1_u8_u2_n171 ) );
  INV_X1 u1_u8_u2_U17 (.A( u1_u8_u2_n120 ) , .ZN( u1_u8_u2_n188 ) );
  NAND2_X1 u1_u8_u2_U18 (.A2( u1_u8_u2_n122 ) , .ZN( u1_u8_u2_n150 ) , .A1( u1_u8_u2_n152 ) );
  INV_X1 u1_u8_u2_U19 (.A( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n170 ) );
  INV_X1 u1_u8_u2_U20 (.A( u1_u8_u2_n137 ) , .ZN( u1_u8_u2_n173 ) );
  NAND2_X1 u1_u8_u2_U21 (.A1( u1_u8_u2_n132 ) , .A2( u1_u8_u2_n139 ) , .ZN( u1_u8_u2_n157 ) );
  INV_X1 u1_u8_u2_U22 (.A( u1_u8_u2_n113 ) , .ZN( u1_u8_u2_n178 ) );
  INV_X1 u1_u8_u2_U23 (.A( u1_u8_u2_n139 ) , .ZN( u1_u8_u2_n175 ) );
  INV_X1 u1_u8_u2_U24 (.A( u1_u8_u2_n155 ) , .ZN( u1_u8_u2_n181 ) );
  INV_X1 u1_u8_u2_U25 (.A( u1_u8_u2_n119 ) , .ZN( u1_u8_u2_n177 ) );
  INV_X1 u1_u8_u2_U26 (.A( u1_u8_u2_n116 ) , .ZN( u1_u8_u2_n180 ) );
  INV_X1 u1_u8_u2_U27 (.A( u1_u8_u2_n131 ) , .ZN( u1_u8_u2_n179 ) );
  INV_X1 u1_u8_u2_U28 (.A( u1_u8_u2_n154 ) , .ZN( u1_u8_u2_n176 ) );
  NAND2_X1 u1_u8_u2_U29 (.A2( u1_u8_u2_n116 ) , .A1( u1_u8_u2_n117 ) , .ZN( u1_u8_u2_n118 ) );
  NOR2_X1 u1_u8_u2_U3 (.ZN( u1_u8_u2_n121 ) , .A2( u1_u8_u2_n177 ) , .A1( u1_u8_u2_n180 ) );
  INV_X1 u1_u8_u2_U30 (.A( u1_u8_u2_n132 ) , .ZN( u1_u8_u2_n182 ) );
  INV_X1 u1_u8_u2_U31 (.A( u1_u8_u2_n158 ) , .ZN( u1_u8_u2_n183 ) );
  OAI21_X1 u1_u8_u2_U32 (.A( u1_u8_u2_n156 ) , .B1( u1_u8_u2_n157 ) , .ZN( u1_u8_u2_n158 ) , .B2( u1_u8_u2_n179 ) );
  NOR2_X1 u1_u8_u2_U33 (.ZN( u1_u8_u2_n156 ) , .A1( u1_u8_u2_n166 ) , .A2( u1_u8_u2_n169 ) );
  NOR2_X1 u1_u8_u2_U34 (.A2( u1_u8_u2_n114 ) , .ZN( u1_u8_u2_n137 ) , .A1( u1_u8_u2_n140 ) );
  NOR2_X1 u1_u8_u2_U35 (.A2( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n153 ) , .A1( u1_u8_u2_n156 ) );
  AOI211_X1 u1_u8_u2_U36 (.ZN( u1_u8_u2_n130 ) , .C1( u1_u8_u2_n138 ) , .C2( u1_u8_u2_n179 ) , .B( u1_u8_u2_n96 ) , .A( u1_u8_u2_n97 ) );
  OAI22_X1 u1_u8_u2_U37 (.B1( u1_u8_u2_n133 ) , .A2( u1_u8_u2_n137 ) , .A1( u1_u8_u2_n152 ) , .B2( u1_u8_u2_n168 ) , .ZN( u1_u8_u2_n97 ) );
  OAI221_X1 u1_u8_u2_U38 (.B1( u1_u8_u2_n113 ) , .C1( u1_u8_u2_n132 ) , .A( u1_u8_u2_n149 ) , .B2( u1_u8_u2_n171 ) , .C2( u1_u8_u2_n172 ) , .ZN( u1_u8_u2_n96 ) );
  OAI221_X1 u1_u8_u2_U39 (.A( u1_u8_u2_n115 ) , .C2( u1_u8_u2_n123 ) , .B2( u1_u8_u2_n143 ) , .B1( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n163 ) , .C1( u1_u8_u2_n168 ) );
  INV_X1 u1_u8_u2_U4 (.A( u1_u8_u2_n134 ) , .ZN( u1_u8_u2_n185 ) );
  OAI21_X1 u1_u8_u2_U40 (.A( u1_u8_u2_n114 ) , .ZN( u1_u8_u2_n115 ) , .B1( u1_u8_u2_n176 ) , .B2( u1_u8_u2_n178 ) );
  OAI221_X1 u1_u8_u2_U41 (.A( u1_u8_u2_n135 ) , .B2( u1_u8_u2_n136 ) , .B1( u1_u8_u2_n137 ) , .ZN( u1_u8_u2_n162 ) , .C2( u1_u8_u2_n167 ) , .C1( u1_u8_u2_n185 ) );
  AND3_X1 u1_u8_u2_U42 (.A3( u1_u8_u2_n131 ) , .A2( u1_u8_u2_n132 ) , .A1( u1_u8_u2_n133 ) , .ZN( u1_u8_u2_n136 ) );
  AOI22_X1 u1_u8_u2_U43 (.ZN( u1_u8_u2_n135 ) , .B1( u1_u8_u2_n140 ) , .A1( u1_u8_u2_n156 ) , .B2( u1_u8_u2_n180 ) , .A2( u1_u8_u2_n188 ) );
  AOI21_X1 u1_u8_u2_U44 (.ZN( u1_u8_u2_n149 ) , .B1( u1_u8_u2_n173 ) , .B2( u1_u8_u2_n188 ) , .A( u1_u8_u2_n95 ) );
  AND3_X1 u1_u8_u2_U45 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n104 ) , .A3( u1_u8_u2_n156 ) , .ZN( u1_u8_u2_n95 ) );
  OAI21_X1 u1_u8_u2_U46 (.A( u1_u8_u2_n101 ) , .B2( u1_u8_u2_n121 ) , .B1( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n164 ) );
  NAND2_X1 u1_u8_u2_U47 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n107 ) , .ZN( u1_u8_u2_n155 ) );
  NAND2_X1 u1_u8_u2_U48 (.A2( u1_u8_u2_n105 ) , .A1( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n143 ) );
  NAND2_X1 u1_u8_u2_U49 (.A1( u1_u8_u2_n104 ) , .A2( u1_u8_u2_n106 ) , .ZN( u1_u8_u2_n152 ) );
  NOR4_X1 u1_u8_u2_U5 (.A4( u1_u8_u2_n124 ) , .A3( u1_u8_u2_n125 ) , .A2( u1_u8_u2_n126 ) , .A1( u1_u8_u2_n127 ) , .ZN( u1_u8_u2_n128 ) );
  NAND2_X1 u1_u8_u2_U50 (.A1( u1_u8_u2_n100 ) , .A2( u1_u8_u2_n105 ) , .ZN( u1_u8_u2_n132 ) );
  INV_X1 u1_u8_u2_U51 (.A( u1_u8_u2_n140 ) , .ZN( u1_u8_u2_n168 ) );
  INV_X1 u1_u8_u2_U52 (.A( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n167 ) );
  OAI21_X1 u1_u8_u2_U53 (.A( u1_u8_u2_n141 ) , .B2( u1_u8_u2_n142 ) , .ZN( u1_u8_u2_n146 ) , .B1( u1_u8_u2_n153 ) );
  OAI21_X1 u1_u8_u2_U54 (.A( u1_u8_u2_n140 ) , .ZN( u1_u8_u2_n141 ) , .B1( u1_u8_u2_n176 ) , .B2( u1_u8_u2_n177 ) );
  NOR3_X1 u1_u8_u2_U55 (.ZN( u1_u8_u2_n142 ) , .A3( u1_u8_u2_n175 ) , .A2( u1_u8_u2_n178 ) , .A1( u1_u8_u2_n181 ) );
  NAND2_X1 u1_u8_u2_U56 (.A1( u1_u8_u2_n102 ) , .A2( u1_u8_u2_n106 ) , .ZN( u1_u8_u2_n113 ) );
  NAND2_X1 u1_u8_u2_U57 (.A1( u1_u8_u2_n106 ) , .A2( u1_u8_u2_n107 ) , .ZN( u1_u8_u2_n131 ) );
  NAND2_X1 u1_u8_u2_U58 (.A1( u1_u8_u2_n103 ) , .A2( u1_u8_u2_n107 ) , .ZN( u1_u8_u2_n139 ) );
  NAND2_X1 u1_u8_u2_U59 (.A1( u1_u8_u2_n103 ) , .A2( u1_u8_u2_n105 ) , .ZN( u1_u8_u2_n133 ) );
  AOI21_X1 u1_u8_u2_U6 (.B2( u1_u8_u2_n119 ) , .ZN( u1_u8_u2_n127 ) , .A( u1_u8_u2_n137 ) , .B1( u1_u8_u2_n155 ) );
  NAND2_X1 u1_u8_u2_U60 (.A1( u1_u8_u2_n102 ) , .A2( u1_u8_u2_n103 ) , .ZN( u1_u8_u2_n154 ) );
  NAND2_X1 u1_u8_u2_U61 (.A2( u1_u8_u2_n103 ) , .A1( u1_u8_u2_n104 ) , .ZN( u1_u8_u2_n119 ) );
  NAND2_X1 u1_u8_u2_U62 (.A2( u1_u8_u2_n107 ) , .A1( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n123 ) );
  NAND2_X1 u1_u8_u2_U63 (.A1( u1_u8_u2_n104 ) , .A2( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n122 ) );
  INV_X1 u1_u8_u2_U64 (.A( u1_u8_u2_n114 ) , .ZN( u1_u8_u2_n172 ) );
  NAND2_X1 u1_u8_u2_U65 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n102 ) , .ZN( u1_u8_u2_n116 ) );
  NAND2_X1 u1_u8_u2_U66 (.A1( u1_u8_u2_n102 ) , .A2( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n120 ) );
  NAND2_X1 u1_u8_u2_U67 (.A2( u1_u8_u2_n105 ) , .A1( u1_u8_u2_n106 ) , .ZN( u1_u8_u2_n117 ) );
  INV_X1 u1_u8_u2_U68 (.ZN( u1_u8_u2_n187 ) , .A( u1_u8_u2_n99 ) );
  OAI21_X1 u1_u8_u2_U69 (.B1( u1_u8_u2_n137 ) , .B2( u1_u8_u2_n143 ) , .A( u1_u8_u2_n98 ) , .ZN( u1_u8_u2_n99 ) );
  AOI21_X1 u1_u8_u2_U7 (.ZN( u1_u8_u2_n124 ) , .B1( u1_u8_u2_n131 ) , .B2( u1_u8_u2_n143 ) , .A( u1_u8_u2_n172 ) );
  NOR2_X1 u1_u8_u2_U70 (.A2( u1_u8_X_16 ) , .ZN( u1_u8_u2_n140 ) , .A1( u1_u8_u2_n166 ) );
  NOR2_X1 u1_u8_u2_U71 (.A2( u1_u8_X_13 ) , .A1( u1_u8_X_14 ) , .ZN( u1_u8_u2_n100 ) );
  NOR2_X1 u1_u8_u2_U72 (.A2( u1_u8_X_16 ) , .A1( u1_u8_X_17 ) , .ZN( u1_u8_u2_n138 ) );
  NOR2_X1 u1_u8_u2_U73 (.A2( u1_u8_X_15 ) , .A1( u1_u8_X_18 ) , .ZN( u1_u8_u2_n104 ) );
  NOR2_X1 u1_u8_u2_U74 (.A2( u1_u8_X_14 ) , .ZN( u1_u8_u2_n103 ) , .A1( u1_u8_u2_n174 ) );
  NOR2_X1 u1_u8_u2_U75 (.A2( u1_u8_X_15 ) , .ZN( u1_u8_u2_n102 ) , .A1( u1_u8_u2_n165 ) );
  NOR2_X1 u1_u8_u2_U76 (.A2( u1_u8_X_17 ) , .ZN( u1_u8_u2_n114 ) , .A1( u1_u8_u2_n169 ) );
  AND2_X1 u1_u8_u2_U77 (.A1( u1_u8_X_15 ) , .ZN( u1_u8_u2_n105 ) , .A2( u1_u8_u2_n165 ) );
  AND2_X1 u1_u8_u2_U78 (.A2( u1_u8_X_15 ) , .A1( u1_u8_X_18 ) , .ZN( u1_u8_u2_n107 ) );
  AND2_X1 u1_u8_u2_U79 (.A1( u1_u8_X_14 ) , .ZN( u1_u8_u2_n106 ) , .A2( u1_u8_u2_n174 ) );
  AOI21_X1 u1_u8_u2_U8 (.B2( u1_u8_u2_n120 ) , .B1( u1_u8_u2_n121 ) , .ZN( u1_u8_u2_n126 ) , .A( u1_u8_u2_n167 ) );
  AND2_X1 u1_u8_u2_U80 (.A1( u1_u8_X_13 ) , .A2( u1_u8_X_14 ) , .ZN( u1_u8_u2_n108 ) );
  INV_X1 u1_u8_u2_U81 (.A( u1_u8_X_16 ) , .ZN( u1_u8_u2_n169 ) );
  INV_X1 u1_u8_u2_U82 (.A( u1_u8_X_17 ) , .ZN( u1_u8_u2_n166 ) );
  INV_X1 u1_u8_u2_U83 (.A( u1_u8_X_13 ) , .ZN( u1_u8_u2_n174 ) );
  INV_X1 u1_u8_u2_U84 (.A( u1_u8_X_18 ) , .ZN( u1_u8_u2_n165 ) );
  NAND4_X1 u1_u8_u2_U85 (.ZN( u1_out8_30 ) , .A4( u1_u8_u2_n147 ) , .A3( u1_u8_u2_n148 ) , .A2( u1_u8_u2_n149 ) , .A1( u1_u8_u2_n187 ) );
  NOR3_X1 u1_u8_u2_U86 (.A3( u1_u8_u2_n144 ) , .A2( u1_u8_u2_n145 ) , .A1( u1_u8_u2_n146 ) , .ZN( u1_u8_u2_n147 ) );
  AOI21_X1 u1_u8_u2_U87 (.B2( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n148 ) , .A( u1_u8_u2_n162 ) , .B1( u1_u8_u2_n182 ) );
  NAND4_X1 u1_u8_u2_U88 (.ZN( u1_out8_24 ) , .A4( u1_u8_u2_n111 ) , .A3( u1_u8_u2_n112 ) , .A1( u1_u8_u2_n130 ) , .A2( u1_u8_u2_n187 ) );
  AOI221_X1 u1_u8_u2_U89 (.A( u1_u8_u2_n109 ) , .B1( u1_u8_u2_n110 ) , .ZN( u1_u8_u2_n111 ) , .C1( u1_u8_u2_n134 ) , .C2( u1_u8_u2_n170 ) , .B2( u1_u8_u2_n173 ) );
  OAI22_X1 u1_u8_u2_U9 (.ZN( u1_u8_u2_n109 ) , .A2( u1_u8_u2_n113 ) , .B2( u1_u8_u2_n133 ) , .B1( u1_u8_u2_n167 ) , .A1( u1_u8_u2_n168 ) );
  AOI21_X1 u1_u8_u2_U90 (.ZN( u1_u8_u2_n112 ) , .B2( u1_u8_u2_n156 ) , .A( u1_u8_u2_n164 ) , .B1( u1_u8_u2_n181 ) );
  NAND4_X1 u1_u8_u2_U91 (.ZN( u1_out8_16 ) , .A4( u1_u8_u2_n128 ) , .A3( u1_u8_u2_n129 ) , .A1( u1_u8_u2_n130 ) , .A2( u1_u8_u2_n186 ) );
  AOI22_X1 u1_u8_u2_U92 (.A2( u1_u8_u2_n118 ) , .ZN( u1_u8_u2_n129 ) , .A1( u1_u8_u2_n140 ) , .B1( u1_u8_u2_n157 ) , .B2( u1_u8_u2_n170 ) );
  INV_X1 u1_u8_u2_U93 (.A( u1_u8_u2_n163 ) , .ZN( u1_u8_u2_n186 ) );
  OR4_X1 u1_u8_u2_U94 (.ZN( u1_out8_6 ) , .A4( u1_u8_u2_n161 ) , .A3( u1_u8_u2_n162 ) , .A2( u1_u8_u2_n163 ) , .A1( u1_u8_u2_n164 ) );
  OR3_X1 u1_u8_u2_U95 (.A2( u1_u8_u2_n159 ) , .A1( u1_u8_u2_n160 ) , .ZN( u1_u8_u2_n161 ) , .A3( u1_u8_u2_n183 ) );
  AOI21_X1 u1_u8_u2_U96 (.B2( u1_u8_u2_n154 ) , .B1( u1_u8_u2_n155 ) , .ZN( u1_u8_u2_n159 ) , .A( u1_u8_u2_n167 ) );
  NAND3_X1 u1_u8_u2_U97 (.A2( u1_u8_u2_n117 ) , .A1( u1_u8_u2_n122 ) , .A3( u1_u8_u2_n123 ) , .ZN( u1_u8_u2_n134 ) );
  NAND3_X1 u1_u8_u2_U98 (.ZN( u1_u8_u2_n110 ) , .A2( u1_u8_u2_n131 ) , .A3( u1_u8_u2_n139 ) , .A1( u1_u8_u2_n154 ) );
  NAND3_X1 u1_u8_u2_U99 (.A2( u1_u8_u2_n100 ) , .ZN( u1_u8_u2_n101 ) , .A1( u1_u8_u2_n104 ) , .A3( u1_u8_u2_n114 ) );
  OAI22_X1 u1_u8_u3_U10 (.B1( u1_u8_u3_n113 ) , .A2( u1_u8_u3_n135 ) , .A1( u1_u8_u3_n150 ) , .B2( u1_u8_u3_n164 ) , .ZN( u1_u8_u3_n98 ) );
  OAI211_X1 u1_u8_u3_U11 (.B( u1_u8_u3_n106 ) , .ZN( u1_u8_u3_n119 ) , .C2( u1_u8_u3_n128 ) , .C1( u1_u8_u3_n167 ) , .A( u1_u8_u3_n181 ) );
  AOI221_X1 u1_u8_u3_U12 (.C1( u1_u8_u3_n105 ) , .ZN( u1_u8_u3_n106 ) , .A( u1_u8_u3_n131 ) , .B2( u1_u8_u3_n132 ) , .C2( u1_u8_u3_n133 ) , .B1( u1_u8_u3_n169 ) );
  INV_X1 u1_u8_u3_U13 (.ZN( u1_u8_u3_n181 ) , .A( u1_u8_u3_n98 ) );
  NAND2_X1 u1_u8_u3_U14 (.ZN( u1_u8_u3_n105 ) , .A2( u1_u8_u3_n130 ) , .A1( u1_u8_u3_n155 ) );
  AOI22_X1 u1_u8_u3_U15 (.B1( u1_u8_u3_n115 ) , .A2( u1_u8_u3_n116 ) , .ZN( u1_u8_u3_n123 ) , .B2( u1_u8_u3_n133 ) , .A1( u1_u8_u3_n169 ) );
  NAND2_X1 u1_u8_u3_U16 (.ZN( u1_u8_u3_n116 ) , .A2( u1_u8_u3_n151 ) , .A1( u1_u8_u3_n182 ) );
  NOR2_X1 u1_u8_u3_U17 (.ZN( u1_u8_u3_n126 ) , .A2( u1_u8_u3_n150 ) , .A1( u1_u8_u3_n164 ) );
  AOI21_X1 u1_u8_u3_U18 (.ZN( u1_u8_u3_n112 ) , .B2( u1_u8_u3_n146 ) , .B1( u1_u8_u3_n155 ) , .A( u1_u8_u3_n167 ) );
  NAND2_X1 u1_u8_u3_U19 (.A1( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n142 ) , .A2( u1_u8_u3_n164 ) );
  NAND2_X1 u1_u8_u3_U20 (.ZN( u1_u8_u3_n132 ) , .A2( u1_u8_u3_n152 ) , .A1( u1_u8_u3_n156 ) );
  AND2_X1 u1_u8_u3_U21 (.A2( u1_u8_u3_n113 ) , .A1( u1_u8_u3_n114 ) , .ZN( u1_u8_u3_n151 ) );
  INV_X1 u1_u8_u3_U22 (.A( u1_u8_u3_n133 ) , .ZN( u1_u8_u3_n165 ) );
  INV_X1 u1_u8_u3_U23 (.A( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n170 ) );
  NAND2_X1 u1_u8_u3_U24 (.A1( u1_u8_u3_n107 ) , .A2( u1_u8_u3_n108 ) , .ZN( u1_u8_u3_n140 ) );
  NAND2_X1 u1_u8_u3_U25 (.ZN( u1_u8_u3_n117 ) , .A1( u1_u8_u3_n124 ) , .A2( u1_u8_u3_n148 ) );
  NAND2_X1 u1_u8_u3_U26 (.ZN( u1_u8_u3_n143 ) , .A1( u1_u8_u3_n165 ) , .A2( u1_u8_u3_n167 ) );
  INV_X1 u1_u8_u3_U27 (.A( u1_u8_u3_n130 ) , .ZN( u1_u8_u3_n177 ) );
  INV_X1 u1_u8_u3_U28 (.A( u1_u8_u3_n128 ) , .ZN( u1_u8_u3_n176 ) );
  INV_X1 u1_u8_u3_U29 (.A( u1_u8_u3_n155 ) , .ZN( u1_u8_u3_n174 ) );
  INV_X1 u1_u8_u3_U3 (.A( u1_u8_u3_n129 ) , .ZN( u1_u8_u3_n183 ) );
  INV_X1 u1_u8_u3_U30 (.A( u1_u8_u3_n139 ) , .ZN( u1_u8_u3_n185 ) );
  NOR2_X1 u1_u8_u3_U31 (.ZN( u1_u8_u3_n135 ) , .A2( u1_u8_u3_n141 ) , .A1( u1_u8_u3_n169 ) );
  OAI222_X1 u1_u8_u3_U32 (.C2( u1_u8_u3_n107 ) , .A2( u1_u8_u3_n108 ) , .B1( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n138 ) , .B2( u1_u8_u3_n146 ) , .C1( u1_u8_u3_n154 ) , .A1( u1_u8_u3_n164 ) );
  NOR4_X1 u1_u8_u3_U33 (.A4( u1_u8_u3_n157 ) , .A3( u1_u8_u3_n158 ) , .A2( u1_u8_u3_n159 ) , .A1( u1_u8_u3_n160 ) , .ZN( u1_u8_u3_n161 ) );
  AOI21_X1 u1_u8_u3_U34 (.B2( u1_u8_u3_n152 ) , .B1( u1_u8_u3_n153 ) , .ZN( u1_u8_u3_n158 ) , .A( u1_u8_u3_n164 ) );
  AOI21_X1 u1_u8_u3_U35 (.A( u1_u8_u3_n149 ) , .B2( u1_u8_u3_n150 ) , .B1( u1_u8_u3_n151 ) , .ZN( u1_u8_u3_n159 ) );
  AOI21_X1 u1_u8_u3_U36 (.A( u1_u8_u3_n154 ) , .B2( u1_u8_u3_n155 ) , .B1( u1_u8_u3_n156 ) , .ZN( u1_u8_u3_n157 ) );
  AOI211_X1 u1_u8_u3_U37 (.ZN( u1_u8_u3_n109 ) , .A( u1_u8_u3_n119 ) , .C2( u1_u8_u3_n129 ) , .B( u1_u8_u3_n138 ) , .C1( u1_u8_u3_n141 ) );
  AOI211_X1 u1_u8_u3_U38 (.B( u1_u8_u3_n119 ) , .A( u1_u8_u3_n120 ) , .C2( u1_u8_u3_n121 ) , .ZN( u1_u8_u3_n122 ) , .C1( u1_u8_u3_n179 ) );
  INV_X1 u1_u8_u3_U39 (.A( u1_u8_u3_n156 ) , .ZN( u1_u8_u3_n179 ) );
  INV_X1 u1_u8_u3_U4 (.A( u1_u8_u3_n140 ) , .ZN( u1_u8_u3_n182 ) );
  OAI22_X1 u1_u8_u3_U40 (.B1( u1_u8_u3_n118 ) , .ZN( u1_u8_u3_n120 ) , .A1( u1_u8_u3_n135 ) , .B2( u1_u8_u3_n154 ) , .A2( u1_u8_u3_n178 ) );
  AND3_X1 u1_u8_u3_U41 (.ZN( u1_u8_u3_n118 ) , .A2( u1_u8_u3_n124 ) , .A1( u1_u8_u3_n144 ) , .A3( u1_u8_u3_n152 ) );
  INV_X1 u1_u8_u3_U42 (.A( u1_u8_u3_n121 ) , .ZN( u1_u8_u3_n164 ) );
  NAND2_X1 u1_u8_u3_U43 (.ZN( u1_u8_u3_n133 ) , .A1( u1_u8_u3_n154 ) , .A2( u1_u8_u3_n164 ) );
  OAI211_X1 u1_u8_u3_U44 (.B( u1_u8_u3_n127 ) , .ZN( u1_u8_u3_n139 ) , .C1( u1_u8_u3_n150 ) , .C2( u1_u8_u3_n154 ) , .A( u1_u8_u3_n184 ) );
  INV_X1 u1_u8_u3_U45 (.A( u1_u8_u3_n125 ) , .ZN( u1_u8_u3_n184 ) );
  AOI221_X1 u1_u8_u3_U46 (.A( u1_u8_u3_n126 ) , .ZN( u1_u8_u3_n127 ) , .C2( u1_u8_u3_n132 ) , .C1( u1_u8_u3_n169 ) , .B2( u1_u8_u3_n170 ) , .B1( u1_u8_u3_n174 ) );
  OAI22_X1 u1_u8_u3_U47 (.A1( u1_u8_u3_n124 ) , .ZN( u1_u8_u3_n125 ) , .B2( u1_u8_u3_n145 ) , .A2( u1_u8_u3_n165 ) , .B1( u1_u8_u3_n167 ) );
  NOR2_X1 u1_u8_u3_U48 (.A1( u1_u8_u3_n113 ) , .ZN( u1_u8_u3_n131 ) , .A2( u1_u8_u3_n154 ) );
  NAND2_X1 u1_u8_u3_U49 (.A1( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n150 ) , .A2( u1_u8_u3_n99 ) );
  INV_X1 u1_u8_u3_U5 (.A( u1_u8_u3_n117 ) , .ZN( u1_u8_u3_n178 ) );
  NAND2_X1 u1_u8_u3_U50 (.A2( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n155 ) , .A1( u1_u8_u3_n97 ) );
  INV_X1 u1_u8_u3_U51 (.A( u1_u8_u3_n141 ) , .ZN( u1_u8_u3_n167 ) );
  AOI21_X1 u1_u8_u3_U52 (.B2( u1_u8_u3_n114 ) , .B1( u1_u8_u3_n146 ) , .A( u1_u8_u3_n154 ) , .ZN( u1_u8_u3_n94 ) );
  AOI21_X1 u1_u8_u3_U53 (.ZN( u1_u8_u3_n110 ) , .B2( u1_u8_u3_n142 ) , .B1( u1_u8_u3_n186 ) , .A( u1_u8_u3_n95 ) );
  INV_X1 u1_u8_u3_U54 (.A( u1_u8_u3_n145 ) , .ZN( u1_u8_u3_n186 ) );
  AOI21_X1 u1_u8_u3_U55 (.B1( u1_u8_u3_n124 ) , .A( u1_u8_u3_n149 ) , .B2( u1_u8_u3_n155 ) , .ZN( u1_u8_u3_n95 ) );
  INV_X1 u1_u8_u3_U56 (.A( u1_u8_u3_n149 ) , .ZN( u1_u8_u3_n169 ) );
  NAND2_X1 u1_u8_u3_U57 (.ZN( u1_u8_u3_n124 ) , .A1( u1_u8_u3_n96 ) , .A2( u1_u8_u3_n97 ) );
  NAND2_X1 u1_u8_u3_U58 (.A2( u1_u8_u3_n100 ) , .ZN( u1_u8_u3_n146 ) , .A1( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U59 (.A1( u1_u8_u3_n101 ) , .ZN( u1_u8_u3_n145 ) , .A2( u1_u8_u3_n99 ) );
  AOI221_X1 u1_u8_u3_U6 (.A( u1_u8_u3_n131 ) , .C2( u1_u8_u3_n132 ) , .C1( u1_u8_u3_n133 ) , .ZN( u1_u8_u3_n134 ) , .B1( u1_u8_u3_n143 ) , .B2( u1_u8_u3_n177 ) );
  NAND2_X1 u1_u8_u3_U60 (.A1( u1_u8_u3_n100 ) , .ZN( u1_u8_u3_n156 ) , .A2( u1_u8_u3_n99 ) );
  NAND2_X1 u1_u8_u3_U61 (.A2( u1_u8_u3_n101 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n148 ) );
  NAND2_X1 u1_u8_u3_U62 (.A1( u1_u8_u3_n100 ) , .A2( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n128 ) );
  NAND2_X1 u1_u8_u3_U63 (.A2( u1_u8_u3_n101 ) , .A1( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n152 ) );
  NAND2_X1 u1_u8_u3_U64 (.A2( u1_u8_u3_n101 ) , .ZN( u1_u8_u3_n114 ) , .A1( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U65 (.ZN( u1_u8_u3_n107 ) , .A1( u1_u8_u3_n97 ) , .A2( u1_u8_u3_n99 ) );
  NAND2_X1 u1_u8_u3_U66 (.A2( u1_u8_u3_n100 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n113 ) );
  NAND2_X1 u1_u8_u3_U67 (.A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n153 ) , .A2( u1_u8_u3_n97 ) );
  NAND2_X1 u1_u8_u3_U68 (.A2( u1_u8_u3_n103 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n130 ) );
  NAND2_X1 u1_u8_u3_U69 (.A2( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n144 ) , .A1( u1_u8_u3_n96 ) );
  OAI22_X1 u1_u8_u3_U7 (.B2( u1_u8_u3_n147 ) , .A2( u1_u8_u3_n148 ) , .ZN( u1_u8_u3_n160 ) , .B1( u1_u8_u3_n165 ) , .A1( u1_u8_u3_n168 ) );
  NAND2_X1 u1_u8_u3_U70 (.A1( u1_u8_u3_n102 ) , .A2( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n108 ) );
  NOR2_X1 u1_u8_u3_U71 (.A2( u1_u8_X_19 ) , .A1( u1_u8_X_20 ) , .ZN( u1_u8_u3_n99 ) );
  NOR2_X1 u1_u8_u3_U72 (.A2( u1_u8_X_21 ) , .A1( u1_u8_X_24 ) , .ZN( u1_u8_u3_n103 ) );
  NOR2_X1 u1_u8_u3_U73 (.A2( u1_u8_X_24 ) , .A1( u1_u8_u3_n171 ) , .ZN( u1_u8_u3_n97 ) );
  NOR2_X1 u1_u8_u3_U74 (.A2( u1_u8_X_23 ) , .ZN( u1_u8_u3_n141 ) , .A1( u1_u8_u3_n166 ) );
  NOR2_X1 u1_u8_u3_U75 (.A2( u1_u8_X_19 ) , .A1( u1_u8_u3_n172 ) , .ZN( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U76 (.A1( u1_u8_X_22 ) , .A2( u1_u8_X_23 ) , .ZN( u1_u8_u3_n154 ) );
  NAND2_X1 u1_u8_u3_U77 (.A1( u1_u8_X_23 ) , .ZN( u1_u8_u3_n149 ) , .A2( u1_u8_u3_n166 ) );
  NOR2_X1 u1_u8_u3_U78 (.A2( u1_u8_X_22 ) , .A1( u1_u8_X_23 ) , .ZN( u1_u8_u3_n121 ) );
  AND2_X1 u1_u8_u3_U79 (.A1( u1_u8_X_24 ) , .ZN( u1_u8_u3_n101 ) , .A2( u1_u8_u3_n171 ) );
  AND3_X1 u1_u8_u3_U8 (.A3( u1_u8_u3_n144 ) , .A2( u1_u8_u3_n145 ) , .A1( u1_u8_u3_n146 ) , .ZN( u1_u8_u3_n147 ) );
  AND2_X1 u1_u8_u3_U80 (.A1( u1_u8_X_19 ) , .ZN( u1_u8_u3_n102 ) , .A2( u1_u8_u3_n172 ) );
  AND2_X1 u1_u8_u3_U81 (.A1( u1_u8_X_21 ) , .A2( u1_u8_X_24 ) , .ZN( u1_u8_u3_n100 ) );
  AND2_X1 u1_u8_u3_U82 (.A2( u1_u8_X_19 ) , .A1( u1_u8_X_20 ) , .ZN( u1_u8_u3_n104 ) );
  INV_X1 u1_u8_u3_U83 (.A( u1_u8_X_22 ) , .ZN( u1_u8_u3_n166 ) );
  INV_X1 u1_u8_u3_U84 (.A( u1_u8_X_21 ) , .ZN( u1_u8_u3_n171 ) );
  INV_X1 u1_u8_u3_U85 (.A( u1_u8_X_20 ) , .ZN( u1_u8_u3_n172 ) );
  OR4_X1 u1_u8_u3_U86 (.ZN( u1_out8_10 ) , .A4( u1_u8_u3_n136 ) , .A3( u1_u8_u3_n137 ) , .A1( u1_u8_u3_n138 ) , .A2( u1_u8_u3_n139 ) );
  OAI222_X1 u1_u8_u3_U87 (.C1( u1_u8_u3_n128 ) , .ZN( u1_u8_u3_n137 ) , .B1( u1_u8_u3_n148 ) , .A2( u1_u8_u3_n150 ) , .B2( u1_u8_u3_n154 ) , .C2( u1_u8_u3_n164 ) , .A1( u1_u8_u3_n167 ) );
  OAI221_X1 u1_u8_u3_U88 (.A( u1_u8_u3_n134 ) , .B2( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n136 ) , .C1( u1_u8_u3_n149 ) , .B1( u1_u8_u3_n151 ) , .C2( u1_u8_u3_n183 ) );
  NAND4_X1 u1_u8_u3_U89 (.ZN( u1_out8_26 ) , .A4( u1_u8_u3_n109 ) , .A3( u1_u8_u3_n110 ) , .A2( u1_u8_u3_n111 ) , .A1( u1_u8_u3_n173 ) );
  INV_X1 u1_u8_u3_U9 (.A( u1_u8_u3_n143 ) , .ZN( u1_u8_u3_n168 ) );
  INV_X1 u1_u8_u3_U90 (.ZN( u1_u8_u3_n173 ) , .A( u1_u8_u3_n94 ) );
  OAI21_X1 u1_u8_u3_U91 (.ZN( u1_u8_u3_n111 ) , .B2( u1_u8_u3_n117 ) , .A( u1_u8_u3_n133 ) , .B1( u1_u8_u3_n176 ) );
  NAND4_X1 u1_u8_u3_U92 (.ZN( u1_out8_20 ) , .A4( u1_u8_u3_n122 ) , .A3( u1_u8_u3_n123 ) , .A1( u1_u8_u3_n175 ) , .A2( u1_u8_u3_n180 ) );
  INV_X1 u1_u8_u3_U93 (.A( u1_u8_u3_n126 ) , .ZN( u1_u8_u3_n180 ) );
  INV_X1 u1_u8_u3_U94 (.A( u1_u8_u3_n112 ) , .ZN( u1_u8_u3_n175 ) );
  NAND4_X1 u1_u8_u3_U95 (.ZN( u1_out8_1 ) , .A4( u1_u8_u3_n161 ) , .A3( u1_u8_u3_n162 ) , .A2( u1_u8_u3_n163 ) , .A1( u1_u8_u3_n185 ) );
  NAND2_X1 u1_u8_u3_U96 (.ZN( u1_u8_u3_n163 ) , .A2( u1_u8_u3_n170 ) , .A1( u1_u8_u3_n176 ) );
  AOI22_X1 u1_u8_u3_U97 (.B2( u1_u8_u3_n140 ) , .B1( u1_u8_u3_n141 ) , .A2( u1_u8_u3_n142 ) , .ZN( u1_u8_u3_n162 ) , .A1( u1_u8_u3_n177 ) );
  NAND3_X1 u1_u8_u3_U98 (.A1( u1_u8_u3_n114 ) , .ZN( u1_u8_u3_n115 ) , .A2( u1_u8_u3_n145 ) , .A3( u1_u8_u3_n153 ) );
  NAND3_X1 u1_u8_u3_U99 (.ZN( u1_u8_u3_n129 ) , .A2( u1_u8_u3_n144 ) , .A1( u1_u8_u3_n153 ) , .A3( u1_u8_u3_n182 ) );
  XOR2_X1 u1_u9_U10 (.B( u1_K10_45 ) , .A( u1_R8_30 ) , .Z( u1_u9_X_45 ) );
  XOR2_X1 u1_u9_U11 (.B( u1_K10_44 ) , .A( u1_R8_29 ) , .Z( u1_u9_X_44 ) );
  XOR2_X1 u1_u9_U12 (.B( u1_K10_43 ) , .A( u1_R8_28 ) , .Z( u1_u9_X_43 ) );
  XOR2_X1 u1_u9_U7 (.B( u1_K10_48 ) , .A( u1_R8_1 ) , .Z( u1_u9_X_48 ) );
  XOR2_X1 u1_u9_U8 (.B( u1_K10_47 ) , .A( u1_R8_32 ) , .Z( u1_u9_X_47 ) );
  XOR2_X1 u1_u9_U9 (.B( u1_K10_46 ) , .A( u1_R8_31 ) , .Z( u1_u9_X_46 ) );
  AND3_X1 u1_u9_u7_U10 (.A3( u1_u9_u7_n110 ) , .A2( u1_u9_u7_n127 ) , .A1( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U11 (.A( u1_u9_u7_n161 ) , .B1( u1_u9_u7_n168 ) , .B2( u1_u9_u7_n173 ) , .ZN( u1_u9_u7_n91 ) );
  AOI211_X1 u1_u9_u7_U12 (.A( u1_u9_u7_n117 ) , .ZN( u1_u9_u7_n118 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n177 ) , .B( u1_u9_u7_n180 ) );
  OAI22_X1 u1_u9_u7_U13 (.B1( u1_u9_u7_n115 ) , .ZN( u1_u9_u7_n117 ) , .A2( u1_u9_u7_n133 ) , .A1( u1_u9_u7_n137 ) , .B2( u1_u9_u7_n162 ) );
  INV_X1 u1_u9_u7_U14 (.A( u1_u9_u7_n116 ) , .ZN( u1_u9_u7_n180 ) );
  NOR3_X1 u1_u9_u7_U15 (.ZN( u1_u9_u7_n115 ) , .A3( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n168 ) , .A1( u1_u9_u7_n169 ) );
  OAI211_X1 u1_u9_u7_U16 (.B( u1_u9_u7_n122 ) , .A( u1_u9_u7_n123 ) , .C2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n154 ) , .C1( u1_u9_u7_n162 ) );
  AOI222_X1 u1_u9_u7_U17 (.ZN( u1_u9_u7_n122 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n161 ) , .A2( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n170 ) , .A1( u1_u9_u7_n176 ) );
  INV_X1 u1_u9_u7_U18 (.A( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n176 ) );
  NOR3_X1 u1_u9_u7_U19 (.A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n135 ) , .ZN( u1_u9_u7_n136 ) , .A3( u1_u9_u7_n171 ) );
  NOR2_X1 u1_u9_u7_U20 (.A1( u1_u9_u7_n130 ) , .A2( u1_u9_u7_n134 ) , .ZN( u1_u9_u7_n153 ) );
  INV_X1 u1_u9_u7_U21 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n165 ) );
  NOR2_X1 u1_u9_u7_U22 (.ZN( u1_u9_u7_n111 ) , .A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n169 ) );
  AOI21_X1 u1_u9_u7_U23 (.ZN( u1_u9_u7_n104 ) , .B2( u1_u9_u7_n112 ) , .B1( u1_u9_u7_n127 ) , .A( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U24 (.ZN( u1_u9_u7_n106 ) , .B1( u1_u9_u7_n133 ) , .B2( u1_u9_u7_n146 ) , .A( u1_u9_u7_n162 ) );
  AOI21_X1 u1_u9_u7_U25 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n107 ) , .B2( u1_u9_u7_n128 ) , .B1( u1_u9_u7_n175 ) );
  INV_X1 u1_u9_u7_U26 (.A( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n171 ) );
  INV_X1 u1_u9_u7_U27 (.A( u1_u9_u7_n131 ) , .ZN( u1_u9_u7_n177 ) );
  INV_X1 u1_u9_u7_U28 (.A( u1_u9_u7_n110 ) , .ZN( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U29 (.A1( u1_u9_u7_n129 ) , .A2( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n149 ) );
  OAI21_X1 u1_u9_u7_U3 (.ZN( u1_u9_u7_n159 ) , .A( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n171 ) , .B1( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U30 (.A1( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n130 ) );
  INV_X1 u1_u9_u7_U31 (.A( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n173 ) );
  INV_X1 u1_u9_u7_U32 (.A( u1_u9_u7_n128 ) , .ZN( u1_u9_u7_n168 ) );
  INV_X1 u1_u9_u7_U33 (.A( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n169 ) );
  INV_X1 u1_u9_u7_U34 (.A( u1_u9_u7_n127 ) , .ZN( u1_u9_u7_n179 ) );
  NOR2_X1 u1_u9_u7_U35 (.ZN( u1_u9_u7_n101 ) , .A2( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n156 ) );
  AOI211_X1 u1_u9_u7_U36 (.B( u1_u9_u7_n154 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n156 ) , .ZN( u1_u9_u7_n157 ) , .C2( u1_u9_u7_n172 ) );
  INV_X1 u1_u9_u7_U37 (.A( u1_u9_u7_n153 ) , .ZN( u1_u9_u7_n172 ) );
  AOI211_X1 u1_u9_u7_U38 (.B( u1_u9_u7_n139 ) , .A( u1_u9_u7_n140 ) , .C2( u1_u9_u7_n141 ) , .ZN( u1_u9_u7_n142 ) , .C1( u1_u9_u7_n156 ) );
  NAND4_X1 u1_u9_u7_U39 (.A3( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n141 ) , .A4( u1_u9_u7_n147 ) );
  INV_X1 u1_u9_u7_U4 (.A( u1_u9_u7_n111 ) , .ZN( u1_u9_u7_n170 ) );
  AOI21_X1 u1_u9_u7_U40 (.A( u1_u9_u7_n137 ) , .B1( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n139 ) , .B2( u1_u9_u7_n146 ) );
  OAI22_X1 u1_u9_u7_U41 (.B1( u1_u9_u7_n136 ) , .ZN( u1_u9_u7_n140 ) , .A1( u1_u9_u7_n153 ) , .B2( u1_u9_u7_n162 ) , .A2( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U42 (.ZN( u1_u9_u7_n123 ) , .B1( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n177 ) , .A( u1_u9_u7_n97 ) );
  AOI21_X1 u1_u9_u7_U43 (.B2( u1_u9_u7_n113 ) , .B1( u1_u9_u7_n124 ) , .A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n97 ) );
  INV_X1 u1_u9_u7_U44 (.A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U45 (.A( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n162 ) );
  AOI22_X1 u1_u9_u7_U46 (.A2( u1_u9_u7_n114 ) , .ZN( u1_u9_u7_n119 ) , .B1( u1_u9_u7_n130 ) , .A1( u1_u9_u7_n156 ) , .B2( u1_u9_u7_n165 ) );
  NAND2_X1 u1_u9_u7_U47 (.A2( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n114 ) , .A1( u1_u9_u7_n175 ) );
  AND2_X1 u1_u9_u7_U48 (.ZN( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n98 ) , .A1( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U49 (.ZN( u1_u9_u7_n137 ) , .A1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U5 (.A( u1_u9_u7_n149 ) , .ZN( u1_u9_u7_n175 ) );
  AOI21_X1 u1_u9_u7_U50 (.ZN( u1_u9_u7_n105 ) , .B2( u1_u9_u7_n110 ) , .A( u1_u9_u7_n125 ) , .B1( u1_u9_u7_n147 ) );
  NAND2_X1 u1_u9_u7_U51 (.ZN( u1_u9_u7_n146 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U52 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U53 (.A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n99 ) );
  OR2_X1 u1_u9_u7_U54 (.ZN( u1_u9_u7_n126 ) , .A2( u1_u9_u7_n152 ) , .A1( u1_u9_u7_n156 ) );
  NAND2_X1 u1_u9_u7_U55 (.A2( u1_u9_u7_n102 ) , .A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n133 ) );
  NAND2_X1 u1_u9_u7_U56 (.ZN( u1_u9_u7_n112 ) , .A2( u1_u9_u7_n96 ) , .A1( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U57 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U58 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U59 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n124 ) , .A1( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U6 (.A( u1_u9_u7_n154 ) , .ZN( u1_u9_u7_n178 ) );
  NAND2_X1 u1_u9_u7_U60 (.ZN( u1_u9_u7_n110 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U61 (.A( u1_u9_u7_n150 ) , .ZN( u1_u9_u7_n164 ) );
  AND2_X1 u1_u9_u7_U62 (.ZN( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U63 (.A1( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n129 ) );
  NAND2_X1 u1_u9_u7_U64 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n131 ) , .A1( u1_u9_u7_n95 ) );
  NAND2_X1 u1_u9_u7_U65 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n138 ) , .A2( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U66 (.ZN( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n96 ) );
  NAND2_X1 u1_u9_u7_U67 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n148 ) , .A2( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U68 (.A2( u1_u9_X_47 ) , .ZN( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n163 ) );
  NOR2_X1 u1_u9_u7_U69 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n103 ) );
  AOI211_X1 u1_u9_u7_U7 (.ZN( u1_u9_u7_n116 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n161 ) , .C2( u1_u9_u7_n171 ) , .B( u1_u9_u7_n94 ) );
  NOR2_X1 u1_u9_u7_U70 (.A2( u1_u9_X_48 ) , .A1( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U71 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U72 (.A2( u1_u9_X_44 ) , .A1( u1_u9_u7_n167 ) , .ZN( u1_u9_u7_n98 ) );
  NOR2_X1 u1_u9_u7_U73 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n152 ) );
  AND2_X1 u1_u9_u7_U74 (.A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n156 ) , .A2( u1_u9_u7_n163 ) );
  NAND2_X1 u1_u9_u7_U75 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n125 ) );
  AND2_X1 u1_u9_u7_U76 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n102 ) );
  AND2_X1 u1_u9_u7_U77 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n96 ) );
  AND2_X1 u1_u9_u7_U78 (.A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n167 ) );
  AND2_X1 u1_u9_u7_U79 (.A1( u1_u9_X_48 ) , .A2( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n93 ) );
  OAI222_X1 u1_u9_u7_U8 (.C2( u1_u9_u7_n101 ) , .B2( u1_u9_u7_n111 ) , .A1( u1_u9_u7_n113 ) , .C1( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n162 ) , .B1( u1_u9_u7_n164 ) , .ZN( u1_u9_u7_n94 ) );
  INV_X1 u1_u9_u7_U80 (.A( u1_u9_X_46 ) , .ZN( u1_u9_u7_n163 ) );
  INV_X1 u1_u9_u7_U81 (.A( u1_u9_X_43 ) , .ZN( u1_u9_u7_n167 ) );
  INV_X1 u1_u9_u7_U82 (.A( u1_u9_X_45 ) , .ZN( u1_u9_u7_n166 ) );
  NAND4_X1 u1_u9_u7_U83 (.ZN( u1_out9_5 ) , .A4( u1_u9_u7_n108 ) , .A3( u1_u9_u7_n109 ) , .A1( u1_u9_u7_n116 ) , .A2( u1_u9_u7_n123 ) );
  AOI22_X1 u1_u9_u7_U84 (.ZN( u1_u9_u7_n109 ) , .A2( u1_u9_u7_n126 ) , .B2( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n156 ) , .A1( u1_u9_u7_n171 ) );
  NOR4_X1 u1_u9_u7_U85 (.A4( u1_u9_u7_n104 ) , .A3( u1_u9_u7_n105 ) , .A2( u1_u9_u7_n106 ) , .A1( u1_u9_u7_n107 ) , .ZN( u1_u9_u7_n108 ) );
  NAND4_X1 u1_u9_u7_U86 (.ZN( u1_out9_27 ) , .A4( u1_u9_u7_n118 ) , .A3( u1_u9_u7_n119 ) , .A2( u1_u9_u7_n120 ) , .A1( u1_u9_u7_n121 ) );
  OAI21_X1 u1_u9_u7_U87 (.ZN( u1_u9_u7_n121 ) , .B2( u1_u9_u7_n145 ) , .A( u1_u9_u7_n150 ) , .B1( u1_u9_u7_n174 ) );
  OAI21_X1 u1_u9_u7_U88 (.ZN( u1_u9_u7_n120 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n170 ) , .B1( u1_u9_u7_n179 ) );
  NAND4_X1 u1_u9_u7_U89 (.ZN( u1_out9_21 ) , .A4( u1_u9_u7_n157 ) , .A3( u1_u9_u7_n158 ) , .A2( u1_u9_u7_n159 ) , .A1( u1_u9_u7_n160 ) );
  OAI221_X1 u1_u9_u7_U9 (.C1( u1_u9_u7_n101 ) , .C2( u1_u9_u7_n147 ) , .ZN( u1_u9_u7_n155 ) , .B2( u1_u9_u7_n162 ) , .A( u1_u9_u7_n91 ) , .B1( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U90 (.B1( u1_u9_u7_n145 ) , .ZN( u1_u9_u7_n160 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n177 ) );
  AOI22_X1 u1_u9_u7_U91 (.B2( u1_u9_u7_n149 ) , .B1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n151 ) , .A1( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n158 ) );
  NAND4_X1 u1_u9_u7_U92 (.ZN( u1_out9_15 ) , .A4( u1_u9_u7_n142 ) , .A3( u1_u9_u7_n143 ) , .A2( u1_u9_u7_n144 ) , .A1( u1_u9_u7_n178 ) );
  OR2_X1 u1_u9_u7_U93 (.A2( u1_u9_u7_n125 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n144 ) );
  AOI22_X1 u1_u9_u7_U94 (.A2( u1_u9_u7_n126 ) , .ZN( u1_u9_u7_n143 ) , .B2( u1_u9_u7_n165 ) , .B1( u1_u9_u7_n173 ) , .A1( u1_u9_u7_n174 ) );
  NAND3_X1 u1_u9_u7_U95 (.A3( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n151 ) );
  NAND3_X1 u1_u9_u7_U96 (.A3( u1_u9_u7_n131 ) , .A2( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n135 ) );
  OAI21_X1 u1_uk_U1000 (.ZN( u1_K6_23 ) , .A( u1_uk_n1093 ) , .B2( u1_uk_n1472 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1001 (.A1( u1_uk_K_r4_27 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1093 ) );
  OAI22_X1 u1_uk_U101 (.ZN( u1_K15_41 ) , .B2( u1_uk_n1865 ) , .A2( u1_uk_n1883 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1026 (.ZN( u1_K1_37 ) , .A( u1_uk_n1013 ) , .B2( u1_uk_n1174 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U1027 (.A1( u1_key_r_50 ) , .ZN( u1_uk_n1013 ) , .A2( u1_uk_n162 ) );
  OAI21_X1 u1_uk_U1046 (.ZN( u1_K6_41 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1099 ) , .B2( u1_uk_n1475 ) );
  NAND2_X1 u1_uk_U1047 (.A1( u1_uk_K_r4_31 ) , .ZN( u1_uk_n1099 ) , .A2( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1054 (.ZN( u1_K9_14 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1151 ) , .B2( u1_uk_n1604 ) );
  NAND2_X1 u1_uk_U1055 (.A1( u1_uk_K_r7_34 ) , .A2( u1_uk_n100 ) , .ZN( u1_uk_n1151 ) );
  OAI21_X1 u1_uk_U1066 (.ZN( u1_K15_32 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1855 ) , .A( u1_uk_n971 ) );
  NAND2_X1 u1_uk_U1067 (.A1( u1_uk_K_r13_36 ) , .A2( u1_uk_n147 ) , .ZN( u1_uk_n971 ) );
  INV_X1 u1_uk_U1078 (.A( u1_key_r_9 ) , .ZN( u1_uk_n1179 ) );
  INV_X1 u1_uk_U1079 (.A( u1_key_r_7 ) , .ZN( u1_uk_n1177 ) );
  INV_X1 u1_uk_U1083 (.A( u1_key_r_23 ) , .ZN( u1_uk_n1188 ) );
  INV_X1 u1_uk_U1086 (.A( u1_key_r_30 ) , .ZN( u1_uk_n1195 ) );
  INV_X1 u1_uk_U1092 (.A( u1_key_r_37 ) , .ZN( u1_uk_n1201 ) );
  INV_X1 u1_uk_U1093 (.A( u1_key_r_52 ) , .ZN( u1_uk_n1213 ) );
  INV_X1 u1_uk_U1094 (.A( u1_key_r_0 ) , .ZN( u1_uk_n1172 ) );
  INV_X1 u1_uk_U1095 (.A( u1_key_r_16 ) , .ZN( u1_uk_n1182 ) );
  INV_X1 u1_uk_U1097 (.A( u1_key_r_1 ) , .ZN( u1_uk_n1173 ) );
  INV_X1 u1_uk_U1098 (.A( u1_key_r_2 ) , .ZN( u1_uk_n1174 ) );
  INV_X1 u1_uk_U1119 (.ZN( u1_K9_11 ) , .A( u1_uk_n1148 ) );
  AOI22_X1 u1_uk_U1120 (.B2( u1_uk_K_r7_48 ) , .A2( u1_uk_K_r7_55 ) , .B1( u1_uk_n109 ) , .ZN( u1_uk_n1148 ) , .A1( u1_uk_n220 ) );
  INV_X1 u1_uk_U1127 (.ZN( u1_K1_41 ) , .A( u1_uk_n1015 ) );
  AOI22_X1 u1_uk_U1128 (.B2( u1_key_r_35 ) , .A2( u1_key_r_42 ) , .ZN( u1_uk_n1015 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n298 ) );
  INV_X1 u1_uk_U1145 (.ZN( u1_K9_20 ) , .A( u1_uk_n1156 ) );
  AOI22_X1 u1_uk_U1146 (.B2( u1_uk_K_r7_32 ) , .A2( u1_uk_K_r7_39 ) , .B1( u1_uk_n11 ) , .ZN( u1_uk_n1156 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U115 (.ZN( u1_K9_5 ) , .B2( u1_uk_n1610 ) , .A2( u1_uk_n1616 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n188 ) );
  INV_X1 u1_uk_U1151 (.ZN( u1_K1_32 ) , .A( u1_uk_n1010 ) );
  AOI22_X1 u1_uk_U1152 (.B2( u1_key_r_22 ) , .A2( u1_key_r_29 ) , .ZN( u1_uk_n1010 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) );
  INV_X1 u1_uk_U1155 (.ZN( u1_K6_2 ) , .A( u1_uk_n1096 ) );
  AOI22_X1 u1_uk_U1156 (.B2( u1_uk_K_r4_17 ) , .A2( u1_uk_K_r4_55 ) , .ZN( u1_uk_n1096 ) , .B1( u1_uk_n257 ) , .A1( u1_uk_n27 ) );
  AOI22_X1 u1_uk_U1165 (.B1( n116 ) , .A2( u1_uk_K_r13_2 ) , .B2( u1_uk_K_r13_23 ) , .A1( u1_uk_n286 ) , .ZN( u1_uk_n974 ) );
  INV_X1 u1_uk_U1166 (.ZN( u1_K15_43 ) , .A( u1_uk_n974 ) );
  INV_X1 u1_uk_U1170 (.ZN( u1_K9_2 ) , .A( u1_uk_n1160 ) );
  OAI22_X1 u1_uk_U128 (.ZN( u1_K10_47 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1624 ) , .B2( u1_uk_n1639 ) , .B1( u1_uk_n223 ) );
  INV_X1 u1_uk_U15 (.A( u1_uk_n188 ) , .ZN( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U150 (.ZN( u1_K6_19 ) , .A( u1_uk_n1091 ) , .B2( u1_uk_n1444 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U151 (.A1( u1_uk_K_r4_48 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1091 ) );
  INV_X1 u1_uk_U163 (.ZN( u1_K9_19 ) , .A( u1_uk_n1154 ) );
  AOI22_X1 u1_uk_U164 (.B1( u1_uk_K_r7_13 ) , .A2( u1_uk_K_r7_20 ) , .ZN( u1_uk_n1154 ) , .A1( u1_uk_n291 ) , .B2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U194 (.ZN( u1_K6_14 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1440 ) , .B2( u1_uk_n1446 ) , .B1( u1_uk_n257 ) );
  OAI21_X1 u1_uk_U209 (.ZN( u1_K1_30 ) , .A( u1_uk_n1009 ) , .B2( u1_uk_n1213 ) , .B1( u1_uk_n93 ) );
  NAND2_X1 u1_uk_U210 (.A1( u1_key_r_45 ) , .ZN( u1_uk_n1009 ) , .A2( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U220 (.ZN( u1_K1_31 ) , .A2( u1_uk_n1177 ) , .B2( u1_uk_n1181 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U221 (.A( u1_key_r_14 ) , .ZN( u1_uk_n1181 ) );
  OAI22_X1 u1_uk_U236 (.ZN( u1_K6_31 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1455 ) , .A2( u1_uk_n1460 ) , .A1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U238 (.ZN( u1_K5_31 ) , .B1( u1_uk_n100 ) , .A( u1_uk_n1077 ) , .B2( u1_uk_n1401 ) );
  NAND2_X1 u1_uk_U239 (.A1( u1_uk_K_r3_44 ) , .ZN( u1_uk_n1077 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U240 (.ZN( u1_K15_31 ) , .B2( u1_uk_n1843 ) , .A2( u1_uk_n1860 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U241 (.ZN( u1_K1_39 ) , .A( u1_uk_n1014 ) , .B2( u1_uk_n1187 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U242 (.A1( u1_key_r_15 ) , .ZN( u1_uk_n1014 ) , .A2( u1_uk_n155 ) );
  INV_X1 u1_uk_U243 (.A( u1_key_r_22 ) , .ZN( u1_uk_n1187 ) );
  OAI22_X1 u1_uk_U246 (.ZN( u1_K15_39 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1848 ) , .B2( u1_uk_n1866 ) , .B1( u1_uk_n214 ) );
  INV_X1 u1_uk_U259 (.ZN( u1_K1_48 ) , .A( u1_uk_n1019 ) );
  AOI22_X1 u1_uk_U260 (.B2( u1_key_r_21 ) , .A2( u1_key_r_28 ) , .ZN( u1_uk_n1019 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n291 ) );
  INV_X1 u1_uk_U261 (.ZN( u1_K1_44 ) , .A( u1_uk_n1017 ) );
  AOI22_X1 u1_uk_U262 (.B2( u1_key_r_36 ) , .A2( u1_key_r_43 ) , .ZN( u1_uk_n1017 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U263 (.ZN( u1_K15_44 ) , .B2( u1_uk_n1866 ) , .A2( u1_uk_n1884 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U264 (.ZN( u1_K15_48 ) , .B1( u1_uk_n10 ) , .B2( u1_uk_n1854 ) , .A( u1_uk_n975 ) );
  NAND2_X1 u1_uk_U265 (.A1( u1_uk_K_r13_35 ) , .A2( u1_uk_n148 ) , .ZN( u1_uk_n975 ) );
  OAI22_X1 u1_uk_U274 (.ZN( u1_K10_44 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1627 ) , .A2( u1_uk_n1647 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U275 (.ZN( u1_K10_48 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1640 ) , .A2( u1_uk_n1656 ) , .A1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U290 (.ZN( u1_K6_6 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1474 ) , .A2( u1_uk_n1478 ) , .A1( u1_uk_n231 ) );
  INV_X1 u1_uk_U306 (.ZN( u1_K4_8 ) , .A( u1_uk_n1070 ) );
  AOI22_X1 u1_uk_U307 (.B2( u1_uk_K_r2_41 ) , .A2( u1_uk_K_r2_46 ) , .ZN( u1_uk_n1070 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U312 (.ZN( u1_K1_26 ) , .A( u1_uk_n1006 ) );
  AOI22_X1 u1_uk_U313 (.B2( u1_key_r_31 ) , .A2( u1_key_r_51 ) , .ZN( u1_uk_n1006 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n240 ) );
  OAI21_X1 u1_uk_U321 (.ZN( u1_K6_26 ) , .A( u1_uk_n1094 ) , .B2( u1_uk_n1469 ) , .B1( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U322 (.A1( u1_uk_K_r4_35 ) , .ZN( u1_uk_n1094 ) , .A2( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U336 (.ZN( u1_K15_46 ) , .A2( u1_uk_n1848 ) , .B2( u1_uk_n1875 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U343 (.ZN( u1_K1_46 ) , .A( u1_uk_n1018 ) , .B2( u1_uk_n1173 ) , .B1( u1_uk_n17 ) );
  NAND2_X1 u1_uk_U344 (.A1( u1_key_r_49 ) , .ZN( u1_uk_n1018 ) , .A2( u1_uk_n142 ) );
  INV_X1 u1_uk_U351 (.ZN( u1_K6_4 ) , .A( u1_uk_n1101 ) );
  AOI22_X1 u1_uk_U352 (.B2( u1_uk_K_r4_41 ) , .A2( u1_uk_K_r4_47 ) , .ZN( u1_uk_n1101 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U357 (.ZN( u1_K1_40 ) , .B2( u1_uk_n1172 ) , .A2( u1_uk_n1213 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U362 (.ZN( u1_K15_40 ) , .A2( u1_uk_n1847 ) , .B2( u1_uk_n1879 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U364 (.ZN( u1_K6_40 ) , .A2( u1_uk_n1442 ) , .B2( u1_uk_n1450 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n240 ) );
  BUF_X1 u1_uk_U37 (.Z( u1_uk_n213 ) , .A( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U378 (.ZN( u1_K15_33 ) , .B2( u1_uk_n1870 ) , .B1( u1_uk_n83 ) , .A( u1_uk_n972 ) );
  NAND2_X1 u1_uk_U379 (.A1( u1_uk_K_r13_31 ) , .A2( u1_uk_n60 ) , .ZN( u1_uk_n972 ) );
  OAI22_X1 u1_uk_U382 (.ZN( u1_K1_28 ) , .B2( u1_uk_n1173 ) , .A2( u1_uk_n1178 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U383 (.A( u1_key_r_8 ) , .ZN( u1_uk_n1178 ) );
  OAI22_X1 u1_uk_U386 (.ZN( u1_K6_28 ) , .B2( u1_uk_n1450 ) , .A2( u1_uk_n1477 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n250 ) );
  OAI21_X1 u1_uk_U388 (.ZN( u1_K5_33 ) , .A( u1_uk_n1078 ) , .B2( u1_uk_n1431 ) , .B1( u1_uk_n214 ) );
  NAND2_X1 u1_uk_U389 (.A1( u1_uk_K_r3_14 ) , .ZN( u1_uk_n1078 ) , .A2( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U407 (.ZN( u1_K9_16 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1578 ) , .A2( u1_uk_n1585 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U411 (.ZN( u1_K6_16 ) , .B2( u1_uk_n1466 ) , .A2( u1_uk_n1472 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U425 (.ZN( u1_K4_9 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1359 ) , .A2( u1_uk_n1369 ) , .B1( u1_uk_n231 ) );
  INV_X1 u1_uk_U447 (.ZN( u1_K9_9 ) , .A( u1_uk_n1171 ) );
  AOI22_X1 u1_uk_U448 (.B2( u1_uk_K_r7_13 ) , .A1( u1_uk_K_r7_6 ) , .ZN( u1_uk_n1171 ) , .A2( u1_uk_n148 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U465 (.ZN( u1_K1_33 ) , .A( u1_uk_n1011 ) );
  AOI22_X1 u1_uk_U466 (.B2( u1_key_r_44 ) , .A2( u1_key_r_51 ) , .ZN( u1_uk_n1011 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U468 (.ZN( u1_K6_33 ) , .B2( u1_uk_n1458 ) , .A2( u1_uk_n1463 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U470 (.ZN( u1_K15_37 ) , .A2( u1_uk_n1849 ) , .B2( u1_uk_n1876 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U477 (.ZN( u1_K6_37 ) , .A( u1_uk_n1098 ) , .B2( u1_uk_n1468 ) , .B1( u1_uk_n271 ) );
  NAND2_X1 u1_uk_U478 (.A1( u1_uk_K_r4_38 ) , .ZN( u1_uk_n1098 ) , .A2( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U480 (.ZN( u1_K1_29 ) , .B2( u1_uk_n1182 ) , .A2( u1_uk_n1188 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U499 (.ZN( u1_K6_29 ) , .A( u1_uk_n1095 ) , .B2( u1_uk_n1442 ) , .B1( u1_uk_n213 ) );
  NAND2_X1 u1_uk_U500 (.A1( u1_uk_K_r4_0 ) , .ZN( u1_uk_n1095 ) , .A2( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U514 (.ZN( u1_K9_12 ) , .A( u1_uk_n1149 ) , .B2( u1_uk_n1573 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U515 (.A1( u1_uk_K_r7_53 ) , .ZN( u1_uk_n1149 ) , .A2( u1_uk_n142 ) );
  OAI21_X1 u1_uk_U521 (.ZN( u1_K9_17 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1152 ) , .B2( u1_uk_n1598 ) );
  NAND2_X1 u1_uk_U522 (.A1( u1_uk_K_r7_26 ) , .ZN( u1_uk_n1152 ) , .A2( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U542 (.ZN( u1_K4_12 ) , .B2( u1_uk_n1371 ) , .A2( u1_uk_n1391 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U545 (.ZN( u1_K1_36 ) , .B2( u1_uk_n1188 ) , .A2( u1_uk_n1195 ) , .A1( u1_uk_n148 ) , .B1( u1_uk_n223 ) );
  INV_X1 u1_uk_U554 (.ZN( u1_K6_17 ) , .A( u1_uk_n1089 ) );
  AOI22_X1 u1_uk_U555 (.B2( u1_uk_K_r4_4 ) , .A2( u1_uk_K_r4_55 ) , .ZN( u1_uk_n1089 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U556 (.ZN( u1_K15_36 ) , .B2( u1_uk_n1856 ) , .A2( u1_uk_n1870 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U561 (.ZN( u1_K1_38 ) , .B2( u1_uk_n1195 ) , .A2( u1_uk_n1201 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n202 ) );
  INV_X1 u1_uk_U570 (.ZN( u1_K5_36 ) , .A( u1_uk_n1080 ) );
  AOI22_X1 u1_uk_U571 (.B2( u1_uk_K_r3_29 ) , .A2( u1_uk_K_r3_52 ) , .ZN( u1_uk_n1080 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U572 (.ZN( u1_K15_38 ) , .A( u1_uk_n973 ) );
  AOI22_X1 u1_uk_U573 (.B2( u1_uk_K_r13_23 ) , .A2( u1_uk_K_r13_44 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n220 ) , .ZN( u1_uk_n973 ) );
  OAI22_X1 u1_uk_U577 (.ZN( u1_K6_38 ) , .B2( u1_uk_n1448 ) , .B1( u1_uk_n145 ) , .A2( u1_uk_n1455 ) , .A1( u1_uk_n213 ) );
  INV_X1 u1_uk_U587 (.ZN( u1_K9_10 ) , .A( u1_uk_n1147 ) );
  AOI22_X1 u1_uk_U588 (.B1( n116 ) , .B2( u1_uk_K_r7_25 ) , .A2( u1_uk_K_r7_32 ) , .ZN( u1_uk_n1147 ) , .A1( u1_uk_n208 ) );
  INV_X1 u1_uk_U592 (.ZN( u1_K4_10 ) , .A( u1_uk_n1050 ) );
  AOI22_X1 u1_uk_U593 (.B2( u1_uk_K_r2_26 ) , .A2( u1_uk_K_r2_6 ) , .ZN( u1_uk_n1050 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U605 (.ZN( u1_K9_22 ) , .A( u1_uk_n1157 ) );
  AOI22_X1 u1_uk_U606 (.B2( u1_uk_K_r7_41 ) , .A2( u1_uk_K_r7_48 ) , .ZN( u1_uk_n1157 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U617 (.ZN( u1_K15_35 ) , .B2( u1_uk_n1860 ) , .A2( u1_uk_n1875 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U626 (.ZN( u1_K6_35 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1469 ) , .A2( u1_uk_n1476 ) , .A1( u1_uk_n203 ) );
  INV_X1 u1_uk_U627 (.ZN( u1_K5_35 ) , .A( u1_uk_n1079 ) );
  AOI22_X1 u1_uk_U628 (.B2( u1_uk_K_r3_29 ) , .A2( u1_uk_K_r3_38 ) , .ZN( u1_uk_n1079 ) , .B1( u1_uk_n251 ) , .A1( u1_uk_n31 ) );
  INV_X1 u1_uk_U631 (.ZN( u1_K1_35 ) , .A( u1_uk_n1012 ) );
  AOI22_X1 u1_uk_U632 (.B2( u1_key_r_28 ) , .A2( u1_key_r_35 ) , .ZN( u1_uk_n1012 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U653 (.ZN( u1_K1_45 ) , .B2( u1_uk_n1201 ) , .A2( u1_uk_n1208 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n242 ) );
  INV_X1 u1_uk_U654 (.A( u1_key_r_44 ) , .ZN( u1_uk_n1208 ) );
  OAI22_X1 u1_uk_U663 (.ZN( u1_K4_7 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1353 ) , .B2( u1_uk_n1357 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U676 (.ZN( u1_K10_43 ) , .A2( u1_uk_n1623 ) , .B2( u1_uk_n1651 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U677 (.ZN( u1_K10_45 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1628 ) , .A2( u1_uk_n1644 ) , .A1( u1_uk_n238 ) );
  INV_X1 u1_uk_U713 (.ZN( u1_K1_25 ) , .A( u1_uk_n1005 ) );
  AOI22_X1 u1_uk_U714 (.B2( u1_key_r_29 ) , .A2( u1_key_r_36 ) , .ZN( u1_uk_n1005 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U727 (.ZN( u1_K6_32 ) , .B2( u1_uk_n1448 ) , .A2( u1_uk_n1464 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U729 (.ZN( u1_K5_32 ) , .B2( u1_uk_n1408 ) , .A2( u1_uk_n1412 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U732 (.ZN( u1_K15_42 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1879 ) , .A2( u1_uk_n1885 ) , .B1( u1_uk_n231 ) );
  INV_X1 u1_uk_U746 (.ZN( u1_K1_42 ) , .A( u1_uk_n1016 ) );
  AOI22_X1 u1_uk_U747 (.B2( u1_key_r_31 ) , .A2( u1_key_r_38 ) , .ZN( u1_uk_n1016 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U75 (.ZN( u1_K15_34 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1856 ) , .A2( u1_uk_n1884 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U758 (.ZN( u1_K6_13 ) , .B2( u1_uk_n1462 ) , .A2( u1_uk_n1466 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U761 (.ZN( u1_K9_13 ) , .A( u1_uk_n1150 ) , .B2( u1_uk_n1579 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U762 (.A1( u1_uk_K_r7_5 ) , .ZN( u1_uk_n1150 ) , .A2( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U768 (.ZN( u1_K9_21 ) , .B2( u1_uk_n1598 ) , .A2( u1_uk_n1603 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n83 ) );
  INV_X1 u1_uk_U785 (.ZN( u1_K6_21 ) , .A( u1_uk_n1092 ) );
  AOI22_X1 u1_uk_U786 (.B2( u1_uk_K_r4_11 ) , .A2( u1_uk_K_r4_5 ) , .ZN( u1_uk_n1092 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U789 (.ZN( u1_K6_27 ) , .B2( u1_uk_n1459 ) , .A2( u1_uk_n1464 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U79 (.ZN( u1_K6_34 ) , .A( u1_uk_n1097 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1471 ) );
  INV_X1 u1_uk_U798 (.ZN( u1_K1_27 ) , .A( u1_uk_n1007 ) );
  AOI22_X1 u1_uk_U799 (.B2( u1_key_r_14 ) , .A2( u1_key_r_21 ) , .ZN( u1_uk_n1007 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n257 ) );
  NAND2_X1 u1_uk_U80 (.A1( u1_uk_K_r4_49 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1097 ) );
  OAI22_X1 u1_uk_U805 (.ZN( u1_K6_1 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1462 ) , .A2( u1_uk_n1478 ) , .B1( u1_uk_n188 ) );
  INV_X1 u1_uk_U806 (.ZN( u1_K9_1 ) , .A( u1_uk_n1155 ) );
  AOI22_X1 u1_uk_U807 (.B2( u1_uk_K_r7_24 ) , .A2( u1_uk_K_r7_6 ) , .ZN( u1_uk_n1155 ) , .B1( u1_uk_n155 ) , .A1( u1_uk_n250 ) );
  INV_X1 u1_uk_U831 (.ZN( u1_K9_18 ) , .A( u1_uk_n1153 ) );
  AOI22_X1 u1_uk_U832 (.B2( u1_uk_K_r7_39 ) , .A2( u1_uk_K_r7_46 ) , .ZN( u1_uk_n1153 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n230 ) );
  INV_X1 u1_uk_U833 (.ZN( u1_K6_18 ) , .A( u1_uk_n1090 ) );
  AOI22_X1 u1_uk_U834 (.B2( u1_uk_K_r4_11 ) , .A2( u1_uk_K_r4_17 ) , .ZN( u1_uk_n1090 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U846 (.ZN( u1_K1_43 ) , .A2( u1_uk_n1179 ) , .B2( u1_uk_n1182 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n60 ) );
  AOI22_X1 u1_uk_U859 (.B2( u1_uk_K_r7_20 ) , .A2( u1_uk_K_r7_27 ) , .ZN( u1_uk_n1160 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U871 (.ZN( u1_K6_22 ) , .B2( u1_uk_n1447 ) , .A2( u1_uk_n1452 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U876 (.ZN( u1_K5_34 ) , .B1( u1_uk_n118 ) , .A2( u1_uk_n1401 ) , .B2( u1_uk_n1414 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U879 (.ZN( u1_K6_5 ) , .B2( u1_uk_n1452 ) , .A2( u1_uk_n1456 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U883 (.B1( n116 ) , .ZN( u1_K4_11 ) , .B2( u1_uk_n1363 ) , .A2( u1_uk_n1391 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U885 (.ZN( u1_K15_45 ) , .B2( u1_uk_n1867 ) , .A2( u1_uk_n1885 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U893 (.ZN( u1_K9_3 ) , .B1( u1_uk_n147 ) , .A2( u1_uk_n1573 ) , .B2( u1_uk_n1577 ) , .A1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U894 (.ZN( u1_K9_7 ) , .B1( u1_uk_n146 ) , .A2( u1_uk_n1574 ) , .B2( u1_uk_n1578 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U900 (.ZN( u1_K6_24 ) , .B2( u1_uk_n1457 ) , .A2( u1_uk_n1461 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U903 (.ZN( u1_K9_24 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1574 ) , .A2( u1_uk_n1616 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U917 (.ZN( u1_K6_30 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1438 ) , .A2( u1_uk_n1443 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U922 (.ZN( u1_K6_42 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1468 ) , .A2( u1_uk_n1475 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U923 (.ZN( u1_K6_39 ) , .A2( u1_uk_n1441 ) , .B2( u1_uk_n1460 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U929 (.ZN( u1_K9_23 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1584 ) , .A2( u1_uk_n1592 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U935 (.ZN( u1_K9_6 ) , .B2( u1_uk_n1585 ) , .A2( u1_uk_n1593 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U936 (.ZN( u1_K9_8 ) , .B2( u1_uk_n1603 ) , .A2( u1_uk_n1610 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U945 (.ZN( u1_K15_47 ) , .B2( u1_uk_n1854 ) , .A2( u1_uk_n1886 ) , .B1( u1_uk_n208 ) , .A1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U947 (.ZN( u1_K10_46 ) , .B2( u1_uk_n1632 ) , .A2( u1_uk_n1641 ) , .B1( u1_uk_n279 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U952 (.ZN( u1_K9_4 ) , .A1( u1_uk_n10 ) , .B2( u1_uk_n1579 ) , .A2( u1_uk_n1586 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U957 (.ZN( u1_K6_20 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1439 ) , .B2( u1_uk_n1444 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U965 (.ZN( u1_K6_36 ) , .A1( u1_uk_n11 ) , .A2( u1_uk_n1441 ) , .B2( u1_uk_n1449 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U981 (.ZN( u1_K6_3 ) , .B2( u1_uk_n1447 ) , .A2( u1_uk_n1461 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U986 (.ZN( u1_K9_15 ) , .B2( u1_uk_n1577 ) , .A2( u1_uk_n1584 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U987 (.ZN( u1_K6_15 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1453 ) , .A2( u1_uk_n1465 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U988 (.ZN( u1_K6_25 ) , .B2( u1_uk_n1454 ) , .A2( u1_uk_n1470 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U991 (.ZN( u1_K1_34 ) , .B2( u1_uk_n1174 ) , .A2( u1_uk_n1179 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U992 (.ZN( u1_K1_47 ) , .B2( u1_uk_n1172 ) , .A2( u1_uk_n1177 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n242 ) );
  XOR2_X1 u2_U181 (.B( u2_L0_6 ) , .Z( u2_N37 ) , .A( u2_out1_6 ) );
  XOR2_X1 u2_U273 (.B( u2_L7_32 ) , .Z( u2_N287 ) , .A( u2_out8_32 ) );
  XOR2_X1 u2_U276 (.B( u2_L7_29 ) , .Z( u2_N284 ) , .A( u2_out8_29 ) );
  XOR2_X1 u2_U284 (.B( u2_L7_22 ) , .Z( u2_N277 ) , .A( u2_out8_22 ) );
  XOR2_X1 u2_U287 (.B( u2_L7_19 ) , .Z( u2_N274 ) , .A( u2_out8_19 ) );
  XOR2_X1 u2_U295 (.B( u2_L7_12 ) , .Z( u2_N267 ) , .A( u2_out8_12 ) );
  XOR2_X1 u2_U296 (.B( u2_L7_11 ) , .Z( u2_N266 ) , .A( u2_out8_11 ) );
  XOR2_X1 u2_U300 (.B( u2_L7_7 ) , .Z( u2_N262 ) , .A( u2_out8_7 ) );
  XOR2_X1 u2_U304 (.B( u2_L7_4 ) , .Z( u2_N259 ) , .A( u2_out8_4 ) );
  XOR2_X1 u2_U44 (.B( u2_L0_30 ) , .Z( u2_N61 ) , .A( u2_out1_30 ) );
  XOR2_X1 u2_U51 (.B( u2_L0_24 ) , .Z( u2_N55 ) , .A( u2_out1_24 ) );
  XOR2_X1 u2_U70 (.B( u2_L0_16 ) , .Z( u2_N47 ) , .A( u2_out1_16 ) );
  XOR2_X1 u2_u1_U40 (.B( u2_K2_18 ) , .A( u2_R0_13 ) , .Z( u2_u1_X_18 ) );
  XOR2_X1 u2_u1_U41 (.B( u2_K2_17 ) , .A( u2_R0_12 ) , .Z( u2_u1_X_17 ) );
  XOR2_X1 u2_u1_U42 (.B( u2_K2_16 ) , .A( u2_R0_11 ) , .Z( u2_u1_X_16 ) );
  XOR2_X1 u2_u1_U43 (.B( u2_K2_15 ) , .A( u2_R0_10 ) , .Z( u2_u1_X_15 ) );
  XOR2_X1 u2_u1_U44 (.B( u2_K2_14 ) , .A( u2_R0_9 ) , .Z( u2_u1_X_14 ) );
  XOR2_X1 u2_u1_U45 (.B( u2_K2_13 ) , .A( u2_R0_8 ) , .Z( u2_u1_X_13 ) );
  OAI22_X1 u2_u1_u2_U10 (.ZN( u2_u1_u2_n109 ) , .A2( u2_u1_u2_n113 ) , .B2( u2_u1_u2_n133 ) , .B1( u2_u1_u2_n167 ) , .A1( u2_u1_u2_n168 ) );
  NAND3_X1 u2_u1_u2_U100 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n104 ) , .A3( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n98 ) );
  OAI22_X1 u2_u1_u2_U11 (.B1( u2_u1_u2_n151 ) , .A2( u2_u1_u2_n152 ) , .A1( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n160 ) , .B2( u2_u1_u2_n168 ) );
  NOR3_X1 u2_u1_u2_U12 (.A1( u2_u1_u2_n150 ) , .ZN( u2_u1_u2_n151 ) , .A3( u2_u1_u2_n175 ) , .A2( u2_u1_u2_n188 ) );
  AOI21_X1 u2_u1_u2_U13 (.ZN( u2_u1_u2_n144 ) , .B2( u2_u1_u2_n155 ) , .A( u2_u1_u2_n172 ) , .B1( u2_u1_u2_n185 ) );
  AOI21_X1 u2_u1_u2_U14 (.B2( u2_u1_u2_n143 ) , .ZN( u2_u1_u2_n145 ) , .B1( u2_u1_u2_n152 ) , .A( u2_u1_u2_n171 ) );
  AOI21_X1 u2_u1_u2_U15 (.B2( u2_u1_u2_n120 ) , .B1( u2_u1_u2_n121 ) , .ZN( u2_u1_u2_n126 ) , .A( u2_u1_u2_n167 ) );
  INV_X1 u2_u1_u2_U16 (.A( u2_u1_u2_n156 ) , .ZN( u2_u1_u2_n171 ) );
  INV_X1 u2_u1_u2_U17 (.A( u2_u1_u2_n120 ) , .ZN( u2_u1_u2_n188 ) );
  NAND2_X1 u2_u1_u2_U18 (.A2( u2_u1_u2_n122 ) , .ZN( u2_u1_u2_n150 ) , .A1( u2_u1_u2_n152 ) );
  INV_X1 u2_u1_u2_U19 (.A( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n170 ) );
  INV_X1 u2_u1_u2_U20 (.A( u2_u1_u2_n137 ) , .ZN( u2_u1_u2_n173 ) );
  NAND2_X1 u2_u1_u2_U21 (.A1( u2_u1_u2_n132 ) , .A2( u2_u1_u2_n139 ) , .ZN( u2_u1_u2_n157 ) );
  INV_X1 u2_u1_u2_U22 (.A( u2_u1_u2_n113 ) , .ZN( u2_u1_u2_n178 ) );
  INV_X1 u2_u1_u2_U23 (.A( u2_u1_u2_n139 ) , .ZN( u2_u1_u2_n175 ) );
  INV_X1 u2_u1_u2_U24 (.A( u2_u1_u2_n155 ) , .ZN( u2_u1_u2_n181 ) );
  INV_X1 u2_u1_u2_U25 (.A( u2_u1_u2_n119 ) , .ZN( u2_u1_u2_n177 ) );
  INV_X1 u2_u1_u2_U26 (.A( u2_u1_u2_n116 ) , .ZN( u2_u1_u2_n180 ) );
  INV_X1 u2_u1_u2_U27 (.A( u2_u1_u2_n131 ) , .ZN( u2_u1_u2_n179 ) );
  INV_X1 u2_u1_u2_U28 (.A( u2_u1_u2_n154 ) , .ZN( u2_u1_u2_n176 ) );
  NAND2_X1 u2_u1_u2_U29 (.A2( u2_u1_u2_n116 ) , .A1( u2_u1_u2_n117 ) , .ZN( u2_u1_u2_n118 ) );
  NOR2_X1 u2_u1_u2_U3 (.ZN( u2_u1_u2_n121 ) , .A2( u2_u1_u2_n177 ) , .A1( u2_u1_u2_n180 ) );
  INV_X1 u2_u1_u2_U30 (.A( u2_u1_u2_n132 ) , .ZN( u2_u1_u2_n182 ) );
  INV_X1 u2_u1_u2_U31 (.A( u2_u1_u2_n158 ) , .ZN( u2_u1_u2_n183 ) );
  OAI21_X1 u2_u1_u2_U32 (.A( u2_u1_u2_n156 ) , .B1( u2_u1_u2_n157 ) , .ZN( u2_u1_u2_n158 ) , .B2( u2_u1_u2_n179 ) );
  NOR2_X1 u2_u1_u2_U33 (.ZN( u2_u1_u2_n156 ) , .A1( u2_u1_u2_n166 ) , .A2( u2_u1_u2_n169 ) );
  NOR2_X1 u2_u1_u2_U34 (.A2( u2_u1_u2_n114 ) , .ZN( u2_u1_u2_n137 ) , .A1( u2_u1_u2_n140 ) );
  NOR2_X1 u2_u1_u2_U35 (.A2( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n153 ) , .A1( u2_u1_u2_n156 ) );
  AOI211_X1 u2_u1_u2_U36 (.ZN( u2_u1_u2_n130 ) , .C1( u2_u1_u2_n138 ) , .C2( u2_u1_u2_n179 ) , .B( u2_u1_u2_n96 ) , .A( u2_u1_u2_n97 ) );
  OAI22_X1 u2_u1_u2_U37 (.B1( u2_u1_u2_n133 ) , .A2( u2_u1_u2_n137 ) , .A1( u2_u1_u2_n152 ) , .B2( u2_u1_u2_n168 ) , .ZN( u2_u1_u2_n97 ) );
  OAI221_X1 u2_u1_u2_U38 (.B1( u2_u1_u2_n113 ) , .C1( u2_u1_u2_n132 ) , .A( u2_u1_u2_n149 ) , .B2( u2_u1_u2_n171 ) , .C2( u2_u1_u2_n172 ) , .ZN( u2_u1_u2_n96 ) );
  OAI221_X1 u2_u1_u2_U39 (.A( u2_u1_u2_n115 ) , .C2( u2_u1_u2_n123 ) , .B2( u2_u1_u2_n143 ) , .B1( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n163 ) , .C1( u2_u1_u2_n168 ) );
  INV_X1 u2_u1_u2_U4 (.A( u2_u1_u2_n134 ) , .ZN( u2_u1_u2_n185 ) );
  OAI21_X1 u2_u1_u2_U40 (.A( u2_u1_u2_n114 ) , .ZN( u2_u1_u2_n115 ) , .B1( u2_u1_u2_n176 ) , .B2( u2_u1_u2_n178 ) );
  OAI221_X1 u2_u1_u2_U41 (.A( u2_u1_u2_n135 ) , .B2( u2_u1_u2_n136 ) , .B1( u2_u1_u2_n137 ) , .ZN( u2_u1_u2_n162 ) , .C2( u2_u1_u2_n167 ) , .C1( u2_u1_u2_n185 ) );
  AND3_X1 u2_u1_u2_U42 (.A3( u2_u1_u2_n131 ) , .A2( u2_u1_u2_n132 ) , .A1( u2_u1_u2_n133 ) , .ZN( u2_u1_u2_n136 ) );
  AOI22_X1 u2_u1_u2_U43 (.ZN( u2_u1_u2_n135 ) , .B1( u2_u1_u2_n140 ) , .A1( u2_u1_u2_n156 ) , .B2( u2_u1_u2_n180 ) , .A2( u2_u1_u2_n188 ) );
  AOI21_X1 u2_u1_u2_U44 (.ZN( u2_u1_u2_n149 ) , .B1( u2_u1_u2_n173 ) , .B2( u2_u1_u2_n188 ) , .A( u2_u1_u2_n95 ) );
  AND3_X1 u2_u1_u2_U45 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n104 ) , .A3( u2_u1_u2_n156 ) , .ZN( u2_u1_u2_n95 ) );
  OAI21_X1 u2_u1_u2_U46 (.A( u2_u1_u2_n101 ) , .B2( u2_u1_u2_n121 ) , .B1( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n164 ) );
  NAND2_X1 u2_u1_u2_U47 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n107 ) , .ZN( u2_u1_u2_n155 ) );
  NAND2_X1 u2_u1_u2_U48 (.A2( u2_u1_u2_n105 ) , .A1( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n143 ) );
  NAND2_X1 u2_u1_u2_U49 (.A1( u2_u1_u2_n104 ) , .A2( u2_u1_u2_n106 ) , .ZN( u2_u1_u2_n152 ) );
  INV_X1 u2_u1_u2_U5 (.A( u2_u1_u2_n150 ) , .ZN( u2_u1_u2_n184 ) );
  NAND2_X1 u2_u1_u2_U50 (.A1( u2_u1_u2_n100 ) , .A2( u2_u1_u2_n105 ) , .ZN( u2_u1_u2_n132 ) );
  INV_X1 u2_u1_u2_U51 (.A( u2_u1_u2_n140 ) , .ZN( u2_u1_u2_n168 ) );
  INV_X1 u2_u1_u2_U52 (.A( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n167 ) );
  OAI21_X1 u2_u1_u2_U53 (.A( u2_u1_u2_n141 ) , .B2( u2_u1_u2_n142 ) , .ZN( u2_u1_u2_n146 ) , .B1( u2_u1_u2_n153 ) );
  OAI21_X1 u2_u1_u2_U54 (.A( u2_u1_u2_n140 ) , .ZN( u2_u1_u2_n141 ) , .B1( u2_u1_u2_n176 ) , .B2( u2_u1_u2_n177 ) );
  NOR3_X1 u2_u1_u2_U55 (.ZN( u2_u1_u2_n142 ) , .A3( u2_u1_u2_n175 ) , .A2( u2_u1_u2_n178 ) , .A1( u2_u1_u2_n181 ) );
  NAND2_X1 u2_u1_u2_U56 (.A1( u2_u1_u2_n102 ) , .A2( u2_u1_u2_n106 ) , .ZN( u2_u1_u2_n113 ) );
  NAND2_X1 u2_u1_u2_U57 (.A1( u2_u1_u2_n106 ) , .A2( u2_u1_u2_n107 ) , .ZN( u2_u1_u2_n131 ) );
  NAND2_X1 u2_u1_u2_U58 (.A1( u2_u1_u2_n103 ) , .A2( u2_u1_u2_n107 ) , .ZN( u2_u1_u2_n139 ) );
  NAND2_X1 u2_u1_u2_U59 (.A1( u2_u1_u2_n103 ) , .A2( u2_u1_u2_n105 ) , .ZN( u2_u1_u2_n133 ) );
  NOR4_X1 u2_u1_u2_U6 (.A4( u2_u1_u2_n124 ) , .A3( u2_u1_u2_n125 ) , .A2( u2_u1_u2_n126 ) , .A1( u2_u1_u2_n127 ) , .ZN( u2_u1_u2_n128 ) );
  NAND2_X1 u2_u1_u2_U60 (.A1( u2_u1_u2_n102 ) , .A2( u2_u1_u2_n103 ) , .ZN( u2_u1_u2_n154 ) );
  NAND2_X1 u2_u1_u2_U61 (.A2( u2_u1_u2_n103 ) , .A1( u2_u1_u2_n104 ) , .ZN( u2_u1_u2_n119 ) );
  NAND2_X1 u2_u1_u2_U62 (.A2( u2_u1_u2_n107 ) , .A1( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n123 ) );
  NAND2_X1 u2_u1_u2_U63 (.A1( u2_u1_u2_n104 ) , .A2( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n122 ) );
  INV_X1 u2_u1_u2_U64 (.A( u2_u1_u2_n114 ) , .ZN( u2_u1_u2_n172 ) );
  NAND2_X1 u2_u1_u2_U65 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n102 ) , .ZN( u2_u1_u2_n116 ) );
  NAND2_X1 u2_u1_u2_U66 (.A1( u2_u1_u2_n102 ) , .A2( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n120 ) );
  NAND2_X1 u2_u1_u2_U67 (.A2( u2_u1_u2_n105 ) , .A1( u2_u1_u2_n106 ) , .ZN( u2_u1_u2_n117 ) );
  INV_X1 u2_u1_u2_U68 (.ZN( u2_u1_u2_n187 ) , .A( u2_u1_u2_n99 ) );
  OAI21_X1 u2_u1_u2_U69 (.B1( u2_u1_u2_n137 ) , .B2( u2_u1_u2_n143 ) , .A( u2_u1_u2_n98 ) , .ZN( u2_u1_u2_n99 ) );
  AOI21_X1 u2_u1_u2_U7 (.B2( u2_u1_u2_n119 ) , .ZN( u2_u1_u2_n127 ) , .A( u2_u1_u2_n137 ) , .B1( u2_u1_u2_n155 ) );
  NOR2_X1 u2_u1_u2_U70 (.A2( u2_u1_X_16 ) , .ZN( u2_u1_u2_n140 ) , .A1( u2_u1_u2_n166 ) );
  NOR2_X1 u2_u1_u2_U71 (.A2( u2_u1_X_13 ) , .A1( u2_u1_X_14 ) , .ZN( u2_u1_u2_n100 ) );
  NOR2_X1 u2_u1_u2_U72 (.A2( u2_u1_X_16 ) , .A1( u2_u1_X_17 ) , .ZN( u2_u1_u2_n138 ) );
  NOR2_X1 u2_u1_u2_U73 (.A2( u2_u1_X_15 ) , .A1( u2_u1_X_18 ) , .ZN( u2_u1_u2_n104 ) );
  NOR2_X1 u2_u1_u2_U74 (.A2( u2_u1_X_14 ) , .ZN( u2_u1_u2_n103 ) , .A1( u2_u1_u2_n174 ) );
  NOR2_X1 u2_u1_u2_U75 (.A2( u2_u1_X_15 ) , .ZN( u2_u1_u2_n102 ) , .A1( u2_u1_u2_n165 ) );
  NOR2_X1 u2_u1_u2_U76 (.A2( u2_u1_X_17 ) , .ZN( u2_u1_u2_n114 ) , .A1( u2_u1_u2_n169 ) );
  AND2_X1 u2_u1_u2_U77 (.A1( u2_u1_X_15 ) , .ZN( u2_u1_u2_n105 ) , .A2( u2_u1_u2_n165 ) );
  AND2_X1 u2_u1_u2_U78 (.A2( u2_u1_X_15 ) , .A1( u2_u1_X_18 ) , .ZN( u2_u1_u2_n107 ) );
  AND2_X1 u2_u1_u2_U79 (.A1( u2_u1_X_14 ) , .ZN( u2_u1_u2_n106 ) , .A2( u2_u1_u2_n174 ) );
  AOI21_X1 u2_u1_u2_U8 (.ZN( u2_u1_u2_n124 ) , .B1( u2_u1_u2_n131 ) , .B2( u2_u1_u2_n143 ) , .A( u2_u1_u2_n172 ) );
  AND2_X1 u2_u1_u2_U80 (.A1( u2_u1_X_13 ) , .A2( u2_u1_X_14 ) , .ZN( u2_u1_u2_n108 ) );
  INV_X1 u2_u1_u2_U81 (.A( u2_u1_X_16 ) , .ZN( u2_u1_u2_n169 ) );
  INV_X1 u2_u1_u2_U82 (.A( u2_u1_X_17 ) , .ZN( u2_u1_u2_n166 ) );
  INV_X1 u2_u1_u2_U83 (.A( u2_u1_X_13 ) , .ZN( u2_u1_u2_n174 ) );
  INV_X1 u2_u1_u2_U84 (.A( u2_u1_X_18 ) , .ZN( u2_u1_u2_n165 ) );
  NAND4_X1 u2_u1_u2_U85 (.ZN( u2_out1_30 ) , .A4( u2_u1_u2_n147 ) , .A3( u2_u1_u2_n148 ) , .A2( u2_u1_u2_n149 ) , .A1( u2_u1_u2_n187 ) );
  NOR3_X1 u2_u1_u2_U86 (.A3( u2_u1_u2_n144 ) , .A2( u2_u1_u2_n145 ) , .A1( u2_u1_u2_n146 ) , .ZN( u2_u1_u2_n147 ) );
  AOI21_X1 u2_u1_u2_U87 (.B2( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n148 ) , .A( u2_u1_u2_n162 ) , .B1( u2_u1_u2_n182 ) );
  NAND4_X1 u2_u1_u2_U88 (.ZN( u2_out1_24 ) , .A4( u2_u1_u2_n111 ) , .A3( u2_u1_u2_n112 ) , .A1( u2_u1_u2_n130 ) , .A2( u2_u1_u2_n187 ) );
  AOI221_X1 u2_u1_u2_U89 (.A( u2_u1_u2_n109 ) , .B1( u2_u1_u2_n110 ) , .ZN( u2_u1_u2_n111 ) , .C1( u2_u1_u2_n134 ) , .C2( u2_u1_u2_n170 ) , .B2( u2_u1_u2_n173 ) );
  AOI21_X1 u2_u1_u2_U9 (.B2( u2_u1_u2_n123 ) , .ZN( u2_u1_u2_n125 ) , .A( u2_u1_u2_n171 ) , .B1( u2_u1_u2_n184 ) );
  AOI21_X1 u2_u1_u2_U90 (.ZN( u2_u1_u2_n112 ) , .B2( u2_u1_u2_n156 ) , .A( u2_u1_u2_n164 ) , .B1( u2_u1_u2_n181 ) );
  NAND4_X1 u2_u1_u2_U91 (.ZN( u2_out1_16 ) , .A4( u2_u1_u2_n128 ) , .A3( u2_u1_u2_n129 ) , .A1( u2_u1_u2_n130 ) , .A2( u2_u1_u2_n186 ) );
  AOI22_X1 u2_u1_u2_U92 (.A2( u2_u1_u2_n118 ) , .ZN( u2_u1_u2_n129 ) , .A1( u2_u1_u2_n140 ) , .B1( u2_u1_u2_n157 ) , .B2( u2_u1_u2_n170 ) );
  INV_X1 u2_u1_u2_U93 (.A( u2_u1_u2_n163 ) , .ZN( u2_u1_u2_n186 ) );
  OR4_X1 u2_u1_u2_U94 (.ZN( u2_out1_6 ) , .A4( u2_u1_u2_n161 ) , .A3( u2_u1_u2_n162 ) , .A2( u2_u1_u2_n163 ) , .A1( u2_u1_u2_n164 ) );
  OR3_X1 u2_u1_u2_U95 (.A2( u2_u1_u2_n159 ) , .A1( u2_u1_u2_n160 ) , .ZN( u2_u1_u2_n161 ) , .A3( u2_u1_u2_n183 ) );
  AOI21_X1 u2_u1_u2_U96 (.B2( u2_u1_u2_n154 ) , .B1( u2_u1_u2_n155 ) , .ZN( u2_u1_u2_n159 ) , .A( u2_u1_u2_n167 ) );
  NAND3_X1 u2_u1_u2_U97 (.A2( u2_u1_u2_n117 ) , .A1( u2_u1_u2_n122 ) , .A3( u2_u1_u2_n123 ) , .ZN( u2_u1_u2_n134 ) );
  NAND3_X1 u2_u1_u2_U98 (.ZN( u2_u1_u2_n110 ) , .A2( u2_u1_u2_n131 ) , .A3( u2_u1_u2_n139 ) , .A1( u2_u1_u2_n154 ) );
  NAND3_X1 u2_u1_u2_U99 (.A2( u2_u1_u2_n100 ) , .ZN( u2_u1_u2_n101 ) , .A1( u2_u1_u2_n104 ) , .A3( u2_u1_u2_n114 ) );
  XOR2_X1 u2_u8_U13 (.B( u2_K9_42 ) , .A( u2_R7_29 ) , .Z( u2_u8_X_42 ) );
  XOR2_X1 u2_u8_U14 (.B( u2_K9_41 ) , .A( u2_R7_28 ) , .Z( u2_u8_X_41 ) );
  XOR2_X1 u2_u8_U15 (.B( u2_K9_40 ) , .A( u2_R7_27 ) , .Z( u2_u8_X_40 ) );
  XOR2_X1 u2_u8_U17 (.B( u2_K9_39 ) , .A( u2_R7_26 ) , .Z( u2_u8_X_39 ) );
  XOR2_X1 u2_u8_U18 (.B( u2_K9_38 ) , .A( u2_R7_25 ) , .Z( u2_u8_X_38 ) );
  XOR2_X1 u2_u8_U19 (.B( u2_K9_37 ) , .A( u2_R7_24 ) , .Z( u2_u8_X_37 ) );
  XOR2_X1 u2_u8_U20 (.B( u2_K9_36 ) , .A( u2_R7_25 ) , .Z( u2_u8_X_36 ) );
  XOR2_X1 u2_u8_U21 (.B( u2_K9_35 ) , .A( u2_R7_24 ) , .Z( u2_u8_X_35 ) );
  XOR2_X1 u2_u8_U22 (.B( u2_K9_34 ) , .A( u2_R7_23 ) , .Z( u2_u8_X_34 ) );
  XOR2_X1 u2_u8_U23 (.B( u2_K9_33 ) , .A( u2_R7_22 ) , .Z( u2_u8_X_33 ) );
  XOR2_X1 u2_u8_U24 (.B( u2_K9_32 ) , .A( u2_R7_21 ) , .Z( u2_u8_X_32 ) );
  XOR2_X1 u2_u8_U25 (.B( u2_K9_31 ) , .A( u2_R7_20 ) , .Z( u2_u8_X_31 ) );
  NOR2_X1 u2_u8_u5_U10 (.ZN( u2_u8_u5_n135 ) , .A1( u2_u8_u5_n173 ) , .A2( u2_u8_u5_n176 ) );
  NOR3_X1 u2_u8_u5_U100 (.A3( u2_u8_u5_n141 ) , .A1( u2_u8_u5_n142 ) , .ZN( u2_u8_u5_n143 ) , .A2( u2_u8_u5_n191 ) );
  NAND4_X1 u2_u8_u5_U101 (.ZN( u2_out8_4 ) , .A4( u2_u8_u5_n112 ) , .A2( u2_u8_u5_n113 ) , .A1( u2_u8_u5_n114 ) , .A3( u2_u8_u5_n195 ) );
  AOI211_X1 u2_u8_u5_U102 (.A( u2_u8_u5_n110 ) , .C1( u2_u8_u5_n111 ) , .ZN( u2_u8_u5_n112 ) , .B( u2_u8_u5_n118 ) , .C2( u2_u8_u5_n177 ) );
  INV_X1 u2_u8_u5_U103 (.A( u2_u8_u5_n102 ) , .ZN( u2_u8_u5_n195 ) );
  NAND3_X1 u2_u8_u5_U104 (.A2( u2_u8_u5_n154 ) , .A3( u2_u8_u5_n158 ) , .A1( u2_u8_u5_n161 ) , .ZN( u2_u8_u5_n99 ) );
  INV_X1 u2_u8_u5_U11 (.A( u2_u8_u5_n121 ) , .ZN( u2_u8_u5_n177 ) );
  NOR2_X1 u2_u8_u5_U12 (.ZN( u2_u8_u5_n160 ) , .A2( u2_u8_u5_n173 ) , .A1( u2_u8_u5_n177 ) );
  INV_X1 u2_u8_u5_U13 (.A( u2_u8_u5_n150 ) , .ZN( u2_u8_u5_n174 ) );
  AOI21_X1 u2_u8_u5_U14 (.A( u2_u8_u5_n160 ) , .B2( u2_u8_u5_n161 ) , .ZN( u2_u8_u5_n162 ) , .B1( u2_u8_u5_n192 ) );
  INV_X1 u2_u8_u5_U15 (.A( u2_u8_u5_n159 ) , .ZN( u2_u8_u5_n192 ) );
  AOI21_X1 u2_u8_u5_U16 (.A( u2_u8_u5_n156 ) , .B2( u2_u8_u5_n157 ) , .B1( u2_u8_u5_n158 ) , .ZN( u2_u8_u5_n163 ) );
  AOI21_X1 u2_u8_u5_U17 (.B2( u2_u8_u5_n139 ) , .B1( u2_u8_u5_n140 ) , .ZN( u2_u8_u5_n141 ) , .A( u2_u8_u5_n150 ) );
  OAI21_X1 u2_u8_u5_U18 (.A( u2_u8_u5_n133 ) , .B2( u2_u8_u5_n134 ) , .B1( u2_u8_u5_n135 ) , .ZN( u2_u8_u5_n142 ) );
  OAI21_X1 u2_u8_u5_U19 (.ZN( u2_u8_u5_n133 ) , .B2( u2_u8_u5_n147 ) , .A( u2_u8_u5_n173 ) , .B1( u2_u8_u5_n188 ) );
  NAND2_X1 u2_u8_u5_U20 (.A2( u2_u8_u5_n119 ) , .A1( u2_u8_u5_n123 ) , .ZN( u2_u8_u5_n137 ) );
  INV_X1 u2_u8_u5_U21 (.A( u2_u8_u5_n155 ) , .ZN( u2_u8_u5_n194 ) );
  NAND2_X1 u2_u8_u5_U22 (.A1( u2_u8_u5_n121 ) , .ZN( u2_u8_u5_n132 ) , .A2( u2_u8_u5_n172 ) );
  NAND2_X1 u2_u8_u5_U23 (.A2( u2_u8_u5_n122 ) , .ZN( u2_u8_u5_n136 ) , .A1( u2_u8_u5_n154 ) );
  NAND2_X1 u2_u8_u5_U24 (.A2( u2_u8_u5_n119 ) , .A1( u2_u8_u5_n120 ) , .ZN( u2_u8_u5_n159 ) );
  INV_X1 u2_u8_u5_U25 (.A( u2_u8_u5_n156 ) , .ZN( u2_u8_u5_n175 ) );
  INV_X1 u2_u8_u5_U26 (.A( u2_u8_u5_n158 ) , .ZN( u2_u8_u5_n188 ) );
  INV_X1 u2_u8_u5_U27 (.A( u2_u8_u5_n152 ) , .ZN( u2_u8_u5_n179 ) );
  INV_X1 u2_u8_u5_U28 (.A( u2_u8_u5_n140 ) , .ZN( u2_u8_u5_n182 ) );
  INV_X1 u2_u8_u5_U29 (.A( u2_u8_u5_n151 ) , .ZN( u2_u8_u5_n183 ) );
  NOR2_X1 u2_u8_u5_U3 (.ZN( u2_u8_u5_n134 ) , .A1( u2_u8_u5_n183 ) , .A2( u2_u8_u5_n190 ) );
  INV_X1 u2_u8_u5_U30 (.A( u2_u8_u5_n123 ) , .ZN( u2_u8_u5_n185 ) );
  INV_X1 u2_u8_u5_U31 (.A( u2_u8_u5_n161 ) , .ZN( u2_u8_u5_n184 ) );
  INV_X1 u2_u8_u5_U32 (.A( u2_u8_u5_n139 ) , .ZN( u2_u8_u5_n189 ) );
  INV_X1 u2_u8_u5_U33 (.A( u2_u8_u5_n157 ) , .ZN( u2_u8_u5_n190 ) );
  INV_X1 u2_u8_u5_U34 (.A( u2_u8_u5_n120 ) , .ZN( u2_u8_u5_n193 ) );
  NAND2_X1 u2_u8_u5_U35 (.ZN( u2_u8_u5_n111 ) , .A1( u2_u8_u5_n140 ) , .A2( u2_u8_u5_n155 ) );
  NOR2_X1 u2_u8_u5_U36 (.ZN( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n170 ) , .A2( u2_u8_u5_n180 ) );
  INV_X1 u2_u8_u5_U37 (.A( u2_u8_u5_n117 ) , .ZN( u2_u8_u5_n196 ) );
  OAI221_X1 u2_u8_u5_U38 (.A( u2_u8_u5_n116 ) , .ZN( u2_u8_u5_n117 ) , .B2( u2_u8_u5_n119 ) , .C1( u2_u8_u5_n153 ) , .C2( u2_u8_u5_n158 ) , .B1( u2_u8_u5_n172 ) );
  AOI222_X1 u2_u8_u5_U39 (.ZN( u2_u8_u5_n116 ) , .B2( u2_u8_u5_n145 ) , .C1( u2_u8_u5_n148 ) , .A2( u2_u8_u5_n174 ) , .C2( u2_u8_u5_n177 ) , .B1( u2_u8_u5_n187 ) , .A1( u2_u8_u5_n193 ) );
  INV_X1 u2_u8_u5_U4 (.A( u2_u8_u5_n138 ) , .ZN( u2_u8_u5_n191 ) );
  INV_X1 u2_u8_u5_U40 (.A( u2_u8_u5_n115 ) , .ZN( u2_u8_u5_n187 ) );
  OAI221_X1 u2_u8_u5_U41 (.A( u2_u8_u5_n101 ) , .ZN( u2_u8_u5_n102 ) , .C2( u2_u8_u5_n115 ) , .C1( u2_u8_u5_n126 ) , .B1( u2_u8_u5_n134 ) , .B2( u2_u8_u5_n160 ) );
  OAI21_X1 u2_u8_u5_U42 (.ZN( u2_u8_u5_n101 ) , .B1( u2_u8_u5_n137 ) , .A( u2_u8_u5_n146 ) , .B2( u2_u8_u5_n147 ) );
  AOI22_X1 u2_u8_u5_U43 (.B2( u2_u8_u5_n131 ) , .A2( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n169 ) , .B1( u2_u8_u5_n174 ) , .A1( u2_u8_u5_n185 ) );
  NOR2_X1 u2_u8_u5_U44 (.A1( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n150 ) , .A2( u2_u8_u5_n173 ) );
  AOI21_X1 u2_u8_u5_U45 (.A( u2_u8_u5_n118 ) , .B2( u2_u8_u5_n145 ) , .ZN( u2_u8_u5_n168 ) , .B1( u2_u8_u5_n186 ) );
  INV_X1 u2_u8_u5_U46 (.A( u2_u8_u5_n122 ) , .ZN( u2_u8_u5_n186 ) );
  NOR2_X1 u2_u8_u5_U47 (.A1( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n152 ) , .A2( u2_u8_u5_n176 ) );
  NOR2_X1 u2_u8_u5_U48 (.A1( u2_u8_u5_n115 ) , .ZN( u2_u8_u5_n118 ) , .A2( u2_u8_u5_n153 ) );
  NOR2_X1 u2_u8_u5_U49 (.A2( u2_u8_u5_n145 ) , .ZN( u2_u8_u5_n156 ) , .A1( u2_u8_u5_n174 ) );
  OAI21_X1 u2_u8_u5_U5 (.B2( u2_u8_u5_n136 ) , .B1( u2_u8_u5_n137 ) , .ZN( u2_u8_u5_n138 ) , .A( u2_u8_u5_n177 ) );
  NOR2_X1 u2_u8_u5_U50 (.ZN( u2_u8_u5_n121 ) , .A2( u2_u8_u5_n145 ) , .A1( u2_u8_u5_n176 ) );
  AOI22_X1 u2_u8_u5_U51 (.ZN( u2_u8_u5_n114 ) , .A2( u2_u8_u5_n137 ) , .A1( u2_u8_u5_n145 ) , .B2( u2_u8_u5_n175 ) , .B1( u2_u8_u5_n193 ) );
  OAI211_X1 u2_u8_u5_U52 (.B( u2_u8_u5_n124 ) , .A( u2_u8_u5_n125 ) , .C2( u2_u8_u5_n126 ) , .C1( u2_u8_u5_n127 ) , .ZN( u2_u8_u5_n128 ) );
  NOR3_X1 u2_u8_u5_U53 (.ZN( u2_u8_u5_n127 ) , .A1( u2_u8_u5_n136 ) , .A3( u2_u8_u5_n148 ) , .A2( u2_u8_u5_n182 ) );
  OAI21_X1 u2_u8_u5_U54 (.ZN( u2_u8_u5_n124 ) , .A( u2_u8_u5_n177 ) , .B2( u2_u8_u5_n183 ) , .B1( u2_u8_u5_n189 ) );
  OAI21_X1 u2_u8_u5_U55 (.ZN( u2_u8_u5_n125 ) , .A( u2_u8_u5_n174 ) , .B2( u2_u8_u5_n185 ) , .B1( u2_u8_u5_n190 ) );
  AOI21_X1 u2_u8_u5_U56 (.A( u2_u8_u5_n153 ) , .B2( u2_u8_u5_n154 ) , .B1( u2_u8_u5_n155 ) , .ZN( u2_u8_u5_n164 ) );
  AOI21_X1 u2_u8_u5_U57 (.ZN( u2_u8_u5_n110 ) , .B1( u2_u8_u5_n122 ) , .B2( u2_u8_u5_n139 ) , .A( u2_u8_u5_n153 ) );
  INV_X1 u2_u8_u5_U58 (.A( u2_u8_u5_n153 ) , .ZN( u2_u8_u5_n176 ) );
  INV_X1 u2_u8_u5_U59 (.A( u2_u8_u5_n126 ) , .ZN( u2_u8_u5_n173 ) );
  AOI222_X1 u2_u8_u5_U6 (.ZN( u2_u8_u5_n113 ) , .A1( u2_u8_u5_n131 ) , .C1( u2_u8_u5_n148 ) , .B2( u2_u8_u5_n174 ) , .C2( u2_u8_u5_n178 ) , .A2( u2_u8_u5_n179 ) , .B1( u2_u8_u5_n99 ) );
  AND2_X1 u2_u8_u5_U60 (.A2( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n107 ) , .ZN( u2_u8_u5_n147 ) );
  AND2_X1 u2_u8_u5_U61 (.A2( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n108 ) , .ZN( u2_u8_u5_n148 ) );
  NAND2_X1 u2_u8_u5_U62 (.A1( u2_u8_u5_n105 ) , .A2( u2_u8_u5_n106 ) , .ZN( u2_u8_u5_n158 ) );
  NAND2_X1 u2_u8_u5_U63 (.A2( u2_u8_u5_n108 ) , .A1( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n139 ) );
  NAND2_X1 u2_u8_u5_U64 (.A1( u2_u8_u5_n106 ) , .A2( u2_u8_u5_n108 ) , .ZN( u2_u8_u5_n119 ) );
  NAND2_X1 u2_u8_u5_U65 (.A2( u2_u8_u5_n103 ) , .A1( u2_u8_u5_n105 ) , .ZN( u2_u8_u5_n140 ) );
  NAND2_X1 u2_u8_u5_U66 (.A2( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n105 ) , .ZN( u2_u8_u5_n155 ) );
  NAND2_X1 u2_u8_u5_U67 (.A2( u2_u8_u5_n106 ) , .A1( u2_u8_u5_n107 ) , .ZN( u2_u8_u5_n122 ) );
  NAND2_X1 u2_u8_u5_U68 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n106 ) , .ZN( u2_u8_u5_n115 ) );
  NAND2_X1 u2_u8_u5_U69 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n103 ) , .ZN( u2_u8_u5_n161 ) );
  INV_X1 u2_u8_u5_U7 (.A( u2_u8_u5_n135 ) , .ZN( u2_u8_u5_n178 ) );
  NAND2_X1 u2_u8_u5_U70 (.A1( u2_u8_u5_n105 ) , .A2( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n154 ) );
  INV_X1 u2_u8_u5_U71 (.A( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n172 ) );
  NAND2_X1 u2_u8_u5_U72 (.A1( u2_u8_u5_n103 ) , .A2( u2_u8_u5_n108 ) , .ZN( u2_u8_u5_n123 ) );
  NAND2_X1 u2_u8_u5_U73 (.A2( u2_u8_u5_n103 ) , .A1( u2_u8_u5_n107 ) , .ZN( u2_u8_u5_n151 ) );
  NAND2_X1 u2_u8_u5_U74 (.A2( u2_u8_u5_n107 ) , .A1( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n120 ) );
  NAND2_X1 u2_u8_u5_U75 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n109 ) , .ZN( u2_u8_u5_n157 ) );
  AND2_X1 u2_u8_u5_U76 (.A2( u2_u8_u5_n100 ) , .A1( u2_u8_u5_n104 ) , .ZN( u2_u8_u5_n131 ) );
  NOR2_X1 u2_u8_u5_U77 (.A2( u2_u8_X_34 ) , .A1( u2_u8_X_35 ) , .ZN( u2_u8_u5_n145 ) );
  NOR2_X1 u2_u8_u5_U78 (.A2( u2_u8_X_34 ) , .ZN( u2_u8_u5_n146 ) , .A1( u2_u8_u5_n171 ) );
  NOR2_X1 u2_u8_u5_U79 (.A2( u2_u8_X_31 ) , .A1( u2_u8_X_32 ) , .ZN( u2_u8_u5_n103 ) );
  OAI22_X1 u2_u8_u5_U8 (.B2( u2_u8_u5_n149 ) , .B1( u2_u8_u5_n150 ) , .A2( u2_u8_u5_n151 ) , .A1( u2_u8_u5_n152 ) , .ZN( u2_u8_u5_n165 ) );
  NOR2_X1 u2_u8_u5_U80 (.A2( u2_u8_X_36 ) , .ZN( u2_u8_u5_n105 ) , .A1( u2_u8_u5_n180 ) );
  NOR2_X1 u2_u8_u5_U81 (.A2( u2_u8_X_33 ) , .ZN( u2_u8_u5_n108 ) , .A1( u2_u8_u5_n170 ) );
  NOR2_X1 u2_u8_u5_U82 (.A2( u2_u8_X_33 ) , .A1( u2_u8_X_36 ) , .ZN( u2_u8_u5_n107 ) );
  NOR2_X1 u2_u8_u5_U83 (.A2( u2_u8_X_31 ) , .ZN( u2_u8_u5_n104 ) , .A1( u2_u8_u5_n181 ) );
  NAND2_X1 u2_u8_u5_U84 (.A2( u2_u8_X_34 ) , .A1( u2_u8_X_35 ) , .ZN( u2_u8_u5_n153 ) );
  NAND2_X1 u2_u8_u5_U85 (.A1( u2_u8_X_34 ) , .ZN( u2_u8_u5_n126 ) , .A2( u2_u8_u5_n171 ) );
  AND2_X1 u2_u8_u5_U86 (.A1( u2_u8_X_31 ) , .A2( u2_u8_X_32 ) , .ZN( u2_u8_u5_n106 ) );
  AND2_X1 u2_u8_u5_U87 (.A1( u2_u8_X_31 ) , .ZN( u2_u8_u5_n109 ) , .A2( u2_u8_u5_n181 ) );
  INV_X1 u2_u8_u5_U88 (.A( u2_u8_X_33 ) , .ZN( u2_u8_u5_n180 ) );
  INV_X1 u2_u8_u5_U89 (.A( u2_u8_X_35 ) , .ZN( u2_u8_u5_n171 ) );
  NOR3_X1 u2_u8_u5_U9 (.A2( u2_u8_u5_n147 ) , .A1( u2_u8_u5_n148 ) , .ZN( u2_u8_u5_n149 ) , .A3( u2_u8_u5_n194 ) );
  INV_X1 u2_u8_u5_U90 (.A( u2_u8_X_36 ) , .ZN( u2_u8_u5_n170 ) );
  INV_X1 u2_u8_u5_U91 (.A( u2_u8_X_32 ) , .ZN( u2_u8_u5_n181 ) );
  NAND4_X1 u2_u8_u5_U92 (.ZN( u2_out8_29 ) , .A4( u2_u8_u5_n129 ) , .A3( u2_u8_u5_n130 ) , .A2( u2_u8_u5_n168 ) , .A1( u2_u8_u5_n196 ) );
  AOI221_X1 u2_u8_u5_U93 (.A( u2_u8_u5_n128 ) , .ZN( u2_u8_u5_n129 ) , .C2( u2_u8_u5_n132 ) , .B2( u2_u8_u5_n159 ) , .B1( u2_u8_u5_n176 ) , .C1( u2_u8_u5_n184 ) );
  AOI222_X1 u2_u8_u5_U94 (.ZN( u2_u8_u5_n130 ) , .A2( u2_u8_u5_n146 ) , .B1( u2_u8_u5_n147 ) , .C2( u2_u8_u5_n175 ) , .B2( u2_u8_u5_n179 ) , .A1( u2_u8_u5_n188 ) , .C1( u2_u8_u5_n194 ) );
  NAND4_X1 u2_u8_u5_U95 (.ZN( u2_out8_19 ) , .A4( u2_u8_u5_n166 ) , .A3( u2_u8_u5_n167 ) , .A2( u2_u8_u5_n168 ) , .A1( u2_u8_u5_n169 ) );
  AOI22_X1 u2_u8_u5_U96 (.B2( u2_u8_u5_n145 ) , .A2( u2_u8_u5_n146 ) , .ZN( u2_u8_u5_n167 ) , .B1( u2_u8_u5_n182 ) , .A1( u2_u8_u5_n189 ) );
  NOR4_X1 u2_u8_u5_U97 (.A4( u2_u8_u5_n162 ) , .A3( u2_u8_u5_n163 ) , .A2( u2_u8_u5_n164 ) , .A1( u2_u8_u5_n165 ) , .ZN( u2_u8_u5_n166 ) );
  NAND4_X1 u2_u8_u5_U98 (.ZN( u2_out8_11 ) , .A4( u2_u8_u5_n143 ) , .A3( u2_u8_u5_n144 ) , .A2( u2_u8_u5_n169 ) , .A1( u2_u8_u5_n196 ) );
  AOI22_X1 u2_u8_u5_U99 (.A2( u2_u8_u5_n132 ) , .ZN( u2_u8_u5_n144 ) , .B2( u2_u8_u5_n145 ) , .B1( u2_u8_u5_n184 ) , .A1( u2_u8_u5_n194 ) );
  AOI22_X1 u2_u8_u6_U10 (.A2( u2_u8_u6_n151 ) , .B2( u2_u8_u6_n161 ) , .A1( u2_u8_u6_n167 ) , .B1( u2_u8_u6_n170 ) , .ZN( u2_u8_u6_n89 ) );
  AOI21_X1 u2_u8_u6_U11 (.B1( u2_u8_u6_n107 ) , .B2( u2_u8_u6_n132 ) , .A( u2_u8_u6_n158 ) , .ZN( u2_u8_u6_n88 ) );
  AOI21_X1 u2_u8_u6_U12 (.B2( u2_u8_u6_n147 ) , .B1( u2_u8_u6_n148 ) , .ZN( u2_u8_u6_n149 ) , .A( u2_u8_u6_n158 ) );
  AOI21_X1 u2_u8_u6_U13 (.ZN( u2_u8_u6_n106 ) , .A( u2_u8_u6_n142 ) , .B2( u2_u8_u6_n159 ) , .B1( u2_u8_u6_n164 ) );
  INV_X1 u2_u8_u6_U14 (.A( u2_u8_u6_n155 ) , .ZN( u2_u8_u6_n161 ) );
  INV_X1 u2_u8_u6_U15 (.A( u2_u8_u6_n128 ) , .ZN( u2_u8_u6_n164 ) );
  NAND2_X1 u2_u8_u6_U16 (.ZN( u2_u8_u6_n110 ) , .A1( u2_u8_u6_n122 ) , .A2( u2_u8_u6_n129 ) );
  NAND2_X1 u2_u8_u6_U17 (.ZN( u2_u8_u6_n124 ) , .A2( u2_u8_u6_n146 ) , .A1( u2_u8_u6_n148 ) );
  INV_X1 u2_u8_u6_U18 (.A( u2_u8_u6_n132 ) , .ZN( u2_u8_u6_n171 ) );
  AND2_X1 u2_u8_u6_U19 (.A1( u2_u8_u6_n100 ) , .ZN( u2_u8_u6_n130 ) , .A2( u2_u8_u6_n147 ) );
  INV_X1 u2_u8_u6_U20 (.A( u2_u8_u6_n127 ) , .ZN( u2_u8_u6_n173 ) );
  INV_X1 u2_u8_u6_U21 (.A( u2_u8_u6_n121 ) , .ZN( u2_u8_u6_n167 ) );
  INV_X1 u2_u8_u6_U22 (.A( u2_u8_u6_n100 ) , .ZN( u2_u8_u6_n169 ) );
  INV_X1 u2_u8_u6_U23 (.A( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n170 ) );
  INV_X1 u2_u8_u6_U24 (.A( u2_u8_u6_n113 ) , .ZN( u2_u8_u6_n168 ) );
  AND2_X1 u2_u8_u6_U25 (.A1( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n119 ) , .ZN( u2_u8_u6_n133 ) );
  AND2_X1 u2_u8_u6_U26 (.A2( u2_u8_u6_n121 ) , .A1( u2_u8_u6_n122 ) , .ZN( u2_u8_u6_n131 ) );
  AND3_X1 u2_u8_u6_U27 (.ZN( u2_u8_u6_n120 ) , .A2( u2_u8_u6_n127 ) , .A1( u2_u8_u6_n132 ) , .A3( u2_u8_u6_n145 ) );
  INV_X1 u2_u8_u6_U28 (.A( u2_u8_u6_n146 ) , .ZN( u2_u8_u6_n163 ) );
  AOI222_X1 u2_u8_u6_U29 (.ZN( u2_u8_u6_n114 ) , .A1( u2_u8_u6_n118 ) , .A2( u2_u8_u6_n126 ) , .B2( u2_u8_u6_n151 ) , .C2( u2_u8_u6_n159 ) , .C1( u2_u8_u6_n168 ) , .B1( u2_u8_u6_n169 ) );
  INV_X1 u2_u8_u6_U3 (.A( u2_u8_u6_n110 ) , .ZN( u2_u8_u6_n166 ) );
  NOR2_X1 u2_u8_u6_U30 (.A1( u2_u8_u6_n162 ) , .A2( u2_u8_u6_n165 ) , .ZN( u2_u8_u6_n98 ) );
  AOI211_X1 u2_u8_u6_U31 (.B( u2_u8_u6_n134 ) , .A( u2_u8_u6_n135 ) , .C1( u2_u8_u6_n136 ) , .ZN( u2_u8_u6_n137 ) , .C2( u2_u8_u6_n151 ) );
  AOI21_X1 u2_u8_u6_U32 (.B2( u2_u8_u6_n132 ) , .B1( u2_u8_u6_n133 ) , .ZN( u2_u8_u6_n134 ) , .A( u2_u8_u6_n158 ) );
  NAND4_X1 u2_u8_u6_U33 (.A4( u2_u8_u6_n127 ) , .A3( u2_u8_u6_n128 ) , .A2( u2_u8_u6_n129 ) , .A1( u2_u8_u6_n130 ) , .ZN( u2_u8_u6_n136 ) );
  AOI21_X1 u2_u8_u6_U34 (.B1( u2_u8_u6_n131 ) , .ZN( u2_u8_u6_n135 ) , .A( u2_u8_u6_n144 ) , .B2( u2_u8_u6_n146 ) );
  NAND2_X1 u2_u8_u6_U35 (.A1( u2_u8_u6_n144 ) , .ZN( u2_u8_u6_n151 ) , .A2( u2_u8_u6_n158 ) );
  NAND2_X1 u2_u8_u6_U36 (.ZN( u2_u8_u6_n132 ) , .A1( u2_u8_u6_n91 ) , .A2( u2_u8_u6_n97 ) );
  AOI22_X1 u2_u8_u6_U37 (.B2( u2_u8_u6_n110 ) , .B1( u2_u8_u6_n111 ) , .A1( u2_u8_u6_n112 ) , .ZN( u2_u8_u6_n115 ) , .A2( u2_u8_u6_n161 ) );
  NAND4_X1 u2_u8_u6_U38 (.A3( u2_u8_u6_n109 ) , .ZN( u2_u8_u6_n112 ) , .A4( u2_u8_u6_n132 ) , .A2( u2_u8_u6_n147 ) , .A1( u2_u8_u6_n166 ) );
  NOR2_X1 u2_u8_u6_U39 (.ZN( u2_u8_u6_n109 ) , .A1( u2_u8_u6_n170 ) , .A2( u2_u8_u6_n173 ) );
  INV_X1 u2_u8_u6_U4 (.A( u2_u8_u6_n142 ) , .ZN( u2_u8_u6_n174 ) );
  NOR2_X1 u2_u8_u6_U40 (.A2( u2_u8_u6_n126 ) , .ZN( u2_u8_u6_n155 ) , .A1( u2_u8_u6_n160 ) );
  NAND2_X1 u2_u8_u6_U41 (.ZN( u2_u8_u6_n146 ) , .A2( u2_u8_u6_n94 ) , .A1( u2_u8_u6_n99 ) );
  AOI21_X1 u2_u8_u6_U42 (.A( u2_u8_u6_n144 ) , .B2( u2_u8_u6_n145 ) , .B1( u2_u8_u6_n146 ) , .ZN( u2_u8_u6_n150 ) );
  INV_X1 u2_u8_u6_U43 (.A( u2_u8_u6_n111 ) , .ZN( u2_u8_u6_n158 ) );
  NAND2_X1 u2_u8_u6_U44 (.ZN( u2_u8_u6_n127 ) , .A1( u2_u8_u6_n91 ) , .A2( u2_u8_u6_n92 ) );
  NAND2_X1 u2_u8_u6_U45 (.ZN( u2_u8_u6_n129 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n96 ) );
  INV_X1 u2_u8_u6_U46 (.A( u2_u8_u6_n144 ) , .ZN( u2_u8_u6_n159 ) );
  NAND2_X1 u2_u8_u6_U47 (.ZN( u2_u8_u6_n145 ) , .A2( u2_u8_u6_n97 ) , .A1( u2_u8_u6_n98 ) );
  NAND2_X1 u2_u8_u6_U48 (.ZN( u2_u8_u6_n148 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n94 ) );
  NAND2_X1 u2_u8_u6_U49 (.ZN( u2_u8_u6_n108 ) , .A2( u2_u8_u6_n139 ) , .A1( u2_u8_u6_n144 ) );
  NAND2_X1 u2_u8_u6_U5 (.A2( u2_u8_u6_n143 ) , .ZN( u2_u8_u6_n152 ) , .A1( u2_u8_u6_n166 ) );
  NAND2_X1 u2_u8_u6_U50 (.ZN( u2_u8_u6_n121 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n97 ) );
  NAND2_X1 u2_u8_u6_U51 (.ZN( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n95 ) );
  AND2_X1 u2_u8_u6_U52 (.ZN( u2_u8_u6_n118 ) , .A2( u2_u8_u6_n91 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U53 (.ZN( u2_u8_u6_n147 ) , .A2( u2_u8_u6_n98 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U54 (.ZN( u2_u8_u6_n128 ) , .A1( u2_u8_u6_n94 ) , .A2( u2_u8_u6_n96 ) );
  NAND2_X1 u2_u8_u6_U55 (.ZN( u2_u8_u6_n119 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U56 (.ZN( u2_u8_u6_n123 ) , .A2( u2_u8_u6_n91 ) , .A1( u2_u8_u6_n96 ) );
  NAND2_X1 u2_u8_u6_U57 (.ZN( u2_u8_u6_n100 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n98 ) );
  NAND2_X1 u2_u8_u6_U58 (.ZN( u2_u8_u6_n122 ) , .A1( u2_u8_u6_n94 ) , .A2( u2_u8_u6_n97 ) );
  INV_X1 u2_u8_u6_U59 (.A( u2_u8_u6_n139 ) , .ZN( u2_u8_u6_n160 ) );
  AOI22_X1 u2_u8_u6_U6 (.B2( u2_u8_u6_n101 ) , .A1( u2_u8_u6_n102 ) , .ZN( u2_u8_u6_n103 ) , .B1( u2_u8_u6_n160 ) , .A2( u2_u8_u6_n161 ) );
  NAND2_X1 u2_u8_u6_U60 (.ZN( u2_u8_u6_n113 ) , .A1( u2_u8_u6_n96 ) , .A2( u2_u8_u6_n98 ) );
  NOR2_X1 u2_u8_u6_U61 (.A2( u2_u8_X_40 ) , .A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n126 ) );
  NOR2_X1 u2_u8_u6_U62 (.A2( u2_u8_X_39 ) , .A1( u2_u8_X_42 ) , .ZN( u2_u8_u6_n92 ) );
  NOR2_X1 u2_u8_u6_U63 (.A2( u2_u8_X_39 ) , .A1( u2_u8_u6_n156 ) , .ZN( u2_u8_u6_n97 ) );
  NOR2_X1 u2_u8_u6_U64 (.A2( u2_u8_X_38 ) , .A1( u2_u8_u6_n165 ) , .ZN( u2_u8_u6_n95 ) );
  NOR2_X1 u2_u8_u6_U65 (.A2( u2_u8_X_41 ) , .ZN( u2_u8_u6_n111 ) , .A1( u2_u8_u6_n157 ) );
  NOR2_X1 u2_u8_u6_U66 (.A2( u2_u8_X_37 ) , .A1( u2_u8_u6_n162 ) , .ZN( u2_u8_u6_n94 ) );
  NOR2_X1 u2_u8_u6_U67 (.A2( u2_u8_X_37 ) , .A1( u2_u8_X_38 ) , .ZN( u2_u8_u6_n91 ) );
  NAND2_X1 u2_u8_u6_U68 (.A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n144 ) , .A2( u2_u8_u6_n157 ) );
  NAND2_X1 u2_u8_u6_U69 (.A2( u2_u8_X_40 ) , .A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n139 ) );
  NOR2_X1 u2_u8_u6_U7 (.A1( u2_u8_u6_n118 ) , .ZN( u2_u8_u6_n143 ) , .A2( u2_u8_u6_n168 ) );
  AND2_X1 u2_u8_u6_U70 (.A1( u2_u8_X_39 ) , .A2( u2_u8_u6_n156 ) , .ZN( u2_u8_u6_n96 ) );
  AND2_X1 u2_u8_u6_U71 (.A1( u2_u8_X_39 ) , .A2( u2_u8_X_42 ) , .ZN( u2_u8_u6_n99 ) );
  INV_X1 u2_u8_u6_U72 (.A( u2_u8_X_40 ) , .ZN( u2_u8_u6_n157 ) );
  INV_X1 u2_u8_u6_U73 (.A( u2_u8_X_37 ) , .ZN( u2_u8_u6_n165 ) );
  INV_X1 u2_u8_u6_U74 (.A( u2_u8_X_38 ) , .ZN( u2_u8_u6_n162 ) );
  INV_X1 u2_u8_u6_U75 (.A( u2_u8_X_42 ) , .ZN( u2_u8_u6_n156 ) );
  NAND4_X1 u2_u8_u6_U76 (.ZN( u2_out8_32 ) , .A4( u2_u8_u6_n103 ) , .A3( u2_u8_u6_n104 ) , .A2( u2_u8_u6_n105 ) , .A1( u2_u8_u6_n106 ) );
  AOI22_X1 u2_u8_u6_U77 (.ZN( u2_u8_u6_n105 ) , .A2( u2_u8_u6_n108 ) , .A1( u2_u8_u6_n118 ) , .B2( u2_u8_u6_n126 ) , .B1( u2_u8_u6_n171 ) );
  AOI22_X1 u2_u8_u6_U78 (.ZN( u2_u8_u6_n104 ) , .A1( u2_u8_u6_n111 ) , .B1( u2_u8_u6_n124 ) , .B2( u2_u8_u6_n151 ) , .A2( u2_u8_u6_n93 ) );
  NAND4_X1 u2_u8_u6_U79 (.ZN( u2_out8_12 ) , .A4( u2_u8_u6_n114 ) , .A3( u2_u8_u6_n115 ) , .A2( u2_u8_u6_n116 ) , .A1( u2_u8_u6_n117 ) );
  OAI21_X1 u2_u8_u6_U8 (.A( u2_u8_u6_n159 ) , .B1( u2_u8_u6_n169 ) , .B2( u2_u8_u6_n173 ) , .ZN( u2_u8_u6_n90 ) );
  OAI22_X1 u2_u8_u6_U80 (.B2( u2_u8_u6_n111 ) , .ZN( u2_u8_u6_n116 ) , .B1( u2_u8_u6_n126 ) , .A2( u2_u8_u6_n164 ) , .A1( u2_u8_u6_n167 ) );
  OAI21_X1 u2_u8_u6_U81 (.A( u2_u8_u6_n108 ) , .ZN( u2_u8_u6_n117 ) , .B2( u2_u8_u6_n141 ) , .B1( u2_u8_u6_n163 ) );
  OAI211_X1 u2_u8_u6_U82 (.ZN( u2_out8_7 ) , .B( u2_u8_u6_n153 ) , .C2( u2_u8_u6_n154 ) , .C1( u2_u8_u6_n155 ) , .A( u2_u8_u6_n174 ) );
  NOR3_X1 u2_u8_u6_U83 (.A1( u2_u8_u6_n141 ) , .ZN( u2_u8_u6_n154 ) , .A3( u2_u8_u6_n164 ) , .A2( u2_u8_u6_n171 ) );
  AOI211_X1 u2_u8_u6_U84 (.B( u2_u8_u6_n149 ) , .A( u2_u8_u6_n150 ) , .C2( u2_u8_u6_n151 ) , .C1( u2_u8_u6_n152 ) , .ZN( u2_u8_u6_n153 ) );
  OAI211_X1 u2_u8_u6_U85 (.ZN( u2_out8_22 ) , .B( u2_u8_u6_n137 ) , .A( u2_u8_u6_n138 ) , .C2( u2_u8_u6_n139 ) , .C1( u2_u8_u6_n140 ) );
  AOI22_X1 u2_u8_u6_U86 (.B1( u2_u8_u6_n124 ) , .A2( u2_u8_u6_n125 ) , .A1( u2_u8_u6_n126 ) , .ZN( u2_u8_u6_n138 ) , .B2( u2_u8_u6_n161 ) );
  AND4_X1 u2_u8_u6_U87 (.A3( u2_u8_u6_n119 ) , .A1( u2_u8_u6_n120 ) , .A4( u2_u8_u6_n129 ) , .ZN( u2_u8_u6_n140 ) , .A2( u2_u8_u6_n143 ) );
  NAND3_X1 u2_u8_u6_U88 (.A2( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n125 ) , .A1( u2_u8_u6_n130 ) , .A3( u2_u8_u6_n131 ) );
  NAND3_X1 u2_u8_u6_U89 (.A3( u2_u8_u6_n133 ) , .ZN( u2_u8_u6_n141 ) , .A1( u2_u8_u6_n145 ) , .A2( u2_u8_u6_n148 ) );
  INV_X1 u2_u8_u6_U9 (.ZN( u2_u8_u6_n172 ) , .A( u2_u8_u6_n88 ) );
  NAND3_X1 u2_u8_u6_U90 (.ZN( u2_u8_u6_n101 ) , .A3( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n121 ) , .A1( u2_u8_u6_n127 ) );
  NAND3_X1 u2_u8_u6_U91 (.ZN( u2_u8_u6_n102 ) , .A3( u2_u8_u6_n130 ) , .A2( u2_u8_u6_n145 ) , .A1( u2_u8_u6_n166 ) );
  NAND3_X1 u2_u8_u6_U92 (.A3( u2_u8_u6_n113 ) , .A1( u2_u8_u6_n119 ) , .A2( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n93 ) );
  NAND3_X1 u2_u8_u6_U93 (.ZN( u2_u8_u6_n142 ) , .A2( u2_u8_u6_n172 ) , .A3( u2_u8_u6_n89 ) , .A1( u2_u8_u6_n90 ) );
  OAI21_X1 u2_uk_U1009 (.ZN( u2_K9_39 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1135 ) , .B2( u2_uk_n1571 ) );
  NAND2_X1 u2_uk_U1010 (.A1( u2_uk_K_r7_31 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n1135 ) );
  OAI21_X1 u2_uk_U139 (.ZN( u2_K2_15 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1261 ) , .A( u2_uk_n994 ) );
  INV_X1 u2_uk_U184 (.ZN( u2_K2_14 ) , .A( u2_uk_n993 ) );
  AOI22_X1 u2_uk_U185 (.B2( u2_uk_K_r0_11 ) , .A2( u2_uk_K_r0_32 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n993 ) );
  OAI22_X1 u2_uk_U236 (.ZN( u2_K9_31 ) , .B2( u2_uk_n1542 ) , .A2( u2_uk_n1583 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U444 (.ZN( u2_K9_33 ) , .A( u2_uk_n1132 ) );
  OAI21_X1 u2_uk_U466 (.ZN( u2_K9_37 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1134 ) , .B2( u2_uk_n1551 ) );
  INV_X1 u2_uk_U616 (.ZN( u2_K9_35 ) , .A( u2_uk_n1133 ) );
  AOI22_X1 u2_uk_U617 (.B2( u2_uk_K_r7_16 ) , .A2( u2_uk_K_r7_23 ) , .B1( u2_uk_n102 ) , .ZN( u2_uk_n1133 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U752 (.ZN( u2_K2_13 ) , .A2( u2_uk_n1231 ) , .B2( u2_uk_n1260 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U894 (.ZN( u2_K2_17 ) , .A2( u2_uk_n1231 ) , .B2( u2_uk_n1247 ) , .A1( u2_uk_n145 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U927 (.ZN( u2_K9_34 ) , .A1( u2_uk_n100 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1551 ) , .A2( u2_uk_n1558 ) );
  INV_X1 u2_uk_U968 (.ZN( u2_K9_41 ) , .A( u2_uk_n1136 ) );
  INV_X1 u2_uk_U972 (.ZN( u2_K9_42 ) , .A( u2_uk_n1137 ) );
endmodule

