module aes_aes_die_6 ( sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa21_0, 
       sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa23_sr_0, 
        sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7 );
  input sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa21_0, 
        sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7;
  output sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa23_sr_0, 
        sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7;
  wire us12_n438, us12_n439, us12_n440, us12_n441, us12_n442, us12_n443, us12_n444, us12_n445, us12_n446, 
       us12_n447, us12_n448, us12_n449, us12_n450, us12_n451, us12_n452, us12_n453, us12_n454, us12_n455, 
       us12_n456, us12_n457, us12_n458, us12_n459, us12_n460, us12_n461, us12_n462, us12_n463, us12_n464, 
       us12_n465, us12_n466, us12_n467, us12_n468, us12_n469, us12_n470, us12_n471, us12_n472, us12_n473, 
       us12_n474, us12_n475, us12_n476, us12_n477, us12_n478, us12_n479, us12_n480, us12_n481, us12_n482, 
       us12_n483, us12_n484, us12_n485, us12_n486, us12_n487, us12_n488, us12_n489, us12_n490, us12_n491, 
       us12_n492, us12_n493, us12_n494, us12_n495, us12_n496, us12_n497, us12_n498, us12_n499, us12_n500, 
       us12_n501, us12_n502, us12_n503, us12_n504, us12_n505, us12_n506, us12_n507, us12_n508, us12_n509, 
       us12_n510, us12_n511, us12_n512, us12_n513, us12_n514, us12_n515, us12_n516, us12_n517, us12_n518, 
       us12_n519, us12_n520, us12_n521, us12_n522, us12_n523, us12_n524, us12_n525, us12_n526, us12_n527, 
       us12_n528, us12_n529, us12_n530, us12_n531, us12_n532, us12_n533, us12_n534, us12_n535, us12_n536, 
       us12_n537, us12_n538, us12_n539, us12_n540, us12_n541, us12_n542, us12_n543, us12_n544, us12_n545, 
       us12_n546, us12_n547, us12_n548, us12_n549, us12_n550, us12_n551, us12_n552, us12_n553, us12_n554, 
       us12_n555, us12_n556, us12_n557, us12_n558, us12_n559, us12_n560, us12_n561, us12_n562, us12_n563, 
       us12_n564, us12_n565, us12_n566, us12_n567, us12_n568, us12_n569, us12_n570, us12_n571, us12_n572, 
       us12_n573, us12_n574, us12_n575, us12_n576, us12_n577, us12_n578, us12_n579, us12_n580, us12_n581, 
       us12_n582, us12_n583, us12_n584, us12_n585, us12_n586, us12_n587, us12_n588, us12_n589, us12_n590, 
       us12_n591, us12_n592, us12_n593, us12_n594, us12_n595, us12_n596, us12_n597, us12_n598, us12_n599, 
       us12_n600, us12_n601, us12_n602, us12_n603, us12_n604, us12_n605, us12_n606, us12_n607, us12_n608, 
       us12_n609, us12_n610, us12_n611, us12_n612, us12_n613, us12_n614, us12_n615, us12_n616, us12_n617, 
       us12_n618, us12_n619, us12_n620, us12_n621, us12_n622, us12_n623, us12_n624, us12_n625, us12_n626, 
       us12_n627, us12_n628, us12_n629, us12_n630, us12_n631, us12_n632, us12_n633, us12_n634, us12_n635, 
       us12_n636, us12_n637, us12_n638, us12_n639, us12_n640, us12_n641, us12_n642, us12_n643, us12_n644, 
       us12_n645, us12_n646, us12_n647, us12_n648, us12_n649, us12_n650, us12_n651, us12_n652, us12_n653, 
       us12_n654, us12_n655, us12_n656, us12_n657, us12_n658, us12_n659, us12_n660, us12_n661, us12_n662, 
       us12_n663, us12_n664, us12_n665, us12_n666, us12_n667, us12_n668, us12_n669, us12_n670, us12_n671, 
       us12_n672, us12_n673, us12_n674, us12_n675, us12_n676, us12_n677, us12_n678, us12_n679, us12_n680, 
       us12_n681, us12_n682, us12_n683, us12_n684, us12_n685, us12_n686, us12_n687, us12_n688, us12_n689, 
       us12_n690, us12_n691, us12_n692, us12_n693, us12_n694, us12_n695, us12_n696, us12_n697, us12_n698, 
       us12_n699, us12_n700, us12_n701, us12_n702, us12_n703, us12_n704, us12_n705, us12_n706, us12_n707, 
       us12_n708, us12_n709, us12_n710, us12_n711, us12_n712, us12_n713, us12_n714, us12_n715, us12_n716, 
       us12_n717, us12_n718, us12_n719, us12_n720, us12_n721, us12_n722, us12_n723, us12_n724, us12_n725, 
       us12_n726, us12_n727, us12_n728, us12_n729, us12_n730, us12_n731, us12_n732, us12_n733, us12_n734, 
       us12_n735, us12_n736, us12_n737, us12_n738, us12_n739, us12_n740, us12_n741, us12_n742, us12_n743, 
       us12_n744, us12_n745, us12_n746, us12_n747, us12_n748, us12_n749, us12_n750, us12_n751, us12_n752, 
       us12_n753, us12_n754, us12_n755, us12_n756, us12_n757, us12_n758, us12_n759, us12_n760, us12_n761, 
       us12_n762, us12_n763, us12_n764, us12_n765, us12_n766, us12_n767, us12_n768, us12_n769, us12_n770, 
       us12_n771, us12_n772, us12_n773, us12_n774, us12_n775, us12_n776, us12_n777, us12_n778, us12_n779, 
       us12_n780, us12_n781, us12_n782, us12_n783, us12_n784, us12_n785, us12_n786, us12_n787, us12_n788, 
       us12_n789, us12_n790, us12_n791, us12_n792, us12_n793, us12_n794, us12_n795, us12_n796, us12_n797, 
       us12_n798, us12_n799, us12_n800, us12_n801, us12_n802, us12_n803, us12_n804, us12_n805, us12_n806, 
       us12_n807, us12_n808, us12_n809, us12_n810, us12_n811, us12_n812, us12_n813, us12_n814, us12_n815, 
       us12_n816, us12_n817, us12_n818, us12_n819, us12_n820, us12_n821, us12_n822, us12_n823, us12_n824, 
       us12_n825, us12_n826, us12_n827, us12_n828, us12_n829, us12_n830, us12_n831, us12_n832, us12_n833, 
       us12_n834, us12_n835, us12_n836, us12_n837, us12_n838, us12_n839, us12_n840, us12_n841, us12_n842, 
       us12_n843, us12_n844, us12_n845, us12_n846, us12_n847, us12_n848, us12_n849, us12_n850, us12_n851, 
       us12_n852, us12_n853, us12_n854, us12_n855, us12_n856, us12_n857, us12_n858, us12_n859, us12_n860, 
       us12_n861, us12_n862, us12_n863, us12_n864, us12_n865, us12_n866, us12_n867, us12_n868, us12_n869, 
       us12_n870, us12_n871, us12_n872, us12_n873, us12_n874, us12_n875, us12_n876, us21_n438, us21_n439, 
       us21_n440, us21_n441, us21_n442, us21_n443, us21_n444, us21_n445, us21_n446, us21_n447, us21_n448, 
       us21_n449, us21_n450, us21_n451, us21_n452, us21_n453, us21_n454, us21_n455, us21_n456, us21_n457, 
       us21_n458, us21_n459, us21_n460, us21_n461, us21_n462, us21_n463, us21_n464, us21_n465, us21_n466, 
       us21_n467, us21_n468, us21_n469, us21_n470, us21_n471, us21_n472, us21_n473, us21_n474, us21_n475, 
       us21_n476, us21_n477, us21_n478, us21_n479, us21_n480, us21_n481, us21_n482, us21_n483, us21_n484, 
       us21_n485, us21_n486, us21_n487, us21_n488, us21_n489, us21_n490, us21_n491, us21_n492, us21_n493, 
       us21_n494, us21_n495, us21_n496, us21_n497, us21_n498, us21_n499, us21_n500, us21_n501, us21_n502, 
       us21_n503, us21_n504, us21_n505, us21_n506, us21_n507, us21_n508, us21_n509, us21_n510, us21_n511, 
       us21_n512, us21_n513, us21_n514, us21_n515, us21_n516, us21_n517, us21_n518, us21_n519, us21_n520, 
       us21_n521, us21_n522, us21_n523, us21_n524, us21_n525, us21_n526, us21_n527, us21_n528, us21_n529, 
       us21_n530, us21_n531, us21_n532, us21_n533, us21_n534, us21_n535, us21_n536, us21_n537, us21_n538, 
       us21_n539, us21_n540, us21_n541, us21_n542, us21_n543, us21_n544, us21_n545, us21_n546, us21_n547, 
       us21_n548, us21_n549, us21_n550, us21_n551, us21_n552, us21_n553, us21_n554, us21_n555, us21_n556, 
       us21_n557, us21_n558, us21_n559, us21_n560, us21_n561, us21_n562, us21_n563, us21_n564, us21_n565, 
       us21_n566, us21_n567, us21_n568, us21_n569, us21_n570, us21_n571, us21_n572, us21_n573, us21_n574, 
       us21_n575, us21_n576, us21_n577, us21_n578, us21_n579, us21_n580, us21_n581, us21_n582, us21_n583, 
       us21_n584, us21_n585, us21_n586, us21_n587, us21_n588, us21_n589, us21_n590, us21_n591, us21_n592, 
       us21_n593, us21_n594, us21_n595, us21_n596, us21_n597, us21_n598, us21_n599, us21_n600, us21_n601, 
       us21_n602, us21_n603, us21_n604, us21_n605, us21_n606, us21_n607, us21_n608, us21_n609, us21_n610, 
       us21_n611, us21_n612, us21_n613, us21_n614, us21_n615, us21_n616, us21_n617, us21_n618, us21_n619, 
       us21_n620, us21_n621, us21_n622, us21_n623, us21_n624, us21_n625, us21_n626, us21_n627, us21_n628, 
       us21_n629, us21_n630, us21_n631, us21_n632, us21_n633, us21_n634, us21_n635, us21_n636, us21_n637, 
       us21_n638, us21_n639, us21_n640, us21_n641, us21_n642, us21_n643, us21_n644, us21_n645, us21_n646, 
       us21_n647, us21_n648, us21_n649, us21_n650, us21_n651, us21_n652, us21_n653, us21_n654, us21_n655, 
       us21_n656, us21_n657, us21_n658, us21_n659, us21_n660, us21_n661, us21_n662, us21_n663, us21_n664, 
       us21_n665, us21_n666, us21_n667, us21_n668, us21_n669, us21_n670, us21_n671, us21_n672, us21_n673, 
       us21_n674, us21_n675, us21_n676, us21_n677, us21_n678, us21_n679, us21_n680, us21_n681, us21_n682, 
       us21_n683, us21_n684, us21_n685, us21_n686, us21_n687, us21_n688, us21_n689, us21_n690, us21_n691, 
       us21_n692, us21_n693, us21_n694, us21_n695, us21_n696, us21_n697, us21_n698, us21_n699, us21_n700, 
       us21_n701, us21_n702, us21_n703, us21_n704, us21_n705, us21_n706, us21_n707, us21_n708, us21_n709, 
       us21_n710, us21_n711, us21_n712, us21_n713, us21_n714, us21_n715, us21_n716, us21_n717, us21_n718, 
       us21_n719, us21_n720, us21_n721, us21_n722, us21_n723, us21_n724, us21_n725, us21_n726, us21_n727, 
       us21_n728, us21_n729, us21_n730, us21_n731, us21_n732, us21_n733, us21_n734, us21_n735, us21_n736, 
       us21_n737, us21_n738, us21_n739, us21_n740, us21_n741, us21_n742, us21_n743, us21_n744, us21_n745, 
       us21_n746, us21_n747, us21_n748, us21_n749, us21_n750, us21_n751, us21_n752, us21_n753, us21_n754, 
       us21_n755, us21_n756, us21_n757, us21_n758, us21_n759, us21_n760, us21_n761, us21_n762, us21_n763, 
       us21_n764, us21_n765, us21_n766, us21_n767, us21_n768, us21_n769, us21_n770, us21_n771, us21_n772, 
       us21_n773, us21_n774, us21_n775, us21_n776, us21_n777, us21_n778, us21_n779, us21_n780, us21_n781, 
       us21_n782, us21_n783, us21_n784, us21_n785, us21_n786, us21_n787, us21_n788, us21_n789, us21_n790, 
       us21_n791, us21_n792, us21_n793, us21_n794, us21_n795, us21_n796, us21_n797, us21_n798, us21_n799, 
       us21_n800, us21_n801, us21_n802, us21_n803, us21_n804, us21_n805, us21_n806, us21_n807, us21_n808, 
       us21_n809, us21_n810, us21_n811, us21_n812, us21_n813, us21_n814, us21_n815, us21_n816, us21_n817, 
       us21_n818, us21_n819, us21_n820, us21_n821, us21_n822, us21_n823, us21_n824, us21_n825, us21_n826, 
       us21_n827, us21_n828, us21_n829, us21_n830, us21_n831, us21_n832, us21_n833, us21_n834, us21_n835, 
       us21_n836, us21_n837, us21_n838, us21_n839, us21_n840, us21_n841, us21_n842, us21_n843, us21_n844, 
       us21_n845, us21_n846, us21_n847, us21_n848, us21_n849, us21_n850, us21_n851, us21_n852, us21_n853, 
       us21_n854, us21_n855, us21_n856, us21_n857, us21_n858, us21_n859, us21_n860, us21_n861, us21_n862, 
       us21_n863, us21_n864, us21_n865, us21_n866, us21_n867, us21_n868, us21_n869, us21_n870, us21_n871, 
       us21_n872, us21_n873,  us21_n874;
  NOR3_X1 us12_U10 (.ZN( us12_n504 ) , .A2( us12_n679 ) , .A3( us12_n777 ) , .A1( us12_n876 ) );
  NOR4_X1 us12_U100 (.A4( us12_n529 ) , .A3( us12_n530 ) , .ZN( us12_n537 ) , .A2( us12_n684 ) , .A1( us12_n794 ) );
  NAND4_X1 us12_U101 (.A4( us12_n479 ) , .A3( us12_n480 ) , .A2( us12_n481 ) , .A1( us12_n482 ) , .ZN( us12_n694 ) );
  NOR3_X1 us12_U102 (.ZN( us12_n480 ) , .A2( us12_n508 ) , .A3( us12_n601 ) , .A1( us12_n610 ) );
  AOI211_X1 us12_U103 (.B( us12_n477 ) , .A( us12_n478 ) , .ZN( us12_n482 ) , .C2( us12_n833 ) , .C1( us12_n861 ) );
  NOR4_X1 us12_U104 (.ZN( us12_n481 ) , .A3( us12_n532 ) , .A4( us12_n545 ) , .A2( us12_n567 ) , .A1( us12_n717 ) );
  NAND4_X1 us12_U105 (.A4( us12_n548 ) , .A3( us12_n549 ) , .A2( us12_n550 ) , .A1( us12_n551 ) , .ZN( us12_n745 ) );
  NOR3_X1 us12_U106 (.ZN( us12_n549 ) , .A2( us12_n651 ) , .A1( us12_n667 ) , .A3( us12_n771 ) );
  AOI211_X1 us12_U107 (.B( us12_n539 ) , .A( us12_n540 ) , .ZN( us12_n551 ) , .C2( us12_n839 ) , .C1( us12_n851 ) );
  NOR4_X1 us12_U108 (.A4( us12_n541 ) , .A3( us12_n542 ) , .A2( us12_n543 ) , .ZN( us12_n550 ) , .A1( us12_n688 ) );
  NOR4_X1 us12_U109 (.ZN( us12_n620 ) , .A1( us12_n656 ) , .A3( us12_n666 ) , .A4( us12_n682 ) , .A2( us12_n766 ) );
  INV_X1 us12_U11 (.A( us12_n706 ) , .ZN( us12_n876 ) );
  NOR4_X1 us12_U110 (.A4( us12_n609 ) , .A3( us12_n610 ) , .A2( us12_n611 ) , .A1( us12_n612 ) , .ZN( us12_n619 ) );
  NOR4_X1 us12_U111 (.A4( us12_n614 ) , .A3( us12_n615 ) , .A2( us12_n616 ) , .A1( us12_n617 ) , .ZN( us12_n618 ) );
  NOR2_X1 us12_U112 (.ZN( us12_n686 ) , .A1( us12_n831 ) , .A2( us12_n832 ) );
  NAND4_X1 us12_U113 (.A4( us12_n485 ) , .A3( us12_n486 ) , .A2( us12_n487 ) , .A1( us12_n488 ) , .ZN( us12_n778 ) );
  NOR4_X1 us12_U114 (.A4( us12_n484 ) , .ZN( us12_n487 ) , .A1( us12_n566 ) , .A2( us12_n581 ) , .A3( us12_n602 ) );
  NOR4_X1 us12_U115 (.ZN( us12_n486 ) , .A1( us12_n507 ) , .A2( us12_n519 ) , .A4( us12_n546 ) , .A3( us12_n611 ) );
  NOR4_X1 us12_U116 (.ZN( us12_n485 ) , .A2( us12_n533 ) , .A1( us12_n558 ) , .A3( us12_n631 ) , .A4( us12_n718 ) );
  NAND4_X1 us12_U117 (.A4( us12_n691 ) , .A3( us12_n692 ) , .A1( us12_n693 ) , .ZN( us12_n776 ) , .A2( us12_n872 ) );
  AOI221_X1 us12_U118 (.A( us12_n681 ) , .ZN( us12_n692 ) , .B2( us12_n840 ) , .C1( us12_n842 ) , .C2( us12_n862 ) , .B1( us12_n865 ) );
  INV_X1 us12_U119 (.A( us12_n679 ) , .ZN( us12_n872 ) );
  NOR3_X1 us12_U12 (.A3( us12_n621 ) , .A2( us12_n622 ) , .ZN( us12_n636 ) , .A1( us12_n725 ) );
  NOR4_X1 us12_U120 (.A4( us12_n687 ) , .A3( us12_n688 ) , .A2( us12_n689 ) , .A1( us12_n690 ) , .ZN( us12_n691 ) );
  NAND4_X1 us12_U121 (.A4( us12_n719 ) , .A3( us12_n720 ) , .A2( us12_n721 ) , .ZN( us12_n741 ) , .A1( us12_n857 ) );
  INV_X1 us12_U122 (.A( us12_n709 ) , .ZN( us12_n857 ) );
  AOI221_X1 us12_U123 (.A( us12_n710 ) , .ZN( us12_n721 ) , .C2( us12_n844 ) , .B2( us12_n845 ) , .C1( us12_n861 ) , .B1( us12_n862 ) );
  NOR4_X1 us12_U124 (.A4( us12_n715 ) , .A3( us12_n716 ) , .A2( us12_n717 ) , .A1( us12_n718 ) , .ZN( us12_n719 ) );
  NAND4_X1 us12_U125 (.A4( us12_n473 ) , .A3( us12_n474 ) , .A2( us12_n475 ) , .A1( us12_n476 ) , .ZN( us12_n678 ) );
  NOR4_X1 us12_U126 (.ZN( us12_n475 ) , .A1( us12_n531 ) , .A3( us12_n568 ) , .A4( us12_n600 ) , .A2( us12_n642 ) );
  NOR4_X1 us12_U127 (.A4( us12_n470 ) , .ZN( us12_n476 ) , .A3( us12_n556 ) , .A1( us12_n735 ) , .A2( us12_n755 ) );
  NOR4_X1 us12_U128 (.ZN( us12_n474 ) , .A1( us12_n506 ) , .A3( us12_n544 ) , .A2( us12_n583 ) , .A4( us12_n716 ) );
  NOR2_X1 us12_U129 (.ZN( us12_n733 ) , .A2( us12_n832 ) , .A1( us12_n845 ) );
  NOR2_X1 us12_U13 (.ZN( us12_n495 ) , .A1( us12_n678 ) , .A2( us12_n694 ) );
  NOR2_X1 us12_U130 (.ZN( us12_n789 ) , .A2( us12_n862 ) , .A1( us12_n868 ) );
  NAND4_X1 us12_U131 (.A4( us12_n573 ) , .A3( us12_n574 ) , .A1( us12_n575 ) , .ZN( us12_n723 ) , .A2( us12_n874 ) );
  NOR4_X1 us12_U132 (.A4( us12_n569 ) , .A3( us12_n570 ) , .A2( us12_n571 ) , .A1( us12_n572 ) , .ZN( us12_n573 ) );
  AOI221_X1 us12_U133 (.A( us12_n564 ) , .C2( us12_n565 ) , .ZN( us12_n574 ) , .B2( us12_n845 ) , .B1( us12_n852 ) , .C1( us12_n853 ) );
  NOR2_X1 us12_U134 (.ZN( us12_n575 ) , .A1( us12_n622 ) , .A2( us12_n745 ) );
  NAND4_X1 us12_U135 (.A4( us12_n633 ) , .A3( us12_n634 ) , .A2( us12_n635 ) , .A1( us12_n636 ) , .ZN( us12_n743 ) );
  AOI211_X1 us12_U136 (.B( us12_n623 ) , .A( us12_n624 ) , .ZN( us12_n635 ) , .C2( us12_n836 ) , .C1( us12_n863 ) );
  NOR4_X1 us12_U137 (.A4( us12_n629 ) , .A3( us12_n630 ) , .A2( us12_n631 ) , .A1( us12_n632 ) , .ZN( us12_n633 ) );
  NOR4_X1 us12_U138 (.A4( us12_n626 ) , .A3( us12_n627 ) , .A2( us12_n628 ) , .ZN( us12_n634 ) , .A1( us12_n664 ) );
  NAND4_X1 us12_U139 (.A4( us12_n493 ) , .A3( us12_n494 ) , .A1( us12_n495 ) , .ZN( us12_n802 ) , .A2( us12_n867 ) );
  NOR2_X1 us12_U14 (.A1( us12_n678 ) , .ZN( us12_n693 ) , .A2( us12_n807 ) );
  AOI221_X1 us12_U140 (.A( us12_n489 ) , .ZN( us12_n494 ) , .B2( us12_n836 ) , .C2( us12_n841 ) , .C1( us12_n851 ) , .B1( us12_n860 ) );
  INV_X1 us12_U141 (.A( us12_n778 ) , .ZN( us12_n867 ) );
  NOR4_X1 us12_U142 (.A2( us12_n491 ) , .A1( us12_n492 ) , .ZN( us12_n493 ) , .A3( us12_n580 ) , .A4( us12_n612 ) );
  NOR4_X1 us12_U143 (.A3( us12_n755 ) , .A2( us12_n756 ) , .A1( us12_n757 ) , .ZN( us12_n758 ) , .A4( us12_n869 ) );
  AOI211_X1 us12_U144 (.B( us12_n745 ) , .A( us12_n746 ) , .ZN( us12_n759 ) , .C1( us12_n832 ) , .C2( us12_n853 ) );
  NOR3_X1 us12_U145 (.A3( us12_n741 ) , .A2( us12_n742 ) , .A1( us12_n743 ) , .ZN( us12_n760 ) );
  NOR2_X1 us12_U146 (.ZN( us12_n647 ) , .A1( us12_n854 ) , .A2( us12_n868 ) );
  INV_X1 us12_U147 (.A( us12_n762 ) , .ZN( us12_n830 ) );
  INV_X1 us12_U148 (.A( us12_n754 ) , .ZN( us12_n869 ) );
  OAI21_X1 us12_U149 (.B1( us12_n753 ) , .ZN( us12_n754 ) , .A( us12_n845 ) , .B2( us12_n868 ) );
  INV_X1 us12_U15 (.A( us12_n607 ) , .ZN( us12_n874 ) );
  OR4_X1 us12_U150 (.ZN( us12_n466 ) , .A4( us12_n518 ) , .A3( us12_n529 ) , .A2( us12_n578 ) , .A1( us12_n712 ) );
  OR4_X1 us12_U151 (.A4( us12_n566 ) , .A3( us12_n567 ) , .A2( us12_n568 ) , .ZN( us12_n572 ) , .A1( us12_n665 ) );
  OR4_X1 us12_U152 (.ZN( us12_n492 ) , .A4( us12_n534 ) , .A2( us12_n547 ) , .A1( us12_n559 ) , .A3( us12_n632 ) );
  OR4_X1 us12_U153 (.A4( us12_n518 ) , .A2( us12_n519 ) , .A1( us12_n520 ) , .ZN( us12_n522 ) , .A3( us12_n821 ) );
  OR4_X1 us12_U154 (.A4( us12_n682 ) , .A3( us12_n683 ) , .A2( us12_n684 ) , .A1( us12_n685 ) , .ZN( us12_n690 ) );
  OR4_X1 us12_U155 (.A4( us12_n580 ) , .A3( us12_n581 ) , .A2( us12_n582 ) , .A1( us12_n583 ) , .ZN( us12_n584 ) );
  NAND2_X1 us12_U156 (.ZN( us12_n613 ) , .A2( us12_n837 ) , .A1( us12_n873 ) );
  OR3_X1 us12_U157 (.A3( us12_n506 ) , .A2( us12_n507 ) , .A1( us12_n508 ) , .ZN( us12_n511 ) );
  INV_X1 us12_U158 (.A( us12_n463 ) , .ZN( us12_n864 ) );
  OAI21_X1 us12_U159 (.ZN( us12_n463 ) , .B1( us12_n809 ) , .A( us12_n834 ) , .B2( us12_n851 ) );
  INV_X1 us12_U16 (.A( us12_n680 ) , .ZN( us12_n840 ) );
  INV_X1 us12_U160 (.A( us12_n672 ) , .ZN( us12_n859 ) );
  AOI21_X1 us12_U161 (.A( us12_n670 ) , .B1( us12_n671 ) , .ZN( us12_n672 ) , .B2( us12_n856 ) );
  OAI222_X1 us12_U162 (.B2( us12_n708 ) , .ZN( us12_n709 ) , .C2( us12_n724 ) , .B1( us12_n747 ) , .A1( us12_n806 ) , .C1( us12_n814 ) , .A2( us12_n815 ) );
  AOI22_X1 us12_U163 (.ZN( us12_n696 ) , .A1( us12_n830 ) , .B2( us12_n843 ) , .A2( us12_n865 ) , .B1( us12_n868 ) );
  INV_X1 us12_U164 (.A( us12_n730 ) , .ZN( us12_n839 ) );
  NAND2_X1 us12_U165 (.A1( us12_n447 ) , .A2( us12_n465 ) , .ZN( us12_n749 ) );
  AOI221_X1 us12_U166 (.A( us12_n483 ) , .ZN( us12_n488 ) , .B1( us12_n831 ) , .C2( us12_n844 ) , .C1( us12_n852 ) , .B2( us12_n862 ) );
  OAI22_X1 us12_U167 (.ZN( us12_n483 ) , .A1( us12_n708 ) , .B2( us12_n785 ) , .A2( us12_n806 ) , .B1( us12_n812 ) );
  INV_X1 us12_U168 (.A( us12_n790 ) , .ZN( us12_n832 ) );
  NAND2_X1 us12_U169 (.A1( us12_n451 ) , .A2( us12_n453 ) , .ZN( us12_n762 ) );
  NOR4_X1 us12_U17 (.A4( us12_n445 ) , .A3( us12_n446 ) , .A2( us12_n516 ) , .A1( us12_n541 ) , .ZN( us12_n706 ) );
  AOI211_X1 us12_U170 (.A( us12_n637 ) , .ZN( us12_n645 ) , .B( us12_n743 ) , .C2( us12_n839 ) , .C1( us12_n854 ) );
  OAI22_X1 us12_U171 (.ZN( us12_n637 ) , .A1( us12_n699 ) , .B2( us12_n728 ) , .A2( us12_n762 ) , .B1( us12_n816 ) );
  INV_X1 us12_U172 (.A( us12_n786 ) , .ZN( us12_n862 ) );
  OAI22_X1 us12_U173 (.B2( us12_n779 ) , .B1( us12_n780 ) , .ZN( us12_n781 ) , .A2( us12_n814 ) , .A1( us12_n815 ) );
  OAI22_X1 us12_U174 (.ZN( us12_n489 ) , .A1( us12_n724 ) , .B2( us12_n728 ) , .B1( us12_n730 ) , .A2( us12_n779 ) );
  INV_X1 us12_U175 (.A( us12_n788 ) , .ZN( us12_n845 ) );
  INV_X1 us12_U176 (.A( us12_n816 ) , .ZN( us12_n831 ) );
  OAI22_X1 us12_U177 (.A1( us12_n724 ) , .ZN( us12_n726 ) , .B2( us12_n750 ) , .B1( us12_n812 ) , .A2( us12_n816 ) );
  OAI22_X1 us12_U178 (.B2( us12_n803 ) , .B1( us12_n804 ) , .A2( us12_n805 ) , .A1( us12_n806 ) , .ZN( us12_n808 ) );
  OAI22_X1 us12_U179 (.ZN( us12_n496 ) , .A2( us12_n744 ) , .A1( us12_n780 ) , .B1( us12_n791 ) , .B2( us12_n806 ) );
  OR3_X1 us12_U18 (.ZN( us12_n446 ) , .A1( us12_n528 ) , .A3( us12_n577 ) , .A2( us12_n875 ) );
  INV_X1 us12_U180 (.A( us12_n814 ) , .ZN( us12_n833 ) );
  INV_X1 us12_U181 (.A( us12_n805 ) , .ZN( us12_n860 ) );
  OAI22_X1 us12_U182 (.ZN( us12_n710 ) , .A2( us12_n728 ) , .B2( us12_n729 ) , .A1( us12_n744 ) , .B1( us12_n813 ) );
  INV_X1 us12_U183 (.A( us12_n750 ) , .ZN( us12_n842 ) );
  OAI22_X1 us12_U184 (.B1( us12_n490 ) , .ZN( us12_n491 ) , .A1( us12_n686 ) , .A2( us12_n763 ) , .B2( us12_n817 ) );
  NOR3_X1 us12_U185 (.ZN( us12_n490 ) , .A1( us12_n782 ) , .A2( us12_n850 ) , .A3( us12_n863 ) );
  OAI22_X1 us12_U186 (.ZN( us12_n695 ) , .A2( us12_n730 ) , .A1( us12_n780 ) , .B1( us12_n791 ) , .B2( us12_n817 ) );
  OAI22_X1 us12_U187 (.B2( us12_n744 ) , .ZN( us12_n746 ) , .A2( us12_n762 ) , .B1( us12_n780 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U188 (.ZN( us12_n532 ) , .A2( us12_n749 ) , .A1( us12_n750 ) );
  INV_X1 us12_U189 (.A( us12_n744 ) , .ZN( us12_n837 ) );
  OR4_X1 us12_U19 (.A4( us12_n442 ) , .A2( us12_n443 ) , .A1( us12_n444 ) , .ZN( us12_n445 ) , .A3( us12_n553 ) );
  NOR2_X1 us12_U190 (.ZN( us12_n666 ) , .A1( us12_n728 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U191 (.ZN( us12_n615 ) , .A1( us12_n785 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U192 (.ZN( us12_n629 ) , .A2( us12_n728 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U193 (.ZN( us12_n715 ) , .A1( us12_n805 ) , .A2( us12_n817 ) );
  NOR2_X1 us12_U194 (.ZN( us12_n570 ) , .A1( us12_n728 ) , .A2( us12_n806 ) );
  NOR2_X1 us12_U195 (.A2( us12_n708 ) , .A1( us12_n750 ) , .ZN( us12_n771 ) );
  NOR2_X1 us12_U196 (.ZN( us12_n611 ) , .A2( us12_n780 ) , .A1( us12_n806 ) );
  NOR2_X1 us12_U197 (.ZN( us12_n601 ) , .A2( us12_n780 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U198 (.ZN( us12_n667 ) , .A1( us12_n750 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U199 (.ZN( us12_n555 ) , .A1( us12_n750 ) , .A2( us12_n791 ) );
  INV_X1 us12_U20 (.A( us12_n613 ) , .ZN( us12_n875 ) );
  NOR2_X1 us12_U200 (.ZN( us12_n654 ) , .A1( us12_n728 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U201 (.ZN( us12_n528 ) , .A2( us12_n724 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U202 (.ZN( us12_n546 ) , .A2( us12_n780 ) , .A1( us12_n814 ) );
  NOR2_X1 us12_U203 (.ZN( us12_n577 ) , .A2( us12_n699 ) , .A1( us12_n814 ) );
  NOR2_X1 us12_U204 (.ZN( us12_n508 ) , .A2( us12_n780 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U205 (.ZN( us12_n543 ) , .A2( us12_n708 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U206 (.ZN( us12_n664 ) , .A1( us12_n785 ) , .A2( us12_n791 ) );
  NOR2_X1 us12_U207 (.A2( us12_n744 ) , .ZN( us12_n755 ) , .A1( us12_n805 ) );
  NOR2_X1 us12_U208 (.ZN( us12_n735 ) , .A2( us12_n803 ) , .A1( us12_n805 ) );
  INV_X1 us12_U209 (.A( us12_n792 ) , .ZN( us12_n851 ) );
  INV_X1 us12_U21 (.A( us12_n749 ) , .ZN( us12_n863 ) );
  INV_X1 us12_U210 (.A( us12_n728 ) , .ZN( us12_n852 ) );
  NOR2_X1 us12_U211 (.A2( us12_n744 ) , .ZN( us12_n769 ) , .A1( us12_n812 ) );
  INV_X1 us12_U212 (.A( us12_n747 ) , .ZN( us12_n834 ) );
  NOR2_X1 us12_U213 (.A1( us12_n699 ) , .ZN( us12_n768 ) , .A2( us12_n813 ) );
  INV_X1 us12_U214 (.A( us12_n806 ) , .ZN( us12_n841 ) );
  NOR2_X1 us12_U215 (.ZN( us12_n531 ) , .A2( us12_n780 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U216 (.ZN( us12_n509 ) , .A1( us12_n729 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U217 (.ZN( us12_n599 ) , .A2( us12_n791 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U218 (.ZN( us12_n661 ) , .A1( us12_n729 ) , .A2( us12_n790 ) );
  NOR2_X1 us12_U219 (.ZN( us12_n507 ) , .A1( us12_n812 ) , .A2( us12_n817 ) );
  AOI222_X1 us12_U22 (.ZN( us12_n605 ) , .B2( us12_n671 ) , .B1( us12_n753 ) , .C2( us12_n831 ) , .A1( us12_n833 ) , .A2( us12_n862 ) , .C1( us12_n863 ) );
  NOR2_X1 us12_U220 (.ZN( us12_n544 ) , .A2( us12_n785 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U221 (.A1( us12_n749 ) , .ZN( us12_n767 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U222 (.ZN( us12_n545 ) , .A1( us12_n749 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U223 (.ZN( us12_n557 ) , .A1( us12_n792 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U224 (.ZN( us12_n556 ) , .A1( us12_n762 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U225 (.ZN( us12_n609 ) , .A2( us12_n724 ) , .A1( us12_n817 ) );
  NOR2_X1 us12_U226 (.ZN( us12_n663 ) , .A1( us12_n729 ) , .A2( us12_n785 ) );
  NOR2_X1 us12_U227 (.ZN( us12_n517 ) , .A1( us12_n708 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U228 (.ZN( us12_n506 ) , .A2( us12_n728 ) , .A1( us12_n762 ) );
  OAI22_X1 us12_U229 (.B1( us12_n440 ) , .ZN( us12_n444 ) , .A2( us12_n728 ) , .A1( us12_n744 ) , .B2( us12_n749 ) );
  AOI222_X1 us12_U23 (.ZN( us12_n563 ) , .B1( us12_n830 ) , .C1( us12_n841 ) , .A2( us12_n843 ) , .A1( us12_n854 ) , .B2( us12_n863 ) , .C2( us12_n873 ) );
  NOR3_X1 us12_U230 (.ZN( us12_n440 ) , .A2( us12_n836 ) , .A3( us12_n837 ) , .A1( us12_n846 ) );
  NOR2_X1 us12_U231 (.ZN( us12_n614 ) , .A1( us12_n762 ) , .A2( us12_n812 ) );
  NOR2_X1 us12_U232 (.ZN( us12_n533 ) , .A2( us12_n724 ) , .A1( us12_n730 ) );
  NOR2_X1 us12_U233 (.ZN( us12_n579 ) , .A2( us12_n708 ) , .A1( us12_n730 ) );
  NOR2_X1 us12_U234 (.ZN( us12_n521 ) , .A1( us12_n790 ) , .A2( us12_n812 ) );
  NOR2_X1 us12_U235 (.ZN( us12_n558 ) , .A1( us12_n708 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U236 (.ZN( us12_n655 ) , .A1( us12_n790 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U237 (.ZN( us12_n670 ) , .A1( us12_n790 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U238 (.ZN( us12_n668 ) , .A2( us12_n708 ) , .A1( us12_n790 ) );
  NOR2_X1 us12_U239 (.ZN( us12_n530 ) , .A2( us12_n744 ) , .A1( us12_n792 ) );
  AOI222_X1 us12_U24 (.ZN( us12_n660 ) , .A2( us12_n839 ) , .B1( us12_n841 ) , .C2( us12_n845 ) , .A1( us12_n860 ) , .C1( us12_n863 ) , .B2( us12_n870 ) );
  NOR2_X1 us12_U240 (.ZN( us12_n631 ) , .A1( us12_n724 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U241 (.ZN( us12_n630 ) , .A1( us12_n747 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U242 (.ZN( us12_n542 ) , .A1( us12_n762 ) , .A2( us12_n791 ) );
  INV_X1 us12_U243 (.A( us12_n763 ) , .ZN( us12_n866 ) );
  AOI21_X1 us12_U244 (.ZN( us12_n515 ) , .A( us12_n729 ) , .B1( us12_n750 ) , .B2( us12_n803 ) );
  NOR2_X1 us12_U245 (.ZN( us12_n718 ) , .A2( us12_n724 ) , .A1( us12_n744 ) );
  NOR2_X1 us12_U246 (.ZN( us12_n516 ) , .A1( us12_n708 ) , .A2( us12_n744 ) );
  INV_X1 us12_U247 (.A( us12_n729 ) , .ZN( us12_n868 ) );
  NOR2_X1 us12_U248 (.ZN( us12_n656 ) , .A1( us12_n747 ) , .A2( us12_n780 ) );
  AOI21_X1 us12_U249 (.ZN( us12_n540 ) , .A( us12_n763 ) , .B2( us12_n779 ) , .B1( us12_n817 ) );
  INV_X1 us12_U25 (.A( us12_n647 ) , .ZN( us12_n870 ) );
  NOR2_X1 us12_U250 (.ZN( us12_n559 ) , .A2( us12_n791 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U251 (.A2( us12_n708 ) , .A1( us12_n762 ) , .ZN( us12_n794 ) );
  NOR2_X1 us12_U252 (.ZN( us12_n642 ) , .A2( us12_n788 ) , .A1( us12_n791 ) );
  NOR2_X1 us12_U253 (.ZN( us12_n683 ) , .A2( us12_n699 ) , .A1( us12_n803 ) );
  AOI21_X1 us12_U254 (.B1( us12_n625 ) , .ZN( us12_n627 ) , .A( us12_n763 ) , .B2( us12_n814 ) );
  AOI21_X1 us12_U255 (.A( us12_n815 ) , .B2( us12_n816 ) , .B1( us12_n817 ) , .ZN( us12_n818 ) );
  AOI21_X1 us12_U256 (.ZN( us12_n650 ) , .A( us12_n779 ) , .B1( us12_n792 ) , .B2( us12_n805 ) );
  AOI21_X1 us12_U257 (.ZN( us12_n499 ) , .B1( us12_n680 ) , .A( us12_n812 ) , .B2( us12_n816 ) );
  NOR2_X1 us12_U258 (.ZN( us12_n520 ) , .A2( us12_n708 ) , .A1( us12_n814 ) );
  AOI21_X1 us12_U259 (.ZN( us12_n569 ) , .B1( us12_n750 ) , .B2( us12_n762 ) , .A( us12_n780 ) );
  NOR4_X1 us12_U26 (.ZN( us12_n473 ) , .A2( us12_n521 ) , .A4( us12_n594 ) , .A1( us12_n609 ) , .A3( us12_n629 ) );
  OAI221_X1 us12_U260 (.A( us12_n727 ) , .C2( us12_n728 ) , .B2( us12_n729 ) , .B1( us12_n730 ) , .ZN( us12_n737 ) , .C1( us12_n817 ) );
  AOI22_X1 us12_U261 (.ZN( us12_n727 ) , .B1( us12_n832 ) , .A2( us12_n838 ) , .A1( us12_n863 ) , .B2( us12_n866 ) );
  AOI21_X1 us12_U262 (.ZN( us12_n589 ) , .B2( us12_n699 ) , .B1( us12_n815 ) , .A( us12_n817 ) );
  NOR2_X1 us12_U263 (.ZN( us12_n519 ) , .A2( us12_n699 ) , .A1( us12_n816 ) );
  AOI21_X1 us12_U264 (.ZN( us12_n539 ) , .B2( us12_n812 ) , .A( us12_n814 ) , .B1( us12_n815 ) );
  AOI21_X1 us12_U265 (.ZN( us12_n640 ) , .B2( us12_n747 ) , .A( us12_n792 ) , .B1( us12_n803 ) );
  AOI21_X1 us12_U266 (.ZN( us12_n514 ) , .A( us12_n779 ) , .B2( us12_n792 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U267 (.B1( us12_n699 ) , .ZN( us12_n700 ) , .A( us12_n732 ) , .B2( us12_n763 ) );
  AOI21_X1 us12_U268 (.ZN( us12_n591 ) , .B2( us12_n763 ) , .A( us12_n785 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U269 (.ZN( us12_n593 ) , .B1( us12_n750 ) , .A( us12_n792 ) , .B2( us12_n813 ) );
  NOR4_X1 us12_U27 (.A4( us12_n544 ) , .A3( us12_n545 ) , .A2( us12_n546 ) , .A1( us12_n547 ) , .ZN( us12_n548 ) );
  NOR2_X1 us12_U270 (.ZN( us12_n547 ) , .A1( us12_n699 ) , .A2( us12_n744 ) );
  INV_X1 us12_U271 (.A( us12_n791 ) , .ZN( us12_n873 ) );
  AOI21_X1 us12_U272 (.ZN( us12_n564 ) , .B1( us12_n724 ) , .A( us12_n779 ) , .B2( us12_n791 ) );
  AOI21_X1 us12_U273 (.ZN( us12_n497 ) , .A( us12_n779 ) , .B2( us12_n791 ) , .B1( us12_n804 ) );
  AOI21_X1 us12_U274 (.ZN( us12_n498 ) , .A( us12_n724 ) , .B2( us12_n762 ) , .B1( us12_n814 ) );
  AOI21_X1 us12_U275 (.ZN( us12_n649 ) , .B1( us12_n729 ) , .B2( us12_n763 ) , .A( us12_n813 ) );
  NOR2_X1 us12_U276 (.ZN( us12_n529 ) , .A1( us12_n708 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U277 (.ZN( us12_n685 ) , .A1( us12_n729 ) , .A2( us12_n816 ) );
  AOI21_X1 us12_U278 (.B1( us12_n686 ) , .ZN( us12_n687 ) , .A( us12_n728 ) , .B2( us12_n761 ) );
  AOI21_X1 us12_U279 (.A( us12_n812 ) , .B2( us12_n813 ) , .B1( us12_n814 ) , .ZN( us12_n819 ) );
  NOR4_X1 us12_U28 (.A4( us12_n532 ) , .A3( us12_n533 ) , .A2( us12_n534 ) , .ZN( us12_n535 ) , .A1( us12_n820 ) );
  AOI21_X1 us12_U280 (.ZN( us12_n450 ) , .B2( us12_n792 ) , .A( us12_n803 ) , .B1( us12_n815 ) );
  NOR2_X1 us12_U281 (.ZN( us12_n568 ) , .A1( us12_n729 ) , .A2( us12_n762 ) );
  NOR2_X1 us12_U282 (.ZN( us12_n682 ) , .A2( us12_n708 ) , .A1( us12_n817 ) );
  AOI21_X1 us12_U283 (.ZN( us12_n641 ) , .B1( us12_n680 ) , .A( us12_n791 ) , .B2( us12_n817 ) );
  INV_X1 us12_U284 (.A( us12_n699 ) , .ZN( us12_n853 ) );
  AOI21_X1 us12_U285 (.ZN( us12_n689 ) , .B2( us12_n749 ) , .B1( us12_n763 ) , .A( us12_n806 ) );
  AOI21_X1 us12_U286 (.ZN( us12_n639 ) , .B2( us12_n749 ) , .A( us12_n788 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U287 (.A( us12_n790 ) , .B2( us12_n791 ) , .B1( us12_n792 ) , .ZN( us12_n793 ) );
  AOI21_X1 us12_U288 (.A( us12_n733 ) , .ZN( us12_n734 ) , .B2( us12_n780 ) , .B1( us12_n792 ) );
  NOR2_X1 us12_U289 (.ZN( us12_n567 ) , .A1( us12_n747 ) , .A2( us12_n805 ) );
  NOR4_X1 us12_U29 (.ZN( us12_n479 ) , .A1( us12_n520 ) , .A4( us12_n557 ) , .A3( us12_n582 ) , .A2( us12_n630 ) );
  NAND2_X1 us12_U290 (.ZN( us12_n753 ) , .A1( us12_n763 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U291 (.A2( us12_n813 ) , .A1( us12_n815 ) , .ZN( us12_n821 ) );
  NOR2_X1 us12_U292 (.ZN( us12_n578 ) , .A1( us12_n708 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U293 (.ZN( us12_n665 ) , .A1( us12_n780 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U294 (.ZN( us12_n711 ) , .A1( us12_n762 ) , .A2( us12_n763 ) );
  NOR2_X1 us12_U295 (.ZN( us12_n583 ) , .A1( us12_n792 ) , .A2( us12_n817 ) );
  AOI21_X1 us12_U296 (.ZN( us12_n442 ) , .A( us12_n699 ) , .B1( us12_n733 ) , .B2( us12_n750 ) );
  NOR2_X1 us12_U297 (.ZN( us12_n534 ) , .A1( us12_n724 ) , .A2( us12_n788 ) );
  NOR2_X1 us12_U298 (.ZN( us12_n582 ) , .A1( us12_n744 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U299 (.ZN( us12_n684 ) , .A1( us12_n791 ) , .A2( us12_n813 ) );
  NAND2_X1 us12_U3 (.A1( us12_n449 ) , .A2( us12_n460 ) , .ZN( us12_n792 ) );
  NOR4_X1 us12_U30 (.ZN( us12_n456 ) , .A2( us12_n517 ) , .A1( us12_n543 ) , .A3( us12_n579 ) , .A4( us12_n615 ) );
  OAI21_X1 us12_U300 (.A( us12_n698 ) , .ZN( us12_n702 ) , .B2( us12_n750 ) , .B1( us12_n804 ) );
  OAI21_X1 us12_U301 (.ZN( us12_n698 ) , .B2( us12_n833 ) , .B1( us12_n838 ) , .A( us12_n860 ) );
  INV_X1 us12_U302 (.A( us12_n815 ) , .ZN( us12_n855 ) );
  INV_X1 us12_U303 (.A( us12_n785 ) , .ZN( us12_n846 ) );
  OAI21_X1 us12_U304 (.A( us12_n731 ) , .B1( us12_n732 ) , .ZN( us12_n736 ) , .B2( us12_n805 ) );
  OAI21_X1 us12_U305 (.ZN( us12_n731 ) , .A( us12_n833 ) , .B2( us12_n852 ) , .B1( us12_n873 ) );
  INV_X1 us12_U306 (.A( us12_n780 ) , .ZN( us12_n850 ) );
  INV_X1 us12_U307 (.A( us12_n813 ) , .ZN( us12_n836 ) );
  OAI221_X1 us12_U308 (.A( us12_n783 ) , .C2( us12_n784 ) , .B2( us12_n785 ) , .B1( us12_n786 ) , .ZN( us12_n796 ) , .C1( us12_n813 ) );
  AOI22_X1 us12_U309 (.A2( us12_n782 ) , .ZN( us12_n783 ) , .B2( us12_n831 ) , .A1( us12_n834 ) , .B1( us12_n863 ) );
  AOI221_X1 us12_U31 (.A( us12_n713 ) , .B2( us12_n714 ) , .ZN( us12_n720 ) , .C1( us12_n832 ) , .B1( us12_n839 ) , .C2( us12_n863 ) );
  OAI21_X1 us12_U310 (.A( us12_n787 ) , .B2( us12_n788 ) , .B1( us12_n789 ) , .ZN( us12_n795 ) );
  OAI21_X1 us12_U311 (.ZN( us12_n787 ) , .A( us12_n839 ) , .B1( us12_n863 ) , .B2( us12_n873 ) );
  NAND2_X1 us12_U312 (.A2( us12_n762 ) , .A1( us12_n806 ) , .ZN( us12_n810 ) );
  NOR2_X1 us12_U313 (.ZN( us12_n470 ) , .A2( us12_n779 ) , .A1( us12_n815 ) );
  NOR2_X1 us12_U314 (.ZN( us12_n484 ) , .A1( us12_n788 ) , .A2( us12_n805 ) );
  NAND2_X1 us12_U315 (.ZN( us12_n714 ) , .A1( us12_n728 ) , .A2( us12_n780 ) );
  NAND2_X1 us12_U316 (.ZN( us12_n671 ) , .A1( us12_n806 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U317 (.ZN( us12_n526 ) , .A1( us12_n724 ) , .A2( us12_n750 ) );
  AOI21_X1 us12_U318 (.ZN( us12_n443 ) , .B1( us12_n789 ) , .B2( us12_n791 ) , .A( us12_n814 ) );
  INV_X1 us12_U319 (.A( us12_n817 ) , .ZN( us12_n844 ) );
  OR2_X1 us12_U32 (.A2( us12_n711 ) , .A1( us12_n712 ) , .ZN( us12_n713 ) );
  NOR2_X1 us12_U320 (.ZN( us12_n712 ) , .A2( us12_n724 ) , .A1( us12_n790 ) );
  NAND2_X1 us12_U321 (.A1( us12_n699 ) , .A2( us12_n729 ) , .ZN( us12_n782 ) );
  NOR2_X1 us12_U322 (.ZN( us12_n518 ) , .A1( us12_n708 ) , .A2( us12_n788 ) );
  OAI22_X1 us12_U323 (.B2( us12_n750 ) , .B1( us12_n751 ) , .A1( us12_n752 ) , .ZN( us12_n756 ) , .A2( us12_n806 ) );
  NOR3_X1 us12_U324 (.ZN( us12_n752 ) , .A2( us12_n853 ) , .A1( us12_n863 ) , .A3( us12_n865 ) );
  NOR2_X1 us12_U325 (.ZN( us12_n751 ) , .A2( us12_n852 ) , .A1( us12_n860 ) );
  INV_X1 us12_U326 (.A( us12_n724 ) , .ZN( us12_n856 ) );
  NAND2_X2 us12_U327 (.A2( us12_n454 ) , .A1( us12_n472 ) , .ZN( us12_n779 ) );
  AND2_X1 us12_U328 (.ZN( us12_n732 ) , .A1( us12_n779 ) , .A2( us12_n785 ) );
  AOI221_X1 us12_U329 (.A( us12_n764 ) , .ZN( us12_n774 ) , .C2( us12_n810 ) , .B2( us12_n835 ) , .C1( us12_n855 ) , .B1( us12_n866 ) );
  NOR2_X1 us12_U33 (.ZN( us12_n680 ) , .A2( us12_n834 ) , .A1( us12_n839 ) );
  AOI21_X1 us12_U330 (.B2( us12_n763 ) , .ZN( us12_n764 ) , .A( us12_n788 ) , .B1( us12_n792 ) );
  INV_X1 us12_U331 (.A( us12_n761 ) , .ZN( us12_n835 ) );
  NAND2_X1 us12_U332 (.A2( us12_n448 ) , .A1( us12_n460 ) , .ZN( us12_n728 ) );
  NAND2_X1 us12_U333 (.A1( us12_n451 ) , .A2( us12_n454 ) , .ZN( us12_n814 ) );
  NAND2_X1 us12_U334 (.A1( us12_n447 ) , .A2( us12_n449 ) , .ZN( us12_n805 ) );
  NAND2_X1 us12_U335 (.A1( us12_n451 ) , .A2( us12_n471 ) , .ZN( us12_n816 ) );
  NAND2_X1 us12_U336 (.A2( us12_n453 ) , .A1( us12_n455 ) , .ZN( us12_n806 ) );
  NAND2_X1 us12_U337 (.A2( us12_n464 ) , .A1( us12_n465 ) , .ZN( us12_n812 ) );
  NAND2_X1 us12_U338 (.A1( us12_n441 ) , .A2( us12_n460 ) , .ZN( us12_n699 ) );
  NAND2_X1 us12_U339 (.A2( us12_n449 ) , .A1( us12_n452 ) , .ZN( us12_n763 ) );
  AOI222_X1 us12_U34 (.ZN( us12_n469 ) , .B1( us12_n832 ) , .A1( us12_n839 ) , .C1( us12_n842 ) , .C2( us12_n851 ) , .A2( us12_n855 ) , .B2( us12_n865 ) );
  NAND2_X2 us12_U340 (.A1( us12_n455 ) , .A2( us12_n462 ) , .ZN( us12_n750 ) );
  NAND2_X1 us12_U341 (.A2( us12_n448 ) , .A1( us12_n452 ) , .ZN( us12_n729 ) );
  NOR2_X1 us12_U342 (.ZN( us12_n453 ) , .A1( us12_n826 ) , .A2( us12_n827 ) );
  NOR2_X1 us12_U343 (.ZN( us12_n465 ) , .A2( us12_n847 ) , .A1( us12_n848 ) );
  NOR2_X1 us12_U344 (.ZN( us12_n451 ) , .A1( us12_n828 ) , .A2( us12_n829 ) );
  NAND2_X1 us12_U345 (.A1( us12_n462 ) , .A2( us12_n472 ) , .ZN( us12_n788 ) );
  NAND2_X1 us12_U346 (.A2( us12_n461 ) , .A1( us12_n471 ) , .ZN( us12_n697 ) );
  NAND2_X1 us12_U347 (.A2( us12_n461 ) , .A1( us12_n462 ) , .ZN( us12_n747 ) );
  NAND2_X1 us12_U348 (.A1( us12_n451 ) , .A2( us12_n462 ) , .ZN( us12_n790 ) );
  NAND2_X1 us12_U349 (.A1( us12_n452 ) , .A2( us12_n465 ) , .ZN( us12_n669 ) );
  NOR4_X1 us12_U35 (.A1( us12_n466 ) , .ZN( us12_n467 ) , .A4( us12_n542 ) , .A2( us12_n554 ) , .A3( us12_n614 ) );
  NAND2_X1 us12_U350 (.A2( us12_n441 ) , .A1( us12_n447 ) , .ZN( us12_n784 ) );
  NAND2_X2 us12_U351 (.A1( us12_n441 ) , .A2( us12_n464 ) , .ZN( us12_n708 ) );
  NAND2_X1 us12_U352 (.A2( us12_n471 ) , .A1( us12_n472 ) , .ZN( us12_n817 ) );
  NAND2_X1 us12_U353 (.A2( us12_n454 ) , .A1( us12_n455 ) , .ZN( us12_n730 ) );
  NOR2_X1 us12_U354 (.ZN( us12_n447 ) , .A2( us12_n849 ) , .A1( us12_n858 ) );
  NAND2_X1 us12_U355 (.A1( us12_n447 ) , .A2( us12_n448 ) , .ZN( us12_n786 ) );
  NAND2_X1 us12_U356 (.A1( us12_n454 ) , .A2( us12_n461 ) , .ZN( us12_n813 ) );
  NAND2_X2 us12_U357 (.A1( us12_n453 ) , .A2( us12_n472 ) , .ZN( us12_n785 ) );
  NAND2_X1 us12_U358 (.A1( us12_n453 ) , .A2( us12_n461 ) , .ZN( us12_n744 ) );
  NOR2_X1 us12_U359 (.A2( sa12_6 ) , .A1( sa12_7 ) , .ZN( us12_n464 ) );
  AOI221_X1 us12_U36 (.ZN( us12_n468 ) , .C2( us12_n714 ) , .B2( us12_n831 ) , .C1( us12_n845 ) , .B1( us12_n860 ) , .A( us12_n864 ) );
  NOR2_X1 us12_U360 (.A2( sa12_2 ) , .ZN( us12_n461 ) , .A1( us12_n829 ) );
  NOR2_X1 us12_U361 (.A2( sa12_7 ) , .ZN( us12_n460 ) , .A1( us12_n849 ) );
  NOR2_X1 us12_U362 (.A2( sa12_4 ) , .ZN( us12_n449 ) , .A1( us12_n848 ) );
  NOR2_X1 us12_U363 (.A2( sa12_4 ) , .A1( sa12_5 ) , .ZN( us12_n441 ) );
  NOR2_X1 us12_U364 (.A2( sa12_5 ) , .ZN( us12_n448 ) , .A1( us12_n847 ) );
  NOR2_X1 us12_U365 (.A2( sa12_0 ) , .ZN( us12_n454 ) , .A1( us12_n827 ) );
  NOR2_X1 us12_U366 (.A2( sa12_1 ) , .ZN( us12_n471 ) , .A1( us12_n826 ) );
  NOR2_X1 us12_U367 (.A2( sa12_6 ) , .ZN( us12_n452 ) , .A1( us12_n858 ) );
  NOR2_X1 us12_U368 (.A2( sa12_0 ) , .A1( sa12_1 ) , .ZN( us12_n462 ) );
  INV_X1 us12_U369 (.A( sa12_6 ) , .ZN( us12_n849 ) );
  NOR4_X1 us12_U37 (.A4( us12_n577 ) , .A3( us12_n578 ) , .A2( us12_n579 ) , .ZN( us12_n586 ) , .A1( us12_n683 ) );
  INV_X1 us12_U370 (.A( sa12_4 ) , .ZN( us12_n847 ) );
  INV_X1 us12_U371 (.A( sa12_1 ) , .ZN( us12_n827 ) );
  NAND2_X2 us12_U372 (.A1( us12_n455 ) , .A2( us12_n471 ) , .ZN( us12_n803 ) );
  INV_X1 us12_U373 (.A( sa12_0 ) , .ZN( us12_n826 ) );
  INV_X1 us12_U374 (.A( sa12_7 ) , .ZN( us12_n858 ) );
  INV_X1 us12_U375 (.A( sa12_5 ) , .ZN( us12_n848 ) );
  INV_X1 us12_U376 (.A( sa12_2 ) , .ZN( us12_n828 ) );
  AOI21_X1 us12_U377 (.ZN( us12_n510 ) , .B2( us12_n669 ) , .A( us12_n730 ) , .B1( us12_n815 ) );
  OAI22_X1 us12_U378 (.ZN( us12_n624 ) , .B1( us12_n669 ) , .B2( us12_n747 ) , .A1( us12_n815 ) , .A2( us12_n816 ) );
  AOI21_X1 us12_U379 (.ZN( us12_n626 ) , .B2( us12_n669 ) , .A( us12_n790 ) , .B1( us12_n791 ) );
  NOR4_X1 us12_U38 (.A1( us12_n584 ) , .ZN( us12_n585 ) , .A3( us12_n652 ) , .A2( us12_n662 ) , .A4( us12_n767 ) );
  INV_X1 us12_U380 (.A( us12_n669 ) , .ZN( us12_n865 ) );
  NOR2_X1 us12_U381 (.A1( us12_n669 ) , .ZN( us12_n766 ) , .A2( us12_n813 ) );
  AOI21_X1 us12_U382 (.ZN( us12_n477 ) , .A( us12_n669 ) , .B1( us12_n750 ) , .B2( us12_n806 ) );
  NOR2_X1 us12_U383 (.A1( us12_n669 ) , .ZN( us12_n673 ) , .A2( us12_n744 ) );
  NOR2_X1 us12_U384 (.ZN( us12_n602 ) , .A1( us12_n669 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U385 (.A1( us12_n669 ) , .ZN( us12_n688 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U386 (.ZN( us12_n527 ) , .A1( us12_n669 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U387 (.ZN( us12_n652 ) , .A1( us12_n669 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U388 (.ZN( us12_n628 ) , .A2( us12_n669 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U389 (.ZN( us12_n581 ) , .A1( us12_n669 ) , .A2( us12_n788 ) );
  NOR4_X1 us12_U39 (.A4( us12_n661 ) , .A3( us12_n662 ) , .A2( us12_n663 ) , .A1( us12_n664 ) , .ZN( us12_n677 ) );
  OAI22_X1 us12_U390 (.ZN( us12_n590 ) , .B1( us12_n730 ) , .B2( us12_n749 ) , .A2( us12_n786 ) , .A1( us12_n803 ) );
  NAND2_X1 us12_U391 (.A2( us12_n749 ) , .A1( us12_n786 ) , .ZN( us12_n809 ) );
  NOR2_X1 us12_U392 (.ZN( us12_n612 ) , .A1( us12_n779 ) , .A2( us12_n786 ) );
  NOR2_X1 us12_U393 (.ZN( us12_n717 ) , .A2( us12_n744 ) , .A1( us12_n786 ) );
  NOR2_X1 us12_U394 (.ZN( us12_n653 ) , .A1( us12_n762 ) , .A2( us12_n786 ) );
  NOR2_X1 us12_U395 (.ZN( us12_n554 ) , .A1( us12_n786 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U396 (.ZN( us12_n701 ) , .A2( us12_n786 ) , .A1( us12_n817 ) );
  OAI222_X1 us12_U397 (.ZN( us12_n617 ) , .B1( us12_n697 ) , .C1( us12_n724 ) , .C2( us12_n747 ) , .B2( us12_n786 ) , .A2( us12_n792 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U398 (.A1( us12_n730 ) , .ZN( us12_n765 ) , .A2( us12_n786 ) );
  NAND2_X1 us12_U399 (.A1( us12_n729 ) , .A2( us12_n784 ) , .ZN( us12_n811 ) );
  NAND2_X1 us12_U4 (.A1( us12_n449 ) , .A2( us12_n464 ) , .ZN( us12_n724 ) );
  NOR4_X1 us12_U40 (.A4( us12_n665 ) , .A3( us12_n666 ) , .A2( us12_n667 ) , .A1( us12_n668 ) , .ZN( us12_n676 ) );
  OAI22_X1 us12_U400 (.ZN( us12_n588 ) , .A2( us12_n747 ) , .B2( us12_n762 ) , .A1( us12_n763 ) , .B1( us12_n784 ) );
  OAI221_X1 us12_U401 (.A( us12_n696 ) , .ZN( us12_n703 ) , .C2( us12_n784 ) , .C1( us12_n785 ) , .B1( us12_n786 ) , .B2( us12_n806 ) );
  AOI21_X1 us12_U402 (.ZN( us12_n592 ) , .B1( us12_n728 ) , .B2( us12_n784 ) , .A( us12_n790 ) );
  AOI21_X1 us12_U403 (.ZN( us12_n648 ) , .A( us12_n762 ) , .B2( us12_n784 ) , .B1( us12_n792 ) );
  AOI21_X1 us12_U404 (.ZN( us12_n623 ) , .B1( us12_n699 ) , .A( us12_n779 ) , .B2( us12_n784 ) );
  OAI22_X1 us12_U405 (.ZN( us12_n681 ) , .A1( us12_n699 ) , .A2( us12_n730 ) , .B2( us12_n784 ) , .B1( us12_n817 ) );
  OAI21_X1 us12_U406 (.A( us12_n613 ) , .ZN( us12_n616 ) , .B1( us12_n625 ) , .B2( us12_n784 ) );
  NOR2_X1 us12_U407 (.ZN( us12_n610 ) , .A1( us12_n784 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U408 (.ZN( us12_n651 ) , .A1( us12_n784 ) , .A2( us12_n788 ) );
  OAI222_X1 us12_U409 (.A2( us12_n669 ) , .ZN( us12_n674 ) , .B1( us12_n747 ) , .B2( us12_n784 ) , .C2( us12_n788 ) , .C1( us12_n815 ) , .A1( us12_n817 ) );
  NOR4_X1 us12_U41 (.A3( us12_n673 ) , .A1( us12_n674 ) , .ZN( us12_n675 ) , .A4( us12_n715 ) , .A2( us12_n859 ) );
  NOR2_X1 us12_U410 (.ZN( us12_n553 ) , .A2( us12_n744 ) , .A1( us12_n784 ) );
  INV_X1 us12_U411 (.A( us12_n784 ) , .ZN( us12_n861 ) );
  AOI21_X1 us12_U412 (.ZN( us12_n500 ) , .A( us12_n697 ) , .B1( us12_n708 ) , .B2( us12_n786 ) );
  INV_X1 us12_U413 (.A( us12_n697 ) , .ZN( us12_n838 ) );
  NOR2_X1 us12_U414 (.A1( us12_n697 ) , .ZN( us12_n770 ) , .A2( us12_n815 ) );
  AOI21_X1 us12_U415 (.ZN( us12_n571 ) , .B2( us12_n697 ) , .B1( us12_n806 ) , .A( us12_n812 ) );
  NOR2_X1 us12_U416 (.ZN( us12_n632 ) , .A2( us12_n697 ) , .A1( us12_n724 ) );
  AOI21_X1 us12_U417 (.ZN( us12_n478 ) , .B2( us12_n697 ) , .A( us12_n749 ) , .B1( us12_n779 ) );
  NOR2_X1 us12_U418 (.A2( us12_n697 ) , .A1( us12_n780 ) , .ZN( us12_n820 ) );
  NOR2_X1 us12_U419 (.ZN( us12_n662 ) , .A2( us12_n697 ) , .A1( us12_n729 ) );
  AOI221_X1 us12_U42 (.A( us12_n781 ) , .ZN( us12_n798 ) , .C2( us12_n837 ) , .B2( us12_n838 ) , .B1( us12_n865 ) , .C1( us12_n866 ) );
  NOR2_X1 us12_U420 (.ZN( us12_n566 ) , .A2( us12_n697 ) , .A1( us12_n763 ) );
  NOR2_X1 us12_U421 (.ZN( us12_n600 ) , .A2( us12_n697 ) , .A1( us12_n784 ) );
  NOR2_X1 us12_U422 (.A2( us12_n697 ) , .ZN( us12_n716 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U423 (.ZN( us12_n594 ) , .A2( us12_n697 ) , .A1( us12_n728 ) );
  AOI21_X1 us12_U424 (.ZN( us12_n552 ) , .B1( us12_n669 ) , .A( us12_n697 ) , .B2( us12_n805 ) );
  NOR2_X1 us12_U425 (.ZN( us12_n541 ) , .A2( us12_n697 ) , .A1( us12_n699 ) );
  NOR2_X1 us12_U426 (.ZN( us12_n580 ) , .A2( us12_n697 ) , .A1( us12_n791 ) );
  NOR2_X1 us12_U427 (.A2( sa12_2 ) , .A1( sa12_3 ) , .ZN( us12_n472 ) );
  NOR2_X1 us12_U428 (.A2( sa12_3 ) , .ZN( us12_n455 ) , .A1( us12_n828 ) );
  INV_X1 us12_U429 (.A( sa12_3 ) , .ZN( us12_n829 ) );
  NOR4_X1 us12_U43 (.A4( us12_n793 ) , .A3( us12_n794 ) , .A2( us12_n795 ) , .A1( us12_n796 ) , .ZN( us12_n797 ) );
  OAI222_X1 us12_U430 (.ZN( us12_n505 ) , .C2( us12_n625 ) , .B2( us12_n647 ) , .B1( us12_n747 ) , .A2( us12_n748 ) , .C1( us12_n805 ) , .A1( us12_n806 ) );
  OAI222_X1 us12_U431 (.B2( us12_n747 ) , .B1( us12_n748 ) , .A2( us12_n749 ) , .ZN( us12_n757 ) , .C2( us12_n805 ) , .C1( us12_n814 ) , .A1( us12_n817 ) );
  NOR2_X1 us12_U432 (.ZN( us12_n748 ) , .A1( us12_n861 ) , .A2( us12_n862 ) );
  AND2_X1 us12_U433 (.ZN( us12_n438 ) , .A2( us12_n831 ) , .A1( us12_n854 ) );
  AND2_X1 us12_U434 (.ZN( us12_n439 ) , .A2( us12_n843 ) , .A1( us12_n861 ) );
  NOR3_X1 us12_U435 (.A1( us12_n438 ) , .A2( us12_n439 ) , .A3( us12_n576 ) , .ZN( us12_n587 ) );
  INV_X1 us12_U436 (.A( us12_n812 ) , .ZN( us12_n854 ) );
  NAND3_X1 us12_U437 (.ZN( sa11_sr_6 ) , .A3( us12_n797 ) , .A2( us12_n798 ) , .A1( us12_n799 ) );
  NAND3_X1 us12_U438 (.ZN( sa11_sr_5 ) , .A3( us12_n758 ) , .A2( us12_n759 ) , .A1( us12_n760 ) );
  NAND3_X1 us12_U439 (.ZN( sa11_sr_4 ) , .A3( us12_n738 ) , .A2( us12_n739 ) , .A1( us12_n740 ) );
  NOR4_X1 us12_U44 (.A4( us12_n776 ) , .A3( us12_n777 ) , .A1( us12_n778 ) , .ZN( us12_n799 ) , .A2( us12_n801 ) );
  NAND3_X1 us12_U440 (.A3( us12_n675 ) , .A2( us12_n676 ) , .A1( us12_n677 ) , .ZN( us12_n807 ) );
  NAND3_X1 us12_U441 (.ZN( us12_n638 ) , .A3( us12_n708 ) , .A2( us12_n724 ) , .A1( us12_n792 ) );
  NAND3_X1 us12_U442 (.A3( us12_n618 ) , .A2( us12_n619 ) , .A1( us12_n620 ) , .ZN( us12_n725 ) );
  NAND3_X1 us12_U443 (.A3( us12_n585 ) , .A2( us12_n586 ) , .A1( us12_n587 ) , .ZN( us12_n621 ) );
  NAND3_X1 us12_U444 (.ZN( us12_n565 ) , .A3( us12_n680 ) , .A2( us12_n750 ) , .A1( us12_n785 ) );
  NAND3_X1 us12_U445 (.A3( us12_n523 ) , .A2( us12_n524 ) , .A1( us12_n525 ) , .ZN( us12_n742 ) );
  NAND3_X1 us12_U446 (.A3( us12_n512 ) , .A1( us12_n513 ) , .ZN( us12_n608 ) , .A2( us12_n871 ) );
  NAND3_X1 us12_U447 (.A3( us12_n467 ) , .A2( us12_n468 ) , .A1( us12_n469 ) , .ZN( us12_n777 ) );
  INV_X1 us12_U448 (.A( us12_n803 ) , .ZN( us12_n843 ) );
  AOI21_X1 us12_U449 (.ZN( us12_n576 ) , .B2( us12_n724 ) , .B1( us12_n748 ) , .A( us12_n785 ) );
  NOR4_X1 us12_U45 (.A4( us12_n734 ) , .A3( us12_n735 ) , .A2( us12_n736 ) , .A1( us12_n737 ) , .ZN( us12_n738 ) );
  AOI211_X1 us12_U46 (.B( us12_n725 ) , .A( us12_n726 ) , .ZN( us12_n739 ) , .C1( us12_n843 ) , .C2( us12_n855 ) );
  NOR3_X1 us12_U47 (.A3( us12_n722 ) , .A1( us12_n723 ) , .ZN( us12_n740 ) , .A2( us12_n741 ) );
  NAND4_X1 us12_U48 (.ZN( sa11_sr_3 ) , .A4( us12_n704 ) , .A3( us12_n705 ) , .A2( us12_n706 ) , .A1( us12_n707 ) );
  NOR4_X1 us12_U49 (.A4( us12_n700 ) , .A3( us12_n701 ) , .A2( us12_n702 ) , .A1( us12_n703 ) , .ZN( us12_n704 ) );
  NAND2_X1 us12_U5 (.A2( us12_n448 ) , .A1( us12_n464 ) , .ZN( us12_n815 ) );
  AOI211_X1 us12_U50 (.B( us12_n694 ) , .A( us12_n695 ) , .ZN( us12_n705 ) , .C2( us12_n831 ) , .C1( us12_n851 ) );
  NOR2_X1 us12_U51 (.ZN( us12_n707 ) , .A2( us12_n776 ) , .A1( us12_n800 ) );
  NOR2_X1 us12_U52 (.ZN( us12_n804 ) , .A1( us12_n854 ) , .A2( us12_n861 ) );
  NAND4_X1 us12_U53 (.ZN( sa11_sr_0 ) , .A4( us12_n501 ) , .A3( us12_n502 ) , .A2( us12_n503 ) , .A1( us12_n504 ) );
  AOI221_X1 us12_U54 (.A( us12_n497 ) , .ZN( us12_n502 ) , .B2( us12_n843 ) , .C1( us12_n846 ) , .C2( us12_n860 ) , .B1( us12_n862 ) );
  NOR4_X1 us12_U55 (.A4( us12_n498 ) , .A3( us12_n499 ) , .A2( us12_n500 ) , .ZN( us12_n501 ) , .A1( us12_n527 ) );
  AOI211_X1 us12_U56 (.A( us12_n496 ) , .ZN( us12_n503 ) , .B( us12_n802 ) , .C2( us12_n839 ) , .C1( us12_n851 ) );
  NAND4_X1 us12_U57 (.ZN( sa11_sr_1 ) , .A4( us12_n595 ) , .A3( us12_n596 ) , .A2( us12_n597 ) , .A1( us12_n598 ) );
  AOI211_X1 us12_U58 (.B( us12_n589 ) , .A( us12_n590 ) , .ZN( us12_n596 ) , .C2( us12_n811 ) , .C1( us12_n833 ) );
  NOR4_X1 us12_U59 (.A4( us12_n591 ) , .A3( us12_n592 ) , .A2( us12_n593 ) , .A1( us12_n594 ) , .ZN( us12_n595 ) );
  NAND2_X1 us12_U6 (.A2( us12_n441 ) , .A1( us12_n452 ) , .ZN( us12_n791 ) );
  AOI211_X1 us12_U60 (.A( us12_n588 ) , .ZN( us12_n597 ) , .B( us12_n621 ) , .C1( us12_n845 ) , .C2( us12_n855 ) );
  NAND4_X1 us12_U61 (.ZN( sa11_sr_7 ) , .A4( us12_n822 ) , .A3( us12_n823 ) , .A2( us12_n824 ) , .A1( us12_n825 ) );
  NOR4_X1 us12_U62 (.A4( us12_n818 ) , .A3( us12_n819 ) , .A2( us12_n820 ) , .A1( us12_n821 ) , .ZN( us12_n822 ) );
  AOI222_X1 us12_U63 (.C2( us12_n809 ) , .B2( us12_n810 ) , .A2( us12_n811 ) , .ZN( us12_n823 ) , .C1( us12_n832 ) , .A1( us12_n839 ) , .B1( us12_n853 ) );
  AOI211_X1 us12_U64 (.B( us12_n807 ) , .A( us12_n808 ) , .ZN( us12_n824 ) , .C1( us12_n842 ) , .C2( us12_n850 ) );
  NAND4_X1 us12_U65 (.ZN( sa11_sr_2 ) , .A4( us12_n643 ) , .A3( us12_n644 ) , .A2( us12_n645 ) , .A1( us12_n646 ) );
  AOI222_X1 us12_U66 (.B2( us12_n638 ) , .ZN( us12_n644 ) , .B1( us12_n841 ) , .A1( us12_n842 ) , .C2( us12_n846 ) , .C1( us12_n863 ) , .A2( us12_n865 ) );
  NOR4_X1 us12_U67 (.A4( us12_n639 ) , .A3( us12_n640 ) , .A2( us12_n641 ) , .A1( us12_n642 ) , .ZN( us12_n643 ) );
  NOR3_X1 us12_U68 (.A2( us12_n607 ) , .A1( us12_n608 ) , .ZN( us12_n646 ) , .A3( us12_n722 ) );
  NAND4_X1 us12_U69 (.A4( us12_n603 ) , .A3( us12_n604 ) , .A2( us12_n605 ) , .A1( us12_n606 ) , .ZN( us12_n722 ) );
  NAND2_X1 us12_U7 (.A2( us12_n460 ) , .A1( us12_n465 ) , .ZN( us12_n780 ) );
  NOR3_X1 us12_U70 (.A1( us12_n599 ) , .ZN( us12_n604 ) , .A3( us12_n663 ) , .A2( us12_n770 ) );
  NOR4_X1 us12_U71 (.A3( us12_n600 ) , .A2( us12_n601 ) , .A1( us12_n602 ) , .ZN( us12_n603 ) , .A4( us12_n655 ) );
  AOI222_X1 us12_U72 (.ZN( us12_n606 ) , .A1( us12_n830 ) , .C2( us12_n837 ) , .B1( us12_n842 ) , .A2( us12_n856 ) , .B2( us12_n861 ) , .C1( us12_n868 ) );
  NOR4_X1 us12_U73 (.A4( us12_n514 ) , .A3( us12_n515 ) , .A2( us12_n516 ) , .A1( us12_n517 ) , .ZN( us12_n524 ) );
  AOI222_X1 us12_U74 (.ZN( us12_n525 ) , .A1( us12_n834 ) , .B2( us12_n837 ) , .C1( us12_n844 ) , .C2( us12_n850 ) , .A2( us12_n852 ) , .B1( us12_n866 ) );
  NOR4_X1 us12_U75 (.A3( us12_n521 ) , .A1( us12_n522 ) , .ZN( us12_n523 ) , .A2( us12_n673 ) , .A4( us12_n769 ) );
  NAND4_X1 us12_U76 (.A4( us12_n657 ) , .A3( us12_n658 ) , .A2( us12_n659 ) , .A1( us12_n660 ) , .ZN( us12_n800 ) );
  NOR3_X1 us12_U77 (.A3( us12_n648 ) , .A2( us12_n649 ) , .A1( us12_n650 ) , .ZN( us12_n659 ) );
  NOR3_X1 us12_U78 (.A3( us12_n651 ) , .A2( us12_n652 ) , .A1( us12_n653 ) , .ZN( us12_n658 ) );
  NOR3_X1 us12_U79 (.A3( us12_n654 ) , .A2( us12_n655 ) , .A1( us12_n656 ) , .ZN( us12_n657 ) );
  NOR3_X1 us12_U8 (.ZN( us12_n598 ) , .A1( us12_n608 ) , .A3( us12_n723 ) , .A2( us12_n742 ) );
  NAND4_X1 us12_U80 (.A4( us12_n560 ) , .A3( us12_n561 ) , .A2( us12_n562 ) , .A1( us12_n563 ) , .ZN( us12_n607 ) );
  NOR4_X1 us12_U81 (.A4( us12_n552 ) , .A3( us12_n553 ) , .A2( us12_n554 ) , .A1( us12_n555 ) , .ZN( us12_n562 ) );
  NOR4_X1 us12_U82 (.ZN( us12_n561 ) , .A1( us12_n653 ) , .A3( us12_n661 ) , .A4( us12_n685 ) , .A2( us12_n768 ) );
  NOR4_X1 us12_U83 (.A4( us12_n556 ) , .A3( us12_n557 ) , .A2( us12_n558 ) , .A1( us12_n559 ) , .ZN( us12_n560 ) );
  NAND4_X1 us12_U84 (.A4( us12_n772 ) , .A3( us12_n773 ) , .A2( us12_n774 ) , .A1( us12_n775 ) , .ZN( us12_n801 ) );
  NOR3_X1 us12_U85 (.A3( us12_n765 ) , .A2( us12_n766 ) , .A1( us12_n767 ) , .ZN( us12_n773 ) );
  NOR4_X1 us12_U86 (.A4( us12_n768 ) , .A3( us12_n769 ) , .A2( us12_n770 ) , .A1( us12_n771 ) , .ZN( us12_n772 ) );
  AOI222_X1 us12_U87 (.ZN( us12_n775 ) , .A1( us12_n830 ) , .C1( us12_n834 ) , .B2( us12_n841 ) , .A2( us12_n850 ) , .B1( us12_n861 ) , .C2( us12_n873 ) );
  NOR2_X1 us12_U88 (.ZN( us12_n625 ) , .A2( us12_n836 ) , .A1( us12_n839 ) );
  NOR2_X1 us12_U89 (.ZN( us12_n761 ) , .A1( us12_n833 ) , .A2( us12_n834 ) );
  NOR3_X1 us12_U9 (.A3( us12_n800 ) , .A2( us12_n801 ) , .A1( us12_n802 ) , .ZN( us12_n825 ) );
  AOI222_X1 us12_U90 (.ZN( us12_n513 ) , .C1( us12_n832 ) , .B2( us12_n837 ) , .A2( us12_n843 ) , .C2( us12_n862 ) , .B1( us12_n863 ) , .A1( us12_n866 ) );
  NOR4_X1 us12_U91 (.A4( us12_n509 ) , .A2( us12_n510 ) , .A1( us12_n511 ) , .ZN( us12_n512 ) , .A3( us12_n670 ) );
  INV_X1 us12_U92 (.A( us12_n505 ) , .ZN( us12_n871 ) );
  NAND4_X1 us12_U93 (.A4( us12_n456 ) , .A3( us12_n457 ) , .A2( us12_n458 ) , .A1( us12_n459 ) , .ZN( us12_n679 ) );
  NOR3_X1 us12_U94 (.ZN( us12_n457 ) , .A3( us12_n530 ) , .A1( us12_n555 ) , .A2( us12_n570 ) );
  AOI221_X1 us12_U95 (.A( us12_n450 ) , .ZN( us12_n459 ) , .C2( us12_n753 ) , .B1( us12_n832 ) , .C1( us12_n842 ) , .B2( us12_n861 ) );
  NOR4_X1 us12_U96 (.ZN( us12_n458 ) , .A2( us12_n509 ) , .A1( us12_n599 ) , .A4( us12_n628 ) , .A3( us12_n711 ) );
  NAND4_X1 us12_U97 (.A4( us12_n535 ) , .A3( us12_n536 ) , .A2( us12_n537 ) , .A1( us12_n538 ) , .ZN( us12_n622 ) );
  NOR4_X1 us12_U98 (.A4( us12_n526 ) , .A2( us12_n527 ) , .A1( us12_n528 ) , .ZN( us12_n538 ) , .A3( us12_n701 ) );
  NOR4_X1 us12_U99 (.A1( us12_n531 ) , .ZN( us12_n536 ) , .A2( us12_n654 ) , .A4( us12_n668 ) , .A3( us12_n765 ) );
  NOR3_X1 us21_U10 (.A3( us21_n619 ) , .A2( us21_n620 ) , .ZN( us21_n634 ) , .A1( us21_n723 ) );
  NOR4_X1 us21_U100 (.A4( us21_n524 ) , .A2( us21_n525 ) , .A1( us21_n526 ) , .ZN( us21_n536 ) , .A3( us21_n699 ) );
  NOR4_X1 us21_U101 (.A1( us21_n529 ) , .ZN( us21_n534 ) , .A2( us21_n652 ) , .A4( us21_n666 ) , .A3( us21_n763 ) );
  NOR4_X1 us21_U102 (.A4( us21_n527 ) , .A3( us21_n528 ) , .ZN( us21_n535 ) , .A2( us21_n682 ) , .A1( us21_n792 ) );
  NAND4_X1 us21_U103 (.A4( us21_n546 ) , .A3( us21_n547 ) , .A2( us21_n548 ) , .A1( us21_n549 ) , .ZN( us21_n743 ) );
  NOR3_X1 us21_U104 (.ZN( us21_n547 ) , .A2( us21_n649 ) , .A1( us21_n665 ) , .A3( us21_n769 ) );
  AOI211_X1 us21_U105 (.B( us21_n537 ) , .A( us21_n538 ) , .ZN( us21_n549 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NOR4_X1 us21_U106 (.A4( us21_n539 ) , .A3( us21_n540 ) , .A2( us21_n541 ) , .ZN( us21_n548 ) , .A1( us21_n686 ) );
  NAND4_X1 us21_U107 (.A4( us21_n477 ) , .A3( us21_n478 ) , .A2( us21_n479 ) , .A1( us21_n480 ) , .ZN( us21_n692 ) );
  NOR3_X1 us21_U108 (.ZN( us21_n478 ) , .A2( us21_n506 ) , .A3( us21_n599 ) , .A1( us21_n608 ) );
  AOI211_X1 us21_U109 (.B( us21_n475 ) , .A( us21_n476 ) , .ZN( us21_n480 ) , .C2( us21_n831 ) , .C1( us21_n859 ) );
  NOR2_X1 us21_U11 (.ZN( us21_n493 ) , .A1( us21_n676 ) , .A2( us21_n692 ) );
  NOR4_X1 us21_U110 (.ZN( us21_n479 ) , .A3( us21_n530 ) , .A4( us21_n543 ) , .A2( us21_n565 ) , .A1( us21_n715 ) );
  NOR4_X1 us21_U111 (.A4( us21_n607 ) , .A3( us21_n608 ) , .A2( us21_n609 ) , .A1( us21_n610 ) , .ZN( us21_n617 ) );
  NOR4_X1 us21_U112 (.ZN( us21_n618 ) , .A1( us21_n654 ) , .A3( us21_n664 ) , .A4( us21_n680 ) , .A2( us21_n764 ) );
  NOR4_X1 us21_U113 (.A4( us21_n612 ) , .A3( us21_n613 ) , .A2( us21_n614 ) , .A1( us21_n615 ) , .ZN( us21_n616 ) );
  NOR2_X1 us21_U114 (.ZN( us21_n684 ) , .A1( us21_n829 ) , .A2( us21_n830 ) );
  NAND4_X1 us21_U115 (.A4( us21_n471 ) , .A3( us21_n472 ) , .A2( us21_n473 ) , .A1( us21_n474 ) , .ZN( us21_n676 ) );
  NOR4_X1 us21_U116 (.A4( us21_n468 ) , .ZN( us21_n474 ) , .A3( us21_n554 ) , .A1( us21_n733 ) , .A2( us21_n753 ) );
  NOR4_X1 us21_U117 (.ZN( us21_n473 ) , .A1( us21_n529 ) , .A3( us21_n566 ) , .A4( us21_n598 ) , .A2( us21_n640 ) );
  NOR4_X1 us21_U118 (.ZN( us21_n472 ) , .A1( us21_n504 ) , .A3( us21_n542 ) , .A2( us21_n581 ) , .A4( us21_n714 ) );
  NAND4_X1 us21_U119 (.A4( us21_n689 ) , .A3( us21_n690 ) , .A1( us21_n691 ) , .ZN( us21_n774 ) , .A2( us21_n870 ) );
  NOR2_X1 us21_U12 (.A1( us21_n676 ) , .ZN( us21_n691 ) , .A2( us21_n805 ) );
  INV_X1 us21_U120 (.A( us21_n677 ) , .ZN( us21_n870 ) );
  AOI221_X1 us21_U121 (.A( us21_n679 ) , .ZN( us21_n690 ) , .B2( us21_n838 ) , .C1( us21_n840 ) , .C2( us21_n860 ) , .B1( us21_n863 ) );
  NOR4_X1 us21_U122 (.A4( us21_n685 ) , .A3( us21_n686 ) , .A2( us21_n687 ) , .A1( us21_n688 ) , .ZN( us21_n689 ) );
  NOR2_X1 us21_U123 (.ZN( us21_n731 ) , .A2( us21_n830 ) , .A1( us21_n843 ) );
  NAND4_X1 us21_U124 (.A4( us21_n717 ) , .A3( us21_n718 ) , .A2( us21_n719 ) , .ZN( us21_n739 ) , .A1( us21_n855 ) );
  INV_X1 us21_U125 (.A( us21_n707 ) , .ZN( us21_n855 ) );
  NOR4_X1 us21_U126 (.A4( us21_n713 ) , .A3( us21_n714 ) , .A2( us21_n715 ) , .A1( us21_n716 ) , .ZN( us21_n717 ) );
  AOI221_X1 us21_U127 (.A( us21_n708 ) , .ZN( us21_n719 ) , .C2( us21_n842 ) , .B2( us21_n843 ) , .C1( us21_n859 ) , .B1( us21_n860 ) );
  NAND4_X1 us21_U128 (.A4( us21_n571 ) , .A3( us21_n572 ) , .A1( us21_n573 ) , .ZN( us21_n721 ) , .A2( us21_n872 ) );
  NOR4_X1 us21_U129 (.A4( us21_n567 ) , .A3( us21_n568 ) , .A2( us21_n569 ) , .A1( us21_n570 ) , .ZN( us21_n571 ) );
  INV_X1 us21_U13 (.A( us21_n605 ) , .ZN( us21_n872 ) );
  AOI221_X1 us21_U130 (.A( us21_n562 ) , .C2( us21_n563 ) , .ZN( us21_n572 ) , .B2( us21_n843 ) , .B1( us21_n850 ) , .C1( us21_n851 ) );
  NOR2_X1 us21_U131 (.ZN( us21_n573 ) , .A1( us21_n620 ) , .A2( us21_n743 ) );
  NAND4_X1 us21_U132 (.A4( us21_n491 ) , .A3( us21_n492 ) , .A1( us21_n493 ) , .ZN( us21_n800 ) , .A2( us21_n865 ) );
  AOI221_X1 us21_U133 (.A( us21_n487 ) , .ZN( us21_n492 ) , .B2( us21_n834 ) , .C2( us21_n839 ) , .C1( us21_n849 ) , .B1( us21_n858 ) );
  INV_X1 us21_U134 (.A( us21_n776 ) , .ZN( us21_n865 ) );
  NOR4_X1 us21_U135 (.A2( us21_n489 ) , .A1( us21_n490 ) , .ZN( us21_n491 ) , .A3( us21_n578 ) , .A4( us21_n610 ) );
  INV_X1 us21_U136 (.A( us21_n760 ) , .ZN( us21_n828 ) );
  NOR2_X1 us21_U137 (.ZN( us21_n645 ) , .A1( us21_n852 ) , .A2( us21_n866 ) );
  INV_X1 us21_U138 (.A( us21_n461 ) , .ZN( us21_n862 ) );
  OAI21_X1 us21_U139 (.ZN( us21_n461 ) , .B1( us21_n807 ) , .A( us21_n832 ) , .B2( us21_n849 ) );
  INV_X1 us21_U14 (.A( us21_n678 ) , .ZN( us21_n838 ) );
  OR4_X1 us21_U140 (.ZN( us21_n490 ) , .A4( us21_n532 ) , .A2( us21_n545 ) , .A1( us21_n557 ) , .A3( us21_n630 ) );
  OR4_X1 us21_U141 (.A4( us21_n564 ) , .A3( us21_n565 ) , .A2( us21_n566 ) , .ZN( us21_n570 ) , .A1( us21_n663 ) );
  OR4_X1 us21_U142 (.A4( us21_n680 ) , .A3( us21_n681 ) , .A2( us21_n682 ) , .A1( us21_n683 ) , .ZN( us21_n688 ) );
  OR4_X1 us21_U143 (.ZN( us21_n464 ) , .A4( us21_n516 ) , .A3( us21_n527 ) , .A2( us21_n576 ) , .A1( us21_n710 ) );
  OR4_X1 us21_U144 (.A4( us21_n516 ) , .A2( us21_n517 ) , .A1( us21_n518 ) , .ZN( us21_n520 ) , .A3( us21_n819 ) );
  OR4_X1 us21_U145 (.A4( us21_n578 ) , .A3( us21_n579 ) , .A2( us21_n580 ) , .A1( us21_n581 ) , .ZN( us21_n582 ) );
  NAND2_X1 us21_U146 (.ZN( us21_n611 ) , .A2( us21_n835 ) , .A1( us21_n871 ) );
  OR3_X1 us21_U147 (.A3( us21_n504 ) , .A2( us21_n505 ) , .A1( us21_n506 ) , .ZN( us21_n509 ) );
  AOI221_X1 us21_U148 (.A( us21_n711 ) , .B2( us21_n712 ) , .ZN( us21_n718 ) , .C1( us21_n830 ) , .B1( us21_n837 ) , .C2( us21_n861 ) );
  OR2_X1 us21_U149 (.A2( us21_n709 ) , .A1( us21_n710 ) , .ZN( us21_n711 ) );
  NOR4_X1 us21_U15 (.A4( us21_n443 ) , .A3( us21_n444 ) , .A2( us21_n514 ) , .A1( us21_n539 ) , .ZN( us21_n704 ) );
  INV_X1 us21_U150 (.A( us21_n752 ) , .ZN( us21_n867 ) );
  OAI21_X1 us21_U151 (.B1( us21_n751 ) , .ZN( us21_n752 ) , .A( us21_n843 ) , .B2( us21_n866 ) );
  INV_X1 us21_U152 (.A( us21_n670 ) , .ZN( us21_n857 ) );
  AOI21_X1 us21_U153 (.A( us21_n668 ) , .B1( us21_n669 ) , .ZN( us21_n670 ) , .B2( us21_n854 ) );
  AOI222_X1 us21_U154 (.ZN( us21_n658 ) , .A2( us21_n837 ) , .B1( us21_n839 ) , .C2( us21_n843 ) , .A1( us21_n858 ) , .C1( us21_n861 ) , .B2( us21_n868 ) );
  INV_X1 us21_U155 (.A( us21_n645 ) , .ZN( us21_n868 ) );
  OAI22_X1 us21_U156 (.ZN( us21_n481 ) , .A1( us21_n706 ) , .B2( us21_n783 ) , .A2( us21_n804 ) , .B1( us21_n810 ) );
  OAI22_X1 us21_U157 (.ZN( us21_n635 ) , .A1( us21_n697 ) , .B2( us21_n726 ) , .A2( us21_n760 ) , .B1( us21_n814 ) );
  OAI222_X1 us21_U158 (.B2( us21_n706 ) , .ZN( us21_n707 ) , .C2( us21_n722 ) , .B1( us21_n745 ) , .A1( us21_n804 ) , .C1( us21_n812 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U159 (.A1( us21_n445 ) , .A2( us21_n463 ) , .ZN( us21_n747 ) );
  OR3_X1 us21_U16 (.ZN( us21_n444 ) , .A1( us21_n526 ) , .A3( us21_n575 ) , .A2( us21_n873 ) );
  AOI22_X1 us21_U160 (.ZN( us21_n694 ) , .A1( us21_n828 ) , .B2( us21_n841 ) , .A2( us21_n863 ) , .B1( us21_n866 ) );
  INV_X1 us21_U161 (.A( us21_n728 ) , .ZN( us21_n837 ) );
  NAND2_X1 us21_U162 (.A1( us21_n449 ) , .A2( us21_n451 ) , .ZN( us21_n760 ) );
  INV_X1 us21_U163 (.A( us21_n788 ) , .ZN( us21_n830 ) );
  OAI221_X1 us21_U164 (.A( us21_n725 ) , .C2( us21_n726 ) , .B2( us21_n727 ) , .B1( us21_n728 ) , .ZN( us21_n735 ) , .C1( us21_n815 ) );
  AOI22_X1 us21_U165 (.ZN( us21_n725 ) , .B1( us21_n830 ) , .A2( us21_n836 ) , .A1( us21_n861 ) , .B2( us21_n864 ) );
  AND2_X1 us21_U166 (.ZN( us21_n746 ) , .A1( us21_n782 ) , .A2( us21_n784 ) );
  OAI22_X1 us21_U167 (.ZN( us21_n487 ) , .A1( us21_n722 ) , .B2( us21_n726 ) , .B1( us21_n728 ) , .A2( us21_n777 ) );
  OAI22_X1 us21_U168 (.ZN( us21_n622 ) , .B1( us21_n667 ) , .B2( us21_n745 ) , .A1( us21_n813 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U169 (.B2( us21_n777 ) , .B1( us21_n778 ) , .ZN( us21_n779 ) , .A2( us21_n812 ) , .A1( us21_n813 ) );
  OR4_X1 us21_U17 (.A4( us21_n440 ) , .A2( us21_n441 ) , .A1( us21_n442 ) , .ZN( us21_n443 ) , .A3( us21_n551 ) );
  OAI22_X1 us21_U170 (.A1( us21_n722 ) , .ZN( us21_n724 ) , .B2( us21_n748 ) , .B1( us21_n810 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U171 (.B2( us21_n742 ) , .ZN( us21_n744 ) , .A2( us21_n760 ) , .B1( us21_n778 ) , .A1( us21_n790 ) );
  OAI22_X1 us21_U172 (.B2( us21_n801 ) , .B1( us21_n802 ) , .A2( us21_n803 ) , .A1( us21_n804 ) , .ZN( us21_n806 ) );
  OAI22_X1 us21_U173 (.ZN( us21_n494 ) , .A2( us21_n742 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n804 ) );
  INV_X1 us21_U174 (.A( us21_n742 ) , .ZN( us21_n835 ) );
  INV_X1 us21_U175 (.A( us21_n786 ) , .ZN( us21_n843 ) );
  INV_X1 us21_U176 (.A( us21_n814 ) , .ZN( us21_n829 ) );
  OAI22_X1 us21_U177 (.B1( us21_n488 ) , .ZN( us21_n489 ) , .A1( us21_n684 ) , .A2( us21_n761 ) , .B2( us21_n815 ) );
  NOR3_X1 us21_U178 (.ZN( us21_n488 ) , .A1( us21_n780 ) , .A2( us21_n848 ) , .A3( us21_n861 ) );
  OAI22_X1 us21_U179 (.ZN( us21_n588 ) , .B1( us21_n728 ) , .B2( us21_n747 ) , .A2( us21_n784 ) , .A1( us21_n801 ) );
  INV_X1 us21_U18 (.A( us21_n611 ) , .ZN( us21_n873 ) );
  OAI22_X1 us21_U180 (.ZN( us21_n693 ) , .A2( us21_n728 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n815 ) );
  OAI22_X1 us21_U181 (.ZN( us21_n708 ) , .A2( us21_n726 ) , .B2( us21_n727 ) , .A1( us21_n742 ) , .B1( us21_n811 ) );
  INV_X1 us21_U182 (.A( us21_n812 ) , .ZN( us21_n831 ) );
  INV_X1 us21_U183 (.A( us21_n667 ) , .ZN( us21_n863 ) );
  NOR2_X1 us21_U184 (.ZN( us21_n716 ) , .A2( us21_n722 ) , .A1( us21_n742 ) );
  NOR2_X1 us21_U185 (.ZN( us21_n664 ) , .A1( us21_n726 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U186 (.ZN( us21_n568 ) , .A1( us21_n726 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U187 (.ZN( us21_n544 ) , .A2( us21_n778 ) , .A1( us21_n812 ) );
  INV_X1 us21_U188 (.A( us21_n748 ) , .ZN( us21_n840 ) );
  NOR2_X1 us21_U189 (.ZN( us21_n530 ) , .A2( us21_n747 ) , .A1( us21_n748 ) );
  INV_X1 us21_U19 (.A( us21_n747 ) , .ZN( us21_n861 ) );
  NOR2_X1 us21_U190 (.ZN( us21_n575 ) , .A2( us21_n697 ) , .A1( us21_n812 ) );
  NOR2_X1 us21_U191 (.ZN( us21_n652 ) , .A1( us21_n726 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U192 (.ZN( us21_n613 ) , .A1( us21_n783 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U193 (.ZN( us21_n627 ) , .A2( us21_n726 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U194 (.ZN( us21_n599 ) , .A2( us21_n778 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U195 (.ZN( us21_n610 ) , .A1( us21_n777 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U196 (.ZN( us21_n526 ) , .A2( us21_n722 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U197 (.ZN( us21_n626 ) , .A2( us21_n667 ) , .A1( us21_n783 ) );
  INV_X1 us21_U198 (.A( us21_n790 ) , .ZN( us21_n849 ) );
  NOR2_X1 us21_U199 (.A2( us21_n742 ) , .ZN( us21_n767 ) , .A1( us21_n810 ) );
  AOI222_X1 us21_U20 (.ZN( us21_n561 ) , .B1( us21_n828 ) , .C1( us21_n839 ) , .A2( us21_n841 ) , .A1( us21_n852 ) , .B2( us21_n861 ) , .C2( us21_n871 ) );
  NOR2_X1 us21_U200 (.ZN( us21_n529 ) , .A2( us21_n778 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U201 (.A2( us21_n706 ) , .A1( us21_n748 ) , .ZN( us21_n769 ) );
  NOR2_X1 us21_U202 (.ZN( us21_n597 ) , .A2( us21_n789 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U203 (.ZN( us21_n609 ) , .A2( us21_n778 ) , .A1( us21_n804 ) );
  NOR2_X1 us21_U204 (.ZN( us21_n650 ) , .A1( us21_n667 ) , .A2( us21_n812 ) );
  INV_X1 us21_U205 (.A( us21_n745 ) , .ZN( us21_n832 ) );
  NOR2_X1 us21_U206 (.A1( us21_n667 ) , .ZN( us21_n671 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U207 (.ZN( us21_n600 ) , .A1( us21_n667 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U208 (.A1( us21_n667 ) , .ZN( us21_n686 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U209 (.ZN( us21_n665 ) , .A1( us21_n748 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U21 (.ZN( us21_n471 ) , .A2( us21_n519 ) , .A4( us21_n592 ) , .A1( us21_n607 ) , .A3( us21_n627 ) );
  NOR2_X1 us21_U210 (.ZN( us21_n553 ) , .A1( us21_n748 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U211 (.ZN( us21_n506 ) , .A2( us21_n778 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U212 (.ZN( us21_n541 ) , .A2( us21_n706 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U213 (.ZN( us21_n662 ) , .A1( us21_n783 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U214 (.A1( us21_n667 ) , .ZN( us21_n764 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U215 (.A1( us21_n697 ) , .ZN( us21_n766 ) , .A2( us21_n811 ) );
  OAI22_X1 us21_U216 (.B1( us21_n438 ) , .ZN( us21_n442 ) , .A2( us21_n726 ) , .A1( us21_n742 ) , .B2( us21_n747 ) );
  NOR3_X1 us21_U217 (.ZN( us21_n438 ) , .A2( us21_n834 ) , .A3( us21_n835 ) , .A1( us21_n844 ) );
  NOR2_X1 us21_U218 (.ZN( us21_n525 ) , .A1( us21_n667 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U219 (.ZN( us21_n505 ) , .A1( us21_n810 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U22 (.A4( us21_n542 ) , .A3( us21_n543 ) , .A2( us21_n544 ) , .A1( us21_n545 ) , .ZN( us21_n546 ) );
  NOR2_X1 us21_U220 (.ZN( us21_n659 ) , .A1( us21_n727 ) , .A2( us21_n788 ) );
  INV_X1 us21_U221 (.A( us21_n801 ) , .ZN( us21_n841 ) );
  NOR2_X1 us21_U222 (.ZN( us21_n555 ) , .A1( us21_n790 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U223 (.ZN( us21_n543 ) , .A1( us21_n747 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U224 (.ZN( us21_n507 ) , .A1( us21_n727 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U225 (.ZN( us21_n528 ) , .A2( us21_n742 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U226 (.A1( us21_n747 ) , .ZN( us21_n765 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U227 (.A2( us21_n742 ) , .ZN( us21_n753 ) , .A1( us21_n803 ) );
  OAI22_X1 us21_U228 (.B2( us21_n748 ) , .B1( us21_n749 ) , .A1( us21_n750 ) , .ZN( us21_n754 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U229 (.ZN( us21_n749 ) , .A2( us21_n850 ) , .A1( us21_n858 ) );
  NOR4_X1 us21_U23 (.ZN( us21_n477 ) , .A1( us21_n518 ) , .A4( us21_n555 ) , .A3( us21_n580 ) , .A2( us21_n628 ) );
  NOR3_X1 us21_U230 (.ZN( us21_n750 ) , .A2( us21_n851 ) , .A1( us21_n861 ) , .A3( us21_n863 ) );
  NOR2_X1 us21_U231 (.ZN( us21_n542 ) , .A2( us21_n783 ) , .A1( us21_n790 ) );
  INV_X1 us21_U232 (.A( us21_n804 ) , .ZN( us21_n839 ) );
  NOR2_X1 us21_U233 (.ZN( us21_n629 ) , .A1( us21_n722 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U234 (.ZN( us21_n733 ) , .A2( us21_n801 ) , .A1( us21_n803 ) );
  NOR2_X1 us21_U235 (.ZN( us21_n514 ) , .A1( us21_n706 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U236 (.ZN( us21_n661 ) , .A1( us21_n727 ) , .A2( us21_n783 ) );
  NOR2_X1 us21_U237 (.ZN( us21_n715 ) , .A2( us21_n742 ) , .A1( us21_n784 ) );
  NOR2_X1 us21_U238 (.ZN( us21_n612 ) , .A1( us21_n760 ) , .A2( us21_n810 ) );
  INV_X1 us21_U239 (.A( us21_n726 ) , .ZN( us21_n850 ) );
  NOR4_X1 us21_U24 (.ZN( us21_n454 ) , .A2( us21_n515 ) , .A1( us21_n541 ) , .A3( us21_n577 ) , .A4( us21_n613 ) );
  NOR2_X1 us21_U240 (.ZN( us21_n552 ) , .A1( us21_n784 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U241 (.ZN( us21_n515 ) , .A1( us21_n706 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U242 (.ZN( us21_n504 ) , .A2( us21_n726 ) , .A1( us21_n760 ) );
  NOR2_X1 us21_U243 (.ZN( us21_n556 ) , .A1( us21_n706 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U244 (.ZN( us21_n519 ) , .A1( us21_n788 ) , .A2( us21_n810 ) );
  INV_X1 us21_U245 (.A( us21_n803 ) , .ZN( us21_n858 ) );
  NOR2_X1 us21_U246 (.ZN( us21_n713 ) , .A1( us21_n803 ) , .A2( us21_n815 ) );
  NOR2_X1 us21_U247 (.ZN( us21_n653 ) , .A1( us21_n788 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U248 (.ZN( us21_n666 ) , .A2( us21_n706 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U249 (.ZN( us21_n628 ) , .A1( us21_n745 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U25 (.A4( us21_n530 ) , .A3( us21_n531 ) , .A2( us21_n532 ) , .ZN( us21_n533 ) , .A1( us21_n818 ) );
  NOR2_X1 us21_U250 (.ZN( us21_n554 ) , .A1( us21_n760 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U251 (.ZN( us21_n540 ) , .A1( us21_n760 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U252 (.ZN( us21_n699 ) , .A2( us21_n784 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U253 (.A1( us21_n728 ) , .ZN( us21_n763 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U254 (.ZN( us21_n607 ) , .A2( us21_n722 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U255 (.ZN( us21_n577 ) , .A2( us21_n706 ) , .A1( us21_n728 ) );
  NOR2_X1 us21_U256 (.ZN( us21_n531 ) , .A2( us21_n722 ) , .A1( us21_n728 ) );
  AOI21_X1 us21_U257 (.A( us21_n810 ) , .B2( us21_n811 ) , .B1( us21_n812 ) , .ZN( us21_n817 ) );
  AOI21_X1 us21_U258 (.ZN( us21_n513 ) , .A( us21_n727 ) , .B1( us21_n748 ) , .B2( us21_n801 ) );
  NOR2_X1 us21_U259 (.ZN( us21_n654 ) , .A1( us21_n745 ) , .A2( us21_n778 ) );
  NOR2_X1 us21_U26 (.ZN( us21_n678 ) , .A2( us21_n832 ) , .A1( us21_n837 ) );
  AOI21_X1 us21_U260 (.A( us21_n813 ) , .B2( us21_n814 ) , .B1( us21_n815 ) , .ZN( us21_n816 ) );
  NOR2_X1 us21_U261 (.ZN( us21_n580 ) , .A1( us21_n742 ) , .A2( us21_n813 ) );
  AOI21_X1 us21_U262 (.ZN( us21_n591 ) , .B1( us21_n748 ) , .A( us21_n790 ) , .B2( us21_n811 ) );
  AOI21_X1 us21_U263 (.B1( us21_n623 ) , .ZN( us21_n625 ) , .A( us21_n761 ) , .B2( us21_n812 ) );
  NOR2_X1 us21_U264 (.A2( us21_n706 ) , .A1( us21_n760 ) , .ZN( us21_n792 ) );
  NOR2_X1 us21_U265 (.ZN( us21_n640 ) , .A2( us21_n786 ) , .A1( us21_n789 ) );
  AOI21_X1 us21_U266 (.ZN( us21_n497 ) , .B1( us21_n678 ) , .A( us21_n810 ) , .B2( us21_n814 ) );
  NOR2_X1 us21_U267 (.ZN( us21_n668 ) , .A1( us21_n788 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U268 (.ZN( us21_n557 ) , .A2( us21_n789 ) , .A1( us21_n801 ) );
  AOI21_X1 us21_U269 (.ZN( us21_n624 ) , .B2( us21_n667 ) , .A( us21_n788 ) , .B1( us21_n789 ) );
  NOR4_X1 us21_U27 (.A4( us21_n575 ) , .A3( us21_n576 ) , .A2( us21_n577 ) , .ZN( us21_n584 ) , .A1( us21_n681 ) );
  NOR2_X1 us21_U270 (.ZN( us21_n681 ) , .A2( us21_n697 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U271 (.ZN( us21_n651 ) , .A1( us21_n760 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U272 (.ZN( us21_n518 ) , .A2( us21_n706 ) , .A1( us21_n812 ) );
  INV_X1 us21_U273 (.A( us21_n811 ) , .ZN( us21_n834 ) );
  NOR2_X1 us21_U274 (.ZN( us21_n517 ) , .A2( us21_n697 ) , .A1( us21_n814 ) );
  AOI21_X1 us21_U275 (.ZN( us21_n475 ) , .A( us21_n667 ) , .B1( us21_n748 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U276 (.ZN( us21_n508 ) , .B2( us21_n667 ) , .A( us21_n728 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U277 (.ZN( us21_n537 ) , .B2( us21_n810 ) , .A( us21_n812 ) , .B1( us21_n813 ) );
  INV_X1 us21_U278 (.A( us21_n761 ) , .ZN( us21_n864 ) );
  AOI21_X1 us21_U279 (.ZN( us21_n538 ) , .A( us21_n761 ) , .B2( us21_n777 ) , .B1( us21_n815 ) );
  NOR4_X1 us21_U28 (.A1( us21_n582 ) , .ZN( us21_n583 ) , .A3( us21_n650 ) , .A2( us21_n660 ) , .A4( us21_n765 ) );
  NOR2_X1 us21_U280 (.ZN( us21_n579 ) , .A1( us21_n667 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U281 (.ZN( us21_n587 ) , .B2( us21_n697 ) , .B1( us21_n813 ) , .A( us21_n815 ) );
  AOI21_X1 us21_U282 (.ZN( us21_n589 ) , .B2( us21_n761 ) , .A( us21_n783 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U283 (.B1( us21_n697 ) , .ZN( us21_n698 ) , .A( us21_n730 ) , .B2( us21_n761 ) );
  AOI21_X1 us21_U284 (.ZN( us21_n638 ) , .B2( us21_n745 ) , .A( us21_n790 ) , .B1( us21_n801 ) );
  AOI21_X1 us21_U285 (.ZN( us21_n496 ) , .A( us21_n722 ) , .B2( us21_n760 ) , .B1( us21_n812 ) );
  INV_X1 us21_U286 (.A( us21_n789 ) , .ZN( us21_n871 ) );
  NOR2_X1 us21_U287 (.ZN( us21_n545 ) , .A1( us21_n697 ) , .A2( us21_n742 ) );
  INV_X1 us21_U288 (.A( us21_n727 ) , .ZN( us21_n866 ) );
  AOI21_X1 us21_U289 (.ZN( us21_n647 ) , .B1( us21_n727 ) , .B2( us21_n761 ) , .A( us21_n811 ) );
  AOI221_X1 us21_U29 (.A( us21_n779 ) , .ZN( us21_n796 ) , .C2( us21_n835 ) , .B2( us21_n836 ) , .B1( us21_n863 ) , .C1( us21_n864 ) );
  AOI21_X1 us21_U290 (.ZN( us21_n567 ) , .B1( us21_n748 ) , .B2( us21_n760 ) , .A( us21_n778 ) );
  INV_X1 us21_U291 (.A( us21_n810 ) , .ZN( us21_n852 ) );
  NOR2_X1 us21_U292 (.ZN( us21_n683 ) , .A1( us21_n727 ) , .A2( us21_n814 ) );
  AOI21_X1 us21_U293 (.B1( us21_n684 ) , .ZN( us21_n685 ) , .A( us21_n726 ) , .B2( us21_n759 ) );
  NOR2_X1 us21_U294 (.ZN( us21_n566 ) , .A1( us21_n727 ) , .A2( us21_n760 ) );
  NOR2_X1 us21_U295 (.ZN( us21_n663 ) , .A1( us21_n778 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U296 (.ZN( us21_n448 ) , .B2( us21_n790 ) , .A( us21_n801 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U297 (.ZN( us21_n512 ) , .A( us21_n777 ) , .B2( us21_n790 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U298 (.ZN( us21_n637 ) , .B2( us21_n747 ) , .A( us21_n786 ) , .B1( us21_n810 ) );
  INV_X1 us21_U299 (.A( us21_n697 ) , .ZN( us21_n851 ) );
  NAND2_X2 us21_U3 (.A2( us21_n458 ) , .A1( us21_n463 ) , .ZN( us21_n778 ) );
  NOR4_X1 us21_U30 (.A4( us21_n791 ) , .A3( us21_n792 ) , .A2( us21_n793 ) , .A1( us21_n794 ) , .ZN( us21_n795 ) );
  AOI21_X1 us21_U300 (.ZN( us21_n562 ) , .B1( us21_n722 ) , .A( us21_n777 ) , .B2( us21_n789 ) );
  NOR2_X1 us21_U301 (.ZN( us21_n576 ) , .A1( us21_n706 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U302 (.ZN( us21_n527 ) , .A1( us21_n706 ) , .A2( us21_n777 ) );
  AOI21_X1 us21_U303 (.ZN( us21_n687 ) , .B2( us21_n747 ) , .B1( us21_n761 ) , .A( us21_n804 ) );
  NOR2_X1 us21_U304 (.ZN( us21_n682 ) , .A1( us21_n789 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U305 (.ZN( us21_n648 ) , .A( us21_n777 ) , .B1( us21_n790 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U306 (.A2( us21_n811 ) , .A1( us21_n813 ) , .ZN( us21_n819 ) );
  AOI21_X1 us21_U307 (.A( us21_n788 ) , .B2( us21_n789 ) , .B1( us21_n790 ) , .ZN( us21_n791 ) );
  AOI21_X1 us21_U308 (.A( us21_n731 ) , .ZN( us21_n732 ) , .B2( us21_n778 ) , .B1( us21_n790 ) );
  NOR2_X1 us21_U309 (.ZN( us21_n581 ) , .A1( us21_n790 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U31 (.A4( us21_n774 ) , .A3( us21_n775 ) , .A1( us21_n776 ) , .ZN( us21_n797 ) , .A2( us21_n799 ) );
  NOR2_X1 us21_U310 (.ZN( us21_n532 ) , .A1( us21_n722 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U311 (.ZN( us21_n639 ) , .B1( us21_n678 ) , .A( us21_n789 ) , .B2( us21_n815 ) );
  NOR2_X1 us21_U312 (.ZN( us21_n709 ) , .A1( us21_n760 ) , .A2( us21_n761 ) );
  NOR2_X1 us21_U313 (.ZN( us21_n565 ) , .A1( us21_n745 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U314 (.ZN( us21_n680 ) , .A2( us21_n706 ) , .A1( us21_n815 ) );
  INV_X1 us21_U315 (.A( us21_n813 ) , .ZN( us21_n853 ) );
  AOI21_X1 us21_U316 (.ZN( us21_n440 ) , .A( us21_n697 ) , .B1( us21_n731 ) , .B2( us21_n748 ) );
  INV_X1 us21_U317 (.A( us21_n778 ) , .ZN( us21_n848 ) );
  AOI22_X1 us21_U318 (.A2( us21_n780 ) , .ZN( us21_n781 ) , .B2( us21_n829 ) , .A1( us21_n832 ) , .B1( us21_n861 ) );
  NAND2_X1 us21_U319 (.ZN( us21_n712 ) , .A1( us21_n726 ) , .A2( us21_n778 ) );
  NOR4_X1 us21_U32 (.A3( us21_n753 ) , .A2( us21_n754 ) , .A1( us21_n755 ) , .ZN( us21_n756 ) , .A4( us21_n867 ) );
  NAND2_X1 us21_U320 (.ZN( us21_n751 ) , .A1( us21_n761 ) , .A2( us21_n803 ) );
  AOI21_X1 us21_U321 (.ZN( us21_n441 ) , .B1( us21_n787 ) , .B2( us21_n789 ) , .A( us21_n812 ) );
  INV_X1 us21_U322 (.A( us21_n783 ) , .ZN( us21_n844 ) );
  AOI21_X1 us21_U323 (.ZN( us21_n495 ) , .A( us21_n777 ) , .B2( us21_n789 ) , .B1( us21_n802 ) );
  NAND2_X1 us21_U324 (.A2( us21_n760 ) , .A1( us21_n804 ) , .ZN( us21_n808 ) );
  NOR2_X1 us21_U325 (.ZN( us21_n468 ) , .A2( us21_n777 ) , .A1( us21_n813 ) );
  NOR2_X1 us21_U326 (.ZN( us21_n710 ) , .A2( us21_n722 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U327 (.ZN( us21_n482 ) , .A1( us21_n786 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U328 (.ZN( us21_n524 ) , .A1( us21_n722 ) , .A2( us21_n748 ) );
  OAI21_X1 us21_U329 (.A( us21_n729 ) , .B1( us21_n730 ) , .ZN( us21_n734 ) , .B2( us21_n803 ) );
  AOI211_X1 us21_U33 (.B( us21_n743 ) , .A( us21_n744 ) , .ZN( us21_n757 ) , .C1( us21_n830 ) , .C2( us21_n851 ) );
  OAI21_X1 us21_U330 (.ZN( us21_n729 ) , .A( us21_n831 ) , .B2( us21_n850 ) , .B1( us21_n871 ) );
  OAI21_X1 us21_U331 (.A( us21_n785 ) , .B2( us21_n786 ) , .B1( us21_n787 ) , .ZN( us21_n793 ) );
  OAI21_X1 us21_U332 (.ZN( us21_n785 ) , .A( us21_n837 ) , .B1( us21_n861 ) , .B2( us21_n871 ) );
  NAND2_X1 us21_U333 (.A1( us21_n697 ) , .A2( us21_n727 ) , .ZN( us21_n780 ) );
  NOR2_X1 us21_U334 (.ZN( us21_n516 ) , .A1( us21_n706 ) , .A2( us21_n786 ) );
  NAND2_X1 us21_U335 (.ZN( us21_n669 ) , .A1( us21_n804 ) , .A2( us21_n814 ) );
  OAI21_X1 us21_U336 (.A( us21_n696 ) , .ZN( us21_n700 ) , .B2( us21_n748 ) , .B1( us21_n802 ) );
  OAI21_X1 us21_U337 (.ZN( us21_n696 ) , .B2( us21_n831 ) , .B1( us21_n836 ) , .A( us21_n858 ) );
  NAND2_X1 us21_U338 (.A2( us21_n747 ) , .A1( us21_n784 ) , .ZN( us21_n807 ) );
  INV_X1 us21_U339 (.A( us21_n722 ) , .ZN( us21_n854 ) );
  NOR3_X1 us21_U34 (.A3( us21_n739 ) , .A2( us21_n740 ) , .A1( us21_n741 ) , .ZN( us21_n758 ) );
  INV_X1 us21_U340 (.A( us21_n815 ) , .ZN( us21_n842 ) );
  AND2_X1 us21_U341 (.ZN( us21_n730 ) , .A1( us21_n777 ) , .A2( us21_n783 ) );
  OAI222_X1 us21_U342 (.ZN( us21_n615 ) , .B1( us21_n695 ) , .C1( us21_n722 ) , .C2( us21_n745 ) , .B2( us21_n784 ) , .A2( us21_n790 ) , .A1( us21_n814 ) );
  AOI221_X1 us21_U343 (.A( us21_n762 ) , .ZN( us21_n772 ) , .C2( us21_n808 ) , .B2( us21_n833 ) , .C1( us21_n853 ) , .B1( us21_n864 ) );
  AOI21_X1 us21_U344 (.B2( us21_n761 ) , .ZN( us21_n762 ) , .A( us21_n786 ) , .B1( us21_n790 ) );
  INV_X1 us21_U345 (.A( us21_n759 ) , .ZN( us21_n833 ) );
  NAND2_X2 us21_U346 (.A2( us21_n439 ) , .A1( us21_n445 ) , .ZN( us21_n782 ) );
  NAND2_X1 us21_U347 (.A1( us21_n453 ) , .A2( us21_n469 ) , .ZN( us21_n801 ) );
  NAND2_X1 us21_U348 (.A1( us21_n452 ) , .A2( us21_n459 ) , .ZN( us21_n811 ) );
  NAND2_X1 us21_U349 (.A1( us21_n451 ) , .A2( us21_n459 ) , .ZN( us21_n742 ) );
  NOR4_X1 us21_U35 (.A4( us21_n732 ) , .A3( us21_n733 ) , .A2( us21_n734 ) , .A1( us21_n735 ) , .ZN( us21_n736 ) );
  NAND2_X1 us21_U350 (.A1( us21_n449 ) , .A2( us21_n452 ) , .ZN( us21_n812 ) );
  NAND2_X1 us21_U351 (.A1( us21_n453 ) , .A2( us21_n460 ) , .ZN( us21_n748 ) );
  NAND2_X1 us21_U352 (.A1( us21_n449 ) , .A2( us21_n469 ) , .ZN( us21_n814 ) );
  NAND2_X1 us21_U353 (.A1( us21_n450 ) , .A2( us21_n463 ) , .ZN( us21_n667 ) );
  NAND2_X1 us21_U354 (.A2( us21_n446 ) , .A1( us21_n458 ) , .ZN( us21_n726 ) );
  NAND2_X1 us21_U355 (.A1( us21_n451 ) , .A2( us21_n470 ) , .ZN( us21_n783 ) );
  NAND2_X1 us21_U356 (.A2( us21_n452 ) , .A1( us21_n470 ) , .ZN( us21_n777 ) );
  NAND2_X1 us21_U357 (.A2( us21_n451 ) , .A1( us21_n453 ) , .ZN( us21_n804 ) );
  NAND2_X1 us21_U358 (.A2( us21_n462 ) , .A1( us21_n463 ) , .ZN( us21_n810 ) );
  NAND2_X1 us21_U359 (.A1( us21_n439 ) , .A2( us21_n458 ) , .ZN( us21_n697 ) );
  AOI211_X1 us21_U36 (.B( us21_n723 ) , .A( us21_n724 ) , .ZN( us21_n737 ) , .C1( us21_n841 ) , .C2( us21_n853 ) );
  NAND2_X1 us21_U360 (.A2( us21_n447 ) , .A1( us21_n450 ) , .ZN( us21_n761 ) );
  NAND2_X1 us21_U361 (.A2( us21_n446 ) , .A1( us21_n450 ) , .ZN( us21_n727 ) );
  NOR2_X1 us21_U362 (.ZN( us21_n445 ) , .A2( us21_n847 ) , .A1( us21_n856 ) );
  NAND2_X1 us21_U363 (.A1( us21_n460 ) , .A2( us21_n470 ) , .ZN( us21_n786 ) );
  NOR2_X1 us21_U364 (.ZN( us21_n463 ) , .A2( us21_n845 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U365 (.ZN( us21_n451 ) , .A1( us21_n824 ) , .A2( us21_n825 ) );
  NAND2_X1 us21_U366 (.A2( us21_n459 ) , .A1( us21_n460 ) , .ZN( us21_n745 ) );
  NOR2_X1 us21_U367 (.ZN( us21_n449 ) , .A1( us21_n826 ) , .A2( us21_n827 ) );
  NAND2_X1 us21_U368 (.A2( us21_n459 ) , .A1( us21_n469 ) , .ZN( us21_n695 ) );
  NAND2_X1 us21_U369 (.A2( us21_n452 ) , .A1( us21_n453 ) , .ZN( us21_n728 ) );
  NOR3_X1 us21_U37 (.A3( us21_n720 ) , .A1( us21_n721 ) , .ZN( us21_n738 ) , .A2( us21_n739 ) );
  NAND2_X1 us21_U370 (.A1( us21_n449 ) , .A2( us21_n460 ) , .ZN( us21_n788 ) );
  NAND2_X2 us21_U371 (.A2( us21_n446 ) , .A1( us21_n462 ) , .ZN( us21_n813 ) );
  NAND2_X2 us21_U372 (.A2( us21_n439 ) , .A1( us21_n450 ) , .ZN( us21_n789 ) );
  NAND2_X2 us21_U373 (.A1( us21_n447 ) , .A2( us21_n458 ) , .ZN( us21_n790 ) );
  NAND2_X2 us21_U374 (.A1( us21_n439 ) , .A2( us21_n462 ) , .ZN( us21_n706 ) );
  NAND2_X2 us21_U375 (.A2( us21_n469 ) , .A1( us21_n470 ) , .ZN( us21_n815 ) );
  NAND2_X2 us21_U376 (.A1( us21_n445 ) , .A2( us21_n446 ) , .ZN( us21_n784 ) );
  NOR2_X1 us21_U377 (.A2( sa21_6 ) , .A1( sa21_7 ) , .ZN( us21_n462 ) );
  NOR2_X1 us21_U378 (.A2( sa21_4 ) , .ZN( us21_n447 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U379 (.A2( sa21_5 ) , .ZN( us21_n446 ) , .A1( us21_n845 ) );
  NAND4_X1 us21_U38 (.ZN( sa23_sr_3 ) , .A4( us21_n702 ) , .A3( us21_n703 ) , .A2( us21_n704 ) , .A1( us21_n705 ) );
  NOR2_X1 us21_U380 (.A2( sa21_7 ) , .ZN( us21_n458 ) , .A1( us21_n847 ) );
  NOR2_X1 us21_U381 (.A2( sa21_4 ) , .A1( sa21_5 ) , .ZN( us21_n439 ) );
  NOR2_X1 us21_U382 (.A2( sa21_1 ) , .ZN( us21_n469 ) , .A1( us21_n824 ) );
  NOR2_X1 us21_U383 (.A2( sa21_2 ) , .A1( sa21_3 ) , .ZN( us21_n470 ) );
  NOR2_X1 us21_U384 (.A2( sa21_6 ) , .ZN( us21_n450 ) , .A1( us21_n856 ) );
  NOR2_X1 us21_U385 (.A2( sa21_2 ) , .ZN( us21_n459 ) , .A1( us21_n827 ) );
  NOR2_X1 us21_U386 (.A2( sa21_0 ) , .ZN( us21_n452 ) , .A1( us21_n825 ) );
  NOR2_X1 us21_U387 (.A2( sa21_0 ) , .A1( sa21_1 ) , .ZN( us21_n460 ) );
  NOR2_X1 us21_U388 (.A2( sa21_3 ) , .ZN( us21_n453 ) , .A1( us21_n826 ) );
  INV_X1 us21_U389 (.A( sa21_6 ) , .ZN( us21_n847 ) );
  NOR4_X1 us21_U39 (.A4( us21_n698 ) , .A3( us21_n699 ) , .A2( us21_n700 ) , .A1( us21_n701 ) , .ZN( us21_n702 ) );
  INV_X1 us21_U390 (.A( sa21_3 ) , .ZN( us21_n827 ) );
  INV_X1 us21_U391 (.A( sa21_1 ) , .ZN( us21_n825 ) );
  INV_X1 us21_U392 (.A( sa21_0 ) , .ZN( us21_n824 ) );
  INV_X1 us21_U393 (.A( sa21_2 ) , .ZN( us21_n826 ) );
  INV_X1 us21_U394 (.A( sa21_5 ) , .ZN( us21_n846 ) );
  INV_X1 us21_U395 (.A( sa21_7 ) , .ZN( us21_n856 ) );
  INV_X1 us21_U396 (.A( us21_n784 ) , .ZN( us21_n860 ) );
  AOI21_X1 us21_U397 (.ZN( us21_n498 ) , .A( us21_n695 ) , .B1( us21_n706 ) , .B2( us21_n784 ) );
  INV_X1 us21_U398 (.A( us21_n695 ) , .ZN( us21_n836 ) );
  NOR2_X1 us21_U399 (.A1( us21_n695 ) , .ZN( us21_n768 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U4 (.A1( us21_n447 ) , .A2( us21_n462 ) , .ZN( us21_n722 ) );
  AOI211_X1 us21_U40 (.B( us21_n692 ) , .A( us21_n693 ) , .ZN( us21_n703 ) , .C2( us21_n829 ) , .C1( us21_n849 ) );
  AOI21_X1 us21_U400 (.ZN( us21_n569 ) , .B2( us21_n695 ) , .B1( us21_n804 ) , .A( us21_n810 ) );
  NOR2_X1 us21_U401 (.ZN( us21_n630 ) , .A2( us21_n695 ) , .A1( us21_n722 ) );
  AOI21_X1 us21_U402 (.ZN( us21_n476 ) , .B2( us21_n695 ) , .A( us21_n747 ) , .B1( us21_n777 ) );
  NOR2_X1 us21_U403 (.ZN( us21_n660 ) , .A2( us21_n695 ) , .A1( us21_n727 ) );
  NOR2_X1 us21_U404 (.A2( us21_n695 ) , .A1( us21_n778 ) , .ZN( us21_n818 ) );
  NOR2_X1 us21_U405 (.A2( us21_n695 ) , .ZN( us21_n714 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U406 (.ZN( us21_n564 ) , .A2( us21_n695 ) , .A1( us21_n761 ) );
  NOR2_X1 us21_U407 (.ZN( us21_n592 ) , .A2( us21_n695 ) , .A1( us21_n726 ) );
  AOI21_X1 us21_U408 (.ZN( us21_n550 ) , .B1( us21_n667 ) , .A( us21_n695 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U409 (.ZN( us21_n539 ) , .A2( us21_n695 ) , .A1( us21_n697 ) );
  NOR2_X1 us21_U41 (.ZN( us21_n705 ) , .A2( us21_n774 ) , .A1( us21_n798 ) );
  NOR2_X1 us21_U410 (.ZN( us21_n578 ) , .A2( us21_n695 ) , .A1( us21_n789 ) );
  OAI222_X1 us21_U411 (.B2( us21_n745 ) , .B1( us21_n746 ) , .A2( us21_n747 ) , .ZN( us21_n755 ) , .C2( us21_n803 ) , .C1( us21_n812 ) , .A1( us21_n815 ) );
  OAI222_X1 us21_U412 (.ZN( us21_n503 ) , .C2( us21_n623 ) , .B2( us21_n645 ) , .B1( us21_n745 ) , .A2( us21_n746 ) , .C1( us21_n803 ) , .A1( us21_n804 ) );
  AOI222_X1 us21_U413 (.ZN( us21_n511 ) , .C1( us21_n830 ) , .B2( us21_n835 ) , .A2( us21_n841 ) , .C2( us21_n860 ) , .B1( us21_n861 ) , .A1( us21_n864 ) );
  AOI222_X1 us21_U414 (.ZN( us21_n603 ) , .B2( us21_n669 ) , .B1( us21_n751 ) , .C2( us21_n829 ) , .A1( us21_n831 ) , .A2( us21_n860 ) , .C1( us21_n861 ) );
  AOI221_X1 us21_U415 (.A( us21_n481 ) , .ZN( us21_n486 ) , .B1( us21_n829 ) , .C2( us21_n842 ) , .C1( us21_n850 ) , .B2( us21_n860 ) );
  NOR2_X1 us21_U416 (.ZN( us21_n787 ) , .A2( us21_n860 ) , .A1( us21_n866 ) );
  OAI221_X1 us21_U417 (.A( us21_n781 ) , .C2( us21_n782 ) , .B2( us21_n783 ) , .B1( us21_n784 ) , .ZN( us21_n794 ) , .C1( us21_n811 ) );
  NAND2_X1 us21_U418 (.A1( us21_n727 ) , .A2( us21_n782 ) , .ZN( us21_n809 ) );
  OAI22_X1 us21_U419 (.ZN( us21_n586 ) , .A2( us21_n745 ) , .B2( us21_n760 ) , .A1( us21_n761 ) , .B1( us21_n782 ) );
  NOR2_X1 us21_U42 (.ZN( us21_n802 ) , .A1( us21_n852 ) , .A2( us21_n859 ) );
  OAI221_X1 us21_U420 (.A( us21_n694 ) , .ZN( us21_n701 ) , .C2( us21_n782 ) , .C1( us21_n783 ) , .B1( us21_n784 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U421 (.ZN( us21_n590 ) , .B1( us21_n726 ) , .B2( us21_n782 ) , .A( us21_n788 ) );
  AOI21_X1 us21_U422 (.ZN( us21_n646 ) , .A( us21_n760 ) , .B2( us21_n782 ) , .B1( us21_n790 ) );
  AOI21_X1 us21_U423 (.ZN( us21_n621 ) , .B1( us21_n697 ) , .A( us21_n777 ) , .B2( us21_n782 ) );
  OAI22_X1 us21_U424 (.ZN( us21_n679 ) , .A1( us21_n697 ) , .A2( us21_n728 ) , .B2( us21_n782 ) , .B1( us21_n815 ) );
  OAI21_X1 us21_U425 (.A( us21_n611 ) , .ZN( us21_n614 ) , .B1( us21_n623 ) , .B2( us21_n782 ) );
  NOR2_X1 us21_U426 (.ZN( us21_n608 ) , .A1( us21_n782 ) , .A2( us21_n814 ) );
  OAI222_X1 us21_U427 (.A2( us21_n667 ) , .ZN( us21_n672 ) , .B1( us21_n745 ) , .B2( us21_n782 ) , .C2( us21_n786 ) , .C1( us21_n813 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U428 (.ZN( us21_n649 ) , .A1( us21_n782 ) , .A2( us21_n786 ) );
  NOR2_X1 us21_U429 (.ZN( us21_n598 ) , .A2( us21_n695 ) , .A1( us21_n782 ) );
  NAND4_X1 us21_U43 (.ZN( sa23_sr_2 ) , .A4( us21_n641 ) , .A3( us21_n642 ) , .A2( us21_n643 ) , .A1( us21_n644 ) );
  NOR2_X1 us21_U430 (.ZN( us21_n551 ) , .A2( us21_n742 ) , .A1( us21_n782 ) );
  INV_X1 us21_U431 (.A( us21_n782 ) , .ZN( us21_n859 ) );
  AOI221_X1 us21_U432 (.A( us21_n574 ) , .ZN( us21_n585 ) , .B2( us21_n829 ) , .C2( us21_n841 ) , .B1( us21_n852 ) , .C1( us21_n859 ) );
  AOI21_X1 us21_U433 (.ZN( us21_n574 ) , .B2( us21_n722 ) , .B1( us21_n746 ) , .A( us21_n783 ) );
  INV_X1 us21_U434 (.A( sa21_4 ) , .ZN( us21_n845 ) );
  AOI211_X1 us21_U435 (.A( us21_n635 ) , .ZN( us21_n643 ) , .B( us21_n741 ) , .C2( us21_n837 ) , .C1( us21_n852 ) );
  NAND4_X1 us21_U436 (.A4( us21_n631 ) , .A3( us21_n632 ) , .A2( us21_n633 ) , .A1( us21_n634 ) , .ZN( us21_n741 ) );
  NAND3_X1 us21_U437 (.ZN( sa23_sr_6 ) , .A3( us21_n795 ) , .A2( us21_n796 ) , .A1( us21_n797 ) );
  NAND3_X1 us21_U438 (.ZN( sa23_sr_5 ) , .A3( us21_n756 ) , .A2( us21_n757 ) , .A1( us21_n758 ) );
  NAND3_X1 us21_U439 (.ZN( sa23_sr_4 ) , .A3( us21_n736 ) , .A2( us21_n737 ) , .A1( us21_n738 ) );
  AOI222_X1 us21_U44 (.B2( us21_n636 ) , .ZN( us21_n642 ) , .B1( us21_n839 ) , .A1( us21_n840 ) , .C2( us21_n844 ) , .C1( us21_n861 ) , .A2( us21_n863 ) );
  NAND3_X1 us21_U440 (.A3( us21_n673 ) , .A2( us21_n674 ) , .A1( us21_n675 ) , .ZN( us21_n805 ) );
  NAND3_X1 us21_U441 (.ZN( us21_n636 ) , .A3( us21_n706 ) , .A2( us21_n722 ) , .A1( us21_n790 ) );
  NAND3_X1 us21_U442 (.A3( us21_n616 ) , .A2( us21_n617 ) , .A1( us21_n618 ) , .ZN( us21_n723 ) );
  NAND3_X1 us21_U443 (.A3( us21_n583 ) , .A2( us21_n584 ) , .A1( us21_n585 ) , .ZN( us21_n619 ) );
  NAND3_X1 us21_U444 (.ZN( us21_n563 ) , .A3( us21_n678 ) , .A2( us21_n748 ) , .A1( us21_n783 ) );
  NAND3_X1 us21_U445 (.A3( us21_n521 ) , .A2( us21_n522 ) , .A1( us21_n523 ) , .ZN( us21_n740 ) );
  NAND3_X1 us21_U446 (.A3( us21_n510 ) , .A1( us21_n511 ) , .ZN( us21_n606 ) , .A2( us21_n869 ) );
  NAND3_X1 us21_U447 (.A3( us21_n465 ) , .A2( us21_n466 ) , .A1( us21_n467 ) , .ZN( us21_n775 ) );
  NOR4_X1 us21_U45 (.A4( us21_n637 ) , .A3( us21_n638 ) , .A2( us21_n639 ) , .A1( us21_n640 ) , .ZN( us21_n641 ) );
  NOR3_X1 us21_U46 (.A2( us21_n605 ) , .A1( us21_n606 ) , .ZN( us21_n644 ) , .A3( us21_n720 ) );
  NAND4_X1 us21_U47 (.ZN( sa23_sr_0 ) , .A4( us21_n499 ) , .A3( us21_n500 ) , .A2( us21_n501 ) , .A1( us21_n502 ) );
  NOR4_X1 us21_U48 (.A4( us21_n496 ) , .A3( us21_n497 ) , .A2( us21_n498 ) , .ZN( us21_n499 ) , .A1( us21_n525 ) );
  AOI221_X1 us21_U49 (.A( us21_n495 ) , .ZN( us21_n500 ) , .B2( us21_n841 ) , .C1( us21_n844 ) , .C2( us21_n858 ) , .B1( us21_n860 ) );
  NAND2_X1 us21_U5 (.A1( us21_n445 ) , .A2( us21_n447 ) , .ZN( us21_n803 ) );
  AOI211_X1 us21_U50 (.A( us21_n494 ) , .ZN( us21_n501 ) , .B( us21_n800 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NAND4_X1 us21_U51 (.ZN( sa23_sr_1 ) , .A4( us21_n593 ) , .A3( us21_n594 ) , .A2( us21_n595 ) , .A1( us21_n596 ) );
  AOI211_X1 us21_U52 (.B( us21_n587 ) , .A( us21_n588 ) , .ZN( us21_n594 ) , .C2( us21_n809 ) , .C1( us21_n831 ) );
  NOR4_X1 us21_U53 (.A4( us21_n589 ) , .A3( us21_n590 ) , .A2( us21_n591 ) , .A1( us21_n592 ) , .ZN( us21_n593 ) );
  AOI211_X1 us21_U54 (.A( us21_n586 ) , .ZN( us21_n595 ) , .B( us21_n619 ) , .C1( us21_n843 ) , .C2( us21_n853 ) );
  NAND4_X1 us21_U55 (.A4( us21_n601 ) , .A3( us21_n602 ) , .A2( us21_n603 ) , .A1( us21_n604 ) , .ZN( us21_n720 ) );
  NOR3_X1 us21_U56 (.A1( us21_n597 ) , .ZN( us21_n602 ) , .A3( us21_n661 ) , .A2( us21_n768 ) );
  NOR4_X1 us21_U57 (.A3( us21_n598 ) , .A2( us21_n599 ) , .A1( us21_n600 ) , .ZN( us21_n601 ) , .A4( us21_n653 ) );
  AOI222_X1 us21_U58 (.ZN( us21_n604 ) , .A1( us21_n828 ) , .C2( us21_n835 ) , .B1( us21_n840 ) , .A2( us21_n854 ) , .B2( us21_n859 ) , .C1( us21_n866 ) );
  AOI222_X1 us21_U59 (.ZN( us21_n467 ) , .B1( us21_n830 ) , .A1( us21_n837 ) , .C1( us21_n840 ) , .C2( us21_n849 ) , .A2( us21_n853 ) , .B2( us21_n863 ) );
  NOR3_X1 us21_U6 (.ZN( us21_n596 ) , .A1( us21_n606 ) , .A3( us21_n721 ) , .A2( us21_n740 ) );
  NOR4_X1 us21_U60 (.A1( us21_n464 ) , .ZN( us21_n465 ) , .A4( us21_n540 ) , .A2( us21_n552 ) , .A3( us21_n612 ) );
  AOI221_X1 us21_U61 (.ZN( us21_n466 ) , .C2( us21_n712 ) , .B2( us21_n829 ) , .C1( us21_n843 ) , .B1( us21_n858 ) , .A( us21_n862 ) );
  NAND4_X1 us21_U62 (.A4( us21_n483 ) , .A3( us21_n484 ) , .A2( us21_n485 ) , .A1( us21_n486 ) , .ZN( us21_n776 ) );
  NOR4_X1 us21_U63 (.ZN( us21_n484 ) , .A1( us21_n505 ) , .A2( us21_n517 ) , .A4( us21_n544 ) , .A3( us21_n609 ) );
  NOR4_X1 us21_U64 (.A4( us21_n482 ) , .ZN( us21_n485 ) , .A1( us21_n564 ) , .A2( us21_n579 ) , .A3( us21_n600 ) );
  NOR4_X1 us21_U65 (.ZN( us21_n483 ) , .A2( us21_n531 ) , .A1( us21_n556 ) , .A3( us21_n629 ) , .A4( us21_n716 ) );
  AOI211_X1 us21_U66 (.B( us21_n621 ) , .A( us21_n622 ) , .ZN( us21_n633 ) , .C2( us21_n834 ) , .C1( us21_n861 ) );
  NOR4_X1 us21_U67 (.A4( us21_n627 ) , .A3( us21_n628 ) , .A2( us21_n629 ) , .A1( us21_n630 ) , .ZN( us21_n631 ) );
  NOR4_X1 us21_U68 (.A4( us21_n624 ) , .A3( us21_n625 ) , .A2( us21_n626 ) , .ZN( us21_n632 ) , .A1( us21_n662 ) );
  NOR4_X1 us21_U69 (.A4( us21_n512 ) , .A3( us21_n513 ) , .A2( us21_n514 ) , .A1( us21_n515 ) , .ZN( us21_n522 ) );
  NOR3_X1 us21_U7 (.A3( us21_n798 ) , .A2( us21_n799 ) , .A1( us21_n800 ) , .ZN( us21_n823 ) );
  AOI222_X1 us21_U70 (.ZN( us21_n523 ) , .A1( us21_n832 ) , .B2( us21_n835 ) , .C1( us21_n842 ) , .C2( us21_n848 ) , .A2( us21_n850 ) , .B1( us21_n864 ) );
  NOR4_X1 us21_U71 (.A3( us21_n519 ) , .A1( us21_n520 ) , .ZN( us21_n521 ) , .A2( us21_n671 ) , .A4( us21_n767 ) );
  NAND4_X1 us21_U72 (.A4( us21_n655 ) , .A3( us21_n656 ) , .A2( us21_n657 ) , .A1( us21_n658 ) , .ZN( us21_n798 ) );
  NOR3_X1 us21_U73 (.A3( us21_n646 ) , .A2( us21_n647 ) , .A1( us21_n648 ) , .ZN( us21_n657 ) );
  NOR3_X1 us21_U74 (.A3( us21_n649 ) , .A2( us21_n650 ) , .A1( us21_n651 ) , .ZN( us21_n656 ) );
  NOR3_X1 us21_U75 (.A3( us21_n652 ) , .A2( us21_n653 ) , .A1( us21_n654 ) , .ZN( us21_n655 ) );
  NAND4_X1 us21_U76 (.A4( us21_n558 ) , .A3( us21_n559 ) , .A2( us21_n560 ) , .A1( us21_n561 ) , .ZN( us21_n605 ) );
  NOR4_X1 us21_U77 (.A4( us21_n550 ) , .A3( us21_n551 ) , .A2( us21_n552 ) , .A1( us21_n553 ) , .ZN( us21_n560 ) );
  NOR4_X1 us21_U78 (.A4( us21_n554 ) , .A3( us21_n555 ) , .A2( us21_n556 ) , .A1( us21_n557 ) , .ZN( us21_n558 ) );
  NOR4_X1 us21_U79 (.ZN( us21_n559 ) , .A1( us21_n651 ) , .A3( us21_n659 ) , .A4( us21_n683 ) , .A2( us21_n766 ) );
  NOR3_X1 us21_U8 (.ZN( us21_n502 ) , .A2( us21_n677 ) , .A3( us21_n775 ) , .A1( us21_n874 ) );
  NAND4_X1 us21_U80 (.A4( us21_n770 ) , .A3( us21_n771 ) , .A2( us21_n772 ) , .A1( us21_n773 ) , .ZN( us21_n799 ) );
  NOR3_X1 us21_U81 (.A3( us21_n763 ) , .A2( us21_n764 ) , .A1( us21_n765 ) , .ZN( us21_n771 ) );
  NOR4_X1 us21_U82 (.A4( us21_n766 ) , .A3( us21_n767 ) , .A2( us21_n768 ) , .A1( us21_n769 ) , .ZN( us21_n770 ) );
  AOI222_X1 us21_U83 (.ZN( us21_n773 ) , .A1( us21_n828 ) , .C1( us21_n832 ) , .B2( us21_n839 ) , .A2( us21_n848 ) , .B1( us21_n859 ) , .C2( us21_n871 ) );
  NOR4_X1 us21_U84 (.A4( us21_n507 ) , .A2( us21_n508 ) , .A1( us21_n509 ) , .ZN( us21_n510 ) , .A3( us21_n668 ) );
  INV_X1 us21_U85 (.A( us21_n503 ) , .ZN( us21_n869 ) );
  NOR4_X1 us21_U86 (.A4( us21_n659 ) , .A3( us21_n660 ) , .A2( us21_n661 ) , .A1( us21_n662 ) , .ZN( us21_n675 ) );
  NOR4_X1 us21_U87 (.A4( us21_n663 ) , .A3( us21_n664 ) , .A2( us21_n665 ) , .A1( us21_n666 ) , .ZN( us21_n674 ) );
  NOR4_X1 us21_U88 (.A3( us21_n671 ) , .A1( us21_n672 ) , .ZN( us21_n673 ) , .A4( us21_n713 ) , .A2( us21_n857 ) );
  NOR2_X1 us21_U89 (.ZN( us21_n623 ) , .A2( us21_n834 ) , .A1( us21_n837 ) );
  INV_X1 us21_U9 (.A( us21_n704 ) , .ZN( us21_n874 ) );
  NOR2_X1 us21_U90 (.ZN( us21_n759 ) , .A1( us21_n831 ) , .A2( us21_n832 ) );
  NAND4_X1 us21_U91 (.A4( us21_n454 ) , .A3( us21_n455 ) , .A2( us21_n456 ) , .A1( us21_n457 ) , .ZN( us21_n677 ) );
  NOR3_X1 us21_U92 (.ZN( us21_n455 ) , .A3( us21_n528 ) , .A1( us21_n553 ) , .A2( us21_n568 ) );
  AOI221_X1 us21_U93 (.A( us21_n448 ) , .ZN( us21_n457 ) , .C2( us21_n751 ) , .B1( us21_n830 ) , .C1( us21_n840 ) , .B2( us21_n859 ) );
  NOR4_X1 us21_U94 (.ZN( us21_n456 ) , .A2( us21_n507 ) , .A1( us21_n597 ) , .A4( us21_n626 ) , .A3( us21_n709 ) );
  NAND4_X1 us21_U95 (.ZN( sa23_sr_7 ) , .A4( us21_n820 ) , .A3( us21_n821 ) , .A2( us21_n822 ) , .A1( us21_n823 ) );
  NOR4_X1 us21_U96 (.A4( us21_n816 ) , .A3( us21_n817 ) , .A2( us21_n818 ) , .A1( us21_n819 ) , .ZN( us21_n820 ) );
  AOI222_X1 us21_U97 (.C2( us21_n807 ) , .B2( us21_n808 ) , .A2( us21_n809 ) , .ZN( us21_n821 ) , .C1( us21_n830 ) , .A1( us21_n837 ) , .B1( us21_n851 ) );
  AOI211_X1 us21_U98 (.B( us21_n805 ) , .A( us21_n806 ) , .ZN( us21_n822 ) , .C1( us21_n840 ) , .C2( us21_n848 ) );
  NAND4_X1 us21_U99 (.A4( us21_n533 ) , .A3( us21_n534 ) , .A2( us21_n535 ) , .A1( us21_n536 ) , .ZN( us21_n620 ) );
endmodule

