module aes_aes_die_5 ( sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7 );
  input sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, sa32_7;
  output sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7;
  wire us32_n438, us32_n439, us32_n440, us32_n441, us32_n442, us32_n443, us32_n444, us32_n445, us32_n446, 
       us32_n447, us32_n448, us32_n449, us32_n450, us32_n451, us32_n452, us32_n453, us32_n454, us32_n455, 
       us32_n456, us32_n457, us32_n458, us32_n459, us32_n460, us32_n461, us32_n462, us32_n463, us32_n464, 
       us32_n465, us32_n466, us32_n467, us32_n468, us32_n469, us32_n470, us32_n471, us32_n472, us32_n473, 
       us32_n474, us32_n475, us32_n476, us32_n477, us32_n478, us32_n479, us32_n480, us32_n481, us32_n482, 
       us32_n483, us32_n484, us32_n485, us32_n486, us32_n487, us32_n488, us32_n489, us32_n490, us32_n491, 
       us32_n492, us32_n493, us32_n494, us32_n495, us32_n496, us32_n497, us32_n498, us32_n499, us32_n500, 
       us32_n501, us32_n502, us32_n503, us32_n504, us32_n505, us32_n506, us32_n507, us32_n508, us32_n509, 
       us32_n510, us32_n511, us32_n512, us32_n513, us32_n514, us32_n515, us32_n516, us32_n517, us32_n518, 
       us32_n519, us32_n520, us32_n521, us32_n522, us32_n523, us32_n524, us32_n525, us32_n526, us32_n527, 
       us32_n528, us32_n529, us32_n530, us32_n531, us32_n532, us32_n533, us32_n534, us32_n535, us32_n536, 
       us32_n537, us32_n538, us32_n539, us32_n540, us32_n541, us32_n542, us32_n543, us32_n544, us32_n545, 
       us32_n546, us32_n547, us32_n548, us32_n549, us32_n550, us32_n551, us32_n552, us32_n553, us32_n554, 
       us32_n555, us32_n556, us32_n557, us32_n558, us32_n559, us32_n560, us32_n561, us32_n562, us32_n563, 
       us32_n564, us32_n565, us32_n566, us32_n567, us32_n568, us32_n569, us32_n570, us32_n571, us32_n572, 
       us32_n573, us32_n574, us32_n575, us32_n576, us32_n577, us32_n578, us32_n579, us32_n580, us32_n581, 
       us32_n582, us32_n583, us32_n584, us32_n585, us32_n586, us32_n587, us32_n588, us32_n589, us32_n590, 
       us32_n591, us32_n592, us32_n593, us32_n594, us32_n595, us32_n596, us32_n597, us32_n598, us32_n599, 
       us32_n600, us32_n601, us32_n602, us32_n603, us32_n604, us32_n605, us32_n606, us32_n607, us32_n608, 
       us32_n609, us32_n610, us32_n611, us32_n612, us32_n613, us32_n614, us32_n615, us32_n616, us32_n617, 
       us32_n618, us32_n619, us32_n620, us32_n621, us32_n622, us32_n623, us32_n624, us32_n625, us32_n626, 
       us32_n627, us32_n628, us32_n629, us32_n630, us32_n631, us32_n632, us32_n633, us32_n634, us32_n635, 
       us32_n636, us32_n637, us32_n638, us32_n639, us32_n640, us32_n641, us32_n642, us32_n643, us32_n644, 
       us32_n645, us32_n646, us32_n647, us32_n648, us32_n649, us32_n650, us32_n651, us32_n652, us32_n653, 
       us32_n654, us32_n655, us32_n656, us32_n657, us32_n658, us32_n659, us32_n660, us32_n661, us32_n662, 
       us32_n663, us32_n664, us32_n665, us32_n666, us32_n667, us32_n668, us32_n669, us32_n670, us32_n671, 
       us32_n672, us32_n673, us32_n674, us32_n675, us32_n676, us32_n677, us32_n678, us32_n679, us32_n680, 
       us32_n681, us32_n682, us32_n683, us32_n684, us32_n685, us32_n686, us32_n687, us32_n688, us32_n689, 
       us32_n690, us32_n691, us32_n692, us32_n693, us32_n694, us32_n695, us32_n696, us32_n697, us32_n698, 
       us32_n699, us32_n700, us32_n701, us32_n702, us32_n703, us32_n704, us32_n705, us32_n706, us32_n707, 
       us32_n708, us32_n709, us32_n710, us32_n711, us32_n712, us32_n713, us32_n714, us32_n715, us32_n716, 
       us32_n717, us32_n718, us32_n719, us32_n720, us32_n721, us32_n722, us32_n723, us32_n724, us32_n725, 
       us32_n726, us32_n727, us32_n728, us32_n729, us32_n730, us32_n731, us32_n732, us32_n733, us32_n734, 
       us32_n735, us32_n736, us32_n737, us32_n738, us32_n739, us32_n740, us32_n741, us32_n742, us32_n743, 
       us32_n744, us32_n745, us32_n746, us32_n747, us32_n748, us32_n749, us32_n750, us32_n751, us32_n752, 
       us32_n753, us32_n754, us32_n755, us32_n756, us32_n757, us32_n758, us32_n759, us32_n760, us32_n761, 
       us32_n762, us32_n763, us32_n764, us32_n765, us32_n766, us32_n767, us32_n768, us32_n769, us32_n770, 
       us32_n771, us32_n772, us32_n773, us32_n774, us32_n775, us32_n776, us32_n777, us32_n778, us32_n779, 
       us32_n780, us32_n781, us32_n782, us32_n783, us32_n784, us32_n785, us32_n786, us32_n787, us32_n788, 
       us32_n789, us32_n790, us32_n791, us32_n792, us32_n793, us32_n794, us32_n795, us32_n796, us32_n797, 
       us32_n798, us32_n799, us32_n800, us32_n801, us32_n802, us32_n803, us32_n804, us32_n805, us32_n806, 
       us32_n807, us32_n808, us32_n809, us32_n810, us32_n811, us32_n812, us32_n813, us32_n814, us32_n815, 
       us32_n816, us32_n817, us32_n818, us32_n819, us32_n820, us32_n821, us32_n822, us32_n823, us32_n824, 
       us32_n825, us32_n826, us32_n827, us32_n828, us32_n829, us32_n830, us32_n831, us32_n832, us32_n833, 
       us32_n834, us32_n835, us32_n836, us32_n837, us32_n838, us32_n839, us32_n840, us32_n841, us32_n842, 
       us32_n843, us32_n844, us32_n845, us32_n846, us32_n847, us32_n848, us32_n849, us32_n850, us32_n851, 
       us32_n852, us32_n853, us32_n854, us32_n855, us32_n856, us32_n857, us32_n858, us32_n859, us32_n860, 
       us32_n861, us32_n862, us32_n863, us32_n864, us32_n865, us32_n866, us32_n867, us32_n868, us32_n869, 
       us32_n870, us32_n871, us32_n872, us32_n873, us32_n874, us32_n875,  us32_n876;
  NOR2_X1 us32_U10 (.A1( us32_n678 ) , .ZN( us32_n693 ) , .A2( us32_n807 ) );
  AOI211_X1 us32_U100 (.B( us32_n477 ) , .A( us32_n478 ) , .ZN( us32_n482 ) , .C2( us32_n833 ) , .C1( us32_n861 ) );
  NOR4_X1 us32_U101 (.ZN( us32_n481 ) , .A3( us32_n532 ) , .A4( us32_n545 ) , .A2( us32_n567 ) , .A1( us32_n717 ) );
  NAND4_X1 us32_U102 (.A4( us32_n548 ) , .A3( us32_n549 ) , .A2( us32_n550 ) , .A1( us32_n551 ) , .ZN( us32_n745 ) );
  NOR3_X1 us32_U103 (.ZN( us32_n549 ) , .A2( us32_n651 ) , .A1( us32_n667 ) , .A3( us32_n771 ) );
  AOI211_X1 us32_U104 (.B( us32_n539 ) , .A( us32_n540 ) , .ZN( us32_n551 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NOR4_X1 us32_U105 (.A4( us32_n541 ) , .A3( us32_n542 ) , .A2( us32_n543 ) , .ZN( us32_n550 ) , .A1( us32_n688 ) );
  NOR4_X1 us32_U106 (.ZN( us32_n620 ) , .A1( us32_n656 ) , .A3( us32_n666 ) , .A4( us32_n682 ) , .A2( us32_n766 ) );
  NOR4_X1 us32_U107 (.A4( us32_n609 ) , .A3( us32_n610 ) , .A2( us32_n611 ) , .A1( us32_n612 ) , .ZN( us32_n619 ) );
  NOR4_X1 us32_U108 (.A4( us32_n614 ) , .A3( us32_n615 ) , .A2( us32_n616 ) , .A1( us32_n617 ) , .ZN( us32_n618 ) );
  NOR2_X1 us32_U109 (.ZN( us32_n686 ) , .A1( us32_n831 ) , .A2( us32_n832 ) );
  NOR3_X1 us32_U11 (.ZN( us32_n504 ) , .A2( us32_n679 ) , .A3( us32_n777 ) , .A1( us32_n876 ) );
  NAND4_X1 us32_U110 (.A4( us32_n485 ) , .A3( us32_n486 ) , .A2( us32_n487 ) , .A1( us32_n488 ) , .ZN( us32_n778 ) );
  NOR4_X1 us32_U111 (.A4( us32_n484 ) , .ZN( us32_n487 ) , .A1( us32_n566 ) , .A2( us32_n581 ) , .A3( us32_n602 ) );
  NOR4_X1 us32_U112 (.ZN( us32_n486 ) , .A1( us32_n507 ) , .A2( us32_n519 ) , .A4( us32_n546 ) , .A3( us32_n611 ) );
  NOR4_X1 us32_U113 (.ZN( us32_n485 ) , .A2( us32_n533 ) , .A1( us32_n558 ) , .A3( us32_n631 ) , .A4( us32_n718 ) );
  NAND4_X1 us32_U114 (.A4( us32_n691 ) , .A3( us32_n692 ) , .A1( us32_n693 ) , .ZN( us32_n776 ) , .A2( us32_n872 ) );
  AOI221_X1 us32_U115 (.A( us32_n681 ) , .ZN( us32_n692 ) , .B2( us32_n840 ) , .C1( us32_n842 ) , .C2( us32_n862 ) , .B1( us32_n865 ) );
  INV_X1 us32_U116 (.A( us32_n679 ) , .ZN( us32_n872 ) );
  NOR4_X1 us32_U117 (.A4( us32_n687 ) , .A3( us32_n688 ) , .A2( us32_n689 ) , .A1( us32_n690 ) , .ZN( us32_n691 ) );
  NAND4_X1 us32_U118 (.A4( us32_n473 ) , .A3( us32_n474 ) , .A2( us32_n475 ) , .A1( us32_n476 ) , .ZN( us32_n678 ) );
  NOR4_X1 us32_U119 (.ZN( us32_n475 ) , .A1( us32_n531 ) , .A3( us32_n568 ) , .A4( us32_n600 ) , .A2( us32_n642 ) );
  INV_X1 us32_U12 (.A( us32_n706 ) , .ZN( us32_n876 ) );
  NOR4_X1 us32_U120 (.A4( us32_n470 ) , .ZN( us32_n476 ) , .A3( us32_n556 ) , .A1( us32_n735 ) , .A2( us32_n755 ) );
  NOR4_X1 us32_U121 (.ZN( us32_n473 ) , .A2( us32_n521 ) , .A4( us32_n594 ) , .A1( us32_n609 ) , .A3( us32_n629 ) );
  NAND4_X1 us32_U122 (.A4( us32_n719 ) , .A3( us32_n720 ) , .A2( us32_n721 ) , .ZN( us32_n741 ) , .A1( us32_n857 ) );
  INV_X1 us32_U123 (.A( us32_n709 ) , .ZN( us32_n857 ) );
  AOI221_X1 us32_U124 (.A( us32_n710 ) , .ZN( us32_n721 ) , .C2( us32_n844 ) , .B2( us32_n845 ) , .C1( us32_n861 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U125 (.A4( us32_n715 ) , .A3( us32_n716 ) , .A2( us32_n717 ) , .A1( us32_n718 ) , .ZN( us32_n719 ) );
  NOR2_X1 us32_U126 (.ZN( us32_n733 ) , .A2( us32_n832 ) , .A1( us32_n845 ) );
  NOR2_X1 us32_U127 (.ZN( us32_n789 ) , .A2( us32_n862 ) , .A1( us32_n868 ) );
  NAND4_X1 us32_U128 (.A4( us32_n573 ) , .A3( us32_n574 ) , .A1( us32_n575 ) , .ZN( us32_n723 ) , .A2( us32_n874 ) );
  AOI221_X1 us32_U129 (.A( us32_n564 ) , .C2( us32_n565 ) , .ZN( us32_n574 ) , .B2( us32_n845 ) , .B1( us32_n852 ) , .C1( us32_n853 ) );
  INV_X1 us32_U13 (.A( us32_n607 ) , .ZN( us32_n874 ) );
  NOR4_X1 us32_U130 (.A4( us32_n569 ) , .A3( us32_n570 ) , .A2( us32_n571 ) , .A1( us32_n572 ) , .ZN( us32_n573 ) );
  NOR2_X1 us32_U131 (.ZN( us32_n575 ) , .A1( us32_n622 ) , .A2( us32_n745 ) );
  NOR2_X1 us32_U132 (.ZN( us32_n748 ) , .A1( us32_n861 ) , .A2( us32_n862 ) );
  NAND4_X1 us32_U133 (.A4( us32_n633 ) , .A3( us32_n634 ) , .A2( us32_n635 ) , .A1( us32_n636 ) , .ZN( us32_n743 ) );
  AOI211_X1 us32_U134 (.B( us32_n623 ) , .A( us32_n624 ) , .ZN( us32_n635 ) , .C2( us32_n836 ) , .C1( us32_n863 ) );
  NOR4_X1 us32_U135 (.A4( us32_n629 ) , .A3( us32_n630 ) , .A2( us32_n631 ) , .A1( us32_n632 ) , .ZN( us32_n633 ) );
  NOR4_X1 us32_U136 (.A4( us32_n626 ) , .A3( us32_n627 ) , .A2( us32_n628 ) , .ZN( us32_n634 ) , .A1( us32_n664 ) );
  NAND4_X1 us32_U137 (.A4( us32_n493 ) , .A3( us32_n494 ) , .A1( us32_n495 ) , .ZN( us32_n802 ) , .A2( us32_n867 ) );
  AOI221_X1 us32_U138 (.A( us32_n489 ) , .ZN( us32_n494 ) , .B2( us32_n836 ) , .C2( us32_n841 ) , .C1( us32_n851 ) , .B1( us32_n860 ) );
  INV_X1 us32_U139 (.A( us32_n778 ) , .ZN( us32_n867 ) );
  INV_X1 us32_U14 (.A( us32_n680 ) , .ZN( us32_n840 ) );
  NOR4_X1 us32_U140 (.A2( us32_n491 ) , .A1( us32_n492 ) , .ZN( us32_n493 ) , .A3( us32_n580 ) , .A4( us32_n612 ) );
  NOR4_X1 us32_U141 (.A4( us32_n734 ) , .A3( us32_n735 ) , .A2( us32_n736 ) , .A1( us32_n737 ) , .ZN( us32_n738 ) );
  AOI211_X1 us32_U142 (.B( us32_n725 ) , .A( us32_n726 ) , .ZN( us32_n739 ) , .C1( us32_n843 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U143 (.A3( us32_n722 ) , .A1( us32_n723 ) , .ZN( us32_n740 ) , .A2( us32_n741 ) );
  NOR2_X1 us32_U144 (.ZN( us32_n647 ) , .A1( us32_n854 ) , .A2( us32_n868 ) );
  INV_X1 us32_U145 (.A( us32_n762 ) , .ZN( us32_n830 ) );
  INV_X1 us32_U146 (.A( us32_n754 ) , .ZN( us32_n869 ) );
  OAI21_X1 us32_U147 (.B1( us32_n753 ) , .ZN( us32_n754 ) , .A( us32_n845 ) , .B2( us32_n868 ) );
  INV_X1 us32_U148 (.A( us32_n697 ) , .ZN( us32_n838 ) );
  OR4_X1 us32_U149 (.ZN( us32_n492 ) , .A4( us32_n534 ) , .A2( us32_n547 ) , .A1( us32_n559 ) , .A3( us32_n632 ) );
  NOR4_X1 us32_U15 (.A4( us32_n445 ) , .A3( us32_n446 ) , .A2( us32_n516 ) , .A1( us32_n541 ) , .ZN( us32_n706 ) );
  OR4_X1 us32_U150 (.A4( us32_n566 ) , .A3( us32_n567 ) , .A2( us32_n568 ) , .ZN( us32_n572 ) , .A1( us32_n665 ) );
  OR4_X1 us32_U151 (.A4( us32_n682 ) , .A3( us32_n683 ) , .A2( us32_n684 ) , .A1( us32_n685 ) , .ZN( us32_n690 ) );
  OR4_X1 us32_U152 (.ZN( us32_n466 ) , .A4( us32_n518 ) , .A3( us32_n529 ) , .A2( us32_n578 ) , .A1( us32_n712 ) );
  OR4_X1 us32_U153 (.A4( us32_n518 ) , .A2( us32_n519 ) , .A1( us32_n520 ) , .ZN( us32_n522 ) , .A3( us32_n821 ) );
  OR4_X1 us32_U154 (.A4( us32_n580 ) , .A3( us32_n581 ) , .A2( us32_n582 ) , .A1( us32_n583 ) , .ZN( us32_n584 ) );
  NAND2_X1 us32_U155 (.ZN( us32_n613 ) , .A2( us32_n837 ) , .A1( us32_n873 ) );
  OR3_X1 us32_U156 (.A3( us32_n506 ) , .A2( us32_n507 ) , .A1( us32_n508 ) , .ZN( us32_n511 ) );
  INV_X1 us32_U157 (.A( us32_n672 ) , .ZN( us32_n859 ) );
  AOI21_X1 us32_U158 (.A( us32_n670 ) , .B1( us32_n671 ) , .ZN( us32_n672 ) , .B2( us32_n856 ) );
  INV_X1 us32_U159 (.A( us32_n463 ) , .ZN( us32_n864 ) );
  OR3_X1 us32_U16 (.ZN( us32_n446 ) , .A1( us32_n528 ) , .A3( us32_n577 ) , .A2( us32_n875 ) );
  OAI21_X1 us32_U160 (.ZN( us32_n463 ) , .B1( us32_n809 ) , .A( us32_n834 ) , .B2( us32_n851 ) );
  OAI222_X1 us32_U161 (.B2( us32_n708 ) , .ZN( us32_n709 ) , .C2( us32_n724 ) , .B1( us32_n747 ) , .A1( us32_n806 ) , .C1( us32_n814 ) , .A2( us32_n815 ) );
  NAND2_X1 us32_U162 (.A1( us32_n447 ) , .A2( us32_n465 ) , .ZN( us32_n749 ) );
  AOI22_X1 us32_U163 (.A2( us32_n782 ) , .ZN( us32_n783 ) , .B2( us32_n831 ) , .A1( us32_n834 ) , .B1( us32_n863 ) );
  AOI22_X1 us32_U164 (.ZN( us32_n696 ) , .A1( us32_n830 ) , .B2( us32_n843 ) , .A2( us32_n865 ) , .B1( us32_n868 ) );
  INV_X1 us32_U165 (.A( us32_n730 ) , .ZN( us32_n839 ) );
  AOI221_X1 us32_U166 (.A( us32_n483 ) , .ZN( us32_n488 ) , .B1( us32_n831 ) , .C2( us32_n844 ) , .C1( us32_n852 ) , .B2( us32_n862 ) );
  OAI22_X1 us32_U167 (.ZN( us32_n483 ) , .A1( us32_n708 ) , .B2( us32_n785 ) , .A2( us32_n806 ) , .B1( us32_n812 ) );
  INV_X1 us32_U168 (.A( us32_n790 ) , .ZN( us32_n832 ) );
  OAI221_X1 us32_U169 (.A( us32_n727 ) , .C2( us32_n728 ) , .B2( us32_n729 ) , .B1( us32_n730 ) , .ZN( us32_n737 ) , .C1( us32_n817 ) );
  OR4_X1 us32_U17 (.A4( us32_n442 ) , .A2( us32_n443 ) , .A1( us32_n444 ) , .ZN( us32_n445 ) , .A3( us32_n553 ) );
  AOI22_X1 us32_U170 (.ZN( us32_n727 ) , .B1( us32_n832 ) , .A2( us32_n838 ) , .A1( us32_n863 ) , .B2( us32_n866 ) );
  NAND2_X1 us32_U171 (.A1( us32_n451 ) , .A2( us32_n453 ) , .ZN( us32_n762 ) );
  INV_X1 us32_U172 (.A( us32_n786 ) , .ZN( us32_n862 ) );
  OAI22_X1 us32_U173 (.ZN( us32_n710 ) , .A2( us32_n728 ) , .B2( us32_n729 ) , .A1( us32_n744 ) , .B1( us32_n813 ) );
  INV_X1 us32_U174 (.A( us32_n816 ) , .ZN( us32_n831 ) );
  OAI22_X1 us32_U175 (.ZN( us32_n489 ) , .A1( us32_n724 ) , .B2( us32_n728 ) , .B1( us32_n730 ) , .A2( us32_n779 ) );
  OAI22_X1 us32_U176 (.ZN( us32_n624 ) , .B1( us32_n669 ) , .B2( us32_n747 ) , .A1( us32_n815 ) , .A2( us32_n816 ) );
  INV_X1 us32_U177 (.A( us32_n788 ) , .ZN( us32_n845 ) );
  OAI22_X1 us32_U178 (.A1( us32_n724 ) , .ZN( us32_n726 ) , .B2( us32_n750 ) , .B1( us32_n812 ) , .A2( us32_n816 ) );
  INV_X1 us32_U179 (.A( us32_n744 ) , .ZN( us32_n837 ) );
  INV_X1 us32_U18 (.A( us32_n613 ) , .ZN( us32_n875 ) );
  OAI22_X1 us32_U180 (.B2( us32_n779 ) , .B1( us32_n780 ) , .ZN( us32_n781 ) , .A2( us32_n814 ) , .A1( us32_n815 ) );
  INV_X1 us32_U181 (.A( us32_n814 ) , .ZN( us32_n833 ) );
  INV_X1 us32_U182 (.A( us32_n669 ) , .ZN( us32_n865 ) );
  OAI22_X1 us32_U183 (.B2( us32_n744 ) , .ZN( us32_n746 ) , .A2( us32_n762 ) , .B1( us32_n780 ) , .A1( us32_n792 ) );
  OAI22_X1 us32_U184 (.ZN( us32_n496 ) , .A2( us32_n744 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n806 ) );
  AOI211_X1 us32_U185 (.A( us32_n637 ) , .ZN( us32_n645 ) , .B( us32_n743 ) , .C2( us32_n839 ) , .C1( us32_n854 ) );
  OAI22_X1 us32_U186 (.ZN( us32_n637 ) , .A1( us32_n699 ) , .B2( us32_n728 ) , .A2( us32_n762 ) , .B1( us32_n816 ) );
  INV_X1 us32_U187 (.A( us32_n750 ) , .ZN( us32_n842 ) );
  OAI22_X1 us32_U188 (.B1( us32_n490 ) , .ZN( us32_n491 ) , .A1( us32_n686 ) , .A2( us32_n763 ) , .B2( us32_n817 ) );
  NOR3_X1 us32_U189 (.ZN( us32_n490 ) , .A1( us32_n782 ) , .A2( us32_n850 ) , .A3( us32_n863 ) );
  INV_X1 us32_U19 (.A( us32_n749 ) , .ZN( us32_n863 ) );
  OAI22_X1 us32_U190 (.ZN( us32_n695 ) , .A2( us32_n730 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U191 (.ZN( us32_n666 ) , .A1( us32_n728 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U192 (.ZN( us32_n594 ) , .A2( us32_n697 ) , .A1( us32_n728 ) );
  NOR2_X1 us32_U193 (.ZN( us32_n570 ) , .A1( us32_n728 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U194 (.ZN( us32_n654 ) , .A1( us32_n728 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U195 (.ZN( us32_n546 ) , .A2( us32_n780 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U196 (.ZN( us32_n532 ) , .A2( us32_n749 ) , .A1( us32_n750 ) );
  NOR2_X1 us32_U197 (.ZN( us32_n577 ) , .A2( us32_n699 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U198 (.ZN( us32_n615 ) , .A1( us32_n785 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U199 (.ZN( us32_n629 ) , .A2( us32_n728 ) , .A1( us32_n785 ) );
  AOI222_X1 us32_U20 (.ZN( us32_n605 ) , .B2( us32_n671 ) , .B1( us32_n753 ) , .C2( us32_n831 ) , .A1( us32_n833 ) , .A2( us32_n862 ) , .C1( us32_n863 ) );
  NOR2_X1 us32_U200 (.ZN( us32_n718 ) , .A2( us32_n724 ) , .A1( us32_n744 ) );
  NOR2_X1 us32_U201 (.ZN( us32_n628 ) , .A2( us32_n669 ) , .A1( us32_n785 ) );
  INV_X1 us32_U202 (.A( us32_n728 ) , .ZN( us32_n852 ) );
  NOR2_X1 us32_U203 (.A2( us32_n744 ) , .ZN( us32_n769 ) , .A1( us32_n812 ) );
  NOR2_X1 us32_U204 (.ZN( us32_n531 ) , .A2( us32_n780 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U205 (.A2( us32_n708 ) , .A1( us32_n750 ) , .ZN( us32_n771 ) );
  NOR2_X1 us32_U206 (.ZN( us32_n599 ) , .A2( us32_n791 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U207 (.ZN( us32_n611 ) , .A2( us32_n780 ) , .A1( us32_n806 ) );
  NOR2_X1 us32_U208 (.ZN( us32_n652 ) , .A1( us32_n669 ) , .A2( us32_n814 ) );
  INV_X1 us32_U209 (.A( us32_n792 ) , .ZN( us32_n851 ) );
  AOI222_X1 us32_U21 (.ZN( us32_n563 ) , .B1( us32_n830 ) , .C1( us32_n841 ) , .A2( us32_n843 ) , .A1( us32_n854 ) , .B2( us32_n863 ) , .C2( us32_n873 ) );
  NOR2_X1 us32_U210 (.A1( us32_n699 ) , .ZN( us32_n768 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U211 (.A1( us32_n669 ) , .ZN( us32_n673 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U212 (.ZN( us32_n541 ) , .A2( us32_n697 ) , .A1( us32_n699 ) );
  NOR2_X1 us32_U213 (.ZN( us32_n602 ) , .A1( us32_n669 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U214 (.A1( us32_n669 ) , .ZN( us32_n688 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U215 (.ZN( us32_n667 ) , .A1( us32_n750 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U216 (.ZN( us32_n555 ) , .A1( us32_n750 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U217 (.ZN( us32_n508 ) , .A2( us32_n780 ) , .A1( us32_n785 ) );
  NOR2_X1 us32_U218 (.ZN( us32_n543 ) , .A2( us32_n708 ) , .A1( us32_n785 ) );
  INV_X1 us32_U219 (.A( us32_n747 ) , .ZN( us32_n834 ) );
  AOI222_X1 us32_U22 (.ZN( us32_n660 ) , .A2( us32_n839 ) , .B1( us32_n841 ) , .C2( us32_n845 ) , .A1( us32_n860 ) , .C1( us32_n863 ) , .B2( us32_n870 ) );
  NOR2_X1 us32_U220 (.ZN( us32_n664 ) , .A1( us32_n785 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U221 (.A1( us32_n669 ) , .ZN( us32_n766 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U222 (.ZN( us32_n527 ) , .A1( us32_n669 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U223 (.ZN( us32_n661 ) , .A1( us32_n729 ) , .A2( us32_n790 ) );
  NOR2_X1 us32_U224 (.ZN( us32_n601 ) , .A2( us32_n780 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U225 (.ZN( us32_n507 ) , .A1( us32_n812 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U226 (.ZN( us32_n528 ) , .A2( us32_n724 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U227 (.ZN( us32_n509 ) , .A1( us32_n729 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U228 (.ZN( us32_n557 ) , .A1( us32_n792 ) , .A2( us32_n814 ) );
  NOR2_X1 us32_U229 (.ZN( us32_n545 ) , .A1( us32_n749 ) , .A2( us32_n814 ) );
  INV_X1 us32_U23 (.A( us32_n647 ) , .ZN( us32_n870 ) );
  OAI22_X1 us32_U230 (.B1( us32_n440 ) , .ZN( us32_n444 ) , .A2( us32_n728 ) , .A1( us32_n744 ) , .B2( us32_n749 ) );
  NOR3_X1 us32_U231 (.ZN( us32_n440 ) , .A2( us32_n836 ) , .A3( us32_n837 ) , .A1( us32_n846 ) );
  NOR2_X1 us32_U232 (.ZN( us32_n662 ) , .A2( us32_n697 ) , .A1( us32_n729 ) );
  OAI22_X1 us32_U233 (.B2( us32_n750 ) , .B1( us32_n751 ) , .A1( us32_n752 ) , .ZN( us32_n756 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U234 (.ZN( us32_n751 ) , .A2( us32_n852 ) , .A1( us32_n860 ) );
  NOR3_X1 us32_U235 (.ZN( us32_n752 ) , .A2( us32_n853 ) , .A1( us32_n863 ) , .A3( us32_n865 ) );
  NOR2_X1 us32_U236 (.ZN( us32_n544 ) , .A2( us32_n785 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U237 (.ZN( us32_n663 ) , .A1( us32_n729 ) , .A2( us32_n785 ) );
  INV_X1 us32_U238 (.A( us32_n806 ) , .ZN( us32_n841 ) );
  NOR2_X1 us32_U239 (.ZN( us32_n506 ) , .A2( us32_n728 ) , .A1( us32_n762 ) );
  NOR4_X1 us32_U24 (.A4( us32_n544 ) , .A3( us32_n545 ) , .A2( us32_n546 ) , .A1( us32_n547 ) , .ZN( us32_n548 ) );
  NOR2_X1 us32_U240 (.ZN( us32_n631 ) , .A1( us32_n724 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U241 (.ZN( us32_n614 ) , .A1( us32_n762 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U242 (.ZN( us32_n530 ) , .A2( us32_n744 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U243 (.ZN( us32_n558 ) , .A1( us32_n708 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U244 (.ZN( us32_n516 ) , .A1( us32_n708 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U245 (.A2( us32_n697 ) , .ZN( us32_n716 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U246 (.A1( us32_n749 ) , .ZN( us32_n767 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U247 (.ZN( us32_n521 ) , .A1( us32_n790 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U248 (.ZN( us32_n655 ) , .A1( us32_n790 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U249 (.ZN( us32_n668 ) , .A2( us32_n708 ) , .A1( us32_n790 ) );
  NOR4_X1 us32_U25 (.ZN( us32_n479 ) , .A1( us32_n520 ) , .A4( us32_n557 ) , .A3( us32_n582 ) , .A2( us32_n630 ) );
  NOR2_X1 us32_U250 (.ZN( us32_n517 ) , .A1( us32_n708 ) , .A2( us32_n803 ) );
  INV_X1 us32_U251 (.A( us32_n763 ) , .ZN( us32_n866 ) );
  NOR2_X1 us32_U252 (.ZN( us32_n542 ) , .A1( us32_n762 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U253 (.ZN( us32_n630 ) , .A1( us32_n747 ) , .A2( us32_n815 ) );
  INV_X1 us32_U254 (.A( us32_n729 ) , .ZN( us32_n868 ) );
  NOR2_X1 us32_U255 (.ZN( us32_n609 ) , .A2( us32_n724 ) , .A1( us32_n817 ) );
  AOI21_X1 us32_U256 (.A( us32_n815 ) , .B2( us32_n816 ) , .B1( us32_n817 ) , .ZN( us32_n818 ) );
  NOR2_X1 us32_U257 (.ZN( us32_n579 ) , .A2( us32_n708 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U258 (.ZN( us32_n533 ) , .A2( us32_n724 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U259 (.ZN( us32_n642 ) , .A2( us32_n788 ) , .A1( us32_n791 ) );
  NOR4_X1 us32_U26 (.ZN( us32_n456 ) , .A2( us32_n517 ) , .A1( us32_n543 ) , .A3( us32_n579 ) , .A4( us32_n615 ) );
  AOI21_X1 us32_U260 (.B1( us32_n625 ) , .ZN( us32_n627 ) , .A( us32_n763 ) , .B2( us32_n814 ) );
  NOR2_X1 us32_U261 (.ZN( us32_n656 ) , .A1( us32_n747 ) , .A2( us32_n780 ) );
  AOI21_X1 us32_U262 (.A( us32_n812 ) , .B2( us32_n813 ) , .B1( us32_n814 ) , .ZN( us32_n819 ) );
  NOR2_X1 us32_U263 (.A2( us32_n697 ) , .A1( us32_n780 ) , .ZN( us32_n820 ) );
  AOI21_X1 us32_U264 (.ZN( us32_n499 ) , .B1( us32_n680 ) , .A( us32_n812 ) , .B2( us32_n816 ) );
  NOR2_X1 us32_U265 (.A2( us32_n708 ) , .A1( us32_n762 ) , .ZN( us32_n794 ) );
  AOI21_X1 us32_U266 (.ZN( us32_n593 ) , .B1( us32_n750 ) , .A( us32_n792 ) , .B2( us32_n813 ) );
  AOI21_X1 us32_U267 (.ZN( us32_n626 ) , .B2( us32_n669 ) , .A( us32_n790 ) , .B1( us32_n791 ) );
  NOR2_X1 us32_U268 (.ZN( us32_n520 ) , .A2( us32_n708 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U269 (.A1( us32_n697 ) , .ZN( us32_n770 ) , .A2( us32_n815 ) );
  NOR4_X1 us32_U27 (.A4( us32_n532 ) , .A3( us32_n533 ) , .A2( us32_n534 ) , .ZN( us32_n535 ) , .A1( us32_n820 ) );
  NOR2_X1 us32_U270 (.ZN( us32_n582 ) , .A1( us32_n744 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U271 (.ZN( us32_n519 ) , .A2( us32_n699 ) , .A1( us32_n816 ) );
  AOI21_X1 us32_U272 (.ZN( us32_n477 ) , .A( us32_n669 ) , .B1( us32_n750 ) , .B2( us32_n806 ) );
  AOI21_X1 us32_U273 (.ZN( us32_n510 ) , .B2( us32_n669 ) , .A( us32_n730 ) , .B1( us32_n815 ) );
  INV_X1 us32_U274 (.A( us32_n813 ) , .ZN( us32_n836 ) );
  AOI21_X1 us32_U275 (.ZN( us32_n589 ) , .B2( us32_n699 ) , .B1( us32_n815 ) , .A( us32_n817 ) );
  AOI21_X1 us32_U276 (.ZN( us32_n515 ) , .A( us32_n729 ) , .B1( us32_n750 ) , .B2( us32_n803 ) );
  AOI21_X1 us32_U277 (.ZN( us32_n539 ) , .B2( us32_n812 ) , .A( us32_n814 ) , .B1( us32_n815 ) );
  NOR2_X1 us32_U278 (.ZN( us32_n581 ) , .A1( us32_n669 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U279 (.ZN( us32_n547 ) , .A1( us32_n699 ) , .A2( us32_n744 ) );
  NOR4_X1 us32_U28 (.ZN( us32_n474 ) , .A1( us32_n506 ) , .A3( us32_n544 ) , .A2( us32_n583 ) , .A4( us32_n716 ) );
  AOI21_X1 us32_U280 (.ZN( us32_n540 ) , .A( us32_n763 ) , .B2( us32_n779 ) , .B1( us32_n817 ) );
  AOI21_X1 us32_U281 (.B1( us32_n699 ) , .ZN( us32_n700 ) , .A( us32_n732 ) , .B2( us32_n763 ) );
  AOI21_X1 us32_U282 (.ZN( us32_n591 ) , .B2( us32_n763 ) , .A( us32_n785 ) , .B1( us32_n812 ) );
  INV_X1 us32_U283 (.A( us32_n791 ) , .ZN( us32_n873 ) );
  NOR2_X1 us32_U284 (.ZN( us32_n559 ) , .A2( us32_n791 ) , .A1( us32_n803 ) );
  AOI21_X1 us32_U285 (.ZN( us32_n498 ) , .A( us32_n724 ) , .B2( us32_n762 ) , .B1( us32_n814 ) );
  NOR2_X1 us32_U286 (.ZN( us32_n683 ) , .A2( us32_n699 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U287 (.ZN( us32_n685 ) , .A1( us32_n729 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U288 (.B1( us32_n686 ) , .ZN( us32_n687 ) , .A( us32_n728 ) , .B2( us32_n761 ) );
  AOI21_X1 us32_U289 (.ZN( us32_n569 ) , .B1( us32_n750 ) , .B2( us32_n762 ) , .A( us32_n780 ) );
  AOI221_X1 us32_U29 (.A( us32_n713 ) , .B2( us32_n714 ) , .ZN( us32_n720 ) , .C1( us32_n832 ) , .B1( us32_n839 ) , .C2( us32_n863 ) );
  AOI21_X1 us32_U290 (.ZN( us32_n649 ) , .B1( us32_n729 ) , .B2( us32_n763 ) , .A( us32_n813 ) );
  NOR2_X1 us32_U291 (.ZN( us32_n568 ) , .A1( us32_n729 ) , .A2( us32_n762 ) );
  INV_X1 us32_U292 (.A( us32_n699 ) , .ZN( us32_n853 ) );
  NOR2_X1 us32_U293 (.ZN( us32_n566 ) , .A2( us32_n697 ) , .A1( us32_n763 ) );
  AOI21_X1 us32_U294 (.ZN( us32_n514 ) , .A( us32_n779 ) , .B2( us32_n792 ) , .B1( us32_n812 ) );
  AOI21_X1 us32_U295 (.ZN( us32_n639 ) , .B2( us32_n749 ) , .A( us32_n788 ) , .B1( us32_n812 ) );
  NOR2_X1 us32_U296 (.ZN( us32_n665 ) , .A1( us32_n780 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U297 (.ZN( us32_n571 ) , .B2( us32_n697 ) , .B1( us32_n806 ) , .A( us32_n812 ) );
  AOI21_X1 us32_U298 (.ZN( us32_n564 ) , .B1( us32_n724 ) , .A( us32_n779 ) , .B2( us32_n791 ) );
  AOI21_X1 us32_U299 (.ZN( us32_n497 ) , .A( us32_n779 ) , .B2( us32_n791 ) , .B1( us32_n804 ) );
  NAND2_X1 us32_U3 (.A1( us32_n449 ) , .A2( us32_n464 ) , .ZN( us32_n724 ) );
  OR2_X1 us32_U30 (.A2( us32_n711 ) , .A1( us32_n712 ) , .ZN( us32_n713 ) );
  AOI21_X1 us32_U300 (.ZN( us32_n640 ) , .B2( us32_n747 ) , .A( us32_n792 ) , .B1( us32_n803 ) );
  NOR2_X1 us32_U301 (.ZN( us32_n578 ) , .A1( us32_n708 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U302 (.ZN( us32_n529 ) , .A1( us32_n708 ) , .A2( us32_n779 ) );
  AOI21_X1 us32_U303 (.ZN( us32_n689 ) , .B2( us32_n749 ) , .B1( us32_n763 ) , .A( us32_n806 ) );
  AOI21_X1 us32_U304 (.A( us32_n790 ) , .B2( us32_n791 ) , .B1( us32_n792 ) , .ZN( us32_n793 ) );
  AOI21_X1 us32_U305 (.ZN( us32_n478 ) , .B2( us32_n697 ) , .A( us32_n749 ) , .B1( us32_n779 ) );
  NOR2_X1 us32_U306 (.ZN( us32_n684 ) , .A1( us32_n791 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U307 (.ZN( us32_n450 ) , .B2( us32_n792 ) , .A( us32_n803 ) , .B1( us32_n815 ) );
  AOI21_X1 us32_U308 (.A( us32_n733 ) , .ZN( us32_n734 ) , .B2( us32_n780 ) , .B1( us32_n792 ) );
  NOR2_X1 us32_U309 (.A2( us32_n813 ) , .A1( us32_n815 ) , .ZN( us32_n821 ) );
  NOR2_X1 us32_U31 (.ZN( us32_n680 ) , .A2( us32_n834 ) , .A1( us32_n839 ) );
  AOI21_X1 us32_U310 (.ZN( us32_n641 ) , .B1( us32_n680 ) , .A( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U311 (.ZN( us32_n583 ) , .A1( us32_n792 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U312 (.ZN( us32_n711 ) , .A1( us32_n762 ) , .A2( us32_n763 ) );
  NOR2_X1 us32_U313 (.ZN( us32_n534 ) , .A1( us32_n724 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U314 (.ZN( us32_n632 ) , .A2( us32_n697 ) , .A1( us32_n724 ) );
  NOR2_X1 us32_U315 (.ZN( us32_n580 ) , .A2( us32_n697 ) , .A1( us32_n791 ) );
  NOR2_X1 us32_U316 (.ZN( us32_n682 ) , .A2( us32_n708 ) , .A1( us32_n817 ) );
  INV_X1 us32_U317 (.A( us32_n815 ) , .ZN( us32_n855 ) );
  AOI21_X1 us32_U318 (.ZN( us32_n442 ) , .A( us32_n699 ) , .B1( us32_n733 ) , .B2( us32_n750 ) );
  INV_X1 us32_U319 (.A( us32_n780 ) , .ZN( us32_n850 ) );
  NOR4_X1 us32_U32 (.A4( us32_n514 ) , .A3( us32_n515 ) , .A2( us32_n516 ) , .A1( us32_n517 ) , .ZN( us32_n524 ) );
  INV_X1 us32_U320 (.A( us32_n785 ) , .ZN( us32_n846 ) );
  NAND2_X1 us32_U321 (.ZN( us32_n714 ) , .A1( us32_n728 ) , .A2( us32_n780 ) );
  NAND2_X1 us32_U322 (.ZN( us32_n671 ) , .A1( us32_n806 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U323 (.ZN( us32_n443 ) , .B1( us32_n789 ) , .B2( us32_n791 ) , .A( us32_n814 ) );
  NOR2_X1 us32_U324 (.ZN( us32_n470 ) , .A2( us32_n779 ) , .A1( us32_n815 ) );
  NAND2_X1 us32_U325 (.A2( us32_n762 ) , .A1( us32_n806 ) , .ZN( us32_n810 ) );
  NOR2_X1 us32_U326 (.ZN( us32_n526 ) , .A1( us32_n724 ) , .A2( us32_n750 ) );
  OAI21_X1 us32_U327 (.A( us32_n787 ) , .B2( us32_n788 ) , .B1( us32_n789 ) , .ZN( us32_n795 ) );
  OAI21_X1 us32_U328 (.ZN( us32_n787 ) , .A( us32_n839 ) , .B1( us32_n863 ) , .B2( us32_n873 ) );
  NAND2_X1 us32_U329 (.A1( us32_n699 ) , .A2( us32_n729 ) , .ZN( us32_n782 ) );
  AOI222_X1 us32_U33 (.ZN( us32_n525 ) , .A1( us32_n834 ) , .B2( us32_n837 ) , .C1( us32_n844 ) , .C2( us32_n850 ) , .A2( us32_n852 ) , .B1( us32_n866 ) );
  NOR2_X1 us32_U330 (.ZN( us32_n712 ) , .A2( us32_n724 ) , .A1( us32_n790 ) );
  NOR2_X1 us32_U331 (.ZN( us32_n518 ) , .A1( us32_n708 ) , .A2( us32_n788 ) );
  OAI21_X1 us32_U332 (.A( us32_n698 ) , .ZN( us32_n702 ) , .B2( us32_n750 ) , .B1( us32_n804 ) );
  OAI21_X1 us32_U333 (.ZN( us32_n698 ) , .B2( us32_n833 ) , .B1( us32_n838 ) , .A( us32_n860 ) );
  INV_X1 us32_U334 (.A( us32_n817 ) , .ZN( us32_n844 ) );
  INV_X1 us32_U335 (.A( us32_n724 ) , .ZN( us32_n856 ) );
  OAI21_X1 us32_U336 (.ZN( us32_n731 ) , .A( us32_n833 ) , .B2( us32_n852 ) , .B1( us32_n873 ) );
  AND2_X1 us32_U337 (.ZN( us32_n732 ) , .A1( us32_n779 ) , .A2( us32_n785 ) );
  AOI221_X1 us32_U338 (.A( us32_n764 ) , .ZN( us32_n774 ) , .C2( us32_n810 ) , .B2( us32_n835 ) , .C1( us32_n855 ) , .B1( us32_n866 ) );
  AOI21_X1 us32_U339 (.B2( us32_n763 ) , .ZN( us32_n764 ) , .A( us32_n788 ) , .B1( us32_n792 ) );
  NOR4_X1 us32_U34 (.A3( us32_n521 ) , .A1( us32_n522 ) , .ZN( us32_n523 ) , .A2( us32_n673 ) , .A4( us32_n769 ) );
  INV_X1 us32_U340 (.A( us32_n761 ) , .ZN( us32_n835 ) );
  NAND2_X1 us32_U341 (.A2( us32_n448 ) , .A1( us32_n460 ) , .ZN( us32_n728 ) );
  NAND2_X1 us32_U342 (.A1( us32_n451 ) , .A2( us32_n454 ) , .ZN( us32_n814 ) );
  NAND2_X1 us32_U343 (.A1( us32_n455 ) , .A2( us32_n462 ) , .ZN( us32_n750 ) );
  NAND2_X1 us32_U344 (.A1( us32_n451 ) , .A2( us32_n471 ) , .ZN( us32_n816 ) );
  NAND2_X1 us32_U345 (.A1( us32_n454 ) , .A2( us32_n461 ) , .ZN( us32_n813 ) );
  NAND2_X1 us32_U346 (.A1( us32_n452 ) , .A2( us32_n465 ) , .ZN( us32_n669 ) );
  NAND2_X1 us32_U347 (.A1( us32_n453 ) , .A2( us32_n472 ) , .ZN( us32_n785 ) );
  NAND2_X1 us32_U348 (.A1( us32_n453 ) , .A2( us32_n461 ) , .ZN( us32_n744 ) );
  NAND2_X1 us32_U349 (.A2( us32_n453 ) , .A1( us32_n455 ) , .ZN( us32_n806 ) );
  AOI221_X1 us32_U35 (.A( us32_n781 ) , .ZN( us32_n798 ) , .C2( us32_n837 ) , .B2( us32_n838 ) , .B1( us32_n865 ) , .C1( us32_n866 ) );
  NAND2_X1 us32_U350 (.A1( us32_n455 ) , .A2( us32_n471 ) , .ZN( us32_n803 ) );
  NAND2_X1 us32_U351 (.A2( us32_n454 ) , .A1( us32_n472 ) , .ZN( us32_n779 ) );
  NAND2_X1 us32_U352 (.A2( us32_n464 ) , .A1( us32_n465 ) , .ZN( us32_n812 ) );
  NAND2_X1 us32_U353 (.A1( us32_n441 ) , .A2( us32_n460 ) , .ZN( us32_n699 ) );
  NAND2_X1 us32_U354 (.A2( us32_n448 ) , .A1( us32_n452 ) , .ZN( us32_n729 ) );
  NAND2_X1 us32_U355 (.A2( us32_n449 ) , .A1( us32_n452 ) , .ZN( us32_n763 ) );
  NOR2_X1 us32_U356 (.ZN( us32_n465 ) , .A2( us32_n847 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U357 (.ZN( us32_n453 ) , .A1( us32_n826 ) , .A2( us32_n827 ) );
  NAND2_X1 us32_U358 (.A1( us32_n462 ) , .A2( us32_n472 ) , .ZN( us32_n788 ) );
  NOR2_X1 us32_U359 (.ZN( us32_n451 ) , .A1( us32_n828 ) , .A2( us32_n829 ) );
  NOR4_X1 us32_U36 (.A4( us32_n793 ) , .A3( us32_n794 ) , .A2( us32_n795 ) , .A1( us32_n796 ) , .ZN( us32_n797 ) );
  NAND2_X1 us32_U360 (.A2( us32_n461 ) , .A1( us32_n462 ) , .ZN( us32_n747 ) );
  NAND2_X1 us32_U361 (.A1( us32_n451 ) , .A2( us32_n462 ) , .ZN( us32_n790 ) );
  NAND2_X2 us32_U362 (.A2( us32_n448 ) , .A1( us32_n464 ) , .ZN( us32_n815 ) );
  NAND2_X1 us32_U363 (.A2( us32_n441 ) , .A1( us32_n447 ) , .ZN( us32_n784 ) );
  NAND2_X1 us32_U364 (.A1( us32_n447 ) , .A2( us32_n449 ) , .ZN( us32_n805 ) );
  NAND2_X1 us32_U365 (.A2( us32_n454 ) , .A1( us32_n455 ) , .ZN( us32_n730 ) );
  NAND2_X2 us32_U366 (.A1( us32_n449 ) , .A2( us32_n460 ) , .ZN( us32_n792 ) );
  NAND2_X2 us32_U367 (.A2( us32_n460 ) , .A1( us32_n465 ) , .ZN( us32_n780 ) );
  NOR2_X1 us32_U368 (.ZN( us32_n447 ) , .A2( us32_n849 ) , .A1( us32_n858 ) );
  NAND2_X1 us32_U369 (.A1( us32_n447 ) , .A2( us32_n448 ) , .ZN( us32_n786 ) );
  NOR4_X1 us32_U37 (.A4( us32_n776 ) , .A3( us32_n777 ) , .A1( us32_n778 ) , .ZN( us32_n799 ) , .A2( us32_n801 ) );
  NAND2_X1 us32_U370 (.A2( us32_n471 ) , .A1( us32_n472 ) , .ZN( us32_n817 ) );
  NOR2_X1 us32_U371 (.A2( sa32_6 ) , .A1( sa32_7 ) , .ZN( us32_n464 ) );
  NOR2_X1 us32_U372 (.A2( sa32_7 ) , .ZN( us32_n460 ) , .A1( us32_n849 ) );
  NOR2_X1 us32_U373 (.A2( sa32_4 ) , .ZN( us32_n449 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U374 (.A2( sa32_4 ) , .A1( sa32_5 ) , .ZN( us32_n441 ) );
  NOR2_X1 us32_U375 (.A2( sa32_5 ) , .ZN( us32_n448 ) , .A1( us32_n847 ) );
  NOR2_X1 us32_U376 (.A2( sa32_2 ) , .A1( sa32_3 ) , .ZN( us32_n472 ) );
  NOR2_X1 us32_U377 (.A2( sa32_6 ) , .ZN( us32_n452 ) , .A1( us32_n858 ) );
  NOR2_X1 us32_U378 (.A2( sa32_1 ) , .ZN( us32_n471 ) , .A1( us32_n826 ) );
  NOR2_X1 us32_U379 (.A2( sa32_0 ) , .ZN( us32_n454 ) , .A1( us32_n827 ) );
  NOR4_X1 us32_U38 (.A3( us32_n755 ) , .A2( us32_n756 ) , .A1( us32_n757 ) , .ZN( us32_n758 ) , .A4( us32_n869 ) );
  NOR2_X1 us32_U380 (.A2( sa32_0 ) , .A1( sa32_1 ) , .ZN( us32_n462 ) );
  NOR2_X1 us32_U381 (.A2( sa32_3 ) , .ZN( us32_n455 ) , .A1( us32_n828 ) );
  NOR2_X1 us32_U382 (.A2( sa32_2 ) , .ZN( us32_n461 ) , .A1( us32_n829 ) );
  INV_X1 us32_U383 (.A( sa32_4 ) , .ZN( us32_n847 ) );
  INV_X1 us32_U384 (.A( sa32_6 ) , .ZN( us32_n849 ) );
  INV_X1 us32_U385 (.A( sa32_3 ) , .ZN( us32_n829 ) );
  INV_X1 us32_U386 (.A( sa32_1 ) , .ZN( us32_n827 ) );
  INV_X1 us32_U387 (.A( sa32_0 ) , .ZN( us32_n826 ) );
  INV_X1 us32_U388 (.A( sa32_2 ) , .ZN( us32_n828 ) );
  INV_X1 us32_U389 (.A( sa32_5 ) , .ZN( us32_n848 ) );
  AOI211_X1 us32_U39 (.B( us32_n745 ) , .A( us32_n746 ) , .ZN( us32_n759 ) , .C1( us32_n832 ) , .C2( us32_n853 ) );
  INV_X1 us32_U390 (.A( sa32_7 ) , .ZN( us32_n858 ) );
  NAND2_X1 us32_U391 (.A2( us32_n461 ) , .A1( us32_n471 ) , .ZN( us32_n697 ) );
  OAI222_X1 us32_U392 (.B2( us32_n747 ) , .B1( us32_n748 ) , .A2( us32_n749 ) , .ZN( us32_n757 ) , .C2( us32_n805 ) , .C1( us32_n814 ) , .A1( us32_n817 ) );
  OAI22_X1 us32_U393 (.B2( us32_n803 ) , .B1( us32_n804 ) , .A2( us32_n805 ) , .A1( us32_n806 ) , .ZN( us32_n808 ) );
  OAI21_X1 us32_U394 (.A( us32_n731 ) , .B1( us32_n732 ) , .ZN( us32_n736 ) , .B2( us32_n805 ) );
  OAI222_X1 us32_U395 (.ZN( us32_n505 ) , .C2( us32_n625 ) , .B2( us32_n647 ) , .B1( us32_n747 ) , .A2( us32_n748 ) , .C1( us32_n805 ) , .A1( us32_n806 ) );
  AOI21_X1 us32_U396 (.ZN( us32_n650 ) , .A( us32_n779 ) , .B1( us32_n792 ) , .B2( us32_n805 ) );
  INV_X1 us32_U397 (.A( us32_n805 ) , .ZN( us32_n860 ) );
  NOR2_X1 us32_U398 (.ZN( us32_n735 ) , .A2( us32_n803 ) , .A1( us32_n805 ) );
  NOR2_X1 us32_U399 (.ZN( us32_n484 ) , .A1( us32_n788 ) , .A2( us32_n805 ) );
  NAND2_X1 us32_U4 (.A1( us32_n441 ) , .A2( us32_n464 ) , .ZN( us32_n708 ) );
  NOR3_X1 us32_U40 (.A3( us32_n741 ) , .A2( us32_n742 ) , .A1( us32_n743 ) , .ZN( us32_n760 ) );
  NOR2_X1 us32_U400 (.A2( us32_n744 ) , .ZN( us32_n755 ) , .A1( us32_n805 ) );
  NAND2_X1 us32_U401 (.ZN( us32_n753 ) , .A1( us32_n763 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U402 (.ZN( us32_n715 ) , .A1( us32_n805 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U403 (.ZN( us32_n567 ) , .A1( us32_n747 ) , .A2( us32_n805 ) );
  AOI21_X1 us32_U404 (.ZN( us32_n552 ) , .B1( us32_n669 ) , .A( us32_n697 ) , .B2( us32_n805 ) );
  NOR2_X1 us32_U405 (.ZN( us32_n556 ) , .A1( us32_n762 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U406 (.ZN( us32_n670 ) , .A1( us32_n790 ) , .A2( us32_n805 ) );
  OAI221_X1 us32_U407 (.A( us32_n783 ) , .C2( us32_n784 ) , .B2( us32_n785 ) , .B1( us32_n786 ) , .ZN( us32_n796 ) , .C1( us32_n813 ) );
  NAND2_X1 us32_U408 (.A1( us32_n729 ) , .A2( us32_n784 ) , .ZN( us32_n811 ) );
  OAI22_X1 us32_U409 (.ZN( us32_n588 ) , .A2( us32_n747 ) , .B2( us32_n762 ) , .A1( us32_n763 ) , .B1( us32_n784 ) );
  NAND4_X1 us32_U41 (.ZN( sa33_sr_3 ) , .A4( us32_n704 ) , .A3( us32_n705 ) , .A2( us32_n706 ) , .A1( us32_n707 ) );
  AOI21_X1 us32_U410 (.ZN( us32_n592 ) , .B1( us32_n728 ) , .B2( us32_n784 ) , .A( us32_n790 ) );
  AOI21_X1 us32_U411 (.ZN( us32_n623 ) , .B1( us32_n699 ) , .A( us32_n779 ) , .B2( us32_n784 ) );
  AOI21_X1 us32_U412 (.ZN( us32_n648 ) , .A( us32_n762 ) , .B2( us32_n784 ) , .B1( us32_n792 ) );
  OAI22_X1 us32_U413 (.ZN( us32_n681 ) , .A1( us32_n699 ) , .A2( us32_n730 ) , .B2( us32_n784 ) , .B1( us32_n817 ) );
  OAI21_X1 us32_U414 (.A( us32_n613 ) , .ZN( us32_n616 ) , .B1( us32_n625 ) , .B2( us32_n784 ) );
  NOR2_X1 us32_U415 (.ZN( us32_n610 ) , .A1( us32_n784 ) , .A2( us32_n816 ) );
  OAI222_X1 us32_U416 (.A2( us32_n669 ) , .ZN( us32_n674 ) , .B1( us32_n747 ) , .B2( us32_n784 ) , .C2( us32_n788 ) , .C1( us32_n815 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U417 (.ZN( us32_n651 ) , .A1( us32_n784 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U418 (.ZN( us32_n600 ) , .A2( us32_n697 ) , .A1( us32_n784 ) );
  NOR2_X1 us32_U419 (.ZN( us32_n553 ) , .A2( us32_n744 ) , .A1( us32_n784 ) );
  NOR4_X1 us32_U42 (.A4( us32_n700 ) , .A3( us32_n701 ) , .A2( us32_n702 ) , .A1( us32_n703 ) , .ZN( us32_n704 ) );
  INV_X1 us32_U420 (.A( us32_n784 ) , .ZN( us32_n861 ) );
  AOI21_X1 us32_U421 (.ZN( us32_n500 ) , .A( us32_n697 ) , .B1( us32_n708 ) , .B2( us32_n786 ) );
  OAI221_X1 us32_U422 (.A( us32_n696 ) , .ZN( us32_n703 ) , .C2( us32_n784 ) , .C1( us32_n785 ) , .B1( us32_n786 ) , .B2( us32_n806 ) );
  OAI22_X1 us32_U423 (.ZN( us32_n590 ) , .B1( us32_n730 ) , .B2( us32_n749 ) , .A2( us32_n786 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U424 (.ZN( us32_n612 ) , .A1( us32_n779 ) , .A2( us32_n786 ) );
  NAND2_X1 us32_U425 (.A2( us32_n749 ) , .A1( us32_n786 ) , .ZN( us32_n809 ) );
  OAI222_X1 us32_U426 (.ZN( us32_n617 ) , .B1( us32_n697 ) , .C1( us32_n724 ) , .C2( us32_n747 ) , .B2( us32_n786 ) , .A2( us32_n792 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U427 (.ZN( us32_n717 ) , .A2( us32_n744 ) , .A1( us32_n786 ) );
  NOR2_X1 us32_U428 (.ZN( us32_n653 ) , .A1( us32_n762 ) , .A2( us32_n786 ) );
  NOR2_X1 us32_U429 (.ZN( us32_n554 ) , .A1( us32_n786 ) , .A2( us32_n813 ) );
  AOI211_X1 us32_U43 (.B( us32_n694 ) , .A( us32_n695 ) , .ZN( us32_n705 ) , .C2( us32_n831 ) , .C1( us32_n851 ) );
  NOR2_X1 us32_U430 (.ZN( us32_n701 ) , .A2( us32_n786 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U431 (.A1( us32_n730 ) , .ZN( us32_n765 ) , .A2( us32_n786 ) );
  AND2_X1 us32_U432 (.ZN( us32_n438 ) , .A2( us32_n831 ) , .A1( us32_n854 ) );
  AND2_X1 us32_U433 (.ZN( us32_n439 ) , .A2( us32_n843 ) , .A1( us32_n861 ) );
  NOR3_X1 us32_U434 (.A1( us32_n438 ) , .A2( us32_n439 ) , .A3( us32_n576 ) , .ZN( us32_n587 ) );
  NAND4_X1 us32_U435 (.ZN( sa33_sr_2 ) , .A4( us32_n643 ) , .A3( us32_n644 ) , .A2( us32_n645 ) , .A1( us32_n646 ) );
  INV_X1 us32_U436 (.A( us32_n812 ) , .ZN( us32_n854 ) );
  NAND3_X1 us32_U437 (.ZN( sa33_sr_6 ) , .A3( us32_n797 ) , .A2( us32_n798 ) , .A1( us32_n799 ) );
  NAND3_X1 us32_U438 (.ZN( sa33_sr_5 ) , .A3( us32_n758 ) , .A2( us32_n759 ) , .A1( us32_n760 ) );
  NAND3_X1 us32_U439 (.ZN( sa33_sr_4 ) , .A3( us32_n738 ) , .A2( us32_n739 ) , .A1( us32_n740 ) );
  NOR2_X1 us32_U44 (.ZN( us32_n707 ) , .A2( us32_n776 ) , .A1( us32_n800 ) );
  NAND3_X1 us32_U440 (.A3( us32_n675 ) , .A2( us32_n676 ) , .A1( us32_n677 ) , .ZN( us32_n807 ) );
  NAND3_X1 us32_U441 (.ZN( us32_n638 ) , .A3( us32_n708 ) , .A2( us32_n724 ) , .A1( us32_n792 ) );
  NAND3_X1 us32_U442 (.A3( us32_n618 ) , .A2( us32_n619 ) , .A1( us32_n620 ) , .ZN( us32_n725 ) );
  NAND3_X1 us32_U443 (.A3( us32_n585 ) , .A2( us32_n586 ) , .A1( us32_n587 ) , .ZN( us32_n621 ) );
  NAND3_X1 us32_U444 (.ZN( us32_n565 ) , .A3( us32_n680 ) , .A2( us32_n750 ) , .A1( us32_n785 ) );
  NAND3_X1 us32_U445 (.A3( us32_n523 ) , .A2( us32_n524 ) , .A1( us32_n525 ) , .ZN( us32_n742 ) );
  NAND3_X1 us32_U446 (.A3( us32_n512 ) , .A1( us32_n513 ) , .ZN( us32_n608 ) , .A2( us32_n871 ) );
  NAND3_X1 us32_U447 (.A3( us32_n467 ) , .A2( us32_n468 ) , .A1( us32_n469 ) , .ZN( us32_n777 ) );
  INV_X1 us32_U448 (.A( us32_n803 ) , .ZN( us32_n843 ) );
  AOI21_X1 us32_U449 (.ZN( us32_n576 ) , .B2( us32_n724 ) , .B1( us32_n748 ) , .A( us32_n785 ) );
  AOI222_X1 us32_U45 (.B2( us32_n638 ) , .ZN( us32_n644 ) , .B1( us32_n841 ) , .A1( us32_n842 ) , .C2( us32_n846 ) , .C1( us32_n863 ) , .A2( us32_n865 ) );
  NOR4_X1 us32_U46 (.A4( us32_n639 ) , .A3( us32_n640 ) , .A2( us32_n641 ) , .A1( us32_n642 ) , .ZN( us32_n643 ) );
  NOR3_X1 us32_U47 (.A2( us32_n607 ) , .A1( us32_n608 ) , .ZN( us32_n646 ) , .A3( us32_n722 ) );
  NAND4_X1 us32_U48 (.ZN( sa33_sr_7 ) , .A4( us32_n822 ) , .A3( us32_n823 ) , .A2( us32_n824 ) , .A1( us32_n825 ) );
  NOR4_X1 us32_U49 (.A4( us32_n818 ) , .A3( us32_n819 ) , .A2( us32_n820 ) , .A1( us32_n821 ) , .ZN( us32_n822 ) );
  NAND2_X1 us32_U5 (.A2( us32_n441 ) , .A1( us32_n452 ) , .ZN( us32_n791 ) );
  AOI222_X1 us32_U50 (.C2( us32_n809 ) , .B2( us32_n810 ) , .A2( us32_n811 ) , .ZN( us32_n823 ) , .C1( us32_n832 ) , .A1( us32_n839 ) , .B1( us32_n853 ) );
  AOI211_X1 us32_U51 (.B( us32_n807 ) , .A( us32_n808 ) , .ZN( us32_n824 ) , .C1( us32_n842 ) , .C2( us32_n850 ) );
  NAND4_X1 us32_U52 (.ZN( sa33_sr_0 ) , .A4( us32_n501 ) , .A3( us32_n502 ) , .A2( us32_n503 ) , .A1( us32_n504 ) );
  AOI221_X1 us32_U53 (.A( us32_n497 ) , .ZN( us32_n502 ) , .B2( us32_n843 ) , .C1( us32_n846 ) , .C2( us32_n860 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U54 (.A4( us32_n498 ) , .A3( us32_n499 ) , .A2( us32_n500 ) , .ZN( us32_n501 ) , .A1( us32_n527 ) );
  AOI211_X1 us32_U55 (.A( us32_n496 ) , .ZN( us32_n503 ) , .B( us32_n802 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NAND4_X1 us32_U56 (.ZN( sa33_sr_1 ) , .A4( us32_n595 ) , .A3( us32_n596 ) , .A2( us32_n597 ) , .A1( us32_n598 ) );
  NOR4_X1 us32_U57 (.A4( us32_n591 ) , .A3( us32_n592 ) , .A2( us32_n593 ) , .A1( us32_n594 ) , .ZN( us32_n595 ) );
  AOI211_X1 us32_U58 (.B( us32_n589 ) , .A( us32_n590 ) , .ZN( us32_n596 ) , .C2( us32_n811 ) , .C1( us32_n833 ) );
  AOI211_X1 us32_U59 (.A( us32_n588 ) , .ZN( us32_n597 ) , .B( us32_n621 ) , .C1( us32_n845 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U6 (.ZN( us32_n598 ) , .A1( us32_n608 ) , .A3( us32_n723 ) , .A2( us32_n742 ) );
  NOR2_X1 us32_U60 (.ZN( us32_n804 ) , .A1( us32_n854 ) , .A2( us32_n861 ) );
  AOI222_X1 us32_U61 (.ZN( us32_n469 ) , .B1( us32_n832 ) , .A1( us32_n839 ) , .C1( us32_n842 ) , .C2( us32_n851 ) , .A2( us32_n855 ) , .B2( us32_n865 ) );
  NOR4_X1 us32_U62 (.A1( us32_n466 ) , .ZN( us32_n467 ) , .A4( us32_n542 ) , .A2( us32_n554 ) , .A3( us32_n614 ) );
  AOI221_X1 us32_U63 (.ZN( us32_n468 ) , .C2( us32_n714 ) , .B2( us32_n831 ) , .C1( us32_n845 ) , .B1( us32_n860 ) , .A( us32_n864 ) );
  NAND4_X1 us32_U64 (.A4( us32_n603 ) , .A3( us32_n604 ) , .A2( us32_n605 ) , .A1( us32_n606 ) , .ZN( us32_n722 ) );
  NOR3_X1 us32_U65 (.A1( us32_n599 ) , .ZN( us32_n604 ) , .A3( us32_n663 ) , .A2( us32_n770 ) );
  NOR4_X1 us32_U66 (.A3( us32_n600 ) , .A2( us32_n601 ) , .A1( us32_n602 ) , .ZN( us32_n603 ) , .A4( us32_n655 ) );
  AOI222_X1 us32_U67 (.ZN( us32_n606 ) , .A1( us32_n830 ) , .C2( us32_n837 ) , .B1( us32_n842 ) , .A2( us32_n856 ) , .B2( us32_n861 ) , .C1( us32_n868 ) );
  NAND4_X1 us32_U68 (.A4( us32_n657 ) , .A3( us32_n658 ) , .A2( us32_n659 ) , .A1( us32_n660 ) , .ZN( us32_n800 ) );
  NOR3_X1 us32_U69 (.A3( us32_n648 ) , .A2( us32_n649 ) , .A1( us32_n650 ) , .ZN( us32_n659 ) );
  NOR3_X1 us32_U7 (.A3( us32_n800 ) , .A2( us32_n801 ) , .A1( us32_n802 ) , .ZN( us32_n825 ) );
  NOR3_X1 us32_U70 (.A3( us32_n651 ) , .A2( us32_n652 ) , .A1( us32_n653 ) , .ZN( us32_n658 ) );
  NOR3_X1 us32_U71 (.A3( us32_n654 ) , .A2( us32_n655 ) , .A1( us32_n656 ) , .ZN( us32_n657 ) );
  NAND4_X1 us32_U72 (.A4( us32_n560 ) , .A3( us32_n561 ) , .A2( us32_n562 ) , .A1( us32_n563 ) , .ZN( us32_n607 ) );
  NOR4_X1 us32_U73 (.A4( us32_n556 ) , .A3( us32_n557 ) , .A2( us32_n558 ) , .A1( us32_n559 ) , .ZN( us32_n560 ) );
  NOR4_X1 us32_U74 (.ZN( us32_n561 ) , .A1( us32_n653 ) , .A3( us32_n661 ) , .A4( us32_n685 ) , .A2( us32_n768 ) );
  NOR4_X1 us32_U75 (.A4( us32_n552 ) , .A3( us32_n553 ) , .A2( us32_n554 ) , .A1( us32_n555 ) , .ZN( us32_n562 ) );
  NAND4_X1 us32_U76 (.A4( us32_n772 ) , .A3( us32_n773 ) , .A2( us32_n774 ) , .A1( us32_n775 ) , .ZN( us32_n801 ) );
  NOR3_X1 us32_U77 (.A3( us32_n765 ) , .A2( us32_n766 ) , .A1( us32_n767 ) , .ZN( us32_n773 ) );
  NOR4_X1 us32_U78 (.A4( us32_n768 ) , .A3( us32_n769 ) , .A2( us32_n770 ) , .A1( us32_n771 ) , .ZN( us32_n772 ) );
  AOI222_X1 us32_U79 (.ZN( us32_n775 ) , .A1( us32_n830 ) , .C1( us32_n834 ) , .B2( us32_n841 ) , .A2( us32_n850 ) , .B1( us32_n861 ) , .C2( us32_n873 ) );
  NOR3_X1 us32_U8 (.A3( us32_n621 ) , .A2( us32_n622 ) , .ZN( us32_n636 ) , .A1( us32_n725 ) );
  NOR4_X1 us32_U80 (.A4( us32_n665 ) , .A3( us32_n666 ) , .A2( us32_n667 ) , .A1( us32_n668 ) , .ZN( us32_n676 ) );
  NOR4_X1 us32_U81 (.A4( us32_n661 ) , .A3( us32_n662 ) , .A2( us32_n663 ) , .A1( us32_n664 ) , .ZN( us32_n677 ) );
  NOR4_X1 us32_U82 (.A3( us32_n673 ) , .A1( us32_n674 ) , .ZN( us32_n675 ) , .A4( us32_n715 ) , .A2( us32_n859 ) );
  NOR2_X1 us32_U83 (.ZN( us32_n625 ) , .A2( us32_n836 ) , .A1( us32_n839 ) );
  NOR2_X1 us32_U84 (.ZN( us32_n761 ) , .A1( us32_n833 ) , .A2( us32_n834 ) );
  NOR4_X1 us32_U85 (.A4( us32_n577 ) , .A3( us32_n578 ) , .A2( us32_n579 ) , .ZN( us32_n586 ) , .A1( us32_n683 ) );
  NOR4_X1 us32_U86 (.A1( us32_n584 ) , .ZN( us32_n585 ) , .A3( us32_n652 ) , .A2( us32_n662 ) , .A4( us32_n767 ) );
  AOI222_X1 us32_U87 (.ZN( us32_n513 ) , .C1( us32_n832 ) , .B2( us32_n837 ) , .A2( us32_n843 ) , .C2( us32_n862 ) , .B1( us32_n863 ) , .A1( us32_n866 ) );
  NOR4_X1 us32_U88 (.A4( us32_n509 ) , .A2( us32_n510 ) , .A1( us32_n511 ) , .ZN( us32_n512 ) , .A3( us32_n670 ) );
  INV_X1 us32_U89 (.A( us32_n505 ) , .ZN( us32_n871 ) );
  NOR2_X1 us32_U9 (.ZN( us32_n495 ) , .A1( us32_n678 ) , .A2( us32_n694 ) );
  NAND4_X1 us32_U90 (.A4( us32_n456 ) , .A3( us32_n457 ) , .A2( us32_n458 ) , .A1( us32_n459 ) , .ZN( us32_n679 ) );
  NOR3_X1 us32_U91 (.ZN( us32_n457 ) , .A3( us32_n530 ) , .A1( us32_n555 ) , .A2( us32_n570 ) );
  AOI221_X1 us32_U92 (.A( us32_n450 ) , .ZN( us32_n459 ) , .C2( us32_n753 ) , .B1( us32_n832 ) , .C1( us32_n842 ) , .B2( us32_n861 ) );
  NOR4_X1 us32_U93 (.ZN( us32_n458 ) , .A2( us32_n509 ) , .A1( us32_n599 ) , .A4( us32_n628 ) , .A3( us32_n711 ) );
  NAND4_X1 us32_U94 (.A4( us32_n535 ) , .A3( us32_n536 ) , .A2( us32_n537 ) , .A1( us32_n538 ) , .ZN( us32_n622 ) );
  NOR4_X1 us32_U95 (.A4( us32_n526 ) , .A2( us32_n527 ) , .A1( us32_n528 ) , .ZN( us32_n538 ) , .A3( us32_n701 ) );
  NOR4_X1 us32_U96 (.A1( us32_n531 ) , .ZN( us32_n536 ) , .A2( us32_n654 ) , .A4( us32_n668 ) , .A3( us32_n765 ) );
  NOR4_X1 us32_U97 (.A4( us32_n529 ) , .A3( us32_n530 ) , .ZN( us32_n537 ) , .A2( us32_n684 ) , .A1( us32_n794 ) );
  NAND4_X1 us32_U98 (.A4( us32_n479 ) , .A3( us32_n480 ) , .A2( us32_n481 ) , .A1( us32_n482 ) , .ZN( us32_n694 ) );
  NOR3_X1 us32_U99 (.ZN( us32_n480 ) , .A2( us32_n508 ) , .A3( us32_n601 ) , .A1( us32_n610 ) );
endmodule

