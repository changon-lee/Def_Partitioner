module des_des_die_3 ( u0_K15_47, u0_L13_12, u0_L13_15, u0_L13_21, u0_L13_22, u0_L13_27, u0_L13_32, u0_L13_5, u0_L13_7, 
       u0_R13_1, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
       u0_R13_32, u0_key_r_18, u0_uk_K_r0_52, u0_uk_K_r13_2, u0_uk_K_r13_23, u0_uk_K_r13_35, u0_uk_K_r9_5, u0_uk_n10, u0_uk_n12, 
       u0_uk_n128, u0_uk_n13, u0_uk_n141, u0_uk_n155, u0_uk_n163, u0_uk_n17, u0_uk_n187, u0_uk_n21, u0_uk_n22, 
       u0_uk_n220, u0_uk_n23, u0_uk_n27, u0_uk_n3, u0_uk_n34, u0_uk_n39, u0_uk_n4, u0_uk_n40, u0_uk_n41, 
       u0_uk_n5, u0_uk_n9, u0_uk_n916, u0_uk_n93, u1_FP_40, u1_FP_41, u1_FP_42, u1_FP_43, u1_FP_44, 
       u1_FP_45, u1_L0_13, u1_L0_16, u1_L0_18, u1_L0_2, u1_L0_24, u1_L0_28, u1_L0_30, u1_L0_6, 
       u1_L11_1, u1_L11_10, u1_L11_13, u1_L11_17, u1_L11_18, u1_L11_2, u1_L11_20, u1_L11_23, u1_L11_26, 
       u1_L11_28, u1_L11_31, u1_L11_9, u1_L14_16, u1_L14_24, u1_L14_30, u1_L14_6, u1_L3_13, u1_L3_18, 
       u1_L3_2, u1_L3_28, u1_L8_13, u1_L8_16, u1_L8_17, u1_L8_18, u1_L8_2, u1_L8_23, u1_L8_24, 
       u1_L8_28, u1_L8_30, u1_L8_31, u1_L8_6, u1_L8_9, u1_L9_11, u1_L9_13, u1_L9_16, u1_L9_17, 
       u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_23, u1_L9_24, u1_L9_28, u1_L9_29, u1_L9_30, u1_L9_31, 
       u1_L9_4, u1_L9_6, u1_L9_9, u1_R0_10, u1_R0_11, u1_R0_12, u1_R0_13, u1_R0_4, u1_R0_5, 
       u1_R0_6, u1_R0_7, u1_R0_8, u1_R0_9, u1_R11_1, u1_R11_12, u1_R11_13, u1_R11_14, u1_R11_15, 
       u1_R11_16, u1_R11_17, u1_R11_2, u1_R11_3, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_6, u1_R11_7, 
       u1_R11_8, u1_R11_9, u1_R3_4, u1_R3_5, u1_R3_6, u1_R3_7, u1_R3_8, u1_R3_9, u1_R8_1, 
       u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_2, u1_R8_3, u1_R8_32, u1_R8_4, u1_R8_5, 
       u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_10, u1_R9_11, u1_R9_12, u1_R9_13, 
       u1_R9_2, u1_R9_20, u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_3, u1_R9_32, 
       u1_R9_4, u1_R9_5, u1_R9_6, u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_10, u1_desIn_r_12, u1_desIn_r_13, 
       u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_2, u1_desIn_r_21, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_26, u1_desIn_r_29, u1_desIn_r_3, 
       u1_desIn_r_31, u1_desIn_r_36, u1_desIn_r_37, u1_desIn_r_39, u1_desIn_r_4, u1_desIn_r_40, u1_desIn_r_45, u1_desIn_r_46, u1_desIn_r_47, 
       u1_desIn_r_48, u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_53, u1_desIn_r_55, u1_desIn_r_57, u1_desIn_r_58, u1_desIn_r_6, u1_desIn_r_60, 
       u1_desIn_r_61, u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_8, u1_key_r_10, u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_17, 
       u1_key_r_18, u1_key_r_19, u1_key_r_20, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, u1_key_r_3, u1_key_r_32, 
       u1_key_r_33, u1_key_r_34, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_46, u1_key_r_47, u1_key_r_48, 
       u1_key_r_5, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_uk_K_r0_11, u1_uk_K_r0_13, u1_uk_K_r0_17, u1_uk_K_r0_19, 
       u1_uk_K_r0_25, u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_55, u1_uk_K_r11_10, u1_uk_K_r11_17, u1_uk_K_r11_19, u1_uk_K_r11_24, u1_uk_K_r11_25, 
       u1_uk_K_r11_26, u1_uk_K_r11_33, u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, 
       u1_uk_K_r11_53, u1_uk_K_r11_54, u1_uk_K_r11_6, u1_uk_K_r14_10, u1_uk_K_r14_18, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r3_11, u1_uk_K_r3_19, 
       u1_uk_K_r8_10, u1_uk_K_r8_17, u1_uk_K_r8_27, u1_uk_K_r8_32, u1_uk_K_r8_39, u1_uk_K_r8_41, u1_uk_K_r8_48, u1_uk_K_r9_12, u1_uk_K_r9_15, 
       u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_25, u1_uk_K_r9_30, u1_uk_K_r9_33, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_49, 
       u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, 
       u1_uk_n110, u1_uk_n117, u1_uk_n1227, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1243, u1_uk_n1244, u1_uk_n1257, 
       u1_uk_n1259, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1269, u1_uk_n1270, u1_uk_n1274, u1_uk_n1277, u1_uk_n1278, 
       u1_uk_n129, u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1297, u1_uk_n1300, u1_uk_n1399, u1_uk_n1403, u1_uk_n1405, 
       u1_uk_n141, u1_uk_n1415, u1_uk_n1423, u1_uk_n1427, u1_uk_n1435, u1_uk_n1437, u1_uk_n145, u1_uk_n146, u1_uk_n147, 
       u1_uk_n148, u1_uk_n155, u1_uk_n161, u1_uk_n162, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1625, u1_uk_n1626, 
       u1_uk_n163, u1_uk_n1630, u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n164, u1_uk_n1642, u1_uk_n1643, u1_uk_n1649, 
       u1_uk_n1653, u1_uk_n1654, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1663, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, 
       u1_uk_n1673, u1_uk_n1676, u1_uk_n1682, u1_uk_n1683, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, 
       u1_uk_n1692, u1_uk_n1693, u1_uk_n1695, u1_uk_n1698, u1_uk_n1699, u1_uk_n17, u1_uk_n1703, u1_uk_n1705, u1_uk_n1707, 
       u1_uk_n1756, u1_uk_n1757, u1_uk_n1761, u1_uk_n1762, u1_uk_n1767, u1_uk_n1773, u1_uk_n1781, u1_uk_n1787, u1_uk_n1797, 
       u1_uk_n182, u1_uk_n187, u1_uk_n188, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, u1_uk_n209, 
       u1_uk_n213, u1_uk_n214, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n231, u1_uk_n238, u1_uk_n240, 
       u1_uk_n242, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, 
       u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n83, u1_uk_n93, 
       u1_uk_n94, u1_uk_n99, u2_FP_48, u2_FP_49, u2_FP_50, u2_FP_51, u2_FP_52, u2_FP_53, u2_K16_26, 
       u2_K3_13, u2_K3_15, u2_K3_16, u2_L14_14, u2_L14_25, u2_L14_3, u2_L14_8, u2_L1_16, u2_L1_17, 
       u2_L1_23, u2_L1_24, u2_L1_30, u2_L1_31, u2_L1_6, u2_L1_9, u2_R1_1, u2_R1_10, u2_R1_11, 
       u2_R1_12, u2_R1_13, u2_R1_2, u2_R1_3, u2_R1_32, u2_R1_4, u2_R1_5, u2_R1_8, u2_R1_9, 
       u2_uk_K_r14_45, u2_uk_K_r1_47, u2_uk_n10, u2_uk_n100, u2_uk_n1018, u2_uk_n102, u2_uk_n11, u2_uk_n1189, u2_uk_n1195, 
       u2_uk_n1200, u2_uk_n1209, u2_uk_n1216, u2_uk_n1226, u2_uk_n1282, u2_uk_n1285, u2_uk_n1287, u2_uk_n129, u2_uk_n1290, 
       u2_uk_n1293, u2_uk_n1295, u2_uk_n1301, u2_uk_n1302, u2_uk_n1306, u2_uk_n1310, u2_uk_n1317, u2_uk_n1318, u2_uk_n148, 
       u2_uk_n182, u2_uk_n187, u2_uk_n202, u2_uk_n208, u2_uk_n213, u2_uk_n214, u2_uk_n220, u2_uk_n222, u2_uk_n231, 
       u2_uk_n27, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n954, u2_uk_n955, u0_N452, u0_N454, u0_N459, u0_N462, u0_N468, u0_N469, u0_N474, u0_N479, u0_uk_n856, 
        u0_uk_n889, u0_uk_n998, u1_FP_16, u1_FP_24, u1_FP_30, u1_FP_6, u1_N0, u1_N1, u1_N12, 
        u1_N129, u1_N140, u1_N145, u1_N15, u1_N155, u1_N16, u1_N17, u1_N19, u1_N22, 
        u1_N23, u1_N25, u1_N27, u1_N289, u1_N29, u1_N293, u1_N296, u1_N30, u1_N300, 
        u1_N303, u1_N304, u1_N305, u1_N310, u1_N311, u1_N315, u1_N317, u1_N318, u1_N321, 
        u1_N323, u1_N325, u1_N328, u1_N33, u1_N330, u1_N332, u1_N335, u1_N336, u1_N337, 
        u1_N338, u1_N342, u1_N343, u1_N347, u1_N348, u1_N349, u1_N350, u1_N37, u1_N384, 
        u1_N385, u1_N392, u1_N393, u1_N396, u1_N400, u1_N401, u1_N403, u1_N406, u1_N409, 
        u1_N411, u1_N414, u1_N44, u1_N47, u1_N49, u1_N5, u1_N55, u1_N59, u1_N61, 
        u1_N8, u1_N9, u1_uk_n118, u1_uk_n128, u1_uk_n142, u1_uk_n250, u2_FP_14, u2_FP_25, u2_FP_3, 
        u2_FP_8, u2_N69, u2_N72, u2_N79, u2_N80, u2_N86, u2_N87, u2_N93, u2_N94 );
  input u0_K15_47, u0_L13_12, u0_L13_15, u0_L13_21, u0_L13_22, u0_L13_27, u0_L13_32, u0_L13_5, u0_L13_7, 
        u0_R13_1, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, 
        u0_R13_32, u0_key_r_18, u0_uk_K_r0_52, u0_uk_K_r13_2, u0_uk_K_r13_23, u0_uk_K_r13_35, u0_uk_K_r9_5, u0_uk_n10, u0_uk_n12, 
        u0_uk_n128, u0_uk_n13, u0_uk_n141, u0_uk_n155, u0_uk_n163, u0_uk_n17, u0_uk_n187, u0_uk_n21, u0_uk_n22, 
        u0_uk_n220, u0_uk_n23, u0_uk_n27, u0_uk_n3, u0_uk_n34, u0_uk_n39, u0_uk_n4, u0_uk_n40, u0_uk_n41, 
        u0_uk_n5, u0_uk_n9, u0_uk_n916, u0_uk_n93, u1_FP_40, u1_FP_41, u1_FP_42, u1_FP_43, u1_FP_44, 
        u1_FP_45, u1_L0_13, u1_L0_16, u1_L0_18, u1_L0_2, u1_L0_24, u1_L0_28, u1_L0_30, u1_L0_6, 
        u1_L11_1, u1_L11_10, u1_L11_13, u1_L11_17, u1_L11_18, u1_L11_2, u1_L11_20, u1_L11_23, u1_L11_26, 
        u1_L11_28, u1_L11_31, u1_L11_9, u1_L14_16, u1_L14_24, u1_L14_30, u1_L14_6, u1_L3_13, u1_L3_18, 
        u1_L3_2, u1_L3_28, u1_L8_13, u1_L8_16, u1_L8_17, u1_L8_18, u1_L8_2, u1_L8_23, u1_L8_24, 
        u1_L8_28, u1_L8_30, u1_L8_31, u1_L8_6, u1_L8_9, u1_L9_11, u1_L9_13, u1_L9_16, u1_L9_17, 
        u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_23, u1_L9_24, u1_L9_28, u1_L9_29, u1_L9_30, u1_L9_31, 
        u1_L9_4, u1_L9_6, u1_L9_9, u1_R0_10, u1_R0_11, u1_R0_12, u1_R0_13, u1_R0_4, u1_R0_5, 
        u1_R0_6, u1_R0_7, u1_R0_8, u1_R0_9, u1_R11_1, u1_R11_12, u1_R11_13, u1_R11_14, u1_R11_15, 
        u1_R11_16, u1_R11_17, u1_R11_2, u1_R11_3, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_6, u1_R11_7, 
        u1_R11_8, u1_R11_9, u1_R3_4, u1_R3_5, u1_R3_6, u1_R3_7, u1_R3_8, u1_R3_9, u1_R8_1, 
        u1_R8_10, u1_R8_11, u1_R8_12, u1_R8_13, u1_R8_2, u1_R8_3, u1_R8_32, u1_R8_4, u1_R8_5, 
        u1_R8_6, u1_R8_7, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_10, u1_R9_11, u1_R9_12, u1_R9_13, 
        u1_R9_2, u1_R9_20, u1_R9_21, u1_R9_22, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_3, u1_R9_32, 
        u1_R9_4, u1_R9_5, u1_R9_6, u1_R9_7, u1_R9_8, u1_R9_9, u1_desIn_r_10, u1_desIn_r_12, u1_desIn_r_13, 
        u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_2, u1_desIn_r_21, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_26, u1_desIn_r_29, u1_desIn_r_3, 
        u1_desIn_r_31, u1_desIn_r_36, u1_desIn_r_37, u1_desIn_r_39, u1_desIn_r_4, u1_desIn_r_40, u1_desIn_r_45, u1_desIn_r_46, u1_desIn_r_47, 
        u1_desIn_r_48, u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_53, u1_desIn_r_55, u1_desIn_r_57, u1_desIn_r_58, u1_desIn_r_6, u1_desIn_r_60, 
        u1_desIn_r_61, u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_8, u1_key_r_10, u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_17, 
        u1_key_r_18, u1_key_r_19, u1_key_r_20, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, u1_key_r_3, u1_key_r_32, 
        u1_key_r_33, u1_key_r_34, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_46, u1_key_r_47, u1_key_r_48, 
        u1_key_r_5, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_uk_K_r0_11, u1_uk_K_r0_13, u1_uk_K_r0_17, u1_uk_K_r0_19, 
        u1_uk_K_r0_25, u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_55, u1_uk_K_r11_10, u1_uk_K_r11_17, u1_uk_K_r11_19, u1_uk_K_r11_24, u1_uk_K_r11_25, 
        u1_uk_K_r11_26, u1_uk_K_r11_33, u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, 
        u1_uk_K_r11_53, u1_uk_K_r11_54, u1_uk_K_r11_6, u1_uk_K_r14_10, u1_uk_K_r14_18, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r3_11, u1_uk_K_r3_19, 
        u1_uk_K_r8_10, u1_uk_K_r8_17, u1_uk_K_r8_27, u1_uk_K_r8_32, u1_uk_K_r8_39, u1_uk_K_r8_41, u1_uk_K_r8_48, u1_uk_K_r9_12, u1_uk_K_r9_15, 
        u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_25, u1_uk_K_r9_30, u1_uk_K_r9_33, u1_uk_K_r9_4, u1_uk_K_r9_45, u1_uk_K_r9_49, 
        u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, 
        u1_uk_n110, u1_uk_n117, u1_uk_n1227, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1243, u1_uk_n1244, u1_uk_n1257, 
        u1_uk_n1259, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1269, u1_uk_n1270, u1_uk_n1274, u1_uk_n1277, u1_uk_n1278, 
        u1_uk_n129, u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1297, u1_uk_n1300, u1_uk_n1399, u1_uk_n1403, u1_uk_n1405, 
        u1_uk_n141, u1_uk_n1415, u1_uk_n1423, u1_uk_n1427, u1_uk_n1435, u1_uk_n1437, u1_uk_n145, u1_uk_n146, u1_uk_n147, 
        u1_uk_n148, u1_uk_n155, u1_uk_n161, u1_uk_n162, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1625, u1_uk_n1626, 
        u1_uk_n163, u1_uk_n1630, u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n164, u1_uk_n1642, u1_uk_n1643, u1_uk_n1649, 
        u1_uk_n1653, u1_uk_n1654, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1663, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, 
        u1_uk_n1673, u1_uk_n1676, u1_uk_n1682, u1_uk_n1683, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, 
        u1_uk_n1692, u1_uk_n1693, u1_uk_n1695, u1_uk_n1698, u1_uk_n1699, u1_uk_n17, u1_uk_n1703, u1_uk_n1705, u1_uk_n1707, 
        u1_uk_n1756, u1_uk_n1757, u1_uk_n1761, u1_uk_n1762, u1_uk_n1767, u1_uk_n1773, u1_uk_n1781, u1_uk_n1787, u1_uk_n1797, 
        u1_uk_n182, u1_uk_n187, u1_uk_n188, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, u1_uk_n209, 
        u1_uk_n213, u1_uk_n214, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n231, u1_uk_n238, u1_uk_n240, 
        u1_uk_n242, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, 
        u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n83, u1_uk_n93, 
        u1_uk_n94, u1_uk_n99, u2_FP_48, u2_FP_49, u2_FP_50, u2_FP_51, u2_FP_52, u2_FP_53, u2_K16_26, 
        u2_K3_13, u2_K3_15, u2_K3_16, u2_L14_14, u2_L14_25, u2_L14_3, u2_L14_8, u2_L1_16, u2_L1_17, 
        u2_L1_23, u2_L1_24, u2_L1_30, u2_L1_31, u2_L1_6, u2_L1_9, u2_R1_1, u2_R1_10, u2_R1_11, 
        u2_R1_12, u2_R1_13, u2_R1_2, u2_R1_3, u2_R1_32, u2_R1_4, u2_R1_5, u2_R1_8, u2_R1_9, 
        u2_uk_K_r14_45, u2_uk_K_r1_47, u2_uk_n10, u2_uk_n100, u2_uk_n1018, u2_uk_n102, u2_uk_n11, u2_uk_n1189, u2_uk_n1195, 
        u2_uk_n1200, u2_uk_n1209, u2_uk_n1216, u2_uk_n1226, u2_uk_n1282, u2_uk_n1285, u2_uk_n1287, u2_uk_n129, u2_uk_n1290, 
        u2_uk_n1293, u2_uk_n1295, u2_uk_n1301, u2_uk_n1302, u2_uk_n1306, u2_uk_n1310, u2_uk_n1317, u2_uk_n1318, u2_uk_n148, 
        u2_uk_n182, u2_uk_n187, u2_uk_n202, u2_uk_n208, u2_uk_n213, u2_uk_n214, u2_uk_n220, u2_uk_n222, u2_uk_n231, 
        u2_uk_n27, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n954, u2_uk_n955;
  output u0_N452, u0_N454, u0_N459, u0_N462, u0_N468, u0_N469, u0_N474, u0_N479, u0_uk_n856, 
        u0_uk_n889, u0_uk_n998, u1_FP_16, u1_FP_24, u1_FP_30, u1_FP_6, u1_N0, u1_N1, u1_N12, 
        u1_N129, u1_N140, u1_N145, u1_N15, u1_N155, u1_N16, u1_N17, u1_N19, u1_N22, 
        u1_N23, u1_N25, u1_N27, u1_N289, u1_N29, u1_N293, u1_N296, u1_N30, u1_N300, 
        u1_N303, u1_N304, u1_N305, u1_N310, u1_N311, u1_N315, u1_N317, u1_N318, u1_N321, 
        u1_N323, u1_N325, u1_N328, u1_N33, u1_N330, u1_N332, u1_N335, u1_N336, u1_N337, 
        u1_N338, u1_N342, u1_N343, u1_N347, u1_N348, u1_N349, u1_N350, u1_N37, u1_N384, 
        u1_N385, u1_N392, u1_N393, u1_N396, u1_N400, u1_N401, u1_N403, u1_N406, u1_N409, 
        u1_N411, u1_N414, u1_N44, u1_N47, u1_N49, u1_N5, u1_N55, u1_N59, u1_N61, 
        u1_N8, u1_N9, u1_uk_n118, u1_uk_n128, u1_uk_n142, u1_uk_n250, u2_FP_14, u2_FP_25, u2_FP_3, 
        u2_FP_8, u2_N69, u2_N72, u2_N79, u2_N80, u2_N86, u2_N87, u2_N93, u2_N94;
  wire u0_K15_37, u0_K15_38, u0_K15_39, u0_K15_40, u0_K15_41, u0_K15_42, u0_K15_43, u0_K15_44, u0_K15_45, 
       u0_K15_46, u0_K15_48, u0_out14_12, u0_out14_15, u0_out14_21, u0_out14_22, u0_out14_27, u0_out14_32, u0_out14_5, 
       u0_out14_7, u0_u14_X_37, u0_u14_X_38, u0_u14_X_39, u0_u14_X_40, u0_u14_X_41, u0_u14_X_42, u0_u14_X_43, u0_u14_X_44, 
       u0_u14_X_45, u0_u14_X_46, u0_u14_X_47, u0_u14_X_48, u0_u14_u6_n100, u0_u14_u6_n101, u0_u14_u6_n102, u0_u14_u6_n103, u0_u14_u6_n104, 
       u0_u14_u6_n105, u0_u14_u6_n106, u0_u14_u6_n107, u0_u14_u6_n108, u0_u14_u6_n109, u0_u14_u6_n110, u0_u14_u6_n111, u0_u14_u6_n112, u0_u14_u6_n113, 
       u0_u14_u6_n114, u0_u14_u6_n115, u0_u14_u6_n116, u0_u14_u6_n117, u0_u14_u6_n118, u0_u14_u6_n119, u0_u14_u6_n120, u0_u14_u6_n121, u0_u14_u6_n122, 
       u0_u14_u6_n123, u0_u14_u6_n124, u0_u14_u6_n125, u0_u14_u6_n126, u0_u14_u6_n127, u0_u14_u6_n128, u0_u14_u6_n129, u0_u14_u6_n130, u0_u14_u6_n131, 
       u0_u14_u6_n132, u0_u14_u6_n133, u0_u14_u6_n134, u0_u14_u6_n135, u0_u14_u6_n136, u0_u14_u6_n137, u0_u14_u6_n138, u0_u14_u6_n139, u0_u14_u6_n140, 
       u0_u14_u6_n141, u0_u14_u6_n142, u0_u14_u6_n143, u0_u14_u6_n144, u0_u14_u6_n145, u0_u14_u6_n146, u0_u14_u6_n147, u0_u14_u6_n148, u0_u14_u6_n149, 
       u0_u14_u6_n150, u0_u14_u6_n151, u0_u14_u6_n152, u0_u14_u6_n153, u0_u14_u6_n154, u0_u14_u6_n155, u0_u14_u6_n156, u0_u14_u6_n157, u0_u14_u6_n158, 
       u0_u14_u6_n159, u0_u14_u6_n160, u0_u14_u6_n161, u0_u14_u6_n162, u0_u14_u6_n163, u0_u14_u6_n164, u0_u14_u6_n165, u0_u14_u6_n166, u0_u14_u6_n167, 
       u0_u14_u6_n168, u0_u14_u6_n169, u0_u14_u6_n170, u0_u14_u6_n171, u0_u14_u6_n172, u0_u14_u6_n173, u0_u14_u6_n174, u0_u14_u6_n88, u0_u14_u6_n89, 
       u0_u14_u6_n90, u0_u14_u6_n91, u0_u14_u6_n92, u0_u14_u6_n93, u0_u14_u6_n94, u0_u14_u6_n95, u0_u14_u6_n96, u0_u14_u6_n97, u0_u14_u6_n98, 
       u0_u14_u6_n99, u0_u14_u7_n100, u0_u14_u7_n101, u0_u14_u7_n102, u0_u14_u7_n103, u0_u14_u7_n104, u0_u14_u7_n105, u0_u14_u7_n106, u0_u14_u7_n107, 
       u0_u14_u7_n108, u0_u14_u7_n109, u0_u14_u7_n110, u0_u14_u7_n111, u0_u14_u7_n112, u0_u14_u7_n113, u0_u14_u7_n114, u0_u14_u7_n115, u0_u14_u7_n116, 
       u0_u14_u7_n117, u0_u14_u7_n118, u0_u14_u7_n119, u0_u14_u7_n120, u0_u14_u7_n121, u0_u14_u7_n122, u0_u14_u7_n123, u0_u14_u7_n124, u0_u14_u7_n125, 
       u0_u14_u7_n126, u0_u14_u7_n127, u0_u14_u7_n128, u0_u14_u7_n129, u0_u14_u7_n130, u0_u14_u7_n131, u0_u14_u7_n132, u0_u14_u7_n133, u0_u14_u7_n134, 
       u0_u14_u7_n135, u0_u14_u7_n136, u0_u14_u7_n137, u0_u14_u7_n138, u0_u14_u7_n139, u0_u14_u7_n140, u0_u14_u7_n141, u0_u14_u7_n142, u0_u14_u7_n143, 
       u0_u14_u7_n144, u0_u14_u7_n145, u0_u14_u7_n146, u0_u14_u7_n147, u0_u14_u7_n148, u0_u14_u7_n149, u0_u14_u7_n150, u0_u14_u7_n151, u0_u14_u7_n152, 
       u0_u14_u7_n153, u0_u14_u7_n154, u0_u14_u7_n155, u0_u14_u7_n156, u0_u14_u7_n157, u0_u14_u7_n158, u0_u14_u7_n159, u0_u14_u7_n160, u0_u14_u7_n161, 
       u0_u14_u7_n162, u0_u14_u7_n163, u0_u14_u7_n164, u0_u14_u7_n165, u0_u14_u7_n166, u0_u14_u7_n167, u0_u14_u7_n168, u0_u14_u7_n169, u0_u14_u7_n170, 
       u0_u14_u7_n171, u0_u14_u7_n172, u0_u14_u7_n173, u0_u14_u7_n174, u0_u14_u7_n175, u0_u14_u7_n176, u0_u14_u7_n177, u0_u14_u7_n178, u0_u14_u7_n179, 
       u0_u14_u7_n180, u0_u14_u7_n91, u0_u14_u7_n92, u0_u14_u7_n93, u0_u14_u7_n94, u0_u14_u7_n95, u0_u14_u7_n96, u0_u14_u7_n97, u0_u14_u7_n98, 
       u0_u14_u7_n99, u0_uk_n914, u0_uk_n915, u1_K10_1, u1_K10_10, u1_K10_11, u1_K10_12, u1_K10_13, u1_K10_14, 
       u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_2, u1_K10_3, u1_K10_4, u1_K10_5, u1_K10_6, 
       u1_K10_7, u1_K10_8, u1_K10_9, u1_K11_1, u1_K11_10, u1_K11_11, u1_K11_12, u1_K11_13, u1_K11_14, 
       u1_K11_15, u1_K11_16, u1_K11_17, u1_K11_18, u1_K11_2, u1_K11_3, u1_K11_31, u1_K11_32, u1_K11_33, 
       u1_K11_34, u1_K11_35, u1_K11_36, u1_K11_4, u1_K11_5, u1_K11_6, u1_K11_7, u1_K11_8, u1_K11_9, 
       u1_K13_1, u1_K13_10, u1_K13_11, u1_K13_12, u1_K13_19, u1_K13_2, u1_K13_20, u1_K13_21, u1_K13_22, 
       u1_K13_23, u1_K13_24, u1_K13_3, u1_K13_4, u1_K13_5, u1_K13_6, u1_K13_7, u1_K13_8, u1_K13_9, 
       u1_K16_13, u1_K16_14, u1_K16_15, u1_K16_16, u1_K16_17, u1_K16_18, u1_K1_1, u1_K1_10, u1_K1_11, 
       u1_K1_12, u1_K1_13, u1_K1_14, u1_K1_15, u1_K1_16, u1_K1_17, u1_K1_18, u1_K1_19, u1_K1_2, 
       u1_K1_20, u1_K1_21, u1_K1_22, u1_K1_23, u1_K1_24, u1_K1_3, u1_K1_4, u1_K1_5, u1_K1_6, 
       u1_K1_7, u1_K1_8, u1_K1_9, u1_K2_10, u1_K2_11, u1_K2_12, u1_K2_13, u1_K2_14, u1_K2_15, 
       u1_K2_16, u1_K2_17, u1_K2_18, u1_K2_7, u1_K2_8, u1_K2_9, u1_K5_10, u1_K5_11, u1_K5_12, 
       u1_K5_7, u1_K5_8, u1_K5_9, u1_out0_1, u1_out0_10, u1_out0_13, u1_out0_16, u1_out0_17, u1_out0_18, 
       u1_out0_2, u1_out0_20, u1_out0_23, u1_out0_24, u1_out0_26, u1_out0_28, u1_out0_30, u1_out0_31, u1_out0_6, 
       u1_out0_9, u1_out10_11, u1_out10_13, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_23, 
       u1_out10_24, u1_out10_28, u1_out10_29, u1_out10_30, u1_out10_31, u1_out10_4, u1_out10_6, u1_out10_9, u1_out12_1, 
       u1_out12_10, u1_out12_13, u1_out12_17, u1_out12_18, u1_out12_2, u1_out12_20, u1_out12_23, u1_out12_26, u1_out12_28, 
       u1_out12_31, u1_out12_9, u1_out15_16, u1_out15_24, u1_out15_30, u1_out15_6, u1_out1_13, u1_out1_16, u1_out1_18, 
       u1_out1_2, u1_out1_24, u1_out1_28, u1_out1_30, u1_out1_6, u1_out4_13, u1_out4_18, u1_out4_2, u1_out4_28, 
       u1_out9_13, u1_out9_16, u1_out9_17, u1_out9_18, u1_out9_2, u1_out9_23, u1_out9_24, u1_out9_28, u1_out9_30, 
       u1_out9_31, u1_out9_6, u1_out9_9, u1_u0_X_1, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_13, u1_u0_X_14, 
       u1_u0_X_15, u1_u0_X_16, u1_u0_X_17, u1_u0_X_18, u1_u0_X_19, u1_u0_X_2, u1_u0_X_20, u1_u0_X_21, u1_u0_X_22, 
       u1_u0_X_23, u1_u0_X_24, u1_u0_X_3, u1_u0_X_4, u1_u0_X_5, u1_u0_X_6, u1_u0_X_7, u1_u0_X_8, u1_u0_X_9, 
       u1_u0_u0_n100, u1_u0_u0_n101, u1_u0_u0_n102, u1_u0_u0_n103, u1_u0_u0_n104, u1_u0_u0_n105, u1_u0_u0_n106, u1_u0_u0_n107, u1_u0_u0_n108, 
       u1_u0_u0_n109, u1_u0_u0_n110, u1_u0_u0_n111, u1_u0_u0_n112, u1_u0_u0_n113, u1_u0_u0_n114, u1_u0_u0_n115, u1_u0_u0_n116, u1_u0_u0_n117, 
       u1_u0_u0_n118, u1_u0_u0_n119, u1_u0_u0_n120, u1_u0_u0_n121, u1_u0_u0_n122, u1_u0_u0_n123, u1_u0_u0_n124, u1_u0_u0_n125, u1_u0_u0_n126, 
       u1_u0_u0_n127, u1_u0_u0_n128, u1_u0_u0_n129, u1_u0_u0_n130, u1_u0_u0_n131, u1_u0_u0_n132, u1_u0_u0_n133, u1_u0_u0_n134, u1_u0_u0_n135, 
       u1_u0_u0_n136, u1_u0_u0_n137, u1_u0_u0_n138, u1_u0_u0_n139, u1_u0_u0_n140, u1_u0_u0_n141, u1_u0_u0_n142, u1_u0_u0_n143, u1_u0_u0_n144, 
       u1_u0_u0_n145, u1_u0_u0_n146, u1_u0_u0_n147, u1_u0_u0_n148, u1_u0_u0_n149, u1_u0_u0_n150, u1_u0_u0_n151, u1_u0_u0_n152, u1_u0_u0_n153, 
       u1_u0_u0_n154, u1_u0_u0_n155, u1_u0_u0_n156, u1_u0_u0_n157, u1_u0_u0_n158, u1_u0_u0_n159, u1_u0_u0_n160, u1_u0_u0_n161, u1_u0_u0_n162, 
       u1_u0_u0_n163, u1_u0_u0_n164, u1_u0_u0_n165, u1_u0_u0_n166, u1_u0_u0_n167, u1_u0_u0_n168, u1_u0_u0_n169, u1_u0_u0_n170, u1_u0_u0_n171, 
       u1_u0_u0_n172, u1_u0_u0_n173, u1_u0_u0_n174, u1_u0_u0_n88, u1_u0_u0_n89, u1_u0_u0_n90, u1_u0_u0_n91, u1_u0_u0_n92, u1_u0_u0_n93, 
       u1_u0_u0_n94, u1_u0_u0_n95, u1_u0_u0_n96, u1_u0_u0_n97, u1_u0_u0_n98, u1_u0_u0_n99, u1_u0_u1_n100, u1_u0_u1_n101, u1_u0_u1_n102, 
       u1_u0_u1_n103, u1_u0_u1_n104, u1_u0_u1_n105, u1_u0_u1_n106, u1_u0_u1_n107, u1_u0_u1_n108, u1_u0_u1_n109, u1_u0_u1_n110, u1_u0_u1_n111, 
       u1_u0_u1_n112, u1_u0_u1_n113, u1_u0_u1_n114, u1_u0_u1_n115, u1_u0_u1_n116, u1_u0_u1_n117, u1_u0_u1_n118, u1_u0_u1_n119, u1_u0_u1_n120, 
       u1_u0_u1_n121, u1_u0_u1_n122, u1_u0_u1_n123, u1_u0_u1_n124, u1_u0_u1_n125, u1_u0_u1_n126, u1_u0_u1_n127, u1_u0_u1_n128, u1_u0_u1_n129, 
       u1_u0_u1_n130, u1_u0_u1_n131, u1_u0_u1_n132, u1_u0_u1_n133, u1_u0_u1_n134, u1_u0_u1_n135, u1_u0_u1_n136, u1_u0_u1_n137, u1_u0_u1_n138, 
       u1_u0_u1_n139, u1_u0_u1_n140, u1_u0_u1_n141, u1_u0_u1_n142, u1_u0_u1_n143, u1_u0_u1_n144, u1_u0_u1_n145, u1_u0_u1_n146, u1_u0_u1_n147, 
       u1_u0_u1_n148, u1_u0_u1_n149, u1_u0_u1_n150, u1_u0_u1_n151, u1_u0_u1_n152, u1_u0_u1_n153, u1_u0_u1_n154, u1_u0_u1_n155, u1_u0_u1_n156, 
       u1_u0_u1_n157, u1_u0_u1_n158, u1_u0_u1_n159, u1_u0_u1_n160, u1_u0_u1_n161, u1_u0_u1_n162, u1_u0_u1_n163, u1_u0_u1_n164, u1_u0_u1_n165, 
       u1_u0_u1_n166, u1_u0_u1_n167, u1_u0_u1_n168, u1_u0_u1_n169, u1_u0_u1_n170, u1_u0_u1_n171, u1_u0_u1_n172, u1_u0_u1_n173, u1_u0_u1_n174, 
       u1_u0_u1_n175, u1_u0_u1_n176, u1_u0_u1_n177, u1_u0_u1_n178, u1_u0_u1_n179, u1_u0_u1_n180, u1_u0_u1_n181, u1_u0_u1_n182, u1_u0_u1_n183, 
       u1_u0_u1_n184, u1_u0_u1_n185, u1_u0_u1_n186, u1_u0_u1_n187, u1_u0_u1_n188, u1_u0_u1_n95, u1_u0_u1_n96, u1_u0_u1_n97, u1_u0_u1_n98, 
       u1_u0_u1_n99, u1_u0_u2_n100, u1_u0_u2_n101, u1_u0_u2_n102, u1_u0_u2_n103, u1_u0_u2_n104, u1_u0_u2_n105, u1_u0_u2_n106, u1_u0_u2_n107, 
       u1_u0_u2_n108, u1_u0_u2_n109, u1_u0_u2_n110, u1_u0_u2_n111, u1_u0_u2_n112, u1_u0_u2_n113, u1_u0_u2_n114, u1_u0_u2_n115, u1_u0_u2_n116, 
       u1_u0_u2_n117, u1_u0_u2_n118, u1_u0_u2_n119, u1_u0_u2_n120, u1_u0_u2_n121, u1_u0_u2_n122, u1_u0_u2_n123, u1_u0_u2_n124, u1_u0_u2_n125, 
       u1_u0_u2_n126, u1_u0_u2_n127, u1_u0_u2_n128, u1_u0_u2_n129, u1_u0_u2_n130, u1_u0_u2_n131, u1_u0_u2_n132, u1_u0_u2_n133, u1_u0_u2_n134, 
       u1_u0_u2_n135, u1_u0_u2_n136, u1_u0_u2_n137, u1_u0_u2_n138, u1_u0_u2_n139, u1_u0_u2_n140, u1_u0_u2_n141, u1_u0_u2_n142, u1_u0_u2_n143, 
       u1_u0_u2_n144, u1_u0_u2_n145, u1_u0_u2_n146, u1_u0_u2_n147, u1_u0_u2_n148, u1_u0_u2_n149, u1_u0_u2_n150, u1_u0_u2_n151, u1_u0_u2_n152, 
       u1_u0_u2_n153, u1_u0_u2_n154, u1_u0_u2_n155, u1_u0_u2_n156, u1_u0_u2_n157, u1_u0_u2_n158, u1_u0_u2_n159, u1_u0_u2_n160, u1_u0_u2_n161, 
       u1_u0_u2_n162, u1_u0_u2_n163, u1_u0_u2_n164, u1_u0_u2_n165, u1_u0_u2_n166, u1_u0_u2_n167, u1_u0_u2_n168, u1_u0_u2_n169, u1_u0_u2_n170, 
       u1_u0_u2_n171, u1_u0_u2_n172, u1_u0_u2_n173, u1_u0_u2_n174, u1_u0_u2_n175, u1_u0_u2_n176, u1_u0_u2_n177, u1_u0_u2_n178, u1_u0_u2_n179, 
       u1_u0_u2_n180, u1_u0_u2_n181, u1_u0_u2_n182, u1_u0_u2_n183, u1_u0_u2_n184, u1_u0_u2_n185, u1_u0_u2_n186, u1_u0_u2_n187, u1_u0_u2_n188, 
       u1_u0_u2_n95, u1_u0_u2_n96, u1_u0_u2_n97, u1_u0_u2_n98, u1_u0_u2_n99, u1_u0_u3_n100, u1_u0_u3_n101, u1_u0_u3_n102, u1_u0_u3_n103, 
       u1_u0_u3_n104, u1_u0_u3_n105, u1_u0_u3_n106, u1_u0_u3_n107, u1_u0_u3_n108, u1_u0_u3_n109, u1_u0_u3_n110, u1_u0_u3_n111, u1_u0_u3_n112, 
       u1_u0_u3_n113, u1_u0_u3_n114, u1_u0_u3_n115, u1_u0_u3_n116, u1_u0_u3_n117, u1_u0_u3_n118, u1_u0_u3_n119, u1_u0_u3_n120, u1_u0_u3_n121, 
       u1_u0_u3_n122, u1_u0_u3_n123, u1_u0_u3_n124, u1_u0_u3_n125, u1_u0_u3_n126, u1_u0_u3_n127, u1_u0_u3_n128, u1_u0_u3_n129, u1_u0_u3_n130, 
       u1_u0_u3_n131, u1_u0_u3_n132, u1_u0_u3_n133, u1_u0_u3_n134, u1_u0_u3_n135, u1_u0_u3_n136, u1_u0_u3_n137, u1_u0_u3_n138, u1_u0_u3_n139, 
       u1_u0_u3_n140, u1_u0_u3_n141, u1_u0_u3_n142, u1_u0_u3_n143, u1_u0_u3_n144, u1_u0_u3_n145, u1_u0_u3_n146, u1_u0_u3_n147, u1_u0_u3_n148, 
       u1_u0_u3_n149, u1_u0_u3_n150, u1_u0_u3_n151, u1_u0_u3_n152, u1_u0_u3_n153, u1_u0_u3_n154, u1_u0_u3_n155, u1_u0_u3_n156, u1_u0_u3_n157, 
       u1_u0_u3_n158, u1_u0_u3_n159, u1_u0_u3_n160, u1_u0_u3_n161, u1_u0_u3_n162, u1_u0_u3_n163, u1_u0_u3_n164, u1_u0_u3_n165, u1_u0_u3_n166, 
       u1_u0_u3_n167, u1_u0_u3_n168, u1_u0_u3_n169, u1_u0_u3_n170, u1_u0_u3_n171, u1_u0_u3_n172, u1_u0_u3_n173, u1_u0_u3_n174, u1_u0_u3_n175, 
       u1_u0_u3_n176, u1_u0_u3_n177, u1_u0_u3_n178, u1_u0_u3_n179, u1_u0_u3_n180, u1_u0_u3_n181, u1_u0_u3_n182, u1_u0_u3_n183, u1_u0_u3_n184, 
       u1_u0_u3_n185, u1_u0_u3_n186, u1_u0_u3_n94, u1_u0_u3_n95, u1_u0_u3_n96, u1_u0_u3_n97, u1_u0_u3_n98, u1_u0_u3_n99, u1_u10_X_1, 
       u1_u10_X_10, u1_u10_X_11, u1_u10_X_12, u1_u10_X_13, u1_u10_X_14, u1_u10_X_15, u1_u10_X_16, u1_u10_X_17, u1_u10_X_18, 
       u1_u10_X_2, u1_u10_X_3, u1_u10_X_31, u1_u10_X_32, u1_u10_X_33, u1_u10_X_34, u1_u10_X_35, u1_u10_X_36, u1_u10_X_4, 
       u1_u10_X_5, u1_u10_X_6, u1_u10_X_7, u1_u10_X_8, u1_u10_X_9, u1_u10_u0_n100, u1_u10_u0_n101, u1_u10_u0_n102, u1_u10_u0_n103, 
       u1_u10_u0_n104, u1_u10_u0_n105, u1_u10_u0_n106, u1_u10_u0_n107, u1_u10_u0_n108, u1_u10_u0_n109, u1_u10_u0_n110, u1_u10_u0_n111, u1_u10_u0_n112, 
       u1_u10_u0_n113, u1_u10_u0_n114, u1_u10_u0_n115, u1_u10_u0_n116, u1_u10_u0_n117, u1_u10_u0_n118, u1_u10_u0_n119, u1_u10_u0_n120, u1_u10_u0_n121, 
       u1_u10_u0_n122, u1_u10_u0_n123, u1_u10_u0_n124, u1_u10_u0_n125, u1_u10_u0_n126, u1_u10_u0_n127, u1_u10_u0_n128, u1_u10_u0_n129, u1_u10_u0_n130, 
       u1_u10_u0_n131, u1_u10_u0_n132, u1_u10_u0_n133, u1_u10_u0_n134, u1_u10_u0_n135, u1_u10_u0_n136, u1_u10_u0_n137, u1_u10_u0_n138, u1_u10_u0_n139, 
       u1_u10_u0_n140, u1_u10_u0_n141, u1_u10_u0_n142, u1_u10_u0_n143, u1_u10_u0_n144, u1_u10_u0_n145, u1_u10_u0_n146, u1_u10_u0_n147, u1_u10_u0_n148, 
       u1_u10_u0_n149, u1_u10_u0_n150, u1_u10_u0_n151, u1_u10_u0_n152, u1_u10_u0_n153, u1_u10_u0_n154, u1_u10_u0_n155, u1_u10_u0_n156, u1_u10_u0_n157, 
       u1_u10_u0_n158, u1_u10_u0_n159, u1_u10_u0_n160, u1_u10_u0_n161, u1_u10_u0_n162, u1_u10_u0_n163, u1_u10_u0_n164, u1_u10_u0_n165, u1_u10_u0_n166, 
       u1_u10_u0_n167, u1_u10_u0_n168, u1_u10_u0_n169, u1_u10_u0_n170, u1_u10_u0_n171, u1_u10_u0_n172, u1_u10_u0_n173, u1_u10_u0_n174, u1_u10_u0_n88, 
       u1_u10_u0_n89, u1_u10_u0_n90, u1_u10_u0_n91, u1_u10_u0_n92, u1_u10_u0_n93, u1_u10_u0_n94, u1_u10_u0_n95, u1_u10_u0_n96, u1_u10_u0_n97, 
       u1_u10_u0_n98, u1_u10_u0_n99, u1_u10_u1_n100, u1_u10_u1_n101, u1_u10_u1_n102, u1_u10_u1_n103, u1_u10_u1_n104, u1_u10_u1_n105, u1_u10_u1_n106, 
       u1_u10_u1_n107, u1_u10_u1_n108, u1_u10_u1_n109, u1_u10_u1_n110, u1_u10_u1_n111, u1_u10_u1_n112, u1_u10_u1_n113, u1_u10_u1_n114, u1_u10_u1_n115, 
       u1_u10_u1_n116, u1_u10_u1_n117, u1_u10_u1_n118, u1_u10_u1_n119, u1_u10_u1_n120, u1_u10_u1_n121, u1_u10_u1_n122, u1_u10_u1_n123, u1_u10_u1_n124, 
       u1_u10_u1_n125, u1_u10_u1_n126, u1_u10_u1_n127, u1_u10_u1_n128, u1_u10_u1_n129, u1_u10_u1_n130, u1_u10_u1_n131, u1_u10_u1_n132, u1_u10_u1_n133, 
       u1_u10_u1_n134, u1_u10_u1_n135, u1_u10_u1_n136, u1_u10_u1_n137, u1_u10_u1_n138, u1_u10_u1_n139, u1_u10_u1_n140, u1_u10_u1_n141, u1_u10_u1_n142, 
       u1_u10_u1_n143, u1_u10_u1_n144, u1_u10_u1_n145, u1_u10_u1_n146, u1_u10_u1_n147, u1_u10_u1_n148, u1_u10_u1_n149, u1_u10_u1_n150, u1_u10_u1_n151, 
       u1_u10_u1_n152, u1_u10_u1_n153, u1_u10_u1_n154, u1_u10_u1_n155, u1_u10_u1_n156, u1_u10_u1_n157, u1_u10_u1_n158, u1_u10_u1_n159, u1_u10_u1_n160, 
       u1_u10_u1_n161, u1_u10_u1_n162, u1_u10_u1_n163, u1_u10_u1_n164, u1_u10_u1_n165, u1_u10_u1_n166, u1_u10_u1_n167, u1_u10_u1_n168, u1_u10_u1_n169, 
       u1_u10_u1_n170, u1_u10_u1_n171, u1_u10_u1_n172, u1_u10_u1_n173, u1_u10_u1_n174, u1_u10_u1_n175, u1_u10_u1_n176, u1_u10_u1_n177, u1_u10_u1_n178, 
       u1_u10_u1_n179, u1_u10_u1_n180, u1_u10_u1_n181, u1_u10_u1_n182, u1_u10_u1_n183, u1_u10_u1_n184, u1_u10_u1_n185, u1_u10_u1_n186, u1_u10_u1_n187, 
       u1_u10_u1_n188, u1_u10_u1_n95, u1_u10_u1_n96, u1_u10_u1_n97, u1_u10_u1_n98, u1_u10_u1_n99, u1_u10_u2_n100, u1_u10_u2_n101, u1_u10_u2_n102, 
       u1_u10_u2_n103, u1_u10_u2_n104, u1_u10_u2_n105, u1_u10_u2_n106, u1_u10_u2_n107, u1_u10_u2_n108, u1_u10_u2_n109, u1_u10_u2_n110, u1_u10_u2_n111, 
       u1_u10_u2_n112, u1_u10_u2_n113, u1_u10_u2_n114, u1_u10_u2_n115, u1_u10_u2_n116, u1_u10_u2_n117, u1_u10_u2_n118, u1_u10_u2_n119, u1_u10_u2_n120, 
       u1_u10_u2_n121, u1_u10_u2_n122, u1_u10_u2_n123, u1_u10_u2_n124, u1_u10_u2_n125, u1_u10_u2_n126, u1_u10_u2_n127, u1_u10_u2_n128, u1_u10_u2_n129, 
       u1_u10_u2_n130, u1_u10_u2_n131, u1_u10_u2_n132, u1_u10_u2_n133, u1_u10_u2_n134, u1_u10_u2_n135, u1_u10_u2_n136, u1_u10_u2_n137, u1_u10_u2_n138, 
       u1_u10_u2_n139, u1_u10_u2_n140, u1_u10_u2_n141, u1_u10_u2_n142, u1_u10_u2_n143, u1_u10_u2_n144, u1_u10_u2_n145, u1_u10_u2_n146, u1_u10_u2_n147, 
       u1_u10_u2_n148, u1_u10_u2_n149, u1_u10_u2_n150, u1_u10_u2_n151, u1_u10_u2_n152, u1_u10_u2_n153, u1_u10_u2_n154, u1_u10_u2_n155, u1_u10_u2_n156, 
       u1_u10_u2_n157, u1_u10_u2_n158, u1_u10_u2_n159, u1_u10_u2_n160, u1_u10_u2_n161, u1_u10_u2_n162, u1_u10_u2_n163, u1_u10_u2_n164, u1_u10_u2_n165, 
       u1_u10_u2_n166, u1_u10_u2_n167, u1_u10_u2_n168, u1_u10_u2_n169, u1_u10_u2_n170, u1_u10_u2_n171, u1_u10_u2_n172, u1_u10_u2_n173, u1_u10_u2_n174, 
       u1_u10_u2_n175, u1_u10_u2_n176, u1_u10_u2_n177, u1_u10_u2_n178, u1_u10_u2_n179, u1_u10_u2_n180, u1_u10_u2_n181, u1_u10_u2_n182, u1_u10_u2_n183, 
       u1_u10_u2_n184, u1_u10_u2_n185, u1_u10_u2_n186, u1_u10_u2_n187, u1_u10_u2_n188, u1_u10_u2_n95, u1_u10_u2_n96, u1_u10_u2_n97, u1_u10_u2_n98, 
       u1_u10_u2_n99, u1_u10_u5_n100, u1_u10_u5_n101, u1_u10_u5_n102, u1_u10_u5_n103, u1_u10_u5_n104, u1_u10_u5_n105, u1_u10_u5_n106, u1_u10_u5_n107, 
       u1_u10_u5_n108, u1_u10_u5_n109, u1_u10_u5_n110, u1_u10_u5_n111, u1_u10_u5_n112, u1_u10_u5_n113, u1_u10_u5_n114, u1_u10_u5_n115, u1_u10_u5_n116, 
       u1_u10_u5_n117, u1_u10_u5_n118, u1_u10_u5_n119, u1_u10_u5_n120, u1_u10_u5_n121, u1_u10_u5_n122, u1_u10_u5_n123, u1_u10_u5_n124, u1_u10_u5_n125, 
       u1_u10_u5_n126, u1_u10_u5_n127, u1_u10_u5_n128, u1_u10_u5_n129, u1_u10_u5_n130, u1_u10_u5_n131, u1_u10_u5_n132, u1_u10_u5_n133, u1_u10_u5_n134, 
       u1_u10_u5_n135, u1_u10_u5_n136, u1_u10_u5_n137, u1_u10_u5_n138, u1_u10_u5_n139, u1_u10_u5_n140, u1_u10_u5_n141, u1_u10_u5_n142, u1_u10_u5_n143, 
       u1_u10_u5_n144, u1_u10_u5_n145, u1_u10_u5_n146, u1_u10_u5_n147, u1_u10_u5_n148, u1_u10_u5_n149, u1_u10_u5_n150, u1_u10_u5_n151, u1_u10_u5_n152, 
       u1_u10_u5_n153, u1_u10_u5_n154, u1_u10_u5_n155, u1_u10_u5_n156, u1_u10_u5_n157, u1_u10_u5_n158, u1_u10_u5_n159, u1_u10_u5_n160, u1_u10_u5_n161, 
       u1_u10_u5_n162, u1_u10_u5_n163, u1_u10_u5_n164, u1_u10_u5_n165, u1_u10_u5_n166, u1_u10_u5_n167, u1_u10_u5_n168, u1_u10_u5_n169, u1_u10_u5_n170, 
       u1_u10_u5_n171, u1_u10_u5_n172, u1_u10_u5_n173, u1_u10_u5_n174, u1_u10_u5_n175, u1_u10_u5_n176, u1_u10_u5_n177, u1_u10_u5_n178, u1_u10_u5_n179, 
       u1_u10_u5_n180, u1_u10_u5_n181, u1_u10_u5_n182, u1_u10_u5_n183, u1_u10_u5_n184, u1_u10_u5_n185, u1_u10_u5_n186, u1_u10_u5_n187, u1_u10_u5_n188, 
       u1_u10_u5_n189, u1_u10_u5_n190, u1_u10_u5_n191, u1_u10_u5_n192, u1_u10_u5_n193, u1_u10_u5_n194, u1_u10_u5_n195, u1_u10_u5_n196, u1_u10_u5_n99, 
       u1_u12_X_1, u1_u12_X_10, u1_u12_X_11, u1_u12_X_12, u1_u12_X_19, u1_u12_X_2, u1_u12_X_20, u1_u12_X_21, u1_u12_X_22, 
       u1_u12_X_23, u1_u12_X_24, u1_u12_X_3, u1_u12_X_4, u1_u12_X_5, u1_u12_X_6, u1_u12_X_7, u1_u12_X_8, u1_u12_X_9, 
       u1_u12_u0_n100, u1_u12_u0_n101, u1_u12_u0_n102, u1_u12_u0_n103, u1_u12_u0_n104, u1_u12_u0_n105, u1_u12_u0_n106, u1_u12_u0_n107, u1_u12_u0_n108, 
       u1_u12_u0_n109, u1_u12_u0_n110, u1_u12_u0_n111, u1_u12_u0_n112, u1_u12_u0_n113, u1_u12_u0_n114, u1_u12_u0_n115, u1_u12_u0_n116, u1_u12_u0_n117, 
       u1_u12_u0_n118, u1_u12_u0_n119, u1_u12_u0_n120, u1_u12_u0_n121, u1_u12_u0_n122, u1_u12_u0_n123, u1_u12_u0_n124, u1_u12_u0_n125, u1_u12_u0_n126, 
       u1_u12_u0_n127, u1_u12_u0_n128, u1_u12_u0_n129, u1_u12_u0_n130, u1_u12_u0_n131, u1_u12_u0_n132, u1_u12_u0_n133, u1_u12_u0_n134, u1_u12_u0_n135, 
       u1_u12_u0_n136, u1_u12_u0_n137, u1_u12_u0_n138, u1_u12_u0_n139, u1_u12_u0_n140, u1_u12_u0_n141, u1_u12_u0_n142, u1_u12_u0_n143, u1_u12_u0_n144, 
       u1_u12_u0_n145, u1_u12_u0_n146, u1_u12_u0_n147, u1_u12_u0_n148, u1_u12_u0_n149, u1_u12_u0_n150, u1_u12_u0_n151, u1_u12_u0_n152, u1_u12_u0_n153, 
       u1_u12_u0_n154, u1_u12_u0_n155, u1_u12_u0_n156, u1_u12_u0_n157, u1_u12_u0_n158, u1_u12_u0_n159, u1_u12_u0_n160, u1_u12_u0_n161, u1_u12_u0_n162, 
       u1_u12_u0_n163, u1_u12_u0_n164, u1_u12_u0_n165, u1_u12_u0_n166, u1_u12_u0_n167, u1_u12_u0_n168, u1_u12_u0_n169, u1_u12_u0_n170, u1_u12_u0_n171, 
       u1_u12_u0_n172, u1_u12_u0_n173, u1_u12_u0_n174, u1_u12_u0_n88, u1_u12_u0_n89, u1_u12_u0_n90, u1_u12_u0_n91, u1_u12_u0_n92, u1_u12_u0_n93, 
       u1_u12_u0_n94, u1_u12_u0_n95, u1_u12_u0_n96, u1_u12_u0_n97, u1_u12_u0_n98, u1_u12_u0_n99, u1_u12_u1_n100, u1_u12_u1_n101, u1_u12_u1_n102, 
       u1_u12_u1_n103, u1_u12_u1_n104, u1_u12_u1_n105, u1_u12_u1_n106, u1_u12_u1_n107, u1_u12_u1_n108, u1_u12_u1_n109, u1_u12_u1_n110, u1_u12_u1_n111, 
       u1_u12_u1_n112, u1_u12_u1_n113, u1_u12_u1_n114, u1_u12_u1_n115, u1_u12_u1_n116, u1_u12_u1_n117, u1_u12_u1_n118, u1_u12_u1_n119, u1_u12_u1_n120, 
       u1_u12_u1_n121, u1_u12_u1_n122, u1_u12_u1_n123, u1_u12_u1_n124, u1_u12_u1_n125, u1_u12_u1_n126, u1_u12_u1_n127, u1_u12_u1_n128, u1_u12_u1_n129, 
       u1_u12_u1_n130, u1_u12_u1_n131, u1_u12_u1_n132, u1_u12_u1_n133, u1_u12_u1_n134, u1_u12_u1_n135, u1_u12_u1_n136, u1_u12_u1_n137, u1_u12_u1_n138, 
       u1_u12_u1_n139, u1_u12_u1_n140, u1_u12_u1_n141, u1_u12_u1_n142, u1_u12_u1_n143, u1_u12_u1_n144, u1_u12_u1_n145, u1_u12_u1_n146, u1_u12_u1_n147, 
       u1_u12_u1_n148, u1_u12_u1_n149, u1_u12_u1_n150, u1_u12_u1_n151, u1_u12_u1_n152, u1_u12_u1_n153, u1_u12_u1_n154, u1_u12_u1_n155, u1_u12_u1_n156, 
       u1_u12_u1_n157, u1_u12_u1_n158, u1_u12_u1_n159, u1_u12_u1_n160, u1_u12_u1_n161, u1_u12_u1_n162, u1_u12_u1_n163, u1_u12_u1_n164, u1_u12_u1_n165, 
       u1_u12_u1_n166, u1_u12_u1_n167, u1_u12_u1_n168, u1_u12_u1_n169, u1_u12_u1_n170, u1_u12_u1_n171, u1_u12_u1_n172, u1_u12_u1_n173, u1_u12_u1_n174, 
       u1_u12_u1_n175, u1_u12_u1_n176, u1_u12_u1_n177, u1_u12_u1_n178, u1_u12_u1_n179, u1_u12_u1_n180, u1_u12_u1_n181, u1_u12_u1_n182, u1_u12_u1_n183, 
       u1_u12_u1_n184, u1_u12_u1_n185, u1_u12_u1_n186, u1_u12_u1_n187, u1_u12_u1_n188, u1_u12_u1_n95, u1_u12_u1_n96, u1_u12_u1_n97, u1_u12_u1_n98, 
       u1_u12_u1_n99, u1_u12_u3_n100, u1_u12_u3_n101, u1_u12_u3_n102, u1_u12_u3_n103, u1_u12_u3_n104, u1_u12_u3_n105, u1_u12_u3_n106, u1_u12_u3_n107, 
       u1_u12_u3_n108, u1_u12_u3_n109, u1_u12_u3_n110, u1_u12_u3_n111, u1_u12_u3_n112, u1_u12_u3_n113, u1_u12_u3_n114, u1_u12_u3_n115, u1_u12_u3_n116, 
       u1_u12_u3_n117, u1_u12_u3_n118, u1_u12_u3_n119, u1_u12_u3_n120, u1_u12_u3_n121, u1_u12_u3_n122, u1_u12_u3_n123, u1_u12_u3_n124, u1_u12_u3_n125, 
       u1_u12_u3_n126, u1_u12_u3_n127, u1_u12_u3_n128, u1_u12_u3_n129, u1_u12_u3_n130, u1_u12_u3_n131, u1_u12_u3_n132, u1_u12_u3_n133, u1_u12_u3_n134, 
       u1_u12_u3_n135, u1_u12_u3_n136, u1_u12_u3_n137, u1_u12_u3_n138, u1_u12_u3_n139, u1_u12_u3_n140, u1_u12_u3_n141, u1_u12_u3_n142, u1_u12_u3_n143, 
       u1_u12_u3_n144, u1_u12_u3_n145, u1_u12_u3_n146, u1_u12_u3_n147, u1_u12_u3_n148, u1_u12_u3_n149, u1_u12_u3_n150, u1_u12_u3_n151, u1_u12_u3_n152, 
       u1_u12_u3_n153, u1_u12_u3_n154, u1_u12_u3_n155, u1_u12_u3_n156, u1_u12_u3_n157, u1_u12_u3_n158, u1_u12_u3_n159, u1_u12_u3_n160, u1_u12_u3_n161, 
       u1_u12_u3_n162, u1_u12_u3_n163, u1_u12_u3_n164, u1_u12_u3_n165, u1_u12_u3_n166, u1_u12_u3_n167, u1_u12_u3_n168, u1_u12_u3_n169, u1_u12_u3_n170, 
       u1_u12_u3_n171, u1_u12_u3_n172, u1_u12_u3_n173, u1_u12_u3_n174, u1_u12_u3_n175, u1_u12_u3_n176, u1_u12_u3_n177, u1_u12_u3_n178, u1_u12_u3_n179, 
       u1_u12_u3_n180, u1_u12_u3_n181, u1_u12_u3_n182, u1_u12_u3_n183, u1_u12_u3_n184, u1_u12_u3_n185, u1_u12_u3_n186, u1_u12_u3_n94, u1_u12_u3_n95, 
       u1_u12_u3_n96, u1_u12_u3_n97, u1_u12_u3_n98, u1_u12_u3_n99, u1_u15_X_13, u1_u15_X_14, u1_u15_X_15, u1_u15_X_16, u1_u15_X_17, 
       u1_u15_X_18, u1_u15_u2_n100, u1_u15_u2_n101, u1_u15_u2_n102, u1_u15_u2_n103, u1_u15_u2_n104, u1_u15_u2_n105, u1_u15_u2_n106, u1_u15_u2_n107, 
       u1_u15_u2_n108, u1_u15_u2_n109, u1_u15_u2_n110, u1_u15_u2_n111, u1_u15_u2_n112, u1_u15_u2_n113, u1_u15_u2_n114, u1_u15_u2_n115, u1_u15_u2_n116, 
       u1_u15_u2_n117, u1_u15_u2_n118, u1_u15_u2_n119, u1_u15_u2_n120, u1_u15_u2_n121, u1_u15_u2_n122, u1_u15_u2_n123, u1_u15_u2_n124, u1_u15_u2_n125, 
       u1_u15_u2_n126, u1_u15_u2_n127, u1_u15_u2_n128, u1_u15_u2_n129, u1_u15_u2_n130, u1_u15_u2_n131, u1_u15_u2_n132, u1_u15_u2_n133, u1_u15_u2_n134, 
       u1_u15_u2_n135, u1_u15_u2_n136, u1_u15_u2_n137, u1_u15_u2_n138, u1_u15_u2_n139, u1_u15_u2_n140, u1_u15_u2_n141, u1_u15_u2_n142, u1_u15_u2_n143, 
       u1_u15_u2_n144, u1_u15_u2_n145, u1_u15_u2_n146, u1_u15_u2_n147, u1_u15_u2_n148, u1_u15_u2_n149, u1_u15_u2_n150, u1_u15_u2_n151, u1_u15_u2_n152, 
       u1_u15_u2_n153, u1_u15_u2_n154, u1_u15_u2_n155, u1_u15_u2_n156, u1_u15_u2_n157, u1_u15_u2_n158, u1_u15_u2_n159, u1_u15_u2_n160, u1_u15_u2_n161, 
       u1_u15_u2_n162, u1_u15_u2_n163, u1_u15_u2_n164, u1_u15_u2_n165, u1_u15_u2_n166, u1_u15_u2_n167, u1_u15_u2_n168, u1_u15_u2_n169, u1_u15_u2_n170, 
       u1_u15_u2_n171, u1_u15_u2_n172, u1_u15_u2_n173, u1_u15_u2_n174, u1_u15_u2_n175, u1_u15_u2_n176, u1_u15_u2_n177, u1_u15_u2_n178, u1_u15_u2_n179, 
       u1_u15_u2_n180, u1_u15_u2_n181, u1_u15_u2_n182, u1_u15_u2_n183, u1_u15_u2_n184, u1_u15_u2_n185, u1_u15_u2_n186, u1_u15_u2_n187, u1_u15_u2_n188, 
       u1_u15_u2_n95, u1_u15_u2_n96, u1_u15_u2_n97, u1_u15_u2_n98, u1_u15_u2_n99, u1_u1_X_10, u1_u1_X_11, u1_u1_X_12, u1_u1_X_13, 
       u1_u1_X_14, u1_u1_X_15, u1_u1_X_16, u1_u1_X_17, u1_u1_X_18, u1_u1_X_7, u1_u1_X_8, u1_u1_X_9, u1_u1_u1_n100, 
       u1_u1_u1_n101, u1_u1_u1_n102, u1_u1_u1_n103, u1_u1_u1_n104, u1_u1_u1_n105, u1_u1_u1_n106, u1_u1_u1_n107, u1_u1_u1_n108, u1_u1_u1_n109, 
       u1_u1_u1_n110, u1_u1_u1_n111, u1_u1_u1_n112, u1_u1_u1_n113, u1_u1_u1_n114, u1_u1_u1_n115, u1_u1_u1_n116, u1_u1_u1_n117, u1_u1_u1_n118, 
       u1_u1_u1_n119, u1_u1_u1_n120, u1_u1_u1_n121, u1_u1_u1_n122, u1_u1_u1_n123, u1_u1_u1_n124, u1_u1_u1_n125, u1_u1_u1_n126, u1_u1_u1_n127, 
       u1_u1_u1_n128, u1_u1_u1_n129, u1_u1_u1_n130, u1_u1_u1_n131, u1_u1_u1_n132, u1_u1_u1_n133, u1_u1_u1_n134, u1_u1_u1_n135, u1_u1_u1_n136, 
       u1_u1_u1_n137, u1_u1_u1_n138, u1_u1_u1_n139, u1_u1_u1_n140, u1_u1_u1_n141, u1_u1_u1_n142, u1_u1_u1_n143, u1_u1_u1_n144, u1_u1_u1_n145, 
       u1_u1_u1_n146, u1_u1_u1_n147, u1_u1_u1_n148, u1_u1_u1_n149, u1_u1_u1_n150, u1_u1_u1_n151, u1_u1_u1_n152, u1_u1_u1_n153, u1_u1_u1_n154, 
       u1_u1_u1_n155, u1_u1_u1_n156, u1_u1_u1_n157, u1_u1_u1_n158, u1_u1_u1_n159, u1_u1_u1_n160, u1_u1_u1_n161, u1_u1_u1_n162, u1_u1_u1_n163, 
       u1_u1_u1_n164, u1_u1_u1_n165, u1_u1_u1_n166, u1_u1_u1_n167, u1_u1_u1_n168, u1_u1_u1_n169, u1_u1_u1_n170, u1_u1_u1_n171, u1_u1_u1_n172, 
       u1_u1_u1_n173, u1_u1_u1_n174, u1_u1_u1_n175, u1_u1_u1_n176, u1_u1_u1_n177, u1_u1_u1_n178, u1_u1_u1_n179, u1_u1_u1_n180, u1_u1_u1_n181, 
       u1_u1_u1_n182, u1_u1_u1_n183, u1_u1_u1_n184, u1_u1_u1_n185, u1_u1_u1_n186, u1_u1_u1_n187, u1_u1_u1_n188, u1_u1_u1_n95, u1_u1_u1_n96, 
       u1_u1_u1_n97, u1_u1_u1_n98, u1_u1_u1_n99, u1_u1_u2_n100, u1_u1_u2_n101, u1_u1_u2_n102, u1_u1_u2_n103, u1_u1_u2_n104, u1_u1_u2_n105, 
       u1_u1_u2_n106, u1_u1_u2_n107, u1_u1_u2_n108, u1_u1_u2_n109, u1_u1_u2_n110, u1_u1_u2_n111, u1_u1_u2_n112, u1_u1_u2_n113, u1_u1_u2_n114, 
       u1_u1_u2_n115, u1_u1_u2_n116, u1_u1_u2_n117, u1_u1_u2_n118, u1_u1_u2_n119, u1_u1_u2_n120, u1_u1_u2_n121, u1_u1_u2_n122, u1_u1_u2_n123, 
       u1_u1_u2_n124, u1_u1_u2_n125, u1_u1_u2_n126, u1_u1_u2_n127, u1_u1_u2_n128, u1_u1_u2_n129, u1_u1_u2_n130, u1_u1_u2_n131, u1_u1_u2_n132, 
       u1_u1_u2_n133, u1_u1_u2_n134, u1_u1_u2_n135, u1_u1_u2_n136, u1_u1_u2_n137, u1_u1_u2_n138, u1_u1_u2_n139, u1_u1_u2_n140, u1_u1_u2_n141, 
       u1_u1_u2_n142, u1_u1_u2_n143, u1_u1_u2_n144, u1_u1_u2_n145, u1_u1_u2_n146, u1_u1_u2_n147, u1_u1_u2_n148, u1_u1_u2_n149, u1_u1_u2_n150, 
       u1_u1_u2_n151, u1_u1_u2_n152, u1_u1_u2_n153, u1_u1_u2_n154, u1_u1_u2_n155, u1_u1_u2_n156, u1_u1_u2_n157, u1_u1_u2_n158, u1_u1_u2_n159, 
       u1_u1_u2_n160, u1_u1_u2_n161, u1_u1_u2_n162, u1_u1_u2_n163, u1_u1_u2_n164, u1_u1_u2_n165, u1_u1_u2_n166, u1_u1_u2_n167, u1_u1_u2_n168, 
       u1_u1_u2_n169, u1_u1_u2_n170, u1_u1_u2_n171, u1_u1_u2_n172, u1_u1_u2_n173, u1_u1_u2_n174, u1_u1_u2_n175, u1_u1_u2_n176, u1_u1_u2_n177, 
       u1_u1_u2_n178, u1_u1_u2_n179, u1_u1_u2_n180, u1_u1_u2_n181, u1_u1_u2_n182, u1_u1_u2_n183, u1_u1_u2_n184, u1_u1_u2_n185, u1_u1_u2_n186, 
       u1_u1_u2_n187, u1_u1_u2_n188, u1_u1_u2_n95, u1_u1_u2_n96, u1_u1_u2_n97, u1_u1_u2_n98, u1_u1_u2_n99, u1_u4_X_10, u1_u4_X_11, 
       u1_u4_X_12, u1_u4_X_7, u1_u4_X_8, u1_u4_X_9, u1_u4_u1_n100, u1_u4_u1_n101, u1_u4_u1_n102, u1_u4_u1_n103, u1_u4_u1_n104, 
       u1_u4_u1_n105, u1_u4_u1_n106, u1_u4_u1_n107, u1_u4_u1_n108, u1_u4_u1_n109, u1_u4_u1_n110, u1_u4_u1_n111, u1_u4_u1_n112, u1_u4_u1_n113, 
       u1_u4_u1_n114, u1_u4_u1_n115, u1_u4_u1_n116, u1_u4_u1_n117, u1_u4_u1_n118, u1_u4_u1_n119, u1_u4_u1_n120, u1_u4_u1_n121, u1_u4_u1_n122, 
       u1_u4_u1_n123, u1_u4_u1_n124, u1_u4_u1_n125, u1_u4_u1_n126, u1_u4_u1_n127, u1_u4_u1_n128, u1_u4_u1_n129, u1_u4_u1_n130, u1_u4_u1_n131, 
       u1_u4_u1_n132, u1_u4_u1_n133, u1_u4_u1_n134, u1_u4_u1_n135, u1_u4_u1_n136, u1_u4_u1_n137, u1_u4_u1_n138, u1_u4_u1_n139, u1_u4_u1_n140, 
       u1_u4_u1_n141, u1_u4_u1_n142, u1_u4_u1_n143, u1_u4_u1_n144, u1_u4_u1_n145, u1_u4_u1_n146, u1_u4_u1_n147, u1_u4_u1_n148, u1_u4_u1_n149, 
       u1_u4_u1_n150, u1_u4_u1_n151, u1_u4_u1_n152, u1_u4_u1_n153, u1_u4_u1_n154, u1_u4_u1_n155, u1_u4_u1_n156, u1_u4_u1_n157, u1_u4_u1_n158, 
       u1_u4_u1_n159, u1_u4_u1_n160, u1_u4_u1_n161, u1_u4_u1_n162, u1_u4_u1_n163, u1_u4_u1_n164, u1_u4_u1_n165, u1_u4_u1_n166, u1_u4_u1_n167, 
       u1_u4_u1_n168, u1_u4_u1_n169, u1_u4_u1_n170, u1_u4_u1_n171, u1_u4_u1_n172, u1_u4_u1_n173, u1_u4_u1_n174, u1_u4_u1_n175, u1_u4_u1_n176, 
       u1_u4_u1_n177, u1_u4_u1_n178, u1_u4_u1_n179, u1_u4_u1_n180, u1_u4_u1_n181, u1_u4_u1_n182, u1_u4_u1_n183, u1_u4_u1_n184, u1_u4_u1_n185, 
       u1_u4_u1_n186, u1_u4_u1_n187, u1_u4_u1_n188, u1_u4_u1_n95, u1_u4_u1_n96, u1_u4_u1_n97, u1_u4_u1_n98, u1_u4_u1_n99, u1_u9_X_1, 
       u1_u9_X_10, u1_u9_X_11, u1_u9_X_12, u1_u9_X_13, u1_u9_X_14, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_18, 
       u1_u9_X_2, u1_u9_X_3, u1_u9_X_4, u1_u9_X_5, u1_u9_X_6, u1_u9_X_7, u1_u9_X_8, u1_u9_X_9, u1_u9_u0_n100, 
       u1_u9_u0_n101, u1_u9_u0_n102, u1_u9_u0_n103, u1_u9_u0_n104, u1_u9_u0_n105, u1_u9_u0_n106, u1_u9_u0_n107, u1_u9_u0_n108, u1_u9_u0_n109, 
       u1_u9_u0_n110, u1_u9_u0_n111, u1_u9_u0_n112, u1_u9_u0_n113, u1_u9_u0_n114, u1_u9_u0_n115, u1_u9_u0_n116, u1_u9_u0_n117, u1_u9_u0_n118, 
       u1_u9_u0_n119, u1_u9_u0_n120, u1_u9_u0_n121, u1_u9_u0_n122, u1_u9_u0_n123, u1_u9_u0_n124, u1_u9_u0_n125, u1_u9_u0_n126, u1_u9_u0_n127, 
       u1_u9_u0_n128, u1_u9_u0_n129, u1_u9_u0_n130, u1_u9_u0_n131, u1_u9_u0_n132, u1_u9_u0_n133, u1_u9_u0_n134, u1_u9_u0_n135, u1_u9_u0_n136, 
       u1_u9_u0_n137, u1_u9_u0_n138, u1_u9_u0_n139, u1_u9_u0_n140, u1_u9_u0_n141, u1_u9_u0_n142, u1_u9_u0_n143, u1_u9_u0_n144, u1_u9_u0_n145, 
       u1_u9_u0_n146, u1_u9_u0_n147, u1_u9_u0_n148, u1_u9_u0_n149, u1_u9_u0_n150, u1_u9_u0_n151, u1_u9_u0_n152, u1_u9_u0_n153, u1_u9_u0_n154, 
       u1_u9_u0_n155, u1_u9_u0_n156, u1_u9_u0_n157, u1_u9_u0_n158, u1_u9_u0_n159, u1_u9_u0_n160, u1_u9_u0_n161, u1_u9_u0_n162, u1_u9_u0_n163, 
       u1_u9_u0_n164, u1_u9_u0_n165, u1_u9_u0_n166, u1_u9_u0_n167, u1_u9_u0_n168, u1_u9_u0_n169, u1_u9_u0_n170, u1_u9_u0_n171, u1_u9_u0_n172, 
       u1_u9_u0_n173, u1_u9_u0_n174, u1_u9_u0_n88, u1_u9_u0_n89, u1_u9_u0_n90, u1_u9_u0_n91, u1_u9_u0_n92, u1_u9_u0_n93, u1_u9_u0_n94, 
       u1_u9_u0_n95, u1_u9_u0_n96, u1_u9_u0_n97, u1_u9_u0_n98, u1_u9_u0_n99, u1_u9_u1_n100, u1_u9_u1_n101, u1_u9_u1_n102, u1_u9_u1_n103, 
       u1_u9_u1_n104, u1_u9_u1_n105, u1_u9_u1_n106, u1_u9_u1_n107, u1_u9_u1_n108, u1_u9_u1_n109, u1_u9_u1_n110, u1_u9_u1_n111, u1_u9_u1_n112, 
       u1_u9_u1_n113, u1_u9_u1_n114, u1_u9_u1_n115, u1_u9_u1_n116, u1_u9_u1_n117, u1_u9_u1_n118, u1_u9_u1_n119, u1_u9_u1_n120, u1_u9_u1_n121, 
       u1_u9_u1_n122, u1_u9_u1_n123, u1_u9_u1_n124, u1_u9_u1_n125, u1_u9_u1_n126, u1_u9_u1_n127, u1_u9_u1_n128, u1_u9_u1_n129, u1_u9_u1_n130, 
       u1_u9_u1_n131, u1_u9_u1_n132, u1_u9_u1_n133, u1_u9_u1_n134, u1_u9_u1_n135, u1_u9_u1_n136, u1_u9_u1_n137, u1_u9_u1_n138, u1_u9_u1_n139, 
       u1_u9_u1_n140, u1_u9_u1_n141, u1_u9_u1_n142, u1_u9_u1_n143, u1_u9_u1_n144, u1_u9_u1_n145, u1_u9_u1_n146, u1_u9_u1_n147, u1_u9_u1_n148, 
       u1_u9_u1_n149, u1_u9_u1_n150, u1_u9_u1_n151, u1_u9_u1_n152, u1_u9_u1_n153, u1_u9_u1_n154, u1_u9_u1_n155, u1_u9_u1_n156, u1_u9_u1_n157, 
       u1_u9_u1_n158, u1_u9_u1_n159, u1_u9_u1_n160, u1_u9_u1_n161, u1_u9_u1_n162, u1_u9_u1_n163, u1_u9_u1_n164, u1_u9_u1_n165, u1_u9_u1_n166, 
       u1_u9_u1_n167, u1_u9_u1_n168, u1_u9_u1_n169, u1_u9_u1_n170, u1_u9_u1_n171, u1_u9_u1_n172, u1_u9_u1_n173, u1_u9_u1_n174, u1_u9_u1_n175, 
       u1_u9_u1_n176, u1_u9_u1_n177, u1_u9_u1_n178, u1_u9_u1_n179, u1_u9_u1_n180, u1_u9_u1_n181, u1_u9_u1_n182, u1_u9_u1_n183, u1_u9_u1_n184, 
       u1_u9_u1_n185, u1_u9_u1_n186, u1_u9_u1_n187, u1_u9_u1_n188, u1_u9_u1_n95, u1_u9_u1_n96, u1_u9_u1_n97, u1_u9_u1_n98, u1_u9_u1_n99, 
       u1_u9_u2_n100, u1_u9_u2_n101, u1_u9_u2_n102, u1_u9_u2_n103, u1_u9_u2_n104, u1_u9_u2_n105, u1_u9_u2_n106, u1_u9_u2_n107, u1_u9_u2_n108, 
       u1_u9_u2_n109, u1_u9_u2_n110, u1_u9_u2_n111, u1_u9_u2_n112, u1_u9_u2_n113, u1_u9_u2_n114, u1_u9_u2_n115, u1_u9_u2_n116, u1_u9_u2_n117, 
       u1_u9_u2_n118, u1_u9_u2_n119, u1_u9_u2_n120, u1_u9_u2_n121, u1_u9_u2_n122, u1_u9_u2_n123, u1_u9_u2_n124, u1_u9_u2_n125, u1_u9_u2_n126, 
       u1_u9_u2_n127, u1_u9_u2_n128, u1_u9_u2_n129, u1_u9_u2_n130, u1_u9_u2_n131, u1_u9_u2_n132, u1_u9_u2_n133, u1_u9_u2_n134, u1_u9_u2_n135, 
       u1_u9_u2_n136, u1_u9_u2_n137, u1_u9_u2_n138, u1_u9_u2_n139, u1_u9_u2_n140, u1_u9_u2_n141, u1_u9_u2_n142, u1_u9_u2_n143, u1_u9_u2_n144, 
       u1_u9_u2_n145, u1_u9_u2_n146, u1_u9_u2_n147, u1_u9_u2_n148, u1_u9_u2_n149, u1_u9_u2_n150, u1_u9_u2_n151, u1_u9_u2_n152, u1_u9_u2_n153, 
       u1_u9_u2_n154, u1_u9_u2_n155, u1_u9_u2_n156, u1_u9_u2_n157, u1_u9_u2_n158, u1_u9_u2_n159, u1_u9_u2_n160, u1_u9_u2_n161, u1_u9_u2_n162, 
       u1_u9_u2_n163, u1_u9_u2_n164, u1_u9_u2_n165, u1_u9_u2_n166, u1_u9_u2_n167, u1_u9_u2_n168, u1_u9_u2_n169, u1_u9_u2_n170, u1_u9_u2_n171, 
       u1_u9_u2_n172, u1_u9_u2_n173, u1_u9_u2_n174, u1_u9_u2_n175, u1_u9_u2_n176, u1_u9_u2_n177, u1_u9_u2_n178, u1_u9_u2_n179, u1_u9_u2_n180, 
       u1_u9_u2_n181, u1_u9_u2_n182, u1_u9_u2_n183, u1_u9_u2_n184, u1_u9_u2_n185, u1_u9_u2_n186, u1_u9_u2_n187, u1_u9_u2_n188, u1_u9_u2_n95, 
       u1_u9_u2_n96, u1_u9_u2_n97, u1_u9_u2_n98, u1_u9_u2_n99, u1_uk_n1000, u1_uk_n1001, u1_uk_n1002, u1_uk_n1003, u1_uk_n1004, 
       u1_uk_n1008, u1_uk_n1020, u1_uk_n1021, u1_uk_n1022, u1_uk_n1023, u1_uk_n1024, u1_uk_n1034, u1_uk_n1035, u1_uk_n1071, 
       u1_uk_n1087, u1_uk_n1175, u1_uk_n1176, u1_uk_n1180, u1_uk_n1183, u1_uk_n1184, u1_uk_n1185, u1_uk_n1189, u1_uk_n1190, 
       u1_uk_n1191, u1_uk_n1192, u1_uk_n1197, u1_uk_n1198, u1_uk_n1204, u1_uk_n1205, u1_uk_n1209, u1_uk_n1214, u1_uk_n1215, 
       u1_uk_n299, u1_uk_n301, u1_uk_n305, u1_uk_n306, u1_uk_n338, u1_uk_n376, u1_uk_n377, u1_uk_n379, u1_uk_n382, 
       u1_uk_n385, u1_uk_n437, u1_uk_n443, u1_uk_n454, u1_uk_n496, u1_uk_n500, u1_uk_n501, u1_uk_n671, u1_uk_n672, 
       u1_uk_n676, u1_uk_n685, u1_uk_n686, u1_uk_n688, u1_uk_n689, u1_uk_n692, u1_uk_n702, u1_uk_n945, u1_uk_n948, 
       u1_uk_n949, u1_uk_n950, u1_uk_n980, u1_uk_n981, u1_uk_n982, u1_uk_n983, u1_uk_n996, u1_uk_n997, u1_uk_n998, 
       u1_uk_n999, u2_K16_25, u2_K16_27, u2_K16_28, u2_K16_29, u2_K16_30, u2_K3_1, u2_K3_14, u2_K3_17, 
       u2_K3_18, u2_K3_2, u2_K3_3, u2_K3_4, u2_K3_5, u2_K3_6, u2_out15_14, u2_out15_25, u2_out15_3, 
       u2_out15_8, u2_out2_16, u2_out2_17, u2_out2_23, u2_out2_24, u2_out2_30, u2_out2_31, u2_out2_6, u2_out2_9, 
       u2_u15_X_25, u2_u15_X_26, u2_u15_X_27, u2_u15_X_28, u2_u15_X_29, u2_u15_X_30, u2_u15_u4_n100, u2_u15_u4_n101, u2_u15_u4_n102, 
       u2_u15_u4_n103, u2_u15_u4_n104, u2_u15_u4_n105, u2_u15_u4_n106, u2_u15_u4_n107, u2_u15_u4_n108, u2_u15_u4_n109, u2_u15_u4_n110, u2_u15_u4_n111, 
       u2_u15_u4_n112, u2_u15_u4_n113, u2_u15_u4_n114, u2_u15_u4_n115, u2_u15_u4_n116, u2_u15_u4_n117, u2_u15_u4_n118, u2_u15_u4_n119, u2_u15_u4_n120, 
       u2_u15_u4_n121, u2_u15_u4_n122, u2_u15_u4_n123, u2_u15_u4_n124, u2_u15_u4_n125, u2_u15_u4_n126, u2_u15_u4_n127, u2_u15_u4_n128, u2_u15_u4_n129, 
       u2_u15_u4_n130, u2_u15_u4_n131, u2_u15_u4_n132, u2_u15_u4_n133, u2_u15_u4_n134, u2_u15_u4_n135, u2_u15_u4_n136, u2_u15_u4_n137, u2_u15_u4_n138, 
       u2_u15_u4_n139, u2_u15_u4_n140, u2_u15_u4_n141, u2_u15_u4_n142, u2_u15_u4_n143, u2_u15_u4_n144, u2_u15_u4_n145, u2_u15_u4_n146, u2_u15_u4_n147, 
       u2_u15_u4_n148, u2_u15_u4_n149, u2_u15_u4_n150, u2_u15_u4_n151, u2_u15_u4_n152, u2_u15_u4_n153, u2_u15_u4_n154, u2_u15_u4_n155, u2_u15_u4_n156, 
       u2_u15_u4_n157, u2_u15_u4_n158, u2_u15_u4_n159, u2_u15_u4_n160, u2_u15_u4_n161, u2_u15_u4_n162, u2_u15_u4_n163, u2_u15_u4_n164, u2_u15_u4_n165, 
       u2_u15_u4_n166, u2_u15_u4_n167, u2_u15_u4_n168, u2_u15_u4_n169, u2_u15_u4_n170, u2_u15_u4_n171, u2_u15_u4_n172, u2_u15_u4_n173, u2_u15_u4_n174, 
       u2_u15_u4_n175, u2_u15_u4_n176, u2_u15_u4_n177, u2_u15_u4_n178, u2_u15_u4_n179, u2_u15_u4_n180, u2_u15_u4_n181, u2_u15_u4_n182, u2_u15_u4_n183, 
       u2_u15_u4_n184, u2_u15_u4_n185, u2_u15_u4_n186, u2_u15_u4_n94, u2_u15_u4_n95, u2_u15_u4_n96, u2_u15_u4_n97, u2_u15_u4_n98, u2_u15_u4_n99, 
       u2_u2_X_1, u2_u2_X_13, u2_u2_X_14, u2_u2_X_15, u2_u2_X_16, u2_u2_X_17, u2_u2_X_18, u2_u2_X_2, u2_u2_X_3, 
       u2_u2_X_4, u2_u2_X_5, u2_u2_X_6, u2_u2_u0_n100, u2_u2_u0_n101, u2_u2_u0_n102, u2_u2_u0_n103, u2_u2_u0_n104, u2_u2_u0_n105, 
       u2_u2_u0_n106, u2_u2_u0_n107, u2_u2_u0_n108, u2_u2_u0_n109, u2_u2_u0_n110, u2_u2_u0_n111, u2_u2_u0_n112, u2_u2_u0_n113, u2_u2_u0_n114, 
       u2_u2_u0_n115, u2_u2_u0_n116, u2_u2_u0_n117, u2_u2_u0_n118, u2_u2_u0_n119, u2_u2_u0_n120, u2_u2_u0_n121, u2_u2_u0_n122, u2_u2_u0_n123, 
       u2_u2_u0_n124, u2_u2_u0_n125, u2_u2_u0_n126, u2_u2_u0_n127, u2_u2_u0_n128, u2_u2_u0_n129, u2_u2_u0_n130, u2_u2_u0_n131, u2_u2_u0_n132, 
       u2_u2_u0_n133, u2_u2_u0_n134, u2_u2_u0_n135, u2_u2_u0_n136, u2_u2_u0_n137, u2_u2_u0_n138, u2_u2_u0_n139, u2_u2_u0_n140, u2_u2_u0_n141, 
       u2_u2_u0_n142, u2_u2_u0_n143, u2_u2_u0_n144, u2_u2_u0_n145, u2_u2_u0_n146, u2_u2_u0_n147, u2_u2_u0_n148, u2_u2_u0_n149, u2_u2_u0_n150, 
       u2_u2_u0_n151, u2_u2_u0_n152, u2_u2_u0_n153, u2_u2_u0_n154, u2_u2_u0_n155, u2_u2_u0_n156, u2_u2_u0_n157, u2_u2_u0_n158, u2_u2_u0_n159, 
       u2_u2_u0_n160, u2_u2_u0_n161, u2_u2_u0_n162, u2_u2_u0_n163, u2_u2_u0_n164, u2_u2_u0_n165, u2_u2_u0_n166, u2_u2_u0_n167, u2_u2_u0_n168, 
       u2_u2_u0_n169, u2_u2_u0_n170, u2_u2_u0_n171, u2_u2_u0_n172, u2_u2_u0_n173, u2_u2_u0_n174, u2_u2_u0_n88, u2_u2_u0_n89, u2_u2_u0_n90, 
       u2_u2_u0_n91, u2_u2_u0_n92, u2_u2_u0_n93, u2_u2_u0_n94, u2_u2_u0_n95, u2_u2_u0_n96, u2_u2_u0_n97, u2_u2_u0_n98, u2_u2_u0_n99, 
       u2_u2_u2_n100, u2_u2_u2_n101, u2_u2_u2_n102, u2_u2_u2_n103, u2_u2_u2_n104, u2_u2_u2_n105, u2_u2_u2_n106, u2_u2_u2_n107, u2_u2_u2_n108, 
       u2_u2_u2_n109, u2_u2_u2_n110, u2_u2_u2_n111, u2_u2_u2_n112, u2_u2_u2_n113, u2_u2_u2_n114, u2_u2_u2_n115, u2_u2_u2_n116, u2_u2_u2_n117, 
       u2_u2_u2_n118, u2_u2_u2_n119, u2_u2_u2_n120, u2_u2_u2_n121, u2_u2_u2_n122, u2_u2_u2_n123, u2_u2_u2_n124, u2_u2_u2_n125, u2_u2_u2_n126, 
       u2_u2_u2_n127, u2_u2_u2_n128, u2_u2_u2_n129, u2_u2_u2_n130, u2_u2_u2_n131, u2_u2_u2_n132, u2_u2_u2_n133, u2_u2_u2_n134, u2_u2_u2_n135, 
       u2_u2_u2_n136, u2_u2_u2_n137, u2_u2_u2_n138, u2_u2_u2_n139, u2_u2_u2_n140, u2_u2_u2_n141, u2_u2_u2_n142, u2_u2_u2_n143, u2_u2_u2_n144, 
       u2_u2_u2_n145, u2_u2_u2_n146, u2_u2_u2_n147, u2_u2_u2_n148, u2_u2_u2_n149, u2_u2_u2_n150, u2_u2_u2_n151, u2_u2_u2_n152, u2_u2_u2_n153, 
       u2_u2_u2_n154, u2_u2_u2_n155, u2_u2_u2_n156, u2_u2_u2_n157, u2_u2_u2_n158, u2_u2_u2_n159, u2_u2_u2_n160, u2_u2_u2_n161, u2_u2_u2_n162, 
       u2_u2_u2_n163, u2_u2_u2_n164, u2_u2_u2_n165, u2_u2_u2_n166, u2_u2_u2_n167, u2_u2_u2_n168, u2_u2_u2_n169, u2_u2_u2_n170, u2_u2_u2_n171, 
       u2_u2_u2_n172, u2_u2_u2_n173, u2_u2_u2_n174, u2_u2_u2_n175, u2_u2_u2_n176, u2_u2_u2_n177, u2_u2_u2_n178, u2_u2_u2_n179, u2_u2_u2_n180, 
       u2_u2_u2_n181, u2_u2_u2_n182, u2_u2_u2_n183, u2_u2_u2_n184, u2_u2_u2_n185, u2_u2_u2_n186, u2_u2_u2_n187, u2_u2_u2_n188, u2_u2_u2_n95, 
       u2_u2_u2_n96, u2_u2_u2_n97, u2_u2_u2_n98, u2_u2_u2_n99, u2_uk_n1013,  u2_uk_n957;
  XOR2_X1 u0_U60 (.B( u0_L13_32 ) , .Z( u0_N479 ) , .A( u0_out14_32 ) );
  XOR2_X1 u0_U65 (.B( u0_L13_27 ) , .Z( u0_N474 ) , .A( u0_out14_27 ) );
  XOR2_X1 u0_U71 (.B( u0_L13_22 ) , .Z( u0_N469 ) , .A( u0_out14_22 ) );
  XOR2_X1 u0_U72 (.B( u0_L13_21 ) , .Z( u0_N468 ) , .A( u0_out14_21 ) );
  XOR2_X1 u0_U78 (.B( u0_L13_15 ) , .Z( u0_N462 ) , .A( u0_out14_15 ) );
  XOR2_X1 u0_U82 (.B( u0_L13_12 ) , .Z( u0_N459 ) , .A( u0_out14_12 ) );
  XOR2_X1 u0_U87 (.B( u0_L13_7 ) , .Z( u0_N454 ) , .A( u0_out14_7 ) );
  XOR2_X1 u0_U89 (.B( u0_L13_5 ) , .Z( u0_N452 ) , .A( u0_out14_5 ) );
  XOR2_X1 u0_u14_U10 (.B( u0_K15_45 ) , .A( u0_R13_30 ) , .Z( u0_u14_X_45 ) );
  XOR2_X1 u0_u14_U11 (.B( u0_K15_44 ) , .A( u0_R13_29 ) , .Z( u0_u14_X_44 ) );
  XOR2_X1 u0_u14_U12 (.B( u0_K15_43 ) , .A( u0_R13_28 ) , .Z( u0_u14_X_43 ) );
  XOR2_X1 u0_u14_U13 (.B( u0_K15_42 ) , .A( u0_R13_29 ) , .Z( u0_u14_X_42 ) );
  XOR2_X1 u0_u14_U14 (.B( u0_K15_41 ) , .A( u0_R13_28 ) , .Z( u0_u14_X_41 ) );
  XOR2_X1 u0_u14_U15 (.B( u0_K15_40 ) , .A( u0_R13_27 ) , .Z( u0_u14_X_40 ) );
  XOR2_X1 u0_u14_U17 (.B( u0_K15_39 ) , .A( u0_R13_26 ) , .Z( u0_u14_X_39 ) );
  XOR2_X1 u0_u14_U18 (.B( u0_K15_38 ) , .A( u0_R13_25 ) , .Z( u0_u14_X_38 ) );
  XOR2_X1 u0_u14_U19 (.B( u0_K15_37 ) , .A( u0_R13_24 ) , .Z( u0_u14_X_37 ) );
  XOR2_X1 u0_u14_U7 (.B( u0_K15_48 ) , .A( u0_R13_1 ) , .Z( u0_u14_X_48 ) );
  XOR2_X1 u0_u14_U8 (.B( u0_K15_47 ) , .A( u0_R13_32 ) , .Z( u0_u14_X_47 ) );
  XOR2_X1 u0_u14_U9 (.B( u0_K15_46 ) , .A( u0_R13_31 ) , .Z( u0_u14_X_46 ) );
  AOI21_X1 u0_u14_u6_U10 (.ZN( u0_u14_u6_n106 ) , .A( u0_u14_u6_n142 ) , .B2( u0_u14_u6_n159 ) , .B1( u0_u14_u6_n164 ) );
  INV_X1 u0_u14_u6_U11 (.A( u0_u14_u6_n155 ) , .ZN( u0_u14_u6_n161 ) );
  INV_X1 u0_u14_u6_U12 (.A( u0_u14_u6_n128 ) , .ZN( u0_u14_u6_n164 ) );
  NAND2_X1 u0_u14_u6_U13 (.ZN( u0_u14_u6_n110 ) , .A1( u0_u14_u6_n122 ) , .A2( u0_u14_u6_n129 ) );
  NAND2_X1 u0_u14_u6_U14 (.ZN( u0_u14_u6_n124 ) , .A2( u0_u14_u6_n146 ) , .A1( u0_u14_u6_n148 ) );
  INV_X1 u0_u14_u6_U15 (.A( u0_u14_u6_n132 ) , .ZN( u0_u14_u6_n171 ) );
  AND2_X1 u0_u14_u6_U16 (.A1( u0_u14_u6_n100 ) , .ZN( u0_u14_u6_n130 ) , .A2( u0_u14_u6_n147 ) );
  INV_X1 u0_u14_u6_U17 (.A( u0_u14_u6_n127 ) , .ZN( u0_u14_u6_n173 ) );
  INV_X1 u0_u14_u6_U18 (.A( u0_u14_u6_n121 ) , .ZN( u0_u14_u6_n167 ) );
  INV_X1 u0_u14_u6_U19 (.A( u0_u14_u6_n100 ) , .ZN( u0_u14_u6_n169 ) );
  INV_X1 u0_u14_u6_U20 (.A( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n170 ) );
  INV_X1 u0_u14_u6_U21 (.A( u0_u14_u6_n113 ) , .ZN( u0_u14_u6_n168 ) );
  AND2_X1 u0_u14_u6_U22 (.A1( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n119 ) , .ZN( u0_u14_u6_n133 ) );
  AND2_X1 u0_u14_u6_U23 (.A2( u0_u14_u6_n121 ) , .A1( u0_u14_u6_n122 ) , .ZN( u0_u14_u6_n131 ) );
  AND3_X1 u0_u14_u6_U24 (.ZN( u0_u14_u6_n120 ) , .A2( u0_u14_u6_n127 ) , .A1( u0_u14_u6_n132 ) , .A3( u0_u14_u6_n145 ) );
  INV_X1 u0_u14_u6_U25 (.A( u0_u14_u6_n146 ) , .ZN( u0_u14_u6_n163 ) );
  AOI222_X1 u0_u14_u6_U26 (.ZN( u0_u14_u6_n114 ) , .A1( u0_u14_u6_n118 ) , .A2( u0_u14_u6_n126 ) , .B2( u0_u14_u6_n151 ) , .C2( u0_u14_u6_n159 ) , .C1( u0_u14_u6_n168 ) , .B1( u0_u14_u6_n169 ) );
  NOR2_X1 u0_u14_u6_U27 (.A1( u0_u14_u6_n162 ) , .A2( u0_u14_u6_n165 ) , .ZN( u0_u14_u6_n98 ) );
  AOI211_X1 u0_u14_u6_U28 (.B( u0_u14_u6_n149 ) , .A( u0_u14_u6_n150 ) , .C2( u0_u14_u6_n151 ) , .C1( u0_u14_u6_n152 ) , .ZN( u0_u14_u6_n153 ) );
  AOI21_X1 u0_u14_u6_U29 (.B2( u0_u14_u6_n147 ) , .B1( u0_u14_u6_n148 ) , .ZN( u0_u14_u6_n149 ) , .A( u0_u14_u6_n158 ) );
  INV_X1 u0_u14_u6_U3 (.A( u0_u14_u6_n110 ) , .ZN( u0_u14_u6_n166 ) );
  AOI21_X1 u0_u14_u6_U30 (.A( u0_u14_u6_n144 ) , .B2( u0_u14_u6_n145 ) , .B1( u0_u14_u6_n146 ) , .ZN( u0_u14_u6_n150 ) );
  NAND2_X1 u0_u14_u6_U31 (.A2( u0_u14_u6_n143 ) , .ZN( u0_u14_u6_n152 ) , .A1( u0_u14_u6_n166 ) );
  NAND2_X1 u0_u14_u6_U32 (.A1( u0_u14_u6_n144 ) , .ZN( u0_u14_u6_n151 ) , .A2( u0_u14_u6_n158 ) );
  NAND2_X1 u0_u14_u6_U33 (.ZN( u0_u14_u6_n132 ) , .A1( u0_u14_u6_n91 ) , .A2( u0_u14_u6_n97 ) );
  AOI22_X1 u0_u14_u6_U34 (.B2( u0_u14_u6_n110 ) , .B1( u0_u14_u6_n111 ) , .A1( u0_u14_u6_n112 ) , .ZN( u0_u14_u6_n115 ) , .A2( u0_u14_u6_n161 ) );
  NAND4_X1 u0_u14_u6_U35 (.A3( u0_u14_u6_n109 ) , .ZN( u0_u14_u6_n112 ) , .A4( u0_u14_u6_n132 ) , .A2( u0_u14_u6_n147 ) , .A1( u0_u14_u6_n166 ) );
  NOR2_X1 u0_u14_u6_U36 (.ZN( u0_u14_u6_n109 ) , .A1( u0_u14_u6_n170 ) , .A2( u0_u14_u6_n173 ) );
  NOR2_X1 u0_u14_u6_U37 (.A2( u0_u14_u6_n126 ) , .ZN( u0_u14_u6_n155 ) , .A1( u0_u14_u6_n160 ) );
  NAND2_X1 u0_u14_u6_U38 (.ZN( u0_u14_u6_n146 ) , .A2( u0_u14_u6_n94 ) , .A1( u0_u14_u6_n99 ) );
  AOI211_X1 u0_u14_u6_U39 (.B( u0_u14_u6_n134 ) , .A( u0_u14_u6_n135 ) , .C1( u0_u14_u6_n136 ) , .ZN( u0_u14_u6_n137 ) , .C2( u0_u14_u6_n151 ) );
  AOI22_X1 u0_u14_u6_U4 (.B2( u0_u14_u6_n101 ) , .A1( u0_u14_u6_n102 ) , .ZN( u0_u14_u6_n103 ) , .B1( u0_u14_u6_n160 ) , .A2( u0_u14_u6_n161 ) );
  AOI21_X1 u0_u14_u6_U40 (.B2( u0_u14_u6_n132 ) , .B1( u0_u14_u6_n133 ) , .ZN( u0_u14_u6_n134 ) , .A( u0_u14_u6_n158 ) );
  NAND4_X1 u0_u14_u6_U41 (.A4( u0_u14_u6_n127 ) , .A3( u0_u14_u6_n128 ) , .A2( u0_u14_u6_n129 ) , .A1( u0_u14_u6_n130 ) , .ZN( u0_u14_u6_n136 ) );
  AOI21_X1 u0_u14_u6_U42 (.B1( u0_u14_u6_n131 ) , .ZN( u0_u14_u6_n135 ) , .A( u0_u14_u6_n144 ) , .B2( u0_u14_u6_n146 ) );
  INV_X1 u0_u14_u6_U43 (.A( u0_u14_u6_n111 ) , .ZN( u0_u14_u6_n158 ) );
  NAND2_X1 u0_u14_u6_U44 (.ZN( u0_u14_u6_n127 ) , .A1( u0_u14_u6_n91 ) , .A2( u0_u14_u6_n92 ) );
  NAND2_X1 u0_u14_u6_U45 (.ZN( u0_u14_u6_n129 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n96 ) );
  INV_X1 u0_u14_u6_U46 (.A( u0_u14_u6_n144 ) , .ZN( u0_u14_u6_n159 ) );
  NAND2_X1 u0_u14_u6_U47 (.ZN( u0_u14_u6_n145 ) , .A2( u0_u14_u6_n97 ) , .A1( u0_u14_u6_n98 ) );
  NAND2_X1 u0_u14_u6_U48 (.ZN( u0_u14_u6_n148 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n94 ) );
  NAND2_X1 u0_u14_u6_U49 (.ZN( u0_u14_u6_n108 ) , .A2( u0_u14_u6_n139 ) , .A1( u0_u14_u6_n144 ) );
  NOR2_X1 u0_u14_u6_U5 (.A1( u0_u14_u6_n118 ) , .ZN( u0_u14_u6_n143 ) , .A2( u0_u14_u6_n168 ) );
  NAND2_X1 u0_u14_u6_U50 (.ZN( u0_u14_u6_n121 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n97 ) );
  NAND2_X1 u0_u14_u6_U51 (.ZN( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n95 ) );
  AND2_X1 u0_u14_u6_U52 (.ZN( u0_u14_u6_n118 ) , .A2( u0_u14_u6_n91 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U53 (.ZN( u0_u14_u6_n147 ) , .A2( u0_u14_u6_n98 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U54 (.ZN( u0_u14_u6_n128 ) , .A1( u0_u14_u6_n94 ) , .A2( u0_u14_u6_n96 ) );
  NAND2_X1 u0_u14_u6_U55 (.ZN( u0_u14_u6_n119 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U56 (.ZN( u0_u14_u6_n123 ) , .A2( u0_u14_u6_n91 ) , .A1( u0_u14_u6_n96 ) );
  NAND2_X1 u0_u14_u6_U57 (.ZN( u0_u14_u6_n100 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n98 ) );
  NAND2_X1 u0_u14_u6_U58 (.ZN( u0_u14_u6_n122 ) , .A1( u0_u14_u6_n94 ) , .A2( u0_u14_u6_n97 ) );
  INV_X1 u0_u14_u6_U59 (.A( u0_u14_u6_n139 ) , .ZN( u0_u14_u6_n160 ) );
  INV_X1 u0_u14_u6_U6 (.ZN( u0_u14_u6_n172 ) , .A( u0_u14_u6_n88 ) );
  NAND2_X1 u0_u14_u6_U60 (.ZN( u0_u14_u6_n113 ) , .A1( u0_u14_u6_n96 ) , .A2( u0_u14_u6_n98 ) );
  NOR2_X1 u0_u14_u6_U61 (.A2( u0_u14_X_40 ) , .A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n126 ) );
  NOR2_X1 u0_u14_u6_U62 (.A2( u0_u14_X_39 ) , .A1( u0_u14_X_42 ) , .ZN( u0_u14_u6_n92 ) );
  NOR2_X1 u0_u14_u6_U63 (.A2( u0_u14_X_39 ) , .A1( u0_u14_u6_n156 ) , .ZN( u0_u14_u6_n97 ) );
  NOR2_X1 u0_u14_u6_U64 (.A2( u0_u14_X_38 ) , .A1( u0_u14_u6_n165 ) , .ZN( u0_u14_u6_n95 ) );
  NOR2_X1 u0_u14_u6_U65 (.A2( u0_u14_X_41 ) , .ZN( u0_u14_u6_n111 ) , .A1( u0_u14_u6_n157 ) );
  NOR2_X1 u0_u14_u6_U66 (.A2( u0_u14_X_37 ) , .A1( u0_u14_u6_n162 ) , .ZN( u0_u14_u6_n94 ) );
  NOR2_X1 u0_u14_u6_U67 (.A2( u0_u14_X_37 ) , .A1( u0_u14_X_38 ) , .ZN( u0_u14_u6_n91 ) );
  NAND2_X1 u0_u14_u6_U68 (.A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n144 ) , .A2( u0_u14_u6_n157 ) );
  NAND2_X1 u0_u14_u6_U69 (.A2( u0_u14_X_40 ) , .A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n139 ) );
  OAI21_X1 u0_u14_u6_U7 (.A( u0_u14_u6_n159 ) , .B1( u0_u14_u6_n169 ) , .B2( u0_u14_u6_n173 ) , .ZN( u0_u14_u6_n90 ) );
  AND2_X1 u0_u14_u6_U70 (.A1( u0_u14_X_39 ) , .A2( u0_u14_u6_n156 ) , .ZN( u0_u14_u6_n96 ) );
  AND2_X1 u0_u14_u6_U71 (.A1( u0_u14_X_39 ) , .A2( u0_u14_X_42 ) , .ZN( u0_u14_u6_n99 ) );
  INV_X1 u0_u14_u6_U72 (.A( u0_u14_X_40 ) , .ZN( u0_u14_u6_n157 ) );
  INV_X1 u0_u14_u6_U73 (.A( u0_u14_X_37 ) , .ZN( u0_u14_u6_n165 ) );
  INV_X1 u0_u14_u6_U74 (.A( u0_u14_X_38 ) , .ZN( u0_u14_u6_n162 ) );
  INV_X1 u0_u14_u6_U75 (.A( u0_u14_X_42 ) , .ZN( u0_u14_u6_n156 ) );
  NAND4_X1 u0_u14_u6_U76 (.ZN( u0_out14_32 ) , .A4( u0_u14_u6_n103 ) , .A3( u0_u14_u6_n104 ) , .A2( u0_u14_u6_n105 ) , .A1( u0_u14_u6_n106 ) );
  AOI22_X1 u0_u14_u6_U77 (.ZN( u0_u14_u6_n105 ) , .A2( u0_u14_u6_n108 ) , .A1( u0_u14_u6_n118 ) , .B2( u0_u14_u6_n126 ) , .B1( u0_u14_u6_n171 ) );
  AOI22_X1 u0_u14_u6_U78 (.ZN( u0_u14_u6_n104 ) , .A1( u0_u14_u6_n111 ) , .B1( u0_u14_u6_n124 ) , .B2( u0_u14_u6_n151 ) , .A2( u0_u14_u6_n93 ) );
  NAND4_X1 u0_u14_u6_U79 (.ZN( u0_out14_12 ) , .A4( u0_u14_u6_n114 ) , .A3( u0_u14_u6_n115 ) , .A2( u0_u14_u6_n116 ) , .A1( u0_u14_u6_n117 ) );
  AOI22_X1 u0_u14_u6_U8 (.A2( u0_u14_u6_n151 ) , .B2( u0_u14_u6_n161 ) , .A1( u0_u14_u6_n167 ) , .B1( u0_u14_u6_n170 ) , .ZN( u0_u14_u6_n89 ) );
  OAI22_X1 u0_u14_u6_U80 (.B2( u0_u14_u6_n111 ) , .ZN( u0_u14_u6_n116 ) , .B1( u0_u14_u6_n126 ) , .A2( u0_u14_u6_n164 ) , .A1( u0_u14_u6_n167 ) );
  OAI21_X1 u0_u14_u6_U81 (.A( u0_u14_u6_n108 ) , .ZN( u0_u14_u6_n117 ) , .B2( u0_u14_u6_n141 ) , .B1( u0_u14_u6_n163 ) );
  OAI211_X1 u0_u14_u6_U82 (.ZN( u0_out14_22 ) , .B( u0_u14_u6_n137 ) , .A( u0_u14_u6_n138 ) , .C2( u0_u14_u6_n139 ) , .C1( u0_u14_u6_n140 ) );
  AOI22_X1 u0_u14_u6_U83 (.B1( u0_u14_u6_n124 ) , .A2( u0_u14_u6_n125 ) , .A1( u0_u14_u6_n126 ) , .ZN( u0_u14_u6_n138 ) , .B2( u0_u14_u6_n161 ) );
  AND4_X1 u0_u14_u6_U84 (.A3( u0_u14_u6_n119 ) , .A1( u0_u14_u6_n120 ) , .A4( u0_u14_u6_n129 ) , .ZN( u0_u14_u6_n140 ) , .A2( u0_u14_u6_n143 ) );
  OAI211_X1 u0_u14_u6_U85 (.ZN( u0_out14_7 ) , .B( u0_u14_u6_n153 ) , .C2( u0_u14_u6_n154 ) , .C1( u0_u14_u6_n155 ) , .A( u0_u14_u6_n174 ) );
  NOR3_X1 u0_u14_u6_U86 (.A1( u0_u14_u6_n141 ) , .ZN( u0_u14_u6_n154 ) , .A3( u0_u14_u6_n164 ) , .A2( u0_u14_u6_n171 ) );
  INV_X1 u0_u14_u6_U87 (.A( u0_u14_u6_n142 ) , .ZN( u0_u14_u6_n174 ) );
  NAND3_X1 u0_u14_u6_U88 (.A2( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n125 ) , .A1( u0_u14_u6_n130 ) , .A3( u0_u14_u6_n131 ) );
  NAND3_X1 u0_u14_u6_U89 (.A3( u0_u14_u6_n133 ) , .ZN( u0_u14_u6_n141 ) , .A1( u0_u14_u6_n145 ) , .A2( u0_u14_u6_n148 ) );
  AOI21_X1 u0_u14_u6_U9 (.B1( u0_u14_u6_n107 ) , .B2( u0_u14_u6_n132 ) , .A( u0_u14_u6_n158 ) , .ZN( u0_u14_u6_n88 ) );
  NAND3_X1 u0_u14_u6_U90 (.ZN( u0_u14_u6_n101 ) , .A3( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n121 ) , .A1( u0_u14_u6_n127 ) );
  NAND3_X1 u0_u14_u6_U91 (.ZN( u0_u14_u6_n102 ) , .A3( u0_u14_u6_n130 ) , .A2( u0_u14_u6_n145 ) , .A1( u0_u14_u6_n166 ) );
  NAND3_X1 u0_u14_u6_U92 (.A3( u0_u14_u6_n113 ) , .A1( u0_u14_u6_n119 ) , .A2( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n93 ) );
  NAND3_X1 u0_u14_u6_U93 (.ZN( u0_u14_u6_n142 ) , .A2( u0_u14_u6_n172 ) , .A3( u0_u14_u6_n89 ) , .A1( u0_u14_u6_n90 ) );
  AND3_X1 u0_u14_u7_U10 (.A3( u0_u14_u7_n110 ) , .A2( u0_u14_u7_n127 ) , .A1( u0_u14_u7_n132 ) , .ZN( u0_u14_u7_n92 ) );
  OAI21_X1 u0_u14_u7_U11 (.A( u0_u14_u7_n161 ) , .B1( u0_u14_u7_n168 ) , .B2( u0_u14_u7_n173 ) , .ZN( u0_u14_u7_n91 ) );
  AOI211_X1 u0_u14_u7_U12 (.A( u0_u14_u7_n117 ) , .ZN( u0_u14_u7_n118 ) , .C2( u0_u14_u7_n126 ) , .C1( u0_u14_u7_n177 ) , .B( u0_u14_u7_n180 ) );
  OAI22_X1 u0_u14_u7_U13 (.B1( u0_u14_u7_n115 ) , .ZN( u0_u14_u7_n117 ) , .A2( u0_u14_u7_n133 ) , .A1( u0_u14_u7_n137 ) , .B2( u0_u14_u7_n162 ) );
  INV_X1 u0_u14_u7_U14 (.A( u0_u14_u7_n116 ) , .ZN( u0_u14_u7_n180 ) );
  NOR3_X1 u0_u14_u7_U15 (.ZN( u0_u14_u7_n115 ) , .A3( u0_u14_u7_n145 ) , .A2( u0_u14_u7_n168 ) , .A1( u0_u14_u7_n169 ) );
  NOR3_X1 u0_u14_u7_U16 (.A2( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n135 ) , .ZN( u0_u14_u7_n136 ) , .A3( u0_u14_u7_n171 ) );
  NOR2_X1 u0_u14_u7_U17 (.A1( u0_u14_u7_n130 ) , .A2( u0_u14_u7_n134 ) , .ZN( u0_u14_u7_n153 ) );
  NOR2_X1 u0_u14_u7_U18 (.ZN( u0_u14_u7_n111 ) , .A2( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n169 ) );
  AOI21_X1 u0_u14_u7_U19 (.ZN( u0_u14_u7_n104 ) , .B2( u0_u14_u7_n112 ) , .B1( u0_u14_u7_n127 ) , .A( u0_u14_u7_n164 ) );
  AOI21_X1 u0_u14_u7_U20 (.ZN( u0_u14_u7_n106 ) , .B1( u0_u14_u7_n133 ) , .B2( u0_u14_u7_n146 ) , .A( u0_u14_u7_n162 ) );
  AOI21_X1 u0_u14_u7_U21 (.A( u0_u14_u7_n101 ) , .ZN( u0_u14_u7_n107 ) , .B2( u0_u14_u7_n128 ) , .B1( u0_u14_u7_n175 ) );
  INV_X1 u0_u14_u7_U22 (.A( u0_u14_u7_n101 ) , .ZN( u0_u14_u7_n165 ) );
  INV_X1 u0_u14_u7_U23 (.A( u0_u14_u7_n138 ) , .ZN( u0_u14_u7_n171 ) );
  INV_X1 u0_u14_u7_U24 (.A( u0_u14_u7_n131 ) , .ZN( u0_u14_u7_n177 ) );
  INV_X1 u0_u14_u7_U25 (.A( u0_u14_u7_n110 ) , .ZN( u0_u14_u7_n174 ) );
  NAND2_X1 u0_u14_u7_U26 (.A1( u0_u14_u7_n129 ) , .A2( u0_u14_u7_n132 ) , .ZN( u0_u14_u7_n149 ) );
  NAND2_X1 u0_u14_u7_U27 (.A1( u0_u14_u7_n113 ) , .A2( u0_u14_u7_n124 ) , .ZN( u0_u14_u7_n130 ) );
  INV_X1 u0_u14_u7_U28 (.A( u0_u14_u7_n128 ) , .ZN( u0_u14_u7_n168 ) );
  INV_X1 u0_u14_u7_U29 (.A( u0_u14_u7_n148 ) , .ZN( u0_u14_u7_n169 ) );
  INV_X1 u0_u14_u7_U3 (.A( u0_u14_u7_n149 ) , .ZN( u0_u14_u7_n175 ) );
  INV_X1 u0_u14_u7_U30 (.A( u0_u14_u7_n112 ) , .ZN( u0_u14_u7_n173 ) );
  INV_X1 u0_u14_u7_U31 (.A( u0_u14_u7_n127 ) , .ZN( u0_u14_u7_n179 ) );
  NOR2_X1 u0_u14_u7_U32 (.ZN( u0_u14_u7_n101 ) , .A2( u0_u14_u7_n150 ) , .A1( u0_u14_u7_n156 ) );
  AOI211_X1 u0_u14_u7_U33 (.B( u0_u14_u7_n154 ) , .A( u0_u14_u7_n155 ) , .C1( u0_u14_u7_n156 ) , .ZN( u0_u14_u7_n157 ) , .C2( u0_u14_u7_n172 ) );
  INV_X1 u0_u14_u7_U34 (.A( u0_u14_u7_n153 ) , .ZN( u0_u14_u7_n172 ) );
  AOI211_X1 u0_u14_u7_U35 (.B( u0_u14_u7_n139 ) , .A( u0_u14_u7_n140 ) , .C2( u0_u14_u7_n141 ) , .ZN( u0_u14_u7_n142 ) , .C1( u0_u14_u7_n156 ) );
  NAND4_X1 u0_u14_u7_U36 (.A3( u0_u14_u7_n127 ) , .A2( u0_u14_u7_n128 ) , .A1( u0_u14_u7_n129 ) , .ZN( u0_u14_u7_n141 ) , .A4( u0_u14_u7_n147 ) );
  AOI21_X1 u0_u14_u7_U37 (.A( u0_u14_u7_n137 ) , .B1( u0_u14_u7_n138 ) , .ZN( u0_u14_u7_n139 ) , .B2( u0_u14_u7_n146 ) );
  OAI22_X1 u0_u14_u7_U38 (.B1( u0_u14_u7_n136 ) , .ZN( u0_u14_u7_n140 ) , .A1( u0_u14_u7_n153 ) , .B2( u0_u14_u7_n162 ) , .A2( u0_u14_u7_n164 ) );
  INV_X1 u0_u14_u7_U39 (.A( u0_u14_u7_n125 ) , .ZN( u0_u14_u7_n161 ) );
  INV_X1 u0_u14_u7_U4 (.A( u0_u14_u7_n154 ) , .ZN( u0_u14_u7_n178 ) );
  AOI21_X1 u0_u14_u7_U40 (.ZN( u0_u14_u7_n123 ) , .B1( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n177 ) , .A( u0_u14_u7_n97 ) );
  AOI21_X1 u0_u14_u7_U41 (.B2( u0_u14_u7_n113 ) , .B1( u0_u14_u7_n124 ) , .A( u0_u14_u7_n125 ) , .ZN( u0_u14_u7_n97 ) );
  INV_X1 u0_u14_u7_U42 (.A( u0_u14_u7_n152 ) , .ZN( u0_u14_u7_n162 ) );
  AOI22_X1 u0_u14_u7_U43 (.A2( u0_u14_u7_n114 ) , .ZN( u0_u14_u7_n119 ) , .B1( u0_u14_u7_n130 ) , .A1( u0_u14_u7_n156 ) , .B2( u0_u14_u7_n165 ) );
  NAND2_X1 u0_u14_u7_U44 (.A2( u0_u14_u7_n112 ) , .ZN( u0_u14_u7_n114 ) , .A1( u0_u14_u7_n175 ) );
  AOI22_X1 u0_u14_u7_U45 (.B2( u0_u14_u7_n149 ) , .B1( u0_u14_u7_n150 ) , .A2( u0_u14_u7_n151 ) , .A1( u0_u14_u7_n152 ) , .ZN( u0_u14_u7_n158 ) );
  NOR2_X1 u0_u14_u7_U46 (.ZN( u0_u14_u7_n137 ) , .A1( u0_u14_u7_n150 ) , .A2( u0_u14_u7_n161 ) );
  AND2_X1 u0_u14_u7_U47 (.ZN( u0_u14_u7_n145 ) , .A2( u0_u14_u7_n98 ) , .A1( u0_u14_u7_n99 ) );
  AOI21_X1 u0_u14_u7_U48 (.ZN( u0_u14_u7_n105 ) , .B2( u0_u14_u7_n110 ) , .A( u0_u14_u7_n125 ) , .B1( u0_u14_u7_n147 ) );
  NAND2_X1 u0_u14_u7_U49 (.ZN( u0_u14_u7_n146 ) , .A1( u0_u14_u7_n95 ) , .A2( u0_u14_u7_n98 ) );
  INV_X1 u0_u14_u7_U5 (.A( u0_u14_u7_n111 ) , .ZN( u0_u14_u7_n170 ) );
  NAND2_X1 u0_u14_u7_U50 (.A2( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n147 ) , .A1( u0_u14_u7_n93 ) );
  NAND2_X1 u0_u14_u7_U51 (.A1( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n127 ) , .A2( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U52 (.A2( u0_u14_u7_n102 ) , .A1( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n133 ) );
  OR2_X1 u0_u14_u7_U53 (.ZN( u0_u14_u7_n126 ) , .A2( u0_u14_u7_n152 ) , .A1( u0_u14_u7_n156 ) );
  NAND2_X1 u0_u14_u7_U54 (.ZN( u0_u14_u7_n112 ) , .A2( u0_u14_u7_n96 ) , .A1( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U55 (.A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n128 ) , .A1( u0_u14_u7_n98 ) );
  INV_X1 u0_u14_u7_U56 (.A( u0_u14_u7_n150 ) , .ZN( u0_u14_u7_n164 ) );
  AND2_X1 u0_u14_u7_U57 (.ZN( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n93 ) , .A2( u0_u14_u7_n98 ) );
  NAND2_X1 u0_u14_u7_U58 (.ZN( u0_u14_u7_n110 ) , .A1( u0_u14_u7_n95 ) , .A2( u0_u14_u7_n96 ) );
  NAND2_X1 u0_u14_u7_U59 (.A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n124 ) , .A1( u0_u14_u7_n96 ) );
  AOI211_X1 u0_u14_u7_U6 (.ZN( u0_u14_u7_n116 ) , .A( u0_u14_u7_n155 ) , .C1( u0_u14_u7_n161 ) , .C2( u0_u14_u7_n171 ) , .B( u0_u14_u7_n94 ) );
  NAND2_X1 u0_u14_u7_U60 (.ZN( u0_u14_u7_n132 ) , .A1( u0_u14_u7_n93 ) , .A2( u0_u14_u7_n96 ) );
  NAND2_X1 u0_u14_u7_U61 (.A2( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n131 ) , .A1( u0_u14_u7_n95 ) );
  NOR2_X1 u0_u14_u7_U62 (.A2( u0_u14_X_47 ) , .ZN( u0_u14_u7_n150 ) , .A1( u0_u14_u7_n163 ) );
  NOR2_X1 u0_u14_u7_U63 (.A2( u0_u14_X_43 ) , .A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n103 ) );
  NOR2_X1 u0_u14_u7_U64 (.A2( u0_u14_X_48 ) , .A1( u0_u14_u7_n166 ) , .ZN( u0_u14_u7_n95 ) );
  NOR2_X1 u0_u14_u7_U65 (.A2( u0_u14_X_44 ) , .A1( u0_u14_u7_n167 ) , .ZN( u0_u14_u7_n98 ) );
  NOR2_X1 u0_u14_u7_U66 (.A2( u0_u14_X_45 ) , .A1( u0_u14_X_48 ) , .ZN( u0_u14_u7_n99 ) );
  NOR2_X1 u0_u14_u7_U67 (.A2( u0_u14_X_46 ) , .A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n152 ) );
  AND2_X1 u0_u14_u7_U68 (.A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n156 ) , .A2( u0_u14_u7_n163 ) );
  NAND2_X1 u0_u14_u7_U69 (.A2( u0_u14_X_46 ) , .A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n125 ) );
  OAI222_X1 u0_u14_u7_U7 (.C2( u0_u14_u7_n101 ) , .B2( u0_u14_u7_n111 ) , .A1( u0_u14_u7_n113 ) , .C1( u0_u14_u7_n146 ) , .A2( u0_u14_u7_n162 ) , .B1( u0_u14_u7_n164 ) , .ZN( u0_u14_u7_n94 ) );
  AND2_X1 u0_u14_u7_U70 (.A2( u0_u14_X_43 ) , .A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n96 ) );
  AND2_X1 u0_u14_u7_U71 (.A2( u0_u14_X_45 ) , .A1( u0_u14_X_48 ) , .ZN( u0_u14_u7_n102 ) );
  AND2_X1 u0_u14_u7_U72 (.A1( u0_u14_X_48 ) , .A2( u0_u14_u7_n166 ) , .ZN( u0_u14_u7_n93 ) );
  INV_X1 u0_u14_u7_U73 (.A( u0_u14_X_46 ) , .ZN( u0_u14_u7_n163 ) );
  AND2_X1 u0_u14_u7_U74 (.A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n100 ) , .A2( u0_u14_u7_n167 ) );
  INV_X1 u0_u14_u7_U75 (.A( u0_u14_X_43 ) , .ZN( u0_u14_u7_n167 ) );
  INV_X1 u0_u14_u7_U76 (.A( u0_u14_X_45 ) , .ZN( u0_u14_u7_n166 ) );
  NAND4_X1 u0_u14_u7_U77 (.ZN( u0_out14_27 ) , .A4( u0_u14_u7_n118 ) , .A3( u0_u14_u7_n119 ) , .A2( u0_u14_u7_n120 ) , .A1( u0_u14_u7_n121 ) );
  OAI21_X1 u0_u14_u7_U78 (.ZN( u0_u14_u7_n121 ) , .B2( u0_u14_u7_n145 ) , .A( u0_u14_u7_n150 ) , .B1( u0_u14_u7_n174 ) );
  OAI21_X1 u0_u14_u7_U79 (.ZN( u0_u14_u7_n120 ) , .A( u0_u14_u7_n161 ) , .B2( u0_u14_u7_n170 ) , .B1( u0_u14_u7_n179 ) );
  INV_X1 u0_u14_u7_U8 (.A( u0_u14_u7_n133 ) , .ZN( u0_u14_u7_n176 ) );
  NAND4_X1 u0_u14_u7_U80 (.ZN( u0_out14_21 ) , .A4( u0_u14_u7_n157 ) , .A3( u0_u14_u7_n158 ) , .A2( u0_u14_u7_n159 ) , .A1( u0_u14_u7_n160 ) );
  OAI21_X1 u0_u14_u7_U81 (.B1( u0_u14_u7_n145 ) , .ZN( u0_u14_u7_n160 ) , .A( u0_u14_u7_n161 ) , .B2( u0_u14_u7_n177 ) );
  OAI21_X1 u0_u14_u7_U82 (.ZN( u0_u14_u7_n159 ) , .A( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n171 ) , .B1( u0_u14_u7_n174 ) );
  NAND4_X1 u0_u14_u7_U83 (.ZN( u0_out14_15 ) , .A4( u0_u14_u7_n142 ) , .A3( u0_u14_u7_n143 ) , .A2( u0_u14_u7_n144 ) , .A1( u0_u14_u7_n178 ) );
  OR2_X1 u0_u14_u7_U84 (.A2( u0_u14_u7_n125 ) , .A1( u0_u14_u7_n129 ) , .ZN( u0_u14_u7_n144 ) );
  AOI22_X1 u0_u14_u7_U85 (.A2( u0_u14_u7_n126 ) , .ZN( u0_u14_u7_n143 ) , .B2( u0_u14_u7_n165 ) , .B1( u0_u14_u7_n173 ) , .A1( u0_u14_u7_n174 ) );
  NAND4_X1 u0_u14_u7_U86 (.ZN( u0_out14_5 ) , .A4( u0_u14_u7_n108 ) , .A3( u0_u14_u7_n109 ) , .A1( u0_u14_u7_n116 ) , .A2( u0_u14_u7_n123 ) );
  AOI22_X1 u0_u14_u7_U87 (.ZN( u0_u14_u7_n109 ) , .A2( u0_u14_u7_n126 ) , .B2( u0_u14_u7_n145 ) , .B1( u0_u14_u7_n156 ) , .A1( u0_u14_u7_n171 ) );
  NOR4_X1 u0_u14_u7_U88 (.A4( u0_u14_u7_n104 ) , .A3( u0_u14_u7_n105 ) , .A2( u0_u14_u7_n106 ) , .A1( u0_u14_u7_n107 ) , .ZN( u0_u14_u7_n108 ) );
  NAND2_X1 u0_u14_u7_U89 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n148 ) , .A2( u0_u14_u7_n95 ) );
  OAI221_X1 u0_u14_u7_U9 (.C1( u0_u14_u7_n101 ) , .C2( u0_u14_u7_n147 ) , .ZN( u0_u14_u7_n155 ) , .B2( u0_u14_u7_n162 ) , .A( u0_u14_u7_n91 ) , .B1( u0_u14_u7_n92 ) );
  NAND2_X1 u0_u14_u7_U90 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n113 ) , .A2( u0_u14_u7_n93 ) );
  NAND2_X1 u0_u14_u7_U91 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n138 ) , .A2( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U92 (.A1( u0_u14_u7_n100 ) , .A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n129 ) );
  OAI211_X1 u0_u14_u7_U93 (.B( u0_u14_u7_n122 ) , .A( u0_u14_u7_n123 ) , .C2( u0_u14_u7_n124 ) , .ZN( u0_u14_u7_n154 ) , .C1( u0_u14_u7_n162 ) );
  AOI222_X1 u0_u14_u7_U94 (.ZN( u0_u14_u7_n122 ) , .C2( u0_u14_u7_n126 ) , .C1( u0_u14_u7_n145 ) , .B1( u0_u14_u7_n161 ) , .A2( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n170 ) , .A1( u0_u14_u7_n176 ) );
  NAND3_X1 u0_u14_u7_U95 (.A3( u0_u14_u7_n146 ) , .A2( u0_u14_u7_n147 ) , .A1( u0_u14_u7_n148 ) , .ZN( u0_u14_u7_n151 ) );
  NAND3_X1 u0_u14_u7_U96 (.A3( u0_u14_u7_n131 ) , .A2( u0_u14_u7_n132 ) , .A1( u0_u14_u7_n133 ) , .ZN( u0_u14_u7_n135 ) );
  NAND2_X1 u0_uk_U125 (.A1( u0_uk_K_r0_52 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n856 ) );
  NAND2_X1 u0_uk_U171 (.A1( u0_key_r_18 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n889 ) );
  OAI22_X1 u0_uk_U236 (.ZN( u0_K15_39 ) , .A1( u0_uk_n128 ) , .B2( u0_uk_n22 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n40 ) );
  OAI22_X1 u0_uk_U244 (.ZN( u0_K15_44 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n22 ) , .A2( u0_uk_n4 ) );
  OAI21_X1 u0_uk_U245 (.ZN( u0_K15_48 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n34 ) , .A( u0_uk_n914 ) );
  NAND2_X1 u0_uk_U246 (.A1( u0_uk_K_r13_35 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n914 ) );
  OAI22_X1 u0_uk_U320 (.ZN( u0_K15_46 ) , .B2( u0_uk_n13 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n40 ) );
  OAI22_X1 u0_uk_U360 (.ZN( u0_K15_40 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n41 ) , .B2( u0_uk_n9 ) );
  OAI22_X1 u0_uk_U454 (.ZN( u0_K15_37 ) , .B2( u0_uk_n12 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n39 ) );
  INV_X1 u0_uk_U562 (.ZN( u0_K15_38 ) , .A( u0_uk_n916 ) );
  INV_X1 u0_uk_U660 (.ZN( u0_K15_43 ) , .A( u0_uk_n915 ) );
  AOI22_X1 u0_uk_U661 (.A2( u0_uk_K_r13_2 ) , .B2( u0_uk_K_r13_23 ) , .A1( u0_uk_n163 ) , .ZN( u0_uk_n915 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U726 (.ZN( u0_K15_42 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n3 ) , .B2( u0_uk_n9 ) );
  NAND2_X1 u0_uk_U763 (.A1( u0_uk_K_r9_5 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n998 ) );
  OAI22_X1 u0_uk_U88 (.ZN( u0_K15_41 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n23 ) , .A2( u0_uk_n5 ) );
  OAI22_X1 u0_uk_U886 (.ZN( u0_K15_45 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n21 ) , .A2( u0_uk_n3 ) );
  XOR2_X1 u1_U103 (.B( u1_L0_13 ) , .Z( u1_N44 ) , .A( u1_out1_13 ) );
  XOR2_X1 u1_U13 (.Z( u1_N9 ) , .B( u1_desIn_r_12 ) , .A( u1_out0_10 ) );
  XOR2_X1 u1_U131 (.B( u1_L11_31 ) , .Z( u1_N414 ) , .A( u1_out12_31 ) );
  XOR2_X1 u1_U134 (.B( u1_L11_28 ) , .Z( u1_N411 ) , .A( u1_out12_28 ) );
  XOR2_X1 u1_U137 (.B( u1_L11_26 ) , .Z( u1_N409 ) , .A( u1_out12_26 ) );
  XOR2_X1 u1_U140 (.B( u1_L11_23 ) , .Z( u1_N406 ) , .A( u1_out12_23 ) );
  XOR2_X1 u1_U143 (.B( u1_L11_20 ) , .Z( u1_N403 ) , .A( u1_out12_20 ) );
  XOR2_X1 u1_U145 (.B( u1_L11_18 ) , .Z( u1_N401 ) , .A( u1_out12_18 ) );
  XOR2_X1 u1_U146 (.B( u1_L11_17 ) , .Z( u1_N400 ) , .A( u1_out12_17 ) );
  XOR2_X1 u1_U152 (.B( u1_L11_13 ) , .Z( u1_N396 ) , .A( u1_out12_13 ) );
  XOR2_X1 u1_U155 (.B( u1_L11_10 ) , .Z( u1_N393 ) , .A( u1_out12_10 ) );
  XOR2_X1 u1_U156 (.B( u1_L11_9 ) , .Z( u1_N392 ) , .A( u1_out12_9 ) );
  XOR2_X1 u1_U164 (.B( u1_L11_2 ) , .Z( u1_N385 ) , .A( u1_out12_2 ) );
  XOR2_X1 u1_U165 (.B( u1_L11_1 ) , .Z( u1_N384 ) , .A( u1_out12_1 ) );
  XOR2_X1 u1_U181 (.B( u1_L0_6 ) , .Z( u1_N37 ) , .A( u1_out1_6 ) );
  XOR2_X1 u1_U202 (.B( u1_L9_31 ) , .Z( u1_N350 ) , .A( u1_out10_31 ) );
  XOR2_X1 u1_U204 (.B( u1_L9_30 ) , .Z( u1_N349 ) , .A( u1_out10_30 ) );
  XOR2_X1 u1_U205 (.B( u1_L9_29 ) , .Z( u1_N348 ) , .A( u1_out10_29 ) );
  XOR2_X1 u1_U206 (.B( u1_L9_28 ) , .Z( u1_N347 ) , .A( u1_out10_28 ) );
  XOR2_X1 u1_U210 (.B( u1_L9_24 ) , .Z( u1_N343 ) , .A( u1_out10_24 ) );
  XOR2_X1 u1_U211 (.B( u1_L9_23 ) , .Z( u1_N342 ) , .A( u1_out10_23 ) );
  XOR2_X1 u1_U216 (.B( u1_L9_19 ) , .Z( u1_N338 ) , .A( u1_out10_19 ) );
  XOR2_X1 u1_U217 (.B( u1_L9_18 ) , .Z( u1_N337 ) , .A( u1_out10_18 ) );
  XOR2_X1 u1_U218 (.B( u1_L9_17 ) , .Z( u1_N336 ) , .A( u1_out10_17 ) );
  XOR2_X1 u1_U219 (.B( u1_L9_16 ) , .Z( u1_N335 ) , .A( u1_out10_16 ) );
  XOR2_X1 u1_U222 (.B( u1_L9_13 ) , .Z( u1_N332 ) , .A( u1_out10_13 ) );
  XOR2_X1 u1_U224 (.B( u1_L9_11 ) , .Z( u1_N330 ) , .A( u1_out10_11 ) );
  XOR2_X1 u1_U225 (.B( u1_L0_2 ) , .Z( u1_N33 ) , .A( u1_out1_2 ) );
  XOR2_X1 u1_U227 (.B( u1_L9_9 ) , .Z( u1_N328 ) , .A( u1_out10_9 ) );
  XOR2_X1 u1_U230 (.B( u1_L9_6 ) , .Z( u1_N325 ) , .A( u1_out10_6 ) );
  XOR2_X1 u1_U232 (.B( u1_L9_4 ) , .Z( u1_N323 ) , .A( u1_out10_4 ) );
  XOR2_X1 u1_U234 (.B( u1_L9_2 ) , .Z( u1_N321 ) , .A( u1_out10_2 ) );
  XOR2_X1 u1_U238 (.B( u1_L8_31 ) , .Z( u1_N318 ) , .A( u1_out9_31 ) );
  XOR2_X1 u1_U239 (.B( u1_L8_30 ) , .Z( u1_N317 ) , .A( u1_out9_30 ) );
  XOR2_X1 u1_U24 (.Z( u1_N8 ) , .B( u1_desIn_r_4 ) , .A( u1_out0_9 ) );
  XOR2_X1 u1_U241 (.B( u1_L8_28 ) , .Z( u1_N315 ) , .A( u1_out9_28 ) );
  XOR2_X1 u1_U245 (.B( u1_L8_24 ) , .Z( u1_N311 ) , .A( u1_out9_24 ) );
  XOR2_X1 u1_U246 (.B( u1_L8_23 ) , .Z( u1_N310 ) , .A( u1_out9_23 ) );
  XOR2_X1 u1_U252 (.B( u1_L8_18 ) , .Z( u1_N305 ) , .A( u1_out9_18 ) );
  XOR2_X1 u1_U253 (.B( u1_L8_17 ) , .Z( u1_N304 ) , .A( u1_out9_17 ) );
  XOR2_X1 u1_U254 (.B( u1_L8_16 ) , .Z( u1_N303 ) , .A( u1_out9_16 ) );
  XOR2_X1 u1_U257 (.B( u1_L8_13 ) , .Z( u1_N300 ) , .A( u1_out9_13 ) );
  XOR2_X1 u1_U258 (.Z( u1_N30 ) , .B( u1_desIn_r_48 ) , .A( u1_out0_31 ) );
  XOR2_X1 u1_U263 (.B( u1_L8_9 ) , .Z( u1_N296 ) , .A( u1_out9_9 ) );
  XOR2_X1 u1_U266 (.B( u1_L8_6 ) , .Z( u1_N293 ) , .A( u1_out9_6 ) );
  XOR2_X1 u1_U270 (.Z( u1_N29 ) , .B( u1_desIn_r_40 ) , .A( u1_out0_30 ) );
  XOR2_X1 u1_U271 (.B( u1_L8_2 ) , .Z( u1_N289 ) , .A( u1_out9_2 ) );
  XOR2_X1 u1_U292 (.Z( u1_N27 ) , .B( u1_desIn_r_24 ) , .A( u1_out0_28 ) );
  XOR2_X1 u1_U314 (.Z( u1_N25 ) , .B( u1_desIn_r_8 ) , .A( u1_out0_26 ) );
  XOR2_X1 u1_U336 (.Z( u1_N23 ) , .B( u1_desIn_r_58 ) , .A( u1_out0_24 ) );
  XOR2_X1 u1_U347 (.Z( u1_N22 ) , .B( u1_desIn_r_50 ) , .A( u1_out0_23 ) );
  XOR2_X1 u1_U381 (.Z( u1_N19 ) , .B( u1_desIn_r_26 ) , .A( u1_out0_20 ) );
  XOR2_X1 u1_U403 (.Z( u1_N17 ) , .B( u1_desIn_r_10 ) , .A( u1_out0_18 ) );
  XOR2_X1 u1_U414 (.Z( u1_N16 ) , .B( u1_desIn_r_2 ) , .A( u1_out0_17 ) );
  XOR2_X1 u1_U419 (.B( u1_L3_28 ) , .Z( u1_N155 ) , .A( u1_out4_28 ) );
  XOR2_X1 u1_U425 (.Z( u1_N15 ) , .B( u1_desIn_r_60 ) , .A( u1_out0_16 ) );
  XOR2_X1 u1_U430 (.B( u1_L3_18 ) , .Z( u1_N145 ) , .A( u1_out4_18 ) );
  XOR2_X1 u1_U435 (.B( u1_L3_13 ) , .Z( u1_N140 ) , .A( u1_out4_13 ) );
  XOR2_X1 u1_U44 (.B( u1_L0_30 ) , .Z( u1_N61 ) , .A( u1_out1_30 ) );
  XOR2_X1 u1_U448 (.B( u1_L3_2 ) , .Z( u1_N129 ) , .A( u1_out4_2 ) );
  XOR2_X1 u1_U458 (.Z( u1_N12 ) , .B( u1_desIn_r_36 ) , .A( u1_out0_13 ) );
  XOR2_X1 u1_U47 (.B( u1_L0_28 ) , .Z( u1_N59 ) , .A( u1_out1_28 ) );
  XOR2_X1 u1_U481 (.Z( u1_N1 ) , .B( u1_desIn_r_14 ) , .A( u1_out0_2 ) );
  XOR2_X1 u1_U482 (.Z( u1_N0 ) , .B( u1_desIn_r_6 ) , .A( u1_out0_1 ) );
  XOR2_X1 u1_U486 (.Z( u1_FP_6 ) , .B( u1_L14_6 ) , .A( u1_out15_6 ) );
  XOR2_X1 u1_U492 (.Z( u1_FP_30 ) , .B( u1_L14_30 ) , .A( u1_out15_30 ) );
  XOR2_X1 u1_U499 (.Z( u1_FP_24 ) , .B( u1_L14_24 ) , .A( u1_out15_24 ) );
  XOR2_X1 u1_U508 (.Z( u1_FP_16 ) , .B( u1_L14_16 ) , .A( u1_out15_16 ) );
  XOR2_X1 u1_U51 (.B( u1_L0_24 ) , .Z( u1_N55 ) , .A( u1_out1_24 ) );
  XOR2_X1 u1_U57 (.Z( u1_N5 ) , .B( u1_desIn_r_46 ) , .A( u1_out0_6 ) );
  XOR2_X1 u1_U58 (.B( u1_L0_18 ) , .Z( u1_N49 ) , .A( u1_out1_18 ) );
  XOR2_X1 u1_U70 (.B( u1_L0_16 ) , .Z( u1_N47 ) , .A( u1_out1_16 ) );
  XOR2_X1 u1_u0_U1 (.B( u1_K1_9 ) , .A( u1_desIn_r_47 ) , .Z( u1_u0_X_9 ) );
  XOR2_X1 u1_u0_U16 (.B( u1_K1_3 ) , .A( u1_desIn_r_15 ) , .Z( u1_u0_X_3 ) );
  XOR2_X1 u1_u0_U2 (.B( u1_K1_8 ) , .A( u1_desIn_r_39 ) , .Z( u1_u0_X_8 ) );
  XOR2_X1 u1_u0_U27 (.B( u1_K1_2 ) , .A( u1_desIn_r_7 ) , .Z( u1_u0_X_2 ) );
  XOR2_X1 u1_u0_U3 (.B( u1_K1_7 ) , .A( u1_desIn_r_31 ) , .Z( u1_u0_X_7 ) );
  XOR2_X1 u1_u0_U33 (.B( u1_K1_24 ) , .A( u1_desIn_r_3 ) , .Z( u1_u0_X_24 ) );
  XOR2_X1 u1_u0_U34 (.B( u1_K1_23 ) , .A( u1_desIn_r_61 ) , .Z( u1_u0_X_23 ) );
  XOR2_X1 u1_u0_U35 (.B( u1_K1_22 ) , .A( u1_desIn_r_53 ) , .Z( u1_u0_X_22 ) );
  XOR2_X1 u1_u0_U36 (.B( u1_K1_21 ) , .A( u1_desIn_r_45 ) , .Z( u1_u0_X_21 ) );
  XOR2_X1 u1_u0_U37 (.B( u1_K1_20 ) , .A( u1_desIn_r_37 ) , .Z( u1_u0_X_20 ) );
  XOR2_X1 u1_u0_U38 (.B( u1_K1_1 ) , .A( u1_desIn_r_57 ) , .Z( u1_u0_X_1 ) );
  XOR2_X1 u1_u0_U39 (.B( u1_K1_19 ) , .A( u1_desIn_r_29 ) , .Z( u1_u0_X_19 ) );
  XOR2_X1 u1_u0_U4 (.B( u1_K1_6 ) , .A( u1_desIn_r_39 ) , .Z( u1_u0_X_6 ) );
  XOR2_X1 u1_u0_U40 (.B( u1_K1_18 ) , .A( u1_desIn_r_37 ) , .Z( u1_u0_X_18 ) );
  XOR2_X1 u1_u0_U41 (.B( u1_K1_17 ) , .A( u1_desIn_r_29 ) , .Z( u1_u0_X_17 ) );
  XOR2_X1 u1_u0_U42 (.B( u1_K1_16 ) , .A( u1_desIn_r_21 ) , .Z( u1_u0_X_16 ) );
  XOR2_X1 u1_u0_U43 (.B( u1_K1_15 ) , .A( u1_desIn_r_13 ) , .Z( u1_u0_X_15 ) );
  XOR2_X1 u1_u0_U44 (.B( u1_K1_14 ) , .A( u1_desIn_r_5 ) , .Z( u1_u0_X_14 ) );
  XOR2_X1 u1_u0_U45 (.B( u1_K1_13 ) , .A( u1_desIn_r_63 ) , .Z( u1_u0_X_13 ) );
  XOR2_X1 u1_u0_U46 (.B( u1_K1_12 ) , .A( u1_desIn_r_5 ) , .Z( u1_u0_X_12 ) );
  XOR2_X1 u1_u0_U47 (.B( u1_K1_11 ) , .A( u1_desIn_r_63 ) , .Z( u1_u0_X_11 ) );
  XOR2_X1 u1_u0_U48 (.B( u1_K1_10 ) , .A( u1_desIn_r_55 ) , .Z( u1_u0_X_10 ) );
  XOR2_X1 u1_u0_U5 (.B( u1_K1_5 ) , .A( u1_desIn_r_31 ) , .Z( u1_u0_X_5 ) );
  XOR2_X1 u1_u0_U6 (.B( u1_K1_4 ) , .A( u1_desIn_r_23 ) , .Z( u1_u0_X_4 ) );
  NAND2_X1 u1_u0_u0_U10 (.ZN( u1_u0_u0_n113 ) , .A1( u1_u0_u0_n139 ) , .A2( u1_u0_u0_n149 ) );
  AND3_X1 u1_u0_u0_U11 (.A2( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n127 ) , .A3( u1_u0_u0_n130 ) , .A1( u1_u0_u0_n148 ) );
  AND2_X1 u1_u0_u0_U12 (.ZN( u1_u0_u0_n107 ) , .A1( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n140 ) );
  AND2_X1 u1_u0_u0_U13 (.A2( u1_u0_u0_n129 ) , .A1( u1_u0_u0_n130 ) , .ZN( u1_u0_u0_n151 ) );
  AND2_X1 u1_u0_u0_U14 (.A1( u1_u0_u0_n108 ) , .A2( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U15 (.A( u1_u0_u0_n143 ) , .ZN( u1_u0_u0_n173 ) );
  NOR2_X1 u1_u0_u0_U16 (.A2( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n147 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U17 (.ZN( u1_u0_u0_n172 ) , .A( u1_u0_u0_n88 ) );
  OAI222_X1 u1_u0_u0_U18 (.C1( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n125 ) , .B2( u1_u0_u0_n128 ) , .B1( u1_u0_u0_n144 ) , .A2( u1_u0_u0_n158 ) , .C2( u1_u0_u0_n161 ) , .ZN( u1_u0_u0_n88 ) );
  AOI21_X1 u1_u0_u0_U19 (.B1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n132 ) , .A( u1_u0_u0_n165 ) , .B2( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U20 (.A( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n165 ) );
  OAI22_X1 u1_u0_u0_U21 (.B1( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n126 ) , .A1( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n146 ) , .B2( u1_u0_u0_n147 ) );
  OAI22_X1 u1_u0_u0_U22 (.B1( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n147 ) , .A2( u1_u0_u0_n90 ) , .ZN( u1_u0_u0_n91 ) );
  AND3_X1 u1_u0_u0_U23 (.A3( u1_u0_u0_n121 ) , .A2( u1_u0_u0_n125 ) , .A1( u1_u0_u0_n148 ) , .ZN( u1_u0_u0_n90 ) );
  INV_X1 u1_u0_u0_U24 (.A( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n161 ) );
  AOI22_X1 u1_u0_u0_U25 (.B2( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n110 ) , .ZN( u1_u0_u0_n111 ) , .B1( u1_u0_u0_n118 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U26 (.A( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U27 (.B1( u1_u0_u0_n127 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n96 ) );
  AOI21_X1 u1_u0_u0_U28 (.ZN( u1_u0_u0_n104 ) , .B1( u1_u0_u0_n107 ) , .B2( u1_u0_u0_n141 ) , .A( u1_u0_u0_n144 ) );
  NAND2_X1 u1_u0_u0_U29 (.A1( u1_u0_u0_n100 ) , .A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n125 ) );
  INV_X1 u1_u0_u0_U3 (.A( u1_u0_u0_n113 ) , .ZN( u1_u0_u0_n166 ) );
  NAND2_X1 u1_u0_u0_U30 (.A2( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n92 ) );
  NAND2_X1 u1_u0_u0_U31 (.A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n114 ) , .A1( u1_u0_u0_n92 ) );
  NOR2_X1 u1_u0_u0_U32 (.A1( u1_u0_u0_n120 ) , .ZN( u1_u0_u0_n143 ) , .A2( u1_u0_u0_n167 ) );
  OAI221_X1 u1_u0_u0_U33 (.C1( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n120 ) , .B1( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n141 ) , .C2( u1_u0_u0_n147 ) , .A( u1_u0_u0_n172 ) );
  AOI21_X1 u1_u0_u0_U34 (.ZN( u1_u0_u0_n116 ) , .B2( u1_u0_u0_n142 ) , .A( u1_u0_u0_n144 ) , .B1( u1_u0_u0_n166 ) );
  INV_X1 u1_u0_u0_U35 (.A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n160 ) );
  NAND2_X1 u1_u0_u0_U36 (.A2( u1_u0_u0_n102 ) , .A1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n149 ) );
  NAND2_X1 u1_u0_u0_U37 (.ZN( u1_u0_u0_n112 ) , .A2( u1_u0_u0_n92 ) , .A1( u1_u0_u0_n93 ) );
  OR3_X1 u1_u0_u0_U38 (.A3( u1_u0_u0_n152 ) , .A2( u1_u0_u0_n153 ) , .A1( u1_u0_u0_n154 ) , .ZN( u1_u0_u0_n155 ) );
  AOI21_X1 u1_u0_u0_U39 (.B2( u1_u0_u0_n150 ) , .B1( u1_u0_u0_n151 ) , .ZN( u1_u0_u0_n152 ) , .A( u1_u0_u0_n158 ) );
  NOR2_X1 u1_u0_u0_U4 (.A1( u1_u0_u0_n108 ) , .ZN( u1_u0_u0_n123 ) , .A2( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U40 (.A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n145 ) , .B1( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n154 ) );
  AOI21_X1 u1_u0_u0_U41 (.A( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n148 ) , .B1( u1_u0_u0_n149 ) , .ZN( u1_u0_u0_n153 ) );
  INV_X1 u1_u0_u0_U42 (.ZN( u1_u0_u0_n171 ) , .A( u1_u0_u0_n99 ) );
  OAI211_X1 u1_u0_u0_U43 (.C2( u1_u0_u0_n140 ) , .C1( u1_u0_u0_n161 ) , .A( u1_u0_u0_n169 ) , .B( u1_u0_u0_n98 ) , .ZN( u1_u0_u0_n99 ) );
  AOI211_X1 u1_u0_u0_U44 (.C1( u1_u0_u0_n118 ) , .A( u1_u0_u0_n123 ) , .B( u1_u0_u0_n96 ) , .C2( u1_u0_u0_n97 ) , .ZN( u1_u0_u0_n98 ) );
  INV_X1 u1_u0_u0_U45 (.ZN( u1_u0_u0_n169 ) , .A( u1_u0_u0_n91 ) );
  NOR2_X1 u1_u0_u0_U46 (.A2( u1_u0_X_2 ) , .ZN( u1_u0_u0_n103 ) , .A1( u1_u0_u0_n164 ) );
  NOR2_X1 u1_u0_u0_U47 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n118 ) );
  NAND2_X1 u1_u0_u0_U48 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n144 ) );
  NOR2_X1 u1_u0_u0_U49 (.A2( u1_u0_X_5 ) , .ZN( u1_u0_u0_n136 ) , .A1( u1_u0_u0_n159 ) );
  AOI21_X1 u1_u0_u0_U5 (.B2( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n134 ) , .B1( u1_u0_u0_n151 ) , .A( u1_u0_u0_n158 ) );
  NAND2_X1 u1_u0_u0_U50 (.A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n159 ) );
  AND2_X1 u1_u0_u0_U51 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n102 ) );
  AND2_X1 u1_u0_u0_U52 (.A1( u1_u0_X_6 ) , .A2( u1_u0_u0_n162 ) , .ZN( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U53 (.A( u1_u0_X_4 ) , .ZN( u1_u0_u0_n159 ) );
  INV_X1 u1_u0_u0_U54 (.A( u1_u0_X_2 ) , .ZN( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U55 (.A( u1_u0_X_3 ) , .ZN( u1_u0_u0_n162 ) );
  INV_X1 u1_u0_u0_U56 (.A( u1_u0_u0_n126 ) , .ZN( u1_u0_u0_n168 ) );
  AOI211_X1 u1_u0_u0_U57 (.B( u1_u0_u0_n133 ) , .A( u1_u0_u0_n134 ) , .C2( u1_u0_u0_n135 ) , .C1( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n137 ) );
  OR4_X1 u1_u0_u0_U58 (.ZN( u1_out0_17 ) , .A4( u1_u0_u0_n122 ) , .A2( u1_u0_u0_n123 ) , .A1( u1_u0_u0_n124 ) , .A3( u1_u0_u0_n170 ) );
  AOI21_X1 u1_u0_u0_U59 (.B2( u1_u0_u0_n107 ) , .ZN( u1_u0_u0_n124 ) , .B1( u1_u0_u0_n128 ) , .A( u1_u0_u0_n161 ) );
  OAI21_X1 u1_u0_u0_U6 (.B1( u1_u0_u0_n150 ) , .B2( u1_u0_u0_n158 ) , .A( u1_u0_u0_n172 ) , .ZN( u1_u0_u0_n89 ) );
  INV_X1 u1_u0_u0_U60 (.A( u1_u0_u0_n111 ) , .ZN( u1_u0_u0_n170 ) );
  OR4_X1 u1_u0_u0_U61 (.ZN( u1_out0_31 ) , .A4( u1_u0_u0_n155 ) , .A2( u1_u0_u0_n156 ) , .A1( u1_u0_u0_n157 ) , .A3( u1_u0_u0_n173 ) );
  AOI21_X1 u1_u0_u0_U62 (.A( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n139 ) , .B1( u1_u0_u0_n140 ) , .ZN( u1_u0_u0_n157 ) );
  AOI21_X1 u1_u0_u0_U63 (.B2( u1_u0_u0_n141 ) , .B1( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n156 ) , .A( u1_u0_u0_n161 ) );
  INV_X1 u1_u0_u0_U64 (.ZN( u1_u0_u0_n174 ) , .A( u1_u0_u0_n89 ) );
  AOI211_X1 u1_u0_u0_U65 (.B( u1_u0_u0_n104 ) , .A( u1_u0_u0_n105 ) , .ZN( u1_u0_u0_n106 ) , .C2( u1_u0_u0_n113 ) , .C1( u1_u0_u0_n160 ) );
  AOI211_X1 u1_u0_u0_U66 (.B( u1_u0_u0_n115 ) , .A( u1_u0_u0_n116 ) , .C2( u1_u0_u0_n117 ) , .C1( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n119 ) );
  NAND2_X1 u1_u0_u0_U67 (.A2( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n121 ) , .A1( u1_u0_u0_n93 ) );
  NAND2_X1 u1_u0_u0_U68 (.A1( u1_u0_u0_n101 ) , .A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n150 ) );
  NOR2_X1 u1_u0_u0_U69 (.A2( u1_u0_X_1 ) , .A1( u1_u0_X_2 ) , .ZN( u1_u0_u0_n92 ) );
  AOI21_X1 u1_u0_u0_U7 (.B1( u1_u0_u0_n114 ) , .ZN( u1_u0_u0_n115 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n161 ) );
  NAND2_X1 u1_u0_u0_U70 (.A2( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n139 ) );
  NOR2_X1 u1_u0_u0_U71 (.A2( u1_u0_X_1 ) , .ZN( u1_u0_u0_n101 ) , .A1( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U72 (.A( u1_u0_X_1 ) , .ZN( u1_u0_u0_n164 ) );
  NAND2_X1 u1_u0_u0_U73 (.A1( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n128 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U74 (.A1( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n129 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U75 (.ZN( u1_u0_u0_n148 ) , .A1( u1_u0_u0_n93 ) , .A2( u1_u0_u0_n95 ) );
  OAI221_X1 u1_u0_u0_U76 (.C1( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n122 ) , .B2( u1_u0_u0_n127 ) , .A( u1_u0_u0_n143 ) , .B1( u1_u0_u0_n144 ) , .C2( u1_u0_u0_n147 ) );
  NOR2_X1 u1_u0_u0_U77 (.A1( u1_u0_u0_n163 ) , .A2( u1_u0_u0_n164 ) , .ZN( u1_u0_u0_n95 ) );
  AOI21_X1 u1_u0_u0_U78 (.B1( u1_u0_u0_n132 ) , .ZN( u1_u0_u0_n133 ) , .A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n166 ) );
  OAI22_X1 u1_u0_u0_U79 (.ZN( u1_u0_u0_n105 ) , .A2( u1_u0_u0_n132 ) , .B1( u1_u0_u0_n146 ) , .A1( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n161 ) );
  AND2_X1 u1_u0_u0_U8 (.A1( u1_u0_u0_n114 ) , .A2( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n146 ) );
  NAND2_X1 u1_u0_u0_U80 (.ZN( u1_u0_u0_n110 ) , .A2( u1_u0_u0_n132 ) , .A1( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U81 (.A( u1_u0_u0_n119 ) , .ZN( u1_u0_u0_n167 ) );
  NAND2_X1 u1_u0_u0_U82 (.A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U83 (.A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U84 (.ZN( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n92 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U85 (.ZN( u1_u0_u0_n142 ) , .A1( u1_u0_u0_n94 ) , .A2( u1_u0_u0_n95 ) );
  NOR2_X1 u1_u0_u0_U86 (.A2( u1_u0_X_6 ) , .ZN( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n162 ) );
  NOR2_X1 u1_u0_u0_U87 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n94 ) );
  NAND3_X1 u1_u0_u0_U88 (.ZN( u1_out0_23 ) , .A3( u1_u0_u0_n137 ) , .A1( u1_u0_u0_n168 ) , .A2( u1_u0_u0_n171 ) );
  NAND3_X1 u1_u0_u0_U89 (.A3( u1_u0_u0_n127 ) , .A2( u1_u0_u0_n128 ) , .ZN( u1_u0_u0_n135 ) , .A1( u1_u0_u0_n150 ) );
  AND2_X1 u1_u0_u0_U9 (.A1( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n141 ) , .A2( u1_u0_u0_n150 ) );
  NAND3_X1 u1_u0_u0_U90 (.ZN( u1_u0_u0_n117 ) , .A3( u1_u0_u0_n132 ) , .A2( u1_u0_u0_n139 ) , .A1( u1_u0_u0_n148 ) );
  NAND3_X1 u1_u0_u0_U91 (.ZN( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n114 ) , .A3( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n149 ) );
  NAND3_X1 u1_u0_u0_U92 (.ZN( u1_out0_9 ) , .A3( u1_u0_u0_n106 ) , .A2( u1_u0_u0_n171 ) , .A1( u1_u0_u0_n174 ) );
  NAND3_X1 u1_u0_u0_U93 (.A2( u1_u0_u0_n128 ) , .A1( u1_u0_u0_n132 ) , .A3( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n97 ) );
  AOI21_X1 u1_u0_u1_U10 (.B2( u1_u0_u1_n155 ) , .B1( u1_u0_u1_n156 ) , .ZN( u1_u0_u1_n157 ) , .A( u1_u0_u1_n174 ) );
  NAND3_X1 u1_u0_u1_U100 (.ZN( u1_u0_u1_n113 ) , .A1( u1_u0_u1_n120 ) , .A3( u1_u0_u1_n133 ) , .A2( u1_u0_u1_n155 ) );
  NAND2_X1 u1_u0_u1_U11 (.ZN( u1_u0_u1_n140 ) , .A2( u1_u0_u1_n150 ) , .A1( u1_u0_u1_n155 ) );
  NAND2_X1 u1_u0_u1_U12 (.A1( u1_u0_u1_n131 ) , .ZN( u1_u0_u1_n147 ) , .A2( u1_u0_u1_n153 ) );
  AOI22_X1 u1_u0_u1_U13 (.B2( u1_u0_u1_n136 ) , .A2( u1_u0_u1_n137 ) , .ZN( u1_u0_u1_n143 ) , .A1( u1_u0_u1_n171 ) , .B1( u1_u0_u1_n173 ) );
  INV_X1 u1_u0_u1_U14 (.A( u1_u0_u1_n147 ) , .ZN( u1_u0_u1_n181 ) );
  INV_X1 u1_u0_u1_U15 (.A( u1_u0_u1_n139 ) , .ZN( u1_u0_u1_n174 ) );
  OR4_X1 u1_u0_u1_U16 (.A4( u1_u0_u1_n106 ) , .A3( u1_u0_u1_n107 ) , .ZN( u1_u0_u1_n108 ) , .A1( u1_u0_u1_n117 ) , .A2( u1_u0_u1_n184 ) );
  AOI21_X1 u1_u0_u1_U17 (.ZN( u1_u0_u1_n106 ) , .A( u1_u0_u1_n112 ) , .B1( u1_u0_u1_n154 ) , .B2( u1_u0_u1_n156 ) );
  AOI21_X1 u1_u0_u1_U18 (.ZN( u1_u0_u1_n107 ) , .B1( u1_u0_u1_n134 ) , .B2( u1_u0_u1_n149 ) , .A( u1_u0_u1_n174 ) );
  INV_X1 u1_u0_u1_U19 (.A( u1_u0_u1_n101 ) , .ZN( u1_u0_u1_n184 ) );
  INV_X1 u1_u0_u1_U20 (.A( u1_u0_u1_n112 ) , .ZN( u1_u0_u1_n171 ) );
  NAND2_X1 u1_u0_u1_U21 (.ZN( u1_u0_u1_n141 ) , .A1( u1_u0_u1_n153 ) , .A2( u1_u0_u1_n156 ) );
  AND2_X1 u1_u0_u1_U22 (.A1( u1_u0_u1_n123 ) , .ZN( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n161 ) );
  NAND2_X1 u1_u0_u1_U23 (.A2( u1_u0_u1_n115 ) , .A1( u1_u0_u1_n116 ) , .ZN( u1_u0_u1_n148 ) );
  NAND2_X1 u1_u0_u1_U24 (.A2( u1_u0_u1_n133 ) , .A1( u1_u0_u1_n135 ) , .ZN( u1_u0_u1_n159 ) );
  NAND2_X1 u1_u0_u1_U25 (.A2( u1_u0_u1_n115 ) , .A1( u1_u0_u1_n120 ) , .ZN( u1_u0_u1_n132 ) );
  INV_X1 u1_u0_u1_U26 (.A( u1_u0_u1_n154 ) , .ZN( u1_u0_u1_n178 ) );
  INV_X1 u1_u0_u1_U27 (.A( u1_u0_u1_n151 ) , .ZN( u1_u0_u1_n183 ) );
  AND2_X1 u1_u0_u1_U28 (.A1( u1_u0_u1_n129 ) , .A2( u1_u0_u1_n133 ) , .ZN( u1_u0_u1_n149 ) );
  INV_X1 u1_u0_u1_U29 (.A( u1_u0_u1_n131 ) , .ZN( u1_u0_u1_n180 ) );
  INV_X1 u1_u0_u1_U3 (.A( u1_u0_u1_n159 ) , .ZN( u1_u0_u1_n182 ) );
  AOI221_X1 u1_u0_u1_U30 (.B1( u1_u0_u1_n140 ) , .ZN( u1_u0_u1_n167 ) , .B2( u1_u0_u1_n172 ) , .C2( u1_u0_u1_n175 ) , .C1( u1_u0_u1_n178 ) , .A( u1_u0_u1_n188 ) );
  INV_X1 u1_u0_u1_U31 (.ZN( u1_u0_u1_n188 ) , .A( u1_u0_u1_n97 ) );
  AOI211_X1 u1_u0_u1_U32 (.A( u1_u0_u1_n118 ) , .C1( u1_u0_u1_n132 ) , .C2( u1_u0_u1_n139 ) , .B( u1_u0_u1_n96 ) , .ZN( u1_u0_u1_n97 ) );
  AOI21_X1 u1_u0_u1_U33 (.B2( u1_u0_u1_n121 ) , .B1( u1_u0_u1_n135 ) , .A( u1_u0_u1_n152 ) , .ZN( u1_u0_u1_n96 ) );
  OAI221_X1 u1_u0_u1_U34 (.A( u1_u0_u1_n119 ) , .C2( u1_u0_u1_n129 ) , .ZN( u1_u0_u1_n138 ) , .B2( u1_u0_u1_n152 ) , .C1( u1_u0_u1_n174 ) , .B1( u1_u0_u1_n187 ) );
  INV_X1 u1_u0_u1_U35 (.A( u1_u0_u1_n148 ) , .ZN( u1_u0_u1_n187 ) );
  AOI211_X1 u1_u0_u1_U36 (.B( u1_u0_u1_n117 ) , .A( u1_u0_u1_n118 ) , .ZN( u1_u0_u1_n119 ) , .C2( u1_u0_u1_n146 ) , .C1( u1_u0_u1_n159 ) );
  NOR2_X1 u1_u0_u1_U37 (.A1( u1_u0_u1_n168 ) , .A2( u1_u0_u1_n176 ) , .ZN( u1_u0_u1_n98 ) );
  AOI211_X1 u1_u0_u1_U38 (.B( u1_u0_u1_n162 ) , .A( u1_u0_u1_n163 ) , .C2( u1_u0_u1_n164 ) , .ZN( u1_u0_u1_n165 ) , .C1( u1_u0_u1_n171 ) );
  AOI21_X1 u1_u0_u1_U39 (.A( u1_u0_u1_n160 ) , .B2( u1_u0_u1_n161 ) , .ZN( u1_u0_u1_n162 ) , .B1( u1_u0_u1_n182 ) );
  AOI221_X1 u1_u0_u1_U4 (.A( u1_u0_u1_n138 ) , .C2( u1_u0_u1_n139 ) , .C1( u1_u0_u1_n140 ) , .B2( u1_u0_u1_n141 ) , .ZN( u1_u0_u1_n142 ) , .B1( u1_u0_u1_n175 ) );
  OR2_X1 u1_u0_u1_U40 (.A2( u1_u0_u1_n157 ) , .A1( u1_u0_u1_n158 ) , .ZN( u1_u0_u1_n163 ) );
  OAI21_X1 u1_u0_u1_U41 (.B2( u1_u0_u1_n123 ) , .ZN( u1_u0_u1_n145 ) , .B1( u1_u0_u1_n160 ) , .A( u1_u0_u1_n185 ) );
  INV_X1 u1_u0_u1_U42 (.A( u1_u0_u1_n122 ) , .ZN( u1_u0_u1_n185 ) );
  AOI21_X1 u1_u0_u1_U43 (.B2( u1_u0_u1_n120 ) , .B1( u1_u0_u1_n121 ) , .ZN( u1_u0_u1_n122 ) , .A( u1_u0_u1_n128 ) );
  NAND2_X1 u1_u0_u1_U44 (.A1( u1_u0_u1_n128 ) , .ZN( u1_u0_u1_n146 ) , .A2( u1_u0_u1_n160 ) );
  NAND2_X1 u1_u0_u1_U45 (.A2( u1_u0_u1_n112 ) , .ZN( u1_u0_u1_n139 ) , .A1( u1_u0_u1_n152 ) );
  NAND2_X1 u1_u0_u1_U46 (.A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n156 ) , .A2( u1_u0_u1_n99 ) );
  NOR2_X1 u1_u0_u1_U47 (.ZN( u1_u0_u1_n117 ) , .A1( u1_u0_u1_n121 ) , .A2( u1_u0_u1_n160 ) );
  AOI21_X1 u1_u0_u1_U48 (.A( u1_u0_u1_n128 ) , .B2( u1_u0_u1_n129 ) , .ZN( u1_u0_u1_n130 ) , .B1( u1_u0_u1_n150 ) );
  NAND2_X1 u1_u0_u1_U49 (.ZN( u1_u0_u1_n112 ) , .A1( u1_u0_u1_n169 ) , .A2( u1_u0_u1_n170 ) );
  AOI211_X1 u1_u0_u1_U5 (.ZN( u1_u0_u1_n124 ) , .A( u1_u0_u1_n138 ) , .C2( u1_u0_u1_n139 ) , .B( u1_u0_u1_n145 ) , .C1( u1_u0_u1_n147 ) );
  NAND2_X1 u1_u0_u1_U50 (.ZN( u1_u0_u1_n129 ) , .A2( u1_u0_u1_n95 ) , .A1( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U51 (.A1( u1_u0_u1_n102 ) , .ZN( u1_u0_u1_n154 ) , .A2( u1_u0_u1_n99 ) );
  NAND2_X1 u1_u0_u1_U52 (.A2( u1_u0_u1_n100 ) , .ZN( u1_u0_u1_n135 ) , .A1( u1_u0_u1_n99 ) );
  AOI21_X1 u1_u0_u1_U53 (.A( u1_u0_u1_n152 ) , .B2( u1_u0_u1_n153 ) , .B1( u1_u0_u1_n154 ) , .ZN( u1_u0_u1_n158 ) );
  INV_X1 u1_u0_u1_U54 (.A( u1_u0_u1_n160 ) , .ZN( u1_u0_u1_n175 ) );
  NAND2_X1 u1_u0_u1_U55 (.A1( u1_u0_u1_n100 ) , .ZN( u1_u0_u1_n116 ) , .A2( u1_u0_u1_n95 ) );
  NAND2_X1 u1_u0_u1_U56 (.A1( u1_u0_u1_n102 ) , .ZN( u1_u0_u1_n131 ) , .A2( u1_u0_u1_n95 ) );
  NAND2_X1 u1_u0_u1_U57 (.A2( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n121 ) , .A1( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U58 (.A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n153 ) , .A2( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U59 (.A2( u1_u0_u1_n104 ) , .A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n133 ) );
  AOI22_X1 u1_u0_u1_U6 (.B2( u1_u0_u1_n113 ) , .A2( u1_u0_u1_n114 ) , .ZN( u1_u0_u1_n125 ) , .A1( u1_u0_u1_n171 ) , .B1( u1_u0_u1_n173 ) );
  NAND2_X1 u1_u0_u1_U60 (.ZN( u1_u0_u1_n150 ) , .A2( u1_u0_u1_n98 ) , .A1( u1_u0_u1_n99 ) );
  NAND2_X1 u1_u0_u1_U61 (.A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n155 ) , .A2( u1_u0_u1_n95 ) );
  OAI21_X1 u1_u0_u1_U62 (.ZN( u1_u0_u1_n109 ) , .B1( u1_u0_u1_n129 ) , .B2( u1_u0_u1_n160 ) , .A( u1_u0_u1_n167 ) );
  NAND2_X1 u1_u0_u1_U63 (.A2( u1_u0_u1_n100 ) , .A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n120 ) );
  NAND2_X1 u1_u0_u1_U64 (.A1( u1_u0_u1_n102 ) , .A2( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n115 ) );
  NAND2_X1 u1_u0_u1_U65 (.A2( u1_u0_u1_n100 ) , .A1( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n151 ) );
  NAND2_X1 u1_u0_u1_U66 (.A2( u1_u0_u1_n103 ) , .A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n161 ) );
  INV_X1 u1_u0_u1_U67 (.A( u1_u0_u1_n152 ) , .ZN( u1_u0_u1_n173 ) );
  INV_X1 u1_u0_u1_U68 (.A( u1_u0_u1_n128 ) , .ZN( u1_u0_u1_n172 ) );
  NAND2_X1 u1_u0_u1_U69 (.A2( u1_u0_u1_n102 ) , .A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n123 ) );
  NAND2_X1 u1_u0_u1_U7 (.ZN( u1_u0_u1_n114 ) , .A1( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n156 ) );
  NOR2_X1 u1_u0_u1_U70 (.A2( u1_u0_X_7 ) , .A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n95 ) );
  NOR2_X1 u1_u0_u1_U71 (.A1( u1_u0_X_12 ) , .A2( u1_u0_X_9 ) , .ZN( u1_u0_u1_n100 ) );
  NOR2_X1 u1_u0_u1_U72 (.A2( u1_u0_X_8 ) , .A1( u1_u0_u1_n177 ) , .ZN( u1_u0_u1_n99 ) );
  NOR2_X1 u1_u0_u1_U73 (.A2( u1_u0_X_12 ) , .ZN( u1_u0_u1_n102 ) , .A1( u1_u0_u1_n176 ) );
  NOR2_X1 u1_u0_u1_U74 (.A2( u1_u0_X_9 ) , .ZN( u1_u0_u1_n105 ) , .A1( u1_u0_u1_n168 ) );
  NAND2_X1 u1_u0_u1_U75 (.A1( u1_u0_X_10 ) , .ZN( u1_u0_u1_n160 ) , .A2( u1_u0_u1_n169 ) );
  NAND2_X1 u1_u0_u1_U76 (.A2( u1_u0_X_10 ) , .A1( u1_u0_X_11 ) , .ZN( u1_u0_u1_n152 ) );
  NAND2_X1 u1_u0_u1_U77 (.A1( u1_u0_X_11 ) , .ZN( u1_u0_u1_n128 ) , .A2( u1_u0_u1_n170 ) );
  AND2_X1 u1_u0_u1_U78 (.A2( u1_u0_X_7 ) , .A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n104 ) );
  AND2_X1 u1_u0_u1_U79 (.A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n103 ) , .A2( u1_u0_u1_n177 ) );
  NOR2_X1 u1_u0_u1_U8 (.A1( u1_u0_u1_n112 ) , .A2( u1_u0_u1_n116 ) , .ZN( u1_u0_u1_n118 ) );
  INV_X1 u1_u0_u1_U80 (.A( u1_u0_X_10 ) , .ZN( u1_u0_u1_n170 ) );
  INV_X1 u1_u0_u1_U81 (.A( u1_u0_X_9 ) , .ZN( u1_u0_u1_n176 ) );
  INV_X1 u1_u0_u1_U82 (.A( u1_u0_X_11 ) , .ZN( u1_u0_u1_n169 ) );
  INV_X1 u1_u0_u1_U83 (.A( u1_u0_X_12 ) , .ZN( u1_u0_u1_n168 ) );
  INV_X1 u1_u0_u1_U84 (.A( u1_u0_X_7 ) , .ZN( u1_u0_u1_n177 ) );
  NAND4_X1 u1_u0_u1_U85 (.ZN( u1_out0_28 ) , .A4( u1_u0_u1_n124 ) , .A3( u1_u0_u1_n125 ) , .A2( u1_u0_u1_n126 ) , .A1( u1_u0_u1_n127 ) );
  OAI21_X1 u1_u0_u1_U86 (.ZN( u1_u0_u1_n127 ) , .B2( u1_u0_u1_n139 ) , .B1( u1_u0_u1_n175 ) , .A( u1_u0_u1_n183 ) );
  OAI21_X1 u1_u0_u1_U87 (.ZN( u1_u0_u1_n126 ) , .B2( u1_u0_u1_n140 ) , .A( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n178 ) );
  NAND4_X1 u1_u0_u1_U88 (.ZN( u1_out0_18 ) , .A4( u1_u0_u1_n165 ) , .A3( u1_u0_u1_n166 ) , .A1( u1_u0_u1_n167 ) , .A2( u1_u0_u1_n186 ) );
  AOI22_X1 u1_u0_u1_U89 (.B2( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n147 ) , .A2( u1_u0_u1_n148 ) , .ZN( u1_u0_u1_n166 ) , .A1( u1_u0_u1_n172 ) );
  OAI21_X1 u1_u0_u1_U9 (.ZN( u1_u0_u1_n101 ) , .B1( u1_u0_u1_n141 ) , .A( u1_u0_u1_n146 ) , .B2( u1_u0_u1_n183 ) );
  INV_X1 u1_u0_u1_U90 (.A( u1_u0_u1_n145 ) , .ZN( u1_u0_u1_n186 ) );
  NAND4_X1 u1_u0_u1_U91 (.ZN( u1_out0_2 ) , .A4( u1_u0_u1_n142 ) , .A3( u1_u0_u1_n143 ) , .A2( u1_u0_u1_n144 ) , .A1( u1_u0_u1_n179 ) );
  OAI21_X1 u1_u0_u1_U92 (.B2( u1_u0_u1_n132 ) , .ZN( u1_u0_u1_n144 ) , .A( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n180 ) );
  INV_X1 u1_u0_u1_U93 (.A( u1_u0_u1_n130 ) , .ZN( u1_u0_u1_n179 ) );
  OR4_X1 u1_u0_u1_U94 (.ZN( u1_out0_13 ) , .A4( u1_u0_u1_n108 ) , .A3( u1_u0_u1_n109 ) , .A2( u1_u0_u1_n110 ) , .A1( u1_u0_u1_n111 ) );
  AOI21_X1 u1_u0_u1_U95 (.ZN( u1_u0_u1_n111 ) , .A( u1_u0_u1_n128 ) , .B2( u1_u0_u1_n131 ) , .B1( u1_u0_u1_n135 ) );
  AOI21_X1 u1_u0_u1_U96 (.ZN( u1_u0_u1_n110 ) , .A( u1_u0_u1_n116 ) , .B1( u1_u0_u1_n152 ) , .B2( u1_u0_u1_n160 ) );
  NAND3_X1 u1_u0_u1_U97 (.A3( u1_u0_u1_n149 ) , .A2( u1_u0_u1_n150 ) , .A1( u1_u0_u1_n151 ) , .ZN( u1_u0_u1_n164 ) );
  NAND3_X1 u1_u0_u1_U98 (.A3( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n135 ) , .ZN( u1_u0_u1_n136 ) , .A1( u1_u0_u1_n151 ) );
  NAND3_X1 u1_u0_u1_U99 (.A1( u1_u0_u1_n133 ) , .ZN( u1_u0_u1_n137 ) , .A2( u1_u0_u1_n154 ) , .A3( u1_u0_u1_n181 ) );
  OAI22_X1 u1_u0_u2_U10 (.B1( u1_u0_u2_n151 ) , .A2( u1_u0_u2_n152 ) , .A1( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n160 ) , .B2( u1_u0_u2_n168 ) );
  NAND3_X1 u1_u0_u2_U100 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n104 ) , .A3( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n98 ) );
  NOR3_X1 u1_u0_u2_U11 (.A1( u1_u0_u2_n150 ) , .ZN( u1_u0_u2_n151 ) , .A3( u1_u0_u2_n175 ) , .A2( u1_u0_u2_n188 ) );
  AOI21_X1 u1_u0_u2_U12 (.B2( u1_u0_u2_n123 ) , .ZN( u1_u0_u2_n125 ) , .A( u1_u0_u2_n171 ) , .B1( u1_u0_u2_n184 ) );
  INV_X1 u1_u0_u2_U13 (.A( u1_u0_u2_n150 ) , .ZN( u1_u0_u2_n184 ) );
  AOI21_X1 u1_u0_u2_U14 (.ZN( u1_u0_u2_n144 ) , .B2( u1_u0_u2_n155 ) , .A( u1_u0_u2_n172 ) , .B1( u1_u0_u2_n185 ) );
  AOI21_X1 u1_u0_u2_U15 (.B2( u1_u0_u2_n143 ) , .ZN( u1_u0_u2_n145 ) , .B1( u1_u0_u2_n152 ) , .A( u1_u0_u2_n171 ) );
  INV_X1 u1_u0_u2_U16 (.A( u1_u0_u2_n156 ) , .ZN( u1_u0_u2_n171 ) );
  INV_X1 u1_u0_u2_U17 (.A( u1_u0_u2_n120 ) , .ZN( u1_u0_u2_n188 ) );
  NAND2_X1 u1_u0_u2_U18 (.A2( u1_u0_u2_n122 ) , .ZN( u1_u0_u2_n150 ) , .A1( u1_u0_u2_n152 ) );
  INV_X1 u1_u0_u2_U19 (.A( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n170 ) );
  INV_X1 u1_u0_u2_U20 (.A( u1_u0_u2_n137 ) , .ZN( u1_u0_u2_n173 ) );
  NAND2_X1 u1_u0_u2_U21 (.A1( u1_u0_u2_n132 ) , .A2( u1_u0_u2_n139 ) , .ZN( u1_u0_u2_n157 ) );
  INV_X1 u1_u0_u2_U22 (.A( u1_u0_u2_n113 ) , .ZN( u1_u0_u2_n178 ) );
  INV_X1 u1_u0_u2_U23 (.A( u1_u0_u2_n139 ) , .ZN( u1_u0_u2_n175 ) );
  INV_X1 u1_u0_u2_U24 (.A( u1_u0_u2_n155 ) , .ZN( u1_u0_u2_n181 ) );
  INV_X1 u1_u0_u2_U25 (.A( u1_u0_u2_n119 ) , .ZN( u1_u0_u2_n177 ) );
  INV_X1 u1_u0_u2_U26 (.A( u1_u0_u2_n116 ) , .ZN( u1_u0_u2_n180 ) );
  INV_X1 u1_u0_u2_U27 (.A( u1_u0_u2_n131 ) , .ZN( u1_u0_u2_n179 ) );
  INV_X1 u1_u0_u2_U28 (.A( u1_u0_u2_n154 ) , .ZN( u1_u0_u2_n176 ) );
  NAND2_X1 u1_u0_u2_U29 (.A2( u1_u0_u2_n116 ) , .A1( u1_u0_u2_n117 ) , .ZN( u1_u0_u2_n118 ) );
  NOR2_X1 u1_u0_u2_U3 (.ZN( u1_u0_u2_n121 ) , .A2( u1_u0_u2_n177 ) , .A1( u1_u0_u2_n180 ) );
  INV_X1 u1_u0_u2_U30 (.A( u1_u0_u2_n132 ) , .ZN( u1_u0_u2_n182 ) );
  INV_X1 u1_u0_u2_U31 (.A( u1_u0_u2_n158 ) , .ZN( u1_u0_u2_n183 ) );
  OAI21_X1 u1_u0_u2_U32 (.A( u1_u0_u2_n156 ) , .B1( u1_u0_u2_n157 ) , .ZN( u1_u0_u2_n158 ) , .B2( u1_u0_u2_n179 ) );
  NOR2_X1 u1_u0_u2_U33 (.ZN( u1_u0_u2_n156 ) , .A1( u1_u0_u2_n166 ) , .A2( u1_u0_u2_n169 ) );
  NOR2_X1 u1_u0_u2_U34 (.A2( u1_u0_u2_n114 ) , .ZN( u1_u0_u2_n137 ) , .A1( u1_u0_u2_n140 ) );
  NOR2_X1 u1_u0_u2_U35 (.A2( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n153 ) , .A1( u1_u0_u2_n156 ) );
  AOI211_X1 u1_u0_u2_U36 (.ZN( u1_u0_u2_n130 ) , .C1( u1_u0_u2_n138 ) , .C2( u1_u0_u2_n179 ) , .B( u1_u0_u2_n96 ) , .A( u1_u0_u2_n97 ) );
  OAI22_X1 u1_u0_u2_U37 (.B1( u1_u0_u2_n133 ) , .A2( u1_u0_u2_n137 ) , .A1( u1_u0_u2_n152 ) , .B2( u1_u0_u2_n168 ) , .ZN( u1_u0_u2_n97 ) );
  OAI221_X1 u1_u0_u2_U38 (.B1( u1_u0_u2_n113 ) , .C1( u1_u0_u2_n132 ) , .A( u1_u0_u2_n149 ) , .B2( u1_u0_u2_n171 ) , .C2( u1_u0_u2_n172 ) , .ZN( u1_u0_u2_n96 ) );
  OAI221_X1 u1_u0_u2_U39 (.A( u1_u0_u2_n115 ) , .C2( u1_u0_u2_n123 ) , .B2( u1_u0_u2_n143 ) , .B1( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n163 ) , .C1( u1_u0_u2_n168 ) );
  INV_X1 u1_u0_u2_U4 (.A( u1_u0_u2_n134 ) , .ZN( u1_u0_u2_n185 ) );
  OAI21_X1 u1_u0_u2_U40 (.A( u1_u0_u2_n114 ) , .ZN( u1_u0_u2_n115 ) , .B1( u1_u0_u2_n176 ) , .B2( u1_u0_u2_n178 ) );
  OAI221_X1 u1_u0_u2_U41 (.A( u1_u0_u2_n135 ) , .B2( u1_u0_u2_n136 ) , .B1( u1_u0_u2_n137 ) , .ZN( u1_u0_u2_n162 ) , .C2( u1_u0_u2_n167 ) , .C1( u1_u0_u2_n185 ) );
  AND3_X1 u1_u0_u2_U42 (.A3( u1_u0_u2_n131 ) , .A2( u1_u0_u2_n132 ) , .A1( u1_u0_u2_n133 ) , .ZN( u1_u0_u2_n136 ) );
  AOI22_X1 u1_u0_u2_U43 (.ZN( u1_u0_u2_n135 ) , .B1( u1_u0_u2_n140 ) , .A1( u1_u0_u2_n156 ) , .B2( u1_u0_u2_n180 ) , .A2( u1_u0_u2_n188 ) );
  AOI21_X1 u1_u0_u2_U44 (.ZN( u1_u0_u2_n149 ) , .B1( u1_u0_u2_n173 ) , .B2( u1_u0_u2_n188 ) , .A( u1_u0_u2_n95 ) );
  AND3_X1 u1_u0_u2_U45 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n104 ) , .A3( u1_u0_u2_n156 ) , .ZN( u1_u0_u2_n95 ) );
  OAI21_X1 u1_u0_u2_U46 (.A( u1_u0_u2_n101 ) , .B2( u1_u0_u2_n121 ) , .B1( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n164 ) );
  NAND2_X1 u1_u0_u2_U47 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n107 ) , .ZN( u1_u0_u2_n155 ) );
  NAND2_X1 u1_u0_u2_U48 (.A2( u1_u0_u2_n105 ) , .A1( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n143 ) );
  NAND2_X1 u1_u0_u2_U49 (.A1( u1_u0_u2_n104 ) , .A2( u1_u0_u2_n106 ) , .ZN( u1_u0_u2_n152 ) );
  NOR4_X1 u1_u0_u2_U5 (.A4( u1_u0_u2_n124 ) , .A3( u1_u0_u2_n125 ) , .A2( u1_u0_u2_n126 ) , .A1( u1_u0_u2_n127 ) , .ZN( u1_u0_u2_n128 ) );
  NAND2_X1 u1_u0_u2_U50 (.A1( u1_u0_u2_n100 ) , .A2( u1_u0_u2_n105 ) , .ZN( u1_u0_u2_n132 ) );
  INV_X1 u1_u0_u2_U51 (.A( u1_u0_u2_n140 ) , .ZN( u1_u0_u2_n168 ) );
  INV_X1 u1_u0_u2_U52 (.A( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n167 ) );
  OAI21_X1 u1_u0_u2_U53 (.A( u1_u0_u2_n141 ) , .B2( u1_u0_u2_n142 ) , .ZN( u1_u0_u2_n146 ) , .B1( u1_u0_u2_n153 ) );
  OAI21_X1 u1_u0_u2_U54 (.A( u1_u0_u2_n140 ) , .ZN( u1_u0_u2_n141 ) , .B1( u1_u0_u2_n176 ) , .B2( u1_u0_u2_n177 ) );
  NOR3_X1 u1_u0_u2_U55 (.ZN( u1_u0_u2_n142 ) , .A3( u1_u0_u2_n175 ) , .A2( u1_u0_u2_n178 ) , .A1( u1_u0_u2_n181 ) );
  NAND2_X1 u1_u0_u2_U56 (.A1( u1_u0_u2_n102 ) , .A2( u1_u0_u2_n106 ) , .ZN( u1_u0_u2_n113 ) );
  NAND2_X1 u1_u0_u2_U57 (.A1( u1_u0_u2_n106 ) , .A2( u1_u0_u2_n107 ) , .ZN( u1_u0_u2_n131 ) );
  NAND2_X1 u1_u0_u2_U58 (.A1( u1_u0_u2_n103 ) , .A2( u1_u0_u2_n107 ) , .ZN( u1_u0_u2_n139 ) );
  NAND2_X1 u1_u0_u2_U59 (.A1( u1_u0_u2_n103 ) , .A2( u1_u0_u2_n105 ) , .ZN( u1_u0_u2_n133 ) );
  AOI21_X1 u1_u0_u2_U6 (.B2( u1_u0_u2_n119 ) , .ZN( u1_u0_u2_n127 ) , .A( u1_u0_u2_n137 ) , .B1( u1_u0_u2_n155 ) );
  NAND2_X1 u1_u0_u2_U60 (.A1( u1_u0_u2_n102 ) , .A2( u1_u0_u2_n103 ) , .ZN( u1_u0_u2_n154 ) );
  NAND2_X1 u1_u0_u2_U61 (.A2( u1_u0_u2_n103 ) , .A1( u1_u0_u2_n104 ) , .ZN( u1_u0_u2_n119 ) );
  NAND2_X1 u1_u0_u2_U62 (.A2( u1_u0_u2_n107 ) , .A1( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n123 ) );
  NAND2_X1 u1_u0_u2_U63 (.A1( u1_u0_u2_n104 ) , .A2( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n122 ) );
  INV_X1 u1_u0_u2_U64 (.A( u1_u0_u2_n114 ) , .ZN( u1_u0_u2_n172 ) );
  NAND2_X1 u1_u0_u2_U65 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n102 ) , .ZN( u1_u0_u2_n116 ) );
  NAND2_X1 u1_u0_u2_U66 (.A1( u1_u0_u2_n102 ) , .A2( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n120 ) );
  NAND2_X1 u1_u0_u2_U67 (.A2( u1_u0_u2_n105 ) , .A1( u1_u0_u2_n106 ) , .ZN( u1_u0_u2_n117 ) );
  INV_X1 u1_u0_u2_U68 (.ZN( u1_u0_u2_n187 ) , .A( u1_u0_u2_n99 ) );
  OAI21_X1 u1_u0_u2_U69 (.B1( u1_u0_u2_n137 ) , .B2( u1_u0_u2_n143 ) , .A( u1_u0_u2_n98 ) , .ZN( u1_u0_u2_n99 ) );
  AOI21_X1 u1_u0_u2_U7 (.ZN( u1_u0_u2_n124 ) , .B1( u1_u0_u2_n131 ) , .B2( u1_u0_u2_n143 ) , .A( u1_u0_u2_n172 ) );
  NOR2_X1 u1_u0_u2_U70 (.A2( u1_u0_X_16 ) , .ZN( u1_u0_u2_n140 ) , .A1( u1_u0_u2_n166 ) );
  NOR2_X1 u1_u0_u2_U71 (.A2( u1_u0_X_13 ) , .A1( u1_u0_X_14 ) , .ZN( u1_u0_u2_n100 ) );
  NOR2_X1 u1_u0_u2_U72 (.A2( u1_u0_X_16 ) , .A1( u1_u0_X_17 ) , .ZN( u1_u0_u2_n138 ) );
  NOR2_X1 u1_u0_u2_U73 (.A2( u1_u0_X_15 ) , .A1( u1_u0_X_18 ) , .ZN( u1_u0_u2_n104 ) );
  NOR2_X1 u1_u0_u2_U74 (.A2( u1_u0_X_14 ) , .ZN( u1_u0_u2_n103 ) , .A1( u1_u0_u2_n174 ) );
  NOR2_X1 u1_u0_u2_U75 (.A2( u1_u0_X_15 ) , .ZN( u1_u0_u2_n102 ) , .A1( u1_u0_u2_n165 ) );
  NOR2_X1 u1_u0_u2_U76 (.A2( u1_u0_X_17 ) , .ZN( u1_u0_u2_n114 ) , .A1( u1_u0_u2_n169 ) );
  AND2_X1 u1_u0_u2_U77 (.A1( u1_u0_X_15 ) , .ZN( u1_u0_u2_n105 ) , .A2( u1_u0_u2_n165 ) );
  AND2_X1 u1_u0_u2_U78 (.A2( u1_u0_X_15 ) , .A1( u1_u0_X_18 ) , .ZN( u1_u0_u2_n107 ) );
  AND2_X1 u1_u0_u2_U79 (.A1( u1_u0_X_14 ) , .ZN( u1_u0_u2_n106 ) , .A2( u1_u0_u2_n174 ) );
  AOI21_X1 u1_u0_u2_U8 (.B2( u1_u0_u2_n120 ) , .B1( u1_u0_u2_n121 ) , .ZN( u1_u0_u2_n126 ) , .A( u1_u0_u2_n167 ) );
  AND2_X1 u1_u0_u2_U80 (.A1( u1_u0_X_13 ) , .A2( u1_u0_X_14 ) , .ZN( u1_u0_u2_n108 ) );
  INV_X1 u1_u0_u2_U81 (.A( u1_u0_X_16 ) , .ZN( u1_u0_u2_n169 ) );
  INV_X1 u1_u0_u2_U82 (.A( u1_u0_X_17 ) , .ZN( u1_u0_u2_n166 ) );
  INV_X1 u1_u0_u2_U83 (.A( u1_u0_X_13 ) , .ZN( u1_u0_u2_n174 ) );
  INV_X1 u1_u0_u2_U84 (.A( u1_u0_X_18 ) , .ZN( u1_u0_u2_n165 ) );
  NAND4_X1 u1_u0_u2_U85 (.ZN( u1_out0_30 ) , .A4( u1_u0_u2_n147 ) , .A3( u1_u0_u2_n148 ) , .A2( u1_u0_u2_n149 ) , .A1( u1_u0_u2_n187 ) );
  NOR3_X1 u1_u0_u2_U86 (.A3( u1_u0_u2_n144 ) , .A2( u1_u0_u2_n145 ) , .A1( u1_u0_u2_n146 ) , .ZN( u1_u0_u2_n147 ) );
  AOI21_X1 u1_u0_u2_U87 (.B2( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n148 ) , .A( u1_u0_u2_n162 ) , .B1( u1_u0_u2_n182 ) );
  NAND4_X1 u1_u0_u2_U88 (.ZN( u1_out0_24 ) , .A4( u1_u0_u2_n111 ) , .A3( u1_u0_u2_n112 ) , .A1( u1_u0_u2_n130 ) , .A2( u1_u0_u2_n187 ) );
  AOI221_X1 u1_u0_u2_U89 (.A( u1_u0_u2_n109 ) , .B1( u1_u0_u2_n110 ) , .ZN( u1_u0_u2_n111 ) , .C1( u1_u0_u2_n134 ) , .C2( u1_u0_u2_n170 ) , .B2( u1_u0_u2_n173 ) );
  OAI22_X1 u1_u0_u2_U9 (.ZN( u1_u0_u2_n109 ) , .A2( u1_u0_u2_n113 ) , .B2( u1_u0_u2_n133 ) , .B1( u1_u0_u2_n167 ) , .A1( u1_u0_u2_n168 ) );
  AOI21_X1 u1_u0_u2_U90 (.ZN( u1_u0_u2_n112 ) , .B2( u1_u0_u2_n156 ) , .A( u1_u0_u2_n164 ) , .B1( u1_u0_u2_n181 ) );
  NAND4_X1 u1_u0_u2_U91 (.ZN( u1_out0_16 ) , .A4( u1_u0_u2_n128 ) , .A3( u1_u0_u2_n129 ) , .A1( u1_u0_u2_n130 ) , .A2( u1_u0_u2_n186 ) );
  AOI22_X1 u1_u0_u2_U92 (.A2( u1_u0_u2_n118 ) , .ZN( u1_u0_u2_n129 ) , .A1( u1_u0_u2_n140 ) , .B1( u1_u0_u2_n157 ) , .B2( u1_u0_u2_n170 ) );
  INV_X1 u1_u0_u2_U93 (.A( u1_u0_u2_n163 ) , .ZN( u1_u0_u2_n186 ) );
  OR4_X1 u1_u0_u2_U94 (.ZN( u1_out0_6 ) , .A4( u1_u0_u2_n161 ) , .A3( u1_u0_u2_n162 ) , .A2( u1_u0_u2_n163 ) , .A1( u1_u0_u2_n164 ) );
  OR3_X1 u1_u0_u2_U95 (.A2( u1_u0_u2_n159 ) , .A1( u1_u0_u2_n160 ) , .ZN( u1_u0_u2_n161 ) , .A3( u1_u0_u2_n183 ) );
  AOI21_X1 u1_u0_u2_U96 (.B2( u1_u0_u2_n154 ) , .B1( u1_u0_u2_n155 ) , .ZN( u1_u0_u2_n159 ) , .A( u1_u0_u2_n167 ) );
  NAND3_X1 u1_u0_u2_U97 (.A2( u1_u0_u2_n117 ) , .A1( u1_u0_u2_n122 ) , .A3( u1_u0_u2_n123 ) , .ZN( u1_u0_u2_n134 ) );
  NAND3_X1 u1_u0_u2_U98 (.ZN( u1_u0_u2_n110 ) , .A2( u1_u0_u2_n131 ) , .A3( u1_u0_u2_n139 ) , .A1( u1_u0_u2_n154 ) );
  NAND3_X1 u1_u0_u2_U99 (.A2( u1_u0_u2_n100 ) , .ZN( u1_u0_u2_n101 ) , .A1( u1_u0_u2_n104 ) , .A3( u1_u0_u2_n114 ) );
  OAI22_X1 u1_u0_u3_U10 (.B1( u1_u0_u3_n113 ) , .A2( u1_u0_u3_n135 ) , .A1( u1_u0_u3_n150 ) , .B2( u1_u0_u3_n164 ) , .ZN( u1_u0_u3_n98 ) );
  OAI211_X1 u1_u0_u3_U11 (.B( u1_u0_u3_n106 ) , .ZN( u1_u0_u3_n119 ) , .C2( u1_u0_u3_n128 ) , .C1( u1_u0_u3_n167 ) , .A( u1_u0_u3_n181 ) );
  AOI221_X1 u1_u0_u3_U12 (.C1( u1_u0_u3_n105 ) , .ZN( u1_u0_u3_n106 ) , .A( u1_u0_u3_n131 ) , .B2( u1_u0_u3_n132 ) , .C2( u1_u0_u3_n133 ) , .B1( u1_u0_u3_n169 ) );
  INV_X1 u1_u0_u3_U13 (.ZN( u1_u0_u3_n181 ) , .A( u1_u0_u3_n98 ) );
  NAND2_X1 u1_u0_u3_U14 (.ZN( u1_u0_u3_n105 ) , .A2( u1_u0_u3_n130 ) , .A1( u1_u0_u3_n155 ) );
  AOI22_X1 u1_u0_u3_U15 (.B1( u1_u0_u3_n115 ) , .A2( u1_u0_u3_n116 ) , .ZN( u1_u0_u3_n123 ) , .B2( u1_u0_u3_n133 ) , .A1( u1_u0_u3_n169 ) );
  NAND2_X1 u1_u0_u3_U16 (.ZN( u1_u0_u3_n116 ) , .A2( u1_u0_u3_n151 ) , .A1( u1_u0_u3_n182 ) );
  NOR2_X1 u1_u0_u3_U17 (.ZN( u1_u0_u3_n126 ) , .A2( u1_u0_u3_n150 ) , .A1( u1_u0_u3_n164 ) );
  AOI21_X1 u1_u0_u3_U18 (.ZN( u1_u0_u3_n112 ) , .B2( u1_u0_u3_n146 ) , .B1( u1_u0_u3_n155 ) , .A( u1_u0_u3_n167 ) );
  NAND2_X1 u1_u0_u3_U19 (.A1( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n142 ) , .A2( u1_u0_u3_n164 ) );
  NAND2_X1 u1_u0_u3_U20 (.ZN( u1_u0_u3_n132 ) , .A2( u1_u0_u3_n152 ) , .A1( u1_u0_u3_n156 ) );
  INV_X1 u1_u0_u3_U21 (.A( u1_u0_u3_n133 ) , .ZN( u1_u0_u3_n165 ) );
  AND2_X1 u1_u0_u3_U22 (.A2( u1_u0_u3_n113 ) , .A1( u1_u0_u3_n114 ) , .ZN( u1_u0_u3_n151 ) );
  INV_X1 u1_u0_u3_U23 (.A( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n170 ) );
  NAND2_X1 u1_u0_u3_U24 (.A1( u1_u0_u3_n107 ) , .A2( u1_u0_u3_n108 ) , .ZN( u1_u0_u3_n140 ) );
  NAND2_X1 u1_u0_u3_U25 (.ZN( u1_u0_u3_n117 ) , .A1( u1_u0_u3_n124 ) , .A2( u1_u0_u3_n148 ) );
  NAND2_X1 u1_u0_u3_U26 (.ZN( u1_u0_u3_n143 ) , .A1( u1_u0_u3_n165 ) , .A2( u1_u0_u3_n167 ) );
  INV_X1 u1_u0_u3_U27 (.A( u1_u0_u3_n130 ) , .ZN( u1_u0_u3_n177 ) );
  INV_X1 u1_u0_u3_U28 (.A( u1_u0_u3_n128 ) , .ZN( u1_u0_u3_n176 ) );
  INV_X1 u1_u0_u3_U29 (.A( u1_u0_u3_n155 ) , .ZN( u1_u0_u3_n174 ) );
  INV_X1 u1_u0_u3_U3 (.A( u1_u0_u3_n140 ) , .ZN( u1_u0_u3_n182 ) );
  INV_X1 u1_u0_u3_U30 (.A( u1_u0_u3_n139 ) , .ZN( u1_u0_u3_n185 ) );
  NOR2_X1 u1_u0_u3_U31 (.ZN( u1_u0_u3_n135 ) , .A2( u1_u0_u3_n141 ) , .A1( u1_u0_u3_n169 ) );
  OAI222_X1 u1_u0_u3_U32 (.C2( u1_u0_u3_n107 ) , .A2( u1_u0_u3_n108 ) , .B1( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n138 ) , .B2( u1_u0_u3_n146 ) , .C1( u1_u0_u3_n154 ) , .A1( u1_u0_u3_n164 ) );
  NOR4_X1 u1_u0_u3_U33 (.A4( u1_u0_u3_n157 ) , .A3( u1_u0_u3_n158 ) , .A2( u1_u0_u3_n159 ) , .A1( u1_u0_u3_n160 ) , .ZN( u1_u0_u3_n161 ) );
  AOI21_X1 u1_u0_u3_U34 (.B2( u1_u0_u3_n152 ) , .B1( u1_u0_u3_n153 ) , .ZN( u1_u0_u3_n158 ) , .A( u1_u0_u3_n164 ) );
  AOI21_X1 u1_u0_u3_U35 (.A( u1_u0_u3_n154 ) , .B2( u1_u0_u3_n155 ) , .B1( u1_u0_u3_n156 ) , .ZN( u1_u0_u3_n157 ) );
  AOI21_X1 u1_u0_u3_U36 (.A( u1_u0_u3_n149 ) , .B2( u1_u0_u3_n150 ) , .B1( u1_u0_u3_n151 ) , .ZN( u1_u0_u3_n159 ) );
  OAI211_X1 u1_u0_u3_U37 (.B( u1_u0_u3_n127 ) , .ZN( u1_u0_u3_n139 ) , .C1( u1_u0_u3_n150 ) , .C2( u1_u0_u3_n154 ) , .A( u1_u0_u3_n184 ) );
  INV_X1 u1_u0_u3_U38 (.A( u1_u0_u3_n125 ) , .ZN( u1_u0_u3_n184 ) );
  AOI221_X1 u1_u0_u3_U39 (.A( u1_u0_u3_n126 ) , .ZN( u1_u0_u3_n127 ) , .C2( u1_u0_u3_n132 ) , .C1( u1_u0_u3_n169 ) , .B2( u1_u0_u3_n170 ) , .B1( u1_u0_u3_n174 ) );
  INV_X1 u1_u0_u3_U4 (.A( u1_u0_u3_n129 ) , .ZN( u1_u0_u3_n183 ) );
  OAI22_X1 u1_u0_u3_U40 (.A1( u1_u0_u3_n124 ) , .ZN( u1_u0_u3_n125 ) , .B2( u1_u0_u3_n145 ) , .A2( u1_u0_u3_n165 ) , .B1( u1_u0_u3_n167 ) );
  AOI211_X1 u1_u0_u3_U41 (.ZN( u1_u0_u3_n109 ) , .A( u1_u0_u3_n119 ) , .C2( u1_u0_u3_n129 ) , .B( u1_u0_u3_n138 ) , .C1( u1_u0_u3_n141 ) );
  AOI211_X1 u1_u0_u3_U42 (.B( u1_u0_u3_n119 ) , .A( u1_u0_u3_n120 ) , .C2( u1_u0_u3_n121 ) , .ZN( u1_u0_u3_n122 ) , .C1( u1_u0_u3_n179 ) );
  INV_X1 u1_u0_u3_U43 (.A( u1_u0_u3_n156 ) , .ZN( u1_u0_u3_n179 ) );
  OAI22_X1 u1_u0_u3_U44 (.B1( u1_u0_u3_n118 ) , .ZN( u1_u0_u3_n120 ) , .A1( u1_u0_u3_n135 ) , .B2( u1_u0_u3_n154 ) , .A2( u1_u0_u3_n178 ) );
  AND3_X1 u1_u0_u3_U45 (.ZN( u1_u0_u3_n118 ) , .A2( u1_u0_u3_n124 ) , .A1( u1_u0_u3_n144 ) , .A3( u1_u0_u3_n152 ) );
  INV_X1 u1_u0_u3_U46 (.A( u1_u0_u3_n121 ) , .ZN( u1_u0_u3_n164 ) );
  NAND2_X1 u1_u0_u3_U47 (.ZN( u1_u0_u3_n133 ) , .A1( u1_u0_u3_n154 ) , .A2( u1_u0_u3_n164 ) );
  NOR2_X1 u1_u0_u3_U48 (.A1( u1_u0_u3_n113 ) , .ZN( u1_u0_u3_n131 ) , .A2( u1_u0_u3_n154 ) );
  NAND2_X1 u1_u0_u3_U49 (.A1( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n150 ) , .A2( u1_u0_u3_n99 ) );
  INV_X1 u1_u0_u3_U5 (.A( u1_u0_u3_n117 ) , .ZN( u1_u0_u3_n178 ) );
  NAND2_X1 u1_u0_u3_U50 (.A2( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n155 ) , .A1( u1_u0_u3_n97 ) );
  INV_X1 u1_u0_u3_U51 (.A( u1_u0_u3_n141 ) , .ZN( u1_u0_u3_n167 ) );
  AOI21_X1 u1_u0_u3_U52 (.B2( u1_u0_u3_n114 ) , .B1( u1_u0_u3_n146 ) , .A( u1_u0_u3_n154 ) , .ZN( u1_u0_u3_n94 ) );
  AOI21_X1 u1_u0_u3_U53 (.ZN( u1_u0_u3_n110 ) , .B2( u1_u0_u3_n142 ) , .B1( u1_u0_u3_n186 ) , .A( u1_u0_u3_n95 ) );
  INV_X1 u1_u0_u3_U54 (.A( u1_u0_u3_n145 ) , .ZN( u1_u0_u3_n186 ) );
  AOI21_X1 u1_u0_u3_U55 (.B1( u1_u0_u3_n124 ) , .A( u1_u0_u3_n149 ) , .B2( u1_u0_u3_n155 ) , .ZN( u1_u0_u3_n95 ) );
  INV_X1 u1_u0_u3_U56 (.A( u1_u0_u3_n149 ) , .ZN( u1_u0_u3_n169 ) );
  NAND2_X1 u1_u0_u3_U57 (.ZN( u1_u0_u3_n124 ) , .A1( u1_u0_u3_n96 ) , .A2( u1_u0_u3_n97 ) );
  NAND2_X1 u1_u0_u3_U58 (.A2( u1_u0_u3_n100 ) , .ZN( u1_u0_u3_n146 ) , .A1( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U59 (.A1( u1_u0_u3_n101 ) , .ZN( u1_u0_u3_n145 ) , .A2( u1_u0_u3_n99 ) );
  AOI221_X1 u1_u0_u3_U6 (.A( u1_u0_u3_n131 ) , .C2( u1_u0_u3_n132 ) , .C1( u1_u0_u3_n133 ) , .ZN( u1_u0_u3_n134 ) , .B1( u1_u0_u3_n143 ) , .B2( u1_u0_u3_n177 ) );
  NAND2_X1 u1_u0_u3_U60 (.A1( u1_u0_u3_n100 ) , .ZN( u1_u0_u3_n156 ) , .A2( u1_u0_u3_n99 ) );
  NAND2_X1 u1_u0_u3_U61 (.A2( u1_u0_u3_n101 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n148 ) );
  NAND2_X1 u1_u0_u3_U62 (.A1( u1_u0_u3_n100 ) , .A2( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n128 ) );
  NAND2_X1 u1_u0_u3_U63 (.A2( u1_u0_u3_n101 ) , .A1( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n152 ) );
  NAND2_X1 u1_u0_u3_U64 (.A2( u1_u0_u3_n101 ) , .ZN( u1_u0_u3_n114 ) , .A1( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U65 (.ZN( u1_u0_u3_n107 ) , .A1( u1_u0_u3_n97 ) , .A2( u1_u0_u3_n99 ) );
  NAND2_X1 u1_u0_u3_U66 (.A2( u1_u0_u3_n100 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n113 ) );
  NAND2_X1 u1_u0_u3_U67 (.A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n153 ) , .A2( u1_u0_u3_n97 ) );
  NAND2_X1 u1_u0_u3_U68 (.A2( u1_u0_u3_n103 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n130 ) );
  NAND2_X1 u1_u0_u3_U69 (.A2( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n144 ) , .A1( u1_u0_u3_n96 ) );
  OAI22_X1 u1_u0_u3_U7 (.B2( u1_u0_u3_n147 ) , .A2( u1_u0_u3_n148 ) , .ZN( u1_u0_u3_n160 ) , .B1( u1_u0_u3_n165 ) , .A1( u1_u0_u3_n168 ) );
  NAND2_X1 u1_u0_u3_U70 (.A1( u1_u0_u3_n102 ) , .A2( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n108 ) );
  NOR2_X1 u1_u0_u3_U71 (.A2( u1_u0_X_19 ) , .A1( u1_u0_X_20 ) , .ZN( u1_u0_u3_n99 ) );
  NOR2_X1 u1_u0_u3_U72 (.A2( u1_u0_X_21 ) , .A1( u1_u0_X_24 ) , .ZN( u1_u0_u3_n103 ) );
  NOR2_X1 u1_u0_u3_U73 (.A2( u1_u0_X_24 ) , .A1( u1_u0_u3_n171 ) , .ZN( u1_u0_u3_n97 ) );
  NOR2_X1 u1_u0_u3_U74 (.A2( u1_u0_X_23 ) , .ZN( u1_u0_u3_n141 ) , .A1( u1_u0_u3_n166 ) );
  NOR2_X1 u1_u0_u3_U75 (.A2( u1_u0_X_19 ) , .A1( u1_u0_u3_n172 ) , .ZN( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U76 (.A1( u1_u0_X_22 ) , .A2( u1_u0_X_23 ) , .ZN( u1_u0_u3_n154 ) );
  NAND2_X1 u1_u0_u3_U77 (.A1( u1_u0_X_23 ) , .ZN( u1_u0_u3_n149 ) , .A2( u1_u0_u3_n166 ) );
  NOR2_X1 u1_u0_u3_U78 (.A2( u1_u0_X_22 ) , .A1( u1_u0_X_23 ) , .ZN( u1_u0_u3_n121 ) );
  AND2_X1 u1_u0_u3_U79 (.A1( u1_u0_X_24 ) , .ZN( u1_u0_u3_n101 ) , .A2( u1_u0_u3_n171 ) );
  AND3_X1 u1_u0_u3_U8 (.A3( u1_u0_u3_n144 ) , .A2( u1_u0_u3_n145 ) , .A1( u1_u0_u3_n146 ) , .ZN( u1_u0_u3_n147 ) );
  AND2_X1 u1_u0_u3_U80 (.A1( u1_u0_X_19 ) , .ZN( u1_u0_u3_n102 ) , .A2( u1_u0_u3_n172 ) );
  AND2_X1 u1_u0_u3_U81 (.A1( u1_u0_X_21 ) , .A2( u1_u0_X_24 ) , .ZN( u1_u0_u3_n100 ) );
  AND2_X1 u1_u0_u3_U82 (.A2( u1_u0_X_19 ) , .A1( u1_u0_X_20 ) , .ZN( u1_u0_u3_n104 ) );
  INV_X1 u1_u0_u3_U83 (.A( u1_u0_X_22 ) , .ZN( u1_u0_u3_n166 ) );
  INV_X1 u1_u0_u3_U84 (.A( u1_u0_X_21 ) , .ZN( u1_u0_u3_n171 ) );
  INV_X1 u1_u0_u3_U85 (.A( u1_u0_X_20 ) , .ZN( u1_u0_u3_n172 ) );
  NAND4_X1 u1_u0_u3_U86 (.ZN( u1_out0_26 ) , .A4( u1_u0_u3_n109 ) , .A3( u1_u0_u3_n110 ) , .A2( u1_u0_u3_n111 ) , .A1( u1_u0_u3_n173 ) );
  INV_X1 u1_u0_u3_U87 (.ZN( u1_u0_u3_n173 ) , .A( u1_u0_u3_n94 ) );
  OAI21_X1 u1_u0_u3_U88 (.ZN( u1_u0_u3_n111 ) , .B2( u1_u0_u3_n117 ) , .A( u1_u0_u3_n133 ) , .B1( u1_u0_u3_n176 ) );
  NAND4_X1 u1_u0_u3_U89 (.ZN( u1_out0_20 ) , .A4( u1_u0_u3_n122 ) , .A3( u1_u0_u3_n123 ) , .A1( u1_u0_u3_n175 ) , .A2( u1_u0_u3_n180 ) );
  INV_X1 u1_u0_u3_U9 (.A( u1_u0_u3_n143 ) , .ZN( u1_u0_u3_n168 ) );
  INV_X1 u1_u0_u3_U90 (.A( u1_u0_u3_n126 ) , .ZN( u1_u0_u3_n180 ) );
  INV_X1 u1_u0_u3_U91 (.A( u1_u0_u3_n112 ) , .ZN( u1_u0_u3_n175 ) );
  NAND4_X1 u1_u0_u3_U92 (.ZN( u1_out0_1 ) , .A4( u1_u0_u3_n161 ) , .A3( u1_u0_u3_n162 ) , .A2( u1_u0_u3_n163 ) , .A1( u1_u0_u3_n185 ) );
  NAND2_X1 u1_u0_u3_U93 (.ZN( u1_u0_u3_n163 ) , .A2( u1_u0_u3_n170 ) , .A1( u1_u0_u3_n176 ) );
  AOI22_X1 u1_u0_u3_U94 (.B2( u1_u0_u3_n140 ) , .B1( u1_u0_u3_n141 ) , .A2( u1_u0_u3_n142 ) , .ZN( u1_u0_u3_n162 ) , .A1( u1_u0_u3_n177 ) );
  OR4_X1 u1_u0_u3_U95 (.ZN( u1_out0_10 ) , .A4( u1_u0_u3_n136 ) , .A3( u1_u0_u3_n137 ) , .A1( u1_u0_u3_n138 ) , .A2( u1_u0_u3_n139 ) );
  OAI222_X1 u1_u0_u3_U96 (.C1( u1_u0_u3_n128 ) , .ZN( u1_u0_u3_n137 ) , .B1( u1_u0_u3_n148 ) , .A2( u1_u0_u3_n150 ) , .B2( u1_u0_u3_n154 ) , .C2( u1_u0_u3_n164 ) , .A1( u1_u0_u3_n167 ) );
  OAI221_X1 u1_u0_u3_U97 (.A( u1_u0_u3_n134 ) , .B2( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n136 ) , .C1( u1_u0_u3_n149 ) , .B1( u1_u0_u3_n151 ) , .C2( u1_u0_u3_n183 ) );
  NAND3_X1 u1_u0_u3_U98 (.A1( u1_u0_u3_n114 ) , .ZN( u1_u0_u3_n115 ) , .A2( u1_u0_u3_n145 ) , .A3( u1_u0_u3_n153 ) );
  NAND3_X1 u1_u0_u3_U99 (.ZN( u1_u0_u3_n129 ) , .A2( u1_u0_u3_n144 ) , .A1( u1_u0_u3_n153 ) , .A3( u1_u0_u3_n182 ) );
  XOR2_X1 u1_u10_U1 (.B( u1_K11_9 ) , .A( u1_R9_6 ) , .Z( u1_u10_X_9 ) );
  XOR2_X1 u1_u10_U16 (.B( u1_K11_3 ) , .A( u1_R9_2 ) , .Z( u1_u10_X_3 ) );
  XOR2_X1 u1_u10_U2 (.B( u1_K11_8 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_8 ) );
  XOR2_X1 u1_u10_U20 (.B( u1_K11_36 ) , .A( u1_R9_25 ) , .Z( u1_u10_X_36 ) );
  XOR2_X1 u1_u10_U21 (.B( u1_K11_35 ) , .A( u1_R9_24 ) , .Z( u1_u10_X_35 ) );
  XOR2_X1 u1_u10_U22 (.B( u1_K11_34 ) , .A( u1_R9_23 ) , .Z( u1_u10_X_34 ) );
  XOR2_X1 u1_u10_U23 (.B( u1_K11_33 ) , .A( u1_R9_22 ) , .Z( u1_u10_X_33 ) );
  XOR2_X1 u1_u10_U24 (.B( u1_K11_32 ) , .A( u1_R9_21 ) , .Z( u1_u10_X_32 ) );
  XOR2_X1 u1_u10_U25 (.B( u1_K11_31 ) , .A( u1_R9_20 ) , .Z( u1_u10_X_31 ) );
  XOR2_X1 u1_u10_U27 (.B( u1_K11_2 ) , .A( u1_R9_1 ) , .Z( u1_u10_X_2 ) );
  XOR2_X1 u1_u10_U3 (.B( u1_K11_7 ) , .A( u1_R9_4 ) , .Z( u1_u10_X_7 ) );
  XOR2_X1 u1_u10_U38 (.B( u1_K11_1 ) , .A( u1_R9_32 ) , .Z( u1_u10_X_1 ) );
  XOR2_X1 u1_u10_U4 (.B( u1_K11_6 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_6 ) );
  XOR2_X1 u1_u10_U40 (.B( u1_K11_18 ) , .A( u1_R9_13 ) , .Z( u1_u10_X_18 ) );
  XOR2_X1 u1_u10_U41 (.B( u1_K11_17 ) , .A( u1_R9_12 ) , .Z( u1_u10_X_17 ) );
  XOR2_X1 u1_u10_U42 (.B( u1_K11_16 ) , .A( u1_R9_11 ) , .Z( u1_u10_X_16 ) );
  XOR2_X1 u1_u10_U43 (.B( u1_K11_15 ) , .A( u1_R9_10 ) , .Z( u1_u10_X_15 ) );
  XOR2_X1 u1_u10_U44 (.B( u1_K11_14 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_14 ) );
  XOR2_X1 u1_u10_U45 (.B( u1_K11_13 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_13 ) );
  XOR2_X1 u1_u10_U46 (.B( u1_K11_12 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_12 ) );
  XOR2_X1 u1_u10_U47 (.B( u1_K11_11 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_11 ) );
  XOR2_X1 u1_u10_U48 (.B( u1_K11_10 ) , .A( u1_R9_7 ) , .Z( u1_u10_X_10 ) );
  XOR2_X1 u1_u10_U5 (.B( u1_K11_5 ) , .A( u1_R9_4 ) , .Z( u1_u10_X_5 ) );
  XOR2_X1 u1_u10_U6 (.B( u1_K11_4 ) , .A( u1_R9_3 ) , .Z( u1_u10_X_4 ) );
  AND3_X1 u1_u10_u0_U10 (.A2( u1_u10_u0_n112 ) , .ZN( u1_u10_u0_n127 ) , .A3( u1_u10_u0_n130 ) , .A1( u1_u10_u0_n148 ) );
  NAND2_X1 u1_u10_u0_U11 (.ZN( u1_u10_u0_n113 ) , .A1( u1_u10_u0_n139 ) , .A2( u1_u10_u0_n149 ) );
  AND2_X1 u1_u10_u0_U12 (.ZN( u1_u10_u0_n107 ) , .A1( u1_u10_u0_n130 ) , .A2( u1_u10_u0_n140 ) );
  AND2_X1 u1_u10_u0_U13 (.A2( u1_u10_u0_n129 ) , .A1( u1_u10_u0_n130 ) , .ZN( u1_u10_u0_n151 ) );
  AND2_X1 u1_u10_u0_U14 (.A1( u1_u10_u0_n108 ) , .A2( u1_u10_u0_n125 ) , .ZN( u1_u10_u0_n145 ) );
  INV_X1 u1_u10_u0_U15 (.A( u1_u10_u0_n143 ) , .ZN( u1_u10_u0_n173 ) );
  NOR2_X1 u1_u10_u0_U16 (.A2( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n147 ) , .A1( u1_u10_u0_n160 ) );
  NOR2_X1 u1_u10_u0_U17 (.A1( u1_u10_u0_n163 ) , .A2( u1_u10_u0_n164 ) , .ZN( u1_u10_u0_n95 ) );
  AOI21_X1 u1_u10_u0_U18 (.B1( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n132 ) , .A( u1_u10_u0_n165 ) , .B2( u1_u10_u0_n93 ) );
  INV_X1 u1_u10_u0_U19 (.A( u1_u10_u0_n142 ) , .ZN( u1_u10_u0_n165 ) );
  OAI221_X1 u1_u10_u0_U20 (.C1( u1_u10_u0_n121 ) , .ZN( u1_u10_u0_n122 ) , .B2( u1_u10_u0_n127 ) , .A( u1_u10_u0_n143 ) , .B1( u1_u10_u0_n144 ) , .C2( u1_u10_u0_n147 ) );
  OAI22_X1 u1_u10_u0_U21 (.B1( u1_u10_u0_n125 ) , .ZN( u1_u10_u0_n126 ) , .A1( u1_u10_u0_n138 ) , .A2( u1_u10_u0_n146 ) , .B2( u1_u10_u0_n147 ) );
  OAI22_X1 u1_u10_u0_U22 (.B1( u1_u10_u0_n131 ) , .A1( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n147 ) , .A2( u1_u10_u0_n90 ) , .ZN( u1_u10_u0_n91 ) );
  AND3_X1 u1_u10_u0_U23 (.A3( u1_u10_u0_n121 ) , .A2( u1_u10_u0_n125 ) , .A1( u1_u10_u0_n148 ) , .ZN( u1_u10_u0_n90 ) );
  INV_X1 u1_u10_u0_U24 (.A( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n161 ) );
  NOR2_X1 u1_u10_u0_U25 (.A1( u1_u10_u0_n120 ) , .ZN( u1_u10_u0_n143 ) , .A2( u1_u10_u0_n167 ) );
  OAI221_X1 u1_u10_u0_U26 (.C1( u1_u10_u0_n112 ) , .ZN( u1_u10_u0_n120 ) , .B1( u1_u10_u0_n138 ) , .B2( u1_u10_u0_n141 ) , .C2( u1_u10_u0_n147 ) , .A( u1_u10_u0_n172 ) );
  AOI22_X1 u1_u10_u0_U27 (.B2( u1_u10_u0_n109 ) , .A2( u1_u10_u0_n110 ) , .ZN( u1_u10_u0_n111 ) , .B1( u1_u10_u0_n118 ) , .A1( u1_u10_u0_n160 ) );
  INV_X1 u1_u10_u0_U28 (.A( u1_u10_u0_n118 ) , .ZN( u1_u10_u0_n158 ) );
  AOI21_X1 u1_u10_u0_U29 (.B1( u1_u10_u0_n132 ) , .ZN( u1_u10_u0_n133 ) , .A( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n166 ) );
  INV_X1 u1_u10_u0_U3 (.A( u1_u10_u0_n113 ) , .ZN( u1_u10_u0_n166 ) );
  AOI21_X1 u1_u10_u0_U30 (.ZN( u1_u10_u0_n104 ) , .B1( u1_u10_u0_n107 ) , .B2( u1_u10_u0_n141 ) , .A( u1_u10_u0_n144 ) );
  AOI21_X1 u1_u10_u0_U31 (.B1( u1_u10_u0_n127 ) , .B2( u1_u10_u0_n129 ) , .A( u1_u10_u0_n138 ) , .ZN( u1_u10_u0_n96 ) );
  AOI21_X1 u1_u10_u0_U32 (.ZN( u1_u10_u0_n116 ) , .B2( u1_u10_u0_n142 ) , .A( u1_u10_u0_n144 ) , .B1( u1_u10_u0_n166 ) );
  NAND2_X1 u1_u10_u0_U33 (.A1( u1_u10_u0_n100 ) , .A2( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n125 ) );
  NAND2_X1 u1_u10_u0_U34 (.A2( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n140 ) , .A1( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U35 (.A1( u1_u10_u0_n101 ) , .A2( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n150 ) );
  INV_X1 u1_u10_u0_U36 (.A( u1_u10_u0_n138 ) , .ZN( u1_u10_u0_n160 ) );
  NAND2_X1 u1_u10_u0_U37 (.ZN( u1_u10_u0_n142 ) , .A1( u1_u10_u0_n94 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U38 (.A1( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n128 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U39 (.A2( u1_u10_u0_n102 ) , .A1( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n149 ) );
  AOI21_X1 u1_u10_u0_U4 (.B2( u1_u10_u0_n131 ) , .ZN( u1_u10_u0_n134 ) , .B1( u1_u10_u0_n151 ) , .A( u1_u10_u0_n158 ) );
  NAND2_X1 u1_u10_u0_U40 (.A1( u1_u10_u0_n100 ) , .ZN( u1_u10_u0_n129 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U41 (.A2( u1_u10_u0_n100 ) , .A1( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n139 ) );
  NAND2_X1 u1_u10_u0_U42 (.A2( u1_u10_u0_n100 ) , .ZN( u1_u10_u0_n131 ) , .A1( u1_u10_u0_n92 ) );
  NAND2_X1 u1_u10_u0_U43 (.ZN( u1_u10_u0_n108 ) , .A1( u1_u10_u0_n92 ) , .A2( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U44 (.ZN( u1_u10_u0_n148 ) , .A1( u1_u10_u0_n93 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U45 (.A2( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n114 ) , .A1( u1_u10_u0_n92 ) );
  NAND2_X1 u1_u10_u0_U46 (.A1( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n130 ) , .A2( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U47 (.A2( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n121 ) , .A1( u1_u10_u0_n93 ) );
  INV_X1 u1_u10_u0_U48 (.ZN( u1_u10_u0_n172 ) , .A( u1_u10_u0_n88 ) );
  OAI222_X1 u1_u10_u0_U49 (.C1( u1_u10_u0_n108 ) , .A1( u1_u10_u0_n125 ) , .B2( u1_u10_u0_n128 ) , .B1( u1_u10_u0_n144 ) , .A2( u1_u10_u0_n158 ) , .C2( u1_u10_u0_n161 ) , .ZN( u1_u10_u0_n88 ) );
  NOR2_X1 u1_u10_u0_U5 (.A1( u1_u10_u0_n108 ) , .ZN( u1_u10_u0_n123 ) , .A2( u1_u10_u0_n158 ) );
  NAND2_X1 u1_u10_u0_U50 (.ZN( u1_u10_u0_n112 ) , .A2( u1_u10_u0_n92 ) , .A1( u1_u10_u0_n93 ) );
  OR3_X1 u1_u10_u0_U51 (.A3( u1_u10_u0_n152 ) , .A2( u1_u10_u0_n153 ) , .A1( u1_u10_u0_n154 ) , .ZN( u1_u10_u0_n155 ) );
  AOI21_X1 u1_u10_u0_U52 (.A( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n145 ) , .B1( u1_u10_u0_n146 ) , .ZN( u1_u10_u0_n154 ) );
  AOI21_X1 u1_u10_u0_U53 (.B2( u1_u10_u0_n150 ) , .B1( u1_u10_u0_n151 ) , .ZN( u1_u10_u0_n152 ) , .A( u1_u10_u0_n158 ) );
  AOI21_X1 u1_u10_u0_U54 (.A( u1_u10_u0_n147 ) , .B2( u1_u10_u0_n148 ) , .B1( u1_u10_u0_n149 ) , .ZN( u1_u10_u0_n153 ) );
  INV_X1 u1_u10_u0_U55 (.ZN( u1_u10_u0_n171 ) , .A( u1_u10_u0_n99 ) );
  OAI211_X1 u1_u10_u0_U56 (.C2( u1_u10_u0_n140 ) , .C1( u1_u10_u0_n161 ) , .A( u1_u10_u0_n169 ) , .B( u1_u10_u0_n98 ) , .ZN( u1_u10_u0_n99 ) );
  INV_X1 u1_u10_u0_U57 (.ZN( u1_u10_u0_n169 ) , .A( u1_u10_u0_n91 ) );
  AOI211_X1 u1_u10_u0_U58 (.C1( u1_u10_u0_n118 ) , .A( u1_u10_u0_n123 ) , .B( u1_u10_u0_n96 ) , .C2( u1_u10_u0_n97 ) , .ZN( u1_u10_u0_n98 ) );
  NOR2_X1 u1_u10_u0_U59 (.A2( u1_u10_X_2 ) , .ZN( u1_u10_u0_n103 ) , .A1( u1_u10_u0_n164 ) );
  OAI21_X1 u1_u10_u0_U6 (.B1( u1_u10_u0_n150 ) , .B2( u1_u10_u0_n158 ) , .A( u1_u10_u0_n172 ) , .ZN( u1_u10_u0_n89 ) );
  NOR2_X1 u1_u10_u0_U60 (.A2( u1_u10_X_3 ) , .A1( u1_u10_X_6 ) , .ZN( u1_u10_u0_n94 ) );
  NOR2_X1 u1_u10_u0_U61 (.A2( u1_u10_X_6 ) , .ZN( u1_u10_u0_n100 ) , .A1( u1_u10_u0_n162 ) );
  NOR2_X1 u1_u10_u0_U62 (.A2( u1_u10_X_1 ) , .A1( u1_u10_X_2 ) , .ZN( u1_u10_u0_n92 ) );
  NOR2_X1 u1_u10_u0_U63 (.A2( u1_u10_X_1 ) , .ZN( u1_u10_u0_n101 ) , .A1( u1_u10_u0_n163 ) );
  NOR2_X1 u1_u10_u0_U64 (.A2( u1_u10_X_4 ) , .A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n118 ) );
  NAND2_X1 u1_u10_u0_U65 (.A2( u1_u10_X_4 ) , .A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n144 ) );
  NOR2_X1 u1_u10_u0_U66 (.A2( u1_u10_X_5 ) , .ZN( u1_u10_u0_n136 ) , .A1( u1_u10_u0_n159 ) );
  NAND2_X1 u1_u10_u0_U67 (.A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n138 ) , .A2( u1_u10_u0_n159 ) );
  AND2_X1 u1_u10_u0_U68 (.A2( u1_u10_X_3 ) , .A1( u1_u10_X_6 ) , .ZN( u1_u10_u0_n102 ) );
  AND2_X1 u1_u10_u0_U69 (.A1( u1_u10_X_6 ) , .A2( u1_u10_u0_n162 ) , .ZN( u1_u10_u0_n93 ) );
  AOI21_X1 u1_u10_u0_U7 (.B1( u1_u10_u0_n114 ) , .ZN( u1_u10_u0_n115 ) , .B2( u1_u10_u0_n129 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U70 (.A( u1_u10_X_4 ) , .ZN( u1_u10_u0_n159 ) );
  INV_X1 u1_u10_u0_U71 (.A( u1_u10_X_1 ) , .ZN( u1_u10_u0_n164 ) );
  INV_X1 u1_u10_u0_U72 (.A( u1_u10_X_2 ) , .ZN( u1_u10_u0_n163 ) );
  INV_X1 u1_u10_u0_U73 (.A( u1_u10_X_3 ) , .ZN( u1_u10_u0_n162 ) );
  INV_X1 u1_u10_u0_U74 (.ZN( u1_u10_u0_n174 ) , .A( u1_u10_u0_n89 ) );
  AOI211_X1 u1_u10_u0_U75 (.B( u1_u10_u0_n104 ) , .A( u1_u10_u0_n105 ) , .ZN( u1_u10_u0_n106 ) , .C2( u1_u10_u0_n113 ) , .C1( u1_u10_u0_n160 ) );
  OR4_X1 u1_u10_u0_U76 (.ZN( u1_out10_17 ) , .A4( u1_u10_u0_n122 ) , .A2( u1_u10_u0_n123 ) , .A1( u1_u10_u0_n124 ) , .A3( u1_u10_u0_n170 ) );
  AOI21_X1 u1_u10_u0_U77 (.B2( u1_u10_u0_n107 ) , .ZN( u1_u10_u0_n124 ) , .B1( u1_u10_u0_n128 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U78 (.A( u1_u10_u0_n111 ) , .ZN( u1_u10_u0_n170 ) );
  OR4_X1 u1_u10_u0_U79 (.ZN( u1_out10_31 ) , .A4( u1_u10_u0_n155 ) , .A2( u1_u10_u0_n156 ) , .A1( u1_u10_u0_n157 ) , .A3( u1_u10_u0_n173 ) );
  AND2_X1 u1_u10_u0_U8 (.A1( u1_u10_u0_n114 ) , .A2( u1_u10_u0_n121 ) , .ZN( u1_u10_u0_n146 ) );
  AOI21_X1 u1_u10_u0_U80 (.A( u1_u10_u0_n138 ) , .B2( u1_u10_u0_n139 ) , .B1( u1_u10_u0_n140 ) , .ZN( u1_u10_u0_n157 ) );
  AOI21_X1 u1_u10_u0_U81 (.B2( u1_u10_u0_n141 ) , .B1( u1_u10_u0_n142 ) , .ZN( u1_u10_u0_n156 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U82 (.A( u1_u10_u0_n126 ) , .ZN( u1_u10_u0_n168 ) );
  AOI211_X1 u1_u10_u0_U83 (.B( u1_u10_u0_n133 ) , .A( u1_u10_u0_n134 ) , .C2( u1_u10_u0_n135 ) , .C1( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n137 ) );
  AOI211_X1 u1_u10_u0_U84 (.B( u1_u10_u0_n115 ) , .A( u1_u10_u0_n116 ) , .C2( u1_u10_u0_n117 ) , .C1( u1_u10_u0_n118 ) , .ZN( u1_u10_u0_n119 ) );
  INV_X1 u1_u10_u0_U85 (.A( u1_u10_u0_n119 ) , .ZN( u1_u10_u0_n167 ) );
  NAND2_X1 u1_u10_u0_U86 (.ZN( u1_u10_u0_n110 ) , .A2( u1_u10_u0_n132 ) , .A1( u1_u10_u0_n145 ) );
  OAI22_X1 u1_u10_u0_U87 (.ZN( u1_u10_u0_n105 ) , .A2( u1_u10_u0_n132 ) , .B1( u1_u10_u0_n146 ) , .A1( u1_u10_u0_n147 ) , .B2( u1_u10_u0_n161 ) );
  NAND3_X1 u1_u10_u0_U88 (.ZN( u1_out10_23 ) , .A3( u1_u10_u0_n137 ) , .A1( u1_u10_u0_n168 ) , .A2( u1_u10_u0_n171 ) );
  NAND3_X1 u1_u10_u0_U89 (.A3( u1_u10_u0_n127 ) , .A2( u1_u10_u0_n128 ) , .ZN( u1_u10_u0_n135 ) , .A1( u1_u10_u0_n150 ) );
  AND2_X1 u1_u10_u0_U9 (.A1( u1_u10_u0_n131 ) , .ZN( u1_u10_u0_n141 ) , .A2( u1_u10_u0_n150 ) );
  NAND3_X1 u1_u10_u0_U90 (.ZN( u1_u10_u0_n117 ) , .A3( u1_u10_u0_n132 ) , .A2( u1_u10_u0_n139 ) , .A1( u1_u10_u0_n148 ) );
  NAND3_X1 u1_u10_u0_U91 (.ZN( u1_u10_u0_n109 ) , .A2( u1_u10_u0_n114 ) , .A3( u1_u10_u0_n140 ) , .A1( u1_u10_u0_n149 ) );
  NAND3_X1 u1_u10_u0_U92 (.ZN( u1_out10_9 ) , .A3( u1_u10_u0_n106 ) , .A2( u1_u10_u0_n171 ) , .A1( u1_u10_u0_n174 ) );
  NAND3_X1 u1_u10_u0_U93 (.A2( u1_u10_u0_n128 ) , .A1( u1_u10_u0_n132 ) , .A3( u1_u10_u0_n146 ) , .ZN( u1_u10_u0_n97 ) );
  AOI21_X1 u1_u10_u1_U10 (.B2( u1_u10_u1_n155 ) , .B1( u1_u10_u1_n156 ) , .ZN( u1_u10_u1_n157 ) , .A( u1_u10_u1_n174 ) );
  NAND3_X1 u1_u10_u1_U100 (.ZN( u1_u10_u1_n113 ) , .A1( u1_u10_u1_n120 ) , .A3( u1_u10_u1_n133 ) , .A2( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U11 (.ZN( u1_u10_u1_n140 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U12 (.A1( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n153 ) );
  AOI22_X1 u1_u10_u1_U13 (.B2( u1_u10_u1_n136 ) , .A2( u1_u10_u1_n137 ) , .ZN( u1_u10_u1_n143 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U14 (.A( u1_u10_u1_n147 ) , .ZN( u1_u10_u1_n181 ) );
  INV_X1 u1_u10_u1_U15 (.A( u1_u10_u1_n139 ) , .ZN( u1_u10_u1_n174 ) );
  OR4_X1 u1_u10_u1_U16 (.A4( u1_u10_u1_n106 ) , .A3( u1_u10_u1_n107 ) , .ZN( u1_u10_u1_n108 ) , .A1( u1_u10_u1_n117 ) , .A2( u1_u10_u1_n184 ) );
  AOI21_X1 u1_u10_u1_U17 (.ZN( u1_u10_u1_n106 ) , .A( u1_u10_u1_n112 ) , .B1( u1_u10_u1_n154 ) , .B2( u1_u10_u1_n156 ) );
  AOI21_X1 u1_u10_u1_U18 (.ZN( u1_u10_u1_n107 ) , .B1( u1_u10_u1_n134 ) , .B2( u1_u10_u1_n149 ) , .A( u1_u10_u1_n174 ) );
  INV_X1 u1_u10_u1_U19 (.A( u1_u10_u1_n101 ) , .ZN( u1_u10_u1_n184 ) );
  INV_X1 u1_u10_u1_U20 (.A( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n171 ) );
  NAND2_X1 u1_u10_u1_U21 (.ZN( u1_u10_u1_n141 ) , .A1( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n156 ) );
  AND2_X1 u1_u10_u1_U22 (.A1( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n161 ) );
  NAND2_X1 u1_u10_u1_U23 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n148 ) );
  NAND2_X1 u1_u10_u1_U24 (.A2( u1_u10_u1_n133 ) , .A1( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n159 ) );
  NAND2_X1 u1_u10_u1_U25 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n120 ) , .ZN( u1_u10_u1_n132 ) );
  INV_X1 u1_u10_u1_U26 (.A( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n178 ) );
  INV_X1 u1_u10_u1_U27 (.A( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n183 ) );
  AND2_X1 u1_u10_u1_U28 (.A1( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n149 ) );
  INV_X1 u1_u10_u1_U29 (.A( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n180 ) );
  INV_X1 u1_u10_u1_U3 (.A( u1_u10_u1_n159 ) , .ZN( u1_u10_u1_n182 ) );
  OAI221_X1 u1_u10_u1_U30 (.A( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n138 ) , .B2( u1_u10_u1_n152 ) , .C1( u1_u10_u1_n174 ) , .B1( u1_u10_u1_n187 ) );
  INV_X1 u1_u10_u1_U31 (.A( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n187 ) );
  AOI211_X1 u1_u10_u1_U32 (.B( u1_u10_u1_n117 ) , .A( u1_u10_u1_n118 ) , .ZN( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n146 ) , .C1( u1_u10_u1_n159 ) );
  NOR2_X1 u1_u10_u1_U33 (.A1( u1_u10_u1_n168 ) , .A2( u1_u10_u1_n176 ) , .ZN( u1_u10_u1_n98 ) );
  AOI211_X1 u1_u10_u1_U34 (.B( u1_u10_u1_n162 ) , .A( u1_u10_u1_n163 ) , .C2( u1_u10_u1_n164 ) , .ZN( u1_u10_u1_n165 ) , .C1( u1_u10_u1_n171 ) );
  AOI21_X1 u1_u10_u1_U35 (.A( u1_u10_u1_n160 ) , .B2( u1_u10_u1_n161 ) , .ZN( u1_u10_u1_n162 ) , .B1( u1_u10_u1_n182 ) );
  OR2_X1 u1_u10_u1_U36 (.A2( u1_u10_u1_n157 ) , .A1( u1_u10_u1_n158 ) , .ZN( u1_u10_u1_n163 ) );
  OAI21_X1 u1_u10_u1_U37 (.B2( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n145 ) , .B1( u1_u10_u1_n160 ) , .A( u1_u10_u1_n185 ) );
  INV_X1 u1_u10_u1_U38 (.A( u1_u10_u1_n122 ) , .ZN( u1_u10_u1_n185 ) );
  AOI21_X1 u1_u10_u1_U39 (.B2( u1_u10_u1_n120 ) , .B1( u1_u10_u1_n121 ) , .ZN( u1_u10_u1_n122 ) , .A( u1_u10_u1_n128 ) );
  AOI221_X1 u1_u10_u1_U4 (.A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .C1( u1_u10_u1_n140 ) , .B2( u1_u10_u1_n141 ) , .ZN( u1_u10_u1_n142 ) , .B1( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U40 (.A1( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n146 ) , .A2( u1_u10_u1_n160 ) );
  NAND2_X1 u1_u10_u1_U41 (.A2( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n139 ) , .A1( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U42 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n156 ) , .A2( u1_u10_u1_n99 ) );
  AOI221_X1 u1_u10_u1_U43 (.B1( u1_u10_u1_n140 ) , .ZN( u1_u10_u1_n167 ) , .B2( u1_u10_u1_n172 ) , .C2( u1_u10_u1_n175 ) , .C1( u1_u10_u1_n178 ) , .A( u1_u10_u1_n188 ) );
  INV_X1 u1_u10_u1_U44 (.ZN( u1_u10_u1_n188 ) , .A( u1_u10_u1_n97 ) );
  AOI211_X1 u1_u10_u1_U45 (.A( u1_u10_u1_n118 ) , .C1( u1_u10_u1_n132 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n96 ) , .ZN( u1_u10_u1_n97 ) );
  AOI21_X1 u1_u10_u1_U46 (.B2( u1_u10_u1_n121 ) , .B1( u1_u10_u1_n135 ) , .A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n96 ) );
  NOR2_X1 u1_u10_u1_U47 (.ZN( u1_u10_u1_n117 ) , .A1( u1_u10_u1_n121 ) , .A2( u1_u10_u1_n160 ) );
  AOI21_X1 u1_u10_u1_U48 (.A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n130 ) , .B1( u1_u10_u1_n150 ) );
  NAND2_X1 u1_u10_u1_U49 (.ZN( u1_u10_u1_n112 ) , .A1( u1_u10_u1_n169 ) , .A2( u1_u10_u1_n170 ) );
  AOI211_X1 u1_u10_u1_U5 (.ZN( u1_u10_u1_n124 ) , .A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n145 ) , .C1( u1_u10_u1_n147 ) );
  NAND2_X1 u1_u10_u1_U50 (.ZN( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n95 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U51 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n154 ) , .A2( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U52 (.A2( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n135 ) , .A1( u1_u10_u1_n99 ) );
  AOI21_X1 u1_u10_u1_U53 (.A( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n153 ) , .B1( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n158 ) );
  INV_X1 u1_u10_u1_U54 (.A( u1_u10_u1_n160 ) , .ZN( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U55 (.A1( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n116 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U56 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n131 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U57 (.A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n121 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U58 (.A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U59 (.A2( u1_u10_u1_n104 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n133 ) );
  AOI22_X1 u1_u10_u1_U6 (.B2( u1_u10_u1_n113 ) , .A2( u1_u10_u1_n114 ) , .ZN( u1_u10_u1_n125 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  NAND2_X1 u1_u10_u1_U60 (.ZN( u1_u10_u1_n150 ) , .A2( u1_u10_u1_n98 ) , .A1( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U61 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n155 ) , .A2( u1_u10_u1_n95 ) );
  OAI21_X1 u1_u10_u1_U62 (.ZN( u1_u10_u1_n109 ) , .B1( u1_u10_u1_n129 ) , .B2( u1_u10_u1_n160 ) , .A( u1_u10_u1_n167 ) );
  NAND2_X1 u1_u10_u1_U63 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n120 ) );
  NAND2_X1 u1_u10_u1_U64 (.A1( u1_u10_u1_n102 ) , .A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n115 ) );
  NAND2_X1 u1_u10_u1_U65 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n151 ) );
  NAND2_X1 u1_u10_u1_U66 (.A2( u1_u10_u1_n103 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n161 ) );
  INV_X1 u1_u10_u1_U67 (.A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U68 (.A( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n172 ) );
  NAND2_X1 u1_u10_u1_U69 (.A2( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n123 ) );
  NAND2_X1 u1_u10_u1_U7 (.ZN( u1_u10_u1_n114 ) , .A1( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n156 ) );
  NOR2_X1 u1_u10_u1_U70 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n95 ) );
  NOR2_X1 u1_u10_u1_U71 (.A1( u1_u10_X_12 ) , .A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n100 ) );
  NOR2_X1 u1_u10_u1_U72 (.A2( u1_u10_X_8 ) , .A1( u1_u10_u1_n177 ) , .ZN( u1_u10_u1_n99 ) );
  NOR2_X1 u1_u10_u1_U73 (.A2( u1_u10_X_12 ) , .ZN( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n176 ) );
  NOR2_X1 u1_u10_u1_U74 (.A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n105 ) , .A1( u1_u10_u1_n168 ) );
  NAND2_X1 u1_u10_u1_U75 (.A1( u1_u10_X_10 ) , .ZN( u1_u10_u1_n160 ) , .A2( u1_u10_u1_n169 ) );
  NAND2_X1 u1_u10_u1_U76 (.A2( u1_u10_X_10 ) , .A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U77 (.A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n128 ) , .A2( u1_u10_u1_n170 ) );
  AND2_X1 u1_u10_u1_U78 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n104 ) );
  AND2_X1 u1_u10_u1_U79 (.A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n103 ) , .A2( u1_u10_u1_n177 ) );
  NOR2_X1 u1_u10_u1_U8 (.A1( u1_u10_u1_n112 ) , .A2( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n118 ) );
  INV_X1 u1_u10_u1_U80 (.A( u1_u10_X_10 ) , .ZN( u1_u10_u1_n170 ) );
  INV_X1 u1_u10_u1_U81 (.A( u1_u10_X_9 ) , .ZN( u1_u10_u1_n176 ) );
  INV_X1 u1_u10_u1_U82 (.A( u1_u10_X_11 ) , .ZN( u1_u10_u1_n169 ) );
  INV_X1 u1_u10_u1_U83 (.A( u1_u10_X_12 ) , .ZN( u1_u10_u1_n168 ) );
  INV_X1 u1_u10_u1_U84 (.A( u1_u10_X_7 ) , .ZN( u1_u10_u1_n177 ) );
  NAND4_X1 u1_u10_u1_U85 (.ZN( u1_out10_18 ) , .A4( u1_u10_u1_n165 ) , .A3( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n167 ) , .A2( u1_u10_u1_n186 ) );
  AOI22_X1 u1_u10_u1_U86 (.B2( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n172 ) );
  INV_X1 u1_u10_u1_U87 (.A( u1_u10_u1_n145 ) , .ZN( u1_u10_u1_n186 ) );
  NAND4_X1 u1_u10_u1_U88 (.ZN( u1_out10_2 ) , .A4( u1_u10_u1_n142 ) , .A3( u1_u10_u1_n143 ) , .A2( u1_u10_u1_n144 ) , .A1( u1_u10_u1_n179 ) );
  OAI21_X1 u1_u10_u1_U89 (.B2( u1_u10_u1_n132 ) , .ZN( u1_u10_u1_n144 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n180 ) );
  OAI21_X1 u1_u10_u1_U9 (.ZN( u1_u10_u1_n101 ) , .B1( u1_u10_u1_n141 ) , .A( u1_u10_u1_n146 ) , .B2( u1_u10_u1_n183 ) );
  INV_X1 u1_u10_u1_U90 (.A( u1_u10_u1_n130 ) , .ZN( u1_u10_u1_n179 ) );
  OR4_X1 u1_u10_u1_U91 (.ZN( u1_out10_13 ) , .A4( u1_u10_u1_n108 ) , .A3( u1_u10_u1_n109 ) , .A2( u1_u10_u1_n110 ) , .A1( u1_u10_u1_n111 ) );
  AOI21_X1 u1_u10_u1_U92 (.ZN( u1_u10_u1_n111 ) , .A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n131 ) , .B1( u1_u10_u1_n135 ) );
  AOI21_X1 u1_u10_u1_U93 (.ZN( u1_u10_u1_n110 ) , .A( u1_u10_u1_n116 ) , .B1( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n160 ) );
  NAND4_X1 u1_u10_u1_U94 (.ZN( u1_out10_28 ) , .A4( u1_u10_u1_n124 ) , .A3( u1_u10_u1_n125 ) , .A2( u1_u10_u1_n126 ) , .A1( u1_u10_u1_n127 ) );
  OAI21_X1 u1_u10_u1_U95 (.ZN( u1_u10_u1_n127 ) , .B2( u1_u10_u1_n139 ) , .B1( u1_u10_u1_n175 ) , .A( u1_u10_u1_n183 ) );
  OAI21_X1 u1_u10_u1_U96 (.ZN( u1_u10_u1_n126 ) , .B2( u1_u10_u1_n140 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n178 ) );
  NAND3_X1 u1_u10_u1_U97 (.A3( u1_u10_u1_n149 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n164 ) );
  NAND3_X1 u1_u10_u1_U98 (.A3( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n136 ) , .A1( u1_u10_u1_n151 ) );
  NAND3_X1 u1_u10_u1_U99 (.A1( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n137 ) , .A2( u1_u10_u1_n154 ) , .A3( u1_u10_u1_n181 ) );
  OAI22_X1 u1_u10_u2_U10 (.ZN( u1_u10_u2_n109 ) , .A2( u1_u10_u2_n113 ) , .B2( u1_u10_u2_n133 ) , .B1( u1_u10_u2_n167 ) , .A1( u1_u10_u2_n168 ) );
  NAND3_X1 u1_u10_u2_U100 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n98 ) );
  OAI22_X1 u1_u10_u2_U11 (.B1( u1_u10_u2_n151 ) , .A2( u1_u10_u2_n152 ) , .A1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n160 ) , .B2( u1_u10_u2_n168 ) );
  NOR3_X1 u1_u10_u2_U12 (.A1( u1_u10_u2_n150 ) , .ZN( u1_u10_u2_n151 ) , .A3( u1_u10_u2_n175 ) , .A2( u1_u10_u2_n188 ) );
  AOI21_X1 u1_u10_u2_U13 (.ZN( u1_u10_u2_n144 ) , .B2( u1_u10_u2_n155 ) , .A( u1_u10_u2_n172 ) , .B1( u1_u10_u2_n185 ) );
  AOI21_X1 u1_u10_u2_U14 (.B2( u1_u10_u2_n143 ) , .ZN( u1_u10_u2_n145 ) , .B1( u1_u10_u2_n152 ) , .A( u1_u10_u2_n171 ) );
  AOI21_X1 u1_u10_u2_U15 (.B2( u1_u10_u2_n120 ) , .B1( u1_u10_u2_n121 ) , .ZN( u1_u10_u2_n126 ) , .A( u1_u10_u2_n167 ) );
  INV_X1 u1_u10_u2_U16 (.A( u1_u10_u2_n156 ) , .ZN( u1_u10_u2_n171 ) );
  INV_X1 u1_u10_u2_U17 (.A( u1_u10_u2_n120 ) , .ZN( u1_u10_u2_n188 ) );
  NAND2_X1 u1_u10_u2_U18 (.A2( u1_u10_u2_n122 ) , .ZN( u1_u10_u2_n150 ) , .A1( u1_u10_u2_n152 ) );
  INV_X1 u1_u10_u2_U19 (.A( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n170 ) );
  INV_X1 u1_u10_u2_U20 (.A( u1_u10_u2_n137 ) , .ZN( u1_u10_u2_n173 ) );
  NAND2_X1 u1_u10_u2_U21 (.A1( u1_u10_u2_n132 ) , .A2( u1_u10_u2_n139 ) , .ZN( u1_u10_u2_n157 ) );
  INV_X1 u1_u10_u2_U22 (.A( u1_u10_u2_n113 ) , .ZN( u1_u10_u2_n178 ) );
  INV_X1 u1_u10_u2_U23 (.A( u1_u10_u2_n139 ) , .ZN( u1_u10_u2_n175 ) );
  INV_X1 u1_u10_u2_U24 (.A( u1_u10_u2_n155 ) , .ZN( u1_u10_u2_n181 ) );
  INV_X1 u1_u10_u2_U25 (.A( u1_u10_u2_n119 ) , .ZN( u1_u10_u2_n177 ) );
  INV_X1 u1_u10_u2_U26 (.A( u1_u10_u2_n116 ) , .ZN( u1_u10_u2_n180 ) );
  INV_X1 u1_u10_u2_U27 (.A( u1_u10_u2_n131 ) , .ZN( u1_u10_u2_n179 ) );
  INV_X1 u1_u10_u2_U28 (.A( u1_u10_u2_n154 ) , .ZN( u1_u10_u2_n176 ) );
  NAND2_X1 u1_u10_u2_U29 (.A2( u1_u10_u2_n116 ) , .A1( u1_u10_u2_n117 ) , .ZN( u1_u10_u2_n118 ) );
  NOR2_X1 u1_u10_u2_U3 (.ZN( u1_u10_u2_n121 ) , .A2( u1_u10_u2_n177 ) , .A1( u1_u10_u2_n180 ) );
  INV_X1 u1_u10_u2_U30 (.A( u1_u10_u2_n132 ) , .ZN( u1_u10_u2_n182 ) );
  INV_X1 u1_u10_u2_U31 (.A( u1_u10_u2_n158 ) , .ZN( u1_u10_u2_n183 ) );
  OAI21_X1 u1_u10_u2_U32 (.A( u1_u10_u2_n156 ) , .B1( u1_u10_u2_n157 ) , .ZN( u1_u10_u2_n158 ) , .B2( u1_u10_u2_n179 ) );
  NOR2_X1 u1_u10_u2_U33 (.ZN( u1_u10_u2_n156 ) , .A1( u1_u10_u2_n166 ) , .A2( u1_u10_u2_n169 ) );
  NOR2_X1 u1_u10_u2_U34 (.A2( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n137 ) , .A1( u1_u10_u2_n140 ) );
  NOR2_X1 u1_u10_u2_U35 (.A2( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n153 ) , .A1( u1_u10_u2_n156 ) );
  AOI211_X1 u1_u10_u2_U36 (.ZN( u1_u10_u2_n130 ) , .C1( u1_u10_u2_n138 ) , .C2( u1_u10_u2_n179 ) , .B( u1_u10_u2_n96 ) , .A( u1_u10_u2_n97 ) );
  OAI22_X1 u1_u10_u2_U37 (.B1( u1_u10_u2_n133 ) , .A2( u1_u10_u2_n137 ) , .A1( u1_u10_u2_n152 ) , .B2( u1_u10_u2_n168 ) , .ZN( u1_u10_u2_n97 ) );
  OAI221_X1 u1_u10_u2_U38 (.B1( u1_u10_u2_n113 ) , .C1( u1_u10_u2_n132 ) , .A( u1_u10_u2_n149 ) , .B2( u1_u10_u2_n171 ) , .C2( u1_u10_u2_n172 ) , .ZN( u1_u10_u2_n96 ) );
  OAI221_X1 u1_u10_u2_U39 (.A( u1_u10_u2_n115 ) , .C2( u1_u10_u2_n123 ) , .B2( u1_u10_u2_n143 ) , .B1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n163 ) , .C1( u1_u10_u2_n168 ) );
  INV_X1 u1_u10_u2_U4 (.A( u1_u10_u2_n134 ) , .ZN( u1_u10_u2_n185 ) );
  OAI21_X1 u1_u10_u2_U40 (.A( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n115 ) , .B1( u1_u10_u2_n176 ) , .B2( u1_u10_u2_n178 ) );
  OAI221_X1 u1_u10_u2_U41 (.A( u1_u10_u2_n135 ) , .B2( u1_u10_u2_n136 ) , .B1( u1_u10_u2_n137 ) , .ZN( u1_u10_u2_n162 ) , .C2( u1_u10_u2_n167 ) , .C1( u1_u10_u2_n185 ) );
  AND3_X1 u1_u10_u2_U42 (.A3( u1_u10_u2_n131 ) , .A2( u1_u10_u2_n132 ) , .A1( u1_u10_u2_n133 ) , .ZN( u1_u10_u2_n136 ) );
  AOI22_X1 u1_u10_u2_U43 (.ZN( u1_u10_u2_n135 ) , .B1( u1_u10_u2_n140 ) , .A1( u1_u10_u2_n156 ) , .B2( u1_u10_u2_n180 ) , .A2( u1_u10_u2_n188 ) );
  AOI21_X1 u1_u10_u2_U44 (.ZN( u1_u10_u2_n149 ) , .B1( u1_u10_u2_n173 ) , .B2( u1_u10_u2_n188 ) , .A( u1_u10_u2_n95 ) );
  AND3_X1 u1_u10_u2_U45 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n156 ) , .ZN( u1_u10_u2_n95 ) );
  OAI21_X1 u1_u10_u2_U46 (.A( u1_u10_u2_n101 ) , .B2( u1_u10_u2_n121 ) , .B1( u1_u10_u2_n153 ) , .ZN( u1_u10_u2_n164 ) );
  NAND2_X1 u1_u10_u2_U47 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n155 ) );
  NAND2_X1 u1_u10_u2_U48 (.A2( u1_u10_u2_n105 ) , .A1( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n143 ) );
  NAND2_X1 u1_u10_u2_U49 (.A1( u1_u10_u2_n104 ) , .A2( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n152 ) );
  INV_X1 u1_u10_u2_U5 (.A( u1_u10_u2_n150 ) , .ZN( u1_u10_u2_n184 ) );
  NAND2_X1 u1_u10_u2_U50 (.A1( u1_u10_u2_n100 ) , .A2( u1_u10_u2_n105 ) , .ZN( u1_u10_u2_n132 ) );
  INV_X1 u1_u10_u2_U51 (.A( u1_u10_u2_n140 ) , .ZN( u1_u10_u2_n168 ) );
  INV_X1 u1_u10_u2_U52 (.A( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n167 ) );
  OAI21_X1 u1_u10_u2_U53 (.A( u1_u10_u2_n141 ) , .B2( u1_u10_u2_n142 ) , .ZN( u1_u10_u2_n146 ) , .B1( u1_u10_u2_n153 ) );
  OAI21_X1 u1_u10_u2_U54 (.A( u1_u10_u2_n140 ) , .ZN( u1_u10_u2_n141 ) , .B1( u1_u10_u2_n176 ) , .B2( u1_u10_u2_n177 ) );
  NOR3_X1 u1_u10_u2_U55 (.ZN( u1_u10_u2_n142 ) , .A3( u1_u10_u2_n175 ) , .A2( u1_u10_u2_n178 ) , .A1( u1_u10_u2_n181 ) );
  NAND2_X1 u1_u10_u2_U56 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n113 ) );
  NAND2_X1 u1_u10_u2_U57 (.A1( u1_u10_u2_n106 ) , .A2( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n131 ) );
  NAND2_X1 u1_u10_u2_U58 (.A1( u1_u10_u2_n103 ) , .A2( u1_u10_u2_n107 ) , .ZN( u1_u10_u2_n139 ) );
  NAND2_X1 u1_u10_u2_U59 (.A1( u1_u10_u2_n103 ) , .A2( u1_u10_u2_n105 ) , .ZN( u1_u10_u2_n133 ) );
  NOR4_X1 u1_u10_u2_U6 (.A4( u1_u10_u2_n124 ) , .A3( u1_u10_u2_n125 ) , .A2( u1_u10_u2_n126 ) , .A1( u1_u10_u2_n127 ) , .ZN( u1_u10_u2_n128 ) );
  NAND2_X1 u1_u10_u2_U60 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n103 ) , .ZN( u1_u10_u2_n154 ) );
  NAND2_X1 u1_u10_u2_U61 (.A2( u1_u10_u2_n103 ) , .A1( u1_u10_u2_n104 ) , .ZN( u1_u10_u2_n119 ) );
  NAND2_X1 u1_u10_u2_U62 (.A2( u1_u10_u2_n107 ) , .A1( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n123 ) );
  NAND2_X1 u1_u10_u2_U63 (.A1( u1_u10_u2_n104 ) , .A2( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n122 ) );
  INV_X1 u1_u10_u2_U64 (.A( u1_u10_u2_n114 ) , .ZN( u1_u10_u2_n172 ) );
  NAND2_X1 u1_u10_u2_U65 (.A2( u1_u10_u2_n100 ) , .A1( u1_u10_u2_n102 ) , .ZN( u1_u10_u2_n116 ) );
  NAND2_X1 u1_u10_u2_U66 (.A1( u1_u10_u2_n102 ) , .A2( u1_u10_u2_n108 ) , .ZN( u1_u10_u2_n120 ) );
  NAND2_X1 u1_u10_u2_U67 (.A2( u1_u10_u2_n105 ) , .A1( u1_u10_u2_n106 ) , .ZN( u1_u10_u2_n117 ) );
  INV_X1 u1_u10_u2_U68 (.ZN( u1_u10_u2_n187 ) , .A( u1_u10_u2_n99 ) );
  OAI21_X1 u1_u10_u2_U69 (.B1( u1_u10_u2_n137 ) , .B2( u1_u10_u2_n143 ) , .A( u1_u10_u2_n98 ) , .ZN( u1_u10_u2_n99 ) );
  AOI21_X1 u1_u10_u2_U7 (.ZN( u1_u10_u2_n124 ) , .B1( u1_u10_u2_n131 ) , .B2( u1_u10_u2_n143 ) , .A( u1_u10_u2_n172 ) );
  NOR2_X1 u1_u10_u2_U70 (.A2( u1_u10_X_16 ) , .ZN( u1_u10_u2_n140 ) , .A1( u1_u10_u2_n166 ) );
  NOR2_X1 u1_u10_u2_U71 (.A2( u1_u10_X_13 ) , .A1( u1_u10_X_14 ) , .ZN( u1_u10_u2_n100 ) );
  NOR2_X1 u1_u10_u2_U72 (.A2( u1_u10_X_16 ) , .A1( u1_u10_X_17 ) , .ZN( u1_u10_u2_n138 ) );
  NOR2_X1 u1_u10_u2_U73 (.A2( u1_u10_X_15 ) , .A1( u1_u10_X_18 ) , .ZN( u1_u10_u2_n104 ) );
  NOR2_X1 u1_u10_u2_U74 (.A2( u1_u10_X_14 ) , .ZN( u1_u10_u2_n103 ) , .A1( u1_u10_u2_n174 ) );
  NOR2_X1 u1_u10_u2_U75 (.A2( u1_u10_X_15 ) , .ZN( u1_u10_u2_n102 ) , .A1( u1_u10_u2_n165 ) );
  NOR2_X1 u1_u10_u2_U76 (.A2( u1_u10_X_17 ) , .ZN( u1_u10_u2_n114 ) , .A1( u1_u10_u2_n169 ) );
  AND2_X1 u1_u10_u2_U77 (.A1( u1_u10_X_15 ) , .ZN( u1_u10_u2_n105 ) , .A2( u1_u10_u2_n165 ) );
  AND2_X1 u1_u10_u2_U78 (.A2( u1_u10_X_15 ) , .A1( u1_u10_X_18 ) , .ZN( u1_u10_u2_n107 ) );
  AND2_X1 u1_u10_u2_U79 (.A1( u1_u10_X_14 ) , .ZN( u1_u10_u2_n106 ) , .A2( u1_u10_u2_n174 ) );
  AOI21_X1 u1_u10_u2_U8 (.B2( u1_u10_u2_n119 ) , .ZN( u1_u10_u2_n127 ) , .A( u1_u10_u2_n137 ) , .B1( u1_u10_u2_n155 ) );
  AND2_X1 u1_u10_u2_U80 (.A1( u1_u10_X_13 ) , .A2( u1_u10_X_14 ) , .ZN( u1_u10_u2_n108 ) );
  INV_X1 u1_u10_u2_U81 (.A( u1_u10_X_16 ) , .ZN( u1_u10_u2_n169 ) );
  INV_X1 u1_u10_u2_U82 (.A( u1_u10_X_17 ) , .ZN( u1_u10_u2_n166 ) );
  INV_X1 u1_u10_u2_U83 (.A( u1_u10_X_13 ) , .ZN( u1_u10_u2_n174 ) );
  INV_X1 u1_u10_u2_U84 (.A( u1_u10_X_18 ) , .ZN( u1_u10_u2_n165 ) );
  NAND4_X1 u1_u10_u2_U85 (.ZN( u1_out10_30 ) , .A4( u1_u10_u2_n147 ) , .A3( u1_u10_u2_n148 ) , .A2( u1_u10_u2_n149 ) , .A1( u1_u10_u2_n187 ) );
  NOR3_X1 u1_u10_u2_U86 (.A3( u1_u10_u2_n144 ) , .A2( u1_u10_u2_n145 ) , .A1( u1_u10_u2_n146 ) , .ZN( u1_u10_u2_n147 ) );
  AOI21_X1 u1_u10_u2_U87 (.B2( u1_u10_u2_n138 ) , .ZN( u1_u10_u2_n148 ) , .A( u1_u10_u2_n162 ) , .B1( u1_u10_u2_n182 ) );
  NAND4_X1 u1_u10_u2_U88 (.ZN( u1_out10_24 ) , .A4( u1_u10_u2_n111 ) , .A3( u1_u10_u2_n112 ) , .A1( u1_u10_u2_n130 ) , .A2( u1_u10_u2_n187 ) );
  AOI221_X1 u1_u10_u2_U89 (.A( u1_u10_u2_n109 ) , .B1( u1_u10_u2_n110 ) , .ZN( u1_u10_u2_n111 ) , .C1( u1_u10_u2_n134 ) , .C2( u1_u10_u2_n170 ) , .B2( u1_u10_u2_n173 ) );
  AOI21_X1 u1_u10_u2_U9 (.B2( u1_u10_u2_n123 ) , .ZN( u1_u10_u2_n125 ) , .A( u1_u10_u2_n171 ) , .B1( u1_u10_u2_n184 ) );
  AOI21_X1 u1_u10_u2_U90 (.ZN( u1_u10_u2_n112 ) , .B2( u1_u10_u2_n156 ) , .A( u1_u10_u2_n164 ) , .B1( u1_u10_u2_n181 ) );
  NAND4_X1 u1_u10_u2_U91 (.ZN( u1_out10_16 ) , .A4( u1_u10_u2_n128 ) , .A3( u1_u10_u2_n129 ) , .A1( u1_u10_u2_n130 ) , .A2( u1_u10_u2_n186 ) );
  AOI22_X1 u1_u10_u2_U92 (.A2( u1_u10_u2_n118 ) , .ZN( u1_u10_u2_n129 ) , .A1( u1_u10_u2_n140 ) , .B1( u1_u10_u2_n157 ) , .B2( u1_u10_u2_n170 ) );
  INV_X1 u1_u10_u2_U93 (.A( u1_u10_u2_n163 ) , .ZN( u1_u10_u2_n186 ) );
  OR4_X1 u1_u10_u2_U94 (.ZN( u1_out10_6 ) , .A4( u1_u10_u2_n161 ) , .A3( u1_u10_u2_n162 ) , .A2( u1_u10_u2_n163 ) , .A1( u1_u10_u2_n164 ) );
  OR3_X1 u1_u10_u2_U95 (.A2( u1_u10_u2_n159 ) , .A1( u1_u10_u2_n160 ) , .ZN( u1_u10_u2_n161 ) , .A3( u1_u10_u2_n183 ) );
  AOI21_X1 u1_u10_u2_U96 (.B2( u1_u10_u2_n154 ) , .B1( u1_u10_u2_n155 ) , .ZN( u1_u10_u2_n159 ) , .A( u1_u10_u2_n167 ) );
  NAND3_X1 u1_u10_u2_U97 (.A2( u1_u10_u2_n117 ) , .A1( u1_u10_u2_n122 ) , .A3( u1_u10_u2_n123 ) , .ZN( u1_u10_u2_n134 ) );
  NAND3_X1 u1_u10_u2_U98 (.ZN( u1_u10_u2_n110 ) , .A2( u1_u10_u2_n131 ) , .A3( u1_u10_u2_n139 ) , .A1( u1_u10_u2_n154 ) );
  NAND3_X1 u1_u10_u2_U99 (.A2( u1_u10_u2_n100 ) , .ZN( u1_u10_u2_n101 ) , .A1( u1_u10_u2_n104 ) , .A3( u1_u10_u2_n114 ) );
  INV_X1 u1_u10_u5_U10 (.A( u1_u10_u5_n121 ) , .ZN( u1_u10_u5_n177 ) );
  NOR3_X1 u1_u10_u5_U100 (.A3( u1_u10_u5_n141 ) , .A1( u1_u10_u5_n142 ) , .ZN( u1_u10_u5_n143 ) , .A2( u1_u10_u5_n191 ) );
  NAND4_X1 u1_u10_u5_U101 (.ZN( u1_out10_4 ) , .A4( u1_u10_u5_n112 ) , .A2( u1_u10_u5_n113 ) , .A1( u1_u10_u5_n114 ) , .A3( u1_u10_u5_n195 ) );
  AOI211_X1 u1_u10_u5_U102 (.A( u1_u10_u5_n110 ) , .C1( u1_u10_u5_n111 ) , .ZN( u1_u10_u5_n112 ) , .B( u1_u10_u5_n118 ) , .C2( u1_u10_u5_n177 ) );
  AOI222_X1 u1_u10_u5_U103 (.ZN( u1_u10_u5_n113 ) , .A1( u1_u10_u5_n131 ) , .C1( u1_u10_u5_n148 ) , .B2( u1_u10_u5_n174 ) , .C2( u1_u10_u5_n178 ) , .A2( u1_u10_u5_n179 ) , .B1( u1_u10_u5_n99 ) );
  NAND3_X1 u1_u10_u5_U104 (.A2( u1_u10_u5_n154 ) , .A3( u1_u10_u5_n158 ) , .A1( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n99 ) );
  NOR2_X1 u1_u10_u5_U11 (.ZN( u1_u10_u5_n160 ) , .A2( u1_u10_u5_n173 ) , .A1( u1_u10_u5_n177 ) );
  INV_X1 u1_u10_u5_U12 (.A( u1_u10_u5_n150 ) , .ZN( u1_u10_u5_n174 ) );
  AOI21_X1 u1_u10_u5_U13 (.A( u1_u10_u5_n160 ) , .B2( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n162 ) , .B1( u1_u10_u5_n192 ) );
  INV_X1 u1_u10_u5_U14 (.A( u1_u10_u5_n159 ) , .ZN( u1_u10_u5_n192 ) );
  AOI21_X1 u1_u10_u5_U15 (.A( u1_u10_u5_n156 ) , .B2( u1_u10_u5_n157 ) , .B1( u1_u10_u5_n158 ) , .ZN( u1_u10_u5_n163 ) );
  AOI21_X1 u1_u10_u5_U16 (.B2( u1_u10_u5_n139 ) , .B1( u1_u10_u5_n140 ) , .ZN( u1_u10_u5_n141 ) , .A( u1_u10_u5_n150 ) );
  OAI21_X1 u1_u10_u5_U17 (.A( u1_u10_u5_n133 ) , .B2( u1_u10_u5_n134 ) , .B1( u1_u10_u5_n135 ) , .ZN( u1_u10_u5_n142 ) );
  OAI21_X1 u1_u10_u5_U18 (.ZN( u1_u10_u5_n133 ) , .B2( u1_u10_u5_n147 ) , .A( u1_u10_u5_n173 ) , .B1( u1_u10_u5_n188 ) );
  NAND2_X1 u1_u10_u5_U19 (.A2( u1_u10_u5_n119 ) , .A1( u1_u10_u5_n123 ) , .ZN( u1_u10_u5_n137 ) );
  INV_X1 u1_u10_u5_U20 (.A( u1_u10_u5_n155 ) , .ZN( u1_u10_u5_n194 ) );
  NAND2_X1 u1_u10_u5_U21 (.A1( u1_u10_u5_n121 ) , .ZN( u1_u10_u5_n132 ) , .A2( u1_u10_u5_n172 ) );
  NAND2_X1 u1_u10_u5_U22 (.A2( u1_u10_u5_n122 ) , .ZN( u1_u10_u5_n136 ) , .A1( u1_u10_u5_n154 ) );
  NAND2_X1 u1_u10_u5_U23 (.A2( u1_u10_u5_n119 ) , .A1( u1_u10_u5_n120 ) , .ZN( u1_u10_u5_n159 ) );
  INV_X1 u1_u10_u5_U24 (.A( u1_u10_u5_n156 ) , .ZN( u1_u10_u5_n175 ) );
  INV_X1 u1_u10_u5_U25 (.A( u1_u10_u5_n158 ) , .ZN( u1_u10_u5_n188 ) );
  INV_X1 u1_u10_u5_U26 (.A( u1_u10_u5_n152 ) , .ZN( u1_u10_u5_n179 ) );
  INV_X1 u1_u10_u5_U27 (.A( u1_u10_u5_n140 ) , .ZN( u1_u10_u5_n182 ) );
  INV_X1 u1_u10_u5_U28 (.A( u1_u10_u5_n151 ) , .ZN( u1_u10_u5_n183 ) );
  INV_X1 u1_u10_u5_U29 (.A( u1_u10_u5_n123 ) , .ZN( u1_u10_u5_n185 ) );
  NOR2_X1 u1_u10_u5_U3 (.ZN( u1_u10_u5_n134 ) , .A1( u1_u10_u5_n183 ) , .A2( u1_u10_u5_n190 ) );
  INV_X1 u1_u10_u5_U30 (.A( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n184 ) );
  INV_X1 u1_u10_u5_U31 (.A( u1_u10_u5_n139 ) , .ZN( u1_u10_u5_n189 ) );
  INV_X1 u1_u10_u5_U32 (.A( u1_u10_u5_n157 ) , .ZN( u1_u10_u5_n190 ) );
  INV_X1 u1_u10_u5_U33 (.A( u1_u10_u5_n120 ) , .ZN( u1_u10_u5_n193 ) );
  NAND2_X1 u1_u10_u5_U34 (.ZN( u1_u10_u5_n111 ) , .A1( u1_u10_u5_n140 ) , .A2( u1_u10_u5_n155 ) );
  INV_X1 u1_u10_u5_U35 (.A( u1_u10_u5_n117 ) , .ZN( u1_u10_u5_n196 ) );
  OAI221_X1 u1_u10_u5_U36 (.A( u1_u10_u5_n116 ) , .ZN( u1_u10_u5_n117 ) , .B2( u1_u10_u5_n119 ) , .C1( u1_u10_u5_n153 ) , .C2( u1_u10_u5_n158 ) , .B1( u1_u10_u5_n172 ) );
  AOI222_X1 u1_u10_u5_U37 (.ZN( u1_u10_u5_n116 ) , .B2( u1_u10_u5_n145 ) , .C1( u1_u10_u5_n148 ) , .A2( u1_u10_u5_n174 ) , .C2( u1_u10_u5_n177 ) , .B1( u1_u10_u5_n187 ) , .A1( u1_u10_u5_n193 ) );
  INV_X1 u1_u10_u5_U38 (.A( u1_u10_u5_n115 ) , .ZN( u1_u10_u5_n187 ) );
  NOR2_X1 u1_u10_u5_U39 (.ZN( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n170 ) , .A2( u1_u10_u5_n180 ) );
  INV_X1 u1_u10_u5_U4 (.A( u1_u10_u5_n138 ) , .ZN( u1_u10_u5_n191 ) );
  AOI22_X1 u1_u10_u5_U40 (.B2( u1_u10_u5_n131 ) , .A2( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n169 ) , .B1( u1_u10_u5_n174 ) , .A1( u1_u10_u5_n185 ) );
  NOR2_X1 u1_u10_u5_U41 (.A1( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n150 ) , .A2( u1_u10_u5_n173 ) );
  AOI21_X1 u1_u10_u5_U42 (.A( u1_u10_u5_n118 ) , .B2( u1_u10_u5_n145 ) , .ZN( u1_u10_u5_n168 ) , .B1( u1_u10_u5_n186 ) );
  INV_X1 u1_u10_u5_U43 (.A( u1_u10_u5_n122 ) , .ZN( u1_u10_u5_n186 ) );
  NOR2_X1 u1_u10_u5_U44 (.A1( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n152 ) , .A2( u1_u10_u5_n176 ) );
  NOR2_X1 u1_u10_u5_U45 (.A1( u1_u10_u5_n115 ) , .ZN( u1_u10_u5_n118 ) , .A2( u1_u10_u5_n153 ) );
  NOR2_X1 u1_u10_u5_U46 (.A2( u1_u10_u5_n145 ) , .ZN( u1_u10_u5_n156 ) , .A1( u1_u10_u5_n174 ) );
  NOR2_X1 u1_u10_u5_U47 (.ZN( u1_u10_u5_n121 ) , .A2( u1_u10_u5_n145 ) , .A1( u1_u10_u5_n176 ) );
  AOI22_X1 u1_u10_u5_U48 (.ZN( u1_u10_u5_n114 ) , .A2( u1_u10_u5_n137 ) , .A1( u1_u10_u5_n145 ) , .B2( u1_u10_u5_n175 ) , .B1( u1_u10_u5_n193 ) );
  OAI211_X1 u1_u10_u5_U49 (.B( u1_u10_u5_n124 ) , .A( u1_u10_u5_n125 ) , .C2( u1_u10_u5_n126 ) , .C1( u1_u10_u5_n127 ) , .ZN( u1_u10_u5_n128 ) );
  OAI21_X1 u1_u10_u5_U5 (.B2( u1_u10_u5_n136 ) , .B1( u1_u10_u5_n137 ) , .ZN( u1_u10_u5_n138 ) , .A( u1_u10_u5_n177 ) );
  NOR3_X1 u1_u10_u5_U50 (.ZN( u1_u10_u5_n127 ) , .A1( u1_u10_u5_n136 ) , .A3( u1_u10_u5_n148 ) , .A2( u1_u10_u5_n182 ) );
  OAI21_X1 u1_u10_u5_U51 (.ZN( u1_u10_u5_n124 ) , .A( u1_u10_u5_n177 ) , .B2( u1_u10_u5_n183 ) , .B1( u1_u10_u5_n189 ) );
  OAI21_X1 u1_u10_u5_U52 (.ZN( u1_u10_u5_n125 ) , .A( u1_u10_u5_n174 ) , .B2( u1_u10_u5_n185 ) , .B1( u1_u10_u5_n190 ) );
  AOI21_X1 u1_u10_u5_U53 (.A( u1_u10_u5_n153 ) , .B2( u1_u10_u5_n154 ) , .B1( u1_u10_u5_n155 ) , .ZN( u1_u10_u5_n164 ) );
  AOI21_X1 u1_u10_u5_U54 (.ZN( u1_u10_u5_n110 ) , .B1( u1_u10_u5_n122 ) , .B2( u1_u10_u5_n139 ) , .A( u1_u10_u5_n153 ) );
  INV_X1 u1_u10_u5_U55 (.A( u1_u10_u5_n153 ) , .ZN( u1_u10_u5_n176 ) );
  INV_X1 u1_u10_u5_U56 (.A( u1_u10_u5_n126 ) , .ZN( u1_u10_u5_n173 ) );
  AND2_X1 u1_u10_u5_U57 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n147 ) );
  AND2_X1 u1_u10_u5_U58 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n148 ) );
  NAND2_X1 u1_u10_u5_U59 (.A1( u1_u10_u5_n105 ) , .A2( u1_u10_u5_n106 ) , .ZN( u1_u10_u5_n158 ) );
  INV_X1 u1_u10_u5_U6 (.A( u1_u10_u5_n135 ) , .ZN( u1_u10_u5_n178 ) );
  NAND2_X1 u1_u10_u5_U60 (.A2( u1_u10_u5_n108 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n139 ) );
  NAND2_X1 u1_u10_u5_U61 (.A1( u1_u10_u5_n106 ) , .A2( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n119 ) );
  NAND2_X1 u1_u10_u5_U62 (.A2( u1_u10_u5_n103 ) , .A1( u1_u10_u5_n105 ) , .ZN( u1_u10_u5_n140 ) );
  NAND2_X1 u1_u10_u5_U63 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n105 ) , .ZN( u1_u10_u5_n155 ) );
  NAND2_X1 u1_u10_u5_U64 (.A2( u1_u10_u5_n106 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n122 ) );
  NAND2_X1 u1_u10_u5_U65 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n106 ) , .ZN( u1_u10_u5_n115 ) );
  NAND2_X1 u1_u10_u5_U66 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n103 ) , .ZN( u1_u10_u5_n161 ) );
  NAND2_X1 u1_u10_u5_U67 (.A1( u1_u10_u5_n105 ) , .A2( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n154 ) );
  INV_X1 u1_u10_u5_U68 (.A( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n172 ) );
  NAND2_X1 u1_u10_u5_U69 (.A1( u1_u10_u5_n103 ) , .A2( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n123 ) );
  OAI22_X1 u1_u10_u5_U7 (.B2( u1_u10_u5_n149 ) , .B1( u1_u10_u5_n150 ) , .A2( u1_u10_u5_n151 ) , .A1( u1_u10_u5_n152 ) , .ZN( u1_u10_u5_n165 ) );
  NAND2_X1 u1_u10_u5_U70 (.A2( u1_u10_u5_n103 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n151 ) );
  NAND2_X1 u1_u10_u5_U71 (.A2( u1_u10_u5_n107 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n120 ) );
  NAND2_X1 u1_u10_u5_U72 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n157 ) );
  AND2_X1 u1_u10_u5_U73 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n104 ) , .ZN( u1_u10_u5_n131 ) );
  INV_X1 u1_u10_u5_U74 (.A( u1_u10_u5_n102 ) , .ZN( u1_u10_u5_n195 ) );
  OAI221_X1 u1_u10_u5_U75 (.A( u1_u10_u5_n101 ) , .ZN( u1_u10_u5_n102 ) , .C2( u1_u10_u5_n115 ) , .C1( u1_u10_u5_n126 ) , .B1( u1_u10_u5_n134 ) , .B2( u1_u10_u5_n160 ) );
  OAI21_X1 u1_u10_u5_U76 (.ZN( u1_u10_u5_n101 ) , .B1( u1_u10_u5_n137 ) , .A( u1_u10_u5_n146 ) , .B2( u1_u10_u5_n147 ) );
  NOR2_X1 u1_u10_u5_U77 (.A2( u1_u10_X_34 ) , .A1( u1_u10_X_35 ) , .ZN( u1_u10_u5_n145 ) );
  NOR2_X1 u1_u10_u5_U78 (.A2( u1_u10_X_34 ) , .ZN( u1_u10_u5_n146 ) , .A1( u1_u10_u5_n171 ) );
  NOR2_X1 u1_u10_u5_U79 (.A2( u1_u10_X_31 ) , .A1( u1_u10_X_32 ) , .ZN( u1_u10_u5_n103 ) );
  NOR3_X1 u1_u10_u5_U8 (.A2( u1_u10_u5_n147 ) , .A1( u1_u10_u5_n148 ) , .ZN( u1_u10_u5_n149 ) , .A3( u1_u10_u5_n194 ) );
  NOR2_X1 u1_u10_u5_U80 (.A2( u1_u10_X_36 ) , .ZN( u1_u10_u5_n105 ) , .A1( u1_u10_u5_n180 ) );
  NOR2_X1 u1_u10_u5_U81 (.A2( u1_u10_X_33 ) , .ZN( u1_u10_u5_n108 ) , .A1( u1_u10_u5_n170 ) );
  NOR2_X1 u1_u10_u5_U82 (.A2( u1_u10_X_33 ) , .A1( u1_u10_X_36 ) , .ZN( u1_u10_u5_n107 ) );
  NOR2_X1 u1_u10_u5_U83 (.A2( u1_u10_X_31 ) , .ZN( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n181 ) );
  NAND2_X1 u1_u10_u5_U84 (.A2( u1_u10_X_34 ) , .A1( u1_u10_X_35 ) , .ZN( u1_u10_u5_n153 ) );
  NAND2_X1 u1_u10_u5_U85 (.A1( u1_u10_X_34 ) , .ZN( u1_u10_u5_n126 ) , .A2( u1_u10_u5_n171 ) );
  AND2_X1 u1_u10_u5_U86 (.A1( u1_u10_X_31 ) , .A2( u1_u10_X_32 ) , .ZN( u1_u10_u5_n106 ) );
  AND2_X1 u1_u10_u5_U87 (.A1( u1_u10_X_31 ) , .ZN( u1_u10_u5_n109 ) , .A2( u1_u10_u5_n181 ) );
  INV_X1 u1_u10_u5_U88 (.A( u1_u10_X_33 ) , .ZN( u1_u10_u5_n180 ) );
  INV_X1 u1_u10_u5_U89 (.A( u1_u10_X_35 ) , .ZN( u1_u10_u5_n171 ) );
  NOR2_X1 u1_u10_u5_U9 (.ZN( u1_u10_u5_n135 ) , .A1( u1_u10_u5_n173 ) , .A2( u1_u10_u5_n176 ) );
  INV_X1 u1_u10_u5_U90 (.A( u1_u10_X_36 ) , .ZN( u1_u10_u5_n170 ) );
  INV_X1 u1_u10_u5_U91 (.A( u1_u10_X_32 ) , .ZN( u1_u10_u5_n181 ) );
  NAND4_X1 u1_u10_u5_U92 (.ZN( u1_out10_29 ) , .A4( u1_u10_u5_n129 ) , .A3( u1_u10_u5_n130 ) , .A2( u1_u10_u5_n168 ) , .A1( u1_u10_u5_n196 ) );
  AOI221_X1 u1_u10_u5_U93 (.A( u1_u10_u5_n128 ) , .ZN( u1_u10_u5_n129 ) , .C2( u1_u10_u5_n132 ) , .B2( u1_u10_u5_n159 ) , .B1( u1_u10_u5_n176 ) , .C1( u1_u10_u5_n184 ) );
  AOI222_X1 u1_u10_u5_U94 (.ZN( u1_u10_u5_n130 ) , .A2( u1_u10_u5_n146 ) , .B1( u1_u10_u5_n147 ) , .C2( u1_u10_u5_n175 ) , .B2( u1_u10_u5_n179 ) , .A1( u1_u10_u5_n188 ) , .C1( u1_u10_u5_n194 ) );
  NAND4_X1 u1_u10_u5_U95 (.ZN( u1_out10_19 ) , .A4( u1_u10_u5_n166 ) , .A3( u1_u10_u5_n167 ) , .A2( u1_u10_u5_n168 ) , .A1( u1_u10_u5_n169 ) );
  AOI22_X1 u1_u10_u5_U96 (.B2( u1_u10_u5_n145 ) , .A2( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n167 ) , .B1( u1_u10_u5_n182 ) , .A1( u1_u10_u5_n189 ) );
  NOR4_X1 u1_u10_u5_U97 (.A4( u1_u10_u5_n162 ) , .A3( u1_u10_u5_n163 ) , .A2( u1_u10_u5_n164 ) , .A1( u1_u10_u5_n165 ) , .ZN( u1_u10_u5_n166 ) );
  NAND4_X1 u1_u10_u5_U98 (.ZN( u1_out10_11 ) , .A4( u1_u10_u5_n143 ) , .A3( u1_u10_u5_n144 ) , .A2( u1_u10_u5_n169 ) , .A1( u1_u10_u5_n196 ) );
  AOI22_X1 u1_u10_u5_U99 (.A2( u1_u10_u5_n132 ) , .ZN( u1_u10_u5_n144 ) , .B2( u1_u10_u5_n145 ) , .B1( u1_u10_u5_n184 ) , .A1( u1_u10_u5_n194 ) );
  XOR2_X1 u1_u12_U1 (.B( u1_K13_9 ) , .A( u1_R11_6 ) , .Z( u1_u12_X_9 ) );
  XOR2_X1 u1_u12_U16 (.B( u1_K13_3 ) , .A( u1_R11_2 ) , .Z( u1_u12_X_3 ) );
  XOR2_X1 u1_u12_U2 (.B( u1_K13_8 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_8 ) );
  XOR2_X1 u1_u12_U27 (.B( u1_K13_2 ) , .A( u1_R11_1 ) , .Z( u1_u12_X_2 ) );
  XOR2_X1 u1_u12_U3 (.B( u1_K13_7 ) , .A( u1_R11_4 ) , .Z( u1_u12_X_7 ) );
  XOR2_X1 u1_u12_U33 (.B( u1_K13_24 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_24 ) );
  XOR2_X1 u1_u12_U34 (.B( u1_K13_23 ) , .A( u1_R11_16 ) , .Z( u1_u12_X_23 ) );
  XOR2_X1 u1_u12_U35 (.B( u1_K13_22 ) , .A( u1_R11_15 ) , .Z( u1_u12_X_22 ) );
  XOR2_X1 u1_u12_U36 (.B( u1_K13_21 ) , .A( u1_R11_14 ) , .Z( u1_u12_X_21 ) );
  XOR2_X1 u1_u12_U37 (.B( u1_K13_20 ) , .A( u1_R11_13 ) , .Z( u1_u12_X_20 ) );
  XOR2_X1 u1_u12_U38 (.B( u1_K13_1 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_1 ) );
  XOR2_X1 u1_u12_U39 (.B( u1_K13_19 ) , .A( u1_R11_12 ) , .Z( u1_u12_X_19 ) );
  XOR2_X1 u1_u12_U4 (.B( u1_K13_6 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_6 ) );
  XOR2_X1 u1_u12_U46 (.B( u1_K13_12 ) , .A( u1_R11_9 ) , .Z( u1_u12_X_12 ) );
  XOR2_X1 u1_u12_U47 (.B( u1_K13_11 ) , .A( u1_R11_8 ) , .Z( u1_u12_X_11 ) );
  XOR2_X1 u1_u12_U48 (.B( u1_K13_10 ) , .A( u1_R11_7 ) , .Z( u1_u12_X_10 ) );
  XOR2_X1 u1_u12_U5 (.B( u1_K13_5 ) , .A( u1_R11_4 ) , .Z( u1_u12_X_5 ) );
  XOR2_X1 u1_u12_U6 (.B( u1_K13_4 ) , .A( u1_R11_3 ) , .Z( u1_u12_X_4 ) );
  NAND2_X1 u1_u12_u0_U10 (.ZN( u1_u12_u0_n113 ) , .A1( u1_u12_u0_n139 ) , .A2( u1_u12_u0_n149 ) );
  AND3_X1 u1_u12_u0_U11 (.A2( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n127 ) , .A3( u1_u12_u0_n130 ) , .A1( u1_u12_u0_n148 ) );
  AND2_X1 u1_u12_u0_U12 (.ZN( u1_u12_u0_n107 ) , .A1( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n140 ) );
  AND2_X1 u1_u12_u0_U13 (.A2( u1_u12_u0_n129 ) , .A1( u1_u12_u0_n130 ) , .ZN( u1_u12_u0_n151 ) );
  AND2_X1 u1_u12_u0_U14 (.A1( u1_u12_u0_n108 ) , .A2( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n145 ) );
  INV_X1 u1_u12_u0_U15 (.A( u1_u12_u0_n143 ) , .ZN( u1_u12_u0_n173 ) );
  NOR2_X1 u1_u12_u0_U16 (.A2( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n147 ) , .A1( u1_u12_u0_n160 ) );
  AOI21_X1 u1_u12_u0_U17 (.B1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n132 ) , .A( u1_u12_u0_n165 ) , .B2( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U18 (.A( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n165 ) );
  OAI22_X1 u1_u12_u0_U19 (.B1( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n147 ) , .A2( u1_u12_u0_n90 ) , .ZN( u1_u12_u0_n91 ) );
  AND3_X1 u1_u12_u0_U20 (.A3( u1_u12_u0_n121 ) , .A2( u1_u12_u0_n125 ) , .A1( u1_u12_u0_n148 ) , .ZN( u1_u12_u0_n90 ) );
  OAI22_X1 u1_u12_u0_U21 (.B1( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n126 ) , .A1( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n146 ) , .B2( u1_u12_u0_n147 ) );
  INV_X1 u1_u12_u0_U22 (.A( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n161 ) );
  AOI22_X1 u1_u12_u0_U23 (.B2( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n110 ) , .ZN( u1_u12_u0_n111 ) , .B1( u1_u12_u0_n118 ) , .A1( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U24 (.A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U25 (.A2( u1_u12_u0_n102 ) , .A1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n149 ) );
  INV_X1 u1_u12_u0_U26 (.A( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n158 ) );
  NAND2_X1 u1_u12_u0_U27 (.A2( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U28 (.ZN( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n92 ) , .A2( u1_u12_u0_n94 ) );
  AOI21_X1 u1_u12_u0_U29 (.ZN( u1_u12_u0_n104 ) , .B1( u1_u12_u0_n107 ) , .B2( u1_u12_u0_n141 ) , .A( u1_u12_u0_n144 ) );
  INV_X1 u1_u12_u0_U3 (.A( u1_u12_u0_n113 ) , .ZN( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U30 (.ZN( u1_u12_u0_n116 ) , .B2( u1_u12_u0_n142 ) , .A( u1_u12_u0_n144 ) , .B1( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U31 (.B1( u1_u12_u0_n127 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n96 ) );
  NAND2_X1 u1_u12_u0_U32 (.A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n114 ) , .A1( u1_u12_u0_n92 ) );
  NOR2_X1 u1_u12_u0_U33 (.A1( u1_u12_u0_n120 ) , .ZN( u1_u12_u0_n143 ) , .A2( u1_u12_u0_n167 ) );
  OAI221_X1 u1_u12_u0_U34 (.C1( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n120 ) , .B1( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n141 ) , .C2( u1_u12_u0_n147 ) , .A( u1_u12_u0_n172 ) );
  AOI211_X1 u1_u12_u0_U35 (.B( u1_u12_u0_n115 ) , .A( u1_u12_u0_n116 ) , .C2( u1_u12_u0_n117 ) , .C1( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n119 ) );
  NAND2_X1 u1_u12_u0_U36 (.A1( u1_u12_u0_n100 ) , .A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n125 ) );
  NAND2_X1 u1_u12_u0_U37 (.A1( u1_u12_u0_n101 ) , .A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n150 ) );
  INV_X1 u1_u12_u0_U38 (.A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U39 (.A2( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n139 ) );
  AOI21_X1 u1_u12_u0_U4 (.B1( u1_u12_u0_n114 ) , .ZN( u1_u12_u0_n115 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U40 (.A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U41 (.ZN( u1_u12_u0_n112 ) , .A2( u1_u12_u0_n92 ) , .A1( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U42 (.ZN( u1_u12_u0_n172 ) , .A( u1_u12_u0_n88 ) );
  OAI222_X1 u1_u12_u0_U43 (.C1( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n125 ) , .B2( u1_u12_u0_n128 ) , .B1( u1_u12_u0_n144 ) , .A2( u1_u12_u0_n158 ) , .C2( u1_u12_u0_n161 ) , .ZN( u1_u12_u0_n88 ) );
  NAND2_X1 u1_u12_u0_U44 (.A2( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n121 ) , .A1( u1_u12_u0_n93 ) );
  OR3_X1 u1_u12_u0_U45 (.A3( u1_u12_u0_n152 ) , .A2( u1_u12_u0_n153 ) , .A1( u1_u12_u0_n154 ) , .ZN( u1_u12_u0_n155 ) );
  AOI21_X1 u1_u12_u0_U46 (.B2( u1_u12_u0_n150 ) , .B1( u1_u12_u0_n151 ) , .ZN( u1_u12_u0_n152 ) , .A( u1_u12_u0_n158 ) );
  AOI21_X1 u1_u12_u0_U47 (.A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n145 ) , .B1( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n154 ) );
  AOI21_X1 u1_u12_u0_U48 (.A( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n148 ) , .B1( u1_u12_u0_n149 ) , .ZN( u1_u12_u0_n153 ) );
  INV_X1 u1_u12_u0_U49 (.ZN( u1_u12_u0_n171 ) , .A( u1_u12_u0_n99 ) );
  AOI21_X1 u1_u12_u0_U5 (.B2( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n134 ) , .B1( u1_u12_u0_n151 ) , .A( u1_u12_u0_n158 ) );
  OAI211_X1 u1_u12_u0_U50 (.C2( u1_u12_u0_n140 ) , .C1( u1_u12_u0_n161 ) , .A( u1_u12_u0_n169 ) , .B( u1_u12_u0_n98 ) , .ZN( u1_u12_u0_n99 ) );
  INV_X1 u1_u12_u0_U51 (.ZN( u1_u12_u0_n169 ) , .A( u1_u12_u0_n91 ) );
  AOI211_X1 u1_u12_u0_U52 (.C1( u1_u12_u0_n118 ) , .A( u1_u12_u0_n123 ) , .B( u1_u12_u0_n96 ) , .C2( u1_u12_u0_n97 ) , .ZN( u1_u12_u0_n98 ) );
  NOR2_X1 u1_u12_u0_U53 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n118 ) );
  NOR2_X1 u1_u12_u0_U54 (.A2( u1_u12_X_1 ) , .ZN( u1_u12_u0_n101 ) , .A1( u1_u12_u0_n163 ) );
  NOR2_X1 u1_u12_u0_U55 (.A2( u1_u12_X_6 ) , .ZN( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n162 ) );
  NAND2_X1 u1_u12_u0_U56 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n144 ) );
  NOR2_X1 u1_u12_u0_U57 (.A2( u1_u12_X_5 ) , .ZN( u1_u12_u0_n136 ) , .A1( u1_u12_u0_n159 ) );
  NAND2_X1 u1_u12_u0_U58 (.A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n159 ) );
  AND2_X1 u1_u12_u0_U59 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n102 ) );
  NOR2_X1 u1_u12_u0_U6 (.A1( u1_u12_u0_n108 ) , .ZN( u1_u12_u0_n123 ) , .A2( u1_u12_u0_n158 ) );
  AND2_X1 u1_u12_u0_U60 (.A1( u1_u12_X_6 ) , .A2( u1_u12_u0_n162 ) , .ZN( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U61 (.A( u1_u12_X_4 ) , .ZN( u1_u12_u0_n159 ) );
  INV_X1 u1_u12_u0_U62 (.A( u1_u12_X_1 ) , .ZN( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U63 (.A( u1_u12_X_3 ) , .ZN( u1_u12_u0_n162 ) );
  OR4_X1 u1_u12_u0_U64 (.ZN( u1_out12_17 ) , .A4( u1_u12_u0_n122 ) , .A2( u1_u12_u0_n123 ) , .A1( u1_u12_u0_n124 ) , .A3( u1_u12_u0_n170 ) );
  AOI21_X1 u1_u12_u0_U65 (.B2( u1_u12_u0_n107 ) , .ZN( u1_u12_u0_n124 ) , .B1( u1_u12_u0_n128 ) , .A( u1_u12_u0_n161 ) );
  INV_X1 u1_u12_u0_U66 (.A( u1_u12_u0_n111 ) , .ZN( u1_u12_u0_n170 ) );
  OR4_X1 u1_u12_u0_U67 (.ZN( u1_out12_31 ) , .A4( u1_u12_u0_n155 ) , .A2( u1_u12_u0_n156 ) , .A1( u1_u12_u0_n157 ) , .A3( u1_u12_u0_n173 ) );
  AOI21_X1 u1_u12_u0_U68 (.A( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n139 ) , .B1( u1_u12_u0_n140 ) , .ZN( u1_u12_u0_n157 ) );
  AOI21_X1 u1_u12_u0_U69 (.B2( u1_u12_u0_n141 ) , .B1( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n156 ) , .A( u1_u12_u0_n161 ) );
  OAI21_X1 u1_u12_u0_U7 (.B1( u1_u12_u0_n150 ) , .B2( u1_u12_u0_n158 ) , .A( u1_u12_u0_n172 ) , .ZN( u1_u12_u0_n89 ) );
  INV_X1 u1_u12_u0_U70 (.ZN( u1_u12_u0_n174 ) , .A( u1_u12_u0_n89 ) );
  AOI211_X1 u1_u12_u0_U71 (.B( u1_u12_u0_n104 ) , .A( u1_u12_u0_n105 ) , .ZN( u1_u12_u0_n106 ) , .C2( u1_u12_u0_n113 ) , .C1( u1_u12_u0_n160 ) );
  INV_X1 u1_u12_u0_U72 (.A( u1_u12_u0_n126 ) , .ZN( u1_u12_u0_n168 ) );
  AOI211_X1 u1_u12_u0_U73 (.B( u1_u12_u0_n133 ) , .A( u1_u12_u0_n134 ) , .C2( u1_u12_u0_n135 ) , .C1( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n137 ) );
  NOR2_X1 u1_u12_u0_U74 (.A1( u1_u12_u0_n163 ) , .A2( u1_u12_u0_n164 ) , .ZN( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U75 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n94 ) );
  OAI221_X1 u1_u12_u0_U76 (.C1( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n122 ) , .B2( u1_u12_u0_n127 ) , .A( u1_u12_u0_n143 ) , .B1( u1_u12_u0_n144 ) , .C2( u1_u12_u0_n147 ) );
  AOI21_X1 u1_u12_u0_U77 (.B1( u1_u12_u0_n132 ) , .ZN( u1_u12_u0_n133 ) , .A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n166 ) );
  OAI22_X1 u1_u12_u0_U78 (.ZN( u1_u12_u0_n105 ) , .A2( u1_u12_u0_n132 ) , .B1( u1_u12_u0_n146 ) , .A1( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U79 (.ZN( u1_u12_u0_n110 ) , .A2( u1_u12_u0_n132 ) , .A1( u1_u12_u0_n145 ) );
  AND2_X1 u1_u12_u0_U8 (.A1( u1_u12_u0_n114 ) , .A2( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n146 ) );
  INV_X1 u1_u12_u0_U80 (.A( u1_u12_u0_n119 ) , .ZN( u1_u12_u0_n167 ) );
  NAND2_X1 u1_u12_u0_U81 (.ZN( u1_u12_u0_n148 ) , .A1( u1_u12_u0_n93 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U82 (.A1( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n129 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U83 (.A1( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n128 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U84 (.A2( u1_u12_X_1 ) , .A1( u1_u12_X_2 ) , .ZN( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U85 (.ZN( u1_u12_u0_n142 ) , .A1( u1_u12_u0_n94 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U86 (.A2( u1_u12_X_2 ) , .ZN( u1_u12_u0_n103 ) , .A1( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U87 (.A( u1_u12_X_2 ) , .ZN( u1_u12_u0_n163 ) );
  NAND3_X1 u1_u12_u0_U88 (.ZN( u1_out12_23 ) , .A3( u1_u12_u0_n137 ) , .A1( u1_u12_u0_n168 ) , .A2( u1_u12_u0_n171 ) );
  NAND3_X1 u1_u12_u0_U89 (.A3( u1_u12_u0_n127 ) , .A2( u1_u12_u0_n128 ) , .ZN( u1_u12_u0_n135 ) , .A1( u1_u12_u0_n150 ) );
  AND2_X1 u1_u12_u0_U9 (.A1( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n141 ) , .A2( u1_u12_u0_n150 ) );
  NAND3_X1 u1_u12_u0_U90 (.ZN( u1_u12_u0_n117 ) , .A3( u1_u12_u0_n132 ) , .A2( u1_u12_u0_n139 ) , .A1( u1_u12_u0_n148 ) );
  NAND3_X1 u1_u12_u0_U91 (.ZN( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n114 ) , .A3( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n149 ) );
  NAND3_X1 u1_u12_u0_U92 (.ZN( u1_out12_9 ) , .A3( u1_u12_u0_n106 ) , .A2( u1_u12_u0_n171 ) , .A1( u1_u12_u0_n174 ) );
  NAND3_X1 u1_u12_u0_U93 (.A2( u1_u12_u0_n128 ) , .A1( u1_u12_u0_n132 ) , .A3( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n97 ) );
  NOR2_X1 u1_u12_u1_U10 (.A1( u1_u12_u1_n112 ) , .A2( u1_u12_u1_n116 ) , .ZN( u1_u12_u1_n118 ) );
  NAND3_X1 u1_u12_u1_U100 (.ZN( u1_u12_u1_n113 ) , .A1( u1_u12_u1_n120 ) , .A3( u1_u12_u1_n133 ) , .A2( u1_u12_u1_n155 ) );
  OAI21_X1 u1_u12_u1_U11 (.ZN( u1_u12_u1_n101 ) , .B1( u1_u12_u1_n141 ) , .A( u1_u12_u1_n146 ) , .B2( u1_u12_u1_n183 ) );
  AOI21_X1 u1_u12_u1_U12 (.B2( u1_u12_u1_n155 ) , .B1( u1_u12_u1_n156 ) , .ZN( u1_u12_u1_n157 ) , .A( u1_u12_u1_n174 ) );
  NAND2_X1 u1_u12_u1_U13 (.ZN( u1_u12_u1_n140 ) , .A2( u1_u12_u1_n150 ) , .A1( u1_u12_u1_n155 ) );
  NAND2_X1 u1_u12_u1_U14 (.A1( u1_u12_u1_n131 ) , .ZN( u1_u12_u1_n147 ) , .A2( u1_u12_u1_n153 ) );
  INV_X1 u1_u12_u1_U15 (.A( u1_u12_u1_n139 ) , .ZN( u1_u12_u1_n174 ) );
  OR4_X1 u1_u12_u1_U16 (.A4( u1_u12_u1_n106 ) , .A3( u1_u12_u1_n107 ) , .ZN( u1_u12_u1_n108 ) , .A1( u1_u12_u1_n117 ) , .A2( u1_u12_u1_n184 ) );
  AOI21_X1 u1_u12_u1_U17 (.ZN( u1_u12_u1_n106 ) , .A( u1_u12_u1_n112 ) , .B1( u1_u12_u1_n154 ) , .B2( u1_u12_u1_n156 ) );
  INV_X1 u1_u12_u1_U18 (.A( u1_u12_u1_n101 ) , .ZN( u1_u12_u1_n184 ) );
  AOI21_X1 u1_u12_u1_U19 (.ZN( u1_u12_u1_n107 ) , .B1( u1_u12_u1_n134 ) , .B2( u1_u12_u1_n149 ) , .A( u1_u12_u1_n174 ) );
  INV_X1 u1_u12_u1_U20 (.A( u1_u12_u1_n112 ) , .ZN( u1_u12_u1_n171 ) );
  NAND2_X1 u1_u12_u1_U21 (.ZN( u1_u12_u1_n141 ) , .A1( u1_u12_u1_n153 ) , .A2( u1_u12_u1_n156 ) );
  AND2_X1 u1_u12_u1_U22 (.A1( u1_u12_u1_n123 ) , .ZN( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n161 ) );
  NAND2_X1 u1_u12_u1_U23 (.A2( u1_u12_u1_n115 ) , .A1( u1_u12_u1_n116 ) , .ZN( u1_u12_u1_n148 ) );
  NAND2_X1 u1_u12_u1_U24 (.A2( u1_u12_u1_n133 ) , .A1( u1_u12_u1_n135 ) , .ZN( u1_u12_u1_n159 ) );
  NAND2_X1 u1_u12_u1_U25 (.A2( u1_u12_u1_n115 ) , .A1( u1_u12_u1_n120 ) , .ZN( u1_u12_u1_n132 ) );
  INV_X1 u1_u12_u1_U26 (.A( u1_u12_u1_n154 ) , .ZN( u1_u12_u1_n178 ) );
  INV_X1 u1_u12_u1_U27 (.A( u1_u12_u1_n151 ) , .ZN( u1_u12_u1_n183 ) );
  AND2_X1 u1_u12_u1_U28 (.A1( u1_u12_u1_n129 ) , .A2( u1_u12_u1_n133 ) , .ZN( u1_u12_u1_n149 ) );
  INV_X1 u1_u12_u1_U29 (.A( u1_u12_u1_n131 ) , .ZN( u1_u12_u1_n180 ) );
  INV_X1 u1_u12_u1_U3 (.A( u1_u12_u1_n159 ) , .ZN( u1_u12_u1_n182 ) );
  AOI221_X1 u1_u12_u1_U30 (.B1( u1_u12_u1_n140 ) , .ZN( u1_u12_u1_n167 ) , .B2( u1_u12_u1_n172 ) , .C2( u1_u12_u1_n175 ) , .C1( u1_u12_u1_n178 ) , .A( u1_u12_u1_n188 ) );
  INV_X1 u1_u12_u1_U31 (.ZN( u1_u12_u1_n188 ) , .A( u1_u12_u1_n97 ) );
  AOI211_X1 u1_u12_u1_U32 (.A( u1_u12_u1_n118 ) , .C1( u1_u12_u1_n132 ) , .C2( u1_u12_u1_n139 ) , .B( u1_u12_u1_n96 ) , .ZN( u1_u12_u1_n97 ) );
  AOI21_X1 u1_u12_u1_U33 (.B2( u1_u12_u1_n121 ) , .B1( u1_u12_u1_n135 ) , .A( u1_u12_u1_n152 ) , .ZN( u1_u12_u1_n96 ) );
  OAI221_X1 u1_u12_u1_U34 (.A( u1_u12_u1_n119 ) , .C2( u1_u12_u1_n129 ) , .ZN( u1_u12_u1_n138 ) , .B2( u1_u12_u1_n152 ) , .C1( u1_u12_u1_n174 ) , .B1( u1_u12_u1_n187 ) );
  INV_X1 u1_u12_u1_U35 (.A( u1_u12_u1_n148 ) , .ZN( u1_u12_u1_n187 ) );
  AOI211_X1 u1_u12_u1_U36 (.B( u1_u12_u1_n117 ) , .A( u1_u12_u1_n118 ) , .ZN( u1_u12_u1_n119 ) , .C2( u1_u12_u1_n146 ) , .C1( u1_u12_u1_n159 ) );
  NOR2_X1 u1_u12_u1_U37 (.A1( u1_u12_u1_n168 ) , .A2( u1_u12_u1_n176 ) , .ZN( u1_u12_u1_n98 ) );
  AOI211_X1 u1_u12_u1_U38 (.B( u1_u12_u1_n162 ) , .A( u1_u12_u1_n163 ) , .C2( u1_u12_u1_n164 ) , .ZN( u1_u12_u1_n165 ) , .C1( u1_u12_u1_n171 ) );
  AOI21_X1 u1_u12_u1_U39 (.A( u1_u12_u1_n160 ) , .B2( u1_u12_u1_n161 ) , .ZN( u1_u12_u1_n162 ) , .B1( u1_u12_u1_n182 ) );
  AOI221_X1 u1_u12_u1_U4 (.A( u1_u12_u1_n138 ) , .C2( u1_u12_u1_n139 ) , .C1( u1_u12_u1_n140 ) , .B2( u1_u12_u1_n141 ) , .ZN( u1_u12_u1_n142 ) , .B1( u1_u12_u1_n175 ) );
  OR2_X1 u1_u12_u1_U40 (.A2( u1_u12_u1_n157 ) , .A1( u1_u12_u1_n158 ) , .ZN( u1_u12_u1_n163 ) );
  NAND2_X1 u1_u12_u1_U41 (.A1( u1_u12_u1_n128 ) , .ZN( u1_u12_u1_n146 ) , .A2( u1_u12_u1_n160 ) );
  NAND2_X1 u1_u12_u1_U42 (.A2( u1_u12_u1_n112 ) , .ZN( u1_u12_u1_n139 ) , .A1( u1_u12_u1_n152 ) );
  NAND2_X1 u1_u12_u1_U43 (.A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n156 ) , .A2( u1_u12_u1_n99 ) );
  NOR2_X1 u1_u12_u1_U44 (.ZN( u1_u12_u1_n117 ) , .A1( u1_u12_u1_n121 ) , .A2( u1_u12_u1_n160 ) );
  OAI21_X1 u1_u12_u1_U45 (.B2( u1_u12_u1_n123 ) , .ZN( u1_u12_u1_n145 ) , .B1( u1_u12_u1_n160 ) , .A( u1_u12_u1_n185 ) );
  INV_X1 u1_u12_u1_U46 (.A( u1_u12_u1_n122 ) , .ZN( u1_u12_u1_n185 ) );
  AOI21_X1 u1_u12_u1_U47 (.B2( u1_u12_u1_n120 ) , .B1( u1_u12_u1_n121 ) , .ZN( u1_u12_u1_n122 ) , .A( u1_u12_u1_n128 ) );
  AOI21_X1 u1_u12_u1_U48 (.A( u1_u12_u1_n128 ) , .B2( u1_u12_u1_n129 ) , .ZN( u1_u12_u1_n130 ) , .B1( u1_u12_u1_n150 ) );
  NAND2_X1 u1_u12_u1_U49 (.ZN( u1_u12_u1_n112 ) , .A1( u1_u12_u1_n169 ) , .A2( u1_u12_u1_n170 ) );
  AOI211_X1 u1_u12_u1_U5 (.ZN( u1_u12_u1_n124 ) , .A( u1_u12_u1_n138 ) , .C2( u1_u12_u1_n139 ) , .B( u1_u12_u1_n145 ) , .C1( u1_u12_u1_n147 ) );
  NAND2_X1 u1_u12_u1_U50 (.ZN( u1_u12_u1_n129 ) , .A2( u1_u12_u1_n95 ) , .A1( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U51 (.A1( u1_u12_u1_n102 ) , .ZN( u1_u12_u1_n154 ) , .A2( u1_u12_u1_n99 ) );
  NAND2_X1 u1_u12_u1_U52 (.A2( u1_u12_u1_n100 ) , .ZN( u1_u12_u1_n135 ) , .A1( u1_u12_u1_n99 ) );
  AOI21_X1 u1_u12_u1_U53 (.A( u1_u12_u1_n152 ) , .B2( u1_u12_u1_n153 ) , .B1( u1_u12_u1_n154 ) , .ZN( u1_u12_u1_n158 ) );
  INV_X1 u1_u12_u1_U54 (.A( u1_u12_u1_n160 ) , .ZN( u1_u12_u1_n175 ) );
  NAND2_X1 u1_u12_u1_U55 (.A1( u1_u12_u1_n100 ) , .ZN( u1_u12_u1_n116 ) , .A2( u1_u12_u1_n95 ) );
  NAND2_X1 u1_u12_u1_U56 (.A1( u1_u12_u1_n102 ) , .ZN( u1_u12_u1_n131 ) , .A2( u1_u12_u1_n95 ) );
  NAND2_X1 u1_u12_u1_U57 (.A2( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n121 ) , .A1( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U58 (.A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n153 ) , .A2( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U59 (.A2( u1_u12_u1_n104 ) , .A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n133 ) );
  AOI22_X1 u1_u12_u1_U6 (.B2( u1_u12_u1_n113 ) , .A2( u1_u12_u1_n114 ) , .ZN( u1_u12_u1_n125 ) , .A1( u1_u12_u1_n171 ) , .B1( u1_u12_u1_n173 ) );
  NAND2_X1 u1_u12_u1_U60 (.ZN( u1_u12_u1_n150 ) , .A2( u1_u12_u1_n98 ) , .A1( u1_u12_u1_n99 ) );
  NAND2_X1 u1_u12_u1_U61 (.A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n155 ) , .A2( u1_u12_u1_n95 ) );
  OAI21_X1 u1_u12_u1_U62 (.ZN( u1_u12_u1_n109 ) , .B1( u1_u12_u1_n129 ) , .B2( u1_u12_u1_n160 ) , .A( u1_u12_u1_n167 ) );
  NAND2_X1 u1_u12_u1_U63 (.A2( u1_u12_u1_n100 ) , .A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n120 ) );
  NAND2_X1 u1_u12_u1_U64 (.A1( u1_u12_u1_n102 ) , .A2( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n115 ) );
  NAND2_X1 u1_u12_u1_U65 (.A2( u1_u12_u1_n100 ) , .A1( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n151 ) );
  NAND2_X1 u1_u12_u1_U66 (.A2( u1_u12_u1_n103 ) , .A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n161 ) );
  INV_X1 u1_u12_u1_U67 (.A( u1_u12_u1_n152 ) , .ZN( u1_u12_u1_n173 ) );
  INV_X1 u1_u12_u1_U68 (.A( u1_u12_u1_n128 ) , .ZN( u1_u12_u1_n172 ) );
  NAND2_X1 u1_u12_u1_U69 (.A2( u1_u12_u1_n102 ) , .A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n123 ) );
  NAND2_X1 u1_u12_u1_U7 (.ZN( u1_u12_u1_n114 ) , .A1( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n156 ) );
  NOR2_X1 u1_u12_u1_U70 (.A2( u1_u12_X_7 ) , .A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n95 ) );
  NOR2_X1 u1_u12_u1_U71 (.A1( u1_u12_X_12 ) , .A2( u1_u12_X_9 ) , .ZN( u1_u12_u1_n100 ) );
  NOR2_X1 u1_u12_u1_U72 (.A2( u1_u12_X_8 ) , .A1( u1_u12_u1_n177 ) , .ZN( u1_u12_u1_n99 ) );
  NOR2_X1 u1_u12_u1_U73 (.A2( u1_u12_X_12 ) , .ZN( u1_u12_u1_n102 ) , .A1( u1_u12_u1_n176 ) );
  NOR2_X1 u1_u12_u1_U74 (.A2( u1_u12_X_9 ) , .ZN( u1_u12_u1_n105 ) , .A1( u1_u12_u1_n168 ) );
  NAND2_X1 u1_u12_u1_U75 (.A1( u1_u12_X_10 ) , .ZN( u1_u12_u1_n160 ) , .A2( u1_u12_u1_n169 ) );
  NAND2_X1 u1_u12_u1_U76 (.A2( u1_u12_X_10 ) , .A1( u1_u12_X_11 ) , .ZN( u1_u12_u1_n152 ) );
  NAND2_X1 u1_u12_u1_U77 (.A1( u1_u12_X_11 ) , .ZN( u1_u12_u1_n128 ) , .A2( u1_u12_u1_n170 ) );
  AND2_X1 u1_u12_u1_U78 (.A2( u1_u12_X_7 ) , .A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n104 ) );
  AND2_X1 u1_u12_u1_U79 (.A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n103 ) , .A2( u1_u12_u1_n177 ) );
  AOI22_X1 u1_u12_u1_U8 (.B2( u1_u12_u1_n136 ) , .A2( u1_u12_u1_n137 ) , .ZN( u1_u12_u1_n143 ) , .A1( u1_u12_u1_n171 ) , .B1( u1_u12_u1_n173 ) );
  INV_X1 u1_u12_u1_U80 (.A( u1_u12_X_10 ) , .ZN( u1_u12_u1_n170 ) );
  INV_X1 u1_u12_u1_U81 (.A( u1_u12_X_9 ) , .ZN( u1_u12_u1_n176 ) );
  INV_X1 u1_u12_u1_U82 (.A( u1_u12_X_11 ) , .ZN( u1_u12_u1_n169 ) );
  INV_X1 u1_u12_u1_U83 (.A( u1_u12_X_12 ) , .ZN( u1_u12_u1_n168 ) );
  INV_X1 u1_u12_u1_U84 (.A( u1_u12_X_7 ) , .ZN( u1_u12_u1_n177 ) );
  NAND4_X1 u1_u12_u1_U85 (.ZN( u1_out12_28 ) , .A4( u1_u12_u1_n124 ) , .A3( u1_u12_u1_n125 ) , .A2( u1_u12_u1_n126 ) , .A1( u1_u12_u1_n127 ) );
  OAI21_X1 u1_u12_u1_U86 (.ZN( u1_u12_u1_n127 ) , .B2( u1_u12_u1_n139 ) , .B1( u1_u12_u1_n175 ) , .A( u1_u12_u1_n183 ) );
  OAI21_X1 u1_u12_u1_U87 (.ZN( u1_u12_u1_n126 ) , .B2( u1_u12_u1_n140 ) , .A( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n178 ) );
  NAND4_X1 u1_u12_u1_U88 (.ZN( u1_out12_18 ) , .A4( u1_u12_u1_n165 ) , .A3( u1_u12_u1_n166 ) , .A1( u1_u12_u1_n167 ) , .A2( u1_u12_u1_n186 ) );
  AOI22_X1 u1_u12_u1_U89 (.B2( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n147 ) , .A2( u1_u12_u1_n148 ) , .ZN( u1_u12_u1_n166 ) , .A1( u1_u12_u1_n172 ) );
  INV_X1 u1_u12_u1_U9 (.A( u1_u12_u1_n147 ) , .ZN( u1_u12_u1_n181 ) );
  INV_X1 u1_u12_u1_U90 (.A( u1_u12_u1_n145 ) , .ZN( u1_u12_u1_n186 ) );
  NAND4_X1 u1_u12_u1_U91 (.ZN( u1_out12_2 ) , .A4( u1_u12_u1_n142 ) , .A3( u1_u12_u1_n143 ) , .A2( u1_u12_u1_n144 ) , .A1( u1_u12_u1_n179 ) );
  OAI21_X1 u1_u12_u1_U92 (.B2( u1_u12_u1_n132 ) , .ZN( u1_u12_u1_n144 ) , .A( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n180 ) );
  INV_X1 u1_u12_u1_U93 (.A( u1_u12_u1_n130 ) , .ZN( u1_u12_u1_n179 ) );
  OR4_X1 u1_u12_u1_U94 (.ZN( u1_out12_13 ) , .A4( u1_u12_u1_n108 ) , .A3( u1_u12_u1_n109 ) , .A2( u1_u12_u1_n110 ) , .A1( u1_u12_u1_n111 ) );
  AOI21_X1 u1_u12_u1_U95 (.ZN( u1_u12_u1_n111 ) , .A( u1_u12_u1_n128 ) , .B2( u1_u12_u1_n131 ) , .B1( u1_u12_u1_n135 ) );
  AOI21_X1 u1_u12_u1_U96 (.ZN( u1_u12_u1_n110 ) , .A( u1_u12_u1_n116 ) , .B1( u1_u12_u1_n152 ) , .B2( u1_u12_u1_n160 ) );
  NAND3_X1 u1_u12_u1_U97 (.A3( u1_u12_u1_n149 ) , .A2( u1_u12_u1_n150 ) , .A1( u1_u12_u1_n151 ) , .ZN( u1_u12_u1_n164 ) );
  NAND3_X1 u1_u12_u1_U98 (.A3( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n135 ) , .ZN( u1_u12_u1_n136 ) , .A1( u1_u12_u1_n151 ) );
  NAND3_X1 u1_u12_u1_U99 (.A1( u1_u12_u1_n133 ) , .ZN( u1_u12_u1_n137 ) , .A2( u1_u12_u1_n154 ) , .A3( u1_u12_u1_n181 ) );
  OAI22_X1 u1_u12_u3_U10 (.B1( u1_u12_u3_n113 ) , .A2( u1_u12_u3_n135 ) , .A1( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n164 ) , .ZN( u1_u12_u3_n98 ) );
  OAI211_X1 u1_u12_u3_U11 (.B( u1_u12_u3_n106 ) , .ZN( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n128 ) , .C1( u1_u12_u3_n167 ) , .A( u1_u12_u3_n181 ) );
  AOI221_X1 u1_u12_u3_U12 (.C1( u1_u12_u3_n105 ) , .ZN( u1_u12_u3_n106 ) , .A( u1_u12_u3_n131 ) , .B2( u1_u12_u3_n132 ) , .C2( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n169 ) );
  INV_X1 u1_u12_u3_U13 (.ZN( u1_u12_u3_n181 ) , .A( u1_u12_u3_n98 ) );
  NAND2_X1 u1_u12_u3_U14 (.ZN( u1_u12_u3_n105 ) , .A2( u1_u12_u3_n130 ) , .A1( u1_u12_u3_n155 ) );
  AOI22_X1 u1_u12_u3_U15 (.B1( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n116 ) , .ZN( u1_u12_u3_n123 ) , .B2( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U16 (.ZN( u1_u12_u3_n116 ) , .A2( u1_u12_u3_n151 ) , .A1( u1_u12_u3_n182 ) );
  NOR2_X1 u1_u12_u3_U17 (.ZN( u1_u12_u3_n126 ) , .A2( u1_u12_u3_n150 ) , .A1( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U18 (.ZN( u1_u12_u3_n112 ) , .B2( u1_u12_u3_n146 ) , .B1( u1_u12_u3_n155 ) , .A( u1_u12_u3_n167 ) );
  NAND2_X1 u1_u12_u3_U19 (.A1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n142 ) , .A2( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U20 (.ZN( u1_u12_u3_n132 ) , .A2( u1_u12_u3_n152 ) , .A1( u1_u12_u3_n156 ) );
  AND2_X1 u1_u12_u3_U21 (.A2( u1_u12_u3_n113 ) , .A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n151 ) );
  INV_X1 u1_u12_u3_U22 (.A( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n165 ) );
  INV_X1 u1_u12_u3_U23 (.A( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n170 ) );
  NAND2_X1 u1_u12_u3_U24 (.A1( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .ZN( u1_u12_u3_n140 ) );
  NAND2_X1 u1_u12_u3_U25 (.ZN( u1_u12_u3_n117 ) , .A1( u1_u12_u3_n124 ) , .A2( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U26 (.ZN( u1_u12_u3_n143 ) , .A1( u1_u12_u3_n165 ) , .A2( u1_u12_u3_n167 ) );
  INV_X1 u1_u12_u3_U27 (.A( u1_u12_u3_n130 ) , .ZN( u1_u12_u3_n177 ) );
  INV_X1 u1_u12_u3_U28 (.A( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n176 ) );
  INV_X1 u1_u12_u3_U29 (.A( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n174 ) );
  INV_X1 u1_u12_u3_U3 (.A( u1_u12_u3_n129 ) , .ZN( u1_u12_u3_n183 ) );
  INV_X1 u1_u12_u3_U30 (.A( u1_u12_u3_n139 ) , .ZN( u1_u12_u3_n185 ) );
  NOR2_X1 u1_u12_u3_U31 (.ZN( u1_u12_u3_n135 ) , .A2( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n169 ) );
  OAI222_X1 u1_u12_u3_U32 (.C2( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .B1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n138 ) , .B2( u1_u12_u3_n146 ) , .C1( u1_u12_u3_n154 ) , .A1( u1_u12_u3_n164 ) );
  NOR4_X1 u1_u12_u3_U33 (.A4( u1_u12_u3_n157 ) , .A3( u1_u12_u3_n158 ) , .A2( u1_u12_u3_n159 ) , .A1( u1_u12_u3_n160 ) , .ZN( u1_u12_u3_n161 ) );
  AOI21_X1 u1_u12_u3_U34 (.B2( u1_u12_u3_n152 ) , .B1( u1_u12_u3_n153 ) , .ZN( u1_u12_u3_n158 ) , .A( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U35 (.A( u1_u12_u3_n154 ) , .B2( u1_u12_u3_n155 ) , .B1( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n157 ) );
  AOI21_X1 u1_u12_u3_U36 (.A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n150 ) , .B1( u1_u12_u3_n151 ) , .ZN( u1_u12_u3_n159 ) );
  AOI211_X1 u1_u12_u3_U37 (.ZN( u1_u12_u3_n109 ) , .A( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n129 ) , .B( u1_u12_u3_n138 ) , .C1( u1_u12_u3_n141 ) );
  AOI211_X1 u1_u12_u3_U38 (.B( u1_u12_u3_n119 ) , .A( u1_u12_u3_n120 ) , .C2( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n122 ) , .C1( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U39 (.A( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U4 (.A( u1_u12_u3_n140 ) , .ZN( u1_u12_u3_n182 ) );
  OAI22_X1 u1_u12_u3_U40 (.B1( u1_u12_u3_n118 ) , .ZN( u1_u12_u3_n120 ) , .A1( u1_u12_u3_n135 ) , .B2( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n178 ) );
  AND3_X1 u1_u12_u3_U41 (.ZN( u1_u12_u3_n118 ) , .A2( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n144 ) , .A3( u1_u12_u3_n152 ) );
  INV_X1 u1_u12_u3_U42 (.A( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U43 (.ZN( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n164 ) );
  OAI211_X1 u1_u12_u3_U44 (.B( u1_u12_u3_n127 ) , .ZN( u1_u12_u3_n139 ) , .C1( u1_u12_u3_n150 ) , .C2( u1_u12_u3_n154 ) , .A( u1_u12_u3_n184 ) );
  INV_X1 u1_u12_u3_U45 (.A( u1_u12_u3_n125 ) , .ZN( u1_u12_u3_n184 ) );
  AOI221_X1 u1_u12_u3_U46 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n127 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n169 ) , .B2( u1_u12_u3_n170 ) , .B1( u1_u12_u3_n174 ) );
  OAI22_X1 u1_u12_u3_U47 (.A1( u1_u12_u3_n124 ) , .ZN( u1_u12_u3_n125 ) , .B2( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n165 ) , .B1( u1_u12_u3_n167 ) );
  NOR2_X1 u1_u12_u3_U48 (.A1( u1_u12_u3_n113 ) , .ZN( u1_u12_u3_n131 ) , .A2( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U49 (.A1( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n150 ) , .A2( u1_u12_u3_n99 ) );
  INV_X1 u1_u12_u3_U5 (.A( u1_u12_u3_n117 ) , .ZN( u1_u12_u3_n178 ) );
  NAND2_X1 u1_u12_u3_U50 (.A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n155 ) , .A1( u1_u12_u3_n97 ) );
  INV_X1 u1_u12_u3_U51 (.A( u1_u12_u3_n141 ) , .ZN( u1_u12_u3_n167 ) );
  AOI21_X1 u1_u12_u3_U52 (.B2( u1_u12_u3_n114 ) , .B1( u1_u12_u3_n146 ) , .A( u1_u12_u3_n154 ) , .ZN( u1_u12_u3_n94 ) );
  AOI21_X1 u1_u12_u3_U53 (.ZN( u1_u12_u3_n110 ) , .B2( u1_u12_u3_n142 ) , .B1( u1_u12_u3_n186 ) , .A( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U54 (.A( u1_u12_u3_n145 ) , .ZN( u1_u12_u3_n186 ) );
  AOI21_X1 u1_u12_u3_U55 (.B1( u1_u12_u3_n124 ) , .A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U56 (.A( u1_u12_u3_n149 ) , .ZN( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U57 (.ZN( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n96 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U58 (.A2( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n146 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U59 (.A1( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n99 ) );
  AOI221_X1 u1_u12_u3_U6 (.A( u1_u12_u3_n131 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n134 ) , .B1( u1_u12_u3_n143 ) , .B2( u1_u12_u3_n177 ) );
  NAND2_X1 u1_u12_u3_U60 (.A1( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n156 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U61 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U62 (.A1( u1_u12_u3_n100 ) , .A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n128 ) );
  NAND2_X1 u1_u12_u3_U63 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n152 ) );
  NAND2_X1 u1_u12_u3_U64 (.A2( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n114 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U65 (.ZN( u1_u12_u3_n107 ) , .A1( u1_u12_u3_n97 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U66 (.A2( u1_u12_u3_n100 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n113 ) );
  NAND2_X1 u1_u12_u3_U67 (.A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n153 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U68 (.A2( u1_u12_u3_n103 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n130 ) );
  NAND2_X1 u1_u12_u3_U69 (.A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n96 ) );
  OAI22_X1 u1_u12_u3_U7 (.B2( u1_u12_u3_n147 ) , .A2( u1_u12_u3_n148 ) , .ZN( u1_u12_u3_n160 ) , .B1( u1_u12_u3_n165 ) , .A1( u1_u12_u3_n168 ) );
  NAND2_X1 u1_u12_u3_U70 (.A1( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n108 ) );
  NOR2_X1 u1_u12_u3_U71 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n99 ) );
  NOR2_X1 u1_u12_u3_U72 (.A2( u1_u12_X_21 ) , .A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n103 ) );
  NOR2_X1 u1_u12_u3_U73 (.A2( u1_u12_X_24 ) , .A1( u1_u12_u3_n171 ) , .ZN( u1_u12_u3_n97 ) );
  NOR2_X1 u1_u12_u3_U74 (.A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U75 (.A2( u1_u12_X_19 ) , .A1( u1_u12_u3_n172 ) , .ZN( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U76 (.A1( u1_u12_X_22 ) , .A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U77 (.A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n149 ) , .A2( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U78 (.A2( u1_u12_X_22 ) , .A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n121 ) );
  AND2_X1 u1_u12_u3_U79 (.A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n101 ) , .A2( u1_u12_u3_n171 ) );
  AND3_X1 u1_u12_u3_U8 (.A3( u1_u12_u3_n144 ) , .A2( u1_u12_u3_n145 ) , .A1( u1_u12_u3_n146 ) , .ZN( u1_u12_u3_n147 ) );
  AND2_X1 u1_u12_u3_U80 (.A1( u1_u12_X_19 ) , .ZN( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n172 ) );
  AND2_X1 u1_u12_u3_U81 (.A1( u1_u12_X_21 ) , .A2( u1_u12_X_24 ) , .ZN( u1_u12_u3_n100 ) );
  AND2_X1 u1_u12_u3_U82 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n104 ) );
  INV_X1 u1_u12_u3_U83 (.A( u1_u12_X_22 ) , .ZN( u1_u12_u3_n166 ) );
  INV_X1 u1_u12_u3_U84 (.A( u1_u12_X_21 ) , .ZN( u1_u12_u3_n171 ) );
  INV_X1 u1_u12_u3_U85 (.A( u1_u12_X_20 ) , .ZN( u1_u12_u3_n172 ) );
  NAND4_X1 u1_u12_u3_U86 (.ZN( u1_out12_26 ) , .A4( u1_u12_u3_n109 ) , .A3( u1_u12_u3_n110 ) , .A2( u1_u12_u3_n111 ) , .A1( u1_u12_u3_n173 ) );
  INV_X1 u1_u12_u3_U87 (.ZN( u1_u12_u3_n173 ) , .A( u1_u12_u3_n94 ) );
  OAI21_X1 u1_u12_u3_U88 (.ZN( u1_u12_u3_n111 ) , .B2( u1_u12_u3_n117 ) , .A( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n176 ) );
  NAND4_X1 u1_u12_u3_U89 (.ZN( u1_out12_20 ) , .A4( u1_u12_u3_n122 ) , .A3( u1_u12_u3_n123 ) , .A1( u1_u12_u3_n175 ) , .A2( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U9 (.A( u1_u12_u3_n143 ) , .ZN( u1_u12_u3_n168 ) );
  INV_X1 u1_u12_u3_U90 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U91 (.A( u1_u12_u3_n112 ) , .ZN( u1_u12_u3_n175 ) );
  NAND4_X1 u1_u12_u3_U92 (.ZN( u1_out12_1 ) , .A4( u1_u12_u3_n161 ) , .A3( u1_u12_u3_n162 ) , .A2( u1_u12_u3_n163 ) , .A1( u1_u12_u3_n185 ) );
  NAND2_X1 u1_u12_u3_U93 (.ZN( u1_u12_u3_n163 ) , .A2( u1_u12_u3_n170 ) , .A1( u1_u12_u3_n176 ) );
  AOI22_X1 u1_u12_u3_U94 (.B2( u1_u12_u3_n140 ) , .B1( u1_u12_u3_n141 ) , .A2( u1_u12_u3_n142 ) , .ZN( u1_u12_u3_n162 ) , .A1( u1_u12_u3_n177 ) );
  OR4_X1 u1_u12_u3_U95 (.ZN( u1_out12_10 ) , .A4( u1_u12_u3_n136 ) , .A3( u1_u12_u3_n137 ) , .A1( u1_u12_u3_n138 ) , .A2( u1_u12_u3_n139 ) );
  OAI222_X1 u1_u12_u3_U96 (.C1( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n137 ) , .B1( u1_u12_u3_n148 ) , .A2( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n154 ) , .C2( u1_u12_u3_n164 ) , .A1( u1_u12_u3_n167 ) );
  OAI221_X1 u1_u12_u3_U97 (.A( u1_u12_u3_n134 ) , .B2( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n136 ) , .C1( u1_u12_u3_n149 ) , .B1( u1_u12_u3_n151 ) , .C2( u1_u12_u3_n183 ) );
  NAND3_X1 u1_u12_u3_U98 (.A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n145 ) , .A3( u1_u12_u3_n153 ) );
  NAND3_X1 u1_u12_u3_U99 (.ZN( u1_u12_u3_n129 ) , .A2( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n153 ) , .A3( u1_u12_u3_n182 ) );
  XOR2_X1 u1_u15_U40 (.A( u1_FP_45 ) , .B( u1_K16_18 ) , .Z( u1_u15_X_18 ) );
  XOR2_X1 u1_u15_U41 (.A( u1_FP_44 ) , .B( u1_K16_17 ) , .Z( u1_u15_X_17 ) );
  XOR2_X1 u1_u15_U42 (.A( u1_FP_43 ) , .B( u1_K16_16 ) , .Z( u1_u15_X_16 ) );
  XOR2_X1 u1_u15_U43 (.A( u1_FP_42 ) , .B( u1_K16_15 ) , .Z( u1_u15_X_15 ) );
  XOR2_X1 u1_u15_U44 (.A( u1_FP_41 ) , .B( u1_K16_14 ) , .Z( u1_u15_X_14 ) );
  XOR2_X1 u1_u15_U45 (.A( u1_FP_40 ) , .B( u1_K16_13 ) , .Z( u1_u15_X_13 ) );
  OAI22_X1 u1_u15_u2_U10 (.B1( u1_u15_u2_n151 ) , .A2( u1_u15_u2_n152 ) , .A1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n160 ) , .B2( u1_u15_u2_n168 ) );
  NAND3_X1 u1_u15_u2_U100 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n98 ) );
  NOR3_X1 u1_u15_u2_U11 (.A1( u1_u15_u2_n150 ) , .ZN( u1_u15_u2_n151 ) , .A3( u1_u15_u2_n175 ) , .A2( u1_u15_u2_n188 ) );
  AOI21_X1 u1_u15_u2_U12 (.B2( u1_u15_u2_n123 ) , .ZN( u1_u15_u2_n125 ) , .A( u1_u15_u2_n171 ) , .B1( u1_u15_u2_n184 ) );
  INV_X1 u1_u15_u2_U13 (.A( u1_u15_u2_n150 ) , .ZN( u1_u15_u2_n184 ) );
  AOI21_X1 u1_u15_u2_U14 (.ZN( u1_u15_u2_n144 ) , .B2( u1_u15_u2_n155 ) , .A( u1_u15_u2_n172 ) , .B1( u1_u15_u2_n185 ) );
  AOI21_X1 u1_u15_u2_U15 (.B2( u1_u15_u2_n143 ) , .ZN( u1_u15_u2_n145 ) , .B1( u1_u15_u2_n152 ) , .A( u1_u15_u2_n171 ) );
  INV_X1 u1_u15_u2_U16 (.A( u1_u15_u2_n156 ) , .ZN( u1_u15_u2_n171 ) );
  INV_X1 u1_u15_u2_U17 (.A( u1_u15_u2_n120 ) , .ZN( u1_u15_u2_n188 ) );
  NAND2_X1 u1_u15_u2_U18 (.A2( u1_u15_u2_n122 ) , .ZN( u1_u15_u2_n150 ) , .A1( u1_u15_u2_n152 ) );
  INV_X1 u1_u15_u2_U19 (.A( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n170 ) );
  INV_X1 u1_u15_u2_U20 (.A( u1_u15_u2_n137 ) , .ZN( u1_u15_u2_n173 ) );
  NAND2_X1 u1_u15_u2_U21 (.A1( u1_u15_u2_n132 ) , .A2( u1_u15_u2_n139 ) , .ZN( u1_u15_u2_n157 ) );
  INV_X1 u1_u15_u2_U22 (.A( u1_u15_u2_n113 ) , .ZN( u1_u15_u2_n178 ) );
  INV_X1 u1_u15_u2_U23 (.A( u1_u15_u2_n139 ) , .ZN( u1_u15_u2_n175 ) );
  INV_X1 u1_u15_u2_U24 (.A( u1_u15_u2_n155 ) , .ZN( u1_u15_u2_n181 ) );
  INV_X1 u1_u15_u2_U25 (.A( u1_u15_u2_n119 ) , .ZN( u1_u15_u2_n177 ) );
  INV_X1 u1_u15_u2_U26 (.A( u1_u15_u2_n116 ) , .ZN( u1_u15_u2_n180 ) );
  INV_X1 u1_u15_u2_U27 (.A( u1_u15_u2_n131 ) , .ZN( u1_u15_u2_n179 ) );
  INV_X1 u1_u15_u2_U28 (.A( u1_u15_u2_n154 ) , .ZN( u1_u15_u2_n176 ) );
  NAND2_X1 u1_u15_u2_U29 (.A2( u1_u15_u2_n116 ) , .A1( u1_u15_u2_n117 ) , .ZN( u1_u15_u2_n118 ) );
  NOR2_X1 u1_u15_u2_U3 (.ZN( u1_u15_u2_n121 ) , .A2( u1_u15_u2_n177 ) , .A1( u1_u15_u2_n180 ) );
  INV_X1 u1_u15_u2_U30 (.A( u1_u15_u2_n132 ) , .ZN( u1_u15_u2_n182 ) );
  INV_X1 u1_u15_u2_U31 (.A( u1_u15_u2_n158 ) , .ZN( u1_u15_u2_n183 ) );
  OAI21_X1 u1_u15_u2_U32 (.A( u1_u15_u2_n156 ) , .B1( u1_u15_u2_n157 ) , .ZN( u1_u15_u2_n158 ) , .B2( u1_u15_u2_n179 ) );
  NOR2_X1 u1_u15_u2_U33 (.ZN( u1_u15_u2_n156 ) , .A1( u1_u15_u2_n166 ) , .A2( u1_u15_u2_n169 ) );
  NOR2_X1 u1_u15_u2_U34 (.A2( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n137 ) , .A1( u1_u15_u2_n140 ) );
  NOR2_X1 u1_u15_u2_U35 (.A2( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n153 ) , .A1( u1_u15_u2_n156 ) );
  AOI211_X1 u1_u15_u2_U36 (.ZN( u1_u15_u2_n130 ) , .C1( u1_u15_u2_n138 ) , .C2( u1_u15_u2_n179 ) , .B( u1_u15_u2_n96 ) , .A( u1_u15_u2_n97 ) );
  OAI22_X1 u1_u15_u2_U37 (.B1( u1_u15_u2_n133 ) , .A2( u1_u15_u2_n137 ) , .A1( u1_u15_u2_n152 ) , .B2( u1_u15_u2_n168 ) , .ZN( u1_u15_u2_n97 ) );
  OAI221_X1 u1_u15_u2_U38 (.B1( u1_u15_u2_n113 ) , .C1( u1_u15_u2_n132 ) , .A( u1_u15_u2_n149 ) , .B2( u1_u15_u2_n171 ) , .C2( u1_u15_u2_n172 ) , .ZN( u1_u15_u2_n96 ) );
  OAI221_X1 u1_u15_u2_U39 (.A( u1_u15_u2_n115 ) , .C2( u1_u15_u2_n123 ) , .B2( u1_u15_u2_n143 ) , .B1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n163 ) , .C1( u1_u15_u2_n168 ) );
  INV_X1 u1_u15_u2_U4 (.A( u1_u15_u2_n134 ) , .ZN( u1_u15_u2_n185 ) );
  OAI21_X1 u1_u15_u2_U40 (.A( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n115 ) , .B1( u1_u15_u2_n176 ) , .B2( u1_u15_u2_n178 ) );
  OAI221_X1 u1_u15_u2_U41 (.A( u1_u15_u2_n135 ) , .B2( u1_u15_u2_n136 ) , .B1( u1_u15_u2_n137 ) , .ZN( u1_u15_u2_n162 ) , .C2( u1_u15_u2_n167 ) , .C1( u1_u15_u2_n185 ) );
  AND3_X1 u1_u15_u2_U42 (.A3( u1_u15_u2_n131 ) , .A2( u1_u15_u2_n132 ) , .A1( u1_u15_u2_n133 ) , .ZN( u1_u15_u2_n136 ) );
  AOI22_X1 u1_u15_u2_U43 (.ZN( u1_u15_u2_n135 ) , .B1( u1_u15_u2_n140 ) , .A1( u1_u15_u2_n156 ) , .B2( u1_u15_u2_n180 ) , .A2( u1_u15_u2_n188 ) );
  AOI21_X1 u1_u15_u2_U44 (.ZN( u1_u15_u2_n149 ) , .B1( u1_u15_u2_n173 ) , .B2( u1_u15_u2_n188 ) , .A( u1_u15_u2_n95 ) );
  AND3_X1 u1_u15_u2_U45 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n156 ) , .ZN( u1_u15_u2_n95 ) );
  OAI21_X1 u1_u15_u2_U46 (.A( u1_u15_u2_n101 ) , .B2( u1_u15_u2_n121 ) , .B1( u1_u15_u2_n153 ) , .ZN( u1_u15_u2_n164 ) );
  NAND2_X1 u1_u15_u2_U47 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n155 ) );
  NAND2_X1 u1_u15_u2_U48 (.A2( u1_u15_u2_n105 ) , .A1( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n143 ) );
  NAND2_X1 u1_u15_u2_U49 (.A1( u1_u15_u2_n104 ) , .A2( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n152 ) );
  NOR4_X1 u1_u15_u2_U5 (.A4( u1_u15_u2_n124 ) , .A3( u1_u15_u2_n125 ) , .A2( u1_u15_u2_n126 ) , .A1( u1_u15_u2_n127 ) , .ZN( u1_u15_u2_n128 ) );
  NAND2_X1 u1_u15_u2_U50 (.A1( u1_u15_u2_n100 ) , .A2( u1_u15_u2_n105 ) , .ZN( u1_u15_u2_n132 ) );
  INV_X1 u1_u15_u2_U51 (.A( u1_u15_u2_n140 ) , .ZN( u1_u15_u2_n168 ) );
  INV_X1 u1_u15_u2_U52 (.A( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n167 ) );
  OAI21_X1 u1_u15_u2_U53 (.A( u1_u15_u2_n141 ) , .B2( u1_u15_u2_n142 ) , .ZN( u1_u15_u2_n146 ) , .B1( u1_u15_u2_n153 ) );
  OAI21_X1 u1_u15_u2_U54 (.A( u1_u15_u2_n140 ) , .ZN( u1_u15_u2_n141 ) , .B1( u1_u15_u2_n176 ) , .B2( u1_u15_u2_n177 ) );
  NOR3_X1 u1_u15_u2_U55 (.ZN( u1_u15_u2_n142 ) , .A3( u1_u15_u2_n175 ) , .A2( u1_u15_u2_n178 ) , .A1( u1_u15_u2_n181 ) );
  INV_X1 u1_u15_u2_U56 (.ZN( u1_u15_u2_n187 ) , .A( u1_u15_u2_n99 ) );
  OAI21_X1 u1_u15_u2_U57 (.B1( u1_u15_u2_n137 ) , .B2( u1_u15_u2_n143 ) , .A( u1_u15_u2_n98 ) , .ZN( u1_u15_u2_n99 ) );
  NAND2_X1 u1_u15_u2_U58 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n113 ) );
  NAND2_X1 u1_u15_u2_U59 (.A1( u1_u15_u2_n106 ) , .A2( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n131 ) );
  AOI21_X1 u1_u15_u2_U6 (.B2( u1_u15_u2_n119 ) , .ZN( u1_u15_u2_n127 ) , .A( u1_u15_u2_n137 ) , .B1( u1_u15_u2_n155 ) );
  NAND2_X1 u1_u15_u2_U60 (.A1( u1_u15_u2_n103 ) , .A2( u1_u15_u2_n107 ) , .ZN( u1_u15_u2_n139 ) );
  NAND2_X1 u1_u15_u2_U61 (.A1( u1_u15_u2_n103 ) , .A2( u1_u15_u2_n105 ) , .ZN( u1_u15_u2_n133 ) );
  NAND2_X1 u1_u15_u2_U62 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n103 ) , .ZN( u1_u15_u2_n154 ) );
  NAND2_X1 u1_u15_u2_U63 (.A2( u1_u15_u2_n103 ) , .A1( u1_u15_u2_n104 ) , .ZN( u1_u15_u2_n119 ) );
  NAND2_X1 u1_u15_u2_U64 (.A2( u1_u15_u2_n107 ) , .A1( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n123 ) );
  NAND2_X1 u1_u15_u2_U65 (.A1( u1_u15_u2_n104 ) , .A2( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n122 ) );
  INV_X1 u1_u15_u2_U66 (.A( u1_u15_u2_n114 ) , .ZN( u1_u15_u2_n172 ) );
  NAND2_X1 u1_u15_u2_U67 (.A2( u1_u15_u2_n100 ) , .A1( u1_u15_u2_n102 ) , .ZN( u1_u15_u2_n116 ) );
  NAND2_X1 u1_u15_u2_U68 (.A1( u1_u15_u2_n102 ) , .A2( u1_u15_u2_n108 ) , .ZN( u1_u15_u2_n120 ) );
  NAND2_X1 u1_u15_u2_U69 (.A2( u1_u15_u2_n105 ) , .A1( u1_u15_u2_n106 ) , .ZN( u1_u15_u2_n117 ) );
  AOI21_X1 u1_u15_u2_U7 (.ZN( u1_u15_u2_n124 ) , .B1( u1_u15_u2_n131 ) , .B2( u1_u15_u2_n143 ) , .A( u1_u15_u2_n172 ) );
  NOR2_X1 u1_u15_u2_U70 (.A2( u1_u15_X_16 ) , .ZN( u1_u15_u2_n140 ) , .A1( u1_u15_u2_n166 ) );
  NOR2_X1 u1_u15_u2_U71 (.A2( u1_u15_X_13 ) , .A1( u1_u15_X_14 ) , .ZN( u1_u15_u2_n100 ) );
  NOR2_X1 u1_u15_u2_U72 (.A2( u1_u15_X_16 ) , .A1( u1_u15_X_17 ) , .ZN( u1_u15_u2_n138 ) );
  NOR2_X1 u1_u15_u2_U73 (.A2( u1_u15_X_15 ) , .A1( u1_u15_X_18 ) , .ZN( u1_u15_u2_n104 ) );
  NOR2_X1 u1_u15_u2_U74 (.A2( u1_u15_X_14 ) , .ZN( u1_u15_u2_n103 ) , .A1( u1_u15_u2_n174 ) );
  NOR2_X1 u1_u15_u2_U75 (.A2( u1_u15_X_15 ) , .ZN( u1_u15_u2_n102 ) , .A1( u1_u15_u2_n165 ) );
  NOR2_X1 u1_u15_u2_U76 (.A2( u1_u15_X_17 ) , .ZN( u1_u15_u2_n114 ) , .A1( u1_u15_u2_n169 ) );
  AND2_X1 u1_u15_u2_U77 (.A1( u1_u15_X_15 ) , .ZN( u1_u15_u2_n105 ) , .A2( u1_u15_u2_n165 ) );
  AND2_X1 u1_u15_u2_U78 (.A2( u1_u15_X_15 ) , .A1( u1_u15_X_18 ) , .ZN( u1_u15_u2_n107 ) );
  AND2_X1 u1_u15_u2_U79 (.A1( u1_u15_X_14 ) , .ZN( u1_u15_u2_n106 ) , .A2( u1_u15_u2_n174 ) );
  AOI21_X1 u1_u15_u2_U8 (.B2( u1_u15_u2_n120 ) , .B1( u1_u15_u2_n121 ) , .ZN( u1_u15_u2_n126 ) , .A( u1_u15_u2_n167 ) );
  AND2_X1 u1_u15_u2_U80 (.A1( u1_u15_X_13 ) , .A2( u1_u15_X_14 ) , .ZN( u1_u15_u2_n108 ) );
  INV_X1 u1_u15_u2_U81 (.A( u1_u15_X_16 ) , .ZN( u1_u15_u2_n169 ) );
  INV_X1 u1_u15_u2_U82 (.A( u1_u15_X_17 ) , .ZN( u1_u15_u2_n166 ) );
  INV_X1 u1_u15_u2_U83 (.A( u1_u15_X_13 ) , .ZN( u1_u15_u2_n174 ) );
  INV_X1 u1_u15_u2_U84 (.A( u1_u15_X_18 ) , .ZN( u1_u15_u2_n165 ) );
  NAND4_X1 u1_u15_u2_U85 (.ZN( u1_out15_30 ) , .A4( u1_u15_u2_n147 ) , .A3( u1_u15_u2_n148 ) , .A2( u1_u15_u2_n149 ) , .A1( u1_u15_u2_n187 ) );
  NOR3_X1 u1_u15_u2_U86 (.A3( u1_u15_u2_n144 ) , .A2( u1_u15_u2_n145 ) , .A1( u1_u15_u2_n146 ) , .ZN( u1_u15_u2_n147 ) );
  AOI21_X1 u1_u15_u2_U87 (.B2( u1_u15_u2_n138 ) , .ZN( u1_u15_u2_n148 ) , .A( u1_u15_u2_n162 ) , .B1( u1_u15_u2_n182 ) );
  NAND4_X1 u1_u15_u2_U88 (.ZN( u1_out15_24 ) , .A4( u1_u15_u2_n111 ) , .A3( u1_u15_u2_n112 ) , .A1( u1_u15_u2_n130 ) , .A2( u1_u15_u2_n187 ) );
  AOI221_X1 u1_u15_u2_U89 (.A( u1_u15_u2_n109 ) , .B1( u1_u15_u2_n110 ) , .ZN( u1_u15_u2_n111 ) , .C1( u1_u15_u2_n134 ) , .C2( u1_u15_u2_n170 ) , .B2( u1_u15_u2_n173 ) );
  OAI22_X1 u1_u15_u2_U9 (.ZN( u1_u15_u2_n109 ) , .A2( u1_u15_u2_n113 ) , .B2( u1_u15_u2_n133 ) , .B1( u1_u15_u2_n167 ) , .A1( u1_u15_u2_n168 ) );
  AOI21_X1 u1_u15_u2_U90 (.ZN( u1_u15_u2_n112 ) , .B2( u1_u15_u2_n156 ) , .A( u1_u15_u2_n164 ) , .B1( u1_u15_u2_n181 ) );
  NAND4_X1 u1_u15_u2_U91 (.ZN( u1_out15_16 ) , .A4( u1_u15_u2_n128 ) , .A3( u1_u15_u2_n129 ) , .A1( u1_u15_u2_n130 ) , .A2( u1_u15_u2_n186 ) );
  AOI22_X1 u1_u15_u2_U92 (.A2( u1_u15_u2_n118 ) , .ZN( u1_u15_u2_n129 ) , .A1( u1_u15_u2_n140 ) , .B1( u1_u15_u2_n157 ) , .B2( u1_u15_u2_n170 ) );
  INV_X1 u1_u15_u2_U93 (.A( u1_u15_u2_n163 ) , .ZN( u1_u15_u2_n186 ) );
  OR4_X1 u1_u15_u2_U94 (.ZN( u1_out15_6 ) , .A4( u1_u15_u2_n161 ) , .A3( u1_u15_u2_n162 ) , .A2( u1_u15_u2_n163 ) , .A1( u1_u15_u2_n164 ) );
  OR3_X1 u1_u15_u2_U95 (.A2( u1_u15_u2_n159 ) , .A1( u1_u15_u2_n160 ) , .ZN( u1_u15_u2_n161 ) , .A3( u1_u15_u2_n183 ) );
  AOI21_X1 u1_u15_u2_U96 (.B2( u1_u15_u2_n154 ) , .B1( u1_u15_u2_n155 ) , .ZN( u1_u15_u2_n159 ) , .A( u1_u15_u2_n167 ) );
  NAND3_X1 u1_u15_u2_U97 (.A2( u1_u15_u2_n117 ) , .A1( u1_u15_u2_n122 ) , .A3( u1_u15_u2_n123 ) , .ZN( u1_u15_u2_n134 ) );
  NAND3_X1 u1_u15_u2_U98 (.ZN( u1_u15_u2_n110 ) , .A2( u1_u15_u2_n131 ) , .A3( u1_u15_u2_n139 ) , .A1( u1_u15_u2_n154 ) );
  NAND3_X1 u1_u15_u2_U99 (.A2( u1_u15_u2_n100 ) , .ZN( u1_u15_u2_n101 ) , .A1( u1_u15_u2_n104 ) , .A3( u1_u15_u2_n114 ) );
  XOR2_X1 u1_u1_U1 (.B( u1_K2_9 ) , .A( u1_R0_6 ) , .Z( u1_u1_X_9 ) );
  XOR2_X1 u1_u1_U2 (.B( u1_K2_8 ) , .A( u1_R0_5 ) , .Z( u1_u1_X_8 ) );
  XOR2_X1 u1_u1_U3 (.B( u1_K2_7 ) , .A( u1_R0_4 ) , .Z( u1_u1_X_7 ) );
  XOR2_X1 u1_u1_U40 (.B( u1_K2_18 ) , .A( u1_R0_13 ) , .Z( u1_u1_X_18 ) );
  XOR2_X1 u1_u1_U41 (.B( u1_K2_17 ) , .A( u1_R0_12 ) , .Z( u1_u1_X_17 ) );
  XOR2_X1 u1_u1_U42 (.B( u1_K2_16 ) , .A( u1_R0_11 ) , .Z( u1_u1_X_16 ) );
  XOR2_X1 u1_u1_U43 (.B( u1_K2_15 ) , .A( u1_R0_10 ) , .Z( u1_u1_X_15 ) );
  XOR2_X1 u1_u1_U44 (.B( u1_K2_14 ) , .A( u1_R0_9 ) , .Z( u1_u1_X_14 ) );
  XOR2_X1 u1_u1_U45 (.B( u1_K2_13 ) , .A( u1_R0_8 ) , .Z( u1_u1_X_13 ) );
  XOR2_X1 u1_u1_U46 (.B( u1_K2_12 ) , .A( u1_R0_9 ) , .Z( u1_u1_X_12 ) );
  XOR2_X1 u1_u1_U47 (.B( u1_K2_11 ) , .A( u1_R0_8 ) , .Z( u1_u1_X_11 ) );
  XOR2_X1 u1_u1_U48 (.B( u1_K2_10 ) , .A( u1_R0_7 ) , .Z( u1_u1_X_10 ) );
  NOR2_X1 u1_u1_u1_U10 (.A1( u1_u1_u1_n112 ) , .A2( u1_u1_u1_n116 ) , .ZN( u1_u1_u1_n118 ) );
  NAND3_X1 u1_u1_u1_U100 (.ZN( u1_u1_u1_n113 ) , .A1( u1_u1_u1_n120 ) , .A3( u1_u1_u1_n133 ) , .A2( u1_u1_u1_n155 ) );
  OAI21_X1 u1_u1_u1_U11 (.ZN( u1_u1_u1_n101 ) , .B1( u1_u1_u1_n141 ) , .A( u1_u1_u1_n146 ) , .B2( u1_u1_u1_n183 ) );
  AOI21_X1 u1_u1_u1_U12 (.B2( u1_u1_u1_n155 ) , .B1( u1_u1_u1_n156 ) , .ZN( u1_u1_u1_n157 ) , .A( u1_u1_u1_n174 ) );
  NAND2_X1 u1_u1_u1_U13 (.ZN( u1_u1_u1_n140 ) , .A2( u1_u1_u1_n150 ) , .A1( u1_u1_u1_n155 ) );
  NAND2_X1 u1_u1_u1_U14 (.A1( u1_u1_u1_n131 ) , .ZN( u1_u1_u1_n147 ) , .A2( u1_u1_u1_n153 ) );
  INV_X1 u1_u1_u1_U15 (.A( u1_u1_u1_n139 ) , .ZN( u1_u1_u1_n174 ) );
  OR4_X1 u1_u1_u1_U16 (.A4( u1_u1_u1_n106 ) , .A3( u1_u1_u1_n107 ) , .ZN( u1_u1_u1_n108 ) , .A1( u1_u1_u1_n117 ) , .A2( u1_u1_u1_n184 ) );
  AOI21_X1 u1_u1_u1_U17 (.ZN( u1_u1_u1_n106 ) , .A( u1_u1_u1_n112 ) , .B1( u1_u1_u1_n154 ) , .B2( u1_u1_u1_n156 ) );
  INV_X1 u1_u1_u1_U18 (.A( u1_u1_u1_n101 ) , .ZN( u1_u1_u1_n184 ) );
  AOI21_X1 u1_u1_u1_U19 (.ZN( u1_u1_u1_n107 ) , .B1( u1_u1_u1_n134 ) , .B2( u1_u1_u1_n149 ) , .A( u1_u1_u1_n174 ) );
  INV_X1 u1_u1_u1_U20 (.A( u1_u1_u1_n112 ) , .ZN( u1_u1_u1_n171 ) );
  NAND2_X1 u1_u1_u1_U21 (.ZN( u1_u1_u1_n141 ) , .A1( u1_u1_u1_n153 ) , .A2( u1_u1_u1_n156 ) );
  AND2_X1 u1_u1_u1_U22 (.A1( u1_u1_u1_n123 ) , .ZN( u1_u1_u1_n134 ) , .A2( u1_u1_u1_n161 ) );
  NAND2_X1 u1_u1_u1_U23 (.A2( u1_u1_u1_n115 ) , .A1( u1_u1_u1_n116 ) , .ZN( u1_u1_u1_n148 ) );
  NAND2_X1 u1_u1_u1_U24 (.A2( u1_u1_u1_n133 ) , .A1( u1_u1_u1_n135 ) , .ZN( u1_u1_u1_n159 ) );
  NAND2_X1 u1_u1_u1_U25 (.A2( u1_u1_u1_n115 ) , .A1( u1_u1_u1_n120 ) , .ZN( u1_u1_u1_n132 ) );
  INV_X1 u1_u1_u1_U26 (.A( u1_u1_u1_n154 ) , .ZN( u1_u1_u1_n178 ) );
  INV_X1 u1_u1_u1_U27 (.A( u1_u1_u1_n151 ) , .ZN( u1_u1_u1_n183 ) );
  AND2_X1 u1_u1_u1_U28 (.A1( u1_u1_u1_n129 ) , .A2( u1_u1_u1_n133 ) , .ZN( u1_u1_u1_n149 ) );
  INV_X1 u1_u1_u1_U29 (.A( u1_u1_u1_n131 ) , .ZN( u1_u1_u1_n180 ) );
  INV_X1 u1_u1_u1_U3 (.A( u1_u1_u1_n159 ) , .ZN( u1_u1_u1_n182 ) );
  AOI221_X1 u1_u1_u1_U30 (.B1( u1_u1_u1_n140 ) , .ZN( u1_u1_u1_n167 ) , .B2( u1_u1_u1_n172 ) , .C2( u1_u1_u1_n175 ) , .C1( u1_u1_u1_n178 ) , .A( u1_u1_u1_n188 ) );
  INV_X1 u1_u1_u1_U31 (.ZN( u1_u1_u1_n188 ) , .A( u1_u1_u1_n97 ) );
  AOI211_X1 u1_u1_u1_U32 (.A( u1_u1_u1_n118 ) , .C1( u1_u1_u1_n132 ) , .C2( u1_u1_u1_n139 ) , .B( u1_u1_u1_n96 ) , .ZN( u1_u1_u1_n97 ) );
  AOI21_X1 u1_u1_u1_U33 (.B2( u1_u1_u1_n121 ) , .B1( u1_u1_u1_n135 ) , .A( u1_u1_u1_n152 ) , .ZN( u1_u1_u1_n96 ) );
  OAI221_X1 u1_u1_u1_U34 (.A( u1_u1_u1_n119 ) , .C2( u1_u1_u1_n129 ) , .ZN( u1_u1_u1_n138 ) , .B2( u1_u1_u1_n152 ) , .C1( u1_u1_u1_n174 ) , .B1( u1_u1_u1_n187 ) );
  INV_X1 u1_u1_u1_U35 (.A( u1_u1_u1_n148 ) , .ZN( u1_u1_u1_n187 ) );
  AOI211_X1 u1_u1_u1_U36 (.B( u1_u1_u1_n117 ) , .A( u1_u1_u1_n118 ) , .ZN( u1_u1_u1_n119 ) , .C2( u1_u1_u1_n146 ) , .C1( u1_u1_u1_n159 ) );
  NOR2_X1 u1_u1_u1_U37 (.A1( u1_u1_u1_n168 ) , .A2( u1_u1_u1_n176 ) , .ZN( u1_u1_u1_n98 ) );
  AOI211_X1 u1_u1_u1_U38 (.B( u1_u1_u1_n162 ) , .A( u1_u1_u1_n163 ) , .C2( u1_u1_u1_n164 ) , .ZN( u1_u1_u1_n165 ) , .C1( u1_u1_u1_n171 ) );
  AOI21_X1 u1_u1_u1_U39 (.A( u1_u1_u1_n160 ) , .B2( u1_u1_u1_n161 ) , .ZN( u1_u1_u1_n162 ) , .B1( u1_u1_u1_n182 ) );
  AOI221_X1 u1_u1_u1_U4 (.A( u1_u1_u1_n138 ) , .C2( u1_u1_u1_n139 ) , .C1( u1_u1_u1_n140 ) , .B2( u1_u1_u1_n141 ) , .ZN( u1_u1_u1_n142 ) , .B1( u1_u1_u1_n175 ) );
  OR2_X1 u1_u1_u1_U40 (.A2( u1_u1_u1_n157 ) , .A1( u1_u1_u1_n158 ) , .ZN( u1_u1_u1_n163 ) );
  OAI21_X1 u1_u1_u1_U41 (.B2( u1_u1_u1_n123 ) , .ZN( u1_u1_u1_n145 ) , .B1( u1_u1_u1_n160 ) , .A( u1_u1_u1_n185 ) );
  INV_X1 u1_u1_u1_U42 (.A( u1_u1_u1_n122 ) , .ZN( u1_u1_u1_n185 ) );
  AOI21_X1 u1_u1_u1_U43 (.B2( u1_u1_u1_n120 ) , .B1( u1_u1_u1_n121 ) , .ZN( u1_u1_u1_n122 ) , .A( u1_u1_u1_n128 ) );
  NAND2_X1 u1_u1_u1_U44 (.A1( u1_u1_u1_n128 ) , .ZN( u1_u1_u1_n146 ) , .A2( u1_u1_u1_n160 ) );
  NAND2_X1 u1_u1_u1_U45 (.A2( u1_u1_u1_n112 ) , .ZN( u1_u1_u1_n139 ) , .A1( u1_u1_u1_n152 ) );
  NAND2_X1 u1_u1_u1_U46 (.A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n156 ) , .A2( u1_u1_u1_n99 ) );
  NOR2_X1 u1_u1_u1_U47 (.ZN( u1_u1_u1_n117 ) , .A1( u1_u1_u1_n121 ) , .A2( u1_u1_u1_n160 ) );
  AOI21_X1 u1_u1_u1_U48 (.A( u1_u1_u1_n128 ) , .B2( u1_u1_u1_n129 ) , .ZN( u1_u1_u1_n130 ) , .B1( u1_u1_u1_n150 ) );
  NAND2_X1 u1_u1_u1_U49 (.ZN( u1_u1_u1_n112 ) , .A1( u1_u1_u1_n169 ) , .A2( u1_u1_u1_n170 ) );
  AOI211_X1 u1_u1_u1_U5 (.ZN( u1_u1_u1_n124 ) , .A( u1_u1_u1_n138 ) , .C2( u1_u1_u1_n139 ) , .B( u1_u1_u1_n145 ) , .C1( u1_u1_u1_n147 ) );
  NAND2_X1 u1_u1_u1_U50 (.ZN( u1_u1_u1_n129 ) , .A2( u1_u1_u1_n95 ) , .A1( u1_u1_u1_n98 ) );
  NAND2_X1 u1_u1_u1_U51 (.A1( u1_u1_u1_n102 ) , .ZN( u1_u1_u1_n154 ) , .A2( u1_u1_u1_n99 ) );
  NAND2_X1 u1_u1_u1_U52 (.A2( u1_u1_u1_n100 ) , .ZN( u1_u1_u1_n135 ) , .A1( u1_u1_u1_n99 ) );
  AOI21_X1 u1_u1_u1_U53 (.A( u1_u1_u1_n152 ) , .B2( u1_u1_u1_n153 ) , .B1( u1_u1_u1_n154 ) , .ZN( u1_u1_u1_n158 ) );
  INV_X1 u1_u1_u1_U54 (.A( u1_u1_u1_n160 ) , .ZN( u1_u1_u1_n175 ) );
  NAND2_X1 u1_u1_u1_U55 (.A1( u1_u1_u1_n100 ) , .ZN( u1_u1_u1_n116 ) , .A2( u1_u1_u1_n95 ) );
  NAND2_X1 u1_u1_u1_U56 (.A1( u1_u1_u1_n102 ) , .ZN( u1_u1_u1_n131 ) , .A2( u1_u1_u1_n95 ) );
  NAND2_X1 u1_u1_u1_U57 (.A2( u1_u1_u1_n104 ) , .ZN( u1_u1_u1_n121 ) , .A1( u1_u1_u1_n98 ) );
  NAND2_X1 u1_u1_u1_U58 (.A1( u1_u1_u1_n103 ) , .ZN( u1_u1_u1_n153 ) , .A2( u1_u1_u1_n98 ) );
  NAND2_X1 u1_u1_u1_U59 (.A2( u1_u1_u1_n104 ) , .A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n133 ) );
  AOI22_X1 u1_u1_u1_U6 (.B2( u1_u1_u1_n113 ) , .A2( u1_u1_u1_n114 ) , .ZN( u1_u1_u1_n125 ) , .A1( u1_u1_u1_n171 ) , .B1( u1_u1_u1_n173 ) );
  NAND2_X1 u1_u1_u1_U60 (.ZN( u1_u1_u1_n150 ) , .A2( u1_u1_u1_n98 ) , .A1( u1_u1_u1_n99 ) );
  NAND2_X1 u1_u1_u1_U61 (.A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n155 ) , .A2( u1_u1_u1_n95 ) );
  OAI21_X1 u1_u1_u1_U62 (.ZN( u1_u1_u1_n109 ) , .B1( u1_u1_u1_n129 ) , .B2( u1_u1_u1_n160 ) , .A( u1_u1_u1_n167 ) );
  NAND2_X1 u1_u1_u1_U63 (.A2( u1_u1_u1_n100 ) , .A1( u1_u1_u1_n103 ) , .ZN( u1_u1_u1_n120 ) );
  NAND2_X1 u1_u1_u1_U64 (.A1( u1_u1_u1_n102 ) , .A2( u1_u1_u1_n104 ) , .ZN( u1_u1_u1_n115 ) );
  NAND2_X1 u1_u1_u1_U65 (.A2( u1_u1_u1_n100 ) , .A1( u1_u1_u1_n104 ) , .ZN( u1_u1_u1_n151 ) );
  NAND2_X1 u1_u1_u1_U66 (.A2( u1_u1_u1_n103 ) , .A1( u1_u1_u1_n105 ) , .ZN( u1_u1_u1_n161 ) );
  INV_X1 u1_u1_u1_U67 (.A( u1_u1_u1_n152 ) , .ZN( u1_u1_u1_n173 ) );
  INV_X1 u1_u1_u1_U68 (.A( u1_u1_u1_n128 ) , .ZN( u1_u1_u1_n172 ) );
  NAND2_X1 u1_u1_u1_U69 (.A2( u1_u1_u1_n102 ) , .A1( u1_u1_u1_n103 ) , .ZN( u1_u1_u1_n123 ) );
  NAND2_X1 u1_u1_u1_U7 (.ZN( u1_u1_u1_n114 ) , .A1( u1_u1_u1_n134 ) , .A2( u1_u1_u1_n156 ) );
  NOR2_X1 u1_u1_u1_U70 (.A2( u1_u1_X_7 ) , .A1( u1_u1_X_8 ) , .ZN( u1_u1_u1_n95 ) );
  NOR2_X1 u1_u1_u1_U71 (.A1( u1_u1_X_12 ) , .A2( u1_u1_X_9 ) , .ZN( u1_u1_u1_n100 ) );
  NOR2_X1 u1_u1_u1_U72 (.A2( u1_u1_X_8 ) , .A1( u1_u1_u1_n177 ) , .ZN( u1_u1_u1_n99 ) );
  NOR2_X1 u1_u1_u1_U73 (.A2( u1_u1_X_12 ) , .ZN( u1_u1_u1_n102 ) , .A1( u1_u1_u1_n176 ) );
  NOR2_X1 u1_u1_u1_U74 (.A2( u1_u1_X_9 ) , .ZN( u1_u1_u1_n105 ) , .A1( u1_u1_u1_n168 ) );
  NAND2_X1 u1_u1_u1_U75 (.A1( u1_u1_X_10 ) , .ZN( u1_u1_u1_n160 ) , .A2( u1_u1_u1_n169 ) );
  NAND2_X1 u1_u1_u1_U76 (.A2( u1_u1_X_10 ) , .A1( u1_u1_X_11 ) , .ZN( u1_u1_u1_n152 ) );
  NAND2_X1 u1_u1_u1_U77 (.A1( u1_u1_X_11 ) , .ZN( u1_u1_u1_n128 ) , .A2( u1_u1_u1_n170 ) );
  AND2_X1 u1_u1_u1_U78 (.A2( u1_u1_X_7 ) , .A1( u1_u1_X_8 ) , .ZN( u1_u1_u1_n104 ) );
  AND2_X1 u1_u1_u1_U79 (.A1( u1_u1_X_8 ) , .ZN( u1_u1_u1_n103 ) , .A2( u1_u1_u1_n177 ) );
  AOI22_X1 u1_u1_u1_U8 (.B2( u1_u1_u1_n136 ) , .A2( u1_u1_u1_n137 ) , .ZN( u1_u1_u1_n143 ) , .A1( u1_u1_u1_n171 ) , .B1( u1_u1_u1_n173 ) );
  INV_X1 u1_u1_u1_U80 (.A( u1_u1_X_10 ) , .ZN( u1_u1_u1_n170 ) );
  INV_X1 u1_u1_u1_U81 (.A( u1_u1_X_9 ) , .ZN( u1_u1_u1_n176 ) );
  INV_X1 u1_u1_u1_U82 (.A( u1_u1_X_11 ) , .ZN( u1_u1_u1_n169 ) );
  INV_X1 u1_u1_u1_U83 (.A( u1_u1_X_12 ) , .ZN( u1_u1_u1_n168 ) );
  INV_X1 u1_u1_u1_U84 (.A( u1_u1_X_7 ) , .ZN( u1_u1_u1_n177 ) );
  NAND4_X1 u1_u1_u1_U85 (.ZN( u1_out1_28 ) , .A4( u1_u1_u1_n124 ) , .A3( u1_u1_u1_n125 ) , .A2( u1_u1_u1_n126 ) , .A1( u1_u1_u1_n127 ) );
  OAI21_X1 u1_u1_u1_U86 (.ZN( u1_u1_u1_n127 ) , .B2( u1_u1_u1_n139 ) , .B1( u1_u1_u1_n175 ) , .A( u1_u1_u1_n183 ) );
  OAI21_X1 u1_u1_u1_U87 (.ZN( u1_u1_u1_n126 ) , .B2( u1_u1_u1_n140 ) , .A( u1_u1_u1_n146 ) , .B1( u1_u1_u1_n178 ) );
  NAND4_X1 u1_u1_u1_U88 (.ZN( u1_out1_18 ) , .A4( u1_u1_u1_n165 ) , .A3( u1_u1_u1_n166 ) , .A1( u1_u1_u1_n167 ) , .A2( u1_u1_u1_n186 ) );
  AOI22_X1 u1_u1_u1_U89 (.B2( u1_u1_u1_n146 ) , .B1( u1_u1_u1_n147 ) , .A2( u1_u1_u1_n148 ) , .ZN( u1_u1_u1_n166 ) , .A1( u1_u1_u1_n172 ) );
  INV_X1 u1_u1_u1_U9 (.A( u1_u1_u1_n147 ) , .ZN( u1_u1_u1_n181 ) );
  INV_X1 u1_u1_u1_U90 (.A( u1_u1_u1_n145 ) , .ZN( u1_u1_u1_n186 ) );
  NAND4_X1 u1_u1_u1_U91 (.ZN( u1_out1_2 ) , .A4( u1_u1_u1_n142 ) , .A3( u1_u1_u1_n143 ) , .A2( u1_u1_u1_n144 ) , .A1( u1_u1_u1_n179 ) );
  INV_X1 u1_u1_u1_U92 (.A( u1_u1_u1_n130 ) , .ZN( u1_u1_u1_n179 ) );
  OAI21_X1 u1_u1_u1_U93 (.B2( u1_u1_u1_n132 ) , .ZN( u1_u1_u1_n144 ) , .A( u1_u1_u1_n146 ) , .B1( u1_u1_u1_n180 ) );
  OR4_X1 u1_u1_u1_U94 (.ZN( u1_out1_13 ) , .A4( u1_u1_u1_n108 ) , .A3( u1_u1_u1_n109 ) , .A2( u1_u1_u1_n110 ) , .A1( u1_u1_u1_n111 ) );
  AOI21_X1 u1_u1_u1_U95 (.ZN( u1_u1_u1_n111 ) , .A( u1_u1_u1_n128 ) , .B2( u1_u1_u1_n131 ) , .B1( u1_u1_u1_n135 ) );
  AOI21_X1 u1_u1_u1_U96 (.ZN( u1_u1_u1_n110 ) , .A( u1_u1_u1_n116 ) , .B1( u1_u1_u1_n152 ) , .B2( u1_u1_u1_n160 ) );
  NAND3_X1 u1_u1_u1_U97 (.A3( u1_u1_u1_n149 ) , .A2( u1_u1_u1_n150 ) , .A1( u1_u1_u1_n151 ) , .ZN( u1_u1_u1_n164 ) );
  NAND3_X1 u1_u1_u1_U98 (.A3( u1_u1_u1_n134 ) , .A2( u1_u1_u1_n135 ) , .ZN( u1_u1_u1_n136 ) , .A1( u1_u1_u1_n151 ) );
  NAND3_X1 u1_u1_u1_U99 (.A1( u1_u1_u1_n133 ) , .ZN( u1_u1_u1_n137 ) , .A2( u1_u1_u1_n154 ) , .A3( u1_u1_u1_n181 ) );
  OAI22_X1 u1_u1_u2_U10 (.ZN( u1_u1_u2_n109 ) , .A2( u1_u1_u2_n113 ) , .B2( u1_u1_u2_n133 ) , .B1( u1_u1_u2_n167 ) , .A1( u1_u1_u2_n168 ) );
  NAND3_X1 u1_u1_u2_U100 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n104 ) , .A3( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n98 ) );
  OAI22_X1 u1_u1_u2_U11 (.B1( u1_u1_u2_n151 ) , .A2( u1_u1_u2_n152 ) , .A1( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n160 ) , .B2( u1_u1_u2_n168 ) );
  NOR3_X1 u1_u1_u2_U12 (.A1( u1_u1_u2_n150 ) , .ZN( u1_u1_u2_n151 ) , .A3( u1_u1_u2_n175 ) , .A2( u1_u1_u2_n188 ) );
  AOI21_X1 u1_u1_u2_U13 (.ZN( u1_u1_u2_n144 ) , .B2( u1_u1_u2_n155 ) , .A( u1_u1_u2_n172 ) , .B1( u1_u1_u2_n185 ) );
  AOI21_X1 u1_u1_u2_U14 (.B2( u1_u1_u2_n143 ) , .ZN( u1_u1_u2_n145 ) , .B1( u1_u1_u2_n152 ) , .A( u1_u1_u2_n171 ) );
  AOI21_X1 u1_u1_u2_U15 (.B2( u1_u1_u2_n120 ) , .B1( u1_u1_u2_n121 ) , .ZN( u1_u1_u2_n126 ) , .A( u1_u1_u2_n167 ) );
  INV_X1 u1_u1_u2_U16 (.A( u1_u1_u2_n156 ) , .ZN( u1_u1_u2_n171 ) );
  INV_X1 u1_u1_u2_U17 (.A( u1_u1_u2_n120 ) , .ZN( u1_u1_u2_n188 ) );
  NAND2_X1 u1_u1_u2_U18 (.A2( u1_u1_u2_n122 ) , .ZN( u1_u1_u2_n150 ) , .A1( u1_u1_u2_n152 ) );
  INV_X1 u1_u1_u2_U19 (.A( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n170 ) );
  INV_X1 u1_u1_u2_U20 (.A( u1_u1_u2_n137 ) , .ZN( u1_u1_u2_n173 ) );
  NAND2_X1 u1_u1_u2_U21 (.A1( u1_u1_u2_n132 ) , .A2( u1_u1_u2_n139 ) , .ZN( u1_u1_u2_n157 ) );
  INV_X1 u1_u1_u2_U22 (.A( u1_u1_u2_n113 ) , .ZN( u1_u1_u2_n178 ) );
  INV_X1 u1_u1_u2_U23 (.A( u1_u1_u2_n139 ) , .ZN( u1_u1_u2_n175 ) );
  INV_X1 u1_u1_u2_U24 (.A( u1_u1_u2_n155 ) , .ZN( u1_u1_u2_n181 ) );
  INV_X1 u1_u1_u2_U25 (.A( u1_u1_u2_n119 ) , .ZN( u1_u1_u2_n177 ) );
  INV_X1 u1_u1_u2_U26 (.A( u1_u1_u2_n116 ) , .ZN( u1_u1_u2_n180 ) );
  INV_X1 u1_u1_u2_U27 (.A( u1_u1_u2_n131 ) , .ZN( u1_u1_u2_n179 ) );
  INV_X1 u1_u1_u2_U28 (.A( u1_u1_u2_n154 ) , .ZN( u1_u1_u2_n176 ) );
  NAND2_X1 u1_u1_u2_U29 (.A2( u1_u1_u2_n116 ) , .A1( u1_u1_u2_n117 ) , .ZN( u1_u1_u2_n118 ) );
  NOR2_X1 u1_u1_u2_U3 (.ZN( u1_u1_u2_n121 ) , .A2( u1_u1_u2_n177 ) , .A1( u1_u1_u2_n180 ) );
  INV_X1 u1_u1_u2_U30 (.A( u1_u1_u2_n132 ) , .ZN( u1_u1_u2_n182 ) );
  INV_X1 u1_u1_u2_U31 (.A( u1_u1_u2_n158 ) , .ZN( u1_u1_u2_n183 ) );
  OAI21_X1 u1_u1_u2_U32 (.A( u1_u1_u2_n156 ) , .B1( u1_u1_u2_n157 ) , .ZN( u1_u1_u2_n158 ) , .B2( u1_u1_u2_n179 ) );
  NOR2_X1 u1_u1_u2_U33 (.ZN( u1_u1_u2_n156 ) , .A1( u1_u1_u2_n166 ) , .A2( u1_u1_u2_n169 ) );
  NOR2_X1 u1_u1_u2_U34 (.A2( u1_u1_u2_n114 ) , .ZN( u1_u1_u2_n137 ) , .A1( u1_u1_u2_n140 ) );
  NOR2_X1 u1_u1_u2_U35 (.A2( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n153 ) , .A1( u1_u1_u2_n156 ) );
  AOI211_X1 u1_u1_u2_U36 (.ZN( u1_u1_u2_n130 ) , .C1( u1_u1_u2_n138 ) , .C2( u1_u1_u2_n179 ) , .B( u1_u1_u2_n96 ) , .A( u1_u1_u2_n97 ) );
  OAI22_X1 u1_u1_u2_U37 (.B1( u1_u1_u2_n133 ) , .A2( u1_u1_u2_n137 ) , .A1( u1_u1_u2_n152 ) , .B2( u1_u1_u2_n168 ) , .ZN( u1_u1_u2_n97 ) );
  OAI221_X1 u1_u1_u2_U38 (.B1( u1_u1_u2_n113 ) , .C1( u1_u1_u2_n132 ) , .A( u1_u1_u2_n149 ) , .B2( u1_u1_u2_n171 ) , .C2( u1_u1_u2_n172 ) , .ZN( u1_u1_u2_n96 ) );
  OAI221_X1 u1_u1_u2_U39 (.A( u1_u1_u2_n115 ) , .C2( u1_u1_u2_n123 ) , .B2( u1_u1_u2_n143 ) , .B1( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n163 ) , .C1( u1_u1_u2_n168 ) );
  INV_X1 u1_u1_u2_U4 (.A( u1_u1_u2_n134 ) , .ZN( u1_u1_u2_n185 ) );
  OAI21_X1 u1_u1_u2_U40 (.A( u1_u1_u2_n114 ) , .ZN( u1_u1_u2_n115 ) , .B1( u1_u1_u2_n176 ) , .B2( u1_u1_u2_n178 ) );
  OAI221_X1 u1_u1_u2_U41 (.A( u1_u1_u2_n135 ) , .B2( u1_u1_u2_n136 ) , .B1( u1_u1_u2_n137 ) , .ZN( u1_u1_u2_n162 ) , .C2( u1_u1_u2_n167 ) , .C1( u1_u1_u2_n185 ) );
  AND3_X1 u1_u1_u2_U42 (.A3( u1_u1_u2_n131 ) , .A2( u1_u1_u2_n132 ) , .A1( u1_u1_u2_n133 ) , .ZN( u1_u1_u2_n136 ) );
  AOI22_X1 u1_u1_u2_U43 (.ZN( u1_u1_u2_n135 ) , .B1( u1_u1_u2_n140 ) , .A1( u1_u1_u2_n156 ) , .B2( u1_u1_u2_n180 ) , .A2( u1_u1_u2_n188 ) );
  AOI21_X1 u1_u1_u2_U44 (.ZN( u1_u1_u2_n149 ) , .B1( u1_u1_u2_n173 ) , .B2( u1_u1_u2_n188 ) , .A( u1_u1_u2_n95 ) );
  AND3_X1 u1_u1_u2_U45 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n104 ) , .A3( u1_u1_u2_n156 ) , .ZN( u1_u1_u2_n95 ) );
  OAI21_X1 u1_u1_u2_U46 (.A( u1_u1_u2_n101 ) , .B2( u1_u1_u2_n121 ) , .B1( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n164 ) );
  NAND2_X1 u1_u1_u2_U47 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n107 ) , .ZN( u1_u1_u2_n155 ) );
  NAND2_X1 u1_u1_u2_U48 (.A2( u1_u1_u2_n105 ) , .A1( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n143 ) );
  NAND2_X1 u1_u1_u2_U49 (.A1( u1_u1_u2_n104 ) , .A2( u1_u1_u2_n106 ) , .ZN( u1_u1_u2_n152 ) );
  INV_X1 u1_u1_u2_U5 (.A( u1_u1_u2_n150 ) , .ZN( u1_u1_u2_n184 ) );
  NAND2_X1 u1_u1_u2_U50 (.A1( u1_u1_u2_n100 ) , .A2( u1_u1_u2_n105 ) , .ZN( u1_u1_u2_n132 ) );
  INV_X1 u1_u1_u2_U51 (.A( u1_u1_u2_n140 ) , .ZN( u1_u1_u2_n168 ) );
  INV_X1 u1_u1_u2_U52 (.A( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n167 ) );
  OAI21_X1 u1_u1_u2_U53 (.A( u1_u1_u2_n141 ) , .B2( u1_u1_u2_n142 ) , .ZN( u1_u1_u2_n146 ) , .B1( u1_u1_u2_n153 ) );
  OAI21_X1 u1_u1_u2_U54 (.A( u1_u1_u2_n140 ) , .ZN( u1_u1_u2_n141 ) , .B1( u1_u1_u2_n176 ) , .B2( u1_u1_u2_n177 ) );
  NOR3_X1 u1_u1_u2_U55 (.ZN( u1_u1_u2_n142 ) , .A3( u1_u1_u2_n175 ) , .A2( u1_u1_u2_n178 ) , .A1( u1_u1_u2_n181 ) );
  NAND2_X1 u1_u1_u2_U56 (.A1( u1_u1_u2_n102 ) , .A2( u1_u1_u2_n106 ) , .ZN( u1_u1_u2_n113 ) );
  NAND2_X1 u1_u1_u2_U57 (.A1( u1_u1_u2_n106 ) , .A2( u1_u1_u2_n107 ) , .ZN( u1_u1_u2_n131 ) );
  NAND2_X1 u1_u1_u2_U58 (.A1( u1_u1_u2_n103 ) , .A2( u1_u1_u2_n107 ) , .ZN( u1_u1_u2_n139 ) );
  NAND2_X1 u1_u1_u2_U59 (.A1( u1_u1_u2_n103 ) , .A2( u1_u1_u2_n105 ) , .ZN( u1_u1_u2_n133 ) );
  NOR4_X1 u1_u1_u2_U6 (.A4( u1_u1_u2_n124 ) , .A3( u1_u1_u2_n125 ) , .A2( u1_u1_u2_n126 ) , .A1( u1_u1_u2_n127 ) , .ZN( u1_u1_u2_n128 ) );
  NAND2_X1 u1_u1_u2_U60 (.A1( u1_u1_u2_n102 ) , .A2( u1_u1_u2_n103 ) , .ZN( u1_u1_u2_n154 ) );
  NAND2_X1 u1_u1_u2_U61 (.A2( u1_u1_u2_n103 ) , .A1( u1_u1_u2_n104 ) , .ZN( u1_u1_u2_n119 ) );
  NAND2_X1 u1_u1_u2_U62 (.A2( u1_u1_u2_n107 ) , .A1( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n123 ) );
  NAND2_X1 u1_u1_u2_U63 (.A1( u1_u1_u2_n104 ) , .A2( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n122 ) );
  INV_X1 u1_u1_u2_U64 (.A( u1_u1_u2_n114 ) , .ZN( u1_u1_u2_n172 ) );
  NAND2_X1 u1_u1_u2_U65 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n102 ) , .ZN( u1_u1_u2_n116 ) );
  NAND2_X1 u1_u1_u2_U66 (.A1( u1_u1_u2_n102 ) , .A2( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n120 ) );
  NAND2_X1 u1_u1_u2_U67 (.A2( u1_u1_u2_n105 ) , .A1( u1_u1_u2_n106 ) , .ZN( u1_u1_u2_n117 ) );
  INV_X1 u1_u1_u2_U68 (.ZN( u1_u1_u2_n187 ) , .A( u1_u1_u2_n99 ) );
  OAI21_X1 u1_u1_u2_U69 (.B1( u1_u1_u2_n137 ) , .B2( u1_u1_u2_n143 ) , .A( u1_u1_u2_n98 ) , .ZN( u1_u1_u2_n99 ) );
  AOI21_X1 u1_u1_u2_U7 (.B2( u1_u1_u2_n119 ) , .ZN( u1_u1_u2_n127 ) , .A( u1_u1_u2_n137 ) , .B1( u1_u1_u2_n155 ) );
  NOR2_X1 u1_u1_u2_U70 (.A2( u1_u1_X_16 ) , .ZN( u1_u1_u2_n140 ) , .A1( u1_u1_u2_n166 ) );
  NOR2_X1 u1_u1_u2_U71 (.A2( u1_u1_X_13 ) , .A1( u1_u1_X_14 ) , .ZN( u1_u1_u2_n100 ) );
  NOR2_X1 u1_u1_u2_U72 (.A2( u1_u1_X_16 ) , .A1( u1_u1_X_17 ) , .ZN( u1_u1_u2_n138 ) );
  NOR2_X1 u1_u1_u2_U73 (.A2( u1_u1_X_15 ) , .A1( u1_u1_X_18 ) , .ZN( u1_u1_u2_n104 ) );
  NOR2_X1 u1_u1_u2_U74 (.A2( u1_u1_X_14 ) , .ZN( u1_u1_u2_n103 ) , .A1( u1_u1_u2_n174 ) );
  NOR2_X1 u1_u1_u2_U75 (.A2( u1_u1_X_15 ) , .ZN( u1_u1_u2_n102 ) , .A1( u1_u1_u2_n165 ) );
  NOR2_X1 u1_u1_u2_U76 (.A2( u1_u1_X_17 ) , .ZN( u1_u1_u2_n114 ) , .A1( u1_u1_u2_n169 ) );
  AND2_X1 u1_u1_u2_U77 (.A1( u1_u1_X_15 ) , .ZN( u1_u1_u2_n105 ) , .A2( u1_u1_u2_n165 ) );
  AND2_X1 u1_u1_u2_U78 (.A2( u1_u1_X_15 ) , .A1( u1_u1_X_18 ) , .ZN( u1_u1_u2_n107 ) );
  AND2_X1 u1_u1_u2_U79 (.A1( u1_u1_X_14 ) , .ZN( u1_u1_u2_n106 ) , .A2( u1_u1_u2_n174 ) );
  AOI21_X1 u1_u1_u2_U8 (.ZN( u1_u1_u2_n124 ) , .B1( u1_u1_u2_n131 ) , .B2( u1_u1_u2_n143 ) , .A( u1_u1_u2_n172 ) );
  AND2_X1 u1_u1_u2_U80 (.A1( u1_u1_X_13 ) , .A2( u1_u1_X_14 ) , .ZN( u1_u1_u2_n108 ) );
  INV_X1 u1_u1_u2_U81 (.A( u1_u1_X_16 ) , .ZN( u1_u1_u2_n169 ) );
  INV_X1 u1_u1_u2_U82 (.A( u1_u1_X_17 ) , .ZN( u1_u1_u2_n166 ) );
  INV_X1 u1_u1_u2_U83 (.A( u1_u1_X_13 ) , .ZN( u1_u1_u2_n174 ) );
  INV_X1 u1_u1_u2_U84 (.A( u1_u1_X_18 ) , .ZN( u1_u1_u2_n165 ) );
  NAND4_X1 u1_u1_u2_U85 (.ZN( u1_out1_30 ) , .A4( u1_u1_u2_n147 ) , .A3( u1_u1_u2_n148 ) , .A2( u1_u1_u2_n149 ) , .A1( u1_u1_u2_n187 ) );
  NOR3_X1 u1_u1_u2_U86 (.A3( u1_u1_u2_n144 ) , .A2( u1_u1_u2_n145 ) , .A1( u1_u1_u2_n146 ) , .ZN( u1_u1_u2_n147 ) );
  AOI21_X1 u1_u1_u2_U87 (.B2( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n148 ) , .A( u1_u1_u2_n162 ) , .B1( u1_u1_u2_n182 ) );
  NAND4_X1 u1_u1_u2_U88 (.ZN( u1_out1_24 ) , .A4( u1_u1_u2_n111 ) , .A3( u1_u1_u2_n112 ) , .A1( u1_u1_u2_n130 ) , .A2( u1_u1_u2_n187 ) );
  AOI221_X1 u1_u1_u2_U89 (.A( u1_u1_u2_n109 ) , .B1( u1_u1_u2_n110 ) , .ZN( u1_u1_u2_n111 ) , .C1( u1_u1_u2_n134 ) , .C2( u1_u1_u2_n170 ) , .B2( u1_u1_u2_n173 ) );
  AOI21_X1 u1_u1_u2_U9 (.B2( u1_u1_u2_n123 ) , .ZN( u1_u1_u2_n125 ) , .A( u1_u1_u2_n171 ) , .B1( u1_u1_u2_n184 ) );
  AOI21_X1 u1_u1_u2_U90 (.ZN( u1_u1_u2_n112 ) , .B2( u1_u1_u2_n156 ) , .A( u1_u1_u2_n164 ) , .B1( u1_u1_u2_n181 ) );
  NAND4_X1 u1_u1_u2_U91 (.ZN( u1_out1_16 ) , .A4( u1_u1_u2_n128 ) , .A3( u1_u1_u2_n129 ) , .A1( u1_u1_u2_n130 ) , .A2( u1_u1_u2_n186 ) );
  AOI22_X1 u1_u1_u2_U92 (.A2( u1_u1_u2_n118 ) , .ZN( u1_u1_u2_n129 ) , .A1( u1_u1_u2_n140 ) , .B1( u1_u1_u2_n157 ) , .B2( u1_u1_u2_n170 ) );
  INV_X1 u1_u1_u2_U93 (.A( u1_u1_u2_n163 ) , .ZN( u1_u1_u2_n186 ) );
  OR4_X1 u1_u1_u2_U94 (.ZN( u1_out1_6 ) , .A4( u1_u1_u2_n161 ) , .A3( u1_u1_u2_n162 ) , .A2( u1_u1_u2_n163 ) , .A1( u1_u1_u2_n164 ) );
  OR3_X1 u1_u1_u2_U95 (.A2( u1_u1_u2_n159 ) , .A1( u1_u1_u2_n160 ) , .ZN( u1_u1_u2_n161 ) , .A3( u1_u1_u2_n183 ) );
  AOI21_X1 u1_u1_u2_U96 (.B2( u1_u1_u2_n154 ) , .B1( u1_u1_u2_n155 ) , .ZN( u1_u1_u2_n159 ) , .A( u1_u1_u2_n167 ) );
  NAND3_X1 u1_u1_u2_U97 (.A2( u1_u1_u2_n117 ) , .A1( u1_u1_u2_n122 ) , .A3( u1_u1_u2_n123 ) , .ZN( u1_u1_u2_n134 ) );
  NAND3_X1 u1_u1_u2_U98 (.ZN( u1_u1_u2_n110 ) , .A2( u1_u1_u2_n131 ) , .A3( u1_u1_u2_n139 ) , .A1( u1_u1_u2_n154 ) );
  NAND3_X1 u1_u1_u2_U99 (.A2( u1_u1_u2_n100 ) , .ZN( u1_u1_u2_n101 ) , .A1( u1_u1_u2_n104 ) , .A3( u1_u1_u2_n114 ) );
  XOR2_X1 u1_u4_U1 (.B( u1_K5_9 ) , .A( u1_R3_6 ) , .Z( u1_u4_X_9 ) );
  XOR2_X1 u1_u4_U2 (.B( u1_K5_8 ) , .A( u1_R3_5 ) , .Z( u1_u4_X_8 ) );
  XOR2_X1 u1_u4_U3 (.B( u1_K5_7 ) , .A( u1_R3_4 ) , .Z( u1_u4_X_7 ) );
  XOR2_X1 u1_u4_U46 (.B( u1_K5_12 ) , .A( u1_R3_9 ) , .Z( u1_u4_X_12 ) );
  XOR2_X1 u1_u4_U47 (.B( u1_K5_11 ) , .A( u1_R3_8 ) , .Z( u1_u4_X_11 ) );
  XOR2_X1 u1_u4_U48 (.B( u1_K5_10 ) , .A( u1_R3_7 ) , .Z( u1_u4_X_10 ) );
  NOR2_X1 u1_u4_u1_U10 (.A1( u1_u4_u1_n112 ) , .A2( u1_u4_u1_n116 ) , .ZN( u1_u4_u1_n118 ) );
  NAND3_X1 u1_u4_u1_U100 (.ZN( u1_u4_u1_n113 ) , .A1( u1_u4_u1_n120 ) , .A3( u1_u4_u1_n133 ) , .A2( u1_u4_u1_n155 ) );
  OAI21_X1 u1_u4_u1_U11 (.ZN( u1_u4_u1_n101 ) , .B1( u1_u4_u1_n141 ) , .A( u1_u4_u1_n146 ) , .B2( u1_u4_u1_n183 ) );
  AOI21_X1 u1_u4_u1_U12 (.B2( u1_u4_u1_n155 ) , .B1( u1_u4_u1_n156 ) , .ZN( u1_u4_u1_n157 ) , .A( u1_u4_u1_n174 ) );
  NAND2_X1 u1_u4_u1_U13 (.ZN( u1_u4_u1_n140 ) , .A2( u1_u4_u1_n150 ) , .A1( u1_u4_u1_n155 ) );
  NAND2_X1 u1_u4_u1_U14 (.A1( u1_u4_u1_n131 ) , .ZN( u1_u4_u1_n147 ) , .A2( u1_u4_u1_n153 ) );
  INV_X1 u1_u4_u1_U15 (.A( u1_u4_u1_n139 ) , .ZN( u1_u4_u1_n174 ) );
  OR4_X1 u1_u4_u1_U16 (.A4( u1_u4_u1_n106 ) , .A3( u1_u4_u1_n107 ) , .ZN( u1_u4_u1_n108 ) , .A1( u1_u4_u1_n117 ) , .A2( u1_u4_u1_n184 ) );
  AOI21_X1 u1_u4_u1_U17 (.ZN( u1_u4_u1_n106 ) , .A( u1_u4_u1_n112 ) , .B1( u1_u4_u1_n154 ) , .B2( u1_u4_u1_n156 ) );
  AOI21_X1 u1_u4_u1_U18 (.ZN( u1_u4_u1_n107 ) , .B1( u1_u4_u1_n134 ) , .B2( u1_u4_u1_n149 ) , .A( u1_u4_u1_n174 ) );
  INV_X1 u1_u4_u1_U19 (.A( u1_u4_u1_n101 ) , .ZN( u1_u4_u1_n184 ) );
  INV_X1 u1_u4_u1_U20 (.A( u1_u4_u1_n112 ) , .ZN( u1_u4_u1_n171 ) );
  NAND2_X1 u1_u4_u1_U21 (.ZN( u1_u4_u1_n141 ) , .A1( u1_u4_u1_n153 ) , .A2( u1_u4_u1_n156 ) );
  AND2_X1 u1_u4_u1_U22 (.A1( u1_u4_u1_n123 ) , .ZN( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n161 ) );
  NAND2_X1 u1_u4_u1_U23 (.A2( u1_u4_u1_n115 ) , .A1( u1_u4_u1_n116 ) , .ZN( u1_u4_u1_n148 ) );
  NAND2_X1 u1_u4_u1_U24 (.A2( u1_u4_u1_n133 ) , .A1( u1_u4_u1_n135 ) , .ZN( u1_u4_u1_n159 ) );
  NAND2_X1 u1_u4_u1_U25 (.A2( u1_u4_u1_n115 ) , .A1( u1_u4_u1_n120 ) , .ZN( u1_u4_u1_n132 ) );
  INV_X1 u1_u4_u1_U26 (.A( u1_u4_u1_n154 ) , .ZN( u1_u4_u1_n178 ) );
  INV_X1 u1_u4_u1_U27 (.A( u1_u4_u1_n151 ) , .ZN( u1_u4_u1_n183 ) );
  AND2_X1 u1_u4_u1_U28 (.A1( u1_u4_u1_n129 ) , .A2( u1_u4_u1_n133 ) , .ZN( u1_u4_u1_n149 ) );
  INV_X1 u1_u4_u1_U29 (.A( u1_u4_u1_n131 ) , .ZN( u1_u4_u1_n180 ) );
  INV_X1 u1_u4_u1_U3 (.A( u1_u4_u1_n159 ) , .ZN( u1_u4_u1_n182 ) );
  OAI221_X1 u1_u4_u1_U30 (.A( u1_u4_u1_n119 ) , .C2( u1_u4_u1_n129 ) , .ZN( u1_u4_u1_n138 ) , .B2( u1_u4_u1_n152 ) , .C1( u1_u4_u1_n174 ) , .B1( u1_u4_u1_n187 ) );
  INV_X1 u1_u4_u1_U31 (.A( u1_u4_u1_n148 ) , .ZN( u1_u4_u1_n187 ) );
  AOI211_X1 u1_u4_u1_U32 (.B( u1_u4_u1_n117 ) , .A( u1_u4_u1_n118 ) , .ZN( u1_u4_u1_n119 ) , .C2( u1_u4_u1_n146 ) , .C1( u1_u4_u1_n159 ) );
  NOR2_X1 u1_u4_u1_U33 (.A1( u1_u4_u1_n168 ) , .A2( u1_u4_u1_n176 ) , .ZN( u1_u4_u1_n98 ) );
  AOI211_X1 u1_u4_u1_U34 (.B( u1_u4_u1_n162 ) , .A( u1_u4_u1_n163 ) , .C2( u1_u4_u1_n164 ) , .ZN( u1_u4_u1_n165 ) , .C1( u1_u4_u1_n171 ) );
  AOI21_X1 u1_u4_u1_U35 (.A( u1_u4_u1_n160 ) , .B2( u1_u4_u1_n161 ) , .ZN( u1_u4_u1_n162 ) , .B1( u1_u4_u1_n182 ) );
  OR2_X1 u1_u4_u1_U36 (.A2( u1_u4_u1_n157 ) , .A1( u1_u4_u1_n158 ) , .ZN( u1_u4_u1_n163 ) );
  NAND2_X1 u1_u4_u1_U37 (.A1( u1_u4_u1_n128 ) , .ZN( u1_u4_u1_n146 ) , .A2( u1_u4_u1_n160 ) );
  NAND2_X1 u1_u4_u1_U38 (.A2( u1_u4_u1_n112 ) , .ZN( u1_u4_u1_n139 ) , .A1( u1_u4_u1_n152 ) );
  NAND2_X1 u1_u4_u1_U39 (.A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n156 ) , .A2( u1_u4_u1_n99 ) );
  AOI221_X1 u1_u4_u1_U4 (.A( u1_u4_u1_n138 ) , .C2( u1_u4_u1_n139 ) , .C1( u1_u4_u1_n140 ) , .B2( u1_u4_u1_n141 ) , .ZN( u1_u4_u1_n142 ) , .B1( u1_u4_u1_n175 ) );
  AOI221_X1 u1_u4_u1_U40 (.B1( u1_u4_u1_n140 ) , .ZN( u1_u4_u1_n167 ) , .B2( u1_u4_u1_n172 ) , .C2( u1_u4_u1_n175 ) , .C1( u1_u4_u1_n178 ) , .A( u1_u4_u1_n188 ) );
  INV_X1 u1_u4_u1_U41 (.ZN( u1_u4_u1_n188 ) , .A( u1_u4_u1_n97 ) );
  AOI211_X1 u1_u4_u1_U42 (.A( u1_u4_u1_n118 ) , .C1( u1_u4_u1_n132 ) , .C2( u1_u4_u1_n139 ) , .B( u1_u4_u1_n96 ) , .ZN( u1_u4_u1_n97 ) );
  AOI21_X1 u1_u4_u1_U43 (.B2( u1_u4_u1_n121 ) , .B1( u1_u4_u1_n135 ) , .A( u1_u4_u1_n152 ) , .ZN( u1_u4_u1_n96 ) );
  NOR2_X1 u1_u4_u1_U44 (.ZN( u1_u4_u1_n117 ) , .A1( u1_u4_u1_n121 ) , .A2( u1_u4_u1_n160 ) );
  OAI21_X1 u1_u4_u1_U45 (.B2( u1_u4_u1_n123 ) , .ZN( u1_u4_u1_n145 ) , .B1( u1_u4_u1_n160 ) , .A( u1_u4_u1_n185 ) );
  INV_X1 u1_u4_u1_U46 (.A( u1_u4_u1_n122 ) , .ZN( u1_u4_u1_n185 ) );
  AOI21_X1 u1_u4_u1_U47 (.B2( u1_u4_u1_n120 ) , .B1( u1_u4_u1_n121 ) , .ZN( u1_u4_u1_n122 ) , .A( u1_u4_u1_n128 ) );
  AOI21_X1 u1_u4_u1_U48 (.A( u1_u4_u1_n128 ) , .B2( u1_u4_u1_n129 ) , .ZN( u1_u4_u1_n130 ) , .B1( u1_u4_u1_n150 ) );
  NAND2_X1 u1_u4_u1_U49 (.ZN( u1_u4_u1_n112 ) , .A1( u1_u4_u1_n169 ) , .A2( u1_u4_u1_n170 ) );
  AOI211_X1 u1_u4_u1_U5 (.ZN( u1_u4_u1_n124 ) , .A( u1_u4_u1_n138 ) , .C2( u1_u4_u1_n139 ) , .B( u1_u4_u1_n145 ) , .C1( u1_u4_u1_n147 ) );
  NAND2_X1 u1_u4_u1_U50 (.ZN( u1_u4_u1_n129 ) , .A2( u1_u4_u1_n95 ) , .A1( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U51 (.A1( u1_u4_u1_n102 ) , .ZN( u1_u4_u1_n154 ) , .A2( u1_u4_u1_n99 ) );
  NAND2_X1 u1_u4_u1_U52 (.A2( u1_u4_u1_n100 ) , .ZN( u1_u4_u1_n135 ) , .A1( u1_u4_u1_n99 ) );
  AOI21_X1 u1_u4_u1_U53 (.A( u1_u4_u1_n152 ) , .B2( u1_u4_u1_n153 ) , .B1( u1_u4_u1_n154 ) , .ZN( u1_u4_u1_n158 ) );
  INV_X1 u1_u4_u1_U54 (.A( u1_u4_u1_n160 ) , .ZN( u1_u4_u1_n175 ) );
  NAND2_X1 u1_u4_u1_U55 (.A1( u1_u4_u1_n100 ) , .ZN( u1_u4_u1_n116 ) , .A2( u1_u4_u1_n95 ) );
  NAND2_X1 u1_u4_u1_U56 (.A1( u1_u4_u1_n102 ) , .ZN( u1_u4_u1_n131 ) , .A2( u1_u4_u1_n95 ) );
  NAND2_X1 u1_u4_u1_U57 (.A2( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n121 ) , .A1( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U58 (.A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n153 ) , .A2( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U59 (.A2( u1_u4_u1_n104 ) , .A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n133 ) );
  AOI22_X1 u1_u4_u1_U6 (.B2( u1_u4_u1_n113 ) , .A2( u1_u4_u1_n114 ) , .ZN( u1_u4_u1_n125 ) , .A1( u1_u4_u1_n171 ) , .B1( u1_u4_u1_n173 ) );
  NAND2_X1 u1_u4_u1_U60 (.ZN( u1_u4_u1_n150 ) , .A2( u1_u4_u1_n98 ) , .A1( u1_u4_u1_n99 ) );
  NAND2_X1 u1_u4_u1_U61 (.A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n155 ) , .A2( u1_u4_u1_n95 ) );
  OAI21_X1 u1_u4_u1_U62 (.ZN( u1_u4_u1_n109 ) , .B1( u1_u4_u1_n129 ) , .B2( u1_u4_u1_n160 ) , .A( u1_u4_u1_n167 ) );
  NAND2_X1 u1_u4_u1_U63 (.A2( u1_u4_u1_n100 ) , .A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n120 ) );
  NAND2_X1 u1_u4_u1_U64 (.A1( u1_u4_u1_n102 ) , .A2( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n115 ) );
  NAND2_X1 u1_u4_u1_U65 (.A2( u1_u4_u1_n100 ) , .A1( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n151 ) );
  NAND2_X1 u1_u4_u1_U66 (.A2( u1_u4_u1_n103 ) , .A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n161 ) );
  INV_X1 u1_u4_u1_U67 (.A( u1_u4_u1_n152 ) , .ZN( u1_u4_u1_n173 ) );
  INV_X1 u1_u4_u1_U68 (.A( u1_u4_u1_n128 ) , .ZN( u1_u4_u1_n172 ) );
  NAND2_X1 u1_u4_u1_U69 (.A2( u1_u4_u1_n102 ) , .A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n123 ) );
  NAND2_X1 u1_u4_u1_U7 (.ZN( u1_u4_u1_n114 ) , .A1( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n156 ) );
  NOR2_X1 u1_u4_u1_U70 (.A2( u1_u4_X_7 ) , .A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n95 ) );
  NOR2_X1 u1_u4_u1_U71 (.A1( u1_u4_X_12 ) , .A2( u1_u4_X_9 ) , .ZN( u1_u4_u1_n100 ) );
  NOR2_X1 u1_u4_u1_U72 (.A2( u1_u4_X_8 ) , .A1( u1_u4_u1_n177 ) , .ZN( u1_u4_u1_n99 ) );
  NOR2_X1 u1_u4_u1_U73 (.A2( u1_u4_X_12 ) , .ZN( u1_u4_u1_n102 ) , .A1( u1_u4_u1_n176 ) );
  NOR2_X1 u1_u4_u1_U74 (.A2( u1_u4_X_9 ) , .ZN( u1_u4_u1_n105 ) , .A1( u1_u4_u1_n168 ) );
  NAND2_X1 u1_u4_u1_U75 (.A1( u1_u4_X_10 ) , .ZN( u1_u4_u1_n160 ) , .A2( u1_u4_u1_n169 ) );
  NAND2_X1 u1_u4_u1_U76 (.A2( u1_u4_X_10 ) , .A1( u1_u4_X_11 ) , .ZN( u1_u4_u1_n152 ) );
  NAND2_X1 u1_u4_u1_U77 (.A1( u1_u4_X_11 ) , .ZN( u1_u4_u1_n128 ) , .A2( u1_u4_u1_n170 ) );
  AND2_X1 u1_u4_u1_U78 (.A2( u1_u4_X_7 ) , .A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n104 ) );
  AND2_X1 u1_u4_u1_U79 (.A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n103 ) , .A2( u1_u4_u1_n177 ) );
  AOI22_X1 u1_u4_u1_U8 (.B2( u1_u4_u1_n136 ) , .A2( u1_u4_u1_n137 ) , .ZN( u1_u4_u1_n143 ) , .A1( u1_u4_u1_n171 ) , .B1( u1_u4_u1_n173 ) );
  INV_X1 u1_u4_u1_U80 (.A( u1_u4_X_10 ) , .ZN( u1_u4_u1_n170 ) );
  INV_X1 u1_u4_u1_U81 (.A( u1_u4_X_9 ) , .ZN( u1_u4_u1_n176 ) );
  INV_X1 u1_u4_u1_U82 (.A( u1_u4_X_11 ) , .ZN( u1_u4_u1_n169 ) );
  INV_X1 u1_u4_u1_U83 (.A( u1_u4_X_12 ) , .ZN( u1_u4_u1_n168 ) );
  INV_X1 u1_u4_u1_U84 (.A( u1_u4_X_7 ) , .ZN( u1_u4_u1_n177 ) );
  NAND4_X1 u1_u4_u1_U85 (.ZN( u1_out4_18 ) , .A4( u1_u4_u1_n165 ) , .A3( u1_u4_u1_n166 ) , .A1( u1_u4_u1_n167 ) , .A2( u1_u4_u1_n186 ) );
  AOI22_X1 u1_u4_u1_U86 (.B2( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n147 ) , .A2( u1_u4_u1_n148 ) , .ZN( u1_u4_u1_n166 ) , .A1( u1_u4_u1_n172 ) );
  INV_X1 u1_u4_u1_U87 (.A( u1_u4_u1_n145 ) , .ZN( u1_u4_u1_n186 ) );
  NAND4_X1 u1_u4_u1_U88 (.ZN( u1_out4_2 ) , .A4( u1_u4_u1_n142 ) , .A3( u1_u4_u1_n143 ) , .A2( u1_u4_u1_n144 ) , .A1( u1_u4_u1_n179 ) );
  OAI21_X1 u1_u4_u1_U89 (.B2( u1_u4_u1_n132 ) , .ZN( u1_u4_u1_n144 ) , .A( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n180 ) );
  INV_X1 u1_u4_u1_U9 (.A( u1_u4_u1_n147 ) , .ZN( u1_u4_u1_n181 ) );
  INV_X1 u1_u4_u1_U90 (.A( u1_u4_u1_n130 ) , .ZN( u1_u4_u1_n179 ) );
  NAND4_X1 u1_u4_u1_U91 (.ZN( u1_out4_28 ) , .A4( u1_u4_u1_n124 ) , .A3( u1_u4_u1_n125 ) , .A2( u1_u4_u1_n126 ) , .A1( u1_u4_u1_n127 ) );
  OAI21_X1 u1_u4_u1_U92 (.ZN( u1_u4_u1_n127 ) , .B2( u1_u4_u1_n139 ) , .B1( u1_u4_u1_n175 ) , .A( u1_u4_u1_n183 ) );
  OAI21_X1 u1_u4_u1_U93 (.ZN( u1_u4_u1_n126 ) , .B2( u1_u4_u1_n140 ) , .A( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n178 ) );
  OR4_X1 u1_u4_u1_U94 (.ZN( u1_out4_13 ) , .A4( u1_u4_u1_n108 ) , .A3( u1_u4_u1_n109 ) , .A2( u1_u4_u1_n110 ) , .A1( u1_u4_u1_n111 ) );
  AOI21_X1 u1_u4_u1_U95 (.ZN( u1_u4_u1_n111 ) , .A( u1_u4_u1_n128 ) , .B2( u1_u4_u1_n131 ) , .B1( u1_u4_u1_n135 ) );
  AOI21_X1 u1_u4_u1_U96 (.ZN( u1_u4_u1_n110 ) , .A( u1_u4_u1_n116 ) , .B1( u1_u4_u1_n152 ) , .B2( u1_u4_u1_n160 ) );
  NAND3_X1 u1_u4_u1_U97 (.A3( u1_u4_u1_n149 ) , .A2( u1_u4_u1_n150 ) , .A1( u1_u4_u1_n151 ) , .ZN( u1_u4_u1_n164 ) );
  NAND3_X1 u1_u4_u1_U98 (.A3( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n135 ) , .ZN( u1_u4_u1_n136 ) , .A1( u1_u4_u1_n151 ) );
  NAND3_X1 u1_u4_u1_U99 (.A1( u1_u4_u1_n133 ) , .ZN( u1_u4_u1_n137 ) , .A2( u1_u4_u1_n154 ) , .A3( u1_u4_u1_n181 ) );
  XOR2_X1 u1_u9_U1 (.B( u1_K10_9 ) , .A( u1_R8_6 ) , .Z( u1_u9_X_9 ) );
  XOR2_X1 u1_u9_U16 (.B( u1_K10_3 ) , .A( u1_R8_2 ) , .Z( u1_u9_X_3 ) );
  XOR2_X1 u1_u9_U2 (.B( u1_K10_8 ) , .A( u1_R8_5 ) , .Z( u1_u9_X_8 ) );
  XOR2_X1 u1_u9_U27 (.B( u1_K10_2 ) , .A( u1_R8_1 ) , .Z( u1_u9_X_2 ) );
  XOR2_X1 u1_u9_U3 (.B( u1_K10_7 ) , .A( u1_R8_4 ) , .Z( u1_u9_X_7 ) );
  XOR2_X1 u1_u9_U38 (.B( u1_K10_1 ) , .A( u1_R8_32 ) , .Z( u1_u9_X_1 ) );
  XOR2_X1 u1_u9_U4 (.B( u1_K10_6 ) , .A( u1_R8_5 ) , .Z( u1_u9_X_6 ) );
  XOR2_X1 u1_u9_U40 (.B( u1_K10_18 ) , .A( u1_R8_13 ) , .Z( u1_u9_X_18 ) );
  XOR2_X1 u1_u9_U41 (.B( u1_K10_17 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_17 ) );
  XOR2_X1 u1_u9_U42 (.B( u1_K10_16 ) , .A( u1_R8_11 ) , .Z( u1_u9_X_16 ) );
  XOR2_X1 u1_u9_U43 (.B( u1_K10_15 ) , .A( u1_R8_10 ) , .Z( u1_u9_X_15 ) );
  XOR2_X1 u1_u9_U44 (.B( u1_K10_14 ) , .A( u1_R8_9 ) , .Z( u1_u9_X_14 ) );
  XOR2_X1 u1_u9_U45 (.B( u1_K10_13 ) , .A( u1_R8_8 ) , .Z( u1_u9_X_13 ) );
  XOR2_X1 u1_u9_U46 (.B( u1_K10_12 ) , .A( u1_R8_9 ) , .Z( u1_u9_X_12 ) );
  XOR2_X1 u1_u9_U47 (.B( u1_K10_11 ) , .A( u1_R8_8 ) , .Z( u1_u9_X_11 ) );
  XOR2_X1 u1_u9_U48 (.B( u1_K10_10 ) , .A( u1_R8_7 ) , .Z( u1_u9_X_10 ) );
  XOR2_X1 u1_u9_U5 (.B( u1_K10_5 ) , .A( u1_R8_4 ) , .Z( u1_u9_X_5 ) );
  XOR2_X1 u1_u9_U6 (.B( u1_K10_4 ) , .A( u1_R8_3 ) , .Z( u1_u9_X_4 ) );
  AND3_X1 u1_u9_u0_U10 (.A2( u1_u9_u0_n112 ) , .ZN( u1_u9_u0_n127 ) , .A3( u1_u9_u0_n130 ) , .A1( u1_u9_u0_n148 ) );
  NAND2_X1 u1_u9_u0_U11 (.ZN( u1_u9_u0_n113 ) , .A1( u1_u9_u0_n139 ) , .A2( u1_u9_u0_n149 ) );
  AND2_X1 u1_u9_u0_U12 (.ZN( u1_u9_u0_n107 ) , .A1( u1_u9_u0_n130 ) , .A2( u1_u9_u0_n140 ) );
  AND2_X1 u1_u9_u0_U13 (.A2( u1_u9_u0_n129 ) , .A1( u1_u9_u0_n130 ) , .ZN( u1_u9_u0_n151 ) );
  AND2_X1 u1_u9_u0_U14 (.A1( u1_u9_u0_n108 ) , .A2( u1_u9_u0_n125 ) , .ZN( u1_u9_u0_n145 ) );
  INV_X1 u1_u9_u0_U15 (.A( u1_u9_u0_n143 ) , .ZN( u1_u9_u0_n173 ) );
  NOR2_X1 u1_u9_u0_U16 (.A2( u1_u9_u0_n136 ) , .ZN( u1_u9_u0_n147 ) , .A1( u1_u9_u0_n160 ) );
  AOI21_X1 u1_u9_u0_U17 (.B1( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n132 ) , .A( u1_u9_u0_n165 ) , .B2( u1_u9_u0_n93 ) );
  INV_X1 u1_u9_u0_U18 (.A( u1_u9_u0_n142 ) , .ZN( u1_u9_u0_n165 ) );
  OAI221_X1 u1_u9_u0_U19 (.C1( u1_u9_u0_n121 ) , .ZN( u1_u9_u0_n122 ) , .B2( u1_u9_u0_n127 ) , .A( u1_u9_u0_n143 ) , .B1( u1_u9_u0_n144 ) , .C2( u1_u9_u0_n147 ) );
  OAI22_X1 u1_u9_u0_U20 (.B1( u1_u9_u0_n131 ) , .A1( u1_u9_u0_n144 ) , .B2( u1_u9_u0_n147 ) , .A2( u1_u9_u0_n90 ) , .ZN( u1_u9_u0_n91 ) );
  AND3_X1 u1_u9_u0_U21 (.A3( u1_u9_u0_n121 ) , .A2( u1_u9_u0_n125 ) , .A1( u1_u9_u0_n148 ) , .ZN( u1_u9_u0_n90 ) );
  OAI22_X1 u1_u9_u0_U22 (.B1( u1_u9_u0_n125 ) , .ZN( u1_u9_u0_n126 ) , .A1( u1_u9_u0_n138 ) , .A2( u1_u9_u0_n146 ) , .B2( u1_u9_u0_n147 ) );
  NOR2_X1 u1_u9_u0_U23 (.A1( u1_u9_u0_n163 ) , .A2( u1_u9_u0_n164 ) , .ZN( u1_u9_u0_n95 ) );
  INV_X1 u1_u9_u0_U24 (.A( u1_u9_u0_n136 ) , .ZN( u1_u9_u0_n161 ) );
  NOR2_X1 u1_u9_u0_U25 (.A1( u1_u9_u0_n120 ) , .ZN( u1_u9_u0_n143 ) , .A2( u1_u9_u0_n167 ) );
  OAI221_X1 u1_u9_u0_U26 (.C1( u1_u9_u0_n112 ) , .ZN( u1_u9_u0_n120 ) , .B1( u1_u9_u0_n138 ) , .B2( u1_u9_u0_n141 ) , .C2( u1_u9_u0_n147 ) , .A( u1_u9_u0_n172 ) );
  AOI211_X1 u1_u9_u0_U27 (.B( u1_u9_u0_n115 ) , .A( u1_u9_u0_n116 ) , .C2( u1_u9_u0_n117 ) , .C1( u1_u9_u0_n118 ) , .ZN( u1_u9_u0_n119 ) );
  NAND2_X1 u1_u9_u0_U28 (.A1( u1_u9_u0_n101 ) , .A2( u1_u9_u0_n102 ) , .ZN( u1_u9_u0_n150 ) );
  AOI22_X1 u1_u9_u0_U29 (.B2( u1_u9_u0_n109 ) , .A2( u1_u9_u0_n110 ) , .ZN( u1_u9_u0_n111 ) , .B1( u1_u9_u0_n118 ) , .A1( u1_u9_u0_n160 ) );
  INV_X1 u1_u9_u0_U3 (.A( u1_u9_u0_n113 ) , .ZN( u1_u9_u0_n166 ) );
  INV_X1 u1_u9_u0_U30 (.A( u1_u9_u0_n118 ) , .ZN( u1_u9_u0_n158 ) );
  NAND2_X1 u1_u9_u0_U31 (.A2( u1_u9_u0_n100 ) , .A1( u1_u9_u0_n101 ) , .ZN( u1_u9_u0_n139 ) );
  NAND2_X1 u1_u9_u0_U32 (.A2( u1_u9_u0_n100 ) , .ZN( u1_u9_u0_n131 ) , .A1( u1_u9_u0_n92 ) );
  NAND2_X1 u1_u9_u0_U33 (.ZN( u1_u9_u0_n108 ) , .A1( u1_u9_u0_n92 ) , .A2( u1_u9_u0_n94 ) );
  AOI21_X1 u1_u9_u0_U34 (.ZN( u1_u9_u0_n104 ) , .B1( u1_u9_u0_n107 ) , .B2( u1_u9_u0_n141 ) , .A( u1_u9_u0_n144 ) );
  AOI21_X1 u1_u9_u0_U35 (.B1( u1_u9_u0_n127 ) , .B2( u1_u9_u0_n129 ) , .A( u1_u9_u0_n138 ) , .ZN( u1_u9_u0_n96 ) );
  NAND2_X1 u1_u9_u0_U36 (.A2( u1_u9_u0_n102 ) , .ZN( u1_u9_u0_n114 ) , .A1( u1_u9_u0_n92 ) );
  AOI21_X1 u1_u9_u0_U37 (.ZN( u1_u9_u0_n116 ) , .B2( u1_u9_u0_n142 ) , .A( u1_u9_u0_n144 ) , .B1( u1_u9_u0_n166 ) );
  NAND2_X1 u1_u9_u0_U38 (.A1( u1_u9_u0_n101 ) , .ZN( u1_u9_u0_n130 ) , .A2( u1_u9_u0_n94 ) );
  NAND2_X1 u1_u9_u0_U39 (.A1( u1_u9_u0_n100 ) , .A2( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n125 ) );
  AOI21_X1 u1_u9_u0_U4 (.B1( u1_u9_u0_n114 ) , .ZN( u1_u9_u0_n115 ) , .B2( u1_u9_u0_n129 ) , .A( u1_u9_u0_n161 ) );
  NAND2_X1 u1_u9_u0_U40 (.A2( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n140 ) , .A1( u1_u9_u0_n94 ) );
  INV_X1 u1_u9_u0_U41 (.A( u1_u9_u0_n138 ) , .ZN( u1_u9_u0_n160 ) );
  NAND2_X1 u1_u9_u0_U42 (.A2( u1_u9_u0_n102 ) , .A1( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n149 ) );
  NAND2_X1 u1_u9_u0_U43 (.A2( u1_u9_u0_n101 ) , .ZN( u1_u9_u0_n121 ) , .A1( u1_u9_u0_n93 ) );
  NAND2_X1 u1_u9_u0_U44 (.ZN( u1_u9_u0_n112 ) , .A2( u1_u9_u0_n92 ) , .A1( u1_u9_u0_n93 ) );
  INV_X1 u1_u9_u0_U45 (.ZN( u1_u9_u0_n172 ) , .A( u1_u9_u0_n88 ) );
  OAI222_X1 u1_u9_u0_U46 (.C1( u1_u9_u0_n108 ) , .A1( u1_u9_u0_n125 ) , .B2( u1_u9_u0_n128 ) , .B1( u1_u9_u0_n144 ) , .A2( u1_u9_u0_n158 ) , .C2( u1_u9_u0_n161 ) , .ZN( u1_u9_u0_n88 ) );
  OR3_X1 u1_u9_u0_U47 (.A3( u1_u9_u0_n152 ) , .A2( u1_u9_u0_n153 ) , .A1( u1_u9_u0_n154 ) , .ZN( u1_u9_u0_n155 ) );
  AOI21_X1 u1_u9_u0_U48 (.A( u1_u9_u0_n144 ) , .B2( u1_u9_u0_n145 ) , .B1( u1_u9_u0_n146 ) , .ZN( u1_u9_u0_n154 ) );
  AOI21_X1 u1_u9_u0_U49 (.B2( u1_u9_u0_n150 ) , .B1( u1_u9_u0_n151 ) , .ZN( u1_u9_u0_n152 ) , .A( u1_u9_u0_n158 ) );
  AOI21_X1 u1_u9_u0_U5 (.B2( u1_u9_u0_n131 ) , .ZN( u1_u9_u0_n134 ) , .B1( u1_u9_u0_n151 ) , .A( u1_u9_u0_n158 ) );
  AOI21_X1 u1_u9_u0_U50 (.A( u1_u9_u0_n147 ) , .B2( u1_u9_u0_n148 ) , .B1( u1_u9_u0_n149 ) , .ZN( u1_u9_u0_n153 ) );
  INV_X1 u1_u9_u0_U51 (.ZN( u1_u9_u0_n171 ) , .A( u1_u9_u0_n99 ) );
  OAI211_X1 u1_u9_u0_U52 (.C2( u1_u9_u0_n140 ) , .C1( u1_u9_u0_n161 ) , .A( u1_u9_u0_n169 ) , .B( u1_u9_u0_n98 ) , .ZN( u1_u9_u0_n99 ) );
  INV_X1 u1_u9_u0_U53 (.ZN( u1_u9_u0_n169 ) , .A( u1_u9_u0_n91 ) );
  AOI211_X1 u1_u9_u0_U54 (.C1( u1_u9_u0_n118 ) , .A( u1_u9_u0_n123 ) , .B( u1_u9_u0_n96 ) , .C2( u1_u9_u0_n97 ) , .ZN( u1_u9_u0_n98 ) );
  NOR2_X1 u1_u9_u0_U55 (.A2( u1_u9_X_2 ) , .ZN( u1_u9_u0_n103 ) , .A1( u1_u9_u0_n164 ) );
  NOR2_X1 u1_u9_u0_U56 (.A2( u1_u9_X_4 ) , .A1( u1_u9_X_5 ) , .ZN( u1_u9_u0_n118 ) );
  NOR2_X1 u1_u9_u0_U57 (.A2( u1_u9_X_3 ) , .A1( u1_u9_X_6 ) , .ZN( u1_u9_u0_n94 ) );
  NOR2_X1 u1_u9_u0_U58 (.A2( u1_u9_X_6 ) , .ZN( u1_u9_u0_n100 ) , .A1( u1_u9_u0_n162 ) );
  NAND2_X1 u1_u9_u0_U59 (.A2( u1_u9_X_4 ) , .A1( u1_u9_X_5 ) , .ZN( u1_u9_u0_n144 ) );
  NOR2_X1 u1_u9_u0_U6 (.A1( u1_u9_u0_n108 ) , .ZN( u1_u9_u0_n123 ) , .A2( u1_u9_u0_n158 ) );
  NOR2_X1 u1_u9_u0_U60 (.A2( u1_u9_X_5 ) , .ZN( u1_u9_u0_n136 ) , .A1( u1_u9_u0_n159 ) );
  NAND2_X1 u1_u9_u0_U61 (.A1( u1_u9_X_5 ) , .ZN( u1_u9_u0_n138 ) , .A2( u1_u9_u0_n159 ) );
  AND2_X1 u1_u9_u0_U62 (.A2( u1_u9_X_3 ) , .A1( u1_u9_X_6 ) , .ZN( u1_u9_u0_n102 ) );
  AND2_X1 u1_u9_u0_U63 (.A1( u1_u9_X_6 ) , .A2( u1_u9_u0_n162 ) , .ZN( u1_u9_u0_n93 ) );
  INV_X1 u1_u9_u0_U64 (.A( u1_u9_X_4 ) , .ZN( u1_u9_u0_n159 ) );
  INV_X1 u1_u9_u0_U65 (.A( u1_u9_X_3 ) , .ZN( u1_u9_u0_n162 ) );
  INV_X1 u1_u9_u0_U66 (.A( u1_u9_X_2 ) , .ZN( u1_u9_u0_n163 ) );
  INV_X1 u1_u9_u0_U67 (.A( u1_u9_u0_n126 ) , .ZN( u1_u9_u0_n168 ) );
  AOI211_X1 u1_u9_u0_U68 (.B( u1_u9_u0_n133 ) , .A( u1_u9_u0_n134 ) , .C2( u1_u9_u0_n135 ) , .C1( u1_u9_u0_n136 ) , .ZN( u1_u9_u0_n137 ) );
  INV_X1 u1_u9_u0_U69 (.ZN( u1_u9_u0_n174 ) , .A( u1_u9_u0_n89 ) );
  OAI21_X1 u1_u9_u0_U7 (.B1( u1_u9_u0_n150 ) , .B2( u1_u9_u0_n158 ) , .A( u1_u9_u0_n172 ) , .ZN( u1_u9_u0_n89 ) );
  AOI211_X1 u1_u9_u0_U70 (.B( u1_u9_u0_n104 ) , .A( u1_u9_u0_n105 ) , .ZN( u1_u9_u0_n106 ) , .C2( u1_u9_u0_n113 ) , .C1( u1_u9_u0_n160 ) );
  OR4_X1 u1_u9_u0_U71 (.ZN( u1_out9_17 ) , .A4( u1_u9_u0_n122 ) , .A2( u1_u9_u0_n123 ) , .A1( u1_u9_u0_n124 ) , .A3( u1_u9_u0_n170 ) );
  AOI21_X1 u1_u9_u0_U72 (.B2( u1_u9_u0_n107 ) , .ZN( u1_u9_u0_n124 ) , .B1( u1_u9_u0_n128 ) , .A( u1_u9_u0_n161 ) );
  INV_X1 u1_u9_u0_U73 (.A( u1_u9_u0_n111 ) , .ZN( u1_u9_u0_n170 ) );
  OR4_X1 u1_u9_u0_U74 (.ZN( u1_out9_31 ) , .A4( u1_u9_u0_n155 ) , .A2( u1_u9_u0_n156 ) , .A1( u1_u9_u0_n157 ) , .A3( u1_u9_u0_n173 ) );
  AOI21_X1 u1_u9_u0_U75 (.A( u1_u9_u0_n138 ) , .B2( u1_u9_u0_n139 ) , .B1( u1_u9_u0_n140 ) , .ZN( u1_u9_u0_n157 ) );
  AOI21_X1 u1_u9_u0_U76 (.B2( u1_u9_u0_n141 ) , .B1( u1_u9_u0_n142 ) , .ZN( u1_u9_u0_n156 ) , .A( u1_u9_u0_n161 ) );
  AOI21_X1 u1_u9_u0_U77 (.B1( u1_u9_u0_n132 ) , .ZN( u1_u9_u0_n133 ) , .A( u1_u9_u0_n144 ) , .B2( u1_u9_u0_n166 ) );
  OAI22_X1 u1_u9_u0_U78 (.ZN( u1_u9_u0_n105 ) , .A2( u1_u9_u0_n132 ) , .B1( u1_u9_u0_n146 ) , .A1( u1_u9_u0_n147 ) , .B2( u1_u9_u0_n161 ) );
  NAND2_X1 u1_u9_u0_U79 (.ZN( u1_u9_u0_n110 ) , .A2( u1_u9_u0_n132 ) , .A1( u1_u9_u0_n145 ) );
  AND2_X1 u1_u9_u0_U8 (.A1( u1_u9_u0_n114 ) , .A2( u1_u9_u0_n121 ) , .ZN( u1_u9_u0_n146 ) );
  INV_X1 u1_u9_u0_U80 (.A( u1_u9_u0_n119 ) , .ZN( u1_u9_u0_n167 ) );
  NAND2_X1 u1_u9_u0_U81 (.ZN( u1_u9_u0_n148 ) , .A1( u1_u9_u0_n93 ) , .A2( u1_u9_u0_n95 ) );
  NAND2_X1 u1_u9_u0_U82 (.A1( u1_u9_u0_n100 ) , .ZN( u1_u9_u0_n129 ) , .A2( u1_u9_u0_n95 ) );
  NAND2_X1 u1_u9_u0_U83 (.A1( u1_u9_u0_n102 ) , .ZN( u1_u9_u0_n128 ) , .A2( u1_u9_u0_n95 ) );
  NOR2_X1 u1_u9_u0_U84 (.A2( u1_u9_X_1 ) , .A1( u1_u9_X_2 ) , .ZN( u1_u9_u0_n92 ) );
  NAND2_X1 u1_u9_u0_U85 (.ZN( u1_u9_u0_n142 ) , .A1( u1_u9_u0_n94 ) , .A2( u1_u9_u0_n95 ) );
  NOR2_X1 u1_u9_u0_U86 (.A2( u1_u9_X_1 ) , .ZN( u1_u9_u0_n101 ) , .A1( u1_u9_u0_n163 ) );
  INV_X1 u1_u9_u0_U87 (.A( u1_u9_X_1 ) , .ZN( u1_u9_u0_n164 ) );
  NAND3_X1 u1_u9_u0_U88 (.ZN( u1_out9_23 ) , .A3( u1_u9_u0_n137 ) , .A1( u1_u9_u0_n168 ) , .A2( u1_u9_u0_n171 ) );
  NAND3_X1 u1_u9_u0_U89 (.A3( u1_u9_u0_n127 ) , .A2( u1_u9_u0_n128 ) , .ZN( u1_u9_u0_n135 ) , .A1( u1_u9_u0_n150 ) );
  AND2_X1 u1_u9_u0_U9 (.A1( u1_u9_u0_n131 ) , .ZN( u1_u9_u0_n141 ) , .A2( u1_u9_u0_n150 ) );
  NAND3_X1 u1_u9_u0_U90 (.ZN( u1_u9_u0_n117 ) , .A3( u1_u9_u0_n132 ) , .A2( u1_u9_u0_n139 ) , .A1( u1_u9_u0_n148 ) );
  NAND3_X1 u1_u9_u0_U91 (.ZN( u1_u9_u0_n109 ) , .A2( u1_u9_u0_n114 ) , .A3( u1_u9_u0_n140 ) , .A1( u1_u9_u0_n149 ) );
  NAND3_X1 u1_u9_u0_U92 (.ZN( u1_out9_9 ) , .A3( u1_u9_u0_n106 ) , .A2( u1_u9_u0_n171 ) , .A1( u1_u9_u0_n174 ) );
  NAND3_X1 u1_u9_u0_U93 (.A2( u1_u9_u0_n128 ) , .A1( u1_u9_u0_n132 ) , .A3( u1_u9_u0_n146 ) , .ZN( u1_u9_u0_n97 ) );
  NOR2_X1 u1_u9_u1_U10 (.A1( u1_u9_u1_n112 ) , .A2( u1_u9_u1_n116 ) , .ZN( u1_u9_u1_n118 ) );
  NAND3_X1 u1_u9_u1_U100 (.ZN( u1_u9_u1_n113 ) , .A1( u1_u9_u1_n120 ) , .A3( u1_u9_u1_n133 ) , .A2( u1_u9_u1_n155 ) );
  OAI21_X1 u1_u9_u1_U11 (.ZN( u1_u9_u1_n101 ) , .B1( u1_u9_u1_n141 ) , .A( u1_u9_u1_n146 ) , .B2( u1_u9_u1_n183 ) );
  AOI21_X1 u1_u9_u1_U12 (.B2( u1_u9_u1_n155 ) , .B1( u1_u9_u1_n156 ) , .ZN( u1_u9_u1_n157 ) , .A( u1_u9_u1_n174 ) );
  NAND2_X1 u1_u9_u1_U13 (.ZN( u1_u9_u1_n140 ) , .A2( u1_u9_u1_n150 ) , .A1( u1_u9_u1_n155 ) );
  NAND2_X1 u1_u9_u1_U14 (.A1( u1_u9_u1_n131 ) , .ZN( u1_u9_u1_n147 ) , .A2( u1_u9_u1_n153 ) );
  INV_X1 u1_u9_u1_U15 (.A( u1_u9_u1_n139 ) , .ZN( u1_u9_u1_n174 ) );
  OR4_X1 u1_u9_u1_U16 (.A4( u1_u9_u1_n106 ) , .A3( u1_u9_u1_n107 ) , .ZN( u1_u9_u1_n108 ) , .A1( u1_u9_u1_n117 ) , .A2( u1_u9_u1_n184 ) );
  AOI21_X1 u1_u9_u1_U17 (.ZN( u1_u9_u1_n106 ) , .A( u1_u9_u1_n112 ) , .B1( u1_u9_u1_n154 ) , .B2( u1_u9_u1_n156 ) );
  AOI21_X1 u1_u9_u1_U18 (.ZN( u1_u9_u1_n107 ) , .B1( u1_u9_u1_n134 ) , .B2( u1_u9_u1_n149 ) , .A( u1_u9_u1_n174 ) );
  INV_X1 u1_u9_u1_U19 (.A( u1_u9_u1_n101 ) , .ZN( u1_u9_u1_n184 ) );
  INV_X1 u1_u9_u1_U20 (.A( u1_u9_u1_n112 ) , .ZN( u1_u9_u1_n171 ) );
  NAND2_X1 u1_u9_u1_U21 (.ZN( u1_u9_u1_n141 ) , .A1( u1_u9_u1_n153 ) , .A2( u1_u9_u1_n156 ) );
  AND2_X1 u1_u9_u1_U22 (.A1( u1_u9_u1_n123 ) , .ZN( u1_u9_u1_n134 ) , .A2( u1_u9_u1_n161 ) );
  NAND2_X1 u1_u9_u1_U23 (.A2( u1_u9_u1_n115 ) , .A1( u1_u9_u1_n116 ) , .ZN( u1_u9_u1_n148 ) );
  NAND2_X1 u1_u9_u1_U24 (.A2( u1_u9_u1_n133 ) , .A1( u1_u9_u1_n135 ) , .ZN( u1_u9_u1_n159 ) );
  NAND2_X1 u1_u9_u1_U25 (.A2( u1_u9_u1_n115 ) , .A1( u1_u9_u1_n120 ) , .ZN( u1_u9_u1_n132 ) );
  INV_X1 u1_u9_u1_U26 (.A( u1_u9_u1_n154 ) , .ZN( u1_u9_u1_n178 ) );
  INV_X1 u1_u9_u1_U27 (.A( u1_u9_u1_n151 ) , .ZN( u1_u9_u1_n183 ) );
  AND2_X1 u1_u9_u1_U28 (.A1( u1_u9_u1_n129 ) , .A2( u1_u9_u1_n133 ) , .ZN( u1_u9_u1_n149 ) );
  INV_X1 u1_u9_u1_U29 (.A( u1_u9_u1_n131 ) , .ZN( u1_u9_u1_n180 ) );
  INV_X1 u1_u9_u1_U3 (.A( u1_u9_u1_n159 ) , .ZN( u1_u9_u1_n182 ) );
  OAI221_X1 u1_u9_u1_U30 (.A( u1_u9_u1_n119 ) , .C2( u1_u9_u1_n129 ) , .ZN( u1_u9_u1_n138 ) , .B2( u1_u9_u1_n152 ) , .C1( u1_u9_u1_n174 ) , .B1( u1_u9_u1_n187 ) );
  INV_X1 u1_u9_u1_U31 (.A( u1_u9_u1_n148 ) , .ZN( u1_u9_u1_n187 ) );
  AOI211_X1 u1_u9_u1_U32 (.B( u1_u9_u1_n117 ) , .A( u1_u9_u1_n118 ) , .ZN( u1_u9_u1_n119 ) , .C2( u1_u9_u1_n146 ) , .C1( u1_u9_u1_n159 ) );
  NOR2_X1 u1_u9_u1_U33 (.A1( u1_u9_u1_n168 ) , .A2( u1_u9_u1_n176 ) , .ZN( u1_u9_u1_n98 ) );
  AOI211_X1 u1_u9_u1_U34 (.B( u1_u9_u1_n162 ) , .A( u1_u9_u1_n163 ) , .C2( u1_u9_u1_n164 ) , .ZN( u1_u9_u1_n165 ) , .C1( u1_u9_u1_n171 ) );
  AOI21_X1 u1_u9_u1_U35 (.A( u1_u9_u1_n160 ) , .B2( u1_u9_u1_n161 ) , .ZN( u1_u9_u1_n162 ) , .B1( u1_u9_u1_n182 ) );
  OR2_X1 u1_u9_u1_U36 (.A2( u1_u9_u1_n157 ) , .A1( u1_u9_u1_n158 ) , .ZN( u1_u9_u1_n163 ) );
  NAND2_X1 u1_u9_u1_U37 (.A1( u1_u9_u1_n128 ) , .ZN( u1_u9_u1_n146 ) , .A2( u1_u9_u1_n160 ) );
  NAND2_X1 u1_u9_u1_U38 (.A2( u1_u9_u1_n112 ) , .ZN( u1_u9_u1_n139 ) , .A1( u1_u9_u1_n152 ) );
  NAND2_X1 u1_u9_u1_U39 (.A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n156 ) , .A2( u1_u9_u1_n99 ) );
  AOI221_X1 u1_u9_u1_U4 (.A( u1_u9_u1_n138 ) , .C2( u1_u9_u1_n139 ) , .C1( u1_u9_u1_n140 ) , .B2( u1_u9_u1_n141 ) , .ZN( u1_u9_u1_n142 ) , .B1( u1_u9_u1_n175 ) );
  AOI221_X1 u1_u9_u1_U40 (.B1( u1_u9_u1_n140 ) , .ZN( u1_u9_u1_n167 ) , .B2( u1_u9_u1_n172 ) , .C2( u1_u9_u1_n175 ) , .C1( u1_u9_u1_n178 ) , .A( u1_u9_u1_n188 ) );
  INV_X1 u1_u9_u1_U41 (.ZN( u1_u9_u1_n188 ) , .A( u1_u9_u1_n97 ) );
  AOI211_X1 u1_u9_u1_U42 (.A( u1_u9_u1_n118 ) , .C1( u1_u9_u1_n132 ) , .C2( u1_u9_u1_n139 ) , .B( u1_u9_u1_n96 ) , .ZN( u1_u9_u1_n97 ) );
  AOI21_X1 u1_u9_u1_U43 (.B2( u1_u9_u1_n121 ) , .B1( u1_u9_u1_n135 ) , .A( u1_u9_u1_n152 ) , .ZN( u1_u9_u1_n96 ) );
  NOR2_X1 u1_u9_u1_U44 (.ZN( u1_u9_u1_n117 ) , .A1( u1_u9_u1_n121 ) , .A2( u1_u9_u1_n160 ) );
  OAI21_X1 u1_u9_u1_U45 (.B2( u1_u9_u1_n123 ) , .ZN( u1_u9_u1_n145 ) , .B1( u1_u9_u1_n160 ) , .A( u1_u9_u1_n185 ) );
  INV_X1 u1_u9_u1_U46 (.A( u1_u9_u1_n122 ) , .ZN( u1_u9_u1_n185 ) );
  AOI21_X1 u1_u9_u1_U47 (.B2( u1_u9_u1_n120 ) , .B1( u1_u9_u1_n121 ) , .ZN( u1_u9_u1_n122 ) , .A( u1_u9_u1_n128 ) );
  AOI21_X1 u1_u9_u1_U48 (.A( u1_u9_u1_n128 ) , .B2( u1_u9_u1_n129 ) , .ZN( u1_u9_u1_n130 ) , .B1( u1_u9_u1_n150 ) );
  NAND2_X1 u1_u9_u1_U49 (.ZN( u1_u9_u1_n112 ) , .A1( u1_u9_u1_n169 ) , .A2( u1_u9_u1_n170 ) );
  AOI211_X1 u1_u9_u1_U5 (.ZN( u1_u9_u1_n124 ) , .A( u1_u9_u1_n138 ) , .C2( u1_u9_u1_n139 ) , .B( u1_u9_u1_n145 ) , .C1( u1_u9_u1_n147 ) );
  NAND2_X1 u1_u9_u1_U50 (.ZN( u1_u9_u1_n129 ) , .A2( u1_u9_u1_n95 ) , .A1( u1_u9_u1_n98 ) );
  NAND2_X1 u1_u9_u1_U51 (.A1( u1_u9_u1_n102 ) , .ZN( u1_u9_u1_n154 ) , .A2( u1_u9_u1_n99 ) );
  NAND2_X1 u1_u9_u1_U52 (.A2( u1_u9_u1_n100 ) , .ZN( u1_u9_u1_n135 ) , .A1( u1_u9_u1_n99 ) );
  AOI21_X1 u1_u9_u1_U53 (.A( u1_u9_u1_n152 ) , .B2( u1_u9_u1_n153 ) , .B1( u1_u9_u1_n154 ) , .ZN( u1_u9_u1_n158 ) );
  INV_X1 u1_u9_u1_U54 (.A( u1_u9_u1_n160 ) , .ZN( u1_u9_u1_n175 ) );
  NAND2_X1 u1_u9_u1_U55 (.A1( u1_u9_u1_n100 ) , .ZN( u1_u9_u1_n116 ) , .A2( u1_u9_u1_n95 ) );
  NAND2_X1 u1_u9_u1_U56 (.A1( u1_u9_u1_n102 ) , .ZN( u1_u9_u1_n131 ) , .A2( u1_u9_u1_n95 ) );
  NAND2_X1 u1_u9_u1_U57 (.A2( u1_u9_u1_n104 ) , .ZN( u1_u9_u1_n121 ) , .A1( u1_u9_u1_n98 ) );
  NAND2_X1 u1_u9_u1_U58 (.A1( u1_u9_u1_n103 ) , .ZN( u1_u9_u1_n153 ) , .A2( u1_u9_u1_n98 ) );
  NAND2_X1 u1_u9_u1_U59 (.A2( u1_u9_u1_n104 ) , .A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n133 ) );
  AOI22_X1 u1_u9_u1_U6 (.B2( u1_u9_u1_n136 ) , .A2( u1_u9_u1_n137 ) , .ZN( u1_u9_u1_n143 ) , .A1( u1_u9_u1_n171 ) , .B1( u1_u9_u1_n173 ) );
  NAND2_X1 u1_u9_u1_U60 (.ZN( u1_u9_u1_n150 ) , .A2( u1_u9_u1_n98 ) , .A1( u1_u9_u1_n99 ) );
  NAND2_X1 u1_u9_u1_U61 (.A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n155 ) , .A2( u1_u9_u1_n95 ) );
  OAI21_X1 u1_u9_u1_U62 (.ZN( u1_u9_u1_n109 ) , .B1( u1_u9_u1_n129 ) , .B2( u1_u9_u1_n160 ) , .A( u1_u9_u1_n167 ) );
  NAND2_X1 u1_u9_u1_U63 (.A2( u1_u9_u1_n100 ) , .A1( u1_u9_u1_n103 ) , .ZN( u1_u9_u1_n120 ) );
  NAND2_X1 u1_u9_u1_U64 (.A1( u1_u9_u1_n102 ) , .A2( u1_u9_u1_n104 ) , .ZN( u1_u9_u1_n115 ) );
  NAND2_X1 u1_u9_u1_U65 (.A2( u1_u9_u1_n100 ) , .A1( u1_u9_u1_n104 ) , .ZN( u1_u9_u1_n151 ) );
  NAND2_X1 u1_u9_u1_U66 (.A2( u1_u9_u1_n103 ) , .A1( u1_u9_u1_n105 ) , .ZN( u1_u9_u1_n161 ) );
  INV_X1 u1_u9_u1_U67 (.A( u1_u9_u1_n152 ) , .ZN( u1_u9_u1_n173 ) );
  INV_X1 u1_u9_u1_U68 (.A( u1_u9_u1_n128 ) , .ZN( u1_u9_u1_n172 ) );
  NAND2_X1 u1_u9_u1_U69 (.A2( u1_u9_u1_n102 ) , .A1( u1_u9_u1_n103 ) , .ZN( u1_u9_u1_n123 ) );
  INV_X1 u1_u9_u1_U7 (.A( u1_u9_u1_n147 ) , .ZN( u1_u9_u1_n181 ) );
  NOR2_X1 u1_u9_u1_U70 (.A2( u1_u9_X_7 ) , .A1( u1_u9_X_8 ) , .ZN( u1_u9_u1_n95 ) );
  NOR2_X1 u1_u9_u1_U71 (.A1( u1_u9_X_12 ) , .A2( u1_u9_X_9 ) , .ZN( u1_u9_u1_n100 ) );
  NOR2_X1 u1_u9_u1_U72 (.A2( u1_u9_X_8 ) , .A1( u1_u9_u1_n177 ) , .ZN( u1_u9_u1_n99 ) );
  NOR2_X1 u1_u9_u1_U73 (.A2( u1_u9_X_12 ) , .ZN( u1_u9_u1_n102 ) , .A1( u1_u9_u1_n176 ) );
  NOR2_X1 u1_u9_u1_U74 (.A2( u1_u9_X_9 ) , .ZN( u1_u9_u1_n105 ) , .A1( u1_u9_u1_n168 ) );
  NAND2_X1 u1_u9_u1_U75 (.A1( u1_u9_X_10 ) , .ZN( u1_u9_u1_n160 ) , .A2( u1_u9_u1_n169 ) );
  NAND2_X1 u1_u9_u1_U76 (.A2( u1_u9_X_10 ) , .A1( u1_u9_X_11 ) , .ZN( u1_u9_u1_n152 ) );
  NAND2_X1 u1_u9_u1_U77 (.A1( u1_u9_X_11 ) , .ZN( u1_u9_u1_n128 ) , .A2( u1_u9_u1_n170 ) );
  AND2_X1 u1_u9_u1_U78 (.A2( u1_u9_X_7 ) , .A1( u1_u9_X_8 ) , .ZN( u1_u9_u1_n104 ) );
  AND2_X1 u1_u9_u1_U79 (.A1( u1_u9_X_8 ) , .ZN( u1_u9_u1_n103 ) , .A2( u1_u9_u1_n177 ) );
  AOI22_X1 u1_u9_u1_U8 (.B2( u1_u9_u1_n113 ) , .A2( u1_u9_u1_n114 ) , .ZN( u1_u9_u1_n125 ) , .A1( u1_u9_u1_n171 ) , .B1( u1_u9_u1_n173 ) );
  INV_X1 u1_u9_u1_U80 (.A( u1_u9_X_10 ) , .ZN( u1_u9_u1_n170 ) );
  INV_X1 u1_u9_u1_U81 (.A( u1_u9_X_9 ) , .ZN( u1_u9_u1_n176 ) );
  INV_X1 u1_u9_u1_U82 (.A( u1_u9_X_11 ) , .ZN( u1_u9_u1_n169 ) );
  INV_X1 u1_u9_u1_U83 (.A( u1_u9_X_12 ) , .ZN( u1_u9_u1_n168 ) );
  INV_X1 u1_u9_u1_U84 (.A( u1_u9_X_7 ) , .ZN( u1_u9_u1_n177 ) );
  NAND4_X1 u1_u9_u1_U85 (.ZN( u1_out9_18 ) , .A4( u1_u9_u1_n165 ) , .A3( u1_u9_u1_n166 ) , .A1( u1_u9_u1_n167 ) , .A2( u1_u9_u1_n186 ) );
  AOI22_X1 u1_u9_u1_U86 (.B2( u1_u9_u1_n146 ) , .B1( u1_u9_u1_n147 ) , .A2( u1_u9_u1_n148 ) , .ZN( u1_u9_u1_n166 ) , .A1( u1_u9_u1_n172 ) );
  INV_X1 u1_u9_u1_U87 (.A( u1_u9_u1_n145 ) , .ZN( u1_u9_u1_n186 ) );
  NAND4_X1 u1_u9_u1_U88 (.ZN( u1_out9_2 ) , .A4( u1_u9_u1_n142 ) , .A3( u1_u9_u1_n143 ) , .A2( u1_u9_u1_n144 ) , .A1( u1_u9_u1_n179 ) );
  OAI21_X1 u1_u9_u1_U89 (.B2( u1_u9_u1_n132 ) , .ZN( u1_u9_u1_n144 ) , .A( u1_u9_u1_n146 ) , .B1( u1_u9_u1_n180 ) );
  NAND2_X1 u1_u9_u1_U9 (.ZN( u1_u9_u1_n114 ) , .A1( u1_u9_u1_n134 ) , .A2( u1_u9_u1_n156 ) );
  INV_X1 u1_u9_u1_U90 (.A( u1_u9_u1_n130 ) , .ZN( u1_u9_u1_n179 ) );
  NAND4_X1 u1_u9_u1_U91 (.ZN( u1_out9_28 ) , .A4( u1_u9_u1_n124 ) , .A3( u1_u9_u1_n125 ) , .A2( u1_u9_u1_n126 ) , .A1( u1_u9_u1_n127 ) );
  OAI21_X1 u1_u9_u1_U92 (.ZN( u1_u9_u1_n127 ) , .B2( u1_u9_u1_n139 ) , .B1( u1_u9_u1_n175 ) , .A( u1_u9_u1_n183 ) );
  OAI21_X1 u1_u9_u1_U93 (.ZN( u1_u9_u1_n126 ) , .B2( u1_u9_u1_n140 ) , .A( u1_u9_u1_n146 ) , .B1( u1_u9_u1_n178 ) );
  OR4_X1 u1_u9_u1_U94 (.ZN( u1_out9_13 ) , .A4( u1_u9_u1_n108 ) , .A3( u1_u9_u1_n109 ) , .A2( u1_u9_u1_n110 ) , .A1( u1_u9_u1_n111 ) );
  AOI21_X1 u1_u9_u1_U95 (.ZN( u1_u9_u1_n110 ) , .A( u1_u9_u1_n116 ) , .B1( u1_u9_u1_n152 ) , .B2( u1_u9_u1_n160 ) );
  AOI21_X1 u1_u9_u1_U96 (.ZN( u1_u9_u1_n111 ) , .A( u1_u9_u1_n128 ) , .B2( u1_u9_u1_n131 ) , .B1( u1_u9_u1_n135 ) );
  NAND3_X1 u1_u9_u1_U97 (.A3( u1_u9_u1_n149 ) , .A2( u1_u9_u1_n150 ) , .A1( u1_u9_u1_n151 ) , .ZN( u1_u9_u1_n164 ) );
  NAND3_X1 u1_u9_u1_U98 (.A3( u1_u9_u1_n134 ) , .A2( u1_u9_u1_n135 ) , .ZN( u1_u9_u1_n136 ) , .A1( u1_u9_u1_n151 ) );
  NAND3_X1 u1_u9_u1_U99 (.A1( u1_u9_u1_n133 ) , .ZN( u1_u9_u1_n137 ) , .A2( u1_u9_u1_n154 ) , .A3( u1_u9_u1_n181 ) );
  OAI22_X1 u1_u9_u2_U10 (.B1( u1_u9_u2_n151 ) , .A2( u1_u9_u2_n152 ) , .A1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n160 ) , .B2( u1_u9_u2_n168 ) );
  NAND3_X1 u1_u9_u2_U100 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n98 ) );
  NOR3_X1 u1_u9_u2_U11 (.A1( u1_u9_u2_n150 ) , .ZN( u1_u9_u2_n151 ) , .A3( u1_u9_u2_n175 ) , .A2( u1_u9_u2_n188 ) );
  AOI21_X1 u1_u9_u2_U12 (.B2( u1_u9_u2_n123 ) , .ZN( u1_u9_u2_n125 ) , .A( u1_u9_u2_n171 ) , .B1( u1_u9_u2_n184 ) );
  INV_X1 u1_u9_u2_U13 (.A( u1_u9_u2_n150 ) , .ZN( u1_u9_u2_n184 ) );
  AOI21_X1 u1_u9_u2_U14 (.ZN( u1_u9_u2_n144 ) , .B2( u1_u9_u2_n155 ) , .A( u1_u9_u2_n172 ) , .B1( u1_u9_u2_n185 ) );
  AOI21_X1 u1_u9_u2_U15 (.B2( u1_u9_u2_n143 ) , .ZN( u1_u9_u2_n145 ) , .B1( u1_u9_u2_n152 ) , .A( u1_u9_u2_n171 ) );
  INV_X1 u1_u9_u2_U16 (.A( u1_u9_u2_n156 ) , .ZN( u1_u9_u2_n171 ) );
  INV_X1 u1_u9_u2_U17 (.A( u1_u9_u2_n120 ) , .ZN( u1_u9_u2_n188 ) );
  NAND2_X1 u1_u9_u2_U18 (.A2( u1_u9_u2_n122 ) , .ZN( u1_u9_u2_n150 ) , .A1( u1_u9_u2_n152 ) );
  INV_X1 u1_u9_u2_U19 (.A( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n170 ) );
  INV_X1 u1_u9_u2_U20 (.A( u1_u9_u2_n137 ) , .ZN( u1_u9_u2_n173 ) );
  NAND2_X1 u1_u9_u2_U21 (.A1( u1_u9_u2_n132 ) , .A2( u1_u9_u2_n139 ) , .ZN( u1_u9_u2_n157 ) );
  INV_X1 u1_u9_u2_U22 (.A( u1_u9_u2_n113 ) , .ZN( u1_u9_u2_n178 ) );
  INV_X1 u1_u9_u2_U23 (.A( u1_u9_u2_n139 ) , .ZN( u1_u9_u2_n175 ) );
  INV_X1 u1_u9_u2_U24 (.A( u1_u9_u2_n155 ) , .ZN( u1_u9_u2_n181 ) );
  INV_X1 u1_u9_u2_U25 (.A( u1_u9_u2_n119 ) , .ZN( u1_u9_u2_n177 ) );
  INV_X1 u1_u9_u2_U26 (.A( u1_u9_u2_n116 ) , .ZN( u1_u9_u2_n180 ) );
  INV_X1 u1_u9_u2_U27 (.A( u1_u9_u2_n131 ) , .ZN( u1_u9_u2_n179 ) );
  INV_X1 u1_u9_u2_U28 (.A( u1_u9_u2_n154 ) , .ZN( u1_u9_u2_n176 ) );
  NAND2_X1 u1_u9_u2_U29 (.A2( u1_u9_u2_n116 ) , .A1( u1_u9_u2_n117 ) , .ZN( u1_u9_u2_n118 ) );
  NOR2_X1 u1_u9_u2_U3 (.ZN( u1_u9_u2_n121 ) , .A2( u1_u9_u2_n177 ) , .A1( u1_u9_u2_n180 ) );
  INV_X1 u1_u9_u2_U30 (.A( u1_u9_u2_n132 ) , .ZN( u1_u9_u2_n182 ) );
  INV_X1 u1_u9_u2_U31 (.A( u1_u9_u2_n158 ) , .ZN( u1_u9_u2_n183 ) );
  OAI21_X1 u1_u9_u2_U32 (.A( u1_u9_u2_n156 ) , .B1( u1_u9_u2_n157 ) , .ZN( u1_u9_u2_n158 ) , .B2( u1_u9_u2_n179 ) );
  NOR2_X1 u1_u9_u2_U33 (.ZN( u1_u9_u2_n156 ) , .A1( u1_u9_u2_n166 ) , .A2( u1_u9_u2_n169 ) );
  NOR2_X1 u1_u9_u2_U34 (.A2( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n137 ) , .A1( u1_u9_u2_n140 ) );
  NOR2_X1 u1_u9_u2_U35 (.A2( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n153 ) , .A1( u1_u9_u2_n156 ) );
  AOI211_X1 u1_u9_u2_U36 (.ZN( u1_u9_u2_n130 ) , .C1( u1_u9_u2_n138 ) , .C2( u1_u9_u2_n179 ) , .B( u1_u9_u2_n96 ) , .A( u1_u9_u2_n97 ) );
  OAI22_X1 u1_u9_u2_U37 (.B1( u1_u9_u2_n133 ) , .A2( u1_u9_u2_n137 ) , .A1( u1_u9_u2_n152 ) , .B2( u1_u9_u2_n168 ) , .ZN( u1_u9_u2_n97 ) );
  OAI221_X1 u1_u9_u2_U38 (.B1( u1_u9_u2_n113 ) , .C1( u1_u9_u2_n132 ) , .A( u1_u9_u2_n149 ) , .B2( u1_u9_u2_n171 ) , .C2( u1_u9_u2_n172 ) , .ZN( u1_u9_u2_n96 ) );
  OAI221_X1 u1_u9_u2_U39 (.A( u1_u9_u2_n115 ) , .C2( u1_u9_u2_n123 ) , .B2( u1_u9_u2_n143 ) , .B1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n163 ) , .C1( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U4 (.A( u1_u9_u2_n134 ) , .ZN( u1_u9_u2_n185 ) );
  OAI21_X1 u1_u9_u2_U40 (.A( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n115 ) , .B1( u1_u9_u2_n176 ) , .B2( u1_u9_u2_n178 ) );
  OAI221_X1 u1_u9_u2_U41 (.A( u1_u9_u2_n135 ) , .B2( u1_u9_u2_n136 ) , .B1( u1_u9_u2_n137 ) , .ZN( u1_u9_u2_n162 ) , .C2( u1_u9_u2_n167 ) , .C1( u1_u9_u2_n185 ) );
  AND3_X1 u1_u9_u2_U42 (.A3( u1_u9_u2_n131 ) , .A2( u1_u9_u2_n132 ) , .A1( u1_u9_u2_n133 ) , .ZN( u1_u9_u2_n136 ) );
  AOI22_X1 u1_u9_u2_U43 (.ZN( u1_u9_u2_n135 ) , .B1( u1_u9_u2_n140 ) , .A1( u1_u9_u2_n156 ) , .B2( u1_u9_u2_n180 ) , .A2( u1_u9_u2_n188 ) );
  AOI21_X1 u1_u9_u2_U44 (.ZN( u1_u9_u2_n149 ) , .B1( u1_u9_u2_n173 ) , .B2( u1_u9_u2_n188 ) , .A( u1_u9_u2_n95 ) );
  AND3_X1 u1_u9_u2_U45 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n156 ) , .ZN( u1_u9_u2_n95 ) );
  OAI21_X1 u1_u9_u2_U46 (.A( u1_u9_u2_n101 ) , .B2( u1_u9_u2_n121 ) , .B1( u1_u9_u2_n153 ) , .ZN( u1_u9_u2_n164 ) );
  NAND2_X1 u1_u9_u2_U47 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n155 ) );
  NAND2_X1 u1_u9_u2_U48 (.A2( u1_u9_u2_n105 ) , .A1( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n143 ) );
  NAND2_X1 u1_u9_u2_U49 (.A1( u1_u9_u2_n104 ) , .A2( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n152 ) );
  NOR4_X1 u1_u9_u2_U5 (.A4( u1_u9_u2_n124 ) , .A3( u1_u9_u2_n125 ) , .A2( u1_u9_u2_n126 ) , .A1( u1_u9_u2_n127 ) , .ZN( u1_u9_u2_n128 ) );
  NAND2_X1 u1_u9_u2_U50 (.A1( u1_u9_u2_n100 ) , .A2( u1_u9_u2_n105 ) , .ZN( u1_u9_u2_n132 ) );
  INV_X1 u1_u9_u2_U51 (.A( u1_u9_u2_n140 ) , .ZN( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U52 (.A( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n167 ) );
  OAI21_X1 u1_u9_u2_U53 (.A( u1_u9_u2_n141 ) , .B2( u1_u9_u2_n142 ) , .ZN( u1_u9_u2_n146 ) , .B1( u1_u9_u2_n153 ) );
  OAI21_X1 u1_u9_u2_U54 (.A( u1_u9_u2_n140 ) , .ZN( u1_u9_u2_n141 ) , .B1( u1_u9_u2_n176 ) , .B2( u1_u9_u2_n177 ) );
  NOR3_X1 u1_u9_u2_U55 (.ZN( u1_u9_u2_n142 ) , .A3( u1_u9_u2_n175 ) , .A2( u1_u9_u2_n178 ) , .A1( u1_u9_u2_n181 ) );
  NAND2_X1 u1_u9_u2_U56 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n113 ) );
  NAND2_X1 u1_u9_u2_U57 (.A1( u1_u9_u2_n106 ) , .A2( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n131 ) );
  NAND2_X1 u1_u9_u2_U58 (.A1( u1_u9_u2_n103 ) , .A2( u1_u9_u2_n107 ) , .ZN( u1_u9_u2_n139 ) );
  NAND2_X1 u1_u9_u2_U59 (.A1( u1_u9_u2_n103 ) , .A2( u1_u9_u2_n105 ) , .ZN( u1_u9_u2_n133 ) );
  AOI21_X1 u1_u9_u2_U6 (.B2( u1_u9_u2_n119 ) , .ZN( u1_u9_u2_n127 ) , .A( u1_u9_u2_n137 ) , .B1( u1_u9_u2_n155 ) );
  NAND2_X1 u1_u9_u2_U60 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n103 ) , .ZN( u1_u9_u2_n154 ) );
  NAND2_X1 u1_u9_u2_U61 (.A2( u1_u9_u2_n103 ) , .A1( u1_u9_u2_n104 ) , .ZN( u1_u9_u2_n119 ) );
  NAND2_X1 u1_u9_u2_U62 (.A2( u1_u9_u2_n107 ) , .A1( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n123 ) );
  NAND2_X1 u1_u9_u2_U63 (.A1( u1_u9_u2_n104 ) , .A2( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n122 ) );
  INV_X1 u1_u9_u2_U64 (.A( u1_u9_u2_n114 ) , .ZN( u1_u9_u2_n172 ) );
  NAND2_X1 u1_u9_u2_U65 (.A2( u1_u9_u2_n100 ) , .A1( u1_u9_u2_n102 ) , .ZN( u1_u9_u2_n116 ) );
  NAND2_X1 u1_u9_u2_U66 (.A1( u1_u9_u2_n102 ) , .A2( u1_u9_u2_n108 ) , .ZN( u1_u9_u2_n120 ) );
  NAND2_X1 u1_u9_u2_U67 (.A2( u1_u9_u2_n105 ) , .A1( u1_u9_u2_n106 ) , .ZN( u1_u9_u2_n117 ) );
  INV_X1 u1_u9_u2_U68 (.ZN( u1_u9_u2_n187 ) , .A( u1_u9_u2_n99 ) );
  OAI21_X1 u1_u9_u2_U69 (.B1( u1_u9_u2_n137 ) , .B2( u1_u9_u2_n143 ) , .A( u1_u9_u2_n98 ) , .ZN( u1_u9_u2_n99 ) );
  AOI21_X1 u1_u9_u2_U7 (.ZN( u1_u9_u2_n124 ) , .B1( u1_u9_u2_n131 ) , .B2( u1_u9_u2_n143 ) , .A( u1_u9_u2_n172 ) );
  NOR2_X1 u1_u9_u2_U70 (.A2( u1_u9_X_16 ) , .ZN( u1_u9_u2_n140 ) , .A1( u1_u9_u2_n166 ) );
  NOR2_X1 u1_u9_u2_U71 (.A2( u1_u9_X_13 ) , .A1( u1_u9_X_14 ) , .ZN( u1_u9_u2_n100 ) );
  NOR2_X1 u1_u9_u2_U72 (.A2( u1_u9_X_16 ) , .A1( u1_u9_X_17 ) , .ZN( u1_u9_u2_n138 ) );
  NOR2_X1 u1_u9_u2_U73 (.A2( u1_u9_X_15 ) , .A1( u1_u9_X_18 ) , .ZN( u1_u9_u2_n104 ) );
  NOR2_X1 u1_u9_u2_U74 (.A2( u1_u9_X_14 ) , .ZN( u1_u9_u2_n103 ) , .A1( u1_u9_u2_n174 ) );
  NOR2_X1 u1_u9_u2_U75 (.A2( u1_u9_X_15 ) , .ZN( u1_u9_u2_n102 ) , .A1( u1_u9_u2_n165 ) );
  NOR2_X1 u1_u9_u2_U76 (.A2( u1_u9_X_17 ) , .ZN( u1_u9_u2_n114 ) , .A1( u1_u9_u2_n169 ) );
  AND2_X1 u1_u9_u2_U77 (.A1( u1_u9_X_15 ) , .ZN( u1_u9_u2_n105 ) , .A2( u1_u9_u2_n165 ) );
  AND2_X1 u1_u9_u2_U78 (.A2( u1_u9_X_15 ) , .A1( u1_u9_X_18 ) , .ZN( u1_u9_u2_n107 ) );
  AND2_X1 u1_u9_u2_U79 (.A1( u1_u9_X_14 ) , .ZN( u1_u9_u2_n106 ) , .A2( u1_u9_u2_n174 ) );
  AOI21_X1 u1_u9_u2_U8 (.B2( u1_u9_u2_n120 ) , .B1( u1_u9_u2_n121 ) , .ZN( u1_u9_u2_n126 ) , .A( u1_u9_u2_n167 ) );
  AND2_X1 u1_u9_u2_U80 (.A1( u1_u9_X_13 ) , .A2( u1_u9_X_14 ) , .ZN( u1_u9_u2_n108 ) );
  INV_X1 u1_u9_u2_U81 (.A( u1_u9_X_16 ) , .ZN( u1_u9_u2_n169 ) );
  INV_X1 u1_u9_u2_U82 (.A( u1_u9_X_17 ) , .ZN( u1_u9_u2_n166 ) );
  INV_X1 u1_u9_u2_U83 (.A( u1_u9_X_13 ) , .ZN( u1_u9_u2_n174 ) );
  INV_X1 u1_u9_u2_U84 (.A( u1_u9_X_18 ) , .ZN( u1_u9_u2_n165 ) );
  NAND4_X1 u1_u9_u2_U85 (.ZN( u1_out9_24 ) , .A4( u1_u9_u2_n111 ) , .A3( u1_u9_u2_n112 ) , .A1( u1_u9_u2_n130 ) , .A2( u1_u9_u2_n187 ) );
  AOI221_X1 u1_u9_u2_U86 (.A( u1_u9_u2_n109 ) , .B1( u1_u9_u2_n110 ) , .ZN( u1_u9_u2_n111 ) , .C1( u1_u9_u2_n134 ) , .C2( u1_u9_u2_n170 ) , .B2( u1_u9_u2_n173 ) );
  AOI21_X1 u1_u9_u2_U87 (.ZN( u1_u9_u2_n112 ) , .B2( u1_u9_u2_n156 ) , .A( u1_u9_u2_n164 ) , .B1( u1_u9_u2_n181 ) );
  NAND4_X1 u1_u9_u2_U88 (.ZN( u1_out9_16 ) , .A4( u1_u9_u2_n128 ) , .A3( u1_u9_u2_n129 ) , .A1( u1_u9_u2_n130 ) , .A2( u1_u9_u2_n186 ) );
  AOI22_X1 u1_u9_u2_U89 (.A2( u1_u9_u2_n118 ) , .ZN( u1_u9_u2_n129 ) , .A1( u1_u9_u2_n140 ) , .B1( u1_u9_u2_n157 ) , .B2( u1_u9_u2_n170 ) );
  OAI22_X1 u1_u9_u2_U9 (.ZN( u1_u9_u2_n109 ) , .A2( u1_u9_u2_n113 ) , .B2( u1_u9_u2_n133 ) , .B1( u1_u9_u2_n167 ) , .A1( u1_u9_u2_n168 ) );
  INV_X1 u1_u9_u2_U90 (.A( u1_u9_u2_n163 ) , .ZN( u1_u9_u2_n186 ) );
  NAND4_X1 u1_u9_u2_U91 (.ZN( u1_out9_30 ) , .A4( u1_u9_u2_n147 ) , .A3( u1_u9_u2_n148 ) , .A2( u1_u9_u2_n149 ) , .A1( u1_u9_u2_n187 ) );
  AOI21_X1 u1_u9_u2_U92 (.B2( u1_u9_u2_n138 ) , .ZN( u1_u9_u2_n148 ) , .A( u1_u9_u2_n162 ) , .B1( u1_u9_u2_n182 ) );
  NOR3_X1 u1_u9_u2_U93 (.A3( u1_u9_u2_n144 ) , .A2( u1_u9_u2_n145 ) , .A1( u1_u9_u2_n146 ) , .ZN( u1_u9_u2_n147 ) );
  OR4_X1 u1_u9_u2_U94 (.ZN( u1_out9_6 ) , .A4( u1_u9_u2_n161 ) , .A3( u1_u9_u2_n162 ) , .A2( u1_u9_u2_n163 ) , .A1( u1_u9_u2_n164 ) );
  OR3_X1 u1_u9_u2_U95 (.A2( u1_u9_u2_n159 ) , .A1( u1_u9_u2_n160 ) , .ZN( u1_u9_u2_n161 ) , .A3( u1_u9_u2_n183 ) );
  AOI21_X1 u1_u9_u2_U96 (.B2( u1_u9_u2_n154 ) , .B1( u1_u9_u2_n155 ) , .ZN( u1_u9_u2_n159 ) , .A( u1_u9_u2_n167 ) );
  NAND3_X1 u1_u9_u2_U97 (.A2( u1_u9_u2_n117 ) , .A1( u1_u9_u2_n122 ) , .A3( u1_u9_u2_n123 ) , .ZN( u1_u9_u2_n134 ) );
  NAND3_X1 u1_u9_u2_U98 (.ZN( u1_u9_u2_n110 ) , .A2( u1_u9_u2_n131 ) , .A3( u1_u9_u2_n139 ) , .A1( u1_u9_u2_n154 ) );
  NAND3_X1 u1_u9_u2_U99 (.A2( u1_u9_u2_n100 ) , .ZN( u1_u9_u2_n101 ) , .A1( u1_u9_u2_n104 ) , .A3( u1_u9_u2_n114 ) );
  OAI21_X1 u1_uk_U1020 (.ZN( u1_K1_13 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1214 ) , .A( u1_uk_n999 ) );
  NAND2_X1 u1_uk_U1021 (.A1( u1_key_r_46 ) , .A2( u1_uk_n146 ) , .ZN( u1_uk_n999 ) );
  OAI21_X1 u1_uk_U1022 (.ZN( u1_K1_17 ) , .A( u1_uk_n1001 ) , .B2( u1_uk_n1183 ) , .B1( u1_uk_n129 ) );
  NAND2_X1 u1_uk_U1023 (.A1( u1_key_r_10 ) , .ZN( u1_uk_n1001 ) , .A2( u1_uk_n187 ) );
  OAI21_X1 u1_uk_U1038 (.ZN( u1_K10_13 ) , .B2( u1_uk_n1635 ) , .A( u1_uk_n301 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1039 (.A1( u1_uk_K_r8_48 ) , .ZN( u1_uk_n301 ) , .A2( u1_uk_n31 ) );
  INV_X1 u1_uk_U105 (.ZN( u1_K11_5 ) , .A( u1_uk_n496 ) );
  AOI22_X1 u1_uk_U106 (.B2( u1_uk_K_r9_19 ) , .A2( u1_uk_K_r9_25 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n250 ) , .ZN( u1_uk_n496 ) );
  OAI22_X1 u1_uk_U107 (.ZN( u1_K1_5 ) , .A2( u1_uk_n1176 ) , .B2( u1_uk_n1180 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U1080 (.A( u1_key_r_6 ) , .ZN( u1_uk_n1176 ) );
  INV_X1 u1_uk_U1081 (.A( u1_key_r_54 ) , .ZN( u1_uk_n1215 ) );
  INV_X1 u1_uk_U1082 (.A( u1_key_r_33 ) , .ZN( u1_uk_n1197 ) );
  INV_X1 u1_uk_U1084 (.A( u1_key_r_26 ) , .ZN( u1_uk_n1191 ) );
  INV_X1 u1_uk_U1085 (.A( u1_key_r_40 ) , .ZN( u1_uk_n1204 ) );
  INV_X1 u1_uk_U1087 (.A( u1_key_r_47 ) , .ZN( u1_uk_n1209 ) );
  INV_X1 u1_uk_U1088 (.A( u1_key_r_34 ) , .ZN( u1_uk_n1198 ) );
  INV_X1 u1_uk_U1089 (.A( u1_key_r_27 ) , .ZN( u1_uk_n1192 ) );
  INV_X1 u1_uk_U1090 (.A( u1_key_r_24 ) , .ZN( u1_uk_n1189 ) );
  INV_X1 u1_uk_U1091 (.A( u1_key_r_20 ) , .ZN( u1_uk_n1185 ) );
  INV_X1 u1_uk_U1096 (.A( u1_key_r_13 ) , .ZN( u1_uk_n1180 ) );
  INV_X1 u1_uk_U1099 (.A( u1_key_r_19 ) , .ZN( u1_uk_n1184 ) );
  INV_X1 u1_uk_U1100 (.A( u1_key_r_4 ) , .ZN( u1_uk_n1175 ) );
  INV_X1 u1_uk_U1101 (.A( u1_key_r_17 ) , .ZN( u1_uk_n1183 ) );
  INV_X1 u1_uk_U1102 (.A( u1_key_r_53 ) , .ZN( u1_uk_n1214 ) );
  OAI21_X1 u1_uk_U1107 (.ZN( u1_K16_14 ) , .B2( u1_uk_n1235 ) , .B1( u1_uk_n252 ) , .A( u1_uk_n981 ) );
  NAND2_X1 u1_uk_U1108 (.A1( u1_uk_K_r14_18 ) , .A2( u1_uk_n291 ) , .ZN( u1_uk_n981 ) );
  INV_X1 u1_uk_U1117 (.ZN( u1_K13_10 ) , .A( u1_uk_n671 ) );
  AOI22_X1 u1_uk_U1118 (.B2( u1_uk_K_r11_26 ) , .A2( u1_uk_K_r11_6 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n203 ) , .ZN( u1_uk_n671 ) );
  INV_X1 u1_uk_U112 (.ZN( u1_K13_5 ) , .A( u1_uk_n948 ) );
  INV_X1 u1_uk_U1121 (.ZN( u1_K2_10 ) , .A( u1_uk_n1021 ) );
  AOI22_X1 u1_uk_U1122 (.B2( u1_uk_K_r0_34 ) , .A2( u1_uk_K_r0_55 ) , .ZN( u1_uk_n1021 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) );
  INV_X1 u1_uk_U1123 (.ZN( u1_K1_11 ) , .A( u1_uk_n997 ) );
  AOI22_X1 u1_uk_U1124 (.B2( u1_key_r_32 ) , .A2( u1_key_r_39 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n277 ) , .ZN( u1_uk_n997 ) );
  INV_X1 u1_uk_U1125 (.ZN( u1_K1_18 ) , .A( u1_uk_n1002 ) );
  AOI22_X1 u1_uk_U1126 (.A2( u1_key_r_5 ) , .B2( u1_key_r_55 ) , .ZN( u1_uk_n1002 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n294 ) );
  INV_X1 u1_uk_U1129 (.ZN( u1_K11_8 ) , .A( u1_uk_n501 ) );
  AOI22_X1 u1_uk_U113 (.B2( u1_uk_K_r11_48 ) , .A2( u1_uk_K_r11_53 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n223 ) , .ZN( u1_uk_n948 ) );
  AOI22_X1 u1_uk_U1130 (.B2( u1_uk_K_r9_12 ) , .A2( u1_uk_K_r9_18 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n501 ) );
  INV_X1 u1_uk_U1131 (.ZN( u1_K11_12 ) , .A( u1_uk_n379 ) );
  AOI22_X1 u1_uk_U1132 (.B2( u1_uk_K_r9_25 ) , .A2( u1_uk_K_r9_6 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n291 ) , .ZN( u1_uk_n379 ) );
  INV_X1 u1_uk_U1135 (.ZN( u1_K2_7 ) , .A( u1_uk_n1034 ) );
  AOI22_X1 u1_uk_U1136 (.B2( u1_uk_K_r0_13 ) , .A2( u1_uk_K_r0_34 ) , .ZN( u1_uk_n1034 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n27 ) );
  INV_X1 u1_uk_U1137 (.ZN( u1_K1_20 ) , .A( u1_uk_n1003 ) );
  AOI22_X1 u1_uk_U1138 (.B2( u1_key_r_48 ) , .A2( u1_key_r_55 ) , .ZN( u1_uk_n1003 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n250 ) );
  INV_X1 u1_uk_U1157 (.ZN( u1_K10_12 ) , .A( u1_uk_n299 ) );
  AOI22_X1 u1_uk_U1158 (.B2( u1_uk_K_r8_17 ) , .A2( u1_uk_K_r8_39 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n297 ) , .ZN( u1_uk_n299 ) );
  INV_X1 u1_uk_U1163 (.ZN( u1_K13_12 ) , .A( u1_uk_n676 ) );
  AOI22_X1 u1_uk_U1164 (.B2( u1_uk_K_r11_34 ) , .A2( u1_uk_K_r11_54 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n252 ) , .ZN( u1_uk_n676 ) );
  AOI22_X1 u1_uk_U1167 (.B2( u1_uk_K_r11_26 ) , .A2( u1_uk_K_r11_46 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n27 ) , .ZN( u1_uk_n702 ) );
  INV_X1 u1_uk_U1168 (.ZN( u1_K13_2 ) , .A( u1_uk_n702 ) );
  INV_X1 u1_uk_U1172 (.ZN( u1_K13_6 ) , .A( u1_uk_n949 ) );
  OAI22_X1 u1_uk_U137 (.ZN( u1_K1_15 ) , .B2( u1_uk_n1191 ) , .A2( u1_uk_n1197 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U147 (.ZN( u1_K13_19 ) , .A( u1_uk_n685 ) );
  AOI22_X1 u1_uk_U148 (.B2( u1_uk_K_r11_19 ) , .A2( u1_uk_K_r11_39 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n252 ) , .ZN( u1_uk_n685 ) );
  OAI22_X1 u1_uk_U149 (.ZN( u1_K11_15 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1676 ) , .A2( u1_uk_n1691 ) , .A1( u1_uk_n297 ) );
  OAI21_X1 u1_uk_U152 (.ZN( u1_K2_15 ) , .A( u1_uk_n1024 ) , .B2( u1_uk_n1291 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U153 (.A1( u1_uk_K_r0_19 ) , .ZN( u1_uk_n1024 ) , .A2( u1_uk_n118 ) );
  OAI22_X1 u1_uk_U154 (.ZN( u1_K1_19 ) , .B2( u1_uk_n1175 ) , .A2( u1_uk_n1215 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U155 (.ZN( u1_K16_15 ) , .B2( u1_uk_n1236 ) , .A2( u1_uk_n1243 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U156 (.ZN( u1_K10_15 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1622 ) , .B2( u1_uk_n1659 ) , .B1( u1_uk_n286 ) );
  INV_X1 u1_uk_U18 (.ZN( u1_uk_n118 ) , .A( u1_uk_n220 ) );
  OAI21_X1 u1_uk_U181 (.ZN( u1_K1_14 ) , .A( u1_uk_n1000 ) , .B2( u1_uk_n1190 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U182 (.A1( u1_key_r_18 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1000 ) );
  INV_X1 u1_uk_U183 (.A( u1_key_r_25 ) , .ZN( u1_uk_n1190 ) );
  INV_X1 u1_uk_U190 (.ZN( u1_K11_14 ) , .A( u1_uk_n382 ) );
  AOI22_X1 u1_uk_U191 (.B2( u1_uk_K_r9_12 ) , .A2( u1_uk_K_r9_6 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n207 ) , .ZN( u1_uk_n382 ) );
  INV_X1 u1_uk_U195 (.ZN( u1_K2_14 ) , .A( u1_uk_n1023 ) );
  AOI22_X1 u1_uk_U196 (.B2( u1_uk_K_r0_11 ) , .A2( u1_uk_K_r0_32 ) , .ZN( u1_uk_n1023 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U197 (.ZN( u1_K1_24 ) , .B2( u1_uk_n1180 ) , .A2( u1_uk_n1185 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U198 (.ZN( u1_K10_14 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1630 ) , .A2( u1_uk_n1661 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U20 (.ZN( u1_uk_n142 ) , .A( u1_uk_n251 ) );
  INV_X1 u1_uk_U21 (.ZN( u1_uk_n128 ) , .A( u1_uk_n297 ) );
  INV_X1 u1_uk_U226 (.ZN( u1_K11_31 ) , .A( u1_uk_n437 ) );
  AOI22_X1 u1_uk_U227 (.B2( u1_uk_K_r9_22 ) , .A2( u1_uk_K_r9_30 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n251 ) , .ZN( u1_uk_n437 ) );
  OAI22_X1 u1_uk_U288 (.ZN( u1_K10_6 ) , .B1( u1_uk_n129 ) , .A2( u1_uk_n1621 ) , .B2( u1_uk_n1649 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U298 (.ZN( u1_K1_8 ) , .A1( u1_uk_n100 ) , .A2( u1_uk_n1176 ) , .B2( u1_uk_n1189 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U305 (.ZN( u1_K5_8 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1415 ) , .A2( u1_uk_n1437 ) , .B1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U309 (.ZN( u1_K2_8 ) , .A( u1_uk_n1035 ) , .B2( u1_uk_n1270 ) , .B1( u1_uk_n148 ) );
  NAND2_X1 u1_uk_U310 (.A1( u1_uk_K_r0_17 ) , .ZN( u1_uk_n1035 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U345 (.ZN( u1_K11_4 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1693 ) , .A2( u1_uk_n1699 ) , .B1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U349 (.ZN( u1_K1_4 ) , .A( u1_uk_n1020 ) , .B2( u1_uk_n1214 ) , .B1( u1_uk_n250 ) );
  NAND2_X1 u1_uk_U350 (.A1( u1_key_r_3 ) , .ZN( u1_uk_n1020 ) , .A2( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U361 (.ZN( u1_K10_4 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1642 ) , .A2( u1_uk_n1661 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U397 (.ZN( u1_K11_1 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1688 ) , .A2( u1_uk_n1705 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U403 (.ZN( u1_K1_9 ) , .B2( u1_uk_n1209 ) , .A2( u1_uk_n1215 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U405 (.ZN( u1_K10_16 ) , .B2( u1_uk_n1660 ) , .B1( u1_uk_n286 ) , .A( u1_uk_n305 ) );
  NAND2_X1 u1_uk_U406 (.A1( u1_uk_K_r8_32 ) , .A2( u1_uk_n203 ) , .ZN( u1_uk_n305 ) );
  OAI22_X1 u1_uk_U415 (.ZN( u1_K1_16 ) , .B2( u1_uk_n1192 ) , .A2( u1_uk_n1198 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U420 (.ZN( u1_K13_9 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1761 ) , .A2( u1_uk_n1773 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U422 (.ZN( u1_K11_9 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1663 ) , .A2( u1_uk_n1693 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U424 (.ZN( u1_K5_9 ) , .B2( u1_uk_n1427 ) , .A2( u1_uk_n1437 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U428 (.ZN( u1_K2_9 ) , .A2( u1_uk_n1262 ) , .B2( u1_uk_n1291 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U432 (.ZN( u1_K16_16 ) , .B2( u1_uk_n1237 ) , .A2( u1_uk_n1244 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U435 (.ZN( u1_K2_16 ) , .B2( u1_uk_n1274 ) , .A2( u1_uk_n1292 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U445 (.ZN( u1_K10_9 ) , .A( u1_uk_n376 ) );
  AOI22_X1 u1_uk_U446 (.B2( u1_uk_K_r8_17 ) , .A2( u1_uk_K_r8_27 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n297 ) , .ZN( u1_uk_n376 ) );
  OAI22_X1 u1_uk_U458 (.ZN( u1_K11_33 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1683 ) , .A2( u1_uk_n1689 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U506 (.ZN( u1_K11_2 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1673 ) , .A2( u1_uk_n1707 ) , .B1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U516 (.ZN( u1_K1_12 ) , .B2( u1_uk_n1184 ) , .B1( u1_uk_n148 ) , .A( u1_uk_n998 ) );
  NAND2_X1 u1_uk_U517 (.A1( u1_key_r_12 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n998 ) );
  OAI22_X1 u1_uk_U520 (.ZN( u1_K10_17 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1626 ) , .A2( u1_uk_n1654 ) , .B1( u1_uk_n251 ) );
  INV_X1 u1_uk_U536 (.ZN( u1_K11_17 ) , .A( u1_uk_n385 ) );
  AOI22_X1 u1_uk_U537 (.B2( u1_uk_K_r9_4 ) , .A2( u1_uk_K_r9_55 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n188 ) , .ZN( u1_uk_n385 ) );
  BUF_X1 u1_uk_U54 (.Z( u1_uk_n250 ) , .A( u1_uk_n257 ) );
  OAI21_X1 u1_uk_U540 (.ZN( u1_K5_12 ) , .A( u1_uk_n1071 ) , .B2( u1_uk_n1405 ) , .B1( u1_uk_n230 ) );
  NAND2_X1 u1_uk_U541 (.A1( u1_uk_K_r3_11 ) , .ZN( u1_uk_n1071 ) , .A2( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U544 (.ZN( u1_K2_12 ) , .A2( u1_uk_n1263 ) , .B2( u1_uk_n1278 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U548 (.ZN( u1_K16_17 ) , .B2( u1_uk_n1227 ) , .B1( u1_uk_n202 ) , .A( u1_uk_n982 ) );
  NAND2_X1 u1_uk_U549 (.A1( u1_uk_K_r14_10 ) , .A2( u1_uk_n257 ) , .ZN( u1_uk_n982 ) );
  INV_X1 u1_uk_U568 (.ZN( u1_K11_36 ) , .A( u1_uk_n454 ) );
  AOI22_X1 u1_uk_U569 (.B2( u1_uk_K_r9_15 ) , .A2( u1_uk_K_r9_7 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n202 ) , .ZN( u1_uk_n454 ) );
  OAI21_X1 u1_uk_U583 (.ZN( u1_K11_10 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1663 ) , .A( u1_uk_n377 ) );
  NAND2_X1 u1_uk_U584 (.A1( u1_uk_K_r9_54 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n377 ) );
  OAI22_X1 u1_uk_U585 (.ZN( u1_K10_10 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1625 ) , .A2( u1_uk_n1653 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U586 (.ZN( u1_K5_10 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1403 ) , .A2( u1_uk_n1423 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U594 (.ZN( u1_K1_10 ) , .A( u1_uk_n996 ) );
  AOI22_X1 u1_uk_U595 (.B2( u1_key_r_41 ) , .A2( u1_key_r_48 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n298 ) , .ZN( u1_uk_n996 ) );
  INV_X1 u1_uk_U599 (.ZN( u1_K13_22 ) , .A( u1_uk_n692 ) );
  AOI22_X1 u1_uk_U600 (.B2( u1_uk_K_r11_10 ) , .A2( u1_uk_K_r11_47 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n238 ) , .ZN( u1_uk_n692 ) );
  INV_X1 u1_uk_U610 (.ZN( u1_K1_22 ) , .A( u1_uk_n1004 ) );
  AOI22_X1 u1_uk_U611 (.B2( u1_key_r_25 ) , .A2( u1_key_r_32 ) , .ZN( u1_uk_n1004 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U613 (.ZN( u1_K11_35 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1695 ) , .A2( u1_uk_n1703 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U638 (.ZN( u1_K11_11 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1676 ) , .A2( u1_uk_n1682 ) , .B1( u1_uk_n251 ) );
  OAI21_X1 u1_uk_U640 (.ZN( u1_K2_11 ) , .A( u1_uk_n1022 ) , .B2( u1_uk_n1297 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U641 (.A1( u1_uk_K_r0_25 ) , .ZN( u1_uk_n1022 ) , .A2( u1_uk_n141 ) );
  INV_X1 u1_uk_U642 (.ZN( u1_K13_11 ) , .A( u1_uk_n672 ) );
  AOI22_X1 u1_uk_U643 (.B2( u1_uk_K_r11_17 ) , .A2( u1_uk_K_r11_54 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n191 ) , .ZN( u1_uk_n672 ) );
  OAI22_X1 u1_uk_U644 (.ZN( u1_K10_11 ) , .B2( u1_uk_n1626 ) , .A2( u1_uk_n1643 ) , .A1( u1_uk_n214 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U649 (.ZN( u1_K5_11 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1399 ) , .B2( u1_uk_n1423 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U661 (.ZN( u1_K11_3 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1669 ) , .A2( u1_uk_n1687 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U662 (.ZN( u1_K1_7 ) , .B2( u1_uk_n1185 ) , .A2( u1_uk_n1192 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U681 (.ZN( u1_K10_7 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1634 ) , .A2( u1_uk_n1654 ) , .A1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U686 (.ZN( u1_K11_7 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1691 ) , .A( u1_uk_n500 ) );
  NAND2_X1 u1_uk_U687 (.A1( u1_uk_K_r9_33 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n500 ) );
  INV_X1 u1_uk_U69 (.ZN( u1_K11_34 ) , .A( u1_uk_n443 ) );
  AOI22_X1 u1_uk_U70 (.B2( u1_uk_K_r9_45 ) , .A2( u1_uk_K_r9_49 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n443 ) );
  INV_X1 u1_uk_U709 (.ZN( u1_K13_7 ) , .A( u1_uk_n950 ) );
  AOI22_X1 u1_uk_U710 (.B2( u1_uk_K_r11_10 ) , .A2( u1_uk_K_r11_5 ) , .B1( u1_uk_n207 ) , .A1( u1_uk_n93 ) , .ZN( u1_uk_n950 ) );
  OAI21_X1 u1_uk_U711 (.ZN( u1_K5_7 ) , .A( u1_uk_n1087 ) , .B2( u1_uk_n1435 ) , .B1( u1_uk_n250 ) );
  NAND2_X1 u1_uk_U712 (.A1( u1_uk_K_r3_19 ) , .ZN( u1_uk_n1087 ) , .A2( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U718 (.ZN( u1_K10_2 ) , .B2( u1_uk_n1622 ) , .B1( u1_uk_n257 ) , .A( u1_uk_n338 ) );
  NAND2_X1 u1_uk_U719 (.A1( u1_uk_K_r8_41 ) , .A2( u1_uk_n188 ) , .ZN( u1_uk_n338 ) );
  OAI21_X1 u1_uk_U720 (.ZN( u1_K1_2 ) , .A( u1_uk_n1008 ) , .B2( u1_uk_n1175 ) , .B1( u1_uk_n242 ) );
  NAND2_X1 u1_uk_U721 (.A1( u1_key_r_11 ) , .ZN( u1_uk_n1008 ) , .A2( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U725 (.ZN( u1_K11_32 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1670 ) , .A2( u1_uk_n1690 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U756 (.ZN( u1_K11_13 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1688 ) , .A2( u1_uk_n1692 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U759 (.ZN( u1_K2_13 ) , .A2( u1_uk_n1261 ) , .B2( u1_uk_n1290 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U760 (.ZN( u1_K1_21 ) , .B2( u1_uk_n1183 ) , .A2( u1_uk_n1189 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n222 ) );
  INV_X1 u1_uk_U783 (.ZN( u1_K13_21 ) , .A( u1_uk_n689 ) );
  AOI22_X1 u1_uk_U784 (.B2( u1_uk_K_r11_34 ) , .A2( u1_uk_K_r11_39 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n230 ) , .ZN( u1_uk_n689 ) );
  OAI21_X1 u1_uk_U787 (.ZN( u1_K16_13 ) , .B2( u1_uk_n1257 ) , .B1( u1_uk_n297 ) , .A( u1_uk_n980 ) );
  NAND2_X1 u1_uk_U788 (.A1( u1_uk_K_r14_46 ) , .A2( u1_uk_n242 ) , .ZN( u1_uk_n980 ) );
  OAI21_X1 u1_uk_U803 (.ZN( u1_K13_1 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1757 ) , .A( u1_uk_n686 ) );
  NAND2_X1 u1_uk_U804 (.A1( u1_uk_K_r11_25 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n686 ) );
  OAI21_X1 u1_uk_U813 (.ZN( u1_K13_20 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1762 ) , .A( u1_uk_n688 ) );
  NAND2_X1 u1_uk_U814 (.A1( u1_uk_K_r11_33 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n688 ) );
  OAI22_X1 u1_uk_U820 (.ZN( u1_K2_18 ) , .B2( u1_uk_n1269 ) , .A2( u1_uk_n1300 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U821 (.ZN( u1_K16_18 ) , .B2( u1_uk_n1259 ) , .B1( u1_uk_n94 ) , .A( u1_uk_n983 ) );
  NAND2_X1 u1_uk_U822 (.A1( u1_uk_K_r14_5 ) , .A2( u1_uk_n118 ) , .ZN( u1_uk_n983 ) );
  OAI22_X1 u1_uk_U823 (.ZN( u1_K10_18 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1620 ) , .B2( u1_uk_n1634 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U843 (.ZN( u1_K1_6 ) , .B2( u1_uk_n1198 ) , .A2( u1_uk_n1205 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n240 ) );
  INV_X1 u1_uk_U844 (.A( u1_key_r_41 ) , .ZN( u1_uk_n1205 ) );
  OAI21_X1 u1_uk_U847 (.ZN( u1_K13_3 ) , .B2( u1_uk_n1781 ) , .B1( u1_uk_n27 ) , .A( u1_uk_n945 ) );
  NAND2_X1 u1_uk_U848 (.A1( u1_uk_K_r11_4 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n945 ) );
  OAI21_X1 u1_uk_U861 (.ZN( u1_K10_1 ) , .B2( u1_uk_n1630 ) , .A( u1_uk_n306 ) , .B1( u1_uk_n31 ) );
  NAND2_X1 u1_uk_U862 (.A1( u1_uk_K_r8_10 ) , .A2( u1_uk_n118 ) , .ZN( u1_uk_n306 ) );
  OAI22_X1 u1_uk_U863 (.ZN( u1_K1_1 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1204 ) , .A2( u1_uk_n1209 ) , .B1( u1_uk_n240 ) );
  AOI22_X1 u1_uk_U865 (.B2( u1_uk_K_r11_19 ) , .A2( u1_uk_K_r11_24 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) , .ZN( u1_uk_n949 ) );
  OAI22_X1 u1_uk_U868 (.ZN( u1_K10_5 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1625 ) , .A2( u1_uk_n1642 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U892 (.ZN( u1_K10_3 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1633 ) , .A2( u1_uk_n1653 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U899 (.ZN( u1_K13_24 ) , .B2( u1_uk_n1756 ) , .A2( u1_uk_n1797 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U916 (.ZN( u1_K2_17 ) , .A2( u1_uk_n1261 ) , .B2( u1_uk_n1277 ) , .A1( u1_uk_n291 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U928 (.ZN( u1_K13_23 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1767 ) , .A2( u1_uk_n1797 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U932 (.ZN( u1_K11_16 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1692 ) , .A2( u1_uk_n1698 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U934 (.ZN( u1_K11_6 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1699 ) , .A2( u1_uk_n1705 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U951 (.ZN( u1_K13_4 ) , .A1( u1_uk_n155 ) , .B2( u1_uk_n1762 ) , .A2( u1_uk_n1767 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U955 (.ZN( u1_K10_8 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1621 ) , .B2( u1_uk_n1635 ) , .B1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U956 (.ZN( u1_K13_8 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1781 ) , .A2( u1_uk_n1787 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U958 (.ZN( u1_K11_18 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1667 ) , .A2( u1_uk_n1673 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U990 (.ZN( u1_K1_23 ) , .B2( u1_uk_n1197 ) , .A2( u1_uk_n1204 ) , .A1( u1_uk_n128 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U993 (.ZN( u1_K1_3 ) , .B2( u1_uk_n1184 ) , .A2( u1_uk_n1191 ) , .A1( u1_uk_n128 ) , .B1( u1_uk_n238 ) );
  XOR2_X1 u2_U16 (.B( u2_L1_24 ) , .Z( u2_N87 ) , .A( u2_out2_24 ) );
  XOR2_X1 u2_U17 (.B( u2_L1_23 ) , .Z( u2_N86 ) , .A( u2_out2_23 ) );
  XOR2_X1 u2_U23 (.B( u2_L1_17 ) , .Z( u2_N80 ) , .A( u2_out2_17 ) );
  XOR2_X1 u2_U25 (.B( u2_L1_16 ) , .Z( u2_N79 ) , .A( u2_out2_16 ) );
  XOR2_X1 u2_U32 (.B( u2_L1_9 ) , .Z( u2_N72 ) , .A( u2_out2_9 ) );
  XOR2_X1 u2_U36 (.B( u2_L1_6 ) , .Z( u2_N69 ) , .A( u2_out2_6 ) );
  XOR2_X1 u2_U484 (.Z( u2_FP_8 ) , .B( u2_L14_8 ) , .A( u2_out15_8 ) );
  XOR2_X1 u2_U489 (.Z( u2_FP_3 ) , .B( u2_L14_3 ) , .A( u2_out15_3 ) );
  XOR2_X1 u2_U498 (.Z( u2_FP_25 ) , .B( u2_L14_25 ) , .A( u2_out15_25 ) );
  XOR2_X1 u2_U510 (.Z( u2_FP_14 ) , .B( u2_L14_14 ) , .A( u2_out15_14 ) );
  XOR2_X1 u2_U8 (.B( u2_L1_31 ) , .Z( u2_N94 ) , .A( u2_out2_31 ) );
  XOR2_X1 u2_U9 (.B( u2_L1_30 ) , .Z( u2_N93 ) , .A( u2_out2_30 ) );
  XOR2_X1 u2_u15_U26 (.A( u2_FP_53 ) , .B( u2_K16_30 ) , .Z( u2_u15_X_30 ) );
  XOR2_X1 u2_u15_U28 (.A( u2_FP_52 ) , .B( u2_K16_29 ) , .Z( u2_u15_X_29 ) );
  XOR2_X1 u2_u15_U29 (.A( u2_FP_51 ) , .B( u2_K16_28 ) , .Z( u2_u15_X_28 ) );
  XOR2_X1 u2_u15_U30 (.A( u2_FP_50 ) , .B( u2_K16_27 ) , .Z( u2_u15_X_27 ) );
  XOR2_X1 u2_u15_U31 (.A( u2_FP_49 ) , .B( u2_K16_26 ) , .Z( u2_u15_X_26 ) );
  XOR2_X1 u2_u15_U32 (.A( u2_FP_48 ) , .B( u2_K16_25 ) , .Z( u2_u15_X_25 ) );
  OAI22_X1 u2_u15_u4_U10 (.B2( u2_u15_u4_n135 ) , .ZN( u2_u15_u4_n137 ) , .B1( u2_u15_u4_n153 ) , .A1( u2_u15_u4_n155 ) , .A2( u2_u15_u4_n171 ) );
  AND3_X1 u2_u15_u4_U11 (.A2( u2_u15_u4_n134 ) , .ZN( u2_u15_u4_n135 ) , .A3( u2_u15_u4_n145 ) , .A1( u2_u15_u4_n157 ) );
  OR3_X1 u2_u15_u4_U12 (.A3( u2_u15_u4_n114 ) , .A2( u2_u15_u4_n115 ) , .A1( u2_u15_u4_n116 ) , .ZN( u2_u15_u4_n136 ) );
  AOI21_X1 u2_u15_u4_U13 (.A( u2_u15_u4_n113 ) , .ZN( u2_u15_u4_n116 ) , .B2( u2_u15_u4_n173 ) , .B1( u2_u15_u4_n174 ) );
  AOI21_X1 u2_u15_u4_U14 (.ZN( u2_u15_u4_n115 ) , .B2( u2_u15_u4_n145 ) , .B1( u2_u15_u4_n146 ) , .A( u2_u15_u4_n156 ) );
  OAI22_X1 u2_u15_u4_U15 (.ZN( u2_u15_u4_n114 ) , .A2( u2_u15_u4_n121 ) , .B1( u2_u15_u4_n160 ) , .B2( u2_u15_u4_n170 ) , .A1( u2_u15_u4_n171 ) );
  NAND2_X1 u2_u15_u4_U16 (.ZN( u2_u15_u4_n132 ) , .A2( u2_u15_u4_n170 ) , .A1( u2_u15_u4_n173 ) );
  AOI21_X1 u2_u15_u4_U17 (.B2( u2_u15_u4_n160 ) , .B1( u2_u15_u4_n161 ) , .ZN( u2_u15_u4_n162 ) , .A( u2_u15_u4_n170 ) );
  AOI21_X1 u2_u15_u4_U18 (.ZN( u2_u15_u4_n107 ) , .B2( u2_u15_u4_n143 ) , .A( u2_u15_u4_n174 ) , .B1( u2_u15_u4_n184 ) );
  AOI21_X1 u2_u15_u4_U19 (.B2( u2_u15_u4_n158 ) , .B1( u2_u15_u4_n159 ) , .ZN( u2_u15_u4_n163 ) , .A( u2_u15_u4_n174 ) );
  AOI21_X1 u2_u15_u4_U20 (.A( u2_u15_u4_n153 ) , .B2( u2_u15_u4_n154 ) , .B1( u2_u15_u4_n155 ) , .ZN( u2_u15_u4_n165 ) );
  AOI21_X1 u2_u15_u4_U21 (.A( u2_u15_u4_n156 ) , .B2( u2_u15_u4_n157 ) , .ZN( u2_u15_u4_n164 ) , .B1( u2_u15_u4_n184 ) );
  INV_X1 u2_u15_u4_U22 (.A( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n170 ) );
  AND2_X1 u2_u15_u4_U23 (.A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n155 ) , .A1( u2_u15_u4_n160 ) );
  INV_X1 u2_u15_u4_U24 (.A( u2_u15_u4_n156 ) , .ZN( u2_u15_u4_n175 ) );
  NAND2_X1 u2_u15_u4_U25 (.A2( u2_u15_u4_n118 ) , .ZN( u2_u15_u4_n131 ) , .A1( u2_u15_u4_n147 ) );
  NAND2_X1 u2_u15_u4_U26 (.A1( u2_u15_u4_n119 ) , .A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n130 ) );
  NAND2_X1 u2_u15_u4_U27 (.ZN( u2_u15_u4_n117 ) , .A2( u2_u15_u4_n118 ) , .A1( u2_u15_u4_n148 ) );
  NAND2_X1 u2_u15_u4_U28 (.ZN( u2_u15_u4_n129 ) , .A1( u2_u15_u4_n134 ) , .A2( u2_u15_u4_n148 ) );
  AND3_X1 u2_u15_u4_U29 (.A1( u2_u15_u4_n119 ) , .A2( u2_u15_u4_n143 ) , .A3( u2_u15_u4_n154 ) , .ZN( u2_u15_u4_n161 ) );
  NOR2_X1 u2_u15_u4_U3 (.ZN( u2_u15_u4_n121 ) , .A1( u2_u15_u4_n181 ) , .A2( u2_u15_u4_n182 ) );
  AND2_X1 u2_u15_u4_U30 (.A1( u2_u15_u4_n145 ) , .A2( u2_u15_u4_n147 ) , .ZN( u2_u15_u4_n159 ) );
  INV_X1 u2_u15_u4_U31 (.A( u2_u15_u4_n158 ) , .ZN( u2_u15_u4_n182 ) );
  INV_X1 u2_u15_u4_U32 (.ZN( u2_u15_u4_n181 ) , .A( u2_u15_u4_n96 ) );
  INV_X1 u2_u15_u4_U33 (.A( u2_u15_u4_n144 ) , .ZN( u2_u15_u4_n179 ) );
  INV_X1 u2_u15_u4_U34 (.A( u2_u15_u4_n157 ) , .ZN( u2_u15_u4_n178 ) );
  NAND2_X1 u2_u15_u4_U35 (.A2( u2_u15_u4_n154 ) , .A1( u2_u15_u4_n96 ) , .ZN( u2_u15_u4_n97 ) );
  INV_X1 u2_u15_u4_U36 (.ZN( u2_u15_u4_n186 ) , .A( u2_u15_u4_n95 ) );
  OAI221_X1 u2_u15_u4_U37 (.C1( u2_u15_u4_n134 ) , .B1( u2_u15_u4_n158 ) , .B2( u2_u15_u4_n171 ) , .C2( u2_u15_u4_n173 ) , .A( u2_u15_u4_n94 ) , .ZN( u2_u15_u4_n95 ) );
  AOI222_X1 u2_u15_u4_U38 (.B2( u2_u15_u4_n132 ) , .A1( u2_u15_u4_n138 ) , .C2( u2_u15_u4_n175 ) , .A2( u2_u15_u4_n179 ) , .C1( u2_u15_u4_n181 ) , .B1( u2_u15_u4_n185 ) , .ZN( u2_u15_u4_n94 ) );
  INV_X1 u2_u15_u4_U39 (.A( u2_u15_u4_n113 ) , .ZN( u2_u15_u4_n185 ) );
  INV_X1 u2_u15_u4_U4 (.A( u2_u15_u4_n117 ) , .ZN( u2_u15_u4_n184 ) );
  INV_X1 u2_u15_u4_U40 (.A( u2_u15_u4_n143 ) , .ZN( u2_u15_u4_n183 ) );
  NOR2_X1 u2_u15_u4_U41 (.ZN( u2_u15_u4_n138 ) , .A1( u2_u15_u4_n168 ) , .A2( u2_u15_u4_n169 ) );
  NOR2_X1 u2_u15_u4_U42 (.A1( u2_u15_u4_n150 ) , .A2( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n153 ) );
  NOR2_X1 u2_u15_u4_U43 (.A2( u2_u15_u4_n128 ) , .A1( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n156 ) );
  AOI22_X1 u2_u15_u4_U44 (.B2( u2_u15_u4_n122 ) , .A1( u2_u15_u4_n123 ) , .ZN( u2_u15_u4_n124 ) , .B1( u2_u15_u4_n128 ) , .A2( u2_u15_u4_n172 ) );
  NAND2_X1 u2_u15_u4_U45 (.A2( u2_u15_u4_n120 ) , .ZN( u2_u15_u4_n123 ) , .A1( u2_u15_u4_n161 ) );
  INV_X1 u2_u15_u4_U46 (.A( u2_u15_u4_n153 ) , .ZN( u2_u15_u4_n172 ) );
  AOI22_X1 u2_u15_u4_U47 (.B2( u2_u15_u4_n132 ) , .A2( u2_u15_u4_n133 ) , .ZN( u2_u15_u4_n140 ) , .A1( u2_u15_u4_n150 ) , .B1( u2_u15_u4_n179 ) );
  NAND2_X1 u2_u15_u4_U48 (.ZN( u2_u15_u4_n133 ) , .A2( u2_u15_u4_n146 ) , .A1( u2_u15_u4_n154 ) );
  NAND2_X1 u2_u15_u4_U49 (.A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n154 ) , .A2( u2_u15_u4_n98 ) );
  NOR4_X1 u2_u15_u4_U5 (.A4( u2_u15_u4_n106 ) , .A3( u2_u15_u4_n107 ) , .A2( u2_u15_u4_n108 ) , .A1( u2_u15_u4_n109 ) , .ZN( u2_u15_u4_n110 ) );
  NAND2_X1 u2_u15_u4_U50 (.A1( u2_u15_u4_n101 ) , .ZN( u2_u15_u4_n158 ) , .A2( u2_u15_u4_n99 ) );
  AOI21_X1 u2_u15_u4_U51 (.ZN( u2_u15_u4_n127 ) , .A( u2_u15_u4_n136 ) , .B2( u2_u15_u4_n150 ) , .B1( u2_u15_u4_n180 ) );
  INV_X1 u2_u15_u4_U52 (.A( u2_u15_u4_n160 ) , .ZN( u2_u15_u4_n180 ) );
  NAND2_X1 u2_u15_u4_U53 (.A2( u2_u15_u4_n104 ) , .A1( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n146 ) );
  NAND2_X1 u2_u15_u4_U54 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n160 ) );
  NAND2_X1 u2_u15_u4_U55 (.ZN( u2_u15_u4_n134 ) , .A1( u2_u15_u4_n98 ) , .A2( u2_u15_u4_n99 ) );
  NAND2_X1 u2_u15_u4_U56 (.A1( u2_u15_u4_n103 ) , .A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n143 ) );
  NAND2_X1 u2_u15_u4_U57 (.A2( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n145 ) , .A1( u2_u15_u4_n98 ) );
  NAND2_X1 u2_u15_u4_U58 (.A1( u2_u15_u4_n100 ) , .A2( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n120 ) );
  NAND2_X1 u2_u15_u4_U59 (.A1( u2_u15_u4_n102 ) , .A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n148 ) );
  AOI21_X1 u2_u15_u4_U6 (.ZN( u2_u15_u4_n106 ) , .B2( u2_u15_u4_n146 ) , .B1( u2_u15_u4_n158 ) , .A( u2_u15_u4_n170 ) );
  NAND2_X1 u2_u15_u4_U60 (.A2( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n157 ) );
  INV_X1 u2_u15_u4_U61 (.A( u2_u15_u4_n150 ) , .ZN( u2_u15_u4_n173 ) );
  INV_X1 u2_u15_u4_U62 (.A( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n171 ) );
  NAND2_X1 u2_u15_u4_U63 (.A1( u2_u15_u4_n100 ) , .ZN( u2_u15_u4_n118 ) , .A2( u2_u15_u4_n99 ) );
  NAND2_X1 u2_u15_u4_U64 (.A2( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n144 ) );
  NAND2_X1 u2_u15_u4_U65 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n105 ) , .ZN( u2_u15_u4_n96 ) );
  INV_X1 u2_u15_u4_U66 (.A( u2_u15_u4_n128 ) , .ZN( u2_u15_u4_n174 ) );
  NAND2_X1 u2_u15_u4_U67 (.A2( u2_u15_u4_n102 ) , .ZN( u2_u15_u4_n119 ) , .A1( u2_u15_u4_n98 ) );
  NAND2_X1 u2_u15_u4_U68 (.A2( u2_u15_u4_n101 ) , .A1( u2_u15_u4_n103 ) , .ZN( u2_u15_u4_n147 ) );
  NAND2_X1 u2_u15_u4_U69 (.A2( u2_u15_u4_n104 ) , .ZN( u2_u15_u4_n113 ) , .A1( u2_u15_u4_n99 ) );
  AOI21_X1 u2_u15_u4_U7 (.ZN( u2_u15_u4_n108 ) , .B2( u2_u15_u4_n134 ) , .B1( u2_u15_u4_n155 ) , .A( u2_u15_u4_n156 ) );
  NOR2_X1 u2_u15_u4_U70 (.A2( u2_u15_X_28 ) , .ZN( u2_u15_u4_n150 ) , .A1( u2_u15_u4_n168 ) );
  NOR2_X1 u2_u15_u4_U71 (.A2( u2_u15_X_29 ) , .ZN( u2_u15_u4_n152 ) , .A1( u2_u15_u4_n169 ) );
  NOR2_X1 u2_u15_u4_U72 (.A2( u2_u15_X_26 ) , .ZN( u2_u15_u4_n100 ) , .A1( u2_u15_u4_n177 ) );
  NOR2_X1 u2_u15_u4_U73 (.A2( u2_u15_X_30 ) , .ZN( u2_u15_u4_n105 ) , .A1( u2_u15_u4_n176 ) );
  NOR2_X1 u2_u15_u4_U74 (.A2( u2_u15_X_28 ) , .A1( u2_u15_X_29 ) , .ZN( u2_u15_u4_n128 ) );
  NOR2_X1 u2_u15_u4_U75 (.A2( u2_u15_X_25 ) , .A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n98 ) );
  NOR2_X1 u2_u15_u4_U76 (.A2( u2_u15_X_27 ) , .A1( u2_u15_X_30 ) , .ZN( u2_u15_u4_n102 ) );
  AND2_X1 u2_u15_u4_U77 (.A2( u2_u15_X_25 ) , .A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n104 ) );
  AND2_X1 u2_u15_u4_U78 (.A1( u2_u15_X_30 ) , .A2( u2_u15_u4_n176 ) , .ZN( u2_u15_u4_n99 ) );
  AND2_X1 u2_u15_u4_U79 (.A1( u2_u15_X_26 ) , .ZN( u2_u15_u4_n101 ) , .A2( u2_u15_u4_n177 ) );
  AOI21_X1 u2_u15_u4_U8 (.ZN( u2_u15_u4_n109 ) , .A( u2_u15_u4_n153 ) , .B1( u2_u15_u4_n159 ) , .B2( u2_u15_u4_n184 ) );
  AND2_X1 u2_u15_u4_U80 (.A1( u2_u15_X_27 ) , .A2( u2_u15_X_30 ) , .ZN( u2_u15_u4_n103 ) );
  INV_X1 u2_u15_u4_U81 (.A( u2_u15_X_28 ) , .ZN( u2_u15_u4_n169 ) );
  INV_X1 u2_u15_u4_U82 (.A( u2_u15_X_29 ) , .ZN( u2_u15_u4_n168 ) );
  INV_X1 u2_u15_u4_U83 (.A( u2_u15_X_25 ) , .ZN( u2_u15_u4_n177 ) );
  INV_X1 u2_u15_u4_U84 (.A( u2_u15_X_27 ) , .ZN( u2_u15_u4_n176 ) );
  NAND4_X1 u2_u15_u4_U85 (.ZN( u2_out15_14 ) , .A4( u2_u15_u4_n124 ) , .A3( u2_u15_u4_n125 ) , .A2( u2_u15_u4_n126 ) , .A1( u2_u15_u4_n127 ) );
  AOI22_X1 u2_u15_u4_U86 (.B2( u2_u15_u4_n117 ) , .ZN( u2_u15_u4_n126 ) , .A1( u2_u15_u4_n129 ) , .B1( u2_u15_u4_n152 ) , .A2( u2_u15_u4_n175 ) );
  AOI22_X1 u2_u15_u4_U87 (.ZN( u2_u15_u4_n125 ) , .B2( u2_u15_u4_n131 ) , .A2( u2_u15_u4_n132 ) , .B1( u2_u15_u4_n138 ) , .A1( u2_u15_u4_n178 ) );
  AOI22_X1 u2_u15_u4_U88 (.B2( u2_u15_u4_n149 ) , .B1( u2_u15_u4_n150 ) , .A2( u2_u15_u4_n151 ) , .A1( u2_u15_u4_n152 ) , .ZN( u2_u15_u4_n167 ) );
  NOR4_X1 u2_u15_u4_U89 (.A4( u2_u15_u4_n162 ) , .A3( u2_u15_u4_n163 ) , .A2( u2_u15_u4_n164 ) , .A1( u2_u15_u4_n165 ) , .ZN( u2_u15_u4_n166 ) );
  AOI211_X1 u2_u15_u4_U9 (.B( u2_u15_u4_n136 ) , .A( u2_u15_u4_n137 ) , .C2( u2_u15_u4_n138 ) , .ZN( u2_u15_u4_n139 ) , .C1( u2_u15_u4_n182 ) );
  NAND4_X1 u2_u15_u4_U90 (.ZN( u2_out15_8 ) , .A4( u2_u15_u4_n110 ) , .A3( u2_u15_u4_n111 ) , .A2( u2_u15_u4_n112 ) , .A1( u2_u15_u4_n186 ) );
  NAND2_X1 u2_u15_u4_U91 (.ZN( u2_u15_u4_n112 ) , .A2( u2_u15_u4_n130 ) , .A1( u2_u15_u4_n150 ) );
  AOI22_X1 u2_u15_u4_U92 (.ZN( u2_u15_u4_n111 ) , .B2( u2_u15_u4_n132 ) , .A1( u2_u15_u4_n152 ) , .B1( u2_u15_u4_n178 ) , .A2( u2_u15_u4_n97 ) );
  NAND4_X1 u2_u15_u4_U93 (.ZN( u2_out15_25 ) , .A4( u2_u15_u4_n139 ) , .A3( u2_u15_u4_n140 ) , .A2( u2_u15_u4_n141 ) , .A1( u2_u15_u4_n142 ) );
  OAI21_X1 u2_u15_u4_U94 (.A( u2_u15_u4_n128 ) , .B2( u2_u15_u4_n129 ) , .B1( u2_u15_u4_n130 ) , .ZN( u2_u15_u4_n142 ) );
  OAI21_X1 u2_u15_u4_U95 (.B2( u2_u15_u4_n131 ) , .ZN( u2_u15_u4_n141 ) , .A( u2_u15_u4_n175 ) , .B1( u2_u15_u4_n183 ) );
  NAND3_X1 u2_u15_u4_U96 (.ZN( u2_out15_3 ) , .A3( u2_u15_u4_n166 ) , .A1( u2_u15_u4_n167 ) , .A2( u2_u15_u4_n186 ) );
  NAND3_X1 u2_u15_u4_U97 (.A3( u2_u15_u4_n146 ) , .A2( u2_u15_u4_n147 ) , .A1( u2_u15_u4_n148 ) , .ZN( u2_u15_u4_n149 ) );
  NAND3_X1 u2_u15_u4_U98 (.A3( u2_u15_u4_n143 ) , .A2( u2_u15_u4_n144 ) , .A1( u2_u15_u4_n145 ) , .ZN( u2_u15_u4_n151 ) );
  NAND3_X1 u2_u15_u4_U99 (.A3( u2_u15_u4_n121 ) , .ZN( u2_u15_u4_n122 ) , .A2( u2_u15_u4_n144 ) , .A1( u2_u15_u4_n154 ) );
  XOR2_X1 u2_u2_U16 (.B( u2_K3_3 ) , .A( u2_R1_2 ) , .Z( u2_u2_X_3 ) );
  XOR2_X1 u2_u2_U27 (.B( u2_K3_2 ) , .A( u2_R1_1 ) , .Z( u2_u2_X_2 ) );
  XOR2_X1 u2_u2_U38 (.B( u2_K3_1 ) , .A( u2_R1_32 ) , .Z( u2_u2_X_1 ) );
  XOR2_X1 u2_u2_U4 (.B( u2_K3_6 ) , .A( u2_R1_5 ) , .Z( u2_u2_X_6 ) );
  XOR2_X1 u2_u2_U40 (.B( u2_K3_18 ) , .A( u2_R1_13 ) , .Z( u2_u2_X_18 ) );
  XOR2_X1 u2_u2_U41 (.B( u2_K3_17 ) , .A( u2_R1_12 ) , .Z( u2_u2_X_17 ) );
  XOR2_X1 u2_u2_U42 (.B( u2_K3_16 ) , .A( u2_R1_11 ) , .Z( u2_u2_X_16 ) );
  XOR2_X1 u2_u2_U43 (.B( u2_K3_15 ) , .A( u2_R1_10 ) , .Z( u2_u2_X_15 ) );
  XOR2_X1 u2_u2_U44 (.B( u2_K3_14 ) , .A( u2_R1_9 ) , .Z( u2_u2_X_14 ) );
  XOR2_X1 u2_u2_U45 (.B( u2_K3_13 ) , .A( u2_R1_8 ) , .Z( u2_u2_X_13 ) );
  XOR2_X1 u2_u2_U5 (.B( u2_K3_5 ) , .A( u2_R1_4 ) , .Z( u2_u2_X_5 ) );
  XOR2_X1 u2_u2_U6 (.B( u2_K3_4 ) , .A( u2_R1_3 ) , .Z( u2_u2_X_4 ) );
  AND3_X1 u2_u2_u0_U10 (.A2( u2_u2_u0_n112 ) , .ZN( u2_u2_u0_n127 ) , .A3( u2_u2_u0_n130 ) , .A1( u2_u2_u0_n148 ) );
  NAND2_X1 u2_u2_u0_U11 (.ZN( u2_u2_u0_n113 ) , .A1( u2_u2_u0_n139 ) , .A2( u2_u2_u0_n149 ) );
  AND2_X1 u2_u2_u0_U12 (.ZN( u2_u2_u0_n107 ) , .A1( u2_u2_u0_n130 ) , .A2( u2_u2_u0_n140 ) );
  AND2_X1 u2_u2_u0_U13 (.A2( u2_u2_u0_n129 ) , .A1( u2_u2_u0_n130 ) , .ZN( u2_u2_u0_n151 ) );
  AND2_X1 u2_u2_u0_U14 (.A1( u2_u2_u0_n108 ) , .A2( u2_u2_u0_n125 ) , .ZN( u2_u2_u0_n145 ) );
  INV_X1 u2_u2_u0_U15 (.A( u2_u2_u0_n143 ) , .ZN( u2_u2_u0_n173 ) );
  NOR2_X1 u2_u2_u0_U16 (.A2( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n147 ) , .A1( u2_u2_u0_n160 ) );
  INV_X1 u2_u2_u0_U17 (.ZN( u2_u2_u0_n172 ) , .A( u2_u2_u0_n88 ) );
  OAI222_X1 u2_u2_u0_U18 (.C1( u2_u2_u0_n108 ) , .A1( u2_u2_u0_n125 ) , .B2( u2_u2_u0_n128 ) , .B1( u2_u2_u0_n144 ) , .A2( u2_u2_u0_n158 ) , .C2( u2_u2_u0_n161 ) , .ZN( u2_u2_u0_n88 ) );
  NOR2_X1 u2_u2_u0_U19 (.A1( u2_u2_u0_n163 ) , .A2( u2_u2_u0_n164 ) , .ZN( u2_u2_u0_n95 ) );
  AOI21_X1 u2_u2_u0_U20 (.B1( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n132 ) , .A( u2_u2_u0_n165 ) , .B2( u2_u2_u0_n93 ) );
  INV_X1 u2_u2_u0_U21 (.A( u2_u2_u0_n142 ) , .ZN( u2_u2_u0_n165 ) );
  OAI221_X1 u2_u2_u0_U22 (.C1( u2_u2_u0_n121 ) , .ZN( u2_u2_u0_n122 ) , .B2( u2_u2_u0_n127 ) , .A( u2_u2_u0_n143 ) , .B1( u2_u2_u0_n144 ) , .C2( u2_u2_u0_n147 ) );
  OAI22_X1 u2_u2_u0_U23 (.B1( u2_u2_u0_n125 ) , .ZN( u2_u2_u0_n126 ) , .A1( u2_u2_u0_n138 ) , .A2( u2_u2_u0_n146 ) , .B2( u2_u2_u0_n147 ) );
  OAI22_X1 u2_u2_u0_U24 (.B1( u2_u2_u0_n131 ) , .A1( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n147 ) , .A2( u2_u2_u0_n90 ) , .ZN( u2_u2_u0_n91 ) );
  AND3_X1 u2_u2_u0_U25 (.A3( u2_u2_u0_n121 ) , .A2( u2_u2_u0_n125 ) , .A1( u2_u2_u0_n148 ) , .ZN( u2_u2_u0_n90 ) );
  INV_X1 u2_u2_u0_U26 (.A( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n161 ) );
  NOR2_X1 u2_u2_u0_U27 (.A1( u2_u2_u0_n120 ) , .ZN( u2_u2_u0_n143 ) , .A2( u2_u2_u0_n167 ) );
  OAI221_X1 u2_u2_u0_U28 (.C1( u2_u2_u0_n112 ) , .ZN( u2_u2_u0_n120 ) , .B1( u2_u2_u0_n138 ) , .B2( u2_u2_u0_n141 ) , .C2( u2_u2_u0_n147 ) , .A( u2_u2_u0_n172 ) );
  AOI211_X1 u2_u2_u0_U29 (.B( u2_u2_u0_n115 ) , .A( u2_u2_u0_n116 ) , .C2( u2_u2_u0_n117 ) , .C1( u2_u2_u0_n118 ) , .ZN( u2_u2_u0_n119 ) );
  INV_X1 u2_u2_u0_U3 (.A( u2_u2_u0_n113 ) , .ZN( u2_u2_u0_n166 ) );
  AOI22_X1 u2_u2_u0_U30 (.B2( u2_u2_u0_n109 ) , .A2( u2_u2_u0_n110 ) , .ZN( u2_u2_u0_n111 ) , .B1( u2_u2_u0_n118 ) , .A1( u2_u2_u0_n160 ) );
  INV_X1 u2_u2_u0_U31 (.A( u2_u2_u0_n118 ) , .ZN( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U32 (.ZN( u2_u2_u0_n104 ) , .B1( u2_u2_u0_n107 ) , .B2( u2_u2_u0_n141 ) , .A( u2_u2_u0_n144 ) );
  AOI21_X1 u2_u2_u0_U33 (.B1( u2_u2_u0_n127 ) , .B2( u2_u2_u0_n129 ) , .A( u2_u2_u0_n138 ) , .ZN( u2_u2_u0_n96 ) );
  AOI21_X1 u2_u2_u0_U34 (.ZN( u2_u2_u0_n116 ) , .B2( u2_u2_u0_n142 ) , .A( u2_u2_u0_n144 ) , .B1( u2_u2_u0_n166 ) );
  NAND2_X1 u2_u2_u0_U35 (.A1( u2_u2_u0_n100 ) , .A2( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n125 ) );
  NAND2_X1 u2_u2_u0_U36 (.A1( u2_u2_u0_n101 ) , .A2( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n150 ) );
  INV_X1 u2_u2_u0_U37 (.A( u2_u2_u0_n138 ) , .ZN( u2_u2_u0_n160 ) );
  NAND2_X1 u2_u2_u0_U38 (.A1( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n128 ) , .A2( u2_u2_u0_n95 ) );
  NAND2_X1 u2_u2_u0_U39 (.A1( u2_u2_u0_n100 ) , .ZN( u2_u2_u0_n129 ) , .A2( u2_u2_u0_n95 ) );
  AOI21_X1 u2_u2_u0_U4 (.B1( u2_u2_u0_n114 ) , .ZN( u2_u2_u0_n115 ) , .B2( u2_u2_u0_n129 ) , .A( u2_u2_u0_n161 ) );
  NAND2_X1 u2_u2_u0_U40 (.A2( u2_u2_u0_n100 ) , .ZN( u2_u2_u0_n131 ) , .A1( u2_u2_u0_n92 ) );
  NAND2_X1 u2_u2_u0_U41 (.A2( u2_u2_u0_n100 ) , .A1( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n139 ) );
  NAND2_X1 u2_u2_u0_U42 (.ZN( u2_u2_u0_n148 ) , .A1( u2_u2_u0_n93 ) , .A2( u2_u2_u0_n95 ) );
  NAND2_X1 u2_u2_u0_U43 (.A2( u2_u2_u0_n102 ) , .A1( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n149 ) );
  NAND2_X1 u2_u2_u0_U44 (.A2( u2_u2_u0_n102 ) , .ZN( u2_u2_u0_n114 ) , .A1( u2_u2_u0_n92 ) );
  NAND2_X1 u2_u2_u0_U45 (.A2( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n121 ) , .A1( u2_u2_u0_n93 ) );
  NAND2_X1 u2_u2_u0_U46 (.ZN( u2_u2_u0_n112 ) , .A2( u2_u2_u0_n92 ) , .A1( u2_u2_u0_n93 ) );
  OR3_X1 u2_u2_u0_U47 (.A3( u2_u2_u0_n152 ) , .A2( u2_u2_u0_n153 ) , .A1( u2_u2_u0_n154 ) , .ZN( u2_u2_u0_n155 ) );
  AOI21_X1 u2_u2_u0_U48 (.B2( u2_u2_u0_n150 ) , .B1( u2_u2_u0_n151 ) , .ZN( u2_u2_u0_n152 ) , .A( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U49 (.A( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n145 ) , .B1( u2_u2_u0_n146 ) , .ZN( u2_u2_u0_n154 ) );
  AOI21_X1 u2_u2_u0_U5 (.B2( u2_u2_u0_n131 ) , .ZN( u2_u2_u0_n134 ) , .B1( u2_u2_u0_n151 ) , .A( u2_u2_u0_n158 ) );
  AOI21_X1 u2_u2_u0_U50 (.A( u2_u2_u0_n147 ) , .B2( u2_u2_u0_n148 ) , .B1( u2_u2_u0_n149 ) , .ZN( u2_u2_u0_n153 ) );
  INV_X1 u2_u2_u0_U51 (.ZN( u2_u2_u0_n171 ) , .A( u2_u2_u0_n99 ) );
  OAI211_X1 u2_u2_u0_U52 (.C2( u2_u2_u0_n140 ) , .C1( u2_u2_u0_n161 ) , .A( u2_u2_u0_n169 ) , .B( u2_u2_u0_n98 ) , .ZN( u2_u2_u0_n99 ) );
  INV_X1 u2_u2_u0_U53 (.ZN( u2_u2_u0_n169 ) , .A( u2_u2_u0_n91 ) );
  AOI211_X1 u2_u2_u0_U54 (.C1( u2_u2_u0_n118 ) , .A( u2_u2_u0_n123 ) , .B( u2_u2_u0_n96 ) , .C2( u2_u2_u0_n97 ) , .ZN( u2_u2_u0_n98 ) );
  NOR2_X1 u2_u2_u0_U55 (.A2( u2_u2_X_6 ) , .ZN( u2_u2_u0_n100 ) , .A1( u2_u2_u0_n162 ) );
  NOR2_X1 u2_u2_u0_U56 (.A2( u2_u2_X_4 ) , .A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n118 ) );
  NOR2_X1 u2_u2_u0_U57 (.A2( u2_u2_X_2 ) , .ZN( u2_u2_u0_n103 ) , .A1( u2_u2_u0_n164 ) );
  NOR2_X1 u2_u2_u0_U58 (.A2( u2_u2_X_1 ) , .A1( u2_u2_X_2 ) , .ZN( u2_u2_u0_n92 ) );
  NOR2_X1 u2_u2_u0_U59 (.A2( u2_u2_X_1 ) , .ZN( u2_u2_u0_n101 ) , .A1( u2_u2_u0_n163 ) );
  NOR2_X1 u2_u2_u0_U6 (.A1( u2_u2_u0_n108 ) , .ZN( u2_u2_u0_n123 ) , .A2( u2_u2_u0_n158 ) );
  NAND2_X1 u2_u2_u0_U60 (.A2( u2_u2_X_4 ) , .A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n144 ) );
  NOR2_X1 u2_u2_u0_U61 (.A2( u2_u2_X_5 ) , .ZN( u2_u2_u0_n136 ) , .A1( u2_u2_u0_n159 ) );
  NAND2_X1 u2_u2_u0_U62 (.A1( u2_u2_X_5 ) , .ZN( u2_u2_u0_n138 ) , .A2( u2_u2_u0_n159 ) );
  NOR2_X1 u2_u2_u0_U63 (.A2( u2_u2_X_3 ) , .A1( u2_u2_X_6 ) , .ZN( u2_u2_u0_n94 ) );
  AND2_X1 u2_u2_u0_U64 (.A2( u2_u2_X_3 ) , .A1( u2_u2_X_6 ) , .ZN( u2_u2_u0_n102 ) );
  AND2_X1 u2_u2_u0_U65 (.A1( u2_u2_X_6 ) , .A2( u2_u2_u0_n162 ) , .ZN( u2_u2_u0_n93 ) );
  INV_X1 u2_u2_u0_U66 (.A( u2_u2_X_4 ) , .ZN( u2_u2_u0_n159 ) );
  INV_X1 u2_u2_u0_U67 (.A( u2_u2_X_1 ) , .ZN( u2_u2_u0_n164 ) );
  INV_X1 u2_u2_u0_U68 (.A( u2_u2_X_2 ) , .ZN( u2_u2_u0_n163 ) );
  INV_X1 u2_u2_u0_U69 (.A( u2_u2_X_3 ) , .ZN( u2_u2_u0_n162 ) );
  OAI21_X1 u2_u2_u0_U7 (.B1( u2_u2_u0_n150 ) , .B2( u2_u2_u0_n158 ) , .A( u2_u2_u0_n172 ) , .ZN( u2_u2_u0_n89 ) );
  INV_X1 u2_u2_u0_U70 (.A( u2_u2_u0_n126 ) , .ZN( u2_u2_u0_n168 ) );
  AOI211_X1 u2_u2_u0_U71 (.B( u2_u2_u0_n133 ) , .A( u2_u2_u0_n134 ) , .C2( u2_u2_u0_n135 ) , .C1( u2_u2_u0_n136 ) , .ZN( u2_u2_u0_n137 ) );
  INV_X1 u2_u2_u0_U72 (.ZN( u2_u2_u0_n174 ) , .A( u2_u2_u0_n89 ) );
  AOI211_X1 u2_u2_u0_U73 (.B( u2_u2_u0_n104 ) , .A( u2_u2_u0_n105 ) , .ZN( u2_u2_u0_n106 ) , .C2( u2_u2_u0_n113 ) , .C1( u2_u2_u0_n160 ) );
  OR4_X1 u2_u2_u0_U74 (.ZN( u2_out2_17 ) , .A4( u2_u2_u0_n122 ) , .A2( u2_u2_u0_n123 ) , .A1( u2_u2_u0_n124 ) , .A3( u2_u2_u0_n170 ) );
  AOI21_X1 u2_u2_u0_U75 (.B2( u2_u2_u0_n107 ) , .ZN( u2_u2_u0_n124 ) , .B1( u2_u2_u0_n128 ) , .A( u2_u2_u0_n161 ) );
  INV_X1 u2_u2_u0_U76 (.A( u2_u2_u0_n111 ) , .ZN( u2_u2_u0_n170 ) );
  OR4_X1 u2_u2_u0_U77 (.ZN( u2_out2_31 ) , .A4( u2_u2_u0_n155 ) , .A2( u2_u2_u0_n156 ) , .A1( u2_u2_u0_n157 ) , .A3( u2_u2_u0_n173 ) );
  AOI21_X1 u2_u2_u0_U78 (.A( u2_u2_u0_n138 ) , .B2( u2_u2_u0_n139 ) , .B1( u2_u2_u0_n140 ) , .ZN( u2_u2_u0_n157 ) );
  AOI21_X1 u2_u2_u0_U79 (.B2( u2_u2_u0_n141 ) , .B1( u2_u2_u0_n142 ) , .ZN( u2_u2_u0_n156 ) , .A( u2_u2_u0_n161 ) );
  AND2_X1 u2_u2_u0_U8 (.A1( u2_u2_u0_n114 ) , .A2( u2_u2_u0_n121 ) , .ZN( u2_u2_u0_n146 ) );
  AOI21_X1 u2_u2_u0_U80 (.B1( u2_u2_u0_n132 ) , .ZN( u2_u2_u0_n133 ) , .A( u2_u2_u0_n144 ) , .B2( u2_u2_u0_n166 ) );
  OAI22_X1 u2_u2_u0_U81 (.ZN( u2_u2_u0_n105 ) , .A2( u2_u2_u0_n132 ) , .B1( u2_u2_u0_n146 ) , .A1( u2_u2_u0_n147 ) , .B2( u2_u2_u0_n161 ) );
  NAND2_X1 u2_u2_u0_U82 (.ZN( u2_u2_u0_n110 ) , .A2( u2_u2_u0_n132 ) , .A1( u2_u2_u0_n145 ) );
  INV_X1 u2_u2_u0_U83 (.A( u2_u2_u0_n119 ) , .ZN( u2_u2_u0_n167 ) );
  NAND2_X1 u2_u2_u0_U84 (.A2( u2_u2_u0_n103 ) , .ZN( u2_u2_u0_n140 ) , .A1( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U85 (.A1( u2_u2_u0_n101 ) , .ZN( u2_u2_u0_n130 ) , .A2( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U86 (.ZN( u2_u2_u0_n108 ) , .A1( u2_u2_u0_n92 ) , .A2( u2_u2_u0_n94 ) );
  NAND2_X1 u2_u2_u0_U87 (.ZN( u2_u2_u0_n142 ) , .A1( u2_u2_u0_n94 ) , .A2( u2_u2_u0_n95 ) );
  NAND3_X1 u2_u2_u0_U88 (.ZN( u2_out2_23 ) , .A3( u2_u2_u0_n137 ) , .A1( u2_u2_u0_n168 ) , .A2( u2_u2_u0_n171 ) );
  NAND3_X1 u2_u2_u0_U89 (.A3( u2_u2_u0_n127 ) , .A2( u2_u2_u0_n128 ) , .ZN( u2_u2_u0_n135 ) , .A1( u2_u2_u0_n150 ) );
  AND2_X1 u2_u2_u0_U9 (.A1( u2_u2_u0_n131 ) , .ZN( u2_u2_u0_n141 ) , .A2( u2_u2_u0_n150 ) );
  NAND3_X1 u2_u2_u0_U90 (.ZN( u2_u2_u0_n117 ) , .A3( u2_u2_u0_n132 ) , .A2( u2_u2_u0_n139 ) , .A1( u2_u2_u0_n148 ) );
  NAND3_X1 u2_u2_u0_U91 (.ZN( u2_u2_u0_n109 ) , .A2( u2_u2_u0_n114 ) , .A3( u2_u2_u0_n140 ) , .A1( u2_u2_u0_n149 ) );
  NAND3_X1 u2_u2_u0_U92 (.ZN( u2_out2_9 ) , .A3( u2_u2_u0_n106 ) , .A2( u2_u2_u0_n171 ) , .A1( u2_u2_u0_n174 ) );
  NAND3_X1 u2_u2_u0_U93 (.A2( u2_u2_u0_n128 ) , .A1( u2_u2_u0_n132 ) , .A3( u2_u2_u0_n146 ) , .ZN( u2_u2_u0_n97 ) );
  OAI22_X1 u2_u2_u2_U10 (.B1( u2_u2_u2_n151 ) , .A2( u2_u2_u2_n152 ) , .A1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n160 ) , .B2( u2_u2_u2_n168 ) );
  NAND3_X1 u2_u2_u2_U100 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n98 ) );
  NOR3_X1 u2_u2_u2_U11 (.A1( u2_u2_u2_n150 ) , .ZN( u2_u2_u2_n151 ) , .A3( u2_u2_u2_n175 ) , .A2( u2_u2_u2_n188 ) );
  AOI21_X1 u2_u2_u2_U12 (.B2( u2_u2_u2_n123 ) , .ZN( u2_u2_u2_n125 ) , .A( u2_u2_u2_n171 ) , .B1( u2_u2_u2_n184 ) );
  INV_X1 u2_u2_u2_U13 (.A( u2_u2_u2_n150 ) , .ZN( u2_u2_u2_n184 ) );
  AOI21_X1 u2_u2_u2_U14 (.ZN( u2_u2_u2_n144 ) , .B2( u2_u2_u2_n155 ) , .A( u2_u2_u2_n172 ) , .B1( u2_u2_u2_n185 ) );
  AOI21_X1 u2_u2_u2_U15 (.B2( u2_u2_u2_n143 ) , .ZN( u2_u2_u2_n145 ) , .B1( u2_u2_u2_n152 ) , .A( u2_u2_u2_n171 ) );
  INV_X1 u2_u2_u2_U16 (.A( u2_u2_u2_n156 ) , .ZN( u2_u2_u2_n171 ) );
  INV_X1 u2_u2_u2_U17 (.A( u2_u2_u2_n120 ) , .ZN( u2_u2_u2_n188 ) );
  NAND2_X1 u2_u2_u2_U18 (.A2( u2_u2_u2_n122 ) , .ZN( u2_u2_u2_n150 ) , .A1( u2_u2_u2_n152 ) );
  INV_X1 u2_u2_u2_U19 (.A( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n170 ) );
  INV_X1 u2_u2_u2_U20 (.A( u2_u2_u2_n137 ) , .ZN( u2_u2_u2_n173 ) );
  NAND2_X1 u2_u2_u2_U21 (.A1( u2_u2_u2_n132 ) , .A2( u2_u2_u2_n139 ) , .ZN( u2_u2_u2_n157 ) );
  INV_X1 u2_u2_u2_U22 (.A( u2_u2_u2_n113 ) , .ZN( u2_u2_u2_n178 ) );
  INV_X1 u2_u2_u2_U23 (.A( u2_u2_u2_n139 ) , .ZN( u2_u2_u2_n175 ) );
  INV_X1 u2_u2_u2_U24 (.A( u2_u2_u2_n155 ) , .ZN( u2_u2_u2_n181 ) );
  INV_X1 u2_u2_u2_U25 (.A( u2_u2_u2_n119 ) , .ZN( u2_u2_u2_n177 ) );
  INV_X1 u2_u2_u2_U26 (.A( u2_u2_u2_n116 ) , .ZN( u2_u2_u2_n180 ) );
  INV_X1 u2_u2_u2_U27 (.A( u2_u2_u2_n131 ) , .ZN( u2_u2_u2_n179 ) );
  INV_X1 u2_u2_u2_U28 (.A( u2_u2_u2_n154 ) , .ZN( u2_u2_u2_n176 ) );
  NAND2_X1 u2_u2_u2_U29 (.A2( u2_u2_u2_n116 ) , .A1( u2_u2_u2_n117 ) , .ZN( u2_u2_u2_n118 ) );
  NOR2_X1 u2_u2_u2_U3 (.ZN( u2_u2_u2_n121 ) , .A2( u2_u2_u2_n177 ) , .A1( u2_u2_u2_n180 ) );
  INV_X1 u2_u2_u2_U30 (.A( u2_u2_u2_n132 ) , .ZN( u2_u2_u2_n182 ) );
  INV_X1 u2_u2_u2_U31 (.A( u2_u2_u2_n158 ) , .ZN( u2_u2_u2_n183 ) );
  OAI21_X1 u2_u2_u2_U32 (.A( u2_u2_u2_n156 ) , .B1( u2_u2_u2_n157 ) , .ZN( u2_u2_u2_n158 ) , .B2( u2_u2_u2_n179 ) );
  NOR2_X1 u2_u2_u2_U33 (.ZN( u2_u2_u2_n156 ) , .A1( u2_u2_u2_n166 ) , .A2( u2_u2_u2_n169 ) );
  NOR2_X1 u2_u2_u2_U34 (.A2( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n137 ) , .A1( u2_u2_u2_n140 ) );
  NOR2_X1 u2_u2_u2_U35 (.A2( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n153 ) , .A1( u2_u2_u2_n156 ) );
  AOI211_X1 u2_u2_u2_U36 (.ZN( u2_u2_u2_n130 ) , .C1( u2_u2_u2_n138 ) , .C2( u2_u2_u2_n179 ) , .B( u2_u2_u2_n96 ) , .A( u2_u2_u2_n97 ) );
  OAI22_X1 u2_u2_u2_U37 (.B1( u2_u2_u2_n133 ) , .A2( u2_u2_u2_n137 ) , .A1( u2_u2_u2_n152 ) , .B2( u2_u2_u2_n168 ) , .ZN( u2_u2_u2_n97 ) );
  OAI221_X1 u2_u2_u2_U38 (.B1( u2_u2_u2_n113 ) , .C1( u2_u2_u2_n132 ) , .A( u2_u2_u2_n149 ) , .B2( u2_u2_u2_n171 ) , .C2( u2_u2_u2_n172 ) , .ZN( u2_u2_u2_n96 ) );
  OAI221_X1 u2_u2_u2_U39 (.A( u2_u2_u2_n115 ) , .C2( u2_u2_u2_n123 ) , .B2( u2_u2_u2_n143 ) , .B1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n163 ) , .C1( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U4 (.A( u2_u2_u2_n134 ) , .ZN( u2_u2_u2_n185 ) );
  OAI21_X1 u2_u2_u2_U40 (.A( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n115 ) , .B1( u2_u2_u2_n176 ) , .B2( u2_u2_u2_n178 ) );
  OAI221_X1 u2_u2_u2_U41 (.A( u2_u2_u2_n135 ) , .B2( u2_u2_u2_n136 ) , .B1( u2_u2_u2_n137 ) , .ZN( u2_u2_u2_n162 ) , .C2( u2_u2_u2_n167 ) , .C1( u2_u2_u2_n185 ) );
  AND3_X1 u2_u2_u2_U42 (.A3( u2_u2_u2_n131 ) , .A2( u2_u2_u2_n132 ) , .A1( u2_u2_u2_n133 ) , .ZN( u2_u2_u2_n136 ) );
  AOI22_X1 u2_u2_u2_U43 (.ZN( u2_u2_u2_n135 ) , .B1( u2_u2_u2_n140 ) , .A1( u2_u2_u2_n156 ) , .B2( u2_u2_u2_n180 ) , .A2( u2_u2_u2_n188 ) );
  AOI21_X1 u2_u2_u2_U44 (.ZN( u2_u2_u2_n149 ) , .B1( u2_u2_u2_n173 ) , .B2( u2_u2_u2_n188 ) , .A( u2_u2_u2_n95 ) );
  AND3_X1 u2_u2_u2_U45 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n156 ) , .ZN( u2_u2_u2_n95 ) );
  OAI21_X1 u2_u2_u2_U46 (.A( u2_u2_u2_n141 ) , .B2( u2_u2_u2_n142 ) , .ZN( u2_u2_u2_n146 ) , .B1( u2_u2_u2_n153 ) );
  OAI21_X1 u2_u2_u2_U47 (.A( u2_u2_u2_n140 ) , .ZN( u2_u2_u2_n141 ) , .B1( u2_u2_u2_n176 ) , .B2( u2_u2_u2_n177 ) );
  NOR3_X1 u2_u2_u2_U48 (.ZN( u2_u2_u2_n142 ) , .A3( u2_u2_u2_n175 ) , .A2( u2_u2_u2_n178 ) , .A1( u2_u2_u2_n181 ) );
  OAI21_X1 u2_u2_u2_U49 (.A( u2_u2_u2_n101 ) , .B2( u2_u2_u2_n121 ) , .B1( u2_u2_u2_n153 ) , .ZN( u2_u2_u2_n164 ) );
  NOR4_X1 u2_u2_u2_U5 (.A4( u2_u2_u2_n124 ) , .A3( u2_u2_u2_n125 ) , .A2( u2_u2_u2_n126 ) , .A1( u2_u2_u2_n127 ) , .ZN( u2_u2_u2_n128 ) );
  NAND2_X1 u2_u2_u2_U50 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n155 ) );
  NAND2_X1 u2_u2_u2_U51 (.A2( u2_u2_u2_n105 ) , .A1( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n143 ) );
  NAND2_X1 u2_u2_u2_U52 (.A1( u2_u2_u2_n104 ) , .A2( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n152 ) );
  NAND2_X1 u2_u2_u2_U53 (.A1( u2_u2_u2_n100 ) , .A2( u2_u2_u2_n105 ) , .ZN( u2_u2_u2_n132 ) );
  INV_X1 u2_u2_u2_U54 (.A( u2_u2_u2_n140 ) , .ZN( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U55 (.A( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n167 ) );
  INV_X1 u2_u2_u2_U56 (.ZN( u2_u2_u2_n187 ) , .A( u2_u2_u2_n99 ) );
  OAI21_X1 u2_u2_u2_U57 (.B1( u2_u2_u2_n137 ) , .B2( u2_u2_u2_n143 ) , .A( u2_u2_u2_n98 ) , .ZN( u2_u2_u2_n99 ) );
  NAND2_X1 u2_u2_u2_U58 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n113 ) );
  NAND2_X1 u2_u2_u2_U59 (.A1( u2_u2_u2_n106 ) , .A2( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n131 ) );
  AOI21_X1 u2_u2_u2_U6 (.B2( u2_u2_u2_n119 ) , .ZN( u2_u2_u2_n127 ) , .A( u2_u2_u2_n137 ) , .B1( u2_u2_u2_n155 ) );
  NAND2_X1 u2_u2_u2_U60 (.A1( u2_u2_u2_n103 ) , .A2( u2_u2_u2_n107 ) , .ZN( u2_u2_u2_n139 ) );
  NAND2_X1 u2_u2_u2_U61 (.A1( u2_u2_u2_n103 ) , .A2( u2_u2_u2_n105 ) , .ZN( u2_u2_u2_n133 ) );
  NAND2_X1 u2_u2_u2_U62 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n103 ) , .ZN( u2_u2_u2_n154 ) );
  NAND2_X1 u2_u2_u2_U63 (.A2( u2_u2_u2_n103 ) , .A1( u2_u2_u2_n104 ) , .ZN( u2_u2_u2_n119 ) );
  NAND2_X1 u2_u2_u2_U64 (.A2( u2_u2_u2_n107 ) , .A1( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n123 ) );
  NAND2_X1 u2_u2_u2_U65 (.A1( u2_u2_u2_n104 ) , .A2( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n122 ) );
  INV_X1 u2_u2_u2_U66 (.A( u2_u2_u2_n114 ) , .ZN( u2_u2_u2_n172 ) );
  NAND2_X1 u2_u2_u2_U67 (.A2( u2_u2_u2_n100 ) , .A1( u2_u2_u2_n102 ) , .ZN( u2_u2_u2_n116 ) );
  NAND2_X1 u2_u2_u2_U68 (.A1( u2_u2_u2_n102 ) , .A2( u2_u2_u2_n108 ) , .ZN( u2_u2_u2_n120 ) );
  NAND2_X1 u2_u2_u2_U69 (.A2( u2_u2_u2_n105 ) , .A1( u2_u2_u2_n106 ) , .ZN( u2_u2_u2_n117 ) );
  AOI21_X1 u2_u2_u2_U7 (.ZN( u2_u2_u2_n124 ) , .B1( u2_u2_u2_n131 ) , .B2( u2_u2_u2_n143 ) , .A( u2_u2_u2_n172 ) );
  NOR2_X1 u2_u2_u2_U70 (.A2( u2_u2_X_16 ) , .ZN( u2_u2_u2_n140 ) , .A1( u2_u2_u2_n166 ) );
  NOR2_X1 u2_u2_u2_U71 (.A2( u2_u2_X_13 ) , .A1( u2_u2_X_14 ) , .ZN( u2_u2_u2_n100 ) );
  NOR2_X1 u2_u2_u2_U72 (.A2( u2_u2_X_16 ) , .A1( u2_u2_X_17 ) , .ZN( u2_u2_u2_n138 ) );
  NOR2_X1 u2_u2_u2_U73 (.A2( u2_u2_X_15 ) , .A1( u2_u2_X_18 ) , .ZN( u2_u2_u2_n104 ) );
  NOR2_X1 u2_u2_u2_U74 (.A2( u2_u2_X_14 ) , .ZN( u2_u2_u2_n103 ) , .A1( u2_u2_u2_n174 ) );
  NOR2_X1 u2_u2_u2_U75 (.A2( u2_u2_X_15 ) , .ZN( u2_u2_u2_n102 ) , .A1( u2_u2_u2_n165 ) );
  NOR2_X1 u2_u2_u2_U76 (.A2( u2_u2_X_17 ) , .ZN( u2_u2_u2_n114 ) , .A1( u2_u2_u2_n169 ) );
  AND2_X1 u2_u2_u2_U77 (.A1( u2_u2_X_15 ) , .ZN( u2_u2_u2_n105 ) , .A2( u2_u2_u2_n165 ) );
  AND2_X1 u2_u2_u2_U78 (.A2( u2_u2_X_15 ) , .A1( u2_u2_X_18 ) , .ZN( u2_u2_u2_n107 ) );
  AND2_X1 u2_u2_u2_U79 (.A1( u2_u2_X_14 ) , .ZN( u2_u2_u2_n106 ) , .A2( u2_u2_u2_n174 ) );
  AOI21_X1 u2_u2_u2_U8 (.B2( u2_u2_u2_n120 ) , .B1( u2_u2_u2_n121 ) , .ZN( u2_u2_u2_n126 ) , .A( u2_u2_u2_n167 ) );
  AND2_X1 u2_u2_u2_U80 (.A1( u2_u2_X_13 ) , .A2( u2_u2_X_14 ) , .ZN( u2_u2_u2_n108 ) );
  INV_X1 u2_u2_u2_U81 (.A( u2_u2_X_16 ) , .ZN( u2_u2_u2_n169 ) );
  INV_X1 u2_u2_u2_U82 (.A( u2_u2_X_17 ) , .ZN( u2_u2_u2_n166 ) );
  INV_X1 u2_u2_u2_U83 (.A( u2_u2_X_13 ) , .ZN( u2_u2_u2_n174 ) );
  INV_X1 u2_u2_u2_U84 (.A( u2_u2_X_18 ) , .ZN( u2_u2_u2_n165 ) );
  NAND4_X1 u2_u2_u2_U85 (.ZN( u2_out2_24 ) , .A4( u2_u2_u2_n111 ) , .A3( u2_u2_u2_n112 ) , .A1( u2_u2_u2_n130 ) , .A2( u2_u2_u2_n187 ) );
  AOI21_X1 u2_u2_u2_U86 (.ZN( u2_u2_u2_n112 ) , .B2( u2_u2_u2_n156 ) , .A( u2_u2_u2_n164 ) , .B1( u2_u2_u2_n181 ) );
  AOI221_X1 u2_u2_u2_U87 (.A( u2_u2_u2_n109 ) , .B1( u2_u2_u2_n110 ) , .ZN( u2_u2_u2_n111 ) , .C1( u2_u2_u2_n134 ) , .C2( u2_u2_u2_n170 ) , .B2( u2_u2_u2_n173 ) );
  NAND4_X1 u2_u2_u2_U88 (.ZN( u2_out2_16 ) , .A4( u2_u2_u2_n128 ) , .A3( u2_u2_u2_n129 ) , .A1( u2_u2_u2_n130 ) , .A2( u2_u2_u2_n186 ) );
  AOI22_X1 u2_u2_u2_U89 (.A2( u2_u2_u2_n118 ) , .ZN( u2_u2_u2_n129 ) , .A1( u2_u2_u2_n140 ) , .B1( u2_u2_u2_n157 ) , .B2( u2_u2_u2_n170 ) );
  OAI22_X1 u2_u2_u2_U9 (.ZN( u2_u2_u2_n109 ) , .A2( u2_u2_u2_n113 ) , .B2( u2_u2_u2_n133 ) , .B1( u2_u2_u2_n167 ) , .A1( u2_u2_u2_n168 ) );
  INV_X1 u2_u2_u2_U90 (.A( u2_u2_u2_n163 ) , .ZN( u2_u2_u2_n186 ) );
  NAND4_X1 u2_u2_u2_U91 (.ZN( u2_out2_30 ) , .A4( u2_u2_u2_n147 ) , .A3( u2_u2_u2_n148 ) , .A2( u2_u2_u2_n149 ) , .A1( u2_u2_u2_n187 ) );
  NOR3_X1 u2_u2_u2_U92 (.A3( u2_u2_u2_n144 ) , .A2( u2_u2_u2_n145 ) , .A1( u2_u2_u2_n146 ) , .ZN( u2_u2_u2_n147 ) );
  AOI21_X1 u2_u2_u2_U93 (.B2( u2_u2_u2_n138 ) , .ZN( u2_u2_u2_n148 ) , .A( u2_u2_u2_n162 ) , .B1( u2_u2_u2_n182 ) );
  OR4_X1 u2_u2_u2_U94 (.ZN( u2_out2_6 ) , .A4( u2_u2_u2_n161 ) , .A3( u2_u2_u2_n162 ) , .A2( u2_u2_u2_n163 ) , .A1( u2_u2_u2_n164 ) );
  OR3_X1 u2_u2_u2_U95 (.A2( u2_u2_u2_n159 ) , .A1( u2_u2_u2_n160 ) , .ZN( u2_u2_u2_n161 ) , .A3( u2_u2_u2_n183 ) );
  AOI21_X1 u2_u2_u2_U96 (.B2( u2_u2_u2_n154 ) , .B1( u2_u2_u2_n155 ) , .ZN( u2_u2_u2_n159 ) , .A( u2_u2_u2_n167 ) );
  NAND3_X1 u2_u2_u2_U97 (.A2( u2_u2_u2_n117 ) , .A1( u2_u2_u2_n122 ) , .A3( u2_u2_u2_n123 ) , .ZN( u2_u2_u2_n134 ) );
  NAND3_X1 u2_u2_u2_U98 (.ZN( u2_u2_u2_n110 ) , .A2( u2_u2_u2_n131 ) , .A3( u2_u2_u2_n139 ) , .A1( u2_u2_u2_n154 ) );
  NAND3_X1 u2_u2_u2_U99 (.A2( u2_u2_u2_n100 ) , .ZN( u2_u2_u2_n101 ) , .A1( u2_u2_u2_n104 ) , .A3( u2_u2_u2_n114 ) );
  OAI21_X1 u2_uk_U173 (.ZN( u2_K16_30 ) , .B2( u2_uk_n1226 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n957 ) );
  NAND2_X1 u2_uk_U174 (.A1( u2_uk_K_r14_45 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n957 ) );
  OAI22_X1 u2_uk_U208 (.ZN( u2_K3_14 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1310 ) , .A2( u2_uk_n1317 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U283 (.ZN( u2_K3_6 ) , .A2( u2_uk_n1282 ) , .B2( u2_uk_n1287 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U342 (.ZN( u2_K3_4 ) , .B2( u2_uk_n1293 ) , .A2( u2_uk_n1301 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U368 (.ZN( u2_K16_28 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1189 ) , .A( u2_uk_n954 ) );
  OAI22_X1 u2_uk_U390 (.ZN( u2_K3_1 ) , .B2( u2_uk_n1285 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1290 ) , .B1( u2_uk_n27 ) );
  INV_X1 u2_uk_U481 (.ZN( u2_K16_29 ) , .A( u2_uk_n955 ) );
  OAI22_X1 u2_uk_U502 (.ZN( u2_K3_2 ) , .B2( u2_uk_n1301 ) , .A2( u2_uk_n1306 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U519 (.ZN( u2_K3_17 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1287 ) , .A2( u2_uk_n1310 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U682 (.ZN( u2_K3_3 ) , .A( u2_uk_n1013 ) , .B2( u2_uk_n1318 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U683 (.A1( u2_uk_K_r1_47 ) , .ZN( u2_uk_n1013 ) , .A2( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U709 (.ZN( u2_K16_25 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1209 ) , .A2( u2_uk_n1216 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U747 (.ZN( u2_K16_27 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1195 ) , .A2( u2_uk_n1200 ) , .A1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U845 (.ZN( u2_K3_18 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1295 ) , .A2( u2_uk_n1302 ) , .A1( u2_uk_n220 ) );
  OAI21_X1 u2_uk_U993 (.ZN( u2_K3_5 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1018 ) , .B2( u2_uk_n1302 ) );
endmodule

