module aes_aes_die_12 ( sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7 );
  input sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7;
  output sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7;
  wire us13_n438, us13_n439, us13_n440, us13_n441, us13_n442, us13_n443, us13_n444, us13_n445, us13_n446, 
       us13_n447, us13_n448, us13_n449, us13_n450, us13_n451, us13_n452, us13_n453, us13_n454, us13_n455, 
       us13_n456, us13_n457, us13_n458, us13_n459, us13_n460, us13_n461, us13_n462, us13_n463, us13_n464, 
       us13_n465, us13_n466, us13_n467, us13_n468, us13_n469, us13_n470, us13_n471, us13_n472, us13_n473, 
       us13_n474, us13_n475, us13_n476, us13_n477, us13_n478, us13_n479, us13_n480, us13_n481, us13_n482, 
       us13_n483, us13_n484, us13_n485, us13_n486, us13_n487, us13_n488, us13_n489, us13_n490, us13_n491, 
       us13_n492, us13_n493, us13_n494, us13_n495, us13_n496, us13_n497, us13_n498, us13_n499, us13_n500, 
       us13_n501, us13_n502, us13_n503, us13_n504, us13_n505, us13_n506, us13_n507, us13_n508, us13_n509, 
       us13_n510, us13_n511, us13_n512, us13_n513, us13_n514, us13_n515, us13_n516, us13_n517, us13_n518, 
       us13_n519, us13_n520, us13_n521, us13_n522, us13_n523, us13_n524, us13_n525, us13_n526, us13_n527, 
       us13_n528, us13_n529, us13_n530, us13_n531, us13_n532, us13_n533, us13_n534, us13_n535, us13_n536, 
       us13_n537, us13_n538, us13_n539, us13_n540, us13_n541, us13_n542, us13_n543, us13_n544, us13_n545, 
       us13_n546, us13_n547, us13_n548, us13_n549, us13_n550, us13_n551, us13_n552, us13_n553, us13_n554, 
       us13_n555, us13_n556, us13_n557, us13_n558, us13_n559, us13_n560, us13_n561, us13_n562, us13_n563, 
       us13_n564, us13_n565, us13_n566, us13_n567, us13_n568, us13_n569, us13_n570, us13_n571, us13_n572, 
       us13_n573, us13_n574, us13_n575, us13_n576, us13_n577, us13_n578, us13_n579, us13_n580, us13_n581, 
       us13_n582, us13_n583, us13_n584, us13_n585, us13_n586, us13_n587, us13_n588, us13_n589, us13_n590, 
       us13_n591, us13_n592, us13_n593, us13_n594, us13_n595, us13_n596, us13_n597, us13_n598, us13_n599, 
       us13_n600, us13_n601, us13_n602, us13_n603, us13_n604, us13_n605, us13_n606, us13_n607, us13_n608, 
       us13_n609, us13_n610, us13_n611, us13_n612, us13_n613, us13_n614, us13_n615, us13_n616, us13_n617, 
       us13_n618, us13_n619, us13_n620, us13_n621, us13_n622, us13_n623, us13_n624, us13_n625, us13_n626, 
       us13_n627, us13_n628, us13_n629, us13_n630, us13_n631, us13_n632, us13_n633, us13_n634, us13_n635, 
       us13_n636, us13_n637, us13_n638, us13_n639, us13_n640, us13_n641, us13_n642, us13_n643, us13_n644, 
       us13_n645, us13_n646, us13_n647, us13_n648, us13_n649, us13_n650, us13_n651, us13_n652, us13_n653, 
       us13_n654, us13_n655, us13_n656, us13_n657, us13_n658, us13_n659, us13_n660, us13_n661, us13_n662, 
       us13_n663, us13_n664, us13_n665, us13_n666, us13_n667, us13_n668, us13_n669, us13_n670, us13_n671, 
       us13_n672, us13_n673, us13_n674, us13_n675, us13_n676, us13_n677, us13_n678, us13_n679, us13_n680, 
       us13_n681, us13_n682, us13_n683, us13_n684, us13_n685, us13_n686, us13_n687, us13_n688, us13_n689, 
       us13_n690, us13_n691, us13_n692, us13_n693, us13_n694, us13_n695, us13_n696, us13_n697, us13_n698, 
       us13_n699, us13_n700, us13_n701, us13_n702, us13_n703, us13_n704, us13_n705, us13_n706, us13_n707, 
       us13_n708, us13_n709, us13_n710, us13_n711, us13_n712, us13_n713, us13_n714, us13_n715, us13_n716, 
       us13_n717, us13_n718, us13_n719, us13_n720, us13_n721, us13_n722, us13_n723, us13_n724, us13_n725, 
       us13_n726, us13_n727, us13_n728, us13_n729, us13_n730, us13_n731, us13_n732, us13_n733, us13_n734, 
       us13_n735, us13_n736, us13_n737, us13_n738, us13_n739, us13_n740, us13_n741, us13_n742, us13_n743, 
       us13_n744, us13_n745, us13_n746, us13_n747, us13_n748, us13_n749, us13_n750, us13_n751, us13_n752, 
       us13_n753, us13_n754, us13_n755, us13_n756, us13_n757, us13_n758, us13_n759, us13_n760, us13_n761, 
       us13_n762, us13_n763, us13_n764, us13_n765, us13_n766, us13_n767, us13_n768, us13_n769, us13_n770, 
       us13_n771, us13_n772, us13_n773, us13_n774, us13_n775, us13_n776, us13_n777, us13_n778, us13_n779, 
       us13_n780, us13_n781, us13_n782, us13_n783, us13_n784, us13_n785, us13_n786, us13_n787, us13_n788, 
       us13_n789, us13_n790, us13_n791, us13_n792, us13_n793, us13_n794, us13_n795, us13_n796, us13_n797, 
       us13_n798, us13_n799, us13_n800, us13_n801, us13_n802, us13_n803, us13_n804, us13_n805, us13_n806, 
       us13_n807, us13_n808, us13_n809, us13_n810, us13_n811, us13_n812, us13_n813, us13_n814, us13_n815, 
       us13_n816, us13_n817, us13_n818, us13_n819, us13_n820, us13_n821, us13_n822, us13_n823, us13_n824, 
       us13_n825, us13_n826, us13_n827, us13_n828, us13_n829, us13_n830, us13_n831, us13_n832, us13_n833, 
       us13_n834, us13_n835, us13_n836, us13_n837, us13_n838, us13_n839, us13_n840, us13_n841, us13_n842, 
       us13_n843, us13_n844, us13_n845, us13_n846, us13_n847, us13_n848, us13_n849, us13_n850, us13_n851, 
       us13_n852, us13_n853, us13_n854, us13_n855, us13_n856, us13_n857, us13_n858, us13_n859, us13_n860, 
       us13_n861, us13_n862, us13_n863, us13_n864, us13_n865, us13_n866, us13_n867, us13_n868, us13_n869, 
       us13_n870, us13_n871, us13_n872, us13_n873, us13_n874, us13_n875,  us13_n876;
  NOR3_X1 us13_U10 (.A3( us13_n621 ) , .A2( us13_n622 ) , .ZN( us13_n636 ) , .A1( us13_n725 ) );
  NOR4_X1 us13_U100 (.ZN( us13_n458 ) , .A2( us13_n509 ) , .A1( us13_n599 ) , .A4( us13_n628 ) , .A3( us13_n711 ) );
  NAND4_X1 us13_U101 (.A4( us13_n535 ) , .A3( us13_n536 ) , .A2( us13_n537 ) , .A1( us13_n538 ) , .ZN( us13_n622 ) );
  NOR4_X1 us13_U102 (.A4( us13_n526 ) , .A2( us13_n527 ) , .A1( us13_n528 ) , .ZN( us13_n538 ) , .A3( us13_n701 ) );
  NOR4_X1 us13_U103 (.A4( us13_n529 ) , .A3( us13_n530 ) , .ZN( us13_n537 ) , .A2( us13_n684 ) , .A1( us13_n794 ) );
  NOR4_X1 us13_U104 (.A4( us13_n532 ) , .A3( us13_n533 ) , .A2( us13_n534 ) , .ZN( us13_n535 ) , .A1( us13_n820 ) );
  NAND4_X1 us13_U105 (.A4( us13_n548 ) , .A3( us13_n549 ) , .A2( us13_n550 ) , .A1( us13_n551 ) , .ZN( us13_n745 ) );
  NOR3_X1 us13_U106 (.ZN( us13_n549 ) , .A2( us13_n651 ) , .A1( us13_n667 ) , .A3( us13_n771 ) );
  AOI211_X1 us13_U107 (.B( us13_n539 ) , .A( us13_n540 ) , .ZN( us13_n551 ) , .C2( us13_n839 ) , .C1( us13_n851 ) );
  NOR4_X1 us13_U108 (.A4( us13_n541 ) , .A3( us13_n542 ) , .A2( us13_n543 ) , .ZN( us13_n550 ) , .A1( us13_n688 ) );
  NAND4_X1 us13_U109 (.A4( us13_n479 ) , .A3( us13_n480 ) , .A2( us13_n481 ) , .A1( us13_n482 ) , .ZN( us13_n694 ) );
  NOR2_X1 us13_U11 (.A1( us13_n678 ) , .ZN( us13_n693 ) , .A2( us13_n807 ) );
  NOR3_X1 us13_U110 (.ZN( us13_n480 ) , .A2( us13_n508 ) , .A3( us13_n601 ) , .A1( us13_n610 ) );
  AOI211_X1 us13_U111 (.B( us13_n477 ) , .A( us13_n478 ) , .ZN( us13_n482 ) , .C2( us13_n833 ) , .C1( us13_n861 ) );
  NOR4_X1 us13_U112 (.ZN( us13_n481 ) , .A3( us13_n532 ) , .A4( us13_n545 ) , .A2( us13_n567 ) , .A1( us13_n717 ) );
  NOR2_X1 us13_U113 (.ZN( us13_n647 ) , .A1( us13_n854 ) , .A2( us13_n868 ) );
  NOR4_X1 us13_U114 (.ZN( us13_n620 ) , .A1( us13_n656 ) , .A3( us13_n666 ) , .A4( us13_n682 ) , .A2( us13_n766 ) );
  NOR4_X1 us13_U115 (.A4( us13_n609 ) , .A3( us13_n610 ) , .A2( us13_n611 ) , .A1( us13_n612 ) , .ZN( us13_n619 ) );
  NOR4_X1 us13_U116 (.A4( us13_n614 ) , .A3( us13_n615 ) , .A2( us13_n616 ) , .A1( us13_n617 ) , .ZN( us13_n618 ) );
  NOR2_X1 us13_U117 (.ZN( us13_n686 ) , .A1( us13_n831 ) , .A2( us13_n832 ) );
  NAND4_X1 us13_U118 (.A4( us13_n473 ) , .A3( us13_n474 ) , .A2( us13_n475 ) , .A1( us13_n476 ) , .ZN( us13_n678 ) );
  NOR4_X1 us13_U119 (.ZN( us13_n475 ) , .A1( us13_n531 ) , .A3( us13_n568 ) , .A4( us13_n600 ) , .A2( us13_n642 ) );
  INV_X1 us13_U12 (.A( us13_n607 ) , .ZN( us13_n874 ) );
  NOR4_X1 us13_U120 (.A4( us13_n470 ) , .ZN( us13_n476 ) , .A3( us13_n556 ) , .A1( us13_n735 ) , .A2( us13_n755 ) );
  NOR4_X1 us13_U121 (.ZN( us13_n474 ) , .A1( us13_n506 ) , .A3( us13_n544 ) , .A2( us13_n583 ) , .A4( us13_n716 ) );
  NOR2_X1 us13_U122 (.ZN( us13_n733 ) , .A2( us13_n832 ) , .A1( us13_n845 ) );
  NAND4_X1 us13_U123 (.A4( us13_n719 ) , .A3( us13_n720 ) , .A2( us13_n721 ) , .ZN( us13_n741 ) , .A1( us13_n857 ) );
  INV_X1 us13_U124 (.A( us13_n709 ) , .ZN( us13_n857 ) );
  NOR4_X1 us13_U125 (.A4( us13_n715 ) , .A3( us13_n716 ) , .A2( us13_n717 ) , .A1( us13_n718 ) , .ZN( us13_n719 ) );
  AOI221_X1 us13_U126 (.A( us13_n710 ) , .ZN( us13_n721 ) , .C2( us13_n844 ) , .B2( us13_n845 ) , .C1( us13_n861 ) , .B1( us13_n862 ) );
  NAND4_X1 us13_U127 (.A4( us13_n573 ) , .A3( us13_n574 ) , .A1( us13_n575 ) , .ZN( us13_n723 ) , .A2( us13_n874 ) );
  NOR4_X1 us13_U128 (.A4( us13_n569 ) , .A3( us13_n570 ) , .A2( us13_n571 ) , .A1( us13_n572 ) , .ZN( us13_n573 ) );
  AOI221_X1 us13_U129 (.A( us13_n564 ) , .C2( us13_n565 ) , .ZN( us13_n574 ) , .B2( us13_n845 ) , .B1( us13_n852 ) , .C1( us13_n853 ) );
  INV_X1 us13_U13 (.A( us13_n680 ) , .ZN( us13_n840 ) );
  NOR2_X1 us13_U130 (.ZN( us13_n575 ) , .A1( us13_n622 ) , .A2( us13_n745 ) );
  NAND4_X1 us13_U131 (.A4( us13_n633 ) , .A3( us13_n634 ) , .A2( us13_n635 ) , .A1( us13_n636 ) , .ZN( us13_n743 ) );
  AOI211_X1 us13_U132 (.B( us13_n623 ) , .A( us13_n624 ) , .ZN( us13_n635 ) , .C2( us13_n836 ) , .C1( us13_n863 ) );
  NOR4_X1 us13_U133 (.A4( us13_n629 ) , .A3( us13_n630 ) , .A2( us13_n631 ) , .A1( us13_n632 ) , .ZN( us13_n633 ) );
  NOR4_X1 us13_U134 (.A4( us13_n626 ) , .A3( us13_n627 ) , .A2( us13_n628 ) , .ZN( us13_n634 ) , .A1( us13_n664 ) );
  NAND4_X1 us13_U135 (.A4( us13_n493 ) , .A3( us13_n494 ) , .A1( us13_n495 ) , .ZN( us13_n802 ) , .A2( us13_n867 ) );
  AOI221_X1 us13_U136 (.A( us13_n489 ) , .ZN( us13_n494 ) , .B2( us13_n836 ) , .C2( us13_n841 ) , .C1( us13_n851 ) , .B1( us13_n860 ) );
  INV_X1 us13_U137 (.A( us13_n778 ) , .ZN( us13_n867 ) );
  NOR2_X1 us13_U138 (.ZN( us13_n495 ) , .A1( us13_n678 ) , .A2( us13_n694 ) );
  INV_X1 us13_U139 (.A( us13_n762 ) , .ZN( us13_n830 ) );
  NOR4_X1 us13_U14 (.A4( us13_n445 ) , .A3( us13_n446 ) , .A2( us13_n516 ) , .A1( us13_n541 ) , .ZN( us13_n706 ) );
  OR4_X1 us13_U140 (.A4( us13_n566 ) , .A3( us13_n567 ) , .A2( us13_n568 ) , .ZN( us13_n572 ) , .A1( us13_n665 ) );
  OR4_X1 us13_U141 (.A4( us13_n518 ) , .A2( us13_n519 ) , .A1( us13_n520 ) , .ZN( us13_n522 ) , .A3( us13_n821 ) );
  OR4_X1 us13_U142 (.ZN( us13_n466 ) , .A4( us13_n518 ) , .A3( us13_n529 ) , .A2( us13_n578 ) , .A1( us13_n712 ) );
  OR4_X1 us13_U143 (.A4( us13_n682 ) , .A3( us13_n683 ) , .A2( us13_n684 ) , .A1( us13_n685 ) , .ZN( us13_n690 ) );
  OR4_X1 us13_U144 (.A4( us13_n580 ) , .A3( us13_n581 ) , .A2( us13_n582 ) , .A1( us13_n583 ) , .ZN( us13_n584 ) );
  NAND2_X1 us13_U145 (.ZN( us13_n613 ) , .A2( us13_n837 ) , .A1( us13_n873 ) );
  OR3_X1 us13_U146 (.A3( us13_n506 ) , .A2( us13_n507 ) , .A1( us13_n508 ) , .ZN( us13_n511 ) );
  AOI221_X1 us13_U147 (.A( us13_n713 ) , .B2( us13_n714 ) , .ZN( us13_n720 ) , .C1( us13_n832 ) , .B1( us13_n839 ) , .C2( us13_n863 ) );
  OR2_X1 us13_U148 (.A2( us13_n711 ) , .A1( us13_n712 ) , .ZN( us13_n713 ) );
  INV_X1 us13_U149 (.A( us13_n463 ) , .ZN( us13_n864 ) );
  OR3_X1 us13_U15 (.ZN( us13_n446 ) , .A1( us13_n528 ) , .A3( us13_n577 ) , .A2( us13_n875 ) );
  OAI21_X1 us13_U150 (.ZN( us13_n463 ) , .B1( us13_n809 ) , .A( us13_n834 ) , .B2( us13_n851 ) );
  INV_X1 us13_U151 (.A( us13_n754 ) , .ZN( us13_n869 ) );
  OAI21_X1 us13_U152 (.B1( us13_n753 ) , .ZN( us13_n754 ) , .A( us13_n845 ) , .B2( us13_n868 ) );
  INV_X1 us13_U153 (.A( us13_n672 ) , .ZN( us13_n859 ) );
  AOI21_X1 us13_U154 (.A( us13_n670 ) , .B1( us13_n671 ) , .ZN( us13_n672 ) , .B2( us13_n856 ) );
  NAND2_X1 us13_U155 (.A1( us13_n447 ) , .A2( us13_n465 ) , .ZN( us13_n749 ) );
  OAI222_X1 us13_U156 (.B2( us13_n747 ) , .B1( us13_n748 ) , .A2( us13_n749 ) , .ZN( us13_n757 ) , .C2( us13_n805 ) , .C1( us13_n814 ) , .A1( us13_n817 ) );
  OAI222_X1 us13_U157 (.B2( us13_n708 ) , .ZN( us13_n709 ) , .C2( us13_n724 ) , .B1( us13_n747 ) , .A1( us13_n806 ) , .C1( us13_n814 ) , .A2( us13_n815 ) );
  OAI222_X1 us13_U158 (.ZN( us13_n505 ) , .C2( us13_n625 ) , .B2( us13_n647 ) , .B1( us13_n747 ) , .A2( us13_n748 ) , .C1( us13_n805 ) , .A1( us13_n806 ) );
  NOR4_X1 us13_U159 (.A2( us13_n491 ) , .A1( us13_n492 ) , .ZN( us13_n493 ) , .A3( us13_n580 ) , .A4( us13_n612 ) );
  OR4_X1 us13_U16 (.A4( us13_n442 ) , .A2( us13_n443 ) , .A1( us13_n444 ) , .ZN( us13_n445 ) , .A3( us13_n553 ) );
  OR4_X1 us13_U160 (.ZN( us13_n492 ) , .A4( us13_n534 ) , .A2( us13_n547 ) , .A1( us13_n559 ) , .A3( us13_n632 ) );
  OAI22_X1 us13_U161 (.B1( us13_n490 ) , .ZN( us13_n491 ) , .A1( us13_n686 ) , .A2( us13_n763 ) , .B2( us13_n817 ) );
  NOR3_X1 us13_U162 (.ZN( us13_n490 ) , .A1( us13_n782 ) , .A2( us13_n850 ) , .A3( us13_n863 ) );
  INV_X1 us13_U163 (.A( us13_n730 ) , .ZN( us13_n839 ) );
  INV_X1 us13_U164 (.A( us13_n790 ) , .ZN( us13_n832 ) );
  NAND2_X1 us13_U165 (.A1( us13_n451 ) , .A2( us13_n453 ) , .ZN( us13_n762 ) );
  AOI211_X1 us13_U166 (.A( us13_n637 ) , .ZN( us13_n645 ) , .B( us13_n743 ) , .C2( us13_n839 ) , .C1( us13_n854 ) );
  OAI22_X1 us13_U167 (.ZN( us13_n637 ) , .A1( us13_n699 ) , .B2( us13_n728 ) , .A2( us13_n762 ) , .B1( us13_n816 ) );
  OAI221_X1 us13_U168 (.A( us13_n727 ) , .C2( us13_n728 ) , .B2( us13_n729 ) , .B1( us13_n730 ) , .ZN( us13_n737 ) , .C1( us13_n817 ) );
  AOI22_X1 us13_U169 (.ZN( us13_n727 ) , .B1( us13_n832 ) , .A2( us13_n838 ) , .A1( us13_n863 ) , .B2( us13_n866 ) );
  INV_X1 us13_U17 (.A( us13_n613 ) , .ZN( us13_n875 ) );
  INV_X1 us13_U170 (.A( us13_n744 ) , .ZN( us13_n837 ) );
  OAI22_X1 us13_U171 (.ZN( us13_n489 ) , .A1( us13_n724 ) , .B2( us13_n728 ) , .B1( us13_n730 ) , .A2( us13_n779 ) );
  OAI22_X1 us13_U172 (.ZN( us13_n624 ) , .B1( us13_n669 ) , .B2( us13_n747 ) , .A1( us13_n815 ) , .A2( us13_n816 ) );
  OAI22_X1 us13_U173 (.B2( us13_n779 ) , .B1( us13_n780 ) , .ZN( us13_n781 ) , .A2( us13_n814 ) , .A1( us13_n815 ) );
  OAI22_X1 us13_U174 (.A1( us13_n724 ) , .ZN( us13_n726 ) , .B2( us13_n750 ) , .B1( us13_n812 ) , .A2( us13_n816 ) );
  INV_X1 us13_U175 (.A( us13_n805 ) , .ZN( us13_n860 ) );
  OAI22_X1 us13_U176 (.B2( us13_n744 ) , .ZN( us13_n746 ) , .A2( us13_n762 ) , .B1( us13_n780 ) , .A1( us13_n792 ) );
  OAI22_X1 us13_U177 (.B2( us13_n803 ) , .B1( us13_n804 ) , .A2( us13_n805 ) , .A1( us13_n806 ) , .ZN( us13_n808 ) );
  OAI22_X1 us13_U178 (.ZN( us13_n496 ) , .A2( us13_n744 ) , .A1( us13_n780 ) , .B1( us13_n791 ) , .B2( us13_n806 ) );
  OAI22_X1 us13_U179 (.ZN( us13_n710 ) , .A2( us13_n728 ) , .B2( us13_n729 ) , .A1( us13_n744 ) , .B1( us13_n813 ) );
  INV_X1 us13_U18 (.A( us13_n749 ) , .ZN( us13_n863 ) );
  INV_X1 us13_U180 (.A( us13_n788 ) , .ZN( us13_n845 ) );
  INV_X1 us13_U181 (.A( us13_n814 ) , .ZN( us13_n833 ) );
  OAI22_X1 us13_U182 (.ZN( us13_n590 ) , .B1( us13_n730 ) , .B2( us13_n749 ) , .A2( us13_n786 ) , .A1( us13_n803 ) );
  OAI22_X1 us13_U183 (.ZN( us13_n695 ) , .A2( us13_n730 ) , .A1( us13_n780 ) , .B1( us13_n791 ) , .B2( us13_n817 ) );
  INV_X1 us13_U184 (.A( us13_n816 ) , .ZN( us13_n831 ) );
  INV_X1 us13_U185 (.A( us13_n669 ) , .ZN( us13_n865 ) );
  NOR2_X1 us13_U186 (.ZN( us13_n715 ) , .A1( us13_n805 ) , .A2( us13_n817 ) );
  NOR2_X1 us13_U187 (.ZN( us13_n718 ) , .A2( us13_n724 ) , .A1( us13_n744 ) );
  NOR2_X1 us13_U188 (.ZN( us13_n666 ) , .A1( us13_n728 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U189 (.ZN( us13_n546 ) , .A2( us13_n780 ) , .A1( us13_n814 ) );
  AOI222_X1 us13_U19 (.ZN( us13_n563 ) , .B1( us13_n830 ) , .C1( us13_n841 ) , .A2( us13_n843 ) , .A1( us13_n854 ) , .B2( us13_n863 ) , .C2( us13_n873 ) );
  NOR2_X1 us13_U190 (.ZN( us13_n577 ) , .A2( us13_n699 ) , .A1( us13_n814 ) );
  NOR2_X1 us13_U191 (.ZN( us13_n570 ) , .A1( us13_n728 ) , .A2( us13_n806 ) );
  NOR2_X1 us13_U192 (.A2( us13_n744 ) , .ZN( us13_n755 ) , .A1( us13_n805 ) );
  INV_X1 us13_U193 (.A( us13_n750 ) , .ZN( us13_n842 ) );
  NOR2_X1 us13_U194 (.ZN( us13_n735 ) , .A2( us13_n803 ) , .A1( us13_n805 ) );
  NOR2_X1 us13_U195 (.ZN( us13_n532 ) , .A2( us13_n749 ) , .A1( us13_n750 ) );
  NOR2_X1 us13_U196 (.ZN( us13_n654 ) , .A1( us13_n728 ) , .A2( us13_n813 ) );
  OAI22_X1 us13_U197 (.ZN( us13_n483 ) , .A1( us13_n708 ) , .B2( us13_n785 ) , .A2( us13_n806 ) , .B1( us13_n812 ) );
  NOR2_X1 us13_U198 (.ZN( us13_n629 ) , .A2( us13_n728 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U199 (.ZN( us13_n615 ) , .A1( us13_n785 ) , .A2( us13_n815 ) );
  AOI222_X1 us13_U20 (.ZN( us13_n660 ) , .A2( us13_n839 ) , .B1( us13_n841 ) , .C2( us13_n845 ) , .A1( us13_n860 ) , .C1( us13_n863 ) , .B2( us13_n870 ) );
  NOR2_X1 us13_U200 (.ZN( us13_n612 ) , .A1( us13_n779 ) , .A2( us13_n786 ) );
  NOR2_X1 us13_U201 (.ZN( us13_n628 ) , .A2( us13_n669 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U202 (.ZN( us13_n611 ) , .A2( us13_n780 ) , .A1( us13_n806 ) );
  NOR2_X1 us13_U203 (.ZN( us13_n601 ) , .A2( us13_n780 ) , .A1( us13_n803 ) );
  INV_X1 us13_U204 (.A( us13_n747 ) , .ZN( us13_n834 ) );
  NOR2_X1 us13_U205 (.ZN( us13_n528 ) , .A2( us13_n724 ) , .A1( us13_n803 ) );
  NOR2_X1 us13_U206 (.ZN( us13_n531 ) , .A2( us13_n780 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U207 (.A2( us13_n708 ) , .A1( us13_n750 ) , .ZN( us13_n771 ) );
  NOR2_X1 us13_U208 (.ZN( us13_n599 ) , .A2( us13_n791 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U209 (.ZN( us13_n652 ) , .A1( us13_n669 ) , .A2( us13_n814 ) );
  INV_X1 us13_U21 (.A( us13_n647 ) , .ZN( us13_n870 ) );
  INV_X1 us13_U210 (.A( us13_n792 ) , .ZN( us13_n851 ) );
  NOR2_X1 us13_U211 (.A1( us13_n669 ) , .ZN( us13_n673 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U212 (.ZN( us13_n602 ) , .A1( us13_n669 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U213 (.A1( us13_n669 ) , .ZN( us13_n688 ) , .A2( us13_n816 ) );
  NOR2_X1 us13_U214 (.ZN( us13_n667 ) , .A1( us13_n750 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U215 (.A2( us13_n744 ) , .ZN( us13_n769 ) , .A1( us13_n812 ) );
  NOR2_X1 us13_U216 (.ZN( us13_n555 ) , .A1( us13_n750 ) , .A2( us13_n791 ) );
  NOR2_X1 us13_U217 (.ZN( us13_n508 ) , .A2( us13_n780 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U218 (.ZN( us13_n543 ) , .A2( us13_n708 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U219 (.ZN( us13_n664 ) , .A1( us13_n785 ) , .A2( us13_n791 ) );
  NOR4_X1 us13_U22 (.ZN( us13_n473 ) , .A2( us13_n521 ) , .A4( us13_n594 ) , .A1( us13_n609 ) , .A3( us13_n629 ) );
  NOR2_X1 us13_U220 (.A1( us13_n669 ) , .ZN( us13_n766 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U221 (.A1( us13_n699 ) , .ZN( us13_n768 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U222 (.ZN( us13_n527 ) , .A1( us13_n669 ) , .A2( us13_n779 ) );
  NOR2_X1 us13_U223 (.ZN( us13_n557 ) , .A1( us13_n792 ) , .A2( us13_n814 ) );
  NOR2_X1 us13_U224 (.ZN( us13_n545 ) , .A1( us13_n749 ) , .A2( us13_n814 ) );
  NOR2_X1 us13_U225 (.ZN( us13_n556 ) , .A1( us13_n762 ) , .A2( us13_n805 ) );
  NOR2_X1 us13_U226 (.ZN( us13_n661 ) , .A1( us13_n729 ) , .A2( us13_n790 ) );
  NOR2_X1 us13_U227 (.ZN( us13_n507 ) , .A1( us13_n812 ) , .A2( us13_n817 ) );
  INV_X1 us13_U228 (.A( us13_n806 ) , .ZN( us13_n841 ) );
  NOR2_X1 us13_U229 (.ZN( us13_n554 ) , .A1( us13_n786 ) , .A2( us13_n813 ) );
  NOR4_X1 us13_U23 (.A4( us13_n544 ) , .A3( us13_n545 ) , .A2( us13_n546 ) , .A1( us13_n547 ) , .ZN( us13_n548 ) );
  NOR2_X1 us13_U230 (.ZN( us13_n509 ) , .A1( us13_n729 ) , .A2( us13_n779 ) );
  NOR2_X1 us13_U231 (.ZN( us13_n530 ) , .A2( us13_n744 ) , .A1( us13_n792 ) );
  OAI22_X1 us13_U232 (.B2( us13_n750 ) , .B1( us13_n751 ) , .A1( us13_n752 ) , .ZN( us13_n756 ) , .A2( us13_n806 ) );
  NOR2_X1 us13_U233 (.ZN( us13_n751 ) , .A2( us13_n852 ) , .A1( us13_n860 ) );
  NOR3_X1 us13_U234 (.ZN( us13_n752 ) , .A2( us13_n853 ) , .A1( us13_n863 ) , .A3( us13_n865 ) );
  NOR2_X1 us13_U235 (.ZN( us13_n544 ) , .A2( us13_n785 ) , .A1( us13_n792 ) );
  NOR2_X1 us13_U236 (.A1( us13_n749 ) , .ZN( us13_n767 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U237 (.ZN( us13_n516 ) , .A1( us13_n708 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U238 (.ZN( us13_n663 ) , .A1( us13_n729 ) , .A2( us13_n785 ) );
  OAI22_X1 us13_U239 (.B1( us13_n440 ) , .ZN( us13_n444 ) , .A2( us13_n728 ) , .A1( us13_n744 ) , .B2( us13_n749 ) );
  NOR4_X1 us13_U24 (.ZN( us13_n479 ) , .A1( us13_n520 ) , .A4( us13_n557 ) , .A3( us13_n582 ) , .A2( us13_n630 ) );
  NOR3_X1 us13_U240 (.ZN( us13_n440 ) , .A2( us13_n836 ) , .A3( us13_n837 ) , .A1( us13_n846 ) );
  NOR2_X1 us13_U241 (.ZN( us13_n717 ) , .A2( us13_n744 ) , .A1( us13_n786 ) );
  INV_X1 us13_U242 (.A( us13_n728 ) , .ZN( us13_n852 ) );
  NOR2_X1 us13_U243 (.ZN( us13_n506 ) , .A2( us13_n728 ) , .A1( us13_n762 ) );
  NOR2_X1 us13_U244 (.ZN( us13_n614 ) , .A1( us13_n762 ) , .A2( us13_n812 ) );
  NOR2_X1 us13_U245 (.ZN( us13_n517 ) , .A1( us13_n708 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U246 (.ZN( us13_n558 ) , .A1( us13_n708 ) , .A2( us13_n816 ) );
  AOI21_X1 us13_U247 (.A( us13_n812 ) , .B2( us13_n813 ) , .B1( us13_n814 ) , .ZN( us13_n819 ) );
  NOR2_X1 us13_U248 (.ZN( us13_n670 ) , .A1( us13_n790 ) , .A2( us13_n805 ) );
  NOR2_X1 us13_U249 (.ZN( us13_n630 ) , .A1( us13_n747 ) , .A2( us13_n815 ) );
  NOR4_X1 us13_U25 (.ZN( us13_n456 ) , .A2( us13_n517 ) , .A1( us13_n543 ) , .A3( us13_n579 ) , .A4( us13_n615 ) );
  NOR2_X1 us13_U250 (.ZN( us13_n655 ) , .A1( us13_n790 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U251 (.ZN( us13_n521 ) , .A1( us13_n790 ) , .A2( us13_n812 ) );
  NOR2_X1 us13_U252 (.ZN( us13_n668 ) , .A2( us13_n708 ) , .A1( us13_n790 ) );
  NOR2_X1 us13_U253 (.ZN( us13_n542 ) , .A1( us13_n762 ) , .A2( us13_n791 ) );
  NOR2_X1 us13_U254 (.ZN( us13_n701 ) , .A2( us13_n786 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U255 (.ZN( us13_n631 ) , .A1( us13_n724 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U256 (.ZN( us13_n656 ) , .A1( us13_n747 ) , .A2( us13_n780 ) );
  INV_X1 us13_U257 (.A( us13_n763 ) , .ZN( us13_n866 ) );
  NOR2_X1 us13_U258 (.ZN( us13_n609 ) , .A2( us13_n724 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U259 (.A1( us13_n730 ) , .ZN( us13_n765 ) , .A2( us13_n786 ) );
  NOR4_X1 us13_U26 (.ZN( us13_n485 ) , .A2( us13_n533 ) , .A1( us13_n558 ) , .A3( us13_n631 ) , .A4( us13_n718 ) );
  NOR2_X1 us13_U260 (.ZN( us13_n533 ) , .A2( us13_n724 ) , .A1( us13_n730 ) );
  NOR2_X1 us13_U261 (.ZN( us13_n579 ) , .A2( us13_n708 ) , .A1( us13_n730 ) );
  AOI21_X1 us13_U262 (.B1( us13_n625 ) , .ZN( us13_n627 ) , .A( us13_n763 ) , .B2( us13_n814 ) );
  AOI21_X1 us13_U263 (.A( us13_n815 ) , .B2( us13_n816 ) , .B1( us13_n817 ) , .ZN( us13_n818 ) );
  NOR2_X1 us13_U264 (.ZN( us13_n582 ) , .A1( us13_n744 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U265 (.A2( us13_n708 ) , .A1( us13_n762 ) , .ZN( us13_n794 ) );
  AOI21_X1 us13_U266 (.ZN( us13_n515 ) , .A( us13_n729 ) , .B1( us13_n750 ) , .B2( us13_n803 ) );
  NOR2_X1 us13_U267 (.ZN( us13_n642 ) , .A2( us13_n788 ) , .A1( us13_n791 ) );
  AOI21_X1 us13_U268 (.ZN( us13_n499 ) , .B1( us13_n680 ) , .A( us13_n812 ) , .B2( us13_n816 ) );
  AOI21_X1 us13_U269 (.ZN( us13_n650 ) , .A( us13_n779 ) , .B1( us13_n792 ) , .B2( us13_n805 ) );
  NOR4_X1 us13_U27 (.A1( us13_n531 ) , .ZN( us13_n536 ) , .A2( us13_n654 ) , .A4( us13_n668 ) , .A3( us13_n765 ) );
  NOR2_X1 us13_U270 (.ZN( us13_n520 ) , .A2( us13_n708 ) , .A1( us13_n814 ) );
  AOI21_X1 us13_U271 (.ZN( us13_n626 ) , .B2( us13_n669 ) , .A( us13_n790 ) , .B1( us13_n791 ) );
  NOR2_X1 us13_U272 (.ZN( us13_n653 ) , .A1( us13_n762 ) , .A2( us13_n786 ) );
  AOI21_X1 us13_U273 (.ZN( us13_n477 ) , .A( us13_n669 ) , .B1( us13_n750 ) , .B2( us13_n806 ) );
  NOR2_X1 us13_U274 (.ZN( us13_n559 ) , .A2( us13_n791 ) , .A1( us13_n803 ) );
  NOR2_X1 us13_U275 (.ZN( us13_n519 ) , .A2( us13_n699 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U276 (.ZN( us13_n683 ) , .A2( us13_n699 ) , .A1( us13_n803 ) );
  AOI21_X1 us13_U277 (.ZN( us13_n510 ) , .B2( us13_n669 ) , .A( us13_n730 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U278 (.ZN( us13_n540 ) , .A( us13_n763 ) , .B2( us13_n779 ) , .B1( us13_n817 ) );
  NOR2_X1 us13_U279 (.ZN( us13_n581 ) , .A1( us13_n669 ) , .A2( us13_n788 ) );
  NOR2_X1 us13_U28 (.ZN( us13_n680 ) , .A2( us13_n834 ) , .A1( us13_n839 ) );
  AOI21_X1 us13_U280 (.ZN( us13_n589 ) , .B2( us13_n699 ) , .B1( us13_n815 ) , .A( us13_n817 ) );
  AOI21_X1 us13_U281 (.ZN( us13_n498 ) , .A( us13_n724 ) , .B2( us13_n762 ) , .B1( us13_n814 ) );
  AOI21_X1 us13_U282 (.ZN( us13_n539 ) , .B2( us13_n812 ) , .A( us13_n814 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U283 (.B1( us13_n699 ) , .ZN( us13_n700 ) , .A( us13_n732 ) , .B2( us13_n763 ) );
  AOI21_X1 us13_U284 (.ZN( us13_n591 ) , .B2( us13_n763 ) , .A( us13_n785 ) , .B1( us13_n812 ) );
  INV_X1 us13_U285 (.A( us13_n791 ) , .ZN( us13_n873 ) );
  NOR2_X1 us13_U286 (.ZN( us13_n547 ) , .A1( us13_n699 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U287 (.ZN( us13_n665 ) , .A1( us13_n780 ) , .A2( us13_n813 ) );
  INV_X1 us13_U288 (.A( us13_n729 ) , .ZN( us13_n868 ) );
  AOI21_X1 us13_U289 (.ZN( us13_n640 ) , .B2( us13_n747 ) , .A( us13_n792 ) , .B1( us13_n803 ) );
  AOI221_X1 us13_U29 (.A( us13_n781 ) , .ZN( us13_n798 ) , .C2( us13_n837 ) , .B2( us13_n838 ) , .B1( us13_n865 ) , .C1( us13_n866 ) );
  AOI21_X1 us13_U290 (.ZN( us13_n569 ) , .B1( us13_n750 ) , .B2( us13_n762 ) , .A( us13_n780 ) );
  AOI21_X1 us13_U291 (.ZN( us13_n649 ) , .B1( us13_n729 ) , .B2( us13_n763 ) , .A( us13_n813 ) );
  NOR2_X1 us13_U292 (.ZN( us13_n685 ) , .A1( us13_n729 ) , .A2( us13_n816 ) );
  AOI21_X1 us13_U293 (.B1( us13_n686 ) , .ZN( us13_n687 ) , .A( us13_n728 ) , .B2( us13_n761 ) );
  NOR2_X1 us13_U294 (.ZN( us13_n568 ) , .A1( us13_n729 ) , .A2( us13_n762 ) );
  NOR2_X1 us13_U295 (.ZN( us13_n684 ) , .A1( us13_n791 ) , .A2( us13_n813 ) );
  AOI21_X1 us13_U296 (.ZN( us13_n514 ) , .A( us13_n779 ) , .B2( us13_n792 ) , .B1( us13_n812 ) );
  AOI21_X1 us13_U297 (.ZN( us13_n593 ) , .B1( us13_n750 ) , .A( us13_n792 ) , .B2( us13_n813 ) );
  AOI21_X1 us13_U298 (.ZN( us13_n450 ) , .B2( us13_n792 ) , .A( us13_n803 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U299 (.ZN( us13_n639 ) , .B2( us13_n749 ) , .A( us13_n788 ) , .B1( us13_n812 ) );
  NAND4_X1 us13_U3 (.ZN( sa12_sr_2 ) , .A4( us13_n643 ) , .A3( us13_n644 ) , .A2( us13_n645 ) , .A1( us13_n646 ) );
  NOR4_X1 us13_U30 (.A4( us13_n793 ) , .A3( us13_n794 ) , .A2( us13_n795 ) , .A1( us13_n796 ) , .ZN( us13_n797 ) );
  INV_X1 us13_U300 (.A( us13_n699 ) , .ZN( us13_n853 ) );
  AOI21_X1 us13_U301 (.ZN( us13_n564 ) , .B1( us13_n724 ) , .A( us13_n779 ) , .B2( us13_n791 ) );
  AOI21_X1 us13_U302 (.ZN( us13_n497 ) , .A( us13_n779 ) , .B2( us13_n791 ) , .B1( us13_n804 ) );
  NOR2_X1 us13_U303 (.ZN( us13_n529 ) , .A1( us13_n708 ) , .A2( us13_n779 ) );
  AOI21_X1 us13_U304 (.ZN( us13_n689 ) , .B2( us13_n749 ) , .B1( us13_n763 ) , .A( us13_n806 ) );
  NOR2_X1 us13_U305 (.ZN( us13_n567 ) , .A1( us13_n747 ) , .A2( us13_n805 ) );
  AOI21_X1 us13_U306 (.A( us13_n790 ) , .B2( us13_n791 ) , .B1( us13_n792 ) , .ZN( us13_n793 ) );
  AOI21_X1 us13_U307 (.A( us13_n733 ) , .ZN( us13_n734 ) , .B2( us13_n780 ) , .B1( us13_n792 ) );
  NOR2_X1 us13_U308 (.A2( us13_n813 ) , .A1( us13_n815 ) , .ZN( us13_n821 ) );
  AOI21_X1 us13_U309 (.ZN( us13_n641 ) , .B1( us13_n680 ) , .A( us13_n791 ) , .B2( us13_n817 ) );
  NOR4_X1 us13_U31 (.A4( us13_n776 ) , .A3( us13_n777 ) , .A1( us13_n778 ) , .ZN( us13_n799 ) , .A2( us13_n801 ) );
  NOR2_X1 us13_U310 (.ZN( us13_n578 ) , .A1( us13_n708 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U311 (.ZN( us13_n682 ) , .A2( us13_n708 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U312 (.ZN( us13_n711 ) , .A1( us13_n762 ) , .A2( us13_n763 ) );
  NOR2_X1 us13_U313 (.ZN( us13_n583 ) , .A1( us13_n792 ) , .A2( us13_n817 ) );
  NOR2_X1 us13_U314 (.ZN( us13_n534 ) , .A1( us13_n724 ) , .A2( us13_n788 ) );
  NAND2_X1 us13_U315 (.ZN( us13_n753 ) , .A1( us13_n763 ) , .A2( us13_n805 ) );
  INV_X1 us13_U316 (.A( us13_n815 ) , .ZN( us13_n855 ) );
  AOI21_X1 us13_U317 (.ZN( us13_n442 ) , .A( us13_n699 ) , .B1( us13_n733 ) , .B2( us13_n750 ) );
  OAI21_X1 us13_U318 (.A( us13_n731 ) , .B1( us13_n732 ) , .ZN( us13_n736 ) , .B2( us13_n805 ) );
  OAI21_X1 us13_U319 (.ZN( us13_n731 ) , .A( us13_n833 ) , .B2( us13_n852 ) , .B1( us13_n873 ) );
  NOR4_X1 us13_U32 (.A3( us13_n755 ) , .A2( us13_n756 ) , .A1( us13_n757 ) , .ZN( us13_n758 ) , .A4( us13_n869 ) );
  INV_X1 us13_U320 (.A( us13_n780 ) , .ZN( us13_n850 ) );
  INV_X1 us13_U321 (.A( us13_n785 ) , .ZN( us13_n846 ) );
  AOI22_X1 us13_U322 (.ZN( us13_n696 ) , .A1( us13_n830 ) , .B2( us13_n843 ) , .A2( us13_n865 ) , .B1( us13_n868 ) );
  AOI22_X1 us13_U323 (.A2( us13_n782 ) , .ZN( us13_n783 ) , .B2( us13_n831 ) , .A1( us13_n834 ) , .B1( us13_n863 ) );
  AOI21_X1 us13_U324 (.ZN( us13_n443 ) , .B1( us13_n789 ) , .B2( us13_n791 ) , .A( us13_n814 ) );
  NAND2_X1 us13_U325 (.ZN( us13_n714 ) , .A1( us13_n728 ) , .A2( us13_n780 ) );
  OAI21_X1 us13_U326 (.A( us13_n787 ) , .B2( us13_n788 ) , .B1( us13_n789 ) , .ZN( us13_n795 ) );
  OAI21_X1 us13_U327 (.ZN( us13_n787 ) , .A( us13_n839 ) , .B1( us13_n863 ) , .B2( us13_n873 ) );
  NAND2_X1 us13_U328 (.A2( us13_n762 ) , .A1( us13_n806 ) , .ZN( us13_n810 ) );
  NOR2_X1 us13_U329 (.ZN( us13_n484 ) , .A1( us13_n788 ) , .A2( us13_n805 ) );
  AOI211_X1 us13_U33 (.B( us13_n745 ) , .A( us13_n746 ) , .ZN( us13_n759 ) , .C1( us13_n832 ) , .C2( us13_n853 ) );
  NOR2_X1 us13_U330 (.ZN( us13_n470 ) , .A2( us13_n779 ) , .A1( us13_n815 ) );
  NOR2_X1 us13_U331 (.ZN( us13_n712 ) , .A2( us13_n724 ) , .A1( us13_n790 ) );
  NOR2_X1 us13_U332 (.ZN( us13_n526 ) , .A1( us13_n724 ) , .A2( us13_n750 ) );
  NAND2_X1 us13_U333 (.A1( us13_n699 ) , .A2( us13_n729 ) , .ZN( us13_n782 ) );
  NOR2_X1 us13_U334 (.ZN( us13_n518 ) , .A1( us13_n708 ) , .A2( us13_n788 ) );
  INV_X1 us13_U335 (.A( us13_n813 ) , .ZN( us13_n836 ) );
  NAND2_X1 us13_U336 (.ZN( us13_n671 ) , .A1( us13_n806 ) , .A2( us13_n816 ) );
  OAI21_X1 us13_U337 (.A( us13_n698 ) , .ZN( us13_n702 ) , .B2( us13_n750 ) , .B1( us13_n804 ) );
  OAI21_X1 us13_U338 (.ZN( us13_n698 ) , .B2( us13_n833 ) , .B1( us13_n838 ) , .A( us13_n860 ) );
  NAND2_X1 us13_U339 (.A2( us13_n749 ) , .A1( us13_n786 ) , .ZN( us13_n809 ) );
  NOR3_X1 us13_U34 (.A3( us13_n741 ) , .A2( us13_n742 ) , .A1( us13_n743 ) , .ZN( us13_n760 ) );
  INV_X1 us13_U340 (.A( us13_n724 ) , .ZN( us13_n856 ) );
  INV_X1 us13_U341 (.A( us13_n817 ) , .ZN( us13_n844 ) );
  NAND2_X2 us13_U342 (.A1( us13_n451 ) , .A2( us13_n462 ) , .ZN( us13_n790 ) );
  AND2_X1 us13_U343 (.ZN( us13_n732 ) , .A1( us13_n779 ) , .A2( us13_n785 ) );
  OAI222_X1 us13_U344 (.ZN( us13_n617 ) , .B1( us13_n697 ) , .C1( us13_n724 ) , .C2( us13_n747 ) , .B2( us13_n786 ) , .A2( us13_n792 ) , .A1( us13_n816 ) );
  AOI221_X1 us13_U345 (.A( us13_n764 ) , .ZN( us13_n774 ) , .C2( us13_n810 ) , .B2( us13_n835 ) , .C1( us13_n855 ) , .B1( us13_n866 ) );
  AOI21_X1 us13_U346 (.B2( us13_n763 ) , .ZN( us13_n764 ) , .A( us13_n788 ) , .B1( us13_n792 ) );
  INV_X1 us13_U347 (.A( us13_n761 ) , .ZN( us13_n835 ) );
  NAND2_X1 us13_U348 (.A1( us13_n451 ) , .A2( us13_n454 ) , .ZN( us13_n814 ) );
  NAND2_X1 us13_U349 (.A1( us13_n447 ) , .A2( us13_n449 ) , .ZN( us13_n805 ) );
  NOR4_X1 us13_U35 (.A4( us13_n734 ) , .A3( us13_n735 ) , .A2( us13_n736 ) , .A1( us13_n737 ) , .ZN( us13_n738 ) );
  NAND2_X1 us13_U350 (.A1( us13_n453 ) , .A2( us13_n461 ) , .ZN( us13_n744 ) );
  NAND2_X1 us13_U351 (.A1( us13_n455 ) , .A2( us13_n471 ) , .ZN( us13_n803 ) );
  NAND2_X1 us13_U352 (.A1( us13_n455 ) , .A2( us13_n462 ) , .ZN( us13_n750 ) );
  NAND2_X1 us13_U353 (.A1( us13_n451 ) , .A2( us13_n471 ) , .ZN( us13_n816 ) );
  NAND2_X1 us13_U354 (.A1( us13_n452 ) , .A2( us13_n465 ) , .ZN( us13_n669 ) );
  NAND2_X1 us13_U355 (.A2( us13_n448 ) , .A1( us13_n460 ) , .ZN( us13_n728 ) );
  NAND2_X1 us13_U356 (.A2( us13_n453 ) , .A1( us13_n455 ) , .ZN( us13_n806 ) );
  NAND2_X1 us13_U357 (.A1( us13_n453 ) , .A2( us13_n472 ) , .ZN( us13_n785 ) );
  NAND2_X1 us13_U358 (.A2( us13_n454 ) , .A1( us13_n472 ) , .ZN( us13_n779 ) );
  NAND2_X1 us13_U359 (.A2( us13_n464 ) , .A1( us13_n465 ) , .ZN( us13_n812 ) );
  AOI211_X1 us13_U36 (.B( us13_n725 ) , .A( us13_n726 ) , .ZN( us13_n739 ) , .C1( us13_n843 ) , .C2( us13_n855 ) );
  NAND2_X1 us13_U360 (.A1( us13_n441 ) , .A2( us13_n460 ) , .ZN( us13_n699 ) );
  NAND2_X1 us13_U361 (.A2( us13_n449 ) , .A1( us13_n452 ) , .ZN( us13_n763 ) );
  NAND2_X1 us13_U362 (.A2( us13_n448 ) , .A1( us13_n452 ) , .ZN( us13_n729 ) );
  NAND2_X1 us13_U363 (.A1( us13_n447 ) , .A2( us13_n448 ) , .ZN( us13_n786 ) );
  NAND2_X1 us13_U364 (.A2( us13_n461 ) , .A1( us13_n462 ) , .ZN( us13_n747 ) );
  NAND2_X1 us13_U365 (.A1( us13_n462 ) , .A2( us13_n472 ) , .ZN( us13_n788 ) );
  NOR2_X1 us13_U366 (.ZN( us13_n465 ) , .A2( us13_n847 ) , .A1( us13_n848 ) );
  NOR2_X1 us13_U367 (.ZN( us13_n453 ) , .A1( us13_n826 ) , .A2( us13_n827 ) );
  NOR2_X1 us13_U368 (.ZN( us13_n451 ) , .A1( us13_n828 ) , .A2( us13_n829 ) );
  NAND2_X1 us13_U369 (.A2( us13_n461 ) , .A1( us13_n471 ) , .ZN( us13_n697 ) );
  NOR3_X1 us13_U37 (.A3( us13_n722 ) , .A1( us13_n723 ) , .ZN( us13_n740 ) , .A2( us13_n741 ) );
  NAND2_X1 us13_U370 (.A2( us13_n454 ) , .A1( us13_n455 ) , .ZN( us13_n730 ) );
  NAND2_X1 us13_U371 (.A2( us13_n441 ) , .A1( us13_n447 ) , .ZN( us13_n784 ) );
  NAND2_X2 us13_U372 (.A2( us13_n448 ) , .A1( us13_n464 ) , .ZN( us13_n815 ) );
  NAND2_X2 us13_U373 (.A2( us13_n441 ) , .A1( us13_n452 ) , .ZN( us13_n791 ) );
  NAND2_X2 us13_U374 (.A1( us13_n449 ) , .A2( us13_n460 ) , .ZN( us13_n792 ) );
  NAND2_X2 us13_U375 (.A1( us13_n441 ) , .A2( us13_n464 ) , .ZN( us13_n708 ) );
  NAND2_X2 us13_U376 (.A2( us13_n460 ) , .A1( us13_n465 ) , .ZN( us13_n780 ) );
  NOR2_X1 us13_U377 (.ZN( us13_n447 ) , .A2( us13_n849 ) , .A1( us13_n858 ) );
  NOR2_X1 us13_U378 (.A2( sa13_6 ) , .A1( sa13_7 ) , .ZN( us13_n464 ) );
  NOR2_X1 us13_U379 (.A2( sa13_7 ) , .ZN( us13_n460 ) , .A1( us13_n849 ) );
  NAND4_X1 us13_U38 (.ZN( sa12_sr_3 ) , .A4( us13_n704 ) , .A3( us13_n705 ) , .A2( us13_n706 ) , .A1( us13_n707 ) );
  NOR2_X1 us13_U380 (.A2( sa13_4 ) , .ZN( us13_n449 ) , .A1( us13_n848 ) );
  NOR2_X1 us13_U381 (.A2( sa13_4 ) , .A1( sa13_5 ) , .ZN( us13_n441 ) );
  NOR2_X1 us13_U382 (.A2( sa13_5 ) , .ZN( us13_n448 ) , .A1( us13_n847 ) );
  NOR2_X1 us13_U383 (.A2( sa13_1 ) , .ZN( us13_n471 ) , .A1( us13_n826 ) );
  NOR2_X1 us13_U384 (.A2( sa13_2 ) , .A1( sa13_3 ) , .ZN( us13_n472 ) );
  NOR2_X1 us13_U385 (.A2( sa13_6 ) , .ZN( us13_n452 ) , .A1( us13_n858 ) );
  NOR2_X1 us13_U386 (.A2( sa13_0 ) , .A1( sa13_1 ) , .ZN( us13_n462 ) );
  NOR2_X1 us13_U387 (.A2( sa13_3 ) , .ZN( us13_n455 ) , .A1( us13_n828 ) );
  NOR2_X1 us13_U388 (.A2( sa13_2 ) , .ZN( us13_n461 ) , .A1( us13_n829 ) );
  NOR2_X1 us13_U389 (.A2( sa13_0 ) , .ZN( us13_n454 ) , .A1( us13_n827 ) );
  NOR4_X1 us13_U39 (.A4( us13_n700 ) , .A3( us13_n701 ) , .A2( us13_n702 ) , .A1( us13_n703 ) , .ZN( us13_n704 ) );
  INV_X1 us13_U390 (.A( sa13_4 ) , .ZN( us13_n847 ) );
  INV_X1 us13_U391 (.A( sa13_6 ) , .ZN( us13_n849 ) );
  INV_X1 us13_U392 (.A( sa13_1 ) , .ZN( us13_n827 ) );
  INV_X1 us13_U393 (.A( sa13_3 ) , .ZN( us13_n829 ) );
  INV_X1 us13_U394 (.A( sa13_0 ) , .ZN( us13_n826 ) );
  INV_X1 us13_U395 (.A( sa13_2 ) , .ZN( us13_n828 ) );
  INV_X1 us13_U396 (.A( sa13_7 ) , .ZN( us13_n858 ) );
  INV_X1 us13_U397 (.A( sa13_5 ) , .ZN( us13_n848 ) );
  AOI21_X1 us13_U398 (.ZN( us13_n500 ) , .A( us13_n697 ) , .B1( us13_n708 ) , .B2( us13_n786 ) );
  INV_X1 us13_U399 (.A( us13_n697 ) , .ZN( us13_n838 ) );
  NAND2_X1 us13_U4 (.A1( us13_n449 ) , .A2( us13_n464 ) , .ZN( us13_n724 ) );
  AOI211_X1 us13_U40 (.B( us13_n694 ) , .A( us13_n695 ) , .ZN( us13_n705 ) , .C2( us13_n831 ) , .C1( us13_n851 ) );
  AOI21_X1 us13_U400 (.ZN( us13_n571 ) , .B2( us13_n697 ) , .B1( us13_n806 ) , .A( us13_n812 ) );
  NOR2_X1 us13_U401 (.A1( us13_n697 ) , .ZN( us13_n770 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U402 (.ZN( us13_n566 ) , .A2( us13_n697 ) , .A1( us13_n763 ) );
  AOI21_X1 us13_U403 (.ZN( us13_n552 ) , .B1( us13_n669 ) , .A( us13_n697 ) , .B2( us13_n805 ) );
  NOR2_X1 us13_U404 (.ZN( us13_n632 ) , .A2( us13_n697 ) , .A1( us13_n724 ) );
  NOR2_X1 us13_U405 (.ZN( us13_n541 ) , .A2( us13_n697 ) , .A1( us13_n699 ) );
  AOI21_X1 us13_U406 (.ZN( us13_n478 ) , .B2( us13_n697 ) , .A( us13_n749 ) , .B1( us13_n779 ) );
  NOR2_X1 us13_U407 (.A2( us13_n697 ) , .A1( us13_n780 ) , .ZN( us13_n820 ) );
  NOR2_X1 us13_U408 (.ZN( us13_n662 ) , .A2( us13_n697 ) , .A1( us13_n729 ) );
  NOR2_X1 us13_U409 (.A2( us13_n697 ) , .ZN( us13_n716 ) , .A1( us13_n792 ) );
  NOR2_X1 us13_U41 (.ZN( us13_n707 ) , .A2( us13_n776 ) , .A1( us13_n800 ) );
  NOR2_X1 us13_U410 (.ZN( us13_n594 ) , .A2( us13_n697 ) , .A1( us13_n728 ) );
  NOR2_X1 us13_U411 (.ZN( us13_n580 ) , .A2( us13_n697 ) , .A1( us13_n791 ) );
  OAI221_X1 us13_U412 (.A( us13_n783 ) , .C2( us13_n784 ) , .B2( us13_n785 ) , .B1( us13_n786 ) , .ZN( us13_n796 ) , .C1( us13_n813 ) );
  OAI22_X1 us13_U413 (.ZN( us13_n588 ) , .A2( us13_n747 ) , .B2( us13_n762 ) , .A1( us13_n763 ) , .B1( us13_n784 ) );
  AOI21_X1 us13_U414 (.ZN( us13_n592 ) , .B1( us13_n728 ) , .B2( us13_n784 ) , .A( us13_n790 ) );
  OAI221_X1 us13_U415 (.A( us13_n696 ) , .ZN( us13_n703 ) , .C2( us13_n784 ) , .C1( us13_n785 ) , .B1( us13_n786 ) , .B2( us13_n806 ) );
  NAND2_X1 us13_U416 (.A1( us13_n729 ) , .A2( us13_n784 ) , .ZN( us13_n811 ) );
  AOI21_X1 us13_U417 (.ZN( us13_n623 ) , .B1( us13_n699 ) , .A( us13_n779 ) , .B2( us13_n784 ) );
  AOI21_X1 us13_U418 (.ZN( us13_n648 ) , .A( us13_n762 ) , .B2( us13_n784 ) , .B1( us13_n792 ) );
  OAI22_X1 us13_U419 (.ZN( us13_n681 ) , .A1( us13_n699 ) , .A2( us13_n730 ) , .B2( us13_n784 ) , .B1( us13_n817 ) );
  NOR2_X1 us13_U42 (.ZN( us13_n804 ) , .A1( us13_n854 ) , .A2( us13_n861 ) );
  NOR2_X1 us13_U420 (.ZN( us13_n651 ) , .A1( us13_n784 ) , .A2( us13_n788 ) );
  NOR2_X1 us13_U421 (.ZN( us13_n553 ) , .A2( us13_n744 ) , .A1( us13_n784 ) );
  OAI21_X1 us13_U422 (.A( us13_n613 ) , .ZN( us13_n616 ) , .B1( us13_n625 ) , .B2( us13_n784 ) );
  NOR2_X1 us13_U423 (.ZN( us13_n610 ) , .A1( us13_n784 ) , .A2( us13_n816 ) );
  OAI222_X1 us13_U424 (.A2( us13_n669 ) , .ZN( us13_n674 ) , .B1( us13_n747 ) , .B2( us13_n784 ) , .C2( us13_n788 ) , .C1( us13_n815 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U425 (.ZN( us13_n600 ) , .A2( us13_n697 ) , .A1( us13_n784 ) );
  INV_X1 us13_U426 (.A( us13_n784 ) , .ZN( us13_n861 ) );
  NAND2_X1 us13_U427 (.A1( us13_n454 ) , .A2( us13_n461 ) , .ZN( us13_n813 ) );
  NOR2_X1 us13_U428 (.ZN( us13_n789 ) , .A2( us13_n862 ) , .A1( us13_n868 ) );
  AOI221_X1 us13_U429 (.A( us13_n483 ) , .ZN( us13_n488 ) , .B1( us13_n831 ) , .C2( us13_n844 ) , .C1( us13_n852 ) , .B2( us13_n862 ) );
  AOI222_X1 us13_U43 (.B2( us13_n638 ) , .ZN( us13_n644 ) , .B1( us13_n841 ) , .A1( us13_n842 ) , .C2( us13_n846 ) , .C1( us13_n863 ) , .A2( us13_n865 ) );
  AOI221_X1 us13_U430 (.A( us13_n681 ) , .ZN( us13_n692 ) , .B2( us13_n840 ) , .C1( us13_n842 ) , .C2( us13_n862 ) , .B1( us13_n865 ) );
  AOI222_X1 us13_U431 (.ZN( us13_n605 ) , .B2( us13_n671 ) , .B1( us13_n753 ) , .C2( us13_n831 ) , .A1( us13_n833 ) , .A2( us13_n862 ) , .C1( us13_n863 ) );
  INV_X1 us13_U432 (.A( us13_n786 ) , .ZN( us13_n862 ) );
  AND2_X1 us13_U433 (.ZN( us13_n438 ) , .A2( us13_n831 ) , .A1( us13_n854 ) );
  AND2_X1 us13_U434 (.ZN( us13_n439 ) , .A2( us13_n843 ) , .A1( us13_n861 ) );
  NOR3_X1 us13_U435 (.A1( us13_n438 ) , .A2( us13_n439 ) , .A3( us13_n576 ) , .ZN( us13_n587 ) );
  INV_X1 us13_U436 (.A( us13_n812 ) , .ZN( us13_n854 ) );
  NAND3_X1 us13_U437 (.ZN( sa12_sr_6 ) , .A3( us13_n797 ) , .A2( us13_n798 ) , .A1( us13_n799 ) );
  NAND3_X1 us13_U438 (.ZN( sa12_sr_5 ) , .A3( us13_n758 ) , .A2( us13_n759 ) , .A1( us13_n760 ) );
  NAND3_X1 us13_U439 (.ZN( sa12_sr_4 ) , .A3( us13_n738 ) , .A2( us13_n739 ) , .A1( us13_n740 ) );
  NOR4_X1 us13_U44 (.A4( us13_n639 ) , .A3( us13_n640 ) , .A2( us13_n641 ) , .A1( us13_n642 ) , .ZN( us13_n643 ) );
  NAND3_X1 us13_U440 (.A3( us13_n675 ) , .A2( us13_n676 ) , .A1( us13_n677 ) , .ZN( us13_n807 ) );
  NAND3_X1 us13_U441 (.ZN( us13_n638 ) , .A3( us13_n708 ) , .A2( us13_n724 ) , .A1( us13_n792 ) );
  NAND3_X1 us13_U442 (.A3( us13_n618 ) , .A2( us13_n619 ) , .A1( us13_n620 ) , .ZN( us13_n725 ) );
  NAND3_X1 us13_U443 (.A3( us13_n585 ) , .A2( us13_n586 ) , .A1( us13_n587 ) , .ZN( us13_n621 ) );
  NAND3_X1 us13_U444 (.ZN( us13_n565 ) , .A3( us13_n680 ) , .A2( us13_n750 ) , .A1( us13_n785 ) );
  NAND3_X1 us13_U445 (.A3( us13_n523 ) , .A2( us13_n524 ) , .A1( us13_n525 ) , .ZN( us13_n742 ) );
  NAND3_X1 us13_U446 (.A3( us13_n512 ) , .A1( us13_n513 ) , .ZN( us13_n608 ) , .A2( us13_n871 ) );
  NAND3_X1 us13_U447 (.A3( us13_n467 ) , .A2( us13_n468 ) , .A1( us13_n469 ) , .ZN( us13_n777 ) );
  INV_X1 us13_U448 (.A( us13_n803 ) , .ZN( us13_n843 ) );
  AOI21_X1 us13_U449 (.ZN( us13_n576 ) , .B2( us13_n724 ) , .B1( us13_n748 ) , .A( us13_n785 ) );
  NOR3_X1 us13_U45 (.A2( us13_n607 ) , .A1( us13_n608 ) , .ZN( us13_n646 ) , .A3( us13_n722 ) );
  NAND4_X1 us13_U46 (.ZN( sa12_sr_0 ) , .A4( us13_n501 ) , .A3( us13_n502 ) , .A2( us13_n503 ) , .A1( us13_n504 ) );
  AOI221_X1 us13_U47 (.A( us13_n497 ) , .ZN( us13_n502 ) , .B2( us13_n843 ) , .C1( us13_n846 ) , .C2( us13_n860 ) , .B1( us13_n862 ) );
  NOR4_X1 us13_U48 (.A4( us13_n498 ) , .A3( us13_n499 ) , .A2( us13_n500 ) , .ZN( us13_n501 ) , .A1( us13_n527 ) );
  AOI211_X1 us13_U49 (.A( us13_n496 ) , .ZN( us13_n503 ) , .B( us13_n802 ) , .C2( us13_n839 ) , .C1( us13_n851 ) );
  NAND2_X1 us13_U5 (.A2( us13_n471 ) , .A1( us13_n472 ) , .ZN( us13_n817 ) );
  NAND4_X1 us13_U50 (.ZN( sa12_sr_1 ) , .A4( us13_n595 ) , .A3( us13_n596 ) , .A2( us13_n597 ) , .A1( us13_n598 ) );
  AOI211_X1 us13_U51 (.B( us13_n589 ) , .A( us13_n590 ) , .ZN( us13_n596 ) , .C2( us13_n811 ) , .C1( us13_n833 ) );
  NOR4_X1 us13_U52 (.A4( us13_n591 ) , .A3( us13_n592 ) , .A2( us13_n593 ) , .A1( us13_n594 ) , .ZN( us13_n595 ) );
  AOI211_X1 us13_U53 (.A( us13_n588 ) , .ZN( us13_n597 ) , .B( us13_n621 ) , .C1( us13_n845 ) , .C2( us13_n855 ) );
  NOR2_X1 us13_U54 (.ZN( us13_n748 ) , .A1( us13_n861 ) , .A2( us13_n862 ) );
  NAND4_X1 us13_U55 (.ZN( sa12_sr_7 ) , .A4( us13_n822 ) , .A3( us13_n823 ) , .A2( us13_n824 ) , .A1( us13_n825 ) );
  AOI222_X1 us13_U56 (.C2( us13_n809 ) , .B2( us13_n810 ) , .A2( us13_n811 ) , .ZN( us13_n823 ) , .C1( us13_n832 ) , .A1( us13_n839 ) , .B1( us13_n853 ) );
  NOR4_X1 us13_U57 (.A4( us13_n818 ) , .A3( us13_n819 ) , .A2( us13_n820 ) , .A1( us13_n821 ) , .ZN( us13_n822 ) );
  AOI211_X1 us13_U58 (.B( us13_n807 ) , .A( us13_n808 ) , .ZN( us13_n824 ) , .C1( us13_n842 ) , .C2( us13_n850 ) );
  NOR2_X1 us13_U59 (.ZN( us13_n625 ) , .A2( us13_n836 ) , .A1( us13_n839 ) );
  NOR3_X1 us13_U6 (.ZN( us13_n598 ) , .A1( us13_n608 ) , .A3( us13_n723 ) , .A2( us13_n742 ) );
  NAND4_X1 us13_U60 (.A4( us13_n603 ) , .A3( us13_n604 ) , .A2( us13_n605 ) , .A1( us13_n606 ) , .ZN( us13_n722 ) );
  NOR3_X1 us13_U61 (.A1( us13_n599 ) , .ZN( us13_n604 ) , .A3( us13_n663 ) , .A2( us13_n770 ) );
  NOR4_X1 us13_U62 (.A3( us13_n600 ) , .A2( us13_n601 ) , .A1( us13_n602 ) , .ZN( us13_n603 ) , .A4( us13_n655 ) );
  AOI222_X1 us13_U63 (.ZN( us13_n606 ) , .A1( us13_n830 ) , .C2( us13_n837 ) , .B1( us13_n842 ) , .A2( us13_n856 ) , .B2( us13_n861 ) , .C1( us13_n868 ) );
  AOI222_X1 us13_U64 (.ZN( us13_n469 ) , .B1( us13_n832 ) , .A1( us13_n839 ) , .C1( us13_n842 ) , .C2( us13_n851 ) , .A2( us13_n855 ) , .B2( us13_n865 ) );
  NOR4_X1 us13_U65 (.A1( us13_n466 ) , .ZN( us13_n467 ) , .A4( us13_n542 ) , .A2( us13_n554 ) , .A3( us13_n614 ) );
  AOI221_X1 us13_U66 (.ZN( us13_n468 ) , .C2( us13_n714 ) , .B2( us13_n831 ) , .C1( us13_n845 ) , .B1( us13_n860 ) , .A( us13_n864 ) );
  NAND4_X1 us13_U67 (.A4( us13_n485 ) , .A3( us13_n486 ) , .A2( us13_n487 ) , .A1( us13_n488 ) , .ZN( us13_n778 ) );
  NOR4_X1 us13_U68 (.A4( us13_n484 ) , .ZN( us13_n487 ) , .A1( us13_n566 ) , .A2( us13_n581 ) , .A3( us13_n602 ) );
  NOR4_X1 us13_U69 (.ZN( us13_n486 ) , .A1( us13_n507 ) , .A2( us13_n519 ) , .A4( us13_n546 ) , .A3( us13_n611 ) );
  NOR3_X1 us13_U7 (.A3( us13_n800 ) , .A2( us13_n801 ) , .A1( us13_n802 ) , .ZN( us13_n825 ) );
  NOR4_X1 us13_U70 (.A4( us13_n514 ) , .A3( us13_n515 ) , .A2( us13_n516 ) , .A1( us13_n517 ) , .ZN( us13_n524 ) );
  AOI222_X1 us13_U71 (.ZN( us13_n525 ) , .A1( us13_n834 ) , .B2( us13_n837 ) , .C1( us13_n844 ) , .C2( us13_n850 ) , .A2( us13_n852 ) , .B1( us13_n866 ) );
  NOR4_X1 us13_U72 (.A3( us13_n521 ) , .A1( us13_n522 ) , .ZN( us13_n523 ) , .A2( us13_n673 ) , .A4( us13_n769 ) );
  NAND4_X1 us13_U73 (.A4( us13_n657 ) , .A3( us13_n658 ) , .A2( us13_n659 ) , .A1( us13_n660 ) , .ZN( us13_n800 ) );
  NOR3_X1 us13_U74 (.A3( us13_n651 ) , .A2( us13_n652 ) , .A1( us13_n653 ) , .ZN( us13_n658 ) );
  NOR3_X1 us13_U75 (.A3( us13_n648 ) , .A2( us13_n649 ) , .A1( us13_n650 ) , .ZN( us13_n659 ) );
  NOR3_X1 us13_U76 (.A3( us13_n654 ) , .A2( us13_n655 ) , .A1( us13_n656 ) , .ZN( us13_n657 ) );
  NAND4_X1 us13_U77 (.A4( us13_n560 ) , .A3( us13_n561 ) , .A2( us13_n562 ) , .A1( us13_n563 ) , .ZN( us13_n607 ) );
  NOR4_X1 us13_U78 (.A4( us13_n552 ) , .A3( us13_n553 ) , .A2( us13_n554 ) , .A1( us13_n555 ) , .ZN( us13_n562 ) );
  NOR4_X1 us13_U79 (.ZN( us13_n561 ) , .A1( us13_n653 ) , .A3( us13_n661 ) , .A4( us13_n685 ) , .A2( us13_n768 ) );
  NOR3_X1 us13_U8 (.ZN( us13_n504 ) , .A2( us13_n679 ) , .A3( us13_n777 ) , .A1( us13_n876 ) );
  NOR4_X1 us13_U80 (.A4( us13_n556 ) , .A3( us13_n557 ) , .A2( us13_n558 ) , .A1( us13_n559 ) , .ZN( us13_n560 ) );
  NAND4_X1 us13_U81 (.A4( us13_n772 ) , .A3( us13_n773 ) , .A2( us13_n774 ) , .A1( us13_n775 ) , .ZN( us13_n801 ) );
  NOR3_X1 us13_U82 (.A3( us13_n765 ) , .A2( us13_n766 ) , .A1( us13_n767 ) , .ZN( us13_n773 ) );
  AOI222_X1 us13_U83 (.ZN( us13_n775 ) , .A1( us13_n830 ) , .C1( us13_n834 ) , .B2( us13_n841 ) , .A2( us13_n850 ) , .B1( us13_n861 ) , .C2( us13_n873 ) );
  NOR4_X1 us13_U84 (.A4( us13_n768 ) , .A3( us13_n769 ) , .A2( us13_n770 ) , .A1( us13_n771 ) , .ZN( us13_n772 ) );
  NAND4_X1 us13_U85 (.A4( us13_n691 ) , .A3( us13_n692 ) , .A1( us13_n693 ) , .ZN( us13_n776 ) , .A2( us13_n872 ) );
  INV_X1 us13_U86 (.A( us13_n679 ) , .ZN( us13_n872 ) );
  NOR4_X1 us13_U87 (.A4( us13_n687 ) , .A3( us13_n688 ) , .A2( us13_n689 ) , .A1( us13_n690 ) , .ZN( us13_n691 ) );
  NOR4_X1 us13_U88 (.A4( us13_n661 ) , .A3( us13_n662 ) , .A2( us13_n663 ) , .A1( us13_n664 ) , .ZN( us13_n677 ) );
  NOR4_X1 us13_U89 (.A4( us13_n665 ) , .A3( us13_n666 ) , .A2( us13_n667 ) , .A1( us13_n668 ) , .ZN( us13_n676 ) );
  INV_X1 us13_U9 (.A( us13_n706 ) , .ZN( us13_n876 ) );
  NOR4_X1 us13_U90 (.A3( us13_n673 ) , .A1( us13_n674 ) , .ZN( us13_n675 ) , .A4( us13_n715 ) , .A2( us13_n859 ) );
  NOR2_X1 us13_U91 (.ZN( us13_n761 ) , .A1( us13_n833 ) , .A2( us13_n834 ) );
  NOR4_X1 us13_U92 (.A4( us13_n577 ) , .A3( us13_n578 ) , .A2( us13_n579 ) , .ZN( us13_n586 ) , .A1( us13_n683 ) );
  NOR4_X1 us13_U93 (.A1( us13_n584 ) , .ZN( us13_n585 ) , .A3( us13_n652 ) , .A2( us13_n662 ) , .A4( us13_n767 ) );
  AOI222_X1 us13_U94 (.ZN( us13_n513 ) , .C1( us13_n832 ) , .B2( us13_n837 ) , .A2( us13_n843 ) , .C2( us13_n862 ) , .B1( us13_n863 ) , .A1( us13_n866 ) );
  NOR4_X1 us13_U95 (.A4( us13_n509 ) , .A2( us13_n510 ) , .A1( us13_n511 ) , .ZN( us13_n512 ) , .A3( us13_n670 ) );
  INV_X1 us13_U96 (.A( us13_n505 ) , .ZN( us13_n871 ) );
  NAND4_X1 us13_U97 (.A4( us13_n456 ) , .A3( us13_n457 ) , .A2( us13_n458 ) , .A1( us13_n459 ) , .ZN( us13_n679 ) );
  NOR3_X1 us13_U98 (.ZN( us13_n457 ) , .A3( us13_n530 ) , .A1( us13_n555 ) , .A2( us13_n570 ) );
  AOI221_X1 us13_U99 (.A( us13_n450 ) , .ZN( us13_n459 ) , .C2( us13_n753 ) , .B1( us13_n832 ) , .C1( us13_n842 ) , .B2( us13_n861 ) );
endmodule

