module aes_aes_die_6 ( sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa22_0, 
       sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, u0_n268, u0_n270, 
       u0_n272, u0_n274, w3_10, w3_11, w3_8, w3_9, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa20_sr_0, 
        sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, u0_subword_16, u0_subword_17, 
        u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23 );
  input sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa22_0, 
        sa22_1, sa22_2, sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, u0_n268, u0_n270, 
        u0_n272, u0_n274, w3_10, w3_11, w3_8, w3_9;
  output sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa20_sr_0, 
        sa20_sr_1, sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, u0_subword_16, u0_subword_17, 
        u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23;
  wire u0_u1_n41, u0_u1_n438, u0_u1_n439, u0_u1_n440, u0_u1_n441, u0_u1_n442, u0_u1_n443, u0_u1_n444, u0_u1_n445, 
       u0_u1_n446, u0_u1_n447, u0_u1_n448, u0_u1_n449, u0_u1_n450, u0_u1_n451, u0_u1_n452, u0_u1_n453, u0_u1_n454, 
       u0_u1_n455, u0_u1_n456, u0_u1_n457, u0_u1_n458, u0_u1_n459, u0_u1_n460, u0_u1_n461, u0_u1_n462, u0_u1_n463, 
       u0_u1_n464, u0_u1_n465, u0_u1_n466, u0_u1_n467, u0_u1_n468, u0_u1_n469, u0_u1_n470, u0_u1_n471, u0_u1_n472, 
       u0_u1_n473, u0_u1_n474, u0_u1_n475, u0_u1_n476, u0_u1_n477, u0_u1_n478, u0_u1_n479, u0_u1_n480, u0_u1_n481, 
       u0_u1_n482, u0_u1_n483, u0_u1_n484, u0_u1_n485, u0_u1_n486, u0_u1_n487, u0_u1_n488, u0_u1_n489, u0_u1_n490, 
       u0_u1_n491, u0_u1_n492, u0_u1_n493, u0_u1_n494, u0_u1_n495, u0_u1_n496, u0_u1_n497, u0_u1_n498, u0_u1_n499, 
       u0_u1_n500, u0_u1_n501, u0_u1_n502, u0_u1_n503, u0_u1_n504, u0_u1_n505, u0_u1_n506, u0_u1_n507, u0_u1_n508, 
       u0_u1_n509, u0_u1_n510, u0_u1_n511, u0_u1_n512, u0_u1_n513, u0_u1_n514, u0_u1_n515, u0_u1_n516, u0_u1_n517, 
       u0_u1_n518, u0_u1_n519, u0_u1_n520, u0_u1_n521, u0_u1_n522, u0_u1_n523, u0_u1_n524, u0_u1_n525, u0_u1_n526, 
       u0_u1_n527, u0_u1_n528, u0_u1_n529, u0_u1_n530, u0_u1_n531, u0_u1_n532, u0_u1_n533, u0_u1_n534, u0_u1_n535, 
       u0_u1_n536, u0_u1_n537, u0_u1_n538, u0_u1_n539, u0_u1_n540, u0_u1_n541, u0_u1_n542, u0_u1_n543, u0_u1_n544, 
       u0_u1_n545, u0_u1_n546, u0_u1_n547, u0_u1_n548, u0_u1_n549, u0_u1_n550, u0_u1_n551, u0_u1_n552, u0_u1_n553, 
       u0_u1_n554, u0_u1_n555, u0_u1_n556, u0_u1_n557, u0_u1_n558, u0_u1_n559, u0_u1_n560, u0_u1_n561, u0_u1_n562, 
       u0_u1_n563, u0_u1_n564, u0_u1_n565, u0_u1_n566, u0_u1_n567, u0_u1_n568, u0_u1_n569, u0_u1_n570, u0_u1_n571, 
       u0_u1_n572, u0_u1_n573, u0_u1_n574, u0_u1_n575, u0_u1_n576, u0_u1_n577, u0_u1_n578, u0_u1_n579, u0_u1_n580, 
       u0_u1_n581, u0_u1_n582, u0_u1_n583, u0_u1_n584, u0_u1_n585, u0_u1_n586, u0_u1_n587, u0_u1_n588, u0_u1_n589, 
       u0_u1_n590, u0_u1_n591, u0_u1_n592, u0_u1_n593, u0_u1_n594, u0_u1_n595, u0_u1_n596, u0_u1_n597, u0_u1_n598, 
       u0_u1_n599, u0_u1_n600, u0_u1_n601, u0_u1_n602, u0_u1_n603, u0_u1_n604, u0_u1_n605, u0_u1_n606, u0_u1_n607, 
       u0_u1_n608, u0_u1_n609, u0_u1_n610, u0_u1_n611, u0_u1_n612, u0_u1_n613, u0_u1_n614, u0_u1_n615, u0_u1_n616, 
       u0_u1_n617, u0_u1_n618, u0_u1_n619, u0_u1_n620, u0_u1_n621, u0_u1_n622, u0_u1_n623, u0_u1_n624, u0_u1_n625, 
       u0_u1_n626, u0_u1_n627, u0_u1_n628, u0_u1_n629, u0_u1_n630, u0_u1_n631, u0_u1_n632, u0_u1_n633, u0_u1_n634, 
       u0_u1_n635, u0_u1_n636, u0_u1_n637, u0_u1_n638, u0_u1_n639, u0_u1_n640, u0_u1_n641, u0_u1_n642, u0_u1_n643, 
       u0_u1_n644, u0_u1_n645, u0_u1_n646, u0_u1_n647, u0_u1_n648, u0_u1_n649, u0_u1_n650, u0_u1_n651, u0_u1_n652, 
       u0_u1_n653, u0_u1_n654, u0_u1_n655, u0_u1_n656, u0_u1_n657, u0_u1_n658, u0_u1_n659, u0_u1_n660, u0_u1_n661, 
       u0_u1_n662, u0_u1_n663, u0_u1_n664, u0_u1_n665, u0_u1_n666, u0_u1_n667, u0_u1_n668, u0_u1_n669, u0_u1_n670, 
       u0_u1_n671, u0_u1_n672, u0_u1_n673, u0_u1_n674, u0_u1_n675, u0_u1_n676, u0_u1_n677, u0_u1_n678, u0_u1_n679, 
       u0_u1_n680, u0_u1_n681, u0_u1_n682, u0_u1_n683, u0_u1_n684, u0_u1_n685, u0_u1_n686, u0_u1_n687, u0_u1_n688, 
       u0_u1_n689, u0_u1_n690, u0_u1_n691, u0_u1_n692, u0_u1_n693, u0_u1_n694, u0_u1_n695, u0_u1_n696, u0_u1_n697, 
       u0_u1_n698, u0_u1_n699, u0_u1_n700, u0_u1_n701, u0_u1_n702, u0_u1_n703, u0_u1_n704, u0_u1_n705, u0_u1_n706, 
       u0_u1_n707, u0_u1_n708, u0_u1_n709, u0_u1_n710, u0_u1_n711, u0_u1_n712, u0_u1_n713, u0_u1_n714, u0_u1_n715, 
       u0_u1_n716, u0_u1_n717, u0_u1_n718, u0_u1_n719, u0_u1_n720, u0_u1_n721, u0_u1_n722, u0_u1_n723, u0_u1_n724, 
       u0_u1_n725, u0_u1_n726, u0_u1_n727, u0_u1_n728, u0_u1_n729, u0_u1_n730, u0_u1_n731, u0_u1_n732, u0_u1_n733, 
       u0_u1_n734, u0_u1_n735, u0_u1_n736, u0_u1_n737, u0_u1_n738, u0_u1_n739, u0_u1_n740, u0_u1_n741, u0_u1_n742, 
       u0_u1_n743, u0_u1_n744, u0_u1_n745, u0_u1_n746, u0_u1_n747, u0_u1_n748, u0_u1_n749, u0_u1_n750, u0_u1_n751, 
       u0_u1_n752, u0_u1_n753, u0_u1_n754, u0_u1_n755, u0_u1_n756, u0_u1_n757, u0_u1_n758, u0_u1_n759, u0_u1_n760, 
       u0_u1_n761, u0_u1_n762, u0_u1_n763, u0_u1_n764, u0_u1_n765, u0_u1_n766, u0_u1_n767, u0_u1_n768, u0_u1_n769, 
       u0_u1_n770, u0_u1_n771, u0_u1_n772, u0_u1_n773, u0_u1_n774, u0_u1_n775, u0_u1_n776, u0_u1_n777, u0_u1_n778, 
       u0_u1_n779, u0_u1_n780, u0_u1_n781, u0_u1_n782, u0_u1_n783, u0_u1_n784, u0_u1_n785, u0_u1_n786, u0_u1_n787, 
       u0_u1_n788, u0_u1_n789, u0_u1_n790, u0_u1_n791, u0_u1_n792, u0_u1_n793, u0_u1_n794, u0_u1_n795, u0_u1_n796, 
       u0_u1_n797, u0_u1_n798, u0_u1_n799, u0_u1_n800, u0_u1_n801, u0_u1_n802, u0_u1_n803, u0_u1_n804, u0_u1_n805, 
       u0_u1_n806, u0_u1_n807, u0_u1_n808, u0_u1_n809, u0_u1_n810, u0_u1_n811, u0_u1_n812, u0_u1_n813, u0_u1_n814, 
       u0_u1_n815, u0_u1_n816, u0_u1_n817, u0_u1_n818, u0_u1_n819, u0_u1_n820, u0_u1_n821, u0_u1_n822, u0_u1_n823, 
       u0_u1_n824, u0_u1_n825, u0_u1_n826, u0_u1_n827, u0_u1_n828, u0_u1_n829, u0_u1_n830, u0_u1_n831, u0_u1_n832, 
       u0_u1_n833, u0_u1_n834, u0_u1_n835, u0_u1_n836, u0_u1_n837, u0_u1_n838, u0_u1_n839, u0_u1_n840, u0_u1_n841, 
       u0_u1_n842, u0_u1_n843, u0_u1_n844, u0_u1_n845, u0_u1_n846, u0_u1_n847, u0_u1_n848, u0_u1_n849, u0_u1_n850, 
       u0_u1_n851, u0_u1_n852, u0_u1_n853, u0_u1_n854, u0_u1_n855, u0_u1_n856, u0_u1_n857, u0_u1_n858, u0_u1_n859, 
       u0_u1_n860, u0_u1_n861, u0_u1_n862, u0_u1_n863, u0_u1_n864, u0_u1_n865, u0_u1_n866, u0_u1_n867, u0_u1_n868, 
       u0_u1_n869, u0_u1_n870, u0_u1_n871, u0_u1_n872, u0_u1_n873, u0_u1_n874, u0_u1_n875, u0_u1_n876, u0_u1_n877, 
       us11_n438, us11_n439, us11_n440, us11_n441, us11_n442, us11_n443, us11_n444, us11_n445, us11_n446, 
       us11_n447, us11_n448, us11_n449, us11_n450, us11_n451, us11_n452, us11_n453, us11_n454, us11_n455, 
       us11_n456, us11_n457, us11_n458, us11_n459, us11_n460, us11_n461, us11_n462, us11_n463, us11_n464, 
       us11_n465, us11_n466, us11_n467, us11_n468, us11_n469, us11_n470, us11_n471, us11_n472, us11_n473, 
       us11_n474, us11_n475, us11_n476, us11_n477, us11_n478, us11_n479, us11_n480, us11_n481, us11_n482, 
       us11_n483, us11_n484, us11_n485, us11_n486, us11_n487, us11_n488, us11_n489, us11_n490, us11_n491, 
       us11_n492, us11_n493, us11_n494, us11_n495, us11_n496, us11_n497, us11_n498, us11_n499, us11_n500, 
       us11_n501, us11_n502, us11_n503, us11_n504, us11_n505, us11_n506, us11_n507, us11_n508, us11_n509, 
       us11_n510, us11_n511, us11_n512, us11_n513, us11_n514, us11_n515, us11_n516, us11_n517, us11_n518, 
       us11_n519, us11_n520, us11_n521, us11_n522, us11_n523, us11_n524, us11_n525, us11_n526, us11_n527, 
       us11_n528, us11_n529, us11_n530, us11_n531, us11_n532, us11_n533, us11_n534, us11_n535, us11_n536, 
       us11_n537, us11_n538, us11_n539, us11_n540, us11_n541, us11_n542, us11_n543, us11_n544, us11_n545, 
       us11_n546, us11_n547, us11_n548, us11_n549, us11_n550, us11_n551, us11_n552, us11_n553, us11_n554, 
       us11_n555, us11_n556, us11_n557, us11_n558, us11_n559, us11_n560, us11_n561, us11_n562, us11_n563, 
       us11_n564, us11_n565, us11_n566, us11_n567, us11_n568, us11_n569, us11_n570, us11_n571, us11_n572, 
       us11_n573, us11_n574, us11_n575, us11_n576, us11_n577, us11_n578, us11_n579, us11_n580, us11_n581, 
       us11_n582, us11_n583, us11_n584, us11_n585, us11_n586, us11_n587, us11_n588, us11_n589, us11_n590, 
       us11_n591, us11_n592, us11_n593, us11_n594, us11_n595, us11_n596, us11_n597, us11_n598, us11_n599, 
       us11_n600, us11_n601, us11_n602, us11_n603, us11_n604, us11_n605, us11_n606, us11_n607, us11_n608, 
       us11_n609, us11_n610, us11_n611, us11_n612, us11_n613, us11_n614, us11_n615, us11_n616, us11_n617, 
       us11_n618, us11_n619, us11_n620, us11_n621, us11_n622, us11_n623, us11_n624, us11_n625, us11_n626, 
       us11_n627, us11_n628, us11_n629, us11_n630, us11_n631, us11_n632, us11_n633, us11_n634, us11_n635, 
       us11_n636, us11_n637, us11_n638, us11_n639, us11_n640, us11_n641, us11_n642, us11_n643, us11_n644, 
       us11_n645, us11_n646, us11_n647, us11_n648, us11_n649, us11_n650, us11_n651, us11_n652, us11_n653, 
       us11_n654, us11_n655, us11_n656, us11_n657, us11_n658, us11_n659, us11_n660, us11_n661, us11_n662, 
       us11_n663, us11_n664, us11_n665, us11_n666, us11_n667, us11_n668, us11_n669, us11_n670, us11_n671, 
       us11_n672, us11_n673, us11_n674, us11_n675, us11_n676, us11_n677, us11_n678, us11_n679, us11_n680, 
       us11_n681, us11_n682, us11_n683, us11_n684, us11_n685, us11_n686, us11_n687, us11_n688, us11_n689, 
       us11_n690, us11_n691, us11_n692, us11_n693, us11_n694, us11_n695, us11_n696, us11_n697, us11_n698, 
       us11_n699, us11_n700, us11_n701, us11_n702, us11_n703, us11_n704, us11_n705, us11_n706, us11_n707, 
       us11_n708, us11_n709, us11_n710, us11_n711, us11_n712, us11_n713, us11_n714, us11_n715, us11_n716, 
       us11_n717, us11_n718, us11_n719, us11_n720, us11_n721, us11_n722, us11_n723, us11_n724, us11_n725, 
       us11_n726, us11_n727, us11_n728, us11_n729, us11_n730, us11_n731, us11_n732, us11_n733, us11_n734, 
       us11_n735, us11_n736, us11_n737, us11_n738, us11_n739, us11_n740, us11_n741, us11_n742, us11_n743, 
       us11_n744, us11_n745, us11_n746, us11_n747, us11_n748, us11_n749, us11_n750, us11_n751, us11_n752, 
       us11_n753, us11_n754, us11_n755, us11_n756, us11_n757, us11_n758, us11_n759, us11_n760, us11_n761, 
       us11_n762, us11_n763, us11_n764, us11_n765, us11_n766, us11_n767, us11_n768, us11_n769, us11_n770, 
       us11_n771, us11_n772, us11_n773, us11_n774, us11_n775, us11_n776, us11_n777, us11_n778, us11_n779, 
       us11_n780, us11_n781, us11_n782, us11_n783, us11_n784, us11_n785, us11_n786, us11_n787, us11_n788, 
       us11_n789, us11_n790, us11_n791, us11_n792, us11_n793, us11_n794, us11_n795, us11_n796, us11_n797, 
       us11_n798, us11_n799, us11_n800, us11_n801, us11_n802, us11_n803, us11_n804, us11_n805, us11_n806, 
       us11_n807, us11_n808, us11_n809, us11_n810, us11_n811, us11_n812, us11_n813, us11_n814, us11_n815, 
       us11_n816, us11_n817, us11_n818, us11_n819, us11_n820, us11_n821, us11_n822, us11_n823, us11_n824, 
       us11_n825, us11_n826, us11_n827, us11_n828, us11_n829, us11_n830, us11_n831, us11_n832, us11_n833, 
       us11_n834, us11_n835, us11_n836, us11_n837, us11_n838, us11_n839, us11_n840, us11_n841, us11_n842, 
       us11_n843, us11_n844, us11_n845, us11_n846, us11_n847, us11_n848, us11_n849, us11_n850, us11_n851, 
       us11_n852, us11_n853, us11_n854, us11_n855, us11_n856, us11_n857, us11_n858, us11_n859, us11_n860, 
       us11_n861, us11_n862, us11_n863, us11_n864, us11_n865, us11_n866, us11_n867, us11_n868, us11_n869, 
       us11_n870, us11_n871, us11_n872, us11_n873, us11_n874, us11_n875, us11_n876, us22_n438, us22_n439, 
       us22_n440, us22_n441, us22_n442, us22_n443, us22_n444, us22_n445, us22_n446, us22_n447, us22_n448, 
       us22_n449, us22_n450, us22_n451, us22_n452, us22_n453, us22_n454, us22_n455, us22_n456, us22_n457, 
       us22_n458, us22_n459, us22_n460, us22_n461, us22_n462, us22_n463, us22_n464, us22_n465, us22_n466, 
       us22_n467, us22_n468, us22_n469, us22_n470, us22_n471, us22_n472, us22_n473, us22_n474, us22_n475, 
       us22_n476, us22_n477, us22_n478, us22_n479, us22_n480, us22_n481, us22_n482, us22_n483, us22_n484, 
       us22_n485, us22_n486, us22_n487, us22_n488, us22_n489, us22_n490, us22_n491, us22_n492, us22_n493, 
       us22_n494, us22_n495, us22_n496, us22_n497, us22_n498, us22_n499, us22_n500, us22_n501, us22_n502, 
       us22_n503, us22_n504, us22_n505, us22_n506, us22_n507, us22_n508, us22_n509, us22_n510, us22_n511, 
       us22_n512, us22_n513, us22_n514, us22_n515, us22_n516, us22_n517, us22_n518, us22_n519, us22_n520, 
       us22_n521, us22_n522, us22_n523, us22_n524, us22_n525, us22_n526, us22_n527, us22_n528, us22_n529, 
       us22_n530, us22_n531, us22_n532, us22_n533, us22_n534, us22_n535, us22_n536, us22_n537, us22_n538, 
       us22_n539, us22_n540, us22_n541, us22_n542, us22_n543, us22_n544, us22_n545, us22_n546, us22_n547, 
       us22_n548, us22_n549, us22_n550, us22_n551, us22_n552, us22_n553, us22_n554, us22_n555, us22_n556, 
       us22_n557, us22_n558, us22_n559, us22_n560, us22_n561, us22_n562, us22_n563, us22_n564, us22_n565, 
       us22_n566, us22_n567, us22_n568, us22_n569, us22_n570, us22_n571, us22_n572, us22_n573, us22_n574, 
       us22_n575, us22_n576, us22_n577, us22_n578, us22_n579, us22_n580, us22_n581, us22_n582, us22_n583, 
       us22_n584, us22_n585, us22_n586, us22_n587, us22_n588, us22_n589, us22_n590, us22_n591, us22_n592, 
       us22_n593, us22_n594, us22_n595, us22_n596, us22_n597, us22_n598, us22_n599, us22_n600, us22_n601, 
       us22_n602, us22_n603, us22_n604, us22_n605, us22_n606, us22_n607, us22_n608, us22_n609, us22_n610, 
       us22_n611, us22_n612, us22_n613, us22_n614, us22_n615, us22_n616, us22_n617, us22_n618, us22_n619, 
       us22_n620, us22_n621, us22_n622, us22_n623, us22_n624, us22_n625, us22_n626, us22_n627, us22_n628, 
       us22_n629, us22_n630, us22_n631, us22_n632, us22_n633, us22_n634, us22_n635, us22_n636, us22_n637, 
       us22_n638, us22_n639, us22_n640, us22_n641, us22_n642, us22_n643, us22_n644, us22_n645, us22_n646, 
       us22_n647, us22_n648, us22_n649, us22_n650, us22_n651, us22_n652, us22_n653, us22_n654, us22_n655, 
       us22_n656, us22_n657, us22_n658, us22_n659, us22_n660, us22_n661, us22_n662, us22_n663, us22_n664, 
       us22_n665, us22_n666, us22_n667, us22_n668, us22_n669, us22_n670, us22_n671, us22_n672, us22_n673, 
       us22_n674, us22_n675, us22_n676, us22_n677, us22_n678, us22_n679, us22_n680, us22_n681, us22_n682, 
       us22_n683, us22_n684, us22_n685, us22_n686, us22_n687, us22_n688, us22_n689, us22_n690, us22_n691, 
       us22_n692, us22_n693, us22_n694, us22_n695, us22_n696, us22_n697, us22_n698, us22_n699, us22_n700, 
       us22_n701, us22_n702, us22_n703, us22_n704, us22_n705, us22_n706, us22_n707, us22_n708, us22_n709, 
       us22_n710, us22_n711, us22_n712, us22_n713, us22_n714, us22_n715, us22_n716, us22_n717, us22_n718, 
       us22_n719, us22_n720, us22_n721, us22_n722, us22_n723, us22_n724, us22_n725, us22_n726, us22_n727, 
       us22_n728, us22_n729, us22_n730, us22_n731, us22_n732, us22_n733, us22_n734, us22_n735, us22_n736, 
       us22_n737, us22_n738, us22_n739, us22_n740, us22_n741, us22_n742, us22_n743, us22_n744, us22_n745, 
       us22_n746, us22_n747, us22_n748, us22_n749, us22_n750, us22_n751, us22_n752, us22_n753, us22_n754, 
       us22_n755, us22_n756, us22_n757, us22_n758, us22_n759, us22_n760, us22_n761, us22_n762, us22_n763, 
       us22_n764, us22_n765, us22_n766, us22_n767, us22_n768, us22_n769, us22_n770, us22_n771, us22_n772, 
       us22_n773, us22_n774, us22_n775, us22_n776, us22_n777, us22_n778, us22_n779, us22_n780, us22_n781, 
       us22_n782, us22_n783, us22_n784, us22_n785, us22_n786, us22_n787, us22_n788, us22_n789, us22_n790, 
       us22_n791, us22_n792, us22_n793, us22_n794, us22_n795, us22_n796, us22_n797, us22_n798, us22_n799, 
       us22_n800, us22_n801, us22_n802, us22_n803, us22_n804, us22_n805, us22_n806, us22_n807, us22_n808, 
       us22_n809, us22_n810, us22_n811, us22_n812, us22_n813, us22_n814, us22_n815, us22_n816, us22_n817, 
       us22_n818, us22_n819, us22_n820, us22_n821, us22_n822, us22_n823, us22_n824, us22_n825, us22_n826, 
       us22_n827, us22_n828, us22_n829, us22_n830, us22_n831, us22_n832, us22_n833, us22_n834, us22_n835, 
       us22_n836, us22_n837, us22_n838, us22_n839, us22_n840, us22_n841, us22_n842, us22_n843, us22_n844, 
       us22_n845, us22_n846, us22_n847, us22_n848, us22_n849, us22_n850, us22_n851, us22_n852, us22_n853, 
       us22_n854, us22_n855, us22_n856, us22_n857, us22_n858, us22_n859, us22_n860, us22_n861, us22_n862, 
       us22_n863, us22_n864, us22_n865, us22_n866, us22_n867, us22_n868, us22_n869, us22_n870, us22_n871, 
       us22_n872, us22_n873,  us22_n874;
  NOR2_X1 u0_u1_U10 (.ZN( u0_u1_n709 ) , .A2( u0_u1_n778 ) , .A1( u0_u1_n802 ) );
  INV_X1 u0_u1_U100 (.A( u0_u1_n819 ) , .ZN( u0_u1_n845 ) );
  INV_X1 u0_u1_U101 (.A( u0_u1_n674 ) , .ZN( u0_u1_n860 ) );
  AOI21_X1 u0_u1_U102 (.A( u0_u1_n672 ) , .B1( u0_u1_n673 ) , .ZN( u0_u1_n674 ) , .B2( u0_u1_n857 ) );
  INV_X1 u0_u1_U103 (.A( u0_u1_n756 ) , .ZN( u0_u1_n870 ) );
  OAI21_X1 u0_u1_U104 (.B1( u0_u1_n755 ) , .ZN( u0_u1_n756 ) , .A( u0_u1_n846 ) , .B2( u0_u1_n869 ) );
  AOI221_X1 u0_u1_U105 (.A( u0_u1_n715 ) , .B2( u0_u1_n716 ) , .ZN( u0_u1_n722 ) , .C1( u0_u1_n834 ) , .B1( u0_u1_n840 ) , .C2( u0_u1_n864 ) );
  OR2_X1 u0_u1_U106 (.A2( u0_u1_n713 ) , .A1( u0_u1_n714 ) , .ZN( u0_u1_n715 ) );
  NAND2_X1 u0_u1_U107 (.A1( u0_u1_n449 ) , .A2( u0_u1_n451 ) , .ZN( u0_u1_n807 ) );
  NOR3_X1 u0_u1_U108 (.ZN( u0_u1_n754 ) , .A2( u0_u1_n854 ) , .A1( u0_u1_n864 ) , .A3( u0_u1_n866 ) );
  NOR2_X1 u0_u1_U109 (.ZN( u0_u1_n753 ) , .A2( u0_u1_n853 ) , .A1( u0_u1_n861 ) );
  NOR2_X1 u0_u1_U11 (.A1( u0_u1_n680 ) , .ZN( u0_u1_n695 ) , .A2( u0_u1_n809 ) );
  INV_X1 u0_u1_U110 (.A( u0_u1_n440 ) , .ZN( u0_u1_n815 ) );
  NAND2_X1 u0_u1_U111 (.A1( u0_u1_n449 ) , .A2( u0_u1_n467 ) , .ZN( u0_u1_n751 ) );
  AOI211_X1 u0_u1_U112 (.B( u0_u1_n809 ) , .A( u0_u1_n810 ) , .ZN( u0_u1_n826 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n851 ) );
  NOR2_X1 u0_u1_U113 (.ZN( u0_u1_n509 ) , .A1( u0_u1_n814 ) , .A2( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U114 (.B1( u0_u1_n492 ) , .ZN( u0_u1_n493 ) , .A1( u0_u1_n688 ) , .A2( u0_u1_n765 ) , .B2( u0_u1_n819 ) );
  NOR3_X1 u0_u1_U115 (.ZN( u0_u1_n492 ) , .A1( u0_u1_n784 ) , .A2( u0_u1_n851 ) , .A3( u0_u1_n864 ) );
  NOR2_X1 u0_u1_U116 (.ZN( u0_u1_n579 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U117 (.ZN( u0_u1_n548 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U118 (.ZN( u0_u1_n508 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n764 ) );
  INV_X1 u0_u1_U119 (.A( u0_u1_n814 ) , .ZN( u0_u1_n855 ) );
  INV_X1 u0_u1_U12 (.A( u0_u1_n609 ) , .ZN( u0_u1_n875 ) );
  NOR2_X1 u0_u1_U120 (.ZN( u0_u1_n534 ) , .A2( u0_u1_n751 ) , .A1( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U121 (.ZN( u0_u1_n603 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U122 (.ZN( u0_u1_n530 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n805 ) );
  INV_X1 u0_u1_U123 (.A( u0_u1_n816 ) , .ZN( u0_u1_n835 ) );
  AOI21_X1 u0_u1_U124 (.B1( u0_u1_n701 ) , .ZN( u0_u1_n702 ) , .A( u0_u1_n734 ) , .B2( u0_u1_n765 ) );
  NOR2_X1 u0_u1_U125 (.ZN( u0_u1_n557 ) , .A1( u0_u1_n752 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U126 (.ZN( u0_u1_n668 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U127 (.ZN( u0_u1_n547 ) , .A1( u0_u1_n751 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U128 (.ZN( u0_u1_n511 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U129 (.A1( u0_u1_n751 ) , .ZN( u0_u1_n769 ) , .A2( u0_u1_n805 ) );
  INV_X1 u0_u1_U13 (.A( u0_u1_n649 ) , .ZN( u0_u1_n871 ) );
  NOR2_X1 u0_u1_U130 (.ZN( u0_u1_n654 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U131 (.ZN( u0_u1_n604 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U132 (.ZN( u0_u1_n658 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n782 ) );
  NOR2_X1 u0_u1_U133 (.ZN( u0_u1_n529 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n781 ) );
  INV_X1 u0_u1_U134 (.A( u0_u1_n701 ) , .ZN( u0_u1_n854 ) );
  NOR2_X1 u0_u1_U135 (.ZN( u0_u1_n611 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n819 ) );
  AOI21_X1 u0_u1_U136 (.ZN( u0_u1_n571 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n764 ) , .A( u0_u1_n782 ) );
  AOI21_X1 u0_u1_U137 (.ZN( u0_u1_n500 ) , .A( u0_u1_n726 ) , .B2( u0_u1_n764 ) , .B1( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U138 (.ZN( u0_u1_n685 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U139 (.ZN( u0_u1_n713 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n765 ) );
  NOR4_X1 u0_u1_U14 (.ZN( u0_u1_n458 ) , .A2( u0_u1_n519 ) , .A1( u0_u1_n545 ) , .A3( u0_u1_n581 ) , .A4( u0_u1_n617 ) );
  INV_X1 u0_u1_U140 (.A( u0_u1_n805 ) , .ZN( u0_u1_n844 ) );
  AOI21_X1 u0_u1_U141 (.ZN( u0_u1_n517 ) , .A( u0_u1_n731 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U142 (.B1( u0_u1_n627 ) , .ZN( u0_u1_n629 ) , .A( u0_u1_n765 ) , .B2( u0_u1_n816 ) );
  INV_X1 u0_u1_U143 (.A( u0_u1_n792 ) , .ZN( u0_u1_n834 ) );
  NOR2_X1 u0_u1_U144 (.ZN( u0_u1_n616 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U145 (.ZN( u0_u1_n561 ) , .A2( u0_u1_n793 ) , .A1( u0_u1_n805 ) );
  NAND2_X1 u0_u1_U146 (.A1( u0_u1_n701 ) , .A2( u0_u1_n731 ) , .ZN( u0_u1_n784 ) );
  INV_X1 u0_u1_U147 (.A( u0_u1_n749 ) , .ZN( u0_u1_n836 ) );
  INV_X1 u0_u1_U148 (.A( u0_u1_n752 ) , .ZN( u0_u1_n843 ) );
  NOR2_X1 u0_u1_U149 (.ZN( u0_u1_n570 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n764 ) );
  NOR4_X1 u0_u1_U15 (.ZN( u0_u1_n487 ) , .A2( u0_u1_n535 ) , .A1( u0_u1_n560 ) , .A3( u0_u1_n633 ) , .A4( u0_u1_n720 ) );
  INV_X1 u0_u1_U150 (.A( u0_u1_n730 ) , .ZN( u0_u1_n853 ) );
  AOI21_X1 u0_u1_U151 (.ZN( u0_u1_n566 ) , .B1( u0_u1_n726 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U152 (.B1( u0_u1_n688 ) , .ZN( u0_u1_n689 ) , .A( u0_u1_n730 ) , .B2( u0_u1_n763 ) );
  INV_X1 u0_u1_U153 (.A( u0_u1_n731 ) , .ZN( u0_u1_n869 ) );
  AOI211_X1 u0_u1_U154 (.C2( u0_u1_n440 ) , .B( u0_u1_n625 ) , .A( u0_u1_n626 ) , .ZN( u0_u1_n637 ) , .C1( u0_u1_n864 ) );
  NOR4_X1 u0_u1_U155 (.A4( u0_u1_n631 ) , .A3( u0_u1_n632 ) , .A2( u0_u1_n633 ) , .A1( u0_u1_n634 ) , .ZN( u0_u1_n635 ) );
  NOR4_X1 u0_u1_U156 (.A4( u0_u1_n628 ) , .A3( u0_u1_n629 ) , .A2( u0_u1_n630 ) , .ZN( u0_u1_n636 ) , .A1( u0_u1_n666 ) );
  AOI21_X1 u0_u1_U157 (.ZN( u0_u1_n542 ) , .A( u0_u1_n765 ) , .B2( u0_u1_n781 ) , .B1( u0_u1_n819 ) );
  OAI21_X1 u0_u1_U158 (.A( u0_u1_n700 ) , .ZN( u0_u1_n704 ) , .B2( u0_u1_n752 ) , .B1( u0_u1_n806 ) );
  OAI21_X1 u0_u1_U159 (.ZN( u0_u1_n700 ) , .B2( u0_u1_n835 ) , .B1( u0_u1_n839 ) , .A( u0_u1_n861 ) );
  NOR4_X1 u0_u1_U16 (.A4( u0_u1_n447 ) , .A3( u0_u1_n448 ) , .A2( u0_u1_n518 ) , .A1( u0_u1_n543 ) , .ZN( u0_u1_n708 ) );
  INV_X1 u0_u1_U160 (.A( u0_u1_n765 ) , .ZN( u0_u1_n867 ) );
  NOR2_X1 u0_u1_U161 (.ZN( u0_u1_n528 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n752 ) );
  AOI21_X1 u0_u1_U162 (.ZN( u0_u1_n445 ) , .B1( u0_u1_n791 ) , .B2( u0_u1_n793 ) , .A( u0_u1_n816 ) );
  NAND4_X1 u0_u1_U163 (.A4( u0_u1_n495 ) , .A3( u0_u1_n496 ) , .A1( u0_u1_n497 ) , .ZN( u0_u1_n804 ) , .A2( u0_u1_n868 ) );
  AOI221_X1 u0_u1_U164 (.B2( u0_u1_n440 ) , .A( u0_u1_n491 ) , .ZN( u0_u1_n496 ) , .C2( u0_u1_n842 ) , .C1( u0_u1_n852 ) , .B1( u0_u1_n861 ) );
  NOR4_X1 u0_u1_U165 (.A3( u0_u1_n439 ) , .A2( u0_u1_n493 ) , .A1( u0_u1_n494 ) , .ZN( u0_u1_n495 ) , .A4( u0_u1_n614 ) );
  INV_X1 u0_u1_U166 (.A( u0_u1_n780 ) , .ZN( u0_u1_n868 ) );
  AOI21_X1 u0_u1_U167 (.ZN( u0_u1_n499 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n793 ) , .B1( u0_u1_n806 ) );
  INV_X1 u0_u1_U168 (.A( u0_u1_n782 ) , .ZN( u0_u1_n851 ) );
  NAND2_X1 u0_u1_U169 (.ZN( u0_u1_n716 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n782 ) );
  OR3_X1 u0_u1_U17 (.ZN( u0_u1_n448 ) , .A1( u0_u1_n530 ) , .A3( u0_u1_n579 ) , .A2( u0_u1_n876 ) );
  BUF_X2 u0_u1_U170 (.Z( u0_u1_n41 ) , .A( u0_u1_n699 ) );
  OR4_X1 u0_u1_U171 (.A4( u0_u1_n582 ) , .A3( u0_u1_n583 ) , .A2( u0_u1_n584 ) , .A1( u0_u1_n585 ) , .ZN( u0_u1_n586 ) );
  INV_X1 u0_u1_U172 (.A( u0_u1_n726 ) , .ZN( u0_u1_n857 ) );
  OAI222_X1 u0_u1_U173 (.B2( u0_u1_n710 ) , .ZN( u0_u1_n711 ) , .C2( u0_u1_n726 ) , .B1( u0_u1_n749 ) , .A1( u0_u1_n808 ) , .C1( u0_u1_n816 ) , .A2( u0_u1_n817 ) );
  AOI221_X1 u0_u1_U174 (.A( u0_u1_n766 ) , .ZN( u0_u1_n776 ) , .C2( u0_u1_n812 ) , .B2( u0_u1_n837 ) , .C1( u0_u1_n856 ) , .B1( u0_u1_n867 ) );
  INV_X1 u0_u1_U175 (.A( u0_u1_n763 ) , .ZN( u0_u1_n837 ) );
  OAI221_X1 u0_u1_U176 (.A( u0_u1_n729 ) , .C2( u0_u1_n730 ) , .B2( u0_u1_n731 ) , .B1( u0_u1_n732 ) , .ZN( u0_u1_n739 ) , .C1( u0_u1_n819 ) );
  OAI221_X1 u0_u1_U177 (.C2( u0_u1_n441 ) , .A( u0_u1_n785 ) , .B2( u0_u1_n787 ) , .B1( u0_u1_n788 ) , .ZN( u0_u1_n798 ) , .C1( u0_u1_n815 ) );
  AOI22_X1 u0_u1_U178 (.A2( u0_u1_n784 ) , .ZN( u0_u1_n785 ) , .B2( u0_u1_n833 ) , .A1( u0_u1_n836 ) , .B1( u0_u1_n864 ) );
  OAI221_X1 u0_u1_U179 (.C2( u0_u1_n441 ) , .A( u0_u1_n698 ) , .ZN( u0_u1_n705 ) , .C1( u0_u1_n787 ) , .B1( u0_u1_n788 ) , .B2( u0_u1_n808 ) );
  OR4_X1 u0_u1_U18 (.A4( u0_u1_n444 ) , .A2( u0_u1_n445 ) , .A1( u0_u1_n446 ) , .ZN( u0_u1_n447 ) , .A3( u0_u1_n555 ) );
  AOI22_X1 u0_u1_U180 (.ZN( u0_u1_n698 ) , .A1( u0_u1_n832 ) , .B2( u0_u1_n844 ) , .A2( u0_u1_n866 ) , .B1( u0_u1_n869 ) );
  OAI222_X1 u0_u1_U181 (.B1( u0_u1_n41 ) , .ZN( u0_u1_n619 ) , .C1( u0_u1_n726 ) , .C2( u0_u1_n749 ) , .B2( u0_u1_n788 ) , .A2( u0_u1_n794 ) , .A1( u0_u1_n818 ) );
  NAND2_X1 u0_u1_U182 (.A2( u0_u1_n450 ) , .A1( u0_u1_n466 ) , .ZN( u0_u1_n817 ) );
  NAND2_X1 u0_u1_U183 (.A2( u0_u1_n456 ) , .A1( u0_u1_n474 ) , .ZN( u0_u1_n781 ) );
  NAND2_X1 u0_u1_U184 (.A2( u0_u1_n450 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n731 ) );
  NAND2_X1 u0_u1_U185 (.A1( u0_u1_n455 ) , .A2( u0_u1_n474 ) , .ZN( u0_u1_n787 ) );
  NAND2_X1 u0_u1_U186 (.A1( u0_u1_n455 ) , .A2( u0_u1_n463 ) , .ZN( u0_u1_n746 ) );
  NAND2_X1 u0_u1_U187 (.A1( u0_u1_n453 ) , .A2( u0_u1_n473 ) , .ZN( u0_u1_n818 ) );
  NAND2_X1 u0_u1_U188 (.A2( u0_u1_n455 ) , .A1( u0_u1_n457 ) , .ZN( u0_u1_n808 ) );
  NOR2_X1 u0_u1_U189 (.ZN( u0_u1_n467 ) , .A2( u0_u1_n848 ) , .A1( u0_u1_n849 ) );
  INV_X1 u0_u1_U19 (.A( u0_u1_n615 ) , .ZN( u0_u1_n876 ) );
  NAND2_X1 u0_u1_U190 (.A1( u0_u1_n449 ) , .A2( u0_u1_n450 ) , .ZN( u0_u1_n788 ) );
  NAND2_X1 u0_u1_U191 (.A2( u0_u1_n463 ) , .A1( u0_u1_n464 ) , .ZN( u0_u1_n749 ) );
  NAND2_X1 u0_u1_U192 (.A1( u0_u1_n464 ) , .A2( u0_u1_n474 ) , .ZN( u0_u1_n790 ) );
  NAND2_X1 u0_u1_U193 (.A1( u0_u1_n453 ) , .A2( u0_u1_n464 ) , .ZN( u0_u1_n792 ) );
  AND2_X1 u0_u1_U194 (.ZN( u0_u1_n440 ) , .A1( u0_u1_n456 ) , .A2( u0_u1_n463 ) );
  NOR2_X1 u0_u1_U195 (.A2( u0_n268 ) , .ZN( u0_u1_n462 ) , .A1( u0_u1_n850 ) );
  AOI222_X1 u0_u1_U196 (.B2( u0_u1_n640 ) , .ZN( u0_u1_n646 ) , .B1( u0_u1_n842 ) , .A1( u0_u1_n843 ) , .C2( u0_u1_n847 ) , .C1( u0_u1_n864 ) , .A2( u0_u1_n866 ) );
  NOR4_X1 u0_u1_U197 (.A4( u0_u1_n641 ) , .A3( u0_u1_n642 ) , .A2( u0_u1_n643 ) , .A1( u0_u1_n644 ) , .ZN( u0_u1_n645 ) );
  NOR4_X1 u0_u1_U198 (.A4( u0_u1_n500 ) , .A3( u0_u1_n501 ) , .A2( u0_u1_n502 ) , .ZN( u0_u1_n503 ) , .A1( u0_u1_n529 ) );
  AOI221_X1 u0_u1_U199 (.A( u0_u1_n499 ) , .ZN( u0_u1_n504 ) , .B2( u0_u1_n844 ) , .C1( u0_u1_n847 ) , .C2( u0_u1_n861 ) , .B1( u0_u1_n863 ) );
  NOR4_X1 u0_u1_U20 (.ZN( u0_u1_n622 ) , .A1( u0_u1_n658 ) , .A3( u0_u1_n668 ) , .A4( u0_u1_n684 ) , .A2( u0_u1_n768 ) );
  AOI221_X1 u0_u1_U200 (.A( u0_u1_n783 ) , .ZN( u0_u1_n800 ) , .C2( u0_u1_n838 ) , .B2( u0_u1_n839 ) , .B1( u0_u1_n866 ) , .C1( u0_u1_n867 ) );
  NOR4_X1 u0_u1_U201 (.A4( u0_u1_n795 ) , .A3( u0_u1_n796 ) , .A2( u0_u1_n797 ) , .A1( u0_u1_n798 ) , .ZN( u0_u1_n799 ) );
  NAND4_X1 u0_u1_U202 (.ZN( u0_subword_23 ) , .A4( u0_u1_n824 ) , .A3( u0_u1_n825 ) , .A2( u0_u1_n826 ) , .A1( u0_u1_n827 ) );
  NOR4_X1 u0_u1_U203 (.A4( u0_u1_n820 ) , .A3( u0_u1_n821 ) , .A2( u0_u1_n822 ) , .A1( u0_u1_n823 ) , .ZN( u0_u1_n824 ) );
  NOR4_X1 u0_u1_U204 (.A4( u0_u1_n736 ) , .A3( u0_u1_n737 ) , .A2( u0_u1_n738 ) , .A1( u0_u1_n739 ) , .ZN( u0_u1_n740 ) );
  NOR4_X1 u0_u1_U205 (.A3( u0_u1_n757 ) , .A2( u0_u1_n758 ) , .A1( u0_u1_n759 ) , .ZN( u0_u1_n760 ) , .A4( u0_u1_n870 ) );
  AOI211_X1 u0_u1_U206 (.B( u0_u1_n747 ) , .A( u0_u1_n748 ) , .ZN( u0_u1_n761 ) , .C1( u0_u1_n834 ) , .C2( u0_u1_n854 ) );
  NOR4_X1 u0_u1_U207 (.A4( u0_u1_n702 ) , .A3( u0_u1_n703 ) , .A2( u0_u1_n704 ) , .A1( u0_u1_n705 ) , .ZN( u0_u1_n706 ) );
  AOI211_X1 u0_u1_U208 (.B( u0_u1_n696 ) , .A( u0_u1_n697 ) , .ZN( u0_u1_n707 ) , .C2( u0_u1_n833 ) , .C1( u0_u1_n852 ) );
  NAND4_X1 u0_u1_U209 (.ZN( u0_subword_17 ) , .A4( u0_u1_n597 ) , .A3( u0_u1_n598 ) , .A2( u0_u1_n599 ) , .A1( u0_u1_n600 ) );
  NOR4_X1 u0_u1_U21 (.A4( u0_u1_n611 ) , .A3( u0_u1_n612 ) , .A2( u0_u1_n613 ) , .A1( u0_u1_n614 ) , .ZN( u0_u1_n621 ) );
  NOR4_X1 u0_u1_U210 (.A4( u0_u1_n593 ) , .A3( u0_u1_n594 ) , .A2( u0_u1_n595 ) , .A1( u0_u1_n596 ) , .ZN( u0_u1_n597 ) );
  AOI211_X1 u0_u1_U211 (.B( u0_u1_n591 ) , .A( u0_u1_n592 ) , .ZN( u0_u1_n598 ) , .C2( u0_u1_n813 ) , .C1( u0_u1_n835 ) );
  NAND2_X1 u0_u1_U212 (.A2( u0_u1_n443 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U213 (.ZN( u0_u1_n642 ) , .B2( u0_u1_n749 ) , .A( u0_u1_n794 ) , .B1( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U214 (.ZN( u0_u1_n516 ) , .A( u0_u1_n781 ) , .B2( u0_u1_n794 ) , .B1( u0_u1_n814 ) );
  INV_X1 u0_u1_U215 (.A( u0_u1_n794 ) , .ZN( u0_u1_n852 ) );
  NOR2_X1 u0_u1_U216 (.ZN( u0_u1_n559 ) , .A1( u0_u1_n794 ) , .A2( u0_u1_n816 ) );
  NOR2_X1 u0_u1_U217 (.ZN( u0_u1_n585 ) , .A1( u0_u1_n794 ) , .A2( u0_u1_n819 ) );
  NAND2_X2 u0_u1_U218 (.A1( u0_u1_n453 ) , .A2( u0_u1_n455 ) , .ZN( u0_u1_n764 ) );
  NAND2_X2 u0_u1_U219 (.A1( u0_u1_n453 ) , .A2( u0_u1_n456 ) , .ZN( u0_u1_n816 ) );
  NOR4_X1 u0_u1_U22 (.ZN( u0_u1_n563 ) , .A1( u0_u1_n655 ) , .A3( u0_u1_n663 ) , .A4( u0_u1_n687 ) , .A2( u0_u1_n770 ) );
  NOR2_X1 u0_u1_U220 (.ZN( u0_u1_n453 ) , .A1( u0_u1_n830 ) , .A2( u0_u1_n831 ) );
  NAND2_X1 u0_u1_U221 (.A1( u0_u1_n454 ) , .A2( u0_u1_n467 ) , .ZN( u0_u1_n671 ) );
  NAND2_X1 u0_u1_U222 (.A1( u0_u1_n443 ) , .A2( u0_u1_n462 ) , .ZN( u0_u1_n701 ) );
  NOR2_X1 u0_u1_U223 (.ZN( u0_u1_n455 ) , .A1( u0_u1_n828 ) , .A2( u0_u1_n829 ) );
  AOI211_X1 u0_u1_U224 (.B( u0_u1_n727 ) , .A( u0_u1_n728 ) , .ZN( u0_u1_n741 ) , .C1( u0_u1_n844 ) , .C2( u0_u1_n856 ) );
  NOR2_X1 u0_u1_U225 (.A2( u0_u1_n710 ) , .A1( u0_u1_n764 ) , .ZN( u0_u1_n796 ) );
  NOR2_X1 u0_u1_U226 (.ZN( u0_u1_n519 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n805 ) );
  NOR2_X1 u0_u1_U227 (.ZN( u0_u1_n684 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U228 (.A2( u0_u1_n710 ) , .A1( u0_u1_n752 ) , .ZN( u0_u1_n773 ) );
  NOR2_X1 u0_u1_U229 (.ZN( u0_u1_n522 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n816 ) );
  NOR4_X1 u0_u1_U23 (.ZN( u0_u1_n477 ) , .A1( u0_u1_n533 ) , .A3( u0_u1_n570 ) , .A4( u0_u1_n602 ) , .A2( u0_u1_n644 ) );
  NOR2_X1 u0_u1_U230 (.ZN( u0_u1_n531 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n781 ) );
  INV_X1 u0_u1_U231 (.A( u0_u1_n682 ) , .ZN( u0_u1_n841 ) );
  AOI21_X1 u0_u1_U232 (.ZN( u0_u1_n643 ) , .B1( u0_u1_n682 ) , .A( u0_u1_n793 ) , .B2( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U233 (.B2( u0_u1_n781 ) , .B1( u0_u1_n782 ) , .ZN( u0_u1_n783 ) , .A2( u0_u1_n816 ) , .A1( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U234 (.ZN( u0_u1_n591 ) , .B2( u0_u1_n701 ) , .B1( u0_u1_n817 ) , .A( u0_u1_n819 ) );
  INV_X1 u0_u1_U235 (.A( u0_u1_n817 ) , .ZN( u0_u1_n856 ) );
  NOR2_X1 u0_u1_U236 (.ZN( u0_u1_n669 ) , .A1( u0_u1_n752 ) , .A2( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U237 (.ZN( u0_u1_n541 ) , .B2( u0_u1_n814 ) , .A( u0_u1_n816 ) , .B1( u0_u1_n817 ) );
  AOI21_X1 u0_u1_U238 (.ZN( u0_u1_n452 ) , .B2( u0_u1_n794 ) , .A( u0_u1_n805 ) , .B1( u0_u1_n817 ) );
  NOR2_X1 u0_u1_U239 (.ZN( u0_u1_n472 ) , .A2( u0_u1_n781 ) , .A1( u0_u1_n817 ) );
  NOR4_X1 u0_u1_U24 (.ZN( u0_u1_n483 ) , .A3( u0_u1_n534 ) , .A4( u0_u1_n547 ) , .A2( u0_u1_n569 ) , .A1( u0_u1_n719 ) );
  OAI222_X1 u0_u1_U240 (.A2( u0_u1_n671 ) , .ZN( u0_u1_n676 ) , .B1( u0_u1_n749 ) , .B2( u0_u1_n786 ) , .C2( u0_u1_n790 ) , .C1( u0_u1_n817 ) , .A1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U241 (.ZN( u0_u1_n632 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n817 ) );
  NAND2_X1 u0_u1_U242 (.A1( u0_u1_n443 ) , .A2( u0_u1_n466 ) , .ZN( u0_u1_n710 ) );
  NAND2_X1 u0_u1_U243 (.A2( u0_u1_n463 ) , .A1( u0_u1_n473 ) , .ZN( u0_u1_n699 ) );
  INV_X1 u0_u1_U244 (.ZN( u0_u1_n438 ) , .A( u0_u1_n788 ) );
  INV_X1 u0_u1_U245 (.ZN( u0_u1_n828 ) , .A( w3_8 ) );
  NOR2_X1 u0_u1_U246 (.ZN( u0_u1_n456 ) , .A1( u0_u1_n829 ) , .A2( w3_8 ) );
  NOR2_X1 u0_u1_U247 (.A2( u0_n270 ) , .ZN( u0_u1_n454 ) , .A1( u0_u1_n859 ) );
  OAI21_X1 u0_u1_U248 (.A( u0_u1_n789 ) , .B2( u0_u1_n790 ) , .B1( u0_u1_n791 ) , .ZN( u0_u1_n797 ) );
  AOI21_X1 u0_u1_U249 (.ZN( u0_u1_n641 ) , .B2( u0_u1_n751 ) , .A( u0_u1_n790 ) , .B1( u0_u1_n814 ) );
  INV_X1 u0_u1_U25 (.A( u0_u1_n751 ) , .ZN( u0_u1_n864 ) );
  AOI21_X1 u0_u1_U250 (.A( u0_u1_n735 ) , .ZN( u0_u1_n736 ) , .B2( u0_u1_n782 ) , .B1( u0_u1_n794 ) );
  AOI21_X1 u0_u1_U251 (.B2( u0_u1_n765 ) , .ZN( u0_u1_n766 ) , .A( u0_u1_n790 ) , .B1( u0_u1_n794 ) );
  AOI21_X1 u0_u1_U252 (.ZN( u0_u1_n444 ) , .A( u0_u1_n701 ) , .B1( u0_u1_n735 ) , .B2( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U253 (.ZN( u0_u1_n520 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n790 ) );
  NOR2_X1 u0_u1_U254 (.ZN( u0_u1_n536 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n790 ) );
  NOR2_X1 u0_u1_U255 (.ZN( u0_u1_n644 ) , .A2( u0_u1_n790 ) , .A1( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U256 (.ZN( u0_u1_n583 ) , .A1( u0_u1_n671 ) , .A2( u0_u1_n790 ) );
  INV_X1 u0_u1_U257 (.A( u0_u1_n790 ) , .ZN( u0_u1_n846 ) );
  AOI222_X1 u0_u1_U258 (.ZN( u0_u1_n527 ) , .A1( u0_u1_n836 ) , .B2( u0_u1_n838 ) , .C1( u0_u1_n845 ) , .C2( u0_u1_n851 ) , .A2( u0_u1_n853 ) , .B1( u0_u1_n867 ) );
  NOR3_X1 u0_u1_U259 (.A2( u0_u1_n440 ) , .ZN( u0_u1_n442 ) , .A3( u0_u1_n838 ) , .A1( u0_u1_n847 ) );
  NOR4_X1 u0_u1_U26 (.A1( u0_u1_n533 ) , .ZN( u0_u1_n538 ) , .A2( u0_u1_n656 ) , .A4( u0_u1_n670 ) , .A3( u0_u1_n767 ) );
  NAND2_X1 u0_u1_U260 (.ZN( u0_u1_n615 ) , .A2( u0_u1_n838 ) , .A1( u0_u1_n874 ) );
  AND2_X1 u0_u1_U261 (.ZN( u0_u1_n627 ) , .A1( u0_u1_n732 ) , .A2( u0_u1_n815 ) );
  NAND2_X1 u0_u1_U262 (.A2( u0_u1_n456 ) , .A1( u0_u1_n457 ) , .ZN( u0_u1_n732 ) );
  NOR2_X1 u0_u1_U263 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n439 ) , .A1( u0_u1_n793 ) );
  AOI21_X1 u0_u1_U264 (.ZN( u0_u1_n593 ) , .B2( u0_u1_n765 ) , .A( u0_u1_n787 ) , .B1( u0_u1_n814 ) );
  AND2_X1 u0_u1_U265 (.ZN( u0_u1_n734 ) , .A1( u0_u1_n781 ) , .A2( u0_u1_n787 ) );
  NAND4_X1 u0_u1_U266 (.A4( u0_u1_n550 ) , .A3( u0_u1_n551 ) , .A2( u0_u1_n552 ) , .A1( u0_u1_n553 ) , .ZN( u0_u1_n747 ) );
  NOR2_X1 u0_u1_U267 (.ZN( u0_u1_n666 ) , .A1( u0_u1_n787 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U268 (.ZN( u0_u1_n665 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U269 (.ZN( u0_u1_n510 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n787 ) );
  NOR4_X1 u0_u1_U27 (.A4( u0_u1_n543 ) , .A3( u0_u1_n544 ) , .A2( u0_u1_n545 ) , .ZN( u0_u1_n552 ) , .A1( u0_u1_n690 ) );
  NOR2_X1 u0_u1_U270 (.ZN( u0_u1_n630 ) , .A2( u0_u1_n671 ) , .A1( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U271 (.ZN( u0_u1_n617 ) , .A1( u0_u1_n787 ) , .A2( u0_u1_n817 ) );
  INV_X1 u0_u1_U272 (.A( u0_u1_n787 ) , .ZN( u0_u1_n847 ) );
  NOR2_X1 u0_u1_U273 (.ZN( u0_u1_n545 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n787 ) );
  NOR2_X1 u0_u1_U274 (.ZN( u0_u1_n546 ) , .A2( u0_u1_n787 ) , .A1( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U275 (.A2( u0_u1_n473 ) , .A1( u0_u1_n474 ) , .ZN( u0_u1_n819 ) );
  AOI222_X1 u0_u1_U276 (.C2( u0_u1_n811 ) , .B2( u0_u1_n812 ) , .A2( u0_u1_n813 ) , .ZN( u0_u1_n825 ) , .C1( u0_u1_n834 ) , .A1( u0_u1_n840 ) , .B1( u0_u1_n854 ) );
  AOI22_X1 u0_u1_U277 (.ZN( u0_u1_n729 ) , .B1( u0_u1_n834 ) , .A2( u0_u1_n839 ) , .A1( u0_u1_n864 ) , .B2( u0_u1_n867 ) );
  AOI222_X1 u0_u1_U278 (.ZN( u0_u1_n471 ) , .B1( u0_u1_n834 ) , .A1( u0_u1_n840 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n852 ) , .A2( u0_u1_n856 ) , .B2( u0_u1_n866 ) );
  NOR2_X1 u0_u1_U279 (.ZN( u0_u1_n688 ) , .A1( u0_u1_n833 ) , .A2( u0_u1_n834 ) );
  NOR2_X1 u0_u1_U28 (.ZN( u0_u1_n544 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U280 (.ZN( u0_u1_n735 ) , .A2( u0_u1_n834 ) , .A1( u0_u1_n846 ) );
  NAND4_X1 u0_u1_U281 (.A4( u0_u1_n537 ) , .A3( u0_u1_n538 ) , .A2( u0_u1_n539 ) , .A1( u0_u1_n540 ) , .ZN( u0_u1_n624 ) );
  NAND2_X2 u0_u1_U282 (.A1( u0_u1_n451 ) , .A2( u0_u1_n462 ) , .ZN( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U283 (.A2( u0_u1_n466 ) , .A1( u0_u1_n467 ) , .ZN( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U284 (.ZN( u0_u1_n631 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n787 ) );
  NAND2_X2 u0_u1_U285 (.A2( u0_u1_n450 ) , .A1( u0_u1_n462 ) , .ZN( u0_u1_n730 ) );
  NOR2_X1 u0_u1_U286 (.A2( u0_n274 ) , .ZN( u0_u1_n451 ) , .A1( u0_u1_n849 ) );
  NOR2_X1 u0_u1_U287 (.A1( u0_n272 ) , .A2( u0_n274 ) , .ZN( u0_u1_n443 ) );
  OAI22_X1 u0_u1_U288 (.ZN( u0_u1_n697 ) , .A2( u0_u1_n732 ) , .A1( u0_u1_n782 ) , .B1( u0_u1_n793 ) , .B2( u0_u1_n819 ) );
  AOI21_X1 u0_u1_U289 (.ZN( u0_u1_n512 ) , .B2( u0_u1_n671 ) , .A( u0_u1_n732 ) , .B1( u0_u1_n817 ) );
  NAND4_X1 u0_u1_U29 (.A4( u0_u1_n605 ) , .A3( u0_u1_n606 ) , .A2( u0_u1_n607 ) , .A1( u0_u1_n608 ) , .ZN( u0_u1_n724 ) );
  OAI22_X1 u0_u1_U290 (.ZN( u0_u1_n491 ) , .A1( u0_u1_n726 ) , .B2( u0_u1_n730 ) , .B1( u0_u1_n732 ) , .A2( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U291 (.ZN( u0_u1_n581 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n732 ) );
  NOR2_X1 u0_u1_U292 (.ZN( u0_u1_n535 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n732 ) );
  INV_X1 u0_u1_U293 (.A( u0_u1_n732 ) , .ZN( u0_u1_n840 ) );
  AOI211_X1 u0_u1_U294 (.A( u0_u1_n498 ) , .ZN( u0_u1_n505 ) , .B( u0_u1_n804 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n852 ) );
  OAI21_X1 u0_u1_U295 (.ZN( u0_u1_n789 ) , .A( u0_u1_n840 ) , .B1( u0_u1_n864 ) , .B2( u0_u1_n874 ) );
  AOI222_X1 u0_u1_U296 (.ZN( u0_u1_n662 ) , .A2( u0_u1_n840 ) , .B1( u0_u1_n842 ) , .C2( u0_u1_n846 ) , .A1( u0_u1_n861 ) , .C1( u0_u1_n864 ) , .B2( u0_u1_n871 ) );
  AOI211_X1 u0_u1_U297 (.B( u0_u1_n541 ) , .A( u0_u1_n542 ) , .ZN( u0_u1_n553 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n852 ) );
  NOR2_X1 u0_u1_U298 (.ZN( u0_u1_n682 ) , .A2( u0_u1_n836 ) , .A1( u0_u1_n840 ) );
  NAND4_X1 u0_u1_U299 (.ZN( u0_subword_16 ) , .A4( u0_u1_n503 ) , .A3( u0_u1_n504 ) , .A2( u0_u1_n505 ) , .A1( u0_u1_n506 ) );
  NAND2_X1 u0_u1_U3 (.A1( u0_u1_n451 ) , .A2( u0_u1_n466 ) , .ZN( u0_u1_n726 ) );
  NOR4_X1 u0_u1_U30 (.A3( u0_u1_n602 ) , .A2( u0_u1_n603 ) , .A1( u0_u1_n604 ) , .ZN( u0_u1_n605 ) , .A4( u0_u1_n657 ) );
  AOI21_X1 u0_u1_U300 (.A( u0_u1_n792 ) , .B2( u0_u1_n793 ) , .B1( u0_u1_n794 ) , .ZN( u0_u1_n795 ) );
  AOI21_X1 u0_u1_U301 (.ZN( u0_u1_n628 ) , .B2( u0_u1_n671 ) , .A( u0_u1_n792 ) , .B1( u0_u1_n793 ) );
  NOR2_X1 u0_u1_U302 (.ZN( u0_u1_n657 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n817 ) );
  NOR2_X1 u0_u1_U303 (.ZN( u0_u1_n714 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n792 ) );
  NOR2_X1 u0_u1_U304 (.ZN( u0_u1_n523 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U305 (.ZN( u0_u1_n663 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n792 ) );
  NOR2_X1 u0_u1_U306 (.ZN( u0_u1_n670 ) , .A2( u0_u1_n710 ) , .A1( u0_u1_n792 ) );
  NOR3_X1 u0_u1_U307 (.A3( u0_u1_n743 ) , .A2( u0_u1_n744 ) , .A1( u0_u1_n745 ) , .ZN( u0_u1_n762 ) );
  NAND2_X2 u0_u1_U308 (.A2( u0_u1_n451 ) , .A1( u0_u1_n454 ) , .ZN( u0_u1_n765 ) );
  OAI22_X1 u0_u1_U309 (.ZN( u0_u1_n639 ) , .A1( u0_u1_n701 ) , .B2( u0_u1_n730 ) , .A2( u0_u1_n764 ) , .B1( u0_u1_n818 ) );
  NOR3_X1 u0_u1_U31 (.A1( u0_u1_n601 ) , .ZN( u0_u1_n606 ) , .A3( u0_u1_n665 ) , .A2( u0_u1_n772 ) );
  AOI21_X1 u0_u1_U310 (.ZN( u0_u1_n501 ) , .B1( u0_u1_n682 ) , .A( u0_u1_n814 ) , .B2( u0_u1_n818 ) );
  OAI22_X1 u0_u1_U311 (.A1( u0_u1_n726 ) , .ZN( u0_u1_n728 ) , .B2( u0_u1_n752 ) , .B1( u0_u1_n814 ) , .A2( u0_u1_n818 ) );
  AOI21_X1 u0_u1_U312 (.A( u0_u1_n817 ) , .B2( u0_u1_n818 ) , .B1( u0_u1_n819 ) , .ZN( u0_u1_n820 ) );
  OAI22_X1 u0_u1_U313 (.ZN( u0_u1_n626 ) , .B1( u0_u1_n671 ) , .B2( u0_u1_n749 ) , .A1( u0_u1_n817 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U314 (.ZN( u0_u1_n601 ) , .A2( u0_u1_n793 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U315 (.ZN( u0_u1_n533 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U316 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n690 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U317 (.ZN( u0_u1_n521 ) , .A2( u0_u1_n701 ) , .A1( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U318 (.ZN( u0_u1_n560 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U319 (.ZN( u0_u1_n687 ) , .A1( u0_u1_n731 ) , .A2( u0_u1_n818 ) );
  NOR3_X1 u0_u1_U32 (.ZN( u0_u1_n551 ) , .A2( u0_u1_n653 ) , .A1( u0_u1_n669 ) , .A3( u0_u1_n773 ) );
  INV_X1 u0_u1_U320 (.A( u0_u1_n818 ) , .ZN( u0_u1_n833 ) );
  BUF_X2 u0_u1_U321 (.Z( u0_u1_n441 ) , .A( u0_u1_n786 ) );
  NAND2_X1 u0_u1_U322 (.A2( u0_u1_n443 ) , .A1( u0_u1_n449 ) , .ZN( u0_u1_n786 ) );
  AOI222_X1 u0_u1_U323 (.ZN( u0_u1_n777 ) , .A1( u0_u1_n832 ) , .C1( u0_u1_n836 ) , .B2( u0_u1_n842 ) , .A2( u0_u1_n851 ) , .B1( u0_u1_n862 ) , .C2( u0_u1_n874 ) );
  INV_X1 u0_u1_U324 (.A( u0_n268 ) , .ZN( u0_u1_n859 ) );
  INV_X1 u0_u1_U325 (.A( u0_n274 ) , .ZN( u0_u1_n848 ) );
  INV_X1 u0_u1_U326 (.A( u0_u1_n786 ) , .ZN( u0_u1_n862 ) );
  OAI22_X1 u0_u1_U327 (.B2( u0_u1_n752 ) , .B1( u0_u1_n753 ) , .A1( u0_u1_n754 ) , .ZN( u0_u1_n758 ) , .A2( u0_u1_n808 ) );
  OAI222_X1 u0_u1_U328 (.ZN( u0_u1_n507 ) , .C2( u0_u1_n627 ) , .B2( u0_u1_n649 ) , .B1( u0_u1_n749 ) , .A2( u0_u1_n750 ) , .C1( u0_u1_n807 ) , .A1( u0_u1_n808 ) );
  AOI21_X1 u0_u1_U329 (.ZN( u0_u1_n691 ) , .B2( u0_u1_n751 ) , .B1( u0_u1_n765 ) , .A( u0_u1_n808 ) );
  NOR4_X1 u0_u1_U33 (.A4( u0_u1_n546 ) , .A3( u0_u1_n547 ) , .A2( u0_u1_n548 ) , .A1( u0_u1_n549 ) , .ZN( u0_u1_n550 ) );
  NAND2_X1 u0_u1_U330 (.A2( u0_u1_n764 ) , .A1( u0_u1_n808 ) , .ZN( u0_u1_n812 ) );
  NOR2_X1 u0_u1_U331 (.ZN( u0_u1_n572 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n808 ) );
  AOI21_X1 u0_u1_U332 (.ZN( u0_u1_n479 ) , .A( u0_u1_n671 ) , .B1( u0_u1_n752 ) , .B2( u0_u1_n808 ) );
  OAI22_X1 u0_u1_U333 (.ZN( u0_u1_n485 ) , .A1( u0_u1_n710 ) , .B2( u0_u1_n787 ) , .A2( u0_u1_n808 ) , .B1( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U334 (.ZN( u0_u1_n613 ) , .A2( u0_u1_n782 ) , .A1( u0_u1_n808 ) );
  INV_X1 u0_u1_U335 (.A( u0_u1_n808 ) , .ZN( u0_u1_n842 ) );
  NAND2_X1 u0_u1_U336 (.ZN( u0_u1_n673 ) , .A1( u0_u1_n808 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U337 (.ZN( u0_u1_n464 ) , .A2( w3_8 ) , .A1( w3_9 ) );
  NOR2_X1 u0_u1_U338 (.ZN( u0_u1_n473 ) , .A1( u0_u1_n828 ) , .A2( w3_9 ) );
  INV_X1 u0_u1_U339 (.ZN( u0_u1_n829 ) , .A( w3_9 ) );
  NOR2_X1 u0_u1_U34 (.ZN( u0_u1_n806 ) , .A1( u0_u1_n855 ) , .A2( u0_u1_n862 ) );
  NAND2_X2 u0_u1_U340 (.A1( u0_u1_n457 ) , .A2( u0_u1_n464 ) , .ZN( u0_u1_n752 ) );
  NOR2_X1 u0_u1_U341 (.ZN( u0_u1_n463 ) , .A1( u0_u1_n831 ) , .A2( w3_10 ) );
  INV_X1 u0_u1_U342 (.ZN( u0_u1_n830 ) , .A( w3_10 ) );
  AOI211_X1 u0_u1_U343 (.A( u0_u1_n590 ) , .ZN( u0_u1_n599 ) , .B( u0_u1_n623 ) , .C1( u0_u1_n846 ) , .C2( u0_u1_n856 ) );
  NOR3_X1 u0_u1_U344 (.A3( u0_u1_n623 ) , .A2( u0_u1_n624 ) , .ZN( u0_u1_n638 ) , .A1( u0_u1_n727 ) );
  AOI211_X1 u0_u1_U345 (.B( u0_u1_n479 ) , .A( u0_u1_n480 ) , .ZN( u0_u1_n484 ) , .C2( u0_u1_n835 ) , .C1( u0_u1_n862 ) );
  AOI222_X1 u0_u1_U346 (.ZN( u0_u1_n608 ) , .A1( u0_u1_n832 ) , .C2( u0_u1_n838 ) , .B1( u0_u1_n843 ) , .A2( u0_u1_n857 ) , .B2( u0_u1_n862 ) , .C1( u0_u1_n869 ) );
  AOI21_X1 u0_u1_U347 (.ZN( u0_u1_n595 ) , .B1( u0_u1_n752 ) , .A( u0_u1_n794 ) , .B2( u0_u1_n815 ) );
  AOI21_X1 u0_u1_U348 (.A( u0_u1_n814 ) , .B2( u0_u1_n815 ) , .B1( u0_u1_n816 ) , .ZN( u0_u1_n821 ) );
  AOI21_X1 u0_u1_U349 (.ZN( u0_u1_n651 ) , .B1( u0_u1_n731 ) , .B2( u0_u1_n765 ) , .A( u0_u1_n815 ) );
  NAND4_X1 u0_u1_U35 (.A4( u0_u1_n659 ) , .A3( u0_u1_n660 ) , .A2( u0_u1_n661 ) , .A1( u0_u1_n662 ) , .ZN( u0_u1_n802 ) );
  NOR4_X1 u0_u1_U350 (.A4( u0_u1_n616 ) , .A3( u0_u1_n617 ) , .A2( u0_u1_n618 ) , .A1( u0_u1_n619 ) , .ZN( u0_u1_n620 ) );
  NOR2_X1 u0_u1_U351 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n768 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U352 (.A2( u0_u1_n815 ) , .A1( u0_u1_n817 ) , .ZN( u0_u1_n823 ) );
  NOR2_X1 u0_u1_U353 (.ZN( u0_u1_n580 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U354 (.ZN( u0_u1_n667 ) , .A1( u0_u1_n782 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U355 (.ZN( u0_u1_n686 ) , .A1( u0_u1_n793 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U356 (.A1( u0_u1_n701 ) , .ZN( u0_u1_n770 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U357 (.ZN( u0_u1_n656 ) , .A1( u0_u1_n730 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U358 (.ZN( u0_u1_n633 ) , .A1( u0_u1_n726 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U359 (.ZN( u0_u1_n457 ) , .A1( u0_u1_n830 ) , .A2( w3_11 ) );
  NOR3_X1 u0_u1_U36 (.A3( u0_u1_n650 ) , .A2( u0_u1_n651 ) , .A1( u0_u1_n652 ) , .ZN( u0_u1_n661 ) );
  NOR2_X1 u0_u1_U360 (.ZN( u0_u1_n474 ) , .A2( w3_10 ) , .A1( w3_11 ) );
  INV_X1 u0_u1_U361 (.ZN( u0_u1_n831 ) , .A( w3_11 ) );
  INV_X1 u0_u1_U362 (.A( u0_n270 ) , .ZN( u0_u1_n850 ) );
  NOR2_X1 u0_u1_U363 (.A1( u0_n268 ) , .A2( u0_n270 ) , .ZN( u0_u1_n466 ) );
  NOR2_X1 u0_u1_U364 (.ZN( u0_u1_n449 ) , .A2( u0_u1_n850 ) , .A1( u0_u1_n859 ) );
  INV_X1 u0_u1_U365 (.A( u0_n272 ) , .ZN( u0_u1_n849 ) );
  NOR2_X1 u0_u1_U366 (.A2( u0_n272 ) , .ZN( u0_u1_n450 ) , .A1( u0_u1_n848 ) );
  NOR2_X1 u0_u1_U367 (.A2( u0_u1_n438 ) , .ZN( u0_u1_n750 ) , .A1( u0_u1_n862 ) );
  NOR4_X1 u0_u1_U368 (.A4( u0_u1_n778 ) , .A3( u0_u1_n779 ) , .A1( u0_u1_n780 ) , .ZN( u0_u1_n801 ) , .A2( u0_u1_n803 ) );
  NAND4_X1 u0_u1_U369 (.A4( u0_u1_n693 ) , .A3( u0_u1_n694 ) , .A1( u0_u1_n695 ) , .ZN( u0_u1_n778 ) , .A2( u0_u1_n873 ) );
  NOR3_X1 u0_u1_U37 (.A3( u0_u1_n653 ) , .A2( u0_u1_n654 ) , .A1( u0_u1_n655 ) , .ZN( u0_u1_n660 ) );
  INV_X1 u0_u1_U370 (.A( u0_u1_n41 ) , .ZN( u0_u1_n839 ) );
  NOR2_X1 u0_u1_U371 (.A1( u0_u1_n41 ) , .ZN( u0_u1_n772 ) , .A2( u0_u1_n817 ) );
  NAND2_X2 u0_u1_U372 (.A1( u0_u1_n457 ) , .A2( u0_u1_n473 ) , .ZN( u0_u1_n805 ) );
  AOI21_X1 u0_u1_U373 (.B2( u0_u1_n41 ) , .ZN( u0_u1_n573 ) , .B1( u0_u1_n808 ) , .A( u0_u1_n814 ) );
  NOR2_X1 u0_u1_U374 (.A2( u0_u1_n41 ) , .A1( u0_u1_n782 ) , .ZN( u0_u1_n822 ) );
  NOR2_X1 u0_u1_U375 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n634 ) , .A1( u0_u1_n726 ) );
  NOR2_X1 u0_u1_U376 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n568 ) , .A1( u0_u1_n765 ) );
  NOR2_X1 u0_u1_U377 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n664 ) , .A1( u0_u1_n731 ) );
  AOI21_X1 u0_u1_U378 (.B2( u0_u1_n41 ) , .ZN( u0_u1_n480 ) , .A( u0_u1_n751 ) , .B1( u0_u1_n781 ) );
  NOR2_X1 u0_u1_U379 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n718 ) , .A1( u0_u1_n794 ) );
  NOR3_X1 u0_u1_U38 (.A3( u0_u1_n656 ) , .A2( u0_u1_n657 ) , .A1( u0_u1_n658 ) , .ZN( u0_u1_n659 ) );
  NOR2_X1 u0_u1_U380 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n596 ) , .A1( u0_u1_n730 ) );
  NOR2_X1 u0_u1_U381 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n543 ) , .A1( u0_u1_n701 ) );
  NOR2_X1 u0_u1_U382 (.ZN( u0_u1_n582 ) , .A2( u0_u1_n699 ) , .A1( u0_u1_n793 ) );
  NAND4_X1 u0_u1_U383 (.ZN( u0_subword_18 ) , .A4( u0_u1_n645 ) , .A3( u0_u1_n646 ) , .A2( u0_u1_n647 ) , .A1( u0_u1_n648 ) );
  OAI21_X1 u0_u1_U384 (.A( u0_u1_n733 ) , .B1( u0_u1_n734 ) , .ZN( u0_u1_n738 ) , .B2( u0_u1_n807 ) );
  OAI222_X1 u0_u1_U385 (.B2( u0_u1_n749 ) , .B1( u0_u1_n750 ) , .A2( u0_u1_n751 ) , .ZN( u0_u1_n759 ) , .C2( u0_u1_n807 ) , .C1( u0_u1_n816 ) , .A1( u0_u1_n819 ) );
  OAI22_X1 u0_u1_U386 (.B2( u0_u1_n805 ) , .B1( u0_u1_n806 ) , .A2( u0_u1_n807 ) , .A1( u0_u1_n808 ) , .ZN( u0_u1_n810 ) );
  AOI21_X1 u0_u1_U387 (.ZN( u0_u1_n652 ) , .A( u0_u1_n781 ) , .B1( u0_u1_n794 ) , .B2( u0_u1_n807 ) );
  INV_X1 u0_u1_U388 (.A( u0_u1_n807 ) , .ZN( u0_u1_n861 ) );
  NOR2_X1 u0_u1_U389 (.ZN( u0_u1_n737 ) , .A2( u0_u1_n805 ) , .A1( u0_u1_n807 ) );
  OAI21_X1 u0_u1_U39 (.ZN( u0_u1_n733 ) , .A( u0_u1_n835 ) , .B2( u0_u1_n853 ) , .B1( u0_u1_n874 ) );
  NOR2_X1 u0_u1_U390 (.ZN( u0_u1_n486 ) , .A1( u0_u1_n790 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U391 (.ZN( u0_u1_n569 ) , .A1( u0_u1_n749 ) , .A2( u0_u1_n807 ) );
  AOI21_X1 u0_u1_U392 (.A( u0_u1_n41 ) , .ZN( u0_u1_n554 ) , .B1( u0_u1_n671 ) , .B2( u0_u1_n807 ) );
  NAND2_X1 u0_u1_U393 (.ZN( u0_u1_n755 ) , .A1( u0_u1_n765 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U394 (.ZN( u0_u1_n717 ) , .A1( u0_u1_n807 ) , .A2( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U395 (.ZN( u0_u1_n558 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U396 (.ZN( u0_u1_n672 ) , .A1( u0_u1_n792 ) , .A2( u0_u1_n807 ) );
  NAND4_X1 u0_u1_U397 (.ZN( u0_subword_19 ) , .A4( u0_u1_n706 ) , .A3( u0_u1_n707 ) , .A2( u0_u1_n708 ) , .A1( u0_u1_n709 ) );
  INV_X1 u0_u1_U398 (.A( u0_u1_n708 ) , .ZN( u0_u1_n877 ) );
  OAI22_X1 u0_u1_U399 (.B2( u0_u1_n746 ) , .ZN( u0_u1_n748 ) , .A2( u0_u1_n764 ) , .B1( u0_u1_n782 ) , .A1( u0_u1_n794 ) );
  NAND2_X1 u0_u1_U4 (.A2( u0_u1_n462 ) , .A1( u0_u1_n467 ) , .ZN( u0_u1_n782 ) );
  INV_X1 u0_u1_U40 (.A( u0_u1_n681 ) , .ZN( u0_u1_n873 ) );
  OAI22_X1 u0_u1_U400 (.ZN( u0_u1_n498 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n782 ) , .B1( u0_u1_n793 ) , .B2( u0_u1_n808 ) );
  NOR2_X1 u0_u1_U401 (.ZN( u0_u1_n518 ) , .A1( u0_u1_n710 ) , .A2( u0_u1_n746 ) );
  OAI22_X1 u0_u1_U402 (.ZN( u0_u1_n712 ) , .A2( u0_u1_n730 ) , .B2( u0_u1_n731 ) , .A1( u0_u1_n746 ) , .B1( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U403 (.A2( u0_u1_n746 ) , .ZN( u0_u1_n771 ) , .A1( u0_u1_n814 ) );
  OAI22_X1 u0_u1_U404 (.B1( u0_u1_n442 ) , .ZN( u0_u1_n446 ) , .A2( u0_u1_n730 ) , .A1( u0_u1_n746 ) , .B2( u0_u1_n751 ) );
  NOR2_X1 u0_u1_U405 (.ZN( u0_u1_n549 ) , .A1( u0_u1_n701 ) , .A2( u0_u1_n746 ) );
  NOR2_X1 u0_u1_U406 (.ZN( u0_u1_n532 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n794 ) );
  NOR2_X1 u0_u1_U407 (.A2( u0_u1_n746 ) , .ZN( u0_u1_n757 ) , .A1( u0_u1_n807 ) );
  NOR2_X1 u0_u1_U408 (.A1( u0_u1_n671 ) , .ZN( u0_u1_n675 ) , .A2( u0_u1_n746 ) );
  NOR2_X1 u0_u1_U409 (.ZN( u0_u1_n720 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n746 ) );
  NOR4_X1 u0_u1_U41 (.A4( u0_u1_n689 ) , .A3( u0_u1_n690 ) , .A2( u0_u1_n691 ) , .A1( u0_u1_n692 ) , .ZN( u0_u1_n693 ) );
  NOR2_X1 u0_u1_U410 (.ZN( u0_u1_n584 ) , .A1( u0_u1_n746 ) , .A2( u0_u1_n817 ) );
  INV_X1 u0_u1_U411 (.A( u0_u1_n746 ) , .ZN( u0_u1_n838 ) );
  AOI221_X1 u0_u1_U412 (.A( u0_u1_n578 ) , .ZN( u0_u1_n589 ) , .B2( u0_u1_n833 ) , .C2( u0_u1_n844 ) , .B1( u0_u1_n855 ) , .C1( u0_u1_n862 ) );
  AOI21_X1 u0_u1_U413 (.ZN( u0_u1_n578 ) , .B2( u0_u1_n726 ) , .B1( u0_u1_n750 ) , .A( u0_u1_n787 ) );
  AOI211_X1 u0_u1_U414 (.A( u0_u1_n639 ) , .ZN( u0_u1_n647 ) , .B( u0_u1_n745 ) , .C2( u0_u1_n840 ) , .C1( u0_u1_n855 ) );
  NAND4_X1 u0_u1_U415 (.A4( u0_u1_n635 ) , .A3( u0_u1_n636 ) , .A2( u0_u1_n637 ) , .A1( u0_u1_n638 ) , .ZN( u0_u1_n745 ) );
  OAI22_X1 u0_u1_U416 (.B1( u0_u1_n441 ) , .ZN( u0_u1_n590 ) , .A2( u0_u1_n749 ) , .B2( u0_u1_n764 ) , .A1( u0_u1_n765 ) );
  NAND2_X1 u0_u1_U417 (.A2( u0_u1_n441 ) , .A1( u0_u1_n731 ) , .ZN( u0_u1_n813 ) );
  AOI21_X1 u0_u1_U418 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n594 ) , .B1( u0_u1_n730 ) , .A( u0_u1_n792 ) );
  AOI21_X1 u0_u1_U419 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n650 ) , .A( u0_u1_n764 ) , .B1( u0_u1_n794 ) );
  AOI221_X1 u0_u1_U42 (.A( u0_u1_n683 ) , .ZN( u0_u1_n694 ) , .B2( u0_u1_n841 ) , .C1( u0_u1_n843 ) , .C2( u0_u1_n863 ) , .B1( u0_u1_n866 ) );
  AOI21_X1 u0_u1_U420 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n625 ) , .B1( u0_u1_n701 ) , .A( u0_u1_n781 ) );
  OAI22_X1 u0_u1_U421 (.B2( u0_u1_n441 ) , .ZN( u0_u1_n683 ) , .A1( u0_u1_n701 ) , .A2( u0_u1_n732 ) , .B1( u0_u1_n819 ) );
  NOR2_X1 u0_u1_U422 (.ZN( u0_u1_n653 ) , .A1( u0_u1_n786 ) , .A2( u0_u1_n790 ) );
  OAI21_X1 u0_u1_U423 (.B2( u0_u1_n441 ) , .A( u0_u1_n615 ) , .ZN( u0_u1_n618 ) , .B1( u0_u1_n627 ) );
  NOR2_X1 u0_u1_U424 (.A1( u0_u1_n441 ) , .ZN( u0_u1_n612 ) , .A2( u0_u1_n818 ) );
  NOR2_X1 u0_u1_U425 (.ZN( u0_u1_n555 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n786 ) );
  NOR2_X1 u0_u1_U426 (.A2( u0_u1_n41 ) , .ZN( u0_u1_n602 ) , .A1( u0_u1_n786 ) );
  AOI21_X1 u0_u1_U427 (.A( u0_u1_n41 ) , .ZN( u0_u1_n502 ) , .B1( u0_u1_n710 ) , .B2( u0_u1_n788 ) );
  OAI22_X1 u0_u1_U428 (.ZN( u0_u1_n592 ) , .B1( u0_u1_n732 ) , .B2( u0_u1_n751 ) , .A2( u0_u1_n788 ) , .A1( u0_u1_n805 ) );
  AOI222_X1 u0_u1_U429 (.ZN( u0_u1_n515 ) , .C1( u0_u1_n834 ) , .B2( u0_u1_n838 ) , .A2( u0_u1_n844 ) , .C2( u0_u1_n863 ) , .B1( u0_u1_n864 ) , .A1( u0_u1_n867 ) );
  NOR4_X1 u0_u1_U43 (.A4( u0_u1_n528 ) , .A2( u0_u1_n529 ) , .A1( u0_u1_n530 ) , .ZN( u0_u1_n540 ) , .A3( u0_u1_n703 ) );
  AOI222_X1 u0_u1_U430 (.ZN( u0_u1_n607 ) , .B2( u0_u1_n673 ) , .B1( u0_u1_n755 ) , .C2( u0_u1_n833 ) , .A1( u0_u1_n835 ) , .A2( u0_u1_n863 ) , .C1( u0_u1_n864 ) );
  AOI221_X1 u0_u1_U431 (.A( u0_u1_n485 ) , .ZN( u0_u1_n490 ) , .B1( u0_u1_n833 ) , .C2( u0_u1_n845 ) , .C1( u0_u1_n853 ) , .B2( u0_u1_n863 ) );
  NOR2_X1 u0_u1_U432 (.ZN( u0_u1_n655 ) , .A1( u0_u1_n764 ) , .A2( u0_u1_n788 ) );
  NAND2_X1 u0_u1_U433 (.A2( u0_u1_n751 ) , .A1( u0_u1_n788 ) , .ZN( u0_u1_n811 ) );
  NOR2_X1 u0_u1_U434 (.ZN( u0_u1_n556 ) , .A1( u0_u1_n788 ) , .A2( u0_u1_n815 ) );
  NOR2_X1 u0_u1_U435 (.ZN( u0_u1_n614 ) , .A1( u0_u1_n781 ) , .A2( u0_u1_n788 ) );
  NOR2_X1 u0_u1_U436 (.ZN( u0_u1_n719 ) , .A2( u0_u1_n746 ) , .A1( u0_u1_n788 ) );
  NAND3_X1 u0_u1_U437 (.ZN( u0_subword_22 ) , .A3( u0_u1_n799 ) , .A2( u0_u1_n800 ) , .A1( u0_u1_n801 ) );
  NAND3_X1 u0_u1_U438 (.ZN( u0_subword_21 ) , .A3( u0_u1_n760 ) , .A2( u0_u1_n761 ) , .A1( u0_u1_n762 ) );
  NAND3_X1 u0_u1_U439 (.ZN( u0_subword_20 ) , .A3( u0_u1_n740 ) , .A2( u0_u1_n741 ) , .A1( u0_u1_n742 ) );
  NOR4_X1 u0_u1_U44 (.A4( u0_u1_n534 ) , .A3( u0_u1_n535 ) , .A2( u0_u1_n536 ) , .ZN( u0_u1_n537 ) , .A1( u0_u1_n822 ) );
  NAND3_X1 u0_u1_U440 (.A3( u0_u1_n677 ) , .A2( u0_u1_n678 ) , .A1( u0_u1_n679 ) , .ZN( u0_u1_n809 ) );
  NAND3_X1 u0_u1_U441 (.ZN( u0_u1_n640 ) , .A3( u0_u1_n710 ) , .A2( u0_u1_n726 ) , .A1( u0_u1_n794 ) );
  NAND3_X1 u0_u1_U442 (.A3( u0_u1_n620 ) , .A2( u0_u1_n621 ) , .A1( u0_u1_n622 ) , .ZN( u0_u1_n727 ) );
  NAND3_X1 u0_u1_U443 (.A3( u0_u1_n587 ) , .A2( u0_u1_n588 ) , .A1( u0_u1_n589 ) , .ZN( u0_u1_n623 ) );
  NAND3_X1 u0_u1_U444 (.ZN( u0_u1_n567 ) , .A3( u0_u1_n682 ) , .A2( u0_u1_n752 ) , .A1( u0_u1_n787 ) );
  NAND3_X1 u0_u1_U445 (.A3( u0_u1_n525 ) , .A2( u0_u1_n526 ) , .A1( u0_u1_n527 ) , .ZN( u0_u1_n744 ) );
  NAND3_X1 u0_u1_U446 (.A3( u0_u1_n514 ) , .A1( u0_u1_n515 ) , .ZN( u0_u1_n610 ) , .A2( u0_u1_n872 ) );
  NAND3_X1 u0_u1_U447 (.A3( u0_u1_n469 ) , .A2( u0_u1_n470 ) , .A1( u0_u1_n471 ) , .ZN( u0_u1_n779 ) );
  NOR2_X1 u0_u1_U448 (.ZN( u0_u1_n791 ) , .A2( u0_u1_n863 ) , .A1( u0_u1_n869 ) );
  NOR2_X1 u0_u1_U449 (.ZN( u0_u1_n703 ) , .A2( u0_u1_n788 ) , .A1( u0_u1_n819 ) );
  NOR4_X1 u0_u1_U45 (.A4( u0_u1_n531 ) , .A3( u0_u1_n532 ) , .ZN( u0_u1_n539 ) , .A2( u0_u1_n686 ) , .A1( u0_u1_n796 ) );
  NOR2_X1 u0_u1_U450 (.A1( u0_u1_n732 ) , .ZN( u0_u1_n767 ) , .A2( u0_u1_n788 ) );
  INV_X1 u0_u1_U451 (.A( u0_u1_n788 ) , .ZN( u0_u1_n863 ) );
  NOR3_X1 u0_u1_U46 (.A3( u0_u1_n802 ) , .A2( u0_u1_n803 ) , .A1( u0_u1_n804 ) , .ZN( u0_u1_n827 ) );
  NAND4_X1 u0_u1_U47 (.A4( u0_u1_n481 ) , .A3( u0_u1_n482 ) , .A2( u0_u1_n483 ) , .A1( u0_u1_n484 ) , .ZN( u0_u1_n696 ) );
  NOR3_X1 u0_u1_U48 (.ZN( u0_u1_n482 ) , .A2( u0_u1_n510 ) , .A3( u0_u1_n603 ) , .A1( u0_u1_n612 ) );
  NOR4_X1 u0_u1_U49 (.ZN( u0_u1_n481 ) , .A1( u0_u1_n522 ) , .A4( u0_u1_n559 ) , .A3( u0_u1_n584 ) , .A2( u0_u1_n632 ) );
  NOR3_X1 u0_u1_U5 (.ZN( u0_u1_n600 ) , .A1( u0_u1_n610 ) , .A3( u0_u1_n725 ) , .A2( u0_u1_n744 ) );
  NAND4_X1 u0_u1_U50 (.A4( u0_u1_n774 ) , .A3( u0_u1_n775 ) , .A2( u0_u1_n776 ) , .A1( u0_u1_n777 ) , .ZN( u0_u1_n803 ) );
  NOR3_X1 u0_u1_U51 (.A3( u0_u1_n767 ) , .A2( u0_u1_n768 ) , .A1( u0_u1_n769 ) , .ZN( u0_u1_n775 ) );
  NOR4_X1 u0_u1_U52 (.A4( u0_u1_n770 ) , .A3( u0_u1_n771 ) , .A2( u0_u1_n772 ) , .A1( u0_u1_n773 ) , .ZN( u0_u1_n774 ) );
  NAND4_X1 u0_u1_U53 (.A4( u0_u1_n562 ) , .A3( u0_u1_n563 ) , .A2( u0_u1_n564 ) , .A1( u0_u1_n565 ) , .ZN( u0_u1_n609 ) );
  NOR4_X1 u0_u1_U54 (.A4( u0_u1_n554 ) , .A3( u0_u1_n555 ) , .A2( u0_u1_n556 ) , .A1( u0_u1_n557 ) , .ZN( u0_u1_n564 ) );
  AOI222_X1 u0_u1_U55 (.ZN( u0_u1_n565 ) , .B1( u0_u1_n832 ) , .C1( u0_u1_n842 ) , .A2( u0_u1_n844 ) , .A1( u0_u1_n855 ) , .B2( u0_u1_n864 ) , .C2( u0_u1_n874 ) );
  NOR4_X1 u0_u1_U56 (.A4( u0_u1_n558 ) , .A3( u0_u1_n559 ) , .A2( u0_u1_n560 ) , .A1( u0_u1_n561 ) , .ZN( u0_u1_n562 ) );
  INV_X1 u0_u1_U57 (.A( u0_u1_n507 ) , .ZN( u0_u1_n872 ) );
  NOR4_X1 u0_u1_U58 (.A4( u0_u1_n511 ) , .A2( u0_u1_n512 ) , .A1( u0_u1_n513 ) , .ZN( u0_u1_n514 ) , .A3( u0_u1_n672 ) );
  NOR4_X1 u0_u1_U59 (.A4( u0_u1_n663 ) , .A3( u0_u1_n664 ) , .A2( u0_u1_n665 ) , .A1( u0_u1_n666 ) , .ZN( u0_u1_n679 ) );
  NOR3_X1 u0_u1_U6 (.A2( u0_u1_n609 ) , .A1( u0_u1_n610 ) , .ZN( u0_u1_n648 ) , .A3( u0_u1_n724 ) );
  NOR4_X1 u0_u1_U60 (.A4( u0_u1_n667 ) , .A3( u0_u1_n668 ) , .A2( u0_u1_n669 ) , .A1( u0_u1_n670 ) , .ZN( u0_u1_n678 ) );
  NOR4_X1 u0_u1_U61 (.A3( u0_u1_n675 ) , .A1( u0_u1_n676 ) , .ZN( u0_u1_n677 ) , .A4( u0_u1_n717 ) , .A2( u0_u1_n860 ) );
  AOI221_X1 u0_u1_U62 (.ZN( u0_u1_n470 ) , .C2( u0_u1_n716 ) , .B2( u0_u1_n833 ) , .C1( u0_u1_n846 ) , .B1( u0_u1_n861 ) , .A( u0_u1_n865 ) );
  NOR4_X1 u0_u1_U63 (.A1( u0_u1_n468 ) , .ZN( u0_u1_n469 ) , .A4( u0_u1_n544 ) , .A2( u0_u1_n556 ) , .A3( u0_u1_n616 ) );
  NAND4_X1 u0_u1_U64 (.A4( u0_u1_n487 ) , .A3( u0_u1_n488 ) , .A2( u0_u1_n489 ) , .A1( u0_u1_n490 ) , .ZN( u0_u1_n780 ) );
  NOR4_X1 u0_u1_U65 (.A4( u0_u1_n486 ) , .ZN( u0_u1_n489 ) , .A1( u0_u1_n568 ) , .A2( u0_u1_n583 ) , .A3( u0_u1_n604 ) );
  NOR4_X1 u0_u1_U66 (.ZN( u0_u1_n488 ) , .A1( u0_u1_n509 ) , .A2( u0_u1_n521 ) , .A4( u0_u1_n548 ) , .A3( u0_u1_n613 ) );
  NOR2_X1 u0_u1_U67 (.ZN( u0_u1_n763 ) , .A1( u0_u1_n835 ) , .A2( u0_u1_n836 ) );
  NOR4_X1 u0_u1_U68 (.A4( u0_u1_n516 ) , .A3( u0_u1_n517 ) , .A2( u0_u1_n518 ) , .A1( u0_u1_n519 ) , .ZN( u0_u1_n526 ) );
  NOR4_X1 u0_u1_U69 (.A3( u0_u1_n523 ) , .A1( u0_u1_n524 ) , .ZN( u0_u1_n525 ) , .A2( u0_u1_n675 ) , .A4( u0_u1_n771 ) );
  NOR3_X1 u0_u1_U7 (.A3( u0_u1_n724 ) , .A1( u0_u1_n725 ) , .ZN( u0_u1_n742 ) , .A2( u0_u1_n743 ) );
  NAND4_X1 u0_u1_U70 (.A4( u0_u1_n475 ) , .A3( u0_u1_n476 ) , .A2( u0_u1_n477 ) , .A1( u0_u1_n478 ) , .ZN( u0_u1_n680 ) );
  NOR4_X1 u0_u1_U71 (.ZN( u0_u1_n476 ) , .A1( u0_u1_n508 ) , .A3( u0_u1_n546 ) , .A2( u0_u1_n585 ) , .A4( u0_u1_n718 ) );
  NOR4_X1 u0_u1_U72 (.ZN( u0_u1_n475 ) , .A2( u0_u1_n523 ) , .A4( u0_u1_n596 ) , .A1( u0_u1_n611 ) , .A3( u0_u1_n631 ) );
  NOR4_X1 u0_u1_U73 (.A4( u0_u1_n472 ) , .ZN( u0_u1_n478 ) , .A3( u0_u1_n558 ) , .A1( u0_u1_n737 ) , .A2( u0_u1_n757 ) );
  NAND4_X1 u0_u1_U74 (.A4( u0_u1_n458 ) , .A3( u0_u1_n459 ) , .A2( u0_u1_n460 ) , .A1( u0_u1_n461 ) , .ZN( u0_u1_n681 ) );
  NOR3_X1 u0_u1_U75 (.ZN( u0_u1_n459 ) , .A3( u0_u1_n532 ) , .A1( u0_u1_n557 ) , .A2( u0_u1_n572 ) );
  AOI221_X1 u0_u1_U76 (.A( u0_u1_n452 ) , .ZN( u0_u1_n461 ) , .C2( u0_u1_n755 ) , .B1( u0_u1_n834 ) , .C1( u0_u1_n843 ) , .B2( u0_u1_n862 ) );
  NOR4_X1 u0_u1_U77 (.ZN( u0_u1_n460 ) , .A2( u0_u1_n511 ) , .A1( u0_u1_n601 ) , .A4( u0_u1_n630 ) , .A3( u0_u1_n713 ) );
  INV_X1 u0_u1_U78 (.A( u0_u1_n671 ) , .ZN( u0_u1_n866 ) );
  NAND4_X1 u0_u1_U79 (.A4( u0_u1_n575 ) , .A3( u0_u1_n576 ) , .A1( u0_u1_n577 ) , .ZN( u0_u1_n725 ) , .A2( u0_u1_n875 ) );
  NOR3_X1 u0_u1_U8 (.ZN( u0_u1_n506 ) , .A2( u0_u1_n681 ) , .A3( u0_u1_n779 ) , .A1( u0_u1_n877 ) );
  NOR4_X1 u0_u1_U80 (.A4( u0_u1_n571 ) , .A3( u0_u1_n572 ) , .A2( u0_u1_n573 ) , .A1( u0_u1_n574 ) , .ZN( u0_u1_n575 ) );
  AOI221_X1 u0_u1_U81 (.A( u0_u1_n566 ) , .C2( u0_u1_n567 ) , .ZN( u0_u1_n576 ) , .B2( u0_u1_n846 ) , .B1( u0_u1_n853 ) , .C1( u0_u1_n854 ) );
  NOR2_X1 u0_u1_U82 (.ZN( u0_u1_n577 ) , .A1( u0_u1_n624 ) , .A2( u0_u1_n747 ) );
  INV_X1 u0_u1_U83 (.A( u0_u1_n764 ) , .ZN( u0_u1_n832 ) );
  NOR2_X1 u0_u1_U84 (.ZN( u0_u1_n649 ) , .A1( u0_u1_n855 ) , .A2( u0_u1_n869 ) );
  NOR4_X1 u0_u1_U85 (.A4( u0_u1_n579 ) , .A3( u0_u1_n580 ) , .A2( u0_u1_n581 ) , .ZN( u0_u1_n588 ) , .A1( u0_u1_n685 ) );
  NOR4_X1 u0_u1_U86 (.A1( u0_u1_n586 ) , .ZN( u0_u1_n587 ) , .A3( u0_u1_n654 ) , .A2( u0_u1_n664 ) , .A4( u0_u1_n769 ) );
  NAND4_X1 u0_u1_U87 (.A4( u0_u1_n721 ) , .A3( u0_u1_n722 ) , .A2( u0_u1_n723 ) , .ZN( u0_u1_n743 ) , .A1( u0_u1_n858 ) );
  NOR4_X1 u0_u1_U88 (.A4( u0_u1_n717 ) , .A3( u0_u1_n718 ) , .A2( u0_u1_n719 ) , .A1( u0_u1_n720 ) , .ZN( u0_u1_n721 ) );
  INV_X1 u0_u1_U89 (.A( u0_u1_n711 ) , .ZN( u0_u1_n858 ) );
  NOR2_X1 u0_u1_U9 (.ZN( u0_u1_n497 ) , .A1( u0_u1_n680 ) , .A2( u0_u1_n696 ) );
  AOI221_X1 u0_u1_U90 (.A( u0_u1_n712 ) , .ZN( u0_u1_n723 ) , .C2( u0_u1_n845 ) , .B2( u0_u1_n846 ) , .C1( u0_u1_n862 ) , .B1( u0_u1_n863 ) );
  INV_X1 u0_u1_U91 (.A( u0_u1_n465 ) , .ZN( u0_u1_n865 ) );
  OAI21_X1 u0_u1_U92 (.ZN( u0_u1_n465 ) , .B1( u0_u1_n811 ) , .A( u0_u1_n836 ) , .B2( u0_u1_n852 ) );
  INV_X1 u0_u1_U93 (.A( u0_u1_n793 ) , .ZN( u0_u1_n874 ) );
  OR4_X1 u0_u1_U94 (.A4( u0_u1_n568 ) , .A3( u0_u1_n569 ) , .A2( u0_u1_n570 ) , .ZN( u0_u1_n574 ) , .A1( u0_u1_n667 ) );
  OR4_X1 u0_u1_U95 (.A4( u0_u1_n520 ) , .A2( u0_u1_n521 ) , .A1( u0_u1_n522 ) , .ZN( u0_u1_n524 ) , .A3( u0_u1_n823 ) );
  OR4_X1 u0_u1_U96 (.ZN( u0_u1_n494 ) , .A4( u0_u1_n536 ) , .A2( u0_u1_n549 ) , .A1( u0_u1_n561 ) , .A3( u0_u1_n634 ) );
  OR4_X1 u0_u1_U97 (.ZN( u0_u1_n468 ) , .A4( u0_u1_n520 ) , .A3( u0_u1_n531 ) , .A2( u0_u1_n580 ) , .A1( u0_u1_n714 ) );
  OR4_X1 u0_u1_U98 (.A4( u0_u1_n684 ) , .A3( u0_u1_n685 ) , .A2( u0_u1_n686 ) , .A1( u0_u1_n687 ) , .ZN( u0_u1_n692 ) );
  OR3_X1 u0_u1_U99 (.A3( u0_u1_n508 ) , .A2( u0_u1_n509 ) , .A1( u0_u1_n510 ) , .ZN( u0_u1_n513 ) );
  NOR3_X1 us11_U10 (.ZN( us11_n504 ) , .A2( us11_n679 ) , .A3( us11_n777 ) , .A1( us11_n876 ) );
  NOR4_X1 us11_U100 (.A4( us11_n529 ) , .A3( us11_n530 ) , .ZN( us11_n537 ) , .A2( us11_n684 ) , .A1( us11_n794 ) );
  NAND4_X1 us11_U101 (.A4( us11_n479 ) , .A3( us11_n480 ) , .A2( us11_n481 ) , .A1( us11_n482 ) , .ZN( us11_n694 ) );
  NOR3_X1 us11_U102 (.ZN( us11_n480 ) , .A2( us11_n508 ) , .A3( us11_n601 ) , .A1( us11_n610 ) );
  AOI211_X1 us11_U103 (.B( us11_n477 ) , .A( us11_n478 ) , .ZN( us11_n482 ) , .C2( us11_n833 ) , .C1( us11_n861 ) );
  NOR4_X1 us11_U104 (.ZN( us11_n481 ) , .A3( us11_n532 ) , .A4( us11_n545 ) , .A2( us11_n567 ) , .A1( us11_n717 ) );
  NAND4_X1 us11_U105 (.A4( us11_n548 ) , .A3( us11_n549 ) , .A2( us11_n550 ) , .A1( us11_n551 ) , .ZN( us11_n745 ) );
  NOR3_X1 us11_U106 (.ZN( us11_n549 ) , .A2( us11_n651 ) , .A1( us11_n667 ) , .A3( us11_n771 ) );
  AOI211_X1 us11_U107 (.B( us11_n539 ) , .A( us11_n540 ) , .ZN( us11_n551 ) , .C2( us11_n839 ) , .C1( us11_n851 ) );
  NOR4_X1 us11_U108 (.A4( us11_n544 ) , .A3( us11_n545 ) , .A2( us11_n546 ) , .A1( us11_n547 ) , .ZN( us11_n548 ) );
  NOR4_X1 us11_U109 (.ZN( us11_n620 ) , .A1( us11_n656 ) , .A3( us11_n666 ) , .A4( us11_n682 ) , .A2( us11_n766 ) );
  INV_X1 us11_U11 (.A( us11_n706 ) , .ZN( us11_n876 ) );
  NOR4_X1 us11_U110 (.A4( us11_n609 ) , .A3( us11_n610 ) , .A2( us11_n611 ) , .A1( us11_n612 ) , .ZN( us11_n619 ) );
  NOR4_X1 us11_U111 (.A4( us11_n614 ) , .A3( us11_n615 ) , .A2( us11_n616 ) , .A1( us11_n617 ) , .ZN( us11_n618 ) );
  NOR2_X1 us11_U112 (.ZN( us11_n686 ) , .A1( us11_n831 ) , .A2( us11_n832 ) );
  NAND4_X1 us11_U113 (.A4( us11_n473 ) , .A3( us11_n474 ) , .A2( us11_n475 ) , .A1( us11_n476 ) , .ZN( us11_n678 ) );
  NOR4_X1 us11_U114 (.A4( us11_n470 ) , .ZN( us11_n476 ) , .A3( us11_n556 ) , .A1( us11_n735 ) , .A2( us11_n755 ) );
  NOR4_X1 us11_U115 (.ZN( us11_n475 ) , .A1( us11_n531 ) , .A3( us11_n568 ) , .A4( us11_n600 ) , .A2( us11_n642 ) );
  NOR4_X1 us11_U116 (.ZN( us11_n474 ) , .A1( us11_n506 ) , .A3( us11_n544 ) , .A2( us11_n583 ) , .A4( us11_n716 ) );
  NAND4_X1 us11_U117 (.A4( us11_n691 ) , .A3( us11_n692 ) , .A1( us11_n693 ) , .ZN( us11_n776 ) , .A2( us11_n872 ) );
  INV_X1 us11_U118 (.A( us11_n679 ) , .ZN( us11_n872 ) );
  NOR4_X1 us11_U119 (.A4( us11_n687 ) , .A3( us11_n688 ) , .A2( us11_n689 ) , .A1( us11_n690 ) , .ZN( us11_n691 ) );
  NOR3_X1 us11_U12 (.A3( us11_n621 ) , .A2( us11_n622 ) , .ZN( us11_n636 ) , .A1( us11_n725 ) );
  AOI221_X1 us11_U120 (.A( us11_n681 ) , .ZN( us11_n692 ) , .B2( us11_n840 ) , .C1( us11_n842 ) , .C2( us11_n862 ) , .B1( us11_n865 ) );
  NOR2_X1 us11_U121 (.ZN( us11_n733 ) , .A2( us11_n832 ) , .A1( us11_n845 ) );
  NAND4_X1 us11_U122 (.A4( us11_n719 ) , .A3( us11_n720 ) , .A2( us11_n721 ) , .ZN( us11_n741 ) , .A1( us11_n857 ) );
  AOI221_X1 us11_U123 (.A( us11_n710 ) , .ZN( us11_n721 ) , .C2( us11_n844 ) , .B2( us11_n845 ) , .C1( us11_n861 ) , .B1( us11_n862 ) );
  INV_X1 us11_U124 (.A( us11_n709 ) , .ZN( us11_n857 ) );
  NOR4_X1 us11_U125 (.A4( us11_n715 ) , .A3( us11_n716 ) , .A2( us11_n717 ) , .A1( us11_n718 ) , .ZN( us11_n719 ) );
  NAND4_X1 us11_U126 (.A4( us11_n573 ) , .A3( us11_n574 ) , .A1( us11_n575 ) , .ZN( us11_n723 ) , .A2( us11_n874 ) );
  NOR4_X1 us11_U127 (.A4( us11_n569 ) , .A3( us11_n570 ) , .A2( us11_n571 ) , .A1( us11_n572 ) , .ZN( us11_n573 ) );
  INV_X1 us11_U128 (.A( us11_n607 ) , .ZN( us11_n874 ) );
  NOR2_X1 us11_U129 (.ZN( us11_n575 ) , .A1( us11_n622 ) , .A2( us11_n745 ) );
  NOR2_X1 us11_U13 (.ZN( us11_n495 ) , .A1( us11_n678 ) , .A2( us11_n694 ) );
  NAND4_X1 us11_U130 (.A4( us11_n493 ) , .A3( us11_n494 ) , .A1( us11_n495 ) , .ZN( us11_n802 ) , .A2( us11_n867 ) );
  AOI221_X1 us11_U131 (.A( us11_n489 ) , .ZN( us11_n494 ) , .B2( us11_n836 ) , .C2( us11_n841 ) , .C1( us11_n851 ) , .B1( us11_n860 ) );
  INV_X1 us11_U132 (.A( us11_n778 ) , .ZN( us11_n867 ) );
  NOR4_X1 us11_U133 (.A2( us11_n491 ) , .A1( us11_n492 ) , .ZN( us11_n493 ) , .A3( us11_n580 ) , .A4( us11_n612 ) );
  NOR2_X1 us11_U134 (.ZN( us11_n647 ) , .A1( us11_n854 ) , .A2( us11_n868 ) );
  INV_X1 us11_U135 (.A( us11_n762 ) , .ZN( us11_n830 ) );
  NAND4_X1 us11_U136 (.A4( us11_n633 ) , .A3( us11_n634 ) , .A2( us11_n635 ) , .A1( us11_n636 ) , .ZN( us11_n743 ) );
  AOI211_X1 us11_U137 (.B( us11_n623 ) , .A( us11_n624 ) , .ZN( us11_n635 ) , .C2( us11_n836 ) , .C1( us11_n863 ) );
  NOR4_X1 us11_U138 (.A4( us11_n629 ) , .A3( us11_n630 ) , .A2( us11_n631 ) , .A1( us11_n632 ) , .ZN( us11_n633 ) );
  NOR4_X1 us11_U139 (.A4( us11_n626 ) , .A3( us11_n627 ) , .A2( us11_n628 ) , .ZN( us11_n634 ) , .A1( us11_n664 ) );
  NOR2_X1 us11_U14 (.A1( us11_n678 ) , .ZN( us11_n693 ) , .A2( us11_n807 ) );
  OR4_X1 us11_U140 (.A4( us11_n566 ) , .A3( us11_n567 ) , .A2( us11_n568 ) , .ZN( us11_n572 ) , .A1( us11_n665 ) );
  OR4_X1 us11_U141 (.A4( us11_n518 ) , .A2( us11_n519 ) , .A1( us11_n520 ) , .ZN( us11_n522 ) , .A3( us11_n821 ) );
  OR4_X1 us11_U142 (.ZN( us11_n492 ) , .A4( us11_n534 ) , .A2( us11_n547 ) , .A1( us11_n559 ) , .A3( us11_n632 ) );
  OR4_X1 us11_U143 (.A4( us11_n682 ) , .A3( us11_n683 ) , .A2( us11_n684 ) , .A1( us11_n685 ) , .ZN( us11_n690 ) );
  OR4_X1 us11_U144 (.ZN( us11_n466 ) , .A4( us11_n518 ) , .A3( us11_n529 ) , .A2( us11_n578 ) , .A1( us11_n712 ) );
  INV_X1 us11_U145 (.A( us11_n697 ) , .ZN( us11_n838 ) );
  OR4_X1 us11_U146 (.A4( us11_n580 ) , .A3( us11_n581 ) , .A2( us11_n582 ) , .A1( us11_n583 ) , .ZN( us11_n584 ) );
  NAND2_X1 us11_U147 (.ZN( us11_n613 ) , .A2( us11_n837 ) , .A1( us11_n873 ) );
  OR3_X1 us11_U148 (.A3( us11_n506 ) , .A2( us11_n507 ) , .A1( us11_n508 ) , .ZN( us11_n511 ) );
  INV_X1 us11_U149 (.A( us11_n463 ) , .ZN( us11_n864 ) );
  INV_X1 us11_U15 (.A( us11_n680 ) , .ZN( us11_n840 ) );
  OAI21_X1 us11_U150 (.ZN( us11_n463 ) , .B1( us11_n809 ) , .A( us11_n834 ) , .B2( us11_n851 ) );
  INV_X1 us11_U151 (.A( us11_n754 ) , .ZN( us11_n869 ) );
  OAI21_X1 us11_U152 (.B1( us11_n753 ) , .ZN( us11_n754 ) , .A( us11_n845 ) , .B2( us11_n868 ) );
  INV_X1 us11_U153 (.A( us11_n672 ) , .ZN( us11_n859 ) );
  AOI21_X1 us11_U154 (.A( us11_n670 ) , .B1( us11_n671 ) , .ZN( us11_n672 ) , .B2( us11_n856 ) );
  AOI222_X1 us11_U155 (.ZN( us11_n660 ) , .A2( us11_n839 ) , .B1( us11_n841 ) , .C2( us11_n845 ) , .A1( us11_n860 ) , .C1( us11_n863 ) , .B2( us11_n870 ) );
  INV_X1 us11_U156 (.A( us11_n647 ) , .ZN( us11_n870 ) );
  NAND2_X1 us11_U157 (.A1( us11_n447 ) , .A2( us11_n465 ) , .ZN( us11_n749 ) );
  OAI222_X1 us11_U158 (.ZN( us11_n617 ) , .B1( us11_n697 ) , .C1( us11_n724 ) , .C2( us11_n747 ) , .B2( us11_n786 ) , .A2( us11_n792 ) , .A1( us11_n816 ) );
  OAI222_X1 us11_U159 (.B2( us11_n708 ) , .ZN( us11_n709 ) , .C2( us11_n724 ) , .B1( us11_n747 ) , .A1( us11_n806 ) , .C1( us11_n814 ) , .A2( us11_n815 ) );
  NOR4_X1 us11_U16 (.A4( us11_n445 ) , .A3( us11_n446 ) , .A2( us11_n516 ) , .A1( us11_n541 ) , .ZN( us11_n706 ) );
  AOI22_X1 us11_U160 (.ZN( us11_n696 ) , .A1( us11_n830 ) , .B2( us11_n843 ) , .A2( us11_n865 ) , .B1( us11_n868 ) );
  AOI22_X1 us11_U161 (.A2( us11_n782 ) , .ZN( us11_n783 ) , .B2( us11_n831 ) , .A1( us11_n834 ) , .B1( us11_n863 ) );
  INV_X1 us11_U162 (.A( us11_n730 ) , .ZN( us11_n839 ) );
  AOI221_X1 us11_U163 (.A( us11_n564 ) , .C2( us11_n565 ) , .ZN( us11_n574 ) , .B2( us11_n845 ) , .B1( us11_n852 ) , .C1( us11_n853 ) );
  AOI21_X1 us11_U164 (.ZN( us11_n564 ) , .B1( us11_n724 ) , .A( us11_n779 ) , .B2( us11_n791 ) );
  NAND2_X1 us11_U165 (.A1( us11_n451 ) , .A2( us11_n453 ) , .ZN( us11_n762 ) );
  INV_X1 us11_U166 (.A( us11_n790 ) , .ZN( us11_n832 ) );
  OAI22_X1 us11_U167 (.ZN( us11_n637 ) , .A1( us11_n699 ) , .B2( us11_n728 ) , .A2( us11_n762 ) , .B1( us11_n816 ) );
  OAI221_X1 us11_U168 (.A( us11_n727 ) , .C2( us11_n728 ) , .B2( us11_n729 ) , .B1( us11_n730 ) , .ZN( us11_n737 ) , .C1( us11_n817 ) );
  AOI22_X1 us11_U169 (.ZN( us11_n727 ) , .B1( us11_n832 ) , .A2( us11_n838 ) , .A1( us11_n863 ) , .B2( us11_n866 ) );
  OR3_X1 us11_U17 (.ZN( us11_n446 ) , .A1( us11_n528 ) , .A3( us11_n577 ) , .A2( us11_n875 ) );
  INV_X1 us11_U170 (.A( us11_n747 ) , .ZN( us11_n834 ) );
  OAI22_X1 us11_U171 (.ZN( us11_n624 ) , .B1( us11_n669 ) , .B2( us11_n747 ) , .A1( us11_n815 ) , .A2( us11_n816 ) );
  OAI22_X1 us11_U172 (.ZN( us11_n489 ) , .A1( us11_n724 ) , .B2( us11_n728 ) , .B1( us11_n730 ) , .A2( us11_n779 ) );
  OAI22_X1 us11_U173 (.B2( us11_n779 ) , .B1( us11_n780 ) , .ZN( us11_n781 ) , .A2( us11_n814 ) , .A1( us11_n815 ) );
  OAI22_X1 us11_U174 (.A1( us11_n724 ) , .ZN( us11_n726 ) , .B2( us11_n750 ) , .B1( us11_n812 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U175 (.ZN( us11_n630 ) , .A1( us11_n747 ) , .A2( us11_n815 ) );
  OAI22_X1 us11_U176 (.B2( us11_n750 ) , .B1( us11_n751 ) , .A1( us11_n752 ) , .ZN( us11_n756 ) , .A2( us11_n806 ) );
  NOR3_X1 us11_U177 (.ZN( us11_n752 ) , .A2( us11_n853 ) , .A1( us11_n863 ) , .A3( us11_n865 ) );
  NOR2_X1 us11_U178 (.ZN( us11_n751 ) , .A2( us11_n852 ) , .A1( us11_n860 ) );
  OAI22_X1 us11_U179 (.B2( us11_n803 ) , .B1( us11_n804 ) , .A2( us11_n805 ) , .A1( us11_n806 ) , .ZN( us11_n808 ) );
  OR4_X1 us11_U18 (.A4( us11_n442 ) , .A2( us11_n443 ) , .A1( us11_n444 ) , .ZN( us11_n445 ) , .A3( us11_n553 ) );
  NOR2_X1 us11_U180 (.ZN( us11_n656 ) , .A1( us11_n747 ) , .A2( us11_n780 ) );
  OAI22_X1 us11_U181 (.B2( us11_n744 ) , .ZN( us11_n746 ) , .A2( us11_n762 ) , .B1( us11_n780 ) , .A1( us11_n792 ) );
  OAI22_X1 us11_U182 (.ZN( us11_n496 ) , .A2( us11_n744 ) , .A1( us11_n780 ) , .B1( us11_n791 ) , .B2( us11_n806 ) );
  OAI22_X1 us11_U183 (.ZN( us11_n695 ) , .A2( us11_n730 ) , .A1( us11_n780 ) , .B1( us11_n791 ) , .B2( us11_n817 ) );
  INV_X1 us11_U184 (.A( us11_n744 ) , .ZN( us11_n837 ) );
  INV_X1 us11_U185 (.A( us11_n805 ) , .ZN( us11_n860 ) );
  INV_X1 us11_U186 (.A( us11_n816 ) , .ZN( us11_n831 ) );
  INV_X1 us11_U187 (.A( us11_n788 ) , .ZN( us11_n845 ) );
  OAI22_X1 us11_U188 (.ZN( us11_n590 ) , .B1( us11_n730 ) , .B2( us11_n749 ) , .A2( us11_n786 ) , .A1( us11_n803 ) );
  OAI22_X1 us11_U189 (.B1( us11_n490 ) , .ZN( us11_n491 ) , .A1( us11_n686 ) , .A2( us11_n763 ) , .B2( us11_n817 ) );
  INV_X1 us11_U19 (.A( us11_n613 ) , .ZN( us11_n875 ) );
  NOR3_X1 us11_U190 (.ZN( us11_n490 ) , .A1( us11_n782 ) , .A2( us11_n850 ) , .A3( us11_n863 ) );
  OAI22_X1 us11_U191 (.ZN( us11_n710 ) , .A2( us11_n728 ) , .B2( us11_n729 ) , .A1( us11_n744 ) , .B1( us11_n813 ) );
  INV_X1 us11_U192 (.A( us11_n792 ) , .ZN( us11_n851 ) );
  NOR2_X1 us11_U193 (.ZN( us11_n715 ) , .A1( us11_n805 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U194 (.A1( us11_n699 ) , .ZN( us11_n768 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U195 (.ZN( us11_n541 ) , .A2( us11_n697 ) , .A1( us11_n699 ) );
  INV_X1 us11_U196 (.A( us11_n814 ) , .ZN( us11_n833 ) );
  NOR2_X1 us11_U197 (.A1( us11_n669 ) , .ZN( us11_n673 ) , .A2( us11_n744 ) );
  NOR2_X1 us11_U198 (.ZN( us11_n602 ) , .A1( us11_n669 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U199 (.A1( us11_n669 ) , .ZN( us11_n688 ) , .A2( us11_n816 ) );
  INV_X1 us11_U20 (.A( us11_n749 ) , .ZN( us11_n863 ) );
  NOR2_X1 us11_U200 (.A2( us11_n744 ) , .ZN( us11_n755 ) , .A1( us11_n805 ) );
  NOR2_X1 us11_U201 (.ZN( us11_n735 ) , .A2( us11_n803 ) , .A1( us11_n805 ) );
  NOR2_X1 us11_U202 (.A1( us11_n669 ) , .ZN( us11_n766 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U203 (.ZN( us11_n527 ) , .A1( us11_n669 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U204 (.ZN( us11_n666 ) , .A1( us11_n728 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U205 (.ZN( us11_n594 ) , .A2( us11_n697 ) , .A1( us11_n728 ) );
  NOR2_X1 us11_U206 (.ZN( us11_n718 ) , .A2( us11_n724 ) , .A1( us11_n744 ) );
  NOR2_X1 us11_U207 (.ZN( us11_n570 ) , .A1( us11_n728 ) , .A2( us11_n806 ) );
  NOR2_X1 us11_U208 (.ZN( us11_n661 ) , .A1( us11_n729 ) , .A2( us11_n790 ) );
  OAI22_X1 us11_U209 (.ZN( us11_n483 ) , .A1( us11_n708 ) , .B2( us11_n785 ) , .A2( us11_n806 ) , .B1( us11_n812 ) );
  AOI222_X1 us11_U21 (.ZN( us11_n563 ) , .B1( us11_n830 ) , .C1( us11_n841 ) , .A2( us11_n843 ) , .A1( us11_n854 ) , .B2( us11_n863 ) , .C2( us11_n873 ) );
  NOR2_X1 us11_U210 (.ZN( us11_n601 ) , .A2( us11_n780 ) , .A1( us11_n803 ) );
  NOR2_X1 us11_U211 (.ZN( us11_n531 ) , .A2( us11_n780 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U212 (.ZN( us11_n654 ) , .A1( us11_n728 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U213 (.ZN( us11_n509 ) , .A1( us11_n729 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U214 (.ZN( us11_n599 ) , .A2( us11_n791 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U215 (.ZN( us11_n612 ) , .A1( us11_n779 ) , .A2( us11_n786 ) );
  NOR2_X1 us11_U216 (.ZN( us11_n546 ) , .A2( us11_n780 ) , .A1( us11_n814 ) );
  INV_X1 us11_U217 (.A( us11_n750 ) , .ZN( us11_n842 ) );
  NOR2_X1 us11_U218 (.ZN( us11_n532 ) , .A2( us11_n749 ) , .A1( us11_n750 ) );
  NOR2_X1 us11_U219 (.ZN( us11_n528 ) , .A2( us11_n724 ) , .A1( us11_n803 ) );
  NOR4_X1 us11_U22 (.ZN( us11_n479 ) , .A1( us11_n520 ) , .A4( us11_n557 ) , .A3( us11_n582 ) , .A2( us11_n630 ) );
  NOR2_X1 us11_U220 (.ZN( us11_n577 ) , .A2( us11_n699 ) , .A1( us11_n814 ) );
  AOI21_X1 us11_U221 (.ZN( us11_n640 ) , .B2( us11_n747 ) , .A( us11_n792 ) , .B1( us11_n803 ) );
  NOR2_X1 us11_U222 (.ZN( us11_n615 ) , .A1( us11_n785 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U223 (.ZN( us11_n629 ) , .A2( us11_n728 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U224 (.ZN( us11_n663 ) , .A1( us11_n729 ) , .A2( us11_n785 ) );
  NOR2_X1 us11_U225 (.ZN( us11_n628 ) , .A2( us11_n669 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U226 (.ZN( us11_n611 ) , .A2( us11_n780 ) , .A1( us11_n806 ) );
  NOR2_X1 us11_U227 (.A2( us11_n744 ) , .ZN( us11_n769 ) , .A1( us11_n812 ) );
  NOR2_X1 us11_U228 (.ZN( us11_n567 ) , .A1( us11_n747 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U229 (.A2( us11_n708 ) , .A1( us11_n750 ) , .ZN( us11_n771 ) );
  NOR4_X1 us11_U23 (.ZN( us11_n473 ) , .A2( us11_n521 ) , .A4( us11_n594 ) , .A1( us11_n609 ) , .A3( us11_n629 ) );
  NOR2_X1 us11_U230 (.ZN( us11_n557 ) , .A1( us11_n792 ) , .A2( us11_n814 ) );
  NOR2_X1 us11_U231 (.A2( us11_n697 ) , .ZN( us11_n716 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U232 (.ZN( us11_n544 ) , .A2( us11_n785 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U233 (.ZN( us11_n667 ) , .A1( us11_n750 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U234 (.ZN( us11_n555 ) , .A1( us11_n750 ) , .A2( us11_n791 ) );
  NOR2_X1 us11_U235 (.ZN( us11_n508 ) , .A2( us11_n780 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U236 (.ZN( us11_n543 ) , .A2( us11_n708 ) , .A1( us11_n785 ) );
  NOR2_X1 us11_U237 (.ZN( us11_n664 ) , .A1( us11_n785 ) , .A2( us11_n791 ) );
  OAI22_X1 us11_U238 (.B1( us11_n440 ) , .ZN( us11_n444 ) , .A2( us11_n728 ) , .A1( us11_n744 ) , .B2( us11_n749 ) );
  NOR3_X1 us11_U239 (.ZN( us11_n440 ) , .A2( us11_n836 ) , .A3( us11_n837 ) , .A1( us11_n846 ) );
  NOR4_X1 us11_U24 (.ZN( us11_n485 ) , .A2( us11_n533 ) , .A1( us11_n558 ) , .A3( us11_n631 ) , .A4( us11_n718 ) );
  NOR2_X1 us11_U240 (.ZN( us11_n631 ) , .A1( us11_n724 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U241 (.ZN( us11_n556 ) , .A1( us11_n762 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U242 (.ZN( us11_n530 ) , .A2( us11_n744 ) , .A1( us11_n792 ) );
  NOR2_X1 us11_U243 (.ZN( us11_n507 ) , .A1( us11_n812 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U244 (.ZN( us11_n516 ) , .A1( us11_n708 ) , .A2( us11_n744 ) );
  NOR2_X1 us11_U245 (.ZN( us11_n558 ) , .A1( us11_n708 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U246 (.ZN( us11_n517 ) , .A1( us11_n708 ) , .A2( us11_n803 ) );
  INV_X1 us11_U247 (.A( us11_n806 ) , .ZN( us11_n841 ) );
  NOR2_X1 us11_U248 (.ZN( us11_n545 ) , .A1( us11_n749 ) , .A2( us11_n814 ) );
  INV_X1 us11_U249 (.A( us11_n728 ) , .ZN( us11_n852 ) );
  NOR4_X1 us11_U25 (.A4( us11_n532 ) , .A3( us11_n533 ) , .A2( us11_n534 ) , .ZN( us11_n535 ) , .A1( us11_n820 ) );
  NOR2_X1 us11_U250 (.ZN( us11_n554 ) , .A1( us11_n786 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U251 (.ZN( us11_n670 ) , .A1( us11_n790 ) , .A2( us11_n805 ) );
  NOR2_X1 us11_U252 (.ZN( us11_n717 ) , .A2( us11_n744 ) , .A1( us11_n786 ) );
  NOR2_X1 us11_U253 (.ZN( us11_n506 ) , .A2( us11_n728 ) , .A1( us11_n762 ) );
  NOR2_X1 us11_U254 (.ZN( us11_n642 ) , .A2( us11_n788 ) , .A1( us11_n791 ) );
  NOR2_X1 us11_U255 (.ZN( us11_n614 ) , .A1( us11_n762 ) , .A2( us11_n812 ) );
  AOI21_X1 us11_U256 (.ZN( us11_n626 ) , .B2( us11_n669 ) , .A( us11_n790 ) , .B1( us11_n791 ) );
  AOI21_X1 us11_U257 (.ZN( us11_n552 ) , .B1( us11_n669 ) , .A( us11_n697 ) , .B2( us11_n805 ) );
  AOI21_X1 us11_U258 (.ZN( us11_n589 ) , .B2( us11_n699 ) , .B1( us11_n815 ) , .A( us11_n817 ) );
  INV_X1 us11_U259 (.A( us11_n763 ) , .ZN( us11_n866 ) );
  NOR4_X1 us11_U26 (.ZN( us11_n456 ) , .A2( us11_n517 ) , .A1( us11_n543 ) , .A3( us11_n579 ) , .A4( us11_n615 ) );
  NOR2_X1 us11_U260 (.ZN( us11_n609 ) , .A2( us11_n724 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U261 (.ZN( us11_n668 ) , .A2( us11_n708 ) , .A1( us11_n790 ) );
  NOR2_X1 us11_U262 (.ZN( us11_n533 ) , .A2( us11_n724 ) , .A1( us11_n730 ) );
  NOR2_X1 us11_U263 (.ZN( us11_n521 ) , .A1( us11_n790 ) , .A2( us11_n812 ) );
  AOI21_X1 us11_U264 (.A( us11_n815 ) , .B2( us11_n816 ) , .B1( us11_n817 ) , .ZN( us11_n818 ) );
  NOR2_X1 us11_U265 (.ZN( us11_n547 ) , .A1( us11_n699 ) , .A2( us11_n744 ) );
  AOI21_X1 us11_U266 (.ZN( us11_n510 ) , .B2( us11_n669 ) , .A( us11_n730 ) , .B1( us11_n815 ) );
  NOR2_X1 us11_U267 (.ZN( us11_n655 ) , .A1( us11_n790 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U268 (.ZN( us11_n579 ) , .A2( us11_n708 ) , .A1( us11_n730 ) );
  INV_X1 us11_U269 (.A( us11_n729 ) , .ZN( us11_n868 ) );
  NOR4_X1 us11_U27 (.A4( us11_n577 ) , .A3( us11_n578 ) , .A2( us11_n579 ) , .ZN( us11_n586 ) , .A1( us11_n683 ) );
  NOR2_X1 us11_U270 (.ZN( us11_n542 ) , .A1( us11_n762 ) , .A2( us11_n791 ) );
  NOR2_X1 us11_U271 (.ZN( us11_n701 ) , .A2( us11_n786 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U272 (.A2( us11_n708 ) , .A1( us11_n762 ) , .ZN( us11_n794 ) );
  AOI21_X1 us11_U273 (.ZN( us11_n499 ) , .B1( us11_n680 ) , .A( us11_n812 ) , .B2( us11_n816 ) );
  AOI21_X1 us11_U274 (.ZN( us11_n650 ) , .A( us11_n779 ) , .B1( us11_n792 ) , .B2( us11_n805 ) );
  INV_X1 us11_U275 (.A( us11_n699 ) , .ZN( us11_n853 ) );
  NOR2_X1 us11_U276 (.ZN( us11_n652 ) , .A1( us11_n669 ) , .A2( us11_n814 ) );
  NOR2_X1 us11_U277 (.ZN( us11_n581 ) , .A1( us11_n669 ) , .A2( us11_n788 ) );
  AOI21_X1 us11_U278 (.ZN( us11_n515 ) , .A( us11_n729 ) , .B1( us11_n750 ) , .B2( us11_n803 ) );
  AOI21_X1 us11_U279 (.B1( us11_n699 ) , .ZN( us11_n700 ) , .A( us11_n732 ) , .B2( us11_n763 ) );
  AOI222_X1 us11_U28 (.B2( us11_n638 ) , .ZN( us11_n644 ) , .B1( us11_n841 ) , .A1( us11_n842 ) , .C2( us11_n846 ) , .C1( us11_n863 ) , .A2( us11_n865 ) );
  AOI21_X1 us11_U280 (.ZN( us11_n591 ) , .B2( us11_n763 ) , .A( us11_n785 ) , .B1( us11_n812 ) );
  AOI21_X1 us11_U281 (.A( us11_n812 ) , .B2( us11_n813 ) , .B1( us11_n814 ) , .ZN( us11_n819 ) );
  NOR2_X1 us11_U282 (.A1( us11_n730 ) , .ZN( us11_n765 ) , .A2( us11_n786 ) );
  INV_X1 us11_U283 (.A( us11_n791 ) , .ZN( us11_n873 ) );
  AOI21_X1 us11_U284 (.ZN( us11_n593 ) , .B1( us11_n750 ) , .A( us11_n792 ) , .B2( us11_n813 ) );
  NOR2_X1 us11_U285 (.ZN( us11_n582 ) , .A1( us11_n744 ) , .A2( us11_n815 ) );
  NOR2_X1 us11_U286 (.ZN( us11_n519 ) , .A2( us11_n699 ) , .A1( us11_n816 ) );
  NOR2_X1 us11_U287 (.ZN( us11_n685 ) , .A1( us11_n729 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U288 (.ZN( us11_n559 ) , .A2( us11_n791 ) , .A1( us11_n803 ) );
  AOI21_X1 us11_U289 (.ZN( us11_n649 ) , .B1( us11_n729 ) , .B2( us11_n763 ) , .A( us11_n813 ) );
  NOR4_X1 us11_U29 (.A4( us11_n639 ) , .A3( us11_n640 ) , .A2( us11_n641 ) , .A1( us11_n642 ) , .ZN( us11_n643 ) );
  AOI21_X1 us11_U290 (.B1( us11_n625 ) , .ZN( us11_n627 ) , .A( us11_n763 ) , .B2( us11_n814 ) );
  NOR2_X1 us11_U291 (.ZN( us11_n683 ) , .A2( us11_n699 ) , .A1( us11_n803 ) );
  NOR2_X1 us11_U292 (.A2( us11_n697 ) , .A1( us11_n780 ) , .ZN( us11_n820 ) );
  NOR2_X1 us11_U293 (.ZN( us11_n653 ) , .A1( us11_n762 ) , .A2( us11_n786 ) );
  NOR2_X1 us11_U294 (.ZN( us11_n568 ) , .A1( us11_n729 ) , .A2( us11_n762 ) );
  NOR2_X1 us11_U295 (.ZN( us11_n662 ) , .A2( us11_n697 ) , .A1( us11_n729 ) );
  INV_X1 us11_U296 (.A( us11_n813 ) , .ZN( us11_n836 ) );
  NOR2_X1 us11_U297 (.ZN( us11_n566 ) , .A2( us11_n697 ) , .A1( us11_n763 ) );
  NOR2_X1 us11_U298 (.ZN( us11_n520 ) , .A2( us11_n708 ) , .A1( us11_n814 ) );
  AOI21_X1 us11_U299 (.ZN( us11_n477 ) , .A( us11_n669 ) , .B1( us11_n750 ) , .B2( us11_n806 ) );
  NAND2_X2 us11_U3 (.A2( us11_n460 ) , .A1( us11_n465 ) , .ZN( us11_n780 ) );
  NOR3_X1 us11_U30 (.A2( us11_n607 ) , .A1( us11_n608 ) , .ZN( us11_n646 ) , .A3( us11_n722 ) );
  NOR2_X1 us11_U300 (.A1( us11_n697 ) , .ZN( us11_n770 ) , .A2( us11_n815 ) );
  AOI21_X1 us11_U301 (.ZN( us11_n514 ) , .A( us11_n779 ) , .B2( us11_n792 ) , .B1( us11_n812 ) );
  INV_X1 us11_U302 (.A( us11_n786 ) , .ZN( us11_n862 ) );
  AOI21_X1 us11_U303 (.ZN( us11_n540 ) , .A( us11_n763 ) , .B2( us11_n779 ) , .B1( us11_n817 ) );
  AOI21_X1 us11_U304 (.ZN( us11_n450 ) , .B2( us11_n792 ) , .A( us11_n803 ) , .B1( us11_n815 ) );
  AOI21_X1 us11_U305 (.ZN( us11_n539 ) , .B2( us11_n812 ) , .A( us11_n814 ) , .B1( us11_n815 ) );
  NOR2_X1 us11_U306 (.ZN( us11_n529 ) , .A1( us11_n708 ) , .A2( us11_n779 ) );
  NOR2_X1 us11_U307 (.ZN( us11_n578 ) , .A1( us11_n708 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U308 (.ZN( us11_n583 ) , .A1( us11_n792 ) , .A2( us11_n817 ) );
  NOR2_X1 us11_U309 (.ZN( us11_n534 ) , .A1( us11_n724 ) , .A2( us11_n788 ) );
  NOR4_X1 us11_U31 (.A4( us11_n541 ) , .A3( us11_n542 ) , .A2( us11_n543 ) , .ZN( us11_n550 ) , .A1( us11_n688 ) );
  NOR2_X1 us11_U310 (.ZN( us11_n632 ) , .A2( us11_n697 ) , .A1( us11_n724 ) );
  AOI21_X1 us11_U311 (.ZN( us11_n498 ) , .A( us11_n724 ) , .B2( us11_n762 ) , .B1( us11_n814 ) );
  AOI21_X1 us11_U312 (.A( us11_n790 ) , .B2( us11_n791 ) , .B1( us11_n792 ) , .ZN( us11_n793 ) );
  AOI21_X1 us11_U313 (.ZN( us11_n689 ) , .B2( us11_n749 ) , .B1( us11_n763 ) , .A( us11_n806 ) );
  AOI21_X1 us11_U314 (.B1( us11_n686 ) , .ZN( us11_n687 ) , .A( us11_n728 ) , .B2( us11_n761 ) );
  AOI21_X1 us11_U315 (.ZN( us11_n569 ) , .B1( us11_n750 ) , .B2( us11_n762 ) , .A( us11_n780 ) );
  AOI21_X1 us11_U316 (.ZN( us11_n500 ) , .A( us11_n697 ) , .B1( us11_n708 ) , .B2( us11_n786 ) );
  NOR2_X1 us11_U317 (.ZN( us11_n665 ) , .A1( us11_n780 ) , .A2( us11_n813 ) );
  NOR2_X1 us11_U318 (.ZN( us11_n580 ) , .A2( us11_n697 ) , .A1( us11_n791 ) );
  AOI21_X1 us11_U319 (.ZN( us11_n571 ) , .B2( us11_n697 ) , .B1( us11_n806 ) , .A( us11_n812 ) );
  AOI221_X1 us11_U32 (.A( us11_n713 ) , .B2( us11_n714 ) , .ZN( us11_n720 ) , .C1( us11_n832 ) , .B1( us11_n839 ) , .C2( us11_n863 ) );
  NOR2_X1 us11_U320 (.ZN( us11_n684 ) , .A1( us11_n791 ) , .A2( us11_n813 ) );
  AOI21_X1 us11_U321 (.ZN( us11_n639 ) , .B2( us11_n749 ) , .A( us11_n788 ) , .B1( us11_n812 ) );
  AOI21_X1 us11_U322 (.A( us11_n733 ) , .ZN( us11_n734 ) , .B2( us11_n780 ) , .B1( us11_n792 ) );
  NAND2_X2 us11_U323 (.A1( us11_n452 ) , .A2( us11_n465 ) , .ZN( us11_n669 ) );
  NOR2_X1 us11_U324 (.ZN( us11_n711 ) , .A1( us11_n762 ) , .A2( us11_n763 ) );
  AOI21_X1 us11_U325 (.ZN( us11_n478 ) , .B2( us11_n697 ) , .A( us11_n749 ) , .B1( us11_n779 ) );
  NOR2_X1 us11_U326 (.A2( us11_n813 ) , .A1( us11_n815 ) , .ZN( us11_n821 ) );
  NOR2_X1 us11_U327 (.A1( us11_n749 ) , .ZN( us11_n767 ) , .A2( us11_n803 ) );
  NOR2_X1 us11_U328 (.ZN( us11_n682 ) , .A2( us11_n708 ) , .A1( us11_n817 ) );
  NAND2_X2 us11_U329 (.A1( us11_n451 ) , .A2( us11_n471 ) , .ZN( us11_n816 ) );
  OR2_X1 us11_U33 (.A2( us11_n711 ) , .A1( us11_n712 ) , .ZN( us11_n713 ) );
  AOI21_X1 us11_U330 (.ZN( us11_n641 ) , .B1( us11_n680 ) , .A( us11_n791 ) , .B2( us11_n817 ) );
  NAND2_X1 us11_U331 (.ZN( us11_n753 ) , .A1( us11_n763 ) , .A2( us11_n805 ) );
  OAI21_X1 us11_U332 (.A( us11_n731 ) , .B1( us11_n732 ) , .ZN( us11_n736 ) , .B2( us11_n805 ) );
  OAI21_X1 us11_U333 (.ZN( us11_n731 ) , .A( us11_n833 ) , .B2( us11_n852 ) , .B1( us11_n873 ) );
  INV_X1 us11_U334 (.A( us11_n815 ) , .ZN( us11_n855 ) );
  NAND2_X2 us11_U335 (.A1( us11_n447 ) , .A2( us11_n449 ) , .ZN( us11_n805 ) );
  NAND2_X2 us11_U336 (.A2( us11_n449 ) , .A1( us11_n452 ) , .ZN( us11_n763 ) );
  AOI21_X1 us11_U337 (.ZN( us11_n442 ) , .A( us11_n699 ) , .B1( us11_n733 ) , .B2( us11_n750 ) );
  OAI21_X1 us11_U338 (.A( us11_n698 ) , .ZN( us11_n702 ) , .B2( us11_n750 ) , .B1( us11_n804 ) );
  OAI21_X1 us11_U339 (.ZN( us11_n698 ) , .B2( us11_n833 ) , .B1( us11_n838 ) , .A( us11_n860 ) );
  NOR2_X1 us11_U34 (.ZN( us11_n680 ) , .A2( us11_n834 ) , .A1( us11_n839 ) );
  NAND2_X1 us11_U340 (.A1( us11_n699 ) , .A2( us11_n729 ) , .ZN( us11_n782 ) );
  NOR2_X1 us11_U341 (.ZN( us11_n526 ) , .A1( us11_n724 ) , .A2( us11_n750 ) );
  INV_X1 us11_U342 (.A( us11_n780 ) , .ZN( us11_n850 ) );
  NOR2_X1 us11_U343 (.ZN( us11_n518 ) , .A1( us11_n708 ) , .A2( us11_n788 ) );
  AOI21_X1 us11_U344 (.ZN( us11_n443 ) , .B1( us11_n789 ) , .B2( us11_n791 ) , .A( us11_n814 ) );
  AOI21_X1 us11_U345 (.ZN( us11_n497 ) , .A( us11_n779 ) , .B2( us11_n791 ) , .B1( us11_n804 ) );
  NAND2_X2 us11_U346 (.A2( us11_n441 ) , .A1( us11_n447 ) , .ZN( us11_n784 ) );
  NAND2_X1 us11_U347 (.ZN( us11_n714 ) , .A1( us11_n728 ) , .A2( us11_n780 ) );
  NOR2_X1 us11_U348 (.ZN( us11_n484 ) , .A1( us11_n788 ) , .A2( us11_n805 ) );
  OAI21_X1 us11_U349 (.A( us11_n787 ) , .B2( us11_n788 ) , .B1( us11_n789 ) , .ZN( us11_n795 ) );
  AOI222_X1 us11_U35 (.ZN( us11_n469 ) , .B1( us11_n832 ) , .A1( us11_n839 ) , .C1( us11_n842 ) , .C2( us11_n851 ) , .A2( us11_n855 ) , .B2( us11_n865 ) );
  NAND2_X2 us11_U350 (.A2( us11_n448 ) , .A1( us11_n452 ) , .ZN( us11_n729 ) );
  OAI21_X1 us11_U351 (.ZN( us11_n787 ) , .A( us11_n839 ) , .B1( us11_n863 ) , .B2( us11_n873 ) );
  NAND2_X1 us11_U352 (.A2( us11_n762 ) , .A1( us11_n806 ) , .ZN( us11_n810 ) );
  INV_X1 us11_U353 (.A( us11_n785 ) , .ZN( us11_n846 ) );
  NOR2_X1 us11_U354 (.ZN( us11_n470 ) , .A2( us11_n779 ) , .A1( us11_n815 ) );
  NOR2_X1 us11_U355 (.ZN( us11_n712 ) , .A2( us11_n724 ) , .A1( us11_n790 ) );
  NAND2_X1 us11_U356 (.ZN( us11_n671 ) , .A1( us11_n806 ) , .A2( us11_n816 ) );
  NAND2_X1 us11_U357 (.A2( us11_n749 ) , .A1( us11_n786 ) , .ZN( us11_n809 ) );
  INV_X1 us11_U358 (.A( us11_n724 ) , .ZN( us11_n856 ) );
  INV_X1 us11_U359 (.A( us11_n817 ) , .ZN( us11_n844 ) );
  NOR4_X1 us11_U36 (.A1( us11_n466 ) , .ZN( us11_n467 ) , .A4( us11_n542 ) , .A2( us11_n554 ) , .A3( us11_n614 ) );
  AND2_X1 us11_U360 (.ZN( us11_n732 ) , .A1( us11_n779 ) , .A2( us11_n785 ) );
  AOI221_X1 us11_U361 (.A( us11_n764 ) , .ZN( us11_n774 ) , .C2( us11_n810 ) , .B2( us11_n835 ) , .C1( us11_n855 ) , .B1( us11_n866 ) );
  AOI21_X1 us11_U362 (.B2( us11_n763 ) , .ZN( us11_n764 ) , .A( us11_n788 ) , .B1( us11_n792 ) );
  INV_X1 us11_U363 (.A( us11_n761 ) , .ZN( us11_n835 ) );
  NAND2_X1 us11_U364 (.A2( us11_n448 ) , .A1( us11_n460 ) , .ZN( us11_n728 ) );
  NAND2_X1 us11_U365 (.A1( us11_n451 ) , .A2( us11_n454 ) , .ZN( us11_n814 ) );
  NAND2_X1 us11_U366 (.A1( us11_n455 ) , .A2( us11_n462 ) , .ZN( us11_n750 ) );
  NAND2_X1 us11_U367 (.A2( us11_n454 ) , .A1( us11_n472 ) , .ZN( us11_n779 ) );
  NAND2_X1 us11_U368 (.A2( us11_n453 ) , .A1( us11_n455 ) , .ZN( us11_n806 ) );
  NAND2_X1 us11_U369 (.A1( us11_n453 ) , .A2( us11_n472 ) , .ZN( us11_n785 ) );
  AOI221_X1 us11_U37 (.ZN( us11_n468 ) , .C2( us11_n714 ) , .B2( us11_n831 ) , .C1( us11_n845 ) , .B1( us11_n860 ) , .A( us11_n864 ) );
  NAND2_X1 us11_U370 (.A2( us11_n464 ) , .A1( us11_n465 ) , .ZN( us11_n812 ) );
  NAND2_X1 us11_U371 (.A1( us11_n447 ) , .A2( us11_n448 ) , .ZN( us11_n786 ) );
  NAND2_X2 us11_U372 (.A1( us11_n455 ) , .A2( us11_n471 ) , .ZN( us11_n803 ) );
  NAND2_X1 us11_U373 (.A1( us11_n462 ) , .A2( us11_n472 ) , .ZN( us11_n788 ) );
  NOR2_X1 us11_U374 (.ZN( us11_n465 ) , .A2( us11_n847 ) , .A1( us11_n848 ) );
  NAND2_X2 us11_U375 (.A1( us11_n453 ) , .A2( us11_n461 ) , .ZN( us11_n744 ) );
  NOR2_X1 us11_U376 (.ZN( us11_n453 ) , .A1( us11_n826 ) , .A2( us11_n827 ) );
  NOR2_X1 us11_U377 (.ZN( us11_n451 ) , .A1( us11_n828 ) , .A2( us11_n829 ) );
  NAND2_X1 us11_U378 (.A2( us11_n454 ) , .A1( us11_n455 ) , .ZN( us11_n730 ) );
  NAND2_X1 us11_U379 (.A1( us11_n451 ) , .A2( us11_n462 ) , .ZN( us11_n790 ) );
  NOR4_X1 us11_U38 (.A4( us11_n514 ) , .A3( us11_n515 ) , .A2( us11_n516 ) , .A1( us11_n517 ) , .ZN( us11_n524 ) );
  NAND2_X2 us11_U380 (.A1( us11_n449 ) , .A2( us11_n460 ) , .ZN( us11_n792 ) );
  NAND2_X2 us11_U381 (.A2( us11_n448 ) , .A1( us11_n464 ) , .ZN( us11_n815 ) );
  NAND2_X2 us11_U382 (.A2( us11_n471 ) , .A1( us11_n472 ) , .ZN( us11_n817 ) );
  NAND2_X2 us11_U383 (.A1( us11_n441 ) , .A2( us11_n460 ) , .ZN( us11_n699 ) );
  NOR2_X1 us11_U384 (.ZN( us11_n447 ) , .A2( us11_n849 ) , .A1( us11_n858 ) );
  NOR2_X1 us11_U385 (.A2( sa11_6 ) , .A1( sa11_7 ) , .ZN( us11_n464 ) );
  NOR2_X1 us11_U386 (.A2( sa11_7 ) , .ZN( us11_n460 ) , .A1( us11_n849 ) );
  NOR2_X1 us11_U387 (.A2( sa11_5 ) , .ZN( us11_n448 ) , .A1( us11_n847 ) );
  NOR2_X1 us11_U388 (.A2( sa11_2 ) , .A1( sa11_3 ) , .ZN( us11_n472 ) );
  NOR2_X1 us11_U389 (.A2( sa11_0 ) , .ZN( us11_n454 ) , .A1( us11_n827 ) );
  AOI222_X1 us11_U39 (.ZN( us11_n525 ) , .A1( us11_n834 ) , .B2( us11_n837 ) , .C1( us11_n844 ) , .C2( us11_n850 ) , .A2( us11_n852 ) , .B1( us11_n866 ) );
  NOR2_X1 us11_U390 (.A2( sa11_3 ) , .ZN( us11_n455 ) , .A1( us11_n828 ) );
  NOR2_X1 us11_U391 (.A2( sa11_0 ) , .A1( sa11_1 ) , .ZN( us11_n462 ) );
  INV_X1 us11_U392 (.A( sa11_6 ) , .ZN( us11_n849 ) );
  INV_X1 us11_U393 (.A( sa11_1 ) , .ZN( us11_n827 ) );
  INV_X1 us11_U394 (.A( sa11_2 ) , .ZN( us11_n828 ) );
  INV_X1 us11_U395 (.A( sa11_5 ) , .ZN( us11_n848 ) );
  NAND2_X1 us11_U396 (.A2( us11_n461 ) , .A1( us11_n471 ) , .ZN( us11_n697 ) );
  NOR2_X1 us11_U397 (.A2( sa11_6 ) , .ZN( us11_n452 ) , .A1( us11_n858 ) );
  INV_X1 us11_U398 (.A( sa11_7 ) , .ZN( us11_n858 ) );
  NAND2_X1 us11_U399 (.A2( us11_n461 ) , .A1( us11_n462 ) , .ZN( us11_n747 ) );
  NAND2_X2 us11_U4 (.A1( us11_n441 ) , .A2( us11_n464 ) , .ZN( us11_n708 ) );
  NOR4_X1 us11_U40 (.A3( us11_n521 ) , .A1( us11_n522 ) , .ZN( us11_n523 ) , .A2( us11_n673 ) , .A4( us11_n769 ) );
  NAND2_X2 us11_U400 (.A1( us11_n454 ) , .A2( us11_n461 ) , .ZN( us11_n813 ) );
  NOR2_X1 us11_U401 (.A2( sa11_1 ) , .ZN( us11_n471 ) , .A1( us11_n826 ) );
  INV_X1 us11_U402 (.A( sa11_0 ) , .ZN( us11_n826 ) );
  OAI221_X1 us11_U403 (.A( us11_n783 ) , .C2( us11_n784 ) , .B2( us11_n785 ) , .B1( us11_n786 ) , .ZN( us11_n796 ) , .C1( us11_n813 ) );
  NAND2_X1 us11_U404 (.A1( us11_n729 ) , .A2( us11_n784 ) , .ZN( us11_n811 ) );
  OAI22_X1 us11_U405 (.ZN( us11_n588 ) , .A2( us11_n747 ) , .B2( us11_n762 ) , .A1( us11_n763 ) , .B1( us11_n784 ) );
  OAI221_X1 us11_U406 (.A( us11_n696 ) , .ZN( us11_n703 ) , .C2( us11_n784 ) , .C1( us11_n785 ) , .B1( us11_n786 ) , .B2( us11_n806 ) );
  AOI21_X1 us11_U407 (.ZN( us11_n592 ) , .B1( us11_n728 ) , .B2( us11_n784 ) , .A( us11_n790 ) );
  AOI21_X1 us11_U408 (.ZN( us11_n648 ) , .A( us11_n762 ) , .B2( us11_n784 ) , .B1( us11_n792 ) );
  AOI21_X1 us11_U409 (.ZN( us11_n623 ) , .B1( us11_n699 ) , .A( us11_n779 ) , .B2( us11_n784 ) );
  AOI221_X1 us11_U41 (.A( us11_n781 ) , .ZN( us11_n798 ) , .C2( us11_n837 ) , .B2( us11_n838 ) , .B1( us11_n865 ) , .C1( us11_n866 ) );
  OAI22_X1 us11_U410 (.ZN( us11_n681 ) , .A1( us11_n699 ) , .A2( us11_n730 ) , .B2( us11_n784 ) , .B1( us11_n817 ) );
  OAI21_X1 us11_U411 (.A( us11_n613 ) , .ZN( us11_n616 ) , .B1( us11_n625 ) , .B2( us11_n784 ) );
  NOR2_X1 us11_U412 (.ZN( us11_n610 ) , .A1( us11_n784 ) , .A2( us11_n816 ) );
  NOR2_X1 us11_U413 (.ZN( us11_n651 ) , .A1( us11_n784 ) , .A2( us11_n788 ) );
  OAI222_X1 us11_U414 (.A2( us11_n669 ) , .ZN( us11_n674 ) , .B1( us11_n747 ) , .B2( us11_n784 ) , .C2( us11_n788 ) , .C1( us11_n815 ) , .A1( us11_n817 ) );
  NOR2_X1 us11_U415 (.ZN( us11_n600 ) , .A2( us11_n697 ) , .A1( us11_n784 ) );
  NOR2_X1 us11_U416 (.ZN( us11_n553 ) , .A2( us11_n744 ) , .A1( us11_n784 ) );
  INV_X1 us11_U417 (.A( us11_n784 ) , .ZN( us11_n861 ) );
  NAND4_X1 us11_U418 (.ZN( sa10_sr_2 ) , .A4( us11_n643 ) , .A3( us11_n644 ) , .A2( us11_n645 ) , .A1( us11_n646 ) );
  AOI211_X1 us11_U419 (.A( us11_n637 ) , .ZN( us11_n645 ) , .B( us11_n743 ) , .C2( us11_n839 ) , .C1( us11_n854 ) );
  NOR4_X1 us11_U42 (.A4( us11_n793 ) , .A3( us11_n794 ) , .A2( us11_n795 ) , .A1( us11_n796 ) , .ZN( us11_n797 ) );
  NOR4_X1 us11_U420 (.A1( us11_n584 ) , .ZN( us11_n585 ) , .A3( us11_n652 ) , .A2( us11_n662 ) , .A4( us11_n767 ) );
  NOR2_X1 us11_U421 (.A2( sa11_2 ) , .ZN( us11_n461 ) , .A1( us11_n829 ) );
  INV_X1 us11_U422 (.A( sa11_3 ) , .ZN( us11_n829 ) );
  OAI222_X1 us11_U423 (.B2( us11_n747 ) , .B1( us11_n748 ) , .A2( us11_n749 ) , .ZN( us11_n757 ) , .C2( us11_n805 ) , .C1( us11_n814 ) , .A1( us11_n817 ) );
  OAI222_X1 us11_U424 (.ZN( us11_n505 ) , .C2( us11_n625 ) , .B2( us11_n647 ) , .B1( us11_n747 ) , .A2( us11_n748 ) , .C1( us11_n805 ) , .A1( us11_n806 ) );
  AOI222_X1 us11_U425 (.ZN( us11_n605 ) , .B2( us11_n671 ) , .B1( us11_n753 ) , .C2( us11_n831 ) , .A1( us11_n833 ) , .A2( us11_n862 ) , .C1( us11_n863 ) );
  AOI222_X1 us11_U426 (.ZN( us11_n513 ) , .C1( us11_n832 ) , .B2( us11_n837 ) , .A2( us11_n843 ) , .C2( us11_n862 ) , .B1( us11_n863 ) , .A1( us11_n866 ) );
  AOI221_X1 us11_U427 (.A( us11_n483 ) , .ZN( us11_n488 ) , .B1( us11_n831 ) , .C2( us11_n844 ) , .C1( us11_n852 ) , .B2( us11_n862 ) );
  NOR2_X1 us11_U428 (.ZN( us11_n789 ) , .A2( us11_n862 ) , .A1( us11_n868 ) );
  NOR2_X1 us11_U429 (.ZN( us11_n748 ) , .A1( us11_n861 ) , .A2( us11_n862 ) );
  NOR4_X1 us11_U43 (.A4( us11_n776 ) , .A3( us11_n777 ) , .A1( us11_n778 ) , .ZN( us11_n799 ) , .A2( us11_n801 ) );
  NOR2_X1 us11_U430 (.A2( sa11_4 ) , .ZN( us11_n449 ) , .A1( us11_n848 ) );
  NOR2_X1 us11_U431 (.A2( sa11_4 ) , .A1( sa11_5 ) , .ZN( us11_n441 ) );
  INV_X1 us11_U432 (.A( sa11_4 ) , .ZN( us11_n847 ) );
  AND2_X1 us11_U433 (.ZN( us11_n438 ) , .A2( us11_n831 ) , .A1( us11_n854 ) );
  AND2_X1 us11_U434 (.ZN( us11_n439 ) , .A2( us11_n843 ) , .A1( us11_n861 ) );
  NOR3_X1 us11_U435 (.A1( us11_n438 ) , .A2( us11_n439 ) , .A3( us11_n576 ) , .ZN( us11_n587 ) );
  INV_X1 us11_U436 (.A( us11_n812 ) , .ZN( us11_n854 ) );
  NAND3_X1 us11_U437 (.ZN( sa10_sr_6 ) , .A3( us11_n797 ) , .A2( us11_n798 ) , .A1( us11_n799 ) );
  NAND3_X1 us11_U438 (.ZN( sa10_sr_5 ) , .A3( us11_n758 ) , .A2( us11_n759 ) , .A1( us11_n760 ) );
  NAND3_X1 us11_U439 (.ZN( sa10_sr_4 ) , .A3( us11_n738 ) , .A2( us11_n739 ) , .A1( us11_n740 ) );
  NOR4_X1 us11_U44 (.A4( us11_n734 ) , .A3( us11_n735 ) , .A2( us11_n736 ) , .A1( us11_n737 ) , .ZN( us11_n738 ) );
  NAND3_X1 us11_U440 (.A3( us11_n675 ) , .A2( us11_n676 ) , .A1( us11_n677 ) , .ZN( us11_n807 ) );
  NAND3_X1 us11_U441 (.ZN( us11_n638 ) , .A3( us11_n708 ) , .A2( us11_n724 ) , .A1( us11_n792 ) );
  NAND3_X1 us11_U442 (.A3( us11_n618 ) , .A2( us11_n619 ) , .A1( us11_n620 ) , .ZN( us11_n725 ) );
  NAND3_X1 us11_U443 (.A3( us11_n585 ) , .A2( us11_n586 ) , .A1( us11_n587 ) , .ZN( us11_n621 ) );
  NAND3_X1 us11_U444 (.ZN( us11_n565 ) , .A3( us11_n680 ) , .A2( us11_n750 ) , .A1( us11_n785 ) );
  NAND3_X1 us11_U445 (.A3( us11_n523 ) , .A2( us11_n524 ) , .A1( us11_n525 ) , .ZN( us11_n742 ) );
  NAND3_X1 us11_U446 (.A3( us11_n512 ) , .A1( us11_n513 ) , .ZN( us11_n608 ) , .A2( us11_n871 ) );
  NAND3_X1 us11_U447 (.A3( us11_n467 ) , .A2( us11_n468 ) , .A1( us11_n469 ) , .ZN( us11_n777 ) );
  INV_X1 us11_U448 (.A( us11_n803 ) , .ZN( us11_n843 ) );
  AOI21_X1 us11_U449 (.ZN( us11_n576 ) , .B2( us11_n724 ) , .B1( us11_n748 ) , .A( us11_n785 ) );
  AOI211_X1 us11_U45 (.B( us11_n725 ) , .A( us11_n726 ) , .ZN( us11_n739 ) , .C1( us11_n843 ) , .C2( us11_n855 ) );
  NOR3_X1 us11_U46 (.A3( us11_n722 ) , .A1( us11_n723 ) , .ZN( us11_n740 ) , .A2( us11_n741 ) );
  NOR4_X1 us11_U47 (.A3( us11_n755 ) , .A2( us11_n756 ) , .A1( us11_n757 ) , .ZN( us11_n758 ) , .A4( us11_n869 ) );
  AOI211_X1 us11_U48 (.B( us11_n745 ) , .A( us11_n746 ) , .ZN( us11_n759 ) , .C1( us11_n832 ) , .C2( us11_n853 ) );
  NOR3_X1 us11_U49 (.A3( us11_n741 ) , .A2( us11_n742 ) , .A1( us11_n743 ) , .ZN( us11_n760 ) );
  NAND2_X2 us11_U5 (.A2( us11_n441 ) , .A1( us11_n452 ) , .ZN( us11_n791 ) );
  NAND4_X1 us11_U50 (.ZN( sa10_sr_3 ) , .A4( us11_n704 ) , .A3( us11_n705 ) , .A2( us11_n706 ) , .A1( us11_n707 ) );
  NOR4_X1 us11_U51 (.A4( us11_n700 ) , .A3( us11_n701 ) , .A2( us11_n702 ) , .A1( us11_n703 ) , .ZN( us11_n704 ) );
  AOI211_X1 us11_U52 (.B( us11_n694 ) , .A( us11_n695 ) , .ZN( us11_n705 ) , .C2( us11_n831 ) , .C1( us11_n851 ) );
  NOR2_X1 us11_U53 (.ZN( us11_n707 ) , .A2( us11_n776 ) , .A1( us11_n800 ) );
  NOR2_X1 us11_U54 (.ZN( us11_n804 ) , .A1( us11_n854 ) , .A2( us11_n861 ) );
  NAND4_X1 us11_U55 (.ZN( sa10_sr_1 ) , .A4( us11_n595 ) , .A3( us11_n596 ) , .A2( us11_n597 ) , .A1( us11_n598 ) );
  AOI211_X1 us11_U56 (.B( us11_n589 ) , .A( us11_n590 ) , .ZN( us11_n596 ) , .C2( us11_n811 ) , .C1( us11_n833 ) );
  NOR4_X1 us11_U57 (.A4( us11_n591 ) , .A3( us11_n592 ) , .A2( us11_n593 ) , .A1( us11_n594 ) , .ZN( us11_n595 ) );
  AOI211_X1 us11_U58 (.A( us11_n588 ) , .ZN( us11_n597 ) , .B( us11_n621 ) , .C1( us11_n845 ) , .C2( us11_n855 ) );
  NAND4_X1 us11_U59 (.ZN( sa10_sr_0 ) , .A4( us11_n501 ) , .A3( us11_n502 ) , .A2( us11_n503 ) , .A1( us11_n504 ) );
  INV_X1 us11_U6 (.A( us11_n669 ) , .ZN( us11_n865 ) );
  AOI221_X1 us11_U60 (.A( us11_n497 ) , .ZN( us11_n502 ) , .B2( us11_n843 ) , .C1( us11_n846 ) , .C2( us11_n860 ) , .B1( us11_n862 ) );
  NOR4_X1 us11_U61 (.A4( us11_n498 ) , .A3( us11_n499 ) , .A2( us11_n500 ) , .ZN( us11_n501 ) , .A1( us11_n527 ) );
  AOI211_X1 us11_U62 (.A( us11_n496 ) , .ZN( us11_n503 ) , .B( us11_n802 ) , .C2( us11_n839 ) , .C1( us11_n851 ) );
  NAND4_X1 us11_U63 (.ZN( sa10_sr_7 ) , .A4( us11_n822 ) , .A3( us11_n823 ) , .A2( us11_n824 ) , .A1( us11_n825 ) );
  AOI222_X1 us11_U64 (.C2( us11_n809 ) , .B2( us11_n810 ) , .A2( us11_n811 ) , .ZN( us11_n823 ) , .C1( us11_n832 ) , .A1( us11_n839 ) , .B1( us11_n853 ) );
  NOR4_X1 us11_U65 (.A4( us11_n818 ) , .A3( us11_n819 ) , .A2( us11_n820 ) , .A1( us11_n821 ) , .ZN( us11_n822 ) );
  AOI211_X1 us11_U66 (.B( us11_n807 ) , .A( us11_n808 ) , .ZN( us11_n824 ) , .C1( us11_n842 ) , .C2( us11_n850 ) );
  NAND4_X1 us11_U67 (.A4( us11_n603 ) , .A3( us11_n604 ) , .A2( us11_n605 ) , .A1( us11_n606 ) , .ZN( us11_n722 ) );
  NOR3_X1 us11_U68 (.A1( us11_n599 ) , .ZN( us11_n604 ) , .A3( us11_n663 ) , .A2( us11_n770 ) );
  NOR4_X1 us11_U69 (.A3( us11_n600 ) , .A2( us11_n601 ) , .A1( us11_n602 ) , .ZN( us11_n603 ) , .A4( us11_n655 ) );
  NAND2_X1 us11_U7 (.A1( us11_n449 ) , .A2( us11_n464 ) , .ZN( us11_n724 ) );
  AOI222_X1 us11_U70 (.ZN( us11_n606 ) , .A1( us11_n830 ) , .C2( us11_n837 ) , .B1( us11_n842 ) , .A2( us11_n856 ) , .B2( us11_n861 ) , .C1( us11_n868 ) );
  NAND4_X1 us11_U71 (.A4( us11_n485 ) , .A3( us11_n486 ) , .A2( us11_n487 ) , .A1( us11_n488 ) , .ZN( us11_n778 ) );
  NOR4_X1 us11_U72 (.A4( us11_n484 ) , .ZN( us11_n487 ) , .A1( us11_n566 ) , .A2( us11_n581 ) , .A3( us11_n602 ) );
  NOR4_X1 us11_U73 (.ZN( us11_n486 ) , .A1( us11_n507 ) , .A2( us11_n519 ) , .A4( us11_n546 ) , .A3( us11_n611 ) );
  NAND4_X1 us11_U74 (.A4( us11_n657 ) , .A3( us11_n658 ) , .A2( us11_n659 ) , .A1( us11_n660 ) , .ZN( us11_n800 ) );
  NOR3_X1 us11_U75 (.A3( us11_n654 ) , .A2( us11_n655 ) , .A1( us11_n656 ) , .ZN( us11_n657 ) );
  NOR3_X1 us11_U76 (.A3( us11_n651 ) , .A2( us11_n652 ) , .A1( us11_n653 ) , .ZN( us11_n658 ) );
  NOR3_X1 us11_U77 (.A3( us11_n648 ) , .A2( us11_n649 ) , .A1( us11_n650 ) , .ZN( us11_n659 ) );
  NAND4_X1 us11_U78 (.A4( us11_n560 ) , .A3( us11_n561 ) , .A2( us11_n562 ) , .A1( us11_n563 ) , .ZN( us11_n607 ) );
  NOR4_X1 us11_U79 (.ZN( us11_n561 ) , .A1( us11_n653 ) , .A3( us11_n661 ) , .A4( us11_n685 ) , .A2( us11_n768 ) );
  NOR3_X1 us11_U8 (.ZN( us11_n598 ) , .A1( us11_n608 ) , .A3( us11_n723 ) , .A2( us11_n742 ) );
  NOR4_X1 us11_U80 (.A4( us11_n552 ) , .A3( us11_n553 ) , .A2( us11_n554 ) , .A1( us11_n555 ) , .ZN( us11_n562 ) );
  NOR4_X1 us11_U81 (.A4( us11_n556 ) , .A3( us11_n557 ) , .A2( us11_n558 ) , .A1( us11_n559 ) , .ZN( us11_n560 ) );
  NAND4_X1 us11_U82 (.A4( us11_n772 ) , .A3( us11_n773 ) , .A2( us11_n774 ) , .A1( us11_n775 ) , .ZN( us11_n801 ) );
  NOR3_X1 us11_U83 (.A3( us11_n765 ) , .A2( us11_n766 ) , .A1( us11_n767 ) , .ZN( us11_n773 ) );
  NOR4_X1 us11_U84 (.A4( us11_n768 ) , .A3( us11_n769 ) , .A2( us11_n770 ) , .A1( us11_n771 ) , .ZN( us11_n772 ) );
  AOI222_X1 us11_U85 (.ZN( us11_n775 ) , .A1( us11_n830 ) , .C1( us11_n834 ) , .B2( us11_n841 ) , .A2( us11_n850 ) , .B1( us11_n861 ) , .C2( us11_n873 ) );
  NOR4_X1 us11_U86 (.A4( us11_n509 ) , .A2( us11_n510 ) , .A1( us11_n511 ) , .ZN( us11_n512 ) , .A3( us11_n670 ) );
  INV_X1 us11_U87 (.A( us11_n505 ) , .ZN( us11_n871 ) );
  NOR4_X1 us11_U88 (.A4( us11_n665 ) , .A3( us11_n666 ) , .A2( us11_n667 ) , .A1( us11_n668 ) , .ZN( us11_n676 ) );
  NOR4_X1 us11_U89 (.A4( us11_n661 ) , .A3( us11_n662 ) , .A2( us11_n663 ) , .A1( us11_n664 ) , .ZN( us11_n677 ) );
  NOR3_X1 us11_U9 (.A3( us11_n800 ) , .A2( us11_n801 ) , .A1( us11_n802 ) , .ZN( us11_n825 ) );
  NOR4_X1 us11_U90 (.A3( us11_n673 ) , .A1( us11_n674 ) , .ZN( us11_n675 ) , .A4( us11_n715 ) , .A2( us11_n859 ) );
  NOR2_X1 us11_U91 (.ZN( us11_n625 ) , .A2( us11_n836 ) , .A1( us11_n839 ) );
  NOR2_X1 us11_U92 (.ZN( us11_n761 ) , .A1( us11_n833 ) , .A2( us11_n834 ) );
  NAND4_X1 us11_U93 (.A4( us11_n456 ) , .A3( us11_n457 ) , .A2( us11_n458 ) , .A1( us11_n459 ) , .ZN( us11_n679 ) );
  AOI221_X1 us11_U94 (.A( us11_n450 ) , .ZN( us11_n459 ) , .C2( us11_n753 ) , .B1( us11_n832 ) , .C1( us11_n842 ) , .B2( us11_n861 ) );
  NOR3_X1 us11_U95 (.ZN( us11_n457 ) , .A3( us11_n530 ) , .A1( us11_n555 ) , .A2( us11_n570 ) );
  NOR4_X1 us11_U96 (.ZN( us11_n458 ) , .A2( us11_n509 ) , .A1( us11_n599 ) , .A4( us11_n628 ) , .A3( us11_n711 ) );
  NAND4_X1 us11_U97 (.A4( us11_n535 ) , .A3( us11_n536 ) , .A2( us11_n537 ) , .A1( us11_n538 ) , .ZN( us11_n622 ) );
  NOR4_X1 us11_U98 (.A1( us11_n531 ) , .ZN( us11_n536 ) , .A2( us11_n654 ) , .A4( us11_n668 ) , .A3( us11_n765 ) );
  NOR4_X1 us11_U99 (.A4( us11_n526 ) , .A2( us11_n527 ) , .A1( us11_n528 ) , .ZN( us11_n538 ) , .A3( us11_n701 ) );
  NOR2_X1 us22_U10 (.ZN( us22_n573 ) , .A1( us22_n620 ) , .A2( us22_n743 ) );
  NOR4_X1 us22_U100 (.A4( us22_n527 ) , .A3( us22_n528 ) , .ZN( us22_n535 ) , .A2( us22_n682 ) , .A1( us22_n792 ) );
  NAND4_X1 us22_U101 (.A4( us22_n477 ) , .A3( us22_n478 ) , .A2( us22_n479 ) , .A1( us22_n480 ) , .ZN( us22_n692 ) );
  NOR3_X1 us22_U102 (.ZN( us22_n478 ) , .A2( us22_n506 ) , .A3( us22_n599 ) , .A1( us22_n608 ) );
  AOI211_X1 us22_U103 (.B( us22_n475 ) , .A( us22_n476 ) , .ZN( us22_n480 ) , .C2( us22_n831 ) , .C1( us22_n859 ) );
  NOR4_X1 us22_U104 (.ZN( us22_n479 ) , .A3( us22_n530 ) , .A4( us22_n543 ) , .A2( us22_n565 ) , .A1( us22_n715 ) );
  NAND4_X1 us22_U105 (.A4( us22_n546 ) , .A3( us22_n547 ) , .A2( us22_n548 ) , .A1( us22_n549 ) , .ZN( us22_n743 ) );
  NOR3_X1 us22_U106 (.ZN( us22_n547 ) , .A2( us22_n649 ) , .A1( us22_n665 ) , .A3( us22_n769 ) );
  AOI211_X1 us22_U107 (.B( us22_n537 ) , .A( us22_n538 ) , .ZN( us22_n549 ) , .C2( us22_n837 ) , .C1( us22_n849 ) );
  NOR4_X1 us22_U108 (.A4( us22_n542 ) , .A3( us22_n543 ) , .A2( us22_n544 ) , .A1( us22_n545 ) , .ZN( us22_n546 ) );
  NOR2_X1 us22_U109 (.ZN( us22_n684 ) , .A1( us22_n829 ) , .A2( us22_n830 ) );
  NOR2_X1 us22_U11 (.A1( us22_n676 ) , .ZN( us22_n691 ) , .A2( us22_n805 ) );
  NOR4_X1 us22_U110 (.ZN( us22_n618 ) , .A1( us22_n654 ) , .A3( us22_n664 ) , .A4( us22_n680 ) , .A2( us22_n764 ) );
  NOR4_X1 us22_U111 (.A4( us22_n607 ) , .A3( us22_n608 ) , .A2( us22_n609 ) , .A1( us22_n610 ) , .ZN( us22_n617 ) );
  NOR4_X1 us22_U112 (.A4( us22_n612 ) , .A3( us22_n613 ) , .A2( us22_n614 ) , .A1( us22_n615 ) , .ZN( us22_n616 ) );
  NAND4_X1 us22_U113 (.A4( us22_n483 ) , .A3( us22_n484 ) , .A2( us22_n485 ) , .A1( us22_n486 ) , .ZN( us22_n776 ) );
  NOR4_X1 us22_U114 (.A4( us22_n482 ) , .ZN( us22_n485 ) , .A1( us22_n564 ) , .A2( us22_n579 ) , .A3( us22_n600 ) );
  NOR4_X1 us22_U115 (.ZN( us22_n484 ) , .A1( us22_n505 ) , .A2( us22_n517 ) , .A4( us22_n544 ) , .A3( us22_n609 ) );
  NOR4_X1 us22_U116 (.ZN( us22_n483 ) , .A2( us22_n531 ) , .A1( us22_n556 ) , .A3( us22_n629 ) , .A4( us22_n716 ) );
  NAND4_X1 us22_U117 (.A4( us22_n689 ) , .A3( us22_n690 ) , .A1( us22_n691 ) , .ZN( us22_n774 ) , .A2( us22_n870 ) );
  AOI221_X1 us22_U118 (.A( us22_n679 ) , .ZN( us22_n690 ) , .B2( us22_n838 ) , .C1( us22_n840 ) , .C2( us22_n860 ) , .B1( us22_n863 ) );
  INV_X1 us22_U119 (.A( us22_n677 ) , .ZN( us22_n870 ) );
  INV_X1 us22_U12 (.A( us22_n678 ) , .ZN( us22_n838 ) );
  NOR4_X1 us22_U120 (.A4( us22_n685 ) , .A3( us22_n686 ) , .A2( us22_n687 ) , .A1( us22_n688 ) , .ZN( us22_n689 ) );
  NAND4_X1 us22_U121 (.A4( us22_n717 ) , .A3( us22_n718 ) , .A2( us22_n719 ) , .ZN( us22_n739 ) , .A1( us22_n855 ) );
  INV_X1 us22_U122 (.A( us22_n707 ) , .ZN( us22_n855 ) );
  AOI221_X1 us22_U123 (.A( us22_n708 ) , .ZN( us22_n719 ) , .C2( us22_n842 ) , .B2( us22_n843 ) , .C1( us22_n859 ) , .B1( us22_n860 ) );
  NOR4_X1 us22_U124 (.A4( us22_n713 ) , .A3( us22_n714 ) , .A2( us22_n715 ) , .A1( us22_n716 ) , .ZN( us22_n717 ) );
  NAND4_X1 us22_U125 (.A4( us22_n471 ) , .A3( us22_n472 ) , .A2( us22_n473 ) , .A1( us22_n474 ) , .ZN( us22_n676 ) );
  NOR4_X1 us22_U126 (.A4( us22_n468 ) , .ZN( us22_n474 ) , .A3( us22_n554 ) , .A1( us22_n733 ) , .A2( us22_n753 ) );
  NOR4_X1 us22_U127 (.ZN( us22_n473 ) , .A1( us22_n529 ) , .A3( us22_n566 ) , .A4( us22_n598 ) , .A2( us22_n640 ) );
  NOR4_X1 us22_U128 (.ZN( us22_n472 ) , .A1( us22_n504 ) , .A3( us22_n542 ) , .A2( us22_n581 ) , .A4( us22_n714 ) );
  NOR2_X1 us22_U129 (.ZN( us22_n731 ) , .A2( us22_n830 ) , .A1( us22_n843 ) );
  NOR4_X1 us22_U13 (.A4( us22_n443 ) , .A3( us22_n444 ) , .A2( us22_n514 ) , .A1( us22_n539 ) , .ZN( us22_n704 ) );
  NOR2_X1 us22_U130 (.ZN( us22_n787 ) , .A2( us22_n860 ) , .A1( us22_n866 ) );
  NOR2_X1 us22_U131 (.ZN( us22_n645 ) , .A1( us22_n852 ) , .A2( us22_n866 ) );
  NAND4_X1 us22_U132 (.A4( us22_n571 ) , .A3( us22_n572 ) , .A1( us22_n573 ) , .ZN( us22_n721 ) , .A2( us22_n872 ) );
  NOR4_X1 us22_U133 (.A4( us22_n567 ) , .A3( us22_n568 ) , .A2( us22_n569 ) , .A1( us22_n570 ) , .ZN( us22_n571 ) );
  AOI221_X1 us22_U134 (.A( us22_n562 ) , .C2( us22_n563 ) , .ZN( us22_n572 ) , .B2( us22_n843 ) , .B1( us22_n850 ) , .C1( us22_n851 ) );
  INV_X1 us22_U135 (.A( us22_n605 ) , .ZN( us22_n872 ) );
  NAND4_X1 us22_U136 (.A4( us22_n491 ) , .A3( us22_n492 ) , .A1( us22_n493 ) , .ZN( us22_n800 ) , .A2( us22_n865 ) );
  AOI221_X1 us22_U137 (.A( us22_n487 ) , .ZN( us22_n492 ) , .B2( us22_n834 ) , .C2( us22_n839 ) , .C1( us22_n849 ) , .B1( us22_n858 ) );
  INV_X1 us22_U138 (.A( us22_n776 ) , .ZN( us22_n865 ) );
  NOR2_X1 us22_U139 (.ZN( us22_n493 ) , .A1( us22_n676 ) , .A2( us22_n692 ) );
  OR3_X1 us22_U14 (.ZN( us22_n444 ) , .A1( us22_n526 ) , .A3( us22_n575 ) , .A2( us22_n873 ) );
  INV_X1 us22_U140 (.A( us22_n760 ) , .ZN( us22_n828 ) );
  INV_X1 us22_U141 (.A( us22_n461 ) , .ZN( us22_n862 ) );
  OAI21_X1 us22_U142 (.ZN( us22_n461 ) , .B1( us22_n807 ) , .A( us22_n832 ) , .B2( us22_n849 ) );
  OR4_X1 us22_U143 (.A4( us22_n578 ) , .A3( us22_n579 ) , .A2( us22_n580 ) , .A1( us22_n581 ) , .ZN( us22_n582 ) );
  OR4_X1 us22_U144 (.A4( us22_n680 ) , .A3( us22_n681 ) , .A2( us22_n682 ) , .A1( us22_n683 ) , .ZN( us22_n688 ) );
  OR4_X1 us22_U145 (.A4( us22_n564 ) , .A3( us22_n565 ) , .A2( us22_n566 ) , .ZN( us22_n570 ) , .A1( us22_n663 ) );
  OR4_X1 us22_U146 (.A4( us22_n516 ) , .A2( us22_n517 ) , .A1( us22_n518 ) , .ZN( us22_n520 ) , .A3( us22_n819 ) );
  OR4_X1 us22_U147 (.ZN( us22_n464 ) , .A4( us22_n516 ) , .A3( us22_n527 ) , .A2( us22_n576 ) , .A1( us22_n710 ) );
  NAND2_X1 us22_U148 (.ZN( us22_n611 ) , .A2( us22_n835 ) , .A1( us22_n871 ) );
  OR3_X1 us22_U149 (.A3( us22_n504 ) , .A2( us22_n505 ) , .A1( us22_n506 ) , .ZN( us22_n509 ) );
  OR4_X1 us22_U15 (.A4( us22_n440 ) , .A2( us22_n441 ) , .A1( us22_n442 ) , .ZN( us22_n443 ) , .A3( us22_n551 ) );
  AOI221_X1 us22_U150 (.A( us22_n711 ) , .B2( us22_n712 ) , .ZN( us22_n718 ) , .C1( us22_n830 ) , .B1( us22_n837 ) , .C2( us22_n861 ) );
  OR2_X1 us22_U151 (.A2( us22_n709 ) , .A1( us22_n710 ) , .ZN( us22_n711 ) );
  INV_X1 us22_U152 (.A( us22_n752 ) , .ZN( us22_n867 ) );
  OAI21_X1 us22_U153 (.B1( us22_n751 ) , .ZN( us22_n752 ) , .A( us22_n843 ) , .B2( us22_n866 ) );
  INV_X1 us22_U154 (.A( us22_n670 ) , .ZN( us22_n857 ) );
  AOI21_X1 us22_U155 (.A( us22_n668 ) , .B1( us22_n669 ) , .ZN( us22_n670 ) , .B2( us22_n854 ) );
  NAND2_X1 us22_U156 (.A1( us22_n445 ) , .A2( us22_n463 ) , .ZN( us22_n747 ) );
  OAI222_X1 us22_U157 (.B2( us22_n745 ) , .B1( us22_n746 ) , .A2( us22_n747 ) , .ZN( us22_n755 ) , .C2( us22_n803 ) , .C1( us22_n812 ) , .A1( us22_n815 ) );
  OAI222_X1 us22_U158 (.B2( us22_n706 ) , .ZN( us22_n707 ) , .C2( us22_n722 ) , .B1( us22_n745 ) , .A1( us22_n804 ) , .C1( us22_n812 ) , .A2( us22_n813 ) );
  OAI222_X1 us22_U159 (.ZN( us22_n615 ) , .B1( us22_n695 ) , .C1( us22_n722 ) , .C2( us22_n745 ) , .B2( us22_n784 ) , .A2( us22_n790 ) , .A1( us22_n814 ) );
  INV_X1 us22_U16 (.A( us22_n611 ) , .ZN( us22_n873 ) );
  OAI222_X1 us22_U160 (.ZN( us22_n503 ) , .C2( us22_n623 ) , .B2( us22_n645 ) , .B1( us22_n745 ) , .A2( us22_n746 ) , .C1( us22_n803 ) , .A1( us22_n804 ) );
  NOR4_X1 us22_U161 (.A2( us22_n489 ) , .A1( us22_n490 ) , .ZN( us22_n491 ) , .A3( us22_n578 ) , .A4( us22_n610 ) );
  OR4_X1 us22_U162 (.ZN( us22_n490 ) , .A4( us22_n532 ) , .A2( us22_n545 ) , .A1( us22_n557 ) , .A3( us22_n630 ) );
  OAI22_X1 us22_U163 (.B1( us22_n488 ) , .ZN( us22_n489 ) , .A1( us22_n684 ) , .A2( us22_n761 ) , .B2( us22_n815 ) );
  NOR3_X1 us22_U164 (.ZN( us22_n488 ) , .A1( us22_n780 ) , .A2( us22_n848 ) , .A3( us22_n861 ) );
  AOI22_X1 us22_U165 (.ZN( us22_n694 ) , .A1( us22_n828 ) , .B2( us22_n841 ) , .A2( us22_n863 ) , .B1( us22_n866 ) );
  AOI22_X1 us22_U166 (.A2( us22_n780 ) , .ZN( us22_n781 ) , .B2( us22_n829 ) , .A1( us22_n832 ) , .B1( us22_n861 ) );
  INV_X1 us22_U167 (.A( us22_n728 ) , .ZN( us22_n837 ) );
  AOI221_X1 us22_U168 (.A( us22_n481 ) , .ZN( us22_n486 ) , .B1( us22_n829 ) , .C2( us22_n842 ) , .C1( us22_n850 ) , .B2( us22_n860 ) );
  OAI22_X1 us22_U169 (.ZN( us22_n481 ) , .A1( us22_n706 ) , .B2( us22_n783 ) , .A2( us22_n804 ) , .B1( us22_n810 ) );
  INV_X1 us22_U17 (.A( us22_n747 ) , .ZN( us22_n861 ) );
  INV_X1 us22_U170 (.A( us22_n788 ) , .ZN( us22_n830 ) );
  NAND2_X1 us22_U171 (.A1( us22_n449 ) , .A2( us22_n451 ) , .ZN( us22_n760 ) );
  OAI22_X1 us22_U172 (.ZN( us22_n635 ) , .A1( us22_n697 ) , .B2( us22_n726 ) , .A2( us22_n760 ) , .B1( us22_n814 ) );
  OAI221_X1 us22_U173 (.A( us22_n725 ) , .C2( us22_n726 ) , .B2( us22_n727 ) , .B1( us22_n728 ) , .ZN( us22_n735 ) , .C1( us22_n815 ) );
  AOI22_X1 us22_U174 (.ZN( us22_n725 ) , .B1( us22_n830 ) , .A2( us22_n836 ) , .A1( us22_n861 ) , .B2( us22_n864 ) );
  OAI22_X1 us22_U175 (.ZN( us22_n708 ) , .A2( us22_n726 ) , .B2( us22_n727 ) , .A1( us22_n742 ) , .B1( us22_n811 ) );
  INV_X1 us22_U176 (.A( us22_n814 ) , .ZN( us22_n829 ) );
  OAI22_X1 us22_U177 (.ZN( us22_n487 ) , .A1( us22_n722 ) , .B2( us22_n726 ) , .B1( us22_n728 ) , .A2( us22_n777 ) );
  OAI22_X1 us22_U178 (.ZN( us22_n622 ) , .B1( us22_n667 ) , .B2( us22_n745 ) , .A1( us22_n813 ) , .A2( us22_n814 ) );
  INV_X1 us22_U179 (.A( us22_n742 ) , .ZN( us22_n835 ) );
  AOI222_X1 us22_U18 (.ZN( us22_n603 ) , .B2( us22_n669 ) , .B1( us22_n751 ) , .C2( us22_n829 ) , .A1( us22_n831 ) , .A2( us22_n860 ) , .C1( us22_n861 ) );
  OAI22_X1 us22_U180 (.A1( us22_n722 ) , .ZN( us22_n724 ) , .B2( us22_n748 ) , .B1( us22_n810 ) , .A2( us22_n814 ) );
  OAI22_X1 us22_U181 (.B2( us22_n777 ) , .B1( us22_n778 ) , .ZN( us22_n779 ) , .A2( us22_n812 ) , .A1( us22_n813 ) );
  INV_X1 us22_U182 (.A( us22_n786 ) , .ZN( us22_n843 ) );
  INV_X1 us22_U183 (.A( us22_n812 ) , .ZN( us22_n831 ) );
  OAI22_X1 us22_U184 (.B2( us22_n742 ) , .ZN( us22_n744 ) , .A2( us22_n760 ) , .B1( us22_n778 ) , .A1( us22_n790 ) );
  OAI22_X1 us22_U185 (.B2( us22_n801 ) , .B1( us22_n802 ) , .A2( us22_n803 ) , .A1( us22_n804 ) , .ZN( us22_n806 ) );
  INV_X1 us22_U186 (.A( us22_n667 ) , .ZN( us22_n863 ) );
  OAI22_X1 us22_U187 (.ZN( us22_n494 ) , .A2( us22_n742 ) , .A1( us22_n778 ) , .B1( us22_n789 ) , .B2( us22_n804 ) );
  INV_X1 us22_U188 (.A( us22_n748 ) , .ZN( us22_n840 ) );
  OAI22_X1 us22_U189 (.ZN( us22_n588 ) , .B1( us22_n728 ) , .B2( us22_n747 ) , .A2( us22_n784 ) , .A1( us22_n801 ) );
  AOI222_X1 us22_U19 (.ZN( us22_n561 ) , .B1( us22_n828 ) , .C1( us22_n839 ) , .A2( us22_n841 ) , .A1( us22_n852 ) , .B2( us22_n861 ) , .C2( us22_n871 ) );
  OAI22_X1 us22_U190 (.ZN( us22_n693 ) , .A2( us22_n728 ) , .A1( us22_n778 ) , .B1( us22_n789 ) , .B2( us22_n815 ) );
  INV_X1 us22_U191 (.A( us22_n801 ) , .ZN( us22_n841 ) );
  NOR2_X1 us22_U192 (.A1( us22_n695 ) , .ZN( us22_n768 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U193 (.ZN( us22_n664 ) , .A1( us22_n726 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U194 (.ZN( us22_n592 ) , .A2( us22_n695 ) , .A1( us22_n726 ) );
  NOR2_X1 us22_U195 (.ZN( us22_n568 ) , .A1( us22_n726 ) , .A2( us22_n804 ) );
  NOR2_X1 us22_U196 (.ZN( us22_n716 ) , .A2( us22_n722 ) , .A1( us22_n742 ) );
  NOR2_X1 us22_U197 (.ZN( us22_n544 ) , .A2( us22_n778 ) , .A1( us22_n812 ) );
  NOR2_X1 us22_U198 (.ZN( us22_n575 ) , .A2( us22_n697 ) , .A1( us22_n812 ) );
  NOR2_X1 us22_U199 (.ZN( us22_n652 ) , .A1( us22_n726 ) , .A2( us22_n811 ) );
  AOI222_X1 us22_U20 (.ZN( us22_n658 ) , .A2( us22_n837 ) , .B1( us22_n839 ) , .C2( us22_n843 ) , .A1( us22_n858 ) , .C1( us22_n861 ) , .B2( us22_n868 ) );
  NOR2_X1 us22_U200 (.ZN( us22_n610 ) , .A1( us22_n777 ) , .A2( us22_n784 ) );
  NOR2_X1 us22_U201 (.ZN( us22_n530 ) , .A2( us22_n747 ) , .A1( us22_n748 ) );
  NOR2_X1 us22_U202 (.ZN( us22_n627 ) , .A2( us22_n726 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U203 (.ZN( us22_n613 ) , .A1( us22_n783 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U204 (.ZN( us22_n599 ) , .A2( us22_n778 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U205 (.ZN( us22_n609 ) , .A2( us22_n778 ) , .A1( us22_n804 ) );
  INV_X1 us22_U206 (.A( us22_n745 ) , .ZN( us22_n832 ) );
  NOR2_X1 us22_U207 (.A2( us22_n742 ) , .ZN( us22_n767 ) , .A1( us22_n810 ) );
  NOR2_X1 us22_U208 (.ZN( us22_n526 ) , .A2( us22_n722 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U209 (.ZN( us22_n529 ) , .A2( us22_n778 ) , .A1( us22_n814 ) );
  INV_X1 us22_U21 (.A( us22_n645 ) , .ZN( us22_n868 ) );
  NOR2_X1 us22_U210 (.ZN( us22_n626 ) , .A2( us22_n667 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U211 (.ZN( us22_n597 ) , .A2( us22_n789 ) , .A1( us22_n814 ) );
  INV_X1 us22_U212 (.A( us22_n790 ) , .ZN( us22_n849 ) );
  INV_X1 us22_U213 (.A( us22_n726 ) , .ZN( us22_n850 ) );
  NOR2_X1 us22_U214 (.ZN( us22_n650 ) , .A1( us22_n667 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U215 (.A1( us22_n667 ) , .ZN( us22_n671 ) , .A2( us22_n742 ) );
  INV_X1 us22_U216 (.A( us22_n803 ) , .ZN( us22_n858 ) );
  NOR2_X1 us22_U217 (.ZN( us22_n600 ) , .A1( us22_n667 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U218 (.A1( us22_n667 ) , .ZN( us22_n686 ) , .A2( us22_n814 ) );
  NOR2_X1 us22_U219 (.A2( us22_n706 ) , .A1( us22_n748 ) , .ZN( us22_n769 ) );
  NOR4_X1 us22_U22 (.ZN( us22_n471 ) , .A2( us22_n519 ) , .A4( us22_n592 ) , .A1( us22_n607 ) , .A3( us22_n627 ) );
  NOR2_X1 us22_U220 (.A1( us22_n667 ) , .ZN( us22_n764 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U221 (.A1( us22_n697 ) , .ZN( us22_n766 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U222 (.ZN( us22_n539 ) , .A2( us22_n695 ) , .A1( us22_n697 ) );
  NOR2_X1 us22_U223 (.ZN( us22_n525 ) , .A1( us22_n667 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U224 (.ZN( us22_n665 ) , .A1( us22_n748 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U225 (.ZN( us22_n553 ) , .A1( us22_n748 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U226 (.ZN( us22_n506 ) , .A2( us22_n778 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U227 (.ZN( us22_n541 ) , .A2( us22_n706 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U228 (.ZN( us22_n662 ) , .A1( us22_n783 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U229 (.A2( us22_n695 ) , .ZN( us22_n714 ) , .A1( us22_n790 ) );
  NOR4_X1 us22_U23 (.ZN( us22_n477 ) , .A1( us22_n518 ) , .A4( us22_n555 ) , .A3( us22_n580 ) , .A2( us22_n628 ) );
  NOR2_X1 us22_U230 (.ZN( us22_n505 ) , .A1( us22_n810 ) , .A2( us22_n815 ) );
  INV_X1 us22_U231 (.A( us22_n804 ) , .ZN( us22_n839 ) );
  NOR2_X1 us22_U232 (.ZN( us22_n659 ) , .A1( us22_n727 ) , .A2( us22_n788 ) );
  NOR2_X1 us22_U233 (.ZN( us22_n660 ) , .A2( us22_n695 ) , .A1( us22_n727 ) );
  NOR2_X1 us22_U234 (.ZN( us22_n555 ) , .A1( us22_n790 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U235 (.ZN( us22_n543 ) , .A1( us22_n747 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U236 (.ZN( us22_n507 ) , .A1( us22_n727 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U237 (.A2( us22_n695 ) , .A1( us22_n778 ) , .ZN( us22_n818 ) );
  OAI22_X1 us22_U238 (.B2( us22_n748 ) , .B1( us22_n749 ) , .A1( us22_n750 ) , .ZN( us22_n754 ) , .A2( us22_n804 ) );
  NOR2_X1 us22_U239 (.ZN( us22_n749 ) , .A2( us22_n850 ) , .A1( us22_n858 ) );
  NOR4_X1 us22_U24 (.ZN( us22_n454 ) , .A2( us22_n515 ) , .A1( us22_n541 ) , .A3( us22_n577 ) , .A4( us22_n613 ) );
  NOR3_X1 us22_U240 (.ZN( us22_n750 ) , .A2( us22_n851 ) , .A1( us22_n861 ) , .A3( us22_n863 ) );
  NOR2_X1 us22_U241 (.ZN( us22_n528 ) , .A2( us22_n742 ) , .A1( us22_n790 ) );
  NOR2_X1 us22_U242 (.A1( us22_n747 ) , .ZN( us22_n765 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U243 (.A2( us22_n742 ) , .ZN( us22_n753 ) , .A1( us22_n803 ) );
  NOR2_X1 us22_U244 (.ZN( us22_n542 ) , .A2( us22_n783 ) , .A1( us22_n790 ) );
  NOR2_X1 us22_U245 (.ZN( us22_n661 ) , .A1( us22_n727 ) , .A2( us22_n783 ) );
  NOR2_X1 us22_U246 (.ZN( us22_n629 ) , .A1( us22_n722 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U247 (.ZN( us22_n733 ) , .A2( us22_n801 ) , .A1( us22_n803 ) );
  NOR2_X1 us22_U248 (.ZN( us22_n612 ) , .A1( us22_n760 ) , .A2( us22_n810 ) );
  OAI22_X1 us22_U249 (.B1( us22_n438 ) , .ZN( us22_n442 ) , .A2( us22_n726 ) , .A1( us22_n742 ) , .B2( us22_n747 ) );
  NOR4_X1 us22_U25 (.A4( us22_n530 ) , .A3( us22_n531 ) , .A2( us22_n532 ) , .ZN( us22_n533 ) , .A1( us22_n818 ) );
  NOR3_X1 us22_U250 (.ZN( us22_n438 ) , .A2( us22_n834 ) , .A3( us22_n835 ) , .A1( us22_n844 ) );
  NOR2_X1 us22_U251 (.ZN( us22_n504 ) , .A2( us22_n726 ) , .A1( us22_n760 ) );
  NOR2_X1 us22_U252 (.ZN( us22_n514 ) , .A1( us22_n706 ) , .A2( us22_n742 ) );
  NOR2_X1 us22_U253 (.ZN( us22_n715 ) , .A2( us22_n742 ) , .A1( us22_n784 ) );
  NOR2_X1 us22_U254 (.ZN( us22_n552 ) , .A1( us22_n784 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U255 (.ZN( us22_n515 ) , .A1( us22_n706 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U256 (.ZN( us22_n556 ) , .A1( us22_n706 ) , .A2( us22_n814 ) );
  NOR2_X1 us22_U257 (.ZN( us22_n519 ) , .A1( us22_n788 ) , .A2( us22_n810 ) );
  NOR2_X1 us22_U258 (.ZN( us22_n628 ) , .A1( us22_n745 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U259 (.ZN( us22_n713 ) , .A1( us22_n803 ) , .A2( us22_n815 ) );
  NOR4_X1 us22_U26 (.A4( us22_n539 ) , .A3( us22_n540 ) , .A2( us22_n541 ) , .ZN( us22_n548 ) , .A1( us22_n686 ) );
  AOI21_X1 us22_U260 (.ZN( us22_n569 ) , .B2( us22_n695 ) , .B1( us22_n804 ) , .A( us22_n810 ) );
  INV_X1 us22_U261 (.A( us22_n761 ) , .ZN( us22_n864 ) );
  NOR2_X1 us22_U262 (.ZN( us22_n653 ) , .A1( us22_n788 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U263 (.ZN( us22_n666 ) , .A2( us22_n706 ) , .A1( us22_n788 ) );
  NOR2_X1 us22_U264 (.ZN( us22_n654 ) , .A1( us22_n745 ) , .A2( us22_n778 ) );
  NOR2_X1 us22_U265 (.ZN( us22_n554 ) , .A1( us22_n760 ) , .A2( us22_n803 ) );
  NOR2_X1 us22_U266 (.ZN( us22_n540 ) , .A1( us22_n760 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U267 (.ZN( us22_n699 ) , .A2( us22_n784 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U268 (.ZN( us22_n607 ) , .A2( us22_n722 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U269 (.A1( us22_n728 ) , .ZN( us22_n763 ) , .A2( us22_n784 ) );
  NOR2_X1 us22_U27 (.ZN( us22_n678 ) , .A2( us22_n832 ) , .A1( us22_n837 ) );
  AOI21_X1 us22_U270 (.A( us22_n813 ) , .B2( us22_n814 ) , .B1( us22_n815 ) , .ZN( us22_n816 ) );
  INV_X1 us22_U271 (.A( us22_n727 ) , .ZN( us22_n866 ) );
  NOR2_X1 us22_U272 (.ZN( us22_n577 ) , .A2( us22_n706 ) , .A1( us22_n728 ) );
  NOR2_X1 us22_U273 (.ZN( us22_n531 ) , .A2( us22_n722 ) , .A1( us22_n728 ) );
  AOI21_X1 us22_U274 (.B1( us22_n623 ) , .ZN( us22_n625 ) , .A( us22_n761 ) , .B2( us22_n812 ) );
  AOI21_X1 us22_U275 (.A( us22_n810 ) , .B2( us22_n811 ) , .B1( us22_n812 ) , .ZN( us22_n817 ) );
  AOI21_X1 us22_U276 (.ZN( us22_n513 ) , .A( us22_n727 ) , .B1( us22_n748 ) , .B2( us22_n801 ) );
  AOI21_X1 us22_U277 (.ZN( us22_n497 ) , .B1( us22_n678 ) , .A( us22_n810 ) , .B2( us22_n814 ) );
  AOI21_X1 us22_U278 (.ZN( us22_n476 ) , .B2( us22_n695 ) , .A( us22_n747 ) , .B1( us22_n777 ) );
  NOR2_X1 us22_U279 (.ZN( us22_n580 ) , .A1( us22_n742 ) , .A2( us22_n813 ) );
  NOR4_X1 us22_U28 (.A4( us22_n512 ) , .A3( us22_n513 ) , .A2( us22_n514 ) , .A1( us22_n515 ) , .ZN( us22_n522 ) );
  NOR2_X1 us22_U280 (.ZN( us22_n640 ) , .A2( us22_n786 ) , .A1( us22_n789 ) );
  AOI21_X1 us22_U281 (.ZN( us22_n591 ) , .B1( us22_n748 ) , .A( us22_n790 ) , .B2( us22_n811 ) );
  NOR2_X1 us22_U282 (.A2( us22_n706 ) , .A1( us22_n760 ) , .ZN( us22_n792 ) );
  AOI21_X1 us22_U283 (.ZN( us22_n624 ) , .B2( us22_n667 ) , .A( us22_n788 ) , .B1( us22_n789 ) );
  NOR2_X1 us22_U284 (.ZN( us22_n668 ) , .A1( us22_n788 ) , .A2( us22_n803 ) );
  NOR2_X1 us22_U285 (.ZN( us22_n518 ) , .A2( us22_n706 ) , .A1( us22_n812 ) );
  AOI21_X1 us22_U286 (.ZN( us22_n475 ) , .A( us22_n667 ) , .B1( us22_n748 ) , .B2( us22_n804 ) );
  NOR2_X1 us22_U287 (.ZN( us22_n557 ) , .A2( us22_n789 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U288 (.ZN( us22_n517 ) , .A2( us22_n697 ) , .A1( us22_n814 ) );
  NOR2_X1 us22_U289 (.ZN( us22_n681 ) , .A2( us22_n697 ) , .A1( us22_n801 ) );
  AOI222_X1 us22_U29 (.ZN( us22_n523 ) , .A1( us22_n832 ) , .B2( us22_n835 ) , .C1( us22_n842 ) , .C2( us22_n848 ) , .A2( us22_n850 ) , .B1( us22_n864 ) );
  NOR2_X1 us22_U290 (.ZN( us22_n651 ) , .A1( us22_n760 ) , .A2( us22_n784 ) );
  INV_X1 us22_U291 (.A( us22_n811 ) , .ZN( us22_n834 ) );
  AOI21_X1 us22_U292 (.ZN( us22_n508 ) , .B2( us22_n667 ) , .A( us22_n728 ) , .B1( us22_n813 ) );
  AOI21_X1 us22_U293 (.ZN( us22_n537 ) , .B2( us22_n810 ) , .A( us22_n812 ) , .B1( us22_n813 ) );
  AOI21_X1 us22_U294 (.ZN( us22_n538 ) , .A( us22_n761 ) , .B2( us22_n777 ) , .B1( us22_n815 ) );
  NOR2_X1 us22_U295 (.ZN( us22_n579 ) , .A1( us22_n667 ) , .A2( us22_n786 ) );
  AOI21_X1 us22_U296 (.ZN( us22_n587 ) , .B2( us22_n697 ) , .B1( us22_n813 ) , .A( us22_n815 ) );
  AOI21_X1 us22_U297 (.B1( us22_n697 ) , .ZN( us22_n698 ) , .A( us22_n730 ) , .B2( us22_n761 ) );
  AOI21_X1 us22_U298 (.ZN( us22_n589 ) , .B2( us22_n761 ) , .A( us22_n783 ) , .B1( us22_n810 ) );
  AOI21_X1 us22_U299 (.ZN( us22_n496 ) , .A( us22_n722 ) , .B2( us22_n760 ) , .B1( us22_n812 ) );
  NAND2_X2 us22_U3 (.A1( us22_n445 ) , .A2( us22_n446 ) , .ZN( us22_n784 ) );
  NOR4_X1 us22_U30 (.A3( us22_n519 ) , .A1( us22_n520 ) , .ZN( us22_n521 ) , .A2( us22_n671 ) , .A4( us22_n767 ) );
  AOI21_X1 us22_U300 (.ZN( us22_n550 ) , .B1( us22_n667 ) , .A( us22_n695 ) , .B2( us22_n803 ) );
  NOR2_X1 us22_U301 (.ZN( us22_n545 ) , .A1( us22_n697 ) , .A2( us22_n742 ) );
  INV_X1 us22_U302 (.A( us22_n789 ) , .ZN( us22_n871 ) );
  INV_X1 us22_U303 (.A( us22_n810 ) , .ZN( us22_n852 ) );
  AOI21_X1 us22_U304 (.ZN( us22_n638 ) , .B2( us22_n745 ) , .A( us22_n790 ) , .B1( us22_n801 ) );
  AOI21_X1 us22_U305 (.ZN( us22_n647 ) , .B1( us22_n727 ) , .B2( us22_n761 ) , .A( us22_n811 ) );
  NOR2_X1 us22_U306 (.ZN( us22_n683 ) , .A1( us22_n727 ) , .A2( us22_n814 ) );
  AOI21_X1 us22_U307 (.B1( us22_n684 ) , .ZN( us22_n685 ) , .A( us22_n726 ) , .B2( us22_n759 ) );
  AOI21_X1 us22_U308 (.ZN( us22_n567 ) , .B1( us22_n748 ) , .B2( us22_n760 ) , .A( us22_n778 ) );
  AOI21_X1 us22_U309 (.ZN( us22_n498 ) , .A( us22_n695 ) , .B1( us22_n706 ) , .B2( us22_n784 ) );
  AOI221_X1 us22_U31 (.A( us22_n779 ) , .ZN( us22_n796 ) , .C2( us22_n835 ) , .B2( us22_n836 ) , .B1( us22_n863 ) , .C1( us22_n864 ) );
  NOR2_X1 us22_U310 (.ZN( us22_n566 ) , .A1( us22_n727 ) , .A2( us22_n760 ) );
  AOI21_X1 us22_U311 (.ZN( us22_n637 ) , .B2( us22_n747 ) , .A( us22_n786 ) , .B1( us22_n810 ) );
  NOR2_X1 us22_U312 (.ZN( us22_n564 ) , .A2( us22_n695 ) , .A1( us22_n761 ) );
  NOR2_X1 us22_U313 (.ZN( us22_n578 ) , .A2( us22_n695 ) , .A1( us22_n789 ) );
  AOI21_X1 us22_U314 (.ZN( us22_n512 ) , .A( us22_n777 ) , .B2( us22_n790 ) , .B1( us22_n810 ) );
  INV_X1 us22_U315 (.A( us22_n697 ) , .ZN( us22_n851 ) );
  NOR2_X1 us22_U316 (.ZN( us22_n663 ) , .A1( us22_n778 ) , .A2( us22_n811 ) );
  AOI21_X1 us22_U317 (.ZN( us22_n448 ) , .B2( us22_n790 ) , .A( us22_n801 ) , .B1( us22_n813 ) );
  NOR2_X1 us22_U318 (.ZN( us22_n630 ) , .A2( us22_n695 ) , .A1( us22_n722 ) );
  AOI21_X1 us22_U319 (.ZN( us22_n562 ) , .B1( us22_n722 ) , .A( us22_n777 ) , .B2( us22_n789 ) );
  NOR4_X1 us22_U32 (.A4( us22_n791 ) , .A3( us22_n792 ) , .A2( us22_n793 ) , .A1( us22_n794 ) , .ZN( us22_n795 ) );
  AOI21_X1 us22_U320 (.ZN( us22_n495 ) , .A( us22_n777 ) , .B2( us22_n789 ) , .B1( us22_n802 ) );
  AOI21_X1 us22_U321 (.ZN( us22_n687 ) , .B2( us22_n747 ) , .B1( us22_n761 ) , .A( us22_n804 ) );
  NOR2_X1 us22_U322 (.ZN( us22_n527 ) , .A1( us22_n706 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U323 (.ZN( us22_n576 ) , .A1( us22_n706 ) , .A2( us22_n811 ) );
  AOI21_X1 us22_U324 (.ZN( us22_n648 ) , .A( us22_n777 ) , .B1( us22_n790 ) , .B2( us22_n803 ) );
  NOR2_X1 us22_U325 (.ZN( us22_n682 ) , .A1( us22_n789 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U326 (.A2( us22_n811 ) , .A1( us22_n813 ) , .ZN( us22_n819 ) );
  AOI21_X1 us22_U327 (.A( us22_n788 ) , .B2( us22_n789 ) , .B1( us22_n790 ) , .ZN( us22_n791 ) );
  AOI21_X1 us22_U328 (.A( us22_n731 ) , .ZN( us22_n732 ) , .B2( us22_n778 ) , .B1( us22_n790 ) );
  NOR2_X1 us22_U329 (.ZN( us22_n565 ) , .A1( us22_n745 ) , .A2( us22_n803 ) );
  NOR4_X1 us22_U33 (.A4( us22_n774 ) , .A3( us22_n775 ) , .A1( us22_n776 ) , .ZN( us22_n797 ) , .A2( us22_n799 ) );
  NOR2_X1 us22_U330 (.ZN( us22_n581 ) , .A1( us22_n790 ) , .A2( us22_n815 ) );
  NOR2_X1 us22_U331 (.ZN( us22_n532 ) , .A1( us22_n722 ) , .A2( us22_n786 ) );
  AOI21_X1 us22_U332 (.ZN( us22_n639 ) , .B1( us22_n678 ) , .A( us22_n789 ) , .B2( us22_n815 ) );
  NOR2_X1 us22_U333 (.ZN( us22_n709 ) , .A1( us22_n760 ) , .A2( us22_n761 ) );
  NOR2_X1 us22_U334 (.ZN( us22_n680 ) , .A2( us22_n706 ) , .A1( us22_n815 ) );
  INV_X1 us22_U335 (.A( us22_n695 ) , .ZN( us22_n836 ) );
  INV_X1 us22_U336 (.A( us22_n813 ) , .ZN( us22_n853 ) );
  AOI21_X1 us22_U337 (.ZN( us22_n440 ) , .A( us22_n697 ) , .B1( us22_n731 ) , .B2( us22_n748 ) );
  OAI21_X1 us22_U338 (.A( us22_n696 ) , .ZN( us22_n700 ) , .B2( us22_n748 ) , .B1( us22_n802 ) );
  OAI21_X1 us22_U339 (.ZN( us22_n696 ) , .B2( us22_n831 ) , .B1( us22_n836 ) , .A( us22_n858 ) );
  NOR4_X1 us22_U34 (.A3( us22_n753 ) , .A2( us22_n754 ) , .A1( us22_n755 ) , .ZN( us22_n756 ) , .A4( us22_n867 ) );
  NAND2_X1 us22_U340 (.ZN( us22_n751 ) , .A1( us22_n761 ) , .A2( us22_n803 ) );
  INV_X1 us22_U341 (.A( us22_n778 ) , .ZN( us22_n848 ) );
  INV_X1 us22_U342 (.A( us22_n783 ) , .ZN( us22_n844 ) );
  NAND2_X1 us22_U343 (.ZN( us22_n669 ) , .A1( us22_n804 ) , .A2( us22_n814 ) );
  NAND2_X1 us22_U344 (.ZN( us22_n712 ) , .A1( us22_n726 ) , .A2( us22_n778 ) );
  NAND2_X1 us22_U345 (.A2( us22_n760 ) , .A1( us22_n804 ) , .ZN( us22_n808 ) );
  NAND2_X2 us22_U346 (.A2( us22_n439 ) , .A1( us22_n445 ) , .ZN( us22_n782 ) );
  AOI21_X1 us22_U347 (.ZN( us22_n441 ) , .B1( us22_n787 ) , .B2( us22_n789 ) , .A( us22_n812 ) );
  NOR2_X1 us22_U348 (.ZN( us22_n468 ) , .A2( us22_n777 ) , .A1( us22_n813 ) );
  OAI21_X1 us22_U349 (.A( us22_n785 ) , .B2( us22_n786 ) , .B1( us22_n787 ) , .ZN( us22_n793 ) );
  AOI211_X1 us22_U35 (.B( us22_n743 ) , .A( us22_n744 ) , .ZN( us22_n757 ) , .C1( us22_n830 ) , .C2( us22_n851 ) );
  OAI21_X1 us22_U350 (.ZN( us22_n785 ) , .A( us22_n837 ) , .B1( us22_n861 ) , .B2( us22_n871 ) );
  NOR2_X1 us22_U351 (.ZN( us22_n524 ) , .A1( us22_n722 ) , .A2( us22_n748 ) );
  NOR2_X1 us22_U352 (.ZN( us22_n710 ) , .A2( us22_n722 ) , .A1( us22_n788 ) );
  NOR2_X1 us22_U353 (.ZN( us22_n482 ) , .A1( us22_n786 ) , .A2( us22_n803 ) );
  NAND2_X1 us22_U354 (.A1( us22_n697 ) , .A2( us22_n727 ) , .ZN( us22_n780 ) );
  NOR2_X1 us22_U355 (.ZN( us22_n516 ) , .A1( us22_n706 ) , .A2( us22_n786 ) );
  NAND2_X1 us22_U356 (.A2( us22_n747 ) , .A1( us22_n784 ) , .ZN( us22_n807 ) );
  OAI21_X1 us22_U357 (.A( us22_n729 ) , .B1( us22_n730 ) , .ZN( us22_n734 ) , .B2( us22_n803 ) );
  OAI21_X1 us22_U358 (.ZN( us22_n729 ) , .A( us22_n831 ) , .B2( us22_n850 ) , .B1( us22_n871 ) );
  INV_X1 us22_U359 (.A( us22_n815 ) , .ZN( us22_n842 ) );
  NOR3_X1 us22_U36 (.A3( us22_n739 ) , .A2( us22_n740 ) , .A1( us22_n741 ) , .ZN( us22_n758 ) );
  INV_X1 us22_U360 (.A( us22_n722 ) , .ZN( us22_n854 ) );
  AND2_X1 us22_U361 (.ZN( us22_n730 ) , .A1( us22_n777 ) , .A2( us22_n783 ) );
  AOI221_X1 us22_U362 (.A( us22_n762 ) , .ZN( us22_n772 ) , .C2( us22_n808 ) , .B2( us22_n833 ) , .C1( us22_n853 ) , .B1( us22_n864 ) );
  AOI21_X1 us22_U363 (.B2( us22_n761 ) , .ZN( us22_n762 ) , .A( us22_n786 ) , .B1( us22_n790 ) );
  INV_X1 us22_U364 (.A( us22_n759 ) , .ZN( us22_n833 ) );
  NAND2_X1 us22_U365 (.A1( us22_n453 ) , .A2( us22_n469 ) , .ZN( us22_n801 ) );
  NAND2_X1 us22_U366 (.A1( us22_n449 ) , .A2( us22_n452 ) , .ZN( us22_n812 ) );
  NAND2_X1 us22_U367 (.A1( us22_n449 ) , .A2( us22_n469 ) , .ZN( us22_n814 ) );
  NAND2_X1 us22_U368 (.A1( us22_n452 ) , .A2( us22_n459 ) , .ZN( us22_n811 ) );
  NAND2_X1 us22_U369 (.A1( us22_n451 ) , .A2( us22_n459 ) , .ZN( us22_n742 ) );
  NOR4_X1 us22_U37 (.A4( us22_n732 ) , .A3( us22_n733 ) , .A2( us22_n734 ) , .A1( us22_n735 ) , .ZN( us22_n736 ) );
  NAND2_X1 us22_U370 (.A1( us22_n450 ) , .A2( us22_n463 ) , .ZN( us22_n667 ) );
  NAND2_X1 us22_U371 (.A2( us22_n446 ) , .A1( us22_n458 ) , .ZN( us22_n726 ) );
  NAND2_X1 us22_U372 (.A1( us22_n453 ) , .A2( us22_n460 ) , .ZN( us22_n748 ) );
  NAND2_X1 us22_U373 (.A2( us22_n451 ) , .A1( us22_n453 ) , .ZN( us22_n804 ) );
  NAND2_X1 us22_U374 (.A2( us22_n452 ) , .A1( us22_n470 ) , .ZN( us22_n777 ) );
  NAND2_X1 us22_U375 (.A1( us22_n451 ) , .A2( us22_n470 ) , .ZN( us22_n783 ) );
  NAND2_X1 us22_U376 (.A2( us22_n462 ) , .A1( us22_n463 ) , .ZN( us22_n810 ) );
  NAND2_X1 us22_U377 (.A1( us22_n439 ) , .A2( us22_n458 ) , .ZN( us22_n697 ) );
  NAND2_X1 us22_U378 (.A2( us22_n447 ) , .A1( us22_n450 ) , .ZN( us22_n761 ) );
  NAND2_X1 us22_U379 (.A2( us22_n446 ) , .A1( us22_n450 ) , .ZN( us22_n727 ) );
  AOI211_X1 us22_U38 (.B( us22_n723 ) , .A( us22_n724 ) , .ZN( us22_n737 ) , .C1( us22_n841 ) , .C2( us22_n853 ) );
  NAND2_X2 us22_U380 (.A2( us22_n459 ) , .A1( us22_n469 ) , .ZN( us22_n695 ) );
  NOR2_X1 us22_U381 (.ZN( us22_n445 ) , .A2( us22_n847 ) , .A1( us22_n856 ) );
  NAND2_X1 us22_U382 (.A2( us22_n459 ) , .A1( us22_n460 ) , .ZN( us22_n745 ) );
  NAND2_X1 us22_U383 (.A1( us22_n460 ) , .A2( us22_n470 ) , .ZN( us22_n786 ) );
  NOR2_X1 us22_U384 (.ZN( us22_n463 ) , .A2( us22_n845 ) , .A1( us22_n846 ) );
  NOR2_X1 us22_U385 (.ZN( us22_n451 ) , .A1( us22_n824 ) , .A2( us22_n825 ) );
  NOR2_X1 us22_U386 (.ZN( us22_n449 ) , .A1( us22_n826 ) , .A2( us22_n827 ) );
  NAND2_X1 us22_U387 (.A2( us22_n452 ) , .A1( us22_n453 ) , .ZN( us22_n728 ) );
  NAND2_X1 us22_U388 (.A1( us22_n449 ) , .A2( us22_n460 ) , .ZN( us22_n788 ) );
  NAND2_X2 us22_U389 (.A2( us22_n446 ) , .A1( us22_n462 ) , .ZN( us22_n813 ) );
  NOR3_X1 us22_U39 (.A3( us22_n720 ) , .A1( us22_n721 ) , .ZN( us22_n738 ) , .A2( us22_n739 ) );
  NAND2_X2 us22_U390 (.A2( us22_n439 ) , .A1( us22_n450 ) , .ZN( us22_n789 ) );
  NAND2_X2 us22_U391 (.A1( us22_n447 ) , .A2( us22_n462 ) , .ZN( us22_n722 ) );
  NAND2_X2 us22_U392 (.A1( us22_n447 ) , .A2( us22_n458 ) , .ZN( us22_n790 ) );
  NAND2_X2 us22_U393 (.A1( us22_n439 ) , .A2( us22_n462 ) , .ZN( us22_n706 ) );
  NAND2_X2 us22_U394 (.A2( us22_n469 ) , .A1( us22_n470 ) , .ZN( us22_n815 ) );
  NAND2_X2 us22_U395 (.A2( us22_n458 ) , .A1( us22_n463 ) , .ZN( us22_n778 ) );
  NAND2_X1 us22_U396 (.A1( us22_n445 ) , .A2( us22_n447 ) , .ZN( us22_n803 ) );
  NOR2_X1 us22_U397 (.A2( sa22_6 ) , .A1( sa22_7 ) , .ZN( us22_n462 ) );
  NOR2_X1 us22_U398 (.A2( sa22_4 ) , .ZN( us22_n447 ) , .A1( us22_n846 ) );
  NOR2_X1 us22_U399 (.A2( sa22_5 ) , .ZN( us22_n446 ) , .A1( us22_n845 ) );
  INV_X1 us22_U4 (.A( us22_n784 ) , .ZN( us22_n860 ) );
  NAND4_X1 us22_U40 (.ZN( sa20_sr_3 ) , .A4( us22_n702 ) , .A3( us22_n703 ) , .A2( us22_n704 ) , .A1( us22_n705 ) );
  NOR2_X1 us22_U400 (.A2( sa22_7 ) , .ZN( us22_n458 ) , .A1( us22_n847 ) );
  NOR2_X1 us22_U401 (.A2( sa22_4 ) , .A1( sa22_5 ) , .ZN( us22_n439 ) );
  NOR2_X1 us22_U402 (.A2( sa22_1 ) , .ZN( us22_n469 ) , .A1( us22_n824 ) );
  NOR2_X1 us22_U403 (.A2( sa22_2 ) , .A1( sa22_3 ) , .ZN( us22_n470 ) );
  NOR2_X1 us22_U404 (.A2( sa22_6 ) , .ZN( us22_n450 ) , .A1( us22_n856 ) );
  NOR2_X1 us22_U405 (.A2( sa22_2 ) , .ZN( us22_n459 ) , .A1( us22_n827 ) );
  NOR2_X1 us22_U406 (.A2( sa22_0 ) , .ZN( us22_n452 ) , .A1( us22_n825 ) );
  NOR2_X1 us22_U407 (.A2( sa22_0 ) , .A1( sa22_1 ) , .ZN( us22_n460 ) );
  NOR2_X1 us22_U408 (.A2( sa22_3 ) , .ZN( us22_n453 ) , .A1( us22_n826 ) );
  INV_X1 us22_U409 (.A( sa22_6 ) , .ZN( us22_n847 ) );
  NOR4_X1 us22_U41 (.A4( us22_n698 ) , .A3( us22_n699 ) , .A2( us22_n700 ) , .A1( us22_n701 ) , .ZN( us22_n702 ) );
  INV_X1 us22_U410 (.A( sa22_3 ) , .ZN( us22_n827 ) );
  INV_X1 us22_U411 (.A( sa22_1 ) , .ZN( us22_n825 ) );
  INV_X1 us22_U412 (.A( sa22_2 ) , .ZN( us22_n826 ) );
  INV_X1 us22_U413 (.A( sa22_0 ) , .ZN( us22_n824 ) );
  INV_X1 us22_U414 (.A( sa22_7 ) , .ZN( us22_n856 ) );
  INV_X1 us22_U415 (.A( sa22_5 ) , .ZN( us22_n846 ) );
  OAI221_X1 us22_U416 (.A( us22_n781 ) , .C2( us22_n782 ) , .B2( us22_n783 ) , .B1( us22_n784 ) , .ZN( us22_n794 ) , .C1( us22_n811 ) );
  NAND2_X1 us22_U417 (.A1( us22_n727 ) , .A2( us22_n782 ) , .ZN( us22_n809 ) );
  OAI22_X1 us22_U418 (.ZN( us22_n586 ) , .A2( us22_n745 ) , .B2( us22_n760 ) , .A1( us22_n761 ) , .B1( us22_n782 ) );
  OAI221_X1 us22_U419 (.A( us22_n694 ) , .ZN( us22_n701 ) , .C2( us22_n782 ) , .C1( us22_n783 ) , .B1( us22_n784 ) , .B2( us22_n804 ) );
  AOI211_X1 us22_U42 (.B( us22_n692 ) , .A( us22_n693 ) , .ZN( us22_n703 ) , .C2( us22_n829 ) , .C1( us22_n849 ) );
  AOI21_X1 us22_U420 (.ZN( us22_n590 ) , .B1( us22_n726 ) , .B2( us22_n782 ) , .A( us22_n788 ) );
  AOI21_X1 us22_U421 (.ZN( us22_n621 ) , .B1( us22_n697 ) , .A( us22_n777 ) , .B2( us22_n782 ) );
  AOI21_X1 us22_U422 (.ZN( us22_n646 ) , .A( us22_n760 ) , .B2( us22_n782 ) , .B1( us22_n790 ) );
  OAI22_X1 us22_U423 (.ZN( us22_n679 ) , .A1( us22_n697 ) , .A2( us22_n728 ) , .B2( us22_n782 ) , .B1( us22_n815 ) );
  OAI21_X1 us22_U424 (.A( us22_n611 ) , .ZN( us22_n614 ) , .B1( us22_n623 ) , .B2( us22_n782 ) );
  NOR2_X1 us22_U425 (.ZN( us22_n608 ) , .A1( us22_n782 ) , .A2( us22_n814 ) );
  OAI222_X1 us22_U426 (.A2( us22_n667 ) , .ZN( us22_n672 ) , .B1( us22_n745 ) , .B2( us22_n782 ) , .C2( us22_n786 ) , .C1( us22_n813 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U427 (.ZN( us22_n649 ) , .A1( us22_n782 ) , .A2( us22_n786 ) );
  NOR2_X1 us22_U428 (.ZN( us22_n598 ) , .A2( us22_n695 ) , .A1( us22_n782 ) );
  NOR2_X1 us22_U429 (.ZN( us22_n551 ) , .A2( us22_n742 ) , .A1( us22_n782 ) );
  NOR2_X1 us22_U43 (.ZN( us22_n705 ) , .A2( us22_n774 ) , .A1( us22_n798 ) );
  INV_X1 us22_U430 (.A( us22_n782 ) , .ZN( us22_n859 ) );
  NAND4_X1 us22_U431 (.ZN( sa20_sr_2 ) , .A4( us22_n641 ) , .A3( us22_n642 ) , .A1( us22_n643 ) , .A2( us22_n644 ) );
  AOI221_X1 us22_U432 (.A( us22_n574 ) , .ZN( us22_n585 ) , .B2( us22_n829 ) , .C2( us22_n841 ) , .B1( us22_n852 ) , .C1( us22_n859 ) );
  AOI21_X1 us22_U433 (.ZN( us22_n574 ) , .B2( us22_n722 ) , .B1( us22_n746 ) , .A( us22_n783 ) );
  AOI211_X1 us22_U434 (.A( us22_n635 ) , .ZN( us22_n643 ) , .B( us22_n741 ) , .C2( us22_n837 ) , .C1( us22_n852 ) );
  NAND4_X1 us22_U435 (.A4( us22_n631 ) , .A3( us22_n632 ) , .A2( us22_n633 ) , .A1( us22_n634 ) , .ZN( us22_n741 ) );
  INV_X1 us22_U436 (.A( sa22_4 ) , .ZN( us22_n845 ) );
  NAND3_X1 us22_U437 (.ZN( sa20_sr_6 ) , .A3( us22_n795 ) , .A2( us22_n796 ) , .A1( us22_n797 ) );
  NAND3_X1 us22_U438 (.ZN( sa20_sr_5 ) , .A3( us22_n756 ) , .A2( us22_n757 ) , .A1( us22_n758 ) );
  NAND3_X1 us22_U439 (.ZN( sa20_sr_4 ) , .A3( us22_n736 ) , .A2( us22_n737 ) , .A1( us22_n738 ) );
  AOI222_X1 us22_U44 (.B2( us22_n636 ) , .ZN( us22_n642 ) , .B1( us22_n839 ) , .A1( us22_n840 ) , .C2( us22_n844 ) , .C1( us22_n861 ) , .A2( us22_n863 ) );
  NAND3_X1 us22_U440 (.A3( us22_n673 ) , .A2( us22_n674 ) , .A1( us22_n675 ) , .ZN( us22_n805 ) );
  NAND3_X1 us22_U441 (.ZN( us22_n636 ) , .A3( us22_n706 ) , .A2( us22_n722 ) , .A1( us22_n790 ) );
  NAND3_X1 us22_U442 (.A3( us22_n616 ) , .A2( us22_n617 ) , .A1( us22_n618 ) , .ZN( us22_n723 ) );
  NAND3_X1 us22_U443 (.A3( us22_n583 ) , .A2( us22_n584 ) , .A1( us22_n585 ) , .ZN( us22_n619 ) );
  NAND3_X1 us22_U444 (.ZN( us22_n563 ) , .A3( us22_n678 ) , .A2( us22_n748 ) , .A1( us22_n783 ) );
  NAND3_X1 us22_U445 (.A3( us22_n521 ) , .A2( us22_n522 ) , .A1( us22_n523 ) , .ZN( us22_n740 ) );
  NAND3_X1 us22_U446 (.A3( us22_n510 ) , .A1( us22_n511 ) , .ZN( us22_n606 ) , .A2( us22_n869 ) );
  NAND3_X1 us22_U447 (.A3( us22_n465 ) , .A2( us22_n466 ) , .A1( us22_n467 ) , .ZN( us22_n775 ) );
  NOR4_X1 us22_U45 (.A4( us22_n637 ) , .A3( us22_n638 ) , .A2( us22_n639 ) , .A1( us22_n640 ) , .ZN( us22_n641 ) );
  NOR3_X1 us22_U46 (.A2( us22_n605 ) , .A1( us22_n606 ) , .ZN( us22_n644 ) , .A3( us22_n720 ) );
  NOR2_X1 us22_U47 (.ZN( us22_n802 ) , .A1( us22_n852 ) , .A2( us22_n859 ) );
  NAND4_X1 us22_U48 (.ZN( sa20_sr_7 ) , .A4( us22_n820 ) , .A3( us22_n821 ) , .A2( us22_n822 ) , .A1( us22_n823 ) );
  NOR4_X1 us22_U49 (.A4( us22_n816 ) , .A3( us22_n817 ) , .A2( us22_n818 ) , .A1( us22_n819 ) , .ZN( us22_n820 ) );
  NOR3_X1 us22_U5 (.ZN( us22_n596 ) , .A1( us22_n606 ) , .A3( us22_n721 ) , .A2( us22_n740 ) );
  AOI222_X1 us22_U50 (.C2( us22_n807 ) , .B2( us22_n808 ) , .A2( us22_n809 ) , .ZN( us22_n821 ) , .C1( us22_n830 ) , .A1( us22_n837 ) , .B1( us22_n851 ) );
  AOI211_X1 us22_U51 (.B( us22_n805 ) , .A( us22_n806 ) , .ZN( us22_n822 ) , .C1( us22_n840 ) , .C2( us22_n848 ) );
  NAND4_X1 us22_U52 (.ZN( sa20_sr_0 ) , .A4( us22_n499 ) , .A3( us22_n500 ) , .A2( us22_n501 ) , .A1( us22_n502 ) );
  AOI221_X1 us22_U53 (.A( us22_n495 ) , .ZN( us22_n500 ) , .B2( us22_n841 ) , .C1( us22_n844 ) , .C2( us22_n858 ) , .B1( us22_n860 ) );
  NOR4_X1 us22_U54 (.A4( us22_n496 ) , .A3( us22_n497 ) , .A2( us22_n498 ) , .ZN( us22_n499 ) , .A1( us22_n525 ) );
  AOI211_X1 us22_U55 (.A( us22_n494 ) , .ZN( us22_n501 ) , .B( us22_n800 ) , .C2( us22_n837 ) , .C1( us22_n849 ) );
  NOR2_X1 us22_U56 (.ZN( us22_n746 ) , .A1( us22_n859 ) , .A2( us22_n860 ) );
  NAND4_X1 us22_U57 (.ZN( sa20_sr_1 ) , .A4( us22_n593 ) , .A3( us22_n594 ) , .A2( us22_n595 ) , .A1( us22_n596 ) );
  NOR4_X1 us22_U58 (.A4( us22_n589 ) , .A3( us22_n590 ) , .A2( us22_n591 ) , .A1( us22_n592 ) , .ZN( us22_n593 ) );
  AOI211_X1 us22_U59 (.B( us22_n587 ) , .A( us22_n588 ) , .ZN( us22_n594 ) , .C2( us22_n809 ) , .C1( us22_n831 ) );
  NOR3_X1 us22_U6 (.A3( us22_n798 ) , .A2( us22_n799 ) , .A1( us22_n800 ) , .ZN( us22_n823 ) );
  AOI211_X1 us22_U60 (.A( us22_n586 ) , .ZN( us22_n595 ) , .B( us22_n619 ) , .C1( us22_n843 ) , .C2( us22_n853 ) );
  NOR2_X1 us22_U61 (.ZN( us22_n623 ) , .A2( us22_n834 ) , .A1( us22_n837 ) );
  AOI222_X1 us22_U62 (.ZN( us22_n467 ) , .B1( us22_n830 ) , .A1( us22_n837 ) , .C1( us22_n840 ) , .C2( us22_n849 ) , .A2( us22_n853 ) , .B2( us22_n863 ) );
  NOR4_X1 us22_U63 (.A1( us22_n464 ) , .ZN( us22_n465 ) , .A4( us22_n540 ) , .A2( us22_n552 ) , .A3( us22_n612 ) );
  AOI221_X1 us22_U64 (.ZN( us22_n466 ) , .C2( us22_n712 ) , .B2( us22_n829 ) , .C1( us22_n843 ) , .B1( us22_n858 ) , .A( us22_n862 ) );
  NAND4_X1 us22_U65 (.A4( us22_n601 ) , .A3( us22_n602 ) , .A2( us22_n603 ) , .A1( us22_n604 ) , .ZN( us22_n720 ) );
  NOR3_X1 us22_U66 (.A1( us22_n597 ) , .ZN( us22_n602 ) , .A3( us22_n661 ) , .A2( us22_n768 ) );
  NOR4_X1 us22_U67 (.A3( us22_n598 ) , .A2( us22_n599 ) , .A1( us22_n600 ) , .ZN( us22_n601 ) , .A4( us22_n653 ) );
  AOI222_X1 us22_U68 (.ZN( us22_n604 ) , .A1( us22_n828 ) , .C2( us22_n835 ) , .B1( us22_n840 ) , .A2( us22_n854 ) , .B2( us22_n859 ) , .C1( us22_n866 ) );
  NOR4_X1 us22_U69 (.A4( us22_n575 ) , .A3( us22_n576 ) , .A2( us22_n577 ) , .ZN( us22_n584 ) , .A1( us22_n681 ) );
  NOR3_X1 us22_U7 (.ZN( us22_n502 ) , .A2( us22_n677 ) , .A3( us22_n775 ) , .A1( us22_n874 ) );
  NOR4_X1 us22_U70 (.A1( us22_n582 ) , .ZN( us22_n583 ) , .A3( us22_n650 ) , .A2( us22_n660 ) , .A4( us22_n765 ) );
  AOI211_X1 us22_U71 (.B( us22_n621 ) , .A( us22_n622 ) , .ZN( us22_n633 ) , .C2( us22_n834 ) , .C1( us22_n861 ) );
  NOR4_X1 us22_U72 (.A4( us22_n627 ) , .A3( us22_n628 ) , .A2( us22_n629 ) , .A1( us22_n630 ) , .ZN( us22_n631 ) );
  NOR4_X1 us22_U73 (.A4( us22_n624 ) , .A3( us22_n625 ) , .A2( us22_n626 ) , .ZN( us22_n632 ) , .A1( us22_n662 ) );
  NAND4_X1 us22_U74 (.A4( us22_n655 ) , .A3( us22_n656 ) , .A2( us22_n657 ) , .A1( us22_n658 ) , .ZN( us22_n798 ) );
  NOR3_X1 us22_U75 (.A3( us22_n646 ) , .A2( us22_n647 ) , .A1( us22_n648 ) , .ZN( us22_n657 ) );
  NOR3_X1 us22_U76 (.A3( us22_n649 ) , .A2( us22_n650 ) , .A1( us22_n651 ) , .ZN( us22_n656 ) );
  NOR3_X1 us22_U77 (.A3( us22_n652 ) , .A2( us22_n653 ) , .A1( us22_n654 ) , .ZN( us22_n655 ) );
  NAND4_X1 us22_U78 (.A4( us22_n558 ) , .A3( us22_n559 ) , .A2( us22_n560 ) , .A1( us22_n561 ) , .ZN( us22_n605 ) );
  NOR4_X1 us22_U79 (.A4( us22_n554 ) , .A3( us22_n555 ) , .A2( us22_n556 ) , .A1( us22_n557 ) , .ZN( us22_n558 ) );
  INV_X1 us22_U8 (.A( us22_n704 ) , .ZN( us22_n874 ) );
  NOR4_X1 us22_U80 (.ZN( us22_n559 ) , .A1( us22_n651 ) , .A3( us22_n659 ) , .A4( us22_n683 ) , .A2( us22_n766 ) );
  NOR4_X1 us22_U81 (.A4( us22_n550 ) , .A3( us22_n551 ) , .A2( us22_n552 ) , .A1( us22_n553 ) , .ZN( us22_n560 ) );
  NAND4_X1 us22_U82 (.A4( us22_n770 ) , .A3( us22_n771 ) , .A2( us22_n772 ) , .A1( us22_n773 ) , .ZN( us22_n799 ) );
  NOR3_X1 us22_U83 (.A3( us22_n763 ) , .A2( us22_n764 ) , .A1( us22_n765 ) , .ZN( us22_n771 ) );
  NOR4_X1 us22_U84 (.A4( us22_n766 ) , .A3( us22_n767 ) , .A2( us22_n768 ) , .A1( us22_n769 ) , .ZN( us22_n770 ) );
  AOI222_X1 us22_U85 (.ZN( us22_n773 ) , .A1( us22_n828 ) , .C1( us22_n832 ) , .B2( us22_n839 ) , .A2( us22_n848 ) , .B1( us22_n859 ) , .C2( us22_n871 ) );
  NOR4_X1 us22_U86 (.A4( us22_n663 ) , .A3( us22_n664 ) , .A2( us22_n665 ) , .A1( us22_n666 ) , .ZN( us22_n674 ) );
  NOR4_X1 us22_U87 (.A4( us22_n659 ) , .A3( us22_n660 ) , .A2( us22_n661 ) , .A1( us22_n662 ) , .ZN( us22_n675 ) );
  NOR4_X1 us22_U88 (.A3( us22_n671 ) , .A1( us22_n672 ) , .ZN( us22_n673 ) , .A4( us22_n713 ) , .A2( us22_n857 ) );
  NOR2_X1 us22_U89 (.ZN( us22_n759 ) , .A1( us22_n831 ) , .A2( us22_n832 ) );
  NOR3_X1 us22_U9 (.A3( us22_n619 ) , .A2( us22_n620 ) , .ZN( us22_n634 ) , .A1( us22_n723 ) );
  AOI222_X1 us22_U90 (.ZN( us22_n511 ) , .C1( us22_n830 ) , .B2( us22_n835 ) , .A2( us22_n841 ) , .C2( us22_n860 ) , .B1( us22_n861 ) , .A1( us22_n864 ) );
  NOR4_X1 us22_U91 (.A4( us22_n507 ) , .A2( us22_n508 ) , .A1( us22_n509 ) , .ZN( us22_n510 ) , .A3( us22_n668 ) );
  INV_X1 us22_U92 (.A( us22_n503 ) , .ZN( us22_n869 ) );
  NAND4_X1 us22_U93 (.A4( us22_n454 ) , .A3( us22_n455 ) , .A2( us22_n456 ) , .A1( us22_n457 ) , .ZN( us22_n677 ) );
  NOR3_X1 us22_U94 (.ZN( us22_n455 ) , .A3( us22_n528 ) , .A1( us22_n553 ) , .A2( us22_n568 ) );
  AOI221_X1 us22_U95 (.A( us22_n448 ) , .ZN( us22_n457 ) , .C2( us22_n751 ) , .B1( us22_n830 ) , .C1( us22_n840 ) , .B2( us22_n859 ) );
  NOR4_X1 us22_U96 (.ZN( us22_n456 ) , .A2( us22_n507 ) , .A1( us22_n597 ) , .A4( us22_n626 ) , .A3( us22_n709 ) );
  NAND4_X1 us22_U97 (.A4( us22_n533 ) , .A3( us22_n534 ) , .A2( us22_n535 ) , .A1( us22_n536 ) , .ZN( us22_n620 ) );
  NOR4_X1 us22_U98 (.A4( us22_n524 ) , .A2( us22_n525 ) , .A1( us22_n526 ) , .ZN( us22_n536 ) , .A3( us22_n699 ) );
  NOR4_X1 us22_U99 (.A1( us22_n529 ) , .ZN( us22_n534 ) , .A2( us22_n652 ) , .A4( us22_n666 ) , .A3( us22_n763 ) );
endmodule

