module des_des_die_2 ( u0_K10_19, u0_K10_20, u0_K11_21, u0_K11_37, u0_K11_48, u0_K2_11, u0_K2_12, u0_K2_25, u0_K2_30, 
       u0_K2_34, u0_K2_35, u0_K2_4, u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_10, u0_K3_12, u0_K3_14, 
       u0_K3_15, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_5, u0_K4_24, u0_K4_27, u0_K4_28, 
       u0_K4_35, u0_K4_6, u0_K6_19, u0_K6_20, u0_K6_22, u0_K6_23, u0_K6_24, u0_K6_27, u0_K6_41, 
       u0_K7_2, u0_K7_22, u0_K7_23, u0_K8_45, u0_L0_11, u0_L0_12, u0_L0_13, u0_L0_14, u0_L0_17, 
       u0_L0_18, u0_L0_19, u0_L0_2, u0_L0_22, u0_L0_23, u0_L0_25, u0_L0_28, u0_L0_29, u0_L0_3, 
       u0_L0_31, u0_L0_32, u0_L0_4, u0_L0_7, u0_L0_8, u0_L0_9, u0_L11_1, u0_L11_10, u0_L11_13, 
       u0_L11_16, u0_L11_18, u0_L11_2, u0_L11_20, u0_L11_24, u0_L11_26, u0_L11_28, u0_L11_30, u0_L11_6, 
       u0_L13_14, u0_L13_25, u0_L13_3, u0_L13_8, u0_L1_1, u0_L1_10, u0_L1_13, u0_L1_16, u0_L1_17, 
       u0_L1_18, u0_L1_2, u0_L1_20, u0_L1_23, u0_L1_24, u0_L1_26, u0_L1_28, u0_L1_30, u0_L1_31, 
       u0_L1_6, u0_L1_9, u0_L2_1, u0_L2_10, u0_L2_11, u0_L2_13, u0_L2_14, u0_L2_16, u0_L2_17, 
       u0_L2_18, u0_L2_19, u0_L2_2, u0_L2_20, u0_L2_23, u0_L2_24, u0_L2_25, u0_L2_26, u0_L2_28, 
       u0_L2_29, u0_L2_3, u0_L2_30, u0_L2_31, u0_L2_4, u0_L2_6, u0_L2_8, u0_L2_9, u0_L4_1, 
       u0_L4_10, u0_L4_11, u0_L4_12, u0_L4_14, u0_L4_19, u0_L4_20, u0_L4_22, u0_L4_25, u0_L4_26, 
       u0_L4_29, u0_L4_3, u0_L4_32, u0_L4_4, u0_L4_7, u0_L4_8, u0_L5_1, u0_L5_10, u0_L5_13, 
       u0_L5_15, u0_L5_16, u0_L5_17, u0_L5_18, u0_L5_2, u0_L5_20, u0_L5_21, u0_L5_23, u0_L5_24, 
       u0_L5_26, u0_L5_27, u0_L5_28, u0_L5_30, u0_L5_31, u0_L5_5, u0_L5_6, u0_L5_9, u0_L6_15, 
       u0_L6_21, u0_L6_27, u0_L6_5, u0_L8_1, u0_L8_10, u0_L8_20, u0_L8_26, u0_L9_1, u0_L9_10, 
       u0_L9_11, u0_L9_12, u0_L9_13, u0_L9_15, u0_L9_16, u0_L9_18, u0_L9_19, u0_L9_2, u0_L9_20, 
       u0_L9_21, u0_L9_22, u0_L9_24, u0_L9_26, u0_L9_27, u0_L9_28, u0_L9_29, u0_L9_30, u0_L9_32, 
       u0_L9_4, u0_L9_5, u0_L9_6, u0_L9_7, u0_R0_1, u0_R0_16, u0_R0_17, u0_R0_18, u0_R0_19, 
       u0_R0_2, u0_R0_20, u0_R0_21, u0_R0_22, u0_R0_23, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, 
       u0_R0_28, u0_R0_29, u0_R0_3, u0_R0_32, u0_R0_4, u0_R0_5, u0_R0_6, u0_R0_7, u0_R0_8, 
       u0_R0_9, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_17, 
       u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, u0_R11_9, u0_R13_16, u0_R13_17, u0_R13_18, 
       u0_R13_19, u0_R13_20, u0_R13_21, u0_R1_1, u0_R1_10, u0_R1_11, u0_R1_12, u0_R1_13, u0_R1_14, 
       u0_R1_15, u0_R1_16, u0_R1_17, u0_R1_2, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_6, 
       u0_R1_7, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, 
       u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_18, u0_R2_19, u0_R2_2, u0_R2_20, u0_R2_21, u0_R2_22, 
       u0_R2_23, u0_R2_24, u0_R2_25, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, 
       u0_R2_8, u0_R2_9, u0_R4_12, u0_R4_13, u0_R4_14, u0_R4_15, u0_R4_16, u0_R4_17, u0_R4_18, 
       u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_23, u0_R4_24, u0_R4_25, u0_R4_26, u0_R4_27, 
       u0_R4_28, u0_R4_29, u0_R5_1, u0_R5_10, u0_R5_11, u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_15, 
       u0_R5_16, u0_R5_17, u0_R5_2, u0_R5_28, u0_R5_29, u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, 
       u0_R5_4, u0_R5_5, u0_R5_6, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_1, u0_R6_28, u0_R6_29, 
       u0_R6_30, u0_R6_31, u0_R6_32, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, u0_R8_17, 
       u0_R9_1, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_14, u0_R9_15, u0_R9_16, u0_R9_17, 
       u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_28, 
       u0_R9_29, u0_R9_30, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, 
       u0_R9_9, u0_key_r_33, u0_key_r_46, u0_uk_K_r0_15, u0_uk_K_r0_22, u0_uk_K_r0_25, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_34, 
       u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_55, u0_uk_K_r0_7, u0_uk_K_r10_16, u0_uk_K_r11_10, u0_uk_K_r11_11, u0_uk_K_r11_17, u0_uk_K_r11_19, 
       u0_uk_K_r11_20, u0_uk_K_r11_27, u0_uk_K_r11_28, u0_uk_K_r11_33, u0_uk_K_r11_34, u0_uk_K_r11_39, u0_uk_K_r11_47, u0_uk_K_r11_48, u0_uk_K_r11_54, 
       u0_uk_K_r11_6, u0_uk_K_r12_42, u0_uk_K_r13_0, u0_uk_K_r13_22, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_36, 
       u0_uk_K_r1_41, u0_uk_K_r1_47, u0_uk_K_r2_13, u0_uk_K_r2_16, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, 
       u0_uk_K_r2_28, u0_uk_K_r2_31, u0_uk_K_r2_33, u0_uk_K_r2_36, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_53, u0_uk_K_r2_55, 
       u0_uk_K_r2_7, u0_uk_K_r3_4, u0_uk_K_r4_0, u0_uk_K_r4_11, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_48, u0_uk_K_r4_49, u0_uk_K_r4_5, 
       u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_18, u0_uk_K_r5_19, u0_uk_K_r5_26, u0_uk_K_r5_32, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_40, 
       u0_uk_K_r5_41, u0_uk_K_r5_48, u0_uk_K_r5_5, u0_uk_K_r6_0, u0_uk_K_r6_37, u0_uk_K_r8_13, u0_uk_K_r8_21, u0_uk_K_r8_40, u0_uk_K_r8_43, 
       u0_uk_K_r9_10, u0_uk_K_r9_12, u0_uk_K_r9_13, u0_uk_K_r9_15, u0_uk_K_r9_18, u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_23, u0_uk_K_r9_25, 
       u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_31, u0_uk_K_r9_33, u0_uk_K_r9_45, u0_uk_K_r9_48, u0_uk_K_r9_49, u0_uk_K_r9_6, u0_uk_K_r9_7, 
       u0_uk_K_r9_9, u0_uk_n10, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n101, u0_uk_n1019, u0_uk_n1020, u0_uk_n107, 
       u0_uk_n108, u0_uk_n115, u0_uk_n117, u0_uk_n12, u0_uk_n121, u0_uk_n122, u0_uk_n126, u0_uk_n127, u0_uk_n132, 
       u0_uk_n141, u0_uk_n163, u0_uk_n17, u0_uk_n184, u0_uk_n185, u0_uk_n186, u0_uk_n188, u0_uk_n190, u0_uk_n191, 
       u0_uk_n193, u0_uk_n194, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n200, u0_uk_n201, 
       u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n208, u0_uk_n21, u0_uk_n210, u0_uk_n211, u0_uk_n212, u0_uk_n215, 
       u0_uk_n216, u0_uk_n218, u0_uk_n221, u0_uk_n224, u0_uk_n225, u0_uk_n226, u0_uk_n228, u0_uk_n23, u0_uk_n230, 
       u0_uk_n231, u0_uk_n257, u0_uk_n259, u0_uk_n268, u0_uk_n27, u0_uk_n320, u0_uk_n321, u0_uk_n326, u0_uk_n327, 
       u0_uk_n33, u0_uk_n347, u0_uk_n354, u0_uk_n361, u0_uk_n362, u0_uk_n364, u0_uk_n367, u0_uk_n370, u0_uk_n371, 
       u0_uk_n374, u0_uk_n378, u0_uk_n381, u0_uk_n383, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n39, u0_uk_n390, 
       u0_uk_n392, u0_uk_n393, u0_uk_n396, u0_uk_n397, u0_uk_n398, u0_uk_n399, u0_uk_n400, u0_uk_n401, u0_uk_n402, 
       u0_uk_n403, u0_uk_n404, u0_uk_n405, u0_uk_n41, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n417, u0_uk_n418, 
       u0_uk_n419, u0_uk_n420, u0_uk_n424, u0_uk_n425, u0_uk_n428, u0_uk_n430, u0_uk_n433, u0_uk_n434, u0_uk_n438, 
       u0_uk_n439, u0_uk_n440, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n450, u0_uk_n497, u0_uk_n5, u0_uk_n502, 
       u0_uk_n506, u0_uk_n507, u0_uk_n508, u0_uk_n510, u0_uk_n511, u0_uk_n512, u0_uk_n513, u0_uk_n517, u0_uk_n519, 
       u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, u0_uk_n535, 
       u0_uk_n536, u0_uk_n539, u0_uk_n540, u0_uk_n542, u0_uk_n547, u0_uk_n552, u0_uk_n557, u0_uk_n562, u0_uk_n563, 
       u0_uk_n564, u0_uk_n565, u0_uk_n567, u0_uk_n568, u0_uk_n569, u0_uk_n571, u0_uk_n573, u0_uk_n576, u0_uk_n577, 
       u0_uk_n578, u0_uk_n583, u0_uk_n584, u0_uk_n592, u0_uk_n593, u0_uk_n594, u0_uk_n597, u0_uk_n599, u0_uk_n600, 
       u0_uk_n604, u0_uk_n606, u0_uk_n607, u0_uk_n612, u0_uk_n613, u0_uk_n615, u0_uk_n616, u0_uk_n619, u0_uk_n621, 
       u0_uk_n622, u0_uk_n623, u0_uk_n626, u0_uk_n628, u0_uk_n63, u0_uk_n746, u0_uk_n763, u0_uk_n765, u0_uk_n780, 
       u0_uk_n826, u0_uk_n83, u0_uk_n832, u0_uk_n834, u0_uk_n839, u0_uk_n853, u0_uk_n855, u0_uk_n91, u0_uk_n92, 
       u0_uk_n93, u0_uk_n939, u0_uk_n950, u0_uk_n960, u0_uk_n99, u0_uk_n990, u0_uk_n999, u1_L0_1, u1_L0_10, 
       u1_L0_20, u1_L0_26, u1_R0_12, u1_R0_13, u1_R0_14, u1_R0_15, u1_R0_16, u1_R0_17, u1_uk_K_r0_11, 
       u1_uk_K_r0_47, u1_uk_n1263, u1_uk_n1264, u1_uk_n1268, u1_uk_n1273, u1_uk_n1278, u1_uk_n1279, u1_uk_n1290, u1_uk_n1292, 
       u1_uk_n1299, u1_uk_n141, u1_uk_n142, u1_uk_n163, u1_uk_n164, u1_uk_n191, u1_uk_n220, u1_uk_n222, u1_uk_n223, 
       u1_uk_n231, u1_uk_n31, u1_uk_n60, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, u2_FP_38, 
       u2_FP_39, u2_FP_40, u2_FP_41, u2_FP_42, u2_FP_43, u2_FP_44, u2_FP_45, u2_FP_46, u2_FP_47, 
       u2_FP_48, u2_FP_49, u2_FP_64, u2_K10_10, u2_K10_11, u2_K10_15, u2_K10_17, u2_K11_38, u2_K11_42, 
       u2_K12_25, u2_K12_26, u2_K12_27, u2_K12_29, u2_K12_34, u2_K12_37, u2_K12_41, u2_K12_46, u2_K12_47, 
       u2_K15_1, u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_21, u2_K15_23, u2_K15_5, 
       u2_K16_5, u2_K16_6, u2_K16_8, u2_K16_9, u2_K1_15, u2_K1_16, u2_K1_5, u2_K1_9, u2_K2_1, 
       u2_K6_13, u2_K6_14, u2_K6_15, u2_K6_16, u2_K6_20, u2_K6_22, u2_K6_24, u2_K6_32, u2_K6_34, 
       u2_K6_36, u2_K6_40, u2_K7_3, u2_K7_4, u2_K7_5, u2_K7_7, u2_L0_13, u2_L0_17, u2_L0_18, 
       u2_L0_2, u2_L0_23, u2_L0_28, u2_L0_31, u2_L0_9, u2_L10_11, u2_L10_12, u2_L10_14, u2_L10_15, 
       u2_L10_19, u2_L10_21, u2_L10_22, u2_L10_25, u2_L10_27, u2_L10_29, u2_L10_3, u2_L10_32, u2_L10_4, 
       u2_L10_5, u2_L10_7, u2_L10_8, u2_L13_1, u2_L13_10, u2_L13_13, u2_L13_16, u2_L13_17, u2_L13_18, 
       u2_L13_2, u2_L13_20, u2_L13_23, u2_L13_24, u2_L13_26, u2_L13_28, u2_L13_30, u2_L13_31, u2_L13_6, 
       u2_L13_9, u2_L14_1, u2_L14_10, u2_L14_13, u2_L14_16, u2_L14_17, u2_L14_18, u2_L14_2, u2_L14_20, 
       u2_L14_23, u2_L14_24, u2_L14_26, u2_L14_28, u2_L14_30, u2_L14_31, u2_L14_6, u2_L14_9, u2_L4_1, 
       u2_L4_10, u2_L4_11, u2_L4_12, u2_L4_16, u2_L4_19, u2_L4_20, u2_L4_22, u2_L4_24, u2_L4_26, 
       u2_L4_29, u2_L4_30, u2_L4_32, u2_L4_4, u2_L4_6, u2_L4_7, u2_L5_13, u2_L5_16, u2_L5_17, 
       u2_L5_18, u2_L5_2, u2_L5_23, u2_L5_24, u2_L5_28, u2_L5_30, u2_L5_31, u2_L5_6, u2_L5_9, 
       u2_L8_13, u2_L8_16, u2_L8_18, u2_L8_2, u2_L8_24, u2_L8_28, u2_L8_30, u2_L8_6, u2_L9_11, 
       u2_L9_12, u2_L9_19, u2_L9_22, u2_L9_29, u2_L9_32, u2_L9_4, u2_L9_7, u2_R0_1, u2_R0_2, 
       u2_R0_3, u2_R0_32, u2_R0_4, u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, 
       u2_R10_16, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_20, u2_R10_21, u2_R10_22, u2_R10_23, u2_R10_24, 
       u2_R10_25, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_29, u2_R10_30, u2_R10_31, u2_R10_32, u2_R13_1, 
       u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_14, u2_R13_15, u2_R13_16, u2_R13_17, u2_R13_2, 
       u2_R13_3, u2_R13_32, u2_R13_4, u2_R13_5, u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R4_10, 
       u2_R4_11, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_15, u2_R4_16, u2_R4_17, u2_R4_20, u2_R4_21, 
       u2_R4_22, u2_R4_23, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_27, u2_R4_28, u2_R4_29, u2_R4_8, 
       u2_R4_9, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_2, u2_R5_3, u2_R5_32, 
       u2_R5_4, u2_R5_5, u2_R5_6, u2_R5_7, u2_R5_8, u2_R5_9, u2_R8_10, u2_R8_11, u2_R8_12, 
       u2_R8_13, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_7, u2_R8_8, u2_R8_9, u2_R9_20, u2_R9_21, 
       u2_R9_22, u2_R9_23, u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_desIn_r_10, 
       u2_desIn_r_13, u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_2, u2_desIn_r_21, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_29, u2_desIn_r_31, 
       u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_5, 
       u2_desIn_r_50, u2_desIn_r_55, u2_desIn_r_58, u2_desIn_r_60, u2_desIn_r_63, u2_desIn_r_7, u2_key_r_10, u2_key_r_11, u2_key_r_12, 
       u2_key_r_13, u2_key_r_17, u2_key_r_19, u2_key_r_20, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_27, u2_key_r_3, 
       u2_key_r_34, u2_key_r_4, u2_key_r_41, u2_key_r_46, u2_key_r_48, u2_key_r_53, u2_key_r_54, u2_key_r_6, u2_key_r_8, 
       u2_u0_X_1, u2_uk_K_r0_13, u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_34, u2_uk_K_r0_55, u2_uk_K_r10_16, u2_uk_K_r10_43, u2_uk_K_r10_44, 
       u2_uk_K_r10_49, u2_uk_K_r11_7, u2_uk_K_r13_13, u2_uk_K_r13_17, u2_uk_K_r13_19, u2_uk_K_r13_25, u2_uk_K_r13_32, u2_uk_K_r13_55, u2_uk_K_r14_10, 
       u2_uk_K_r14_12, u2_uk_K_r14_18, u2_uk_K_r14_3, u2_uk_K_r14_46, u2_uk_K_r14_5, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_38, u2_uk_K_r4_4, 
       u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_16, u2_uk_K_r5_17, u2_uk_K_r5_26, u2_uk_K_r5_37, u2_uk_K_r5_39, u2_uk_K_r5_4, 
       u2_uk_K_r5_41, u2_uk_K_r5_48, u2_uk_K_r6_46, u2_uk_K_r8_17, u2_uk_K_r8_21, u2_uk_K_r8_27, u2_uk_K_r8_32, u2_uk_K_r8_48, u2_uk_K_r9_0, 
       u2_uk_K_r9_31, u2_uk_K_r9_45, u2_uk_K_r9_49, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n1061, u2_uk_n1063, u2_uk_n1069, 
       u2_uk_n1077, u2_uk_n109, u2_uk_n1096, u2_uk_n117, u2_uk_n118, u2_uk_n1190, u2_uk_n1194, u2_uk_n1197, u2_uk_n1198, 
       u2_uk_n1199, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1212, u2_uk_n1213, u2_uk_n1214, u2_uk_n1218, 
       u2_uk_n1219, u2_uk_n1221, u2_uk_n1222, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, u2_uk_n1232, u2_uk_n1233, u2_uk_n1238, 
       u2_uk_n1239, u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1254, u2_uk_n1261, 
       u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, u2_uk_n128, u2_uk_n141, u2_uk_n1411, u2_uk_n1414, u2_uk_n1418, u2_uk_n142, 
       u2_uk_n1425, u2_uk_n1428, u2_uk_n1430, u2_uk_n1433, u2_uk_n1438, u2_uk_n1439, u2_uk_n1442, u2_uk_n1445, u2_uk_n1446, 
       u2_uk_n145, u2_uk_n1453, u2_uk_n1454, u2_uk_n1457, u2_uk_n1458, u2_uk_n146, u2_uk_n1461, u2_uk_n1462, u2_uk_n1466, 
       u2_uk_n1468, u2_uk_n1475, u2_uk_n148, u2_uk_n1487, u2_uk_n1488, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n155, 
       u2_uk_n1590, u2_uk_n1591, u2_uk_n1600, u2_uk_n1604, u2_uk_n1605, u2_uk_n161, u2_uk_n162, u2_uk_n1624, u2_uk_n1630, 
       u2_uk_n1631, u2_uk_n1634, u2_uk_n164, u2_uk_n1640, u2_uk_n1642, u2_uk_n1653, u2_uk_n1659, u2_uk_n1660, u2_uk_n1664, 
       u2_uk_n1665, u2_uk_n1672, u2_uk_n1673, u2_uk_n1678, u2_uk_n1680, u2_uk_n1684, u2_uk_n1685, u2_uk_n1687, u2_uk_n1690, 
       u2_uk_n1691, u2_uk_n1698, u2_uk_n1699, u2_uk_n17, u2_uk_n1700, u2_uk_n1705, u2_uk_n1707, u2_uk_n1718, u2_uk_n1814, 
       u2_uk_n1815, u2_uk_n1816, u2_uk_n182, u2_uk_n1820, u2_uk_n1821, u2_uk_n1822, u2_uk_n1823, u2_uk_n1828, u2_uk_n1832, 
       u2_uk_n1833, u2_uk_n1834, u2_uk_n1838, u2_uk_n1839, u2_uk_n1842, u2_uk_n1843, u2_uk_n1850, u2_uk_n1851, u2_uk_n1852, 
       u2_uk_n187, u2_uk_n203, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, 
       u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n240, u2_uk_n27, u2_uk_n31, u2_uk_n373, u2_uk_n376, 
       u2_uk_n377, u2_uk_n379, u2_uk_n456, u2_uk_n467, u2_uk_n468, u2_uk_n472, u2_uk_n503, u2_uk_n504, u2_uk_n63, 
       u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n947, u2_uk_n948, u2_uk_n956, u2_uk_n967, u2_uk_n970, 
       u2_uk_n972, u2_uk_n99, u0_N101, u0_N103, u0_N104, u0_N105, u0_N106, u0_N108, u0_N109, u0_N111, u0_N112, 
        u0_N113, u0_N114, u0_N115, u0_N118, u0_N119, u0_N120, u0_N121, u0_N123, u0_N124, 
        u0_N125, u0_N126, u0_N160, u0_N162, u0_N163, u0_N166, u0_N167, u0_N169, u0_N170, 
        u0_N171, u0_N173, u0_N178, u0_N179, u0_N181, u0_N184, u0_N185, u0_N188, u0_N191, 
        u0_N192, u0_N193, u0_N196, u0_N197, u0_N200, u0_N201, u0_N204, u0_N206, u0_N207, 
        u0_N208, u0_N209, u0_N211, u0_N212, u0_N214, u0_N215, u0_N217, u0_N218, u0_N219, 
        u0_N221, u0_N222, u0_N228, u0_N238, u0_N244, u0_N250, u0_N288, u0_N297, u0_N307, 
        u0_N313, u0_N320, u0_N321, u0_N323, u0_N324, u0_N325, u0_N326, u0_N329, u0_N33, 
        u0_N330, u0_N331, u0_N332, u0_N334, u0_N335, u0_N337, u0_N338, u0_N339, u0_N34, 
        u0_N340, u0_N341, u0_N343, u0_N345, u0_N346, u0_N347, u0_N348, u0_N349, u0_N35, 
        u0_N351, u0_N38, u0_N384, u0_N385, u0_N389, u0_N39, u0_N393, u0_N396, u0_N399, 
        u0_N40, u0_N401, u0_N403, u0_N407, u0_N409, u0_N411, u0_N413, u0_N42, u0_N43, 
        u0_N44, u0_N45, u0_N450, u0_N455, u0_N461, u0_N472, u0_N48, u0_N49, u0_N50, 
        u0_N53, u0_N54, u0_N56, u0_N59, u0_N60, u0_N62, u0_N63, u0_N64, u0_N65, 
        u0_N69, u0_N72, u0_N73, u0_N76, u0_N79, u0_N80, u0_N81, u0_N83, u0_N86, 
        u0_N87, u0_N89, u0_N91, u0_N93, u0_N94, u0_N96, u0_N97, u0_N98, u0_N99, 
        u0_uk_n100, u0_uk_n1010, u0_uk_n1016, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n118, u0_uk_n128, 
        u0_uk_n129, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n161, u0_uk_n162, u0_uk_n164, 
        u0_uk_n182, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, 
        u0_uk_n222, u0_uk_n223, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n31, 
        u0_uk_n60, u0_uk_n691, u0_uk_n773, u0_uk_n778, u0_uk_n798, u0_uk_n804, u0_uk_n848, u0_uk_n863, u0_uk_n867, 
        u0_uk_n890, u0_uk_n936, u0_uk_n94, u0_uk_n945, u0_uk_n969, u1_N32, u1_N41, u1_N51, u1_N57, 
        u2_FP_1, u2_FP_10, u2_FP_13, u2_FP_16, u2_FP_17, u2_FP_18, u2_FP_2, u2_FP_20, u2_FP_23, 
        u2_FP_24, u2_FP_26, u2_FP_28, u2_FP_30, u2_FP_31, u2_FP_6, u2_FP_9, u2_K1_21, u2_N1, 
        u2_N12, u2_N15, u2_N16, u2_N160, u2_N163, u2_N165, u2_N166, u2_N169, u2_N17, 
        u2_N170, u2_N171, u2_N175, u2_N178, u2_N179, u2_N181, u2_N183, u2_N185, u2_N188, 
        u2_N189, u2_N191, u2_N193, u2_N197, u2_N200, u2_N204, u2_N207, u2_N208, u2_N209, 
        u2_N214, u2_N215, u2_N219, u2_N22, u2_N221, u2_N222, u2_N23, u2_N27, u2_N289, 
        u2_N29, u2_N293, u2_N30, u2_N300, u2_N303, u2_N305, u2_N311, u2_N315, u2_N317, 
        u2_N323, u2_N326, u2_N33, u2_N330, u2_N331, u2_N338, u2_N341, u2_N348, u2_N351, 
        u2_N354, u2_N355, u2_N356, u2_N358, u2_N359, u2_N362, u2_N363, u2_N365, u2_N366, 
        u2_N370, u2_N372, u2_N373, u2_N376, u2_N378, u2_N380, u2_N383, u2_N40, u2_N44, 
        u2_N448, u2_N449, u2_N453, u2_N456, u2_N457, u2_N460, u2_N463, u2_N464, u2_N465, 
        u2_N467, u2_N470, u2_N471, u2_N473, u2_N475, u2_N477, u2_N478, u2_N48, u2_N49, 
        u2_N5, u2_N54, u2_N59, u2_N62, u2_N8, u2_uk_n1087, u2_uk_n1090, u2_uk_n11, u2_uk_n110, 
        u2_uk_n1102, u2_uk_n1145, u2_uk_n1146, u2_uk_n1148, u2_uk_n1150, u2_uk_n1155, u2_uk_n1161, u2_uk_n1162, u2_uk_n1168, 
        u2_uk_n1185, u2_uk_n129, u2_uk_n147, u2_uk_n163, u2_uk_n188, u2_uk_n191, u2_uk_n207, u2_uk_n298, u2_uk_n366, 
        u2_uk_n60, u2_uk_n656 );
  input u0_K10_19, u0_K10_20, u0_K11_21, u0_K11_37, u0_K11_48, u0_K2_11, u0_K2_12, u0_K2_25, u0_K2_30, 
        u0_K2_34, u0_K2_35, u0_K2_4, u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_10, u0_K3_12, u0_K3_14, 
        u0_K3_15, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_5, u0_K4_24, u0_K4_27, u0_K4_28, 
        u0_K4_35, u0_K4_6, u0_K6_19, u0_K6_20, u0_K6_22, u0_K6_23, u0_K6_24, u0_K6_27, u0_K6_41, 
        u0_K7_2, u0_K7_22, u0_K7_23, u0_K8_45, u0_L0_11, u0_L0_12, u0_L0_13, u0_L0_14, u0_L0_17, 
        u0_L0_18, u0_L0_19, u0_L0_2, u0_L0_22, u0_L0_23, u0_L0_25, u0_L0_28, u0_L0_29, u0_L0_3, 
        u0_L0_31, u0_L0_32, u0_L0_4, u0_L0_7, u0_L0_8, u0_L0_9, u0_L11_1, u0_L11_10, u0_L11_13, 
        u0_L11_16, u0_L11_18, u0_L11_2, u0_L11_20, u0_L11_24, u0_L11_26, u0_L11_28, u0_L11_30, u0_L11_6, 
        u0_L13_14, u0_L13_25, u0_L13_3, u0_L13_8, u0_L1_1, u0_L1_10, u0_L1_13, u0_L1_16, u0_L1_17, 
        u0_L1_18, u0_L1_2, u0_L1_20, u0_L1_23, u0_L1_24, u0_L1_26, u0_L1_28, u0_L1_30, u0_L1_31, 
        u0_L1_6, u0_L1_9, u0_L2_1, u0_L2_10, u0_L2_11, u0_L2_13, u0_L2_14, u0_L2_16, u0_L2_17, 
        u0_L2_18, u0_L2_19, u0_L2_2, u0_L2_20, u0_L2_23, u0_L2_24, u0_L2_25, u0_L2_26, u0_L2_28, 
        u0_L2_29, u0_L2_3, u0_L2_30, u0_L2_31, u0_L2_4, u0_L2_6, u0_L2_8, u0_L2_9, u0_L4_1, 
        u0_L4_10, u0_L4_11, u0_L4_12, u0_L4_14, u0_L4_19, u0_L4_20, u0_L4_22, u0_L4_25, u0_L4_26, 
        u0_L4_29, u0_L4_3, u0_L4_32, u0_L4_4, u0_L4_7, u0_L4_8, u0_L5_1, u0_L5_10, u0_L5_13, 
        u0_L5_15, u0_L5_16, u0_L5_17, u0_L5_18, u0_L5_2, u0_L5_20, u0_L5_21, u0_L5_23, u0_L5_24, 
        u0_L5_26, u0_L5_27, u0_L5_28, u0_L5_30, u0_L5_31, u0_L5_5, u0_L5_6, u0_L5_9, u0_L6_15, 
        u0_L6_21, u0_L6_27, u0_L6_5, u0_L8_1, u0_L8_10, u0_L8_20, u0_L8_26, u0_L9_1, u0_L9_10, 
        u0_L9_11, u0_L9_12, u0_L9_13, u0_L9_15, u0_L9_16, u0_L9_18, u0_L9_19, u0_L9_2, u0_L9_20, 
        u0_L9_21, u0_L9_22, u0_L9_24, u0_L9_26, u0_L9_27, u0_L9_28, u0_L9_29, u0_L9_30, u0_L9_32, 
        u0_L9_4, u0_L9_5, u0_L9_6, u0_L9_7, u0_R0_1, u0_R0_16, u0_R0_17, u0_R0_18, u0_R0_19, 
        u0_R0_2, u0_R0_20, u0_R0_21, u0_R0_22, u0_R0_23, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, 
        u0_R0_28, u0_R0_29, u0_R0_3, u0_R0_32, u0_R0_4, u0_R0_5, u0_R0_6, u0_R0_7, u0_R0_8, 
        u0_R0_9, u0_R11_10, u0_R11_11, u0_R11_12, u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_17, 
        u0_R11_4, u0_R11_5, u0_R11_6, u0_R11_7, u0_R11_8, u0_R11_9, u0_R13_16, u0_R13_17, u0_R13_18, 
        u0_R13_19, u0_R13_20, u0_R13_21, u0_R1_1, u0_R1_10, u0_R1_11, u0_R1_12, u0_R1_13, u0_R1_14, 
        u0_R1_15, u0_R1_16, u0_R1_17, u0_R1_2, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_6, 
        u0_R1_7, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, 
        u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_18, u0_R2_19, u0_R2_2, u0_R2_20, u0_R2_21, u0_R2_22, 
        u0_R2_23, u0_R2_24, u0_R2_25, u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, 
        u0_R2_8, u0_R2_9, u0_R4_12, u0_R4_13, u0_R4_14, u0_R4_15, u0_R4_16, u0_R4_17, u0_R4_18, 
        u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_23, u0_R4_24, u0_R4_25, u0_R4_26, u0_R4_27, 
        u0_R4_28, u0_R4_29, u0_R5_1, u0_R5_10, u0_R5_11, u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_15, 
        u0_R5_16, u0_R5_17, u0_R5_2, u0_R5_28, u0_R5_29, u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, 
        u0_R5_4, u0_R5_5, u0_R5_6, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_1, u0_R6_28, u0_R6_29, 
        u0_R6_30, u0_R6_31, u0_R6_32, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, u0_R8_17, 
        u0_R9_1, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_14, u0_R9_15, u0_R9_16, u0_R9_17, 
        u0_R9_20, u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_28, 
        u0_R9_29, u0_R9_30, u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, 
        u0_R9_9, u0_key_r_33, u0_key_r_46, u0_uk_K_r0_15, u0_uk_K_r0_22, u0_uk_K_r0_25, u0_uk_K_r0_28, u0_uk_K_r0_31, u0_uk_K_r0_34, 
        u0_uk_K_r0_36, u0_uk_K_r0_49, u0_uk_K_r0_55, u0_uk_K_r0_7, u0_uk_K_r10_16, u0_uk_K_r11_10, u0_uk_K_r11_11, u0_uk_K_r11_17, u0_uk_K_r11_19, 
        u0_uk_K_r11_20, u0_uk_K_r11_27, u0_uk_K_r11_28, u0_uk_K_r11_33, u0_uk_K_r11_34, u0_uk_K_r11_39, u0_uk_K_r11_47, u0_uk_K_r11_48, u0_uk_K_r11_54, 
        u0_uk_K_r11_6, u0_uk_K_r12_42, u0_uk_K_r13_0, u0_uk_K_r13_22, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_36, 
        u0_uk_K_r1_41, u0_uk_K_r1_47, u0_uk_K_r2_13, u0_uk_K_r2_16, u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, 
        u0_uk_K_r2_28, u0_uk_K_r2_31, u0_uk_K_r2_33, u0_uk_K_r2_36, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_53, u0_uk_K_r2_55, 
        u0_uk_K_r2_7, u0_uk_K_r3_4, u0_uk_K_r4_0, u0_uk_K_r4_11, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r4_48, u0_uk_K_r4_49, u0_uk_K_r4_5, 
        u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_18, u0_uk_K_r5_19, u0_uk_K_r5_26, u0_uk_K_r5_32, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r5_40, 
        u0_uk_K_r5_41, u0_uk_K_r5_48, u0_uk_K_r5_5, u0_uk_K_r6_0, u0_uk_K_r6_37, u0_uk_K_r8_13, u0_uk_K_r8_21, u0_uk_K_r8_40, u0_uk_K_r8_43, 
        u0_uk_K_r9_10, u0_uk_K_r9_12, u0_uk_K_r9_13, u0_uk_K_r9_15, u0_uk_K_r9_18, u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_23, u0_uk_K_r9_25, 
        u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_31, u0_uk_K_r9_33, u0_uk_K_r9_45, u0_uk_K_r9_48, u0_uk_K_r9_49, u0_uk_K_r9_6, u0_uk_K_r9_7, 
        u0_uk_K_r9_9, u0_uk_n10, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n101, u0_uk_n1019, u0_uk_n1020, u0_uk_n107, 
        u0_uk_n108, u0_uk_n115, u0_uk_n117, u0_uk_n12, u0_uk_n121, u0_uk_n122, u0_uk_n126, u0_uk_n127, u0_uk_n132, 
        u0_uk_n141, u0_uk_n163, u0_uk_n17, u0_uk_n184, u0_uk_n185, u0_uk_n186, u0_uk_n188, u0_uk_n190, u0_uk_n191, 
        u0_uk_n193, u0_uk_n194, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n200, u0_uk_n201, 
        u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n208, u0_uk_n21, u0_uk_n210, u0_uk_n211, u0_uk_n212, u0_uk_n215, 
        u0_uk_n216, u0_uk_n218, u0_uk_n221, u0_uk_n224, u0_uk_n225, u0_uk_n226, u0_uk_n228, u0_uk_n23, u0_uk_n230, 
        u0_uk_n231, u0_uk_n257, u0_uk_n259, u0_uk_n268, u0_uk_n27, u0_uk_n320, u0_uk_n321, u0_uk_n326, u0_uk_n327, 
        u0_uk_n33, u0_uk_n347, u0_uk_n354, u0_uk_n361, u0_uk_n362, u0_uk_n364, u0_uk_n367, u0_uk_n370, u0_uk_n371, 
        u0_uk_n374, u0_uk_n378, u0_uk_n381, u0_uk_n383, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n39, u0_uk_n390, 
        u0_uk_n392, u0_uk_n393, u0_uk_n396, u0_uk_n397, u0_uk_n398, u0_uk_n399, u0_uk_n400, u0_uk_n401, u0_uk_n402, 
        u0_uk_n403, u0_uk_n404, u0_uk_n405, u0_uk_n41, u0_uk_n411, u0_uk_n412, u0_uk_n413, u0_uk_n417, u0_uk_n418, 
        u0_uk_n419, u0_uk_n420, u0_uk_n424, u0_uk_n425, u0_uk_n428, u0_uk_n430, u0_uk_n433, u0_uk_n434, u0_uk_n438, 
        u0_uk_n439, u0_uk_n440, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n450, u0_uk_n497, u0_uk_n5, u0_uk_n502, 
        u0_uk_n506, u0_uk_n507, u0_uk_n508, u0_uk_n510, u0_uk_n511, u0_uk_n512, u0_uk_n513, u0_uk_n517, u0_uk_n519, 
        u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n532, u0_uk_n534, u0_uk_n535, 
        u0_uk_n536, u0_uk_n539, u0_uk_n540, u0_uk_n542, u0_uk_n547, u0_uk_n552, u0_uk_n557, u0_uk_n562, u0_uk_n563, 
        u0_uk_n564, u0_uk_n565, u0_uk_n567, u0_uk_n568, u0_uk_n569, u0_uk_n571, u0_uk_n573, u0_uk_n576, u0_uk_n577, 
        u0_uk_n578, u0_uk_n583, u0_uk_n584, u0_uk_n592, u0_uk_n593, u0_uk_n594, u0_uk_n597, u0_uk_n599, u0_uk_n600, 
        u0_uk_n604, u0_uk_n606, u0_uk_n607, u0_uk_n612, u0_uk_n613, u0_uk_n615, u0_uk_n616, u0_uk_n619, u0_uk_n621, 
        u0_uk_n622, u0_uk_n623, u0_uk_n626, u0_uk_n628, u0_uk_n63, u0_uk_n746, u0_uk_n763, u0_uk_n765, u0_uk_n780, 
        u0_uk_n826, u0_uk_n83, u0_uk_n832, u0_uk_n834, u0_uk_n839, u0_uk_n853, u0_uk_n855, u0_uk_n91, u0_uk_n92, 
        u0_uk_n93, u0_uk_n939, u0_uk_n950, u0_uk_n960, u0_uk_n99, u0_uk_n990, u0_uk_n999, u1_L0_1, u1_L0_10, 
        u1_L0_20, u1_L0_26, u1_R0_12, u1_R0_13, u1_R0_14, u1_R0_15, u1_R0_16, u1_R0_17, u1_uk_K_r0_11, 
        u1_uk_K_r0_47, u1_uk_n1263, u1_uk_n1264, u1_uk_n1268, u1_uk_n1273, u1_uk_n1278, u1_uk_n1279, u1_uk_n1290, u1_uk_n1292, 
        u1_uk_n1299, u1_uk_n141, u1_uk_n142, u1_uk_n163, u1_uk_n164, u1_uk_n191, u1_uk_n220, u1_uk_n222, u1_uk_n223, 
        u1_uk_n231, u1_uk_n31, u1_uk_n60, u2_FP_33, u2_FP_34, u2_FP_35, u2_FP_36, u2_FP_37, u2_FP_38, 
        u2_FP_39, u2_FP_40, u2_FP_41, u2_FP_42, u2_FP_43, u2_FP_44, u2_FP_45, u2_FP_46, u2_FP_47, 
        u2_FP_48, u2_FP_49, u2_FP_64, u2_K10_10, u2_K10_11, u2_K10_15, u2_K10_17, u2_K11_38, u2_K11_42, 
        u2_K12_25, u2_K12_26, u2_K12_27, u2_K12_29, u2_K12_34, u2_K12_37, u2_K12_41, u2_K12_46, u2_K12_47, 
        u2_K15_1, u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_2, u2_K15_20, u2_K15_21, u2_K15_23, u2_K15_5, 
        u2_K16_5, u2_K16_6, u2_K16_8, u2_K16_9, u2_K1_15, u2_K1_16, u2_K1_5, u2_K1_9, u2_K2_1, 
        u2_K6_13, u2_K6_14, u2_K6_15, u2_K6_16, u2_K6_20, u2_K6_22, u2_K6_24, u2_K6_32, u2_K6_34, 
        u2_K6_36, u2_K6_40, u2_K7_3, u2_K7_4, u2_K7_5, u2_K7_7, u2_L0_13, u2_L0_17, u2_L0_18, 
        u2_L0_2, u2_L0_23, u2_L0_28, u2_L0_31, u2_L0_9, u2_L10_11, u2_L10_12, u2_L10_14, u2_L10_15, 
        u2_L10_19, u2_L10_21, u2_L10_22, u2_L10_25, u2_L10_27, u2_L10_29, u2_L10_3, u2_L10_32, u2_L10_4, 
        u2_L10_5, u2_L10_7, u2_L10_8, u2_L13_1, u2_L13_10, u2_L13_13, u2_L13_16, u2_L13_17, u2_L13_18, 
        u2_L13_2, u2_L13_20, u2_L13_23, u2_L13_24, u2_L13_26, u2_L13_28, u2_L13_30, u2_L13_31, u2_L13_6, 
        u2_L13_9, u2_L14_1, u2_L14_10, u2_L14_13, u2_L14_16, u2_L14_17, u2_L14_18, u2_L14_2, u2_L14_20, 
        u2_L14_23, u2_L14_24, u2_L14_26, u2_L14_28, u2_L14_30, u2_L14_31, u2_L14_6, u2_L14_9, u2_L4_1, 
        u2_L4_10, u2_L4_11, u2_L4_12, u2_L4_16, u2_L4_19, u2_L4_20, u2_L4_22, u2_L4_24, u2_L4_26, 
        u2_L4_29, u2_L4_30, u2_L4_32, u2_L4_4, u2_L4_6, u2_L4_7, u2_L5_13, u2_L5_16, u2_L5_17, 
        u2_L5_18, u2_L5_2, u2_L5_23, u2_L5_24, u2_L5_28, u2_L5_30, u2_L5_31, u2_L5_6, u2_L5_9, 
        u2_L8_13, u2_L8_16, u2_L8_18, u2_L8_2, u2_L8_24, u2_L8_28, u2_L8_30, u2_L8_6, u2_L9_11, 
        u2_L9_12, u2_L9_19, u2_L9_22, u2_L9_29, u2_L9_32, u2_L9_4, u2_L9_7, u2_R0_1, u2_R0_2, 
        u2_R0_3, u2_R0_32, u2_R0_4, u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, 
        u2_R10_16, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_20, u2_R10_21, u2_R10_22, u2_R10_23, u2_R10_24, 
        u2_R10_25, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_29, u2_R10_30, u2_R10_31, u2_R10_32, u2_R13_1, 
        u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_14, u2_R13_15, u2_R13_16, u2_R13_17, u2_R13_2, 
        u2_R13_3, u2_R13_32, u2_R13_4, u2_R13_5, u2_R13_6, u2_R13_7, u2_R13_8, u2_R13_9, u2_R4_10, 
        u2_R4_11, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_15, u2_R4_16, u2_R4_17, u2_R4_20, u2_R4_21, 
        u2_R4_22, u2_R4_23, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_27, u2_R4_28, u2_R4_29, u2_R4_8, 
        u2_R4_9, u2_R5_1, u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_2, u2_R5_3, u2_R5_32, 
        u2_R5_4, u2_R5_5, u2_R5_6, u2_R5_7, u2_R5_8, u2_R5_9, u2_R8_10, u2_R8_11, u2_R8_12, 
        u2_R8_13, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_7, u2_R8_8, u2_R8_9, u2_R9_20, u2_R9_21, 
        u2_R9_22, u2_R9_23, u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_desIn_r_10, 
        u2_desIn_r_13, u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_2, u2_desIn_r_21, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_29, u2_desIn_r_31, 
        u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_5, 
        u2_desIn_r_50, u2_desIn_r_55, u2_desIn_r_58, u2_desIn_r_60, u2_desIn_r_63, u2_desIn_r_7, u2_key_r_10, u2_key_r_11, u2_key_r_12, 
        u2_key_r_13, u2_key_r_17, u2_key_r_19, u2_key_r_20, u2_key_r_24, u2_key_r_25, u2_key_r_26, u2_key_r_27, u2_key_r_3, 
        u2_key_r_34, u2_key_r_4, u2_key_r_41, u2_key_r_46, u2_key_r_48, u2_key_r_53, u2_key_r_54, u2_key_r_6, u2_key_r_8, 
        u2_u0_X_1, u2_uk_K_r0_13, u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_34, u2_uk_K_r0_55, u2_uk_K_r10_16, u2_uk_K_r10_43, u2_uk_K_r10_44, 
        u2_uk_K_r10_49, u2_uk_K_r11_7, u2_uk_K_r13_13, u2_uk_K_r13_17, u2_uk_K_r13_19, u2_uk_K_r13_25, u2_uk_K_r13_32, u2_uk_K_r13_55, u2_uk_K_r14_10, 
        u2_uk_K_r14_12, u2_uk_K_r14_18, u2_uk_K_r14_3, u2_uk_K_r14_46, u2_uk_K_r14_5, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_38, u2_uk_K_r4_4, 
        u2_uk_K_r4_5, u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_16, u2_uk_K_r5_17, u2_uk_K_r5_26, u2_uk_K_r5_37, u2_uk_K_r5_39, u2_uk_K_r5_4, 
        u2_uk_K_r5_41, u2_uk_K_r5_48, u2_uk_K_r6_46, u2_uk_K_r8_17, u2_uk_K_r8_21, u2_uk_K_r8_27, u2_uk_K_r8_32, u2_uk_K_r8_48, u2_uk_K_r9_0, 
        u2_uk_K_r9_31, u2_uk_K_r9_45, u2_uk_K_r9_49, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n1061, u2_uk_n1063, u2_uk_n1069, 
        u2_uk_n1077, u2_uk_n109, u2_uk_n1096, u2_uk_n117, u2_uk_n118, u2_uk_n1190, u2_uk_n1194, u2_uk_n1197, u2_uk_n1198, 
        u2_uk_n1199, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1212, u2_uk_n1213, u2_uk_n1214, u2_uk_n1218, 
        u2_uk_n1219, u2_uk_n1221, u2_uk_n1222, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, u2_uk_n1232, u2_uk_n1233, u2_uk_n1238, 
        u2_uk_n1239, u2_uk_n1240, u2_uk_n1243, u2_uk_n1244, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1254, u2_uk_n1261, 
        u2_uk_n1267, u2_uk_n1270, u2_uk_n1275, u2_uk_n128, u2_uk_n141, u2_uk_n1411, u2_uk_n1414, u2_uk_n1418, u2_uk_n142, 
        u2_uk_n1425, u2_uk_n1428, u2_uk_n1430, u2_uk_n1433, u2_uk_n1438, u2_uk_n1439, u2_uk_n1442, u2_uk_n1445, u2_uk_n1446, 
        u2_uk_n145, u2_uk_n1453, u2_uk_n1454, u2_uk_n1457, u2_uk_n1458, u2_uk_n146, u2_uk_n1461, u2_uk_n1462, u2_uk_n1466, 
        u2_uk_n1468, u2_uk_n1475, u2_uk_n148, u2_uk_n1487, u2_uk_n1488, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n155, 
        u2_uk_n1590, u2_uk_n1591, u2_uk_n1600, u2_uk_n1604, u2_uk_n1605, u2_uk_n161, u2_uk_n162, u2_uk_n1624, u2_uk_n1630, 
        u2_uk_n1631, u2_uk_n1634, u2_uk_n164, u2_uk_n1640, u2_uk_n1642, u2_uk_n1653, u2_uk_n1659, u2_uk_n1660, u2_uk_n1664, 
        u2_uk_n1665, u2_uk_n1672, u2_uk_n1673, u2_uk_n1678, u2_uk_n1680, u2_uk_n1684, u2_uk_n1685, u2_uk_n1687, u2_uk_n1690, 
        u2_uk_n1691, u2_uk_n1698, u2_uk_n1699, u2_uk_n17, u2_uk_n1700, u2_uk_n1705, u2_uk_n1707, u2_uk_n1718, u2_uk_n1814, 
        u2_uk_n1815, u2_uk_n1816, u2_uk_n182, u2_uk_n1820, u2_uk_n1821, u2_uk_n1822, u2_uk_n1823, u2_uk_n1828, u2_uk_n1832, 
        u2_uk_n1833, u2_uk_n1834, u2_uk_n1838, u2_uk_n1839, u2_uk_n1842, u2_uk_n1843, u2_uk_n1850, u2_uk_n1851, u2_uk_n1852, 
        u2_uk_n187, u2_uk_n203, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n222, 
        u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n238, u2_uk_n240, u2_uk_n27, u2_uk_n31, u2_uk_n373, u2_uk_n376, 
        u2_uk_n377, u2_uk_n379, u2_uk_n456, u2_uk_n467, u2_uk_n468, u2_uk_n472, u2_uk_n503, u2_uk_n504, u2_uk_n63, 
        u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n947, u2_uk_n948, u2_uk_n956, u2_uk_n967, u2_uk_n970, 
        u2_uk_n972, u2_uk_n99;
  output u0_N101, u0_N103, u0_N104, u0_N105, u0_N106, u0_N108, u0_N109, u0_N111, u0_N112, 
        u0_N113, u0_N114, u0_N115, u0_N118, u0_N119, u0_N120, u0_N121, u0_N123, u0_N124, 
        u0_N125, u0_N126, u0_N160, u0_N162, u0_N163, u0_N166, u0_N167, u0_N169, u0_N170, 
        u0_N171, u0_N173, u0_N178, u0_N179, u0_N181, u0_N184, u0_N185, u0_N188, u0_N191, 
        u0_N192, u0_N193, u0_N196, u0_N197, u0_N200, u0_N201, u0_N204, u0_N206, u0_N207, 
        u0_N208, u0_N209, u0_N211, u0_N212, u0_N214, u0_N215, u0_N217, u0_N218, u0_N219, 
        u0_N221, u0_N222, u0_N228, u0_N238, u0_N244, u0_N250, u0_N288, u0_N297, u0_N307, 
        u0_N313, u0_N320, u0_N321, u0_N323, u0_N324, u0_N325, u0_N326, u0_N329, u0_N33, 
        u0_N330, u0_N331, u0_N332, u0_N334, u0_N335, u0_N337, u0_N338, u0_N339, u0_N34, 
        u0_N340, u0_N341, u0_N343, u0_N345, u0_N346, u0_N347, u0_N348, u0_N349, u0_N35, 
        u0_N351, u0_N38, u0_N384, u0_N385, u0_N389, u0_N39, u0_N393, u0_N396, u0_N399, 
        u0_N40, u0_N401, u0_N403, u0_N407, u0_N409, u0_N411, u0_N413, u0_N42, u0_N43, 
        u0_N44, u0_N45, u0_N450, u0_N455, u0_N461, u0_N472, u0_N48, u0_N49, u0_N50, 
        u0_N53, u0_N54, u0_N56, u0_N59, u0_N60, u0_N62, u0_N63, u0_N64, u0_N65, 
        u0_N69, u0_N72, u0_N73, u0_N76, u0_N79, u0_N80, u0_N81, u0_N83, u0_N86, 
        u0_N87, u0_N89, u0_N91, u0_N93, u0_N94, u0_N96, u0_N97, u0_N98, u0_N99, 
        u0_uk_n100, u0_uk_n1010, u0_uk_n1016, u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n118, u0_uk_n128, 
        u0_uk_n129, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n161, u0_uk_n162, u0_uk_n164, 
        u0_uk_n182, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, 
        u0_uk_n222, u0_uk_n223, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n31, 
        u0_uk_n60, u0_uk_n691, u0_uk_n773, u0_uk_n778, u0_uk_n798, u0_uk_n804, u0_uk_n848, u0_uk_n863, u0_uk_n867, 
        u0_uk_n890, u0_uk_n936, u0_uk_n94, u0_uk_n945, u0_uk_n969, u1_N32, u1_N41, u1_N51, u1_N57, 
        u2_FP_1, u2_FP_10, u2_FP_13, u2_FP_16, u2_FP_17, u2_FP_18, u2_FP_2, u2_FP_20, u2_FP_23, 
        u2_FP_24, u2_FP_26, u2_FP_28, u2_FP_30, u2_FP_31, u2_FP_6, u2_FP_9, u2_K1_21, u2_N1, 
        u2_N12, u2_N15, u2_N16, u2_N160, u2_N163, u2_N165, u2_N166, u2_N169, u2_N17, 
        u2_N170, u2_N171, u2_N175, u2_N178, u2_N179, u2_N181, u2_N183, u2_N185, u2_N188, 
        u2_N189, u2_N191, u2_N193, u2_N197, u2_N200, u2_N204, u2_N207, u2_N208, u2_N209, 
        u2_N214, u2_N215, u2_N219, u2_N22, u2_N221, u2_N222, u2_N23, u2_N27, u2_N289, 
        u2_N29, u2_N293, u2_N30, u2_N300, u2_N303, u2_N305, u2_N311, u2_N315, u2_N317, 
        u2_N323, u2_N326, u2_N33, u2_N330, u2_N331, u2_N338, u2_N341, u2_N348, u2_N351, 
        u2_N354, u2_N355, u2_N356, u2_N358, u2_N359, u2_N362, u2_N363, u2_N365, u2_N366, 
        u2_N370, u2_N372, u2_N373, u2_N376, u2_N378, u2_N380, u2_N383, u2_N40, u2_N44, 
        u2_N448, u2_N449, u2_N453, u2_N456, u2_N457, u2_N460, u2_N463, u2_N464, u2_N465, 
        u2_N467, u2_N470, u2_N471, u2_N473, u2_N475, u2_N477, u2_N478, u2_N48, u2_N49, 
        u2_N5, u2_N54, u2_N59, u2_N62, u2_N8, u2_uk_n1087, u2_uk_n1090, u2_uk_n11, u2_uk_n110, 
        u2_uk_n1102, u2_uk_n1145, u2_uk_n1146, u2_uk_n1148, u2_uk_n1150, u2_uk_n1155, u2_uk_n1161, u2_uk_n1162, u2_uk_n1168, 
        u2_uk_n1185, u2_uk_n129, u2_uk_n147, u2_uk_n163, u2_uk_n188, u2_uk_n191, u2_uk_n207, u2_uk_n298, u2_uk_n366, 
        u2_uk_n60, u2_uk_n656;
  wire u0_K10_21, u0_K10_22, u0_K10_23, u0_K10_24, u0_K11_10, u0_K11_11, u0_K11_12, u0_K11_13, u0_K11_14, 
       u0_K11_15, u0_K11_16, u0_K11_17, u0_K11_18, u0_K11_19, u0_K11_20, u0_K11_22, u0_K11_23, u0_K11_24, 
       u0_K11_31, u0_K11_32, u0_K11_33, u0_K11_34, u0_K11_35, u0_K11_36, u0_K11_38, u0_K11_39, u0_K11_40, 
       u0_K11_41, u0_K11_42, u0_K11_43, u0_K11_44, u0_K11_45, u0_K11_46, u0_K11_47, u0_K11_7, u0_K11_8, 
       u0_K11_9, u0_K13_10, u0_K13_11, u0_K13_12, u0_K13_13, u0_K13_14, u0_K13_15, u0_K13_16, u0_K13_17, 
       u0_K13_18, u0_K13_19, u0_K13_20, u0_K13_21, u0_K13_22, u0_K13_23, u0_K13_24, u0_K13_7, u0_K13_8, 
       u0_K13_9, u0_K15_25, u0_K15_26, u0_K15_27, u0_K15_28, u0_K15_29, u0_K15_30, u0_K2_1, u0_K2_10, 
       u0_K2_2, u0_K2_26, u0_K2_27, u0_K2_28, u0_K2_29, u0_K2_3, u0_K2_31, u0_K2_32, u0_K2_33, 
       u0_K2_36, u0_K2_37, u0_K2_38, u0_K2_39, u0_K2_40, u0_K2_41, u0_K2_42, u0_K2_7, u0_K2_9, 
       u0_K3_1, u0_K3_11, u0_K3_13, u0_K3_16, u0_K3_2, u0_K3_20, u0_K3_21, u0_K3_22, u0_K3_24, 
       u0_K3_3, u0_K3_4, u0_K3_6, u0_K3_7, u0_K3_8, u0_K3_9, u0_K4_1, u0_K4_10, u0_K4_11, 
       u0_K4_12, u0_K4_13, u0_K4_14, u0_K4_15, u0_K4_16, u0_K4_17, u0_K4_18, u0_K4_19, u0_K4_2, 
       u0_K4_20, u0_K4_21, u0_K4_22, u0_K4_23, u0_K4_25, u0_K4_26, u0_K4_29, u0_K4_3, u0_K4_30, 
       u0_K4_31, u0_K4_32, u0_K4_33, u0_K4_34, u0_K4_36, u0_K4_4, u0_K4_5, u0_K4_7, u0_K4_8, 
       u0_K4_9, u0_K6_21, u0_K6_25, u0_K6_26, u0_K6_28, u0_K6_29, u0_K6_30, u0_K6_31, u0_K6_32, 
       u0_K6_33, u0_K6_34, u0_K6_35, u0_K6_36, u0_K6_37, u0_K6_38, u0_K6_39, u0_K6_40, u0_K6_42, 
       u0_K7_1, u0_K7_10, u0_K7_11, u0_K7_12, u0_K7_13, u0_K7_14, u0_K7_15, u0_K7_16, u0_K7_17, 
       u0_K7_18, u0_K7_19, u0_K7_20, u0_K7_21, u0_K7_24, u0_K7_3, u0_K7_4, u0_K7_43, u0_K7_44, 
       u0_K7_45, u0_K7_46, u0_K7_47, u0_K7_48, u0_K7_5, u0_K7_6, u0_K7_7, u0_K7_8, u0_K7_9, 
       u0_K8_43, u0_K8_44, u0_K8_46, u0_K8_47, u0_K8_48, u0_out10_1, u0_out10_10, u0_out10_11, u0_out10_12, 
       u0_out10_13, u0_out10_15, u0_out10_16, u0_out10_18, u0_out10_19, u0_out10_2, u0_out10_20, u0_out10_21, u0_out10_22, 
       u0_out10_24, u0_out10_26, u0_out10_27, u0_out10_28, u0_out10_29, u0_out10_30, u0_out10_32, u0_out10_4, u0_out10_5, 
       u0_out10_6, u0_out10_7, u0_out12_1, u0_out12_10, u0_out12_13, u0_out12_16, u0_out12_18, u0_out12_2, u0_out12_20, 
       u0_out12_24, u0_out12_26, u0_out12_28, u0_out12_30, u0_out12_6, u0_out14_14, u0_out14_25, u0_out14_3, u0_out14_8, 
       u0_out1_11, u0_out1_12, u0_out1_13, u0_out1_14, u0_out1_17, u0_out1_18, u0_out1_19, u0_out1_2, u0_out1_22, 
       u0_out1_23, u0_out1_25, u0_out1_28, u0_out1_29, u0_out1_3, u0_out1_31, u0_out1_32, u0_out1_4, u0_out1_7, 
       u0_out1_8, u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_13, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_2, 
       u0_out2_20, u0_out2_23, u0_out2_24, u0_out2_26, u0_out2_28, u0_out2_30, u0_out2_31, u0_out2_6, u0_out2_9, 
       u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_13, u0_out3_14, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, 
       u0_out3_2, u0_out3_20, u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_28, u0_out3_29, u0_out3_3, 
       u0_out3_30, u0_out3_31, u0_out3_4, u0_out3_6, u0_out3_8, u0_out3_9, u0_out5_1, u0_out5_10, u0_out5_11, 
       u0_out5_12, u0_out5_14, u0_out5_19, u0_out5_20, u0_out5_22, u0_out5_25, u0_out5_26, u0_out5_29, u0_out5_3, 
       u0_out5_32, u0_out5_4, u0_out5_7, u0_out5_8, u0_out6_1, u0_out6_10, u0_out6_13, u0_out6_15, u0_out6_16, 
       u0_out6_17, u0_out6_18, u0_out6_2, u0_out6_20, u0_out6_21, u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_27, 
       u0_out6_28, u0_out6_30, u0_out6_31, u0_out6_5, u0_out6_6, u0_out6_9, u0_out7_15, u0_out7_21, u0_out7_27, 
       u0_out7_5, u0_out9_1, u0_out9_10, u0_out9_20, u0_out9_26, u0_u10_X_10, u0_u10_X_11, u0_u10_X_12, u0_u10_X_13, 
       u0_u10_X_14, u0_u10_X_15, u0_u10_X_16, u0_u10_X_17, u0_u10_X_18, u0_u10_X_19, u0_u10_X_20, u0_u10_X_21, u0_u10_X_22, 
       u0_u10_X_23, u0_u10_X_24, u0_u10_X_31, u0_u10_X_32, u0_u10_X_33, u0_u10_X_34, u0_u10_X_35, u0_u10_X_36, u0_u10_X_37, 
       u0_u10_X_38, u0_u10_X_39, u0_u10_X_40, u0_u10_X_41, u0_u10_X_42, u0_u10_X_43, u0_u10_X_44, u0_u10_X_45, u0_u10_X_46, 
       u0_u10_X_47, u0_u10_X_48, u0_u10_X_7, u0_u10_X_8, u0_u10_X_9, u0_u10_u1_n100, u0_u10_u1_n101, u0_u10_u1_n102, u0_u10_u1_n103, 
       u0_u10_u1_n104, u0_u10_u1_n105, u0_u10_u1_n106, u0_u10_u1_n107, u0_u10_u1_n108, u0_u10_u1_n109, u0_u10_u1_n110, u0_u10_u1_n111, u0_u10_u1_n112, 
       u0_u10_u1_n113, u0_u10_u1_n114, u0_u10_u1_n115, u0_u10_u1_n116, u0_u10_u1_n117, u0_u10_u1_n118, u0_u10_u1_n119, u0_u10_u1_n120, u0_u10_u1_n121, 
       u0_u10_u1_n122, u0_u10_u1_n123, u0_u10_u1_n124, u0_u10_u1_n125, u0_u10_u1_n126, u0_u10_u1_n127, u0_u10_u1_n128, u0_u10_u1_n129, u0_u10_u1_n130, 
       u0_u10_u1_n131, u0_u10_u1_n132, u0_u10_u1_n133, u0_u10_u1_n134, u0_u10_u1_n135, u0_u10_u1_n136, u0_u10_u1_n137, u0_u10_u1_n138, u0_u10_u1_n139, 
       u0_u10_u1_n140, u0_u10_u1_n141, u0_u10_u1_n142, u0_u10_u1_n143, u0_u10_u1_n144, u0_u10_u1_n145, u0_u10_u1_n146, u0_u10_u1_n147, u0_u10_u1_n148, 
       u0_u10_u1_n149, u0_u10_u1_n150, u0_u10_u1_n151, u0_u10_u1_n152, u0_u10_u1_n153, u0_u10_u1_n154, u0_u10_u1_n155, u0_u10_u1_n156, u0_u10_u1_n157, 
       u0_u10_u1_n158, u0_u10_u1_n159, u0_u10_u1_n160, u0_u10_u1_n161, u0_u10_u1_n162, u0_u10_u1_n163, u0_u10_u1_n164, u0_u10_u1_n165, u0_u10_u1_n166, 
       u0_u10_u1_n167, u0_u10_u1_n168, u0_u10_u1_n169, u0_u10_u1_n170, u0_u10_u1_n171, u0_u10_u1_n172, u0_u10_u1_n173, u0_u10_u1_n174, u0_u10_u1_n175, 
       u0_u10_u1_n176, u0_u10_u1_n177, u0_u10_u1_n178, u0_u10_u1_n179, u0_u10_u1_n180, u0_u10_u1_n181, u0_u10_u1_n182, u0_u10_u1_n183, u0_u10_u1_n184, 
       u0_u10_u1_n185, u0_u10_u1_n186, u0_u10_u1_n187, u0_u10_u1_n188, u0_u10_u1_n95, u0_u10_u1_n96, u0_u10_u1_n97, u0_u10_u1_n98, u0_u10_u1_n99, 
       u0_u10_u2_n100, u0_u10_u2_n101, u0_u10_u2_n102, u0_u10_u2_n103, u0_u10_u2_n104, u0_u10_u2_n105, u0_u10_u2_n106, u0_u10_u2_n107, u0_u10_u2_n108, 
       u0_u10_u2_n109, u0_u10_u2_n110, u0_u10_u2_n111, u0_u10_u2_n112, u0_u10_u2_n113, u0_u10_u2_n114, u0_u10_u2_n115, u0_u10_u2_n116, u0_u10_u2_n117, 
       u0_u10_u2_n118, u0_u10_u2_n119, u0_u10_u2_n120, u0_u10_u2_n121, u0_u10_u2_n122, u0_u10_u2_n123, u0_u10_u2_n124, u0_u10_u2_n125, u0_u10_u2_n126, 
       u0_u10_u2_n127, u0_u10_u2_n128, u0_u10_u2_n129, u0_u10_u2_n130, u0_u10_u2_n131, u0_u10_u2_n132, u0_u10_u2_n133, u0_u10_u2_n134, u0_u10_u2_n135, 
       u0_u10_u2_n136, u0_u10_u2_n137, u0_u10_u2_n138, u0_u10_u2_n139, u0_u10_u2_n140, u0_u10_u2_n141, u0_u10_u2_n142, u0_u10_u2_n143, u0_u10_u2_n144, 
       u0_u10_u2_n145, u0_u10_u2_n146, u0_u10_u2_n147, u0_u10_u2_n148, u0_u10_u2_n149, u0_u10_u2_n150, u0_u10_u2_n151, u0_u10_u2_n152, u0_u10_u2_n153, 
       u0_u10_u2_n154, u0_u10_u2_n155, u0_u10_u2_n156, u0_u10_u2_n157, u0_u10_u2_n158, u0_u10_u2_n159, u0_u10_u2_n160, u0_u10_u2_n161, u0_u10_u2_n162, 
       u0_u10_u2_n163, u0_u10_u2_n164, u0_u10_u2_n165, u0_u10_u2_n166, u0_u10_u2_n167, u0_u10_u2_n168, u0_u10_u2_n169, u0_u10_u2_n170, u0_u10_u2_n171, 
       u0_u10_u2_n172, u0_u10_u2_n173, u0_u10_u2_n174, u0_u10_u2_n175, u0_u10_u2_n176, u0_u10_u2_n177, u0_u10_u2_n178, u0_u10_u2_n179, u0_u10_u2_n180, 
       u0_u10_u2_n181, u0_u10_u2_n182, u0_u10_u2_n183, u0_u10_u2_n184, u0_u10_u2_n185, u0_u10_u2_n186, u0_u10_u2_n187, u0_u10_u2_n188, u0_u10_u2_n95, 
       u0_u10_u2_n96, u0_u10_u2_n97, u0_u10_u2_n98, u0_u10_u2_n99, u0_u10_u3_n100, u0_u10_u3_n101, u0_u10_u3_n102, u0_u10_u3_n103, u0_u10_u3_n104, 
       u0_u10_u3_n105, u0_u10_u3_n106, u0_u10_u3_n107, u0_u10_u3_n108, u0_u10_u3_n109, u0_u10_u3_n110, u0_u10_u3_n111, u0_u10_u3_n112, u0_u10_u3_n113, 
       u0_u10_u3_n114, u0_u10_u3_n115, u0_u10_u3_n116, u0_u10_u3_n117, u0_u10_u3_n118, u0_u10_u3_n119, u0_u10_u3_n120, u0_u10_u3_n121, u0_u10_u3_n122, 
       u0_u10_u3_n123, u0_u10_u3_n124, u0_u10_u3_n125, u0_u10_u3_n126, u0_u10_u3_n127, u0_u10_u3_n128, u0_u10_u3_n129, u0_u10_u3_n130, u0_u10_u3_n131, 
       u0_u10_u3_n132, u0_u10_u3_n133, u0_u10_u3_n134, u0_u10_u3_n135, u0_u10_u3_n136, u0_u10_u3_n137, u0_u10_u3_n138, u0_u10_u3_n139, u0_u10_u3_n140, 
       u0_u10_u3_n141, u0_u10_u3_n142, u0_u10_u3_n143, u0_u10_u3_n144, u0_u10_u3_n145, u0_u10_u3_n146, u0_u10_u3_n147, u0_u10_u3_n148, u0_u10_u3_n149, 
       u0_u10_u3_n150, u0_u10_u3_n151, u0_u10_u3_n152, u0_u10_u3_n153, u0_u10_u3_n154, u0_u10_u3_n155, u0_u10_u3_n156, u0_u10_u3_n157, u0_u10_u3_n158, 
       u0_u10_u3_n159, u0_u10_u3_n160, u0_u10_u3_n161, u0_u10_u3_n162, u0_u10_u3_n163, u0_u10_u3_n164, u0_u10_u3_n165, u0_u10_u3_n166, u0_u10_u3_n167, 
       u0_u10_u3_n168, u0_u10_u3_n169, u0_u10_u3_n170, u0_u10_u3_n171, u0_u10_u3_n172, u0_u10_u3_n173, u0_u10_u3_n174, u0_u10_u3_n175, u0_u10_u3_n176, 
       u0_u10_u3_n177, u0_u10_u3_n178, u0_u10_u3_n179, u0_u10_u3_n180, u0_u10_u3_n181, u0_u10_u3_n182, u0_u10_u3_n183, u0_u10_u3_n184, u0_u10_u3_n185, 
       u0_u10_u3_n186, u0_u10_u3_n94, u0_u10_u3_n95, u0_u10_u3_n96, u0_u10_u3_n97, u0_u10_u3_n98, u0_u10_u3_n99, u0_u10_u5_n100, u0_u10_u5_n101, 
       u0_u10_u5_n102, u0_u10_u5_n103, u0_u10_u5_n104, u0_u10_u5_n105, u0_u10_u5_n106, u0_u10_u5_n107, u0_u10_u5_n108, u0_u10_u5_n109, u0_u10_u5_n110, 
       u0_u10_u5_n111, u0_u10_u5_n112, u0_u10_u5_n113, u0_u10_u5_n114, u0_u10_u5_n115, u0_u10_u5_n116, u0_u10_u5_n117, u0_u10_u5_n118, u0_u10_u5_n119, 
       u0_u10_u5_n120, u0_u10_u5_n121, u0_u10_u5_n122, u0_u10_u5_n123, u0_u10_u5_n124, u0_u10_u5_n125, u0_u10_u5_n126, u0_u10_u5_n127, u0_u10_u5_n128, 
       u0_u10_u5_n129, u0_u10_u5_n130, u0_u10_u5_n131, u0_u10_u5_n132, u0_u10_u5_n133, u0_u10_u5_n134, u0_u10_u5_n135, u0_u10_u5_n136, u0_u10_u5_n137, 
       u0_u10_u5_n138, u0_u10_u5_n139, u0_u10_u5_n140, u0_u10_u5_n141, u0_u10_u5_n142, u0_u10_u5_n143, u0_u10_u5_n144, u0_u10_u5_n145, u0_u10_u5_n146, 
       u0_u10_u5_n147, u0_u10_u5_n148, u0_u10_u5_n149, u0_u10_u5_n150, u0_u10_u5_n151, u0_u10_u5_n152, u0_u10_u5_n153, u0_u10_u5_n154, u0_u10_u5_n155, 
       u0_u10_u5_n156, u0_u10_u5_n157, u0_u10_u5_n158, u0_u10_u5_n159, u0_u10_u5_n160, u0_u10_u5_n161, u0_u10_u5_n162, u0_u10_u5_n163, u0_u10_u5_n164, 
       u0_u10_u5_n165, u0_u10_u5_n166, u0_u10_u5_n167, u0_u10_u5_n168, u0_u10_u5_n169, u0_u10_u5_n170, u0_u10_u5_n171, u0_u10_u5_n172, u0_u10_u5_n173, 
       u0_u10_u5_n174, u0_u10_u5_n175, u0_u10_u5_n176, u0_u10_u5_n177, u0_u10_u5_n178, u0_u10_u5_n179, u0_u10_u5_n180, u0_u10_u5_n181, u0_u10_u5_n182, 
       u0_u10_u5_n183, u0_u10_u5_n184, u0_u10_u5_n185, u0_u10_u5_n186, u0_u10_u5_n187, u0_u10_u5_n188, u0_u10_u5_n189, u0_u10_u5_n190, u0_u10_u5_n191, 
       u0_u10_u5_n192, u0_u10_u5_n193, u0_u10_u5_n194, u0_u10_u5_n195, u0_u10_u5_n196, u0_u10_u5_n99, u0_u10_u6_n100, u0_u10_u6_n101, u0_u10_u6_n102, 
       u0_u10_u6_n103, u0_u10_u6_n104, u0_u10_u6_n105, u0_u10_u6_n106, u0_u10_u6_n107, u0_u10_u6_n108, u0_u10_u6_n109, u0_u10_u6_n110, u0_u10_u6_n111, 
       u0_u10_u6_n112, u0_u10_u6_n113, u0_u10_u6_n114, u0_u10_u6_n115, u0_u10_u6_n116, u0_u10_u6_n117, u0_u10_u6_n118, u0_u10_u6_n119, u0_u10_u6_n120, 
       u0_u10_u6_n121, u0_u10_u6_n122, u0_u10_u6_n123, u0_u10_u6_n124, u0_u10_u6_n125, u0_u10_u6_n126, u0_u10_u6_n127, u0_u10_u6_n128, u0_u10_u6_n129, 
       u0_u10_u6_n130, u0_u10_u6_n131, u0_u10_u6_n132, u0_u10_u6_n133, u0_u10_u6_n134, u0_u10_u6_n135, u0_u10_u6_n136, u0_u10_u6_n137, u0_u10_u6_n138, 
       u0_u10_u6_n139, u0_u10_u6_n140, u0_u10_u6_n141, u0_u10_u6_n142, u0_u10_u6_n143, u0_u10_u6_n144, u0_u10_u6_n145, u0_u10_u6_n146, u0_u10_u6_n147, 
       u0_u10_u6_n148, u0_u10_u6_n149, u0_u10_u6_n150, u0_u10_u6_n151, u0_u10_u6_n152, u0_u10_u6_n153, u0_u10_u6_n154, u0_u10_u6_n155, u0_u10_u6_n156, 
       u0_u10_u6_n157, u0_u10_u6_n158, u0_u10_u6_n159, u0_u10_u6_n160, u0_u10_u6_n161, u0_u10_u6_n162, u0_u10_u6_n163, u0_u10_u6_n164, u0_u10_u6_n165, 
       u0_u10_u6_n166, u0_u10_u6_n167, u0_u10_u6_n168, u0_u10_u6_n169, u0_u10_u6_n170, u0_u10_u6_n171, u0_u10_u6_n172, u0_u10_u6_n173, u0_u10_u6_n174, 
       u0_u10_u6_n88, u0_u10_u6_n89, u0_u10_u6_n90, u0_u10_u6_n91, u0_u10_u6_n92, u0_u10_u6_n93, u0_u10_u6_n94, u0_u10_u6_n95, u0_u10_u6_n96, 
       u0_u10_u6_n97, u0_u10_u6_n98, u0_u10_u6_n99, u0_u10_u7_n100, u0_u10_u7_n101, u0_u10_u7_n102, u0_u10_u7_n103, u0_u10_u7_n104, u0_u10_u7_n105, 
       u0_u10_u7_n106, u0_u10_u7_n107, u0_u10_u7_n108, u0_u10_u7_n109, u0_u10_u7_n110, u0_u10_u7_n111, u0_u10_u7_n112, u0_u10_u7_n113, u0_u10_u7_n114, 
       u0_u10_u7_n115, u0_u10_u7_n116, u0_u10_u7_n117, u0_u10_u7_n118, u0_u10_u7_n119, u0_u10_u7_n120, u0_u10_u7_n121, u0_u10_u7_n122, u0_u10_u7_n123, 
       u0_u10_u7_n124, u0_u10_u7_n125, u0_u10_u7_n126, u0_u10_u7_n127, u0_u10_u7_n128, u0_u10_u7_n129, u0_u10_u7_n130, u0_u10_u7_n131, u0_u10_u7_n132, 
       u0_u10_u7_n133, u0_u10_u7_n134, u0_u10_u7_n135, u0_u10_u7_n136, u0_u10_u7_n137, u0_u10_u7_n138, u0_u10_u7_n139, u0_u10_u7_n140, u0_u10_u7_n141, 
       u0_u10_u7_n142, u0_u10_u7_n143, u0_u10_u7_n144, u0_u10_u7_n145, u0_u10_u7_n146, u0_u10_u7_n147, u0_u10_u7_n148, u0_u10_u7_n149, u0_u10_u7_n150, 
       u0_u10_u7_n151, u0_u10_u7_n152, u0_u10_u7_n153, u0_u10_u7_n154, u0_u10_u7_n155, u0_u10_u7_n156, u0_u10_u7_n157, u0_u10_u7_n158, u0_u10_u7_n159, 
       u0_u10_u7_n160, u0_u10_u7_n161, u0_u10_u7_n162, u0_u10_u7_n163, u0_u10_u7_n164, u0_u10_u7_n165, u0_u10_u7_n166, u0_u10_u7_n167, u0_u10_u7_n168, 
       u0_u10_u7_n169, u0_u10_u7_n170, u0_u10_u7_n171, u0_u10_u7_n172, u0_u10_u7_n173, u0_u10_u7_n174, u0_u10_u7_n175, u0_u10_u7_n176, u0_u10_u7_n177, 
       u0_u10_u7_n178, u0_u10_u7_n179, u0_u10_u7_n180, u0_u10_u7_n91, u0_u10_u7_n92, u0_u10_u7_n93, u0_u10_u7_n94, u0_u10_u7_n95, u0_u10_u7_n96, 
       u0_u10_u7_n97, u0_u10_u7_n98, u0_u10_u7_n99, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, u0_u12_X_15, 
       u0_u12_X_16, u0_u12_X_17, u0_u12_X_18, u0_u12_X_19, u0_u12_X_20, u0_u12_X_21, u0_u12_X_22, u0_u12_X_23, u0_u12_X_24, 
       u0_u12_X_7, u0_u12_X_8, u0_u12_X_9, u0_u12_u1_n100, u0_u12_u1_n101, u0_u12_u1_n102, u0_u12_u1_n103, u0_u12_u1_n104, u0_u12_u1_n105, 
       u0_u12_u1_n106, u0_u12_u1_n107, u0_u12_u1_n108, u0_u12_u1_n109, u0_u12_u1_n110, u0_u12_u1_n111, u0_u12_u1_n112, u0_u12_u1_n113, u0_u12_u1_n114, 
       u0_u12_u1_n115, u0_u12_u1_n116, u0_u12_u1_n117, u0_u12_u1_n118, u0_u12_u1_n119, u0_u12_u1_n120, u0_u12_u1_n121, u0_u12_u1_n122, u0_u12_u1_n123, 
       u0_u12_u1_n124, u0_u12_u1_n125, u0_u12_u1_n126, u0_u12_u1_n127, u0_u12_u1_n128, u0_u12_u1_n129, u0_u12_u1_n130, u0_u12_u1_n131, u0_u12_u1_n132, 
       u0_u12_u1_n133, u0_u12_u1_n134, u0_u12_u1_n135, u0_u12_u1_n136, u0_u12_u1_n137, u0_u12_u1_n138, u0_u12_u1_n139, u0_u12_u1_n140, u0_u12_u1_n141, 
       u0_u12_u1_n142, u0_u12_u1_n143, u0_u12_u1_n144, u0_u12_u1_n145, u0_u12_u1_n146, u0_u12_u1_n147, u0_u12_u1_n148, u0_u12_u1_n149, u0_u12_u1_n150, 
       u0_u12_u1_n151, u0_u12_u1_n152, u0_u12_u1_n153, u0_u12_u1_n154, u0_u12_u1_n155, u0_u12_u1_n156, u0_u12_u1_n157, u0_u12_u1_n158, u0_u12_u1_n159, 
       u0_u12_u1_n160, u0_u12_u1_n161, u0_u12_u1_n162, u0_u12_u1_n163, u0_u12_u1_n164, u0_u12_u1_n165, u0_u12_u1_n166, u0_u12_u1_n167, u0_u12_u1_n168, 
       u0_u12_u1_n169, u0_u12_u1_n170, u0_u12_u1_n171, u0_u12_u1_n172, u0_u12_u1_n173, u0_u12_u1_n174, u0_u12_u1_n175, u0_u12_u1_n176, u0_u12_u1_n177, 
       u0_u12_u1_n178, u0_u12_u1_n179, u0_u12_u1_n180, u0_u12_u1_n181, u0_u12_u1_n182, u0_u12_u1_n183, u0_u12_u1_n184, u0_u12_u1_n185, u0_u12_u1_n186, 
       u0_u12_u1_n187, u0_u12_u1_n188, u0_u12_u1_n95, u0_u12_u1_n96, u0_u12_u1_n97, u0_u12_u1_n98, u0_u12_u1_n99, u0_u12_u2_n100, u0_u12_u2_n101, 
       u0_u12_u2_n102, u0_u12_u2_n103, u0_u12_u2_n104, u0_u12_u2_n105, u0_u12_u2_n106, u0_u12_u2_n107, u0_u12_u2_n108, u0_u12_u2_n109, u0_u12_u2_n110, 
       u0_u12_u2_n111, u0_u12_u2_n112, u0_u12_u2_n113, u0_u12_u2_n114, u0_u12_u2_n115, u0_u12_u2_n116, u0_u12_u2_n117, u0_u12_u2_n118, u0_u12_u2_n119, 
       u0_u12_u2_n120, u0_u12_u2_n121, u0_u12_u2_n122, u0_u12_u2_n123, u0_u12_u2_n124, u0_u12_u2_n125, u0_u12_u2_n126, u0_u12_u2_n127, u0_u12_u2_n128, 
       u0_u12_u2_n129, u0_u12_u2_n130, u0_u12_u2_n131, u0_u12_u2_n132, u0_u12_u2_n133, u0_u12_u2_n134, u0_u12_u2_n135, u0_u12_u2_n136, u0_u12_u2_n137, 
       u0_u12_u2_n138, u0_u12_u2_n139, u0_u12_u2_n140, u0_u12_u2_n141, u0_u12_u2_n142, u0_u12_u2_n143, u0_u12_u2_n144, u0_u12_u2_n145, u0_u12_u2_n146, 
       u0_u12_u2_n147, u0_u12_u2_n148, u0_u12_u2_n149, u0_u12_u2_n150, u0_u12_u2_n151, u0_u12_u2_n152, u0_u12_u2_n153, u0_u12_u2_n154, u0_u12_u2_n155, 
       u0_u12_u2_n156, u0_u12_u2_n157, u0_u12_u2_n158, u0_u12_u2_n159, u0_u12_u2_n160, u0_u12_u2_n161, u0_u12_u2_n162, u0_u12_u2_n163, u0_u12_u2_n164, 
       u0_u12_u2_n165, u0_u12_u2_n166, u0_u12_u2_n167, u0_u12_u2_n168, u0_u12_u2_n169, u0_u12_u2_n170, u0_u12_u2_n171, u0_u12_u2_n172, u0_u12_u2_n173, 
       u0_u12_u2_n174, u0_u12_u2_n175, u0_u12_u2_n176, u0_u12_u2_n177, u0_u12_u2_n178, u0_u12_u2_n179, u0_u12_u2_n180, u0_u12_u2_n181, u0_u12_u2_n182, 
       u0_u12_u2_n183, u0_u12_u2_n184, u0_u12_u2_n185, u0_u12_u2_n186, u0_u12_u2_n187, u0_u12_u2_n188, u0_u12_u2_n95, u0_u12_u2_n96, u0_u12_u2_n97, 
       u0_u12_u2_n98, u0_u12_u2_n99, u0_u12_u3_n100, u0_u12_u3_n101, u0_u12_u3_n102, u0_u12_u3_n103, u0_u12_u3_n104, u0_u12_u3_n105, u0_u12_u3_n106, 
       u0_u12_u3_n107, u0_u12_u3_n108, u0_u12_u3_n109, u0_u12_u3_n110, u0_u12_u3_n111, u0_u12_u3_n112, u0_u12_u3_n113, u0_u12_u3_n114, u0_u12_u3_n115, 
       u0_u12_u3_n116, u0_u12_u3_n117, u0_u12_u3_n118, u0_u12_u3_n119, u0_u12_u3_n120, u0_u12_u3_n121, u0_u12_u3_n122, u0_u12_u3_n123, u0_u12_u3_n124, 
       u0_u12_u3_n125, u0_u12_u3_n126, u0_u12_u3_n127, u0_u12_u3_n128, u0_u12_u3_n129, u0_u12_u3_n130, u0_u12_u3_n131, u0_u12_u3_n132, u0_u12_u3_n133, 
       u0_u12_u3_n134, u0_u12_u3_n135, u0_u12_u3_n136, u0_u12_u3_n137, u0_u12_u3_n138, u0_u12_u3_n139, u0_u12_u3_n140, u0_u12_u3_n141, u0_u12_u3_n142, 
       u0_u12_u3_n143, u0_u12_u3_n144, u0_u12_u3_n145, u0_u12_u3_n146, u0_u12_u3_n147, u0_u12_u3_n148, u0_u12_u3_n149, u0_u12_u3_n150, u0_u12_u3_n151, 
       u0_u12_u3_n152, u0_u12_u3_n153, u0_u12_u3_n154, u0_u12_u3_n155, u0_u12_u3_n156, u0_u12_u3_n157, u0_u12_u3_n158, u0_u12_u3_n159, u0_u12_u3_n160, 
       u0_u12_u3_n161, u0_u12_u3_n162, u0_u12_u3_n163, u0_u12_u3_n164, u0_u12_u3_n165, u0_u12_u3_n166, u0_u12_u3_n167, u0_u12_u3_n168, u0_u12_u3_n169, 
       u0_u12_u3_n170, u0_u12_u3_n171, u0_u12_u3_n172, u0_u12_u3_n173, u0_u12_u3_n174, u0_u12_u3_n175, u0_u12_u3_n176, u0_u12_u3_n177, u0_u12_u3_n178, 
       u0_u12_u3_n179, u0_u12_u3_n180, u0_u12_u3_n181, u0_u12_u3_n182, u0_u12_u3_n183, u0_u12_u3_n184, u0_u12_u3_n185, u0_u12_u3_n186, u0_u12_u3_n94, 
       u0_u12_u3_n95, u0_u12_u3_n96, u0_u12_u3_n97, u0_u12_u3_n98, u0_u12_u3_n99, u0_u14_X_25, u0_u14_X_26, u0_u14_X_27, u0_u14_X_28, 
       u0_u14_X_29, u0_u14_X_30, u0_u14_u4_n100, u0_u14_u4_n101, u0_u14_u4_n102, u0_u14_u4_n103, u0_u14_u4_n104, u0_u14_u4_n105, u0_u14_u4_n106, 
       u0_u14_u4_n107, u0_u14_u4_n108, u0_u14_u4_n109, u0_u14_u4_n110, u0_u14_u4_n111, u0_u14_u4_n112, u0_u14_u4_n113, u0_u14_u4_n114, u0_u14_u4_n115, 
       u0_u14_u4_n116, u0_u14_u4_n117, u0_u14_u4_n118, u0_u14_u4_n119, u0_u14_u4_n120, u0_u14_u4_n121, u0_u14_u4_n122, u0_u14_u4_n123, u0_u14_u4_n124, 
       u0_u14_u4_n125, u0_u14_u4_n126, u0_u14_u4_n127, u0_u14_u4_n128, u0_u14_u4_n129, u0_u14_u4_n130, u0_u14_u4_n131, u0_u14_u4_n132, u0_u14_u4_n133, 
       u0_u14_u4_n134, u0_u14_u4_n135, u0_u14_u4_n136, u0_u14_u4_n137, u0_u14_u4_n138, u0_u14_u4_n139, u0_u14_u4_n140, u0_u14_u4_n141, u0_u14_u4_n142, 
       u0_u14_u4_n143, u0_u14_u4_n144, u0_u14_u4_n145, u0_u14_u4_n146, u0_u14_u4_n147, u0_u14_u4_n148, u0_u14_u4_n149, u0_u14_u4_n150, u0_u14_u4_n151, 
       u0_u14_u4_n152, u0_u14_u4_n153, u0_u14_u4_n154, u0_u14_u4_n155, u0_u14_u4_n156, u0_u14_u4_n157, u0_u14_u4_n158, u0_u14_u4_n159, u0_u14_u4_n160, 
       u0_u14_u4_n161, u0_u14_u4_n162, u0_u14_u4_n163, u0_u14_u4_n164, u0_u14_u4_n165, u0_u14_u4_n166, u0_u14_u4_n167, u0_u14_u4_n168, u0_u14_u4_n169, 
       u0_u14_u4_n170, u0_u14_u4_n171, u0_u14_u4_n172, u0_u14_u4_n173, u0_u14_u4_n174, u0_u14_u4_n175, u0_u14_u4_n176, u0_u14_u4_n177, u0_u14_u4_n178, 
       u0_u14_u4_n179, u0_u14_u4_n180, u0_u14_u4_n181, u0_u14_u4_n182, u0_u14_u4_n183, u0_u14_u4_n184, u0_u14_u4_n185, u0_u14_u4_n186, u0_u14_u4_n94, 
       u0_u14_u4_n95, u0_u14_u4_n96, u0_u14_u4_n97, u0_u14_u4_n98, u0_u14_u4_n99, u0_u1_X_1, u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, 
       u0_u1_X_2, u0_u1_X_25, u0_u1_X_26, u0_u1_X_27, u0_u1_X_28, u0_u1_X_29, u0_u1_X_3, u0_u1_X_30, u0_u1_X_31, 
       u0_u1_X_32, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, u0_u1_X_36, u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_4, 
       u0_u1_X_40, u0_u1_X_41, u0_u1_X_42, u0_u1_X_5, u0_u1_X_6, u0_u1_X_7, u0_u1_X_8, u0_u1_X_9, u0_u1_u0_n100, 
       u0_u1_u0_n101, u0_u1_u0_n102, u0_u1_u0_n103, u0_u1_u0_n104, u0_u1_u0_n105, u0_u1_u0_n106, u0_u1_u0_n107, u0_u1_u0_n108, u0_u1_u0_n109, 
       u0_u1_u0_n110, u0_u1_u0_n111, u0_u1_u0_n112, u0_u1_u0_n113, u0_u1_u0_n114, u0_u1_u0_n115, u0_u1_u0_n116, u0_u1_u0_n117, u0_u1_u0_n118, 
       u0_u1_u0_n119, u0_u1_u0_n120, u0_u1_u0_n121, u0_u1_u0_n122, u0_u1_u0_n123, u0_u1_u0_n124, u0_u1_u0_n125, u0_u1_u0_n126, u0_u1_u0_n127, 
       u0_u1_u0_n128, u0_u1_u0_n129, u0_u1_u0_n130, u0_u1_u0_n131, u0_u1_u0_n132, u0_u1_u0_n133, u0_u1_u0_n134, u0_u1_u0_n135, u0_u1_u0_n136, 
       u0_u1_u0_n137, u0_u1_u0_n138, u0_u1_u0_n139, u0_u1_u0_n140, u0_u1_u0_n141, u0_u1_u0_n142, u0_u1_u0_n143, u0_u1_u0_n144, u0_u1_u0_n145, 
       u0_u1_u0_n146, u0_u1_u0_n147, u0_u1_u0_n148, u0_u1_u0_n149, u0_u1_u0_n150, u0_u1_u0_n151, u0_u1_u0_n152, u0_u1_u0_n153, u0_u1_u0_n154, 
       u0_u1_u0_n155, u0_u1_u0_n156, u0_u1_u0_n157, u0_u1_u0_n158, u0_u1_u0_n159, u0_u1_u0_n160, u0_u1_u0_n161, u0_u1_u0_n162, u0_u1_u0_n163, 
       u0_u1_u0_n164, u0_u1_u0_n165, u0_u1_u0_n166, u0_u1_u0_n167, u0_u1_u0_n168, u0_u1_u0_n169, u0_u1_u0_n170, u0_u1_u0_n171, u0_u1_u0_n172, 
       u0_u1_u0_n173, u0_u1_u0_n174, u0_u1_u0_n88, u0_u1_u0_n89, u0_u1_u0_n90, u0_u1_u0_n91, u0_u1_u0_n92, u0_u1_u0_n93, u0_u1_u0_n94, 
       u0_u1_u0_n95, u0_u1_u0_n96, u0_u1_u0_n97, u0_u1_u0_n98, u0_u1_u0_n99, u0_u1_u1_n100, u0_u1_u1_n101, u0_u1_u1_n102, u0_u1_u1_n103, 
       u0_u1_u1_n104, u0_u1_u1_n105, u0_u1_u1_n106, u0_u1_u1_n107, u0_u1_u1_n108, u0_u1_u1_n109, u0_u1_u1_n110, u0_u1_u1_n111, u0_u1_u1_n112, 
       u0_u1_u1_n113, u0_u1_u1_n114, u0_u1_u1_n115, u0_u1_u1_n116, u0_u1_u1_n117, u0_u1_u1_n118, u0_u1_u1_n119, u0_u1_u1_n120, u0_u1_u1_n121, 
       u0_u1_u1_n122, u0_u1_u1_n123, u0_u1_u1_n124, u0_u1_u1_n125, u0_u1_u1_n126, u0_u1_u1_n127, u0_u1_u1_n128, u0_u1_u1_n129, u0_u1_u1_n130, 
       u0_u1_u1_n131, u0_u1_u1_n132, u0_u1_u1_n133, u0_u1_u1_n134, u0_u1_u1_n135, u0_u1_u1_n136, u0_u1_u1_n137, u0_u1_u1_n138, u0_u1_u1_n139, 
       u0_u1_u1_n140, u0_u1_u1_n141, u0_u1_u1_n142, u0_u1_u1_n143, u0_u1_u1_n144, u0_u1_u1_n145, u0_u1_u1_n146, u0_u1_u1_n147, u0_u1_u1_n148, 
       u0_u1_u1_n149, u0_u1_u1_n150, u0_u1_u1_n151, u0_u1_u1_n152, u0_u1_u1_n153, u0_u1_u1_n154, u0_u1_u1_n155, u0_u1_u1_n156, u0_u1_u1_n157, 
       u0_u1_u1_n158, u0_u1_u1_n159, u0_u1_u1_n160, u0_u1_u1_n161, u0_u1_u1_n162, u0_u1_u1_n163, u0_u1_u1_n164, u0_u1_u1_n165, u0_u1_u1_n166, 
       u0_u1_u1_n167, u0_u1_u1_n168, u0_u1_u1_n169, u0_u1_u1_n170, u0_u1_u1_n171, u0_u1_u1_n172, u0_u1_u1_n173, u0_u1_u1_n174, u0_u1_u1_n175, 
       u0_u1_u1_n176, u0_u1_u1_n177, u0_u1_u1_n178, u0_u1_u1_n179, u0_u1_u1_n180, u0_u1_u1_n181, u0_u1_u1_n182, u0_u1_u1_n183, u0_u1_u1_n184, 
       u0_u1_u1_n185, u0_u1_u1_n186, u0_u1_u1_n187, u0_u1_u1_n188, u0_u1_u1_n95, u0_u1_u1_n96, u0_u1_u1_n97, u0_u1_u1_n98, u0_u1_u1_n99, 
       u0_u1_u4_n100, u0_u1_u4_n101, u0_u1_u4_n102, u0_u1_u4_n103, u0_u1_u4_n104, u0_u1_u4_n105, u0_u1_u4_n106, u0_u1_u4_n107, u0_u1_u4_n108, 
       u0_u1_u4_n109, u0_u1_u4_n110, u0_u1_u4_n111, u0_u1_u4_n112, u0_u1_u4_n113, u0_u1_u4_n114, u0_u1_u4_n115, u0_u1_u4_n116, u0_u1_u4_n117, 
       u0_u1_u4_n118, u0_u1_u4_n119, u0_u1_u4_n120, u0_u1_u4_n121, u0_u1_u4_n122, u0_u1_u4_n123, u0_u1_u4_n124, u0_u1_u4_n125, u0_u1_u4_n126, 
       u0_u1_u4_n127, u0_u1_u4_n128, u0_u1_u4_n129, u0_u1_u4_n130, u0_u1_u4_n131, u0_u1_u4_n132, u0_u1_u4_n133, u0_u1_u4_n134, u0_u1_u4_n135, 
       u0_u1_u4_n136, u0_u1_u4_n137, u0_u1_u4_n138, u0_u1_u4_n139, u0_u1_u4_n140, u0_u1_u4_n141, u0_u1_u4_n142, u0_u1_u4_n143, u0_u1_u4_n144, 
       u0_u1_u4_n145, u0_u1_u4_n146, u0_u1_u4_n147, u0_u1_u4_n148, u0_u1_u4_n149, u0_u1_u4_n150, u0_u1_u4_n151, u0_u1_u4_n152, u0_u1_u4_n153, 
       u0_u1_u4_n154, u0_u1_u4_n155, u0_u1_u4_n156, u0_u1_u4_n157, u0_u1_u4_n158, u0_u1_u4_n159, u0_u1_u4_n160, u0_u1_u4_n161, u0_u1_u4_n162, 
       u0_u1_u4_n163, u0_u1_u4_n164, u0_u1_u4_n165, u0_u1_u4_n166, u0_u1_u4_n167, u0_u1_u4_n168, u0_u1_u4_n169, u0_u1_u4_n170, u0_u1_u4_n171, 
       u0_u1_u4_n172, u0_u1_u4_n173, u0_u1_u4_n174, u0_u1_u4_n175, u0_u1_u4_n176, u0_u1_u4_n177, u0_u1_u4_n178, u0_u1_u4_n179, u0_u1_u4_n180, 
       u0_u1_u4_n181, u0_u1_u4_n182, u0_u1_u4_n183, u0_u1_u4_n184, u0_u1_u4_n185, u0_u1_u4_n186, u0_u1_u4_n94, u0_u1_u4_n95, u0_u1_u4_n96, 
       u0_u1_u4_n97, u0_u1_u4_n98, u0_u1_u4_n99, u0_u1_u5_n100, u0_u1_u5_n101, u0_u1_u5_n102, u0_u1_u5_n103, u0_u1_u5_n104, u0_u1_u5_n105, 
       u0_u1_u5_n106, u0_u1_u5_n107, u0_u1_u5_n108, u0_u1_u5_n109, u0_u1_u5_n110, u0_u1_u5_n111, u0_u1_u5_n112, u0_u1_u5_n113, u0_u1_u5_n114, 
       u0_u1_u5_n115, u0_u1_u5_n116, u0_u1_u5_n117, u0_u1_u5_n118, u0_u1_u5_n119, u0_u1_u5_n120, u0_u1_u5_n121, u0_u1_u5_n122, u0_u1_u5_n123, 
       u0_u1_u5_n124, u0_u1_u5_n125, u0_u1_u5_n126, u0_u1_u5_n127, u0_u1_u5_n128, u0_u1_u5_n129, u0_u1_u5_n130, u0_u1_u5_n131, u0_u1_u5_n132, 
       u0_u1_u5_n133, u0_u1_u5_n134, u0_u1_u5_n135, u0_u1_u5_n136, u0_u1_u5_n137, u0_u1_u5_n138, u0_u1_u5_n139, u0_u1_u5_n140, u0_u1_u5_n141, 
       u0_u1_u5_n142, u0_u1_u5_n143, u0_u1_u5_n144, u0_u1_u5_n145, u0_u1_u5_n146, u0_u1_u5_n147, u0_u1_u5_n148, u0_u1_u5_n149, u0_u1_u5_n150, 
       u0_u1_u5_n151, u0_u1_u5_n152, u0_u1_u5_n153, u0_u1_u5_n154, u0_u1_u5_n155, u0_u1_u5_n156, u0_u1_u5_n157, u0_u1_u5_n158, u0_u1_u5_n159, 
       u0_u1_u5_n160, u0_u1_u5_n161, u0_u1_u5_n162, u0_u1_u5_n163, u0_u1_u5_n164, u0_u1_u5_n165, u0_u1_u5_n166, u0_u1_u5_n167, u0_u1_u5_n168, 
       u0_u1_u5_n169, u0_u1_u5_n170, u0_u1_u5_n171, u0_u1_u5_n172, u0_u1_u5_n173, u0_u1_u5_n174, u0_u1_u5_n175, u0_u1_u5_n176, u0_u1_u5_n177, 
       u0_u1_u5_n178, u0_u1_u5_n179, u0_u1_u5_n180, u0_u1_u5_n181, u0_u1_u5_n182, u0_u1_u5_n183, u0_u1_u5_n184, u0_u1_u5_n185, u0_u1_u5_n186, 
       u0_u1_u5_n187, u0_u1_u5_n188, u0_u1_u5_n189, u0_u1_u5_n190, u0_u1_u5_n191, u0_u1_u5_n192, u0_u1_u5_n193, u0_u1_u5_n194, u0_u1_u5_n195, 
       u0_u1_u5_n196, u0_u1_u5_n99, u0_u1_u6_n100, u0_u1_u6_n101, u0_u1_u6_n102, u0_u1_u6_n103, u0_u1_u6_n104, u0_u1_u6_n105, u0_u1_u6_n106, 
       u0_u1_u6_n107, u0_u1_u6_n108, u0_u1_u6_n109, u0_u1_u6_n110, u0_u1_u6_n111, u0_u1_u6_n112, u0_u1_u6_n113, u0_u1_u6_n114, u0_u1_u6_n115, 
       u0_u1_u6_n116, u0_u1_u6_n117, u0_u1_u6_n118, u0_u1_u6_n119, u0_u1_u6_n120, u0_u1_u6_n121, u0_u1_u6_n122, u0_u1_u6_n123, u0_u1_u6_n124, 
       u0_u1_u6_n125, u0_u1_u6_n126, u0_u1_u6_n127, u0_u1_u6_n128, u0_u1_u6_n129, u0_u1_u6_n130, u0_u1_u6_n131, u0_u1_u6_n132, u0_u1_u6_n133, 
       u0_u1_u6_n134, u0_u1_u6_n135, u0_u1_u6_n136, u0_u1_u6_n137, u0_u1_u6_n138, u0_u1_u6_n139, u0_u1_u6_n140, u0_u1_u6_n141, u0_u1_u6_n142, 
       u0_u1_u6_n143, u0_u1_u6_n144, u0_u1_u6_n145, u0_u1_u6_n146, u0_u1_u6_n147, u0_u1_u6_n148, u0_u1_u6_n149, u0_u1_u6_n150, u0_u1_u6_n151, 
       u0_u1_u6_n152, u0_u1_u6_n153, u0_u1_u6_n154, u0_u1_u6_n155, u0_u1_u6_n156, u0_u1_u6_n157, u0_u1_u6_n158, u0_u1_u6_n159, u0_u1_u6_n160, 
       u0_u1_u6_n161, u0_u1_u6_n162, u0_u1_u6_n163, u0_u1_u6_n164, u0_u1_u6_n165, u0_u1_u6_n166, u0_u1_u6_n167, u0_u1_u6_n168, u0_u1_u6_n169, 
       u0_u1_u6_n170, u0_u1_u6_n171, u0_u1_u6_n172, u0_u1_u6_n173, u0_u1_u6_n174, u0_u1_u6_n88, u0_u1_u6_n89, u0_u1_u6_n90, u0_u1_u6_n91, 
       u0_u1_u6_n92, u0_u1_u6_n93, u0_u1_u6_n94, u0_u1_u6_n95, u0_u1_u6_n96, u0_u1_u6_n97, u0_u1_u6_n98, u0_u1_u6_n99, u0_u2_X_1, 
       u0_u2_X_10, u0_u2_X_11, u0_u2_X_12, u0_u2_X_13, u0_u2_X_14, u0_u2_X_15, u0_u2_X_16, u0_u2_X_17, u0_u2_X_18, 
       u0_u2_X_19, u0_u2_X_2, u0_u2_X_20, u0_u2_X_21, u0_u2_X_22, u0_u2_X_23, u0_u2_X_24, u0_u2_X_3, u0_u2_X_4, 
       u0_u2_X_5, u0_u2_X_6, u0_u2_X_7, u0_u2_X_8, u0_u2_X_9, u0_u2_u0_n100, u0_u2_u0_n101, u0_u2_u0_n102, u0_u2_u0_n103, 
       u0_u2_u0_n104, u0_u2_u0_n105, u0_u2_u0_n106, u0_u2_u0_n107, u0_u2_u0_n108, u0_u2_u0_n109, u0_u2_u0_n110, u0_u2_u0_n111, u0_u2_u0_n112, 
       u0_u2_u0_n113, u0_u2_u0_n114, u0_u2_u0_n115, u0_u2_u0_n116, u0_u2_u0_n117, u0_u2_u0_n118, u0_u2_u0_n119, u0_u2_u0_n120, u0_u2_u0_n121, 
       u0_u2_u0_n122, u0_u2_u0_n123, u0_u2_u0_n124, u0_u2_u0_n125, u0_u2_u0_n126, u0_u2_u0_n127, u0_u2_u0_n128, u0_u2_u0_n129, u0_u2_u0_n130, 
       u0_u2_u0_n131, u0_u2_u0_n132, u0_u2_u0_n133, u0_u2_u0_n134, u0_u2_u0_n135, u0_u2_u0_n136, u0_u2_u0_n137, u0_u2_u0_n138, u0_u2_u0_n139, 
       u0_u2_u0_n140, u0_u2_u0_n141, u0_u2_u0_n142, u0_u2_u0_n143, u0_u2_u0_n144, u0_u2_u0_n145, u0_u2_u0_n146, u0_u2_u0_n147, u0_u2_u0_n148, 
       u0_u2_u0_n149, u0_u2_u0_n150, u0_u2_u0_n151, u0_u2_u0_n152, u0_u2_u0_n153, u0_u2_u0_n154, u0_u2_u0_n155, u0_u2_u0_n156, u0_u2_u0_n157, 
       u0_u2_u0_n158, u0_u2_u0_n159, u0_u2_u0_n160, u0_u2_u0_n161, u0_u2_u0_n162, u0_u2_u0_n163, u0_u2_u0_n164, u0_u2_u0_n165, u0_u2_u0_n166, 
       u0_u2_u0_n167, u0_u2_u0_n168, u0_u2_u0_n169, u0_u2_u0_n170, u0_u2_u0_n171, u0_u2_u0_n172, u0_u2_u0_n173, u0_u2_u0_n174, u0_u2_u0_n88, 
       u0_u2_u0_n89, u0_u2_u0_n90, u0_u2_u0_n91, u0_u2_u0_n92, u0_u2_u0_n93, u0_u2_u0_n94, u0_u2_u0_n95, u0_u2_u0_n96, u0_u2_u0_n97, 
       u0_u2_u0_n98, u0_u2_u0_n99, u0_u2_u1_n100, u0_u2_u1_n101, u0_u2_u1_n102, u0_u2_u1_n103, u0_u2_u1_n104, u0_u2_u1_n105, u0_u2_u1_n106, 
       u0_u2_u1_n107, u0_u2_u1_n108, u0_u2_u1_n109, u0_u2_u1_n110, u0_u2_u1_n111, u0_u2_u1_n112, u0_u2_u1_n113, u0_u2_u1_n114, u0_u2_u1_n115, 
       u0_u2_u1_n116, u0_u2_u1_n117, u0_u2_u1_n118, u0_u2_u1_n119, u0_u2_u1_n120, u0_u2_u1_n121, u0_u2_u1_n122, u0_u2_u1_n123, u0_u2_u1_n124, 
       u0_u2_u1_n125, u0_u2_u1_n126, u0_u2_u1_n127, u0_u2_u1_n128, u0_u2_u1_n129, u0_u2_u1_n130, u0_u2_u1_n131, u0_u2_u1_n132, u0_u2_u1_n133, 
       u0_u2_u1_n134, u0_u2_u1_n135, u0_u2_u1_n136, u0_u2_u1_n137, u0_u2_u1_n138, u0_u2_u1_n139, u0_u2_u1_n140, u0_u2_u1_n141, u0_u2_u1_n142, 
       u0_u2_u1_n143, u0_u2_u1_n144, u0_u2_u1_n145, u0_u2_u1_n146, u0_u2_u1_n147, u0_u2_u1_n148, u0_u2_u1_n149, u0_u2_u1_n150, u0_u2_u1_n151, 
       u0_u2_u1_n152, u0_u2_u1_n153, u0_u2_u1_n154, u0_u2_u1_n155, u0_u2_u1_n156, u0_u2_u1_n157, u0_u2_u1_n158, u0_u2_u1_n159, u0_u2_u1_n160, 
       u0_u2_u1_n161, u0_u2_u1_n162, u0_u2_u1_n163, u0_u2_u1_n164, u0_u2_u1_n165, u0_u2_u1_n166, u0_u2_u1_n167, u0_u2_u1_n168, u0_u2_u1_n169, 
       u0_u2_u1_n170, u0_u2_u1_n171, u0_u2_u1_n172, u0_u2_u1_n173, u0_u2_u1_n174, u0_u2_u1_n175, u0_u2_u1_n176, u0_u2_u1_n177, u0_u2_u1_n178, 
       u0_u2_u1_n179, u0_u2_u1_n180, u0_u2_u1_n181, u0_u2_u1_n182, u0_u2_u1_n183, u0_u2_u1_n184, u0_u2_u1_n185, u0_u2_u1_n186, u0_u2_u1_n187, 
       u0_u2_u1_n188, u0_u2_u1_n95, u0_u2_u1_n96, u0_u2_u1_n97, u0_u2_u1_n98, u0_u2_u1_n99, u0_u2_u2_n100, u0_u2_u2_n101, u0_u2_u2_n102, 
       u0_u2_u2_n103, u0_u2_u2_n104, u0_u2_u2_n105, u0_u2_u2_n106, u0_u2_u2_n107, u0_u2_u2_n108, u0_u2_u2_n109, u0_u2_u2_n110, u0_u2_u2_n111, 
       u0_u2_u2_n112, u0_u2_u2_n113, u0_u2_u2_n114, u0_u2_u2_n115, u0_u2_u2_n116, u0_u2_u2_n117, u0_u2_u2_n118, u0_u2_u2_n119, u0_u2_u2_n120, 
       u0_u2_u2_n121, u0_u2_u2_n122, u0_u2_u2_n123, u0_u2_u2_n124, u0_u2_u2_n125, u0_u2_u2_n126, u0_u2_u2_n127, u0_u2_u2_n128, u0_u2_u2_n129, 
       u0_u2_u2_n130, u0_u2_u2_n131, u0_u2_u2_n132, u0_u2_u2_n133, u0_u2_u2_n134, u0_u2_u2_n135, u0_u2_u2_n136, u0_u2_u2_n137, u0_u2_u2_n138, 
       u0_u2_u2_n139, u0_u2_u2_n140, u0_u2_u2_n141, u0_u2_u2_n142, u0_u2_u2_n143, u0_u2_u2_n144, u0_u2_u2_n145, u0_u2_u2_n146, u0_u2_u2_n147, 
       u0_u2_u2_n148, u0_u2_u2_n149, u0_u2_u2_n150, u0_u2_u2_n151, u0_u2_u2_n152, u0_u2_u2_n153, u0_u2_u2_n154, u0_u2_u2_n155, u0_u2_u2_n156, 
       u0_u2_u2_n157, u0_u2_u2_n158, u0_u2_u2_n159, u0_u2_u2_n160, u0_u2_u2_n161, u0_u2_u2_n162, u0_u2_u2_n163, u0_u2_u2_n164, u0_u2_u2_n165, 
       u0_u2_u2_n166, u0_u2_u2_n167, u0_u2_u2_n168, u0_u2_u2_n169, u0_u2_u2_n170, u0_u2_u2_n171, u0_u2_u2_n172, u0_u2_u2_n173, u0_u2_u2_n174, 
       u0_u2_u2_n175, u0_u2_u2_n176, u0_u2_u2_n177, u0_u2_u2_n178, u0_u2_u2_n179, u0_u2_u2_n180, u0_u2_u2_n181, u0_u2_u2_n182, u0_u2_u2_n183, 
       u0_u2_u2_n184, u0_u2_u2_n185, u0_u2_u2_n186, u0_u2_u2_n187, u0_u2_u2_n188, u0_u2_u2_n95, u0_u2_u2_n96, u0_u2_u2_n97, u0_u2_u2_n98, 
       u0_u2_u2_n99, u0_u2_u3_n100, u0_u2_u3_n101, u0_u2_u3_n102, u0_u2_u3_n103, u0_u2_u3_n104, u0_u2_u3_n105, u0_u2_u3_n106, u0_u2_u3_n107, 
       u0_u2_u3_n108, u0_u2_u3_n109, u0_u2_u3_n110, u0_u2_u3_n111, u0_u2_u3_n112, u0_u2_u3_n113, u0_u2_u3_n114, u0_u2_u3_n115, u0_u2_u3_n116, 
       u0_u2_u3_n117, u0_u2_u3_n118, u0_u2_u3_n119, u0_u2_u3_n120, u0_u2_u3_n121, u0_u2_u3_n122, u0_u2_u3_n123, u0_u2_u3_n124, u0_u2_u3_n125, 
       u0_u2_u3_n126, u0_u2_u3_n127, u0_u2_u3_n128, u0_u2_u3_n129, u0_u2_u3_n130, u0_u2_u3_n131, u0_u2_u3_n132, u0_u2_u3_n133, u0_u2_u3_n134, 
       u0_u2_u3_n135, u0_u2_u3_n136, u0_u2_u3_n137, u0_u2_u3_n138, u0_u2_u3_n139, u0_u2_u3_n140, u0_u2_u3_n141, u0_u2_u3_n142, u0_u2_u3_n143, 
       u0_u2_u3_n144, u0_u2_u3_n145, u0_u2_u3_n146, u0_u2_u3_n147, u0_u2_u3_n148, u0_u2_u3_n149, u0_u2_u3_n150, u0_u2_u3_n151, u0_u2_u3_n152, 
       u0_u2_u3_n153, u0_u2_u3_n154, u0_u2_u3_n155, u0_u2_u3_n156, u0_u2_u3_n157, u0_u2_u3_n158, u0_u2_u3_n159, u0_u2_u3_n160, u0_u2_u3_n161, 
       u0_u2_u3_n162, u0_u2_u3_n163, u0_u2_u3_n164, u0_u2_u3_n165, u0_u2_u3_n166, u0_u2_u3_n167, u0_u2_u3_n168, u0_u2_u3_n169, u0_u2_u3_n170, 
       u0_u2_u3_n171, u0_u2_u3_n172, u0_u2_u3_n173, u0_u2_u3_n174, u0_u2_u3_n175, u0_u2_u3_n176, u0_u2_u3_n177, u0_u2_u3_n178, u0_u2_u3_n179, 
       u0_u2_u3_n180, u0_u2_u3_n181, u0_u2_u3_n182, u0_u2_u3_n183, u0_u2_u3_n184, u0_u2_u3_n185, u0_u2_u3_n186, u0_u2_u3_n94, u0_u2_u3_n95, 
       u0_u2_u3_n96, u0_u2_u3_n97, u0_u2_u3_n98, u0_u2_u3_n99, u0_u3_X_1, u0_u3_X_10, u0_u3_X_11, u0_u3_X_12, u0_u3_X_13, 
       u0_u3_X_14, u0_u3_X_15, u0_u3_X_16, u0_u3_X_17, u0_u3_X_18, u0_u3_X_19, u0_u3_X_2, u0_u3_X_20, u0_u3_X_21, 
       u0_u3_X_22, u0_u3_X_23, u0_u3_X_24, u0_u3_X_25, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, u0_u3_X_3, 
       u0_u3_X_30, u0_u3_X_31, u0_u3_X_32, u0_u3_X_33, u0_u3_X_34, u0_u3_X_35, u0_u3_X_36, u0_u3_X_4, u0_u3_X_5, 
       u0_u3_X_6, u0_u3_X_7, u0_u3_X_8, u0_u3_X_9, u0_u3_u0_n100, u0_u3_u0_n101, u0_u3_u0_n102, u0_u3_u0_n103, u0_u3_u0_n104, 
       u0_u3_u0_n105, u0_u3_u0_n106, u0_u3_u0_n107, u0_u3_u0_n108, u0_u3_u0_n109, u0_u3_u0_n110, u0_u3_u0_n111, u0_u3_u0_n112, u0_u3_u0_n113, 
       u0_u3_u0_n114, u0_u3_u0_n115, u0_u3_u0_n116, u0_u3_u0_n117, u0_u3_u0_n118, u0_u3_u0_n119, u0_u3_u0_n120, u0_u3_u0_n121, u0_u3_u0_n122, 
       u0_u3_u0_n123, u0_u3_u0_n124, u0_u3_u0_n125, u0_u3_u0_n126, u0_u3_u0_n127, u0_u3_u0_n128, u0_u3_u0_n129, u0_u3_u0_n130, u0_u3_u0_n131, 
       u0_u3_u0_n132, u0_u3_u0_n133, u0_u3_u0_n134, u0_u3_u0_n135, u0_u3_u0_n136, u0_u3_u0_n137, u0_u3_u0_n138, u0_u3_u0_n139, u0_u3_u0_n140, 
       u0_u3_u0_n141, u0_u3_u0_n142, u0_u3_u0_n143, u0_u3_u0_n144, u0_u3_u0_n145, u0_u3_u0_n146, u0_u3_u0_n147, u0_u3_u0_n148, u0_u3_u0_n149, 
       u0_u3_u0_n150, u0_u3_u0_n151, u0_u3_u0_n152, u0_u3_u0_n153, u0_u3_u0_n154, u0_u3_u0_n155, u0_u3_u0_n156, u0_u3_u0_n157, u0_u3_u0_n158, 
       u0_u3_u0_n159, u0_u3_u0_n160, u0_u3_u0_n161, u0_u3_u0_n162, u0_u3_u0_n163, u0_u3_u0_n164, u0_u3_u0_n165, u0_u3_u0_n166, u0_u3_u0_n167, 
       u0_u3_u0_n168, u0_u3_u0_n169, u0_u3_u0_n170, u0_u3_u0_n171, u0_u3_u0_n172, u0_u3_u0_n173, u0_u3_u0_n174, u0_u3_u0_n175, u0_u3_u0_n176, 
       u0_u3_u0_n88, u0_u3_u0_n89, u0_u3_u0_n90, u0_u3_u0_n91, u0_u3_u0_n92, u0_u3_u0_n93, u0_u3_u0_n94, u0_u3_u0_n95, u0_u3_u0_n96, 
       u0_u3_u0_n97, u0_u3_u0_n98, u0_u3_u0_n99, u0_u3_u1_n100, u0_u3_u1_n101, u0_u3_u1_n102, u0_u3_u1_n103, u0_u3_u1_n104, u0_u3_u1_n105, 
       u0_u3_u1_n106, u0_u3_u1_n107, u0_u3_u1_n108, u0_u3_u1_n109, u0_u3_u1_n110, u0_u3_u1_n111, u0_u3_u1_n112, u0_u3_u1_n113, u0_u3_u1_n114, 
       u0_u3_u1_n115, u0_u3_u1_n116, u0_u3_u1_n117, u0_u3_u1_n118, u0_u3_u1_n119, u0_u3_u1_n120, u0_u3_u1_n121, u0_u3_u1_n122, u0_u3_u1_n123, 
       u0_u3_u1_n124, u0_u3_u1_n125, u0_u3_u1_n126, u0_u3_u1_n127, u0_u3_u1_n128, u0_u3_u1_n129, u0_u3_u1_n130, u0_u3_u1_n131, u0_u3_u1_n132, 
       u0_u3_u1_n133, u0_u3_u1_n134, u0_u3_u1_n135, u0_u3_u1_n136, u0_u3_u1_n137, u0_u3_u1_n138, u0_u3_u1_n139, u0_u3_u1_n140, u0_u3_u1_n141, 
       u0_u3_u1_n142, u0_u3_u1_n143, u0_u3_u1_n144, u0_u3_u1_n145, u0_u3_u1_n146, u0_u3_u1_n147, u0_u3_u1_n148, u0_u3_u1_n149, u0_u3_u1_n150, 
       u0_u3_u1_n151, u0_u3_u1_n152, u0_u3_u1_n153, u0_u3_u1_n154, u0_u3_u1_n155, u0_u3_u1_n156, u0_u3_u1_n157, u0_u3_u1_n158, u0_u3_u1_n159, 
       u0_u3_u1_n160, u0_u3_u1_n161, u0_u3_u1_n162, u0_u3_u1_n163, u0_u3_u1_n164, u0_u3_u1_n165, u0_u3_u1_n166, u0_u3_u1_n167, u0_u3_u1_n168, 
       u0_u3_u1_n169, u0_u3_u1_n170, u0_u3_u1_n171, u0_u3_u1_n172, u0_u3_u1_n173, u0_u3_u1_n174, u0_u3_u1_n175, u0_u3_u1_n176, u0_u3_u1_n177, 
       u0_u3_u1_n178, u0_u3_u1_n179, u0_u3_u1_n180, u0_u3_u1_n181, u0_u3_u1_n182, u0_u3_u1_n183, u0_u3_u1_n184, u0_u3_u1_n185, u0_u3_u1_n186, 
       u0_u3_u1_n187, u0_u3_u1_n188, u0_u3_u1_n95, u0_u3_u1_n96, u0_u3_u1_n97, u0_u3_u1_n98, u0_u3_u1_n99, u0_u3_u2_n100, u0_u3_u2_n101, 
       u0_u3_u2_n102, u0_u3_u2_n103, u0_u3_u2_n104, u0_u3_u2_n105, u0_u3_u2_n106, u0_u3_u2_n107, u0_u3_u2_n108, u0_u3_u2_n109, u0_u3_u2_n110, 
       u0_u3_u2_n111, u0_u3_u2_n112, u0_u3_u2_n113, u0_u3_u2_n114, u0_u3_u2_n115, u0_u3_u2_n116, u0_u3_u2_n117, u0_u3_u2_n118, u0_u3_u2_n119, 
       u0_u3_u2_n120, u0_u3_u2_n121, u0_u3_u2_n122, u0_u3_u2_n123, u0_u3_u2_n124, u0_u3_u2_n125, u0_u3_u2_n126, u0_u3_u2_n127, u0_u3_u2_n128, 
       u0_u3_u2_n129, u0_u3_u2_n130, u0_u3_u2_n131, u0_u3_u2_n132, u0_u3_u2_n133, u0_u3_u2_n134, u0_u3_u2_n135, u0_u3_u2_n136, u0_u3_u2_n137, 
       u0_u3_u2_n138, u0_u3_u2_n139, u0_u3_u2_n140, u0_u3_u2_n141, u0_u3_u2_n142, u0_u3_u2_n143, u0_u3_u2_n144, u0_u3_u2_n145, u0_u3_u2_n146, 
       u0_u3_u2_n147, u0_u3_u2_n148, u0_u3_u2_n149, u0_u3_u2_n150, u0_u3_u2_n151, u0_u3_u2_n152, u0_u3_u2_n153, u0_u3_u2_n154, u0_u3_u2_n155, 
       u0_u3_u2_n156, u0_u3_u2_n157, u0_u3_u2_n158, u0_u3_u2_n159, u0_u3_u2_n160, u0_u3_u2_n161, u0_u3_u2_n162, u0_u3_u2_n163, u0_u3_u2_n164, 
       u0_u3_u2_n165, u0_u3_u2_n166, u0_u3_u2_n167, u0_u3_u2_n168, u0_u3_u2_n169, u0_u3_u2_n170, u0_u3_u2_n171, u0_u3_u2_n172, u0_u3_u2_n173, 
       u0_u3_u2_n174, u0_u3_u2_n175, u0_u3_u2_n176, u0_u3_u2_n177, u0_u3_u2_n178, u0_u3_u2_n179, u0_u3_u2_n180, u0_u3_u2_n181, u0_u3_u2_n182, 
       u0_u3_u2_n183, u0_u3_u2_n184, u0_u3_u2_n185, u0_u3_u2_n186, u0_u3_u2_n187, u0_u3_u2_n188, u0_u3_u2_n95, u0_u3_u2_n96, u0_u3_u2_n97, 
       u0_u3_u2_n98, u0_u3_u2_n99, u0_u3_u3_n100, u0_u3_u3_n101, u0_u3_u3_n102, u0_u3_u3_n103, u0_u3_u3_n104, u0_u3_u3_n105, u0_u3_u3_n106, 
       u0_u3_u3_n107, u0_u3_u3_n108, u0_u3_u3_n109, u0_u3_u3_n110, u0_u3_u3_n111, u0_u3_u3_n112, u0_u3_u3_n113, u0_u3_u3_n114, u0_u3_u3_n115, 
       u0_u3_u3_n116, u0_u3_u3_n117, u0_u3_u3_n118, u0_u3_u3_n119, u0_u3_u3_n120, u0_u3_u3_n121, u0_u3_u3_n122, u0_u3_u3_n123, u0_u3_u3_n124, 
       u0_u3_u3_n125, u0_u3_u3_n126, u0_u3_u3_n127, u0_u3_u3_n128, u0_u3_u3_n129, u0_u3_u3_n130, u0_u3_u3_n131, u0_u3_u3_n132, u0_u3_u3_n133, 
       u0_u3_u3_n134, u0_u3_u3_n135, u0_u3_u3_n136, u0_u3_u3_n137, u0_u3_u3_n138, u0_u3_u3_n139, u0_u3_u3_n140, u0_u3_u3_n141, u0_u3_u3_n142, 
       u0_u3_u3_n143, u0_u3_u3_n144, u0_u3_u3_n145, u0_u3_u3_n146, u0_u3_u3_n147, u0_u3_u3_n148, u0_u3_u3_n149, u0_u3_u3_n150, u0_u3_u3_n151, 
       u0_u3_u3_n152, u0_u3_u3_n153, u0_u3_u3_n154, u0_u3_u3_n155, u0_u3_u3_n156, u0_u3_u3_n157, u0_u3_u3_n158, u0_u3_u3_n159, u0_u3_u3_n160, 
       u0_u3_u3_n161, u0_u3_u3_n162, u0_u3_u3_n163, u0_u3_u3_n164, u0_u3_u3_n165, u0_u3_u3_n166, u0_u3_u3_n167, u0_u3_u3_n168, u0_u3_u3_n169, 
       u0_u3_u3_n170, u0_u3_u3_n171, u0_u3_u3_n172, u0_u3_u3_n173, u0_u3_u3_n174, u0_u3_u3_n175, u0_u3_u3_n176, u0_u3_u3_n177, u0_u3_u3_n178, 
       u0_u3_u3_n179, u0_u3_u3_n180, u0_u3_u3_n181, u0_u3_u3_n182, u0_u3_u3_n183, u0_u3_u3_n184, u0_u3_u3_n185, u0_u3_u3_n186, u0_u3_u3_n94, 
       u0_u3_u3_n95, u0_u3_u3_n96, u0_u3_u3_n97, u0_u3_u3_n98, u0_u3_u3_n99, u0_u3_u4_n100, u0_u3_u4_n101, u0_u3_u4_n102, u0_u3_u4_n103, 
       u0_u3_u4_n104, u0_u3_u4_n105, u0_u3_u4_n106, u0_u3_u4_n107, u0_u3_u4_n108, u0_u3_u4_n109, u0_u3_u4_n110, u0_u3_u4_n111, u0_u3_u4_n112, 
       u0_u3_u4_n113, u0_u3_u4_n114, u0_u3_u4_n115, u0_u3_u4_n116, u0_u3_u4_n117, u0_u3_u4_n118, u0_u3_u4_n119, u0_u3_u4_n120, u0_u3_u4_n121, 
       u0_u3_u4_n122, u0_u3_u4_n123, u0_u3_u4_n124, u0_u3_u4_n125, u0_u3_u4_n126, u0_u3_u4_n127, u0_u3_u4_n128, u0_u3_u4_n129, u0_u3_u4_n130, 
       u0_u3_u4_n131, u0_u3_u4_n132, u0_u3_u4_n133, u0_u3_u4_n134, u0_u3_u4_n135, u0_u3_u4_n136, u0_u3_u4_n137, u0_u3_u4_n138, u0_u3_u4_n139, 
       u0_u3_u4_n140, u0_u3_u4_n141, u0_u3_u4_n142, u0_u3_u4_n143, u0_u3_u4_n144, u0_u3_u4_n145, u0_u3_u4_n146, u0_u3_u4_n147, u0_u3_u4_n148, 
       u0_u3_u4_n149, u0_u3_u4_n150, u0_u3_u4_n151, u0_u3_u4_n152, u0_u3_u4_n153, u0_u3_u4_n154, u0_u3_u4_n155, u0_u3_u4_n156, u0_u3_u4_n157, 
       u0_u3_u4_n158, u0_u3_u4_n159, u0_u3_u4_n160, u0_u3_u4_n161, u0_u3_u4_n162, u0_u3_u4_n163, u0_u3_u4_n164, u0_u3_u4_n165, u0_u3_u4_n166, 
       u0_u3_u4_n167, u0_u3_u4_n168, u0_u3_u4_n169, u0_u3_u4_n170, u0_u3_u4_n171, u0_u3_u4_n172, u0_u3_u4_n173, u0_u3_u4_n174, u0_u3_u4_n175, 
       u0_u3_u4_n176, u0_u3_u4_n177, u0_u3_u4_n178, u0_u3_u4_n179, u0_u3_u4_n180, u0_u3_u4_n181, u0_u3_u4_n182, u0_u3_u4_n183, u0_u3_u4_n184, 
       u0_u3_u4_n185, u0_u3_u4_n186, u0_u3_u4_n94, u0_u3_u4_n95, u0_u3_u4_n96, u0_u3_u4_n97, u0_u3_u4_n98, u0_u3_u4_n99, u0_u3_u5_n100, 
       u0_u3_u5_n101, u0_u3_u5_n102, u0_u3_u5_n103, u0_u3_u5_n104, u0_u3_u5_n105, u0_u3_u5_n106, u0_u3_u5_n107, u0_u3_u5_n108, u0_u3_u5_n109, 
       u0_u3_u5_n110, u0_u3_u5_n111, u0_u3_u5_n112, u0_u3_u5_n113, u0_u3_u5_n114, u0_u3_u5_n115, u0_u3_u5_n116, u0_u3_u5_n117, u0_u3_u5_n118, 
       u0_u3_u5_n119, u0_u3_u5_n120, u0_u3_u5_n121, u0_u3_u5_n122, u0_u3_u5_n123, u0_u3_u5_n124, u0_u3_u5_n125, u0_u3_u5_n126, u0_u3_u5_n127, 
       u0_u3_u5_n128, u0_u3_u5_n129, u0_u3_u5_n130, u0_u3_u5_n131, u0_u3_u5_n132, u0_u3_u5_n133, u0_u3_u5_n134, u0_u3_u5_n135, u0_u3_u5_n136, 
       u0_u3_u5_n137, u0_u3_u5_n138, u0_u3_u5_n139, u0_u3_u5_n140, u0_u3_u5_n141, u0_u3_u5_n142, u0_u3_u5_n143, u0_u3_u5_n144, u0_u3_u5_n145, 
       u0_u3_u5_n146, u0_u3_u5_n147, u0_u3_u5_n148, u0_u3_u5_n149, u0_u3_u5_n150, u0_u3_u5_n151, u0_u3_u5_n152, u0_u3_u5_n153, u0_u3_u5_n154, 
       u0_u3_u5_n155, u0_u3_u5_n156, u0_u3_u5_n157, u0_u3_u5_n158, u0_u3_u5_n159, u0_u3_u5_n160, u0_u3_u5_n161, u0_u3_u5_n162, u0_u3_u5_n163, 
       u0_u3_u5_n164, u0_u3_u5_n165, u0_u3_u5_n166, u0_u3_u5_n167, u0_u3_u5_n168, u0_u3_u5_n169, u0_u3_u5_n170, u0_u3_u5_n171, u0_u3_u5_n172, 
       u0_u3_u5_n173, u0_u3_u5_n174, u0_u3_u5_n175, u0_u3_u5_n176, u0_u3_u5_n177, u0_u3_u5_n178, u0_u3_u5_n179, u0_u3_u5_n180, u0_u3_u5_n181, 
       u0_u3_u5_n182, u0_u3_u5_n183, u0_u3_u5_n184, u0_u3_u5_n185, u0_u3_u5_n186, u0_u3_u5_n187, u0_u3_u5_n188, u0_u3_u5_n189, u0_u3_u5_n190, 
       u0_u3_u5_n191, u0_u3_u5_n192, u0_u3_u5_n193, u0_u3_u5_n194, u0_u3_u5_n195, u0_u3_u5_n196, u0_u3_u5_n99, u0_u5_X_19, u0_u5_X_20, 
       u0_u5_X_21, u0_u5_X_22, u0_u5_X_23, u0_u5_X_24, u0_u5_X_25, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, 
       u0_u5_X_30, u0_u5_X_31, u0_u5_X_32, u0_u5_X_33, u0_u5_X_34, u0_u5_X_35, u0_u5_X_36, u0_u5_X_37, u0_u5_X_38, 
       u0_u5_X_39, u0_u5_X_40, u0_u5_X_41, u0_u5_X_42, u0_u5_u3_n100, u0_u5_u3_n101, u0_u5_u3_n102, u0_u5_u3_n103, u0_u5_u3_n104, 
       u0_u5_u3_n105, u0_u5_u3_n106, u0_u5_u3_n107, u0_u5_u3_n108, u0_u5_u3_n109, u0_u5_u3_n110, u0_u5_u3_n111, u0_u5_u3_n112, u0_u5_u3_n113, 
       u0_u5_u3_n114, u0_u5_u3_n115, u0_u5_u3_n116, u0_u5_u3_n117, u0_u5_u3_n118, u0_u5_u3_n119, u0_u5_u3_n120, u0_u5_u3_n121, u0_u5_u3_n122, 
       u0_u5_u3_n123, u0_u5_u3_n124, u0_u5_u3_n125, u0_u5_u3_n126, u0_u5_u3_n127, u0_u5_u3_n128, u0_u5_u3_n129, u0_u5_u3_n130, u0_u5_u3_n131, 
       u0_u5_u3_n132, u0_u5_u3_n133, u0_u5_u3_n134, u0_u5_u3_n135, u0_u5_u3_n136, u0_u5_u3_n137, u0_u5_u3_n138, u0_u5_u3_n139, u0_u5_u3_n140, 
       u0_u5_u3_n141, u0_u5_u3_n142, u0_u5_u3_n143, u0_u5_u3_n144, u0_u5_u3_n145, u0_u5_u3_n146, u0_u5_u3_n147, u0_u5_u3_n148, u0_u5_u3_n149, 
       u0_u5_u3_n150, u0_u5_u3_n151, u0_u5_u3_n152, u0_u5_u3_n153, u0_u5_u3_n154, u0_u5_u3_n155, u0_u5_u3_n156, u0_u5_u3_n157, u0_u5_u3_n158, 
       u0_u5_u3_n159, u0_u5_u3_n160, u0_u5_u3_n161, u0_u5_u3_n162, u0_u5_u3_n163, u0_u5_u3_n164, u0_u5_u3_n165, u0_u5_u3_n166, u0_u5_u3_n167, 
       u0_u5_u3_n168, u0_u5_u3_n169, u0_u5_u3_n170, u0_u5_u3_n171, u0_u5_u3_n172, u0_u5_u3_n173, u0_u5_u3_n174, u0_u5_u3_n175, u0_u5_u3_n176, 
       u0_u5_u3_n177, u0_u5_u3_n178, u0_u5_u3_n179, u0_u5_u3_n180, u0_u5_u3_n181, u0_u5_u3_n182, u0_u5_u3_n183, u0_u5_u3_n184, u0_u5_u3_n185, 
       u0_u5_u3_n186, u0_u5_u3_n94, u0_u5_u3_n95, u0_u5_u3_n96, u0_u5_u3_n97, u0_u5_u3_n98, u0_u5_u3_n99, u0_u5_u4_n100, u0_u5_u4_n101, 
       u0_u5_u4_n102, u0_u5_u4_n103, u0_u5_u4_n104, u0_u5_u4_n105, u0_u5_u4_n106, u0_u5_u4_n107, u0_u5_u4_n108, u0_u5_u4_n109, u0_u5_u4_n110, 
       u0_u5_u4_n111, u0_u5_u4_n112, u0_u5_u4_n113, u0_u5_u4_n114, u0_u5_u4_n115, u0_u5_u4_n116, u0_u5_u4_n117, u0_u5_u4_n118, u0_u5_u4_n119, 
       u0_u5_u4_n120, u0_u5_u4_n121, u0_u5_u4_n122, u0_u5_u4_n123, u0_u5_u4_n124, u0_u5_u4_n125, u0_u5_u4_n126, u0_u5_u4_n127, u0_u5_u4_n128, 
       u0_u5_u4_n129, u0_u5_u4_n130, u0_u5_u4_n131, u0_u5_u4_n132, u0_u5_u4_n133, u0_u5_u4_n134, u0_u5_u4_n135, u0_u5_u4_n136, u0_u5_u4_n137, 
       u0_u5_u4_n138, u0_u5_u4_n139, u0_u5_u4_n140, u0_u5_u4_n141, u0_u5_u4_n142, u0_u5_u4_n143, u0_u5_u4_n144, u0_u5_u4_n145, u0_u5_u4_n146, 
       u0_u5_u4_n147, u0_u5_u4_n148, u0_u5_u4_n149, u0_u5_u4_n150, u0_u5_u4_n151, u0_u5_u4_n152, u0_u5_u4_n153, u0_u5_u4_n154, u0_u5_u4_n155, 
       u0_u5_u4_n156, u0_u5_u4_n157, u0_u5_u4_n158, u0_u5_u4_n159, u0_u5_u4_n160, u0_u5_u4_n161, u0_u5_u4_n162, u0_u5_u4_n163, u0_u5_u4_n164, 
       u0_u5_u4_n165, u0_u5_u4_n166, u0_u5_u4_n167, u0_u5_u4_n168, u0_u5_u4_n169, u0_u5_u4_n170, u0_u5_u4_n171, u0_u5_u4_n172, u0_u5_u4_n173, 
       u0_u5_u4_n174, u0_u5_u4_n175, u0_u5_u4_n176, u0_u5_u4_n177, u0_u5_u4_n178, u0_u5_u4_n179, u0_u5_u4_n180, u0_u5_u4_n181, u0_u5_u4_n182, 
       u0_u5_u4_n183, u0_u5_u4_n184, u0_u5_u4_n185, u0_u5_u4_n186, u0_u5_u4_n94, u0_u5_u4_n95, u0_u5_u4_n96, u0_u5_u4_n97, u0_u5_u4_n98, 
       u0_u5_u4_n99, u0_u5_u5_n100, u0_u5_u5_n101, u0_u5_u5_n102, u0_u5_u5_n103, u0_u5_u5_n104, u0_u5_u5_n105, u0_u5_u5_n106, u0_u5_u5_n107, 
       u0_u5_u5_n108, u0_u5_u5_n109, u0_u5_u5_n110, u0_u5_u5_n111, u0_u5_u5_n112, u0_u5_u5_n113, u0_u5_u5_n114, u0_u5_u5_n115, u0_u5_u5_n116, 
       u0_u5_u5_n117, u0_u5_u5_n118, u0_u5_u5_n119, u0_u5_u5_n120, u0_u5_u5_n121, u0_u5_u5_n122, u0_u5_u5_n123, u0_u5_u5_n124, u0_u5_u5_n125, 
       u0_u5_u5_n126, u0_u5_u5_n127, u0_u5_u5_n128, u0_u5_u5_n129, u0_u5_u5_n130, u0_u5_u5_n131, u0_u5_u5_n132, u0_u5_u5_n133, u0_u5_u5_n134, 
       u0_u5_u5_n135, u0_u5_u5_n136, u0_u5_u5_n137, u0_u5_u5_n138, u0_u5_u5_n139, u0_u5_u5_n140, u0_u5_u5_n141, u0_u5_u5_n142, u0_u5_u5_n143, 
       u0_u5_u5_n144, u0_u5_u5_n145, u0_u5_u5_n146, u0_u5_u5_n147, u0_u5_u5_n148, u0_u5_u5_n149, u0_u5_u5_n150, u0_u5_u5_n151, u0_u5_u5_n152, 
       u0_u5_u5_n153, u0_u5_u5_n154, u0_u5_u5_n155, u0_u5_u5_n156, u0_u5_u5_n157, u0_u5_u5_n158, u0_u5_u5_n159, u0_u5_u5_n160, u0_u5_u5_n161, 
       u0_u5_u5_n162, u0_u5_u5_n163, u0_u5_u5_n164, u0_u5_u5_n165, u0_u5_u5_n166, u0_u5_u5_n167, u0_u5_u5_n168, u0_u5_u5_n169, u0_u5_u5_n170, 
       u0_u5_u5_n171, u0_u5_u5_n172, u0_u5_u5_n173, u0_u5_u5_n174, u0_u5_u5_n175, u0_u5_u5_n176, u0_u5_u5_n177, u0_u5_u5_n178, u0_u5_u5_n179, 
       u0_u5_u5_n180, u0_u5_u5_n181, u0_u5_u5_n182, u0_u5_u5_n183, u0_u5_u5_n184, u0_u5_u5_n185, u0_u5_u5_n186, u0_u5_u5_n187, u0_u5_u5_n188, 
       u0_u5_u5_n189, u0_u5_u5_n190, u0_u5_u5_n191, u0_u5_u5_n192, u0_u5_u5_n193, u0_u5_u5_n194, u0_u5_u5_n195, u0_u5_u5_n196, u0_u5_u5_n99, 
       u0_u5_u6_n100, u0_u5_u6_n101, u0_u5_u6_n102, u0_u5_u6_n103, u0_u5_u6_n104, u0_u5_u6_n105, u0_u5_u6_n106, u0_u5_u6_n107, u0_u5_u6_n108, 
       u0_u5_u6_n109, u0_u5_u6_n110, u0_u5_u6_n111, u0_u5_u6_n112, u0_u5_u6_n113, u0_u5_u6_n114, u0_u5_u6_n115, u0_u5_u6_n116, u0_u5_u6_n117, 
       u0_u5_u6_n118, u0_u5_u6_n119, u0_u5_u6_n120, u0_u5_u6_n121, u0_u5_u6_n122, u0_u5_u6_n123, u0_u5_u6_n124, u0_u5_u6_n125, u0_u5_u6_n126, 
       u0_u5_u6_n127, u0_u5_u6_n128, u0_u5_u6_n129, u0_u5_u6_n130, u0_u5_u6_n131, u0_u5_u6_n132, u0_u5_u6_n133, u0_u5_u6_n134, u0_u5_u6_n135, 
       u0_u5_u6_n136, u0_u5_u6_n137, u0_u5_u6_n138, u0_u5_u6_n139, u0_u5_u6_n140, u0_u5_u6_n141, u0_u5_u6_n142, u0_u5_u6_n143, u0_u5_u6_n144, 
       u0_u5_u6_n145, u0_u5_u6_n146, u0_u5_u6_n147, u0_u5_u6_n148, u0_u5_u6_n149, u0_u5_u6_n150, u0_u5_u6_n151, u0_u5_u6_n152, u0_u5_u6_n153, 
       u0_u5_u6_n154, u0_u5_u6_n155, u0_u5_u6_n156, u0_u5_u6_n157, u0_u5_u6_n158, u0_u5_u6_n159, u0_u5_u6_n160, u0_u5_u6_n161, u0_u5_u6_n162, 
       u0_u5_u6_n163, u0_u5_u6_n164, u0_u5_u6_n165, u0_u5_u6_n166, u0_u5_u6_n167, u0_u5_u6_n168, u0_u5_u6_n169, u0_u5_u6_n170, u0_u5_u6_n171, 
       u0_u5_u6_n172, u0_u5_u6_n173, u0_u5_u6_n174, u0_u5_u6_n88, u0_u5_u6_n89, u0_u5_u6_n90, u0_u5_u6_n91, u0_u5_u6_n92, u0_u5_u6_n93, 
       u0_u5_u6_n94, u0_u5_u6_n95, u0_u5_u6_n96, u0_u5_u6_n97, u0_u5_u6_n98, u0_u5_u6_n99, u0_u6_X_1, u0_u6_X_10, u0_u6_X_11, 
       u0_u6_X_12, u0_u6_X_13, u0_u6_X_14, u0_u6_X_15, u0_u6_X_16, u0_u6_X_17, u0_u6_X_18, u0_u6_X_19, u0_u6_X_2, 
       u0_u6_X_20, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_3, u0_u6_X_4, u0_u6_X_43, u0_u6_X_44, 
       u0_u6_X_45, u0_u6_X_46, u0_u6_X_47, u0_u6_X_48, u0_u6_X_5, u0_u6_X_6, u0_u6_X_7, u0_u6_X_8, u0_u6_X_9, 
       u0_u6_u0_n100, u0_u6_u0_n101, u0_u6_u0_n102, u0_u6_u0_n103, u0_u6_u0_n104, u0_u6_u0_n105, u0_u6_u0_n106, u0_u6_u0_n107, u0_u6_u0_n108, 
       u0_u6_u0_n109, u0_u6_u0_n110, u0_u6_u0_n111, u0_u6_u0_n112, u0_u6_u0_n113, u0_u6_u0_n114, u0_u6_u0_n115, u0_u6_u0_n116, u0_u6_u0_n117, 
       u0_u6_u0_n118, u0_u6_u0_n119, u0_u6_u0_n120, u0_u6_u0_n121, u0_u6_u0_n122, u0_u6_u0_n123, u0_u6_u0_n124, u0_u6_u0_n125, u0_u6_u0_n126, 
       u0_u6_u0_n127, u0_u6_u0_n128, u0_u6_u0_n129, u0_u6_u0_n130, u0_u6_u0_n131, u0_u6_u0_n132, u0_u6_u0_n133, u0_u6_u0_n134, u0_u6_u0_n135, 
       u0_u6_u0_n136, u0_u6_u0_n137, u0_u6_u0_n138, u0_u6_u0_n139, u0_u6_u0_n140, u0_u6_u0_n141, u0_u6_u0_n142, u0_u6_u0_n143, u0_u6_u0_n144, 
       u0_u6_u0_n145, u0_u6_u0_n146, u0_u6_u0_n147, u0_u6_u0_n148, u0_u6_u0_n149, u0_u6_u0_n150, u0_u6_u0_n151, u0_u6_u0_n152, u0_u6_u0_n153, 
       u0_u6_u0_n154, u0_u6_u0_n155, u0_u6_u0_n156, u0_u6_u0_n157, u0_u6_u0_n158, u0_u6_u0_n159, u0_u6_u0_n160, u0_u6_u0_n161, u0_u6_u0_n162, 
       u0_u6_u0_n163, u0_u6_u0_n164, u0_u6_u0_n165, u0_u6_u0_n166, u0_u6_u0_n167, u0_u6_u0_n168, u0_u6_u0_n169, u0_u6_u0_n170, u0_u6_u0_n171, 
       u0_u6_u0_n172, u0_u6_u0_n173, u0_u6_u0_n174, u0_u6_u0_n88, u0_u6_u0_n89, u0_u6_u0_n90, u0_u6_u0_n91, u0_u6_u0_n92, u0_u6_u0_n93, 
       u0_u6_u0_n94, u0_u6_u0_n95, u0_u6_u0_n96, u0_u6_u0_n97, u0_u6_u0_n98, u0_u6_u0_n99, u0_u6_u1_n100, u0_u6_u1_n101, u0_u6_u1_n102, 
       u0_u6_u1_n103, u0_u6_u1_n104, u0_u6_u1_n105, u0_u6_u1_n106, u0_u6_u1_n107, u0_u6_u1_n108, u0_u6_u1_n109, u0_u6_u1_n110, u0_u6_u1_n111, 
       u0_u6_u1_n112, u0_u6_u1_n113, u0_u6_u1_n114, u0_u6_u1_n115, u0_u6_u1_n116, u0_u6_u1_n117, u0_u6_u1_n118, u0_u6_u1_n119, u0_u6_u1_n120, 
       u0_u6_u1_n121, u0_u6_u1_n122, u0_u6_u1_n123, u0_u6_u1_n124, u0_u6_u1_n125, u0_u6_u1_n126, u0_u6_u1_n127, u0_u6_u1_n128, u0_u6_u1_n129, 
       u0_u6_u1_n130, u0_u6_u1_n131, u0_u6_u1_n132, u0_u6_u1_n133, u0_u6_u1_n134, u0_u6_u1_n135, u0_u6_u1_n136, u0_u6_u1_n137, u0_u6_u1_n138, 
       u0_u6_u1_n139, u0_u6_u1_n140, u0_u6_u1_n141, u0_u6_u1_n142, u0_u6_u1_n143, u0_u6_u1_n144, u0_u6_u1_n145, u0_u6_u1_n146, u0_u6_u1_n147, 
       u0_u6_u1_n148, u0_u6_u1_n149, u0_u6_u1_n150, u0_u6_u1_n151, u0_u6_u1_n152, u0_u6_u1_n153, u0_u6_u1_n154, u0_u6_u1_n155, u0_u6_u1_n156, 
       u0_u6_u1_n157, u0_u6_u1_n158, u0_u6_u1_n159, u0_u6_u1_n160, u0_u6_u1_n161, u0_u6_u1_n162, u0_u6_u1_n163, u0_u6_u1_n164, u0_u6_u1_n165, 
       u0_u6_u1_n166, u0_u6_u1_n167, u0_u6_u1_n168, u0_u6_u1_n169, u0_u6_u1_n170, u0_u6_u1_n171, u0_u6_u1_n172, u0_u6_u1_n173, u0_u6_u1_n174, 
       u0_u6_u1_n175, u0_u6_u1_n176, u0_u6_u1_n177, u0_u6_u1_n178, u0_u6_u1_n179, u0_u6_u1_n180, u0_u6_u1_n181, u0_u6_u1_n182, u0_u6_u1_n183, 
       u0_u6_u1_n184, u0_u6_u1_n185, u0_u6_u1_n186, u0_u6_u1_n187, u0_u6_u1_n188, u0_u6_u1_n95, u0_u6_u1_n96, u0_u6_u1_n97, u0_u6_u1_n98, 
       u0_u6_u1_n99, u0_u6_u2_n100, u0_u6_u2_n101, u0_u6_u2_n102, u0_u6_u2_n103, u0_u6_u2_n104, u0_u6_u2_n105, u0_u6_u2_n106, u0_u6_u2_n107, 
       u0_u6_u2_n108, u0_u6_u2_n109, u0_u6_u2_n110, u0_u6_u2_n111, u0_u6_u2_n112, u0_u6_u2_n113, u0_u6_u2_n114, u0_u6_u2_n115, u0_u6_u2_n116, 
       u0_u6_u2_n117, u0_u6_u2_n118, u0_u6_u2_n119, u0_u6_u2_n120, u0_u6_u2_n121, u0_u6_u2_n122, u0_u6_u2_n123, u0_u6_u2_n124, u0_u6_u2_n125, 
       u0_u6_u2_n126, u0_u6_u2_n127, u0_u6_u2_n128, u0_u6_u2_n129, u0_u6_u2_n130, u0_u6_u2_n131, u0_u6_u2_n132, u0_u6_u2_n133, u0_u6_u2_n134, 
       u0_u6_u2_n135, u0_u6_u2_n136, u0_u6_u2_n137, u0_u6_u2_n138, u0_u6_u2_n139, u0_u6_u2_n140, u0_u6_u2_n141, u0_u6_u2_n142, u0_u6_u2_n143, 
       u0_u6_u2_n144, u0_u6_u2_n145, u0_u6_u2_n146, u0_u6_u2_n147, u0_u6_u2_n148, u0_u6_u2_n149, u0_u6_u2_n150, u0_u6_u2_n151, u0_u6_u2_n152, 
       u0_u6_u2_n153, u0_u6_u2_n154, u0_u6_u2_n155, u0_u6_u2_n156, u0_u6_u2_n157, u0_u6_u2_n158, u0_u6_u2_n159, u0_u6_u2_n160, u0_u6_u2_n161, 
       u0_u6_u2_n162, u0_u6_u2_n163, u0_u6_u2_n164, u0_u6_u2_n165, u0_u6_u2_n166, u0_u6_u2_n167, u0_u6_u2_n168, u0_u6_u2_n169, u0_u6_u2_n170, 
       u0_u6_u2_n171, u0_u6_u2_n172, u0_u6_u2_n173, u0_u6_u2_n174, u0_u6_u2_n175, u0_u6_u2_n176, u0_u6_u2_n177, u0_u6_u2_n178, u0_u6_u2_n179, 
       u0_u6_u2_n180, u0_u6_u2_n181, u0_u6_u2_n182, u0_u6_u2_n183, u0_u6_u2_n184, u0_u6_u2_n185, u0_u6_u2_n186, u0_u6_u2_n187, u0_u6_u2_n188, 
       u0_u6_u2_n95, u0_u6_u2_n96, u0_u6_u2_n97, u0_u6_u2_n98, u0_u6_u2_n99, u0_u6_u3_n100, u0_u6_u3_n101, u0_u6_u3_n102, u0_u6_u3_n103, 
       u0_u6_u3_n104, u0_u6_u3_n105, u0_u6_u3_n106, u0_u6_u3_n107, u0_u6_u3_n108, u0_u6_u3_n109, u0_u6_u3_n110, u0_u6_u3_n111, u0_u6_u3_n112, 
       u0_u6_u3_n113, u0_u6_u3_n114, u0_u6_u3_n115, u0_u6_u3_n116, u0_u6_u3_n117, u0_u6_u3_n118, u0_u6_u3_n119, u0_u6_u3_n120, u0_u6_u3_n121, 
       u0_u6_u3_n122, u0_u6_u3_n123, u0_u6_u3_n124, u0_u6_u3_n125, u0_u6_u3_n126, u0_u6_u3_n127, u0_u6_u3_n128, u0_u6_u3_n129, u0_u6_u3_n130, 
       u0_u6_u3_n131, u0_u6_u3_n132, u0_u6_u3_n133, u0_u6_u3_n134, u0_u6_u3_n135, u0_u6_u3_n136, u0_u6_u3_n137, u0_u6_u3_n138, u0_u6_u3_n139, 
       u0_u6_u3_n140, u0_u6_u3_n141, u0_u6_u3_n142, u0_u6_u3_n143, u0_u6_u3_n144, u0_u6_u3_n145, u0_u6_u3_n146, u0_u6_u3_n147, u0_u6_u3_n148, 
       u0_u6_u3_n149, u0_u6_u3_n150, u0_u6_u3_n151, u0_u6_u3_n152, u0_u6_u3_n153, u0_u6_u3_n154, u0_u6_u3_n155, u0_u6_u3_n156, u0_u6_u3_n157, 
       u0_u6_u3_n158, u0_u6_u3_n159, u0_u6_u3_n160, u0_u6_u3_n161, u0_u6_u3_n162, u0_u6_u3_n163, u0_u6_u3_n164, u0_u6_u3_n165, u0_u6_u3_n166, 
       u0_u6_u3_n167, u0_u6_u3_n168, u0_u6_u3_n169, u0_u6_u3_n170, u0_u6_u3_n171, u0_u6_u3_n172, u0_u6_u3_n173, u0_u6_u3_n174, u0_u6_u3_n175, 
       u0_u6_u3_n176, u0_u6_u3_n177, u0_u6_u3_n178, u0_u6_u3_n179, u0_u6_u3_n180, u0_u6_u3_n181, u0_u6_u3_n182, u0_u6_u3_n183, u0_u6_u3_n184, 
       u0_u6_u3_n185, u0_u6_u3_n186, u0_u6_u3_n94, u0_u6_u3_n95, u0_u6_u3_n96, u0_u6_u3_n97, u0_u6_u3_n98, u0_u6_u3_n99, u0_u6_u7_n100, 
       u0_u6_u7_n101, u0_u6_u7_n102, u0_u6_u7_n103, u0_u6_u7_n104, u0_u6_u7_n105, u0_u6_u7_n106, u0_u6_u7_n107, u0_u6_u7_n108, u0_u6_u7_n109, 
       u0_u6_u7_n110, u0_u6_u7_n111, u0_u6_u7_n112, u0_u6_u7_n113, u0_u6_u7_n114, u0_u6_u7_n115, u0_u6_u7_n116, u0_u6_u7_n117, u0_u6_u7_n118, 
       u0_u6_u7_n119, u0_u6_u7_n120, u0_u6_u7_n121, u0_u6_u7_n122, u0_u6_u7_n123, u0_u6_u7_n124, u0_u6_u7_n125, u0_u6_u7_n126, u0_u6_u7_n127, 
       u0_u6_u7_n128, u0_u6_u7_n129, u0_u6_u7_n130, u0_u6_u7_n131, u0_u6_u7_n132, u0_u6_u7_n133, u0_u6_u7_n134, u0_u6_u7_n135, u0_u6_u7_n136, 
       u0_u6_u7_n137, u0_u6_u7_n138, u0_u6_u7_n139, u0_u6_u7_n140, u0_u6_u7_n141, u0_u6_u7_n142, u0_u6_u7_n143, u0_u6_u7_n144, u0_u6_u7_n145, 
       u0_u6_u7_n146, u0_u6_u7_n147, u0_u6_u7_n148, u0_u6_u7_n149, u0_u6_u7_n150, u0_u6_u7_n151, u0_u6_u7_n152, u0_u6_u7_n153, u0_u6_u7_n154, 
       u0_u6_u7_n155, u0_u6_u7_n156, u0_u6_u7_n157, u0_u6_u7_n158, u0_u6_u7_n159, u0_u6_u7_n160, u0_u6_u7_n161, u0_u6_u7_n162, u0_u6_u7_n163, 
       u0_u6_u7_n164, u0_u6_u7_n165, u0_u6_u7_n166, u0_u6_u7_n167, u0_u6_u7_n168, u0_u6_u7_n169, u0_u6_u7_n170, u0_u6_u7_n171, u0_u6_u7_n172, 
       u0_u6_u7_n173, u0_u6_u7_n174, u0_u6_u7_n175, u0_u6_u7_n176, u0_u6_u7_n177, u0_u6_u7_n178, u0_u6_u7_n179, u0_u6_u7_n180, u0_u6_u7_n91, 
       u0_u6_u7_n92, u0_u6_u7_n93, u0_u6_u7_n94, u0_u6_u7_n95, u0_u6_u7_n96, u0_u6_u7_n97, u0_u6_u7_n98, u0_u6_u7_n99, u0_u7_X_43, 
       u0_u7_X_44, u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, u0_u7_u7_n100, u0_u7_u7_n101, u0_u7_u7_n102, u0_u7_u7_n103, 
       u0_u7_u7_n104, u0_u7_u7_n105, u0_u7_u7_n106, u0_u7_u7_n107, u0_u7_u7_n108, u0_u7_u7_n109, u0_u7_u7_n110, u0_u7_u7_n111, u0_u7_u7_n112, 
       u0_u7_u7_n113, u0_u7_u7_n114, u0_u7_u7_n115, u0_u7_u7_n116, u0_u7_u7_n117, u0_u7_u7_n118, u0_u7_u7_n119, u0_u7_u7_n120, u0_u7_u7_n121, 
       u0_u7_u7_n122, u0_u7_u7_n123, u0_u7_u7_n124, u0_u7_u7_n125, u0_u7_u7_n126, u0_u7_u7_n127, u0_u7_u7_n128, u0_u7_u7_n129, u0_u7_u7_n130, 
       u0_u7_u7_n131, u0_u7_u7_n132, u0_u7_u7_n133, u0_u7_u7_n134, u0_u7_u7_n135, u0_u7_u7_n136, u0_u7_u7_n137, u0_u7_u7_n138, u0_u7_u7_n139, 
       u0_u7_u7_n140, u0_u7_u7_n141, u0_u7_u7_n142, u0_u7_u7_n143, u0_u7_u7_n144, u0_u7_u7_n145, u0_u7_u7_n146, u0_u7_u7_n147, u0_u7_u7_n148, 
       u0_u7_u7_n149, u0_u7_u7_n150, u0_u7_u7_n151, u0_u7_u7_n152, u0_u7_u7_n153, u0_u7_u7_n154, u0_u7_u7_n155, u0_u7_u7_n156, u0_u7_u7_n157, 
       u0_u7_u7_n158, u0_u7_u7_n159, u0_u7_u7_n160, u0_u7_u7_n161, u0_u7_u7_n162, u0_u7_u7_n163, u0_u7_u7_n164, u0_u7_u7_n165, u0_u7_u7_n166, 
       u0_u7_u7_n167, u0_u7_u7_n168, u0_u7_u7_n169, u0_u7_u7_n170, u0_u7_u7_n171, u0_u7_u7_n172, u0_u7_u7_n173, u0_u7_u7_n174, u0_u7_u7_n175, 
       u0_u7_u7_n176, u0_u7_u7_n177, u0_u7_u7_n178, u0_u7_u7_n179, u0_u7_u7_n180, u0_u7_u7_n91, u0_u7_u7_n92, u0_u7_u7_n93, u0_u7_u7_n94, 
       u0_u7_u7_n95, u0_u7_u7_n96, u0_u7_u7_n97, u0_u7_u7_n98, u0_u7_u7_n99, u0_u9_X_19, u0_u9_X_20, u0_u9_X_21, u0_u9_X_22, 
       u0_u9_X_23, u0_u9_X_24, u0_u9_u3_n100, u0_u9_u3_n101, u0_u9_u3_n102, u0_u9_u3_n103, u0_u9_u3_n104, u0_u9_u3_n105, u0_u9_u3_n106, 
       u0_u9_u3_n107, u0_u9_u3_n108, u0_u9_u3_n109, u0_u9_u3_n110, u0_u9_u3_n111, u0_u9_u3_n112, u0_u9_u3_n113, u0_u9_u3_n114, u0_u9_u3_n115, 
       u0_u9_u3_n116, u0_u9_u3_n117, u0_u9_u3_n118, u0_u9_u3_n119, u0_u9_u3_n120, u0_u9_u3_n121, u0_u9_u3_n122, u0_u9_u3_n123, u0_u9_u3_n124, 
       u0_u9_u3_n125, u0_u9_u3_n126, u0_u9_u3_n127, u0_u9_u3_n128, u0_u9_u3_n129, u0_u9_u3_n130, u0_u9_u3_n131, u0_u9_u3_n132, u0_u9_u3_n133, 
       u0_u9_u3_n134, u0_u9_u3_n135, u0_u9_u3_n136, u0_u9_u3_n137, u0_u9_u3_n138, u0_u9_u3_n139, u0_u9_u3_n140, u0_u9_u3_n141, u0_u9_u3_n142, 
       u0_u9_u3_n143, u0_u9_u3_n144, u0_u9_u3_n145, u0_u9_u3_n146, u0_u9_u3_n147, u0_u9_u3_n148, u0_u9_u3_n149, u0_u9_u3_n150, u0_u9_u3_n151, 
       u0_u9_u3_n152, u0_u9_u3_n153, u0_u9_u3_n154, u0_u9_u3_n155, u0_u9_u3_n156, u0_u9_u3_n157, u0_u9_u3_n158, u0_u9_u3_n159, u0_u9_u3_n160, 
       u0_u9_u3_n161, u0_u9_u3_n162, u0_u9_u3_n163, u0_u9_u3_n164, u0_u9_u3_n165, u0_u9_u3_n166, u0_u9_u3_n167, u0_u9_u3_n168, u0_u9_u3_n169, 
       u0_u9_u3_n170, u0_u9_u3_n171, u0_u9_u3_n172, u0_u9_u3_n173, u0_u9_u3_n174, u0_u9_u3_n175, u0_u9_u3_n176, u0_u9_u3_n177, u0_u9_u3_n178, 
       u0_u9_u3_n179, u0_u9_u3_n180, u0_u9_u3_n181, u0_u9_u3_n182, u0_u9_u3_n183, u0_u9_u3_n184, u0_u9_u3_n185, u0_u9_u3_n186, u0_u9_u3_n94, 
       u0_u9_u3_n95, u0_u9_u3_n96, u0_u9_u3_n97, u0_u9_u3_n98, u0_u9_u3_n99, u0_uk_n1000, u0_uk_n1003, u0_uk_n1017, u0_uk_n1018, 
       u0_uk_n744, u0_uk_n745, u0_uk_n764, u0_uk_n776, u0_uk_n779, u0_uk_n781, u0_uk_n782, u0_uk_n783, u0_uk_n784, 
       u0_uk_n791, u0_uk_n792, u0_uk_n794, u0_uk_n795, u0_uk_n797, u0_uk_n819, u0_uk_n821, u0_uk_n822, u0_uk_n824, 
       u0_uk_n827, u0_uk_n828, u0_uk_n829, u0_uk_n831, u0_uk_n833, u0_uk_n835, u0_uk_n836, u0_uk_n837, u0_uk_n838, 
       u0_uk_n840, u0_uk_n846, u0_uk_n851, u0_uk_n858, u0_uk_n859, u0_uk_n860, u0_uk_n861, u0_uk_n862, u0_uk_n868, 
       u0_uk_n919, u0_uk_n920, u0_uk_n921, u0_uk_n949, u0_uk_n951, u0_uk_n953, u0_uk_n954, u0_uk_n955, u0_uk_n956, 
       u0_uk_n957, u0_uk_n958, u0_uk_n959, u0_uk_n982, u0_uk_n983, u0_uk_n985, u0_uk_n986, u0_uk_n987, u0_uk_n988, 
       u0_uk_n991, u0_uk_n992, u0_uk_n996, u0_uk_n997, u1_K2_19, u1_K2_20, u1_K2_21, u1_K2_22, u1_K2_23, 
       u1_K2_24, u1_out1_1, u1_out1_10, u1_out1_20, u1_out1_26, u1_u1_X_19, u1_u1_X_20, u1_u1_X_21, u1_u1_X_22, 
       u1_u1_X_23, u1_u1_X_24, u1_u1_u3_n100, u1_u1_u3_n101, u1_u1_u3_n102, u1_u1_u3_n103, u1_u1_u3_n104, u1_u1_u3_n105, u1_u1_u3_n106, 
       u1_u1_u3_n107, u1_u1_u3_n108, u1_u1_u3_n109, u1_u1_u3_n110, u1_u1_u3_n111, u1_u1_u3_n112, u1_u1_u3_n113, u1_u1_u3_n114, u1_u1_u3_n115, 
       u1_u1_u3_n116, u1_u1_u3_n117, u1_u1_u3_n118, u1_u1_u3_n119, u1_u1_u3_n120, u1_u1_u3_n121, u1_u1_u3_n122, u1_u1_u3_n123, u1_u1_u3_n124, 
       u1_u1_u3_n125, u1_u1_u3_n126, u1_u1_u3_n127, u1_u1_u3_n128, u1_u1_u3_n129, u1_u1_u3_n130, u1_u1_u3_n131, u1_u1_u3_n132, u1_u1_u3_n133, 
       u1_u1_u3_n134, u1_u1_u3_n135, u1_u1_u3_n136, u1_u1_u3_n137, u1_u1_u3_n138, u1_u1_u3_n139, u1_u1_u3_n140, u1_u1_u3_n141, u1_u1_u3_n142, 
       u1_u1_u3_n143, u1_u1_u3_n144, u1_u1_u3_n145, u1_u1_u3_n146, u1_u1_u3_n147, u1_u1_u3_n148, u1_u1_u3_n149, u1_u1_u3_n150, u1_u1_u3_n151, 
       u1_u1_u3_n152, u1_u1_u3_n153, u1_u1_u3_n154, u1_u1_u3_n155, u1_u1_u3_n156, u1_u1_u3_n157, u1_u1_u3_n158, u1_u1_u3_n159, u1_u1_u3_n160, 
       u1_u1_u3_n161, u1_u1_u3_n162, u1_u1_u3_n163, u1_u1_u3_n164, u1_u1_u3_n165, u1_u1_u3_n166, u1_u1_u3_n167, u1_u1_u3_n168, u1_u1_u3_n169, 
       u1_u1_u3_n170, u1_u1_u3_n171, u1_u1_u3_n172, u1_u1_u3_n173, u1_u1_u3_n174, u1_u1_u3_n175, u1_u1_u3_n176, u1_u1_u3_n177, u1_u1_u3_n178, 
       u1_u1_u3_n179, u1_u1_u3_n180, u1_u1_u3_n181, u1_u1_u3_n182, u1_u1_u3_n183, u1_u1_u3_n184, u1_u1_u3_n185, u1_u1_u3_n186, u1_u1_u3_n94, 
       u1_u1_u3_n95, u1_u1_u3_n96, u1_u1_u3_n97, u1_u1_u3_n98, u1_u1_u3_n99, u1_uk_n1025, u2_K10_12, u2_K10_13, u2_K10_14, 
       u2_K10_16, u2_K10_18, u2_K10_7, u2_K10_8, u2_K10_9, u2_K11_31, u2_K11_32, u2_K11_33, u2_K11_34, 
       u2_K11_35, u2_K11_36, u2_K11_37, u2_K11_39, u2_K11_40, u2_K11_41, u2_K12_28, u2_K12_30, u2_K12_31, 
       u2_K12_32, u2_K12_33, u2_K12_35, u2_K12_36, u2_K12_38, u2_K12_39, u2_K12_40, u2_K12_42, u2_K12_43, 
       u2_K12_44, u2_K12_45, u2_K12_48, u2_K15_10, u2_K15_11, u2_K15_12, u2_K15_14, u2_K15_15, u2_K15_17, 
       u2_K15_19, u2_K15_22, u2_K15_24, u2_K15_3, u2_K15_4, u2_K15_6, u2_K15_7, u2_K15_8, u2_K15_9, 
       u2_K16_1, u2_K16_10, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_15, u2_K16_16, u2_K16_17, 
       u2_K16_18, u2_K16_19, u2_K16_2, u2_K16_20, u2_K16_21, u2_K16_22, u2_K16_23, u2_K16_24, u2_K16_3, 
       u2_K16_4, u2_K16_7, u2_K1_10, u2_K1_11, u2_K1_12, u2_K1_13, u2_K1_14, u2_K1_17, u2_K1_18, 
       u2_K1_2, u2_K1_3, u2_K1_4, u2_K1_6, u2_K1_7, u2_K1_8, u2_K2_10, u2_K2_11, u2_K2_12, 
       u2_K2_2, u2_K2_3, u2_K2_4, u2_K2_5, u2_K2_6, u2_K2_7, u2_K2_8, u2_K2_9, u2_K6_17, 
       u2_K6_18, u2_K6_19, u2_K6_21, u2_K6_23, u2_K6_31, u2_K6_33, u2_K6_35, u2_K6_37, u2_K6_38, 
       u2_K6_39, u2_K6_41, u2_K6_42, u2_K7_1, u2_K7_10, u2_K7_11, u2_K7_12, u2_K7_13, u2_K7_14, 
       u2_K7_15, u2_K7_16, u2_K7_17, u2_K7_18, u2_K7_2, u2_K7_6, u2_K7_8, u2_K7_9, u2_out0_13, 
       u2_out0_16, u2_out0_17, u2_out0_18, u2_out0_2, u2_out0_23, u2_out0_24, u2_out0_28, u2_out0_30, u2_out0_31, 
       u2_out0_6, u2_out0_9, u2_out10_11, u2_out10_12, u2_out10_19, u2_out10_22, u2_out10_29, u2_out10_32, u2_out10_4, 
       u2_out10_7, u2_out11_11, u2_out11_12, u2_out11_14, u2_out11_15, u2_out11_19, u2_out11_21, u2_out11_22, u2_out11_25, 
       u2_out11_27, u2_out11_29, u2_out11_3, u2_out11_32, u2_out11_4, u2_out11_5, u2_out11_7, u2_out11_8, u2_out14_1, 
       u2_out14_10, u2_out14_13, u2_out14_16, u2_out14_17, u2_out14_18, u2_out14_2, u2_out14_20, u2_out14_23, u2_out14_24, 
       u2_out14_26, u2_out14_28, u2_out14_30, u2_out14_31, u2_out14_6, u2_out14_9, u2_out15_1, u2_out15_10, u2_out15_13, 
       u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_2, u2_out15_20, u2_out15_23, u2_out15_24, u2_out15_26, u2_out15_28, 
       u2_out15_30, u2_out15_31, u2_out15_6, u2_out15_9, u2_out1_13, u2_out1_17, u2_out1_18, u2_out1_2, u2_out1_23, 
       u2_out1_28, u2_out1_31, u2_out1_9, u2_out5_1, u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_16, u2_out5_19, 
       u2_out5_20, u2_out5_22, u2_out5_24, u2_out5_26, u2_out5_29, u2_out5_30, u2_out5_32, u2_out5_4, u2_out5_6, 
       u2_out5_7, u2_out6_13, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_2, u2_out6_23, u2_out6_24, u2_out6_28, 
       u2_out6_30, u2_out6_31, u2_out6_6, u2_out6_9, u2_out9_13, u2_out9_16, u2_out9_18, u2_out9_2, u2_out9_24, 
       u2_out9_28, u2_out9_30, u2_out9_6, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, u2_u0_X_13, u2_u0_X_14, u2_u0_X_15, 
       u2_u0_X_16, u2_u0_X_17, u2_u0_X_18, u2_u0_X_2, u2_u0_X_3, u2_u0_X_4, u2_u0_X_5, u2_u0_X_6, u2_u0_X_7, 
       u2_u0_X_8, u2_u0_X_9, u2_u0_u0_n100, u2_u0_u0_n101, u2_u0_u0_n102, u2_u0_u0_n103, u2_u0_u0_n104, u2_u0_u0_n105, u2_u0_u0_n106, 
       u2_u0_u0_n107, u2_u0_u0_n108, u2_u0_u0_n109, u2_u0_u0_n110, u2_u0_u0_n111, u2_u0_u0_n112, u2_u0_u0_n113, u2_u0_u0_n114, u2_u0_u0_n115, 
       u2_u0_u0_n116, u2_u0_u0_n117, u2_u0_u0_n118, u2_u0_u0_n119, u2_u0_u0_n120, u2_u0_u0_n121, u2_u0_u0_n122, u2_u0_u0_n123, u2_u0_u0_n124, 
       u2_u0_u0_n125, u2_u0_u0_n126, u2_u0_u0_n127, u2_u0_u0_n128, u2_u0_u0_n129, u2_u0_u0_n130, u2_u0_u0_n131, u2_u0_u0_n132, u2_u0_u0_n133, 
       u2_u0_u0_n134, u2_u0_u0_n135, u2_u0_u0_n136, u2_u0_u0_n137, u2_u0_u0_n138, u2_u0_u0_n139, u2_u0_u0_n140, u2_u0_u0_n141, u2_u0_u0_n142, 
       u2_u0_u0_n143, u2_u0_u0_n144, u2_u0_u0_n145, u2_u0_u0_n146, u2_u0_u0_n147, u2_u0_u0_n148, u2_u0_u0_n149, u2_u0_u0_n150, u2_u0_u0_n151, 
       u2_u0_u0_n152, u2_u0_u0_n153, u2_u0_u0_n154, u2_u0_u0_n155, u2_u0_u0_n156, u2_u0_u0_n157, u2_u0_u0_n158, u2_u0_u0_n159, u2_u0_u0_n160, 
       u2_u0_u0_n161, u2_u0_u0_n162, u2_u0_u0_n163, u2_u0_u0_n164, u2_u0_u0_n165, u2_u0_u0_n166, u2_u0_u0_n167, u2_u0_u0_n168, u2_u0_u0_n169, 
       u2_u0_u0_n170, u2_u0_u0_n171, u2_u0_u0_n172, u2_u0_u0_n173, u2_u0_u0_n174, u2_u0_u0_n88, u2_u0_u0_n89, u2_u0_u0_n90, u2_u0_u0_n91, 
       u2_u0_u0_n92, u2_u0_u0_n93, u2_u0_u0_n94, u2_u0_u0_n95, u2_u0_u0_n96, u2_u0_u0_n97, u2_u0_u0_n98, u2_u0_u0_n99, u2_u0_u1_n100, 
       u2_u0_u1_n101, u2_u0_u1_n102, u2_u0_u1_n103, u2_u0_u1_n104, u2_u0_u1_n105, u2_u0_u1_n106, u2_u0_u1_n107, u2_u0_u1_n108, u2_u0_u1_n109, 
       u2_u0_u1_n110, u2_u0_u1_n111, u2_u0_u1_n112, u2_u0_u1_n113, u2_u0_u1_n114, u2_u0_u1_n115, u2_u0_u1_n116, u2_u0_u1_n117, u2_u0_u1_n118, 
       u2_u0_u1_n119, u2_u0_u1_n120, u2_u0_u1_n121, u2_u0_u1_n122, u2_u0_u1_n123, u2_u0_u1_n124, u2_u0_u1_n125, u2_u0_u1_n126, u2_u0_u1_n127, 
       u2_u0_u1_n128, u2_u0_u1_n129, u2_u0_u1_n130, u2_u0_u1_n131, u2_u0_u1_n132, u2_u0_u1_n133, u2_u0_u1_n134, u2_u0_u1_n135, u2_u0_u1_n136, 
       u2_u0_u1_n137, u2_u0_u1_n138, u2_u0_u1_n139, u2_u0_u1_n140, u2_u0_u1_n141, u2_u0_u1_n142, u2_u0_u1_n143, u2_u0_u1_n144, u2_u0_u1_n145, 
       u2_u0_u1_n146, u2_u0_u1_n147, u2_u0_u1_n148, u2_u0_u1_n149, u2_u0_u1_n150, u2_u0_u1_n151, u2_u0_u1_n152, u2_u0_u1_n153, u2_u0_u1_n154, 
       u2_u0_u1_n155, u2_u0_u1_n156, u2_u0_u1_n157, u2_u0_u1_n158, u2_u0_u1_n159, u2_u0_u1_n160, u2_u0_u1_n161, u2_u0_u1_n162, u2_u0_u1_n163, 
       u2_u0_u1_n164, u2_u0_u1_n165, u2_u0_u1_n166, u2_u0_u1_n167, u2_u0_u1_n168, u2_u0_u1_n169, u2_u0_u1_n170, u2_u0_u1_n171, u2_u0_u1_n172, 
       u2_u0_u1_n173, u2_u0_u1_n174, u2_u0_u1_n175, u2_u0_u1_n176, u2_u0_u1_n177, u2_u0_u1_n178, u2_u0_u1_n179, u2_u0_u1_n180, u2_u0_u1_n181, 
       u2_u0_u1_n182, u2_u0_u1_n183, u2_u0_u1_n184, u2_u0_u1_n185, u2_u0_u1_n186, u2_u0_u1_n187, u2_u0_u1_n188, u2_u0_u1_n95, u2_u0_u1_n96, 
       u2_u0_u1_n97, u2_u0_u1_n98, u2_u0_u1_n99, u2_u0_u2_n100, u2_u0_u2_n101, u2_u0_u2_n102, u2_u0_u2_n103, u2_u0_u2_n104, u2_u0_u2_n105, 
       u2_u0_u2_n106, u2_u0_u2_n107, u2_u0_u2_n108, u2_u0_u2_n109, u2_u0_u2_n110, u2_u0_u2_n111, u2_u0_u2_n112, u2_u0_u2_n113, u2_u0_u2_n114, 
       u2_u0_u2_n115, u2_u0_u2_n116, u2_u0_u2_n117, u2_u0_u2_n118, u2_u0_u2_n119, u2_u0_u2_n120, u2_u0_u2_n121, u2_u0_u2_n122, u2_u0_u2_n123, 
       u2_u0_u2_n124, u2_u0_u2_n125, u2_u0_u2_n126, u2_u0_u2_n127, u2_u0_u2_n128, u2_u0_u2_n129, u2_u0_u2_n130, u2_u0_u2_n131, u2_u0_u2_n132, 
       u2_u0_u2_n133, u2_u0_u2_n134, u2_u0_u2_n135, u2_u0_u2_n136, u2_u0_u2_n137, u2_u0_u2_n138, u2_u0_u2_n139, u2_u0_u2_n140, u2_u0_u2_n141, 
       u2_u0_u2_n142, u2_u0_u2_n143, u2_u0_u2_n144, u2_u0_u2_n145, u2_u0_u2_n146, u2_u0_u2_n147, u2_u0_u2_n148, u2_u0_u2_n149, u2_u0_u2_n150, 
       u2_u0_u2_n151, u2_u0_u2_n152, u2_u0_u2_n153, u2_u0_u2_n154, u2_u0_u2_n155, u2_u0_u2_n156, u2_u0_u2_n157, u2_u0_u2_n158, u2_u0_u2_n159, 
       u2_u0_u2_n160, u2_u0_u2_n161, u2_u0_u2_n162, u2_u0_u2_n163, u2_u0_u2_n164, u2_u0_u2_n165, u2_u0_u2_n166, u2_u0_u2_n167, u2_u0_u2_n168, 
       u2_u0_u2_n169, u2_u0_u2_n170, u2_u0_u2_n171, u2_u0_u2_n172, u2_u0_u2_n173, u2_u0_u2_n174, u2_u0_u2_n175, u2_u0_u2_n176, u2_u0_u2_n177, 
       u2_u0_u2_n178, u2_u0_u2_n179, u2_u0_u2_n180, u2_u0_u2_n181, u2_u0_u2_n182, u2_u0_u2_n183, u2_u0_u2_n184, u2_u0_u2_n185, u2_u0_u2_n186, 
       u2_u0_u2_n187, u2_u0_u2_n188, u2_u0_u2_n95, u2_u0_u2_n96, u2_u0_u2_n97, u2_u0_u2_n98, u2_u0_u2_n99, u2_u10_X_31, u2_u10_X_32, 
       u2_u10_X_33, u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, 
       u2_u10_X_42, u2_u10_u5_n100, u2_u10_u5_n101, u2_u10_u5_n102, u2_u10_u5_n103, u2_u10_u5_n104, u2_u10_u5_n105, u2_u10_u5_n106, u2_u10_u5_n107, 
       u2_u10_u5_n108, u2_u10_u5_n109, u2_u10_u5_n110, u2_u10_u5_n111, u2_u10_u5_n112, u2_u10_u5_n113, u2_u10_u5_n114, u2_u10_u5_n115, u2_u10_u5_n116, 
       u2_u10_u5_n117, u2_u10_u5_n118, u2_u10_u5_n119, u2_u10_u5_n120, u2_u10_u5_n121, u2_u10_u5_n122, u2_u10_u5_n123, u2_u10_u5_n124, u2_u10_u5_n125, 
       u2_u10_u5_n126, u2_u10_u5_n127, u2_u10_u5_n128, u2_u10_u5_n129, u2_u10_u5_n130, u2_u10_u5_n131, u2_u10_u5_n132, u2_u10_u5_n133, u2_u10_u5_n134, 
       u2_u10_u5_n135, u2_u10_u5_n136, u2_u10_u5_n137, u2_u10_u5_n138, u2_u10_u5_n139, u2_u10_u5_n140, u2_u10_u5_n141, u2_u10_u5_n142, u2_u10_u5_n143, 
       u2_u10_u5_n144, u2_u10_u5_n145, u2_u10_u5_n146, u2_u10_u5_n147, u2_u10_u5_n148, u2_u10_u5_n149, u2_u10_u5_n150, u2_u10_u5_n151, u2_u10_u5_n152, 
       u2_u10_u5_n153, u2_u10_u5_n154, u2_u10_u5_n155, u2_u10_u5_n156, u2_u10_u5_n157, u2_u10_u5_n158, u2_u10_u5_n159, u2_u10_u5_n160, u2_u10_u5_n161, 
       u2_u10_u5_n162, u2_u10_u5_n163, u2_u10_u5_n164, u2_u10_u5_n165, u2_u10_u5_n166, u2_u10_u5_n167, u2_u10_u5_n168, u2_u10_u5_n169, u2_u10_u5_n170, 
       u2_u10_u5_n171, u2_u10_u5_n172, u2_u10_u5_n173, u2_u10_u5_n174, u2_u10_u5_n175, u2_u10_u5_n176, u2_u10_u5_n177, u2_u10_u5_n178, u2_u10_u5_n179, 
       u2_u10_u5_n180, u2_u10_u5_n181, u2_u10_u5_n182, u2_u10_u5_n183, u2_u10_u5_n184, u2_u10_u5_n185, u2_u10_u5_n186, u2_u10_u5_n187, u2_u10_u5_n188, 
       u2_u10_u5_n189, u2_u10_u5_n190, u2_u10_u5_n191, u2_u10_u5_n192, u2_u10_u5_n193, u2_u10_u5_n194, u2_u10_u5_n195, u2_u10_u5_n196, u2_u10_u5_n99, 
       u2_u10_u6_n100, u2_u10_u6_n101, u2_u10_u6_n102, u2_u10_u6_n103, u2_u10_u6_n104, u2_u10_u6_n105, u2_u10_u6_n106, u2_u10_u6_n107, u2_u10_u6_n108, 
       u2_u10_u6_n109, u2_u10_u6_n110, u2_u10_u6_n111, u2_u10_u6_n112, u2_u10_u6_n113, u2_u10_u6_n114, u2_u10_u6_n115, u2_u10_u6_n116, u2_u10_u6_n117, 
       u2_u10_u6_n118, u2_u10_u6_n119, u2_u10_u6_n120, u2_u10_u6_n121, u2_u10_u6_n122, u2_u10_u6_n123, u2_u10_u6_n124, u2_u10_u6_n125, u2_u10_u6_n126, 
       u2_u10_u6_n127, u2_u10_u6_n128, u2_u10_u6_n129, u2_u10_u6_n130, u2_u10_u6_n131, u2_u10_u6_n132, u2_u10_u6_n133, u2_u10_u6_n134, u2_u10_u6_n135, 
       u2_u10_u6_n136, u2_u10_u6_n137, u2_u10_u6_n138, u2_u10_u6_n139, u2_u10_u6_n140, u2_u10_u6_n141, u2_u10_u6_n142, u2_u10_u6_n143, u2_u10_u6_n144, 
       u2_u10_u6_n145, u2_u10_u6_n146, u2_u10_u6_n147, u2_u10_u6_n148, u2_u10_u6_n149, u2_u10_u6_n150, u2_u10_u6_n151, u2_u10_u6_n152, u2_u10_u6_n153, 
       u2_u10_u6_n154, u2_u10_u6_n155, u2_u10_u6_n156, u2_u10_u6_n157, u2_u10_u6_n158, u2_u10_u6_n159, u2_u10_u6_n160, u2_u10_u6_n161, u2_u10_u6_n162, 
       u2_u10_u6_n163, u2_u10_u6_n164, u2_u10_u6_n165, u2_u10_u6_n166, u2_u10_u6_n167, u2_u10_u6_n168, u2_u10_u6_n169, u2_u10_u6_n170, u2_u10_u6_n171, 
       u2_u10_u6_n172, u2_u10_u6_n173, u2_u10_u6_n174, u2_u10_u6_n88, u2_u10_u6_n89, u2_u10_u6_n90, u2_u10_u6_n91, u2_u10_u6_n92, u2_u10_u6_n93, 
       u2_u10_u6_n94, u2_u10_u6_n95, u2_u10_u6_n96, u2_u10_u6_n97, u2_u10_u6_n98, u2_u10_u6_n99, u2_u11_X_25, u2_u11_X_26, u2_u11_X_27, 
       u2_u11_X_28, u2_u11_X_29, u2_u11_X_30, u2_u11_X_31, u2_u11_X_32, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_36, 
       u2_u11_X_37, u2_u11_X_38, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, u2_u11_X_42, u2_u11_X_43, u2_u11_X_44, u2_u11_X_45, 
       u2_u11_X_46, u2_u11_X_47, u2_u11_X_48, u2_u11_u4_n100, u2_u11_u4_n101, u2_u11_u4_n102, u2_u11_u4_n103, u2_u11_u4_n104, u2_u11_u4_n105, 
       u2_u11_u4_n106, u2_u11_u4_n107, u2_u11_u4_n108, u2_u11_u4_n109, u2_u11_u4_n110, u2_u11_u4_n111, u2_u11_u4_n112, u2_u11_u4_n113, u2_u11_u4_n114, 
       u2_u11_u4_n115, u2_u11_u4_n116, u2_u11_u4_n117, u2_u11_u4_n118, u2_u11_u4_n119, u2_u11_u4_n120, u2_u11_u4_n121, u2_u11_u4_n122, u2_u11_u4_n123, 
       u2_u11_u4_n124, u2_u11_u4_n125, u2_u11_u4_n126, u2_u11_u4_n127, u2_u11_u4_n128, u2_u11_u4_n129, u2_u11_u4_n130, u2_u11_u4_n131, u2_u11_u4_n132, 
       u2_u11_u4_n133, u2_u11_u4_n134, u2_u11_u4_n135, u2_u11_u4_n136, u2_u11_u4_n137, u2_u11_u4_n138, u2_u11_u4_n139, u2_u11_u4_n140, u2_u11_u4_n141, 
       u2_u11_u4_n142, u2_u11_u4_n143, u2_u11_u4_n144, u2_u11_u4_n145, u2_u11_u4_n146, u2_u11_u4_n147, u2_u11_u4_n148, u2_u11_u4_n149, u2_u11_u4_n150, 
       u2_u11_u4_n151, u2_u11_u4_n152, u2_u11_u4_n153, u2_u11_u4_n154, u2_u11_u4_n155, u2_u11_u4_n156, u2_u11_u4_n157, u2_u11_u4_n158, u2_u11_u4_n159, 
       u2_u11_u4_n160, u2_u11_u4_n161, u2_u11_u4_n162, u2_u11_u4_n163, u2_u11_u4_n164, u2_u11_u4_n165, u2_u11_u4_n166, u2_u11_u4_n167, u2_u11_u4_n168, 
       u2_u11_u4_n169, u2_u11_u4_n170, u2_u11_u4_n171, u2_u11_u4_n172, u2_u11_u4_n173, u2_u11_u4_n174, u2_u11_u4_n175, u2_u11_u4_n176, u2_u11_u4_n177, 
       u2_u11_u4_n178, u2_u11_u4_n179, u2_u11_u4_n180, u2_u11_u4_n181, u2_u11_u4_n182, u2_u11_u4_n183, u2_u11_u4_n184, u2_u11_u4_n185, u2_u11_u4_n186, 
       u2_u11_u4_n94, u2_u11_u4_n95, u2_u11_u4_n96, u2_u11_u4_n97, u2_u11_u4_n98, u2_u11_u4_n99, u2_u11_u5_n100, u2_u11_u5_n101, u2_u11_u5_n102, 
       u2_u11_u5_n103, u2_u11_u5_n104, u2_u11_u5_n105, u2_u11_u5_n106, u2_u11_u5_n107, u2_u11_u5_n108, u2_u11_u5_n109, u2_u11_u5_n110, u2_u11_u5_n111, 
       u2_u11_u5_n112, u2_u11_u5_n113, u2_u11_u5_n114, u2_u11_u5_n115, u2_u11_u5_n116, u2_u11_u5_n117, u2_u11_u5_n118, u2_u11_u5_n119, u2_u11_u5_n120, 
       u2_u11_u5_n121, u2_u11_u5_n122, u2_u11_u5_n123, u2_u11_u5_n124, u2_u11_u5_n125, u2_u11_u5_n126, u2_u11_u5_n127, u2_u11_u5_n128, u2_u11_u5_n129, 
       u2_u11_u5_n130, u2_u11_u5_n131, u2_u11_u5_n132, u2_u11_u5_n133, u2_u11_u5_n134, u2_u11_u5_n135, u2_u11_u5_n136, u2_u11_u5_n137, u2_u11_u5_n138, 
       u2_u11_u5_n139, u2_u11_u5_n140, u2_u11_u5_n141, u2_u11_u5_n142, u2_u11_u5_n143, u2_u11_u5_n144, u2_u11_u5_n145, u2_u11_u5_n146, u2_u11_u5_n147, 
       u2_u11_u5_n148, u2_u11_u5_n149, u2_u11_u5_n150, u2_u11_u5_n151, u2_u11_u5_n152, u2_u11_u5_n153, u2_u11_u5_n154, u2_u11_u5_n155, u2_u11_u5_n156, 
       u2_u11_u5_n157, u2_u11_u5_n158, u2_u11_u5_n159, u2_u11_u5_n160, u2_u11_u5_n161, u2_u11_u5_n162, u2_u11_u5_n163, u2_u11_u5_n164, u2_u11_u5_n165, 
       u2_u11_u5_n166, u2_u11_u5_n167, u2_u11_u5_n168, u2_u11_u5_n169, u2_u11_u5_n170, u2_u11_u5_n171, u2_u11_u5_n172, u2_u11_u5_n173, u2_u11_u5_n174, 
       u2_u11_u5_n175, u2_u11_u5_n176, u2_u11_u5_n177, u2_u11_u5_n178, u2_u11_u5_n179, u2_u11_u5_n180, u2_u11_u5_n181, u2_u11_u5_n182, u2_u11_u5_n183, 
       u2_u11_u5_n184, u2_u11_u5_n185, u2_u11_u5_n186, u2_u11_u5_n187, u2_u11_u5_n188, u2_u11_u5_n189, u2_u11_u5_n190, u2_u11_u5_n191, u2_u11_u5_n192, 
       u2_u11_u5_n193, u2_u11_u5_n194, u2_u11_u5_n195, u2_u11_u5_n196, u2_u11_u5_n99, u2_u11_u6_n100, u2_u11_u6_n101, u2_u11_u6_n102, u2_u11_u6_n103, 
       u2_u11_u6_n104, u2_u11_u6_n105, u2_u11_u6_n106, u2_u11_u6_n107, u2_u11_u6_n108, u2_u11_u6_n109, u2_u11_u6_n110, u2_u11_u6_n111, u2_u11_u6_n112, 
       u2_u11_u6_n113, u2_u11_u6_n114, u2_u11_u6_n115, u2_u11_u6_n116, u2_u11_u6_n117, u2_u11_u6_n118, u2_u11_u6_n119, u2_u11_u6_n120, u2_u11_u6_n121, 
       u2_u11_u6_n122, u2_u11_u6_n123, u2_u11_u6_n124, u2_u11_u6_n125, u2_u11_u6_n126, u2_u11_u6_n127, u2_u11_u6_n128, u2_u11_u6_n129, u2_u11_u6_n130, 
       u2_u11_u6_n131, u2_u11_u6_n132, u2_u11_u6_n133, u2_u11_u6_n134, u2_u11_u6_n135, u2_u11_u6_n136, u2_u11_u6_n137, u2_u11_u6_n138, u2_u11_u6_n139, 
       u2_u11_u6_n140, u2_u11_u6_n141, u2_u11_u6_n142, u2_u11_u6_n143, u2_u11_u6_n144, u2_u11_u6_n145, u2_u11_u6_n146, u2_u11_u6_n147, u2_u11_u6_n148, 
       u2_u11_u6_n149, u2_u11_u6_n150, u2_u11_u6_n151, u2_u11_u6_n152, u2_u11_u6_n153, u2_u11_u6_n154, u2_u11_u6_n155, u2_u11_u6_n156, u2_u11_u6_n157, 
       u2_u11_u6_n158, u2_u11_u6_n159, u2_u11_u6_n160, u2_u11_u6_n161, u2_u11_u6_n162, u2_u11_u6_n163, u2_u11_u6_n164, u2_u11_u6_n165, u2_u11_u6_n166, 
       u2_u11_u6_n167, u2_u11_u6_n168, u2_u11_u6_n169, u2_u11_u6_n170, u2_u11_u6_n171, u2_u11_u6_n172, u2_u11_u6_n173, u2_u11_u6_n174, u2_u11_u6_n88, 
       u2_u11_u6_n89, u2_u11_u6_n90, u2_u11_u6_n91, u2_u11_u6_n92, u2_u11_u6_n93, u2_u11_u6_n94, u2_u11_u6_n95, u2_u11_u6_n96, u2_u11_u6_n97, 
       u2_u11_u6_n98, u2_u11_u6_n99, u2_u11_u7_n100, u2_u11_u7_n101, u2_u11_u7_n102, u2_u11_u7_n103, u2_u11_u7_n104, u2_u11_u7_n105, u2_u11_u7_n106, 
       u2_u11_u7_n107, u2_u11_u7_n108, u2_u11_u7_n109, u2_u11_u7_n110, u2_u11_u7_n111, u2_u11_u7_n112, u2_u11_u7_n113, u2_u11_u7_n114, u2_u11_u7_n115, 
       u2_u11_u7_n116, u2_u11_u7_n117, u2_u11_u7_n118, u2_u11_u7_n119, u2_u11_u7_n120, u2_u11_u7_n121, u2_u11_u7_n122, u2_u11_u7_n123, u2_u11_u7_n124, 
       u2_u11_u7_n125, u2_u11_u7_n126, u2_u11_u7_n127, u2_u11_u7_n128, u2_u11_u7_n129, u2_u11_u7_n130, u2_u11_u7_n131, u2_u11_u7_n132, u2_u11_u7_n133, 
       u2_u11_u7_n134, u2_u11_u7_n135, u2_u11_u7_n136, u2_u11_u7_n137, u2_u11_u7_n138, u2_u11_u7_n139, u2_u11_u7_n140, u2_u11_u7_n141, u2_u11_u7_n142, 
       u2_u11_u7_n143, u2_u11_u7_n144, u2_u11_u7_n145, u2_u11_u7_n146, u2_u11_u7_n147, u2_u11_u7_n148, u2_u11_u7_n149, u2_u11_u7_n150, u2_u11_u7_n151, 
       u2_u11_u7_n152, u2_u11_u7_n153, u2_u11_u7_n154, u2_u11_u7_n155, u2_u11_u7_n156, u2_u11_u7_n157, u2_u11_u7_n158, u2_u11_u7_n159, u2_u11_u7_n160, 
       u2_u11_u7_n161, u2_u11_u7_n162, u2_u11_u7_n163, u2_u11_u7_n164, u2_u11_u7_n165, u2_u11_u7_n166, u2_u11_u7_n167, u2_u11_u7_n168, u2_u11_u7_n169, 
       u2_u11_u7_n170, u2_u11_u7_n171, u2_u11_u7_n172, u2_u11_u7_n173, u2_u11_u7_n174, u2_u11_u7_n175, u2_u11_u7_n176, u2_u11_u7_n177, u2_u11_u7_n178, 
       u2_u11_u7_n179, u2_u11_u7_n180, u2_u11_u7_n91, u2_u11_u7_n92, u2_u11_u7_n93, u2_u11_u7_n94, u2_u11_u7_n95, u2_u11_u7_n96, u2_u11_u7_n97, 
       u2_u11_u7_n98, u2_u11_u7_n99, u2_u14_X_1, u2_u14_X_10, u2_u14_X_11, u2_u14_X_12, u2_u14_X_13, u2_u14_X_14, u2_u14_X_15, 
       u2_u14_X_16, u2_u14_X_17, u2_u14_X_18, u2_u14_X_19, u2_u14_X_2, u2_u14_X_20, u2_u14_X_21, u2_u14_X_22, u2_u14_X_23, 
       u2_u14_X_24, u2_u14_X_3, u2_u14_X_4, u2_u14_X_5, u2_u14_X_6, u2_u14_X_7, u2_u14_X_8, u2_u14_X_9, u2_u14_u0_n100, 
       u2_u14_u0_n101, u2_u14_u0_n102, u2_u14_u0_n103, u2_u14_u0_n104, u2_u14_u0_n105, u2_u14_u0_n106, u2_u14_u0_n107, u2_u14_u0_n108, u2_u14_u0_n109, 
       u2_u14_u0_n110, u2_u14_u0_n111, u2_u14_u0_n112, u2_u14_u0_n113, u2_u14_u0_n114, u2_u14_u0_n115, u2_u14_u0_n116, u2_u14_u0_n117, u2_u14_u0_n118, 
       u2_u14_u0_n119, u2_u14_u0_n120, u2_u14_u0_n121, u2_u14_u0_n122, u2_u14_u0_n123, u2_u14_u0_n124, u2_u14_u0_n125, u2_u14_u0_n126, u2_u14_u0_n127, 
       u2_u14_u0_n128, u2_u14_u0_n129, u2_u14_u0_n130, u2_u14_u0_n131, u2_u14_u0_n132, u2_u14_u0_n133, u2_u14_u0_n134, u2_u14_u0_n135, u2_u14_u0_n136, 
       u2_u14_u0_n137, u2_u14_u0_n138, u2_u14_u0_n139, u2_u14_u0_n140, u2_u14_u0_n141, u2_u14_u0_n142, u2_u14_u0_n143, u2_u14_u0_n144, u2_u14_u0_n145, 
       u2_u14_u0_n146, u2_u14_u0_n147, u2_u14_u0_n148, u2_u14_u0_n149, u2_u14_u0_n150, u2_u14_u0_n151, u2_u14_u0_n152, u2_u14_u0_n153, u2_u14_u0_n154, 
       u2_u14_u0_n155, u2_u14_u0_n156, u2_u14_u0_n157, u2_u14_u0_n158, u2_u14_u0_n159, u2_u14_u0_n160, u2_u14_u0_n161, u2_u14_u0_n162, u2_u14_u0_n163, 
       u2_u14_u0_n164, u2_u14_u0_n165, u2_u14_u0_n166, u2_u14_u0_n167, u2_u14_u0_n168, u2_u14_u0_n169, u2_u14_u0_n170, u2_u14_u0_n171, u2_u14_u0_n172, 
       u2_u14_u0_n173, u2_u14_u0_n174, u2_u14_u0_n88, u2_u14_u0_n89, u2_u14_u0_n90, u2_u14_u0_n91, u2_u14_u0_n92, u2_u14_u0_n93, u2_u14_u0_n94, 
       u2_u14_u0_n95, u2_u14_u0_n96, u2_u14_u0_n97, u2_u14_u0_n98, u2_u14_u0_n99, u2_u14_u1_n100, u2_u14_u1_n101, u2_u14_u1_n102, u2_u14_u1_n103, 
       u2_u14_u1_n104, u2_u14_u1_n105, u2_u14_u1_n106, u2_u14_u1_n107, u2_u14_u1_n108, u2_u14_u1_n109, u2_u14_u1_n110, u2_u14_u1_n111, u2_u14_u1_n112, 
       u2_u14_u1_n113, u2_u14_u1_n114, u2_u14_u1_n115, u2_u14_u1_n116, u2_u14_u1_n117, u2_u14_u1_n118, u2_u14_u1_n119, u2_u14_u1_n120, u2_u14_u1_n121, 
       u2_u14_u1_n122, u2_u14_u1_n123, u2_u14_u1_n124, u2_u14_u1_n125, u2_u14_u1_n126, u2_u14_u1_n127, u2_u14_u1_n128, u2_u14_u1_n129, u2_u14_u1_n130, 
       u2_u14_u1_n131, u2_u14_u1_n132, u2_u14_u1_n133, u2_u14_u1_n134, u2_u14_u1_n135, u2_u14_u1_n136, u2_u14_u1_n137, u2_u14_u1_n138, u2_u14_u1_n139, 
       u2_u14_u1_n140, u2_u14_u1_n141, u2_u14_u1_n142, u2_u14_u1_n143, u2_u14_u1_n144, u2_u14_u1_n145, u2_u14_u1_n146, u2_u14_u1_n147, u2_u14_u1_n148, 
       u2_u14_u1_n149, u2_u14_u1_n150, u2_u14_u1_n151, u2_u14_u1_n152, u2_u14_u1_n153, u2_u14_u1_n154, u2_u14_u1_n155, u2_u14_u1_n156, u2_u14_u1_n157, 
       u2_u14_u1_n158, u2_u14_u1_n159, u2_u14_u1_n160, u2_u14_u1_n161, u2_u14_u1_n162, u2_u14_u1_n163, u2_u14_u1_n164, u2_u14_u1_n165, u2_u14_u1_n166, 
       u2_u14_u1_n167, u2_u14_u1_n168, u2_u14_u1_n169, u2_u14_u1_n170, u2_u14_u1_n171, u2_u14_u1_n172, u2_u14_u1_n173, u2_u14_u1_n174, u2_u14_u1_n175, 
       u2_u14_u1_n176, u2_u14_u1_n177, u2_u14_u1_n178, u2_u14_u1_n179, u2_u14_u1_n180, u2_u14_u1_n181, u2_u14_u1_n182, u2_u14_u1_n183, u2_u14_u1_n184, 
       u2_u14_u1_n185, u2_u14_u1_n186, u2_u14_u1_n187, u2_u14_u1_n188, u2_u14_u1_n95, u2_u14_u1_n96, u2_u14_u1_n97, u2_u14_u1_n98, u2_u14_u1_n99, 
       u2_u14_u2_n100, u2_u14_u2_n101, u2_u14_u2_n102, u2_u14_u2_n103, u2_u14_u2_n104, u2_u14_u2_n105, u2_u14_u2_n106, u2_u14_u2_n107, u2_u14_u2_n108, 
       u2_u14_u2_n109, u2_u14_u2_n110, u2_u14_u2_n111, u2_u14_u2_n112, u2_u14_u2_n113, u2_u14_u2_n114, u2_u14_u2_n115, u2_u14_u2_n116, u2_u14_u2_n117, 
       u2_u14_u2_n118, u2_u14_u2_n119, u2_u14_u2_n120, u2_u14_u2_n121, u2_u14_u2_n122, u2_u14_u2_n123, u2_u14_u2_n124, u2_u14_u2_n125, u2_u14_u2_n126, 
       u2_u14_u2_n127, u2_u14_u2_n128, u2_u14_u2_n129, u2_u14_u2_n130, u2_u14_u2_n131, u2_u14_u2_n132, u2_u14_u2_n133, u2_u14_u2_n134, u2_u14_u2_n135, 
       u2_u14_u2_n136, u2_u14_u2_n137, u2_u14_u2_n138, u2_u14_u2_n139, u2_u14_u2_n140, u2_u14_u2_n141, u2_u14_u2_n142, u2_u14_u2_n143, u2_u14_u2_n144, 
       u2_u14_u2_n145, u2_u14_u2_n146, u2_u14_u2_n147, u2_u14_u2_n148, u2_u14_u2_n149, u2_u14_u2_n150, u2_u14_u2_n151, u2_u14_u2_n152, u2_u14_u2_n153, 
       u2_u14_u2_n154, u2_u14_u2_n155, u2_u14_u2_n156, u2_u14_u2_n157, u2_u14_u2_n158, u2_u14_u2_n159, u2_u14_u2_n160, u2_u14_u2_n161, u2_u14_u2_n162, 
       u2_u14_u2_n163, u2_u14_u2_n164, u2_u14_u2_n165, u2_u14_u2_n166, u2_u14_u2_n167, u2_u14_u2_n168, u2_u14_u2_n169, u2_u14_u2_n170, u2_u14_u2_n171, 
       u2_u14_u2_n172, u2_u14_u2_n173, u2_u14_u2_n174, u2_u14_u2_n175, u2_u14_u2_n176, u2_u14_u2_n177, u2_u14_u2_n178, u2_u14_u2_n179, u2_u14_u2_n180, 
       u2_u14_u2_n181, u2_u14_u2_n182, u2_u14_u2_n183, u2_u14_u2_n184, u2_u14_u2_n185, u2_u14_u2_n186, u2_u14_u2_n187, u2_u14_u2_n188, u2_u14_u2_n95, 
       u2_u14_u2_n96, u2_u14_u2_n97, u2_u14_u2_n98, u2_u14_u2_n99, u2_u14_u3_n100, u2_u14_u3_n101, u2_u14_u3_n102, u2_u14_u3_n103, u2_u14_u3_n104, 
       u2_u14_u3_n105, u2_u14_u3_n106, u2_u14_u3_n107, u2_u14_u3_n108, u2_u14_u3_n109, u2_u14_u3_n110, u2_u14_u3_n111, u2_u14_u3_n112, u2_u14_u3_n113, 
       u2_u14_u3_n114, u2_u14_u3_n115, u2_u14_u3_n116, u2_u14_u3_n117, u2_u14_u3_n118, u2_u14_u3_n119, u2_u14_u3_n120, u2_u14_u3_n121, u2_u14_u3_n122, 
       u2_u14_u3_n123, u2_u14_u3_n124, u2_u14_u3_n125, u2_u14_u3_n126, u2_u14_u3_n127, u2_u14_u3_n128, u2_u14_u3_n129, u2_u14_u3_n130, u2_u14_u3_n131, 
       u2_u14_u3_n132, u2_u14_u3_n133, u2_u14_u3_n134, u2_u14_u3_n135, u2_u14_u3_n136, u2_u14_u3_n137, u2_u14_u3_n138, u2_u14_u3_n139, u2_u14_u3_n140, 
       u2_u14_u3_n141, u2_u14_u3_n142, u2_u14_u3_n143, u2_u14_u3_n144, u2_u14_u3_n145, u2_u14_u3_n146, u2_u14_u3_n147, u2_u14_u3_n148, u2_u14_u3_n149, 
       u2_u14_u3_n150, u2_u14_u3_n151, u2_u14_u3_n152, u2_u14_u3_n153, u2_u14_u3_n154, u2_u14_u3_n155, u2_u14_u3_n156, u2_u14_u3_n157, u2_u14_u3_n158, 
       u2_u14_u3_n159, u2_u14_u3_n160, u2_u14_u3_n161, u2_u14_u3_n162, u2_u14_u3_n163, u2_u14_u3_n164, u2_u14_u3_n165, u2_u14_u3_n166, u2_u14_u3_n167, 
       u2_u14_u3_n168, u2_u14_u3_n169, u2_u14_u3_n170, u2_u14_u3_n171, u2_u14_u3_n172, u2_u14_u3_n173, u2_u14_u3_n174, u2_u14_u3_n175, u2_u14_u3_n176, 
       u2_u14_u3_n177, u2_u14_u3_n178, u2_u14_u3_n179, u2_u14_u3_n180, u2_u14_u3_n181, u2_u14_u3_n182, u2_u14_u3_n183, u2_u14_u3_n184, u2_u14_u3_n185, 
       u2_u14_u3_n186, u2_u14_u3_n94, u2_u14_u3_n95, u2_u14_u3_n96, u2_u14_u3_n97, u2_u14_u3_n98, u2_u14_u3_n99, u2_u15_X_1, u2_u15_X_10, 
       u2_u15_X_11, u2_u15_X_12, u2_u15_X_13, u2_u15_X_14, u2_u15_X_15, u2_u15_X_16, u2_u15_X_17, u2_u15_X_18, u2_u15_X_19, 
       u2_u15_X_2, u2_u15_X_20, u2_u15_X_21, u2_u15_X_22, u2_u15_X_23, u2_u15_X_24, u2_u15_X_3, u2_u15_X_4, u2_u15_X_5, 
       u2_u15_X_6, u2_u15_X_7, u2_u15_X_8, u2_u15_X_9, u2_u15_u0_n100, u2_u15_u0_n101, u2_u15_u0_n102, u2_u15_u0_n103, u2_u15_u0_n104, 
       u2_u15_u0_n105, u2_u15_u0_n106, u2_u15_u0_n107, u2_u15_u0_n108, u2_u15_u0_n109, u2_u15_u0_n110, u2_u15_u0_n111, u2_u15_u0_n112, u2_u15_u0_n113, 
       u2_u15_u0_n114, u2_u15_u0_n115, u2_u15_u0_n116, u2_u15_u0_n117, u2_u15_u0_n118, u2_u15_u0_n119, u2_u15_u0_n120, u2_u15_u0_n121, u2_u15_u0_n122, 
       u2_u15_u0_n123, u2_u15_u0_n124, u2_u15_u0_n125, u2_u15_u0_n126, u2_u15_u0_n127, u2_u15_u0_n128, u2_u15_u0_n129, u2_u15_u0_n130, u2_u15_u0_n131, 
       u2_u15_u0_n132, u2_u15_u0_n133, u2_u15_u0_n134, u2_u15_u0_n135, u2_u15_u0_n136, u2_u15_u0_n137, u2_u15_u0_n138, u2_u15_u0_n139, u2_u15_u0_n140, 
       u2_u15_u0_n141, u2_u15_u0_n142, u2_u15_u0_n143, u2_u15_u0_n144, u2_u15_u0_n145, u2_u15_u0_n146, u2_u15_u0_n147, u2_u15_u0_n148, u2_u15_u0_n149, 
       u2_u15_u0_n150, u2_u15_u0_n151, u2_u15_u0_n152, u2_u15_u0_n153, u2_u15_u0_n154, u2_u15_u0_n155, u2_u15_u0_n156, u2_u15_u0_n157, u2_u15_u0_n158, 
       u2_u15_u0_n159, u2_u15_u0_n160, u2_u15_u0_n161, u2_u15_u0_n162, u2_u15_u0_n163, u2_u15_u0_n164, u2_u15_u0_n165, u2_u15_u0_n166, u2_u15_u0_n167, 
       u2_u15_u0_n168, u2_u15_u0_n169, u2_u15_u0_n170, u2_u15_u0_n171, u2_u15_u0_n172, u2_u15_u0_n173, u2_u15_u0_n174, u2_u15_u0_n88, u2_u15_u0_n89, 
       u2_u15_u0_n90, u2_u15_u0_n91, u2_u15_u0_n92, u2_u15_u0_n93, u2_u15_u0_n94, u2_u15_u0_n95, u2_u15_u0_n96, u2_u15_u0_n97, u2_u15_u0_n98, 
       u2_u15_u0_n99, u2_u15_u1_n100, u2_u15_u1_n101, u2_u15_u1_n102, u2_u15_u1_n103, u2_u15_u1_n104, u2_u15_u1_n105, u2_u15_u1_n106, u2_u15_u1_n107, 
       u2_u15_u1_n108, u2_u15_u1_n109, u2_u15_u1_n110, u2_u15_u1_n111, u2_u15_u1_n112, u2_u15_u1_n113, u2_u15_u1_n114, u2_u15_u1_n115, u2_u15_u1_n116, 
       u2_u15_u1_n117, u2_u15_u1_n118, u2_u15_u1_n119, u2_u15_u1_n120, u2_u15_u1_n121, u2_u15_u1_n122, u2_u15_u1_n123, u2_u15_u1_n124, u2_u15_u1_n125, 
       u2_u15_u1_n126, u2_u15_u1_n127, u2_u15_u1_n128, u2_u15_u1_n129, u2_u15_u1_n130, u2_u15_u1_n131, u2_u15_u1_n132, u2_u15_u1_n133, u2_u15_u1_n134, 
       u2_u15_u1_n135, u2_u15_u1_n136, u2_u15_u1_n137, u2_u15_u1_n138, u2_u15_u1_n139, u2_u15_u1_n140, u2_u15_u1_n141, u2_u15_u1_n142, u2_u15_u1_n143, 
       u2_u15_u1_n144, u2_u15_u1_n145, u2_u15_u1_n146, u2_u15_u1_n147, u2_u15_u1_n148, u2_u15_u1_n149, u2_u15_u1_n150, u2_u15_u1_n151, u2_u15_u1_n152, 
       u2_u15_u1_n153, u2_u15_u1_n154, u2_u15_u1_n155, u2_u15_u1_n156, u2_u15_u1_n157, u2_u15_u1_n158, u2_u15_u1_n159, u2_u15_u1_n160, u2_u15_u1_n161, 
       u2_u15_u1_n162, u2_u15_u1_n163, u2_u15_u1_n164, u2_u15_u1_n165, u2_u15_u1_n166, u2_u15_u1_n167, u2_u15_u1_n168, u2_u15_u1_n169, u2_u15_u1_n170, 
       u2_u15_u1_n171, u2_u15_u1_n172, u2_u15_u1_n173, u2_u15_u1_n174, u2_u15_u1_n175, u2_u15_u1_n176, u2_u15_u1_n177, u2_u15_u1_n178, u2_u15_u1_n179, 
       u2_u15_u1_n180, u2_u15_u1_n181, u2_u15_u1_n182, u2_u15_u1_n183, u2_u15_u1_n184, u2_u15_u1_n185, u2_u15_u1_n186, u2_u15_u1_n187, u2_u15_u1_n188, 
       u2_u15_u1_n95, u2_u15_u1_n96, u2_u15_u1_n97, u2_u15_u1_n98, u2_u15_u1_n99, u2_u15_u2_n100, u2_u15_u2_n101, u2_u15_u2_n102, u2_u15_u2_n103, 
       u2_u15_u2_n104, u2_u15_u2_n105, u2_u15_u2_n106, u2_u15_u2_n107, u2_u15_u2_n108, u2_u15_u2_n109, u2_u15_u2_n110, u2_u15_u2_n111, u2_u15_u2_n112, 
       u2_u15_u2_n113, u2_u15_u2_n114, u2_u15_u2_n115, u2_u15_u2_n116, u2_u15_u2_n117, u2_u15_u2_n118, u2_u15_u2_n119, u2_u15_u2_n120, u2_u15_u2_n121, 
       u2_u15_u2_n122, u2_u15_u2_n123, u2_u15_u2_n124, u2_u15_u2_n125, u2_u15_u2_n126, u2_u15_u2_n127, u2_u15_u2_n128, u2_u15_u2_n129, u2_u15_u2_n130, 
       u2_u15_u2_n131, u2_u15_u2_n132, u2_u15_u2_n133, u2_u15_u2_n134, u2_u15_u2_n135, u2_u15_u2_n136, u2_u15_u2_n137, u2_u15_u2_n138, u2_u15_u2_n139, 
       u2_u15_u2_n140, u2_u15_u2_n141, u2_u15_u2_n142, u2_u15_u2_n143, u2_u15_u2_n144, u2_u15_u2_n145, u2_u15_u2_n146, u2_u15_u2_n147, u2_u15_u2_n148, 
       u2_u15_u2_n149, u2_u15_u2_n150, u2_u15_u2_n151, u2_u15_u2_n152, u2_u15_u2_n153, u2_u15_u2_n154, u2_u15_u2_n155, u2_u15_u2_n156, u2_u15_u2_n157, 
       u2_u15_u2_n158, u2_u15_u2_n159, u2_u15_u2_n160, u2_u15_u2_n161, u2_u15_u2_n162, u2_u15_u2_n163, u2_u15_u2_n164, u2_u15_u2_n165, u2_u15_u2_n166, 
       u2_u15_u2_n167, u2_u15_u2_n168, u2_u15_u2_n169, u2_u15_u2_n170, u2_u15_u2_n171, u2_u15_u2_n172, u2_u15_u2_n173, u2_u15_u2_n174, u2_u15_u2_n175, 
       u2_u15_u2_n176, u2_u15_u2_n177, u2_u15_u2_n178, u2_u15_u2_n179, u2_u15_u2_n180, u2_u15_u2_n181, u2_u15_u2_n182, u2_u15_u2_n183, u2_u15_u2_n184, 
       u2_u15_u2_n185, u2_u15_u2_n186, u2_u15_u2_n187, u2_u15_u2_n188, u2_u15_u2_n95, u2_u15_u2_n96, u2_u15_u2_n97, u2_u15_u2_n98, u2_u15_u2_n99, 
       u2_u15_u3_n100, u2_u15_u3_n101, u2_u15_u3_n102, u2_u15_u3_n103, u2_u15_u3_n104, u2_u15_u3_n105, u2_u15_u3_n106, u2_u15_u3_n107, u2_u15_u3_n108, 
       u2_u15_u3_n109, u2_u15_u3_n110, u2_u15_u3_n111, u2_u15_u3_n112, u2_u15_u3_n113, u2_u15_u3_n114, u2_u15_u3_n115, u2_u15_u3_n116, u2_u15_u3_n117, 
       u2_u15_u3_n118, u2_u15_u3_n119, u2_u15_u3_n120, u2_u15_u3_n121, u2_u15_u3_n122, u2_u15_u3_n123, u2_u15_u3_n124, u2_u15_u3_n125, u2_u15_u3_n126, 
       u2_u15_u3_n127, u2_u15_u3_n128, u2_u15_u3_n129, u2_u15_u3_n130, u2_u15_u3_n131, u2_u15_u3_n132, u2_u15_u3_n133, u2_u15_u3_n134, u2_u15_u3_n135, 
       u2_u15_u3_n136, u2_u15_u3_n137, u2_u15_u3_n138, u2_u15_u3_n139, u2_u15_u3_n140, u2_u15_u3_n141, u2_u15_u3_n142, u2_u15_u3_n143, u2_u15_u3_n144, 
       u2_u15_u3_n145, u2_u15_u3_n146, u2_u15_u3_n147, u2_u15_u3_n148, u2_u15_u3_n149, u2_u15_u3_n150, u2_u15_u3_n151, u2_u15_u3_n152, u2_u15_u3_n153, 
       u2_u15_u3_n154, u2_u15_u3_n155, u2_u15_u3_n156, u2_u15_u3_n157, u2_u15_u3_n158, u2_u15_u3_n159, u2_u15_u3_n160, u2_u15_u3_n161, u2_u15_u3_n162, 
       u2_u15_u3_n163, u2_u15_u3_n164, u2_u15_u3_n165, u2_u15_u3_n166, u2_u15_u3_n167, u2_u15_u3_n168, u2_u15_u3_n169, u2_u15_u3_n170, u2_u15_u3_n171, 
       u2_u15_u3_n172, u2_u15_u3_n173, u2_u15_u3_n174, u2_u15_u3_n175, u2_u15_u3_n176, u2_u15_u3_n177, u2_u15_u3_n178, u2_u15_u3_n179, u2_u15_u3_n180, 
       u2_u15_u3_n181, u2_u15_u3_n182, u2_u15_u3_n183, u2_u15_u3_n184, u2_u15_u3_n185, u2_u15_u3_n186, u2_u15_u3_n94, u2_u15_u3_n95, u2_u15_u3_n96, 
       u2_u15_u3_n97, u2_u15_u3_n98, u2_u15_u3_n99, u2_u1_X_1, u2_u1_X_10, u2_u1_X_11, u2_u1_X_12, u2_u1_X_2, u2_u1_X_3, 
       u2_u1_X_4, u2_u1_X_5, u2_u1_X_6, u2_u1_X_7, u2_u1_X_8, u2_u1_X_9, u2_u1_u0_n100, u2_u1_u0_n101, u2_u1_u0_n102, 
       u2_u1_u0_n103, u2_u1_u0_n104, u2_u1_u0_n105, u2_u1_u0_n106, u2_u1_u0_n107, u2_u1_u0_n108, u2_u1_u0_n109, u2_u1_u0_n110, u2_u1_u0_n111, 
       u2_u1_u0_n112, u2_u1_u0_n113, u2_u1_u0_n114, u2_u1_u0_n115, u2_u1_u0_n116, u2_u1_u0_n117, u2_u1_u0_n118, u2_u1_u0_n119, u2_u1_u0_n120, 
       u2_u1_u0_n121, u2_u1_u0_n122, u2_u1_u0_n123, u2_u1_u0_n124, u2_u1_u0_n125, u2_u1_u0_n126, u2_u1_u0_n127, u2_u1_u0_n128, u2_u1_u0_n129, 
       u2_u1_u0_n130, u2_u1_u0_n131, u2_u1_u0_n132, u2_u1_u0_n133, u2_u1_u0_n134, u2_u1_u0_n135, u2_u1_u0_n136, u2_u1_u0_n137, u2_u1_u0_n138, 
       u2_u1_u0_n139, u2_u1_u0_n140, u2_u1_u0_n141, u2_u1_u0_n142, u2_u1_u0_n143, u2_u1_u0_n144, u2_u1_u0_n145, u2_u1_u0_n146, u2_u1_u0_n147, 
       u2_u1_u0_n148, u2_u1_u0_n149, u2_u1_u0_n150, u2_u1_u0_n151, u2_u1_u0_n152, u2_u1_u0_n153, u2_u1_u0_n154, u2_u1_u0_n155, u2_u1_u0_n156, 
       u2_u1_u0_n157, u2_u1_u0_n158, u2_u1_u0_n159, u2_u1_u0_n160, u2_u1_u0_n161, u2_u1_u0_n162, u2_u1_u0_n163, u2_u1_u0_n164, u2_u1_u0_n165, 
       u2_u1_u0_n166, u2_u1_u0_n167, u2_u1_u0_n168, u2_u1_u0_n169, u2_u1_u0_n170, u2_u1_u0_n171, u2_u1_u0_n172, u2_u1_u0_n173, u2_u1_u0_n174, 
       u2_u1_u0_n88, u2_u1_u0_n89, u2_u1_u0_n90, u2_u1_u0_n91, u2_u1_u0_n92, u2_u1_u0_n93, u2_u1_u0_n94, u2_u1_u0_n95, u2_u1_u0_n96, 
       u2_u1_u0_n97, u2_u1_u0_n98, u2_u1_u0_n99, u2_u1_u1_n100, u2_u1_u1_n101, u2_u1_u1_n102, u2_u1_u1_n103, u2_u1_u1_n104, u2_u1_u1_n105, 
       u2_u1_u1_n106, u2_u1_u1_n107, u2_u1_u1_n108, u2_u1_u1_n109, u2_u1_u1_n110, u2_u1_u1_n111, u2_u1_u1_n112, u2_u1_u1_n113, u2_u1_u1_n114, 
       u2_u1_u1_n115, u2_u1_u1_n116, u2_u1_u1_n117, u2_u1_u1_n118, u2_u1_u1_n119, u2_u1_u1_n120, u2_u1_u1_n121, u2_u1_u1_n122, u2_u1_u1_n123, 
       u2_u1_u1_n124, u2_u1_u1_n125, u2_u1_u1_n126, u2_u1_u1_n127, u2_u1_u1_n128, u2_u1_u1_n129, u2_u1_u1_n130, u2_u1_u1_n131, u2_u1_u1_n132, 
       u2_u1_u1_n133, u2_u1_u1_n134, u2_u1_u1_n135, u2_u1_u1_n136, u2_u1_u1_n137, u2_u1_u1_n138, u2_u1_u1_n139, u2_u1_u1_n140, u2_u1_u1_n141, 
       u2_u1_u1_n142, u2_u1_u1_n143, u2_u1_u1_n144, u2_u1_u1_n145, u2_u1_u1_n146, u2_u1_u1_n147, u2_u1_u1_n148, u2_u1_u1_n149, u2_u1_u1_n150, 
       u2_u1_u1_n151, u2_u1_u1_n152, u2_u1_u1_n153, u2_u1_u1_n154, u2_u1_u1_n155, u2_u1_u1_n156, u2_u1_u1_n157, u2_u1_u1_n158, u2_u1_u1_n159, 
       u2_u1_u1_n160, u2_u1_u1_n161, u2_u1_u1_n162, u2_u1_u1_n163, u2_u1_u1_n164, u2_u1_u1_n165, u2_u1_u1_n166, u2_u1_u1_n167, u2_u1_u1_n168, 
       u2_u1_u1_n169, u2_u1_u1_n170, u2_u1_u1_n171, u2_u1_u1_n172, u2_u1_u1_n173, u2_u1_u1_n174, u2_u1_u1_n175, u2_u1_u1_n176, u2_u1_u1_n177, 
       u2_u1_u1_n178, u2_u1_u1_n179, u2_u1_u1_n180, u2_u1_u1_n181, u2_u1_u1_n182, u2_u1_u1_n183, u2_u1_u1_n184, u2_u1_u1_n185, u2_u1_u1_n186, 
       u2_u1_u1_n187, u2_u1_u1_n188, u2_u1_u1_n95, u2_u1_u1_n96, u2_u1_u1_n97, u2_u1_u1_n98, u2_u1_u1_n99, u2_u5_X_13, u2_u5_X_14, 
       u2_u5_X_15, u2_u5_X_16, u2_u5_X_17, u2_u5_X_18, u2_u5_X_19, u2_u5_X_20, u2_u5_X_21, u2_u5_X_22, u2_u5_X_23, 
       u2_u5_X_24, u2_u5_X_31, u2_u5_X_32, u2_u5_X_33, u2_u5_X_34, u2_u5_X_35, u2_u5_X_36, u2_u5_X_37, u2_u5_X_38, 
       u2_u5_X_39, u2_u5_X_40, u2_u5_X_41, u2_u5_X_42, u2_u5_u2_n100, u2_u5_u2_n101, u2_u5_u2_n102, u2_u5_u2_n103, u2_u5_u2_n104, 
       u2_u5_u2_n105, u2_u5_u2_n106, u2_u5_u2_n107, u2_u5_u2_n108, u2_u5_u2_n109, u2_u5_u2_n110, u2_u5_u2_n111, u2_u5_u2_n112, u2_u5_u2_n113, 
       u2_u5_u2_n114, u2_u5_u2_n115, u2_u5_u2_n116, u2_u5_u2_n117, u2_u5_u2_n118, u2_u5_u2_n119, u2_u5_u2_n120, u2_u5_u2_n121, u2_u5_u2_n122, 
       u2_u5_u2_n123, u2_u5_u2_n124, u2_u5_u2_n125, u2_u5_u2_n126, u2_u5_u2_n127, u2_u5_u2_n128, u2_u5_u2_n129, u2_u5_u2_n130, u2_u5_u2_n131, 
       u2_u5_u2_n132, u2_u5_u2_n133, u2_u5_u2_n134, u2_u5_u2_n135, u2_u5_u2_n136, u2_u5_u2_n137, u2_u5_u2_n138, u2_u5_u2_n139, u2_u5_u2_n140, 
       u2_u5_u2_n141, u2_u5_u2_n142, u2_u5_u2_n143, u2_u5_u2_n144, u2_u5_u2_n145, u2_u5_u2_n146, u2_u5_u2_n147, u2_u5_u2_n148, u2_u5_u2_n149, 
       u2_u5_u2_n150, u2_u5_u2_n151, u2_u5_u2_n152, u2_u5_u2_n153, u2_u5_u2_n154, u2_u5_u2_n155, u2_u5_u2_n156, u2_u5_u2_n157, u2_u5_u2_n158, 
       u2_u5_u2_n159, u2_u5_u2_n160, u2_u5_u2_n161, u2_u5_u2_n162, u2_u5_u2_n163, u2_u5_u2_n164, u2_u5_u2_n165, u2_u5_u2_n166, u2_u5_u2_n167, 
       u2_u5_u2_n168, u2_u5_u2_n169, u2_u5_u2_n170, u2_u5_u2_n171, u2_u5_u2_n172, u2_u5_u2_n173, u2_u5_u2_n174, u2_u5_u2_n175, u2_u5_u2_n176, 
       u2_u5_u2_n177, u2_u5_u2_n178, u2_u5_u2_n179, u2_u5_u2_n180, u2_u5_u2_n181, u2_u5_u2_n182, u2_u5_u2_n183, u2_u5_u2_n184, u2_u5_u2_n185, 
       u2_u5_u2_n186, u2_u5_u2_n187, u2_u5_u2_n188, u2_u5_u2_n95, u2_u5_u2_n96, u2_u5_u2_n97, u2_u5_u2_n98, u2_u5_u2_n99, u2_u5_u3_n100, 
       u2_u5_u3_n101, u2_u5_u3_n102, u2_u5_u3_n103, u2_u5_u3_n104, u2_u5_u3_n105, u2_u5_u3_n106, u2_u5_u3_n107, u2_u5_u3_n108, u2_u5_u3_n109, 
       u2_u5_u3_n110, u2_u5_u3_n111, u2_u5_u3_n112, u2_u5_u3_n113, u2_u5_u3_n114, u2_u5_u3_n115, u2_u5_u3_n116, u2_u5_u3_n117, u2_u5_u3_n118, 
       u2_u5_u3_n119, u2_u5_u3_n120, u2_u5_u3_n121, u2_u5_u3_n122, u2_u5_u3_n123, u2_u5_u3_n124, u2_u5_u3_n125, u2_u5_u3_n126, u2_u5_u3_n127, 
       u2_u5_u3_n128, u2_u5_u3_n129, u2_u5_u3_n130, u2_u5_u3_n131, u2_u5_u3_n132, u2_u5_u3_n133, u2_u5_u3_n134, u2_u5_u3_n135, u2_u5_u3_n136, 
       u2_u5_u3_n137, u2_u5_u3_n138, u2_u5_u3_n139, u2_u5_u3_n140, u2_u5_u3_n141, u2_u5_u3_n142, u2_u5_u3_n143, u2_u5_u3_n144, u2_u5_u3_n145, 
       u2_u5_u3_n146, u2_u5_u3_n147, u2_u5_u3_n148, u2_u5_u3_n149, u2_u5_u3_n150, u2_u5_u3_n151, u2_u5_u3_n152, u2_u5_u3_n153, u2_u5_u3_n154, 
       u2_u5_u3_n155, u2_u5_u3_n156, u2_u5_u3_n157, u2_u5_u3_n158, u2_u5_u3_n159, u2_u5_u3_n160, u2_u5_u3_n161, u2_u5_u3_n162, u2_u5_u3_n163, 
       u2_u5_u3_n164, u2_u5_u3_n165, u2_u5_u3_n166, u2_u5_u3_n167, u2_u5_u3_n168, u2_u5_u3_n169, u2_u5_u3_n170, u2_u5_u3_n171, u2_u5_u3_n172, 
       u2_u5_u3_n173, u2_u5_u3_n174, u2_u5_u3_n175, u2_u5_u3_n176, u2_u5_u3_n177, u2_u5_u3_n178, u2_u5_u3_n179, u2_u5_u3_n180, u2_u5_u3_n181, 
       u2_u5_u3_n182, u2_u5_u3_n183, u2_u5_u3_n184, u2_u5_u3_n185, u2_u5_u3_n186, u2_u5_u3_n94, u2_u5_u3_n95, u2_u5_u3_n96, u2_u5_u3_n97, 
       u2_u5_u3_n98, u2_u5_u3_n99, u2_u5_u5_n100, u2_u5_u5_n101, u2_u5_u5_n102, u2_u5_u5_n103, u2_u5_u5_n104, u2_u5_u5_n105, u2_u5_u5_n106, 
       u2_u5_u5_n107, u2_u5_u5_n108, u2_u5_u5_n109, u2_u5_u5_n110, u2_u5_u5_n111, u2_u5_u5_n112, u2_u5_u5_n113, u2_u5_u5_n114, u2_u5_u5_n115, 
       u2_u5_u5_n116, u2_u5_u5_n117, u2_u5_u5_n118, u2_u5_u5_n119, u2_u5_u5_n120, u2_u5_u5_n121, u2_u5_u5_n122, u2_u5_u5_n123, u2_u5_u5_n124, 
       u2_u5_u5_n125, u2_u5_u5_n126, u2_u5_u5_n127, u2_u5_u5_n128, u2_u5_u5_n129, u2_u5_u5_n130, u2_u5_u5_n131, u2_u5_u5_n132, u2_u5_u5_n133, 
       u2_u5_u5_n134, u2_u5_u5_n135, u2_u5_u5_n136, u2_u5_u5_n137, u2_u5_u5_n138, u2_u5_u5_n139, u2_u5_u5_n140, u2_u5_u5_n141, u2_u5_u5_n142, 
       u2_u5_u5_n143, u2_u5_u5_n144, u2_u5_u5_n145, u2_u5_u5_n146, u2_u5_u5_n147, u2_u5_u5_n148, u2_u5_u5_n149, u2_u5_u5_n150, u2_u5_u5_n151, 
       u2_u5_u5_n152, u2_u5_u5_n153, u2_u5_u5_n154, u2_u5_u5_n155, u2_u5_u5_n156, u2_u5_u5_n157, u2_u5_u5_n158, u2_u5_u5_n159, u2_u5_u5_n160, 
       u2_u5_u5_n161, u2_u5_u5_n162, u2_u5_u5_n163, u2_u5_u5_n164, u2_u5_u5_n165, u2_u5_u5_n166, u2_u5_u5_n167, u2_u5_u5_n168, u2_u5_u5_n169, 
       u2_u5_u5_n170, u2_u5_u5_n171, u2_u5_u5_n172, u2_u5_u5_n173, u2_u5_u5_n174, u2_u5_u5_n175, u2_u5_u5_n176, u2_u5_u5_n177, u2_u5_u5_n178, 
       u2_u5_u5_n179, u2_u5_u5_n180, u2_u5_u5_n181, u2_u5_u5_n182, u2_u5_u5_n183, u2_u5_u5_n184, u2_u5_u5_n185, u2_u5_u5_n186, u2_u5_u5_n187, 
       u2_u5_u5_n188, u2_u5_u5_n189, u2_u5_u5_n190, u2_u5_u5_n191, u2_u5_u5_n192, u2_u5_u5_n193, u2_u5_u5_n194, u2_u5_u5_n195, u2_u5_u5_n196, 
       u2_u5_u5_n99, u2_u5_u6_n100, u2_u5_u6_n101, u2_u5_u6_n102, u2_u5_u6_n103, u2_u5_u6_n104, u2_u5_u6_n105, u2_u5_u6_n106, u2_u5_u6_n107, 
       u2_u5_u6_n108, u2_u5_u6_n109, u2_u5_u6_n110, u2_u5_u6_n111, u2_u5_u6_n112, u2_u5_u6_n113, u2_u5_u6_n114, u2_u5_u6_n115, u2_u5_u6_n116, 
       u2_u5_u6_n117, u2_u5_u6_n118, u2_u5_u6_n119, u2_u5_u6_n120, u2_u5_u6_n121, u2_u5_u6_n122, u2_u5_u6_n123, u2_u5_u6_n124, u2_u5_u6_n125, 
       u2_u5_u6_n126, u2_u5_u6_n127, u2_u5_u6_n128, u2_u5_u6_n129, u2_u5_u6_n130, u2_u5_u6_n131, u2_u5_u6_n132, u2_u5_u6_n133, u2_u5_u6_n134, 
       u2_u5_u6_n135, u2_u5_u6_n136, u2_u5_u6_n137, u2_u5_u6_n138, u2_u5_u6_n139, u2_u5_u6_n140, u2_u5_u6_n141, u2_u5_u6_n142, u2_u5_u6_n143, 
       u2_u5_u6_n144, u2_u5_u6_n145, u2_u5_u6_n146, u2_u5_u6_n147, u2_u5_u6_n148, u2_u5_u6_n149, u2_u5_u6_n150, u2_u5_u6_n151, u2_u5_u6_n152, 
       u2_u5_u6_n153, u2_u5_u6_n154, u2_u5_u6_n155, u2_u5_u6_n156, u2_u5_u6_n157, u2_u5_u6_n158, u2_u5_u6_n159, u2_u5_u6_n160, u2_u5_u6_n161, 
       u2_u5_u6_n162, u2_u5_u6_n163, u2_u5_u6_n164, u2_u5_u6_n165, u2_u5_u6_n166, u2_u5_u6_n167, u2_u5_u6_n168, u2_u5_u6_n169, u2_u5_u6_n170, 
       u2_u5_u6_n171, u2_u5_u6_n172, u2_u5_u6_n173, u2_u5_u6_n174, u2_u5_u6_n88, u2_u5_u6_n89, u2_u5_u6_n90, u2_u5_u6_n91, u2_u5_u6_n92, 
       u2_u5_u6_n93, u2_u5_u6_n94, u2_u5_u6_n95, u2_u5_u6_n96, u2_u5_u6_n97, u2_u5_u6_n98, u2_u5_u6_n99, u2_u6_X_1, u2_u6_X_10, 
       u2_u6_X_11, u2_u6_X_12, u2_u6_X_13, u2_u6_X_14, u2_u6_X_15, u2_u6_X_16, u2_u6_X_17, u2_u6_X_18, u2_u6_X_2, 
       u2_u6_X_3, u2_u6_X_4, u2_u6_X_5, u2_u6_X_6, u2_u6_X_7, u2_u6_X_8, u2_u6_X_9, u2_u6_u0_n100, u2_u6_u0_n101, 
       u2_u6_u0_n102, u2_u6_u0_n103, u2_u6_u0_n104, u2_u6_u0_n105, u2_u6_u0_n106, u2_u6_u0_n107, u2_u6_u0_n108, u2_u6_u0_n109, u2_u6_u0_n110, 
       u2_u6_u0_n111, u2_u6_u0_n112, u2_u6_u0_n113, u2_u6_u0_n114, u2_u6_u0_n115, u2_u6_u0_n116, u2_u6_u0_n117, u2_u6_u0_n118, u2_u6_u0_n119, 
       u2_u6_u0_n120, u2_u6_u0_n121, u2_u6_u0_n122, u2_u6_u0_n123, u2_u6_u0_n124, u2_u6_u0_n125, u2_u6_u0_n126, u2_u6_u0_n127, u2_u6_u0_n128, 
       u2_u6_u0_n129, u2_u6_u0_n130, u2_u6_u0_n131, u2_u6_u0_n132, u2_u6_u0_n133, u2_u6_u0_n134, u2_u6_u0_n135, u2_u6_u0_n136, u2_u6_u0_n137, 
       u2_u6_u0_n138, u2_u6_u0_n139, u2_u6_u0_n140, u2_u6_u0_n141, u2_u6_u0_n142, u2_u6_u0_n143, u2_u6_u0_n144, u2_u6_u0_n145, u2_u6_u0_n146, 
       u2_u6_u0_n147, u2_u6_u0_n148, u2_u6_u0_n149, u2_u6_u0_n150, u2_u6_u0_n151, u2_u6_u0_n152, u2_u6_u0_n153, u2_u6_u0_n154, u2_u6_u0_n155, 
       u2_u6_u0_n156, u2_u6_u0_n157, u2_u6_u0_n158, u2_u6_u0_n159, u2_u6_u0_n160, u2_u6_u0_n161, u2_u6_u0_n162, u2_u6_u0_n163, u2_u6_u0_n164, 
       u2_u6_u0_n165, u2_u6_u0_n166, u2_u6_u0_n167, u2_u6_u0_n168, u2_u6_u0_n169, u2_u6_u0_n170, u2_u6_u0_n171, u2_u6_u0_n172, u2_u6_u0_n173, 
       u2_u6_u0_n174, u2_u6_u0_n88, u2_u6_u0_n89, u2_u6_u0_n90, u2_u6_u0_n91, u2_u6_u0_n92, u2_u6_u0_n93, u2_u6_u0_n94, u2_u6_u0_n95, 
       u2_u6_u0_n96, u2_u6_u0_n97, u2_u6_u0_n98, u2_u6_u0_n99, u2_u6_u1_n100, u2_u6_u1_n101, u2_u6_u1_n102, u2_u6_u1_n103, u2_u6_u1_n104, 
       u2_u6_u1_n105, u2_u6_u1_n106, u2_u6_u1_n107, u2_u6_u1_n108, u2_u6_u1_n109, u2_u6_u1_n110, u2_u6_u1_n111, u2_u6_u1_n112, u2_u6_u1_n113, 
       u2_u6_u1_n114, u2_u6_u1_n115, u2_u6_u1_n116, u2_u6_u1_n117, u2_u6_u1_n118, u2_u6_u1_n119, u2_u6_u1_n120, u2_u6_u1_n121, u2_u6_u1_n122, 
       u2_u6_u1_n123, u2_u6_u1_n124, u2_u6_u1_n125, u2_u6_u1_n126, u2_u6_u1_n127, u2_u6_u1_n128, u2_u6_u1_n129, u2_u6_u1_n130, u2_u6_u1_n131, 
       u2_u6_u1_n132, u2_u6_u1_n133, u2_u6_u1_n134, u2_u6_u1_n135, u2_u6_u1_n136, u2_u6_u1_n137, u2_u6_u1_n138, u2_u6_u1_n139, u2_u6_u1_n140, 
       u2_u6_u1_n141, u2_u6_u1_n142, u2_u6_u1_n143, u2_u6_u1_n144, u2_u6_u1_n145, u2_u6_u1_n146, u2_u6_u1_n147, u2_u6_u1_n148, u2_u6_u1_n149, 
       u2_u6_u1_n150, u2_u6_u1_n151, u2_u6_u1_n152, u2_u6_u1_n153, u2_u6_u1_n154, u2_u6_u1_n155, u2_u6_u1_n156, u2_u6_u1_n157, u2_u6_u1_n158, 
       u2_u6_u1_n159, u2_u6_u1_n160, u2_u6_u1_n161, u2_u6_u1_n162, u2_u6_u1_n163, u2_u6_u1_n164, u2_u6_u1_n165, u2_u6_u1_n166, u2_u6_u1_n167, 
       u2_u6_u1_n168, u2_u6_u1_n169, u2_u6_u1_n170, u2_u6_u1_n171, u2_u6_u1_n172, u2_u6_u1_n173, u2_u6_u1_n174, u2_u6_u1_n175, u2_u6_u1_n176, 
       u2_u6_u1_n177, u2_u6_u1_n178, u2_u6_u1_n179, u2_u6_u1_n180, u2_u6_u1_n181, u2_u6_u1_n182, u2_u6_u1_n183, u2_u6_u1_n184, u2_u6_u1_n185, 
       u2_u6_u1_n186, u2_u6_u1_n187, u2_u6_u1_n188, u2_u6_u1_n95, u2_u6_u1_n96, u2_u6_u1_n97, u2_u6_u1_n98, u2_u6_u1_n99, u2_u6_u2_n100, 
       u2_u6_u2_n101, u2_u6_u2_n102, u2_u6_u2_n103, u2_u6_u2_n104, u2_u6_u2_n105, u2_u6_u2_n106, u2_u6_u2_n107, u2_u6_u2_n108, u2_u6_u2_n109, 
       u2_u6_u2_n110, u2_u6_u2_n111, u2_u6_u2_n112, u2_u6_u2_n113, u2_u6_u2_n114, u2_u6_u2_n115, u2_u6_u2_n116, u2_u6_u2_n117, u2_u6_u2_n118, 
       u2_u6_u2_n119, u2_u6_u2_n120, u2_u6_u2_n121, u2_u6_u2_n122, u2_u6_u2_n123, u2_u6_u2_n124, u2_u6_u2_n125, u2_u6_u2_n126, u2_u6_u2_n127, 
       u2_u6_u2_n128, u2_u6_u2_n129, u2_u6_u2_n130, u2_u6_u2_n131, u2_u6_u2_n132, u2_u6_u2_n133, u2_u6_u2_n134, u2_u6_u2_n135, u2_u6_u2_n136, 
       u2_u6_u2_n137, u2_u6_u2_n138, u2_u6_u2_n139, u2_u6_u2_n140, u2_u6_u2_n141, u2_u6_u2_n142, u2_u6_u2_n143, u2_u6_u2_n144, u2_u6_u2_n145, 
       u2_u6_u2_n146, u2_u6_u2_n147, u2_u6_u2_n148, u2_u6_u2_n149, u2_u6_u2_n150, u2_u6_u2_n151, u2_u6_u2_n152, u2_u6_u2_n153, u2_u6_u2_n154, 
       u2_u6_u2_n155, u2_u6_u2_n156, u2_u6_u2_n157, u2_u6_u2_n158, u2_u6_u2_n159, u2_u6_u2_n160, u2_u6_u2_n161, u2_u6_u2_n162, u2_u6_u2_n163, 
       u2_u6_u2_n164, u2_u6_u2_n165, u2_u6_u2_n166, u2_u6_u2_n167, u2_u6_u2_n168, u2_u6_u2_n169, u2_u6_u2_n170, u2_u6_u2_n171, u2_u6_u2_n172, 
       u2_u6_u2_n173, u2_u6_u2_n174, u2_u6_u2_n175, u2_u6_u2_n176, u2_u6_u2_n177, u2_u6_u2_n178, u2_u6_u2_n179, u2_u6_u2_n180, u2_u6_u2_n181, 
       u2_u6_u2_n182, u2_u6_u2_n183, u2_u6_u2_n184, u2_u6_u2_n185, u2_u6_u2_n186, u2_u6_u2_n187, u2_u6_u2_n188, u2_u6_u2_n95, u2_u6_u2_n96, 
       u2_u6_u2_n97, u2_u6_u2_n98, u2_u6_u2_n99, u2_u9_X_10, u2_u9_X_11, u2_u9_X_12, u2_u9_X_13, u2_u9_X_14, u2_u9_X_15, 
       u2_u9_X_16, u2_u9_X_17, u2_u9_X_18, u2_u9_X_7, u2_u9_X_8, u2_u9_X_9, u2_u9_u1_n100, u2_u9_u1_n101, u2_u9_u1_n102, 
       u2_u9_u1_n103, u2_u9_u1_n104, u2_u9_u1_n105, u2_u9_u1_n106, u2_u9_u1_n107, u2_u9_u1_n108, u2_u9_u1_n109, u2_u9_u1_n110, u2_u9_u1_n111, 
       u2_u9_u1_n112, u2_u9_u1_n113, u2_u9_u1_n114, u2_u9_u1_n115, u2_u9_u1_n116, u2_u9_u1_n117, u2_u9_u1_n118, u2_u9_u1_n119, u2_u9_u1_n120, 
       u2_u9_u1_n121, u2_u9_u1_n122, u2_u9_u1_n123, u2_u9_u1_n124, u2_u9_u1_n125, u2_u9_u1_n126, u2_u9_u1_n127, u2_u9_u1_n128, u2_u9_u1_n129, 
       u2_u9_u1_n130, u2_u9_u1_n131, u2_u9_u1_n132, u2_u9_u1_n133, u2_u9_u1_n134, u2_u9_u1_n135, u2_u9_u1_n136, u2_u9_u1_n137, u2_u9_u1_n138, 
       u2_u9_u1_n139, u2_u9_u1_n140, u2_u9_u1_n141, u2_u9_u1_n142, u2_u9_u1_n143, u2_u9_u1_n144, u2_u9_u1_n145, u2_u9_u1_n146, u2_u9_u1_n147, 
       u2_u9_u1_n148, u2_u9_u1_n149, u2_u9_u1_n150, u2_u9_u1_n151, u2_u9_u1_n152, u2_u9_u1_n153, u2_u9_u1_n154, u2_u9_u1_n155, u2_u9_u1_n156, 
       u2_u9_u1_n157, u2_u9_u1_n158, u2_u9_u1_n159, u2_u9_u1_n160, u2_u9_u1_n161, u2_u9_u1_n162, u2_u9_u1_n163, u2_u9_u1_n164, u2_u9_u1_n165, 
       u2_u9_u1_n166, u2_u9_u1_n167, u2_u9_u1_n168, u2_u9_u1_n169, u2_u9_u1_n170, u2_u9_u1_n171, u2_u9_u1_n172, u2_u9_u1_n173, u2_u9_u1_n174, 
       u2_u9_u1_n175, u2_u9_u1_n176, u2_u9_u1_n177, u2_u9_u1_n178, u2_u9_u1_n179, u2_u9_u1_n180, u2_u9_u1_n181, u2_u9_u1_n182, u2_u9_u1_n183, 
       u2_u9_u1_n184, u2_u9_u1_n185, u2_u9_u1_n186, u2_u9_u1_n187, u2_u9_u1_n188, u2_u9_u1_n95, u2_u9_u1_n96, u2_u9_u1_n97, u2_u9_u1_n98, 
       u2_u9_u1_n99, u2_u9_u2_n100, u2_u9_u2_n101, u2_u9_u2_n102, u2_u9_u2_n103, u2_u9_u2_n104, u2_u9_u2_n105, u2_u9_u2_n106, u2_u9_u2_n107, 
       u2_u9_u2_n108, u2_u9_u2_n109, u2_u9_u2_n110, u2_u9_u2_n111, u2_u9_u2_n112, u2_u9_u2_n113, u2_u9_u2_n114, u2_u9_u2_n115, u2_u9_u2_n116, 
       u2_u9_u2_n117, u2_u9_u2_n118, u2_u9_u2_n119, u2_u9_u2_n120, u2_u9_u2_n121, u2_u9_u2_n122, u2_u9_u2_n123, u2_u9_u2_n124, u2_u9_u2_n125, 
       u2_u9_u2_n126, u2_u9_u2_n127, u2_u9_u2_n128, u2_u9_u2_n129, u2_u9_u2_n130, u2_u9_u2_n131, u2_u9_u2_n132, u2_u9_u2_n133, u2_u9_u2_n134, 
       u2_u9_u2_n135, u2_u9_u2_n136, u2_u9_u2_n137, u2_u9_u2_n138, u2_u9_u2_n139, u2_u9_u2_n140, u2_u9_u2_n141, u2_u9_u2_n142, u2_u9_u2_n143, 
       u2_u9_u2_n144, u2_u9_u2_n145, u2_u9_u2_n146, u2_u9_u2_n147, u2_u9_u2_n148, u2_u9_u2_n149, u2_u9_u2_n150, u2_u9_u2_n151, u2_u9_u2_n152, 
       u2_u9_u2_n153, u2_u9_u2_n154, u2_u9_u2_n155, u2_u9_u2_n156, u2_u9_u2_n157, u2_u9_u2_n158, u2_u9_u2_n159, u2_u9_u2_n160, u2_u9_u2_n161, 
       u2_u9_u2_n162, u2_u9_u2_n163, u2_u9_u2_n164, u2_u9_u2_n165, u2_u9_u2_n166, u2_u9_u2_n167, u2_u9_u2_n168, u2_u9_u2_n169, u2_u9_u2_n170, 
       u2_u9_u2_n171, u2_u9_u2_n172, u2_u9_u2_n173, u2_u9_u2_n174, u2_u9_u2_n175, u2_u9_u2_n176, u2_u9_u2_n177, u2_u9_u2_n178, u2_u9_u2_n179, 
       u2_u9_u2_n180, u2_u9_u2_n181, u2_u9_u2_n182, u2_u9_u2_n183, u2_u9_u2_n184, u2_u9_u2_n185, u2_u9_u2_n186, u2_u9_u2_n187, u2_u9_u2_n188, 
       u2_u9_u2_n95, u2_u9_u2_n96, u2_u9_u2_n97, u2_u9_u2_n98, u2_u9_u2_n99, u2_uk_n1004, u2_uk_n1005, u2_uk_n1059, u2_uk_n1060, 
       u2_uk_n1062, u2_uk_n1068, u2_uk_n1075, u2_uk_n1076, u2_uk_n1078, u2_uk_n1086, u2_uk_n1095, u2_uk_n1153, u2_uk_n1154, 
       u2_uk_n1159, u2_uk_n1160, u2_uk_n1175, u2_uk_n1184, u2_uk_n242, u2_uk_n250, u2_uk_n308, u2_uk_n375, u2_uk_n382, 
       u2_uk_n460, u2_uk_n496, u2_uk_n501, u2_uk_n509, u2_uk_n934, u2_uk_n935, u2_uk_n936, u2_uk_n937, u2_uk_n946, 
       u2_uk_n949, u2_uk_n950, u2_uk_n951, u2_uk_n952, u2_uk_n953, u2_uk_n965, u2_uk_n966, u2_uk_n968, u2_uk_n969, 
       u2_uk_n971, u2_uk_n978, u2_uk_n990, u2_uk_n991,  u2_uk_n992;
  XOR2_X1 u0_U103 (.B( u0_L0_13 ) , .Z( u0_N44 ) , .A( u0_out1_13 ) );
  XOR2_X1 u0_U11 (.B( u0_L1_28 ) , .Z( u0_N91 ) , .A( u0_out2_28 ) );
  XOR2_X1 u0_U114 (.B( u0_L0_12 ) , .Z( u0_N43 ) , .A( u0_out1_12 ) );
  XOR2_X1 u0_U125 (.B( u0_L0_11 ) , .Z( u0_N42 ) , .A( u0_out1_11 ) );
  XOR2_X1 u0_U132 (.B( u0_L11_30 ) , .Z( u0_N413 ) , .A( u0_out12_30 ) );
  XOR2_X1 u0_U134 (.B( u0_L11_28 ) , .Z( u0_N411 ) , .A( u0_out12_28 ) );
  XOR2_X1 u0_U137 (.B( u0_L11_26 ) , .Z( u0_N409 ) , .A( u0_out12_26 ) );
  XOR2_X1 u0_U139 (.B( u0_L11_24 ) , .Z( u0_N407 ) , .A( u0_out12_24 ) );
  XOR2_X1 u0_U14 (.B( u0_L1_26 ) , .Z( u0_N89 ) , .A( u0_out2_26 ) );
  XOR2_X1 u0_U143 (.B( u0_L11_20 ) , .Z( u0_N403 ) , .A( u0_out12_20 ) );
  XOR2_X1 u0_U145 (.B( u0_L11_18 ) , .Z( u0_N401 ) , .A( u0_out12_18 ) );
  XOR2_X1 u0_U147 (.B( u0_L0_9 ) , .Z( u0_N40 ) , .A( u0_out1_9 ) );
  XOR2_X1 u0_U149 (.B( u0_L11_16 ) , .Z( u0_N399 ) , .A( u0_out12_16 ) );
  XOR2_X1 u0_U152 (.B( u0_L11_13 ) , .Z( u0_N396 ) , .A( u0_out12_13 ) );
  XOR2_X1 u0_U155 (.B( u0_L11_10 ) , .Z( u0_N393 ) , .A( u0_out12_10 ) );
  XOR2_X1 u0_U159 (.B( u0_L0_8 ) , .Z( u0_N39 ) , .A( u0_out1_8 ) );
  XOR2_X1 u0_U16 (.B( u0_L1_24 ) , .Z( u0_N87 ) , .A( u0_out2_24 ) );
  XOR2_X1 u0_U160 (.B( u0_L11_6 ) , .Z( u0_N389 ) , .A( u0_out12_6 ) );
  XOR2_X1 u0_U164 (.B( u0_L11_2 ) , .Z( u0_N385 ) , .A( u0_out12_2 ) );
  XOR2_X1 u0_U165 (.B( u0_L11_1 ) , .Z( u0_N384 ) , .A( u0_out12_1 ) );
  XOR2_X1 u0_U17 (.B( u0_L1_23 ) , .Z( u0_N86 ) , .A( u0_out2_23 ) );
  XOR2_X1 u0_U170 (.B( u0_L0_7 ) , .Z( u0_N38 ) , .A( u0_out1_7 ) );
  XOR2_X1 u0_U20 (.B( u0_L1_20 ) , .Z( u0_N83 ) , .A( u0_out2_20 ) );
  XOR2_X1 u0_U201 (.B( u0_L9_32 ) , .Z( u0_N351 ) , .A( u0_out10_32 ) );
  XOR2_X1 u0_U203 (.B( u0_L0_4 ) , .Z( u0_N35 ) , .A( u0_out1_4 ) );
  XOR2_X1 u0_U204 (.B( u0_L9_30 ) , .Z( u0_N349 ) , .A( u0_out10_30 ) );
  XOR2_X1 u0_U205 (.B( u0_L9_29 ) , .Z( u0_N348 ) , .A( u0_out10_29 ) );
  XOR2_X1 u0_U206 (.B( u0_L9_28 ) , .Z( u0_N347 ) , .A( u0_out10_28 ) );
  XOR2_X1 u0_U207 (.B( u0_L9_27 ) , .Z( u0_N346 ) , .A( u0_out10_27 ) );
  XOR2_X1 u0_U208 (.B( u0_L9_26 ) , .Z( u0_N345 ) , .A( u0_out10_26 ) );
  XOR2_X1 u0_U210 (.B( u0_L9_24 ) , .Z( u0_N343 ) , .A( u0_out10_24 ) );
  XOR2_X1 u0_U212 (.B( u0_L9_22 ) , .Z( u0_N341 ) , .A( u0_out10_22 ) );
  XOR2_X1 u0_U213 (.B( u0_L9_21 ) , .Z( u0_N340 ) , .A( u0_out10_21 ) );
  XOR2_X1 u0_U214 (.B( u0_L0_3 ) , .Z( u0_N34 ) , .A( u0_out1_3 ) );
  XOR2_X1 u0_U215 (.B( u0_L9_20 ) , .Z( u0_N339 ) , .A( u0_out10_20 ) );
  XOR2_X1 u0_U216 (.B( u0_L9_19 ) , .Z( u0_N338 ) , .A( u0_out10_19 ) );
  XOR2_X1 u0_U217 (.B( u0_L9_18 ) , .Z( u0_N337 ) , .A( u0_out10_18 ) );
  XOR2_X1 u0_U219 (.B( u0_L9_16 ) , .Z( u0_N335 ) , .A( u0_out10_16 ) );
  XOR2_X1 u0_U22 (.B( u0_L1_18 ) , .Z( u0_N81 ) , .A( u0_out2_18 ) );
  XOR2_X1 u0_U220 (.B( u0_L9_15 ) , .Z( u0_N334 ) , .A( u0_out10_15 ) );
  XOR2_X1 u0_U222 (.B( u0_L9_13 ) , .Z( u0_N332 ) , .A( u0_out10_13 ) );
  XOR2_X1 u0_U223 (.B( u0_L9_12 ) , .Z( u0_N331 ) , .A( u0_out10_12 ) );
  XOR2_X1 u0_U224 (.B( u0_L9_11 ) , .Z( u0_N330 ) , .A( u0_out10_11 ) );
  XOR2_X1 u0_U225 (.B( u0_L0_2 ) , .Z( u0_N33 ) , .A( u0_out1_2 ) );
  XOR2_X1 u0_U226 (.B( u0_L9_10 ) , .Z( u0_N329 ) , .A( u0_out10_10 ) );
  XOR2_X1 u0_U229 (.B( u0_L9_7 ) , .Z( u0_N326 ) , .A( u0_out10_7 ) );
  XOR2_X1 u0_U23 (.B( u0_L1_17 ) , .Z( u0_N80 ) , .A( u0_out2_17 ) );
  XOR2_X1 u0_U230 (.B( u0_L9_6 ) , .Z( u0_N325 ) , .A( u0_out10_6 ) );
  XOR2_X1 u0_U231 (.B( u0_L9_5 ) , .Z( u0_N324 ) , .A( u0_out10_5 ) );
  XOR2_X1 u0_U232 (.B( u0_L9_4 ) , .Z( u0_N323 ) , .A( u0_out10_4 ) );
  XOR2_X1 u0_U234 (.B( u0_L9_2 ) , .Z( u0_N321 ) , .A( u0_out10_2 ) );
  XOR2_X1 u0_U235 (.B( u0_L9_1 ) , .Z( u0_N320 ) , .A( u0_out10_1 ) );
  XOR2_X1 u0_U243 (.B( u0_L8_26 ) , .Z( u0_N313 ) , .A( u0_out9_26 ) );
  XOR2_X1 u0_U25 (.B( u0_L1_16 ) , .Z( u0_N79 ) , .A( u0_out2_16 ) );
  XOR2_X1 u0_U250 (.B( u0_L8_20 ) , .Z( u0_N307 ) , .A( u0_out9_20 ) );
  XOR2_X1 u0_U262 (.B( u0_L8_10 ) , .Z( u0_N297 ) , .A( u0_out9_10 ) );
  XOR2_X1 u0_U272 (.B( u0_L8_1 ) , .Z( u0_N288 ) , .A( u0_out9_1 ) );
  XOR2_X1 u0_U28 (.B( u0_L1_13 ) , .Z( u0_N76 ) , .A( u0_out2_13 ) );
  XOR2_X1 u0_U3 (.B( u0_L2_4 ) , .Z( u0_N99 ) , .A( u0_out3_4 ) );
  XOR2_X1 u0_U31 (.B( u0_L1_10 ) , .Z( u0_N73 ) , .A( u0_out2_10 ) );
  XOR2_X1 u0_U313 (.B( u0_L6_27 ) , .Z( u0_N250 ) , .A( u0_out7_27 ) );
  XOR2_X1 u0_U32 (.B( u0_L1_9 ) , .Z( u0_N72 ) , .A( u0_out2_9 ) );
  XOR2_X1 u0_U320 (.B( u0_L6_21 ) , .Z( u0_N244 ) , .A( u0_out7_21 ) );
  XOR2_X1 u0_U327 (.B( u0_L6_15 ) , .Z( u0_N238 ) , .A( u0_out7_15 ) );
  XOR2_X1 u0_U338 (.B( u0_L6_5 ) , .Z( u0_N228 ) , .A( u0_out7_5 ) );
  XOR2_X1 u0_U344 (.B( u0_L5_31 ) , .Z( u0_N222 ) , .A( u0_out6_31 ) );
  XOR2_X1 u0_U345 (.B( u0_L5_30 ) , .Z( u0_N221 ) , .A( u0_out6_30 ) );
  XOR2_X1 u0_U348 (.B( u0_L5_28 ) , .Z( u0_N219 ) , .A( u0_out6_28 ) );
  XOR2_X1 u0_U349 (.B( u0_L5_27 ) , .Z( u0_N218 ) , .A( u0_out6_27 ) );
  XOR2_X1 u0_U350 (.B( u0_L5_26 ) , .Z( u0_N217 ) , .A( u0_out6_26 ) );
  XOR2_X1 u0_U352 (.B( u0_L5_24 ) , .Z( u0_N215 ) , .A( u0_out6_24 ) );
  XOR2_X1 u0_U353 (.B( u0_L5_23 ) , .Z( u0_N214 ) , .A( u0_out6_23 ) );
  XOR2_X1 u0_U355 (.B( u0_L5_21 ) , .Z( u0_N212 ) , .A( u0_out6_21 ) );
  XOR2_X1 u0_U356 (.B( u0_L5_20 ) , .Z( u0_N211 ) , .A( u0_out6_20 ) );
  XOR2_X1 u0_U359 (.B( u0_L5_18 ) , .Z( u0_N209 ) , .A( u0_out6_18 ) );
  XOR2_X1 u0_U36 (.B( u0_L1_6 ) , .Z( u0_N69 ) , .A( u0_out2_6 ) );
  XOR2_X1 u0_U360 (.B( u0_L5_17 ) , .Z( u0_N208 ) , .A( u0_out6_17 ) );
  XOR2_X1 u0_U361 (.B( u0_L5_16 ) , .Z( u0_N207 ) , .A( u0_out6_16 ) );
  XOR2_X1 u0_U362 (.B( u0_L5_15 ) , .Z( u0_N206 ) , .A( u0_out6_15 ) );
  XOR2_X1 u0_U364 (.B( u0_L5_13 ) , .Z( u0_N204 ) , .A( u0_out6_13 ) );
  XOR2_X1 u0_U367 (.B( u0_L5_10 ) , .Z( u0_N201 ) , .A( u0_out6_10 ) );
  XOR2_X1 u0_U368 (.B( u0_L5_9 ) , .Z( u0_N200 ) , .A( u0_out6_9 ) );
  XOR2_X1 u0_U373 (.B( u0_L5_6 ) , .Z( u0_N197 ) , .A( u0_out6_6 ) );
  XOR2_X1 u0_U374 (.B( u0_L5_5 ) , .Z( u0_N196 ) , .A( u0_out6_5 ) );
  XOR2_X1 u0_U377 (.B( u0_L5_2 ) , .Z( u0_N193 ) , .A( u0_out6_2 ) );
  XOR2_X1 u0_U378 (.B( u0_L5_1 ) , .Z( u0_N192 ) , .A( u0_out6_1 ) );
  XOR2_X1 u0_U379 (.B( u0_L4_32 ) , .Z( u0_N191 ) , .A( u0_out5_32 ) );
  XOR2_X1 u0_U383 (.B( u0_L4_29 ) , .Z( u0_N188 ) , .A( u0_out5_29 ) );
  XOR2_X1 u0_U386 (.B( u0_L4_26 ) , .Z( u0_N185 ) , .A( u0_out5_26 ) );
  XOR2_X1 u0_U387 (.B( u0_L4_25 ) , .Z( u0_N184 ) , .A( u0_out5_25 ) );
  XOR2_X1 u0_U390 (.B( u0_L4_22 ) , .Z( u0_N181 ) , .A( u0_out5_22 ) );
  XOR2_X1 u0_U393 (.B( u0_L4_20 ) , .Z( u0_N179 ) , .A( u0_out5_20 ) );
  XOR2_X1 u0_U394 (.B( u0_L4_19 ) , .Z( u0_N178 ) , .A( u0_out5_19 ) );
  XOR2_X1 u0_U399 (.B( u0_L4_14 ) , .Z( u0_N173 ) , .A( u0_out5_14 ) );
  XOR2_X1 u0_U4 (.B( u0_L2_3 ) , .Z( u0_N98 ) , .A( u0_out3_3 ) );
  XOR2_X1 u0_U40 (.B( u0_L1_2 ) , .Z( u0_N65 ) , .A( u0_out2_2 ) );
  XOR2_X1 u0_U401 (.B( u0_L4_12 ) , .Z( u0_N171 ) , .A( u0_out5_12 ) );
  XOR2_X1 u0_U402 (.B( u0_L4_11 ) , .Z( u0_N170 ) , .A( u0_out5_11 ) );
  XOR2_X1 u0_U404 (.B( u0_L4_10 ) , .Z( u0_N169 ) , .A( u0_out5_10 ) );
  XOR2_X1 u0_U406 (.B( u0_L4_8 ) , .Z( u0_N167 ) , .A( u0_out5_8 ) );
  XOR2_X1 u0_U407 (.B( u0_L4_7 ) , .Z( u0_N166 ) , .A( u0_out5_7 ) );
  XOR2_X1 u0_U41 (.B( u0_L1_1 ) , .Z( u0_N64 ) , .A( u0_out2_1 ) );
  XOR2_X1 u0_U410 (.B( u0_L4_4 ) , .Z( u0_N163 ) , .A( u0_out5_4 ) );
  XOR2_X1 u0_U411 (.B( u0_L4_3 ) , .Z( u0_N162 ) , .A( u0_out5_3 ) );
  XOR2_X1 u0_U413 (.B( u0_L4_1 ) , .Z( u0_N160 ) , .A( u0_out5_1 ) );
  XOR2_X1 u0_U42 (.B( u0_L0_32 ) , .Z( u0_N63 ) , .A( u0_out1_32 ) );
  XOR2_X1 u0_U43 (.B( u0_L0_31 ) , .Z( u0_N62 ) , .A( u0_out1_31 ) );
  XOR2_X1 u0_U45 (.B( u0_L0_29 ) , .Z( u0_N60 ) , .A( u0_out1_29 ) );
  XOR2_X1 u0_U451 (.B( u0_L2_31 ) , .Z( u0_N126 ) , .A( u0_out3_31 ) );
  XOR2_X1 u0_U452 (.B( u0_L2_30 ) , .Z( u0_N125 ) , .A( u0_out3_30 ) );
  XOR2_X1 u0_U453 (.B( u0_L2_29 ) , .Z( u0_N124 ) , .A( u0_out3_29 ) );
  XOR2_X1 u0_U454 (.B( u0_L2_28 ) , .Z( u0_N123 ) , .A( u0_out3_28 ) );
  XOR2_X1 u0_U456 (.B( u0_L2_26 ) , .Z( u0_N121 ) , .A( u0_out3_26 ) );
  XOR2_X1 u0_U457 (.B( u0_L2_25 ) , .Z( u0_N120 ) , .A( u0_out3_25 ) );
  XOR2_X1 u0_U459 (.B( u0_L2_24 ) , .Z( u0_N119 ) , .A( u0_out3_24 ) );
  XOR2_X1 u0_U460 (.B( u0_L2_23 ) , .Z( u0_N118 ) , .A( u0_out3_23 ) );
  XOR2_X1 u0_U463 (.B( u0_L2_20 ) , .Z( u0_N115 ) , .A( u0_out3_20 ) );
  XOR2_X1 u0_U464 (.B( u0_L2_19 ) , .Z( u0_N114 ) , .A( u0_out3_19 ) );
  XOR2_X1 u0_U465 (.B( u0_L2_18 ) , .Z( u0_N113 ) , .A( u0_out3_18 ) );
  XOR2_X1 u0_U466 (.B( u0_L2_17 ) , .Z( u0_N112 ) , .A( u0_out3_17 ) );
  XOR2_X1 u0_U467 (.B( u0_L2_16 ) , .Z( u0_N111 ) , .A( u0_out3_16 ) );
  XOR2_X1 u0_U47 (.B( u0_L0_28 ) , .Z( u0_N59 ) , .A( u0_out1_28 ) );
  XOR2_X1 u0_U470 (.B( u0_L2_14 ) , .Z( u0_N109 ) , .A( u0_out3_14 ) );
  XOR2_X1 u0_U471 (.B( u0_L2_13 ) , .Z( u0_N108 ) , .A( u0_out3_13 ) );
  XOR2_X1 u0_U473 (.B( u0_L2_11 ) , .Z( u0_N106 ) , .A( u0_out3_11 ) );
  XOR2_X1 u0_U474 (.B( u0_L2_10 ) , .Z( u0_N105 ) , .A( u0_out3_10 ) );
  XOR2_X1 u0_U475 (.B( u0_L2_9 ) , .Z( u0_N104 ) , .A( u0_out3_9 ) );
  XOR2_X1 u0_U476 (.B( u0_L2_8 ) , .Z( u0_N103 ) , .A( u0_out3_8 ) );
  XOR2_X1 u0_U478 (.B( u0_L2_6 ) , .Z( u0_N101 ) , .A( u0_out3_6 ) );
  XOR2_X1 u0_U5 (.B( u0_L2_2 ) , .Z( u0_N97 ) , .A( u0_out3_2 ) );
  XOR2_X1 u0_U50 (.B( u0_L0_25 ) , .Z( u0_N56 ) , .A( u0_out1_25 ) );
  XOR2_X1 u0_U52 (.B( u0_L0_23 ) , .Z( u0_N54 ) , .A( u0_out1_23 ) );
  XOR2_X1 u0_U53 (.B( u0_L0_22 ) , .Z( u0_N53 ) , .A( u0_out1_22 ) );
  XOR2_X1 u0_U56 (.B( u0_L0_19 ) , .Z( u0_N50 ) , .A( u0_out1_19 ) );
  XOR2_X1 u0_U58 (.B( u0_L0_18 ) , .Z( u0_N49 ) , .A( u0_out1_18 ) );
  XOR2_X1 u0_U59 (.B( u0_L0_17 ) , .Z( u0_N48 ) , .A( u0_out1_17 ) );
  XOR2_X1 u0_U6 (.B( u0_L2_1 ) , .Z( u0_N96 ) , .A( u0_out3_1 ) );
  XOR2_X1 u0_U67 (.B( u0_L13_25 ) , .Z( u0_N472 ) , .A( u0_out14_25 ) );
  XOR2_X1 u0_U79 (.B( u0_L13_14 ) , .Z( u0_N461 ) , .A( u0_out14_14 ) );
  XOR2_X1 u0_U8 (.B( u0_L1_31 ) , .Z( u0_N94 ) , .A( u0_out2_31 ) );
  XOR2_X1 u0_U86 (.B( u0_L13_8 ) , .Z( u0_N455 ) , .A( u0_out14_8 ) );
  XOR2_X1 u0_U9 (.B( u0_L1_30 ) , .Z( u0_N93 ) , .A( u0_out2_30 ) );
  XOR2_X1 u0_U91 (.B( u0_L13_3 ) , .Z( u0_N450 ) , .A( u0_out14_3 ) );
  XOR2_X1 u0_U92 (.B( u0_L0_14 ) , .Z( u0_N45 ) , .A( u0_out1_14 ) );
  XOR2_X1 u0_u10_U1 (.B( u0_K11_9 ) , .A( u0_R9_6 ) , .Z( u0_u10_X_9 ) );
  XOR2_X1 u0_u10_U10 (.B( u0_K11_45 ) , .A( u0_R9_30 ) , .Z( u0_u10_X_45 ) );
  XOR2_X1 u0_u10_U11 (.B( u0_K11_44 ) , .A( u0_R9_29 ) , .Z( u0_u10_X_44 ) );
  XOR2_X1 u0_u10_U12 (.B( u0_K11_43 ) , .A( u0_R9_28 ) , .Z( u0_u10_X_43 ) );
  XOR2_X1 u0_u10_U13 (.B( u0_K11_42 ) , .A( u0_R9_29 ) , .Z( u0_u10_X_42 ) );
  XOR2_X1 u0_u10_U14 (.B( u0_K11_41 ) , .A( u0_R9_28 ) , .Z( u0_u10_X_41 ) );
  XOR2_X1 u0_u10_U15 (.B( u0_K11_40 ) , .A( u0_R9_27 ) , .Z( u0_u10_X_40 ) );
  XOR2_X1 u0_u10_U17 (.B( u0_K11_39 ) , .A( u0_R9_26 ) , .Z( u0_u10_X_39 ) );
  XOR2_X1 u0_u10_U18 (.B( u0_K11_38 ) , .A( u0_R9_25 ) , .Z( u0_u10_X_38 ) );
  XOR2_X1 u0_u10_U19 (.B( u0_K11_37 ) , .A( u0_R9_24 ) , .Z( u0_u10_X_37 ) );
  XOR2_X1 u0_u10_U2 (.B( u0_K11_8 ) , .A( u0_R9_5 ) , .Z( u0_u10_X_8 ) );
  XOR2_X1 u0_u10_U20 (.B( u0_K11_36 ) , .A( u0_R9_25 ) , .Z( u0_u10_X_36 ) );
  XOR2_X1 u0_u10_U21 (.B( u0_K11_35 ) , .A( u0_R9_24 ) , .Z( u0_u10_X_35 ) );
  XOR2_X1 u0_u10_U22 (.B( u0_K11_34 ) , .A( u0_R9_23 ) , .Z( u0_u10_X_34 ) );
  XOR2_X1 u0_u10_U23 (.B( u0_K11_33 ) , .A( u0_R9_22 ) , .Z( u0_u10_X_33 ) );
  XOR2_X1 u0_u10_U24 (.B( u0_K11_32 ) , .A( u0_R9_21 ) , .Z( u0_u10_X_32 ) );
  XOR2_X1 u0_u10_U25 (.B( u0_K11_31 ) , .A( u0_R9_20 ) , .Z( u0_u10_X_31 ) );
  XOR2_X1 u0_u10_U3 (.B( u0_K11_7 ) , .A( u0_R9_4 ) , .Z( u0_u10_X_7 ) );
  XOR2_X1 u0_u10_U33 (.B( u0_K11_24 ) , .A( u0_R9_17 ) , .Z( u0_u10_X_24 ) );
  XOR2_X1 u0_u10_U34 (.B( u0_K11_23 ) , .A( u0_R9_16 ) , .Z( u0_u10_X_23 ) );
  XOR2_X1 u0_u10_U35 (.B( u0_K11_22 ) , .A( u0_R9_15 ) , .Z( u0_u10_X_22 ) );
  XOR2_X1 u0_u10_U36 (.B( u0_K11_21 ) , .A( u0_R9_14 ) , .Z( u0_u10_X_21 ) );
  XOR2_X1 u0_u10_U37 (.B( u0_K11_20 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_20 ) );
  XOR2_X1 u0_u10_U39 (.B( u0_K11_19 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_19 ) );
  XOR2_X1 u0_u10_U40 (.B( u0_K11_18 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_18 ) );
  XOR2_X1 u0_u10_U41 (.B( u0_K11_17 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_17 ) );
  XOR2_X1 u0_u10_U42 (.B( u0_K11_16 ) , .A( u0_R9_11 ) , .Z( u0_u10_X_16 ) );
  XOR2_X1 u0_u10_U43 (.B( u0_K11_15 ) , .A( u0_R9_10 ) , .Z( u0_u10_X_15 ) );
  XOR2_X1 u0_u10_U44 (.B( u0_K11_14 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_14 ) );
  XOR2_X1 u0_u10_U45 (.B( u0_K11_13 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_13 ) );
  XOR2_X1 u0_u10_U46 (.B( u0_K11_12 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_12 ) );
  XOR2_X1 u0_u10_U47 (.B( u0_K11_11 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_11 ) );
  XOR2_X1 u0_u10_U48 (.B( u0_K11_10 ) , .A( u0_R9_7 ) , .Z( u0_u10_X_10 ) );
  XOR2_X1 u0_u10_U7 (.B( u0_K11_48 ) , .A( u0_R9_1 ) , .Z( u0_u10_X_48 ) );
  XOR2_X1 u0_u10_U8 (.B( u0_K11_47 ) , .A( u0_R9_32 ) , .Z( u0_u10_X_47 ) );
  XOR2_X1 u0_u10_U9 (.B( u0_K11_46 ) , .A( u0_R9_31 ) , .Z( u0_u10_X_46 ) );
  AOI21_X1 u0_u10_u1_U10 (.B2( u0_u10_u1_n155 ) , .B1( u0_u10_u1_n156 ) , .ZN( u0_u10_u1_n157 ) , .A( u0_u10_u1_n174 ) );
  NAND3_X1 u0_u10_u1_U100 (.ZN( u0_u10_u1_n113 ) , .A1( u0_u10_u1_n120 ) , .A3( u0_u10_u1_n133 ) , .A2( u0_u10_u1_n155 ) );
  NAND2_X1 u0_u10_u1_U11 (.ZN( u0_u10_u1_n140 ) , .A2( u0_u10_u1_n150 ) , .A1( u0_u10_u1_n155 ) );
  NAND2_X1 u0_u10_u1_U12 (.A1( u0_u10_u1_n131 ) , .ZN( u0_u10_u1_n147 ) , .A2( u0_u10_u1_n153 ) );
  AOI22_X1 u0_u10_u1_U13 (.B2( u0_u10_u1_n136 ) , .A2( u0_u10_u1_n137 ) , .ZN( u0_u10_u1_n143 ) , .A1( u0_u10_u1_n171 ) , .B1( u0_u10_u1_n173 ) );
  INV_X1 u0_u10_u1_U14 (.A( u0_u10_u1_n147 ) , .ZN( u0_u10_u1_n181 ) );
  INV_X1 u0_u10_u1_U15 (.A( u0_u10_u1_n139 ) , .ZN( u0_u10_u1_n174 ) );
  OR4_X1 u0_u10_u1_U16 (.A4( u0_u10_u1_n106 ) , .A3( u0_u10_u1_n107 ) , .ZN( u0_u10_u1_n108 ) , .A1( u0_u10_u1_n117 ) , .A2( u0_u10_u1_n184 ) );
  AOI21_X1 u0_u10_u1_U17 (.ZN( u0_u10_u1_n106 ) , .A( u0_u10_u1_n112 ) , .B1( u0_u10_u1_n154 ) , .B2( u0_u10_u1_n156 ) );
  AOI21_X1 u0_u10_u1_U18 (.ZN( u0_u10_u1_n107 ) , .B1( u0_u10_u1_n134 ) , .B2( u0_u10_u1_n149 ) , .A( u0_u10_u1_n174 ) );
  INV_X1 u0_u10_u1_U19 (.A( u0_u10_u1_n101 ) , .ZN( u0_u10_u1_n184 ) );
  INV_X1 u0_u10_u1_U20 (.A( u0_u10_u1_n112 ) , .ZN( u0_u10_u1_n171 ) );
  NAND2_X1 u0_u10_u1_U21 (.ZN( u0_u10_u1_n141 ) , .A1( u0_u10_u1_n153 ) , .A2( u0_u10_u1_n156 ) );
  AND2_X1 u0_u10_u1_U22 (.A1( u0_u10_u1_n123 ) , .ZN( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n161 ) );
  NAND2_X1 u0_u10_u1_U23 (.A2( u0_u10_u1_n115 ) , .A1( u0_u10_u1_n116 ) , .ZN( u0_u10_u1_n148 ) );
  NAND2_X1 u0_u10_u1_U24 (.A2( u0_u10_u1_n133 ) , .A1( u0_u10_u1_n135 ) , .ZN( u0_u10_u1_n159 ) );
  NAND2_X1 u0_u10_u1_U25 (.A2( u0_u10_u1_n115 ) , .A1( u0_u10_u1_n120 ) , .ZN( u0_u10_u1_n132 ) );
  INV_X1 u0_u10_u1_U26 (.A( u0_u10_u1_n154 ) , .ZN( u0_u10_u1_n178 ) );
  INV_X1 u0_u10_u1_U27 (.A( u0_u10_u1_n151 ) , .ZN( u0_u10_u1_n183 ) );
  AND2_X1 u0_u10_u1_U28 (.A1( u0_u10_u1_n129 ) , .A2( u0_u10_u1_n133 ) , .ZN( u0_u10_u1_n149 ) );
  INV_X1 u0_u10_u1_U29 (.A( u0_u10_u1_n131 ) , .ZN( u0_u10_u1_n180 ) );
  INV_X1 u0_u10_u1_U3 (.A( u0_u10_u1_n159 ) , .ZN( u0_u10_u1_n182 ) );
  OAI221_X1 u0_u10_u1_U30 (.A( u0_u10_u1_n119 ) , .C2( u0_u10_u1_n129 ) , .ZN( u0_u10_u1_n138 ) , .B2( u0_u10_u1_n152 ) , .C1( u0_u10_u1_n174 ) , .B1( u0_u10_u1_n187 ) );
  INV_X1 u0_u10_u1_U31 (.A( u0_u10_u1_n148 ) , .ZN( u0_u10_u1_n187 ) );
  AOI211_X1 u0_u10_u1_U32 (.B( u0_u10_u1_n117 ) , .A( u0_u10_u1_n118 ) , .ZN( u0_u10_u1_n119 ) , .C2( u0_u10_u1_n146 ) , .C1( u0_u10_u1_n159 ) );
  NOR2_X1 u0_u10_u1_U33 (.A1( u0_u10_u1_n168 ) , .A2( u0_u10_u1_n176 ) , .ZN( u0_u10_u1_n98 ) );
  OAI21_X1 u0_u10_u1_U34 (.B2( u0_u10_u1_n123 ) , .ZN( u0_u10_u1_n145 ) , .B1( u0_u10_u1_n160 ) , .A( u0_u10_u1_n185 ) );
  INV_X1 u0_u10_u1_U35 (.A( u0_u10_u1_n122 ) , .ZN( u0_u10_u1_n185 ) );
  AOI21_X1 u0_u10_u1_U36 (.B2( u0_u10_u1_n120 ) , .B1( u0_u10_u1_n121 ) , .ZN( u0_u10_u1_n122 ) , .A( u0_u10_u1_n128 ) );
  NAND2_X1 u0_u10_u1_U37 (.A1( u0_u10_u1_n128 ) , .ZN( u0_u10_u1_n146 ) , .A2( u0_u10_u1_n160 ) );
  NAND2_X1 u0_u10_u1_U38 (.A2( u0_u10_u1_n112 ) , .ZN( u0_u10_u1_n139 ) , .A1( u0_u10_u1_n152 ) );
  NAND2_X1 u0_u10_u1_U39 (.A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n156 ) , .A2( u0_u10_u1_n99 ) );
  AOI221_X1 u0_u10_u1_U4 (.A( u0_u10_u1_n138 ) , .C2( u0_u10_u1_n139 ) , .C1( u0_u10_u1_n140 ) , .B2( u0_u10_u1_n141 ) , .ZN( u0_u10_u1_n142 ) , .B1( u0_u10_u1_n175 ) );
  AOI221_X1 u0_u10_u1_U40 (.B1( u0_u10_u1_n140 ) , .ZN( u0_u10_u1_n167 ) , .B2( u0_u10_u1_n172 ) , .C2( u0_u10_u1_n175 ) , .C1( u0_u10_u1_n178 ) , .A( u0_u10_u1_n188 ) );
  INV_X1 u0_u10_u1_U41 (.ZN( u0_u10_u1_n188 ) , .A( u0_u10_u1_n97 ) );
  AOI211_X1 u0_u10_u1_U42 (.A( u0_u10_u1_n118 ) , .C1( u0_u10_u1_n132 ) , .C2( u0_u10_u1_n139 ) , .B( u0_u10_u1_n96 ) , .ZN( u0_u10_u1_n97 ) );
  AOI21_X1 u0_u10_u1_U43 (.B2( u0_u10_u1_n121 ) , .B1( u0_u10_u1_n135 ) , .A( u0_u10_u1_n152 ) , .ZN( u0_u10_u1_n96 ) );
  NOR2_X1 u0_u10_u1_U44 (.ZN( u0_u10_u1_n117 ) , .A1( u0_u10_u1_n121 ) , .A2( u0_u10_u1_n160 ) );
  AOI21_X1 u0_u10_u1_U45 (.A( u0_u10_u1_n128 ) , .B2( u0_u10_u1_n129 ) , .ZN( u0_u10_u1_n130 ) , .B1( u0_u10_u1_n150 ) );
  NAND2_X1 u0_u10_u1_U46 (.ZN( u0_u10_u1_n112 ) , .A1( u0_u10_u1_n169 ) , .A2( u0_u10_u1_n170 ) );
  NAND2_X1 u0_u10_u1_U47 (.ZN( u0_u10_u1_n129 ) , .A2( u0_u10_u1_n95 ) , .A1( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U48 (.A1( u0_u10_u1_n102 ) , .ZN( u0_u10_u1_n154 ) , .A2( u0_u10_u1_n99 ) );
  NAND2_X1 u0_u10_u1_U49 (.A2( u0_u10_u1_n100 ) , .ZN( u0_u10_u1_n135 ) , .A1( u0_u10_u1_n99 ) );
  AOI211_X1 u0_u10_u1_U5 (.ZN( u0_u10_u1_n124 ) , .A( u0_u10_u1_n138 ) , .C2( u0_u10_u1_n139 ) , .B( u0_u10_u1_n145 ) , .C1( u0_u10_u1_n147 ) );
  AOI21_X1 u0_u10_u1_U50 (.A( u0_u10_u1_n152 ) , .B2( u0_u10_u1_n153 ) , .B1( u0_u10_u1_n154 ) , .ZN( u0_u10_u1_n158 ) );
  INV_X1 u0_u10_u1_U51 (.A( u0_u10_u1_n160 ) , .ZN( u0_u10_u1_n175 ) );
  NAND2_X1 u0_u10_u1_U52 (.A1( u0_u10_u1_n100 ) , .ZN( u0_u10_u1_n116 ) , .A2( u0_u10_u1_n95 ) );
  NAND2_X1 u0_u10_u1_U53 (.A1( u0_u10_u1_n102 ) , .ZN( u0_u10_u1_n131 ) , .A2( u0_u10_u1_n95 ) );
  NAND2_X1 u0_u10_u1_U54 (.A2( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n121 ) , .A1( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U55 (.A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n153 ) , .A2( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U56 (.A2( u0_u10_u1_n104 ) , .A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n133 ) );
  NAND2_X1 u0_u10_u1_U57 (.ZN( u0_u10_u1_n150 ) , .A2( u0_u10_u1_n98 ) , .A1( u0_u10_u1_n99 ) );
  NAND2_X1 u0_u10_u1_U58 (.A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n155 ) , .A2( u0_u10_u1_n95 ) );
  OAI21_X1 u0_u10_u1_U59 (.ZN( u0_u10_u1_n109 ) , .B1( u0_u10_u1_n129 ) , .B2( u0_u10_u1_n160 ) , .A( u0_u10_u1_n167 ) );
  AOI22_X1 u0_u10_u1_U6 (.B2( u0_u10_u1_n113 ) , .A2( u0_u10_u1_n114 ) , .ZN( u0_u10_u1_n125 ) , .A1( u0_u10_u1_n171 ) , .B1( u0_u10_u1_n173 ) );
  NAND2_X1 u0_u10_u1_U60 (.A2( u0_u10_u1_n100 ) , .A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n120 ) );
  NAND2_X1 u0_u10_u1_U61 (.A1( u0_u10_u1_n102 ) , .A2( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n115 ) );
  NAND2_X1 u0_u10_u1_U62 (.A2( u0_u10_u1_n100 ) , .A1( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n151 ) );
  NAND2_X1 u0_u10_u1_U63 (.A2( u0_u10_u1_n103 ) , .A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n161 ) );
  INV_X1 u0_u10_u1_U64 (.A( u0_u10_u1_n152 ) , .ZN( u0_u10_u1_n173 ) );
  INV_X1 u0_u10_u1_U65 (.A( u0_u10_u1_n128 ) , .ZN( u0_u10_u1_n172 ) );
  NAND2_X1 u0_u10_u1_U66 (.A2( u0_u10_u1_n102 ) , .A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n123 ) );
  AOI211_X1 u0_u10_u1_U67 (.B( u0_u10_u1_n162 ) , .A( u0_u10_u1_n163 ) , .C2( u0_u10_u1_n164 ) , .ZN( u0_u10_u1_n165 ) , .C1( u0_u10_u1_n171 ) );
  AOI21_X1 u0_u10_u1_U68 (.A( u0_u10_u1_n160 ) , .B2( u0_u10_u1_n161 ) , .ZN( u0_u10_u1_n162 ) , .B1( u0_u10_u1_n182 ) );
  OR2_X1 u0_u10_u1_U69 (.A2( u0_u10_u1_n157 ) , .A1( u0_u10_u1_n158 ) , .ZN( u0_u10_u1_n163 ) );
  NAND2_X1 u0_u10_u1_U7 (.ZN( u0_u10_u1_n114 ) , .A1( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n156 ) );
  NOR2_X1 u0_u10_u1_U70 (.A2( u0_u10_X_7 ) , .A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n95 ) );
  NOR2_X1 u0_u10_u1_U71 (.A1( u0_u10_X_12 ) , .A2( u0_u10_X_9 ) , .ZN( u0_u10_u1_n100 ) );
  NOR2_X1 u0_u10_u1_U72 (.A2( u0_u10_X_8 ) , .A1( u0_u10_u1_n177 ) , .ZN( u0_u10_u1_n99 ) );
  NOR2_X1 u0_u10_u1_U73 (.A2( u0_u10_X_12 ) , .ZN( u0_u10_u1_n102 ) , .A1( u0_u10_u1_n176 ) );
  NOR2_X1 u0_u10_u1_U74 (.A2( u0_u10_X_9 ) , .ZN( u0_u10_u1_n105 ) , .A1( u0_u10_u1_n168 ) );
  NAND2_X1 u0_u10_u1_U75 (.A1( u0_u10_X_10 ) , .ZN( u0_u10_u1_n160 ) , .A2( u0_u10_u1_n169 ) );
  NAND2_X1 u0_u10_u1_U76 (.A2( u0_u10_X_10 ) , .A1( u0_u10_X_11 ) , .ZN( u0_u10_u1_n152 ) );
  NAND2_X1 u0_u10_u1_U77 (.A1( u0_u10_X_11 ) , .ZN( u0_u10_u1_n128 ) , .A2( u0_u10_u1_n170 ) );
  AND2_X1 u0_u10_u1_U78 (.A2( u0_u10_X_7 ) , .A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n104 ) );
  AND2_X1 u0_u10_u1_U79 (.A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n103 ) , .A2( u0_u10_u1_n177 ) );
  NOR2_X1 u0_u10_u1_U8 (.A1( u0_u10_u1_n112 ) , .A2( u0_u10_u1_n116 ) , .ZN( u0_u10_u1_n118 ) );
  INV_X1 u0_u10_u1_U80 (.A( u0_u10_X_10 ) , .ZN( u0_u10_u1_n170 ) );
  INV_X1 u0_u10_u1_U81 (.A( u0_u10_X_9 ) , .ZN( u0_u10_u1_n176 ) );
  INV_X1 u0_u10_u1_U82 (.A( u0_u10_X_11 ) , .ZN( u0_u10_u1_n169 ) );
  INV_X1 u0_u10_u1_U83 (.A( u0_u10_X_12 ) , .ZN( u0_u10_u1_n168 ) );
  INV_X1 u0_u10_u1_U84 (.A( u0_u10_X_7 ) , .ZN( u0_u10_u1_n177 ) );
  NAND4_X1 u0_u10_u1_U85 (.ZN( u0_out10_28 ) , .A4( u0_u10_u1_n124 ) , .A3( u0_u10_u1_n125 ) , .A2( u0_u10_u1_n126 ) , .A1( u0_u10_u1_n127 ) );
  OAI21_X1 u0_u10_u1_U86 (.ZN( u0_u10_u1_n127 ) , .B2( u0_u10_u1_n139 ) , .B1( u0_u10_u1_n175 ) , .A( u0_u10_u1_n183 ) );
  OAI21_X1 u0_u10_u1_U87 (.ZN( u0_u10_u1_n126 ) , .B2( u0_u10_u1_n140 ) , .A( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n178 ) );
  NAND4_X1 u0_u10_u1_U88 (.ZN( u0_out10_18 ) , .A4( u0_u10_u1_n165 ) , .A3( u0_u10_u1_n166 ) , .A1( u0_u10_u1_n167 ) , .A2( u0_u10_u1_n186 ) );
  AOI22_X1 u0_u10_u1_U89 (.B2( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n147 ) , .A2( u0_u10_u1_n148 ) , .ZN( u0_u10_u1_n166 ) , .A1( u0_u10_u1_n172 ) );
  OAI21_X1 u0_u10_u1_U9 (.ZN( u0_u10_u1_n101 ) , .B1( u0_u10_u1_n141 ) , .A( u0_u10_u1_n146 ) , .B2( u0_u10_u1_n183 ) );
  INV_X1 u0_u10_u1_U90 (.A( u0_u10_u1_n145 ) , .ZN( u0_u10_u1_n186 ) );
  NAND4_X1 u0_u10_u1_U91 (.ZN( u0_out10_2 ) , .A4( u0_u10_u1_n142 ) , .A3( u0_u10_u1_n143 ) , .A2( u0_u10_u1_n144 ) , .A1( u0_u10_u1_n179 ) );
  OAI21_X1 u0_u10_u1_U92 (.B2( u0_u10_u1_n132 ) , .ZN( u0_u10_u1_n144 ) , .A( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n180 ) );
  INV_X1 u0_u10_u1_U93 (.A( u0_u10_u1_n130 ) , .ZN( u0_u10_u1_n179 ) );
  OR4_X1 u0_u10_u1_U94 (.ZN( u0_out10_13 ) , .A4( u0_u10_u1_n108 ) , .A3( u0_u10_u1_n109 ) , .A2( u0_u10_u1_n110 ) , .A1( u0_u10_u1_n111 ) );
  AOI21_X1 u0_u10_u1_U95 (.ZN( u0_u10_u1_n111 ) , .A( u0_u10_u1_n128 ) , .B2( u0_u10_u1_n131 ) , .B1( u0_u10_u1_n135 ) );
  AOI21_X1 u0_u10_u1_U96 (.ZN( u0_u10_u1_n110 ) , .A( u0_u10_u1_n116 ) , .B1( u0_u10_u1_n152 ) , .B2( u0_u10_u1_n160 ) );
  NAND3_X1 u0_u10_u1_U97 (.A3( u0_u10_u1_n149 ) , .A2( u0_u10_u1_n150 ) , .A1( u0_u10_u1_n151 ) , .ZN( u0_u10_u1_n164 ) );
  NAND3_X1 u0_u10_u1_U98 (.A3( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n135 ) , .ZN( u0_u10_u1_n136 ) , .A1( u0_u10_u1_n151 ) );
  NAND3_X1 u0_u10_u1_U99 (.A1( u0_u10_u1_n133 ) , .ZN( u0_u10_u1_n137 ) , .A2( u0_u10_u1_n154 ) , .A3( u0_u10_u1_n181 ) );
  OAI22_X1 u0_u10_u2_U10 (.ZN( u0_u10_u2_n109 ) , .A2( u0_u10_u2_n113 ) , .B2( u0_u10_u2_n133 ) , .B1( u0_u10_u2_n167 ) , .A1( u0_u10_u2_n168 ) );
  NAND3_X1 u0_u10_u2_U100 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n98 ) );
  OAI22_X1 u0_u10_u2_U11 (.B1( u0_u10_u2_n151 ) , .A2( u0_u10_u2_n152 ) , .A1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n160 ) , .B2( u0_u10_u2_n168 ) );
  NOR3_X1 u0_u10_u2_U12 (.A1( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n151 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U13 (.ZN( u0_u10_u2_n144 ) , .B2( u0_u10_u2_n155 ) , .A( u0_u10_u2_n172 ) , .B1( u0_u10_u2_n185 ) );
  AOI21_X1 u0_u10_u2_U14 (.B2( u0_u10_u2_n143 ) , .ZN( u0_u10_u2_n145 ) , .B1( u0_u10_u2_n152 ) , .A( u0_u10_u2_n171 ) );
  AOI21_X1 u0_u10_u2_U15 (.B2( u0_u10_u2_n120 ) , .B1( u0_u10_u2_n121 ) , .ZN( u0_u10_u2_n126 ) , .A( u0_u10_u2_n167 ) );
  INV_X1 u0_u10_u2_U16 (.A( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n171 ) );
  INV_X1 u0_u10_u2_U17 (.A( u0_u10_u2_n120 ) , .ZN( u0_u10_u2_n188 ) );
  NAND2_X1 u0_u10_u2_U18 (.A2( u0_u10_u2_n122 ) , .ZN( u0_u10_u2_n150 ) , .A1( u0_u10_u2_n152 ) );
  INV_X1 u0_u10_u2_U19 (.A( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U20 (.A( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n173 ) );
  NAND2_X1 u0_u10_u2_U21 (.A1( u0_u10_u2_n132 ) , .A2( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n157 ) );
  INV_X1 u0_u10_u2_U22 (.A( u0_u10_u2_n113 ) , .ZN( u0_u10_u2_n178 ) );
  INV_X1 u0_u10_u2_U23 (.A( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n175 ) );
  INV_X1 u0_u10_u2_U24 (.A( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n181 ) );
  INV_X1 u0_u10_u2_U25 (.A( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n177 ) );
  INV_X1 u0_u10_u2_U26 (.A( u0_u10_u2_n116 ) , .ZN( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U27 (.A( u0_u10_u2_n131 ) , .ZN( u0_u10_u2_n179 ) );
  INV_X1 u0_u10_u2_U28 (.A( u0_u10_u2_n154 ) , .ZN( u0_u10_u2_n176 ) );
  NAND2_X1 u0_u10_u2_U29 (.A2( u0_u10_u2_n116 ) , .A1( u0_u10_u2_n117 ) , .ZN( u0_u10_u2_n118 ) );
  NOR2_X1 u0_u10_u2_U3 (.ZN( u0_u10_u2_n121 ) , .A2( u0_u10_u2_n177 ) , .A1( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U30 (.A( u0_u10_u2_n132 ) , .ZN( u0_u10_u2_n182 ) );
  INV_X1 u0_u10_u2_U31 (.A( u0_u10_u2_n158 ) , .ZN( u0_u10_u2_n183 ) );
  OAI21_X1 u0_u10_u2_U32 (.A( u0_u10_u2_n156 ) , .B1( u0_u10_u2_n157 ) , .ZN( u0_u10_u2_n158 ) , .B2( u0_u10_u2_n179 ) );
  NOR2_X1 u0_u10_u2_U33 (.ZN( u0_u10_u2_n156 ) , .A1( u0_u10_u2_n166 ) , .A2( u0_u10_u2_n169 ) );
  NOR2_X1 u0_u10_u2_U34 (.A2( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n140 ) );
  NOR2_X1 u0_u10_u2_U35 (.A2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n153 ) , .A1( u0_u10_u2_n156 ) );
  AOI211_X1 u0_u10_u2_U36 (.ZN( u0_u10_u2_n130 ) , .C1( u0_u10_u2_n138 ) , .C2( u0_u10_u2_n179 ) , .B( u0_u10_u2_n96 ) , .A( u0_u10_u2_n97 ) );
  OAI22_X1 u0_u10_u2_U37 (.B1( u0_u10_u2_n133 ) , .A2( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n152 ) , .B2( u0_u10_u2_n168 ) , .ZN( u0_u10_u2_n97 ) );
  OAI221_X1 u0_u10_u2_U38 (.B1( u0_u10_u2_n113 ) , .C1( u0_u10_u2_n132 ) , .A( u0_u10_u2_n149 ) , .B2( u0_u10_u2_n171 ) , .C2( u0_u10_u2_n172 ) , .ZN( u0_u10_u2_n96 ) );
  OAI221_X1 u0_u10_u2_U39 (.A( u0_u10_u2_n115 ) , .C2( u0_u10_u2_n123 ) , .B2( u0_u10_u2_n143 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n163 ) , .C1( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U4 (.A( u0_u10_u2_n134 ) , .ZN( u0_u10_u2_n185 ) );
  OAI21_X1 u0_u10_u2_U40 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n115 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n178 ) );
  OAI221_X1 u0_u10_u2_U41 (.A( u0_u10_u2_n135 ) , .B2( u0_u10_u2_n136 ) , .B1( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n162 ) , .C2( u0_u10_u2_n167 ) , .C1( u0_u10_u2_n185 ) );
  AND3_X1 u0_u10_u2_U42 (.A3( u0_u10_u2_n131 ) , .A2( u0_u10_u2_n132 ) , .A1( u0_u10_u2_n133 ) , .ZN( u0_u10_u2_n136 ) );
  AOI22_X1 u0_u10_u2_U43 (.ZN( u0_u10_u2_n135 ) , .B1( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n156 ) , .B2( u0_u10_u2_n180 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U44 (.ZN( u0_u10_u2_n149 ) , .B1( u0_u10_u2_n173 ) , .B2( u0_u10_u2_n188 ) , .A( u0_u10_u2_n95 ) );
  AND3_X1 u0_u10_u2_U45 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n95 ) );
  OAI21_X1 u0_u10_u2_U46 (.A( u0_u10_u2_n141 ) , .B2( u0_u10_u2_n142 ) , .ZN( u0_u10_u2_n146 ) , .B1( u0_u10_u2_n153 ) );
  OAI21_X1 u0_u10_u2_U47 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n141 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n177 ) );
  NOR3_X1 u0_u10_u2_U48 (.ZN( u0_u10_u2_n142 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n178 ) , .A1( u0_u10_u2_n181 ) );
  OAI21_X1 u0_u10_u2_U49 (.A( u0_u10_u2_n101 ) , .B2( u0_u10_u2_n121 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n164 ) );
  INV_X1 u0_u10_u2_U5 (.A( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n184 ) );
  NAND2_X1 u0_u10_u2_U50 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n155 ) );
  NAND2_X1 u0_u10_u2_U51 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n143 ) );
  NAND2_X1 u0_u10_u2_U52 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n152 ) );
  NAND2_X1 u0_u10_u2_U53 (.A1( u0_u10_u2_n100 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n132 ) );
  INV_X1 u0_u10_u2_U54 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U55 (.A( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n167 ) );
  NAND2_X1 u0_u10_u2_U56 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n113 ) );
  NAND2_X1 u0_u10_u2_U57 (.A1( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n131 ) );
  NAND2_X1 u0_u10_u2_U58 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n139 ) );
  NAND2_X1 u0_u10_u2_U59 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n133 ) );
  NOR4_X1 u0_u10_u2_U6 (.A4( u0_u10_u2_n124 ) , .A3( u0_u10_u2_n125 ) , .A2( u0_u10_u2_n126 ) , .A1( u0_u10_u2_n127 ) , .ZN( u0_u10_u2_n128 ) );
  NAND2_X1 u0_u10_u2_U60 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n103 ) , .ZN( u0_u10_u2_n154 ) );
  NAND2_X1 u0_u10_u2_U61 (.A2( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n104 ) , .ZN( u0_u10_u2_n119 ) );
  NAND2_X1 u0_u10_u2_U62 (.A2( u0_u10_u2_n107 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n123 ) );
  NAND2_X1 u0_u10_u2_U63 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n122 ) );
  INV_X1 u0_u10_u2_U64 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n172 ) );
  NAND2_X1 u0_u10_u2_U65 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n102 ) , .ZN( u0_u10_u2_n116 ) );
  NAND2_X1 u0_u10_u2_U66 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n120 ) );
  NAND2_X1 u0_u10_u2_U67 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n117 ) );
  INV_X1 u0_u10_u2_U68 (.ZN( u0_u10_u2_n187 ) , .A( u0_u10_u2_n99 ) );
  OAI21_X1 u0_u10_u2_U69 (.B1( u0_u10_u2_n137 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n98 ) , .ZN( u0_u10_u2_n99 ) );
  AOI21_X1 u0_u10_u2_U7 (.ZN( u0_u10_u2_n124 ) , .B1( u0_u10_u2_n131 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n172 ) );
  NOR2_X1 u0_u10_u2_U70 (.A2( u0_u10_X_16 ) , .ZN( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n166 ) );
  NOR2_X1 u0_u10_u2_U71 (.A2( u0_u10_X_13 ) , .A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n100 ) );
  NOR2_X1 u0_u10_u2_U72 (.A2( u0_u10_X_16 ) , .A1( u0_u10_X_17 ) , .ZN( u0_u10_u2_n138 ) );
  NOR2_X1 u0_u10_u2_U73 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n104 ) );
  NOR2_X1 u0_u10_u2_U74 (.A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n174 ) );
  NOR2_X1 u0_u10_u2_U75 (.A2( u0_u10_X_15 ) , .ZN( u0_u10_u2_n102 ) , .A1( u0_u10_u2_n165 ) );
  NOR2_X1 u0_u10_u2_U76 (.A2( u0_u10_X_17 ) , .ZN( u0_u10_u2_n114 ) , .A1( u0_u10_u2_n169 ) );
  AND2_X1 u0_u10_u2_U77 (.A1( u0_u10_X_15 ) , .ZN( u0_u10_u2_n105 ) , .A2( u0_u10_u2_n165 ) );
  AND2_X1 u0_u10_u2_U78 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n107 ) );
  AND2_X1 u0_u10_u2_U79 (.A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n174 ) );
  AOI21_X1 u0_u10_u2_U8 (.B2( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n127 ) , .A( u0_u10_u2_n137 ) , .B1( u0_u10_u2_n155 ) );
  AND2_X1 u0_u10_u2_U80 (.A1( u0_u10_X_13 ) , .A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n108 ) );
  INV_X1 u0_u10_u2_U81 (.A( u0_u10_X_16 ) , .ZN( u0_u10_u2_n169 ) );
  INV_X1 u0_u10_u2_U82 (.A( u0_u10_X_17 ) , .ZN( u0_u10_u2_n166 ) );
  INV_X1 u0_u10_u2_U83 (.A( u0_u10_X_13 ) , .ZN( u0_u10_u2_n174 ) );
  INV_X1 u0_u10_u2_U84 (.A( u0_u10_X_18 ) , .ZN( u0_u10_u2_n165 ) );
  NAND4_X1 u0_u10_u2_U85 (.ZN( u0_out10_30 ) , .A4( u0_u10_u2_n147 ) , .A3( u0_u10_u2_n148 ) , .A2( u0_u10_u2_n149 ) , .A1( u0_u10_u2_n187 ) );
  NOR3_X1 u0_u10_u2_U86 (.A3( u0_u10_u2_n144 ) , .A2( u0_u10_u2_n145 ) , .A1( u0_u10_u2_n146 ) , .ZN( u0_u10_u2_n147 ) );
  AOI21_X1 u0_u10_u2_U87 (.B2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n148 ) , .A( u0_u10_u2_n162 ) , .B1( u0_u10_u2_n182 ) );
  NAND4_X1 u0_u10_u2_U88 (.ZN( u0_out10_24 ) , .A4( u0_u10_u2_n111 ) , .A3( u0_u10_u2_n112 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n187 ) );
  AOI221_X1 u0_u10_u2_U89 (.A( u0_u10_u2_n109 ) , .B1( u0_u10_u2_n110 ) , .ZN( u0_u10_u2_n111 ) , .C1( u0_u10_u2_n134 ) , .C2( u0_u10_u2_n170 ) , .B2( u0_u10_u2_n173 ) );
  AOI21_X1 u0_u10_u2_U9 (.B2( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n125 ) , .A( u0_u10_u2_n171 ) , .B1( u0_u10_u2_n184 ) );
  AOI21_X1 u0_u10_u2_U90 (.ZN( u0_u10_u2_n112 ) , .B2( u0_u10_u2_n156 ) , .A( u0_u10_u2_n164 ) , .B1( u0_u10_u2_n181 ) );
  NAND4_X1 u0_u10_u2_U91 (.ZN( u0_out10_16 ) , .A4( u0_u10_u2_n128 ) , .A3( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n186 ) );
  AOI22_X1 u0_u10_u2_U92 (.A2( u0_u10_u2_n118 ) , .ZN( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n140 ) , .B1( u0_u10_u2_n157 ) , .B2( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U93 (.A( u0_u10_u2_n163 ) , .ZN( u0_u10_u2_n186 ) );
  OR4_X1 u0_u10_u2_U94 (.ZN( u0_out10_6 ) , .A4( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n162 ) , .A2( u0_u10_u2_n163 ) , .A1( u0_u10_u2_n164 ) );
  OR3_X1 u0_u10_u2_U95 (.A2( u0_u10_u2_n159 ) , .A1( u0_u10_u2_n160 ) , .ZN( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n183 ) );
  AOI21_X1 u0_u10_u2_U96 (.B2( u0_u10_u2_n154 ) , .B1( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n159 ) , .A( u0_u10_u2_n167 ) );
  NAND3_X1 u0_u10_u2_U97 (.A2( u0_u10_u2_n117 ) , .A1( u0_u10_u2_n122 ) , .A3( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n134 ) );
  NAND3_X1 u0_u10_u2_U98 (.ZN( u0_u10_u2_n110 ) , .A2( u0_u10_u2_n131 ) , .A3( u0_u10_u2_n139 ) , .A1( u0_u10_u2_n154 ) );
  NAND3_X1 u0_u10_u2_U99 (.A2( u0_u10_u2_n100 ) , .ZN( u0_u10_u2_n101 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n114 ) );
  OAI22_X1 u0_u10_u3_U10 (.B1( u0_u10_u3_n113 ) , .A2( u0_u10_u3_n135 ) , .A1( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n164 ) , .ZN( u0_u10_u3_n98 ) );
  OAI211_X1 u0_u10_u3_U11 (.B( u0_u10_u3_n106 ) , .ZN( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n128 ) , .C1( u0_u10_u3_n167 ) , .A( u0_u10_u3_n181 ) );
  AOI221_X1 u0_u10_u3_U12 (.C1( u0_u10_u3_n105 ) , .ZN( u0_u10_u3_n106 ) , .A( u0_u10_u3_n131 ) , .B2( u0_u10_u3_n132 ) , .C2( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n169 ) );
  INV_X1 u0_u10_u3_U13 (.ZN( u0_u10_u3_n181 ) , .A( u0_u10_u3_n98 ) );
  NAND2_X1 u0_u10_u3_U14 (.ZN( u0_u10_u3_n105 ) , .A2( u0_u10_u3_n130 ) , .A1( u0_u10_u3_n155 ) );
  AOI22_X1 u0_u10_u3_U15 (.B1( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n116 ) , .ZN( u0_u10_u3_n123 ) , .B2( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U16 (.ZN( u0_u10_u3_n116 ) , .A2( u0_u10_u3_n151 ) , .A1( u0_u10_u3_n182 ) );
  NOR2_X1 u0_u10_u3_U17 (.ZN( u0_u10_u3_n126 ) , .A2( u0_u10_u3_n150 ) , .A1( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U18 (.ZN( u0_u10_u3_n112 ) , .B2( u0_u10_u3_n146 ) , .B1( u0_u10_u3_n155 ) , .A( u0_u10_u3_n167 ) );
  NAND2_X1 u0_u10_u3_U19 (.A1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n142 ) , .A2( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U20 (.ZN( u0_u10_u3_n132 ) , .A2( u0_u10_u3_n152 ) , .A1( u0_u10_u3_n156 ) );
  AND2_X1 u0_u10_u3_U21 (.A2( u0_u10_u3_n113 ) , .A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n151 ) );
  INV_X1 u0_u10_u3_U22 (.A( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n165 ) );
  INV_X1 u0_u10_u3_U23 (.A( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n170 ) );
  NAND2_X1 u0_u10_u3_U24 (.A1( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .ZN( u0_u10_u3_n140 ) );
  NAND2_X1 u0_u10_u3_U25 (.ZN( u0_u10_u3_n117 ) , .A1( u0_u10_u3_n124 ) , .A2( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U26 (.ZN( u0_u10_u3_n143 ) , .A1( u0_u10_u3_n165 ) , .A2( u0_u10_u3_n167 ) );
  INV_X1 u0_u10_u3_U27 (.A( u0_u10_u3_n130 ) , .ZN( u0_u10_u3_n177 ) );
  INV_X1 u0_u10_u3_U28 (.A( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n176 ) );
  INV_X1 u0_u10_u3_U29 (.A( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n174 ) );
  INV_X1 u0_u10_u3_U3 (.A( u0_u10_u3_n129 ) , .ZN( u0_u10_u3_n183 ) );
  INV_X1 u0_u10_u3_U30 (.A( u0_u10_u3_n139 ) , .ZN( u0_u10_u3_n185 ) );
  NOR2_X1 u0_u10_u3_U31 (.ZN( u0_u10_u3_n135 ) , .A2( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n169 ) );
  OAI222_X1 u0_u10_u3_U32 (.C2( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .B1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n138 ) , .B2( u0_u10_u3_n146 ) , .C1( u0_u10_u3_n154 ) , .A1( u0_u10_u3_n164 ) );
  NOR4_X1 u0_u10_u3_U33 (.A4( u0_u10_u3_n157 ) , .A3( u0_u10_u3_n158 ) , .A2( u0_u10_u3_n159 ) , .A1( u0_u10_u3_n160 ) , .ZN( u0_u10_u3_n161 ) );
  AOI21_X1 u0_u10_u3_U34 (.B2( u0_u10_u3_n152 ) , .B1( u0_u10_u3_n153 ) , .ZN( u0_u10_u3_n158 ) , .A( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U35 (.A( u0_u10_u3_n154 ) , .B2( u0_u10_u3_n155 ) , .B1( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n157 ) );
  AOI21_X1 u0_u10_u3_U36 (.A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n150 ) , .B1( u0_u10_u3_n151 ) , .ZN( u0_u10_u3_n159 ) );
  AOI211_X1 u0_u10_u3_U37 (.ZN( u0_u10_u3_n109 ) , .A( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n129 ) , .B( u0_u10_u3_n138 ) , .C1( u0_u10_u3_n141 ) );
  AOI211_X1 u0_u10_u3_U38 (.B( u0_u10_u3_n119 ) , .A( u0_u10_u3_n120 ) , .C2( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n122 ) , .C1( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U39 (.A( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U4 (.A( u0_u10_u3_n140 ) , .ZN( u0_u10_u3_n182 ) );
  OAI22_X1 u0_u10_u3_U40 (.B1( u0_u10_u3_n118 ) , .ZN( u0_u10_u3_n120 ) , .A1( u0_u10_u3_n135 ) , .B2( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n178 ) );
  AND3_X1 u0_u10_u3_U41 (.ZN( u0_u10_u3_n118 ) , .A2( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n144 ) , .A3( u0_u10_u3_n152 ) );
  INV_X1 u0_u10_u3_U42 (.A( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U43 (.ZN( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n164 ) );
  OAI211_X1 u0_u10_u3_U44 (.B( u0_u10_u3_n127 ) , .ZN( u0_u10_u3_n139 ) , .C1( u0_u10_u3_n150 ) , .C2( u0_u10_u3_n154 ) , .A( u0_u10_u3_n184 ) );
  INV_X1 u0_u10_u3_U45 (.A( u0_u10_u3_n125 ) , .ZN( u0_u10_u3_n184 ) );
  AOI221_X1 u0_u10_u3_U46 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n127 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n169 ) , .B2( u0_u10_u3_n170 ) , .B1( u0_u10_u3_n174 ) );
  OAI22_X1 u0_u10_u3_U47 (.A1( u0_u10_u3_n124 ) , .ZN( u0_u10_u3_n125 ) , .B2( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n165 ) , .B1( u0_u10_u3_n167 ) );
  NOR2_X1 u0_u10_u3_U48 (.A1( u0_u10_u3_n113 ) , .ZN( u0_u10_u3_n131 ) , .A2( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U49 (.A1( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n150 ) , .A2( u0_u10_u3_n99 ) );
  INV_X1 u0_u10_u3_U5 (.A( u0_u10_u3_n117 ) , .ZN( u0_u10_u3_n178 ) );
  NAND2_X1 u0_u10_u3_U50 (.A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n155 ) , .A1( u0_u10_u3_n97 ) );
  INV_X1 u0_u10_u3_U51 (.A( u0_u10_u3_n141 ) , .ZN( u0_u10_u3_n167 ) );
  AOI21_X1 u0_u10_u3_U52 (.B2( u0_u10_u3_n114 ) , .B1( u0_u10_u3_n146 ) , .A( u0_u10_u3_n154 ) , .ZN( u0_u10_u3_n94 ) );
  AOI21_X1 u0_u10_u3_U53 (.ZN( u0_u10_u3_n110 ) , .B2( u0_u10_u3_n142 ) , .B1( u0_u10_u3_n186 ) , .A( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U54 (.A( u0_u10_u3_n145 ) , .ZN( u0_u10_u3_n186 ) );
  AOI21_X1 u0_u10_u3_U55 (.B1( u0_u10_u3_n124 ) , .A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U56 (.A( u0_u10_u3_n149 ) , .ZN( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U57 (.ZN( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n96 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U58 (.A2( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n146 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U59 (.A1( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n99 ) );
  AOI221_X1 u0_u10_u3_U6 (.A( u0_u10_u3_n131 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n134 ) , .B1( u0_u10_u3_n143 ) , .B2( u0_u10_u3_n177 ) );
  NAND2_X1 u0_u10_u3_U60 (.A1( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n156 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U61 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U62 (.A1( u0_u10_u3_n100 ) , .A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n128 ) );
  NAND2_X1 u0_u10_u3_U63 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n152 ) );
  NAND2_X1 u0_u10_u3_U64 (.A2( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n114 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U65 (.ZN( u0_u10_u3_n107 ) , .A1( u0_u10_u3_n97 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U66 (.A2( u0_u10_u3_n100 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n113 ) );
  NAND2_X1 u0_u10_u3_U67 (.A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n153 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U68 (.A2( u0_u10_u3_n103 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n130 ) );
  NAND2_X1 u0_u10_u3_U69 (.A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n96 ) );
  OAI22_X1 u0_u10_u3_U7 (.B2( u0_u10_u3_n147 ) , .A2( u0_u10_u3_n148 ) , .ZN( u0_u10_u3_n160 ) , .B1( u0_u10_u3_n165 ) , .A1( u0_u10_u3_n168 ) );
  NAND2_X1 u0_u10_u3_U70 (.A1( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n108 ) );
  NOR2_X1 u0_u10_u3_U71 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n99 ) );
  NOR2_X1 u0_u10_u3_U72 (.A2( u0_u10_X_21 ) , .A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n103 ) );
  NOR2_X1 u0_u10_u3_U73 (.A2( u0_u10_X_24 ) , .A1( u0_u10_u3_n171 ) , .ZN( u0_u10_u3_n97 ) );
  NOR2_X1 u0_u10_u3_U74 (.A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U75 (.A2( u0_u10_X_19 ) , .A1( u0_u10_u3_n172 ) , .ZN( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U76 (.A1( u0_u10_X_22 ) , .A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U77 (.A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n149 ) , .A2( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U78 (.A2( u0_u10_X_22 ) , .A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n121 ) );
  AND2_X1 u0_u10_u3_U79 (.A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n101 ) , .A2( u0_u10_u3_n171 ) );
  AND3_X1 u0_u10_u3_U8 (.A3( u0_u10_u3_n144 ) , .A2( u0_u10_u3_n145 ) , .A1( u0_u10_u3_n146 ) , .ZN( u0_u10_u3_n147 ) );
  AND2_X1 u0_u10_u3_U80 (.A1( u0_u10_X_19 ) , .ZN( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n172 ) );
  AND2_X1 u0_u10_u3_U81 (.A1( u0_u10_X_21 ) , .A2( u0_u10_X_24 ) , .ZN( u0_u10_u3_n100 ) );
  AND2_X1 u0_u10_u3_U82 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n104 ) );
  INV_X1 u0_u10_u3_U83 (.A( u0_u10_X_22 ) , .ZN( u0_u10_u3_n166 ) );
  INV_X1 u0_u10_u3_U84 (.A( u0_u10_X_21 ) , .ZN( u0_u10_u3_n171 ) );
  INV_X1 u0_u10_u3_U85 (.A( u0_u10_X_20 ) , .ZN( u0_u10_u3_n172 ) );
  OR4_X1 u0_u10_u3_U86 (.ZN( u0_out10_10 ) , .A4( u0_u10_u3_n136 ) , .A3( u0_u10_u3_n137 ) , .A1( u0_u10_u3_n138 ) , .A2( u0_u10_u3_n139 ) );
  OAI222_X1 u0_u10_u3_U87 (.C1( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n137 ) , .B1( u0_u10_u3_n148 ) , .A2( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n154 ) , .C2( u0_u10_u3_n164 ) , .A1( u0_u10_u3_n167 ) );
  OAI221_X1 u0_u10_u3_U88 (.A( u0_u10_u3_n134 ) , .B2( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n136 ) , .C1( u0_u10_u3_n149 ) , .B1( u0_u10_u3_n151 ) , .C2( u0_u10_u3_n183 ) );
  NAND4_X1 u0_u10_u3_U89 (.ZN( u0_out10_26 ) , .A4( u0_u10_u3_n109 ) , .A3( u0_u10_u3_n110 ) , .A2( u0_u10_u3_n111 ) , .A1( u0_u10_u3_n173 ) );
  INV_X1 u0_u10_u3_U9 (.A( u0_u10_u3_n143 ) , .ZN( u0_u10_u3_n168 ) );
  INV_X1 u0_u10_u3_U90 (.ZN( u0_u10_u3_n173 ) , .A( u0_u10_u3_n94 ) );
  OAI21_X1 u0_u10_u3_U91 (.ZN( u0_u10_u3_n111 ) , .B2( u0_u10_u3_n117 ) , .A( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n176 ) );
  NAND4_X1 u0_u10_u3_U92 (.ZN( u0_out10_20 ) , .A4( u0_u10_u3_n122 ) , .A3( u0_u10_u3_n123 ) , .A1( u0_u10_u3_n175 ) , .A2( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U93 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U94 (.A( u0_u10_u3_n112 ) , .ZN( u0_u10_u3_n175 ) );
  NAND4_X1 u0_u10_u3_U95 (.ZN( u0_out10_1 ) , .A4( u0_u10_u3_n161 ) , .A3( u0_u10_u3_n162 ) , .A2( u0_u10_u3_n163 ) , .A1( u0_u10_u3_n185 ) );
  NAND2_X1 u0_u10_u3_U96 (.ZN( u0_u10_u3_n163 ) , .A2( u0_u10_u3_n170 ) , .A1( u0_u10_u3_n176 ) );
  AOI22_X1 u0_u10_u3_U97 (.B2( u0_u10_u3_n140 ) , .B1( u0_u10_u3_n141 ) , .A2( u0_u10_u3_n142 ) , .ZN( u0_u10_u3_n162 ) , .A1( u0_u10_u3_n177 ) );
  NAND3_X1 u0_u10_u3_U98 (.A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n145 ) , .A3( u0_u10_u3_n153 ) );
  NAND3_X1 u0_u10_u3_U99 (.ZN( u0_u10_u3_n129 ) , .A2( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n153 ) , .A3( u0_u10_u3_n182 ) );
  INV_X1 u0_u10_u5_U10 (.A( u0_u10_u5_n121 ) , .ZN( u0_u10_u5_n177 ) );
  NOR3_X1 u0_u10_u5_U100 (.A3( u0_u10_u5_n141 ) , .A1( u0_u10_u5_n142 ) , .ZN( u0_u10_u5_n143 ) , .A2( u0_u10_u5_n191 ) );
  NAND4_X1 u0_u10_u5_U101 (.ZN( u0_out10_4 ) , .A4( u0_u10_u5_n112 ) , .A2( u0_u10_u5_n113 ) , .A1( u0_u10_u5_n114 ) , .A3( u0_u10_u5_n195 ) );
  AOI211_X1 u0_u10_u5_U102 (.A( u0_u10_u5_n110 ) , .C1( u0_u10_u5_n111 ) , .ZN( u0_u10_u5_n112 ) , .B( u0_u10_u5_n118 ) , .C2( u0_u10_u5_n177 ) );
  AOI222_X1 u0_u10_u5_U103 (.ZN( u0_u10_u5_n113 ) , .A1( u0_u10_u5_n131 ) , .C1( u0_u10_u5_n148 ) , .B2( u0_u10_u5_n174 ) , .C2( u0_u10_u5_n178 ) , .A2( u0_u10_u5_n179 ) , .B1( u0_u10_u5_n99 ) );
  NAND3_X1 u0_u10_u5_U104 (.A2( u0_u10_u5_n154 ) , .A3( u0_u10_u5_n158 ) , .A1( u0_u10_u5_n161 ) , .ZN( u0_u10_u5_n99 ) );
  NOR2_X1 u0_u10_u5_U11 (.ZN( u0_u10_u5_n160 ) , .A2( u0_u10_u5_n173 ) , .A1( u0_u10_u5_n177 ) );
  INV_X1 u0_u10_u5_U12 (.A( u0_u10_u5_n150 ) , .ZN( u0_u10_u5_n174 ) );
  AOI21_X1 u0_u10_u5_U13 (.A( u0_u10_u5_n160 ) , .B2( u0_u10_u5_n161 ) , .ZN( u0_u10_u5_n162 ) , .B1( u0_u10_u5_n192 ) );
  INV_X1 u0_u10_u5_U14 (.A( u0_u10_u5_n159 ) , .ZN( u0_u10_u5_n192 ) );
  AOI21_X1 u0_u10_u5_U15 (.A( u0_u10_u5_n156 ) , .B2( u0_u10_u5_n157 ) , .B1( u0_u10_u5_n158 ) , .ZN( u0_u10_u5_n163 ) );
  AOI21_X1 u0_u10_u5_U16 (.B2( u0_u10_u5_n139 ) , .B1( u0_u10_u5_n140 ) , .ZN( u0_u10_u5_n141 ) , .A( u0_u10_u5_n150 ) );
  OAI21_X1 u0_u10_u5_U17 (.A( u0_u10_u5_n133 ) , .B2( u0_u10_u5_n134 ) , .B1( u0_u10_u5_n135 ) , .ZN( u0_u10_u5_n142 ) );
  OAI21_X1 u0_u10_u5_U18 (.ZN( u0_u10_u5_n133 ) , .B2( u0_u10_u5_n147 ) , .A( u0_u10_u5_n173 ) , .B1( u0_u10_u5_n188 ) );
  NAND2_X1 u0_u10_u5_U19 (.A2( u0_u10_u5_n119 ) , .A1( u0_u10_u5_n123 ) , .ZN( u0_u10_u5_n137 ) );
  INV_X1 u0_u10_u5_U20 (.A( u0_u10_u5_n155 ) , .ZN( u0_u10_u5_n194 ) );
  NAND2_X1 u0_u10_u5_U21 (.A1( u0_u10_u5_n121 ) , .ZN( u0_u10_u5_n132 ) , .A2( u0_u10_u5_n172 ) );
  NAND2_X1 u0_u10_u5_U22 (.A2( u0_u10_u5_n122 ) , .ZN( u0_u10_u5_n136 ) , .A1( u0_u10_u5_n154 ) );
  NAND2_X1 u0_u10_u5_U23 (.A2( u0_u10_u5_n119 ) , .A1( u0_u10_u5_n120 ) , .ZN( u0_u10_u5_n159 ) );
  INV_X1 u0_u10_u5_U24 (.A( u0_u10_u5_n156 ) , .ZN( u0_u10_u5_n175 ) );
  INV_X1 u0_u10_u5_U25 (.A( u0_u10_u5_n158 ) , .ZN( u0_u10_u5_n188 ) );
  INV_X1 u0_u10_u5_U26 (.A( u0_u10_u5_n152 ) , .ZN( u0_u10_u5_n179 ) );
  INV_X1 u0_u10_u5_U27 (.A( u0_u10_u5_n140 ) , .ZN( u0_u10_u5_n182 ) );
  INV_X1 u0_u10_u5_U28 (.A( u0_u10_u5_n151 ) , .ZN( u0_u10_u5_n183 ) );
  INV_X1 u0_u10_u5_U29 (.A( u0_u10_u5_n123 ) , .ZN( u0_u10_u5_n185 ) );
  NOR2_X1 u0_u10_u5_U3 (.ZN( u0_u10_u5_n134 ) , .A1( u0_u10_u5_n183 ) , .A2( u0_u10_u5_n190 ) );
  INV_X1 u0_u10_u5_U30 (.A( u0_u10_u5_n161 ) , .ZN( u0_u10_u5_n184 ) );
  INV_X1 u0_u10_u5_U31 (.A( u0_u10_u5_n139 ) , .ZN( u0_u10_u5_n189 ) );
  INV_X1 u0_u10_u5_U32 (.A( u0_u10_u5_n157 ) , .ZN( u0_u10_u5_n190 ) );
  INV_X1 u0_u10_u5_U33 (.A( u0_u10_u5_n120 ) , .ZN( u0_u10_u5_n193 ) );
  NAND2_X1 u0_u10_u5_U34 (.ZN( u0_u10_u5_n111 ) , .A1( u0_u10_u5_n140 ) , .A2( u0_u10_u5_n155 ) );
  NOR2_X1 u0_u10_u5_U35 (.ZN( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n170 ) , .A2( u0_u10_u5_n180 ) );
  INV_X1 u0_u10_u5_U36 (.A( u0_u10_u5_n117 ) , .ZN( u0_u10_u5_n196 ) );
  OAI221_X1 u0_u10_u5_U37 (.A( u0_u10_u5_n116 ) , .ZN( u0_u10_u5_n117 ) , .B2( u0_u10_u5_n119 ) , .C1( u0_u10_u5_n153 ) , .C2( u0_u10_u5_n158 ) , .B1( u0_u10_u5_n172 ) );
  AOI222_X1 u0_u10_u5_U38 (.ZN( u0_u10_u5_n116 ) , .B2( u0_u10_u5_n145 ) , .C1( u0_u10_u5_n148 ) , .A2( u0_u10_u5_n174 ) , .C2( u0_u10_u5_n177 ) , .B1( u0_u10_u5_n187 ) , .A1( u0_u10_u5_n193 ) );
  INV_X1 u0_u10_u5_U39 (.A( u0_u10_u5_n115 ) , .ZN( u0_u10_u5_n187 ) );
  INV_X1 u0_u10_u5_U4 (.A( u0_u10_u5_n138 ) , .ZN( u0_u10_u5_n191 ) );
  AOI22_X1 u0_u10_u5_U40 (.B2( u0_u10_u5_n131 ) , .A2( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n169 ) , .B1( u0_u10_u5_n174 ) , .A1( u0_u10_u5_n185 ) );
  NOR2_X1 u0_u10_u5_U41 (.A1( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n150 ) , .A2( u0_u10_u5_n173 ) );
  AOI21_X1 u0_u10_u5_U42 (.A( u0_u10_u5_n118 ) , .B2( u0_u10_u5_n145 ) , .ZN( u0_u10_u5_n168 ) , .B1( u0_u10_u5_n186 ) );
  INV_X1 u0_u10_u5_U43 (.A( u0_u10_u5_n122 ) , .ZN( u0_u10_u5_n186 ) );
  NOR2_X1 u0_u10_u5_U44 (.A1( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n152 ) , .A2( u0_u10_u5_n176 ) );
  NOR2_X1 u0_u10_u5_U45 (.A1( u0_u10_u5_n115 ) , .ZN( u0_u10_u5_n118 ) , .A2( u0_u10_u5_n153 ) );
  NOR2_X1 u0_u10_u5_U46 (.A2( u0_u10_u5_n145 ) , .ZN( u0_u10_u5_n156 ) , .A1( u0_u10_u5_n174 ) );
  NOR2_X1 u0_u10_u5_U47 (.ZN( u0_u10_u5_n121 ) , .A2( u0_u10_u5_n145 ) , .A1( u0_u10_u5_n176 ) );
  AOI22_X1 u0_u10_u5_U48 (.ZN( u0_u10_u5_n114 ) , .A2( u0_u10_u5_n137 ) , .A1( u0_u10_u5_n145 ) , .B2( u0_u10_u5_n175 ) , .B1( u0_u10_u5_n193 ) );
  OAI211_X1 u0_u10_u5_U49 (.B( u0_u10_u5_n124 ) , .A( u0_u10_u5_n125 ) , .C2( u0_u10_u5_n126 ) , .C1( u0_u10_u5_n127 ) , .ZN( u0_u10_u5_n128 ) );
  OAI21_X1 u0_u10_u5_U5 (.B2( u0_u10_u5_n136 ) , .B1( u0_u10_u5_n137 ) , .ZN( u0_u10_u5_n138 ) , .A( u0_u10_u5_n177 ) );
  NOR3_X1 u0_u10_u5_U50 (.ZN( u0_u10_u5_n127 ) , .A1( u0_u10_u5_n136 ) , .A3( u0_u10_u5_n148 ) , .A2( u0_u10_u5_n182 ) );
  OAI21_X1 u0_u10_u5_U51 (.ZN( u0_u10_u5_n124 ) , .A( u0_u10_u5_n177 ) , .B2( u0_u10_u5_n183 ) , .B1( u0_u10_u5_n189 ) );
  OAI21_X1 u0_u10_u5_U52 (.ZN( u0_u10_u5_n125 ) , .A( u0_u10_u5_n174 ) , .B2( u0_u10_u5_n185 ) , .B1( u0_u10_u5_n190 ) );
  AOI21_X1 u0_u10_u5_U53 (.A( u0_u10_u5_n153 ) , .B2( u0_u10_u5_n154 ) , .B1( u0_u10_u5_n155 ) , .ZN( u0_u10_u5_n164 ) );
  AOI21_X1 u0_u10_u5_U54 (.ZN( u0_u10_u5_n110 ) , .B1( u0_u10_u5_n122 ) , .B2( u0_u10_u5_n139 ) , .A( u0_u10_u5_n153 ) );
  INV_X1 u0_u10_u5_U55 (.A( u0_u10_u5_n153 ) , .ZN( u0_u10_u5_n176 ) );
  INV_X1 u0_u10_u5_U56 (.A( u0_u10_u5_n126 ) , .ZN( u0_u10_u5_n173 ) );
  AND2_X1 u0_u10_u5_U57 (.A2( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n107 ) , .ZN( u0_u10_u5_n147 ) );
  AND2_X1 u0_u10_u5_U58 (.A2( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n108 ) , .ZN( u0_u10_u5_n148 ) );
  NAND2_X1 u0_u10_u5_U59 (.A1( u0_u10_u5_n105 ) , .A2( u0_u10_u5_n106 ) , .ZN( u0_u10_u5_n158 ) );
  INV_X1 u0_u10_u5_U6 (.A( u0_u10_u5_n135 ) , .ZN( u0_u10_u5_n178 ) );
  NAND2_X1 u0_u10_u5_U60 (.A2( u0_u10_u5_n108 ) , .A1( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n139 ) );
  NAND2_X1 u0_u10_u5_U61 (.A1( u0_u10_u5_n106 ) , .A2( u0_u10_u5_n108 ) , .ZN( u0_u10_u5_n119 ) );
  NAND2_X1 u0_u10_u5_U62 (.A2( u0_u10_u5_n103 ) , .A1( u0_u10_u5_n105 ) , .ZN( u0_u10_u5_n140 ) );
  NAND2_X1 u0_u10_u5_U63 (.A2( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n105 ) , .ZN( u0_u10_u5_n155 ) );
  NAND2_X1 u0_u10_u5_U64 (.A2( u0_u10_u5_n106 ) , .A1( u0_u10_u5_n107 ) , .ZN( u0_u10_u5_n122 ) );
  NAND2_X1 u0_u10_u5_U65 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n106 ) , .ZN( u0_u10_u5_n115 ) );
  NAND2_X1 u0_u10_u5_U66 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n103 ) , .ZN( u0_u10_u5_n161 ) );
  NAND2_X1 u0_u10_u5_U67 (.A1( u0_u10_u5_n105 ) , .A2( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n154 ) );
  INV_X1 u0_u10_u5_U68 (.A( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n172 ) );
  NAND2_X1 u0_u10_u5_U69 (.A1( u0_u10_u5_n103 ) , .A2( u0_u10_u5_n108 ) , .ZN( u0_u10_u5_n123 ) );
  OAI22_X1 u0_u10_u5_U7 (.B2( u0_u10_u5_n149 ) , .B1( u0_u10_u5_n150 ) , .A2( u0_u10_u5_n151 ) , .A1( u0_u10_u5_n152 ) , .ZN( u0_u10_u5_n165 ) );
  NAND2_X1 u0_u10_u5_U70 (.A2( u0_u10_u5_n103 ) , .A1( u0_u10_u5_n107 ) , .ZN( u0_u10_u5_n151 ) );
  NAND2_X1 u0_u10_u5_U71 (.A2( u0_u10_u5_n107 ) , .A1( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n120 ) );
  NAND2_X1 u0_u10_u5_U72 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n157 ) );
  AND2_X1 u0_u10_u5_U73 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n104 ) , .ZN( u0_u10_u5_n131 ) );
  INV_X1 u0_u10_u5_U74 (.A( u0_u10_u5_n102 ) , .ZN( u0_u10_u5_n195 ) );
  OAI221_X1 u0_u10_u5_U75 (.A( u0_u10_u5_n101 ) , .ZN( u0_u10_u5_n102 ) , .C2( u0_u10_u5_n115 ) , .C1( u0_u10_u5_n126 ) , .B1( u0_u10_u5_n134 ) , .B2( u0_u10_u5_n160 ) );
  OAI21_X1 u0_u10_u5_U76 (.ZN( u0_u10_u5_n101 ) , .B1( u0_u10_u5_n137 ) , .A( u0_u10_u5_n146 ) , .B2( u0_u10_u5_n147 ) );
  NOR2_X1 u0_u10_u5_U77 (.A2( u0_u10_X_34 ) , .A1( u0_u10_X_35 ) , .ZN( u0_u10_u5_n145 ) );
  NOR2_X1 u0_u10_u5_U78 (.A2( u0_u10_X_34 ) , .ZN( u0_u10_u5_n146 ) , .A1( u0_u10_u5_n171 ) );
  NOR2_X1 u0_u10_u5_U79 (.A2( u0_u10_X_31 ) , .A1( u0_u10_X_32 ) , .ZN( u0_u10_u5_n103 ) );
  NOR3_X1 u0_u10_u5_U8 (.A2( u0_u10_u5_n147 ) , .A1( u0_u10_u5_n148 ) , .ZN( u0_u10_u5_n149 ) , .A3( u0_u10_u5_n194 ) );
  NOR2_X1 u0_u10_u5_U80 (.A2( u0_u10_X_36 ) , .ZN( u0_u10_u5_n105 ) , .A1( u0_u10_u5_n180 ) );
  NOR2_X1 u0_u10_u5_U81 (.A2( u0_u10_X_33 ) , .ZN( u0_u10_u5_n108 ) , .A1( u0_u10_u5_n170 ) );
  NOR2_X1 u0_u10_u5_U82 (.A2( u0_u10_X_33 ) , .A1( u0_u10_X_36 ) , .ZN( u0_u10_u5_n107 ) );
  NOR2_X1 u0_u10_u5_U83 (.A2( u0_u10_X_31 ) , .ZN( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n181 ) );
  NAND2_X1 u0_u10_u5_U84 (.A2( u0_u10_X_34 ) , .A1( u0_u10_X_35 ) , .ZN( u0_u10_u5_n153 ) );
  NAND2_X1 u0_u10_u5_U85 (.A1( u0_u10_X_34 ) , .ZN( u0_u10_u5_n126 ) , .A2( u0_u10_u5_n171 ) );
  AND2_X1 u0_u10_u5_U86 (.A1( u0_u10_X_31 ) , .A2( u0_u10_X_32 ) , .ZN( u0_u10_u5_n106 ) );
  AND2_X1 u0_u10_u5_U87 (.A1( u0_u10_X_31 ) , .ZN( u0_u10_u5_n109 ) , .A2( u0_u10_u5_n181 ) );
  INV_X1 u0_u10_u5_U88 (.A( u0_u10_X_33 ) , .ZN( u0_u10_u5_n180 ) );
  INV_X1 u0_u10_u5_U89 (.A( u0_u10_X_35 ) , .ZN( u0_u10_u5_n171 ) );
  NOR2_X1 u0_u10_u5_U9 (.ZN( u0_u10_u5_n135 ) , .A1( u0_u10_u5_n173 ) , .A2( u0_u10_u5_n176 ) );
  INV_X1 u0_u10_u5_U90 (.A( u0_u10_X_36 ) , .ZN( u0_u10_u5_n170 ) );
  INV_X1 u0_u10_u5_U91 (.A( u0_u10_X_32 ) , .ZN( u0_u10_u5_n181 ) );
  NAND4_X1 u0_u10_u5_U92 (.ZN( u0_out10_29 ) , .A4( u0_u10_u5_n129 ) , .A3( u0_u10_u5_n130 ) , .A2( u0_u10_u5_n168 ) , .A1( u0_u10_u5_n196 ) );
  AOI221_X1 u0_u10_u5_U93 (.A( u0_u10_u5_n128 ) , .ZN( u0_u10_u5_n129 ) , .C2( u0_u10_u5_n132 ) , .B2( u0_u10_u5_n159 ) , .B1( u0_u10_u5_n176 ) , .C1( u0_u10_u5_n184 ) );
  AOI222_X1 u0_u10_u5_U94 (.ZN( u0_u10_u5_n130 ) , .A2( u0_u10_u5_n146 ) , .B1( u0_u10_u5_n147 ) , .C2( u0_u10_u5_n175 ) , .B2( u0_u10_u5_n179 ) , .A1( u0_u10_u5_n188 ) , .C1( u0_u10_u5_n194 ) );
  NAND4_X1 u0_u10_u5_U95 (.ZN( u0_out10_19 ) , .A4( u0_u10_u5_n166 ) , .A3( u0_u10_u5_n167 ) , .A2( u0_u10_u5_n168 ) , .A1( u0_u10_u5_n169 ) );
  AOI22_X1 u0_u10_u5_U96 (.B2( u0_u10_u5_n145 ) , .A2( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n167 ) , .B1( u0_u10_u5_n182 ) , .A1( u0_u10_u5_n189 ) );
  NOR4_X1 u0_u10_u5_U97 (.A4( u0_u10_u5_n162 ) , .A3( u0_u10_u5_n163 ) , .A2( u0_u10_u5_n164 ) , .A1( u0_u10_u5_n165 ) , .ZN( u0_u10_u5_n166 ) );
  NAND4_X1 u0_u10_u5_U98 (.ZN( u0_out10_11 ) , .A4( u0_u10_u5_n143 ) , .A3( u0_u10_u5_n144 ) , .A2( u0_u10_u5_n169 ) , .A1( u0_u10_u5_n196 ) );
  AOI22_X1 u0_u10_u5_U99 (.A2( u0_u10_u5_n132 ) , .ZN( u0_u10_u5_n144 ) , .B2( u0_u10_u5_n145 ) , .B1( u0_u10_u5_n184 ) , .A1( u0_u10_u5_n194 ) );
  AOI22_X1 u0_u10_u6_U10 (.A2( u0_u10_u6_n151 ) , .B2( u0_u10_u6_n161 ) , .A1( u0_u10_u6_n167 ) , .B1( u0_u10_u6_n170 ) , .ZN( u0_u10_u6_n89 ) );
  AOI21_X1 u0_u10_u6_U11 (.B1( u0_u10_u6_n107 ) , .B2( u0_u10_u6_n132 ) , .A( u0_u10_u6_n158 ) , .ZN( u0_u10_u6_n88 ) );
  AOI21_X1 u0_u10_u6_U12 (.B2( u0_u10_u6_n147 ) , .B1( u0_u10_u6_n148 ) , .ZN( u0_u10_u6_n149 ) , .A( u0_u10_u6_n158 ) );
  AOI21_X1 u0_u10_u6_U13 (.ZN( u0_u10_u6_n106 ) , .A( u0_u10_u6_n142 ) , .B2( u0_u10_u6_n159 ) , .B1( u0_u10_u6_n164 ) );
  INV_X1 u0_u10_u6_U14 (.A( u0_u10_u6_n155 ) , .ZN( u0_u10_u6_n161 ) );
  INV_X1 u0_u10_u6_U15 (.A( u0_u10_u6_n128 ) , .ZN( u0_u10_u6_n164 ) );
  NAND2_X1 u0_u10_u6_U16 (.ZN( u0_u10_u6_n110 ) , .A1( u0_u10_u6_n122 ) , .A2( u0_u10_u6_n129 ) );
  NAND2_X1 u0_u10_u6_U17 (.ZN( u0_u10_u6_n124 ) , .A2( u0_u10_u6_n146 ) , .A1( u0_u10_u6_n148 ) );
  INV_X1 u0_u10_u6_U18 (.A( u0_u10_u6_n132 ) , .ZN( u0_u10_u6_n171 ) );
  AND2_X1 u0_u10_u6_U19 (.A1( u0_u10_u6_n100 ) , .ZN( u0_u10_u6_n130 ) , .A2( u0_u10_u6_n147 ) );
  INV_X1 u0_u10_u6_U20 (.A( u0_u10_u6_n127 ) , .ZN( u0_u10_u6_n173 ) );
  INV_X1 u0_u10_u6_U21 (.A( u0_u10_u6_n121 ) , .ZN( u0_u10_u6_n167 ) );
  INV_X1 u0_u10_u6_U22 (.A( u0_u10_u6_n100 ) , .ZN( u0_u10_u6_n169 ) );
  INV_X1 u0_u10_u6_U23 (.A( u0_u10_u6_n123 ) , .ZN( u0_u10_u6_n170 ) );
  INV_X1 u0_u10_u6_U24 (.A( u0_u10_u6_n113 ) , .ZN( u0_u10_u6_n168 ) );
  AND2_X1 u0_u10_u6_U25 (.A1( u0_u10_u6_n107 ) , .A2( u0_u10_u6_n119 ) , .ZN( u0_u10_u6_n133 ) );
  AND2_X1 u0_u10_u6_U26 (.A2( u0_u10_u6_n121 ) , .A1( u0_u10_u6_n122 ) , .ZN( u0_u10_u6_n131 ) );
  AND3_X1 u0_u10_u6_U27 (.ZN( u0_u10_u6_n120 ) , .A2( u0_u10_u6_n127 ) , .A1( u0_u10_u6_n132 ) , .A3( u0_u10_u6_n145 ) );
  INV_X1 u0_u10_u6_U28 (.A( u0_u10_u6_n146 ) , .ZN( u0_u10_u6_n163 ) );
  AOI222_X1 u0_u10_u6_U29 (.ZN( u0_u10_u6_n114 ) , .A1( u0_u10_u6_n118 ) , .A2( u0_u10_u6_n126 ) , .B2( u0_u10_u6_n151 ) , .C2( u0_u10_u6_n159 ) , .C1( u0_u10_u6_n168 ) , .B1( u0_u10_u6_n169 ) );
  INV_X1 u0_u10_u6_U3 (.A( u0_u10_u6_n110 ) , .ZN( u0_u10_u6_n166 ) );
  NOR2_X1 u0_u10_u6_U30 (.A1( u0_u10_u6_n162 ) , .A2( u0_u10_u6_n165 ) , .ZN( u0_u10_u6_n98 ) );
  AOI211_X1 u0_u10_u6_U31 (.B( u0_u10_u6_n134 ) , .A( u0_u10_u6_n135 ) , .C1( u0_u10_u6_n136 ) , .ZN( u0_u10_u6_n137 ) , .C2( u0_u10_u6_n151 ) );
  NAND4_X1 u0_u10_u6_U32 (.A4( u0_u10_u6_n127 ) , .A3( u0_u10_u6_n128 ) , .A2( u0_u10_u6_n129 ) , .A1( u0_u10_u6_n130 ) , .ZN( u0_u10_u6_n136 ) );
  AOI21_X1 u0_u10_u6_U33 (.B2( u0_u10_u6_n132 ) , .B1( u0_u10_u6_n133 ) , .ZN( u0_u10_u6_n134 ) , .A( u0_u10_u6_n158 ) );
  AOI21_X1 u0_u10_u6_U34 (.B1( u0_u10_u6_n131 ) , .ZN( u0_u10_u6_n135 ) , .A( u0_u10_u6_n144 ) , .B2( u0_u10_u6_n146 ) );
  NAND2_X1 u0_u10_u6_U35 (.A1( u0_u10_u6_n144 ) , .ZN( u0_u10_u6_n151 ) , .A2( u0_u10_u6_n158 ) );
  NAND2_X1 u0_u10_u6_U36 (.ZN( u0_u10_u6_n132 ) , .A1( u0_u10_u6_n91 ) , .A2( u0_u10_u6_n97 ) );
  AOI22_X1 u0_u10_u6_U37 (.B2( u0_u10_u6_n110 ) , .B1( u0_u10_u6_n111 ) , .A1( u0_u10_u6_n112 ) , .ZN( u0_u10_u6_n115 ) , .A2( u0_u10_u6_n161 ) );
  NAND4_X1 u0_u10_u6_U38 (.A3( u0_u10_u6_n109 ) , .ZN( u0_u10_u6_n112 ) , .A4( u0_u10_u6_n132 ) , .A2( u0_u10_u6_n147 ) , .A1( u0_u10_u6_n166 ) );
  NOR2_X1 u0_u10_u6_U39 (.ZN( u0_u10_u6_n109 ) , .A1( u0_u10_u6_n170 ) , .A2( u0_u10_u6_n173 ) );
  INV_X1 u0_u10_u6_U4 (.A( u0_u10_u6_n142 ) , .ZN( u0_u10_u6_n174 ) );
  NOR2_X1 u0_u10_u6_U40 (.A2( u0_u10_u6_n126 ) , .ZN( u0_u10_u6_n155 ) , .A1( u0_u10_u6_n160 ) );
  NAND2_X1 u0_u10_u6_U41 (.ZN( u0_u10_u6_n146 ) , .A2( u0_u10_u6_n94 ) , .A1( u0_u10_u6_n99 ) );
  AOI21_X1 u0_u10_u6_U42 (.A( u0_u10_u6_n144 ) , .B2( u0_u10_u6_n145 ) , .B1( u0_u10_u6_n146 ) , .ZN( u0_u10_u6_n150 ) );
  INV_X1 u0_u10_u6_U43 (.A( u0_u10_u6_n111 ) , .ZN( u0_u10_u6_n158 ) );
  NAND2_X1 u0_u10_u6_U44 (.ZN( u0_u10_u6_n127 ) , .A1( u0_u10_u6_n91 ) , .A2( u0_u10_u6_n92 ) );
  NAND2_X1 u0_u10_u6_U45 (.ZN( u0_u10_u6_n129 ) , .A2( u0_u10_u6_n95 ) , .A1( u0_u10_u6_n96 ) );
  INV_X1 u0_u10_u6_U46 (.A( u0_u10_u6_n144 ) , .ZN( u0_u10_u6_n159 ) );
  NAND2_X1 u0_u10_u6_U47 (.ZN( u0_u10_u6_n145 ) , .A2( u0_u10_u6_n97 ) , .A1( u0_u10_u6_n98 ) );
  NAND2_X1 u0_u10_u6_U48 (.ZN( u0_u10_u6_n148 ) , .A2( u0_u10_u6_n92 ) , .A1( u0_u10_u6_n94 ) );
  NAND2_X1 u0_u10_u6_U49 (.ZN( u0_u10_u6_n108 ) , .A2( u0_u10_u6_n139 ) , .A1( u0_u10_u6_n144 ) );
  NAND2_X1 u0_u10_u6_U5 (.A2( u0_u10_u6_n143 ) , .ZN( u0_u10_u6_n152 ) , .A1( u0_u10_u6_n166 ) );
  NAND2_X1 u0_u10_u6_U50 (.ZN( u0_u10_u6_n121 ) , .A2( u0_u10_u6_n95 ) , .A1( u0_u10_u6_n97 ) );
  NAND2_X1 u0_u10_u6_U51 (.ZN( u0_u10_u6_n107 ) , .A2( u0_u10_u6_n92 ) , .A1( u0_u10_u6_n95 ) );
  AND2_X1 u0_u10_u6_U52 (.ZN( u0_u10_u6_n118 ) , .A2( u0_u10_u6_n91 ) , .A1( u0_u10_u6_n99 ) );
  NAND2_X1 u0_u10_u6_U53 (.ZN( u0_u10_u6_n147 ) , .A2( u0_u10_u6_n98 ) , .A1( u0_u10_u6_n99 ) );
  NAND2_X1 u0_u10_u6_U54 (.ZN( u0_u10_u6_n128 ) , .A1( u0_u10_u6_n94 ) , .A2( u0_u10_u6_n96 ) );
  NAND2_X1 u0_u10_u6_U55 (.ZN( u0_u10_u6_n119 ) , .A2( u0_u10_u6_n95 ) , .A1( u0_u10_u6_n99 ) );
  NAND2_X1 u0_u10_u6_U56 (.ZN( u0_u10_u6_n123 ) , .A2( u0_u10_u6_n91 ) , .A1( u0_u10_u6_n96 ) );
  NAND2_X1 u0_u10_u6_U57 (.ZN( u0_u10_u6_n100 ) , .A2( u0_u10_u6_n92 ) , .A1( u0_u10_u6_n98 ) );
  NAND2_X1 u0_u10_u6_U58 (.ZN( u0_u10_u6_n122 ) , .A1( u0_u10_u6_n94 ) , .A2( u0_u10_u6_n97 ) );
  INV_X1 u0_u10_u6_U59 (.A( u0_u10_u6_n139 ) , .ZN( u0_u10_u6_n160 ) );
  AOI22_X1 u0_u10_u6_U6 (.B2( u0_u10_u6_n101 ) , .A1( u0_u10_u6_n102 ) , .ZN( u0_u10_u6_n103 ) , .B1( u0_u10_u6_n160 ) , .A2( u0_u10_u6_n161 ) );
  NAND2_X1 u0_u10_u6_U60 (.ZN( u0_u10_u6_n113 ) , .A1( u0_u10_u6_n96 ) , .A2( u0_u10_u6_n98 ) );
  NOR2_X1 u0_u10_u6_U61 (.A2( u0_u10_X_40 ) , .A1( u0_u10_X_41 ) , .ZN( u0_u10_u6_n126 ) );
  NOR2_X1 u0_u10_u6_U62 (.A2( u0_u10_X_39 ) , .A1( u0_u10_X_42 ) , .ZN( u0_u10_u6_n92 ) );
  NOR2_X1 u0_u10_u6_U63 (.A2( u0_u10_X_39 ) , .A1( u0_u10_u6_n156 ) , .ZN( u0_u10_u6_n97 ) );
  NOR2_X1 u0_u10_u6_U64 (.A2( u0_u10_X_38 ) , .A1( u0_u10_u6_n165 ) , .ZN( u0_u10_u6_n95 ) );
  NOR2_X1 u0_u10_u6_U65 (.A2( u0_u10_X_41 ) , .ZN( u0_u10_u6_n111 ) , .A1( u0_u10_u6_n157 ) );
  NOR2_X1 u0_u10_u6_U66 (.A2( u0_u10_X_37 ) , .A1( u0_u10_u6_n162 ) , .ZN( u0_u10_u6_n94 ) );
  NOR2_X1 u0_u10_u6_U67 (.A2( u0_u10_X_37 ) , .A1( u0_u10_X_38 ) , .ZN( u0_u10_u6_n91 ) );
  NAND2_X1 u0_u10_u6_U68 (.A1( u0_u10_X_41 ) , .ZN( u0_u10_u6_n144 ) , .A2( u0_u10_u6_n157 ) );
  NAND2_X1 u0_u10_u6_U69 (.A2( u0_u10_X_40 ) , .A1( u0_u10_X_41 ) , .ZN( u0_u10_u6_n139 ) );
  NOR2_X1 u0_u10_u6_U7 (.A1( u0_u10_u6_n118 ) , .ZN( u0_u10_u6_n143 ) , .A2( u0_u10_u6_n168 ) );
  AND2_X1 u0_u10_u6_U70 (.A1( u0_u10_X_39 ) , .A2( u0_u10_u6_n156 ) , .ZN( u0_u10_u6_n96 ) );
  AND2_X1 u0_u10_u6_U71 (.A1( u0_u10_X_39 ) , .A2( u0_u10_X_42 ) , .ZN( u0_u10_u6_n99 ) );
  INV_X1 u0_u10_u6_U72 (.A( u0_u10_X_40 ) , .ZN( u0_u10_u6_n157 ) );
  INV_X1 u0_u10_u6_U73 (.A( u0_u10_X_37 ) , .ZN( u0_u10_u6_n165 ) );
  INV_X1 u0_u10_u6_U74 (.A( u0_u10_X_38 ) , .ZN( u0_u10_u6_n162 ) );
  INV_X1 u0_u10_u6_U75 (.A( u0_u10_X_42 ) , .ZN( u0_u10_u6_n156 ) );
  NAND4_X1 u0_u10_u6_U76 (.ZN( u0_out10_32 ) , .A4( u0_u10_u6_n103 ) , .A3( u0_u10_u6_n104 ) , .A2( u0_u10_u6_n105 ) , .A1( u0_u10_u6_n106 ) );
  AOI22_X1 u0_u10_u6_U77 (.ZN( u0_u10_u6_n105 ) , .A2( u0_u10_u6_n108 ) , .A1( u0_u10_u6_n118 ) , .B2( u0_u10_u6_n126 ) , .B1( u0_u10_u6_n171 ) );
  AOI22_X1 u0_u10_u6_U78 (.ZN( u0_u10_u6_n104 ) , .A1( u0_u10_u6_n111 ) , .B1( u0_u10_u6_n124 ) , .B2( u0_u10_u6_n151 ) , .A2( u0_u10_u6_n93 ) );
  NAND4_X1 u0_u10_u6_U79 (.ZN( u0_out10_12 ) , .A4( u0_u10_u6_n114 ) , .A3( u0_u10_u6_n115 ) , .A2( u0_u10_u6_n116 ) , .A1( u0_u10_u6_n117 ) );
  INV_X1 u0_u10_u6_U8 (.ZN( u0_u10_u6_n172 ) , .A( u0_u10_u6_n88 ) );
  OAI22_X1 u0_u10_u6_U80 (.B2( u0_u10_u6_n111 ) , .ZN( u0_u10_u6_n116 ) , .B1( u0_u10_u6_n126 ) , .A2( u0_u10_u6_n164 ) , .A1( u0_u10_u6_n167 ) );
  OAI21_X1 u0_u10_u6_U81 (.A( u0_u10_u6_n108 ) , .ZN( u0_u10_u6_n117 ) , .B2( u0_u10_u6_n141 ) , .B1( u0_u10_u6_n163 ) );
  OAI211_X1 u0_u10_u6_U82 (.ZN( u0_out10_7 ) , .B( u0_u10_u6_n153 ) , .C2( u0_u10_u6_n154 ) , .C1( u0_u10_u6_n155 ) , .A( u0_u10_u6_n174 ) );
  NOR3_X1 u0_u10_u6_U83 (.A1( u0_u10_u6_n141 ) , .ZN( u0_u10_u6_n154 ) , .A3( u0_u10_u6_n164 ) , .A2( u0_u10_u6_n171 ) );
  AOI211_X1 u0_u10_u6_U84 (.B( u0_u10_u6_n149 ) , .A( u0_u10_u6_n150 ) , .C2( u0_u10_u6_n151 ) , .C1( u0_u10_u6_n152 ) , .ZN( u0_u10_u6_n153 ) );
  OAI211_X1 u0_u10_u6_U85 (.ZN( u0_out10_22 ) , .B( u0_u10_u6_n137 ) , .A( u0_u10_u6_n138 ) , .C2( u0_u10_u6_n139 ) , .C1( u0_u10_u6_n140 ) );
  AOI22_X1 u0_u10_u6_U86 (.B1( u0_u10_u6_n124 ) , .A2( u0_u10_u6_n125 ) , .A1( u0_u10_u6_n126 ) , .ZN( u0_u10_u6_n138 ) , .B2( u0_u10_u6_n161 ) );
  AND4_X1 u0_u10_u6_U87 (.A3( u0_u10_u6_n119 ) , .A1( u0_u10_u6_n120 ) , .A4( u0_u10_u6_n129 ) , .ZN( u0_u10_u6_n140 ) , .A2( u0_u10_u6_n143 ) );
  NAND3_X1 u0_u10_u6_U88 (.A2( u0_u10_u6_n123 ) , .ZN( u0_u10_u6_n125 ) , .A1( u0_u10_u6_n130 ) , .A3( u0_u10_u6_n131 ) );
  NAND3_X1 u0_u10_u6_U89 (.A3( u0_u10_u6_n133 ) , .ZN( u0_u10_u6_n141 ) , .A1( u0_u10_u6_n145 ) , .A2( u0_u10_u6_n148 ) );
  OAI21_X1 u0_u10_u6_U9 (.A( u0_u10_u6_n159 ) , .B1( u0_u10_u6_n169 ) , .B2( u0_u10_u6_n173 ) , .ZN( u0_u10_u6_n90 ) );
  NAND3_X1 u0_u10_u6_U90 (.ZN( u0_u10_u6_n101 ) , .A3( u0_u10_u6_n107 ) , .A2( u0_u10_u6_n121 ) , .A1( u0_u10_u6_n127 ) );
  NAND3_X1 u0_u10_u6_U91 (.ZN( u0_u10_u6_n102 ) , .A3( u0_u10_u6_n130 ) , .A2( u0_u10_u6_n145 ) , .A1( u0_u10_u6_n166 ) );
  NAND3_X1 u0_u10_u6_U92 (.A3( u0_u10_u6_n113 ) , .A1( u0_u10_u6_n119 ) , .A2( u0_u10_u6_n123 ) , .ZN( u0_u10_u6_n93 ) );
  NAND3_X1 u0_u10_u6_U93 (.ZN( u0_u10_u6_n142 ) , .A2( u0_u10_u6_n172 ) , .A3( u0_u10_u6_n89 ) , .A1( u0_u10_u6_n90 ) );
  AND3_X1 u0_u10_u7_U10 (.A3( u0_u10_u7_n110 ) , .A2( u0_u10_u7_n127 ) , .A1( u0_u10_u7_n132 ) , .ZN( u0_u10_u7_n92 ) );
  OAI21_X1 u0_u10_u7_U11 (.A( u0_u10_u7_n161 ) , .B1( u0_u10_u7_n168 ) , .B2( u0_u10_u7_n173 ) , .ZN( u0_u10_u7_n91 ) );
  AOI211_X1 u0_u10_u7_U12 (.A( u0_u10_u7_n117 ) , .ZN( u0_u10_u7_n118 ) , .C2( u0_u10_u7_n126 ) , .C1( u0_u10_u7_n177 ) , .B( u0_u10_u7_n180 ) );
  OAI22_X1 u0_u10_u7_U13 (.B1( u0_u10_u7_n115 ) , .ZN( u0_u10_u7_n117 ) , .A2( u0_u10_u7_n133 ) , .A1( u0_u10_u7_n137 ) , .B2( u0_u10_u7_n162 ) );
  INV_X1 u0_u10_u7_U14 (.A( u0_u10_u7_n116 ) , .ZN( u0_u10_u7_n180 ) );
  NOR3_X1 u0_u10_u7_U15 (.ZN( u0_u10_u7_n115 ) , .A3( u0_u10_u7_n145 ) , .A2( u0_u10_u7_n168 ) , .A1( u0_u10_u7_n169 ) );
  OAI211_X1 u0_u10_u7_U16 (.B( u0_u10_u7_n122 ) , .A( u0_u10_u7_n123 ) , .C2( u0_u10_u7_n124 ) , .ZN( u0_u10_u7_n154 ) , .C1( u0_u10_u7_n162 ) );
  AOI222_X1 u0_u10_u7_U17 (.ZN( u0_u10_u7_n122 ) , .C2( u0_u10_u7_n126 ) , .C1( u0_u10_u7_n145 ) , .B1( u0_u10_u7_n161 ) , .A2( u0_u10_u7_n165 ) , .B2( u0_u10_u7_n170 ) , .A1( u0_u10_u7_n176 ) );
  INV_X1 u0_u10_u7_U18 (.A( u0_u10_u7_n133 ) , .ZN( u0_u10_u7_n176 ) );
  NOR3_X1 u0_u10_u7_U19 (.A2( u0_u10_u7_n134 ) , .A1( u0_u10_u7_n135 ) , .ZN( u0_u10_u7_n136 ) , .A3( u0_u10_u7_n171 ) );
  NOR2_X1 u0_u10_u7_U20 (.A1( u0_u10_u7_n130 ) , .A2( u0_u10_u7_n134 ) , .ZN( u0_u10_u7_n153 ) );
  INV_X1 u0_u10_u7_U21 (.A( u0_u10_u7_n101 ) , .ZN( u0_u10_u7_n165 ) );
  NOR2_X1 u0_u10_u7_U22 (.ZN( u0_u10_u7_n111 ) , .A2( u0_u10_u7_n134 ) , .A1( u0_u10_u7_n169 ) );
  AOI21_X1 u0_u10_u7_U23 (.ZN( u0_u10_u7_n104 ) , .B2( u0_u10_u7_n112 ) , .B1( u0_u10_u7_n127 ) , .A( u0_u10_u7_n164 ) );
  AOI21_X1 u0_u10_u7_U24 (.ZN( u0_u10_u7_n106 ) , .B1( u0_u10_u7_n133 ) , .B2( u0_u10_u7_n146 ) , .A( u0_u10_u7_n162 ) );
  AOI21_X1 u0_u10_u7_U25 (.A( u0_u10_u7_n101 ) , .ZN( u0_u10_u7_n107 ) , .B2( u0_u10_u7_n128 ) , .B1( u0_u10_u7_n175 ) );
  INV_X1 u0_u10_u7_U26 (.A( u0_u10_u7_n138 ) , .ZN( u0_u10_u7_n171 ) );
  INV_X1 u0_u10_u7_U27 (.A( u0_u10_u7_n131 ) , .ZN( u0_u10_u7_n177 ) );
  INV_X1 u0_u10_u7_U28 (.A( u0_u10_u7_n110 ) , .ZN( u0_u10_u7_n174 ) );
  NAND2_X1 u0_u10_u7_U29 (.A1( u0_u10_u7_n129 ) , .A2( u0_u10_u7_n132 ) , .ZN( u0_u10_u7_n149 ) );
  OAI21_X1 u0_u10_u7_U3 (.ZN( u0_u10_u7_n159 ) , .A( u0_u10_u7_n165 ) , .B2( u0_u10_u7_n171 ) , .B1( u0_u10_u7_n174 ) );
  NAND2_X1 u0_u10_u7_U30 (.A1( u0_u10_u7_n113 ) , .A2( u0_u10_u7_n124 ) , .ZN( u0_u10_u7_n130 ) );
  INV_X1 u0_u10_u7_U31 (.A( u0_u10_u7_n112 ) , .ZN( u0_u10_u7_n173 ) );
  INV_X1 u0_u10_u7_U32 (.A( u0_u10_u7_n128 ) , .ZN( u0_u10_u7_n168 ) );
  INV_X1 u0_u10_u7_U33 (.A( u0_u10_u7_n148 ) , .ZN( u0_u10_u7_n169 ) );
  INV_X1 u0_u10_u7_U34 (.A( u0_u10_u7_n127 ) , .ZN( u0_u10_u7_n179 ) );
  NOR2_X1 u0_u10_u7_U35 (.ZN( u0_u10_u7_n101 ) , .A2( u0_u10_u7_n150 ) , .A1( u0_u10_u7_n156 ) );
  AOI211_X1 u0_u10_u7_U36 (.B( u0_u10_u7_n154 ) , .A( u0_u10_u7_n155 ) , .C1( u0_u10_u7_n156 ) , .ZN( u0_u10_u7_n157 ) , .C2( u0_u10_u7_n172 ) );
  INV_X1 u0_u10_u7_U37 (.A( u0_u10_u7_n153 ) , .ZN( u0_u10_u7_n172 ) );
  AOI211_X1 u0_u10_u7_U38 (.B( u0_u10_u7_n139 ) , .A( u0_u10_u7_n140 ) , .C2( u0_u10_u7_n141 ) , .ZN( u0_u10_u7_n142 ) , .C1( u0_u10_u7_n156 ) );
  NAND4_X1 u0_u10_u7_U39 (.A3( u0_u10_u7_n127 ) , .A2( u0_u10_u7_n128 ) , .A1( u0_u10_u7_n129 ) , .ZN( u0_u10_u7_n141 ) , .A4( u0_u10_u7_n147 ) );
  INV_X1 u0_u10_u7_U4 (.A( u0_u10_u7_n111 ) , .ZN( u0_u10_u7_n170 ) );
  AOI21_X1 u0_u10_u7_U40 (.A( u0_u10_u7_n137 ) , .B1( u0_u10_u7_n138 ) , .ZN( u0_u10_u7_n139 ) , .B2( u0_u10_u7_n146 ) );
  OAI22_X1 u0_u10_u7_U41 (.B1( u0_u10_u7_n136 ) , .ZN( u0_u10_u7_n140 ) , .A1( u0_u10_u7_n153 ) , .B2( u0_u10_u7_n162 ) , .A2( u0_u10_u7_n164 ) );
  AOI21_X1 u0_u10_u7_U42 (.ZN( u0_u10_u7_n123 ) , .B1( u0_u10_u7_n165 ) , .B2( u0_u10_u7_n177 ) , .A( u0_u10_u7_n97 ) );
  AOI21_X1 u0_u10_u7_U43 (.B2( u0_u10_u7_n113 ) , .B1( u0_u10_u7_n124 ) , .A( u0_u10_u7_n125 ) , .ZN( u0_u10_u7_n97 ) );
  INV_X1 u0_u10_u7_U44 (.A( u0_u10_u7_n125 ) , .ZN( u0_u10_u7_n161 ) );
  INV_X1 u0_u10_u7_U45 (.A( u0_u10_u7_n152 ) , .ZN( u0_u10_u7_n162 ) );
  AOI22_X1 u0_u10_u7_U46 (.A2( u0_u10_u7_n114 ) , .ZN( u0_u10_u7_n119 ) , .B1( u0_u10_u7_n130 ) , .A1( u0_u10_u7_n156 ) , .B2( u0_u10_u7_n165 ) );
  NAND2_X1 u0_u10_u7_U47 (.A2( u0_u10_u7_n112 ) , .ZN( u0_u10_u7_n114 ) , .A1( u0_u10_u7_n175 ) );
  AND2_X1 u0_u10_u7_U48 (.ZN( u0_u10_u7_n145 ) , .A2( u0_u10_u7_n98 ) , .A1( u0_u10_u7_n99 ) );
  NOR2_X1 u0_u10_u7_U49 (.ZN( u0_u10_u7_n137 ) , .A1( u0_u10_u7_n150 ) , .A2( u0_u10_u7_n161 ) );
  INV_X1 u0_u10_u7_U5 (.A( u0_u10_u7_n149 ) , .ZN( u0_u10_u7_n175 ) );
  AOI21_X1 u0_u10_u7_U50 (.ZN( u0_u10_u7_n105 ) , .B2( u0_u10_u7_n110 ) , .A( u0_u10_u7_n125 ) , .B1( u0_u10_u7_n147 ) );
  NAND2_X1 u0_u10_u7_U51 (.ZN( u0_u10_u7_n146 ) , .A1( u0_u10_u7_n95 ) , .A2( u0_u10_u7_n98 ) );
  NAND2_X1 u0_u10_u7_U52 (.A2( u0_u10_u7_n103 ) , .ZN( u0_u10_u7_n147 ) , .A1( u0_u10_u7_n93 ) );
  NAND2_X1 u0_u10_u7_U53 (.A1( u0_u10_u7_n103 ) , .ZN( u0_u10_u7_n127 ) , .A2( u0_u10_u7_n99 ) );
  OR2_X1 u0_u10_u7_U54 (.ZN( u0_u10_u7_n126 ) , .A2( u0_u10_u7_n152 ) , .A1( u0_u10_u7_n156 ) );
  NAND2_X1 u0_u10_u7_U55 (.A2( u0_u10_u7_n102 ) , .A1( u0_u10_u7_n103 ) , .ZN( u0_u10_u7_n133 ) );
  NAND2_X1 u0_u10_u7_U56 (.ZN( u0_u10_u7_n112 ) , .A2( u0_u10_u7_n96 ) , .A1( u0_u10_u7_n99 ) );
  NAND2_X1 u0_u10_u7_U57 (.A2( u0_u10_u7_n102 ) , .ZN( u0_u10_u7_n128 ) , .A1( u0_u10_u7_n98 ) );
  NAND2_X1 u0_u10_u7_U58 (.A1( u0_u10_u7_n100 ) , .ZN( u0_u10_u7_n113 ) , .A2( u0_u10_u7_n93 ) );
  NAND2_X1 u0_u10_u7_U59 (.A2( u0_u10_u7_n102 ) , .ZN( u0_u10_u7_n124 ) , .A1( u0_u10_u7_n96 ) );
  INV_X1 u0_u10_u7_U6 (.A( u0_u10_u7_n154 ) , .ZN( u0_u10_u7_n178 ) );
  NAND2_X1 u0_u10_u7_U60 (.ZN( u0_u10_u7_n110 ) , .A1( u0_u10_u7_n95 ) , .A2( u0_u10_u7_n96 ) );
  INV_X1 u0_u10_u7_U61 (.A( u0_u10_u7_n150 ) , .ZN( u0_u10_u7_n164 ) );
  AND2_X1 u0_u10_u7_U62 (.ZN( u0_u10_u7_n134 ) , .A1( u0_u10_u7_n93 ) , .A2( u0_u10_u7_n98 ) );
  NAND2_X1 u0_u10_u7_U63 (.A1( u0_u10_u7_n100 ) , .A2( u0_u10_u7_n102 ) , .ZN( u0_u10_u7_n129 ) );
  NAND2_X1 u0_u10_u7_U64 (.A2( u0_u10_u7_n103 ) , .ZN( u0_u10_u7_n131 ) , .A1( u0_u10_u7_n95 ) );
  NAND2_X1 u0_u10_u7_U65 (.A1( u0_u10_u7_n100 ) , .ZN( u0_u10_u7_n138 ) , .A2( u0_u10_u7_n99 ) );
  NAND2_X1 u0_u10_u7_U66 (.ZN( u0_u10_u7_n132 ) , .A1( u0_u10_u7_n93 ) , .A2( u0_u10_u7_n96 ) );
  NAND2_X1 u0_u10_u7_U67 (.A1( u0_u10_u7_n100 ) , .ZN( u0_u10_u7_n148 ) , .A2( u0_u10_u7_n95 ) );
  NOR2_X1 u0_u10_u7_U68 (.A2( u0_u10_X_47 ) , .ZN( u0_u10_u7_n150 ) , .A1( u0_u10_u7_n163 ) );
  NOR2_X1 u0_u10_u7_U69 (.A2( u0_u10_X_43 ) , .A1( u0_u10_X_44 ) , .ZN( u0_u10_u7_n103 ) );
  AOI211_X1 u0_u10_u7_U7 (.ZN( u0_u10_u7_n116 ) , .A( u0_u10_u7_n155 ) , .C1( u0_u10_u7_n161 ) , .C2( u0_u10_u7_n171 ) , .B( u0_u10_u7_n94 ) );
  NOR2_X1 u0_u10_u7_U70 (.A2( u0_u10_X_48 ) , .A1( u0_u10_u7_n166 ) , .ZN( u0_u10_u7_n95 ) );
  NOR2_X1 u0_u10_u7_U71 (.A2( u0_u10_X_45 ) , .A1( u0_u10_X_48 ) , .ZN( u0_u10_u7_n99 ) );
  NOR2_X1 u0_u10_u7_U72 (.A2( u0_u10_X_44 ) , .A1( u0_u10_u7_n167 ) , .ZN( u0_u10_u7_n98 ) );
  NOR2_X1 u0_u10_u7_U73 (.A2( u0_u10_X_46 ) , .A1( u0_u10_X_47 ) , .ZN( u0_u10_u7_n152 ) );
  AND2_X1 u0_u10_u7_U74 (.A1( u0_u10_X_47 ) , .ZN( u0_u10_u7_n156 ) , .A2( u0_u10_u7_n163 ) );
  NAND2_X1 u0_u10_u7_U75 (.A2( u0_u10_X_46 ) , .A1( u0_u10_X_47 ) , .ZN( u0_u10_u7_n125 ) );
  AND2_X1 u0_u10_u7_U76 (.A2( u0_u10_X_45 ) , .A1( u0_u10_X_48 ) , .ZN( u0_u10_u7_n102 ) );
  AND2_X1 u0_u10_u7_U77 (.A2( u0_u10_X_43 ) , .A1( u0_u10_X_44 ) , .ZN( u0_u10_u7_n96 ) );
  AND2_X1 u0_u10_u7_U78 (.A1( u0_u10_X_44 ) , .ZN( u0_u10_u7_n100 ) , .A2( u0_u10_u7_n167 ) );
  AND2_X1 u0_u10_u7_U79 (.A1( u0_u10_X_48 ) , .A2( u0_u10_u7_n166 ) , .ZN( u0_u10_u7_n93 ) );
  OAI222_X1 u0_u10_u7_U8 (.C2( u0_u10_u7_n101 ) , .B2( u0_u10_u7_n111 ) , .A1( u0_u10_u7_n113 ) , .C1( u0_u10_u7_n146 ) , .A2( u0_u10_u7_n162 ) , .B1( u0_u10_u7_n164 ) , .ZN( u0_u10_u7_n94 ) );
  INV_X1 u0_u10_u7_U80 (.A( u0_u10_X_46 ) , .ZN( u0_u10_u7_n163 ) );
  INV_X1 u0_u10_u7_U81 (.A( u0_u10_X_43 ) , .ZN( u0_u10_u7_n167 ) );
  INV_X1 u0_u10_u7_U82 (.A( u0_u10_X_45 ) , .ZN( u0_u10_u7_n166 ) );
  NAND4_X1 u0_u10_u7_U83 (.ZN( u0_out10_27 ) , .A4( u0_u10_u7_n118 ) , .A3( u0_u10_u7_n119 ) , .A2( u0_u10_u7_n120 ) , .A1( u0_u10_u7_n121 ) );
  OAI21_X1 u0_u10_u7_U84 (.ZN( u0_u10_u7_n121 ) , .B2( u0_u10_u7_n145 ) , .A( u0_u10_u7_n150 ) , .B1( u0_u10_u7_n174 ) );
  OAI21_X1 u0_u10_u7_U85 (.ZN( u0_u10_u7_n120 ) , .A( u0_u10_u7_n161 ) , .B2( u0_u10_u7_n170 ) , .B1( u0_u10_u7_n179 ) );
  NAND4_X1 u0_u10_u7_U86 (.ZN( u0_out10_21 ) , .A4( u0_u10_u7_n157 ) , .A3( u0_u10_u7_n158 ) , .A2( u0_u10_u7_n159 ) , .A1( u0_u10_u7_n160 ) );
  OAI21_X1 u0_u10_u7_U87 (.B1( u0_u10_u7_n145 ) , .ZN( u0_u10_u7_n160 ) , .A( u0_u10_u7_n161 ) , .B2( u0_u10_u7_n177 ) );
  AOI22_X1 u0_u10_u7_U88 (.B2( u0_u10_u7_n149 ) , .B1( u0_u10_u7_n150 ) , .A2( u0_u10_u7_n151 ) , .A1( u0_u10_u7_n152 ) , .ZN( u0_u10_u7_n158 ) );
  NAND4_X1 u0_u10_u7_U89 (.ZN( u0_out10_15 ) , .A4( u0_u10_u7_n142 ) , .A3( u0_u10_u7_n143 ) , .A2( u0_u10_u7_n144 ) , .A1( u0_u10_u7_n178 ) );
  OAI221_X1 u0_u10_u7_U9 (.C1( u0_u10_u7_n101 ) , .C2( u0_u10_u7_n147 ) , .ZN( u0_u10_u7_n155 ) , .B2( u0_u10_u7_n162 ) , .A( u0_u10_u7_n91 ) , .B1( u0_u10_u7_n92 ) );
  OR2_X1 u0_u10_u7_U90 (.A2( u0_u10_u7_n125 ) , .A1( u0_u10_u7_n129 ) , .ZN( u0_u10_u7_n144 ) );
  AOI22_X1 u0_u10_u7_U91 (.A2( u0_u10_u7_n126 ) , .ZN( u0_u10_u7_n143 ) , .B2( u0_u10_u7_n165 ) , .B1( u0_u10_u7_n173 ) , .A1( u0_u10_u7_n174 ) );
  NAND4_X1 u0_u10_u7_U92 (.ZN( u0_out10_5 ) , .A4( u0_u10_u7_n108 ) , .A3( u0_u10_u7_n109 ) , .A1( u0_u10_u7_n116 ) , .A2( u0_u10_u7_n123 ) );
  AOI22_X1 u0_u10_u7_U93 (.ZN( u0_u10_u7_n109 ) , .A2( u0_u10_u7_n126 ) , .B2( u0_u10_u7_n145 ) , .B1( u0_u10_u7_n156 ) , .A1( u0_u10_u7_n171 ) );
  NOR4_X1 u0_u10_u7_U94 (.A4( u0_u10_u7_n104 ) , .A3( u0_u10_u7_n105 ) , .A2( u0_u10_u7_n106 ) , .A1( u0_u10_u7_n107 ) , .ZN( u0_u10_u7_n108 ) );
  NAND3_X1 u0_u10_u7_U95 (.A3( u0_u10_u7_n146 ) , .A2( u0_u10_u7_n147 ) , .A1( u0_u10_u7_n148 ) , .ZN( u0_u10_u7_n151 ) );
  NAND3_X1 u0_u10_u7_U96 (.A3( u0_u10_u7_n131 ) , .A2( u0_u10_u7_n132 ) , .A1( u0_u10_u7_n133 ) , .ZN( u0_u10_u7_n135 ) );
  XOR2_X1 u0_u12_U1 (.B( u0_K13_9 ) , .A( u0_R11_6 ) , .Z( u0_u12_X_9 ) );
  XOR2_X1 u0_u12_U2 (.B( u0_K13_8 ) , .A( u0_R11_5 ) , .Z( u0_u12_X_8 ) );
  XOR2_X1 u0_u12_U3 (.B( u0_K13_7 ) , .A( u0_R11_4 ) , .Z( u0_u12_X_7 ) );
  XOR2_X1 u0_u12_U33 (.B( u0_K13_24 ) , .A( u0_R11_17 ) , .Z( u0_u12_X_24 ) );
  XOR2_X1 u0_u12_U34 (.B( u0_K13_23 ) , .A( u0_R11_16 ) , .Z( u0_u12_X_23 ) );
  XOR2_X1 u0_u12_U35 (.B( u0_K13_22 ) , .A( u0_R11_15 ) , .Z( u0_u12_X_22 ) );
  XOR2_X1 u0_u12_U36 (.B( u0_K13_21 ) , .A( u0_R11_14 ) , .Z( u0_u12_X_21 ) );
  XOR2_X1 u0_u12_U37 (.B( u0_K13_20 ) , .A( u0_R11_13 ) , .Z( u0_u12_X_20 ) );
  XOR2_X1 u0_u12_U39 (.B( u0_K13_19 ) , .A( u0_R11_12 ) , .Z( u0_u12_X_19 ) );
  XOR2_X1 u0_u12_U40 (.B( u0_K13_18 ) , .A( u0_R11_13 ) , .Z( u0_u12_X_18 ) );
  XOR2_X1 u0_u12_U41 (.B( u0_K13_17 ) , .A( u0_R11_12 ) , .Z( u0_u12_X_17 ) );
  XOR2_X1 u0_u12_U42 (.B( u0_K13_16 ) , .A( u0_R11_11 ) , .Z( u0_u12_X_16 ) );
  XOR2_X1 u0_u12_U43 (.B( u0_K13_15 ) , .A( u0_R11_10 ) , .Z( u0_u12_X_15 ) );
  XOR2_X1 u0_u12_U44 (.B( u0_K13_14 ) , .A( u0_R11_9 ) , .Z( u0_u12_X_14 ) );
  XOR2_X1 u0_u12_U45 (.B( u0_K13_13 ) , .A( u0_R11_8 ) , .Z( u0_u12_X_13 ) );
  XOR2_X1 u0_u12_U46 (.B( u0_K13_12 ) , .A( u0_R11_9 ) , .Z( u0_u12_X_12 ) );
  XOR2_X1 u0_u12_U47 (.B( u0_K13_11 ) , .A( u0_R11_8 ) , .Z( u0_u12_X_11 ) );
  XOR2_X1 u0_u12_U48 (.B( u0_K13_10 ) , .A( u0_R11_7 ) , .Z( u0_u12_X_10 ) );
  NOR2_X1 u0_u12_u1_U10 (.A1( u0_u12_u1_n112 ) , .A2( u0_u12_u1_n116 ) , .ZN( u0_u12_u1_n118 ) );
  NAND3_X1 u0_u12_u1_U100 (.ZN( u0_u12_u1_n113 ) , .A1( u0_u12_u1_n120 ) , .A3( u0_u12_u1_n133 ) , .A2( u0_u12_u1_n155 ) );
  OAI21_X1 u0_u12_u1_U11 (.ZN( u0_u12_u1_n101 ) , .B1( u0_u12_u1_n141 ) , .A( u0_u12_u1_n146 ) , .B2( u0_u12_u1_n183 ) );
  AOI21_X1 u0_u12_u1_U12 (.B2( u0_u12_u1_n155 ) , .B1( u0_u12_u1_n156 ) , .ZN( u0_u12_u1_n157 ) , .A( u0_u12_u1_n174 ) );
  OR4_X1 u0_u12_u1_U13 (.A4( u0_u12_u1_n106 ) , .A3( u0_u12_u1_n107 ) , .ZN( u0_u12_u1_n108 ) , .A1( u0_u12_u1_n117 ) , .A2( u0_u12_u1_n184 ) );
  AOI21_X1 u0_u12_u1_U14 (.ZN( u0_u12_u1_n106 ) , .A( u0_u12_u1_n112 ) , .B1( u0_u12_u1_n154 ) , .B2( u0_u12_u1_n156 ) );
  INV_X1 u0_u12_u1_U15 (.A( u0_u12_u1_n101 ) , .ZN( u0_u12_u1_n184 ) );
  AOI21_X1 u0_u12_u1_U16 (.ZN( u0_u12_u1_n107 ) , .B1( u0_u12_u1_n134 ) , .B2( u0_u12_u1_n149 ) , .A( u0_u12_u1_n174 ) );
  NAND2_X1 u0_u12_u1_U17 (.ZN( u0_u12_u1_n140 ) , .A2( u0_u12_u1_n150 ) , .A1( u0_u12_u1_n155 ) );
  NAND2_X1 u0_u12_u1_U18 (.A1( u0_u12_u1_n131 ) , .ZN( u0_u12_u1_n147 ) , .A2( u0_u12_u1_n153 ) );
  INV_X1 u0_u12_u1_U19 (.A( u0_u12_u1_n139 ) , .ZN( u0_u12_u1_n174 ) );
  INV_X1 u0_u12_u1_U20 (.A( u0_u12_u1_n112 ) , .ZN( u0_u12_u1_n171 ) );
  NAND2_X1 u0_u12_u1_U21 (.ZN( u0_u12_u1_n141 ) , .A1( u0_u12_u1_n153 ) , .A2( u0_u12_u1_n156 ) );
  AND2_X1 u0_u12_u1_U22 (.A1( u0_u12_u1_n123 ) , .ZN( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n161 ) );
  NAND2_X1 u0_u12_u1_U23 (.A2( u0_u12_u1_n115 ) , .A1( u0_u12_u1_n116 ) , .ZN( u0_u12_u1_n148 ) );
  NAND2_X1 u0_u12_u1_U24 (.A2( u0_u12_u1_n133 ) , .A1( u0_u12_u1_n135 ) , .ZN( u0_u12_u1_n159 ) );
  NAND2_X1 u0_u12_u1_U25 (.A2( u0_u12_u1_n115 ) , .A1( u0_u12_u1_n120 ) , .ZN( u0_u12_u1_n132 ) );
  INV_X1 u0_u12_u1_U26 (.A( u0_u12_u1_n154 ) , .ZN( u0_u12_u1_n178 ) );
  INV_X1 u0_u12_u1_U27 (.A( u0_u12_u1_n151 ) , .ZN( u0_u12_u1_n183 ) );
  AND2_X1 u0_u12_u1_U28 (.A1( u0_u12_u1_n129 ) , .A2( u0_u12_u1_n133 ) , .ZN( u0_u12_u1_n149 ) );
  INV_X1 u0_u12_u1_U29 (.A( u0_u12_u1_n131 ) , .ZN( u0_u12_u1_n180 ) );
  INV_X1 u0_u12_u1_U3 (.A( u0_u12_u1_n159 ) , .ZN( u0_u12_u1_n182 ) );
  AOI221_X1 u0_u12_u1_U30 (.B1( u0_u12_u1_n140 ) , .ZN( u0_u12_u1_n167 ) , .B2( u0_u12_u1_n172 ) , .C2( u0_u12_u1_n175 ) , .C1( u0_u12_u1_n178 ) , .A( u0_u12_u1_n188 ) );
  INV_X1 u0_u12_u1_U31 (.ZN( u0_u12_u1_n188 ) , .A( u0_u12_u1_n97 ) );
  AOI211_X1 u0_u12_u1_U32 (.A( u0_u12_u1_n118 ) , .C1( u0_u12_u1_n132 ) , .C2( u0_u12_u1_n139 ) , .B( u0_u12_u1_n96 ) , .ZN( u0_u12_u1_n97 ) );
  AOI21_X1 u0_u12_u1_U33 (.B2( u0_u12_u1_n121 ) , .B1( u0_u12_u1_n135 ) , .A( u0_u12_u1_n152 ) , .ZN( u0_u12_u1_n96 ) );
  OAI221_X1 u0_u12_u1_U34 (.A( u0_u12_u1_n119 ) , .C2( u0_u12_u1_n129 ) , .ZN( u0_u12_u1_n138 ) , .B2( u0_u12_u1_n152 ) , .C1( u0_u12_u1_n174 ) , .B1( u0_u12_u1_n187 ) );
  INV_X1 u0_u12_u1_U35 (.A( u0_u12_u1_n148 ) , .ZN( u0_u12_u1_n187 ) );
  AOI211_X1 u0_u12_u1_U36 (.B( u0_u12_u1_n117 ) , .A( u0_u12_u1_n118 ) , .ZN( u0_u12_u1_n119 ) , .C2( u0_u12_u1_n146 ) , .C1( u0_u12_u1_n159 ) );
  NOR2_X1 u0_u12_u1_U37 (.A1( u0_u12_u1_n168 ) , .A2( u0_u12_u1_n176 ) , .ZN( u0_u12_u1_n98 ) );
  AOI211_X1 u0_u12_u1_U38 (.B( u0_u12_u1_n162 ) , .A( u0_u12_u1_n163 ) , .C2( u0_u12_u1_n164 ) , .ZN( u0_u12_u1_n165 ) , .C1( u0_u12_u1_n171 ) );
  AOI21_X1 u0_u12_u1_U39 (.A( u0_u12_u1_n160 ) , .B2( u0_u12_u1_n161 ) , .ZN( u0_u12_u1_n162 ) , .B1( u0_u12_u1_n182 ) );
  AOI221_X1 u0_u12_u1_U4 (.A( u0_u12_u1_n138 ) , .C2( u0_u12_u1_n139 ) , .C1( u0_u12_u1_n140 ) , .B2( u0_u12_u1_n141 ) , .ZN( u0_u12_u1_n142 ) , .B1( u0_u12_u1_n175 ) );
  OR2_X1 u0_u12_u1_U40 (.A2( u0_u12_u1_n157 ) , .A1( u0_u12_u1_n158 ) , .ZN( u0_u12_u1_n163 ) );
  NAND2_X1 u0_u12_u1_U41 (.A1( u0_u12_u1_n128 ) , .ZN( u0_u12_u1_n146 ) , .A2( u0_u12_u1_n160 ) );
  NAND2_X1 u0_u12_u1_U42 (.A2( u0_u12_u1_n112 ) , .ZN( u0_u12_u1_n139 ) , .A1( u0_u12_u1_n152 ) );
  NAND2_X1 u0_u12_u1_U43 (.A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n156 ) , .A2( u0_u12_u1_n99 ) );
  NOR2_X1 u0_u12_u1_U44 (.ZN( u0_u12_u1_n117 ) , .A1( u0_u12_u1_n121 ) , .A2( u0_u12_u1_n160 ) );
  OAI21_X1 u0_u12_u1_U45 (.B2( u0_u12_u1_n123 ) , .ZN( u0_u12_u1_n145 ) , .B1( u0_u12_u1_n160 ) , .A( u0_u12_u1_n185 ) );
  INV_X1 u0_u12_u1_U46 (.A( u0_u12_u1_n122 ) , .ZN( u0_u12_u1_n185 ) );
  AOI21_X1 u0_u12_u1_U47 (.B2( u0_u12_u1_n120 ) , .B1( u0_u12_u1_n121 ) , .ZN( u0_u12_u1_n122 ) , .A( u0_u12_u1_n128 ) );
  AOI21_X1 u0_u12_u1_U48 (.A( u0_u12_u1_n128 ) , .B2( u0_u12_u1_n129 ) , .ZN( u0_u12_u1_n130 ) , .B1( u0_u12_u1_n150 ) );
  NAND2_X1 u0_u12_u1_U49 (.ZN( u0_u12_u1_n112 ) , .A1( u0_u12_u1_n169 ) , .A2( u0_u12_u1_n170 ) );
  AOI211_X1 u0_u12_u1_U5 (.ZN( u0_u12_u1_n124 ) , .A( u0_u12_u1_n138 ) , .C2( u0_u12_u1_n139 ) , .B( u0_u12_u1_n145 ) , .C1( u0_u12_u1_n147 ) );
  NAND2_X1 u0_u12_u1_U50 (.ZN( u0_u12_u1_n129 ) , .A2( u0_u12_u1_n95 ) , .A1( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U51 (.A1( u0_u12_u1_n102 ) , .ZN( u0_u12_u1_n154 ) , .A2( u0_u12_u1_n99 ) );
  NAND2_X1 u0_u12_u1_U52 (.A2( u0_u12_u1_n100 ) , .ZN( u0_u12_u1_n135 ) , .A1( u0_u12_u1_n99 ) );
  AOI21_X1 u0_u12_u1_U53 (.A( u0_u12_u1_n152 ) , .B2( u0_u12_u1_n153 ) , .B1( u0_u12_u1_n154 ) , .ZN( u0_u12_u1_n158 ) );
  INV_X1 u0_u12_u1_U54 (.A( u0_u12_u1_n160 ) , .ZN( u0_u12_u1_n175 ) );
  NAND2_X1 u0_u12_u1_U55 (.A1( u0_u12_u1_n100 ) , .ZN( u0_u12_u1_n116 ) , .A2( u0_u12_u1_n95 ) );
  NAND2_X1 u0_u12_u1_U56 (.A1( u0_u12_u1_n102 ) , .ZN( u0_u12_u1_n131 ) , .A2( u0_u12_u1_n95 ) );
  NAND2_X1 u0_u12_u1_U57 (.A2( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n121 ) , .A1( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U58 (.A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n153 ) , .A2( u0_u12_u1_n98 ) );
  NAND2_X1 u0_u12_u1_U59 (.A2( u0_u12_u1_n104 ) , .A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n133 ) );
  AOI22_X1 u0_u12_u1_U6 (.B2( u0_u12_u1_n113 ) , .A2( u0_u12_u1_n114 ) , .ZN( u0_u12_u1_n125 ) , .A1( u0_u12_u1_n171 ) , .B1( u0_u12_u1_n173 ) );
  NAND2_X1 u0_u12_u1_U60 (.ZN( u0_u12_u1_n150 ) , .A2( u0_u12_u1_n98 ) , .A1( u0_u12_u1_n99 ) );
  NAND2_X1 u0_u12_u1_U61 (.A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n155 ) , .A2( u0_u12_u1_n95 ) );
  OAI21_X1 u0_u12_u1_U62 (.ZN( u0_u12_u1_n109 ) , .B1( u0_u12_u1_n129 ) , .B2( u0_u12_u1_n160 ) , .A( u0_u12_u1_n167 ) );
  NAND2_X1 u0_u12_u1_U63 (.A2( u0_u12_u1_n100 ) , .A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n120 ) );
  NAND2_X1 u0_u12_u1_U64 (.A1( u0_u12_u1_n102 ) , .A2( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n115 ) );
  NAND2_X1 u0_u12_u1_U65 (.A2( u0_u12_u1_n100 ) , .A1( u0_u12_u1_n104 ) , .ZN( u0_u12_u1_n151 ) );
  NAND2_X1 u0_u12_u1_U66 (.A2( u0_u12_u1_n103 ) , .A1( u0_u12_u1_n105 ) , .ZN( u0_u12_u1_n161 ) );
  INV_X1 u0_u12_u1_U67 (.A( u0_u12_u1_n152 ) , .ZN( u0_u12_u1_n173 ) );
  INV_X1 u0_u12_u1_U68 (.A( u0_u12_u1_n128 ) , .ZN( u0_u12_u1_n172 ) );
  NAND2_X1 u0_u12_u1_U69 (.A2( u0_u12_u1_n102 ) , .A1( u0_u12_u1_n103 ) , .ZN( u0_u12_u1_n123 ) );
  NAND2_X1 u0_u12_u1_U7 (.ZN( u0_u12_u1_n114 ) , .A1( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n156 ) );
  NOR2_X1 u0_u12_u1_U70 (.A2( u0_u12_X_7 ) , .A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n95 ) );
  NOR2_X1 u0_u12_u1_U71 (.A1( u0_u12_X_12 ) , .A2( u0_u12_X_9 ) , .ZN( u0_u12_u1_n100 ) );
  NOR2_X1 u0_u12_u1_U72 (.A2( u0_u12_X_8 ) , .A1( u0_u12_u1_n177 ) , .ZN( u0_u12_u1_n99 ) );
  NOR2_X1 u0_u12_u1_U73 (.A2( u0_u12_X_12 ) , .ZN( u0_u12_u1_n102 ) , .A1( u0_u12_u1_n176 ) );
  NOR2_X1 u0_u12_u1_U74 (.A2( u0_u12_X_9 ) , .ZN( u0_u12_u1_n105 ) , .A1( u0_u12_u1_n168 ) );
  NAND2_X1 u0_u12_u1_U75 (.A1( u0_u12_X_10 ) , .ZN( u0_u12_u1_n160 ) , .A2( u0_u12_u1_n169 ) );
  NAND2_X1 u0_u12_u1_U76 (.A2( u0_u12_X_10 ) , .A1( u0_u12_X_11 ) , .ZN( u0_u12_u1_n152 ) );
  NAND2_X1 u0_u12_u1_U77 (.A1( u0_u12_X_11 ) , .ZN( u0_u12_u1_n128 ) , .A2( u0_u12_u1_n170 ) );
  AND2_X1 u0_u12_u1_U78 (.A2( u0_u12_X_7 ) , .A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n104 ) );
  AND2_X1 u0_u12_u1_U79 (.A1( u0_u12_X_8 ) , .ZN( u0_u12_u1_n103 ) , .A2( u0_u12_u1_n177 ) );
  AOI22_X1 u0_u12_u1_U8 (.B2( u0_u12_u1_n136 ) , .A2( u0_u12_u1_n137 ) , .ZN( u0_u12_u1_n143 ) , .A1( u0_u12_u1_n171 ) , .B1( u0_u12_u1_n173 ) );
  INV_X1 u0_u12_u1_U80 (.A( u0_u12_X_10 ) , .ZN( u0_u12_u1_n170 ) );
  INV_X1 u0_u12_u1_U81 (.A( u0_u12_X_9 ) , .ZN( u0_u12_u1_n176 ) );
  INV_X1 u0_u12_u1_U82 (.A( u0_u12_X_11 ) , .ZN( u0_u12_u1_n169 ) );
  INV_X1 u0_u12_u1_U83 (.A( u0_u12_X_12 ) , .ZN( u0_u12_u1_n168 ) );
  INV_X1 u0_u12_u1_U84 (.A( u0_u12_X_7 ) , .ZN( u0_u12_u1_n177 ) );
  NAND4_X1 u0_u12_u1_U85 (.ZN( u0_out12_28 ) , .A4( u0_u12_u1_n124 ) , .A3( u0_u12_u1_n125 ) , .A2( u0_u12_u1_n126 ) , .A1( u0_u12_u1_n127 ) );
  OAI21_X1 u0_u12_u1_U86 (.ZN( u0_u12_u1_n127 ) , .B2( u0_u12_u1_n139 ) , .B1( u0_u12_u1_n175 ) , .A( u0_u12_u1_n183 ) );
  OAI21_X1 u0_u12_u1_U87 (.ZN( u0_u12_u1_n126 ) , .B2( u0_u12_u1_n140 ) , .A( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n178 ) );
  NAND4_X1 u0_u12_u1_U88 (.ZN( u0_out12_18 ) , .A4( u0_u12_u1_n165 ) , .A3( u0_u12_u1_n166 ) , .A1( u0_u12_u1_n167 ) , .A2( u0_u12_u1_n186 ) );
  AOI22_X1 u0_u12_u1_U89 (.B2( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n147 ) , .A2( u0_u12_u1_n148 ) , .ZN( u0_u12_u1_n166 ) , .A1( u0_u12_u1_n172 ) );
  INV_X1 u0_u12_u1_U9 (.A( u0_u12_u1_n147 ) , .ZN( u0_u12_u1_n181 ) );
  INV_X1 u0_u12_u1_U90 (.A( u0_u12_u1_n145 ) , .ZN( u0_u12_u1_n186 ) );
  NAND4_X1 u0_u12_u1_U91 (.ZN( u0_out12_2 ) , .A4( u0_u12_u1_n142 ) , .A3( u0_u12_u1_n143 ) , .A2( u0_u12_u1_n144 ) , .A1( u0_u12_u1_n179 ) );
  OAI21_X1 u0_u12_u1_U92 (.B2( u0_u12_u1_n132 ) , .ZN( u0_u12_u1_n144 ) , .A( u0_u12_u1_n146 ) , .B1( u0_u12_u1_n180 ) );
  INV_X1 u0_u12_u1_U93 (.A( u0_u12_u1_n130 ) , .ZN( u0_u12_u1_n179 ) );
  OR4_X1 u0_u12_u1_U94 (.ZN( u0_out12_13 ) , .A4( u0_u12_u1_n108 ) , .A3( u0_u12_u1_n109 ) , .A2( u0_u12_u1_n110 ) , .A1( u0_u12_u1_n111 ) );
  AOI21_X1 u0_u12_u1_U95 (.ZN( u0_u12_u1_n111 ) , .A( u0_u12_u1_n128 ) , .B2( u0_u12_u1_n131 ) , .B1( u0_u12_u1_n135 ) );
  AOI21_X1 u0_u12_u1_U96 (.ZN( u0_u12_u1_n110 ) , .A( u0_u12_u1_n116 ) , .B1( u0_u12_u1_n152 ) , .B2( u0_u12_u1_n160 ) );
  NAND3_X1 u0_u12_u1_U97 (.A3( u0_u12_u1_n149 ) , .A2( u0_u12_u1_n150 ) , .A1( u0_u12_u1_n151 ) , .ZN( u0_u12_u1_n164 ) );
  NAND3_X1 u0_u12_u1_U98 (.A3( u0_u12_u1_n134 ) , .A2( u0_u12_u1_n135 ) , .ZN( u0_u12_u1_n136 ) , .A1( u0_u12_u1_n151 ) );
  NAND3_X1 u0_u12_u1_U99 (.A1( u0_u12_u1_n133 ) , .ZN( u0_u12_u1_n137 ) , .A2( u0_u12_u1_n154 ) , .A3( u0_u12_u1_n181 ) );
  OAI22_X1 u0_u12_u2_U10 (.B1( u0_u12_u2_n151 ) , .A2( u0_u12_u2_n152 ) , .A1( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n160 ) , .B2( u0_u12_u2_n168 ) );
  NAND3_X1 u0_u12_u2_U100 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n104 ) , .A3( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n98 ) );
  NOR3_X1 u0_u12_u2_U11 (.A1( u0_u12_u2_n150 ) , .ZN( u0_u12_u2_n151 ) , .A3( u0_u12_u2_n175 ) , .A2( u0_u12_u2_n188 ) );
  AOI21_X1 u0_u12_u2_U12 (.B2( u0_u12_u2_n123 ) , .ZN( u0_u12_u2_n125 ) , .A( u0_u12_u2_n171 ) , .B1( u0_u12_u2_n184 ) );
  INV_X1 u0_u12_u2_U13 (.A( u0_u12_u2_n150 ) , .ZN( u0_u12_u2_n184 ) );
  AOI21_X1 u0_u12_u2_U14 (.ZN( u0_u12_u2_n144 ) , .B2( u0_u12_u2_n155 ) , .A( u0_u12_u2_n172 ) , .B1( u0_u12_u2_n185 ) );
  AOI21_X1 u0_u12_u2_U15 (.B2( u0_u12_u2_n143 ) , .ZN( u0_u12_u2_n145 ) , .B1( u0_u12_u2_n152 ) , .A( u0_u12_u2_n171 ) );
  INV_X1 u0_u12_u2_U16 (.A( u0_u12_u2_n156 ) , .ZN( u0_u12_u2_n171 ) );
  INV_X1 u0_u12_u2_U17 (.A( u0_u12_u2_n120 ) , .ZN( u0_u12_u2_n188 ) );
  NAND2_X1 u0_u12_u2_U18 (.A2( u0_u12_u2_n122 ) , .ZN( u0_u12_u2_n150 ) , .A1( u0_u12_u2_n152 ) );
  INV_X1 u0_u12_u2_U19 (.A( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n170 ) );
  INV_X1 u0_u12_u2_U20 (.A( u0_u12_u2_n137 ) , .ZN( u0_u12_u2_n173 ) );
  NAND2_X1 u0_u12_u2_U21 (.A1( u0_u12_u2_n132 ) , .A2( u0_u12_u2_n139 ) , .ZN( u0_u12_u2_n157 ) );
  INV_X1 u0_u12_u2_U22 (.A( u0_u12_u2_n113 ) , .ZN( u0_u12_u2_n178 ) );
  INV_X1 u0_u12_u2_U23 (.A( u0_u12_u2_n139 ) , .ZN( u0_u12_u2_n175 ) );
  INV_X1 u0_u12_u2_U24 (.A( u0_u12_u2_n155 ) , .ZN( u0_u12_u2_n181 ) );
  INV_X1 u0_u12_u2_U25 (.A( u0_u12_u2_n119 ) , .ZN( u0_u12_u2_n177 ) );
  INV_X1 u0_u12_u2_U26 (.A( u0_u12_u2_n116 ) , .ZN( u0_u12_u2_n180 ) );
  INV_X1 u0_u12_u2_U27 (.A( u0_u12_u2_n131 ) , .ZN( u0_u12_u2_n179 ) );
  INV_X1 u0_u12_u2_U28 (.A( u0_u12_u2_n154 ) , .ZN( u0_u12_u2_n176 ) );
  NAND2_X1 u0_u12_u2_U29 (.A2( u0_u12_u2_n116 ) , .A1( u0_u12_u2_n117 ) , .ZN( u0_u12_u2_n118 ) );
  NOR2_X1 u0_u12_u2_U3 (.ZN( u0_u12_u2_n121 ) , .A2( u0_u12_u2_n177 ) , .A1( u0_u12_u2_n180 ) );
  INV_X1 u0_u12_u2_U30 (.A( u0_u12_u2_n132 ) , .ZN( u0_u12_u2_n182 ) );
  INV_X1 u0_u12_u2_U31 (.A( u0_u12_u2_n158 ) , .ZN( u0_u12_u2_n183 ) );
  OAI21_X1 u0_u12_u2_U32 (.A( u0_u12_u2_n156 ) , .B1( u0_u12_u2_n157 ) , .ZN( u0_u12_u2_n158 ) , .B2( u0_u12_u2_n179 ) );
  NOR2_X1 u0_u12_u2_U33 (.ZN( u0_u12_u2_n156 ) , .A1( u0_u12_u2_n166 ) , .A2( u0_u12_u2_n169 ) );
  NOR2_X1 u0_u12_u2_U34 (.A2( u0_u12_u2_n114 ) , .ZN( u0_u12_u2_n137 ) , .A1( u0_u12_u2_n140 ) );
  NOR2_X1 u0_u12_u2_U35 (.A2( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n153 ) , .A1( u0_u12_u2_n156 ) );
  AOI211_X1 u0_u12_u2_U36 (.ZN( u0_u12_u2_n130 ) , .C1( u0_u12_u2_n138 ) , .C2( u0_u12_u2_n179 ) , .B( u0_u12_u2_n96 ) , .A( u0_u12_u2_n97 ) );
  OAI22_X1 u0_u12_u2_U37 (.B1( u0_u12_u2_n133 ) , .A2( u0_u12_u2_n137 ) , .A1( u0_u12_u2_n152 ) , .B2( u0_u12_u2_n168 ) , .ZN( u0_u12_u2_n97 ) );
  OAI221_X1 u0_u12_u2_U38 (.B1( u0_u12_u2_n113 ) , .C1( u0_u12_u2_n132 ) , .A( u0_u12_u2_n149 ) , .B2( u0_u12_u2_n171 ) , .C2( u0_u12_u2_n172 ) , .ZN( u0_u12_u2_n96 ) );
  OAI221_X1 u0_u12_u2_U39 (.A( u0_u12_u2_n115 ) , .C2( u0_u12_u2_n123 ) , .B2( u0_u12_u2_n143 ) , .B1( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n163 ) , .C1( u0_u12_u2_n168 ) );
  INV_X1 u0_u12_u2_U4 (.A( u0_u12_u2_n134 ) , .ZN( u0_u12_u2_n185 ) );
  OAI21_X1 u0_u12_u2_U40 (.A( u0_u12_u2_n114 ) , .ZN( u0_u12_u2_n115 ) , .B1( u0_u12_u2_n176 ) , .B2( u0_u12_u2_n178 ) );
  OAI221_X1 u0_u12_u2_U41 (.A( u0_u12_u2_n135 ) , .B2( u0_u12_u2_n136 ) , .B1( u0_u12_u2_n137 ) , .ZN( u0_u12_u2_n162 ) , .C2( u0_u12_u2_n167 ) , .C1( u0_u12_u2_n185 ) );
  AND3_X1 u0_u12_u2_U42 (.A3( u0_u12_u2_n131 ) , .A2( u0_u12_u2_n132 ) , .A1( u0_u12_u2_n133 ) , .ZN( u0_u12_u2_n136 ) );
  AOI22_X1 u0_u12_u2_U43 (.ZN( u0_u12_u2_n135 ) , .B1( u0_u12_u2_n140 ) , .A1( u0_u12_u2_n156 ) , .B2( u0_u12_u2_n180 ) , .A2( u0_u12_u2_n188 ) );
  AOI21_X1 u0_u12_u2_U44 (.ZN( u0_u12_u2_n149 ) , .B1( u0_u12_u2_n173 ) , .B2( u0_u12_u2_n188 ) , .A( u0_u12_u2_n95 ) );
  AND3_X1 u0_u12_u2_U45 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n104 ) , .A3( u0_u12_u2_n156 ) , .ZN( u0_u12_u2_n95 ) );
  OAI21_X1 u0_u12_u2_U46 (.A( u0_u12_u2_n101 ) , .B2( u0_u12_u2_n121 ) , .B1( u0_u12_u2_n153 ) , .ZN( u0_u12_u2_n164 ) );
  NAND2_X1 u0_u12_u2_U47 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n107 ) , .ZN( u0_u12_u2_n155 ) );
  NAND2_X1 u0_u12_u2_U48 (.A2( u0_u12_u2_n105 ) , .A1( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n143 ) );
  NAND2_X1 u0_u12_u2_U49 (.A1( u0_u12_u2_n104 ) , .A2( u0_u12_u2_n106 ) , .ZN( u0_u12_u2_n152 ) );
  NOR4_X1 u0_u12_u2_U5 (.A4( u0_u12_u2_n124 ) , .A3( u0_u12_u2_n125 ) , .A2( u0_u12_u2_n126 ) , .A1( u0_u12_u2_n127 ) , .ZN( u0_u12_u2_n128 ) );
  NAND2_X1 u0_u12_u2_U50 (.A1( u0_u12_u2_n100 ) , .A2( u0_u12_u2_n105 ) , .ZN( u0_u12_u2_n132 ) );
  INV_X1 u0_u12_u2_U51 (.A( u0_u12_u2_n140 ) , .ZN( u0_u12_u2_n168 ) );
  INV_X1 u0_u12_u2_U52 (.A( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n167 ) );
  OAI21_X1 u0_u12_u2_U53 (.A( u0_u12_u2_n141 ) , .B2( u0_u12_u2_n142 ) , .ZN( u0_u12_u2_n146 ) , .B1( u0_u12_u2_n153 ) );
  OAI21_X1 u0_u12_u2_U54 (.A( u0_u12_u2_n140 ) , .ZN( u0_u12_u2_n141 ) , .B1( u0_u12_u2_n176 ) , .B2( u0_u12_u2_n177 ) );
  NOR3_X1 u0_u12_u2_U55 (.ZN( u0_u12_u2_n142 ) , .A3( u0_u12_u2_n175 ) , .A2( u0_u12_u2_n178 ) , .A1( u0_u12_u2_n181 ) );
  NAND2_X1 u0_u12_u2_U56 (.A1( u0_u12_u2_n102 ) , .A2( u0_u12_u2_n106 ) , .ZN( u0_u12_u2_n113 ) );
  NAND2_X1 u0_u12_u2_U57 (.A1( u0_u12_u2_n106 ) , .A2( u0_u12_u2_n107 ) , .ZN( u0_u12_u2_n131 ) );
  NAND2_X1 u0_u12_u2_U58 (.A1( u0_u12_u2_n103 ) , .A2( u0_u12_u2_n107 ) , .ZN( u0_u12_u2_n139 ) );
  NAND2_X1 u0_u12_u2_U59 (.A1( u0_u12_u2_n103 ) , .A2( u0_u12_u2_n105 ) , .ZN( u0_u12_u2_n133 ) );
  AOI21_X1 u0_u12_u2_U6 (.B2( u0_u12_u2_n119 ) , .ZN( u0_u12_u2_n127 ) , .A( u0_u12_u2_n137 ) , .B1( u0_u12_u2_n155 ) );
  NAND2_X1 u0_u12_u2_U60 (.A1( u0_u12_u2_n102 ) , .A2( u0_u12_u2_n103 ) , .ZN( u0_u12_u2_n154 ) );
  NAND2_X1 u0_u12_u2_U61 (.A2( u0_u12_u2_n103 ) , .A1( u0_u12_u2_n104 ) , .ZN( u0_u12_u2_n119 ) );
  NAND2_X1 u0_u12_u2_U62 (.A2( u0_u12_u2_n107 ) , .A1( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n123 ) );
  NAND2_X1 u0_u12_u2_U63 (.A1( u0_u12_u2_n104 ) , .A2( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n122 ) );
  INV_X1 u0_u12_u2_U64 (.A( u0_u12_u2_n114 ) , .ZN( u0_u12_u2_n172 ) );
  NAND2_X1 u0_u12_u2_U65 (.A2( u0_u12_u2_n100 ) , .A1( u0_u12_u2_n102 ) , .ZN( u0_u12_u2_n116 ) );
  NAND2_X1 u0_u12_u2_U66 (.A1( u0_u12_u2_n102 ) , .A2( u0_u12_u2_n108 ) , .ZN( u0_u12_u2_n120 ) );
  NAND2_X1 u0_u12_u2_U67 (.A2( u0_u12_u2_n105 ) , .A1( u0_u12_u2_n106 ) , .ZN( u0_u12_u2_n117 ) );
  INV_X1 u0_u12_u2_U68 (.ZN( u0_u12_u2_n187 ) , .A( u0_u12_u2_n99 ) );
  OAI21_X1 u0_u12_u2_U69 (.B1( u0_u12_u2_n137 ) , .B2( u0_u12_u2_n143 ) , .A( u0_u12_u2_n98 ) , .ZN( u0_u12_u2_n99 ) );
  AOI21_X1 u0_u12_u2_U7 (.ZN( u0_u12_u2_n124 ) , .B1( u0_u12_u2_n131 ) , .B2( u0_u12_u2_n143 ) , .A( u0_u12_u2_n172 ) );
  NOR2_X1 u0_u12_u2_U70 (.A2( u0_u12_X_16 ) , .ZN( u0_u12_u2_n140 ) , .A1( u0_u12_u2_n166 ) );
  NOR2_X1 u0_u12_u2_U71 (.A2( u0_u12_X_13 ) , .A1( u0_u12_X_14 ) , .ZN( u0_u12_u2_n100 ) );
  NOR2_X1 u0_u12_u2_U72 (.A2( u0_u12_X_16 ) , .A1( u0_u12_X_17 ) , .ZN( u0_u12_u2_n138 ) );
  NOR2_X1 u0_u12_u2_U73 (.A2( u0_u12_X_15 ) , .A1( u0_u12_X_18 ) , .ZN( u0_u12_u2_n104 ) );
  NOR2_X1 u0_u12_u2_U74 (.A2( u0_u12_X_14 ) , .ZN( u0_u12_u2_n103 ) , .A1( u0_u12_u2_n174 ) );
  NOR2_X1 u0_u12_u2_U75 (.A2( u0_u12_X_15 ) , .ZN( u0_u12_u2_n102 ) , .A1( u0_u12_u2_n165 ) );
  NOR2_X1 u0_u12_u2_U76 (.A2( u0_u12_X_17 ) , .ZN( u0_u12_u2_n114 ) , .A1( u0_u12_u2_n169 ) );
  AND2_X1 u0_u12_u2_U77 (.A1( u0_u12_X_15 ) , .ZN( u0_u12_u2_n105 ) , .A2( u0_u12_u2_n165 ) );
  AND2_X1 u0_u12_u2_U78 (.A2( u0_u12_X_15 ) , .A1( u0_u12_X_18 ) , .ZN( u0_u12_u2_n107 ) );
  AND2_X1 u0_u12_u2_U79 (.A1( u0_u12_X_14 ) , .ZN( u0_u12_u2_n106 ) , .A2( u0_u12_u2_n174 ) );
  AOI21_X1 u0_u12_u2_U8 (.B2( u0_u12_u2_n120 ) , .B1( u0_u12_u2_n121 ) , .ZN( u0_u12_u2_n126 ) , .A( u0_u12_u2_n167 ) );
  AND2_X1 u0_u12_u2_U80 (.A1( u0_u12_X_13 ) , .A2( u0_u12_X_14 ) , .ZN( u0_u12_u2_n108 ) );
  INV_X1 u0_u12_u2_U81 (.A( u0_u12_X_16 ) , .ZN( u0_u12_u2_n169 ) );
  INV_X1 u0_u12_u2_U82 (.A( u0_u12_X_17 ) , .ZN( u0_u12_u2_n166 ) );
  INV_X1 u0_u12_u2_U83 (.A( u0_u12_X_13 ) , .ZN( u0_u12_u2_n174 ) );
  INV_X1 u0_u12_u2_U84 (.A( u0_u12_X_18 ) , .ZN( u0_u12_u2_n165 ) );
  NAND4_X1 u0_u12_u2_U85 (.ZN( u0_out12_30 ) , .A4( u0_u12_u2_n147 ) , .A3( u0_u12_u2_n148 ) , .A2( u0_u12_u2_n149 ) , .A1( u0_u12_u2_n187 ) );
  AOI21_X1 u0_u12_u2_U86 (.B2( u0_u12_u2_n138 ) , .ZN( u0_u12_u2_n148 ) , .A( u0_u12_u2_n162 ) , .B1( u0_u12_u2_n182 ) );
  NOR3_X1 u0_u12_u2_U87 (.A3( u0_u12_u2_n144 ) , .A2( u0_u12_u2_n145 ) , .A1( u0_u12_u2_n146 ) , .ZN( u0_u12_u2_n147 ) );
  NAND4_X1 u0_u12_u2_U88 (.ZN( u0_out12_24 ) , .A4( u0_u12_u2_n111 ) , .A3( u0_u12_u2_n112 ) , .A1( u0_u12_u2_n130 ) , .A2( u0_u12_u2_n187 ) );
  AOI221_X1 u0_u12_u2_U89 (.A( u0_u12_u2_n109 ) , .B1( u0_u12_u2_n110 ) , .ZN( u0_u12_u2_n111 ) , .C1( u0_u12_u2_n134 ) , .C2( u0_u12_u2_n170 ) , .B2( u0_u12_u2_n173 ) );
  OAI22_X1 u0_u12_u2_U9 (.ZN( u0_u12_u2_n109 ) , .A2( u0_u12_u2_n113 ) , .B2( u0_u12_u2_n133 ) , .B1( u0_u12_u2_n167 ) , .A1( u0_u12_u2_n168 ) );
  AOI21_X1 u0_u12_u2_U90 (.ZN( u0_u12_u2_n112 ) , .B2( u0_u12_u2_n156 ) , .A( u0_u12_u2_n164 ) , .B1( u0_u12_u2_n181 ) );
  NAND4_X1 u0_u12_u2_U91 (.ZN( u0_out12_16 ) , .A4( u0_u12_u2_n128 ) , .A3( u0_u12_u2_n129 ) , .A1( u0_u12_u2_n130 ) , .A2( u0_u12_u2_n186 ) );
  AOI22_X1 u0_u12_u2_U92 (.A2( u0_u12_u2_n118 ) , .ZN( u0_u12_u2_n129 ) , .A1( u0_u12_u2_n140 ) , .B1( u0_u12_u2_n157 ) , .B2( u0_u12_u2_n170 ) );
  INV_X1 u0_u12_u2_U93 (.A( u0_u12_u2_n163 ) , .ZN( u0_u12_u2_n186 ) );
  OR4_X1 u0_u12_u2_U94 (.ZN( u0_out12_6 ) , .A4( u0_u12_u2_n161 ) , .A3( u0_u12_u2_n162 ) , .A2( u0_u12_u2_n163 ) , .A1( u0_u12_u2_n164 ) );
  OR3_X1 u0_u12_u2_U95 (.A2( u0_u12_u2_n159 ) , .A1( u0_u12_u2_n160 ) , .ZN( u0_u12_u2_n161 ) , .A3( u0_u12_u2_n183 ) );
  AOI21_X1 u0_u12_u2_U96 (.B2( u0_u12_u2_n154 ) , .B1( u0_u12_u2_n155 ) , .ZN( u0_u12_u2_n159 ) , .A( u0_u12_u2_n167 ) );
  NAND3_X1 u0_u12_u2_U97 (.A2( u0_u12_u2_n117 ) , .A1( u0_u12_u2_n122 ) , .A3( u0_u12_u2_n123 ) , .ZN( u0_u12_u2_n134 ) );
  NAND3_X1 u0_u12_u2_U98 (.ZN( u0_u12_u2_n110 ) , .A2( u0_u12_u2_n131 ) , .A3( u0_u12_u2_n139 ) , .A1( u0_u12_u2_n154 ) );
  NAND3_X1 u0_u12_u2_U99 (.A2( u0_u12_u2_n100 ) , .ZN( u0_u12_u2_n101 ) , .A1( u0_u12_u2_n104 ) , .A3( u0_u12_u2_n114 ) );
  OAI22_X1 u0_u12_u3_U10 (.B1( u0_u12_u3_n113 ) , .A2( u0_u12_u3_n135 ) , .A1( u0_u12_u3_n150 ) , .B2( u0_u12_u3_n164 ) , .ZN( u0_u12_u3_n98 ) );
  OAI211_X1 u0_u12_u3_U11 (.B( u0_u12_u3_n106 ) , .ZN( u0_u12_u3_n119 ) , .C2( u0_u12_u3_n128 ) , .C1( u0_u12_u3_n167 ) , .A( u0_u12_u3_n181 ) );
  AOI221_X1 u0_u12_u3_U12 (.C1( u0_u12_u3_n105 ) , .ZN( u0_u12_u3_n106 ) , .A( u0_u12_u3_n131 ) , .B2( u0_u12_u3_n132 ) , .C2( u0_u12_u3_n133 ) , .B1( u0_u12_u3_n169 ) );
  INV_X1 u0_u12_u3_U13 (.ZN( u0_u12_u3_n181 ) , .A( u0_u12_u3_n98 ) );
  NAND2_X1 u0_u12_u3_U14 (.ZN( u0_u12_u3_n105 ) , .A2( u0_u12_u3_n130 ) , .A1( u0_u12_u3_n155 ) );
  AOI22_X1 u0_u12_u3_U15 (.B1( u0_u12_u3_n115 ) , .A2( u0_u12_u3_n116 ) , .ZN( u0_u12_u3_n123 ) , .B2( u0_u12_u3_n133 ) , .A1( u0_u12_u3_n169 ) );
  NAND2_X1 u0_u12_u3_U16 (.ZN( u0_u12_u3_n116 ) , .A2( u0_u12_u3_n151 ) , .A1( u0_u12_u3_n182 ) );
  NOR2_X1 u0_u12_u3_U17 (.ZN( u0_u12_u3_n126 ) , .A2( u0_u12_u3_n150 ) , .A1( u0_u12_u3_n164 ) );
  AOI21_X1 u0_u12_u3_U18 (.ZN( u0_u12_u3_n112 ) , .B2( u0_u12_u3_n146 ) , .B1( u0_u12_u3_n155 ) , .A( u0_u12_u3_n167 ) );
  NAND2_X1 u0_u12_u3_U19 (.A1( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n142 ) , .A2( u0_u12_u3_n164 ) );
  NAND2_X1 u0_u12_u3_U20 (.ZN( u0_u12_u3_n132 ) , .A2( u0_u12_u3_n152 ) , .A1( u0_u12_u3_n156 ) );
  AND2_X1 u0_u12_u3_U21 (.A2( u0_u12_u3_n113 ) , .A1( u0_u12_u3_n114 ) , .ZN( u0_u12_u3_n151 ) );
  INV_X1 u0_u12_u3_U22 (.A( u0_u12_u3_n133 ) , .ZN( u0_u12_u3_n165 ) );
  INV_X1 u0_u12_u3_U23 (.A( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n170 ) );
  NAND2_X1 u0_u12_u3_U24 (.A1( u0_u12_u3_n107 ) , .A2( u0_u12_u3_n108 ) , .ZN( u0_u12_u3_n140 ) );
  NAND2_X1 u0_u12_u3_U25 (.ZN( u0_u12_u3_n117 ) , .A1( u0_u12_u3_n124 ) , .A2( u0_u12_u3_n148 ) );
  NAND2_X1 u0_u12_u3_U26 (.ZN( u0_u12_u3_n143 ) , .A1( u0_u12_u3_n165 ) , .A2( u0_u12_u3_n167 ) );
  INV_X1 u0_u12_u3_U27 (.A( u0_u12_u3_n130 ) , .ZN( u0_u12_u3_n177 ) );
  INV_X1 u0_u12_u3_U28 (.A( u0_u12_u3_n128 ) , .ZN( u0_u12_u3_n176 ) );
  INV_X1 u0_u12_u3_U29 (.A( u0_u12_u3_n155 ) , .ZN( u0_u12_u3_n174 ) );
  INV_X1 u0_u12_u3_U3 (.A( u0_u12_u3_n129 ) , .ZN( u0_u12_u3_n183 ) );
  INV_X1 u0_u12_u3_U30 (.A( u0_u12_u3_n139 ) , .ZN( u0_u12_u3_n185 ) );
  NOR2_X1 u0_u12_u3_U31 (.ZN( u0_u12_u3_n135 ) , .A2( u0_u12_u3_n141 ) , .A1( u0_u12_u3_n169 ) );
  OAI222_X1 u0_u12_u3_U32 (.C2( u0_u12_u3_n107 ) , .A2( u0_u12_u3_n108 ) , .B1( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n138 ) , .B2( u0_u12_u3_n146 ) , .C1( u0_u12_u3_n154 ) , .A1( u0_u12_u3_n164 ) );
  NOR4_X1 u0_u12_u3_U33 (.A4( u0_u12_u3_n157 ) , .A3( u0_u12_u3_n158 ) , .A2( u0_u12_u3_n159 ) , .A1( u0_u12_u3_n160 ) , .ZN( u0_u12_u3_n161 ) );
  AOI21_X1 u0_u12_u3_U34 (.B2( u0_u12_u3_n152 ) , .B1( u0_u12_u3_n153 ) , .ZN( u0_u12_u3_n158 ) , .A( u0_u12_u3_n164 ) );
  AOI21_X1 u0_u12_u3_U35 (.A( u0_u12_u3_n154 ) , .B2( u0_u12_u3_n155 ) , .B1( u0_u12_u3_n156 ) , .ZN( u0_u12_u3_n157 ) );
  AOI21_X1 u0_u12_u3_U36 (.A( u0_u12_u3_n149 ) , .B2( u0_u12_u3_n150 ) , .B1( u0_u12_u3_n151 ) , .ZN( u0_u12_u3_n159 ) );
  AOI211_X1 u0_u12_u3_U37 (.ZN( u0_u12_u3_n109 ) , .A( u0_u12_u3_n119 ) , .C2( u0_u12_u3_n129 ) , .B( u0_u12_u3_n138 ) , .C1( u0_u12_u3_n141 ) );
  AOI211_X1 u0_u12_u3_U38 (.B( u0_u12_u3_n119 ) , .A( u0_u12_u3_n120 ) , .C2( u0_u12_u3_n121 ) , .ZN( u0_u12_u3_n122 ) , .C1( u0_u12_u3_n179 ) );
  INV_X1 u0_u12_u3_U39 (.A( u0_u12_u3_n156 ) , .ZN( u0_u12_u3_n179 ) );
  INV_X1 u0_u12_u3_U4 (.A( u0_u12_u3_n140 ) , .ZN( u0_u12_u3_n182 ) );
  OAI22_X1 u0_u12_u3_U40 (.B1( u0_u12_u3_n118 ) , .ZN( u0_u12_u3_n120 ) , .A1( u0_u12_u3_n135 ) , .B2( u0_u12_u3_n154 ) , .A2( u0_u12_u3_n178 ) );
  AND3_X1 u0_u12_u3_U41 (.ZN( u0_u12_u3_n118 ) , .A2( u0_u12_u3_n124 ) , .A1( u0_u12_u3_n144 ) , .A3( u0_u12_u3_n152 ) );
  INV_X1 u0_u12_u3_U42 (.A( u0_u12_u3_n121 ) , .ZN( u0_u12_u3_n164 ) );
  NAND2_X1 u0_u12_u3_U43 (.ZN( u0_u12_u3_n133 ) , .A1( u0_u12_u3_n154 ) , .A2( u0_u12_u3_n164 ) );
  OAI211_X1 u0_u12_u3_U44 (.B( u0_u12_u3_n127 ) , .ZN( u0_u12_u3_n139 ) , .C1( u0_u12_u3_n150 ) , .C2( u0_u12_u3_n154 ) , .A( u0_u12_u3_n184 ) );
  INV_X1 u0_u12_u3_U45 (.A( u0_u12_u3_n125 ) , .ZN( u0_u12_u3_n184 ) );
  AOI221_X1 u0_u12_u3_U46 (.A( u0_u12_u3_n126 ) , .ZN( u0_u12_u3_n127 ) , .C2( u0_u12_u3_n132 ) , .C1( u0_u12_u3_n169 ) , .B2( u0_u12_u3_n170 ) , .B1( u0_u12_u3_n174 ) );
  OAI22_X1 u0_u12_u3_U47 (.A1( u0_u12_u3_n124 ) , .ZN( u0_u12_u3_n125 ) , .B2( u0_u12_u3_n145 ) , .A2( u0_u12_u3_n165 ) , .B1( u0_u12_u3_n167 ) );
  NOR2_X1 u0_u12_u3_U48 (.A1( u0_u12_u3_n113 ) , .ZN( u0_u12_u3_n131 ) , .A2( u0_u12_u3_n154 ) );
  NAND2_X1 u0_u12_u3_U49 (.A1( u0_u12_u3_n103 ) , .ZN( u0_u12_u3_n150 ) , .A2( u0_u12_u3_n99 ) );
  INV_X1 u0_u12_u3_U5 (.A( u0_u12_u3_n117 ) , .ZN( u0_u12_u3_n178 ) );
  NAND2_X1 u0_u12_u3_U50 (.A2( u0_u12_u3_n102 ) , .ZN( u0_u12_u3_n155 ) , .A1( u0_u12_u3_n97 ) );
  INV_X1 u0_u12_u3_U51 (.A( u0_u12_u3_n141 ) , .ZN( u0_u12_u3_n167 ) );
  AOI21_X1 u0_u12_u3_U52 (.B2( u0_u12_u3_n114 ) , .B1( u0_u12_u3_n146 ) , .A( u0_u12_u3_n154 ) , .ZN( u0_u12_u3_n94 ) );
  AOI21_X1 u0_u12_u3_U53 (.ZN( u0_u12_u3_n110 ) , .B2( u0_u12_u3_n142 ) , .B1( u0_u12_u3_n186 ) , .A( u0_u12_u3_n95 ) );
  INV_X1 u0_u12_u3_U54 (.A( u0_u12_u3_n145 ) , .ZN( u0_u12_u3_n186 ) );
  AOI21_X1 u0_u12_u3_U55 (.B1( u0_u12_u3_n124 ) , .A( u0_u12_u3_n149 ) , .B2( u0_u12_u3_n155 ) , .ZN( u0_u12_u3_n95 ) );
  INV_X1 u0_u12_u3_U56 (.A( u0_u12_u3_n149 ) , .ZN( u0_u12_u3_n169 ) );
  NAND2_X1 u0_u12_u3_U57 (.ZN( u0_u12_u3_n124 ) , .A1( u0_u12_u3_n96 ) , .A2( u0_u12_u3_n97 ) );
  NAND2_X1 u0_u12_u3_U58 (.A2( u0_u12_u3_n100 ) , .ZN( u0_u12_u3_n146 ) , .A1( u0_u12_u3_n96 ) );
  NAND2_X1 u0_u12_u3_U59 (.A1( u0_u12_u3_n101 ) , .ZN( u0_u12_u3_n145 ) , .A2( u0_u12_u3_n99 ) );
  AOI221_X1 u0_u12_u3_U6 (.A( u0_u12_u3_n131 ) , .C2( u0_u12_u3_n132 ) , .C1( u0_u12_u3_n133 ) , .ZN( u0_u12_u3_n134 ) , .B1( u0_u12_u3_n143 ) , .B2( u0_u12_u3_n177 ) );
  NAND2_X1 u0_u12_u3_U60 (.A1( u0_u12_u3_n100 ) , .ZN( u0_u12_u3_n156 ) , .A2( u0_u12_u3_n99 ) );
  NAND2_X1 u0_u12_u3_U61 (.A2( u0_u12_u3_n101 ) , .A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n148 ) );
  NAND2_X1 u0_u12_u3_U62 (.A1( u0_u12_u3_n100 ) , .A2( u0_u12_u3_n102 ) , .ZN( u0_u12_u3_n128 ) );
  NAND2_X1 u0_u12_u3_U63 (.A2( u0_u12_u3_n101 ) , .A1( u0_u12_u3_n102 ) , .ZN( u0_u12_u3_n152 ) );
  NAND2_X1 u0_u12_u3_U64 (.A2( u0_u12_u3_n101 ) , .ZN( u0_u12_u3_n114 ) , .A1( u0_u12_u3_n96 ) );
  NAND2_X1 u0_u12_u3_U65 (.ZN( u0_u12_u3_n107 ) , .A1( u0_u12_u3_n97 ) , .A2( u0_u12_u3_n99 ) );
  NAND2_X1 u0_u12_u3_U66 (.A2( u0_u12_u3_n100 ) , .A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n113 ) );
  NAND2_X1 u0_u12_u3_U67 (.A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n153 ) , .A2( u0_u12_u3_n97 ) );
  NAND2_X1 u0_u12_u3_U68 (.A2( u0_u12_u3_n103 ) , .A1( u0_u12_u3_n104 ) , .ZN( u0_u12_u3_n130 ) );
  NAND2_X1 u0_u12_u3_U69 (.A2( u0_u12_u3_n103 ) , .ZN( u0_u12_u3_n144 ) , .A1( u0_u12_u3_n96 ) );
  OAI22_X1 u0_u12_u3_U7 (.B2( u0_u12_u3_n147 ) , .A2( u0_u12_u3_n148 ) , .ZN( u0_u12_u3_n160 ) , .B1( u0_u12_u3_n165 ) , .A1( u0_u12_u3_n168 ) );
  NAND2_X1 u0_u12_u3_U70 (.A1( u0_u12_u3_n102 ) , .A2( u0_u12_u3_n103 ) , .ZN( u0_u12_u3_n108 ) );
  NOR2_X1 u0_u12_u3_U71 (.A2( u0_u12_X_19 ) , .A1( u0_u12_X_20 ) , .ZN( u0_u12_u3_n99 ) );
  NOR2_X1 u0_u12_u3_U72 (.A2( u0_u12_X_21 ) , .A1( u0_u12_X_24 ) , .ZN( u0_u12_u3_n103 ) );
  NOR2_X1 u0_u12_u3_U73 (.A2( u0_u12_X_24 ) , .A1( u0_u12_u3_n171 ) , .ZN( u0_u12_u3_n97 ) );
  NOR2_X1 u0_u12_u3_U74 (.A2( u0_u12_X_23 ) , .ZN( u0_u12_u3_n141 ) , .A1( u0_u12_u3_n166 ) );
  NOR2_X1 u0_u12_u3_U75 (.A2( u0_u12_X_19 ) , .A1( u0_u12_u3_n172 ) , .ZN( u0_u12_u3_n96 ) );
  NAND2_X1 u0_u12_u3_U76 (.A1( u0_u12_X_22 ) , .A2( u0_u12_X_23 ) , .ZN( u0_u12_u3_n154 ) );
  NAND2_X1 u0_u12_u3_U77 (.A1( u0_u12_X_23 ) , .ZN( u0_u12_u3_n149 ) , .A2( u0_u12_u3_n166 ) );
  NOR2_X1 u0_u12_u3_U78 (.A2( u0_u12_X_22 ) , .A1( u0_u12_X_23 ) , .ZN( u0_u12_u3_n121 ) );
  AND2_X1 u0_u12_u3_U79 (.A1( u0_u12_X_24 ) , .ZN( u0_u12_u3_n101 ) , .A2( u0_u12_u3_n171 ) );
  AND3_X1 u0_u12_u3_U8 (.A3( u0_u12_u3_n144 ) , .A2( u0_u12_u3_n145 ) , .A1( u0_u12_u3_n146 ) , .ZN( u0_u12_u3_n147 ) );
  AND2_X1 u0_u12_u3_U80 (.A1( u0_u12_X_19 ) , .ZN( u0_u12_u3_n102 ) , .A2( u0_u12_u3_n172 ) );
  AND2_X1 u0_u12_u3_U81 (.A1( u0_u12_X_21 ) , .A2( u0_u12_X_24 ) , .ZN( u0_u12_u3_n100 ) );
  AND2_X1 u0_u12_u3_U82 (.A2( u0_u12_X_19 ) , .A1( u0_u12_X_20 ) , .ZN( u0_u12_u3_n104 ) );
  INV_X1 u0_u12_u3_U83 (.A( u0_u12_X_22 ) , .ZN( u0_u12_u3_n166 ) );
  INV_X1 u0_u12_u3_U84 (.A( u0_u12_X_21 ) , .ZN( u0_u12_u3_n171 ) );
  INV_X1 u0_u12_u3_U85 (.A( u0_u12_X_20 ) , .ZN( u0_u12_u3_n172 ) );
  OR4_X1 u0_u12_u3_U86 (.ZN( u0_out12_10 ) , .A4( u0_u12_u3_n136 ) , .A3( u0_u12_u3_n137 ) , .A1( u0_u12_u3_n138 ) , .A2( u0_u12_u3_n139 ) );
  OAI222_X1 u0_u12_u3_U87 (.C1( u0_u12_u3_n128 ) , .ZN( u0_u12_u3_n137 ) , .B1( u0_u12_u3_n148 ) , .A2( u0_u12_u3_n150 ) , .B2( u0_u12_u3_n154 ) , .C2( u0_u12_u3_n164 ) , .A1( u0_u12_u3_n167 ) );
  OAI221_X1 u0_u12_u3_U88 (.A( u0_u12_u3_n134 ) , .B2( u0_u12_u3_n135 ) , .ZN( u0_u12_u3_n136 ) , .C1( u0_u12_u3_n149 ) , .B1( u0_u12_u3_n151 ) , .C2( u0_u12_u3_n183 ) );
  NAND4_X1 u0_u12_u3_U89 (.ZN( u0_out12_26 ) , .A4( u0_u12_u3_n109 ) , .A3( u0_u12_u3_n110 ) , .A2( u0_u12_u3_n111 ) , .A1( u0_u12_u3_n173 ) );
  INV_X1 u0_u12_u3_U9 (.A( u0_u12_u3_n143 ) , .ZN( u0_u12_u3_n168 ) );
  INV_X1 u0_u12_u3_U90 (.ZN( u0_u12_u3_n173 ) , .A( u0_u12_u3_n94 ) );
  OAI21_X1 u0_u12_u3_U91 (.ZN( u0_u12_u3_n111 ) , .B2( u0_u12_u3_n117 ) , .A( u0_u12_u3_n133 ) , .B1( u0_u12_u3_n176 ) );
  NAND4_X1 u0_u12_u3_U92 (.ZN( u0_out12_20 ) , .A4( u0_u12_u3_n122 ) , .A3( u0_u12_u3_n123 ) , .A1( u0_u12_u3_n175 ) , .A2( u0_u12_u3_n180 ) );
  INV_X1 u0_u12_u3_U93 (.A( u0_u12_u3_n126 ) , .ZN( u0_u12_u3_n180 ) );
  INV_X1 u0_u12_u3_U94 (.A( u0_u12_u3_n112 ) , .ZN( u0_u12_u3_n175 ) );
  NAND4_X1 u0_u12_u3_U95 (.ZN( u0_out12_1 ) , .A4( u0_u12_u3_n161 ) , .A3( u0_u12_u3_n162 ) , .A2( u0_u12_u3_n163 ) , .A1( u0_u12_u3_n185 ) );
  NAND2_X1 u0_u12_u3_U96 (.ZN( u0_u12_u3_n163 ) , .A2( u0_u12_u3_n170 ) , .A1( u0_u12_u3_n176 ) );
  AOI22_X1 u0_u12_u3_U97 (.B2( u0_u12_u3_n140 ) , .B1( u0_u12_u3_n141 ) , .A2( u0_u12_u3_n142 ) , .ZN( u0_u12_u3_n162 ) , .A1( u0_u12_u3_n177 ) );
  NAND3_X1 u0_u12_u3_U98 (.A1( u0_u12_u3_n114 ) , .ZN( u0_u12_u3_n115 ) , .A2( u0_u12_u3_n145 ) , .A3( u0_u12_u3_n153 ) );
  NAND3_X1 u0_u12_u3_U99 (.ZN( u0_u12_u3_n129 ) , .A2( u0_u12_u3_n144 ) , .A1( u0_u12_u3_n153 ) , .A3( u0_u12_u3_n182 ) );
  XOR2_X1 u0_u14_U26 (.B( u0_K15_30 ) , .A( u0_R13_21 ) , .Z( u0_u14_X_30 ) );
  XOR2_X1 u0_u14_U28 (.B( u0_K15_29 ) , .A( u0_R13_20 ) , .Z( u0_u14_X_29 ) );
  XOR2_X1 u0_u14_U29 (.B( u0_K15_28 ) , .A( u0_R13_19 ) , .Z( u0_u14_X_28 ) );
  XOR2_X1 u0_u14_U30 (.B( u0_K15_27 ) , .A( u0_R13_18 ) , .Z( u0_u14_X_27 ) );
  XOR2_X1 u0_u14_U31 (.B( u0_K15_26 ) , .A( u0_R13_17 ) , .Z( u0_u14_X_26 ) );
  XOR2_X1 u0_u14_U32 (.B( u0_K15_25 ) , .A( u0_R13_16 ) , .Z( u0_u14_X_25 ) );
  OAI22_X1 u0_u14_u4_U10 (.B2( u0_u14_u4_n135 ) , .ZN( u0_u14_u4_n137 ) , .B1( u0_u14_u4_n153 ) , .A1( u0_u14_u4_n155 ) , .A2( u0_u14_u4_n171 ) );
  AND3_X1 u0_u14_u4_U11 (.A2( u0_u14_u4_n134 ) , .ZN( u0_u14_u4_n135 ) , .A3( u0_u14_u4_n145 ) , .A1( u0_u14_u4_n157 ) );
  NAND2_X1 u0_u14_u4_U12 (.ZN( u0_u14_u4_n132 ) , .A2( u0_u14_u4_n170 ) , .A1( u0_u14_u4_n173 ) );
  AOI21_X1 u0_u14_u4_U13 (.B2( u0_u14_u4_n160 ) , .B1( u0_u14_u4_n161 ) , .ZN( u0_u14_u4_n162 ) , .A( u0_u14_u4_n170 ) );
  AOI21_X1 u0_u14_u4_U14 (.ZN( u0_u14_u4_n107 ) , .B2( u0_u14_u4_n143 ) , .A( u0_u14_u4_n174 ) , .B1( u0_u14_u4_n184 ) );
  AOI21_X1 u0_u14_u4_U15 (.B2( u0_u14_u4_n158 ) , .B1( u0_u14_u4_n159 ) , .ZN( u0_u14_u4_n163 ) , .A( u0_u14_u4_n174 ) );
  AOI21_X1 u0_u14_u4_U16 (.A( u0_u14_u4_n153 ) , .B2( u0_u14_u4_n154 ) , .B1( u0_u14_u4_n155 ) , .ZN( u0_u14_u4_n165 ) );
  AOI21_X1 u0_u14_u4_U17 (.A( u0_u14_u4_n156 ) , .B2( u0_u14_u4_n157 ) , .ZN( u0_u14_u4_n164 ) , .B1( u0_u14_u4_n184 ) );
  INV_X1 u0_u14_u4_U18 (.A( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n170 ) );
  AND2_X1 u0_u14_u4_U19 (.A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n155 ) , .A1( u0_u14_u4_n160 ) );
  INV_X1 u0_u14_u4_U20 (.A( u0_u14_u4_n156 ) , .ZN( u0_u14_u4_n175 ) );
  NAND2_X1 u0_u14_u4_U21 (.A2( u0_u14_u4_n118 ) , .ZN( u0_u14_u4_n131 ) , .A1( u0_u14_u4_n147 ) );
  NAND2_X1 u0_u14_u4_U22 (.A1( u0_u14_u4_n119 ) , .A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n130 ) );
  NAND2_X1 u0_u14_u4_U23 (.ZN( u0_u14_u4_n117 ) , .A2( u0_u14_u4_n118 ) , .A1( u0_u14_u4_n148 ) );
  NAND2_X1 u0_u14_u4_U24 (.ZN( u0_u14_u4_n129 ) , .A1( u0_u14_u4_n134 ) , .A2( u0_u14_u4_n148 ) );
  AND3_X1 u0_u14_u4_U25 (.A1( u0_u14_u4_n119 ) , .A2( u0_u14_u4_n143 ) , .A3( u0_u14_u4_n154 ) , .ZN( u0_u14_u4_n161 ) );
  AND2_X1 u0_u14_u4_U26 (.A1( u0_u14_u4_n145 ) , .A2( u0_u14_u4_n147 ) , .ZN( u0_u14_u4_n159 ) );
  OR3_X1 u0_u14_u4_U27 (.A3( u0_u14_u4_n114 ) , .A2( u0_u14_u4_n115 ) , .A1( u0_u14_u4_n116 ) , .ZN( u0_u14_u4_n136 ) );
  AOI21_X1 u0_u14_u4_U28 (.A( u0_u14_u4_n113 ) , .ZN( u0_u14_u4_n116 ) , .B2( u0_u14_u4_n173 ) , .B1( u0_u14_u4_n174 ) );
  AOI21_X1 u0_u14_u4_U29 (.ZN( u0_u14_u4_n115 ) , .B2( u0_u14_u4_n145 ) , .B1( u0_u14_u4_n146 ) , .A( u0_u14_u4_n156 ) );
  NOR2_X1 u0_u14_u4_U3 (.ZN( u0_u14_u4_n121 ) , .A1( u0_u14_u4_n181 ) , .A2( u0_u14_u4_n182 ) );
  OAI22_X1 u0_u14_u4_U30 (.ZN( u0_u14_u4_n114 ) , .A2( u0_u14_u4_n121 ) , .B1( u0_u14_u4_n160 ) , .B2( u0_u14_u4_n170 ) , .A1( u0_u14_u4_n171 ) );
  INV_X1 u0_u14_u4_U31 (.A( u0_u14_u4_n158 ) , .ZN( u0_u14_u4_n182 ) );
  INV_X1 u0_u14_u4_U32 (.ZN( u0_u14_u4_n181 ) , .A( u0_u14_u4_n96 ) );
  INV_X1 u0_u14_u4_U33 (.A( u0_u14_u4_n144 ) , .ZN( u0_u14_u4_n179 ) );
  INV_X1 u0_u14_u4_U34 (.A( u0_u14_u4_n157 ) , .ZN( u0_u14_u4_n178 ) );
  NAND2_X1 u0_u14_u4_U35 (.A2( u0_u14_u4_n154 ) , .A1( u0_u14_u4_n96 ) , .ZN( u0_u14_u4_n97 ) );
  INV_X1 u0_u14_u4_U36 (.ZN( u0_u14_u4_n186 ) , .A( u0_u14_u4_n95 ) );
  OAI221_X1 u0_u14_u4_U37 (.C1( u0_u14_u4_n134 ) , .B1( u0_u14_u4_n158 ) , .B2( u0_u14_u4_n171 ) , .C2( u0_u14_u4_n173 ) , .A( u0_u14_u4_n94 ) , .ZN( u0_u14_u4_n95 ) );
  AOI222_X1 u0_u14_u4_U38 (.B2( u0_u14_u4_n132 ) , .A1( u0_u14_u4_n138 ) , .C2( u0_u14_u4_n175 ) , .A2( u0_u14_u4_n179 ) , .C1( u0_u14_u4_n181 ) , .B1( u0_u14_u4_n185 ) , .ZN( u0_u14_u4_n94 ) );
  INV_X1 u0_u14_u4_U39 (.A( u0_u14_u4_n113 ) , .ZN( u0_u14_u4_n185 ) );
  INV_X1 u0_u14_u4_U4 (.A( u0_u14_u4_n117 ) , .ZN( u0_u14_u4_n184 ) );
  INV_X1 u0_u14_u4_U40 (.A( u0_u14_u4_n143 ) , .ZN( u0_u14_u4_n183 ) );
  NOR2_X1 u0_u14_u4_U41 (.ZN( u0_u14_u4_n138 ) , .A1( u0_u14_u4_n168 ) , .A2( u0_u14_u4_n169 ) );
  NOR2_X1 u0_u14_u4_U42 (.A1( u0_u14_u4_n150 ) , .A2( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n153 ) );
  NOR2_X1 u0_u14_u4_U43 (.A2( u0_u14_u4_n128 ) , .A1( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n156 ) );
  AOI22_X1 u0_u14_u4_U44 (.B2( u0_u14_u4_n122 ) , .A1( u0_u14_u4_n123 ) , .ZN( u0_u14_u4_n124 ) , .B1( u0_u14_u4_n128 ) , .A2( u0_u14_u4_n172 ) );
  INV_X1 u0_u14_u4_U45 (.A( u0_u14_u4_n153 ) , .ZN( u0_u14_u4_n172 ) );
  NAND2_X1 u0_u14_u4_U46 (.A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n123 ) , .A1( u0_u14_u4_n161 ) );
  AOI22_X1 u0_u14_u4_U47 (.B2( u0_u14_u4_n132 ) , .A2( u0_u14_u4_n133 ) , .ZN( u0_u14_u4_n140 ) , .A1( u0_u14_u4_n150 ) , .B1( u0_u14_u4_n179 ) );
  NAND2_X1 u0_u14_u4_U48 (.ZN( u0_u14_u4_n133 ) , .A2( u0_u14_u4_n146 ) , .A1( u0_u14_u4_n154 ) );
  NAND2_X1 u0_u14_u4_U49 (.A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n154 ) , .A2( u0_u14_u4_n98 ) );
  NOR4_X1 u0_u14_u4_U5 (.A4( u0_u14_u4_n106 ) , .A3( u0_u14_u4_n107 ) , .A2( u0_u14_u4_n108 ) , .A1( u0_u14_u4_n109 ) , .ZN( u0_u14_u4_n110 ) );
  NAND2_X1 u0_u14_u4_U50 (.A1( u0_u14_u4_n101 ) , .ZN( u0_u14_u4_n158 ) , .A2( u0_u14_u4_n99 ) );
  AOI21_X1 u0_u14_u4_U51 (.ZN( u0_u14_u4_n127 ) , .A( u0_u14_u4_n136 ) , .B2( u0_u14_u4_n150 ) , .B1( u0_u14_u4_n180 ) );
  INV_X1 u0_u14_u4_U52 (.A( u0_u14_u4_n160 ) , .ZN( u0_u14_u4_n180 ) );
  NAND2_X1 u0_u14_u4_U53 (.A2( u0_u14_u4_n104 ) , .A1( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n146 ) );
  NAND2_X1 u0_u14_u4_U54 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n160 ) );
  NAND2_X1 u0_u14_u4_U55 (.ZN( u0_u14_u4_n134 ) , .A1( u0_u14_u4_n98 ) , .A2( u0_u14_u4_n99 ) );
  NAND2_X1 u0_u14_u4_U56 (.A1( u0_u14_u4_n103 ) , .A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n143 ) );
  NAND2_X1 u0_u14_u4_U57 (.A2( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n145 ) , .A1( u0_u14_u4_n98 ) );
  NAND2_X1 u0_u14_u4_U58 (.A1( u0_u14_u4_n100 ) , .A2( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n120 ) );
  NAND2_X1 u0_u14_u4_U59 (.A1( u0_u14_u4_n102 ) , .A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n148 ) );
  AOI21_X1 u0_u14_u4_U6 (.ZN( u0_u14_u4_n106 ) , .B2( u0_u14_u4_n146 ) , .B1( u0_u14_u4_n158 ) , .A( u0_u14_u4_n170 ) );
  NAND2_X1 u0_u14_u4_U60 (.A2( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n157 ) );
  INV_X1 u0_u14_u4_U61 (.A( u0_u14_u4_n150 ) , .ZN( u0_u14_u4_n173 ) );
  INV_X1 u0_u14_u4_U62 (.A( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n171 ) );
  NAND2_X1 u0_u14_u4_U63 (.A1( u0_u14_u4_n100 ) , .ZN( u0_u14_u4_n118 ) , .A2( u0_u14_u4_n99 ) );
  NAND2_X1 u0_u14_u4_U64 (.A2( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n144 ) );
  NAND2_X1 u0_u14_u4_U65 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n96 ) );
  INV_X1 u0_u14_u4_U66 (.A( u0_u14_u4_n128 ) , .ZN( u0_u14_u4_n174 ) );
  NAND2_X1 u0_u14_u4_U67 (.A2( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n119 ) , .A1( u0_u14_u4_n98 ) );
  NAND2_X1 u0_u14_u4_U68 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n147 ) );
  NAND2_X1 u0_u14_u4_U69 (.A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n113 ) , .A1( u0_u14_u4_n99 ) );
  AOI21_X1 u0_u14_u4_U7 (.ZN( u0_u14_u4_n108 ) , .B2( u0_u14_u4_n134 ) , .B1( u0_u14_u4_n155 ) , .A( u0_u14_u4_n156 ) );
  NOR2_X1 u0_u14_u4_U70 (.A2( u0_u14_X_28 ) , .ZN( u0_u14_u4_n150 ) , .A1( u0_u14_u4_n168 ) );
  NOR2_X1 u0_u14_u4_U71 (.A2( u0_u14_X_29 ) , .ZN( u0_u14_u4_n152 ) , .A1( u0_u14_u4_n169 ) );
  NOR2_X1 u0_u14_u4_U72 (.A2( u0_u14_X_30 ) , .ZN( u0_u14_u4_n105 ) , .A1( u0_u14_u4_n176 ) );
  NOR2_X1 u0_u14_u4_U73 (.A2( u0_u14_X_26 ) , .ZN( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n177 ) );
  NOR2_X1 u0_u14_u4_U74 (.A2( u0_u14_X_28 ) , .A1( u0_u14_X_29 ) , .ZN( u0_u14_u4_n128 ) );
  NOR2_X1 u0_u14_u4_U75 (.A2( u0_u14_X_27 ) , .A1( u0_u14_X_30 ) , .ZN( u0_u14_u4_n102 ) );
  NOR2_X1 u0_u14_u4_U76 (.A2( u0_u14_X_25 ) , .A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n98 ) );
  AND2_X1 u0_u14_u4_U77 (.A2( u0_u14_X_25 ) , .A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n104 ) );
  AND2_X1 u0_u14_u4_U78 (.A1( u0_u14_X_30 ) , .A2( u0_u14_u4_n176 ) , .ZN( u0_u14_u4_n99 ) );
  AND2_X1 u0_u14_u4_U79 (.A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n101 ) , .A2( u0_u14_u4_n177 ) );
  AOI21_X1 u0_u14_u4_U8 (.ZN( u0_u14_u4_n109 ) , .A( u0_u14_u4_n153 ) , .B1( u0_u14_u4_n159 ) , .B2( u0_u14_u4_n184 ) );
  AND2_X1 u0_u14_u4_U80 (.A1( u0_u14_X_27 ) , .A2( u0_u14_X_30 ) , .ZN( u0_u14_u4_n103 ) );
  INV_X1 u0_u14_u4_U81 (.A( u0_u14_X_28 ) , .ZN( u0_u14_u4_n169 ) );
  INV_X1 u0_u14_u4_U82 (.A( u0_u14_X_29 ) , .ZN( u0_u14_u4_n168 ) );
  INV_X1 u0_u14_u4_U83 (.A( u0_u14_X_25 ) , .ZN( u0_u14_u4_n177 ) );
  INV_X1 u0_u14_u4_U84 (.A( u0_u14_X_27 ) , .ZN( u0_u14_u4_n176 ) );
  NAND4_X1 u0_u14_u4_U85 (.ZN( u0_out14_25 ) , .A4( u0_u14_u4_n139 ) , .A3( u0_u14_u4_n140 ) , .A2( u0_u14_u4_n141 ) , .A1( u0_u14_u4_n142 ) );
  OAI21_X1 u0_u14_u4_U86 (.A( u0_u14_u4_n128 ) , .B2( u0_u14_u4_n129 ) , .B1( u0_u14_u4_n130 ) , .ZN( u0_u14_u4_n142 ) );
  OAI21_X1 u0_u14_u4_U87 (.B2( u0_u14_u4_n131 ) , .ZN( u0_u14_u4_n141 ) , .A( u0_u14_u4_n175 ) , .B1( u0_u14_u4_n183 ) );
  NAND4_X1 u0_u14_u4_U88 (.ZN( u0_out14_14 ) , .A4( u0_u14_u4_n124 ) , .A3( u0_u14_u4_n125 ) , .A2( u0_u14_u4_n126 ) , .A1( u0_u14_u4_n127 ) );
  AOI22_X1 u0_u14_u4_U89 (.B2( u0_u14_u4_n117 ) , .ZN( u0_u14_u4_n126 ) , .A1( u0_u14_u4_n129 ) , .B1( u0_u14_u4_n152 ) , .A2( u0_u14_u4_n175 ) );
  AOI211_X1 u0_u14_u4_U9 (.B( u0_u14_u4_n136 ) , .A( u0_u14_u4_n137 ) , .C2( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n139 ) , .C1( u0_u14_u4_n182 ) );
  AOI22_X1 u0_u14_u4_U90 (.ZN( u0_u14_u4_n125 ) , .B2( u0_u14_u4_n131 ) , .A2( u0_u14_u4_n132 ) , .B1( u0_u14_u4_n138 ) , .A1( u0_u14_u4_n178 ) );
  NAND4_X1 u0_u14_u4_U91 (.ZN( u0_out14_8 ) , .A4( u0_u14_u4_n110 ) , .A3( u0_u14_u4_n111 ) , .A2( u0_u14_u4_n112 ) , .A1( u0_u14_u4_n186 ) );
  NAND2_X1 u0_u14_u4_U92 (.ZN( u0_u14_u4_n112 ) , .A2( u0_u14_u4_n130 ) , .A1( u0_u14_u4_n150 ) );
  AOI22_X1 u0_u14_u4_U93 (.ZN( u0_u14_u4_n111 ) , .B2( u0_u14_u4_n132 ) , .A1( u0_u14_u4_n152 ) , .B1( u0_u14_u4_n178 ) , .A2( u0_u14_u4_n97 ) );
  AOI22_X1 u0_u14_u4_U94 (.B2( u0_u14_u4_n149 ) , .B1( u0_u14_u4_n150 ) , .A2( u0_u14_u4_n151 ) , .A1( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n167 ) );
  NOR4_X1 u0_u14_u4_U95 (.A4( u0_u14_u4_n162 ) , .A3( u0_u14_u4_n163 ) , .A2( u0_u14_u4_n164 ) , .A1( u0_u14_u4_n165 ) , .ZN( u0_u14_u4_n166 ) );
  NAND3_X1 u0_u14_u4_U96 (.ZN( u0_out14_3 ) , .A3( u0_u14_u4_n166 ) , .A1( u0_u14_u4_n167 ) , .A2( u0_u14_u4_n186 ) );
  NAND3_X1 u0_u14_u4_U97 (.A3( u0_u14_u4_n146 ) , .A2( u0_u14_u4_n147 ) , .A1( u0_u14_u4_n148 ) , .ZN( u0_u14_u4_n149 ) );
  NAND3_X1 u0_u14_u4_U98 (.A3( u0_u14_u4_n143 ) , .A2( u0_u14_u4_n144 ) , .A1( u0_u14_u4_n145 ) , .ZN( u0_u14_u4_n151 ) );
  NAND3_X1 u0_u14_u4_U99 (.A3( u0_u14_u4_n121 ) , .ZN( u0_u14_u4_n122 ) , .A2( u0_u14_u4_n144 ) , .A1( u0_u14_u4_n154 ) );
  XOR2_X1 u0_u1_U1 (.B( u0_K2_9 ) , .A( u0_R0_6 ) , .Z( u0_u1_X_9 ) );
  XOR2_X1 u0_u1_U13 (.B( u0_K2_42 ) , .A( u0_R0_29 ) , .Z( u0_u1_X_42 ) );
  XOR2_X1 u0_u1_U14 (.B( u0_K2_41 ) , .A( u0_R0_28 ) , .Z( u0_u1_X_41 ) );
  XOR2_X1 u0_u1_U15 (.B( u0_K2_40 ) , .A( u0_R0_27 ) , .Z( u0_u1_X_40 ) );
  XOR2_X1 u0_u1_U16 (.B( u0_K2_3 ) , .A( u0_R0_2 ) , .Z( u0_u1_X_3 ) );
  XOR2_X1 u0_u1_U17 (.B( u0_K2_39 ) , .A( u0_R0_26 ) , .Z( u0_u1_X_39 ) );
  XOR2_X1 u0_u1_U18 (.B( u0_K2_38 ) , .A( u0_R0_25 ) , .Z( u0_u1_X_38 ) );
  XOR2_X1 u0_u1_U19 (.B( u0_K2_37 ) , .A( u0_R0_24 ) , .Z( u0_u1_X_37 ) );
  XOR2_X1 u0_u1_U2 (.B( u0_K2_8 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_8 ) );
  XOR2_X1 u0_u1_U20 (.B( u0_K2_36 ) , .A( u0_R0_25 ) , .Z( u0_u1_X_36 ) );
  XOR2_X1 u0_u1_U21 (.B( u0_K2_35 ) , .A( u0_R0_24 ) , .Z( u0_u1_X_35 ) );
  XOR2_X1 u0_u1_U22 (.B( u0_K2_34 ) , .A( u0_R0_23 ) , .Z( u0_u1_X_34 ) );
  XOR2_X1 u0_u1_U23 (.B( u0_K2_33 ) , .A( u0_R0_22 ) , .Z( u0_u1_X_33 ) );
  XOR2_X1 u0_u1_U24 (.B( u0_K2_32 ) , .A( u0_R0_21 ) , .Z( u0_u1_X_32 ) );
  XOR2_X1 u0_u1_U25 (.B( u0_K2_31 ) , .A( u0_R0_20 ) , .Z( u0_u1_X_31 ) );
  XOR2_X1 u0_u1_U26 (.B( u0_K2_30 ) , .A( u0_R0_21 ) , .Z( u0_u1_X_30 ) );
  XOR2_X1 u0_u1_U27 (.B( u0_K2_2 ) , .A( u0_R0_1 ) , .Z( u0_u1_X_2 ) );
  XOR2_X1 u0_u1_U28 (.B( u0_K2_29 ) , .A( u0_R0_20 ) , .Z( u0_u1_X_29 ) );
  XOR2_X1 u0_u1_U29 (.B( u0_K2_28 ) , .A( u0_R0_19 ) , .Z( u0_u1_X_28 ) );
  XOR2_X1 u0_u1_U3 (.B( u0_K2_7 ) , .A( u0_R0_4 ) , .Z( u0_u1_X_7 ) );
  XOR2_X1 u0_u1_U30 (.B( u0_K2_27 ) , .A( u0_R0_18 ) , .Z( u0_u1_X_27 ) );
  XOR2_X1 u0_u1_U31 (.B( u0_K2_26 ) , .A( u0_R0_17 ) , .Z( u0_u1_X_26 ) );
  XOR2_X1 u0_u1_U32 (.B( u0_K2_25 ) , .A( u0_R0_16 ) , .Z( u0_u1_X_25 ) );
  XOR2_X1 u0_u1_U38 (.B( u0_K2_1 ) , .A( u0_R0_32 ) , .Z( u0_u1_X_1 ) );
  XOR2_X1 u0_u1_U4 (.B( u0_K2_6 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_6 ) );
  XOR2_X1 u0_u1_U46 (.B( u0_K2_12 ) , .A( u0_R0_9 ) , .Z( u0_u1_X_12 ) );
  XOR2_X1 u0_u1_U47 (.B( u0_K2_11 ) , .A( u0_R0_8 ) , .Z( u0_u1_X_11 ) );
  XOR2_X1 u0_u1_U48 (.B( u0_K2_10 ) , .A( u0_R0_7 ) , .Z( u0_u1_X_10 ) );
  XOR2_X1 u0_u1_U5 (.B( u0_K2_5 ) , .A( u0_R0_4 ) , .Z( u0_u1_X_5 ) );
  XOR2_X1 u0_u1_U6 (.B( u0_K2_4 ) , .A( u0_R0_3 ) , .Z( u0_u1_X_4 ) );
  AND3_X1 u0_u1_u0_U10 (.A2( u0_u1_u0_n112 ) , .ZN( u0_u1_u0_n127 ) , .A3( u0_u1_u0_n130 ) , .A1( u0_u1_u0_n148 ) );
  NAND2_X1 u0_u1_u0_U11 (.ZN( u0_u1_u0_n113 ) , .A1( u0_u1_u0_n139 ) , .A2( u0_u1_u0_n149 ) );
  AND2_X1 u0_u1_u0_U12 (.ZN( u0_u1_u0_n107 ) , .A1( u0_u1_u0_n130 ) , .A2( u0_u1_u0_n140 ) );
  AND2_X1 u0_u1_u0_U13 (.A2( u0_u1_u0_n129 ) , .A1( u0_u1_u0_n130 ) , .ZN( u0_u1_u0_n151 ) );
  AND2_X1 u0_u1_u0_U14 (.A1( u0_u1_u0_n108 ) , .A2( u0_u1_u0_n125 ) , .ZN( u0_u1_u0_n145 ) );
  INV_X1 u0_u1_u0_U15 (.A( u0_u1_u0_n143 ) , .ZN( u0_u1_u0_n173 ) );
  NOR2_X1 u0_u1_u0_U16 (.A2( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n147 ) , .A1( u0_u1_u0_n160 ) );
  NOR2_X1 u0_u1_u0_U17 (.A1( u0_u1_u0_n163 ) , .A2( u0_u1_u0_n164 ) , .ZN( u0_u1_u0_n95 ) );
  AOI21_X1 u0_u1_u0_U18 (.B1( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n132 ) , .A( u0_u1_u0_n165 ) , .B2( u0_u1_u0_n93 ) );
  INV_X1 u0_u1_u0_U19 (.A( u0_u1_u0_n142 ) , .ZN( u0_u1_u0_n165 ) );
  OAI221_X1 u0_u1_u0_U20 (.C1( u0_u1_u0_n121 ) , .ZN( u0_u1_u0_n122 ) , .B2( u0_u1_u0_n127 ) , .A( u0_u1_u0_n143 ) , .B1( u0_u1_u0_n144 ) , .C2( u0_u1_u0_n147 ) );
  OAI22_X1 u0_u1_u0_U21 (.B1( u0_u1_u0_n125 ) , .ZN( u0_u1_u0_n126 ) , .A1( u0_u1_u0_n138 ) , .A2( u0_u1_u0_n146 ) , .B2( u0_u1_u0_n147 ) );
  OAI22_X1 u0_u1_u0_U22 (.B1( u0_u1_u0_n131 ) , .A1( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n147 ) , .A2( u0_u1_u0_n90 ) , .ZN( u0_u1_u0_n91 ) );
  AND3_X1 u0_u1_u0_U23 (.A3( u0_u1_u0_n121 ) , .A2( u0_u1_u0_n125 ) , .A1( u0_u1_u0_n148 ) , .ZN( u0_u1_u0_n90 ) );
  INV_X1 u0_u1_u0_U24 (.A( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n161 ) );
  NOR2_X1 u0_u1_u0_U25 (.A1( u0_u1_u0_n120 ) , .ZN( u0_u1_u0_n143 ) , .A2( u0_u1_u0_n167 ) );
  OAI221_X1 u0_u1_u0_U26 (.C1( u0_u1_u0_n112 ) , .ZN( u0_u1_u0_n120 ) , .B1( u0_u1_u0_n138 ) , .B2( u0_u1_u0_n141 ) , .C2( u0_u1_u0_n147 ) , .A( u0_u1_u0_n172 ) );
  AOI211_X1 u0_u1_u0_U27 (.B( u0_u1_u0_n115 ) , .A( u0_u1_u0_n116 ) , .C2( u0_u1_u0_n117 ) , .C1( u0_u1_u0_n118 ) , .ZN( u0_u1_u0_n119 ) );
  AOI22_X1 u0_u1_u0_U28 (.B2( u0_u1_u0_n109 ) , .A2( u0_u1_u0_n110 ) , .ZN( u0_u1_u0_n111 ) , .B1( u0_u1_u0_n118 ) , .A1( u0_u1_u0_n160 ) );
  INV_X1 u0_u1_u0_U29 (.A( u0_u1_u0_n118 ) , .ZN( u0_u1_u0_n158 ) );
  INV_X1 u0_u1_u0_U3 (.A( u0_u1_u0_n113 ) , .ZN( u0_u1_u0_n166 ) );
  AOI21_X1 u0_u1_u0_U30 (.ZN( u0_u1_u0_n104 ) , .B1( u0_u1_u0_n107 ) , .B2( u0_u1_u0_n141 ) , .A( u0_u1_u0_n144 ) );
  AOI21_X1 u0_u1_u0_U31 (.B1( u0_u1_u0_n127 ) , .B2( u0_u1_u0_n129 ) , .A( u0_u1_u0_n138 ) , .ZN( u0_u1_u0_n96 ) );
  AOI21_X1 u0_u1_u0_U32 (.ZN( u0_u1_u0_n116 ) , .B2( u0_u1_u0_n142 ) , .A( u0_u1_u0_n144 ) , .B1( u0_u1_u0_n166 ) );
  NAND2_X1 u0_u1_u0_U33 (.A1( u0_u1_u0_n100 ) , .A2( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n125 ) );
  NAND2_X1 u0_u1_u0_U34 (.A2( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n140 ) , .A1( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U35 (.A1( u0_u1_u0_n101 ) , .A2( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n150 ) );
  INV_X1 u0_u1_u0_U36 (.A( u0_u1_u0_n138 ) , .ZN( u0_u1_u0_n160 ) );
  NAND2_X1 u0_u1_u0_U37 (.ZN( u0_u1_u0_n142 ) , .A1( u0_u1_u0_n94 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U38 (.A1( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n128 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U39 (.A2( u0_u1_u0_n102 ) , .A1( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n149 ) );
  AOI21_X1 u0_u1_u0_U4 (.B1( u0_u1_u0_n114 ) , .ZN( u0_u1_u0_n115 ) , .B2( u0_u1_u0_n129 ) , .A( u0_u1_u0_n161 ) );
  NAND2_X1 u0_u1_u0_U40 (.A1( u0_u1_u0_n100 ) , .ZN( u0_u1_u0_n129 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U41 (.A2( u0_u1_u0_n100 ) , .A1( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n139 ) );
  NAND2_X1 u0_u1_u0_U42 (.A2( u0_u1_u0_n100 ) , .ZN( u0_u1_u0_n131 ) , .A1( u0_u1_u0_n92 ) );
  NAND2_X1 u0_u1_u0_U43 (.ZN( u0_u1_u0_n108 ) , .A1( u0_u1_u0_n92 ) , .A2( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U44 (.ZN( u0_u1_u0_n148 ) , .A1( u0_u1_u0_n93 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U45 (.A2( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n114 ) , .A1( u0_u1_u0_n92 ) );
  NAND2_X1 u0_u1_u0_U46 (.A1( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n130 ) , .A2( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U47 (.A2( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n121 ) , .A1( u0_u1_u0_n93 ) );
  INV_X1 u0_u1_u0_U48 (.ZN( u0_u1_u0_n172 ) , .A( u0_u1_u0_n88 ) );
  OAI222_X1 u0_u1_u0_U49 (.C1( u0_u1_u0_n108 ) , .A1( u0_u1_u0_n125 ) , .B2( u0_u1_u0_n128 ) , .B1( u0_u1_u0_n144 ) , .A2( u0_u1_u0_n158 ) , .C2( u0_u1_u0_n161 ) , .ZN( u0_u1_u0_n88 ) );
  AOI21_X1 u0_u1_u0_U5 (.B2( u0_u1_u0_n131 ) , .ZN( u0_u1_u0_n134 ) , .B1( u0_u1_u0_n151 ) , .A( u0_u1_u0_n158 ) );
  NAND2_X1 u0_u1_u0_U50 (.ZN( u0_u1_u0_n112 ) , .A2( u0_u1_u0_n92 ) , .A1( u0_u1_u0_n93 ) );
  OR3_X1 u0_u1_u0_U51 (.A3( u0_u1_u0_n152 ) , .A2( u0_u1_u0_n153 ) , .A1( u0_u1_u0_n154 ) , .ZN( u0_u1_u0_n155 ) );
  AOI21_X1 u0_u1_u0_U52 (.B2( u0_u1_u0_n150 ) , .B1( u0_u1_u0_n151 ) , .ZN( u0_u1_u0_n152 ) , .A( u0_u1_u0_n158 ) );
  AOI21_X1 u0_u1_u0_U53 (.A( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n145 ) , .B1( u0_u1_u0_n146 ) , .ZN( u0_u1_u0_n154 ) );
  AOI21_X1 u0_u1_u0_U54 (.A( u0_u1_u0_n147 ) , .B2( u0_u1_u0_n148 ) , .B1( u0_u1_u0_n149 ) , .ZN( u0_u1_u0_n153 ) );
  INV_X1 u0_u1_u0_U55 (.ZN( u0_u1_u0_n171 ) , .A( u0_u1_u0_n99 ) );
  OAI211_X1 u0_u1_u0_U56 (.C2( u0_u1_u0_n140 ) , .C1( u0_u1_u0_n161 ) , .A( u0_u1_u0_n169 ) , .B( u0_u1_u0_n98 ) , .ZN( u0_u1_u0_n99 ) );
  INV_X1 u0_u1_u0_U57 (.ZN( u0_u1_u0_n169 ) , .A( u0_u1_u0_n91 ) );
  AOI211_X1 u0_u1_u0_U58 (.C1( u0_u1_u0_n118 ) , .A( u0_u1_u0_n123 ) , .B( u0_u1_u0_n96 ) , .C2( u0_u1_u0_n97 ) , .ZN( u0_u1_u0_n98 ) );
  NOR2_X1 u0_u1_u0_U59 (.A2( u0_u1_X_2 ) , .ZN( u0_u1_u0_n103 ) , .A1( u0_u1_u0_n164 ) );
  NOR2_X1 u0_u1_u0_U6 (.A1( u0_u1_u0_n108 ) , .ZN( u0_u1_u0_n123 ) , .A2( u0_u1_u0_n158 ) );
  NOR2_X1 u0_u1_u0_U60 (.A2( u0_u1_X_3 ) , .A1( u0_u1_X_6 ) , .ZN( u0_u1_u0_n94 ) );
  NOR2_X1 u0_u1_u0_U61 (.A2( u0_u1_X_6 ) , .ZN( u0_u1_u0_n100 ) , .A1( u0_u1_u0_n162 ) );
  NOR2_X1 u0_u1_u0_U62 (.A2( u0_u1_X_4 ) , .A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n118 ) );
  NOR2_X1 u0_u1_u0_U63 (.A2( u0_u1_X_1 ) , .A1( u0_u1_X_2 ) , .ZN( u0_u1_u0_n92 ) );
  NOR2_X1 u0_u1_u0_U64 (.A2( u0_u1_X_1 ) , .ZN( u0_u1_u0_n101 ) , .A1( u0_u1_u0_n163 ) );
  NAND2_X1 u0_u1_u0_U65 (.A2( u0_u1_X_4 ) , .A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n144 ) );
  NOR2_X1 u0_u1_u0_U66 (.A2( u0_u1_X_5 ) , .ZN( u0_u1_u0_n136 ) , .A1( u0_u1_u0_n159 ) );
  NAND2_X1 u0_u1_u0_U67 (.A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n138 ) , .A2( u0_u1_u0_n159 ) );
  AND2_X1 u0_u1_u0_U68 (.A2( u0_u1_X_3 ) , .A1( u0_u1_X_6 ) , .ZN( u0_u1_u0_n102 ) );
  AND2_X1 u0_u1_u0_U69 (.A1( u0_u1_X_6 ) , .A2( u0_u1_u0_n162 ) , .ZN( u0_u1_u0_n93 ) );
  OAI21_X1 u0_u1_u0_U7 (.B1( u0_u1_u0_n150 ) , .B2( u0_u1_u0_n158 ) , .A( u0_u1_u0_n172 ) , .ZN( u0_u1_u0_n89 ) );
  INV_X1 u0_u1_u0_U70 (.A( u0_u1_X_4 ) , .ZN( u0_u1_u0_n159 ) );
  INV_X1 u0_u1_u0_U71 (.A( u0_u1_X_1 ) , .ZN( u0_u1_u0_n164 ) );
  INV_X1 u0_u1_u0_U72 (.A( u0_u1_X_2 ) , .ZN( u0_u1_u0_n163 ) );
  INV_X1 u0_u1_u0_U73 (.A( u0_u1_X_3 ) , .ZN( u0_u1_u0_n162 ) );
  INV_X1 u0_u1_u0_U74 (.ZN( u0_u1_u0_n174 ) , .A( u0_u1_u0_n89 ) );
  AOI211_X1 u0_u1_u0_U75 (.B( u0_u1_u0_n104 ) , .A( u0_u1_u0_n105 ) , .ZN( u0_u1_u0_n106 ) , .C2( u0_u1_u0_n113 ) , .C1( u0_u1_u0_n160 ) );
  INV_X1 u0_u1_u0_U76 (.A( u0_u1_u0_n126 ) , .ZN( u0_u1_u0_n168 ) );
  AOI211_X1 u0_u1_u0_U77 (.B( u0_u1_u0_n133 ) , .A( u0_u1_u0_n134 ) , .C2( u0_u1_u0_n135 ) , .C1( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n137 ) );
  OR4_X1 u0_u1_u0_U78 (.ZN( u0_out1_31 ) , .A4( u0_u1_u0_n155 ) , .A2( u0_u1_u0_n156 ) , .A1( u0_u1_u0_n157 ) , .A3( u0_u1_u0_n173 ) );
  AOI21_X1 u0_u1_u0_U79 (.A( u0_u1_u0_n138 ) , .B2( u0_u1_u0_n139 ) , .B1( u0_u1_u0_n140 ) , .ZN( u0_u1_u0_n157 ) );
  AND2_X1 u0_u1_u0_U8 (.A1( u0_u1_u0_n114 ) , .A2( u0_u1_u0_n121 ) , .ZN( u0_u1_u0_n146 ) );
  AOI21_X1 u0_u1_u0_U80 (.B2( u0_u1_u0_n141 ) , .B1( u0_u1_u0_n142 ) , .ZN( u0_u1_u0_n156 ) , .A( u0_u1_u0_n161 ) );
  OR4_X1 u0_u1_u0_U81 (.ZN( u0_out1_17 ) , .A4( u0_u1_u0_n122 ) , .A2( u0_u1_u0_n123 ) , .A1( u0_u1_u0_n124 ) , .A3( u0_u1_u0_n170 ) );
  AOI21_X1 u0_u1_u0_U82 (.B2( u0_u1_u0_n107 ) , .ZN( u0_u1_u0_n124 ) , .B1( u0_u1_u0_n128 ) , .A( u0_u1_u0_n161 ) );
  INV_X1 u0_u1_u0_U83 (.A( u0_u1_u0_n111 ) , .ZN( u0_u1_u0_n170 ) );
  AOI21_X1 u0_u1_u0_U84 (.B1( u0_u1_u0_n132 ) , .ZN( u0_u1_u0_n133 ) , .A( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n166 ) );
  OAI22_X1 u0_u1_u0_U85 (.ZN( u0_u1_u0_n105 ) , .A2( u0_u1_u0_n132 ) , .B1( u0_u1_u0_n146 ) , .A1( u0_u1_u0_n147 ) , .B2( u0_u1_u0_n161 ) );
  NAND2_X1 u0_u1_u0_U86 (.ZN( u0_u1_u0_n110 ) , .A2( u0_u1_u0_n132 ) , .A1( u0_u1_u0_n145 ) );
  INV_X1 u0_u1_u0_U87 (.A( u0_u1_u0_n119 ) , .ZN( u0_u1_u0_n167 ) );
  NAND3_X1 u0_u1_u0_U88 (.ZN( u0_out1_23 ) , .A3( u0_u1_u0_n137 ) , .A1( u0_u1_u0_n168 ) , .A2( u0_u1_u0_n171 ) );
  NAND3_X1 u0_u1_u0_U89 (.A3( u0_u1_u0_n127 ) , .A2( u0_u1_u0_n128 ) , .ZN( u0_u1_u0_n135 ) , .A1( u0_u1_u0_n150 ) );
  AND2_X1 u0_u1_u0_U9 (.A1( u0_u1_u0_n131 ) , .ZN( u0_u1_u0_n141 ) , .A2( u0_u1_u0_n150 ) );
  NAND3_X1 u0_u1_u0_U90 (.ZN( u0_u1_u0_n117 ) , .A3( u0_u1_u0_n132 ) , .A2( u0_u1_u0_n139 ) , .A1( u0_u1_u0_n148 ) );
  NAND3_X1 u0_u1_u0_U91 (.ZN( u0_u1_u0_n109 ) , .A2( u0_u1_u0_n114 ) , .A3( u0_u1_u0_n140 ) , .A1( u0_u1_u0_n149 ) );
  NAND3_X1 u0_u1_u0_U92 (.ZN( u0_out1_9 ) , .A3( u0_u1_u0_n106 ) , .A2( u0_u1_u0_n171 ) , .A1( u0_u1_u0_n174 ) );
  NAND3_X1 u0_u1_u0_U93 (.A2( u0_u1_u0_n128 ) , .A1( u0_u1_u0_n132 ) , .A3( u0_u1_u0_n146 ) , .ZN( u0_u1_u0_n97 ) );
  NOR2_X1 u0_u1_u1_U10 (.A1( u0_u1_u1_n112 ) , .A2( u0_u1_u1_n116 ) , .ZN( u0_u1_u1_n118 ) );
  NAND3_X1 u0_u1_u1_U100 (.ZN( u0_u1_u1_n113 ) , .A1( u0_u1_u1_n120 ) , .A3( u0_u1_u1_n133 ) , .A2( u0_u1_u1_n155 ) );
  OAI21_X1 u0_u1_u1_U11 (.ZN( u0_u1_u1_n101 ) , .B1( u0_u1_u1_n141 ) , .A( u0_u1_u1_n146 ) , .B2( u0_u1_u1_n183 ) );
  AOI21_X1 u0_u1_u1_U12 (.B2( u0_u1_u1_n155 ) , .B1( u0_u1_u1_n156 ) , .ZN( u0_u1_u1_n157 ) , .A( u0_u1_u1_n174 ) );
  OR4_X1 u0_u1_u1_U13 (.A4( u0_u1_u1_n106 ) , .A3( u0_u1_u1_n107 ) , .ZN( u0_u1_u1_n108 ) , .A1( u0_u1_u1_n117 ) , .A2( u0_u1_u1_n184 ) );
  AOI21_X1 u0_u1_u1_U14 (.ZN( u0_u1_u1_n106 ) , .A( u0_u1_u1_n112 ) , .B1( u0_u1_u1_n154 ) , .B2( u0_u1_u1_n156 ) );
  INV_X1 u0_u1_u1_U15 (.A( u0_u1_u1_n101 ) , .ZN( u0_u1_u1_n184 ) );
  AOI21_X1 u0_u1_u1_U16 (.ZN( u0_u1_u1_n107 ) , .B1( u0_u1_u1_n134 ) , .B2( u0_u1_u1_n149 ) , .A( u0_u1_u1_n174 ) );
  NAND2_X1 u0_u1_u1_U17 (.ZN( u0_u1_u1_n140 ) , .A2( u0_u1_u1_n150 ) , .A1( u0_u1_u1_n155 ) );
  NAND2_X1 u0_u1_u1_U18 (.A1( u0_u1_u1_n131 ) , .ZN( u0_u1_u1_n147 ) , .A2( u0_u1_u1_n153 ) );
  INV_X1 u0_u1_u1_U19 (.A( u0_u1_u1_n139 ) , .ZN( u0_u1_u1_n174 ) );
  INV_X1 u0_u1_u1_U20 (.A( u0_u1_u1_n112 ) , .ZN( u0_u1_u1_n171 ) );
  NAND2_X1 u0_u1_u1_U21 (.ZN( u0_u1_u1_n141 ) , .A1( u0_u1_u1_n153 ) , .A2( u0_u1_u1_n156 ) );
  AND2_X1 u0_u1_u1_U22 (.A1( u0_u1_u1_n123 ) , .ZN( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n161 ) );
  NAND2_X1 u0_u1_u1_U23 (.A2( u0_u1_u1_n115 ) , .A1( u0_u1_u1_n116 ) , .ZN( u0_u1_u1_n148 ) );
  NAND2_X1 u0_u1_u1_U24 (.A2( u0_u1_u1_n133 ) , .A1( u0_u1_u1_n135 ) , .ZN( u0_u1_u1_n159 ) );
  NAND2_X1 u0_u1_u1_U25 (.A2( u0_u1_u1_n115 ) , .A1( u0_u1_u1_n120 ) , .ZN( u0_u1_u1_n132 ) );
  INV_X1 u0_u1_u1_U26 (.A( u0_u1_u1_n154 ) , .ZN( u0_u1_u1_n178 ) );
  INV_X1 u0_u1_u1_U27 (.A( u0_u1_u1_n151 ) , .ZN( u0_u1_u1_n183 ) );
  AND2_X1 u0_u1_u1_U28 (.A1( u0_u1_u1_n129 ) , .A2( u0_u1_u1_n133 ) , .ZN( u0_u1_u1_n149 ) );
  INV_X1 u0_u1_u1_U29 (.A( u0_u1_u1_n131 ) , .ZN( u0_u1_u1_n180 ) );
  INV_X1 u0_u1_u1_U3 (.A( u0_u1_u1_n159 ) , .ZN( u0_u1_u1_n182 ) );
  AOI221_X1 u0_u1_u1_U30 (.B1( u0_u1_u1_n140 ) , .ZN( u0_u1_u1_n167 ) , .B2( u0_u1_u1_n172 ) , .C2( u0_u1_u1_n175 ) , .C1( u0_u1_u1_n178 ) , .A( u0_u1_u1_n188 ) );
  INV_X1 u0_u1_u1_U31 (.ZN( u0_u1_u1_n188 ) , .A( u0_u1_u1_n97 ) );
  AOI211_X1 u0_u1_u1_U32 (.A( u0_u1_u1_n118 ) , .C1( u0_u1_u1_n132 ) , .C2( u0_u1_u1_n139 ) , .B( u0_u1_u1_n96 ) , .ZN( u0_u1_u1_n97 ) );
  AOI21_X1 u0_u1_u1_U33 (.B2( u0_u1_u1_n121 ) , .B1( u0_u1_u1_n135 ) , .A( u0_u1_u1_n152 ) , .ZN( u0_u1_u1_n96 ) );
  OAI221_X1 u0_u1_u1_U34 (.A( u0_u1_u1_n119 ) , .C2( u0_u1_u1_n129 ) , .ZN( u0_u1_u1_n138 ) , .B2( u0_u1_u1_n152 ) , .C1( u0_u1_u1_n174 ) , .B1( u0_u1_u1_n187 ) );
  INV_X1 u0_u1_u1_U35 (.A( u0_u1_u1_n148 ) , .ZN( u0_u1_u1_n187 ) );
  AOI211_X1 u0_u1_u1_U36 (.B( u0_u1_u1_n117 ) , .A( u0_u1_u1_n118 ) , .ZN( u0_u1_u1_n119 ) , .C2( u0_u1_u1_n146 ) , .C1( u0_u1_u1_n159 ) );
  NOR2_X1 u0_u1_u1_U37 (.A1( u0_u1_u1_n168 ) , .A2( u0_u1_u1_n176 ) , .ZN( u0_u1_u1_n98 ) );
  AOI211_X1 u0_u1_u1_U38 (.B( u0_u1_u1_n162 ) , .A( u0_u1_u1_n163 ) , .C2( u0_u1_u1_n164 ) , .ZN( u0_u1_u1_n165 ) , .C1( u0_u1_u1_n171 ) );
  AOI21_X1 u0_u1_u1_U39 (.A( u0_u1_u1_n160 ) , .B2( u0_u1_u1_n161 ) , .ZN( u0_u1_u1_n162 ) , .B1( u0_u1_u1_n182 ) );
  AOI221_X1 u0_u1_u1_U4 (.A( u0_u1_u1_n138 ) , .C2( u0_u1_u1_n139 ) , .C1( u0_u1_u1_n140 ) , .B2( u0_u1_u1_n141 ) , .ZN( u0_u1_u1_n142 ) , .B1( u0_u1_u1_n175 ) );
  OR2_X1 u0_u1_u1_U40 (.A2( u0_u1_u1_n157 ) , .A1( u0_u1_u1_n158 ) , .ZN( u0_u1_u1_n163 ) );
  OAI21_X1 u0_u1_u1_U41 (.B2( u0_u1_u1_n123 ) , .ZN( u0_u1_u1_n145 ) , .B1( u0_u1_u1_n160 ) , .A( u0_u1_u1_n185 ) );
  INV_X1 u0_u1_u1_U42 (.A( u0_u1_u1_n122 ) , .ZN( u0_u1_u1_n185 ) );
  AOI21_X1 u0_u1_u1_U43 (.B2( u0_u1_u1_n120 ) , .B1( u0_u1_u1_n121 ) , .ZN( u0_u1_u1_n122 ) , .A( u0_u1_u1_n128 ) );
  NAND2_X1 u0_u1_u1_U44 (.A1( u0_u1_u1_n128 ) , .ZN( u0_u1_u1_n146 ) , .A2( u0_u1_u1_n160 ) );
  NAND2_X1 u0_u1_u1_U45 (.A2( u0_u1_u1_n112 ) , .ZN( u0_u1_u1_n139 ) , .A1( u0_u1_u1_n152 ) );
  NAND2_X1 u0_u1_u1_U46 (.A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n156 ) , .A2( u0_u1_u1_n99 ) );
  NOR2_X1 u0_u1_u1_U47 (.ZN( u0_u1_u1_n117 ) , .A1( u0_u1_u1_n121 ) , .A2( u0_u1_u1_n160 ) );
  AOI21_X1 u0_u1_u1_U48 (.A( u0_u1_u1_n128 ) , .B2( u0_u1_u1_n129 ) , .ZN( u0_u1_u1_n130 ) , .B1( u0_u1_u1_n150 ) );
  NAND2_X1 u0_u1_u1_U49 (.ZN( u0_u1_u1_n112 ) , .A1( u0_u1_u1_n169 ) , .A2( u0_u1_u1_n170 ) );
  AOI211_X1 u0_u1_u1_U5 (.ZN( u0_u1_u1_n124 ) , .A( u0_u1_u1_n138 ) , .C2( u0_u1_u1_n139 ) , .B( u0_u1_u1_n145 ) , .C1( u0_u1_u1_n147 ) );
  NAND2_X1 u0_u1_u1_U50 (.ZN( u0_u1_u1_n129 ) , .A2( u0_u1_u1_n95 ) , .A1( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U51 (.A1( u0_u1_u1_n102 ) , .ZN( u0_u1_u1_n154 ) , .A2( u0_u1_u1_n99 ) );
  NAND2_X1 u0_u1_u1_U52 (.A2( u0_u1_u1_n100 ) , .ZN( u0_u1_u1_n135 ) , .A1( u0_u1_u1_n99 ) );
  AOI21_X1 u0_u1_u1_U53 (.A( u0_u1_u1_n152 ) , .B2( u0_u1_u1_n153 ) , .B1( u0_u1_u1_n154 ) , .ZN( u0_u1_u1_n158 ) );
  INV_X1 u0_u1_u1_U54 (.A( u0_u1_u1_n160 ) , .ZN( u0_u1_u1_n175 ) );
  NAND2_X1 u0_u1_u1_U55 (.A1( u0_u1_u1_n100 ) , .ZN( u0_u1_u1_n116 ) , .A2( u0_u1_u1_n95 ) );
  NAND2_X1 u0_u1_u1_U56 (.A1( u0_u1_u1_n102 ) , .ZN( u0_u1_u1_n131 ) , .A2( u0_u1_u1_n95 ) );
  NAND2_X1 u0_u1_u1_U57 (.A2( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n121 ) , .A1( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U58 (.A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n153 ) , .A2( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U59 (.A2( u0_u1_u1_n104 ) , .A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n133 ) );
  AOI22_X1 u0_u1_u1_U6 (.B2( u0_u1_u1_n113 ) , .A2( u0_u1_u1_n114 ) , .ZN( u0_u1_u1_n125 ) , .A1( u0_u1_u1_n171 ) , .B1( u0_u1_u1_n173 ) );
  NAND2_X1 u0_u1_u1_U60 (.ZN( u0_u1_u1_n150 ) , .A2( u0_u1_u1_n98 ) , .A1( u0_u1_u1_n99 ) );
  NAND2_X1 u0_u1_u1_U61 (.A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n155 ) , .A2( u0_u1_u1_n95 ) );
  OAI21_X1 u0_u1_u1_U62 (.ZN( u0_u1_u1_n109 ) , .B1( u0_u1_u1_n129 ) , .B2( u0_u1_u1_n160 ) , .A( u0_u1_u1_n167 ) );
  NAND2_X1 u0_u1_u1_U63 (.A2( u0_u1_u1_n100 ) , .A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n120 ) );
  NAND2_X1 u0_u1_u1_U64 (.A1( u0_u1_u1_n102 ) , .A2( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n115 ) );
  NAND2_X1 u0_u1_u1_U65 (.A2( u0_u1_u1_n100 ) , .A1( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n151 ) );
  NAND2_X1 u0_u1_u1_U66 (.A2( u0_u1_u1_n103 ) , .A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n161 ) );
  INV_X1 u0_u1_u1_U67 (.A( u0_u1_u1_n152 ) , .ZN( u0_u1_u1_n173 ) );
  INV_X1 u0_u1_u1_U68 (.A( u0_u1_u1_n128 ) , .ZN( u0_u1_u1_n172 ) );
  NAND2_X1 u0_u1_u1_U69 (.A2( u0_u1_u1_n102 ) , .A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n123 ) );
  NAND2_X1 u0_u1_u1_U7 (.ZN( u0_u1_u1_n114 ) , .A1( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n156 ) );
  NOR2_X1 u0_u1_u1_U70 (.A2( u0_u1_X_7 ) , .A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n95 ) );
  NOR2_X1 u0_u1_u1_U71 (.A1( u0_u1_X_12 ) , .A2( u0_u1_X_9 ) , .ZN( u0_u1_u1_n100 ) );
  NOR2_X1 u0_u1_u1_U72 (.A2( u0_u1_X_8 ) , .A1( u0_u1_u1_n177 ) , .ZN( u0_u1_u1_n99 ) );
  NOR2_X1 u0_u1_u1_U73 (.A2( u0_u1_X_12 ) , .ZN( u0_u1_u1_n102 ) , .A1( u0_u1_u1_n176 ) );
  NOR2_X1 u0_u1_u1_U74 (.A2( u0_u1_X_9 ) , .ZN( u0_u1_u1_n105 ) , .A1( u0_u1_u1_n168 ) );
  NAND2_X1 u0_u1_u1_U75 (.A1( u0_u1_X_10 ) , .ZN( u0_u1_u1_n160 ) , .A2( u0_u1_u1_n169 ) );
  NAND2_X1 u0_u1_u1_U76 (.A2( u0_u1_X_10 ) , .A1( u0_u1_X_11 ) , .ZN( u0_u1_u1_n152 ) );
  NAND2_X1 u0_u1_u1_U77 (.A1( u0_u1_X_11 ) , .ZN( u0_u1_u1_n128 ) , .A2( u0_u1_u1_n170 ) );
  AND2_X1 u0_u1_u1_U78 (.A2( u0_u1_X_7 ) , .A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n104 ) );
  AND2_X1 u0_u1_u1_U79 (.A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n103 ) , .A2( u0_u1_u1_n177 ) );
  AOI22_X1 u0_u1_u1_U8 (.B2( u0_u1_u1_n136 ) , .A2( u0_u1_u1_n137 ) , .ZN( u0_u1_u1_n143 ) , .A1( u0_u1_u1_n171 ) , .B1( u0_u1_u1_n173 ) );
  INV_X1 u0_u1_u1_U80 (.A( u0_u1_X_10 ) , .ZN( u0_u1_u1_n170 ) );
  INV_X1 u0_u1_u1_U81 (.A( u0_u1_X_9 ) , .ZN( u0_u1_u1_n176 ) );
  INV_X1 u0_u1_u1_U82 (.A( u0_u1_X_11 ) , .ZN( u0_u1_u1_n169 ) );
  INV_X1 u0_u1_u1_U83 (.A( u0_u1_X_12 ) , .ZN( u0_u1_u1_n168 ) );
  INV_X1 u0_u1_u1_U84 (.A( u0_u1_X_7 ) , .ZN( u0_u1_u1_n177 ) );
  NAND4_X1 u0_u1_u1_U85 (.ZN( u0_out1_28 ) , .A4( u0_u1_u1_n124 ) , .A3( u0_u1_u1_n125 ) , .A2( u0_u1_u1_n126 ) , .A1( u0_u1_u1_n127 ) );
  OAI21_X1 u0_u1_u1_U86 (.ZN( u0_u1_u1_n127 ) , .B2( u0_u1_u1_n139 ) , .B1( u0_u1_u1_n175 ) , .A( u0_u1_u1_n183 ) );
  OAI21_X1 u0_u1_u1_U87 (.ZN( u0_u1_u1_n126 ) , .B2( u0_u1_u1_n140 ) , .A( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n178 ) );
  NAND4_X1 u0_u1_u1_U88 (.ZN( u0_out1_18 ) , .A4( u0_u1_u1_n165 ) , .A3( u0_u1_u1_n166 ) , .A1( u0_u1_u1_n167 ) , .A2( u0_u1_u1_n186 ) );
  AOI22_X1 u0_u1_u1_U89 (.B2( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n147 ) , .A2( u0_u1_u1_n148 ) , .ZN( u0_u1_u1_n166 ) , .A1( u0_u1_u1_n172 ) );
  INV_X1 u0_u1_u1_U9 (.A( u0_u1_u1_n147 ) , .ZN( u0_u1_u1_n181 ) );
  INV_X1 u0_u1_u1_U90 (.A( u0_u1_u1_n145 ) , .ZN( u0_u1_u1_n186 ) );
  NAND4_X1 u0_u1_u1_U91 (.ZN( u0_out1_2 ) , .A4( u0_u1_u1_n142 ) , .A3( u0_u1_u1_n143 ) , .A2( u0_u1_u1_n144 ) , .A1( u0_u1_u1_n179 ) );
  INV_X1 u0_u1_u1_U92 (.A( u0_u1_u1_n130 ) , .ZN( u0_u1_u1_n179 ) );
  OAI21_X1 u0_u1_u1_U93 (.B2( u0_u1_u1_n132 ) , .ZN( u0_u1_u1_n144 ) , .A( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n180 ) );
  OR4_X1 u0_u1_u1_U94 (.ZN( u0_out1_13 ) , .A4( u0_u1_u1_n108 ) , .A3( u0_u1_u1_n109 ) , .A2( u0_u1_u1_n110 ) , .A1( u0_u1_u1_n111 ) );
  AOI21_X1 u0_u1_u1_U95 (.ZN( u0_u1_u1_n111 ) , .A( u0_u1_u1_n128 ) , .B2( u0_u1_u1_n131 ) , .B1( u0_u1_u1_n135 ) );
  AOI21_X1 u0_u1_u1_U96 (.ZN( u0_u1_u1_n110 ) , .A( u0_u1_u1_n116 ) , .B1( u0_u1_u1_n152 ) , .B2( u0_u1_u1_n160 ) );
  NAND3_X1 u0_u1_u1_U97 (.A3( u0_u1_u1_n149 ) , .A2( u0_u1_u1_n150 ) , .A1( u0_u1_u1_n151 ) , .ZN( u0_u1_u1_n164 ) );
  NAND3_X1 u0_u1_u1_U98 (.A3( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n135 ) , .ZN( u0_u1_u1_n136 ) , .A1( u0_u1_u1_n151 ) );
  NAND3_X1 u0_u1_u1_U99 (.A1( u0_u1_u1_n133 ) , .ZN( u0_u1_u1_n137 ) , .A2( u0_u1_u1_n154 ) , .A3( u0_u1_u1_n181 ) );
  OAI22_X1 u0_u1_u4_U10 (.B2( u0_u1_u4_n135 ) , .ZN( u0_u1_u4_n137 ) , .B1( u0_u1_u4_n153 ) , .A1( u0_u1_u4_n155 ) , .A2( u0_u1_u4_n171 ) );
  AND3_X1 u0_u1_u4_U11 (.A2( u0_u1_u4_n134 ) , .ZN( u0_u1_u4_n135 ) , .A3( u0_u1_u4_n145 ) , .A1( u0_u1_u4_n157 ) );
  NAND2_X1 u0_u1_u4_U12 (.ZN( u0_u1_u4_n132 ) , .A2( u0_u1_u4_n170 ) , .A1( u0_u1_u4_n173 ) );
  AOI21_X1 u0_u1_u4_U13 (.B2( u0_u1_u4_n160 ) , .B1( u0_u1_u4_n161 ) , .ZN( u0_u1_u4_n162 ) , .A( u0_u1_u4_n170 ) );
  AOI21_X1 u0_u1_u4_U14 (.ZN( u0_u1_u4_n107 ) , .B2( u0_u1_u4_n143 ) , .A( u0_u1_u4_n174 ) , .B1( u0_u1_u4_n184 ) );
  AOI21_X1 u0_u1_u4_U15 (.B2( u0_u1_u4_n158 ) , .B1( u0_u1_u4_n159 ) , .ZN( u0_u1_u4_n163 ) , .A( u0_u1_u4_n174 ) );
  AOI21_X1 u0_u1_u4_U16 (.A( u0_u1_u4_n153 ) , .B2( u0_u1_u4_n154 ) , .B1( u0_u1_u4_n155 ) , .ZN( u0_u1_u4_n165 ) );
  AOI21_X1 u0_u1_u4_U17 (.A( u0_u1_u4_n156 ) , .B2( u0_u1_u4_n157 ) , .ZN( u0_u1_u4_n164 ) , .B1( u0_u1_u4_n184 ) );
  INV_X1 u0_u1_u4_U18 (.A( u0_u1_u4_n138 ) , .ZN( u0_u1_u4_n170 ) );
  AND2_X1 u0_u1_u4_U19 (.A2( u0_u1_u4_n120 ) , .ZN( u0_u1_u4_n155 ) , .A1( u0_u1_u4_n160 ) );
  INV_X1 u0_u1_u4_U20 (.A( u0_u1_u4_n156 ) , .ZN( u0_u1_u4_n175 ) );
  NAND2_X1 u0_u1_u4_U21 (.A2( u0_u1_u4_n118 ) , .ZN( u0_u1_u4_n131 ) , .A1( u0_u1_u4_n147 ) );
  NAND2_X1 u0_u1_u4_U22 (.A1( u0_u1_u4_n119 ) , .A2( u0_u1_u4_n120 ) , .ZN( u0_u1_u4_n130 ) );
  NAND2_X1 u0_u1_u4_U23 (.ZN( u0_u1_u4_n117 ) , .A2( u0_u1_u4_n118 ) , .A1( u0_u1_u4_n148 ) );
  NAND2_X1 u0_u1_u4_U24 (.ZN( u0_u1_u4_n129 ) , .A1( u0_u1_u4_n134 ) , .A2( u0_u1_u4_n148 ) );
  AND3_X1 u0_u1_u4_U25 (.A1( u0_u1_u4_n119 ) , .A2( u0_u1_u4_n143 ) , .A3( u0_u1_u4_n154 ) , .ZN( u0_u1_u4_n161 ) );
  AND2_X1 u0_u1_u4_U26 (.A1( u0_u1_u4_n145 ) , .A2( u0_u1_u4_n147 ) , .ZN( u0_u1_u4_n159 ) );
  OR3_X1 u0_u1_u4_U27 (.A3( u0_u1_u4_n114 ) , .A2( u0_u1_u4_n115 ) , .A1( u0_u1_u4_n116 ) , .ZN( u0_u1_u4_n136 ) );
  AOI21_X1 u0_u1_u4_U28 (.A( u0_u1_u4_n113 ) , .ZN( u0_u1_u4_n116 ) , .B2( u0_u1_u4_n173 ) , .B1( u0_u1_u4_n174 ) );
  AOI21_X1 u0_u1_u4_U29 (.ZN( u0_u1_u4_n115 ) , .B2( u0_u1_u4_n145 ) , .B1( u0_u1_u4_n146 ) , .A( u0_u1_u4_n156 ) );
  NOR2_X1 u0_u1_u4_U3 (.ZN( u0_u1_u4_n121 ) , .A1( u0_u1_u4_n181 ) , .A2( u0_u1_u4_n182 ) );
  OAI22_X1 u0_u1_u4_U30 (.ZN( u0_u1_u4_n114 ) , .A2( u0_u1_u4_n121 ) , .B1( u0_u1_u4_n160 ) , .B2( u0_u1_u4_n170 ) , .A1( u0_u1_u4_n171 ) );
  INV_X1 u0_u1_u4_U31 (.A( u0_u1_u4_n158 ) , .ZN( u0_u1_u4_n182 ) );
  INV_X1 u0_u1_u4_U32 (.ZN( u0_u1_u4_n181 ) , .A( u0_u1_u4_n96 ) );
  INV_X1 u0_u1_u4_U33 (.A( u0_u1_u4_n144 ) , .ZN( u0_u1_u4_n179 ) );
  INV_X1 u0_u1_u4_U34 (.A( u0_u1_u4_n157 ) , .ZN( u0_u1_u4_n178 ) );
  NAND2_X1 u0_u1_u4_U35 (.A2( u0_u1_u4_n154 ) , .A1( u0_u1_u4_n96 ) , .ZN( u0_u1_u4_n97 ) );
  INV_X1 u0_u1_u4_U36 (.ZN( u0_u1_u4_n186 ) , .A( u0_u1_u4_n95 ) );
  OAI221_X1 u0_u1_u4_U37 (.C1( u0_u1_u4_n134 ) , .B1( u0_u1_u4_n158 ) , .B2( u0_u1_u4_n171 ) , .C2( u0_u1_u4_n173 ) , .A( u0_u1_u4_n94 ) , .ZN( u0_u1_u4_n95 ) );
  AOI222_X1 u0_u1_u4_U38 (.B2( u0_u1_u4_n132 ) , .A1( u0_u1_u4_n138 ) , .C2( u0_u1_u4_n175 ) , .A2( u0_u1_u4_n179 ) , .C1( u0_u1_u4_n181 ) , .B1( u0_u1_u4_n185 ) , .ZN( u0_u1_u4_n94 ) );
  INV_X1 u0_u1_u4_U39 (.A( u0_u1_u4_n113 ) , .ZN( u0_u1_u4_n185 ) );
  INV_X1 u0_u1_u4_U4 (.A( u0_u1_u4_n117 ) , .ZN( u0_u1_u4_n184 ) );
  INV_X1 u0_u1_u4_U40 (.A( u0_u1_u4_n143 ) , .ZN( u0_u1_u4_n183 ) );
  NOR2_X1 u0_u1_u4_U41 (.ZN( u0_u1_u4_n138 ) , .A1( u0_u1_u4_n168 ) , .A2( u0_u1_u4_n169 ) );
  NOR2_X1 u0_u1_u4_U42 (.A1( u0_u1_u4_n150 ) , .A2( u0_u1_u4_n152 ) , .ZN( u0_u1_u4_n153 ) );
  NOR2_X1 u0_u1_u4_U43 (.A2( u0_u1_u4_n128 ) , .A1( u0_u1_u4_n138 ) , .ZN( u0_u1_u4_n156 ) );
  AOI22_X1 u0_u1_u4_U44 (.B2( u0_u1_u4_n122 ) , .A1( u0_u1_u4_n123 ) , .ZN( u0_u1_u4_n124 ) , .B1( u0_u1_u4_n128 ) , .A2( u0_u1_u4_n172 ) );
  NAND2_X1 u0_u1_u4_U45 (.A2( u0_u1_u4_n120 ) , .ZN( u0_u1_u4_n123 ) , .A1( u0_u1_u4_n161 ) );
  INV_X1 u0_u1_u4_U46 (.A( u0_u1_u4_n153 ) , .ZN( u0_u1_u4_n172 ) );
  AOI22_X1 u0_u1_u4_U47 (.B2( u0_u1_u4_n132 ) , .A2( u0_u1_u4_n133 ) , .ZN( u0_u1_u4_n140 ) , .A1( u0_u1_u4_n150 ) , .B1( u0_u1_u4_n179 ) );
  NAND2_X1 u0_u1_u4_U48 (.ZN( u0_u1_u4_n133 ) , .A2( u0_u1_u4_n146 ) , .A1( u0_u1_u4_n154 ) );
  NAND2_X1 u0_u1_u4_U49 (.A1( u0_u1_u4_n103 ) , .ZN( u0_u1_u4_n154 ) , .A2( u0_u1_u4_n98 ) );
  NOR4_X1 u0_u1_u4_U5 (.A4( u0_u1_u4_n106 ) , .A3( u0_u1_u4_n107 ) , .A2( u0_u1_u4_n108 ) , .A1( u0_u1_u4_n109 ) , .ZN( u0_u1_u4_n110 ) );
  NAND2_X1 u0_u1_u4_U50 (.A1( u0_u1_u4_n101 ) , .ZN( u0_u1_u4_n158 ) , .A2( u0_u1_u4_n99 ) );
  AOI21_X1 u0_u1_u4_U51 (.ZN( u0_u1_u4_n127 ) , .A( u0_u1_u4_n136 ) , .B2( u0_u1_u4_n150 ) , .B1( u0_u1_u4_n180 ) );
  INV_X1 u0_u1_u4_U52 (.A( u0_u1_u4_n160 ) , .ZN( u0_u1_u4_n180 ) );
  NAND2_X1 u0_u1_u4_U53 (.A2( u0_u1_u4_n104 ) , .A1( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n146 ) );
  NAND2_X1 u0_u1_u4_U54 (.A2( u0_u1_u4_n101 ) , .A1( u0_u1_u4_n102 ) , .ZN( u0_u1_u4_n160 ) );
  NAND2_X1 u0_u1_u4_U55 (.ZN( u0_u1_u4_n134 ) , .A1( u0_u1_u4_n98 ) , .A2( u0_u1_u4_n99 ) );
  NAND2_X1 u0_u1_u4_U56 (.A1( u0_u1_u4_n103 ) , .A2( u0_u1_u4_n104 ) , .ZN( u0_u1_u4_n143 ) );
  NAND2_X1 u0_u1_u4_U57 (.A2( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n145 ) , .A1( u0_u1_u4_n98 ) );
  NAND2_X1 u0_u1_u4_U58 (.A1( u0_u1_u4_n100 ) , .A2( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n120 ) );
  NAND2_X1 u0_u1_u4_U59 (.A1( u0_u1_u4_n102 ) , .A2( u0_u1_u4_n104 ) , .ZN( u0_u1_u4_n148 ) );
  AOI21_X1 u0_u1_u4_U6 (.ZN( u0_u1_u4_n106 ) , .B2( u0_u1_u4_n146 ) , .B1( u0_u1_u4_n158 ) , .A( u0_u1_u4_n170 ) );
  NAND2_X1 u0_u1_u4_U60 (.A2( u0_u1_u4_n100 ) , .A1( u0_u1_u4_n103 ) , .ZN( u0_u1_u4_n157 ) );
  INV_X1 u0_u1_u4_U61 (.A( u0_u1_u4_n150 ) , .ZN( u0_u1_u4_n173 ) );
  INV_X1 u0_u1_u4_U62 (.A( u0_u1_u4_n152 ) , .ZN( u0_u1_u4_n171 ) );
  NAND2_X1 u0_u1_u4_U63 (.A1( u0_u1_u4_n100 ) , .ZN( u0_u1_u4_n118 ) , .A2( u0_u1_u4_n99 ) );
  NAND2_X1 u0_u1_u4_U64 (.A2( u0_u1_u4_n100 ) , .A1( u0_u1_u4_n102 ) , .ZN( u0_u1_u4_n144 ) );
  NAND2_X1 u0_u1_u4_U65 (.A2( u0_u1_u4_n101 ) , .A1( u0_u1_u4_n105 ) , .ZN( u0_u1_u4_n96 ) );
  INV_X1 u0_u1_u4_U66 (.A( u0_u1_u4_n128 ) , .ZN( u0_u1_u4_n174 ) );
  NAND2_X1 u0_u1_u4_U67 (.A2( u0_u1_u4_n102 ) , .ZN( u0_u1_u4_n119 ) , .A1( u0_u1_u4_n98 ) );
  NAND2_X1 u0_u1_u4_U68 (.A2( u0_u1_u4_n101 ) , .A1( u0_u1_u4_n103 ) , .ZN( u0_u1_u4_n147 ) );
  NAND2_X1 u0_u1_u4_U69 (.A2( u0_u1_u4_n104 ) , .ZN( u0_u1_u4_n113 ) , .A1( u0_u1_u4_n99 ) );
  AOI21_X1 u0_u1_u4_U7 (.ZN( u0_u1_u4_n108 ) , .B2( u0_u1_u4_n134 ) , .B1( u0_u1_u4_n155 ) , .A( u0_u1_u4_n156 ) );
  NOR2_X1 u0_u1_u4_U70 (.A2( u0_u1_X_28 ) , .ZN( u0_u1_u4_n150 ) , .A1( u0_u1_u4_n168 ) );
  NOR2_X1 u0_u1_u4_U71 (.A2( u0_u1_X_29 ) , .ZN( u0_u1_u4_n152 ) , .A1( u0_u1_u4_n169 ) );
  NOR2_X1 u0_u1_u4_U72 (.A2( u0_u1_X_30 ) , .ZN( u0_u1_u4_n105 ) , .A1( u0_u1_u4_n176 ) );
  NOR2_X1 u0_u1_u4_U73 (.A2( u0_u1_X_26 ) , .ZN( u0_u1_u4_n100 ) , .A1( u0_u1_u4_n177 ) );
  NOR2_X1 u0_u1_u4_U74 (.A2( u0_u1_X_28 ) , .A1( u0_u1_X_29 ) , .ZN( u0_u1_u4_n128 ) );
  NOR2_X1 u0_u1_u4_U75 (.A2( u0_u1_X_27 ) , .A1( u0_u1_X_30 ) , .ZN( u0_u1_u4_n102 ) );
  NOR2_X1 u0_u1_u4_U76 (.A2( u0_u1_X_25 ) , .A1( u0_u1_X_26 ) , .ZN( u0_u1_u4_n98 ) );
  AND2_X1 u0_u1_u4_U77 (.A2( u0_u1_X_25 ) , .A1( u0_u1_X_26 ) , .ZN( u0_u1_u4_n104 ) );
  AND2_X1 u0_u1_u4_U78 (.A1( u0_u1_X_30 ) , .A2( u0_u1_u4_n176 ) , .ZN( u0_u1_u4_n99 ) );
  AND2_X1 u0_u1_u4_U79 (.A1( u0_u1_X_26 ) , .ZN( u0_u1_u4_n101 ) , .A2( u0_u1_u4_n177 ) );
  AOI21_X1 u0_u1_u4_U8 (.ZN( u0_u1_u4_n109 ) , .A( u0_u1_u4_n153 ) , .B1( u0_u1_u4_n159 ) , .B2( u0_u1_u4_n184 ) );
  AND2_X1 u0_u1_u4_U80 (.A1( u0_u1_X_27 ) , .A2( u0_u1_X_30 ) , .ZN( u0_u1_u4_n103 ) );
  INV_X1 u0_u1_u4_U81 (.A( u0_u1_X_28 ) , .ZN( u0_u1_u4_n169 ) );
  INV_X1 u0_u1_u4_U82 (.A( u0_u1_X_29 ) , .ZN( u0_u1_u4_n168 ) );
  INV_X1 u0_u1_u4_U83 (.A( u0_u1_X_25 ) , .ZN( u0_u1_u4_n177 ) );
  INV_X1 u0_u1_u4_U84 (.A( u0_u1_X_27 ) , .ZN( u0_u1_u4_n176 ) );
  NAND4_X1 u0_u1_u4_U85 (.ZN( u0_out1_25 ) , .A4( u0_u1_u4_n139 ) , .A3( u0_u1_u4_n140 ) , .A2( u0_u1_u4_n141 ) , .A1( u0_u1_u4_n142 ) );
  OAI21_X1 u0_u1_u4_U86 (.A( u0_u1_u4_n128 ) , .B2( u0_u1_u4_n129 ) , .B1( u0_u1_u4_n130 ) , .ZN( u0_u1_u4_n142 ) );
  OAI21_X1 u0_u1_u4_U87 (.B2( u0_u1_u4_n131 ) , .ZN( u0_u1_u4_n141 ) , .A( u0_u1_u4_n175 ) , .B1( u0_u1_u4_n183 ) );
  NAND4_X1 u0_u1_u4_U88 (.ZN( u0_out1_14 ) , .A4( u0_u1_u4_n124 ) , .A3( u0_u1_u4_n125 ) , .A2( u0_u1_u4_n126 ) , .A1( u0_u1_u4_n127 ) );
  AOI22_X1 u0_u1_u4_U89 (.B2( u0_u1_u4_n117 ) , .ZN( u0_u1_u4_n126 ) , .A1( u0_u1_u4_n129 ) , .B1( u0_u1_u4_n152 ) , .A2( u0_u1_u4_n175 ) );
  AOI211_X1 u0_u1_u4_U9 (.B( u0_u1_u4_n136 ) , .A( u0_u1_u4_n137 ) , .C2( u0_u1_u4_n138 ) , .ZN( u0_u1_u4_n139 ) , .C1( u0_u1_u4_n182 ) );
  AOI22_X1 u0_u1_u4_U90 (.ZN( u0_u1_u4_n125 ) , .B2( u0_u1_u4_n131 ) , .A2( u0_u1_u4_n132 ) , .B1( u0_u1_u4_n138 ) , .A1( u0_u1_u4_n178 ) );
  NAND4_X1 u0_u1_u4_U91 (.ZN( u0_out1_8 ) , .A4( u0_u1_u4_n110 ) , .A3( u0_u1_u4_n111 ) , .A2( u0_u1_u4_n112 ) , .A1( u0_u1_u4_n186 ) );
  NAND2_X1 u0_u1_u4_U92 (.ZN( u0_u1_u4_n112 ) , .A2( u0_u1_u4_n130 ) , .A1( u0_u1_u4_n150 ) );
  AOI22_X1 u0_u1_u4_U93 (.ZN( u0_u1_u4_n111 ) , .B2( u0_u1_u4_n132 ) , .A1( u0_u1_u4_n152 ) , .B1( u0_u1_u4_n178 ) , .A2( u0_u1_u4_n97 ) );
  AOI22_X1 u0_u1_u4_U94 (.B2( u0_u1_u4_n149 ) , .B1( u0_u1_u4_n150 ) , .A2( u0_u1_u4_n151 ) , .A1( u0_u1_u4_n152 ) , .ZN( u0_u1_u4_n167 ) );
  NOR4_X1 u0_u1_u4_U95 (.A4( u0_u1_u4_n162 ) , .A3( u0_u1_u4_n163 ) , .A2( u0_u1_u4_n164 ) , .A1( u0_u1_u4_n165 ) , .ZN( u0_u1_u4_n166 ) );
  NAND3_X1 u0_u1_u4_U96 (.ZN( u0_out1_3 ) , .A3( u0_u1_u4_n166 ) , .A1( u0_u1_u4_n167 ) , .A2( u0_u1_u4_n186 ) );
  NAND3_X1 u0_u1_u4_U97 (.A3( u0_u1_u4_n146 ) , .A2( u0_u1_u4_n147 ) , .A1( u0_u1_u4_n148 ) , .ZN( u0_u1_u4_n149 ) );
  NAND3_X1 u0_u1_u4_U98 (.A3( u0_u1_u4_n143 ) , .A2( u0_u1_u4_n144 ) , .A1( u0_u1_u4_n145 ) , .ZN( u0_u1_u4_n151 ) );
  NAND3_X1 u0_u1_u4_U99 (.A3( u0_u1_u4_n121 ) , .ZN( u0_u1_u4_n122 ) , .A2( u0_u1_u4_n144 ) , .A1( u0_u1_u4_n154 ) );
  INV_X1 u0_u1_u5_U10 (.A( u0_u1_u5_n121 ) , .ZN( u0_u1_u5_n177 ) );
  NOR3_X1 u0_u1_u5_U100 (.A3( u0_u1_u5_n141 ) , .A1( u0_u1_u5_n142 ) , .ZN( u0_u1_u5_n143 ) , .A2( u0_u1_u5_n191 ) );
  NAND4_X1 u0_u1_u5_U101 (.ZN( u0_out1_4 ) , .A4( u0_u1_u5_n112 ) , .A2( u0_u1_u5_n113 ) , .A1( u0_u1_u5_n114 ) , .A3( u0_u1_u5_n195 ) );
  AOI211_X1 u0_u1_u5_U102 (.A( u0_u1_u5_n110 ) , .C1( u0_u1_u5_n111 ) , .ZN( u0_u1_u5_n112 ) , .B( u0_u1_u5_n118 ) , .C2( u0_u1_u5_n177 ) );
  AOI222_X1 u0_u1_u5_U103 (.ZN( u0_u1_u5_n113 ) , .A1( u0_u1_u5_n131 ) , .C1( u0_u1_u5_n148 ) , .B2( u0_u1_u5_n174 ) , .C2( u0_u1_u5_n178 ) , .A2( u0_u1_u5_n179 ) , .B1( u0_u1_u5_n99 ) );
  NAND3_X1 u0_u1_u5_U104 (.A2( u0_u1_u5_n154 ) , .A3( u0_u1_u5_n158 ) , .A1( u0_u1_u5_n161 ) , .ZN( u0_u1_u5_n99 ) );
  NOR2_X1 u0_u1_u5_U11 (.ZN( u0_u1_u5_n160 ) , .A2( u0_u1_u5_n173 ) , .A1( u0_u1_u5_n177 ) );
  INV_X1 u0_u1_u5_U12 (.A( u0_u1_u5_n150 ) , .ZN( u0_u1_u5_n174 ) );
  AOI21_X1 u0_u1_u5_U13 (.A( u0_u1_u5_n160 ) , .B2( u0_u1_u5_n161 ) , .ZN( u0_u1_u5_n162 ) , .B1( u0_u1_u5_n192 ) );
  INV_X1 u0_u1_u5_U14 (.A( u0_u1_u5_n159 ) , .ZN( u0_u1_u5_n192 ) );
  AOI21_X1 u0_u1_u5_U15 (.A( u0_u1_u5_n156 ) , .B2( u0_u1_u5_n157 ) , .B1( u0_u1_u5_n158 ) , .ZN( u0_u1_u5_n163 ) );
  AOI21_X1 u0_u1_u5_U16 (.B2( u0_u1_u5_n139 ) , .B1( u0_u1_u5_n140 ) , .ZN( u0_u1_u5_n141 ) , .A( u0_u1_u5_n150 ) );
  OAI21_X1 u0_u1_u5_U17 (.A( u0_u1_u5_n133 ) , .B2( u0_u1_u5_n134 ) , .B1( u0_u1_u5_n135 ) , .ZN( u0_u1_u5_n142 ) );
  OAI21_X1 u0_u1_u5_U18 (.ZN( u0_u1_u5_n133 ) , .B2( u0_u1_u5_n147 ) , .A( u0_u1_u5_n173 ) , .B1( u0_u1_u5_n188 ) );
  NAND2_X1 u0_u1_u5_U19 (.A2( u0_u1_u5_n119 ) , .A1( u0_u1_u5_n123 ) , .ZN( u0_u1_u5_n137 ) );
  INV_X1 u0_u1_u5_U20 (.A( u0_u1_u5_n155 ) , .ZN( u0_u1_u5_n194 ) );
  NAND2_X1 u0_u1_u5_U21 (.A1( u0_u1_u5_n121 ) , .ZN( u0_u1_u5_n132 ) , .A2( u0_u1_u5_n172 ) );
  NAND2_X1 u0_u1_u5_U22 (.A2( u0_u1_u5_n122 ) , .ZN( u0_u1_u5_n136 ) , .A1( u0_u1_u5_n154 ) );
  NAND2_X1 u0_u1_u5_U23 (.A2( u0_u1_u5_n119 ) , .A1( u0_u1_u5_n120 ) , .ZN( u0_u1_u5_n159 ) );
  INV_X1 u0_u1_u5_U24 (.A( u0_u1_u5_n156 ) , .ZN( u0_u1_u5_n175 ) );
  INV_X1 u0_u1_u5_U25 (.A( u0_u1_u5_n158 ) , .ZN( u0_u1_u5_n188 ) );
  INV_X1 u0_u1_u5_U26 (.A( u0_u1_u5_n152 ) , .ZN( u0_u1_u5_n179 ) );
  INV_X1 u0_u1_u5_U27 (.A( u0_u1_u5_n140 ) , .ZN( u0_u1_u5_n182 ) );
  INV_X1 u0_u1_u5_U28 (.A( u0_u1_u5_n151 ) , .ZN( u0_u1_u5_n183 ) );
  INV_X1 u0_u1_u5_U29 (.A( u0_u1_u5_n123 ) , .ZN( u0_u1_u5_n185 ) );
  NOR2_X1 u0_u1_u5_U3 (.ZN( u0_u1_u5_n134 ) , .A1( u0_u1_u5_n183 ) , .A2( u0_u1_u5_n190 ) );
  INV_X1 u0_u1_u5_U30 (.A( u0_u1_u5_n161 ) , .ZN( u0_u1_u5_n184 ) );
  INV_X1 u0_u1_u5_U31 (.A( u0_u1_u5_n139 ) , .ZN( u0_u1_u5_n189 ) );
  INV_X1 u0_u1_u5_U32 (.A( u0_u1_u5_n157 ) , .ZN( u0_u1_u5_n190 ) );
  INV_X1 u0_u1_u5_U33 (.A( u0_u1_u5_n120 ) , .ZN( u0_u1_u5_n193 ) );
  NAND2_X1 u0_u1_u5_U34 (.ZN( u0_u1_u5_n111 ) , .A1( u0_u1_u5_n140 ) , .A2( u0_u1_u5_n155 ) );
  INV_X1 u0_u1_u5_U35 (.A( u0_u1_u5_n117 ) , .ZN( u0_u1_u5_n196 ) );
  OAI221_X1 u0_u1_u5_U36 (.A( u0_u1_u5_n116 ) , .ZN( u0_u1_u5_n117 ) , .B2( u0_u1_u5_n119 ) , .C1( u0_u1_u5_n153 ) , .C2( u0_u1_u5_n158 ) , .B1( u0_u1_u5_n172 ) );
  AOI222_X1 u0_u1_u5_U37 (.ZN( u0_u1_u5_n116 ) , .B2( u0_u1_u5_n145 ) , .C1( u0_u1_u5_n148 ) , .A2( u0_u1_u5_n174 ) , .C2( u0_u1_u5_n177 ) , .B1( u0_u1_u5_n187 ) , .A1( u0_u1_u5_n193 ) );
  INV_X1 u0_u1_u5_U38 (.A( u0_u1_u5_n115 ) , .ZN( u0_u1_u5_n187 ) );
  NOR2_X1 u0_u1_u5_U39 (.ZN( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n170 ) , .A2( u0_u1_u5_n180 ) );
  INV_X1 u0_u1_u5_U4 (.A( u0_u1_u5_n138 ) , .ZN( u0_u1_u5_n191 ) );
  AOI22_X1 u0_u1_u5_U40 (.B2( u0_u1_u5_n131 ) , .A2( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n169 ) , .B1( u0_u1_u5_n174 ) , .A1( u0_u1_u5_n185 ) );
  NOR2_X1 u0_u1_u5_U41 (.A1( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n150 ) , .A2( u0_u1_u5_n173 ) );
  AOI21_X1 u0_u1_u5_U42 (.A( u0_u1_u5_n118 ) , .B2( u0_u1_u5_n145 ) , .ZN( u0_u1_u5_n168 ) , .B1( u0_u1_u5_n186 ) );
  INV_X1 u0_u1_u5_U43 (.A( u0_u1_u5_n122 ) , .ZN( u0_u1_u5_n186 ) );
  NOR2_X1 u0_u1_u5_U44 (.A1( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n152 ) , .A2( u0_u1_u5_n176 ) );
  NOR2_X1 u0_u1_u5_U45 (.A1( u0_u1_u5_n115 ) , .ZN( u0_u1_u5_n118 ) , .A2( u0_u1_u5_n153 ) );
  NOR2_X1 u0_u1_u5_U46 (.A2( u0_u1_u5_n145 ) , .ZN( u0_u1_u5_n156 ) , .A1( u0_u1_u5_n174 ) );
  NOR2_X1 u0_u1_u5_U47 (.ZN( u0_u1_u5_n121 ) , .A2( u0_u1_u5_n145 ) , .A1( u0_u1_u5_n176 ) );
  AOI22_X1 u0_u1_u5_U48 (.ZN( u0_u1_u5_n114 ) , .A2( u0_u1_u5_n137 ) , .A1( u0_u1_u5_n145 ) , .B2( u0_u1_u5_n175 ) , .B1( u0_u1_u5_n193 ) );
  OAI211_X1 u0_u1_u5_U49 (.B( u0_u1_u5_n124 ) , .A( u0_u1_u5_n125 ) , .C2( u0_u1_u5_n126 ) , .C1( u0_u1_u5_n127 ) , .ZN( u0_u1_u5_n128 ) );
  OAI21_X1 u0_u1_u5_U5 (.B2( u0_u1_u5_n136 ) , .B1( u0_u1_u5_n137 ) , .ZN( u0_u1_u5_n138 ) , .A( u0_u1_u5_n177 ) );
  OAI21_X1 u0_u1_u5_U50 (.ZN( u0_u1_u5_n124 ) , .A( u0_u1_u5_n177 ) , .B2( u0_u1_u5_n183 ) , .B1( u0_u1_u5_n189 ) );
  NOR3_X1 u0_u1_u5_U51 (.ZN( u0_u1_u5_n127 ) , .A1( u0_u1_u5_n136 ) , .A3( u0_u1_u5_n148 ) , .A2( u0_u1_u5_n182 ) );
  OAI21_X1 u0_u1_u5_U52 (.ZN( u0_u1_u5_n125 ) , .A( u0_u1_u5_n174 ) , .B2( u0_u1_u5_n185 ) , .B1( u0_u1_u5_n190 ) );
  AOI21_X1 u0_u1_u5_U53 (.A( u0_u1_u5_n153 ) , .B2( u0_u1_u5_n154 ) , .B1( u0_u1_u5_n155 ) , .ZN( u0_u1_u5_n164 ) );
  AOI21_X1 u0_u1_u5_U54 (.ZN( u0_u1_u5_n110 ) , .B1( u0_u1_u5_n122 ) , .B2( u0_u1_u5_n139 ) , .A( u0_u1_u5_n153 ) );
  INV_X1 u0_u1_u5_U55 (.A( u0_u1_u5_n153 ) , .ZN( u0_u1_u5_n176 ) );
  INV_X1 u0_u1_u5_U56 (.A( u0_u1_u5_n126 ) , .ZN( u0_u1_u5_n173 ) );
  AND2_X1 u0_u1_u5_U57 (.A2( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n107 ) , .ZN( u0_u1_u5_n147 ) );
  AND2_X1 u0_u1_u5_U58 (.A2( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n108 ) , .ZN( u0_u1_u5_n148 ) );
  NAND2_X1 u0_u1_u5_U59 (.A1( u0_u1_u5_n105 ) , .A2( u0_u1_u5_n106 ) , .ZN( u0_u1_u5_n158 ) );
  INV_X1 u0_u1_u5_U6 (.A( u0_u1_u5_n135 ) , .ZN( u0_u1_u5_n178 ) );
  NAND2_X1 u0_u1_u5_U60 (.A2( u0_u1_u5_n108 ) , .A1( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n139 ) );
  NAND2_X1 u0_u1_u5_U61 (.A1( u0_u1_u5_n106 ) , .A2( u0_u1_u5_n108 ) , .ZN( u0_u1_u5_n119 ) );
  NAND2_X1 u0_u1_u5_U62 (.A2( u0_u1_u5_n103 ) , .A1( u0_u1_u5_n105 ) , .ZN( u0_u1_u5_n140 ) );
  NAND2_X1 u0_u1_u5_U63 (.A2( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n105 ) , .ZN( u0_u1_u5_n155 ) );
  NAND2_X1 u0_u1_u5_U64 (.A2( u0_u1_u5_n106 ) , .A1( u0_u1_u5_n107 ) , .ZN( u0_u1_u5_n122 ) );
  NAND2_X1 u0_u1_u5_U65 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n106 ) , .ZN( u0_u1_u5_n115 ) );
  NAND2_X1 u0_u1_u5_U66 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n103 ) , .ZN( u0_u1_u5_n161 ) );
  NAND2_X1 u0_u1_u5_U67 (.A1( u0_u1_u5_n105 ) , .A2( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n154 ) );
  INV_X1 u0_u1_u5_U68 (.A( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n172 ) );
  NAND2_X1 u0_u1_u5_U69 (.A1( u0_u1_u5_n103 ) , .A2( u0_u1_u5_n108 ) , .ZN( u0_u1_u5_n123 ) );
  OAI22_X1 u0_u1_u5_U7 (.B2( u0_u1_u5_n149 ) , .B1( u0_u1_u5_n150 ) , .A2( u0_u1_u5_n151 ) , .A1( u0_u1_u5_n152 ) , .ZN( u0_u1_u5_n165 ) );
  NAND2_X1 u0_u1_u5_U70 (.A2( u0_u1_u5_n103 ) , .A1( u0_u1_u5_n107 ) , .ZN( u0_u1_u5_n151 ) );
  NAND2_X1 u0_u1_u5_U71 (.A2( u0_u1_u5_n107 ) , .A1( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n120 ) );
  NAND2_X1 u0_u1_u5_U72 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n109 ) , .ZN( u0_u1_u5_n157 ) );
  AND2_X1 u0_u1_u5_U73 (.A2( u0_u1_u5_n100 ) , .A1( u0_u1_u5_n104 ) , .ZN( u0_u1_u5_n131 ) );
  INV_X1 u0_u1_u5_U74 (.A( u0_u1_u5_n102 ) , .ZN( u0_u1_u5_n195 ) );
  OAI221_X1 u0_u1_u5_U75 (.A( u0_u1_u5_n101 ) , .ZN( u0_u1_u5_n102 ) , .C2( u0_u1_u5_n115 ) , .C1( u0_u1_u5_n126 ) , .B1( u0_u1_u5_n134 ) , .B2( u0_u1_u5_n160 ) );
  OAI21_X1 u0_u1_u5_U76 (.ZN( u0_u1_u5_n101 ) , .B1( u0_u1_u5_n137 ) , .A( u0_u1_u5_n146 ) , .B2( u0_u1_u5_n147 ) );
  NOR2_X1 u0_u1_u5_U77 (.A2( u0_u1_X_34 ) , .A1( u0_u1_X_35 ) , .ZN( u0_u1_u5_n145 ) );
  NOR2_X1 u0_u1_u5_U78 (.A2( u0_u1_X_34 ) , .ZN( u0_u1_u5_n146 ) , .A1( u0_u1_u5_n171 ) );
  NOR2_X1 u0_u1_u5_U79 (.A2( u0_u1_X_31 ) , .A1( u0_u1_X_32 ) , .ZN( u0_u1_u5_n103 ) );
  NOR3_X1 u0_u1_u5_U8 (.A2( u0_u1_u5_n147 ) , .A1( u0_u1_u5_n148 ) , .ZN( u0_u1_u5_n149 ) , .A3( u0_u1_u5_n194 ) );
  NOR2_X1 u0_u1_u5_U80 (.A2( u0_u1_X_36 ) , .ZN( u0_u1_u5_n105 ) , .A1( u0_u1_u5_n180 ) );
  NOR2_X1 u0_u1_u5_U81 (.A2( u0_u1_X_33 ) , .ZN( u0_u1_u5_n108 ) , .A1( u0_u1_u5_n170 ) );
  NOR2_X1 u0_u1_u5_U82 (.A2( u0_u1_X_33 ) , .A1( u0_u1_X_36 ) , .ZN( u0_u1_u5_n107 ) );
  NOR2_X1 u0_u1_u5_U83 (.A2( u0_u1_X_31 ) , .ZN( u0_u1_u5_n104 ) , .A1( u0_u1_u5_n181 ) );
  NAND2_X1 u0_u1_u5_U84 (.A2( u0_u1_X_34 ) , .A1( u0_u1_X_35 ) , .ZN( u0_u1_u5_n153 ) );
  NAND2_X1 u0_u1_u5_U85 (.A1( u0_u1_X_34 ) , .ZN( u0_u1_u5_n126 ) , .A2( u0_u1_u5_n171 ) );
  AND2_X1 u0_u1_u5_U86 (.A1( u0_u1_X_31 ) , .A2( u0_u1_X_32 ) , .ZN( u0_u1_u5_n106 ) );
  AND2_X1 u0_u1_u5_U87 (.A1( u0_u1_X_31 ) , .ZN( u0_u1_u5_n109 ) , .A2( u0_u1_u5_n181 ) );
  INV_X1 u0_u1_u5_U88 (.A( u0_u1_X_33 ) , .ZN( u0_u1_u5_n180 ) );
  INV_X1 u0_u1_u5_U89 (.A( u0_u1_X_35 ) , .ZN( u0_u1_u5_n171 ) );
  NOR2_X1 u0_u1_u5_U9 (.ZN( u0_u1_u5_n135 ) , .A1( u0_u1_u5_n173 ) , .A2( u0_u1_u5_n176 ) );
  INV_X1 u0_u1_u5_U90 (.A( u0_u1_X_36 ) , .ZN( u0_u1_u5_n170 ) );
  INV_X1 u0_u1_u5_U91 (.A( u0_u1_X_32 ) , .ZN( u0_u1_u5_n181 ) );
  NAND4_X1 u0_u1_u5_U92 (.ZN( u0_out1_29 ) , .A4( u0_u1_u5_n129 ) , .A3( u0_u1_u5_n130 ) , .A2( u0_u1_u5_n168 ) , .A1( u0_u1_u5_n196 ) );
  AOI221_X1 u0_u1_u5_U93 (.A( u0_u1_u5_n128 ) , .ZN( u0_u1_u5_n129 ) , .C2( u0_u1_u5_n132 ) , .B2( u0_u1_u5_n159 ) , .B1( u0_u1_u5_n176 ) , .C1( u0_u1_u5_n184 ) );
  AOI222_X1 u0_u1_u5_U94 (.ZN( u0_u1_u5_n130 ) , .A2( u0_u1_u5_n146 ) , .B1( u0_u1_u5_n147 ) , .C2( u0_u1_u5_n175 ) , .B2( u0_u1_u5_n179 ) , .A1( u0_u1_u5_n188 ) , .C1( u0_u1_u5_n194 ) );
  NAND4_X1 u0_u1_u5_U95 (.ZN( u0_out1_19 ) , .A4( u0_u1_u5_n166 ) , .A3( u0_u1_u5_n167 ) , .A2( u0_u1_u5_n168 ) , .A1( u0_u1_u5_n169 ) );
  AOI22_X1 u0_u1_u5_U96 (.B2( u0_u1_u5_n145 ) , .A2( u0_u1_u5_n146 ) , .ZN( u0_u1_u5_n167 ) , .B1( u0_u1_u5_n182 ) , .A1( u0_u1_u5_n189 ) );
  NOR4_X1 u0_u1_u5_U97 (.A4( u0_u1_u5_n162 ) , .A3( u0_u1_u5_n163 ) , .A2( u0_u1_u5_n164 ) , .A1( u0_u1_u5_n165 ) , .ZN( u0_u1_u5_n166 ) );
  NAND4_X1 u0_u1_u5_U98 (.ZN( u0_out1_11 ) , .A4( u0_u1_u5_n143 ) , .A3( u0_u1_u5_n144 ) , .A2( u0_u1_u5_n169 ) , .A1( u0_u1_u5_n196 ) );
  AOI22_X1 u0_u1_u5_U99 (.A2( u0_u1_u5_n132 ) , .ZN( u0_u1_u5_n144 ) , .B2( u0_u1_u5_n145 ) , .B1( u0_u1_u5_n184 ) , .A1( u0_u1_u5_n194 ) );
  AOI22_X1 u0_u1_u6_U10 (.A2( u0_u1_u6_n151 ) , .B2( u0_u1_u6_n161 ) , .A1( u0_u1_u6_n167 ) , .B1( u0_u1_u6_n170 ) , .ZN( u0_u1_u6_n89 ) );
  AOI21_X1 u0_u1_u6_U11 (.B1( u0_u1_u6_n107 ) , .B2( u0_u1_u6_n132 ) , .A( u0_u1_u6_n158 ) , .ZN( u0_u1_u6_n88 ) );
  AOI21_X1 u0_u1_u6_U12 (.B2( u0_u1_u6_n147 ) , .B1( u0_u1_u6_n148 ) , .ZN( u0_u1_u6_n149 ) , .A( u0_u1_u6_n158 ) );
  AOI21_X1 u0_u1_u6_U13 (.ZN( u0_u1_u6_n106 ) , .A( u0_u1_u6_n142 ) , .B2( u0_u1_u6_n159 ) , .B1( u0_u1_u6_n164 ) );
  INV_X1 u0_u1_u6_U14 (.A( u0_u1_u6_n155 ) , .ZN( u0_u1_u6_n161 ) );
  INV_X1 u0_u1_u6_U15 (.A( u0_u1_u6_n128 ) , .ZN( u0_u1_u6_n164 ) );
  NAND2_X1 u0_u1_u6_U16 (.ZN( u0_u1_u6_n110 ) , .A1( u0_u1_u6_n122 ) , .A2( u0_u1_u6_n129 ) );
  NAND2_X1 u0_u1_u6_U17 (.ZN( u0_u1_u6_n124 ) , .A2( u0_u1_u6_n146 ) , .A1( u0_u1_u6_n148 ) );
  INV_X1 u0_u1_u6_U18 (.A( u0_u1_u6_n132 ) , .ZN( u0_u1_u6_n171 ) );
  AND2_X1 u0_u1_u6_U19 (.A1( u0_u1_u6_n100 ) , .ZN( u0_u1_u6_n130 ) , .A2( u0_u1_u6_n147 ) );
  INV_X1 u0_u1_u6_U20 (.A( u0_u1_u6_n127 ) , .ZN( u0_u1_u6_n173 ) );
  INV_X1 u0_u1_u6_U21 (.A( u0_u1_u6_n121 ) , .ZN( u0_u1_u6_n167 ) );
  INV_X1 u0_u1_u6_U22 (.A( u0_u1_u6_n100 ) , .ZN( u0_u1_u6_n169 ) );
  INV_X1 u0_u1_u6_U23 (.A( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n170 ) );
  INV_X1 u0_u1_u6_U24 (.A( u0_u1_u6_n113 ) , .ZN( u0_u1_u6_n168 ) );
  AND2_X1 u0_u1_u6_U25 (.A1( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n119 ) , .ZN( u0_u1_u6_n133 ) );
  AND2_X1 u0_u1_u6_U26 (.A2( u0_u1_u6_n121 ) , .A1( u0_u1_u6_n122 ) , .ZN( u0_u1_u6_n131 ) );
  AND3_X1 u0_u1_u6_U27 (.ZN( u0_u1_u6_n120 ) , .A2( u0_u1_u6_n127 ) , .A1( u0_u1_u6_n132 ) , .A3( u0_u1_u6_n145 ) );
  INV_X1 u0_u1_u6_U28 (.A( u0_u1_u6_n146 ) , .ZN( u0_u1_u6_n163 ) );
  AOI222_X1 u0_u1_u6_U29 (.ZN( u0_u1_u6_n114 ) , .A1( u0_u1_u6_n118 ) , .A2( u0_u1_u6_n126 ) , .B2( u0_u1_u6_n151 ) , .C2( u0_u1_u6_n159 ) , .C1( u0_u1_u6_n168 ) , .B1( u0_u1_u6_n169 ) );
  INV_X1 u0_u1_u6_U3 (.A( u0_u1_u6_n110 ) , .ZN( u0_u1_u6_n166 ) );
  NOR2_X1 u0_u1_u6_U30 (.A1( u0_u1_u6_n162 ) , .A2( u0_u1_u6_n165 ) , .ZN( u0_u1_u6_n98 ) );
  AOI211_X1 u0_u1_u6_U31 (.B( u0_u1_u6_n134 ) , .A( u0_u1_u6_n135 ) , .C1( u0_u1_u6_n136 ) , .ZN( u0_u1_u6_n137 ) , .C2( u0_u1_u6_n151 ) );
  AOI21_X1 u0_u1_u6_U32 (.B1( u0_u1_u6_n131 ) , .ZN( u0_u1_u6_n135 ) , .A( u0_u1_u6_n144 ) , .B2( u0_u1_u6_n146 ) );
  NAND4_X1 u0_u1_u6_U33 (.A4( u0_u1_u6_n127 ) , .A3( u0_u1_u6_n128 ) , .A2( u0_u1_u6_n129 ) , .A1( u0_u1_u6_n130 ) , .ZN( u0_u1_u6_n136 ) );
  AOI21_X1 u0_u1_u6_U34 (.B2( u0_u1_u6_n132 ) , .B1( u0_u1_u6_n133 ) , .ZN( u0_u1_u6_n134 ) , .A( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U35 (.A1( u0_u1_u6_n144 ) , .ZN( u0_u1_u6_n151 ) , .A2( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U36 (.ZN( u0_u1_u6_n132 ) , .A1( u0_u1_u6_n91 ) , .A2( u0_u1_u6_n97 ) );
  AOI22_X1 u0_u1_u6_U37 (.B2( u0_u1_u6_n110 ) , .B1( u0_u1_u6_n111 ) , .A1( u0_u1_u6_n112 ) , .ZN( u0_u1_u6_n115 ) , .A2( u0_u1_u6_n161 ) );
  NAND4_X1 u0_u1_u6_U38 (.A3( u0_u1_u6_n109 ) , .ZN( u0_u1_u6_n112 ) , .A4( u0_u1_u6_n132 ) , .A2( u0_u1_u6_n147 ) , .A1( u0_u1_u6_n166 ) );
  NOR2_X1 u0_u1_u6_U39 (.ZN( u0_u1_u6_n109 ) , .A1( u0_u1_u6_n170 ) , .A2( u0_u1_u6_n173 ) );
  INV_X1 u0_u1_u6_U4 (.A( u0_u1_u6_n142 ) , .ZN( u0_u1_u6_n174 ) );
  NOR2_X1 u0_u1_u6_U40 (.A2( u0_u1_u6_n126 ) , .ZN( u0_u1_u6_n155 ) , .A1( u0_u1_u6_n160 ) );
  NAND2_X1 u0_u1_u6_U41 (.ZN( u0_u1_u6_n146 ) , .A2( u0_u1_u6_n94 ) , .A1( u0_u1_u6_n99 ) );
  AOI21_X1 u0_u1_u6_U42 (.A( u0_u1_u6_n144 ) , .B2( u0_u1_u6_n145 ) , .B1( u0_u1_u6_n146 ) , .ZN( u0_u1_u6_n150 ) );
  INV_X1 u0_u1_u6_U43 (.A( u0_u1_u6_n111 ) , .ZN( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U44 (.ZN( u0_u1_u6_n127 ) , .A1( u0_u1_u6_n91 ) , .A2( u0_u1_u6_n92 ) );
  NAND2_X1 u0_u1_u6_U45 (.ZN( u0_u1_u6_n129 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n96 ) );
  INV_X1 u0_u1_u6_U46 (.A( u0_u1_u6_n144 ) , .ZN( u0_u1_u6_n159 ) );
  NAND2_X1 u0_u1_u6_U47 (.ZN( u0_u1_u6_n145 ) , .A2( u0_u1_u6_n97 ) , .A1( u0_u1_u6_n98 ) );
  NAND2_X1 u0_u1_u6_U48 (.ZN( u0_u1_u6_n148 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n94 ) );
  NAND2_X1 u0_u1_u6_U49 (.ZN( u0_u1_u6_n108 ) , .A2( u0_u1_u6_n139 ) , .A1( u0_u1_u6_n144 ) );
  NAND2_X1 u0_u1_u6_U5 (.A2( u0_u1_u6_n143 ) , .ZN( u0_u1_u6_n152 ) , .A1( u0_u1_u6_n166 ) );
  NAND2_X1 u0_u1_u6_U50 (.ZN( u0_u1_u6_n121 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n97 ) );
  NAND2_X1 u0_u1_u6_U51 (.ZN( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n95 ) );
  AND2_X1 u0_u1_u6_U52 (.ZN( u0_u1_u6_n118 ) , .A2( u0_u1_u6_n91 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U53 (.ZN( u0_u1_u6_n147 ) , .A2( u0_u1_u6_n98 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U54 (.ZN( u0_u1_u6_n128 ) , .A1( u0_u1_u6_n94 ) , .A2( u0_u1_u6_n96 ) );
  NAND2_X1 u0_u1_u6_U55 (.ZN( u0_u1_u6_n119 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U56 (.ZN( u0_u1_u6_n123 ) , .A2( u0_u1_u6_n91 ) , .A1( u0_u1_u6_n96 ) );
  NAND2_X1 u0_u1_u6_U57 (.ZN( u0_u1_u6_n100 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n98 ) );
  NAND2_X1 u0_u1_u6_U58 (.ZN( u0_u1_u6_n122 ) , .A1( u0_u1_u6_n94 ) , .A2( u0_u1_u6_n97 ) );
  INV_X1 u0_u1_u6_U59 (.A( u0_u1_u6_n139 ) , .ZN( u0_u1_u6_n160 ) );
  AOI22_X1 u0_u1_u6_U6 (.B2( u0_u1_u6_n101 ) , .A1( u0_u1_u6_n102 ) , .ZN( u0_u1_u6_n103 ) , .B1( u0_u1_u6_n160 ) , .A2( u0_u1_u6_n161 ) );
  NAND2_X1 u0_u1_u6_U60 (.ZN( u0_u1_u6_n113 ) , .A1( u0_u1_u6_n96 ) , .A2( u0_u1_u6_n98 ) );
  NOR2_X1 u0_u1_u6_U61 (.A2( u0_u1_X_40 ) , .A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n126 ) );
  NOR2_X1 u0_u1_u6_U62 (.A2( u0_u1_X_39 ) , .A1( u0_u1_X_42 ) , .ZN( u0_u1_u6_n92 ) );
  NOR2_X1 u0_u1_u6_U63 (.A2( u0_u1_X_39 ) , .A1( u0_u1_u6_n156 ) , .ZN( u0_u1_u6_n97 ) );
  NOR2_X1 u0_u1_u6_U64 (.A2( u0_u1_X_38 ) , .A1( u0_u1_u6_n165 ) , .ZN( u0_u1_u6_n95 ) );
  NOR2_X1 u0_u1_u6_U65 (.A2( u0_u1_X_41 ) , .ZN( u0_u1_u6_n111 ) , .A1( u0_u1_u6_n157 ) );
  NOR2_X1 u0_u1_u6_U66 (.A2( u0_u1_X_37 ) , .A1( u0_u1_u6_n162 ) , .ZN( u0_u1_u6_n94 ) );
  NOR2_X1 u0_u1_u6_U67 (.A2( u0_u1_X_37 ) , .A1( u0_u1_X_38 ) , .ZN( u0_u1_u6_n91 ) );
  NAND2_X1 u0_u1_u6_U68 (.A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n144 ) , .A2( u0_u1_u6_n157 ) );
  NAND2_X1 u0_u1_u6_U69 (.A2( u0_u1_X_40 ) , .A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n139 ) );
  NOR2_X1 u0_u1_u6_U7 (.A1( u0_u1_u6_n118 ) , .ZN( u0_u1_u6_n143 ) , .A2( u0_u1_u6_n168 ) );
  AND2_X1 u0_u1_u6_U70 (.A1( u0_u1_X_39 ) , .A2( u0_u1_u6_n156 ) , .ZN( u0_u1_u6_n96 ) );
  AND2_X1 u0_u1_u6_U71 (.A1( u0_u1_X_39 ) , .A2( u0_u1_X_42 ) , .ZN( u0_u1_u6_n99 ) );
  INV_X1 u0_u1_u6_U72 (.A( u0_u1_X_40 ) , .ZN( u0_u1_u6_n157 ) );
  INV_X1 u0_u1_u6_U73 (.A( u0_u1_X_37 ) , .ZN( u0_u1_u6_n165 ) );
  INV_X1 u0_u1_u6_U74 (.A( u0_u1_X_38 ) , .ZN( u0_u1_u6_n162 ) );
  INV_X1 u0_u1_u6_U75 (.A( u0_u1_X_42 ) , .ZN( u0_u1_u6_n156 ) );
  NAND4_X1 u0_u1_u6_U76 (.ZN( u0_out1_12 ) , .A4( u0_u1_u6_n114 ) , .A3( u0_u1_u6_n115 ) , .A2( u0_u1_u6_n116 ) , .A1( u0_u1_u6_n117 ) );
  OAI22_X1 u0_u1_u6_U77 (.B2( u0_u1_u6_n111 ) , .ZN( u0_u1_u6_n116 ) , .B1( u0_u1_u6_n126 ) , .A2( u0_u1_u6_n164 ) , .A1( u0_u1_u6_n167 ) );
  OAI21_X1 u0_u1_u6_U78 (.A( u0_u1_u6_n108 ) , .ZN( u0_u1_u6_n117 ) , .B2( u0_u1_u6_n141 ) , .B1( u0_u1_u6_n163 ) );
  NAND4_X1 u0_u1_u6_U79 (.ZN( u0_out1_32 ) , .A4( u0_u1_u6_n103 ) , .A3( u0_u1_u6_n104 ) , .A2( u0_u1_u6_n105 ) , .A1( u0_u1_u6_n106 ) );
  OAI21_X1 u0_u1_u6_U8 (.A( u0_u1_u6_n159 ) , .B1( u0_u1_u6_n169 ) , .B2( u0_u1_u6_n173 ) , .ZN( u0_u1_u6_n90 ) );
  AOI22_X1 u0_u1_u6_U80 (.ZN( u0_u1_u6_n105 ) , .A2( u0_u1_u6_n108 ) , .A1( u0_u1_u6_n118 ) , .B2( u0_u1_u6_n126 ) , .B1( u0_u1_u6_n171 ) );
  AOI22_X1 u0_u1_u6_U81 (.ZN( u0_u1_u6_n104 ) , .A1( u0_u1_u6_n111 ) , .B1( u0_u1_u6_n124 ) , .B2( u0_u1_u6_n151 ) , .A2( u0_u1_u6_n93 ) );
  OAI211_X1 u0_u1_u6_U82 (.ZN( u0_out1_22 ) , .B( u0_u1_u6_n137 ) , .A( u0_u1_u6_n138 ) , .C2( u0_u1_u6_n139 ) , .C1( u0_u1_u6_n140 ) );
  AND4_X1 u0_u1_u6_U83 (.A3( u0_u1_u6_n119 ) , .A1( u0_u1_u6_n120 ) , .A4( u0_u1_u6_n129 ) , .ZN( u0_u1_u6_n140 ) , .A2( u0_u1_u6_n143 ) );
  AOI22_X1 u0_u1_u6_U84 (.B1( u0_u1_u6_n124 ) , .A2( u0_u1_u6_n125 ) , .A1( u0_u1_u6_n126 ) , .ZN( u0_u1_u6_n138 ) , .B2( u0_u1_u6_n161 ) );
  OAI211_X1 u0_u1_u6_U85 (.ZN( u0_out1_7 ) , .B( u0_u1_u6_n153 ) , .C2( u0_u1_u6_n154 ) , .C1( u0_u1_u6_n155 ) , .A( u0_u1_u6_n174 ) );
  NOR3_X1 u0_u1_u6_U86 (.A1( u0_u1_u6_n141 ) , .ZN( u0_u1_u6_n154 ) , .A3( u0_u1_u6_n164 ) , .A2( u0_u1_u6_n171 ) );
  AOI211_X1 u0_u1_u6_U87 (.B( u0_u1_u6_n149 ) , .A( u0_u1_u6_n150 ) , .C2( u0_u1_u6_n151 ) , .C1( u0_u1_u6_n152 ) , .ZN( u0_u1_u6_n153 ) );
  NAND3_X1 u0_u1_u6_U88 (.A2( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n125 ) , .A1( u0_u1_u6_n130 ) , .A3( u0_u1_u6_n131 ) );
  NAND3_X1 u0_u1_u6_U89 (.A3( u0_u1_u6_n133 ) , .ZN( u0_u1_u6_n141 ) , .A1( u0_u1_u6_n145 ) , .A2( u0_u1_u6_n148 ) );
  INV_X1 u0_u1_u6_U9 (.ZN( u0_u1_u6_n172 ) , .A( u0_u1_u6_n88 ) );
  NAND3_X1 u0_u1_u6_U90 (.ZN( u0_u1_u6_n101 ) , .A3( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n121 ) , .A1( u0_u1_u6_n127 ) );
  NAND3_X1 u0_u1_u6_U91 (.ZN( u0_u1_u6_n102 ) , .A3( u0_u1_u6_n130 ) , .A2( u0_u1_u6_n145 ) , .A1( u0_u1_u6_n166 ) );
  NAND3_X1 u0_u1_u6_U92 (.A3( u0_u1_u6_n113 ) , .A1( u0_u1_u6_n119 ) , .A2( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n93 ) );
  NAND3_X1 u0_u1_u6_U93 (.ZN( u0_u1_u6_n142 ) , .A2( u0_u1_u6_n172 ) , .A3( u0_u1_u6_n89 ) , .A1( u0_u1_u6_n90 ) );
  XOR2_X1 u0_u2_U1 (.B( u0_K3_9 ) , .A( u0_R1_6 ) , .Z( u0_u2_X_9 ) );
  XOR2_X1 u0_u2_U16 (.B( u0_K3_3 ) , .A( u0_R1_2 ) , .Z( u0_u2_X_3 ) );
  XOR2_X1 u0_u2_U2 (.B( u0_K3_8 ) , .A( u0_R1_5 ) , .Z( u0_u2_X_8 ) );
  XOR2_X1 u0_u2_U27 (.B( u0_K3_2 ) , .A( u0_R1_1 ) , .Z( u0_u2_X_2 ) );
  XOR2_X1 u0_u2_U3 (.B( u0_K3_7 ) , .A( u0_R1_4 ) , .Z( u0_u2_X_7 ) );
  XOR2_X1 u0_u2_U33 (.B( u0_K3_24 ) , .A( u0_R1_17 ) , .Z( u0_u2_X_24 ) );
  XOR2_X1 u0_u2_U34 (.B( u0_K3_23 ) , .A( u0_R1_16 ) , .Z( u0_u2_X_23 ) );
  XOR2_X1 u0_u2_U35 (.B( u0_K3_22 ) , .A( u0_R1_15 ) , .Z( u0_u2_X_22 ) );
  XOR2_X1 u0_u2_U36 (.B( u0_K3_21 ) , .A( u0_R1_14 ) , .Z( u0_u2_X_21 ) );
  XOR2_X1 u0_u2_U37 (.B( u0_K3_20 ) , .A( u0_R1_13 ) , .Z( u0_u2_X_20 ) );
  XOR2_X1 u0_u2_U38 (.B( u0_K3_1 ) , .A( u0_R1_32 ) , .Z( u0_u2_X_1 ) );
  XOR2_X1 u0_u2_U39 (.B( u0_K3_19 ) , .A( u0_R1_12 ) , .Z( u0_u2_X_19 ) );
  XOR2_X1 u0_u2_U4 (.B( u0_K3_6 ) , .A( u0_R1_5 ) , .Z( u0_u2_X_6 ) );
  XOR2_X1 u0_u2_U40 (.B( u0_K3_18 ) , .A( u0_R1_13 ) , .Z( u0_u2_X_18 ) );
  XOR2_X1 u0_u2_U41 (.B( u0_K3_17 ) , .A( u0_R1_12 ) , .Z( u0_u2_X_17 ) );
  XOR2_X1 u0_u2_U42 (.B( u0_K3_16 ) , .A( u0_R1_11 ) , .Z( u0_u2_X_16 ) );
  XOR2_X1 u0_u2_U43 (.B( u0_K3_15 ) , .A( u0_R1_10 ) , .Z( u0_u2_X_15 ) );
  XOR2_X1 u0_u2_U44 (.B( u0_K3_14 ) , .A( u0_R1_9 ) , .Z( u0_u2_X_14 ) );
  XOR2_X1 u0_u2_U45 (.B( u0_K3_13 ) , .A( u0_R1_8 ) , .Z( u0_u2_X_13 ) );
  XOR2_X1 u0_u2_U46 (.B( u0_K3_12 ) , .A( u0_R1_9 ) , .Z( u0_u2_X_12 ) );
  XOR2_X1 u0_u2_U47 (.B( u0_K3_11 ) , .A( u0_R1_8 ) , .Z( u0_u2_X_11 ) );
  XOR2_X1 u0_u2_U48 (.B( u0_K3_10 ) , .A( u0_R1_7 ) , .Z( u0_u2_X_10 ) );
  XOR2_X1 u0_u2_U5 (.B( u0_K3_5 ) , .A( u0_R1_4 ) , .Z( u0_u2_X_5 ) );
  XOR2_X1 u0_u2_U6 (.B( u0_K3_4 ) , .A( u0_R1_3 ) , .Z( u0_u2_X_4 ) );
  AND3_X1 u0_u2_u0_U10 (.A2( u0_u2_u0_n112 ) , .ZN( u0_u2_u0_n127 ) , .A3( u0_u2_u0_n130 ) , .A1( u0_u2_u0_n148 ) );
  NAND2_X1 u0_u2_u0_U11 (.ZN( u0_u2_u0_n113 ) , .A1( u0_u2_u0_n139 ) , .A2( u0_u2_u0_n149 ) );
  AND2_X1 u0_u2_u0_U12 (.ZN( u0_u2_u0_n107 ) , .A1( u0_u2_u0_n130 ) , .A2( u0_u2_u0_n140 ) );
  AND2_X1 u0_u2_u0_U13 (.A2( u0_u2_u0_n129 ) , .A1( u0_u2_u0_n130 ) , .ZN( u0_u2_u0_n151 ) );
  AND2_X1 u0_u2_u0_U14 (.A1( u0_u2_u0_n108 ) , .A2( u0_u2_u0_n125 ) , .ZN( u0_u2_u0_n145 ) );
  INV_X1 u0_u2_u0_U15 (.A( u0_u2_u0_n143 ) , .ZN( u0_u2_u0_n173 ) );
  NOR2_X1 u0_u2_u0_U16 (.A2( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n147 ) , .A1( u0_u2_u0_n160 ) );
  INV_X1 u0_u2_u0_U17 (.ZN( u0_u2_u0_n172 ) , .A( u0_u2_u0_n88 ) );
  OAI222_X1 u0_u2_u0_U18 (.C1( u0_u2_u0_n108 ) , .A1( u0_u2_u0_n125 ) , .B2( u0_u2_u0_n128 ) , .B1( u0_u2_u0_n144 ) , .A2( u0_u2_u0_n158 ) , .C2( u0_u2_u0_n161 ) , .ZN( u0_u2_u0_n88 ) );
  NOR2_X1 u0_u2_u0_U19 (.A1( u0_u2_u0_n163 ) , .A2( u0_u2_u0_n164 ) , .ZN( u0_u2_u0_n95 ) );
  AOI21_X1 u0_u2_u0_U20 (.B1( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n132 ) , .A( u0_u2_u0_n165 ) , .B2( u0_u2_u0_n93 ) );
  INV_X1 u0_u2_u0_U21 (.A( u0_u2_u0_n142 ) , .ZN( u0_u2_u0_n165 ) );
  OAI221_X1 u0_u2_u0_U22 (.C1( u0_u2_u0_n121 ) , .ZN( u0_u2_u0_n122 ) , .B2( u0_u2_u0_n127 ) , .A( u0_u2_u0_n143 ) , .B1( u0_u2_u0_n144 ) , .C2( u0_u2_u0_n147 ) );
  OAI22_X1 u0_u2_u0_U23 (.B1( u0_u2_u0_n125 ) , .ZN( u0_u2_u0_n126 ) , .A1( u0_u2_u0_n138 ) , .A2( u0_u2_u0_n146 ) , .B2( u0_u2_u0_n147 ) );
  OAI22_X1 u0_u2_u0_U24 (.B1( u0_u2_u0_n131 ) , .A1( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n147 ) , .A2( u0_u2_u0_n90 ) , .ZN( u0_u2_u0_n91 ) );
  AND3_X1 u0_u2_u0_U25 (.A3( u0_u2_u0_n121 ) , .A2( u0_u2_u0_n125 ) , .A1( u0_u2_u0_n148 ) , .ZN( u0_u2_u0_n90 ) );
  INV_X1 u0_u2_u0_U26 (.A( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n161 ) );
  NOR2_X1 u0_u2_u0_U27 (.A1( u0_u2_u0_n120 ) , .ZN( u0_u2_u0_n143 ) , .A2( u0_u2_u0_n167 ) );
  OAI221_X1 u0_u2_u0_U28 (.C1( u0_u2_u0_n112 ) , .ZN( u0_u2_u0_n120 ) , .B1( u0_u2_u0_n138 ) , .B2( u0_u2_u0_n141 ) , .C2( u0_u2_u0_n147 ) , .A( u0_u2_u0_n172 ) );
  AOI211_X1 u0_u2_u0_U29 (.B( u0_u2_u0_n115 ) , .A( u0_u2_u0_n116 ) , .C2( u0_u2_u0_n117 ) , .C1( u0_u2_u0_n118 ) , .ZN( u0_u2_u0_n119 ) );
  INV_X1 u0_u2_u0_U3 (.A( u0_u2_u0_n113 ) , .ZN( u0_u2_u0_n166 ) );
  AOI22_X1 u0_u2_u0_U30 (.B2( u0_u2_u0_n109 ) , .A2( u0_u2_u0_n110 ) , .ZN( u0_u2_u0_n111 ) , .B1( u0_u2_u0_n118 ) , .A1( u0_u2_u0_n160 ) );
  INV_X1 u0_u2_u0_U31 (.A( u0_u2_u0_n118 ) , .ZN( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U32 (.ZN( u0_u2_u0_n104 ) , .B1( u0_u2_u0_n107 ) , .B2( u0_u2_u0_n141 ) , .A( u0_u2_u0_n144 ) );
  AOI21_X1 u0_u2_u0_U33 (.B1( u0_u2_u0_n127 ) , .B2( u0_u2_u0_n129 ) , .A( u0_u2_u0_n138 ) , .ZN( u0_u2_u0_n96 ) );
  AOI21_X1 u0_u2_u0_U34 (.ZN( u0_u2_u0_n116 ) , .B2( u0_u2_u0_n142 ) , .A( u0_u2_u0_n144 ) , .B1( u0_u2_u0_n166 ) );
  NAND2_X1 u0_u2_u0_U35 (.A1( u0_u2_u0_n100 ) , .A2( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n125 ) );
  NAND2_X1 u0_u2_u0_U36 (.A1( u0_u2_u0_n101 ) , .A2( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n150 ) );
  INV_X1 u0_u2_u0_U37 (.A( u0_u2_u0_n138 ) , .ZN( u0_u2_u0_n160 ) );
  NAND2_X1 u0_u2_u0_U38 (.A1( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n128 ) , .A2( u0_u2_u0_n95 ) );
  NAND2_X1 u0_u2_u0_U39 (.A1( u0_u2_u0_n100 ) , .ZN( u0_u2_u0_n129 ) , .A2( u0_u2_u0_n95 ) );
  AOI21_X1 u0_u2_u0_U4 (.B1( u0_u2_u0_n114 ) , .ZN( u0_u2_u0_n115 ) , .B2( u0_u2_u0_n129 ) , .A( u0_u2_u0_n161 ) );
  NAND2_X1 u0_u2_u0_U40 (.A2( u0_u2_u0_n100 ) , .ZN( u0_u2_u0_n131 ) , .A1( u0_u2_u0_n92 ) );
  NAND2_X1 u0_u2_u0_U41 (.A2( u0_u2_u0_n100 ) , .A1( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n139 ) );
  NAND2_X1 u0_u2_u0_U42 (.ZN( u0_u2_u0_n148 ) , .A1( u0_u2_u0_n93 ) , .A2( u0_u2_u0_n95 ) );
  NAND2_X1 u0_u2_u0_U43 (.A2( u0_u2_u0_n102 ) , .A1( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n149 ) );
  NAND2_X1 u0_u2_u0_U44 (.A2( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n114 ) , .A1( u0_u2_u0_n92 ) );
  NAND2_X1 u0_u2_u0_U45 (.A2( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n121 ) , .A1( u0_u2_u0_n93 ) );
  NAND2_X1 u0_u2_u0_U46 (.ZN( u0_u2_u0_n112 ) , .A2( u0_u2_u0_n92 ) , .A1( u0_u2_u0_n93 ) );
  OR3_X1 u0_u2_u0_U47 (.A3( u0_u2_u0_n152 ) , .A2( u0_u2_u0_n153 ) , .A1( u0_u2_u0_n154 ) , .ZN( u0_u2_u0_n155 ) );
  AOI21_X1 u0_u2_u0_U48 (.B2( u0_u2_u0_n150 ) , .B1( u0_u2_u0_n151 ) , .ZN( u0_u2_u0_n152 ) , .A( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U49 (.A( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n145 ) , .B1( u0_u2_u0_n146 ) , .ZN( u0_u2_u0_n154 ) );
  AOI21_X1 u0_u2_u0_U5 (.B2( u0_u2_u0_n131 ) , .ZN( u0_u2_u0_n134 ) , .B1( u0_u2_u0_n151 ) , .A( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U50 (.A( u0_u2_u0_n147 ) , .B2( u0_u2_u0_n148 ) , .B1( u0_u2_u0_n149 ) , .ZN( u0_u2_u0_n153 ) );
  INV_X1 u0_u2_u0_U51 (.ZN( u0_u2_u0_n171 ) , .A( u0_u2_u0_n99 ) );
  OAI211_X1 u0_u2_u0_U52 (.C2( u0_u2_u0_n140 ) , .C1( u0_u2_u0_n161 ) , .A( u0_u2_u0_n169 ) , .B( u0_u2_u0_n98 ) , .ZN( u0_u2_u0_n99 ) );
  AOI211_X1 u0_u2_u0_U53 (.C1( u0_u2_u0_n118 ) , .A( u0_u2_u0_n123 ) , .B( u0_u2_u0_n96 ) , .C2( u0_u2_u0_n97 ) , .ZN( u0_u2_u0_n98 ) );
  INV_X1 u0_u2_u0_U54 (.ZN( u0_u2_u0_n169 ) , .A( u0_u2_u0_n91 ) );
  NOR2_X1 u0_u2_u0_U55 (.A2( u0_u2_X_6 ) , .ZN( u0_u2_u0_n100 ) , .A1( u0_u2_u0_n162 ) );
  NOR2_X1 u0_u2_u0_U56 (.A2( u0_u2_X_4 ) , .A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n118 ) );
  NOR2_X1 u0_u2_u0_U57 (.A2( u0_u2_X_2 ) , .ZN( u0_u2_u0_n103 ) , .A1( u0_u2_u0_n164 ) );
  NOR2_X1 u0_u2_u0_U58 (.A2( u0_u2_X_1 ) , .A1( u0_u2_X_2 ) , .ZN( u0_u2_u0_n92 ) );
  NOR2_X1 u0_u2_u0_U59 (.A2( u0_u2_X_1 ) , .ZN( u0_u2_u0_n101 ) , .A1( u0_u2_u0_n163 ) );
  NOR2_X1 u0_u2_u0_U6 (.A1( u0_u2_u0_n108 ) , .ZN( u0_u2_u0_n123 ) , .A2( u0_u2_u0_n158 ) );
  NAND2_X1 u0_u2_u0_U60 (.A2( u0_u2_X_4 ) , .A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n144 ) );
  NOR2_X1 u0_u2_u0_U61 (.A2( u0_u2_X_5 ) , .ZN( u0_u2_u0_n136 ) , .A1( u0_u2_u0_n159 ) );
  NAND2_X1 u0_u2_u0_U62 (.A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n138 ) , .A2( u0_u2_u0_n159 ) );
  AND2_X1 u0_u2_u0_U63 (.A2( u0_u2_X_3 ) , .A1( u0_u2_X_6 ) , .ZN( u0_u2_u0_n102 ) );
  AND2_X1 u0_u2_u0_U64 (.A1( u0_u2_X_6 ) , .A2( u0_u2_u0_n162 ) , .ZN( u0_u2_u0_n93 ) );
  INV_X1 u0_u2_u0_U65 (.A( u0_u2_X_4 ) , .ZN( u0_u2_u0_n159 ) );
  INV_X1 u0_u2_u0_U66 (.A( u0_u2_X_1 ) , .ZN( u0_u2_u0_n164 ) );
  INV_X1 u0_u2_u0_U67 (.A( u0_u2_X_2 ) , .ZN( u0_u2_u0_n163 ) );
  INV_X1 u0_u2_u0_U68 (.ZN( u0_u2_u0_n174 ) , .A( u0_u2_u0_n89 ) );
  AOI211_X1 u0_u2_u0_U69 (.B( u0_u2_u0_n104 ) , .A( u0_u2_u0_n105 ) , .ZN( u0_u2_u0_n106 ) , .C2( u0_u2_u0_n113 ) , .C1( u0_u2_u0_n160 ) );
  OAI21_X1 u0_u2_u0_U7 (.B1( u0_u2_u0_n150 ) , .B2( u0_u2_u0_n158 ) , .A( u0_u2_u0_n172 ) , .ZN( u0_u2_u0_n89 ) );
  INV_X1 u0_u2_u0_U70 (.A( u0_u2_u0_n126 ) , .ZN( u0_u2_u0_n168 ) );
  AOI211_X1 u0_u2_u0_U71 (.B( u0_u2_u0_n133 ) , .A( u0_u2_u0_n134 ) , .C2( u0_u2_u0_n135 ) , .C1( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n137 ) );
  OR4_X1 u0_u2_u0_U72 (.ZN( u0_out2_31 ) , .A4( u0_u2_u0_n155 ) , .A2( u0_u2_u0_n156 ) , .A1( u0_u2_u0_n157 ) , .A3( u0_u2_u0_n173 ) );
  AOI21_X1 u0_u2_u0_U73 (.A( u0_u2_u0_n138 ) , .B2( u0_u2_u0_n139 ) , .B1( u0_u2_u0_n140 ) , .ZN( u0_u2_u0_n157 ) );
  AOI21_X1 u0_u2_u0_U74 (.B2( u0_u2_u0_n141 ) , .B1( u0_u2_u0_n142 ) , .ZN( u0_u2_u0_n156 ) , .A( u0_u2_u0_n161 ) );
  OR4_X1 u0_u2_u0_U75 (.ZN( u0_out2_17 ) , .A4( u0_u2_u0_n122 ) , .A2( u0_u2_u0_n123 ) , .A1( u0_u2_u0_n124 ) , .A3( u0_u2_u0_n170 ) );
  AOI21_X1 u0_u2_u0_U76 (.B2( u0_u2_u0_n107 ) , .ZN( u0_u2_u0_n124 ) , .B1( u0_u2_u0_n128 ) , .A( u0_u2_u0_n161 ) );
  INV_X1 u0_u2_u0_U77 (.A( u0_u2_u0_n111 ) , .ZN( u0_u2_u0_n170 ) );
  AOI21_X1 u0_u2_u0_U78 (.B1( u0_u2_u0_n132 ) , .ZN( u0_u2_u0_n133 ) , .A( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n166 ) );
  OAI22_X1 u0_u2_u0_U79 (.ZN( u0_u2_u0_n105 ) , .A2( u0_u2_u0_n132 ) , .B1( u0_u2_u0_n146 ) , .A1( u0_u2_u0_n147 ) , .B2( u0_u2_u0_n161 ) );
  AND2_X1 u0_u2_u0_U8 (.A1( u0_u2_u0_n114 ) , .A2( u0_u2_u0_n121 ) , .ZN( u0_u2_u0_n146 ) );
  NAND2_X1 u0_u2_u0_U80 (.ZN( u0_u2_u0_n110 ) , .A2( u0_u2_u0_n132 ) , .A1( u0_u2_u0_n145 ) );
  INV_X1 u0_u2_u0_U81 (.A( u0_u2_u0_n119 ) , .ZN( u0_u2_u0_n167 ) );
  NAND2_X1 u0_u2_u0_U82 (.A2( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n140 ) , .A1( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U83 (.A1( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n130 ) , .A2( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U84 (.ZN( u0_u2_u0_n108 ) , .A1( u0_u2_u0_n92 ) , .A2( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U85 (.ZN( u0_u2_u0_n142 ) , .A1( u0_u2_u0_n94 ) , .A2( u0_u2_u0_n95 ) );
  INV_X1 u0_u2_u0_U86 (.A( u0_u2_X_3 ) , .ZN( u0_u2_u0_n162 ) );
  NOR2_X1 u0_u2_u0_U87 (.A2( u0_u2_X_3 ) , .A1( u0_u2_X_6 ) , .ZN( u0_u2_u0_n94 ) );
  NAND3_X1 u0_u2_u0_U88 (.ZN( u0_out2_23 ) , .A3( u0_u2_u0_n137 ) , .A1( u0_u2_u0_n168 ) , .A2( u0_u2_u0_n171 ) );
  NAND3_X1 u0_u2_u0_U89 (.A3( u0_u2_u0_n127 ) , .A2( u0_u2_u0_n128 ) , .ZN( u0_u2_u0_n135 ) , .A1( u0_u2_u0_n150 ) );
  AND2_X1 u0_u2_u0_U9 (.A1( u0_u2_u0_n131 ) , .ZN( u0_u2_u0_n141 ) , .A2( u0_u2_u0_n150 ) );
  NAND3_X1 u0_u2_u0_U90 (.ZN( u0_u2_u0_n117 ) , .A3( u0_u2_u0_n132 ) , .A2( u0_u2_u0_n139 ) , .A1( u0_u2_u0_n148 ) );
  NAND3_X1 u0_u2_u0_U91 (.ZN( u0_u2_u0_n109 ) , .A2( u0_u2_u0_n114 ) , .A3( u0_u2_u0_n140 ) , .A1( u0_u2_u0_n149 ) );
  NAND3_X1 u0_u2_u0_U92 (.ZN( u0_out2_9 ) , .A3( u0_u2_u0_n106 ) , .A2( u0_u2_u0_n171 ) , .A1( u0_u2_u0_n174 ) );
  NAND3_X1 u0_u2_u0_U93 (.A2( u0_u2_u0_n128 ) , .A1( u0_u2_u0_n132 ) , .A3( u0_u2_u0_n146 ) , .ZN( u0_u2_u0_n97 ) );
  NOR2_X1 u0_u2_u1_U10 (.A1( u0_u2_u1_n112 ) , .A2( u0_u2_u1_n116 ) , .ZN( u0_u2_u1_n118 ) );
  NAND3_X1 u0_u2_u1_U100 (.ZN( u0_u2_u1_n113 ) , .A1( u0_u2_u1_n120 ) , .A3( u0_u2_u1_n133 ) , .A2( u0_u2_u1_n155 ) );
  OAI21_X1 u0_u2_u1_U11 (.ZN( u0_u2_u1_n101 ) , .B1( u0_u2_u1_n141 ) , .A( u0_u2_u1_n146 ) , .B2( u0_u2_u1_n183 ) );
  AOI21_X1 u0_u2_u1_U12 (.B2( u0_u2_u1_n155 ) , .B1( u0_u2_u1_n156 ) , .ZN( u0_u2_u1_n157 ) , .A( u0_u2_u1_n174 ) );
  OR4_X1 u0_u2_u1_U13 (.A4( u0_u2_u1_n106 ) , .A3( u0_u2_u1_n107 ) , .ZN( u0_u2_u1_n108 ) , .A1( u0_u2_u1_n117 ) , .A2( u0_u2_u1_n184 ) );
  AOI21_X1 u0_u2_u1_U14 (.ZN( u0_u2_u1_n106 ) , .A( u0_u2_u1_n112 ) , .B1( u0_u2_u1_n154 ) , .B2( u0_u2_u1_n156 ) );
  INV_X1 u0_u2_u1_U15 (.A( u0_u2_u1_n101 ) , .ZN( u0_u2_u1_n184 ) );
  AOI21_X1 u0_u2_u1_U16 (.ZN( u0_u2_u1_n107 ) , .B1( u0_u2_u1_n134 ) , .B2( u0_u2_u1_n149 ) , .A( u0_u2_u1_n174 ) );
  NAND2_X1 u0_u2_u1_U17 (.ZN( u0_u2_u1_n140 ) , .A2( u0_u2_u1_n150 ) , .A1( u0_u2_u1_n155 ) );
  NAND2_X1 u0_u2_u1_U18 (.A1( u0_u2_u1_n131 ) , .ZN( u0_u2_u1_n147 ) , .A2( u0_u2_u1_n153 ) );
  INV_X1 u0_u2_u1_U19 (.A( u0_u2_u1_n139 ) , .ZN( u0_u2_u1_n174 ) );
  INV_X1 u0_u2_u1_U20 (.A( u0_u2_u1_n112 ) , .ZN( u0_u2_u1_n171 ) );
  NAND2_X1 u0_u2_u1_U21 (.ZN( u0_u2_u1_n141 ) , .A1( u0_u2_u1_n153 ) , .A2( u0_u2_u1_n156 ) );
  AND2_X1 u0_u2_u1_U22 (.A1( u0_u2_u1_n123 ) , .ZN( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n161 ) );
  NAND2_X1 u0_u2_u1_U23 (.A2( u0_u2_u1_n115 ) , .A1( u0_u2_u1_n116 ) , .ZN( u0_u2_u1_n148 ) );
  NAND2_X1 u0_u2_u1_U24 (.A2( u0_u2_u1_n133 ) , .A1( u0_u2_u1_n135 ) , .ZN( u0_u2_u1_n159 ) );
  NAND2_X1 u0_u2_u1_U25 (.A2( u0_u2_u1_n115 ) , .A1( u0_u2_u1_n120 ) , .ZN( u0_u2_u1_n132 ) );
  INV_X1 u0_u2_u1_U26 (.A( u0_u2_u1_n154 ) , .ZN( u0_u2_u1_n178 ) );
  INV_X1 u0_u2_u1_U27 (.A( u0_u2_u1_n151 ) , .ZN( u0_u2_u1_n183 ) );
  AND2_X1 u0_u2_u1_U28 (.A1( u0_u2_u1_n129 ) , .A2( u0_u2_u1_n133 ) , .ZN( u0_u2_u1_n149 ) );
  INV_X1 u0_u2_u1_U29 (.A( u0_u2_u1_n131 ) , .ZN( u0_u2_u1_n180 ) );
  INV_X1 u0_u2_u1_U3 (.A( u0_u2_u1_n159 ) , .ZN( u0_u2_u1_n182 ) );
  OAI221_X1 u0_u2_u1_U30 (.A( u0_u2_u1_n119 ) , .C2( u0_u2_u1_n129 ) , .ZN( u0_u2_u1_n138 ) , .B2( u0_u2_u1_n152 ) , .C1( u0_u2_u1_n174 ) , .B1( u0_u2_u1_n187 ) );
  INV_X1 u0_u2_u1_U31 (.A( u0_u2_u1_n148 ) , .ZN( u0_u2_u1_n187 ) );
  AOI211_X1 u0_u2_u1_U32 (.B( u0_u2_u1_n117 ) , .A( u0_u2_u1_n118 ) , .ZN( u0_u2_u1_n119 ) , .C2( u0_u2_u1_n146 ) , .C1( u0_u2_u1_n159 ) );
  NOR2_X1 u0_u2_u1_U33 (.A1( u0_u2_u1_n168 ) , .A2( u0_u2_u1_n176 ) , .ZN( u0_u2_u1_n98 ) );
  AOI211_X1 u0_u2_u1_U34 (.B( u0_u2_u1_n162 ) , .A( u0_u2_u1_n163 ) , .C2( u0_u2_u1_n164 ) , .ZN( u0_u2_u1_n165 ) , .C1( u0_u2_u1_n171 ) );
  AOI21_X1 u0_u2_u1_U35 (.A( u0_u2_u1_n160 ) , .B2( u0_u2_u1_n161 ) , .ZN( u0_u2_u1_n162 ) , .B1( u0_u2_u1_n182 ) );
  OR2_X1 u0_u2_u1_U36 (.A2( u0_u2_u1_n157 ) , .A1( u0_u2_u1_n158 ) , .ZN( u0_u2_u1_n163 ) );
  OAI21_X1 u0_u2_u1_U37 (.B2( u0_u2_u1_n123 ) , .ZN( u0_u2_u1_n145 ) , .B1( u0_u2_u1_n160 ) , .A( u0_u2_u1_n185 ) );
  INV_X1 u0_u2_u1_U38 (.A( u0_u2_u1_n122 ) , .ZN( u0_u2_u1_n185 ) );
  AOI21_X1 u0_u2_u1_U39 (.B2( u0_u2_u1_n120 ) , .B1( u0_u2_u1_n121 ) , .ZN( u0_u2_u1_n122 ) , .A( u0_u2_u1_n128 ) );
  AOI221_X1 u0_u2_u1_U4 (.A( u0_u2_u1_n138 ) , .C2( u0_u2_u1_n139 ) , .C1( u0_u2_u1_n140 ) , .B2( u0_u2_u1_n141 ) , .ZN( u0_u2_u1_n142 ) , .B1( u0_u2_u1_n175 ) );
  NAND2_X1 u0_u2_u1_U40 (.A1( u0_u2_u1_n128 ) , .ZN( u0_u2_u1_n146 ) , .A2( u0_u2_u1_n160 ) );
  NAND2_X1 u0_u2_u1_U41 (.A2( u0_u2_u1_n112 ) , .ZN( u0_u2_u1_n139 ) , .A1( u0_u2_u1_n152 ) );
  NAND2_X1 u0_u2_u1_U42 (.A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n156 ) , .A2( u0_u2_u1_n99 ) );
  AOI221_X1 u0_u2_u1_U43 (.B1( u0_u2_u1_n140 ) , .ZN( u0_u2_u1_n167 ) , .B2( u0_u2_u1_n172 ) , .C2( u0_u2_u1_n175 ) , .C1( u0_u2_u1_n178 ) , .A( u0_u2_u1_n188 ) );
  INV_X1 u0_u2_u1_U44 (.ZN( u0_u2_u1_n188 ) , .A( u0_u2_u1_n97 ) );
  AOI211_X1 u0_u2_u1_U45 (.A( u0_u2_u1_n118 ) , .C1( u0_u2_u1_n132 ) , .C2( u0_u2_u1_n139 ) , .B( u0_u2_u1_n96 ) , .ZN( u0_u2_u1_n97 ) );
  AOI21_X1 u0_u2_u1_U46 (.B2( u0_u2_u1_n121 ) , .B1( u0_u2_u1_n135 ) , .A( u0_u2_u1_n152 ) , .ZN( u0_u2_u1_n96 ) );
  NOR2_X1 u0_u2_u1_U47 (.ZN( u0_u2_u1_n117 ) , .A1( u0_u2_u1_n121 ) , .A2( u0_u2_u1_n160 ) );
  AOI21_X1 u0_u2_u1_U48 (.A( u0_u2_u1_n128 ) , .B2( u0_u2_u1_n129 ) , .ZN( u0_u2_u1_n130 ) , .B1( u0_u2_u1_n150 ) );
  NAND2_X1 u0_u2_u1_U49 (.ZN( u0_u2_u1_n112 ) , .A1( u0_u2_u1_n169 ) , .A2( u0_u2_u1_n170 ) );
  AOI211_X1 u0_u2_u1_U5 (.ZN( u0_u2_u1_n124 ) , .A( u0_u2_u1_n138 ) , .C2( u0_u2_u1_n139 ) , .B( u0_u2_u1_n145 ) , .C1( u0_u2_u1_n147 ) );
  NAND2_X1 u0_u2_u1_U50 (.ZN( u0_u2_u1_n129 ) , .A2( u0_u2_u1_n95 ) , .A1( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U51 (.A1( u0_u2_u1_n102 ) , .ZN( u0_u2_u1_n154 ) , .A2( u0_u2_u1_n99 ) );
  NAND2_X1 u0_u2_u1_U52 (.A2( u0_u2_u1_n100 ) , .ZN( u0_u2_u1_n135 ) , .A1( u0_u2_u1_n99 ) );
  AOI21_X1 u0_u2_u1_U53 (.A( u0_u2_u1_n152 ) , .B2( u0_u2_u1_n153 ) , .B1( u0_u2_u1_n154 ) , .ZN( u0_u2_u1_n158 ) );
  INV_X1 u0_u2_u1_U54 (.A( u0_u2_u1_n160 ) , .ZN( u0_u2_u1_n175 ) );
  NAND2_X1 u0_u2_u1_U55 (.A1( u0_u2_u1_n100 ) , .ZN( u0_u2_u1_n116 ) , .A2( u0_u2_u1_n95 ) );
  NAND2_X1 u0_u2_u1_U56 (.A1( u0_u2_u1_n102 ) , .ZN( u0_u2_u1_n131 ) , .A2( u0_u2_u1_n95 ) );
  NAND2_X1 u0_u2_u1_U57 (.A2( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n121 ) , .A1( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U58 (.A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n153 ) , .A2( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U59 (.A2( u0_u2_u1_n104 ) , .A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n133 ) );
  AOI22_X1 u0_u2_u1_U6 (.B2( u0_u2_u1_n113 ) , .A2( u0_u2_u1_n114 ) , .ZN( u0_u2_u1_n125 ) , .A1( u0_u2_u1_n171 ) , .B1( u0_u2_u1_n173 ) );
  NAND2_X1 u0_u2_u1_U60 (.ZN( u0_u2_u1_n150 ) , .A2( u0_u2_u1_n98 ) , .A1( u0_u2_u1_n99 ) );
  NAND2_X1 u0_u2_u1_U61 (.A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n155 ) , .A2( u0_u2_u1_n95 ) );
  OAI21_X1 u0_u2_u1_U62 (.ZN( u0_u2_u1_n109 ) , .B1( u0_u2_u1_n129 ) , .B2( u0_u2_u1_n160 ) , .A( u0_u2_u1_n167 ) );
  NAND2_X1 u0_u2_u1_U63 (.A2( u0_u2_u1_n100 ) , .A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n120 ) );
  NAND2_X1 u0_u2_u1_U64 (.A1( u0_u2_u1_n102 ) , .A2( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n115 ) );
  NAND2_X1 u0_u2_u1_U65 (.A2( u0_u2_u1_n100 ) , .A1( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n151 ) );
  NAND2_X1 u0_u2_u1_U66 (.A2( u0_u2_u1_n103 ) , .A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n161 ) );
  INV_X1 u0_u2_u1_U67 (.A( u0_u2_u1_n152 ) , .ZN( u0_u2_u1_n173 ) );
  INV_X1 u0_u2_u1_U68 (.A( u0_u2_u1_n128 ) , .ZN( u0_u2_u1_n172 ) );
  NAND2_X1 u0_u2_u1_U69 (.A2( u0_u2_u1_n102 ) , .A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n123 ) );
  NAND2_X1 u0_u2_u1_U7 (.ZN( u0_u2_u1_n114 ) , .A1( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n156 ) );
  NOR2_X1 u0_u2_u1_U70 (.A2( u0_u2_X_7 ) , .A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n95 ) );
  NOR2_X1 u0_u2_u1_U71 (.A1( u0_u2_X_12 ) , .A2( u0_u2_X_9 ) , .ZN( u0_u2_u1_n100 ) );
  NOR2_X1 u0_u2_u1_U72 (.A2( u0_u2_X_8 ) , .A1( u0_u2_u1_n177 ) , .ZN( u0_u2_u1_n99 ) );
  NOR2_X1 u0_u2_u1_U73 (.A2( u0_u2_X_12 ) , .ZN( u0_u2_u1_n102 ) , .A1( u0_u2_u1_n176 ) );
  NOR2_X1 u0_u2_u1_U74 (.A2( u0_u2_X_9 ) , .ZN( u0_u2_u1_n105 ) , .A1( u0_u2_u1_n168 ) );
  NAND2_X1 u0_u2_u1_U75 (.A1( u0_u2_X_10 ) , .ZN( u0_u2_u1_n160 ) , .A2( u0_u2_u1_n169 ) );
  NAND2_X1 u0_u2_u1_U76 (.A2( u0_u2_X_10 ) , .A1( u0_u2_X_11 ) , .ZN( u0_u2_u1_n152 ) );
  NAND2_X1 u0_u2_u1_U77 (.A1( u0_u2_X_11 ) , .ZN( u0_u2_u1_n128 ) , .A2( u0_u2_u1_n170 ) );
  AND2_X1 u0_u2_u1_U78 (.A2( u0_u2_X_7 ) , .A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n104 ) );
  AND2_X1 u0_u2_u1_U79 (.A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n103 ) , .A2( u0_u2_u1_n177 ) );
  AOI22_X1 u0_u2_u1_U8 (.B2( u0_u2_u1_n136 ) , .A2( u0_u2_u1_n137 ) , .ZN( u0_u2_u1_n143 ) , .A1( u0_u2_u1_n171 ) , .B1( u0_u2_u1_n173 ) );
  INV_X1 u0_u2_u1_U80 (.A( u0_u2_X_10 ) , .ZN( u0_u2_u1_n170 ) );
  INV_X1 u0_u2_u1_U81 (.A( u0_u2_X_9 ) , .ZN( u0_u2_u1_n176 ) );
  INV_X1 u0_u2_u1_U82 (.A( u0_u2_X_11 ) , .ZN( u0_u2_u1_n169 ) );
  INV_X1 u0_u2_u1_U83 (.A( u0_u2_X_12 ) , .ZN( u0_u2_u1_n168 ) );
  INV_X1 u0_u2_u1_U84 (.A( u0_u2_X_7 ) , .ZN( u0_u2_u1_n177 ) );
  NAND4_X1 u0_u2_u1_U85 (.ZN( u0_out2_28 ) , .A4( u0_u2_u1_n124 ) , .A3( u0_u2_u1_n125 ) , .A2( u0_u2_u1_n126 ) , .A1( u0_u2_u1_n127 ) );
  OAI21_X1 u0_u2_u1_U86 (.ZN( u0_u2_u1_n127 ) , .B2( u0_u2_u1_n139 ) , .B1( u0_u2_u1_n175 ) , .A( u0_u2_u1_n183 ) );
  OAI21_X1 u0_u2_u1_U87 (.ZN( u0_u2_u1_n126 ) , .B2( u0_u2_u1_n140 ) , .A( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n178 ) );
  NAND4_X1 u0_u2_u1_U88 (.ZN( u0_out2_18 ) , .A4( u0_u2_u1_n165 ) , .A3( u0_u2_u1_n166 ) , .A1( u0_u2_u1_n167 ) , .A2( u0_u2_u1_n186 ) );
  AOI22_X1 u0_u2_u1_U89 (.B2( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n147 ) , .A2( u0_u2_u1_n148 ) , .ZN( u0_u2_u1_n166 ) , .A1( u0_u2_u1_n172 ) );
  INV_X1 u0_u2_u1_U9 (.A( u0_u2_u1_n147 ) , .ZN( u0_u2_u1_n181 ) );
  INV_X1 u0_u2_u1_U90 (.A( u0_u2_u1_n145 ) , .ZN( u0_u2_u1_n186 ) );
  NAND4_X1 u0_u2_u1_U91 (.ZN( u0_out2_2 ) , .A4( u0_u2_u1_n142 ) , .A3( u0_u2_u1_n143 ) , .A2( u0_u2_u1_n144 ) , .A1( u0_u2_u1_n179 ) );
  OAI21_X1 u0_u2_u1_U92 (.B2( u0_u2_u1_n132 ) , .ZN( u0_u2_u1_n144 ) , .A( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n180 ) );
  INV_X1 u0_u2_u1_U93 (.A( u0_u2_u1_n130 ) , .ZN( u0_u2_u1_n179 ) );
  OR4_X1 u0_u2_u1_U94 (.ZN( u0_out2_13 ) , .A4( u0_u2_u1_n108 ) , .A3( u0_u2_u1_n109 ) , .A2( u0_u2_u1_n110 ) , .A1( u0_u2_u1_n111 ) );
  AOI21_X1 u0_u2_u1_U95 (.ZN( u0_u2_u1_n111 ) , .A( u0_u2_u1_n128 ) , .B2( u0_u2_u1_n131 ) , .B1( u0_u2_u1_n135 ) );
  AOI21_X1 u0_u2_u1_U96 (.ZN( u0_u2_u1_n110 ) , .A( u0_u2_u1_n116 ) , .B1( u0_u2_u1_n152 ) , .B2( u0_u2_u1_n160 ) );
  NAND3_X1 u0_u2_u1_U97 (.A3( u0_u2_u1_n149 ) , .A2( u0_u2_u1_n150 ) , .A1( u0_u2_u1_n151 ) , .ZN( u0_u2_u1_n164 ) );
  NAND3_X1 u0_u2_u1_U98 (.A3( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n135 ) , .ZN( u0_u2_u1_n136 ) , .A1( u0_u2_u1_n151 ) );
  NAND3_X1 u0_u2_u1_U99 (.A1( u0_u2_u1_n133 ) , .ZN( u0_u2_u1_n137 ) , .A2( u0_u2_u1_n154 ) , .A3( u0_u2_u1_n181 ) );
  OAI22_X1 u0_u2_u2_U10 (.B1( u0_u2_u2_n151 ) , .A2( u0_u2_u2_n152 ) , .A1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n160 ) , .B2( u0_u2_u2_n168 ) );
  NAND3_X1 u0_u2_u2_U100 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n98 ) );
  NOR3_X1 u0_u2_u2_U11 (.A1( u0_u2_u2_n150 ) , .ZN( u0_u2_u2_n151 ) , .A3( u0_u2_u2_n175 ) , .A2( u0_u2_u2_n188 ) );
  AOI21_X1 u0_u2_u2_U12 (.B2( u0_u2_u2_n123 ) , .ZN( u0_u2_u2_n125 ) , .A( u0_u2_u2_n171 ) , .B1( u0_u2_u2_n184 ) );
  INV_X1 u0_u2_u2_U13 (.A( u0_u2_u2_n150 ) , .ZN( u0_u2_u2_n184 ) );
  AOI21_X1 u0_u2_u2_U14 (.ZN( u0_u2_u2_n144 ) , .B2( u0_u2_u2_n155 ) , .A( u0_u2_u2_n172 ) , .B1( u0_u2_u2_n185 ) );
  AOI21_X1 u0_u2_u2_U15 (.B2( u0_u2_u2_n143 ) , .ZN( u0_u2_u2_n145 ) , .B1( u0_u2_u2_n152 ) , .A( u0_u2_u2_n171 ) );
  INV_X1 u0_u2_u2_U16 (.A( u0_u2_u2_n156 ) , .ZN( u0_u2_u2_n171 ) );
  INV_X1 u0_u2_u2_U17 (.A( u0_u2_u2_n120 ) , .ZN( u0_u2_u2_n188 ) );
  NAND2_X1 u0_u2_u2_U18 (.A2( u0_u2_u2_n122 ) , .ZN( u0_u2_u2_n150 ) , .A1( u0_u2_u2_n152 ) );
  INV_X1 u0_u2_u2_U19 (.A( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n170 ) );
  INV_X1 u0_u2_u2_U20 (.A( u0_u2_u2_n137 ) , .ZN( u0_u2_u2_n173 ) );
  NAND2_X1 u0_u2_u2_U21 (.A1( u0_u2_u2_n132 ) , .A2( u0_u2_u2_n139 ) , .ZN( u0_u2_u2_n157 ) );
  INV_X1 u0_u2_u2_U22 (.A( u0_u2_u2_n113 ) , .ZN( u0_u2_u2_n178 ) );
  INV_X1 u0_u2_u2_U23 (.A( u0_u2_u2_n139 ) , .ZN( u0_u2_u2_n175 ) );
  INV_X1 u0_u2_u2_U24 (.A( u0_u2_u2_n155 ) , .ZN( u0_u2_u2_n181 ) );
  INV_X1 u0_u2_u2_U25 (.A( u0_u2_u2_n119 ) , .ZN( u0_u2_u2_n177 ) );
  INV_X1 u0_u2_u2_U26 (.A( u0_u2_u2_n116 ) , .ZN( u0_u2_u2_n180 ) );
  INV_X1 u0_u2_u2_U27 (.A( u0_u2_u2_n131 ) , .ZN( u0_u2_u2_n179 ) );
  INV_X1 u0_u2_u2_U28 (.A( u0_u2_u2_n154 ) , .ZN( u0_u2_u2_n176 ) );
  NAND2_X1 u0_u2_u2_U29 (.A2( u0_u2_u2_n116 ) , .A1( u0_u2_u2_n117 ) , .ZN( u0_u2_u2_n118 ) );
  NOR2_X1 u0_u2_u2_U3 (.ZN( u0_u2_u2_n121 ) , .A2( u0_u2_u2_n177 ) , .A1( u0_u2_u2_n180 ) );
  INV_X1 u0_u2_u2_U30 (.A( u0_u2_u2_n132 ) , .ZN( u0_u2_u2_n182 ) );
  INV_X1 u0_u2_u2_U31 (.A( u0_u2_u2_n158 ) , .ZN( u0_u2_u2_n183 ) );
  OAI21_X1 u0_u2_u2_U32 (.A( u0_u2_u2_n156 ) , .B1( u0_u2_u2_n157 ) , .ZN( u0_u2_u2_n158 ) , .B2( u0_u2_u2_n179 ) );
  NOR2_X1 u0_u2_u2_U33 (.ZN( u0_u2_u2_n156 ) , .A1( u0_u2_u2_n166 ) , .A2( u0_u2_u2_n169 ) );
  NOR2_X1 u0_u2_u2_U34 (.A2( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n137 ) , .A1( u0_u2_u2_n140 ) );
  NOR2_X1 u0_u2_u2_U35 (.A2( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n153 ) , .A1( u0_u2_u2_n156 ) );
  AOI211_X1 u0_u2_u2_U36 (.ZN( u0_u2_u2_n130 ) , .C1( u0_u2_u2_n138 ) , .C2( u0_u2_u2_n179 ) , .B( u0_u2_u2_n96 ) , .A( u0_u2_u2_n97 ) );
  OAI22_X1 u0_u2_u2_U37 (.B1( u0_u2_u2_n133 ) , .A2( u0_u2_u2_n137 ) , .A1( u0_u2_u2_n152 ) , .B2( u0_u2_u2_n168 ) , .ZN( u0_u2_u2_n97 ) );
  OAI221_X1 u0_u2_u2_U38 (.B1( u0_u2_u2_n113 ) , .C1( u0_u2_u2_n132 ) , .A( u0_u2_u2_n149 ) , .B2( u0_u2_u2_n171 ) , .C2( u0_u2_u2_n172 ) , .ZN( u0_u2_u2_n96 ) );
  OAI221_X1 u0_u2_u2_U39 (.A( u0_u2_u2_n115 ) , .C2( u0_u2_u2_n123 ) , .B2( u0_u2_u2_n143 ) , .B1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n163 ) , .C1( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U4 (.A( u0_u2_u2_n134 ) , .ZN( u0_u2_u2_n185 ) );
  OAI21_X1 u0_u2_u2_U40 (.A( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n115 ) , .B1( u0_u2_u2_n176 ) , .B2( u0_u2_u2_n178 ) );
  OAI221_X1 u0_u2_u2_U41 (.A( u0_u2_u2_n135 ) , .B2( u0_u2_u2_n136 ) , .B1( u0_u2_u2_n137 ) , .ZN( u0_u2_u2_n162 ) , .C2( u0_u2_u2_n167 ) , .C1( u0_u2_u2_n185 ) );
  AND3_X1 u0_u2_u2_U42 (.A3( u0_u2_u2_n131 ) , .A2( u0_u2_u2_n132 ) , .A1( u0_u2_u2_n133 ) , .ZN( u0_u2_u2_n136 ) );
  AOI22_X1 u0_u2_u2_U43 (.ZN( u0_u2_u2_n135 ) , .B1( u0_u2_u2_n140 ) , .A1( u0_u2_u2_n156 ) , .B2( u0_u2_u2_n180 ) , .A2( u0_u2_u2_n188 ) );
  AOI21_X1 u0_u2_u2_U44 (.ZN( u0_u2_u2_n149 ) , .B1( u0_u2_u2_n173 ) , .B2( u0_u2_u2_n188 ) , .A( u0_u2_u2_n95 ) );
  AND3_X1 u0_u2_u2_U45 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n156 ) , .ZN( u0_u2_u2_n95 ) );
  OAI21_X1 u0_u2_u2_U46 (.A( u0_u2_u2_n141 ) , .B2( u0_u2_u2_n142 ) , .ZN( u0_u2_u2_n146 ) , .B1( u0_u2_u2_n153 ) );
  OAI21_X1 u0_u2_u2_U47 (.A( u0_u2_u2_n140 ) , .ZN( u0_u2_u2_n141 ) , .B1( u0_u2_u2_n176 ) , .B2( u0_u2_u2_n177 ) );
  NOR3_X1 u0_u2_u2_U48 (.ZN( u0_u2_u2_n142 ) , .A3( u0_u2_u2_n175 ) , .A2( u0_u2_u2_n178 ) , .A1( u0_u2_u2_n181 ) );
  OAI21_X1 u0_u2_u2_U49 (.A( u0_u2_u2_n101 ) , .B2( u0_u2_u2_n121 ) , .B1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n164 ) );
  NOR4_X1 u0_u2_u2_U5 (.A4( u0_u2_u2_n124 ) , .A3( u0_u2_u2_n125 ) , .A2( u0_u2_u2_n126 ) , .A1( u0_u2_u2_n127 ) , .ZN( u0_u2_u2_n128 ) );
  NAND2_X1 u0_u2_u2_U50 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n155 ) );
  NAND2_X1 u0_u2_u2_U51 (.A2( u0_u2_u2_n105 ) , .A1( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n143 ) );
  NAND2_X1 u0_u2_u2_U52 (.A1( u0_u2_u2_n104 ) , .A2( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n152 ) );
  NAND2_X1 u0_u2_u2_U53 (.A1( u0_u2_u2_n100 ) , .A2( u0_u2_u2_n105 ) , .ZN( u0_u2_u2_n132 ) );
  INV_X1 u0_u2_u2_U54 (.A( u0_u2_u2_n140 ) , .ZN( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U55 (.A( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n167 ) );
  INV_X1 u0_u2_u2_U56 (.ZN( u0_u2_u2_n187 ) , .A( u0_u2_u2_n99 ) );
  OAI21_X1 u0_u2_u2_U57 (.B1( u0_u2_u2_n137 ) , .B2( u0_u2_u2_n143 ) , .A( u0_u2_u2_n98 ) , .ZN( u0_u2_u2_n99 ) );
  NAND2_X1 u0_u2_u2_U58 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n113 ) );
  NAND2_X1 u0_u2_u2_U59 (.A1( u0_u2_u2_n106 ) , .A2( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n131 ) );
  AOI21_X1 u0_u2_u2_U6 (.B2( u0_u2_u2_n119 ) , .ZN( u0_u2_u2_n127 ) , .A( u0_u2_u2_n137 ) , .B1( u0_u2_u2_n155 ) );
  NAND2_X1 u0_u2_u2_U60 (.A1( u0_u2_u2_n103 ) , .A2( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n139 ) );
  NAND2_X1 u0_u2_u2_U61 (.A1( u0_u2_u2_n103 ) , .A2( u0_u2_u2_n105 ) , .ZN( u0_u2_u2_n133 ) );
  NAND2_X1 u0_u2_u2_U62 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n103 ) , .ZN( u0_u2_u2_n154 ) );
  NAND2_X1 u0_u2_u2_U63 (.A2( u0_u2_u2_n103 ) , .A1( u0_u2_u2_n104 ) , .ZN( u0_u2_u2_n119 ) );
  NAND2_X1 u0_u2_u2_U64 (.A2( u0_u2_u2_n107 ) , .A1( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n123 ) );
  NAND2_X1 u0_u2_u2_U65 (.A1( u0_u2_u2_n104 ) , .A2( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n122 ) );
  INV_X1 u0_u2_u2_U66 (.A( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n172 ) );
  NAND2_X1 u0_u2_u2_U67 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n102 ) , .ZN( u0_u2_u2_n116 ) );
  NAND2_X1 u0_u2_u2_U68 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n120 ) );
  NAND2_X1 u0_u2_u2_U69 (.A2( u0_u2_u2_n105 ) , .A1( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n117 ) );
  AOI21_X1 u0_u2_u2_U7 (.ZN( u0_u2_u2_n124 ) , .B1( u0_u2_u2_n131 ) , .B2( u0_u2_u2_n143 ) , .A( u0_u2_u2_n172 ) );
  NOR2_X1 u0_u2_u2_U70 (.A2( u0_u2_X_16 ) , .ZN( u0_u2_u2_n140 ) , .A1( u0_u2_u2_n166 ) );
  NOR2_X1 u0_u2_u2_U71 (.A2( u0_u2_X_13 ) , .A1( u0_u2_X_14 ) , .ZN( u0_u2_u2_n100 ) );
  NOR2_X1 u0_u2_u2_U72 (.A2( u0_u2_X_16 ) , .A1( u0_u2_X_17 ) , .ZN( u0_u2_u2_n138 ) );
  NOR2_X1 u0_u2_u2_U73 (.A2( u0_u2_X_15 ) , .A1( u0_u2_X_18 ) , .ZN( u0_u2_u2_n104 ) );
  NOR2_X1 u0_u2_u2_U74 (.A2( u0_u2_X_14 ) , .ZN( u0_u2_u2_n103 ) , .A1( u0_u2_u2_n174 ) );
  NOR2_X1 u0_u2_u2_U75 (.A2( u0_u2_X_15 ) , .ZN( u0_u2_u2_n102 ) , .A1( u0_u2_u2_n165 ) );
  NOR2_X1 u0_u2_u2_U76 (.A2( u0_u2_X_17 ) , .ZN( u0_u2_u2_n114 ) , .A1( u0_u2_u2_n169 ) );
  AND2_X1 u0_u2_u2_U77 (.A1( u0_u2_X_15 ) , .ZN( u0_u2_u2_n105 ) , .A2( u0_u2_u2_n165 ) );
  AND2_X1 u0_u2_u2_U78 (.A2( u0_u2_X_15 ) , .A1( u0_u2_X_18 ) , .ZN( u0_u2_u2_n107 ) );
  AND2_X1 u0_u2_u2_U79 (.A1( u0_u2_X_14 ) , .ZN( u0_u2_u2_n106 ) , .A2( u0_u2_u2_n174 ) );
  AOI21_X1 u0_u2_u2_U8 (.B2( u0_u2_u2_n120 ) , .B1( u0_u2_u2_n121 ) , .ZN( u0_u2_u2_n126 ) , .A( u0_u2_u2_n167 ) );
  AND2_X1 u0_u2_u2_U80 (.A1( u0_u2_X_13 ) , .A2( u0_u2_X_14 ) , .ZN( u0_u2_u2_n108 ) );
  INV_X1 u0_u2_u2_U81 (.A( u0_u2_X_16 ) , .ZN( u0_u2_u2_n169 ) );
  INV_X1 u0_u2_u2_U82 (.A( u0_u2_X_17 ) , .ZN( u0_u2_u2_n166 ) );
  INV_X1 u0_u2_u2_U83 (.A( u0_u2_X_13 ) , .ZN( u0_u2_u2_n174 ) );
  INV_X1 u0_u2_u2_U84 (.A( u0_u2_X_18 ) , .ZN( u0_u2_u2_n165 ) );
  NAND4_X1 u0_u2_u2_U85 (.ZN( u0_out2_24 ) , .A4( u0_u2_u2_n111 ) , .A3( u0_u2_u2_n112 ) , .A1( u0_u2_u2_n130 ) , .A2( u0_u2_u2_n187 ) );
  AOI21_X1 u0_u2_u2_U86 (.ZN( u0_u2_u2_n112 ) , .B2( u0_u2_u2_n156 ) , .A( u0_u2_u2_n164 ) , .B1( u0_u2_u2_n181 ) );
  AOI221_X1 u0_u2_u2_U87 (.A( u0_u2_u2_n109 ) , .B1( u0_u2_u2_n110 ) , .ZN( u0_u2_u2_n111 ) , .C1( u0_u2_u2_n134 ) , .C2( u0_u2_u2_n170 ) , .B2( u0_u2_u2_n173 ) );
  NAND4_X1 u0_u2_u2_U88 (.ZN( u0_out2_16 ) , .A4( u0_u2_u2_n128 ) , .A3( u0_u2_u2_n129 ) , .A1( u0_u2_u2_n130 ) , .A2( u0_u2_u2_n186 ) );
  AOI22_X1 u0_u2_u2_U89 (.A2( u0_u2_u2_n118 ) , .ZN( u0_u2_u2_n129 ) , .A1( u0_u2_u2_n140 ) , .B1( u0_u2_u2_n157 ) , .B2( u0_u2_u2_n170 ) );
  OAI22_X1 u0_u2_u2_U9 (.ZN( u0_u2_u2_n109 ) , .A2( u0_u2_u2_n113 ) , .B2( u0_u2_u2_n133 ) , .B1( u0_u2_u2_n167 ) , .A1( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U90 (.A( u0_u2_u2_n163 ) , .ZN( u0_u2_u2_n186 ) );
  NAND4_X1 u0_u2_u2_U91 (.ZN( u0_out2_30 ) , .A4( u0_u2_u2_n147 ) , .A3( u0_u2_u2_n148 ) , .A2( u0_u2_u2_n149 ) , .A1( u0_u2_u2_n187 ) );
  NOR3_X1 u0_u2_u2_U92 (.A3( u0_u2_u2_n144 ) , .A2( u0_u2_u2_n145 ) , .A1( u0_u2_u2_n146 ) , .ZN( u0_u2_u2_n147 ) );
  AOI21_X1 u0_u2_u2_U93 (.B2( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n148 ) , .A( u0_u2_u2_n162 ) , .B1( u0_u2_u2_n182 ) );
  OR4_X1 u0_u2_u2_U94 (.ZN( u0_out2_6 ) , .A4( u0_u2_u2_n161 ) , .A3( u0_u2_u2_n162 ) , .A2( u0_u2_u2_n163 ) , .A1( u0_u2_u2_n164 ) );
  OR3_X1 u0_u2_u2_U95 (.A2( u0_u2_u2_n159 ) , .A1( u0_u2_u2_n160 ) , .ZN( u0_u2_u2_n161 ) , .A3( u0_u2_u2_n183 ) );
  AOI21_X1 u0_u2_u2_U96 (.B2( u0_u2_u2_n154 ) , .B1( u0_u2_u2_n155 ) , .ZN( u0_u2_u2_n159 ) , .A( u0_u2_u2_n167 ) );
  NAND3_X1 u0_u2_u2_U97 (.A2( u0_u2_u2_n117 ) , .A1( u0_u2_u2_n122 ) , .A3( u0_u2_u2_n123 ) , .ZN( u0_u2_u2_n134 ) );
  NAND3_X1 u0_u2_u2_U98 (.ZN( u0_u2_u2_n110 ) , .A2( u0_u2_u2_n131 ) , .A3( u0_u2_u2_n139 ) , .A1( u0_u2_u2_n154 ) );
  NAND3_X1 u0_u2_u2_U99 (.A2( u0_u2_u2_n100 ) , .ZN( u0_u2_u2_n101 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n114 ) );
  OAI22_X1 u0_u2_u3_U10 (.B1( u0_u2_u3_n113 ) , .A2( u0_u2_u3_n135 ) , .A1( u0_u2_u3_n150 ) , .B2( u0_u2_u3_n164 ) , .ZN( u0_u2_u3_n98 ) );
  OAI211_X1 u0_u2_u3_U11 (.B( u0_u2_u3_n106 ) , .ZN( u0_u2_u3_n119 ) , .C2( u0_u2_u3_n128 ) , .C1( u0_u2_u3_n167 ) , .A( u0_u2_u3_n181 ) );
  AOI221_X1 u0_u2_u3_U12 (.C1( u0_u2_u3_n105 ) , .ZN( u0_u2_u3_n106 ) , .A( u0_u2_u3_n131 ) , .B2( u0_u2_u3_n132 ) , .C2( u0_u2_u3_n133 ) , .B1( u0_u2_u3_n169 ) );
  INV_X1 u0_u2_u3_U13 (.ZN( u0_u2_u3_n181 ) , .A( u0_u2_u3_n98 ) );
  NAND2_X1 u0_u2_u3_U14 (.ZN( u0_u2_u3_n105 ) , .A2( u0_u2_u3_n130 ) , .A1( u0_u2_u3_n155 ) );
  AOI22_X1 u0_u2_u3_U15 (.B1( u0_u2_u3_n115 ) , .A2( u0_u2_u3_n116 ) , .ZN( u0_u2_u3_n123 ) , .B2( u0_u2_u3_n133 ) , .A1( u0_u2_u3_n169 ) );
  NAND2_X1 u0_u2_u3_U16 (.ZN( u0_u2_u3_n116 ) , .A2( u0_u2_u3_n151 ) , .A1( u0_u2_u3_n182 ) );
  NOR2_X1 u0_u2_u3_U17 (.ZN( u0_u2_u3_n126 ) , .A2( u0_u2_u3_n150 ) , .A1( u0_u2_u3_n164 ) );
  AOI21_X1 u0_u2_u3_U18 (.ZN( u0_u2_u3_n112 ) , .B2( u0_u2_u3_n146 ) , .B1( u0_u2_u3_n155 ) , .A( u0_u2_u3_n167 ) );
  NAND2_X1 u0_u2_u3_U19 (.A1( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n142 ) , .A2( u0_u2_u3_n164 ) );
  NAND2_X1 u0_u2_u3_U20 (.ZN( u0_u2_u3_n132 ) , .A2( u0_u2_u3_n152 ) , .A1( u0_u2_u3_n156 ) );
  AND2_X1 u0_u2_u3_U21 (.A2( u0_u2_u3_n113 ) , .A1( u0_u2_u3_n114 ) , .ZN( u0_u2_u3_n151 ) );
  INV_X1 u0_u2_u3_U22 (.A( u0_u2_u3_n133 ) , .ZN( u0_u2_u3_n165 ) );
  INV_X1 u0_u2_u3_U23 (.A( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n170 ) );
  NAND2_X1 u0_u2_u3_U24 (.A1( u0_u2_u3_n107 ) , .A2( u0_u2_u3_n108 ) , .ZN( u0_u2_u3_n140 ) );
  NAND2_X1 u0_u2_u3_U25 (.ZN( u0_u2_u3_n117 ) , .A1( u0_u2_u3_n124 ) , .A2( u0_u2_u3_n148 ) );
  NAND2_X1 u0_u2_u3_U26 (.ZN( u0_u2_u3_n143 ) , .A1( u0_u2_u3_n165 ) , .A2( u0_u2_u3_n167 ) );
  INV_X1 u0_u2_u3_U27 (.A( u0_u2_u3_n130 ) , .ZN( u0_u2_u3_n177 ) );
  INV_X1 u0_u2_u3_U28 (.A( u0_u2_u3_n128 ) , .ZN( u0_u2_u3_n176 ) );
  INV_X1 u0_u2_u3_U29 (.A( u0_u2_u3_n155 ) , .ZN( u0_u2_u3_n174 ) );
  INV_X1 u0_u2_u3_U3 (.A( u0_u2_u3_n129 ) , .ZN( u0_u2_u3_n183 ) );
  INV_X1 u0_u2_u3_U30 (.A( u0_u2_u3_n139 ) , .ZN( u0_u2_u3_n185 ) );
  NOR2_X1 u0_u2_u3_U31 (.ZN( u0_u2_u3_n135 ) , .A2( u0_u2_u3_n141 ) , .A1( u0_u2_u3_n169 ) );
  OAI222_X1 u0_u2_u3_U32 (.C2( u0_u2_u3_n107 ) , .A2( u0_u2_u3_n108 ) , .B1( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n138 ) , .B2( u0_u2_u3_n146 ) , .C1( u0_u2_u3_n154 ) , .A1( u0_u2_u3_n164 ) );
  NOR4_X1 u0_u2_u3_U33 (.A4( u0_u2_u3_n157 ) , .A3( u0_u2_u3_n158 ) , .A2( u0_u2_u3_n159 ) , .A1( u0_u2_u3_n160 ) , .ZN( u0_u2_u3_n161 ) );
  AOI21_X1 u0_u2_u3_U34 (.B2( u0_u2_u3_n152 ) , .B1( u0_u2_u3_n153 ) , .ZN( u0_u2_u3_n158 ) , .A( u0_u2_u3_n164 ) );
  AOI21_X1 u0_u2_u3_U35 (.A( u0_u2_u3_n154 ) , .B2( u0_u2_u3_n155 ) , .B1( u0_u2_u3_n156 ) , .ZN( u0_u2_u3_n157 ) );
  AOI21_X1 u0_u2_u3_U36 (.A( u0_u2_u3_n149 ) , .B2( u0_u2_u3_n150 ) , .B1( u0_u2_u3_n151 ) , .ZN( u0_u2_u3_n159 ) );
  AOI211_X1 u0_u2_u3_U37 (.ZN( u0_u2_u3_n109 ) , .A( u0_u2_u3_n119 ) , .C2( u0_u2_u3_n129 ) , .B( u0_u2_u3_n138 ) , .C1( u0_u2_u3_n141 ) );
  AOI211_X1 u0_u2_u3_U38 (.B( u0_u2_u3_n119 ) , .A( u0_u2_u3_n120 ) , .C2( u0_u2_u3_n121 ) , .ZN( u0_u2_u3_n122 ) , .C1( u0_u2_u3_n179 ) );
  INV_X1 u0_u2_u3_U39 (.A( u0_u2_u3_n156 ) , .ZN( u0_u2_u3_n179 ) );
  INV_X1 u0_u2_u3_U4 (.A( u0_u2_u3_n140 ) , .ZN( u0_u2_u3_n182 ) );
  OAI22_X1 u0_u2_u3_U40 (.B1( u0_u2_u3_n118 ) , .ZN( u0_u2_u3_n120 ) , .A1( u0_u2_u3_n135 ) , .B2( u0_u2_u3_n154 ) , .A2( u0_u2_u3_n178 ) );
  AND3_X1 u0_u2_u3_U41 (.ZN( u0_u2_u3_n118 ) , .A2( u0_u2_u3_n124 ) , .A1( u0_u2_u3_n144 ) , .A3( u0_u2_u3_n152 ) );
  INV_X1 u0_u2_u3_U42 (.A( u0_u2_u3_n121 ) , .ZN( u0_u2_u3_n164 ) );
  NAND2_X1 u0_u2_u3_U43 (.ZN( u0_u2_u3_n133 ) , .A1( u0_u2_u3_n154 ) , .A2( u0_u2_u3_n164 ) );
  OAI211_X1 u0_u2_u3_U44 (.B( u0_u2_u3_n127 ) , .ZN( u0_u2_u3_n139 ) , .C1( u0_u2_u3_n150 ) , .C2( u0_u2_u3_n154 ) , .A( u0_u2_u3_n184 ) );
  INV_X1 u0_u2_u3_U45 (.A( u0_u2_u3_n125 ) , .ZN( u0_u2_u3_n184 ) );
  AOI221_X1 u0_u2_u3_U46 (.A( u0_u2_u3_n126 ) , .ZN( u0_u2_u3_n127 ) , .C2( u0_u2_u3_n132 ) , .C1( u0_u2_u3_n169 ) , .B2( u0_u2_u3_n170 ) , .B1( u0_u2_u3_n174 ) );
  OAI22_X1 u0_u2_u3_U47 (.A1( u0_u2_u3_n124 ) , .ZN( u0_u2_u3_n125 ) , .B2( u0_u2_u3_n145 ) , .A2( u0_u2_u3_n165 ) , .B1( u0_u2_u3_n167 ) );
  NOR2_X1 u0_u2_u3_U48 (.A1( u0_u2_u3_n113 ) , .ZN( u0_u2_u3_n131 ) , .A2( u0_u2_u3_n154 ) );
  NAND2_X1 u0_u2_u3_U49 (.A1( u0_u2_u3_n103 ) , .ZN( u0_u2_u3_n150 ) , .A2( u0_u2_u3_n99 ) );
  INV_X1 u0_u2_u3_U5 (.A( u0_u2_u3_n117 ) , .ZN( u0_u2_u3_n178 ) );
  NAND2_X1 u0_u2_u3_U50 (.A2( u0_u2_u3_n102 ) , .ZN( u0_u2_u3_n155 ) , .A1( u0_u2_u3_n97 ) );
  INV_X1 u0_u2_u3_U51 (.A( u0_u2_u3_n141 ) , .ZN( u0_u2_u3_n167 ) );
  AOI21_X1 u0_u2_u3_U52 (.B2( u0_u2_u3_n114 ) , .B1( u0_u2_u3_n146 ) , .A( u0_u2_u3_n154 ) , .ZN( u0_u2_u3_n94 ) );
  AOI21_X1 u0_u2_u3_U53 (.ZN( u0_u2_u3_n110 ) , .B2( u0_u2_u3_n142 ) , .B1( u0_u2_u3_n186 ) , .A( u0_u2_u3_n95 ) );
  INV_X1 u0_u2_u3_U54 (.A( u0_u2_u3_n145 ) , .ZN( u0_u2_u3_n186 ) );
  AOI21_X1 u0_u2_u3_U55 (.B1( u0_u2_u3_n124 ) , .A( u0_u2_u3_n149 ) , .B2( u0_u2_u3_n155 ) , .ZN( u0_u2_u3_n95 ) );
  INV_X1 u0_u2_u3_U56 (.A( u0_u2_u3_n149 ) , .ZN( u0_u2_u3_n169 ) );
  NAND2_X1 u0_u2_u3_U57 (.ZN( u0_u2_u3_n124 ) , .A1( u0_u2_u3_n96 ) , .A2( u0_u2_u3_n97 ) );
  NAND2_X1 u0_u2_u3_U58 (.A2( u0_u2_u3_n100 ) , .ZN( u0_u2_u3_n146 ) , .A1( u0_u2_u3_n96 ) );
  NAND2_X1 u0_u2_u3_U59 (.A1( u0_u2_u3_n101 ) , .ZN( u0_u2_u3_n145 ) , .A2( u0_u2_u3_n99 ) );
  AOI221_X1 u0_u2_u3_U6 (.A( u0_u2_u3_n131 ) , .C2( u0_u2_u3_n132 ) , .C1( u0_u2_u3_n133 ) , .ZN( u0_u2_u3_n134 ) , .B1( u0_u2_u3_n143 ) , .B2( u0_u2_u3_n177 ) );
  NAND2_X1 u0_u2_u3_U60 (.A1( u0_u2_u3_n100 ) , .ZN( u0_u2_u3_n156 ) , .A2( u0_u2_u3_n99 ) );
  NAND2_X1 u0_u2_u3_U61 (.A2( u0_u2_u3_n101 ) , .A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n148 ) );
  NAND2_X1 u0_u2_u3_U62 (.A1( u0_u2_u3_n100 ) , .A2( u0_u2_u3_n102 ) , .ZN( u0_u2_u3_n128 ) );
  NAND2_X1 u0_u2_u3_U63 (.A2( u0_u2_u3_n101 ) , .A1( u0_u2_u3_n102 ) , .ZN( u0_u2_u3_n152 ) );
  NAND2_X1 u0_u2_u3_U64 (.A2( u0_u2_u3_n101 ) , .ZN( u0_u2_u3_n114 ) , .A1( u0_u2_u3_n96 ) );
  NAND2_X1 u0_u2_u3_U65 (.ZN( u0_u2_u3_n107 ) , .A1( u0_u2_u3_n97 ) , .A2( u0_u2_u3_n99 ) );
  NAND2_X1 u0_u2_u3_U66 (.A2( u0_u2_u3_n100 ) , .A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n113 ) );
  NAND2_X1 u0_u2_u3_U67 (.A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n153 ) , .A2( u0_u2_u3_n97 ) );
  NAND2_X1 u0_u2_u3_U68 (.A2( u0_u2_u3_n103 ) , .A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n130 ) );
  NAND2_X1 u0_u2_u3_U69 (.A2( u0_u2_u3_n103 ) , .ZN( u0_u2_u3_n144 ) , .A1( u0_u2_u3_n96 ) );
  OAI22_X1 u0_u2_u3_U7 (.B2( u0_u2_u3_n147 ) , .A2( u0_u2_u3_n148 ) , .ZN( u0_u2_u3_n160 ) , .B1( u0_u2_u3_n165 ) , .A1( u0_u2_u3_n168 ) );
  NAND2_X1 u0_u2_u3_U70 (.A1( u0_u2_u3_n102 ) , .A2( u0_u2_u3_n103 ) , .ZN( u0_u2_u3_n108 ) );
  NOR2_X1 u0_u2_u3_U71 (.A2( u0_u2_X_19 ) , .A1( u0_u2_X_20 ) , .ZN( u0_u2_u3_n99 ) );
  NOR2_X1 u0_u2_u3_U72 (.A2( u0_u2_X_21 ) , .A1( u0_u2_X_24 ) , .ZN( u0_u2_u3_n103 ) );
  NOR2_X1 u0_u2_u3_U73 (.A2( u0_u2_X_24 ) , .A1( u0_u2_u3_n171 ) , .ZN( u0_u2_u3_n97 ) );
  NOR2_X1 u0_u2_u3_U74 (.A2( u0_u2_X_23 ) , .ZN( u0_u2_u3_n141 ) , .A1( u0_u2_u3_n166 ) );
  NOR2_X1 u0_u2_u3_U75 (.A2( u0_u2_X_19 ) , .A1( u0_u2_u3_n172 ) , .ZN( u0_u2_u3_n96 ) );
  NAND2_X1 u0_u2_u3_U76 (.A1( u0_u2_X_22 ) , .A2( u0_u2_X_23 ) , .ZN( u0_u2_u3_n154 ) );
  NAND2_X1 u0_u2_u3_U77 (.A1( u0_u2_X_23 ) , .ZN( u0_u2_u3_n149 ) , .A2( u0_u2_u3_n166 ) );
  NOR2_X1 u0_u2_u3_U78 (.A2( u0_u2_X_22 ) , .A1( u0_u2_X_23 ) , .ZN( u0_u2_u3_n121 ) );
  AND2_X1 u0_u2_u3_U79 (.A1( u0_u2_X_24 ) , .ZN( u0_u2_u3_n101 ) , .A2( u0_u2_u3_n171 ) );
  AND3_X1 u0_u2_u3_U8 (.A3( u0_u2_u3_n144 ) , .A2( u0_u2_u3_n145 ) , .A1( u0_u2_u3_n146 ) , .ZN( u0_u2_u3_n147 ) );
  AND2_X1 u0_u2_u3_U80 (.A1( u0_u2_X_19 ) , .ZN( u0_u2_u3_n102 ) , .A2( u0_u2_u3_n172 ) );
  AND2_X1 u0_u2_u3_U81 (.A1( u0_u2_X_21 ) , .A2( u0_u2_X_24 ) , .ZN( u0_u2_u3_n100 ) );
  AND2_X1 u0_u2_u3_U82 (.A2( u0_u2_X_19 ) , .A1( u0_u2_X_20 ) , .ZN( u0_u2_u3_n104 ) );
  INV_X1 u0_u2_u3_U83 (.A( u0_u2_X_22 ) , .ZN( u0_u2_u3_n166 ) );
  INV_X1 u0_u2_u3_U84 (.A( u0_u2_X_21 ) , .ZN( u0_u2_u3_n171 ) );
  INV_X1 u0_u2_u3_U85 (.A( u0_u2_X_20 ) , .ZN( u0_u2_u3_n172 ) );
  OR4_X1 u0_u2_u3_U86 (.ZN( u0_out2_10 ) , .A4( u0_u2_u3_n136 ) , .A3( u0_u2_u3_n137 ) , .A1( u0_u2_u3_n138 ) , .A2( u0_u2_u3_n139 ) );
  OAI222_X1 u0_u2_u3_U87 (.C1( u0_u2_u3_n128 ) , .ZN( u0_u2_u3_n137 ) , .B1( u0_u2_u3_n148 ) , .A2( u0_u2_u3_n150 ) , .B2( u0_u2_u3_n154 ) , .C2( u0_u2_u3_n164 ) , .A1( u0_u2_u3_n167 ) );
  OAI221_X1 u0_u2_u3_U88 (.A( u0_u2_u3_n134 ) , .B2( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n136 ) , .C1( u0_u2_u3_n149 ) , .B1( u0_u2_u3_n151 ) , .C2( u0_u2_u3_n183 ) );
  NAND4_X1 u0_u2_u3_U89 (.ZN( u0_out2_26 ) , .A4( u0_u2_u3_n109 ) , .A3( u0_u2_u3_n110 ) , .A2( u0_u2_u3_n111 ) , .A1( u0_u2_u3_n173 ) );
  INV_X1 u0_u2_u3_U9 (.A( u0_u2_u3_n143 ) , .ZN( u0_u2_u3_n168 ) );
  INV_X1 u0_u2_u3_U90 (.ZN( u0_u2_u3_n173 ) , .A( u0_u2_u3_n94 ) );
  OAI21_X1 u0_u2_u3_U91 (.ZN( u0_u2_u3_n111 ) , .B2( u0_u2_u3_n117 ) , .A( u0_u2_u3_n133 ) , .B1( u0_u2_u3_n176 ) );
  NAND4_X1 u0_u2_u3_U92 (.ZN( u0_out2_20 ) , .A4( u0_u2_u3_n122 ) , .A3( u0_u2_u3_n123 ) , .A1( u0_u2_u3_n175 ) , .A2( u0_u2_u3_n180 ) );
  INV_X1 u0_u2_u3_U93 (.A( u0_u2_u3_n112 ) , .ZN( u0_u2_u3_n175 ) );
  INV_X1 u0_u2_u3_U94 (.A( u0_u2_u3_n126 ) , .ZN( u0_u2_u3_n180 ) );
  NAND4_X1 u0_u2_u3_U95 (.ZN( u0_out2_1 ) , .A4( u0_u2_u3_n161 ) , .A3( u0_u2_u3_n162 ) , .A2( u0_u2_u3_n163 ) , .A1( u0_u2_u3_n185 ) );
  NAND2_X1 u0_u2_u3_U96 (.ZN( u0_u2_u3_n163 ) , .A2( u0_u2_u3_n170 ) , .A1( u0_u2_u3_n176 ) );
  AOI22_X1 u0_u2_u3_U97 (.B2( u0_u2_u3_n140 ) , .B1( u0_u2_u3_n141 ) , .A2( u0_u2_u3_n142 ) , .ZN( u0_u2_u3_n162 ) , .A1( u0_u2_u3_n177 ) );
  NAND3_X1 u0_u2_u3_U98 (.A1( u0_u2_u3_n114 ) , .ZN( u0_u2_u3_n115 ) , .A2( u0_u2_u3_n145 ) , .A3( u0_u2_u3_n153 ) );
  NAND3_X1 u0_u2_u3_U99 (.ZN( u0_u2_u3_n129 ) , .A2( u0_u2_u3_n144 ) , .A1( u0_u2_u3_n153 ) , .A3( u0_u2_u3_n182 ) );
  XOR2_X1 u0_u3_U1 (.B( u0_K4_9 ) , .A( u0_R2_6 ) , .Z( u0_u3_X_9 ) );
  XOR2_X1 u0_u3_U16 (.B( u0_K4_3 ) , .A( u0_R2_2 ) , .Z( u0_u3_X_3 ) );
  XOR2_X1 u0_u3_U2 (.B( u0_K4_8 ) , .A( u0_R2_5 ) , .Z( u0_u3_X_8 ) );
  XOR2_X1 u0_u3_U20 (.B( u0_K4_36 ) , .A( u0_R2_25 ) , .Z( u0_u3_X_36 ) );
  XOR2_X1 u0_u3_U21 (.B( u0_K4_35 ) , .A( u0_R2_24 ) , .Z( u0_u3_X_35 ) );
  XOR2_X1 u0_u3_U22 (.B( u0_K4_34 ) , .A( u0_R2_23 ) , .Z( u0_u3_X_34 ) );
  XOR2_X1 u0_u3_U23 (.B( u0_K4_33 ) , .A( u0_R2_22 ) , .Z( u0_u3_X_33 ) );
  XOR2_X1 u0_u3_U24 (.B( u0_K4_32 ) , .A( u0_R2_21 ) , .Z( u0_u3_X_32 ) );
  XOR2_X1 u0_u3_U25 (.B( u0_K4_31 ) , .A( u0_R2_20 ) , .Z( u0_u3_X_31 ) );
  XOR2_X1 u0_u3_U26 (.B( u0_K4_30 ) , .A( u0_R2_21 ) , .Z( u0_u3_X_30 ) );
  XOR2_X1 u0_u3_U27 (.B( u0_K4_2 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_2 ) );
  XOR2_X1 u0_u3_U28 (.B( u0_K4_29 ) , .A( u0_R2_20 ) , .Z( u0_u3_X_29 ) );
  XOR2_X1 u0_u3_U29 (.B( u0_K4_28 ) , .A( u0_R2_19 ) , .Z( u0_u3_X_28 ) );
  XOR2_X1 u0_u3_U3 (.B( u0_K4_7 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_7 ) );
  XOR2_X1 u0_u3_U30 (.B( u0_K4_27 ) , .A( u0_R2_18 ) , .Z( u0_u3_X_27 ) );
  XOR2_X1 u0_u3_U31 (.B( u0_K4_26 ) , .A( u0_R2_17 ) , .Z( u0_u3_X_26 ) );
  XOR2_X1 u0_u3_U32 (.B( u0_K4_25 ) , .A( u0_R2_16 ) , .Z( u0_u3_X_25 ) );
  XOR2_X1 u0_u3_U33 (.B( u0_K4_24 ) , .A( u0_R2_17 ) , .Z( u0_u3_X_24 ) );
  XOR2_X1 u0_u3_U34 (.B( u0_K4_23 ) , .A( u0_R2_16 ) , .Z( u0_u3_X_23 ) );
  XOR2_X1 u0_u3_U35 (.B( u0_K4_22 ) , .A( u0_R2_15 ) , .Z( u0_u3_X_22 ) );
  XOR2_X1 u0_u3_U36 (.B( u0_K4_21 ) , .A( u0_R2_14 ) , .Z( u0_u3_X_21 ) );
  XOR2_X1 u0_u3_U37 (.B( u0_K4_20 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_20 ) );
  XOR2_X1 u0_u3_U38 (.B( u0_K4_1 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_1 ) );
  XOR2_X1 u0_u3_U39 (.B( u0_K4_19 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_19 ) );
  XOR2_X1 u0_u3_U4 (.B( u0_K4_6 ) , .A( u0_R2_5 ) , .Z( u0_u3_X_6 ) );
  XOR2_X1 u0_u3_U40 (.B( u0_K4_18 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_18 ) );
  XOR2_X1 u0_u3_U41 (.B( u0_K4_17 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_17 ) );
  XOR2_X1 u0_u3_U42 (.B( u0_K4_16 ) , .A( u0_R2_11 ) , .Z( u0_u3_X_16 ) );
  XOR2_X1 u0_u3_U43 (.B( u0_K4_15 ) , .A( u0_R2_10 ) , .Z( u0_u3_X_15 ) );
  XOR2_X1 u0_u3_U44 (.B( u0_K4_14 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_14 ) );
  XOR2_X1 u0_u3_U45 (.B( u0_K4_13 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_13 ) );
  XOR2_X1 u0_u3_U46 (.B( u0_K4_12 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_12 ) );
  XOR2_X1 u0_u3_U47 (.B( u0_K4_11 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_11 ) );
  XOR2_X1 u0_u3_U48 (.B( u0_K4_10 ) , .A( u0_R2_7 ) , .Z( u0_u3_X_10 ) );
  XOR2_X1 u0_u3_U5 (.B( u0_K4_5 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_5 ) );
  XOR2_X1 u0_u3_U6 (.B( u0_K4_4 ) , .A( u0_R2_3 ) , .Z( u0_u3_X_4 ) );
  AND2_X1 u0_u3_u0_U10 (.A1( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n143 ) , .A2( u0_u3_u0_n152 ) );
  AND2_X1 u0_u3_u0_U11 (.ZN( u0_u3_u0_n109 ) , .A1( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n142 ) );
  AND2_X1 u0_u3_u0_U12 (.A2( u0_u3_u0_n131 ) , .A1( u0_u3_u0_n132 ) , .ZN( u0_u3_u0_n153 ) );
  AND2_X1 u0_u3_u0_U13 (.A1( u0_u3_u0_n110 ) , .A2( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U14 (.A( u0_u3_u0_n145 ) , .ZN( u0_u3_u0_n175 ) );
  NOR2_X1 u0_u3_u0_U15 (.A2( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n149 ) , .A1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U16 (.B1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n134 ) , .A( u0_u3_u0_n167 ) , .B2( u0_u3_u0_n95 ) );
  OAI22_X1 u0_u3_u0_U17 (.B1( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n149 ) , .A2( u0_u3_u0_n92 ) , .ZN( u0_u3_u0_n93 ) );
  AND3_X1 u0_u3_u0_U18 (.A3( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n127 ) , .A1( u0_u3_u0_n150 ) , .ZN( u0_u3_u0_n92 ) );
  OAI22_X1 u0_u3_u0_U19 (.B1( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n128 ) , .A1( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n148 ) , .B2( u0_u3_u0_n149 ) );
  NOR2_X1 u0_u3_u0_U20 (.A1( u0_u3_u0_n165 ) , .A2( u0_u3_u0_n166 ) , .ZN( u0_u3_u0_n97 ) );
  AOI22_X1 u0_u3_u0_U21 (.B2( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n112 ) , .ZN( u0_u3_u0_n113 ) , .B1( u0_u3_u0_n120 ) , .A1( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U22 (.A2( u0_u3_u0_n104 ) , .A1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n151 ) );
  INV_X1 u0_u3_u0_U23 (.A( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U24 (.A( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n160 ) );
  NAND2_X1 u0_u3_u0_U25 (.A2( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n94 ) );
  NAND2_X1 u0_u3_u0_U26 (.ZN( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n94 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U27 (.ZN( u0_u3_u0_n106 ) , .B1( u0_u3_u0_n109 ) , .B2( u0_u3_u0_n143 ) , .A( u0_u3_u0_n146 ) );
  AOI21_X1 u0_u3_u0_U28 (.B1( u0_u3_u0_n129 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n98 ) );
  NAND2_X1 u0_u3_u0_U29 (.A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n116 ) , .A1( u0_u3_u0_n94 ) );
  INV_X1 u0_u3_u0_U3 (.A( u0_u3_u0_n115 ) , .ZN( u0_u3_u0_n168 ) );
  NOR2_X1 u0_u3_u0_U30 (.A1( u0_u3_u0_n122 ) , .ZN( u0_u3_u0_n145 ) , .A2( u0_u3_u0_n169 ) );
  OAI221_X1 u0_u3_u0_U31 (.C1( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n122 ) , .B1( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n143 ) , .C2( u0_u3_u0_n149 ) , .A( u0_u3_u0_n174 ) );
  AOI211_X1 u0_u3_u0_U32 (.B( u0_u3_u0_n117 ) , .A( u0_u3_u0_n118 ) , .C2( u0_u3_u0_n119 ) , .C1( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n121 ) );
  NAND2_X1 u0_u3_u0_U33 (.A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n96 ) );
  NAND2_X1 u0_u3_u0_U34 (.A1( u0_u3_u0_n102 ) , .A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n127 ) );
  NAND2_X1 u0_u3_u0_U35 (.A1( u0_u3_u0_n103 ) , .A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n152 ) );
  INV_X1 u0_u3_u0_U36 (.A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U37 (.A2( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n141 ) );
  NAND2_X1 u0_u3_u0_U38 (.ZN( u0_u3_u0_n114 ) , .A2( u0_u3_u0_n94 ) , .A1( u0_u3_u0_n95 ) );
  NAND2_X1 u0_u3_u0_U39 (.A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U4 (.B1( u0_u3_u0_n116 ) , .ZN( u0_u3_u0_n117 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U40 (.ZN( u0_u3_u0_n174 ) , .A( u0_u3_u0_n90 ) );
  OAI222_X1 u0_u3_u0_U41 (.C1( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n127 ) , .B2( u0_u3_u0_n130 ) , .B1( u0_u3_u0_n146 ) , .A2( u0_u3_u0_n160 ) , .C2( u0_u3_u0_n163 ) , .ZN( u0_u3_u0_n90 ) );
  OR3_X1 u0_u3_u0_U42 (.A3( u0_u3_u0_n154 ) , .A2( u0_u3_u0_n155 ) , .A1( u0_u3_u0_n156 ) , .ZN( u0_u3_u0_n157 ) );
  AOI21_X1 u0_u3_u0_U43 (.A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n147 ) , .B1( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n156 ) );
  AOI21_X1 u0_u3_u0_U44 (.B2( u0_u3_u0_n152 ) , .B1( u0_u3_u0_n153 ) , .ZN( u0_u3_u0_n154 ) , .A( u0_u3_u0_n160 ) );
  AOI21_X1 u0_u3_u0_U45 (.A( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n150 ) , .B1( u0_u3_u0_n151 ) , .ZN( u0_u3_u0_n155 ) );
  INV_X1 u0_u3_u0_U46 (.A( u0_u3_u0_n101 ) , .ZN( u0_u3_u0_n173 ) );
  OAI211_X1 u0_u3_u0_U47 (.B( u0_u3_u0_n100 ) , .ZN( u0_u3_u0_n101 ) , .C2( u0_u3_u0_n142 ) , .C1( u0_u3_u0_n163 ) , .A( u0_u3_u0_n171 ) );
  INV_X1 u0_u3_u0_U48 (.ZN( u0_u3_u0_n171 ) , .A( u0_u3_u0_n93 ) );
  AOI211_X1 u0_u3_u0_U49 (.ZN( u0_u3_u0_n100 ) , .C1( u0_u3_u0_n120 ) , .A( u0_u3_u0_n125 ) , .B( u0_u3_u0_n98 ) , .C2( u0_u3_u0_n99 ) );
  AOI21_X1 u0_u3_u0_U5 (.B2( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n136 ) , .B1( u0_u3_u0_n153 ) , .A( u0_u3_u0_n160 ) );
  NOR2_X1 u0_u3_u0_U50 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n120 ) );
  NOR2_X1 u0_u3_u0_U51 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n96 ) );
  NOR2_X1 u0_u3_u0_U52 (.A2( u0_u3_X_6 ) , .ZN( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n164 ) );
  NOR2_X1 u0_u3_u0_U53 (.A2( u0_u3_X_1 ) , .ZN( u0_u3_u0_n103 ) , .A1( u0_u3_u0_n165 ) );
  NAND2_X1 u0_u3_u0_U54 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n146 ) );
  NOR2_X1 u0_u3_u0_U55 (.A2( u0_u3_X_5 ) , .ZN( u0_u3_u0_n138 ) , .A1( u0_u3_u0_n161 ) );
  NAND2_X1 u0_u3_u0_U56 (.A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n161 ) );
  AND2_X1 u0_u3_u0_U57 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n104 ) );
  AND2_X1 u0_u3_u0_U58 (.A1( u0_u3_X_6 ) , .A2( u0_u3_u0_n164 ) , .ZN( u0_u3_u0_n95 ) );
  INV_X1 u0_u3_u0_U59 (.A( u0_u3_X_4 ) , .ZN( u0_u3_u0_n161 ) );
  NOR2_X1 u0_u3_u0_U6 (.A1( u0_u3_u0_n110 ) , .ZN( u0_u3_u0_n125 ) , .A2( u0_u3_u0_n160 ) );
  INV_X1 u0_u3_u0_U60 (.A( u0_u3_X_1 ) , .ZN( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U61 (.A( u0_u3_X_3 ) , .ZN( u0_u3_u0_n164 ) );
  INV_X1 u0_u3_u0_U62 (.A( u0_u3_u0_n128 ) , .ZN( u0_u3_u0_n170 ) );
  AOI211_X1 u0_u3_u0_U63 (.B( u0_u3_u0_n135 ) , .A( u0_u3_u0_n136 ) , .C2( u0_u3_u0_n137 ) , .C1( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n139 ) );
  OR4_X1 u0_u3_u0_U64 (.ZN( u0_out3_31 ) , .A4( u0_u3_u0_n157 ) , .A2( u0_u3_u0_n158 ) , .A1( u0_u3_u0_n159 ) , .A3( u0_u3_u0_n175 ) );
  AOI21_X1 u0_u3_u0_U65 (.A( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n141 ) , .B1( u0_u3_u0_n142 ) , .ZN( u0_u3_u0_n159 ) );
  OR4_X1 u0_u3_u0_U66 (.ZN( u0_out3_17 ) , .A4( u0_u3_u0_n124 ) , .A2( u0_u3_u0_n125 ) , .A1( u0_u3_u0_n126 ) , .A3( u0_u3_u0_n172 ) );
  AOI21_X1 u0_u3_u0_U67 (.B2( u0_u3_u0_n109 ) , .ZN( u0_u3_u0_n126 ) , .B1( u0_u3_u0_n130 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U68 (.A( u0_u3_u0_n113 ) , .ZN( u0_u3_u0_n172 ) );
  INV_X1 u0_u3_u0_U69 (.ZN( u0_u3_u0_n176 ) , .A( u0_u3_u0_n91 ) );
  OAI21_X1 u0_u3_u0_U7 (.B1( u0_u3_u0_n152 ) , .B2( u0_u3_u0_n160 ) , .A( u0_u3_u0_n174 ) , .ZN( u0_u3_u0_n91 ) );
  AOI211_X1 u0_u3_u0_U70 (.B( u0_u3_u0_n106 ) , .A( u0_u3_u0_n107 ) , .ZN( u0_u3_u0_n108 ) , .C2( u0_u3_u0_n115 ) , .C1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U71 (.B2( u0_u3_u0_n143 ) , .B1( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n158 ) , .A( u0_u3_u0_n163 ) );
  AOI21_X1 u0_u3_u0_U72 (.ZN( u0_u3_u0_n118 ) , .B2( u0_u3_u0_n144 ) , .A( u0_u3_u0_n146 ) , .B1( u0_u3_u0_n168 ) );
  INV_X1 u0_u3_u0_U73 (.A( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n167 ) );
  NOR2_X1 u0_u3_u0_U74 (.A2( u0_u3_X_1 ) , .A1( u0_u3_X_2 ) , .ZN( u0_u3_u0_n94 ) );
  NOR2_X1 u0_u3_u0_U75 (.A2( u0_u3_X_2 ) , .ZN( u0_u3_u0_n105 ) , .A1( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U76 (.A( u0_u3_X_2 ) , .ZN( u0_u3_u0_n165 ) );
  OR2_X1 u0_u3_u0_U77 (.A2( u0_u3_u0_n129 ) , .A1( u0_u3_u0_n146 ) , .ZN( u0_u3_u0_n88 ) );
  OR2_X1 u0_u3_u0_U78 (.A1( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n149 ) , .ZN( u0_u3_u0_n89 ) );
  NAND3_X1 u0_u3_u0_U79 (.ZN( u0_u3_u0_n124 ) , .A3( u0_u3_u0_n145 ) , .A1( u0_u3_u0_n88 ) , .A2( u0_u3_u0_n89 ) );
  AND2_X1 u0_u3_u0_U8 (.A1( u0_u3_u0_n116 ) , .A2( u0_u3_u0_n123 ) , .ZN( u0_u3_u0_n148 ) );
  AND3_X1 u0_u3_u0_U80 (.A2( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n129 ) , .A3( u0_u3_u0_n132 ) , .A1( u0_u3_u0_n150 ) );
  NAND2_X1 u0_u3_u0_U81 (.A2( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n123 ) , .A1( u0_u3_u0_n95 ) );
  AOI21_X1 u0_u3_u0_U82 (.B1( u0_u3_u0_n134 ) , .ZN( u0_u3_u0_n135 ) , .A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n168 ) );
  OAI22_X1 u0_u3_u0_U83 (.ZN( u0_u3_u0_n107 ) , .A2( u0_u3_u0_n134 ) , .B1( u0_u3_u0_n148 ) , .A1( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n163 ) );
  NAND2_X1 u0_u3_u0_U84 (.ZN( u0_u3_u0_n112 ) , .A2( u0_u3_u0_n134 ) , .A1( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U85 (.A( u0_u3_u0_n121 ) , .ZN( u0_u3_u0_n169 ) );
  NAND2_X1 u0_u3_u0_U86 (.ZN( u0_u3_u0_n150 ) , .A1( u0_u3_u0_n95 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U87 (.A1( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n131 ) , .A2( u0_u3_u0_n97 ) );
  NAND3_X1 u0_u3_u0_U88 (.ZN( u0_out3_23 ) , .A3( u0_u3_u0_n139 ) , .A1( u0_u3_u0_n170 ) , .A2( u0_u3_u0_n173 ) );
  NAND3_X1 u0_u3_u0_U89 (.A3( u0_u3_u0_n129 ) , .A2( u0_u3_u0_n130 ) , .ZN( u0_u3_u0_n137 ) , .A1( u0_u3_u0_n152 ) );
  NAND2_X1 u0_u3_u0_U9 (.ZN( u0_u3_u0_n115 ) , .A1( u0_u3_u0_n141 ) , .A2( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U90 (.ZN( u0_u3_u0_n119 ) , .A3( u0_u3_u0_n134 ) , .A2( u0_u3_u0_n141 ) , .A1( u0_u3_u0_n150 ) );
  NAND3_X1 u0_u3_u0_U91 (.ZN( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n116 ) , .A3( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U92 (.ZN( u0_out3_9 ) , .A3( u0_u3_u0_n108 ) , .A2( u0_u3_u0_n173 ) , .A1( u0_u3_u0_n176 ) );
  NAND3_X1 u0_u3_u0_U93 (.A2( u0_u3_u0_n130 ) , .A1( u0_u3_u0_n134 ) , .A3( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n99 ) );
  NAND2_X1 u0_u3_u0_U94 (.A1( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n130 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U95 (.ZN( u0_u3_u0_n144 ) , .A1( u0_u3_u0_n96 ) , .A2( u0_u3_u0_n97 ) );
  NOR2_X1 u0_u3_u1_U10 (.A1( u0_u3_u1_n112 ) , .A2( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n118 ) );
  NAND3_X1 u0_u3_u1_U100 (.ZN( u0_u3_u1_n113 ) , .A1( u0_u3_u1_n120 ) , .A3( u0_u3_u1_n133 ) , .A2( u0_u3_u1_n155 ) );
  OAI21_X1 u0_u3_u1_U11 (.ZN( u0_u3_u1_n101 ) , .B1( u0_u3_u1_n141 ) , .A( u0_u3_u1_n146 ) , .B2( u0_u3_u1_n183 ) );
  AOI21_X1 u0_u3_u1_U12 (.B2( u0_u3_u1_n155 ) , .B1( u0_u3_u1_n156 ) , .ZN( u0_u3_u1_n157 ) , .A( u0_u3_u1_n174 ) );
  NAND2_X1 u0_u3_u1_U13 (.ZN( u0_u3_u1_n140 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n155 ) );
  NAND2_X1 u0_u3_u1_U14 (.A1( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n153 ) );
  INV_X1 u0_u3_u1_U15 (.A( u0_u3_u1_n139 ) , .ZN( u0_u3_u1_n174 ) );
  OR4_X1 u0_u3_u1_U16 (.A4( u0_u3_u1_n106 ) , .A3( u0_u3_u1_n107 ) , .ZN( u0_u3_u1_n108 ) , .A1( u0_u3_u1_n117 ) , .A2( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U17 (.ZN( u0_u3_u1_n106 ) , .A( u0_u3_u1_n112 ) , .B1( u0_u3_u1_n154 ) , .B2( u0_u3_u1_n156 ) );
  INV_X1 u0_u3_u1_U18 (.A( u0_u3_u1_n101 ) , .ZN( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U19 (.ZN( u0_u3_u1_n107 ) , .B1( u0_u3_u1_n134 ) , .B2( u0_u3_u1_n149 ) , .A( u0_u3_u1_n174 ) );
  INV_X1 u0_u3_u1_U20 (.A( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n171 ) );
  NAND2_X1 u0_u3_u1_U21 (.ZN( u0_u3_u1_n141 ) , .A1( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n156 ) );
  AND2_X1 u0_u3_u1_U22 (.A1( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n161 ) );
  NAND2_X1 u0_u3_u1_U23 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n148 ) );
  NAND2_X1 u0_u3_u1_U24 (.A2( u0_u3_u1_n133 ) , .A1( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n159 ) );
  NAND2_X1 u0_u3_u1_U25 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n120 ) , .ZN( u0_u3_u1_n132 ) );
  INV_X1 u0_u3_u1_U26 (.A( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n178 ) );
  INV_X1 u0_u3_u1_U27 (.A( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n183 ) );
  AND2_X1 u0_u3_u1_U28 (.A1( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n149 ) );
  INV_X1 u0_u3_u1_U29 (.A( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n180 ) );
  INV_X1 u0_u3_u1_U3 (.A( u0_u3_u1_n159 ) , .ZN( u0_u3_u1_n182 ) );
  AOI221_X1 u0_u3_u1_U30 (.B1( u0_u3_u1_n140 ) , .ZN( u0_u3_u1_n167 ) , .B2( u0_u3_u1_n172 ) , .C2( u0_u3_u1_n175 ) , .C1( u0_u3_u1_n178 ) , .A( u0_u3_u1_n188 ) );
  INV_X1 u0_u3_u1_U31 (.ZN( u0_u3_u1_n188 ) , .A( u0_u3_u1_n97 ) );
  AOI211_X1 u0_u3_u1_U32 (.A( u0_u3_u1_n118 ) , .C1( u0_u3_u1_n132 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n96 ) , .ZN( u0_u3_u1_n97 ) );
  AOI21_X1 u0_u3_u1_U33 (.B2( u0_u3_u1_n121 ) , .B1( u0_u3_u1_n135 ) , .A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n96 ) );
  OAI221_X1 u0_u3_u1_U34 (.A( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n138 ) , .B2( u0_u3_u1_n152 ) , .C1( u0_u3_u1_n174 ) , .B1( u0_u3_u1_n187 ) );
  INV_X1 u0_u3_u1_U35 (.A( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n187 ) );
  AOI211_X1 u0_u3_u1_U36 (.B( u0_u3_u1_n117 ) , .A( u0_u3_u1_n118 ) , .ZN( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n146 ) , .C1( u0_u3_u1_n159 ) );
  NOR2_X1 u0_u3_u1_U37 (.A1( u0_u3_u1_n168 ) , .A2( u0_u3_u1_n176 ) , .ZN( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U38 (.A1( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n146 ) , .A2( u0_u3_u1_n160 ) );
  NAND2_X1 u0_u3_u1_U39 (.A2( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n139 ) , .A1( u0_u3_u1_n152 ) );
  AOI221_X1 u0_u3_u1_U4 (.A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .C1( u0_u3_u1_n140 ) , .B2( u0_u3_u1_n141 ) , .ZN( u0_u3_u1_n142 ) , .B1( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U40 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n156 ) , .A2( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U41 (.ZN( u0_u3_u1_n117 ) , .A1( u0_u3_u1_n121 ) , .A2( u0_u3_u1_n160 ) );
  OAI21_X1 u0_u3_u1_U42 (.B2( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n145 ) , .B1( u0_u3_u1_n160 ) , .A( u0_u3_u1_n185 ) );
  INV_X1 u0_u3_u1_U43 (.A( u0_u3_u1_n122 ) , .ZN( u0_u3_u1_n185 ) );
  AOI21_X1 u0_u3_u1_U44 (.B2( u0_u3_u1_n120 ) , .B1( u0_u3_u1_n121 ) , .ZN( u0_u3_u1_n122 ) , .A( u0_u3_u1_n128 ) );
  AOI21_X1 u0_u3_u1_U45 (.A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n130 ) , .B1( u0_u3_u1_n150 ) );
  NAND2_X1 u0_u3_u1_U46 (.ZN( u0_u3_u1_n112 ) , .A1( u0_u3_u1_n169 ) , .A2( u0_u3_u1_n170 ) );
  NAND2_X1 u0_u3_u1_U47 (.ZN( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n95 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U48 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n154 ) , .A2( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U49 (.A2( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n135 ) , .A1( u0_u3_u1_n99 ) );
  AOI211_X1 u0_u3_u1_U5 (.ZN( u0_u3_u1_n124 ) , .A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n145 ) , .C1( u0_u3_u1_n147 ) );
  AOI21_X1 u0_u3_u1_U50 (.A( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n153 ) , .B1( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n158 ) );
  INV_X1 u0_u3_u1_U51 (.A( u0_u3_u1_n160 ) , .ZN( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U52 (.A1( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n116 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U53 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n131 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U54 (.A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n121 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U55 (.A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U56 (.A2( u0_u3_u1_n104 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n133 ) );
  NAND2_X1 u0_u3_u1_U57 (.ZN( u0_u3_u1_n150 ) , .A2( u0_u3_u1_n98 ) , .A1( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U58 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n155 ) , .A2( u0_u3_u1_n95 ) );
  OAI21_X1 u0_u3_u1_U59 (.ZN( u0_u3_u1_n109 ) , .B1( u0_u3_u1_n129 ) , .B2( u0_u3_u1_n160 ) , .A( u0_u3_u1_n167 ) );
  AOI22_X1 u0_u3_u1_U6 (.B2( u0_u3_u1_n113 ) , .A2( u0_u3_u1_n114 ) , .ZN( u0_u3_u1_n125 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  NAND2_X1 u0_u3_u1_U60 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n120 ) );
  NAND2_X1 u0_u3_u1_U61 (.A1( u0_u3_u1_n102 ) , .A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n115 ) );
  NAND2_X1 u0_u3_u1_U62 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n151 ) );
  NAND2_X1 u0_u3_u1_U63 (.A2( u0_u3_u1_n103 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n161 ) );
  INV_X1 u0_u3_u1_U64 (.A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U65 (.A( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n172 ) );
  NAND2_X1 u0_u3_u1_U66 (.A2( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n123 ) );
  AOI211_X1 u0_u3_u1_U67 (.B( u0_u3_u1_n162 ) , .A( u0_u3_u1_n163 ) , .C2( u0_u3_u1_n164 ) , .ZN( u0_u3_u1_n165 ) , .C1( u0_u3_u1_n171 ) );
  AOI21_X1 u0_u3_u1_U68 (.A( u0_u3_u1_n160 ) , .B2( u0_u3_u1_n161 ) , .ZN( u0_u3_u1_n162 ) , .B1( u0_u3_u1_n182 ) );
  OR2_X1 u0_u3_u1_U69 (.A2( u0_u3_u1_n157 ) , .A1( u0_u3_u1_n158 ) , .ZN( u0_u3_u1_n163 ) );
  NAND2_X1 u0_u3_u1_U7 (.ZN( u0_u3_u1_n114 ) , .A1( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n156 ) );
  NOR2_X1 u0_u3_u1_U70 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n95 ) );
  NOR2_X1 u0_u3_u1_U71 (.A1( u0_u3_X_12 ) , .A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n100 ) );
  NOR2_X1 u0_u3_u1_U72 (.A2( u0_u3_X_8 ) , .A1( u0_u3_u1_n177 ) , .ZN( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U73 (.A2( u0_u3_X_12 ) , .ZN( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n176 ) );
  NOR2_X1 u0_u3_u1_U74 (.A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n105 ) , .A1( u0_u3_u1_n168 ) );
  NAND2_X1 u0_u3_u1_U75 (.A1( u0_u3_X_10 ) , .ZN( u0_u3_u1_n160 ) , .A2( u0_u3_u1_n169 ) );
  NAND2_X1 u0_u3_u1_U76 (.A2( u0_u3_X_10 ) , .A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n152 ) );
  NAND2_X1 u0_u3_u1_U77 (.A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n128 ) , .A2( u0_u3_u1_n170 ) );
  AND2_X1 u0_u3_u1_U78 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n104 ) );
  AND2_X1 u0_u3_u1_U79 (.A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n103 ) , .A2( u0_u3_u1_n177 ) );
  AOI22_X1 u0_u3_u1_U8 (.B2( u0_u3_u1_n136 ) , .A2( u0_u3_u1_n137 ) , .ZN( u0_u3_u1_n143 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U80 (.A( u0_u3_X_10 ) , .ZN( u0_u3_u1_n170 ) );
  INV_X1 u0_u3_u1_U81 (.A( u0_u3_X_9 ) , .ZN( u0_u3_u1_n176 ) );
  INV_X1 u0_u3_u1_U82 (.A( u0_u3_X_11 ) , .ZN( u0_u3_u1_n169 ) );
  INV_X1 u0_u3_u1_U83 (.A( u0_u3_X_12 ) , .ZN( u0_u3_u1_n168 ) );
  INV_X1 u0_u3_u1_U84 (.A( u0_u3_X_7 ) , .ZN( u0_u3_u1_n177 ) );
  NAND4_X1 u0_u3_u1_U85 (.ZN( u0_out3_28 ) , .A4( u0_u3_u1_n124 ) , .A3( u0_u3_u1_n125 ) , .A2( u0_u3_u1_n126 ) , .A1( u0_u3_u1_n127 ) );
  OAI21_X1 u0_u3_u1_U86 (.ZN( u0_u3_u1_n127 ) , .B2( u0_u3_u1_n139 ) , .B1( u0_u3_u1_n175 ) , .A( u0_u3_u1_n183 ) );
  OAI21_X1 u0_u3_u1_U87 (.ZN( u0_u3_u1_n126 ) , .B2( u0_u3_u1_n140 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n178 ) );
  NAND4_X1 u0_u3_u1_U88 (.ZN( u0_out3_18 ) , .A4( u0_u3_u1_n165 ) , .A3( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n167 ) , .A2( u0_u3_u1_n186 ) );
  AOI22_X1 u0_u3_u1_U89 (.B2( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n172 ) );
  INV_X1 u0_u3_u1_U9 (.A( u0_u3_u1_n147 ) , .ZN( u0_u3_u1_n181 ) );
  INV_X1 u0_u3_u1_U90 (.A( u0_u3_u1_n145 ) , .ZN( u0_u3_u1_n186 ) );
  NAND4_X1 u0_u3_u1_U91 (.ZN( u0_out3_2 ) , .A4( u0_u3_u1_n142 ) , .A3( u0_u3_u1_n143 ) , .A2( u0_u3_u1_n144 ) , .A1( u0_u3_u1_n179 ) );
  INV_X1 u0_u3_u1_U92 (.A( u0_u3_u1_n130 ) , .ZN( u0_u3_u1_n179 ) );
  OAI21_X1 u0_u3_u1_U93 (.B2( u0_u3_u1_n132 ) , .ZN( u0_u3_u1_n144 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n180 ) );
  OR4_X1 u0_u3_u1_U94 (.ZN( u0_out3_13 ) , .A4( u0_u3_u1_n108 ) , .A3( u0_u3_u1_n109 ) , .A2( u0_u3_u1_n110 ) , .A1( u0_u3_u1_n111 ) );
  AOI21_X1 u0_u3_u1_U95 (.ZN( u0_u3_u1_n111 ) , .A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n131 ) , .B1( u0_u3_u1_n135 ) );
  AOI21_X1 u0_u3_u1_U96 (.ZN( u0_u3_u1_n110 ) , .A( u0_u3_u1_n116 ) , .B1( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n160 ) );
  NAND3_X1 u0_u3_u1_U97 (.A3( u0_u3_u1_n149 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n164 ) );
  NAND3_X1 u0_u3_u1_U98 (.A3( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n136 ) , .A1( u0_u3_u1_n151 ) );
  NAND3_X1 u0_u3_u1_U99 (.A1( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n137 ) , .A2( u0_u3_u1_n154 ) , .A3( u0_u3_u1_n181 ) );
  OAI22_X1 u0_u3_u2_U10 (.B1( u0_u3_u2_n151 ) , .A2( u0_u3_u2_n152 ) , .A1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n160 ) , .B2( u0_u3_u2_n168 ) );
  NAND3_X1 u0_u3_u2_U100 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n98 ) );
  NOR3_X1 u0_u3_u2_U11 (.A1( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n151 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U12 (.B2( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n125 ) , .A( u0_u3_u2_n171 ) , .B1( u0_u3_u2_n184 ) );
  INV_X1 u0_u3_u2_U13 (.A( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n184 ) );
  AOI21_X1 u0_u3_u2_U14 (.ZN( u0_u3_u2_n144 ) , .B2( u0_u3_u2_n155 ) , .A( u0_u3_u2_n172 ) , .B1( u0_u3_u2_n185 ) );
  AOI21_X1 u0_u3_u2_U15 (.B2( u0_u3_u2_n143 ) , .ZN( u0_u3_u2_n145 ) , .B1( u0_u3_u2_n152 ) , .A( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U16 (.A( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U17 (.A( u0_u3_u2_n120 ) , .ZN( u0_u3_u2_n188 ) );
  NAND2_X1 u0_u3_u2_U18 (.A2( u0_u3_u2_n122 ) , .ZN( u0_u3_u2_n150 ) , .A1( u0_u3_u2_n152 ) );
  INV_X1 u0_u3_u2_U19 (.A( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n170 ) );
  INV_X1 u0_u3_u2_U20 (.A( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n173 ) );
  NAND2_X1 u0_u3_u2_U21 (.A1( u0_u3_u2_n132 ) , .A2( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n157 ) );
  INV_X1 u0_u3_u2_U22 (.A( u0_u3_u2_n113 ) , .ZN( u0_u3_u2_n178 ) );
  INV_X1 u0_u3_u2_U23 (.A( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n175 ) );
  INV_X1 u0_u3_u2_U24 (.A( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n181 ) );
  INV_X1 u0_u3_u2_U25 (.A( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n177 ) );
  INV_X1 u0_u3_u2_U26 (.A( u0_u3_u2_n116 ) , .ZN( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U27 (.A( u0_u3_u2_n131 ) , .ZN( u0_u3_u2_n179 ) );
  INV_X1 u0_u3_u2_U28 (.A( u0_u3_u2_n154 ) , .ZN( u0_u3_u2_n176 ) );
  NAND2_X1 u0_u3_u2_U29 (.A2( u0_u3_u2_n116 ) , .A1( u0_u3_u2_n117 ) , .ZN( u0_u3_u2_n118 ) );
  NOR2_X1 u0_u3_u2_U3 (.ZN( u0_u3_u2_n121 ) , .A2( u0_u3_u2_n177 ) , .A1( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U30 (.A( u0_u3_u2_n132 ) , .ZN( u0_u3_u2_n182 ) );
  INV_X1 u0_u3_u2_U31 (.A( u0_u3_u2_n158 ) , .ZN( u0_u3_u2_n183 ) );
  OAI21_X1 u0_u3_u2_U32 (.A( u0_u3_u2_n156 ) , .B1( u0_u3_u2_n157 ) , .ZN( u0_u3_u2_n158 ) , .B2( u0_u3_u2_n179 ) );
  NOR2_X1 u0_u3_u2_U33 (.ZN( u0_u3_u2_n156 ) , .A1( u0_u3_u2_n166 ) , .A2( u0_u3_u2_n169 ) );
  NOR2_X1 u0_u3_u2_U34 (.A2( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n140 ) );
  NOR2_X1 u0_u3_u2_U35 (.A2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n153 ) , .A1( u0_u3_u2_n156 ) );
  AOI211_X1 u0_u3_u2_U36 (.ZN( u0_u3_u2_n130 ) , .C1( u0_u3_u2_n138 ) , .C2( u0_u3_u2_n179 ) , .B( u0_u3_u2_n96 ) , .A( u0_u3_u2_n97 ) );
  OAI22_X1 u0_u3_u2_U37 (.B1( u0_u3_u2_n133 ) , .A2( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n152 ) , .B2( u0_u3_u2_n168 ) , .ZN( u0_u3_u2_n97 ) );
  OAI221_X1 u0_u3_u2_U38 (.B1( u0_u3_u2_n113 ) , .C1( u0_u3_u2_n132 ) , .A( u0_u3_u2_n149 ) , .B2( u0_u3_u2_n171 ) , .C2( u0_u3_u2_n172 ) , .ZN( u0_u3_u2_n96 ) );
  OAI221_X1 u0_u3_u2_U39 (.A( u0_u3_u2_n115 ) , .C2( u0_u3_u2_n123 ) , .B2( u0_u3_u2_n143 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n163 ) , .C1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U4 (.A( u0_u3_u2_n134 ) , .ZN( u0_u3_u2_n185 ) );
  OAI21_X1 u0_u3_u2_U40 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n115 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n178 ) );
  OAI221_X1 u0_u3_u2_U41 (.A( u0_u3_u2_n135 ) , .B2( u0_u3_u2_n136 ) , .B1( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n162 ) , .C2( u0_u3_u2_n167 ) , .C1( u0_u3_u2_n185 ) );
  AND3_X1 u0_u3_u2_U42 (.A3( u0_u3_u2_n131 ) , .A2( u0_u3_u2_n132 ) , .A1( u0_u3_u2_n133 ) , .ZN( u0_u3_u2_n136 ) );
  AOI22_X1 u0_u3_u2_U43 (.ZN( u0_u3_u2_n135 ) , .B1( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n156 ) , .B2( u0_u3_u2_n180 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U44 (.ZN( u0_u3_u2_n149 ) , .B1( u0_u3_u2_n173 ) , .B2( u0_u3_u2_n188 ) , .A( u0_u3_u2_n95 ) );
  AND3_X1 u0_u3_u2_U45 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n95 ) );
  OAI21_X1 u0_u3_u2_U46 (.A( u0_u3_u2_n141 ) , .B2( u0_u3_u2_n142 ) , .ZN( u0_u3_u2_n146 ) , .B1( u0_u3_u2_n153 ) );
  OAI21_X1 u0_u3_u2_U47 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n141 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n177 ) );
  NOR3_X1 u0_u3_u2_U48 (.ZN( u0_u3_u2_n142 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n178 ) , .A1( u0_u3_u2_n181 ) );
  OAI21_X1 u0_u3_u2_U49 (.A( u0_u3_u2_n101 ) , .B2( u0_u3_u2_n121 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n164 ) );
  NOR4_X1 u0_u3_u2_U5 (.A4( u0_u3_u2_n124 ) , .A3( u0_u3_u2_n125 ) , .A2( u0_u3_u2_n126 ) , .A1( u0_u3_u2_n127 ) , .ZN( u0_u3_u2_n128 ) );
  NAND2_X1 u0_u3_u2_U50 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U51 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n143 ) );
  NAND2_X1 u0_u3_u2_U52 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n152 ) );
  NAND2_X1 u0_u3_u2_U53 (.A1( u0_u3_u2_n100 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n132 ) );
  INV_X1 u0_u3_u2_U54 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U55 (.A( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n167 ) );
  INV_X1 u0_u3_u2_U56 (.ZN( u0_u3_u2_n187 ) , .A( u0_u3_u2_n99 ) );
  OAI21_X1 u0_u3_u2_U57 (.B1( u0_u3_u2_n137 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n98 ) , .ZN( u0_u3_u2_n99 ) );
  NAND2_X1 u0_u3_u2_U58 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n113 ) );
  NAND2_X1 u0_u3_u2_U59 (.A1( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n131 ) );
  AOI21_X1 u0_u3_u2_U6 (.B2( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n127 ) , .A( u0_u3_u2_n137 ) , .B1( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U60 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n139 ) );
  NAND2_X1 u0_u3_u2_U61 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n133 ) );
  NAND2_X1 u0_u3_u2_U62 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n103 ) , .ZN( u0_u3_u2_n154 ) );
  NAND2_X1 u0_u3_u2_U63 (.A2( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n104 ) , .ZN( u0_u3_u2_n119 ) );
  NAND2_X1 u0_u3_u2_U64 (.A2( u0_u3_u2_n107 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n123 ) );
  NAND2_X1 u0_u3_u2_U65 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n122 ) );
  INV_X1 u0_u3_u2_U66 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n172 ) );
  NAND2_X1 u0_u3_u2_U67 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n102 ) , .ZN( u0_u3_u2_n116 ) );
  NAND2_X1 u0_u3_u2_U68 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n120 ) );
  NAND2_X1 u0_u3_u2_U69 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n117 ) );
  AOI21_X1 u0_u3_u2_U7 (.ZN( u0_u3_u2_n124 ) , .B1( u0_u3_u2_n131 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n172 ) );
  NOR2_X1 u0_u3_u2_U70 (.A2( u0_u3_X_16 ) , .ZN( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n166 ) );
  NOR2_X1 u0_u3_u2_U71 (.A2( u0_u3_X_13 ) , .A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n100 ) );
  NOR2_X1 u0_u3_u2_U72 (.A2( u0_u3_X_16 ) , .A1( u0_u3_X_17 ) , .ZN( u0_u3_u2_n138 ) );
  NOR2_X1 u0_u3_u2_U73 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n104 ) );
  NOR2_X1 u0_u3_u2_U74 (.A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n174 ) );
  NOR2_X1 u0_u3_u2_U75 (.A2( u0_u3_X_15 ) , .ZN( u0_u3_u2_n102 ) , .A1( u0_u3_u2_n165 ) );
  NOR2_X1 u0_u3_u2_U76 (.A2( u0_u3_X_17 ) , .ZN( u0_u3_u2_n114 ) , .A1( u0_u3_u2_n169 ) );
  AND2_X1 u0_u3_u2_U77 (.A1( u0_u3_X_15 ) , .ZN( u0_u3_u2_n105 ) , .A2( u0_u3_u2_n165 ) );
  AND2_X1 u0_u3_u2_U78 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n107 ) );
  AND2_X1 u0_u3_u2_U79 (.A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n174 ) );
  AOI21_X1 u0_u3_u2_U8 (.B2( u0_u3_u2_n120 ) , .B1( u0_u3_u2_n121 ) , .ZN( u0_u3_u2_n126 ) , .A( u0_u3_u2_n167 ) );
  AND2_X1 u0_u3_u2_U80 (.A1( u0_u3_X_13 ) , .A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n108 ) );
  INV_X1 u0_u3_u2_U81 (.A( u0_u3_X_16 ) , .ZN( u0_u3_u2_n169 ) );
  INV_X1 u0_u3_u2_U82 (.A( u0_u3_X_17 ) , .ZN( u0_u3_u2_n166 ) );
  INV_X1 u0_u3_u2_U83 (.A( u0_u3_X_13 ) , .ZN( u0_u3_u2_n174 ) );
  INV_X1 u0_u3_u2_U84 (.A( u0_u3_X_18 ) , .ZN( u0_u3_u2_n165 ) );
  NAND4_X1 u0_u3_u2_U85 (.ZN( u0_out3_24 ) , .A4( u0_u3_u2_n111 ) , .A3( u0_u3_u2_n112 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n187 ) );
  AOI221_X1 u0_u3_u2_U86 (.A( u0_u3_u2_n109 ) , .B1( u0_u3_u2_n110 ) , .ZN( u0_u3_u2_n111 ) , .C1( u0_u3_u2_n134 ) , .C2( u0_u3_u2_n170 ) , .B2( u0_u3_u2_n173 ) );
  AOI21_X1 u0_u3_u2_U87 (.ZN( u0_u3_u2_n112 ) , .B2( u0_u3_u2_n156 ) , .A( u0_u3_u2_n164 ) , .B1( u0_u3_u2_n181 ) );
  NAND4_X1 u0_u3_u2_U88 (.ZN( u0_out3_16 ) , .A4( u0_u3_u2_n128 ) , .A3( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n186 ) );
  AOI22_X1 u0_u3_u2_U89 (.A2( u0_u3_u2_n118 ) , .ZN( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n140 ) , .B1( u0_u3_u2_n157 ) , .B2( u0_u3_u2_n170 ) );
  OAI22_X1 u0_u3_u2_U9 (.ZN( u0_u3_u2_n109 ) , .A2( u0_u3_u2_n113 ) , .B2( u0_u3_u2_n133 ) , .B1( u0_u3_u2_n167 ) , .A1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U90 (.A( u0_u3_u2_n163 ) , .ZN( u0_u3_u2_n186 ) );
  NAND4_X1 u0_u3_u2_U91 (.ZN( u0_out3_30 ) , .A4( u0_u3_u2_n147 ) , .A3( u0_u3_u2_n148 ) , .A2( u0_u3_u2_n149 ) , .A1( u0_u3_u2_n187 ) );
  AOI21_X1 u0_u3_u2_U92 (.B2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n148 ) , .A( u0_u3_u2_n162 ) , .B1( u0_u3_u2_n182 ) );
  NOR3_X1 u0_u3_u2_U93 (.A3( u0_u3_u2_n144 ) , .A2( u0_u3_u2_n145 ) , .A1( u0_u3_u2_n146 ) , .ZN( u0_u3_u2_n147 ) );
  OR4_X1 u0_u3_u2_U94 (.ZN( u0_out3_6 ) , .A4( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n162 ) , .A2( u0_u3_u2_n163 ) , .A1( u0_u3_u2_n164 ) );
  OR3_X1 u0_u3_u2_U95 (.A2( u0_u3_u2_n159 ) , .A1( u0_u3_u2_n160 ) , .ZN( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n183 ) );
  AOI21_X1 u0_u3_u2_U96 (.B2( u0_u3_u2_n154 ) , .B1( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n159 ) , .A( u0_u3_u2_n167 ) );
  NAND3_X1 u0_u3_u2_U97 (.A2( u0_u3_u2_n117 ) , .A1( u0_u3_u2_n122 ) , .A3( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n134 ) );
  NAND3_X1 u0_u3_u2_U98 (.ZN( u0_u3_u2_n110 ) , .A2( u0_u3_u2_n131 ) , .A3( u0_u3_u2_n139 ) , .A1( u0_u3_u2_n154 ) );
  NAND3_X1 u0_u3_u2_U99 (.A2( u0_u3_u2_n100 ) , .ZN( u0_u3_u2_n101 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n114 ) );
  OAI22_X1 u0_u3_u3_U10 (.B1( u0_u3_u3_n113 ) , .A2( u0_u3_u3_n135 ) , .A1( u0_u3_u3_n150 ) , .B2( u0_u3_u3_n164 ) , .ZN( u0_u3_u3_n98 ) );
  OAI211_X1 u0_u3_u3_U11 (.B( u0_u3_u3_n106 ) , .ZN( u0_u3_u3_n119 ) , .C2( u0_u3_u3_n128 ) , .C1( u0_u3_u3_n167 ) , .A( u0_u3_u3_n181 ) );
  AOI221_X1 u0_u3_u3_U12 (.C1( u0_u3_u3_n105 ) , .ZN( u0_u3_u3_n106 ) , .A( u0_u3_u3_n131 ) , .B2( u0_u3_u3_n132 ) , .C2( u0_u3_u3_n133 ) , .B1( u0_u3_u3_n169 ) );
  INV_X1 u0_u3_u3_U13 (.ZN( u0_u3_u3_n181 ) , .A( u0_u3_u3_n98 ) );
  NAND2_X1 u0_u3_u3_U14 (.ZN( u0_u3_u3_n105 ) , .A2( u0_u3_u3_n130 ) , .A1( u0_u3_u3_n155 ) );
  AOI22_X1 u0_u3_u3_U15 (.B1( u0_u3_u3_n115 ) , .A2( u0_u3_u3_n116 ) , .ZN( u0_u3_u3_n123 ) , .B2( u0_u3_u3_n133 ) , .A1( u0_u3_u3_n169 ) );
  NAND2_X1 u0_u3_u3_U16 (.ZN( u0_u3_u3_n116 ) , .A2( u0_u3_u3_n151 ) , .A1( u0_u3_u3_n182 ) );
  NOR2_X1 u0_u3_u3_U17 (.ZN( u0_u3_u3_n126 ) , .A2( u0_u3_u3_n150 ) , .A1( u0_u3_u3_n164 ) );
  AOI21_X1 u0_u3_u3_U18 (.ZN( u0_u3_u3_n112 ) , .B2( u0_u3_u3_n146 ) , .B1( u0_u3_u3_n155 ) , .A( u0_u3_u3_n167 ) );
  NAND2_X1 u0_u3_u3_U19 (.A1( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n142 ) , .A2( u0_u3_u3_n164 ) );
  NAND2_X1 u0_u3_u3_U20 (.ZN( u0_u3_u3_n132 ) , .A2( u0_u3_u3_n152 ) , .A1( u0_u3_u3_n156 ) );
  INV_X1 u0_u3_u3_U21 (.A( u0_u3_u3_n133 ) , .ZN( u0_u3_u3_n165 ) );
  NAND2_X1 u0_u3_u3_U22 (.ZN( u0_u3_u3_n143 ) , .A1( u0_u3_u3_n165 ) , .A2( u0_u3_u3_n167 ) );
  AND2_X1 u0_u3_u3_U23 (.A2( u0_u3_u3_n113 ) , .A1( u0_u3_u3_n114 ) , .ZN( u0_u3_u3_n151 ) );
  INV_X1 u0_u3_u3_U24 (.A( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n170 ) );
  NAND2_X1 u0_u3_u3_U25 (.A1( u0_u3_u3_n107 ) , .A2( u0_u3_u3_n108 ) , .ZN( u0_u3_u3_n140 ) );
  NAND2_X1 u0_u3_u3_U26 (.ZN( u0_u3_u3_n117 ) , .A1( u0_u3_u3_n124 ) , .A2( u0_u3_u3_n148 ) );
  INV_X1 u0_u3_u3_U27 (.A( u0_u3_u3_n130 ) , .ZN( u0_u3_u3_n177 ) );
  INV_X1 u0_u3_u3_U28 (.A( u0_u3_u3_n128 ) , .ZN( u0_u3_u3_n176 ) );
  INV_X1 u0_u3_u3_U29 (.A( u0_u3_u3_n155 ) , .ZN( u0_u3_u3_n174 ) );
  INV_X1 u0_u3_u3_U3 (.A( u0_u3_u3_n140 ) , .ZN( u0_u3_u3_n182 ) );
  INV_X1 u0_u3_u3_U30 (.A( u0_u3_u3_n139 ) , .ZN( u0_u3_u3_n185 ) );
  NOR2_X1 u0_u3_u3_U31 (.ZN( u0_u3_u3_n135 ) , .A2( u0_u3_u3_n141 ) , .A1( u0_u3_u3_n169 ) );
  INV_X1 u0_u3_u3_U32 (.A( u0_u3_u3_n156 ) , .ZN( u0_u3_u3_n179 ) );
  OAI22_X1 u0_u3_u3_U33 (.B1( u0_u3_u3_n118 ) , .ZN( u0_u3_u3_n120 ) , .A1( u0_u3_u3_n135 ) , .B2( u0_u3_u3_n154 ) , .A2( u0_u3_u3_n178 ) );
  AND3_X1 u0_u3_u3_U34 (.ZN( u0_u3_u3_n118 ) , .A2( u0_u3_u3_n124 ) , .A1( u0_u3_u3_n144 ) , .A3( u0_u3_u3_n152 ) );
  OAI222_X1 u0_u3_u3_U35 (.C2( u0_u3_u3_n107 ) , .A2( u0_u3_u3_n108 ) , .B1( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n138 ) , .B2( u0_u3_u3_n146 ) , .C1( u0_u3_u3_n154 ) , .A1( u0_u3_u3_n164 ) );
  NOR4_X1 u0_u3_u3_U36 (.A4( u0_u3_u3_n157 ) , .A3( u0_u3_u3_n158 ) , .A2( u0_u3_u3_n159 ) , .A1( u0_u3_u3_n160 ) , .ZN( u0_u3_u3_n161 ) );
  AOI21_X1 u0_u3_u3_U37 (.B2( u0_u3_u3_n152 ) , .B1( u0_u3_u3_n153 ) , .ZN( u0_u3_u3_n158 ) , .A( u0_u3_u3_n164 ) );
  AOI21_X1 u0_u3_u3_U38 (.A( u0_u3_u3_n149 ) , .B2( u0_u3_u3_n150 ) , .B1( u0_u3_u3_n151 ) , .ZN( u0_u3_u3_n159 ) );
  AOI21_X1 u0_u3_u3_U39 (.A( u0_u3_u3_n154 ) , .B2( u0_u3_u3_n155 ) , .B1( u0_u3_u3_n156 ) , .ZN( u0_u3_u3_n157 ) );
  INV_X1 u0_u3_u3_U4 (.A( u0_u3_u3_n129 ) , .ZN( u0_u3_u3_n183 ) );
  AOI211_X1 u0_u3_u3_U40 (.ZN( u0_u3_u3_n109 ) , .A( u0_u3_u3_n119 ) , .C2( u0_u3_u3_n129 ) , .B( u0_u3_u3_n138 ) , .C1( u0_u3_u3_n141 ) );
  INV_X1 u0_u3_u3_U41 (.A( u0_u3_u3_n121 ) , .ZN( u0_u3_u3_n164 ) );
  NAND2_X1 u0_u3_u3_U42 (.ZN( u0_u3_u3_n133 ) , .A1( u0_u3_u3_n154 ) , .A2( u0_u3_u3_n164 ) );
  OAI211_X1 u0_u3_u3_U43 (.B( u0_u3_u3_n127 ) , .ZN( u0_u3_u3_n139 ) , .C1( u0_u3_u3_n150 ) , .C2( u0_u3_u3_n154 ) , .A( u0_u3_u3_n184 ) );
  INV_X1 u0_u3_u3_U44 (.A( u0_u3_u3_n125 ) , .ZN( u0_u3_u3_n184 ) );
  AOI221_X1 u0_u3_u3_U45 (.A( u0_u3_u3_n126 ) , .ZN( u0_u3_u3_n127 ) , .C2( u0_u3_u3_n132 ) , .C1( u0_u3_u3_n169 ) , .B2( u0_u3_u3_n170 ) , .B1( u0_u3_u3_n174 ) );
  OAI22_X1 u0_u3_u3_U46 (.A1( u0_u3_u3_n124 ) , .ZN( u0_u3_u3_n125 ) , .B2( u0_u3_u3_n145 ) , .A2( u0_u3_u3_n165 ) , .B1( u0_u3_u3_n167 ) );
  NOR2_X1 u0_u3_u3_U47 (.A1( u0_u3_u3_n113 ) , .ZN( u0_u3_u3_n131 ) , .A2( u0_u3_u3_n154 ) );
  NAND2_X1 u0_u3_u3_U48 (.A1( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n150 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U49 (.A2( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n155 ) , .A1( u0_u3_u3_n97 ) );
  INV_X1 u0_u3_u3_U5 (.A( u0_u3_u3_n117 ) , .ZN( u0_u3_u3_n178 ) );
  INV_X1 u0_u3_u3_U50 (.A( u0_u3_u3_n141 ) , .ZN( u0_u3_u3_n167 ) );
  AOI21_X1 u0_u3_u3_U51 (.B2( u0_u3_u3_n114 ) , .B1( u0_u3_u3_n146 ) , .A( u0_u3_u3_n154 ) , .ZN( u0_u3_u3_n94 ) );
  AOI21_X1 u0_u3_u3_U52 (.ZN( u0_u3_u3_n110 ) , .B2( u0_u3_u3_n142 ) , .B1( u0_u3_u3_n186 ) , .A( u0_u3_u3_n95 ) );
  INV_X1 u0_u3_u3_U53 (.A( u0_u3_u3_n145 ) , .ZN( u0_u3_u3_n186 ) );
  AOI21_X1 u0_u3_u3_U54 (.B1( u0_u3_u3_n124 ) , .A( u0_u3_u3_n149 ) , .B2( u0_u3_u3_n155 ) , .ZN( u0_u3_u3_n95 ) );
  INV_X1 u0_u3_u3_U55 (.A( u0_u3_u3_n149 ) , .ZN( u0_u3_u3_n169 ) );
  NAND2_X1 u0_u3_u3_U56 (.ZN( u0_u3_u3_n124 ) , .A1( u0_u3_u3_n96 ) , .A2( u0_u3_u3_n97 ) );
  NAND2_X1 u0_u3_u3_U57 (.A2( u0_u3_u3_n100 ) , .ZN( u0_u3_u3_n146 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U58 (.A1( u0_u3_u3_n101 ) , .ZN( u0_u3_u3_n145 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U59 (.A1( u0_u3_u3_n100 ) , .ZN( u0_u3_u3_n156 ) , .A2( u0_u3_u3_n99 ) );
  AOI221_X1 u0_u3_u3_U6 (.A( u0_u3_u3_n131 ) , .C2( u0_u3_u3_n132 ) , .C1( u0_u3_u3_n133 ) , .ZN( u0_u3_u3_n134 ) , .B1( u0_u3_u3_n143 ) , .B2( u0_u3_u3_n177 ) );
  NAND2_X1 u0_u3_u3_U60 (.A2( u0_u3_u3_n101 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n148 ) );
  NAND2_X1 u0_u3_u3_U61 (.A1( u0_u3_u3_n100 ) , .A2( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n128 ) );
  NAND2_X1 u0_u3_u3_U62 (.A2( u0_u3_u3_n101 ) , .A1( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n152 ) );
  NAND2_X1 u0_u3_u3_U63 (.A2( u0_u3_u3_n101 ) , .ZN( u0_u3_u3_n114 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U64 (.ZN( u0_u3_u3_n107 ) , .A1( u0_u3_u3_n97 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U65 (.A2( u0_u3_u3_n100 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n113 ) );
  NAND2_X1 u0_u3_u3_U66 (.A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n153 ) , .A2( u0_u3_u3_n97 ) );
  NAND2_X1 u0_u3_u3_U67 (.A2( u0_u3_u3_n103 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n130 ) );
  NAND2_X1 u0_u3_u3_U68 (.A2( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n144 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U69 (.A1( u0_u3_u3_n102 ) , .A2( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n108 ) );
  OAI22_X1 u0_u3_u3_U7 (.B2( u0_u3_u3_n147 ) , .A2( u0_u3_u3_n148 ) , .ZN( u0_u3_u3_n160 ) , .B1( u0_u3_u3_n165 ) , .A1( u0_u3_u3_n168 ) );
  NOR2_X1 u0_u3_u3_U70 (.A2( u0_u3_X_19 ) , .A1( u0_u3_X_20 ) , .ZN( u0_u3_u3_n99 ) );
  NOR2_X1 u0_u3_u3_U71 (.A2( u0_u3_X_21 ) , .A1( u0_u3_X_24 ) , .ZN( u0_u3_u3_n103 ) );
  NOR2_X1 u0_u3_u3_U72 (.A2( u0_u3_X_24 ) , .A1( u0_u3_u3_n171 ) , .ZN( u0_u3_u3_n97 ) );
  NOR2_X1 u0_u3_u3_U73 (.A2( u0_u3_X_19 ) , .A1( u0_u3_u3_n172 ) , .ZN( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U74 (.A1( u0_u3_X_22 ) , .A2( u0_u3_X_23 ) , .ZN( u0_u3_u3_n154 ) );
  AND2_X1 u0_u3_u3_U75 (.A1( u0_u3_X_24 ) , .ZN( u0_u3_u3_n101 ) , .A2( u0_u3_u3_n171 ) );
  AND2_X1 u0_u3_u3_U76 (.A1( u0_u3_X_19 ) , .ZN( u0_u3_u3_n102 ) , .A2( u0_u3_u3_n172 ) );
  AND2_X1 u0_u3_u3_U77 (.A1( u0_u3_X_21 ) , .A2( u0_u3_X_24 ) , .ZN( u0_u3_u3_n100 ) );
  AND2_X1 u0_u3_u3_U78 (.A2( u0_u3_X_19 ) , .A1( u0_u3_X_20 ) , .ZN( u0_u3_u3_n104 ) );
  INV_X1 u0_u3_u3_U79 (.A( u0_u3_X_21 ) , .ZN( u0_u3_u3_n171 ) );
  AND3_X1 u0_u3_u3_U8 (.A3( u0_u3_u3_n144 ) , .A2( u0_u3_u3_n145 ) , .A1( u0_u3_u3_n146 ) , .ZN( u0_u3_u3_n147 ) );
  INV_X1 u0_u3_u3_U80 (.A( u0_u3_X_20 ) , .ZN( u0_u3_u3_n172 ) );
  INV_X1 u0_u3_u3_U81 (.A( u0_u3_X_22 ) , .ZN( u0_u3_u3_n166 ) );
  NAND4_X1 u0_u3_u3_U82 (.ZN( u0_out3_26 ) , .A4( u0_u3_u3_n109 ) , .A3( u0_u3_u3_n110 ) , .A2( u0_u3_u3_n111 ) , .A1( u0_u3_u3_n173 ) );
  INV_X1 u0_u3_u3_U83 (.ZN( u0_u3_u3_n173 ) , .A( u0_u3_u3_n94 ) );
  OAI21_X1 u0_u3_u3_U84 (.ZN( u0_u3_u3_n111 ) , .B2( u0_u3_u3_n117 ) , .A( u0_u3_u3_n133 ) , .B1( u0_u3_u3_n176 ) );
  NAND4_X1 u0_u3_u3_U85 (.ZN( u0_out3_1 ) , .A4( u0_u3_u3_n161 ) , .A3( u0_u3_u3_n162 ) , .A2( u0_u3_u3_n163 ) , .A1( u0_u3_u3_n185 ) );
  NAND2_X1 u0_u3_u3_U86 (.ZN( u0_u3_u3_n163 ) , .A2( u0_u3_u3_n170 ) , .A1( u0_u3_u3_n176 ) );
  AOI22_X1 u0_u3_u3_U87 (.B2( u0_u3_u3_n140 ) , .B1( u0_u3_u3_n141 ) , .A2( u0_u3_u3_n142 ) , .ZN( u0_u3_u3_n162 ) , .A1( u0_u3_u3_n177 ) );
  NAND4_X1 u0_u3_u3_U88 (.ZN( u0_out3_20 ) , .A4( u0_u3_u3_n122 ) , .A3( u0_u3_u3_n123 ) , .A1( u0_u3_u3_n175 ) , .A2( u0_u3_u3_n180 ) );
  INV_X1 u0_u3_u3_U89 (.A( u0_u3_u3_n126 ) , .ZN( u0_u3_u3_n180 ) );
  INV_X1 u0_u3_u3_U9 (.A( u0_u3_u3_n143 ) , .ZN( u0_u3_u3_n168 ) );
  INV_X1 u0_u3_u3_U90 (.A( u0_u3_u3_n112 ) , .ZN( u0_u3_u3_n175 ) );
  OR4_X1 u0_u3_u3_U91 (.ZN( u0_out3_10 ) , .A4( u0_u3_u3_n136 ) , .A3( u0_u3_u3_n137 ) , .A1( u0_u3_u3_n138 ) , .A2( u0_u3_u3_n139 ) );
  OAI222_X1 u0_u3_u3_U92 (.C1( u0_u3_u3_n128 ) , .ZN( u0_u3_u3_n137 ) , .B1( u0_u3_u3_n148 ) , .A2( u0_u3_u3_n150 ) , .B2( u0_u3_u3_n154 ) , .C2( u0_u3_u3_n164 ) , .A1( u0_u3_u3_n167 ) );
  AOI211_X1 u0_u3_u3_U93 (.B( u0_u3_u3_n119 ) , .A( u0_u3_u3_n120 ) , .C2( u0_u3_u3_n121 ) , .ZN( u0_u3_u3_n122 ) , .C1( u0_u3_u3_n179 ) );
  OAI221_X1 u0_u3_u3_U94 (.A( u0_u3_u3_n134 ) , .B2( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n136 ) , .C1( u0_u3_u3_n149 ) , .B1( u0_u3_u3_n151 ) , .C2( u0_u3_u3_n183 ) );
  NOR2_X1 u0_u3_u3_U95 (.A2( u0_u3_X_23 ) , .ZN( u0_u3_u3_n141 ) , .A1( u0_u3_u3_n166 ) );
  NAND2_X1 u0_u3_u3_U96 (.A1( u0_u3_X_23 ) , .ZN( u0_u3_u3_n149 ) , .A2( u0_u3_u3_n166 ) );
  NOR2_X1 u0_u3_u3_U97 (.A2( u0_u3_X_22 ) , .A1( u0_u3_X_23 ) , .ZN( u0_u3_u3_n121 ) );
  NAND3_X1 u0_u3_u3_U98 (.A1( u0_u3_u3_n114 ) , .ZN( u0_u3_u3_n115 ) , .A2( u0_u3_u3_n145 ) , .A3( u0_u3_u3_n153 ) );
  NAND3_X1 u0_u3_u3_U99 (.ZN( u0_u3_u3_n129 ) , .A2( u0_u3_u3_n144 ) , .A1( u0_u3_u3_n153 ) , .A3( u0_u3_u3_n182 ) );
  OAI22_X1 u0_u3_u4_U10 (.B2( u0_u3_u4_n135 ) , .ZN( u0_u3_u4_n137 ) , .B1( u0_u3_u4_n153 ) , .A1( u0_u3_u4_n155 ) , .A2( u0_u3_u4_n171 ) );
  AND3_X1 u0_u3_u4_U11 (.A2( u0_u3_u4_n134 ) , .ZN( u0_u3_u4_n135 ) , .A3( u0_u3_u4_n145 ) , .A1( u0_u3_u4_n157 ) );
  OR3_X1 u0_u3_u4_U12 (.A3( u0_u3_u4_n114 ) , .A2( u0_u3_u4_n115 ) , .A1( u0_u3_u4_n116 ) , .ZN( u0_u3_u4_n136 ) );
  AOI21_X1 u0_u3_u4_U13 (.A( u0_u3_u4_n113 ) , .ZN( u0_u3_u4_n116 ) , .B2( u0_u3_u4_n173 ) , .B1( u0_u3_u4_n174 ) );
  AOI21_X1 u0_u3_u4_U14 (.ZN( u0_u3_u4_n115 ) , .B2( u0_u3_u4_n145 ) , .B1( u0_u3_u4_n146 ) , .A( u0_u3_u4_n156 ) );
  OAI22_X1 u0_u3_u4_U15 (.ZN( u0_u3_u4_n114 ) , .A2( u0_u3_u4_n121 ) , .B1( u0_u3_u4_n160 ) , .B2( u0_u3_u4_n170 ) , .A1( u0_u3_u4_n171 ) );
  NAND2_X1 u0_u3_u4_U16 (.ZN( u0_u3_u4_n132 ) , .A2( u0_u3_u4_n170 ) , .A1( u0_u3_u4_n173 ) );
  AOI21_X1 u0_u3_u4_U17 (.B2( u0_u3_u4_n160 ) , .B1( u0_u3_u4_n161 ) , .ZN( u0_u3_u4_n162 ) , .A( u0_u3_u4_n170 ) );
  AOI21_X1 u0_u3_u4_U18 (.ZN( u0_u3_u4_n107 ) , .B2( u0_u3_u4_n143 ) , .A( u0_u3_u4_n174 ) , .B1( u0_u3_u4_n184 ) );
  AOI21_X1 u0_u3_u4_U19 (.B2( u0_u3_u4_n158 ) , .B1( u0_u3_u4_n159 ) , .ZN( u0_u3_u4_n163 ) , .A( u0_u3_u4_n174 ) );
  AOI21_X1 u0_u3_u4_U20 (.A( u0_u3_u4_n153 ) , .B2( u0_u3_u4_n154 ) , .B1( u0_u3_u4_n155 ) , .ZN( u0_u3_u4_n165 ) );
  AOI21_X1 u0_u3_u4_U21 (.A( u0_u3_u4_n156 ) , .B2( u0_u3_u4_n157 ) , .ZN( u0_u3_u4_n164 ) , .B1( u0_u3_u4_n184 ) );
  INV_X1 u0_u3_u4_U22 (.A( u0_u3_u4_n138 ) , .ZN( u0_u3_u4_n170 ) );
  AND2_X1 u0_u3_u4_U23 (.A2( u0_u3_u4_n120 ) , .ZN( u0_u3_u4_n155 ) , .A1( u0_u3_u4_n160 ) );
  INV_X1 u0_u3_u4_U24 (.A( u0_u3_u4_n156 ) , .ZN( u0_u3_u4_n175 ) );
  NAND2_X1 u0_u3_u4_U25 (.A2( u0_u3_u4_n118 ) , .ZN( u0_u3_u4_n131 ) , .A1( u0_u3_u4_n147 ) );
  NAND2_X1 u0_u3_u4_U26 (.A1( u0_u3_u4_n119 ) , .A2( u0_u3_u4_n120 ) , .ZN( u0_u3_u4_n130 ) );
  NAND2_X1 u0_u3_u4_U27 (.ZN( u0_u3_u4_n117 ) , .A2( u0_u3_u4_n118 ) , .A1( u0_u3_u4_n148 ) );
  NAND2_X1 u0_u3_u4_U28 (.ZN( u0_u3_u4_n129 ) , .A1( u0_u3_u4_n134 ) , .A2( u0_u3_u4_n148 ) );
  AND3_X1 u0_u3_u4_U29 (.A1( u0_u3_u4_n119 ) , .A2( u0_u3_u4_n143 ) , .A3( u0_u3_u4_n154 ) , .ZN( u0_u3_u4_n161 ) );
  NOR2_X1 u0_u3_u4_U3 (.ZN( u0_u3_u4_n121 ) , .A1( u0_u3_u4_n181 ) , .A2( u0_u3_u4_n182 ) );
  AND2_X1 u0_u3_u4_U30 (.A1( u0_u3_u4_n145 ) , .A2( u0_u3_u4_n147 ) , .ZN( u0_u3_u4_n159 ) );
  INV_X1 u0_u3_u4_U31 (.A( u0_u3_u4_n158 ) , .ZN( u0_u3_u4_n182 ) );
  INV_X1 u0_u3_u4_U32 (.ZN( u0_u3_u4_n181 ) , .A( u0_u3_u4_n96 ) );
  INV_X1 u0_u3_u4_U33 (.A( u0_u3_u4_n144 ) , .ZN( u0_u3_u4_n179 ) );
  INV_X1 u0_u3_u4_U34 (.A( u0_u3_u4_n157 ) , .ZN( u0_u3_u4_n178 ) );
  NAND2_X1 u0_u3_u4_U35 (.A2( u0_u3_u4_n154 ) , .A1( u0_u3_u4_n96 ) , .ZN( u0_u3_u4_n97 ) );
  INV_X1 u0_u3_u4_U36 (.ZN( u0_u3_u4_n186 ) , .A( u0_u3_u4_n95 ) );
  OAI221_X1 u0_u3_u4_U37 (.C1( u0_u3_u4_n134 ) , .B1( u0_u3_u4_n158 ) , .B2( u0_u3_u4_n171 ) , .C2( u0_u3_u4_n173 ) , .A( u0_u3_u4_n94 ) , .ZN( u0_u3_u4_n95 ) );
  AOI222_X1 u0_u3_u4_U38 (.B2( u0_u3_u4_n132 ) , .A1( u0_u3_u4_n138 ) , .C2( u0_u3_u4_n175 ) , .A2( u0_u3_u4_n179 ) , .C1( u0_u3_u4_n181 ) , .B1( u0_u3_u4_n185 ) , .ZN( u0_u3_u4_n94 ) );
  INV_X1 u0_u3_u4_U39 (.A( u0_u3_u4_n113 ) , .ZN( u0_u3_u4_n185 ) );
  INV_X1 u0_u3_u4_U4 (.A( u0_u3_u4_n117 ) , .ZN( u0_u3_u4_n184 ) );
  INV_X1 u0_u3_u4_U40 (.A( u0_u3_u4_n143 ) , .ZN( u0_u3_u4_n183 ) );
  NOR2_X1 u0_u3_u4_U41 (.ZN( u0_u3_u4_n138 ) , .A1( u0_u3_u4_n168 ) , .A2( u0_u3_u4_n169 ) );
  NOR2_X1 u0_u3_u4_U42 (.A1( u0_u3_u4_n150 ) , .A2( u0_u3_u4_n152 ) , .ZN( u0_u3_u4_n153 ) );
  NOR2_X1 u0_u3_u4_U43 (.A2( u0_u3_u4_n128 ) , .A1( u0_u3_u4_n138 ) , .ZN( u0_u3_u4_n156 ) );
  AOI22_X1 u0_u3_u4_U44 (.B2( u0_u3_u4_n122 ) , .A1( u0_u3_u4_n123 ) , .ZN( u0_u3_u4_n124 ) , .B1( u0_u3_u4_n128 ) , .A2( u0_u3_u4_n172 ) );
  INV_X1 u0_u3_u4_U45 (.A( u0_u3_u4_n153 ) , .ZN( u0_u3_u4_n172 ) );
  NAND2_X1 u0_u3_u4_U46 (.A2( u0_u3_u4_n120 ) , .ZN( u0_u3_u4_n123 ) , .A1( u0_u3_u4_n161 ) );
  AOI22_X1 u0_u3_u4_U47 (.B2( u0_u3_u4_n132 ) , .A2( u0_u3_u4_n133 ) , .ZN( u0_u3_u4_n140 ) , .A1( u0_u3_u4_n150 ) , .B1( u0_u3_u4_n179 ) );
  NAND2_X1 u0_u3_u4_U48 (.ZN( u0_u3_u4_n133 ) , .A2( u0_u3_u4_n146 ) , .A1( u0_u3_u4_n154 ) );
  NAND2_X1 u0_u3_u4_U49 (.A1( u0_u3_u4_n103 ) , .ZN( u0_u3_u4_n154 ) , .A2( u0_u3_u4_n98 ) );
  NOR4_X1 u0_u3_u4_U5 (.A4( u0_u3_u4_n106 ) , .A3( u0_u3_u4_n107 ) , .A2( u0_u3_u4_n108 ) , .A1( u0_u3_u4_n109 ) , .ZN( u0_u3_u4_n110 ) );
  NAND2_X1 u0_u3_u4_U50 (.A1( u0_u3_u4_n101 ) , .ZN( u0_u3_u4_n158 ) , .A2( u0_u3_u4_n99 ) );
  AOI21_X1 u0_u3_u4_U51 (.ZN( u0_u3_u4_n127 ) , .A( u0_u3_u4_n136 ) , .B2( u0_u3_u4_n150 ) , .B1( u0_u3_u4_n180 ) );
  INV_X1 u0_u3_u4_U52 (.A( u0_u3_u4_n160 ) , .ZN( u0_u3_u4_n180 ) );
  NAND2_X1 u0_u3_u4_U53 (.A2( u0_u3_u4_n104 ) , .A1( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n146 ) );
  NAND2_X1 u0_u3_u4_U54 (.A2( u0_u3_u4_n101 ) , .A1( u0_u3_u4_n102 ) , .ZN( u0_u3_u4_n160 ) );
  NAND2_X1 u0_u3_u4_U55 (.ZN( u0_u3_u4_n134 ) , .A1( u0_u3_u4_n98 ) , .A2( u0_u3_u4_n99 ) );
  NAND2_X1 u0_u3_u4_U56 (.A1( u0_u3_u4_n103 ) , .A2( u0_u3_u4_n104 ) , .ZN( u0_u3_u4_n143 ) );
  NAND2_X1 u0_u3_u4_U57 (.A2( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n145 ) , .A1( u0_u3_u4_n98 ) );
  NAND2_X1 u0_u3_u4_U58 (.A1( u0_u3_u4_n100 ) , .A2( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n120 ) );
  NAND2_X1 u0_u3_u4_U59 (.A1( u0_u3_u4_n102 ) , .A2( u0_u3_u4_n104 ) , .ZN( u0_u3_u4_n148 ) );
  AOI21_X1 u0_u3_u4_U6 (.ZN( u0_u3_u4_n106 ) , .B2( u0_u3_u4_n146 ) , .B1( u0_u3_u4_n158 ) , .A( u0_u3_u4_n170 ) );
  NAND2_X1 u0_u3_u4_U60 (.A2( u0_u3_u4_n100 ) , .A1( u0_u3_u4_n103 ) , .ZN( u0_u3_u4_n157 ) );
  INV_X1 u0_u3_u4_U61 (.A( u0_u3_u4_n150 ) , .ZN( u0_u3_u4_n173 ) );
  INV_X1 u0_u3_u4_U62 (.A( u0_u3_u4_n152 ) , .ZN( u0_u3_u4_n171 ) );
  NAND2_X1 u0_u3_u4_U63 (.A1( u0_u3_u4_n100 ) , .ZN( u0_u3_u4_n118 ) , .A2( u0_u3_u4_n99 ) );
  NAND2_X1 u0_u3_u4_U64 (.A2( u0_u3_u4_n100 ) , .A1( u0_u3_u4_n102 ) , .ZN( u0_u3_u4_n144 ) );
  NAND2_X1 u0_u3_u4_U65 (.A2( u0_u3_u4_n101 ) , .A1( u0_u3_u4_n105 ) , .ZN( u0_u3_u4_n96 ) );
  INV_X1 u0_u3_u4_U66 (.A( u0_u3_u4_n128 ) , .ZN( u0_u3_u4_n174 ) );
  NAND2_X1 u0_u3_u4_U67 (.A2( u0_u3_u4_n102 ) , .ZN( u0_u3_u4_n119 ) , .A1( u0_u3_u4_n98 ) );
  NAND2_X1 u0_u3_u4_U68 (.A2( u0_u3_u4_n101 ) , .A1( u0_u3_u4_n103 ) , .ZN( u0_u3_u4_n147 ) );
  NAND2_X1 u0_u3_u4_U69 (.A2( u0_u3_u4_n104 ) , .ZN( u0_u3_u4_n113 ) , .A1( u0_u3_u4_n99 ) );
  AOI21_X1 u0_u3_u4_U7 (.ZN( u0_u3_u4_n109 ) , .A( u0_u3_u4_n153 ) , .B1( u0_u3_u4_n159 ) , .B2( u0_u3_u4_n184 ) );
  NOR2_X1 u0_u3_u4_U70 (.A2( u0_u3_X_28 ) , .ZN( u0_u3_u4_n150 ) , .A1( u0_u3_u4_n168 ) );
  NOR2_X1 u0_u3_u4_U71 (.A2( u0_u3_X_29 ) , .ZN( u0_u3_u4_n152 ) , .A1( u0_u3_u4_n169 ) );
  NOR2_X1 u0_u3_u4_U72 (.A2( u0_u3_X_30 ) , .ZN( u0_u3_u4_n105 ) , .A1( u0_u3_u4_n176 ) );
  NOR2_X1 u0_u3_u4_U73 (.A2( u0_u3_X_26 ) , .ZN( u0_u3_u4_n100 ) , .A1( u0_u3_u4_n177 ) );
  NOR2_X1 u0_u3_u4_U74 (.A2( u0_u3_X_28 ) , .A1( u0_u3_X_29 ) , .ZN( u0_u3_u4_n128 ) );
  NOR2_X1 u0_u3_u4_U75 (.A2( u0_u3_X_27 ) , .A1( u0_u3_X_30 ) , .ZN( u0_u3_u4_n102 ) );
  NOR2_X1 u0_u3_u4_U76 (.A2( u0_u3_X_25 ) , .A1( u0_u3_X_26 ) , .ZN( u0_u3_u4_n98 ) );
  AND2_X1 u0_u3_u4_U77 (.A2( u0_u3_X_25 ) , .A1( u0_u3_X_26 ) , .ZN( u0_u3_u4_n104 ) );
  AND2_X1 u0_u3_u4_U78 (.A1( u0_u3_X_30 ) , .A2( u0_u3_u4_n176 ) , .ZN( u0_u3_u4_n99 ) );
  AND2_X1 u0_u3_u4_U79 (.A1( u0_u3_X_26 ) , .ZN( u0_u3_u4_n101 ) , .A2( u0_u3_u4_n177 ) );
  AOI21_X1 u0_u3_u4_U8 (.ZN( u0_u3_u4_n108 ) , .B2( u0_u3_u4_n134 ) , .B1( u0_u3_u4_n155 ) , .A( u0_u3_u4_n156 ) );
  AND2_X1 u0_u3_u4_U80 (.A1( u0_u3_X_27 ) , .A2( u0_u3_X_30 ) , .ZN( u0_u3_u4_n103 ) );
  INV_X1 u0_u3_u4_U81 (.A( u0_u3_X_28 ) , .ZN( u0_u3_u4_n169 ) );
  INV_X1 u0_u3_u4_U82 (.A( u0_u3_X_29 ) , .ZN( u0_u3_u4_n168 ) );
  INV_X1 u0_u3_u4_U83 (.A( u0_u3_X_25 ) , .ZN( u0_u3_u4_n177 ) );
  INV_X1 u0_u3_u4_U84 (.A( u0_u3_X_27 ) , .ZN( u0_u3_u4_n176 ) );
  NAND4_X1 u0_u3_u4_U85 (.ZN( u0_out3_25 ) , .A4( u0_u3_u4_n139 ) , .A3( u0_u3_u4_n140 ) , .A2( u0_u3_u4_n141 ) , .A1( u0_u3_u4_n142 ) );
  OAI21_X1 u0_u3_u4_U86 (.A( u0_u3_u4_n128 ) , .B2( u0_u3_u4_n129 ) , .B1( u0_u3_u4_n130 ) , .ZN( u0_u3_u4_n142 ) );
  OAI21_X1 u0_u3_u4_U87 (.B2( u0_u3_u4_n131 ) , .ZN( u0_u3_u4_n141 ) , .A( u0_u3_u4_n175 ) , .B1( u0_u3_u4_n183 ) );
  NAND4_X1 u0_u3_u4_U88 (.ZN( u0_out3_14 ) , .A4( u0_u3_u4_n124 ) , .A3( u0_u3_u4_n125 ) , .A2( u0_u3_u4_n126 ) , .A1( u0_u3_u4_n127 ) );
  AOI22_X1 u0_u3_u4_U89 (.B2( u0_u3_u4_n117 ) , .ZN( u0_u3_u4_n126 ) , .A1( u0_u3_u4_n129 ) , .B1( u0_u3_u4_n152 ) , .A2( u0_u3_u4_n175 ) );
  AOI211_X1 u0_u3_u4_U9 (.B( u0_u3_u4_n136 ) , .A( u0_u3_u4_n137 ) , .C2( u0_u3_u4_n138 ) , .ZN( u0_u3_u4_n139 ) , .C1( u0_u3_u4_n182 ) );
  AOI22_X1 u0_u3_u4_U90 (.ZN( u0_u3_u4_n125 ) , .B2( u0_u3_u4_n131 ) , .A2( u0_u3_u4_n132 ) , .B1( u0_u3_u4_n138 ) , .A1( u0_u3_u4_n178 ) );
  AOI22_X1 u0_u3_u4_U91 (.B2( u0_u3_u4_n149 ) , .B1( u0_u3_u4_n150 ) , .A2( u0_u3_u4_n151 ) , .A1( u0_u3_u4_n152 ) , .ZN( u0_u3_u4_n167 ) );
  NOR4_X1 u0_u3_u4_U92 (.A4( u0_u3_u4_n162 ) , .A3( u0_u3_u4_n163 ) , .A2( u0_u3_u4_n164 ) , .A1( u0_u3_u4_n165 ) , .ZN( u0_u3_u4_n166 ) );
  NAND4_X1 u0_u3_u4_U93 (.ZN( u0_out3_8 ) , .A4( u0_u3_u4_n110 ) , .A3( u0_u3_u4_n111 ) , .A2( u0_u3_u4_n112 ) , .A1( u0_u3_u4_n186 ) );
  NAND2_X1 u0_u3_u4_U94 (.ZN( u0_u3_u4_n112 ) , .A2( u0_u3_u4_n130 ) , .A1( u0_u3_u4_n150 ) );
  AOI22_X1 u0_u3_u4_U95 (.ZN( u0_u3_u4_n111 ) , .B2( u0_u3_u4_n132 ) , .A1( u0_u3_u4_n152 ) , .B1( u0_u3_u4_n178 ) , .A2( u0_u3_u4_n97 ) );
  NAND3_X1 u0_u3_u4_U96 (.ZN( u0_out3_3 ) , .A3( u0_u3_u4_n166 ) , .A1( u0_u3_u4_n167 ) , .A2( u0_u3_u4_n186 ) );
  NAND3_X1 u0_u3_u4_U97 (.A3( u0_u3_u4_n146 ) , .A2( u0_u3_u4_n147 ) , .A1( u0_u3_u4_n148 ) , .ZN( u0_u3_u4_n149 ) );
  NAND3_X1 u0_u3_u4_U98 (.A3( u0_u3_u4_n143 ) , .A2( u0_u3_u4_n144 ) , .A1( u0_u3_u4_n145 ) , .ZN( u0_u3_u4_n151 ) );
  NAND3_X1 u0_u3_u4_U99 (.A3( u0_u3_u4_n121 ) , .ZN( u0_u3_u4_n122 ) , .A2( u0_u3_u4_n144 ) , .A1( u0_u3_u4_n154 ) );
  INV_X1 u0_u3_u5_U10 (.A( u0_u3_u5_n121 ) , .ZN( u0_u3_u5_n177 ) );
  NOR3_X1 u0_u3_u5_U100 (.A3( u0_u3_u5_n141 ) , .A1( u0_u3_u5_n142 ) , .ZN( u0_u3_u5_n143 ) , .A2( u0_u3_u5_n191 ) );
  NAND4_X1 u0_u3_u5_U101 (.ZN( u0_out3_4 ) , .A4( u0_u3_u5_n112 ) , .A2( u0_u3_u5_n113 ) , .A1( u0_u3_u5_n114 ) , .A3( u0_u3_u5_n195 ) );
  AOI211_X1 u0_u3_u5_U102 (.A( u0_u3_u5_n110 ) , .C1( u0_u3_u5_n111 ) , .ZN( u0_u3_u5_n112 ) , .B( u0_u3_u5_n118 ) , .C2( u0_u3_u5_n177 ) );
  AOI222_X1 u0_u3_u5_U103 (.ZN( u0_u3_u5_n113 ) , .A1( u0_u3_u5_n131 ) , .C1( u0_u3_u5_n148 ) , .B2( u0_u3_u5_n174 ) , .C2( u0_u3_u5_n178 ) , .A2( u0_u3_u5_n179 ) , .B1( u0_u3_u5_n99 ) );
  NAND3_X1 u0_u3_u5_U104 (.A2( u0_u3_u5_n154 ) , .A3( u0_u3_u5_n158 ) , .A1( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n99 ) );
  NOR2_X1 u0_u3_u5_U11 (.ZN( u0_u3_u5_n160 ) , .A2( u0_u3_u5_n173 ) , .A1( u0_u3_u5_n177 ) );
  INV_X1 u0_u3_u5_U12 (.A( u0_u3_u5_n150 ) , .ZN( u0_u3_u5_n174 ) );
  AOI21_X1 u0_u3_u5_U13 (.A( u0_u3_u5_n160 ) , .B2( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n162 ) , .B1( u0_u3_u5_n192 ) );
  INV_X1 u0_u3_u5_U14 (.A( u0_u3_u5_n159 ) , .ZN( u0_u3_u5_n192 ) );
  AOI21_X1 u0_u3_u5_U15 (.A( u0_u3_u5_n156 ) , .B2( u0_u3_u5_n157 ) , .B1( u0_u3_u5_n158 ) , .ZN( u0_u3_u5_n163 ) );
  AOI21_X1 u0_u3_u5_U16 (.B2( u0_u3_u5_n139 ) , .B1( u0_u3_u5_n140 ) , .ZN( u0_u3_u5_n141 ) , .A( u0_u3_u5_n150 ) );
  OAI21_X1 u0_u3_u5_U17 (.A( u0_u3_u5_n133 ) , .B2( u0_u3_u5_n134 ) , .B1( u0_u3_u5_n135 ) , .ZN( u0_u3_u5_n142 ) );
  OAI21_X1 u0_u3_u5_U18 (.ZN( u0_u3_u5_n133 ) , .B2( u0_u3_u5_n147 ) , .A( u0_u3_u5_n173 ) , .B1( u0_u3_u5_n188 ) );
  NAND2_X1 u0_u3_u5_U19 (.A2( u0_u3_u5_n119 ) , .A1( u0_u3_u5_n123 ) , .ZN( u0_u3_u5_n137 ) );
  INV_X1 u0_u3_u5_U20 (.A( u0_u3_u5_n155 ) , .ZN( u0_u3_u5_n194 ) );
  NAND2_X1 u0_u3_u5_U21 (.A1( u0_u3_u5_n121 ) , .ZN( u0_u3_u5_n132 ) , .A2( u0_u3_u5_n172 ) );
  NAND2_X1 u0_u3_u5_U22 (.A2( u0_u3_u5_n122 ) , .ZN( u0_u3_u5_n136 ) , .A1( u0_u3_u5_n154 ) );
  NAND2_X1 u0_u3_u5_U23 (.A2( u0_u3_u5_n119 ) , .A1( u0_u3_u5_n120 ) , .ZN( u0_u3_u5_n159 ) );
  INV_X1 u0_u3_u5_U24 (.A( u0_u3_u5_n156 ) , .ZN( u0_u3_u5_n175 ) );
  INV_X1 u0_u3_u5_U25 (.A( u0_u3_u5_n158 ) , .ZN( u0_u3_u5_n188 ) );
  INV_X1 u0_u3_u5_U26 (.A( u0_u3_u5_n152 ) , .ZN( u0_u3_u5_n179 ) );
  INV_X1 u0_u3_u5_U27 (.A( u0_u3_u5_n140 ) , .ZN( u0_u3_u5_n182 ) );
  INV_X1 u0_u3_u5_U28 (.A( u0_u3_u5_n151 ) , .ZN( u0_u3_u5_n183 ) );
  INV_X1 u0_u3_u5_U29 (.A( u0_u3_u5_n123 ) , .ZN( u0_u3_u5_n185 ) );
  NOR2_X1 u0_u3_u5_U3 (.ZN( u0_u3_u5_n134 ) , .A1( u0_u3_u5_n183 ) , .A2( u0_u3_u5_n190 ) );
  INV_X1 u0_u3_u5_U30 (.A( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n184 ) );
  INV_X1 u0_u3_u5_U31 (.A( u0_u3_u5_n139 ) , .ZN( u0_u3_u5_n189 ) );
  INV_X1 u0_u3_u5_U32 (.A( u0_u3_u5_n157 ) , .ZN( u0_u3_u5_n190 ) );
  INV_X1 u0_u3_u5_U33 (.A( u0_u3_u5_n120 ) , .ZN( u0_u3_u5_n193 ) );
  NAND2_X1 u0_u3_u5_U34 (.ZN( u0_u3_u5_n111 ) , .A1( u0_u3_u5_n140 ) , .A2( u0_u3_u5_n155 ) );
  INV_X1 u0_u3_u5_U35 (.A( u0_u3_u5_n117 ) , .ZN( u0_u3_u5_n196 ) );
  OAI221_X1 u0_u3_u5_U36 (.A( u0_u3_u5_n116 ) , .ZN( u0_u3_u5_n117 ) , .B2( u0_u3_u5_n119 ) , .C1( u0_u3_u5_n153 ) , .C2( u0_u3_u5_n158 ) , .B1( u0_u3_u5_n172 ) );
  AOI222_X1 u0_u3_u5_U37 (.ZN( u0_u3_u5_n116 ) , .B2( u0_u3_u5_n145 ) , .C1( u0_u3_u5_n148 ) , .A2( u0_u3_u5_n174 ) , .C2( u0_u3_u5_n177 ) , .B1( u0_u3_u5_n187 ) , .A1( u0_u3_u5_n193 ) );
  INV_X1 u0_u3_u5_U38 (.A( u0_u3_u5_n115 ) , .ZN( u0_u3_u5_n187 ) );
  NOR2_X1 u0_u3_u5_U39 (.ZN( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n170 ) , .A2( u0_u3_u5_n180 ) );
  INV_X1 u0_u3_u5_U4 (.A( u0_u3_u5_n138 ) , .ZN( u0_u3_u5_n191 ) );
  AOI22_X1 u0_u3_u5_U40 (.B2( u0_u3_u5_n131 ) , .A2( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n169 ) , .B1( u0_u3_u5_n174 ) , .A1( u0_u3_u5_n185 ) );
  NOR2_X1 u0_u3_u5_U41 (.A1( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n150 ) , .A2( u0_u3_u5_n173 ) );
  AOI21_X1 u0_u3_u5_U42 (.A( u0_u3_u5_n118 ) , .B2( u0_u3_u5_n145 ) , .ZN( u0_u3_u5_n168 ) , .B1( u0_u3_u5_n186 ) );
  INV_X1 u0_u3_u5_U43 (.A( u0_u3_u5_n122 ) , .ZN( u0_u3_u5_n186 ) );
  NOR2_X1 u0_u3_u5_U44 (.A1( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n152 ) , .A2( u0_u3_u5_n176 ) );
  NOR2_X1 u0_u3_u5_U45 (.A1( u0_u3_u5_n115 ) , .ZN( u0_u3_u5_n118 ) , .A2( u0_u3_u5_n153 ) );
  NOR2_X1 u0_u3_u5_U46 (.A2( u0_u3_u5_n145 ) , .ZN( u0_u3_u5_n156 ) , .A1( u0_u3_u5_n174 ) );
  NOR2_X1 u0_u3_u5_U47 (.ZN( u0_u3_u5_n121 ) , .A2( u0_u3_u5_n145 ) , .A1( u0_u3_u5_n176 ) );
  AOI22_X1 u0_u3_u5_U48 (.ZN( u0_u3_u5_n114 ) , .A2( u0_u3_u5_n137 ) , .A1( u0_u3_u5_n145 ) , .B2( u0_u3_u5_n175 ) , .B1( u0_u3_u5_n193 ) );
  OAI211_X1 u0_u3_u5_U49 (.B( u0_u3_u5_n124 ) , .A( u0_u3_u5_n125 ) , .C2( u0_u3_u5_n126 ) , .C1( u0_u3_u5_n127 ) , .ZN( u0_u3_u5_n128 ) );
  OAI21_X1 u0_u3_u5_U5 (.B2( u0_u3_u5_n136 ) , .B1( u0_u3_u5_n137 ) , .ZN( u0_u3_u5_n138 ) , .A( u0_u3_u5_n177 ) );
  NOR3_X1 u0_u3_u5_U50 (.ZN( u0_u3_u5_n127 ) , .A1( u0_u3_u5_n136 ) , .A3( u0_u3_u5_n148 ) , .A2( u0_u3_u5_n182 ) );
  OAI21_X1 u0_u3_u5_U51 (.ZN( u0_u3_u5_n124 ) , .A( u0_u3_u5_n177 ) , .B2( u0_u3_u5_n183 ) , .B1( u0_u3_u5_n189 ) );
  OAI21_X1 u0_u3_u5_U52 (.ZN( u0_u3_u5_n125 ) , .A( u0_u3_u5_n174 ) , .B2( u0_u3_u5_n185 ) , .B1( u0_u3_u5_n190 ) );
  AOI21_X1 u0_u3_u5_U53 (.A( u0_u3_u5_n153 ) , .B2( u0_u3_u5_n154 ) , .B1( u0_u3_u5_n155 ) , .ZN( u0_u3_u5_n164 ) );
  AOI21_X1 u0_u3_u5_U54 (.ZN( u0_u3_u5_n110 ) , .B1( u0_u3_u5_n122 ) , .B2( u0_u3_u5_n139 ) , .A( u0_u3_u5_n153 ) );
  INV_X1 u0_u3_u5_U55 (.A( u0_u3_u5_n153 ) , .ZN( u0_u3_u5_n176 ) );
  INV_X1 u0_u3_u5_U56 (.A( u0_u3_u5_n126 ) , .ZN( u0_u3_u5_n173 ) );
  AND2_X1 u0_u3_u5_U57 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n147 ) );
  AND2_X1 u0_u3_u5_U58 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n148 ) );
  NAND2_X1 u0_u3_u5_U59 (.A1( u0_u3_u5_n105 ) , .A2( u0_u3_u5_n106 ) , .ZN( u0_u3_u5_n158 ) );
  INV_X1 u0_u3_u5_U6 (.A( u0_u3_u5_n135 ) , .ZN( u0_u3_u5_n178 ) );
  NAND2_X1 u0_u3_u5_U60 (.A2( u0_u3_u5_n108 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n139 ) );
  NAND2_X1 u0_u3_u5_U61 (.A1( u0_u3_u5_n106 ) , .A2( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n119 ) );
  NAND2_X1 u0_u3_u5_U62 (.A2( u0_u3_u5_n103 ) , .A1( u0_u3_u5_n105 ) , .ZN( u0_u3_u5_n140 ) );
  NAND2_X1 u0_u3_u5_U63 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n105 ) , .ZN( u0_u3_u5_n155 ) );
  NAND2_X1 u0_u3_u5_U64 (.A2( u0_u3_u5_n106 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n122 ) );
  NAND2_X1 u0_u3_u5_U65 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n106 ) , .ZN( u0_u3_u5_n115 ) );
  NAND2_X1 u0_u3_u5_U66 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n103 ) , .ZN( u0_u3_u5_n161 ) );
  NAND2_X1 u0_u3_u5_U67 (.A1( u0_u3_u5_n105 ) , .A2( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n154 ) );
  INV_X1 u0_u3_u5_U68 (.A( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n172 ) );
  NAND2_X1 u0_u3_u5_U69 (.A1( u0_u3_u5_n103 ) , .A2( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n123 ) );
  OAI22_X1 u0_u3_u5_U7 (.B2( u0_u3_u5_n149 ) , .B1( u0_u3_u5_n150 ) , .A2( u0_u3_u5_n151 ) , .A1( u0_u3_u5_n152 ) , .ZN( u0_u3_u5_n165 ) );
  NAND2_X1 u0_u3_u5_U70 (.A2( u0_u3_u5_n103 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n151 ) );
  NAND2_X1 u0_u3_u5_U71 (.A2( u0_u3_u5_n107 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n120 ) );
  NAND2_X1 u0_u3_u5_U72 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n157 ) );
  AND2_X1 u0_u3_u5_U73 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n104 ) , .ZN( u0_u3_u5_n131 ) );
  INV_X1 u0_u3_u5_U74 (.A( u0_u3_u5_n102 ) , .ZN( u0_u3_u5_n195 ) );
  OAI221_X1 u0_u3_u5_U75 (.A( u0_u3_u5_n101 ) , .ZN( u0_u3_u5_n102 ) , .C2( u0_u3_u5_n115 ) , .C1( u0_u3_u5_n126 ) , .B1( u0_u3_u5_n134 ) , .B2( u0_u3_u5_n160 ) );
  OAI21_X1 u0_u3_u5_U76 (.ZN( u0_u3_u5_n101 ) , .B1( u0_u3_u5_n137 ) , .A( u0_u3_u5_n146 ) , .B2( u0_u3_u5_n147 ) );
  NOR2_X1 u0_u3_u5_U77 (.A2( u0_u3_X_34 ) , .A1( u0_u3_X_35 ) , .ZN( u0_u3_u5_n145 ) );
  NOR2_X1 u0_u3_u5_U78 (.A2( u0_u3_X_34 ) , .ZN( u0_u3_u5_n146 ) , .A1( u0_u3_u5_n171 ) );
  NOR2_X1 u0_u3_u5_U79 (.A2( u0_u3_X_31 ) , .A1( u0_u3_X_32 ) , .ZN( u0_u3_u5_n103 ) );
  NOR3_X1 u0_u3_u5_U8 (.A2( u0_u3_u5_n147 ) , .A1( u0_u3_u5_n148 ) , .ZN( u0_u3_u5_n149 ) , .A3( u0_u3_u5_n194 ) );
  NOR2_X1 u0_u3_u5_U80 (.A2( u0_u3_X_36 ) , .ZN( u0_u3_u5_n105 ) , .A1( u0_u3_u5_n180 ) );
  NOR2_X1 u0_u3_u5_U81 (.A2( u0_u3_X_33 ) , .ZN( u0_u3_u5_n108 ) , .A1( u0_u3_u5_n170 ) );
  NOR2_X1 u0_u3_u5_U82 (.A2( u0_u3_X_33 ) , .A1( u0_u3_X_36 ) , .ZN( u0_u3_u5_n107 ) );
  NOR2_X1 u0_u3_u5_U83 (.A2( u0_u3_X_31 ) , .ZN( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n181 ) );
  NAND2_X1 u0_u3_u5_U84 (.A2( u0_u3_X_34 ) , .A1( u0_u3_X_35 ) , .ZN( u0_u3_u5_n153 ) );
  NAND2_X1 u0_u3_u5_U85 (.A1( u0_u3_X_34 ) , .ZN( u0_u3_u5_n126 ) , .A2( u0_u3_u5_n171 ) );
  AND2_X1 u0_u3_u5_U86 (.A1( u0_u3_X_31 ) , .A2( u0_u3_X_32 ) , .ZN( u0_u3_u5_n106 ) );
  AND2_X1 u0_u3_u5_U87 (.A1( u0_u3_X_31 ) , .ZN( u0_u3_u5_n109 ) , .A2( u0_u3_u5_n181 ) );
  INV_X1 u0_u3_u5_U88 (.A( u0_u3_X_33 ) , .ZN( u0_u3_u5_n180 ) );
  INV_X1 u0_u3_u5_U89 (.A( u0_u3_X_35 ) , .ZN( u0_u3_u5_n171 ) );
  NOR2_X1 u0_u3_u5_U9 (.ZN( u0_u3_u5_n135 ) , .A1( u0_u3_u5_n173 ) , .A2( u0_u3_u5_n176 ) );
  INV_X1 u0_u3_u5_U90 (.A( u0_u3_X_36 ) , .ZN( u0_u3_u5_n170 ) );
  INV_X1 u0_u3_u5_U91 (.A( u0_u3_X_32 ) , .ZN( u0_u3_u5_n181 ) );
  NAND4_X1 u0_u3_u5_U92 (.ZN( u0_out3_29 ) , .A4( u0_u3_u5_n129 ) , .A3( u0_u3_u5_n130 ) , .A2( u0_u3_u5_n168 ) , .A1( u0_u3_u5_n196 ) );
  AOI221_X1 u0_u3_u5_U93 (.A( u0_u3_u5_n128 ) , .ZN( u0_u3_u5_n129 ) , .C2( u0_u3_u5_n132 ) , .B2( u0_u3_u5_n159 ) , .B1( u0_u3_u5_n176 ) , .C1( u0_u3_u5_n184 ) );
  AOI222_X1 u0_u3_u5_U94 (.ZN( u0_u3_u5_n130 ) , .A2( u0_u3_u5_n146 ) , .B1( u0_u3_u5_n147 ) , .C2( u0_u3_u5_n175 ) , .B2( u0_u3_u5_n179 ) , .A1( u0_u3_u5_n188 ) , .C1( u0_u3_u5_n194 ) );
  NAND4_X1 u0_u3_u5_U95 (.ZN( u0_out3_19 ) , .A4( u0_u3_u5_n166 ) , .A3( u0_u3_u5_n167 ) , .A2( u0_u3_u5_n168 ) , .A1( u0_u3_u5_n169 ) );
  AOI22_X1 u0_u3_u5_U96 (.B2( u0_u3_u5_n145 ) , .A2( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n167 ) , .B1( u0_u3_u5_n182 ) , .A1( u0_u3_u5_n189 ) );
  NOR4_X1 u0_u3_u5_U97 (.A4( u0_u3_u5_n162 ) , .A3( u0_u3_u5_n163 ) , .A2( u0_u3_u5_n164 ) , .A1( u0_u3_u5_n165 ) , .ZN( u0_u3_u5_n166 ) );
  NAND4_X1 u0_u3_u5_U98 (.ZN( u0_out3_11 ) , .A4( u0_u3_u5_n143 ) , .A3( u0_u3_u5_n144 ) , .A2( u0_u3_u5_n169 ) , .A1( u0_u3_u5_n196 ) );
  AOI22_X1 u0_u3_u5_U99 (.A2( u0_u3_u5_n132 ) , .ZN( u0_u3_u5_n144 ) , .B2( u0_u3_u5_n145 ) , .B1( u0_u3_u5_n184 ) , .A1( u0_u3_u5_n194 ) );
  XOR2_X1 u0_u5_U13 (.B( u0_K6_42 ) , .A( u0_R4_29 ) , .Z( u0_u5_X_42 ) );
  XOR2_X1 u0_u5_U14 (.B( u0_K6_41 ) , .A( u0_R4_28 ) , .Z( u0_u5_X_41 ) );
  XOR2_X1 u0_u5_U15 (.B( u0_K6_40 ) , .A( u0_R4_27 ) , .Z( u0_u5_X_40 ) );
  XOR2_X1 u0_u5_U17 (.B( u0_K6_39 ) , .A( u0_R4_26 ) , .Z( u0_u5_X_39 ) );
  XOR2_X1 u0_u5_U18 (.B( u0_K6_38 ) , .A( u0_R4_25 ) , .Z( u0_u5_X_38 ) );
  XOR2_X1 u0_u5_U19 (.B( u0_K6_37 ) , .A( u0_R4_24 ) , .Z( u0_u5_X_37 ) );
  XOR2_X1 u0_u5_U20 (.B( u0_K6_36 ) , .A( u0_R4_25 ) , .Z( u0_u5_X_36 ) );
  XOR2_X1 u0_u5_U21 (.B( u0_K6_35 ) , .A( u0_R4_24 ) , .Z( u0_u5_X_35 ) );
  XOR2_X1 u0_u5_U22 (.B( u0_K6_34 ) , .A( u0_R4_23 ) , .Z( u0_u5_X_34 ) );
  XOR2_X1 u0_u5_U23 (.B( u0_K6_33 ) , .A( u0_R4_22 ) , .Z( u0_u5_X_33 ) );
  XOR2_X1 u0_u5_U24 (.B( u0_K6_32 ) , .A( u0_R4_21 ) , .Z( u0_u5_X_32 ) );
  XOR2_X1 u0_u5_U25 (.B( u0_K6_31 ) , .A( u0_R4_20 ) , .Z( u0_u5_X_31 ) );
  XOR2_X1 u0_u5_U26 (.B( u0_K6_30 ) , .A( u0_R4_21 ) , .Z( u0_u5_X_30 ) );
  XOR2_X1 u0_u5_U28 (.B( u0_K6_29 ) , .A( u0_R4_20 ) , .Z( u0_u5_X_29 ) );
  XOR2_X1 u0_u5_U29 (.B( u0_K6_28 ) , .A( u0_R4_19 ) , .Z( u0_u5_X_28 ) );
  XOR2_X1 u0_u5_U30 (.B( u0_K6_27 ) , .A( u0_R4_18 ) , .Z( u0_u5_X_27 ) );
  XOR2_X1 u0_u5_U31 (.B( u0_K6_26 ) , .A( u0_R4_17 ) , .Z( u0_u5_X_26 ) );
  XOR2_X1 u0_u5_U32 (.B( u0_K6_25 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_25 ) );
  XOR2_X1 u0_u5_U33 (.B( u0_K6_24 ) , .A( u0_R4_17 ) , .Z( u0_u5_X_24 ) );
  XOR2_X1 u0_u5_U34 (.B( u0_K6_23 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_23 ) );
  XOR2_X1 u0_u5_U35 (.B( u0_K6_22 ) , .A( u0_R4_15 ) , .Z( u0_u5_X_22 ) );
  XOR2_X1 u0_u5_U36 (.B( u0_K6_21 ) , .A( u0_R4_14 ) , .Z( u0_u5_X_21 ) );
  XOR2_X1 u0_u5_U37 (.B( u0_K6_20 ) , .A( u0_R4_13 ) , .Z( u0_u5_X_20 ) );
  XOR2_X1 u0_u5_U39 (.B( u0_K6_19 ) , .A( u0_R4_12 ) , .Z( u0_u5_X_19 ) );
  OAI22_X1 u0_u5_u3_U10 (.B1( u0_u5_u3_n113 ) , .A2( u0_u5_u3_n135 ) , .A1( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n164 ) , .ZN( u0_u5_u3_n98 ) );
  OAI211_X1 u0_u5_u3_U11 (.B( u0_u5_u3_n106 ) , .ZN( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n128 ) , .C1( u0_u5_u3_n167 ) , .A( u0_u5_u3_n181 ) );
  AOI221_X1 u0_u5_u3_U12 (.C1( u0_u5_u3_n105 ) , .ZN( u0_u5_u3_n106 ) , .A( u0_u5_u3_n131 ) , .B2( u0_u5_u3_n132 ) , .C2( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n169 ) );
  INV_X1 u0_u5_u3_U13 (.ZN( u0_u5_u3_n181 ) , .A( u0_u5_u3_n98 ) );
  NAND2_X1 u0_u5_u3_U14 (.ZN( u0_u5_u3_n105 ) , .A2( u0_u5_u3_n130 ) , .A1( u0_u5_u3_n155 ) );
  AOI22_X1 u0_u5_u3_U15 (.B1( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n116 ) , .ZN( u0_u5_u3_n123 ) , .B2( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U16 (.ZN( u0_u5_u3_n116 ) , .A2( u0_u5_u3_n151 ) , .A1( u0_u5_u3_n182 ) );
  NOR2_X1 u0_u5_u3_U17 (.ZN( u0_u5_u3_n126 ) , .A2( u0_u5_u3_n150 ) , .A1( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U18 (.ZN( u0_u5_u3_n112 ) , .B2( u0_u5_u3_n146 ) , .B1( u0_u5_u3_n155 ) , .A( u0_u5_u3_n167 ) );
  NAND2_X1 u0_u5_u3_U19 (.A1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n142 ) , .A2( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U20 (.ZN( u0_u5_u3_n132 ) , .A2( u0_u5_u3_n152 ) , .A1( u0_u5_u3_n156 ) );
  AND2_X1 u0_u5_u3_U21 (.A2( u0_u5_u3_n113 ) , .A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n151 ) );
  INV_X1 u0_u5_u3_U22 (.A( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n165 ) );
  INV_X1 u0_u5_u3_U23 (.A( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n170 ) );
  NAND2_X1 u0_u5_u3_U24 (.A1( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .ZN( u0_u5_u3_n140 ) );
  NAND2_X1 u0_u5_u3_U25 (.ZN( u0_u5_u3_n117 ) , .A1( u0_u5_u3_n124 ) , .A2( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U26 (.ZN( u0_u5_u3_n143 ) , .A1( u0_u5_u3_n165 ) , .A2( u0_u5_u3_n167 ) );
  INV_X1 u0_u5_u3_U27 (.A( u0_u5_u3_n130 ) , .ZN( u0_u5_u3_n177 ) );
  INV_X1 u0_u5_u3_U28 (.A( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n176 ) );
  INV_X1 u0_u5_u3_U29 (.A( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n174 ) );
  INV_X1 u0_u5_u3_U3 (.A( u0_u5_u3_n129 ) , .ZN( u0_u5_u3_n183 ) );
  INV_X1 u0_u5_u3_U30 (.A( u0_u5_u3_n139 ) , .ZN( u0_u5_u3_n185 ) );
  NOR2_X1 u0_u5_u3_U31 (.ZN( u0_u5_u3_n135 ) , .A2( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n169 ) );
  OAI222_X1 u0_u5_u3_U32 (.C2( u0_u5_u3_n107 ) , .A2( u0_u5_u3_n108 ) , .B1( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n138 ) , .B2( u0_u5_u3_n146 ) , .C1( u0_u5_u3_n154 ) , .A1( u0_u5_u3_n164 ) );
  NOR4_X1 u0_u5_u3_U33 (.A4( u0_u5_u3_n157 ) , .A3( u0_u5_u3_n158 ) , .A2( u0_u5_u3_n159 ) , .A1( u0_u5_u3_n160 ) , .ZN( u0_u5_u3_n161 ) );
  AOI21_X1 u0_u5_u3_U34 (.B2( u0_u5_u3_n152 ) , .B1( u0_u5_u3_n153 ) , .ZN( u0_u5_u3_n158 ) , .A( u0_u5_u3_n164 ) );
  AOI21_X1 u0_u5_u3_U35 (.A( u0_u5_u3_n154 ) , .B2( u0_u5_u3_n155 ) , .B1( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n157 ) );
  AOI21_X1 u0_u5_u3_U36 (.A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n150 ) , .B1( u0_u5_u3_n151 ) , .ZN( u0_u5_u3_n159 ) );
  AOI211_X1 u0_u5_u3_U37 (.ZN( u0_u5_u3_n109 ) , .A( u0_u5_u3_n119 ) , .C2( u0_u5_u3_n129 ) , .B( u0_u5_u3_n138 ) , .C1( u0_u5_u3_n141 ) );
  AOI211_X1 u0_u5_u3_U38 (.B( u0_u5_u3_n119 ) , .A( u0_u5_u3_n120 ) , .C2( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n122 ) , .C1( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U39 (.A( u0_u5_u3_n156 ) , .ZN( u0_u5_u3_n179 ) );
  INV_X1 u0_u5_u3_U4 (.A( u0_u5_u3_n140 ) , .ZN( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u3_U40 (.B1( u0_u5_u3_n118 ) , .ZN( u0_u5_u3_n120 ) , .A1( u0_u5_u3_n135 ) , .B2( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n178 ) );
  AND3_X1 u0_u5_u3_U41 (.ZN( u0_u5_u3_n118 ) , .A2( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n144 ) , .A3( u0_u5_u3_n152 ) );
  INV_X1 u0_u5_u3_U42 (.A( u0_u5_u3_n121 ) , .ZN( u0_u5_u3_n164 ) );
  NAND2_X1 u0_u5_u3_U43 (.ZN( u0_u5_u3_n133 ) , .A1( u0_u5_u3_n154 ) , .A2( u0_u5_u3_n164 ) );
  OAI211_X1 u0_u5_u3_U44 (.B( u0_u5_u3_n127 ) , .ZN( u0_u5_u3_n139 ) , .C1( u0_u5_u3_n150 ) , .C2( u0_u5_u3_n154 ) , .A( u0_u5_u3_n184 ) );
  INV_X1 u0_u5_u3_U45 (.A( u0_u5_u3_n125 ) , .ZN( u0_u5_u3_n184 ) );
  AOI221_X1 u0_u5_u3_U46 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n127 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n169 ) , .B2( u0_u5_u3_n170 ) , .B1( u0_u5_u3_n174 ) );
  OAI22_X1 u0_u5_u3_U47 (.A1( u0_u5_u3_n124 ) , .ZN( u0_u5_u3_n125 ) , .B2( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n165 ) , .B1( u0_u5_u3_n167 ) );
  NOR2_X1 u0_u5_u3_U48 (.A1( u0_u5_u3_n113 ) , .ZN( u0_u5_u3_n131 ) , .A2( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U49 (.A1( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n150 ) , .A2( u0_u5_u3_n99 ) );
  INV_X1 u0_u5_u3_U5 (.A( u0_u5_u3_n117 ) , .ZN( u0_u5_u3_n178 ) );
  NAND2_X1 u0_u5_u3_U50 (.A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n155 ) , .A1( u0_u5_u3_n97 ) );
  INV_X1 u0_u5_u3_U51 (.A( u0_u5_u3_n141 ) , .ZN( u0_u5_u3_n167 ) );
  AOI21_X1 u0_u5_u3_U52 (.B2( u0_u5_u3_n114 ) , .B1( u0_u5_u3_n146 ) , .A( u0_u5_u3_n154 ) , .ZN( u0_u5_u3_n94 ) );
  AOI21_X1 u0_u5_u3_U53 (.ZN( u0_u5_u3_n110 ) , .B2( u0_u5_u3_n142 ) , .B1( u0_u5_u3_n186 ) , .A( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U54 (.A( u0_u5_u3_n145 ) , .ZN( u0_u5_u3_n186 ) );
  AOI21_X1 u0_u5_u3_U55 (.B1( u0_u5_u3_n124 ) , .A( u0_u5_u3_n149 ) , .B2( u0_u5_u3_n155 ) , .ZN( u0_u5_u3_n95 ) );
  INV_X1 u0_u5_u3_U56 (.A( u0_u5_u3_n149 ) , .ZN( u0_u5_u3_n169 ) );
  NAND2_X1 u0_u5_u3_U57 (.ZN( u0_u5_u3_n124 ) , .A1( u0_u5_u3_n96 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U58 (.A2( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n146 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U59 (.A1( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n145 ) , .A2( u0_u5_u3_n99 ) );
  AOI221_X1 u0_u5_u3_U6 (.A( u0_u5_u3_n131 ) , .C2( u0_u5_u3_n132 ) , .C1( u0_u5_u3_n133 ) , .ZN( u0_u5_u3_n134 ) , .B1( u0_u5_u3_n143 ) , .B2( u0_u5_u3_n177 ) );
  NAND2_X1 u0_u5_u3_U60 (.A1( u0_u5_u3_n100 ) , .ZN( u0_u5_u3_n156 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U61 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n148 ) );
  NAND2_X1 u0_u5_u3_U62 (.A1( u0_u5_u3_n100 ) , .A2( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n128 ) );
  NAND2_X1 u0_u5_u3_U63 (.A2( u0_u5_u3_n101 ) , .A1( u0_u5_u3_n102 ) , .ZN( u0_u5_u3_n152 ) );
  NAND2_X1 u0_u5_u3_U64 (.A2( u0_u5_u3_n101 ) , .ZN( u0_u5_u3_n114 ) , .A1( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U65 (.ZN( u0_u5_u3_n107 ) , .A1( u0_u5_u3_n97 ) , .A2( u0_u5_u3_n99 ) );
  NAND2_X1 u0_u5_u3_U66 (.A2( u0_u5_u3_n100 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n113 ) );
  NAND2_X1 u0_u5_u3_U67 (.A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n153 ) , .A2( u0_u5_u3_n97 ) );
  NAND2_X1 u0_u5_u3_U68 (.A2( u0_u5_u3_n103 ) , .A1( u0_u5_u3_n104 ) , .ZN( u0_u5_u3_n130 ) );
  NAND2_X1 u0_u5_u3_U69 (.A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n96 ) );
  OAI22_X1 u0_u5_u3_U7 (.B2( u0_u5_u3_n147 ) , .A2( u0_u5_u3_n148 ) , .ZN( u0_u5_u3_n160 ) , .B1( u0_u5_u3_n165 ) , .A1( u0_u5_u3_n168 ) );
  NAND2_X1 u0_u5_u3_U70 (.A1( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n103 ) , .ZN( u0_u5_u3_n108 ) );
  NOR2_X1 u0_u5_u3_U71 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n99 ) );
  NOR2_X1 u0_u5_u3_U72 (.A2( u0_u5_X_21 ) , .A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n103 ) );
  NOR2_X1 u0_u5_u3_U73 (.A2( u0_u5_X_24 ) , .A1( u0_u5_u3_n171 ) , .ZN( u0_u5_u3_n97 ) );
  NOR2_X1 u0_u5_u3_U74 (.A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n141 ) , .A1( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U75 (.A2( u0_u5_X_19 ) , .A1( u0_u5_u3_n172 ) , .ZN( u0_u5_u3_n96 ) );
  NAND2_X1 u0_u5_u3_U76 (.A1( u0_u5_X_22 ) , .A2( u0_u5_X_23 ) , .ZN( u0_u5_u3_n154 ) );
  NAND2_X1 u0_u5_u3_U77 (.A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n149 ) , .A2( u0_u5_u3_n166 ) );
  NOR2_X1 u0_u5_u3_U78 (.A2( u0_u5_X_22 ) , .A1( u0_u5_X_23 ) , .ZN( u0_u5_u3_n121 ) );
  AND2_X1 u0_u5_u3_U79 (.A1( u0_u5_X_24 ) , .ZN( u0_u5_u3_n101 ) , .A2( u0_u5_u3_n171 ) );
  AND3_X1 u0_u5_u3_U8 (.A3( u0_u5_u3_n144 ) , .A2( u0_u5_u3_n145 ) , .A1( u0_u5_u3_n146 ) , .ZN( u0_u5_u3_n147 ) );
  AND2_X1 u0_u5_u3_U80 (.A1( u0_u5_X_19 ) , .ZN( u0_u5_u3_n102 ) , .A2( u0_u5_u3_n172 ) );
  AND2_X1 u0_u5_u3_U81 (.A1( u0_u5_X_21 ) , .A2( u0_u5_X_24 ) , .ZN( u0_u5_u3_n100 ) );
  AND2_X1 u0_u5_u3_U82 (.A2( u0_u5_X_19 ) , .A1( u0_u5_X_20 ) , .ZN( u0_u5_u3_n104 ) );
  INV_X1 u0_u5_u3_U83 (.A( u0_u5_X_22 ) , .ZN( u0_u5_u3_n166 ) );
  INV_X1 u0_u5_u3_U84 (.A( u0_u5_X_21 ) , .ZN( u0_u5_u3_n171 ) );
  INV_X1 u0_u5_u3_U85 (.A( u0_u5_X_20 ) , .ZN( u0_u5_u3_n172 ) );
  NAND4_X1 u0_u5_u3_U86 (.ZN( u0_out5_26 ) , .A4( u0_u5_u3_n109 ) , .A3( u0_u5_u3_n110 ) , .A2( u0_u5_u3_n111 ) , .A1( u0_u5_u3_n173 ) );
  INV_X1 u0_u5_u3_U87 (.ZN( u0_u5_u3_n173 ) , .A( u0_u5_u3_n94 ) );
  OAI21_X1 u0_u5_u3_U88 (.ZN( u0_u5_u3_n111 ) , .B2( u0_u5_u3_n117 ) , .A( u0_u5_u3_n133 ) , .B1( u0_u5_u3_n176 ) );
  NAND4_X1 u0_u5_u3_U89 (.ZN( u0_out5_20 ) , .A4( u0_u5_u3_n122 ) , .A3( u0_u5_u3_n123 ) , .A1( u0_u5_u3_n175 ) , .A2( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U9 (.A( u0_u5_u3_n143 ) , .ZN( u0_u5_u3_n168 ) );
  INV_X1 u0_u5_u3_U90 (.A( u0_u5_u3_n126 ) , .ZN( u0_u5_u3_n180 ) );
  INV_X1 u0_u5_u3_U91 (.A( u0_u5_u3_n112 ) , .ZN( u0_u5_u3_n175 ) );
  NAND4_X1 u0_u5_u3_U92 (.ZN( u0_out5_1 ) , .A4( u0_u5_u3_n161 ) , .A3( u0_u5_u3_n162 ) , .A2( u0_u5_u3_n163 ) , .A1( u0_u5_u3_n185 ) );
  NAND2_X1 u0_u5_u3_U93 (.ZN( u0_u5_u3_n163 ) , .A2( u0_u5_u3_n170 ) , .A1( u0_u5_u3_n176 ) );
  AOI22_X1 u0_u5_u3_U94 (.B2( u0_u5_u3_n140 ) , .B1( u0_u5_u3_n141 ) , .A2( u0_u5_u3_n142 ) , .ZN( u0_u5_u3_n162 ) , .A1( u0_u5_u3_n177 ) );
  OR4_X1 u0_u5_u3_U95 (.ZN( u0_out5_10 ) , .A4( u0_u5_u3_n136 ) , .A3( u0_u5_u3_n137 ) , .A1( u0_u5_u3_n138 ) , .A2( u0_u5_u3_n139 ) );
  OAI222_X1 u0_u5_u3_U96 (.C1( u0_u5_u3_n128 ) , .ZN( u0_u5_u3_n137 ) , .B1( u0_u5_u3_n148 ) , .A2( u0_u5_u3_n150 ) , .B2( u0_u5_u3_n154 ) , .C2( u0_u5_u3_n164 ) , .A1( u0_u5_u3_n167 ) );
  OAI221_X1 u0_u5_u3_U97 (.A( u0_u5_u3_n134 ) , .B2( u0_u5_u3_n135 ) , .ZN( u0_u5_u3_n136 ) , .C1( u0_u5_u3_n149 ) , .B1( u0_u5_u3_n151 ) , .C2( u0_u5_u3_n183 ) );
  NAND3_X1 u0_u5_u3_U98 (.A1( u0_u5_u3_n114 ) , .ZN( u0_u5_u3_n115 ) , .A2( u0_u5_u3_n145 ) , .A3( u0_u5_u3_n153 ) );
  NAND3_X1 u0_u5_u3_U99 (.ZN( u0_u5_u3_n129 ) , .A2( u0_u5_u3_n144 ) , .A1( u0_u5_u3_n153 ) , .A3( u0_u5_u3_n182 ) );
  OAI22_X1 u0_u5_u4_U10 (.B2( u0_u5_u4_n135 ) , .ZN( u0_u5_u4_n137 ) , .B1( u0_u5_u4_n153 ) , .A1( u0_u5_u4_n155 ) , .A2( u0_u5_u4_n171 ) );
  AND3_X1 u0_u5_u4_U11 (.A2( u0_u5_u4_n134 ) , .ZN( u0_u5_u4_n135 ) , .A3( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n157 ) );
  NAND2_X1 u0_u5_u4_U12 (.ZN( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n173 ) );
  AOI21_X1 u0_u5_u4_U13 (.B2( u0_u5_u4_n160 ) , .B1( u0_u5_u4_n161 ) , .ZN( u0_u5_u4_n162 ) , .A( u0_u5_u4_n170 ) );
  AOI21_X1 u0_u5_u4_U14 (.ZN( u0_u5_u4_n107 ) , .B2( u0_u5_u4_n143 ) , .A( u0_u5_u4_n174 ) , .B1( u0_u5_u4_n184 ) );
  AOI21_X1 u0_u5_u4_U15 (.B2( u0_u5_u4_n158 ) , .B1( u0_u5_u4_n159 ) , .ZN( u0_u5_u4_n163 ) , .A( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U16 (.A( u0_u5_u4_n153 ) , .B2( u0_u5_u4_n154 ) , .B1( u0_u5_u4_n155 ) , .ZN( u0_u5_u4_n165 ) );
  AOI21_X1 u0_u5_u4_U17 (.A( u0_u5_u4_n156 ) , .B2( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n164 ) , .B1( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U18 (.A( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n170 ) );
  AND2_X1 u0_u5_u4_U19 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n155 ) , .A1( u0_u5_u4_n160 ) );
  INV_X1 u0_u5_u4_U20 (.A( u0_u5_u4_n156 ) , .ZN( u0_u5_u4_n175 ) );
  NAND2_X1 u0_u5_u4_U21 (.A2( u0_u5_u4_n118 ) , .ZN( u0_u5_u4_n131 ) , .A1( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U22 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n130 ) );
  NAND2_X1 u0_u5_u4_U23 (.ZN( u0_u5_u4_n117 ) , .A2( u0_u5_u4_n118 ) , .A1( u0_u5_u4_n148 ) );
  NAND2_X1 u0_u5_u4_U24 (.ZN( u0_u5_u4_n129 ) , .A1( u0_u5_u4_n134 ) , .A2( u0_u5_u4_n148 ) );
  AND3_X1 u0_u5_u4_U25 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n143 ) , .A3( u0_u5_u4_n154 ) , .ZN( u0_u5_u4_n161 ) );
  AND2_X1 u0_u5_u4_U26 (.A1( u0_u5_u4_n145 ) , .A2( u0_u5_u4_n147 ) , .ZN( u0_u5_u4_n159 ) );
  OR3_X1 u0_u5_u4_U27 (.A3( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n115 ) , .A1( u0_u5_u4_n116 ) , .ZN( u0_u5_u4_n136 ) );
  AOI21_X1 u0_u5_u4_U28 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n116 ) , .B2( u0_u5_u4_n173 ) , .B1( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U29 (.ZN( u0_u5_u4_n115 ) , .B2( u0_u5_u4_n145 ) , .B1( u0_u5_u4_n146 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U3 (.ZN( u0_u5_u4_n121 ) , .A1( u0_u5_u4_n181 ) , .A2( u0_u5_u4_n182 ) );
  OAI22_X1 u0_u5_u4_U30 (.ZN( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n121 ) , .B1( u0_u5_u4_n160 ) , .B2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n171 ) );
  INV_X1 u0_u5_u4_U31 (.A( u0_u5_u4_n158 ) , .ZN( u0_u5_u4_n182 ) );
  INV_X1 u0_u5_u4_U32 (.ZN( u0_u5_u4_n181 ) , .A( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U33 (.A( u0_u5_u4_n144 ) , .ZN( u0_u5_u4_n179 ) );
  INV_X1 u0_u5_u4_U34 (.A( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n178 ) );
  NAND2_X1 u0_u5_u4_U35 (.A2( u0_u5_u4_n154 ) , .A1( u0_u5_u4_n96 ) , .ZN( u0_u5_u4_n97 ) );
  INV_X1 u0_u5_u4_U36 (.ZN( u0_u5_u4_n186 ) , .A( u0_u5_u4_n95 ) );
  OAI221_X1 u0_u5_u4_U37 (.C1( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n158 ) , .B2( u0_u5_u4_n171 ) , .C2( u0_u5_u4_n173 ) , .A( u0_u5_u4_n94 ) , .ZN( u0_u5_u4_n95 ) );
  AOI222_X1 u0_u5_u4_U38 (.B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n138 ) , .C2( u0_u5_u4_n175 ) , .A2( u0_u5_u4_n179 ) , .C1( u0_u5_u4_n181 ) , .B1( u0_u5_u4_n185 ) , .ZN( u0_u5_u4_n94 ) );
  INV_X1 u0_u5_u4_U39 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n185 ) );
  INV_X1 u0_u5_u4_U4 (.A( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U40 (.A( u0_u5_u4_n143 ) , .ZN( u0_u5_u4_n183 ) );
  NOR2_X1 u0_u5_u4_U41 (.ZN( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n168 ) , .A2( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U42 (.A1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n153 ) );
  NOR2_X1 u0_u5_u4_U43 (.A2( u0_u5_u4_n128 ) , .A1( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n156 ) );
  AOI22_X1 u0_u5_u4_U44 (.B2( u0_u5_u4_n122 ) , .A1( u0_u5_u4_n123 ) , .ZN( u0_u5_u4_n124 ) , .B1( u0_u5_u4_n128 ) , .A2( u0_u5_u4_n172 ) );
  INV_X1 u0_u5_u4_U45 (.A( u0_u5_u4_n153 ) , .ZN( u0_u5_u4_n172 ) );
  NAND2_X1 u0_u5_u4_U46 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n123 ) , .A1( u0_u5_u4_n161 ) );
  AOI22_X1 u0_u5_u4_U47 (.B2( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n133 ) , .ZN( u0_u5_u4_n140 ) , .A1( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n179 ) );
  NAND2_X1 u0_u5_u4_U48 (.ZN( u0_u5_u4_n133 ) , .A2( u0_u5_u4_n146 ) , .A1( u0_u5_u4_n154 ) );
  NAND2_X1 u0_u5_u4_U49 (.A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n154 ) , .A2( u0_u5_u4_n98 ) );
  NOR4_X1 u0_u5_u4_U5 (.A4( u0_u5_u4_n106 ) , .A3( u0_u5_u4_n107 ) , .A2( u0_u5_u4_n108 ) , .A1( u0_u5_u4_n109 ) , .ZN( u0_u5_u4_n110 ) );
  NAND2_X1 u0_u5_u4_U50 (.A1( u0_u5_u4_n101 ) , .ZN( u0_u5_u4_n158 ) , .A2( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U51 (.ZN( u0_u5_u4_n127 ) , .A( u0_u5_u4_n136 ) , .B2( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n180 ) );
  INV_X1 u0_u5_u4_U52 (.A( u0_u5_u4_n160 ) , .ZN( u0_u5_u4_n180 ) );
  NAND2_X1 u0_u5_u4_U53 (.A2( u0_u5_u4_n104 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n146 ) );
  NAND2_X1 u0_u5_u4_U54 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n160 ) );
  NAND2_X1 u0_u5_u4_U55 (.ZN( u0_u5_u4_n134 ) , .A1( u0_u5_u4_n98 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U56 (.A1( u0_u5_u4_n103 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n143 ) );
  NAND2_X1 u0_u5_u4_U57 (.A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U58 (.A1( u0_u5_u4_n100 ) , .A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n120 ) );
  NAND2_X1 u0_u5_u4_U59 (.A1( u0_u5_u4_n102 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n148 ) );
  AOI21_X1 u0_u5_u4_U6 (.ZN( u0_u5_u4_n106 ) , .B2( u0_u5_u4_n146 ) , .B1( u0_u5_u4_n158 ) , .A( u0_u5_u4_n170 ) );
  NAND2_X1 u0_u5_u4_U60 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n157 ) );
  INV_X1 u0_u5_u4_U61 (.A( u0_u5_u4_n150 ) , .ZN( u0_u5_u4_n173 ) );
  INV_X1 u0_u5_u4_U62 (.A( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n171 ) );
  NAND2_X1 u0_u5_u4_U63 (.A1( u0_u5_u4_n100 ) , .ZN( u0_u5_u4_n118 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U64 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n144 ) );
  NAND2_X1 u0_u5_u4_U65 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U66 (.A( u0_u5_u4_n128 ) , .ZN( u0_u5_u4_n174 ) );
  NAND2_X1 u0_u5_u4_U67 (.A2( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n119 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U68 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U69 (.A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n113 ) , .A1( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U7 (.ZN( u0_u5_u4_n108 ) , .B2( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n155 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U70 (.A2( u0_u5_X_28 ) , .ZN( u0_u5_u4_n150 ) , .A1( u0_u5_u4_n168 ) );
  NOR2_X1 u0_u5_u4_U71 (.A2( u0_u5_X_29 ) , .ZN( u0_u5_u4_n152 ) , .A1( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U72 (.A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n105 ) , .A1( u0_u5_u4_n176 ) );
  NOR2_X1 u0_u5_u4_U73 (.A2( u0_u5_X_26 ) , .ZN( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n177 ) );
  NOR2_X1 u0_u5_u4_U74 (.A2( u0_u5_X_28 ) , .A1( u0_u5_X_29 ) , .ZN( u0_u5_u4_n128 ) );
  NOR2_X1 u0_u5_u4_U75 (.A2( u0_u5_X_27 ) , .A1( u0_u5_X_30 ) , .ZN( u0_u5_u4_n102 ) );
  NOR2_X1 u0_u5_u4_U76 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n98 ) );
  AND2_X1 u0_u5_u4_U77 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n104 ) );
  AND2_X1 u0_u5_u4_U78 (.A1( u0_u5_X_30 ) , .A2( u0_u5_u4_n176 ) , .ZN( u0_u5_u4_n99 ) );
  AND2_X1 u0_u5_u4_U79 (.A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n101 ) , .A2( u0_u5_u4_n177 ) );
  AOI21_X1 u0_u5_u4_U8 (.ZN( u0_u5_u4_n109 ) , .A( u0_u5_u4_n153 ) , .B1( u0_u5_u4_n159 ) , .B2( u0_u5_u4_n184 ) );
  AND2_X1 u0_u5_u4_U80 (.A1( u0_u5_X_27 ) , .A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n103 ) );
  INV_X1 u0_u5_u4_U81 (.A( u0_u5_X_28 ) , .ZN( u0_u5_u4_n169 ) );
  INV_X1 u0_u5_u4_U82 (.A( u0_u5_X_29 ) , .ZN( u0_u5_u4_n168 ) );
  INV_X1 u0_u5_u4_U83 (.A( u0_u5_X_25 ) , .ZN( u0_u5_u4_n177 ) );
  INV_X1 u0_u5_u4_U84 (.A( u0_u5_X_27 ) , .ZN( u0_u5_u4_n176 ) );
  NAND4_X1 u0_u5_u4_U85 (.ZN( u0_out5_25 ) , .A4( u0_u5_u4_n139 ) , .A3( u0_u5_u4_n140 ) , .A2( u0_u5_u4_n141 ) , .A1( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U86 (.A( u0_u5_u4_n128 ) , .B2( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n130 ) , .ZN( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U87 (.B2( u0_u5_u4_n131 ) , .ZN( u0_u5_u4_n141 ) , .A( u0_u5_u4_n175 ) , .B1( u0_u5_u4_n183 ) );
  NAND4_X1 u0_u5_u4_U88 (.ZN( u0_out5_14 ) , .A4( u0_u5_u4_n124 ) , .A3( u0_u5_u4_n125 ) , .A2( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n127 ) );
  AOI22_X1 u0_u5_u4_U89 (.B2( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n152 ) , .A2( u0_u5_u4_n175 ) );
  AOI211_X1 u0_u5_u4_U9 (.B( u0_u5_u4_n136 ) , .A( u0_u5_u4_n137 ) , .C2( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n139 ) , .C1( u0_u5_u4_n182 ) );
  AOI22_X1 u0_u5_u4_U90 (.ZN( u0_u5_u4_n125 ) , .B2( u0_u5_u4_n131 ) , .A2( u0_u5_u4_n132 ) , .B1( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n178 ) );
  NAND4_X1 u0_u5_u4_U91 (.ZN( u0_out5_8 ) , .A4( u0_u5_u4_n110 ) , .A3( u0_u5_u4_n111 ) , .A2( u0_u5_u4_n112 ) , .A1( u0_u5_u4_n186 ) );
  NAND2_X1 u0_u5_u4_U92 (.ZN( u0_u5_u4_n112 ) , .A2( u0_u5_u4_n130 ) , .A1( u0_u5_u4_n150 ) );
  AOI22_X1 u0_u5_u4_U93 (.ZN( u0_u5_u4_n111 ) , .B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n152 ) , .B1( u0_u5_u4_n178 ) , .A2( u0_u5_u4_n97 ) );
  AOI22_X1 u0_u5_u4_U94 (.B2( u0_u5_u4_n149 ) , .B1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n151 ) , .A1( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n167 ) );
  NOR4_X1 u0_u5_u4_U95 (.A4( u0_u5_u4_n162 ) , .A3( u0_u5_u4_n163 ) , .A2( u0_u5_u4_n164 ) , .A1( u0_u5_u4_n165 ) , .ZN( u0_u5_u4_n166 ) );
  NAND3_X1 u0_u5_u4_U96 (.ZN( u0_out5_3 ) , .A3( u0_u5_u4_n166 ) , .A1( u0_u5_u4_n167 ) , .A2( u0_u5_u4_n186 ) );
  NAND3_X1 u0_u5_u4_U97 (.A3( u0_u5_u4_n146 ) , .A2( u0_u5_u4_n147 ) , .A1( u0_u5_u4_n148 ) , .ZN( u0_u5_u4_n149 ) );
  NAND3_X1 u0_u5_u4_U98 (.A3( u0_u5_u4_n143 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n145 ) , .ZN( u0_u5_u4_n151 ) );
  NAND3_X1 u0_u5_u4_U99 (.A3( u0_u5_u4_n121 ) , .ZN( u0_u5_u4_n122 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n154 ) );
  INV_X1 u0_u5_u5_U10 (.A( u0_u5_u5_n121 ) , .ZN( u0_u5_u5_n177 ) );
  NOR3_X1 u0_u5_u5_U100 (.A3( u0_u5_u5_n141 ) , .A1( u0_u5_u5_n142 ) , .ZN( u0_u5_u5_n143 ) , .A2( u0_u5_u5_n191 ) );
  NAND4_X1 u0_u5_u5_U101 (.ZN( u0_out5_4 ) , .A4( u0_u5_u5_n112 ) , .A2( u0_u5_u5_n113 ) , .A1( u0_u5_u5_n114 ) , .A3( u0_u5_u5_n195 ) );
  AOI211_X1 u0_u5_u5_U102 (.A( u0_u5_u5_n110 ) , .C1( u0_u5_u5_n111 ) , .ZN( u0_u5_u5_n112 ) , .B( u0_u5_u5_n118 ) , .C2( u0_u5_u5_n177 ) );
  AOI222_X1 u0_u5_u5_U103 (.ZN( u0_u5_u5_n113 ) , .A1( u0_u5_u5_n131 ) , .C1( u0_u5_u5_n148 ) , .B2( u0_u5_u5_n174 ) , .C2( u0_u5_u5_n178 ) , .A2( u0_u5_u5_n179 ) , .B1( u0_u5_u5_n99 ) );
  NAND3_X1 u0_u5_u5_U104 (.A2( u0_u5_u5_n154 ) , .A3( u0_u5_u5_n158 ) , .A1( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n99 ) );
  NOR2_X1 u0_u5_u5_U11 (.ZN( u0_u5_u5_n160 ) , .A2( u0_u5_u5_n173 ) , .A1( u0_u5_u5_n177 ) );
  INV_X1 u0_u5_u5_U12 (.A( u0_u5_u5_n150 ) , .ZN( u0_u5_u5_n174 ) );
  AOI21_X1 u0_u5_u5_U13 (.A( u0_u5_u5_n160 ) , .B2( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n162 ) , .B1( u0_u5_u5_n192 ) );
  INV_X1 u0_u5_u5_U14 (.A( u0_u5_u5_n159 ) , .ZN( u0_u5_u5_n192 ) );
  AOI21_X1 u0_u5_u5_U15 (.A( u0_u5_u5_n156 ) , .B2( u0_u5_u5_n157 ) , .B1( u0_u5_u5_n158 ) , .ZN( u0_u5_u5_n163 ) );
  AOI21_X1 u0_u5_u5_U16 (.B2( u0_u5_u5_n139 ) , .B1( u0_u5_u5_n140 ) , .ZN( u0_u5_u5_n141 ) , .A( u0_u5_u5_n150 ) );
  OAI21_X1 u0_u5_u5_U17 (.A( u0_u5_u5_n133 ) , .B2( u0_u5_u5_n134 ) , .B1( u0_u5_u5_n135 ) , .ZN( u0_u5_u5_n142 ) );
  OAI21_X1 u0_u5_u5_U18 (.ZN( u0_u5_u5_n133 ) , .B2( u0_u5_u5_n147 ) , .A( u0_u5_u5_n173 ) , .B1( u0_u5_u5_n188 ) );
  NAND2_X1 u0_u5_u5_U19 (.A2( u0_u5_u5_n119 ) , .A1( u0_u5_u5_n123 ) , .ZN( u0_u5_u5_n137 ) );
  INV_X1 u0_u5_u5_U20 (.A( u0_u5_u5_n155 ) , .ZN( u0_u5_u5_n194 ) );
  NAND2_X1 u0_u5_u5_U21 (.A1( u0_u5_u5_n121 ) , .ZN( u0_u5_u5_n132 ) , .A2( u0_u5_u5_n172 ) );
  NAND2_X1 u0_u5_u5_U22 (.A2( u0_u5_u5_n122 ) , .ZN( u0_u5_u5_n136 ) , .A1( u0_u5_u5_n154 ) );
  NAND2_X1 u0_u5_u5_U23 (.A2( u0_u5_u5_n119 ) , .A1( u0_u5_u5_n120 ) , .ZN( u0_u5_u5_n159 ) );
  INV_X1 u0_u5_u5_U24 (.A( u0_u5_u5_n156 ) , .ZN( u0_u5_u5_n175 ) );
  INV_X1 u0_u5_u5_U25 (.A( u0_u5_u5_n158 ) , .ZN( u0_u5_u5_n188 ) );
  INV_X1 u0_u5_u5_U26 (.A( u0_u5_u5_n152 ) , .ZN( u0_u5_u5_n179 ) );
  INV_X1 u0_u5_u5_U27 (.A( u0_u5_u5_n140 ) , .ZN( u0_u5_u5_n182 ) );
  INV_X1 u0_u5_u5_U28 (.A( u0_u5_u5_n151 ) , .ZN( u0_u5_u5_n183 ) );
  INV_X1 u0_u5_u5_U29 (.A( u0_u5_u5_n123 ) , .ZN( u0_u5_u5_n185 ) );
  NOR2_X1 u0_u5_u5_U3 (.ZN( u0_u5_u5_n134 ) , .A1( u0_u5_u5_n183 ) , .A2( u0_u5_u5_n190 ) );
  INV_X1 u0_u5_u5_U30 (.A( u0_u5_u5_n161 ) , .ZN( u0_u5_u5_n184 ) );
  INV_X1 u0_u5_u5_U31 (.A( u0_u5_u5_n139 ) , .ZN( u0_u5_u5_n189 ) );
  INV_X1 u0_u5_u5_U32 (.A( u0_u5_u5_n157 ) , .ZN( u0_u5_u5_n190 ) );
  INV_X1 u0_u5_u5_U33 (.A( u0_u5_u5_n120 ) , .ZN( u0_u5_u5_n193 ) );
  NAND2_X1 u0_u5_u5_U34 (.ZN( u0_u5_u5_n111 ) , .A1( u0_u5_u5_n140 ) , .A2( u0_u5_u5_n155 ) );
  NOR2_X1 u0_u5_u5_U35 (.ZN( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n170 ) , .A2( u0_u5_u5_n180 ) );
  INV_X1 u0_u5_u5_U36 (.A( u0_u5_u5_n117 ) , .ZN( u0_u5_u5_n196 ) );
  OAI221_X1 u0_u5_u5_U37 (.A( u0_u5_u5_n116 ) , .ZN( u0_u5_u5_n117 ) , .B2( u0_u5_u5_n119 ) , .C1( u0_u5_u5_n153 ) , .C2( u0_u5_u5_n158 ) , .B1( u0_u5_u5_n172 ) );
  AOI222_X1 u0_u5_u5_U38 (.ZN( u0_u5_u5_n116 ) , .B2( u0_u5_u5_n145 ) , .C1( u0_u5_u5_n148 ) , .A2( u0_u5_u5_n174 ) , .C2( u0_u5_u5_n177 ) , .B1( u0_u5_u5_n187 ) , .A1( u0_u5_u5_n193 ) );
  INV_X1 u0_u5_u5_U39 (.A( u0_u5_u5_n115 ) , .ZN( u0_u5_u5_n187 ) );
  INV_X1 u0_u5_u5_U4 (.A( u0_u5_u5_n138 ) , .ZN( u0_u5_u5_n191 ) );
  AOI22_X1 u0_u5_u5_U40 (.B2( u0_u5_u5_n131 ) , .A2( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n169 ) , .B1( u0_u5_u5_n174 ) , .A1( u0_u5_u5_n185 ) );
  NOR2_X1 u0_u5_u5_U41 (.A1( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n150 ) , .A2( u0_u5_u5_n173 ) );
  AOI21_X1 u0_u5_u5_U42 (.A( u0_u5_u5_n118 ) , .B2( u0_u5_u5_n145 ) , .ZN( u0_u5_u5_n168 ) , .B1( u0_u5_u5_n186 ) );
  INV_X1 u0_u5_u5_U43 (.A( u0_u5_u5_n122 ) , .ZN( u0_u5_u5_n186 ) );
  NOR2_X1 u0_u5_u5_U44 (.A1( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n152 ) , .A2( u0_u5_u5_n176 ) );
  NOR2_X1 u0_u5_u5_U45 (.A1( u0_u5_u5_n115 ) , .ZN( u0_u5_u5_n118 ) , .A2( u0_u5_u5_n153 ) );
  NOR2_X1 u0_u5_u5_U46 (.A2( u0_u5_u5_n145 ) , .ZN( u0_u5_u5_n156 ) , .A1( u0_u5_u5_n174 ) );
  NOR2_X1 u0_u5_u5_U47 (.ZN( u0_u5_u5_n121 ) , .A2( u0_u5_u5_n145 ) , .A1( u0_u5_u5_n176 ) );
  AOI22_X1 u0_u5_u5_U48 (.ZN( u0_u5_u5_n114 ) , .A2( u0_u5_u5_n137 ) , .A1( u0_u5_u5_n145 ) , .B2( u0_u5_u5_n175 ) , .B1( u0_u5_u5_n193 ) );
  OAI211_X1 u0_u5_u5_U49 (.B( u0_u5_u5_n124 ) , .A( u0_u5_u5_n125 ) , .C2( u0_u5_u5_n126 ) , .C1( u0_u5_u5_n127 ) , .ZN( u0_u5_u5_n128 ) );
  OAI21_X1 u0_u5_u5_U5 (.B2( u0_u5_u5_n136 ) , .B1( u0_u5_u5_n137 ) , .ZN( u0_u5_u5_n138 ) , .A( u0_u5_u5_n177 ) );
  NOR3_X1 u0_u5_u5_U50 (.ZN( u0_u5_u5_n127 ) , .A1( u0_u5_u5_n136 ) , .A3( u0_u5_u5_n148 ) , .A2( u0_u5_u5_n182 ) );
  OAI21_X1 u0_u5_u5_U51 (.ZN( u0_u5_u5_n124 ) , .A( u0_u5_u5_n177 ) , .B2( u0_u5_u5_n183 ) , .B1( u0_u5_u5_n189 ) );
  OAI21_X1 u0_u5_u5_U52 (.ZN( u0_u5_u5_n125 ) , .A( u0_u5_u5_n174 ) , .B2( u0_u5_u5_n185 ) , .B1( u0_u5_u5_n190 ) );
  AOI21_X1 u0_u5_u5_U53 (.A( u0_u5_u5_n153 ) , .B2( u0_u5_u5_n154 ) , .B1( u0_u5_u5_n155 ) , .ZN( u0_u5_u5_n164 ) );
  AOI21_X1 u0_u5_u5_U54 (.ZN( u0_u5_u5_n110 ) , .B1( u0_u5_u5_n122 ) , .B2( u0_u5_u5_n139 ) , .A( u0_u5_u5_n153 ) );
  INV_X1 u0_u5_u5_U55 (.A( u0_u5_u5_n153 ) , .ZN( u0_u5_u5_n176 ) );
  INV_X1 u0_u5_u5_U56 (.A( u0_u5_u5_n126 ) , .ZN( u0_u5_u5_n173 ) );
  AND2_X1 u0_u5_u5_U57 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n147 ) );
  AND2_X1 u0_u5_u5_U58 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n148 ) );
  NAND2_X1 u0_u5_u5_U59 (.A1( u0_u5_u5_n105 ) , .A2( u0_u5_u5_n106 ) , .ZN( u0_u5_u5_n158 ) );
  INV_X1 u0_u5_u5_U6 (.A( u0_u5_u5_n135 ) , .ZN( u0_u5_u5_n178 ) );
  NAND2_X1 u0_u5_u5_U60 (.A2( u0_u5_u5_n108 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n139 ) );
  NAND2_X1 u0_u5_u5_U61 (.A1( u0_u5_u5_n106 ) , .A2( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n119 ) );
  NAND2_X1 u0_u5_u5_U62 (.A2( u0_u5_u5_n103 ) , .A1( u0_u5_u5_n105 ) , .ZN( u0_u5_u5_n140 ) );
  NAND2_X1 u0_u5_u5_U63 (.A2( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n105 ) , .ZN( u0_u5_u5_n155 ) );
  NAND2_X1 u0_u5_u5_U64 (.A2( u0_u5_u5_n106 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n122 ) );
  NAND2_X1 u0_u5_u5_U65 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n106 ) , .ZN( u0_u5_u5_n115 ) );
  NAND2_X1 u0_u5_u5_U66 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n103 ) , .ZN( u0_u5_u5_n161 ) );
  NAND2_X1 u0_u5_u5_U67 (.A1( u0_u5_u5_n105 ) , .A2( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n154 ) );
  INV_X1 u0_u5_u5_U68 (.A( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n172 ) );
  NAND2_X1 u0_u5_u5_U69 (.A1( u0_u5_u5_n103 ) , .A2( u0_u5_u5_n108 ) , .ZN( u0_u5_u5_n123 ) );
  OAI22_X1 u0_u5_u5_U7 (.B2( u0_u5_u5_n149 ) , .B1( u0_u5_u5_n150 ) , .A2( u0_u5_u5_n151 ) , .A1( u0_u5_u5_n152 ) , .ZN( u0_u5_u5_n165 ) );
  NAND2_X1 u0_u5_u5_U70 (.A2( u0_u5_u5_n103 ) , .A1( u0_u5_u5_n107 ) , .ZN( u0_u5_u5_n151 ) );
  NAND2_X1 u0_u5_u5_U71 (.A2( u0_u5_u5_n107 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n120 ) );
  NAND2_X1 u0_u5_u5_U72 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n109 ) , .ZN( u0_u5_u5_n157 ) );
  AND2_X1 u0_u5_u5_U73 (.A2( u0_u5_u5_n100 ) , .A1( u0_u5_u5_n104 ) , .ZN( u0_u5_u5_n131 ) );
  INV_X1 u0_u5_u5_U74 (.A( u0_u5_u5_n102 ) , .ZN( u0_u5_u5_n195 ) );
  OAI221_X1 u0_u5_u5_U75 (.A( u0_u5_u5_n101 ) , .ZN( u0_u5_u5_n102 ) , .C2( u0_u5_u5_n115 ) , .C1( u0_u5_u5_n126 ) , .B1( u0_u5_u5_n134 ) , .B2( u0_u5_u5_n160 ) );
  OAI21_X1 u0_u5_u5_U76 (.ZN( u0_u5_u5_n101 ) , .B1( u0_u5_u5_n137 ) , .A( u0_u5_u5_n146 ) , .B2( u0_u5_u5_n147 ) );
  NOR2_X1 u0_u5_u5_U77 (.A2( u0_u5_X_34 ) , .A1( u0_u5_X_35 ) , .ZN( u0_u5_u5_n145 ) );
  NOR2_X1 u0_u5_u5_U78 (.A2( u0_u5_X_34 ) , .ZN( u0_u5_u5_n146 ) , .A1( u0_u5_u5_n171 ) );
  NOR2_X1 u0_u5_u5_U79 (.A2( u0_u5_X_31 ) , .A1( u0_u5_X_32 ) , .ZN( u0_u5_u5_n103 ) );
  NOR3_X1 u0_u5_u5_U8 (.A2( u0_u5_u5_n147 ) , .A1( u0_u5_u5_n148 ) , .ZN( u0_u5_u5_n149 ) , .A3( u0_u5_u5_n194 ) );
  NOR2_X1 u0_u5_u5_U80 (.A2( u0_u5_X_36 ) , .ZN( u0_u5_u5_n105 ) , .A1( u0_u5_u5_n180 ) );
  NOR2_X1 u0_u5_u5_U81 (.A2( u0_u5_X_33 ) , .ZN( u0_u5_u5_n108 ) , .A1( u0_u5_u5_n170 ) );
  NOR2_X1 u0_u5_u5_U82 (.A2( u0_u5_X_33 ) , .A1( u0_u5_X_36 ) , .ZN( u0_u5_u5_n107 ) );
  NOR2_X1 u0_u5_u5_U83 (.A2( u0_u5_X_31 ) , .ZN( u0_u5_u5_n104 ) , .A1( u0_u5_u5_n181 ) );
  NAND2_X1 u0_u5_u5_U84 (.A2( u0_u5_X_34 ) , .A1( u0_u5_X_35 ) , .ZN( u0_u5_u5_n153 ) );
  NAND2_X1 u0_u5_u5_U85 (.A1( u0_u5_X_34 ) , .ZN( u0_u5_u5_n126 ) , .A2( u0_u5_u5_n171 ) );
  AND2_X1 u0_u5_u5_U86 (.A1( u0_u5_X_31 ) , .A2( u0_u5_X_32 ) , .ZN( u0_u5_u5_n106 ) );
  AND2_X1 u0_u5_u5_U87 (.A1( u0_u5_X_31 ) , .ZN( u0_u5_u5_n109 ) , .A2( u0_u5_u5_n181 ) );
  INV_X1 u0_u5_u5_U88 (.A( u0_u5_X_33 ) , .ZN( u0_u5_u5_n180 ) );
  INV_X1 u0_u5_u5_U89 (.A( u0_u5_X_35 ) , .ZN( u0_u5_u5_n171 ) );
  NOR2_X1 u0_u5_u5_U9 (.ZN( u0_u5_u5_n135 ) , .A1( u0_u5_u5_n173 ) , .A2( u0_u5_u5_n176 ) );
  INV_X1 u0_u5_u5_U90 (.A( u0_u5_X_36 ) , .ZN( u0_u5_u5_n170 ) );
  INV_X1 u0_u5_u5_U91 (.A( u0_u5_X_32 ) , .ZN( u0_u5_u5_n181 ) );
  NAND4_X1 u0_u5_u5_U92 (.ZN( u0_out5_29 ) , .A4( u0_u5_u5_n129 ) , .A3( u0_u5_u5_n130 ) , .A2( u0_u5_u5_n168 ) , .A1( u0_u5_u5_n196 ) );
  AOI221_X1 u0_u5_u5_U93 (.A( u0_u5_u5_n128 ) , .ZN( u0_u5_u5_n129 ) , .C2( u0_u5_u5_n132 ) , .B2( u0_u5_u5_n159 ) , .B1( u0_u5_u5_n176 ) , .C1( u0_u5_u5_n184 ) );
  AOI222_X1 u0_u5_u5_U94 (.ZN( u0_u5_u5_n130 ) , .A2( u0_u5_u5_n146 ) , .B1( u0_u5_u5_n147 ) , .C2( u0_u5_u5_n175 ) , .B2( u0_u5_u5_n179 ) , .A1( u0_u5_u5_n188 ) , .C1( u0_u5_u5_n194 ) );
  NAND4_X1 u0_u5_u5_U95 (.ZN( u0_out5_19 ) , .A4( u0_u5_u5_n166 ) , .A3( u0_u5_u5_n167 ) , .A2( u0_u5_u5_n168 ) , .A1( u0_u5_u5_n169 ) );
  AOI22_X1 u0_u5_u5_U96 (.B2( u0_u5_u5_n145 ) , .A2( u0_u5_u5_n146 ) , .ZN( u0_u5_u5_n167 ) , .B1( u0_u5_u5_n182 ) , .A1( u0_u5_u5_n189 ) );
  NOR4_X1 u0_u5_u5_U97 (.A4( u0_u5_u5_n162 ) , .A3( u0_u5_u5_n163 ) , .A2( u0_u5_u5_n164 ) , .A1( u0_u5_u5_n165 ) , .ZN( u0_u5_u5_n166 ) );
  NAND4_X1 u0_u5_u5_U98 (.ZN( u0_out5_11 ) , .A4( u0_u5_u5_n143 ) , .A3( u0_u5_u5_n144 ) , .A2( u0_u5_u5_n169 ) , .A1( u0_u5_u5_n196 ) );
  AOI22_X1 u0_u5_u5_U99 (.A2( u0_u5_u5_n132 ) , .ZN( u0_u5_u5_n144 ) , .B2( u0_u5_u5_n145 ) , .B1( u0_u5_u5_n184 ) , .A1( u0_u5_u5_n194 ) );
  OAI21_X1 u0_u5_u6_U10 (.A( u0_u5_u6_n159 ) , .B1( u0_u5_u6_n169 ) , .B2( u0_u5_u6_n173 ) , .ZN( u0_u5_u6_n90 ) );
  INV_X1 u0_u5_u6_U11 (.ZN( u0_u5_u6_n172 ) , .A( u0_u5_u6_n88 ) );
  AOI22_X1 u0_u5_u6_U12 (.A2( u0_u5_u6_n151 ) , .B2( u0_u5_u6_n161 ) , .A1( u0_u5_u6_n167 ) , .B1( u0_u5_u6_n170 ) , .ZN( u0_u5_u6_n89 ) );
  AOI21_X1 u0_u5_u6_U13 (.ZN( u0_u5_u6_n106 ) , .A( u0_u5_u6_n142 ) , .B2( u0_u5_u6_n159 ) , .B1( u0_u5_u6_n164 ) );
  INV_X1 u0_u5_u6_U14 (.A( u0_u5_u6_n155 ) , .ZN( u0_u5_u6_n161 ) );
  INV_X1 u0_u5_u6_U15 (.A( u0_u5_u6_n128 ) , .ZN( u0_u5_u6_n164 ) );
  NAND2_X1 u0_u5_u6_U16 (.ZN( u0_u5_u6_n110 ) , .A1( u0_u5_u6_n122 ) , .A2( u0_u5_u6_n129 ) );
  NAND2_X1 u0_u5_u6_U17 (.ZN( u0_u5_u6_n124 ) , .A2( u0_u5_u6_n146 ) , .A1( u0_u5_u6_n148 ) );
  INV_X1 u0_u5_u6_U18 (.A( u0_u5_u6_n132 ) , .ZN( u0_u5_u6_n171 ) );
  AND2_X1 u0_u5_u6_U19 (.A1( u0_u5_u6_n100 ) , .ZN( u0_u5_u6_n130 ) , .A2( u0_u5_u6_n147 ) );
  INV_X1 u0_u5_u6_U20 (.A( u0_u5_u6_n127 ) , .ZN( u0_u5_u6_n173 ) );
  INV_X1 u0_u5_u6_U21 (.A( u0_u5_u6_n121 ) , .ZN( u0_u5_u6_n167 ) );
  INV_X1 u0_u5_u6_U22 (.A( u0_u5_u6_n100 ) , .ZN( u0_u5_u6_n169 ) );
  INV_X1 u0_u5_u6_U23 (.A( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n170 ) );
  INV_X1 u0_u5_u6_U24 (.A( u0_u5_u6_n113 ) , .ZN( u0_u5_u6_n168 ) );
  AND2_X1 u0_u5_u6_U25 (.A1( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n119 ) , .ZN( u0_u5_u6_n133 ) );
  AND2_X1 u0_u5_u6_U26 (.A2( u0_u5_u6_n121 ) , .A1( u0_u5_u6_n122 ) , .ZN( u0_u5_u6_n131 ) );
  AND3_X1 u0_u5_u6_U27 (.ZN( u0_u5_u6_n120 ) , .A2( u0_u5_u6_n127 ) , .A1( u0_u5_u6_n132 ) , .A3( u0_u5_u6_n145 ) );
  INV_X1 u0_u5_u6_U28 (.A( u0_u5_u6_n146 ) , .ZN( u0_u5_u6_n163 ) );
  AOI222_X1 u0_u5_u6_U29 (.ZN( u0_u5_u6_n114 ) , .A1( u0_u5_u6_n118 ) , .A2( u0_u5_u6_n126 ) , .B2( u0_u5_u6_n151 ) , .C2( u0_u5_u6_n159 ) , .C1( u0_u5_u6_n168 ) , .B1( u0_u5_u6_n169 ) );
  INV_X1 u0_u5_u6_U3 (.A( u0_u5_u6_n110 ) , .ZN( u0_u5_u6_n166 ) );
  NOR2_X1 u0_u5_u6_U30 (.A1( u0_u5_u6_n162 ) , .A2( u0_u5_u6_n165 ) , .ZN( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U31 (.A1( u0_u5_u6_n144 ) , .ZN( u0_u5_u6_n151 ) , .A2( u0_u5_u6_n158 ) );
  NAND2_X1 u0_u5_u6_U32 (.ZN( u0_u5_u6_n132 ) , .A1( u0_u5_u6_n91 ) , .A2( u0_u5_u6_n97 ) );
  NOR2_X1 u0_u5_u6_U33 (.A2( u0_u5_u6_n126 ) , .ZN( u0_u5_u6_n155 ) , .A1( u0_u5_u6_n160 ) );
  NAND2_X1 u0_u5_u6_U34 (.ZN( u0_u5_u6_n146 ) , .A2( u0_u5_u6_n94 ) , .A1( u0_u5_u6_n99 ) );
  AOI21_X1 u0_u5_u6_U35 (.A( u0_u5_u6_n144 ) , .B2( u0_u5_u6_n145 ) , .B1( u0_u5_u6_n146 ) , .ZN( u0_u5_u6_n150 ) );
  INV_X1 u0_u5_u6_U36 (.A( u0_u5_u6_n111 ) , .ZN( u0_u5_u6_n158 ) );
  NAND2_X1 u0_u5_u6_U37 (.ZN( u0_u5_u6_n127 ) , .A1( u0_u5_u6_n91 ) , .A2( u0_u5_u6_n92 ) );
  NAND2_X1 u0_u5_u6_U38 (.ZN( u0_u5_u6_n129 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n96 ) );
  INV_X1 u0_u5_u6_U39 (.A( u0_u5_u6_n144 ) , .ZN( u0_u5_u6_n159 ) );
  INV_X1 u0_u5_u6_U4 (.A( u0_u5_u6_n142 ) , .ZN( u0_u5_u6_n174 ) );
  NAND2_X1 u0_u5_u6_U40 (.ZN( u0_u5_u6_n145 ) , .A2( u0_u5_u6_n97 ) , .A1( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U41 (.ZN( u0_u5_u6_n148 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n94 ) );
  NAND2_X1 u0_u5_u6_U42 (.ZN( u0_u5_u6_n108 ) , .A2( u0_u5_u6_n139 ) , .A1( u0_u5_u6_n144 ) );
  NAND2_X1 u0_u5_u6_U43 (.ZN( u0_u5_u6_n121 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n97 ) );
  NAND2_X1 u0_u5_u6_U44 (.ZN( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n95 ) );
  AND2_X1 u0_u5_u6_U45 (.ZN( u0_u5_u6_n118 ) , .A2( u0_u5_u6_n91 ) , .A1( u0_u5_u6_n99 ) );
  AOI22_X1 u0_u5_u6_U46 (.B2( u0_u5_u6_n110 ) , .B1( u0_u5_u6_n111 ) , .A1( u0_u5_u6_n112 ) , .ZN( u0_u5_u6_n115 ) , .A2( u0_u5_u6_n161 ) );
  NAND4_X1 u0_u5_u6_U47 (.A3( u0_u5_u6_n109 ) , .ZN( u0_u5_u6_n112 ) , .A4( u0_u5_u6_n132 ) , .A2( u0_u5_u6_n147 ) , .A1( u0_u5_u6_n166 ) );
  NOR2_X1 u0_u5_u6_U48 (.ZN( u0_u5_u6_n109 ) , .A1( u0_u5_u6_n170 ) , .A2( u0_u5_u6_n173 ) );
  NAND2_X1 u0_u5_u6_U49 (.ZN( u0_u5_u6_n147 ) , .A2( u0_u5_u6_n98 ) , .A1( u0_u5_u6_n99 ) );
  NAND2_X1 u0_u5_u6_U5 (.A2( u0_u5_u6_n143 ) , .ZN( u0_u5_u6_n152 ) , .A1( u0_u5_u6_n166 ) );
  NAND2_X1 u0_u5_u6_U50 (.ZN( u0_u5_u6_n128 ) , .A1( u0_u5_u6_n94 ) , .A2( u0_u5_u6_n96 ) );
  AOI211_X1 u0_u5_u6_U51 (.B( u0_u5_u6_n134 ) , .A( u0_u5_u6_n135 ) , .C1( u0_u5_u6_n136 ) , .ZN( u0_u5_u6_n137 ) , .C2( u0_u5_u6_n151 ) );
  AOI21_X1 u0_u5_u6_U52 (.B2( u0_u5_u6_n132 ) , .B1( u0_u5_u6_n133 ) , .ZN( u0_u5_u6_n134 ) , .A( u0_u5_u6_n158 ) );
  AOI21_X1 u0_u5_u6_U53 (.B1( u0_u5_u6_n131 ) , .ZN( u0_u5_u6_n135 ) , .A( u0_u5_u6_n144 ) , .B2( u0_u5_u6_n146 ) );
  NAND4_X1 u0_u5_u6_U54 (.A4( u0_u5_u6_n127 ) , .A3( u0_u5_u6_n128 ) , .A2( u0_u5_u6_n129 ) , .A1( u0_u5_u6_n130 ) , .ZN( u0_u5_u6_n136 ) );
  NAND2_X1 u0_u5_u6_U55 (.ZN( u0_u5_u6_n119 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n99 ) );
  NAND2_X1 u0_u5_u6_U56 (.ZN( u0_u5_u6_n123 ) , .A2( u0_u5_u6_n91 ) , .A1( u0_u5_u6_n96 ) );
  NAND2_X1 u0_u5_u6_U57 (.ZN( u0_u5_u6_n100 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U58 (.ZN( u0_u5_u6_n122 ) , .A1( u0_u5_u6_n94 ) , .A2( u0_u5_u6_n97 ) );
  INV_X1 u0_u5_u6_U59 (.A( u0_u5_u6_n139 ) , .ZN( u0_u5_u6_n160 ) );
  AOI22_X1 u0_u5_u6_U6 (.B2( u0_u5_u6_n101 ) , .A1( u0_u5_u6_n102 ) , .ZN( u0_u5_u6_n103 ) , .B1( u0_u5_u6_n160 ) , .A2( u0_u5_u6_n161 ) );
  NAND2_X1 u0_u5_u6_U60 (.ZN( u0_u5_u6_n113 ) , .A1( u0_u5_u6_n96 ) , .A2( u0_u5_u6_n98 ) );
  NOR2_X1 u0_u5_u6_U61 (.A2( u0_u5_X_40 ) , .A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n126 ) );
  NOR2_X1 u0_u5_u6_U62 (.A2( u0_u5_X_39 ) , .A1( u0_u5_X_42 ) , .ZN( u0_u5_u6_n92 ) );
  NOR2_X1 u0_u5_u6_U63 (.A2( u0_u5_X_39 ) , .A1( u0_u5_u6_n156 ) , .ZN( u0_u5_u6_n97 ) );
  NOR2_X1 u0_u5_u6_U64 (.A2( u0_u5_X_38 ) , .A1( u0_u5_u6_n165 ) , .ZN( u0_u5_u6_n95 ) );
  NOR2_X1 u0_u5_u6_U65 (.A2( u0_u5_X_41 ) , .ZN( u0_u5_u6_n111 ) , .A1( u0_u5_u6_n157 ) );
  NOR2_X1 u0_u5_u6_U66 (.A2( u0_u5_X_37 ) , .A1( u0_u5_u6_n162 ) , .ZN( u0_u5_u6_n94 ) );
  NOR2_X1 u0_u5_u6_U67 (.A2( u0_u5_X_37 ) , .A1( u0_u5_X_38 ) , .ZN( u0_u5_u6_n91 ) );
  NAND2_X1 u0_u5_u6_U68 (.A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n144 ) , .A2( u0_u5_u6_n157 ) );
  NAND2_X1 u0_u5_u6_U69 (.A2( u0_u5_X_40 ) , .A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n139 ) );
  NOR2_X1 u0_u5_u6_U7 (.A1( u0_u5_u6_n118 ) , .ZN( u0_u5_u6_n143 ) , .A2( u0_u5_u6_n168 ) );
  AND2_X1 u0_u5_u6_U70 (.A1( u0_u5_X_39 ) , .A2( u0_u5_u6_n156 ) , .ZN( u0_u5_u6_n96 ) );
  AND2_X1 u0_u5_u6_U71 (.A1( u0_u5_X_39 ) , .A2( u0_u5_X_42 ) , .ZN( u0_u5_u6_n99 ) );
  INV_X1 u0_u5_u6_U72 (.A( u0_u5_X_40 ) , .ZN( u0_u5_u6_n157 ) );
  INV_X1 u0_u5_u6_U73 (.A( u0_u5_X_37 ) , .ZN( u0_u5_u6_n165 ) );
  INV_X1 u0_u5_u6_U74 (.A( u0_u5_X_38 ) , .ZN( u0_u5_u6_n162 ) );
  INV_X1 u0_u5_u6_U75 (.A( u0_u5_X_42 ) , .ZN( u0_u5_u6_n156 ) );
  NAND4_X1 u0_u5_u6_U76 (.ZN( u0_out5_32 ) , .A4( u0_u5_u6_n103 ) , .A3( u0_u5_u6_n104 ) , .A2( u0_u5_u6_n105 ) , .A1( u0_u5_u6_n106 ) );
  AOI22_X1 u0_u5_u6_U77 (.ZN( u0_u5_u6_n105 ) , .A2( u0_u5_u6_n108 ) , .A1( u0_u5_u6_n118 ) , .B2( u0_u5_u6_n126 ) , .B1( u0_u5_u6_n171 ) );
  AOI22_X1 u0_u5_u6_U78 (.ZN( u0_u5_u6_n104 ) , .A1( u0_u5_u6_n111 ) , .B1( u0_u5_u6_n124 ) , .B2( u0_u5_u6_n151 ) , .A2( u0_u5_u6_n93 ) );
  NAND4_X1 u0_u5_u6_U79 (.ZN( u0_out5_12 ) , .A4( u0_u5_u6_n114 ) , .A3( u0_u5_u6_n115 ) , .A2( u0_u5_u6_n116 ) , .A1( u0_u5_u6_n117 ) );
  AOI21_X1 u0_u5_u6_U8 (.B1( u0_u5_u6_n107 ) , .B2( u0_u5_u6_n132 ) , .A( u0_u5_u6_n158 ) , .ZN( u0_u5_u6_n88 ) );
  OAI22_X1 u0_u5_u6_U80 (.B2( u0_u5_u6_n111 ) , .ZN( u0_u5_u6_n116 ) , .B1( u0_u5_u6_n126 ) , .A2( u0_u5_u6_n164 ) , .A1( u0_u5_u6_n167 ) );
  OAI21_X1 u0_u5_u6_U81 (.A( u0_u5_u6_n108 ) , .ZN( u0_u5_u6_n117 ) , .B2( u0_u5_u6_n141 ) , .B1( u0_u5_u6_n163 ) );
  OAI211_X1 u0_u5_u6_U82 (.ZN( u0_out5_22 ) , .B( u0_u5_u6_n137 ) , .A( u0_u5_u6_n138 ) , .C2( u0_u5_u6_n139 ) , .C1( u0_u5_u6_n140 ) );
  AOI22_X1 u0_u5_u6_U83 (.B1( u0_u5_u6_n124 ) , .A2( u0_u5_u6_n125 ) , .A1( u0_u5_u6_n126 ) , .ZN( u0_u5_u6_n138 ) , .B2( u0_u5_u6_n161 ) );
  AND4_X1 u0_u5_u6_U84 (.A3( u0_u5_u6_n119 ) , .A1( u0_u5_u6_n120 ) , .A4( u0_u5_u6_n129 ) , .ZN( u0_u5_u6_n140 ) , .A2( u0_u5_u6_n143 ) );
  OAI211_X1 u0_u5_u6_U85 (.ZN( u0_out5_7 ) , .B( u0_u5_u6_n153 ) , .C2( u0_u5_u6_n154 ) , .C1( u0_u5_u6_n155 ) , .A( u0_u5_u6_n174 ) );
  NOR3_X1 u0_u5_u6_U86 (.A1( u0_u5_u6_n141 ) , .ZN( u0_u5_u6_n154 ) , .A3( u0_u5_u6_n164 ) , .A2( u0_u5_u6_n171 ) );
  AOI211_X1 u0_u5_u6_U87 (.B( u0_u5_u6_n149 ) , .A( u0_u5_u6_n150 ) , .C2( u0_u5_u6_n151 ) , .C1( u0_u5_u6_n152 ) , .ZN( u0_u5_u6_n153 ) );
  NAND3_X1 u0_u5_u6_U88 (.A2( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n125 ) , .A1( u0_u5_u6_n130 ) , .A3( u0_u5_u6_n131 ) );
  NAND3_X1 u0_u5_u6_U89 (.A3( u0_u5_u6_n133 ) , .ZN( u0_u5_u6_n141 ) , .A1( u0_u5_u6_n145 ) , .A2( u0_u5_u6_n148 ) );
  AOI21_X1 u0_u5_u6_U9 (.B2( u0_u5_u6_n147 ) , .B1( u0_u5_u6_n148 ) , .ZN( u0_u5_u6_n149 ) , .A( u0_u5_u6_n158 ) );
  NAND3_X1 u0_u5_u6_U90 (.ZN( u0_u5_u6_n101 ) , .A3( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n121 ) , .A1( u0_u5_u6_n127 ) );
  NAND3_X1 u0_u5_u6_U91 (.ZN( u0_u5_u6_n102 ) , .A3( u0_u5_u6_n130 ) , .A2( u0_u5_u6_n145 ) , .A1( u0_u5_u6_n166 ) );
  NAND3_X1 u0_u5_u6_U92 (.A3( u0_u5_u6_n113 ) , .A1( u0_u5_u6_n119 ) , .A2( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n93 ) );
  NAND3_X1 u0_u5_u6_U93 (.ZN( u0_u5_u6_n142 ) , .A2( u0_u5_u6_n172 ) , .A3( u0_u5_u6_n89 ) , .A1( u0_u5_u6_n90 ) );
  XOR2_X1 u0_u6_U1 (.B( u0_K7_9 ) , .A( u0_R5_6 ) , .Z( u0_u6_X_9 ) );
  XOR2_X1 u0_u6_U10 (.B( u0_K7_45 ) , .A( u0_R5_30 ) , .Z( u0_u6_X_45 ) );
  XOR2_X1 u0_u6_U11 (.B( u0_K7_44 ) , .A( u0_R5_29 ) , .Z( u0_u6_X_44 ) );
  XOR2_X1 u0_u6_U12 (.B( u0_K7_43 ) , .A( u0_R5_28 ) , .Z( u0_u6_X_43 ) );
  XOR2_X1 u0_u6_U16 (.B( u0_K7_3 ) , .A( u0_R5_2 ) , .Z( u0_u6_X_3 ) );
  XOR2_X1 u0_u6_U2 (.B( u0_K7_8 ) , .A( u0_R5_5 ) , .Z( u0_u6_X_8 ) );
  XOR2_X1 u0_u6_U27 (.B( u0_K7_2 ) , .A( u0_R5_1 ) , .Z( u0_u6_X_2 ) );
  XOR2_X1 u0_u6_U3 (.B( u0_K7_7 ) , .A( u0_R5_4 ) , .Z( u0_u6_X_7 ) );
  XOR2_X1 u0_u6_U33 (.B( u0_K7_24 ) , .A( u0_R5_17 ) , .Z( u0_u6_X_24 ) );
  XOR2_X1 u0_u6_U34 (.B( u0_K7_23 ) , .A( u0_R5_16 ) , .Z( u0_u6_X_23 ) );
  XOR2_X1 u0_u6_U35 (.B( u0_K7_22 ) , .A( u0_R5_15 ) , .Z( u0_u6_X_22 ) );
  XOR2_X1 u0_u6_U36 (.B( u0_K7_21 ) , .A( u0_R5_14 ) , .Z( u0_u6_X_21 ) );
  XOR2_X1 u0_u6_U37 (.B( u0_K7_20 ) , .A( u0_R5_13 ) , .Z( u0_u6_X_20 ) );
  XOR2_X1 u0_u6_U38 (.B( u0_K7_1 ) , .A( u0_R5_32 ) , .Z( u0_u6_X_1 ) );
  XOR2_X1 u0_u6_U39 (.B( u0_K7_19 ) , .A( u0_R5_12 ) , .Z( u0_u6_X_19 ) );
  XOR2_X1 u0_u6_U4 (.B( u0_K7_6 ) , .A( u0_R5_5 ) , .Z( u0_u6_X_6 ) );
  XOR2_X1 u0_u6_U40 (.B( u0_K7_18 ) , .A( u0_R5_13 ) , .Z( u0_u6_X_18 ) );
  XOR2_X1 u0_u6_U41 (.B( u0_K7_17 ) , .A( u0_R5_12 ) , .Z( u0_u6_X_17 ) );
  XOR2_X1 u0_u6_U42 (.B( u0_K7_16 ) , .A( u0_R5_11 ) , .Z( u0_u6_X_16 ) );
  XOR2_X1 u0_u6_U43 (.B( u0_K7_15 ) , .A( u0_R5_10 ) , .Z( u0_u6_X_15 ) );
  XOR2_X1 u0_u6_U44 (.B( u0_K7_14 ) , .A( u0_R5_9 ) , .Z( u0_u6_X_14 ) );
  XOR2_X1 u0_u6_U45 (.B( u0_K7_13 ) , .A( u0_R5_8 ) , .Z( u0_u6_X_13 ) );
  XOR2_X1 u0_u6_U46 (.B( u0_K7_12 ) , .A( u0_R5_9 ) , .Z( u0_u6_X_12 ) );
  XOR2_X1 u0_u6_U47 (.B( u0_K7_11 ) , .A( u0_R5_8 ) , .Z( u0_u6_X_11 ) );
  XOR2_X1 u0_u6_U48 (.B( u0_K7_10 ) , .A( u0_R5_7 ) , .Z( u0_u6_X_10 ) );
  XOR2_X1 u0_u6_U5 (.B( u0_K7_5 ) , .A( u0_R5_4 ) , .Z( u0_u6_X_5 ) );
  XOR2_X1 u0_u6_U6 (.B( u0_K7_4 ) , .A( u0_R5_3 ) , .Z( u0_u6_X_4 ) );
  XOR2_X1 u0_u6_U7 (.B( u0_K7_48 ) , .A( u0_R5_1 ) , .Z( u0_u6_X_48 ) );
  XOR2_X1 u0_u6_U8 (.B( u0_K7_47 ) , .A( u0_R5_32 ) , .Z( u0_u6_X_47 ) );
  XOR2_X1 u0_u6_U9 (.B( u0_K7_46 ) , .A( u0_R5_31 ) , .Z( u0_u6_X_46 ) );
  NAND2_X1 u0_u6_u0_U10 (.ZN( u0_u6_u0_n113 ) , .A1( u0_u6_u0_n139 ) , .A2( u0_u6_u0_n149 ) );
  AND2_X1 u0_u6_u0_U11 (.A1( u0_u6_u0_n131 ) , .ZN( u0_u6_u0_n141 ) , .A2( u0_u6_u0_n150 ) );
  AND2_X1 u0_u6_u0_U12 (.ZN( u0_u6_u0_n107 ) , .A1( u0_u6_u0_n130 ) , .A2( u0_u6_u0_n140 ) );
  AND2_X1 u0_u6_u0_U13 (.A2( u0_u6_u0_n129 ) , .A1( u0_u6_u0_n130 ) , .ZN( u0_u6_u0_n151 ) );
  AND2_X1 u0_u6_u0_U14 (.A1( u0_u6_u0_n108 ) , .A2( u0_u6_u0_n125 ) , .ZN( u0_u6_u0_n145 ) );
  INV_X1 u0_u6_u0_U15 (.A( u0_u6_u0_n143 ) , .ZN( u0_u6_u0_n173 ) );
  NOR2_X1 u0_u6_u0_U16 (.A2( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n147 ) , .A1( u0_u6_u0_n160 ) );
  AOI21_X1 u0_u6_u0_U17 (.B1( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n132 ) , .A( u0_u6_u0_n165 ) , .B2( u0_u6_u0_n93 ) );
  OAI221_X1 u0_u6_u0_U18 (.C1( u0_u6_u0_n121 ) , .ZN( u0_u6_u0_n122 ) , .B2( u0_u6_u0_n127 ) , .A( u0_u6_u0_n143 ) , .B1( u0_u6_u0_n144 ) , .C2( u0_u6_u0_n147 ) );
  OAI22_X1 u0_u6_u0_U19 (.B1( u0_u6_u0_n125 ) , .ZN( u0_u6_u0_n126 ) , .A1( u0_u6_u0_n138 ) , .A2( u0_u6_u0_n146 ) , .B2( u0_u6_u0_n147 ) );
  OAI22_X1 u0_u6_u0_U20 (.B1( u0_u6_u0_n131 ) , .A1( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n147 ) , .A2( u0_u6_u0_n90 ) , .ZN( u0_u6_u0_n91 ) );
  AND3_X1 u0_u6_u0_U21 (.A3( u0_u6_u0_n121 ) , .A2( u0_u6_u0_n125 ) , .A1( u0_u6_u0_n148 ) , .ZN( u0_u6_u0_n90 ) );
  NOR2_X1 u0_u6_u0_U22 (.A1( u0_u6_u0_n163 ) , .A2( u0_u6_u0_n164 ) , .ZN( u0_u6_u0_n95 ) );
  NOR2_X1 u0_u6_u0_U23 (.A1( u0_u6_u0_n120 ) , .ZN( u0_u6_u0_n143 ) , .A2( u0_u6_u0_n167 ) );
  OAI221_X1 u0_u6_u0_U24 (.C1( u0_u6_u0_n112 ) , .ZN( u0_u6_u0_n120 ) , .B1( u0_u6_u0_n138 ) , .B2( u0_u6_u0_n141 ) , .C2( u0_u6_u0_n147 ) , .A( u0_u6_u0_n172 ) );
  AOI211_X1 u0_u6_u0_U25 (.B( u0_u6_u0_n115 ) , .A( u0_u6_u0_n116 ) , .C2( u0_u6_u0_n117 ) , .C1( u0_u6_u0_n118 ) , .ZN( u0_u6_u0_n119 ) );
  AOI22_X1 u0_u6_u0_U26 (.B2( u0_u6_u0_n109 ) , .A2( u0_u6_u0_n110 ) , .ZN( u0_u6_u0_n111 ) , .B1( u0_u6_u0_n118 ) , .A1( u0_u6_u0_n160 ) );
  NAND2_X1 u0_u6_u0_U27 (.A1( u0_u6_u0_n100 ) , .A2( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n125 ) );
  INV_X1 u0_u6_u0_U28 (.A( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U29 (.A( u0_u6_u0_n118 ) , .ZN( u0_u6_u0_n158 ) );
  INV_X1 u0_u6_u0_U3 (.A( u0_u6_u0_n113 ) , .ZN( u0_u6_u0_n166 ) );
  AOI21_X1 u0_u6_u0_U30 (.B1( u0_u6_u0_n127 ) , .B2( u0_u6_u0_n129 ) , .A( u0_u6_u0_n138 ) , .ZN( u0_u6_u0_n96 ) );
  AOI21_X1 u0_u6_u0_U31 (.ZN( u0_u6_u0_n104 ) , .B1( u0_u6_u0_n107 ) , .B2( u0_u6_u0_n141 ) , .A( u0_u6_u0_n144 ) );
  NAND2_X1 u0_u6_u0_U32 (.A2( u0_u6_u0_n102 ) , .A1( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n149 ) );
  NAND2_X1 u0_u6_u0_U33 (.A2( u0_u6_u0_n100 ) , .ZN( u0_u6_u0_n131 ) , .A1( u0_u6_u0_n92 ) );
  NAND2_X1 u0_u6_u0_U34 (.A2( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n114 ) , .A1( u0_u6_u0_n92 ) );
  NAND2_X1 u0_u6_u0_U35 (.A1( u0_u6_u0_n101 ) , .A2( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n150 ) );
  INV_X1 u0_u6_u0_U36 (.A( u0_u6_u0_n138 ) , .ZN( u0_u6_u0_n160 ) );
  NAND2_X1 u0_u6_u0_U37 (.A2( u0_u6_u0_n100 ) , .A1( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n139 ) );
  NAND2_X1 u0_u6_u0_U38 (.ZN( u0_u6_u0_n112 ) , .A2( u0_u6_u0_n92 ) , .A1( u0_u6_u0_n93 ) );
  NAND2_X1 u0_u6_u0_U39 (.A2( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n121 ) , .A1( u0_u6_u0_n93 ) );
  AOI21_X1 u0_u6_u0_U4 (.B1( u0_u6_u0_n114 ) , .ZN( u0_u6_u0_n115 ) , .B2( u0_u6_u0_n129 ) , .A( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U40 (.ZN( u0_u6_u0_n172 ) , .A( u0_u6_u0_n88 ) );
  OAI222_X1 u0_u6_u0_U41 (.C1( u0_u6_u0_n108 ) , .A1( u0_u6_u0_n125 ) , .B2( u0_u6_u0_n128 ) , .B1( u0_u6_u0_n144 ) , .A2( u0_u6_u0_n158 ) , .C2( u0_u6_u0_n161 ) , .ZN( u0_u6_u0_n88 ) );
  OR3_X1 u0_u6_u0_U42 (.A3( u0_u6_u0_n152 ) , .A2( u0_u6_u0_n153 ) , .A1( u0_u6_u0_n154 ) , .ZN( u0_u6_u0_n155 ) );
  AOI21_X1 u0_u6_u0_U43 (.A( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n145 ) , .B1( u0_u6_u0_n146 ) , .ZN( u0_u6_u0_n154 ) );
  AOI21_X1 u0_u6_u0_U44 (.B2( u0_u6_u0_n150 ) , .B1( u0_u6_u0_n151 ) , .ZN( u0_u6_u0_n152 ) , .A( u0_u6_u0_n158 ) );
  AOI21_X1 u0_u6_u0_U45 (.A( u0_u6_u0_n147 ) , .B2( u0_u6_u0_n148 ) , .B1( u0_u6_u0_n149 ) , .ZN( u0_u6_u0_n153 ) );
  INV_X1 u0_u6_u0_U46 (.ZN( u0_u6_u0_n171 ) , .A( u0_u6_u0_n99 ) );
  OAI211_X1 u0_u6_u0_U47 (.C2( u0_u6_u0_n140 ) , .C1( u0_u6_u0_n161 ) , .A( u0_u6_u0_n169 ) , .B( u0_u6_u0_n98 ) , .ZN( u0_u6_u0_n99 ) );
  AOI211_X1 u0_u6_u0_U48 (.C1( u0_u6_u0_n118 ) , .A( u0_u6_u0_n123 ) , .B( u0_u6_u0_n96 ) , .C2( u0_u6_u0_n97 ) , .ZN( u0_u6_u0_n98 ) );
  INV_X1 u0_u6_u0_U49 (.ZN( u0_u6_u0_n169 ) , .A( u0_u6_u0_n91 ) );
  NOR2_X1 u0_u6_u0_U5 (.A1( u0_u6_u0_n108 ) , .ZN( u0_u6_u0_n123 ) , .A2( u0_u6_u0_n158 ) );
  NOR2_X1 u0_u6_u0_U50 (.A2( u0_u6_X_4 ) , .A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n118 ) );
  NOR2_X1 u0_u6_u0_U51 (.A2( u0_u6_X_1 ) , .ZN( u0_u6_u0_n101 ) , .A1( u0_u6_u0_n163 ) );
  NAND2_X1 u0_u6_u0_U52 (.A2( u0_u6_X_4 ) , .A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n144 ) );
  NOR2_X1 u0_u6_u0_U53 (.A2( u0_u6_X_5 ) , .ZN( u0_u6_u0_n136 ) , .A1( u0_u6_u0_n159 ) );
  NAND2_X1 u0_u6_u0_U54 (.A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n138 ) , .A2( u0_u6_u0_n159 ) );
  AND2_X1 u0_u6_u0_U55 (.A2( u0_u6_X_3 ) , .A1( u0_u6_X_6 ) , .ZN( u0_u6_u0_n102 ) );
  INV_X1 u0_u6_u0_U56 (.A( u0_u6_X_4 ) , .ZN( u0_u6_u0_n159 ) );
  INV_X1 u0_u6_u0_U57 (.A( u0_u6_X_1 ) , .ZN( u0_u6_u0_n164 ) );
  INV_X1 u0_u6_u0_U58 (.A( u0_u6_X_3 ) , .ZN( u0_u6_u0_n162 ) );
  INV_X1 u0_u6_u0_U59 (.A( u0_u6_u0_n126 ) , .ZN( u0_u6_u0_n168 ) );
  AOI21_X1 u0_u6_u0_U6 (.B2( u0_u6_u0_n131 ) , .ZN( u0_u6_u0_n134 ) , .B1( u0_u6_u0_n151 ) , .A( u0_u6_u0_n158 ) );
  AOI211_X1 u0_u6_u0_U60 (.B( u0_u6_u0_n133 ) , .A( u0_u6_u0_n134 ) , .C2( u0_u6_u0_n135 ) , .C1( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n137 ) );
  INV_X1 u0_u6_u0_U61 (.ZN( u0_u6_u0_n174 ) , .A( u0_u6_u0_n89 ) );
  AOI211_X1 u0_u6_u0_U62 (.B( u0_u6_u0_n104 ) , .A( u0_u6_u0_n105 ) , .ZN( u0_u6_u0_n106 ) , .C2( u0_u6_u0_n113 ) , .C1( u0_u6_u0_n160 ) );
  OR4_X1 u0_u6_u0_U63 (.ZN( u0_out6_31 ) , .A4( u0_u6_u0_n155 ) , .A2( u0_u6_u0_n156 ) , .A1( u0_u6_u0_n157 ) , .A3( u0_u6_u0_n173 ) );
  AOI21_X1 u0_u6_u0_U64 (.A( u0_u6_u0_n138 ) , .B2( u0_u6_u0_n139 ) , .B1( u0_u6_u0_n140 ) , .ZN( u0_u6_u0_n157 ) );
  OR4_X1 u0_u6_u0_U65 (.ZN( u0_out6_17 ) , .A4( u0_u6_u0_n122 ) , .A2( u0_u6_u0_n123 ) , .A1( u0_u6_u0_n124 ) , .A3( u0_u6_u0_n170 ) );
  AOI21_X1 u0_u6_u0_U66 (.B2( u0_u6_u0_n107 ) , .ZN( u0_u6_u0_n124 ) , .B1( u0_u6_u0_n128 ) , .A( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U67 (.A( u0_u6_u0_n111 ) , .ZN( u0_u6_u0_n170 ) );
  AOI21_X1 u0_u6_u0_U68 (.B2( u0_u6_u0_n141 ) , .B1( u0_u6_u0_n142 ) , .ZN( u0_u6_u0_n156 ) , .A( u0_u6_u0_n161 ) );
  AOI21_X1 u0_u6_u0_U69 (.ZN( u0_u6_u0_n116 ) , .B2( u0_u6_u0_n142 ) , .A( u0_u6_u0_n144 ) , .B1( u0_u6_u0_n166 ) );
  OAI21_X1 u0_u6_u0_U7 (.B1( u0_u6_u0_n150 ) , .B2( u0_u6_u0_n158 ) , .A( u0_u6_u0_n172 ) , .ZN( u0_u6_u0_n89 ) );
  NAND2_X1 u0_u6_u0_U70 (.ZN( u0_u6_u0_n148 ) , .A1( u0_u6_u0_n93 ) , .A2( u0_u6_u0_n95 ) );
  NAND2_X1 u0_u6_u0_U71 (.A1( u0_u6_u0_n100 ) , .ZN( u0_u6_u0_n129 ) , .A2( u0_u6_u0_n95 ) );
  NAND2_X1 u0_u6_u0_U72 (.A1( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n128 ) , .A2( u0_u6_u0_n95 ) );
  INV_X1 u0_u6_u0_U73 (.A( u0_u6_u0_n142 ) , .ZN( u0_u6_u0_n165 ) );
  NOR2_X1 u0_u6_u0_U74 (.A2( u0_u6_X_1 ) , .A1( u0_u6_X_2 ) , .ZN( u0_u6_u0_n92 ) );
  NOR2_X1 u0_u6_u0_U75 (.A2( u0_u6_X_2 ) , .ZN( u0_u6_u0_n103 ) , .A1( u0_u6_u0_n164 ) );
  INV_X1 u0_u6_u0_U76 (.A( u0_u6_X_2 ) , .ZN( u0_u6_u0_n163 ) );
  AOI21_X1 u0_u6_u0_U77 (.B1( u0_u6_u0_n132 ) , .ZN( u0_u6_u0_n133 ) , .A( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n166 ) );
  OAI22_X1 u0_u6_u0_U78 (.ZN( u0_u6_u0_n105 ) , .A2( u0_u6_u0_n132 ) , .B1( u0_u6_u0_n146 ) , .A1( u0_u6_u0_n147 ) , .B2( u0_u6_u0_n161 ) );
  NAND2_X1 u0_u6_u0_U79 (.ZN( u0_u6_u0_n110 ) , .A2( u0_u6_u0_n132 ) , .A1( u0_u6_u0_n145 ) );
  AND2_X1 u0_u6_u0_U8 (.A1( u0_u6_u0_n114 ) , .A2( u0_u6_u0_n121 ) , .ZN( u0_u6_u0_n146 ) );
  INV_X1 u0_u6_u0_U80 (.A( u0_u6_u0_n119 ) , .ZN( u0_u6_u0_n167 ) );
  NAND2_X1 u0_u6_u0_U81 (.A2( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n140 ) , .A1( u0_u6_u0_n94 ) );
  NAND2_X1 u0_u6_u0_U82 (.A1( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n130 ) , .A2( u0_u6_u0_n94 ) );
  NAND2_X1 u0_u6_u0_U83 (.ZN( u0_u6_u0_n108 ) , .A1( u0_u6_u0_n92 ) , .A2( u0_u6_u0_n94 ) );
  AND2_X1 u0_u6_u0_U84 (.A1( u0_u6_X_6 ) , .A2( u0_u6_u0_n162 ) , .ZN( u0_u6_u0_n93 ) );
  NAND2_X1 u0_u6_u0_U85 (.ZN( u0_u6_u0_n142 ) , .A1( u0_u6_u0_n94 ) , .A2( u0_u6_u0_n95 ) );
  NOR2_X1 u0_u6_u0_U86 (.A2( u0_u6_X_6 ) , .ZN( u0_u6_u0_n100 ) , .A1( u0_u6_u0_n162 ) );
  NOR2_X1 u0_u6_u0_U87 (.A2( u0_u6_X_3 ) , .A1( u0_u6_X_6 ) , .ZN( u0_u6_u0_n94 ) );
  NAND3_X1 u0_u6_u0_U88 (.ZN( u0_out6_23 ) , .A3( u0_u6_u0_n137 ) , .A1( u0_u6_u0_n168 ) , .A2( u0_u6_u0_n171 ) );
  NAND3_X1 u0_u6_u0_U89 (.A3( u0_u6_u0_n127 ) , .A2( u0_u6_u0_n128 ) , .ZN( u0_u6_u0_n135 ) , .A1( u0_u6_u0_n150 ) );
  AND3_X1 u0_u6_u0_U9 (.A2( u0_u6_u0_n112 ) , .ZN( u0_u6_u0_n127 ) , .A3( u0_u6_u0_n130 ) , .A1( u0_u6_u0_n148 ) );
  NAND3_X1 u0_u6_u0_U90 (.ZN( u0_u6_u0_n117 ) , .A3( u0_u6_u0_n132 ) , .A2( u0_u6_u0_n139 ) , .A1( u0_u6_u0_n148 ) );
  NAND3_X1 u0_u6_u0_U91 (.ZN( u0_u6_u0_n109 ) , .A2( u0_u6_u0_n114 ) , .A3( u0_u6_u0_n140 ) , .A1( u0_u6_u0_n149 ) );
  NAND3_X1 u0_u6_u0_U92 (.ZN( u0_out6_9 ) , .A3( u0_u6_u0_n106 ) , .A2( u0_u6_u0_n171 ) , .A1( u0_u6_u0_n174 ) );
  NAND3_X1 u0_u6_u0_U93 (.A2( u0_u6_u0_n128 ) , .A1( u0_u6_u0_n132 ) , .A3( u0_u6_u0_n146 ) , .ZN( u0_u6_u0_n97 ) );
  AOI21_X1 u0_u6_u1_U10 (.B2( u0_u6_u1_n155 ) , .B1( u0_u6_u1_n156 ) , .ZN( u0_u6_u1_n157 ) , .A( u0_u6_u1_n174 ) );
  NAND3_X1 u0_u6_u1_U100 (.ZN( u0_u6_u1_n113 ) , .A1( u0_u6_u1_n120 ) , .A3( u0_u6_u1_n133 ) , .A2( u0_u6_u1_n155 ) );
  NAND2_X1 u0_u6_u1_U11 (.ZN( u0_u6_u1_n140 ) , .A2( u0_u6_u1_n150 ) , .A1( u0_u6_u1_n155 ) );
  NAND2_X1 u0_u6_u1_U12 (.A1( u0_u6_u1_n131 ) , .ZN( u0_u6_u1_n147 ) , .A2( u0_u6_u1_n153 ) );
  INV_X1 u0_u6_u1_U13 (.A( u0_u6_u1_n139 ) , .ZN( u0_u6_u1_n174 ) );
  OR4_X1 u0_u6_u1_U14 (.A4( u0_u6_u1_n106 ) , .A3( u0_u6_u1_n107 ) , .ZN( u0_u6_u1_n108 ) , .A1( u0_u6_u1_n117 ) , .A2( u0_u6_u1_n184 ) );
  AOI21_X1 u0_u6_u1_U15 (.ZN( u0_u6_u1_n106 ) , .A( u0_u6_u1_n112 ) , .B1( u0_u6_u1_n154 ) , .B2( u0_u6_u1_n156 ) );
  AOI21_X1 u0_u6_u1_U16 (.ZN( u0_u6_u1_n107 ) , .B1( u0_u6_u1_n134 ) , .B2( u0_u6_u1_n149 ) , .A( u0_u6_u1_n174 ) );
  INV_X1 u0_u6_u1_U17 (.A( u0_u6_u1_n101 ) , .ZN( u0_u6_u1_n184 ) );
  INV_X1 u0_u6_u1_U18 (.A( u0_u6_u1_n112 ) , .ZN( u0_u6_u1_n171 ) );
  NAND2_X1 u0_u6_u1_U19 (.ZN( u0_u6_u1_n141 ) , .A1( u0_u6_u1_n153 ) , .A2( u0_u6_u1_n156 ) );
  AND2_X1 u0_u6_u1_U20 (.A1( u0_u6_u1_n123 ) , .ZN( u0_u6_u1_n134 ) , .A2( u0_u6_u1_n161 ) );
  NAND2_X1 u0_u6_u1_U21 (.A2( u0_u6_u1_n115 ) , .A1( u0_u6_u1_n116 ) , .ZN( u0_u6_u1_n148 ) );
  NAND2_X1 u0_u6_u1_U22 (.A2( u0_u6_u1_n133 ) , .A1( u0_u6_u1_n135 ) , .ZN( u0_u6_u1_n159 ) );
  NAND2_X1 u0_u6_u1_U23 (.A2( u0_u6_u1_n115 ) , .A1( u0_u6_u1_n120 ) , .ZN( u0_u6_u1_n132 ) );
  INV_X1 u0_u6_u1_U24 (.A( u0_u6_u1_n154 ) , .ZN( u0_u6_u1_n178 ) );
  AOI22_X1 u0_u6_u1_U25 (.B2( u0_u6_u1_n113 ) , .A2( u0_u6_u1_n114 ) , .ZN( u0_u6_u1_n125 ) , .A1( u0_u6_u1_n171 ) , .B1( u0_u6_u1_n173 ) );
  NAND2_X1 u0_u6_u1_U26 (.ZN( u0_u6_u1_n114 ) , .A1( u0_u6_u1_n134 ) , .A2( u0_u6_u1_n156 ) );
  INV_X1 u0_u6_u1_U27 (.A( u0_u6_u1_n151 ) , .ZN( u0_u6_u1_n183 ) );
  AND2_X1 u0_u6_u1_U28 (.A1( u0_u6_u1_n129 ) , .A2( u0_u6_u1_n133 ) , .ZN( u0_u6_u1_n149 ) );
  INV_X1 u0_u6_u1_U29 (.A( u0_u6_u1_n131 ) , .ZN( u0_u6_u1_n180 ) );
  INV_X1 u0_u6_u1_U3 (.A( u0_u6_u1_n159 ) , .ZN( u0_u6_u1_n182 ) );
  AOI221_X1 u0_u6_u1_U30 (.B1( u0_u6_u1_n140 ) , .ZN( u0_u6_u1_n167 ) , .B2( u0_u6_u1_n172 ) , .C2( u0_u6_u1_n175 ) , .C1( u0_u6_u1_n178 ) , .A( u0_u6_u1_n188 ) );
  INV_X1 u0_u6_u1_U31 (.ZN( u0_u6_u1_n188 ) , .A( u0_u6_u1_n97 ) );
  AOI211_X1 u0_u6_u1_U32 (.A( u0_u6_u1_n118 ) , .C1( u0_u6_u1_n132 ) , .C2( u0_u6_u1_n139 ) , .B( u0_u6_u1_n96 ) , .ZN( u0_u6_u1_n97 ) );
  AOI21_X1 u0_u6_u1_U33 (.B2( u0_u6_u1_n121 ) , .B1( u0_u6_u1_n135 ) , .A( u0_u6_u1_n152 ) , .ZN( u0_u6_u1_n96 ) );
  OAI221_X1 u0_u6_u1_U34 (.A( u0_u6_u1_n119 ) , .C2( u0_u6_u1_n129 ) , .ZN( u0_u6_u1_n138 ) , .B2( u0_u6_u1_n152 ) , .C1( u0_u6_u1_n174 ) , .B1( u0_u6_u1_n187 ) );
  INV_X1 u0_u6_u1_U35 (.A( u0_u6_u1_n148 ) , .ZN( u0_u6_u1_n187 ) );
  AOI211_X1 u0_u6_u1_U36 (.B( u0_u6_u1_n117 ) , .A( u0_u6_u1_n118 ) , .ZN( u0_u6_u1_n119 ) , .C2( u0_u6_u1_n146 ) , .C1( u0_u6_u1_n159 ) );
  NOR2_X1 u0_u6_u1_U37 (.A1( u0_u6_u1_n168 ) , .A2( u0_u6_u1_n176 ) , .ZN( u0_u6_u1_n98 ) );
  AOI211_X1 u0_u6_u1_U38 (.B( u0_u6_u1_n162 ) , .A( u0_u6_u1_n163 ) , .C2( u0_u6_u1_n164 ) , .ZN( u0_u6_u1_n165 ) , .C1( u0_u6_u1_n171 ) );
  AOI21_X1 u0_u6_u1_U39 (.A( u0_u6_u1_n160 ) , .B2( u0_u6_u1_n161 ) , .ZN( u0_u6_u1_n162 ) , .B1( u0_u6_u1_n182 ) );
  AOI221_X1 u0_u6_u1_U4 (.A( u0_u6_u1_n138 ) , .C2( u0_u6_u1_n139 ) , .C1( u0_u6_u1_n140 ) , .B2( u0_u6_u1_n141 ) , .ZN( u0_u6_u1_n142 ) , .B1( u0_u6_u1_n175 ) );
  OR2_X1 u0_u6_u1_U40 (.A2( u0_u6_u1_n157 ) , .A1( u0_u6_u1_n158 ) , .ZN( u0_u6_u1_n163 ) );
  NAND2_X1 u0_u6_u1_U41 (.A1( u0_u6_u1_n128 ) , .ZN( u0_u6_u1_n146 ) , .A2( u0_u6_u1_n160 ) );
  NAND2_X1 u0_u6_u1_U42 (.A2( u0_u6_u1_n112 ) , .ZN( u0_u6_u1_n139 ) , .A1( u0_u6_u1_n152 ) );
  NAND2_X1 u0_u6_u1_U43 (.A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n156 ) , .A2( u0_u6_u1_n99 ) );
  NOR2_X1 u0_u6_u1_U44 (.ZN( u0_u6_u1_n117 ) , .A1( u0_u6_u1_n121 ) , .A2( u0_u6_u1_n160 ) );
  OAI21_X1 u0_u6_u1_U45 (.B2( u0_u6_u1_n123 ) , .ZN( u0_u6_u1_n145 ) , .B1( u0_u6_u1_n160 ) , .A( u0_u6_u1_n185 ) );
  INV_X1 u0_u6_u1_U46 (.A( u0_u6_u1_n122 ) , .ZN( u0_u6_u1_n185 ) );
  AOI21_X1 u0_u6_u1_U47 (.B2( u0_u6_u1_n120 ) , .B1( u0_u6_u1_n121 ) , .ZN( u0_u6_u1_n122 ) , .A( u0_u6_u1_n128 ) );
  AOI21_X1 u0_u6_u1_U48 (.A( u0_u6_u1_n128 ) , .B2( u0_u6_u1_n129 ) , .ZN( u0_u6_u1_n130 ) , .B1( u0_u6_u1_n150 ) );
  NAND2_X1 u0_u6_u1_U49 (.ZN( u0_u6_u1_n112 ) , .A1( u0_u6_u1_n169 ) , .A2( u0_u6_u1_n170 ) );
  AOI211_X1 u0_u6_u1_U5 (.ZN( u0_u6_u1_n124 ) , .A( u0_u6_u1_n138 ) , .C2( u0_u6_u1_n139 ) , .B( u0_u6_u1_n145 ) , .C1( u0_u6_u1_n147 ) );
  NAND2_X1 u0_u6_u1_U50 (.ZN( u0_u6_u1_n129 ) , .A2( u0_u6_u1_n95 ) , .A1( u0_u6_u1_n98 ) );
  NAND2_X1 u0_u6_u1_U51 (.A1( u0_u6_u1_n102 ) , .ZN( u0_u6_u1_n154 ) , .A2( u0_u6_u1_n99 ) );
  NAND2_X1 u0_u6_u1_U52 (.A2( u0_u6_u1_n100 ) , .ZN( u0_u6_u1_n135 ) , .A1( u0_u6_u1_n99 ) );
  AOI21_X1 u0_u6_u1_U53 (.A( u0_u6_u1_n152 ) , .B2( u0_u6_u1_n153 ) , .B1( u0_u6_u1_n154 ) , .ZN( u0_u6_u1_n158 ) );
  INV_X1 u0_u6_u1_U54 (.A( u0_u6_u1_n160 ) , .ZN( u0_u6_u1_n175 ) );
  NAND2_X1 u0_u6_u1_U55 (.A1( u0_u6_u1_n100 ) , .ZN( u0_u6_u1_n116 ) , .A2( u0_u6_u1_n95 ) );
  NAND2_X1 u0_u6_u1_U56 (.A1( u0_u6_u1_n102 ) , .ZN( u0_u6_u1_n131 ) , .A2( u0_u6_u1_n95 ) );
  NAND2_X1 u0_u6_u1_U57 (.A2( u0_u6_u1_n104 ) , .ZN( u0_u6_u1_n121 ) , .A1( u0_u6_u1_n98 ) );
  NAND2_X1 u0_u6_u1_U58 (.A1( u0_u6_u1_n103 ) , .ZN( u0_u6_u1_n153 ) , .A2( u0_u6_u1_n98 ) );
  NAND2_X1 u0_u6_u1_U59 (.A2( u0_u6_u1_n104 ) , .A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n133 ) );
  AOI22_X1 u0_u6_u1_U6 (.B2( u0_u6_u1_n136 ) , .A2( u0_u6_u1_n137 ) , .ZN( u0_u6_u1_n143 ) , .A1( u0_u6_u1_n171 ) , .B1( u0_u6_u1_n173 ) );
  NAND2_X1 u0_u6_u1_U60 (.ZN( u0_u6_u1_n150 ) , .A2( u0_u6_u1_n98 ) , .A1( u0_u6_u1_n99 ) );
  NAND2_X1 u0_u6_u1_U61 (.A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n155 ) , .A2( u0_u6_u1_n95 ) );
  OAI21_X1 u0_u6_u1_U62 (.ZN( u0_u6_u1_n109 ) , .B1( u0_u6_u1_n129 ) , .B2( u0_u6_u1_n160 ) , .A( u0_u6_u1_n167 ) );
  NAND2_X1 u0_u6_u1_U63 (.A2( u0_u6_u1_n100 ) , .A1( u0_u6_u1_n103 ) , .ZN( u0_u6_u1_n120 ) );
  NAND2_X1 u0_u6_u1_U64 (.A1( u0_u6_u1_n102 ) , .A2( u0_u6_u1_n104 ) , .ZN( u0_u6_u1_n115 ) );
  NAND2_X1 u0_u6_u1_U65 (.A2( u0_u6_u1_n100 ) , .A1( u0_u6_u1_n104 ) , .ZN( u0_u6_u1_n151 ) );
  NAND2_X1 u0_u6_u1_U66 (.A2( u0_u6_u1_n103 ) , .A1( u0_u6_u1_n105 ) , .ZN( u0_u6_u1_n161 ) );
  INV_X1 u0_u6_u1_U67 (.A( u0_u6_u1_n152 ) , .ZN( u0_u6_u1_n173 ) );
  INV_X1 u0_u6_u1_U68 (.A( u0_u6_u1_n128 ) , .ZN( u0_u6_u1_n172 ) );
  NAND2_X1 u0_u6_u1_U69 (.A2( u0_u6_u1_n102 ) , .A1( u0_u6_u1_n103 ) , .ZN( u0_u6_u1_n123 ) );
  INV_X1 u0_u6_u1_U7 (.A( u0_u6_u1_n147 ) , .ZN( u0_u6_u1_n181 ) );
  NOR2_X1 u0_u6_u1_U70 (.A2( u0_u6_X_7 ) , .A1( u0_u6_X_8 ) , .ZN( u0_u6_u1_n95 ) );
  NOR2_X1 u0_u6_u1_U71 (.A1( u0_u6_X_12 ) , .A2( u0_u6_X_9 ) , .ZN( u0_u6_u1_n100 ) );
  NOR2_X1 u0_u6_u1_U72 (.A2( u0_u6_X_8 ) , .A1( u0_u6_u1_n177 ) , .ZN( u0_u6_u1_n99 ) );
  NOR2_X1 u0_u6_u1_U73 (.A2( u0_u6_X_12 ) , .ZN( u0_u6_u1_n102 ) , .A1( u0_u6_u1_n176 ) );
  NOR2_X1 u0_u6_u1_U74 (.A2( u0_u6_X_9 ) , .ZN( u0_u6_u1_n105 ) , .A1( u0_u6_u1_n168 ) );
  NAND2_X1 u0_u6_u1_U75 (.A1( u0_u6_X_10 ) , .ZN( u0_u6_u1_n160 ) , .A2( u0_u6_u1_n169 ) );
  NAND2_X1 u0_u6_u1_U76 (.A2( u0_u6_X_10 ) , .A1( u0_u6_X_11 ) , .ZN( u0_u6_u1_n152 ) );
  NAND2_X1 u0_u6_u1_U77 (.A1( u0_u6_X_11 ) , .ZN( u0_u6_u1_n128 ) , .A2( u0_u6_u1_n170 ) );
  AND2_X1 u0_u6_u1_U78 (.A2( u0_u6_X_7 ) , .A1( u0_u6_X_8 ) , .ZN( u0_u6_u1_n104 ) );
  AND2_X1 u0_u6_u1_U79 (.A1( u0_u6_X_8 ) , .ZN( u0_u6_u1_n103 ) , .A2( u0_u6_u1_n177 ) );
  NOR2_X1 u0_u6_u1_U8 (.A1( u0_u6_u1_n112 ) , .A2( u0_u6_u1_n116 ) , .ZN( u0_u6_u1_n118 ) );
  INV_X1 u0_u6_u1_U80 (.A( u0_u6_X_10 ) , .ZN( u0_u6_u1_n170 ) );
  INV_X1 u0_u6_u1_U81 (.A( u0_u6_X_9 ) , .ZN( u0_u6_u1_n176 ) );
  INV_X1 u0_u6_u1_U82 (.A( u0_u6_X_11 ) , .ZN( u0_u6_u1_n169 ) );
  INV_X1 u0_u6_u1_U83 (.A( u0_u6_X_12 ) , .ZN( u0_u6_u1_n168 ) );
  INV_X1 u0_u6_u1_U84 (.A( u0_u6_X_7 ) , .ZN( u0_u6_u1_n177 ) );
  NAND4_X1 u0_u6_u1_U85 (.ZN( u0_out6_28 ) , .A4( u0_u6_u1_n124 ) , .A3( u0_u6_u1_n125 ) , .A2( u0_u6_u1_n126 ) , .A1( u0_u6_u1_n127 ) );
  OAI21_X1 u0_u6_u1_U86 (.ZN( u0_u6_u1_n127 ) , .B2( u0_u6_u1_n139 ) , .B1( u0_u6_u1_n175 ) , .A( u0_u6_u1_n183 ) );
  OAI21_X1 u0_u6_u1_U87 (.ZN( u0_u6_u1_n126 ) , .B2( u0_u6_u1_n140 ) , .A( u0_u6_u1_n146 ) , .B1( u0_u6_u1_n178 ) );
  NAND4_X1 u0_u6_u1_U88 (.ZN( u0_out6_18 ) , .A4( u0_u6_u1_n165 ) , .A3( u0_u6_u1_n166 ) , .A1( u0_u6_u1_n167 ) , .A2( u0_u6_u1_n186 ) );
  AOI22_X1 u0_u6_u1_U89 (.B2( u0_u6_u1_n146 ) , .B1( u0_u6_u1_n147 ) , .A2( u0_u6_u1_n148 ) , .ZN( u0_u6_u1_n166 ) , .A1( u0_u6_u1_n172 ) );
  OAI21_X1 u0_u6_u1_U9 (.ZN( u0_u6_u1_n101 ) , .B1( u0_u6_u1_n141 ) , .A( u0_u6_u1_n146 ) , .B2( u0_u6_u1_n183 ) );
  INV_X1 u0_u6_u1_U90 (.A( u0_u6_u1_n145 ) , .ZN( u0_u6_u1_n186 ) );
  NAND4_X1 u0_u6_u1_U91 (.ZN( u0_out6_2 ) , .A4( u0_u6_u1_n142 ) , .A3( u0_u6_u1_n143 ) , .A2( u0_u6_u1_n144 ) , .A1( u0_u6_u1_n179 ) );
  OAI21_X1 u0_u6_u1_U92 (.B2( u0_u6_u1_n132 ) , .ZN( u0_u6_u1_n144 ) , .A( u0_u6_u1_n146 ) , .B1( u0_u6_u1_n180 ) );
  INV_X1 u0_u6_u1_U93 (.A( u0_u6_u1_n130 ) , .ZN( u0_u6_u1_n179 ) );
  OR4_X1 u0_u6_u1_U94 (.ZN( u0_out6_13 ) , .A4( u0_u6_u1_n108 ) , .A3( u0_u6_u1_n109 ) , .A2( u0_u6_u1_n110 ) , .A1( u0_u6_u1_n111 ) );
  AOI21_X1 u0_u6_u1_U95 (.ZN( u0_u6_u1_n111 ) , .A( u0_u6_u1_n128 ) , .B2( u0_u6_u1_n131 ) , .B1( u0_u6_u1_n135 ) );
  AOI21_X1 u0_u6_u1_U96 (.ZN( u0_u6_u1_n110 ) , .A( u0_u6_u1_n116 ) , .B1( u0_u6_u1_n152 ) , .B2( u0_u6_u1_n160 ) );
  NAND3_X1 u0_u6_u1_U97 (.A3( u0_u6_u1_n149 ) , .A2( u0_u6_u1_n150 ) , .A1( u0_u6_u1_n151 ) , .ZN( u0_u6_u1_n164 ) );
  NAND3_X1 u0_u6_u1_U98 (.A3( u0_u6_u1_n134 ) , .A2( u0_u6_u1_n135 ) , .ZN( u0_u6_u1_n136 ) , .A1( u0_u6_u1_n151 ) );
  NAND3_X1 u0_u6_u1_U99 (.A1( u0_u6_u1_n133 ) , .ZN( u0_u6_u1_n137 ) , .A2( u0_u6_u1_n154 ) , .A3( u0_u6_u1_n181 ) );
  OAI22_X1 u0_u6_u2_U10 (.B1( u0_u6_u2_n151 ) , .A2( u0_u6_u2_n152 ) , .A1( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n160 ) , .B2( u0_u6_u2_n168 ) );
  NAND3_X1 u0_u6_u2_U100 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n104 ) , .A3( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n98 ) );
  NOR3_X1 u0_u6_u2_U11 (.A1( u0_u6_u2_n150 ) , .ZN( u0_u6_u2_n151 ) , .A3( u0_u6_u2_n175 ) , .A2( u0_u6_u2_n188 ) );
  AOI21_X1 u0_u6_u2_U12 (.B2( u0_u6_u2_n123 ) , .ZN( u0_u6_u2_n125 ) , .A( u0_u6_u2_n171 ) , .B1( u0_u6_u2_n184 ) );
  INV_X1 u0_u6_u2_U13 (.A( u0_u6_u2_n150 ) , .ZN( u0_u6_u2_n184 ) );
  AOI21_X1 u0_u6_u2_U14 (.ZN( u0_u6_u2_n144 ) , .B2( u0_u6_u2_n155 ) , .A( u0_u6_u2_n172 ) , .B1( u0_u6_u2_n185 ) );
  AOI21_X1 u0_u6_u2_U15 (.B2( u0_u6_u2_n143 ) , .ZN( u0_u6_u2_n145 ) , .B1( u0_u6_u2_n152 ) , .A( u0_u6_u2_n171 ) );
  INV_X1 u0_u6_u2_U16 (.A( u0_u6_u2_n156 ) , .ZN( u0_u6_u2_n171 ) );
  INV_X1 u0_u6_u2_U17 (.A( u0_u6_u2_n120 ) , .ZN( u0_u6_u2_n188 ) );
  NAND2_X1 u0_u6_u2_U18 (.A2( u0_u6_u2_n122 ) , .ZN( u0_u6_u2_n150 ) , .A1( u0_u6_u2_n152 ) );
  INV_X1 u0_u6_u2_U19 (.A( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n170 ) );
  INV_X1 u0_u6_u2_U20 (.A( u0_u6_u2_n137 ) , .ZN( u0_u6_u2_n173 ) );
  NAND2_X1 u0_u6_u2_U21 (.A1( u0_u6_u2_n132 ) , .A2( u0_u6_u2_n139 ) , .ZN( u0_u6_u2_n157 ) );
  INV_X1 u0_u6_u2_U22 (.A( u0_u6_u2_n113 ) , .ZN( u0_u6_u2_n178 ) );
  INV_X1 u0_u6_u2_U23 (.A( u0_u6_u2_n139 ) , .ZN( u0_u6_u2_n175 ) );
  INV_X1 u0_u6_u2_U24 (.A( u0_u6_u2_n155 ) , .ZN( u0_u6_u2_n181 ) );
  INV_X1 u0_u6_u2_U25 (.A( u0_u6_u2_n119 ) , .ZN( u0_u6_u2_n177 ) );
  INV_X1 u0_u6_u2_U26 (.A( u0_u6_u2_n116 ) , .ZN( u0_u6_u2_n180 ) );
  INV_X1 u0_u6_u2_U27 (.A( u0_u6_u2_n131 ) , .ZN( u0_u6_u2_n179 ) );
  INV_X1 u0_u6_u2_U28 (.A( u0_u6_u2_n154 ) , .ZN( u0_u6_u2_n176 ) );
  NAND2_X1 u0_u6_u2_U29 (.A2( u0_u6_u2_n116 ) , .A1( u0_u6_u2_n117 ) , .ZN( u0_u6_u2_n118 ) );
  NOR2_X1 u0_u6_u2_U3 (.ZN( u0_u6_u2_n121 ) , .A2( u0_u6_u2_n177 ) , .A1( u0_u6_u2_n180 ) );
  INV_X1 u0_u6_u2_U30 (.A( u0_u6_u2_n132 ) , .ZN( u0_u6_u2_n182 ) );
  INV_X1 u0_u6_u2_U31 (.A( u0_u6_u2_n158 ) , .ZN( u0_u6_u2_n183 ) );
  OAI21_X1 u0_u6_u2_U32 (.A( u0_u6_u2_n156 ) , .B1( u0_u6_u2_n157 ) , .ZN( u0_u6_u2_n158 ) , .B2( u0_u6_u2_n179 ) );
  NOR2_X1 u0_u6_u2_U33 (.ZN( u0_u6_u2_n156 ) , .A1( u0_u6_u2_n166 ) , .A2( u0_u6_u2_n169 ) );
  NOR2_X1 u0_u6_u2_U34 (.A2( u0_u6_u2_n114 ) , .ZN( u0_u6_u2_n137 ) , .A1( u0_u6_u2_n140 ) );
  NOR2_X1 u0_u6_u2_U35 (.A2( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n153 ) , .A1( u0_u6_u2_n156 ) );
  AOI211_X1 u0_u6_u2_U36 (.ZN( u0_u6_u2_n130 ) , .C1( u0_u6_u2_n138 ) , .C2( u0_u6_u2_n179 ) , .B( u0_u6_u2_n96 ) , .A( u0_u6_u2_n97 ) );
  OAI22_X1 u0_u6_u2_U37 (.B1( u0_u6_u2_n133 ) , .A2( u0_u6_u2_n137 ) , .A1( u0_u6_u2_n152 ) , .B2( u0_u6_u2_n168 ) , .ZN( u0_u6_u2_n97 ) );
  OAI221_X1 u0_u6_u2_U38 (.B1( u0_u6_u2_n113 ) , .C1( u0_u6_u2_n132 ) , .A( u0_u6_u2_n149 ) , .B2( u0_u6_u2_n171 ) , .C2( u0_u6_u2_n172 ) , .ZN( u0_u6_u2_n96 ) );
  OAI221_X1 u0_u6_u2_U39 (.A( u0_u6_u2_n115 ) , .C2( u0_u6_u2_n123 ) , .B2( u0_u6_u2_n143 ) , .B1( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n163 ) , .C1( u0_u6_u2_n168 ) );
  INV_X1 u0_u6_u2_U4 (.A( u0_u6_u2_n134 ) , .ZN( u0_u6_u2_n185 ) );
  OAI21_X1 u0_u6_u2_U40 (.A( u0_u6_u2_n114 ) , .ZN( u0_u6_u2_n115 ) , .B1( u0_u6_u2_n176 ) , .B2( u0_u6_u2_n178 ) );
  OAI221_X1 u0_u6_u2_U41 (.A( u0_u6_u2_n135 ) , .B2( u0_u6_u2_n136 ) , .B1( u0_u6_u2_n137 ) , .ZN( u0_u6_u2_n162 ) , .C2( u0_u6_u2_n167 ) , .C1( u0_u6_u2_n185 ) );
  AND3_X1 u0_u6_u2_U42 (.A3( u0_u6_u2_n131 ) , .A2( u0_u6_u2_n132 ) , .A1( u0_u6_u2_n133 ) , .ZN( u0_u6_u2_n136 ) );
  AOI22_X1 u0_u6_u2_U43 (.ZN( u0_u6_u2_n135 ) , .B1( u0_u6_u2_n140 ) , .A1( u0_u6_u2_n156 ) , .B2( u0_u6_u2_n180 ) , .A2( u0_u6_u2_n188 ) );
  AOI21_X1 u0_u6_u2_U44 (.ZN( u0_u6_u2_n149 ) , .B1( u0_u6_u2_n173 ) , .B2( u0_u6_u2_n188 ) , .A( u0_u6_u2_n95 ) );
  AND3_X1 u0_u6_u2_U45 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n104 ) , .A3( u0_u6_u2_n156 ) , .ZN( u0_u6_u2_n95 ) );
  OAI21_X1 u0_u6_u2_U46 (.A( u0_u6_u2_n141 ) , .B2( u0_u6_u2_n142 ) , .ZN( u0_u6_u2_n146 ) , .B1( u0_u6_u2_n153 ) );
  OAI21_X1 u0_u6_u2_U47 (.A( u0_u6_u2_n140 ) , .ZN( u0_u6_u2_n141 ) , .B1( u0_u6_u2_n176 ) , .B2( u0_u6_u2_n177 ) );
  NOR3_X1 u0_u6_u2_U48 (.ZN( u0_u6_u2_n142 ) , .A3( u0_u6_u2_n175 ) , .A2( u0_u6_u2_n178 ) , .A1( u0_u6_u2_n181 ) );
  OAI21_X1 u0_u6_u2_U49 (.A( u0_u6_u2_n101 ) , .B2( u0_u6_u2_n121 ) , .B1( u0_u6_u2_n153 ) , .ZN( u0_u6_u2_n164 ) );
  NOR4_X1 u0_u6_u2_U5 (.A4( u0_u6_u2_n124 ) , .A3( u0_u6_u2_n125 ) , .A2( u0_u6_u2_n126 ) , .A1( u0_u6_u2_n127 ) , .ZN( u0_u6_u2_n128 ) );
  NAND2_X1 u0_u6_u2_U50 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n107 ) , .ZN( u0_u6_u2_n155 ) );
  NAND2_X1 u0_u6_u2_U51 (.A2( u0_u6_u2_n105 ) , .A1( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n143 ) );
  NAND2_X1 u0_u6_u2_U52 (.A1( u0_u6_u2_n104 ) , .A2( u0_u6_u2_n106 ) , .ZN( u0_u6_u2_n152 ) );
  NAND2_X1 u0_u6_u2_U53 (.A1( u0_u6_u2_n100 ) , .A2( u0_u6_u2_n105 ) , .ZN( u0_u6_u2_n132 ) );
  INV_X1 u0_u6_u2_U54 (.A( u0_u6_u2_n140 ) , .ZN( u0_u6_u2_n168 ) );
  INV_X1 u0_u6_u2_U55 (.A( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n167 ) );
  INV_X1 u0_u6_u2_U56 (.ZN( u0_u6_u2_n187 ) , .A( u0_u6_u2_n99 ) );
  OAI21_X1 u0_u6_u2_U57 (.B1( u0_u6_u2_n137 ) , .B2( u0_u6_u2_n143 ) , .A( u0_u6_u2_n98 ) , .ZN( u0_u6_u2_n99 ) );
  NAND2_X1 u0_u6_u2_U58 (.A1( u0_u6_u2_n102 ) , .A2( u0_u6_u2_n106 ) , .ZN( u0_u6_u2_n113 ) );
  NAND2_X1 u0_u6_u2_U59 (.A1( u0_u6_u2_n106 ) , .A2( u0_u6_u2_n107 ) , .ZN( u0_u6_u2_n131 ) );
  AOI21_X1 u0_u6_u2_U6 (.B2( u0_u6_u2_n119 ) , .ZN( u0_u6_u2_n127 ) , .A( u0_u6_u2_n137 ) , .B1( u0_u6_u2_n155 ) );
  NAND2_X1 u0_u6_u2_U60 (.A1( u0_u6_u2_n103 ) , .A2( u0_u6_u2_n107 ) , .ZN( u0_u6_u2_n139 ) );
  NAND2_X1 u0_u6_u2_U61 (.A1( u0_u6_u2_n103 ) , .A2( u0_u6_u2_n105 ) , .ZN( u0_u6_u2_n133 ) );
  NAND2_X1 u0_u6_u2_U62 (.A1( u0_u6_u2_n102 ) , .A2( u0_u6_u2_n103 ) , .ZN( u0_u6_u2_n154 ) );
  NAND2_X1 u0_u6_u2_U63 (.A2( u0_u6_u2_n103 ) , .A1( u0_u6_u2_n104 ) , .ZN( u0_u6_u2_n119 ) );
  NAND2_X1 u0_u6_u2_U64 (.A2( u0_u6_u2_n107 ) , .A1( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n123 ) );
  NAND2_X1 u0_u6_u2_U65 (.A1( u0_u6_u2_n104 ) , .A2( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n122 ) );
  INV_X1 u0_u6_u2_U66 (.A( u0_u6_u2_n114 ) , .ZN( u0_u6_u2_n172 ) );
  NAND2_X1 u0_u6_u2_U67 (.A2( u0_u6_u2_n100 ) , .A1( u0_u6_u2_n102 ) , .ZN( u0_u6_u2_n116 ) );
  NAND2_X1 u0_u6_u2_U68 (.A1( u0_u6_u2_n102 ) , .A2( u0_u6_u2_n108 ) , .ZN( u0_u6_u2_n120 ) );
  NAND2_X1 u0_u6_u2_U69 (.A2( u0_u6_u2_n105 ) , .A1( u0_u6_u2_n106 ) , .ZN( u0_u6_u2_n117 ) );
  AOI21_X1 u0_u6_u2_U7 (.ZN( u0_u6_u2_n124 ) , .B1( u0_u6_u2_n131 ) , .B2( u0_u6_u2_n143 ) , .A( u0_u6_u2_n172 ) );
  NOR2_X1 u0_u6_u2_U70 (.A2( u0_u6_X_16 ) , .ZN( u0_u6_u2_n140 ) , .A1( u0_u6_u2_n166 ) );
  NOR2_X1 u0_u6_u2_U71 (.A2( u0_u6_X_13 ) , .A1( u0_u6_X_14 ) , .ZN( u0_u6_u2_n100 ) );
  NOR2_X1 u0_u6_u2_U72 (.A2( u0_u6_X_16 ) , .A1( u0_u6_X_17 ) , .ZN( u0_u6_u2_n138 ) );
  NOR2_X1 u0_u6_u2_U73 (.A2( u0_u6_X_15 ) , .A1( u0_u6_X_18 ) , .ZN( u0_u6_u2_n104 ) );
  NOR2_X1 u0_u6_u2_U74 (.A2( u0_u6_X_14 ) , .ZN( u0_u6_u2_n103 ) , .A1( u0_u6_u2_n174 ) );
  NOR2_X1 u0_u6_u2_U75 (.A2( u0_u6_X_15 ) , .ZN( u0_u6_u2_n102 ) , .A1( u0_u6_u2_n165 ) );
  NOR2_X1 u0_u6_u2_U76 (.A2( u0_u6_X_17 ) , .ZN( u0_u6_u2_n114 ) , .A1( u0_u6_u2_n169 ) );
  AND2_X1 u0_u6_u2_U77 (.A1( u0_u6_X_15 ) , .ZN( u0_u6_u2_n105 ) , .A2( u0_u6_u2_n165 ) );
  AND2_X1 u0_u6_u2_U78 (.A2( u0_u6_X_15 ) , .A1( u0_u6_X_18 ) , .ZN( u0_u6_u2_n107 ) );
  AND2_X1 u0_u6_u2_U79 (.A1( u0_u6_X_14 ) , .ZN( u0_u6_u2_n106 ) , .A2( u0_u6_u2_n174 ) );
  AOI21_X1 u0_u6_u2_U8 (.B2( u0_u6_u2_n120 ) , .B1( u0_u6_u2_n121 ) , .ZN( u0_u6_u2_n126 ) , .A( u0_u6_u2_n167 ) );
  AND2_X1 u0_u6_u2_U80 (.A1( u0_u6_X_13 ) , .A2( u0_u6_X_14 ) , .ZN( u0_u6_u2_n108 ) );
  INV_X1 u0_u6_u2_U81 (.A( u0_u6_X_16 ) , .ZN( u0_u6_u2_n169 ) );
  INV_X1 u0_u6_u2_U82 (.A( u0_u6_X_17 ) , .ZN( u0_u6_u2_n166 ) );
  INV_X1 u0_u6_u2_U83 (.A( u0_u6_X_13 ) , .ZN( u0_u6_u2_n174 ) );
  INV_X1 u0_u6_u2_U84 (.A( u0_u6_X_18 ) , .ZN( u0_u6_u2_n165 ) );
  NAND4_X1 u0_u6_u2_U85 (.ZN( u0_out6_30 ) , .A4( u0_u6_u2_n147 ) , .A3( u0_u6_u2_n148 ) , .A2( u0_u6_u2_n149 ) , .A1( u0_u6_u2_n187 ) );
  AOI21_X1 u0_u6_u2_U86 (.B2( u0_u6_u2_n138 ) , .ZN( u0_u6_u2_n148 ) , .A( u0_u6_u2_n162 ) , .B1( u0_u6_u2_n182 ) );
  NOR3_X1 u0_u6_u2_U87 (.A3( u0_u6_u2_n144 ) , .A2( u0_u6_u2_n145 ) , .A1( u0_u6_u2_n146 ) , .ZN( u0_u6_u2_n147 ) );
  NAND4_X1 u0_u6_u2_U88 (.ZN( u0_out6_24 ) , .A4( u0_u6_u2_n111 ) , .A3( u0_u6_u2_n112 ) , .A1( u0_u6_u2_n130 ) , .A2( u0_u6_u2_n187 ) );
  AOI221_X1 u0_u6_u2_U89 (.A( u0_u6_u2_n109 ) , .B1( u0_u6_u2_n110 ) , .ZN( u0_u6_u2_n111 ) , .C1( u0_u6_u2_n134 ) , .C2( u0_u6_u2_n170 ) , .B2( u0_u6_u2_n173 ) );
  OAI22_X1 u0_u6_u2_U9 (.ZN( u0_u6_u2_n109 ) , .A2( u0_u6_u2_n113 ) , .B2( u0_u6_u2_n133 ) , .B1( u0_u6_u2_n167 ) , .A1( u0_u6_u2_n168 ) );
  AOI21_X1 u0_u6_u2_U90 (.ZN( u0_u6_u2_n112 ) , .B2( u0_u6_u2_n156 ) , .A( u0_u6_u2_n164 ) , .B1( u0_u6_u2_n181 ) );
  NAND4_X1 u0_u6_u2_U91 (.ZN( u0_out6_16 ) , .A4( u0_u6_u2_n128 ) , .A3( u0_u6_u2_n129 ) , .A1( u0_u6_u2_n130 ) , .A2( u0_u6_u2_n186 ) );
  AOI22_X1 u0_u6_u2_U92 (.A2( u0_u6_u2_n118 ) , .ZN( u0_u6_u2_n129 ) , .A1( u0_u6_u2_n140 ) , .B1( u0_u6_u2_n157 ) , .B2( u0_u6_u2_n170 ) );
  INV_X1 u0_u6_u2_U93 (.A( u0_u6_u2_n163 ) , .ZN( u0_u6_u2_n186 ) );
  OR4_X1 u0_u6_u2_U94 (.ZN( u0_out6_6 ) , .A4( u0_u6_u2_n161 ) , .A3( u0_u6_u2_n162 ) , .A2( u0_u6_u2_n163 ) , .A1( u0_u6_u2_n164 ) );
  OR3_X1 u0_u6_u2_U95 (.A2( u0_u6_u2_n159 ) , .A1( u0_u6_u2_n160 ) , .ZN( u0_u6_u2_n161 ) , .A3( u0_u6_u2_n183 ) );
  AOI21_X1 u0_u6_u2_U96 (.B2( u0_u6_u2_n154 ) , .B1( u0_u6_u2_n155 ) , .ZN( u0_u6_u2_n159 ) , .A( u0_u6_u2_n167 ) );
  NAND3_X1 u0_u6_u2_U97 (.A2( u0_u6_u2_n117 ) , .A1( u0_u6_u2_n122 ) , .A3( u0_u6_u2_n123 ) , .ZN( u0_u6_u2_n134 ) );
  NAND3_X1 u0_u6_u2_U98 (.ZN( u0_u6_u2_n110 ) , .A2( u0_u6_u2_n131 ) , .A3( u0_u6_u2_n139 ) , .A1( u0_u6_u2_n154 ) );
  NAND3_X1 u0_u6_u2_U99 (.A2( u0_u6_u2_n100 ) , .ZN( u0_u6_u2_n101 ) , .A1( u0_u6_u2_n104 ) , .A3( u0_u6_u2_n114 ) );
  OAI22_X1 u0_u6_u3_U10 (.B1( u0_u6_u3_n113 ) , .A2( u0_u6_u3_n135 ) , .A1( u0_u6_u3_n150 ) , .B2( u0_u6_u3_n164 ) , .ZN( u0_u6_u3_n98 ) );
  OAI211_X1 u0_u6_u3_U11 (.B( u0_u6_u3_n106 ) , .ZN( u0_u6_u3_n119 ) , .C2( u0_u6_u3_n128 ) , .C1( u0_u6_u3_n167 ) , .A( u0_u6_u3_n181 ) );
  AOI221_X1 u0_u6_u3_U12 (.C1( u0_u6_u3_n105 ) , .ZN( u0_u6_u3_n106 ) , .A( u0_u6_u3_n131 ) , .B2( u0_u6_u3_n132 ) , .C2( u0_u6_u3_n133 ) , .B1( u0_u6_u3_n169 ) );
  INV_X1 u0_u6_u3_U13 (.ZN( u0_u6_u3_n181 ) , .A( u0_u6_u3_n98 ) );
  NAND2_X1 u0_u6_u3_U14 (.ZN( u0_u6_u3_n105 ) , .A2( u0_u6_u3_n130 ) , .A1( u0_u6_u3_n155 ) );
  NOR2_X1 u0_u6_u3_U15 (.ZN( u0_u6_u3_n126 ) , .A2( u0_u6_u3_n150 ) , .A1( u0_u6_u3_n164 ) );
  AOI21_X1 u0_u6_u3_U16 (.ZN( u0_u6_u3_n112 ) , .B2( u0_u6_u3_n146 ) , .B1( u0_u6_u3_n155 ) , .A( u0_u6_u3_n167 ) );
  NAND2_X1 u0_u6_u3_U17 (.A1( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n142 ) , .A2( u0_u6_u3_n164 ) );
  NAND2_X1 u0_u6_u3_U18 (.ZN( u0_u6_u3_n132 ) , .A2( u0_u6_u3_n152 ) , .A1( u0_u6_u3_n156 ) );
  AND2_X1 u0_u6_u3_U19 (.A2( u0_u6_u3_n113 ) , .A1( u0_u6_u3_n114 ) , .ZN( u0_u6_u3_n151 ) );
  INV_X1 u0_u6_u3_U20 (.A( u0_u6_u3_n133 ) , .ZN( u0_u6_u3_n165 ) );
  INV_X1 u0_u6_u3_U21 (.A( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n170 ) );
  NAND2_X1 u0_u6_u3_U22 (.A1( u0_u6_u3_n107 ) , .A2( u0_u6_u3_n108 ) , .ZN( u0_u6_u3_n140 ) );
  NAND2_X1 u0_u6_u3_U23 (.ZN( u0_u6_u3_n117 ) , .A1( u0_u6_u3_n124 ) , .A2( u0_u6_u3_n148 ) );
  NAND2_X1 u0_u6_u3_U24 (.ZN( u0_u6_u3_n143 ) , .A1( u0_u6_u3_n165 ) , .A2( u0_u6_u3_n167 ) );
  INV_X1 u0_u6_u3_U25 (.A( u0_u6_u3_n130 ) , .ZN( u0_u6_u3_n177 ) );
  INV_X1 u0_u6_u3_U26 (.A( u0_u6_u3_n128 ) , .ZN( u0_u6_u3_n176 ) );
  INV_X1 u0_u6_u3_U27 (.A( u0_u6_u3_n155 ) , .ZN( u0_u6_u3_n174 ) );
  AOI22_X1 u0_u6_u3_U28 (.B1( u0_u6_u3_n115 ) , .A2( u0_u6_u3_n116 ) , .ZN( u0_u6_u3_n123 ) , .B2( u0_u6_u3_n133 ) , .A1( u0_u6_u3_n169 ) );
  NAND2_X1 u0_u6_u3_U29 (.ZN( u0_u6_u3_n116 ) , .A2( u0_u6_u3_n151 ) , .A1( u0_u6_u3_n182 ) );
  INV_X1 u0_u6_u3_U3 (.A( u0_u6_u3_n129 ) , .ZN( u0_u6_u3_n183 ) );
  INV_X1 u0_u6_u3_U30 (.A( u0_u6_u3_n139 ) , .ZN( u0_u6_u3_n185 ) );
  NOR2_X1 u0_u6_u3_U31 (.ZN( u0_u6_u3_n135 ) , .A2( u0_u6_u3_n141 ) , .A1( u0_u6_u3_n169 ) );
  OAI222_X1 u0_u6_u3_U32 (.C2( u0_u6_u3_n107 ) , .A2( u0_u6_u3_n108 ) , .B1( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n138 ) , .B2( u0_u6_u3_n146 ) , .C1( u0_u6_u3_n154 ) , .A1( u0_u6_u3_n164 ) );
  NOR4_X1 u0_u6_u3_U33 (.A4( u0_u6_u3_n157 ) , .A3( u0_u6_u3_n158 ) , .A2( u0_u6_u3_n159 ) , .A1( u0_u6_u3_n160 ) , .ZN( u0_u6_u3_n161 ) );
  AOI21_X1 u0_u6_u3_U34 (.B2( u0_u6_u3_n152 ) , .B1( u0_u6_u3_n153 ) , .ZN( u0_u6_u3_n158 ) , .A( u0_u6_u3_n164 ) );
  AOI21_X1 u0_u6_u3_U35 (.A( u0_u6_u3_n154 ) , .B2( u0_u6_u3_n155 ) , .B1( u0_u6_u3_n156 ) , .ZN( u0_u6_u3_n157 ) );
  AOI21_X1 u0_u6_u3_U36 (.A( u0_u6_u3_n149 ) , .B2( u0_u6_u3_n150 ) , .B1( u0_u6_u3_n151 ) , .ZN( u0_u6_u3_n159 ) );
  AOI211_X1 u0_u6_u3_U37 (.ZN( u0_u6_u3_n109 ) , .A( u0_u6_u3_n119 ) , .C2( u0_u6_u3_n129 ) , .B( u0_u6_u3_n138 ) , .C1( u0_u6_u3_n141 ) );
  AOI211_X1 u0_u6_u3_U38 (.B( u0_u6_u3_n119 ) , .A( u0_u6_u3_n120 ) , .C2( u0_u6_u3_n121 ) , .ZN( u0_u6_u3_n122 ) , .C1( u0_u6_u3_n179 ) );
  INV_X1 u0_u6_u3_U39 (.A( u0_u6_u3_n156 ) , .ZN( u0_u6_u3_n179 ) );
  INV_X1 u0_u6_u3_U4 (.A( u0_u6_u3_n140 ) , .ZN( u0_u6_u3_n182 ) );
  OAI22_X1 u0_u6_u3_U40 (.B1( u0_u6_u3_n118 ) , .ZN( u0_u6_u3_n120 ) , .A1( u0_u6_u3_n135 ) , .B2( u0_u6_u3_n154 ) , .A2( u0_u6_u3_n178 ) );
  AND3_X1 u0_u6_u3_U41 (.ZN( u0_u6_u3_n118 ) , .A2( u0_u6_u3_n124 ) , .A1( u0_u6_u3_n144 ) , .A3( u0_u6_u3_n152 ) );
  INV_X1 u0_u6_u3_U42 (.A( u0_u6_u3_n121 ) , .ZN( u0_u6_u3_n164 ) );
  NAND2_X1 u0_u6_u3_U43 (.ZN( u0_u6_u3_n133 ) , .A1( u0_u6_u3_n154 ) , .A2( u0_u6_u3_n164 ) );
  OAI211_X1 u0_u6_u3_U44 (.B( u0_u6_u3_n127 ) , .ZN( u0_u6_u3_n139 ) , .C1( u0_u6_u3_n150 ) , .C2( u0_u6_u3_n154 ) , .A( u0_u6_u3_n184 ) );
  INV_X1 u0_u6_u3_U45 (.A( u0_u6_u3_n125 ) , .ZN( u0_u6_u3_n184 ) );
  AOI221_X1 u0_u6_u3_U46 (.A( u0_u6_u3_n126 ) , .ZN( u0_u6_u3_n127 ) , .C2( u0_u6_u3_n132 ) , .C1( u0_u6_u3_n169 ) , .B2( u0_u6_u3_n170 ) , .B1( u0_u6_u3_n174 ) );
  OAI22_X1 u0_u6_u3_U47 (.A1( u0_u6_u3_n124 ) , .ZN( u0_u6_u3_n125 ) , .B2( u0_u6_u3_n145 ) , .A2( u0_u6_u3_n165 ) , .B1( u0_u6_u3_n167 ) );
  NOR2_X1 u0_u6_u3_U48 (.A1( u0_u6_u3_n113 ) , .ZN( u0_u6_u3_n131 ) , .A2( u0_u6_u3_n154 ) );
  NAND2_X1 u0_u6_u3_U49 (.A1( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n150 ) , .A2( u0_u6_u3_n99 ) );
  INV_X1 u0_u6_u3_U5 (.A( u0_u6_u3_n117 ) , .ZN( u0_u6_u3_n178 ) );
  NAND2_X1 u0_u6_u3_U50 (.A2( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n155 ) , .A1( u0_u6_u3_n97 ) );
  INV_X1 u0_u6_u3_U51 (.A( u0_u6_u3_n141 ) , .ZN( u0_u6_u3_n167 ) );
  AOI21_X1 u0_u6_u3_U52 (.B2( u0_u6_u3_n114 ) , .B1( u0_u6_u3_n146 ) , .A( u0_u6_u3_n154 ) , .ZN( u0_u6_u3_n94 ) );
  AOI21_X1 u0_u6_u3_U53 (.ZN( u0_u6_u3_n110 ) , .B2( u0_u6_u3_n142 ) , .B1( u0_u6_u3_n186 ) , .A( u0_u6_u3_n95 ) );
  INV_X1 u0_u6_u3_U54 (.A( u0_u6_u3_n145 ) , .ZN( u0_u6_u3_n186 ) );
  AOI21_X1 u0_u6_u3_U55 (.B1( u0_u6_u3_n124 ) , .A( u0_u6_u3_n149 ) , .B2( u0_u6_u3_n155 ) , .ZN( u0_u6_u3_n95 ) );
  INV_X1 u0_u6_u3_U56 (.A( u0_u6_u3_n149 ) , .ZN( u0_u6_u3_n169 ) );
  NAND2_X1 u0_u6_u3_U57 (.ZN( u0_u6_u3_n124 ) , .A1( u0_u6_u3_n96 ) , .A2( u0_u6_u3_n97 ) );
  NAND2_X1 u0_u6_u3_U58 (.A2( u0_u6_u3_n100 ) , .ZN( u0_u6_u3_n146 ) , .A1( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U59 (.A1( u0_u6_u3_n101 ) , .ZN( u0_u6_u3_n145 ) , .A2( u0_u6_u3_n99 ) );
  AOI221_X1 u0_u6_u3_U6 (.A( u0_u6_u3_n131 ) , .C2( u0_u6_u3_n132 ) , .C1( u0_u6_u3_n133 ) , .ZN( u0_u6_u3_n134 ) , .B1( u0_u6_u3_n143 ) , .B2( u0_u6_u3_n177 ) );
  NAND2_X1 u0_u6_u3_U60 (.A1( u0_u6_u3_n100 ) , .ZN( u0_u6_u3_n156 ) , .A2( u0_u6_u3_n99 ) );
  NAND2_X1 u0_u6_u3_U61 (.A2( u0_u6_u3_n101 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n148 ) );
  NAND2_X1 u0_u6_u3_U62 (.A1( u0_u6_u3_n100 ) , .A2( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n128 ) );
  NAND2_X1 u0_u6_u3_U63 (.A2( u0_u6_u3_n101 ) , .A1( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n152 ) );
  NAND2_X1 u0_u6_u3_U64 (.A2( u0_u6_u3_n101 ) , .ZN( u0_u6_u3_n114 ) , .A1( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U65 (.ZN( u0_u6_u3_n107 ) , .A1( u0_u6_u3_n97 ) , .A2( u0_u6_u3_n99 ) );
  NAND2_X1 u0_u6_u3_U66 (.A2( u0_u6_u3_n100 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n113 ) );
  NAND2_X1 u0_u6_u3_U67 (.A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n153 ) , .A2( u0_u6_u3_n97 ) );
  NAND2_X1 u0_u6_u3_U68 (.A2( u0_u6_u3_n103 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n130 ) );
  NAND2_X1 u0_u6_u3_U69 (.A2( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n144 ) , .A1( u0_u6_u3_n96 ) );
  OAI22_X1 u0_u6_u3_U7 (.B2( u0_u6_u3_n147 ) , .A2( u0_u6_u3_n148 ) , .ZN( u0_u6_u3_n160 ) , .B1( u0_u6_u3_n165 ) , .A1( u0_u6_u3_n168 ) );
  NAND2_X1 u0_u6_u3_U70 (.A1( u0_u6_u3_n102 ) , .A2( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n108 ) );
  NOR2_X1 u0_u6_u3_U71 (.A2( u0_u6_X_19 ) , .A1( u0_u6_X_20 ) , .ZN( u0_u6_u3_n99 ) );
  NOR2_X1 u0_u6_u3_U72 (.A2( u0_u6_X_21 ) , .A1( u0_u6_X_24 ) , .ZN( u0_u6_u3_n103 ) );
  NOR2_X1 u0_u6_u3_U73 (.A2( u0_u6_X_24 ) , .A1( u0_u6_u3_n171 ) , .ZN( u0_u6_u3_n97 ) );
  NOR2_X1 u0_u6_u3_U74 (.A2( u0_u6_X_23 ) , .ZN( u0_u6_u3_n141 ) , .A1( u0_u6_u3_n166 ) );
  NOR2_X1 u0_u6_u3_U75 (.A2( u0_u6_X_19 ) , .A1( u0_u6_u3_n172 ) , .ZN( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U76 (.A1( u0_u6_X_22 ) , .A2( u0_u6_X_23 ) , .ZN( u0_u6_u3_n154 ) );
  NAND2_X1 u0_u6_u3_U77 (.A1( u0_u6_X_23 ) , .ZN( u0_u6_u3_n149 ) , .A2( u0_u6_u3_n166 ) );
  NOR2_X1 u0_u6_u3_U78 (.A2( u0_u6_X_22 ) , .A1( u0_u6_X_23 ) , .ZN( u0_u6_u3_n121 ) );
  AND2_X1 u0_u6_u3_U79 (.A1( u0_u6_X_24 ) , .ZN( u0_u6_u3_n101 ) , .A2( u0_u6_u3_n171 ) );
  AND3_X1 u0_u6_u3_U8 (.A3( u0_u6_u3_n144 ) , .A2( u0_u6_u3_n145 ) , .A1( u0_u6_u3_n146 ) , .ZN( u0_u6_u3_n147 ) );
  AND2_X1 u0_u6_u3_U80 (.A1( u0_u6_X_19 ) , .ZN( u0_u6_u3_n102 ) , .A2( u0_u6_u3_n172 ) );
  AND2_X1 u0_u6_u3_U81 (.A1( u0_u6_X_21 ) , .A2( u0_u6_X_24 ) , .ZN( u0_u6_u3_n100 ) );
  AND2_X1 u0_u6_u3_U82 (.A2( u0_u6_X_19 ) , .A1( u0_u6_X_20 ) , .ZN( u0_u6_u3_n104 ) );
  INV_X1 u0_u6_u3_U83 (.A( u0_u6_X_22 ) , .ZN( u0_u6_u3_n166 ) );
  INV_X1 u0_u6_u3_U84 (.A( u0_u6_X_21 ) , .ZN( u0_u6_u3_n171 ) );
  INV_X1 u0_u6_u3_U85 (.A( u0_u6_X_20 ) , .ZN( u0_u6_u3_n172 ) );
  NAND4_X1 u0_u6_u3_U86 (.ZN( u0_out6_26 ) , .A4( u0_u6_u3_n109 ) , .A3( u0_u6_u3_n110 ) , .A2( u0_u6_u3_n111 ) , .A1( u0_u6_u3_n173 ) );
  INV_X1 u0_u6_u3_U87 (.ZN( u0_u6_u3_n173 ) , .A( u0_u6_u3_n94 ) );
  OAI21_X1 u0_u6_u3_U88 (.ZN( u0_u6_u3_n111 ) , .B2( u0_u6_u3_n117 ) , .A( u0_u6_u3_n133 ) , .B1( u0_u6_u3_n176 ) );
  NAND4_X1 u0_u6_u3_U89 (.ZN( u0_out6_20 ) , .A4( u0_u6_u3_n122 ) , .A3( u0_u6_u3_n123 ) , .A1( u0_u6_u3_n175 ) , .A2( u0_u6_u3_n180 ) );
  INV_X1 u0_u6_u3_U9 (.A( u0_u6_u3_n143 ) , .ZN( u0_u6_u3_n168 ) );
  INV_X1 u0_u6_u3_U90 (.A( u0_u6_u3_n126 ) , .ZN( u0_u6_u3_n180 ) );
  INV_X1 u0_u6_u3_U91 (.A( u0_u6_u3_n112 ) , .ZN( u0_u6_u3_n175 ) );
  NAND4_X1 u0_u6_u3_U92 (.ZN( u0_out6_1 ) , .A4( u0_u6_u3_n161 ) , .A3( u0_u6_u3_n162 ) , .A2( u0_u6_u3_n163 ) , .A1( u0_u6_u3_n185 ) );
  NAND2_X1 u0_u6_u3_U93 (.ZN( u0_u6_u3_n163 ) , .A2( u0_u6_u3_n170 ) , .A1( u0_u6_u3_n176 ) );
  AOI22_X1 u0_u6_u3_U94 (.B2( u0_u6_u3_n140 ) , .B1( u0_u6_u3_n141 ) , .A2( u0_u6_u3_n142 ) , .ZN( u0_u6_u3_n162 ) , .A1( u0_u6_u3_n177 ) );
  OR4_X1 u0_u6_u3_U95 (.ZN( u0_out6_10 ) , .A4( u0_u6_u3_n136 ) , .A3( u0_u6_u3_n137 ) , .A1( u0_u6_u3_n138 ) , .A2( u0_u6_u3_n139 ) );
  OAI222_X1 u0_u6_u3_U96 (.C1( u0_u6_u3_n128 ) , .ZN( u0_u6_u3_n137 ) , .B1( u0_u6_u3_n148 ) , .A2( u0_u6_u3_n150 ) , .B2( u0_u6_u3_n154 ) , .C2( u0_u6_u3_n164 ) , .A1( u0_u6_u3_n167 ) );
  OAI221_X1 u0_u6_u3_U97 (.A( u0_u6_u3_n134 ) , .B2( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n136 ) , .C1( u0_u6_u3_n149 ) , .B1( u0_u6_u3_n151 ) , .C2( u0_u6_u3_n183 ) );
  NAND3_X1 u0_u6_u3_U98 (.A1( u0_u6_u3_n114 ) , .ZN( u0_u6_u3_n115 ) , .A2( u0_u6_u3_n145 ) , .A3( u0_u6_u3_n153 ) );
  NAND3_X1 u0_u6_u3_U99 (.ZN( u0_u6_u3_n129 ) , .A2( u0_u6_u3_n144 ) , .A1( u0_u6_u3_n153 ) , .A3( u0_u6_u3_n182 ) );
  AND3_X1 u0_u6_u7_U10 (.A3( u0_u6_u7_n110 ) , .A2( u0_u6_u7_n127 ) , .A1( u0_u6_u7_n132 ) , .ZN( u0_u6_u7_n92 ) );
  OAI21_X1 u0_u6_u7_U11 (.A( u0_u6_u7_n161 ) , .B1( u0_u6_u7_n168 ) , .B2( u0_u6_u7_n173 ) , .ZN( u0_u6_u7_n91 ) );
  AOI211_X1 u0_u6_u7_U12 (.A( u0_u6_u7_n117 ) , .ZN( u0_u6_u7_n118 ) , .C2( u0_u6_u7_n126 ) , .C1( u0_u6_u7_n177 ) , .B( u0_u6_u7_n180 ) );
  OAI22_X1 u0_u6_u7_U13 (.B1( u0_u6_u7_n115 ) , .ZN( u0_u6_u7_n117 ) , .A2( u0_u6_u7_n133 ) , .A1( u0_u6_u7_n137 ) , .B2( u0_u6_u7_n162 ) );
  INV_X1 u0_u6_u7_U14 (.A( u0_u6_u7_n116 ) , .ZN( u0_u6_u7_n180 ) );
  NOR3_X1 u0_u6_u7_U15 (.ZN( u0_u6_u7_n115 ) , .A3( u0_u6_u7_n145 ) , .A2( u0_u6_u7_n168 ) , .A1( u0_u6_u7_n169 ) );
  OAI211_X1 u0_u6_u7_U16 (.B( u0_u6_u7_n122 ) , .A( u0_u6_u7_n123 ) , .C2( u0_u6_u7_n124 ) , .ZN( u0_u6_u7_n154 ) , .C1( u0_u6_u7_n162 ) );
  AOI222_X1 u0_u6_u7_U17 (.ZN( u0_u6_u7_n122 ) , .C2( u0_u6_u7_n126 ) , .C1( u0_u6_u7_n145 ) , .B1( u0_u6_u7_n161 ) , .A2( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n170 ) , .A1( u0_u6_u7_n176 ) );
  INV_X1 u0_u6_u7_U18 (.A( u0_u6_u7_n133 ) , .ZN( u0_u6_u7_n176 ) );
  NOR3_X1 u0_u6_u7_U19 (.A2( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n135 ) , .ZN( u0_u6_u7_n136 ) , .A3( u0_u6_u7_n171 ) );
  NOR2_X1 u0_u6_u7_U20 (.A1( u0_u6_u7_n130 ) , .A2( u0_u6_u7_n134 ) , .ZN( u0_u6_u7_n153 ) );
  INV_X1 u0_u6_u7_U21 (.A( u0_u6_u7_n101 ) , .ZN( u0_u6_u7_n165 ) );
  NOR2_X1 u0_u6_u7_U22 (.ZN( u0_u6_u7_n111 ) , .A2( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n169 ) );
  AOI21_X1 u0_u6_u7_U23 (.ZN( u0_u6_u7_n104 ) , .B2( u0_u6_u7_n112 ) , .B1( u0_u6_u7_n127 ) , .A( u0_u6_u7_n164 ) );
  AOI21_X1 u0_u6_u7_U24 (.ZN( u0_u6_u7_n106 ) , .B1( u0_u6_u7_n133 ) , .B2( u0_u6_u7_n146 ) , .A( u0_u6_u7_n162 ) );
  AOI21_X1 u0_u6_u7_U25 (.A( u0_u6_u7_n101 ) , .ZN( u0_u6_u7_n107 ) , .B2( u0_u6_u7_n128 ) , .B1( u0_u6_u7_n175 ) );
  INV_X1 u0_u6_u7_U26 (.A( u0_u6_u7_n138 ) , .ZN( u0_u6_u7_n171 ) );
  INV_X1 u0_u6_u7_U27 (.A( u0_u6_u7_n131 ) , .ZN( u0_u6_u7_n177 ) );
  INV_X1 u0_u6_u7_U28 (.A( u0_u6_u7_n110 ) , .ZN( u0_u6_u7_n174 ) );
  NAND2_X1 u0_u6_u7_U29 (.A1( u0_u6_u7_n129 ) , .A2( u0_u6_u7_n132 ) , .ZN( u0_u6_u7_n149 ) );
  OAI21_X1 u0_u6_u7_U3 (.ZN( u0_u6_u7_n159 ) , .A( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n171 ) , .B1( u0_u6_u7_n174 ) );
  NAND2_X1 u0_u6_u7_U30 (.A1( u0_u6_u7_n113 ) , .A2( u0_u6_u7_n124 ) , .ZN( u0_u6_u7_n130 ) );
  INV_X1 u0_u6_u7_U31 (.A( u0_u6_u7_n112 ) , .ZN( u0_u6_u7_n173 ) );
  INV_X1 u0_u6_u7_U32 (.A( u0_u6_u7_n128 ) , .ZN( u0_u6_u7_n168 ) );
  INV_X1 u0_u6_u7_U33 (.A( u0_u6_u7_n148 ) , .ZN( u0_u6_u7_n169 ) );
  INV_X1 u0_u6_u7_U34 (.A( u0_u6_u7_n127 ) , .ZN( u0_u6_u7_n179 ) );
  NOR2_X1 u0_u6_u7_U35 (.ZN( u0_u6_u7_n101 ) , .A2( u0_u6_u7_n150 ) , .A1( u0_u6_u7_n156 ) );
  AOI211_X1 u0_u6_u7_U36 (.B( u0_u6_u7_n154 ) , .A( u0_u6_u7_n155 ) , .C1( u0_u6_u7_n156 ) , .ZN( u0_u6_u7_n157 ) , .C2( u0_u6_u7_n172 ) );
  INV_X1 u0_u6_u7_U37 (.A( u0_u6_u7_n153 ) , .ZN( u0_u6_u7_n172 ) );
  AOI211_X1 u0_u6_u7_U38 (.B( u0_u6_u7_n139 ) , .A( u0_u6_u7_n140 ) , .C2( u0_u6_u7_n141 ) , .ZN( u0_u6_u7_n142 ) , .C1( u0_u6_u7_n156 ) );
  NAND4_X1 u0_u6_u7_U39 (.A3( u0_u6_u7_n127 ) , .A2( u0_u6_u7_n128 ) , .A1( u0_u6_u7_n129 ) , .ZN( u0_u6_u7_n141 ) , .A4( u0_u6_u7_n147 ) );
  INV_X1 u0_u6_u7_U4 (.A( u0_u6_u7_n111 ) , .ZN( u0_u6_u7_n170 ) );
  AOI21_X1 u0_u6_u7_U40 (.A( u0_u6_u7_n137 ) , .B1( u0_u6_u7_n138 ) , .ZN( u0_u6_u7_n139 ) , .B2( u0_u6_u7_n146 ) );
  OAI22_X1 u0_u6_u7_U41 (.B1( u0_u6_u7_n136 ) , .ZN( u0_u6_u7_n140 ) , .A1( u0_u6_u7_n153 ) , .B2( u0_u6_u7_n162 ) , .A2( u0_u6_u7_n164 ) );
  AOI21_X1 u0_u6_u7_U42 (.ZN( u0_u6_u7_n123 ) , .B1( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n177 ) , .A( u0_u6_u7_n97 ) );
  AOI21_X1 u0_u6_u7_U43 (.B2( u0_u6_u7_n113 ) , .B1( u0_u6_u7_n124 ) , .A( u0_u6_u7_n125 ) , .ZN( u0_u6_u7_n97 ) );
  INV_X1 u0_u6_u7_U44 (.A( u0_u6_u7_n125 ) , .ZN( u0_u6_u7_n161 ) );
  INV_X1 u0_u6_u7_U45 (.A( u0_u6_u7_n152 ) , .ZN( u0_u6_u7_n162 ) );
  AOI22_X1 u0_u6_u7_U46 (.A2( u0_u6_u7_n114 ) , .ZN( u0_u6_u7_n119 ) , .B1( u0_u6_u7_n130 ) , .A1( u0_u6_u7_n156 ) , .B2( u0_u6_u7_n165 ) );
  NAND2_X1 u0_u6_u7_U47 (.A2( u0_u6_u7_n112 ) , .ZN( u0_u6_u7_n114 ) , .A1( u0_u6_u7_n175 ) );
  AND2_X1 u0_u6_u7_U48 (.ZN( u0_u6_u7_n145 ) , .A2( u0_u6_u7_n98 ) , .A1( u0_u6_u7_n99 ) );
  NOR2_X1 u0_u6_u7_U49 (.ZN( u0_u6_u7_n137 ) , .A1( u0_u6_u7_n150 ) , .A2( u0_u6_u7_n161 ) );
  INV_X1 u0_u6_u7_U5 (.A( u0_u6_u7_n149 ) , .ZN( u0_u6_u7_n175 ) );
  AOI21_X1 u0_u6_u7_U50 (.ZN( u0_u6_u7_n105 ) , .B2( u0_u6_u7_n110 ) , .A( u0_u6_u7_n125 ) , .B1( u0_u6_u7_n147 ) );
  NAND2_X1 u0_u6_u7_U51 (.ZN( u0_u6_u7_n146 ) , .A1( u0_u6_u7_n95 ) , .A2( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U52 (.A2( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n147 ) , .A1( u0_u6_u7_n93 ) );
  NAND2_X1 u0_u6_u7_U53 (.A1( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n127 ) , .A2( u0_u6_u7_n99 ) );
  OR2_X1 u0_u6_u7_U54 (.ZN( u0_u6_u7_n126 ) , .A2( u0_u6_u7_n152 ) , .A1( u0_u6_u7_n156 ) );
  NAND2_X1 u0_u6_u7_U55 (.A2( u0_u6_u7_n102 ) , .A1( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n133 ) );
  NAND2_X1 u0_u6_u7_U56 (.ZN( u0_u6_u7_n112 ) , .A2( u0_u6_u7_n96 ) , .A1( u0_u6_u7_n99 ) );
  NAND2_X1 u0_u6_u7_U57 (.A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n128 ) , .A1( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U58 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n113 ) , .A2( u0_u6_u7_n93 ) );
  NAND2_X1 u0_u6_u7_U59 (.A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n124 ) , .A1( u0_u6_u7_n96 ) );
  INV_X1 u0_u6_u7_U6 (.A( u0_u6_u7_n154 ) , .ZN( u0_u6_u7_n178 ) );
  NAND2_X1 u0_u6_u7_U60 (.ZN( u0_u6_u7_n110 ) , .A1( u0_u6_u7_n95 ) , .A2( u0_u6_u7_n96 ) );
  INV_X1 u0_u6_u7_U61 (.A( u0_u6_u7_n150 ) , .ZN( u0_u6_u7_n164 ) );
  AND2_X1 u0_u6_u7_U62 (.ZN( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n93 ) , .A2( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U63 (.A1( u0_u6_u7_n100 ) , .A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n129 ) );
  NAND2_X1 u0_u6_u7_U64 (.A2( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n131 ) , .A1( u0_u6_u7_n95 ) );
  NAND2_X1 u0_u6_u7_U65 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n138 ) , .A2( u0_u6_u7_n99 ) );
  NAND2_X1 u0_u6_u7_U66 (.ZN( u0_u6_u7_n132 ) , .A1( u0_u6_u7_n93 ) , .A2( u0_u6_u7_n96 ) );
  NAND2_X1 u0_u6_u7_U67 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n148 ) , .A2( u0_u6_u7_n95 ) );
  NOR2_X1 u0_u6_u7_U68 (.A2( u0_u6_X_47 ) , .ZN( u0_u6_u7_n150 ) , .A1( u0_u6_u7_n163 ) );
  NOR2_X1 u0_u6_u7_U69 (.A2( u0_u6_X_43 ) , .A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n103 ) );
  AOI211_X1 u0_u6_u7_U7 (.ZN( u0_u6_u7_n116 ) , .A( u0_u6_u7_n155 ) , .C1( u0_u6_u7_n161 ) , .C2( u0_u6_u7_n171 ) , .B( u0_u6_u7_n94 ) );
  NOR2_X1 u0_u6_u7_U70 (.A2( u0_u6_X_48 ) , .A1( u0_u6_u7_n166 ) , .ZN( u0_u6_u7_n95 ) );
  NOR2_X1 u0_u6_u7_U71 (.A2( u0_u6_X_45 ) , .A1( u0_u6_X_48 ) , .ZN( u0_u6_u7_n99 ) );
  NOR2_X1 u0_u6_u7_U72 (.A2( u0_u6_X_44 ) , .A1( u0_u6_u7_n167 ) , .ZN( u0_u6_u7_n98 ) );
  NOR2_X1 u0_u6_u7_U73 (.A2( u0_u6_X_46 ) , .A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n152 ) );
  AND2_X1 u0_u6_u7_U74 (.A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n156 ) , .A2( u0_u6_u7_n163 ) );
  NAND2_X1 u0_u6_u7_U75 (.A2( u0_u6_X_46 ) , .A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n125 ) );
  AND2_X1 u0_u6_u7_U76 (.A2( u0_u6_X_45 ) , .A1( u0_u6_X_48 ) , .ZN( u0_u6_u7_n102 ) );
  AND2_X1 u0_u6_u7_U77 (.A2( u0_u6_X_43 ) , .A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n96 ) );
  AND2_X1 u0_u6_u7_U78 (.A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n100 ) , .A2( u0_u6_u7_n167 ) );
  AND2_X1 u0_u6_u7_U79 (.A1( u0_u6_X_48 ) , .A2( u0_u6_u7_n166 ) , .ZN( u0_u6_u7_n93 ) );
  OAI222_X1 u0_u6_u7_U8 (.C2( u0_u6_u7_n101 ) , .B2( u0_u6_u7_n111 ) , .A1( u0_u6_u7_n113 ) , .C1( u0_u6_u7_n146 ) , .A2( u0_u6_u7_n162 ) , .B1( u0_u6_u7_n164 ) , .ZN( u0_u6_u7_n94 ) );
  INV_X1 u0_u6_u7_U80 (.A( u0_u6_X_46 ) , .ZN( u0_u6_u7_n163 ) );
  INV_X1 u0_u6_u7_U81 (.A( u0_u6_X_43 ) , .ZN( u0_u6_u7_n167 ) );
  INV_X1 u0_u6_u7_U82 (.A( u0_u6_X_45 ) , .ZN( u0_u6_u7_n166 ) );
  NAND4_X1 u0_u6_u7_U83 (.ZN( u0_out6_5 ) , .A4( u0_u6_u7_n108 ) , .A3( u0_u6_u7_n109 ) , .A1( u0_u6_u7_n116 ) , .A2( u0_u6_u7_n123 ) );
  AOI22_X1 u0_u6_u7_U84 (.ZN( u0_u6_u7_n109 ) , .A2( u0_u6_u7_n126 ) , .B2( u0_u6_u7_n145 ) , .B1( u0_u6_u7_n156 ) , .A1( u0_u6_u7_n171 ) );
  NOR4_X1 u0_u6_u7_U85 (.A4( u0_u6_u7_n104 ) , .A3( u0_u6_u7_n105 ) , .A2( u0_u6_u7_n106 ) , .A1( u0_u6_u7_n107 ) , .ZN( u0_u6_u7_n108 ) );
  NAND4_X1 u0_u6_u7_U86 (.ZN( u0_out6_27 ) , .A4( u0_u6_u7_n118 ) , .A3( u0_u6_u7_n119 ) , .A2( u0_u6_u7_n120 ) , .A1( u0_u6_u7_n121 ) );
  OAI21_X1 u0_u6_u7_U87 (.ZN( u0_u6_u7_n121 ) , .B2( u0_u6_u7_n145 ) , .A( u0_u6_u7_n150 ) , .B1( u0_u6_u7_n174 ) );
  OAI21_X1 u0_u6_u7_U88 (.ZN( u0_u6_u7_n120 ) , .A( u0_u6_u7_n161 ) , .B2( u0_u6_u7_n170 ) , .B1( u0_u6_u7_n179 ) );
  NAND4_X1 u0_u6_u7_U89 (.ZN( u0_out6_21 ) , .A4( u0_u6_u7_n157 ) , .A3( u0_u6_u7_n158 ) , .A2( u0_u6_u7_n159 ) , .A1( u0_u6_u7_n160 ) );
  OAI221_X1 u0_u6_u7_U9 (.C1( u0_u6_u7_n101 ) , .C2( u0_u6_u7_n147 ) , .ZN( u0_u6_u7_n155 ) , .B2( u0_u6_u7_n162 ) , .A( u0_u6_u7_n91 ) , .B1( u0_u6_u7_n92 ) );
  OAI21_X1 u0_u6_u7_U90 (.B1( u0_u6_u7_n145 ) , .ZN( u0_u6_u7_n160 ) , .A( u0_u6_u7_n161 ) , .B2( u0_u6_u7_n177 ) );
  AOI22_X1 u0_u6_u7_U91 (.B2( u0_u6_u7_n149 ) , .B1( u0_u6_u7_n150 ) , .A2( u0_u6_u7_n151 ) , .A1( u0_u6_u7_n152 ) , .ZN( u0_u6_u7_n158 ) );
  NAND4_X1 u0_u6_u7_U92 (.ZN( u0_out6_15 ) , .A4( u0_u6_u7_n142 ) , .A3( u0_u6_u7_n143 ) , .A2( u0_u6_u7_n144 ) , .A1( u0_u6_u7_n178 ) );
  OR2_X1 u0_u6_u7_U93 (.A2( u0_u6_u7_n125 ) , .A1( u0_u6_u7_n129 ) , .ZN( u0_u6_u7_n144 ) );
  AOI22_X1 u0_u6_u7_U94 (.A2( u0_u6_u7_n126 ) , .ZN( u0_u6_u7_n143 ) , .B2( u0_u6_u7_n165 ) , .B1( u0_u6_u7_n173 ) , .A1( u0_u6_u7_n174 ) );
  NAND3_X1 u0_u6_u7_U95 (.A3( u0_u6_u7_n146 ) , .A2( u0_u6_u7_n147 ) , .A1( u0_u6_u7_n148 ) , .ZN( u0_u6_u7_n151 ) );
  NAND3_X1 u0_u6_u7_U96 (.A3( u0_u6_u7_n131 ) , .A2( u0_u6_u7_n132 ) , .A1( u0_u6_u7_n133 ) , .ZN( u0_u6_u7_n135 ) );
  XOR2_X1 u0_u7_U10 (.B( u0_K8_45 ) , .A( u0_R6_30 ) , .Z( u0_u7_X_45 ) );
  XOR2_X1 u0_u7_U11 (.B( u0_K8_44 ) , .A( u0_R6_29 ) , .Z( u0_u7_X_44 ) );
  XOR2_X1 u0_u7_U12 (.B( u0_K8_43 ) , .A( u0_R6_28 ) , .Z( u0_u7_X_43 ) );
  XOR2_X1 u0_u7_U7 (.B( u0_K8_48 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_48 ) );
  XOR2_X1 u0_u7_U8 (.B( u0_K8_47 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_47 ) );
  XOR2_X1 u0_u7_U9 (.B( u0_K8_46 ) , .A( u0_R6_31 ) , .Z( u0_u7_X_46 ) );
  OAI221_X1 u0_u7_u7_U10 (.C1( u0_u7_u7_n101 ) , .C2( u0_u7_u7_n147 ) , .ZN( u0_u7_u7_n155 ) , .B2( u0_u7_u7_n162 ) , .A( u0_u7_u7_n91 ) , .B1( u0_u7_u7_n92 ) );
  AND3_X1 u0_u7_u7_U11 (.A3( u0_u7_u7_n110 ) , .A2( u0_u7_u7_n127 ) , .A1( u0_u7_u7_n132 ) , .ZN( u0_u7_u7_n92 ) );
  OAI21_X1 u0_u7_u7_U12 (.A( u0_u7_u7_n161 ) , .B1( u0_u7_u7_n168 ) , .B2( u0_u7_u7_n173 ) , .ZN( u0_u7_u7_n91 ) );
  AOI211_X1 u0_u7_u7_U13 (.A( u0_u7_u7_n117 ) , .ZN( u0_u7_u7_n118 ) , .C2( u0_u7_u7_n126 ) , .C1( u0_u7_u7_n177 ) , .B( u0_u7_u7_n180 ) );
  OAI22_X1 u0_u7_u7_U14 (.B1( u0_u7_u7_n115 ) , .ZN( u0_u7_u7_n117 ) , .A2( u0_u7_u7_n133 ) , .A1( u0_u7_u7_n137 ) , .B2( u0_u7_u7_n162 ) );
  INV_X1 u0_u7_u7_U15 (.A( u0_u7_u7_n116 ) , .ZN( u0_u7_u7_n180 ) );
  NOR3_X1 u0_u7_u7_U16 (.ZN( u0_u7_u7_n115 ) , .A3( u0_u7_u7_n145 ) , .A2( u0_u7_u7_n168 ) , .A1( u0_u7_u7_n169 ) );
  NOR3_X1 u0_u7_u7_U17 (.A2( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n135 ) , .ZN( u0_u7_u7_n136 ) , .A3( u0_u7_u7_n171 ) );
  NOR2_X1 u0_u7_u7_U18 (.A1( u0_u7_u7_n130 ) , .A2( u0_u7_u7_n134 ) , .ZN( u0_u7_u7_n153 ) );
  NOR2_X1 u0_u7_u7_U19 (.ZN( u0_u7_u7_n111 ) , .A2( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n169 ) );
  AOI21_X1 u0_u7_u7_U20 (.ZN( u0_u7_u7_n104 ) , .B2( u0_u7_u7_n112 ) , .B1( u0_u7_u7_n127 ) , .A( u0_u7_u7_n164 ) );
  AOI21_X1 u0_u7_u7_U21 (.ZN( u0_u7_u7_n106 ) , .B1( u0_u7_u7_n133 ) , .B2( u0_u7_u7_n146 ) , .A( u0_u7_u7_n162 ) );
  AOI21_X1 u0_u7_u7_U22 (.A( u0_u7_u7_n101 ) , .ZN( u0_u7_u7_n107 ) , .B2( u0_u7_u7_n128 ) , .B1( u0_u7_u7_n175 ) );
  INV_X1 u0_u7_u7_U23 (.A( u0_u7_u7_n101 ) , .ZN( u0_u7_u7_n165 ) );
  INV_X1 u0_u7_u7_U24 (.A( u0_u7_u7_n138 ) , .ZN( u0_u7_u7_n171 ) );
  INV_X1 u0_u7_u7_U25 (.A( u0_u7_u7_n131 ) , .ZN( u0_u7_u7_n177 ) );
  INV_X1 u0_u7_u7_U26 (.A( u0_u7_u7_n110 ) , .ZN( u0_u7_u7_n174 ) );
  NAND2_X1 u0_u7_u7_U27 (.A1( u0_u7_u7_n129 ) , .A2( u0_u7_u7_n132 ) , .ZN( u0_u7_u7_n149 ) );
  NAND2_X1 u0_u7_u7_U28 (.A1( u0_u7_u7_n113 ) , .A2( u0_u7_u7_n124 ) , .ZN( u0_u7_u7_n130 ) );
  INV_X1 u0_u7_u7_U29 (.A( u0_u7_u7_n128 ) , .ZN( u0_u7_u7_n168 ) );
  OAI21_X1 u0_u7_u7_U3 (.ZN( u0_u7_u7_n159 ) , .A( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n171 ) , .B1( u0_u7_u7_n174 ) );
  INV_X1 u0_u7_u7_U30 (.A( u0_u7_u7_n148 ) , .ZN( u0_u7_u7_n169 ) );
  INV_X1 u0_u7_u7_U31 (.A( u0_u7_u7_n112 ) , .ZN( u0_u7_u7_n173 ) );
  INV_X1 u0_u7_u7_U32 (.A( u0_u7_u7_n127 ) , .ZN( u0_u7_u7_n179 ) );
  NOR2_X1 u0_u7_u7_U33 (.ZN( u0_u7_u7_n101 ) , .A2( u0_u7_u7_n150 ) , .A1( u0_u7_u7_n156 ) );
  AOI211_X1 u0_u7_u7_U34 (.B( u0_u7_u7_n154 ) , .A( u0_u7_u7_n155 ) , .C1( u0_u7_u7_n156 ) , .ZN( u0_u7_u7_n157 ) , .C2( u0_u7_u7_n172 ) );
  INV_X1 u0_u7_u7_U35 (.A( u0_u7_u7_n153 ) , .ZN( u0_u7_u7_n172 ) );
  AOI211_X1 u0_u7_u7_U36 (.B( u0_u7_u7_n139 ) , .A( u0_u7_u7_n140 ) , .C2( u0_u7_u7_n141 ) , .ZN( u0_u7_u7_n142 ) , .C1( u0_u7_u7_n156 ) );
  NAND4_X1 u0_u7_u7_U37 (.A3( u0_u7_u7_n127 ) , .A2( u0_u7_u7_n128 ) , .A1( u0_u7_u7_n129 ) , .ZN( u0_u7_u7_n141 ) , .A4( u0_u7_u7_n147 ) );
  AOI21_X1 u0_u7_u7_U38 (.A( u0_u7_u7_n137 ) , .B1( u0_u7_u7_n138 ) , .ZN( u0_u7_u7_n139 ) , .B2( u0_u7_u7_n146 ) );
  OAI22_X1 u0_u7_u7_U39 (.B1( u0_u7_u7_n136 ) , .ZN( u0_u7_u7_n140 ) , .A1( u0_u7_u7_n153 ) , .B2( u0_u7_u7_n162 ) , .A2( u0_u7_u7_n164 ) );
  INV_X1 u0_u7_u7_U4 (.A( u0_u7_u7_n149 ) , .ZN( u0_u7_u7_n175 ) );
  INV_X1 u0_u7_u7_U40 (.A( u0_u7_u7_n125 ) , .ZN( u0_u7_u7_n161 ) );
  AOI21_X1 u0_u7_u7_U41 (.ZN( u0_u7_u7_n123 ) , .B1( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n177 ) , .A( u0_u7_u7_n97 ) );
  AOI21_X1 u0_u7_u7_U42 (.B2( u0_u7_u7_n113 ) , .B1( u0_u7_u7_n124 ) , .A( u0_u7_u7_n125 ) , .ZN( u0_u7_u7_n97 ) );
  INV_X1 u0_u7_u7_U43 (.A( u0_u7_u7_n152 ) , .ZN( u0_u7_u7_n162 ) );
  AOI22_X1 u0_u7_u7_U44 (.A2( u0_u7_u7_n114 ) , .ZN( u0_u7_u7_n119 ) , .B1( u0_u7_u7_n130 ) , .A1( u0_u7_u7_n156 ) , .B2( u0_u7_u7_n165 ) );
  NAND2_X1 u0_u7_u7_U45 (.A2( u0_u7_u7_n112 ) , .ZN( u0_u7_u7_n114 ) , .A1( u0_u7_u7_n175 ) );
  NOR2_X1 u0_u7_u7_U46 (.ZN( u0_u7_u7_n137 ) , .A1( u0_u7_u7_n150 ) , .A2( u0_u7_u7_n161 ) );
  AND2_X1 u0_u7_u7_U47 (.ZN( u0_u7_u7_n145 ) , .A2( u0_u7_u7_n98 ) , .A1( u0_u7_u7_n99 ) );
  AOI21_X1 u0_u7_u7_U48 (.ZN( u0_u7_u7_n105 ) , .B2( u0_u7_u7_n110 ) , .A( u0_u7_u7_n125 ) , .B1( u0_u7_u7_n147 ) );
  NAND2_X1 u0_u7_u7_U49 (.ZN( u0_u7_u7_n146 ) , .A1( u0_u7_u7_n95 ) , .A2( u0_u7_u7_n98 ) );
  INV_X1 u0_u7_u7_U5 (.A( u0_u7_u7_n154 ) , .ZN( u0_u7_u7_n178 ) );
  NAND2_X1 u0_u7_u7_U50 (.A2( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n147 ) , .A1( u0_u7_u7_n93 ) );
  NAND2_X1 u0_u7_u7_U51 (.A1( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n127 ) , .A2( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U52 (.A2( u0_u7_u7_n102 ) , .A1( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n133 ) );
  OR2_X1 u0_u7_u7_U53 (.ZN( u0_u7_u7_n126 ) , .A2( u0_u7_u7_n152 ) , .A1( u0_u7_u7_n156 ) );
  NAND2_X1 u0_u7_u7_U54 (.ZN( u0_u7_u7_n112 ) , .A2( u0_u7_u7_n96 ) , .A1( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U55 (.A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n128 ) , .A1( u0_u7_u7_n98 ) );
  INV_X1 u0_u7_u7_U56 (.A( u0_u7_u7_n150 ) , .ZN( u0_u7_u7_n164 ) );
  AND2_X1 u0_u7_u7_U57 (.ZN( u0_u7_u7_n134 ) , .A1( u0_u7_u7_n93 ) , .A2( u0_u7_u7_n98 ) );
  NAND2_X1 u0_u7_u7_U58 (.ZN( u0_u7_u7_n110 ) , .A1( u0_u7_u7_n95 ) , .A2( u0_u7_u7_n96 ) );
  NAND2_X1 u0_u7_u7_U59 (.A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n124 ) , .A1( u0_u7_u7_n96 ) );
  INV_X1 u0_u7_u7_U6 (.A( u0_u7_u7_n111 ) , .ZN( u0_u7_u7_n170 ) );
  NAND2_X1 u0_u7_u7_U60 (.ZN( u0_u7_u7_n132 ) , .A1( u0_u7_u7_n93 ) , .A2( u0_u7_u7_n96 ) );
  NAND2_X1 u0_u7_u7_U61 (.A2( u0_u7_u7_n103 ) , .ZN( u0_u7_u7_n131 ) , .A1( u0_u7_u7_n95 ) );
  NOR2_X1 u0_u7_u7_U62 (.A2( u0_u7_X_47 ) , .ZN( u0_u7_u7_n150 ) , .A1( u0_u7_u7_n163 ) );
  NOR2_X1 u0_u7_u7_U63 (.A2( u0_u7_X_43 ) , .A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n103 ) );
  NOR2_X1 u0_u7_u7_U64 (.A2( u0_u7_X_48 ) , .A1( u0_u7_u7_n166 ) , .ZN( u0_u7_u7_n95 ) );
  NOR2_X1 u0_u7_u7_U65 (.A2( u0_u7_X_44 ) , .A1( u0_u7_u7_n167 ) , .ZN( u0_u7_u7_n98 ) );
  NOR2_X1 u0_u7_u7_U66 (.A2( u0_u7_X_45 ) , .A1( u0_u7_X_48 ) , .ZN( u0_u7_u7_n99 ) );
  NOR2_X1 u0_u7_u7_U67 (.A2( u0_u7_X_46 ) , .A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n152 ) );
  AND2_X1 u0_u7_u7_U68 (.A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n156 ) , .A2( u0_u7_u7_n163 ) );
  NAND2_X1 u0_u7_u7_U69 (.A2( u0_u7_X_46 ) , .A1( u0_u7_X_47 ) , .ZN( u0_u7_u7_n125 ) );
  AOI211_X1 u0_u7_u7_U7 (.ZN( u0_u7_u7_n116 ) , .A( u0_u7_u7_n155 ) , .C1( u0_u7_u7_n161 ) , .C2( u0_u7_u7_n171 ) , .B( u0_u7_u7_n94 ) );
  AND2_X1 u0_u7_u7_U70 (.A2( u0_u7_X_43 ) , .A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n96 ) );
  AND2_X1 u0_u7_u7_U71 (.A2( u0_u7_X_45 ) , .A1( u0_u7_X_48 ) , .ZN( u0_u7_u7_n102 ) );
  AND2_X1 u0_u7_u7_U72 (.A1( u0_u7_X_48 ) , .A2( u0_u7_u7_n166 ) , .ZN( u0_u7_u7_n93 ) );
  INV_X1 u0_u7_u7_U73 (.A( u0_u7_X_46 ) , .ZN( u0_u7_u7_n163 ) );
  AND2_X1 u0_u7_u7_U74 (.A1( u0_u7_X_44 ) , .ZN( u0_u7_u7_n100 ) , .A2( u0_u7_u7_n167 ) );
  INV_X1 u0_u7_u7_U75 (.A( u0_u7_X_45 ) , .ZN( u0_u7_u7_n166 ) );
  INV_X1 u0_u7_u7_U76 (.A( u0_u7_X_43 ) , .ZN( u0_u7_u7_n167 ) );
  NAND4_X1 u0_u7_u7_U77 (.ZN( u0_out7_5 ) , .A4( u0_u7_u7_n108 ) , .A3( u0_u7_u7_n109 ) , .A1( u0_u7_u7_n116 ) , .A2( u0_u7_u7_n123 ) );
  AOI22_X1 u0_u7_u7_U78 (.ZN( u0_u7_u7_n109 ) , .A2( u0_u7_u7_n126 ) , .B2( u0_u7_u7_n145 ) , .B1( u0_u7_u7_n156 ) , .A1( u0_u7_u7_n171 ) );
  NOR4_X1 u0_u7_u7_U79 (.A4( u0_u7_u7_n104 ) , .A3( u0_u7_u7_n105 ) , .A2( u0_u7_u7_n106 ) , .A1( u0_u7_u7_n107 ) , .ZN( u0_u7_u7_n108 ) );
  OAI222_X1 u0_u7_u7_U8 (.C2( u0_u7_u7_n101 ) , .B2( u0_u7_u7_n111 ) , .A1( u0_u7_u7_n113 ) , .C1( u0_u7_u7_n146 ) , .A2( u0_u7_u7_n162 ) , .B1( u0_u7_u7_n164 ) , .ZN( u0_u7_u7_n94 ) );
  NAND4_X1 u0_u7_u7_U80 (.ZN( u0_out7_27 ) , .A4( u0_u7_u7_n118 ) , .A3( u0_u7_u7_n119 ) , .A2( u0_u7_u7_n120 ) , .A1( u0_u7_u7_n121 ) );
  OAI21_X1 u0_u7_u7_U81 (.ZN( u0_u7_u7_n121 ) , .B2( u0_u7_u7_n145 ) , .A( u0_u7_u7_n150 ) , .B1( u0_u7_u7_n174 ) );
  OAI21_X1 u0_u7_u7_U82 (.ZN( u0_u7_u7_n120 ) , .A( u0_u7_u7_n161 ) , .B2( u0_u7_u7_n170 ) , .B1( u0_u7_u7_n179 ) );
  NAND4_X1 u0_u7_u7_U83 (.ZN( u0_out7_21 ) , .A4( u0_u7_u7_n157 ) , .A3( u0_u7_u7_n158 ) , .A2( u0_u7_u7_n159 ) , .A1( u0_u7_u7_n160 ) );
  OAI21_X1 u0_u7_u7_U84 (.B1( u0_u7_u7_n145 ) , .ZN( u0_u7_u7_n160 ) , .A( u0_u7_u7_n161 ) , .B2( u0_u7_u7_n177 ) );
  AOI22_X1 u0_u7_u7_U85 (.B2( u0_u7_u7_n149 ) , .B1( u0_u7_u7_n150 ) , .A2( u0_u7_u7_n151 ) , .A1( u0_u7_u7_n152 ) , .ZN( u0_u7_u7_n158 ) );
  NAND4_X1 u0_u7_u7_U86 (.ZN( u0_out7_15 ) , .A4( u0_u7_u7_n142 ) , .A3( u0_u7_u7_n143 ) , .A2( u0_u7_u7_n144 ) , .A1( u0_u7_u7_n178 ) );
  OR2_X1 u0_u7_u7_U87 (.A2( u0_u7_u7_n125 ) , .A1( u0_u7_u7_n129 ) , .ZN( u0_u7_u7_n144 ) );
  AOI22_X1 u0_u7_u7_U88 (.A2( u0_u7_u7_n126 ) , .ZN( u0_u7_u7_n143 ) , .B2( u0_u7_u7_n165 ) , .B1( u0_u7_u7_n173 ) , .A1( u0_u7_u7_n174 ) );
  NAND2_X1 u0_u7_u7_U89 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n148 ) , .A2( u0_u7_u7_n95 ) );
  INV_X1 u0_u7_u7_U9 (.A( u0_u7_u7_n133 ) , .ZN( u0_u7_u7_n176 ) );
  NAND2_X1 u0_u7_u7_U90 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n113 ) , .A2( u0_u7_u7_n93 ) );
  NAND2_X1 u0_u7_u7_U91 (.A1( u0_u7_u7_n100 ) , .ZN( u0_u7_u7_n138 ) , .A2( u0_u7_u7_n99 ) );
  NAND2_X1 u0_u7_u7_U92 (.A1( u0_u7_u7_n100 ) , .A2( u0_u7_u7_n102 ) , .ZN( u0_u7_u7_n129 ) );
  OAI211_X1 u0_u7_u7_U93 (.B( u0_u7_u7_n122 ) , .A( u0_u7_u7_n123 ) , .C2( u0_u7_u7_n124 ) , .ZN( u0_u7_u7_n154 ) , .C1( u0_u7_u7_n162 ) );
  AOI222_X1 u0_u7_u7_U94 (.ZN( u0_u7_u7_n122 ) , .C2( u0_u7_u7_n126 ) , .C1( u0_u7_u7_n145 ) , .B1( u0_u7_u7_n161 ) , .A2( u0_u7_u7_n165 ) , .B2( u0_u7_u7_n170 ) , .A1( u0_u7_u7_n176 ) );
  NAND3_X1 u0_u7_u7_U95 (.A3( u0_u7_u7_n146 ) , .A2( u0_u7_u7_n147 ) , .A1( u0_u7_u7_n148 ) , .ZN( u0_u7_u7_n151 ) );
  NAND3_X1 u0_u7_u7_U96 (.A3( u0_u7_u7_n131 ) , .A2( u0_u7_u7_n132 ) , .A1( u0_u7_u7_n133 ) , .ZN( u0_u7_u7_n135 ) );
  XOR2_X1 u0_u9_U33 (.B( u0_K10_24 ) , .A( u0_R8_17 ) , .Z( u0_u9_X_24 ) );
  XOR2_X1 u0_u9_U34 (.B( u0_K10_23 ) , .A( u0_R8_16 ) , .Z( u0_u9_X_23 ) );
  XOR2_X1 u0_u9_U35 (.B( u0_K10_22 ) , .A( u0_R8_15 ) , .Z( u0_u9_X_22 ) );
  XOR2_X1 u0_u9_U36 (.B( u0_K10_21 ) , .A( u0_R8_14 ) , .Z( u0_u9_X_21 ) );
  XOR2_X1 u0_u9_U37 (.B( u0_K10_20 ) , .A( u0_R8_13 ) , .Z( u0_u9_X_20 ) );
  XOR2_X1 u0_u9_U39 (.B( u0_K10_19 ) , .A( u0_R8_12 ) , .Z( u0_u9_X_19 ) );
  OAI22_X1 u0_u9_u3_U10 (.B1( u0_u9_u3_n113 ) , .A2( u0_u9_u3_n135 ) , .A1( u0_u9_u3_n150 ) , .B2( u0_u9_u3_n164 ) , .ZN( u0_u9_u3_n98 ) );
  OAI211_X1 u0_u9_u3_U11 (.B( u0_u9_u3_n106 ) , .ZN( u0_u9_u3_n119 ) , .C2( u0_u9_u3_n128 ) , .C1( u0_u9_u3_n167 ) , .A( u0_u9_u3_n181 ) );
  AOI221_X1 u0_u9_u3_U12 (.C1( u0_u9_u3_n105 ) , .ZN( u0_u9_u3_n106 ) , .A( u0_u9_u3_n131 ) , .B2( u0_u9_u3_n132 ) , .C2( u0_u9_u3_n133 ) , .B1( u0_u9_u3_n169 ) );
  INV_X1 u0_u9_u3_U13 (.ZN( u0_u9_u3_n181 ) , .A( u0_u9_u3_n98 ) );
  NAND2_X1 u0_u9_u3_U14 (.ZN( u0_u9_u3_n105 ) , .A2( u0_u9_u3_n130 ) , .A1( u0_u9_u3_n155 ) );
  AOI22_X1 u0_u9_u3_U15 (.B1( u0_u9_u3_n115 ) , .A2( u0_u9_u3_n116 ) , .ZN( u0_u9_u3_n123 ) , .B2( u0_u9_u3_n133 ) , .A1( u0_u9_u3_n169 ) );
  NAND2_X1 u0_u9_u3_U16 (.ZN( u0_u9_u3_n116 ) , .A2( u0_u9_u3_n151 ) , .A1( u0_u9_u3_n182 ) );
  NOR2_X1 u0_u9_u3_U17 (.ZN( u0_u9_u3_n126 ) , .A2( u0_u9_u3_n150 ) , .A1( u0_u9_u3_n164 ) );
  AOI21_X1 u0_u9_u3_U18 (.ZN( u0_u9_u3_n112 ) , .B2( u0_u9_u3_n146 ) , .B1( u0_u9_u3_n155 ) , .A( u0_u9_u3_n167 ) );
  NAND2_X1 u0_u9_u3_U19 (.A1( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n142 ) , .A2( u0_u9_u3_n164 ) );
  NAND2_X1 u0_u9_u3_U20 (.ZN( u0_u9_u3_n132 ) , .A2( u0_u9_u3_n152 ) , .A1( u0_u9_u3_n156 ) );
  AND2_X1 u0_u9_u3_U21 (.A2( u0_u9_u3_n113 ) , .A1( u0_u9_u3_n114 ) , .ZN( u0_u9_u3_n151 ) );
  INV_X1 u0_u9_u3_U22 (.A( u0_u9_u3_n133 ) , .ZN( u0_u9_u3_n165 ) );
  INV_X1 u0_u9_u3_U23 (.A( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n170 ) );
  NAND2_X1 u0_u9_u3_U24 (.A1( u0_u9_u3_n107 ) , .A2( u0_u9_u3_n108 ) , .ZN( u0_u9_u3_n140 ) );
  NAND2_X1 u0_u9_u3_U25 (.ZN( u0_u9_u3_n117 ) , .A1( u0_u9_u3_n124 ) , .A2( u0_u9_u3_n148 ) );
  NAND2_X1 u0_u9_u3_U26 (.ZN( u0_u9_u3_n143 ) , .A1( u0_u9_u3_n165 ) , .A2( u0_u9_u3_n167 ) );
  INV_X1 u0_u9_u3_U27 (.A( u0_u9_u3_n130 ) , .ZN( u0_u9_u3_n177 ) );
  INV_X1 u0_u9_u3_U28 (.A( u0_u9_u3_n128 ) , .ZN( u0_u9_u3_n176 ) );
  INV_X1 u0_u9_u3_U29 (.A( u0_u9_u3_n155 ) , .ZN( u0_u9_u3_n174 ) );
  INV_X1 u0_u9_u3_U3 (.A( u0_u9_u3_n129 ) , .ZN( u0_u9_u3_n183 ) );
  INV_X1 u0_u9_u3_U30 (.A( u0_u9_u3_n139 ) , .ZN( u0_u9_u3_n185 ) );
  NOR2_X1 u0_u9_u3_U31 (.ZN( u0_u9_u3_n135 ) , .A2( u0_u9_u3_n141 ) , .A1( u0_u9_u3_n169 ) );
  OAI222_X1 u0_u9_u3_U32 (.C2( u0_u9_u3_n107 ) , .A2( u0_u9_u3_n108 ) , .B1( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n138 ) , .B2( u0_u9_u3_n146 ) , .C1( u0_u9_u3_n154 ) , .A1( u0_u9_u3_n164 ) );
  NOR4_X1 u0_u9_u3_U33 (.A4( u0_u9_u3_n157 ) , .A3( u0_u9_u3_n158 ) , .A2( u0_u9_u3_n159 ) , .A1( u0_u9_u3_n160 ) , .ZN( u0_u9_u3_n161 ) );
  AOI21_X1 u0_u9_u3_U34 (.B2( u0_u9_u3_n152 ) , .B1( u0_u9_u3_n153 ) , .ZN( u0_u9_u3_n158 ) , .A( u0_u9_u3_n164 ) );
  AOI21_X1 u0_u9_u3_U35 (.A( u0_u9_u3_n154 ) , .B2( u0_u9_u3_n155 ) , .B1( u0_u9_u3_n156 ) , .ZN( u0_u9_u3_n157 ) );
  AOI21_X1 u0_u9_u3_U36 (.A( u0_u9_u3_n149 ) , .B2( u0_u9_u3_n150 ) , .B1( u0_u9_u3_n151 ) , .ZN( u0_u9_u3_n159 ) );
  AOI211_X1 u0_u9_u3_U37 (.ZN( u0_u9_u3_n109 ) , .A( u0_u9_u3_n119 ) , .C2( u0_u9_u3_n129 ) , .B( u0_u9_u3_n138 ) , .C1( u0_u9_u3_n141 ) );
  AOI211_X1 u0_u9_u3_U38 (.B( u0_u9_u3_n119 ) , .A( u0_u9_u3_n120 ) , .C2( u0_u9_u3_n121 ) , .ZN( u0_u9_u3_n122 ) , .C1( u0_u9_u3_n179 ) );
  INV_X1 u0_u9_u3_U39 (.A( u0_u9_u3_n156 ) , .ZN( u0_u9_u3_n179 ) );
  INV_X1 u0_u9_u3_U4 (.A( u0_u9_u3_n140 ) , .ZN( u0_u9_u3_n182 ) );
  OAI22_X1 u0_u9_u3_U40 (.B1( u0_u9_u3_n118 ) , .ZN( u0_u9_u3_n120 ) , .A1( u0_u9_u3_n135 ) , .B2( u0_u9_u3_n154 ) , .A2( u0_u9_u3_n178 ) );
  AND3_X1 u0_u9_u3_U41 (.ZN( u0_u9_u3_n118 ) , .A2( u0_u9_u3_n124 ) , .A1( u0_u9_u3_n144 ) , .A3( u0_u9_u3_n152 ) );
  INV_X1 u0_u9_u3_U42 (.A( u0_u9_u3_n121 ) , .ZN( u0_u9_u3_n164 ) );
  NAND2_X1 u0_u9_u3_U43 (.ZN( u0_u9_u3_n133 ) , .A1( u0_u9_u3_n154 ) , .A2( u0_u9_u3_n164 ) );
  OAI211_X1 u0_u9_u3_U44 (.B( u0_u9_u3_n127 ) , .ZN( u0_u9_u3_n139 ) , .C1( u0_u9_u3_n150 ) , .C2( u0_u9_u3_n154 ) , .A( u0_u9_u3_n184 ) );
  INV_X1 u0_u9_u3_U45 (.A( u0_u9_u3_n125 ) , .ZN( u0_u9_u3_n184 ) );
  AOI221_X1 u0_u9_u3_U46 (.A( u0_u9_u3_n126 ) , .ZN( u0_u9_u3_n127 ) , .C2( u0_u9_u3_n132 ) , .C1( u0_u9_u3_n169 ) , .B2( u0_u9_u3_n170 ) , .B1( u0_u9_u3_n174 ) );
  OAI22_X1 u0_u9_u3_U47 (.A1( u0_u9_u3_n124 ) , .ZN( u0_u9_u3_n125 ) , .B2( u0_u9_u3_n145 ) , .A2( u0_u9_u3_n165 ) , .B1( u0_u9_u3_n167 ) );
  NOR2_X1 u0_u9_u3_U48 (.A1( u0_u9_u3_n113 ) , .ZN( u0_u9_u3_n131 ) , .A2( u0_u9_u3_n154 ) );
  NAND2_X1 u0_u9_u3_U49 (.A1( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n150 ) , .A2( u0_u9_u3_n99 ) );
  INV_X1 u0_u9_u3_U5 (.A( u0_u9_u3_n117 ) , .ZN( u0_u9_u3_n178 ) );
  NAND2_X1 u0_u9_u3_U50 (.A2( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n155 ) , .A1( u0_u9_u3_n97 ) );
  INV_X1 u0_u9_u3_U51 (.A( u0_u9_u3_n141 ) , .ZN( u0_u9_u3_n167 ) );
  AOI21_X1 u0_u9_u3_U52 (.B2( u0_u9_u3_n114 ) , .B1( u0_u9_u3_n146 ) , .A( u0_u9_u3_n154 ) , .ZN( u0_u9_u3_n94 ) );
  AOI21_X1 u0_u9_u3_U53 (.ZN( u0_u9_u3_n110 ) , .B2( u0_u9_u3_n142 ) , .B1( u0_u9_u3_n186 ) , .A( u0_u9_u3_n95 ) );
  INV_X1 u0_u9_u3_U54 (.A( u0_u9_u3_n145 ) , .ZN( u0_u9_u3_n186 ) );
  AOI21_X1 u0_u9_u3_U55 (.B1( u0_u9_u3_n124 ) , .A( u0_u9_u3_n149 ) , .B2( u0_u9_u3_n155 ) , .ZN( u0_u9_u3_n95 ) );
  INV_X1 u0_u9_u3_U56 (.A( u0_u9_u3_n149 ) , .ZN( u0_u9_u3_n169 ) );
  NAND2_X1 u0_u9_u3_U57 (.ZN( u0_u9_u3_n124 ) , .A1( u0_u9_u3_n96 ) , .A2( u0_u9_u3_n97 ) );
  NAND2_X1 u0_u9_u3_U58 (.A2( u0_u9_u3_n100 ) , .ZN( u0_u9_u3_n146 ) , .A1( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U59 (.A1( u0_u9_u3_n101 ) , .ZN( u0_u9_u3_n145 ) , .A2( u0_u9_u3_n99 ) );
  AOI221_X1 u0_u9_u3_U6 (.A( u0_u9_u3_n131 ) , .C2( u0_u9_u3_n132 ) , .C1( u0_u9_u3_n133 ) , .ZN( u0_u9_u3_n134 ) , .B1( u0_u9_u3_n143 ) , .B2( u0_u9_u3_n177 ) );
  NAND2_X1 u0_u9_u3_U60 (.A1( u0_u9_u3_n100 ) , .ZN( u0_u9_u3_n156 ) , .A2( u0_u9_u3_n99 ) );
  NAND2_X1 u0_u9_u3_U61 (.A2( u0_u9_u3_n101 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n148 ) );
  NAND2_X1 u0_u9_u3_U62 (.A1( u0_u9_u3_n100 ) , .A2( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n128 ) );
  NAND2_X1 u0_u9_u3_U63 (.A2( u0_u9_u3_n101 ) , .A1( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n152 ) );
  NAND2_X1 u0_u9_u3_U64 (.A2( u0_u9_u3_n101 ) , .ZN( u0_u9_u3_n114 ) , .A1( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U65 (.ZN( u0_u9_u3_n107 ) , .A1( u0_u9_u3_n97 ) , .A2( u0_u9_u3_n99 ) );
  NAND2_X1 u0_u9_u3_U66 (.A2( u0_u9_u3_n100 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n113 ) );
  NAND2_X1 u0_u9_u3_U67 (.A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n153 ) , .A2( u0_u9_u3_n97 ) );
  NAND2_X1 u0_u9_u3_U68 (.A2( u0_u9_u3_n103 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n130 ) );
  NAND2_X1 u0_u9_u3_U69 (.A2( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n144 ) , .A1( u0_u9_u3_n96 ) );
  OAI22_X1 u0_u9_u3_U7 (.B2( u0_u9_u3_n147 ) , .A2( u0_u9_u3_n148 ) , .ZN( u0_u9_u3_n160 ) , .B1( u0_u9_u3_n165 ) , .A1( u0_u9_u3_n168 ) );
  NAND2_X1 u0_u9_u3_U70 (.A1( u0_u9_u3_n102 ) , .A2( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n108 ) );
  NOR2_X1 u0_u9_u3_U71 (.A2( u0_u9_X_19 ) , .A1( u0_u9_X_20 ) , .ZN( u0_u9_u3_n99 ) );
  NOR2_X1 u0_u9_u3_U72 (.A2( u0_u9_X_21 ) , .A1( u0_u9_X_24 ) , .ZN( u0_u9_u3_n103 ) );
  NOR2_X1 u0_u9_u3_U73 (.A2( u0_u9_X_24 ) , .A1( u0_u9_u3_n171 ) , .ZN( u0_u9_u3_n97 ) );
  NOR2_X1 u0_u9_u3_U74 (.A2( u0_u9_X_23 ) , .ZN( u0_u9_u3_n141 ) , .A1( u0_u9_u3_n166 ) );
  NOR2_X1 u0_u9_u3_U75 (.A2( u0_u9_X_19 ) , .A1( u0_u9_u3_n172 ) , .ZN( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U76 (.A1( u0_u9_X_22 ) , .A2( u0_u9_X_23 ) , .ZN( u0_u9_u3_n154 ) );
  NAND2_X1 u0_u9_u3_U77 (.A1( u0_u9_X_23 ) , .ZN( u0_u9_u3_n149 ) , .A2( u0_u9_u3_n166 ) );
  NOR2_X1 u0_u9_u3_U78 (.A2( u0_u9_X_22 ) , .A1( u0_u9_X_23 ) , .ZN( u0_u9_u3_n121 ) );
  AND2_X1 u0_u9_u3_U79 (.A1( u0_u9_X_24 ) , .ZN( u0_u9_u3_n101 ) , .A2( u0_u9_u3_n171 ) );
  AND3_X1 u0_u9_u3_U8 (.A3( u0_u9_u3_n144 ) , .A2( u0_u9_u3_n145 ) , .A1( u0_u9_u3_n146 ) , .ZN( u0_u9_u3_n147 ) );
  AND2_X1 u0_u9_u3_U80 (.A1( u0_u9_X_19 ) , .ZN( u0_u9_u3_n102 ) , .A2( u0_u9_u3_n172 ) );
  AND2_X1 u0_u9_u3_U81 (.A1( u0_u9_X_21 ) , .A2( u0_u9_X_24 ) , .ZN( u0_u9_u3_n100 ) );
  AND2_X1 u0_u9_u3_U82 (.A2( u0_u9_X_19 ) , .A1( u0_u9_X_20 ) , .ZN( u0_u9_u3_n104 ) );
  INV_X1 u0_u9_u3_U83 (.A( u0_u9_X_22 ) , .ZN( u0_u9_u3_n166 ) );
  INV_X1 u0_u9_u3_U84 (.A( u0_u9_X_21 ) , .ZN( u0_u9_u3_n171 ) );
  INV_X1 u0_u9_u3_U85 (.A( u0_u9_X_20 ) , .ZN( u0_u9_u3_n172 ) );
  OR4_X1 u0_u9_u3_U86 (.ZN( u0_out9_10 ) , .A4( u0_u9_u3_n136 ) , .A3( u0_u9_u3_n137 ) , .A1( u0_u9_u3_n138 ) , .A2( u0_u9_u3_n139 ) );
  OAI222_X1 u0_u9_u3_U87 (.C1( u0_u9_u3_n128 ) , .ZN( u0_u9_u3_n137 ) , .B1( u0_u9_u3_n148 ) , .A2( u0_u9_u3_n150 ) , .B2( u0_u9_u3_n154 ) , .C2( u0_u9_u3_n164 ) , .A1( u0_u9_u3_n167 ) );
  OAI221_X1 u0_u9_u3_U88 (.A( u0_u9_u3_n134 ) , .B2( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n136 ) , .C1( u0_u9_u3_n149 ) , .B1( u0_u9_u3_n151 ) , .C2( u0_u9_u3_n183 ) );
  NAND4_X1 u0_u9_u3_U89 (.ZN( u0_out9_26 ) , .A4( u0_u9_u3_n109 ) , .A3( u0_u9_u3_n110 ) , .A2( u0_u9_u3_n111 ) , .A1( u0_u9_u3_n173 ) );
  INV_X1 u0_u9_u3_U9 (.A( u0_u9_u3_n143 ) , .ZN( u0_u9_u3_n168 ) );
  INV_X1 u0_u9_u3_U90 (.ZN( u0_u9_u3_n173 ) , .A( u0_u9_u3_n94 ) );
  OAI21_X1 u0_u9_u3_U91 (.ZN( u0_u9_u3_n111 ) , .B2( u0_u9_u3_n117 ) , .A( u0_u9_u3_n133 ) , .B1( u0_u9_u3_n176 ) );
  NAND4_X1 u0_u9_u3_U92 (.ZN( u0_out9_20 ) , .A4( u0_u9_u3_n122 ) , .A3( u0_u9_u3_n123 ) , .A1( u0_u9_u3_n175 ) , .A2( u0_u9_u3_n180 ) );
  INV_X1 u0_u9_u3_U93 (.A( u0_u9_u3_n126 ) , .ZN( u0_u9_u3_n180 ) );
  INV_X1 u0_u9_u3_U94 (.A( u0_u9_u3_n112 ) , .ZN( u0_u9_u3_n175 ) );
  NAND4_X1 u0_u9_u3_U95 (.ZN( u0_out9_1 ) , .A4( u0_u9_u3_n161 ) , .A3( u0_u9_u3_n162 ) , .A2( u0_u9_u3_n163 ) , .A1( u0_u9_u3_n185 ) );
  NAND2_X1 u0_u9_u3_U96 (.ZN( u0_u9_u3_n163 ) , .A2( u0_u9_u3_n170 ) , .A1( u0_u9_u3_n176 ) );
  AOI22_X1 u0_u9_u3_U97 (.B2( u0_u9_u3_n140 ) , .B1( u0_u9_u3_n141 ) , .A2( u0_u9_u3_n142 ) , .ZN( u0_u9_u3_n162 ) , .A1( u0_u9_u3_n177 ) );
  NAND3_X1 u0_u9_u3_U98 (.A1( u0_u9_u3_n114 ) , .ZN( u0_u9_u3_n115 ) , .A2( u0_u9_u3_n145 ) , .A3( u0_u9_u3_n153 ) );
  NAND3_X1 u0_u9_u3_U99 (.ZN( u0_u9_u3_n129 ) , .A2( u0_u9_u3_n144 ) , .A1( u0_u9_u3_n153 ) , .A3( u0_u9_u3_n182 ) );
  INV_X1 u0_uk_U10 (.A( u0_uk_n252 ) , .ZN( u0_uk_n31 ) );
  NAND2_X1 u0_uk_U1009 (.A1( u0_key_r_46 ) , .A2( u0_uk_n60 ) , .ZN( u0_uk_n890 ) );
  OAI21_X1 u0_uk_U1012 (.ZN( u0_K10_21 ) , .A( u0_uk_n1020 ) , .B2( u0_uk_n228 ) , .B1( u0_uk_n31 ) );
  OAI22_X1 u0_uk_U102 (.ZN( u0_K7_5 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n384 ) , .B2( u0_uk_n401 ) );
  OAI21_X1 u0_uk_U1024 (.ZN( u0_K8_46 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n326 ) , .A( u0_uk_n744 ) );
  NAND2_X1 u0_uk_U1025 (.A1( u0_uk_K_r6_37 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n744 ) );
  OAI21_X1 u0_uk_U104 (.ZN( u0_K4_5 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n502 ) , .A( u0_uk_n821 ) );
  NAND2_X1 u0_uk_U105 (.A1( u0_uk_K_r2_53 ) , .ZN( u0_uk_n821 ) , .A2( u0_uk_n99 ) );
  INV_X1 u0_uk_U1066 (.A( u0_key_r_33 ) , .ZN( u0_uk_n691 ) );
  INV_X1 u0_uk_U1101 (.ZN( u0_K2_10 ) , .A( u0_uk_n868 ) );
  AOI22_X1 u0_uk_U1102 (.B2( u0_uk_K_r0_34 ) , .A2( u0_uk_K_r0_55 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n868 ) );
  INV_X1 u0_uk_U1109 (.ZN( u0_K11_8 ) , .A( u0_uk_n982 ) );
  AOI22_X1 u0_uk_U1110 (.B2( u0_uk_K_r9_12 ) , .A2( u0_uk_K_r9_18 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n982 ) );
  INV_X1 u0_uk_U1111 (.ZN( u0_K11_12 ) , .A( u0_uk_n1003 ) );
  AOI22_X1 u0_uk_U1112 (.B2( u0_uk_K_r9_25 ) , .A2( u0_uk_K_r9_6 ) , .ZN( u0_uk_n1003 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n207 ) );
  INV_X1 u0_uk_U1119 (.ZN( u0_K2_7 ) , .A( u0_uk_n855 ) );
  INV_X1 u0_uk_U1123 (.ZN( u0_K7_13 ) , .A( u0_uk_n783 ) );
  AOI22_X1 u0_uk_U1124 (.B2( u0_uk_K_r5_26 ) , .A2( u0_uk_K_r5_48 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n188 ) , .ZN( u0_uk_n783 ) );
  INV_X1 u0_uk_U1135 (.ZN( u0_K4_2 ) , .A( u0_uk_n828 ) );
  AOI22_X1 u0_uk_U1136 (.B2( u0_uk_K_r2_26 ) , .A2( u0_uk_K_r2_46 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n148 ) , .ZN( u0_uk_n828 ) );
  INV_X1 u0_uk_U1137 (.ZN( u0_K4_20 ) , .A( u0_uk_n835 ) );
  AOI22_X1 u0_uk_U1138 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_33 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n208 ) , .ZN( u0_uk_n835 ) );
  INV_X1 u0_uk_U1143 (.ZN( u0_K13_12 ) , .A( u0_uk_n958 ) );
  AOI22_X1 u0_uk_U1144 (.B2( u0_uk_K_r11_34 ) , .A2( u0_uk_K_r11_54 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n958 ) );
  INV_X1 u0_uk_U115 (.ZN( u0_K11_47 ) , .A( u0_uk_n985 ) );
  AOI22_X1 u0_uk_U116 (.B2( u0_uk_K_r9_15 ) , .A2( u0_uk_K_r9_23 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n985 ) );
  OAI22_X1 u0_uk_U118 (.ZN( u0_K8_47 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n327 ) );
  OAI22_X1 u0_uk_U119 (.ZN( u0_K7_47 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n388 ) , .A2( u0_uk_n402 ) );
  OAI22_X1 u0_uk_U127 (.ZN( u0_K4_15 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n502 ) , .B2( u0_uk_n530 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U13 (.A( u0_uk_n252 ) , .ZN( u0_uk_n60 ) );
  INV_X1 u0_uk_U130 (.ZN( u0_K13_15 ) , .A( u0_uk_n956 ) );
  AOI22_X1 u0_uk_U131 (.B2( u0_uk_K_r11_11 ) , .A2( u0_uk_K_r11_48 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n956 ) );
  OAI22_X1 u0_uk_U132 (.ZN( u0_K7_15 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n364 ) , .A2( u0_uk_n404 ) );
  INV_X1 u0_uk_U136 (.ZN( u0_K13_19 ) , .A( u0_uk_n953 ) );
  AOI22_X1 u0_uk_U137 (.B2( u0_uk_K_r11_19 ) , .A2( u0_uk_K_r11_39 ) , .B1( u0_uk_n207 ) , .A1( u0_uk_n94 ) , .ZN( u0_uk_n953 ) );
  OAI22_X1 u0_uk_U139 (.ZN( u0_K11_15 ) , .A1( u0_uk_n147 ) , .A2( u0_uk_n197 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U14 (.A( u0_uk_n222 ) , .ZN( u0_uk_n94 ) );
  NAND2_X1 u0_uk_U141 (.A1( u0_uk_K_r4_48 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n798 ) );
  INV_X1 u0_uk_U151 (.ZN( u0_K11_19 ) , .A( u0_uk_n1000 ) );
  AOI22_X1 u0_uk_U152 (.B2( u0_uk_K_r9_10 ) , .A2( u0_uk_K_r9_48 ) , .ZN( u0_uk_n1000 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n220 ) );
  OAI22_X1 u0_uk_U155 (.ZN( u0_K7_19 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n383 ) , .B2( u0_uk_n393 ) );
  OAI22_X1 u0_uk_U156 (.ZN( u0_K4_19 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n511 ) , .B2( u0_uk_n523 ) );
  INV_X1 u0_uk_U16 (.ZN( u0_uk_n110 ) , .A( u0_uk_n222 ) );
  INV_X1 u0_uk_U17 (.ZN( u0_uk_n100 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U177 (.ZN( u0_K13_14 ) , .A2( u0_uk_n108 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n132 ) , .B1( u0_uk_n242 ) );
  INV_X1 u0_uk_U180 (.ZN( u0_K11_14 ) , .A( u0_uk_n1002 ) );
  OAI21_X1 u0_uk_U182 (.ZN( u0_K10_24 ) , .A( u0_uk_n1017 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n259 ) );
  NAND2_X1 u0_uk_U183 (.A1( u0_uk_K_r8_40 ) , .ZN( u0_uk_n1017 ) , .A2( u0_uk_n11 ) );
  INV_X1 u0_uk_U19 (.ZN( u0_uk_n118 ) , .A( u0_uk_n214 ) );
  NAND2_X1 u0_uk_U194 (.A1( u0_uk_K_r11_28 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n945 ) );
  INV_X1 u0_uk_U195 (.ZN( u0_K7_24 ) , .A( u0_uk_n776 ) );
  AOI22_X1 u0_uk_U196 (.B2( u0_uk_K_r5_18 ) , .A2( u0_uk_K_r5_40 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n776 ) );
  INV_X1 u0_uk_U198 (.ZN( u0_K3_24 ) , .A( u0_uk_n851 ) );
  AOI22_X1 u0_uk_U199 (.B2( u0_uk_K_r1_17 ) , .A2( u0_uk_K_r1_41 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n851 ) );
  INV_X1 u0_uk_U20 (.ZN( u0_uk_n109 ) , .A( u0_uk_n214 ) );
  OAI21_X1 u0_uk_U205 (.ZN( u0_K4_30 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n513 ) , .A( u0_uk_n827 ) );
  NAND2_X1 u0_uk_U206 (.A1( u0_uk_K_r2_28 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n827 ) );
  INV_X1 u0_uk_U207 (.ZN( u0_K15_30 ) , .A( u0_uk_n919 ) );
  AOI22_X1 u0_uk_U208 (.B2( u0_uk_K_r13_0 ) , .A2( u0_uk_K_r13_38 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n919 ) );
  INV_X1 u0_uk_U21 (.ZN( u0_uk_n102 ) , .A( u0_uk_n162 ) );
  INV_X1 u0_uk_U210 (.ZN( u0_K4_31 ) , .A( u0_uk_n826 ) );
  INV_X1 u0_uk_U218 (.ZN( u0_K11_31 ) , .A( u0_uk_n992 ) );
  AOI22_X1 u0_uk_U219 (.B2( u0_uk_K_r9_22 ) , .A2( u0_uk_K_r9_30 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n992 ) );
  INV_X1 u0_uk_U22 (.ZN( u0_uk_n128 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U220 (.ZN( u0_K2_31 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n613 ) , .B2( u0_uk_n628 ) );
  INV_X1 u0_uk_U221 (.ZN( u0_K11_39 ) , .A( u0_uk_n988 ) );
  AOI22_X1 u0_uk_U222 (.B2( u0_uk_K_r9_30 ) , .A2( u0_uk_K_r9_7 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n988 ) );
  OAI22_X1 u0_uk_U228 (.ZN( u0_K6_31 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n428 ) , .B2( u0_uk_n433 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U24 (.ZN( u0_uk_n11 ) , .A( u0_uk_n242 ) );
  NAND2_X1 u0_uk_U240 (.A1( u0_uk_K_r10_16 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n969 ) );
  OAI21_X1 u0_uk_U247 (.ZN( u0_K8_44 ) , .B1( u0_uk_n117 ) , .B2( u0_uk_n320 ) , .A( u0_uk_n745 ) );
  NAND2_X1 u0_uk_U248 (.A1( u0_uk_K_r6_0 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n745 ) );
  OAI22_X1 u0_uk_U249 (.ZN( u0_K8_48 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n223 ) , .B2( u0_uk_n347 ) , .A2( u0_uk_n354 ) );
  INV_X1 u0_uk_U25 (.ZN( u0_uk_n146 ) , .A( u0_uk_n148 ) );
  INV_X1 u0_uk_U26 (.ZN( u0_uk_n129 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U261 (.ZN( u0_K11_44 ) , .A2( u0_uk_n185 ) , .B2( u0_uk_n205 ) , .A1( u0_uk_n242 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U266 (.ZN( u0_K7_44 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n378 ) , .B2( u0_uk_n399 ) );
  OAI22_X1 u0_uk_U267 (.ZN( u0_K7_48 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n257 ) , .A2( u0_uk_n367 ) , .B2( u0_uk_n387 ) );
  BUF_X1 u0_uk_U28 (.Z( u0_uk_n147 ) , .A( u0_uk_n250 ) );
  INV_X1 u0_uk_U288 (.ZN( u0_K7_8 ) , .A( u0_uk_n763 ) );
  BUF_X1 u0_uk_U29 (.Z( u0_uk_n162 ) , .A( u0_uk_n217 ) );
  INV_X1 u0_uk_U291 (.ZN( u0_K4_8 ) , .A( u0_uk_n819 ) );
  AOI22_X1 u0_uk_U292 (.B2( u0_uk_K_r2_41 ) , .A2( u0_uk_K_r2_46 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n819 ) );
  OAI22_X1 u0_uk_U293 (.ZN( u0_K3_8 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n562 ) , .A2( u0_uk_n578 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U3 (.ZN( u0_uk_n142 ) , .A( u0_uk_n191 ) );
  BUF_X1 u0_uk_U30 (.Z( u0_uk_n161 ) , .A( u0_uk_n238 ) );
  INV_X1 u0_uk_U302 (.ZN( u0_K4_26 ) , .A( u0_uk_n831 ) );
  AOI22_X1 u0_uk_U303 (.B2( u0_uk_K_r2_16 ) , .A2( u0_uk_K_r2_7 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n831 ) );
  INV_X1 u0_uk_U304 (.ZN( u0_K15_26 ) , .A( u0_uk_n920 ) );
  AOI22_X1 u0_uk_U305 (.B2( u0_uk_K_r13_38 ) , .A2( u0_uk_K_r13_44 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n920 ) );
  OAI21_X1 u0_uk_U306 (.ZN( u0_K6_26 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n419 ) , .A( u0_uk_n795 ) );
  NAND2_X1 u0_uk_U307 (.A1( u0_uk_K_r4_35 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n795 ) );
  OAI22_X1 u0_uk_U313 (.ZN( u0_K2_26 ) , .A1( u0_uk_n164 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n593 ) , .B2( u0_uk_n599 ) );
  BUF_X1 u0_uk_U32 (.Z( u0_uk_n148 ) , .A( u0_uk_n240 ) );
  INV_X1 u0_uk_U333 (.ZN( u0_K7_46 ) , .A( u0_uk_n765 ) );
  BUF_X1 u0_uk_U34 (.Z( u0_uk_n164 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U340 (.ZN( u0_K7_4 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n361 ) , .B2( u0_uk_n384 ) );
  NAND2_X1 u0_uk_U344 (.A1( u0_uk_K_r3_4 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n804 ) );
  INV_X1 u0_uk_U345 (.ZN( u0_K4_4 ) , .A( u0_uk_n822 ) );
  AOI22_X1 u0_uk_U346 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_18 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n822 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U347 (.ZN( u0_K3_4 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n557 ) , .B2( u0_uk_n565 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U352 (.ZN( u0_K6_40 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n438 ) , .A2( u0_uk_n446 ) );
  INV_X1 u0_uk_U353 (.ZN( u0_K11_46 ) , .A( u0_uk_n986 ) );
  AOI22_X1 u0_uk_U354 (.B2( u0_uk_K_r9_45 ) , .A2( u0_uk_K_r9_9 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n208 ) , .ZN( u0_uk_n986 ) );
  OAI22_X1 u0_uk_U362 (.ZN( u0_K11_40 ) , .B2( u0_uk_n216 ) , .A2( u0_uk_n224 ) , .A1( u0_uk_n240 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U366 (.ZN( u0_K2_40 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n592 ) , .A2( u0_uk_n623 ) );
  OAI21_X1 u0_uk_U369 (.ZN( u0_K2_33 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n600 ) , .A( u0_uk_n859 ) );
  BUF_X1 u0_uk_U37 (.Z( u0_uk_n182 ) , .A( u0_uk_n214 ) );
  NAND2_X1 u0_uk_U370 (.A1( u0_uk_K_r0_31 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n859 ) );
  OAI22_X1 u0_uk_U375 (.ZN( u0_K6_28 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n411 ) , .B2( u0_uk_n438 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U38 (.Z( u0_uk_n203 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U381 (.ZN( u0_K15_28 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n33 ) , .A2( u0_uk_n5 ) );
  OAI22_X1 u0_uk_U389 (.ZN( u0_K3_1 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n568 ) , .B2( u0_uk_n573 ) , .B1( u0_uk_n60 ) );
  BUF_X1 u0_uk_U39 (.Z( u0_uk_n202 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U390 (.ZN( u0_K2_1 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n583 ) , .B2( u0_uk_n604 ) );
  OAI22_X1 u0_uk_U392 (.ZN( u0_K13_16 ) , .A1( u0_uk_n118 ) , .A2( u0_uk_n122 ) , .B2( u0_uk_n127 ) , .B1( u0_uk_n242 ) );
  OAI21_X1 u0_uk_U398 (.ZN( u0_K3_16 ) , .B1( u0_uk_n102 ) , .B2( u0_uk_n540 ) , .A( u0_uk_n853 ) );
  INV_X1 u0_uk_U4 (.ZN( u0_uk_n145 ) , .A( u0_uk_n242 ) );
  OAI22_X1 u0_uk_U401 (.ZN( u0_K4_16 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n525 ) , .B2( u0_uk_n529 ) );
  OAI22_X1 u0_uk_U406 (.ZN( u0_K13_9 ) , .A2( u0_uk_n115 ) , .B2( u0_uk_n127 ) , .A1( u0_uk_n230 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U408 (.ZN( u0_K11_9 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n195 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n225 ) );
  BUF_X1 u0_uk_U41 (.Z( u0_uk_n214 ) , .A( u0_uk_n257 ) );
  INV_X1 u0_uk_U410 (.ZN( u0_K2_28 ) , .A( u0_uk_n861 ) );
  AOI22_X1 u0_uk_U411 (.B2( u0_uk_K_r0_15 ) , .A2( u0_uk_K_r0_49 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n861 ) );
  BUF_X1 u0_uk_U42 (.Z( u0_uk_n238 ) , .A( u0_uk_n252 ) );
  OAI22_X1 u0_uk_U420 (.ZN( u0_K7_9 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n390 ) , .B2( u0_uk_n397 ) );
  OAI22_X1 u0_uk_U421 (.ZN( u0_K4_9 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n519 ) , .B2( u0_uk_n529 ) );
  OAI21_X1 u0_uk_U422 (.ZN( u0_K3_9 ) , .B1( u0_uk_n209 ) , .B2( u0_uk_n563 ) , .A( u0_uk_n840 ) );
  NAND2_X1 u0_uk_U423 (.A1( u0_uk_K_r1_18 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n840 ) );
  OAI22_X1 u0_uk_U424 (.ZN( u0_K2_9 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n597 ) , .A2( u0_uk_n626 ) );
  BUF_X1 u0_uk_U43 (.Z( u0_uk_n220 ) , .A( u0_uk_n251 ) );
  OAI21_X1 u0_uk_U432 (.ZN( u0_K7_16 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n362 ) , .A( u0_uk_n782 ) );
  NAND2_X1 u0_uk_U433 (.A1( u0_uk_K_r5_32 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n782 ) );
  OAI22_X1 u0_uk_U436 (.ZN( u0_K11_33 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n199 ) , .B2( u0_uk_n205 ) , .B1( u0_uk_n222 ) );
  BUF_X1 u0_uk_U44 (.Z( u0_uk_n209 ) , .A( u0_uk_n252 ) );
  OAI22_X1 u0_uk_U448 (.ZN( u0_K6_33 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n425 ) , .B2( u0_uk_n430 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U449 (.ZN( u0_K4_33 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n532 ) , .B2( u0_uk_n539 ) );
  BUF_X1 u0_uk_U45 (.A( u0_uk_n238 ) , .Z( u0_uk_n240 ) );
  BUF_X1 u0_uk_U46 (.A( u0_uk_n162 ) , .Z( u0_uk_n223 ) );
  OAI21_X1 u0_uk_U461 (.ZN( u0_K6_37 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n420 ) , .A( u0_uk_n791 ) );
  NAND2_X1 u0_uk_U462 (.A1( u0_uk_K_r4_38 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n791 ) );
  BUF_X1 u0_uk_U47 (.Z( u0_uk_n217 ) , .A( u0_uk_n240 ) );
  NAND2_X1 u0_uk_U471 (.A1( u0_uk_K_r8_21 ) , .ZN( u0_uk_n1010 ) , .A2( u0_uk_n11 ) );
  OAI21_X1 u0_uk_U477 (.ZN( u0_K6_29 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n446 ) , .A( u0_uk_n794 ) );
  NAND2_X1 u0_uk_U478 (.A1( u0_uk_K_r4_0 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n794 ) );
  BUF_X1 u0_uk_U48 (.Z( u0_uk_n222 ) , .A( u0_uk_n250 ) );
  OAI22_X1 u0_uk_U481 (.ZN( u0_K2_29 ) , .A1( u0_uk_n188 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n606 ) , .A2( u0_uk_n621 ) );
  OAI22_X1 u0_uk_U482 (.ZN( u0_K15_29 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n21 ) , .A2( u0_uk_n39 ) );
  OAI22_X1 u0_uk_U491 (.ZN( u0_K3_2 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n552 ) , .B2( u0_uk_n557 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U492 (.ZN( u0_K2_2 ) , .A1( u0_uk_n164 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n583 ) , .B2( u0_uk_n615 ) );
  BUF_X1 u0_uk_U50 (.A( u0_uk_n162 ) , .Z( u0_uk_n213 ) );
  OAI21_X1 u0_uk_U501 (.ZN( u0_K13_17 ) , .B2( u0_uk_n115 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n955 ) );
  NAND2_X1 u0_uk_U502 (.A1( u0_uk_K_r11_27 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n955 ) );
  INV_X1 u0_uk_U508 (.ZN( u0_K11_17 ) , .A( u0_uk_n1001 ) );
  BUF_X1 u0_uk_U51 (.A( u0_uk_n161 ) , .Z( u0_uk_n242 ) );
  OAI22_X1 u0_uk_U512 (.ZN( u0_K7_17 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n370 ) , .B2( u0_uk_n400 ) );
  OAI21_X1 u0_uk_U513 (.ZN( u0_K4_17 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n519 ) , .A( u0_uk_n838 ) );
  NAND2_X1 u0_uk_U514 (.A1( u0_uk_K_r2_27 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n838 ) );
  INV_X1 u0_uk_U516 (.ZN( u0_K4_29 ) , .A( u0_uk_n829 ) );
  AOI22_X1 u0_uk_U517 (.B2( u0_uk_K_r2_31 ) , .A2( u0_uk_K_r2_36 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n829 ) , .A1( u0_uk_n94 ) );
  BUF_X1 u0_uk_U52 (.Z( u0_uk_n207 ) , .A( u0_uk_n217 ) );
  INV_X1 u0_uk_U522 (.ZN( u0_K7_12 ) , .A( u0_uk_n784 ) );
  AOI22_X1 u0_uk_U523 (.B2( u0_uk_K_r5_17 ) , .A2( u0_uk_K_r5_39 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n784 ) );
  OAI22_X1 u0_uk_U526 (.ZN( u0_K4_12 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n517 ) );
  BUF_X1 u0_uk_U54 (.Z( u0_uk_n251 ) , .A( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U548 (.ZN( u0_K2_36 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n250 ) , .A2( u0_uk_n600 ) , .B2( u0_uk_n616 ) );
  BUF_X1 u0_uk_U55 (.A( u0_uk_n250 ) , .Z( u0_uk_n252 ) );
  OAI22_X1 u0_uk_U556 (.ZN( u0_K11_38 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n210 ) , .B2( u0_uk_n218 ) );
  BUF_X1 u0_uk_U56 (.Z( u0_uk_n250 ) , .A( u0_uk_n257 ) );
  INV_X1 u0_uk_U560 (.ZN( u0_K11_36 ) , .A( u0_uk_n990 ) );
  OAI22_X1 u0_uk_U567 (.ZN( u0_K6_38 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n433 ) , .B2( u0_uk_n440 ) , .B1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U575 (.ZN( u0_K11_10 ) , .A( u0_uk_n1004 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n225 ) );
  INV_X1 u0_uk_U577 (.ZN( u0_K13_10 ) , .A( u0_uk_n960 ) );
  INV_X1 u0_uk_U584 (.ZN( u0_K4_10 ) , .A( u0_uk_n839 ) );
  OAI22_X1 u0_uk_U588 (.ZN( u0_K3_22 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n542 ) , .B2( u0_uk_n577 ) );
  INV_X1 u0_uk_U590 (.ZN( u0_K13_22 ) , .A( u0_uk_n949 ) );
  AOI22_X1 u0_uk_U591 (.B2( u0_uk_K_r11_10 ) , .A2( u0_uk_K_r11_47 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n949 ) );
  INV_X1 u0_uk_U592 (.ZN( u0_K11_22 ) , .A( u0_uk_n997 ) );
  AOI22_X1 u0_uk_U593 (.B2( u0_uk_K_r9_13 ) , .A2( u0_uk_K_r9_19 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n997 ) );
  INV_X1 u0_uk_U594 (.ZN( u0_K10_22 ) , .A( u0_uk_n1019 ) );
  INV_X1 u0_uk_U60 (.ZN( u0_K11_34 ) , .A( u0_uk_n991 ) );
  OAI22_X1 u0_uk_U604 (.ZN( u0_K11_35 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n185 ) , .B2( u0_uk_n193 ) , .B1( u0_uk_n222 ) );
  AOI22_X1 u0_uk_U61 (.B2( u0_uk_K_r9_45 ) , .A2( u0_uk_K_r9_49 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n991 ) );
  OAI22_X1 u0_uk_U618 (.ZN( u0_K6_35 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n412 ) , .B2( u0_uk_n419 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U627 (.ZN( u0_K11_11 ) , .A1( u0_uk_n145 ) , .A2( u0_uk_n206 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n214 ) );
  INV_X1 u0_uk_U628 (.ZN( u0_K13_11 ) , .A( u0_uk_n959 ) );
  AOI22_X1 u0_uk_U629 (.B2( u0_uk_K_r11_17 ) , .A2( u0_uk_K_r11_54 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n959 ) );
  OAI22_X1 u0_uk_U633 (.ZN( u0_K7_11 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n383 ) , .B2( u0_uk_n400 ) );
  OAI22_X1 u0_uk_U634 (.ZN( u0_K3_11 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n573 ) , .A2( u0_uk_n578 ) );
  NAND2_X1 u0_uk_U636 (.A1( u0_uk_K_r0_25 ) , .A2( u0_uk_n109 ) , .ZN( u0_uk_n867 ) );
  INV_X1 u0_uk_U643 (.ZN( u0_K4_23 ) , .A( u0_uk_n833 ) );
  AOI22_X1 u0_uk_U644 (.B2( u0_uk_K_r2_18 ) , .A2( u0_uk_K_r2_55 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n833 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U651 (.ZN( u0_K7_43 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n374 ) , .A2( u0_uk_n403 ) );
  OAI22_X1 u0_uk_U668 (.ZN( u0_K11_43 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n184 ) , .B2( u0_uk_n226 ) , .B1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U68 (.ZN( u0_K6_34 ) , .B1( u0_uk_n118 ) , .B2( u0_uk_n417 ) , .A( u0_uk_n792 ) );
  OAI21_X1 u0_uk_U682 (.ZN( u0_K11_7 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n197 ) , .A( u0_uk_n983 ) );
  NAND2_X1 u0_uk_U683 (.A1( u0_uk_K_r9_33 ) , .A2( u0_uk_n146 ) , .ZN( u0_uk_n983 ) );
  OAI22_X1 u0_uk_U684 (.ZN( u0_K4_7 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n531 ) , .A2( u0_uk_n535 ) , .A1( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U686 (.ZN( u0_K15_25 ) , .B2( u0_uk_n12 ) , .B1( u0_uk_n147 ) , .A( u0_uk_n921 ) );
  NAND2_X1 u0_uk_U687 (.A1( u0_uk_K_r13_22 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n921 ) );
  NAND2_X1 u0_uk_U69 (.A1( u0_uk_K_r4_49 ) , .ZN( u0_uk_n792 ) , .A2( u0_uk_n83 ) );
  NAND2_X1 u0_uk_U693 (.A1( u0_uk_K_r0_22 ) , .ZN( u0_uk_n863 ) , .A2( u0_uk_n94 ) );
  INV_X1 u0_uk_U697 (.ZN( u0_K8_43 ) , .A( u0_uk_n746 ) );
  OAI22_X1 u0_uk_U70 (.ZN( u0_K4_34 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n208 ) , .A2( u0_uk_n506 ) , .B2( u0_uk_n522 ) );
  INV_X1 u0_uk_U702 (.ZN( u0_K4_3 ) , .A( u0_uk_n824 ) );
  AOI22_X1 u0_uk_U703 (.A2( u0_uk_K_r2_4 ) , .B2( u0_uk_K_r2_41 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n824 ) , .B1( u0_uk_n99 ) );
  INV_X1 u0_uk_U704 (.ZN( u0_K13_7 ) , .A( u0_uk_n939 ) );
  INV_X1 u0_uk_U712 (.ZN( u0_K4_25 ) , .A( u0_uk_n832 ) );
  OAI22_X1 u0_uk_U716 (.ZN( u0_K4_32 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n508 ) , .A2( u0_uk_n532 ) );
  OAI22_X1 u0_uk_U719 (.ZN( u0_K11_32 ) , .A2( u0_uk_n198 ) , .A1( u0_uk_n208 ) , .B2( u0_uk_n218 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U72 (.A1( u0_uk_K_r1_36 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n848 ) );
  OAI22_X1 u0_uk_U721 (.ZN( u0_K6_32 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n424 ) , .B2( u0_uk_n440 ) );
  OAI22_X1 u0_uk_U729 (.ZN( u0_K11_42 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n186 ) , .B2( u0_uk_n194 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U735 (.ZN( u0_K2_42 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n584 ) , .B2( u0_uk_n592 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U740 (.ZN( u0_K2_32 ) , .A( u0_uk_n860 ) );
  AOI22_X1 u0_uk_U741 (.B2( u0_uk_K_r0_15 ) , .A2( u0_uk_K_r0_36 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n231 ) , .ZN( u0_uk_n860 ) );
  NAND2_X1 u0_uk_U745 (.A1( u0_uk_K_r12_42 ) , .A2( u0_uk_n129 ) , .ZN( u0_uk_n936 ) );
  NAND2_X1 u0_uk_U748 (.A1( u0_uk_K_r8_43 ) , .ZN( u0_uk_n1016 ) , .A2( u0_uk_n11 ) );
  OAI21_X1 u0_uk_U75 (.ZN( u0_K11_23 ) , .B2( u0_uk_n190 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n996 ) );
  OAI22_X1 u0_uk_U752 (.ZN( u0_K11_13 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n196 ) , .B2( u0_uk_n200 ) );
  NAND2_X1 u0_uk_U76 (.A1( u0_uk_K_r9_27 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n996 ) );
  OAI22_X1 u0_uk_U766 (.ZN( u0_K4_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n511 ) , .B2( u0_uk_n517 ) );
  OAI21_X1 u0_uk_U77 (.ZN( u0_K10_23 ) , .A( u0_uk_n1018 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n268 ) );
  OAI22_X1 u0_uk_U771 (.ZN( u0_K15_27 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n23 ) , .A2( u0_uk_n41 ) );
  OAI22_X1 u0_uk_U772 (.ZN( u0_K4_13 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n530 ) , .A2( u0_uk_n534 ) , .A1( u0_uk_n60 ) );
  INV_X1 u0_uk_U776 (.ZN( u0_K2_27 ) , .A( u0_uk_n862 ) );
  AOI22_X1 u0_uk_U777 (.B2( u0_uk_K_r0_28 ) , .A2( u0_uk_K_r0_7 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n862 ) );
  NAND2_X1 u0_uk_U78 (.A1( u0_uk_K_r8_13 ) , .ZN( u0_uk_n1018 ) , .A2( u0_uk_n252 ) );
  INV_X1 u0_uk_U780 (.ZN( u0_K13_13 ) , .A( u0_uk_n957 ) );
  AOI22_X1 u0_uk_U781 (.B2( u0_uk_K_r11_11 ) , .A2( u0_uk_K_r11_6 ) , .B1( u0_uk_n207 ) , .A1( u0_uk_n94 ) , .ZN( u0_uk_n957 ) );
  INV_X1 u0_uk_U782 (.ZN( u0_K13_21 ) , .A( u0_uk_n950 ) );
  INV_X1 u0_uk_U786 (.ZN( u0_K6_21 ) , .A( u0_uk_n797 ) );
  AOI22_X1 u0_uk_U787 (.B2( u0_uk_K_r4_11 ) , .A2( u0_uk_K_r4_5 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n797 ) );
  OAI21_X1 u0_uk_U790 (.ZN( u0_K7_21 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n362 ) , .A( u0_uk_n779 ) );
  NAND2_X1 u0_uk_U791 (.A1( u0_uk_K_r5_19 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n779 ) );
  OAI21_X1 u0_uk_U800 (.ZN( u0_K7_1 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n396 ) , .A( u0_uk_n781 ) );
  NAND2_X1 u0_uk_U801 (.A1( u0_uk_K_r5_10 ) , .A2( u0_uk_n147 ) , .ZN( u0_uk_n781 ) );
  OAI21_X1 u0_uk_U802 (.ZN( u0_K4_1 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n535 ) , .A( u0_uk_n836 ) );
  NAND2_X1 u0_uk_U803 (.A1( u0_uk_K_r2_25 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n836 ) );
  OAI21_X1 u0_uk_U804 (.ZN( u0_K4_18 ) , .B2( u0_uk_n510 ) , .A( u0_uk_n837 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U805 (.A1( u0_uk_K_r2_20 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n837 ) );
  OAI22_X1 u0_uk_U807 (.ZN( u0_K7_18 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n392 ) , .A2( u0_uk_n405 ) );
  OAI21_X1 u0_uk_U808 (.ZN( u0_K13_20 ) , .B2( u0_uk_n126 ) , .B1( u0_uk_n92 ) , .A( u0_uk_n951 ) );
  NAND2_X1 u0_uk_U809 (.A1( u0_uk_K_r11_33 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n951 ) );
  OAI21_X1 u0_uk_U819 (.ZN( u0_K13_18 ) , .B2( u0_uk_n108 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n954 ) );
  NAND2_X1 u0_uk_U820 (.A1( u0_uk_K_r11_20 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n954 ) );
  OAI22_X1 u0_uk_U821 (.ZN( u0_K3_20 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n562 ) , .B2( u0_uk_n568 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U829 (.ZN( u0_K11_20 ) , .A( u0_uk_n999 ) );
  INV_X1 u0_uk_U833 (.ZN( u0_K7_20 ) , .A( u0_uk_n780 ) );
  OAI21_X1 u0_uk_U838 (.ZN( u0_K4_22 ) , .B2( u0_uk_n531 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n834 ) );
  OAI21_X1 u0_uk_U84 (.ZN( u0_K11_41 ) , .B2( u0_uk_n186 ) , .B1( u0_uk_n203 ) , .A( u0_uk_n987 ) );
  OAI22_X1 u0_uk_U849 (.ZN( u0_K7_3 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n371 ) , .B2( u0_uk_n393 ) );
  NAND2_X1 u0_uk_U85 (.A1( u0_uk_K_r9_31 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n987 ) );
  INV_X1 u0_uk_U854 (.ZN( u0_K7_6 ) , .A( u0_uk_n764 ) );
  AOI22_X1 u0_uk_U855 (.B2( u0_uk_K_r5_39 ) , .A2( u0_uk_K_r5_4 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n764 ) );
  OAI21_X1 u0_uk_U858 (.ZN( u0_K3_3 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n540 ) , .A( u0_uk_n846 ) );
  NAND2_X1 u0_uk_U859 (.A1( u0_uk_K_r1_47 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n846 ) );
  INV_X1 u0_uk_U86 (.ZN( u0_K2_41 ) , .A( u0_uk_n858 ) );
  NAND2_X1 u0_uk_U863 (.A1( u0_uk_K_r5_41 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n773 ) );
  AOI22_X1 u0_uk_U87 (.B2( u0_uk_K_r0_28 ) , .A2( u0_uk_K_r0_49 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n858 ) );
  OAI22_X1 u0_uk_U883 (.ZN( u0_K7_10 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n371 ) , .B2( u0_uk_n401 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U884 (.ZN( u0_K4_11 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n525 ) );
  OAI22_X1 u0_uk_U898 (.ZN( u0_K7_14 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n361 ) , .B2( u0_uk_n396 ) );
  OAI22_X1 u0_uk_U900 (.ZN( u0_K13_24 ) , .B2( u0_uk_n132 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n83 ) , .A2( u0_uk_n91 ) );
  OAI22_X1 u0_uk_U903 (.ZN( u0_K3_21 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n542 ) , .B2( u0_uk_n567 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U914 (.ZN( u0_K4_14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n510 ) , .B2( u0_uk_n536 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U915 (.ZN( u0_K3_13 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n564 ) , .B2( u0_uk_n569 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U916 (.ZN( u0_K4_36 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n208 ) , .A2( u0_uk_n507 ) , .B2( u0_uk_n512 ) );
  OAI22_X1 u0_uk_U918 (.ZN( u0_K6_30 ) , .A1( u0_uk_n203 ) , .A2( u0_uk_n445 ) , .B2( u0_uk_n450 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U923 (.ZN( u0_K6_42 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n413 ) , .B2( u0_uk_n420 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U924 (.ZN( u0_K6_39 ) , .A1( u0_uk_n162 ) , .B2( u0_uk_n428 ) , .A2( u0_uk_n447 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U928 (.ZN( u0_K2_39 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n607 ) , .A2( u0_uk_n622 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U929 (.ZN( u0_K13_23 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n121 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n91 ) );
  OAI22_X1 u0_uk_U933 (.ZN( u0_K11_16 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n190 ) , .B2( u0_uk_n196 ) );
  OAI22_X1 u0_uk_U942 (.ZN( u0_K11_24 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n201 ) , .B2( u0_uk_n206 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U957 (.ZN( u0_K13_8 ) , .A2( u0_uk_n101 ) , .B2( u0_uk_n107 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n147 ) );
  OAI22_X1 u0_uk_U959 (.ZN( u0_K11_18 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n215 ) , .B2( u0_uk_n221 ) );
  OAI22_X1 u0_uk_U965 (.ZN( u0_K6_36 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n439 ) , .A2( u0_uk_n447 ) );
  OAI22_X1 u0_uk_U968 (.ZN( u0_K2_38 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n593 ) , .B2( u0_uk_n612 ) );
  OAI22_X1 u0_uk_U970 (.ZN( u0_K2_37 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n594 ) , .A2( u0_uk_n621 ) );
  OAI22_X1 u0_uk_U975 (.ZN( u0_K11_45 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n204 ) , .B2( u0_uk_n211 ) , .B1( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U976 (.ZN( u0_K7_45 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n381 ) , .B2( u0_uk_n398 ) );
  OAI22_X1 u0_uk_U980 (.ZN( u0_K2_3 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n604 ) , .B2( u0_uk_n619 ) );
  OAI22_X1 u0_uk_U982 (.ZN( u0_K3_6 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n571 ) , .A2( u0_uk_n576 ) );
  OAI22_X1 u0_uk_U984 (.ZN( u0_K7_7 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n257 ) , .A2( u0_uk_n370 ) , .B2( u0_uk_n392 ) );
  OAI22_X1 u0_uk_U985 (.ZN( u0_K3_7 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n547 ) , .B2( u0_uk_n565 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U988 (.ZN( u0_K6_25 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n434 ) );
  NAND2_X1 u0_uk_U995 (.A1( u0_uk_K_r5_5 ) , .ZN( u0_uk_n778 ) , .A2( u0_uk_n93 ) );
  XOR2_X1 u1_U136 (.B( u1_L0_10 ) , .Z( u1_N41 ) , .A( u1_out1_10 ) );
  XOR2_X1 u1_U236 (.B( u1_L0_1 ) , .Z( u1_N32 ) , .A( u1_out1_1 ) );
  XOR2_X1 u1_U49 (.B( u1_L0_26 ) , .Z( u1_N57 ) , .A( u1_out1_26 ) );
  XOR2_X1 u1_U55 (.B( u1_L0_20 ) , .Z( u1_N51 ) , .A( u1_out1_20 ) );
  XOR2_X1 u1_u1_U33 (.B( u1_K2_24 ) , .A( u1_R0_17 ) , .Z( u1_u1_X_24 ) );
  XOR2_X1 u1_u1_U34 (.B( u1_K2_23 ) , .A( u1_R0_16 ) , .Z( u1_u1_X_23 ) );
  XOR2_X1 u1_u1_U35 (.B( u1_K2_22 ) , .A( u1_R0_15 ) , .Z( u1_u1_X_22 ) );
  XOR2_X1 u1_u1_U36 (.B( u1_K2_21 ) , .A( u1_R0_14 ) , .Z( u1_u1_X_21 ) );
  XOR2_X1 u1_u1_U37 (.B( u1_K2_20 ) , .A( u1_R0_13 ) , .Z( u1_u1_X_20 ) );
  XOR2_X1 u1_u1_U39 (.B( u1_K2_19 ) , .A( u1_R0_12 ) , .Z( u1_u1_X_19 ) );
  OAI22_X1 u1_u1_u3_U10 (.B1( u1_u1_u3_n113 ) , .A2( u1_u1_u3_n135 ) , .A1( u1_u1_u3_n150 ) , .B2( u1_u1_u3_n164 ) , .ZN( u1_u1_u3_n98 ) );
  OAI211_X1 u1_u1_u3_U11 (.B( u1_u1_u3_n106 ) , .ZN( u1_u1_u3_n119 ) , .C2( u1_u1_u3_n128 ) , .C1( u1_u1_u3_n167 ) , .A( u1_u1_u3_n181 ) );
  AOI221_X1 u1_u1_u3_U12 (.C1( u1_u1_u3_n105 ) , .ZN( u1_u1_u3_n106 ) , .A( u1_u1_u3_n131 ) , .B2( u1_u1_u3_n132 ) , .C2( u1_u1_u3_n133 ) , .B1( u1_u1_u3_n169 ) );
  INV_X1 u1_u1_u3_U13 (.ZN( u1_u1_u3_n181 ) , .A( u1_u1_u3_n98 ) );
  NAND2_X1 u1_u1_u3_U14 (.ZN( u1_u1_u3_n105 ) , .A2( u1_u1_u3_n130 ) , .A1( u1_u1_u3_n155 ) );
  AOI22_X1 u1_u1_u3_U15 (.B1( u1_u1_u3_n115 ) , .A2( u1_u1_u3_n116 ) , .ZN( u1_u1_u3_n123 ) , .B2( u1_u1_u3_n133 ) , .A1( u1_u1_u3_n169 ) );
  NAND2_X1 u1_u1_u3_U16 (.ZN( u1_u1_u3_n116 ) , .A2( u1_u1_u3_n151 ) , .A1( u1_u1_u3_n182 ) );
  NOR2_X1 u1_u1_u3_U17 (.ZN( u1_u1_u3_n126 ) , .A2( u1_u1_u3_n150 ) , .A1( u1_u1_u3_n164 ) );
  AOI21_X1 u1_u1_u3_U18 (.ZN( u1_u1_u3_n112 ) , .B2( u1_u1_u3_n146 ) , .B1( u1_u1_u3_n155 ) , .A( u1_u1_u3_n167 ) );
  NAND2_X1 u1_u1_u3_U19 (.A1( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n142 ) , .A2( u1_u1_u3_n164 ) );
  NAND2_X1 u1_u1_u3_U20 (.ZN( u1_u1_u3_n132 ) , .A2( u1_u1_u3_n152 ) , .A1( u1_u1_u3_n156 ) );
  AND2_X1 u1_u1_u3_U21 (.A2( u1_u1_u3_n113 ) , .A1( u1_u1_u3_n114 ) , .ZN( u1_u1_u3_n151 ) );
  INV_X1 u1_u1_u3_U22 (.A( u1_u1_u3_n133 ) , .ZN( u1_u1_u3_n165 ) );
  INV_X1 u1_u1_u3_U23 (.A( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n170 ) );
  NAND2_X1 u1_u1_u3_U24 (.A1( u1_u1_u3_n107 ) , .A2( u1_u1_u3_n108 ) , .ZN( u1_u1_u3_n140 ) );
  NAND2_X1 u1_u1_u3_U25 (.ZN( u1_u1_u3_n117 ) , .A1( u1_u1_u3_n124 ) , .A2( u1_u1_u3_n148 ) );
  NAND2_X1 u1_u1_u3_U26 (.ZN( u1_u1_u3_n143 ) , .A1( u1_u1_u3_n165 ) , .A2( u1_u1_u3_n167 ) );
  INV_X1 u1_u1_u3_U27 (.A( u1_u1_u3_n130 ) , .ZN( u1_u1_u3_n177 ) );
  INV_X1 u1_u1_u3_U28 (.A( u1_u1_u3_n128 ) , .ZN( u1_u1_u3_n176 ) );
  INV_X1 u1_u1_u3_U29 (.A( u1_u1_u3_n155 ) , .ZN( u1_u1_u3_n174 ) );
  INV_X1 u1_u1_u3_U3 (.A( u1_u1_u3_n129 ) , .ZN( u1_u1_u3_n183 ) );
  INV_X1 u1_u1_u3_U30 (.A( u1_u1_u3_n139 ) , .ZN( u1_u1_u3_n185 ) );
  NOR2_X1 u1_u1_u3_U31 (.ZN( u1_u1_u3_n135 ) , .A2( u1_u1_u3_n141 ) , .A1( u1_u1_u3_n169 ) );
  OAI222_X1 u1_u1_u3_U32 (.C2( u1_u1_u3_n107 ) , .A2( u1_u1_u3_n108 ) , .B1( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n138 ) , .B2( u1_u1_u3_n146 ) , .C1( u1_u1_u3_n154 ) , .A1( u1_u1_u3_n164 ) );
  NOR4_X1 u1_u1_u3_U33 (.A4( u1_u1_u3_n157 ) , .A3( u1_u1_u3_n158 ) , .A2( u1_u1_u3_n159 ) , .A1( u1_u1_u3_n160 ) , .ZN( u1_u1_u3_n161 ) );
  AOI21_X1 u1_u1_u3_U34 (.B2( u1_u1_u3_n152 ) , .B1( u1_u1_u3_n153 ) , .ZN( u1_u1_u3_n158 ) , .A( u1_u1_u3_n164 ) );
  AOI21_X1 u1_u1_u3_U35 (.A( u1_u1_u3_n154 ) , .B2( u1_u1_u3_n155 ) , .B1( u1_u1_u3_n156 ) , .ZN( u1_u1_u3_n157 ) );
  AOI21_X1 u1_u1_u3_U36 (.A( u1_u1_u3_n149 ) , .B2( u1_u1_u3_n150 ) , .B1( u1_u1_u3_n151 ) , .ZN( u1_u1_u3_n159 ) );
  AOI211_X1 u1_u1_u3_U37 (.ZN( u1_u1_u3_n109 ) , .A( u1_u1_u3_n119 ) , .C2( u1_u1_u3_n129 ) , .B( u1_u1_u3_n138 ) , .C1( u1_u1_u3_n141 ) );
  AOI211_X1 u1_u1_u3_U38 (.B( u1_u1_u3_n119 ) , .A( u1_u1_u3_n120 ) , .C2( u1_u1_u3_n121 ) , .ZN( u1_u1_u3_n122 ) , .C1( u1_u1_u3_n179 ) );
  INV_X1 u1_u1_u3_U39 (.A( u1_u1_u3_n156 ) , .ZN( u1_u1_u3_n179 ) );
  INV_X1 u1_u1_u3_U4 (.A( u1_u1_u3_n140 ) , .ZN( u1_u1_u3_n182 ) );
  OAI22_X1 u1_u1_u3_U40 (.B1( u1_u1_u3_n118 ) , .ZN( u1_u1_u3_n120 ) , .A1( u1_u1_u3_n135 ) , .B2( u1_u1_u3_n154 ) , .A2( u1_u1_u3_n178 ) );
  AND3_X1 u1_u1_u3_U41 (.ZN( u1_u1_u3_n118 ) , .A2( u1_u1_u3_n124 ) , .A1( u1_u1_u3_n144 ) , .A3( u1_u1_u3_n152 ) );
  INV_X1 u1_u1_u3_U42 (.A( u1_u1_u3_n121 ) , .ZN( u1_u1_u3_n164 ) );
  NAND2_X1 u1_u1_u3_U43 (.ZN( u1_u1_u3_n133 ) , .A1( u1_u1_u3_n154 ) , .A2( u1_u1_u3_n164 ) );
  OAI211_X1 u1_u1_u3_U44 (.B( u1_u1_u3_n127 ) , .ZN( u1_u1_u3_n139 ) , .C1( u1_u1_u3_n150 ) , .C2( u1_u1_u3_n154 ) , .A( u1_u1_u3_n184 ) );
  INV_X1 u1_u1_u3_U45 (.A( u1_u1_u3_n125 ) , .ZN( u1_u1_u3_n184 ) );
  AOI221_X1 u1_u1_u3_U46 (.A( u1_u1_u3_n126 ) , .ZN( u1_u1_u3_n127 ) , .C2( u1_u1_u3_n132 ) , .C1( u1_u1_u3_n169 ) , .B2( u1_u1_u3_n170 ) , .B1( u1_u1_u3_n174 ) );
  OAI22_X1 u1_u1_u3_U47 (.A1( u1_u1_u3_n124 ) , .ZN( u1_u1_u3_n125 ) , .B2( u1_u1_u3_n145 ) , .A2( u1_u1_u3_n165 ) , .B1( u1_u1_u3_n167 ) );
  NOR2_X1 u1_u1_u3_U48 (.A1( u1_u1_u3_n113 ) , .ZN( u1_u1_u3_n131 ) , .A2( u1_u1_u3_n154 ) );
  NAND2_X1 u1_u1_u3_U49 (.A1( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n150 ) , .A2( u1_u1_u3_n99 ) );
  INV_X1 u1_u1_u3_U5 (.A( u1_u1_u3_n117 ) , .ZN( u1_u1_u3_n178 ) );
  NAND2_X1 u1_u1_u3_U50 (.A2( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n155 ) , .A1( u1_u1_u3_n97 ) );
  INV_X1 u1_u1_u3_U51 (.A( u1_u1_u3_n141 ) , .ZN( u1_u1_u3_n167 ) );
  AOI21_X1 u1_u1_u3_U52 (.B2( u1_u1_u3_n114 ) , .B1( u1_u1_u3_n146 ) , .A( u1_u1_u3_n154 ) , .ZN( u1_u1_u3_n94 ) );
  AOI21_X1 u1_u1_u3_U53 (.ZN( u1_u1_u3_n110 ) , .B2( u1_u1_u3_n142 ) , .B1( u1_u1_u3_n186 ) , .A( u1_u1_u3_n95 ) );
  INV_X1 u1_u1_u3_U54 (.A( u1_u1_u3_n145 ) , .ZN( u1_u1_u3_n186 ) );
  AOI21_X1 u1_u1_u3_U55 (.B1( u1_u1_u3_n124 ) , .A( u1_u1_u3_n149 ) , .B2( u1_u1_u3_n155 ) , .ZN( u1_u1_u3_n95 ) );
  INV_X1 u1_u1_u3_U56 (.A( u1_u1_u3_n149 ) , .ZN( u1_u1_u3_n169 ) );
  NAND2_X1 u1_u1_u3_U57 (.ZN( u1_u1_u3_n124 ) , .A1( u1_u1_u3_n96 ) , .A2( u1_u1_u3_n97 ) );
  NAND2_X1 u1_u1_u3_U58 (.A2( u1_u1_u3_n100 ) , .ZN( u1_u1_u3_n146 ) , .A1( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U59 (.A1( u1_u1_u3_n101 ) , .ZN( u1_u1_u3_n145 ) , .A2( u1_u1_u3_n99 ) );
  AOI221_X1 u1_u1_u3_U6 (.A( u1_u1_u3_n131 ) , .C2( u1_u1_u3_n132 ) , .C1( u1_u1_u3_n133 ) , .ZN( u1_u1_u3_n134 ) , .B1( u1_u1_u3_n143 ) , .B2( u1_u1_u3_n177 ) );
  NAND2_X1 u1_u1_u3_U60 (.A1( u1_u1_u3_n100 ) , .ZN( u1_u1_u3_n156 ) , .A2( u1_u1_u3_n99 ) );
  NAND2_X1 u1_u1_u3_U61 (.A2( u1_u1_u3_n101 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n148 ) );
  NAND2_X1 u1_u1_u3_U62 (.A1( u1_u1_u3_n100 ) , .A2( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n128 ) );
  NAND2_X1 u1_u1_u3_U63 (.A2( u1_u1_u3_n101 ) , .A1( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n152 ) );
  NAND2_X1 u1_u1_u3_U64 (.A2( u1_u1_u3_n101 ) , .ZN( u1_u1_u3_n114 ) , .A1( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U65 (.ZN( u1_u1_u3_n107 ) , .A1( u1_u1_u3_n97 ) , .A2( u1_u1_u3_n99 ) );
  NAND2_X1 u1_u1_u3_U66 (.A2( u1_u1_u3_n100 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n113 ) );
  NAND2_X1 u1_u1_u3_U67 (.A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n153 ) , .A2( u1_u1_u3_n97 ) );
  NAND2_X1 u1_u1_u3_U68 (.A2( u1_u1_u3_n103 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n130 ) );
  NAND2_X1 u1_u1_u3_U69 (.A2( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n144 ) , .A1( u1_u1_u3_n96 ) );
  OAI22_X1 u1_u1_u3_U7 (.B2( u1_u1_u3_n147 ) , .A2( u1_u1_u3_n148 ) , .ZN( u1_u1_u3_n160 ) , .B1( u1_u1_u3_n165 ) , .A1( u1_u1_u3_n168 ) );
  NAND2_X1 u1_u1_u3_U70 (.A1( u1_u1_u3_n102 ) , .A2( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n108 ) );
  NOR2_X1 u1_u1_u3_U71 (.A2( u1_u1_X_19 ) , .A1( u1_u1_X_20 ) , .ZN( u1_u1_u3_n99 ) );
  NOR2_X1 u1_u1_u3_U72 (.A2( u1_u1_X_21 ) , .A1( u1_u1_X_24 ) , .ZN( u1_u1_u3_n103 ) );
  NOR2_X1 u1_u1_u3_U73 (.A2( u1_u1_X_24 ) , .A1( u1_u1_u3_n171 ) , .ZN( u1_u1_u3_n97 ) );
  NOR2_X1 u1_u1_u3_U74 (.A2( u1_u1_X_23 ) , .ZN( u1_u1_u3_n141 ) , .A1( u1_u1_u3_n166 ) );
  NOR2_X1 u1_u1_u3_U75 (.A2( u1_u1_X_19 ) , .A1( u1_u1_u3_n172 ) , .ZN( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U76 (.A1( u1_u1_X_22 ) , .A2( u1_u1_X_23 ) , .ZN( u1_u1_u3_n154 ) );
  NAND2_X1 u1_u1_u3_U77 (.A1( u1_u1_X_23 ) , .ZN( u1_u1_u3_n149 ) , .A2( u1_u1_u3_n166 ) );
  NOR2_X1 u1_u1_u3_U78 (.A2( u1_u1_X_22 ) , .A1( u1_u1_X_23 ) , .ZN( u1_u1_u3_n121 ) );
  AND2_X1 u1_u1_u3_U79 (.A1( u1_u1_X_24 ) , .ZN( u1_u1_u3_n101 ) , .A2( u1_u1_u3_n171 ) );
  AND3_X1 u1_u1_u3_U8 (.A3( u1_u1_u3_n144 ) , .A2( u1_u1_u3_n145 ) , .A1( u1_u1_u3_n146 ) , .ZN( u1_u1_u3_n147 ) );
  AND2_X1 u1_u1_u3_U80 (.A1( u1_u1_X_19 ) , .ZN( u1_u1_u3_n102 ) , .A2( u1_u1_u3_n172 ) );
  AND2_X1 u1_u1_u3_U81 (.A1( u1_u1_X_21 ) , .A2( u1_u1_X_24 ) , .ZN( u1_u1_u3_n100 ) );
  AND2_X1 u1_u1_u3_U82 (.A2( u1_u1_X_19 ) , .A1( u1_u1_X_20 ) , .ZN( u1_u1_u3_n104 ) );
  INV_X1 u1_u1_u3_U83 (.A( u1_u1_X_22 ) , .ZN( u1_u1_u3_n166 ) );
  INV_X1 u1_u1_u3_U84 (.A( u1_u1_X_21 ) , .ZN( u1_u1_u3_n171 ) );
  INV_X1 u1_u1_u3_U85 (.A( u1_u1_X_20 ) , .ZN( u1_u1_u3_n172 ) );
  OR4_X1 u1_u1_u3_U86 (.ZN( u1_out1_10 ) , .A4( u1_u1_u3_n136 ) , .A3( u1_u1_u3_n137 ) , .A1( u1_u1_u3_n138 ) , .A2( u1_u1_u3_n139 ) );
  OAI222_X1 u1_u1_u3_U87 (.C1( u1_u1_u3_n128 ) , .ZN( u1_u1_u3_n137 ) , .B1( u1_u1_u3_n148 ) , .A2( u1_u1_u3_n150 ) , .B2( u1_u1_u3_n154 ) , .C2( u1_u1_u3_n164 ) , .A1( u1_u1_u3_n167 ) );
  OAI221_X1 u1_u1_u3_U88 (.A( u1_u1_u3_n134 ) , .B2( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n136 ) , .C1( u1_u1_u3_n149 ) , .B1( u1_u1_u3_n151 ) , .C2( u1_u1_u3_n183 ) );
  NAND4_X1 u1_u1_u3_U89 (.ZN( u1_out1_26 ) , .A4( u1_u1_u3_n109 ) , .A3( u1_u1_u3_n110 ) , .A2( u1_u1_u3_n111 ) , .A1( u1_u1_u3_n173 ) );
  INV_X1 u1_u1_u3_U9 (.A( u1_u1_u3_n143 ) , .ZN( u1_u1_u3_n168 ) );
  INV_X1 u1_u1_u3_U90 (.ZN( u1_u1_u3_n173 ) , .A( u1_u1_u3_n94 ) );
  OAI21_X1 u1_u1_u3_U91 (.ZN( u1_u1_u3_n111 ) , .B2( u1_u1_u3_n117 ) , .A( u1_u1_u3_n133 ) , .B1( u1_u1_u3_n176 ) );
  NAND4_X1 u1_u1_u3_U92 (.ZN( u1_out1_20 ) , .A4( u1_u1_u3_n122 ) , .A3( u1_u1_u3_n123 ) , .A1( u1_u1_u3_n175 ) , .A2( u1_u1_u3_n180 ) );
  INV_X1 u1_u1_u3_U93 (.A( u1_u1_u3_n112 ) , .ZN( u1_u1_u3_n175 ) );
  INV_X1 u1_u1_u3_U94 (.A( u1_u1_u3_n126 ) , .ZN( u1_u1_u3_n180 ) );
  NAND4_X1 u1_u1_u3_U95 (.ZN( u1_out1_1 ) , .A4( u1_u1_u3_n161 ) , .A3( u1_u1_u3_n162 ) , .A2( u1_u1_u3_n163 ) , .A1( u1_u1_u3_n185 ) );
  NAND2_X1 u1_u1_u3_U96 (.ZN( u1_u1_u3_n163 ) , .A2( u1_u1_u3_n170 ) , .A1( u1_u1_u3_n176 ) );
  AOI22_X1 u1_u1_u3_U97 (.B2( u1_u1_u3_n140 ) , .B1( u1_u1_u3_n141 ) , .A2( u1_u1_u3_n142 ) , .ZN( u1_u1_u3_n162 ) , .A1( u1_u1_u3_n177 ) );
  NAND3_X1 u1_u1_u3_U98 (.A1( u1_u1_u3_n114 ) , .ZN( u1_u1_u3_n115 ) , .A2( u1_u1_u3_n145 ) , .A3( u1_u1_u3_n153 ) );
  NAND3_X1 u1_u1_u3_U99 (.ZN( u1_u1_u3_n129 ) , .A2( u1_u1_u3_n144 ) , .A1( u1_u1_u3_n153 ) , .A3( u1_u1_u3_n182 ) );
  INV_X1 u1_uk_U169 (.ZN( u1_K2_19 ) , .A( u1_uk_n1025 ) );
  AOI22_X1 u1_uk_U170 (.B2( u1_uk_K_r0_11 ) , .A2( u1_uk_K_r0_47 ) , .ZN( u1_uk_n1025 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U770 (.ZN( u1_K2_21 ) , .A2( u1_uk_n1264 ) , .B2( u1_uk_n1268 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U906 (.ZN( u1_K2_24 ) , .A2( u1_uk_n1264 ) , .B2( u1_uk_n1279 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U94 (.ZN( u1_K2_23 ) , .B2( u1_uk_n1278 ) , .A2( u1_uk_n1299 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U940 (.ZN( u1_K2_20 ) , .A2( u1_uk_n1263 ) , .B2( u1_uk_n1292 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U973 (.ZN( u1_K2_22 ) , .B2( u1_uk_n1273 ) , .A2( u1_uk_n1290 ) , .B1( u1_uk_n222 ) , .A1( u1_uk_n31 ) );
  XOR2_X1 u2_U103 (.B( u2_L0_13 ) , .Z( u2_N44 ) , .A( u2_out1_13 ) );
  XOR2_X1 u2_U147 (.B( u2_L0_9 ) , .Z( u2_N40 ) , .A( u2_out1_9 ) );
  XOR2_X1 u2_U166 (.B( u2_L10_32 ) , .Z( u2_N383 ) , .A( u2_out11_32 ) );
  XOR2_X1 u2_U169 (.B( u2_L10_29 ) , .Z( u2_N380 ) , .A( u2_out11_29 ) );
  XOR2_X1 u2_U172 (.B( u2_L10_27 ) , .Z( u2_N378 ) , .A( u2_out11_27 ) );
  XOR2_X1 u2_U174 (.B( u2_L10_25 ) , .Z( u2_N376 ) , .A( u2_out11_25 ) );
  XOR2_X1 u2_U177 (.B( u2_L10_22 ) , .Z( u2_N373 ) , .A( u2_out11_22 ) );
  XOR2_X1 u2_U178 (.B( u2_L10_21 ) , .Z( u2_N372 ) , .A( u2_out11_21 ) );
  XOR2_X1 u2_U180 (.B( u2_L10_19 ) , .Z( u2_N370 ) , .A( u2_out11_19 ) );
  XOR2_X1 u2_U185 (.B( u2_L10_15 ) , .Z( u2_N366 ) , .A( u2_out11_15 ) );
  XOR2_X1 u2_U186 (.B( u2_L10_14 ) , .Z( u2_N365 ) , .A( u2_out11_14 ) );
  XOR2_X1 u2_U188 (.B( u2_L10_12 ) , .Z( u2_N363 ) , .A( u2_out11_12 ) );
  XOR2_X1 u2_U189 (.B( u2_L10_11 ) , .Z( u2_N362 ) , .A( u2_out11_11 ) );
  XOR2_X1 u2_U193 (.B( u2_L10_8 ) , .Z( u2_N359 ) , .A( u2_out11_8 ) );
  XOR2_X1 u2_U194 (.B( u2_L10_7 ) , .Z( u2_N358 ) , .A( u2_out11_7 ) );
  XOR2_X1 u2_U196 (.B( u2_L10_5 ) , .Z( u2_N356 ) , .A( u2_out11_5 ) );
  XOR2_X1 u2_U197 (.B( u2_L10_4 ) , .Z( u2_N355 ) , .A( u2_out11_4 ) );
  XOR2_X1 u2_U198 (.B( u2_L10_3 ) , .Z( u2_N354 ) , .A( u2_out11_3 ) );
  XOR2_X1 u2_U201 (.B( u2_L9_32 ) , .Z( u2_N351 ) , .A( u2_out10_32 ) );
  XOR2_X1 u2_U205 (.B( u2_L9_29 ) , .Z( u2_N348 ) , .A( u2_out10_29 ) );
  XOR2_X1 u2_U212 (.B( u2_L9_22 ) , .Z( u2_N341 ) , .A( u2_out10_22 ) );
  XOR2_X1 u2_U216 (.B( u2_L9_19 ) , .Z( u2_N338 ) , .A( u2_out10_19 ) );
  XOR2_X1 u2_U223 (.B( u2_L9_12 ) , .Z( u2_N331 ) , .A( u2_out10_12 ) );
  XOR2_X1 u2_U224 (.B( u2_L9_11 ) , .Z( u2_N330 ) , .A( u2_out10_11 ) );
  XOR2_X1 u2_U225 (.B( u2_L0_2 ) , .Z( u2_N33 ) , .A( u2_out1_2 ) );
  XOR2_X1 u2_U229 (.B( u2_L9_7 ) , .Z( u2_N326 ) , .A( u2_out10_7 ) );
  XOR2_X1 u2_U232 (.B( u2_L9_4 ) , .Z( u2_N323 ) , .A( u2_out10_4 ) );
  XOR2_X1 u2_U239 (.B( u2_L8_30 ) , .Z( u2_N317 ) , .A( u2_out9_30 ) );
  XOR2_X1 u2_U24 (.Z( u2_N8 ) , .B( u2_desIn_r_4 ) , .A( u2_out0_9 ) );
  XOR2_X1 u2_U241 (.B( u2_L8_28 ) , .Z( u2_N315 ) , .A( u2_out9_28 ) );
  XOR2_X1 u2_U245 (.B( u2_L8_24 ) , .Z( u2_N311 ) , .A( u2_out9_24 ) );
  XOR2_X1 u2_U252 (.B( u2_L8_18 ) , .Z( u2_N305 ) , .A( u2_out9_18 ) );
  XOR2_X1 u2_U254 (.B( u2_L8_16 ) , .Z( u2_N303 ) , .A( u2_out9_16 ) );
  XOR2_X1 u2_U257 (.B( u2_L8_13 ) , .Z( u2_N300 ) , .A( u2_out9_13 ) );
  XOR2_X1 u2_U258 (.Z( u2_N30 ) , .B( u2_desIn_r_48 ) , .A( u2_out0_31 ) );
  XOR2_X1 u2_U266 (.B( u2_L8_6 ) , .Z( u2_N293 ) , .A( u2_out9_6 ) );
  XOR2_X1 u2_U270 (.Z( u2_N29 ) , .B( u2_desIn_r_40 ) , .A( u2_out0_30 ) );
  XOR2_X1 u2_U271 (.B( u2_L8_2 ) , .Z( u2_N289 ) , .A( u2_out9_2 ) );
  XOR2_X1 u2_U292 (.Z( u2_N27 ) , .B( u2_desIn_r_24 ) , .A( u2_out0_28 ) );
  XOR2_X1 u2_U336 (.Z( u2_N23 ) , .B( u2_desIn_r_58 ) , .A( u2_out0_24 ) );
  XOR2_X1 u2_U344 (.B( u2_L5_31 ) , .Z( u2_N222 ) , .A( u2_out6_31 ) );
  XOR2_X1 u2_U345 (.B( u2_L5_30 ) , .Z( u2_N221 ) , .A( u2_out6_30 ) );
  XOR2_X1 u2_U347 (.Z( u2_N22 ) , .B( u2_desIn_r_50 ) , .A( u2_out0_23 ) );
  XOR2_X1 u2_U348 (.B( u2_L5_28 ) , .Z( u2_N219 ) , .A( u2_out6_28 ) );
  XOR2_X1 u2_U352 (.B( u2_L5_24 ) , .Z( u2_N215 ) , .A( u2_out6_24 ) );
  XOR2_X1 u2_U353 (.B( u2_L5_23 ) , .Z( u2_N214 ) , .A( u2_out6_23 ) );
  XOR2_X1 u2_U359 (.B( u2_L5_18 ) , .Z( u2_N209 ) , .A( u2_out6_18 ) );
  XOR2_X1 u2_U360 (.B( u2_L5_17 ) , .Z( u2_N208 ) , .A( u2_out6_17 ) );
  XOR2_X1 u2_U361 (.B( u2_L5_16 ) , .Z( u2_N207 ) , .A( u2_out6_16 ) );
  XOR2_X1 u2_U364 (.B( u2_L5_13 ) , .Z( u2_N204 ) , .A( u2_out6_13 ) );
  XOR2_X1 u2_U368 (.B( u2_L5_9 ) , .Z( u2_N200 ) , .A( u2_out6_9 ) );
  XOR2_X1 u2_U373 (.B( u2_L5_6 ) , .Z( u2_N197 ) , .A( u2_out6_6 ) );
  XOR2_X1 u2_U377 (.B( u2_L5_2 ) , .Z( u2_N193 ) , .A( u2_out6_2 ) );
  XOR2_X1 u2_U379 (.B( u2_L4_32 ) , .Z( u2_N191 ) , .A( u2_out5_32 ) );
  XOR2_X1 u2_U382 (.B( u2_L4_30 ) , .Z( u2_N189 ) , .A( u2_out5_30 ) );
  XOR2_X1 u2_U383 (.B( u2_L4_29 ) , .Z( u2_N188 ) , .A( u2_out5_29 ) );
  XOR2_X1 u2_U386 (.B( u2_L4_26 ) , .Z( u2_N185 ) , .A( u2_out5_26 ) );
  XOR2_X1 u2_U388 (.B( u2_L4_24 ) , .Z( u2_N183 ) , .A( u2_out5_24 ) );
  XOR2_X1 u2_U390 (.B( u2_L4_22 ) , .Z( u2_N181 ) , .A( u2_out5_22 ) );
  XOR2_X1 u2_U393 (.B( u2_L4_20 ) , .Z( u2_N179 ) , .A( u2_out5_20 ) );
  XOR2_X1 u2_U394 (.B( u2_L4_19 ) , .Z( u2_N178 ) , .A( u2_out5_19 ) );
  XOR2_X1 u2_U397 (.B( u2_L4_16 ) , .Z( u2_N175 ) , .A( u2_out5_16 ) );
  XOR2_X1 u2_U401 (.B( u2_L4_12 ) , .Z( u2_N171 ) , .A( u2_out5_12 ) );
  XOR2_X1 u2_U402 (.B( u2_L4_11 ) , .Z( u2_N170 ) , .A( u2_out5_11 ) );
  XOR2_X1 u2_U403 (.Z( u2_N17 ) , .B( u2_desIn_r_10 ) , .A( u2_out0_18 ) );
  XOR2_X1 u2_U404 (.B( u2_L4_10 ) , .Z( u2_N169 ) , .A( u2_out5_10 ) );
  XOR2_X1 u2_U407 (.B( u2_L4_7 ) , .Z( u2_N166 ) , .A( u2_out5_7 ) );
  XOR2_X1 u2_U408 (.B( u2_L4_6 ) , .Z( u2_N165 ) , .A( u2_out5_6 ) );
  XOR2_X1 u2_U410 (.B( u2_L4_4 ) , .Z( u2_N163 ) , .A( u2_out5_4 ) );
  XOR2_X1 u2_U413 (.B( u2_L4_1 ) , .Z( u2_N160 ) , .A( u2_out5_1 ) );
  XOR2_X1 u2_U414 (.Z( u2_N16 ) , .B( u2_desIn_r_2 ) , .A( u2_out0_17 ) );
  XOR2_X1 u2_U425 (.Z( u2_N15 ) , .B( u2_desIn_r_60 ) , .A( u2_out0_16 ) );
  XOR2_X1 u2_U43 (.B( u2_L0_31 ) , .Z( u2_N62 ) , .A( u2_out1_31 ) );
  XOR2_X1 u2_U458 (.Z( u2_N12 ) , .B( u2_desIn_r_36 ) , .A( u2_out0_13 ) );
  XOR2_X1 u2_U47 (.B( u2_L0_28 ) , .Z( u2_N59 ) , .A( u2_out1_28 ) );
  XOR2_X1 u2_U481 (.Z( u2_N1 ) , .B( u2_desIn_r_14 ) , .A( u2_out0_2 ) );
  XOR2_X1 u2_U483 (.Z( u2_FP_9 ) , .B( u2_L14_9 ) , .A( u2_out15_9 ) );
  XOR2_X1 u2_U486 (.Z( u2_FP_6 ) , .B( u2_L14_6 ) , .A( u2_out15_6 ) );
  XOR2_X1 u2_U491 (.Z( u2_FP_31 ) , .B( u2_L14_31 ) , .A( u2_out15_31 ) );
  XOR2_X1 u2_U492 (.Z( u2_FP_30 ) , .B( u2_L14_30 ) , .A( u2_out15_30 ) );
  XOR2_X1 u2_U493 (.Z( u2_FP_2 ) , .B( u2_L14_2 ) , .A( u2_out15_2 ) );
  XOR2_X1 u2_U495 (.Z( u2_FP_28 ) , .B( u2_L14_28 ) , .A( u2_out15_28 ) );
  XOR2_X1 u2_U497 (.Z( u2_FP_26 ) , .B( u2_L14_26 ) , .A( u2_out15_26 ) );
  XOR2_X1 u2_U499 (.Z( u2_FP_24 ) , .B( u2_L14_24 ) , .A( u2_out15_24 ) );
  XOR2_X1 u2_U500 (.Z( u2_FP_23 ) , .B( u2_L14_23 ) , .A( u2_out15_23 ) );
  XOR2_X1 u2_U503 (.Z( u2_FP_20 ) , .B( u2_L14_20 ) , .A( u2_out15_20 ) );
  XOR2_X1 u2_U504 (.Z( u2_FP_1 ) , .B( u2_L14_1 ) , .A( u2_out15_1 ) );
  XOR2_X1 u2_U506 (.Z( u2_FP_18 ) , .B( u2_L14_18 ) , .A( u2_out15_18 ) );
  XOR2_X1 u2_U507 (.Z( u2_FP_17 ) , .B( u2_L14_17 ) , .A( u2_out15_17 ) );
  XOR2_X1 u2_U508 (.Z( u2_FP_16 ) , .B( u2_L14_16 ) , .A( u2_out15_16 ) );
  XOR2_X1 u2_U511 (.Z( u2_FP_13 ) , .B( u2_L14_13 ) , .A( u2_out15_13 ) );
  XOR2_X1 u2_U514 (.Z( u2_FP_10 ) , .B( u2_L14_10 ) , .A( u2_out15_10 ) );
  XOR2_X1 u2_U52 (.B( u2_L0_23 ) , .Z( u2_N54 ) , .A( u2_out1_23 ) );
  XOR2_X1 u2_U57 (.Z( u2_N5 ) , .B( u2_desIn_r_46 ) , .A( u2_out0_6 ) );
  XOR2_X1 u2_U58 (.B( u2_L0_18 ) , .Z( u2_N49 ) , .A( u2_out1_18 ) );
  XOR2_X1 u2_U59 (.B( u2_L0_17 ) , .Z( u2_N48 ) , .A( u2_out1_17 ) );
  XOR2_X1 u2_U61 (.B( u2_L13_31 ) , .Z( u2_N478 ) , .A( u2_out14_31 ) );
  XOR2_X1 u2_U62 (.B( u2_L13_30 ) , .Z( u2_N477 ) , .A( u2_out14_30 ) );
  XOR2_X1 u2_U64 (.B( u2_L13_28 ) , .Z( u2_N475 ) , .A( u2_out14_28 ) );
  XOR2_X1 u2_U66 (.B( u2_L13_26 ) , .Z( u2_N473 ) , .A( u2_out14_26 ) );
  XOR2_X1 u2_U68 (.B( u2_L13_24 ) , .Z( u2_N471 ) , .A( u2_out14_24 ) );
  XOR2_X1 u2_U69 (.B( u2_L13_23 ) , .Z( u2_N470 ) , .A( u2_out14_23 ) );
  XOR2_X1 u2_U73 (.B( u2_L13_20 ) , .Z( u2_N467 ) , .A( u2_out14_20 ) );
  XOR2_X1 u2_U75 (.B( u2_L13_18 ) , .Z( u2_N465 ) , .A( u2_out14_18 ) );
  XOR2_X1 u2_U76 (.B( u2_L13_17 ) , .Z( u2_N464 ) , .A( u2_out14_17 ) );
  XOR2_X1 u2_U77 (.B( u2_L13_16 ) , .Z( u2_N463 ) , .A( u2_out14_16 ) );
  XOR2_X1 u2_U80 (.B( u2_L13_13 ) , .Z( u2_N460 ) , .A( u2_out14_13 ) );
  XOR2_X1 u2_U84 (.B( u2_L13_10 ) , .Z( u2_N457 ) , .A( u2_out14_10 ) );
  XOR2_X1 u2_U85 (.B( u2_L13_9 ) , .Z( u2_N456 ) , .A( u2_out14_9 ) );
  XOR2_X1 u2_U88 (.B( u2_L13_6 ) , .Z( u2_N453 ) , .A( u2_out14_6 ) );
  XOR2_X1 u2_U93 (.B( u2_L13_2 ) , .Z( u2_N449 ) , .A( u2_out14_2 ) );
  XOR2_X1 u2_U94 (.B( u2_L13_1 ) , .Z( u2_N448 ) , .A( u2_out14_1 ) );
  XOR2_X1 u2_u0_U1 (.B( u2_K1_9 ) , .A( u2_desIn_r_47 ) , .Z( u2_u0_X_9 ) );
  XOR2_X1 u2_u0_U16 (.B( u2_K1_3 ) , .A( u2_desIn_r_15 ) , .Z( u2_u0_X_3 ) );
  XOR2_X1 u2_u0_U2 (.B( u2_K1_8 ) , .A( u2_desIn_r_39 ) , .Z( u2_u0_X_8 ) );
  XOR2_X1 u2_u0_U27 (.B( u2_K1_2 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_2 ) );
  XOR2_X1 u2_u0_U3 (.B( u2_K1_7 ) , .A( u2_desIn_r_31 ) , .Z( u2_u0_X_7 ) );
  XOR2_X1 u2_u0_U4 (.B( u2_K1_6 ) , .A( u2_desIn_r_39 ) , .Z( u2_u0_X_6 ) );
  XOR2_X1 u2_u0_U40 (.B( u2_K1_18 ) , .A( u2_desIn_r_37 ) , .Z( u2_u0_X_18 ) );
  XOR2_X1 u2_u0_U41 (.B( u2_K1_17 ) , .A( u2_desIn_r_29 ) , .Z( u2_u0_X_17 ) );
  XOR2_X1 u2_u0_U42 (.B( u2_K1_16 ) , .A( u2_desIn_r_21 ) , .Z( u2_u0_X_16 ) );
  XOR2_X1 u2_u0_U43 (.B( u2_K1_15 ) , .A( u2_desIn_r_13 ) , .Z( u2_u0_X_15 ) );
  XOR2_X1 u2_u0_U44 (.B( u2_K1_14 ) , .A( u2_desIn_r_5 ) , .Z( u2_u0_X_14 ) );
  XOR2_X1 u2_u0_U45 (.B( u2_K1_13 ) , .A( u2_desIn_r_63 ) , .Z( u2_u0_X_13 ) );
  XOR2_X1 u2_u0_U46 (.B( u2_K1_12 ) , .A( u2_desIn_r_5 ) , .Z( u2_u0_X_12 ) );
  XOR2_X1 u2_u0_U47 (.B( u2_K1_11 ) , .A( u2_desIn_r_63 ) , .Z( u2_u0_X_11 ) );
  XOR2_X1 u2_u0_U48 (.B( u2_K1_10 ) , .A( u2_desIn_r_55 ) , .Z( u2_u0_X_10 ) );
  XOR2_X1 u2_u0_U5 (.B( u2_K1_5 ) , .A( u2_desIn_r_31 ) , .Z( u2_u0_X_5 ) );
  XOR2_X1 u2_u0_U6 (.B( u2_K1_4 ) , .A( u2_desIn_r_23 ) , .Z( u2_u0_X_4 ) );
  AND3_X1 u2_u0_u0_U10 (.A2( u2_u0_u0_n112 ) , .ZN( u2_u0_u0_n127 ) , .A3( u2_u0_u0_n130 ) , .A1( u2_u0_u0_n148 ) );
  NAND2_X1 u2_u0_u0_U11 (.ZN( u2_u0_u0_n113 ) , .A1( u2_u0_u0_n139 ) , .A2( u2_u0_u0_n149 ) );
  AND2_X1 u2_u0_u0_U12 (.ZN( u2_u0_u0_n107 ) , .A1( u2_u0_u0_n130 ) , .A2( u2_u0_u0_n140 ) );
  AND2_X1 u2_u0_u0_U13 (.A2( u2_u0_u0_n129 ) , .A1( u2_u0_u0_n130 ) , .ZN( u2_u0_u0_n151 ) );
  AND2_X1 u2_u0_u0_U14 (.A1( u2_u0_u0_n108 ) , .A2( u2_u0_u0_n125 ) , .ZN( u2_u0_u0_n145 ) );
  INV_X1 u2_u0_u0_U15 (.A( u2_u0_u0_n143 ) , .ZN( u2_u0_u0_n173 ) );
  NOR2_X1 u2_u0_u0_U16 (.A2( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n147 ) , .A1( u2_u0_u0_n160 ) );
  OAI22_X1 u2_u0_u0_U17 (.B1( u2_u0_u0_n125 ) , .ZN( u2_u0_u0_n126 ) , .A1( u2_u0_u0_n138 ) , .A2( u2_u0_u0_n146 ) , .B2( u2_u0_u0_n147 ) );
  OAI22_X1 u2_u0_u0_U18 (.B1( u2_u0_u0_n131 ) , .A1( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n147 ) , .A2( u2_u0_u0_n90 ) , .ZN( u2_u0_u0_n91 ) );
  AND3_X1 u2_u0_u0_U19 (.A3( u2_u0_u0_n121 ) , .A2( u2_u0_u0_n125 ) , .A1( u2_u0_u0_n148 ) , .ZN( u2_u0_u0_n90 ) );
  NOR2_X1 u2_u0_u0_U20 (.A1( u2_u0_u0_n163 ) , .A2( u2_u0_u0_n164 ) , .ZN( u2_u0_u0_n95 ) );
  AOI22_X1 u2_u0_u0_U21 (.B2( u2_u0_u0_n109 ) , .A2( u2_u0_u0_n110 ) , .ZN( u2_u0_u0_n111 ) , .B1( u2_u0_u0_n118 ) , .A1( u2_u0_u0_n160 ) );
  NAND2_X1 u2_u0_u0_U22 (.A1( u2_u0_u0_n100 ) , .A2( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n125 ) );
  NAND2_X1 u2_u0_u0_U23 (.A1( u2_u0_u0_n101 ) , .A2( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n150 ) );
  INV_X1 u2_u0_u0_U24 (.A( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n161 ) );
  INV_X1 u2_u0_u0_U25 (.A( u2_u0_u0_n118 ) , .ZN( u2_u0_u0_n158 ) );
  AOI21_X1 u2_u0_u0_U26 (.B1( u2_u0_u0_n127 ) , .B2( u2_u0_u0_n129 ) , .A( u2_u0_u0_n138 ) , .ZN( u2_u0_u0_n96 ) );
  AOI21_X1 u2_u0_u0_U27 (.ZN( u2_u0_u0_n104 ) , .B1( u2_u0_u0_n107 ) , .B2( u2_u0_u0_n141 ) , .A( u2_u0_u0_n144 ) );
  NAND2_X1 u2_u0_u0_U28 (.A2( u2_u0_u0_n100 ) , .A1( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n139 ) );
  NAND2_X1 u2_u0_u0_U29 (.A2( u2_u0_u0_n100 ) , .ZN( u2_u0_u0_n131 ) , .A1( u2_u0_u0_n92 ) );
  INV_X1 u2_u0_u0_U3 (.A( u2_u0_u0_n113 ) , .ZN( u2_u0_u0_n166 ) );
  NAND2_X1 u2_u0_u0_U30 (.A2( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n114 ) , .A1( u2_u0_u0_n92 ) );
  NOR2_X1 u2_u0_u0_U31 (.A1( u2_u0_u0_n120 ) , .ZN( u2_u0_u0_n143 ) , .A2( u2_u0_u0_n167 ) );
  OAI221_X1 u2_u0_u0_U32 (.C1( u2_u0_u0_n112 ) , .ZN( u2_u0_u0_n120 ) , .B1( u2_u0_u0_n138 ) , .B2( u2_u0_u0_n141 ) , .C2( u2_u0_u0_n147 ) , .A( u2_u0_u0_n172 ) );
  AOI211_X1 u2_u0_u0_U33 (.B( u2_u0_u0_n115 ) , .A( u2_u0_u0_n116 ) , .C2( u2_u0_u0_n117 ) , .C1( u2_u0_u0_n118 ) , .ZN( u2_u0_u0_n119 ) );
  INV_X1 u2_u0_u0_U34 (.A( u2_u0_u0_n138 ) , .ZN( u2_u0_u0_n160 ) );
  NAND2_X1 u2_u0_u0_U35 (.A2( u2_u0_u0_n102 ) , .A1( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n149 ) );
  NAND2_X1 u2_u0_u0_U36 (.A2( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n121 ) , .A1( u2_u0_u0_n93 ) );
  NAND2_X1 u2_u0_u0_U37 (.ZN( u2_u0_u0_n112 ) , .A2( u2_u0_u0_n92 ) , .A1( u2_u0_u0_n93 ) );
  INV_X1 u2_u0_u0_U38 (.ZN( u2_u0_u0_n172 ) , .A( u2_u0_u0_n88 ) );
  OAI222_X1 u2_u0_u0_U39 (.C1( u2_u0_u0_n108 ) , .A1( u2_u0_u0_n125 ) , .B2( u2_u0_u0_n128 ) , .B1( u2_u0_u0_n144 ) , .A2( u2_u0_u0_n158 ) , .C2( u2_u0_u0_n161 ) , .ZN( u2_u0_u0_n88 ) );
  AOI21_X1 u2_u0_u0_U4 (.B1( u2_u0_u0_n114 ) , .ZN( u2_u0_u0_n115 ) , .B2( u2_u0_u0_n129 ) , .A( u2_u0_u0_n161 ) );
  AOI21_X1 u2_u0_u0_U40 (.B1( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n132 ) , .A( u2_u0_u0_n165 ) , .B2( u2_u0_u0_n93 ) );
  OR3_X1 u2_u0_u0_U41 (.A3( u2_u0_u0_n152 ) , .A2( u2_u0_u0_n153 ) , .A1( u2_u0_u0_n154 ) , .ZN( u2_u0_u0_n155 ) );
  AOI21_X1 u2_u0_u0_U42 (.B2( u2_u0_u0_n150 ) , .B1( u2_u0_u0_n151 ) , .ZN( u2_u0_u0_n152 ) , .A( u2_u0_u0_n158 ) );
  AOI21_X1 u2_u0_u0_U43 (.A( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n145 ) , .B1( u2_u0_u0_n146 ) , .ZN( u2_u0_u0_n154 ) );
  AOI21_X1 u2_u0_u0_U44 (.A( u2_u0_u0_n147 ) , .B2( u2_u0_u0_n148 ) , .B1( u2_u0_u0_n149 ) , .ZN( u2_u0_u0_n153 ) );
  INV_X1 u2_u0_u0_U45 (.ZN( u2_u0_u0_n171 ) , .A( u2_u0_u0_n99 ) );
  OAI211_X1 u2_u0_u0_U46 (.C2( u2_u0_u0_n140 ) , .C1( u2_u0_u0_n161 ) , .A( u2_u0_u0_n169 ) , .B( u2_u0_u0_n98 ) , .ZN( u2_u0_u0_n99 ) );
  INV_X1 u2_u0_u0_U47 (.ZN( u2_u0_u0_n169 ) , .A( u2_u0_u0_n91 ) );
  AOI211_X1 u2_u0_u0_U48 (.C1( u2_u0_u0_n118 ) , .A( u2_u0_u0_n123 ) , .B( u2_u0_u0_n96 ) , .C2( u2_u0_u0_n97 ) , .ZN( u2_u0_u0_n98 ) );
  NOR2_X1 u2_u0_u0_U49 (.A2( u2_u0_X_4 ) , .A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n118 ) );
  NOR2_X1 u2_u0_u0_U5 (.A1( u2_u0_u0_n108 ) , .ZN( u2_u0_u0_n123 ) , .A2( u2_u0_u0_n158 ) );
  NOR2_X1 u2_u0_u0_U50 (.A2( u2_u0_X_2 ) , .ZN( u2_u0_u0_n103 ) , .A1( u2_u0_u0_n164 ) );
  NAND2_X1 u2_u0_u0_U51 (.A2( u2_u0_X_4 ) , .A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n144 ) );
  NOR2_X1 u2_u0_u0_U52 (.A2( u2_u0_X_5 ) , .ZN( u2_u0_u0_n136 ) , .A1( u2_u0_u0_n159 ) );
  NAND2_X1 u2_u0_u0_U53 (.A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n138 ) , .A2( u2_u0_u0_n159 ) );
  AND2_X1 u2_u0_u0_U54 (.A2( u2_u0_X_3 ) , .A1( u2_u0_X_6 ) , .ZN( u2_u0_u0_n102 ) );
  INV_X1 u2_u0_u0_U55 (.A( u2_u0_X_4 ) , .ZN( u2_u0_u0_n159 ) );
  INV_X1 u2_u0_u0_U56 (.A( u2_u0_X_2 ) , .ZN( u2_u0_u0_n163 ) );
  INV_X1 u2_u0_u0_U57 (.A( u2_u0_X_3 ) , .ZN( u2_u0_u0_n162 ) );
  INV_X1 u2_u0_u0_U58 (.A( u2_u0_u0_n126 ) , .ZN( u2_u0_u0_n168 ) );
  AOI211_X1 u2_u0_u0_U59 (.B( u2_u0_u0_n133 ) , .A( u2_u0_u0_n134 ) , .C2( u2_u0_u0_n135 ) , .C1( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n137 ) );
  AOI21_X1 u2_u0_u0_U6 (.B2( u2_u0_u0_n131 ) , .ZN( u2_u0_u0_n134 ) , .B1( u2_u0_u0_n151 ) , .A( u2_u0_u0_n158 ) );
  OR4_X1 u2_u0_u0_U60 (.ZN( u2_out0_17 ) , .A4( u2_u0_u0_n122 ) , .A2( u2_u0_u0_n123 ) , .A1( u2_u0_u0_n124 ) , .A3( u2_u0_u0_n170 ) );
  AOI21_X1 u2_u0_u0_U61 (.B2( u2_u0_u0_n107 ) , .ZN( u2_u0_u0_n124 ) , .B1( u2_u0_u0_n128 ) , .A( u2_u0_u0_n161 ) );
  INV_X1 u2_u0_u0_U62 (.A( u2_u0_u0_n111 ) , .ZN( u2_u0_u0_n170 ) );
  OR4_X1 u2_u0_u0_U63 (.ZN( u2_out0_31 ) , .A4( u2_u0_u0_n155 ) , .A2( u2_u0_u0_n156 ) , .A1( u2_u0_u0_n157 ) , .A3( u2_u0_u0_n173 ) );
  AOI21_X1 u2_u0_u0_U64 (.A( u2_u0_u0_n138 ) , .B2( u2_u0_u0_n139 ) , .B1( u2_u0_u0_n140 ) , .ZN( u2_u0_u0_n157 ) );
  INV_X1 u2_u0_u0_U65 (.ZN( u2_u0_u0_n174 ) , .A( u2_u0_u0_n89 ) );
  AOI211_X1 u2_u0_u0_U66 (.B( u2_u0_u0_n104 ) , .A( u2_u0_u0_n105 ) , .ZN( u2_u0_u0_n106 ) , .C2( u2_u0_u0_n113 ) , .C1( u2_u0_u0_n160 ) );
  AOI21_X1 u2_u0_u0_U67 (.B2( u2_u0_u0_n141 ) , .B1( u2_u0_u0_n142 ) , .ZN( u2_u0_u0_n156 ) , .A( u2_u0_u0_n161 ) );
  AOI21_X1 u2_u0_u0_U68 (.ZN( u2_u0_u0_n116 ) , .B2( u2_u0_u0_n142 ) , .A( u2_u0_u0_n144 ) , .B1( u2_u0_u0_n166 ) );
  NAND2_X1 u2_u0_u0_U69 (.ZN( u2_u0_u0_n148 ) , .A1( u2_u0_u0_n93 ) , .A2( u2_u0_u0_n95 ) );
  OAI21_X1 u2_u0_u0_U7 (.B1( u2_u0_u0_n150 ) , .B2( u2_u0_u0_n158 ) , .A( u2_u0_u0_n172 ) , .ZN( u2_u0_u0_n89 ) );
  NAND2_X1 u2_u0_u0_U70 (.A1( u2_u0_u0_n100 ) , .ZN( u2_u0_u0_n129 ) , .A2( u2_u0_u0_n95 ) );
  NAND2_X1 u2_u0_u0_U71 (.A1( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n128 ) , .A2( u2_u0_u0_n95 ) );
  INV_X1 u2_u0_u0_U72 (.A( u2_u0_u0_n142 ) , .ZN( u2_u0_u0_n165 ) );
  NOR2_X1 u2_u0_u0_U73 (.A2( u2_u0_X_1 ) , .A1( u2_u0_X_2 ) , .ZN( u2_u0_u0_n92 ) );
  NOR2_X1 u2_u0_u0_U74 (.A2( u2_u0_X_1 ) , .ZN( u2_u0_u0_n101 ) , .A1( u2_u0_u0_n163 ) );
  INV_X1 u2_u0_u0_U75 (.A( u2_u0_X_1 ) , .ZN( u2_u0_u0_n164 ) );
  AND2_X1 u2_u0_u0_U76 (.A1( u2_u0_X_6 ) , .A2( u2_u0_u0_n162 ) , .ZN( u2_u0_u0_n93 ) );
  NOR2_X1 u2_u0_u0_U77 (.A2( u2_u0_X_3 ) , .A1( u2_u0_X_6 ) , .ZN( u2_u0_u0_n94 ) );
  NOR2_X1 u2_u0_u0_U78 (.A2( u2_u0_X_6 ) , .ZN( u2_u0_u0_n100 ) , .A1( u2_u0_u0_n162 ) );
  OAI221_X1 u2_u0_u0_U79 (.C1( u2_u0_u0_n121 ) , .ZN( u2_u0_u0_n122 ) , .B2( u2_u0_u0_n127 ) , .A( u2_u0_u0_n143 ) , .B1( u2_u0_u0_n144 ) , .C2( u2_u0_u0_n147 ) );
  AND2_X1 u2_u0_u0_U8 (.A1( u2_u0_u0_n114 ) , .A2( u2_u0_u0_n121 ) , .ZN( u2_u0_u0_n146 ) );
  AOI21_X1 u2_u0_u0_U80 (.B1( u2_u0_u0_n132 ) , .ZN( u2_u0_u0_n133 ) , .A( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n166 ) );
  OAI22_X1 u2_u0_u0_U81 (.ZN( u2_u0_u0_n105 ) , .A2( u2_u0_u0_n132 ) , .B1( u2_u0_u0_n146 ) , .A1( u2_u0_u0_n147 ) , .B2( u2_u0_u0_n161 ) );
  NAND2_X1 u2_u0_u0_U82 (.ZN( u2_u0_u0_n110 ) , .A2( u2_u0_u0_n132 ) , .A1( u2_u0_u0_n145 ) );
  INV_X1 u2_u0_u0_U83 (.A( u2_u0_u0_n119 ) , .ZN( u2_u0_u0_n167 ) );
  NAND2_X1 u2_u0_u0_U84 (.A2( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n140 ) , .A1( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U85 (.A1( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n130 ) , .A2( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U86 (.ZN( u2_u0_u0_n108 ) , .A1( u2_u0_u0_n92 ) , .A2( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U87 (.ZN( u2_u0_u0_n142 ) , .A1( u2_u0_u0_n94 ) , .A2( u2_u0_u0_n95 ) );
  NAND3_X1 u2_u0_u0_U88 (.ZN( u2_out0_23 ) , .A3( u2_u0_u0_n137 ) , .A1( u2_u0_u0_n168 ) , .A2( u2_u0_u0_n171 ) );
  NAND3_X1 u2_u0_u0_U89 (.A3( u2_u0_u0_n127 ) , .A2( u2_u0_u0_n128 ) , .ZN( u2_u0_u0_n135 ) , .A1( u2_u0_u0_n150 ) );
  AND2_X1 u2_u0_u0_U9 (.A1( u2_u0_u0_n131 ) , .ZN( u2_u0_u0_n141 ) , .A2( u2_u0_u0_n150 ) );
  NAND3_X1 u2_u0_u0_U90 (.ZN( u2_u0_u0_n117 ) , .A3( u2_u0_u0_n132 ) , .A2( u2_u0_u0_n139 ) , .A1( u2_u0_u0_n148 ) );
  NAND3_X1 u2_u0_u0_U91 (.ZN( u2_u0_u0_n109 ) , .A2( u2_u0_u0_n114 ) , .A3( u2_u0_u0_n140 ) , .A1( u2_u0_u0_n149 ) );
  NAND3_X1 u2_u0_u0_U92 (.ZN( u2_out0_9 ) , .A3( u2_u0_u0_n106 ) , .A2( u2_u0_u0_n171 ) , .A1( u2_u0_u0_n174 ) );
  NAND3_X1 u2_u0_u0_U93 (.A2( u2_u0_u0_n128 ) , .A1( u2_u0_u0_n132 ) , .A3( u2_u0_u0_n146 ) , .ZN( u2_u0_u0_n97 ) );
  AOI21_X1 u2_u0_u1_U10 (.B2( u2_u0_u1_n155 ) , .B1( u2_u0_u1_n156 ) , .ZN( u2_u0_u1_n157 ) , .A( u2_u0_u1_n174 ) );
  NAND3_X1 u2_u0_u1_U100 (.ZN( u2_u0_u1_n113 ) , .A1( u2_u0_u1_n120 ) , .A3( u2_u0_u1_n133 ) , .A2( u2_u0_u1_n155 ) );
  NAND2_X1 u2_u0_u1_U11 (.ZN( u2_u0_u1_n140 ) , .A2( u2_u0_u1_n150 ) , .A1( u2_u0_u1_n155 ) );
  NAND2_X1 u2_u0_u1_U12 (.A1( u2_u0_u1_n131 ) , .ZN( u2_u0_u1_n147 ) , .A2( u2_u0_u1_n153 ) );
  AOI22_X1 u2_u0_u1_U13 (.B2( u2_u0_u1_n136 ) , .A2( u2_u0_u1_n137 ) , .ZN( u2_u0_u1_n143 ) , .A1( u2_u0_u1_n171 ) , .B1( u2_u0_u1_n173 ) );
  INV_X1 u2_u0_u1_U14 (.A( u2_u0_u1_n147 ) , .ZN( u2_u0_u1_n181 ) );
  INV_X1 u2_u0_u1_U15 (.A( u2_u0_u1_n139 ) , .ZN( u2_u0_u1_n174 ) );
  OR4_X1 u2_u0_u1_U16 (.A4( u2_u0_u1_n106 ) , .A3( u2_u0_u1_n107 ) , .ZN( u2_u0_u1_n108 ) , .A1( u2_u0_u1_n117 ) , .A2( u2_u0_u1_n184 ) );
  AOI21_X1 u2_u0_u1_U17 (.ZN( u2_u0_u1_n106 ) , .A( u2_u0_u1_n112 ) , .B1( u2_u0_u1_n154 ) , .B2( u2_u0_u1_n156 ) );
  AOI21_X1 u2_u0_u1_U18 (.ZN( u2_u0_u1_n107 ) , .B1( u2_u0_u1_n134 ) , .B2( u2_u0_u1_n149 ) , .A( u2_u0_u1_n174 ) );
  INV_X1 u2_u0_u1_U19 (.A( u2_u0_u1_n101 ) , .ZN( u2_u0_u1_n184 ) );
  INV_X1 u2_u0_u1_U20 (.A( u2_u0_u1_n112 ) , .ZN( u2_u0_u1_n171 ) );
  NAND2_X1 u2_u0_u1_U21 (.ZN( u2_u0_u1_n141 ) , .A1( u2_u0_u1_n153 ) , .A2( u2_u0_u1_n156 ) );
  AND2_X1 u2_u0_u1_U22 (.A1( u2_u0_u1_n123 ) , .ZN( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n161 ) );
  NAND2_X1 u2_u0_u1_U23 (.A2( u2_u0_u1_n115 ) , .A1( u2_u0_u1_n116 ) , .ZN( u2_u0_u1_n148 ) );
  NAND2_X1 u2_u0_u1_U24 (.A2( u2_u0_u1_n133 ) , .A1( u2_u0_u1_n135 ) , .ZN( u2_u0_u1_n159 ) );
  NAND2_X1 u2_u0_u1_U25 (.A2( u2_u0_u1_n115 ) , .A1( u2_u0_u1_n120 ) , .ZN( u2_u0_u1_n132 ) );
  INV_X1 u2_u0_u1_U26 (.A( u2_u0_u1_n154 ) , .ZN( u2_u0_u1_n178 ) );
  INV_X1 u2_u0_u1_U27 (.A( u2_u0_u1_n151 ) , .ZN( u2_u0_u1_n183 ) );
  AND2_X1 u2_u0_u1_U28 (.A1( u2_u0_u1_n129 ) , .A2( u2_u0_u1_n133 ) , .ZN( u2_u0_u1_n149 ) );
  INV_X1 u2_u0_u1_U29 (.A( u2_u0_u1_n131 ) , .ZN( u2_u0_u1_n180 ) );
  INV_X1 u2_u0_u1_U3 (.A( u2_u0_u1_n159 ) , .ZN( u2_u0_u1_n182 ) );
  AOI221_X1 u2_u0_u1_U30 (.B1( u2_u0_u1_n140 ) , .ZN( u2_u0_u1_n167 ) , .B2( u2_u0_u1_n172 ) , .C2( u2_u0_u1_n175 ) , .C1( u2_u0_u1_n178 ) , .A( u2_u0_u1_n188 ) );
  INV_X1 u2_u0_u1_U31 (.ZN( u2_u0_u1_n188 ) , .A( u2_u0_u1_n97 ) );
  AOI211_X1 u2_u0_u1_U32 (.A( u2_u0_u1_n118 ) , .C1( u2_u0_u1_n132 ) , .C2( u2_u0_u1_n139 ) , .B( u2_u0_u1_n96 ) , .ZN( u2_u0_u1_n97 ) );
  AOI21_X1 u2_u0_u1_U33 (.B2( u2_u0_u1_n121 ) , .B1( u2_u0_u1_n135 ) , .A( u2_u0_u1_n152 ) , .ZN( u2_u0_u1_n96 ) );
  OAI221_X1 u2_u0_u1_U34 (.A( u2_u0_u1_n119 ) , .C2( u2_u0_u1_n129 ) , .ZN( u2_u0_u1_n138 ) , .B2( u2_u0_u1_n152 ) , .C1( u2_u0_u1_n174 ) , .B1( u2_u0_u1_n187 ) );
  INV_X1 u2_u0_u1_U35 (.A( u2_u0_u1_n148 ) , .ZN( u2_u0_u1_n187 ) );
  AOI211_X1 u2_u0_u1_U36 (.B( u2_u0_u1_n117 ) , .A( u2_u0_u1_n118 ) , .ZN( u2_u0_u1_n119 ) , .C2( u2_u0_u1_n146 ) , .C1( u2_u0_u1_n159 ) );
  NOR2_X1 u2_u0_u1_U37 (.A1( u2_u0_u1_n168 ) , .A2( u2_u0_u1_n176 ) , .ZN( u2_u0_u1_n98 ) );
  AOI211_X1 u2_u0_u1_U38 (.B( u2_u0_u1_n162 ) , .A( u2_u0_u1_n163 ) , .C2( u2_u0_u1_n164 ) , .ZN( u2_u0_u1_n165 ) , .C1( u2_u0_u1_n171 ) );
  AOI21_X1 u2_u0_u1_U39 (.A( u2_u0_u1_n160 ) , .B2( u2_u0_u1_n161 ) , .ZN( u2_u0_u1_n162 ) , .B1( u2_u0_u1_n182 ) );
  AOI221_X1 u2_u0_u1_U4 (.A( u2_u0_u1_n138 ) , .C2( u2_u0_u1_n139 ) , .C1( u2_u0_u1_n140 ) , .B2( u2_u0_u1_n141 ) , .ZN( u2_u0_u1_n142 ) , .B1( u2_u0_u1_n175 ) );
  OR2_X1 u2_u0_u1_U40 (.A2( u2_u0_u1_n157 ) , .A1( u2_u0_u1_n158 ) , .ZN( u2_u0_u1_n163 ) );
  NAND2_X1 u2_u0_u1_U41 (.A1( u2_u0_u1_n128 ) , .ZN( u2_u0_u1_n146 ) , .A2( u2_u0_u1_n160 ) );
  NAND2_X1 u2_u0_u1_U42 (.A2( u2_u0_u1_n112 ) , .ZN( u2_u0_u1_n139 ) , .A1( u2_u0_u1_n152 ) );
  NAND2_X1 u2_u0_u1_U43 (.A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n156 ) , .A2( u2_u0_u1_n99 ) );
  NOR2_X1 u2_u0_u1_U44 (.ZN( u2_u0_u1_n117 ) , .A1( u2_u0_u1_n121 ) , .A2( u2_u0_u1_n160 ) );
  AOI21_X1 u2_u0_u1_U45 (.A( u2_u0_u1_n128 ) , .B2( u2_u0_u1_n129 ) , .ZN( u2_u0_u1_n130 ) , .B1( u2_u0_u1_n150 ) );
  NAND2_X1 u2_u0_u1_U46 (.ZN( u2_u0_u1_n112 ) , .A1( u2_u0_u1_n169 ) , .A2( u2_u0_u1_n170 ) );
  NAND2_X1 u2_u0_u1_U47 (.ZN( u2_u0_u1_n129 ) , .A2( u2_u0_u1_n95 ) , .A1( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U48 (.A1( u2_u0_u1_n102 ) , .ZN( u2_u0_u1_n154 ) , .A2( u2_u0_u1_n99 ) );
  NAND2_X1 u2_u0_u1_U49 (.A2( u2_u0_u1_n100 ) , .ZN( u2_u0_u1_n135 ) , .A1( u2_u0_u1_n99 ) );
  AOI211_X1 u2_u0_u1_U5 (.ZN( u2_u0_u1_n124 ) , .A( u2_u0_u1_n138 ) , .C2( u2_u0_u1_n139 ) , .B( u2_u0_u1_n145 ) , .C1( u2_u0_u1_n147 ) );
  AOI21_X1 u2_u0_u1_U50 (.A( u2_u0_u1_n152 ) , .B2( u2_u0_u1_n153 ) , .B1( u2_u0_u1_n154 ) , .ZN( u2_u0_u1_n158 ) );
  INV_X1 u2_u0_u1_U51 (.A( u2_u0_u1_n160 ) , .ZN( u2_u0_u1_n175 ) );
  NAND2_X1 u2_u0_u1_U52 (.A1( u2_u0_u1_n100 ) , .ZN( u2_u0_u1_n116 ) , .A2( u2_u0_u1_n95 ) );
  NAND2_X1 u2_u0_u1_U53 (.A1( u2_u0_u1_n102 ) , .ZN( u2_u0_u1_n131 ) , .A2( u2_u0_u1_n95 ) );
  NAND2_X1 u2_u0_u1_U54 (.A2( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n121 ) , .A1( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U55 (.A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n153 ) , .A2( u2_u0_u1_n98 ) );
  NAND2_X1 u2_u0_u1_U56 (.A2( u2_u0_u1_n104 ) , .A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n133 ) );
  NAND2_X1 u2_u0_u1_U57 (.ZN( u2_u0_u1_n150 ) , .A2( u2_u0_u1_n98 ) , .A1( u2_u0_u1_n99 ) );
  NAND2_X1 u2_u0_u1_U58 (.A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n155 ) , .A2( u2_u0_u1_n95 ) );
  OAI21_X1 u2_u0_u1_U59 (.ZN( u2_u0_u1_n109 ) , .B1( u2_u0_u1_n129 ) , .B2( u2_u0_u1_n160 ) , .A( u2_u0_u1_n167 ) );
  AOI22_X1 u2_u0_u1_U6 (.B2( u2_u0_u1_n113 ) , .A2( u2_u0_u1_n114 ) , .ZN( u2_u0_u1_n125 ) , .A1( u2_u0_u1_n171 ) , .B1( u2_u0_u1_n173 ) );
  NAND2_X1 u2_u0_u1_U60 (.A2( u2_u0_u1_n100 ) , .A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n120 ) );
  NAND2_X1 u2_u0_u1_U61 (.A1( u2_u0_u1_n102 ) , .A2( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n115 ) );
  NAND2_X1 u2_u0_u1_U62 (.A2( u2_u0_u1_n100 ) , .A1( u2_u0_u1_n104 ) , .ZN( u2_u0_u1_n151 ) );
  NAND2_X1 u2_u0_u1_U63 (.A2( u2_u0_u1_n103 ) , .A1( u2_u0_u1_n105 ) , .ZN( u2_u0_u1_n161 ) );
  INV_X1 u2_u0_u1_U64 (.A( u2_u0_u1_n152 ) , .ZN( u2_u0_u1_n173 ) );
  INV_X1 u2_u0_u1_U65 (.A( u2_u0_u1_n128 ) , .ZN( u2_u0_u1_n172 ) );
  NAND2_X1 u2_u0_u1_U66 (.A2( u2_u0_u1_n102 ) , .A1( u2_u0_u1_n103 ) , .ZN( u2_u0_u1_n123 ) );
  OAI21_X1 u2_u0_u1_U67 (.B2( u2_u0_u1_n123 ) , .ZN( u2_u0_u1_n145 ) , .B1( u2_u0_u1_n160 ) , .A( u2_u0_u1_n185 ) );
  INV_X1 u2_u0_u1_U68 (.A( u2_u0_u1_n122 ) , .ZN( u2_u0_u1_n185 ) );
  AOI21_X1 u2_u0_u1_U69 (.B2( u2_u0_u1_n120 ) , .B1( u2_u0_u1_n121 ) , .ZN( u2_u0_u1_n122 ) , .A( u2_u0_u1_n128 ) );
  NAND2_X1 u2_u0_u1_U7 (.ZN( u2_u0_u1_n114 ) , .A1( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n156 ) );
  NOR2_X1 u2_u0_u1_U70 (.A2( u2_u0_X_7 ) , .A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n95 ) );
  NOR2_X1 u2_u0_u1_U71 (.A1( u2_u0_X_12 ) , .A2( u2_u0_X_9 ) , .ZN( u2_u0_u1_n100 ) );
  NOR2_X1 u2_u0_u1_U72 (.A2( u2_u0_X_8 ) , .A1( u2_u0_u1_n177 ) , .ZN( u2_u0_u1_n99 ) );
  NOR2_X1 u2_u0_u1_U73 (.A2( u2_u0_X_12 ) , .ZN( u2_u0_u1_n102 ) , .A1( u2_u0_u1_n176 ) );
  NOR2_X1 u2_u0_u1_U74 (.A2( u2_u0_X_9 ) , .ZN( u2_u0_u1_n105 ) , .A1( u2_u0_u1_n168 ) );
  NAND2_X1 u2_u0_u1_U75 (.A1( u2_u0_X_10 ) , .ZN( u2_u0_u1_n160 ) , .A2( u2_u0_u1_n169 ) );
  NAND2_X1 u2_u0_u1_U76 (.A2( u2_u0_X_10 ) , .A1( u2_u0_X_11 ) , .ZN( u2_u0_u1_n152 ) );
  NAND2_X1 u2_u0_u1_U77 (.A1( u2_u0_X_11 ) , .ZN( u2_u0_u1_n128 ) , .A2( u2_u0_u1_n170 ) );
  AND2_X1 u2_u0_u1_U78 (.A2( u2_u0_X_7 ) , .A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n104 ) );
  AND2_X1 u2_u0_u1_U79 (.A1( u2_u0_X_8 ) , .ZN( u2_u0_u1_n103 ) , .A2( u2_u0_u1_n177 ) );
  NOR2_X1 u2_u0_u1_U8 (.A1( u2_u0_u1_n112 ) , .A2( u2_u0_u1_n116 ) , .ZN( u2_u0_u1_n118 ) );
  INV_X1 u2_u0_u1_U80 (.A( u2_u0_X_10 ) , .ZN( u2_u0_u1_n170 ) );
  INV_X1 u2_u0_u1_U81 (.A( u2_u0_X_9 ) , .ZN( u2_u0_u1_n176 ) );
  INV_X1 u2_u0_u1_U82 (.A( u2_u0_X_11 ) , .ZN( u2_u0_u1_n169 ) );
  INV_X1 u2_u0_u1_U83 (.A( u2_u0_X_12 ) , .ZN( u2_u0_u1_n168 ) );
  INV_X1 u2_u0_u1_U84 (.A( u2_u0_X_7 ) , .ZN( u2_u0_u1_n177 ) );
  NAND4_X1 u2_u0_u1_U85 (.ZN( u2_out0_28 ) , .A4( u2_u0_u1_n124 ) , .A3( u2_u0_u1_n125 ) , .A2( u2_u0_u1_n126 ) , .A1( u2_u0_u1_n127 ) );
  OAI21_X1 u2_u0_u1_U86 (.ZN( u2_u0_u1_n127 ) , .B2( u2_u0_u1_n139 ) , .B1( u2_u0_u1_n175 ) , .A( u2_u0_u1_n183 ) );
  OAI21_X1 u2_u0_u1_U87 (.ZN( u2_u0_u1_n126 ) , .B2( u2_u0_u1_n140 ) , .A( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n178 ) );
  NAND4_X1 u2_u0_u1_U88 (.ZN( u2_out0_18 ) , .A4( u2_u0_u1_n165 ) , .A3( u2_u0_u1_n166 ) , .A1( u2_u0_u1_n167 ) , .A2( u2_u0_u1_n186 ) );
  AOI22_X1 u2_u0_u1_U89 (.B2( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n147 ) , .A2( u2_u0_u1_n148 ) , .ZN( u2_u0_u1_n166 ) , .A1( u2_u0_u1_n172 ) );
  OAI21_X1 u2_u0_u1_U9 (.ZN( u2_u0_u1_n101 ) , .B1( u2_u0_u1_n141 ) , .A( u2_u0_u1_n146 ) , .B2( u2_u0_u1_n183 ) );
  INV_X1 u2_u0_u1_U90 (.A( u2_u0_u1_n145 ) , .ZN( u2_u0_u1_n186 ) );
  NAND4_X1 u2_u0_u1_U91 (.ZN( u2_out0_2 ) , .A4( u2_u0_u1_n142 ) , .A3( u2_u0_u1_n143 ) , .A2( u2_u0_u1_n144 ) , .A1( u2_u0_u1_n179 ) );
  OAI21_X1 u2_u0_u1_U92 (.B2( u2_u0_u1_n132 ) , .ZN( u2_u0_u1_n144 ) , .A( u2_u0_u1_n146 ) , .B1( u2_u0_u1_n180 ) );
  INV_X1 u2_u0_u1_U93 (.A( u2_u0_u1_n130 ) , .ZN( u2_u0_u1_n179 ) );
  OR4_X1 u2_u0_u1_U94 (.ZN( u2_out0_13 ) , .A4( u2_u0_u1_n108 ) , .A3( u2_u0_u1_n109 ) , .A2( u2_u0_u1_n110 ) , .A1( u2_u0_u1_n111 ) );
  AOI21_X1 u2_u0_u1_U95 (.ZN( u2_u0_u1_n111 ) , .A( u2_u0_u1_n128 ) , .B2( u2_u0_u1_n131 ) , .B1( u2_u0_u1_n135 ) );
  AOI21_X1 u2_u0_u1_U96 (.ZN( u2_u0_u1_n110 ) , .A( u2_u0_u1_n116 ) , .B1( u2_u0_u1_n152 ) , .B2( u2_u0_u1_n160 ) );
  NAND3_X1 u2_u0_u1_U97 (.A3( u2_u0_u1_n149 ) , .A2( u2_u0_u1_n150 ) , .A1( u2_u0_u1_n151 ) , .ZN( u2_u0_u1_n164 ) );
  NAND3_X1 u2_u0_u1_U98 (.A3( u2_u0_u1_n134 ) , .A2( u2_u0_u1_n135 ) , .ZN( u2_u0_u1_n136 ) , .A1( u2_u0_u1_n151 ) );
  NAND3_X1 u2_u0_u1_U99 (.A1( u2_u0_u1_n133 ) , .ZN( u2_u0_u1_n137 ) , .A2( u2_u0_u1_n154 ) , .A3( u2_u0_u1_n181 ) );
  OAI22_X1 u2_u0_u2_U10 (.B1( u2_u0_u2_n151 ) , .A2( u2_u0_u2_n152 ) , .A1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n160 ) , .B2( u2_u0_u2_n168 ) );
  NAND3_X1 u2_u0_u2_U100 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n98 ) );
  NOR3_X1 u2_u0_u2_U11 (.A1( u2_u0_u2_n150 ) , .ZN( u2_u0_u2_n151 ) , .A3( u2_u0_u2_n175 ) , .A2( u2_u0_u2_n188 ) );
  AOI21_X1 u2_u0_u2_U12 (.B2( u2_u0_u2_n123 ) , .ZN( u2_u0_u2_n125 ) , .A( u2_u0_u2_n171 ) , .B1( u2_u0_u2_n184 ) );
  INV_X1 u2_u0_u2_U13 (.A( u2_u0_u2_n150 ) , .ZN( u2_u0_u2_n184 ) );
  AOI21_X1 u2_u0_u2_U14 (.ZN( u2_u0_u2_n144 ) , .B2( u2_u0_u2_n155 ) , .A( u2_u0_u2_n172 ) , .B1( u2_u0_u2_n185 ) );
  AOI21_X1 u2_u0_u2_U15 (.B2( u2_u0_u2_n143 ) , .ZN( u2_u0_u2_n145 ) , .B1( u2_u0_u2_n152 ) , .A( u2_u0_u2_n171 ) );
  INV_X1 u2_u0_u2_U16 (.A( u2_u0_u2_n156 ) , .ZN( u2_u0_u2_n171 ) );
  INV_X1 u2_u0_u2_U17 (.A( u2_u0_u2_n120 ) , .ZN( u2_u0_u2_n188 ) );
  NAND2_X1 u2_u0_u2_U18 (.A2( u2_u0_u2_n122 ) , .ZN( u2_u0_u2_n150 ) , .A1( u2_u0_u2_n152 ) );
  INV_X1 u2_u0_u2_U19 (.A( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n170 ) );
  INV_X1 u2_u0_u2_U20 (.A( u2_u0_u2_n137 ) , .ZN( u2_u0_u2_n173 ) );
  NAND2_X1 u2_u0_u2_U21 (.A1( u2_u0_u2_n132 ) , .A2( u2_u0_u2_n139 ) , .ZN( u2_u0_u2_n157 ) );
  INV_X1 u2_u0_u2_U22 (.A( u2_u0_u2_n113 ) , .ZN( u2_u0_u2_n178 ) );
  INV_X1 u2_u0_u2_U23 (.A( u2_u0_u2_n139 ) , .ZN( u2_u0_u2_n175 ) );
  INV_X1 u2_u0_u2_U24 (.A( u2_u0_u2_n155 ) , .ZN( u2_u0_u2_n181 ) );
  INV_X1 u2_u0_u2_U25 (.A( u2_u0_u2_n119 ) , .ZN( u2_u0_u2_n177 ) );
  INV_X1 u2_u0_u2_U26 (.A( u2_u0_u2_n116 ) , .ZN( u2_u0_u2_n180 ) );
  INV_X1 u2_u0_u2_U27 (.A( u2_u0_u2_n131 ) , .ZN( u2_u0_u2_n179 ) );
  INV_X1 u2_u0_u2_U28 (.A( u2_u0_u2_n154 ) , .ZN( u2_u0_u2_n176 ) );
  NAND2_X1 u2_u0_u2_U29 (.A2( u2_u0_u2_n116 ) , .A1( u2_u0_u2_n117 ) , .ZN( u2_u0_u2_n118 ) );
  NOR2_X1 u2_u0_u2_U3 (.ZN( u2_u0_u2_n121 ) , .A2( u2_u0_u2_n177 ) , .A1( u2_u0_u2_n180 ) );
  INV_X1 u2_u0_u2_U30 (.A( u2_u0_u2_n132 ) , .ZN( u2_u0_u2_n182 ) );
  INV_X1 u2_u0_u2_U31 (.A( u2_u0_u2_n158 ) , .ZN( u2_u0_u2_n183 ) );
  OAI21_X1 u2_u0_u2_U32 (.A( u2_u0_u2_n156 ) , .B1( u2_u0_u2_n157 ) , .ZN( u2_u0_u2_n158 ) , .B2( u2_u0_u2_n179 ) );
  NOR2_X1 u2_u0_u2_U33 (.ZN( u2_u0_u2_n156 ) , .A1( u2_u0_u2_n166 ) , .A2( u2_u0_u2_n169 ) );
  NOR2_X1 u2_u0_u2_U34 (.A2( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n137 ) , .A1( u2_u0_u2_n140 ) );
  NOR2_X1 u2_u0_u2_U35 (.A2( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n153 ) , .A1( u2_u0_u2_n156 ) );
  AOI211_X1 u2_u0_u2_U36 (.ZN( u2_u0_u2_n130 ) , .C1( u2_u0_u2_n138 ) , .C2( u2_u0_u2_n179 ) , .B( u2_u0_u2_n96 ) , .A( u2_u0_u2_n97 ) );
  OAI22_X1 u2_u0_u2_U37 (.B1( u2_u0_u2_n133 ) , .A2( u2_u0_u2_n137 ) , .A1( u2_u0_u2_n152 ) , .B2( u2_u0_u2_n168 ) , .ZN( u2_u0_u2_n97 ) );
  OAI221_X1 u2_u0_u2_U38 (.B1( u2_u0_u2_n113 ) , .C1( u2_u0_u2_n132 ) , .A( u2_u0_u2_n149 ) , .B2( u2_u0_u2_n171 ) , .C2( u2_u0_u2_n172 ) , .ZN( u2_u0_u2_n96 ) );
  OAI221_X1 u2_u0_u2_U39 (.A( u2_u0_u2_n115 ) , .C2( u2_u0_u2_n123 ) , .B2( u2_u0_u2_n143 ) , .B1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n163 ) , .C1( u2_u0_u2_n168 ) );
  INV_X1 u2_u0_u2_U4 (.A( u2_u0_u2_n134 ) , .ZN( u2_u0_u2_n185 ) );
  OAI21_X1 u2_u0_u2_U40 (.A( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n115 ) , .B1( u2_u0_u2_n176 ) , .B2( u2_u0_u2_n178 ) );
  OAI221_X1 u2_u0_u2_U41 (.A( u2_u0_u2_n135 ) , .B2( u2_u0_u2_n136 ) , .B1( u2_u0_u2_n137 ) , .ZN( u2_u0_u2_n162 ) , .C2( u2_u0_u2_n167 ) , .C1( u2_u0_u2_n185 ) );
  AND3_X1 u2_u0_u2_U42 (.A3( u2_u0_u2_n131 ) , .A2( u2_u0_u2_n132 ) , .A1( u2_u0_u2_n133 ) , .ZN( u2_u0_u2_n136 ) );
  AOI22_X1 u2_u0_u2_U43 (.ZN( u2_u0_u2_n135 ) , .B1( u2_u0_u2_n140 ) , .A1( u2_u0_u2_n156 ) , .B2( u2_u0_u2_n180 ) , .A2( u2_u0_u2_n188 ) );
  AOI21_X1 u2_u0_u2_U44 (.ZN( u2_u0_u2_n149 ) , .B1( u2_u0_u2_n173 ) , .B2( u2_u0_u2_n188 ) , .A( u2_u0_u2_n95 ) );
  AND3_X1 u2_u0_u2_U45 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n156 ) , .ZN( u2_u0_u2_n95 ) );
  OAI21_X1 u2_u0_u2_U46 (.A( u2_u0_u2_n141 ) , .B2( u2_u0_u2_n142 ) , .ZN( u2_u0_u2_n146 ) , .B1( u2_u0_u2_n153 ) );
  OAI21_X1 u2_u0_u2_U47 (.A( u2_u0_u2_n140 ) , .ZN( u2_u0_u2_n141 ) , .B1( u2_u0_u2_n176 ) , .B2( u2_u0_u2_n177 ) );
  NOR3_X1 u2_u0_u2_U48 (.ZN( u2_u0_u2_n142 ) , .A3( u2_u0_u2_n175 ) , .A2( u2_u0_u2_n178 ) , .A1( u2_u0_u2_n181 ) );
  OAI21_X1 u2_u0_u2_U49 (.A( u2_u0_u2_n101 ) , .B2( u2_u0_u2_n121 ) , .B1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n164 ) );
  NOR4_X1 u2_u0_u2_U5 (.A4( u2_u0_u2_n124 ) , .A3( u2_u0_u2_n125 ) , .A2( u2_u0_u2_n126 ) , .A1( u2_u0_u2_n127 ) , .ZN( u2_u0_u2_n128 ) );
  NAND2_X1 u2_u0_u2_U50 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n155 ) );
  NAND2_X1 u2_u0_u2_U51 (.A2( u2_u0_u2_n105 ) , .A1( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n143 ) );
  NAND2_X1 u2_u0_u2_U52 (.A1( u2_u0_u2_n104 ) , .A2( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n152 ) );
  NAND2_X1 u2_u0_u2_U53 (.A1( u2_u0_u2_n100 ) , .A2( u2_u0_u2_n105 ) , .ZN( u2_u0_u2_n132 ) );
  INV_X1 u2_u0_u2_U54 (.A( u2_u0_u2_n140 ) , .ZN( u2_u0_u2_n168 ) );
  INV_X1 u2_u0_u2_U55 (.A( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n167 ) );
  NAND2_X1 u2_u0_u2_U56 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n113 ) );
  NAND2_X1 u2_u0_u2_U57 (.A1( u2_u0_u2_n106 ) , .A2( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n131 ) );
  NAND2_X1 u2_u0_u2_U58 (.A1( u2_u0_u2_n103 ) , .A2( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n139 ) );
  NAND2_X1 u2_u0_u2_U59 (.A1( u2_u0_u2_n103 ) , .A2( u2_u0_u2_n105 ) , .ZN( u2_u0_u2_n133 ) );
  AOI21_X1 u2_u0_u2_U6 (.B2( u2_u0_u2_n119 ) , .ZN( u2_u0_u2_n127 ) , .A( u2_u0_u2_n137 ) , .B1( u2_u0_u2_n155 ) );
  NAND2_X1 u2_u0_u2_U60 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n103 ) , .ZN( u2_u0_u2_n154 ) );
  NAND2_X1 u2_u0_u2_U61 (.A2( u2_u0_u2_n103 ) , .A1( u2_u0_u2_n104 ) , .ZN( u2_u0_u2_n119 ) );
  NAND2_X1 u2_u0_u2_U62 (.A2( u2_u0_u2_n107 ) , .A1( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n123 ) );
  NAND2_X1 u2_u0_u2_U63 (.A1( u2_u0_u2_n104 ) , .A2( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n122 ) );
  INV_X1 u2_u0_u2_U64 (.A( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n172 ) );
  NAND2_X1 u2_u0_u2_U65 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n102 ) , .ZN( u2_u0_u2_n116 ) );
  NAND2_X1 u2_u0_u2_U66 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n120 ) );
  NAND2_X1 u2_u0_u2_U67 (.A2( u2_u0_u2_n105 ) , .A1( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n117 ) );
  INV_X1 u2_u0_u2_U68 (.ZN( u2_u0_u2_n187 ) , .A( u2_u0_u2_n99 ) );
  OAI21_X1 u2_u0_u2_U69 (.B1( u2_u0_u2_n137 ) , .B2( u2_u0_u2_n143 ) , .A( u2_u0_u2_n98 ) , .ZN( u2_u0_u2_n99 ) );
  AOI21_X1 u2_u0_u2_U7 (.ZN( u2_u0_u2_n124 ) , .B1( u2_u0_u2_n131 ) , .B2( u2_u0_u2_n143 ) , .A( u2_u0_u2_n172 ) );
  NOR2_X1 u2_u0_u2_U70 (.A2( u2_u0_X_16 ) , .ZN( u2_u0_u2_n140 ) , .A1( u2_u0_u2_n166 ) );
  NOR2_X1 u2_u0_u2_U71 (.A2( u2_u0_X_13 ) , .A1( u2_u0_X_14 ) , .ZN( u2_u0_u2_n100 ) );
  NOR2_X1 u2_u0_u2_U72 (.A2( u2_u0_X_16 ) , .A1( u2_u0_X_17 ) , .ZN( u2_u0_u2_n138 ) );
  NOR2_X1 u2_u0_u2_U73 (.A2( u2_u0_X_15 ) , .A1( u2_u0_X_18 ) , .ZN( u2_u0_u2_n104 ) );
  NOR2_X1 u2_u0_u2_U74 (.A2( u2_u0_X_14 ) , .ZN( u2_u0_u2_n103 ) , .A1( u2_u0_u2_n174 ) );
  NOR2_X1 u2_u0_u2_U75 (.A2( u2_u0_X_15 ) , .ZN( u2_u0_u2_n102 ) , .A1( u2_u0_u2_n165 ) );
  NOR2_X1 u2_u0_u2_U76 (.A2( u2_u0_X_17 ) , .ZN( u2_u0_u2_n114 ) , .A1( u2_u0_u2_n169 ) );
  AND2_X1 u2_u0_u2_U77 (.A1( u2_u0_X_15 ) , .ZN( u2_u0_u2_n105 ) , .A2( u2_u0_u2_n165 ) );
  AND2_X1 u2_u0_u2_U78 (.A2( u2_u0_X_15 ) , .A1( u2_u0_X_18 ) , .ZN( u2_u0_u2_n107 ) );
  AND2_X1 u2_u0_u2_U79 (.A1( u2_u0_X_14 ) , .ZN( u2_u0_u2_n106 ) , .A2( u2_u0_u2_n174 ) );
  AOI21_X1 u2_u0_u2_U8 (.B2( u2_u0_u2_n120 ) , .B1( u2_u0_u2_n121 ) , .ZN( u2_u0_u2_n126 ) , .A( u2_u0_u2_n167 ) );
  AND2_X1 u2_u0_u2_U80 (.A1( u2_u0_X_13 ) , .A2( u2_u0_X_14 ) , .ZN( u2_u0_u2_n108 ) );
  INV_X1 u2_u0_u2_U81 (.A( u2_u0_X_16 ) , .ZN( u2_u0_u2_n169 ) );
  INV_X1 u2_u0_u2_U82 (.A( u2_u0_X_17 ) , .ZN( u2_u0_u2_n166 ) );
  INV_X1 u2_u0_u2_U83 (.A( u2_u0_X_13 ) , .ZN( u2_u0_u2_n174 ) );
  INV_X1 u2_u0_u2_U84 (.A( u2_u0_X_18 ) , .ZN( u2_u0_u2_n165 ) );
  NAND4_X1 u2_u0_u2_U85 (.ZN( u2_out0_30 ) , .A4( u2_u0_u2_n147 ) , .A3( u2_u0_u2_n148 ) , .A2( u2_u0_u2_n149 ) , .A1( u2_u0_u2_n187 ) );
  NOR3_X1 u2_u0_u2_U86 (.A3( u2_u0_u2_n144 ) , .A2( u2_u0_u2_n145 ) , .A1( u2_u0_u2_n146 ) , .ZN( u2_u0_u2_n147 ) );
  AOI21_X1 u2_u0_u2_U87 (.B2( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n148 ) , .A( u2_u0_u2_n162 ) , .B1( u2_u0_u2_n182 ) );
  NAND4_X1 u2_u0_u2_U88 (.ZN( u2_out0_24 ) , .A4( u2_u0_u2_n111 ) , .A3( u2_u0_u2_n112 ) , .A1( u2_u0_u2_n130 ) , .A2( u2_u0_u2_n187 ) );
  AOI221_X1 u2_u0_u2_U89 (.A( u2_u0_u2_n109 ) , .B1( u2_u0_u2_n110 ) , .ZN( u2_u0_u2_n111 ) , .C1( u2_u0_u2_n134 ) , .C2( u2_u0_u2_n170 ) , .B2( u2_u0_u2_n173 ) );
  OAI22_X1 u2_u0_u2_U9 (.ZN( u2_u0_u2_n109 ) , .A2( u2_u0_u2_n113 ) , .B2( u2_u0_u2_n133 ) , .B1( u2_u0_u2_n167 ) , .A1( u2_u0_u2_n168 ) );
  AOI21_X1 u2_u0_u2_U90 (.ZN( u2_u0_u2_n112 ) , .B2( u2_u0_u2_n156 ) , .A( u2_u0_u2_n164 ) , .B1( u2_u0_u2_n181 ) );
  NAND4_X1 u2_u0_u2_U91 (.ZN( u2_out0_16 ) , .A4( u2_u0_u2_n128 ) , .A3( u2_u0_u2_n129 ) , .A1( u2_u0_u2_n130 ) , .A2( u2_u0_u2_n186 ) );
  AOI22_X1 u2_u0_u2_U92 (.A2( u2_u0_u2_n118 ) , .ZN( u2_u0_u2_n129 ) , .A1( u2_u0_u2_n140 ) , .B1( u2_u0_u2_n157 ) , .B2( u2_u0_u2_n170 ) );
  INV_X1 u2_u0_u2_U93 (.A( u2_u0_u2_n163 ) , .ZN( u2_u0_u2_n186 ) );
  OR4_X1 u2_u0_u2_U94 (.ZN( u2_out0_6 ) , .A4( u2_u0_u2_n161 ) , .A3( u2_u0_u2_n162 ) , .A2( u2_u0_u2_n163 ) , .A1( u2_u0_u2_n164 ) );
  OR3_X1 u2_u0_u2_U95 (.A2( u2_u0_u2_n159 ) , .A1( u2_u0_u2_n160 ) , .ZN( u2_u0_u2_n161 ) , .A3( u2_u0_u2_n183 ) );
  AOI21_X1 u2_u0_u2_U96 (.B2( u2_u0_u2_n154 ) , .B1( u2_u0_u2_n155 ) , .ZN( u2_u0_u2_n159 ) , .A( u2_u0_u2_n167 ) );
  NAND3_X1 u2_u0_u2_U97 (.A2( u2_u0_u2_n117 ) , .A1( u2_u0_u2_n122 ) , .A3( u2_u0_u2_n123 ) , .ZN( u2_u0_u2_n134 ) );
  NAND3_X1 u2_u0_u2_U98 (.ZN( u2_u0_u2_n110 ) , .A2( u2_u0_u2_n131 ) , .A3( u2_u0_u2_n139 ) , .A1( u2_u0_u2_n154 ) );
  NAND3_X1 u2_u0_u2_U99 (.A2( u2_u0_u2_n100 ) , .ZN( u2_u0_u2_n101 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n114 ) );
  XOR2_X1 u2_u10_U13 (.B( u2_K11_42 ) , .A( u2_R9_29 ) , .Z( u2_u10_X_42 ) );
  XOR2_X1 u2_u10_U14 (.B( u2_K11_41 ) , .A( u2_R9_28 ) , .Z( u2_u10_X_41 ) );
  XOR2_X1 u2_u10_U15 (.B( u2_K11_40 ) , .A( u2_R9_27 ) , .Z( u2_u10_X_40 ) );
  XOR2_X1 u2_u10_U17 (.B( u2_K11_39 ) , .A( u2_R9_26 ) , .Z( u2_u10_X_39 ) );
  XOR2_X1 u2_u10_U18 (.B( u2_K11_38 ) , .A( u2_R9_25 ) , .Z( u2_u10_X_38 ) );
  XOR2_X1 u2_u10_U19 (.B( u2_K11_37 ) , .A( u2_R9_24 ) , .Z( u2_u10_X_37 ) );
  XOR2_X1 u2_u10_U20 (.B( u2_K11_36 ) , .A( u2_R9_25 ) , .Z( u2_u10_X_36 ) );
  XOR2_X1 u2_u10_U21 (.B( u2_K11_35 ) , .A( u2_R9_24 ) , .Z( u2_u10_X_35 ) );
  XOR2_X1 u2_u10_U22 (.B( u2_K11_34 ) , .A( u2_R9_23 ) , .Z( u2_u10_X_34 ) );
  XOR2_X1 u2_u10_U23 (.B( u2_K11_33 ) , .A( u2_R9_22 ) , .Z( u2_u10_X_33 ) );
  XOR2_X1 u2_u10_U24 (.B( u2_K11_32 ) , .A( u2_R9_21 ) , .Z( u2_u10_X_32 ) );
  XOR2_X1 u2_u10_U25 (.B( u2_K11_31 ) , .A( u2_R9_20 ) , .Z( u2_u10_X_31 ) );
  INV_X1 u2_u10_u5_U10 (.A( u2_u10_u5_n121 ) , .ZN( u2_u10_u5_n177 ) );
  NOR3_X1 u2_u10_u5_U100 (.A3( u2_u10_u5_n141 ) , .A1( u2_u10_u5_n142 ) , .ZN( u2_u10_u5_n143 ) , .A2( u2_u10_u5_n191 ) );
  NAND4_X1 u2_u10_u5_U101 (.ZN( u2_out10_4 ) , .A4( u2_u10_u5_n112 ) , .A2( u2_u10_u5_n113 ) , .A1( u2_u10_u5_n114 ) , .A3( u2_u10_u5_n195 ) );
  AOI211_X1 u2_u10_u5_U102 (.A( u2_u10_u5_n110 ) , .C1( u2_u10_u5_n111 ) , .ZN( u2_u10_u5_n112 ) , .B( u2_u10_u5_n118 ) , .C2( u2_u10_u5_n177 ) );
  AOI222_X1 u2_u10_u5_U103 (.ZN( u2_u10_u5_n113 ) , .A1( u2_u10_u5_n131 ) , .C1( u2_u10_u5_n148 ) , .B2( u2_u10_u5_n174 ) , .C2( u2_u10_u5_n178 ) , .A2( u2_u10_u5_n179 ) , .B1( u2_u10_u5_n99 ) );
  NAND3_X1 u2_u10_u5_U104 (.A2( u2_u10_u5_n154 ) , .A3( u2_u10_u5_n158 ) , .A1( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n99 ) );
  NOR2_X1 u2_u10_u5_U11 (.ZN( u2_u10_u5_n160 ) , .A2( u2_u10_u5_n173 ) , .A1( u2_u10_u5_n177 ) );
  INV_X1 u2_u10_u5_U12 (.A( u2_u10_u5_n150 ) , .ZN( u2_u10_u5_n174 ) );
  AOI21_X1 u2_u10_u5_U13 (.A( u2_u10_u5_n160 ) , .B2( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n162 ) , .B1( u2_u10_u5_n192 ) );
  INV_X1 u2_u10_u5_U14 (.A( u2_u10_u5_n159 ) , .ZN( u2_u10_u5_n192 ) );
  AOI21_X1 u2_u10_u5_U15 (.A( u2_u10_u5_n156 ) , .B2( u2_u10_u5_n157 ) , .B1( u2_u10_u5_n158 ) , .ZN( u2_u10_u5_n163 ) );
  AOI21_X1 u2_u10_u5_U16 (.B2( u2_u10_u5_n139 ) , .B1( u2_u10_u5_n140 ) , .ZN( u2_u10_u5_n141 ) , .A( u2_u10_u5_n150 ) );
  OAI21_X1 u2_u10_u5_U17 (.A( u2_u10_u5_n133 ) , .B2( u2_u10_u5_n134 ) , .B1( u2_u10_u5_n135 ) , .ZN( u2_u10_u5_n142 ) );
  OAI21_X1 u2_u10_u5_U18 (.ZN( u2_u10_u5_n133 ) , .B2( u2_u10_u5_n147 ) , .A( u2_u10_u5_n173 ) , .B1( u2_u10_u5_n188 ) );
  NAND2_X1 u2_u10_u5_U19 (.A2( u2_u10_u5_n119 ) , .A1( u2_u10_u5_n123 ) , .ZN( u2_u10_u5_n137 ) );
  INV_X1 u2_u10_u5_U20 (.A( u2_u10_u5_n155 ) , .ZN( u2_u10_u5_n194 ) );
  NAND2_X1 u2_u10_u5_U21 (.A1( u2_u10_u5_n121 ) , .ZN( u2_u10_u5_n132 ) , .A2( u2_u10_u5_n172 ) );
  NAND2_X1 u2_u10_u5_U22 (.A2( u2_u10_u5_n122 ) , .ZN( u2_u10_u5_n136 ) , .A1( u2_u10_u5_n154 ) );
  NAND2_X1 u2_u10_u5_U23 (.A2( u2_u10_u5_n119 ) , .A1( u2_u10_u5_n120 ) , .ZN( u2_u10_u5_n159 ) );
  INV_X1 u2_u10_u5_U24 (.A( u2_u10_u5_n156 ) , .ZN( u2_u10_u5_n175 ) );
  INV_X1 u2_u10_u5_U25 (.A( u2_u10_u5_n158 ) , .ZN( u2_u10_u5_n188 ) );
  INV_X1 u2_u10_u5_U26 (.A( u2_u10_u5_n152 ) , .ZN( u2_u10_u5_n179 ) );
  INV_X1 u2_u10_u5_U27 (.A( u2_u10_u5_n140 ) , .ZN( u2_u10_u5_n182 ) );
  INV_X1 u2_u10_u5_U28 (.A( u2_u10_u5_n151 ) , .ZN( u2_u10_u5_n183 ) );
  INV_X1 u2_u10_u5_U29 (.A( u2_u10_u5_n123 ) , .ZN( u2_u10_u5_n185 ) );
  NOR2_X1 u2_u10_u5_U3 (.ZN( u2_u10_u5_n134 ) , .A1( u2_u10_u5_n183 ) , .A2( u2_u10_u5_n190 ) );
  INV_X1 u2_u10_u5_U30 (.A( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n184 ) );
  INV_X1 u2_u10_u5_U31 (.A( u2_u10_u5_n139 ) , .ZN( u2_u10_u5_n189 ) );
  INV_X1 u2_u10_u5_U32 (.A( u2_u10_u5_n157 ) , .ZN( u2_u10_u5_n190 ) );
  INV_X1 u2_u10_u5_U33 (.A( u2_u10_u5_n120 ) , .ZN( u2_u10_u5_n193 ) );
  NAND2_X1 u2_u10_u5_U34 (.ZN( u2_u10_u5_n111 ) , .A1( u2_u10_u5_n140 ) , .A2( u2_u10_u5_n155 ) );
  NOR2_X1 u2_u10_u5_U35 (.ZN( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n170 ) , .A2( u2_u10_u5_n180 ) );
  INV_X1 u2_u10_u5_U36 (.A( u2_u10_u5_n117 ) , .ZN( u2_u10_u5_n196 ) );
  OAI221_X1 u2_u10_u5_U37 (.A( u2_u10_u5_n116 ) , .ZN( u2_u10_u5_n117 ) , .B2( u2_u10_u5_n119 ) , .C1( u2_u10_u5_n153 ) , .C2( u2_u10_u5_n158 ) , .B1( u2_u10_u5_n172 ) );
  AOI222_X1 u2_u10_u5_U38 (.ZN( u2_u10_u5_n116 ) , .B2( u2_u10_u5_n145 ) , .C1( u2_u10_u5_n148 ) , .A2( u2_u10_u5_n174 ) , .C2( u2_u10_u5_n177 ) , .B1( u2_u10_u5_n187 ) , .A1( u2_u10_u5_n193 ) );
  INV_X1 u2_u10_u5_U39 (.A( u2_u10_u5_n115 ) , .ZN( u2_u10_u5_n187 ) );
  INV_X1 u2_u10_u5_U4 (.A( u2_u10_u5_n138 ) , .ZN( u2_u10_u5_n191 ) );
  AOI22_X1 u2_u10_u5_U40 (.B2( u2_u10_u5_n131 ) , .A2( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n169 ) , .B1( u2_u10_u5_n174 ) , .A1( u2_u10_u5_n185 ) );
  NOR2_X1 u2_u10_u5_U41 (.A1( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n150 ) , .A2( u2_u10_u5_n173 ) );
  AOI21_X1 u2_u10_u5_U42 (.A( u2_u10_u5_n118 ) , .B2( u2_u10_u5_n145 ) , .ZN( u2_u10_u5_n168 ) , .B1( u2_u10_u5_n186 ) );
  INV_X1 u2_u10_u5_U43 (.A( u2_u10_u5_n122 ) , .ZN( u2_u10_u5_n186 ) );
  NOR2_X1 u2_u10_u5_U44 (.A1( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n152 ) , .A2( u2_u10_u5_n176 ) );
  NOR2_X1 u2_u10_u5_U45 (.A1( u2_u10_u5_n115 ) , .ZN( u2_u10_u5_n118 ) , .A2( u2_u10_u5_n153 ) );
  NOR2_X1 u2_u10_u5_U46 (.A2( u2_u10_u5_n145 ) , .ZN( u2_u10_u5_n156 ) , .A1( u2_u10_u5_n174 ) );
  NOR2_X1 u2_u10_u5_U47 (.ZN( u2_u10_u5_n121 ) , .A2( u2_u10_u5_n145 ) , .A1( u2_u10_u5_n176 ) );
  AOI22_X1 u2_u10_u5_U48 (.ZN( u2_u10_u5_n114 ) , .A2( u2_u10_u5_n137 ) , .A1( u2_u10_u5_n145 ) , .B2( u2_u10_u5_n175 ) , .B1( u2_u10_u5_n193 ) );
  OAI211_X1 u2_u10_u5_U49 (.B( u2_u10_u5_n124 ) , .A( u2_u10_u5_n125 ) , .C2( u2_u10_u5_n126 ) , .C1( u2_u10_u5_n127 ) , .ZN( u2_u10_u5_n128 ) );
  OAI21_X1 u2_u10_u5_U5 (.B2( u2_u10_u5_n136 ) , .B1( u2_u10_u5_n137 ) , .ZN( u2_u10_u5_n138 ) , .A( u2_u10_u5_n177 ) );
  NOR3_X1 u2_u10_u5_U50 (.ZN( u2_u10_u5_n127 ) , .A1( u2_u10_u5_n136 ) , .A3( u2_u10_u5_n148 ) , .A2( u2_u10_u5_n182 ) );
  OAI21_X1 u2_u10_u5_U51 (.ZN( u2_u10_u5_n124 ) , .A( u2_u10_u5_n177 ) , .B2( u2_u10_u5_n183 ) , .B1( u2_u10_u5_n189 ) );
  OAI21_X1 u2_u10_u5_U52 (.ZN( u2_u10_u5_n125 ) , .A( u2_u10_u5_n174 ) , .B2( u2_u10_u5_n185 ) , .B1( u2_u10_u5_n190 ) );
  AOI21_X1 u2_u10_u5_U53 (.A( u2_u10_u5_n153 ) , .B2( u2_u10_u5_n154 ) , .B1( u2_u10_u5_n155 ) , .ZN( u2_u10_u5_n164 ) );
  AOI21_X1 u2_u10_u5_U54 (.ZN( u2_u10_u5_n110 ) , .B1( u2_u10_u5_n122 ) , .B2( u2_u10_u5_n139 ) , .A( u2_u10_u5_n153 ) );
  INV_X1 u2_u10_u5_U55 (.A( u2_u10_u5_n153 ) , .ZN( u2_u10_u5_n176 ) );
  INV_X1 u2_u10_u5_U56 (.A( u2_u10_u5_n126 ) , .ZN( u2_u10_u5_n173 ) );
  AND2_X1 u2_u10_u5_U57 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n147 ) );
  AND2_X1 u2_u10_u5_U58 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n148 ) );
  NAND2_X1 u2_u10_u5_U59 (.A1( u2_u10_u5_n105 ) , .A2( u2_u10_u5_n106 ) , .ZN( u2_u10_u5_n158 ) );
  INV_X1 u2_u10_u5_U6 (.A( u2_u10_u5_n135 ) , .ZN( u2_u10_u5_n178 ) );
  NAND2_X1 u2_u10_u5_U60 (.A2( u2_u10_u5_n108 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n139 ) );
  NAND2_X1 u2_u10_u5_U61 (.A1( u2_u10_u5_n106 ) , .A2( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n119 ) );
  NAND2_X1 u2_u10_u5_U62 (.A2( u2_u10_u5_n103 ) , .A1( u2_u10_u5_n105 ) , .ZN( u2_u10_u5_n140 ) );
  NAND2_X1 u2_u10_u5_U63 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n105 ) , .ZN( u2_u10_u5_n155 ) );
  NAND2_X1 u2_u10_u5_U64 (.A2( u2_u10_u5_n106 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n122 ) );
  NAND2_X1 u2_u10_u5_U65 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n106 ) , .ZN( u2_u10_u5_n115 ) );
  NAND2_X1 u2_u10_u5_U66 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n103 ) , .ZN( u2_u10_u5_n161 ) );
  NAND2_X1 u2_u10_u5_U67 (.A1( u2_u10_u5_n105 ) , .A2( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n154 ) );
  INV_X1 u2_u10_u5_U68 (.A( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n172 ) );
  NAND2_X1 u2_u10_u5_U69 (.A1( u2_u10_u5_n103 ) , .A2( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n123 ) );
  OAI22_X1 u2_u10_u5_U7 (.B2( u2_u10_u5_n149 ) , .B1( u2_u10_u5_n150 ) , .A2( u2_u10_u5_n151 ) , .A1( u2_u10_u5_n152 ) , .ZN( u2_u10_u5_n165 ) );
  NAND2_X1 u2_u10_u5_U70 (.A2( u2_u10_u5_n103 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n151 ) );
  NAND2_X1 u2_u10_u5_U71 (.A2( u2_u10_u5_n107 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n120 ) );
  NAND2_X1 u2_u10_u5_U72 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n157 ) );
  AND2_X1 u2_u10_u5_U73 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n104 ) , .ZN( u2_u10_u5_n131 ) );
  INV_X1 u2_u10_u5_U74 (.A( u2_u10_u5_n102 ) , .ZN( u2_u10_u5_n195 ) );
  OAI221_X1 u2_u10_u5_U75 (.A( u2_u10_u5_n101 ) , .ZN( u2_u10_u5_n102 ) , .C2( u2_u10_u5_n115 ) , .C1( u2_u10_u5_n126 ) , .B1( u2_u10_u5_n134 ) , .B2( u2_u10_u5_n160 ) );
  OAI21_X1 u2_u10_u5_U76 (.ZN( u2_u10_u5_n101 ) , .B1( u2_u10_u5_n137 ) , .A( u2_u10_u5_n146 ) , .B2( u2_u10_u5_n147 ) );
  NOR2_X1 u2_u10_u5_U77 (.A2( u2_u10_X_34 ) , .A1( u2_u10_X_35 ) , .ZN( u2_u10_u5_n145 ) );
  NOR2_X1 u2_u10_u5_U78 (.A2( u2_u10_X_34 ) , .ZN( u2_u10_u5_n146 ) , .A1( u2_u10_u5_n171 ) );
  NOR2_X1 u2_u10_u5_U79 (.A2( u2_u10_X_31 ) , .A1( u2_u10_X_32 ) , .ZN( u2_u10_u5_n103 ) );
  NOR3_X1 u2_u10_u5_U8 (.A2( u2_u10_u5_n147 ) , .A1( u2_u10_u5_n148 ) , .ZN( u2_u10_u5_n149 ) , .A3( u2_u10_u5_n194 ) );
  NOR2_X1 u2_u10_u5_U80 (.A2( u2_u10_X_36 ) , .ZN( u2_u10_u5_n105 ) , .A1( u2_u10_u5_n180 ) );
  NOR2_X1 u2_u10_u5_U81 (.A2( u2_u10_X_33 ) , .ZN( u2_u10_u5_n108 ) , .A1( u2_u10_u5_n170 ) );
  NOR2_X1 u2_u10_u5_U82 (.A2( u2_u10_X_33 ) , .A1( u2_u10_X_36 ) , .ZN( u2_u10_u5_n107 ) );
  NOR2_X1 u2_u10_u5_U83 (.A2( u2_u10_X_31 ) , .ZN( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n181 ) );
  NAND2_X1 u2_u10_u5_U84 (.A2( u2_u10_X_34 ) , .A1( u2_u10_X_35 ) , .ZN( u2_u10_u5_n153 ) );
  NAND2_X1 u2_u10_u5_U85 (.A1( u2_u10_X_34 ) , .ZN( u2_u10_u5_n126 ) , .A2( u2_u10_u5_n171 ) );
  AND2_X1 u2_u10_u5_U86 (.A1( u2_u10_X_31 ) , .A2( u2_u10_X_32 ) , .ZN( u2_u10_u5_n106 ) );
  AND2_X1 u2_u10_u5_U87 (.A1( u2_u10_X_31 ) , .ZN( u2_u10_u5_n109 ) , .A2( u2_u10_u5_n181 ) );
  INV_X1 u2_u10_u5_U88 (.A( u2_u10_X_33 ) , .ZN( u2_u10_u5_n180 ) );
  INV_X1 u2_u10_u5_U89 (.A( u2_u10_X_35 ) , .ZN( u2_u10_u5_n171 ) );
  NOR2_X1 u2_u10_u5_U9 (.ZN( u2_u10_u5_n135 ) , .A1( u2_u10_u5_n173 ) , .A2( u2_u10_u5_n176 ) );
  INV_X1 u2_u10_u5_U90 (.A( u2_u10_X_36 ) , .ZN( u2_u10_u5_n170 ) );
  INV_X1 u2_u10_u5_U91 (.A( u2_u10_X_32 ) , .ZN( u2_u10_u5_n181 ) );
  NAND4_X1 u2_u10_u5_U92 (.ZN( u2_out10_29 ) , .A4( u2_u10_u5_n129 ) , .A3( u2_u10_u5_n130 ) , .A2( u2_u10_u5_n168 ) , .A1( u2_u10_u5_n196 ) );
  AOI221_X1 u2_u10_u5_U93 (.A( u2_u10_u5_n128 ) , .ZN( u2_u10_u5_n129 ) , .C2( u2_u10_u5_n132 ) , .B2( u2_u10_u5_n159 ) , .B1( u2_u10_u5_n176 ) , .C1( u2_u10_u5_n184 ) );
  AOI222_X1 u2_u10_u5_U94 (.ZN( u2_u10_u5_n130 ) , .A2( u2_u10_u5_n146 ) , .B1( u2_u10_u5_n147 ) , .C2( u2_u10_u5_n175 ) , .B2( u2_u10_u5_n179 ) , .A1( u2_u10_u5_n188 ) , .C1( u2_u10_u5_n194 ) );
  NAND4_X1 u2_u10_u5_U95 (.ZN( u2_out10_19 ) , .A4( u2_u10_u5_n166 ) , .A3( u2_u10_u5_n167 ) , .A2( u2_u10_u5_n168 ) , .A1( u2_u10_u5_n169 ) );
  AOI22_X1 u2_u10_u5_U96 (.B2( u2_u10_u5_n145 ) , .A2( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n167 ) , .B1( u2_u10_u5_n182 ) , .A1( u2_u10_u5_n189 ) );
  NOR4_X1 u2_u10_u5_U97 (.A4( u2_u10_u5_n162 ) , .A3( u2_u10_u5_n163 ) , .A2( u2_u10_u5_n164 ) , .A1( u2_u10_u5_n165 ) , .ZN( u2_u10_u5_n166 ) );
  NAND4_X1 u2_u10_u5_U98 (.ZN( u2_out10_11 ) , .A4( u2_u10_u5_n143 ) , .A3( u2_u10_u5_n144 ) , .A2( u2_u10_u5_n169 ) , .A1( u2_u10_u5_n196 ) );
  AOI22_X1 u2_u10_u5_U99 (.A2( u2_u10_u5_n132 ) , .ZN( u2_u10_u5_n144 ) , .B2( u2_u10_u5_n145 ) , .B1( u2_u10_u5_n184 ) , .A1( u2_u10_u5_n194 ) );
  AOI22_X1 u2_u10_u6_U10 (.A2( u2_u10_u6_n151 ) , .B2( u2_u10_u6_n161 ) , .A1( u2_u10_u6_n167 ) , .B1( u2_u10_u6_n170 ) , .ZN( u2_u10_u6_n89 ) );
  AOI21_X1 u2_u10_u6_U11 (.B1( u2_u10_u6_n107 ) , .B2( u2_u10_u6_n132 ) , .A( u2_u10_u6_n158 ) , .ZN( u2_u10_u6_n88 ) );
  AOI21_X1 u2_u10_u6_U12 (.B2( u2_u10_u6_n147 ) , .B1( u2_u10_u6_n148 ) , .ZN( u2_u10_u6_n149 ) , .A( u2_u10_u6_n158 ) );
  AOI21_X1 u2_u10_u6_U13 (.ZN( u2_u10_u6_n106 ) , .A( u2_u10_u6_n142 ) , .B2( u2_u10_u6_n159 ) , .B1( u2_u10_u6_n164 ) );
  INV_X1 u2_u10_u6_U14 (.A( u2_u10_u6_n155 ) , .ZN( u2_u10_u6_n161 ) );
  INV_X1 u2_u10_u6_U15 (.A( u2_u10_u6_n128 ) , .ZN( u2_u10_u6_n164 ) );
  NAND2_X1 u2_u10_u6_U16 (.ZN( u2_u10_u6_n110 ) , .A1( u2_u10_u6_n122 ) , .A2( u2_u10_u6_n129 ) );
  NAND2_X1 u2_u10_u6_U17 (.ZN( u2_u10_u6_n124 ) , .A2( u2_u10_u6_n146 ) , .A1( u2_u10_u6_n148 ) );
  INV_X1 u2_u10_u6_U18 (.A( u2_u10_u6_n132 ) , .ZN( u2_u10_u6_n171 ) );
  AND2_X1 u2_u10_u6_U19 (.A1( u2_u10_u6_n100 ) , .ZN( u2_u10_u6_n130 ) , .A2( u2_u10_u6_n147 ) );
  INV_X1 u2_u10_u6_U20 (.A( u2_u10_u6_n127 ) , .ZN( u2_u10_u6_n173 ) );
  INV_X1 u2_u10_u6_U21 (.A( u2_u10_u6_n121 ) , .ZN( u2_u10_u6_n167 ) );
  INV_X1 u2_u10_u6_U22 (.A( u2_u10_u6_n100 ) , .ZN( u2_u10_u6_n169 ) );
  INV_X1 u2_u10_u6_U23 (.A( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n170 ) );
  INV_X1 u2_u10_u6_U24 (.A( u2_u10_u6_n113 ) , .ZN( u2_u10_u6_n168 ) );
  AND2_X1 u2_u10_u6_U25 (.A1( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n119 ) , .ZN( u2_u10_u6_n133 ) );
  AND2_X1 u2_u10_u6_U26 (.A2( u2_u10_u6_n121 ) , .A1( u2_u10_u6_n122 ) , .ZN( u2_u10_u6_n131 ) );
  AND3_X1 u2_u10_u6_U27 (.ZN( u2_u10_u6_n120 ) , .A2( u2_u10_u6_n127 ) , .A1( u2_u10_u6_n132 ) , .A3( u2_u10_u6_n145 ) );
  INV_X1 u2_u10_u6_U28 (.A( u2_u10_u6_n146 ) , .ZN( u2_u10_u6_n163 ) );
  AOI222_X1 u2_u10_u6_U29 (.ZN( u2_u10_u6_n114 ) , .A1( u2_u10_u6_n118 ) , .A2( u2_u10_u6_n126 ) , .B2( u2_u10_u6_n151 ) , .C2( u2_u10_u6_n159 ) , .C1( u2_u10_u6_n168 ) , .B1( u2_u10_u6_n169 ) );
  INV_X1 u2_u10_u6_U3 (.A( u2_u10_u6_n110 ) , .ZN( u2_u10_u6_n166 ) );
  NOR2_X1 u2_u10_u6_U30 (.A1( u2_u10_u6_n162 ) , .A2( u2_u10_u6_n165 ) , .ZN( u2_u10_u6_n98 ) );
  AOI211_X1 u2_u10_u6_U31 (.B( u2_u10_u6_n134 ) , .A( u2_u10_u6_n135 ) , .C1( u2_u10_u6_n136 ) , .ZN( u2_u10_u6_n137 ) , .C2( u2_u10_u6_n151 ) );
  NAND4_X1 u2_u10_u6_U32 (.A4( u2_u10_u6_n127 ) , .A3( u2_u10_u6_n128 ) , .A2( u2_u10_u6_n129 ) , .A1( u2_u10_u6_n130 ) , .ZN( u2_u10_u6_n136 ) );
  AOI21_X1 u2_u10_u6_U33 (.B2( u2_u10_u6_n132 ) , .B1( u2_u10_u6_n133 ) , .ZN( u2_u10_u6_n134 ) , .A( u2_u10_u6_n158 ) );
  AOI21_X1 u2_u10_u6_U34 (.B1( u2_u10_u6_n131 ) , .ZN( u2_u10_u6_n135 ) , .A( u2_u10_u6_n144 ) , .B2( u2_u10_u6_n146 ) );
  NAND2_X1 u2_u10_u6_U35 (.A1( u2_u10_u6_n144 ) , .ZN( u2_u10_u6_n151 ) , .A2( u2_u10_u6_n158 ) );
  NAND2_X1 u2_u10_u6_U36 (.ZN( u2_u10_u6_n132 ) , .A1( u2_u10_u6_n91 ) , .A2( u2_u10_u6_n97 ) );
  AOI22_X1 u2_u10_u6_U37 (.B2( u2_u10_u6_n110 ) , .B1( u2_u10_u6_n111 ) , .A1( u2_u10_u6_n112 ) , .ZN( u2_u10_u6_n115 ) , .A2( u2_u10_u6_n161 ) );
  NAND4_X1 u2_u10_u6_U38 (.A3( u2_u10_u6_n109 ) , .ZN( u2_u10_u6_n112 ) , .A4( u2_u10_u6_n132 ) , .A2( u2_u10_u6_n147 ) , .A1( u2_u10_u6_n166 ) );
  NOR2_X1 u2_u10_u6_U39 (.ZN( u2_u10_u6_n109 ) , .A1( u2_u10_u6_n170 ) , .A2( u2_u10_u6_n173 ) );
  INV_X1 u2_u10_u6_U4 (.A( u2_u10_u6_n142 ) , .ZN( u2_u10_u6_n174 ) );
  NOR2_X1 u2_u10_u6_U40 (.A2( u2_u10_u6_n126 ) , .ZN( u2_u10_u6_n155 ) , .A1( u2_u10_u6_n160 ) );
  NAND2_X1 u2_u10_u6_U41 (.ZN( u2_u10_u6_n146 ) , .A2( u2_u10_u6_n94 ) , .A1( u2_u10_u6_n99 ) );
  AOI21_X1 u2_u10_u6_U42 (.A( u2_u10_u6_n144 ) , .B2( u2_u10_u6_n145 ) , .B1( u2_u10_u6_n146 ) , .ZN( u2_u10_u6_n150 ) );
  INV_X1 u2_u10_u6_U43 (.A( u2_u10_u6_n111 ) , .ZN( u2_u10_u6_n158 ) );
  NAND2_X1 u2_u10_u6_U44 (.ZN( u2_u10_u6_n127 ) , .A1( u2_u10_u6_n91 ) , .A2( u2_u10_u6_n92 ) );
  NAND2_X1 u2_u10_u6_U45 (.ZN( u2_u10_u6_n129 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n96 ) );
  INV_X1 u2_u10_u6_U46 (.A( u2_u10_u6_n144 ) , .ZN( u2_u10_u6_n159 ) );
  NAND2_X1 u2_u10_u6_U47 (.ZN( u2_u10_u6_n145 ) , .A2( u2_u10_u6_n97 ) , .A1( u2_u10_u6_n98 ) );
  NAND2_X1 u2_u10_u6_U48 (.ZN( u2_u10_u6_n148 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n94 ) );
  NAND2_X1 u2_u10_u6_U49 (.ZN( u2_u10_u6_n108 ) , .A2( u2_u10_u6_n139 ) , .A1( u2_u10_u6_n144 ) );
  NAND2_X1 u2_u10_u6_U5 (.A2( u2_u10_u6_n143 ) , .ZN( u2_u10_u6_n152 ) , .A1( u2_u10_u6_n166 ) );
  NAND2_X1 u2_u10_u6_U50 (.ZN( u2_u10_u6_n121 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n97 ) );
  NAND2_X1 u2_u10_u6_U51 (.ZN( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n95 ) );
  AND2_X1 u2_u10_u6_U52 (.ZN( u2_u10_u6_n118 ) , .A2( u2_u10_u6_n91 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U53 (.ZN( u2_u10_u6_n147 ) , .A2( u2_u10_u6_n98 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U54 (.ZN( u2_u10_u6_n128 ) , .A1( u2_u10_u6_n94 ) , .A2( u2_u10_u6_n96 ) );
  NAND2_X1 u2_u10_u6_U55 (.ZN( u2_u10_u6_n119 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U56 (.ZN( u2_u10_u6_n123 ) , .A2( u2_u10_u6_n91 ) , .A1( u2_u10_u6_n96 ) );
  NAND2_X1 u2_u10_u6_U57 (.ZN( u2_u10_u6_n100 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n98 ) );
  NAND2_X1 u2_u10_u6_U58 (.ZN( u2_u10_u6_n122 ) , .A1( u2_u10_u6_n94 ) , .A2( u2_u10_u6_n97 ) );
  INV_X1 u2_u10_u6_U59 (.A( u2_u10_u6_n139 ) , .ZN( u2_u10_u6_n160 ) );
  AOI22_X1 u2_u10_u6_U6 (.B2( u2_u10_u6_n101 ) , .A1( u2_u10_u6_n102 ) , .ZN( u2_u10_u6_n103 ) , .B1( u2_u10_u6_n160 ) , .A2( u2_u10_u6_n161 ) );
  NAND2_X1 u2_u10_u6_U60 (.ZN( u2_u10_u6_n113 ) , .A1( u2_u10_u6_n96 ) , .A2( u2_u10_u6_n98 ) );
  NOR2_X1 u2_u10_u6_U61 (.A2( u2_u10_X_40 ) , .A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n126 ) );
  NOR2_X1 u2_u10_u6_U62 (.A2( u2_u10_X_39 ) , .A1( u2_u10_X_42 ) , .ZN( u2_u10_u6_n92 ) );
  NOR2_X1 u2_u10_u6_U63 (.A2( u2_u10_X_39 ) , .A1( u2_u10_u6_n156 ) , .ZN( u2_u10_u6_n97 ) );
  NOR2_X1 u2_u10_u6_U64 (.A2( u2_u10_X_38 ) , .A1( u2_u10_u6_n165 ) , .ZN( u2_u10_u6_n95 ) );
  NOR2_X1 u2_u10_u6_U65 (.A2( u2_u10_X_41 ) , .ZN( u2_u10_u6_n111 ) , .A1( u2_u10_u6_n157 ) );
  NOR2_X1 u2_u10_u6_U66 (.A2( u2_u10_X_37 ) , .A1( u2_u10_u6_n162 ) , .ZN( u2_u10_u6_n94 ) );
  NOR2_X1 u2_u10_u6_U67 (.A2( u2_u10_X_37 ) , .A1( u2_u10_X_38 ) , .ZN( u2_u10_u6_n91 ) );
  NAND2_X1 u2_u10_u6_U68 (.A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n144 ) , .A2( u2_u10_u6_n157 ) );
  NAND2_X1 u2_u10_u6_U69 (.A2( u2_u10_X_40 ) , .A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n139 ) );
  NOR2_X1 u2_u10_u6_U7 (.A1( u2_u10_u6_n118 ) , .ZN( u2_u10_u6_n143 ) , .A2( u2_u10_u6_n168 ) );
  AND2_X1 u2_u10_u6_U70 (.A1( u2_u10_X_39 ) , .A2( u2_u10_u6_n156 ) , .ZN( u2_u10_u6_n96 ) );
  AND2_X1 u2_u10_u6_U71 (.A1( u2_u10_X_39 ) , .A2( u2_u10_X_42 ) , .ZN( u2_u10_u6_n99 ) );
  INV_X1 u2_u10_u6_U72 (.A( u2_u10_X_40 ) , .ZN( u2_u10_u6_n157 ) );
  INV_X1 u2_u10_u6_U73 (.A( u2_u10_X_37 ) , .ZN( u2_u10_u6_n165 ) );
  INV_X1 u2_u10_u6_U74 (.A( u2_u10_X_38 ) , .ZN( u2_u10_u6_n162 ) );
  INV_X1 u2_u10_u6_U75 (.A( u2_u10_X_42 ) , .ZN( u2_u10_u6_n156 ) );
  NAND4_X1 u2_u10_u6_U76 (.ZN( u2_out10_12 ) , .A4( u2_u10_u6_n114 ) , .A3( u2_u10_u6_n115 ) , .A2( u2_u10_u6_n116 ) , .A1( u2_u10_u6_n117 ) );
  OAI22_X1 u2_u10_u6_U77 (.B2( u2_u10_u6_n111 ) , .ZN( u2_u10_u6_n116 ) , .B1( u2_u10_u6_n126 ) , .A2( u2_u10_u6_n164 ) , .A1( u2_u10_u6_n167 ) );
  OAI21_X1 u2_u10_u6_U78 (.A( u2_u10_u6_n108 ) , .ZN( u2_u10_u6_n117 ) , .B2( u2_u10_u6_n141 ) , .B1( u2_u10_u6_n163 ) );
  NAND4_X1 u2_u10_u6_U79 (.ZN( u2_out10_32 ) , .A4( u2_u10_u6_n103 ) , .A3( u2_u10_u6_n104 ) , .A2( u2_u10_u6_n105 ) , .A1( u2_u10_u6_n106 ) );
  INV_X1 u2_u10_u6_U8 (.ZN( u2_u10_u6_n172 ) , .A( u2_u10_u6_n88 ) );
  AOI22_X1 u2_u10_u6_U80 (.ZN( u2_u10_u6_n105 ) , .A2( u2_u10_u6_n108 ) , .A1( u2_u10_u6_n118 ) , .B2( u2_u10_u6_n126 ) , .B1( u2_u10_u6_n171 ) );
  AOI22_X1 u2_u10_u6_U81 (.ZN( u2_u10_u6_n104 ) , .A1( u2_u10_u6_n111 ) , .B1( u2_u10_u6_n124 ) , .B2( u2_u10_u6_n151 ) , .A2( u2_u10_u6_n93 ) );
  OAI211_X1 u2_u10_u6_U82 (.ZN( u2_out10_7 ) , .B( u2_u10_u6_n153 ) , .C2( u2_u10_u6_n154 ) , .C1( u2_u10_u6_n155 ) , .A( u2_u10_u6_n174 ) );
  NOR3_X1 u2_u10_u6_U83 (.A1( u2_u10_u6_n141 ) , .ZN( u2_u10_u6_n154 ) , .A3( u2_u10_u6_n164 ) , .A2( u2_u10_u6_n171 ) );
  AOI211_X1 u2_u10_u6_U84 (.B( u2_u10_u6_n149 ) , .A( u2_u10_u6_n150 ) , .C2( u2_u10_u6_n151 ) , .C1( u2_u10_u6_n152 ) , .ZN( u2_u10_u6_n153 ) );
  OAI211_X1 u2_u10_u6_U85 (.ZN( u2_out10_22 ) , .B( u2_u10_u6_n137 ) , .A( u2_u10_u6_n138 ) , .C2( u2_u10_u6_n139 ) , .C1( u2_u10_u6_n140 ) );
  AOI22_X1 u2_u10_u6_U86 (.B1( u2_u10_u6_n124 ) , .A2( u2_u10_u6_n125 ) , .A1( u2_u10_u6_n126 ) , .ZN( u2_u10_u6_n138 ) , .B2( u2_u10_u6_n161 ) );
  AND4_X1 u2_u10_u6_U87 (.A3( u2_u10_u6_n119 ) , .A1( u2_u10_u6_n120 ) , .A4( u2_u10_u6_n129 ) , .ZN( u2_u10_u6_n140 ) , .A2( u2_u10_u6_n143 ) );
  NAND3_X1 u2_u10_u6_U88 (.A2( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n125 ) , .A1( u2_u10_u6_n130 ) , .A3( u2_u10_u6_n131 ) );
  NAND3_X1 u2_u10_u6_U89 (.A3( u2_u10_u6_n133 ) , .ZN( u2_u10_u6_n141 ) , .A1( u2_u10_u6_n145 ) , .A2( u2_u10_u6_n148 ) );
  OAI21_X1 u2_u10_u6_U9 (.A( u2_u10_u6_n159 ) , .B1( u2_u10_u6_n169 ) , .B2( u2_u10_u6_n173 ) , .ZN( u2_u10_u6_n90 ) );
  NAND3_X1 u2_u10_u6_U90 (.ZN( u2_u10_u6_n101 ) , .A3( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n121 ) , .A1( u2_u10_u6_n127 ) );
  NAND3_X1 u2_u10_u6_U91 (.ZN( u2_u10_u6_n102 ) , .A3( u2_u10_u6_n130 ) , .A2( u2_u10_u6_n145 ) , .A1( u2_u10_u6_n166 ) );
  NAND3_X1 u2_u10_u6_U92 (.A3( u2_u10_u6_n113 ) , .A1( u2_u10_u6_n119 ) , .A2( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n93 ) );
  NAND3_X1 u2_u10_u6_U93 (.ZN( u2_u10_u6_n142 ) , .A2( u2_u10_u6_n172 ) , .A3( u2_u10_u6_n89 ) , .A1( u2_u10_u6_n90 ) );
  XOR2_X1 u2_u11_U10 (.B( u2_K12_45 ) , .A( u2_R10_30 ) , .Z( u2_u11_X_45 ) );
  XOR2_X1 u2_u11_U11 (.B( u2_K12_44 ) , .A( u2_R10_29 ) , .Z( u2_u11_X_44 ) );
  XOR2_X1 u2_u11_U12 (.B( u2_K12_43 ) , .A( u2_R10_28 ) , .Z( u2_u11_X_43 ) );
  XOR2_X1 u2_u11_U13 (.B( u2_K12_42 ) , .A( u2_R10_29 ) , .Z( u2_u11_X_42 ) );
  XOR2_X1 u2_u11_U14 (.B( u2_K12_41 ) , .A( u2_R10_28 ) , .Z( u2_u11_X_41 ) );
  XOR2_X1 u2_u11_U15 (.B( u2_K12_40 ) , .A( u2_R10_27 ) , .Z( u2_u11_X_40 ) );
  XOR2_X1 u2_u11_U17 (.B( u2_K12_39 ) , .A( u2_R10_26 ) , .Z( u2_u11_X_39 ) );
  XOR2_X1 u2_u11_U18 (.B( u2_K12_38 ) , .A( u2_R10_25 ) , .Z( u2_u11_X_38 ) );
  XOR2_X1 u2_u11_U19 (.B( u2_K12_37 ) , .A( u2_R10_24 ) , .Z( u2_u11_X_37 ) );
  XOR2_X1 u2_u11_U20 (.B( u2_K12_36 ) , .A( u2_R10_25 ) , .Z( u2_u11_X_36 ) );
  XOR2_X1 u2_u11_U21 (.B( u2_K12_35 ) , .A( u2_R10_24 ) , .Z( u2_u11_X_35 ) );
  XOR2_X1 u2_u11_U22 (.B( u2_K12_34 ) , .A( u2_R10_23 ) , .Z( u2_u11_X_34 ) );
  XOR2_X1 u2_u11_U23 (.B( u2_K12_33 ) , .A( u2_R10_22 ) , .Z( u2_u11_X_33 ) );
  XOR2_X1 u2_u11_U24 (.B( u2_K12_32 ) , .A( u2_R10_21 ) , .Z( u2_u11_X_32 ) );
  XOR2_X1 u2_u11_U25 (.B( u2_K12_31 ) , .A( u2_R10_20 ) , .Z( u2_u11_X_31 ) );
  XOR2_X1 u2_u11_U26 (.B( u2_K12_30 ) , .A( u2_R10_21 ) , .Z( u2_u11_X_30 ) );
  XOR2_X1 u2_u11_U28 (.B( u2_K12_29 ) , .A( u2_R10_20 ) , .Z( u2_u11_X_29 ) );
  XOR2_X1 u2_u11_U29 (.B( u2_K12_28 ) , .A( u2_R10_19 ) , .Z( u2_u11_X_28 ) );
  XOR2_X1 u2_u11_U30 (.B( u2_K12_27 ) , .A( u2_R10_18 ) , .Z( u2_u11_X_27 ) );
  XOR2_X1 u2_u11_U31 (.B( u2_K12_26 ) , .A( u2_R10_17 ) , .Z( u2_u11_X_26 ) );
  XOR2_X1 u2_u11_U32 (.B( u2_K12_25 ) , .A( u2_R10_16 ) , .Z( u2_u11_X_25 ) );
  XOR2_X1 u2_u11_U7 (.B( u2_K12_48 ) , .A( u2_R10_1 ) , .Z( u2_u11_X_48 ) );
  XOR2_X1 u2_u11_U8 (.B( u2_K12_47 ) , .A( u2_R10_32 ) , .Z( u2_u11_X_47 ) );
  XOR2_X1 u2_u11_U9 (.B( u2_K12_46 ) , .A( u2_R10_31 ) , .Z( u2_u11_X_46 ) );
  OAI22_X1 u2_u11_u4_U10 (.B2( u2_u11_u4_n135 ) , .ZN( u2_u11_u4_n137 ) , .B1( u2_u11_u4_n153 ) , .A1( u2_u11_u4_n155 ) , .A2( u2_u11_u4_n171 ) );
  AND3_X1 u2_u11_u4_U11 (.A2( u2_u11_u4_n134 ) , .ZN( u2_u11_u4_n135 ) , .A3( u2_u11_u4_n145 ) , .A1( u2_u11_u4_n157 ) );
  NAND2_X1 u2_u11_u4_U12 (.ZN( u2_u11_u4_n132 ) , .A2( u2_u11_u4_n170 ) , .A1( u2_u11_u4_n173 ) );
  AOI21_X1 u2_u11_u4_U13 (.B2( u2_u11_u4_n160 ) , .B1( u2_u11_u4_n161 ) , .ZN( u2_u11_u4_n162 ) , .A( u2_u11_u4_n170 ) );
  AOI21_X1 u2_u11_u4_U14 (.ZN( u2_u11_u4_n107 ) , .B2( u2_u11_u4_n143 ) , .A( u2_u11_u4_n174 ) , .B1( u2_u11_u4_n184 ) );
  AOI21_X1 u2_u11_u4_U15 (.B2( u2_u11_u4_n158 ) , .B1( u2_u11_u4_n159 ) , .ZN( u2_u11_u4_n163 ) , .A( u2_u11_u4_n174 ) );
  AOI21_X1 u2_u11_u4_U16 (.A( u2_u11_u4_n153 ) , .B2( u2_u11_u4_n154 ) , .B1( u2_u11_u4_n155 ) , .ZN( u2_u11_u4_n165 ) );
  AOI21_X1 u2_u11_u4_U17 (.A( u2_u11_u4_n156 ) , .B2( u2_u11_u4_n157 ) , .ZN( u2_u11_u4_n164 ) , .B1( u2_u11_u4_n184 ) );
  INV_X1 u2_u11_u4_U18 (.A( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n170 ) );
  AND2_X1 u2_u11_u4_U19 (.A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n155 ) , .A1( u2_u11_u4_n160 ) );
  INV_X1 u2_u11_u4_U20 (.A( u2_u11_u4_n156 ) , .ZN( u2_u11_u4_n175 ) );
  NAND2_X1 u2_u11_u4_U21 (.A2( u2_u11_u4_n118 ) , .ZN( u2_u11_u4_n131 ) , .A1( u2_u11_u4_n147 ) );
  NAND2_X1 u2_u11_u4_U22 (.A1( u2_u11_u4_n119 ) , .A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n130 ) );
  NAND2_X1 u2_u11_u4_U23 (.ZN( u2_u11_u4_n117 ) , .A2( u2_u11_u4_n118 ) , .A1( u2_u11_u4_n148 ) );
  NAND2_X1 u2_u11_u4_U24 (.ZN( u2_u11_u4_n129 ) , .A1( u2_u11_u4_n134 ) , .A2( u2_u11_u4_n148 ) );
  AND3_X1 u2_u11_u4_U25 (.A1( u2_u11_u4_n119 ) , .A2( u2_u11_u4_n143 ) , .A3( u2_u11_u4_n154 ) , .ZN( u2_u11_u4_n161 ) );
  AND2_X1 u2_u11_u4_U26 (.A1( u2_u11_u4_n145 ) , .A2( u2_u11_u4_n147 ) , .ZN( u2_u11_u4_n159 ) );
  OR3_X1 u2_u11_u4_U27 (.A3( u2_u11_u4_n114 ) , .A2( u2_u11_u4_n115 ) , .A1( u2_u11_u4_n116 ) , .ZN( u2_u11_u4_n136 ) );
  AOI21_X1 u2_u11_u4_U28 (.A( u2_u11_u4_n113 ) , .ZN( u2_u11_u4_n116 ) , .B2( u2_u11_u4_n173 ) , .B1( u2_u11_u4_n174 ) );
  AOI21_X1 u2_u11_u4_U29 (.ZN( u2_u11_u4_n115 ) , .B2( u2_u11_u4_n145 ) , .B1( u2_u11_u4_n146 ) , .A( u2_u11_u4_n156 ) );
  NOR2_X1 u2_u11_u4_U3 (.ZN( u2_u11_u4_n121 ) , .A1( u2_u11_u4_n181 ) , .A2( u2_u11_u4_n182 ) );
  OAI22_X1 u2_u11_u4_U30 (.ZN( u2_u11_u4_n114 ) , .A2( u2_u11_u4_n121 ) , .B1( u2_u11_u4_n160 ) , .B2( u2_u11_u4_n170 ) , .A1( u2_u11_u4_n171 ) );
  INV_X1 u2_u11_u4_U31 (.A( u2_u11_u4_n158 ) , .ZN( u2_u11_u4_n182 ) );
  INV_X1 u2_u11_u4_U32 (.ZN( u2_u11_u4_n181 ) , .A( u2_u11_u4_n96 ) );
  INV_X1 u2_u11_u4_U33 (.A( u2_u11_u4_n144 ) , .ZN( u2_u11_u4_n179 ) );
  INV_X1 u2_u11_u4_U34 (.A( u2_u11_u4_n157 ) , .ZN( u2_u11_u4_n178 ) );
  NAND2_X1 u2_u11_u4_U35 (.A2( u2_u11_u4_n154 ) , .A1( u2_u11_u4_n96 ) , .ZN( u2_u11_u4_n97 ) );
  INV_X1 u2_u11_u4_U36 (.ZN( u2_u11_u4_n186 ) , .A( u2_u11_u4_n95 ) );
  OAI221_X1 u2_u11_u4_U37 (.C1( u2_u11_u4_n134 ) , .B1( u2_u11_u4_n158 ) , .B2( u2_u11_u4_n171 ) , .C2( u2_u11_u4_n173 ) , .A( u2_u11_u4_n94 ) , .ZN( u2_u11_u4_n95 ) );
  AOI222_X1 u2_u11_u4_U38 (.B2( u2_u11_u4_n132 ) , .A1( u2_u11_u4_n138 ) , .C2( u2_u11_u4_n175 ) , .A2( u2_u11_u4_n179 ) , .C1( u2_u11_u4_n181 ) , .B1( u2_u11_u4_n185 ) , .ZN( u2_u11_u4_n94 ) );
  INV_X1 u2_u11_u4_U39 (.A( u2_u11_u4_n113 ) , .ZN( u2_u11_u4_n185 ) );
  INV_X1 u2_u11_u4_U4 (.A( u2_u11_u4_n117 ) , .ZN( u2_u11_u4_n184 ) );
  INV_X1 u2_u11_u4_U40 (.A( u2_u11_u4_n143 ) , .ZN( u2_u11_u4_n183 ) );
  NOR2_X1 u2_u11_u4_U41 (.ZN( u2_u11_u4_n138 ) , .A1( u2_u11_u4_n168 ) , .A2( u2_u11_u4_n169 ) );
  NOR2_X1 u2_u11_u4_U42 (.A1( u2_u11_u4_n150 ) , .A2( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n153 ) );
  NOR2_X1 u2_u11_u4_U43 (.A2( u2_u11_u4_n128 ) , .A1( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n156 ) );
  AOI22_X1 u2_u11_u4_U44 (.B2( u2_u11_u4_n122 ) , .A1( u2_u11_u4_n123 ) , .ZN( u2_u11_u4_n124 ) , .B1( u2_u11_u4_n128 ) , .A2( u2_u11_u4_n172 ) );
  INV_X1 u2_u11_u4_U45 (.A( u2_u11_u4_n153 ) , .ZN( u2_u11_u4_n172 ) );
  NAND2_X1 u2_u11_u4_U46 (.A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n123 ) , .A1( u2_u11_u4_n161 ) );
  AOI22_X1 u2_u11_u4_U47 (.B2( u2_u11_u4_n132 ) , .A2( u2_u11_u4_n133 ) , .ZN( u2_u11_u4_n140 ) , .A1( u2_u11_u4_n150 ) , .B1( u2_u11_u4_n179 ) );
  NAND2_X1 u2_u11_u4_U48 (.ZN( u2_u11_u4_n133 ) , .A2( u2_u11_u4_n146 ) , .A1( u2_u11_u4_n154 ) );
  NAND2_X1 u2_u11_u4_U49 (.A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n154 ) , .A2( u2_u11_u4_n98 ) );
  NOR4_X1 u2_u11_u4_U5 (.A4( u2_u11_u4_n106 ) , .A3( u2_u11_u4_n107 ) , .A2( u2_u11_u4_n108 ) , .A1( u2_u11_u4_n109 ) , .ZN( u2_u11_u4_n110 ) );
  NAND2_X1 u2_u11_u4_U50 (.A1( u2_u11_u4_n101 ) , .ZN( u2_u11_u4_n158 ) , .A2( u2_u11_u4_n99 ) );
  AOI21_X1 u2_u11_u4_U51 (.ZN( u2_u11_u4_n127 ) , .A( u2_u11_u4_n136 ) , .B2( u2_u11_u4_n150 ) , .B1( u2_u11_u4_n180 ) );
  INV_X1 u2_u11_u4_U52 (.A( u2_u11_u4_n160 ) , .ZN( u2_u11_u4_n180 ) );
  NAND2_X1 u2_u11_u4_U53 (.A2( u2_u11_u4_n104 ) , .A1( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n146 ) );
  NAND2_X1 u2_u11_u4_U54 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n160 ) );
  NAND2_X1 u2_u11_u4_U55 (.ZN( u2_u11_u4_n134 ) , .A1( u2_u11_u4_n98 ) , .A2( u2_u11_u4_n99 ) );
  NAND2_X1 u2_u11_u4_U56 (.A1( u2_u11_u4_n103 ) , .A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n143 ) );
  NAND2_X1 u2_u11_u4_U57 (.A2( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n145 ) , .A1( u2_u11_u4_n98 ) );
  NAND2_X1 u2_u11_u4_U58 (.A1( u2_u11_u4_n100 ) , .A2( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n120 ) );
  NAND2_X1 u2_u11_u4_U59 (.A1( u2_u11_u4_n102 ) , .A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n148 ) );
  AOI21_X1 u2_u11_u4_U6 (.ZN( u2_u11_u4_n106 ) , .B2( u2_u11_u4_n146 ) , .B1( u2_u11_u4_n158 ) , .A( u2_u11_u4_n170 ) );
  NAND2_X1 u2_u11_u4_U60 (.A2( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n157 ) );
  INV_X1 u2_u11_u4_U61 (.A( u2_u11_u4_n150 ) , .ZN( u2_u11_u4_n173 ) );
  INV_X1 u2_u11_u4_U62 (.A( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n171 ) );
  NAND2_X1 u2_u11_u4_U63 (.A1( u2_u11_u4_n100 ) , .ZN( u2_u11_u4_n118 ) , .A2( u2_u11_u4_n99 ) );
  NAND2_X1 u2_u11_u4_U64 (.A2( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n144 ) );
  NAND2_X1 u2_u11_u4_U65 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n96 ) );
  INV_X1 u2_u11_u4_U66 (.A( u2_u11_u4_n128 ) , .ZN( u2_u11_u4_n174 ) );
  NAND2_X1 u2_u11_u4_U67 (.A2( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n119 ) , .A1( u2_u11_u4_n98 ) );
  NAND2_X1 u2_u11_u4_U68 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n147 ) );
  NAND2_X1 u2_u11_u4_U69 (.A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n113 ) , .A1( u2_u11_u4_n99 ) );
  AOI21_X1 u2_u11_u4_U7 (.ZN( u2_u11_u4_n108 ) , .B2( u2_u11_u4_n134 ) , .B1( u2_u11_u4_n155 ) , .A( u2_u11_u4_n156 ) );
  NOR2_X1 u2_u11_u4_U70 (.A2( u2_u11_X_28 ) , .ZN( u2_u11_u4_n150 ) , .A1( u2_u11_u4_n168 ) );
  NOR2_X1 u2_u11_u4_U71 (.A2( u2_u11_X_29 ) , .ZN( u2_u11_u4_n152 ) , .A1( u2_u11_u4_n169 ) );
  NOR2_X1 u2_u11_u4_U72 (.A2( u2_u11_X_26 ) , .ZN( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n177 ) );
  NOR2_X1 u2_u11_u4_U73 (.A2( u2_u11_X_30 ) , .ZN( u2_u11_u4_n105 ) , .A1( u2_u11_u4_n176 ) );
  NOR2_X1 u2_u11_u4_U74 (.A2( u2_u11_X_28 ) , .A1( u2_u11_X_29 ) , .ZN( u2_u11_u4_n128 ) );
  NOR2_X1 u2_u11_u4_U75 (.A2( u2_u11_X_25 ) , .A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n98 ) );
  NOR2_X1 u2_u11_u4_U76 (.A2( u2_u11_X_27 ) , .A1( u2_u11_X_30 ) , .ZN( u2_u11_u4_n102 ) );
  AND2_X1 u2_u11_u4_U77 (.A2( u2_u11_X_25 ) , .A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n104 ) );
  AND2_X1 u2_u11_u4_U78 (.A1( u2_u11_X_30 ) , .A2( u2_u11_u4_n176 ) , .ZN( u2_u11_u4_n99 ) );
  AND2_X1 u2_u11_u4_U79 (.A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n101 ) , .A2( u2_u11_u4_n177 ) );
  AOI21_X1 u2_u11_u4_U8 (.ZN( u2_u11_u4_n109 ) , .A( u2_u11_u4_n153 ) , .B1( u2_u11_u4_n159 ) , .B2( u2_u11_u4_n184 ) );
  AND2_X1 u2_u11_u4_U80 (.A1( u2_u11_X_27 ) , .A2( u2_u11_X_30 ) , .ZN( u2_u11_u4_n103 ) );
  INV_X1 u2_u11_u4_U81 (.A( u2_u11_X_28 ) , .ZN( u2_u11_u4_n169 ) );
  INV_X1 u2_u11_u4_U82 (.A( u2_u11_X_29 ) , .ZN( u2_u11_u4_n168 ) );
  INV_X1 u2_u11_u4_U83 (.A( u2_u11_X_25 ) , .ZN( u2_u11_u4_n177 ) );
  INV_X1 u2_u11_u4_U84 (.A( u2_u11_X_27 ) , .ZN( u2_u11_u4_n176 ) );
  NAND4_X1 u2_u11_u4_U85 (.ZN( u2_out11_25 ) , .A4( u2_u11_u4_n139 ) , .A3( u2_u11_u4_n140 ) , .A2( u2_u11_u4_n141 ) , .A1( u2_u11_u4_n142 ) );
  OAI21_X1 u2_u11_u4_U86 (.A( u2_u11_u4_n128 ) , .B2( u2_u11_u4_n129 ) , .B1( u2_u11_u4_n130 ) , .ZN( u2_u11_u4_n142 ) );
  OAI21_X1 u2_u11_u4_U87 (.B2( u2_u11_u4_n131 ) , .ZN( u2_u11_u4_n141 ) , .A( u2_u11_u4_n175 ) , .B1( u2_u11_u4_n183 ) );
  NAND4_X1 u2_u11_u4_U88 (.ZN( u2_out11_14 ) , .A4( u2_u11_u4_n124 ) , .A3( u2_u11_u4_n125 ) , .A2( u2_u11_u4_n126 ) , .A1( u2_u11_u4_n127 ) );
  AOI22_X1 u2_u11_u4_U89 (.B2( u2_u11_u4_n117 ) , .ZN( u2_u11_u4_n126 ) , .A1( u2_u11_u4_n129 ) , .B1( u2_u11_u4_n152 ) , .A2( u2_u11_u4_n175 ) );
  AOI211_X1 u2_u11_u4_U9 (.B( u2_u11_u4_n136 ) , .A( u2_u11_u4_n137 ) , .C2( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n139 ) , .C1( u2_u11_u4_n182 ) );
  AOI22_X1 u2_u11_u4_U90 (.ZN( u2_u11_u4_n125 ) , .B2( u2_u11_u4_n131 ) , .A2( u2_u11_u4_n132 ) , .B1( u2_u11_u4_n138 ) , .A1( u2_u11_u4_n178 ) );
  NAND4_X1 u2_u11_u4_U91 (.ZN( u2_out11_8 ) , .A4( u2_u11_u4_n110 ) , .A3( u2_u11_u4_n111 ) , .A2( u2_u11_u4_n112 ) , .A1( u2_u11_u4_n186 ) );
  NAND2_X1 u2_u11_u4_U92 (.ZN( u2_u11_u4_n112 ) , .A2( u2_u11_u4_n130 ) , .A1( u2_u11_u4_n150 ) );
  AOI22_X1 u2_u11_u4_U93 (.ZN( u2_u11_u4_n111 ) , .B2( u2_u11_u4_n132 ) , .A1( u2_u11_u4_n152 ) , .B1( u2_u11_u4_n178 ) , .A2( u2_u11_u4_n97 ) );
  AOI22_X1 u2_u11_u4_U94 (.B2( u2_u11_u4_n149 ) , .B1( u2_u11_u4_n150 ) , .A2( u2_u11_u4_n151 ) , .A1( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n167 ) );
  NOR4_X1 u2_u11_u4_U95 (.A4( u2_u11_u4_n162 ) , .A3( u2_u11_u4_n163 ) , .A2( u2_u11_u4_n164 ) , .A1( u2_u11_u4_n165 ) , .ZN( u2_u11_u4_n166 ) );
  NAND3_X1 u2_u11_u4_U96 (.ZN( u2_out11_3 ) , .A3( u2_u11_u4_n166 ) , .A1( u2_u11_u4_n167 ) , .A2( u2_u11_u4_n186 ) );
  NAND3_X1 u2_u11_u4_U97 (.A3( u2_u11_u4_n146 ) , .A2( u2_u11_u4_n147 ) , .A1( u2_u11_u4_n148 ) , .ZN( u2_u11_u4_n149 ) );
  NAND3_X1 u2_u11_u4_U98 (.A3( u2_u11_u4_n143 ) , .A2( u2_u11_u4_n144 ) , .A1( u2_u11_u4_n145 ) , .ZN( u2_u11_u4_n151 ) );
  NAND3_X1 u2_u11_u4_U99 (.A3( u2_u11_u4_n121 ) , .ZN( u2_u11_u4_n122 ) , .A2( u2_u11_u4_n144 ) , .A1( u2_u11_u4_n154 ) );
  INV_X1 u2_u11_u5_U10 (.A( u2_u11_u5_n121 ) , .ZN( u2_u11_u5_n177 ) );
  NOR3_X1 u2_u11_u5_U100 (.A3( u2_u11_u5_n141 ) , .A1( u2_u11_u5_n142 ) , .ZN( u2_u11_u5_n143 ) , .A2( u2_u11_u5_n191 ) );
  NAND4_X1 u2_u11_u5_U101 (.ZN( u2_out11_4 ) , .A4( u2_u11_u5_n112 ) , .A2( u2_u11_u5_n113 ) , .A1( u2_u11_u5_n114 ) , .A3( u2_u11_u5_n195 ) );
  AOI211_X1 u2_u11_u5_U102 (.A( u2_u11_u5_n110 ) , .C1( u2_u11_u5_n111 ) , .ZN( u2_u11_u5_n112 ) , .B( u2_u11_u5_n118 ) , .C2( u2_u11_u5_n177 ) );
  AOI222_X1 u2_u11_u5_U103 (.ZN( u2_u11_u5_n113 ) , .A1( u2_u11_u5_n131 ) , .C1( u2_u11_u5_n148 ) , .B2( u2_u11_u5_n174 ) , .C2( u2_u11_u5_n178 ) , .A2( u2_u11_u5_n179 ) , .B1( u2_u11_u5_n99 ) );
  NAND3_X1 u2_u11_u5_U104 (.A2( u2_u11_u5_n154 ) , .A3( u2_u11_u5_n158 ) , .A1( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n99 ) );
  NOR2_X1 u2_u11_u5_U11 (.ZN( u2_u11_u5_n160 ) , .A2( u2_u11_u5_n173 ) , .A1( u2_u11_u5_n177 ) );
  INV_X1 u2_u11_u5_U12 (.A( u2_u11_u5_n150 ) , .ZN( u2_u11_u5_n174 ) );
  AOI21_X1 u2_u11_u5_U13 (.A( u2_u11_u5_n160 ) , .B2( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n162 ) , .B1( u2_u11_u5_n192 ) );
  INV_X1 u2_u11_u5_U14 (.A( u2_u11_u5_n159 ) , .ZN( u2_u11_u5_n192 ) );
  AOI21_X1 u2_u11_u5_U15 (.A( u2_u11_u5_n156 ) , .B2( u2_u11_u5_n157 ) , .B1( u2_u11_u5_n158 ) , .ZN( u2_u11_u5_n163 ) );
  AOI21_X1 u2_u11_u5_U16 (.B2( u2_u11_u5_n139 ) , .B1( u2_u11_u5_n140 ) , .ZN( u2_u11_u5_n141 ) , .A( u2_u11_u5_n150 ) );
  OAI21_X1 u2_u11_u5_U17 (.A( u2_u11_u5_n133 ) , .B2( u2_u11_u5_n134 ) , .B1( u2_u11_u5_n135 ) , .ZN( u2_u11_u5_n142 ) );
  OAI21_X1 u2_u11_u5_U18 (.ZN( u2_u11_u5_n133 ) , .B2( u2_u11_u5_n147 ) , .A( u2_u11_u5_n173 ) , .B1( u2_u11_u5_n188 ) );
  NAND2_X1 u2_u11_u5_U19 (.A2( u2_u11_u5_n119 ) , .A1( u2_u11_u5_n123 ) , .ZN( u2_u11_u5_n137 ) );
  INV_X1 u2_u11_u5_U20 (.A( u2_u11_u5_n155 ) , .ZN( u2_u11_u5_n194 ) );
  NAND2_X1 u2_u11_u5_U21 (.A1( u2_u11_u5_n121 ) , .ZN( u2_u11_u5_n132 ) , .A2( u2_u11_u5_n172 ) );
  NAND2_X1 u2_u11_u5_U22 (.A2( u2_u11_u5_n122 ) , .ZN( u2_u11_u5_n136 ) , .A1( u2_u11_u5_n154 ) );
  NAND2_X1 u2_u11_u5_U23 (.A2( u2_u11_u5_n119 ) , .A1( u2_u11_u5_n120 ) , .ZN( u2_u11_u5_n159 ) );
  INV_X1 u2_u11_u5_U24 (.A( u2_u11_u5_n156 ) , .ZN( u2_u11_u5_n175 ) );
  INV_X1 u2_u11_u5_U25 (.A( u2_u11_u5_n158 ) , .ZN( u2_u11_u5_n188 ) );
  INV_X1 u2_u11_u5_U26 (.A( u2_u11_u5_n152 ) , .ZN( u2_u11_u5_n179 ) );
  INV_X1 u2_u11_u5_U27 (.A( u2_u11_u5_n140 ) , .ZN( u2_u11_u5_n182 ) );
  INV_X1 u2_u11_u5_U28 (.A( u2_u11_u5_n151 ) , .ZN( u2_u11_u5_n183 ) );
  INV_X1 u2_u11_u5_U29 (.A( u2_u11_u5_n123 ) , .ZN( u2_u11_u5_n185 ) );
  NOR2_X1 u2_u11_u5_U3 (.ZN( u2_u11_u5_n134 ) , .A1( u2_u11_u5_n183 ) , .A2( u2_u11_u5_n190 ) );
  INV_X1 u2_u11_u5_U30 (.A( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n184 ) );
  INV_X1 u2_u11_u5_U31 (.A( u2_u11_u5_n139 ) , .ZN( u2_u11_u5_n189 ) );
  INV_X1 u2_u11_u5_U32 (.A( u2_u11_u5_n157 ) , .ZN( u2_u11_u5_n190 ) );
  INV_X1 u2_u11_u5_U33 (.A( u2_u11_u5_n120 ) , .ZN( u2_u11_u5_n193 ) );
  NAND2_X1 u2_u11_u5_U34 (.ZN( u2_u11_u5_n111 ) , .A1( u2_u11_u5_n140 ) , .A2( u2_u11_u5_n155 ) );
  NOR2_X1 u2_u11_u5_U35 (.ZN( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n170 ) , .A2( u2_u11_u5_n180 ) );
  INV_X1 u2_u11_u5_U36 (.A( u2_u11_u5_n117 ) , .ZN( u2_u11_u5_n196 ) );
  OAI221_X1 u2_u11_u5_U37 (.A( u2_u11_u5_n116 ) , .ZN( u2_u11_u5_n117 ) , .B2( u2_u11_u5_n119 ) , .C1( u2_u11_u5_n153 ) , .C2( u2_u11_u5_n158 ) , .B1( u2_u11_u5_n172 ) );
  AOI222_X1 u2_u11_u5_U38 (.ZN( u2_u11_u5_n116 ) , .B2( u2_u11_u5_n145 ) , .C1( u2_u11_u5_n148 ) , .A2( u2_u11_u5_n174 ) , .C2( u2_u11_u5_n177 ) , .B1( u2_u11_u5_n187 ) , .A1( u2_u11_u5_n193 ) );
  INV_X1 u2_u11_u5_U39 (.A( u2_u11_u5_n115 ) , .ZN( u2_u11_u5_n187 ) );
  INV_X1 u2_u11_u5_U4 (.A( u2_u11_u5_n138 ) , .ZN( u2_u11_u5_n191 ) );
  AOI22_X1 u2_u11_u5_U40 (.B2( u2_u11_u5_n131 ) , .A2( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n169 ) , .B1( u2_u11_u5_n174 ) , .A1( u2_u11_u5_n185 ) );
  NOR2_X1 u2_u11_u5_U41 (.A1( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n150 ) , .A2( u2_u11_u5_n173 ) );
  AOI21_X1 u2_u11_u5_U42 (.A( u2_u11_u5_n118 ) , .B2( u2_u11_u5_n145 ) , .ZN( u2_u11_u5_n168 ) , .B1( u2_u11_u5_n186 ) );
  INV_X1 u2_u11_u5_U43 (.A( u2_u11_u5_n122 ) , .ZN( u2_u11_u5_n186 ) );
  NOR2_X1 u2_u11_u5_U44 (.A1( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n152 ) , .A2( u2_u11_u5_n176 ) );
  NOR2_X1 u2_u11_u5_U45 (.A1( u2_u11_u5_n115 ) , .ZN( u2_u11_u5_n118 ) , .A2( u2_u11_u5_n153 ) );
  NOR2_X1 u2_u11_u5_U46 (.A2( u2_u11_u5_n145 ) , .ZN( u2_u11_u5_n156 ) , .A1( u2_u11_u5_n174 ) );
  NOR2_X1 u2_u11_u5_U47 (.ZN( u2_u11_u5_n121 ) , .A2( u2_u11_u5_n145 ) , .A1( u2_u11_u5_n176 ) );
  AOI22_X1 u2_u11_u5_U48 (.ZN( u2_u11_u5_n114 ) , .A2( u2_u11_u5_n137 ) , .A1( u2_u11_u5_n145 ) , .B2( u2_u11_u5_n175 ) , .B1( u2_u11_u5_n193 ) );
  OAI211_X1 u2_u11_u5_U49 (.B( u2_u11_u5_n124 ) , .A( u2_u11_u5_n125 ) , .C2( u2_u11_u5_n126 ) , .C1( u2_u11_u5_n127 ) , .ZN( u2_u11_u5_n128 ) );
  OAI21_X1 u2_u11_u5_U5 (.B2( u2_u11_u5_n136 ) , .B1( u2_u11_u5_n137 ) , .ZN( u2_u11_u5_n138 ) , .A( u2_u11_u5_n177 ) );
  OAI21_X1 u2_u11_u5_U50 (.ZN( u2_u11_u5_n124 ) , .A( u2_u11_u5_n177 ) , .B2( u2_u11_u5_n183 ) , .B1( u2_u11_u5_n189 ) );
  NOR3_X1 u2_u11_u5_U51 (.ZN( u2_u11_u5_n127 ) , .A1( u2_u11_u5_n136 ) , .A3( u2_u11_u5_n148 ) , .A2( u2_u11_u5_n182 ) );
  OAI21_X1 u2_u11_u5_U52 (.ZN( u2_u11_u5_n125 ) , .A( u2_u11_u5_n174 ) , .B2( u2_u11_u5_n185 ) , .B1( u2_u11_u5_n190 ) );
  AOI21_X1 u2_u11_u5_U53 (.A( u2_u11_u5_n153 ) , .B2( u2_u11_u5_n154 ) , .B1( u2_u11_u5_n155 ) , .ZN( u2_u11_u5_n164 ) );
  AOI21_X1 u2_u11_u5_U54 (.ZN( u2_u11_u5_n110 ) , .B1( u2_u11_u5_n122 ) , .B2( u2_u11_u5_n139 ) , .A( u2_u11_u5_n153 ) );
  INV_X1 u2_u11_u5_U55 (.A( u2_u11_u5_n153 ) , .ZN( u2_u11_u5_n176 ) );
  INV_X1 u2_u11_u5_U56 (.A( u2_u11_u5_n126 ) , .ZN( u2_u11_u5_n173 ) );
  AND2_X1 u2_u11_u5_U57 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n147 ) );
  AND2_X1 u2_u11_u5_U58 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n148 ) );
  NAND2_X1 u2_u11_u5_U59 (.A1( u2_u11_u5_n105 ) , .A2( u2_u11_u5_n106 ) , .ZN( u2_u11_u5_n158 ) );
  INV_X1 u2_u11_u5_U6 (.A( u2_u11_u5_n135 ) , .ZN( u2_u11_u5_n178 ) );
  NAND2_X1 u2_u11_u5_U60 (.A2( u2_u11_u5_n108 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n139 ) );
  NAND2_X1 u2_u11_u5_U61 (.A1( u2_u11_u5_n106 ) , .A2( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n119 ) );
  NAND2_X1 u2_u11_u5_U62 (.A2( u2_u11_u5_n103 ) , .A1( u2_u11_u5_n105 ) , .ZN( u2_u11_u5_n140 ) );
  NAND2_X1 u2_u11_u5_U63 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n105 ) , .ZN( u2_u11_u5_n155 ) );
  NAND2_X1 u2_u11_u5_U64 (.A2( u2_u11_u5_n106 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n122 ) );
  NAND2_X1 u2_u11_u5_U65 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n106 ) , .ZN( u2_u11_u5_n115 ) );
  NAND2_X1 u2_u11_u5_U66 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n103 ) , .ZN( u2_u11_u5_n161 ) );
  NAND2_X1 u2_u11_u5_U67 (.A1( u2_u11_u5_n105 ) , .A2( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n154 ) );
  INV_X1 u2_u11_u5_U68 (.A( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n172 ) );
  NAND2_X1 u2_u11_u5_U69 (.A1( u2_u11_u5_n103 ) , .A2( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n123 ) );
  OAI22_X1 u2_u11_u5_U7 (.B2( u2_u11_u5_n149 ) , .B1( u2_u11_u5_n150 ) , .A2( u2_u11_u5_n151 ) , .A1( u2_u11_u5_n152 ) , .ZN( u2_u11_u5_n165 ) );
  NAND2_X1 u2_u11_u5_U70 (.A2( u2_u11_u5_n103 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n151 ) );
  NAND2_X1 u2_u11_u5_U71 (.A2( u2_u11_u5_n107 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n120 ) );
  NAND2_X1 u2_u11_u5_U72 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n157 ) );
  AND2_X1 u2_u11_u5_U73 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n104 ) , .ZN( u2_u11_u5_n131 ) );
  INV_X1 u2_u11_u5_U74 (.A( u2_u11_u5_n102 ) , .ZN( u2_u11_u5_n195 ) );
  OAI221_X1 u2_u11_u5_U75 (.A( u2_u11_u5_n101 ) , .ZN( u2_u11_u5_n102 ) , .C2( u2_u11_u5_n115 ) , .C1( u2_u11_u5_n126 ) , .B1( u2_u11_u5_n134 ) , .B2( u2_u11_u5_n160 ) );
  OAI21_X1 u2_u11_u5_U76 (.ZN( u2_u11_u5_n101 ) , .B1( u2_u11_u5_n137 ) , .A( u2_u11_u5_n146 ) , .B2( u2_u11_u5_n147 ) );
  NOR2_X1 u2_u11_u5_U77 (.A2( u2_u11_X_34 ) , .A1( u2_u11_X_35 ) , .ZN( u2_u11_u5_n145 ) );
  NOR2_X1 u2_u11_u5_U78 (.A2( u2_u11_X_34 ) , .ZN( u2_u11_u5_n146 ) , .A1( u2_u11_u5_n171 ) );
  NOR2_X1 u2_u11_u5_U79 (.A2( u2_u11_X_31 ) , .A1( u2_u11_X_32 ) , .ZN( u2_u11_u5_n103 ) );
  NOR3_X1 u2_u11_u5_U8 (.A2( u2_u11_u5_n147 ) , .A1( u2_u11_u5_n148 ) , .ZN( u2_u11_u5_n149 ) , .A3( u2_u11_u5_n194 ) );
  NOR2_X1 u2_u11_u5_U80 (.A2( u2_u11_X_36 ) , .ZN( u2_u11_u5_n105 ) , .A1( u2_u11_u5_n180 ) );
  NOR2_X1 u2_u11_u5_U81 (.A2( u2_u11_X_33 ) , .ZN( u2_u11_u5_n108 ) , .A1( u2_u11_u5_n170 ) );
  NOR2_X1 u2_u11_u5_U82 (.A2( u2_u11_X_33 ) , .A1( u2_u11_X_36 ) , .ZN( u2_u11_u5_n107 ) );
  NOR2_X1 u2_u11_u5_U83 (.A2( u2_u11_X_31 ) , .ZN( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n181 ) );
  NAND2_X1 u2_u11_u5_U84 (.A2( u2_u11_X_34 ) , .A1( u2_u11_X_35 ) , .ZN( u2_u11_u5_n153 ) );
  NAND2_X1 u2_u11_u5_U85 (.A1( u2_u11_X_34 ) , .ZN( u2_u11_u5_n126 ) , .A2( u2_u11_u5_n171 ) );
  AND2_X1 u2_u11_u5_U86 (.A1( u2_u11_X_31 ) , .A2( u2_u11_X_32 ) , .ZN( u2_u11_u5_n106 ) );
  AND2_X1 u2_u11_u5_U87 (.A1( u2_u11_X_31 ) , .ZN( u2_u11_u5_n109 ) , .A2( u2_u11_u5_n181 ) );
  INV_X1 u2_u11_u5_U88 (.A( u2_u11_X_33 ) , .ZN( u2_u11_u5_n180 ) );
  INV_X1 u2_u11_u5_U89 (.A( u2_u11_X_35 ) , .ZN( u2_u11_u5_n171 ) );
  NOR2_X1 u2_u11_u5_U9 (.ZN( u2_u11_u5_n135 ) , .A1( u2_u11_u5_n173 ) , .A2( u2_u11_u5_n176 ) );
  INV_X1 u2_u11_u5_U90 (.A( u2_u11_X_36 ) , .ZN( u2_u11_u5_n170 ) );
  INV_X1 u2_u11_u5_U91 (.A( u2_u11_X_32 ) , .ZN( u2_u11_u5_n181 ) );
  NAND4_X1 u2_u11_u5_U92 (.ZN( u2_out11_29 ) , .A4( u2_u11_u5_n129 ) , .A3( u2_u11_u5_n130 ) , .A2( u2_u11_u5_n168 ) , .A1( u2_u11_u5_n196 ) );
  AOI221_X1 u2_u11_u5_U93 (.A( u2_u11_u5_n128 ) , .ZN( u2_u11_u5_n129 ) , .C2( u2_u11_u5_n132 ) , .B2( u2_u11_u5_n159 ) , .B1( u2_u11_u5_n176 ) , .C1( u2_u11_u5_n184 ) );
  AOI222_X1 u2_u11_u5_U94 (.ZN( u2_u11_u5_n130 ) , .A2( u2_u11_u5_n146 ) , .B1( u2_u11_u5_n147 ) , .C2( u2_u11_u5_n175 ) , .B2( u2_u11_u5_n179 ) , .A1( u2_u11_u5_n188 ) , .C1( u2_u11_u5_n194 ) );
  NAND4_X1 u2_u11_u5_U95 (.ZN( u2_out11_19 ) , .A4( u2_u11_u5_n166 ) , .A3( u2_u11_u5_n167 ) , .A2( u2_u11_u5_n168 ) , .A1( u2_u11_u5_n169 ) );
  AOI22_X1 u2_u11_u5_U96 (.B2( u2_u11_u5_n145 ) , .A2( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n167 ) , .B1( u2_u11_u5_n182 ) , .A1( u2_u11_u5_n189 ) );
  NOR4_X1 u2_u11_u5_U97 (.A4( u2_u11_u5_n162 ) , .A3( u2_u11_u5_n163 ) , .A2( u2_u11_u5_n164 ) , .A1( u2_u11_u5_n165 ) , .ZN( u2_u11_u5_n166 ) );
  NAND4_X1 u2_u11_u5_U98 (.ZN( u2_out11_11 ) , .A4( u2_u11_u5_n143 ) , .A3( u2_u11_u5_n144 ) , .A2( u2_u11_u5_n169 ) , .A1( u2_u11_u5_n196 ) );
  AOI22_X1 u2_u11_u5_U99 (.A2( u2_u11_u5_n132 ) , .ZN( u2_u11_u5_n144 ) , .B2( u2_u11_u5_n145 ) , .B1( u2_u11_u5_n184 ) , .A1( u2_u11_u5_n194 ) );
  OAI21_X1 u2_u11_u6_U10 (.A( u2_u11_u6_n159 ) , .B1( u2_u11_u6_n169 ) , .B2( u2_u11_u6_n173 ) , .ZN( u2_u11_u6_n90 ) );
  INV_X1 u2_u11_u6_U11 (.ZN( u2_u11_u6_n172 ) , .A( u2_u11_u6_n88 ) );
  AOI22_X1 u2_u11_u6_U12 (.A2( u2_u11_u6_n151 ) , .B2( u2_u11_u6_n161 ) , .A1( u2_u11_u6_n167 ) , .B1( u2_u11_u6_n170 ) , .ZN( u2_u11_u6_n89 ) );
  AOI21_X1 u2_u11_u6_U13 (.ZN( u2_u11_u6_n106 ) , .A( u2_u11_u6_n142 ) , .B2( u2_u11_u6_n159 ) , .B1( u2_u11_u6_n164 ) );
  INV_X1 u2_u11_u6_U14 (.A( u2_u11_u6_n155 ) , .ZN( u2_u11_u6_n161 ) );
  INV_X1 u2_u11_u6_U15 (.A( u2_u11_u6_n128 ) , .ZN( u2_u11_u6_n164 ) );
  NAND2_X1 u2_u11_u6_U16 (.ZN( u2_u11_u6_n110 ) , .A1( u2_u11_u6_n122 ) , .A2( u2_u11_u6_n129 ) );
  NAND2_X1 u2_u11_u6_U17 (.ZN( u2_u11_u6_n124 ) , .A2( u2_u11_u6_n146 ) , .A1( u2_u11_u6_n148 ) );
  INV_X1 u2_u11_u6_U18 (.A( u2_u11_u6_n132 ) , .ZN( u2_u11_u6_n171 ) );
  AND2_X1 u2_u11_u6_U19 (.A1( u2_u11_u6_n100 ) , .ZN( u2_u11_u6_n130 ) , .A2( u2_u11_u6_n147 ) );
  INV_X1 u2_u11_u6_U20 (.A( u2_u11_u6_n127 ) , .ZN( u2_u11_u6_n173 ) );
  INV_X1 u2_u11_u6_U21 (.A( u2_u11_u6_n121 ) , .ZN( u2_u11_u6_n167 ) );
  INV_X1 u2_u11_u6_U22 (.A( u2_u11_u6_n100 ) , .ZN( u2_u11_u6_n169 ) );
  INV_X1 u2_u11_u6_U23 (.A( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n170 ) );
  INV_X1 u2_u11_u6_U24 (.A( u2_u11_u6_n113 ) , .ZN( u2_u11_u6_n168 ) );
  AND2_X1 u2_u11_u6_U25 (.A1( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n119 ) , .ZN( u2_u11_u6_n133 ) );
  AND2_X1 u2_u11_u6_U26 (.A2( u2_u11_u6_n121 ) , .A1( u2_u11_u6_n122 ) , .ZN( u2_u11_u6_n131 ) );
  AND3_X1 u2_u11_u6_U27 (.ZN( u2_u11_u6_n120 ) , .A2( u2_u11_u6_n127 ) , .A1( u2_u11_u6_n132 ) , .A3( u2_u11_u6_n145 ) );
  INV_X1 u2_u11_u6_U28 (.A( u2_u11_u6_n146 ) , .ZN( u2_u11_u6_n163 ) );
  AOI222_X1 u2_u11_u6_U29 (.ZN( u2_u11_u6_n114 ) , .A1( u2_u11_u6_n118 ) , .A2( u2_u11_u6_n126 ) , .B2( u2_u11_u6_n151 ) , .C2( u2_u11_u6_n159 ) , .C1( u2_u11_u6_n168 ) , .B1( u2_u11_u6_n169 ) );
  INV_X1 u2_u11_u6_U3 (.A( u2_u11_u6_n110 ) , .ZN( u2_u11_u6_n166 ) );
  NOR2_X1 u2_u11_u6_U30 (.A1( u2_u11_u6_n162 ) , .A2( u2_u11_u6_n165 ) , .ZN( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U31 (.A1( u2_u11_u6_n144 ) , .ZN( u2_u11_u6_n151 ) , .A2( u2_u11_u6_n158 ) );
  NAND2_X1 u2_u11_u6_U32 (.ZN( u2_u11_u6_n132 ) , .A1( u2_u11_u6_n91 ) , .A2( u2_u11_u6_n97 ) );
  AOI22_X1 u2_u11_u6_U33 (.B2( u2_u11_u6_n110 ) , .B1( u2_u11_u6_n111 ) , .A1( u2_u11_u6_n112 ) , .ZN( u2_u11_u6_n115 ) , .A2( u2_u11_u6_n161 ) );
  NAND4_X1 u2_u11_u6_U34 (.A3( u2_u11_u6_n109 ) , .ZN( u2_u11_u6_n112 ) , .A4( u2_u11_u6_n132 ) , .A2( u2_u11_u6_n147 ) , .A1( u2_u11_u6_n166 ) );
  NOR2_X1 u2_u11_u6_U35 (.ZN( u2_u11_u6_n109 ) , .A1( u2_u11_u6_n170 ) , .A2( u2_u11_u6_n173 ) );
  NOR2_X1 u2_u11_u6_U36 (.A2( u2_u11_u6_n126 ) , .ZN( u2_u11_u6_n155 ) , .A1( u2_u11_u6_n160 ) );
  NAND2_X1 u2_u11_u6_U37 (.ZN( u2_u11_u6_n146 ) , .A2( u2_u11_u6_n94 ) , .A1( u2_u11_u6_n99 ) );
  AOI21_X1 u2_u11_u6_U38 (.A( u2_u11_u6_n144 ) , .B2( u2_u11_u6_n145 ) , .B1( u2_u11_u6_n146 ) , .ZN( u2_u11_u6_n150 ) );
  AOI211_X1 u2_u11_u6_U39 (.B( u2_u11_u6_n134 ) , .A( u2_u11_u6_n135 ) , .C1( u2_u11_u6_n136 ) , .ZN( u2_u11_u6_n137 ) , .C2( u2_u11_u6_n151 ) );
  INV_X1 u2_u11_u6_U4 (.A( u2_u11_u6_n142 ) , .ZN( u2_u11_u6_n174 ) );
  NAND4_X1 u2_u11_u6_U40 (.A4( u2_u11_u6_n127 ) , .A3( u2_u11_u6_n128 ) , .A2( u2_u11_u6_n129 ) , .A1( u2_u11_u6_n130 ) , .ZN( u2_u11_u6_n136 ) );
  AOI21_X1 u2_u11_u6_U41 (.B2( u2_u11_u6_n132 ) , .B1( u2_u11_u6_n133 ) , .ZN( u2_u11_u6_n134 ) , .A( u2_u11_u6_n158 ) );
  AOI21_X1 u2_u11_u6_U42 (.B1( u2_u11_u6_n131 ) , .ZN( u2_u11_u6_n135 ) , .A( u2_u11_u6_n144 ) , .B2( u2_u11_u6_n146 ) );
  INV_X1 u2_u11_u6_U43 (.A( u2_u11_u6_n111 ) , .ZN( u2_u11_u6_n158 ) );
  NAND2_X1 u2_u11_u6_U44 (.ZN( u2_u11_u6_n127 ) , .A1( u2_u11_u6_n91 ) , .A2( u2_u11_u6_n92 ) );
  NAND2_X1 u2_u11_u6_U45 (.ZN( u2_u11_u6_n129 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n96 ) );
  INV_X1 u2_u11_u6_U46 (.A( u2_u11_u6_n144 ) , .ZN( u2_u11_u6_n159 ) );
  NAND2_X1 u2_u11_u6_U47 (.ZN( u2_u11_u6_n145 ) , .A2( u2_u11_u6_n97 ) , .A1( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U48 (.ZN( u2_u11_u6_n148 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n94 ) );
  NAND2_X1 u2_u11_u6_U49 (.ZN( u2_u11_u6_n108 ) , .A2( u2_u11_u6_n139 ) , .A1( u2_u11_u6_n144 ) );
  NAND2_X1 u2_u11_u6_U5 (.A2( u2_u11_u6_n143 ) , .ZN( u2_u11_u6_n152 ) , .A1( u2_u11_u6_n166 ) );
  NAND2_X1 u2_u11_u6_U50 (.ZN( u2_u11_u6_n121 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n97 ) );
  NAND2_X1 u2_u11_u6_U51 (.ZN( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n95 ) );
  AND2_X1 u2_u11_u6_U52 (.ZN( u2_u11_u6_n118 ) , .A2( u2_u11_u6_n91 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U53 (.ZN( u2_u11_u6_n147 ) , .A2( u2_u11_u6_n98 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U54 (.ZN( u2_u11_u6_n128 ) , .A1( u2_u11_u6_n94 ) , .A2( u2_u11_u6_n96 ) );
  NAND2_X1 u2_u11_u6_U55 (.ZN( u2_u11_u6_n119 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U56 (.ZN( u2_u11_u6_n123 ) , .A2( u2_u11_u6_n91 ) , .A1( u2_u11_u6_n96 ) );
  NAND2_X1 u2_u11_u6_U57 (.ZN( u2_u11_u6_n100 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U58 (.ZN( u2_u11_u6_n122 ) , .A1( u2_u11_u6_n94 ) , .A2( u2_u11_u6_n97 ) );
  INV_X1 u2_u11_u6_U59 (.A( u2_u11_u6_n139 ) , .ZN( u2_u11_u6_n160 ) );
  AOI22_X1 u2_u11_u6_U6 (.B2( u2_u11_u6_n101 ) , .A1( u2_u11_u6_n102 ) , .ZN( u2_u11_u6_n103 ) , .B1( u2_u11_u6_n160 ) , .A2( u2_u11_u6_n161 ) );
  NAND2_X1 u2_u11_u6_U60 (.ZN( u2_u11_u6_n113 ) , .A1( u2_u11_u6_n96 ) , .A2( u2_u11_u6_n98 ) );
  NOR2_X1 u2_u11_u6_U61 (.A2( u2_u11_X_40 ) , .A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n126 ) );
  NOR2_X1 u2_u11_u6_U62 (.A2( u2_u11_X_39 ) , .A1( u2_u11_X_42 ) , .ZN( u2_u11_u6_n92 ) );
  NOR2_X1 u2_u11_u6_U63 (.A2( u2_u11_X_39 ) , .A1( u2_u11_u6_n156 ) , .ZN( u2_u11_u6_n97 ) );
  NOR2_X1 u2_u11_u6_U64 (.A2( u2_u11_X_38 ) , .A1( u2_u11_u6_n165 ) , .ZN( u2_u11_u6_n95 ) );
  NOR2_X1 u2_u11_u6_U65 (.A2( u2_u11_X_41 ) , .ZN( u2_u11_u6_n111 ) , .A1( u2_u11_u6_n157 ) );
  NOR2_X1 u2_u11_u6_U66 (.A2( u2_u11_X_37 ) , .A1( u2_u11_u6_n162 ) , .ZN( u2_u11_u6_n94 ) );
  NOR2_X1 u2_u11_u6_U67 (.A2( u2_u11_X_37 ) , .A1( u2_u11_X_38 ) , .ZN( u2_u11_u6_n91 ) );
  NAND2_X1 u2_u11_u6_U68 (.A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n144 ) , .A2( u2_u11_u6_n157 ) );
  NAND2_X1 u2_u11_u6_U69 (.A2( u2_u11_X_40 ) , .A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n139 ) );
  NOR2_X1 u2_u11_u6_U7 (.A1( u2_u11_u6_n118 ) , .ZN( u2_u11_u6_n143 ) , .A2( u2_u11_u6_n168 ) );
  AND2_X1 u2_u11_u6_U70 (.A1( u2_u11_X_39 ) , .A2( u2_u11_u6_n156 ) , .ZN( u2_u11_u6_n96 ) );
  AND2_X1 u2_u11_u6_U71 (.A1( u2_u11_X_39 ) , .A2( u2_u11_X_42 ) , .ZN( u2_u11_u6_n99 ) );
  INV_X1 u2_u11_u6_U72 (.A( u2_u11_X_40 ) , .ZN( u2_u11_u6_n157 ) );
  INV_X1 u2_u11_u6_U73 (.A( u2_u11_X_37 ) , .ZN( u2_u11_u6_n165 ) );
  INV_X1 u2_u11_u6_U74 (.A( u2_u11_X_38 ) , .ZN( u2_u11_u6_n162 ) );
  INV_X1 u2_u11_u6_U75 (.A( u2_u11_X_42 ) , .ZN( u2_u11_u6_n156 ) );
  NAND4_X1 u2_u11_u6_U76 (.ZN( u2_out11_32 ) , .A4( u2_u11_u6_n103 ) , .A3( u2_u11_u6_n104 ) , .A2( u2_u11_u6_n105 ) , .A1( u2_u11_u6_n106 ) );
  AOI22_X1 u2_u11_u6_U77 (.ZN( u2_u11_u6_n105 ) , .A2( u2_u11_u6_n108 ) , .A1( u2_u11_u6_n118 ) , .B2( u2_u11_u6_n126 ) , .B1( u2_u11_u6_n171 ) );
  AOI22_X1 u2_u11_u6_U78 (.ZN( u2_u11_u6_n104 ) , .A1( u2_u11_u6_n111 ) , .B1( u2_u11_u6_n124 ) , .B2( u2_u11_u6_n151 ) , .A2( u2_u11_u6_n93 ) );
  NAND4_X1 u2_u11_u6_U79 (.ZN( u2_out11_12 ) , .A4( u2_u11_u6_n114 ) , .A3( u2_u11_u6_n115 ) , .A2( u2_u11_u6_n116 ) , .A1( u2_u11_u6_n117 ) );
  AOI21_X1 u2_u11_u6_U8 (.B1( u2_u11_u6_n107 ) , .B2( u2_u11_u6_n132 ) , .A( u2_u11_u6_n158 ) , .ZN( u2_u11_u6_n88 ) );
  OAI22_X1 u2_u11_u6_U80 (.B2( u2_u11_u6_n111 ) , .ZN( u2_u11_u6_n116 ) , .B1( u2_u11_u6_n126 ) , .A2( u2_u11_u6_n164 ) , .A1( u2_u11_u6_n167 ) );
  OAI21_X1 u2_u11_u6_U81 (.A( u2_u11_u6_n108 ) , .ZN( u2_u11_u6_n117 ) , .B2( u2_u11_u6_n141 ) , .B1( u2_u11_u6_n163 ) );
  OAI211_X1 u2_u11_u6_U82 (.ZN( u2_out11_7 ) , .B( u2_u11_u6_n153 ) , .C2( u2_u11_u6_n154 ) , .C1( u2_u11_u6_n155 ) , .A( u2_u11_u6_n174 ) );
  NOR3_X1 u2_u11_u6_U83 (.A1( u2_u11_u6_n141 ) , .ZN( u2_u11_u6_n154 ) , .A3( u2_u11_u6_n164 ) , .A2( u2_u11_u6_n171 ) );
  AOI211_X1 u2_u11_u6_U84 (.B( u2_u11_u6_n149 ) , .A( u2_u11_u6_n150 ) , .C2( u2_u11_u6_n151 ) , .C1( u2_u11_u6_n152 ) , .ZN( u2_u11_u6_n153 ) );
  OAI211_X1 u2_u11_u6_U85 (.ZN( u2_out11_22 ) , .B( u2_u11_u6_n137 ) , .A( u2_u11_u6_n138 ) , .C2( u2_u11_u6_n139 ) , .C1( u2_u11_u6_n140 ) );
  AOI22_X1 u2_u11_u6_U86 (.B1( u2_u11_u6_n124 ) , .A2( u2_u11_u6_n125 ) , .A1( u2_u11_u6_n126 ) , .ZN( u2_u11_u6_n138 ) , .B2( u2_u11_u6_n161 ) );
  AND4_X1 u2_u11_u6_U87 (.A3( u2_u11_u6_n119 ) , .A1( u2_u11_u6_n120 ) , .A4( u2_u11_u6_n129 ) , .ZN( u2_u11_u6_n140 ) , .A2( u2_u11_u6_n143 ) );
  NAND3_X1 u2_u11_u6_U88 (.A2( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n125 ) , .A1( u2_u11_u6_n130 ) , .A3( u2_u11_u6_n131 ) );
  NAND3_X1 u2_u11_u6_U89 (.A3( u2_u11_u6_n133 ) , .ZN( u2_u11_u6_n141 ) , .A1( u2_u11_u6_n145 ) , .A2( u2_u11_u6_n148 ) );
  AOI21_X1 u2_u11_u6_U9 (.B2( u2_u11_u6_n147 ) , .B1( u2_u11_u6_n148 ) , .ZN( u2_u11_u6_n149 ) , .A( u2_u11_u6_n158 ) );
  NAND3_X1 u2_u11_u6_U90 (.ZN( u2_u11_u6_n101 ) , .A3( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n121 ) , .A1( u2_u11_u6_n127 ) );
  NAND3_X1 u2_u11_u6_U91 (.ZN( u2_u11_u6_n102 ) , .A3( u2_u11_u6_n130 ) , .A2( u2_u11_u6_n145 ) , .A1( u2_u11_u6_n166 ) );
  NAND3_X1 u2_u11_u6_U92 (.A3( u2_u11_u6_n113 ) , .A1( u2_u11_u6_n119 ) , .A2( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n93 ) );
  NAND3_X1 u2_u11_u6_U93 (.ZN( u2_u11_u6_n142 ) , .A2( u2_u11_u6_n172 ) , .A3( u2_u11_u6_n89 ) , .A1( u2_u11_u6_n90 ) );
  AND3_X1 u2_u11_u7_U10 (.A3( u2_u11_u7_n110 ) , .A2( u2_u11_u7_n127 ) , .A1( u2_u11_u7_n132 ) , .ZN( u2_u11_u7_n92 ) );
  OAI21_X1 u2_u11_u7_U11 (.A( u2_u11_u7_n161 ) , .B1( u2_u11_u7_n168 ) , .B2( u2_u11_u7_n173 ) , .ZN( u2_u11_u7_n91 ) );
  AOI211_X1 u2_u11_u7_U12 (.A( u2_u11_u7_n117 ) , .ZN( u2_u11_u7_n118 ) , .C2( u2_u11_u7_n126 ) , .C1( u2_u11_u7_n177 ) , .B( u2_u11_u7_n180 ) );
  OAI22_X1 u2_u11_u7_U13 (.B1( u2_u11_u7_n115 ) , .ZN( u2_u11_u7_n117 ) , .A2( u2_u11_u7_n133 ) , .A1( u2_u11_u7_n137 ) , .B2( u2_u11_u7_n162 ) );
  INV_X1 u2_u11_u7_U14 (.A( u2_u11_u7_n116 ) , .ZN( u2_u11_u7_n180 ) );
  NOR3_X1 u2_u11_u7_U15 (.ZN( u2_u11_u7_n115 ) , .A3( u2_u11_u7_n145 ) , .A2( u2_u11_u7_n168 ) , .A1( u2_u11_u7_n169 ) );
  OAI211_X1 u2_u11_u7_U16 (.B( u2_u11_u7_n122 ) , .A( u2_u11_u7_n123 ) , .C2( u2_u11_u7_n124 ) , .ZN( u2_u11_u7_n154 ) , .C1( u2_u11_u7_n162 ) );
  AOI222_X1 u2_u11_u7_U17 (.ZN( u2_u11_u7_n122 ) , .C2( u2_u11_u7_n126 ) , .C1( u2_u11_u7_n145 ) , .B1( u2_u11_u7_n161 ) , .A2( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n170 ) , .A1( u2_u11_u7_n176 ) );
  INV_X1 u2_u11_u7_U18 (.A( u2_u11_u7_n133 ) , .ZN( u2_u11_u7_n176 ) );
  NOR3_X1 u2_u11_u7_U19 (.A2( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n135 ) , .ZN( u2_u11_u7_n136 ) , .A3( u2_u11_u7_n171 ) );
  NOR2_X1 u2_u11_u7_U20 (.A1( u2_u11_u7_n130 ) , .A2( u2_u11_u7_n134 ) , .ZN( u2_u11_u7_n153 ) );
  INV_X1 u2_u11_u7_U21 (.A( u2_u11_u7_n101 ) , .ZN( u2_u11_u7_n165 ) );
  NOR2_X1 u2_u11_u7_U22 (.ZN( u2_u11_u7_n111 ) , .A2( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n169 ) );
  AOI21_X1 u2_u11_u7_U23 (.ZN( u2_u11_u7_n104 ) , .B2( u2_u11_u7_n112 ) , .B1( u2_u11_u7_n127 ) , .A( u2_u11_u7_n164 ) );
  AOI21_X1 u2_u11_u7_U24 (.ZN( u2_u11_u7_n106 ) , .B1( u2_u11_u7_n133 ) , .B2( u2_u11_u7_n146 ) , .A( u2_u11_u7_n162 ) );
  AOI21_X1 u2_u11_u7_U25 (.A( u2_u11_u7_n101 ) , .ZN( u2_u11_u7_n107 ) , .B2( u2_u11_u7_n128 ) , .B1( u2_u11_u7_n175 ) );
  INV_X1 u2_u11_u7_U26 (.A( u2_u11_u7_n138 ) , .ZN( u2_u11_u7_n171 ) );
  INV_X1 u2_u11_u7_U27 (.A( u2_u11_u7_n131 ) , .ZN( u2_u11_u7_n177 ) );
  INV_X1 u2_u11_u7_U28 (.A( u2_u11_u7_n110 ) , .ZN( u2_u11_u7_n174 ) );
  NAND2_X1 u2_u11_u7_U29 (.A1( u2_u11_u7_n129 ) , .A2( u2_u11_u7_n132 ) , .ZN( u2_u11_u7_n149 ) );
  OAI21_X1 u2_u11_u7_U3 (.ZN( u2_u11_u7_n159 ) , .A( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n171 ) , .B1( u2_u11_u7_n174 ) );
  NAND2_X1 u2_u11_u7_U30 (.A1( u2_u11_u7_n113 ) , .A2( u2_u11_u7_n124 ) , .ZN( u2_u11_u7_n130 ) );
  INV_X1 u2_u11_u7_U31 (.A( u2_u11_u7_n112 ) , .ZN( u2_u11_u7_n173 ) );
  INV_X1 u2_u11_u7_U32 (.A( u2_u11_u7_n128 ) , .ZN( u2_u11_u7_n168 ) );
  INV_X1 u2_u11_u7_U33 (.A( u2_u11_u7_n148 ) , .ZN( u2_u11_u7_n169 ) );
  INV_X1 u2_u11_u7_U34 (.A( u2_u11_u7_n127 ) , .ZN( u2_u11_u7_n179 ) );
  NOR2_X1 u2_u11_u7_U35 (.ZN( u2_u11_u7_n101 ) , .A2( u2_u11_u7_n150 ) , .A1( u2_u11_u7_n156 ) );
  AOI211_X1 u2_u11_u7_U36 (.B( u2_u11_u7_n154 ) , .A( u2_u11_u7_n155 ) , .C1( u2_u11_u7_n156 ) , .ZN( u2_u11_u7_n157 ) , .C2( u2_u11_u7_n172 ) );
  INV_X1 u2_u11_u7_U37 (.A( u2_u11_u7_n153 ) , .ZN( u2_u11_u7_n172 ) );
  AOI211_X1 u2_u11_u7_U38 (.B( u2_u11_u7_n139 ) , .A( u2_u11_u7_n140 ) , .C2( u2_u11_u7_n141 ) , .ZN( u2_u11_u7_n142 ) , .C1( u2_u11_u7_n156 ) );
  AOI21_X1 u2_u11_u7_U39 (.A( u2_u11_u7_n137 ) , .B1( u2_u11_u7_n138 ) , .ZN( u2_u11_u7_n139 ) , .B2( u2_u11_u7_n146 ) );
  INV_X1 u2_u11_u7_U4 (.A( u2_u11_u7_n111 ) , .ZN( u2_u11_u7_n170 ) );
  NAND4_X1 u2_u11_u7_U40 (.A3( u2_u11_u7_n127 ) , .A2( u2_u11_u7_n128 ) , .A1( u2_u11_u7_n129 ) , .ZN( u2_u11_u7_n141 ) , .A4( u2_u11_u7_n147 ) );
  OAI22_X1 u2_u11_u7_U41 (.B1( u2_u11_u7_n136 ) , .ZN( u2_u11_u7_n140 ) , .A1( u2_u11_u7_n153 ) , .B2( u2_u11_u7_n162 ) , .A2( u2_u11_u7_n164 ) );
  AOI21_X1 u2_u11_u7_U42 (.ZN( u2_u11_u7_n123 ) , .B1( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n177 ) , .A( u2_u11_u7_n97 ) );
  AOI21_X1 u2_u11_u7_U43 (.B2( u2_u11_u7_n113 ) , .B1( u2_u11_u7_n124 ) , .A( u2_u11_u7_n125 ) , .ZN( u2_u11_u7_n97 ) );
  INV_X1 u2_u11_u7_U44 (.A( u2_u11_u7_n125 ) , .ZN( u2_u11_u7_n161 ) );
  INV_X1 u2_u11_u7_U45 (.A( u2_u11_u7_n152 ) , .ZN( u2_u11_u7_n162 ) );
  AOI22_X1 u2_u11_u7_U46 (.A2( u2_u11_u7_n114 ) , .ZN( u2_u11_u7_n119 ) , .B1( u2_u11_u7_n130 ) , .A1( u2_u11_u7_n156 ) , .B2( u2_u11_u7_n165 ) );
  NAND2_X1 u2_u11_u7_U47 (.A2( u2_u11_u7_n112 ) , .ZN( u2_u11_u7_n114 ) , .A1( u2_u11_u7_n175 ) );
  AND2_X1 u2_u11_u7_U48 (.ZN( u2_u11_u7_n145 ) , .A2( u2_u11_u7_n98 ) , .A1( u2_u11_u7_n99 ) );
  NOR2_X1 u2_u11_u7_U49 (.ZN( u2_u11_u7_n137 ) , .A1( u2_u11_u7_n150 ) , .A2( u2_u11_u7_n161 ) );
  INV_X1 u2_u11_u7_U5 (.A( u2_u11_u7_n149 ) , .ZN( u2_u11_u7_n175 ) );
  AOI21_X1 u2_u11_u7_U50 (.ZN( u2_u11_u7_n105 ) , .B2( u2_u11_u7_n110 ) , .A( u2_u11_u7_n125 ) , .B1( u2_u11_u7_n147 ) );
  NAND2_X1 u2_u11_u7_U51 (.ZN( u2_u11_u7_n146 ) , .A1( u2_u11_u7_n95 ) , .A2( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U52 (.A2( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n147 ) , .A1( u2_u11_u7_n93 ) );
  NAND2_X1 u2_u11_u7_U53 (.A1( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n127 ) , .A2( u2_u11_u7_n99 ) );
  OR2_X1 u2_u11_u7_U54 (.ZN( u2_u11_u7_n126 ) , .A2( u2_u11_u7_n152 ) , .A1( u2_u11_u7_n156 ) );
  NAND2_X1 u2_u11_u7_U55 (.A2( u2_u11_u7_n102 ) , .A1( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n133 ) );
  NAND2_X1 u2_u11_u7_U56 (.ZN( u2_u11_u7_n112 ) , .A2( u2_u11_u7_n96 ) , .A1( u2_u11_u7_n99 ) );
  NAND2_X1 u2_u11_u7_U57 (.A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n128 ) , .A1( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U58 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n113 ) , .A2( u2_u11_u7_n93 ) );
  NAND2_X1 u2_u11_u7_U59 (.A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n124 ) , .A1( u2_u11_u7_n96 ) );
  INV_X1 u2_u11_u7_U6 (.A( u2_u11_u7_n154 ) , .ZN( u2_u11_u7_n178 ) );
  NAND2_X1 u2_u11_u7_U60 (.ZN( u2_u11_u7_n110 ) , .A1( u2_u11_u7_n95 ) , .A2( u2_u11_u7_n96 ) );
  INV_X1 u2_u11_u7_U61 (.A( u2_u11_u7_n150 ) , .ZN( u2_u11_u7_n164 ) );
  AND2_X1 u2_u11_u7_U62 (.ZN( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n93 ) , .A2( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U63 (.A1( u2_u11_u7_n100 ) , .A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n129 ) );
  NAND2_X1 u2_u11_u7_U64 (.A2( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n131 ) , .A1( u2_u11_u7_n95 ) );
  NAND2_X1 u2_u11_u7_U65 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n138 ) , .A2( u2_u11_u7_n99 ) );
  NAND2_X1 u2_u11_u7_U66 (.ZN( u2_u11_u7_n132 ) , .A1( u2_u11_u7_n93 ) , .A2( u2_u11_u7_n96 ) );
  NAND2_X1 u2_u11_u7_U67 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n148 ) , .A2( u2_u11_u7_n95 ) );
  NOR2_X1 u2_u11_u7_U68 (.A2( u2_u11_X_47 ) , .ZN( u2_u11_u7_n150 ) , .A1( u2_u11_u7_n163 ) );
  NOR2_X1 u2_u11_u7_U69 (.A2( u2_u11_X_43 ) , .A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n103 ) );
  AOI211_X1 u2_u11_u7_U7 (.ZN( u2_u11_u7_n116 ) , .A( u2_u11_u7_n155 ) , .C1( u2_u11_u7_n161 ) , .C2( u2_u11_u7_n171 ) , .B( u2_u11_u7_n94 ) );
  NOR2_X1 u2_u11_u7_U70 (.A2( u2_u11_X_48 ) , .A1( u2_u11_u7_n166 ) , .ZN( u2_u11_u7_n95 ) );
  NOR2_X1 u2_u11_u7_U71 (.A2( u2_u11_X_45 ) , .A1( u2_u11_X_48 ) , .ZN( u2_u11_u7_n99 ) );
  NOR2_X1 u2_u11_u7_U72 (.A2( u2_u11_X_44 ) , .A1( u2_u11_u7_n167 ) , .ZN( u2_u11_u7_n98 ) );
  NOR2_X1 u2_u11_u7_U73 (.A2( u2_u11_X_46 ) , .A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n152 ) );
  AND2_X1 u2_u11_u7_U74 (.A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n156 ) , .A2( u2_u11_u7_n163 ) );
  NAND2_X1 u2_u11_u7_U75 (.A2( u2_u11_X_46 ) , .A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n125 ) );
  AND2_X1 u2_u11_u7_U76 (.A2( u2_u11_X_45 ) , .A1( u2_u11_X_48 ) , .ZN( u2_u11_u7_n102 ) );
  AND2_X1 u2_u11_u7_U77 (.A2( u2_u11_X_43 ) , .A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n96 ) );
  AND2_X1 u2_u11_u7_U78 (.A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n100 ) , .A2( u2_u11_u7_n167 ) );
  AND2_X1 u2_u11_u7_U79 (.A1( u2_u11_X_48 ) , .A2( u2_u11_u7_n166 ) , .ZN( u2_u11_u7_n93 ) );
  OAI222_X1 u2_u11_u7_U8 (.C2( u2_u11_u7_n101 ) , .B2( u2_u11_u7_n111 ) , .A1( u2_u11_u7_n113 ) , .C1( u2_u11_u7_n146 ) , .A2( u2_u11_u7_n162 ) , .B1( u2_u11_u7_n164 ) , .ZN( u2_u11_u7_n94 ) );
  INV_X1 u2_u11_u7_U80 (.A( u2_u11_X_46 ) , .ZN( u2_u11_u7_n163 ) );
  INV_X1 u2_u11_u7_U81 (.A( u2_u11_X_43 ) , .ZN( u2_u11_u7_n167 ) );
  INV_X1 u2_u11_u7_U82 (.A( u2_u11_X_45 ) , .ZN( u2_u11_u7_n166 ) );
  NAND4_X1 u2_u11_u7_U83 (.ZN( u2_out11_27 ) , .A4( u2_u11_u7_n118 ) , .A3( u2_u11_u7_n119 ) , .A2( u2_u11_u7_n120 ) , .A1( u2_u11_u7_n121 ) );
  OAI21_X1 u2_u11_u7_U84 (.ZN( u2_u11_u7_n121 ) , .B2( u2_u11_u7_n145 ) , .A( u2_u11_u7_n150 ) , .B1( u2_u11_u7_n174 ) );
  OAI21_X1 u2_u11_u7_U85 (.ZN( u2_u11_u7_n120 ) , .A( u2_u11_u7_n161 ) , .B2( u2_u11_u7_n170 ) , .B1( u2_u11_u7_n179 ) );
  NAND4_X1 u2_u11_u7_U86 (.ZN( u2_out11_21 ) , .A4( u2_u11_u7_n157 ) , .A3( u2_u11_u7_n158 ) , .A2( u2_u11_u7_n159 ) , .A1( u2_u11_u7_n160 ) );
  OAI21_X1 u2_u11_u7_U87 (.B1( u2_u11_u7_n145 ) , .ZN( u2_u11_u7_n160 ) , .A( u2_u11_u7_n161 ) , .B2( u2_u11_u7_n177 ) );
  AOI22_X1 u2_u11_u7_U88 (.B2( u2_u11_u7_n149 ) , .B1( u2_u11_u7_n150 ) , .A2( u2_u11_u7_n151 ) , .A1( u2_u11_u7_n152 ) , .ZN( u2_u11_u7_n158 ) );
  NAND4_X1 u2_u11_u7_U89 (.ZN( u2_out11_15 ) , .A4( u2_u11_u7_n142 ) , .A3( u2_u11_u7_n143 ) , .A2( u2_u11_u7_n144 ) , .A1( u2_u11_u7_n178 ) );
  OAI221_X1 u2_u11_u7_U9 (.C1( u2_u11_u7_n101 ) , .C2( u2_u11_u7_n147 ) , .ZN( u2_u11_u7_n155 ) , .B2( u2_u11_u7_n162 ) , .A( u2_u11_u7_n91 ) , .B1( u2_u11_u7_n92 ) );
  OR2_X1 u2_u11_u7_U90 (.A2( u2_u11_u7_n125 ) , .A1( u2_u11_u7_n129 ) , .ZN( u2_u11_u7_n144 ) );
  AOI22_X1 u2_u11_u7_U91 (.A2( u2_u11_u7_n126 ) , .ZN( u2_u11_u7_n143 ) , .B2( u2_u11_u7_n165 ) , .B1( u2_u11_u7_n173 ) , .A1( u2_u11_u7_n174 ) );
  NAND4_X1 u2_u11_u7_U92 (.ZN( u2_out11_5 ) , .A4( u2_u11_u7_n108 ) , .A3( u2_u11_u7_n109 ) , .A1( u2_u11_u7_n116 ) , .A2( u2_u11_u7_n123 ) );
  AOI22_X1 u2_u11_u7_U93 (.ZN( u2_u11_u7_n109 ) , .A2( u2_u11_u7_n126 ) , .B2( u2_u11_u7_n145 ) , .B1( u2_u11_u7_n156 ) , .A1( u2_u11_u7_n171 ) );
  NOR4_X1 u2_u11_u7_U94 (.A4( u2_u11_u7_n104 ) , .A3( u2_u11_u7_n105 ) , .A2( u2_u11_u7_n106 ) , .A1( u2_u11_u7_n107 ) , .ZN( u2_u11_u7_n108 ) );
  NAND3_X1 u2_u11_u7_U95 (.A3( u2_u11_u7_n146 ) , .A2( u2_u11_u7_n147 ) , .A1( u2_u11_u7_n148 ) , .ZN( u2_u11_u7_n151 ) );
  NAND3_X1 u2_u11_u7_U96 (.A3( u2_u11_u7_n131 ) , .A2( u2_u11_u7_n132 ) , .A1( u2_u11_u7_n133 ) , .ZN( u2_u11_u7_n135 ) );
  XOR2_X1 u2_u14_U1 (.B( u2_K15_9 ) , .A( u2_R13_6 ) , .Z( u2_u14_X_9 ) );
  XOR2_X1 u2_u14_U16 (.B( u2_K15_3 ) , .A( u2_R13_2 ) , .Z( u2_u14_X_3 ) );
  XOR2_X1 u2_u14_U2 (.B( u2_K15_8 ) , .A( u2_R13_5 ) , .Z( u2_u14_X_8 ) );
  XOR2_X1 u2_u14_U27 (.B( u2_K15_2 ) , .A( u2_R13_1 ) , .Z( u2_u14_X_2 ) );
  XOR2_X1 u2_u14_U3 (.B( u2_K15_7 ) , .A( u2_R13_4 ) , .Z( u2_u14_X_7 ) );
  XOR2_X1 u2_u14_U33 (.B( u2_K15_24 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_24 ) );
  XOR2_X1 u2_u14_U34 (.B( u2_K15_23 ) , .A( u2_R13_16 ) , .Z( u2_u14_X_23 ) );
  XOR2_X1 u2_u14_U35 (.B( u2_K15_22 ) , .A( u2_R13_15 ) , .Z( u2_u14_X_22 ) );
  XOR2_X1 u2_u14_U36 (.B( u2_K15_21 ) , .A( u2_R13_14 ) , .Z( u2_u14_X_21 ) );
  XOR2_X1 u2_u14_U37 (.B( u2_K15_20 ) , .A( u2_R13_13 ) , .Z( u2_u14_X_20 ) );
  XOR2_X1 u2_u14_U38 (.B( u2_K15_1 ) , .A( u2_R13_32 ) , .Z( u2_u14_X_1 ) );
  XOR2_X1 u2_u14_U39 (.B( u2_K15_19 ) , .A( u2_R13_12 ) , .Z( u2_u14_X_19 ) );
  XOR2_X1 u2_u14_U4 (.B( u2_K15_6 ) , .A( u2_R13_5 ) , .Z( u2_u14_X_6 ) );
  XOR2_X1 u2_u14_U40 (.B( u2_K15_18 ) , .A( u2_R13_13 ) , .Z( u2_u14_X_18 ) );
  XOR2_X1 u2_u14_U41 (.B( u2_K15_17 ) , .A( u2_R13_12 ) , .Z( u2_u14_X_17 ) );
  XOR2_X1 u2_u14_U42 (.B( u2_K15_16 ) , .A( u2_R13_11 ) , .Z( u2_u14_X_16 ) );
  XOR2_X1 u2_u14_U43 (.B( u2_K15_15 ) , .A( u2_R13_10 ) , .Z( u2_u14_X_15 ) );
  XOR2_X1 u2_u14_U44 (.B( u2_K15_14 ) , .A( u2_R13_9 ) , .Z( u2_u14_X_14 ) );
  XOR2_X1 u2_u14_U45 (.B( u2_K15_13 ) , .A( u2_R13_8 ) , .Z( u2_u14_X_13 ) );
  XOR2_X1 u2_u14_U46 (.B( u2_K15_12 ) , .A( u2_R13_9 ) , .Z( u2_u14_X_12 ) );
  XOR2_X1 u2_u14_U47 (.B( u2_K15_11 ) , .A( u2_R13_8 ) , .Z( u2_u14_X_11 ) );
  XOR2_X1 u2_u14_U48 (.B( u2_K15_10 ) , .A( u2_R13_7 ) , .Z( u2_u14_X_10 ) );
  XOR2_X1 u2_u14_U5 (.B( u2_K15_5 ) , .A( u2_R13_4 ) , .Z( u2_u14_X_5 ) );
  XOR2_X1 u2_u14_U6 (.B( u2_K15_4 ) , .A( u2_R13_3 ) , .Z( u2_u14_X_4 ) );
  AND3_X1 u2_u14_u0_U10 (.A2( u2_u14_u0_n112 ) , .ZN( u2_u14_u0_n127 ) , .A3( u2_u14_u0_n130 ) , .A1( u2_u14_u0_n148 ) );
  NAND2_X1 u2_u14_u0_U11 (.ZN( u2_u14_u0_n113 ) , .A1( u2_u14_u0_n139 ) , .A2( u2_u14_u0_n149 ) );
  AND2_X1 u2_u14_u0_U12 (.ZN( u2_u14_u0_n107 ) , .A1( u2_u14_u0_n130 ) , .A2( u2_u14_u0_n140 ) );
  AND2_X1 u2_u14_u0_U13 (.A2( u2_u14_u0_n129 ) , .A1( u2_u14_u0_n130 ) , .ZN( u2_u14_u0_n151 ) );
  AND2_X1 u2_u14_u0_U14 (.A1( u2_u14_u0_n108 ) , .A2( u2_u14_u0_n125 ) , .ZN( u2_u14_u0_n145 ) );
  INV_X1 u2_u14_u0_U15 (.A( u2_u14_u0_n143 ) , .ZN( u2_u14_u0_n173 ) );
  NOR2_X1 u2_u14_u0_U16 (.A2( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n147 ) , .A1( u2_u14_u0_n160 ) );
  NOR2_X1 u2_u14_u0_U17 (.A1( u2_u14_u0_n163 ) , .A2( u2_u14_u0_n164 ) , .ZN( u2_u14_u0_n95 ) );
  AOI21_X1 u2_u14_u0_U18 (.B1( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n132 ) , .A( u2_u14_u0_n165 ) , .B2( u2_u14_u0_n93 ) );
  INV_X1 u2_u14_u0_U19 (.A( u2_u14_u0_n142 ) , .ZN( u2_u14_u0_n165 ) );
  OAI221_X1 u2_u14_u0_U20 (.C1( u2_u14_u0_n121 ) , .ZN( u2_u14_u0_n122 ) , .B2( u2_u14_u0_n127 ) , .A( u2_u14_u0_n143 ) , .B1( u2_u14_u0_n144 ) , .C2( u2_u14_u0_n147 ) );
  OAI22_X1 u2_u14_u0_U21 (.B1( u2_u14_u0_n125 ) , .ZN( u2_u14_u0_n126 ) , .A1( u2_u14_u0_n138 ) , .A2( u2_u14_u0_n146 ) , .B2( u2_u14_u0_n147 ) );
  OAI22_X1 u2_u14_u0_U22 (.B1( u2_u14_u0_n131 ) , .A1( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n147 ) , .A2( u2_u14_u0_n90 ) , .ZN( u2_u14_u0_n91 ) );
  AND3_X1 u2_u14_u0_U23 (.A3( u2_u14_u0_n121 ) , .A2( u2_u14_u0_n125 ) , .A1( u2_u14_u0_n148 ) , .ZN( u2_u14_u0_n90 ) );
  INV_X1 u2_u14_u0_U24 (.A( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n161 ) );
  NOR2_X1 u2_u14_u0_U25 (.A1( u2_u14_u0_n120 ) , .ZN( u2_u14_u0_n143 ) , .A2( u2_u14_u0_n167 ) );
  OAI221_X1 u2_u14_u0_U26 (.C1( u2_u14_u0_n112 ) , .ZN( u2_u14_u0_n120 ) , .B1( u2_u14_u0_n138 ) , .B2( u2_u14_u0_n141 ) , .C2( u2_u14_u0_n147 ) , .A( u2_u14_u0_n172 ) );
  AOI211_X1 u2_u14_u0_U27 (.B( u2_u14_u0_n115 ) , .A( u2_u14_u0_n116 ) , .C2( u2_u14_u0_n117 ) , .C1( u2_u14_u0_n118 ) , .ZN( u2_u14_u0_n119 ) );
  AOI22_X1 u2_u14_u0_U28 (.B2( u2_u14_u0_n109 ) , .A2( u2_u14_u0_n110 ) , .ZN( u2_u14_u0_n111 ) , .B1( u2_u14_u0_n118 ) , .A1( u2_u14_u0_n160 ) );
  INV_X1 u2_u14_u0_U29 (.A( u2_u14_u0_n118 ) , .ZN( u2_u14_u0_n158 ) );
  INV_X1 u2_u14_u0_U3 (.A( u2_u14_u0_n113 ) , .ZN( u2_u14_u0_n166 ) );
  AOI21_X1 u2_u14_u0_U30 (.ZN( u2_u14_u0_n104 ) , .B1( u2_u14_u0_n107 ) , .B2( u2_u14_u0_n141 ) , .A( u2_u14_u0_n144 ) );
  AOI21_X1 u2_u14_u0_U31 (.B1( u2_u14_u0_n127 ) , .B2( u2_u14_u0_n129 ) , .A( u2_u14_u0_n138 ) , .ZN( u2_u14_u0_n96 ) );
  AOI21_X1 u2_u14_u0_U32 (.ZN( u2_u14_u0_n116 ) , .B2( u2_u14_u0_n142 ) , .A( u2_u14_u0_n144 ) , .B1( u2_u14_u0_n166 ) );
  NAND2_X1 u2_u14_u0_U33 (.A1( u2_u14_u0_n100 ) , .A2( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n125 ) );
  NAND2_X1 u2_u14_u0_U34 (.A2( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n140 ) , .A1( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U35 (.A1( u2_u14_u0_n101 ) , .A2( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n150 ) );
  INV_X1 u2_u14_u0_U36 (.A( u2_u14_u0_n138 ) , .ZN( u2_u14_u0_n160 ) );
  NAND2_X1 u2_u14_u0_U37 (.ZN( u2_u14_u0_n142 ) , .A1( u2_u14_u0_n94 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U38 (.A1( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n128 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U39 (.A2( u2_u14_u0_n102 ) , .A1( u2_u14_u0_n103 ) , .ZN( u2_u14_u0_n149 ) );
  AOI21_X1 u2_u14_u0_U4 (.B1( u2_u14_u0_n114 ) , .ZN( u2_u14_u0_n115 ) , .B2( u2_u14_u0_n129 ) , .A( u2_u14_u0_n161 ) );
  NAND2_X1 u2_u14_u0_U40 (.A1( u2_u14_u0_n100 ) , .ZN( u2_u14_u0_n129 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U41 (.A2( u2_u14_u0_n100 ) , .A1( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n139 ) );
  NAND2_X1 u2_u14_u0_U42 (.A2( u2_u14_u0_n100 ) , .ZN( u2_u14_u0_n131 ) , .A1( u2_u14_u0_n92 ) );
  NAND2_X1 u2_u14_u0_U43 (.ZN( u2_u14_u0_n108 ) , .A1( u2_u14_u0_n92 ) , .A2( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U44 (.ZN( u2_u14_u0_n148 ) , .A1( u2_u14_u0_n93 ) , .A2( u2_u14_u0_n95 ) );
  NAND2_X1 u2_u14_u0_U45 (.A2( u2_u14_u0_n102 ) , .ZN( u2_u14_u0_n114 ) , .A1( u2_u14_u0_n92 ) );
  NAND2_X1 u2_u14_u0_U46 (.A1( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n130 ) , .A2( u2_u14_u0_n94 ) );
  NAND2_X1 u2_u14_u0_U47 (.A2( u2_u14_u0_n101 ) , .ZN( u2_u14_u0_n121 ) , .A1( u2_u14_u0_n93 ) );
  INV_X1 u2_u14_u0_U48 (.ZN( u2_u14_u0_n172 ) , .A( u2_u14_u0_n88 ) );
  OAI222_X1 u2_u14_u0_U49 (.C1( u2_u14_u0_n108 ) , .A1( u2_u14_u0_n125 ) , .B2( u2_u14_u0_n128 ) , .B1( u2_u14_u0_n144 ) , .A2( u2_u14_u0_n158 ) , .C2( u2_u14_u0_n161 ) , .ZN( u2_u14_u0_n88 ) );
  AOI21_X1 u2_u14_u0_U5 (.B2( u2_u14_u0_n131 ) , .ZN( u2_u14_u0_n134 ) , .B1( u2_u14_u0_n151 ) , .A( u2_u14_u0_n158 ) );
  NAND2_X1 u2_u14_u0_U50 (.ZN( u2_u14_u0_n112 ) , .A2( u2_u14_u0_n92 ) , .A1( u2_u14_u0_n93 ) );
  OR3_X1 u2_u14_u0_U51 (.A3( u2_u14_u0_n152 ) , .A2( u2_u14_u0_n153 ) , .A1( u2_u14_u0_n154 ) , .ZN( u2_u14_u0_n155 ) );
  AOI21_X1 u2_u14_u0_U52 (.B2( u2_u14_u0_n150 ) , .B1( u2_u14_u0_n151 ) , .ZN( u2_u14_u0_n152 ) , .A( u2_u14_u0_n158 ) );
  AOI21_X1 u2_u14_u0_U53 (.A( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n145 ) , .B1( u2_u14_u0_n146 ) , .ZN( u2_u14_u0_n154 ) );
  AOI21_X1 u2_u14_u0_U54 (.A( u2_u14_u0_n147 ) , .B2( u2_u14_u0_n148 ) , .B1( u2_u14_u0_n149 ) , .ZN( u2_u14_u0_n153 ) );
  INV_X1 u2_u14_u0_U55 (.ZN( u2_u14_u0_n171 ) , .A( u2_u14_u0_n99 ) );
  OAI211_X1 u2_u14_u0_U56 (.C2( u2_u14_u0_n140 ) , .C1( u2_u14_u0_n161 ) , .A( u2_u14_u0_n169 ) , .B( u2_u14_u0_n98 ) , .ZN( u2_u14_u0_n99 ) );
  INV_X1 u2_u14_u0_U57 (.ZN( u2_u14_u0_n169 ) , .A( u2_u14_u0_n91 ) );
  AOI211_X1 u2_u14_u0_U58 (.C1( u2_u14_u0_n118 ) , .A( u2_u14_u0_n123 ) , .B( u2_u14_u0_n96 ) , .C2( u2_u14_u0_n97 ) , .ZN( u2_u14_u0_n98 ) );
  NOR2_X1 u2_u14_u0_U59 (.A2( u2_u14_X_2 ) , .ZN( u2_u14_u0_n103 ) , .A1( u2_u14_u0_n164 ) );
  NOR2_X1 u2_u14_u0_U6 (.A1( u2_u14_u0_n108 ) , .ZN( u2_u14_u0_n123 ) , .A2( u2_u14_u0_n158 ) );
  NOR2_X1 u2_u14_u0_U60 (.A2( u2_u14_X_3 ) , .A1( u2_u14_X_6 ) , .ZN( u2_u14_u0_n94 ) );
  NOR2_X1 u2_u14_u0_U61 (.A2( u2_u14_X_6 ) , .ZN( u2_u14_u0_n100 ) , .A1( u2_u14_u0_n162 ) );
  NOR2_X1 u2_u14_u0_U62 (.A2( u2_u14_X_4 ) , .A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n118 ) );
  NOR2_X1 u2_u14_u0_U63 (.A2( u2_u14_X_1 ) , .A1( u2_u14_X_2 ) , .ZN( u2_u14_u0_n92 ) );
  NOR2_X1 u2_u14_u0_U64 (.A2( u2_u14_X_1 ) , .ZN( u2_u14_u0_n101 ) , .A1( u2_u14_u0_n163 ) );
  NAND2_X1 u2_u14_u0_U65 (.A2( u2_u14_X_4 ) , .A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n144 ) );
  NOR2_X1 u2_u14_u0_U66 (.A2( u2_u14_X_5 ) , .ZN( u2_u14_u0_n136 ) , .A1( u2_u14_u0_n159 ) );
  NAND2_X1 u2_u14_u0_U67 (.A1( u2_u14_X_5 ) , .ZN( u2_u14_u0_n138 ) , .A2( u2_u14_u0_n159 ) );
  AND2_X1 u2_u14_u0_U68 (.A2( u2_u14_X_3 ) , .A1( u2_u14_X_6 ) , .ZN( u2_u14_u0_n102 ) );
  AND2_X1 u2_u14_u0_U69 (.A1( u2_u14_X_6 ) , .A2( u2_u14_u0_n162 ) , .ZN( u2_u14_u0_n93 ) );
  OAI21_X1 u2_u14_u0_U7 (.B1( u2_u14_u0_n150 ) , .B2( u2_u14_u0_n158 ) , .A( u2_u14_u0_n172 ) , .ZN( u2_u14_u0_n89 ) );
  INV_X1 u2_u14_u0_U70 (.A( u2_u14_X_4 ) , .ZN( u2_u14_u0_n159 ) );
  INV_X1 u2_u14_u0_U71 (.A( u2_u14_X_1 ) , .ZN( u2_u14_u0_n164 ) );
  INV_X1 u2_u14_u0_U72 (.A( u2_u14_X_2 ) , .ZN( u2_u14_u0_n163 ) );
  INV_X1 u2_u14_u0_U73 (.A( u2_u14_X_3 ) , .ZN( u2_u14_u0_n162 ) );
  INV_X1 u2_u14_u0_U74 (.A( u2_u14_u0_n126 ) , .ZN( u2_u14_u0_n168 ) );
  AOI211_X1 u2_u14_u0_U75 (.B( u2_u14_u0_n133 ) , .A( u2_u14_u0_n134 ) , .C2( u2_u14_u0_n135 ) , .C1( u2_u14_u0_n136 ) , .ZN( u2_u14_u0_n137 ) );
  INV_X1 u2_u14_u0_U76 (.ZN( u2_u14_u0_n174 ) , .A( u2_u14_u0_n89 ) );
  AOI211_X1 u2_u14_u0_U77 (.B( u2_u14_u0_n104 ) , .A( u2_u14_u0_n105 ) , .ZN( u2_u14_u0_n106 ) , .C2( u2_u14_u0_n113 ) , .C1( u2_u14_u0_n160 ) );
  OR4_X1 u2_u14_u0_U78 (.ZN( u2_out14_17 ) , .A4( u2_u14_u0_n122 ) , .A2( u2_u14_u0_n123 ) , .A1( u2_u14_u0_n124 ) , .A3( u2_u14_u0_n170 ) );
  AOI21_X1 u2_u14_u0_U79 (.B2( u2_u14_u0_n107 ) , .ZN( u2_u14_u0_n124 ) , .B1( u2_u14_u0_n128 ) , .A( u2_u14_u0_n161 ) );
  AND2_X1 u2_u14_u0_U8 (.A1( u2_u14_u0_n114 ) , .A2( u2_u14_u0_n121 ) , .ZN( u2_u14_u0_n146 ) );
  INV_X1 u2_u14_u0_U80 (.A( u2_u14_u0_n111 ) , .ZN( u2_u14_u0_n170 ) );
  OR4_X1 u2_u14_u0_U81 (.ZN( u2_out14_31 ) , .A4( u2_u14_u0_n155 ) , .A2( u2_u14_u0_n156 ) , .A1( u2_u14_u0_n157 ) , .A3( u2_u14_u0_n173 ) );
  AOI21_X1 u2_u14_u0_U82 (.A( u2_u14_u0_n138 ) , .B2( u2_u14_u0_n139 ) , .B1( u2_u14_u0_n140 ) , .ZN( u2_u14_u0_n157 ) );
  AOI21_X1 u2_u14_u0_U83 (.B2( u2_u14_u0_n141 ) , .B1( u2_u14_u0_n142 ) , .ZN( u2_u14_u0_n156 ) , .A( u2_u14_u0_n161 ) );
  AOI21_X1 u2_u14_u0_U84 (.B1( u2_u14_u0_n132 ) , .ZN( u2_u14_u0_n133 ) , .A( u2_u14_u0_n144 ) , .B2( u2_u14_u0_n166 ) );
  OAI22_X1 u2_u14_u0_U85 (.ZN( u2_u14_u0_n105 ) , .A2( u2_u14_u0_n132 ) , .B1( u2_u14_u0_n146 ) , .A1( u2_u14_u0_n147 ) , .B2( u2_u14_u0_n161 ) );
  NAND2_X1 u2_u14_u0_U86 (.ZN( u2_u14_u0_n110 ) , .A2( u2_u14_u0_n132 ) , .A1( u2_u14_u0_n145 ) );
  INV_X1 u2_u14_u0_U87 (.A( u2_u14_u0_n119 ) , .ZN( u2_u14_u0_n167 ) );
  NAND3_X1 u2_u14_u0_U88 (.ZN( u2_out14_23 ) , .A3( u2_u14_u0_n137 ) , .A1( u2_u14_u0_n168 ) , .A2( u2_u14_u0_n171 ) );
  NAND3_X1 u2_u14_u0_U89 (.A3( u2_u14_u0_n127 ) , .A2( u2_u14_u0_n128 ) , .ZN( u2_u14_u0_n135 ) , .A1( u2_u14_u0_n150 ) );
  AND2_X1 u2_u14_u0_U9 (.A1( u2_u14_u0_n131 ) , .ZN( u2_u14_u0_n141 ) , .A2( u2_u14_u0_n150 ) );
  NAND3_X1 u2_u14_u0_U90 (.ZN( u2_u14_u0_n117 ) , .A3( u2_u14_u0_n132 ) , .A2( u2_u14_u0_n139 ) , .A1( u2_u14_u0_n148 ) );
  NAND3_X1 u2_u14_u0_U91 (.ZN( u2_u14_u0_n109 ) , .A2( u2_u14_u0_n114 ) , .A3( u2_u14_u0_n140 ) , .A1( u2_u14_u0_n149 ) );
  NAND3_X1 u2_u14_u0_U92 (.ZN( u2_out14_9 ) , .A3( u2_u14_u0_n106 ) , .A2( u2_u14_u0_n171 ) , .A1( u2_u14_u0_n174 ) );
  NAND3_X1 u2_u14_u0_U93 (.A2( u2_u14_u0_n128 ) , .A1( u2_u14_u0_n132 ) , .A3( u2_u14_u0_n146 ) , .ZN( u2_u14_u0_n97 ) );
  AOI21_X1 u2_u14_u1_U10 (.ZN( u2_u14_u1_n106 ) , .A( u2_u14_u1_n112 ) , .B1( u2_u14_u1_n154 ) , .B2( u2_u14_u1_n156 ) );
  NAND3_X1 u2_u14_u1_U100 (.ZN( u2_u14_u1_n113 ) , .A1( u2_u14_u1_n120 ) , .A3( u2_u14_u1_n133 ) , .A2( u2_u14_u1_n155 ) );
  INV_X1 u2_u14_u1_U11 (.A( u2_u14_u1_n101 ) , .ZN( u2_u14_u1_n184 ) );
  AOI21_X1 u2_u14_u1_U12 (.ZN( u2_u14_u1_n107 ) , .B1( u2_u14_u1_n134 ) , .B2( u2_u14_u1_n149 ) , .A( u2_u14_u1_n174 ) );
  NAND2_X1 u2_u14_u1_U13 (.ZN( u2_u14_u1_n140 ) , .A2( u2_u14_u1_n150 ) , .A1( u2_u14_u1_n155 ) );
  NAND2_X1 u2_u14_u1_U14 (.A1( u2_u14_u1_n131 ) , .ZN( u2_u14_u1_n147 ) , .A2( u2_u14_u1_n153 ) );
  AOI22_X1 u2_u14_u1_U15 (.B2( u2_u14_u1_n136 ) , .A2( u2_u14_u1_n137 ) , .ZN( u2_u14_u1_n143 ) , .A1( u2_u14_u1_n171 ) , .B1( u2_u14_u1_n173 ) );
  INV_X1 u2_u14_u1_U16 (.A( u2_u14_u1_n147 ) , .ZN( u2_u14_u1_n181 ) );
  INV_X1 u2_u14_u1_U17 (.A( u2_u14_u1_n139 ) , .ZN( u2_u14_u1_n174 ) );
  INV_X1 u2_u14_u1_U18 (.A( u2_u14_u1_n112 ) , .ZN( u2_u14_u1_n171 ) );
  NAND2_X1 u2_u14_u1_U19 (.ZN( u2_u14_u1_n141 ) , .A1( u2_u14_u1_n153 ) , .A2( u2_u14_u1_n156 ) );
  AND2_X1 u2_u14_u1_U20 (.A1( u2_u14_u1_n123 ) , .ZN( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n161 ) );
  NAND2_X1 u2_u14_u1_U21 (.A2( u2_u14_u1_n115 ) , .A1( u2_u14_u1_n116 ) , .ZN( u2_u14_u1_n148 ) );
  NAND2_X1 u2_u14_u1_U22 (.A2( u2_u14_u1_n133 ) , .A1( u2_u14_u1_n135 ) , .ZN( u2_u14_u1_n159 ) );
  NAND2_X1 u2_u14_u1_U23 (.A2( u2_u14_u1_n115 ) , .A1( u2_u14_u1_n120 ) , .ZN( u2_u14_u1_n132 ) );
  INV_X1 u2_u14_u1_U24 (.A( u2_u14_u1_n154 ) , .ZN( u2_u14_u1_n178 ) );
  AOI22_X1 u2_u14_u1_U25 (.B2( u2_u14_u1_n113 ) , .A2( u2_u14_u1_n114 ) , .ZN( u2_u14_u1_n125 ) , .A1( u2_u14_u1_n171 ) , .B1( u2_u14_u1_n173 ) );
  NAND2_X1 u2_u14_u1_U26 (.ZN( u2_u14_u1_n114 ) , .A1( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n156 ) );
  INV_X1 u2_u14_u1_U27 (.A( u2_u14_u1_n151 ) , .ZN( u2_u14_u1_n183 ) );
  AND2_X1 u2_u14_u1_U28 (.A1( u2_u14_u1_n129 ) , .A2( u2_u14_u1_n133 ) , .ZN( u2_u14_u1_n149 ) );
  INV_X1 u2_u14_u1_U29 (.A( u2_u14_u1_n131 ) , .ZN( u2_u14_u1_n180 ) );
  INV_X1 u2_u14_u1_U3 (.A( u2_u14_u1_n159 ) , .ZN( u2_u14_u1_n182 ) );
  AOI221_X1 u2_u14_u1_U30 (.B1( u2_u14_u1_n140 ) , .ZN( u2_u14_u1_n167 ) , .B2( u2_u14_u1_n172 ) , .C2( u2_u14_u1_n175 ) , .C1( u2_u14_u1_n178 ) , .A( u2_u14_u1_n188 ) );
  INV_X1 u2_u14_u1_U31 (.ZN( u2_u14_u1_n188 ) , .A( u2_u14_u1_n97 ) );
  AOI211_X1 u2_u14_u1_U32 (.A( u2_u14_u1_n118 ) , .C1( u2_u14_u1_n132 ) , .C2( u2_u14_u1_n139 ) , .B( u2_u14_u1_n96 ) , .ZN( u2_u14_u1_n97 ) );
  AOI21_X1 u2_u14_u1_U33 (.B2( u2_u14_u1_n121 ) , .B1( u2_u14_u1_n135 ) , .A( u2_u14_u1_n152 ) , .ZN( u2_u14_u1_n96 ) );
  OAI221_X1 u2_u14_u1_U34 (.A( u2_u14_u1_n119 ) , .C2( u2_u14_u1_n129 ) , .ZN( u2_u14_u1_n138 ) , .B2( u2_u14_u1_n152 ) , .C1( u2_u14_u1_n174 ) , .B1( u2_u14_u1_n187 ) );
  INV_X1 u2_u14_u1_U35 (.A( u2_u14_u1_n148 ) , .ZN( u2_u14_u1_n187 ) );
  AOI211_X1 u2_u14_u1_U36 (.B( u2_u14_u1_n117 ) , .A( u2_u14_u1_n118 ) , .ZN( u2_u14_u1_n119 ) , .C2( u2_u14_u1_n146 ) , .C1( u2_u14_u1_n159 ) );
  NOR2_X1 u2_u14_u1_U37 (.A1( u2_u14_u1_n168 ) , .A2( u2_u14_u1_n176 ) , .ZN( u2_u14_u1_n98 ) );
  AOI211_X1 u2_u14_u1_U38 (.B( u2_u14_u1_n162 ) , .A( u2_u14_u1_n163 ) , .C2( u2_u14_u1_n164 ) , .ZN( u2_u14_u1_n165 ) , .C1( u2_u14_u1_n171 ) );
  AOI21_X1 u2_u14_u1_U39 (.A( u2_u14_u1_n160 ) , .B2( u2_u14_u1_n161 ) , .ZN( u2_u14_u1_n162 ) , .B1( u2_u14_u1_n182 ) );
  AOI221_X1 u2_u14_u1_U4 (.A( u2_u14_u1_n138 ) , .C2( u2_u14_u1_n139 ) , .C1( u2_u14_u1_n140 ) , .B2( u2_u14_u1_n141 ) , .ZN( u2_u14_u1_n142 ) , .B1( u2_u14_u1_n175 ) );
  OR2_X1 u2_u14_u1_U40 (.A2( u2_u14_u1_n157 ) , .A1( u2_u14_u1_n158 ) , .ZN( u2_u14_u1_n163 ) );
  OAI21_X1 u2_u14_u1_U41 (.B2( u2_u14_u1_n123 ) , .ZN( u2_u14_u1_n145 ) , .B1( u2_u14_u1_n160 ) , .A( u2_u14_u1_n185 ) );
  INV_X1 u2_u14_u1_U42 (.A( u2_u14_u1_n122 ) , .ZN( u2_u14_u1_n185 ) );
  AOI21_X1 u2_u14_u1_U43 (.B2( u2_u14_u1_n120 ) , .B1( u2_u14_u1_n121 ) , .ZN( u2_u14_u1_n122 ) , .A( u2_u14_u1_n128 ) );
  NAND2_X1 u2_u14_u1_U44 (.A1( u2_u14_u1_n128 ) , .ZN( u2_u14_u1_n146 ) , .A2( u2_u14_u1_n160 ) );
  NAND2_X1 u2_u14_u1_U45 (.A2( u2_u14_u1_n112 ) , .ZN( u2_u14_u1_n139 ) , .A1( u2_u14_u1_n152 ) );
  NAND2_X1 u2_u14_u1_U46 (.A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n156 ) , .A2( u2_u14_u1_n99 ) );
  NOR2_X1 u2_u14_u1_U47 (.ZN( u2_u14_u1_n117 ) , .A1( u2_u14_u1_n121 ) , .A2( u2_u14_u1_n160 ) );
  AOI21_X1 u2_u14_u1_U48 (.A( u2_u14_u1_n128 ) , .B2( u2_u14_u1_n129 ) , .ZN( u2_u14_u1_n130 ) , .B1( u2_u14_u1_n150 ) );
  NAND2_X1 u2_u14_u1_U49 (.ZN( u2_u14_u1_n112 ) , .A1( u2_u14_u1_n169 ) , .A2( u2_u14_u1_n170 ) );
  AOI211_X1 u2_u14_u1_U5 (.ZN( u2_u14_u1_n124 ) , .A( u2_u14_u1_n138 ) , .C2( u2_u14_u1_n139 ) , .B( u2_u14_u1_n145 ) , .C1( u2_u14_u1_n147 ) );
  NAND2_X1 u2_u14_u1_U50 (.ZN( u2_u14_u1_n129 ) , .A2( u2_u14_u1_n95 ) , .A1( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U51 (.A1( u2_u14_u1_n102 ) , .ZN( u2_u14_u1_n154 ) , .A2( u2_u14_u1_n99 ) );
  NAND2_X1 u2_u14_u1_U52 (.A2( u2_u14_u1_n100 ) , .ZN( u2_u14_u1_n135 ) , .A1( u2_u14_u1_n99 ) );
  AOI21_X1 u2_u14_u1_U53 (.A( u2_u14_u1_n152 ) , .B2( u2_u14_u1_n153 ) , .B1( u2_u14_u1_n154 ) , .ZN( u2_u14_u1_n158 ) );
  INV_X1 u2_u14_u1_U54 (.A( u2_u14_u1_n160 ) , .ZN( u2_u14_u1_n175 ) );
  NAND2_X1 u2_u14_u1_U55 (.A1( u2_u14_u1_n100 ) , .ZN( u2_u14_u1_n116 ) , .A2( u2_u14_u1_n95 ) );
  NAND2_X1 u2_u14_u1_U56 (.A1( u2_u14_u1_n102 ) , .ZN( u2_u14_u1_n131 ) , .A2( u2_u14_u1_n95 ) );
  NAND2_X1 u2_u14_u1_U57 (.A2( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n121 ) , .A1( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U58 (.A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n153 ) , .A2( u2_u14_u1_n98 ) );
  NAND2_X1 u2_u14_u1_U59 (.A2( u2_u14_u1_n104 ) , .A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n133 ) );
  NOR2_X1 u2_u14_u1_U6 (.A1( u2_u14_u1_n112 ) , .A2( u2_u14_u1_n116 ) , .ZN( u2_u14_u1_n118 ) );
  NAND2_X1 u2_u14_u1_U60 (.ZN( u2_u14_u1_n150 ) , .A2( u2_u14_u1_n98 ) , .A1( u2_u14_u1_n99 ) );
  NAND2_X1 u2_u14_u1_U61 (.A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n155 ) , .A2( u2_u14_u1_n95 ) );
  OAI21_X1 u2_u14_u1_U62 (.ZN( u2_u14_u1_n109 ) , .B1( u2_u14_u1_n129 ) , .B2( u2_u14_u1_n160 ) , .A( u2_u14_u1_n167 ) );
  NAND2_X1 u2_u14_u1_U63 (.A2( u2_u14_u1_n100 ) , .A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n120 ) );
  NAND2_X1 u2_u14_u1_U64 (.A1( u2_u14_u1_n102 ) , .A2( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n115 ) );
  NAND2_X1 u2_u14_u1_U65 (.A2( u2_u14_u1_n100 ) , .A1( u2_u14_u1_n104 ) , .ZN( u2_u14_u1_n151 ) );
  NAND2_X1 u2_u14_u1_U66 (.A2( u2_u14_u1_n103 ) , .A1( u2_u14_u1_n105 ) , .ZN( u2_u14_u1_n161 ) );
  INV_X1 u2_u14_u1_U67 (.A( u2_u14_u1_n152 ) , .ZN( u2_u14_u1_n173 ) );
  INV_X1 u2_u14_u1_U68 (.A( u2_u14_u1_n128 ) , .ZN( u2_u14_u1_n172 ) );
  NAND2_X1 u2_u14_u1_U69 (.A2( u2_u14_u1_n102 ) , .A1( u2_u14_u1_n103 ) , .ZN( u2_u14_u1_n123 ) );
  OAI21_X1 u2_u14_u1_U7 (.ZN( u2_u14_u1_n101 ) , .B1( u2_u14_u1_n141 ) , .A( u2_u14_u1_n146 ) , .B2( u2_u14_u1_n183 ) );
  NOR2_X1 u2_u14_u1_U70 (.A2( u2_u14_X_7 ) , .A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n95 ) );
  NOR2_X1 u2_u14_u1_U71 (.A1( u2_u14_X_12 ) , .A2( u2_u14_X_9 ) , .ZN( u2_u14_u1_n100 ) );
  NOR2_X1 u2_u14_u1_U72 (.A2( u2_u14_X_8 ) , .A1( u2_u14_u1_n177 ) , .ZN( u2_u14_u1_n99 ) );
  NOR2_X1 u2_u14_u1_U73 (.A2( u2_u14_X_12 ) , .ZN( u2_u14_u1_n102 ) , .A1( u2_u14_u1_n176 ) );
  NOR2_X1 u2_u14_u1_U74 (.A2( u2_u14_X_9 ) , .ZN( u2_u14_u1_n105 ) , .A1( u2_u14_u1_n168 ) );
  NAND2_X1 u2_u14_u1_U75 (.A1( u2_u14_X_10 ) , .ZN( u2_u14_u1_n160 ) , .A2( u2_u14_u1_n169 ) );
  NAND2_X1 u2_u14_u1_U76 (.A2( u2_u14_X_10 ) , .A1( u2_u14_X_11 ) , .ZN( u2_u14_u1_n152 ) );
  NAND2_X1 u2_u14_u1_U77 (.A1( u2_u14_X_11 ) , .ZN( u2_u14_u1_n128 ) , .A2( u2_u14_u1_n170 ) );
  AND2_X1 u2_u14_u1_U78 (.A2( u2_u14_X_7 ) , .A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n104 ) );
  AND2_X1 u2_u14_u1_U79 (.A1( u2_u14_X_8 ) , .ZN( u2_u14_u1_n103 ) , .A2( u2_u14_u1_n177 ) );
  AOI21_X1 u2_u14_u1_U8 (.B2( u2_u14_u1_n155 ) , .B1( u2_u14_u1_n156 ) , .ZN( u2_u14_u1_n157 ) , .A( u2_u14_u1_n174 ) );
  INV_X1 u2_u14_u1_U80 (.A( u2_u14_X_10 ) , .ZN( u2_u14_u1_n170 ) );
  INV_X1 u2_u14_u1_U81 (.A( u2_u14_X_9 ) , .ZN( u2_u14_u1_n176 ) );
  INV_X1 u2_u14_u1_U82 (.A( u2_u14_X_11 ) , .ZN( u2_u14_u1_n169 ) );
  INV_X1 u2_u14_u1_U83 (.A( u2_u14_X_12 ) , .ZN( u2_u14_u1_n168 ) );
  INV_X1 u2_u14_u1_U84 (.A( u2_u14_X_7 ) , .ZN( u2_u14_u1_n177 ) );
  NAND4_X1 u2_u14_u1_U85 (.ZN( u2_out14_28 ) , .A4( u2_u14_u1_n124 ) , .A3( u2_u14_u1_n125 ) , .A2( u2_u14_u1_n126 ) , .A1( u2_u14_u1_n127 ) );
  OAI21_X1 u2_u14_u1_U86 (.ZN( u2_u14_u1_n127 ) , .B2( u2_u14_u1_n139 ) , .B1( u2_u14_u1_n175 ) , .A( u2_u14_u1_n183 ) );
  OAI21_X1 u2_u14_u1_U87 (.ZN( u2_u14_u1_n126 ) , .B2( u2_u14_u1_n140 ) , .A( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n178 ) );
  NAND4_X1 u2_u14_u1_U88 (.ZN( u2_out14_18 ) , .A4( u2_u14_u1_n165 ) , .A3( u2_u14_u1_n166 ) , .A1( u2_u14_u1_n167 ) , .A2( u2_u14_u1_n186 ) );
  AOI22_X1 u2_u14_u1_U89 (.B2( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n147 ) , .A2( u2_u14_u1_n148 ) , .ZN( u2_u14_u1_n166 ) , .A1( u2_u14_u1_n172 ) );
  OR4_X1 u2_u14_u1_U9 (.A4( u2_u14_u1_n106 ) , .A3( u2_u14_u1_n107 ) , .ZN( u2_u14_u1_n108 ) , .A1( u2_u14_u1_n117 ) , .A2( u2_u14_u1_n184 ) );
  INV_X1 u2_u14_u1_U90 (.A( u2_u14_u1_n145 ) , .ZN( u2_u14_u1_n186 ) );
  NAND4_X1 u2_u14_u1_U91 (.ZN( u2_out14_2 ) , .A4( u2_u14_u1_n142 ) , .A3( u2_u14_u1_n143 ) , .A2( u2_u14_u1_n144 ) , .A1( u2_u14_u1_n179 ) );
  OAI21_X1 u2_u14_u1_U92 (.B2( u2_u14_u1_n132 ) , .ZN( u2_u14_u1_n144 ) , .A( u2_u14_u1_n146 ) , .B1( u2_u14_u1_n180 ) );
  INV_X1 u2_u14_u1_U93 (.A( u2_u14_u1_n130 ) , .ZN( u2_u14_u1_n179 ) );
  OR4_X1 u2_u14_u1_U94 (.ZN( u2_out14_13 ) , .A4( u2_u14_u1_n108 ) , .A3( u2_u14_u1_n109 ) , .A2( u2_u14_u1_n110 ) , .A1( u2_u14_u1_n111 ) );
  AOI21_X1 u2_u14_u1_U95 (.ZN( u2_u14_u1_n111 ) , .A( u2_u14_u1_n128 ) , .B2( u2_u14_u1_n131 ) , .B1( u2_u14_u1_n135 ) );
  AOI21_X1 u2_u14_u1_U96 (.ZN( u2_u14_u1_n110 ) , .A( u2_u14_u1_n116 ) , .B1( u2_u14_u1_n152 ) , .B2( u2_u14_u1_n160 ) );
  NAND3_X1 u2_u14_u1_U97 (.A3( u2_u14_u1_n149 ) , .A2( u2_u14_u1_n150 ) , .A1( u2_u14_u1_n151 ) , .ZN( u2_u14_u1_n164 ) );
  NAND3_X1 u2_u14_u1_U98 (.A3( u2_u14_u1_n134 ) , .A2( u2_u14_u1_n135 ) , .ZN( u2_u14_u1_n136 ) , .A1( u2_u14_u1_n151 ) );
  NAND3_X1 u2_u14_u1_U99 (.A1( u2_u14_u1_n133 ) , .ZN( u2_u14_u1_n137 ) , .A2( u2_u14_u1_n154 ) , .A3( u2_u14_u1_n181 ) );
  OAI22_X1 u2_u14_u2_U10 (.ZN( u2_u14_u2_n109 ) , .A2( u2_u14_u2_n113 ) , .B2( u2_u14_u2_n133 ) , .B1( u2_u14_u2_n167 ) , .A1( u2_u14_u2_n168 ) );
  NAND3_X1 u2_u14_u2_U100 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n98 ) );
  OAI22_X1 u2_u14_u2_U11 (.B1( u2_u14_u2_n151 ) , .A2( u2_u14_u2_n152 ) , .A1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n160 ) , .B2( u2_u14_u2_n168 ) );
  NOR3_X1 u2_u14_u2_U12 (.A1( u2_u14_u2_n150 ) , .ZN( u2_u14_u2_n151 ) , .A3( u2_u14_u2_n175 ) , .A2( u2_u14_u2_n188 ) );
  AOI21_X1 u2_u14_u2_U13 (.ZN( u2_u14_u2_n144 ) , .B2( u2_u14_u2_n155 ) , .A( u2_u14_u2_n172 ) , .B1( u2_u14_u2_n185 ) );
  AOI21_X1 u2_u14_u2_U14 (.B2( u2_u14_u2_n143 ) , .ZN( u2_u14_u2_n145 ) , .B1( u2_u14_u2_n152 ) , .A( u2_u14_u2_n171 ) );
  AOI21_X1 u2_u14_u2_U15 (.B2( u2_u14_u2_n120 ) , .B1( u2_u14_u2_n121 ) , .ZN( u2_u14_u2_n126 ) , .A( u2_u14_u2_n167 ) );
  INV_X1 u2_u14_u2_U16 (.A( u2_u14_u2_n156 ) , .ZN( u2_u14_u2_n171 ) );
  INV_X1 u2_u14_u2_U17 (.A( u2_u14_u2_n120 ) , .ZN( u2_u14_u2_n188 ) );
  NAND2_X1 u2_u14_u2_U18 (.A2( u2_u14_u2_n122 ) , .ZN( u2_u14_u2_n150 ) , .A1( u2_u14_u2_n152 ) );
  INV_X1 u2_u14_u2_U19 (.A( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n170 ) );
  INV_X1 u2_u14_u2_U20 (.A( u2_u14_u2_n137 ) , .ZN( u2_u14_u2_n173 ) );
  NAND2_X1 u2_u14_u2_U21 (.A1( u2_u14_u2_n132 ) , .A2( u2_u14_u2_n139 ) , .ZN( u2_u14_u2_n157 ) );
  INV_X1 u2_u14_u2_U22 (.A( u2_u14_u2_n113 ) , .ZN( u2_u14_u2_n178 ) );
  INV_X1 u2_u14_u2_U23 (.A( u2_u14_u2_n139 ) , .ZN( u2_u14_u2_n175 ) );
  INV_X1 u2_u14_u2_U24 (.A( u2_u14_u2_n155 ) , .ZN( u2_u14_u2_n181 ) );
  INV_X1 u2_u14_u2_U25 (.A( u2_u14_u2_n119 ) , .ZN( u2_u14_u2_n177 ) );
  INV_X1 u2_u14_u2_U26 (.A( u2_u14_u2_n116 ) , .ZN( u2_u14_u2_n180 ) );
  INV_X1 u2_u14_u2_U27 (.A( u2_u14_u2_n131 ) , .ZN( u2_u14_u2_n179 ) );
  INV_X1 u2_u14_u2_U28 (.A( u2_u14_u2_n154 ) , .ZN( u2_u14_u2_n176 ) );
  NAND2_X1 u2_u14_u2_U29 (.A2( u2_u14_u2_n116 ) , .A1( u2_u14_u2_n117 ) , .ZN( u2_u14_u2_n118 ) );
  NOR2_X1 u2_u14_u2_U3 (.ZN( u2_u14_u2_n121 ) , .A2( u2_u14_u2_n177 ) , .A1( u2_u14_u2_n180 ) );
  INV_X1 u2_u14_u2_U30 (.A( u2_u14_u2_n132 ) , .ZN( u2_u14_u2_n182 ) );
  INV_X1 u2_u14_u2_U31 (.A( u2_u14_u2_n158 ) , .ZN( u2_u14_u2_n183 ) );
  OAI21_X1 u2_u14_u2_U32 (.A( u2_u14_u2_n156 ) , .B1( u2_u14_u2_n157 ) , .ZN( u2_u14_u2_n158 ) , .B2( u2_u14_u2_n179 ) );
  NOR2_X1 u2_u14_u2_U33 (.ZN( u2_u14_u2_n156 ) , .A1( u2_u14_u2_n166 ) , .A2( u2_u14_u2_n169 ) );
  NOR2_X1 u2_u14_u2_U34 (.A2( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n137 ) , .A1( u2_u14_u2_n140 ) );
  NOR2_X1 u2_u14_u2_U35 (.A2( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n153 ) , .A1( u2_u14_u2_n156 ) );
  AOI211_X1 u2_u14_u2_U36 (.ZN( u2_u14_u2_n130 ) , .C1( u2_u14_u2_n138 ) , .C2( u2_u14_u2_n179 ) , .B( u2_u14_u2_n96 ) , .A( u2_u14_u2_n97 ) );
  OAI22_X1 u2_u14_u2_U37 (.B1( u2_u14_u2_n133 ) , .A2( u2_u14_u2_n137 ) , .A1( u2_u14_u2_n152 ) , .B2( u2_u14_u2_n168 ) , .ZN( u2_u14_u2_n97 ) );
  OAI221_X1 u2_u14_u2_U38 (.B1( u2_u14_u2_n113 ) , .C1( u2_u14_u2_n132 ) , .A( u2_u14_u2_n149 ) , .B2( u2_u14_u2_n171 ) , .C2( u2_u14_u2_n172 ) , .ZN( u2_u14_u2_n96 ) );
  OAI221_X1 u2_u14_u2_U39 (.A( u2_u14_u2_n115 ) , .C2( u2_u14_u2_n123 ) , .B2( u2_u14_u2_n143 ) , .B1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n163 ) , .C1( u2_u14_u2_n168 ) );
  INV_X1 u2_u14_u2_U4 (.A( u2_u14_u2_n134 ) , .ZN( u2_u14_u2_n185 ) );
  OAI21_X1 u2_u14_u2_U40 (.A( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n115 ) , .B1( u2_u14_u2_n176 ) , .B2( u2_u14_u2_n178 ) );
  OAI221_X1 u2_u14_u2_U41 (.A( u2_u14_u2_n135 ) , .B2( u2_u14_u2_n136 ) , .B1( u2_u14_u2_n137 ) , .ZN( u2_u14_u2_n162 ) , .C2( u2_u14_u2_n167 ) , .C1( u2_u14_u2_n185 ) );
  AND3_X1 u2_u14_u2_U42 (.A3( u2_u14_u2_n131 ) , .A2( u2_u14_u2_n132 ) , .A1( u2_u14_u2_n133 ) , .ZN( u2_u14_u2_n136 ) );
  AOI22_X1 u2_u14_u2_U43 (.ZN( u2_u14_u2_n135 ) , .B1( u2_u14_u2_n140 ) , .A1( u2_u14_u2_n156 ) , .B2( u2_u14_u2_n180 ) , .A2( u2_u14_u2_n188 ) );
  AOI21_X1 u2_u14_u2_U44 (.ZN( u2_u14_u2_n149 ) , .B1( u2_u14_u2_n173 ) , .B2( u2_u14_u2_n188 ) , .A( u2_u14_u2_n95 ) );
  AND3_X1 u2_u14_u2_U45 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n156 ) , .ZN( u2_u14_u2_n95 ) );
  OAI21_X1 u2_u14_u2_U46 (.A( u2_u14_u2_n141 ) , .B2( u2_u14_u2_n142 ) , .ZN( u2_u14_u2_n146 ) , .B1( u2_u14_u2_n153 ) );
  OAI21_X1 u2_u14_u2_U47 (.A( u2_u14_u2_n140 ) , .ZN( u2_u14_u2_n141 ) , .B1( u2_u14_u2_n176 ) , .B2( u2_u14_u2_n177 ) );
  NOR3_X1 u2_u14_u2_U48 (.ZN( u2_u14_u2_n142 ) , .A3( u2_u14_u2_n175 ) , .A2( u2_u14_u2_n178 ) , .A1( u2_u14_u2_n181 ) );
  OAI21_X1 u2_u14_u2_U49 (.A( u2_u14_u2_n101 ) , .B2( u2_u14_u2_n121 ) , .B1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n164 ) );
  INV_X1 u2_u14_u2_U5 (.A( u2_u14_u2_n150 ) , .ZN( u2_u14_u2_n184 ) );
  NAND2_X1 u2_u14_u2_U50 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n155 ) );
  NAND2_X1 u2_u14_u2_U51 (.A2( u2_u14_u2_n105 ) , .A1( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n143 ) );
  NAND2_X1 u2_u14_u2_U52 (.A1( u2_u14_u2_n104 ) , .A2( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n152 ) );
  NAND2_X1 u2_u14_u2_U53 (.A1( u2_u14_u2_n100 ) , .A2( u2_u14_u2_n105 ) , .ZN( u2_u14_u2_n132 ) );
  INV_X1 u2_u14_u2_U54 (.A( u2_u14_u2_n140 ) , .ZN( u2_u14_u2_n168 ) );
  INV_X1 u2_u14_u2_U55 (.A( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n167 ) );
  INV_X1 u2_u14_u2_U56 (.ZN( u2_u14_u2_n187 ) , .A( u2_u14_u2_n99 ) );
  OAI21_X1 u2_u14_u2_U57 (.B1( u2_u14_u2_n137 ) , .B2( u2_u14_u2_n143 ) , .A( u2_u14_u2_n98 ) , .ZN( u2_u14_u2_n99 ) );
  NAND2_X1 u2_u14_u2_U58 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n113 ) );
  NAND2_X1 u2_u14_u2_U59 (.A1( u2_u14_u2_n106 ) , .A2( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n131 ) );
  NOR4_X1 u2_u14_u2_U6 (.A4( u2_u14_u2_n124 ) , .A3( u2_u14_u2_n125 ) , .A2( u2_u14_u2_n126 ) , .A1( u2_u14_u2_n127 ) , .ZN( u2_u14_u2_n128 ) );
  NAND2_X1 u2_u14_u2_U60 (.A1( u2_u14_u2_n103 ) , .A2( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n139 ) );
  NAND2_X1 u2_u14_u2_U61 (.A1( u2_u14_u2_n103 ) , .A2( u2_u14_u2_n105 ) , .ZN( u2_u14_u2_n133 ) );
  NAND2_X1 u2_u14_u2_U62 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n103 ) , .ZN( u2_u14_u2_n154 ) );
  NAND2_X1 u2_u14_u2_U63 (.A2( u2_u14_u2_n103 ) , .A1( u2_u14_u2_n104 ) , .ZN( u2_u14_u2_n119 ) );
  NAND2_X1 u2_u14_u2_U64 (.A2( u2_u14_u2_n107 ) , .A1( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n123 ) );
  NAND2_X1 u2_u14_u2_U65 (.A1( u2_u14_u2_n104 ) , .A2( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n122 ) );
  INV_X1 u2_u14_u2_U66 (.A( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n172 ) );
  NAND2_X1 u2_u14_u2_U67 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n102 ) , .ZN( u2_u14_u2_n116 ) );
  NAND2_X1 u2_u14_u2_U68 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n120 ) );
  NAND2_X1 u2_u14_u2_U69 (.A2( u2_u14_u2_n105 ) , .A1( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n117 ) );
  AOI21_X1 u2_u14_u2_U7 (.B2( u2_u14_u2_n119 ) , .ZN( u2_u14_u2_n127 ) , .A( u2_u14_u2_n137 ) , .B1( u2_u14_u2_n155 ) );
  NOR2_X1 u2_u14_u2_U70 (.A2( u2_u14_X_16 ) , .ZN( u2_u14_u2_n140 ) , .A1( u2_u14_u2_n166 ) );
  NOR2_X1 u2_u14_u2_U71 (.A2( u2_u14_X_13 ) , .A1( u2_u14_X_14 ) , .ZN( u2_u14_u2_n100 ) );
  NOR2_X1 u2_u14_u2_U72 (.A2( u2_u14_X_16 ) , .A1( u2_u14_X_17 ) , .ZN( u2_u14_u2_n138 ) );
  NOR2_X1 u2_u14_u2_U73 (.A2( u2_u14_X_15 ) , .A1( u2_u14_X_18 ) , .ZN( u2_u14_u2_n104 ) );
  NOR2_X1 u2_u14_u2_U74 (.A2( u2_u14_X_14 ) , .ZN( u2_u14_u2_n103 ) , .A1( u2_u14_u2_n174 ) );
  NOR2_X1 u2_u14_u2_U75 (.A2( u2_u14_X_15 ) , .ZN( u2_u14_u2_n102 ) , .A1( u2_u14_u2_n165 ) );
  NOR2_X1 u2_u14_u2_U76 (.A2( u2_u14_X_17 ) , .ZN( u2_u14_u2_n114 ) , .A1( u2_u14_u2_n169 ) );
  AND2_X1 u2_u14_u2_U77 (.A1( u2_u14_X_15 ) , .ZN( u2_u14_u2_n105 ) , .A2( u2_u14_u2_n165 ) );
  AND2_X1 u2_u14_u2_U78 (.A2( u2_u14_X_15 ) , .A1( u2_u14_X_18 ) , .ZN( u2_u14_u2_n107 ) );
  AND2_X1 u2_u14_u2_U79 (.A1( u2_u14_X_14 ) , .ZN( u2_u14_u2_n106 ) , .A2( u2_u14_u2_n174 ) );
  AOI21_X1 u2_u14_u2_U8 (.ZN( u2_u14_u2_n124 ) , .B1( u2_u14_u2_n131 ) , .B2( u2_u14_u2_n143 ) , .A( u2_u14_u2_n172 ) );
  AND2_X1 u2_u14_u2_U80 (.A1( u2_u14_X_13 ) , .A2( u2_u14_X_14 ) , .ZN( u2_u14_u2_n108 ) );
  INV_X1 u2_u14_u2_U81 (.A( u2_u14_X_16 ) , .ZN( u2_u14_u2_n169 ) );
  INV_X1 u2_u14_u2_U82 (.A( u2_u14_X_17 ) , .ZN( u2_u14_u2_n166 ) );
  INV_X1 u2_u14_u2_U83 (.A( u2_u14_X_13 ) , .ZN( u2_u14_u2_n174 ) );
  INV_X1 u2_u14_u2_U84 (.A( u2_u14_X_18 ) , .ZN( u2_u14_u2_n165 ) );
  NAND4_X1 u2_u14_u2_U85 (.ZN( u2_out14_30 ) , .A4( u2_u14_u2_n147 ) , .A3( u2_u14_u2_n148 ) , .A2( u2_u14_u2_n149 ) , .A1( u2_u14_u2_n187 ) );
  NOR3_X1 u2_u14_u2_U86 (.A3( u2_u14_u2_n144 ) , .A2( u2_u14_u2_n145 ) , .A1( u2_u14_u2_n146 ) , .ZN( u2_u14_u2_n147 ) );
  AOI21_X1 u2_u14_u2_U87 (.B2( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n148 ) , .A( u2_u14_u2_n162 ) , .B1( u2_u14_u2_n182 ) );
  NAND4_X1 u2_u14_u2_U88 (.ZN( u2_out14_24 ) , .A4( u2_u14_u2_n111 ) , .A3( u2_u14_u2_n112 ) , .A1( u2_u14_u2_n130 ) , .A2( u2_u14_u2_n187 ) );
  AOI221_X1 u2_u14_u2_U89 (.A( u2_u14_u2_n109 ) , .B1( u2_u14_u2_n110 ) , .ZN( u2_u14_u2_n111 ) , .C1( u2_u14_u2_n134 ) , .C2( u2_u14_u2_n170 ) , .B2( u2_u14_u2_n173 ) );
  AOI21_X1 u2_u14_u2_U9 (.B2( u2_u14_u2_n123 ) , .ZN( u2_u14_u2_n125 ) , .A( u2_u14_u2_n171 ) , .B1( u2_u14_u2_n184 ) );
  AOI21_X1 u2_u14_u2_U90 (.ZN( u2_u14_u2_n112 ) , .B2( u2_u14_u2_n156 ) , .A( u2_u14_u2_n164 ) , .B1( u2_u14_u2_n181 ) );
  NAND4_X1 u2_u14_u2_U91 (.ZN( u2_out14_16 ) , .A4( u2_u14_u2_n128 ) , .A3( u2_u14_u2_n129 ) , .A1( u2_u14_u2_n130 ) , .A2( u2_u14_u2_n186 ) );
  AOI22_X1 u2_u14_u2_U92 (.A2( u2_u14_u2_n118 ) , .ZN( u2_u14_u2_n129 ) , .A1( u2_u14_u2_n140 ) , .B1( u2_u14_u2_n157 ) , .B2( u2_u14_u2_n170 ) );
  INV_X1 u2_u14_u2_U93 (.A( u2_u14_u2_n163 ) , .ZN( u2_u14_u2_n186 ) );
  OR4_X1 u2_u14_u2_U94 (.ZN( u2_out14_6 ) , .A4( u2_u14_u2_n161 ) , .A3( u2_u14_u2_n162 ) , .A2( u2_u14_u2_n163 ) , .A1( u2_u14_u2_n164 ) );
  OR3_X1 u2_u14_u2_U95 (.A2( u2_u14_u2_n159 ) , .A1( u2_u14_u2_n160 ) , .ZN( u2_u14_u2_n161 ) , .A3( u2_u14_u2_n183 ) );
  AOI21_X1 u2_u14_u2_U96 (.B2( u2_u14_u2_n154 ) , .B1( u2_u14_u2_n155 ) , .ZN( u2_u14_u2_n159 ) , .A( u2_u14_u2_n167 ) );
  NAND3_X1 u2_u14_u2_U97 (.A2( u2_u14_u2_n117 ) , .A1( u2_u14_u2_n122 ) , .A3( u2_u14_u2_n123 ) , .ZN( u2_u14_u2_n134 ) );
  NAND3_X1 u2_u14_u2_U98 (.ZN( u2_u14_u2_n110 ) , .A2( u2_u14_u2_n131 ) , .A3( u2_u14_u2_n139 ) , .A1( u2_u14_u2_n154 ) );
  NAND3_X1 u2_u14_u2_U99 (.A2( u2_u14_u2_n100 ) , .ZN( u2_u14_u2_n101 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n114 ) );
  OAI22_X1 u2_u14_u3_U10 (.B1( u2_u14_u3_n113 ) , .A2( u2_u14_u3_n135 ) , .A1( u2_u14_u3_n150 ) , .B2( u2_u14_u3_n164 ) , .ZN( u2_u14_u3_n98 ) );
  OAI211_X1 u2_u14_u3_U11 (.B( u2_u14_u3_n106 ) , .ZN( u2_u14_u3_n119 ) , .C2( u2_u14_u3_n128 ) , .C1( u2_u14_u3_n167 ) , .A( u2_u14_u3_n181 ) );
  AOI221_X1 u2_u14_u3_U12 (.C1( u2_u14_u3_n105 ) , .ZN( u2_u14_u3_n106 ) , .A( u2_u14_u3_n131 ) , .B2( u2_u14_u3_n132 ) , .C2( u2_u14_u3_n133 ) , .B1( u2_u14_u3_n169 ) );
  INV_X1 u2_u14_u3_U13 (.ZN( u2_u14_u3_n181 ) , .A( u2_u14_u3_n98 ) );
  NAND2_X1 u2_u14_u3_U14 (.ZN( u2_u14_u3_n105 ) , .A2( u2_u14_u3_n130 ) , .A1( u2_u14_u3_n155 ) );
  AOI22_X1 u2_u14_u3_U15 (.B1( u2_u14_u3_n115 ) , .A2( u2_u14_u3_n116 ) , .ZN( u2_u14_u3_n123 ) , .B2( u2_u14_u3_n133 ) , .A1( u2_u14_u3_n169 ) );
  NAND2_X1 u2_u14_u3_U16 (.ZN( u2_u14_u3_n116 ) , .A2( u2_u14_u3_n151 ) , .A1( u2_u14_u3_n182 ) );
  NOR2_X1 u2_u14_u3_U17 (.ZN( u2_u14_u3_n126 ) , .A2( u2_u14_u3_n150 ) , .A1( u2_u14_u3_n164 ) );
  AOI21_X1 u2_u14_u3_U18 (.ZN( u2_u14_u3_n112 ) , .B2( u2_u14_u3_n146 ) , .B1( u2_u14_u3_n155 ) , .A( u2_u14_u3_n167 ) );
  NAND2_X1 u2_u14_u3_U19 (.A1( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n142 ) , .A2( u2_u14_u3_n164 ) );
  NAND2_X1 u2_u14_u3_U20 (.ZN( u2_u14_u3_n132 ) , .A2( u2_u14_u3_n152 ) , .A1( u2_u14_u3_n156 ) );
  AND2_X1 u2_u14_u3_U21 (.A2( u2_u14_u3_n113 ) , .A1( u2_u14_u3_n114 ) , .ZN( u2_u14_u3_n151 ) );
  INV_X1 u2_u14_u3_U22 (.A( u2_u14_u3_n133 ) , .ZN( u2_u14_u3_n165 ) );
  INV_X1 u2_u14_u3_U23 (.A( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n170 ) );
  NAND2_X1 u2_u14_u3_U24 (.A1( u2_u14_u3_n107 ) , .A2( u2_u14_u3_n108 ) , .ZN( u2_u14_u3_n140 ) );
  NAND2_X1 u2_u14_u3_U25 (.ZN( u2_u14_u3_n117 ) , .A1( u2_u14_u3_n124 ) , .A2( u2_u14_u3_n148 ) );
  NAND2_X1 u2_u14_u3_U26 (.ZN( u2_u14_u3_n143 ) , .A1( u2_u14_u3_n165 ) , .A2( u2_u14_u3_n167 ) );
  INV_X1 u2_u14_u3_U27 (.A( u2_u14_u3_n130 ) , .ZN( u2_u14_u3_n177 ) );
  INV_X1 u2_u14_u3_U28 (.A( u2_u14_u3_n128 ) , .ZN( u2_u14_u3_n176 ) );
  INV_X1 u2_u14_u3_U29 (.A( u2_u14_u3_n155 ) , .ZN( u2_u14_u3_n174 ) );
  INV_X1 u2_u14_u3_U3 (.A( u2_u14_u3_n129 ) , .ZN( u2_u14_u3_n183 ) );
  INV_X1 u2_u14_u3_U30 (.A( u2_u14_u3_n139 ) , .ZN( u2_u14_u3_n185 ) );
  NOR2_X1 u2_u14_u3_U31 (.ZN( u2_u14_u3_n135 ) , .A2( u2_u14_u3_n141 ) , .A1( u2_u14_u3_n169 ) );
  OAI222_X1 u2_u14_u3_U32 (.C2( u2_u14_u3_n107 ) , .A2( u2_u14_u3_n108 ) , .B1( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n138 ) , .B2( u2_u14_u3_n146 ) , .C1( u2_u14_u3_n154 ) , .A1( u2_u14_u3_n164 ) );
  NOR4_X1 u2_u14_u3_U33 (.A4( u2_u14_u3_n157 ) , .A3( u2_u14_u3_n158 ) , .A2( u2_u14_u3_n159 ) , .A1( u2_u14_u3_n160 ) , .ZN( u2_u14_u3_n161 ) );
  AOI21_X1 u2_u14_u3_U34 (.B2( u2_u14_u3_n152 ) , .B1( u2_u14_u3_n153 ) , .ZN( u2_u14_u3_n158 ) , .A( u2_u14_u3_n164 ) );
  AOI21_X1 u2_u14_u3_U35 (.A( u2_u14_u3_n154 ) , .B2( u2_u14_u3_n155 ) , .B1( u2_u14_u3_n156 ) , .ZN( u2_u14_u3_n157 ) );
  AOI21_X1 u2_u14_u3_U36 (.A( u2_u14_u3_n149 ) , .B2( u2_u14_u3_n150 ) , .B1( u2_u14_u3_n151 ) , .ZN( u2_u14_u3_n159 ) );
  AOI211_X1 u2_u14_u3_U37 (.ZN( u2_u14_u3_n109 ) , .A( u2_u14_u3_n119 ) , .C2( u2_u14_u3_n129 ) , .B( u2_u14_u3_n138 ) , .C1( u2_u14_u3_n141 ) );
  AOI211_X1 u2_u14_u3_U38 (.B( u2_u14_u3_n119 ) , .A( u2_u14_u3_n120 ) , .C2( u2_u14_u3_n121 ) , .ZN( u2_u14_u3_n122 ) , .C1( u2_u14_u3_n179 ) );
  INV_X1 u2_u14_u3_U39 (.A( u2_u14_u3_n156 ) , .ZN( u2_u14_u3_n179 ) );
  INV_X1 u2_u14_u3_U4 (.A( u2_u14_u3_n140 ) , .ZN( u2_u14_u3_n182 ) );
  OAI22_X1 u2_u14_u3_U40 (.B1( u2_u14_u3_n118 ) , .ZN( u2_u14_u3_n120 ) , .A1( u2_u14_u3_n135 ) , .B2( u2_u14_u3_n154 ) , .A2( u2_u14_u3_n178 ) );
  AND3_X1 u2_u14_u3_U41 (.ZN( u2_u14_u3_n118 ) , .A2( u2_u14_u3_n124 ) , .A1( u2_u14_u3_n144 ) , .A3( u2_u14_u3_n152 ) );
  INV_X1 u2_u14_u3_U42 (.A( u2_u14_u3_n121 ) , .ZN( u2_u14_u3_n164 ) );
  NAND2_X1 u2_u14_u3_U43 (.ZN( u2_u14_u3_n133 ) , .A1( u2_u14_u3_n154 ) , .A2( u2_u14_u3_n164 ) );
  OAI211_X1 u2_u14_u3_U44 (.B( u2_u14_u3_n127 ) , .ZN( u2_u14_u3_n139 ) , .C1( u2_u14_u3_n150 ) , .C2( u2_u14_u3_n154 ) , .A( u2_u14_u3_n184 ) );
  INV_X1 u2_u14_u3_U45 (.A( u2_u14_u3_n125 ) , .ZN( u2_u14_u3_n184 ) );
  AOI221_X1 u2_u14_u3_U46 (.A( u2_u14_u3_n126 ) , .ZN( u2_u14_u3_n127 ) , .C2( u2_u14_u3_n132 ) , .C1( u2_u14_u3_n169 ) , .B2( u2_u14_u3_n170 ) , .B1( u2_u14_u3_n174 ) );
  OAI22_X1 u2_u14_u3_U47 (.A1( u2_u14_u3_n124 ) , .ZN( u2_u14_u3_n125 ) , .B2( u2_u14_u3_n145 ) , .A2( u2_u14_u3_n165 ) , .B1( u2_u14_u3_n167 ) );
  NOR2_X1 u2_u14_u3_U48 (.A1( u2_u14_u3_n113 ) , .ZN( u2_u14_u3_n131 ) , .A2( u2_u14_u3_n154 ) );
  NAND2_X1 u2_u14_u3_U49 (.A1( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n150 ) , .A2( u2_u14_u3_n99 ) );
  INV_X1 u2_u14_u3_U5 (.A( u2_u14_u3_n117 ) , .ZN( u2_u14_u3_n178 ) );
  NAND2_X1 u2_u14_u3_U50 (.A2( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n155 ) , .A1( u2_u14_u3_n97 ) );
  INV_X1 u2_u14_u3_U51 (.A( u2_u14_u3_n141 ) , .ZN( u2_u14_u3_n167 ) );
  AOI21_X1 u2_u14_u3_U52 (.B2( u2_u14_u3_n114 ) , .B1( u2_u14_u3_n146 ) , .A( u2_u14_u3_n154 ) , .ZN( u2_u14_u3_n94 ) );
  AOI21_X1 u2_u14_u3_U53 (.ZN( u2_u14_u3_n110 ) , .B2( u2_u14_u3_n142 ) , .B1( u2_u14_u3_n186 ) , .A( u2_u14_u3_n95 ) );
  INV_X1 u2_u14_u3_U54 (.A( u2_u14_u3_n145 ) , .ZN( u2_u14_u3_n186 ) );
  AOI21_X1 u2_u14_u3_U55 (.B1( u2_u14_u3_n124 ) , .A( u2_u14_u3_n149 ) , .B2( u2_u14_u3_n155 ) , .ZN( u2_u14_u3_n95 ) );
  INV_X1 u2_u14_u3_U56 (.A( u2_u14_u3_n149 ) , .ZN( u2_u14_u3_n169 ) );
  NAND2_X1 u2_u14_u3_U57 (.ZN( u2_u14_u3_n124 ) , .A1( u2_u14_u3_n96 ) , .A2( u2_u14_u3_n97 ) );
  NAND2_X1 u2_u14_u3_U58 (.A2( u2_u14_u3_n100 ) , .ZN( u2_u14_u3_n146 ) , .A1( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U59 (.A1( u2_u14_u3_n101 ) , .ZN( u2_u14_u3_n145 ) , .A2( u2_u14_u3_n99 ) );
  AOI221_X1 u2_u14_u3_U6 (.A( u2_u14_u3_n131 ) , .C2( u2_u14_u3_n132 ) , .C1( u2_u14_u3_n133 ) , .ZN( u2_u14_u3_n134 ) , .B1( u2_u14_u3_n143 ) , .B2( u2_u14_u3_n177 ) );
  NAND2_X1 u2_u14_u3_U60 (.A1( u2_u14_u3_n100 ) , .ZN( u2_u14_u3_n156 ) , .A2( u2_u14_u3_n99 ) );
  NAND2_X1 u2_u14_u3_U61 (.A2( u2_u14_u3_n101 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n148 ) );
  NAND2_X1 u2_u14_u3_U62 (.A1( u2_u14_u3_n100 ) , .A2( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n128 ) );
  NAND2_X1 u2_u14_u3_U63 (.A2( u2_u14_u3_n101 ) , .A1( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n152 ) );
  NAND2_X1 u2_u14_u3_U64 (.A2( u2_u14_u3_n101 ) , .ZN( u2_u14_u3_n114 ) , .A1( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U65 (.ZN( u2_u14_u3_n107 ) , .A1( u2_u14_u3_n97 ) , .A2( u2_u14_u3_n99 ) );
  NAND2_X1 u2_u14_u3_U66 (.A2( u2_u14_u3_n100 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n113 ) );
  NAND2_X1 u2_u14_u3_U67 (.A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n153 ) , .A2( u2_u14_u3_n97 ) );
  NAND2_X1 u2_u14_u3_U68 (.A2( u2_u14_u3_n103 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n130 ) );
  NAND2_X1 u2_u14_u3_U69 (.A2( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n144 ) , .A1( u2_u14_u3_n96 ) );
  OAI22_X1 u2_u14_u3_U7 (.B2( u2_u14_u3_n147 ) , .A2( u2_u14_u3_n148 ) , .ZN( u2_u14_u3_n160 ) , .B1( u2_u14_u3_n165 ) , .A1( u2_u14_u3_n168 ) );
  NAND2_X1 u2_u14_u3_U70 (.A1( u2_u14_u3_n102 ) , .A2( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n108 ) );
  NOR2_X1 u2_u14_u3_U71 (.A2( u2_u14_X_19 ) , .A1( u2_u14_X_20 ) , .ZN( u2_u14_u3_n99 ) );
  NOR2_X1 u2_u14_u3_U72 (.A2( u2_u14_X_21 ) , .A1( u2_u14_X_24 ) , .ZN( u2_u14_u3_n103 ) );
  NOR2_X1 u2_u14_u3_U73 (.A2( u2_u14_X_24 ) , .A1( u2_u14_u3_n171 ) , .ZN( u2_u14_u3_n97 ) );
  NOR2_X1 u2_u14_u3_U74 (.A2( u2_u14_X_23 ) , .ZN( u2_u14_u3_n141 ) , .A1( u2_u14_u3_n166 ) );
  NOR2_X1 u2_u14_u3_U75 (.A2( u2_u14_X_19 ) , .A1( u2_u14_u3_n172 ) , .ZN( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U76 (.A1( u2_u14_X_22 ) , .A2( u2_u14_X_23 ) , .ZN( u2_u14_u3_n154 ) );
  NAND2_X1 u2_u14_u3_U77 (.A1( u2_u14_X_23 ) , .ZN( u2_u14_u3_n149 ) , .A2( u2_u14_u3_n166 ) );
  NOR2_X1 u2_u14_u3_U78 (.A2( u2_u14_X_22 ) , .A1( u2_u14_X_23 ) , .ZN( u2_u14_u3_n121 ) );
  AND2_X1 u2_u14_u3_U79 (.A1( u2_u14_X_24 ) , .ZN( u2_u14_u3_n101 ) , .A2( u2_u14_u3_n171 ) );
  AND3_X1 u2_u14_u3_U8 (.A3( u2_u14_u3_n144 ) , .A2( u2_u14_u3_n145 ) , .A1( u2_u14_u3_n146 ) , .ZN( u2_u14_u3_n147 ) );
  AND2_X1 u2_u14_u3_U80 (.A1( u2_u14_X_19 ) , .ZN( u2_u14_u3_n102 ) , .A2( u2_u14_u3_n172 ) );
  AND2_X1 u2_u14_u3_U81 (.A1( u2_u14_X_21 ) , .A2( u2_u14_X_24 ) , .ZN( u2_u14_u3_n100 ) );
  AND2_X1 u2_u14_u3_U82 (.A2( u2_u14_X_19 ) , .A1( u2_u14_X_20 ) , .ZN( u2_u14_u3_n104 ) );
  INV_X1 u2_u14_u3_U83 (.A( u2_u14_X_22 ) , .ZN( u2_u14_u3_n166 ) );
  INV_X1 u2_u14_u3_U84 (.A( u2_u14_X_21 ) , .ZN( u2_u14_u3_n171 ) );
  INV_X1 u2_u14_u3_U85 (.A( u2_u14_X_20 ) , .ZN( u2_u14_u3_n172 ) );
  NAND4_X1 u2_u14_u3_U86 (.ZN( u2_out14_26 ) , .A4( u2_u14_u3_n109 ) , .A3( u2_u14_u3_n110 ) , .A2( u2_u14_u3_n111 ) , .A1( u2_u14_u3_n173 ) );
  INV_X1 u2_u14_u3_U87 (.ZN( u2_u14_u3_n173 ) , .A( u2_u14_u3_n94 ) );
  OAI21_X1 u2_u14_u3_U88 (.ZN( u2_u14_u3_n111 ) , .B2( u2_u14_u3_n117 ) , .A( u2_u14_u3_n133 ) , .B1( u2_u14_u3_n176 ) );
  NAND4_X1 u2_u14_u3_U89 (.ZN( u2_out14_20 ) , .A4( u2_u14_u3_n122 ) , .A3( u2_u14_u3_n123 ) , .A1( u2_u14_u3_n175 ) , .A2( u2_u14_u3_n180 ) );
  INV_X1 u2_u14_u3_U9 (.A( u2_u14_u3_n143 ) , .ZN( u2_u14_u3_n168 ) );
  INV_X1 u2_u14_u3_U90 (.A( u2_u14_u3_n126 ) , .ZN( u2_u14_u3_n180 ) );
  INV_X1 u2_u14_u3_U91 (.A( u2_u14_u3_n112 ) , .ZN( u2_u14_u3_n175 ) );
  NAND4_X1 u2_u14_u3_U92 (.ZN( u2_out14_1 ) , .A4( u2_u14_u3_n161 ) , .A3( u2_u14_u3_n162 ) , .A2( u2_u14_u3_n163 ) , .A1( u2_u14_u3_n185 ) );
  NAND2_X1 u2_u14_u3_U93 (.ZN( u2_u14_u3_n163 ) , .A2( u2_u14_u3_n170 ) , .A1( u2_u14_u3_n176 ) );
  AOI22_X1 u2_u14_u3_U94 (.B2( u2_u14_u3_n140 ) , .B1( u2_u14_u3_n141 ) , .A2( u2_u14_u3_n142 ) , .ZN( u2_u14_u3_n162 ) , .A1( u2_u14_u3_n177 ) );
  OR4_X1 u2_u14_u3_U95 (.ZN( u2_out14_10 ) , .A4( u2_u14_u3_n136 ) , .A3( u2_u14_u3_n137 ) , .A1( u2_u14_u3_n138 ) , .A2( u2_u14_u3_n139 ) );
  OAI222_X1 u2_u14_u3_U96 (.C1( u2_u14_u3_n128 ) , .ZN( u2_u14_u3_n137 ) , .B1( u2_u14_u3_n148 ) , .A2( u2_u14_u3_n150 ) , .B2( u2_u14_u3_n154 ) , .C2( u2_u14_u3_n164 ) , .A1( u2_u14_u3_n167 ) );
  OAI221_X1 u2_u14_u3_U97 (.A( u2_u14_u3_n134 ) , .B2( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n136 ) , .C1( u2_u14_u3_n149 ) , .B1( u2_u14_u3_n151 ) , .C2( u2_u14_u3_n183 ) );
  NAND3_X1 u2_u14_u3_U98 (.A1( u2_u14_u3_n114 ) , .ZN( u2_u14_u3_n115 ) , .A2( u2_u14_u3_n145 ) , .A3( u2_u14_u3_n153 ) );
  NAND3_X1 u2_u14_u3_U99 (.ZN( u2_u14_u3_n129 ) , .A2( u2_u14_u3_n144 ) , .A1( u2_u14_u3_n153 ) , .A3( u2_u14_u3_n182 ) );
  XOR2_X1 u2_u15_U1 (.A( u2_FP_38 ) , .B( u2_K16_9 ) , .Z( u2_u15_X_9 ) );
  XOR2_X1 u2_u15_U16 (.A( u2_FP_34 ) , .B( u2_K16_3 ) , .Z( u2_u15_X_3 ) );
  XOR2_X1 u2_u15_U2 (.A( u2_FP_37 ) , .B( u2_K16_8 ) , .Z( u2_u15_X_8 ) );
  XOR2_X1 u2_u15_U27 (.A( u2_FP_33 ) , .B( u2_K16_2 ) , .Z( u2_u15_X_2 ) );
  XOR2_X1 u2_u15_U3 (.A( u2_FP_36 ) , .B( u2_K16_7 ) , .Z( u2_u15_X_7 ) );
  XOR2_X1 u2_u15_U33 (.A( u2_FP_49 ) , .B( u2_K16_24 ) , .Z( u2_u15_X_24 ) );
  XOR2_X1 u2_u15_U34 (.A( u2_FP_48 ) , .B( u2_K16_23 ) , .Z( u2_u15_X_23 ) );
  XOR2_X1 u2_u15_U35 (.A( u2_FP_47 ) , .B( u2_K16_22 ) , .Z( u2_u15_X_22 ) );
  XOR2_X1 u2_u15_U36 (.A( u2_FP_46 ) , .B( u2_K16_21 ) , .Z( u2_u15_X_21 ) );
  XOR2_X1 u2_u15_U37 (.A( u2_FP_45 ) , .B( u2_K16_20 ) , .Z( u2_u15_X_20 ) );
  XOR2_X1 u2_u15_U38 (.A( u2_FP_64 ) , .B( u2_K16_1 ) , .Z( u2_u15_X_1 ) );
  XOR2_X1 u2_u15_U39 (.A( u2_FP_44 ) , .B( u2_K16_19 ) , .Z( u2_u15_X_19 ) );
  XOR2_X1 u2_u15_U4 (.A( u2_FP_37 ) , .B( u2_K16_6 ) , .Z( u2_u15_X_6 ) );
  XOR2_X1 u2_u15_U40 (.A( u2_FP_45 ) , .B( u2_K16_18 ) , .Z( u2_u15_X_18 ) );
  XOR2_X1 u2_u15_U41 (.A( u2_FP_44 ) , .B( u2_K16_17 ) , .Z( u2_u15_X_17 ) );
  XOR2_X1 u2_u15_U42 (.A( u2_FP_43 ) , .B( u2_K16_16 ) , .Z( u2_u15_X_16 ) );
  XOR2_X1 u2_u15_U43 (.A( u2_FP_42 ) , .B( u2_K16_15 ) , .Z( u2_u15_X_15 ) );
  XOR2_X1 u2_u15_U44 (.A( u2_FP_41 ) , .B( u2_K16_14 ) , .Z( u2_u15_X_14 ) );
  XOR2_X1 u2_u15_U45 (.A( u2_FP_40 ) , .B( u2_K16_13 ) , .Z( u2_u15_X_13 ) );
  XOR2_X1 u2_u15_U46 (.A( u2_FP_41 ) , .B( u2_K16_12 ) , .Z( u2_u15_X_12 ) );
  XOR2_X1 u2_u15_U47 (.A( u2_FP_40 ) , .B( u2_K16_11 ) , .Z( u2_u15_X_11 ) );
  XOR2_X1 u2_u15_U48 (.A( u2_FP_39 ) , .B( u2_K16_10 ) , .Z( u2_u15_X_10 ) );
  XOR2_X1 u2_u15_U5 (.A( u2_FP_36 ) , .B( u2_K16_5 ) , .Z( u2_u15_X_5 ) );
  XOR2_X1 u2_u15_U6 (.A( u2_FP_35 ) , .B( u2_K16_4 ) , .Z( u2_u15_X_4 ) );
  AND3_X1 u2_u15_u0_U10 (.A2( u2_u15_u0_n112 ) , .ZN( u2_u15_u0_n127 ) , .A3( u2_u15_u0_n130 ) , .A1( u2_u15_u0_n148 ) );
  NAND2_X1 u2_u15_u0_U11 (.ZN( u2_u15_u0_n113 ) , .A1( u2_u15_u0_n139 ) , .A2( u2_u15_u0_n149 ) );
  AND2_X1 u2_u15_u0_U12 (.ZN( u2_u15_u0_n107 ) , .A1( u2_u15_u0_n130 ) , .A2( u2_u15_u0_n140 ) );
  AND2_X1 u2_u15_u0_U13 (.A2( u2_u15_u0_n129 ) , .A1( u2_u15_u0_n130 ) , .ZN( u2_u15_u0_n151 ) );
  AND2_X1 u2_u15_u0_U14 (.A1( u2_u15_u0_n108 ) , .A2( u2_u15_u0_n125 ) , .ZN( u2_u15_u0_n145 ) );
  INV_X1 u2_u15_u0_U15 (.A( u2_u15_u0_n143 ) , .ZN( u2_u15_u0_n173 ) );
  NOR2_X1 u2_u15_u0_U16 (.A2( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n147 ) , .A1( u2_u15_u0_n160 ) );
  AOI21_X1 u2_u15_u0_U17 (.B1( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n132 ) , .A( u2_u15_u0_n165 ) , .B2( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U18 (.A( u2_u15_u0_n142 ) , .ZN( u2_u15_u0_n165 ) );
  OAI221_X1 u2_u15_u0_U19 (.C1( u2_u15_u0_n112 ) , .ZN( u2_u15_u0_n120 ) , .B1( u2_u15_u0_n138 ) , .B2( u2_u15_u0_n141 ) , .C2( u2_u15_u0_n147 ) , .A( u2_u15_u0_n172 ) );
  AOI211_X1 u2_u15_u0_U20 (.B( u2_u15_u0_n115 ) , .A( u2_u15_u0_n116 ) , .C2( u2_u15_u0_n117 ) , .C1( u2_u15_u0_n118 ) , .ZN( u2_u15_u0_n119 ) );
  OAI22_X1 u2_u15_u0_U21 (.B1( u2_u15_u0_n125 ) , .ZN( u2_u15_u0_n126 ) , .A1( u2_u15_u0_n138 ) , .A2( u2_u15_u0_n146 ) , .B2( u2_u15_u0_n147 ) );
  OAI22_X1 u2_u15_u0_U22 (.B1( u2_u15_u0_n131 ) , .A1( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n147 ) , .A2( u2_u15_u0_n90 ) , .ZN( u2_u15_u0_n91 ) );
  AND3_X1 u2_u15_u0_U23 (.A3( u2_u15_u0_n121 ) , .A2( u2_u15_u0_n125 ) , .A1( u2_u15_u0_n148 ) , .ZN( u2_u15_u0_n90 ) );
  INV_X1 u2_u15_u0_U24 (.A( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n161 ) );
  AOI22_X1 u2_u15_u0_U25 (.B2( u2_u15_u0_n109 ) , .A2( u2_u15_u0_n110 ) , .ZN( u2_u15_u0_n111 ) , .B1( u2_u15_u0_n118 ) , .A1( u2_u15_u0_n160 ) );
  INV_X1 u2_u15_u0_U26 (.A( u2_u15_u0_n118 ) , .ZN( u2_u15_u0_n158 ) );
  AOI21_X1 u2_u15_u0_U27 (.ZN( u2_u15_u0_n104 ) , .B1( u2_u15_u0_n107 ) , .B2( u2_u15_u0_n141 ) , .A( u2_u15_u0_n144 ) );
  AOI21_X1 u2_u15_u0_U28 (.B1( u2_u15_u0_n127 ) , .B2( u2_u15_u0_n129 ) , .A( u2_u15_u0_n138 ) , .ZN( u2_u15_u0_n96 ) );
  AOI21_X1 u2_u15_u0_U29 (.ZN( u2_u15_u0_n116 ) , .B2( u2_u15_u0_n142 ) , .A( u2_u15_u0_n144 ) , .B1( u2_u15_u0_n166 ) );
  INV_X1 u2_u15_u0_U3 (.A( u2_u15_u0_n113 ) , .ZN( u2_u15_u0_n166 ) );
  NAND2_X1 u2_u15_u0_U30 (.A1( u2_u15_u0_n100 ) , .A2( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n125 ) );
  NAND2_X1 u2_u15_u0_U31 (.A2( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n140 ) , .A1( u2_u15_u0_n94 ) );
  NAND2_X1 u2_u15_u0_U32 (.A1( u2_u15_u0_n101 ) , .A2( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n150 ) );
  INV_X1 u2_u15_u0_U33 (.A( u2_u15_u0_n138 ) , .ZN( u2_u15_u0_n160 ) );
  NAND2_X1 u2_u15_u0_U34 (.A2( u2_u15_u0_n102 ) , .A1( u2_u15_u0_n103 ) , .ZN( u2_u15_u0_n149 ) );
  NAND2_X1 u2_u15_u0_U35 (.A2( u2_u15_u0_n100 ) , .A1( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n139 ) );
  NAND2_X1 u2_u15_u0_U36 (.A2( u2_u15_u0_n100 ) , .ZN( u2_u15_u0_n131 ) , .A1( u2_u15_u0_n92 ) );
  NAND2_X1 u2_u15_u0_U37 (.ZN( u2_u15_u0_n108 ) , .A1( u2_u15_u0_n92 ) , .A2( u2_u15_u0_n94 ) );
  NAND2_X1 u2_u15_u0_U38 (.A2( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n114 ) , .A1( u2_u15_u0_n92 ) );
  NAND2_X1 u2_u15_u0_U39 (.A1( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n130 ) , .A2( u2_u15_u0_n94 ) );
  AOI21_X1 u2_u15_u0_U4 (.B1( u2_u15_u0_n114 ) , .ZN( u2_u15_u0_n115 ) , .B2( u2_u15_u0_n129 ) , .A( u2_u15_u0_n161 ) );
  NAND2_X1 u2_u15_u0_U40 (.A2( u2_u15_u0_n101 ) , .ZN( u2_u15_u0_n121 ) , .A1( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U41 (.ZN( u2_u15_u0_n172 ) , .A( u2_u15_u0_n88 ) );
  OAI222_X1 u2_u15_u0_U42 (.C1( u2_u15_u0_n108 ) , .A1( u2_u15_u0_n125 ) , .B2( u2_u15_u0_n128 ) , .B1( u2_u15_u0_n144 ) , .A2( u2_u15_u0_n158 ) , .C2( u2_u15_u0_n161 ) , .ZN( u2_u15_u0_n88 ) );
  NAND2_X1 u2_u15_u0_U43 (.ZN( u2_u15_u0_n112 ) , .A2( u2_u15_u0_n92 ) , .A1( u2_u15_u0_n93 ) );
  OR3_X1 u2_u15_u0_U44 (.A3( u2_u15_u0_n152 ) , .A2( u2_u15_u0_n153 ) , .A1( u2_u15_u0_n154 ) , .ZN( u2_u15_u0_n155 ) );
  AOI21_X1 u2_u15_u0_U45 (.B2( u2_u15_u0_n150 ) , .B1( u2_u15_u0_n151 ) , .ZN( u2_u15_u0_n152 ) , .A( u2_u15_u0_n158 ) );
  AOI21_X1 u2_u15_u0_U46 (.A( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n145 ) , .B1( u2_u15_u0_n146 ) , .ZN( u2_u15_u0_n154 ) );
  AOI21_X1 u2_u15_u0_U47 (.A( u2_u15_u0_n147 ) , .B2( u2_u15_u0_n148 ) , .B1( u2_u15_u0_n149 ) , .ZN( u2_u15_u0_n153 ) );
  INV_X1 u2_u15_u0_U48 (.ZN( u2_u15_u0_n171 ) , .A( u2_u15_u0_n99 ) );
  OAI211_X1 u2_u15_u0_U49 (.C2( u2_u15_u0_n140 ) , .C1( u2_u15_u0_n161 ) , .A( u2_u15_u0_n169 ) , .B( u2_u15_u0_n98 ) , .ZN( u2_u15_u0_n99 ) );
  AOI21_X1 u2_u15_u0_U5 (.B2( u2_u15_u0_n131 ) , .ZN( u2_u15_u0_n134 ) , .B1( u2_u15_u0_n151 ) , .A( u2_u15_u0_n158 ) );
  AOI211_X1 u2_u15_u0_U50 (.C1( u2_u15_u0_n118 ) , .A( u2_u15_u0_n123 ) , .B( u2_u15_u0_n96 ) , .C2( u2_u15_u0_n97 ) , .ZN( u2_u15_u0_n98 ) );
  INV_X1 u2_u15_u0_U51 (.ZN( u2_u15_u0_n169 ) , .A( u2_u15_u0_n91 ) );
  NOR2_X1 u2_u15_u0_U52 (.A2( u2_u15_X_2 ) , .ZN( u2_u15_u0_n103 ) , .A1( u2_u15_u0_n164 ) );
  NOR2_X1 u2_u15_u0_U53 (.A2( u2_u15_X_4 ) , .A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n118 ) );
  NOR2_X1 u2_u15_u0_U54 (.A2( u2_u15_X_1 ) , .A1( u2_u15_X_2 ) , .ZN( u2_u15_u0_n92 ) );
  NOR2_X1 u2_u15_u0_U55 (.A2( u2_u15_X_1 ) , .ZN( u2_u15_u0_n101 ) , .A1( u2_u15_u0_n163 ) );
  NOR2_X1 u2_u15_u0_U56 (.A2( u2_u15_X_3 ) , .A1( u2_u15_X_6 ) , .ZN( u2_u15_u0_n94 ) );
  NOR2_X1 u2_u15_u0_U57 (.A2( u2_u15_X_6 ) , .ZN( u2_u15_u0_n100 ) , .A1( u2_u15_u0_n162 ) );
  NAND2_X1 u2_u15_u0_U58 (.A2( u2_u15_X_4 ) , .A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n144 ) );
  NOR2_X1 u2_u15_u0_U59 (.A2( u2_u15_X_5 ) , .ZN( u2_u15_u0_n136 ) , .A1( u2_u15_u0_n159 ) );
  NOR2_X1 u2_u15_u0_U6 (.A1( u2_u15_u0_n108 ) , .ZN( u2_u15_u0_n123 ) , .A2( u2_u15_u0_n158 ) );
  NAND2_X1 u2_u15_u0_U60 (.A1( u2_u15_X_5 ) , .ZN( u2_u15_u0_n138 ) , .A2( u2_u15_u0_n159 ) );
  AND2_X1 u2_u15_u0_U61 (.A2( u2_u15_X_3 ) , .A1( u2_u15_X_6 ) , .ZN( u2_u15_u0_n102 ) );
  AND2_X1 u2_u15_u0_U62 (.A1( u2_u15_X_6 ) , .A2( u2_u15_u0_n162 ) , .ZN( u2_u15_u0_n93 ) );
  INV_X1 u2_u15_u0_U63 (.A( u2_u15_X_4 ) , .ZN( u2_u15_u0_n159 ) );
  INV_X1 u2_u15_u0_U64 (.A( u2_u15_X_1 ) , .ZN( u2_u15_u0_n164 ) );
  INV_X1 u2_u15_u0_U65 (.A( u2_u15_X_2 ) , .ZN( u2_u15_u0_n163 ) );
  INV_X1 u2_u15_u0_U66 (.A( u2_u15_X_3 ) , .ZN( u2_u15_u0_n162 ) );
  INV_X1 u2_u15_u0_U67 (.A( u2_u15_u0_n126 ) , .ZN( u2_u15_u0_n168 ) );
  AOI211_X1 u2_u15_u0_U68 (.B( u2_u15_u0_n133 ) , .A( u2_u15_u0_n134 ) , .C2( u2_u15_u0_n135 ) , .C1( u2_u15_u0_n136 ) , .ZN( u2_u15_u0_n137 ) );
  OR4_X1 u2_u15_u0_U69 (.ZN( u2_out15_17 ) , .A4( u2_u15_u0_n122 ) , .A2( u2_u15_u0_n123 ) , .A1( u2_u15_u0_n124 ) , .A3( u2_u15_u0_n170 ) );
  OAI21_X1 u2_u15_u0_U7 (.B1( u2_u15_u0_n150 ) , .B2( u2_u15_u0_n158 ) , .A( u2_u15_u0_n172 ) , .ZN( u2_u15_u0_n89 ) );
  AOI21_X1 u2_u15_u0_U70 (.B2( u2_u15_u0_n107 ) , .ZN( u2_u15_u0_n124 ) , .B1( u2_u15_u0_n128 ) , .A( u2_u15_u0_n161 ) );
  INV_X1 u2_u15_u0_U71 (.A( u2_u15_u0_n111 ) , .ZN( u2_u15_u0_n170 ) );
  OR4_X1 u2_u15_u0_U72 (.ZN( u2_out15_31 ) , .A4( u2_u15_u0_n155 ) , .A2( u2_u15_u0_n156 ) , .A1( u2_u15_u0_n157 ) , .A3( u2_u15_u0_n173 ) );
  AOI21_X1 u2_u15_u0_U73 (.A( u2_u15_u0_n138 ) , .B2( u2_u15_u0_n139 ) , .B1( u2_u15_u0_n140 ) , .ZN( u2_u15_u0_n157 ) );
  AOI21_X1 u2_u15_u0_U74 (.B2( u2_u15_u0_n141 ) , .B1( u2_u15_u0_n142 ) , .ZN( u2_u15_u0_n156 ) , .A( u2_u15_u0_n161 ) );
  INV_X1 u2_u15_u0_U75 (.ZN( u2_u15_u0_n174 ) , .A( u2_u15_u0_n89 ) );
  AOI211_X1 u2_u15_u0_U76 (.B( u2_u15_u0_n104 ) , .A( u2_u15_u0_n105 ) , .ZN( u2_u15_u0_n106 ) , .C2( u2_u15_u0_n113 ) , .C1( u2_u15_u0_n160 ) );
  NOR2_X1 u2_u15_u0_U77 (.A1( u2_u15_u0_n163 ) , .A2( u2_u15_u0_n164 ) , .ZN( u2_u15_u0_n95 ) );
  OAI221_X1 u2_u15_u0_U78 (.C1( u2_u15_u0_n121 ) , .ZN( u2_u15_u0_n122 ) , .B2( u2_u15_u0_n127 ) , .A( u2_u15_u0_n143 ) , .B1( u2_u15_u0_n144 ) , .C2( u2_u15_u0_n147 ) );
  NOR2_X1 u2_u15_u0_U79 (.A1( u2_u15_u0_n120 ) , .ZN( u2_u15_u0_n143 ) , .A2( u2_u15_u0_n167 ) );
  AND2_X1 u2_u15_u0_U8 (.A1( u2_u15_u0_n114 ) , .A2( u2_u15_u0_n121 ) , .ZN( u2_u15_u0_n146 ) );
  AOI21_X1 u2_u15_u0_U80 (.B1( u2_u15_u0_n132 ) , .ZN( u2_u15_u0_n133 ) , .A( u2_u15_u0_n144 ) , .B2( u2_u15_u0_n166 ) );
  OAI22_X1 u2_u15_u0_U81 (.ZN( u2_u15_u0_n105 ) , .A2( u2_u15_u0_n132 ) , .B1( u2_u15_u0_n146 ) , .A1( u2_u15_u0_n147 ) , .B2( u2_u15_u0_n161 ) );
  NAND2_X1 u2_u15_u0_U82 (.ZN( u2_u15_u0_n110 ) , .A2( u2_u15_u0_n132 ) , .A1( u2_u15_u0_n145 ) );
  INV_X1 u2_u15_u0_U83 (.A( u2_u15_u0_n119 ) , .ZN( u2_u15_u0_n167 ) );
  NAND2_X1 u2_u15_u0_U84 (.ZN( u2_u15_u0_n148 ) , .A1( u2_u15_u0_n93 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U85 (.A1( u2_u15_u0_n100 ) , .ZN( u2_u15_u0_n129 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U86 (.A1( u2_u15_u0_n102 ) , .ZN( u2_u15_u0_n128 ) , .A2( u2_u15_u0_n95 ) );
  NAND2_X1 u2_u15_u0_U87 (.ZN( u2_u15_u0_n142 ) , .A1( u2_u15_u0_n94 ) , .A2( u2_u15_u0_n95 ) );
  NAND3_X1 u2_u15_u0_U88 (.ZN( u2_out15_23 ) , .A3( u2_u15_u0_n137 ) , .A1( u2_u15_u0_n168 ) , .A2( u2_u15_u0_n171 ) );
  NAND3_X1 u2_u15_u0_U89 (.A3( u2_u15_u0_n127 ) , .A2( u2_u15_u0_n128 ) , .ZN( u2_u15_u0_n135 ) , .A1( u2_u15_u0_n150 ) );
  AND2_X1 u2_u15_u0_U9 (.A1( u2_u15_u0_n131 ) , .ZN( u2_u15_u0_n141 ) , .A2( u2_u15_u0_n150 ) );
  NAND3_X1 u2_u15_u0_U90 (.ZN( u2_u15_u0_n117 ) , .A3( u2_u15_u0_n132 ) , .A2( u2_u15_u0_n139 ) , .A1( u2_u15_u0_n148 ) );
  NAND3_X1 u2_u15_u0_U91 (.ZN( u2_u15_u0_n109 ) , .A2( u2_u15_u0_n114 ) , .A3( u2_u15_u0_n140 ) , .A1( u2_u15_u0_n149 ) );
  NAND3_X1 u2_u15_u0_U92 (.ZN( u2_out15_9 ) , .A3( u2_u15_u0_n106 ) , .A2( u2_u15_u0_n171 ) , .A1( u2_u15_u0_n174 ) );
  NAND3_X1 u2_u15_u0_U93 (.A2( u2_u15_u0_n128 ) , .A1( u2_u15_u0_n132 ) , .A3( u2_u15_u0_n146 ) , .ZN( u2_u15_u0_n97 ) );
  NOR2_X1 u2_u15_u1_U10 (.A1( u2_u15_u1_n112 ) , .A2( u2_u15_u1_n116 ) , .ZN( u2_u15_u1_n118 ) );
  NAND3_X1 u2_u15_u1_U100 (.ZN( u2_u15_u1_n113 ) , .A1( u2_u15_u1_n120 ) , .A3( u2_u15_u1_n133 ) , .A2( u2_u15_u1_n155 ) );
  OAI21_X1 u2_u15_u1_U11 (.ZN( u2_u15_u1_n101 ) , .B1( u2_u15_u1_n141 ) , .A( u2_u15_u1_n146 ) , .B2( u2_u15_u1_n183 ) );
  AOI21_X1 u2_u15_u1_U12 (.B2( u2_u15_u1_n155 ) , .B1( u2_u15_u1_n156 ) , .ZN( u2_u15_u1_n157 ) , .A( u2_u15_u1_n174 ) );
  NAND2_X1 u2_u15_u1_U13 (.ZN( u2_u15_u1_n140 ) , .A2( u2_u15_u1_n150 ) , .A1( u2_u15_u1_n155 ) );
  NAND2_X1 u2_u15_u1_U14 (.A1( u2_u15_u1_n131 ) , .ZN( u2_u15_u1_n147 ) , .A2( u2_u15_u1_n153 ) );
  INV_X1 u2_u15_u1_U15 (.A( u2_u15_u1_n139 ) , .ZN( u2_u15_u1_n174 ) );
  OR4_X1 u2_u15_u1_U16 (.A4( u2_u15_u1_n106 ) , .A3( u2_u15_u1_n107 ) , .ZN( u2_u15_u1_n108 ) , .A1( u2_u15_u1_n117 ) , .A2( u2_u15_u1_n184 ) );
  AOI21_X1 u2_u15_u1_U17 (.ZN( u2_u15_u1_n106 ) , .A( u2_u15_u1_n112 ) , .B1( u2_u15_u1_n154 ) , .B2( u2_u15_u1_n156 ) );
  AOI21_X1 u2_u15_u1_U18 (.ZN( u2_u15_u1_n107 ) , .B1( u2_u15_u1_n134 ) , .B2( u2_u15_u1_n149 ) , .A( u2_u15_u1_n174 ) );
  INV_X1 u2_u15_u1_U19 (.A( u2_u15_u1_n101 ) , .ZN( u2_u15_u1_n184 ) );
  INV_X1 u2_u15_u1_U20 (.A( u2_u15_u1_n112 ) , .ZN( u2_u15_u1_n171 ) );
  NAND2_X1 u2_u15_u1_U21 (.ZN( u2_u15_u1_n141 ) , .A1( u2_u15_u1_n153 ) , .A2( u2_u15_u1_n156 ) );
  AND2_X1 u2_u15_u1_U22 (.A1( u2_u15_u1_n123 ) , .ZN( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n161 ) );
  NAND2_X1 u2_u15_u1_U23 (.A2( u2_u15_u1_n115 ) , .A1( u2_u15_u1_n116 ) , .ZN( u2_u15_u1_n148 ) );
  NAND2_X1 u2_u15_u1_U24 (.A2( u2_u15_u1_n133 ) , .A1( u2_u15_u1_n135 ) , .ZN( u2_u15_u1_n159 ) );
  NAND2_X1 u2_u15_u1_U25 (.A2( u2_u15_u1_n115 ) , .A1( u2_u15_u1_n120 ) , .ZN( u2_u15_u1_n132 ) );
  INV_X1 u2_u15_u1_U26 (.A( u2_u15_u1_n154 ) , .ZN( u2_u15_u1_n178 ) );
  INV_X1 u2_u15_u1_U27 (.A( u2_u15_u1_n151 ) , .ZN( u2_u15_u1_n183 ) );
  AND2_X1 u2_u15_u1_U28 (.A1( u2_u15_u1_n129 ) , .A2( u2_u15_u1_n133 ) , .ZN( u2_u15_u1_n149 ) );
  INV_X1 u2_u15_u1_U29 (.A( u2_u15_u1_n131 ) , .ZN( u2_u15_u1_n180 ) );
  INV_X1 u2_u15_u1_U3 (.A( u2_u15_u1_n159 ) , .ZN( u2_u15_u1_n182 ) );
  OAI221_X1 u2_u15_u1_U30 (.A( u2_u15_u1_n119 ) , .C2( u2_u15_u1_n129 ) , .ZN( u2_u15_u1_n138 ) , .B2( u2_u15_u1_n152 ) , .C1( u2_u15_u1_n174 ) , .B1( u2_u15_u1_n187 ) );
  INV_X1 u2_u15_u1_U31 (.A( u2_u15_u1_n148 ) , .ZN( u2_u15_u1_n187 ) );
  AOI211_X1 u2_u15_u1_U32 (.B( u2_u15_u1_n117 ) , .A( u2_u15_u1_n118 ) , .ZN( u2_u15_u1_n119 ) , .C2( u2_u15_u1_n146 ) , .C1( u2_u15_u1_n159 ) );
  NOR2_X1 u2_u15_u1_U33 (.A1( u2_u15_u1_n168 ) , .A2( u2_u15_u1_n176 ) , .ZN( u2_u15_u1_n98 ) );
  AOI211_X1 u2_u15_u1_U34 (.B( u2_u15_u1_n162 ) , .A( u2_u15_u1_n163 ) , .C2( u2_u15_u1_n164 ) , .ZN( u2_u15_u1_n165 ) , .C1( u2_u15_u1_n171 ) );
  AOI21_X1 u2_u15_u1_U35 (.A( u2_u15_u1_n160 ) , .B2( u2_u15_u1_n161 ) , .ZN( u2_u15_u1_n162 ) , .B1( u2_u15_u1_n182 ) );
  OR2_X1 u2_u15_u1_U36 (.A2( u2_u15_u1_n157 ) , .A1( u2_u15_u1_n158 ) , .ZN( u2_u15_u1_n163 ) );
  NAND2_X1 u2_u15_u1_U37 (.A1( u2_u15_u1_n128 ) , .ZN( u2_u15_u1_n146 ) , .A2( u2_u15_u1_n160 ) );
  NAND2_X1 u2_u15_u1_U38 (.A2( u2_u15_u1_n112 ) , .ZN( u2_u15_u1_n139 ) , .A1( u2_u15_u1_n152 ) );
  NAND2_X1 u2_u15_u1_U39 (.A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n156 ) , .A2( u2_u15_u1_n99 ) );
  AOI221_X1 u2_u15_u1_U4 (.A( u2_u15_u1_n138 ) , .C2( u2_u15_u1_n139 ) , .C1( u2_u15_u1_n140 ) , .B2( u2_u15_u1_n141 ) , .ZN( u2_u15_u1_n142 ) , .B1( u2_u15_u1_n175 ) );
  AOI221_X1 u2_u15_u1_U40 (.B1( u2_u15_u1_n140 ) , .ZN( u2_u15_u1_n167 ) , .B2( u2_u15_u1_n172 ) , .C2( u2_u15_u1_n175 ) , .C1( u2_u15_u1_n178 ) , .A( u2_u15_u1_n188 ) );
  INV_X1 u2_u15_u1_U41 (.ZN( u2_u15_u1_n188 ) , .A( u2_u15_u1_n97 ) );
  AOI211_X1 u2_u15_u1_U42 (.A( u2_u15_u1_n118 ) , .C1( u2_u15_u1_n132 ) , .C2( u2_u15_u1_n139 ) , .B( u2_u15_u1_n96 ) , .ZN( u2_u15_u1_n97 ) );
  AOI21_X1 u2_u15_u1_U43 (.B2( u2_u15_u1_n121 ) , .B1( u2_u15_u1_n135 ) , .A( u2_u15_u1_n152 ) , .ZN( u2_u15_u1_n96 ) );
  NOR2_X1 u2_u15_u1_U44 (.ZN( u2_u15_u1_n117 ) , .A1( u2_u15_u1_n121 ) , .A2( u2_u15_u1_n160 ) );
  AOI21_X1 u2_u15_u1_U45 (.A( u2_u15_u1_n128 ) , .B2( u2_u15_u1_n129 ) , .ZN( u2_u15_u1_n130 ) , .B1( u2_u15_u1_n150 ) );
  OAI21_X1 u2_u15_u1_U46 (.B2( u2_u15_u1_n123 ) , .ZN( u2_u15_u1_n145 ) , .B1( u2_u15_u1_n160 ) , .A( u2_u15_u1_n185 ) );
  INV_X1 u2_u15_u1_U47 (.A( u2_u15_u1_n122 ) , .ZN( u2_u15_u1_n185 ) );
  AOI21_X1 u2_u15_u1_U48 (.B2( u2_u15_u1_n120 ) , .B1( u2_u15_u1_n121 ) , .ZN( u2_u15_u1_n122 ) , .A( u2_u15_u1_n128 ) );
  NAND2_X1 u2_u15_u1_U49 (.ZN( u2_u15_u1_n112 ) , .A1( u2_u15_u1_n169 ) , .A2( u2_u15_u1_n170 ) );
  AOI211_X1 u2_u15_u1_U5 (.ZN( u2_u15_u1_n124 ) , .A( u2_u15_u1_n138 ) , .C2( u2_u15_u1_n139 ) , .B( u2_u15_u1_n145 ) , .C1( u2_u15_u1_n147 ) );
  NAND2_X1 u2_u15_u1_U50 (.ZN( u2_u15_u1_n129 ) , .A2( u2_u15_u1_n95 ) , .A1( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U51 (.A1( u2_u15_u1_n102 ) , .ZN( u2_u15_u1_n154 ) , .A2( u2_u15_u1_n99 ) );
  NAND2_X1 u2_u15_u1_U52 (.A2( u2_u15_u1_n100 ) , .ZN( u2_u15_u1_n135 ) , .A1( u2_u15_u1_n99 ) );
  AOI21_X1 u2_u15_u1_U53 (.A( u2_u15_u1_n152 ) , .B2( u2_u15_u1_n153 ) , .B1( u2_u15_u1_n154 ) , .ZN( u2_u15_u1_n158 ) );
  INV_X1 u2_u15_u1_U54 (.A( u2_u15_u1_n160 ) , .ZN( u2_u15_u1_n175 ) );
  NAND2_X1 u2_u15_u1_U55 (.A1( u2_u15_u1_n100 ) , .ZN( u2_u15_u1_n116 ) , .A2( u2_u15_u1_n95 ) );
  NAND2_X1 u2_u15_u1_U56 (.A1( u2_u15_u1_n102 ) , .ZN( u2_u15_u1_n131 ) , .A2( u2_u15_u1_n95 ) );
  NAND2_X1 u2_u15_u1_U57 (.A2( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n121 ) , .A1( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U58 (.A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n153 ) , .A2( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U59 (.A2( u2_u15_u1_n104 ) , .A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n133 ) );
  AOI22_X1 u2_u15_u1_U6 (.B2( u2_u15_u1_n136 ) , .A2( u2_u15_u1_n137 ) , .ZN( u2_u15_u1_n143 ) , .A1( u2_u15_u1_n171 ) , .B1( u2_u15_u1_n173 ) );
  NAND2_X1 u2_u15_u1_U60 (.ZN( u2_u15_u1_n150 ) , .A2( u2_u15_u1_n98 ) , .A1( u2_u15_u1_n99 ) );
  NAND2_X1 u2_u15_u1_U61 (.A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n155 ) , .A2( u2_u15_u1_n95 ) );
  OAI21_X1 u2_u15_u1_U62 (.ZN( u2_u15_u1_n109 ) , .B1( u2_u15_u1_n129 ) , .B2( u2_u15_u1_n160 ) , .A( u2_u15_u1_n167 ) );
  NAND2_X1 u2_u15_u1_U63 (.A2( u2_u15_u1_n100 ) , .A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n120 ) );
  NAND2_X1 u2_u15_u1_U64 (.A1( u2_u15_u1_n102 ) , .A2( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n115 ) );
  NAND2_X1 u2_u15_u1_U65 (.A2( u2_u15_u1_n100 ) , .A1( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n151 ) );
  NAND2_X1 u2_u15_u1_U66 (.A2( u2_u15_u1_n103 ) , .A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n161 ) );
  INV_X1 u2_u15_u1_U67 (.A( u2_u15_u1_n152 ) , .ZN( u2_u15_u1_n173 ) );
  INV_X1 u2_u15_u1_U68 (.A( u2_u15_u1_n128 ) , .ZN( u2_u15_u1_n172 ) );
  NAND2_X1 u2_u15_u1_U69 (.A2( u2_u15_u1_n102 ) , .A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n123 ) );
  INV_X1 u2_u15_u1_U7 (.A( u2_u15_u1_n147 ) , .ZN( u2_u15_u1_n181 ) );
  NOR2_X1 u2_u15_u1_U70 (.A2( u2_u15_X_7 ) , .A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n95 ) );
  NOR2_X1 u2_u15_u1_U71 (.A1( u2_u15_X_12 ) , .A2( u2_u15_X_9 ) , .ZN( u2_u15_u1_n100 ) );
  NOR2_X1 u2_u15_u1_U72 (.A2( u2_u15_X_8 ) , .A1( u2_u15_u1_n177 ) , .ZN( u2_u15_u1_n99 ) );
  NOR2_X1 u2_u15_u1_U73 (.A2( u2_u15_X_12 ) , .ZN( u2_u15_u1_n102 ) , .A1( u2_u15_u1_n176 ) );
  NOR2_X1 u2_u15_u1_U74 (.A2( u2_u15_X_9 ) , .ZN( u2_u15_u1_n105 ) , .A1( u2_u15_u1_n168 ) );
  NAND2_X1 u2_u15_u1_U75 (.A1( u2_u15_X_10 ) , .ZN( u2_u15_u1_n160 ) , .A2( u2_u15_u1_n169 ) );
  NAND2_X1 u2_u15_u1_U76 (.A2( u2_u15_X_10 ) , .A1( u2_u15_X_11 ) , .ZN( u2_u15_u1_n152 ) );
  NAND2_X1 u2_u15_u1_U77 (.A1( u2_u15_X_11 ) , .ZN( u2_u15_u1_n128 ) , .A2( u2_u15_u1_n170 ) );
  AND2_X1 u2_u15_u1_U78 (.A2( u2_u15_X_7 ) , .A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n104 ) );
  AND2_X1 u2_u15_u1_U79 (.A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n103 ) , .A2( u2_u15_u1_n177 ) );
  AOI22_X1 u2_u15_u1_U8 (.B2( u2_u15_u1_n113 ) , .A2( u2_u15_u1_n114 ) , .ZN( u2_u15_u1_n125 ) , .A1( u2_u15_u1_n171 ) , .B1( u2_u15_u1_n173 ) );
  INV_X1 u2_u15_u1_U80 (.A( u2_u15_X_10 ) , .ZN( u2_u15_u1_n170 ) );
  INV_X1 u2_u15_u1_U81 (.A( u2_u15_X_9 ) , .ZN( u2_u15_u1_n176 ) );
  INV_X1 u2_u15_u1_U82 (.A( u2_u15_X_11 ) , .ZN( u2_u15_u1_n169 ) );
  INV_X1 u2_u15_u1_U83 (.A( u2_u15_X_12 ) , .ZN( u2_u15_u1_n168 ) );
  INV_X1 u2_u15_u1_U84 (.A( u2_u15_X_7 ) , .ZN( u2_u15_u1_n177 ) );
  NAND4_X1 u2_u15_u1_U85 (.ZN( u2_out15_18 ) , .A4( u2_u15_u1_n165 ) , .A3( u2_u15_u1_n166 ) , .A1( u2_u15_u1_n167 ) , .A2( u2_u15_u1_n186 ) );
  AOI22_X1 u2_u15_u1_U86 (.B2( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n147 ) , .A2( u2_u15_u1_n148 ) , .ZN( u2_u15_u1_n166 ) , .A1( u2_u15_u1_n172 ) );
  INV_X1 u2_u15_u1_U87 (.A( u2_u15_u1_n145 ) , .ZN( u2_u15_u1_n186 ) );
  NAND4_X1 u2_u15_u1_U88 (.ZN( u2_out15_2 ) , .A4( u2_u15_u1_n142 ) , .A3( u2_u15_u1_n143 ) , .A2( u2_u15_u1_n144 ) , .A1( u2_u15_u1_n179 ) );
  OAI21_X1 u2_u15_u1_U89 (.B2( u2_u15_u1_n132 ) , .ZN( u2_u15_u1_n144 ) , .A( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n180 ) );
  NAND2_X1 u2_u15_u1_U9 (.ZN( u2_u15_u1_n114 ) , .A1( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n156 ) );
  INV_X1 u2_u15_u1_U90 (.A( u2_u15_u1_n130 ) , .ZN( u2_u15_u1_n179 ) );
  NAND4_X1 u2_u15_u1_U91 (.ZN( u2_out15_28 ) , .A4( u2_u15_u1_n124 ) , .A3( u2_u15_u1_n125 ) , .A2( u2_u15_u1_n126 ) , .A1( u2_u15_u1_n127 ) );
  OAI21_X1 u2_u15_u1_U92 (.ZN( u2_u15_u1_n127 ) , .B2( u2_u15_u1_n139 ) , .B1( u2_u15_u1_n175 ) , .A( u2_u15_u1_n183 ) );
  OAI21_X1 u2_u15_u1_U93 (.ZN( u2_u15_u1_n126 ) , .B2( u2_u15_u1_n140 ) , .A( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n178 ) );
  OR4_X1 u2_u15_u1_U94 (.ZN( u2_out15_13 ) , .A4( u2_u15_u1_n108 ) , .A3( u2_u15_u1_n109 ) , .A2( u2_u15_u1_n110 ) , .A1( u2_u15_u1_n111 ) );
  AOI21_X1 u2_u15_u1_U95 (.ZN( u2_u15_u1_n111 ) , .A( u2_u15_u1_n128 ) , .B2( u2_u15_u1_n131 ) , .B1( u2_u15_u1_n135 ) );
  AOI21_X1 u2_u15_u1_U96 (.ZN( u2_u15_u1_n110 ) , .A( u2_u15_u1_n116 ) , .B1( u2_u15_u1_n152 ) , .B2( u2_u15_u1_n160 ) );
  NAND3_X1 u2_u15_u1_U97 (.A3( u2_u15_u1_n149 ) , .A2( u2_u15_u1_n150 ) , .A1( u2_u15_u1_n151 ) , .ZN( u2_u15_u1_n164 ) );
  NAND3_X1 u2_u15_u1_U98 (.A3( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n135 ) , .ZN( u2_u15_u1_n136 ) , .A1( u2_u15_u1_n151 ) );
  NAND3_X1 u2_u15_u1_U99 (.A1( u2_u15_u1_n133 ) , .ZN( u2_u15_u1_n137 ) , .A2( u2_u15_u1_n154 ) , .A3( u2_u15_u1_n181 ) );
  OAI22_X1 u2_u15_u2_U10 (.B1( u2_u15_u2_n151 ) , .A2( u2_u15_u2_n152 ) , .A1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n160 ) , .B2( u2_u15_u2_n168 ) );
  NAND3_X1 u2_u15_u2_U100 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n98 ) );
  NOR3_X1 u2_u15_u2_U11 (.A1( u2_u15_u2_n150 ) , .ZN( u2_u15_u2_n151 ) , .A3( u2_u15_u2_n175 ) , .A2( u2_u15_u2_n188 ) );
  AOI21_X1 u2_u15_u2_U12 (.B2( u2_u15_u2_n123 ) , .ZN( u2_u15_u2_n125 ) , .A( u2_u15_u2_n171 ) , .B1( u2_u15_u2_n184 ) );
  INV_X1 u2_u15_u2_U13 (.A( u2_u15_u2_n150 ) , .ZN( u2_u15_u2_n184 ) );
  AOI21_X1 u2_u15_u2_U14 (.ZN( u2_u15_u2_n144 ) , .B2( u2_u15_u2_n155 ) , .A( u2_u15_u2_n172 ) , .B1( u2_u15_u2_n185 ) );
  AOI21_X1 u2_u15_u2_U15 (.B2( u2_u15_u2_n143 ) , .ZN( u2_u15_u2_n145 ) , .B1( u2_u15_u2_n152 ) , .A( u2_u15_u2_n171 ) );
  INV_X1 u2_u15_u2_U16 (.A( u2_u15_u2_n156 ) , .ZN( u2_u15_u2_n171 ) );
  INV_X1 u2_u15_u2_U17 (.A( u2_u15_u2_n120 ) , .ZN( u2_u15_u2_n188 ) );
  NAND2_X1 u2_u15_u2_U18 (.A2( u2_u15_u2_n122 ) , .ZN( u2_u15_u2_n150 ) , .A1( u2_u15_u2_n152 ) );
  INV_X1 u2_u15_u2_U19 (.A( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n170 ) );
  INV_X1 u2_u15_u2_U20 (.A( u2_u15_u2_n137 ) , .ZN( u2_u15_u2_n173 ) );
  NAND2_X1 u2_u15_u2_U21 (.A1( u2_u15_u2_n132 ) , .A2( u2_u15_u2_n139 ) , .ZN( u2_u15_u2_n157 ) );
  INV_X1 u2_u15_u2_U22 (.A( u2_u15_u2_n113 ) , .ZN( u2_u15_u2_n178 ) );
  INV_X1 u2_u15_u2_U23 (.A( u2_u15_u2_n139 ) , .ZN( u2_u15_u2_n175 ) );
  INV_X1 u2_u15_u2_U24 (.A( u2_u15_u2_n155 ) , .ZN( u2_u15_u2_n181 ) );
  INV_X1 u2_u15_u2_U25 (.A( u2_u15_u2_n119 ) , .ZN( u2_u15_u2_n177 ) );
  INV_X1 u2_u15_u2_U26 (.A( u2_u15_u2_n116 ) , .ZN( u2_u15_u2_n180 ) );
  INV_X1 u2_u15_u2_U27 (.A( u2_u15_u2_n131 ) , .ZN( u2_u15_u2_n179 ) );
  INV_X1 u2_u15_u2_U28 (.A( u2_u15_u2_n154 ) , .ZN( u2_u15_u2_n176 ) );
  NAND2_X1 u2_u15_u2_U29 (.A2( u2_u15_u2_n116 ) , .A1( u2_u15_u2_n117 ) , .ZN( u2_u15_u2_n118 ) );
  NOR2_X1 u2_u15_u2_U3 (.ZN( u2_u15_u2_n121 ) , .A2( u2_u15_u2_n177 ) , .A1( u2_u15_u2_n180 ) );
  INV_X1 u2_u15_u2_U30 (.A( u2_u15_u2_n132 ) , .ZN( u2_u15_u2_n182 ) );
  INV_X1 u2_u15_u2_U31 (.A( u2_u15_u2_n158 ) , .ZN( u2_u15_u2_n183 ) );
  OAI21_X1 u2_u15_u2_U32 (.A( u2_u15_u2_n156 ) , .B1( u2_u15_u2_n157 ) , .ZN( u2_u15_u2_n158 ) , .B2( u2_u15_u2_n179 ) );
  NOR2_X1 u2_u15_u2_U33 (.ZN( u2_u15_u2_n156 ) , .A1( u2_u15_u2_n166 ) , .A2( u2_u15_u2_n169 ) );
  NOR2_X1 u2_u15_u2_U34 (.A2( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n137 ) , .A1( u2_u15_u2_n140 ) );
  NOR2_X1 u2_u15_u2_U35 (.A2( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n153 ) , .A1( u2_u15_u2_n156 ) );
  AOI211_X1 u2_u15_u2_U36 (.ZN( u2_u15_u2_n130 ) , .C1( u2_u15_u2_n138 ) , .C2( u2_u15_u2_n179 ) , .B( u2_u15_u2_n96 ) , .A( u2_u15_u2_n97 ) );
  OAI22_X1 u2_u15_u2_U37 (.B1( u2_u15_u2_n133 ) , .A2( u2_u15_u2_n137 ) , .A1( u2_u15_u2_n152 ) , .B2( u2_u15_u2_n168 ) , .ZN( u2_u15_u2_n97 ) );
  OAI221_X1 u2_u15_u2_U38 (.B1( u2_u15_u2_n113 ) , .C1( u2_u15_u2_n132 ) , .A( u2_u15_u2_n149 ) , .B2( u2_u15_u2_n171 ) , .C2( u2_u15_u2_n172 ) , .ZN( u2_u15_u2_n96 ) );
  OAI221_X1 u2_u15_u2_U39 (.A( u2_u15_u2_n115 ) , .C2( u2_u15_u2_n123 ) , .B2( u2_u15_u2_n143 ) , .B1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n163 ) , .C1( u2_u15_u2_n168 ) );
  INV_X1 u2_u15_u2_U4 (.A( u2_u15_u2_n134 ) , .ZN( u2_u15_u2_n185 ) );
  OAI21_X1 u2_u15_u2_U40 (.A( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n115 ) , .B1( u2_u15_u2_n176 ) , .B2( u2_u15_u2_n178 ) );
  OAI221_X1 u2_u15_u2_U41 (.A( u2_u15_u2_n135 ) , .B2( u2_u15_u2_n136 ) , .B1( u2_u15_u2_n137 ) , .ZN( u2_u15_u2_n162 ) , .C2( u2_u15_u2_n167 ) , .C1( u2_u15_u2_n185 ) );
  AND3_X1 u2_u15_u2_U42 (.A3( u2_u15_u2_n131 ) , .A2( u2_u15_u2_n132 ) , .A1( u2_u15_u2_n133 ) , .ZN( u2_u15_u2_n136 ) );
  AOI22_X1 u2_u15_u2_U43 (.ZN( u2_u15_u2_n135 ) , .B1( u2_u15_u2_n140 ) , .A1( u2_u15_u2_n156 ) , .B2( u2_u15_u2_n180 ) , .A2( u2_u15_u2_n188 ) );
  AOI21_X1 u2_u15_u2_U44 (.ZN( u2_u15_u2_n149 ) , .B1( u2_u15_u2_n173 ) , .B2( u2_u15_u2_n188 ) , .A( u2_u15_u2_n95 ) );
  AND3_X1 u2_u15_u2_U45 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n156 ) , .ZN( u2_u15_u2_n95 ) );
  OAI21_X1 u2_u15_u2_U46 (.A( u2_u15_u2_n141 ) , .B2( u2_u15_u2_n142 ) , .ZN( u2_u15_u2_n146 ) , .B1( u2_u15_u2_n153 ) );
  OAI21_X1 u2_u15_u2_U47 (.A( u2_u15_u2_n140 ) , .ZN( u2_u15_u2_n141 ) , .B1( u2_u15_u2_n176 ) , .B2( u2_u15_u2_n177 ) );
  NOR3_X1 u2_u15_u2_U48 (.ZN( u2_u15_u2_n142 ) , .A3( u2_u15_u2_n175 ) , .A2( u2_u15_u2_n178 ) , .A1( u2_u15_u2_n181 ) );
  OAI21_X1 u2_u15_u2_U49 (.A( u2_u15_u2_n101 ) , .B2( u2_u15_u2_n121 ) , .B1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n164 ) );
  NOR4_X1 u2_u15_u2_U5 (.A4( u2_u15_u2_n124 ) , .A3( u2_u15_u2_n125 ) , .A2( u2_u15_u2_n126 ) , .A1( u2_u15_u2_n127 ) , .ZN( u2_u15_u2_n128 ) );
  NAND2_X1 u2_u15_u2_U50 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n155 ) );
  NAND2_X1 u2_u15_u2_U51 (.A2( u2_u15_u2_n105 ) , .A1( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n143 ) );
  NAND2_X1 u2_u15_u2_U52 (.A1( u2_u15_u2_n104 ) , .A2( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n152 ) );
  NAND2_X1 u2_u15_u2_U53 (.A1( u2_u15_u2_n100 ) , .A2( u2_u15_u2_n105 ) , .ZN( u2_u15_u2_n132 ) );
  INV_X1 u2_u15_u2_U54 (.A( u2_u15_u2_n140 ) , .ZN( u2_u15_u2_n168 ) );
  INV_X1 u2_u15_u2_U55 (.A( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n167 ) );
  INV_X1 u2_u15_u2_U56 (.ZN( u2_u15_u2_n187 ) , .A( u2_u15_u2_n99 ) );
  OAI21_X1 u2_u15_u2_U57 (.B1( u2_u15_u2_n137 ) , .B2( u2_u15_u2_n143 ) , .A( u2_u15_u2_n98 ) , .ZN( u2_u15_u2_n99 ) );
  NAND2_X1 u2_u15_u2_U58 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n113 ) );
  NAND2_X1 u2_u15_u2_U59 (.A1( u2_u15_u2_n106 ) , .A2( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n131 ) );
  AOI21_X1 u2_u15_u2_U6 (.B2( u2_u15_u2_n119 ) , .ZN( u2_u15_u2_n127 ) , .A( u2_u15_u2_n137 ) , .B1( u2_u15_u2_n155 ) );
  NAND2_X1 u2_u15_u2_U60 (.A1( u2_u15_u2_n103 ) , .A2( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n139 ) );
  NAND2_X1 u2_u15_u2_U61 (.A1( u2_u15_u2_n103 ) , .A2( u2_u15_u2_n105 ) , .ZN( u2_u15_u2_n133 ) );
  NAND2_X1 u2_u15_u2_U62 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n103 ) , .ZN( u2_u15_u2_n154 ) );
  NAND2_X1 u2_u15_u2_U63 (.A2( u2_u15_u2_n103 ) , .A1( u2_u15_u2_n104 ) , .ZN( u2_u15_u2_n119 ) );
  NAND2_X1 u2_u15_u2_U64 (.A2( u2_u15_u2_n107 ) , .A1( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n123 ) );
  NAND2_X1 u2_u15_u2_U65 (.A1( u2_u15_u2_n104 ) , .A2( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n122 ) );
  INV_X1 u2_u15_u2_U66 (.A( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n172 ) );
  NAND2_X1 u2_u15_u2_U67 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n102 ) , .ZN( u2_u15_u2_n116 ) );
  NAND2_X1 u2_u15_u2_U68 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n120 ) );
  NAND2_X1 u2_u15_u2_U69 (.A2( u2_u15_u2_n105 ) , .A1( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n117 ) );
  AOI21_X1 u2_u15_u2_U7 (.ZN( u2_u15_u2_n124 ) , .B1( u2_u15_u2_n131 ) , .B2( u2_u15_u2_n143 ) , .A( u2_u15_u2_n172 ) );
  NOR2_X1 u2_u15_u2_U70 (.A2( u2_u15_X_16 ) , .ZN( u2_u15_u2_n140 ) , .A1( u2_u15_u2_n166 ) );
  NOR2_X1 u2_u15_u2_U71 (.A2( u2_u15_X_13 ) , .A1( u2_u15_X_14 ) , .ZN( u2_u15_u2_n100 ) );
  NOR2_X1 u2_u15_u2_U72 (.A2( u2_u15_X_16 ) , .A1( u2_u15_X_17 ) , .ZN( u2_u15_u2_n138 ) );
  NOR2_X1 u2_u15_u2_U73 (.A2( u2_u15_X_15 ) , .A1( u2_u15_X_18 ) , .ZN( u2_u15_u2_n104 ) );
  NOR2_X1 u2_u15_u2_U74 (.A2( u2_u15_X_14 ) , .ZN( u2_u15_u2_n103 ) , .A1( u2_u15_u2_n174 ) );
  NOR2_X1 u2_u15_u2_U75 (.A2( u2_u15_X_15 ) , .ZN( u2_u15_u2_n102 ) , .A1( u2_u15_u2_n165 ) );
  NOR2_X1 u2_u15_u2_U76 (.A2( u2_u15_X_17 ) , .ZN( u2_u15_u2_n114 ) , .A1( u2_u15_u2_n169 ) );
  AND2_X1 u2_u15_u2_U77 (.A1( u2_u15_X_15 ) , .ZN( u2_u15_u2_n105 ) , .A2( u2_u15_u2_n165 ) );
  AND2_X1 u2_u15_u2_U78 (.A2( u2_u15_X_15 ) , .A1( u2_u15_X_18 ) , .ZN( u2_u15_u2_n107 ) );
  AND2_X1 u2_u15_u2_U79 (.A1( u2_u15_X_14 ) , .ZN( u2_u15_u2_n106 ) , .A2( u2_u15_u2_n174 ) );
  AOI21_X1 u2_u15_u2_U8 (.B2( u2_u15_u2_n120 ) , .B1( u2_u15_u2_n121 ) , .ZN( u2_u15_u2_n126 ) , .A( u2_u15_u2_n167 ) );
  AND2_X1 u2_u15_u2_U80 (.A1( u2_u15_X_13 ) , .A2( u2_u15_X_14 ) , .ZN( u2_u15_u2_n108 ) );
  INV_X1 u2_u15_u2_U81 (.A( u2_u15_X_16 ) , .ZN( u2_u15_u2_n169 ) );
  INV_X1 u2_u15_u2_U82 (.A( u2_u15_X_17 ) , .ZN( u2_u15_u2_n166 ) );
  INV_X1 u2_u15_u2_U83 (.A( u2_u15_X_13 ) , .ZN( u2_u15_u2_n174 ) );
  INV_X1 u2_u15_u2_U84 (.A( u2_u15_X_18 ) , .ZN( u2_u15_u2_n165 ) );
  NAND4_X1 u2_u15_u2_U85 (.ZN( u2_out15_30 ) , .A4( u2_u15_u2_n147 ) , .A3( u2_u15_u2_n148 ) , .A2( u2_u15_u2_n149 ) , .A1( u2_u15_u2_n187 ) );
  NOR3_X1 u2_u15_u2_U86 (.A3( u2_u15_u2_n144 ) , .A2( u2_u15_u2_n145 ) , .A1( u2_u15_u2_n146 ) , .ZN( u2_u15_u2_n147 ) );
  AOI21_X1 u2_u15_u2_U87 (.B2( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n148 ) , .A( u2_u15_u2_n162 ) , .B1( u2_u15_u2_n182 ) );
  NAND4_X1 u2_u15_u2_U88 (.ZN( u2_out15_24 ) , .A4( u2_u15_u2_n111 ) , .A3( u2_u15_u2_n112 ) , .A1( u2_u15_u2_n130 ) , .A2( u2_u15_u2_n187 ) );
  AOI221_X1 u2_u15_u2_U89 (.A( u2_u15_u2_n109 ) , .B1( u2_u15_u2_n110 ) , .ZN( u2_u15_u2_n111 ) , .C1( u2_u15_u2_n134 ) , .C2( u2_u15_u2_n170 ) , .B2( u2_u15_u2_n173 ) );
  OAI22_X1 u2_u15_u2_U9 (.ZN( u2_u15_u2_n109 ) , .A2( u2_u15_u2_n113 ) , .B2( u2_u15_u2_n133 ) , .B1( u2_u15_u2_n167 ) , .A1( u2_u15_u2_n168 ) );
  AOI21_X1 u2_u15_u2_U90 (.ZN( u2_u15_u2_n112 ) , .B2( u2_u15_u2_n156 ) , .A( u2_u15_u2_n164 ) , .B1( u2_u15_u2_n181 ) );
  NAND4_X1 u2_u15_u2_U91 (.ZN( u2_out15_16 ) , .A4( u2_u15_u2_n128 ) , .A3( u2_u15_u2_n129 ) , .A1( u2_u15_u2_n130 ) , .A2( u2_u15_u2_n186 ) );
  AOI22_X1 u2_u15_u2_U92 (.A2( u2_u15_u2_n118 ) , .ZN( u2_u15_u2_n129 ) , .A1( u2_u15_u2_n140 ) , .B1( u2_u15_u2_n157 ) , .B2( u2_u15_u2_n170 ) );
  INV_X1 u2_u15_u2_U93 (.A( u2_u15_u2_n163 ) , .ZN( u2_u15_u2_n186 ) );
  OR4_X1 u2_u15_u2_U94 (.ZN( u2_out15_6 ) , .A4( u2_u15_u2_n161 ) , .A3( u2_u15_u2_n162 ) , .A2( u2_u15_u2_n163 ) , .A1( u2_u15_u2_n164 ) );
  OR3_X1 u2_u15_u2_U95 (.A2( u2_u15_u2_n159 ) , .A1( u2_u15_u2_n160 ) , .ZN( u2_u15_u2_n161 ) , .A3( u2_u15_u2_n183 ) );
  AOI21_X1 u2_u15_u2_U96 (.B2( u2_u15_u2_n154 ) , .B1( u2_u15_u2_n155 ) , .ZN( u2_u15_u2_n159 ) , .A( u2_u15_u2_n167 ) );
  NAND3_X1 u2_u15_u2_U97 (.A2( u2_u15_u2_n117 ) , .A1( u2_u15_u2_n122 ) , .A3( u2_u15_u2_n123 ) , .ZN( u2_u15_u2_n134 ) );
  NAND3_X1 u2_u15_u2_U98 (.ZN( u2_u15_u2_n110 ) , .A2( u2_u15_u2_n131 ) , .A3( u2_u15_u2_n139 ) , .A1( u2_u15_u2_n154 ) );
  NAND3_X1 u2_u15_u2_U99 (.A2( u2_u15_u2_n100 ) , .ZN( u2_u15_u2_n101 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n114 ) );
  OAI22_X1 u2_u15_u3_U10 (.B1( u2_u15_u3_n113 ) , .A2( u2_u15_u3_n135 ) , .A1( u2_u15_u3_n150 ) , .B2( u2_u15_u3_n164 ) , .ZN( u2_u15_u3_n98 ) );
  OAI211_X1 u2_u15_u3_U11 (.B( u2_u15_u3_n106 ) , .ZN( u2_u15_u3_n119 ) , .C2( u2_u15_u3_n128 ) , .C1( u2_u15_u3_n167 ) , .A( u2_u15_u3_n181 ) );
  AOI221_X1 u2_u15_u3_U12 (.C1( u2_u15_u3_n105 ) , .ZN( u2_u15_u3_n106 ) , .A( u2_u15_u3_n131 ) , .B2( u2_u15_u3_n132 ) , .C2( u2_u15_u3_n133 ) , .B1( u2_u15_u3_n169 ) );
  INV_X1 u2_u15_u3_U13 (.ZN( u2_u15_u3_n181 ) , .A( u2_u15_u3_n98 ) );
  NAND2_X1 u2_u15_u3_U14 (.ZN( u2_u15_u3_n105 ) , .A2( u2_u15_u3_n130 ) , .A1( u2_u15_u3_n155 ) );
  AOI22_X1 u2_u15_u3_U15 (.B1( u2_u15_u3_n115 ) , .A2( u2_u15_u3_n116 ) , .ZN( u2_u15_u3_n123 ) , .B2( u2_u15_u3_n133 ) , .A1( u2_u15_u3_n169 ) );
  NAND2_X1 u2_u15_u3_U16 (.ZN( u2_u15_u3_n116 ) , .A2( u2_u15_u3_n151 ) , .A1( u2_u15_u3_n182 ) );
  NOR2_X1 u2_u15_u3_U17 (.ZN( u2_u15_u3_n126 ) , .A2( u2_u15_u3_n150 ) , .A1( u2_u15_u3_n164 ) );
  AOI21_X1 u2_u15_u3_U18 (.ZN( u2_u15_u3_n112 ) , .B2( u2_u15_u3_n146 ) , .B1( u2_u15_u3_n155 ) , .A( u2_u15_u3_n167 ) );
  NAND2_X1 u2_u15_u3_U19 (.A1( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n142 ) , .A2( u2_u15_u3_n164 ) );
  NAND2_X1 u2_u15_u3_U20 (.ZN( u2_u15_u3_n132 ) , .A2( u2_u15_u3_n152 ) , .A1( u2_u15_u3_n156 ) );
  AND2_X1 u2_u15_u3_U21 (.A2( u2_u15_u3_n113 ) , .A1( u2_u15_u3_n114 ) , .ZN( u2_u15_u3_n151 ) );
  INV_X1 u2_u15_u3_U22 (.A( u2_u15_u3_n133 ) , .ZN( u2_u15_u3_n165 ) );
  INV_X1 u2_u15_u3_U23 (.A( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n170 ) );
  NAND2_X1 u2_u15_u3_U24 (.A1( u2_u15_u3_n107 ) , .A2( u2_u15_u3_n108 ) , .ZN( u2_u15_u3_n140 ) );
  NAND2_X1 u2_u15_u3_U25 (.ZN( u2_u15_u3_n117 ) , .A1( u2_u15_u3_n124 ) , .A2( u2_u15_u3_n148 ) );
  NAND2_X1 u2_u15_u3_U26 (.ZN( u2_u15_u3_n143 ) , .A1( u2_u15_u3_n165 ) , .A2( u2_u15_u3_n167 ) );
  INV_X1 u2_u15_u3_U27 (.A( u2_u15_u3_n130 ) , .ZN( u2_u15_u3_n177 ) );
  INV_X1 u2_u15_u3_U28 (.A( u2_u15_u3_n128 ) , .ZN( u2_u15_u3_n176 ) );
  INV_X1 u2_u15_u3_U29 (.A( u2_u15_u3_n155 ) , .ZN( u2_u15_u3_n174 ) );
  INV_X1 u2_u15_u3_U3 (.A( u2_u15_u3_n129 ) , .ZN( u2_u15_u3_n183 ) );
  INV_X1 u2_u15_u3_U30 (.A( u2_u15_u3_n139 ) , .ZN( u2_u15_u3_n185 ) );
  NOR2_X1 u2_u15_u3_U31 (.ZN( u2_u15_u3_n135 ) , .A2( u2_u15_u3_n141 ) , .A1( u2_u15_u3_n169 ) );
  OAI222_X1 u2_u15_u3_U32 (.C2( u2_u15_u3_n107 ) , .A2( u2_u15_u3_n108 ) , .B1( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n138 ) , .B2( u2_u15_u3_n146 ) , .C1( u2_u15_u3_n154 ) , .A1( u2_u15_u3_n164 ) );
  NOR4_X1 u2_u15_u3_U33 (.A4( u2_u15_u3_n157 ) , .A3( u2_u15_u3_n158 ) , .A2( u2_u15_u3_n159 ) , .A1( u2_u15_u3_n160 ) , .ZN( u2_u15_u3_n161 ) );
  AOI21_X1 u2_u15_u3_U34 (.B2( u2_u15_u3_n152 ) , .B1( u2_u15_u3_n153 ) , .ZN( u2_u15_u3_n158 ) , .A( u2_u15_u3_n164 ) );
  AOI21_X1 u2_u15_u3_U35 (.A( u2_u15_u3_n154 ) , .B2( u2_u15_u3_n155 ) , .B1( u2_u15_u3_n156 ) , .ZN( u2_u15_u3_n157 ) );
  AOI21_X1 u2_u15_u3_U36 (.A( u2_u15_u3_n149 ) , .B2( u2_u15_u3_n150 ) , .B1( u2_u15_u3_n151 ) , .ZN( u2_u15_u3_n159 ) );
  AOI211_X1 u2_u15_u3_U37 (.ZN( u2_u15_u3_n109 ) , .A( u2_u15_u3_n119 ) , .C2( u2_u15_u3_n129 ) , .B( u2_u15_u3_n138 ) , .C1( u2_u15_u3_n141 ) );
  AOI211_X1 u2_u15_u3_U38 (.B( u2_u15_u3_n119 ) , .A( u2_u15_u3_n120 ) , .C2( u2_u15_u3_n121 ) , .ZN( u2_u15_u3_n122 ) , .C1( u2_u15_u3_n179 ) );
  INV_X1 u2_u15_u3_U39 (.A( u2_u15_u3_n156 ) , .ZN( u2_u15_u3_n179 ) );
  INV_X1 u2_u15_u3_U4 (.A( u2_u15_u3_n140 ) , .ZN( u2_u15_u3_n182 ) );
  OAI22_X1 u2_u15_u3_U40 (.B1( u2_u15_u3_n118 ) , .ZN( u2_u15_u3_n120 ) , .A1( u2_u15_u3_n135 ) , .B2( u2_u15_u3_n154 ) , .A2( u2_u15_u3_n178 ) );
  AND3_X1 u2_u15_u3_U41 (.ZN( u2_u15_u3_n118 ) , .A2( u2_u15_u3_n124 ) , .A1( u2_u15_u3_n144 ) , .A3( u2_u15_u3_n152 ) );
  INV_X1 u2_u15_u3_U42 (.A( u2_u15_u3_n121 ) , .ZN( u2_u15_u3_n164 ) );
  NAND2_X1 u2_u15_u3_U43 (.ZN( u2_u15_u3_n133 ) , .A1( u2_u15_u3_n154 ) , .A2( u2_u15_u3_n164 ) );
  OAI211_X1 u2_u15_u3_U44 (.B( u2_u15_u3_n127 ) , .ZN( u2_u15_u3_n139 ) , .C1( u2_u15_u3_n150 ) , .C2( u2_u15_u3_n154 ) , .A( u2_u15_u3_n184 ) );
  INV_X1 u2_u15_u3_U45 (.A( u2_u15_u3_n125 ) , .ZN( u2_u15_u3_n184 ) );
  AOI221_X1 u2_u15_u3_U46 (.A( u2_u15_u3_n126 ) , .ZN( u2_u15_u3_n127 ) , .C2( u2_u15_u3_n132 ) , .C1( u2_u15_u3_n169 ) , .B2( u2_u15_u3_n170 ) , .B1( u2_u15_u3_n174 ) );
  OAI22_X1 u2_u15_u3_U47 (.A1( u2_u15_u3_n124 ) , .ZN( u2_u15_u3_n125 ) , .B2( u2_u15_u3_n145 ) , .A2( u2_u15_u3_n165 ) , .B1( u2_u15_u3_n167 ) );
  NOR2_X1 u2_u15_u3_U48 (.A1( u2_u15_u3_n113 ) , .ZN( u2_u15_u3_n131 ) , .A2( u2_u15_u3_n154 ) );
  NAND2_X1 u2_u15_u3_U49 (.A1( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n150 ) , .A2( u2_u15_u3_n99 ) );
  INV_X1 u2_u15_u3_U5 (.A( u2_u15_u3_n117 ) , .ZN( u2_u15_u3_n178 ) );
  NAND2_X1 u2_u15_u3_U50 (.A2( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n155 ) , .A1( u2_u15_u3_n97 ) );
  INV_X1 u2_u15_u3_U51 (.A( u2_u15_u3_n141 ) , .ZN( u2_u15_u3_n167 ) );
  AOI21_X1 u2_u15_u3_U52 (.B2( u2_u15_u3_n114 ) , .B1( u2_u15_u3_n146 ) , .A( u2_u15_u3_n154 ) , .ZN( u2_u15_u3_n94 ) );
  AOI21_X1 u2_u15_u3_U53 (.ZN( u2_u15_u3_n110 ) , .B2( u2_u15_u3_n142 ) , .B1( u2_u15_u3_n186 ) , .A( u2_u15_u3_n95 ) );
  INV_X1 u2_u15_u3_U54 (.A( u2_u15_u3_n145 ) , .ZN( u2_u15_u3_n186 ) );
  AOI21_X1 u2_u15_u3_U55 (.B1( u2_u15_u3_n124 ) , .A( u2_u15_u3_n149 ) , .B2( u2_u15_u3_n155 ) , .ZN( u2_u15_u3_n95 ) );
  INV_X1 u2_u15_u3_U56 (.A( u2_u15_u3_n149 ) , .ZN( u2_u15_u3_n169 ) );
  NAND2_X1 u2_u15_u3_U57 (.ZN( u2_u15_u3_n124 ) , .A1( u2_u15_u3_n96 ) , .A2( u2_u15_u3_n97 ) );
  NAND2_X1 u2_u15_u3_U58 (.A2( u2_u15_u3_n100 ) , .ZN( u2_u15_u3_n146 ) , .A1( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U59 (.A1( u2_u15_u3_n101 ) , .ZN( u2_u15_u3_n145 ) , .A2( u2_u15_u3_n99 ) );
  AOI221_X1 u2_u15_u3_U6 (.A( u2_u15_u3_n131 ) , .C2( u2_u15_u3_n132 ) , .C1( u2_u15_u3_n133 ) , .ZN( u2_u15_u3_n134 ) , .B1( u2_u15_u3_n143 ) , .B2( u2_u15_u3_n177 ) );
  NAND2_X1 u2_u15_u3_U60 (.A1( u2_u15_u3_n100 ) , .ZN( u2_u15_u3_n156 ) , .A2( u2_u15_u3_n99 ) );
  NAND2_X1 u2_u15_u3_U61 (.A2( u2_u15_u3_n101 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n148 ) );
  NAND2_X1 u2_u15_u3_U62 (.A1( u2_u15_u3_n100 ) , .A2( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n128 ) );
  NAND2_X1 u2_u15_u3_U63 (.A2( u2_u15_u3_n101 ) , .A1( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n152 ) );
  NAND2_X1 u2_u15_u3_U64 (.A2( u2_u15_u3_n101 ) , .ZN( u2_u15_u3_n114 ) , .A1( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U65 (.ZN( u2_u15_u3_n107 ) , .A1( u2_u15_u3_n97 ) , .A2( u2_u15_u3_n99 ) );
  NAND2_X1 u2_u15_u3_U66 (.A2( u2_u15_u3_n100 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n113 ) );
  NAND2_X1 u2_u15_u3_U67 (.A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n153 ) , .A2( u2_u15_u3_n97 ) );
  NAND2_X1 u2_u15_u3_U68 (.A2( u2_u15_u3_n103 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n130 ) );
  NAND2_X1 u2_u15_u3_U69 (.A2( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n144 ) , .A1( u2_u15_u3_n96 ) );
  OAI22_X1 u2_u15_u3_U7 (.B2( u2_u15_u3_n147 ) , .A2( u2_u15_u3_n148 ) , .ZN( u2_u15_u3_n160 ) , .B1( u2_u15_u3_n165 ) , .A1( u2_u15_u3_n168 ) );
  NAND2_X1 u2_u15_u3_U70 (.A1( u2_u15_u3_n102 ) , .A2( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n108 ) );
  NOR2_X1 u2_u15_u3_U71 (.A2( u2_u15_X_19 ) , .A1( u2_u15_X_20 ) , .ZN( u2_u15_u3_n99 ) );
  NOR2_X1 u2_u15_u3_U72 (.A2( u2_u15_X_21 ) , .A1( u2_u15_X_24 ) , .ZN( u2_u15_u3_n103 ) );
  NOR2_X1 u2_u15_u3_U73 (.A2( u2_u15_X_24 ) , .A1( u2_u15_u3_n171 ) , .ZN( u2_u15_u3_n97 ) );
  NOR2_X1 u2_u15_u3_U74 (.A2( u2_u15_X_23 ) , .ZN( u2_u15_u3_n141 ) , .A1( u2_u15_u3_n166 ) );
  NOR2_X1 u2_u15_u3_U75 (.A2( u2_u15_X_19 ) , .A1( u2_u15_u3_n172 ) , .ZN( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U76 (.A1( u2_u15_X_22 ) , .A2( u2_u15_X_23 ) , .ZN( u2_u15_u3_n154 ) );
  NAND2_X1 u2_u15_u3_U77 (.A1( u2_u15_X_23 ) , .ZN( u2_u15_u3_n149 ) , .A2( u2_u15_u3_n166 ) );
  NOR2_X1 u2_u15_u3_U78 (.A2( u2_u15_X_22 ) , .A1( u2_u15_X_23 ) , .ZN( u2_u15_u3_n121 ) );
  AND2_X1 u2_u15_u3_U79 (.A1( u2_u15_X_24 ) , .ZN( u2_u15_u3_n101 ) , .A2( u2_u15_u3_n171 ) );
  AND3_X1 u2_u15_u3_U8 (.A3( u2_u15_u3_n144 ) , .A2( u2_u15_u3_n145 ) , .A1( u2_u15_u3_n146 ) , .ZN( u2_u15_u3_n147 ) );
  AND2_X1 u2_u15_u3_U80 (.A1( u2_u15_X_19 ) , .ZN( u2_u15_u3_n102 ) , .A2( u2_u15_u3_n172 ) );
  AND2_X1 u2_u15_u3_U81 (.A1( u2_u15_X_21 ) , .A2( u2_u15_X_24 ) , .ZN( u2_u15_u3_n100 ) );
  AND2_X1 u2_u15_u3_U82 (.A2( u2_u15_X_19 ) , .A1( u2_u15_X_20 ) , .ZN( u2_u15_u3_n104 ) );
  INV_X1 u2_u15_u3_U83 (.A( u2_u15_X_22 ) , .ZN( u2_u15_u3_n166 ) );
  INV_X1 u2_u15_u3_U84 (.A( u2_u15_X_21 ) , .ZN( u2_u15_u3_n171 ) );
  INV_X1 u2_u15_u3_U85 (.A( u2_u15_X_20 ) , .ZN( u2_u15_u3_n172 ) );
  OR4_X1 u2_u15_u3_U86 (.ZN( u2_out15_10 ) , .A4( u2_u15_u3_n136 ) , .A3( u2_u15_u3_n137 ) , .A1( u2_u15_u3_n138 ) , .A2( u2_u15_u3_n139 ) );
  OAI222_X1 u2_u15_u3_U87 (.C1( u2_u15_u3_n128 ) , .ZN( u2_u15_u3_n137 ) , .B1( u2_u15_u3_n148 ) , .A2( u2_u15_u3_n150 ) , .B2( u2_u15_u3_n154 ) , .C2( u2_u15_u3_n164 ) , .A1( u2_u15_u3_n167 ) );
  OAI221_X1 u2_u15_u3_U88 (.A( u2_u15_u3_n134 ) , .B2( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n136 ) , .C1( u2_u15_u3_n149 ) , .B1( u2_u15_u3_n151 ) , .C2( u2_u15_u3_n183 ) );
  NAND4_X1 u2_u15_u3_U89 (.ZN( u2_out15_1 ) , .A4( u2_u15_u3_n161 ) , .A3( u2_u15_u3_n162 ) , .A2( u2_u15_u3_n163 ) , .A1( u2_u15_u3_n185 ) );
  INV_X1 u2_u15_u3_U9 (.A( u2_u15_u3_n143 ) , .ZN( u2_u15_u3_n168 ) );
  NAND2_X1 u2_u15_u3_U90 (.ZN( u2_u15_u3_n163 ) , .A2( u2_u15_u3_n170 ) , .A1( u2_u15_u3_n176 ) );
  AOI22_X1 u2_u15_u3_U91 (.B2( u2_u15_u3_n140 ) , .B1( u2_u15_u3_n141 ) , .A2( u2_u15_u3_n142 ) , .ZN( u2_u15_u3_n162 ) , .A1( u2_u15_u3_n177 ) );
  NAND4_X1 u2_u15_u3_U92 (.ZN( u2_out15_26 ) , .A4( u2_u15_u3_n109 ) , .A3( u2_u15_u3_n110 ) , .A2( u2_u15_u3_n111 ) , .A1( u2_u15_u3_n173 ) );
  INV_X1 u2_u15_u3_U93 (.ZN( u2_u15_u3_n173 ) , .A( u2_u15_u3_n94 ) );
  OAI21_X1 u2_u15_u3_U94 (.ZN( u2_u15_u3_n111 ) , .B2( u2_u15_u3_n117 ) , .A( u2_u15_u3_n133 ) , .B1( u2_u15_u3_n176 ) );
  NAND4_X1 u2_u15_u3_U95 (.ZN( u2_out15_20 ) , .A4( u2_u15_u3_n122 ) , .A3( u2_u15_u3_n123 ) , .A1( u2_u15_u3_n175 ) , .A2( u2_u15_u3_n180 ) );
  INV_X1 u2_u15_u3_U96 (.A( u2_u15_u3_n126 ) , .ZN( u2_u15_u3_n180 ) );
  INV_X1 u2_u15_u3_U97 (.A( u2_u15_u3_n112 ) , .ZN( u2_u15_u3_n175 ) );
  NAND3_X1 u2_u15_u3_U98 (.A1( u2_u15_u3_n114 ) , .ZN( u2_u15_u3_n115 ) , .A2( u2_u15_u3_n145 ) , .A3( u2_u15_u3_n153 ) );
  NAND3_X1 u2_u15_u3_U99 (.ZN( u2_u15_u3_n129 ) , .A2( u2_u15_u3_n144 ) , .A1( u2_u15_u3_n153 ) , .A3( u2_u15_u3_n182 ) );
  XOR2_X1 u2_u1_U1 (.B( u2_K2_9 ) , .A( u2_R0_6 ) , .Z( u2_u1_X_9 ) );
  XOR2_X1 u2_u1_U16 (.B( u2_K2_3 ) , .A( u2_R0_2 ) , .Z( u2_u1_X_3 ) );
  XOR2_X1 u2_u1_U2 (.B( u2_K2_8 ) , .A( u2_R0_5 ) , .Z( u2_u1_X_8 ) );
  XOR2_X1 u2_u1_U27 (.B( u2_K2_2 ) , .A( u2_R0_1 ) , .Z( u2_u1_X_2 ) );
  XOR2_X1 u2_u1_U3 (.B( u2_K2_7 ) , .A( u2_R0_4 ) , .Z( u2_u1_X_7 ) );
  XOR2_X1 u2_u1_U38 (.B( u2_K2_1 ) , .A( u2_R0_32 ) , .Z( u2_u1_X_1 ) );
  XOR2_X1 u2_u1_U4 (.B( u2_K2_6 ) , .A( u2_R0_5 ) , .Z( u2_u1_X_6 ) );
  XOR2_X1 u2_u1_U46 (.B( u2_K2_12 ) , .A( u2_R0_9 ) , .Z( u2_u1_X_12 ) );
  XOR2_X1 u2_u1_U47 (.B( u2_K2_11 ) , .A( u2_R0_8 ) , .Z( u2_u1_X_11 ) );
  XOR2_X1 u2_u1_U48 (.B( u2_K2_10 ) , .A( u2_R0_7 ) , .Z( u2_u1_X_10 ) );
  XOR2_X1 u2_u1_U5 (.B( u2_K2_5 ) , .A( u2_R0_4 ) , .Z( u2_u1_X_5 ) );
  XOR2_X1 u2_u1_U6 (.B( u2_K2_4 ) , .A( u2_R0_3 ) , .Z( u2_u1_X_4 ) );
  AND3_X1 u2_u1_u0_U10 (.A2( u2_u1_u0_n112 ) , .ZN( u2_u1_u0_n127 ) , .A3( u2_u1_u0_n130 ) , .A1( u2_u1_u0_n148 ) );
  NAND2_X1 u2_u1_u0_U11 (.ZN( u2_u1_u0_n113 ) , .A1( u2_u1_u0_n139 ) , .A2( u2_u1_u0_n149 ) );
  AND2_X1 u2_u1_u0_U12 (.ZN( u2_u1_u0_n107 ) , .A1( u2_u1_u0_n130 ) , .A2( u2_u1_u0_n140 ) );
  AND2_X1 u2_u1_u0_U13 (.A2( u2_u1_u0_n129 ) , .A1( u2_u1_u0_n130 ) , .ZN( u2_u1_u0_n151 ) );
  AND2_X1 u2_u1_u0_U14 (.A1( u2_u1_u0_n108 ) , .A2( u2_u1_u0_n125 ) , .ZN( u2_u1_u0_n145 ) );
  INV_X1 u2_u1_u0_U15 (.A( u2_u1_u0_n143 ) , .ZN( u2_u1_u0_n173 ) );
  NOR2_X1 u2_u1_u0_U16 (.A2( u2_u1_u0_n136 ) , .ZN( u2_u1_u0_n147 ) , .A1( u2_u1_u0_n160 ) );
  NOR2_X1 u2_u1_u0_U17 (.A1( u2_u1_u0_n163 ) , .A2( u2_u1_u0_n164 ) , .ZN( u2_u1_u0_n95 ) );
  AOI21_X1 u2_u1_u0_U18 (.B1( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n132 ) , .A( u2_u1_u0_n165 ) , .B2( u2_u1_u0_n93 ) );
  INV_X1 u2_u1_u0_U19 (.A( u2_u1_u0_n142 ) , .ZN( u2_u1_u0_n165 ) );
  OAI221_X1 u2_u1_u0_U20 (.C1( u2_u1_u0_n121 ) , .ZN( u2_u1_u0_n122 ) , .B2( u2_u1_u0_n127 ) , .A( u2_u1_u0_n143 ) , .B1( u2_u1_u0_n144 ) , .C2( u2_u1_u0_n147 ) );
  OAI22_X1 u2_u1_u0_U21 (.B1( u2_u1_u0_n125 ) , .ZN( u2_u1_u0_n126 ) , .A1( u2_u1_u0_n138 ) , .A2( u2_u1_u0_n146 ) , .B2( u2_u1_u0_n147 ) );
  OAI22_X1 u2_u1_u0_U22 (.B1( u2_u1_u0_n131 ) , .A1( u2_u1_u0_n144 ) , .B2( u2_u1_u0_n147 ) , .A2( u2_u1_u0_n90 ) , .ZN( u2_u1_u0_n91 ) );
  AND3_X1 u2_u1_u0_U23 (.A3( u2_u1_u0_n121 ) , .A2( u2_u1_u0_n125 ) , .A1( u2_u1_u0_n148 ) , .ZN( u2_u1_u0_n90 ) );
  NAND2_X1 u2_u1_u0_U24 (.A1( u2_u1_u0_n100 ) , .A2( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n125 ) );
  INV_X1 u2_u1_u0_U25 (.A( u2_u1_u0_n136 ) , .ZN( u2_u1_u0_n161 ) );
  NOR2_X1 u2_u1_u0_U26 (.A1( u2_u1_u0_n120 ) , .ZN( u2_u1_u0_n143 ) , .A2( u2_u1_u0_n167 ) );
  OAI221_X1 u2_u1_u0_U27 (.C1( u2_u1_u0_n112 ) , .ZN( u2_u1_u0_n120 ) , .B1( u2_u1_u0_n138 ) , .B2( u2_u1_u0_n141 ) , .C2( u2_u1_u0_n147 ) , .A( u2_u1_u0_n172 ) );
  AOI211_X1 u2_u1_u0_U28 (.B( u2_u1_u0_n115 ) , .A( u2_u1_u0_n116 ) , .C2( u2_u1_u0_n117 ) , .C1( u2_u1_u0_n118 ) , .ZN( u2_u1_u0_n119 ) );
  AOI22_X1 u2_u1_u0_U29 (.B2( u2_u1_u0_n109 ) , .A2( u2_u1_u0_n110 ) , .ZN( u2_u1_u0_n111 ) , .B1( u2_u1_u0_n118 ) , .A1( u2_u1_u0_n160 ) );
  INV_X1 u2_u1_u0_U3 (.A( u2_u1_u0_n113 ) , .ZN( u2_u1_u0_n166 ) );
  NAND2_X1 u2_u1_u0_U30 (.A1( u2_u1_u0_n100 ) , .ZN( u2_u1_u0_n129 ) , .A2( u2_u1_u0_n95 ) );
  INV_X1 u2_u1_u0_U31 (.A( u2_u1_u0_n118 ) , .ZN( u2_u1_u0_n158 ) );
  AOI21_X1 u2_u1_u0_U32 (.ZN( u2_u1_u0_n104 ) , .B1( u2_u1_u0_n107 ) , .B2( u2_u1_u0_n141 ) , .A( u2_u1_u0_n144 ) );
  AOI21_X1 u2_u1_u0_U33 (.B1( u2_u1_u0_n127 ) , .B2( u2_u1_u0_n129 ) , .A( u2_u1_u0_n138 ) , .ZN( u2_u1_u0_n96 ) );
  AOI21_X1 u2_u1_u0_U34 (.ZN( u2_u1_u0_n116 ) , .B2( u2_u1_u0_n142 ) , .A( u2_u1_u0_n144 ) , .B1( u2_u1_u0_n166 ) );
  NAND2_X1 u2_u1_u0_U35 (.A2( u2_u1_u0_n100 ) , .A1( u2_u1_u0_n101 ) , .ZN( u2_u1_u0_n139 ) );
  NAND2_X1 u2_u1_u0_U36 (.A2( u2_u1_u0_n100 ) , .ZN( u2_u1_u0_n131 ) , .A1( u2_u1_u0_n92 ) );
  NAND2_X1 u2_u1_u0_U37 (.A1( u2_u1_u0_n101 ) , .A2( u2_u1_u0_n102 ) , .ZN( u2_u1_u0_n150 ) );
  INV_X1 u2_u1_u0_U38 (.A( u2_u1_u0_n138 ) , .ZN( u2_u1_u0_n160 ) );
  NAND2_X1 u2_u1_u0_U39 (.A1( u2_u1_u0_n102 ) , .ZN( u2_u1_u0_n128 ) , .A2( u2_u1_u0_n95 ) );
  AOI21_X1 u2_u1_u0_U4 (.B1( u2_u1_u0_n114 ) , .ZN( u2_u1_u0_n115 ) , .B2( u2_u1_u0_n129 ) , .A( u2_u1_u0_n161 ) );
  NAND2_X1 u2_u1_u0_U40 (.ZN( u2_u1_u0_n148 ) , .A1( u2_u1_u0_n93 ) , .A2( u2_u1_u0_n95 ) );
  NAND2_X1 u2_u1_u0_U41 (.A2( u2_u1_u0_n102 ) , .A1( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n149 ) );
  NAND2_X1 u2_u1_u0_U42 (.A2( u2_u1_u0_n102 ) , .ZN( u2_u1_u0_n114 ) , .A1( u2_u1_u0_n92 ) );
  NAND2_X1 u2_u1_u0_U43 (.A2( u2_u1_u0_n101 ) , .ZN( u2_u1_u0_n121 ) , .A1( u2_u1_u0_n93 ) );
  INV_X1 u2_u1_u0_U44 (.ZN( u2_u1_u0_n172 ) , .A( u2_u1_u0_n88 ) );
  OAI222_X1 u2_u1_u0_U45 (.C1( u2_u1_u0_n108 ) , .A1( u2_u1_u0_n125 ) , .B2( u2_u1_u0_n128 ) , .B1( u2_u1_u0_n144 ) , .A2( u2_u1_u0_n158 ) , .C2( u2_u1_u0_n161 ) , .ZN( u2_u1_u0_n88 ) );
  NAND2_X1 u2_u1_u0_U46 (.ZN( u2_u1_u0_n112 ) , .A2( u2_u1_u0_n92 ) , .A1( u2_u1_u0_n93 ) );
  OR3_X1 u2_u1_u0_U47 (.A3( u2_u1_u0_n152 ) , .A2( u2_u1_u0_n153 ) , .A1( u2_u1_u0_n154 ) , .ZN( u2_u1_u0_n155 ) );
  AOI21_X1 u2_u1_u0_U48 (.B2( u2_u1_u0_n150 ) , .B1( u2_u1_u0_n151 ) , .ZN( u2_u1_u0_n152 ) , .A( u2_u1_u0_n158 ) );
  AOI21_X1 u2_u1_u0_U49 (.A( u2_u1_u0_n144 ) , .B2( u2_u1_u0_n145 ) , .B1( u2_u1_u0_n146 ) , .ZN( u2_u1_u0_n154 ) );
  AOI21_X1 u2_u1_u0_U5 (.B2( u2_u1_u0_n131 ) , .ZN( u2_u1_u0_n134 ) , .B1( u2_u1_u0_n151 ) , .A( u2_u1_u0_n158 ) );
  AOI21_X1 u2_u1_u0_U50 (.A( u2_u1_u0_n147 ) , .B2( u2_u1_u0_n148 ) , .B1( u2_u1_u0_n149 ) , .ZN( u2_u1_u0_n153 ) );
  INV_X1 u2_u1_u0_U51 (.ZN( u2_u1_u0_n171 ) , .A( u2_u1_u0_n99 ) );
  OAI211_X1 u2_u1_u0_U52 (.C2( u2_u1_u0_n140 ) , .C1( u2_u1_u0_n161 ) , .A( u2_u1_u0_n169 ) , .B( u2_u1_u0_n98 ) , .ZN( u2_u1_u0_n99 ) );
  AOI211_X1 u2_u1_u0_U53 (.C1( u2_u1_u0_n118 ) , .A( u2_u1_u0_n123 ) , .B( u2_u1_u0_n96 ) , .C2( u2_u1_u0_n97 ) , .ZN( u2_u1_u0_n98 ) );
  INV_X1 u2_u1_u0_U54 (.ZN( u2_u1_u0_n169 ) , .A( u2_u1_u0_n91 ) );
  NOR2_X1 u2_u1_u0_U55 (.A2( u2_u1_X_4 ) , .A1( u2_u1_X_5 ) , .ZN( u2_u1_u0_n118 ) );
  NOR2_X1 u2_u1_u0_U56 (.A2( u2_u1_X_2 ) , .ZN( u2_u1_u0_n103 ) , .A1( u2_u1_u0_n164 ) );
  NOR2_X1 u2_u1_u0_U57 (.A2( u2_u1_X_1 ) , .A1( u2_u1_X_2 ) , .ZN( u2_u1_u0_n92 ) );
  NOR2_X1 u2_u1_u0_U58 (.A2( u2_u1_X_1 ) , .ZN( u2_u1_u0_n101 ) , .A1( u2_u1_u0_n163 ) );
  NAND2_X1 u2_u1_u0_U59 (.A2( u2_u1_X_4 ) , .A1( u2_u1_X_5 ) , .ZN( u2_u1_u0_n144 ) );
  NOR2_X1 u2_u1_u0_U6 (.A1( u2_u1_u0_n108 ) , .ZN( u2_u1_u0_n123 ) , .A2( u2_u1_u0_n158 ) );
  NOR2_X1 u2_u1_u0_U60 (.A2( u2_u1_X_5 ) , .ZN( u2_u1_u0_n136 ) , .A1( u2_u1_u0_n159 ) );
  NAND2_X1 u2_u1_u0_U61 (.A1( u2_u1_X_5 ) , .ZN( u2_u1_u0_n138 ) , .A2( u2_u1_u0_n159 ) );
  AND2_X1 u2_u1_u0_U62 (.A2( u2_u1_X_3 ) , .A1( u2_u1_X_6 ) , .ZN( u2_u1_u0_n102 ) );
  AND2_X1 u2_u1_u0_U63 (.A1( u2_u1_X_6 ) , .A2( u2_u1_u0_n162 ) , .ZN( u2_u1_u0_n93 ) );
  INV_X1 u2_u1_u0_U64 (.A( u2_u1_X_4 ) , .ZN( u2_u1_u0_n159 ) );
  INV_X1 u2_u1_u0_U65 (.A( u2_u1_X_1 ) , .ZN( u2_u1_u0_n164 ) );
  INV_X1 u2_u1_u0_U66 (.A( u2_u1_X_2 ) , .ZN( u2_u1_u0_n163 ) );
  INV_X1 u2_u1_u0_U67 (.A( u2_u1_X_3 ) , .ZN( u2_u1_u0_n162 ) );
  INV_X1 u2_u1_u0_U68 (.A( u2_u1_u0_n126 ) , .ZN( u2_u1_u0_n168 ) );
  AOI211_X1 u2_u1_u0_U69 (.B( u2_u1_u0_n133 ) , .A( u2_u1_u0_n134 ) , .C2( u2_u1_u0_n135 ) , .C1( u2_u1_u0_n136 ) , .ZN( u2_u1_u0_n137 ) );
  OAI21_X1 u2_u1_u0_U7 (.B1( u2_u1_u0_n150 ) , .B2( u2_u1_u0_n158 ) , .A( u2_u1_u0_n172 ) , .ZN( u2_u1_u0_n89 ) );
  INV_X1 u2_u1_u0_U70 (.ZN( u2_u1_u0_n174 ) , .A( u2_u1_u0_n89 ) );
  AOI211_X1 u2_u1_u0_U71 (.B( u2_u1_u0_n104 ) , .A( u2_u1_u0_n105 ) , .ZN( u2_u1_u0_n106 ) , .C2( u2_u1_u0_n113 ) , .C1( u2_u1_u0_n160 ) );
  OR4_X1 u2_u1_u0_U72 (.ZN( u2_out1_17 ) , .A4( u2_u1_u0_n122 ) , .A2( u2_u1_u0_n123 ) , .A1( u2_u1_u0_n124 ) , .A3( u2_u1_u0_n170 ) );
  AOI21_X1 u2_u1_u0_U73 (.B2( u2_u1_u0_n107 ) , .ZN( u2_u1_u0_n124 ) , .B1( u2_u1_u0_n128 ) , .A( u2_u1_u0_n161 ) );
  INV_X1 u2_u1_u0_U74 (.A( u2_u1_u0_n111 ) , .ZN( u2_u1_u0_n170 ) );
  OR4_X1 u2_u1_u0_U75 (.ZN( u2_out1_31 ) , .A4( u2_u1_u0_n155 ) , .A2( u2_u1_u0_n156 ) , .A1( u2_u1_u0_n157 ) , .A3( u2_u1_u0_n173 ) );
  AOI21_X1 u2_u1_u0_U76 (.A( u2_u1_u0_n138 ) , .B2( u2_u1_u0_n139 ) , .B1( u2_u1_u0_n140 ) , .ZN( u2_u1_u0_n157 ) );
  AOI21_X1 u2_u1_u0_U77 (.B2( u2_u1_u0_n141 ) , .B1( u2_u1_u0_n142 ) , .ZN( u2_u1_u0_n156 ) , .A( u2_u1_u0_n161 ) );
  AOI21_X1 u2_u1_u0_U78 (.B1( u2_u1_u0_n132 ) , .ZN( u2_u1_u0_n133 ) , .A( u2_u1_u0_n144 ) , .B2( u2_u1_u0_n166 ) );
  OAI22_X1 u2_u1_u0_U79 (.ZN( u2_u1_u0_n105 ) , .A2( u2_u1_u0_n132 ) , .B1( u2_u1_u0_n146 ) , .A1( u2_u1_u0_n147 ) , .B2( u2_u1_u0_n161 ) );
  AND2_X1 u2_u1_u0_U8 (.A1( u2_u1_u0_n114 ) , .A2( u2_u1_u0_n121 ) , .ZN( u2_u1_u0_n146 ) );
  NAND2_X1 u2_u1_u0_U80 (.ZN( u2_u1_u0_n110 ) , .A2( u2_u1_u0_n132 ) , .A1( u2_u1_u0_n145 ) );
  INV_X1 u2_u1_u0_U81 (.A( u2_u1_u0_n119 ) , .ZN( u2_u1_u0_n167 ) );
  NAND2_X1 u2_u1_u0_U82 (.A2( u2_u1_u0_n103 ) , .ZN( u2_u1_u0_n140 ) , .A1( u2_u1_u0_n94 ) );
  NAND2_X1 u2_u1_u0_U83 (.A1( u2_u1_u0_n101 ) , .ZN( u2_u1_u0_n130 ) , .A2( u2_u1_u0_n94 ) );
  NAND2_X1 u2_u1_u0_U84 (.ZN( u2_u1_u0_n108 ) , .A1( u2_u1_u0_n92 ) , .A2( u2_u1_u0_n94 ) );
  NAND2_X1 u2_u1_u0_U85 (.ZN( u2_u1_u0_n142 ) , .A1( u2_u1_u0_n94 ) , .A2( u2_u1_u0_n95 ) );
  NOR2_X1 u2_u1_u0_U86 (.A2( u2_u1_X_6 ) , .ZN( u2_u1_u0_n100 ) , .A1( u2_u1_u0_n162 ) );
  NOR2_X1 u2_u1_u0_U87 (.A2( u2_u1_X_3 ) , .A1( u2_u1_X_6 ) , .ZN( u2_u1_u0_n94 ) );
  NAND3_X1 u2_u1_u0_U88 (.ZN( u2_out1_23 ) , .A3( u2_u1_u0_n137 ) , .A1( u2_u1_u0_n168 ) , .A2( u2_u1_u0_n171 ) );
  NAND3_X1 u2_u1_u0_U89 (.A3( u2_u1_u0_n127 ) , .A2( u2_u1_u0_n128 ) , .ZN( u2_u1_u0_n135 ) , .A1( u2_u1_u0_n150 ) );
  AND2_X1 u2_u1_u0_U9 (.A1( u2_u1_u0_n131 ) , .ZN( u2_u1_u0_n141 ) , .A2( u2_u1_u0_n150 ) );
  NAND3_X1 u2_u1_u0_U90 (.ZN( u2_u1_u0_n117 ) , .A3( u2_u1_u0_n132 ) , .A2( u2_u1_u0_n139 ) , .A1( u2_u1_u0_n148 ) );
  NAND3_X1 u2_u1_u0_U91 (.ZN( u2_u1_u0_n109 ) , .A2( u2_u1_u0_n114 ) , .A3( u2_u1_u0_n140 ) , .A1( u2_u1_u0_n149 ) );
  NAND3_X1 u2_u1_u0_U92 (.ZN( u2_out1_9 ) , .A3( u2_u1_u0_n106 ) , .A2( u2_u1_u0_n171 ) , .A1( u2_u1_u0_n174 ) );
  NAND3_X1 u2_u1_u0_U93 (.A2( u2_u1_u0_n128 ) , .A1( u2_u1_u0_n132 ) , .A3( u2_u1_u0_n146 ) , .ZN( u2_u1_u0_n97 ) );
  NOR2_X1 u2_u1_u1_U10 (.A1( u2_u1_u1_n112 ) , .A2( u2_u1_u1_n116 ) , .ZN( u2_u1_u1_n118 ) );
  NAND3_X1 u2_u1_u1_U100 (.ZN( u2_u1_u1_n113 ) , .A1( u2_u1_u1_n120 ) , .A3( u2_u1_u1_n133 ) , .A2( u2_u1_u1_n155 ) );
  OAI21_X1 u2_u1_u1_U11 (.ZN( u2_u1_u1_n101 ) , .B1( u2_u1_u1_n141 ) , .A( u2_u1_u1_n146 ) , .B2( u2_u1_u1_n183 ) );
  AOI21_X1 u2_u1_u1_U12 (.B2( u2_u1_u1_n155 ) , .B1( u2_u1_u1_n156 ) , .ZN( u2_u1_u1_n157 ) , .A( u2_u1_u1_n174 ) );
  OR4_X1 u2_u1_u1_U13 (.A4( u2_u1_u1_n106 ) , .A3( u2_u1_u1_n107 ) , .ZN( u2_u1_u1_n108 ) , .A1( u2_u1_u1_n117 ) , .A2( u2_u1_u1_n184 ) );
  AOI21_X1 u2_u1_u1_U14 (.ZN( u2_u1_u1_n106 ) , .A( u2_u1_u1_n112 ) , .B1( u2_u1_u1_n154 ) , .B2( u2_u1_u1_n156 ) );
  INV_X1 u2_u1_u1_U15 (.A( u2_u1_u1_n101 ) , .ZN( u2_u1_u1_n184 ) );
  AOI21_X1 u2_u1_u1_U16 (.ZN( u2_u1_u1_n107 ) , .B1( u2_u1_u1_n134 ) , .B2( u2_u1_u1_n149 ) , .A( u2_u1_u1_n174 ) );
  NAND2_X1 u2_u1_u1_U17 (.ZN( u2_u1_u1_n140 ) , .A2( u2_u1_u1_n150 ) , .A1( u2_u1_u1_n155 ) );
  NAND2_X1 u2_u1_u1_U18 (.A1( u2_u1_u1_n131 ) , .ZN( u2_u1_u1_n147 ) , .A2( u2_u1_u1_n153 ) );
  INV_X1 u2_u1_u1_U19 (.A( u2_u1_u1_n139 ) , .ZN( u2_u1_u1_n174 ) );
  INV_X1 u2_u1_u1_U20 (.A( u2_u1_u1_n112 ) , .ZN( u2_u1_u1_n171 ) );
  NAND2_X1 u2_u1_u1_U21 (.ZN( u2_u1_u1_n141 ) , .A1( u2_u1_u1_n153 ) , .A2( u2_u1_u1_n156 ) );
  AND2_X1 u2_u1_u1_U22 (.A1( u2_u1_u1_n123 ) , .ZN( u2_u1_u1_n134 ) , .A2( u2_u1_u1_n161 ) );
  NAND2_X1 u2_u1_u1_U23 (.A2( u2_u1_u1_n115 ) , .A1( u2_u1_u1_n116 ) , .ZN( u2_u1_u1_n148 ) );
  NAND2_X1 u2_u1_u1_U24 (.A2( u2_u1_u1_n133 ) , .A1( u2_u1_u1_n135 ) , .ZN( u2_u1_u1_n159 ) );
  NAND2_X1 u2_u1_u1_U25 (.A2( u2_u1_u1_n115 ) , .A1( u2_u1_u1_n120 ) , .ZN( u2_u1_u1_n132 ) );
  INV_X1 u2_u1_u1_U26 (.A( u2_u1_u1_n154 ) , .ZN( u2_u1_u1_n178 ) );
  INV_X1 u2_u1_u1_U27 (.A( u2_u1_u1_n151 ) , .ZN( u2_u1_u1_n183 ) );
  AND2_X1 u2_u1_u1_U28 (.A1( u2_u1_u1_n129 ) , .A2( u2_u1_u1_n133 ) , .ZN( u2_u1_u1_n149 ) );
  INV_X1 u2_u1_u1_U29 (.A( u2_u1_u1_n131 ) , .ZN( u2_u1_u1_n180 ) );
  INV_X1 u2_u1_u1_U3 (.A( u2_u1_u1_n159 ) , .ZN( u2_u1_u1_n182 ) );
  AOI221_X1 u2_u1_u1_U30 (.B1( u2_u1_u1_n140 ) , .ZN( u2_u1_u1_n167 ) , .B2( u2_u1_u1_n172 ) , .C2( u2_u1_u1_n175 ) , .C1( u2_u1_u1_n178 ) , .A( u2_u1_u1_n188 ) );
  INV_X1 u2_u1_u1_U31 (.ZN( u2_u1_u1_n188 ) , .A( u2_u1_u1_n97 ) );
  AOI211_X1 u2_u1_u1_U32 (.A( u2_u1_u1_n118 ) , .C1( u2_u1_u1_n132 ) , .C2( u2_u1_u1_n139 ) , .B( u2_u1_u1_n96 ) , .ZN( u2_u1_u1_n97 ) );
  AOI21_X1 u2_u1_u1_U33 (.B2( u2_u1_u1_n121 ) , .B1( u2_u1_u1_n135 ) , .A( u2_u1_u1_n152 ) , .ZN( u2_u1_u1_n96 ) );
  OAI221_X1 u2_u1_u1_U34 (.A( u2_u1_u1_n119 ) , .C2( u2_u1_u1_n129 ) , .ZN( u2_u1_u1_n138 ) , .B2( u2_u1_u1_n152 ) , .C1( u2_u1_u1_n174 ) , .B1( u2_u1_u1_n187 ) );
  INV_X1 u2_u1_u1_U35 (.A( u2_u1_u1_n148 ) , .ZN( u2_u1_u1_n187 ) );
  AOI211_X1 u2_u1_u1_U36 (.B( u2_u1_u1_n117 ) , .A( u2_u1_u1_n118 ) , .ZN( u2_u1_u1_n119 ) , .C2( u2_u1_u1_n146 ) , .C1( u2_u1_u1_n159 ) );
  NOR2_X1 u2_u1_u1_U37 (.A1( u2_u1_u1_n168 ) , .A2( u2_u1_u1_n176 ) , .ZN( u2_u1_u1_n98 ) );
  AOI211_X1 u2_u1_u1_U38 (.B( u2_u1_u1_n162 ) , .A( u2_u1_u1_n163 ) , .C2( u2_u1_u1_n164 ) , .ZN( u2_u1_u1_n165 ) , .C1( u2_u1_u1_n171 ) );
  AOI21_X1 u2_u1_u1_U39 (.A( u2_u1_u1_n160 ) , .B2( u2_u1_u1_n161 ) , .ZN( u2_u1_u1_n162 ) , .B1( u2_u1_u1_n182 ) );
  AOI221_X1 u2_u1_u1_U4 (.A( u2_u1_u1_n138 ) , .C2( u2_u1_u1_n139 ) , .C1( u2_u1_u1_n140 ) , .B2( u2_u1_u1_n141 ) , .ZN( u2_u1_u1_n142 ) , .B1( u2_u1_u1_n175 ) );
  OR2_X1 u2_u1_u1_U40 (.A2( u2_u1_u1_n157 ) , .A1( u2_u1_u1_n158 ) , .ZN( u2_u1_u1_n163 ) );
  OAI21_X1 u2_u1_u1_U41 (.B2( u2_u1_u1_n123 ) , .ZN( u2_u1_u1_n145 ) , .B1( u2_u1_u1_n160 ) , .A( u2_u1_u1_n185 ) );
  INV_X1 u2_u1_u1_U42 (.A( u2_u1_u1_n122 ) , .ZN( u2_u1_u1_n185 ) );
  AOI21_X1 u2_u1_u1_U43 (.B2( u2_u1_u1_n120 ) , .B1( u2_u1_u1_n121 ) , .ZN( u2_u1_u1_n122 ) , .A( u2_u1_u1_n128 ) );
  NAND2_X1 u2_u1_u1_U44 (.A1( u2_u1_u1_n128 ) , .ZN( u2_u1_u1_n146 ) , .A2( u2_u1_u1_n160 ) );
  NAND2_X1 u2_u1_u1_U45 (.A2( u2_u1_u1_n112 ) , .ZN( u2_u1_u1_n139 ) , .A1( u2_u1_u1_n152 ) );
  NAND2_X1 u2_u1_u1_U46 (.A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n156 ) , .A2( u2_u1_u1_n99 ) );
  NOR2_X1 u2_u1_u1_U47 (.ZN( u2_u1_u1_n117 ) , .A1( u2_u1_u1_n121 ) , .A2( u2_u1_u1_n160 ) );
  AOI21_X1 u2_u1_u1_U48 (.A( u2_u1_u1_n128 ) , .B2( u2_u1_u1_n129 ) , .ZN( u2_u1_u1_n130 ) , .B1( u2_u1_u1_n150 ) );
  NAND2_X1 u2_u1_u1_U49 (.ZN( u2_u1_u1_n112 ) , .A1( u2_u1_u1_n169 ) , .A2( u2_u1_u1_n170 ) );
  AOI211_X1 u2_u1_u1_U5 (.ZN( u2_u1_u1_n124 ) , .A( u2_u1_u1_n138 ) , .C2( u2_u1_u1_n139 ) , .B( u2_u1_u1_n145 ) , .C1( u2_u1_u1_n147 ) );
  NAND2_X1 u2_u1_u1_U50 (.ZN( u2_u1_u1_n129 ) , .A2( u2_u1_u1_n95 ) , .A1( u2_u1_u1_n98 ) );
  NAND2_X1 u2_u1_u1_U51 (.A1( u2_u1_u1_n102 ) , .ZN( u2_u1_u1_n154 ) , .A2( u2_u1_u1_n99 ) );
  NAND2_X1 u2_u1_u1_U52 (.A2( u2_u1_u1_n100 ) , .ZN( u2_u1_u1_n135 ) , .A1( u2_u1_u1_n99 ) );
  AOI21_X1 u2_u1_u1_U53 (.A( u2_u1_u1_n152 ) , .B2( u2_u1_u1_n153 ) , .B1( u2_u1_u1_n154 ) , .ZN( u2_u1_u1_n158 ) );
  INV_X1 u2_u1_u1_U54 (.A( u2_u1_u1_n160 ) , .ZN( u2_u1_u1_n175 ) );
  NAND2_X1 u2_u1_u1_U55 (.A1( u2_u1_u1_n100 ) , .ZN( u2_u1_u1_n116 ) , .A2( u2_u1_u1_n95 ) );
  NAND2_X1 u2_u1_u1_U56 (.A1( u2_u1_u1_n102 ) , .ZN( u2_u1_u1_n131 ) , .A2( u2_u1_u1_n95 ) );
  NAND2_X1 u2_u1_u1_U57 (.A2( u2_u1_u1_n104 ) , .ZN( u2_u1_u1_n121 ) , .A1( u2_u1_u1_n98 ) );
  NAND2_X1 u2_u1_u1_U58 (.A1( u2_u1_u1_n103 ) , .ZN( u2_u1_u1_n153 ) , .A2( u2_u1_u1_n98 ) );
  NAND2_X1 u2_u1_u1_U59 (.A2( u2_u1_u1_n104 ) , .A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n133 ) );
  AOI22_X1 u2_u1_u1_U6 (.B2( u2_u1_u1_n113 ) , .A2( u2_u1_u1_n114 ) , .ZN( u2_u1_u1_n125 ) , .A1( u2_u1_u1_n171 ) , .B1( u2_u1_u1_n173 ) );
  NAND2_X1 u2_u1_u1_U60 (.ZN( u2_u1_u1_n150 ) , .A2( u2_u1_u1_n98 ) , .A1( u2_u1_u1_n99 ) );
  NAND2_X1 u2_u1_u1_U61 (.A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n155 ) , .A2( u2_u1_u1_n95 ) );
  OAI21_X1 u2_u1_u1_U62 (.ZN( u2_u1_u1_n109 ) , .B1( u2_u1_u1_n129 ) , .B2( u2_u1_u1_n160 ) , .A( u2_u1_u1_n167 ) );
  NAND2_X1 u2_u1_u1_U63 (.A2( u2_u1_u1_n100 ) , .A1( u2_u1_u1_n103 ) , .ZN( u2_u1_u1_n120 ) );
  NAND2_X1 u2_u1_u1_U64 (.A1( u2_u1_u1_n102 ) , .A2( u2_u1_u1_n104 ) , .ZN( u2_u1_u1_n115 ) );
  NAND2_X1 u2_u1_u1_U65 (.A2( u2_u1_u1_n100 ) , .A1( u2_u1_u1_n104 ) , .ZN( u2_u1_u1_n151 ) );
  NAND2_X1 u2_u1_u1_U66 (.A2( u2_u1_u1_n103 ) , .A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n161 ) );
  INV_X1 u2_u1_u1_U67 (.A( u2_u1_u1_n152 ) , .ZN( u2_u1_u1_n173 ) );
  INV_X1 u2_u1_u1_U68 (.A( u2_u1_u1_n128 ) , .ZN( u2_u1_u1_n172 ) );
  NAND2_X1 u2_u1_u1_U69 (.A2( u2_u1_u1_n102 ) , .A1( u2_u1_u1_n103 ) , .ZN( u2_u1_u1_n123 ) );
  NAND2_X1 u2_u1_u1_U7 (.ZN( u2_u1_u1_n114 ) , .A1( u2_u1_u1_n134 ) , .A2( u2_u1_u1_n156 ) );
  NOR2_X1 u2_u1_u1_U70 (.A2( u2_u1_X_7 ) , .A1( u2_u1_X_8 ) , .ZN( u2_u1_u1_n95 ) );
  NOR2_X1 u2_u1_u1_U71 (.A1( u2_u1_X_12 ) , .A2( u2_u1_X_9 ) , .ZN( u2_u1_u1_n100 ) );
  NOR2_X1 u2_u1_u1_U72 (.A2( u2_u1_X_8 ) , .A1( u2_u1_u1_n177 ) , .ZN( u2_u1_u1_n99 ) );
  NOR2_X1 u2_u1_u1_U73 (.A2( u2_u1_X_12 ) , .ZN( u2_u1_u1_n102 ) , .A1( u2_u1_u1_n176 ) );
  NOR2_X1 u2_u1_u1_U74 (.A2( u2_u1_X_9 ) , .ZN( u2_u1_u1_n105 ) , .A1( u2_u1_u1_n168 ) );
  NAND2_X1 u2_u1_u1_U75 (.A1( u2_u1_X_10 ) , .ZN( u2_u1_u1_n160 ) , .A2( u2_u1_u1_n169 ) );
  NAND2_X1 u2_u1_u1_U76 (.A2( u2_u1_X_10 ) , .A1( u2_u1_X_11 ) , .ZN( u2_u1_u1_n152 ) );
  NAND2_X1 u2_u1_u1_U77 (.A1( u2_u1_X_11 ) , .ZN( u2_u1_u1_n128 ) , .A2( u2_u1_u1_n170 ) );
  AND2_X1 u2_u1_u1_U78 (.A2( u2_u1_X_7 ) , .A1( u2_u1_X_8 ) , .ZN( u2_u1_u1_n104 ) );
  AND2_X1 u2_u1_u1_U79 (.A1( u2_u1_X_8 ) , .ZN( u2_u1_u1_n103 ) , .A2( u2_u1_u1_n177 ) );
  AOI22_X1 u2_u1_u1_U8 (.B2( u2_u1_u1_n136 ) , .A2( u2_u1_u1_n137 ) , .ZN( u2_u1_u1_n143 ) , .A1( u2_u1_u1_n171 ) , .B1( u2_u1_u1_n173 ) );
  INV_X1 u2_u1_u1_U80 (.A( u2_u1_X_10 ) , .ZN( u2_u1_u1_n170 ) );
  INV_X1 u2_u1_u1_U81 (.A( u2_u1_X_9 ) , .ZN( u2_u1_u1_n176 ) );
  INV_X1 u2_u1_u1_U82 (.A( u2_u1_X_11 ) , .ZN( u2_u1_u1_n169 ) );
  INV_X1 u2_u1_u1_U83 (.A( u2_u1_X_12 ) , .ZN( u2_u1_u1_n168 ) );
  INV_X1 u2_u1_u1_U84 (.A( u2_u1_X_7 ) , .ZN( u2_u1_u1_n177 ) );
  NAND4_X1 u2_u1_u1_U85 (.ZN( u2_out1_18 ) , .A4( u2_u1_u1_n165 ) , .A3( u2_u1_u1_n166 ) , .A1( u2_u1_u1_n167 ) , .A2( u2_u1_u1_n186 ) );
  AOI22_X1 u2_u1_u1_U86 (.B2( u2_u1_u1_n146 ) , .B1( u2_u1_u1_n147 ) , .A2( u2_u1_u1_n148 ) , .ZN( u2_u1_u1_n166 ) , .A1( u2_u1_u1_n172 ) );
  INV_X1 u2_u1_u1_U87 (.A( u2_u1_u1_n145 ) , .ZN( u2_u1_u1_n186 ) );
  NAND4_X1 u2_u1_u1_U88 (.ZN( u2_out1_2 ) , .A4( u2_u1_u1_n142 ) , .A3( u2_u1_u1_n143 ) , .A2( u2_u1_u1_n144 ) , .A1( u2_u1_u1_n179 ) );
  INV_X1 u2_u1_u1_U89 (.A( u2_u1_u1_n130 ) , .ZN( u2_u1_u1_n179 ) );
  INV_X1 u2_u1_u1_U9 (.A( u2_u1_u1_n147 ) , .ZN( u2_u1_u1_n181 ) );
  OAI21_X1 u2_u1_u1_U90 (.B2( u2_u1_u1_n132 ) , .ZN( u2_u1_u1_n144 ) , .A( u2_u1_u1_n146 ) , .B1( u2_u1_u1_n180 ) );
  NAND4_X1 u2_u1_u1_U91 (.ZN( u2_out1_28 ) , .A4( u2_u1_u1_n124 ) , .A3( u2_u1_u1_n125 ) , .A2( u2_u1_u1_n126 ) , .A1( u2_u1_u1_n127 ) );
  OAI21_X1 u2_u1_u1_U92 (.ZN( u2_u1_u1_n127 ) , .B2( u2_u1_u1_n139 ) , .B1( u2_u1_u1_n175 ) , .A( u2_u1_u1_n183 ) );
  OAI21_X1 u2_u1_u1_U93 (.ZN( u2_u1_u1_n126 ) , .B2( u2_u1_u1_n140 ) , .A( u2_u1_u1_n146 ) , .B1( u2_u1_u1_n178 ) );
  OR4_X1 u2_u1_u1_U94 (.ZN( u2_out1_13 ) , .A4( u2_u1_u1_n108 ) , .A3( u2_u1_u1_n109 ) , .A2( u2_u1_u1_n110 ) , .A1( u2_u1_u1_n111 ) );
  AOI21_X1 u2_u1_u1_U95 (.ZN( u2_u1_u1_n111 ) , .A( u2_u1_u1_n128 ) , .B2( u2_u1_u1_n131 ) , .B1( u2_u1_u1_n135 ) );
  AOI21_X1 u2_u1_u1_U96 (.ZN( u2_u1_u1_n110 ) , .A( u2_u1_u1_n116 ) , .B1( u2_u1_u1_n152 ) , .B2( u2_u1_u1_n160 ) );
  NAND3_X1 u2_u1_u1_U97 (.A3( u2_u1_u1_n149 ) , .A2( u2_u1_u1_n150 ) , .A1( u2_u1_u1_n151 ) , .ZN( u2_u1_u1_n164 ) );
  NAND3_X1 u2_u1_u1_U98 (.A3( u2_u1_u1_n134 ) , .A2( u2_u1_u1_n135 ) , .ZN( u2_u1_u1_n136 ) , .A1( u2_u1_u1_n151 ) );
  NAND3_X1 u2_u1_u1_U99 (.A1( u2_u1_u1_n133 ) , .ZN( u2_u1_u1_n137 ) , .A2( u2_u1_u1_n154 ) , .A3( u2_u1_u1_n181 ) );
  XOR2_X1 u2_u5_U13 (.B( u2_K6_42 ) , .A( u2_R4_29 ) , .Z( u2_u5_X_42 ) );
  XOR2_X1 u2_u5_U14 (.B( u2_K6_41 ) , .A( u2_R4_28 ) , .Z( u2_u5_X_41 ) );
  XOR2_X1 u2_u5_U15 (.B( u2_K6_40 ) , .A( u2_R4_27 ) , .Z( u2_u5_X_40 ) );
  XOR2_X1 u2_u5_U17 (.B( u2_K6_39 ) , .A( u2_R4_26 ) , .Z( u2_u5_X_39 ) );
  XOR2_X1 u2_u5_U18 (.B( u2_K6_38 ) , .A( u2_R4_25 ) , .Z( u2_u5_X_38 ) );
  XOR2_X1 u2_u5_U19 (.B( u2_K6_37 ) , .A( u2_R4_24 ) , .Z( u2_u5_X_37 ) );
  XOR2_X1 u2_u5_U20 (.B( u2_K6_36 ) , .A( u2_R4_25 ) , .Z( u2_u5_X_36 ) );
  XOR2_X1 u2_u5_U21 (.B( u2_K6_35 ) , .A( u2_R4_24 ) , .Z( u2_u5_X_35 ) );
  XOR2_X1 u2_u5_U22 (.B( u2_K6_34 ) , .A( u2_R4_23 ) , .Z( u2_u5_X_34 ) );
  XOR2_X1 u2_u5_U23 (.B( u2_K6_33 ) , .A( u2_R4_22 ) , .Z( u2_u5_X_33 ) );
  XOR2_X1 u2_u5_U24 (.B( u2_K6_32 ) , .A( u2_R4_21 ) , .Z( u2_u5_X_32 ) );
  XOR2_X1 u2_u5_U25 (.B( u2_K6_31 ) , .A( u2_R4_20 ) , .Z( u2_u5_X_31 ) );
  XOR2_X1 u2_u5_U33 (.B( u2_K6_24 ) , .A( u2_R4_17 ) , .Z( u2_u5_X_24 ) );
  XOR2_X1 u2_u5_U34 (.B( u2_K6_23 ) , .A( u2_R4_16 ) , .Z( u2_u5_X_23 ) );
  XOR2_X1 u2_u5_U35 (.B( u2_K6_22 ) , .A( u2_R4_15 ) , .Z( u2_u5_X_22 ) );
  XOR2_X1 u2_u5_U36 (.B( u2_K6_21 ) , .A( u2_R4_14 ) , .Z( u2_u5_X_21 ) );
  XOR2_X1 u2_u5_U37 (.B( u2_K6_20 ) , .A( u2_R4_13 ) , .Z( u2_u5_X_20 ) );
  XOR2_X1 u2_u5_U39 (.B( u2_K6_19 ) , .A( u2_R4_12 ) , .Z( u2_u5_X_19 ) );
  XOR2_X1 u2_u5_U40 (.B( u2_K6_18 ) , .A( u2_R4_13 ) , .Z( u2_u5_X_18 ) );
  XOR2_X1 u2_u5_U41 (.B( u2_K6_17 ) , .A( u2_R4_12 ) , .Z( u2_u5_X_17 ) );
  XOR2_X1 u2_u5_U42 (.B( u2_K6_16 ) , .A( u2_R4_11 ) , .Z( u2_u5_X_16 ) );
  XOR2_X1 u2_u5_U43 (.B( u2_K6_15 ) , .A( u2_R4_10 ) , .Z( u2_u5_X_15 ) );
  XOR2_X1 u2_u5_U44 (.B( u2_K6_14 ) , .A( u2_R4_9 ) , .Z( u2_u5_X_14 ) );
  XOR2_X1 u2_u5_U45 (.B( u2_K6_13 ) , .A( u2_R4_8 ) , .Z( u2_u5_X_13 ) );
  OAI22_X1 u2_u5_u2_U10 (.ZN( u2_u5_u2_n109 ) , .A2( u2_u5_u2_n113 ) , .B2( u2_u5_u2_n133 ) , .B1( u2_u5_u2_n167 ) , .A1( u2_u5_u2_n168 ) );
  NAND3_X1 u2_u5_u2_U100 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n98 ) );
  OAI22_X1 u2_u5_u2_U11 (.B1( u2_u5_u2_n151 ) , .A2( u2_u5_u2_n152 ) , .A1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n160 ) , .B2( u2_u5_u2_n168 ) );
  NOR3_X1 u2_u5_u2_U12 (.A1( u2_u5_u2_n150 ) , .ZN( u2_u5_u2_n151 ) , .A3( u2_u5_u2_n175 ) , .A2( u2_u5_u2_n188 ) );
  AOI21_X1 u2_u5_u2_U13 (.ZN( u2_u5_u2_n144 ) , .B2( u2_u5_u2_n155 ) , .A( u2_u5_u2_n172 ) , .B1( u2_u5_u2_n185 ) );
  AOI21_X1 u2_u5_u2_U14 (.B2( u2_u5_u2_n143 ) , .ZN( u2_u5_u2_n145 ) , .B1( u2_u5_u2_n152 ) , .A( u2_u5_u2_n171 ) );
  AOI21_X1 u2_u5_u2_U15 (.B2( u2_u5_u2_n120 ) , .B1( u2_u5_u2_n121 ) , .ZN( u2_u5_u2_n126 ) , .A( u2_u5_u2_n167 ) );
  INV_X1 u2_u5_u2_U16 (.A( u2_u5_u2_n156 ) , .ZN( u2_u5_u2_n171 ) );
  INV_X1 u2_u5_u2_U17 (.A( u2_u5_u2_n120 ) , .ZN( u2_u5_u2_n188 ) );
  NAND2_X1 u2_u5_u2_U18 (.A2( u2_u5_u2_n122 ) , .ZN( u2_u5_u2_n150 ) , .A1( u2_u5_u2_n152 ) );
  INV_X1 u2_u5_u2_U19 (.A( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n170 ) );
  INV_X1 u2_u5_u2_U20 (.A( u2_u5_u2_n137 ) , .ZN( u2_u5_u2_n173 ) );
  NAND2_X1 u2_u5_u2_U21 (.A1( u2_u5_u2_n132 ) , .A2( u2_u5_u2_n139 ) , .ZN( u2_u5_u2_n157 ) );
  INV_X1 u2_u5_u2_U22 (.A( u2_u5_u2_n113 ) , .ZN( u2_u5_u2_n178 ) );
  INV_X1 u2_u5_u2_U23 (.A( u2_u5_u2_n139 ) , .ZN( u2_u5_u2_n175 ) );
  INV_X1 u2_u5_u2_U24 (.A( u2_u5_u2_n155 ) , .ZN( u2_u5_u2_n181 ) );
  INV_X1 u2_u5_u2_U25 (.A( u2_u5_u2_n119 ) , .ZN( u2_u5_u2_n177 ) );
  INV_X1 u2_u5_u2_U26 (.A( u2_u5_u2_n116 ) , .ZN( u2_u5_u2_n180 ) );
  INV_X1 u2_u5_u2_U27 (.A( u2_u5_u2_n131 ) , .ZN( u2_u5_u2_n179 ) );
  INV_X1 u2_u5_u2_U28 (.A( u2_u5_u2_n154 ) , .ZN( u2_u5_u2_n176 ) );
  NAND2_X1 u2_u5_u2_U29 (.A2( u2_u5_u2_n116 ) , .A1( u2_u5_u2_n117 ) , .ZN( u2_u5_u2_n118 ) );
  NOR2_X1 u2_u5_u2_U3 (.ZN( u2_u5_u2_n121 ) , .A2( u2_u5_u2_n177 ) , .A1( u2_u5_u2_n180 ) );
  INV_X1 u2_u5_u2_U30 (.A( u2_u5_u2_n132 ) , .ZN( u2_u5_u2_n182 ) );
  INV_X1 u2_u5_u2_U31 (.A( u2_u5_u2_n158 ) , .ZN( u2_u5_u2_n183 ) );
  OAI21_X1 u2_u5_u2_U32 (.A( u2_u5_u2_n156 ) , .B1( u2_u5_u2_n157 ) , .ZN( u2_u5_u2_n158 ) , .B2( u2_u5_u2_n179 ) );
  NOR2_X1 u2_u5_u2_U33 (.ZN( u2_u5_u2_n156 ) , .A1( u2_u5_u2_n166 ) , .A2( u2_u5_u2_n169 ) );
  NOR2_X1 u2_u5_u2_U34 (.A2( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n137 ) , .A1( u2_u5_u2_n140 ) );
  NOR2_X1 u2_u5_u2_U35 (.A2( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n153 ) , .A1( u2_u5_u2_n156 ) );
  AOI211_X1 u2_u5_u2_U36 (.ZN( u2_u5_u2_n130 ) , .C1( u2_u5_u2_n138 ) , .C2( u2_u5_u2_n179 ) , .B( u2_u5_u2_n96 ) , .A( u2_u5_u2_n97 ) );
  OAI22_X1 u2_u5_u2_U37 (.B1( u2_u5_u2_n133 ) , .A2( u2_u5_u2_n137 ) , .A1( u2_u5_u2_n152 ) , .B2( u2_u5_u2_n168 ) , .ZN( u2_u5_u2_n97 ) );
  OAI221_X1 u2_u5_u2_U38 (.B1( u2_u5_u2_n113 ) , .C1( u2_u5_u2_n132 ) , .A( u2_u5_u2_n149 ) , .B2( u2_u5_u2_n171 ) , .C2( u2_u5_u2_n172 ) , .ZN( u2_u5_u2_n96 ) );
  OAI221_X1 u2_u5_u2_U39 (.A( u2_u5_u2_n115 ) , .C2( u2_u5_u2_n123 ) , .B2( u2_u5_u2_n143 ) , .B1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n163 ) , .C1( u2_u5_u2_n168 ) );
  INV_X1 u2_u5_u2_U4 (.A( u2_u5_u2_n134 ) , .ZN( u2_u5_u2_n185 ) );
  OAI21_X1 u2_u5_u2_U40 (.A( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n115 ) , .B1( u2_u5_u2_n176 ) , .B2( u2_u5_u2_n178 ) );
  OAI221_X1 u2_u5_u2_U41 (.A( u2_u5_u2_n135 ) , .B2( u2_u5_u2_n136 ) , .B1( u2_u5_u2_n137 ) , .ZN( u2_u5_u2_n162 ) , .C2( u2_u5_u2_n167 ) , .C1( u2_u5_u2_n185 ) );
  AND3_X1 u2_u5_u2_U42 (.A3( u2_u5_u2_n131 ) , .A2( u2_u5_u2_n132 ) , .A1( u2_u5_u2_n133 ) , .ZN( u2_u5_u2_n136 ) );
  AOI22_X1 u2_u5_u2_U43 (.ZN( u2_u5_u2_n135 ) , .B1( u2_u5_u2_n140 ) , .A1( u2_u5_u2_n156 ) , .B2( u2_u5_u2_n180 ) , .A2( u2_u5_u2_n188 ) );
  AOI21_X1 u2_u5_u2_U44 (.ZN( u2_u5_u2_n149 ) , .B1( u2_u5_u2_n173 ) , .B2( u2_u5_u2_n188 ) , .A( u2_u5_u2_n95 ) );
  AND3_X1 u2_u5_u2_U45 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n156 ) , .ZN( u2_u5_u2_n95 ) );
  OAI21_X1 u2_u5_u2_U46 (.A( u2_u5_u2_n141 ) , .B2( u2_u5_u2_n142 ) , .ZN( u2_u5_u2_n146 ) , .B1( u2_u5_u2_n153 ) );
  OAI21_X1 u2_u5_u2_U47 (.A( u2_u5_u2_n140 ) , .ZN( u2_u5_u2_n141 ) , .B1( u2_u5_u2_n176 ) , .B2( u2_u5_u2_n177 ) );
  NOR3_X1 u2_u5_u2_U48 (.ZN( u2_u5_u2_n142 ) , .A3( u2_u5_u2_n175 ) , .A2( u2_u5_u2_n178 ) , .A1( u2_u5_u2_n181 ) );
  OAI21_X1 u2_u5_u2_U49 (.A( u2_u5_u2_n101 ) , .B2( u2_u5_u2_n121 ) , .B1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n164 ) );
  INV_X1 u2_u5_u2_U5 (.A( u2_u5_u2_n150 ) , .ZN( u2_u5_u2_n184 ) );
  NAND2_X1 u2_u5_u2_U50 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n155 ) );
  NAND2_X1 u2_u5_u2_U51 (.A2( u2_u5_u2_n105 ) , .A1( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n143 ) );
  NAND2_X1 u2_u5_u2_U52 (.A1( u2_u5_u2_n104 ) , .A2( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n152 ) );
  NAND2_X1 u2_u5_u2_U53 (.A1( u2_u5_u2_n100 ) , .A2( u2_u5_u2_n105 ) , .ZN( u2_u5_u2_n132 ) );
  INV_X1 u2_u5_u2_U54 (.A( u2_u5_u2_n140 ) , .ZN( u2_u5_u2_n168 ) );
  INV_X1 u2_u5_u2_U55 (.A( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n167 ) );
  NAND2_X1 u2_u5_u2_U56 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n113 ) );
  NAND2_X1 u2_u5_u2_U57 (.A1( u2_u5_u2_n106 ) , .A2( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n131 ) );
  NAND2_X1 u2_u5_u2_U58 (.A1( u2_u5_u2_n103 ) , .A2( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n139 ) );
  NAND2_X1 u2_u5_u2_U59 (.A1( u2_u5_u2_n103 ) , .A2( u2_u5_u2_n105 ) , .ZN( u2_u5_u2_n133 ) );
  NOR4_X1 u2_u5_u2_U6 (.A4( u2_u5_u2_n124 ) , .A3( u2_u5_u2_n125 ) , .A2( u2_u5_u2_n126 ) , .A1( u2_u5_u2_n127 ) , .ZN( u2_u5_u2_n128 ) );
  NAND2_X1 u2_u5_u2_U60 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n103 ) , .ZN( u2_u5_u2_n154 ) );
  NAND2_X1 u2_u5_u2_U61 (.A2( u2_u5_u2_n103 ) , .A1( u2_u5_u2_n104 ) , .ZN( u2_u5_u2_n119 ) );
  NAND2_X1 u2_u5_u2_U62 (.A2( u2_u5_u2_n107 ) , .A1( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n123 ) );
  NAND2_X1 u2_u5_u2_U63 (.A1( u2_u5_u2_n104 ) , .A2( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n122 ) );
  INV_X1 u2_u5_u2_U64 (.A( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n172 ) );
  NAND2_X1 u2_u5_u2_U65 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n102 ) , .ZN( u2_u5_u2_n116 ) );
  NAND2_X1 u2_u5_u2_U66 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n120 ) );
  NAND2_X1 u2_u5_u2_U67 (.A2( u2_u5_u2_n105 ) , .A1( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n117 ) );
  INV_X1 u2_u5_u2_U68 (.ZN( u2_u5_u2_n187 ) , .A( u2_u5_u2_n99 ) );
  OAI21_X1 u2_u5_u2_U69 (.B1( u2_u5_u2_n137 ) , .B2( u2_u5_u2_n143 ) , .A( u2_u5_u2_n98 ) , .ZN( u2_u5_u2_n99 ) );
  AOI21_X1 u2_u5_u2_U7 (.B2( u2_u5_u2_n119 ) , .ZN( u2_u5_u2_n127 ) , .A( u2_u5_u2_n137 ) , .B1( u2_u5_u2_n155 ) );
  NOR2_X1 u2_u5_u2_U70 (.A2( u2_u5_X_16 ) , .ZN( u2_u5_u2_n140 ) , .A1( u2_u5_u2_n166 ) );
  NOR2_X1 u2_u5_u2_U71 (.A2( u2_u5_X_13 ) , .A1( u2_u5_X_14 ) , .ZN( u2_u5_u2_n100 ) );
  NOR2_X1 u2_u5_u2_U72 (.A2( u2_u5_X_16 ) , .A1( u2_u5_X_17 ) , .ZN( u2_u5_u2_n138 ) );
  NOR2_X1 u2_u5_u2_U73 (.A2( u2_u5_X_15 ) , .A1( u2_u5_X_18 ) , .ZN( u2_u5_u2_n104 ) );
  NOR2_X1 u2_u5_u2_U74 (.A2( u2_u5_X_14 ) , .ZN( u2_u5_u2_n103 ) , .A1( u2_u5_u2_n174 ) );
  NOR2_X1 u2_u5_u2_U75 (.A2( u2_u5_X_15 ) , .ZN( u2_u5_u2_n102 ) , .A1( u2_u5_u2_n165 ) );
  NOR2_X1 u2_u5_u2_U76 (.A2( u2_u5_X_17 ) , .ZN( u2_u5_u2_n114 ) , .A1( u2_u5_u2_n169 ) );
  AND2_X1 u2_u5_u2_U77 (.A1( u2_u5_X_15 ) , .ZN( u2_u5_u2_n105 ) , .A2( u2_u5_u2_n165 ) );
  AND2_X1 u2_u5_u2_U78 (.A2( u2_u5_X_15 ) , .A1( u2_u5_X_18 ) , .ZN( u2_u5_u2_n107 ) );
  AND2_X1 u2_u5_u2_U79 (.A1( u2_u5_X_14 ) , .ZN( u2_u5_u2_n106 ) , .A2( u2_u5_u2_n174 ) );
  AOI21_X1 u2_u5_u2_U8 (.ZN( u2_u5_u2_n124 ) , .B1( u2_u5_u2_n131 ) , .B2( u2_u5_u2_n143 ) , .A( u2_u5_u2_n172 ) );
  AND2_X1 u2_u5_u2_U80 (.A1( u2_u5_X_13 ) , .A2( u2_u5_X_14 ) , .ZN( u2_u5_u2_n108 ) );
  INV_X1 u2_u5_u2_U81 (.A( u2_u5_X_16 ) , .ZN( u2_u5_u2_n169 ) );
  INV_X1 u2_u5_u2_U82 (.A( u2_u5_X_17 ) , .ZN( u2_u5_u2_n166 ) );
  INV_X1 u2_u5_u2_U83 (.A( u2_u5_X_13 ) , .ZN( u2_u5_u2_n174 ) );
  INV_X1 u2_u5_u2_U84 (.A( u2_u5_X_18 ) , .ZN( u2_u5_u2_n165 ) );
  NAND4_X1 u2_u5_u2_U85 (.ZN( u2_out5_24 ) , .A4( u2_u5_u2_n111 ) , .A3( u2_u5_u2_n112 ) , .A1( u2_u5_u2_n130 ) , .A2( u2_u5_u2_n187 ) );
  AOI221_X1 u2_u5_u2_U86 (.A( u2_u5_u2_n109 ) , .B1( u2_u5_u2_n110 ) , .ZN( u2_u5_u2_n111 ) , .C1( u2_u5_u2_n134 ) , .C2( u2_u5_u2_n170 ) , .B2( u2_u5_u2_n173 ) );
  AOI21_X1 u2_u5_u2_U87 (.ZN( u2_u5_u2_n112 ) , .B2( u2_u5_u2_n156 ) , .A( u2_u5_u2_n164 ) , .B1( u2_u5_u2_n181 ) );
  NAND4_X1 u2_u5_u2_U88 (.ZN( u2_out5_16 ) , .A4( u2_u5_u2_n128 ) , .A3( u2_u5_u2_n129 ) , .A1( u2_u5_u2_n130 ) , .A2( u2_u5_u2_n186 ) );
  AOI22_X1 u2_u5_u2_U89 (.A2( u2_u5_u2_n118 ) , .ZN( u2_u5_u2_n129 ) , .A1( u2_u5_u2_n140 ) , .B1( u2_u5_u2_n157 ) , .B2( u2_u5_u2_n170 ) );
  AOI21_X1 u2_u5_u2_U9 (.B2( u2_u5_u2_n123 ) , .ZN( u2_u5_u2_n125 ) , .A( u2_u5_u2_n171 ) , .B1( u2_u5_u2_n184 ) );
  INV_X1 u2_u5_u2_U90 (.A( u2_u5_u2_n163 ) , .ZN( u2_u5_u2_n186 ) );
  NAND4_X1 u2_u5_u2_U91 (.ZN( u2_out5_30 ) , .A4( u2_u5_u2_n147 ) , .A3( u2_u5_u2_n148 ) , .A2( u2_u5_u2_n149 ) , .A1( u2_u5_u2_n187 ) );
  NOR3_X1 u2_u5_u2_U92 (.A3( u2_u5_u2_n144 ) , .A2( u2_u5_u2_n145 ) , .A1( u2_u5_u2_n146 ) , .ZN( u2_u5_u2_n147 ) );
  AOI21_X1 u2_u5_u2_U93 (.B2( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n148 ) , .A( u2_u5_u2_n162 ) , .B1( u2_u5_u2_n182 ) );
  OR4_X1 u2_u5_u2_U94 (.ZN( u2_out5_6 ) , .A4( u2_u5_u2_n161 ) , .A3( u2_u5_u2_n162 ) , .A2( u2_u5_u2_n163 ) , .A1( u2_u5_u2_n164 ) );
  OR3_X1 u2_u5_u2_U95 (.A2( u2_u5_u2_n159 ) , .A1( u2_u5_u2_n160 ) , .ZN( u2_u5_u2_n161 ) , .A3( u2_u5_u2_n183 ) );
  AOI21_X1 u2_u5_u2_U96 (.B2( u2_u5_u2_n154 ) , .B1( u2_u5_u2_n155 ) , .ZN( u2_u5_u2_n159 ) , .A( u2_u5_u2_n167 ) );
  NAND3_X1 u2_u5_u2_U97 (.A2( u2_u5_u2_n117 ) , .A1( u2_u5_u2_n122 ) , .A3( u2_u5_u2_n123 ) , .ZN( u2_u5_u2_n134 ) );
  NAND3_X1 u2_u5_u2_U98 (.ZN( u2_u5_u2_n110 ) , .A2( u2_u5_u2_n131 ) , .A3( u2_u5_u2_n139 ) , .A1( u2_u5_u2_n154 ) );
  NAND3_X1 u2_u5_u2_U99 (.A2( u2_u5_u2_n100 ) , .ZN( u2_u5_u2_n101 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n114 ) );
  OAI22_X1 u2_u5_u3_U10 (.B1( u2_u5_u3_n113 ) , .A2( u2_u5_u3_n135 ) , .A1( u2_u5_u3_n150 ) , .B2( u2_u5_u3_n164 ) , .ZN( u2_u5_u3_n98 ) );
  OAI211_X1 u2_u5_u3_U11 (.B( u2_u5_u3_n106 ) , .ZN( u2_u5_u3_n119 ) , .C2( u2_u5_u3_n128 ) , .C1( u2_u5_u3_n167 ) , .A( u2_u5_u3_n181 ) );
  AOI221_X1 u2_u5_u3_U12 (.C1( u2_u5_u3_n105 ) , .ZN( u2_u5_u3_n106 ) , .A( u2_u5_u3_n131 ) , .B2( u2_u5_u3_n132 ) , .C2( u2_u5_u3_n133 ) , .B1( u2_u5_u3_n169 ) );
  INV_X1 u2_u5_u3_U13 (.ZN( u2_u5_u3_n181 ) , .A( u2_u5_u3_n98 ) );
  NAND2_X1 u2_u5_u3_U14 (.ZN( u2_u5_u3_n105 ) , .A2( u2_u5_u3_n130 ) , .A1( u2_u5_u3_n155 ) );
  AOI22_X1 u2_u5_u3_U15 (.B1( u2_u5_u3_n115 ) , .A2( u2_u5_u3_n116 ) , .ZN( u2_u5_u3_n123 ) , .B2( u2_u5_u3_n133 ) , .A1( u2_u5_u3_n169 ) );
  NAND2_X1 u2_u5_u3_U16 (.ZN( u2_u5_u3_n116 ) , .A2( u2_u5_u3_n151 ) , .A1( u2_u5_u3_n182 ) );
  NOR2_X1 u2_u5_u3_U17 (.ZN( u2_u5_u3_n126 ) , .A2( u2_u5_u3_n150 ) , .A1( u2_u5_u3_n164 ) );
  AOI21_X1 u2_u5_u3_U18 (.ZN( u2_u5_u3_n112 ) , .B2( u2_u5_u3_n146 ) , .B1( u2_u5_u3_n155 ) , .A( u2_u5_u3_n167 ) );
  NAND2_X1 u2_u5_u3_U19 (.A1( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n142 ) , .A2( u2_u5_u3_n164 ) );
  NAND2_X1 u2_u5_u3_U20 (.ZN( u2_u5_u3_n132 ) , .A2( u2_u5_u3_n152 ) , .A1( u2_u5_u3_n156 ) );
  AND2_X1 u2_u5_u3_U21 (.A2( u2_u5_u3_n113 ) , .A1( u2_u5_u3_n114 ) , .ZN( u2_u5_u3_n151 ) );
  INV_X1 u2_u5_u3_U22 (.A( u2_u5_u3_n133 ) , .ZN( u2_u5_u3_n165 ) );
  INV_X1 u2_u5_u3_U23 (.A( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n170 ) );
  NAND2_X1 u2_u5_u3_U24 (.A1( u2_u5_u3_n107 ) , .A2( u2_u5_u3_n108 ) , .ZN( u2_u5_u3_n140 ) );
  NAND2_X1 u2_u5_u3_U25 (.ZN( u2_u5_u3_n117 ) , .A1( u2_u5_u3_n124 ) , .A2( u2_u5_u3_n148 ) );
  NAND2_X1 u2_u5_u3_U26 (.ZN( u2_u5_u3_n143 ) , .A1( u2_u5_u3_n165 ) , .A2( u2_u5_u3_n167 ) );
  INV_X1 u2_u5_u3_U27 (.A( u2_u5_u3_n130 ) , .ZN( u2_u5_u3_n177 ) );
  INV_X1 u2_u5_u3_U28 (.A( u2_u5_u3_n128 ) , .ZN( u2_u5_u3_n176 ) );
  INV_X1 u2_u5_u3_U29 (.A( u2_u5_u3_n155 ) , .ZN( u2_u5_u3_n174 ) );
  INV_X1 u2_u5_u3_U3 (.A( u2_u5_u3_n129 ) , .ZN( u2_u5_u3_n183 ) );
  INV_X1 u2_u5_u3_U30 (.A( u2_u5_u3_n139 ) , .ZN( u2_u5_u3_n185 ) );
  NOR2_X1 u2_u5_u3_U31 (.ZN( u2_u5_u3_n135 ) , .A2( u2_u5_u3_n141 ) , .A1( u2_u5_u3_n169 ) );
  OAI222_X1 u2_u5_u3_U32 (.C2( u2_u5_u3_n107 ) , .A2( u2_u5_u3_n108 ) , .B1( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n138 ) , .B2( u2_u5_u3_n146 ) , .C1( u2_u5_u3_n154 ) , .A1( u2_u5_u3_n164 ) );
  NOR4_X1 u2_u5_u3_U33 (.A4( u2_u5_u3_n157 ) , .A3( u2_u5_u3_n158 ) , .A2( u2_u5_u3_n159 ) , .A1( u2_u5_u3_n160 ) , .ZN( u2_u5_u3_n161 ) );
  AOI21_X1 u2_u5_u3_U34 (.B2( u2_u5_u3_n152 ) , .B1( u2_u5_u3_n153 ) , .ZN( u2_u5_u3_n158 ) , .A( u2_u5_u3_n164 ) );
  AOI21_X1 u2_u5_u3_U35 (.A( u2_u5_u3_n154 ) , .B2( u2_u5_u3_n155 ) , .B1( u2_u5_u3_n156 ) , .ZN( u2_u5_u3_n157 ) );
  AOI21_X1 u2_u5_u3_U36 (.A( u2_u5_u3_n149 ) , .B2( u2_u5_u3_n150 ) , .B1( u2_u5_u3_n151 ) , .ZN( u2_u5_u3_n159 ) );
  AOI211_X1 u2_u5_u3_U37 (.ZN( u2_u5_u3_n109 ) , .A( u2_u5_u3_n119 ) , .C2( u2_u5_u3_n129 ) , .B( u2_u5_u3_n138 ) , .C1( u2_u5_u3_n141 ) );
  AOI211_X1 u2_u5_u3_U38 (.B( u2_u5_u3_n119 ) , .A( u2_u5_u3_n120 ) , .C2( u2_u5_u3_n121 ) , .ZN( u2_u5_u3_n122 ) , .C1( u2_u5_u3_n179 ) );
  INV_X1 u2_u5_u3_U39 (.A( u2_u5_u3_n156 ) , .ZN( u2_u5_u3_n179 ) );
  INV_X1 u2_u5_u3_U4 (.A( u2_u5_u3_n140 ) , .ZN( u2_u5_u3_n182 ) );
  OAI22_X1 u2_u5_u3_U40 (.B1( u2_u5_u3_n118 ) , .ZN( u2_u5_u3_n120 ) , .A1( u2_u5_u3_n135 ) , .B2( u2_u5_u3_n154 ) , .A2( u2_u5_u3_n178 ) );
  AND3_X1 u2_u5_u3_U41 (.ZN( u2_u5_u3_n118 ) , .A2( u2_u5_u3_n124 ) , .A1( u2_u5_u3_n144 ) , .A3( u2_u5_u3_n152 ) );
  INV_X1 u2_u5_u3_U42 (.A( u2_u5_u3_n121 ) , .ZN( u2_u5_u3_n164 ) );
  NAND2_X1 u2_u5_u3_U43 (.ZN( u2_u5_u3_n133 ) , .A1( u2_u5_u3_n154 ) , .A2( u2_u5_u3_n164 ) );
  OAI211_X1 u2_u5_u3_U44 (.B( u2_u5_u3_n127 ) , .ZN( u2_u5_u3_n139 ) , .C1( u2_u5_u3_n150 ) , .C2( u2_u5_u3_n154 ) , .A( u2_u5_u3_n184 ) );
  INV_X1 u2_u5_u3_U45 (.A( u2_u5_u3_n125 ) , .ZN( u2_u5_u3_n184 ) );
  AOI221_X1 u2_u5_u3_U46 (.A( u2_u5_u3_n126 ) , .ZN( u2_u5_u3_n127 ) , .C2( u2_u5_u3_n132 ) , .C1( u2_u5_u3_n169 ) , .B2( u2_u5_u3_n170 ) , .B1( u2_u5_u3_n174 ) );
  OAI22_X1 u2_u5_u3_U47 (.A1( u2_u5_u3_n124 ) , .ZN( u2_u5_u3_n125 ) , .B2( u2_u5_u3_n145 ) , .A2( u2_u5_u3_n165 ) , .B1( u2_u5_u3_n167 ) );
  NOR2_X1 u2_u5_u3_U48 (.A1( u2_u5_u3_n113 ) , .ZN( u2_u5_u3_n131 ) , .A2( u2_u5_u3_n154 ) );
  NAND2_X1 u2_u5_u3_U49 (.A1( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n150 ) , .A2( u2_u5_u3_n99 ) );
  INV_X1 u2_u5_u3_U5 (.A( u2_u5_u3_n117 ) , .ZN( u2_u5_u3_n178 ) );
  NAND2_X1 u2_u5_u3_U50 (.A2( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n155 ) , .A1( u2_u5_u3_n97 ) );
  INV_X1 u2_u5_u3_U51 (.A( u2_u5_u3_n141 ) , .ZN( u2_u5_u3_n167 ) );
  AOI21_X1 u2_u5_u3_U52 (.B2( u2_u5_u3_n114 ) , .B1( u2_u5_u3_n146 ) , .A( u2_u5_u3_n154 ) , .ZN( u2_u5_u3_n94 ) );
  AOI21_X1 u2_u5_u3_U53 (.ZN( u2_u5_u3_n110 ) , .B2( u2_u5_u3_n142 ) , .B1( u2_u5_u3_n186 ) , .A( u2_u5_u3_n95 ) );
  INV_X1 u2_u5_u3_U54 (.A( u2_u5_u3_n145 ) , .ZN( u2_u5_u3_n186 ) );
  AOI21_X1 u2_u5_u3_U55 (.B1( u2_u5_u3_n124 ) , .A( u2_u5_u3_n149 ) , .B2( u2_u5_u3_n155 ) , .ZN( u2_u5_u3_n95 ) );
  INV_X1 u2_u5_u3_U56 (.A( u2_u5_u3_n149 ) , .ZN( u2_u5_u3_n169 ) );
  NAND2_X1 u2_u5_u3_U57 (.ZN( u2_u5_u3_n124 ) , .A1( u2_u5_u3_n96 ) , .A2( u2_u5_u3_n97 ) );
  NAND2_X1 u2_u5_u3_U58 (.A2( u2_u5_u3_n100 ) , .ZN( u2_u5_u3_n146 ) , .A1( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U59 (.A1( u2_u5_u3_n101 ) , .ZN( u2_u5_u3_n145 ) , .A2( u2_u5_u3_n99 ) );
  AOI221_X1 u2_u5_u3_U6 (.A( u2_u5_u3_n131 ) , .C2( u2_u5_u3_n132 ) , .C1( u2_u5_u3_n133 ) , .ZN( u2_u5_u3_n134 ) , .B1( u2_u5_u3_n143 ) , .B2( u2_u5_u3_n177 ) );
  NAND2_X1 u2_u5_u3_U60 (.A1( u2_u5_u3_n100 ) , .ZN( u2_u5_u3_n156 ) , .A2( u2_u5_u3_n99 ) );
  NAND2_X1 u2_u5_u3_U61 (.A2( u2_u5_u3_n101 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n148 ) );
  NAND2_X1 u2_u5_u3_U62 (.A1( u2_u5_u3_n100 ) , .A2( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n128 ) );
  NAND2_X1 u2_u5_u3_U63 (.A2( u2_u5_u3_n101 ) , .A1( u2_u5_u3_n102 ) , .ZN( u2_u5_u3_n152 ) );
  NAND2_X1 u2_u5_u3_U64 (.A2( u2_u5_u3_n101 ) , .ZN( u2_u5_u3_n114 ) , .A1( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U65 (.ZN( u2_u5_u3_n107 ) , .A1( u2_u5_u3_n97 ) , .A2( u2_u5_u3_n99 ) );
  NAND2_X1 u2_u5_u3_U66 (.A2( u2_u5_u3_n100 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n113 ) );
  NAND2_X1 u2_u5_u3_U67 (.A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n153 ) , .A2( u2_u5_u3_n97 ) );
  NAND2_X1 u2_u5_u3_U68 (.A2( u2_u5_u3_n103 ) , .A1( u2_u5_u3_n104 ) , .ZN( u2_u5_u3_n130 ) );
  NAND2_X1 u2_u5_u3_U69 (.A2( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n144 ) , .A1( u2_u5_u3_n96 ) );
  OAI22_X1 u2_u5_u3_U7 (.B2( u2_u5_u3_n147 ) , .A2( u2_u5_u3_n148 ) , .ZN( u2_u5_u3_n160 ) , .B1( u2_u5_u3_n165 ) , .A1( u2_u5_u3_n168 ) );
  NAND2_X1 u2_u5_u3_U70 (.A1( u2_u5_u3_n102 ) , .A2( u2_u5_u3_n103 ) , .ZN( u2_u5_u3_n108 ) );
  NOR2_X1 u2_u5_u3_U71 (.A2( u2_u5_X_19 ) , .A1( u2_u5_X_20 ) , .ZN( u2_u5_u3_n99 ) );
  NOR2_X1 u2_u5_u3_U72 (.A2( u2_u5_X_21 ) , .A1( u2_u5_X_24 ) , .ZN( u2_u5_u3_n103 ) );
  NOR2_X1 u2_u5_u3_U73 (.A2( u2_u5_X_24 ) , .A1( u2_u5_u3_n171 ) , .ZN( u2_u5_u3_n97 ) );
  NOR2_X1 u2_u5_u3_U74 (.A2( u2_u5_X_23 ) , .ZN( u2_u5_u3_n141 ) , .A1( u2_u5_u3_n166 ) );
  NOR2_X1 u2_u5_u3_U75 (.A2( u2_u5_X_19 ) , .A1( u2_u5_u3_n172 ) , .ZN( u2_u5_u3_n96 ) );
  NAND2_X1 u2_u5_u3_U76 (.A1( u2_u5_X_22 ) , .A2( u2_u5_X_23 ) , .ZN( u2_u5_u3_n154 ) );
  NAND2_X1 u2_u5_u3_U77 (.A1( u2_u5_X_23 ) , .ZN( u2_u5_u3_n149 ) , .A2( u2_u5_u3_n166 ) );
  NOR2_X1 u2_u5_u3_U78 (.A2( u2_u5_X_22 ) , .A1( u2_u5_X_23 ) , .ZN( u2_u5_u3_n121 ) );
  AND2_X1 u2_u5_u3_U79 (.A1( u2_u5_X_24 ) , .ZN( u2_u5_u3_n101 ) , .A2( u2_u5_u3_n171 ) );
  AND3_X1 u2_u5_u3_U8 (.A3( u2_u5_u3_n144 ) , .A2( u2_u5_u3_n145 ) , .A1( u2_u5_u3_n146 ) , .ZN( u2_u5_u3_n147 ) );
  AND2_X1 u2_u5_u3_U80 (.A1( u2_u5_X_19 ) , .ZN( u2_u5_u3_n102 ) , .A2( u2_u5_u3_n172 ) );
  AND2_X1 u2_u5_u3_U81 (.A1( u2_u5_X_21 ) , .A2( u2_u5_X_24 ) , .ZN( u2_u5_u3_n100 ) );
  AND2_X1 u2_u5_u3_U82 (.A2( u2_u5_X_19 ) , .A1( u2_u5_X_20 ) , .ZN( u2_u5_u3_n104 ) );
  INV_X1 u2_u5_u3_U83 (.A( u2_u5_X_22 ) , .ZN( u2_u5_u3_n166 ) );
  INV_X1 u2_u5_u3_U84 (.A( u2_u5_X_21 ) , .ZN( u2_u5_u3_n171 ) );
  INV_X1 u2_u5_u3_U85 (.A( u2_u5_X_20 ) , .ZN( u2_u5_u3_n172 ) );
  NAND4_X1 u2_u5_u3_U86 (.ZN( u2_out5_26 ) , .A4( u2_u5_u3_n109 ) , .A3( u2_u5_u3_n110 ) , .A2( u2_u5_u3_n111 ) , .A1( u2_u5_u3_n173 ) );
  INV_X1 u2_u5_u3_U87 (.ZN( u2_u5_u3_n173 ) , .A( u2_u5_u3_n94 ) );
  OAI21_X1 u2_u5_u3_U88 (.ZN( u2_u5_u3_n111 ) , .B2( u2_u5_u3_n117 ) , .A( u2_u5_u3_n133 ) , .B1( u2_u5_u3_n176 ) );
  NAND4_X1 u2_u5_u3_U89 (.ZN( u2_out5_20 ) , .A4( u2_u5_u3_n122 ) , .A3( u2_u5_u3_n123 ) , .A1( u2_u5_u3_n175 ) , .A2( u2_u5_u3_n180 ) );
  INV_X1 u2_u5_u3_U9 (.A( u2_u5_u3_n143 ) , .ZN( u2_u5_u3_n168 ) );
  INV_X1 u2_u5_u3_U90 (.A( u2_u5_u3_n126 ) , .ZN( u2_u5_u3_n180 ) );
  INV_X1 u2_u5_u3_U91 (.A( u2_u5_u3_n112 ) , .ZN( u2_u5_u3_n175 ) );
  NAND4_X1 u2_u5_u3_U92 (.ZN( u2_out5_1 ) , .A4( u2_u5_u3_n161 ) , .A3( u2_u5_u3_n162 ) , .A2( u2_u5_u3_n163 ) , .A1( u2_u5_u3_n185 ) );
  NAND2_X1 u2_u5_u3_U93 (.ZN( u2_u5_u3_n163 ) , .A2( u2_u5_u3_n170 ) , .A1( u2_u5_u3_n176 ) );
  AOI22_X1 u2_u5_u3_U94 (.B2( u2_u5_u3_n140 ) , .B1( u2_u5_u3_n141 ) , .A2( u2_u5_u3_n142 ) , .ZN( u2_u5_u3_n162 ) , .A1( u2_u5_u3_n177 ) );
  OR4_X1 u2_u5_u3_U95 (.ZN( u2_out5_10 ) , .A4( u2_u5_u3_n136 ) , .A3( u2_u5_u3_n137 ) , .A1( u2_u5_u3_n138 ) , .A2( u2_u5_u3_n139 ) );
  OAI222_X1 u2_u5_u3_U96 (.C1( u2_u5_u3_n128 ) , .ZN( u2_u5_u3_n137 ) , .B1( u2_u5_u3_n148 ) , .A2( u2_u5_u3_n150 ) , .B2( u2_u5_u3_n154 ) , .C2( u2_u5_u3_n164 ) , .A1( u2_u5_u3_n167 ) );
  OAI221_X1 u2_u5_u3_U97 (.A( u2_u5_u3_n134 ) , .B2( u2_u5_u3_n135 ) , .ZN( u2_u5_u3_n136 ) , .C1( u2_u5_u3_n149 ) , .B1( u2_u5_u3_n151 ) , .C2( u2_u5_u3_n183 ) );
  NAND3_X1 u2_u5_u3_U98 (.A1( u2_u5_u3_n114 ) , .ZN( u2_u5_u3_n115 ) , .A2( u2_u5_u3_n145 ) , .A3( u2_u5_u3_n153 ) );
  NAND3_X1 u2_u5_u3_U99 (.ZN( u2_u5_u3_n129 ) , .A2( u2_u5_u3_n144 ) , .A1( u2_u5_u3_n153 ) , .A3( u2_u5_u3_n182 ) );
  INV_X1 u2_u5_u5_U10 (.A( u2_u5_u5_n121 ) , .ZN( u2_u5_u5_n177 ) );
  NOR3_X1 u2_u5_u5_U100 (.A3( u2_u5_u5_n141 ) , .A1( u2_u5_u5_n142 ) , .ZN( u2_u5_u5_n143 ) , .A2( u2_u5_u5_n191 ) );
  NAND4_X1 u2_u5_u5_U101 (.ZN( u2_out5_4 ) , .A4( u2_u5_u5_n112 ) , .A2( u2_u5_u5_n113 ) , .A1( u2_u5_u5_n114 ) , .A3( u2_u5_u5_n195 ) );
  AOI211_X1 u2_u5_u5_U102 (.A( u2_u5_u5_n110 ) , .C1( u2_u5_u5_n111 ) , .ZN( u2_u5_u5_n112 ) , .B( u2_u5_u5_n118 ) , .C2( u2_u5_u5_n177 ) );
  AOI222_X1 u2_u5_u5_U103 (.ZN( u2_u5_u5_n113 ) , .A1( u2_u5_u5_n131 ) , .C1( u2_u5_u5_n148 ) , .B2( u2_u5_u5_n174 ) , .C2( u2_u5_u5_n178 ) , .A2( u2_u5_u5_n179 ) , .B1( u2_u5_u5_n99 ) );
  NAND3_X1 u2_u5_u5_U104 (.A2( u2_u5_u5_n154 ) , .A3( u2_u5_u5_n158 ) , .A1( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n99 ) );
  NOR2_X1 u2_u5_u5_U11 (.ZN( u2_u5_u5_n160 ) , .A2( u2_u5_u5_n173 ) , .A1( u2_u5_u5_n177 ) );
  INV_X1 u2_u5_u5_U12 (.A( u2_u5_u5_n150 ) , .ZN( u2_u5_u5_n174 ) );
  AOI21_X1 u2_u5_u5_U13 (.A( u2_u5_u5_n160 ) , .B2( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n162 ) , .B1( u2_u5_u5_n192 ) );
  INV_X1 u2_u5_u5_U14 (.A( u2_u5_u5_n159 ) , .ZN( u2_u5_u5_n192 ) );
  AOI21_X1 u2_u5_u5_U15 (.A( u2_u5_u5_n156 ) , .B2( u2_u5_u5_n157 ) , .B1( u2_u5_u5_n158 ) , .ZN( u2_u5_u5_n163 ) );
  AOI21_X1 u2_u5_u5_U16 (.B2( u2_u5_u5_n139 ) , .B1( u2_u5_u5_n140 ) , .ZN( u2_u5_u5_n141 ) , .A( u2_u5_u5_n150 ) );
  OAI21_X1 u2_u5_u5_U17 (.A( u2_u5_u5_n133 ) , .B2( u2_u5_u5_n134 ) , .B1( u2_u5_u5_n135 ) , .ZN( u2_u5_u5_n142 ) );
  OAI21_X1 u2_u5_u5_U18 (.ZN( u2_u5_u5_n133 ) , .B2( u2_u5_u5_n147 ) , .A( u2_u5_u5_n173 ) , .B1( u2_u5_u5_n188 ) );
  NAND2_X1 u2_u5_u5_U19 (.A2( u2_u5_u5_n119 ) , .A1( u2_u5_u5_n123 ) , .ZN( u2_u5_u5_n137 ) );
  INV_X1 u2_u5_u5_U20 (.A( u2_u5_u5_n155 ) , .ZN( u2_u5_u5_n194 ) );
  NAND2_X1 u2_u5_u5_U21 (.A1( u2_u5_u5_n121 ) , .ZN( u2_u5_u5_n132 ) , .A2( u2_u5_u5_n172 ) );
  NAND2_X1 u2_u5_u5_U22 (.A2( u2_u5_u5_n122 ) , .ZN( u2_u5_u5_n136 ) , .A1( u2_u5_u5_n154 ) );
  NAND2_X1 u2_u5_u5_U23 (.A2( u2_u5_u5_n119 ) , .A1( u2_u5_u5_n120 ) , .ZN( u2_u5_u5_n159 ) );
  INV_X1 u2_u5_u5_U24 (.A( u2_u5_u5_n156 ) , .ZN( u2_u5_u5_n175 ) );
  INV_X1 u2_u5_u5_U25 (.A( u2_u5_u5_n158 ) , .ZN( u2_u5_u5_n188 ) );
  INV_X1 u2_u5_u5_U26 (.A( u2_u5_u5_n152 ) , .ZN( u2_u5_u5_n179 ) );
  INV_X1 u2_u5_u5_U27 (.A( u2_u5_u5_n140 ) , .ZN( u2_u5_u5_n182 ) );
  INV_X1 u2_u5_u5_U28 (.A( u2_u5_u5_n151 ) , .ZN( u2_u5_u5_n183 ) );
  INV_X1 u2_u5_u5_U29 (.A( u2_u5_u5_n123 ) , .ZN( u2_u5_u5_n185 ) );
  NOR2_X1 u2_u5_u5_U3 (.ZN( u2_u5_u5_n134 ) , .A1( u2_u5_u5_n183 ) , .A2( u2_u5_u5_n190 ) );
  INV_X1 u2_u5_u5_U30 (.A( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n184 ) );
  INV_X1 u2_u5_u5_U31 (.A( u2_u5_u5_n139 ) , .ZN( u2_u5_u5_n189 ) );
  INV_X1 u2_u5_u5_U32 (.A( u2_u5_u5_n157 ) , .ZN( u2_u5_u5_n190 ) );
  INV_X1 u2_u5_u5_U33 (.A( u2_u5_u5_n120 ) , .ZN( u2_u5_u5_n193 ) );
  NAND2_X1 u2_u5_u5_U34 (.ZN( u2_u5_u5_n111 ) , .A1( u2_u5_u5_n140 ) , .A2( u2_u5_u5_n155 ) );
  NOR2_X1 u2_u5_u5_U35 (.ZN( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n170 ) , .A2( u2_u5_u5_n180 ) );
  INV_X1 u2_u5_u5_U36 (.A( u2_u5_u5_n117 ) , .ZN( u2_u5_u5_n196 ) );
  OAI221_X1 u2_u5_u5_U37 (.A( u2_u5_u5_n116 ) , .ZN( u2_u5_u5_n117 ) , .B2( u2_u5_u5_n119 ) , .C1( u2_u5_u5_n153 ) , .C2( u2_u5_u5_n158 ) , .B1( u2_u5_u5_n172 ) );
  AOI222_X1 u2_u5_u5_U38 (.ZN( u2_u5_u5_n116 ) , .B2( u2_u5_u5_n145 ) , .C1( u2_u5_u5_n148 ) , .A2( u2_u5_u5_n174 ) , .C2( u2_u5_u5_n177 ) , .B1( u2_u5_u5_n187 ) , .A1( u2_u5_u5_n193 ) );
  INV_X1 u2_u5_u5_U39 (.A( u2_u5_u5_n115 ) , .ZN( u2_u5_u5_n187 ) );
  INV_X1 u2_u5_u5_U4 (.A( u2_u5_u5_n138 ) , .ZN( u2_u5_u5_n191 ) );
  AOI22_X1 u2_u5_u5_U40 (.B2( u2_u5_u5_n131 ) , .A2( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n169 ) , .B1( u2_u5_u5_n174 ) , .A1( u2_u5_u5_n185 ) );
  NOR2_X1 u2_u5_u5_U41 (.A1( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n150 ) , .A2( u2_u5_u5_n173 ) );
  AOI21_X1 u2_u5_u5_U42 (.A( u2_u5_u5_n118 ) , .B2( u2_u5_u5_n145 ) , .ZN( u2_u5_u5_n168 ) , .B1( u2_u5_u5_n186 ) );
  INV_X1 u2_u5_u5_U43 (.A( u2_u5_u5_n122 ) , .ZN( u2_u5_u5_n186 ) );
  NOR2_X1 u2_u5_u5_U44 (.A1( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n152 ) , .A2( u2_u5_u5_n176 ) );
  NOR2_X1 u2_u5_u5_U45 (.A1( u2_u5_u5_n115 ) , .ZN( u2_u5_u5_n118 ) , .A2( u2_u5_u5_n153 ) );
  NOR2_X1 u2_u5_u5_U46 (.A2( u2_u5_u5_n145 ) , .ZN( u2_u5_u5_n156 ) , .A1( u2_u5_u5_n174 ) );
  NOR2_X1 u2_u5_u5_U47 (.ZN( u2_u5_u5_n121 ) , .A2( u2_u5_u5_n145 ) , .A1( u2_u5_u5_n176 ) );
  AOI22_X1 u2_u5_u5_U48 (.ZN( u2_u5_u5_n114 ) , .A2( u2_u5_u5_n137 ) , .A1( u2_u5_u5_n145 ) , .B2( u2_u5_u5_n175 ) , .B1( u2_u5_u5_n193 ) );
  OAI211_X1 u2_u5_u5_U49 (.B( u2_u5_u5_n124 ) , .A( u2_u5_u5_n125 ) , .C2( u2_u5_u5_n126 ) , .C1( u2_u5_u5_n127 ) , .ZN( u2_u5_u5_n128 ) );
  OAI21_X1 u2_u5_u5_U5 (.B2( u2_u5_u5_n136 ) , .B1( u2_u5_u5_n137 ) , .ZN( u2_u5_u5_n138 ) , .A( u2_u5_u5_n177 ) );
  NOR3_X1 u2_u5_u5_U50 (.ZN( u2_u5_u5_n127 ) , .A1( u2_u5_u5_n136 ) , .A3( u2_u5_u5_n148 ) , .A2( u2_u5_u5_n182 ) );
  OAI21_X1 u2_u5_u5_U51 (.ZN( u2_u5_u5_n124 ) , .A( u2_u5_u5_n177 ) , .B2( u2_u5_u5_n183 ) , .B1( u2_u5_u5_n189 ) );
  OAI21_X1 u2_u5_u5_U52 (.ZN( u2_u5_u5_n125 ) , .A( u2_u5_u5_n174 ) , .B2( u2_u5_u5_n185 ) , .B1( u2_u5_u5_n190 ) );
  AOI21_X1 u2_u5_u5_U53 (.A( u2_u5_u5_n153 ) , .B2( u2_u5_u5_n154 ) , .B1( u2_u5_u5_n155 ) , .ZN( u2_u5_u5_n164 ) );
  AOI21_X1 u2_u5_u5_U54 (.ZN( u2_u5_u5_n110 ) , .B1( u2_u5_u5_n122 ) , .B2( u2_u5_u5_n139 ) , .A( u2_u5_u5_n153 ) );
  INV_X1 u2_u5_u5_U55 (.A( u2_u5_u5_n153 ) , .ZN( u2_u5_u5_n176 ) );
  INV_X1 u2_u5_u5_U56 (.A( u2_u5_u5_n126 ) , .ZN( u2_u5_u5_n173 ) );
  AND2_X1 u2_u5_u5_U57 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n147 ) );
  AND2_X1 u2_u5_u5_U58 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n148 ) );
  NAND2_X1 u2_u5_u5_U59 (.A1( u2_u5_u5_n105 ) , .A2( u2_u5_u5_n106 ) , .ZN( u2_u5_u5_n158 ) );
  INV_X1 u2_u5_u5_U6 (.A( u2_u5_u5_n135 ) , .ZN( u2_u5_u5_n178 ) );
  NAND2_X1 u2_u5_u5_U60 (.A2( u2_u5_u5_n108 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n139 ) );
  NAND2_X1 u2_u5_u5_U61 (.A1( u2_u5_u5_n106 ) , .A2( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n119 ) );
  NAND2_X1 u2_u5_u5_U62 (.A2( u2_u5_u5_n103 ) , .A1( u2_u5_u5_n105 ) , .ZN( u2_u5_u5_n140 ) );
  NAND2_X1 u2_u5_u5_U63 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n105 ) , .ZN( u2_u5_u5_n155 ) );
  NAND2_X1 u2_u5_u5_U64 (.A2( u2_u5_u5_n106 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n122 ) );
  NAND2_X1 u2_u5_u5_U65 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n106 ) , .ZN( u2_u5_u5_n115 ) );
  NAND2_X1 u2_u5_u5_U66 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n103 ) , .ZN( u2_u5_u5_n161 ) );
  NAND2_X1 u2_u5_u5_U67 (.A1( u2_u5_u5_n105 ) , .A2( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n154 ) );
  INV_X1 u2_u5_u5_U68 (.A( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n172 ) );
  NAND2_X1 u2_u5_u5_U69 (.A1( u2_u5_u5_n103 ) , .A2( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n123 ) );
  OAI22_X1 u2_u5_u5_U7 (.B2( u2_u5_u5_n149 ) , .B1( u2_u5_u5_n150 ) , .A2( u2_u5_u5_n151 ) , .A1( u2_u5_u5_n152 ) , .ZN( u2_u5_u5_n165 ) );
  NAND2_X1 u2_u5_u5_U70 (.A2( u2_u5_u5_n103 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n151 ) );
  NAND2_X1 u2_u5_u5_U71 (.A2( u2_u5_u5_n107 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n120 ) );
  NAND2_X1 u2_u5_u5_U72 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n157 ) );
  AND2_X1 u2_u5_u5_U73 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n104 ) , .ZN( u2_u5_u5_n131 ) );
  INV_X1 u2_u5_u5_U74 (.A( u2_u5_u5_n102 ) , .ZN( u2_u5_u5_n195 ) );
  OAI221_X1 u2_u5_u5_U75 (.A( u2_u5_u5_n101 ) , .ZN( u2_u5_u5_n102 ) , .C2( u2_u5_u5_n115 ) , .C1( u2_u5_u5_n126 ) , .B1( u2_u5_u5_n134 ) , .B2( u2_u5_u5_n160 ) );
  OAI21_X1 u2_u5_u5_U76 (.ZN( u2_u5_u5_n101 ) , .B1( u2_u5_u5_n137 ) , .A( u2_u5_u5_n146 ) , .B2( u2_u5_u5_n147 ) );
  NOR2_X1 u2_u5_u5_U77 (.A2( u2_u5_X_34 ) , .A1( u2_u5_X_35 ) , .ZN( u2_u5_u5_n145 ) );
  NOR2_X1 u2_u5_u5_U78 (.A2( u2_u5_X_34 ) , .ZN( u2_u5_u5_n146 ) , .A1( u2_u5_u5_n171 ) );
  NOR2_X1 u2_u5_u5_U79 (.A2( u2_u5_X_31 ) , .A1( u2_u5_X_32 ) , .ZN( u2_u5_u5_n103 ) );
  NOR3_X1 u2_u5_u5_U8 (.A2( u2_u5_u5_n147 ) , .A1( u2_u5_u5_n148 ) , .ZN( u2_u5_u5_n149 ) , .A3( u2_u5_u5_n194 ) );
  NOR2_X1 u2_u5_u5_U80 (.A2( u2_u5_X_36 ) , .ZN( u2_u5_u5_n105 ) , .A1( u2_u5_u5_n180 ) );
  NOR2_X1 u2_u5_u5_U81 (.A2( u2_u5_X_33 ) , .ZN( u2_u5_u5_n108 ) , .A1( u2_u5_u5_n170 ) );
  NOR2_X1 u2_u5_u5_U82 (.A2( u2_u5_X_33 ) , .A1( u2_u5_X_36 ) , .ZN( u2_u5_u5_n107 ) );
  NOR2_X1 u2_u5_u5_U83 (.A2( u2_u5_X_31 ) , .ZN( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n181 ) );
  NAND2_X1 u2_u5_u5_U84 (.A2( u2_u5_X_34 ) , .A1( u2_u5_X_35 ) , .ZN( u2_u5_u5_n153 ) );
  NAND2_X1 u2_u5_u5_U85 (.A1( u2_u5_X_34 ) , .ZN( u2_u5_u5_n126 ) , .A2( u2_u5_u5_n171 ) );
  AND2_X1 u2_u5_u5_U86 (.A1( u2_u5_X_31 ) , .A2( u2_u5_X_32 ) , .ZN( u2_u5_u5_n106 ) );
  AND2_X1 u2_u5_u5_U87 (.A1( u2_u5_X_31 ) , .ZN( u2_u5_u5_n109 ) , .A2( u2_u5_u5_n181 ) );
  INV_X1 u2_u5_u5_U88 (.A( u2_u5_X_33 ) , .ZN( u2_u5_u5_n180 ) );
  INV_X1 u2_u5_u5_U89 (.A( u2_u5_X_35 ) , .ZN( u2_u5_u5_n171 ) );
  NOR2_X1 u2_u5_u5_U9 (.ZN( u2_u5_u5_n135 ) , .A1( u2_u5_u5_n173 ) , .A2( u2_u5_u5_n176 ) );
  INV_X1 u2_u5_u5_U90 (.A( u2_u5_X_36 ) , .ZN( u2_u5_u5_n170 ) );
  INV_X1 u2_u5_u5_U91 (.A( u2_u5_X_32 ) , .ZN( u2_u5_u5_n181 ) );
  NAND4_X1 u2_u5_u5_U92 (.ZN( u2_out5_29 ) , .A4( u2_u5_u5_n129 ) , .A3( u2_u5_u5_n130 ) , .A2( u2_u5_u5_n168 ) , .A1( u2_u5_u5_n196 ) );
  AOI221_X1 u2_u5_u5_U93 (.A( u2_u5_u5_n128 ) , .ZN( u2_u5_u5_n129 ) , .C2( u2_u5_u5_n132 ) , .B2( u2_u5_u5_n159 ) , .B1( u2_u5_u5_n176 ) , .C1( u2_u5_u5_n184 ) );
  AOI222_X1 u2_u5_u5_U94 (.ZN( u2_u5_u5_n130 ) , .A2( u2_u5_u5_n146 ) , .B1( u2_u5_u5_n147 ) , .C2( u2_u5_u5_n175 ) , .B2( u2_u5_u5_n179 ) , .A1( u2_u5_u5_n188 ) , .C1( u2_u5_u5_n194 ) );
  NAND4_X1 u2_u5_u5_U95 (.ZN( u2_out5_19 ) , .A4( u2_u5_u5_n166 ) , .A3( u2_u5_u5_n167 ) , .A2( u2_u5_u5_n168 ) , .A1( u2_u5_u5_n169 ) );
  AOI22_X1 u2_u5_u5_U96 (.B2( u2_u5_u5_n145 ) , .A2( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n167 ) , .B1( u2_u5_u5_n182 ) , .A1( u2_u5_u5_n189 ) );
  NOR4_X1 u2_u5_u5_U97 (.A4( u2_u5_u5_n162 ) , .A3( u2_u5_u5_n163 ) , .A2( u2_u5_u5_n164 ) , .A1( u2_u5_u5_n165 ) , .ZN( u2_u5_u5_n166 ) );
  NAND4_X1 u2_u5_u5_U98 (.ZN( u2_out5_11 ) , .A4( u2_u5_u5_n143 ) , .A3( u2_u5_u5_n144 ) , .A2( u2_u5_u5_n169 ) , .A1( u2_u5_u5_n196 ) );
  AOI22_X1 u2_u5_u5_U99 (.A2( u2_u5_u5_n132 ) , .ZN( u2_u5_u5_n144 ) , .B2( u2_u5_u5_n145 ) , .B1( u2_u5_u5_n184 ) , .A1( u2_u5_u5_n194 ) );
  OAI21_X1 u2_u5_u6_U10 (.A( u2_u5_u6_n159 ) , .B1( u2_u5_u6_n169 ) , .B2( u2_u5_u6_n173 ) , .ZN( u2_u5_u6_n90 ) );
  INV_X1 u2_u5_u6_U11 (.ZN( u2_u5_u6_n172 ) , .A( u2_u5_u6_n88 ) );
  AOI22_X1 u2_u5_u6_U12 (.A2( u2_u5_u6_n151 ) , .B2( u2_u5_u6_n161 ) , .A1( u2_u5_u6_n167 ) , .B1( u2_u5_u6_n170 ) , .ZN( u2_u5_u6_n89 ) );
  AOI21_X1 u2_u5_u6_U13 (.ZN( u2_u5_u6_n106 ) , .A( u2_u5_u6_n142 ) , .B2( u2_u5_u6_n159 ) , .B1( u2_u5_u6_n164 ) );
  INV_X1 u2_u5_u6_U14 (.A( u2_u5_u6_n155 ) , .ZN( u2_u5_u6_n161 ) );
  INV_X1 u2_u5_u6_U15 (.A( u2_u5_u6_n128 ) , .ZN( u2_u5_u6_n164 ) );
  NAND2_X1 u2_u5_u6_U16 (.ZN( u2_u5_u6_n110 ) , .A1( u2_u5_u6_n122 ) , .A2( u2_u5_u6_n129 ) );
  NAND2_X1 u2_u5_u6_U17 (.ZN( u2_u5_u6_n124 ) , .A2( u2_u5_u6_n146 ) , .A1( u2_u5_u6_n148 ) );
  INV_X1 u2_u5_u6_U18 (.A( u2_u5_u6_n132 ) , .ZN( u2_u5_u6_n171 ) );
  AND2_X1 u2_u5_u6_U19 (.A1( u2_u5_u6_n100 ) , .ZN( u2_u5_u6_n130 ) , .A2( u2_u5_u6_n147 ) );
  INV_X1 u2_u5_u6_U20 (.A( u2_u5_u6_n127 ) , .ZN( u2_u5_u6_n173 ) );
  INV_X1 u2_u5_u6_U21 (.A( u2_u5_u6_n121 ) , .ZN( u2_u5_u6_n167 ) );
  INV_X1 u2_u5_u6_U22 (.A( u2_u5_u6_n100 ) , .ZN( u2_u5_u6_n169 ) );
  INV_X1 u2_u5_u6_U23 (.A( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n170 ) );
  INV_X1 u2_u5_u6_U24 (.A( u2_u5_u6_n113 ) , .ZN( u2_u5_u6_n168 ) );
  AND2_X1 u2_u5_u6_U25 (.A1( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n119 ) , .ZN( u2_u5_u6_n133 ) );
  AND2_X1 u2_u5_u6_U26 (.A2( u2_u5_u6_n121 ) , .A1( u2_u5_u6_n122 ) , .ZN( u2_u5_u6_n131 ) );
  AND3_X1 u2_u5_u6_U27 (.ZN( u2_u5_u6_n120 ) , .A2( u2_u5_u6_n127 ) , .A1( u2_u5_u6_n132 ) , .A3( u2_u5_u6_n145 ) );
  INV_X1 u2_u5_u6_U28 (.A( u2_u5_u6_n146 ) , .ZN( u2_u5_u6_n163 ) );
  AOI222_X1 u2_u5_u6_U29 (.ZN( u2_u5_u6_n114 ) , .A1( u2_u5_u6_n118 ) , .A2( u2_u5_u6_n126 ) , .B2( u2_u5_u6_n151 ) , .C2( u2_u5_u6_n159 ) , .C1( u2_u5_u6_n168 ) , .B1( u2_u5_u6_n169 ) );
  INV_X1 u2_u5_u6_U3 (.A( u2_u5_u6_n110 ) , .ZN( u2_u5_u6_n166 ) );
  NOR2_X1 u2_u5_u6_U30 (.A1( u2_u5_u6_n162 ) , .A2( u2_u5_u6_n165 ) , .ZN( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U31 (.A1( u2_u5_u6_n144 ) , .ZN( u2_u5_u6_n151 ) , .A2( u2_u5_u6_n158 ) );
  NAND2_X1 u2_u5_u6_U32 (.ZN( u2_u5_u6_n132 ) , .A1( u2_u5_u6_n91 ) , .A2( u2_u5_u6_n97 ) );
  NOR2_X1 u2_u5_u6_U33 (.A2( u2_u5_u6_n126 ) , .ZN( u2_u5_u6_n155 ) , .A1( u2_u5_u6_n160 ) );
  NAND2_X1 u2_u5_u6_U34 (.ZN( u2_u5_u6_n146 ) , .A2( u2_u5_u6_n94 ) , .A1( u2_u5_u6_n99 ) );
  AOI21_X1 u2_u5_u6_U35 (.A( u2_u5_u6_n144 ) , .B2( u2_u5_u6_n145 ) , .B1( u2_u5_u6_n146 ) , .ZN( u2_u5_u6_n150 ) );
  INV_X1 u2_u5_u6_U36 (.A( u2_u5_u6_n111 ) , .ZN( u2_u5_u6_n158 ) );
  NAND2_X1 u2_u5_u6_U37 (.ZN( u2_u5_u6_n127 ) , .A1( u2_u5_u6_n91 ) , .A2( u2_u5_u6_n92 ) );
  NAND2_X1 u2_u5_u6_U38 (.ZN( u2_u5_u6_n129 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n96 ) );
  INV_X1 u2_u5_u6_U39 (.A( u2_u5_u6_n144 ) , .ZN( u2_u5_u6_n159 ) );
  INV_X1 u2_u5_u6_U4 (.A( u2_u5_u6_n142 ) , .ZN( u2_u5_u6_n174 ) );
  NAND2_X1 u2_u5_u6_U40 (.ZN( u2_u5_u6_n145 ) , .A2( u2_u5_u6_n97 ) , .A1( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U41 (.ZN( u2_u5_u6_n148 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n94 ) );
  NAND2_X1 u2_u5_u6_U42 (.ZN( u2_u5_u6_n108 ) , .A2( u2_u5_u6_n139 ) , .A1( u2_u5_u6_n144 ) );
  NAND2_X1 u2_u5_u6_U43 (.ZN( u2_u5_u6_n121 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n97 ) );
  NAND2_X1 u2_u5_u6_U44 (.ZN( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n95 ) );
  AND2_X1 u2_u5_u6_U45 (.ZN( u2_u5_u6_n118 ) , .A2( u2_u5_u6_n91 ) , .A1( u2_u5_u6_n99 ) );
  AOI22_X1 u2_u5_u6_U46 (.B2( u2_u5_u6_n110 ) , .B1( u2_u5_u6_n111 ) , .A1( u2_u5_u6_n112 ) , .ZN( u2_u5_u6_n115 ) , .A2( u2_u5_u6_n161 ) );
  NAND4_X1 u2_u5_u6_U47 (.A3( u2_u5_u6_n109 ) , .ZN( u2_u5_u6_n112 ) , .A4( u2_u5_u6_n132 ) , .A2( u2_u5_u6_n147 ) , .A1( u2_u5_u6_n166 ) );
  NOR2_X1 u2_u5_u6_U48 (.ZN( u2_u5_u6_n109 ) , .A1( u2_u5_u6_n170 ) , .A2( u2_u5_u6_n173 ) );
  NAND2_X1 u2_u5_u6_U49 (.ZN( u2_u5_u6_n147 ) , .A2( u2_u5_u6_n98 ) , .A1( u2_u5_u6_n99 ) );
  NAND2_X1 u2_u5_u6_U5 (.A2( u2_u5_u6_n143 ) , .ZN( u2_u5_u6_n152 ) , .A1( u2_u5_u6_n166 ) );
  NAND2_X1 u2_u5_u6_U50 (.ZN( u2_u5_u6_n128 ) , .A1( u2_u5_u6_n94 ) , .A2( u2_u5_u6_n96 ) );
  AOI211_X1 u2_u5_u6_U51 (.B( u2_u5_u6_n134 ) , .A( u2_u5_u6_n135 ) , .C1( u2_u5_u6_n136 ) , .ZN( u2_u5_u6_n137 ) , .C2( u2_u5_u6_n151 ) );
  AOI21_X1 u2_u5_u6_U52 (.B2( u2_u5_u6_n132 ) , .B1( u2_u5_u6_n133 ) , .ZN( u2_u5_u6_n134 ) , .A( u2_u5_u6_n158 ) );
  AOI21_X1 u2_u5_u6_U53 (.B1( u2_u5_u6_n131 ) , .ZN( u2_u5_u6_n135 ) , .A( u2_u5_u6_n144 ) , .B2( u2_u5_u6_n146 ) );
  NAND4_X1 u2_u5_u6_U54 (.A4( u2_u5_u6_n127 ) , .A3( u2_u5_u6_n128 ) , .A2( u2_u5_u6_n129 ) , .A1( u2_u5_u6_n130 ) , .ZN( u2_u5_u6_n136 ) );
  NAND2_X1 u2_u5_u6_U55 (.ZN( u2_u5_u6_n119 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n99 ) );
  NAND2_X1 u2_u5_u6_U56 (.ZN( u2_u5_u6_n123 ) , .A2( u2_u5_u6_n91 ) , .A1( u2_u5_u6_n96 ) );
  NAND2_X1 u2_u5_u6_U57 (.ZN( u2_u5_u6_n100 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U58 (.ZN( u2_u5_u6_n122 ) , .A1( u2_u5_u6_n94 ) , .A2( u2_u5_u6_n97 ) );
  INV_X1 u2_u5_u6_U59 (.A( u2_u5_u6_n139 ) , .ZN( u2_u5_u6_n160 ) );
  AOI22_X1 u2_u5_u6_U6 (.B2( u2_u5_u6_n101 ) , .A1( u2_u5_u6_n102 ) , .ZN( u2_u5_u6_n103 ) , .B1( u2_u5_u6_n160 ) , .A2( u2_u5_u6_n161 ) );
  NAND2_X1 u2_u5_u6_U60 (.ZN( u2_u5_u6_n113 ) , .A1( u2_u5_u6_n96 ) , .A2( u2_u5_u6_n98 ) );
  NOR2_X1 u2_u5_u6_U61 (.A2( u2_u5_X_40 ) , .A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n126 ) );
  NOR2_X1 u2_u5_u6_U62 (.A2( u2_u5_X_39 ) , .A1( u2_u5_X_42 ) , .ZN( u2_u5_u6_n92 ) );
  NOR2_X1 u2_u5_u6_U63 (.A2( u2_u5_X_39 ) , .A1( u2_u5_u6_n156 ) , .ZN( u2_u5_u6_n97 ) );
  NOR2_X1 u2_u5_u6_U64 (.A2( u2_u5_X_38 ) , .A1( u2_u5_u6_n165 ) , .ZN( u2_u5_u6_n95 ) );
  NOR2_X1 u2_u5_u6_U65 (.A2( u2_u5_X_41 ) , .ZN( u2_u5_u6_n111 ) , .A1( u2_u5_u6_n157 ) );
  NOR2_X1 u2_u5_u6_U66 (.A2( u2_u5_X_37 ) , .A1( u2_u5_u6_n162 ) , .ZN( u2_u5_u6_n94 ) );
  NOR2_X1 u2_u5_u6_U67 (.A2( u2_u5_X_37 ) , .A1( u2_u5_X_38 ) , .ZN( u2_u5_u6_n91 ) );
  NAND2_X1 u2_u5_u6_U68 (.A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n144 ) , .A2( u2_u5_u6_n157 ) );
  NAND2_X1 u2_u5_u6_U69 (.A2( u2_u5_X_40 ) , .A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n139 ) );
  NOR2_X1 u2_u5_u6_U7 (.A1( u2_u5_u6_n118 ) , .ZN( u2_u5_u6_n143 ) , .A2( u2_u5_u6_n168 ) );
  AND2_X1 u2_u5_u6_U70 (.A1( u2_u5_X_39 ) , .A2( u2_u5_u6_n156 ) , .ZN( u2_u5_u6_n96 ) );
  AND2_X1 u2_u5_u6_U71 (.A1( u2_u5_X_39 ) , .A2( u2_u5_X_42 ) , .ZN( u2_u5_u6_n99 ) );
  INV_X1 u2_u5_u6_U72 (.A( u2_u5_X_40 ) , .ZN( u2_u5_u6_n157 ) );
  INV_X1 u2_u5_u6_U73 (.A( u2_u5_X_37 ) , .ZN( u2_u5_u6_n165 ) );
  INV_X1 u2_u5_u6_U74 (.A( u2_u5_X_38 ) , .ZN( u2_u5_u6_n162 ) );
  INV_X1 u2_u5_u6_U75 (.A( u2_u5_X_42 ) , .ZN( u2_u5_u6_n156 ) );
  NAND4_X1 u2_u5_u6_U76 (.ZN( u2_out5_32 ) , .A4( u2_u5_u6_n103 ) , .A3( u2_u5_u6_n104 ) , .A2( u2_u5_u6_n105 ) , .A1( u2_u5_u6_n106 ) );
  AOI22_X1 u2_u5_u6_U77 (.ZN( u2_u5_u6_n105 ) , .A2( u2_u5_u6_n108 ) , .A1( u2_u5_u6_n118 ) , .B2( u2_u5_u6_n126 ) , .B1( u2_u5_u6_n171 ) );
  AOI22_X1 u2_u5_u6_U78 (.ZN( u2_u5_u6_n104 ) , .A1( u2_u5_u6_n111 ) , .B1( u2_u5_u6_n124 ) , .B2( u2_u5_u6_n151 ) , .A2( u2_u5_u6_n93 ) );
  NAND4_X1 u2_u5_u6_U79 (.ZN( u2_out5_12 ) , .A4( u2_u5_u6_n114 ) , .A3( u2_u5_u6_n115 ) , .A2( u2_u5_u6_n116 ) , .A1( u2_u5_u6_n117 ) );
  AOI21_X1 u2_u5_u6_U8 (.B1( u2_u5_u6_n107 ) , .B2( u2_u5_u6_n132 ) , .A( u2_u5_u6_n158 ) , .ZN( u2_u5_u6_n88 ) );
  OAI22_X1 u2_u5_u6_U80 (.B2( u2_u5_u6_n111 ) , .ZN( u2_u5_u6_n116 ) , .B1( u2_u5_u6_n126 ) , .A2( u2_u5_u6_n164 ) , .A1( u2_u5_u6_n167 ) );
  OAI21_X1 u2_u5_u6_U81 (.A( u2_u5_u6_n108 ) , .ZN( u2_u5_u6_n117 ) , .B2( u2_u5_u6_n141 ) , .B1( u2_u5_u6_n163 ) );
  OAI211_X1 u2_u5_u6_U82 (.ZN( u2_out5_22 ) , .B( u2_u5_u6_n137 ) , .A( u2_u5_u6_n138 ) , .C2( u2_u5_u6_n139 ) , .C1( u2_u5_u6_n140 ) );
  AOI22_X1 u2_u5_u6_U83 (.B1( u2_u5_u6_n124 ) , .A2( u2_u5_u6_n125 ) , .A1( u2_u5_u6_n126 ) , .ZN( u2_u5_u6_n138 ) , .B2( u2_u5_u6_n161 ) );
  AND4_X1 u2_u5_u6_U84 (.A3( u2_u5_u6_n119 ) , .A1( u2_u5_u6_n120 ) , .A4( u2_u5_u6_n129 ) , .ZN( u2_u5_u6_n140 ) , .A2( u2_u5_u6_n143 ) );
  OAI211_X1 u2_u5_u6_U85 (.ZN( u2_out5_7 ) , .B( u2_u5_u6_n153 ) , .C2( u2_u5_u6_n154 ) , .C1( u2_u5_u6_n155 ) , .A( u2_u5_u6_n174 ) );
  NOR3_X1 u2_u5_u6_U86 (.A1( u2_u5_u6_n141 ) , .ZN( u2_u5_u6_n154 ) , .A3( u2_u5_u6_n164 ) , .A2( u2_u5_u6_n171 ) );
  AOI211_X1 u2_u5_u6_U87 (.B( u2_u5_u6_n149 ) , .A( u2_u5_u6_n150 ) , .C2( u2_u5_u6_n151 ) , .C1( u2_u5_u6_n152 ) , .ZN( u2_u5_u6_n153 ) );
  NAND3_X1 u2_u5_u6_U88 (.A2( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n125 ) , .A1( u2_u5_u6_n130 ) , .A3( u2_u5_u6_n131 ) );
  NAND3_X1 u2_u5_u6_U89 (.A3( u2_u5_u6_n133 ) , .ZN( u2_u5_u6_n141 ) , .A1( u2_u5_u6_n145 ) , .A2( u2_u5_u6_n148 ) );
  AOI21_X1 u2_u5_u6_U9 (.B2( u2_u5_u6_n147 ) , .B1( u2_u5_u6_n148 ) , .ZN( u2_u5_u6_n149 ) , .A( u2_u5_u6_n158 ) );
  NAND3_X1 u2_u5_u6_U90 (.ZN( u2_u5_u6_n101 ) , .A3( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n121 ) , .A1( u2_u5_u6_n127 ) );
  NAND3_X1 u2_u5_u6_U91 (.ZN( u2_u5_u6_n102 ) , .A3( u2_u5_u6_n130 ) , .A2( u2_u5_u6_n145 ) , .A1( u2_u5_u6_n166 ) );
  NAND3_X1 u2_u5_u6_U92 (.A3( u2_u5_u6_n113 ) , .A1( u2_u5_u6_n119 ) , .A2( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n93 ) );
  NAND3_X1 u2_u5_u6_U93 (.ZN( u2_u5_u6_n142 ) , .A2( u2_u5_u6_n172 ) , .A3( u2_u5_u6_n89 ) , .A1( u2_u5_u6_n90 ) );
  XOR2_X1 u2_u6_U1 (.B( u2_K7_9 ) , .A( u2_R5_6 ) , .Z( u2_u6_X_9 ) );
  XOR2_X1 u2_u6_U16 (.B( u2_K7_3 ) , .A( u2_R5_2 ) , .Z( u2_u6_X_3 ) );
  XOR2_X1 u2_u6_U2 (.B( u2_K7_8 ) , .A( u2_R5_5 ) , .Z( u2_u6_X_8 ) );
  XOR2_X1 u2_u6_U27 (.B( u2_K7_2 ) , .A( u2_R5_1 ) , .Z( u2_u6_X_2 ) );
  XOR2_X1 u2_u6_U3 (.B( u2_K7_7 ) , .A( u2_R5_4 ) , .Z( u2_u6_X_7 ) );
  XOR2_X1 u2_u6_U38 (.B( u2_K7_1 ) , .A( u2_R5_32 ) , .Z( u2_u6_X_1 ) );
  XOR2_X1 u2_u6_U4 (.B( u2_K7_6 ) , .A( u2_R5_5 ) , .Z( u2_u6_X_6 ) );
  XOR2_X1 u2_u6_U40 (.B( u2_K7_18 ) , .A( u2_R5_13 ) , .Z( u2_u6_X_18 ) );
  XOR2_X1 u2_u6_U41 (.B( u2_K7_17 ) , .A( u2_R5_12 ) , .Z( u2_u6_X_17 ) );
  XOR2_X1 u2_u6_U42 (.B( u2_K7_16 ) , .A( u2_R5_11 ) , .Z( u2_u6_X_16 ) );
  XOR2_X1 u2_u6_U43 (.B( u2_K7_15 ) , .A( u2_R5_10 ) , .Z( u2_u6_X_15 ) );
  XOR2_X1 u2_u6_U44 (.B( u2_K7_14 ) , .A( u2_R5_9 ) , .Z( u2_u6_X_14 ) );
  XOR2_X1 u2_u6_U45 (.B( u2_K7_13 ) , .A( u2_R5_8 ) , .Z( u2_u6_X_13 ) );
  XOR2_X1 u2_u6_U46 (.B( u2_K7_12 ) , .A( u2_R5_9 ) , .Z( u2_u6_X_12 ) );
  XOR2_X1 u2_u6_U47 (.B( u2_K7_11 ) , .A( u2_R5_8 ) , .Z( u2_u6_X_11 ) );
  XOR2_X1 u2_u6_U48 (.B( u2_K7_10 ) , .A( u2_R5_7 ) , .Z( u2_u6_X_10 ) );
  XOR2_X1 u2_u6_U5 (.B( u2_K7_5 ) , .A( u2_R5_4 ) , .Z( u2_u6_X_5 ) );
  XOR2_X1 u2_u6_U6 (.B( u2_K7_4 ) , .A( u2_R5_3 ) , .Z( u2_u6_X_4 ) );
  AND3_X1 u2_u6_u0_U10 (.A2( u2_u6_u0_n112 ) , .ZN( u2_u6_u0_n127 ) , .A3( u2_u6_u0_n130 ) , .A1( u2_u6_u0_n148 ) );
  NAND2_X1 u2_u6_u0_U11 (.ZN( u2_u6_u0_n113 ) , .A1( u2_u6_u0_n139 ) , .A2( u2_u6_u0_n149 ) );
  AND2_X1 u2_u6_u0_U12 (.ZN( u2_u6_u0_n107 ) , .A1( u2_u6_u0_n130 ) , .A2( u2_u6_u0_n140 ) );
  AND2_X1 u2_u6_u0_U13 (.A2( u2_u6_u0_n129 ) , .A1( u2_u6_u0_n130 ) , .ZN( u2_u6_u0_n151 ) );
  AND2_X1 u2_u6_u0_U14 (.A1( u2_u6_u0_n108 ) , .A2( u2_u6_u0_n125 ) , .ZN( u2_u6_u0_n145 ) );
  INV_X1 u2_u6_u0_U15 (.A( u2_u6_u0_n143 ) , .ZN( u2_u6_u0_n173 ) );
  NOR2_X1 u2_u6_u0_U16 (.A2( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n147 ) , .A1( u2_u6_u0_n160 ) );
  NOR2_X1 u2_u6_u0_U17 (.A1( u2_u6_u0_n163 ) , .A2( u2_u6_u0_n164 ) , .ZN( u2_u6_u0_n95 ) );
  AOI21_X1 u2_u6_u0_U18 (.B1( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n132 ) , .A( u2_u6_u0_n165 ) , .B2( u2_u6_u0_n93 ) );
  INV_X1 u2_u6_u0_U19 (.A( u2_u6_u0_n142 ) , .ZN( u2_u6_u0_n165 ) );
  OAI22_X1 u2_u6_u0_U20 (.B1( u2_u6_u0_n125 ) , .ZN( u2_u6_u0_n126 ) , .A1( u2_u6_u0_n138 ) , .A2( u2_u6_u0_n146 ) , .B2( u2_u6_u0_n147 ) );
  OAI22_X1 u2_u6_u0_U21 (.B1( u2_u6_u0_n131 ) , .A1( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n147 ) , .A2( u2_u6_u0_n90 ) , .ZN( u2_u6_u0_n91 ) );
  AND3_X1 u2_u6_u0_U22 (.A3( u2_u6_u0_n121 ) , .A2( u2_u6_u0_n125 ) , .A1( u2_u6_u0_n148 ) , .ZN( u2_u6_u0_n90 ) );
  NAND2_X1 u2_u6_u0_U23 (.A1( u2_u6_u0_n100 ) , .A2( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n125 ) );
  INV_X1 u2_u6_u0_U24 (.A( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n161 ) );
  AOI22_X1 u2_u6_u0_U25 (.B2( u2_u6_u0_n109 ) , .A2( u2_u6_u0_n110 ) , .ZN( u2_u6_u0_n111 ) , .B1( u2_u6_u0_n118 ) , .A1( u2_u6_u0_n160 ) );
  NAND2_X1 u2_u6_u0_U26 (.A1( u2_u6_u0_n100 ) , .ZN( u2_u6_u0_n129 ) , .A2( u2_u6_u0_n95 ) );
  INV_X1 u2_u6_u0_U27 (.A( u2_u6_u0_n118 ) , .ZN( u2_u6_u0_n158 ) );
  AOI21_X1 u2_u6_u0_U28 (.ZN( u2_u6_u0_n104 ) , .B1( u2_u6_u0_n107 ) , .B2( u2_u6_u0_n141 ) , .A( u2_u6_u0_n144 ) );
  AOI21_X1 u2_u6_u0_U29 (.B1( u2_u6_u0_n127 ) , .B2( u2_u6_u0_n129 ) , .A( u2_u6_u0_n138 ) , .ZN( u2_u6_u0_n96 ) );
  INV_X1 u2_u6_u0_U3 (.A( u2_u6_u0_n113 ) , .ZN( u2_u6_u0_n166 ) );
  AOI21_X1 u2_u6_u0_U30 (.ZN( u2_u6_u0_n116 ) , .B2( u2_u6_u0_n142 ) , .A( u2_u6_u0_n144 ) , .B1( u2_u6_u0_n166 ) );
  NOR2_X1 u2_u6_u0_U31 (.A1( u2_u6_u0_n120 ) , .ZN( u2_u6_u0_n143 ) , .A2( u2_u6_u0_n167 ) );
  OAI221_X1 u2_u6_u0_U32 (.C1( u2_u6_u0_n112 ) , .ZN( u2_u6_u0_n120 ) , .B1( u2_u6_u0_n138 ) , .B2( u2_u6_u0_n141 ) , .C2( u2_u6_u0_n147 ) , .A( u2_u6_u0_n172 ) );
  AOI211_X1 u2_u6_u0_U33 (.B( u2_u6_u0_n115 ) , .A( u2_u6_u0_n116 ) , .C2( u2_u6_u0_n117 ) , .C1( u2_u6_u0_n118 ) , .ZN( u2_u6_u0_n119 ) );
  NAND2_X1 u2_u6_u0_U34 (.A2( u2_u6_u0_n100 ) , .A1( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n139 ) );
  NAND2_X1 u2_u6_u0_U35 (.A2( u2_u6_u0_n100 ) , .ZN( u2_u6_u0_n131 ) , .A1( u2_u6_u0_n92 ) );
  NAND2_X1 u2_u6_u0_U36 (.A1( u2_u6_u0_n101 ) , .A2( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n150 ) );
  INV_X1 u2_u6_u0_U37 (.A( u2_u6_u0_n138 ) , .ZN( u2_u6_u0_n160 ) );
  NAND2_X1 u2_u6_u0_U38 (.A1( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n128 ) , .A2( u2_u6_u0_n95 ) );
  NAND2_X1 u2_u6_u0_U39 (.ZN( u2_u6_u0_n148 ) , .A1( u2_u6_u0_n93 ) , .A2( u2_u6_u0_n95 ) );
  AOI21_X1 u2_u6_u0_U4 (.B1( u2_u6_u0_n114 ) , .ZN( u2_u6_u0_n115 ) , .B2( u2_u6_u0_n129 ) , .A( u2_u6_u0_n161 ) );
  NAND2_X1 u2_u6_u0_U40 (.A2( u2_u6_u0_n102 ) , .A1( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n149 ) );
  NAND2_X1 u2_u6_u0_U41 (.A2( u2_u6_u0_n102 ) , .ZN( u2_u6_u0_n114 ) , .A1( u2_u6_u0_n92 ) );
  NAND2_X1 u2_u6_u0_U42 (.A2( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n121 ) , .A1( u2_u6_u0_n93 ) );
  NAND2_X1 u2_u6_u0_U43 (.ZN( u2_u6_u0_n112 ) , .A2( u2_u6_u0_n92 ) , .A1( u2_u6_u0_n93 ) );
  INV_X1 u2_u6_u0_U44 (.ZN( u2_u6_u0_n172 ) , .A( u2_u6_u0_n88 ) );
  OAI222_X1 u2_u6_u0_U45 (.C1( u2_u6_u0_n108 ) , .A1( u2_u6_u0_n125 ) , .B2( u2_u6_u0_n128 ) , .B1( u2_u6_u0_n144 ) , .A2( u2_u6_u0_n158 ) , .C2( u2_u6_u0_n161 ) , .ZN( u2_u6_u0_n88 ) );
  OR3_X1 u2_u6_u0_U46 (.A3( u2_u6_u0_n152 ) , .A2( u2_u6_u0_n153 ) , .A1( u2_u6_u0_n154 ) , .ZN( u2_u6_u0_n155 ) );
  AOI21_X1 u2_u6_u0_U47 (.A( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n145 ) , .B1( u2_u6_u0_n146 ) , .ZN( u2_u6_u0_n154 ) );
  AOI21_X1 u2_u6_u0_U48 (.B2( u2_u6_u0_n150 ) , .B1( u2_u6_u0_n151 ) , .ZN( u2_u6_u0_n152 ) , .A( u2_u6_u0_n158 ) );
  AOI21_X1 u2_u6_u0_U49 (.A( u2_u6_u0_n147 ) , .B2( u2_u6_u0_n148 ) , .B1( u2_u6_u0_n149 ) , .ZN( u2_u6_u0_n153 ) );
  AOI21_X1 u2_u6_u0_U5 (.B2( u2_u6_u0_n131 ) , .ZN( u2_u6_u0_n134 ) , .B1( u2_u6_u0_n151 ) , .A( u2_u6_u0_n158 ) );
  INV_X1 u2_u6_u0_U50 (.ZN( u2_u6_u0_n171 ) , .A( u2_u6_u0_n99 ) );
  OAI211_X1 u2_u6_u0_U51 (.C2( u2_u6_u0_n140 ) , .C1( u2_u6_u0_n161 ) , .A( u2_u6_u0_n169 ) , .B( u2_u6_u0_n98 ) , .ZN( u2_u6_u0_n99 ) );
  INV_X1 u2_u6_u0_U52 (.ZN( u2_u6_u0_n169 ) , .A( u2_u6_u0_n91 ) );
  AOI211_X1 u2_u6_u0_U53 (.C1( u2_u6_u0_n118 ) , .A( u2_u6_u0_n123 ) , .B( u2_u6_u0_n96 ) , .C2( u2_u6_u0_n97 ) , .ZN( u2_u6_u0_n98 ) );
  NOR2_X1 u2_u6_u0_U54 (.A2( u2_u6_X_4 ) , .A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n118 ) );
  NOR2_X1 u2_u6_u0_U55 (.A2( u2_u6_X_2 ) , .ZN( u2_u6_u0_n103 ) , .A1( u2_u6_u0_n164 ) );
  NOR2_X1 u2_u6_u0_U56 (.A2( u2_u6_X_1 ) , .A1( u2_u6_X_2 ) , .ZN( u2_u6_u0_n92 ) );
  NOR2_X1 u2_u6_u0_U57 (.A2( u2_u6_X_1 ) , .ZN( u2_u6_u0_n101 ) , .A1( u2_u6_u0_n163 ) );
  NAND2_X1 u2_u6_u0_U58 (.A2( u2_u6_X_4 ) , .A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n144 ) );
  NOR2_X1 u2_u6_u0_U59 (.A2( u2_u6_X_5 ) , .ZN( u2_u6_u0_n136 ) , .A1( u2_u6_u0_n159 ) );
  NOR2_X1 u2_u6_u0_U6 (.A1( u2_u6_u0_n108 ) , .ZN( u2_u6_u0_n123 ) , .A2( u2_u6_u0_n158 ) );
  NAND2_X1 u2_u6_u0_U60 (.A1( u2_u6_X_5 ) , .ZN( u2_u6_u0_n138 ) , .A2( u2_u6_u0_n159 ) );
  INV_X1 u2_u6_u0_U61 (.A( u2_u6_X_4 ) , .ZN( u2_u6_u0_n159 ) );
  INV_X1 u2_u6_u0_U62 (.A( u2_u6_X_1 ) , .ZN( u2_u6_u0_n164 ) );
  INV_X1 u2_u6_u0_U63 (.A( u2_u6_X_2 ) , .ZN( u2_u6_u0_n163 ) );
  INV_X1 u2_u6_u0_U64 (.A( u2_u6_X_3 ) , .ZN( u2_u6_u0_n162 ) );
  INV_X1 u2_u6_u0_U65 (.A( u2_u6_u0_n126 ) , .ZN( u2_u6_u0_n168 ) );
  AOI211_X1 u2_u6_u0_U66 (.B( u2_u6_u0_n133 ) , .A( u2_u6_u0_n134 ) , .C2( u2_u6_u0_n135 ) , .C1( u2_u6_u0_n136 ) , .ZN( u2_u6_u0_n137 ) );
  OR4_X1 u2_u6_u0_U67 (.ZN( u2_out6_17 ) , .A4( u2_u6_u0_n122 ) , .A2( u2_u6_u0_n123 ) , .A1( u2_u6_u0_n124 ) , .A3( u2_u6_u0_n170 ) );
  AOI21_X1 u2_u6_u0_U68 (.B2( u2_u6_u0_n107 ) , .ZN( u2_u6_u0_n124 ) , .B1( u2_u6_u0_n128 ) , .A( u2_u6_u0_n161 ) );
  INV_X1 u2_u6_u0_U69 (.A( u2_u6_u0_n111 ) , .ZN( u2_u6_u0_n170 ) );
  OAI21_X1 u2_u6_u0_U7 (.B1( u2_u6_u0_n150 ) , .B2( u2_u6_u0_n158 ) , .A( u2_u6_u0_n172 ) , .ZN( u2_u6_u0_n89 ) );
  OR4_X1 u2_u6_u0_U70 (.ZN( u2_out6_31 ) , .A4( u2_u6_u0_n155 ) , .A2( u2_u6_u0_n156 ) , .A1( u2_u6_u0_n157 ) , .A3( u2_u6_u0_n173 ) );
  AOI21_X1 u2_u6_u0_U71 (.A( u2_u6_u0_n138 ) , .B2( u2_u6_u0_n139 ) , .B1( u2_u6_u0_n140 ) , .ZN( u2_u6_u0_n157 ) );
  AOI21_X1 u2_u6_u0_U72 (.B2( u2_u6_u0_n141 ) , .B1( u2_u6_u0_n142 ) , .ZN( u2_u6_u0_n156 ) , .A( u2_u6_u0_n161 ) );
  INV_X1 u2_u6_u0_U73 (.ZN( u2_u6_u0_n174 ) , .A( u2_u6_u0_n89 ) );
  AOI211_X1 u2_u6_u0_U74 (.B( u2_u6_u0_n104 ) , .A( u2_u6_u0_n105 ) , .ZN( u2_u6_u0_n106 ) , .C2( u2_u6_u0_n113 ) , .C1( u2_u6_u0_n160 ) );
  AND2_X1 u2_u6_u0_U75 (.A1( u2_u6_X_6 ) , .A2( u2_u6_u0_n162 ) , .ZN( u2_u6_u0_n93 ) );
  NOR2_X1 u2_u6_u0_U76 (.A2( u2_u6_X_3 ) , .A1( u2_u6_X_6 ) , .ZN( u2_u6_u0_n94 ) );
  NOR2_X1 u2_u6_u0_U77 (.A2( u2_u6_X_6 ) , .ZN( u2_u6_u0_n100 ) , .A1( u2_u6_u0_n162 ) );
  AND2_X1 u2_u6_u0_U78 (.A2( u2_u6_X_3 ) , .A1( u2_u6_X_6 ) , .ZN( u2_u6_u0_n102 ) );
  OAI221_X1 u2_u6_u0_U79 (.C1( u2_u6_u0_n121 ) , .ZN( u2_u6_u0_n122 ) , .B2( u2_u6_u0_n127 ) , .A( u2_u6_u0_n143 ) , .B1( u2_u6_u0_n144 ) , .C2( u2_u6_u0_n147 ) );
  AND2_X1 u2_u6_u0_U8 (.A1( u2_u6_u0_n114 ) , .A2( u2_u6_u0_n121 ) , .ZN( u2_u6_u0_n146 ) );
  AOI21_X1 u2_u6_u0_U80 (.B1( u2_u6_u0_n132 ) , .ZN( u2_u6_u0_n133 ) , .A( u2_u6_u0_n144 ) , .B2( u2_u6_u0_n166 ) );
  OAI22_X1 u2_u6_u0_U81 (.ZN( u2_u6_u0_n105 ) , .A2( u2_u6_u0_n132 ) , .B1( u2_u6_u0_n146 ) , .A1( u2_u6_u0_n147 ) , .B2( u2_u6_u0_n161 ) );
  NAND2_X1 u2_u6_u0_U82 (.ZN( u2_u6_u0_n110 ) , .A2( u2_u6_u0_n132 ) , .A1( u2_u6_u0_n145 ) );
  INV_X1 u2_u6_u0_U83 (.A( u2_u6_u0_n119 ) , .ZN( u2_u6_u0_n167 ) );
  NAND2_X1 u2_u6_u0_U84 (.A2( u2_u6_u0_n103 ) , .ZN( u2_u6_u0_n140 ) , .A1( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U85 (.A1( u2_u6_u0_n101 ) , .ZN( u2_u6_u0_n130 ) , .A2( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U86 (.ZN( u2_u6_u0_n108 ) , .A1( u2_u6_u0_n92 ) , .A2( u2_u6_u0_n94 ) );
  NAND2_X1 u2_u6_u0_U87 (.ZN( u2_u6_u0_n142 ) , .A1( u2_u6_u0_n94 ) , .A2( u2_u6_u0_n95 ) );
  NAND3_X1 u2_u6_u0_U88 (.ZN( u2_out6_23 ) , .A3( u2_u6_u0_n137 ) , .A1( u2_u6_u0_n168 ) , .A2( u2_u6_u0_n171 ) );
  NAND3_X1 u2_u6_u0_U89 (.A3( u2_u6_u0_n127 ) , .A2( u2_u6_u0_n128 ) , .ZN( u2_u6_u0_n135 ) , .A1( u2_u6_u0_n150 ) );
  AND2_X1 u2_u6_u0_U9 (.A1( u2_u6_u0_n131 ) , .ZN( u2_u6_u0_n141 ) , .A2( u2_u6_u0_n150 ) );
  NAND3_X1 u2_u6_u0_U90 (.ZN( u2_u6_u0_n117 ) , .A3( u2_u6_u0_n132 ) , .A2( u2_u6_u0_n139 ) , .A1( u2_u6_u0_n148 ) );
  NAND3_X1 u2_u6_u0_U91 (.ZN( u2_u6_u0_n109 ) , .A2( u2_u6_u0_n114 ) , .A3( u2_u6_u0_n140 ) , .A1( u2_u6_u0_n149 ) );
  NAND3_X1 u2_u6_u0_U92 (.ZN( u2_out6_9 ) , .A3( u2_u6_u0_n106 ) , .A2( u2_u6_u0_n171 ) , .A1( u2_u6_u0_n174 ) );
  NAND3_X1 u2_u6_u0_U93 (.A2( u2_u6_u0_n128 ) , .A1( u2_u6_u0_n132 ) , .A3( u2_u6_u0_n146 ) , .ZN( u2_u6_u0_n97 ) );
  AOI21_X1 u2_u6_u1_U10 (.B2( u2_u6_u1_n155 ) , .B1( u2_u6_u1_n156 ) , .ZN( u2_u6_u1_n157 ) , .A( u2_u6_u1_n174 ) );
  NAND3_X1 u2_u6_u1_U100 (.ZN( u2_u6_u1_n113 ) , .A1( u2_u6_u1_n120 ) , .A3( u2_u6_u1_n133 ) , .A2( u2_u6_u1_n155 ) );
  NAND2_X1 u2_u6_u1_U11 (.ZN( u2_u6_u1_n140 ) , .A2( u2_u6_u1_n150 ) , .A1( u2_u6_u1_n155 ) );
  NAND2_X1 u2_u6_u1_U12 (.A1( u2_u6_u1_n131 ) , .ZN( u2_u6_u1_n147 ) , .A2( u2_u6_u1_n153 ) );
  INV_X1 u2_u6_u1_U13 (.A( u2_u6_u1_n139 ) , .ZN( u2_u6_u1_n174 ) );
  OR4_X1 u2_u6_u1_U14 (.A4( u2_u6_u1_n106 ) , .A3( u2_u6_u1_n107 ) , .ZN( u2_u6_u1_n108 ) , .A1( u2_u6_u1_n117 ) , .A2( u2_u6_u1_n184 ) );
  AOI21_X1 u2_u6_u1_U15 (.ZN( u2_u6_u1_n106 ) , .A( u2_u6_u1_n112 ) , .B1( u2_u6_u1_n154 ) , .B2( u2_u6_u1_n156 ) );
  AOI21_X1 u2_u6_u1_U16 (.ZN( u2_u6_u1_n107 ) , .B1( u2_u6_u1_n134 ) , .B2( u2_u6_u1_n149 ) , .A( u2_u6_u1_n174 ) );
  INV_X1 u2_u6_u1_U17 (.A( u2_u6_u1_n101 ) , .ZN( u2_u6_u1_n184 ) );
  INV_X1 u2_u6_u1_U18 (.A( u2_u6_u1_n112 ) , .ZN( u2_u6_u1_n171 ) );
  NAND2_X1 u2_u6_u1_U19 (.ZN( u2_u6_u1_n141 ) , .A1( u2_u6_u1_n153 ) , .A2( u2_u6_u1_n156 ) );
  AND2_X1 u2_u6_u1_U20 (.A1( u2_u6_u1_n123 ) , .ZN( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n161 ) );
  NAND2_X1 u2_u6_u1_U21 (.A2( u2_u6_u1_n115 ) , .A1( u2_u6_u1_n116 ) , .ZN( u2_u6_u1_n148 ) );
  NAND2_X1 u2_u6_u1_U22 (.A2( u2_u6_u1_n133 ) , .A1( u2_u6_u1_n135 ) , .ZN( u2_u6_u1_n159 ) );
  NAND2_X1 u2_u6_u1_U23 (.A2( u2_u6_u1_n115 ) , .A1( u2_u6_u1_n120 ) , .ZN( u2_u6_u1_n132 ) );
  INV_X1 u2_u6_u1_U24 (.A( u2_u6_u1_n154 ) , .ZN( u2_u6_u1_n178 ) );
  AOI22_X1 u2_u6_u1_U25 (.B2( u2_u6_u1_n113 ) , .A2( u2_u6_u1_n114 ) , .ZN( u2_u6_u1_n125 ) , .A1( u2_u6_u1_n171 ) , .B1( u2_u6_u1_n173 ) );
  NAND2_X1 u2_u6_u1_U26 (.ZN( u2_u6_u1_n114 ) , .A1( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n156 ) );
  INV_X1 u2_u6_u1_U27 (.A( u2_u6_u1_n151 ) , .ZN( u2_u6_u1_n183 ) );
  AND2_X1 u2_u6_u1_U28 (.A1( u2_u6_u1_n129 ) , .A2( u2_u6_u1_n133 ) , .ZN( u2_u6_u1_n149 ) );
  INV_X1 u2_u6_u1_U29 (.A( u2_u6_u1_n131 ) , .ZN( u2_u6_u1_n180 ) );
  INV_X1 u2_u6_u1_U3 (.A( u2_u6_u1_n159 ) , .ZN( u2_u6_u1_n182 ) );
  AOI221_X1 u2_u6_u1_U30 (.B1( u2_u6_u1_n140 ) , .ZN( u2_u6_u1_n167 ) , .B2( u2_u6_u1_n172 ) , .C2( u2_u6_u1_n175 ) , .C1( u2_u6_u1_n178 ) , .A( u2_u6_u1_n188 ) );
  INV_X1 u2_u6_u1_U31 (.ZN( u2_u6_u1_n188 ) , .A( u2_u6_u1_n97 ) );
  AOI211_X1 u2_u6_u1_U32 (.A( u2_u6_u1_n118 ) , .C1( u2_u6_u1_n132 ) , .C2( u2_u6_u1_n139 ) , .B( u2_u6_u1_n96 ) , .ZN( u2_u6_u1_n97 ) );
  AOI21_X1 u2_u6_u1_U33 (.B2( u2_u6_u1_n121 ) , .B1( u2_u6_u1_n135 ) , .A( u2_u6_u1_n152 ) , .ZN( u2_u6_u1_n96 ) );
  OAI221_X1 u2_u6_u1_U34 (.A( u2_u6_u1_n119 ) , .C2( u2_u6_u1_n129 ) , .ZN( u2_u6_u1_n138 ) , .B2( u2_u6_u1_n152 ) , .C1( u2_u6_u1_n174 ) , .B1( u2_u6_u1_n187 ) );
  INV_X1 u2_u6_u1_U35 (.A( u2_u6_u1_n148 ) , .ZN( u2_u6_u1_n187 ) );
  AOI211_X1 u2_u6_u1_U36 (.B( u2_u6_u1_n117 ) , .A( u2_u6_u1_n118 ) , .ZN( u2_u6_u1_n119 ) , .C2( u2_u6_u1_n146 ) , .C1( u2_u6_u1_n159 ) );
  NOR2_X1 u2_u6_u1_U37 (.A1( u2_u6_u1_n168 ) , .A2( u2_u6_u1_n176 ) , .ZN( u2_u6_u1_n98 ) );
  AOI211_X1 u2_u6_u1_U38 (.B( u2_u6_u1_n162 ) , .A( u2_u6_u1_n163 ) , .C2( u2_u6_u1_n164 ) , .ZN( u2_u6_u1_n165 ) , .C1( u2_u6_u1_n171 ) );
  AOI21_X1 u2_u6_u1_U39 (.A( u2_u6_u1_n160 ) , .B2( u2_u6_u1_n161 ) , .ZN( u2_u6_u1_n162 ) , .B1( u2_u6_u1_n182 ) );
  AOI221_X1 u2_u6_u1_U4 (.A( u2_u6_u1_n138 ) , .C2( u2_u6_u1_n139 ) , .C1( u2_u6_u1_n140 ) , .B2( u2_u6_u1_n141 ) , .ZN( u2_u6_u1_n142 ) , .B1( u2_u6_u1_n175 ) );
  OR2_X1 u2_u6_u1_U40 (.A2( u2_u6_u1_n157 ) , .A1( u2_u6_u1_n158 ) , .ZN( u2_u6_u1_n163 ) );
  NAND2_X1 u2_u6_u1_U41 (.A1( u2_u6_u1_n128 ) , .ZN( u2_u6_u1_n146 ) , .A2( u2_u6_u1_n160 ) );
  NAND2_X1 u2_u6_u1_U42 (.A2( u2_u6_u1_n112 ) , .ZN( u2_u6_u1_n139 ) , .A1( u2_u6_u1_n152 ) );
  NAND2_X1 u2_u6_u1_U43 (.A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n156 ) , .A2( u2_u6_u1_n99 ) );
  NOR2_X1 u2_u6_u1_U44 (.ZN( u2_u6_u1_n117 ) , .A1( u2_u6_u1_n121 ) , .A2( u2_u6_u1_n160 ) );
  OAI21_X1 u2_u6_u1_U45 (.B2( u2_u6_u1_n123 ) , .ZN( u2_u6_u1_n145 ) , .B1( u2_u6_u1_n160 ) , .A( u2_u6_u1_n185 ) );
  INV_X1 u2_u6_u1_U46 (.A( u2_u6_u1_n122 ) , .ZN( u2_u6_u1_n185 ) );
  AOI21_X1 u2_u6_u1_U47 (.B2( u2_u6_u1_n120 ) , .B1( u2_u6_u1_n121 ) , .ZN( u2_u6_u1_n122 ) , .A( u2_u6_u1_n128 ) );
  AOI21_X1 u2_u6_u1_U48 (.A( u2_u6_u1_n128 ) , .B2( u2_u6_u1_n129 ) , .ZN( u2_u6_u1_n130 ) , .B1( u2_u6_u1_n150 ) );
  NAND2_X1 u2_u6_u1_U49 (.ZN( u2_u6_u1_n112 ) , .A1( u2_u6_u1_n169 ) , .A2( u2_u6_u1_n170 ) );
  AOI211_X1 u2_u6_u1_U5 (.ZN( u2_u6_u1_n124 ) , .A( u2_u6_u1_n138 ) , .C2( u2_u6_u1_n139 ) , .B( u2_u6_u1_n145 ) , .C1( u2_u6_u1_n147 ) );
  NAND2_X1 u2_u6_u1_U50 (.ZN( u2_u6_u1_n129 ) , .A2( u2_u6_u1_n95 ) , .A1( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U51 (.A1( u2_u6_u1_n102 ) , .ZN( u2_u6_u1_n154 ) , .A2( u2_u6_u1_n99 ) );
  NAND2_X1 u2_u6_u1_U52 (.A2( u2_u6_u1_n100 ) , .ZN( u2_u6_u1_n135 ) , .A1( u2_u6_u1_n99 ) );
  AOI21_X1 u2_u6_u1_U53 (.A( u2_u6_u1_n152 ) , .B2( u2_u6_u1_n153 ) , .B1( u2_u6_u1_n154 ) , .ZN( u2_u6_u1_n158 ) );
  INV_X1 u2_u6_u1_U54 (.A( u2_u6_u1_n160 ) , .ZN( u2_u6_u1_n175 ) );
  NAND2_X1 u2_u6_u1_U55 (.A1( u2_u6_u1_n100 ) , .ZN( u2_u6_u1_n116 ) , .A2( u2_u6_u1_n95 ) );
  NAND2_X1 u2_u6_u1_U56 (.A1( u2_u6_u1_n102 ) , .ZN( u2_u6_u1_n131 ) , .A2( u2_u6_u1_n95 ) );
  NAND2_X1 u2_u6_u1_U57 (.A2( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n121 ) , .A1( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U58 (.A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n153 ) , .A2( u2_u6_u1_n98 ) );
  NAND2_X1 u2_u6_u1_U59 (.A2( u2_u6_u1_n104 ) , .A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n133 ) );
  AOI22_X1 u2_u6_u1_U6 (.B2( u2_u6_u1_n136 ) , .A2( u2_u6_u1_n137 ) , .ZN( u2_u6_u1_n143 ) , .A1( u2_u6_u1_n171 ) , .B1( u2_u6_u1_n173 ) );
  NAND2_X1 u2_u6_u1_U60 (.ZN( u2_u6_u1_n150 ) , .A2( u2_u6_u1_n98 ) , .A1( u2_u6_u1_n99 ) );
  NAND2_X1 u2_u6_u1_U61 (.A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n155 ) , .A2( u2_u6_u1_n95 ) );
  OAI21_X1 u2_u6_u1_U62 (.ZN( u2_u6_u1_n109 ) , .B1( u2_u6_u1_n129 ) , .B2( u2_u6_u1_n160 ) , .A( u2_u6_u1_n167 ) );
  NAND2_X1 u2_u6_u1_U63 (.A2( u2_u6_u1_n100 ) , .A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n120 ) );
  NAND2_X1 u2_u6_u1_U64 (.A1( u2_u6_u1_n102 ) , .A2( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n115 ) );
  NAND2_X1 u2_u6_u1_U65 (.A2( u2_u6_u1_n100 ) , .A1( u2_u6_u1_n104 ) , .ZN( u2_u6_u1_n151 ) );
  NAND2_X1 u2_u6_u1_U66 (.A2( u2_u6_u1_n103 ) , .A1( u2_u6_u1_n105 ) , .ZN( u2_u6_u1_n161 ) );
  INV_X1 u2_u6_u1_U67 (.A( u2_u6_u1_n152 ) , .ZN( u2_u6_u1_n173 ) );
  INV_X1 u2_u6_u1_U68 (.A( u2_u6_u1_n128 ) , .ZN( u2_u6_u1_n172 ) );
  NAND2_X1 u2_u6_u1_U69 (.A2( u2_u6_u1_n102 ) , .A1( u2_u6_u1_n103 ) , .ZN( u2_u6_u1_n123 ) );
  INV_X1 u2_u6_u1_U7 (.A( u2_u6_u1_n147 ) , .ZN( u2_u6_u1_n181 ) );
  NOR2_X1 u2_u6_u1_U70 (.A2( u2_u6_X_7 ) , .A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n95 ) );
  NOR2_X1 u2_u6_u1_U71 (.A1( u2_u6_X_12 ) , .A2( u2_u6_X_9 ) , .ZN( u2_u6_u1_n100 ) );
  NOR2_X1 u2_u6_u1_U72 (.A2( u2_u6_X_8 ) , .A1( u2_u6_u1_n177 ) , .ZN( u2_u6_u1_n99 ) );
  NOR2_X1 u2_u6_u1_U73 (.A2( u2_u6_X_12 ) , .ZN( u2_u6_u1_n102 ) , .A1( u2_u6_u1_n176 ) );
  NOR2_X1 u2_u6_u1_U74 (.A2( u2_u6_X_9 ) , .ZN( u2_u6_u1_n105 ) , .A1( u2_u6_u1_n168 ) );
  NAND2_X1 u2_u6_u1_U75 (.A1( u2_u6_X_10 ) , .ZN( u2_u6_u1_n160 ) , .A2( u2_u6_u1_n169 ) );
  NAND2_X1 u2_u6_u1_U76 (.A2( u2_u6_X_10 ) , .A1( u2_u6_X_11 ) , .ZN( u2_u6_u1_n152 ) );
  NAND2_X1 u2_u6_u1_U77 (.A1( u2_u6_X_11 ) , .ZN( u2_u6_u1_n128 ) , .A2( u2_u6_u1_n170 ) );
  AND2_X1 u2_u6_u1_U78 (.A2( u2_u6_X_7 ) , .A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n104 ) );
  AND2_X1 u2_u6_u1_U79 (.A1( u2_u6_X_8 ) , .ZN( u2_u6_u1_n103 ) , .A2( u2_u6_u1_n177 ) );
  NOR2_X1 u2_u6_u1_U8 (.A1( u2_u6_u1_n112 ) , .A2( u2_u6_u1_n116 ) , .ZN( u2_u6_u1_n118 ) );
  INV_X1 u2_u6_u1_U80 (.A( u2_u6_X_10 ) , .ZN( u2_u6_u1_n170 ) );
  INV_X1 u2_u6_u1_U81 (.A( u2_u6_X_9 ) , .ZN( u2_u6_u1_n176 ) );
  INV_X1 u2_u6_u1_U82 (.A( u2_u6_X_11 ) , .ZN( u2_u6_u1_n169 ) );
  INV_X1 u2_u6_u1_U83 (.A( u2_u6_X_12 ) , .ZN( u2_u6_u1_n168 ) );
  INV_X1 u2_u6_u1_U84 (.A( u2_u6_X_7 ) , .ZN( u2_u6_u1_n177 ) );
  NAND4_X1 u2_u6_u1_U85 (.ZN( u2_out6_28 ) , .A4( u2_u6_u1_n124 ) , .A3( u2_u6_u1_n125 ) , .A2( u2_u6_u1_n126 ) , .A1( u2_u6_u1_n127 ) );
  OAI21_X1 u2_u6_u1_U86 (.ZN( u2_u6_u1_n127 ) , .B2( u2_u6_u1_n139 ) , .B1( u2_u6_u1_n175 ) , .A( u2_u6_u1_n183 ) );
  OAI21_X1 u2_u6_u1_U87 (.ZN( u2_u6_u1_n126 ) , .B2( u2_u6_u1_n140 ) , .A( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n178 ) );
  NAND4_X1 u2_u6_u1_U88 (.ZN( u2_out6_18 ) , .A4( u2_u6_u1_n165 ) , .A3( u2_u6_u1_n166 ) , .A1( u2_u6_u1_n167 ) , .A2( u2_u6_u1_n186 ) );
  AOI22_X1 u2_u6_u1_U89 (.B2( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n147 ) , .A2( u2_u6_u1_n148 ) , .ZN( u2_u6_u1_n166 ) , .A1( u2_u6_u1_n172 ) );
  OAI21_X1 u2_u6_u1_U9 (.ZN( u2_u6_u1_n101 ) , .B1( u2_u6_u1_n141 ) , .A( u2_u6_u1_n146 ) , .B2( u2_u6_u1_n183 ) );
  INV_X1 u2_u6_u1_U90 (.A( u2_u6_u1_n145 ) , .ZN( u2_u6_u1_n186 ) );
  NAND4_X1 u2_u6_u1_U91 (.ZN( u2_out6_2 ) , .A4( u2_u6_u1_n142 ) , .A3( u2_u6_u1_n143 ) , .A2( u2_u6_u1_n144 ) , .A1( u2_u6_u1_n179 ) );
  OAI21_X1 u2_u6_u1_U92 (.B2( u2_u6_u1_n132 ) , .ZN( u2_u6_u1_n144 ) , .A( u2_u6_u1_n146 ) , .B1( u2_u6_u1_n180 ) );
  INV_X1 u2_u6_u1_U93 (.A( u2_u6_u1_n130 ) , .ZN( u2_u6_u1_n179 ) );
  OR4_X1 u2_u6_u1_U94 (.ZN( u2_out6_13 ) , .A4( u2_u6_u1_n108 ) , .A3( u2_u6_u1_n109 ) , .A2( u2_u6_u1_n110 ) , .A1( u2_u6_u1_n111 ) );
  AOI21_X1 u2_u6_u1_U95 (.ZN( u2_u6_u1_n111 ) , .A( u2_u6_u1_n128 ) , .B2( u2_u6_u1_n131 ) , .B1( u2_u6_u1_n135 ) );
  AOI21_X1 u2_u6_u1_U96 (.ZN( u2_u6_u1_n110 ) , .A( u2_u6_u1_n116 ) , .B1( u2_u6_u1_n152 ) , .B2( u2_u6_u1_n160 ) );
  NAND3_X1 u2_u6_u1_U97 (.A3( u2_u6_u1_n149 ) , .A2( u2_u6_u1_n150 ) , .A1( u2_u6_u1_n151 ) , .ZN( u2_u6_u1_n164 ) );
  NAND3_X1 u2_u6_u1_U98 (.A3( u2_u6_u1_n134 ) , .A2( u2_u6_u1_n135 ) , .ZN( u2_u6_u1_n136 ) , .A1( u2_u6_u1_n151 ) );
  NAND3_X1 u2_u6_u1_U99 (.A1( u2_u6_u1_n133 ) , .ZN( u2_u6_u1_n137 ) , .A2( u2_u6_u1_n154 ) , .A3( u2_u6_u1_n181 ) );
  OAI22_X1 u2_u6_u2_U10 (.B1( u2_u6_u2_n151 ) , .A2( u2_u6_u2_n152 ) , .A1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n160 ) , .B2( u2_u6_u2_n168 ) );
  NAND3_X1 u2_u6_u2_U100 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n98 ) );
  NOR3_X1 u2_u6_u2_U11 (.A1( u2_u6_u2_n150 ) , .ZN( u2_u6_u2_n151 ) , .A3( u2_u6_u2_n175 ) , .A2( u2_u6_u2_n188 ) );
  AOI21_X1 u2_u6_u2_U12 (.B2( u2_u6_u2_n123 ) , .ZN( u2_u6_u2_n125 ) , .A( u2_u6_u2_n171 ) , .B1( u2_u6_u2_n184 ) );
  INV_X1 u2_u6_u2_U13 (.A( u2_u6_u2_n150 ) , .ZN( u2_u6_u2_n184 ) );
  AOI21_X1 u2_u6_u2_U14 (.ZN( u2_u6_u2_n144 ) , .B2( u2_u6_u2_n155 ) , .A( u2_u6_u2_n172 ) , .B1( u2_u6_u2_n185 ) );
  AOI21_X1 u2_u6_u2_U15 (.B2( u2_u6_u2_n143 ) , .ZN( u2_u6_u2_n145 ) , .B1( u2_u6_u2_n152 ) , .A( u2_u6_u2_n171 ) );
  INV_X1 u2_u6_u2_U16 (.A( u2_u6_u2_n156 ) , .ZN( u2_u6_u2_n171 ) );
  INV_X1 u2_u6_u2_U17 (.A( u2_u6_u2_n120 ) , .ZN( u2_u6_u2_n188 ) );
  NAND2_X1 u2_u6_u2_U18 (.A2( u2_u6_u2_n122 ) , .ZN( u2_u6_u2_n150 ) , .A1( u2_u6_u2_n152 ) );
  INV_X1 u2_u6_u2_U19 (.A( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n170 ) );
  INV_X1 u2_u6_u2_U20 (.A( u2_u6_u2_n137 ) , .ZN( u2_u6_u2_n173 ) );
  NAND2_X1 u2_u6_u2_U21 (.A1( u2_u6_u2_n132 ) , .A2( u2_u6_u2_n139 ) , .ZN( u2_u6_u2_n157 ) );
  INV_X1 u2_u6_u2_U22 (.A( u2_u6_u2_n113 ) , .ZN( u2_u6_u2_n178 ) );
  INV_X1 u2_u6_u2_U23 (.A( u2_u6_u2_n139 ) , .ZN( u2_u6_u2_n175 ) );
  INV_X1 u2_u6_u2_U24 (.A( u2_u6_u2_n155 ) , .ZN( u2_u6_u2_n181 ) );
  INV_X1 u2_u6_u2_U25 (.A( u2_u6_u2_n119 ) , .ZN( u2_u6_u2_n177 ) );
  INV_X1 u2_u6_u2_U26 (.A( u2_u6_u2_n116 ) , .ZN( u2_u6_u2_n180 ) );
  INV_X1 u2_u6_u2_U27 (.A( u2_u6_u2_n131 ) , .ZN( u2_u6_u2_n179 ) );
  INV_X1 u2_u6_u2_U28 (.A( u2_u6_u2_n154 ) , .ZN( u2_u6_u2_n176 ) );
  NAND2_X1 u2_u6_u2_U29 (.A2( u2_u6_u2_n116 ) , .A1( u2_u6_u2_n117 ) , .ZN( u2_u6_u2_n118 ) );
  NOR2_X1 u2_u6_u2_U3 (.ZN( u2_u6_u2_n121 ) , .A2( u2_u6_u2_n177 ) , .A1( u2_u6_u2_n180 ) );
  INV_X1 u2_u6_u2_U30 (.A( u2_u6_u2_n132 ) , .ZN( u2_u6_u2_n182 ) );
  INV_X1 u2_u6_u2_U31 (.A( u2_u6_u2_n158 ) , .ZN( u2_u6_u2_n183 ) );
  OAI21_X1 u2_u6_u2_U32 (.A( u2_u6_u2_n156 ) , .B1( u2_u6_u2_n157 ) , .ZN( u2_u6_u2_n158 ) , .B2( u2_u6_u2_n179 ) );
  NOR2_X1 u2_u6_u2_U33 (.ZN( u2_u6_u2_n156 ) , .A1( u2_u6_u2_n166 ) , .A2( u2_u6_u2_n169 ) );
  NOR2_X1 u2_u6_u2_U34 (.A2( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n137 ) , .A1( u2_u6_u2_n140 ) );
  NOR2_X1 u2_u6_u2_U35 (.A2( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n153 ) , .A1( u2_u6_u2_n156 ) );
  AOI211_X1 u2_u6_u2_U36 (.ZN( u2_u6_u2_n130 ) , .C1( u2_u6_u2_n138 ) , .C2( u2_u6_u2_n179 ) , .B( u2_u6_u2_n96 ) , .A( u2_u6_u2_n97 ) );
  OAI22_X1 u2_u6_u2_U37 (.B1( u2_u6_u2_n133 ) , .A2( u2_u6_u2_n137 ) , .A1( u2_u6_u2_n152 ) , .B2( u2_u6_u2_n168 ) , .ZN( u2_u6_u2_n97 ) );
  OAI221_X1 u2_u6_u2_U38 (.B1( u2_u6_u2_n113 ) , .C1( u2_u6_u2_n132 ) , .A( u2_u6_u2_n149 ) , .B2( u2_u6_u2_n171 ) , .C2( u2_u6_u2_n172 ) , .ZN( u2_u6_u2_n96 ) );
  OAI221_X1 u2_u6_u2_U39 (.A( u2_u6_u2_n115 ) , .C2( u2_u6_u2_n123 ) , .B2( u2_u6_u2_n143 ) , .B1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n163 ) , .C1( u2_u6_u2_n168 ) );
  INV_X1 u2_u6_u2_U4 (.A( u2_u6_u2_n134 ) , .ZN( u2_u6_u2_n185 ) );
  OAI21_X1 u2_u6_u2_U40 (.A( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n115 ) , .B1( u2_u6_u2_n176 ) , .B2( u2_u6_u2_n178 ) );
  OAI221_X1 u2_u6_u2_U41 (.A( u2_u6_u2_n135 ) , .B2( u2_u6_u2_n136 ) , .B1( u2_u6_u2_n137 ) , .ZN( u2_u6_u2_n162 ) , .C2( u2_u6_u2_n167 ) , .C1( u2_u6_u2_n185 ) );
  AND3_X1 u2_u6_u2_U42 (.A3( u2_u6_u2_n131 ) , .A2( u2_u6_u2_n132 ) , .A1( u2_u6_u2_n133 ) , .ZN( u2_u6_u2_n136 ) );
  AOI22_X1 u2_u6_u2_U43 (.ZN( u2_u6_u2_n135 ) , .B1( u2_u6_u2_n140 ) , .A1( u2_u6_u2_n156 ) , .B2( u2_u6_u2_n180 ) , .A2( u2_u6_u2_n188 ) );
  AOI21_X1 u2_u6_u2_U44 (.ZN( u2_u6_u2_n149 ) , .B1( u2_u6_u2_n173 ) , .B2( u2_u6_u2_n188 ) , .A( u2_u6_u2_n95 ) );
  AND3_X1 u2_u6_u2_U45 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n156 ) , .ZN( u2_u6_u2_n95 ) );
  OAI21_X1 u2_u6_u2_U46 (.A( u2_u6_u2_n141 ) , .B2( u2_u6_u2_n142 ) , .ZN( u2_u6_u2_n146 ) , .B1( u2_u6_u2_n153 ) );
  OAI21_X1 u2_u6_u2_U47 (.A( u2_u6_u2_n140 ) , .ZN( u2_u6_u2_n141 ) , .B1( u2_u6_u2_n176 ) , .B2( u2_u6_u2_n177 ) );
  NOR3_X1 u2_u6_u2_U48 (.ZN( u2_u6_u2_n142 ) , .A3( u2_u6_u2_n175 ) , .A2( u2_u6_u2_n178 ) , .A1( u2_u6_u2_n181 ) );
  OAI21_X1 u2_u6_u2_U49 (.A( u2_u6_u2_n101 ) , .B2( u2_u6_u2_n121 ) , .B1( u2_u6_u2_n153 ) , .ZN( u2_u6_u2_n164 ) );
  NOR4_X1 u2_u6_u2_U5 (.A4( u2_u6_u2_n124 ) , .A3( u2_u6_u2_n125 ) , .A2( u2_u6_u2_n126 ) , .A1( u2_u6_u2_n127 ) , .ZN( u2_u6_u2_n128 ) );
  NAND2_X1 u2_u6_u2_U50 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n155 ) );
  NAND2_X1 u2_u6_u2_U51 (.A2( u2_u6_u2_n105 ) , .A1( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n143 ) );
  NAND2_X1 u2_u6_u2_U52 (.A1( u2_u6_u2_n104 ) , .A2( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n152 ) );
  NAND2_X1 u2_u6_u2_U53 (.A1( u2_u6_u2_n100 ) , .A2( u2_u6_u2_n105 ) , .ZN( u2_u6_u2_n132 ) );
  INV_X1 u2_u6_u2_U54 (.A( u2_u6_u2_n140 ) , .ZN( u2_u6_u2_n168 ) );
  INV_X1 u2_u6_u2_U55 (.A( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n167 ) );
  INV_X1 u2_u6_u2_U56 (.ZN( u2_u6_u2_n187 ) , .A( u2_u6_u2_n99 ) );
  OAI21_X1 u2_u6_u2_U57 (.B1( u2_u6_u2_n137 ) , .B2( u2_u6_u2_n143 ) , .A( u2_u6_u2_n98 ) , .ZN( u2_u6_u2_n99 ) );
  NAND2_X1 u2_u6_u2_U58 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n113 ) );
  NAND2_X1 u2_u6_u2_U59 (.A1( u2_u6_u2_n106 ) , .A2( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n131 ) );
  AOI21_X1 u2_u6_u2_U6 (.B2( u2_u6_u2_n119 ) , .ZN( u2_u6_u2_n127 ) , .A( u2_u6_u2_n137 ) , .B1( u2_u6_u2_n155 ) );
  NAND2_X1 u2_u6_u2_U60 (.A1( u2_u6_u2_n103 ) , .A2( u2_u6_u2_n107 ) , .ZN( u2_u6_u2_n139 ) );
  NAND2_X1 u2_u6_u2_U61 (.A1( u2_u6_u2_n103 ) , .A2( u2_u6_u2_n105 ) , .ZN( u2_u6_u2_n133 ) );
  NAND2_X1 u2_u6_u2_U62 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n103 ) , .ZN( u2_u6_u2_n154 ) );
  NAND2_X1 u2_u6_u2_U63 (.A2( u2_u6_u2_n103 ) , .A1( u2_u6_u2_n104 ) , .ZN( u2_u6_u2_n119 ) );
  NAND2_X1 u2_u6_u2_U64 (.A2( u2_u6_u2_n107 ) , .A1( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n123 ) );
  NAND2_X1 u2_u6_u2_U65 (.A1( u2_u6_u2_n104 ) , .A2( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n122 ) );
  INV_X1 u2_u6_u2_U66 (.A( u2_u6_u2_n114 ) , .ZN( u2_u6_u2_n172 ) );
  NAND2_X1 u2_u6_u2_U67 (.A2( u2_u6_u2_n100 ) , .A1( u2_u6_u2_n102 ) , .ZN( u2_u6_u2_n116 ) );
  NAND2_X1 u2_u6_u2_U68 (.A1( u2_u6_u2_n102 ) , .A2( u2_u6_u2_n108 ) , .ZN( u2_u6_u2_n120 ) );
  NAND2_X1 u2_u6_u2_U69 (.A2( u2_u6_u2_n105 ) , .A1( u2_u6_u2_n106 ) , .ZN( u2_u6_u2_n117 ) );
  AOI21_X1 u2_u6_u2_U7 (.ZN( u2_u6_u2_n124 ) , .B1( u2_u6_u2_n131 ) , .B2( u2_u6_u2_n143 ) , .A( u2_u6_u2_n172 ) );
  NOR2_X1 u2_u6_u2_U70 (.A2( u2_u6_X_16 ) , .ZN( u2_u6_u2_n140 ) , .A1( u2_u6_u2_n166 ) );
  NOR2_X1 u2_u6_u2_U71 (.A2( u2_u6_X_13 ) , .A1( u2_u6_X_14 ) , .ZN( u2_u6_u2_n100 ) );
  NOR2_X1 u2_u6_u2_U72 (.A2( u2_u6_X_16 ) , .A1( u2_u6_X_17 ) , .ZN( u2_u6_u2_n138 ) );
  NOR2_X1 u2_u6_u2_U73 (.A2( u2_u6_X_15 ) , .A1( u2_u6_X_18 ) , .ZN( u2_u6_u2_n104 ) );
  NOR2_X1 u2_u6_u2_U74 (.A2( u2_u6_X_14 ) , .ZN( u2_u6_u2_n103 ) , .A1( u2_u6_u2_n174 ) );
  NOR2_X1 u2_u6_u2_U75 (.A2( u2_u6_X_15 ) , .ZN( u2_u6_u2_n102 ) , .A1( u2_u6_u2_n165 ) );
  NOR2_X1 u2_u6_u2_U76 (.A2( u2_u6_X_17 ) , .ZN( u2_u6_u2_n114 ) , .A1( u2_u6_u2_n169 ) );
  AND2_X1 u2_u6_u2_U77 (.A1( u2_u6_X_15 ) , .ZN( u2_u6_u2_n105 ) , .A2( u2_u6_u2_n165 ) );
  AND2_X1 u2_u6_u2_U78 (.A2( u2_u6_X_15 ) , .A1( u2_u6_X_18 ) , .ZN( u2_u6_u2_n107 ) );
  AND2_X1 u2_u6_u2_U79 (.A1( u2_u6_X_14 ) , .ZN( u2_u6_u2_n106 ) , .A2( u2_u6_u2_n174 ) );
  AOI21_X1 u2_u6_u2_U8 (.B2( u2_u6_u2_n120 ) , .B1( u2_u6_u2_n121 ) , .ZN( u2_u6_u2_n126 ) , .A( u2_u6_u2_n167 ) );
  AND2_X1 u2_u6_u2_U80 (.A1( u2_u6_X_13 ) , .A2( u2_u6_X_14 ) , .ZN( u2_u6_u2_n108 ) );
  INV_X1 u2_u6_u2_U81 (.A( u2_u6_X_16 ) , .ZN( u2_u6_u2_n169 ) );
  INV_X1 u2_u6_u2_U82 (.A( u2_u6_X_17 ) , .ZN( u2_u6_u2_n166 ) );
  INV_X1 u2_u6_u2_U83 (.A( u2_u6_X_13 ) , .ZN( u2_u6_u2_n174 ) );
  INV_X1 u2_u6_u2_U84 (.A( u2_u6_X_18 ) , .ZN( u2_u6_u2_n165 ) );
  NAND4_X1 u2_u6_u2_U85 (.ZN( u2_out6_30 ) , .A4( u2_u6_u2_n147 ) , .A3( u2_u6_u2_n148 ) , .A2( u2_u6_u2_n149 ) , .A1( u2_u6_u2_n187 ) );
  AOI21_X1 u2_u6_u2_U86 (.B2( u2_u6_u2_n138 ) , .ZN( u2_u6_u2_n148 ) , .A( u2_u6_u2_n162 ) , .B1( u2_u6_u2_n182 ) );
  NOR3_X1 u2_u6_u2_U87 (.A3( u2_u6_u2_n144 ) , .A2( u2_u6_u2_n145 ) , .A1( u2_u6_u2_n146 ) , .ZN( u2_u6_u2_n147 ) );
  NAND4_X1 u2_u6_u2_U88 (.ZN( u2_out6_24 ) , .A4( u2_u6_u2_n111 ) , .A3( u2_u6_u2_n112 ) , .A1( u2_u6_u2_n130 ) , .A2( u2_u6_u2_n187 ) );
  AOI221_X1 u2_u6_u2_U89 (.A( u2_u6_u2_n109 ) , .B1( u2_u6_u2_n110 ) , .ZN( u2_u6_u2_n111 ) , .C1( u2_u6_u2_n134 ) , .C2( u2_u6_u2_n170 ) , .B2( u2_u6_u2_n173 ) );
  OAI22_X1 u2_u6_u2_U9 (.ZN( u2_u6_u2_n109 ) , .A2( u2_u6_u2_n113 ) , .B2( u2_u6_u2_n133 ) , .B1( u2_u6_u2_n167 ) , .A1( u2_u6_u2_n168 ) );
  AOI21_X1 u2_u6_u2_U90 (.ZN( u2_u6_u2_n112 ) , .B2( u2_u6_u2_n156 ) , .A( u2_u6_u2_n164 ) , .B1( u2_u6_u2_n181 ) );
  NAND4_X1 u2_u6_u2_U91 (.ZN( u2_out6_16 ) , .A4( u2_u6_u2_n128 ) , .A3( u2_u6_u2_n129 ) , .A1( u2_u6_u2_n130 ) , .A2( u2_u6_u2_n186 ) );
  AOI22_X1 u2_u6_u2_U92 (.A2( u2_u6_u2_n118 ) , .ZN( u2_u6_u2_n129 ) , .A1( u2_u6_u2_n140 ) , .B1( u2_u6_u2_n157 ) , .B2( u2_u6_u2_n170 ) );
  INV_X1 u2_u6_u2_U93 (.A( u2_u6_u2_n163 ) , .ZN( u2_u6_u2_n186 ) );
  OR4_X1 u2_u6_u2_U94 (.ZN( u2_out6_6 ) , .A4( u2_u6_u2_n161 ) , .A3( u2_u6_u2_n162 ) , .A2( u2_u6_u2_n163 ) , .A1( u2_u6_u2_n164 ) );
  OR3_X1 u2_u6_u2_U95 (.A2( u2_u6_u2_n159 ) , .A1( u2_u6_u2_n160 ) , .ZN( u2_u6_u2_n161 ) , .A3( u2_u6_u2_n183 ) );
  AOI21_X1 u2_u6_u2_U96 (.B2( u2_u6_u2_n154 ) , .B1( u2_u6_u2_n155 ) , .ZN( u2_u6_u2_n159 ) , .A( u2_u6_u2_n167 ) );
  NAND3_X1 u2_u6_u2_U97 (.A2( u2_u6_u2_n117 ) , .A1( u2_u6_u2_n122 ) , .A3( u2_u6_u2_n123 ) , .ZN( u2_u6_u2_n134 ) );
  NAND3_X1 u2_u6_u2_U98 (.ZN( u2_u6_u2_n110 ) , .A2( u2_u6_u2_n131 ) , .A3( u2_u6_u2_n139 ) , .A1( u2_u6_u2_n154 ) );
  NAND3_X1 u2_u6_u2_U99 (.A2( u2_u6_u2_n100 ) , .ZN( u2_u6_u2_n101 ) , .A1( u2_u6_u2_n104 ) , .A3( u2_u6_u2_n114 ) );
  XOR2_X1 u2_u9_U1 (.B( u2_K10_9 ) , .A( u2_R8_6 ) , .Z( u2_u9_X_9 ) );
  XOR2_X1 u2_u9_U2 (.B( u2_K10_8 ) , .A( u2_R8_5 ) , .Z( u2_u9_X_8 ) );
  XOR2_X1 u2_u9_U3 (.B( u2_K10_7 ) , .A( u2_R8_4 ) , .Z( u2_u9_X_7 ) );
  XOR2_X1 u2_u9_U40 (.B( u2_K10_18 ) , .A( u2_R8_13 ) , .Z( u2_u9_X_18 ) );
  XOR2_X1 u2_u9_U41 (.B( u2_K10_17 ) , .A( u2_R8_12 ) , .Z( u2_u9_X_17 ) );
  XOR2_X1 u2_u9_U42 (.B( u2_K10_16 ) , .A( u2_R8_11 ) , .Z( u2_u9_X_16 ) );
  XOR2_X1 u2_u9_U43 (.B( u2_K10_15 ) , .A( u2_R8_10 ) , .Z( u2_u9_X_15 ) );
  XOR2_X1 u2_u9_U44 (.B( u2_K10_14 ) , .A( u2_R8_9 ) , .Z( u2_u9_X_14 ) );
  XOR2_X1 u2_u9_U45 (.B( u2_K10_13 ) , .A( u2_R8_8 ) , .Z( u2_u9_X_13 ) );
  XOR2_X1 u2_u9_U46 (.B( u2_K10_12 ) , .A( u2_R8_9 ) , .Z( u2_u9_X_12 ) );
  XOR2_X1 u2_u9_U47 (.B( u2_K10_11 ) , .A( u2_R8_8 ) , .Z( u2_u9_X_11 ) );
  XOR2_X1 u2_u9_U48 (.B( u2_K10_10 ) , .A( u2_R8_7 ) , .Z( u2_u9_X_10 ) );
  NOR2_X1 u2_u9_u1_U10 (.A1( u2_u9_u1_n112 ) , .A2( u2_u9_u1_n116 ) , .ZN( u2_u9_u1_n118 ) );
  NAND3_X1 u2_u9_u1_U100 (.ZN( u2_u9_u1_n113 ) , .A1( u2_u9_u1_n120 ) , .A3( u2_u9_u1_n133 ) , .A2( u2_u9_u1_n155 ) );
  OAI21_X1 u2_u9_u1_U11 (.ZN( u2_u9_u1_n101 ) , .B1( u2_u9_u1_n141 ) , .A( u2_u9_u1_n146 ) , .B2( u2_u9_u1_n183 ) );
  AOI21_X1 u2_u9_u1_U12 (.B2( u2_u9_u1_n155 ) , .B1( u2_u9_u1_n156 ) , .ZN( u2_u9_u1_n157 ) , .A( u2_u9_u1_n174 ) );
  NAND2_X1 u2_u9_u1_U13 (.ZN( u2_u9_u1_n140 ) , .A2( u2_u9_u1_n150 ) , .A1( u2_u9_u1_n155 ) );
  NAND2_X1 u2_u9_u1_U14 (.A1( u2_u9_u1_n131 ) , .ZN( u2_u9_u1_n147 ) , .A2( u2_u9_u1_n153 ) );
  INV_X1 u2_u9_u1_U15 (.A( u2_u9_u1_n139 ) , .ZN( u2_u9_u1_n174 ) );
  OR4_X1 u2_u9_u1_U16 (.A4( u2_u9_u1_n106 ) , .A3( u2_u9_u1_n107 ) , .ZN( u2_u9_u1_n108 ) , .A1( u2_u9_u1_n117 ) , .A2( u2_u9_u1_n184 ) );
  AOI21_X1 u2_u9_u1_U17 (.ZN( u2_u9_u1_n106 ) , .A( u2_u9_u1_n112 ) , .B1( u2_u9_u1_n154 ) , .B2( u2_u9_u1_n156 ) );
  AOI21_X1 u2_u9_u1_U18 (.ZN( u2_u9_u1_n107 ) , .B1( u2_u9_u1_n134 ) , .B2( u2_u9_u1_n149 ) , .A( u2_u9_u1_n174 ) );
  INV_X1 u2_u9_u1_U19 (.A( u2_u9_u1_n101 ) , .ZN( u2_u9_u1_n184 ) );
  INV_X1 u2_u9_u1_U20 (.A( u2_u9_u1_n112 ) , .ZN( u2_u9_u1_n171 ) );
  NAND2_X1 u2_u9_u1_U21 (.ZN( u2_u9_u1_n141 ) , .A1( u2_u9_u1_n153 ) , .A2( u2_u9_u1_n156 ) );
  AND2_X1 u2_u9_u1_U22 (.A1( u2_u9_u1_n123 ) , .ZN( u2_u9_u1_n134 ) , .A2( u2_u9_u1_n161 ) );
  NAND2_X1 u2_u9_u1_U23 (.A2( u2_u9_u1_n115 ) , .A1( u2_u9_u1_n116 ) , .ZN( u2_u9_u1_n148 ) );
  NAND2_X1 u2_u9_u1_U24 (.A2( u2_u9_u1_n133 ) , .A1( u2_u9_u1_n135 ) , .ZN( u2_u9_u1_n159 ) );
  NAND2_X1 u2_u9_u1_U25 (.A2( u2_u9_u1_n115 ) , .A1( u2_u9_u1_n120 ) , .ZN( u2_u9_u1_n132 ) );
  INV_X1 u2_u9_u1_U26 (.A( u2_u9_u1_n154 ) , .ZN( u2_u9_u1_n178 ) );
  INV_X1 u2_u9_u1_U27 (.A( u2_u9_u1_n151 ) , .ZN( u2_u9_u1_n183 ) );
  AND2_X1 u2_u9_u1_U28 (.A1( u2_u9_u1_n129 ) , .A2( u2_u9_u1_n133 ) , .ZN( u2_u9_u1_n149 ) );
  INV_X1 u2_u9_u1_U29 (.A( u2_u9_u1_n131 ) , .ZN( u2_u9_u1_n180 ) );
  INV_X1 u2_u9_u1_U3 (.A( u2_u9_u1_n159 ) , .ZN( u2_u9_u1_n182 ) );
  OAI221_X1 u2_u9_u1_U30 (.A( u2_u9_u1_n119 ) , .C2( u2_u9_u1_n129 ) , .ZN( u2_u9_u1_n138 ) , .B2( u2_u9_u1_n152 ) , .C1( u2_u9_u1_n174 ) , .B1( u2_u9_u1_n187 ) );
  INV_X1 u2_u9_u1_U31 (.A( u2_u9_u1_n148 ) , .ZN( u2_u9_u1_n187 ) );
  AOI211_X1 u2_u9_u1_U32 (.B( u2_u9_u1_n117 ) , .A( u2_u9_u1_n118 ) , .ZN( u2_u9_u1_n119 ) , .C2( u2_u9_u1_n146 ) , .C1( u2_u9_u1_n159 ) );
  NOR2_X1 u2_u9_u1_U33 (.A1( u2_u9_u1_n168 ) , .A2( u2_u9_u1_n176 ) , .ZN( u2_u9_u1_n98 ) );
  AOI211_X1 u2_u9_u1_U34 (.B( u2_u9_u1_n162 ) , .A( u2_u9_u1_n163 ) , .C2( u2_u9_u1_n164 ) , .ZN( u2_u9_u1_n165 ) , .C1( u2_u9_u1_n171 ) );
  AOI21_X1 u2_u9_u1_U35 (.A( u2_u9_u1_n160 ) , .B2( u2_u9_u1_n161 ) , .ZN( u2_u9_u1_n162 ) , .B1( u2_u9_u1_n182 ) );
  OR2_X1 u2_u9_u1_U36 (.A2( u2_u9_u1_n157 ) , .A1( u2_u9_u1_n158 ) , .ZN( u2_u9_u1_n163 ) );
  NAND2_X1 u2_u9_u1_U37 (.A1( u2_u9_u1_n128 ) , .ZN( u2_u9_u1_n146 ) , .A2( u2_u9_u1_n160 ) );
  NAND2_X1 u2_u9_u1_U38 (.A2( u2_u9_u1_n112 ) , .ZN( u2_u9_u1_n139 ) , .A1( u2_u9_u1_n152 ) );
  NAND2_X1 u2_u9_u1_U39 (.A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n156 ) , .A2( u2_u9_u1_n99 ) );
  AOI221_X1 u2_u9_u1_U4 (.A( u2_u9_u1_n138 ) , .C2( u2_u9_u1_n139 ) , .C1( u2_u9_u1_n140 ) , .B2( u2_u9_u1_n141 ) , .ZN( u2_u9_u1_n142 ) , .B1( u2_u9_u1_n175 ) );
  AOI221_X1 u2_u9_u1_U40 (.B1( u2_u9_u1_n140 ) , .ZN( u2_u9_u1_n167 ) , .B2( u2_u9_u1_n172 ) , .C2( u2_u9_u1_n175 ) , .C1( u2_u9_u1_n178 ) , .A( u2_u9_u1_n188 ) );
  INV_X1 u2_u9_u1_U41 (.ZN( u2_u9_u1_n188 ) , .A( u2_u9_u1_n97 ) );
  AOI211_X1 u2_u9_u1_U42 (.A( u2_u9_u1_n118 ) , .C1( u2_u9_u1_n132 ) , .C2( u2_u9_u1_n139 ) , .B( u2_u9_u1_n96 ) , .ZN( u2_u9_u1_n97 ) );
  AOI21_X1 u2_u9_u1_U43 (.B2( u2_u9_u1_n121 ) , .B1( u2_u9_u1_n135 ) , .A( u2_u9_u1_n152 ) , .ZN( u2_u9_u1_n96 ) );
  NOR2_X1 u2_u9_u1_U44 (.ZN( u2_u9_u1_n117 ) , .A1( u2_u9_u1_n121 ) , .A2( u2_u9_u1_n160 ) );
  OAI21_X1 u2_u9_u1_U45 (.B2( u2_u9_u1_n123 ) , .ZN( u2_u9_u1_n145 ) , .B1( u2_u9_u1_n160 ) , .A( u2_u9_u1_n185 ) );
  INV_X1 u2_u9_u1_U46 (.A( u2_u9_u1_n122 ) , .ZN( u2_u9_u1_n185 ) );
  AOI21_X1 u2_u9_u1_U47 (.B2( u2_u9_u1_n120 ) , .B1( u2_u9_u1_n121 ) , .ZN( u2_u9_u1_n122 ) , .A( u2_u9_u1_n128 ) );
  AOI21_X1 u2_u9_u1_U48 (.A( u2_u9_u1_n128 ) , .B2( u2_u9_u1_n129 ) , .ZN( u2_u9_u1_n130 ) , .B1( u2_u9_u1_n150 ) );
  NAND2_X1 u2_u9_u1_U49 (.ZN( u2_u9_u1_n112 ) , .A1( u2_u9_u1_n169 ) , .A2( u2_u9_u1_n170 ) );
  AOI211_X1 u2_u9_u1_U5 (.ZN( u2_u9_u1_n124 ) , .A( u2_u9_u1_n138 ) , .C2( u2_u9_u1_n139 ) , .B( u2_u9_u1_n145 ) , .C1( u2_u9_u1_n147 ) );
  NAND2_X1 u2_u9_u1_U50 (.ZN( u2_u9_u1_n129 ) , .A2( u2_u9_u1_n95 ) , .A1( u2_u9_u1_n98 ) );
  NAND2_X1 u2_u9_u1_U51 (.A1( u2_u9_u1_n102 ) , .ZN( u2_u9_u1_n154 ) , .A2( u2_u9_u1_n99 ) );
  NAND2_X1 u2_u9_u1_U52 (.A2( u2_u9_u1_n100 ) , .ZN( u2_u9_u1_n135 ) , .A1( u2_u9_u1_n99 ) );
  AOI21_X1 u2_u9_u1_U53 (.A( u2_u9_u1_n152 ) , .B2( u2_u9_u1_n153 ) , .B1( u2_u9_u1_n154 ) , .ZN( u2_u9_u1_n158 ) );
  INV_X1 u2_u9_u1_U54 (.A( u2_u9_u1_n160 ) , .ZN( u2_u9_u1_n175 ) );
  NAND2_X1 u2_u9_u1_U55 (.A1( u2_u9_u1_n100 ) , .ZN( u2_u9_u1_n116 ) , .A2( u2_u9_u1_n95 ) );
  NAND2_X1 u2_u9_u1_U56 (.A1( u2_u9_u1_n102 ) , .ZN( u2_u9_u1_n131 ) , .A2( u2_u9_u1_n95 ) );
  NAND2_X1 u2_u9_u1_U57 (.A2( u2_u9_u1_n104 ) , .ZN( u2_u9_u1_n121 ) , .A1( u2_u9_u1_n98 ) );
  NAND2_X1 u2_u9_u1_U58 (.A1( u2_u9_u1_n103 ) , .ZN( u2_u9_u1_n153 ) , .A2( u2_u9_u1_n98 ) );
  NAND2_X1 u2_u9_u1_U59 (.A2( u2_u9_u1_n104 ) , .A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n133 ) );
  AOI22_X1 u2_u9_u1_U6 (.B2( u2_u9_u1_n136 ) , .A2( u2_u9_u1_n137 ) , .ZN( u2_u9_u1_n143 ) , .A1( u2_u9_u1_n171 ) , .B1( u2_u9_u1_n173 ) );
  NAND2_X1 u2_u9_u1_U60 (.ZN( u2_u9_u1_n150 ) , .A2( u2_u9_u1_n98 ) , .A1( u2_u9_u1_n99 ) );
  NAND2_X1 u2_u9_u1_U61 (.A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n155 ) , .A2( u2_u9_u1_n95 ) );
  OAI21_X1 u2_u9_u1_U62 (.ZN( u2_u9_u1_n109 ) , .B1( u2_u9_u1_n129 ) , .B2( u2_u9_u1_n160 ) , .A( u2_u9_u1_n167 ) );
  NAND2_X1 u2_u9_u1_U63 (.A2( u2_u9_u1_n100 ) , .A1( u2_u9_u1_n103 ) , .ZN( u2_u9_u1_n120 ) );
  NAND2_X1 u2_u9_u1_U64 (.A1( u2_u9_u1_n102 ) , .A2( u2_u9_u1_n104 ) , .ZN( u2_u9_u1_n115 ) );
  NAND2_X1 u2_u9_u1_U65 (.A2( u2_u9_u1_n100 ) , .A1( u2_u9_u1_n104 ) , .ZN( u2_u9_u1_n151 ) );
  NAND2_X1 u2_u9_u1_U66 (.A2( u2_u9_u1_n103 ) , .A1( u2_u9_u1_n105 ) , .ZN( u2_u9_u1_n161 ) );
  INV_X1 u2_u9_u1_U67 (.A( u2_u9_u1_n152 ) , .ZN( u2_u9_u1_n173 ) );
  INV_X1 u2_u9_u1_U68 (.A( u2_u9_u1_n128 ) , .ZN( u2_u9_u1_n172 ) );
  NAND2_X1 u2_u9_u1_U69 (.A2( u2_u9_u1_n102 ) , .A1( u2_u9_u1_n103 ) , .ZN( u2_u9_u1_n123 ) );
  INV_X1 u2_u9_u1_U7 (.A( u2_u9_u1_n147 ) , .ZN( u2_u9_u1_n181 ) );
  NOR2_X1 u2_u9_u1_U70 (.A2( u2_u9_X_7 ) , .A1( u2_u9_X_8 ) , .ZN( u2_u9_u1_n95 ) );
  NOR2_X1 u2_u9_u1_U71 (.A1( u2_u9_X_12 ) , .A2( u2_u9_X_9 ) , .ZN( u2_u9_u1_n100 ) );
  NOR2_X1 u2_u9_u1_U72 (.A2( u2_u9_X_8 ) , .A1( u2_u9_u1_n177 ) , .ZN( u2_u9_u1_n99 ) );
  NOR2_X1 u2_u9_u1_U73 (.A2( u2_u9_X_12 ) , .ZN( u2_u9_u1_n102 ) , .A1( u2_u9_u1_n176 ) );
  NOR2_X1 u2_u9_u1_U74 (.A2( u2_u9_X_9 ) , .ZN( u2_u9_u1_n105 ) , .A1( u2_u9_u1_n168 ) );
  NAND2_X1 u2_u9_u1_U75 (.A1( u2_u9_X_10 ) , .ZN( u2_u9_u1_n160 ) , .A2( u2_u9_u1_n169 ) );
  NAND2_X1 u2_u9_u1_U76 (.A2( u2_u9_X_10 ) , .A1( u2_u9_X_11 ) , .ZN( u2_u9_u1_n152 ) );
  NAND2_X1 u2_u9_u1_U77 (.A1( u2_u9_X_11 ) , .ZN( u2_u9_u1_n128 ) , .A2( u2_u9_u1_n170 ) );
  AND2_X1 u2_u9_u1_U78 (.A2( u2_u9_X_7 ) , .A1( u2_u9_X_8 ) , .ZN( u2_u9_u1_n104 ) );
  AND2_X1 u2_u9_u1_U79 (.A1( u2_u9_X_8 ) , .ZN( u2_u9_u1_n103 ) , .A2( u2_u9_u1_n177 ) );
  AOI22_X1 u2_u9_u1_U8 (.B2( u2_u9_u1_n113 ) , .A2( u2_u9_u1_n114 ) , .ZN( u2_u9_u1_n125 ) , .A1( u2_u9_u1_n171 ) , .B1( u2_u9_u1_n173 ) );
  INV_X1 u2_u9_u1_U80 (.A( u2_u9_X_10 ) , .ZN( u2_u9_u1_n170 ) );
  INV_X1 u2_u9_u1_U81 (.A( u2_u9_X_9 ) , .ZN( u2_u9_u1_n176 ) );
  INV_X1 u2_u9_u1_U82 (.A( u2_u9_X_11 ) , .ZN( u2_u9_u1_n169 ) );
  INV_X1 u2_u9_u1_U83 (.A( u2_u9_X_12 ) , .ZN( u2_u9_u1_n168 ) );
  INV_X1 u2_u9_u1_U84 (.A( u2_u9_X_7 ) , .ZN( u2_u9_u1_n177 ) );
  NAND4_X1 u2_u9_u1_U85 (.ZN( u2_out9_28 ) , .A4( u2_u9_u1_n124 ) , .A3( u2_u9_u1_n125 ) , .A2( u2_u9_u1_n126 ) , .A1( u2_u9_u1_n127 ) );
  OAI21_X1 u2_u9_u1_U86 (.ZN( u2_u9_u1_n127 ) , .B2( u2_u9_u1_n139 ) , .B1( u2_u9_u1_n175 ) , .A( u2_u9_u1_n183 ) );
  OAI21_X1 u2_u9_u1_U87 (.ZN( u2_u9_u1_n126 ) , .B2( u2_u9_u1_n140 ) , .A( u2_u9_u1_n146 ) , .B1( u2_u9_u1_n178 ) );
  NAND4_X1 u2_u9_u1_U88 (.ZN( u2_out9_18 ) , .A4( u2_u9_u1_n165 ) , .A3( u2_u9_u1_n166 ) , .A1( u2_u9_u1_n167 ) , .A2( u2_u9_u1_n186 ) );
  AOI22_X1 u2_u9_u1_U89 (.B2( u2_u9_u1_n146 ) , .B1( u2_u9_u1_n147 ) , .A2( u2_u9_u1_n148 ) , .ZN( u2_u9_u1_n166 ) , .A1( u2_u9_u1_n172 ) );
  NAND2_X1 u2_u9_u1_U9 (.ZN( u2_u9_u1_n114 ) , .A1( u2_u9_u1_n134 ) , .A2( u2_u9_u1_n156 ) );
  INV_X1 u2_u9_u1_U90 (.A( u2_u9_u1_n145 ) , .ZN( u2_u9_u1_n186 ) );
  NAND4_X1 u2_u9_u1_U91 (.ZN( u2_out9_2 ) , .A4( u2_u9_u1_n142 ) , .A3( u2_u9_u1_n143 ) , .A2( u2_u9_u1_n144 ) , .A1( u2_u9_u1_n179 ) );
  OAI21_X1 u2_u9_u1_U92 (.B2( u2_u9_u1_n132 ) , .ZN( u2_u9_u1_n144 ) , .A( u2_u9_u1_n146 ) , .B1( u2_u9_u1_n180 ) );
  INV_X1 u2_u9_u1_U93 (.A( u2_u9_u1_n130 ) , .ZN( u2_u9_u1_n179 ) );
  OR4_X1 u2_u9_u1_U94 (.ZN( u2_out9_13 ) , .A4( u2_u9_u1_n108 ) , .A3( u2_u9_u1_n109 ) , .A2( u2_u9_u1_n110 ) , .A1( u2_u9_u1_n111 ) );
  AOI21_X1 u2_u9_u1_U95 (.ZN( u2_u9_u1_n110 ) , .A( u2_u9_u1_n116 ) , .B1( u2_u9_u1_n152 ) , .B2( u2_u9_u1_n160 ) );
  AOI21_X1 u2_u9_u1_U96 (.ZN( u2_u9_u1_n111 ) , .A( u2_u9_u1_n128 ) , .B2( u2_u9_u1_n131 ) , .B1( u2_u9_u1_n135 ) );
  NAND3_X1 u2_u9_u1_U97 (.A3( u2_u9_u1_n149 ) , .A2( u2_u9_u1_n150 ) , .A1( u2_u9_u1_n151 ) , .ZN( u2_u9_u1_n164 ) );
  NAND3_X1 u2_u9_u1_U98 (.A3( u2_u9_u1_n134 ) , .A2( u2_u9_u1_n135 ) , .ZN( u2_u9_u1_n136 ) , .A1( u2_u9_u1_n151 ) );
  NAND3_X1 u2_u9_u1_U99 (.A1( u2_u9_u1_n133 ) , .ZN( u2_u9_u1_n137 ) , .A2( u2_u9_u1_n154 ) , .A3( u2_u9_u1_n181 ) );
  OAI22_X1 u2_u9_u2_U10 (.B1( u2_u9_u2_n151 ) , .A2( u2_u9_u2_n152 ) , .A1( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n160 ) , .B2( u2_u9_u2_n168 ) );
  NAND3_X1 u2_u9_u2_U100 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n104 ) , .A3( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n98 ) );
  NOR3_X1 u2_u9_u2_U11 (.A1( u2_u9_u2_n150 ) , .ZN( u2_u9_u2_n151 ) , .A3( u2_u9_u2_n175 ) , .A2( u2_u9_u2_n188 ) );
  AOI21_X1 u2_u9_u2_U12 (.B2( u2_u9_u2_n123 ) , .ZN( u2_u9_u2_n125 ) , .A( u2_u9_u2_n171 ) , .B1( u2_u9_u2_n184 ) );
  INV_X1 u2_u9_u2_U13 (.A( u2_u9_u2_n150 ) , .ZN( u2_u9_u2_n184 ) );
  AOI21_X1 u2_u9_u2_U14 (.ZN( u2_u9_u2_n144 ) , .B2( u2_u9_u2_n155 ) , .A( u2_u9_u2_n172 ) , .B1( u2_u9_u2_n185 ) );
  AOI21_X1 u2_u9_u2_U15 (.B2( u2_u9_u2_n143 ) , .ZN( u2_u9_u2_n145 ) , .B1( u2_u9_u2_n152 ) , .A( u2_u9_u2_n171 ) );
  INV_X1 u2_u9_u2_U16 (.A( u2_u9_u2_n156 ) , .ZN( u2_u9_u2_n171 ) );
  INV_X1 u2_u9_u2_U17 (.A( u2_u9_u2_n120 ) , .ZN( u2_u9_u2_n188 ) );
  NAND2_X1 u2_u9_u2_U18 (.A2( u2_u9_u2_n122 ) , .ZN( u2_u9_u2_n150 ) , .A1( u2_u9_u2_n152 ) );
  INV_X1 u2_u9_u2_U19 (.A( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n170 ) );
  INV_X1 u2_u9_u2_U20 (.A( u2_u9_u2_n137 ) , .ZN( u2_u9_u2_n173 ) );
  NAND2_X1 u2_u9_u2_U21 (.A1( u2_u9_u2_n132 ) , .A2( u2_u9_u2_n139 ) , .ZN( u2_u9_u2_n157 ) );
  INV_X1 u2_u9_u2_U22 (.A( u2_u9_u2_n113 ) , .ZN( u2_u9_u2_n178 ) );
  INV_X1 u2_u9_u2_U23 (.A( u2_u9_u2_n139 ) , .ZN( u2_u9_u2_n175 ) );
  INV_X1 u2_u9_u2_U24 (.A( u2_u9_u2_n155 ) , .ZN( u2_u9_u2_n181 ) );
  INV_X1 u2_u9_u2_U25 (.A( u2_u9_u2_n119 ) , .ZN( u2_u9_u2_n177 ) );
  INV_X1 u2_u9_u2_U26 (.A( u2_u9_u2_n116 ) , .ZN( u2_u9_u2_n180 ) );
  INV_X1 u2_u9_u2_U27 (.A( u2_u9_u2_n131 ) , .ZN( u2_u9_u2_n179 ) );
  INV_X1 u2_u9_u2_U28 (.A( u2_u9_u2_n154 ) , .ZN( u2_u9_u2_n176 ) );
  NAND2_X1 u2_u9_u2_U29 (.A2( u2_u9_u2_n116 ) , .A1( u2_u9_u2_n117 ) , .ZN( u2_u9_u2_n118 ) );
  NOR2_X1 u2_u9_u2_U3 (.ZN( u2_u9_u2_n121 ) , .A2( u2_u9_u2_n177 ) , .A1( u2_u9_u2_n180 ) );
  INV_X1 u2_u9_u2_U30 (.A( u2_u9_u2_n132 ) , .ZN( u2_u9_u2_n182 ) );
  INV_X1 u2_u9_u2_U31 (.A( u2_u9_u2_n158 ) , .ZN( u2_u9_u2_n183 ) );
  OAI21_X1 u2_u9_u2_U32 (.A( u2_u9_u2_n156 ) , .B1( u2_u9_u2_n157 ) , .ZN( u2_u9_u2_n158 ) , .B2( u2_u9_u2_n179 ) );
  NOR2_X1 u2_u9_u2_U33 (.ZN( u2_u9_u2_n156 ) , .A1( u2_u9_u2_n166 ) , .A2( u2_u9_u2_n169 ) );
  NOR2_X1 u2_u9_u2_U34 (.A2( u2_u9_u2_n114 ) , .ZN( u2_u9_u2_n137 ) , .A1( u2_u9_u2_n140 ) );
  NOR2_X1 u2_u9_u2_U35 (.A2( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n153 ) , .A1( u2_u9_u2_n156 ) );
  AOI211_X1 u2_u9_u2_U36 (.ZN( u2_u9_u2_n130 ) , .C1( u2_u9_u2_n138 ) , .C2( u2_u9_u2_n179 ) , .B( u2_u9_u2_n96 ) , .A( u2_u9_u2_n97 ) );
  OAI22_X1 u2_u9_u2_U37 (.B1( u2_u9_u2_n133 ) , .A2( u2_u9_u2_n137 ) , .A1( u2_u9_u2_n152 ) , .B2( u2_u9_u2_n168 ) , .ZN( u2_u9_u2_n97 ) );
  OAI221_X1 u2_u9_u2_U38 (.B1( u2_u9_u2_n113 ) , .C1( u2_u9_u2_n132 ) , .A( u2_u9_u2_n149 ) , .B2( u2_u9_u2_n171 ) , .C2( u2_u9_u2_n172 ) , .ZN( u2_u9_u2_n96 ) );
  OAI221_X1 u2_u9_u2_U39 (.A( u2_u9_u2_n115 ) , .C2( u2_u9_u2_n123 ) , .B2( u2_u9_u2_n143 ) , .B1( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n163 ) , .C1( u2_u9_u2_n168 ) );
  INV_X1 u2_u9_u2_U4 (.A( u2_u9_u2_n134 ) , .ZN( u2_u9_u2_n185 ) );
  OAI21_X1 u2_u9_u2_U40 (.A( u2_u9_u2_n114 ) , .ZN( u2_u9_u2_n115 ) , .B1( u2_u9_u2_n176 ) , .B2( u2_u9_u2_n178 ) );
  OAI221_X1 u2_u9_u2_U41 (.A( u2_u9_u2_n135 ) , .B2( u2_u9_u2_n136 ) , .B1( u2_u9_u2_n137 ) , .ZN( u2_u9_u2_n162 ) , .C2( u2_u9_u2_n167 ) , .C1( u2_u9_u2_n185 ) );
  AND3_X1 u2_u9_u2_U42 (.A3( u2_u9_u2_n131 ) , .A2( u2_u9_u2_n132 ) , .A1( u2_u9_u2_n133 ) , .ZN( u2_u9_u2_n136 ) );
  AOI22_X1 u2_u9_u2_U43 (.ZN( u2_u9_u2_n135 ) , .B1( u2_u9_u2_n140 ) , .A1( u2_u9_u2_n156 ) , .B2( u2_u9_u2_n180 ) , .A2( u2_u9_u2_n188 ) );
  AOI21_X1 u2_u9_u2_U44 (.ZN( u2_u9_u2_n149 ) , .B1( u2_u9_u2_n173 ) , .B2( u2_u9_u2_n188 ) , .A( u2_u9_u2_n95 ) );
  AND3_X1 u2_u9_u2_U45 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n104 ) , .A3( u2_u9_u2_n156 ) , .ZN( u2_u9_u2_n95 ) );
  OAI21_X1 u2_u9_u2_U46 (.A( u2_u9_u2_n141 ) , .B2( u2_u9_u2_n142 ) , .ZN( u2_u9_u2_n146 ) , .B1( u2_u9_u2_n153 ) );
  OAI21_X1 u2_u9_u2_U47 (.A( u2_u9_u2_n140 ) , .ZN( u2_u9_u2_n141 ) , .B1( u2_u9_u2_n176 ) , .B2( u2_u9_u2_n177 ) );
  NOR3_X1 u2_u9_u2_U48 (.ZN( u2_u9_u2_n142 ) , .A3( u2_u9_u2_n175 ) , .A2( u2_u9_u2_n178 ) , .A1( u2_u9_u2_n181 ) );
  OAI21_X1 u2_u9_u2_U49 (.A( u2_u9_u2_n101 ) , .B2( u2_u9_u2_n121 ) , .B1( u2_u9_u2_n153 ) , .ZN( u2_u9_u2_n164 ) );
  NOR4_X1 u2_u9_u2_U5 (.A4( u2_u9_u2_n124 ) , .A3( u2_u9_u2_n125 ) , .A2( u2_u9_u2_n126 ) , .A1( u2_u9_u2_n127 ) , .ZN( u2_u9_u2_n128 ) );
  NAND2_X1 u2_u9_u2_U50 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n107 ) , .ZN( u2_u9_u2_n155 ) );
  NAND2_X1 u2_u9_u2_U51 (.A2( u2_u9_u2_n105 ) , .A1( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n143 ) );
  NAND2_X1 u2_u9_u2_U52 (.A1( u2_u9_u2_n104 ) , .A2( u2_u9_u2_n106 ) , .ZN( u2_u9_u2_n152 ) );
  NAND2_X1 u2_u9_u2_U53 (.A1( u2_u9_u2_n100 ) , .A2( u2_u9_u2_n105 ) , .ZN( u2_u9_u2_n132 ) );
  INV_X1 u2_u9_u2_U54 (.A( u2_u9_u2_n140 ) , .ZN( u2_u9_u2_n168 ) );
  INV_X1 u2_u9_u2_U55 (.A( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n167 ) );
  NAND2_X1 u2_u9_u2_U56 (.A1( u2_u9_u2_n102 ) , .A2( u2_u9_u2_n106 ) , .ZN( u2_u9_u2_n113 ) );
  NAND2_X1 u2_u9_u2_U57 (.A1( u2_u9_u2_n106 ) , .A2( u2_u9_u2_n107 ) , .ZN( u2_u9_u2_n131 ) );
  NAND2_X1 u2_u9_u2_U58 (.A1( u2_u9_u2_n103 ) , .A2( u2_u9_u2_n107 ) , .ZN( u2_u9_u2_n139 ) );
  NAND2_X1 u2_u9_u2_U59 (.A1( u2_u9_u2_n103 ) , .A2( u2_u9_u2_n105 ) , .ZN( u2_u9_u2_n133 ) );
  AOI21_X1 u2_u9_u2_U6 (.B2( u2_u9_u2_n119 ) , .ZN( u2_u9_u2_n127 ) , .A( u2_u9_u2_n137 ) , .B1( u2_u9_u2_n155 ) );
  NAND2_X1 u2_u9_u2_U60 (.A1( u2_u9_u2_n102 ) , .A2( u2_u9_u2_n103 ) , .ZN( u2_u9_u2_n154 ) );
  NAND2_X1 u2_u9_u2_U61 (.A2( u2_u9_u2_n103 ) , .A1( u2_u9_u2_n104 ) , .ZN( u2_u9_u2_n119 ) );
  NAND2_X1 u2_u9_u2_U62 (.A2( u2_u9_u2_n107 ) , .A1( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n123 ) );
  NAND2_X1 u2_u9_u2_U63 (.A1( u2_u9_u2_n104 ) , .A2( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n122 ) );
  INV_X1 u2_u9_u2_U64 (.A( u2_u9_u2_n114 ) , .ZN( u2_u9_u2_n172 ) );
  NAND2_X1 u2_u9_u2_U65 (.A2( u2_u9_u2_n100 ) , .A1( u2_u9_u2_n102 ) , .ZN( u2_u9_u2_n116 ) );
  NAND2_X1 u2_u9_u2_U66 (.A1( u2_u9_u2_n102 ) , .A2( u2_u9_u2_n108 ) , .ZN( u2_u9_u2_n120 ) );
  NAND2_X1 u2_u9_u2_U67 (.A2( u2_u9_u2_n105 ) , .A1( u2_u9_u2_n106 ) , .ZN( u2_u9_u2_n117 ) );
  INV_X1 u2_u9_u2_U68 (.ZN( u2_u9_u2_n187 ) , .A( u2_u9_u2_n99 ) );
  OAI21_X1 u2_u9_u2_U69 (.B1( u2_u9_u2_n137 ) , .B2( u2_u9_u2_n143 ) , .A( u2_u9_u2_n98 ) , .ZN( u2_u9_u2_n99 ) );
  AOI21_X1 u2_u9_u2_U7 (.ZN( u2_u9_u2_n124 ) , .B1( u2_u9_u2_n131 ) , .B2( u2_u9_u2_n143 ) , .A( u2_u9_u2_n172 ) );
  NOR2_X1 u2_u9_u2_U70 (.A2( u2_u9_X_16 ) , .ZN( u2_u9_u2_n140 ) , .A1( u2_u9_u2_n166 ) );
  NOR2_X1 u2_u9_u2_U71 (.A2( u2_u9_X_13 ) , .A1( u2_u9_X_14 ) , .ZN( u2_u9_u2_n100 ) );
  NOR2_X1 u2_u9_u2_U72 (.A2( u2_u9_X_16 ) , .A1( u2_u9_X_17 ) , .ZN( u2_u9_u2_n138 ) );
  NOR2_X1 u2_u9_u2_U73 (.A2( u2_u9_X_15 ) , .A1( u2_u9_X_18 ) , .ZN( u2_u9_u2_n104 ) );
  NOR2_X1 u2_u9_u2_U74 (.A2( u2_u9_X_14 ) , .ZN( u2_u9_u2_n103 ) , .A1( u2_u9_u2_n174 ) );
  NOR2_X1 u2_u9_u2_U75 (.A2( u2_u9_X_15 ) , .ZN( u2_u9_u2_n102 ) , .A1( u2_u9_u2_n165 ) );
  NOR2_X1 u2_u9_u2_U76 (.A2( u2_u9_X_17 ) , .ZN( u2_u9_u2_n114 ) , .A1( u2_u9_u2_n169 ) );
  AND2_X1 u2_u9_u2_U77 (.A1( u2_u9_X_15 ) , .ZN( u2_u9_u2_n105 ) , .A2( u2_u9_u2_n165 ) );
  AND2_X1 u2_u9_u2_U78 (.A2( u2_u9_X_15 ) , .A1( u2_u9_X_18 ) , .ZN( u2_u9_u2_n107 ) );
  AND2_X1 u2_u9_u2_U79 (.A1( u2_u9_X_14 ) , .ZN( u2_u9_u2_n106 ) , .A2( u2_u9_u2_n174 ) );
  AOI21_X1 u2_u9_u2_U8 (.B2( u2_u9_u2_n120 ) , .B1( u2_u9_u2_n121 ) , .ZN( u2_u9_u2_n126 ) , .A( u2_u9_u2_n167 ) );
  AND2_X1 u2_u9_u2_U80 (.A1( u2_u9_X_13 ) , .A2( u2_u9_X_14 ) , .ZN( u2_u9_u2_n108 ) );
  INV_X1 u2_u9_u2_U81 (.A( u2_u9_X_16 ) , .ZN( u2_u9_u2_n169 ) );
  INV_X1 u2_u9_u2_U82 (.A( u2_u9_X_17 ) , .ZN( u2_u9_u2_n166 ) );
  INV_X1 u2_u9_u2_U83 (.A( u2_u9_X_13 ) , .ZN( u2_u9_u2_n174 ) );
  INV_X1 u2_u9_u2_U84 (.A( u2_u9_X_18 ) , .ZN( u2_u9_u2_n165 ) );
  NAND4_X1 u2_u9_u2_U85 (.ZN( u2_out9_30 ) , .A4( u2_u9_u2_n147 ) , .A3( u2_u9_u2_n148 ) , .A2( u2_u9_u2_n149 ) , .A1( u2_u9_u2_n187 ) );
  AOI21_X1 u2_u9_u2_U86 (.B2( u2_u9_u2_n138 ) , .ZN( u2_u9_u2_n148 ) , .A( u2_u9_u2_n162 ) , .B1( u2_u9_u2_n182 ) );
  NOR3_X1 u2_u9_u2_U87 (.A3( u2_u9_u2_n144 ) , .A2( u2_u9_u2_n145 ) , .A1( u2_u9_u2_n146 ) , .ZN( u2_u9_u2_n147 ) );
  NAND4_X1 u2_u9_u2_U88 (.ZN( u2_out9_24 ) , .A4( u2_u9_u2_n111 ) , .A3( u2_u9_u2_n112 ) , .A1( u2_u9_u2_n130 ) , .A2( u2_u9_u2_n187 ) );
  AOI221_X1 u2_u9_u2_U89 (.A( u2_u9_u2_n109 ) , .B1( u2_u9_u2_n110 ) , .ZN( u2_u9_u2_n111 ) , .C1( u2_u9_u2_n134 ) , .C2( u2_u9_u2_n170 ) , .B2( u2_u9_u2_n173 ) );
  OAI22_X1 u2_u9_u2_U9 (.ZN( u2_u9_u2_n109 ) , .A2( u2_u9_u2_n113 ) , .B2( u2_u9_u2_n133 ) , .B1( u2_u9_u2_n167 ) , .A1( u2_u9_u2_n168 ) );
  AOI21_X1 u2_u9_u2_U90 (.ZN( u2_u9_u2_n112 ) , .B2( u2_u9_u2_n156 ) , .A( u2_u9_u2_n164 ) , .B1( u2_u9_u2_n181 ) );
  NAND4_X1 u2_u9_u2_U91 (.ZN( u2_out9_16 ) , .A4( u2_u9_u2_n128 ) , .A3( u2_u9_u2_n129 ) , .A1( u2_u9_u2_n130 ) , .A2( u2_u9_u2_n186 ) );
  AOI22_X1 u2_u9_u2_U92 (.A2( u2_u9_u2_n118 ) , .ZN( u2_u9_u2_n129 ) , .A1( u2_u9_u2_n140 ) , .B1( u2_u9_u2_n157 ) , .B2( u2_u9_u2_n170 ) );
  INV_X1 u2_u9_u2_U93 (.A( u2_u9_u2_n163 ) , .ZN( u2_u9_u2_n186 ) );
  OR4_X1 u2_u9_u2_U94 (.ZN( u2_out9_6 ) , .A4( u2_u9_u2_n161 ) , .A3( u2_u9_u2_n162 ) , .A2( u2_u9_u2_n163 ) , .A1( u2_u9_u2_n164 ) );
  OR3_X1 u2_u9_u2_U95 (.A2( u2_u9_u2_n159 ) , .A1( u2_u9_u2_n160 ) , .ZN( u2_u9_u2_n161 ) , .A3( u2_u9_u2_n183 ) );
  AOI21_X1 u2_u9_u2_U96 (.B2( u2_u9_u2_n154 ) , .B1( u2_u9_u2_n155 ) , .ZN( u2_u9_u2_n159 ) , .A( u2_u9_u2_n167 ) );
  NAND3_X1 u2_u9_u2_U97 (.A2( u2_u9_u2_n117 ) , .A1( u2_u9_u2_n122 ) , .A3( u2_u9_u2_n123 ) , .ZN( u2_u9_u2_n134 ) );
  NAND3_X1 u2_u9_u2_U98 (.ZN( u2_u9_u2_n110 ) , .A2( u2_u9_u2_n131 ) , .A3( u2_u9_u2_n139 ) , .A1( u2_u9_u2_n154 ) );
  NAND3_X1 u2_u9_u2_U99 (.A2( u2_u9_u2_n100 ) , .ZN( u2_u9_u2_n101 ) , .A1( u2_u9_u2_n104 ) , .A3( u2_u9_u2_n114 ) );
  NAND2_X1 u2_uk_U1000 (.A1( u2_key_r_46 ) , .A2( u2_uk_n100 ) , .ZN( u2_uk_n969 ) );
  OAI21_X1 u2_uk_U1001 (.ZN( u2_K1_17 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1153 ) , .A( u2_uk_n971 ) );
  NAND2_X1 u2_uk_U1002 (.A1( u2_key_r_10 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n971 ) );
  OAI21_X1 u2_uk_U1017 (.ZN( u2_K10_13 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1605 ) , .A( u2_uk_n242 ) );
  NAND2_X1 u2_uk_U1018 (.A1( u2_uk_K_r8_48 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n242 ) );
  OAI21_X1 u2_uk_U1019 (.ZN( u2_K12_36 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1698 ) , .A( u2_uk_n472 ) );
  OAI21_X1 u2_uk_U1021 (.ZN( u2_K6_41 ) , .A( u2_uk_n1069 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1445 ) );
  NAND2_X1 u2_uk_U1028 (.A1( u2_uk_K_r5_16 ) , .ZN( u2_uk_n1087 ) , .A2( u2_uk_n17 ) );
  OAI21_X1 u2_uk_U1029 (.ZN( u2_K12_40 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1699 ) , .A( u2_uk_n501 ) );
  NAND2_X1 u2_uk_U1030 (.A1( u2_uk_K_r10_49 ) , .A2( u2_uk_n102 ) , .ZN( u2_uk_n501 ) );
  OAI21_X1 u2_uk_U1031 (.ZN( u2_K15_14 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1821 ) , .A( u2_uk_n936 ) );
  NAND2_X1 u2_uk_U1032 (.A1( u2_uk_K_r13_32 ) , .A2( u2_uk_n83 ) , .ZN( u2_uk_n936 ) );
  OAI22_X1 u2_uk_U104 (.ZN( u2_K2_5 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1244 ) , .A2( u2_uk_n1247 ) , .A1( u2_uk_n220 ) );
  NAND2_X1 u2_uk_U1042 (.A1( u2_uk_K_r9_0 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n366 ) );
  INV_X1 u2_uk_U1045 (.A( u2_key_r_6 ) , .ZN( u2_uk_n1146 ) );
  INV_X1 u2_uk_U1046 (.A( u2_key_r_54 ) , .ZN( u2_uk_n1185 ) );
  INV_X1 u2_uk_U1048 (.A( u2_key_r_26 ) , .ZN( u2_uk_n1161 ) );
  INV_X1 u2_uk_U1051 (.A( u2_key_r_34 ) , .ZN( u2_uk_n1168 ) );
  INV_X1 u2_uk_U1052 (.A( u2_key_r_27 ) , .ZN( u2_uk_n1162 ) );
  INV_X1 u2_uk_U1053 (.A( u2_key_r_24 ) , .ZN( u2_uk_n1159 ) );
  INV_X1 u2_uk_U1054 (.A( u2_key_r_20 ) , .ZN( u2_uk_n1155 ) );
  INV_X1 u2_uk_U1059 (.A( u2_key_r_13 ) , .ZN( u2_uk_n1150 ) );
  INV_X1 u2_uk_U1062 (.A( u2_key_r_19 ) , .ZN( u2_uk_n1154 ) );
  INV_X1 u2_uk_U1063 (.A( u2_key_r_4 ) , .ZN( u2_uk_n1145 ) );
  INV_X1 u2_uk_U1064 (.A( u2_key_r_17 ) , .ZN( u2_uk_n1153 ) );
  INV_X1 u2_uk_U1065 (.A( u2_key_r_53 ) , .ZN( u2_uk_n1184 ) );
  OAI21_X1 u2_uk_U1070 (.ZN( u2_K16_14 ) , .B2( u2_uk_n1205 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n951 ) );
  NAND2_X1 u2_uk_U1071 (.A1( u2_uk_K_r14_18 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n951 ) );
  INV_X1 u2_uk_U1082 (.ZN( u2_K2_10 ) , .A( u2_uk_n991 ) );
  AOI22_X1 u2_uk_U1083 (.B2( u2_uk_K_r0_34 ) , .A2( u2_uk_K_r0_55 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n147 ) , .ZN( u2_uk_n991 ) );
  INV_X1 u2_uk_U1084 (.ZN( u2_K1_11 ) , .A( u2_uk_n967 ) );
  INV_X1 u2_uk_U1086 (.ZN( u2_K1_18 ) , .A( u2_uk_n972 ) );
  INV_X1 u2_uk_U1090 (.ZN( u2_K7_6 ) , .A( u2_uk_n1095 ) );
  AOI22_X1 u2_uk_U1091 (.B2( u2_uk_K_r5_39 ) , .A2( u2_uk_K_r5_4 ) , .ZN( u2_uk_n1095 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n182 ) );
  INV_X1 u2_uk_U11 (.A( u2_uk_n163 ) , .ZN( u2_uk_n60 ) );
  INV_X1 u2_uk_U1108 (.ZN( u2_K2_7 ) , .A( u2_uk_n1004 ) );
  AOI22_X1 u2_uk_U1109 (.B2( u2_uk_K_r0_13 ) , .A2( u2_uk_K_r0_34 ) , .ZN( u2_uk_n1004 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U1110 (.ZN( u2_K12_32 ) , .A( u2_uk_n467 ) );
  INV_X1 u2_uk_U1116 (.ZN( u2_K7_13 ) , .A( u2_uk_n1076 ) );
  AOI22_X1 u2_uk_U1117 (.B2( u2_uk_K_r5_26 ) , .A2( u2_uk_K_r5_48 ) , .ZN( u2_uk_n1076 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n145 ) );
  INV_X1 u2_uk_U1132 (.ZN( u2_K10_12 ) , .A( u2_uk_n240 ) );
  OAI21_X1 u2_uk_U1140 (.ZN( u2_K16_2 ) , .B2( u2_uk_n1190 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n956 ) );
  OAI22_X1 u2_uk_U130 (.ZN( u2_K7_15 ) , .A2( u2_uk_n1454 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1494 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U137 (.ZN( u2_K6_19 ) , .A( u2_uk_n1061 ) , .B2( u2_uk_n1414 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U142 (.ZN( u2_K16_15 ) , .B2( u2_uk_n1206 ) , .A2( u2_uk_n1213 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U144 (.ZN( u2_K15_15 ) , .B2( u2_uk_n1843 ) , .B1( u2_uk_n188 ) , .A( u2_uk_n937 ) );
  NAND2_X1 u2_uk_U145 (.A1( u2_uk_K_r13_19 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n937 ) );
  OAI22_X1 u2_uk_U158 (.ZN( u2_K16_19 ) , .B2( u2_uk_n1190 ) , .A2( u2_uk_n1228 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U164 (.ZN( u2_K12_30 ) , .A( u2_uk_n456 ) );
  OAI21_X1 u2_uk_U168 (.ZN( u2_K1_14 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1160 ) , .A( u2_uk_n970 ) );
  INV_X1 u2_uk_U170 (.A( u2_key_r_25 ) , .ZN( u2_uk_n1160 ) );
  INV_X1 u2_uk_U18 (.ZN( u2_uk_n110 ) , .A( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U189 (.ZN( u2_K10_14 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1600 ) , .A2( u2_uk_n1631 ) , .B1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U199 (.ZN( u2_K15_24 ) , .A2( u2_uk_n1816 ) , .B2( u2_uk_n1834 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U215 (.ZN( u2_K12_31 ) , .B2( u2_uk_n1685 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n460 ) );
  NAND2_X1 u2_uk_U216 (.A1( u2_uk_K_r10_44 ) , .A2( u2_uk_n217 ) , .ZN( u2_uk_n460 ) );
  INV_X1 u2_uk_U217 (.ZN( u2_K11_31 ) , .A( u2_uk_n373 ) );
  INV_X1 u2_uk_U220 (.ZN( u2_K11_39 ) , .A( u2_uk_n379 ) );
  OAI22_X1 u2_uk_U227 (.ZN( u2_K6_31 ) , .B2( u2_uk_n1425 ) , .A2( u2_uk_n1430 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U240 (.ZN( u2_K12_39 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1690 ) , .A( u2_uk_n496 ) );
  NAND2_X1 u2_uk_U241 (.A1( u2_uk_K_r10_16 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n496 ) );
  INV_X1 u2_uk_U256 (.ZN( u2_K12_44 ) , .A( u2_uk_n504 ) );
  OAI22_X1 u2_uk_U258 (.ZN( u2_K12_48 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1691 ) , .A2( u2_uk_n1700 ) , .B1( u2_uk_n222 ) );
  BUF_X1 u2_uk_U27 (.Z( u2_uk_n129 ) , .A( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U277 (.ZN( u2_K15_6 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1834 ) , .A2( u2_uk_n1852 ) , .A1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U284 (.ZN( u2_K1_8 ) , .A2( u2_uk_n1146 ) , .B2( u2_uk_n1159 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U285 (.ZN( u2_K15_8 ) , .A( u2_uk_n946 ) );
  AOI22_X1 u2_uk_U286 (.B2( u2_uk_K_r13_13 ) , .A2( u2_uk_K_r13_17 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n141 ) , .ZN( u2_uk_n946 ) );
  INV_X1 u2_uk_U289 (.ZN( u2_K7_8 ) , .A( u2_uk_n1096 ) );
  BUF_X1 u2_uk_U29 (.Z( u2_uk_n147 ) , .A( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U295 (.ZN( u2_K2_8 ) , .A( u2_uk_n1005 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1240 ) );
  NAND2_X1 u2_uk_U296 (.A1( u2_uk_K_r0_17 ) , .ZN( u2_uk_n1005 ) , .A2( u2_uk_n93 ) );
  BUF_X1 u2_uk_U31 (.Z( u2_uk_n163 ) , .A( u2_uk_n209 ) );
  NAND2_X1 u2_uk_U312 (.A1( u2_uk_K_r11_7 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n656 ) );
  OAI22_X1 u2_uk_U331 (.ZN( u2_K15_4 ) , .B2( u2_uk_n1820 ) , .A2( u2_uk_n1850 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U343 (.ZN( u2_K2_4 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1238 ) , .A2( u2_uk_n1267 ) , .A1( u2_uk_n129 ) );
  OAI21_X1 u2_uk_U344 (.ZN( u2_K1_4 ) , .B2( u2_uk_n1184 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n990 ) );
  NAND2_X1 u2_uk_U345 (.A1( u2_key_r_3 ) , .A2( u2_uk_n207 ) , .ZN( u2_uk_n990 ) );
  OAI22_X1 u2_uk_U357 (.ZN( u2_K11_40 ) , .A1( u2_uk_n161 ) , .A2( u2_uk_n1634 ) , .B2( u2_uk_n1642 ) , .B1( u2_uk_n63 ) );
  BUF_X1 u2_uk_U36 (.Z( u2_uk_n188 ) , .A( u2_uk_n209 ) );
  INV_X1 u2_uk_U367 (.A( u2_key_r_8 ) , .ZN( u2_uk_n1148 ) );
  OAI22_X1 u2_uk_U377 (.ZN( u2_K12_28 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1680 ) , .A2( u2_uk_n1684 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U391 (.ZN( u2_K16_1 ) , .B2( u2_uk_n1218 ) , .A2( u2_uk_n1221 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n187 ) );
  OAI21_X1 u2_uk_U392 (.ZN( u2_K7_1 ) , .A( u2_uk_n1078 ) , .B2( u2_uk_n1462 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U393 (.A1( u2_uk_K_r5_10 ) , .ZN( u2_uk_n1078 ) , .A2( u2_uk_n129 ) );
  OAI21_X1 u2_uk_U396 (.ZN( u2_K10_16 ) , .B2( u2_uk_n1630 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n250 ) );
  NAND2_X1 u2_uk_U397 (.A1( u2_uk_K_r8_32 ) , .A2( u2_uk_n230 ) , .ZN( u2_uk_n250 ) );
  OAI21_X1 u2_uk_U400 (.ZN( u2_K7_16 ) , .A( u2_uk_n1077 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1496 ) );
  OAI21_X1 u2_uk_U407 (.ZN( u2_K15_9 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1843 ) , .A( u2_uk_n947 ) );
  INV_X1 u2_uk_U420 (.ZN( u2_K10_9 ) , .A( u2_uk_n308 ) );
  AOI22_X1 u2_uk_U421 (.B2( u2_uk_K_r8_17 ) , .A2( u2_uk_K_r8_27 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n308 ) );
  OAI22_X1 u2_uk_U426 (.ZN( u2_K7_9 ) , .B2( u2_uk_n1461 ) , .A2( u2_uk_n1468 ) , .A1( u2_uk_n231 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U430 (.ZN( u2_K2_9 ) , .A2( u2_uk_n1232 ) , .B2( u2_uk_n1261 ) , .B1( u2_uk_n145 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U434 (.ZN( u2_K16_16 ) , .B2( u2_uk_n1207 ) , .A2( u2_uk_n1214 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n17 ) );
  BUF_X1 u2_uk_U45 (.A( u2_uk_n203 ) , .Z( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U450 (.ZN( u2_K12_33 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1718 ) , .A( u2_uk_n468 ) );
  OAI22_X1 u2_uk_U455 (.ZN( u2_K11_33 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1653 ) , .A2( u2_uk_n1659 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U457 (.ZN( u2_K6_33 ) , .B2( u2_uk_n1428 ) , .A2( u2_uk_n1433 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U464 (.ZN( u2_K11_37 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1664 ) , .A( u2_uk_n377 ) );
  OAI21_X1 u2_uk_U468 (.ZN( u2_K6_37 ) , .A( u2_uk_n1068 ) , .B2( u2_uk_n1438 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U469 (.A1( u2_uk_K_r4_38 ) , .ZN( u2_uk_n1068 ) , .A2( u2_uk_n217 ) );
  NAND2_X1 u2_uk_U474 (.A1( u2_uk_K_r8_21 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n298 ) );
  BUF_X1 u2_uk_U48 (.Z( u2_uk_n191 ) , .A( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U503 (.ZN( u2_K7_2 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1086 ) , .B2( u2_uk_n1454 ) );
  NAND2_X1 u2_uk_U504 (.A1( u2_uk_K_r5_41 ) , .ZN( u2_uk_n1086 ) , .A2( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U507 (.ZN( u2_K1_12 ) , .B2( u2_uk_n1154 ) , .B1( u2_uk_n93 ) , .A( u2_uk_n968 ) );
  NAND2_X1 u2_uk_U508 (.A1( u2_key_r_12 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n968 ) );
  OAI22_X1 u2_uk_U516 (.ZN( u2_K7_17 ) , .B2( u2_uk_n1458 ) , .A2( u2_uk_n1488 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U521 (.ZN( u2_K15_12 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1815 ) , .B2( u2_uk_n1833 ) );
  INV_X1 u2_uk_U525 (.ZN( u2_K7_12 ) , .A( u2_uk_n1075 ) );
  AOI22_X1 u2_uk_U526 (.B2( u2_uk_K_r5_17 ) , .A2( u2_uk_K_r5_39 ) , .ZN( u2_uk_n1075 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U531 (.ZN( u2_K2_12 ) , .A2( u2_uk_n1233 ) , .B2( u2_uk_n1248 ) , .A1( u2_uk_n141 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U532 (.ZN( u2_K2_2 ) , .B2( u2_uk_n1243 ) , .A2( u2_uk_n1275 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U534 (.ZN( u2_K16_12 ) , .B2( u2_uk_n1198 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n949 ) );
  NAND2_X1 u2_uk_U535 (.A1( u2_uk_K_r14_12 ) , .A2( u2_uk_n145 ) , .ZN( u2_uk_n949 ) );
  OAI21_X1 u2_uk_U536 (.ZN( u2_K16_17 ) , .B2( u2_uk_n1197 ) , .B1( u2_uk_n188 ) , .A( u2_uk_n952 ) );
  NAND2_X1 u2_uk_U537 (.A1( u2_uk_K_r14_10 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n952 ) );
  OAI22_X1 u2_uk_U539 (.ZN( u2_K15_17 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1814 ) , .B2( u2_uk_n1832 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U54 (.ZN( u2_K11_34 ) , .A( u2_uk_n375 ) );
  INV_X1 u2_uk_U546 (.ZN( u2_K6_17 ) , .A( u2_uk_n1059 ) );
  AOI22_X1 u2_uk_U547 (.B2( u2_uk_K_r4_4 ) , .A2( u2_uk_K_r4_55 ) , .ZN( u2_uk_n1059 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n147 ) );
  AOI22_X1 u2_uk_U55 (.B2( u2_uk_K_r9_45 ) , .A2( u2_uk_K_r9_49 ) , .B1( u2_uk_n10 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n375 ) );
  OAI22_X1 u2_uk_U554 (.ZN( u2_K12_38 ) , .A1( u2_uk_n10 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1678 ) , .A2( u2_uk_n1705 ) );
  INV_X1 u2_uk_U559 (.ZN( u2_K11_36 ) , .A( u2_uk_n376 ) );
  OAI22_X1 u2_uk_U569 (.ZN( u2_K6_38 ) , .B2( u2_uk_n1418 ) , .A2( u2_uk_n1425 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U571 (.ZN( u2_K15_10 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1839 ) , .A( u2_uk_n934 ) );
  NAND2_X1 u2_uk_U572 (.A1( u2_uk_K_r13_55 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n934 ) );
  OAI22_X1 u2_uk_U578 (.ZN( u2_K16_10 ) , .B2( u2_uk_n1219 ) , .A2( u2_uk_n1222 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n217 ) );
  INV_X1 u2_uk_U584 (.ZN( u2_K1_10 ) , .A( u2_uk_n966 ) );
  AOI22_X1 u2_uk_U585 (.B2( u2_key_r_41 ) , .A2( u2_key_r_48 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n161 ) , .ZN( u2_uk_n966 ) );
  OAI22_X1 u2_uk_U588 (.ZN( u2_K16_22 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1205 ) , .A2( u2_uk_n1212 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U605 (.ZN( u2_K11_35 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1665 ) , .A2( u2_uk_n1673 ) , .A1( u2_uk_n93 ) );
  NAND2_X1 u2_uk_U608 (.A1( u2_uk_K_r5_37 ) , .ZN( u2_uk_n1090 ) , .A2( u2_uk_n11 ) );
  OAI22_X1 u2_uk_U611 (.ZN( u2_K12_35 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1698 ) , .A2( u2_uk_n1707 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U618 (.ZN( u2_K6_35 ) , .B2( u2_uk_n1439 ) , .A2( u2_uk_n1446 ) , .A1( u2_uk_n217 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U623 (.ZN( u2_K16_11 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1212 ) , .A( u2_uk_n948 ) );
  OAI22_X1 u2_uk_U625 (.ZN( u2_K7_11 ) , .B2( u2_uk_n1458 ) , .A2( u2_uk_n1475 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U626 (.ZN( u2_K15_11 ) , .B2( u2_uk_n1850 ) , .B1( u2_uk_n231 ) , .A( u2_uk_n935 ) );
  NAND2_X1 u2_uk_U627 (.A1( u2_uk_K_r13_25 ) , .A2( u2_uk_n207 ) , .ZN( u2_uk_n935 ) );
  OAI21_X1 u2_uk_U640 (.ZN( u2_K2_11 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1267 ) , .A( u2_uk_n992 ) );
  NAND2_X1 u2_uk_U641 (.A1( u2_uk_K_r0_25 ) , .A2( u2_uk_n100 ) , .ZN( u2_uk_n992 ) );
  OAI22_X1 u2_uk_U658 (.ZN( u2_K1_7 ) , .B2( u2_uk_n1155 ) , .A2( u2_uk_n1162 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U669 (.ZN( u2_K12_45 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1684 ) , .A( u2_uk_n509 ) );
  NAND2_X1 u2_uk_U670 (.A1( u2_uk_K_r10_43 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n509 ) );
  OAI22_X1 u2_uk_U676 (.ZN( u2_K16_3 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1198 ) , .A2( u2_uk_n1206 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U679 (.ZN( u2_K10_7 ) , .B2( u2_uk_n1604 ) , .A2( u2_uk_n1624 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U684 (.ZN( u2_K15_7 ) , .A1( u2_uk_n163 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1823 ) , .A2( u2_uk_n1839 ) );
  OAI22_X1 u2_uk_U687 (.ZN( u2_K16_7 ) , .B2( u2_uk_n1199 ) , .A2( u2_uk_n1207 ) , .A1( u2_uk_n141 ) , .B1( u2_uk_n17 ) );
  INV_X1 u2_uk_U7 (.ZN( u2_uk_n11 ) , .A( u2_uk_n141 ) );
  OAI22_X1 u2_uk_U70 (.ZN( u2_K16_23 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1213 ) , .A2( u2_uk_n1218 ) , .A1( u2_uk_n164 ) );
  OAI21_X1 u2_uk_U711 (.ZN( u2_K1_2 ) , .B2( u2_uk_n1145 ) , .B1( u2_uk_n220 ) , .A( u2_uk_n978 ) );
  NAND2_X1 u2_uk_U712 (.A1( u2_key_r_11 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n978 ) );
  OAI22_X1 u2_uk_U716 (.ZN( u2_K11_32 ) , .B2( u2_uk_n1640 ) , .A2( u2_uk_n1660 ) , .A1( u2_uk_n203 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U753 (.ZN( u2_K1_21 ) , .B2( u2_uk_n1153 ) , .A2( u2_uk_n1159 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U778 (.ZN( u2_K6_21 ) , .A( u2_uk_n1062 ) );
  AOI22_X1 u2_uk_U779 (.B2( u2_uk_K_r4_11 ) , .A2( u2_uk_K_r4_5 ) , .ZN( u2_uk_n1062 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U780 (.ZN( u2_K16_13 ) , .B2( u2_uk_n1227 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n950 ) );
  NAND2_X1 u2_uk_U781 (.A1( u2_uk_K_r14_46 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n950 ) );
  OAI22_X1 u2_uk_U802 (.ZN( u2_K7_18 ) , .A2( u2_uk_n1453 ) , .B2( u2_uk_n1466 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n31 ) );
  NAND2_X1 u2_uk_U806 (.A1( u2_uk_K_r6_46 ) , .ZN( u2_uk_n1102 ) , .A2( u2_uk_n17 ) );
  OAI21_X1 u2_uk_U808 (.ZN( u2_K16_18 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1229 ) , .A( u2_uk_n953 ) );
  NAND2_X1 u2_uk_U809 (.A1( u2_uk_K_r14_5 ) , .A2( u2_uk_n109 ) , .ZN( u2_uk_n953 ) );
  OAI22_X1 u2_uk_U810 (.ZN( u2_K10_18 ) , .A1( u2_uk_n110 ) , .A2( u2_uk_n1590 ) , .B2( u2_uk_n1604 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U817 (.ZN( u2_K16_20 ) , .B2( u2_uk_n1222 ) , .A2( u2_uk_n1229 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n209 ) );
  OAI21_X1 u2_uk_U82 (.ZN( u2_K11_41 ) , .B2( u2_uk_n1672 ) , .B1( u2_uk_n214 ) , .A( u2_uk_n382 ) );
  INV_X1 u2_uk_U822 (.ZN( u2_K6_18 ) , .A( u2_uk_n1060 ) );
  AOI22_X1 u2_uk_U823 (.B2( u2_uk_K_r4_11 ) , .A2( u2_uk_K_r4_17 ) , .A1( u2_uk_n100 ) , .ZN( u2_uk_n1060 ) , .B1( u2_uk_n155 ) );
  NAND2_X1 u2_uk_U83 (.A1( u2_uk_K_r9_31 ) , .A2( u2_uk_n203 ) , .ZN( u2_uk_n382 ) );
  OAI22_X1 u2_uk_U830 (.ZN( u2_K2_6 ) , .B2( u2_uk_n1249 ) , .A2( u2_uk_n1270 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U836 (.ZN( u2_K2_3 ) , .B2( u2_uk_n1239 ) , .A2( u2_uk_n1254 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U838 (.ZN( u2_K1_6 ) , .B2( u2_uk_n1168 ) , .A2( u2_uk_n1175 ) , .B1( u2_uk_n145 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U839 (.A( u2_key_r_41 ) , .ZN( u2_uk_n1175 ) );
  OAI22_X1 u2_uk_U849 (.ZN( u2_K15_22 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1828 ) , .A2( u2_uk_n1842 ) );
  OAI22_X1 u2_uk_U861 (.ZN( u2_K7_10 ) , .B2( u2_uk_n1457 ) , .A2( u2_uk_n1487 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U866 (.ZN( u2_K12_43 ) , .B2( u2_uk_n1687 ) , .A2( u2_uk_n1707 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U869 (.ZN( u2_K15_3 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1822 ) , .A2( u2_uk_n1838 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U875 (.ZN( u2_K7_14 ) , .B2( u2_uk_n1462 ) , .A2( u2_uk_n1497 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U885 (.ZN( u2_K16_21 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1197 ) , .A2( u2_uk_n1204 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U887 (.ZN( u2_K16_24 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1194 ) , .A2( u2_uk_n1199 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U900 (.ZN( u2_K6_42 ) , .B2( u2_uk_n1438 ) , .A2( u2_uk_n1445 ) , .A1( u2_uk_n163 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U901 (.ZN( u2_K6_39 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1411 ) , .B2( u2_uk_n1430 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U933 (.ZN( u2_K10_8 ) , .A2( u2_uk_n1591 ) , .B2( u2_uk_n1605 ) , .B1( u2_uk_n161 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U939 (.ZN( u2_K15_19 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1821 ) , .A2( u2_uk_n1851 ) , .B1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U967 (.ZN( u2_K1_3 ) , .B2( u2_uk_n1154 ) , .A2( u2_uk_n1161 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n207 ) );
  INV_X1 u2_uk_U970 (.ZN( u2_K12_42 ) , .A( u2_uk_n503 ) );
  OAI21_X1 u2_uk_U979 (.ZN( u2_K6_23 ) , .A( u2_uk_n1063 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1442 ) );
  OAI21_X1 u2_uk_U987 (.ZN( u2_K16_4 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1227 ) , .A( u2_uk_n965 ) );
  NAND2_X1 u2_uk_U988 (.A1( u2_uk_K_r14_3 ) , .A2( u2_uk_n92 ) , .ZN( u2_uk_n965 ) );
  OAI21_X1 u2_uk_U999 (.ZN( u2_K1_13 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1184 ) , .A( u2_uk_n969 ) );
endmodule

