module des_des_die_3 ( u0_K14_42, u0_K14_46, u0_K1_30, u0_K1_31, u0_K1_45, u0_K1_46, u0_K5_1, u0_K5_3, u0_K5_31, 
       u0_K5_32, u0_K5_34, u0_K5_38, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_L12_12, 
       u0_L12_15, u0_L12_21, u0_L12_22, u0_L12_27, u0_L12_32, u0_L12_5, u0_L12_7, u0_L3_11, u0_L3_12, 
       u0_L3_15, u0_L3_17, u0_L3_19, u0_L3_21, u0_L3_22, u0_L3_23, u0_L3_27, u0_L3_29, u0_L3_31, 
       u0_L3_32, u0_L3_4, u0_L3_5, u0_L3_7, u0_L3_9, u0_R12_1, u0_R12_24, u0_R12_25, u0_R12_26, 
       u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_30, u0_R12_31, u0_R12_32, u0_R3_1, u0_R3_2, u0_R3_20, 
       u0_R3_21, u0_R3_22, u0_R3_23, u0_R3_24, u0_R3_25, u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, 
       u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_desIn_r_0, u0_desIn_r_1, u0_desIn_r_11, 
       u0_desIn_r_16, u0_desIn_r_17, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_20, u0_desIn_r_22, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_28, 
       u0_desIn_r_3, u0_desIn_r_30, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_35, u0_desIn_r_38, u0_desIn_r_41, u0_desIn_r_42, 
       u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_49, u0_desIn_r_51, u0_desIn_r_52, u0_desIn_r_54, u0_desIn_r_56, u0_desIn_r_57, u0_desIn_r_59, 
       u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_1, u0_key_r_14, u0_key_r_16, u0_key_r_2, 
       u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, u0_key_r_31, u0_key_r_35, u0_key_r_36, 
       u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, u0_key_r_50, u0_key_r_51, u0_key_r_52, u0_key_r_7, u0_key_r_8, 
       u0_key_r_9, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_21, u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_16, u0_uk_K_r3_29, 
       u0_uk_K_r3_38, u0_uk_K_r3_52, u0_uk_K_r3_9, u0_uk_n10, u0_uk_n100, u0_uk_n109, u0_uk_n110, u0_uk_n117, u0_uk_n118, 
       u0_uk_n128, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n161, u0_uk_n163, u0_uk_n164, 
       u0_uk_n17, u0_uk_n182, u0_uk_n188, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n217, 
       u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
       u0_uk_n251, u0_uk_n252, u0_uk_n27, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n466, u0_uk_n471, u0_uk_n475, 
       u0_uk_n476, u0_uk_n482, u0_uk_n486, u0_uk_n488, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n52, 
       u0_uk_n56, u0_uk_n58, u0_uk_n59, u0_uk_n60, u0_uk_n65, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n77, 
       u0_uk_n805, u0_uk_n81, u0_uk_n810, u0_uk_n82, u0_uk_n875, u0_uk_n878, u0_uk_n90, u0_uk_n92, u0_uk_n93, 
       u0_uk_n99, u2_FP_36, u2_FP_37, u2_FP_38, u2_FP_39, u2_FP_40, u2_FP_41, u2_FP_42, u2_FP_43, 
       u2_FP_44, u2_FP_45, u2_FP_46, u2_FP_47, u2_FP_48, u2_FP_49, u2_K10_25, u2_K10_26, u2_K10_30, 
       u2_K10_32, u2_K10_34, u2_K10_36, u2_K10_42, u2_K11_13, u2_K11_16, u2_K11_18, u2_K11_38, u2_K11_42, 
       u2_K11_45, u2_K11_48, u2_K12_20, u2_K12_22, u2_K12_24, u2_K12_25, u2_K12_26, u2_K12_27, u2_K12_29, 
       u2_K12_34, u2_K12_37, u2_K12_41, u2_K12_46, u2_K12_47, u2_K13_14, u2_K13_20, u2_K13_26, u2_K13_3, 
       u2_K13_31, u2_K13_32, u2_K13_34, u2_K13_8, u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_20, u2_K15_21, 
       u2_K15_23, u2_K16_8, u2_K16_9, u2_K1_28, u2_K1_37, u2_K1_40, u2_K1_43, u2_K1_45, u2_K1_46, 
       u2_K2_16, u2_K2_18, u2_K2_20, u2_K3_30, u2_K4_38, u2_K4_39, u2_K4_42, u2_K4_6, u2_K4_7, 
       u2_K5_25, u2_K5_26, u2_K5_28, u2_K5_31, u2_K5_32, u2_K5_34, u2_K5_38, u2_K5_41, u2_K6_1, 
       u2_K6_11, u2_K6_3, u2_K6_32, u2_K6_34, u2_K6_36, u2_K6_40, u2_K7_31, u2_K7_33, u2_K7_35, 
       u2_K8_26, u2_K8_31, u2_K9_15, u2_K9_23, u2_K9_25, u2_K9_28, u2_K9_29, u2_K9_3, u2_K9_38, 
       u2_K9_40, u2_K9_45, u2_K9_5, u2_L0_1, u2_L0_10, u2_L0_13, u2_L0_16, u2_L0_18, u2_L0_2, 
       u2_L0_20, u2_L0_24, u2_L0_26, u2_L0_28, u2_L0_30, u2_L0_6, u2_L10_1, u2_L10_10, u2_L10_11, 
       u2_L10_12, u2_L10_14, u2_L10_15, u2_L10_19, u2_L10_20, u2_L10_21, u2_L10_22, u2_L10_25, u2_L10_26, 
       u2_L10_27, u2_L10_29, u2_L10_3, u2_L10_32, u2_L10_4, u2_L10_5, u2_L10_7, u2_L10_8, u2_L11_1, 
       u2_L11_10, u2_L11_11, u2_L11_13, u2_L11_14, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_19, u2_L11_2, 
       u2_L11_20, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, u2_L11_28, u2_L11_29, u2_L11_3, u2_L11_30, 
       u2_L11_31, u2_L11_4, u2_L11_6, u2_L11_8, u2_L11_9, u2_L13_1, u2_L13_10, u2_L13_15, u2_L13_16, 
       u2_L13_20, u2_L13_21, u2_L13_24, u2_L13_26, u2_L13_27, u2_L13_30, u2_L13_5, u2_L13_6, u2_L14_1, 
       u2_L14_10, u2_L14_13, u2_L14_16, u2_L14_18, u2_L14_2, u2_L14_20, u2_L14_24, u2_L14_26, u2_L14_28, 
       u2_L14_30, u2_L14_6, u2_L1_14, u2_L1_25, u2_L1_3, u2_L1_8, u2_L2_12, u2_L2_13, u2_L2_15, 
       u2_L2_17, u2_L2_18, u2_L2_2, u2_L2_21, u2_L2_22, u2_L2_23, u2_L2_27, u2_L2_28, u2_L2_31, 
       u2_L2_32, u2_L2_5, u2_L2_7, u2_L2_9, u2_L3_11, u2_L3_12, u2_L3_14, u2_L3_19, u2_L3_22, 
       u2_L3_25, u2_L3_29, u2_L3_3, u2_L3_32, u2_L3_4, u2_L3_7, u2_L3_8, u2_L4_11, u2_L4_12, 
       u2_L4_13, u2_L4_15, u2_L4_17, u2_L4_18, u2_L4_19, u2_L4_2, u2_L4_21, u2_L4_22, u2_L4_23, 
       u2_L4_27, u2_L4_28, u2_L4_29, u2_L4_31, u2_L4_32, u2_L4_4, u2_L4_5, u2_L4_7, u2_L4_9, 
       u2_L5_11, u2_L5_19, u2_L5_29, u2_L5_4, u2_L6_11, u2_L6_14, u2_L6_19, u2_L6_25, u2_L6_29, 
       u2_L6_3, u2_L6_4, u2_L6_8, u2_L7_1, u2_L7_10, u2_L7_12, u2_L7_13, u2_L7_14, u2_L7_15, 
       u2_L7_16, u2_L7_17, u2_L7_18, u2_L7_2, u2_L7_20, u2_L7_21, u2_L7_22, u2_L7_23, u2_L7_24, 
       u2_L7_25, u2_L7_26, u2_L7_27, u2_L7_28, u2_L7_3, u2_L7_30, u2_L7_31, u2_L7_32, u2_L7_5, 
       u2_L7_6, u2_L7_7, u2_L7_8, u2_L7_9, u2_L8_1, u2_L8_10, u2_L8_11, u2_L8_12, u2_L8_14, 
       u2_L8_19, u2_L8_20, u2_L8_22, u2_L8_25, u2_L8_26, u2_L8_29, u2_L8_3, u2_L8_32, u2_L8_4, 
       u2_L8_7, u2_L8_8, u2_L9_11, u2_L9_12, u2_L9_15, u2_L9_16, u2_L9_19, u2_L9_21, u2_L9_22, 
       u2_L9_24, u2_L9_27, u2_L9_29, u2_L9_30, u2_L9_32, u2_L9_4, u2_L9_5, u2_L9_6, u2_L9_7, 
       u2_R0_10, u2_R0_11, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_16, u2_R0_17, u2_R0_4, 
       u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_12, u2_R10_13, u2_R10_14, 
       u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_20, u2_R10_21, u2_R10_22, u2_R10_23, 
       u2_R10_24, u2_R10_25, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_29, u2_R10_30, u2_R10_31, u2_R10_32, 
       u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, u2_R11_17, 
       u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, u2_R11_25, 
       u2_R11_3, u2_R11_32, u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R13_1, 
       u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_14, u2_R13_15, u2_R13_16, u2_R13_17, u2_R13_28, 
       u2_R13_29, u2_R13_30, u2_R13_31, u2_R13_32, u2_R13_8, u2_R13_9, u2_R1_16, u2_R1_17, u2_R1_18, 
       u2_R1_19, u2_R1_20, u2_R1_21, u2_R2_1, u2_R2_2, u2_R2_24, u2_R2_25, u2_R2_26, u2_R2_27, 
       u2_R2_28, u2_R2_29, u2_R2_3, u2_R2_30, u2_R2_31, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, 
       u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_19, u2_R3_20, u2_R3_21, 
       u2_R3_22, u2_R3_23, u2_R3_24, u2_R3_25, u2_R3_26, u2_R3_27, u2_R3_28, u2_R3_29, u2_R4_1, 
       u2_R4_2, u2_R4_20, u2_R4_21, u2_R4_22, u2_R4_23, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_27, 
       u2_R4_28, u2_R4_29, u2_R4_3, u2_R4_30, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, 
       u2_R4_7, u2_R4_8, u2_R4_9, u2_R5_20, u2_R5_21, u2_R5_22, u2_R5_23, u2_R5_24, u2_R5_25, 
       u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_20, u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, 
       u2_R6_25, u2_R7_1, u2_R7_10, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
       u2_R7_17, u2_R7_18, u2_R7_19, u2_R7_2, u2_R7_20, u2_R7_21, u2_R7_24, u2_R7_25, u2_R7_26, 
       u2_R7_27, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_30, u2_R7_31, u2_R7_32, u2_R7_4, u2_R7_5, 
       u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_12, u2_R8_13, u2_R8_14, u2_R8_15, u2_R8_16, 
       u2_R8_17, u2_R8_18, u2_R8_19, u2_R8_20, u2_R8_21, u2_R8_22, u2_R8_23, u2_R8_24, u2_R8_25, 
       u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R9_1, u2_R9_10, u2_R9_11, u2_R9_12, u2_R9_13, 
       u2_R9_20, u2_R9_21, u2_R9_22, u2_R9_23, u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, 
       u2_R9_29, u2_R9_30, u2_R9_31, u2_R9_32, u2_R9_8, u2_R9_9, u2_desIn_r_0, u2_desIn_r_1, u2_desIn_r_11, 
       u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, u2_desIn_r_19, u2_desIn_r_20, u2_desIn_r_22, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_28, 
       u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_32, u2_desIn_r_33, u2_desIn_r_34, u2_desIn_r_35, u2_desIn_r_38, u2_desIn_r_41, u2_desIn_r_42, 
       u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_49, u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_54, u2_desIn_r_56, u2_desIn_r_57, u2_desIn_r_59, 
       u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_7, u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_2, u2_key_r_21, 
       u2_key_r_22, u2_key_r_23, u2_key_r_28, u2_key_r_29, u2_key_r_30, u2_key_r_31, u2_key_r_35, u2_key_r_36, u2_key_r_37, 
       u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_51, u2_key_r_52, u2_key_r_7, u2_key_r_9, u2_uk_K_r0_11, u2_uk_K_r0_13, 
       u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_32, u2_uk_K_r0_34, u2_uk_K_r0_47, u2_uk_K_r0_55, u2_uk_K_r10_16, u2_uk_K_r10_32, u2_uk_K_r10_41, 
       u2_uk_K_r10_43, u2_uk_K_r10_44, u2_uk_K_r10_49, u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, 
       u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, u2_uk_K_r11_28, u2_uk_K_r11_33, u2_uk_K_r11_39, u2_uk_K_r11_4, u2_uk_K_r11_47, u2_uk_K_r11_48, 
       u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r13_19, u2_uk_K_r13_32, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_18, u2_uk_K_r14_46, u2_uk_K_r14_5, 
       u2_uk_K_r1_42, u2_uk_K_r1_44, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_24, u2_uk_K_r2_25, u2_uk_K_r2_26, u2_uk_K_r2_50, u2_uk_K_r2_6, 
       u2_uk_K_r3_10, u2_uk_K_r3_14, u2_uk_K_r3_16, u2_uk_K_r3_29, u2_uk_K_r3_52, u2_uk_K_r3_9, u2_uk_K_r4_17, u2_uk_K_r4_3, u2_uk_K_r4_33, 
       u2_uk_K_r4_38, u2_uk_K_r4_41, u2_uk_K_r4_47, u2_uk_K_r4_54, u2_uk_K_r4_55, u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_21, u2_uk_K_r5_51, 
       u2_uk_K_r6_29, u2_uk_K_r6_51, u2_uk_K_r7_0, u2_uk_K_r7_13, u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_31, 
       u2_uk_K_r7_32, u2_uk_K_r7_37, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_46, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r7_9, u2_uk_K_r8_13, 
       u2_uk_K_r8_16, u2_uk_K_r8_19, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_28, u2_uk_K_r8_37, u2_uk_K_r8_40, u2_uk_K_r8_42, u2_uk_K_r8_43, 
       u2_uk_K_r8_44, u2_uk_K_r8_52, u2_uk_K_r8_8, u2_uk_K_r9_15, u2_uk_K_r9_23, u2_uk_K_r9_31, u2_uk_K_r9_33, u2_uk_K_r9_4, u2_uk_K_r9_45, 
       u2_uk_K_r9_49, u2_uk_K_r9_5, u2_uk_K_r9_55, u2_uk_n10, u2_uk_n100, u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, u2_uk_n1038, 
       u2_uk_n1040, u2_uk_n1046, u2_uk_n1049, u2_uk_n1069, u2_uk_n1070, u2_uk_n1073, u2_uk_n1074, u2_uk_n1089, u2_uk_n11, 
       u2_uk_n1104, u2_uk_n1107, u2_uk_n1119, u2_uk_n1120, u2_uk_n1121, u2_uk_n1125, u2_uk_n1128, u2_uk_n1130, u2_uk_n1131, 
       u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, u2_uk_n1141, u2_uk_n117, u2_uk_n118, u2_uk_n1190, u2_uk_n1194, 
       u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1212, u2_uk_n1213, 
       u2_uk_n1214, u2_uk_n1218, u2_uk_n1219, u2_uk_n1222, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, u2_uk_n1231, u2_uk_n1232, 
       u2_uk_n1233, u2_uk_n1234, u2_uk_n1238, u2_uk_n1240, u2_uk_n1243, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1260, 
       u2_uk_n1261, u2_uk_n1267, u2_uk_n1269, u2_uk_n1279, u2_uk_n1283, u2_uk_n129, u2_uk_n1298, u2_uk_n1299, u2_uk_n1303, 
       u2_uk_n1313, u2_uk_n1315, u2_uk_n1319, u2_uk_n1320, u2_uk_n1321, u2_uk_n1323, u2_uk_n1325, u2_uk_n1329, u2_uk_n1330, 
       u2_uk_n1331, u2_uk_n1333, u2_uk_n1336, u2_uk_n1337, u2_uk_n1339, u2_uk_n1341, u2_uk_n1342, u2_uk_n1344, u2_uk_n1345, 
       u2_uk_n1350, u2_uk_n1352, u2_uk_n1353, u2_uk_n1356, u2_uk_n1359, u2_uk_n1360, u2_uk_n1361, u2_uk_n1365, u2_uk_n1376, 
       u2_uk_n1377, u2_uk_n1378, u2_uk_n1382, u2_uk_n1383, u2_uk_n1395, u2_uk_n1396, u2_uk_n1400, u2_uk_n1401, u2_uk_n1403, 
       u2_uk_n1408, u2_uk_n141, u2_uk_n1410, u2_uk_n1411, u2_uk_n1413, u2_uk_n1416, u2_uk_n1418, u2_uk_n1419, u2_uk_n142, 
       u2_uk_n1422, u2_uk_n1424, u2_uk_n1425, u2_uk_n1426, u2_uk_n1428, u2_uk_n1429, u2_uk_n1430, u2_uk_n1433, u2_uk_n1435, 
       u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, u2_uk_n1444, u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1448, 
       u2_uk_n146, u2_uk_n1498, u2_uk_n1499, u2_uk_n1503, u2_uk_n1504, u2_uk_n1511, u2_uk_n1517, u2_uk_n1524, u2_uk_n1525, 
       u2_uk_n1526, u2_uk_n1530, u2_uk_n1532, u2_uk_n1533, u2_uk_n1538, u2_uk_n1543, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, 
       u2_uk_n1551, u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, u2_uk_n1568, u2_uk_n1570, u2_uk_n1571, 
       u2_uk_n1573, u2_uk_n1574, u2_uk_n1576, u2_uk_n1577, u2_uk_n1580, u2_uk_n1583, u2_uk_n1585, u2_uk_n1586, u2_uk_n1590, 
       u2_uk_n1594, u2_uk_n1597, u2_uk_n1599, u2_uk_n1602, u2_uk_n1603, u2_uk_n161, u2_uk_n1610, u2_uk_n1613, u2_uk_n1615, 
       u2_uk_n1617, u2_uk_n1622, u2_uk_n1625, u2_uk_n1629, u2_uk_n1630, u2_uk_n1632, u2_uk_n1634, u2_uk_n164, u2_uk_n1640, 
       u2_uk_n1642, u2_uk_n1646, u2_uk_n1653, u2_uk_n1659, u2_uk_n1660, u2_uk_n1661, u2_uk_n1664, u2_uk_n1665, u2_uk_n1672, 
       u2_uk_n1673, u2_uk_n1674, u2_uk_n1678, u2_uk_n1680, u2_uk_n1682, u2_uk_n1684, u2_uk_n1685, u2_uk_n1687, u2_uk_n1690, 
       u2_uk_n1691, u2_uk_n1698, u2_uk_n1699, u2_uk_n1700, u2_uk_n1705, u2_uk_n1707, u2_uk_n1718, u2_uk_n1720, u2_uk_n1723, 
       u2_uk_n1724, u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1735, u2_uk_n1736, 
       u2_uk_n1737, u2_uk_n1742, u2_uk_n1743, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, u2_uk_n1753, u2_uk_n1760, 
       u2_uk_n1763, u2_uk_n1767, u2_uk_n1814, u2_uk_n1816, u2_uk_n1818, u2_uk_n182, u2_uk_n1821, u2_uk_n1824, u2_uk_n1828, 
       u2_uk_n1832, u2_uk_n1834, u2_uk_n1836, u2_uk_n1837, u2_uk_n1842, u2_uk_n1843, u2_uk_n1845, u2_uk_n1851, u2_uk_n1854, 
       u2_uk_n1855, u2_uk_n1856, u2_uk_n187, u2_uk_n202, u2_uk_n208, u2_uk_n213, u2_uk_n220, u2_uk_n222, u2_uk_n238, 
       u2_uk_n257, u2_uk_n299, u2_uk_n31, u2_uk_n319, u2_uk_n373, u2_uk_n376, u2_uk_n377, u2_uk_n379, u2_uk_n385, 
       u2_uk_n443, u2_uk_n456, u2_uk_n467, u2_uk_n468, u2_uk_n472, u2_uk_n503, u2_uk_n504, u2_uk_n526, u2_uk_n551, 
       u2_uk_n586, u2_uk_n608, u2_uk_n665, u2_uk_n682, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n944, 
       u2_uk_n945, u2_uk_n948, u2_uk_n979, u2_uk_n984, u2_uk_n986, u2_uk_n994, u0_N10, u0_N11, u0_N13, u0_N131, u0_N132, u0_N134, u0_N136, u0_N138, u0_N139, 
        u0_N14, u0_N142, u0_N144, u0_N146, u0_N148, u0_N149, u0_N150, u0_N154, u0_N156, 
        u0_N158, u0_N159, u0_N18, u0_N2, u0_N20, u0_N21, u0_N24, u0_N26, u0_N28, 
        u0_N3, u0_N31, u0_N4, u0_N420, u0_N422, u0_N427, u0_N430, u0_N436, u0_N437, 
        u0_N442, u0_N447, u0_N6, u0_N7, u0_uk_n675, u0_uk_n687, u0_uk_n707, u0_uk_n711, u0_uk_n715, 
        u2_FP_1, u2_FP_10, u2_FP_13, u2_FP_16, u2_FP_18, u2_FP_2, u2_FP_20, u2_FP_24, u2_FP_26, 
        u2_FP_28, u2_FP_30, u2_FP_6, u2_N10, u2_N100, u2_N102, u2_N104, u2_N107, u2_N108, 
        u2_N11, u2_N110, u2_N112, u2_N113, u2_N116, u2_N117, u2_N118, u2_N122, u2_N123, 
        u2_N126, u2_N127, u2_N13, u2_N130, u2_N131, u2_N134, u2_N135, u2_N138, u2_N139, 
        u2_N14, u2_N141, u2_N146, u2_N149, u2_N152, u2_N156, u2_N159, u2_N161, u2_N163, 
        u2_N164, u2_N166, u2_N168, u2_N170, u2_N171, u2_N172, u2_N174, u2_N176, u2_N177, 
        u2_N178, u2_N18, u2_N180, u2_N181, u2_N182, u2_N186, u2_N187, u2_N188, u2_N190, 
        u2_N191, u2_N195, u2_N2, u2_N20, u2_N202, u2_N21, u2_N210, u2_N220, u2_N226, 
        u2_N227, u2_N231, u2_N234, u2_N237, u2_N24, u2_N242, u2_N248, u2_N252, u2_N256, 
        u2_N257, u2_N258, u2_N26, u2_N260, u2_N261, u2_N262, u2_N263, u2_N264, u2_N265, 
        u2_N267, u2_N268, u2_N269, u2_N270, u2_N271, u2_N272, u2_N273, u2_N275, u2_N276, 
        u2_N277, u2_N278, u2_N279, u2_N28, u2_N280, u2_N281, u2_N282, u2_N283, u2_N285, 
        u2_N286, u2_N287, u2_N288, u2_N290, u2_N291, u2_N294, u2_N295, u2_N297, u2_N298, 
        u2_N299, u2_N3, u2_N301, u2_N306, u2_N307, u2_N309, u2_N31, u2_N312, u2_N313, 
        u2_N316, u2_N319, u2_N32, u2_N323, u2_N324, u2_N325, u2_N326, u2_N33, u2_N330, 
        u2_N331, u2_N334, u2_N335, u2_N338, u2_N340, u2_N341, u2_N343, u2_N346, u2_N348, 
        u2_N349, u2_N351, u2_N352, u2_N354, u2_N355, u2_N356, u2_N358, u2_N359, u2_N361, 
        u2_N362, u2_N363, u2_N365, u2_N366, u2_N37, u2_N370, u2_N371, u2_N372, u2_N373, 
        u2_N376, u2_N377, u2_N378, u2_N380, u2_N383, u2_N384, u2_N385, u2_N386, u2_N387, 
        u2_N389, u2_N391, u2_N392, u2_N393, u2_N394, u2_N396, u2_N397, u2_N399, u2_N4, 
        u2_N400, u2_N401, u2_N402, u2_N403, u2_N406, u2_N407, u2_N408, u2_N409, u2_N41, 
        u2_N411, u2_N412, u2_N413, u2_N414, u2_N44, u2_N448, u2_N452, u2_N453, u2_N457, 
        u2_N462, u2_N463, u2_N467, u2_N468, u2_N47, u2_N471, u2_N473, u2_N474, u2_N477, 
        u2_N49, u2_N51, u2_N55, u2_N57, u2_N59, u2_N6, u2_N61, u2_N66, u2_N7, 
        u2_N71, u2_N77, u2_N88, u2_N97, u2_uk_n102, u2_uk_n1034, u2_uk_n1039, u2_uk_n1056, u2_uk_n109, 
        u2_uk_n110, u2_uk_n1142, u2_uk_n1144, u2_uk_n1149, u2_uk_n1152, u2_uk_n1171, u2_uk_n1178, u2_uk_n1183, u2_uk_n128, 
        u2_uk_n145, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n162, u2_uk_n163, u2_uk_n17, u2_uk_n188, u2_uk_n191, 
        u2_uk_n203, u2_uk_n207, u2_uk_n209, u2_uk_n214, u2_uk_n217, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, 
        u2_uk_n346, u2_uk_n395, u2_uk_n60, u2_uk_n605, u2_uk_n63, u2_uk_n672, u2_uk_n99 );
  input u0_K14_42, u0_K14_46, u0_K1_30, u0_K1_31, u0_K1_45, u0_K1_46, u0_K5_1, u0_K5_3, u0_K5_31, 
        u0_K5_32, u0_K5_34, u0_K5_38, u0_K5_4, u0_K5_41, u0_K5_44, u0_K5_47, u0_K5_48, u0_L12_12, 
        u0_L12_15, u0_L12_21, u0_L12_22, u0_L12_27, u0_L12_32, u0_L12_5, u0_L12_7, u0_L3_11, u0_L3_12, 
        u0_L3_15, u0_L3_17, u0_L3_19, u0_L3_21, u0_L3_22, u0_L3_23, u0_L3_27, u0_L3_29, u0_L3_31, 
        u0_L3_32, u0_L3_4, u0_L3_5, u0_L3_7, u0_L3_9, u0_R12_1, u0_R12_24, u0_R12_25, u0_R12_26, 
        u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_30, u0_R12_31, u0_R12_32, u0_R3_1, u0_R3_2, u0_R3_20, 
        u0_R3_21, u0_R3_22, u0_R3_23, u0_R3_24, u0_R3_25, u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, 
        u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_32, u0_R3_4, u0_R3_5, u0_desIn_r_0, u0_desIn_r_1, u0_desIn_r_11, 
        u0_desIn_r_16, u0_desIn_r_17, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_20, u0_desIn_r_22, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_28, 
        u0_desIn_r_3, u0_desIn_r_30, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_35, u0_desIn_r_38, u0_desIn_r_41, u0_desIn_r_42, 
        u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_49, u0_desIn_r_51, u0_desIn_r_52, u0_desIn_r_54, u0_desIn_r_56, u0_desIn_r_57, u0_desIn_r_59, 
        u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_1, u0_key_r_14, u0_key_r_16, u0_key_r_2, 
        u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, u0_key_r_31, u0_key_r_35, u0_key_r_36, 
        u0_key_r_37, u0_key_r_38, u0_key_r_42, u0_key_r_43, u0_key_r_50, u0_key_r_51, u0_key_r_52, u0_key_r_7, u0_key_r_8, 
        u0_key_r_9, u0_uk_K_r12_15, u0_uk_K_r12_16, u0_uk_K_r12_21, u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r3_15, u0_uk_K_r3_16, u0_uk_K_r3_29, 
        u0_uk_K_r3_38, u0_uk_K_r3_52, u0_uk_K_r3_9, u0_uk_n10, u0_uk_n100, u0_uk_n109, u0_uk_n110, u0_uk_n117, u0_uk_n118, 
        u0_uk_n128, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n161, u0_uk_n163, u0_uk_n164, 
        u0_uk_n17, u0_uk_n182, u0_uk_n188, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n213, u0_uk_n214, u0_uk_n217, 
        u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
        u0_uk_n251, u0_uk_n252, u0_uk_n27, u0_uk_n455, u0_uk_n457, u0_uk_n458, u0_uk_n466, u0_uk_n471, u0_uk_n475, 
        u0_uk_n476, u0_uk_n482, u0_uk_n486, u0_uk_n488, u0_uk_n490, u0_uk_n491, u0_uk_n493, u0_uk_n494, u0_uk_n52, 
        u0_uk_n56, u0_uk_n58, u0_uk_n59, u0_uk_n60, u0_uk_n65, u0_uk_n67, u0_uk_n68, u0_uk_n73, u0_uk_n77, 
        u0_uk_n805, u0_uk_n81, u0_uk_n810, u0_uk_n82, u0_uk_n875, u0_uk_n878, u0_uk_n90, u0_uk_n92, u0_uk_n93, 
        u0_uk_n99, u2_FP_36, u2_FP_37, u2_FP_38, u2_FP_39, u2_FP_40, u2_FP_41, u2_FP_42, u2_FP_43, 
        u2_FP_44, u2_FP_45, u2_FP_46, u2_FP_47, u2_FP_48, u2_FP_49, u2_K10_25, u2_K10_26, u2_K10_30, 
        u2_K10_32, u2_K10_34, u2_K10_36, u2_K10_42, u2_K11_13, u2_K11_16, u2_K11_18, u2_K11_38, u2_K11_42, 
        u2_K11_45, u2_K11_48, u2_K12_20, u2_K12_22, u2_K12_24, u2_K12_25, u2_K12_26, u2_K12_27, u2_K12_29, 
        u2_K12_34, u2_K12_37, u2_K12_41, u2_K12_46, u2_K12_47, u2_K13_14, u2_K13_20, u2_K13_26, u2_K13_3, 
        u2_K13_31, u2_K13_32, u2_K13_34, u2_K13_8, u2_K15_13, u2_K15_16, u2_K15_18, u2_K15_20, u2_K15_21, 
        u2_K15_23, u2_K16_8, u2_K16_9, u2_K1_28, u2_K1_37, u2_K1_40, u2_K1_43, u2_K1_45, u2_K1_46, 
        u2_K2_16, u2_K2_18, u2_K2_20, u2_K3_30, u2_K4_38, u2_K4_39, u2_K4_42, u2_K4_6, u2_K4_7, 
        u2_K5_25, u2_K5_26, u2_K5_28, u2_K5_31, u2_K5_32, u2_K5_34, u2_K5_38, u2_K5_41, u2_K6_1, 
        u2_K6_11, u2_K6_3, u2_K6_32, u2_K6_34, u2_K6_36, u2_K6_40, u2_K7_31, u2_K7_33, u2_K7_35, 
        u2_K8_26, u2_K8_31, u2_K9_15, u2_K9_23, u2_K9_25, u2_K9_28, u2_K9_29, u2_K9_3, u2_K9_38, 
        u2_K9_40, u2_K9_45, u2_K9_5, u2_L0_1, u2_L0_10, u2_L0_13, u2_L0_16, u2_L0_18, u2_L0_2, 
        u2_L0_20, u2_L0_24, u2_L0_26, u2_L0_28, u2_L0_30, u2_L0_6, u2_L10_1, u2_L10_10, u2_L10_11, 
        u2_L10_12, u2_L10_14, u2_L10_15, u2_L10_19, u2_L10_20, u2_L10_21, u2_L10_22, u2_L10_25, u2_L10_26, 
        u2_L10_27, u2_L10_29, u2_L10_3, u2_L10_32, u2_L10_4, u2_L10_5, u2_L10_7, u2_L10_8, u2_L11_1, 
        u2_L11_10, u2_L11_11, u2_L11_13, u2_L11_14, u2_L11_16, u2_L11_17, u2_L11_18, u2_L11_19, u2_L11_2, 
        u2_L11_20, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, u2_L11_28, u2_L11_29, u2_L11_3, u2_L11_30, 
        u2_L11_31, u2_L11_4, u2_L11_6, u2_L11_8, u2_L11_9, u2_L13_1, u2_L13_10, u2_L13_15, u2_L13_16, 
        u2_L13_20, u2_L13_21, u2_L13_24, u2_L13_26, u2_L13_27, u2_L13_30, u2_L13_5, u2_L13_6, u2_L14_1, 
        u2_L14_10, u2_L14_13, u2_L14_16, u2_L14_18, u2_L14_2, u2_L14_20, u2_L14_24, u2_L14_26, u2_L14_28, 
        u2_L14_30, u2_L14_6, u2_L1_14, u2_L1_25, u2_L1_3, u2_L1_8, u2_L2_12, u2_L2_13, u2_L2_15, 
        u2_L2_17, u2_L2_18, u2_L2_2, u2_L2_21, u2_L2_22, u2_L2_23, u2_L2_27, u2_L2_28, u2_L2_31, 
        u2_L2_32, u2_L2_5, u2_L2_7, u2_L2_9, u2_L3_11, u2_L3_12, u2_L3_14, u2_L3_19, u2_L3_22, 
        u2_L3_25, u2_L3_29, u2_L3_3, u2_L3_32, u2_L3_4, u2_L3_7, u2_L3_8, u2_L4_11, u2_L4_12, 
        u2_L4_13, u2_L4_15, u2_L4_17, u2_L4_18, u2_L4_19, u2_L4_2, u2_L4_21, u2_L4_22, u2_L4_23, 
        u2_L4_27, u2_L4_28, u2_L4_29, u2_L4_31, u2_L4_32, u2_L4_4, u2_L4_5, u2_L4_7, u2_L4_9, 
        u2_L5_11, u2_L5_19, u2_L5_29, u2_L5_4, u2_L6_11, u2_L6_14, u2_L6_19, u2_L6_25, u2_L6_29, 
        u2_L6_3, u2_L6_4, u2_L6_8, u2_L7_1, u2_L7_10, u2_L7_12, u2_L7_13, u2_L7_14, u2_L7_15, 
        u2_L7_16, u2_L7_17, u2_L7_18, u2_L7_2, u2_L7_20, u2_L7_21, u2_L7_22, u2_L7_23, u2_L7_24, 
        u2_L7_25, u2_L7_26, u2_L7_27, u2_L7_28, u2_L7_3, u2_L7_30, u2_L7_31, u2_L7_32, u2_L7_5, 
        u2_L7_6, u2_L7_7, u2_L7_8, u2_L7_9, u2_L8_1, u2_L8_10, u2_L8_11, u2_L8_12, u2_L8_14, 
        u2_L8_19, u2_L8_20, u2_L8_22, u2_L8_25, u2_L8_26, u2_L8_29, u2_L8_3, u2_L8_32, u2_L8_4, 
        u2_L8_7, u2_L8_8, u2_L9_11, u2_L9_12, u2_L9_15, u2_L9_16, u2_L9_19, u2_L9_21, u2_L9_22, 
        u2_L9_24, u2_L9_27, u2_L9_29, u2_L9_30, u2_L9_32, u2_L9_4, u2_L9_5, u2_L9_6, u2_L9_7, 
        u2_R0_10, u2_R0_11, u2_R0_12, u2_R0_13, u2_R0_14, u2_R0_15, u2_R0_16, u2_R0_17, u2_R0_4, 
        u2_R0_5, u2_R0_6, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_12, u2_R10_13, u2_R10_14, 
        u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_20, u2_R10_21, u2_R10_22, u2_R10_23, 
        u2_R10_24, u2_R10_25, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_29, u2_R10_30, u2_R10_31, u2_R10_32, 
        u2_R11_1, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, u2_R11_17, 
        u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_21, u2_R11_22, u2_R11_23, u2_R11_24, u2_R11_25, 
        u2_R11_3, u2_R11_32, u2_R11_4, u2_R11_5, u2_R11_6, u2_R11_7, u2_R11_8, u2_R11_9, u2_R13_1, 
        u2_R13_10, u2_R13_11, u2_R13_12, u2_R13_13, u2_R13_14, u2_R13_15, u2_R13_16, u2_R13_17, u2_R13_28, 
        u2_R13_29, u2_R13_30, u2_R13_31, u2_R13_32, u2_R13_8, u2_R13_9, u2_R1_16, u2_R1_17, u2_R1_18, 
        u2_R1_19, u2_R1_20, u2_R1_21, u2_R2_1, u2_R2_2, u2_R2_24, u2_R2_25, u2_R2_26, u2_R2_27, 
        u2_R2_28, u2_R2_29, u2_R2_3, u2_R2_30, u2_R2_31, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, 
        u2_R2_7, u2_R2_8, u2_R2_9, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_19, u2_R3_20, u2_R3_21, 
        u2_R3_22, u2_R3_23, u2_R3_24, u2_R3_25, u2_R3_26, u2_R3_27, u2_R3_28, u2_R3_29, u2_R4_1, 
        u2_R4_2, u2_R4_20, u2_R4_21, u2_R4_22, u2_R4_23, u2_R4_24, u2_R4_25, u2_R4_26, u2_R4_27, 
        u2_R4_28, u2_R4_29, u2_R4_3, u2_R4_30, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, 
        u2_R4_7, u2_R4_8, u2_R4_9, u2_R5_20, u2_R5_21, u2_R5_22, u2_R5_23, u2_R5_24, u2_R5_25, 
        u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_20, u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, 
        u2_R6_25, u2_R7_1, u2_R7_10, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, u2_R7_16, 
        u2_R7_17, u2_R7_18, u2_R7_19, u2_R7_2, u2_R7_20, u2_R7_21, u2_R7_24, u2_R7_25, u2_R7_26, 
        u2_R7_27, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_30, u2_R7_31, u2_R7_32, u2_R7_4, u2_R7_5, 
        u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_12, u2_R8_13, u2_R8_14, u2_R8_15, u2_R8_16, 
        u2_R8_17, u2_R8_18, u2_R8_19, u2_R8_20, u2_R8_21, u2_R8_22, u2_R8_23, u2_R8_24, u2_R8_25, 
        u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_R9_1, u2_R9_10, u2_R9_11, u2_R9_12, u2_R9_13, 
        u2_R9_20, u2_R9_21, u2_R9_22, u2_R9_23, u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, 
        u2_R9_29, u2_R9_30, u2_R9_31, u2_R9_32, u2_R9_8, u2_R9_9, u2_desIn_r_0, u2_desIn_r_1, u2_desIn_r_11, 
        u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, u2_desIn_r_19, u2_desIn_r_20, u2_desIn_r_22, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_28, 
        u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_32, u2_desIn_r_33, u2_desIn_r_34, u2_desIn_r_35, u2_desIn_r_38, u2_desIn_r_41, u2_desIn_r_42, 
        u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_49, u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_54, u2_desIn_r_56, u2_desIn_r_57, u2_desIn_r_59, 
        u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_7, u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_2, u2_key_r_21, 
        u2_key_r_22, u2_key_r_23, u2_key_r_28, u2_key_r_29, u2_key_r_30, u2_key_r_31, u2_key_r_35, u2_key_r_36, u2_key_r_37, 
        u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_51, u2_key_r_52, u2_key_r_7, u2_key_r_9, u2_uk_K_r0_11, u2_uk_K_r0_13, 
        u2_uk_K_r0_17, u2_uk_K_r0_25, u2_uk_K_r0_32, u2_uk_K_r0_34, u2_uk_K_r0_47, u2_uk_K_r0_55, u2_uk_K_r10_16, u2_uk_K_r10_32, u2_uk_K_r10_41, 
        u2_uk_K_r10_43, u2_uk_K_r10_44, u2_uk_K_r10_49, u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_19, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_24, 
        u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, u2_uk_K_r11_28, u2_uk_K_r11_33, u2_uk_K_r11_39, u2_uk_K_r11_4, u2_uk_K_r11_47, u2_uk_K_r11_48, 
        u2_uk_K_r11_53, u2_uk_K_r11_6, u2_uk_K_r13_19, u2_uk_K_r13_32, u2_uk_K_r14_10, u2_uk_K_r14_12, u2_uk_K_r14_18, u2_uk_K_r14_46, u2_uk_K_r14_5, 
        u2_uk_K_r1_42, u2_uk_K_r1_44, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_24, u2_uk_K_r2_25, u2_uk_K_r2_26, u2_uk_K_r2_50, u2_uk_K_r2_6, 
        u2_uk_K_r3_10, u2_uk_K_r3_14, u2_uk_K_r3_16, u2_uk_K_r3_29, u2_uk_K_r3_52, u2_uk_K_r3_9, u2_uk_K_r4_17, u2_uk_K_r4_3, u2_uk_K_r4_33, 
        u2_uk_K_r4_38, u2_uk_K_r4_41, u2_uk_K_r4_47, u2_uk_K_r4_54, u2_uk_K_r4_55, u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_21, u2_uk_K_r5_51, 
        u2_uk_K_r6_29, u2_uk_K_r6_51, u2_uk_K_r7_0, u2_uk_K_r7_13, u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_25, u2_uk_K_r7_26, u2_uk_K_r7_31, 
        u2_uk_K_r7_32, u2_uk_K_r7_37, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_46, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r7_9, u2_uk_K_r8_13, 
        u2_uk_K_r8_16, u2_uk_K_r8_19, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_28, u2_uk_K_r8_37, u2_uk_K_r8_40, u2_uk_K_r8_42, u2_uk_K_r8_43, 
        u2_uk_K_r8_44, u2_uk_K_r8_52, u2_uk_K_r8_8, u2_uk_K_r9_15, u2_uk_K_r9_23, u2_uk_K_r9_31, u2_uk_K_r9_33, u2_uk_K_r9_4, u2_uk_K_r9_45, 
        u2_uk_K_r9_49, u2_uk_K_r9_5, u2_uk_K_r9_55, u2_uk_n10, u2_uk_n100, u2_uk_n1031, u2_uk_n1035, u2_uk_n1036, u2_uk_n1038, 
        u2_uk_n1040, u2_uk_n1046, u2_uk_n1049, u2_uk_n1069, u2_uk_n1070, u2_uk_n1073, u2_uk_n1074, u2_uk_n1089, u2_uk_n11, 
        u2_uk_n1104, u2_uk_n1107, u2_uk_n1119, u2_uk_n1120, u2_uk_n1121, u2_uk_n1125, u2_uk_n1128, u2_uk_n1130, u2_uk_n1131, 
        u2_uk_n1134, u2_uk_n1136, u2_uk_n1137, u2_uk_n1140, u2_uk_n1141, u2_uk_n117, u2_uk_n118, u2_uk_n1190, u2_uk_n1194, 
        u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, u2_uk_n1207, u2_uk_n1212, u2_uk_n1213, 
        u2_uk_n1214, u2_uk_n1218, u2_uk_n1219, u2_uk_n1222, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, u2_uk_n1231, u2_uk_n1232, 
        u2_uk_n1233, u2_uk_n1234, u2_uk_n1238, u2_uk_n1240, u2_uk_n1243, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1260, 
        u2_uk_n1261, u2_uk_n1267, u2_uk_n1269, u2_uk_n1279, u2_uk_n1283, u2_uk_n129, u2_uk_n1298, u2_uk_n1299, u2_uk_n1303, 
        u2_uk_n1313, u2_uk_n1315, u2_uk_n1319, u2_uk_n1320, u2_uk_n1321, u2_uk_n1323, u2_uk_n1325, u2_uk_n1329, u2_uk_n1330, 
        u2_uk_n1331, u2_uk_n1333, u2_uk_n1336, u2_uk_n1337, u2_uk_n1339, u2_uk_n1341, u2_uk_n1342, u2_uk_n1344, u2_uk_n1345, 
        u2_uk_n1350, u2_uk_n1352, u2_uk_n1353, u2_uk_n1356, u2_uk_n1359, u2_uk_n1360, u2_uk_n1361, u2_uk_n1365, u2_uk_n1376, 
        u2_uk_n1377, u2_uk_n1378, u2_uk_n1382, u2_uk_n1383, u2_uk_n1395, u2_uk_n1396, u2_uk_n1400, u2_uk_n1401, u2_uk_n1403, 
        u2_uk_n1408, u2_uk_n141, u2_uk_n1410, u2_uk_n1411, u2_uk_n1413, u2_uk_n1416, u2_uk_n1418, u2_uk_n1419, u2_uk_n142, 
        u2_uk_n1422, u2_uk_n1424, u2_uk_n1425, u2_uk_n1426, u2_uk_n1428, u2_uk_n1429, u2_uk_n1430, u2_uk_n1433, u2_uk_n1435, 
        u2_uk_n1438, u2_uk_n1439, u2_uk_n1440, u2_uk_n1441, u2_uk_n1444, u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1448, 
        u2_uk_n146, u2_uk_n1498, u2_uk_n1499, u2_uk_n1503, u2_uk_n1504, u2_uk_n1511, u2_uk_n1517, u2_uk_n1524, u2_uk_n1525, 
        u2_uk_n1526, u2_uk_n1530, u2_uk_n1532, u2_uk_n1533, u2_uk_n1538, u2_uk_n1543, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, 
        u2_uk_n1551, u2_uk_n1555, u2_uk_n1556, u2_uk_n1558, u2_uk_n1563, u2_uk_n1565, u2_uk_n1568, u2_uk_n1570, u2_uk_n1571, 
        u2_uk_n1573, u2_uk_n1574, u2_uk_n1576, u2_uk_n1577, u2_uk_n1580, u2_uk_n1583, u2_uk_n1585, u2_uk_n1586, u2_uk_n1590, 
        u2_uk_n1594, u2_uk_n1597, u2_uk_n1599, u2_uk_n1602, u2_uk_n1603, u2_uk_n161, u2_uk_n1610, u2_uk_n1613, u2_uk_n1615, 
        u2_uk_n1617, u2_uk_n1622, u2_uk_n1625, u2_uk_n1629, u2_uk_n1630, u2_uk_n1632, u2_uk_n1634, u2_uk_n164, u2_uk_n1640, 
        u2_uk_n1642, u2_uk_n1646, u2_uk_n1653, u2_uk_n1659, u2_uk_n1660, u2_uk_n1661, u2_uk_n1664, u2_uk_n1665, u2_uk_n1672, 
        u2_uk_n1673, u2_uk_n1674, u2_uk_n1678, u2_uk_n1680, u2_uk_n1682, u2_uk_n1684, u2_uk_n1685, u2_uk_n1687, u2_uk_n1690, 
        u2_uk_n1691, u2_uk_n1698, u2_uk_n1699, u2_uk_n1700, u2_uk_n1705, u2_uk_n1707, u2_uk_n1718, u2_uk_n1720, u2_uk_n1723, 
        u2_uk_n1724, u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1734, u2_uk_n1735, u2_uk_n1736, 
        u2_uk_n1737, u2_uk_n1742, u2_uk_n1743, u2_uk_n1745, u2_uk_n1746, u2_uk_n1747, u2_uk_n1750, u2_uk_n1753, u2_uk_n1760, 
        u2_uk_n1763, u2_uk_n1767, u2_uk_n1814, u2_uk_n1816, u2_uk_n1818, u2_uk_n182, u2_uk_n1821, u2_uk_n1824, u2_uk_n1828, 
        u2_uk_n1832, u2_uk_n1834, u2_uk_n1836, u2_uk_n1837, u2_uk_n1842, u2_uk_n1843, u2_uk_n1845, u2_uk_n1851, u2_uk_n1854, 
        u2_uk_n1855, u2_uk_n1856, u2_uk_n187, u2_uk_n202, u2_uk_n208, u2_uk_n213, u2_uk_n220, u2_uk_n222, u2_uk_n238, 
        u2_uk_n257, u2_uk_n299, u2_uk_n31, u2_uk_n319, u2_uk_n373, u2_uk_n376, u2_uk_n377, u2_uk_n379, u2_uk_n385, 
        u2_uk_n443, u2_uk_n456, u2_uk_n467, u2_uk_n468, u2_uk_n472, u2_uk_n503, u2_uk_n504, u2_uk_n526, u2_uk_n551, 
        u2_uk_n586, u2_uk_n608, u2_uk_n665, u2_uk_n682, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n944, 
        u2_uk_n945, u2_uk_n948, u2_uk_n979, u2_uk_n984, u2_uk_n986, u2_uk_n994;
  output u0_N10, u0_N11, u0_N13, u0_N131, u0_N132, u0_N134, u0_N136, u0_N138, u0_N139, 
        u0_N14, u0_N142, u0_N144, u0_N146, u0_N148, u0_N149, u0_N150, u0_N154, u0_N156, 
        u0_N158, u0_N159, u0_N18, u0_N2, u0_N20, u0_N21, u0_N24, u0_N26, u0_N28, 
        u0_N3, u0_N31, u0_N4, u0_N420, u0_N422, u0_N427, u0_N430, u0_N436, u0_N437, 
        u0_N442, u0_N447, u0_N6, u0_N7, u0_uk_n675, u0_uk_n687, u0_uk_n707, u0_uk_n711, u0_uk_n715, 
        u2_FP_1, u2_FP_10, u2_FP_13, u2_FP_16, u2_FP_18, u2_FP_2, u2_FP_20, u2_FP_24, u2_FP_26, 
        u2_FP_28, u2_FP_30, u2_FP_6, u2_N10, u2_N100, u2_N102, u2_N104, u2_N107, u2_N108, 
        u2_N11, u2_N110, u2_N112, u2_N113, u2_N116, u2_N117, u2_N118, u2_N122, u2_N123, 
        u2_N126, u2_N127, u2_N13, u2_N130, u2_N131, u2_N134, u2_N135, u2_N138, u2_N139, 
        u2_N14, u2_N141, u2_N146, u2_N149, u2_N152, u2_N156, u2_N159, u2_N161, u2_N163, 
        u2_N164, u2_N166, u2_N168, u2_N170, u2_N171, u2_N172, u2_N174, u2_N176, u2_N177, 
        u2_N178, u2_N18, u2_N180, u2_N181, u2_N182, u2_N186, u2_N187, u2_N188, u2_N190, 
        u2_N191, u2_N195, u2_N2, u2_N20, u2_N202, u2_N21, u2_N210, u2_N220, u2_N226, 
        u2_N227, u2_N231, u2_N234, u2_N237, u2_N24, u2_N242, u2_N248, u2_N252, u2_N256, 
        u2_N257, u2_N258, u2_N26, u2_N260, u2_N261, u2_N262, u2_N263, u2_N264, u2_N265, 
        u2_N267, u2_N268, u2_N269, u2_N270, u2_N271, u2_N272, u2_N273, u2_N275, u2_N276, 
        u2_N277, u2_N278, u2_N279, u2_N28, u2_N280, u2_N281, u2_N282, u2_N283, u2_N285, 
        u2_N286, u2_N287, u2_N288, u2_N290, u2_N291, u2_N294, u2_N295, u2_N297, u2_N298, 
        u2_N299, u2_N3, u2_N301, u2_N306, u2_N307, u2_N309, u2_N31, u2_N312, u2_N313, 
        u2_N316, u2_N319, u2_N32, u2_N323, u2_N324, u2_N325, u2_N326, u2_N33, u2_N330, 
        u2_N331, u2_N334, u2_N335, u2_N338, u2_N340, u2_N341, u2_N343, u2_N346, u2_N348, 
        u2_N349, u2_N351, u2_N352, u2_N354, u2_N355, u2_N356, u2_N358, u2_N359, u2_N361, 
        u2_N362, u2_N363, u2_N365, u2_N366, u2_N37, u2_N370, u2_N371, u2_N372, u2_N373, 
        u2_N376, u2_N377, u2_N378, u2_N380, u2_N383, u2_N384, u2_N385, u2_N386, u2_N387, 
        u2_N389, u2_N391, u2_N392, u2_N393, u2_N394, u2_N396, u2_N397, u2_N399, u2_N4, 
        u2_N400, u2_N401, u2_N402, u2_N403, u2_N406, u2_N407, u2_N408, u2_N409, u2_N41, 
        u2_N411, u2_N412, u2_N413, u2_N414, u2_N44, u2_N448, u2_N452, u2_N453, u2_N457, 
        u2_N462, u2_N463, u2_N467, u2_N468, u2_N47, u2_N471, u2_N473, u2_N474, u2_N477, 
        u2_N49, u2_N51, u2_N55, u2_N57, u2_N59, u2_N6, u2_N61, u2_N66, u2_N7, 
        u2_N71, u2_N77, u2_N88, u2_N97, u2_uk_n102, u2_uk_n1034, u2_uk_n1039, u2_uk_n1056, u2_uk_n109, 
        u2_uk_n110, u2_uk_n1142, u2_uk_n1144, u2_uk_n1149, u2_uk_n1152, u2_uk_n1171, u2_uk_n1178, u2_uk_n1183, u2_uk_n128, 
        u2_uk_n145, u2_uk_n147, u2_uk_n148, u2_uk_n155, u2_uk_n162, u2_uk_n163, u2_uk_n17, u2_uk_n188, u2_uk_n191, 
        u2_uk_n203, u2_uk_n207, u2_uk_n209, u2_uk_n214, u2_uk_n217, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, 
        u2_uk_n346, u2_uk_n395, u2_uk_n60, u2_uk_n605, u2_uk_n63, u2_uk_n672, u2_uk_n99;
  wire u0_K14_37, u0_K14_38, u0_K14_39, u0_K14_40, u0_K14_41, u0_K14_43, u0_K14_44, u0_K14_45, u0_K14_47, 
       u0_K14_48, u0_K1_25, u0_K1_26, u0_K1_27, u0_K1_28, u0_K1_29, u0_K1_32, u0_K1_33, u0_K1_34, 
       u0_K1_35, u0_K1_36, u0_K1_37, u0_K1_38, u0_K1_39, u0_K1_40, u0_K1_41, u0_K1_42, u0_K1_43, 
       u0_K1_44, u0_K1_47, u0_K1_48, u0_K5_2, u0_K5_33, u0_K5_35, u0_K5_36, u0_K5_37, u0_K5_39, 
       u0_K5_40, u0_K5_42, u0_K5_43, u0_K5_45, u0_K5_46, u0_K5_5, u0_K5_6, u0_out0_11, u0_out0_12, 
       u0_out0_14, u0_out0_15, u0_out0_19, u0_out0_21, u0_out0_22, u0_out0_25, u0_out0_27, u0_out0_29, u0_out0_3, 
       u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_7, u0_out0_8, u0_out13_12, u0_out13_15, u0_out13_21, u0_out13_22, 
       u0_out13_27, u0_out13_32, u0_out13_5, u0_out13_7, u0_out4_11, u0_out4_12, u0_out4_15, u0_out4_17, u0_out4_19, 
       u0_out4_21, u0_out4_22, u0_out4_23, u0_out4_27, u0_out4_29, u0_out4_31, u0_out4_32, u0_out4_4, u0_out4_5, 
       u0_out4_7, u0_out4_9, u0_u0_X_25, u0_u0_X_26, u0_u0_X_27, u0_u0_X_28, u0_u0_X_29, u0_u0_X_30, u0_u0_X_31, 
       u0_u0_X_32, u0_u0_X_33, u0_u0_X_34, u0_u0_X_35, u0_u0_X_36, u0_u0_X_37, u0_u0_X_38, u0_u0_X_39, u0_u0_X_40, 
       u0_u0_X_41, u0_u0_X_42, u0_u0_X_43, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u0_X_47, u0_u0_X_48, u0_u0_u4_n1, 
       u0_u0_u4_n10, u0_u0_u4_n11, u0_u0_u4_n12, u0_u0_u4_n13, u0_u0_u4_n14, u0_u0_u4_n15, u0_u0_u4_n16, u0_u0_u4_n17, u0_u0_u4_n18, 
       u0_u0_u4_n19, u0_u0_u4_n2, u0_u0_u4_n20, u0_u0_u4_n21, u0_u0_u4_n22, u0_u0_u4_n23, u0_u0_u4_n24, u0_u0_u4_n25, u0_u0_u4_n26, 
       u0_u0_u4_n27, u0_u0_u4_n28, u0_u0_u4_n29, u0_u0_u4_n3, u0_u0_u4_n30, u0_u0_u4_n31, u0_u0_u4_n32, u0_u0_u4_n33, u0_u0_u4_n34, 
       u0_u0_u4_n35, u0_u0_u4_n36, u0_u0_u4_n37, u0_u0_u4_n38, u0_u0_u4_n39, u0_u0_u4_n4, u0_u0_u4_n40, u0_u0_u4_n41, u0_u0_u4_n42, 
       u0_u0_u4_n43, u0_u0_u4_n44, u0_u0_u4_n45, u0_u0_u4_n46, u0_u0_u4_n47, u0_u0_u4_n48, u0_u0_u4_n49, u0_u0_u4_n5, u0_u0_u4_n50, 
       u0_u0_u4_n51, u0_u0_u4_n52, u0_u0_u4_n53, u0_u0_u4_n54, u0_u0_u4_n55, u0_u0_u4_n56, u0_u0_u4_n57, u0_u0_u4_n58, u0_u0_u4_n59, 
       u0_u0_u4_n6, u0_u0_u4_n60, u0_u0_u4_n61, u0_u0_u4_n62, u0_u0_u4_n63, u0_u0_u4_n64, u0_u0_u4_n65, u0_u0_u4_n66, u0_u0_u4_n67, 
       u0_u0_u4_n68, u0_u0_u4_n69, u0_u0_u4_n7, u0_u0_u4_n70, u0_u0_u4_n71, u0_u0_u4_n72, u0_u0_u4_n73, u0_u0_u4_n74, u0_u0_u4_n75, 
       u0_u0_u4_n76, u0_u0_u4_n77, u0_u0_u4_n78, u0_u0_u4_n79, u0_u0_u4_n8, u0_u0_u4_n80, u0_u0_u4_n81, u0_u0_u4_n82, u0_u0_u4_n83, 
       u0_u0_u4_n84, u0_u0_u4_n85, u0_u0_u4_n86, u0_u0_u4_n87, u0_u0_u4_n88, u0_u0_u4_n89, u0_u0_u4_n9, u0_u0_u4_n90, u0_u0_u4_n91, 
       u0_u0_u4_n92, u0_u0_u4_n93, u0_u0_u5_n1, u0_u0_u5_n10, u0_u0_u5_n11, u0_u0_u5_n12, u0_u0_u5_n13, u0_u0_u5_n14, u0_u0_u5_n15, 
       u0_u0_u5_n16, u0_u0_u5_n17, u0_u0_u5_n18, u0_u0_u5_n19, u0_u0_u5_n2, u0_u0_u5_n20, u0_u0_u5_n21, u0_u0_u5_n22, u0_u0_u5_n23, 
       u0_u0_u5_n24, u0_u0_u5_n25, u0_u0_u5_n26, u0_u0_u5_n27, u0_u0_u5_n28, u0_u0_u5_n29, u0_u0_u5_n3, u0_u0_u5_n30, u0_u0_u5_n31, 
       u0_u0_u5_n32, u0_u0_u5_n33, u0_u0_u5_n34, u0_u0_u5_n35, u0_u0_u5_n36, u0_u0_u5_n37, u0_u0_u5_n38, u0_u0_u5_n39, u0_u0_u5_n4, 
       u0_u0_u5_n40, u0_u0_u5_n41, u0_u0_u5_n42, u0_u0_u5_n43, u0_u0_u5_n44, u0_u0_u5_n45, u0_u0_u5_n46, u0_u0_u5_n47, u0_u0_u5_n48, 
       u0_u0_u5_n49, u0_u0_u5_n5, u0_u0_u5_n50, u0_u0_u5_n51, u0_u0_u5_n52, u0_u0_u5_n53, u0_u0_u5_n54, u0_u0_u5_n55, u0_u0_u5_n56, 
       u0_u0_u5_n57, u0_u0_u5_n58, u0_u0_u5_n59, u0_u0_u5_n6, u0_u0_u5_n60, u0_u0_u5_n61, u0_u0_u5_n62, u0_u0_u5_n63, u0_u0_u5_n64, 
       u0_u0_u5_n65, u0_u0_u5_n66, u0_u0_u5_n67, u0_u0_u5_n68, u0_u0_u5_n69, u0_u0_u5_n7, u0_u0_u5_n70, u0_u0_u5_n71, u0_u0_u5_n72, 
       u0_u0_u5_n73, u0_u0_u5_n74, u0_u0_u5_n75, u0_u0_u5_n76, u0_u0_u5_n77, u0_u0_u5_n78, u0_u0_u5_n79, u0_u0_u5_n8, u0_u0_u5_n80, 
       u0_u0_u5_n81, u0_u0_u5_n82, u0_u0_u5_n83, u0_u0_u5_n84, u0_u0_u5_n85, u0_u0_u5_n86, u0_u0_u5_n87, u0_u0_u5_n88, u0_u0_u5_n89, 
       u0_u0_u5_n9, u0_u0_u5_n90, u0_u0_u5_n91, u0_u0_u5_n92, u0_u0_u5_n93, u0_u0_u5_n94, u0_u0_u5_n95, u0_u0_u5_n96, u0_u0_u5_n97, 
       u0_u0_u5_n98, u0_u0_u6_n1, u0_u0_u6_n10, u0_u0_u6_n11, u0_u0_u6_n12, u0_u0_u6_n13, u0_u0_u6_n14, u0_u0_u6_n15, u0_u0_u6_n16, 
       u0_u0_u6_n17, u0_u0_u6_n18, u0_u0_u6_n19, u0_u0_u6_n2, u0_u0_u6_n20, u0_u0_u6_n21, u0_u0_u6_n22, u0_u0_u6_n23, u0_u0_u6_n24, 
       u0_u0_u6_n25, u0_u0_u6_n26, u0_u0_u6_n27, u0_u0_u6_n28, u0_u0_u6_n29, u0_u0_u6_n3, u0_u0_u6_n30, u0_u0_u6_n31, u0_u0_u6_n32, 
       u0_u0_u6_n33, u0_u0_u6_n34, u0_u0_u6_n35, u0_u0_u6_n36, u0_u0_u6_n37, u0_u0_u6_n38, u0_u0_u6_n39, u0_u0_u6_n4, u0_u0_u6_n40, 
       u0_u0_u6_n41, u0_u0_u6_n42, u0_u0_u6_n43, u0_u0_u6_n44, u0_u0_u6_n45, u0_u0_u6_n46, u0_u0_u6_n47, u0_u0_u6_n48, u0_u0_u6_n49, 
       u0_u0_u6_n5, u0_u0_u6_n50, u0_u0_u6_n51, u0_u0_u6_n52, u0_u0_u6_n53, u0_u0_u6_n54, u0_u0_u6_n55, u0_u0_u6_n56, u0_u0_u6_n57, 
       u0_u0_u6_n58, u0_u0_u6_n59, u0_u0_u6_n6, u0_u0_u6_n60, u0_u0_u6_n61, u0_u0_u6_n62, u0_u0_u6_n63, u0_u0_u6_n64, u0_u0_u6_n65, 
       u0_u0_u6_n66, u0_u0_u6_n67, u0_u0_u6_n68, u0_u0_u6_n69, u0_u0_u6_n7, u0_u0_u6_n70, u0_u0_u6_n71, u0_u0_u6_n72, u0_u0_u6_n73, 
       u0_u0_u6_n74, u0_u0_u6_n75, u0_u0_u6_n76, u0_u0_u6_n77, u0_u0_u6_n78, u0_u0_u6_n79, u0_u0_u6_n8, u0_u0_u6_n80, u0_u0_u6_n81, 
       u0_u0_u6_n82, u0_u0_u6_n83, u0_u0_u6_n84, u0_u0_u6_n85, u0_u0_u6_n86, u0_u0_u6_n87, u0_u0_u6_n9, u0_u0_u7_n1, u0_u0_u7_n10, 
       u0_u0_u7_n11, u0_u0_u7_n12, u0_u0_u7_n13, u0_u0_u7_n14, u0_u0_u7_n15, u0_u0_u7_n16, u0_u0_u7_n17, u0_u0_u7_n18, u0_u0_u7_n19, 
       u0_u0_u7_n2, u0_u0_u7_n20, u0_u0_u7_n21, u0_u0_u7_n22, u0_u0_u7_n23, u0_u0_u7_n24, u0_u0_u7_n25, u0_u0_u7_n26, u0_u0_u7_n27, 
       u0_u0_u7_n28, u0_u0_u7_n29, u0_u0_u7_n3, u0_u0_u7_n30, u0_u0_u7_n31, u0_u0_u7_n32, u0_u0_u7_n33, u0_u0_u7_n34, u0_u0_u7_n35, 
       u0_u0_u7_n36, u0_u0_u7_n37, u0_u0_u7_n38, u0_u0_u7_n39, u0_u0_u7_n4, u0_u0_u7_n40, u0_u0_u7_n41, u0_u0_u7_n42, u0_u0_u7_n43, 
       u0_u0_u7_n44, u0_u0_u7_n45, u0_u0_u7_n46, u0_u0_u7_n47, u0_u0_u7_n48, u0_u0_u7_n49, u0_u0_u7_n5, u0_u0_u7_n50, u0_u0_u7_n51, 
       u0_u0_u7_n52, u0_u0_u7_n53, u0_u0_u7_n54, u0_u0_u7_n55, u0_u0_u7_n56, u0_u0_u7_n57, u0_u0_u7_n58, u0_u0_u7_n59, u0_u0_u7_n6, 
       u0_u0_u7_n60, u0_u0_u7_n61, u0_u0_u7_n62, u0_u0_u7_n63, u0_u0_u7_n64, u0_u0_u7_n65, u0_u0_u7_n66, u0_u0_u7_n67, u0_u0_u7_n68, 
       u0_u0_u7_n69, u0_u0_u7_n7, u0_u0_u7_n70, u0_u0_u7_n71, u0_u0_u7_n72, u0_u0_u7_n73, u0_u0_u7_n74, u0_u0_u7_n75, u0_u0_u7_n76, 
       u0_u0_u7_n77, u0_u0_u7_n78, u0_u0_u7_n79, u0_u0_u7_n8, u0_u0_u7_n80, u0_u0_u7_n81, u0_u0_u7_n82, u0_u0_u7_n83, u0_u0_u7_n84, 
       u0_u0_u7_n85, u0_u0_u7_n86, u0_u0_u7_n87, u0_u0_u7_n88, u0_u0_u7_n89, u0_u0_u7_n9, u0_u0_u7_n90, u0_u13_X_37, u0_u13_X_38, 
       u0_u13_X_39, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_45, u0_u13_X_46, u0_u13_X_47, 
       u0_u13_X_48, u0_u13_u6_n100, u0_u13_u6_n101, u0_u13_u6_n102, u0_u13_u6_n103, u0_u13_u6_n104, u0_u13_u6_n105, u0_u13_u6_n106, u0_u13_u6_n107, 
       u0_u13_u6_n108, u0_u13_u6_n109, u0_u13_u6_n110, u0_u13_u6_n111, u0_u13_u6_n112, u0_u13_u6_n113, u0_u13_u6_n114, u0_u13_u6_n115, u0_u13_u6_n116, 
       u0_u13_u6_n117, u0_u13_u6_n118, u0_u13_u6_n119, u0_u13_u6_n120, u0_u13_u6_n121, u0_u13_u6_n122, u0_u13_u6_n123, u0_u13_u6_n124, u0_u13_u6_n125, 
       u0_u13_u6_n126, u0_u13_u6_n127, u0_u13_u6_n128, u0_u13_u6_n129, u0_u13_u6_n130, u0_u13_u6_n131, u0_u13_u6_n132, u0_u13_u6_n133, u0_u13_u6_n134, 
       u0_u13_u6_n135, u0_u13_u6_n136, u0_u13_u6_n137, u0_u13_u6_n138, u0_u13_u6_n139, u0_u13_u6_n140, u0_u13_u6_n141, u0_u13_u6_n142, u0_u13_u6_n143, 
       u0_u13_u6_n144, u0_u13_u6_n145, u0_u13_u6_n146, u0_u13_u6_n147, u0_u13_u6_n148, u0_u13_u6_n149, u0_u13_u6_n150, u0_u13_u6_n151, u0_u13_u6_n152, 
       u0_u13_u6_n153, u0_u13_u6_n154, u0_u13_u6_n155, u0_u13_u6_n156, u0_u13_u6_n157, u0_u13_u6_n158, u0_u13_u6_n159, u0_u13_u6_n160, u0_u13_u6_n161, 
       u0_u13_u6_n162, u0_u13_u6_n163, u0_u13_u6_n164, u0_u13_u6_n165, u0_u13_u6_n166, u0_u13_u6_n167, u0_u13_u6_n168, u0_u13_u6_n169, u0_u13_u6_n170, 
       u0_u13_u6_n171, u0_u13_u6_n172, u0_u13_u6_n173, u0_u13_u6_n174, u0_u13_u6_n88, u0_u13_u6_n89, u0_u13_u6_n90, u0_u13_u6_n91, u0_u13_u6_n92, 
       u0_u13_u6_n93, u0_u13_u6_n94, u0_u13_u6_n95, u0_u13_u6_n96, u0_u13_u6_n97, u0_u13_u6_n98, u0_u13_u6_n99, u0_u13_u7_n100, u0_u13_u7_n101, 
       u0_u13_u7_n102, u0_u13_u7_n103, u0_u13_u7_n104, u0_u13_u7_n105, u0_u13_u7_n106, u0_u13_u7_n107, u0_u13_u7_n108, u0_u13_u7_n109, u0_u13_u7_n110, 
       u0_u13_u7_n111, u0_u13_u7_n112, u0_u13_u7_n113, u0_u13_u7_n114, u0_u13_u7_n115, u0_u13_u7_n116, u0_u13_u7_n117, u0_u13_u7_n118, u0_u13_u7_n119, 
       u0_u13_u7_n120, u0_u13_u7_n121, u0_u13_u7_n122, u0_u13_u7_n123, u0_u13_u7_n124, u0_u13_u7_n125, u0_u13_u7_n126, u0_u13_u7_n127, u0_u13_u7_n128, 
       u0_u13_u7_n129, u0_u13_u7_n130, u0_u13_u7_n131, u0_u13_u7_n132, u0_u13_u7_n133, u0_u13_u7_n134, u0_u13_u7_n135, u0_u13_u7_n136, u0_u13_u7_n137, 
       u0_u13_u7_n138, u0_u13_u7_n139, u0_u13_u7_n140, u0_u13_u7_n141, u0_u13_u7_n142, u0_u13_u7_n143, u0_u13_u7_n144, u0_u13_u7_n145, u0_u13_u7_n146, 
       u0_u13_u7_n147, u0_u13_u7_n148, u0_u13_u7_n149, u0_u13_u7_n150, u0_u13_u7_n151, u0_u13_u7_n152, u0_u13_u7_n153, u0_u13_u7_n154, u0_u13_u7_n155, 
       u0_u13_u7_n156, u0_u13_u7_n157, u0_u13_u7_n158, u0_u13_u7_n159, u0_u13_u7_n160, u0_u13_u7_n161, u0_u13_u7_n162, u0_u13_u7_n163, u0_u13_u7_n164, 
       u0_u13_u7_n165, u0_u13_u7_n166, u0_u13_u7_n167, u0_u13_u7_n168, u0_u13_u7_n169, u0_u13_u7_n170, u0_u13_u7_n171, u0_u13_u7_n172, u0_u13_u7_n173, 
       u0_u13_u7_n174, u0_u13_u7_n175, u0_u13_u7_n176, u0_u13_u7_n177, u0_u13_u7_n178, u0_u13_u7_n179, u0_u13_u7_n180, u0_u13_u7_n91, u0_u13_u7_n92, 
       u0_u13_u7_n93, u0_u13_u7_n94, u0_u13_u7_n95, u0_u13_u7_n96, u0_u13_u7_n97, u0_u13_u7_n98, u0_u13_u7_n99, u0_u4_X_1, u0_u4_X_2, 
       u0_u4_X_3, u0_u4_X_31, u0_u4_X_32, u0_u4_X_33, u0_u4_X_34, u0_u4_X_35, u0_u4_X_36, u0_u4_X_37, u0_u4_X_38, 
       u0_u4_X_39, u0_u4_X_4, u0_u4_X_40, u0_u4_X_41, u0_u4_X_42, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, 
       u0_u4_X_47, u0_u4_X_48, u0_u4_X_5, u0_u4_X_6, u0_u4_u0_n100, u0_u4_u0_n101, u0_u4_u0_n102, u0_u4_u0_n103, u0_u4_u0_n104, 
       u0_u4_u0_n105, u0_u4_u0_n106, u0_u4_u0_n107, u0_u4_u0_n108, u0_u4_u0_n109, u0_u4_u0_n110, u0_u4_u0_n111, u0_u4_u0_n112, u0_u4_u0_n113, 
       u0_u4_u0_n114, u0_u4_u0_n115, u0_u4_u0_n116, u0_u4_u0_n117, u0_u4_u0_n118, u0_u4_u0_n119, u0_u4_u0_n120, u0_u4_u0_n121, u0_u4_u0_n122, 
       u0_u4_u0_n123, u0_u4_u0_n124, u0_u4_u0_n125, u0_u4_u0_n126, u0_u4_u0_n127, u0_u4_u0_n128, u0_u4_u0_n129, u0_u4_u0_n130, u0_u4_u0_n131, 
       u0_u4_u0_n132, u0_u4_u0_n133, u0_u4_u0_n134, u0_u4_u0_n135, u0_u4_u0_n136, u0_u4_u0_n137, u0_u4_u0_n138, u0_u4_u0_n139, u0_u4_u0_n140, 
       u0_u4_u0_n141, u0_u4_u0_n142, u0_u4_u0_n143, u0_u4_u0_n144, u0_u4_u0_n145, u0_u4_u0_n146, u0_u4_u0_n147, u0_u4_u0_n148, u0_u4_u0_n149, 
       u0_u4_u0_n150, u0_u4_u0_n151, u0_u4_u0_n152, u0_u4_u0_n153, u0_u4_u0_n154, u0_u4_u0_n155, u0_u4_u0_n156, u0_u4_u0_n157, u0_u4_u0_n158, 
       u0_u4_u0_n159, u0_u4_u0_n160, u0_u4_u0_n161, u0_u4_u0_n162, u0_u4_u0_n163, u0_u4_u0_n164, u0_u4_u0_n165, u0_u4_u0_n166, u0_u4_u0_n167, 
       u0_u4_u0_n168, u0_u4_u0_n169, u0_u4_u0_n170, u0_u4_u0_n171, u0_u4_u0_n172, u0_u4_u0_n173, u0_u4_u0_n174, u0_u4_u0_n88, u0_u4_u0_n89, 
       u0_u4_u0_n90, u0_u4_u0_n91, u0_u4_u0_n92, u0_u4_u0_n93, u0_u4_u0_n94, u0_u4_u0_n95, u0_u4_u0_n96, u0_u4_u0_n97, u0_u4_u0_n98, 
       u0_u4_u0_n99, u0_u4_u5_n100, u0_u4_u5_n101, u0_u4_u5_n102, u0_u4_u5_n103, u0_u4_u5_n104, u0_u4_u5_n105, u0_u4_u5_n106, u0_u4_u5_n107, 
       u0_u4_u5_n108, u0_u4_u5_n109, u0_u4_u5_n110, u0_u4_u5_n111, u0_u4_u5_n112, u0_u4_u5_n113, u0_u4_u5_n114, u0_u4_u5_n115, u0_u4_u5_n116, 
       u0_u4_u5_n117, u0_u4_u5_n118, u0_u4_u5_n119, u0_u4_u5_n120, u0_u4_u5_n121, u0_u4_u5_n122, u0_u4_u5_n123, u0_u4_u5_n124, u0_u4_u5_n125, 
       u0_u4_u5_n126, u0_u4_u5_n127, u0_u4_u5_n128, u0_u4_u5_n129, u0_u4_u5_n130, u0_u4_u5_n131, u0_u4_u5_n132, u0_u4_u5_n133, u0_u4_u5_n134, 
       u0_u4_u5_n135, u0_u4_u5_n136, u0_u4_u5_n137, u0_u4_u5_n138, u0_u4_u5_n139, u0_u4_u5_n140, u0_u4_u5_n141, u0_u4_u5_n142, u0_u4_u5_n143, 
       u0_u4_u5_n144, u0_u4_u5_n145, u0_u4_u5_n146, u0_u4_u5_n147, u0_u4_u5_n148, u0_u4_u5_n149, u0_u4_u5_n150, u0_u4_u5_n151, u0_u4_u5_n152, 
       u0_u4_u5_n153, u0_u4_u5_n154, u0_u4_u5_n155, u0_u4_u5_n156, u0_u4_u5_n157, u0_u4_u5_n158, u0_u4_u5_n159, u0_u4_u5_n160, u0_u4_u5_n161, 
       u0_u4_u5_n162, u0_u4_u5_n163, u0_u4_u5_n164, u0_u4_u5_n165, u0_u4_u5_n166, u0_u4_u5_n167, u0_u4_u5_n168, u0_u4_u5_n169, u0_u4_u5_n170, 
       u0_u4_u5_n171, u0_u4_u5_n172, u0_u4_u5_n173, u0_u4_u5_n174, u0_u4_u5_n175, u0_u4_u5_n176, u0_u4_u5_n177, u0_u4_u5_n178, u0_u4_u5_n179, 
       u0_u4_u5_n180, u0_u4_u5_n181, u0_u4_u5_n182, u0_u4_u5_n183, u0_u4_u5_n184, u0_u4_u5_n185, u0_u4_u5_n186, u0_u4_u5_n187, u0_u4_u5_n188, 
       u0_u4_u5_n189, u0_u4_u5_n190, u0_u4_u5_n191, u0_u4_u5_n192, u0_u4_u5_n193, u0_u4_u5_n194, u0_u4_u5_n195, u0_u4_u5_n196, u0_u4_u5_n99, 
       u0_u4_u6_n100, u0_u4_u6_n101, u0_u4_u6_n102, u0_u4_u6_n103, u0_u4_u6_n104, u0_u4_u6_n105, u0_u4_u6_n106, u0_u4_u6_n107, u0_u4_u6_n108, 
       u0_u4_u6_n109, u0_u4_u6_n110, u0_u4_u6_n111, u0_u4_u6_n112, u0_u4_u6_n113, u0_u4_u6_n114, u0_u4_u6_n115, u0_u4_u6_n116, u0_u4_u6_n117, 
       u0_u4_u6_n118, u0_u4_u6_n119, u0_u4_u6_n120, u0_u4_u6_n121, u0_u4_u6_n122, u0_u4_u6_n123, u0_u4_u6_n124, u0_u4_u6_n125, u0_u4_u6_n126, 
       u0_u4_u6_n127, u0_u4_u6_n128, u0_u4_u6_n129, u0_u4_u6_n130, u0_u4_u6_n131, u0_u4_u6_n132, u0_u4_u6_n133, u0_u4_u6_n134, u0_u4_u6_n135, 
       u0_u4_u6_n136, u0_u4_u6_n137, u0_u4_u6_n138, u0_u4_u6_n139, u0_u4_u6_n140, u0_u4_u6_n141, u0_u4_u6_n142, u0_u4_u6_n143, u0_u4_u6_n144, 
       u0_u4_u6_n145, u0_u4_u6_n146, u0_u4_u6_n147, u0_u4_u6_n148, u0_u4_u6_n149, u0_u4_u6_n150, u0_u4_u6_n151, u0_u4_u6_n152, u0_u4_u6_n153, 
       u0_u4_u6_n154, u0_u4_u6_n155, u0_u4_u6_n156, u0_u4_u6_n157, u0_u4_u6_n158, u0_u4_u6_n159, u0_u4_u6_n160, u0_u4_u6_n161, u0_u4_u6_n162, 
       u0_u4_u6_n163, u0_u4_u6_n164, u0_u4_u6_n165, u0_u4_u6_n166, u0_u4_u6_n167, u0_u4_u6_n168, u0_u4_u6_n169, u0_u4_u6_n170, u0_u4_u6_n171, 
       u0_u4_u6_n172, u0_u4_u6_n173, u0_u4_u6_n174, u0_u4_u6_n88, u0_u4_u6_n89, u0_u4_u6_n90, u0_u4_u6_n91, u0_u4_u6_n92, u0_u4_u6_n93, 
       u0_u4_u6_n94, u0_u4_u6_n95, u0_u4_u6_n96, u0_u4_u6_n97, u0_u4_u6_n98, u0_u4_u6_n99, u0_u4_u7_n100, u0_u4_u7_n101, u0_u4_u7_n102, 
       u0_u4_u7_n103, u0_u4_u7_n104, u0_u4_u7_n105, u0_u4_u7_n106, u0_u4_u7_n107, u0_u4_u7_n108, u0_u4_u7_n109, u0_u4_u7_n110, u0_u4_u7_n111, 
       u0_u4_u7_n112, u0_u4_u7_n113, u0_u4_u7_n114, u0_u4_u7_n115, u0_u4_u7_n116, u0_u4_u7_n117, u0_u4_u7_n118, u0_u4_u7_n119, u0_u4_u7_n120, 
       u0_u4_u7_n121, u0_u4_u7_n122, u0_u4_u7_n123, u0_u4_u7_n124, u0_u4_u7_n125, u0_u4_u7_n126, u0_u4_u7_n127, u0_u4_u7_n128, u0_u4_u7_n129, 
       u0_u4_u7_n130, u0_u4_u7_n131, u0_u4_u7_n132, u0_u4_u7_n133, u0_u4_u7_n134, u0_u4_u7_n135, u0_u4_u7_n136, u0_u4_u7_n137, u0_u4_u7_n138, 
       u0_u4_u7_n139, u0_u4_u7_n140, u0_u4_u7_n141, u0_u4_u7_n142, u0_u4_u7_n143, u0_u4_u7_n144, u0_u4_u7_n145, u0_u4_u7_n146, u0_u4_u7_n147, 
       u0_u4_u7_n148, u0_u4_u7_n149, u0_u4_u7_n150, u0_u4_u7_n151, u0_u4_u7_n152, u0_u4_u7_n153, u0_u4_u7_n154, u0_u4_u7_n155, u0_u4_u7_n156, 
       u0_u4_u7_n157, u0_u4_u7_n158, u0_u4_u7_n159, u0_u4_u7_n160, u0_u4_u7_n161, u0_u4_u7_n162, u0_u4_u7_n163, u0_u4_u7_n164, u0_u4_u7_n165, 
       u0_u4_u7_n166, u0_u4_u7_n167, u0_u4_u7_n168, u0_u4_u7_n169, u0_u4_u7_n170, u0_u4_u7_n171, u0_u4_u7_n172, u0_u4_u7_n173, u0_u4_u7_n174, 
       u0_u4_u7_n175, u0_u4_u7_n176, u0_u4_u7_n177, u0_u4_u7_n178, u0_u4_u7_n179, u0_u4_u7_n180, u0_u4_u7_n91, u0_u4_u7_n92, u0_u4_u7_n93, 
       u0_u4_u7_n94, u0_u4_u7_n95, u0_u4_u7_n96, u0_u4_u7_n97, u0_u4_u7_n98, u0_u4_u7_n99, u0_uk_n693, u0_uk_n700, u0_uk_n701, 
       u0_uk_n706, u0_uk_n709, u0_uk_n710, u0_uk_n714, u0_uk_n716, u0_uk_n803, u0_uk_n806, u0_uk_n807, u0_uk_n808, 
       u0_uk_n809, u0_uk_n811, u0_uk_n870, u0_uk_n872, u0_uk_n873, u0_uk_n874, u0_uk_n876, u0_uk_n877, u0_uk_n879, 
       u0_uk_n882, u0_uk_n883, u0_uk_n884, u0_uk_n929, u0_uk_n930, u0_uk_n931, u2_K10_19, u2_K10_20, u2_K10_21, 
       u2_K10_22, u2_K10_23, u2_K10_24, u2_K10_27, u2_K10_28, u2_K10_29, u2_K10_31, u2_K10_33, u2_K10_35, 
       u2_K10_37, u2_K10_38, u2_K10_39, u2_K10_40, u2_K10_41, u2_K11_14, u2_K11_15, u2_K11_17, u2_K11_31, 
       u2_K11_32, u2_K11_33, u2_K11_34, u2_K11_35, u2_K11_36, u2_K11_37, u2_K11_39, u2_K11_40, u2_K11_41, 
       u2_K11_43, u2_K11_44, u2_K11_46, u2_K11_47, u2_K12_19, u2_K12_21, u2_K12_23, u2_K12_28, u2_K12_30, 
       u2_K12_31, u2_K12_32, u2_K12_33, u2_K12_35, u2_K12_36, u2_K12_38, u2_K12_39, u2_K12_40, u2_K12_42, 
       u2_K12_43, u2_K12_44, u2_K12_45, u2_K12_48, u2_K13_1, u2_K13_10, u2_K13_11, u2_K13_12, u2_K13_13, 
       u2_K13_15, u2_K13_16, u2_K13_17, u2_K13_18, u2_K13_19, u2_K13_2, u2_K13_21, u2_K13_22, u2_K13_23, 
       u2_K13_24, u2_K13_25, u2_K13_27, u2_K13_28, u2_K13_29, u2_K13_30, u2_K13_33, u2_K13_35, u2_K13_36, 
       u2_K13_4, u2_K13_5, u2_K13_6, u2_K13_7, u2_K13_9, u2_K15_14, u2_K15_15, u2_K15_17, u2_K15_19, 
       u2_K15_22, u2_K15_24, u2_K15_43, u2_K15_44, u2_K15_45, u2_K15_46, u2_K15_47, u2_K15_48, u2_K16_10, 
       u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_15, u2_K16_16, u2_K16_17, u2_K16_18, u2_K16_19, 
       u2_K16_20, u2_K16_21, u2_K16_22, u2_K16_23, u2_K16_24, u2_K16_7, u2_K1_25, u2_K1_26, u2_K1_27, 
       u2_K1_29, u2_K1_30, u2_K1_31, u2_K1_32, u2_K1_33, u2_K1_34, u2_K1_35, u2_K1_36, u2_K1_38, 
       u2_K1_39, u2_K1_41, u2_K1_42, u2_K1_44, u2_K1_47, u2_K1_48, u2_K2_10, u2_K2_11, u2_K2_12, 
       u2_K2_13, u2_K2_14, u2_K2_15, u2_K2_17, u2_K2_19, u2_K2_21, u2_K2_22, u2_K2_23, u2_K2_24, 
       u2_K2_7, u2_K2_8, u2_K2_9, u2_K3_25, u2_K3_26, u2_K3_27, u2_K3_28, u2_K3_29, u2_K4_1, 
       u2_K4_10, u2_K4_11, u2_K4_12, u2_K4_2, u2_K4_3, u2_K4_37, u2_K4_4, u2_K4_40, u2_K4_41, 
       u2_K4_43, u2_K4_44, u2_K4_45, u2_K4_46, u2_K4_47, u2_K4_48, u2_K4_5, u2_K4_8, u2_K4_9, 
       u2_K5_27, u2_K5_29, u2_K5_30, u2_K5_33, u2_K5_35, u2_K5_36, u2_K5_37, u2_K5_39, u2_K5_40, 
       u2_K5_42, u2_K6_10, u2_K6_12, u2_K6_2, u2_K6_31, u2_K6_33, u2_K6_35, u2_K6_37, u2_K6_38, 
       u2_K6_39, u2_K6_4, u2_K6_41, u2_K6_42, u2_K6_43, u2_K6_44, u2_K6_45, u2_K6_46, u2_K6_47, 
       u2_K6_48, u2_K6_5, u2_K6_6, u2_K6_7, u2_K6_8, u2_K6_9, u2_K7_32, u2_K7_34, u2_K7_36, 
       u2_K8_25, u2_K8_27, u2_K8_28, u2_K8_29, u2_K8_30, u2_K8_32, u2_K8_33, u2_K8_34, u2_K8_35, 
       u2_K8_36, u2_K9_1, u2_K9_10, u2_K9_11, u2_K9_12, u2_K9_13, u2_K9_14, u2_K9_16, u2_K9_17, 
       u2_K9_18, u2_K9_19, u2_K9_2, u2_K9_20, u2_K9_21, u2_K9_22, u2_K9_24, u2_K9_26, u2_K9_27, 
       u2_K9_30, u2_K9_37, u2_K9_39, u2_K9_4, u2_K9_41, u2_K9_42, u2_K9_43, u2_K9_44, u2_K9_46, 
       u2_K9_47, u2_K9_48, u2_K9_6, u2_K9_7, u2_K9_8, u2_K9_9, u2_out0_11, u2_out0_12, u2_out0_14, 
       u2_out0_15, u2_out0_19, u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, u2_out0_29, u2_out0_3, u2_out0_32, 
       u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, u2_out10_11, u2_out10_12, u2_out10_15, u2_out10_16, u2_out10_19, 
       u2_out10_21, u2_out10_22, u2_out10_24, u2_out10_27, u2_out10_29, u2_out10_30, u2_out10_32, u2_out10_4, u2_out10_5, 
       u2_out10_6, u2_out10_7, u2_out11_1, u2_out11_10, u2_out11_11, u2_out11_12, u2_out11_14, u2_out11_15, u2_out11_19, 
       u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_25, u2_out11_26, u2_out11_27, u2_out11_29, u2_out11_3, u2_out11_32, 
       u2_out11_4, u2_out11_5, u2_out11_7, u2_out11_8, u2_out12_1, u2_out12_10, u2_out12_11, u2_out12_13, u2_out12_14, 
       u2_out12_16, u2_out12_17, u2_out12_18, u2_out12_19, u2_out12_2, u2_out12_20, u2_out12_23, u2_out12_24, u2_out12_25, 
       u2_out12_26, u2_out12_28, u2_out12_29, u2_out12_3, u2_out12_30, u2_out12_31, u2_out12_4, u2_out12_6, u2_out12_8, 
       u2_out12_9, u2_out14_1, u2_out14_10, u2_out14_15, u2_out14_16, u2_out14_20, u2_out14_21, u2_out14_24, u2_out14_26, 
       u2_out14_27, u2_out14_30, u2_out14_5, u2_out14_6, u2_out15_1, u2_out15_10, u2_out15_13, u2_out15_16, u2_out15_18, 
       u2_out15_2, u2_out15_20, u2_out15_24, u2_out15_26, u2_out15_28, u2_out15_30, u2_out15_6, u2_out1_1, u2_out1_10, 
       u2_out1_13, u2_out1_16, u2_out1_18, u2_out1_2, u2_out1_20, u2_out1_24, u2_out1_26, u2_out1_28, u2_out1_30, 
       u2_out1_6, u2_out2_14, u2_out2_25, u2_out2_3, u2_out2_8, u2_out3_12, u2_out3_13, u2_out3_15, u2_out3_17, 
       u2_out3_18, u2_out3_2, u2_out3_21, u2_out3_22, u2_out3_23, u2_out3_27, u2_out3_28, u2_out3_31, u2_out3_32, 
       u2_out3_5, u2_out3_7, u2_out3_9, u2_out4_11, u2_out4_12, u2_out4_14, u2_out4_19, u2_out4_22, u2_out4_25, 
       u2_out4_29, u2_out4_3, u2_out4_32, u2_out4_4, u2_out4_7, u2_out4_8, u2_out5_11, u2_out5_12, u2_out5_13, 
       u2_out5_15, u2_out5_17, u2_out5_18, u2_out5_19, u2_out5_2, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_27, 
       u2_out5_28, u2_out5_29, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, u2_out5_7, u2_out5_9, u2_out6_11, 
       u2_out6_19, u2_out6_29, u2_out6_4, u2_out7_11, u2_out7_14, u2_out7_19, u2_out7_25, u2_out7_29, u2_out7_3, 
       u2_out7_4, u2_out7_8, u2_out8_1, u2_out8_10, u2_out8_12, u2_out8_13, u2_out8_14, u2_out8_15, u2_out8_16, 
       u2_out8_17, u2_out8_18, u2_out8_2, u2_out8_20, u2_out8_21, u2_out8_22, u2_out8_23, u2_out8_24, u2_out8_25, 
       u2_out8_26, u2_out8_27, u2_out8_28, u2_out8_3, u2_out8_30, u2_out8_31, u2_out8_32, u2_out8_5, u2_out8_6, 
       u2_out8_7, u2_out8_8, u2_out8_9, u2_out9_1, u2_out9_10, u2_out9_11, u2_out9_12, u2_out9_14, u2_out9_19, 
       u2_out9_20, u2_out9_22, u2_out9_25, u2_out9_26, u2_out9_29, u2_out9_3, u2_out9_32, u2_out9_4, u2_out9_7, 
       u2_out9_8, u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_29, u2_u0_X_30, u2_u0_X_31, u2_u0_X_32, 
       u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, u2_u0_X_36, u2_u0_X_37, u2_u0_X_38, u2_u0_X_39, u2_u0_X_40, u2_u0_X_41, 
       u2_u0_X_42, u2_u0_X_43, u2_u0_X_44, u2_u0_X_45, u2_u0_X_46, u2_u0_X_47, u2_u0_X_48, u2_u0_u4_n100, u2_u0_u4_n101, 
       u2_u0_u4_n102, u2_u0_u4_n103, u2_u0_u4_n104, u2_u0_u4_n105, u2_u0_u4_n106, u2_u0_u4_n107, u2_u0_u4_n108, u2_u0_u4_n109, u2_u0_u4_n110, 
       u2_u0_u4_n111, u2_u0_u4_n112, u2_u0_u4_n113, u2_u0_u4_n114, u2_u0_u4_n115, u2_u0_u4_n116, u2_u0_u4_n117, u2_u0_u4_n118, u2_u0_u4_n119, 
       u2_u0_u4_n120, u2_u0_u4_n121, u2_u0_u4_n122, u2_u0_u4_n123, u2_u0_u4_n124, u2_u0_u4_n125, u2_u0_u4_n126, u2_u0_u4_n127, u2_u0_u4_n128, 
       u2_u0_u4_n129, u2_u0_u4_n130, u2_u0_u4_n131, u2_u0_u4_n132, u2_u0_u4_n133, u2_u0_u4_n134, u2_u0_u4_n135, u2_u0_u4_n136, u2_u0_u4_n137, 
       u2_u0_u4_n138, u2_u0_u4_n139, u2_u0_u4_n140, u2_u0_u4_n141, u2_u0_u4_n142, u2_u0_u4_n143, u2_u0_u4_n144, u2_u0_u4_n145, u2_u0_u4_n146, 
       u2_u0_u4_n147, u2_u0_u4_n148, u2_u0_u4_n149, u2_u0_u4_n150, u2_u0_u4_n151, u2_u0_u4_n152, u2_u0_u4_n153, u2_u0_u4_n154, u2_u0_u4_n155, 
       u2_u0_u4_n156, u2_u0_u4_n157, u2_u0_u4_n158, u2_u0_u4_n159, u2_u0_u4_n160, u2_u0_u4_n161, u2_u0_u4_n162, u2_u0_u4_n163, u2_u0_u4_n164, 
       u2_u0_u4_n165, u2_u0_u4_n166, u2_u0_u4_n167, u2_u0_u4_n168, u2_u0_u4_n169, u2_u0_u4_n170, u2_u0_u4_n171, u2_u0_u4_n172, u2_u0_u4_n173, 
       u2_u0_u4_n174, u2_u0_u4_n175, u2_u0_u4_n176, u2_u0_u4_n177, u2_u0_u4_n178, u2_u0_u4_n179, u2_u0_u4_n180, u2_u0_u4_n181, u2_u0_u4_n182, 
       u2_u0_u4_n183, u2_u0_u4_n184, u2_u0_u4_n185, u2_u0_u4_n186, u2_u0_u4_n94, u2_u0_u4_n95, u2_u0_u4_n96, u2_u0_u4_n97, u2_u0_u4_n98, 
       u2_u0_u4_n99, u2_u0_u5_n100, u2_u0_u5_n101, u2_u0_u5_n102, u2_u0_u5_n103, u2_u0_u5_n104, u2_u0_u5_n105, u2_u0_u5_n106, u2_u0_u5_n107, 
       u2_u0_u5_n108, u2_u0_u5_n109, u2_u0_u5_n110, u2_u0_u5_n111, u2_u0_u5_n112, u2_u0_u5_n113, u2_u0_u5_n114, u2_u0_u5_n115, u2_u0_u5_n116, 
       u2_u0_u5_n117, u2_u0_u5_n118, u2_u0_u5_n119, u2_u0_u5_n120, u2_u0_u5_n121, u2_u0_u5_n122, u2_u0_u5_n123, u2_u0_u5_n124, u2_u0_u5_n125, 
       u2_u0_u5_n126, u2_u0_u5_n127, u2_u0_u5_n128, u2_u0_u5_n129, u2_u0_u5_n130, u2_u0_u5_n131, u2_u0_u5_n132, u2_u0_u5_n133, u2_u0_u5_n134, 
       u2_u0_u5_n135, u2_u0_u5_n136, u2_u0_u5_n137, u2_u0_u5_n138, u2_u0_u5_n139, u2_u0_u5_n140, u2_u0_u5_n141, u2_u0_u5_n142, u2_u0_u5_n143, 
       u2_u0_u5_n144, u2_u0_u5_n145, u2_u0_u5_n146, u2_u0_u5_n147, u2_u0_u5_n148, u2_u0_u5_n149, u2_u0_u5_n150, u2_u0_u5_n151, u2_u0_u5_n152, 
       u2_u0_u5_n153, u2_u0_u5_n154, u2_u0_u5_n155, u2_u0_u5_n156, u2_u0_u5_n157, u2_u0_u5_n158, u2_u0_u5_n159, u2_u0_u5_n160, u2_u0_u5_n161, 
       u2_u0_u5_n162, u2_u0_u5_n163, u2_u0_u5_n164, u2_u0_u5_n165, u2_u0_u5_n166, u2_u0_u5_n167, u2_u0_u5_n168, u2_u0_u5_n169, u2_u0_u5_n170, 
       u2_u0_u5_n171, u2_u0_u5_n172, u2_u0_u5_n173, u2_u0_u5_n174, u2_u0_u5_n175, u2_u0_u5_n176, u2_u0_u5_n177, u2_u0_u5_n178, u2_u0_u5_n179, 
       u2_u0_u5_n180, u2_u0_u5_n181, u2_u0_u5_n182, u2_u0_u5_n183, u2_u0_u5_n184, u2_u0_u5_n185, u2_u0_u5_n186, u2_u0_u5_n187, u2_u0_u5_n188, 
       u2_u0_u5_n189, u2_u0_u5_n190, u2_u0_u5_n191, u2_u0_u5_n192, u2_u0_u5_n193, u2_u0_u5_n194, u2_u0_u5_n195, u2_u0_u5_n196, u2_u0_u5_n99, 
       u2_u0_u6_n100, u2_u0_u6_n101, u2_u0_u6_n102, u2_u0_u6_n103, u2_u0_u6_n104, u2_u0_u6_n105, u2_u0_u6_n106, u2_u0_u6_n107, u2_u0_u6_n108, 
       u2_u0_u6_n109, u2_u0_u6_n110, u2_u0_u6_n111, u2_u0_u6_n112, u2_u0_u6_n113, u2_u0_u6_n114, u2_u0_u6_n115, u2_u0_u6_n116, u2_u0_u6_n117, 
       u2_u0_u6_n118, u2_u0_u6_n119, u2_u0_u6_n120, u2_u0_u6_n121, u2_u0_u6_n122, u2_u0_u6_n123, u2_u0_u6_n124, u2_u0_u6_n125, u2_u0_u6_n126, 
       u2_u0_u6_n127, u2_u0_u6_n128, u2_u0_u6_n129, u2_u0_u6_n130, u2_u0_u6_n131, u2_u0_u6_n132, u2_u0_u6_n133, u2_u0_u6_n134, u2_u0_u6_n135, 
       u2_u0_u6_n136, u2_u0_u6_n137, u2_u0_u6_n138, u2_u0_u6_n139, u2_u0_u6_n140, u2_u0_u6_n141, u2_u0_u6_n142, u2_u0_u6_n143, u2_u0_u6_n144, 
       u2_u0_u6_n145, u2_u0_u6_n146, u2_u0_u6_n147, u2_u0_u6_n148, u2_u0_u6_n149, u2_u0_u6_n150, u2_u0_u6_n151, u2_u0_u6_n152, u2_u0_u6_n153, 
       u2_u0_u6_n154, u2_u0_u6_n155, u2_u0_u6_n156, u2_u0_u6_n157, u2_u0_u6_n158, u2_u0_u6_n159, u2_u0_u6_n160, u2_u0_u6_n161, u2_u0_u6_n162, 
       u2_u0_u6_n163, u2_u0_u6_n164, u2_u0_u6_n165, u2_u0_u6_n166, u2_u0_u6_n167, u2_u0_u6_n168, u2_u0_u6_n169, u2_u0_u6_n170, u2_u0_u6_n171, 
       u2_u0_u6_n172, u2_u0_u6_n173, u2_u0_u6_n174, u2_u0_u6_n88, u2_u0_u6_n89, u2_u0_u6_n90, u2_u0_u6_n91, u2_u0_u6_n92, u2_u0_u6_n93, 
       u2_u0_u6_n94, u2_u0_u6_n95, u2_u0_u6_n96, u2_u0_u6_n97, u2_u0_u6_n98, u2_u0_u6_n99, u2_u0_u7_n100, u2_u0_u7_n101, u2_u0_u7_n102, 
       u2_u0_u7_n103, u2_u0_u7_n104, u2_u0_u7_n105, u2_u0_u7_n106, u2_u0_u7_n107, u2_u0_u7_n108, u2_u0_u7_n109, u2_u0_u7_n110, u2_u0_u7_n111, 
       u2_u0_u7_n112, u2_u0_u7_n113, u2_u0_u7_n114, u2_u0_u7_n115, u2_u0_u7_n116, u2_u0_u7_n117, u2_u0_u7_n118, u2_u0_u7_n119, u2_u0_u7_n120, 
       u2_u0_u7_n121, u2_u0_u7_n122, u2_u0_u7_n123, u2_u0_u7_n124, u2_u0_u7_n125, u2_u0_u7_n126, u2_u0_u7_n127, u2_u0_u7_n128, u2_u0_u7_n129, 
       u2_u0_u7_n130, u2_u0_u7_n131, u2_u0_u7_n132, u2_u0_u7_n133, u2_u0_u7_n134, u2_u0_u7_n135, u2_u0_u7_n136, u2_u0_u7_n137, u2_u0_u7_n138, 
       u2_u0_u7_n139, u2_u0_u7_n140, u2_u0_u7_n141, u2_u0_u7_n142, u2_u0_u7_n143, u2_u0_u7_n144, u2_u0_u7_n145, u2_u0_u7_n146, u2_u0_u7_n147, 
       u2_u0_u7_n148, u2_u0_u7_n149, u2_u0_u7_n150, u2_u0_u7_n151, u2_u0_u7_n152, u2_u0_u7_n153, u2_u0_u7_n154, u2_u0_u7_n155, u2_u0_u7_n156, 
       u2_u0_u7_n157, u2_u0_u7_n158, u2_u0_u7_n159, u2_u0_u7_n160, u2_u0_u7_n161, u2_u0_u7_n162, u2_u0_u7_n163, u2_u0_u7_n164, u2_u0_u7_n165, 
       u2_u0_u7_n166, u2_u0_u7_n167, u2_u0_u7_n168, u2_u0_u7_n169, u2_u0_u7_n170, u2_u0_u7_n171, u2_u0_u7_n172, u2_u0_u7_n173, u2_u0_u7_n174, 
       u2_u0_u7_n175, u2_u0_u7_n176, u2_u0_u7_n177, u2_u0_u7_n178, u2_u0_u7_n179, u2_u0_u7_n180, u2_u0_u7_n91, u2_u0_u7_n92, u2_u0_u7_n93, 
       u2_u0_u7_n94, u2_u0_u7_n95, u2_u0_u7_n96, u2_u0_u7_n97, u2_u0_u7_n98, u2_u0_u7_n99, u2_u10_X_13, u2_u10_X_14, u2_u10_X_15, 
       u2_u10_X_16, u2_u10_X_17, u2_u10_X_18, u2_u10_X_31, u2_u10_X_32, u2_u10_X_33, u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, 
       u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, 
       u2_u10_X_46, u2_u10_X_47, u2_u10_X_48, u2_u10_u2_n100, u2_u10_u2_n101, u2_u10_u2_n102, u2_u10_u2_n103, u2_u10_u2_n104, u2_u10_u2_n105, 
       u2_u10_u2_n106, u2_u10_u2_n107, u2_u10_u2_n108, u2_u10_u2_n109, u2_u10_u2_n110, u2_u10_u2_n111, u2_u10_u2_n112, u2_u10_u2_n113, u2_u10_u2_n114, 
       u2_u10_u2_n115, u2_u10_u2_n116, u2_u10_u2_n117, u2_u10_u2_n118, u2_u10_u2_n119, u2_u10_u2_n120, u2_u10_u2_n121, u2_u10_u2_n122, u2_u10_u2_n123, 
       u2_u10_u2_n124, u2_u10_u2_n125, u2_u10_u2_n126, u2_u10_u2_n127, u2_u10_u2_n128, u2_u10_u2_n129, u2_u10_u2_n130, u2_u10_u2_n131, u2_u10_u2_n132, 
       u2_u10_u2_n133, u2_u10_u2_n134, u2_u10_u2_n135, u2_u10_u2_n136, u2_u10_u2_n137, u2_u10_u2_n138, u2_u10_u2_n139, u2_u10_u2_n140, u2_u10_u2_n141, 
       u2_u10_u2_n142, u2_u10_u2_n143, u2_u10_u2_n144, u2_u10_u2_n145, u2_u10_u2_n146, u2_u10_u2_n147, u2_u10_u2_n148, u2_u10_u2_n149, u2_u10_u2_n150, 
       u2_u10_u2_n151, u2_u10_u2_n152, u2_u10_u2_n153, u2_u10_u2_n154, u2_u10_u2_n155, u2_u10_u2_n156, u2_u10_u2_n157, u2_u10_u2_n158, u2_u10_u2_n159, 
       u2_u10_u2_n160, u2_u10_u2_n161, u2_u10_u2_n162, u2_u10_u2_n163, u2_u10_u2_n164, u2_u10_u2_n165, u2_u10_u2_n166, u2_u10_u2_n167, u2_u10_u2_n168, 
       u2_u10_u2_n169, u2_u10_u2_n170, u2_u10_u2_n171, u2_u10_u2_n172, u2_u10_u2_n173, u2_u10_u2_n174, u2_u10_u2_n175, u2_u10_u2_n176, u2_u10_u2_n177, 
       u2_u10_u2_n178, u2_u10_u2_n179, u2_u10_u2_n180, u2_u10_u2_n181, u2_u10_u2_n182, u2_u10_u2_n183, u2_u10_u2_n184, u2_u10_u2_n185, u2_u10_u2_n186, 
       u2_u10_u2_n187, u2_u10_u2_n188, u2_u10_u2_n95, u2_u10_u2_n96, u2_u10_u2_n97, u2_u10_u2_n98, u2_u10_u2_n99, u2_u10_u5_n100, u2_u10_u5_n101, 
       u2_u10_u5_n102, u2_u10_u5_n103, u2_u10_u5_n104, u2_u10_u5_n105, u2_u10_u5_n106, u2_u10_u5_n107, u2_u10_u5_n108, u2_u10_u5_n109, u2_u10_u5_n110, 
       u2_u10_u5_n111, u2_u10_u5_n112, u2_u10_u5_n113, u2_u10_u5_n114, u2_u10_u5_n115, u2_u10_u5_n116, u2_u10_u5_n117, u2_u10_u5_n118, u2_u10_u5_n119, 
       u2_u10_u5_n120, u2_u10_u5_n121, u2_u10_u5_n122, u2_u10_u5_n123, u2_u10_u5_n124, u2_u10_u5_n125, u2_u10_u5_n126, u2_u10_u5_n127, u2_u10_u5_n128, 
       u2_u10_u5_n129, u2_u10_u5_n130, u2_u10_u5_n131, u2_u10_u5_n132, u2_u10_u5_n133, u2_u10_u5_n134, u2_u10_u5_n135, u2_u10_u5_n136, u2_u10_u5_n137, 
       u2_u10_u5_n138, u2_u10_u5_n139, u2_u10_u5_n140, u2_u10_u5_n141, u2_u10_u5_n142, u2_u10_u5_n143, u2_u10_u5_n144, u2_u10_u5_n145, u2_u10_u5_n146, 
       u2_u10_u5_n147, u2_u10_u5_n148, u2_u10_u5_n149, u2_u10_u5_n150, u2_u10_u5_n151, u2_u10_u5_n152, u2_u10_u5_n153, u2_u10_u5_n154, u2_u10_u5_n155, 
       u2_u10_u5_n156, u2_u10_u5_n157, u2_u10_u5_n158, u2_u10_u5_n159, u2_u10_u5_n160, u2_u10_u5_n161, u2_u10_u5_n162, u2_u10_u5_n163, u2_u10_u5_n164, 
       u2_u10_u5_n165, u2_u10_u5_n166, u2_u10_u5_n167, u2_u10_u5_n168, u2_u10_u5_n169, u2_u10_u5_n170, u2_u10_u5_n171, u2_u10_u5_n172, u2_u10_u5_n173, 
       u2_u10_u5_n174, u2_u10_u5_n175, u2_u10_u5_n176, u2_u10_u5_n177, u2_u10_u5_n178, u2_u10_u5_n179, u2_u10_u5_n180, u2_u10_u5_n181, u2_u10_u5_n182, 
       u2_u10_u5_n183, u2_u10_u5_n184, u2_u10_u5_n185, u2_u10_u5_n186, u2_u10_u5_n187, u2_u10_u5_n188, u2_u10_u5_n189, u2_u10_u5_n190, u2_u10_u5_n191, 
       u2_u10_u5_n192, u2_u10_u5_n193, u2_u10_u5_n194, u2_u10_u5_n195, u2_u10_u5_n196, u2_u10_u5_n99, u2_u10_u6_n100, u2_u10_u6_n101, u2_u10_u6_n102, 
       u2_u10_u6_n103, u2_u10_u6_n104, u2_u10_u6_n105, u2_u10_u6_n106, u2_u10_u6_n107, u2_u10_u6_n108, u2_u10_u6_n109, u2_u10_u6_n110, u2_u10_u6_n111, 
       u2_u10_u6_n112, u2_u10_u6_n113, u2_u10_u6_n114, u2_u10_u6_n115, u2_u10_u6_n116, u2_u10_u6_n117, u2_u10_u6_n118, u2_u10_u6_n119, u2_u10_u6_n120, 
       u2_u10_u6_n121, u2_u10_u6_n122, u2_u10_u6_n123, u2_u10_u6_n124, u2_u10_u6_n125, u2_u10_u6_n126, u2_u10_u6_n127, u2_u10_u6_n128, u2_u10_u6_n129, 
       u2_u10_u6_n130, u2_u10_u6_n131, u2_u10_u6_n132, u2_u10_u6_n133, u2_u10_u6_n134, u2_u10_u6_n135, u2_u10_u6_n136, u2_u10_u6_n137, u2_u10_u6_n138, 
       u2_u10_u6_n139, u2_u10_u6_n140, u2_u10_u6_n141, u2_u10_u6_n142, u2_u10_u6_n143, u2_u10_u6_n144, u2_u10_u6_n145, u2_u10_u6_n146, u2_u10_u6_n147, 
       u2_u10_u6_n148, u2_u10_u6_n149, u2_u10_u6_n150, u2_u10_u6_n151, u2_u10_u6_n152, u2_u10_u6_n153, u2_u10_u6_n154, u2_u10_u6_n155, u2_u10_u6_n156, 
       u2_u10_u6_n157, u2_u10_u6_n158, u2_u10_u6_n159, u2_u10_u6_n160, u2_u10_u6_n161, u2_u10_u6_n162, u2_u10_u6_n163, u2_u10_u6_n164, u2_u10_u6_n165, 
       u2_u10_u6_n166, u2_u10_u6_n167, u2_u10_u6_n168, u2_u10_u6_n169, u2_u10_u6_n170, u2_u10_u6_n171, u2_u10_u6_n172, u2_u10_u6_n173, u2_u10_u6_n174, 
       u2_u10_u6_n88, u2_u10_u6_n89, u2_u10_u6_n90, u2_u10_u6_n91, u2_u10_u6_n92, u2_u10_u6_n93, u2_u10_u6_n94, u2_u10_u6_n95, u2_u10_u6_n96, 
       u2_u10_u6_n97, u2_u10_u6_n98, u2_u10_u6_n99, u2_u10_u7_n100, u2_u10_u7_n101, u2_u10_u7_n102, u2_u10_u7_n103, u2_u10_u7_n104, u2_u10_u7_n105, 
       u2_u10_u7_n106, u2_u10_u7_n107, u2_u10_u7_n108, u2_u10_u7_n109, u2_u10_u7_n110, u2_u10_u7_n111, u2_u10_u7_n112, u2_u10_u7_n113, u2_u10_u7_n114, 
       u2_u10_u7_n115, u2_u10_u7_n116, u2_u10_u7_n117, u2_u10_u7_n118, u2_u10_u7_n119, u2_u10_u7_n120, u2_u10_u7_n121, u2_u10_u7_n122, u2_u10_u7_n123, 
       u2_u10_u7_n124, u2_u10_u7_n125, u2_u10_u7_n126, u2_u10_u7_n127, u2_u10_u7_n128, u2_u10_u7_n129, u2_u10_u7_n130, u2_u10_u7_n131, u2_u10_u7_n132, 
       u2_u10_u7_n133, u2_u10_u7_n134, u2_u10_u7_n135, u2_u10_u7_n136, u2_u10_u7_n137, u2_u10_u7_n138, u2_u10_u7_n139, u2_u10_u7_n140, u2_u10_u7_n141, 
       u2_u10_u7_n142, u2_u10_u7_n143, u2_u10_u7_n144, u2_u10_u7_n145, u2_u10_u7_n146, u2_u10_u7_n147, u2_u10_u7_n148, u2_u10_u7_n149, u2_u10_u7_n150, 
       u2_u10_u7_n151, u2_u10_u7_n152, u2_u10_u7_n153, u2_u10_u7_n154, u2_u10_u7_n155, u2_u10_u7_n156, u2_u10_u7_n157, u2_u10_u7_n158, u2_u10_u7_n159, 
       u2_u10_u7_n160, u2_u10_u7_n161, u2_u10_u7_n162, u2_u10_u7_n163, u2_u10_u7_n164, u2_u10_u7_n165, u2_u10_u7_n166, u2_u10_u7_n167, u2_u10_u7_n168, 
       u2_u10_u7_n169, u2_u10_u7_n170, u2_u10_u7_n171, u2_u10_u7_n172, u2_u10_u7_n173, u2_u10_u7_n174, u2_u10_u7_n175, u2_u10_u7_n176, u2_u10_u7_n177, 
       u2_u10_u7_n178, u2_u10_u7_n179, u2_u10_u7_n180, u2_u10_u7_n91, u2_u10_u7_n92, u2_u10_u7_n93, u2_u10_u7_n94, u2_u10_u7_n95, u2_u10_u7_n96, 
       u2_u10_u7_n97, u2_u10_u7_n98, u2_u10_u7_n99, u2_u11_X_19, u2_u11_X_20, u2_u11_X_21, u2_u11_X_22, u2_u11_X_23, u2_u11_X_24, 
       u2_u11_X_25, u2_u11_X_26, u2_u11_X_27, u2_u11_X_28, u2_u11_X_29, u2_u11_X_30, u2_u11_X_31, u2_u11_X_32, u2_u11_X_33, 
       u2_u11_X_34, u2_u11_X_35, u2_u11_X_36, u2_u11_X_37, u2_u11_X_38, u2_u11_X_39, u2_u11_X_40, u2_u11_X_41, u2_u11_X_42, 
       u2_u11_X_43, u2_u11_X_44, u2_u11_X_45, u2_u11_X_46, u2_u11_X_47, u2_u11_X_48, u2_u11_u3_n100, u2_u11_u3_n101, u2_u11_u3_n102, 
       u2_u11_u3_n103, u2_u11_u3_n104, u2_u11_u3_n105, u2_u11_u3_n106, u2_u11_u3_n107, u2_u11_u3_n108, u2_u11_u3_n109, u2_u11_u3_n110, u2_u11_u3_n111, 
       u2_u11_u3_n112, u2_u11_u3_n113, u2_u11_u3_n114, u2_u11_u3_n115, u2_u11_u3_n116, u2_u11_u3_n117, u2_u11_u3_n118, u2_u11_u3_n119, u2_u11_u3_n120, 
       u2_u11_u3_n121, u2_u11_u3_n122, u2_u11_u3_n123, u2_u11_u3_n124, u2_u11_u3_n125, u2_u11_u3_n126, u2_u11_u3_n127, u2_u11_u3_n128, u2_u11_u3_n129, 
       u2_u11_u3_n130, u2_u11_u3_n131, u2_u11_u3_n132, u2_u11_u3_n133, u2_u11_u3_n134, u2_u11_u3_n135, u2_u11_u3_n136, u2_u11_u3_n137, u2_u11_u3_n138, 
       u2_u11_u3_n139, u2_u11_u3_n140, u2_u11_u3_n141, u2_u11_u3_n142, u2_u11_u3_n143, u2_u11_u3_n144, u2_u11_u3_n145, u2_u11_u3_n146, u2_u11_u3_n147, 
       u2_u11_u3_n148, u2_u11_u3_n149, u2_u11_u3_n150, u2_u11_u3_n151, u2_u11_u3_n152, u2_u11_u3_n153, u2_u11_u3_n154, u2_u11_u3_n155, u2_u11_u3_n156, 
       u2_u11_u3_n157, u2_u11_u3_n158, u2_u11_u3_n159, u2_u11_u3_n160, u2_u11_u3_n161, u2_u11_u3_n162, u2_u11_u3_n163, u2_u11_u3_n164, u2_u11_u3_n165, 
       u2_u11_u3_n166, u2_u11_u3_n167, u2_u11_u3_n168, u2_u11_u3_n169, u2_u11_u3_n170, u2_u11_u3_n171, u2_u11_u3_n172, u2_u11_u3_n173, u2_u11_u3_n174, 
       u2_u11_u3_n175, u2_u11_u3_n176, u2_u11_u3_n177, u2_u11_u3_n178, u2_u11_u3_n179, u2_u11_u3_n180, u2_u11_u3_n181, u2_u11_u3_n182, u2_u11_u3_n183, 
       u2_u11_u3_n184, u2_u11_u3_n185, u2_u11_u3_n186, u2_u11_u3_n94, u2_u11_u3_n95, u2_u11_u3_n96, u2_u11_u3_n97, u2_u11_u3_n98, u2_u11_u3_n99, 
       u2_u11_u4_n100, u2_u11_u4_n101, u2_u11_u4_n102, u2_u11_u4_n103, u2_u11_u4_n104, u2_u11_u4_n105, u2_u11_u4_n106, u2_u11_u4_n107, u2_u11_u4_n108, 
       u2_u11_u4_n109, u2_u11_u4_n110, u2_u11_u4_n111, u2_u11_u4_n112, u2_u11_u4_n113, u2_u11_u4_n114, u2_u11_u4_n115, u2_u11_u4_n116, u2_u11_u4_n117, 
       u2_u11_u4_n118, u2_u11_u4_n119, u2_u11_u4_n120, u2_u11_u4_n121, u2_u11_u4_n122, u2_u11_u4_n123, u2_u11_u4_n124, u2_u11_u4_n125, u2_u11_u4_n126, 
       u2_u11_u4_n127, u2_u11_u4_n128, u2_u11_u4_n129, u2_u11_u4_n130, u2_u11_u4_n131, u2_u11_u4_n132, u2_u11_u4_n133, u2_u11_u4_n134, u2_u11_u4_n135, 
       u2_u11_u4_n136, u2_u11_u4_n137, u2_u11_u4_n138, u2_u11_u4_n139, u2_u11_u4_n140, u2_u11_u4_n141, u2_u11_u4_n142, u2_u11_u4_n143, u2_u11_u4_n144, 
       u2_u11_u4_n145, u2_u11_u4_n146, u2_u11_u4_n147, u2_u11_u4_n148, u2_u11_u4_n149, u2_u11_u4_n150, u2_u11_u4_n151, u2_u11_u4_n152, u2_u11_u4_n153, 
       u2_u11_u4_n154, u2_u11_u4_n155, u2_u11_u4_n156, u2_u11_u4_n157, u2_u11_u4_n158, u2_u11_u4_n159, u2_u11_u4_n160, u2_u11_u4_n161, u2_u11_u4_n162, 
       u2_u11_u4_n163, u2_u11_u4_n164, u2_u11_u4_n165, u2_u11_u4_n166, u2_u11_u4_n167, u2_u11_u4_n168, u2_u11_u4_n169, u2_u11_u4_n170, u2_u11_u4_n171, 
       u2_u11_u4_n172, u2_u11_u4_n173, u2_u11_u4_n174, u2_u11_u4_n175, u2_u11_u4_n176, u2_u11_u4_n177, u2_u11_u4_n178, u2_u11_u4_n179, u2_u11_u4_n180, 
       u2_u11_u4_n181, u2_u11_u4_n182, u2_u11_u4_n183, u2_u11_u4_n184, u2_u11_u4_n185, u2_u11_u4_n186, u2_u11_u4_n94, u2_u11_u4_n95, u2_u11_u4_n96, 
       u2_u11_u4_n97, u2_u11_u4_n98, u2_u11_u4_n99, u2_u11_u5_n100, u2_u11_u5_n101, u2_u11_u5_n102, u2_u11_u5_n103, u2_u11_u5_n104, u2_u11_u5_n105, 
       u2_u11_u5_n106, u2_u11_u5_n107, u2_u11_u5_n108, u2_u11_u5_n109, u2_u11_u5_n110, u2_u11_u5_n111, u2_u11_u5_n112, u2_u11_u5_n113, u2_u11_u5_n114, 
       u2_u11_u5_n115, u2_u11_u5_n116, u2_u11_u5_n117, u2_u11_u5_n118, u2_u11_u5_n119, u2_u11_u5_n120, u2_u11_u5_n121, u2_u11_u5_n122, u2_u11_u5_n123, 
       u2_u11_u5_n124, u2_u11_u5_n125, u2_u11_u5_n126, u2_u11_u5_n127, u2_u11_u5_n128, u2_u11_u5_n129, u2_u11_u5_n130, u2_u11_u5_n131, u2_u11_u5_n132, 
       u2_u11_u5_n133, u2_u11_u5_n134, u2_u11_u5_n135, u2_u11_u5_n136, u2_u11_u5_n137, u2_u11_u5_n138, u2_u11_u5_n139, u2_u11_u5_n140, u2_u11_u5_n141, 
       u2_u11_u5_n142, u2_u11_u5_n143, u2_u11_u5_n144, u2_u11_u5_n145, u2_u11_u5_n146, u2_u11_u5_n147, u2_u11_u5_n148, u2_u11_u5_n149, u2_u11_u5_n150, 
       u2_u11_u5_n151, u2_u11_u5_n152, u2_u11_u5_n153, u2_u11_u5_n154, u2_u11_u5_n155, u2_u11_u5_n156, u2_u11_u5_n157, u2_u11_u5_n158, u2_u11_u5_n159, 
       u2_u11_u5_n160, u2_u11_u5_n161, u2_u11_u5_n162, u2_u11_u5_n163, u2_u11_u5_n164, u2_u11_u5_n165, u2_u11_u5_n166, u2_u11_u5_n167, u2_u11_u5_n168, 
       u2_u11_u5_n169, u2_u11_u5_n170, u2_u11_u5_n171, u2_u11_u5_n172, u2_u11_u5_n173, u2_u11_u5_n174, u2_u11_u5_n175, u2_u11_u5_n176, u2_u11_u5_n177, 
       u2_u11_u5_n178, u2_u11_u5_n179, u2_u11_u5_n180, u2_u11_u5_n181, u2_u11_u5_n182, u2_u11_u5_n183, u2_u11_u5_n184, u2_u11_u5_n185, u2_u11_u5_n186, 
       u2_u11_u5_n187, u2_u11_u5_n188, u2_u11_u5_n189, u2_u11_u5_n190, u2_u11_u5_n191, u2_u11_u5_n192, u2_u11_u5_n193, u2_u11_u5_n194, u2_u11_u5_n195, 
       u2_u11_u5_n196, u2_u11_u5_n99, u2_u11_u6_n100, u2_u11_u6_n101, u2_u11_u6_n102, u2_u11_u6_n103, u2_u11_u6_n104, u2_u11_u6_n105, u2_u11_u6_n106, 
       u2_u11_u6_n107, u2_u11_u6_n108, u2_u11_u6_n109, u2_u11_u6_n110, u2_u11_u6_n111, u2_u11_u6_n112, u2_u11_u6_n113, u2_u11_u6_n114, u2_u11_u6_n115, 
       u2_u11_u6_n116, u2_u11_u6_n117, u2_u11_u6_n118, u2_u11_u6_n119, u2_u11_u6_n120, u2_u11_u6_n121, u2_u11_u6_n122, u2_u11_u6_n123, u2_u11_u6_n124, 
       u2_u11_u6_n125, u2_u11_u6_n126, u2_u11_u6_n127, u2_u11_u6_n128, u2_u11_u6_n129, u2_u11_u6_n130, u2_u11_u6_n131, u2_u11_u6_n132, u2_u11_u6_n133, 
       u2_u11_u6_n134, u2_u11_u6_n135, u2_u11_u6_n136, u2_u11_u6_n137, u2_u11_u6_n138, u2_u11_u6_n139, u2_u11_u6_n140, u2_u11_u6_n141, u2_u11_u6_n142, 
       u2_u11_u6_n143, u2_u11_u6_n144, u2_u11_u6_n145, u2_u11_u6_n146, u2_u11_u6_n147, u2_u11_u6_n148, u2_u11_u6_n149, u2_u11_u6_n150, u2_u11_u6_n151, 
       u2_u11_u6_n152, u2_u11_u6_n153, u2_u11_u6_n154, u2_u11_u6_n155, u2_u11_u6_n156, u2_u11_u6_n157, u2_u11_u6_n158, u2_u11_u6_n159, u2_u11_u6_n160, 
       u2_u11_u6_n161, u2_u11_u6_n162, u2_u11_u6_n163, u2_u11_u6_n164, u2_u11_u6_n165, u2_u11_u6_n166, u2_u11_u6_n167, u2_u11_u6_n168, u2_u11_u6_n169, 
       u2_u11_u6_n170, u2_u11_u6_n171, u2_u11_u6_n172, u2_u11_u6_n173, u2_u11_u6_n174, u2_u11_u6_n88, u2_u11_u6_n89, u2_u11_u6_n90, u2_u11_u6_n91, 
       u2_u11_u6_n92, u2_u11_u6_n93, u2_u11_u6_n94, u2_u11_u6_n95, u2_u11_u6_n96, u2_u11_u6_n97, u2_u11_u6_n98, u2_u11_u6_n99, u2_u11_u7_n100, 
       u2_u11_u7_n101, u2_u11_u7_n102, u2_u11_u7_n103, u2_u11_u7_n104, u2_u11_u7_n105, u2_u11_u7_n106, u2_u11_u7_n107, u2_u11_u7_n108, u2_u11_u7_n109, 
       u2_u11_u7_n110, u2_u11_u7_n111, u2_u11_u7_n112, u2_u11_u7_n113, u2_u11_u7_n114, u2_u11_u7_n115, u2_u11_u7_n116, u2_u11_u7_n117, u2_u11_u7_n118, 
       u2_u11_u7_n119, u2_u11_u7_n120, u2_u11_u7_n121, u2_u11_u7_n122, u2_u11_u7_n123, u2_u11_u7_n124, u2_u11_u7_n125, u2_u11_u7_n126, u2_u11_u7_n127, 
       u2_u11_u7_n128, u2_u11_u7_n129, u2_u11_u7_n130, u2_u11_u7_n131, u2_u11_u7_n132, u2_u11_u7_n133, u2_u11_u7_n134, u2_u11_u7_n135, u2_u11_u7_n136, 
       u2_u11_u7_n137, u2_u11_u7_n138, u2_u11_u7_n139, u2_u11_u7_n140, u2_u11_u7_n141, u2_u11_u7_n142, u2_u11_u7_n143, u2_u11_u7_n144, u2_u11_u7_n145, 
       u2_u11_u7_n146, u2_u11_u7_n147, u2_u11_u7_n148, u2_u11_u7_n149, u2_u11_u7_n150, u2_u11_u7_n151, u2_u11_u7_n152, u2_u11_u7_n153, u2_u11_u7_n154, 
       u2_u11_u7_n155, u2_u11_u7_n156, u2_u11_u7_n157, u2_u11_u7_n158, u2_u11_u7_n159, u2_u11_u7_n160, u2_u11_u7_n161, u2_u11_u7_n162, u2_u11_u7_n163, 
       u2_u11_u7_n164, u2_u11_u7_n165, u2_u11_u7_n166, u2_u11_u7_n167, u2_u11_u7_n168, u2_u11_u7_n169, u2_u11_u7_n170, u2_u11_u7_n171, u2_u11_u7_n172, 
       u2_u11_u7_n173, u2_u11_u7_n174, u2_u11_u7_n175, u2_u11_u7_n176, u2_u11_u7_n177, u2_u11_u7_n178, u2_u11_u7_n179, u2_u11_u7_n180, u2_u11_u7_n91, 
       u2_u11_u7_n92, u2_u11_u7_n93, u2_u11_u7_n94, u2_u11_u7_n95, u2_u11_u7_n96, u2_u11_u7_n97, u2_u11_u7_n98, u2_u11_u7_n99, u2_u12_X_1, 
       u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_13, u2_u12_X_14, u2_u12_X_15, u2_u12_X_16, u2_u12_X_17, u2_u12_X_18, 
       u2_u12_X_19, u2_u12_X_2, u2_u12_X_20, u2_u12_X_21, u2_u12_X_22, u2_u12_X_23, u2_u12_X_24, u2_u12_X_25, u2_u12_X_26, 
       u2_u12_X_27, u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, u2_u12_X_30, u2_u12_X_31, u2_u12_X_32, u2_u12_X_33, u2_u12_X_34, 
       u2_u12_X_35, u2_u12_X_36, u2_u12_X_4, u2_u12_X_5, u2_u12_X_6, u2_u12_X_7, u2_u12_X_8, u2_u12_X_9, u2_u12_u0_n100, 
       u2_u12_u0_n101, u2_u12_u0_n102, u2_u12_u0_n103, u2_u12_u0_n104, u2_u12_u0_n105, u2_u12_u0_n106, u2_u12_u0_n107, u2_u12_u0_n108, u2_u12_u0_n109, 
       u2_u12_u0_n110, u2_u12_u0_n111, u2_u12_u0_n112, u2_u12_u0_n113, u2_u12_u0_n114, u2_u12_u0_n115, u2_u12_u0_n116, u2_u12_u0_n117, u2_u12_u0_n118, 
       u2_u12_u0_n119, u2_u12_u0_n120, u2_u12_u0_n121, u2_u12_u0_n122, u2_u12_u0_n123, u2_u12_u0_n124, u2_u12_u0_n125, u2_u12_u0_n126, u2_u12_u0_n127, 
       u2_u12_u0_n128, u2_u12_u0_n129, u2_u12_u0_n130, u2_u12_u0_n131, u2_u12_u0_n132, u2_u12_u0_n133, u2_u12_u0_n134, u2_u12_u0_n135, u2_u12_u0_n136, 
       u2_u12_u0_n137, u2_u12_u0_n138, u2_u12_u0_n139, u2_u12_u0_n140, u2_u12_u0_n141, u2_u12_u0_n142, u2_u12_u0_n143, u2_u12_u0_n144, u2_u12_u0_n145, 
       u2_u12_u0_n146, u2_u12_u0_n147, u2_u12_u0_n148, u2_u12_u0_n149, u2_u12_u0_n150, u2_u12_u0_n151, u2_u12_u0_n152, u2_u12_u0_n153, u2_u12_u0_n154, 
       u2_u12_u0_n155, u2_u12_u0_n156, u2_u12_u0_n157, u2_u12_u0_n158, u2_u12_u0_n159, u2_u12_u0_n160, u2_u12_u0_n161, u2_u12_u0_n162, u2_u12_u0_n163, 
       u2_u12_u0_n164, u2_u12_u0_n165, u2_u12_u0_n166, u2_u12_u0_n167, u2_u12_u0_n168, u2_u12_u0_n169, u2_u12_u0_n170, u2_u12_u0_n171, u2_u12_u0_n172, 
       u2_u12_u0_n173, u2_u12_u0_n174, u2_u12_u0_n88, u2_u12_u0_n89, u2_u12_u0_n90, u2_u12_u0_n91, u2_u12_u0_n92, u2_u12_u0_n93, u2_u12_u0_n94, 
       u2_u12_u0_n95, u2_u12_u0_n96, u2_u12_u0_n97, u2_u12_u0_n98, u2_u12_u0_n99, u2_u12_u1_n100, u2_u12_u1_n101, u2_u12_u1_n102, u2_u12_u1_n103, 
       u2_u12_u1_n104, u2_u12_u1_n105, u2_u12_u1_n106, u2_u12_u1_n107, u2_u12_u1_n108, u2_u12_u1_n109, u2_u12_u1_n110, u2_u12_u1_n111, u2_u12_u1_n112, 
       u2_u12_u1_n113, u2_u12_u1_n114, u2_u12_u1_n115, u2_u12_u1_n116, u2_u12_u1_n117, u2_u12_u1_n118, u2_u12_u1_n119, u2_u12_u1_n120, u2_u12_u1_n121, 
       u2_u12_u1_n122, u2_u12_u1_n123, u2_u12_u1_n124, u2_u12_u1_n125, u2_u12_u1_n126, u2_u12_u1_n127, u2_u12_u1_n128, u2_u12_u1_n129, u2_u12_u1_n130, 
       u2_u12_u1_n131, u2_u12_u1_n132, u2_u12_u1_n133, u2_u12_u1_n134, u2_u12_u1_n135, u2_u12_u1_n136, u2_u12_u1_n137, u2_u12_u1_n138, u2_u12_u1_n139, 
       u2_u12_u1_n140, u2_u12_u1_n141, u2_u12_u1_n142, u2_u12_u1_n143, u2_u12_u1_n144, u2_u12_u1_n145, u2_u12_u1_n146, u2_u12_u1_n147, u2_u12_u1_n148, 
       u2_u12_u1_n149, u2_u12_u1_n150, u2_u12_u1_n151, u2_u12_u1_n152, u2_u12_u1_n153, u2_u12_u1_n154, u2_u12_u1_n155, u2_u12_u1_n156, u2_u12_u1_n157, 
       u2_u12_u1_n158, u2_u12_u1_n159, u2_u12_u1_n160, u2_u12_u1_n161, u2_u12_u1_n162, u2_u12_u1_n163, u2_u12_u1_n164, u2_u12_u1_n165, u2_u12_u1_n166, 
       u2_u12_u1_n167, u2_u12_u1_n168, u2_u12_u1_n169, u2_u12_u1_n170, u2_u12_u1_n171, u2_u12_u1_n172, u2_u12_u1_n173, u2_u12_u1_n174, u2_u12_u1_n175, 
       u2_u12_u1_n176, u2_u12_u1_n177, u2_u12_u1_n178, u2_u12_u1_n179, u2_u12_u1_n180, u2_u12_u1_n181, u2_u12_u1_n182, u2_u12_u1_n183, u2_u12_u1_n184, 
       u2_u12_u1_n185, u2_u12_u1_n186, u2_u12_u1_n187, u2_u12_u1_n188, u2_u12_u1_n95, u2_u12_u1_n96, u2_u12_u1_n97, u2_u12_u1_n98, u2_u12_u1_n99, 
       u2_u12_u2_n100, u2_u12_u2_n101, u2_u12_u2_n102, u2_u12_u2_n103, u2_u12_u2_n104, u2_u12_u2_n105, u2_u12_u2_n106, u2_u12_u2_n107, u2_u12_u2_n108, 
       u2_u12_u2_n109, u2_u12_u2_n110, u2_u12_u2_n111, u2_u12_u2_n112, u2_u12_u2_n113, u2_u12_u2_n114, u2_u12_u2_n115, u2_u12_u2_n116, u2_u12_u2_n117, 
       u2_u12_u2_n118, u2_u12_u2_n119, u2_u12_u2_n120, u2_u12_u2_n121, u2_u12_u2_n122, u2_u12_u2_n123, u2_u12_u2_n124, u2_u12_u2_n125, u2_u12_u2_n126, 
       u2_u12_u2_n127, u2_u12_u2_n128, u2_u12_u2_n129, u2_u12_u2_n130, u2_u12_u2_n131, u2_u12_u2_n132, u2_u12_u2_n133, u2_u12_u2_n134, u2_u12_u2_n135, 
       u2_u12_u2_n136, u2_u12_u2_n137, u2_u12_u2_n138, u2_u12_u2_n139, u2_u12_u2_n140, u2_u12_u2_n141, u2_u12_u2_n142, u2_u12_u2_n143, u2_u12_u2_n144, 
       u2_u12_u2_n145, u2_u12_u2_n146, u2_u12_u2_n147, u2_u12_u2_n148, u2_u12_u2_n149, u2_u12_u2_n150, u2_u12_u2_n151, u2_u12_u2_n152, u2_u12_u2_n153, 
       u2_u12_u2_n154, u2_u12_u2_n155, u2_u12_u2_n156, u2_u12_u2_n157, u2_u12_u2_n158, u2_u12_u2_n159, u2_u12_u2_n160, u2_u12_u2_n161, u2_u12_u2_n162, 
       u2_u12_u2_n163, u2_u12_u2_n164, u2_u12_u2_n165, u2_u12_u2_n166, u2_u12_u2_n167, u2_u12_u2_n168, u2_u12_u2_n169, u2_u12_u2_n170, u2_u12_u2_n171, 
       u2_u12_u2_n172, u2_u12_u2_n173, u2_u12_u2_n174, u2_u12_u2_n175, u2_u12_u2_n176, u2_u12_u2_n177, u2_u12_u2_n178, u2_u12_u2_n179, u2_u12_u2_n180, 
       u2_u12_u2_n181, u2_u12_u2_n182, u2_u12_u2_n183, u2_u12_u2_n184, u2_u12_u2_n185, u2_u12_u2_n186, u2_u12_u2_n187, u2_u12_u2_n188, u2_u12_u2_n95, 
       u2_u12_u2_n96, u2_u12_u2_n97, u2_u12_u2_n98, u2_u12_u2_n99, u2_u12_u3_n100, u2_u12_u3_n101, u2_u12_u3_n102, u2_u12_u3_n103, u2_u12_u3_n104, 
       u2_u12_u3_n105, u2_u12_u3_n106, u2_u12_u3_n107, u2_u12_u3_n108, u2_u12_u3_n109, u2_u12_u3_n110, u2_u12_u3_n111, u2_u12_u3_n112, u2_u12_u3_n113, 
       u2_u12_u3_n114, u2_u12_u3_n115, u2_u12_u3_n116, u2_u12_u3_n117, u2_u12_u3_n118, u2_u12_u3_n119, u2_u12_u3_n120, u2_u12_u3_n121, u2_u12_u3_n122, 
       u2_u12_u3_n123, u2_u12_u3_n124, u2_u12_u3_n125, u2_u12_u3_n126, u2_u12_u3_n127, u2_u12_u3_n128, u2_u12_u3_n129, u2_u12_u3_n130, u2_u12_u3_n131, 
       u2_u12_u3_n132, u2_u12_u3_n133, u2_u12_u3_n134, u2_u12_u3_n135, u2_u12_u3_n136, u2_u12_u3_n137, u2_u12_u3_n138, u2_u12_u3_n139, u2_u12_u3_n140, 
       u2_u12_u3_n141, u2_u12_u3_n142, u2_u12_u3_n143, u2_u12_u3_n144, u2_u12_u3_n145, u2_u12_u3_n146, u2_u12_u3_n147, u2_u12_u3_n148, u2_u12_u3_n149, 
       u2_u12_u3_n150, u2_u12_u3_n151, u2_u12_u3_n152, u2_u12_u3_n153, u2_u12_u3_n154, u2_u12_u3_n155, u2_u12_u3_n156, u2_u12_u3_n157, u2_u12_u3_n158, 
       u2_u12_u3_n159, u2_u12_u3_n160, u2_u12_u3_n161, u2_u12_u3_n162, u2_u12_u3_n163, u2_u12_u3_n164, u2_u12_u3_n165, u2_u12_u3_n166, u2_u12_u3_n167, 
       u2_u12_u3_n168, u2_u12_u3_n169, u2_u12_u3_n170, u2_u12_u3_n171, u2_u12_u3_n172, u2_u12_u3_n173, u2_u12_u3_n174, u2_u12_u3_n175, u2_u12_u3_n176, 
       u2_u12_u3_n177, u2_u12_u3_n178, u2_u12_u3_n179, u2_u12_u3_n180, u2_u12_u3_n181, u2_u12_u3_n182, u2_u12_u3_n183, u2_u12_u3_n184, u2_u12_u3_n185, 
       u2_u12_u3_n186, u2_u12_u3_n94, u2_u12_u3_n95, u2_u12_u3_n96, u2_u12_u3_n97, u2_u12_u3_n98, u2_u12_u3_n99, u2_u12_u4_n100, u2_u12_u4_n101, 
       u2_u12_u4_n102, u2_u12_u4_n103, u2_u12_u4_n104, u2_u12_u4_n105, u2_u12_u4_n106, u2_u12_u4_n107, u2_u12_u4_n108, u2_u12_u4_n109, u2_u12_u4_n110, 
       u2_u12_u4_n111, u2_u12_u4_n112, u2_u12_u4_n113, u2_u12_u4_n114, u2_u12_u4_n115, u2_u12_u4_n116, u2_u12_u4_n117, u2_u12_u4_n118, u2_u12_u4_n119, 
       u2_u12_u4_n120, u2_u12_u4_n121, u2_u12_u4_n122, u2_u12_u4_n123, u2_u12_u4_n124, u2_u12_u4_n125, u2_u12_u4_n126, u2_u12_u4_n127, u2_u12_u4_n128, 
       u2_u12_u4_n129, u2_u12_u4_n130, u2_u12_u4_n131, u2_u12_u4_n132, u2_u12_u4_n133, u2_u12_u4_n134, u2_u12_u4_n135, u2_u12_u4_n136, u2_u12_u4_n137, 
       u2_u12_u4_n138, u2_u12_u4_n139, u2_u12_u4_n140, u2_u12_u4_n141, u2_u12_u4_n142, u2_u12_u4_n143, u2_u12_u4_n144, u2_u12_u4_n145, u2_u12_u4_n146, 
       u2_u12_u4_n147, u2_u12_u4_n148, u2_u12_u4_n149, u2_u12_u4_n150, u2_u12_u4_n151, u2_u12_u4_n152, u2_u12_u4_n153, u2_u12_u4_n154, u2_u12_u4_n155, 
       u2_u12_u4_n156, u2_u12_u4_n157, u2_u12_u4_n158, u2_u12_u4_n159, u2_u12_u4_n160, u2_u12_u4_n161, u2_u12_u4_n162, u2_u12_u4_n163, u2_u12_u4_n164, 
       u2_u12_u4_n165, u2_u12_u4_n166, u2_u12_u4_n167, u2_u12_u4_n168, u2_u12_u4_n169, u2_u12_u4_n170, u2_u12_u4_n171, u2_u12_u4_n172, u2_u12_u4_n173, 
       u2_u12_u4_n174, u2_u12_u4_n175, u2_u12_u4_n176, u2_u12_u4_n177, u2_u12_u4_n178, u2_u12_u4_n179, u2_u12_u4_n180, u2_u12_u4_n181, u2_u12_u4_n182, 
       u2_u12_u4_n183, u2_u12_u4_n184, u2_u12_u4_n185, u2_u12_u4_n186, u2_u12_u4_n94, u2_u12_u4_n95, u2_u12_u4_n96, u2_u12_u4_n97, u2_u12_u4_n98, 
       u2_u12_u4_n99, u2_u12_u5_n100, u2_u12_u5_n101, u2_u12_u5_n102, u2_u12_u5_n103, u2_u12_u5_n104, u2_u12_u5_n105, u2_u12_u5_n106, u2_u12_u5_n107, 
       u2_u12_u5_n108, u2_u12_u5_n109, u2_u12_u5_n110, u2_u12_u5_n111, u2_u12_u5_n112, u2_u12_u5_n113, u2_u12_u5_n114, u2_u12_u5_n115, u2_u12_u5_n116, 
       u2_u12_u5_n117, u2_u12_u5_n118, u2_u12_u5_n119, u2_u12_u5_n120, u2_u12_u5_n121, u2_u12_u5_n122, u2_u12_u5_n123, u2_u12_u5_n124, u2_u12_u5_n125, 
       u2_u12_u5_n126, u2_u12_u5_n127, u2_u12_u5_n128, u2_u12_u5_n129, u2_u12_u5_n130, u2_u12_u5_n131, u2_u12_u5_n132, u2_u12_u5_n133, u2_u12_u5_n134, 
       u2_u12_u5_n135, u2_u12_u5_n136, u2_u12_u5_n137, u2_u12_u5_n138, u2_u12_u5_n139, u2_u12_u5_n140, u2_u12_u5_n141, u2_u12_u5_n142, u2_u12_u5_n143, 
       u2_u12_u5_n144, u2_u12_u5_n145, u2_u12_u5_n146, u2_u12_u5_n147, u2_u12_u5_n148, u2_u12_u5_n149, u2_u12_u5_n150, u2_u12_u5_n151, u2_u12_u5_n152, 
       u2_u12_u5_n153, u2_u12_u5_n154, u2_u12_u5_n155, u2_u12_u5_n156, u2_u12_u5_n157, u2_u12_u5_n158, u2_u12_u5_n159, u2_u12_u5_n160, u2_u12_u5_n161, 
       u2_u12_u5_n162, u2_u12_u5_n163, u2_u12_u5_n164, u2_u12_u5_n165, u2_u12_u5_n166, u2_u12_u5_n167, u2_u12_u5_n168, u2_u12_u5_n169, u2_u12_u5_n170, 
       u2_u12_u5_n171, u2_u12_u5_n172, u2_u12_u5_n173, u2_u12_u5_n174, u2_u12_u5_n175, u2_u12_u5_n176, u2_u12_u5_n177, u2_u12_u5_n178, u2_u12_u5_n179, 
       u2_u12_u5_n180, u2_u12_u5_n181, u2_u12_u5_n182, u2_u12_u5_n183, u2_u12_u5_n184, u2_u12_u5_n185, u2_u12_u5_n186, u2_u12_u5_n187, u2_u12_u5_n188, 
       u2_u12_u5_n189, u2_u12_u5_n190, u2_u12_u5_n191, u2_u12_u5_n192, u2_u12_u5_n193, u2_u12_u5_n194, u2_u12_u5_n195, u2_u12_u5_n196, u2_u12_u5_n99, 
       u2_u14_X_13, u2_u14_X_14, u2_u14_X_15, u2_u14_X_16, u2_u14_X_17, u2_u14_X_18, u2_u14_X_19, u2_u14_X_20, u2_u14_X_21, 
       u2_u14_X_22, u2_u14_X_23, u2_u14_X_24, u2_u14_X_43, u2_u14_X_44, u2_u14_X_45, u2_u14_X_46, u2_u14_X_47, u2_u14_X_48, 
       u2_u14_u2_n100, u2_u14_u2_n101, u2_u14_u2_n102, u2_u14_u2_n103, u2_u14_u2_n104, u2_u14_u2_n105, u2_u14_u2_n106, u2_u14_u2_n107, u2_u14_u2_n108, 
       u2_u14_u2_n109, u2_u14_u2_n110, u2_u14_u2_n111, u2_u14_u2_n112, u2_u14_u2_n113, u2_u14_u2_n114, u2_u14_u2_n115, u2_u14_u2_n116, u2_u14_u2_n117, 
       u2_u14_u2_n118, u2_u14_u2_n119, u2_u14_u2_n120, u2_u14_u2_n121, u2_u14_u2_n122, u2_u14_u2_n123, u2_u14_u2_n124, u2_u14_u2_n125, u2_u14_u2_n126, 
       u2_u14_u2_n127, u2_u14_u2_n128, u2_u14_u2_n129, u2_u14_u2_n130, u2_u14_u2_n131, u2_u14_u2_n132, u2_u14_u2_n133, u2_u14_u2_n134, u2_u14_u2_n135, 
       u2_u14_u2_n136, u2_u14_u2_n137, u2_u14_u2_n138, u2_u14_u2_n139, u2_u14_u2_n140, u2_u14_u2_n141, u2_u14_u2_n142, u2_u14_u2_n143, u2_u14_u2_n144, 
       u2_u14_u2_n145, u2_u14_u2_n146, u2_u14_u2_n147, u2_u14_u2_n148, u2_u14_u2_n149, u2_u14_u2_n150, u2_u14_u2_n151, u2_u14_u2_n152, u2_u14_u2_n153, 
       u2_u14_u2_n154, u2_u14_u2_n155, u2_u14_u2_n156, u2_u14_u2_n157, u2_u14_u2_n158, u2_u14_u2_n159, u2_u14_u2_n160, u2_u14_u2_n161, u2_u14_u2_n162, 
       u2_u14_u2_n163, u2_u14_u2_n164, u2_u14_u2_n165, u2_u14_u2_n166, u2_u14_u2_n167, u2_u14_u2_n168, u2_u14_u2_n169, u2_u14_u2_n170, u2_u14_u2_n171, 
       u2_u14_u2_n172, u2_u14_u2_n173, u2_u14_u2_n174, u2_u14_u2_n175, u2_u14_u2_n176, u2_u14_u2_n177, u2_u14_u2_n178, u2_u14_u2_n179, u2_u14_u2_n180, 
       u2_u14_u2_n181, u2_u14_u2_n182, u2_u14_u2_n183, u2_u14_u2_n184, u2_u14_u2_n185, u2_u14_u2_n186, u2_u14_u2_n187, u2_u14_u2_n188, u2_u14_u2_n95, 
       u2_u14_u2_n96, u2_u14_u2_n97, u2_u14_u2_n98, u2_u14_u2_n99, u2_u14_u3_n100, u2_u14_u3_n101, u2_u14_u3_n102, u2_u14_u3_n103, u2_u14_u3_n104, 
       u2_u14_u3_n105, u2_u14_u3_n106, u2_u14_u3_n107, u2_u14_u3_n108, u2_u14_u3_n109, u2_u14_u3_n110, u2_u14_u3_n111, u2_u14_u3_n112, u2_u14_u3_n113, 
       u2_u14_u3_n114, u2_u14_u3_n115, u2_u14_u3_n116, u2_u14_u3_n117, u2_u14_u3_n118, u2_u14_u3_n119, u2_u14_u3_n120, u2_u14_u3_n121, u2_u14_u3_n122, 
       u2_u14_u3_n123, u2_u14_u3_n124, u2_u14_u3_n125, u2_u14_u3_n126, u2_u14_u3_n127, u2_u14_u3_n128, u2_u14_u3_n129, u2_u14_u3_n130, u2_u14_u3_n131, 
       u2_u14_u3_n132, u2_u14_u3_n133, u2_u14_u3_n134, u2_u14_u3_n135, u2_u14_u3_n136, u2_u14_u3_n137, u2_u14_u3_n138, u2_u14_u3_n139, u2_u14_u3_n140, 
       u2_u14_u3_n141, u2_u14_u3_n142, u2_u14_u3_n143, u2_u14_u3_n144, u2_u14_u3_n145, u2_u14_u3_n146, u2_u14_u3_n147, u2_u14_u3_n148, u2_u14_u3_n149, 
       u2_u14_u3_n150, u2_u14_u3_n151, u2_u14_u3_n152, u2_u14_u3_n153, u2_u14_u3_n154, u2_u14_u3_n155, u2_u14_u3_n156, u2_u14_u3_n157, u2_u14_u3_n158, 
       u2_u14_u3_n159, u2_u14_u3_n160, u2_u14_u3_n161, u2_u14_u3_n162, u2_u14_u3_n163, u2_u14_u3_n164, u2_u14_u3_n165, u2_u14_u3_n166, u2_u14_u3_n167, 
       u2_u14_u3_n168, u2_u14_u3_n169, u2_u14_u3_n170, u2_u14_u3_n171, u2_u14_u3_n172, u2_u14_u3_n173, u2_u14_u3_n174, u2_u14_u3_n175, u2_u14_u3_n176, 
       u2_u14_u3_n177, u2_u14_u3_n178, u2_u14_u3_n179, u2_u14_u3_n180, u2_u14_u3_n181, u2_u14_u3_n182, u2_u14_u3_n183, u2_u14_u3_n184, u2_u14_u3_n185, 
       u2_u14_u3_n186, u2_u14_u3_n94, u2_u14_u3_n95, u2_u14_u3_n96, u2_u14_u3_n97, u2_u14_u3_n98, u2_u14_u3_n99, u2_u14_u7_n100, u2_u14_u7_n101, 
       u2_u14_u7_n102, u2_u14_u7_n103, u2_u14_u7_n104, u2_u14_u7_n105, u2_u14_u7_n106, u2_u14_u7_n107, u2_u14_u7_n108, u2_u14_u7_n109, u2_u14_u7_n110, 
       u2_u14_u7_n111, u2_u14_u7_n112, u2_u14_u7_n113, u2_u14_u7_n114, u2_u14_u7_n115, u2_u14_u7_n116, u2_u14_u7_n117, u2_u14_u7_n118, u2_u14_u7_n119, 
       u2_u14_u7_n120, u2_u14_u7_n121, u2_u14_u7_n122, u2_u14_u7_n123, u2_u14_u7_n124, u2_u14_u7_n125, u2_u14_u7_n126, u2_u14_u7_n127, u2_u14_u7_n128, 
       u2_u14_u7_n129, u2_u14_u7_n130, u2_u14_u7_n131, u2_u14_u7_n132, u2_u14_u7_n133, u2_u14_u7_n134, u2_u14_u7_n135, u2_u14_u7_n136, u2_u14_u7_n137, 
       u2_u14_u7_n138, u2_u14_u7_n139, u2_u14_u7_n140, u2_u14_u7_n141, u2_u14_u7_n142, u2_u14_u7_n143, u2_u14_u7_n144, u2_u14_u7_n145, u2_u14_u7_n146, 
       u2_u14_u7_n147, u2_u14_u7_n148, u2_u14_u7_n149, u2_u14_u7_n150, u2_u14_u7_n151, u2_u14_u7_n152, u2_u14_u7_n153, u2_u14_u7_n154, u2_u14_u7_n155, 
       u2_u14_u7_n156, u2_u14_u7_n157, u2_u14_u7_n158, u2_u14_u7_n159, u2_u14_u7_n160, u2_u14_u7_n161, u2_u14_u7_n162, u2_u14_u7_n163, u2_u14_u7_n164, 
       u2_u14_u7_n165, u2_u14_u7_n166, u2_u14_u7_n167, u2_u14_u7_n168, u2_u14_u7_n169, u2_u14_u7_n170, u2_u14_u7_n171, u2_u14_u7_n172, u2_u14_u7_n173, 
       u2_u14_u7_n174, u2_u14_u7_n175, u2_u14_u7_n176, u2_u14_u7_n177, u2_u14_u7_n178, u2_u14_u7_n179, u2_u14_u7_n180, u2_u14_u7_n91, u2_u14_u7_n92, 
       u2_u14_u7_n93, u2_u14_u7_n94, u2_u14_u7_n95, u2_u14_u7_n96, u2_u14_u7_n97, u2_u14_u7_n98, u2_u14_u7_n99, u2_u15_X_10, u2_u15_X_11, 
       u2_u15_X_12, u2_u15_X_13, u2_u15_X_14, u2_u15_X_15, u2_u15_X_16, u2_u15_X_17, u2_u15_X_18, u2_u15_X_19, u2_u15_X_20, 
       u2_u15_X_21, u2_u15_X_22, u2_u15_X_23, u2_u15_X_24, u2_u15_X_7, u2_u15_X_8, u2_u15_X_9, u2_u15_u1_n100, u2_u15_u1_n101, 
       u2_u15_u1_n102, u2_u15_u1_n103, u2_u15_u1_n104, u2_u15_u1_n105, u2_u15_u1_n106, u2_u15_u1_n107, u2_u15_u1_n108, u2_u15_u1_n109, u2_u15_u1_n110, 
       u2_u15_u1_n111, u2_u15_u1_n112, u2_u15_u1_n113, u2_u15_u1_n114, u2_u15_u1_n115, u2_u15_u1_n116, u2_u15_u1_n117, u2_u15_u1_n118, u2_u15_u1_n119, 
       u2_u15_u1_n120, u2_u15_u1_n121, u2_u15_u1_n122, u2_u15_u1_n123, u2_u15_u1_n124, u2_u15_u1_n125, u2_u15_u1_n126, u2_u15_u1_n127, u2_u15_u1_n128, 
       u2_u15_u1_n129, u2_u15_u1_n130, u2_u15_u1_n131, u2_u15_u1_n132, u2_u15_u1_n133, u2_u15_u1_n134, u2_u15_u1_n135, u2_u15_u1_n136, u2_u15_u1_n137, 
       u2_u15_u1_n138, u2_u15_u1_n139, u2_u15_u1_n140, u2_u15_u1_n141, u2_u15_u1_n142, u2_u15_u1_n143, u2_u15_u1_n144, u2_u15_u1_n145, u2_u15_u1_n146, 
       u2_u15_u1_n147, u2_u15_u1_n148, u2_u15_u1_n149, u2_u15_u1_n150, u2_u15_u1_n151, u2_u15_u1_n152, u2_u15_u1_n153, u2_u15_u1_n154, u2_u15_u1_n155, 
       u2_u15_u1_n156, u2_u15_u1_n157, u2_u15_u1_n158, u2_u15_u1_n159, u2_u15_u1_n160, u2_u15_u1_n161, u2_u15_u1_n162, u2_u15_u1_n163, u2_u15_u1_n164, 
       u2_u15_u1_n165, u2_u15_u1_n166, u2_u15_u1_n167, u2_u15_u1_n168, u2_u15_u1_n169, u2_u15_u1_n170, u2_u15_u1_n171, u2_u15_u1_n172, u2_u15_u1_n173, 
       u2_u15_u1_n174, u2_u15_u1_n175, u2_u15_u1_n176, u2_u15_u1_n177, u2_u15_u1_n178, u2_u15_u1_n179, u2_u15_u1_n180, u2_u15_u1_n181, u2_u15_u1_n182, 
       u2_u15_u1_n183, u2_u15_u1_n184, u2_u15_u1_n185, u2_u15_u1_n186, u2_u15_u1_n187, u2_u15_u1_n188, u2_u15_u1_n95, u2_u15_u1_n96, u2_u15_u1_n97, 
       u2_u15_u1_n98, u2_u15_u1_n99, u2_u15_u2_n100, u2_u15_u2_n101, u2_u15_u2_n102, u2_u15_u2_n103, u2_u15_u2_n104, u2_u15_u2_n105, u2_u15_u2_n106, 
       u2_u15_u2_n107, u2_u15_u2_n108, u2_u15_u2_n109, u2_u15_u2_n110, u2_u15_u2_n111, u2_u15_u2_n112, u2_u15_u2_n113, u2_u15_u2_n114, u2_u15_u2_n115, 
       u2_u15_u2_n116, u2_u15_u2_n117, u2_u15_u2_n118, u2_u15_u2_n119, u2_u15_u2_n120, u2_u15_u2_n121, u2_u15_u2_n122, u2_u15_u2_n123, u2_u15_u2_n124, 
       u2_u15_u2_n125, u2_u15_u2_n126, u2_u15_u2_n127, u2_u15_u2_n128, u2_u15_u2_n129, u2_u15_u2_n130, u2_u15_u2_n131, u2_u15_u2_n132, u2_u15_u2_n133, 
       u2_u15_u2_n134, u2_u15_u2_n135, u2_u15_u2_n136, u2_u15_u2_n137, u2_u15_u2_n138, u2_u15_u2_n139, u2_u15_u2_n140, u2_u15_u2_n141, u2_u15_u2_n142, 
       u2_u15_u2_n143, u2_u15_u2_n144, u2_u15_u2_n145, u2_u15_u2_n146, u2_u15_u2_n147, u2_u15_u2_n148, u2_u15_u2_n149, u2_u15_u2_n150, u2_u15_u2_n151, 
       u2_u15_u2_n152, u2_u15_u2_n153, u2_u15_u2_n154, u2_u15_u2_n155, u2_u15_u2_n156, u2_u15_u2_n157, u2_u15_u2_n158, u2_u15_u2_n159, u2_u15_u2_n160, 
       u2_u15_u2_n161, u2_u15_u2_n162, u2_u15_u2_n163, u2_u15_u2_n164, u2_u15_u2_n165, u2_u15_u2_n166, u2_u15_u2_n167, u2_u15_u2_n168, u2_u15_u2_n169, 
       u2_u15_u2_n170, u2_u15_u2_n171, u2_u15_u2_n172, u2_u15_u2_n173, u2_u15_u2_n174, u2_u15_u2_n175, u2_u15_u2_n176, u2_u15_u2_n177, u2_u15_u2_n178, 
       u2_u15_u2_n179, u2_u15_u2_n180, u2_u15_u2_n181, u2_u15_u2_n182, u2_u15_u2_n183, u2_u15_u2_n184, u2_u15_u2_n185, u2_u15_u2_n186, u2_u15_u2_n187, 
       u2_u15_u2_n188, u2_u15_u2_n95, u2_u15_u2_n96, u2_u15_u2_n97, u2_u15_u2_n98, u2_u15_u2_n99, u2_u15_u3_n100, u2_u15_u3_n101, u2_u15_u3_n102, 
       u2_u15_u3_n103, u2_u15_u3_n104, u2_u15_u3_n105, u2_u15_u3_n106, u2_u15_u3_n107, u2_u15_u3_n108, u2_u15_u3_n109, u2_u15_u3_n110, u2_u15_u3_n111, 
       u2_u15_u3_n112, u2_u15_u3_n113, u2_u15_u3_n114, u2_u15_u3_n115, u2_u15_u3_n116, u2_u15_u3_n117, u2_u15_u3_n118, u2_u15_u3_n119, u2_u15_u3_n120, 
       u2_u15_u3_n121, u2_u15_u3_n122, u2_u15_u3_n123, u2_u15_u3_n124, u2_u15_u3_n125, u2_u15_u3_n126, u2_u15_u3_n127, u2_u15_u3_n128, u2_u15_u3_n129, 
       u2_u15_u3_n130, u2_u15_u3_n131, u2_u15_u3_n132, u2_u15_u3_n133, u2_u15_u3_n134, u2_u15_u3_n135, u2_u15_u3_n136, u2_u15_u3_n137, u2_u15_u3_n138, 
       u2_u15_u3_n139, u2_u15_u3_n140, u2_u15_u3_n141, u2_u15_u3_n142, u2_u15_u3_n143, u2_u15_u3_n144, u2_u15_u3_n145, u2_u15_u3_n146, u2_u15_u3_n147, 
       u2_u15_u3_n148, u2_u15_u3_n149, u2_u15_u3_n150, u2_u15_u3_n151, u2_u15_u3_n152, u2_u15_u3_n153, u2_u15_u3_n154, u2_u15_u3_n155, u2_u15_u3_n156, 
       u2_u15_u3_n157, u2_u15_u3_n158, u2_u15_u3_n159, u2_u15_u3_n160, u2_u15_u3_n161, u2_u15_u3_n162, u2_u15_u3_n163, u2_u15_u3_n164, u2_u15_u3_n165, 
       u2_u15_u3_n166, u2_u15_u3_n167, u2_u15_u3_n168, u2_u15_u3_n169, u2_u15_u3_n170, u2_u15_u3_n171, u2_u15_u3_n172, u2_u15_u3_n173, u2_u15_u3_n174, 
       u2_u15_u3_n175, u2_u15_u3_n176, u2_u15_u3_n177, u2_u15_u3_n178, u2_u15_u3_n179, u2_u15_u3_n180, u2_u15_u3_n181, u2_u15_u3_n182, u2_u15_u3_n183, 
       u2_u15_u3_n184, u2_u15_u3_n185, u2_u15_u3_n186, u2_u15_u3_n94, u2_u15_u3_n95, u2_u15_u3_n96, u2_u15_u3_n97, u2_u15_u3_n98, u2_u15_u3_n99, 
       u2_u1_X_10, u2_u1_X_11, u2_u1_X_12, u2_u1_X_13, u2_u1_X_14, u2_u1_X_15, u2_u1_X_16, u2_u1_X_17, u2_u1_X_18, 
       u2_u1_X_19, u2_u1_X_20, u2_u1_X_21, u2_u1_X_22, u2_u1_X_23, u2_u1_X_24, u2_u1_X_7, u2_u1_X_8, u2_u1_X_9, 
       u2_u1_u1_n100, u2_u1_u1_n101, u2_u1_u1_n102, u2_u1_u1_n103, u2_u1_u1_n104, u2_u1_u1_n105, u2_u1_u1_n106, u2_u1_u1_n107, u2_u1_u1_n108, 
       u2_u1_u1_n109, u2_u1_u1_n110, u2_u1_u1_n111, u2_u1_u1_n112, u2_u1_u1_n113, u2_u1_u1_n114, u2_u1_u1_n115, u2_u1_u1_n116, u2_u1_u1_n117, 
       u2_u1_u1_n118, u2_u1_u1_n119, u2_u1_u1_n120, u2_u1_u1_n121, u2_u1_u1_n122, u2_u1_u1_n123, u2_u1_u1_n124, u2_u1_u1_n125, u2_u1_u1_n126, 
       u2_u1_u1_n127, u2_u1_u1_n128, u2_u1_u1_n129, u2_u1_u1_n130, u2_u1_u1_n131, u2_u1_u1_n132, u2_u1_u1_n133, u2_u1_u1_n134, u2_u1_u1_n135, 
       u2_u1_u1_n136, u2_u1_u1_n137, u2_u1_u1_n138, u2_u1_u1_n139, u2_u1_u1_n140, u2_u1_u1_n141, u2_u1_u1_n142, u2_u1_u1_n143, u2_u1_u1_n144, 
       u2_u1_u1_n145, u2_u1_u1_n146, u2_u1_u1_n147, u2_u1_u1_n148, u2_u1_u1_n149, u2_u1_u1_n150, u2_u1_u1_n151, u2_u1_u1_n152, u2_u1_u1_n153, 
       u2_u1_u1_n154, u2_u1_u1_n155, u2_u1_u1_n156, u2_u1_u1_n157, u2_u1_u1_n158, u2_u1_u1_n159, u2_u1_u1_n160, u2_u1_u1_n161, u2_u1_u1_n162, 
       u2_u1_u1_n163, u2_u1_u1_n164, u2_u1_u1_n165, u2_u1_u1_n166, u2_u1_u1_n167, u2_u1_u1_n168, u2_u1_u1_n169, u2_u1_u1_n170, u2_u1_u1_n171, 
       u2_u1_u1_n172, u2_u1_u1_n173, u2_u1_u1_n174, u2_u1_u1_n175, u2_u1_u1_n176, u2_u1_u1_n177, u2_u1_u1_n178, u2_u1_u1_n179, u2_u1_u1_n180, 
       u2_u1_u1_n181, u2_u1_u1_n182, u2_u1_u1_n183, u2_u1_u1_n184, u2_u1_u1_n185, u2_u1_u1_n186, u2_u1_u1_n187, u2_u1_u1_n188, u2_u1_u1_n95, 
       u2_u1_u1_n96, u2_u1_u1_n97, u2_u1_u1_n98, u2_u1_u1_n99, u2_u1_u2_n100, u2_u1_u2_n101, u2_u1_u2_n102, u2_u1_u2_n103, u2_u1_u2_n104, 
       u2_u1_u2_n105, u2_u1_u2_n106, u2_u1_u2_n107, u2_u1_u2_n108, u2_u1_u2_n109, u2_u1_u2_n110, u2_u1_u2_n111, u2_u1_u2_n112, u2_u1_u2_n113, 
       u2_u1_u2_n114, u2_u1_u2_n115, u2_u1_u2_n116, u2_u1_u2_n117, u2_u1_u2_n118, u2_u1_u2_n119, u2_u1_u2_n120, u2_u1_u2_n121, u2_u1_u2_n122, 
       u2_u1_u2_n123, u2_u1_u2_n124, u2_u1_u2_n125, u2_u1_u2_n126, u2_u1_u2_n127, u2_u1_u2_n128, u2_u1_u2_n129, u2_u1_u2_n130, u2_u1_u2_n131, 
       u2_u1_u2_n132, u2_u1_u2_n133, u2_u1_u2_n134, u2_u1_u2_n135, u2_u1_u2_n136, u2_u1_u2_n137, u2_u1_u2_n138, u2_u1_u2_n139, u2_u1_u2_n140, 
       u2_u1_u2_n141, u2_u1_u2_n142, u2_u1_u2_n143, u2_u1_u2_n144, u2_u1_u2_n145, u2_u1_u2_n146, u2_u1_u2_n147, u2_u1_u2_n148, u2_u1_u2_n149, 
       u2_u1_u2_n150, u2_u1_u2_n151, u2_u1_u2_n152, u2_u1_u2_n153, u2_u1_u2_n154, u2_u1_u2_n155, u2_u1_u2_n156, u2_u1_u2_n157, u2_u1_u2_n158, 
       u2_u1_u2_n159, u2_u1_u2_n160, u2_u1_u2_n161, u2_u1_u2_n162, u2_u1_u2_n163, u2_u1_u2_n164, u2_u1_u2_n165, u2_u1_u2_n166, u2_u1_u2_n167, 
       u2_u1_u2_n168, u2_u1_u2_n169, u2_u1_u2_n170, u2_u1_u2_n171, u2_u1_u2_n172, u2_u1_u2_n173, u2_u1_u2_n174, u2_u1_u2_n175, u2_u1_u2_n176, 
       u2_u1_u2_n177, u2_u1_u2_n178, u2_u1_u2_n179, u2_u1_u2_n180, u2_u1_u2_n181, u2_u1_u2_n182, u2_u1_u2_n183, u2_u1_u2_n184, u2_u1_u2_n185, 
       u2_u1_u2_n186, u2_u1_u2_n187, u2_u1_u2_n188, u2_u1_u2_n95, u2_u1_u2_n96, u2_u1_u2_n97, u2_u1_u2_n98, u2_u1_u2_n99, u2_u1_u3_n100, 
       u2_u1_u3_n101, u2_u1_u3_n102, u2_u1_u3_n103, u2_u1_u3_n104, u2_u1_u3_n105, u2_u1_u3_n106, u2_u1_u3_n107, u2_u1_u3_n108, u2_u1_u3_n109, 
       u2_u1_u3_n110, u2_u1_u3_n111, u2_u1_u3_n112, u2_u1_u3_n113, u2_u1_u3_n114, u2_u1_u3_n115, u2_u1_u3_n116, u2_u1_u3_n117, u2_u1_u3_n118, 
       u2_u1_u3_n119, u2_u1_u3_n120, u2_u1_u3_n121, u2_u1_u3_n122, u2_u1_u3_n123, u2_u1_u3_n124, u2_u1_u3_n125, u2_u1_u3_n126, u2_u1_u3_n127, 
       u2_u1_u3_n128, u2_u1_u3_n129, u2_u1_u3_n130, u2_u1_u3_n131, u2_u1_u3_n132, u2_u1_u3_n133, u2_u1_u3_n134, u2_u1_u3_n135, u2_u1_u3_n136, 
       u2_u1_u3_n137, u2_u1_u3_n138, u2_u1_u3_n139, u2_u1_u3_n140, u2_u1_u3_n141, u2_u1_u3_n142, u2_u1_u3_n143, u2_u1_u3_n144, u2_u1_u3_n145, 
       u2_u1_u3_n146, u2_u1_u3_n147, u2_u1_u3_n148, u2_u1_u3_n149, u2_u1_u3_n150, u2_u1_u3_n151, u2_u1_u3_n152, u2_u1_u3_n153, u2_u1_u3_n154, 
       u2_u1_u3_n155, u2_u1_u3_n156, u2_u1_u3_n157, u2_u1_u3_n158, u2_u1_u3_n159, u2_u1_u3_n160, u2_u1_u3_n161, u2_u1_u3_n162, u2_u1_u3_n163, 
       u2_u1_u3_n164, u2_u1_u3_n165, u2_u1_u3_n166, u2_u1_u3_n167, u2_u1_u3_n168, u2_u1_u3_n169, u2_u1_u3_n170, u2_u1_u3_n171, u2_u1_u3_n172, 
       u2_u1_u3_n173, u2_u1_u3_n174, u2_u1_u3_n175, u2_u1_u3_n176, u2_u1_u3_n177, u2_u1_u3_n178, u2_u1_u3_n179, u2_u1_u3_n180, u2_u1_u3_n181, 
       u2_u1_u3_n182, u2_u1_u3_n183, u2_u1_u3_n184, u2_u1_u3_n185, u2_u1_u3_n186, u2_u1_u3_n94, u2_u1_u3_n95, u2_u1_u3_n96, u2_u1_u3_n97, 
       u2_u1_u3_n98, u2_u1_u3_n99, u2_u2_X_25, u2_u2_X_26, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_u4_n100, 
       u2_u2_u4_n101, u2_u2_u4_n102, u2_u2_u4_n103, u2_u2_u4_n104, u2_u2_u4_n105, u2_u2_u4_n106, u2_u2_u4_n107, u2_u2_u4_n108, u2_u2_u4_n109, 
       u2_u2_u4_n110, u2_u2_u4_n111, u2_u2_u4_n112, u2_u2_u4_n113, u2_u2_u4_n114, u2_u2_u4_n115, u2_u2_u4_n116, u2_u2_u4_n117, u2_u2_u4_n118, 
       u2_u2_u4_n119, u2_u2_u4_n120, u2_u2_u4_n121, u2_u2_u4_n122, u2_u2_u4_n123, u2_u2_u4_n124, u2_u2_u4_n125, u2_u2_u4_n126, u2_u2_u4_n127, 
       u2_u2_u4_n128, u2_u2_u4_n129, u2_u2_u4_n130, u2_u2_u4_n131, u2_u2_u4_n132, u2_u2_u4_n133, u2_u2_u4_n134, u2_u2_u4_n135, u2_u2_u4_n136, 
       u2_u2_u4_n137, u2_u2_u4_n138, u2_u2_u4_n139, u2_u2_u4_n140, u2_u2_u4_n141, u2_u2_u4_n142, u2_u2_u4_n143, u2_u2_u4_n144, u2_u2_u4_n145, 
       u2_u2_u4_n146, u2_u2_u4_n147, u2_u2_u4_n148, u2_u2_u4_n149, u2_u2_u4_n150, u2_u2_u4_n151, u2_u2_u4_n152, u2_u2_u4_n153, u2_u2_u4_n154, 
       u2_u2_u4_n155, u2_u2_u4_n156, u2_u2_u4_n157, u2_u2_u4_n158, u2_u2_u4_n159, u2_u2_u4_n160, u2_u2_u4_n161, u2_u2_u4_n162, u2_u2_u4_n163, 
       u2_u2_u4_n164, u2_u2_u4_n165, u2_u2_u4_n166, u2_u2_u4_n167, u2_u2_u4_n168, u2_u2_u4_n169, u2_u2_u4_n170, u2_u2_u4_n171, u2_u2_u4_n172, 
       u2_u2_u4_n173, u2_u2_u4_n174, u2_u2_u4_n175, u2_u2_u4_n176, u2_u2_u4_n177, u2_u2_u4_n178, u2_u2_u4_n179, u2_u2_u4_n180, u2_u2_u4_n181, 
       u2_u2_u4_n182, u2_u2_u4_n183, u2_u2_u4_n184, u2_u2_u4_n185, u2_u2_u4_n186, u2_u2_u4_n94, u2_u2_u4_n95, u2_u2_u4_n96, u2_u2_u4_n97, 
       u2_u2_u4_n98, u2_u2_u4_n99, u2_u3_X_1, u2_u3_X_10, u2_u3_X_11, u2_u3_X_12, u2_u3_X_2, u2_u3_X_3, u2_u3_X_37, 
       u2_u3_X_38, u2_u3_X_39, u2_u3_X_4, u2_u3_X_40, u2_u3_X_41, u2_u3_X_42, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, 
       u2_u3_X_46, u2_u3_X_47, u2_u3_X_48, u2_u3_X_5, u2_u3_X_6, u2_u3_X_7, u2_u3_X_8, u2_u3_X_9, u2_u3_u0_n100, 
       u2_u3_u0_n101, u2_u3_u0_n102, u2_u3_u0_n103, u2_u3_u0_n104, u2_u3_u0_n105, u2_u3_u0_n106, u2_u3_u0_n107, u2_u3_u0_n108, u2_u3_u0_n109, 
       u2_u3_u0_n110, u2_u3_u0_n111, u2_u3_u0_n112, u2_u3_u0_n113, u2_u3_u0_n114, u2_u3_u0_n115, u2_u3_u0_n116, u2_u3_u0_n117, u2_u3_u0_n118, 
       u2_u3_u0_n119, u2_u3_u0_n120, u2_u3_u0_n121, u2_u3_u0_n122, u2_u3_u0_n123, u2_u3_u0_n124, u2_u3_u0_n125, u2_u3_u0_n126, u2_u3_u0_n127, 
       u2_u3_u0_n128, u2_u3_u0_n129, u2_u3_u0_n130, u2_u3_u0_n131, u2_u3_u0_n132, u2_u3_u0_n133, u2_u3_u0_n134, u2_u3_u0_n135, u2_u3_u0_n136, 
       u2_u3_u0_n137, u2_u3_u0_n138, u2_u3_u0_n139, u2_u3_u0_n140, u2_u3_u0_n141, u2_u3_u0_n142, u2_u3_u0_n143, u2_u3_u0_n144, u2_u3_u0_n145, 
       u2_u3_u0_n146, u2_u3_u0_n147, u2_u3_u0_n148, u2_u3_u0_n149, u2_u3_u0_n150, u2_u3_u0_n151, u2_u3_u0_n152, u2_u3_u0_n153, u2_u3_u0_n154, 
       u2_u3_u0_n155, u2_u3_u0_n156, u2_u3_u0_n157, u2_u3_u0_n158, u2_u3_u0_n159, u2_u3_u0_n160, u2_u3_u0_n161, u2_u3_u0_n162, u2_u3_u0_n163, 
       u2_u3_u0_n164, u2_u3_u0_n165, u2_u3_u0_n166, u2_u3_u0_n167, u2_u3_u0_n168, u2_u3_u0_n169, u2_u3_u0_n170, u2_u3_u0_n171, u2_u3_u0_n172, 
       u2_u3_u0_n173, u2_u3_u0_n174, u2_u3_u0_n88, u2_u3_u0_n89, u2_u3_u0_n90, u2_u3_u0_n91, u2_u3_u0_n92, u2_u3_u0_n93, u2_u3_u0_n94, 
       u2_u3_u0_n95, u2_u3_u0_n96, u2_u3_u0_n97, u2_u3_u0_n98, u2_u3_u0_n99, u2_u3_u1_n100, u2_u3_u1_n101, u2_u3_u1_n102, u2_u3_u1_n103, 
       u2_u3_u1_n104, u2_u3_u1_n105, u2_u3_u1_n106, u2_u3_u1_n107, u2_u3_u1_n108, u2_u3_u1_n109, u2_u3_u1_n110, u2_u3_u1_n111, u2_u3_u1_n112, 
       u2_u3_u1_n113, u2_u3_u1_n114, u2_u3_u1_n115, u2_u3_u1_n116, u2_u3_u1_n117, u2_u3_u1_n118, u2_u3_u1_n119, u2_u3_u1_n120, u2_u3_u1_n121, 
       u2_u3_u1_n122, u2_u3_u1_n123, u2_u3_u1_n124, u2_u3_u1_n125, u2_u3_u1_n126, u2_u3_u1_n127, u2_u3_u1_n128, u2_u3_u1_n129, u2_u3_u1_n130, 
       u2_u3_u1_n131, u2_u3_u1_n132, u2_u3_u1_n133, u2_u3_u1_n134, u2_u3_u1_n135, u2_u3_u1_n136, u2_u3_u1_n137, u2_u3_u1_n138, u2_u3_u1_n139, 
       u2_u3_u1_n140, u2_u3_u1_n141, u2_u3_u1_n142, u2_u3_u1_n143, u2_u3_u1_n144, u2_u3_u1_n145, u2_u3_u1_n146, u2_u3_u1_n147, u2_u3_u1_n148, 
       u2_u3_u1_n149, u2_u3_u1_n150, u2_u3_u1_n151, u2_u3_u1_n152, u2_u3_u1_n153, u2_u3_u1_n154, u2_u3_u1_n155, u2_u3_u1_n156, u2_u3_u1_n157, 
       u2_u3_u1_n158, u2_u3_u1_n159, u2_u3_u1_n160, u2_u3_u1_n161, u2_u3_u1_n162, u2_u3_u1_n163, u2_u3_u1_n164, u2_u3_u1_n165, u2_u3_u1_n166, 
       u2_u3_u1_n167, u2_u3_u1_n168, u2_u3_u1_n169, u2_u3_u1_n170, u2_u3_u1_n171, u2_u3_u1_n172, u2_u3_u1_n173, u2_u3_u1_n174, u2_u3_u1_n175, 
       u2_u3_u1_n176, u2_u3_u1_n177, u2_u3_u1_n178, u2_u3_u1_n179, u2_u3_u1_n180, u2_u3_u1_n181, u2_u3_u1_n182, u2_u3_u1_n183, u2_u3_u1_n184, 
       u2_u3_u1_n185, u2_u3_u1_n186, u2_u3_u1_n187, u2_u3_u1_n188, u2_u3_u1_n95, u2_u3_u1_n96, u2_u3_u1_n97, u2_u3_u1_n98, u2_u3_u1_n99, 
       u2_u3_u6_n100, u2_u3_u6_n101, u2_u3_u6_n102, u2_u3_u6_n103, u2_u3_u6_n104, u2_u3_u6_n105, u2_u3_u6_n106, u2_u3_u6_n107, u2_u3_u6_n108, 
       u2_u3_u6_n109, u2_u3_u6_n110, u2_u3_u6_n111, u2_u3_u6_n112, u2_u3_u6_n113, u2_u3_u6_n114, u2_u3_u6_n115, u2_u3_u6_n116, u2_u3_u6_n117, 
       u2_u3_u6_n118, u2_u3_u6_n119, u2_u3_u6_n120, u2_u3_u6_n121, u2_u3_u6_n122, u2_u3_u6_n123, u2_u3_u6_n124, u2_u3_u6_n125, u2_u3_u6_n126, 
       u2_u3_u6_n127, u2_u3_u6_n128, u2_u3_u6_n129, u2_u3_u6_n130, u2_u3_u6_n131, u2_u3_u6_n132, u2_u3_u6_n133, u2_u3_u6_n134, u2_u3_u6_n135, 
       u2_u3_u6_n136, u2_u3_u6_n137, u2_u3_u6_n138, u2_u3_u6_n139, u2_u3_u6_n140, u2_u3_u6_n141, u2_u3_u6_n142, u2_u3_u6_n143, u2_u3_u6_n144, 
       u2_u3_u6_n145, u2_u3_u6_n146, u2_u3_u6_n147, u2_u3_u6_n148, u2_u3_u6_n149, u2_u3_u6_n150, u2_u3_u6_n151, u2_u3_u6_n152, u2_u3_u6_n153, 
       u2_u3_u6_n154, u2_u3_u6_n155, u2_u3_u6_n156, u2_u3_u6_n157, u2_u3_u6_n158, u2_u3_u6_n159, u2_u3_u6_n160, u2_u3_u6_n161, u2_u3_u6_n162, 
       u2_u3_u6_n163, u2_u3_u6_n164, u2_u3_u6_n165, u2_u3_u6_n166, u2_u3_u6_n167, u2_u3_u6_n168, u2_u3_u6_n169, u2_u3_u6_n170, u2_u3_u6_n171, 
       u2_u3_u6_n172, u2_u3_u6_n173, u2_u3_u6_n174, u2_u3_u6_n88, u2_u3_u6_n89, u2_u3_u6_n90, u2_u3_u6_n91, u2_u3_u6_n92, u2_u3_u6_n93, 
       u2_u3_u6_n94, u2_u3_u6_n95, u2_u3_u6_n96, u2_u3_u6_n97, u2_u3_u6_n98, u2_u3_u6_n99, u2_u3_u7_n100, u2_u3_u7_n101, u2_u3_u7_n102, 
       u2_u3_u7_n103, u2_u3_u7_n104, u2_u3_u7_n105, u2_u3_u7_n106, u2_u3_u7_n107, u2_u3_u7_n108, u2_u3_u7_n109, u2_u3_u7_n110, u2_u3_u7_n111, 
       u2_u3_u7_n112, u2_u3_u7_n113, u2_u3_u7_n114, u2_u3_u7_n115, u2_u3_u7_n116, u2_u3_u7_n117, u2_u3_u7_n118, u2_u3_u7_n119, u2_u3_u7_n120, 
       u2_u3_u7_n121, u2_u3_u7_n122, u2_u3_u7_n123, u2_u3_u7_n124, u2_u3_u7_n125, u2_u3_u7_n126, u2_u3_u7_n127, u2_u3_u7_n128, u2_u3_u7_n129, 
       u2_u3_u7_n130, u2_u3_u7_n131, u2_u3_u7_n132, u2_u3_u7_n133, u2_u3_u7_n134, u2_u3_u7_n135, u2_u3_u7_n136, u2_u3_u7_n137, u2_u3_u7_n138, 
       u2_u3_u7_n139, u2_u3_u7_n140, u2_u3_u7_n141, u2_u3_u7_n142, u2_u3_u7_n143, u2_u3_u7_n144, u2_u3_u7_n145, u2_u3_u7_n146, u2_u3_u7_n147, 
       u2_u3_u7_n148, u2_u3_u7_n149, u2_u3_u7_n150, u2_u3_u7_n151, u2_u3_u7_n152, u2_u3_u7_n153, u2_u3_u7_n154, u2_u3_u7_n155, u2_u3_u7_n156, 
       u2_u3_u7_n157, u2_u3_u7_n158, u2_u3_u7_n159, u2_u3_u7_n160, u2_u3_u7_n161, u2_u3_u7_n162, u2_u3_u7_n163, u2_u3_u7_n164, u2_u3_u7_n165, 
       u2_u3_u7_n166, u2_u3_u7_n167, u2_u3_u7_n168, u2_u3_u7_n169, u2_u3_u7_n170, u2_u3_u7_n171, u2_u3_u7_n172, u2_u3_u7_n173, u2_u3_u7_n174, 
       u2_u3_u7_n175, u2_u3_u7_n176, u2_u3_u7_n177, u2_u3_u7_n178, u2_u3_u7_n179, u2_u3_u7_n180, u2_u3_u7_n91, u2_u3_u7_n92, u2_u3_u7_n93, 
       u2_u3_u7_n94, u2_u3_u7_n95, u2_u3_u7_n96, u2_u3_u7_n97, u2_u3_u7_n98, u2_u3_u7_n99, u2_u4_X_25, u2_u4_X_26, u2_u4_X_27, 
       u2_u4_X_28, u2_u4_X_29, u2_u4_X_30, u2_u4_X_31, u2_u4_X_32, u2_u4_X_33, u2_u4_X_34, u2_u4_X_35, u2_u4_X_36, 
       u2_u4_X_37, u2_u4_X_38, u2_u4_X_39, u2_u4_X_40, u2_u4_X_41, u2_u4_X_42, u2_u4_u4_n100, u2_u4_u4_n101, u2_u4_u4_n102, 
       u2_u4_u4_n103, u2_u4_u4_n104, u2_u4_u4_n105, u2_u4_u4_n106, u2_u4_u4_n107, u2_u4_u4_n108, u2_u4_u4_n109, u2_u4_u4_n110, u2_u4_u4_n111, 
       u2_u4_u4_n112, u2_u4_u4_n113, u2_u4_u4_n114, u2_u4_u4_n115, u2_u4_u4_n116, u2_u4_u4_n117, u2_u4_u4_n118, u2_u4_u4_n119, u2_u4_u4_n120, 
       u2_u4_u4_n121, u2_u4_u4_n122, u2_u4_u4_n123, u2_u4_u4_n124, u2_u4_u4_n125, u2_u4_u4_n126, u2_u4_u4_n127, u2_u4_u4_n128, u2_u4_u4_n129, 
       u2_u4_u4_n130, u2_u4_u4_n131, u2_u4_u4_n132, u2_u4_u4_n133, u2_u4_u4_n134, u2_u4_u4_n135, u2_u4_u4_n136, u2_u4_u4_n137, u2_u4_u4_n138, 
       u2_u4_u4_n139, u2_u4_u4_n140, u2_u4_u4_n141, u2_u4_u4_n142, u2_u4_u4_n143, u2_u4_u4_n144, u2_u4_u4_n145, u2_u4_u4_n146, u2_u4_u4_n147, 
       u2_u4_u4_n148, u2_u4_u4_n149, u2_u4_u4_n150, u2_u4_u4_n151, u2_u4_u4_n152, u2_u4_u4_n153, u2_u4_u4_n154, u2_u4_u4_n155, u2_u4_u4_n156, 
       u2_u4_u4_n157, u2_u4_u4_n158, u2_u4_u4_n159, u2_u4_u4_n160, u2_u4_u4_n161, u2_u4_u4_n162, u2_u4_u4_n163, u2_u4_u4_n164, u2_u4_u4_n165, 
       u2_u4_u4_n166, u2_u4_u4_n167, u2_u4_u4_n168, u2_u4_u4_n169, u2_u4_u4_n170, u2_u4_u4_n171, u2_u4_u4_n172, u2_u4_u4_n173, u2_u4_u4_n174, 
       u2_u4_u4_n175, u2_u4_u4_n176, u2_u4_u4_n177, u2_u4_u4_n178, u2_u4_u4_n179, u2_u4_u4_n180, u2_u4_u4_n181, u2_u4_u4_n182, u2_u4_u4_n183, 
       u2_u4_u4_n184, u2_u4_u4_n185, u2_u4_u4_n186, u2_u4_u4_n94, u2_u4_u4_n95, u2_u4_u4_n96, u2_u4_u4_n97, u2_u4_u4_n98, u2_u4_u4_n99, 
       u2_u4_u5_n100, u2_u4_u5_n101, u2_u4_u5_n102, u2_u4_u5_n103, u2_u4_u5_n104, u2_u4_u5_n105, u2_u4_u5_n106, u2_u4_u5_n107, u2_u4_u5_n108, 
       u2_u4_u5_n109, u2_u4_u5_n110, u2_u4_u5_n111, u2_u4_u5_n112, u2_u4_u5_n113, u2_u4_u5_n114, u2_u4_u5_n115, u2_u4_u5_n116, u2_u4_u5_n117, 
       u2_u4_u5_n118, u2_u4_u5_n119, u2_u4_u5_n120, u2_u4_u5_n121, u2_u4_u5_n122, u2_u4_u5_n123, u2_u4_u5_n124, u2_u4_u5_n125, u2_u4_u5_n126, 
       u2_u4_u5_n127, u2_u4_u5_n128, u2_u4_u5_n129, u2_u4_u5_n130, u2_u4_u5_n131, u2_u4_u5_n132, u2_u4_u5_n133, u2_u4_u5_n134, u2_u4_u5_n135, 
       u2_u4_u5_n136, u2_u4_u5_n137, u2_u4_u5_n138, u2_u4_u5_n139, u2_u4_u5_n140, u2_u4_u5_n141, u2_u4_u5_n142, u2_u4_u5_n143, u2_u4_u5_n144, 
       u2_u4_u5_n145, u2_u4_u5_n146, u2_u4_u5_n147, u2_u4_u5_n148, u2_u4_u5_n149, u2_u4_u5_n150, u2_u4_u5_n151, u2_u4_u5_n152, u2_u4_u5_n153, 
       u2_u4_u5_n154, u2_u4_u5_n155, u2_u4_u5_n156, u2_u4_u5_n157, u2_u4_u5_n158, u2_u4_u5_n159, u2_u4_u5_n160, u2_u4_u5_n161, u2_u4_u5_n162, 
       u2_u4_u5_n163, u2_u4_u5_n164, u2_u4_u5_n165, u2_u4_u5_n166, u2_u4_u5_n167, u2_u4_u5_n168, u2_u4_u5_n169, u2_u4_u5_n170, u2_u4_u5_n171, 
       u2_u4_u5_n172, u2_u4_u5_n173, u2_u4_u5_n174, u2_u4_u5_n175, u2_u4_u5_n176, u2_u4_u5_n177, u2_u4_u5_n178, u2_u4_u5_n179, u2_u4_u5_n180, 
       u2_u4_u5_n181, u2_u4_u5_n182, u2_u4_u5_n183, u2_u4_u5_n184, u2_u4_u5_n185, u2_u4_u5_n186, u2_u4_u5_n187, u2_u4_u5_n188, u2_u4_u5_n189, 
       u2_u4_u5_n190, u2_u4_u5_n191, u2_u4_u5_n192, u2_u4_u5_n193, u2_u4_u5_n194, u2_u4_u5_n195, u2_u4_u5_n196, u2_u4_u5_n99, u2_u4_u6_n100, 
       u2_u4_u6_n101, u2_u4_u6_n102, u2_u4_u6_n103, u2_u4_u6_n104, u2_u4_u6_n105, u2_u4_u6_n106, u2_u4_u6_n107, u2_u4_u6_n108, u2_u4_u6_n109, 
       u2_u4_u6_n110, u2_u4_u6_n111, u2_u4_u6_n112, u2_u4_u6_n113, u2_u4_u6_n114, u2_u4_u6_n115, u2_u4_u6_n116, u2_u4_u6_n117, u2_u4_u6_n118, 
       u2_u4_u6_n119, u2_u4_u6_n120, u2_u4_u6_n121, u2_u4_u6_n122, u2_u4_u6_n123, u2_u4_u6_n124, u2_u4_u6_n125, u2_u4_u6_n126, u2_u4_u6_n127, 
       u2_u4_u6_n128, u2_u4_u6_n129, u2_u4_u6_n130, u2_u4_u6_n131, u2_u4_u6_n132, u2_u4_u6_n133, u2_u4_u6_n134, u2_u4_u6_n135, u2_u4_u6_n136, 
       u2_u4_u6_n137, u2_u4_u6_n138, u2_u4_u6_n139, u2_u4_u6_n140, u2_u4_u6_n141, u2_u4_u6_n142, u2_u4_u6_n143, u2_u4_u6_n144, u2_u4_u6_n145, 
       u2_u4_u6_n146, u2_u4_u6_n147, u2_u4_u6_n148, u2_u4_u6_n149, u2_u4_u6_n150, u2_u4_u6_n151, u2_u4_u6_n152, u2_u4_u6_n153, u2_u4_u6_n154, 
       u2_u4_u6_n155, u2_u4_u6_n156, u2_u4_u6_n157, u2_u4_u6_n158, u2_u4_u6_n159, u2_u4_u6_n160, u2_u4_u6_n161, u2_u4_u6_n162, u2_u4_u6_n163, 
       u2_u4_u6_n164, u2_u4_u6_n165, u2_u4_u6_n166, u2_u4_u6_n167, u2_u4_u6_n168, u2_u4_u6_n169, u2_u4_u6_n170, u2_u4_u6_n171, u2_u4_u6_n172, 
       u2_u4_u6_n173, u2_u4_u6_n174, u2_u4_u6_n88, u2_u4_u6_n89, u2_u4_u6_n90, u2_u4_u6_n91, u2_u4_u6_n92, u2_u4_u6_n93, u2_u4_u6_n94, 
       u2_u4_u6_n95, u2_u4_u6_n96, u2_u4_u6_n97, u2_u4_u6_n98, u2_u4_u6_n99, u2_u5_X_1, u2_u5_X_10, u2_u5_X_11, u2_u5_X_12, 
       u2_u5_X_2, u2_u5_X_3, u2_u5_X_31, u2_u5_X_32, u2_u5_X_33, u2_u5_X_34, u2_u5_X_35, u2_u5_X_36, u2_u5_X_37, 
       u2_u5_X_38, u2_u5_X_39, u2_u5_X_4, u2_u5_X_40, u2_u5_X_41, u2_u5_X_42, u2_u5_X_43, u2_u5_X_44, u2_u5_X_45, 
       u2_u5_X_46, u2_u5_X_47, u2_u5_X_48, u2_u5_X_5, u2_u5_X_6, u2_u5_X_7, u2_u5_X_8, u2_u5_X_9, u2_u5_u0_n100, 
       u2_u5_u0_n101, u2_u5_u0_n102, u2_u5_u0_n103, u2_u5_u0_n104, u2_u5_u0_n105, u2_u5_u0_n106, u2_u5_u0_n107, u2_u5_u0_n108, u2_u5_u0_n109, 
       u2_u5_u0_n110, u2_u5_u0_n111, u2_u5_u0_n112, u2_u5_u0_n113, u2_u5_u0_n114, u2_u5_u0_n115, u2_u5_u0_n116, u2_u5_u0_n117, u2_u5_u0_n118, 
       u2_u5_u0_n119, u2_u5_u0_n120, u2_u5_u0_n121, u2_u5_u0_n122, u2_u5_u0_n123, u2_u5_u0_n124, u2_u5_u0_n125, u2_u5_u0_n126, u2_u5_u0_n127, 
       u2_u5_u0_n128, u2_u5_u0_n129, u2_u5_u0_n130, u2_u5_u0_n131, u2_u5_u0_n132, u2_u5_u0_n133, u2_u5_u0_n134, u2_u5_u0_n135, u2_u5_u0_n136, 
       u2_u5_u0_n137, u2_u5_u0_n138, u2_u5_u0_n139, u2_u5_u0_n140, u2_u5_u0_n141, u2_u5_u0_n142, u2_u5_u0_n143, u2_u5_u0_n144, u2_u5_u0_n145, 
       u2_u5_u0_n146, u2_u5_u0_n147, u2_u5_u0_n148, u2_u5_u0_n149, u2_u5_u0_n150, u2_u5_u0_n151, u2_u5_u0_n152, u2_u5_u0_n153, u2_u5_u0_n154, 
       u2_u5_u0_n155, u2_u5_u0_n156, u2_u5_u0_n157, u2_u5_u0_n158, u2_u5_u0_n159, u2_u5_u0_n160, u2_u5_u0_n161, u2_u5_u0_n162, u2_u5_u0_n163, 
       u2_u5_u0_n164, u2_u5_u0_n165, u2_u5_u0_n166, u2_u5_u0_n167, u2_u5_u0_n168, u2_u5_u0_n169, u2_u5_u0_n170, u2_u5_u0_n171, u2_u5_u0_n172, 
       u2_u5_u0_n173, u2_u5_u0_n174, u2_u5_u0_n88, u2_u5_u0_n89, u2_u5_u0_n90, u2_u5_u0_n91, u2_u5_u0_n92, u2_u5_u0_n93, u2_u5_u0_n94, 
       u2_u5_u0_n95, u2_u5_u0_n96, u2_u5_u0_n97, u2_u5_u0_n98, u2_u5_u0_n99, u2_u5_u1_n100, u2_u5_u1_n101, u2_u5_u1_n102, u2_u5_u1_n103, 
       u2_u5_u1_n104, u2_u5_u1_n105, u2_u5_u1_n106, u2_u5_u1_n107, u2_u5_u1_n108, u2_u5_u1_n109, u2_u5_u1_n110, u2_u5_u1_n111, u2_u5_u1_n112, 
       u2_u5_u1_n113, u2_u5_u1_n114, u2_u5_u1_n115, u2_u5_u1_n116, u2_u5_u1_n117, u2_u5_u1_n118, u2_u5_u1_n119, u2_u5_u1_n120, u2_u5_u1_n121, 
       u2_u5_u1_n122, u2_u5_u1_n123, u2_u5_u1_n124, u2_u5_u1_n125, u2_u5_u1_n126, u2_u5_u1_n127, u2_u5_u1_n128, u2_u5_u1_n129, u2_u5_u1_n130, 
       u2_u5_u1_n131, u2_u5_u1_n132, u2_u5_u1_n133, u2_u5_u1_n134, u2_u5_u1_n135, u2_u5_u1_n136, u2_u5_u1_n137, u2_u5_u1_n138, u2_u5_u1_n139, 
       u2_u5_u1_n140, u2_u5_u1_n141, u2_u5_u1_n142, u2_u5_u1_n143, u2_u5_u1_n144, u2_u5_u1_n145, u2_u5_u1_n146, u2_u5_u1_n147, u2_u5_u1_n148, 
       u2_u5_u1_n149, u2_u5_u1_n150, u2_u5_u1_n151, u2_u5_u1_n152, u2_u5_u1_n153, u2_u5_u1_n154, u2_u5_u1_n155, u2_u5_u1_n156, u2_u5_u1_n157, 
       u2_u5_u1_n158, u2_u5_u1_n159, u2_u5_u1_n160, u2_u5_u1_n161, u2_u5_u1_n162, u2_u5_u1_n163, u2_u5_u1_n164, u2_u5_u1_n165, u2_u5_u1_n166, 
       u2_u5_u1_n167, u2_u5_u1_n168, u2_u5_u1_n169, u2_u5_u1_n170, u2_u5_u1_n171, u2_u5_u1_n172, u2_u5_u1_n173, u2_u5_u1_n174, u2_u5_u1_n175, 
       u2_u5_u1_n176, u2_u5_u1_n177, u2_u5_u1_n178, u2_u5_u1_n179, u2_u5_u1_n180, u2_u5_u1_n181, u2_u5_u1_n182, u2_u5_u1_n183, u2_u5_u1_n184, 
       u2_u5_u1_n185, u2_u5_u1_n186, u2_u5_u1_n187, u2_u5_u1_n188, u2_u5_u1_n95, u2_u5_u1_n96, u2_u5_u1_n97, u2_u5_u1_n98, u2_u5_u1_n99, 
       u2_u5_u5_n100, u2_u5_u5_n101, u2_u5_u5_n102, u2_u5_u5_n103, u2_u5_u5_n104, u2_u5_u5_n105, u2_u5_u5_n106, u2_u5_u5_n107, u2_u5_u5_n108, 
       u2_u5_u5_n109, u2_u5_u5_n110, u2_u5_u5_n111, u2_u5_u5_n112, u2_u5_u5_n113, u2_u5_u5_n114, u2_u5_u5_n115, u2_u5_u5_n116, u2_u5_u5_n117, 
       u2_u5_u5_n118, u2_u5_u5_n119, u2_u5_u5_n120, u2_u5_u5_n121, u2_u5_u5_n122, u2_u5_u5_n123, u2_u5_u5_n124, u2_u5_u5_n125, u2_u5_u5_n126, 
       u2_u5_u5_n127, u2_u5_u5_n128, u2_u5_u5_n129, u2_u5_u5_n130, u2_u5_u5_n131, u2_u5_u5_n132, u2_u5_u5_n133, u2_u5_u5_n134, u2_u5_u5_n135, 
       u2_u5_u5_n136, u2_u5_u5_n137, u2_u5_u5_n138, u2_u5_u5_n139, u2_u5_u5_n140, u2_u5_u5_n141, u2_u5_u5_n142, u2_u5_u5_n143, u2_u5_u5_n144, 
       u2_u5_u5_n145, u2_u5_u5_n146, u2_u5_u5_n147, u2_u5_u5_n148, u2_u5_u5_n149, u2_u5_u5_n150, u2_u5_u5_n151, u2_u5_u5_n152, u2_u5_u5_n153, 
       u2_u5_u5_n154, u2_u5_u5_n155, u2_u5_u5_n156, u2_u5_u5_n157, u2_u5_u5_n158, u2_u5_u5_n159, u2_u5_u5_n160, u2_u5_u5_n161, u2_u5_u5_n162, 
       u2_u5_u5_n163, u2_u5_u5_n164, u2_u5_u5_n165, u2_u5_u5_n166, u2_u5_u5_n167, u2_u5_u5_n168, u2_u5_u5_n169, u2_u5_u5_n170, u2_u5_u5_n171, 
       u2_u5_u5_n172, u2_u5_u5_n173, u2_u5_u5_n174, u2_u5_u5_n175, u2_u5_u5_n176, u2_u5_u5_n177, u2_u5_u5_n178, u2_u5_u5_n179, u2_u5_u5_n180, 
       u2_u5_u5_n181, u2_u5_u5_n182, u2_u5_u5_n183, u2_u5_u5_n184, u2_u5_u5_n185, u2_u5_u5_n186, u2_u5_u5_n187, u2_u5_u5_n188, u2_u5_u5_n189, 
       u2_u5_u5_n190, u2_u5_u5_n191, u2_u5_u5_n192, u2_u5_u5_n193, u2_u5_u5_n194, u2_u5_u5_n195, u2_u5_u5_n196, u2_u5_u5_n99, u2_u5_u6_n100, 
       u2_u5_u6_n101, u2_u5_u6_n102, u2_u5_u6_n103, u2_u5_u6_n104, u2_u5_u6_n105, u2_u5_u6_n106, u2_u5_u6_n107, u2_u5_u6_n108, u2_u5_u6_n109, 
       u2_u5_u6_n110, u2_u5_u6_n111, u2_u5_u6_n112, u2_u5_u6_n113, u2_u5_u6_n114, u2_u5_u6_n115, u2_u5_u6_n116, u2_u5_u6_n117, u2_u5_u6_n118, 
       u2_u5_u6_n119, u2_u5_u6_n120, u2_u5_u6_n121, u2_u5_u6_n122, u2_u5_u6_n123, u2_u5_u6_n124, u2_u5_u6_n125, u2_u5_u6_n126, u2_u5_u6_n127, 
       u2_u5_u6_n128, u2_u5_u6_n129, u2_u5_u6_n130, u2_u5_u6_n131, u2_u5_u6_n132, u2_u5_u6_n133, u2_u5_u6_n134, u2_u5_u6_n135, u2_u5_u6_n136, 
       u2_u5_u6_n137, u2_u5_u6_n138, u2_u5_u6_n139, u2_u5_u6_n140, u2_u5_u6_n141, u2_u5_u6_n142, u2_u5_u6_n143, u2_u5_u6_n144, u2_u5_u6_n145, 
       u2_u5_u6_n146, u2_u5_u6_n147, u2_u5_u6_n148, u2_u5_u6_n149, u2_u5_u6_n150, u2_u5_u6_n151, u2_u5_u6_n152, u2_u5_u6_n153, u2_u5_u6_n154, 
       u2_u5_u6_n155, u2_u5_u6_n156, u2_u5_u6_n157, u2_u5_u6_n158, u2_u5_u6_n159, u2_u5_u6_n160, u2_u5_u6_n161, u2_u5_u6_n162, u2_u5_u6_n163, 
       u2_u5_u6_n164, u2_u5_u6_n165, u2_u5_u6_n166, u2_u5_u6_n167, u2_u5_u6_n168, u2_u5_u6_n169, u2_u5_u6_n170, u2_u5_u6_n171, u2_u5_u6_n172, 
       u2_u5_u6_n173, u2_u5_u6_n174, u2_u5_u6_n88, u2_u5_u6_n89, u2_u5_u6_n90, u2_u5_u6_n91, u2_u5_u6_n92, u2_u5_u6_n93, u2_u5_u6_n94, 
       u2_u5_u6_n95, u2_u5_u6_n96, u2_u5_u6_n97, u2_u5_u6_n98, u2_u5_u6_n99, u2_u5_u7_n100, u2_u5_u7_n101, u2_u5_u7_n102, u2_u5_u7_n103, 
       u2_u5_u7_n104, u2_u5_u7_n105, u2_u5_u7_n106, u2_u5_u7_n107, u2_u5_u7_n108, u2_u5_u7_n109, u2_u5_u7_n110, u2_u5_u7_n111, u2_u5_u7_n112, 
       u2_u5_u7_n113, u2_u5_u7_n114, u2_u5_u7_n115, u2_u5_u7_n116, u2_u5_u7_n117, u2_u5_u7_n118, u2_u5_u7_n119, u2_u5_u7_n120, u2_u5_u7_n121, 
       u2_u5_u7_n122, u2_u5_u7_n123, u2_u5_u7_n124, u2_u5_u7_n125, u2_u5_u7_n126, u2_u5_u7_n127, u2_u5_u7_n128, u2_u5_u7_n129, u2_u5_u7_n130, 
       u2_u5_u7_n131, u2_u5_u7_n132, u2_u5_u7_n133, u2_u5_u7_n134, u2_u5_u7_n135, u2_u5_u7_n136, u2_u5_u7_n137, u2_u5_u7_n138, u2_u5_u7_n139, 
       u2_u5_u7_n140, u2_u5_u7_n141, u2_u5_u7_n142, u2_u5_u7_n143, u2_u5_u7_n144, u2_u5_u7_n145, u2_u5_u7_n146, u2_u5_u7_n147, u2_u5_u7_n148, 
       u2_u5_u7_n149, u2_u5_u7_n150, u2_u5_u7_n151, u2_u5_u7_n152, u2_u5_u7_n153, u2_u5_u7_n154, u2_u5_u7_n155, u2_u5_u7_n156, u2_u5_u7_n157, 
       u2_u5_u7_n158, u2_u5_u7_n159, u2_u5_u7_n160, u2_u5_u7_n161, u2_u5_u7_n162, u2_u5_u7_n163, u2_u5_u7_n164, u2_u5_u7_n165, u2_u5_u7_n166, 
       u2_u5_u7_n167, u2_u5_u7_n168, u2_u5_u7_n169, u2_u5_u7_n170, u2_u5_u7_n171, u2_u5_u7_n172, u2_u5_u7_n173, u2_u5_u7_n174, u2_u5_u7_n175, 
       u2_u5_u7_n176, u2_u5_u7_n177, u2_u5_u7_n178, u2_u5_u7_n179, u2_u5_u7_n180, u2_u5_u7_n91, u2_u5_u7_n92, u2_u5_u7_n93, u2_u5_u7_n94, 
       u2_u5_u7_n95, u2_u5_u7_n96, u2_u5_u7_n97, u2_u5_u7_n98, u2_u5_u7_n99, u2_u6_X_31, u2_u6_X_32, u2_u6_X_33, u2_u6_X_34, 
       u2_u6_X_35, u2_u6_X_36, u2_u6_u5_n100, u2_u6_u5_n101, u2_u6_u5_n102, u2_u6_u5_n103, u2_u6_u5_n104, u2_u6_u5_n105, u2_u6_u5_n106, 
       u2_u6_u5_n107, u2_u6_u5_n108, u2_u6_u5_n109, u2_u6_u5_n110, u2_u6_u5_n111, u2_u6_u5_n112, u2_u6_u5_n113, u2_u6_u5_n114, u2_u6_u5_n115, 
       u2_u6_u5_n116, u2_u6_u5_n117, u2_u6_u5_n118, u2_u6_u5_n119, u2_u6_u5_n120, u2_u6_u5_n121, u2_u6_u5_n122, u2_u6_u5_n123, u2_u6_u5_n124, 
       u2_u6_u5_n125, u2_u6_u5_n126, u2_u6_u5_n127, u2_u6_u5_n128, u2_u6_u5_n129, u2_u6_u5_n130, u2_u6_u5_n131, u2_u6_u5_n132, u2_u6_u5_n133, 
       u2_u6_u5_n134, u2_u6_u5_n135, u2_u6_u5_n136, u2_u6_u5_n137, u2_u6_u5_n138, u2_u6_u5_n139, u2_u6_u5_n140, u2_u6_u5_n141, u2_u6_u5_n142, 
       u2_u6_u5_n143, u2_u6_u5_n144, u2_u6_u5_n145, u2_u6_u5_n146, u2_u6_u5_n147, u2_u6_u5_n148, u2_u6_u5_n149, u2_u6_u5_n150, u2_u6_u5_n151, 
       u2_u6_u5_n152, u2_u6_u5_n153, u2_u6_u5_n154, u2_u6_u5_n155, u2_u6_u5_n156, u2_u6_u5_n157, u2_u6_u5_n158, u2_u6_u5_n159, u2_u6_u5_n160, 
       u2_u6_u5_n161, u2_u6_u5_n162, u2_u6_u5_n163, u2_u6_u5_n164, u2_u6_u5_n165, u2_u6_u5_n166, u2_u6_u5_n167, u2_u6_u5_n168, u2_u6_u5_n169, 
       u2_u6_u5_n170, u2_u6_u5_n171, u2_u6_u5_n172, u2_u6_u5_n173, u2_u6_u5_n174, u2_u6_u5_n175, u2_u6_u5_n176, u2_u6_u5_n177, u2_u6_u5_n178, 
       u2_u6_u5_n179, u2_u6_u5_n180, u2_u6_u5_n181, u2_u6_u5_n182, u2_u6_u5_n183, u2_u6_u5_n184, u2_u6_u5_n185, u2_u6_u5_n186, u2_u6_u5_n187, 
       u2_u6_u5_n188, u2_u6_u5_n189, u2_u6_u5_n190, u2_u6_u5_n191, u2_u6_u5_n192, u2_u6_u5_n193, u2_u6_u5_n194, u2_u6_u5_n195, u2_u6_u5_n196, 
       u2_u6_u5_n99, u2_u7_X_25, u2_u7_X_26, u2_u7_X_27, u2_u7_X_28, u2_u7_X_29, u2_u7_X_30, u2_u7_X_31, u2_u7_X_32, 
       u2_u7_X_33, u2_u7_X_34, u2_u7_X_35, u2_u7_X_36, u2_u7_u4_n100, u2_u7_u4_n101, u2_u7_u4_n102, u2_u7_u4_n103, u2_u7_u4_n104, 
       u2_u7_u4_n105, u2_u7_u4_n106, u2_u7_u4_n107, u2_u7_u4_n108, u2_u7_u4_n109, u2_u7_u4_n110, u2_u7_u4_n111, u2_u7_u4_n112, u2_u7_u4_n113, 
       u2_u7_u4_n114, u2_u7_u4_n115, u2_u7_u4_n116, u2_u7_u4_n117, u2_u7_u4_n118, u2_u7_u4_n119, u2_u7_u4_n120, u2_u7_u4_n121, u2_u7_u4_n122, 
       u2_u7_u4_n123, u2_u7_u4_n124, u2_u7_u4_n125, u2_u7_u4_n126, u2_u7_u4_n127, u2_u7_u4_n128, u2_u7_u4_n129, u2_u7_u4_n130, u2_u7_u4_n131, 
       u2_u7_u4_n132, u2_u7_u4_n133, u2_u7_u4_n134, u2_u7_u4_n135, u2_u7_u4_n136, u2_u7_u4_n137, u2_u7_u4_n138, u2_u7_u4_n139, u2_u7_u4_n140, 
       u2_u7_u4_n141, u2_u7_u4_n142, u2_u7_u4_n143, u2_u7_u4_n144, u2_u7_u4_n145, u2_u7_u4_n146, u2_u7_u4_n147, u2_u7_u4_n148, u2_u7_u4_n149, 
       u2_u7_u4_n150, u2_u7_u4_n151, u2_u7_u4_n152, u2_u7_u4_n153, u2_u7_u4_n154, u2_u7_u4_n155, u2_u7_u4_n156, u2_u7_u4_n157, u2_u7_u4_n158, 
       u2_u7_u4_n159, u2_u7_u4_n160, u2_u7_u4_n161, u2_u7_u4_n162, u2_u7_u4_n163, u2_u7_u4_n164, u2_u7_u4_n165, u2_u7_u4_n166, u2_u7_u4_n167, 
       u2_u7_u4_n168, u2_u7_u4_n169, u2_u7_u4_n170, u2_u7_u4_n171, u2_u7_u4_n172, u2_u7_u4_n173, u2_u7_u4_n174, u2_u7_u4_n175, u2_u7_u4_n176, 
       u2_u7_u4_n177, u2_u7_u4_n178, u2_u7_u4_n179, u2_u7_u4_n180, u2_u7_u4_n181, u2_u7_u4_n182, u2_u7_u4_n183, u2_u7_u4_n184, u2_u7_u4_n185, 
       u2_u7_u4_n186, u2_u7_u4_n94, u2_u7_u4_n95, u2_u7_u4_n96, u2_u7_u4_n97, u2_u7_u4_n98, u2_u7_u4_n99, u2_u7_u5_n100, u2_u7_u5_n101, 
       u2_u7_u5_n102, u2_u7_u5_n103, u2_u7_u5_n104, u2_u7_u5_n105, u2_u7_u5_n106, u2_u7_u5_n107, u2_u7_u5_n108, u2_u7_u5_n109, u2_u7_u5_n110, 
       u2_u7_u5_n111, u2_u7_u5_n112, u2_u7_u5_n113, u2_u7_u5_n114, u2_u7_u5_n115, u2_u7_u5_n116, u2_u7_u5_n117, u2_u7_u5_n118, u2_u7_u5_n119, 
       u2_u7_u5_n120, u2_u7_u5_n121, u2_u7_u5_n122, u2_u7_u5_n123, u2_u7_u5_n124, u2_u7_u5_n125, u2_u7_u5_n126, u2_u7_u5_n127, u2_u7_u5_n128, 
       u2_u7_u5_n129, u2_u7_u5_n130, u2_u7_u5_n131, u2_u7_u5_n132, u2_u7_u5_n133, u2_u7_u5_n134, u2_u7_u5_n135, u2_u7_u5_n136, u2_u7_u5_n137, 
       u2_u7_u5_n138, u2_u7_u5_n139, u2_u7_u5_n140, u2_u7_u5_n141, u2_u7_u5_n142, u2_u7_u5_n143, u2_u7_u5_n144, u2_u7_u5_n145, u2_u7_u5_n146, 
       u2_u7_u5_n147, u2_u7_u5_n148, u2_u7_u5_n149, u2_u7_u5_n150, u2_u7_u5_n151, u2_u7_u5_n152, u2_u7_u5_n153, u2_u7_u5_n154, u2_u7_u5_n155, 
       u2_u7_u5_n156, u2_u7_u5_n157, u2_u7_u5_n158, u2_u7_u5_n159, u2_u7_u5_n160, u2_u7_u5_n161, u2_u7_u5_n162, u2_u7_u5_n163, u2_u7_u5_n164, 
       u2_u7_u5_n165, u2_u7_u5_n166, u2_u7_u5_n167, u2_u7_u5_n168, u2_u7_u5_n169, u2_u7_u5_n170, u2_u7_u5_n171, u2_u7_u5_n172, u2_u7_u5_n173, 
       u2_u7_u5_n174, u2_u7_u5_n175, u2_u7_u5_n176, u2_u7_u5_n177, u2_u7_u5_n178, u2_u7_u5_n179, u2_u7_u5_n180, u2_u7_u5_n181, u2_u7_u5_n182, 
       u2_u7_u5_n183, u2_u7_u5_n184, u2_u7_u5_n185, u2_u7_u5_n186, u2_u7_u5_n187, u2_u7_u5_n188, u2_u7_u5_n189, u2_u7_u5_n190, u2_u7_u5_n191, 
       u2_u7_u5_n192, u2_u7_u5_n193, u2_u7_u5_n194, u2_u7_u5_n195, u2_u7_u5_n196, u2_u7_u5_n99, u2_u8_X_1, u2_u8_X_10, u2_u8_X_11, 
       u2_u8_X_12, u2_u8_X_13, u2_u8_X_14, u2_u8_X_15, u2_u8_X_16, u2_u8_X_17, u2_u8_X_18, u2_u8_X_19, u2_u8_X_2, 
       u2_u8_X_20, u2_u8_X_21, u2_u8_X_22, u2_u8_X_23, u2_u8_X_24, u2_u8_X_25, u2_u8_X_26, u2_u8_X_27, u2_u8_X_28, 
       u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u8_X_37, u2_u8_X_38, u2_u8_X_39, u2_u8_X_4, u2_u8_X_40, u2_u8_X_41, 
       u2_u8_X_42, u2_u8_X_43, u2_u8_X_44, u2_u8_X_45, u2_u8_X_46, u2_u8_X_47, u2_u8_X_48, u2_u8_X_5, u2_u8_X_6, 
       u2_u8_X_7, u2_u8_X_8, u2_u8_X_9, u2_u8_u0_n100, u2_u8_u0_n101, u2_u8_u0_n102, u2_u8_u0_n103, u2_u8_u0_n104, u2_u8_u0_n105, 
       u2_u8_u0_n106, u2_u8_u0_n107, u2_u8_u0_n108, u2_u8_u0_n109, u2_u8_u0_n110, u2_u8_u0_n111, u2_u8_u0_n112, u2_u8_u0_n113, u2_u8_u0_n114, 
       u2_u8_u0_n115, u2_u8_u0_n116, u2_u8_u0_n117, u2_u8_u0_n118, u2_u8_u0_n119, u2_u8_u0_n120, u2_u8_u0_n121, u2_u8_u0_n122, u2_u8_u0_n123, 
       u2_u8_u0_n124, u2_u8_u0_n125, u2_u8_u0_n126, u2_u8_u0_n127, u2_u8_u0_n128, u2_u8_u0_n129, u2_u8_u0_n130, u2_u8_u0_n131, u2_u8_u0_n132, 
       u2_u8_u0_n133, u2_u8_u0_n134, u2_u8_u0_n135, u2_u8_u0_n136, u2_u8_u0_n137, u2_u8_u0_n138, u2_u8_u0_n139, u2_u8_u0_n140, u2_u8_u0_n141, 
       u2_u8_u0_n142, u2_u8_u0_n143, u2_u8_u0_n144, u2_u8_u0_n145, u2_u8_u0_n146, u2_u8_u0_n147, u2_u8_u0_n148, u2_u8_u0_n149, u2_u8_u0_n150, 
       u2_u8_u0_n151, u2_u8_u0_n152, u2_u8_u0_n153, u2_u8_u0_n154, u2_u8_u0_n155, u2_u8_u0_n156, u2_u8_u0_n157, u2_u8_u0_n158, u2_u8_u0_n159, 
       u2_u8_u0_n160, u2_u8_u0_n161, u2_u8_u0_n162, u2_u8_u0_n163, u2_u8_u0_n164, u2_u8_u0_n165, u2_u8_u0_n166, u2_u8_u0_n167, u2_u8_u0_n168, 
       u2_u8_u0_n169, u2_u8_u0_n170, u2_u8_u0_n171, u2_u8_u0_n172, u2_u8_u0_n173, u2_u8_u0_n174, u2_u8_u0_n88, u2_u8_u0_n89, u2_u8_u0_n90, 
       u2_u8_u0_n91, u2_u8_u0_n92, u2_u8_u0_n93, u2_u8_u0_n94, u2_u8_u0_n95, u2_u8_u0_n96, u2_u8_u0_n97, u2_u8_u0_n98, u2_u8_u0_n99, 
       u2_u8_u1_n100, u2_u8_u1_n101, u2_u8_u1_n102, u2_u8_u1_n103, u2_u8_u1_n104, u2_u8_u1_n105, u2_u8_u1_n106, u2_u8_u1_n107, u2_u8_u1_n108, 
       u2_u8_u1_n109, u2_u8_u1_n110, u2_u8_u1_n111, u2_u8_u1_n112, u2_u8_u1_n113, u2_u8_u1_n114, u2_u8_u1_n115, u2_u8_u1_n116, u2_u8_u1_n117, 
       u2_u8_u1_n118, u2_u8_u1_n119, u2_u8_u1_n120, u2_u8_u1_n121, u2_u8_u1_n122, u2_u8_u1_n123, u2_u8_u1_n124, u2_u8_u1_n125, u2_u8_u1_n126, 
       u2_u8_u1_n127, u2_u8_u1_n128, u2_u8_u1_n129, u2_u8_u1_n130, u2_u8_u1_n131, u2_u8_u1_n132, u2_u8_u1_n133, u2_u8_u1_n134, u2_u8_u1_n135, 
       u2_u8_u1_n136, u2_u8_u1_n137, u2_u8_u1_n138, u2_u8_u1_n139, u2_u8_u1_n140, u2_u8_u1_n141, u2_u8_u1_n142, u2_u8_u1_n143, u2_u8_u1_n144, 
       u2_u8_u1_n145, u2_u8_u1_n146, u2_u8_u1_n147, u2_u8_u1_n148, u2_u8_u1_n149, u2_u8_u1_n150, u2_u8_u1_n151, u2_u8_u1_n152, u2_u8_u1_n153, 
       u2_u8_u1_n154, u2_u8_u1_n155, u2_u8_u1_n156, u2_u8_u1_n157, u2_u8_u1_n158, u2_u8_u1_n159, u2_u8_u1_n160, u2_u8_u1_n161, u2_u8_u1_n162, 
       u2_u8_u1_n163, u2_u8_u1_n164, u2_u8_u1_n165, u2_u8_u1_n166, u2_u8_u1_n167, u2_u8_u1_n168, u2_u8_u1_n169, u2_u8_u1_n170, u2_u8_u1_n171, 
       u2_u8_u1_n172, u2_u8_u1_n173, u2_u8_u1_n174, u2_u8_u1_n175, u2_u8_u1_n176, u2_u8_u1_n177, u2_u8_u1_n178, u2_u8_u1_n179, u2_u8_u1_n180, 
       u2_u8_u1_n181, u2_u8_u1_n182, u2_u8_u1_n183, u2_u8_u1_n184, u2_u8_u1_n185, u2_u8_u1_n186, u2_u8_u1_n187, u2_u8_u1_n188, u2_u8_u1_n95, 
       u2_u8_u1_n96, u2_u8_u1_n97, u2_u8_u1_n98, u2_u8_u1_n99, u2_u8_u2_n100, u2_u8_u2_n101, u2_u8_u2_n102, u2_u8_u2_n103, u2_u8_u2_n104, 
       u2_u8_u2_n105, u2_u8_u2_n106, u2_u8_u2_n107, u2_u8_u2_n108, u2_u8_u2_n109, u2_u8_u2_n110, u2_u8_u2_n111, u2_u8_u2_n112, u2_u8_u2_n113, 
       u2_u8_u2_n114, u2_u8_u2_n115, u2_u8_u2_n116, u2_u8_u2_n117, u2_u8_u2_n118, u2_u8_u2_n119, u2_u8_u2_n120, u2_u8_u2_n121, u2_u8_u2_n122, 
       u2_u8_u2_n123, u2_u8_u2_n124, u2_u8_u2_n125, u2_u8_u2_n126, u2_u8_u2_n127, u2_u8_u2_n128, u2_u8_u2_n129, u2_u8_u2_n130, u2_u8_u2_n131, 
       u2_u8_u2_n132, u2_u8_u2_n133, u2_u8_u2_n134, u2_u8_u2_n135, u2_u8_u2_n136, u2_u8_u2_n137, u2_u8_u2_n138, u2_u8_u2_n139, u2_u8_u2_n140, 
       u2_u8_u2_n141, u2_u8_u2_n142, u2_u8_u2_n143, u2_u8_u2_n144, u2_u8_u2_n145, u2_u8_u2_n146, u2_u8_u2_n147, u2_u8_u2_n148, u2_u8_u2_n149, 
       u2_u8_u2_n150, u2_u8_u2_n151, u2_u8_u2_n152, u2_u8_u2_n153, u2_u8_u2_n154, u2_u8_u2_n155, u2_u8_u2_n156, u2_u8_u2_n157, u2_u8_u2_n158, 
       u2_u8_u2_n159, u2_u8_u2_n160, u2_u8_u2_n161, u2_u8_u2_n162, u2_u8_u2_n163, u2_u8_u2_n164, u2_u8_u2_n165, u2_u8_u2_n166, u2_u8_u2_n167, 
       u2_u8_u2_n168, u2_u8_u2_n169, u2_u8_u2_n170, u2_u8_u2_n171, u2_u8_u2_n172, u2_u8_u2_n173, u2_u8_u2_n174, u2_u8_u2_n175, u2_u8_u2_n176, 
       u2_u8_u2_n177, u2_u8_u2_n178, u2_u8_u2_n179, u2_u8_u2_n180, u2_u8_u2_n181, u2_u8_u2_n182, u2_u8_u2_n183, u2_u8_u2_n184, u2_u8_u2_n185, 
       u2_u8_u2_n186, u2_u8_u2_n187, u2_u8_u2_n188, u2_u8_u2_n95, u2_u8_u2_n96, u2_u8_u2_n97, u2_u8_u2_n98, u2_u8_u2_n99, u2_u8_u3_n100, 
       u2_u8_u3_n101, u2_u8_u3_n102, u2_u8_u3_n103, u2_u8_u3_n104, u2_u8_u3_n105, u2_u8_u3_n106, u2_u8_u3_n107, u2_u8_u3_n108, u2_u8_u3_n109, 
       u2_u8_u3_n110, u2_u8_u3_n111, u2_u8_u3_n112, u2_u8_u3_n113, u2_u8_u3_n114, u2_u8_u3_n115, u2_u8_u3_n116, u2_u8_u3_n117, u2_u8_u3_n118, 
       u2_u8_u3_n119, u2_u8_u3_n120, u2_u8_u3_n121, u2_u8_u3_n122, u2_u8_u3_n123, u2_u8_u3_n124, u2_u8_u3_n125, u2_u8_u3_n126, u2_u8_u3_n127, 
       u2_u8_u3_n128, u2_u8_u3_n129, u2_u8_u3_n130, u2_u8_u3_n131, u2_u8_u3_n132, u2_u8_u3_n133, u2_u8_u3_n134, u2_u8_u3_n135, u2_u8_u3_n136, 
       u2_u8_u3_n137, u2_u8_u3_n138, u2_u8_u3_n139, u2_u8_u3_n140, u2_u8_u3_n141, u2_u8_u3_n142, u2_u8_u3_n143, u2_u8_u3_n144, u2_u8_u3_n145, 
       u2_u8_u3_n146, u2_u8_u3_n147, u2_u8_u3_n148, u2_u8_u3_n149, u2_u8_u3_n150, u2_u8_u3_n151, u2_u8_u3_n152, u2_u8_u3_n153, u2_u8_u3_n154, 
       u2_u8_u3_n155, u2_u8_u3_n156, u2_u8_u3_n157, u2_u8_u3_n158, u2_u8_u3_n159, u2_u8_u3_n160, u2_u8_u3_n161, u2_u8_u3_n162, u2_u8_u3_n163, 
       u2_u8_u3_n164, u2_u8_u3_n165, u2_u8_u3_n166, u2_u8_u3_n167, u2_u8_u3_n168, u2_u8_u3_n169, u2_u8_u3_n170, u2_u8_u3_n171, u2_u8_u3_n172, 
       u2_u8_u3_n173, u2_u8_u3_n174, u2_u8_u3_n175, u2_u8_u3_n176, u2_u8_u3_n177, u2_u8_u3_n178, u2_u8_u3_n179, u2_u8_u3_n180, u2_u8_u3_n181, 
       u2_u8_u3_n182, u2_u8_u3_n183, u2_u8_u3_n184, u2_u8_u3_n185, u2_u8_u3_n186, u2_u8_u3_n94, u2_u8_u3_n95, u2_u8_u3_n96, u2_u8_u3_n97, 
       u2_u8_u3_n98, u2_u8_u3_n99, u2_u8_u4_n100, u2_u8_u4_n101, u2_u8_u4_n102, u2_u8_u4_n103, u2_u8_u4_n104, u2_u8_u4_n105, u2_u8_u4_n106, 
       u2_u8_u4_n107, u2_u8_u4_n108, u2_u8_u4_n109, u2_u8_u4_n110, u2_u8_u4_n111, u2_u8_u4_n112, u2_u8_u4_n113, u2_u8_u4_n114, u2_u8_u4_n115, 
       u2_u8_u4_n116, u2_u8_u4_n117, u2_u8_u4_n118, u2_u8_u4_n119, u2_u8_u4_n120, u2_u8_u4_n121, u2_u8_u4_n122, u2_u8_u4_n123, u2_u8_u4_n124, 
       u2_u8_u4_n125, u2_u8_u4_n126, u2_u8_u4_n127, u2_u8_u4_n128, u2_u8_u4_n129, u2_u8_u4_n130, u2_u8_u4_n131, u2_u8_u4_n132, u2_u8_u4_n133, 
       u2_u8_u4_n134, u2_u8_u4_n135, u2_u8_u4_n136, u2_u8_u4_n137, u2_u8_u4_n138, u2_u8_u4_n139, u2_u8_u4_n140, u2_u8_u4_n141, u2_u8_u4_n142, 
       u2_u8_u4_n143, u2_u8_u4_n144, u2_u8_u4_n145, u2_u8_u4_n146, u2_u8_u4_n147, u2_u8_u4_n148, u2_u8_u4_n149, u2_u8_u4_n150, u2_u8_u4_n151, 
       u2_u8_u4_n152, u2_u8_u4_n153, u2_u8_u4_n154, u2_u8_u4_n155, u2_u8_u4_n156, u2_u8_u4_n157, u2_u8_u4_n158, u2_u8_u4_n159, u2_u8_u4_n160, 
       u2_u8_u4_n161, u2_u8_u4_n162, u2_u8_u4_n163, u2_u8_u4_n164, u2_u8_u4_n165, u2_u8_u4_n166, u2_u8_u4_n167, u2_u8_u4_n168, u2_u8_u4_n169, 
       u2_u8_u4_n170, u2_u8_u4_n171, u2_u8_u4_n172, u2_u8_u4_n173, u2_u8_u4_n174, u2_u8_u4_n175, u2_u8_u4_n176, u2_u8_u4_n177, u2_u8_u4_n178, 
       u2_u8_u4_n179, u2_u8_u4_n180, u2_u8_u4_n181, u2_u8_u4_n182, u2_u8_u4_n183, u2_u8_u4_n184, u2_u8_u4_n185, u2_u8_u4_n186, u2_u8_u4_n94, 
       u2_u8_u4_n95, u2_u8_u4_n96, u2_u8_u4_n97, u2_u8_u4_n98, u2_u8_u4_n99, u2_u8_u6_n100, u2_u8_u6_n101, u2_u8_u6_n102, u2_u8_u6_n103, 
       u2_u8_u6_n104, u2_u8_u6_n105, u2_u8_u6_n106, u2_u8_u6_n107, u2_u8_u6_n108, u2_u8_u6_n109, u2_u8_u6_n110, u2_u8_u6_n111, u2_u8_u6_n112, 
       u2_u8_u6_n113, u2_u8_u6_n114, u2_u8_u6_n115, u2_u8_u6_n116, u2_u8_u6_n117, u2_u8_u6_n118, u2_u8_u6_n119, u2_u8_u6_n120, u2_u8_u6_n121, 
       u2_u8_u6_n122, u2_u8_u6_n123, u2_u8_u6_n124, u2_u8_u6_n125, u2_u8_u6_n126, u2_u8_u6_n127, u2_u8_u6_n128, u2_u8_u6_n129, u2_u8_u6_n130, 
       u2_u8_u6_n131, u2_u8_u6_n132, u2_u8_u6_n133, u2_u8_u6_n134, u2_u8_u6_n135, u2_u8_u6_n136, u2_u8_u6_n137, u2_u8_u6_n138, u2_u8_u6_n139, 
       u2_u8_u6_n140, u2_u8_u6_n141, u2_u8_u6_n142, u2_u8_u6_n143, u2_u8_u6_n144, u2_u8_u6_n145, u2_u8_u6_n146, u2_u8_u6_n147, u2_u8_u6_n148, 
       u2_u8_u6_n149, u2_u8_u6_n150, u2_u8_u6_n151, u2_u8_u6_n152, u2_u8_u6_n153, u2_u8_u6_n154, u2_u8_u6_n155, u2_u8_u6_n156, u2_u8_u6_n157, 
       u2_u8_u6_n158, u2_u8_u6_n159, u2_u8_u6_n160, u2_u8_u6_n161, u2_u8_u6_n162, u2_u8_u6_n163, u2_u8_u6_n164, u2_u8_u6_n165, u2_u8_u6_n166, 
       u2_u8_u6_n167, u2_u8_u6_n168, u2_u8_u6_n169, u2_u8_u6_n170, u2_u8_u6_n171, u2_u8_u6_n172, u2_u8_u6_n173, u2_u8_u6_n174, u2_u8_u6_n88, 
       u2_u8_u6_n89, u2_u8_u6_n90, u2_u8_u6_n91, u2_u8_u6_n92, u2_u8_u6_n93, u2_u8_u6_n94, u2_u8_u6_n95, u2_u8_u6_n96, u2_u8_u6_n97, 
       u2_u8_u6_n98, u2_u8_u6_n99, u2_u8_u7_n100, u2_u8_u7_n101, u2_u8_u7_n102, u2_u8_u7_n103, u2_u8_u7_n104, u2_u8_u7_n105, u2_u8_u7_n106, 
       u2_u8_u7_n107, u2_u8_u7_n108, u2_u8_u7_n109, u2_u8_u7_n110, u2_u8_u7_n111, u2_u8_u7_n112, u2_u8_u7_n113, u2_u8_u7_n114, u2_u8_u7_n115, 
       u2_u8_u7_n116, u2_u8_u7_n117, u2_u8_u7_n118, u2_u8_u7_n119, u2_u8_u7_n120, u2_u8_u7_n121, u2_u8_u7_n122, u2_u8_u7_n123, u2_u8_u7_n124, 
       u2_u8_u7_n125, u2_u8_u7_n126, u2_u8_u7_n127, u2_u8_u7_n128, u2_u8_u7_n129, u2_u8_u7_n130, u2_u8_u7_n131, u2_u8_u7_n132, u2_u8_u7_n133, 
       u2_u8_u7_n134, u2_u8_u7_n135, u2_u8_u7_n136, u2_u8_u7_n137, u2_u8_u7_n138, u2_u8_u7_n139, u2_u8_u7_n140, u2_u8_u7_n141, u2_u8_u7_n142, 
       u2_u8_u7_n143, u2_u8_u7_n144, u2_u8_u7_n145, u2_u8_u7_n146, u2_u8_u7_n147, u2_u8_u7_n148, u2_u8_u7_n149, u2_u8_u7_n150, u2_u8_u7_n151, 
       u2_u8_u7_n152, u2_u8_u7_n153, u2_u8_u7_n154, u2_u8_u7_n155, u2_u8_u7_n156, u2_u8_u7_n157, u2_u8_u7_n158, u2_u8_u7_n159, u2_u8_u7_n160, 
       u2_u8_u7_n161, u2_u8_u7_n162, u2_u8_u7_n163, u2_u8_u7_n164, u2_u8_u7_n165, u2_u8_u7_n166, u2_u8_u7_n167, u2_u8_u7_n168, u2_u8_u7_n169, 
       u2_u8_u7_n170, u2_u8_u7_n171, u2_u8_u7_n172, u2_u8_u7_n173, u2_u8_u7_n174, u2_u8_u7_n175, u2_u8_u7_n176, u2_u8_u7_n177, u2_u8_u7_n178, 
       u2_u8_u7_n179, u2_u8_u7_n180, u2_u8_u7_n91, u2_u8_u7_n92, u2_u8_u7_n93, u2_u8_u7_n94, u2_u8_u7_n95, u2_u8_u7_n96, u2_u8_u7_n97, 
       u2_u8_u7_n98, u2_u8_u7_n99, u2_u9_X_19, u2_u9_X_20, u2_u9_X_21, u2_u9_X_22, u2_u9_X_23, u2_u9_X_24, u2_u9_X_25, 
       u2_u9_X_26, u2_u9_X_27, u2_u9_X_28, u2_u9_X_29, u2_u9_X_30, u2_u9_X_31, u2_u9_X_32, u2_u9_X_33, u2_u9_X_34, 
       u2_u9_X_35, u2_u9_X_36, u2_u9_X_37, u2_u9_X_38, u2_u9_X_39, u2_u9_X_40, u2_u9_X_41, u2_u9_X_42, u2_u9_u3_n100, 
       u2_u9_u3_n101, u2_u9_u3_n102, u2_u9_u3_n103, u2_u9_u3_n104, u2_u9_u3_n105, u2_u9_u3_n106, u2_u9_u3_n107, u2_u9_u3_n108, u2_u9_u3_n109, 
       u2_u9_u3_n110, u2_u9_u3_n111, u2_u9_u3_n112, u2_u9_u3_n113, u2_u9_u3_n114, u2_u9_u3_n115, u2_u9_u3_n116, u2_u9_u3_n117, u2_u9_u3_n118, 
       u2_u9_u3_n119, u2_u9_u3_n120, u2_u9_u3_n121, u2_u9_u3_n122, u2_u9_u3_n123, u2_u9_u3_n124, u2_u9_u3_n125, u2_u9_u3_n126, u2_u9_u3_n127, 
       u2_u9_u3_n128, u2_u9_u3_n129, u2_u9_u3_n130, u2_u9_u3_n131, u2_u9_u3_n132, u2_u9_u3_n133, u2_u9_u3_n134, u2_u9_u3_n135, u2_u9_u3_n136, 
       u2_u9_u3_n137, u2_u9_u3_n138, u2_u9_u3_n139, u2_u9_u3_n140, u2_u9_u3_n141, u2_u9_u3_n142, u2_u9_u3_n143, u2_u9_u3_n144, u2_u9_u3_n145, 
       u2_u9_u3_n146, u2_u9_u3_n147, u2_u9_u3_n148, u2_u9_u3_n149, u2_u9_u3_n150, u2_u9_u3_n151, u2_u9_u3_n152, u2_u9_u3_n153, u2_u9_u3_n154, 
       u2_u9_u3_n155, u2_u9_u3_n156, u2_u9_u3_n157, u2_u9_u3_n158, u2_u9_u3_n159, u2_u9_u3_n160, u2_u9_u3_n161, u2_u9_u3_n162, u2_u9_u3_n163, 
       u2_u9_u3_n164, u2_u9_u3_n165, u2_u9_u3_n166, u2_u9_u3_n167, u2_u9_u3_n168, u2_u9_u3_n169, u2_u9_u3_n170, u2_u9_u3_n171, u2_u9_u3_n172, 
       u2_u9_u3_n173, u2_u9_u3_n174, u2_u9_u3_n175, u2_u9_u3_n176, u2_u9_u3_n177, u2_u9_u3_n178, u2_u9_u3_n179, u2_u9_u3_n180, u2_u9_u3_n181, 
       u2_u9_u3_n182, u2_u9_u3_n183, u2_u9_u3_n184, u2_u9_u3_n185, u2_u9_u3_n186, u2_u9_u3_n94, u2_u9_u3_n95, u2_u9_u3_n96, u2_u9_u3_n97, 
       u2_u9_u3_n98, u2_u9_u3_n99, u2_u9_u4_n100, u2_u9_u4_n101, u2_u9_u4_n102, u2_u9_u4_n103, u2_u9_u4_n104, u2_u9_u4_n105, u2_u9_u4_n106, 
       u2_u9_u4_n107, u2_u9_u4_n108, u2_u9_u4_n109, u2_u9_u4_n110, u2_u9_u4_n111, u2_u9_u4_n112, u2_u9_u4_n113, u2_u9_u4_n114, u2_u9_u4_n115, 
       u2_u9_u4_n116, u2_u9_u4_n117, u2_u9_u4_n118, u2_u9_u4_n119, u2_u9_u4_n120, u2_u9_u4_n121, u2_u9_u4_n122, u2_u9_u4_n123, u2_u9_u4_n124, 
       u2_u9_u4_n125, u2_u9_u4_n126, u2_u9_u4_n127, u2_u9_u4_n128, u2_u9_u4_n129, u2_u9_u4_n130, u2_u9_u4_n131, u2_u9_u4_n132, u2_u9_u4_n133, 
       u2_u9_u4_n134, u2_u9_u4_n135, u2_u9_u4_n136, u2_u9_u4_n137, u2_u9_u4_n138, u2_u9_u4_n139, u2_u9_u4_n140, u2_u9_u4_n141, u2_u9_u4_n142, 
       u2_u9_u4_n143, u2_u9_u4_n144, u2_u9_u4_n145, u2_u9_u4_n146, u2_u9_u4_n147, u2_u9_u4_n148, u2_u9_u4_n149, u2_u9_u4_n150, u2_u9_u4_n151, 
       u2_u9_u4_n152, u2_u9_u4_n153, u2_u9_u4_n154, u2_u9_u4_n155, u2_u9_u4_n156, u2_u9_u4_n157, u2_u9_u4_n158, u2_u9_u4_n159, u2_u9_u4_n160, 
       u2_u9_u4_n161, u2_u9_u4_n162, u2_u9_u4_n163, u2_u9_u4_n164, u2_u9_u4_n165, u2_u9_u4_n166, u2_u9_u4_n167, u2_u9_u4_n168, u2_u9_u4_n169, 
       u2_u9_u4_n170, u2_u9_u4_n171, u2_u9_u4_n172, u2_u9_u4_n173, u2_u9_u4_n174, u2_u9_u4_n175, u2_u9_u4_n176, u2_u9_u4_n177, u2_u9_u4_n178, 
       u2_u9_u4_n179, u2_u9_u4_n180, u2_u9_u4_n181, u2_u9_u4_n182, u2_u9_u4_n183, u2_u9_u4_n184, u2_u9_u4_n185, u2_u9_u4_n186, u2_u9_u4_n94, 
       u2_u9_u4_n95, u2_u9_u4_n96, u2_u9_u4_n97, u2_u9_u4_n98, u2_u9_u4_n99, u2_u9_u5_n100, u2_u9_u5_n101, u2_u9_u5_n102, u2_u9_u5_n103, 
       u2_u9_u5_n104, u2_u9_u5_n105, u2_u9_u5_n106, u2_u9_u5_n107, u2_u9_u5_n108, u2_u9_u5_n109, u2_u9_u5_n110, u2_u9_u5_n111, u2_u9_u5_n112, 
       u2_u9_u5_n113, u2_u9_u5_n114, u2_u9_u5_n115, u2_u9_u5_n116, u2_u9_u5_n117, u2_u9_u5_n118, u2_u9_u5_n119, u2_u9_u5_n120, u2_u9_u5_n121, 
       u2_u9_u5_n122, u2_u9_u5_n123, u2_u9_u5_n124, u2_u9_u5_n125, u2_u9_u5_n126, u2_u9_u5_n127, u2_u9_u5_n128, u2_u9_u5_n129, u2_u9_u5_n130, 
       u2_u9_u5_n131, u2_u9_u5_n132, u2_u9_u5_n133, u2_u9_u5_n134, u2_u9_u5_n135, u2_u9_u5_n136, u2_u9_u5_n137, u2_u9_u5_n138, u2_u9_u5_n139, 
       u2_u9_u5_n140, u2_u9_u5_n141, u2_u9_u5_n142, u2_u9_u5_n143, u2_u9_u5_n144, u2_u9_u5_n145, u2_u9_u5_n146, u2_u9_u5_n147, u2_u9_u5_n148, 
       u2_u9_u5_n149, u2_u9_u5_n150, u2_u9_u5_n151, u2_u9_u5_n152, u2_u9_u5_n153, u2_u9_u5_n154, u2_u9_u5_n155, u2_u9_u5_n156, u2_u9_u5_n157, 
       u2_u9_u5_n158, u2_u9_u5_n159, u2_u9_u5_n160, u2_u9_u5_n161, u2_u9_u5_n162, u2_u9_u5_n163, u2_u9_u5_n164, u2_u9_u5_n165, u2_u9_u5_n166, 
       u2_u9_u5_n167, u2_u9_u5_n168, u2_u9_u5_n169, u2_u9_u5_n170, u2_u9_u5_n171, u2_u9_u5_n172, u2_u9_u5_n173, u2_u9_u5_n174, u2_u9_u5_n175, 
       u2_u9_u5_n176, u2_u9_u5_n177, u2_u9_u5_n178, u2_u9_u5_n179, u2_u9_u5_n180, u2_u9_u5_n181, u2_u9_u5_n182, u2_u9_u5_n183, u2_u9_u5_n184, 
       u2_u9_u5_n185, u2_u9_u5_n186, u2_u9_u5_n187, u2_u9_u5_n188, u2_u9_u5_n189, u2_u9_u5_n190, u2_u9_u5_n191, u2_u9_u5_n192, u2_u9_u5_n193, 
       u2_u9_u5_n194, u2_u9_u5_n195, u2_u9_u5_n196, u2_u9_u5_n99, u2_u9_u6_n100, u2_u9_u6_n101, u2_u9_u6_n102, u2_u9_u6_n103, u2_u9_u6_n104, 
       u2_u9_u6_n105, u2_u9_u6_n106, u2_u9_u6_n107, u2_u9_u6_n108, u2_u9_u6_n109, u2_u9_u6_n110, u2_u9_u6_n111, u2_u9_u6_n112, u2_u9_u6_n113, 
       u2_u9_u6_n114, u2_u9_u6_n115, u2_u9_u6_n116, u2_u9_u6_n117, u2_u9_u6_n118, u2_u9_u6_n119, u2_u9_u6_n120, u2_u9_u6_n121, u2_u9_u6_n122, 
       u2_u9_u6_n123, u2_u9_u6_n124, u2_u9_u6_n125, u2_u9_u6_n126, u2_u9_u6_n127, u2_u9_u6_n128, u2_u9_u6_n129, u2_u9_u6_n130, u2_u9_u6_n131, 
       u2_u9_u6_n132, u2_u9_u6_n133, u2_u9_u6_n134, u2_u9_u6_n135, u2_u9_u6_n136, u2_u9_u6_n137, u2_u9_u6_n138, u2_u9_u6_n139, u2_u9_u6_n140, 
       u2_u9_u6_n141, u2_u9_u6_n142, u2_u9_u6_n143, u2_u9_u6_n144, u2_u9_u6_n145, u2_u9_u6_n146, u2_u9_u6_n147, u2_u9_u6_n148, u2_u9_u6_n149, 
       u2_u9_u6_n150, u2_u9_u6_n151, u2_u9_u6_n152, u2_u9_u6_n153, u2_u9_u6_n154, u2_u9_u6_n155, u2_u9_u6_n156, u2_u9_u6_n157, u2_u9_u6_n158, 
       u2_u9_u6_n159, u2_u9_u6_n160, u2_u9_u6_n161, u2_u9_u6_n162, u2_u9_u6_n163, u2_u9_u6_n164, u2_u9_u6_n165, u2_u9_u6_n166, u2_u9_u6_n167, 
       u2_u9_u6_n168, u2_u9_u6_n169, u2_u9_u6_n170, u2_u9_u6_n171, u2_u9_u6_n172, u2_u9_u6_n173, u2_u9_u6_n174, u2_u9_u6_n88, u2_u9_u6_n89, 
       u2_u9_u6_n90, u2_u9_u6_n91, u2_u9_u6_n92, u2_u9_u6_n93, u2_u9_u6_n94, u2_u9_u6_n95, u2_u9_u6_n96, u2_u9_u6_n97, u2_u9_u6_n98, 
       u2_u9_u6_n99, u2_uk_n1004, u2_uk_n1005, u2_uk_n1009, u2_uk_n1010, u2_uk_n1020, u2_uk_n1023, u2_uk_n1037, u2_uk_n1048, 
       u2_uk_n1050, u2_uk_n1051, u2_uk_n1052, u2_uk_n1058, u2_uk_n1066, u2_uk_n1068, u2_uk_n1071, u2_uk_n1072, u2_uk_n1088, 
       u2_uk_n1091, u2_uk_n1103, u2_uk_n1106, u2_uk_n1117, u2_uk_n1118, u2_uk_n1122, u2_uk_n1123, u2_uk_n1124, u2_uk_n1126, 
       u2_uk_n1127, u2_uk_n1129, u2_uk_n1135, u2_uk_n1138, u2_uk_n1139, u2_uk_n1147, u2_uk_n1151, u2_uk_n1157, u2_uk_n1158, 
       u2_uk_n1165, u2_uk_n252, u2_uk_n271, u2_uk_n277, u2_uk_n279, u2_uk_n291, u2_uk_n294, u2_uk_n297, u2_uk_n301, 
       u2_uk_n305, u2_uk_n306, u2_uk_n335, u2_uk_n375, u2_uk_n382, u2_uk_n386, u2_uk_n454, u2_uk_n460, u2_uk_n496, 
       u2_uk_n501, u2_uk_n509, u2_uk_n524, u2_uk_n582, u2_uk_n587, u2_uk_n590, u2_uk_n601, u2_uk_n603, u2_uk_n634, 
       u2_uk_n662, u2_uk_n671, u2_uk_n678, u2_uk_n681, u2_uk_n936, u2_uk_n937, u2_uk_n949, u2_uk_n950, u2_uk_n951, 
       u2_uk_n952, u2_uk_n953, u2_uk_n975, u2_uk_n976, u2_uk_n977, u2_uk_n980, u2_uk_n981, u2_uk_n982, u2_uk_n985, 
       u2_uk_n987, u2_uk_n989, u2_uk_n991, u2_uk_n992, u2_uk_n993,  u2_uk_n995;
  XOR2_X1 u0_U100 (.B( u0_L12_27 ) , .Z( u0_N442 ) , .A( u0_out13_27 ) );
  XOR2_X1 u0_U106 (.B( u0_L12_22 ) , .Z( u0_N437 ) , .A( u0_out13_22 ) );
  XOR2_X1 u0_U107 (.B( u0_L12_21 ) , .Z( u0_N436 ) , .A( u0_out13_21 ) );
  XOR2_X1 u0_U113 (.B( u0_L12_15 ) , .Z( u0_N430 ) , .A( u0_out13_15 ) );
  XOR2_X1 u0_U117 (.B( u0_L12_12 ) , .Z( u0_N427 ) , .A( u0_out13_12 ) );
  XOR2_X1 u0_U122 (.B( u0_L12_7 ) , .Z( u0_N422 ) , .A( u0_out13_7 ) );
  XOR2_X1 u0_U124 (.B( u0_L12_5 ) , .Z( u0_N420 ) , .A( u0_out13_5 ) );
  XOR2_X1 u0_U148 (.Z( u0_N4 ) , .B( u0_desIn_r_38 ) , .A( u0_out0_5 ) );
  XOR2_X1 u0_U247 (.Z( u0_N31 ) , .B( u0_desIn_r_56 ) , .A( u0_out0_32 ) );
  XOR2_X1 u0_U259 (.Z( u0_N3 ) , .B( u0_desIn_r_30 ) , .A( u0_out0_4 ) );
  XOR2_X1 u0_U281 (.Z( u0_N28 ) , .B( u0_desIn_r_32 ) , .A( u0_out0_29 ) );
  XOR2_X1 u0_U303 (.Z( u0_N26 ) , .B( u0_desIn_r_16 ) , .A( u0_out0_27 ) );
  XOR2_X1 u0_U325 (.Z( u0_N24 ) , .B( u0_desIn_r_0 ) , .A( u0_out0_25 ) );
  XOR2_X1 u0_U35 (.Z( u0_N7 ) , .B( u0_desIn_r_62 ) , .A( u0_out0_8 ) );
  XOR2_X1 u0_U358 (.Z( u0_N21 ) , .B( u0_desIn_r_42 ) , .A( u0_out0_22 ) );
  XOR2_X1 u0_U369 (.Z( u0_N20 ) , .B( u0_desIn_r_34 ) , .A( u0_out0_21 ) );
  XOR2_X1 u0_U370 (.Z( u0_N2 ) , .B( u0_desIn_r_22 ) , .A( u0_out0_3 ) );
  XOR2_X1 u0_U392 (.Z( u0_N18 ) , .B( u0_desIn_r_18 ) , .A( u0_out0_19 ) );
  XOR2_X1 u0_U415 (.B( u0_L3_32 ) , .Z( u0_N159 ) , .A( u0_out4_32 ) );
  XOR2_X1 u0_U416 (.B( u0_L3_31 ) , .Z( u0_N158 ) , .A( u0_out4_31 ) );
  XOR2_X1 u0_U418 (.B( u0_L3_29 ) , .Z( u0_N156 ) , .A( u0_out4_29 ) );
  XOR2_X1 u0_U420 (.B( u0_L3_27 ) , .Z( u0_N154 ) , .A( u0_out4_27 ) );
  XOR2_X1 u0_U424 (.B( u0_L3_23 ) , .Z( u0_N150 ) , .A( u0_out4_23 ) );
  XOR2_X1 u0_U426 (.B( u0_L3_22 ) , .Z( u0_N149 ) , .A( u0_out4_22 ) );
  XOR2_X1 u0_U427 (.B( u0_L3_21 ) , .Z( u0_N148 ) , .A( u0_out4_21 ) );
  XOR2_X1 u0_U429 (.B( u0_L3_19 ) , .Z( u0_N146 ) , .A( u0_out4_19 ) );
  XOR2_X1 u0_U431 (.B( u0_L3_17 ) , .Z( u0_N144 ) , .A( u0_out4_17 ) );
  XOR2_X1 u0_U433 (.B( u0_L3_15 ) , .Z( u0_N142 ) , .A( u0_out4_15 ) );
  XOR2_X1 u0_U436 (.Z( u0_N14 ) , .B( u0_desIn_r_52 ) , .A( u0_out0_15 ) );
  XOR2_X1 u0_U437 (.B( u0_L3_12 ) , .Z( u0_N139 ) , .A( u0_out4_12 ) );
  XOR2_X1 u0_U438 (.B( u0_L3_11 ) , .Z( u0_N138 ) , .A( u0_out4_11 ) );
  XOR2_X1 u0_U440 (.B( u0_L3_9 ) , .Z( u0_N136 ) , .A( u0_out4_9 ) );
  XOR2_X1 u0_U442 (.B( u0_L3_7 ) , .Z( u0_N134 ) , .A( u0_out4_7 ) );
  XOR2_X1 u0_U444 (.B( u0_L3_5 ) , .Z( u0_N132 ) , .A( u0_out4_5 ) );
  XOR2_X1 u0_U445 (.B( u0_L3_4 ) , .Z( u0_N131 ) , .A( u0_out4_4 ) );
  XOR2_X1 u0_U447 (.Z( u0_N13 ) , .B( u0_desIn_r_44 ) , .A( u0_out0_14 ) );
  XOR2_X1 u0_U46 (.Z( u0_N6 ) , .B( u0_desIn_r_54 ) , .A( u0_out0_7 ) );
  XOR2_X1 u0_U469 (.Z( u0_N11 ) , .B( u0_desIn_r_28 ) , .A( u0_out0_12 ) );
  XOR2_X1 u0_U480 (.Z( u0_N10 ) , .B( u0_desIn_r_20 ) , .A( u0_out0_11 ) );
  XOR2_X1 u0_U95 (.B( u0_L12_32 ) , .Z( u0_N447 ) , .A( u0_out13_32 ) );
  XOR2_X1 u0_u0_U10 (.B( u0_K1_45 ) , .A( u0_desIn_r_41 ) , .Z( u0_u0_X_45 ) );
  XOR2_X1 u0_u0_U11 (.B( u0_K1_44 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_44 ) );
  XOR2_X1 u0_u0_U12 (.B( u0_K1_43 ) , .A( u0_desIn_r_25 ) , .Z( u0_u0_X_43 ) );
  XOR2_X1 u0_u0_U13 (.B( u0_K1_42 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_42 ) );
  XOR2_X1 u0_u0_U14 (.B( u0_K1_41 ) , .A( u0_desIn_r_25 ) , .Z( u0_u0_X_41 ) );
  XOR2_X1 u0_u0_U15 (.B( u0_K1_40 ) , .A( u0_desIn_r_17 ) , .Z( u0_u0_X_40 ) );
  XOR2_X1 u0_u0_U17 (.B( u0_K1_39 ) , .A( u0_desIn_r_9 ) , .Z( u0_u0_X_39 ) );
  XOR2_X1 u0_u0_U18 (.B( u0_K1_38 ) , .A( u0_desIn_r_1 ) , .Z( u0_u0_X_38 ) );
  XOR2_X1 u0_u0_U19 (.B( u0_K1_37 ) , .A( u0_desIn_r_59 ) , .Z( u0_u0_X_37 ) );
  XOR2_X1 u0_u0_U20 (.B( u0_K1_36 ) , .A( u0_desIn_r_1 ) , .Z( u0_u0_X_36 ) );
  XOR2_X1 u0_u0_U21 (.B( u0_K1_35 ) , .A( u0_desIn_r_59 ) , .Z( u0_u0_X_35 ) );
  XOR2_X1 u0_u0_U22 (.B( u0_K1_34 ) , .A( u0_desIn_r_51 ) , .Z( u0_u0_X_34 ) );
  XOR2_X1 u0_u0_U23 (.B( u0_K1_33 ) , .A( u0_desIn_r_43 ) , .Z( u0_u0_X_33 ) );
  XOR2_X1 u0_u0_U24 (.B( u0_K1_32 ) , .A( u0_desIn_r_35 ) , .Z( u0_u0_X_32 ) );
  XOR2_X1 u0_u0_U25 (.B( u0_K1_31 ) , .A( u0_desIn_r_27 ) , .Z( u0_u0_X_31 ) );
  XOR2_X1 u0_u0_U26 (.B( u0_K1_30 ) , .A( u0_desIn_r_35 ) , .Z( u0_u0_X_30 ) );
  XOR2_X1 u0_u0_U28 (.B( u0_K1_29 ) , .A( u0_desIn_r_27 ) , .Z( u0_u0_X_29 ) );
  XOR2_X1 u0_u0_U29 (.B( u0_K1_28 ) , .A( u0_desIn_r_19 ) , .Z( u0_u0_X_28 ) );
  XOR2_X1 u0_u0_U30 (.B( u0_K1_27 ) , .A( u0_desIn_r_11 ) , .Z( u0_u0_X_27 ) );
  XOR2_X1 u0_u0_U31 (.B( u0_K1_26 ) , .A( u0_desIn_r_3 ) , .Z( u0_u0_X_26 ) );
  XOR2_X1 u0_u0_U32 (.B( u0_K1_25 ) , .A( u0_desIn_r_61 ) , .Z( u0_u0_X_25 ) );
  XOR2_X1 u0_u0_U7 (.B( u0_K1_48 ) , .A( u0_desIn_r_7 ) , .Z( u0_u0_X_48 ) );
  XOR2_X1 u0_u0_U8 (.B( u0_K1_47 ) , .A( u0_desIn_r_57 ) , .Z( u0_u0_X_47 ) );
  XOR2_X1 u0_u0_U9 (.B( u0_K1_46 ) , .A( u0_desIn_r_49 ) , .Z( u0_u0_X_46 ) );
  OAI22_X1 u0_u0_u4_U10 (.A2( u0_u0_u4_n16 ) , .A1( u0_u0_u4_n32 ) , .B1( u0_u0_u4_n34 ) , .ZN( u0_u0_u4_n50 ) , .B2( u0_u0_u4_n52 ) );
  AND3_X1 u0_u0_u4_U11 (.A1( u0_u0_u4_n30 ) , .A3( u0_u0_u4_n42 ) , .ZN( u0_u0_u4_n52 ) , .A2( u0_u0_u4_n53 ) );
  NAND2_X1 u0_u0_u4_U12 (.A1( u0_u0_u4_n14 ) , .A2( u0_u0_u4_n17 ) , .ZN( u0_u0_u4_n55 ) );
  AOI21_X1 u0_u0_u4_U13 (.A( u0_u0_u4_n17 ) , .ZN( u0_u0_u4_n25 ) , .B1( u0_u0_u4_n26 ) , .B2( u0_u0_u4_n27 ) );
  AOI21_X1 u0_u0_u4_U14 (.A( u0_u0_u4_n13 ) , .B1( u0_u0_u4_n3 ) , .B2( u0_u0_u4_n44 ) , .ZN( u0_u0_u4_n80 ) );
  AOI21_X1 u0_u0_u4_U15 (.A( u0_u0_u4_n13 ) , .ZN( u0_u0_u4_n24 ) , .B1( u0_u0_u4_n28 ) , .B2( u0_u0_u4_n29 ) );
  AOI21_X1 u0_u0_u4_U16 (.ZN( u0_u0_u4_n22 ) , .B1( u0_u0_u4_n32 ) , .B2( u0_u0_u4_n33 ) , .A( u0_u0_u4_n34 ) );
  AOI21_X1 u0_u0_u4_U17 (.ZN( u0_u0_u4_n23 ) , .B1( u0_u0_u4_n3 ) , .B2( u0_u0_u4_n30 ) , .A( u0_u0_u4_n31 ) );
  INV_X1 u0_u0_u4_U18 (.ZN( u0_u0_u4_n17 ) , .A( u0_u0_u4_n49 ) );
  AND2_X1 u0_u0_u4_U19 (.A1( u0_u0_u4_n27 ) , .ZN( u0_u0_u4_n32 ) , .A2( u0_u0_u4_n67 ) );
  INV_X1 u0_u0_u4_U20 (.ZN( u0_u0_u4_n12 ) , .A( u0_u0_u4_n31 ) );
  NAND2_X1 u0_u0_u4_U21 (.A1( u0_u0_u4_n40 ) , .ZN( u0_u0_u4_n56 ) , .A2( u0_u0_u4_n69 ) );
  NAND2_X1 u0_u0_u4_U22 (.ZN( u0_u0_u4_n57 ) , .A2( u0_u0_u4_n67 ) , .A1( u0_u0_u4_n68 ) );
  NAND2_X1 u0_u0_u4_U23 (.A1( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n69 ) , .ZN( u0_u0_u4_n70 ) );
  NAND2_X1 u0_u0_u4_U24 (.A2( u0_u0_u4_n39 ) , .A1( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n58 ) );
  AND3_X1 u0_u0_u4_U25 (.ZN( u0_u0_u4_n26 ) , .A3( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n44 ) , .A1( u0_u0_u4_n68 ) );
  AND2_X1 u0_u0_u4_U26 (.ZN( u0_u0_u4_n28 ) , .A2( u0_u0_u4_n40 ) , .A1( u0_u0_u4_n42 ) );
  OR3_X1 u0_u0_u4_U27 (.ZN( u0_u0_u4_n51 ) , .A1( u0_u0_u4_n71 ) , .A2( u0_u0_u4_n72 ) , .A3( u0_u0_u4_n73 ) );
  AOI21_X1 u0_u0_u4_U28 (.B1( u0_u0_u4_n13 ) , .B2( u0_u0_u4_n14 ) , .ZN( u0_u0_u4_n71 ) , .A( u0_u0_u4_n74 ) );
  AOI21_X1 u0_u0_u4_U29 (.A( u0_u0_u4_n31 ) , .B1( u0_u0_u4_n41 ) , .B2( u0_u0_u4_n42 ) , .ZN( u0_u0_u4_n72 ) );
  NOR2_X1 u0_u0_u4_U3 (.A2( u0_u0_u4_n5 ) , .A1( u0_u0_u4_n6 ) , .ZN( u0_u0_u4_n66 ) );
  OAI22_X1 u0_u0_u4_U30 (.A1( u0_u0_u4_n16 ) , .B2( u0_u0_u4_n17 ) , .B1( u0_u0_u4_n27 ) , .A2( u0_u0_u4_n66 ) , .ZN( u0_u0_u4_n73 ) );
  INV_X1 u0_u0_u4_U31 (.A( u0_u0_u4_n29 ) , .ZN( u0_u0_u4_n5 ) );
  INV_X1 u0_u0_u4_U32 (.ZN( u0_u0_u4_n6 ) , .A( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U33 (.A( u0_u0_u4_n43 ) , .ZN( u0_u0_u4_n8 ) );
  INV_X1 u0_u0_u4_U34 (.A( u0_u0_u4_n30 ) , .ZN( u0_u0_u4_n9 ) );
  NAND2_X1 u0_u0_u4_U35 (.A2( u0_u0_u4_n33 ) , .ZN( u0_u0_u4_n90 ) , .A1( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U36 (.ZN( u0_u0_u4_n1 ) , .A( u0_u0_u4_n92 ) );
  OAI221_X1 u0_u0_u4_U37 (.C2( u0_u0_u4_n14 ) , .B2( u0_u0_u4_n16 ) , .B1( u0_u0_u4_n29 ) , .C1( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n92 ) , .A( u0_u0_u4_n93 ) );
  AOI222_X1 u0_u0_u4_U38 (.C2( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n2 ) , .A1( u0_u0_u4_n49 ) , .B2( u0_u0_u4_n55 ) , .C1( u0_u0_u4_n6 ) , .A2( u0_u0_u4_n8 ) , .ZN( u0_u0_u4_n93 ) );
  INV_X1 u0_u0_u4_U39 (.ZN( u0_u0_u4_n2 ) , .A( u0_u0_u4_n74 ) );
  INV_X1 u0_u0_u4_U4 (.ZN( u0_u0_u4_n3 ) , .A( u0_u0_u4_n70 ) );
  INV_X1 u0_u0_u4_U40 (.ZN( u0_u0_u4_n4 ) , .A( u0_u0_u4_n44 ) );
  NOR2_X1 u0_u0_u4_U41 (.A2( u0_u0_u4_n18 ) , .A1( u0_u0_u4_n19 ) , .ZN( u0_u0_u4_n49 ) );
  NOR2_X1 u0_u0_u4_U42 (.ZN( u0_u0_u4_n34 ) , .A2( u0_u0_u4_n35 ) , .A1( u0_u0_u4_n37 ) );
  NOR2_X1 u0_u0_u4_U43 (.ZN( u0_u0_u4_n31 ) , .A1( u0_u0_u4_n49 ) , .A2( u0_u0_u4_n59 ) );
  AOI22_X1 u0_u0_u4_U44 (.A2( u0_u0_u4_n15 ) , .B1( u0_u0_u4_n59 ) , .ZN( u0_u0_u4_n63 ) , .A1( u0_u0_u4_n64 ) , .B2( u0_u0_u4_n65 ) );
  INV_X1 u0_u0_u4_U45 (.ZN( u0_u0_u4_n15 ) , .A( u0_u0_u4_n34 ) );
  NAND2_X1 u0_u0_u4_U46 (.A1( u0_u0_u4_n26 ) , .ZN( u0_u0_u4_n64 ) , .A2( u0_u0_u4_n67 ) );
  AOI22_X1 u0_u0_u4_U47 (.A1( u0_u0_u4_n37 ) , .ZN( u0_u0_u4_n47 ) , .A2( u0_u0_u4_n54 ) , .B2( u0_u0_u4_n55 ) , .B1( u0_u0_u4_n8 ) );
  NAND2_X1 u0_u0_u4_U48 (.A1( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n41 ) , .ZN( u0_u0_u4_n54 ) );
  NAND2_X1 u0_u0_u4_U49 (.ZN( u0_u0_u4_n33 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n89 ) );
  NOR4_X1 u0_u0_u4_U5 (.ZN( u0_u0_u4_n77 ) , .A1( u0_u0_u4_n78 ) , .A2( u0_u0_u4_n79 ) , .A3( u0_u0_u4_n80 ) , .A4( u0_u0_u4_n81 ) );
  NAND2_X1 u0_u0_u4_U50 (.ZN( u0_u0_u4_n29 ) , .A1( u0_u0_u4_n86 ) , .A2( u0_u0_u4_n88 ) );
  AOI21_X1 u0_u0_u4_U51 (.B2( u0_u0_u4_n37 ) , .A( u0_u0_u4_n51 ) , .ZN( u0_u0_u4_n60 ) , .B1( u0_u0_u4_n7 ) );
  INV_X1 u0_u0_u4_U52 (.A( u0_u0_u4_n27 ) , .ZN( u0_u0_u4_n7 ) );
  NAND2_X1 u0_u0_u4_U53 (.ZN( u0_u0_u4_n41 ) , .A1( u0_u0_u4_n82 ) , .A2( u0_u0_u4_n83 ) );
  NAND2_X1 u0_u0_u4_U54 (.ZN( u0_u0_u4_n27 ) , .A1( u0_u0_u4_n85 ) , .A2( u0_u0_u4_n86 ) );
  NAND2_X1 u0_u0_u4_U55 (.ZN( u0_u0_u4_n53 ) , .A2( u0_u0_u4_n88 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U56 (.ZN( u0_u0_u4_n44 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n84 ) );
  NAND2_X1 u0_u0_u4_U57 (.ZN( u0_u0_u4_n42 ) , .A2( u0_u0_u4_n82 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U58 (.ZN( u0_u0_u4_n67 ) , .A2( u0_u0_u4_n82 ) , .A1( u0_u0_u4_n87 ) );
  NAND2_X1 u0_u0_u4_U59 (.ZN( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n85 ) );
  AOI21_X1 u0_u0_u4_U6 (.A( u0_u0_u4_n17 ) , .B1( u0_u0_u4_n29 ) , .B2( u0_u0_u4_n41 ) , .ZN( u0_u0_u4_n81 ) );
  NAND2_X1 u0_u0_u4_U60 (.ZN( u0_u0_u4_n30 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n87 ) );
  INV_X1 u0_u0_u4_U61 (.ZN( u0_u0_u4_n14 ) , .A( u0_u0_u4_n37 ) );
  INV_X1 u0_u0_u4_U62 (.ZN( u0_u0_u4_n16 ) , .A( u0_u0_u4_n35 ) );
  NAND2_X1 u0_u0_u4_U63 (.ZN( u0_u0_u4_n69 ) , .A1( u0_u0_u4_n87 ) , .A2( u0_u0_u4_n88 ) );
  NAND2_X1 u0_u0_u4_U64 (.ZN( u0_u0_u4_n43 ) , .A1( u0_u0_u4_n85 ) , .A2( u0_u0_u4_n87 ) );
  NAND2_X1 u0_u0_u4_U65 (.A1( u0_u0_u4_n82 ) , .A2( u0_u0_u4_n86 ) , .ZN( u0_u0_u4_n91 ) );
  INV_X1 u0_u0_u4_U66 (.ZN( u0_u0_u4_n13 ) , .A( u0_u0_u4_n59 ) );
  NAND2_X1 u0_u0_u4_U67 (.ZN( u0_u0_u4_n68 ) , .A2( u0_u0_u4_n85 ) , .A1( u0_u0_u4_n89 ) );
  NAND2_X1 u0_u0_u4_U68 (.ZN( u0_u0_u4_n40 ) , .A1( u0_u0_u4_n84 ) , .A2( u0_u0_u4_n86 ) );
  NAND2_X1 u0_u0_u4_U69 (.ZN( u0_u0_u4_n74 ) , .A2( u0_u0_u4_n83 ) , .A1( u0_u0_u4_n88 ) );
  AOI21_X1 u0_u0_u4_U7 (.A( u0_u0_u4_n31 ) , .B1( u0_u0_u4_n32 ) , .B2( u0_u0_u4_n53 ) , .ZN( u0_u0_u4_n79 ) );
  NOR2_X1 u0_u0_u4_U70 (.A2( u0_u0_X_28 ) , .A1( u0_u0_u4_n19 ) , .ZN( u0_u0_u4_n37 ) );
  NOR2_X1 u0_u0_u4_U71 (.A2( u0_u0_X_29 ) , .A1( u0_u0_u4_n18 ) , .ZN( u0_u0_u4_n35 ) );
  NOR2_X1 u0_u0_u4_U72 (.A2( u0_u0_X_30 ) , .A1( u0_u0_u4_n11 ) , .ZN( u0_u0_u4_n82 ) );
  NOR2_X1 u0_u0_u4_U73 (.A2( u0_u0_X_26 ) , .A1( u0_u0_u4_n10 ) , .ZN( u0_u0_u4_n87 ) );
  NOR2_X1 u0_u0_u4_U74 (.A2( u0_u0_X_28 ) , .A1( u0_u0_X_29 ) , .ZN( u0_u0_u4_n59 ) );
  NOR2_X1 u0_u0_u4_U75 (.A2( u0_u0_X_27 ) , .A1( u0_u0_X_30 ) , .ZN( u0_u0_u4_n85 ) );
  NOR2_X1 u0_u0_u4_U76 (.A2( u0_u0_X_25 ) , .A1( u0_u0_X_26 ) , .ZN( u0_u0_u4_n89 ) );
  AND2_X1 u0_u0_u4_U77 (.A2( u0_u0_X_25 ) , .A1( u0_u0_X_26 ) , .ZN( u0_u0_u4_n83 ) );
  AND2_X1 u0_u0_u4_U78 (.A1( u0_u0_X_30 ) , .A2( u0_u0_u4_n11 ) , .ZN( u0_u0_u4_n88 ) );
  AND2_X1 u0_u0_u4_U79 (.A1( u0_u0_X_26 ) , .A2( u0_u0_u4_n10 ) , .ZN( u0_u0_u4_n86 ) );
  AOI21_X1 u0_u0_u4_U8 (.B1( u0_u0_u4_n28 ) , .B2( u0_u0_u4_n3 ) , .A( u0_u0_u4_n34 ) , .ZN( u0_u0_u4_n78 ) );
  AND2_X1 u0_u0_u4_U80 (.A1( u0_u0_X_27 ) , .A2( u0_u0_X_30 ) , .ZN( u0_u0_u4_n84 ) );
  INV_X1 u0_u0_u4_U81 (.A( u0_u0_X_28 ) , .ZN( u0_u0_u4_n18 ) );
  INV_X1 u0_u0_u4_U82 (.A( u0_u0_X_29 ) , .ZN( u0_u0_u4_n19 ) );
  INV_X1 u0_u0_u4_U83 (.A( u0_u0_X_25 ) , .ZN( u0_u0_u4_n10 ) );
  INV_X1 u0_u0_u4_U84 (.A( u0_u0_X_27 ) , .ZN( u0_u0_u4_n11 ) );
  NAND4_X1 u0_u0_u4_U85 (.ZN( u0_out0_25 ) , .A1( u0_u0_u4_n45 ) , .A2( u0_u0_u4_n46 ) , .A3( u0_u0_u4_n47 ) , .A4( u0_u0_u4_n48 ) );
  OAI21_X1 u0_u0_u4_U86 (.ZN( u0_u0_u4_n45 ) , .B1( u0_u0_u4_n57 ) , .B2( u0_u0_u4_n58 ) , .A( u0_u0_u4_n59 ) );
  OAI21_X1 u0_u0_u4_U87 (.A( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n4 ) , .ZN( u0_u0_u4_n46 ) , .B2( u0_u0_u4_n56 ) );
  NAND4_X1 u0_u0_u4_U88 (.ZN( u0_out0_14 ) , .A1( u0_u0_u4_n60 ) , .A2( u0_u0_u4_n61 ) , .A3( u0_u0_u4_n62 ) , .A4( u0_u0_u4_n63 ) );
  AOI22_X1 u0_u0_u4_U89 (.A2( u0_u0_u4_n12 ) , .B1( u0_u0_u4_n35 ) , .A1( u0_u0_u4_n58 ) , .ZN( u0_u0_u4_n61 ) , .B2( u0_u0_u4_n70 ) );
  AOI211_X1 u0_u0_u4_U9 (.ZN( u0_u0_u4_n48 ) , .C2( u0_u0_u4_n49 ) , .C1( u0_u0_u4_n5 ) , .A( u0_u0_u4_n50 ) , .B( u0_u0_u4_n51 ) );
  AOI22_X1 u0_u0_u4_U90 (.B1( u0_u0_u4_n49 ) , .A2( u0_u0_u4_n55 ) , .B2( u0_u0_u4_n56 ) , .ZN( u0_u0_u4_n62 ) , .A1( u0_u0_u4_n9 ) );
  NAND4_X1 u0_u0_u4_U91 (.ZN( u0_out0_8 ) , .A1( u0_u0_u4_n1 ) , .A2( u0_u0_u4_n75 ) , .A3( u0_u0_u4_n76 ) , .A4( u0_u0_u4_n77 ) );
  NAND2_X1 u0_u0_u4_U92 (.A1( u0_u0_u4_n37 ) , .A2( u0_u0_u4_n57 ) , .ZN( u0_u0_u4_n75 ) );
  AOI22_X1 u0_u0_u4_U93 (.A1( u0_u0_u4_n35 ) , .B2( u0_u0_u4_n55 ) , .ZN( u0_u0_u4_n76 ) , .B1( u0_u0_u4_n9 ) , .A2( u0_u0_u4_n90 ) );
  AOI22_X1 u0_u0_u4_U94 (.ZN( u0_u0_u4_n20 ) , .A1( u0_u0_u4_n35 ) , .A2( u0_u0_u4_n36 ) , .B1( u0_u0_u4_n37 ) , .B2( u0_u0_u4_n38 ) );
  NOR4_X1 u0_u0_u4_U95 (.ZN( u0_u0_u4_n21 ) , .A1( u0_u0_u4_n22 ) , .A2( u0_u0_u4_n23 ) , .A3( u0_u0_u4_n24 ) , .A4( u0_u0_u4_n25 ) );
  NAND3_X1 u0_u0_u4_U96 (.ZN( u0_out0_3 ) , .A2( u0_u0_u4_n1 ) , .A1( u0_u0_u4_n20 ) , .A3( u0_u0_u4_n21 ) );
  NAND3_X1 u0_u0_u4_U97 (.ZN( u0_u0_u4_n38 ) , .A1( u0_u0_u4_n39 ) , .A2( u0_u0_u4_n40 ) , .A3( u0_u0_u4_n41 ) );
  NAND3_X1 u0_u0_u4_U98 (.ZN( u0_u0_u4_n36 ) , .A1( u0_u0_u4_n42 ) , .A2( u0_u0_u4_n43 ) , .A3( u0_u0_u4_n44 ) );
  NAND3_X1 u0_u0_u4_U99 (.A1( u0_u0_u4_n33 ) , .A2( u0_u0_u4_n43 ) , .ZN( u0_u0_u4_n65 ) , .A3( u0_u0_u4_n66 ) );
  INV_X1 u0_u0_u5_U10 (.ZN( u0_u0_u5_n20 ) , .A( u0_u0_u5_n76 ) );
  AOI222_X1 u0_u0_u5_U100 (.A2( u0_u0_u5_n18 ) , .C2( u0_u0_u5_n19 ) , .B2( u0_u0_u5_n23 ) , .C1( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n66 ) , .ZN( u0_u0_u5_n84 ) , .B1( u0_u0_u5_n98 ) );
  NAND4_X1 u0_u0_u5_U101 (.ZN( u0_out0_29 ) , .A1( u0_u0_u5_n1 ) , .A2( u0_u0_u5_n29 ) , .A3( u0_u0_u5_n67 ) , .A4( u0_u0_u5_n68 ) );
  AOI221_X1 u0_u0_u5_U102 (.C1( u0_u0_u5_n13 ) , .B1( u0_u0_u5_n21 ) , .B2( u0_u0_u5_n38 ) , .C2( u0_u0_u5_n65 ) , .ZN( u0_u0_u5_n68 ) , .A( u0_u0_u5_n69 ) );
  AOI222_X1 u0_u0_u5_U103 (.B2( u0_u0_u5_n18 ) , .C2( u0_u0_u5_n22 ) , .C1( u0_u0_u5_n3 ) , .B1( u0_u0_u5_n50 ) , .A2( u0_u0_u5_n51 ) , .ZN( u0_u0_u5_n67 ) , .A1( u0_u0_u5_n9 ) );
  NAND3_X1 u0_u0_u5_U104 (.A1( u0_u0_u5_n36 ) , .A3( u0_u0_u5_n39 ) , .A2( u0_u0_u5_n43 ) , .ZN( u0_u0_u5_n98 ) );
  NOR2_X1 u0_u0_u5_U11 (.A1( u0_u0_u5_n20 ) , .A2( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n37 ) );
  INV_X1 u0_u0_u5_U12 (.ZN( u0_u0_u5_n23 ) , .A( u0_u0_u5_n47 ) );
  AOI21_X1 u0_u0_u5_U13 (.ZN( u0_u0_u5_n35 ) , .B2( u0_u0_u5_n36 ) , .A( u0_u0_u5_n37 ) , .B1( u0_u0_u5_n5 ) );
  INV_X1 u0_u0_u5_U14 (.A( u0_u0_u5_n38 ) , .ZN( u0_u0_u5_n5 ) );
  AOI21_X1 u0_u0_u5_U15 (.ZN( u0_u0_u5_n34 ) , .B1( u0_u0_u5_n39 ) , .B2( u0_u0_u5_n40 ) , .A( u0_u0_u5_n41 ) );
  AOI21_X1 u0_u0_u5_U16 (.A( u0_u0_u5_n47 ) , .ZN( u0_u0_u5_n56 ) , .B1( u0_u0_u5_n57 ) , .B2( u0_u0_u5_n58 ) );
  OAI21_X1 u0_u0_u5_U17 (.ZN( u0_u0_u5_n55 ) , .B1( u0_u0_u5_n62 ) , .B2( u0_u0_u5_n63 ) , .A( u0_u0_u5_n64 ) );
  OAI21_X1 u0_u0_u5_U18 (.A( u0_u0_u5_n24 ) , .B2( u0_u0_u5_n50 ) , .ZN( u0_u0_u5_n64 ) , .B1( u0_u0_u5_n9 ) );
  NAND2_X1 u0_u0_u5_U19 (.ZN( u0_u0_u5_n60 ) , .A1( u0_u0_u5_n74 ) , .A2( u0_u0_u5_n78 ) );
  INV_X1 u0_u0_u5_U20 (.ZN( u0_u0_u5_n3 ) , .A( u0_u0_u5_n42 ) );
  NAND2_X1 u0_u0_u5_U21 (.A2( u0_u0_u5_n25 ) , .ZN( u0_u0_u5_n65 ) , .A1( u0_u0_u5_n76 ) );
  NAND2_X1 u0_u0_u5_U22 (.A1( u0_u0_u5_n43 ) , .ZN( u0_u0_u5_n61 ) , .A2( u0_u0_u5_n75 ) );
  NAND2_X1 u0_u0_u5_U23 (.ZN( u0_u0_u5_n38 ) , .A1( u0_u0_u5_n77 ) , .A2( u0_u0_u5_n78 ) );
  INV_X1 u0_u0_u5_U24 (.ZN( u0_u0_u5_n22 ) , .A( u0_u0_u5_n41 ) );
  INV_X1 u0_u0_u5_U25 (.A( u0_u0_u5_n39 ) , .ZN( u0_u0_u5_n9 ) );
  INV_X1 u0_u0_u5_U26 (.ZN( u0_u0_u5_n18 ) , .A( u0_u0_u5_n45 ) );
  INV_X1 u0_u0_u5_U27 (.ZN( u0_u0_u5_n15 ) , .A( u0_u0_u5_n57 ) );
  INV_X1 u0_u0_u5_U28 (.ZN( u0_u0_u5_n14 ) , .A( u0_u0_u5_n46 ) );
  INV_X1 u0_u0_u5_U29 (.ZN( u0_u0_u5_n12 ) , .A( u0_u0_u5_n74 ) );
  NOR2_X1 u0_u0_u5_U3 (.A1( u0_u0_u5_n14 ) , .ZN( u0_u0_u5_n63 ) , .A2( u0_u0_u5_n7 ) );
  INV_X1 u0_u0_u5_U30 (.ZN( u0_u0_u5_n13 ) , .A( u0_u0_u5_n36 ) );
  INV_X1 u0_u0_u5_U31 (.A( u0_u0_u5_n58 ) , .ZN( u0_u0_u5_n8 ) );
  INV_X1 u0_u0_u5_U32 (.A( u0_u0_u5_n40 ) , .ZN( u0_u0_u5_n7 ) );
  INV_X1 u0_u0_u5_U33 (.ZN( u0_u0_u5_n4 ) , .A( u0_u0_u5_n77 ) );
  NAND2_X1 u0_u0_u5_U34 (.A2( u0_u0_u5_n42 ) , .A1( u0_u0_u5_n57 ) , .ZN( u0_u0_u5_n86 ) );
  NOR2_X1 u0_u0_u5_U35 (.A2( u0_u0_u5_n17 ) , .A1( u0_u0_u5_n27 ) , .ZN( u0_u0_u5_n97 ) );
  INV_X1 u0_u0_u5_U36 (.ZN( u0_u0_u5_n1 ) , .A( u0_u0_u5_n80 ) );
  OAI221_X1 u0_u0_u5_U37 (.B1( u0_u0_u5_n25 ) , .C2( u0_u0_u5_n39 ) , .C1( u0_u0_u5_n44 ) , .B2( u0_u0_u5_n78 ) , .ZN( u0_u0_u5_n80 ) , .A( u0_u0_u5_n81 ) );
  AOI222_X1 u0_u0_u5_U38 (.B1( u0_u0_u5_n10 ) , .C2( u0_u0_u5_n20 ) , .A2( u0_u0_u5_n23 ) , .A1( u0_u0_u5_n4 ) , .C1( u0_u0_u5_n49 ) , .B2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n81 ) );
  INV_X1 u0_u0_u5_U39 (.ZN( u0_u0_u5_n10 ) , .A( u0_u0_u5_n82 ) );
  INV_X1 u0_u0_u5_U4 (.A( u0_u0_u5_n59 ) , .ZN( u0_u0_u5_n6 ) );
  AOI22_X1 u0_u0_u5_U40 (.A1( u0_u0_u5_n12 ) , .B1( u0_u0_u5_n23 ) , .ZN( u0_u0_u5_n28 ) , .A2( u0_u0_u5_n51 ) , .B2( u0_u0_u5_n66 ) );
  NOR2_X1 u0_u0_u5_U41 (.A2( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n47 ) , .A1( u0_u0_u5_n51 ) );
  AOI21_X1 u0_u0_u5_U42 (.B1( u0_u0_u5_n11 ) , .ZN( u0_u0_u5_n29 ) , .B2( u0_u0_u5_n52 ) , .A( u0_u0_u5_n79 ) );
  INV_X1 u0_u0_u5_U43 (.ZN( u0_u0_u5_n11 ) , .A( u0_u0_u5_n75 ) );
  NOR2_X1 u0_u0_u5_U44 (.A2( u0_u0_u5_n21 ) , .ZN( u0_u0_u5_n45 ) , .A1( u0_u0_u5_n51 ) );
  NOR2_X1 u0_u0_u5_U45 (.A2( u0_u0_u5_n44 ) , .ZN( u0_u0_u5_n79 ) , .A1( u0_u0_u5_n82 ) );
  NOR2_X1 u0_u0_u5_U46 (.A1( u0_u0_u5_n23 ) , .ZN( u0_u0_u5_n41 ) , .A2( u0_u0_u5_n52 ) );
  NOR2_X1 u0_u0_u5_U47 (.A1( u0_u0_u5_n21 ) , .A2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n76 ) );
  AOI22_X1 u0_u0_u5_U48 (.B2( u0_u0_u5_n22 ) , .B1( u0_u0_u5_n4 ) , .A1( u0_u0_u5_n52 ) , .A2( u0_u0_u5_n60 ) , .ZN( u0_u0_u5_n83 ) );
  OAI211_X1 u0_u0_u5_U49 (.ZN( u0_u0_u5_n69 ) , .C1( u0_u0_u5_n70 ) , .C2( u0_u0_u5_n71 ) , .A( u0_u0_u5_n72 ) , .B( u0_u0_u5_n73 ) );
  OAI21_X1 u0_u0_u5_U5 (.A( u0_u0_u5_n20 ) , .ZN( u0_u0_u5_n59 ) , .B1( u0_u0_u5_n60 ) , .B2( u0_u0_u5_n61 ) );
  NOR3_X1 u0_u0_u5_U50 (.A2( u0_u0_u5_n15 ) , .A3( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n61 ) , .ZN( u0_u0_u5_n70 ) );
  OAI21_X1 u0_u0_u5_U51 (.B2( u0_u0_u5_n14 ) , .A( u0_u0_u5_n20 ) , .ZN( u0_u0_u5_n73 ) , .B1( u0_u0_u5_n8 ) );
  OAI21_X1 u0_u0_u5_U52 (.B2( u0_u0_u5_n12 ) , .A( u0_u0_u5_n23 ) , .B1( u0_u0_u5_n7 ) , .ZN( u0_u0_u5_n72 ) );
  AOI21_X1 u0_u0_u5_U53 (.ZN( u0_u0_u5_n33 ) , .B1( u0_u0_u5_n42 ) , .B2( u0_u0_u5_n43 ) , .A( u0_u0_u5_n44 ) );
  AOI21_X1 u0_u0_u5_U54 (.A( u0_u0_u5_n44 ) , .B2( u0_u0_u5_n58 ) , .B1( u0_u0_u5_n75 ) , .ZN( u0_u0_u5_n87 ) );
  INV_X1 u0_u0_u5_U55 (.ZN( u0_u0_u5_n21 ) , .A( u0_u0_u5_n44 ) );
  INV_X1 u0_u0_u5_U56 (.ZN( u0_u0_u5_n24 ) , .A( u0_u0_u5_n71 ) );
  AND2_X1 u0_u0_u5_U57 (.ZN( u0_u0_u5_n50 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n93 ) );
  AND2_X1 u0_u0_u5_U58 (.ZN( u0_u0_u5_n49 ) , .A1( u0_u0_u5_n89 ) , .A2( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U59 (.ZN( u0_u0_u5_n39 ) , .A2( u0_u0_u5_n91 ) , .A1( u0_u0_u5_n92 ) );
  INV_X1 u0_u0_u5_U6 (.ZN( u0_u0_u5_n19 ) , .A( u0_u0_u5_n62 ) );
  NAND2_X1 u0_u0_u5_U60 (.ZN( u0_u0_u5_n58 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n89 ) );
  NAND2_X1 u0_u0_u5_U61 (.ZN( u0_u0_u5_n78 ) , .A2( u0_u0_u5_n89 ) , .A1( u0_u0_u5_n91 ) );
  NAND2_X1 u0_u0_u5_U62 (.ZN( u0_u0_u5_n57 ) , .A1( u0_u0_u5_n92 ) , .A2( u0_u0_u5_n94 ) );
  NAND2_X1 u0_u0_u5_U63 (.ZN( u0_u0_u5_n42 ) , .A1( u0_u0_u5_n92 ) , .A2( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U64 (.ZN( u0_u0_u5_n75 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n91 ) );
  NAND2_X1 u0_u0_u5_U65 (.ZN( u0_u0_u5_n82 ) , .A1( u0_u0_u5_n91 ) , .A2( u0_u0_u5_n97 ) );
  NAND2_X1 u0_u0_u5_U66 (.ZN( u0_u0_u5_n36 ) , .A1( u0_u0_u5_n94 ) , .A2( u0_u0_u5_n97 ) );
  NAND2_X1 u0_u0_u5_U67 (.ZN( u0_u0_u5_n43 ) , .A2( u0_u0_u5_n88 ) , .A1( u0_u0_u5_n92 ) );
  INV_X1 u0_u0_u5_U68 (.ZN( u0_u0_u5_n25 ) , .A( u0_u0_u5_n51 ) );
  NAND2_X1 u0_u0_u5_U69 (.ZN( u0_u0_u5_n74 ) , .A2( u0_u0_u5_n89 ) , .A1( u0_u0_u5_n94 ) );
  OAI22_X1 u0_u0_u5_U7 (.ZN( u0_u0_u5_n32 ) , .A1( u0_u0_u5_n45 ) , .A2( u0_u0_u5_n46 ) , .B1( u0_u0_u5_n47 ) , .B2( u0_u0_u5_n48 ) );
  NAND2_X1 u0_u0_u5_U70 (.ZN( u0_u0_u5_n46 ) , .A1( u0_u0_u5_n90 ) , .A2( u0_u0_u5_n94 ) );
  NAND2_X1 u0_u0_u5_U71 (.ZN( u0_u0_u5_n77 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n90 ) );
  NAND2_X1 u0_u0_u5_U72 (.ZN( u0_u0_u5_n40 ) , .A1( u0_u0_u5_n88 ) , .A2( u0_u0_u5_n97 ) );
  AND2_X1 u0_u0_u5_U73 (.ZN( u0_u0_u5_n66 ) , .A1( u0_u0_u5_n93 ) , .A2( u0_u0_u5_n97 ) );
  INV_X1 u0_u0_u5_U74 (.ZN( u0_u0_u5_n2 ) , .A( u0_u0_u5_n95 ) );
  OAI221_X1 u0_u0_u5_U75 (.B2( u0_u0_u5_n37 ) , .B1( u0_u0_u5_n63 ) , .C1( u0_u0_u5_n71 ) , .C2( u0_u0_u5_n82 ) , .ZN( u0_u0_u5_n95 ) , .A( u0_u0_u5_n96 ) );
  OAI21_X1 u0_u0_u5_U76 (.B2( u0_u0_u5_n50 ) , .A( u0_u0_u5_n51 ) , .B1( u0_u0_u5_n60 ) , .ZN( u0_u0_u5_n96 ) );
  NOR2_X1 u0_u0_u5_U77 (.A2( u0_u0_X_34 ) , .A1( u0_u0_X_35 ) , .ZN( u0_u0_u5_n52 ) );
  NOR2_X1 u0_u0_u5_U78 (.A2( u0_u0_X_34 ) , .A1( u0_u0_u5_n26 ) , .ZN( u0_u0_u5_n51 ) );
  NOR2_X1 u0_u0_u5_U79 (.A2( u0_u0_X_31 ) , .A1( u0_u0_X_32 ) , .ZN( u0_u0_u5_n94 ) );
  NOR3_X1 u0_u0_u5_U8 (.A3( u0_u0_u5_n3 ) , .ZN( u0_u0_u5_n48 ) , .A1( u0_u0_u5_n49 ) , .A2( u0_u0_u5_n50 ) );
  NOR2_X1 u0_u0_u5_U80 (.A2( u0_u0_X_36 ) , .A1( u0_u0_u5_n17 ) , .ZN( u0_u0_u5_n92 ) );
  NOR2_X1 u0_u0_u5_U81 (.A2( u0_u0_X_33 ) , .A1( u0_u0_u5_n27 ) , .ZN( u0_u0_u5_n89 ) );
  NOR2_X1 u0_u0_u5_U82 (.A2( u0_u0_X_33 ) , .A1( u0_u0_X_36 ) , .ZN( u0_u0_u5_n90 ) );
  NOR2_X1 u0_u0_u5_U83 (.A2( u0_u0_X_31 ) , .A1( u0_u0_u5_n16 ) , .ZN( u0_u0_u5_n93 ) );
  NAND2_X1 u0_u0_u5_U84 (.A2( u0_u0_X_34 ) , .A1( u0_u0_X_35 ) , .ZN( u0_u0_u5_n44 ) );
  NAND2_X1 u0_u0_u5_U85 (.A1( u0_u0_X_34 ) , .A2( u0_u0_u5_n26 ) , .ZN( u0_u0_u5_n71 ) );
  AND2_X1 u0_u0_u5_U86 (.A1( u0_u0_X_31 ) , .A2( u0_u0_X_32 ) , .ZN( u0_u0_u5_n91 ) );
  AND2_X1 u0_u0_u5_U87 (.A1( u0_u0_X_31 ) , .A2( u0_u0_u5_n16 ) , .ZN( u0_u0_u5_n88 ) );
  INV_X1 u0_u0_u5_U88 (.A( u0_u0_X_33 ) , .ZN( u0_u0_u5_n17 ) );
  INV_X1 u0_u0_u5_U89 (.A( u0_u0_X_35 ) , .ZN( u0_u0_u5_n26 ) );
  NOR2_X1 u0_u0_u5_U9 (.A2( u0_u0_u5_n21 ) , .A1( u0_u0_u5_n24 ) , .ZN( u0_u0_u5_n62 ) );
  INV_X1 u0_u0_u5_U90 (.A( u0_u0_X_36 ) , .ZN( u0_u0_u5_n27 ) );
  INV_X1 u0_u0_u5_U91 (.A( u0_u0_X_32 ) , .ZN( u0_u0_u5_n16 ) );
  NAND4_X1 u0_u0_u5_U92 (.ZN( u0_out0_19 ) , .A1( u0_u0_u5_n28 ) , .A2( u0_u0_u5_n29 ) , .A3( u0_u0_u5_n30 ) , .A4( u0_u0_u5_n31 ) );
  AOI22_X1 u0_u0_u5_U93 (.B1( u0_u0_u5_n15 ) , .ZN( u0_u0_u5_n30 ) , .A2( u0_u0_u5_n51 ) , .B2( u0_u0_u5_n52 ) , .A1( u0_u0_u5_n8 ) );
  NOR4_X1 u0_u0_u5_U94 (.ZN( u0_u0_u5_n31 ) , .A1( u0_u0_u5_n32 ) , .A2( u0_u0_u5_n33 ) , .A3( u0_u0_u5_n34 ) , .A4( u0_u0_u5_n35 ) );
  NAND4_X1 u0_u0_u5_U95 (.ZN( u0_out0_11 ) , .A1( u0_u0_u5_n1 ) , .A2( u0_u0_u5_n28 ) , .A3( u0_u0_u5_n53 ) , .A4( u0_u0_u5_n54 ) );
  AOI22_X1 u0_u0_u5_U96 (.B1( u0_u0_u5_n13 ) , .A1( u0_u0_u5_n3 ) , .B2( u0_u0_u5_n52 ) , .ZN( u0_u0_u5_n53 ) , .A2( u0_u0_u5_n65 ) );
  NOR3_X1 u0_u0_u5_U97 (.ZN( u0_u0_u5_n54 ) , .A1( u0_u0_u5_n55 ) , .A3( u0_u0_u5_n56 ) , .A2( u0_u0_u5_n6 ) );
  NAND4_X1 u0_u0_u5_U98 (.ZN( u0_out0_4 ) , .A3( u0_u0_u5_n2 ) , .A1( u0_u0_u5_n83 ) , .A2( u0_u0_u5_n84 ) , .A4( u0_u0_u5_n85 ) );
  AOI211_X1 u0_u0_u5_U99 (.C2( u0_u0_u5_n20 ) , .B( u0_u0_u5_n79 ) , .ZN( u0_u0_u5_n85 ) , .C1( u0_u0_u5_n86 ) , .A( u0_u0_u5_n87 ) );
  AOI22_X1 u0_u0_u6_U10 (.B2( u0_u0_u6_n14 ) , .A2( u0_u0_u6_n24 ) , .B1( u0_u0_u6_n5 ) , .A1( u0_u0_u6_n8 ) , .ZN( u0_u0_u6_n86 ) );
  AOI21_X1 u0_u0_u6_U11 (.A( u0_u0_u6_n17 ) , .B2( u0_u0_u6_n43 ) , .B1( u0_u0_u6_n68 ) , .ZN( u0_u0_u6_n87 ) );
  AOI21_X1 u0_u0_u6_U12 (.A( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n26 ) , .B1( u0_u0_u6_n27 ) , .B2( u0_u0_u6_n28 ) );
  AOI21_X1 u0_u0_u6_U13 (.B1( u0_u0_u6_n11 ) , .B2( u0_u0_u6_n16 ) , .A( u0_u0_u6_n33 ) , .ZN( u0_u0_u6_n69 ) );
  INV_X1 u0_u0_u6_U14 (.ZN( u0_u0_u6_n14 ) , .A( u0_u0_u6_n20 ) );
  INV_X1 u0_u0_u6_U15 (.ZN( u0_u0_u6_n11 ) , .A( u0_u0_u6_n47 ) );
  NAND2_X1 u0_u0_u6_U16 (.A2( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n53 ) , .ZN( u0_u0_u6_n65 ) );
  NAND2_X1 u0_u0_u6_U17 (.A1( u0_u0_u6_n27 ) , .A2( u0_u0_u6_n29 ) , .ZN( u0_u0_u6_n51 ) );
  INV_X1 u0_u0_u6_U18 (.ZN( u0_u0_u6_n4 ) , .A( u0_u0_u6_n43 ) );
  AND2_X1 u0_u0_u6_U19 (.A2( u0_u0_u6_n28 ) , .ZN( u0_u0_u6_n45 ) , .A1( u0_u0_u6_n75 ) );
  INV_X1 u0_u0_u6_U20 (.ZN( u0_u0_u6_n2 ) , .A( u0_u0_u6_n48 ) );
  INV_X1 u0_u0_u6_U21 (.A( u0_u0_u6_n54 ) , .ZN( u0_u0_u6_n8 ) );
  INV_X1 u0_u0_u6_U22 (.ZN( u0_u0_u6_n6 ) , .A( u0_u0_u6_n75 ) );
  INV_X1 u0_u0_u6_U23 (.ZN( u0_u0_u6_n5 ) , .A( u0_u0_u6_n52 ) );
  INV_X1 u0_u0_u6_U24 (.A( u0_u0_u6_n62 ) , .ZN( u0_u0_u6_n7 ) );
  AND2_X1 u0_u0_u6_U25 (.ZN( u0_u0_u6_n42 ) , .A2( u0_u0_u6_n56 ) , .A1( u0_u0_u6_n68 ) );
  AND2_X1 u0_u0_u6_U26 (.ZN( u0_u0_u6_n44 ) , .A1( u0_u0_u6_n53 ) , .A2( u0_u0_u6_n54 ) );
  AND3_X1 u0_u0_u6_U27 (.A3( u0_u0_u6_n30 ) , .A1( u0_u0_u6_n43 ) , .A2( u0_u0_u6_n48 ) , .ZN( u0_u0_u6_n55 ) );
  INV_X1 u0_u0_u6_U28 (.ZN( u0_u0_u6_n12 ) , .A( u0_u0_u6_n29 ) );
  AOI222_X1 u0_u0_u6_U29 (.C2( u0_u0_u6_n16 ) , .B2( u0_u0_u6_n24 ) , .A2( u0_u0_u6_n49 ) , .A1( u0_u0_u6_n57 ) , .B1( u0_u0_u6_n6 ) , .ZN( u0_u0_u6_n61 ) , .C1( u0_u0_u6_n7 ) );
  INV_X1 u0_u0_u6_U3 (.A( u0_u0_u6_n65 ) , .ZN( u0_u0_u6_n9 ) );
  NOR2_X1 u0_u0_u6_U30 (.A2( u0_u0_u6_n10 ) , .A1( u0_u0_u6_n13 ) , .ZN( u0_u0_u6_n77 ) );
  AOI211_X1 u0_u0_u6_U31 (.C2( u0_u0_u6_n24 ) , .ZN( u0_u0_u6_n38 ) , .C1( u0_u0_u6_n39 ) , .A( u0_u0_u6_n40 ) , .B( u0_u0_u6_n41 ) );
  AOI21_X1 u0_u0_u6_U32 (.A( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n41 ) , .B1( u0_u0_u6_n42 ) , .B2( u0_u0_u6_n43 ) );
  NAND4_X1 u0_u0_u6_U33 (.ZN( u0_u0_u6_n39 ) , .A1( u0_u0_u6_n45 ) , .A2( u0_u0_u6_n46 ) , .A3( u0_u0_u6_n47 ) , .A4( u0_u0_u6_n48 ) );
  AOI21_X1 u0_u0_u6_U34 (.B2( u0_u0_u6_n29 ) , .A( u0_u0_u6_n31 ) , .ZN( u0_u0_u6_n40 ) , .B1( u0_u0_u6_n44 ) );
  NAND2_X1 u0_u0_u6_U35 (.A2( u0_u0_u6_n17 ) , .ZN( u0_u0_u6_n24 ) , .A1( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U36 (.ZN( u0_u0_u6_n43 ) , .A2( u0_u0_u6_n78 ) , .A1( u0_u0_u6_n84 ) );
  AOI22_X1 u0_u0_u6_U37 (.A2( u0_u0_u6_n14 ) , .ZN( u0_u0_u6_n60 ) , .A1( u0_u0_u6_n63 ) , .B1( u0_u0_u6_n64 ) , .B2( u0_u0_u6_n65 ) );
  NAND4_X1 u0_u0_u6_U38 (.A2( u0_u0_u6_n28 ) , .A4( u0_u0_u6_n43 ) , .ZN( u0_u0_u6_n63 ) , .A3( u0_u0_u6_n66 ) , .A1( u0_u0_u6_n9 ) );
  NOR2_X1 u0_u0_u6_U39 (.A2( u0_u0_u6_n2 ) , .A1( u0_u0_u6_n5 ) , .ZN( u0_u0_u6_n66 ) );
  INV_X1 u0_u0_u6_U4 (.ZN( u0_u0_u6_n1 ) , .A( u0_u0_u6_n33 ) );
  NOR2_X1 u0_u0_u6_U40 (.A1( u0_u0_u6_n15 ) , .ZN( u0_u0_u6_n20 ) , .A2( u0_u0_u6_n49 ) );
  NAND2_X1 u0_u0_u6_U41 (.ZN( u0_u0_u6_n29 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n81 ) );
  AOI21_X1 u0_u0_u6_U42 (.ZN( u0_u0_u6_n25 ) , .B1( u0_u0_u6_n29 ) , .B2( u0_u0_u6_n30 ) , .A( u0_u0_u6_n31 ) );
  INV_X1 u0_u0_u6_U43 (.ZN( u0_u0_u6_n17 ) , .A( u0_u0_u6_n64 ) );
  NAND2_X1 u0_u0_u6_U44 (.ZN( u0_u0_u6_n48 ) , .A2( u0_u0_u6_n83 ) , .A1( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U45 (.ZN( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n79 ) , .A2( u0_u0_u6_n80 ) );
  INV_X1 u0_u0_u6_U46 (.ZN( u0_u0_u6_n16 ) , .A( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U47 (.ZN( u0_u0_u6_n30 ) , .A1( u0_u0_u6_n77 ) , .A2( u0_u0_u6_n78 ) );
  NAND2_X1 u0_u0_u6_U48 (.ZN( u0_u0_u6_n27 ) , .A1( u0_u0_u6_n81 ) , .A2( u0_u0_u6_n83 ) );
  NAND2_X1 u0_u0_u6_U49 (.A1( u0_u0_u6_n31 ) , .A2( u0_u0_u6_n36 ) , .ZN( u0_u0_u6_n67 ) );
  NAND2_X1 u0_u0_u6_U5 (.ZN( u0_u0_u6_n23 ) , .A2( u0_u0_u6_n32 ) , .A1( u0_u0_u6_n9 ) );
  NAND2_X1 u0_u0_u6_U50 (.ZN( u0_u0_u6_n54 ) , .A1( u0_u0_u6_n78 ) , .A2( u0_u0_u6_n80 ) );
  NAND2_X1 u0_u0_u6_U51 (.ZN( u0_u0_u6_n68 ) , .A1( u0_u0_u6_n80 ) , .A2( u0_u0_u6_n83 ) );
  AND2_X1 u0_u0_u6_U52 (.ZN( u0_u0_u6_n57 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U53 (.ZN( u0_u0_u6_n28 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n77 ) );
  NAND2_X1 u0_u0_u6_U54 (.ZN( u0_u0_u6_n47 ) , .A2( u0_u0_u6_n79 ) , .A1( u0_u0_u6_n81 ) );
  NAND2_X1 u0_u0_u6_U55 (.ZN( u0_u0_u6_n56 ) , .A1( u0_u0_u6_n76 ) , .A2( u0_u0_u6_n80 ) );
  NAND2_X1 u0_u0_u6_U56 (.ZN( u0_u0_u6_n52 ) , .A1( u0_u0_u6_n79 ) , .A2( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U57 (.ZN( u0_u0_u6_n75 ) , .A1( u0_u0_u6_n77 ) , .A2( u0_u0_u6_n83 ) );
  NAND2_X1 u0_u0_u6_U58 (.ZN( u0_u0_u6_n53 ) , .A2( u0_u0_u6_n78 ) , .A1( u0_u0_u6_n81 ) );
  INV_X1 u0_u0_u6_U59 (.ZN( u0_u0_u6_n15 ) , .A( u0_u0_u6_n36 ) );
  AOI22_X1 u0_u0_u6_U6 (.A2( u0_u0_u6_n14 ) , .B1( u0_u0_u6_n15 ) , .ZN( u0_u0_u6_n72 ) , .A1( u0_u0_u6_n73 ) , .B2( u0_u0_u6_n74 ) );
  NAND2_X1 u0_u0_u6_U60 (.ZN( u0_u0_u6_n62 ) , .A2( u0_u0_u6_n77 ) , .A1( u0_u0_u6_n79 ) );
  NOR2_X1 u0_u0_u6_U61 (.A2( u0_u0_X_40 ) , .A1( u0_u0_X_41 ) , .ZN( u0_u0_u6_n49 ) );
  NOR2_X1 u0_u0_u6_U62 (.A2( u0_u0_X_39 ) , .A1( u0_u0_X_42 ) , .ZN( u0_u0_u6_n83 ) );
  NOR2_X1 u0_u0_u6_U63 (.A2( u0_u0_X_39 ) , .A1( u0_u0_u6_n19 ) , .ZN( u0_u0_u6_n78 ) );
  NOR2_X1 u0_u0_u6_U64 (.A2( u0_u0_X_38 ) , .A1( u0_u0_u6_n10 ) , .ZN( u0_u0_u6_n80 ) );
  NOR2_X1 u0_u0_u6_U65 (.A2( u0_u0_X_41 ) , .A1( u0_u0_u6_n18 ) , .ZN( u0_u0_u6_n64 ) );
  NOR2_X1 u0_u0_u6_U66 (.A2( u0_u0_X_37 ) , .A1( u0_u0_u6_n13 ) , .ZN( u0_u0_u6_n81 ) );
  NOR2_X1 u0_u0_u6_U67 (.A2( u0_u0_X_37 ) , .A1( u0_u0_X_38 ) , .ZN( u0_u0_u6_n84 ) );
  NAND2_X1 u0_u0_u6_U68 (.A1( u0_u0_X_41 ) , .A2( u0_u0_u6_n18 ) , .ZN( u0_u0_u6_n31 ) );
  NAND2_X1 u0_u0_u6_U69 (.A2( u0_u0_X_40 ) , .A1( u0_u0_X_41 ) , .ZN( u0_u0_u6_n36 ) );
  NOR2_X1 u0_u0_u6_U7 (.ZN( u0_u0_u6_n32 ) , .A1( u0_u0_u6_n57 ) , .A2( u0_u0_u6_n7 ) );
  AND2_X1 u0_u0_u6_U70 (.A1( u0_u0_X_39 ) , .A2( u0_u0_u6_n19 ) , .ZN( u0_u0_u6_n79 ) );
  AND2_X1 u0_u0_u6_U71 (.A1( u0_u0_X_39 ) , .A2( u0_u0_X_42 ) , .ZN( u0_u0_u6_n76 ) );
  INV_X1 u0_u0_u6_U72 (.A( u0_u0_X_40 ) , .ZN( u0_u0_u6_n18 ) );
  INV_X1 u0_u0_u6_U73 (.A( u0_u0_X_37 ) , .ZN( u0_u0_u6_n10 ) );
  INV_X1 u0_u0_u6_U74 (.A( u0_u0_X_38 ) , .ZN( u0_u0_u6_n13 ) );
  INV_X1 u0_u0_u6_U75 (.A( u0_u0_X_42 ) , .ZN( u0_u0_u6_n19 ) );
  NAND4_X1 u0_u0_u6_U76 (.ZN( u0_out0_12 ) , .A1( u0_u0_u6_n58 ) , .A2( u0_u0_u6_n59 ) , .A3( u0_u0_u6_n60 ) , .A4( u0_u0_u6_n61 ) );
  OAI22_X1 u0_u0_u6_U77 (.A2( u0_u0_u6_n11 ) , .B1( u0_u0_u6_n49 ) , .ZN( u0_u0_u6_n59 ) , .B2( u0_u0_u6_n64 ) , .A1( u0_u0_u6_n8 ) );
  OAI21_X1 u0_u0_u6_U78 (.B1( u0_u0_u6_n12 ) , .B2( u0_u0_u6_n34 ) , .ZN( u0_u0_u6_n58 ) , .A( u0_u0_u6_n67 ) );
  NAND4_X1 u0_u0_u6_U79 (.ZN( u0_out0_32 ) , .A1( u0_u0_u6_n69 ) , .A2( u0_u0_u6_n70 ) , .A3( u0_u0_u6_n71 ) , .A4( u0_u0_u6_n72 ) );
  OAI21_X1 u0_u0_u6_U8 (.A( u0_u0_u6_n16 ) , .B2( u0_u0_u6_n2 ) , .B1( u0_u0_u6_n6 ) , .ZN( u0_u0_u6_n85 ) );
  AOI22_X1 u0_u0_u6_U80 (.B1( u0_u0_u6_n4 ) , .B2( u0_u0_u6_n49 ) , .A1( u0_u0_u6_n57 ) , .A2( u0_u0_u6_n67 ) , .ZN( u0_u0_u6_n70 ) );
  AOI22_X1 u0_u0_u6_U81 (.B2( u0_u0_u6_n24 ) , .B1( u0_u0_u6_n51 ) , .A1( u0_u0_u6_n64 ) , .ZN( u0_u0_u6_n71 ) , .A2( u0_u0_u6_n82 ) );
  OAI211_X1 u0_u0_u6_U82 (.ZN( u0_out0_7 ) , .A( u0_u0_u6_n1 ) , .C1( u0_u0_u6_n20 ) , .C2( u0_u0_u6_n21 ) , .B( u0_u0_u6_n22 ) );
  NOR3_X1 u0_u0_u6_U83 (.A3( u0_u0_u6_n11 ) , .ZN( u0_u0_u6_n21 ) , .A1( u0_u0_u6_n34 ) , .A2( u0_u0_u6_n4 ) );
  AOI211_X1 u0_u0_u6_U84 (.ZN( u0_u0_u6_n22 ) , .C1( u0_u0_u6_n23 ) , .C2( u0_u0_u6_n24 ) , .A( u0_u0_u6_n25 ) , .B( u0_u0_u6_n26 ) );
  OAI211_X1 u0_u0_u6_U85 (.ZN( u0_out0_22 ) , .C1( u0_u0_u6_n35 ) , .C2( u0_u0_u6_n36 ) , .A( u0_u0_u6_n37 ) , .B( u0_u0_u6_n38 ) );
  AOI22_X1 u0_u0_u6_U86 (.B2( u0_u0_u6_n14 ) , .ZN( u0_u0_u6_n37 ) , .A1( u0_u0_u6_n49 ) , .A2( u0_u0_u6_n50 ) , .B1( u0_u0_u6_n51 ) );
  AND4_X1 u0_u0_u6_U87 (.A2( u0_u0_u6_n32 ) , .ZN( u0_u0_u6_n35 ) , .A4( u0_u0_u6_n46 ) , .A1( u0_u0_u6_n55 ) , .A3( u0_u0_u6_n56 ) );
  NAND3_X1 u0_u0_u6_U88 (.A3( u0_u0_u6_n44 ) , .A1( u0_u0_u6_n45 ) , .ZN( u0_u0_u6_n50 ) , .A2( u0_u0_u6_n52 ) );
  NAND3_X1 u0_u0_u6_U89 (.A2( u0_u0_u6_n27 ) , .A1( u0_u0_u6_n30 ) , .ZN( u0_u0_u6_n34 ) , .A3( u0_u0_u6_n42 ) );
  INV_X1 u0_u0_u6_U9 (.ZN( u0_u0_u6_n3 ) , .A( u0_u0_u6_n87 ) );
  NAND3_X1 u0_u0_u6_U90 (.A1( u0_u0_u6_n48 ) , .A2( u0_u0_u6_n54 ) , .A3( u0_u0_u6_n68 ) , .ZN( u0_u0_u6_n74 ) );
  NAND3_X1 u0_u0_u6_U91 (.A2( u0_u0_u6_n30 ) , .A3( u0_u0_u6_n45 ) , .ZN( u0_u0_u6_n73 ) , .A1( u0_u0_u6_n9 ) );
  NAND3_X1 u0_u0_u6_U92 (.A2( u0_u0_u6_n52 ) , .A1( u0_u0_u6_n56 ) , .A3( u0_u0_u6_n62 ) , .ZN( u0_u0_u6_n82 ) );
  NAND3_X1 u0_u0_u6_U93 (.A2( u0_u0_u6_n3 ) , .ZN( u0_u0_u6_n33 ) , .A1( u0_u0_u6_n85 ) , .A3( u0_u0_u6_n86 ) );
  OAI21_X1 u0_u0_u7_U10 (.B1( u0_u0_u7_n13 ) , .A( u0_u0_u7_n20 ) , .B2( u0_u0_u7_n8 ) , .ZN( u0_u0_u7_n90 ) );
  AOI211_X1 u0_u0_u7_U11 (.B( u0_u0_u7_n1 ) , .C1( u0_u0_u7_n4 ) , .C2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n63 ) , .A( u0_u0_u7_n64 ) );
  OAI22_X1 u0_u0_u7_U12 (.B2( u0_u0_u7_n19 ) , .A1( u0_u0_u7_n44 ) , .A2( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n64 ) , .B1( u0_u0_u7_n66 ) );
  INV_X1 u0_u0_u7_U13 (.ZN( u0_u0_u7_n1 ) , .A( u0_u0_u7_n65 ) );
  NOR3_X1 u0_u0_u7_U14 (.A1( u0_u0_u7_n12 ) , .A2( u0_u0_u7_n13 ) , .A3( u0_u0_u7_n36 ) , .ZN( u0_u0_u7_n66 ) );
  INV_X1 u0_u0_u7_U15 (.A( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n5 ) );
  NOR3_X1 u0_u0_u7_U16 (.A3( u0_u0_u7_n10 ) , .ZN( u0_u0_u7_n45 ) , .A1( u0_u0_u7_n46 ) , .A2( u0_u0_u7_n47 ) );
  NOR2_X1 u0_u0_u7_U17 (.ZN( u0_u0_u7_n28 ) , .A2( u0_u0_u7_n47 ) , .A1( u0_u0_u7_n51 ) );
  AOI21_X1 u0_u0_u7_U18 (.A( u0_u0_u7_n17 ) , .B1( u0_u0_u7_n54 ) , .B2( u0_u0_u7_n69 ) , .ZN( u0_u0_u7_n77 ) );
  AOI21_X1 u0_u0_u7_U19 (.A( u0_u0_u7_n19 ) , .B2( u0_u0_u7_n35 ) , .B1( u0_u0_u7_n48 ) , .ZN( u0_u0_u7_n75 ) );
  AOI21_X1 u0_u0_u7_U20 (.B2( u0_u0_u7_n53 ) , .B1( u0_u0_u7_n6 ) , .ZN( u0_u0_u7_n74 ) , .A( u0_u0_u7_n80 ) );
  INV_X1 u0_u0_u7_U21 (.ZN( u0_u0_u7_n16 ) , .A( u0_u0_u7_n80 ) );
  NOR2_X1 u0_u0_u7_U22 (.A1( u0_u0_u7_n12 ) , .A2( u0_u0_u7_n47 ) , .ZN( u0_u0_u7_n70 ) );
  INV_X1 u0_u0_u7_U23 (.ZN( u0_u0_u7_n10 ) , .A( u0_u0_u7_n43 ) );
  INV_X1 u0_u0_u7_U24 (.ZN( u0_u0_u7_n4 ) , .A( u0_u0_u7_n50 ) );
  INV_X1 u0_u0_u7_U25 (.ZN( u0_u0_u7_n7 ) , .A( u0_u0_u7_n71 ) );
  NAND2_X1 u0_u0_u7_U26 (.ZN( u0_u0_u7_n32 ) , .A2( u0_u0_u7_n49 ) , .A1( u0_u0_u7_n52 ) );
  NAND2_X1 u0_u0_u7_U27 (.ZN( u0_u0_u7_n51 ) , .A2( u0_u0_u7_n57 ) , .A1( u0_u0_u7_n68 ) );
  INV_X1 u0_u0_u7_U28 (.A( u0_u0_u7_n69 ) , .ZN( u0_u0_u7_n8 ) );
  INV_X1 u0_u0_u7_U29 (.ZN( u0_u0_u7_n13 ) , .A( u0_u0_u7_n53 ) );
  OAI21_X1 u0_u0_u7_U3 (.B2( u0_u0_u7_n10 ) , .A( u0_u0_u7_n16 ) , .ZN( u0_u0_u7_n22 ) , .B1( u0_u0_u7_n7 ) );
  INV_X1 u0_u0_u7_U30 (.ZN( u0_u0_u7_n12 ) , .A( u0_u0_u7_n33 ) );
  INV_X1 u0_u0_u7_U31 (.ZN( u0_u0_u7_n2 ) , .A( u0_u0_u7_n54 ) );
  INV_X1 u0_u0_u7_U32 (.A( u0_u0_u7_n28 ) , .ZN( u0_u0_u7_n9 ) );
  NOR2_X1 u0_u0_u7_U33 (.A1( u0_u0_u7_n25 ) , .A2( u0_u0_u7_n31 ) , .ZN( u0_u0_u7_n80 ) );
  AOI211_X1 u0_u0_u7_U34 (.C1( u0_u0_u7_n25 ) , .ZN( u0_u0_u7_n39 ) , .C2( u0_u0_u7_n40 ) , .A( u0_u0_u7_n41 ) , .B( u0_u0_u7_n42 ) );
  NAND4_X1 u0_u0_u7_U35 (.A4( u0_u0_u7_n34 ) , .ZN( u0_u0_u7_n40 ) , .A1( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n53 ) , .A3( u0_u0_u7_n54 ) );
  AOI21_X1 u0_u0_u7_U36 (.B2( u0_u0_u7_n35 ) , .ZN( u0_u0_u7_n42 ) , .B1( u0_u0_u7_n43 ) , .A( u0_u0_u7_n44 ) );
  OAI22_X1 u0_u0_u7_U37 (.A2( u0_u0_u7_n17 ) , .B2( u0_u0_u7_n19 ) , .A1( u0_u0_u7_n28 ) , .ZN( u0_u0_u7_n41 ) , .B1( u0_u0_u7_n45 ) );
  INV_X1 u0_u0_u7_U38 (.ZN( u0_u0_u7_n20 ) , .A( u0_u0_u7_n56 ) );
  AOI21_X1 u0_u0_u7_U39 (.B1( u0_u0_u7_n16 ) , .B2( u0_u0_u7_n4 ) , .ZN( u0_u0_u7_n58 ) , .A( u0_u0_u7_n84 ) );
  INV_X1 u0_u0_u7_U4 (.A( u0_u0_u7_n32 ) , .ZN( u0_u0_u7_n6 ) );
  AOI21_X1 u0_u0_u7_U40 (.A( u0_u0_u7_n56 ) , .B1( u0_u0_u7_n57 ) , .B2( u0_u0_u7_n68 ) , .ZN( u0_u0_u7_n84 ) );
  INV_X1 u0_u0_u7_U41 (.ZN( u0_u0_u7_n19 ) , .A( u0_u0_u7_n29 ) );
  AOI22_X1 u0_u0_u7_U42 (.B2( u0_u0_u7_n16 ) , .A1( u0_u0_u7_n25 ) , .B1( u0_u0_u7_n51 ) , .ZN( u0_u0_u7_n62 ) , .A2( u0_u0_u7_n67 ) );
  NAND2_X1 u0_u0_u7_U43 (.A1( u0_u0_u7_n6 ) , .ZN( u0_u0_u7_n67 ) , .A2( u0_u0_u7_n69 ) );
  NOR2_X1 u0_u0_u7_U44 (.A2( u0_u0_u7_n20 ) , .A1( u0_u0_u7_n31 ) , .ZN( u0_u0_u7_n44 ) );
  AND2_X1 u0_u0_u7_U45 (.ZN( u0_u0_u7_n36 ) , .A1( u0_u0_u7_n82 ) , .A2( u0_u0_u7_n83 ) );
  AOI21_X1 u0_u0_u7_U46 (.B1( u0_u0_u7_n34 ) , .A( u0_u0_u7_n56 ) , .B2( u0_u0_u7_n71 ) , .ZN( u0_u0_u7_n76 ) );
  NAND2_X1 u0_u0_u7_U47 (.ZN( u0_u0_u7_n35 ) , .A2( u0_u0_u7_n83 ) , .A1( u0_u0_u7_n86 ) );
  NAND2_X1 u0_u0_u7_U48 (.ZN( u0_u0_u7_n34 ) , .A2( u0_u0_u7_n78 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U49 (.ZN( u0_u0_u7_n54 ) , .A1( u0_u0_u7_n78 ) , .A2( u0_u0_u7_n82 ) );
  INV_X1 u0_u0_u7_U5 (.A( u0_u0_u7_n27 ) , .ZN( u0_u0_u7_n3 ) );
  NAND2_X1 u0_u0_u7_U50 (.ZN( u0_u0_u7_n48 ) , .A1( u0_u0_u7_n78 ) , .A2( u0_u0_u7_n79 ) );
  OR2_X1 u0_u0_u7_U51 (.A1( u0_u0_u7_n25 ) , .A2( u0_u0_u7_n29 ) , .ZN( u0_u0_u7_n55 ) );
  NAND2_X1 u0_u0_u7_U52 (.ZN( u0_u0_u7_n69 ) , .A1( u0_u0_u7_n82 ) , .A2( u0_u0_u7_n85 ) );
  NAND2_X1 u0_u0_u7_U53 (.ZN( u0_u0_u7_n53 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n83 ) );
  NAND2_X1 u0_u0_u7_U54 (.ZN( u0_u0_u7_n68 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U55 (.ZN( u0_u0_u7_n71 ) , .A2( u0_u0_u7_n85 ) , .A1( u0_u0_u7_n86 ) );
  INV_X1 u0_u0_u7_U56 (.ZN( u0_u0_u7_n17 ) , .A( u0_u0_u7_n31 ) );
  AND2_X1 u0_u0_u7_U57 (.ZN( u0_u0_u7_n47 ) , .A2( u0_u0_u7_n83 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U58 (.ZN( u0_u0_u7_n57 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n85 ) );
  NAND2_X1 u0_u0_u7_U59 (.ZN( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n79 ) , .A1( u0_u0_u7_n81 ) );
  AOI211_X1 u0_u0_u7_U6 (.C2( u0_u0_u7_n10 ) , .C1( u0_u0_u7_n20 ) , .A( u0_u0_u7_n26 ) , .ZN( u0_u0_u7_n65 ) , .B( u0_u0_u7_n87 ) );
  NAND2_X1 u0_u0_u7_U60 (.ZN( u0_u0_u7_n50 ) , .A2( u0_u0_u7_n78 ) , .A1( u0_u0_u7_n86 ) );
  NAND2_X1 u0_u0_u7_U61 (.ZN( u0_u0_u7_n43 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n82 ) );
  NAND2_X1 u0_u0_u7_U62 (.ZN( u0_u0_u7_n49 ) , .A2( u0_u0_u7_n85 ) , .A1( u0_u0_u7_n88 ) );
  NAND2_X1 u0_u0_u7_U63 (.ZN( u0_u0_u7_n33 ) , .A1( u0_u0_u7_n81 ) , .A2( u0_u0_u7_n86 ) );
  NOR2_X1 u0_u0_u7_U64 (.A2( u0_u0_X_47 ) , .A1( u0_u0_u7_n18 ) , .ZN( u0_u0_u7_n31 ) );
  NOR2_X1 u0_u0_u7_U65 (.A2( u0_u0_X_43 ) , .A1( u0_u0_X_44 ) , .ZN( u0_u0_u7_n78 ) );
  NOR2_X1 u0_u0_u7_U66 (.A2( u0_u0_X_48 ) , .A1( u0_u0_u7_n15 ) , .ZN( u0_u0_u7_n86 ) );
  NOR2_X1 u0_u0_u7_U67 (.A2( u0_u0_X_45 ) , .A1( u0_u0_X_48 ) , .ZN( u0_u0_u7_n82 ) );
  NOR2_X1 u0_u0_u7_U68 (.A2( u0_u0_X_44 ) , .A1( u0_u0_u7_n14 ) , .ZN( u0_u0_u7_n83 ) );
  NOR2_X1 u0_u0_u7_U69 (.A2( u0_u0_X_46 ) , .A1( u0_u0_X_47 ) , .ZN( u0_u0_u7_n29 ) );
  OAI222_X1 u0_u0_u7_U7 (.B1( u0_u0_u7_n17 ) , .A2( u0_u0_u7_n19 ) , .C1( u0_u0_u7_n35 ) , .A1( u0_u0_u7_n68 ) , .B2( u0_u0_u7_n70 ) , .C2( u0_u0_u7_n80 ) , .ZN( u0_u0_u7_n87 ) );
  NAND2_X1 u0_u0_u7_U70 (.A2( u0_u0_X_46 ) , .A1( u0_u0_X_47 ) , .ZN( u0_u0_u7_n56 ) );
  AND2_X1 u0_u0_u7_U71 (.A1( u0_u0_X_47 ) , .A2( u0_u0_u7_n18 ) , .ZN( u0_u0_u7_n25 ) );
  AND2_X1 u0_u0_u7_U72 (.A2( u0_u0_X_45 ) , .A1( u0_u0_X_48 ) , .ZN( u0_u0_u7_n79 ) );
  AND2_X1 u0_u0_u7_U73 (.A2( u0_u0_X_43 ) , .A1( u0_u0_X_44 ) , .ZN( u0_u0_u7_n85 ) );
  AND2_X1 u0_u0_u7_U74 (.A1( u0_u0_X_44 ) , .A2( u0_u0_u7_n14 ) , .ZN( u0_u0_u7_n81 ) );
  AND2_X1 u0_u0_u7_U75 (.A1( u0_u0_X_48 ) , .A2( u0_u0_u7_n15 ) , .ZN( u0_u0_u7_n88 ) );
  INV_X1 u0_u0_u7_U76 (.A( u0_u0_X_46 ) , .ZN( u0_u0_u7_n18 ) );
  INV_X1 u0_u0_u7_U77 (.A( u0_u0_X_45 ) , .ZN( u0_u0_u7_n15 ) );
  NAND4_X1 u0_u0_u7_U78 (.ZN( u0_out0_27 ) , .A1( u0_u0_u7_n60 ) , .A2( u0_u0_u7_n61 ) , .A3( u0_u0_u7_n62 ) , .A4( u0_u0_u7_n63 ) );
  OAI21_X1 u0_u0_u7_U79 (.A( u0_u0_u7_n31 ) , .B2( u0_u0_u7_n36 ) , .ZN( u0_u0_u7_n60 ) , .B1( u0_u0_u7_n7 ) );
  OAI221_X1 u0_u0_u7_U8 (.B2( u0_u0_u7_n19 ) , .ZN( u0_u0_u7_n26 ) , .C2( u0_u0_u7_n34 ) , .C1( u0_u0_u7_n80 ) , .B1( u0_u0_u7_n89 ) , .A( u0_u0_u7_n90 ) );
  OAI21_X1 u0_u0_u7_U80 (.B2( u0_u0_u7_n11 ) , .B1( u0_u0_u7_n2 ) , .A( u0_u0_u7_n20 ) , .ZN( u0_u0_u7_n61 ) );
  NAND4_X1 u0_u0_u7_U81 (.ZN( u0_out0_21 ) , .A1( u0_u0_u7_n21 ) , .A2( u0_u0_u7_n22 ) , .A3( u0_u0_u7_n23 ) , .A4( u0_u0_u7_n24 ) );
  OAI21_X1 u0_u0_u7_U82 (.A( u0_u0_u7_n20 ) , .ZN( u0_u0_u7_n21 ) , .B1( u0_u0_u7_n36 ) , .B2( u0_u0_u7_n4 ) );
  AOI22_X1 u0_u0_u7_U83 (.ZN( u0_u0_u7_n23 ) , .A1( u0_u0_u7_n29 ) , .A2( u0_u0_u7_n30 ) , .B1( u0_u0_u7_n31 ) , .B2( u0_u0_u7_n32 ) );
  NAND4_X1 u0_u0_u7_U84 (.ZN( u0_out0_5 ) , .A2( u0_u0_u7_n58 ) , .A1( u0_u0_u7_n65 ) , .A3( u0_u0_u7_n72 ) , .A4( u0_u0_u7_n73 ) );
  AOI22_X1 u0_u0_u7_U85 (.A1( u0_u0_u7_n10 ) , .B1( u0_u0_u7_n25 ) , .B2( u0_u0_u7_n36 ) , .A2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n72 ) );
  NOR4_X1 u0_u0_u7_U86 (.ZN( u0_u0_u7_n73 ) , .A1( u0_u0_u7_n74 ) , .A2( u0_u0_u7_n75 ) , .A3( u0_u0_u7_n76 ) , .A4( u0_u0_u7_n77 ) );
  NAND4_X1 u0_u0_u7_U87 (.ZN( u0_out0_15 ) , .A1( u0_u0_u7_n3 ) , .A2( u0_u0_u7_n37 ) , .A3( u0_u0_u7_n38 ) , .A4( u0_u0_u7_n39 ) );
  OR2_X1 u0_u0_u7_U88 (.ZN( u0_u0_u7_n37 ) , .A1( u0_u0_u7_n52 ) , .A2( u0_u0_u7_n56 ) );
  AOI22_X1 u0_u0_u7_U89 (.B2( u0_u0_u7_n16 ) , .ZN( u0_u0_u7_n38 ) , .A2( u0_u0_u7_n55 ) , .A1( u0_u0_u7_n7 ) , .B1( u0_u0_u7_n8 ) );
  AND3_X1 u0_u0_u7_U9 (.A1( u0_u0_u7_n49 ) , .A2( u0_u0_u7_n54 ) , .A3( u0_u0_u7_n71 ) , .ZN( u0_u0_u7_n89 ) );
  INV_X1 u0_u0_u7_U90 (.A( u0_u0_X_43 ) , .ZN( u0_u0_u7_n14 ) );
  AOI211_X1 u0_u0_u7_U91 (.ZN( u0_u0_u7_n24 ) , .C1( u0_u0_u7_n25 ) , .A( u0_u0_u7_n26 ) , .B( u0_u0_u7_n27 ) , .C2( u0_u0_u7_n9 ) );
  OAI211_X1 u0_u0_u7_U92 (.C1( u0_u0_u7_n19 ) , .ZN( u0_u0_u7_n27 ) , .C2( u0_u0_u7_n57 ) , .A( u0_u0_u7_n58 ) , .B( u0_u0_u7_n59 ) );
  AOI222_X1 u0_u0_u7_U93 (.B2( u0_u0_u7_n11 ) , .A2( u0_u0_u7_n16 ) , .B1( u0_u0_u7_n20 ) , .C1( u0_u0_u7_n36 ) , .A1( u0_u0_u7_n5 ) , .C2( u0_u0_u7_n55 ) , .ZN( u0_u0_u7_n59 ) );
  INV_X1 u0_u0_u7_U94 (.ZN( u0_u0_u7_n11 ) , .A( u0_u0_u7_n70 ) );
  NAND3_X1 u0_u0_u7_U95 (.ZN( u0_u0_u7_n30 ) , .A1( u0_u0_u7_n33 ) , .A2( u0_u0_u7_n34 ) , .A3( u0_u0_u7_n35 ) );
  NAND3_X1 u0_u0_u7_U96 (.ZN( u0_u0_u7_n46 ) , .A1( u0_u0_u7_n48 ) , .A2( u0_u0_u7_n49 ) , .A3( u0_u0_u7_n50 ) );
  XOR2_X1 u0_u13_U10 (.B( u0_K14_45 ) , .A( u0_R12_30 ) , .Z( u0_u13_X_45 ) );
  XOR2_X1 u0_u13_U11 (.B( u0_K14_44 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_44 ) );
  XOR2_X1 u0_u13_U12 (.B( u0_K14_43 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_43 ) );
  XOR2_X1 u0_u13_U13 (.B( u0_K14_42 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_42 ) );
  XOR2_X1 u0_u13_U14 (.B( u0_K14_41 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_41 ) );
  XOR2_X1 u0_u13_U15 (.B( u0_K14_40 ) , .A( u0_R12_27 ) , .Z( u0_u13_X_40 ) );
  XOR2_X1 u0_u13_U17 (.B( u0_K14_39 ) , .A( u0_R12_26 ) , .Z( u0_u13_X_39 ) );
  XOR2_X1 u0_u13_U18 (.B( u0_K14_38 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_38 ) );
  XOR2_X1 u0_u13_U19 (.B( u0_K14_37 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_37 ) );
  XOR2_X1 u0_u13_U7 (.B( u0_K14_48 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_48 ) );
  XOR2_X1 u0_u13_U8 (.B( u0_K14_47 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_47 ) );
  XOR2_X1 u0_u13_U9 (.B( u0_K14_46 ) , .A( u0_R12_31 ) , .Z( u0_u13_X_46 ) );
  AOI22_X1 u0_u13_u6_U10 (.A2( u0_u13_u6_n151 ) , .B2( u0_u13_u6_n161 ) , .A1( u0_u13_u6_n167 ) , .B1( u0_u13_u6_n170 ) , .ZN( u0_u13_u6_n89 ) );
  AOI21_X1 u0_u13_u6_U11 (.B1( u0_u13_u6_n107 ) , .B2( u0_u13_u6_n132 ) , .A( u0_u13_u6_n158 ) , .ZN( u0_u13_u6_n88 ) );
  AOI21_X1 u0_u13_u6_U12 (.B2( u0_u13_u6_n147 ) , .B1( u0_u13_u6_n148 ) , .ZN( u0_u13_u6_n149 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U13 (.ZN( u0_u13_u6_n106 ) , .A( u0_u13_u6_n142 ) , .B2( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n164 ) );
  INV_X1 u0_u13_u6_U14 (.A( u0_u13_u6_n155 ) , .ZN( u0_u13_u6_n161 ) );
  INV_X1 u0_u13_u6_U15 (.A( u0_u13_u6_n128 ) , .ZN( u0_u13_u6_n164 ) );
  NAND2_X1 u0_u13_u6_U16 (.ZN( u0_u13_u6_n110 ) , .A1( u0_u13_u6_n122 ) , .A2( u0_u13_u6_n129 ) );
  NAND2_X1 u0_u13_u6_U17 (.ZN( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n146 ) , .A1( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U18 (.A( u0_u13_u6_n132 ) , .ZN( u0_u13_u6_n171 ) );
  AND2_X1 u0_u13_u6_U19 (.A1( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n147 ) );
  INV_X1 u0_u13_u6_U20 (.A( u0_u13_u6_n127 ) , .ZN( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U21 (.A( u0_u13_u6_n121 ) , .ZN( u0_u13_u6_n167 ) );
  INV_X1 u0_u13_u6_U22 (.A( u0_u13_u6_n100 ) , .ZN( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U23 (.A( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n170 ) );
  INV_X1 u0_u13_u6_U24 (.A( u0_u13_u6_n113 ) , .ZN( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U25 (.A1( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n119 ) , .ZN( u0_u13_u6_n133 ) );
  AND2_X1 u0_u13_u6_U26 (.A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n122 ) , .ZN( u0_u13_u6_n131 ) );
  AND3_X1 u0_u13_u6_U27 (.ZN( u0_u13_u6_n120 ) , .A2( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n132 ) , .A3( u0_u13_u6_n145 ) );
  INV_X1 u0_u13_u6_U28 (.A( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n163 ) );
  AOI222_X1 u0_u13_u6_U29 (.ZN( u0_u13_u6_n114 ) , .A1( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n126 ) , .B2( u0_u13_u6_n151 ) , .C2( u0_u13_u6_n159 ) , .C1( u0_u13_u6_n168 ) , .B1( u0_u13_u6_n169 ) );
  INV_X1 u0_u13_u6_U3 (.A( u0_u13_u6_n110 ) , .ZN( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U30 (.A1( u0_u13_u6_n162 ) , .A2( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n98 ) );
  AOI211_X1 u0_u13_u6_U31 (.B( u0_u13_u6_n134 ) , .A( u0_u13_u6_n135 ) , .C1( u0_u13_u6_n136 ) , .ZN( u0_u13_u6_n137 ) , .C2( u0_u13_u6_n151 ) );
  AOI21_X1 u0_u13_u6_U32 (.B2( u0_u13_u6_n132 ) , .B1( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n134 ) , .A( u0_u13_u6_n158 ) );
  AOI21_X1 u0_u13_u6_U33 (.B1( u0_u13_u6_n131 ) , .ZN( u0_u13_u6_n135 ) , .A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n146 ) );
  NAND4_X1 u0_u13_u6_U34 (.A4( u0_u13_u6_n127 ) , .A3( u0_u13_u6_n128 ) , .A2( u0_u13_u6_n129 ) , .A1( u0_u13_u6_n130 ) , .ZN( u0_u13_u6_n136 ) );
  NAND2_X1 u0_u13_u6_U35 (.A1( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U36 (.ZN( u0_u13_u6_n132 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n97 ) );
  AOI22_X1 u0_u13_u6_U37 (.B2( u0_u13_u6_n110 ) , .B1( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n112 ) , .ZN( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n161 ) );
  NAND4_X1 u0_u13_u6_U38 (.A3( u0_u13_u6_n109 ) , .ZN( u0_u13_u6_n112 ) , .A4( u0_u13_u6_n132 ) , .A2( u0_u13_u6_n147 ) , .A1( u0_u13_u6_n166 ) );
  NOR2_X1 u0_u13_u6_U39 (.ZN( u0_u13_u6_n109 ) , .A1( u0_u13_u6_n170 ) , .A2( u0_u13_u6_n173 ) );
  INV_X1 u0_u13_u6_U4 (.A( u0_u13_u6_n142 ) , .ZN( u0_u13_u6_n174 ) );
  NOR2_X1 u0_u13_u6_U40 (.A2( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n155 ) , .A1( u0_u13_u6_n160 ) );
  NAND2_X1 u0_u13_u6_U41 (.ZN( u0_u13_u6_n146 ) , .A2( u0_u13_u6_n94 ) , .A1( u0_u13_u6_n99 ) );
  AOI21_X1 u0_u13_u6_U42 (.A( u0_u13_u6_n144 ) , .B2( u0_u13_u6_n145 ) , .B1( u0_u13_u6_n146 ) , .ZN( u0_u13_u6_n150 ) );
  INV_X1 u0_u13_u6_U43 (.A( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n158 ) );
  NAND2_X1 u0_u13_u6_U44 (.ZN( u0_u13_u6_n127 ) , .A1( u0_u13_u6_n91 ) , .A2( u0_u13_u6_n92 ) );
  NAND2_X1 u0_u13_u6_U45 (.ZN( u0_u13_u6_n129 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n96 ) );
  INV_X1 u0_u13_u6_U46 (.A( u0_u13_u6_n144 ) , .ZN( u0_u13_u6_n159 ) );
  NAND2_X1 u0_u13_u6_U47 (.ZN( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n97 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U48 (.ZN( u0_u13_u6_n148 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n94 ) );
  NAND2_X1 u0_u13_u6_U49 (.ZN( u0_u13_u6_n108 ) , .A2( u0_u13_u6_n139 ) , .A1( u0_u13_u6_n144 ) );
  NAND2_X1 u0_u13_u6_U5 (.A2( u0_u13_u6_n143 ) , .ZN( u0_u13_u6_n152 ) , .A1( u0_u13_u6_n166 ) );
  NAND2_X1 u0_u13_u6_U50 (.ZN( u0_u13_u6_n121 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n97 ) );
  NAND2_X1 u0_u13_u6_U51 (.ZN( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n95 ) );
  AND2_X1 u0_u13_u6_U52 (.ZN( u0_u13_u6_n118 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U53 (.ZN( u0_u13_u6_n147 ) , .A2( u0_u13_u6_n98 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U54 (.ZN( u0_u13_u6_n128 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U55 (.ZN( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n95 ) , .A1( u0_u13_u6_n99 ) );
  NAND2_X1 u0_u13_u6_U56 (.ZN( u0_u13_u6_n123 ) , .A2( u0_u13_u6_n91 ) , .A1( u0_u13_u6_n96 ) );
  NAND2_X1 u0_u13_u6_U57 (.ZN( u0_u13_u6_n100 ) , .A2( u0_u13_u6_n92 ) , .A1( u0_u13_u6_n98 ) );
  NAND2_X1 u0_u13_u6_U58 (.ZN( u0_u13_u6_n122 ) , .A1( u0_u13_u6_n94 ) , .A2( u0_u13_u6_n97 ) );
  INV_X1 u0_u13_u6_U59 (.A( u0_u13_u6_n139 ) , .ZN( u0_u13_u6_n160 ) );
  AOI22_X1 u0_u13_u6_U6 (.B2( u0_u13_u6_n101 ) , .A1( u0_u13_u6_n102 ) , .ZN( u0_u13_u6_n103 ) , .B1( u0_u13_u6_n160 ) , .A2( u0_u13_u6_n161 ) );
  NAND2_X1 u0_u13_u6_U60 (.ZN( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n96 ) , .A2( u0_u13_u6_n98 ) );
  NOR2_X1 u0_u13_u6_U61 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n126 ) );
  NOR2_X1 u0_u13_u6_U62 (.A2( u0_u13_X_39 ) , .A1( u0_u13_X_42 ) , .ZN( u0_u13_u6_n92 ) );
  NOR2_X1 u0_u13_u6_U63 (.A2( u0_u13_X_39 ) , .A1( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n97 ) );
  NOR2_X1 u0_u13_u6_U64 (.A2( u0_u13_X_38 ) , .A1( u0_u13_u6_n165 ) , .ZN( u0_u13_u6_n95 ) );
  NOR2_X1 u0_u13_u6_U65 (.A2( u0_u13_X_41 ) , .ZN( u0_u13_u6_n111 ) , .A1( u0_u13_u6_n157 ) );
  NOR2_X1 u0_u13_u6_U66 (.A2( u0_u13_X_37 ) , .A1( u0_u13_u6_n162 ) , .ZN( u0_u13_u6_n94 ) );
  NOR2_X1 u0_u13_u6_U67 (.A2( u0_u13_X_37 ) , .A1( u0_u13_X_38 ) , .ZN( u0_u13_u6_n91 ) );
  NAND2_X1 u0_u13_u6_U68 (.A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n144 ) , .A2( u0_u13_u6_n157 ) );
  NAND2_X1 u0_u13_u6_U69 (.A2( u0_u13_X_40 ) , .A1( u0_u13_X_41 ) , .ZN( u0_u13_u6_n139 ) );
  NOR2_X1 u0_u13_u6_U7 (.A1( u0_u13_u6_n118 ) , .ZN( u0_u13_u6_n143 ) , .A2( u0_u13_u6_n168 ) );
  AND2_X1 u0_u13_u6_U70 (.A1( u0_u13_X_39 ) , .A2( u0_u13_u6_n156 ) , .ZN( u0_u13_u6_n96 ) );
  AND2_X1 u0_u13_u6_U71 (.A1( u0_u13_X_39 ) , .A2( u0_u13_X_42 ) , .ZN( u0_u13_u6_n99 ) );
  INV_X1 u0_u13_u6_U72 (.A( u0_u13_X_40 ) , .ZN( u0_u13_u6_n157 ) );
  INV_X1 u0_u13_u6_U73 (.A( u0_u13_X_37 ) , .ZN( u0_u13_u6_n165 ) );
  INV_X1 u0_u13_u6_U74 (.A( u0_u13_X_38 ) , .ZN( u0_u13_u6_n162 ) );
  INV_X1 u0_u13_u6_U75 (.A( u0_u13_X_42 ) , .ZN( u0_u13_u6_n156 ) );
  NAND4_X1 u0_u13_u6_U76 (.ZN( u0_out13_32 ) , .A4( u0_u13_u6_n103 ) , .A3( u0_u13_u6_n104 ) , .A2( u0_u13_u6_n105 ) , .A1( u0_u13_u6_n106 ) );
  AOI22_X1 u0_u13_u6_U77 (.ZN( u0_u13_u6_n105 ) , .A2( u0_u13_u6_n108 ) , .A1( u0_u13_u6_n118 ) , .B2( u0_u13_u6_n126 ) , .B1( u0_u13_u6_n171 ) );
  AOI22_X1 u0_u13_u6_U78 (.ZN( u0_u13_u6_n104 ) , .A1( u0_u13_u6_n111 ) , .B1( u0_u13_u6_n124 ) , .B2( u0_u13_u6_n151 ) , .A2( u0_u13_u6_n93 ) );
  NAND4_X1 u0_u13_u6_U79 (.ZN( u0_out13_12 ) , .A4( u0_u13_u6_n114 ) , .A3( u0_u13_u6_n115 ) , .A2( u0_u13_u6_n116 ) , .A1( u0_u13_u6_n117 ) );
  OAI21_X1 u0_u13_u6_U8 (.A( u0_u13_u6_n159 ) , .B1( u0_u13_u6_n169 ) , .B2( u0_u13_u6_n173 ) , .ZN( u0_u13_u6_n90 ) );
  OAI22_X1 u0_u13_u6_U80 (.B2( u0_u13_u6_n111 ) , .ZN( u0_u13_u6_n116 ) , .B1( u0_u13_u6_n126 ) , .A2( u0_u13_u6_n164 ) , .A1( u0_u13_u6_n167 ) );
  OAI21_X1 u0_u13_u6_U81 (.A( u0_u13_u6_n108 ) , .ZN( u0_u13_u6_n117 ) , .B2( u0_u13_u6_n141 ) , .B1( u0_u13_u6_n163 ) );
  OAI211_X1 u0_u13_u6_U82 (.ZN( u0_out13_7 ) , .B( u0_u13_u6_n153 ) , .C2( u0_u13_u6_n154 ) , .C1( u0_u13_u6_n155 ) , .A( u0_u13_u6_n174 ) );
  NOR3_X1 u0_u13_u6_U83 (.A1( u0_u13_u6_n141 ) , .ZN( u0_u13_u6_n154 ) , .A3( u0_u13_u6_n164 ) , .A2( u0_u13_u6_n171 ) );
  AOI211_X1 u0_u13_u6_U84 (.B( u0_u13_u6_n149 ) , .A( u0_u13_u6_n150 ) , .C2( u0_u13_u6_n151 ) , .C1( u0_u13_u6_n152 ) , .ZN( u0_u13_u6_n153 ) );
  OAI211_X1 u0_u13_u6_U85 (.ZN( u0_out13_22 ) , .B( u0_u13_u6_n137 ) , .A( u0_u13_u6_n138 ) , .C2( u0_u13_u6_n139 ) , .C1( u0_u13_u6_n140 ) );
  AOI22_X1 u0_u13_u6_U86 (.B1( u0_u13_u6_n124 ) , .A2( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n126 ) , .ZN( u0_u13_u6_n138 ) , .B2( u0_u13_u6_n161 ) );
  AND4_X1 u0_u13_u6_U87 (.A3( u0_u13_u6_n119 ) , .A1( u0_u13_u6_n120 ) , .A4( u0_u13_u6_n129 ) , .ZN( u0_u13_u6_n140 ) , .A2( u0_u13_u6_n143 ) );
  NAND3_X1 u0_u13_u6_U88 (.A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n125 ) , .A1( u0_u13_u6_n130 ) , .A3( u0_u13_u6_n131 ) );
  NAND3_X1 u0_u13_u6_U89 (.A3( u0_u13_u6_n133 ) , .ZN( u0_u13_u6_n141 ) , .A1( u0_u13_u6_n145 ) , .A2( u0_u13_u6_n148 ) );
  INV_X1 u0_u13_u6_U9 (.ZN( u0_u13_u6_n172 ) , .A( u0_u13_u6_n88 ) );
  NAND3_X1 u0_u13_u6_U90 (.ZN( u0_u13_u6_n101 ) , .A3( u0_u13_u6_n107 ) , .A2( u0_u13_u6_n121 ) , .A1( u0_u13_u6_n127 ) );
  NAND3_X1 u0_u13_u6_U91 (.ZN( u0_u13_u6_n102 ) , .A3( u0_u13_u6_n130 ) , .A2( u0_u13_u6_n145 ) , .A1( u0_u13_u6_n166 ) );
  NAND3_X1 u0_u13_u6_U92 (.A3( u0_u13_u6_n113 ) , .A1( u0_u13_u6_n119 ) , .A2( u0_u13_u6_n123 ) , .ZN( u0_u13_u6_n93 ) );
  NAND3_X1 u0_u13_u6_U93 (.ZN( u0_u13_u6_n142 ) , .A2( u0_u13_u6_n172 ) , .A3( u0_u13_u6_n89 ) , .A1( u0_u13_u6_n90 ) );
  AND3_X1 u0_u13_u7_U10 (.A3( u0_u13_u7_n110 ) , .A2( u0_u13_u7_n127 ) , .A1( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n92 ) );
  OAI21_X1 u0_u13_u7_U11 (.A( u0_u13_u7_n161 ) , .B1( u0_u13_u7_n168 ) , .B2( u0_u13_u7_n173 ) , .ZN( u0_u13_u7_n91 ) );
  AOI211_X1 u0_u13_u7_U12 (.A( u0_u13_u7_n117 ) , .ZN( u0_u13_u7_n118 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n177 ) , .B( u0_u13_u7_n180 ) );
  OAI22_X1 u0_u13_u7_U13 (.B1( u0_u13_u7_n115 ) , .ZN( u0_u13_u7_n117 ) , .A2( u0_u13_u7_n133 ) , .A1( u0_u13_u7_n137 ) , .B2( u0_u13_u7_n162 ) );
  INV_X1 u0_u13_u7_U14 (.A( u0_u13_u7_n116 ) , .ZN( u0_u13_u7_n180 ) );
  NOR3_X1 u0_u13_u7_U15 (.ZN( u0_u13_u7_n115 ) , .A3( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n168 ) , .A1( u0_u13_u7_n169 ) );
  OAI211_X1 u0_u13_u7_U16 (.B( u0_u13_u7_n122 ) , .A( u0_u13_u7_n123 ) , .C2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n154 ) , .C1( u0_u13_u7_n162 ) );
  AOI222_X1 u0_u13_u7_U17 (.ZN( u0_u13_u7_n122 ) , .C2( u0_u13_u7_n126 ) , .C1( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n161 ) , .A2( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n170 ) , .A1( u0_u13_u7_n176 ) );
  INV_X1 u0_u13_u7_U18 (.A( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n176 ) );
  NOR3_X1 u0_u13_u7_U19 (.A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n135 ) , .ZN( u0_u13_u7_n136 ) , .A3( u0_u13_u7_n171 ) );
  NOR2_X1 u0_u13_u7_U20 (.A1( u0_u13_u7_n130 ) , .A2( u0_u13_u7_n134 ) , .ZN( u0_u13_u7_n153 ) );
  INV_X1 u0_u13_u7_U21 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n165 ) );
  NOR2_X1 u0_u13_u7_U22 (.ZN( u0_u13_u7_n111 ) , .A2( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n169 ) );
  AOI21_X1 u0_u13_u7_U23 (.ZN( u0_u13_u7_n104 ) , .B2( u0_u13_u7_n112 ) , .B1( u0_u13_u7_n127 ) , .A( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U24 (.ZN( u0_u13_u7_n106 ) , .B1( u0_u13_u7_n133 ) , .B2( u0_u13_u7_n146 ) , .A( u0_u13_u7_n162 ) );
  AOI21_X1 u0_u13_u7_U25 (.A( u0_u13_u7_n101 ) , .ZN( u0_u13_u7_n107 ) , .B2( u0_u13_u7_n128 ) , .B1( u0_u13_u7_n175 ) );
  INV_X1 u0_u13_u7_U26 (.A( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n171 ) );
  INV_X1 u0_u13_u7_U27 (.A( u0_u13_u7_n131 ) , .ZN( u0_u13_u7_n177 ) );
  INV_X1 u0_u13_u7_U28 (.A( u0_u13_u7_n110 ) , .ZN( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U29 (.A1( u0_u13_u7_n129 ) , .A2( u0_u13_u7_n132 ) , .ZN( u0_u13_u7_n149 ) );
  OAI21_X1 u0_u13_u7_U3 (.ZN( u0_u13_u7_n159 ) , .A( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n171 ) , .B1( u0_u13_u7_n174 ) );
  NAND2_X1 u0_u13_u7_U30 (.A1( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n124 ) , .ZN( u0_u13_u7_n130 ) );
  INV_X1 u0_u13_u7_U31 (.A( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n173 ) );
  INV_X1 u0_u13_u7_U32 (.A( u0_u13_u7_n128 ) , .ZN( u0_u13_u7_n168 ) );
  INV_X1 u0_u13_u7_U33 (.A( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n169 ) );
  INV_X1 u0_u13_u7_U34 (.A( u0_u13_u7_n127 ) , .ZN( u0_u13_u7_n179 ) );
  NOR2_X1 u0_u13_u7_U35 (.ZN( u0_u13_u7_n101 ) , .A2( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n156 ) );
  AOI211_X1 u0_u13_u7_U36 (.B( u0_u13_u7_n154 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n156 ) , .ZN( u0_u13_u7_n157 ) , .C2( u0_u13_u7_n172 ) );
  INV_X1 u0_u13_u7_U37 (.A( u0_u13_u7_n153 ) , .ZN( u0_u13_u7_n172 ) );
  AOI211_X1 u0_u13_u7_U38 (.B( u0_u13_u7_n139 ) , .A( u0_u13_u7_n140 ) , .C2( u0_u13_u7_n141 ) , .ZN( u0_u13_u7_n142 ) , .C1( u0_u13_u7_n156 ) );
  NAND4_X1 u0_u13_u7_U39 (.A3( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n141 ) , .A4( u0_u13_u7_n147 ) );
  INV_X1 u0_u13_u7_U4 (.A( u0_u13_u7_n111 ) , .ZN( u0_u13_u7_n170 ) );
  AOI21_X1 u0_u13_u7_U40 (.A( u0_u13_u7_n137 ) , .B1( u0_u13_u7_n138 ) , .ZN( u0_u13_u7_n139 ) , .B2( u0_u13_u7_n146 ) );
  OAI22_X1 u0_u13_u7_U41 (.B1( u0_u13_u7_n136 ) , .ZN( u0_u13_u7_n140 ) , .A1( u0_u13_u7_n153 ) , .B2( u0_u13_u7_n162 ) , .A2( u0_u13_u7_n164 ) );
  AOI21_X1 u0_u13_u7_U42 (.ZN( u0_u13_u7_n123 ) , .B1( u0_u13_u7_n165 ) , .B2( u0_u13_u7_n177 ) , .A( u0_u13_u7_n97 ) );
  AOI21_X1 u0_u13_u7_U43 (.B2( u0_u13_u7_n113 ) , .B1( u0_u13_u7_n124 ) , .A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n97 ) );
  INV_X1 u0_u13_u7_U44 (.A( u0_u13_u7_n125 ) , .ZN( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U45 (.A( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n162 ) );
  AOI22_X1 u0_u13_u7_U46 (.A2( u0_u13_u7_n114 ) , .ZN( u0_u13_u7_n119 ) , .B1( u0_u13_u7_n130 ) , .A1( u0_u13_u7_n156 ) , .B2( u0_u13_u7_n165 ) );
  NAND2_X1 u0_u13_u7_U47 (.A2( u0_u13_u7_n112 ) , .ZN( u0_u13_u7_n114 ) , .A1( u0_u13_u7_n175 ) );
  AND2_X1 u0_u13_u7_U48 (.ZN( u0_u13_u7_n145 ) , .A2( u0_u13_u7_n98 ) , .A1( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U49 (.ZN( u0_u13_u7_n137 ) , .A1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n161 ) );
  INV_X1 u0_u13_u7_U5 (.A( u0_u13_u7_n149 ) , .ZN( u0_u13_u7_n175 ) );
  AOI21_X1 u0_u13_u7_U50 (.ZN( u0_u13_u7_n105 ) , .B2( u0_u13_u7_n110 ) , .A( u0_u13_u7_n125 ) , .B1( u0_u13_u7_n147 ) );
  NAND2_X1 u0_u13_u7_U51 (.ZN( u0_u13_u7_n146 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U52 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U53 (.A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n127 ) , .A2( u0_u13_u7_n99 ) );
  OR2_X1 u0_u13_u7_U54 (.ZN( u0_u13_u7_n126 ) , .A2( u0_u13_u7_n152 ) , .A1( u0_u13_u7_n156 ) );
  NAND2_X1 u0_u13_u7_U55 (.A2( u0_u13_u7_n102 ) , .A1( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n133 ) );
  NAND2_X1 u0_u13_u7_U56 (.ZN( u0_u13_u7_n112 ) , .A2( u0_u13_u7_n96 ) , .A1( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U57 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n128 ) , .A1( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U58 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n113 ) , .A2( u0_u13_u7_n93 ) );
  NAND2_X1 u0_u13_u7_U59 (.A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n124 ) , .A1( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U6 (.A( u0_u13_u7_n154 ) , .ZN( u0_u13_u7_n178 ) );
  NAND2_X1 u0_u13_u7_U60 (.ZN( u0_u13_u7_n110 ) , .A1( u0_u13_u7_n95 ) , .A2( u0_u13_u7_n96 ) );
  INV_X1 u0_u13_u7_U61 (.A( u0_u13_u7_n150 ) , .ZN( u0_u13_u7_n164 ) );
  AND2_X1 u0_u13_u7_U62 (.ZN( u0_u13_u7_n134 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n98 ) );
  NAND2_X1 u0_u13_u7_U63 (.A1( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n102 ) , .ZN( u0_u13_u7_n129 ) );
  NAND2_X1 u0_u13_u7_U64 (.A2( u0_u13_u7_n103 ) , .ZN( u0_u13_u7_n131 ) , .A1( u0_u13_u7_n95 ) );
  NAND2_X1 u0_u13_u7_U65 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n138 ) , .A2( u0_u13_u7_n99 ) );
  NAND2_X1 u0_u13_u7_U66 (.ZN( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n93 ) , .A2( u0_u13_u7_n96 ) );
  NAND2_X1 u0_u13_u7_U67 (.A1( u0_u13_u7_n100 ) , .ZN( u0_u13_u7_n148 ) , .A2( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U68 (.A2( u0_u13_X_47 ) , .ZN( u0_u13_u7_n150 ) , .A1( u0_u13_u7_n163 ) );
  NOR2_X1 u0_u13_u7_U69 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n103 ) );
  AOI211_X1 u0_u13_u7_U7 (.ZN( u0_u13_u7_n116 ) , .A( u0_u13_u7_n155 ) , .C1( u0_u13_u7_n161 ) , .C2( u0_u13_u7_n171 ) , .B( u0_u13_u7_n94 ) );
  NOR2_X1 u0_u13_u7_U70 (.A2( u0_u13_X_48 ) , .A1( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n95 ) );
  NOR2_X1 u0_u13_u7_U71 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n99 ) );
  NOR2_X1 u0_u13_u7_U72 (.A2( u0_u13_X_44 ) , .A1( u0_u13_u7_n167 ) , .ZN( u0_u13_u7_n98 ) );
  NOR2_X1 u0_u13_u7_U73 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n152 ) );
  AND2_X1 u0_u13_u7_U74 (.A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n156 ) , .A2( u0_u13_u7_n163 ) );
  NAND2_X1 u0_u13_u7_U75 (.A2( u0_u13_X_46 ) , .A1( u0_u13_X_47 ) , .ZN( u0_u13_u7_n125 ) );
  AND2_X1 u0_u13_u7_U76 (.A2( u0_u13_X_45 ) , .A1( u0_u13_X_48 ) , .ZN( u0_u13_u7_n102 ) );
  AND2_X1 u0_u13_u7_U77 (.A2( u0_u13_X_43 ) , .A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n96 ) );
  AND2_X1 u0_u13_u7_U78 (.A1( u0_u13_X_44 ) , .ZN( u0_u13_u7_n100 ) , .A2( u0_u13_u7_n167 ) );
  AND2_X1 u0_u13_u7_U79 (.A1( u0_u13_X_48 ) , .A2( u0_u13_u7_n166 ) , .ZN( u0_u13_u7_n93 ) );
  OAI222_X1 u0_u13_u7_U8 (.C2( u0_u13_u7_n101 ) , .B2( u0_u13_u7_n111 ) , .A1( u0_u13_u7_n113 ) , .C1( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n162 ) , .B1( u0_u13_u7_n164 ) , .ZN( u0_u13_u7_n94 ) );
  INV_X1 u0_u13_u7_U80 (.A( u0_u13_X_46 ) , .ZN( u0_u13_u7_n163 ) );
  INV_X1 u0_u13_u7_U81 (.A( u0_u13_X_43 ) , .ZN( u0_u13_u7_n167 ) );
  INV_X1 u0_u13_u7_U82 (.A( u0_u13_X_45 ) , .ZN( u0_u13_u7_n166 ) );
  NAND4_X1 u0_u13_u7_U83 (.ZN( u0_out13_27 ) , .A4( u0_u13_u7_n118 ) , .A3( u0_u13_u7_n119 ) , .A2( u0_u13_u7_n120 ) , .A1( u0_u13_u7_n121 ) );
  OAI21_X1 u0_u13_u7_U84 (.ZN( u0_u13_u7_n121 ) , .B2( u0_u13_u7_n145 ) , .A( u0_u13_u7_n150 ) , .B1( u0_u13_u7_n174 ) );
  OAI21_X1 u0_u13_u7_U85 (.ZN( u0_u13_u7_n120 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n170 ) , .B1( u0_u13_u7_n179 ) );
  NAND4_X1 u0_u13_u7_U86 (.ZN( u0_out13_21 ) , .A4( u0_u13_u7_n157 ) , .A3( u0_u13_u7_n158 ) , .A2( u0_u13_u7_n159 ) , .A1( u0_u13_u7_n160 ) );
  OAI21_X1 u0_u13_u7_U87 (.B1( u0_u13_u7_n145 ) , .ZN( u0_u13_u7_n160 ) , .A( u0_u13_u7_n161 ) , .B2( u0_u13_u7_n177 ) );
  AOI22_X1 u0_u13_u7_U88 (.B2( u0_u13_u7_n149 ) , .B1( u0_u13_u7_n150 ) , .A2( u0_u13_u7_n151 ) , .A1( u0_u13_u7_n152 ) , .ZN( u0_u13_u7_n158 ) );
  NAND4_X1 u0_u13_u7_U89 (.ZN( u0_out13_15 ) , .A4( u0_u13_u7_n142 ) , .A3( u0_u13_u7_n143 ) , .A2( u0_u13_u7_n144 ) , .A1( u0_u13_u7_n178 ) );
  OAI221_X1 u0_u13_u7_U9 (.C1( u0_u13_u7_n101 ) , .C2( u0_u13_u7_n147 ) , .ZN( u0_u13_u7_n155 ) , .B2( u0_u13_u7_n162 ) , .A( u0_u13_u7_n91 ) , .B1( u0_u13_u7_n92 ) );
  OR2_X1 u0_u13_u7_U90 (.A2( u0_u13_u7_n125 ) , .A1( u0_u13_u7_n129 ) , .ZN( u0_u13_u7_n144 ) );
  AOI22_X1 u0_u13_u7_U91 (.A2( u0_u13_u7_n126 ) , .ZN( u0_u13_u7_n143 ) , .B2( u0_u13_u7_n165 ) , .B1( u0_u13_u7_n173 ) , .A1( u0_u13_u7_n174 ) );
  NAND4_X1 u0_u13_u7_U92 (.ZN( u0_out13_5 ) , .A4( u0_u13_u7_n108 ) , .A3( u0_u13_u7_n109 ) , .A1( u0_u13_u7_n116 ) , .A2( u0_u13_u7_n123 ) );
  AOI22_X1 u0_u13_u7_U93 (.ZN( u0_u13_u7_n109 ) , .A2( u0_u13_u7_n126 ) , .B2( u0_u13_u7_n145 ) , .B1( u0_u13_u7_n156 ) , .A1( u0_u13_u7_n171 ) );
  NOR4_X1 u0_u13_u7_U94 (.A4( u0_u13_u7_n104 ) , .A3( u0_u13_u7_n105 ) , .A2( u0_u13_u7_n106 ) , .A1( u0_u13_u7_n107 ) , .ZN( u0_u13_u7_n108 ) );
  NAND3_X1 u0_u13_u7_U95 (.A3( u0_u13_u7_n146 ) , .A2( u0_u13_u7_n147 ) , .A1( u0_u13_u7_n148 ) , .ZN( u0_u13_u7_n151 ) );
  NAND3_X1 u0_u13_u7_U96 (.A3( u0_u13_u7_n131 ) , .A2( u0_u13_u7_n132 ) , .A1( u0_u13_u7_n133 ) , .ZN( u0_u13_u7_n135 ) );
  XOR2_X1 u0_u4_U10 (.B( u0_K5_45 ) , .A( u0_R3_30 ) , .Z( u0_u4_X_45 ) );
  XOR2_X1 u0_u4_U11 (.B( u0_K5_44 ) , .A( u0_R3_29 ) , .Z( u0_u4_X_44 ) );
  XOR2_X1 u0_u4_U12 (.B( u0_K5_43 ) , .A( u0_R3_28 ) , .Z( u0_u4_X_43 ) );
  XOR2_X1 u0_u4_U13 (.B( u0_K5_42 ) , .A( u0_R3_29 ) , .Z( u0_u4_X_42 ) );
  XOR2_X1 u0_u4_U14 (.B( u0_K5_41 ) , .A( u0_R3_28 ) , .Z( u0_u4_X_41 ) );
  XOR2_X1 u0_u4_U15 (.B( u0_K5_40 ) , .A( u0_R3_27 ) , .Z( u0_u4_X_40 ) );
  XOR2_X1 u0_u4_U16 (.B( u0_K5_3 ) , .A( u0_R3_2 ) , .Z( u0_u4_X_3 ) );
  XOR2_X1 u0_u4_U17 (.B( u0_K5_39 ) , .A( u0_R3_26 ) , .Z( u0_u4_X_39 ) );
  XOR2_X1 u0_u4_U18 (.B( u0_K5_38 ) , .A( u0_R3_25 ) , .Z( u0_u4_X_38 ) );
  XOR2_X1 u0_u4_U19 (.B( u0_K5_37 ) , .A( u0_R3_24 ) , .Z( u0_u4_X_37 ) );
  XOR2_X1 u0_u4_U20 (.B( u0_K5_36 ) , .A( u0_R3_25 ) , .Z( u0_u4_X_36 ) );
  XOR2_X1 u0_u4_U21 (.B( u0_K5_35 ) , .A( u0_R3_24 ) , .Z( u0_u4_X_35 ) );
  XOR2_X1 u0_u4_U22 (.B( u0_K5_34 ) , .A( u0_R3_23 ) , .Z( u0_u4_X_34 ) );
  XOR2_X1 u0_u4_U23 (.B( u0_K5_33 ) , .A( u0_R3_22 ) , .Z( u0_u4_X_33 ) );
  XOR2_X1 u0_u4_U24 (.B( u0_K5_32 ) , .A( u0_R3_21 ) , .Z( u0_u4_X_32 ) );
  XOR2_X1 u0_u4_U25 (.B( u0_K5_31 ) , .A( u0_R3_20 ) , .Z( u0_u4_X_31 ) );
  XOR2_X1 u0_u4_U27 (.B( u0_K5_2 ) , .A( u0_R3_1 ) , .Z( u0_u4_X_2 ) );
  XOR2_X1 u0_u4_U38 (.B( u0_K5_1 ) , .A( u0_R3_32 ) , .Z( u0_u4_X_1 ) );
  XOR2_X1 u0_u4_U4 (.B( u0_K5_6 ) , .A( u0_R3_5 ) , .Z( u0_u4_X_6 ) );
  XOR2_X1 u0_u4_U5 (.B( u0_K5_5 ) , .A( u0_R3_4 ) , .Z( u0_u4_X_5 ) );
  XOR2_X1 u0_u4_U6 (.B( u0_K5_4 ) , .A( u0_R3_3 ) , .Z( u0_u4_X_4 ) );
  XOR2_X1 u0_u4_U7 (.B( u0_K5_48 ) , .A( u0_R3_1 ) , .Z( u0_u4_X_48 ) );
  XOR2_X1 u0_u4_U8 (.B( u0_K5_47 ) , .A( u0_R3_32 ) , .Z( u0_u4_X_47 ) );
  XOR2_X1 u0_u4_U9 (.B( u0_K5_46 ) , .A( u0_R3_31 ) , .Z( u0_u4_X_46 ) );
  AND3_X1 u0_u4_u0_U10 (.A2( u0_u4_u0_n112 ) , .ZN( u0_u4_u0_n127 ) , .A3( u0_u4_u0_n130 ) , .A1( u0_u4_u0_n148 ) );
  NAND2_X1 u0_u4_u0_U11 (.ZN( u0_u4_u0_n113 ) , .A1( u0_u4_u0_n139 ) , .A2( u0_u4_u0_n149 ) );
  AND2_X1 u0_u4_u0_U12 (.ZN( u0_u4_u0_n107 ) , .A1( u0_u4_u0_n130 ) , .A2( u0_u4_u0_n140 ) );
  AND2_X1 u0_u4_u0_U13 (.A2( u0_u4_u0_n129 ) , .A1( u0_u4_u0_n130 ) , .ZN( u0_u4_u0_n151 ) );
  AND2_X1 u0_u4_u0_U14 (.A1( u0_u4_u0_n108 ) , .A2( u0_u4_u0_n125 ) , .ZN( u0_u4_u0_n145 ) );
  INV_X1 u0_u4_u0_U15 (.A( u0_u4_u0_n143 ) , .ZN( u0_u4_u0_n173 ) );
  NOR2_X1 u0_u4_u0_U16 (.A2( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n147 ) , .A1( u0_u4_u0_n160 ) );
  INV_X1 u0_u4_u0_U17 (.ZN( u0_u4_u0_n172 ) , .A( u0_u4_u0_n88 ) );
  OAI222_X1 u0_u4_u0_U18 (.C1( u0_u4_u0_n108 ) , .A1( u0_u4_u0_n125 ) , .B2( u0_u4_u0_n128 ) , .B1( u0_u4_u0_n144 ) , .A2( u0_u4_u0_n158 ) , .C2( u0_u4_u0_n161 ) , .ZN( u0_u4_u0_n88 ) );
  AOI21_X1 u0_u4_u0_U19 (.B1( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n132 ) , .A( u0_u4_u0_n165 ) , .B2( u0_u4_u0_n93 ) );
  INV_X1 u0_u4_u0_U20 (.A( u0_u4_u0_n142 ) , .ZN( u0_u4_u0_n165 ) );
  OAI221_X1 u0_u4_u0_U21 (.C1( u0_u4_u0_n112 ) , .ZN( u0_u4_u0_n120 ) , .B1( u0_u4_u0_n138 ) , .B2( u0_u4_u0_n141 ) , .C2( u0_u4_u0_n147 ) , .A( u0_u4_u0_n172 ) );
  AOI211_X1 u0_u4_u0_U22 (.B( u0_u4_u0_n115 ) , .A( u0_u4_u0_n116 ) , .C2( u0_u4_u0_n117 ) , .C1( u0_u4_u0_n118 ) , .ZN( u0_u4_u0_n119 ) );
  OAI22_X1 u0_u4_u0_U23 (.B1( u0_u4_u0_n125 ) , .ZN( u0_u4_u0_n126 ) , .A1( u0_u4_u0_n138 ) , .A2( u0_u4_u0_n146 ) , .B2( u0_u4_u0_n147 ) );
  OAI22_X1 u0_u4_u0_U24 (.B1( u0_u4_u0_n131 ) , .A1( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n147 ) , .A2( u0_u4_u0_n90 ) , .ZN( u0_u4_u0_n91 ) );
  AND3_X1 u0_u4_u0_U25 (.A3( u0_u4_u0_n121 ) , .A2( u0_u4_u0_n125 ) , .A1( u0_u4_u0_n148 ) , .ZN( u0_u4_u0_n90 ) );
  INV_X1 u0_u4_u0_U26 (.A( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n161 ) );
  AOI22_X1 u0_u4_u0_U27 (.B2( u0_u4_u0_n109 ) , .A2( u0_u4_u0_n110 ) , .ZN( u0_u4_u0_n111 ) , .B1( u0_u4_u0_n118 ) , .A1( u0_u4_u0_n160 ) );
  INV_X1 u0_u4_u0_U28 (.A( u0_u4_u0_n118 ) , .ZN( u0_u4_u0_n158 ) );
  AOI21_X1 u0_u4_u0_U29 (.ZN( u0_u4_u0_n104 ) , .B1( u0_u4_u0_n107 ) , .B2( u0_u4_u0_n141 ) , .A( u0_u4_u0_n144 ) );
  INV_X1 u0_u4_u0_U3 (.A( u0_u4_u0_n113 ) , .ZN( u0_u4_u0_n166 ) );
  AOI21_X1 u0_u4_u0_U30 (.B1( u0_u4_u0_n127 ) , .B2( u0_u4_u0_n129 ) , .A( u0_u4_u0_n138 ) , .ZN( u0_u4_u0_n96 ) );
  AOI21_X1 u0_u4_u0_U31 (.ZN( u0_u4_u0_n116 ) , .B2( u0_u4_u0_n142 ) , .A( u0_u4_u0_n144 ) , .B1( u0_u4_u0_n166 ) );
  NAND2_X1 u0_u4_u0_U32 (.A1( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n128 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U33 (.A1( u0_u4_u0_n100 ) , .A2( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n125 ) );
  NAND2_X1 u0_u4_u0_U34 (.ZN( u0_u4_u0_n148 ) , .A1( u0_u4_u0_n93 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U35 (.A1( u0_u4_u0_n101 ) , .A2( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n150 ) );
  INV_X1 u0_u4_u0_U36 (.A( u0_u4_u0_n138 ) , .ZN( u0_u4_u0_n160 ) );
  NAND2_X1 u0_u4_u0_U37 (.A1( u0_u4_u0_n100 ) , .ZN( u0_u4_u0_n129 ) , .A2( u0_u4_u0_n95 ) );
  NAND2_X1 u0_u4_u0_U38 (.A2( u0_u4_u0_n102 ) , .A1( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n149 ) );
  NAND2_X1 u0_u4_u0_U39 (.A2( u0_u4_u0_n100 ) , .A1( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n139 ) );
  AOI21_X1 u0_u4_u0_U4 (.B1( u0_u4_u0_n114 ) , .ZN( u0_u4_u0_n115 ) , .B2( u0_u4_u0_n129 ) , .A( u0_u4_u0_n161 ) );
  NAND2_X1 u0_u4_u0_U40 (.A2( u0_u4_u0_n100 ) , .ZN( u0_u4_u0_n131 ) , .A1( u0_u4_u0_n92 ) );
  NAND2_X1 u0_u4_u0_U41 (.A2( u0_u4_u0_n102 ) , .ZN( u0_u4_u0_n114 ) , .A1( u0_u4_u0_n92 ) );
  NAND2_X1 u0_u4_u0_U42 (.A2( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n121 ) , .A1( u0_u4_u0_n93 ) );
  NAND2_X1 u0_u4_u0_U43 (.ZN( u0_u4_u0_n112 ) , .A2( u0_u4_u0_n92 ) , .A1( u0_u4_u0_n93 ) );
  OR3_X1 u0_u4_u0_U44 (.A3( u0_u4_u0_n152 ) , .A2( u0_u4_u0_n153 ) , .A1( u0_u4_u0_n154 ) , .ZN( u0_u4_u0_n155 ) );
  AOI21_X1 u0_u4_u0_U45 (.B2( u0_u4_u0_n150 ) , .B1( u0_u4_u0_n151 ) , .ZN( u0_u4_u0_n152 ) , .A( u0_u4_u0_n158 ) );
  AOI21_X1 u0_u4_u0_U46 (.A( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n145 ) , .B1( u0_u4_u0_n146 ) , .ZN( u0_u4_u0_n154 ) );
  AOI21_X1 u0_u4_u0_U47 (.A( u0_u4_u0_n147 ) , .B2( u0_u4_u0_n148 ) , .B1( u0_u4_u0_n149 ) , .ZN( u0_u4_u0_n153 ) );
  INV_X1 u0_u4_u0_U48 (.ZN( u0_u4_u0_n171 ) , .A( u0_u4_u0_n99 ) );
  OAI211_X1 u0_u4_u0_U49 (.C2( u0_u4_u0_n140 ) , .C1( u0_u4_u0_n161 ) , .A( u0_u4_u0_n169 ) , .B( u0_u4_u0_n98 ) , .ZN( u0_u4_u0_n99 ) );
  AOI21_X1 u0_u4_u0_U5 (.B2( u0_u4_u0_n131 ) , .ZN( u0_u4_u0_n134 ) , .B1( u0_u4_u0_n151 ) , .A( u0_u4_u0_n158 ) );
  AOI211_X1 u0_u4_u0_U50 (.C1( u0_u4_u0_n118 ) , .A( u0_u4_u0_n123 ) , .B( u0_u4_u0_n96 ) , .C2( u0_u4_u0_n97 ) , .ZN( u0_u4_u0_n98 ) );
  INV_X1 u0_u4_u0_U51 (.ZN( u0_u4_u0_n169 ) , .A( u0_u4_u0_n91 ) );
  NOR2_X1 u0_u4_u0_U52 (.A2( u0_u4_X_6 ) , .ZN( u0_u4_u0_n100 ) , .A1( u0_u4_u0_n162 ) );
  NOR2_X1 u0_u4_u0_U53 (.A2( u0_u4_X_4 ) , .A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n118 ) );
  NOR2_X1 u0_u4_u0_U54 (.A2( u0_u4_X_2 ) , .ZN( u0_u4_u0_n103 ) , .A1( u0_u4_u0_n164 ) );
  NOR2_X1 u0_u4_u0_U55 (.A2( u0_u4_X_1 ) , .A1( u0_u4_X_2 ) , .ZN( u0_u4_u0_n92 ) );
  NOR2_X1 u0_u4_u0_U56 (.A2( u0_u4_X_1 ) , .ZN( u0_u4_u0_n101 ) , .A1( u0_u4_u0_n163 ) );
  NAND2_X1 u0_u4_u0_U57 (.A2( u0_u4_X_4 ) , .A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n144 ) );
  NOR2_X1 u0_u4_u0_U58 (.A2( u0_u4_X_5 ) , .ZN( u0_u4_u0_n136 ) , .A1( u0_u4_u0_n159 ) );
  NAND2_X1 u0_u4_u0_U59 (.A1( u0_u4_X_5 ) , .ZN( u0_u4_u0_n138 ) , .A2( u0_u4_u0_n159 ) );
  NOR2_X1 u0_u4_u0_U6 (.A1( u0_u4_u0_n108 ) , .ZN( u0_u4_u0_n123 ) , .A2( u0_u4_u0_n158 ) );
  AND2_X1 u0_u4_u0_U60 (.A2( u0_u4_X_3 ) , .A1( u0_u4_X_6 ) , .ZN( u0_u4_u0_n102 ) );
  AND2_X1 u0_u4_u0_U61 (.A1( u0_u4_X_6 ) , .A2( u0_u4_u0_n162 ) , .ZN( u0_u4_u0_n93 ) );
  INV_X1 u0_u4_u0_U62 (.A( u0_u4_X_4 ) , .ZN( u0_u4_u0_n159 ) );
  INV_X1 u0_u4_u0_U63 (.A( u0_u4_X_1 ) , .ZN( u0_u4_u0_n164 ) );
  INV_X1 u0_u4_u0_U64 (.A( u0_u4_X_2 ) , .ZN( u0_u4_u0_n163 ) );
  INV_X1 u0_u4_u0_U65 (.A( u0_u4_X_3 ) , .ZN( u0_u4_u0_n162 ) );
  INV_X1 u0_u4_u0_U66 (.A( u0_u4_u0_n126 ) , .ZN( u0_u4_u0_n168 ) );
  AOI211_X1 u0_u4_u0_U67 (.B( u0_u4_u0_n133 ) , .A( u0_u4_u0_n134 ) , .C2( u0_u4_u0_n135 ) , .C1( u0_u4_u0_n136 ) , .ZN( u0_u4_u0_n137 ) );
  OR4_X1 u0_u4_u0_U68 (.ZN( u0_out4_17 ) , .A4( u0_u4_u0_n122 ) , .A2( u0_u4_u0_n123 ) , .A1( u0_u4_u0_n124 ) , .A3( u0_u4_u0_n170 ) );
  AOI21_X1 u0_u4_u0_U69 (.B2( u0_u4_u0_n107 ) , .ZN( u0_u4_u0_n124 ) , .B1( u0_u4_u0_n128 ) , .A( u0_u4_u0_n161 ) );
  OAI21_X1 u0_u4_u0_U7 (.B1( u0_u4_u0_n150 ) , .B2( u0_u4_u0_n158 ) , .A( u0_u4_u0_n172 ) , .ZN( u0_u4_u0_n89 ) );
  INV_X1 u0_u4_u0_U70 (.A( u0_u4_u0_n111 ) , .ZN( u0_u4_u0_n170 ) );
  OR4_X1 u0_u4_u0_U71 (.ZN( u0_out4_31 ) , .A4( u0_u4_u0_n155 ) , .A2( u0_u4_u0_n156 ) , .A1( u0_u4_u0_n157 ) , .A3( u0_u4_u0_n173 ) );
  AOI21_X1 u0_u4_u0_U72 (.A( u0_u4_u0_n138 ) , .B2( u0_u4_u0_n139 ) , .B1( u0_u4_u0_n140 ) , .ZN( u0_u4_u0_n157 ) );
  AOI21_X1 u0_u4_u0_U73 (.B2( u0_u4_u0_n141 ) , .B1( u0_u4_u0_n142 ) , .ZN( u0_u4_u0_n156 ) , .A( u0_u4_u0_n161 ) );
  INV_X1 u0_u4_u0_U74 (.ZN( u0_u4_u0_n174 ) , .A( u0_u4_u0_n89 ) );
  AOI211_X1 u0_u4_u0_U75 (.B( u0_u4_u0_n104 ) , .A( u0_u4_u0_n105 ) , .ZN( u0_u4_u0_n106 ) , .C2( u0_u4_u0_n113 ) , .C1( u0_u4_u0_n160 ) );
  NOR2_X1 u0_u4_u0_U76 (.A2( u0_u4_X_3 ) , .A1( u0_u4_X_6 ) , .ZN( u0_u4_u0_n94 ) );
  NOR2_X1 u0_u4_u0_U77 (.A1( u0_u4_u0_n163 ) , .A2( u0_u4_u0_n164 ) , .ZN( u0_u4_u0_n95 ) );
  OAI221_X1 u0_u4_u0_U78 (.C1( u0_u4_u0_n121 ) , .ZN( u0_u4_u0_n122 ) , .B2( u0_u4_u0_n127 ) , .A( u0_u4_u0_n143 ) , .B1( u0_u4_u0_n144 ) , .C2( u0_u4_u0_n147 ) );
  NOR2_X1 u0_u4_u0_U79 (.A1( u0_u4_u0_n120 ) , .ZN( u0_u4_u0_n143 ) , .A2( u0_u4_u0_n167 ) );
  AND2_X1 u0_u4_u0_U8 (.A1( u0_u4_u0_n114 ) , .A2( u0_u4_u0_n121 ) , .ZN( u0_u4_u0_n146 ) );
  AOI21_X1 u0_u4_u0_U80 (.B1( u0_u4_u0_n132 ) , .ZN( u0_u4_u0_n133 ) , .A( u0_u4_u0_n144 ) , .B2( u0_u4_u0_n166 ) );
  OAI22_X1 u0_u4_u0_U81 (.ZN( u0_u4_u0_n105 ) , .A2( u0_u4_u0_n132 ) , .B1( u0_u4_u0_n146 ) , .A1( u0_u4_u0_n147 ) , .B2( u0_u4_u0_n161 ) );
  NAND2_X1 u0_u4_u0_U82 (.ZN( u0_u4_u0_n110 ) , .A2( u0_u4_u0_n132 ) , .A1( u0_u4_u0_n145 ) );
  INV_X1 u0_u4_u0_U83 (.A( u0_u4_u0_n119 ) , .ZN( u0_u4_u0_n167 ) );
  NAND2_X1 u0_u4_u0_U84 (.A2( u0_u4_u0_n103 ) , .ZN( u0_u4_u0_n140 ) , .A1( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U85 (.A1( u0_u4_u0_n101 ) , .ZN( u0_u4_u0_n130 ) , .A2( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U86 (.ZN( u0_u4_u0_n108 ) , .A1( u0_u4_u0_n92 ) , .A2( u0_u4_u0_n94 ) );
  NAND2_X1 u0_u4_u0_U87 (.ZN( u0_u4_u0_n142 ) , .A1( u0_u4_u0_n94 ) , .A2( u0_u4_u0_n95 ) );
  NAND3_X1 u0_u4_u0_U88 (.ZN( u0_out4_23 ) , .A3( u0_u4_u0_n137 ) , .A1( u0_u4_u0_n168 ) , .A2( u0_u4_u0_n171 ) );
  NAND3_X1 u0_u4_u0_U89 (.A3( u0_u4_u0_n127 ) , .A2( u0_u4_u0_n128 ) , .ZN( u0_u4_u0_n135 ) , .A1( u0_u4_u0_n150 ) );
  AND2_X1 u0_u4_u0_U9 (.A1( u0_u4_u0_n131 ) , .ZN( u0_u4_u0_n141 ) , .A2( u0_u4_u0_n150 ) );
  NAND3_X1 u0_u4_u0_U90 (.ZN( u0_u4_u0_n117 ) , .A3( u0_u4_u0_n132 ) , .A2( u0_u4_u0_n139 ) , .A1( u0_u4_u0_n148 ) );
  NAND3_X1 u0_u4_u0_U91 (.ZN( u0_u4_u0_n109 ) , .A2( u0_u4_u0_n114 ) , .A3( u0_u4_u0_n140 ) , .A1( u0_u4_u0_n149 ) );
  NAND3_X1 u0_u4_u0_U92 (.ZN( u0_out4_9 ) , .A3( u0_u4_u0_n106 ) , .A2( u0_u4_u0_n171 ) , .A1( u0_u4_u0_n174 ) );
  NAND3_X1 u0_u4_u0_U93 (.A2( u0_u4_u0_n128 ) , .A1( u0_u4_u0_n132 ) , .A3( u0_u4_u0_n146 ) , .ZN( u0_u4_u0_n97 ) );
  NOR2_X1 u0_u4_u5_U10 (.ZN( u0_u4_u5_n135 ) , .A1( u0_u4_u5_n173 ) , .A2( u0_u4_u5_n176 ) );
  NOR3_X1 u0_u4_u5_U100 (.A3( u0_u4_u5_n141 ) , .A1( u0_u4_u5_n142 ) , .ZN( u0_u4_u5_n143 ) , .A2( u0_u4_u5_n191 ) );
  NAND4_X1 u0_u4_u5_U101 (.ZN( u0_out4_4 ) , .A4( u0_u4_u5_n112 ) , .A2( u0_u4_u5_n113 ) , .A1( u0_u4_u5_n114 ) , .A3( u0_u4_u5_n195 ) );
  AOI211_X1 u0_u4_u5_U102 (.A( u0_u4_u5_n110 ) , .C1( u0_u4_u5_n111 ) , .ZN( u0_u4_u5_n112 ) , .B( u0_u4_u5_n118 ) , .C2( u0_u4_u5_n177 ) );
  INV_X1 u0_u4_u5_U103 (.A( u0_u4_u5_n102 ) , .ZN( u0_u4_u5_n195 ) );
  NAND3_X1 u0_u4_u5_U104 (.A2( u0_u4_u5_n154 ) , .A3( u0_u4_u5_n158 ) , .A1( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n99 ) );
  INV_X1 u0_u4_u5_U11 (.A( u0_u4_u5_n121 ) , .ZN( u0_u4_u5_n177 ) );
  NOR2_X1 u0_u4_u5_U12 (.ZN( u0_u4_u5_n160 ) , .A2( u0_u4_u5_n173 ) , .A1( u0_u4_u5_n177 ) );
  INV_X1 u0_u4_u5_U13 (.A( u0_u4_u5_n150 ) , .ZN( u0_u4_u5_n174 ) );
  AOI21_X1 u0_u4_u5_U14 (.A( u0_u4_u5_n160 ) , .B2( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n162 ) , .B1( u0_u4_u5_n192 ) );
  INV_X1 u0_u4_u5_U15 (.A( u0_u4_u5_n159 ) , .ZN( u0_u4_u5_n192 ) );
  AOI21_X1 u0_u4_u5_U16 (.A( u0_u4_u5_n156 ) , .B2( u0_u4_u5_n157 ) , .B1( u0_u4_u5_n158 ) , .ZN( u0_u4_u5_n163 ) );
  AOI21_X1 u0_u4_u5_U17 (.B2( u0_u4_u5_n139 ) , .B1( u0_u4_u5_n140 ) , .ZN( u0_u4_u5_n141 ) , .A( u0_u4_u5_n150 ) );
  OAI21_X1 u0_u4_u5_U18 (.A( u0_u4_u5_n133 ) , .B2( u0_u4_u5_n134 ) , .B1( u0_u4_u5_n135 ) , .ZN( u0_u4_u5_n142 ) );
  OAI21_X1 u0_u4_u5_U19 (.ZN( u0_u4_u5_n133 ) , .B2( u0_u4_u5_n147 ) , .A( u0_u4_u5_n173 ) , .B1( u0_u4_u5_n188 ) );
  NAND2_X1 u0_u4_u5_U20 (.A2( u0_u4_u5_n119 ) , .A1( u0_u4_u5_n123 ) , .ZN( u0_u4_u5_n137 ) );
  INV_X1 u0_u4_u5_U21 (.A( u0_u4_u5_n155 ) , .ZN( u0_u4_u5_n194 ) );
  NAND2_X1 u0_u4_u5_U22 (.A1( u0_u4_u5_n121 ) , .ZN( u0_u4_u5_n132 ) , .A2( u0_u4_u5_n172 ) );
  NAND2_X1 u0_u4_u5_U23 (.A2( u0_u4_u5_n122 ) , .ZN( u0_u4_u5_n136 ) , .A1( u0_u4_u5_n154 ) );
  NAND2_X1 u0_u4_u5_U24 (.A2( u0_u4_u5_n119 ) , .A1( u0_u4_u5_n120 ) , .ZN( u0_u4_u5_n159 ) );
  INV_X1 u0_u4_u5_U25 (.A( u0_u4_u5_n156 ) , .ZN( u0_u4_u5_n175 ) );
  INV_X1 u0_u4_u5_U26 (.A( u0_u4_u5_n158 ) , .ZN( u0_u4_u5_n188 ) );
  INV_X1 u0_u4_u5_U27 (.A( u0_u4_u5_n152 ) , .ZN( u0_u4_u5_n179 ) );
  INV_X1 u0_u4_u5_U28 (.A( u0_u4_u5_n140 ) , .ZN( u0_u4_u5_n182 ) );
  INV_X1 u0_u4_u5_U29 (.A( u0_u4_u5_n151 ) , .ZN( u0_u4_u5_n183 ) );
  NOR2_X1 u0_u4_u5_U3 (.ZN( u0_u4_u5_n134 ) , .A1( u0_u4_u5_n183 ) , .A2( u0_u4_u5_n190 ) );
  INV_X1 u0_u4_u5_U30 (.A( u0_u4_u5_n123 ) , .ZN( u0_u4_u5_n185 ) );
  INV_X1 u0_u4_u5_U31 (.A( u0_u4_u5_n161 ) , .ZN( u0_u4_u5_n184 ) );
  INV_X1 u0_u4_u5_U32 (.A( u0_u4_u5_n139 ) , .ZN( u0_u4_u5_n189 ) );
  INV_X1 u0_u4_u5_U33 (.A( u0_u4_u5_n157 ) , .ZN( u0_u4_u5_n190 ) );
  INV_X1 u0_u4_u5_U34 (.A( u0_u4_u5_n120 ) , .ZN( u0_u4_u5_n193 ) );
  NAND2_X1 u0_u4_u5_U35 (.ZN( u0_u4_u5_n111 ) , .A1( u0_u4_u5_n140 ) , .A2( u0_u4_u5_n155 ) );
  INV_X1 u0_u4_u5_U36 (.A( u0_u4_u5_n117 ) , .ZN( u0_u4_u5_n196 ) );
  OAI221_X1 u0_u4_u5_U37 (.A( u0_u4_u5_n116 ) , .ZN( u0_u4_u5_n117 ) , .B2( u0_u4_u5_n119 ) , .C1( u0_u4_u5_n153 ) , .C2( u0_u4_u5_n158 ) , .B1( u0_u4_u5_n172 ) );
  AOI222_X1 u0_u4_u5_U38 (.ZN( u0_u4_u5_n116 ) , .B2( u0_u4_u5_n145 ) , .C1( u0_u4_u5_n148 ) , .A2( u0_u4_u5_n174 ) , .C2( u0_u4_u5_n177 ) , .B1( u0_u4_u5_n187 ) , .A1( u0_u4_u5_n193 ) );
  INV_X1 u0_u4_u5_U39 (.A( u0_u4_u5_n115 ) , .ZN( u0_u4_u5_n187 ) );
  INV_X1 u0_u4_u5_U4 (.A( u0_u4_u5_n138 ) , .ZN( u0_u4_u5_n191 ) );
  NOR2_X1 u0_u4_u5_U40 (.ZN( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n170 ) , .A2( u0_u4_u5_n180 ) );
  OAI221_X1 u0_u4_u5_U41 (.A( u0_u4_u5_n101 ) , .ZN( u0_u4_u5_n102 ) , .C2( u0_u4_u5_n115 ) , .C1( u0_u4_u5_n126 ) , .B1( u0_u4_u5_n134 ) , .B2( u0_u4_u5_n160 ) );
  OAI21_X1 u0_u4_u5_U42 (.ZN( u0_u4_u5_n101 ) , .B1( u0_u4_u5_n137 ) , .A( u0_u4_u5_n146 ) , .B2( u0_u4_u5_n147 ) );
  AOI22_X1 u0_u4_u5_U43 (.B2( u0_u4_u5_n131 ) , .A2( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n169 ) , .B1( u0_u4_u5_n174 ) , .A1( u0_u4_u5_n185 ) );
  NOR2_X1 u0_u4_u5_U44 (.A1( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n150 ) , .A2( u0_u4_u5_n173 ) );
  AOI21_X1 u0_u4_u5_U45 (.A( u0_u4_u5_n118 ) , .B2( u0_u4_u5_n145 ) , .ZN( u0_u4_u5_n168 ) , .B1( u0_u4_u5_n186 ) );
  INV_X1 u0_u4_u5_U46 (.A( u0_u4_u5_n122 ) , .ZN( u0_u4_u5_n186 ) );
  NOR2_X1 u0_u4_u5_U47 (.A1( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n152 ) , .A2( u0_u4_u5_n176 ) );
  NOR2_X1 u0_u4_u5_U48 (.A1( u0_u4_u5_n115 ) , .ZN( u0_u4_u5_n118 ) , .A2( u0_u4_u5_n153 ) );
  NOR2_X1 u0_u4_u5_U49 (.A2( u0_u4_u5_n145 ) , .ZN( u0_u4_u5_n156 ) , .A1( u0_u4_u5_n174 ) );
  OAI21_X1 u0_u4_u5_U5 (.B2( u0_u4_u5_n136 ) , .B1( u0_u4_u5_n137 ) , .ZN( u0_u4_u5_n138 ) , .A( u0_u4_u5_n177 ) );
  NOR2_X1 u0_u4_u5_U50 (.ZN( u0_u4_u5_n121 ) , .A2( u0_u4_u5_n145 ) , .A1( u0_u4_u5_n176 ) );
  AOI22_X1 u0_u4_u5_U51 (.ZN( u0_u4_u5_n114 ) , .A2( u0_u4_u5_n137 ) , .A1( u0_u4_u5_n145 ) , .B2( u0_u4_u5_n175 ) , .B1( u0_u4_u5_n193 ) );
  OAI211_X1 u0_u4_u5_U52 (.B( u0_u4_u5_n124 ) , .A( u0_u4_u5_n125 ) , .C2( u0_u4_u5_n126 ) , .C1( u0_u4_u5_n127 ) , .ZN( u0_u4_u5_n128 ) );
  NOR3_X1 u0_u4_u5_U53 (.ZN( u0_u4_u5_n127 ) , .A1( u0_u4_u5_n136 ) , .A3( u0_u4_u5_n148 ) , .A2( u0_u4_u5_n182 ) );
  OAI21_X1 u0_u4_u5_U54 (.ZN( u0_u4_u5_n124 ) , .A( u0_u4_u5_n177 ) , .B2( u0_u4_u5_n183 ) , .B1( u0_u4_u5_n189 ) );
  OAI21_X1 u0_u4_u5_U55 (.ZN( u0_u4_u5_n125 ) , .A( u0_u4_u5_n174 ) , .B2( u0_u4_u5_n185 ) , .B1( u0_u4_u5_n190 ) );
  AOI21_X1 u0_u4_u5_U56 (.A( u0_u4_u5_n153 ) , .B2( u0_u4_u5_n154 ) , .B1( u0_u4_u5_n155 ) , .ZN( u0_u4_u5_n164 ) );
  AOI21_X1 u0_u4_u5_U57 (.ZN( u0_u4_u5_n110 ) , .B1( u0_u4_u5_n122 ) , .B2( u0_u4_u5_n139 ) , .A( u0_u4_u5_n153 ) );
  INV_X1 u0_u4_u5_U58 (.A( u0_u4_u5_n153 ) , .ZN( u0_u4_u5_n176 ) );
  INV_X1 u0_u4_u5_U59 (.A( u0_u4_u5_n126 ) , .ZN( u0_u4_u5_n173 ) );
  AOI222_X1 u0_u4_u5_U6 (.ZN( u0_u4_u5_n113 ) , .A1( u0_u4_u5_n131 ) , .C1( u0_u4_u5_n148 ) , .B2( u0_u4_u5_n174 ) , .C2( u0_u4_u5_n178 ) , .A2( u0_u4_u5_n179 ) , .B1( u0_u4_u5_n99 ) );
  AND2_X1 u0_u4_u5_U60 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n147 ) );
  AND2_X1 u0_u4_u5_U61 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n148 ) );
  NAND2_X1 u0_u4_u5_U62 (.A1( u0_u4_u5_n105 ) , .A2( u0_u4_u5_n106 ) , .ZN( u0_u4_u5_n158 ) );
  NAND2_X1 u0_u4_u5_U63 (.A2( u0_u4_u5_n108 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n139 ) );
  NAND2_X1 u0_u4_u5_U64 (.A1( u0_u4_u5_n106 ) , .A2( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n119 ) );
  NAND2_X1 u0_u4_u5_U65 (.A2( u0_u4_u5_n103 ) , .A1( u0_u4_u5_n105 ) , .ZN( u0_u4_u5_n140 ) );
  NAND2_X1 u0_u4_u5_U66 (.A2( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n105 ) , .ZN( u0_u4_u5_n155 ) );
  NAND2_X1 u0_u4_u5_U67 (.A2( u0_u4_u5_n106 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n122 ) );
  NAND2_X1 u0_u4_u5_U68 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n106 ) , .ZN( u0_u4_u5_n115 ) );
  NAND2_X1 u0_u4_u5_U69 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n103 ) , .ZN( u0_u4_u5_n161 ) );
  INV_X1 u0_u4_u5_U7 (.A( u0_u4_u5_n135 ) , .ZN( u0_u4_u5_n178 ) );
  NAND2_X1 u0_u4_u5_U70 (.A1( u0_u4_u5_n105 ) , .A2( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n154 ) );
  INV_X1 u0_u4_u5_U71 (.A( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n172 ) );
  NAND2_X1 u0_u4_u5_U72 (.A1( u0_u4_u5_n103 ) , .A2( u0_u4_u5_n108 ) , .ZN( u0_u4_u5_n123 ) );
  NAND2_X1 u0_u4_u5_U73 (.A2( u0_u4_u5_n103 ) , .A1( u0_u4_u5_n107 ) , .ZN( u0_u4_u5_n151 ) );
  NAND2_X1 u0_u4_u5_U74 (.A2( u0_u4_u5_n107 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n120 ) );
  NAND2_X1 u0_u4_u5_U75 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n109 ) , .ZN( u0_u4_u5_n157 ) );
  AND2_X1 u0_u4_u5_U76 (.A2( u0_u4_u5_n100 ) , .A1( u0_u4_u5_n104 ) , .ZN( u0_u4_u5_n131 ) );
  NOR2_X1 u0_u4_u5_U77 (.A2( u0_u4_X_34 ) , .A1( u0_u4_X_35 ) , .ZN( u0_u4_u5_n145 ) );
  NOR2_X1 u0_u4_u5_U78 (.A2( u0_u4_X_34 ) , .ZN( u0_u4_u5_n146 ) , .A1( u0_u4_u5_n171 ) );
  NOR2_X1 u0_u4_u5_U79 (.A2( u0_u4_X_31 ) , .A1( u0_u4_X_32 ) , .ZN( u0_u4_u5_n103 ) );
  OAI22_X1 u0_u4_u5_U8 (.B2( u0_u4_u5_n149 ) , .B1( u0_u4_u5_n150 ) , .A2( u0_u4_u5_n151 ) , .A1( u0_u4_u5_n152 ) , .ZN( u0_u4_u5_n165 ) );
  NOR2_X1 u0_u4_u5_U80 (.A2( u0_u4_X_36 ) , .ZN( u0_u4_u5_n105 ) , .A1( u0_u4_u5_n180 ) );
  NOR2_X1 u0_u4_u5_U81 (.A2( u0_u4_X_33 ) , .ZN( u0_u4_u5_n108 ) , .A1( u0_u4_u5_n170 ) );
  NOR2_X1 u0_u4_u5_U82 (.A2( u0_u4_X_33 ) , .A1( u0_u4_X_36 ) , .ZN( u0_u4_u5_n107 ) );
  NOR2_X1 u0_u4_u5_U83 (.A2( u0_u4_X_31 ) , .ZN( u0_u4_u5_n104 ) , .A1( u0_u4_u5_n181 ) );
  NAND2_X1 u0_u4_u5_U84 (.A2( u0_u4_X_34 ) , .A1( u0_u4_X_35 ) , .ZN( u0_u4_u5_n153 ) );
  NAND2_X1 u0_u4_u5_U85 (.A1( u0_u4_X_34 ) , .ZN( u0_u4_u5_n126 ) , .A2( u0_u4_u5_n171 ) );
  AND2_X1 u0_u4_u5_U86 (.A1( u0_u4_X_31 ) , .A2( u0_u4_X_32 ) , .ZN( u0_u4_u5_n106 ) );
  AND2_X1 u0_u4_u5_U87 (.A1( u0_u4_X_31 ) , .ZN( u0_u4_u5_n109 ) , .A2( u0_u4_u5_n181 ) );
  INV_X1 u0_u4_u5_U88 (.A( u0_u4_X_33 ) , .ZN( u0_u4_u5_n180 ) );
  INV_X1 u0_u4_u5_U89 (.A( u0_u4_X_35 ) , .ZN( u0_u4_u5_n171 ) );
  NOR3_X1 u0_u4_u5_U9 (.A2( u0_u4_u5_n147 ) , .A1( u0_u4_u5_n148 ) , .ZN( u0_u4_u5_n149 ) , .A3( u0_u4_u5_n194 ) );
  INV_X1 u0_u4_u5_U90 (.A( u0_u4_X_36 ) , .ZN( u0_u4_u5_n170 ) );
  INV_X1 u0_u4_u5_U91 (.A( u0_u4_X_32 ) , .ZN( u0_u4_u5_n181 ) );
  NAND4_X1 u0_u4_u5_U92 (.ZN( u0_out4_29 ) , .A4( u0_u4_u5_n129 ) , .A3( u0_u4_u5_n130 ) , .A2( u0_u4_u5_n168 ) , .A1( u0_u4_u5_n196 ) );
  AOI221_X1 u0_u4_u5_U93 (.A( u0_u4_u5_n128 ) , .ZN( u0_u4_u5_n129 ) , .C2( u0_u4_u5_n132 ) , .B2( u0_u4_u5_n159 ) , .B1( u0_u4_u5_n176 ) , .C1( u0_u4_u5_n184 ) );
  AOI222_X1 u0_u4_u5_U94 (.ZN( u0_u4_u5_n130 ) , .A2( u0_u4_u5_n146 ) , .B1( u0_u4_u5_n147 ) , .C2( u0_u4_u5_n175 ) , .B2( u0_u4_u5_n179 ) , .A1( u0_u4_u5_n188 ) , .C1( u0_u4_u5_n194 ) );
  NAND4_X1 u0_u4_u5_U95 (.ZN( u0_out4_19 ) , .A4( u0_u4_u5_n166 ) , .A3( u0_u4_u5_n167 ) , .A2( u0_u4_u5_n168 ) , .A1( u0_u4_u5_n169 ) );
  AOI22_X1 u0_u4_u5_U96 (.B2( u0_u4_u5_n145 ) , .A2( u0_u4_u5_n146 ) , .ZN( u0_u4_u5_n167 ) , .B1( u0_u4_u5_n182 ) , .A1( u0_u4_u5_n189 ) );
  NOR4_X1 u0_u4_u5_U97 (.A4( u0_u4_u5_n162 ) , .A3( u0_u4_u5_n163 ) , .A2( u0_u4_u5_n164 ) , .A1( u0_u4_u5_n165 ) , .ZN( u0_u4_u5_n166 ) );
  NAND4_X1 u0_u4_u5_U98 (.ZN( u0_out4_11 ) , .A4( u0_u4_u5_n143 ) , .A3( u0_u4_u5_n144 ) , .A2( u0_u4_u5_n169 ) , .A1( u0_u4_u5_n196 ) );
  AOI22_X1 u0_u4_u5_U99 (.A2( u0_u4_u5_n132 ) , .ZN( u0_u4_u5_n144 ) , .B2( u0_u4_u5_n145 ) , .B1( u0_u4_u5_n184 ) , .A1( u0_u4_u5_n194 ) );
  AOI22_X1 u0_u4_u6_U10 (.A2( u0_u4_u6_n151 ) , .B2( u0_u4_u6_n161 ) , .A1( u0_u4_u6_n167 ) , .B1( u0_u4_u6_n170 ) , .ZN( u0_u4_u6_n89 ) );
  AOI21_X1 u0_u4_u6_U11 (.B1( u0_u4_u6_n107 ) , .B2( u0_u4_u6_n132 ) , .A( u0_u4_u6_n158 ) , .ZN( u0_u4_u6_n88 ) );
  AOI21_X1 u0_u4_u6_U12 (.B2( u0_u4_u6_n147 ) , .B1( u0_u4_u6_n148 ) , .ZN( u0_u4_u6_n149 ) , .A( u0_u4_u6_n158 ) );
  AOI21_X1 u0_u4_u6_U13 (.ZN( u0_u4_u6_n106 ) , .A( u0_u4_u6_n142 ) , .B2( u0_u4_u6_n159 ) , .B1( u0_u4_u6_n164 ) );
  INV_X1 u0_u4_u6_U14 (.A( u0_u4_u6_n155 ) , .ZN( u0_u4_u6_n161 ) );
  INV_X1 u0_u4_u6_U15 (.A( u0_u4_u6_n128 ) , .ZN( u0_u4_u6_n164 ) );
  NAND2_X1 u0_u4_u6_U16 (.ZN( u0_u4_u6_n110 ) , .A1( u0_u4_u6_n122 ) , .A2( u0_u4_u6_n129 ) );
  NAND2_X1 u0_u4_u6_U17 (.ZN( u0_u4_u6_n124 ) , .A2( u0_u4_u6_n146 ) , .A1( u0_u4_u6_n148 ) );
  INV_X1 u0_u4_u6_U18 (.A( u0_u4_u6_n132 ) , .ZN( u0_u4_u6_n171 ) );
  AND2_X1 u0_u4_u6_U19 (.A1( u0_u4_u6_n100 ) , .ZN( u0_u4_u6_n130 ) , .A2( u0_u4_u6_n147 ) );
  INV_X1 u0_u4_u6_U20 (.A( u0_u4_u6_n127 ) , .ZN( u0_u4_u6_n173 ) );
  INV_X1 u0_u4_u6_U21 (.A( u0_u4_u6_n121 ) , .ZN( u0_u4_u6_n167 ) );
  INV_X1 u0_u4_u6_U22 (.A( u0_u4_u6_n100 ) , .ZN( u0_u4_u6_n169 ) );
  INV_X1 u0_u4_u6_U23 (.A( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n170 ) );
  INV_X1 u0_u4_u6_U24 (.A( u0_u4_u6_n113 ) , .ZN( u0_u4_u6_n168 ) );
  AND2_X1 u0_u4_u6_U25 (.A1( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n119 ) , .ZN( u0_u4_u6_n133 ) );
  AND2_X1 u0_u4_u6_U26 (.A2( u0_u4_u6_n121 ) , .A1( u0_u4_u6_n122 ) , .ZN( u0_u4_u6_n131 ) );
  AND3_X1 u0_u4_u6_U27 (.ZN( u0_u4_u6_n120 ) , .A2( u0_u4_u6_n127 ) , .A1( u0_u4_u6_n132 ) , .A3( u0_u4_u6_n145 ) );
  INV_X1 u0_u4_u6_U28 (.A( u0_u4_u6_n146 ) , .ZN( u0_u4_u6_n163 ) );
  AOI222_X1 u0_u4_u6_U29 (.ZN( u0_u4_u6_n114 ) , .A1( u0_u4_u6_n118 ) , .A2( u0_u4_u6_n126 ) , .B2( u0_u4_u6_n151 ) , .C2( u0_u4_u6_n159 ) , .C1( u0_u4_u6_n168 ) , .B1( u0_u4_u6_n169 ) );
  INV_X1 u0_u4_u6_U3 (.A( u0_u4_u6_n110 ) , .ZN( u0_u4_u6_n166 ) );
  NOR2_X1 u0_u4_u6_U30 (.A1( u0_u4_u6_n162 ) , .A2( u0_u4_u6_n165 ) , .ZN( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U31 (.A1( u0_u4_u6_n144 ) , .ZN( u0_u4_u6_n151 ) , .A2( u0_u4_u6_n158 ) );
  NAND2_X1 u0_u4_u6_U32 (.ZN( u0_u4_u6_n132 ) , .A1( u0_u4_u6_n91 ) , .A2( u0_u4_u6_n97 ) );
  AOI22_X1 u0_u4_u6_U33 (.B2( u0_u4_u6_n110 ) , .B1( u0_u4_u6_n111 ) , .A1( u0_u4_u6_n112 ) , .ZN( u0_u4_u6_n115 ) , .A2( u0_u4_u6_n161 ) );
  NAND4_X1 u0_u4_u6_U34 (.A3( u0_u4_u6_n109 ) , .ZN( u0_u4_u6_n112 ) , .A4( u0_u4_u6_n132 ) , .A2( u0_u4_u6_n147 ) , .A1( u0_u4_u6_n166 ) );
  NOR2_X1 u0_u4_u6_U35 (.ZN( u0_u4_u6_n109 ) , .A1( u0_u4_u6_n170 ) , .A2( u0_u4_u6_n173 ) );
  NOR2_X1 u0_u4_u6_U36 (.A2( u0_u4_u6_n126 ) , .ZN( u0_u4_u6_n155 ) , .A1( u0_u4_u6_n160 ) );
  NAND2_X1 u0_u4_u6_U37 (.ZN( u0_u4_u6_n146 ) , .A2( u0_u4_u6_n94 ) , .A1( u0_u4_u6_n99 ) );
  AOI21_X1 u0_u4_u6_U38 (.A( u0_u4_u6_n144 ) , .B2( u0_u4_u6_n145 ) , .B1( u0_u4_u6_n146 ) , .ZN( u0_u4_u6_n150 ) );
  AOI211_X1 u0_u4_u6_U39 (.B( u0_u4_u6_n134 ) , .A( u0_u4_u6_n135 ) , .C1( u0_u4_u6_n136 ) , .ZN( u0_u4_u6_n137 ) , .C2( u0_u4_u6_n151 ) );
  INV_X1 u0_u4_u6_U4 (.A( u0_u4_u6_n142 ) , .ZN( u0_u4_u6_n174 ) );
  NAND4_X1 u0_u4_u6_U40 (.A4( u0_u4_u6_n127 ) , .A3( u0_u4_u6_n128 ) , .A2( u0_u4_u6_n129 ) , .A1( u0_u4_u6_n130 ) , .ZN( u0_u4_u6_n136 ) );
  AOI21_X1 u0_u4_u6_U41 (.B2( u0_u4_u6_n132 ) , .B1( u0_u4_u6_n133 ) , .ZN( u0_u4_u6_n134 ) , .A( u0_u4_u6_n158 ) );
  AOI21_X1 u0_u4_u6_U42 (.B1( u0_u4_u6_n131 ) , .ZN( u0_u4_u6_n135 ) , .A( u0_u4_u6_n144 ) , .B2( u0_u4_u6_n146 ) );
  INV_X1 u0_u4_u6_U43 (.A( u0_u4_u6_n111 ) , .ZN( u0_u4_u6_n158 ) );
  NAND2_X1 u0_u4_u6_U44 (.ZN( u0_u4_u6_n127 ) , .A1( u0_u4_u6_n91 ) , .A2( u0_u4_u6_n92 ) );
  NAND2_X1 u0_u4_u6_U45 (.ZN( u0_u4_u6_n129 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n96 ) );
  INV_X1 u0_u4_u6_U46 (.A( u0_u4_u6_n144 ) , .ZN( u0_u4_u6_n159 ) );
  NAND2_X1 u0_u4_u6_U47 (.ZN( u0_u4_u6_n145 ) , .A2( u0_u4_u6_n97 ) , .A1( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U48 (.ZN( u0_u4_u6_n148 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n94 ) );
  NAND2_X1 u0_u4_u6_U49 (.ZN( u0_u4_u6_n108 ) , .A2( u0_u4_u6_n139 ) , .A1( u0_u4_u6_n144 ) );
  NAND2_X1 u0_u4_u6_U5 (.A2( u0_u4_u6_n143 ) , .ZN( u0_u4_u6_n152 ) , .A1( u0_u4_u6_n166 ) );
  NAND2_X1 u0_u4_u6_U50 (.ZN( u0_u4_u6_n121 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n97 ) );
  NAND2_X1 u0_u4_u6_U51 (.ZN( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n95 ) );
  AND2_X1 u0_u4_u6_U52 (.ZN( u0_u4_u6_n118 ) , .A2( u0_u4_u6_n91 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U53 (.ZN( u0_u4_u6_n147 ) , .A2( u0_u4_u6_n98 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U54 (.ZN( u0_u4_u6_n128 ) , .A1( u0_u4_u6_n94 ) , .A2( u0_u4_u6_n96 ) );
  NAND2_X1 u0_u4_u6_U55 (.ZN( u0_u4_u6_n119 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U56 (.ZN( u0_u4_u6_n123 ) , .A2( u0_u4_u6_n91 ) , .A1( u0_u4_u6_n96 ) );
  NAND2_X1 u0_u4_u6_U57 (.ZN( u0_u4_u6_n100 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U58 (.ZN( u0_u4_u6_n122 ) , .A1( u0_u4_u6_n94 ) , .A2( u0_u4_u6_n97 ) );
  INV_X1 u0_u4_u6_U59 (.A( u0_u4_u6_n139 ) , .ZN( u0_u4_u6_n160 ) );
  AOI22_X1 u0_u4_u6_U6 (.B2( u0_u4_u6_n101 ) , .A1( u0_u4_u6_n102 ) , .ZN( u0_u4_u6_n103 ) , .B1( u0_u4_u6_n160 ) , .A2( u0_u4_u6_n161 ) );
  NAND2_X1 u0_u4_u6_U60 (.ZN( u0_u4_u6_n113 ) , .A1( u0_u4_u6_n96 ) , .A2( u0_u4_u6_n98 ) );
  NOR2_X1 u0_u4_u6_U61 (.A2( u0_u4_X_40 ) , .A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n126 ) );
  NOR2_X1 u0_u4_u6_U62 (.A2( u0_u4_X_39 ) , .A1( u0_u4_X_42 ) , .ZN( u0_u4_u6_n92 ) );
  NOR2_X1 u0_u4_u6_U63 (.A2( u0_u4_X_39 ) , .A1( u0_u4_u6_n156 ) , .ZN( u0_u4_u6_n97 ) );
  NOR2_X1 u0_u4_u6_U64 (.A2( u0_u4_X_38 ) , .A1( u0_u4_u6_n165 ) , .ZN( u0_u4_u6_n95 ) );
  NOR2_X1 u0_u4_u6_U65 (.A2( u0_u4_X_41 ) , .ZN( u0_u4_u6_n111 ) , .A1( u0_u4_u6_n157 ) );
  NOR2_X1 u0_u4_u6_U66 (.A2( u0_u4_X_37 ) , .A1( u0_u4_u6_n162 ) , .ZN( u0_u4_u6_n94 ) );
  NOR2_X1 u0_u4_u6_U67 (.A2( u0_u4_X_37 ) , .A1( u0_u4_X_38 ) , .ZN( u0_u4_u6_n91 ) );
  NAND2_X1 u0_u4_u6_U68 (.A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n144 ) , .A2( u0_u4_u6_n157 ) );
  NAND2_X1 u0_u4_u6_U69 (.A2( u0_u4_X_40 ) , .A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n139 ) );
  NOR2_X1 u0_u4_u6_U7 (.A1( u0_u4_u6_n118 ) , .ZN( u0_u4_u6_n143 ) , .A2( u0_u4_u6_n168 ) );
  AND2_X1 u0_u4_u6_U70 (.A1( u0_u4_X_39 ) , .A2( u0_u4_u6_n156 ) , .ZN( u0_u4_u6_n96 ) );
  AND2_X1 u0_u4_u6_U71 (.A1( u0_u4_X_39 ) , .A2( u0_u4_X_42 ) , .ZN( u0_u4_u6_n99 ) );
  INV_X1 u0_u4_u6_U72 (.A( u0_u4_X_40 ) , .ZN( u0_u4_u6_n157 ) );
  INV_X1 u0_u4_u6_U73 (.A( u0_u4_X_37 ) , .ZN( u0_u4_u6_n165 ) );
  INV_X1 u0_u4_u6_U74 (.A( u0_u4_X_38 ) , .ZN( u0_u4_u6_n162 ) );
  INV_X1 u0_u4_u6_U75 (.A( u0_u4_X_42 ) , .ZN( u0_u4_u6_n156 ) );
  NAND4_X1 u0_u4_u6_U76 (.ZN( u0_out4_32 ) , .A4( u0_u4_u6_n103 ) , .A3( u0_u4_u6_n104 ) , .A2( u0_u4_u6_n105 ) , .A1( u0_u4_u6_n106 ) );
  AOI22_X1 u0_u4_u6_U77 (.ZN( u0_u4_u6_n105 ) , .A2( u0_u4_u6_n108 ) , .A1( u0_u4_u6_n118 ) , .B2( u0_u4_u6_n126 ) , .B1( u0_u4_u6_n171 ) );
  AOI22_X1 u0_u4_u6_U78 (.ZN( u0_u4_u6_n104 ) , .A1( u0_u4_u6_n111 ) , .B1( u0_u4_u6_n124 ) , .B2( u0_u4_u6_n151 ) , .A2( u0_u4_u6_n93 ) );
  NAND4_X1 u0_u4_u6_U79 (.ZN( u0_out4_12 ) , .A4( u0_u4_u6_n114 ) , .A3( u0_u4_u6_n115 ) , .A2( u0_u4_u6_n116 ) , .A1( u0_u4_u6_n117 ) );
  INV_X1 u0_u4_u6_U8 (.ZN( u0_u4_u6_n172 ) , .A( u0_u4_u6_n88 ) );
  OAI22_X1 u0_u4_u6_U80 (.B2( u0_u4_u6_n111 ) , .ZN( u0_u4_u6_n116 ) , .B1( u0_u4_u6_n126 ) , .A2( u0_u4_u6_n164 ) , .A1( u0_u4_u6_n167 ) );
  OAI21_X1 u0_u4_u6_U81 (.A( u0_u4_u6_n108 ) , .ZN( u0_u4_u6_n117 ) , .B2( u0_u4_u6_n141 ) , .B1( u0_u4_u6_n163 ) );
  OAI211_X1 u0_u4_u6_U82 (.ZN( u0_out4_22 ) , .B( u0_u4_u6_n137 ) , .A( u0_u4_u6_n138 ) , .C2( u0_u4_u6_n139 ) , .C1( u0_u4_u6_n140 ) );
  AOI22_X1 u0_u4_u6_U83 (.B1( u0_u4_u6_n124 ) , .A2( u0_u4_u6_n125 ) , .A1( u0_u4_u6_n126 ) , .ZN( u0_u4_u6_n138 ) , .B2( u0_u4_u6_n161 ) );
  AND4_X1 u0_u4_u6_U84 (.A3( u0_u4_u6_n119 ) , .A1( u0_u4_u6_n120 ) , .A4( u0_u4_u6_n129 ) , .ZN( u0_u4_u6_n140 ) , .A2( u0_u4_u6_n143 ) );
  OAI211_X1 u0_u4_u6_U85 (.ZN( u0_out4_7 ) , .B( u0_u4_u6_n153 ) , .C2( u0_u4_u6_n154 ) , .C1( u0_u4_u6_n155 ) , .A( u0_u4_u6_n174 ) );
  NOR3_X1 u0_u4_u6_U86 (.A1( u0_u4_u6_n141 ) , .ZN( u0_u4_u6_n154 ) , .A3( u0_u4_u6_n164 ) , .A2( u0_u4_u6_n171 ) );
  AOI211_X1 u0_u4_u6_U87 (.B( u0_u4_u6_n149 ) , .A( u0_u4_u6_n150 ) , .C2( u0_u4_u6_n151 ) , .C1( u0_u4_u6_n152 ) , .ZN( u0_u4_u6_n153 ) );
  NAND3_X1 u0_u4_u6_U88 (.A2( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n125 ) , .A1( u0_u4_u6_n130 ) , .A3( u0_u4_u6_n131 ) );
  NAND3_X1 u0_u4_u6_U89 (.A3( u0_u4_u6_n133 ) , .ZN( u0_u4_u6_n141 ) , .A1( u0_u4_u6_n145 ) , .A2( u0_u4_u6_n148 ) );
  OAI21_X1 u0_u4_u6_U9 (.A( u0_u4_u6_n159 ) , .B1( u0_u4_u6_n169 ) , .B2( u0_u4_u6_n173 ) , .ZN( u0_u4_u6_n90 ) );
  NAND3_X1 u0_u4_u6_U90 (.ZN( u0_u4_u6_n101 ) , .A3( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n121 ) , .A1( u0_u4_u6_n127 ) );
  NAND3_X1 u0_u4_u6_U91 (.ZN( u0_u4_u6_n102 ) , .A3( u0_u4_u6_n130 ) , .A2( u0_u4_u6_n145 ) , .A1( u0_u4_u6_n166 ) );
  NAND3_X1 u0_u4_u6_U92 (.A3( u0_u4_u6_n113 ) , .A1( u0_u4_u6_n119 ) , .A2( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n93 ) );
  NAND3_X1 u0_u4_u6_U93 (.ZN( u0_u4_u6_n142 ) , .A2( u0_u4_u6_n172 ) , .A3( u0_u4_u6_n89 ) , .A1( u0_u4_u6_n90 ) );
  OAI21_X1 u0_u4_u7_U10 (.A( u0_u4_u7_n161 ) , .B1( u0_u4_u7_n168 ) , .B2( u0_u4_u7_n173 ) , .ZN( u0_u4_u7_n91 ) );
  AOI211_X1 u0_u4_u7_U11 (.A( u0_u4_u7_n117 ) , .ZN( u0_u4_u7_n118 ) , .C2( u0_u4_u7_n126 ) , .C1( u0_u4_u7_n177 ) , .B( u0_u4_u7_n180 ) );
  OAI22_X1 u0_u4_u7_U12 (.B1( u0_u4_u7_n115 ) , .ZN( u0_u4_u7_n117 ) , .A2( u0_u4_u7_n133 ) , .A1( u0_u4_u7_n137 ) , .B2( u0_u4_u7_n162 ) );
  INV_X1 u0_u4_u7_U13 (.A( u0_u4_u7_n116 ) , .ZN( u0_u4_u7_n180 ) );
  NOR3_X1 u0_u4_u7_U14 (.ZN( u0_u4_u7_n115 ) , .A3( u0_u4_u7_n145 ) , .A2( u0_u4_u7_n168 ) , .A1( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U15 (.A( u0_u4_u7_n133 ) , .ZN( u0_u4_u7_n176 ) );
  NOR3_X1 u0_u4_u7_U16 (.A2( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n135 ) , .ZN( u0_u4_u7_n136 ) , .A3( u0_u4_u7_n171 ) );
  NOR2_X1 u0_u4_u7_U17 (.A1( u0_u4_u7_n130 ) , .A2( u0_u4_u7_n134 ) , .ZN( u0_u4_u7_n153 ) );
  AOI21_X1 u0_u4_u7_U18 (.ZN( u0_u4_u7_n104 ) , .B2( u0_u4_u7_n112 ) , .B1( u0_u4_u7_n127 ) , .A( u0_u4_u7_n164 ) );
  AOI21_X1 u0_u4_u7_U19 (.ZN( u0_u4_u7_n106 ) , .B1( u0_u4_u7_n133 ) , .B2( u0_u4_u7_n146 ) , .A( u0_u4_u7_n162 ) );
  AOI21_X1 u0_u4_u7_U20 (.A( u0_u4_u7_n101 ) , .ZN( u0_u4_u7_n107 ) , .B2( u0_u4_u7_n128 ) , .B1( u0_u4_u7_n175 ) );
  INV_X1 u0_u4_u7_U21 (.A( u0_u4_u7_n101 ) , .ZN( u0_u4_u7_n165 ) );
  NOR2_X1 u0_u4_u7_U22 (.ZN( u0_u4_u7_n111 ) , .A2( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U23 (.A( u0_u4_u7_n138 ) , .ZN( u0_u4_u7_n171 ) );
  INV_X1 u0_u4_u7_U24 (.A( u0_u4_u7_n131 ) , .ZN( u0_u4_u7_n177 ) );
  INV_X1 u0_u4_u7_U25 (.A( u0_u4_u7_n110 ) , .ZN( u0_u4_u7_n174 ) );
  NAND2_X1 u0_u4_u7_U26 (.A1( u0_u4_u7_n129 ) , .A2( u0_u4_u7_n132 ) , .ZN( u0_u4_u7_n149 ) );
  NAND2_X1 u0_u4_u7_U27 (.A1( u0_u4_u7_n113 ) , .A2( u0_u4_u7_n124 ) , .ZN( u0_u4_u7_n130 ) );
  INV_X1 u0_u4_u7_U28 (.A( u0_u4_u7_n112 ) , .ZN( u0_u4_u7_n173 ) );
  INV_X1 u0_u4_u7_U29 (.A( u0_u4_u7_n128 ) , .ZN( u0_u4_u7_n168 ) );
  OAI21_X1 u0_u4_u7_U3 (.ZN( u0_u4_u7_n159 ) , .A( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n171 ) , .B1( u0_u4_u7_n174 ) );
  INV_X1 u0_u4_u7_U30 (.A( u0_u4_u7_n148 ) , .ZN( u0_u4_u7_n169 ) );
  INV_X1 u0_u4_u7_U31 (.A( u0_u4_u7_n127 ) , .ZN( u0_u4_u7_n179 ) );
  NOR2_X1 u0_u4_u7_U32 (.ZN( u0_u4_u7_n101 ) , .A2( u0_u4_u7_n150 ) , .A1( u0_u4_u7_n156 ) );
  AOI211_X1 u0_u4_u7_U33 (.B( u0_u4_u7_n139 ) , .A( u0_u4_u7_n140 ) , .C2( u0_u4_u7_n141 ) , .ZN( u0_u4_u7_n142 ) , .C1( u0_u4_u7_n156 ) );
  AOI21_X1 u0_u4_u7_U34 (.A( u0_u4_u7_n137 ) , .B1( u0_u4_u7_n138 ) , .ZN( u0_u4_u7_n139 ) , .B2( u0_u4_u7_n146 ) );
  NAND4_X1 u0_u4_u7_U35 (.A3( u0_u4_u7_n127 ) , .A2( u0_u4_u7_n128 ) , .A1( u0_u4_u7_n129 ) , .ZN( u0_u4_u7_n141 ) , .A4( u0_u4_u7_n147 ) );
  OAI22_X1 u0_u4_u7_U36 (.B1( u0_u4_u7_n136 ) , .ZN( u0_u4_u7_n140 ) , .A1( u0_u4_u7_n153 ) , .B2( u0_u4_u7_n162 ) , .A2( u0_u4_u7_n164 ) );
  INV_X1 u0_u4_u7_U37 (.A( u0_u4_u7_n125 ) , .ZN( u0_u4_u7_n161 ) );
  AOI21_X1 u0_u4_u7_U38 (.ZN( u0_u4_u7_n123 ) , .B1( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n177 ) , .A( u0_u4_u7_n97 ) );
  AOI21_X1 u0_u4_u7_U39 (.B2( u0_u4_u7_n113 ) , .B1( u0_u4_u7_n124 ) , .A( u0_u4_u7_n125 ) , .ZN( u0_u4_u7_n97 ) );
  INV_X1 u0_u4_u7_U4 (.A( u0_u4_u7_n149 ) , .ZN( u0_u4_u7_n175 ) );
  INV_X1 u0_u4_u7_U40 (.A( u0_u4_u7_n152 ) , .ZN( u0_u4_u7_n162 ) );
  AOI22_X1 u0_u4_u7_U41 (.A2( u0_u4_u7_n114 ) , .ZN( u0_u4_u7_n119 ) , .B1( u0_u4_u7_n130 ) , .A1( u0_u4_u7_n156 ) , .B2( u0_u4_u7_n165 ) );
  NAND2_X1 u0_u4_u7_U42 (.A2( u0_u4_u7_n112 ) , .ZN( u0_u4_u7_n114 ) , .A1( u0_u4_u7_n175 ) );
  NOR2_X1 u0_u4_u7_U43 (.ZN( u0_u4_u7_n137 ) , .A1( u0_u4_u7_n150 ) , .A2( u0_u4_u7_n161 ) );
  AND2_X1 u0_u4_u7_U44 (.ZN( u0_u4_u7_n145 ) , .A2( u0_u4_u7_n98 ) , .A1( u0_u4_u7_n99 ) );
  AOI21_X1 u0_u4_u7_U45 (.ZN( u0_u4_u7_n105 ) , .B2( u0_u4_u7_n110 ) , .A( u0_u4_u7_n125 ) , .B1( u0_u4_u7_n147 ) );
  NAND2_X1 u0_u4_u7_U46 (.ZN( u0_u4_u7_n146 ) , .A1( u0_u4_u7_n95 ) , .A2( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U47 (.A2( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n147 ) , .A1( u0_u4_u7_n93 ) );
  NAND2_X1 u0_u4_u7_U48 (.A1( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n127 ) , .A2( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U49 (.A2( u0_u4_u7_n102 ) , .A1( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n133 ) );
  INV_X1 u0_u4_u7_U5 (.A( u0_u4_u7_n154 ) , .ZN( u0_u4_u7_n178 ) );
  OR2_X1 u0_u4_u7_U50 (.ZN( u0_u4_u7_n126 ) , .A2( u0_u4_u7_n152 ) , .A1( u0_u4_u7_n156 ) );
  NAND2_X1 u0_u4_u7_U51 (.ZN( u0_u4_u7_n112 ) , .A2( u0_u4_u7_n96 ) , .A1( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U52 (.A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n128 ) , .A1( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U53 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n113 ) , .A2( u0_u4_u7_n93 ) );
  NAND2_X1 u0_u4_u7_U54 (.ZN( u0_u4_u7_n110 ) , .A1( u0_u4_u7_n95 ) , .A2( u0_u4_u7_n96 ) );
  INV_X1 u0_u4_u7_U55 (.A( u0_u4_u7_n150 ) , .ZN( u0_u4_u7_n164 ) );
  AND2_X1 u0_u4_u7_U56 (.ZN( u0_u4_u7_n134 ) , .A1( u0_u4_u7_n93 ) , .A2( u0_u4_u7_n98 ) );
  NAND2_X1 u0_u4_u7_U57 (.A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n124 ) , .A1( u0_u4_u7_n96 ) );
  NAND2_X1 u0_u4_u7_U58 (.A1( u0_u4_u7_n100 ) , .A2( u0_u4_u7_n102 ) , .ZN( u0_u4_u7_n129 ) );
  NAND2_X1 u0_u4_u7_U59 (.A2( u0_u4_u7_n103 ) , .ZN( u0_u4_u7_n131 ) , .A1( u0_u4_u7_n95 ) );
  AOI211_X1 u0_u4_u7_U6 (.ZN( u0_u4_u7_n116 ) , .A( u0_u4_u7_n155 ) , .C1( u0_u4_u7_n161 ) , .C2( u0_u4_u7_n171 ) , .B( u0_u4_u7_n94 ) );
  NAND2_X1 u0_u4_u7_U60 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n138 ) , .A2( u0_u4_u7_n99 ) );
  NAND2_X1 u0_u4_u7_U61 (.ZN( u0_u4_u7_n132 ) , .A1( u0_u4_u7_n93 ) , .A2( u0_u4_u7_n96 ) );
  NAND2_X1 u0_u4_u7_U62 (.A1( u0_u4_u7_n100 ) , .ZN( u0_u4_u7_n148 ) , .A2( u0_u4_u7_n95 ) );
  AOI211_X1 u0_u4_u7_U63 (.B( u0_u4_u7_n154 ) , .A( u0_u4_u7_n155 ) , .C1( u0_u4_u7_n156 ) , .ZN( u0_u4_u7_n157 ) , .C2( u0_u4_u7_n172 ) );
  INV_X1 u0_u4_u7_U64 (.A( u0_u4_u7_n153 ) , .ZN( u0_u4_u7_n172 ) );
  NOR2_X1 u0_u4_u7_U65 (.A2( u0_u4_X_47 ) , .ZN( u0_u4_u7_n150 ) , .A1( u0_u4_u7_n163 ) );
  NOR2_X1 u0_u4_u7_U66 (.A2( u0_u4_X_43 ) , .A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n103 ) );
  NOR2_X1 u0_u4_u7_U67 (.A2( u0_u4_X_48 ) , .A1( u0_u4_u7_n166 ) , .ZN( u0_u4_u7_n95 ) );
  NOR2_X1 u0_u4_u7_U68 (.A2( u0_u4_X_45 ) , .A1( u0_u4_X_48 ) , .ZN( u0_u4_u7_n99 ) );
  NOR2_X1 u0_u4_u7_U69 (.A2( u0_u4_X_44 ) , .A1( u0_u4_u7_n167 ) , .ZN( u0_u4_u7_n98 ) );
  OAI222_X1 u0_u4_u7_U7 (.C2( u0_u4_u7_n101 ) , .B2( u0_u4_u7_n111 ) , .A1( u0_u4_u7_n113 ) , .C1( u0_u4_u7_n146 ) , .A2( u0_u4_u7_n162 ) , .B1( u0_u4_u7_n164 ) , .ZN( u0_u4_u7_n94 ) );
  NOR2_X1 u0_u4_u7_U70 (.A2( u0_u4_X_46 ) , .A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n152 ) );
  NAND2_X1 u0_u4_u7_U71 (.A2( u0_u4_X_46 ) , .A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n125 ) );
  AND2_X1 u0_u4_u7_U72 (.A1( u0_u4_X_47 ) , .ZN( u0_u4_u7_n156 ) , .A2( u0_u4_u7_n163 ) );
  AND2_X1 u0_u4_u7_U73 (.A2( u0_u4_X_45 ) , .A1( u0_u4_X_48 ) , .ZN( u0_u4_u7_n102 ) );
  AND2_X1 u0_u4_u7_U74 (.A2( u0_u4_X_43 ) , .A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n96 ) );
  AND2_X1 u0_u4_u7_U75 (.A1( u0_u4_X_44 ) , .ZN( u0_u4_u7_n100 ) , .A2( u0_u4_u7_n167 ) );
  AND2_X1 u0_u4_u7_U76 (.A1( u0_u4_X_48 ) , .A2( u0_u4_u7_n166 ) , .ZN( u0_u4_u7_n93 ) );
  INV_X1 u0_u4_u7_U77 (.A( u0_u4_X_46 ) , .ZN( u0_u4_u7_n163 ) );
  INV_X1 u0_u4_u7_U78 (.A( u0_u4_X_43 ) , .ZN( u0_u4_u7_n167 ) );
  INV_X1 u0_u4_u7_U79 (.A( u0_u4_X_45 ) , .ZN( u0_u4_u7_n166 ) );
  OAI221_X1 u0_u4_u7_U8 (.C1( u0_u4_u7_n101 ) , .C2( u0_u4_u7_n147 ) , .ZN( u0_u4_u7_n155 ) , .B2( u0_u4_u7_n162 ) , .A( u0_u4_u7_n91 ) , .B1( u0_u4_u7_n92 ) );
  NAND4_X1 u0_u4_u7_U80 (.ZN( u0_out4_5 ) , .A4( u0_u4_u7_n108 ) , .A3( u0_u4_u7_n109 ) , .A1( u0_u4_u7_n116 ) , .A2( u0_u4_u7_n123 ) );
  AOI22_X1 u0_u4_u7_U81 (.ZN( u0_u4_u7_n109 ) , .A2( u0_u4_u7_n126 ) , .B2( u0_u4_u7_n145 ) , .B1( u0_u4_u7_n156 ) , .A1( u0_u4_u7_n171 ) );
  NOR4_X1 u0_u4_u7_U82 (.A4( u0_u4_u7_n104 ) , .A3( u0_u4_u7_n105 ) , .A2( u0_u4_u7_n106 ) , .A1( u0_u4_u7_n107 ) , .ZN( u0_u4_u7_n108 ) );
  NAND4_X1 u0_u4_u7_U83 (.ZN( u0_out4_27 ) , .A4( u0_u4_u7_n118 ) , .A3( u0_u4_u7_n119 ) , .A2( u0_u4_u7_n120 ) , .A1( u0_u4_u7_n121 ) );
  OAI21_X1 u0_u4_u7_U84 (.ZN( u0_u4_u7_n121 ) , .B2( u0_u4_u7_n145 ) , .A( u0_u4_u7_n150 ) , .B1( u0_u4_u7_n174 ) );
  OAI21_X1 u0_u4_u7_U85 (.ZN( u0_u4_u7_n120 ) , .A( u0_u4_u7_n161 ) , .B2( u0_u4_u7_n170 ) , .B1( u0_u4_u7_n179 ) );
  NAND4_X1 u0_u4_u7_U86 (.ZN( u0_out4_21 ) , .A4( u0_u4_u7_n157 ) , .A3( u0_u4_u7_n158 ) , .A2( u0_u4_u7_n159 ) , .A1( u0_u4_u7_n160 ) );
  OAI21_X1 u0_u4_u7_U87 (.B1( u0_u4_u7_n145 ) , .ZN( u0_u4_u7_n160 ) , .A( u0_u4_u7_n161 ) , .B2( u0_u4_u7_n177 ) );
  AOI22_X1 u0_u4_u7_U88 (.B2( u0_u4_u7_n149 ) , .B1( u0_u4_u7_n150 ) , .A2( u0_u4_u7_n151 ) , .A1( u0_u4_u7_n152 ) , .ZN( u0_u4_u7_n158 ) );
  NAND4_X1 u0_u4_u7_U89 (.ZN( u0_out4_15 ) , .A4( u0_u4_u7_n142 ) , .A3( u0_u4_u7_n143 ) , .A2( u0_u4_u7_n144 ) , .A1( u0_u4_u7_n178 ) );
  AND3_X1 u0_u4_u7_U9 (.A3( u0_u4_u7_n110 ) , .A2( u0_u4_u7_n127 ) , .A1( u0_u4_u7_n132 ) , .ZN( u0_u4_u7_n92 ) );
  OR2_X1 u0_u4_u7_U90 (.A2( u0_u4_u7_n125 ) , .A1( u0_u4_u7_n129 ) , .ZN( u0_u4_u7_n144 ) );
  AOI22_X1 u0_u4_u7_U91 (.A2( u0_u4_u7_n126 ) , .ZN( u0_u4_u7_n143 ) , .B2( u0_u4_u7_n165 ) , .B1( u0_u4_u7_n173 ) , .A1( u0_u4_u7_n174 ) );
  OAI211_X1 u0_u4_u7_U92 (.B( u0_u4_u7_n122 ) , .A( u0_u4_u7_n123 ) , .C2( u0_u4_u7_n124 ) , .ZN( u0_u4_u7_n154 ) , .C1( u0_u4_u7_n162 ) );
  AOI222_X1 u0_u4_u7_U93 (.ZN( u0_u4_u7_n122 ) , .C2( u0_u4_u7_n126 ) , .C1( u0_u4_u7_n145 ) , .B1( u0_u4_u7_n161 ) , .A2( u0_u4_u7_n165 ) , .B2( u0_u4_u7_n170 ) , .A1( u0_u4_u7_n176 ) );
  INV_X1 u0_u4_u7_U94 (.A( u0_u4_u7_n111 ) , .ZN( u0_u4_u7_n170 ) );
  NAND3_X1 u0_u4_u7_U95 (.A3( u0_u4_u7_n146 ) , .A2( u0_u4_u7_n147 ) , .A1( u0_u4_u7_n148 ) , .ZN( u0_u4_u7_n151 ) );
  NAND3_X1 u0_u4_u7_U96 (.A3( u0_u4_u7_n131 ) , .A2( u0_u4_u7_n132 ) , .A1( u0_u4_u7_n133 ) , .ZN( u0_u4_u7_n135 ) );
  OAI21_X1 u0_uk_U1014 (.ZN( u0_K1_37 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n714 ) , .A( u0_uk_n876 ) );
  NAND2_X1 u0_uk_U1015 (.A1( u0_key_r_50 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n876 ) );
  OAI21_X1 u0_uk_U1020 (.ZN( u0_K14_44 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n81 ) , .A( u0_uk_n930 ) );
  NAND2_X1 u0_uk_U1021 (.A1( u0_uk_K_r12_15 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n930 ) );
  OAI22_X1 u0_uk_U103 (.ZN( u0_K5_5 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n466 ) , .A2( u0_uk_n490 ) );
  OAI21_X1 u0_uk_U1042 (.ZN( u0_K14_40 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n65 ) , .A( u0_uk_n931 ) );
  NAND2_X1 u0_uk_U1043 (.A1( u0_uk_K_r12_21 ) , .A2( u0_uk_n110 ) , .ZN( u0_uk_n931 ) );
  INV_X1 u0_uk_U1062 (.A( u0_key_r_9 ) , .ZN( u0_uk_n709 ) );
  INV_X1 u0_uk_U1063 (.A( u0_key_r_7 ) , .ZN( u0_uk_n711 ) );
  INV_X1 u0_uk_U1067 (.A( u0_key_r_23 ) , .ZN( u0_uk_n700 ) );
  INV_X1 u0_uk_U1069 (.A( u0_key_r_30 ) , .ZN( u0_uk_n693 ) );
  INV_X1 u0_uk_U1074 (.A( u0_key_r_37 ) , .ZN( u0_uk_n687 ) );
  INV_X1 u0_uk_U1075 (.A( u0_key_r_52 ) , .ZN( u0_uk_n675 ) );
  INV_X1 u0_uk_U1076 (.A( u0_key_r_0 ) , .ZN( u0_uk_n716 ) );
  INV_X1 u0_uk_U1077 (.A( u0_key_r_16 ) , .ZN( u0_uk_n706 ) );
  INV_X1 u0_uk_U1079 (.A( u0_key_r_1 ) , .ZN( u0_uk_n715 ) );
  INV_X1 u0_uk_U1080 (.A( u0_key_r_2 ) , .ZN( u0_uk_n714 ) );
  OAI22_X1 u0_uk_U109 (.ZN( u0_K14_41 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n77 ) , .A2( u0_uk_n82 ) , .B1( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U1097 (.ZN( u0_K5_39 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n482 ) , .A( u0_uk_n808 ) );
  NAND2_X1 u0_uk_U1098 (.A1( u0_uk_K_r3_16 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n808 ) );
  INV_X1 u0_uk_U1107 (.ZN( u0_K1_41 ) , .A( u0_uk_n874 ) );
  AOI22_X1 u0_uk_U1108 (.B2( u0_key_r_35 ) , .A2( u0_key_r_42 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n874 ) );
  INV_X1 u0_uk_U1125 (.ZN( u0_K1_32 ) , .A( u0_uk_n879 ) );
  AOI22_X1 u0_uk_U1126 (.B2( u0_key_r_22 ) , .A2( u0_key_r_29 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n879 ) );
  INV_X1 u0_uk_U1147 (.ZN( u0_K5_35 ) , .A( u0_uk_n810 ) );
  AOI22_X1 u0_uk_U1149 (.B2( u0_uk_K_r3_15 ) , .A2( u0_uk_K_r3_38 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n230 ) , .ZN( u0_uk_n806 ) );
  INV_X1 u0_uk_U1150 (.ZN( u0_K5_43 ) , .A( u0_uk_n806 ) );
  OAI21_X1 u0_uk_U1151 (.ZN( u0_K5_6 ) , .B1( u0_uk_n109 ) , .B2( u0_uk_n471 ) , .A( u0_uk_n803 ) );
  NAND2_X1 u0_uk_U1152 (.A1( u0_uk_K_r3_10 ) , .ZN( u0_uk_n803 ) , .A2( u0_uk_n93 ) );
  INV_X1 u0_uk_U213 (.A( u0_key_r_14 ) , .ZN( u0_uk_n707 ) );
  OAI21_X1 u0_uk_U231 (.ZN( u0_K1_39 ) , .B1( u0_uk_n118 ) , .B2( u0_uk_n701 ) , .A( u0_uk_n875 ) );
  INV_X1 u0_uk_U233 (.A( u0_key_r_22 ) , .ZN( u0_uk_n701 ) );
  OAI22_X1 u0_uk_U237 (.ZN( u0_K14_39 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n56 ) );
  INV_X1 u0_uk_U250 (.ZN( u0_K1_48 ) , .A( u0_uk_n870 ) );
  AOI22_X1 u0_uk_U251 (.B2( u0_key_r_21 ) , .A2( u0_key_r_28 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n870 ) );
  INV_X1 u0_uk_U252 (.ZN( u0_K1_44 ) , .A( u0_uk_n872 ) );
  AOI22_X1 u0_uk_U253 (.B2( u0_key_r_36 ) , .A2( u0_key_r_43 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n872 ) );
  OAI22_X1 u0_uk_U254 (.ZN( u0_K14_48 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n90 ) );
  INV_X1 u0_uk_U297 (.ZN( u0_K1_26 ) , .A( u0_uk_n883 ) );
  AOI22_X1 u0_uk_U298 (.B2( u0_key_r_31 ) , .A2( u0_key_r_51 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n883 ) );
  OAI22_X1 u0_uk_U325 (.ZN( u0_K5_46 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n457 ) , .B2( u0_uk_n494 ) );
  OAI22_X1 u0_uk_U357 (.ZN( u0_K1_40 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n675 ) , .B2( u0_uk_n716 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U371 (.ZN( u0_K1_28 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n710 ) , .B2( u0_uk_n715 ) );
  INV_X1 u0_uk_U372 (.A( u0_key_r_8 ) , .ZN( u0_uk_n710 ) );
  OAI21_X1 u0_uk_U379 (.ZN( u0_K5_33 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n457 ) , .A( u0_uk_n811 ) );
  NAND2_X1 u0_uk_U380 (.A1( u0_uk_K_r3_14 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n811 ) );
  INV_X1 u0_uk_U426 (.ZN( u0_K1_33 ) , .A( u0_uk_n878 ) );
  OAI22_X1 u0_uk_U451 (.ZN( u0_K14_37 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n67 ) , .B2( u0_uk_n73 ) );
  OAI22_X1 u0_uk_U467 (.ZN( u0_K5_37 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n455 ) , .B2( u0_uk_n493 ) );
  OAI22_X1 u0_uk_U469 (.ZN( u0_K1_29 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n700 ) , .B2( u0_uk_n706 ) );
  OAI22_X1 u0_uk_U530 (.ZN( u0_K5_2 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n486 ) , .A2( u0_uk_n491 ) );
  OAI22_X1 u0_uk_U531 (.ZN( u0_K1_36 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n693 ) , .B2( u0_uk_n700 ) );
  OAI22_X1 u0_uk_U549 (.ZN( u0_K1_38 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n687 ) , .B2( u0_uk_n693 ) );
  INV_X1 u0_uk_U550 (.ZN( u0_K5_36 ) , .A( u0_uk_n809 ) );
  AOI22_X1 u0_uk_U551 (.B2( u0_uk_K_r3_29 ) , .A2( u0_uk_K_r3_52 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n809 ) );
  INV_X1 u0_uk_U620 (.ZN( u0_K1_35 ) , .A( u0_uk_n877 ) );
  AOI22_X1 u0_uk_U621 (.B2( u0_key_r_28 ) , .A2( u0_key_r_35 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n877 ) );
  OAI22_X1 u0_uk_U650 (.ZN( u0_K14_43 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n56 ) , .B2( u0_uk_n59 ) , .A1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U662 (.ZN( u0_K14_45 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n58 ) , .A( u0_uk_n929 ) );
  NAND2_X1 u0_uk_U663 (.A1( u0_uk_K_r12_16 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n929 ) );
  OAI21_X1 u0_uk_U673 (.ZN( u0_K5_45 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n488 ) , .A( u0_uk_n805 ) );
  INV_X1 u0_uk_U710 (.ZN( u0_K1_25 ) , .A( u0_uk_n884 ) );
  AOI22_X1 u0_uk_U711 (.B2( u0_key_r_29 ) , .A2( u0_key_r_36 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n884 ) );
  OAI21_X1 u0_uk_U731 (.ZN( u0_K5_42 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n476 ) , .A( u0_uk_n807 ) );
  NAND2_X1 u0_uk_U732 (.A1( u0_uk_K_r3_9 ) , .ZN( u0_uk_n807 ) , .A2( u0_uk_n92 ) );
  INV_X1 u0_uk_U742 (.ZN( u0_K1_42 ) , .A( u0_uk_n873 ) );
  AOI22_X1 u0_uk_U743 (.B2( u0_key_r_31 ) , .A2( u0_key_r_38 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n873 ) );
  INV_X1 u0_uk_U794 (.ZN( u0_K1_27 ) , .A( u0_uk_n882 ) );
  AOI22_X1 u0_uk_U795 (.B2( u0_key_r_14 ) , .A2( u0_key_r_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n882 ) );
  OAI22_X1 u0_uk_U843 (.ZN( u0_K1_43 ) , .B1( u0_uk_n109 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n706 ) , .A2( u0_uk_n709 ) );
  OAI22_X1 u0_uk_U947 (.ZN( u0_K14_47 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n58 ) , .B2( u0_uk_n68 ) );
  OAI22_X1 u0_uk_U966 (.ZN( u0_K14_38 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n65 ) , .A2( u0_uk_n81 ) );
  OAI22_X1 u0_uk_U972 (.ZN( u0_K5_40 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n458 ) , .B2( u0_uk_n475 ) );
  OAI22_X1 u0_uk_U991 (.ZN( u0_K1_34 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n709 ) , .B2( u0_uk_n714 ) );
  OAI22_X1 u0_uk_U992 (.ZN( u0_K1_47 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n711 ) , .B2( u0_uk_n716 ) );
  XOR2_X1 u2_U103 (.B( u2_L0_13 ) , .Z( u2_N44 ) , .A( u2_out1_13 ) );
  XOR2_X1 u2_U131 (.B( u2_L11_31 ) , .Z( u2_N414 ) , .A( u2_out12_31 ) );
  XOR2_X1 u2_U132 (.B( u2_L11_30 ) , .Z( u2_N413 ) , .A( u2_out12_30 ) );
  XOR2_X1 u2_U133 (.B( u2_L11_29 ) , .Z( u2_N412 ) , .A( u2_out12_29 ) );
  XOR2_X1 u2_U134 (.B( u2_L11_28 ) , .Z( u2_N411 ) , .A( u2_out12_28 ) );
  XOR2_X1 u2_U136 (.B( u2_L0_10 ) , .Z( u2_N41 ) , .A( u2_out1_10 ) );
  XOR2_X1 u2_U137 (.B( u2_L11_26 ) , .Z( u2_N409 ) , .A( u2_out12_26 ) );
  XOR2_X1 u2_U138 (.B( u2_L11_25 ) , .Z( u2_N408 ) , .A( u2_out12_25 ) );
  XOR2_X1 u2_U139 (.B( u2_L11_24 ) , .Z( u2_N407 ) , .A( u2_out12_24 ) );
  XOR2_X1 u2_U140 (.B( u2_L11_23 ) , .Z( u2_N406 ) , .A( u2_out12_23 ) );
  XOR2_X1 u2_U143 (.B( u2_L11_20 ) , .Z( u2_N403 ) , .A( u2_out12_20 ) );
  XOR2_X1 u2_U144 (.B( u2_L11_19 ) , .Z( u2_N402 ) , .A( u2_out12_19 ) );
  XOR2_X1 u2_U145 (.B( u2_L11_18 ) , .Z( u2_N401 ) , .A( u2_out12_18 ) );
  XOR2_X1 u2_U146 (.B( u2_L11_17 ) , .Z( u2_N400 ) , .A( u2_out12_17 ) );
  XOR2_X1 u2_U148 (.Z( u2_N4 ) , .B( u2_desIn_r_38 ) , .A( u2_out0_5 ) );
  XOR2_X1 u2_U149 (.B( u2_L11_16 ) , .Z( u2_N399 ) , .A( u2_out12_16 ) );
  XOR2_X1 u2_U15 (.B( u2_L1_25 ) , .Z( u2_N88 ) , .A( u2_out2_25 ) );
  XOR2_X1 u2_U151 (.B( u2_L11_14 ) , .Z( u2_N397 ) , .A( u2_out12_14 ) );
  XOR2_X1 u2_U152 (.B( u2_L11_13 ) , .Z( u2_N396 ) , .A( u2_out12_13 ) );
  XOR2_X1 u2_U154 (.B( u2_L11_11 ) , .Z( u2_N394 ) , .A( u2_out12_11 ) );
  XOR2_X1 u2_U155 (.B( u2_L11_10 ) , .Z( u2_N393 ) , .A( u2_out12_10 ) );
  XOR2_X1 u2_U156 (.B( u2_L11_9 ) , .Z( u2_N392 ) , .A( u2_out12_9 ) );
  XOR2_X1 u2_U157 (.B( u2_L11_8 ) , .Z( u2_N391 ) , .A( u2_out12_8 ) );
  XOR2_X1 u2_U160 (.B( u2_L11_6 ) , .Z( u2_N389 ) , .A( u2_out12_6 ) );
  XOR2_X1 u2_U162 (.B( u2_L11_4 ) , .Z( u2_N387 ) , .A( u2_out12_4 ) );
  XOR2_X1 u2_U163 (.B( u2_L11_3 ) , .Z( u2_N386 ) , .A( u2_out12_3 ) );
  XOR2_X1 u2_U164 (.B( u2_L11_2 ) , .Z( u2_N385 ) , .A( u2_out12_2 ) );
  XOR2_X1 u2_U165 (.B( u2_L11_1 ) , .Z( u2_N384 ) , .A( u2_out12_1 ) );
  XOR2_X1 u2_U166 (.B( u2_L10_32 ) , .Z( u2_N383 ) , .A( u2_out11_32 ) );
  XOR2_X1 u2_U169 (.B( u2_L10_29 ) , .Z( u2_N380 ) , .A( u2_out11_29 ) );
  XOR2_X1 u2_U172 (.B( u2_L10_27 ) , .Z( u2_N378 ) , .A( u2_out11_27 ) );
  XOR2_X1 u2_U173 (.B( u2_L10_26 ) , .Z( u2_N377 ) , .A( u2_out11_26 ) );
  XOR2_X1 u2_U174 (.B( u2_L10_25 ) , .Z( u2_N376 ) , .A( u2_out11_25 ) );
  XOR2_X1 u2_U177 (.B( u2_L10_22 ) , .Z( u2_N373 ) , .A( u2_out11_22 ) );
  XOR2_X1 u2_U178 (.B( u2_L10_21 ) , .Z( u2_N372 ) , .A( u2_out11_21 ) );
  XOR2_X1 u2_U179 (.B( u2_L10_20 ) , .Z( u2_N371 ) , .A( u2_out11_20 ) );
  XOR2_X1 u2_U180 (.B( u2_L10_19 ) , .Z( u2_N370 ) , .A( u2_out11_19 ) );
  XOR2_X1 u2_U181 (.B( u2_L0_6 ) , .Z( u2_N37 ) , .A( u2_out1_6 ) );
  XOR2_X1 u2_U185 (.B( u2_L10_15 ) , .Z( u2_N366 ) , .A( u2_out11_15 ) );
  XOR2_X1 u2_U186 (.B( u2_L10_14 ) , .Z( u2_N365 ) , .A( u2_out11_14 ) );
  XOR2_X1 u2_U188 (.B( u2_L10_12 ) , .Z( u2_N363 ) , .A( u2_out11_12 ) );
  XOR2_X1 u2_U189 (.B( u2_L10_11 ) , .Z( u2_N362 ) , .A( u2_out11_11 ) );
  XOR2_X1 u2_U190 (.B( u2_L10_10 ) , .Z( u2_N361 ) , .A( u2_out11_10 ) );
  XOR2_X1 u2_U193 (.B( u2_L10_8 ) , .Z( u2_N359 ) , .A( u2_out11_8 ) );
  XOR2_X1 u2_U194 (.B( u2_L10_7 ) , .Z( u2_N358 ) , .A( u2_out11_7 ) );
  XOR2_X1 u2_U196 (.B( u2_L10_5 ) , .Z( u2_N356 ) , .A( u2_out11_5 ) );
  XOR2_X1 u2_U197 (.B( u2_L10_4 ) , .Z( u2_N355 ) , .A( u2_out11_4 ) );
  XOR2_X1 u2_U198 (.B( u2_L10_3 ) , .Z( u2_N354 ) , .A( u2_out11_3 ) );
  XOR2_X1 u2_U200 (.B( u2_L10_1 ) , .Z( u2_N352 ) , .A( u2_out11_1 ) );
  XOR2_X1 u2_U201 (.B( u2_L9_32 ) , .Z( u2_N351 ) , .A( u2_out10_32 ) );
  XOR2_X1 u2_U204 (.B( u2_L9_30 ) , .Z( u2_N349 ) , .A( u2_out10_30 ) );
  XOR2_X1 u2_U205 (.B( u2_L9_29 ) , .Z( u2_N348 ) , .A( u2_out10_29 ) );
  XOR2_X1 u2_U207 (.B( u2_L9_27 ) , .Z( u2_N346 ) , .A( u2_out10_27 ) );
  XOR2_X1 u2_U210 (.B( u2_L9_24 ) , .Z( u2_N343 ) , .A( u2_out10_24 ) );
  XOR2_X1 u2_U212 (.B( u2_L9_22 ) , .Z( u2_N341 ) , .A( u2_out10_22 ) );
  XOR2_X1 u2_U213 (.B( u2_L9_21 ) , .Z( u2_N340 ) , .A( u2_out10_21 ) );
  XOR2_X1 u2_U216 (.B( u2_L9_19 ) , .Z( u2_N338 ) , .A( u2_out10_19 ) );
  XOR2_X1 u2_U219 (.B( u2_L9_16 ) , .Z( u2_N335 ) , .A( u2_out10_16 ) );
  XOR2_X1 u2_U220 (.B( u2_L9_15 ) , .Z( u2_N334 ) , .A( u2_out10_15 ) );
  XOR2_X1 u2_U223 (.B( u2_L9_12 ) , .Z( u2_N331 ) , .A( u2_out10_12 ) );
  XOR2_X1 u2_U224 (.B( u2_L9_11 ) , .Z( u2_N330 ) , .A( u2_out10_11 ) );
  XOR2_X1 u2_U225 (.B( u2_L0_2 ) , .Z( u2_N33 ) , .A( u2_out1_2 ) );
  XOR2_X1 u2_U229 (.B( u2_L9_7 ) , .Z( u2_N326 ) , .A( u2_out10_7 ) );
  XOR2_X1 u2_U230 (.B( u2_L9_6 ) , .Z( u2_N325 ) , .A( u2_out10_6 ) );
  XOR2_X1 u2_U231 (.B( u2_L9_5 ) , .Z( u2_N324 ) , .A( u2_out10_5 ) );
  XOR2_X1 u2_U232 (.B( u2_L9_4 ) , .Z( u2_N323 ) , .A( u2_out10_4 ) );
  XOR2_X1 u2_U236 (.B( u2_L0_1 ) , .Z( u2_N32 ) , .A( u2_out1_1 ) );
  XOR2_X1 u2_U237 (.B( u2_L8_32 ) , .Z( u2_N319 ) , .A( u2_out9_32 ) );
  XOR2_X1 u2_U240 (.B( u2_L8_29 ) , .Z( u2_N316 ) , .A( u2_out9_29 ) );
  XOR2_X1 u2_U243 (.B( u2_L8_26 ) , .Z( u2_N313 ) , .A( u2_out9_26 ) );
  XOR2_X1 u2_U244 (.B( u2_L8_25 ) , .Z( u2_N312 ) , .A( u2_out9_25 ) );
  XOR2_X1 u2_U247 (.Z( u2_N31 ) , .B( u2_desIn_r_56 ) , .A( u2_out0_32 ) );
  XOR2_X1 u2_U248 (.B( u2_L8_22 ) , .Z( u2_N309 ) , .A( u2_out9_22 ) );
  XOR2_X1 u2_U250 (.B( u2_L8_20 ) , .Z( u2_N307 ) , .A( u2_out9_20 ) );
  XOR2_X1 u2_U251 (.B( u2_L8_19 ) , .Z( u2_N306 ) , .A( u2_out9_19 ) );
  XOR2_X1 u2_U256 (.B( u2_L8_14 ) , .Z( u2_N301 ) , .A( u2_out9_14 ) );
  XOR2_X1 u2_U259 (.Z( u2_N3 ) , .B( u2_desIn_r_30 ) , .A( u2_out0_4 ) );
  XOR2_X1 u2_U260 (.B( u2_L8_12 ) , .Z( u2_N299 ) , .A( u2_out9_12 ) );
  XOR2_X1 u2_U261 (.B( u2_L8_11 ) , .Z( u2_N298 ) , .A( u2_out9_11 ) );
  XOR2_X1 u2_U262 (.B( u2_L8_10 ) , .Z( u2_N297 ) , .A( u2_out9_10 ) );
  XOR2_X1 u2_U264 (.B( u2_L8_8 ) , .Z( u2_N295 ) , .A( u2_out9_8 ) );
  XOR2_X1 u2_U265 (.B( u2_L8_7 ) , .Z( u2_N294 ) , .A( u2_out9_7 ) );
  XOR2_X1 u2_U268 (.B( u2_L8_4 ) , .Z( u2_N291 ) , .A( u2_out9_4 ) );
  XOR2_X1 u2_U269 (.B( u2_L8_3 ) , .Z( u2_N290 ) , .A( u2_out9_3 ) );
  XOR2_X1 u2_U27 (.B( u2_L1_14 ) , .Z( u2_N77 ) , .A( u2_out2_14 ) );
  XOR2_X1 u2_U272 (.B( u2_L8_1 ) , .Z( u2_N288 ) , .A( u2_out9_1 ) );
  XOR2_X1 u2_U273 (.B( u2_L7_32 ) , .Z( u2_N287 ) , .A( u2_out8_32 ) );
  XOR2_X1 u2_U274 (.B( u2_L7_31 ) , .Z( u2_N286 ) , .A( u2_out8_31 ) );
  XOR2_X1 u2_U275 (.B( u2_L7_30 ) , .Z( u2_N285 ) , .A( u2_out8_30 ) );
  XOR2_X1 u2_U277 (.B( u2_L7_28 ) , .Z( u2_N283 ) , .A( u2_out8_28 ) );
  XOR2_X1 u2_U278 (.B( u2_L7_27 ) , .Z( u2_N282 ) , .A( u2_out8_27 ) );
  XOR2_X1 u2_U279 (.B( u2_L7_26 ) , .Z( u2_N281 ) , .A( u2_out8_26 ) );
  XOR2_X1 u2_U280 (.B( u2_L7_25 ) , .Z( u2_N280 ) , .A( u2_out8_25 ) );
  XOR2_X1 u2_U281 (.Z( u2_N28 ) , .B( u2_desIn_r_32 ) , .A( u2_out0_29 ) );
  XOR2_X1 u2_U282 (.B( u2_L7_24 ) , .Z( u2_N279 ) , .A( u2_out8_24 ) );
  XOR2_X1 u2_U283 (.B( u2_L7_23 ) , .Z( u2_N278 ) , .A( u2_out8_23 ) );
  XOR2_X1 u2_U284 (.B( u2_L7_22 ) , .Z( u2_N277 ) , .A( u2_out8_22 ) );
  XOR2_X1 u2_U285 (.B( u2_L7_21 ) , .Z( u2_N276 ) , .A( u2_out8_21 ) );
  XOR2_X1 u2_U286 (.B( u2_L7_20 ) , .Z( u2_N275 ) , .A( u2_out8_20 ) );
  XOR2_X1 u2_U288 (.B( u2_L7_18 ) , .Z( u2_N273 ) , .A( u2_out8_18 ) );
  XOR2_X1 u2_U289 (.B( u2_L7_17 ) , .Z( u2_N272 ) , .A( u2_out8_17 ) );
  XOR2_X1 u2_U290 (.B( u2_L7_16 ) , .Z( u2_N271 ) , .A( u2_out8_16 ) );
  XOR2_X1 u2_U291 (.B( u2_L7_15 ) , .Z( u2_N270 ) , .A( u2_out8_15 ) );
  XOR2_X1 u2_U293 (.B( u2_L7_14 ) , .Z( u2_N269 ) , .A( u2_out8_14 ) );
  XOR2_X1 u2_U294 (.B( u2_L7_13 ) , .Z( u2_N268 ) , .A( u2_out8_13 ) );
  XOR2_X1 u2_U295 (.B( u2_L7_12 ) , .Z( u2_N267 ) , .A( u2_out8_12 ) );
  XOR2_X1 u2_U297 (.B( u2_L7_10 ) , .Z( u2_N265 ) , .A( u2_out8_10 ) );
  XOR2_X1 u2_U298 (.B( u2_L7_9 ) , .Z( u2_N264 ) , .A( u2_out8_9 ) );
  XOR2_X1 u2_U299 (.B( u2_L7_8 ) , .Z( u2_N263 ) , .A( u2_out8_8 ) );
  XOR2_X1 u2_U300 (.B( u2_L7_7 ) , .Z( u2_N262 ) , .A( u2_out8_7 ) );
  XOR2_X1 u2_U301 (.B( u2_L7_6 ) , .Z( u2_N261 ) , .A( u2_out8_6 ) );
  XOR2_X1 u2_U302 (.B( u2_L7_5 ) , .Z( u2_N260 ) , .A( u2_out8_5 ) );
  XOR2_X1 u2_U303 (.Z( u2_N26 ) , .B( u2_desIn_r_16 ) , .A( u2_out0_27 ) );
  XOR2_X1 u2_U305 (.B( u2_L7_3 ) , .Z( u2_N258 ) , .A( u2_out8_3 ) );
  XOR2_X1 u2_U306 (.B( u2_L7_2 ) , .Z( u2_N257 ) , .A( u2_out8_2 ) );
  XOR2_X1 u2_U307 (.B( u2_L7_1 ) , .Z( u2_N256 ) , .A( u2_out8_1 ) );
  XOR2_X1 u2_U311 (.B( u2_L6_29 ) , .Z( u2_N252 ) , .A( u2_out7_29 ) );
  XOR2_X1 u2_U316 (.B( u2_L6_25 ) , .Z( u2_N248 ) , .A( u2_out7_25 ) );
  XOR2_X1 u2_U322 (.B( u2_L6_19 ) , .Z( u2_N242 ) , .A( u2_out7_19 ) );
  XOR2_X1 u2_U325 (.Z( u2_N24 ) , .B( u2_desIn_r_0 ) , .A( u2_out0_25 ) );
  XOR2_X1 u2_U328 (.B( u2_L6_14 ) , .Z( u2_N237 ) , .A( u2_out7_14 ) );
  XOR2_X1 u2_U33 (.B( u2_L1_8 ) , .Z( u2_N71 ) , .A( u2_out2_8 ) );
  XOR2_X1 u2_U331 (.B( u2_L6_11 ) , .Z( u2_N234 ) , .A( u2_out7_11 ) );
  XOR2_X1 u2_U334 (.B( u2_L6_8 ) , .Z( u2_N231 ) , .A( u2_out7_8 ) );
  XOR2_X1 u2_U339 (.B( u2_L6_4 ) , .Z( u2_N227 ) , .A( u2_out7_4 ) );
  XOR2_X1 u2_U340 (.B( u2_L6_3 ) , .Z( u2_N226 ) , .A( u2_out7_3 ) );
  XOR2_X1 u2_U346 (.B( u2_L5_29 ) , .Z( u2_N220 ) , .A( u2_out6_29 ) );
  XOR2_X1 u2_U35 (.Z( u2_N7 ) , .B( u2_desIn_r_62 ) , .A( u2_out0_8 ) );
  XOR2_X1 u2_U357 (.B( u2_L5_19 ) , .Z( u2_N210 ) , .A( u2_out6_19 ) );
  XOR2_X1 u2_U358 (.Z( u2_N21 ) , .B( u2_desIn_r_42 ) , .A( u2_out0_22 ) );
  XOR2_X1 u2_U366 (.B( u2_L5_11 ) , .Z( u2_N202 ) , .A( u2_out6_11 ) );
  XOR2_X1 u2_U369 (.Z( u2_N20 ) , .B( u2_desIn_r_34 ) , .A( u2_out0_21 ) );
  XOR2_X1 u2_U370 (.Z( u2_N2 ) , .B( u2_desIn_r_22 ) , .A( u2_out0_3 ) );
  XOR2_X1 u2_U375 (.B( u2_L5_4 ) , .Z( u2_N195 ) , .A( u2_out6_4 ) );
  XOR2_X1 u2_U379 (.B( u2_L4_32 ) , .Z( u2_N191 ) , .A( u2_out5_32 ) );
  XOR2_X1 u2_U380 (.B( u2_L4_31 ) , .Z( u2_N190 ) , .A( u2_out5_31 ) );
  XOR2_X1 u2_U383 (.B( u2_L4_29 ) , .Z( u2_N188 ) , .A( u2_out5_29 ) );
  XOR2_X1 u2_U384 (.B( u2_L4_28 ) , .Z( u2_N187 ) , .A( u2_out5_28 ) );
  XOR2_X1 u2_U385 (.B( u2_L4_27 ) , .Z( u2_N186 ) , .A( u2_out5_27 ) );
  XOR2_X1 u2_U389 (.B( u2_L4_23 ) , .Z( u2_N182 ) , .A( u2_out5_23 ) );
  XOR2_X1 u2_U39 (.B( u2_L1_3 ) , .Z( u2_N66 ) , .A( u2_out2_3 ) );
  XOR2_X1 u2_U390 (.B( u2_L4_22 ) , .Z( u2_N181 ) , .A( u2_out5_22 ) );
  XOR2_X1 u2_U391 (.B( u2_L4_21 ) , .Z( u2_N180 ) , .A( u2_out5_21 ) );
  XOR2_X1 u2_U392 (.Z( u2_N18 ) , .B( u2_desIn_r_18 ) , .A( u2_out0_19 ) );
  XOR2_X1 u2_U394 (.B( u2_L4_19 ) , .Z( u2_N178 ) , .A( u2_out5_19 ) );
  XOR2_X1 u2_U395 (.B( u2_L4_18 ) , .Z( u2_N177 ) , .A( u2_out5_18 ) );
  XOR2_X1 u2_U396 (.B( u2_L4_17 ) , .Z( u2_N176 ) , .A( u2_out5_17 ) );
  XOR2_X1 u2_U398 (.B( u2_L4_15 ) , .Z( u2_N174 ) , .A( u2_out5_15 ) );
  XOR2_X1 u2_U400 (.B( u2_L4_13 ) , .Z( u2_N172 ) , .A( u2_out5_13 ) );
  XOR2_X1 u2_U401 (.B( u2_L4_12 ) , .Z( u2_N171 ) , .A( u2_out5_12 ) );
  XOR2_X1 u2_U402 (.B( u2_L4_11 ) , .Z( u2_N170 ) , .A( u2_out5_11 ) );
  XOR2_X1 u2_U405 (.B( u2_L4_9 ) , .Z( u2_N168 ) , .A( u2_out5_9 ) );
  XOR2_X1 u2_U407 (.B( u2_L4_7 ) , .Z( u2_N166 ) , .A( u2_out5_7 ) );
  XOR2_X1 u2_U409 (.B( u2_L4_5 ) , .Z( u2_N164 ) , .A( u2_out5_5 ) );
  XOR2_X1 u2_U410 (.B( u2_L4_4 ) , .Z( u2_N163 ) , .A( u2_out5_4 ) );
  XOR2_X1 u2_U412 (.B( u2_L4_2 ) , .Z( u2_N161 ) , .A( u2_out5_2 ) );
  XOR2_X1 u2_U415 (.B( u2_L3_32 ) , .Z( u2_N159 ) , .A( u2_out4_32 ) );
  XOR2_X1 u2_U418 (.B( u2_L3_29 ) , .Z( u2_N156 ) , .A( u2_out4_29 ) );
  XOR2_X1 u2_U422 (.B( u2_L3_25 ) , .Z( u2_N152 ) , .A( u2_out4_25 ) );
  XOR2_X1 u2_U426 (.B( u2_L3_22 ) , .Z( u2_N149 ) , .A( u2_out4_22 ) );
  XOR2_X1 u2_U429 (.B( u2_L3_19 ) , .Z( u2_N146 ) , .A( u2_out4_19 ) );
  XOR2_X1 u2_U434 (.B( u2_L3_14 ) , .Z( u2_N141 ) , .A( u2_out4_14 ) );
  XOR2_X1 u2_U436 (.Z( u2_N14 ) , .B( u2_desIn_r_52 ) , .A( u2_out0_15 ) );
  XOR2_X1 u2_U437 (.B( u2_L3_12 ) , .Z( u2_N139 ) , .A( u2_out4_12 ) );
  XOR2_X1 u2_U438 (.B( u2_L3_11 ) , .Z( u2_N138 ) , .A( u2_out4_11 ) );
  XOR2_X1 u2_U44 (.B( u2_L0_30 ) , .Z( u2_N61 ) , .A( u2_out1_30 ) );
  XOR2_X1 u2_U441 (.B( u2_L3_8 ) , .Z( u2_N135 ) , .A( u2_out4_8 ) );
  XOR2_X1 u2_U442 (.B( u2_L3_7 ) , .Z( u2_N134 ) , .A( u2_out4_7 ) );
  XOR2_X1 u2_U445 (.B( u2_L3_4 ) , .Z( u2_N131 ) , .A( u2_out4_4 ) );
  XOR2_X1 u2_U446 (.B( u2_L3_3 ) , .Z( u2_N130 ) , .A( u2_out4_3 ) );
  XOR2_X1 u2_U447 (.Z( u2_N13 ) , .B( u2_desIn_r_44 ) , .A( u2_out0_14 ) );
  XOR2_X1 u2_U450 (.B( u2_L2_32 ) , .Z( u2_N127 ) , .A( u2_out3_32 ) );
  XOR2_X1 u2_U451 (.B( u2_L2_31 ) , .Z( u2_N126 ) , .A( u2_out3_31 ) );
  XOR2_X1 u2_U454 (.B( u2_L2_28 ) , .Z( u2_N123 ) , .A( u2_out3_28 ) );
  XOR2_X1 u2_U455 (.B( u2_L2_27 ) , .Z( u2_N122 ) , .A( u2_out3_27 ) );
  XOR2_X1 u2_U46 (.Z( u2_N6 ) , .B( u2_desIn_r_54 ) , .A( u2_out0_7 ) );
  XOR2_X1 u2_U460 (.B( u2_L2_23 ) , .Z( u2_N118 ) , .A( u2_out3_23 ) );
  XOR2_X1 u2_U461 (.B( u2_L2_22 ) , .Z( u2_N117 ) , .A( u2_out3_22 ) );
  XOR2_X1 u2_U462 (.B( u2_L2_21 ) , .Z( u2_N116 ) , .A( u2_out3_21 ) );
  XOR2_X1 u2_U465 (.B( u2_L2_18 ) , .Z( u2_N113 ) , .A( u2_out3_18 ) );
  XOR2_X1 u2_U466 (.B( u2_L2_17 ) , .Z( u2_N112 ) , .A( u2_out3_17 ) );
  XOR2_X1 u2_U468 (.B( u2_L2_15 ) , .Z( u2_N110 ) , .A( u2_out3_15 ) );
  XOR2_X1 u2_U469 (.Z( u2_N11 ) , .B( u2_desIn_r_28 ) , .A( u2_out0_12 ) );
  XOR2_X1 u2_U47 (.B( u2_L0_28 ) , .Z( u2_N59 ) , .A( u2_out1_28 ) );
  XOR2_X1 u2_U471 (.B( u2_L2_13 ) , .Z( u2_N108 ) , .A( u2_out3_13 ) );
  XOR2_X1 u2_U472 (.B( u2_L2_12 ) , .Z( u2_N107 ) , .A( u2_out3_12 ) );
  XOR2_X1 u2_U475 (.B( u2_L2_9 ) , .Z( u2_N104 ) , .A( u2_out3_9 ) );
  XOR2_X1 u2_U477 (.B( u2_L2_7 ) , .Z( u2_N102 ) , .A( u2_out3_7 ) );
  XOR2_X1 u2_U479 (.B( u2_L2_5 ) , .Z( u2_N100 ) , .A( u2_out3_5 ) );
  XOR2_X1 u2_U480 (.Z( u2_N10 ) , .B( u2_desIn_r_20 ) , .A( u2_out0_11 ) );
  XOR2_X1 u2_U486 (.Z( u2_FP_6 ) , .B( u2_L14_6 ) , .A( u2_out15_6 ) );
  XOR2_X1 u2_U49 (.B( u2_L0_26 ) , .Z( u2_N57 ) , .A( u2_out1_26 ) );
  XOR2_X1 u2_U492 (.Z( u2_FP_30 ) , .B( u2_L14_30 ) , .A( u2_out15_30 ) );
  XOR2_X1 u2_U493 (.Z( u2_FP_2 ) , .B( u2_L14_2 ) , .A( u2_out15_2 ) );
  XOR2_X1 u2_U495 (.Z( u2_FP_28 ) , .B( u2_L14_28 ) , .A( u2_out15_28 ) );
  XOR2_X1 u2_U497 (.Z( u2_FP_26 ) , .B( u2_L14_26 ) , .A( u2_out15_26 ) );
  XOR2_X1 u2_U499 (.Z( u2_FP_24 ) , .B( u2_L14_24 ) , .A( u2_out15_24 ) );
  XOR2_X1 u2_U5 (.B( u2_L2_2 ) , .Z( u2_N97 ) , .A( u2_out3_2 ) );
  XOR2_X1 u2_U503 (.Z( u2_FP_20 ) , .B( u2_L14_20 ) , .A( u2_out15_20 ) );
  XOR2_X1 u2_U504 (.Z( u2_FP_1 ) , .B( u2_L14_1 ) , .A( u2_out15_1 ) );
  XOR2_X1 u2_U506 (.Z( u2_FP_18 ) , .B( u2_L14_18 ) , .A( u2_out15_18 ) );
  XOR2_X1 u2_U508 (.Z( u2_FP_16 ) , .B( u2_L14_16 ) , .A( u2_out15_16 ) );
  XOR2_X1 u2_U51 (.B( u2_L0_24 ) , .Z( u2_N55 ) , .A( u2_out1_24 ) );
  XOR2_X1 u2_U511 (.Z( u2_FP_13 ) , .B( u2_L14_13 ) , .A( u2_out15_13 ) );
  XOR2_X1 u2_U514 (.Z( u2_FP_10 ) , .B( u2_L14_10 ) , .A( u2_out15_10 ) );
  XOR2_X1 u2_U55 (.B( u2_L0_20 ) , .Z( u2_N51 ) , .A( u2_out1_20 ) );
  XOR2_X1 u2_U58 (.B( u2_L0_18 ) , .Z( u2_N49 ) , .A( u2_out1_18 ) );
  XOR2_X1 u2_U62 (.B( u2_L13_30 ) , .Z( u2_N477 ) , .A( u2_out14_30 ) );
  XOR2_X1 u2_U65 (.B( u2_L13_27 ) , .Z( u2_N474 ) , .A( u2_out14_27 ) );
  XOR2_X1 u2_U66 (.B( u2_L13_26 ) , .Z( u2_N473 ) , .A( u2_out14_26 ) );
  XOR2_X1 u2_U68 (.B( u2_L13_24 ) , .Z( u2_N471 ) , .A( u2_out14_24 ) );
  XOR2_X1 u2_U70 (.B( u2_L0_16 ) , .Z( u2_N47 ) , .A( u2_out1_16 ) );
  XOR2_X1 u2_U72 (.B( u2_L13_21 ) , .Z( u2_N468 ) , .A( u2_out14_21 ) );
  XOR2_X1 u2_U73 (.B( u2_L13_20 ) , .Z( u2_N467 ) , .A( u2_out14_20 ) );
  XOR2_X1 u2_U77 (.B( u2_L13_16 ) , .Z( u2_N463 ) , .A( u2_out14_16 ) );
  XOR2_X1 u2_U78 (.B( u2_L13_15 ) , .Z( u2_N462 ) , .A( u2_out14_15 ) );
  XOR2_X1 u2_U84 (.B( u2_L13_10 ) , .Z( u2_N457 ) , .A( u2_out14_10 ) );
  XOR2_X1 u2_U88 (.B( u2_L13_6 ) , .Z( u2_N453 ) , .A( u2_out14_6 ) );
  XOR2_X1 u2_U89 (.B( u2_L13_5 ) , .Z( u2_N452 ) , .A( u2_out14_5 ) );
  XOR2_X1 u2_U94 (.B( u2_L13_1 ) , .Z( u2_N448 ) , .A( u2_out14_1 ) );
  XOR2_X1 u2_u0_U10 (.B( u2_K1_45 ) , .A( u2_desIn_r_41 ) , .Z( u2_u0_X_45 ) );
  XOR2_X1 u2_u0_U11 (.B( u2_K1_44 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_44 ) );
  XOR2_X1 u2_u0_U12 (.B( u2_K1_43 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_43 ) );
  XOR2_X1 u2_u0_U13 (.B( u2_K1_42 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_42 ) );
  XOR2_X1 u2_u0_U14 (.B( u2_K1_41 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_41 ) );
  XOR2_X1 u2_u0_U15 (.B( u2_K1_40 ) , .A( u2_desIn_r_17 ) , .Z( u2_u0_X_40 ) );
  XOR2_X1 u2_u0_U17 (.B( u2_K1_39 ) , .A( u2_desIn_r_9 ) , .Z( u2_u0_X_39 ) );
  XOR2_X1 u2_u0_U18 (.B( u2_K1_38 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_38 ) );
  XOR2_X1 u2_u0_U19 (.B( u2_K1_37 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_37 ) );
  XOR2_X1 u2_u0_U20 (.B( u2_K1_36 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_36 ) );
  XOR2_X1 u2_u0_U21 (.B( u2_K1_35 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_35 ) );
  XOR2_X1 u2_u0_U22 (.B( u2_K1_34 ) , .A( u2_desIn_r_51 ) , .Z( u2_u0_X_34 ) );
  XOR2_X1 u2_u0_U23 (.B( u2_K1_33 ) , .A( u2_desIn_r_43 ) , .Z( u2_u0_X_33 ) );
  XOR2_X1 u2_u0_U24 (.B( u2_K1_32 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_32 ) );
  XOR2_X1 u2_u0_U25 (.B( u2_K1_31 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_31 ) );
  XOR2_X1 u2_u0_U26 (.B( u2_K1_30 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_30 ) );
  XOR2_X1 u2_u0_U28 (.B( u2_K1_29 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_29 ) );
  XOR2_X1 u2_u0_U29 (.B( u2_K1_28 ) , .A( u2_desIn_r_19 ) , .Z( u2_u0_X_28 ) );
  XOR2_X1 u2_u0_U30 (.B( u2_K1_27 ) , .A( u2_desIn_r_11 ) , .Z( u2_u0_X_27 ) );
  XOR2_X1 u2_u0_U31 (.B( u2_K1_26 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_26 ) );
  XOR2_X1 u2_u0_U32 (.B( u2_K1_25 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_25 ) );
  XOR2_X1 u2_u0_U7 (.B( u2_K1_48 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_48 ) );
  XOR2_X1 u2_u0_U8 (.B( u2_K1_47 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_47 ) );
  XOR2_X1 u2_u0_U9 (.B( u2_K1_46 ) , .A( u2_desIn_r_49 ) , .Z( u2_u0_X_46 ) );
  OAI22_X1 u2_u0_u4_U10 (.B2( u2_u0_u4_n135 ) , .ZN( u2_u0_u4_n137 ) , .B1( u2_u0_u4_n153 ) , .A1( u2_u0_u4_n155 ) , .A2( u2_u0_u4_n171 ) );
  AND3_X1 u2_u0_u4_U11 (.A2( u2_u0_u4_n134 ) , .ZN( u2_u0_u4_n135 ) , .A3( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n157 ) );
  NAND2_X1 u2_u0_u4_U12 (.ZN( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n173 ) );
  AOI21_X1 u2_u0_u4_U13 (.B2( u2_u0_u4_n160 ) , .B1( u2_u0_u4_n161 ) , .ZN( u2_u0_u4_n162 ) , .A( u2_u0_u4_n170 ) );
  AOI21_X1 u2_u0_u4_U14 (.ZN( u2_u0_u4_n107 ) , .B2( u2_u0_u4_n143 ) , .A( u2_u0_u4_n174 ) , .B1( u2_u0_u4_n184 ) );
  AOI21_X1 u2_u0_u4_U15 (.B2( u2_u0_u4_n158 ) , .B1( u2_u0_u4_n159 ) , .ZN( u2_u0_u4_n163 ) , .A( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U16 (.A( u2_u0_u4_n153 ) , .B2( u2_u0_u4_n154 ) , .B1( u2_u0_u4_n155 ) , .ZN( u2_u0_u4_n165 ) );
  AOI21_X1 u2_u0_u4_U17 (.A( u2_u0_u4_n156 ) , .B2( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n164 ) , .B1( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U18 (.A( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n170 ) );
  AND2_X1 u2_u0_u4_U19 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n155 ) , .A1( u2_u0_u4_n160 ) );
  INV_X1 u2_u0_u4_U20 (.A( u2_u0_u4_n156 ) , .ZN( u2_u0_u4_n175 ) );
  NAND2_X1 u2_u0_u4_U21 (.A2( u2_u0_u4_n118 ) , .ZN( u2_u0_u4_n131 ) , .A1( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U22 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n130 ) );
  NAND2_X1 u2_u0_u4_U23 (.ZN( u2_u0_u4_n117 ) , .A2( u2_u0_u4_n118 ) , .A1( u2_u0_u4_n148 ) );
  NAND2_X1 u2_u0_u4_U24 (.ZN( u2_u0_u4_n129 ) , .A1( u2_u0_u4_n134 ) , .A2( u2_u0_u4_n148 ) );
  AND3_X1 u2_u0_u4_U25 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n143 ) , .A3( u2_u0_u4_n154 ) , .ZN( u2_u0_u4_n161 ) );
  AND2_X1 u2_u0_u4_U26 (.A1( u2_u0_u4_n145 ) , .A2( u2_u0_u4_n147 ) , .ZN( u2_u0_u4_n159 ) );
  OR3_X1 u2_u0_u4_U27 (.A3( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n115 ) , .A1( u2_u0_u4_n116 ) , .ZN( u2_u0_u4_n136 ) );
  AOI21_X1 u2_u0_u4_U28 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n116 ) , .B2( u2_u0_u4_n173 ) , .B1( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U29 (.ZN( u2_u0_u4_n115 ) , .B2( u2_u0_u4_n145 ) , .B1( u2_u0_u4_n146 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U3 (.ZN( u2_u0_u4_n121 ) , .A1( u2_u0_u4_n181 ) , .A2( u2_u0_u4_n182 ) );
  OAI22_X1 u2_u0_u4_U30 (.ZN( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n121 ) , .B1( u2_u0_u4_n160 ) , .B2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n171 ) );
  INV_X1 u2_u0_u4_U31 (.A( u2_u0_u4_n158 ) , .ZN( u2_u0_u4_n182 ) );
  INV_X1 u2_u0_u4_U32 (.ZN( u2_u0_u4_n181 ) , .A( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U33 (.A( u2_u0_u4_n144 ) , .ZN( u2_u0_u4_n179 ) );
  INV_X1 u2_u0_u4_U34 (.A( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n178 ) );
  NAND2_X1 u2_u0_u4_U35 (.A2( u2_u0_u4_n154 ) , .A1( u2_u0_u4_n96 ) , .ZN( u2_u0_u4_n97 ) );
  INV_X1 u2_u0_u4_U36 (.ZN( u2_u0_u4_n186 ) , .A( u2_u0_u4_n95 ) );
  OAI221_X1 u2_u0_u4_U37 (.C1( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n158 ) , .B2( u2_u0_u4_n171 ) , .C2( u2_u0_u4_n173 ) , .A( u2_u0_u4_n94 ) , .ZN( u2_u0_u4_n95 ) );
  AOI222_X1 u2_u0_u4_U38 (.B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n138 ) , .C2( u2_u0_u4_n175 ) , .A2( u2_u0_u4_n179 ) , .C1( u2_u0_u4_n181 ) , .B1( u2_u0_u4_n185 ) , .ZN( u2_u0_u4_n94 ) );
  INV_X1 u2_u0_u4_U39 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n185 ) );
  INV_X1 u2_u0_u4_U4 (.A( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U40 (.A( u2_u0_u4_n143 ) , .ZN( u2_u0_u4_n183 ) );
  NOR2_X1 u2_u0_u4_U41 (.ZN( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n168 ) , .A2( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U42 (.A1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n153 ) );
  NOR2_X1 u2_u0_u4_U43 (.A2( u2_u0_u4_n128 ) , .A1( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n156 ) );
  AOI22_X1 u2_u0_u4_U44 (.B2( u2_u0_u4_n122 ) , .A1( u2_u0_u4_n123 ) , .ZN( u2_u0_u4_n124 ) , .B1( u2_u0_u4_n128 ) , .A2( u2_u0_u4_n172 ) );
  INV_X1 u2_u0_u4_U45 (.A( u2_u0_u4_n153 ) , .ZN( u2_u0_u4_n172 ) );
  NAND2_X1 u2_u0_u4_U46 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n123 ) , .A1( u2_u0_u4_n161 ) );
  AOI22_X1 u2_u0_u4_U47 (.B2( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n133 ) , .ZN( u2_u0_u4_n140 ) , .A1( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n179 ) );
  NAND2_X1 u2_u0_u4_U48 (.ZN( u2_u0_u4_n133 ) , .A2( u2_u0_u4_n146 ) , .A1( u2_u0_u4_n154 ) );
  NAND2_X1 u2_u0_u4_U49 (.A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n154 ) , .A2( u2_u0_u4_n98 ) );
  NOR4_X1 u2_u0_u4_U5 (.A4( u2_u0_u4_n106 ) , .A3( u2_u0_u4_n107 ) , .A2( u2_u0_u4_n108 ) , .A1( u2_u0_u4_n109 ) , .ZN( u2_u0_u4_n110 ) );
  NAND2_X1 u2_u0_u4_U50 (.A1( u2_u0_u4_n101 ) , .ZN( u2_u0_u4_n158 ) , .A2( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U51 (.ZN( u2_u0_u4_n127 ) , .A( u2_u0_u4_n136 ) , .B2( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n180 ) );
  INV_X1 u2_u0_u4_U52 (.A( u2_u0_u4_n160 ) , .ZN( u2_u0_u4_n180 ) );
  NAND2_X1 u2_u0_u4_U53 (.A2( u2_u0_u4_n104 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n146 ) );
  NAND2_X1 u2_u0_u4_U54 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n160 ) );
  NAND2_X1 u2_u0_u4_U55 (.ZN( u2_u0_u4_n134 ) , .A1( u2_u0_u4_n98 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U56 (.A1( u2_u0_u4_n103 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n143 ) );
  NAND2_X1 u2_u0_u4_U57 (.A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U58 (.A1( u2_u0_u4_n100 ) , .A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n120 ) );
  NAND2_X1 u2_u0_u4_U59 (.A1( u2_u0_u4_n102 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n148 ) );
  AOI21_X1 u2_u0_u4_U6 (.ZN( u2_u0_u4_n106 ) , .B2( u2_u0_u4_n146 ) , .B1( u2_u0_u4_n158 ) , .A( u2_u0_u4_n170 ) );
  NAND2_X1 u2_u0_u4_U60 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n157 ) );
  INV_X1 u2_u0_u4_U61 (.A( u2_u0_u4_n150 ) , .ZN( u2_u0_u4_n173 ) );
  INV_X1 u2_u0_u4_U62 (.A( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n171 ) );
  NAND2_X1 u2_u0_u4_U63 (.A1( u2_u0_u4_n100 ) , .ZN( u2_u0_u4_n118 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U64 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n144 ) );
  NAND2_X1 u2_u0_u4_U65 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U66 (.A( u2_u0_u4_n128 ) , .ZN( u2_u0_u4_n174 ) );
  NAND2_X1 u2_u0_u4_U67 (.A2( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n119 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U68 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U69 (.A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n113 ) , .A1( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U7 (.ZN( u2_u0_u4_n108 ) , .B2( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n155 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U70 (.A2( u2_u0_X_28 ) , .ZN( u2_u0_u4_n150 ) , .A1( u2_u0_u4_n168 ) );
  NOR2_X1 u2_u0_u4_U71 (.A2( u2_u0_X_29 ) , .ZN( u2_u0_u4_n152 ) , .A1( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U72 (.A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n105 ) , .A1( u2_u0_u4_n176 ) );
  NOR2_X1 u2_u0_u4_U73 (.A2( u2_u0_X_26 ) , .ZN( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n177 ) );
  NOR2_X1 u2_u0_u4_U74 (.A2( u2_u0_X_28 ) , .A1( u2_u0_X_29 ) , .ZN( u2_u0_u4_n128 ) );
  NOR2_X1 u2_u0_u4_U75 (.A2( u2_u0_X_27 ) , .A1( u2_u0_X_30 ) , .ZN( u2_u0_u4_n102 ) );
  NOR2_X1 u2_u0_u4_U76 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n98 ) );
  AND2_X1 u2_u0_u4_U77 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n104 ) );
  AND2_X1 u2_u0_u4_U78 (.A1( u2_u0_X_30 ) , .A2( u2_u0_u4_n176 ) , .ZN( u2_u0_u4_n99 ) );
  AND2_X1 u2_u0_u4_U79 (.A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n101 ) , .A2( u2_u0_u4_n177 ) );
  AOI21_X1 u2_u0_u4_U8 (.ZN( u2_u0_u4_n109 ) , .A( u2_u0_u4_n153 ) , .B1( u2_u0_u4_n159 ) , .B2( u2_u0_u4_n184 ) );
  AND2_X1 u2_u0_u4_U80 (.A1( u2_u0_X_27 ) , .A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n103 ) );
  INV_X1 u2_u0_u4_U81 (.A( u2_u0_X_28 ) , .ZN( u2_u0_u4_n169 ) );
  INV_X1 u2_u0_u4_U82 (.A( u2_u0_X_29 ) , .ZN( u2_u0_u4_n168 ) );
  INV_X1 u2_u0_u4_U83 (.A( u2_u0_X_25 ) , .ZN( u2_u0_u4_n177 ) );
  INV_X1 u2_u0_u4_U84 (.A( u2_u0_X_27 ) , .ZN( u2_u0_u4_n176 ) );
  NAND4_X1 u2_u0_u4_U85 (.ZN( u2_out0_25 ) , .A4( u2_u0_u4_n139 ) , .A3( u2_u0_u4_n140 ) , .A2( u2_u0_u4_n141 ) , .A1( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U86 (.A( u2_u0_u4_n128 ) , .B2( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n130 ) , .ZN( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U87 (.B2( u2_u0_u4_n131 ) , .ZN( u2_u0_u4_n141 ) , .A( u2_u0_u4_n175 ) , .B1( u2_u0_u4_n183 ) );
  NAND4_X1 u2_u0_u4_U88 (.ZN( u2_out0_14 ) , .A4( u2_u0_u4_n124 ) , .A3( u2_u0_u4_n125 ) , .A2( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n127 ) );
  AOI22_X1 u2_u0_u4_U89 (.B2( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n152 ) , .A2( u2_u0_u4_n175 ) );
  AOI211_X1 u2_u0_u4_U9 (.B( u2_u0_u4_n136 ) , .A( u2_u0_u4_n137 ) , .C2( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n139 ) , .C1( u2_u0_u4_n182 ) );
  AOI22_X1 u2_u0_u4_U90 (.ZN( u2_u0_u4_n125 ) , .B2( u2_u0_u4_n131 ) , .A2( u2_u0_u4_n132 ) , .B1( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n178 ) );
  NAND4_X1 u2_u0_u4_U91 (.ZN( u2_out0_8 ) , .A4( u2_u0_u4_n110 ) , .A3( u2_u0_u4_n111 ) , .A2( u2_u0_u4_n112 ) , .A1( u2_u0_u4_n186 ) );
  NAND2_X1 u2_u0_u4_U92 (.ZN( u2_u0_u4_n112 ) , .A2( u2_u0_u4_n130 ) , .A1( u2_u0_u4_n150 ) );
  AOI22_X1 u2_u0_u4_U93 (.ZN( u2_u0_u4_n111 ) , .B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n152 ) , .B1( u2_u0_u4_n178 ) , .A2( u2_u0_u4_n97 ) );
  AOI22_X1 u2_u0_u4_U94 (.B2( u2_u0_u4_n149 ) , .B1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n151 ) , .A1( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n167 ) );
  NOR4_X1 u2_u0_u4_U95 (.A4( u2_u0_u4_n162 ) , .A3( u2_u0_u4_n163 ) , .A2( u2_u0_u4_n164 ) , .A1( u2_u0_u4_n165 ) , .ZN( u2_u0_u4_n166 ) );
  NAND3_X1 u2_u0_u4_U96 (.ZN( u2_out0_3 ) , .A3( u2_u0_u4_n166 ) , .A1( u2_u0_u4_n167 ) , .A2( u2_u0_u4_n186 ) );
  NAND3_X1 u2_u0_u4_U97 (.A3( u2_u0_u4_n146 ) , .A2( u2_u0_u4_n147 ) , .A1( u2_u0_u4_n148 ) , .ZN( u2_u0_u4_n149 ) );
  NAND3_X1 u2_u0_u4_U98 (.A3( u2_u0_u4_n143 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n145 ) , .ZN( u2_u0_u4_n151 ) );
  NAND3_X1 u2_u0_u4_U99 (.A3( u2_u0_u4_n121 ) , .ZN( u2_u0_u4_n122 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n154 ) );
  INV_X1 u2_u0_u5_U10 (.A( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U100 (.A3( u2_u0_u5_n141 ) , .A1( u2_u0_u5_n142 ) , .ZN( u2_u0_u5_n143 ) , .A2( u2_u0_u5_n191 ) );
  NAND4_X1 u2_u0_u5_U101 (.ZN( u2_out0_4 ) , .A4( u2_u0_u5_n112 ) , .A2( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n114 ) , .A3( u2_u0_u5_n195 ) );
  AOI211_X1 u2_u0_u5_U102 (.A( u2_u0_u5_n110 ) , .C1( u2_u0_u5_n111 ) , .ZN( u2_u0_u5_n112 ) , .B( u2_u0_u5_n118 ) , .C2( u2_u0_u5_n177 ) );
  AOI222_X1 u2_u0_u5_U103 (.ZN( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n131 ) , .C1( u2_u0_u5_n148 ) , .B2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n178 ) , .A2( u2_u0_u5_n179 ) , .B1( u2_u0_u5_n99 ) );
  NAND3_X1 u2_u0_u5_U104 (.A2( u2_u0_u5_n154 ) , .A3( u2_u0_u5_n158 ) , .A1( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n99 ) );
  NOR2_X1 u2_u0_u5_U11 (.ZN( u2_u0_u5_n160 ) , .A2( u2_u0_u5_n173 ) , .A1( u2_u0_u5_n177 ) );
  INV_X1 u2_u0_u5_U12 (.A( u2_u0_u5_n150 ) , .ZN( u2_u0_u5_n174 ) );
  AOI21_X1 u2_u0_u5_U13 (.A( u2_u0_u5_n160 ) , .B2( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n162 ) , .B1( u2_u0_u5_n192 ) );
  INV_X1 u2_u0_u5_U14 (.A( u2_u0_u5_n159 ) , .ZN( u2_u0_u5_n192 ) );
  AOI21_X1 u2_u0_u5_U15 (.A( u2_u0_u5_n156 ) , .B2( u2_u0_u5_n157 ) , .B1( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n163 ) );
  AOI21_X1 u2_u0_u5_U16 (.B2( u2_u0_u5_n139 ) , .B1( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n141 ) , .A( u2_u0_u5_n150 ) );
  OAI21_X1 u2_u0_u5_U17 (.A( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n134 ) , .B1( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n142 ) );
  OAI21_X1 u2_u0_u5_U18 (.ZN( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n147 ) , .A( u2_u0_u5_n173 ) , .B1( u2_u0_u5_n188 ) );
  NAND2_X1 u2_u0_u5_U19 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n137 ) );
  INV_X1 u2_u0_u5_U20 (.A( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n194 ) );
  NAND2_X1 u2_u0_u5_U21 (.A1( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n132 ) , .A2( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U22 (.A2( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n136 ) , .A1( u2_u0_u5_n154 ) );
  NAND2_X1 u2_u0_u5_U23 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n159 ) );
  INV_X1 u2_u0_u5_U24 (.A( u2_u0_u5_n156 ) , .ZN( u2_u0_u5_n175 ) );
  INV_X1 u2_u0_u5_U25 (.A( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n188 ) );
  INV_X1 u2_u0_u5_U26 (.A( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n179 ) );
  INV_X1 u2_u0_u5_U27 (.A( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n182 ) );
  INV_X1 u2_u0_u5_U28 (.A( u2_u0_u5_n151 ) , .ZN( u2_u0_u5_n183 ) );
  INV_X1 u2_u0_u5_U29 (.A( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U3 (.ZN( u2_u0_u5_n134 ) , .A1( u2_u0_u5_n183 ) , .A2( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U30 (.A( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n184 ) );
  INV_X1 u2_u0_u5_U31 (.A( u2_u0_u5_n139 ) , .ZN( u2_u0_u5_n189 ) );
  INV_X1 u2_u0_u5_U32 (.A( u2_u0_u5_n157 ) , .ZN( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U33 (.A( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n193 ) );
  NAND2_X1 u2_u0_u5_U34 (.ZN( u2_u0_u5_n111 ) , .A1( u2_u0_u5_n140 ) , .A2( u2_u0_u5_n155 ) );
  NOR2_X1 u2_u0_u5_U35 (.ZN( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n170 ) , .A2( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U36 (.A( u2_u0_u5_n117 ) , .ZN( u2_u0_u5_n196 ) );
  OAI221_X1 u2_u0_u5_U37 (.A( u2_u0_u5_n116 ) , .ZN( u2_u0_u5_n117 ) , .B2( u2_u0_u5_n119 ) , .C1( u2_u0_u5_n153 ) , .C2( u2_u0_u5_n158 ) , .B1( u2_u0_u5_n172 ) );
  AOI222_X1 u2_u0_u5_U38 (.ZN( u2_u0_u5_n116 ) , .B2( u2_u0_u5_n145 ) , .C1( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n177 ) , .B1( u2_u0_u5_n187 ) , .A1( u2_u0_u5_n193 ) );
  INV_X1 u2_u0_u5_U39 (.A( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n187 ) );
  INV_X1 u2_u0_u5_U4 (.A( u2_u0_u5_n138 ) , .ZN( u2_u0_u5_n191 ) );
  AOI22_X1 u2_u0_u5_U40 (.B2( u2_u0_u5_n131 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n169 ) , .B1( u2_u0_u5_n174 ) , .A1( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U41 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n173 ) );
  AOI21_X1 u2_u0_u5_U42 (.A( u2_u0_u5_n118 ) , .B2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n168 ) , .B1( u2_u0_u5_n186 ) );
  INV_X1 u2_u0_u5_U43 (.A( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n186 ) );
  NOR2_X1 u2_u0_u5_U44 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n152 ) , .A2( u2_u0_u5_n176 ) );
  NOR2_X1 u2_u0_u5_U45 (.A1( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n118 ) , .A2( u2_u0_u5_n153 ) );
  NOR2_X1 u2_u0_u5_U46 (.A2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n156 ) , .A1( u2_u0_u5_n174 ) );
  NOR2_X1 u2_u0_u5_U47 (.ZN( u2_u0_u5_n121 ) , .A2( u2_u0_u5_n145 ) , .A1( u2_u0_u5_n176 ) );
  AOI22_X1 u2_u0_u5_U48 (.ZN( u2_u0_u5_n114 ) , .A2( u2_u0_u5_n137 ) , .A1( u2_u0_u5_n145 ) , .B2( u2_u0_u5_n175 ) , .B1( u2_u0_u5_n193 ) );
  OAI211_X1 u2_u0_u5_U49 (.B( u2_u0_u5_n124 ) , .A( u2_u0_u5_n125 ) , .C2( u2_u0_u5_n126 ) , .C1( u2_u0_u5_n127 ) , .ZN( u2_u0_u5_n128 ) );
  OAI21_X1 u2_u0_u5_U5 (.B2( u2_u0_u5_n136 ) , .B1( u2_u0_u5_n137 ) , .ZN( u2_u0_u5_n138 ) , .A( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U50 (.ZN( u2_u0_u5_n127 ) , .A1( u2_u0_u5_n136 ) , .A3( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n182 ) );
  OAI21_X1 u2_u0_u5_U51 (.ZN( u2_u0_u5_n124 ) , .A( u2_u0_u5_n177 ) , .B2( u2_u0_u5_n183 ) , .B1( u2_u0_u5_n189 ) );
  OAI21_X1 u2_u0_u5_U52 (.ZN( u2_u0_u5_n125 ) , .A( u2_u0_u5_n174 ) , .B2( u2_u0_u5_n185 ) , .B1( u2_u0_u5_n190 ) );
  AOI21_X1 u2_u0_u5_U53 (.A( u2_u0_u5_n153 ) , .B2( u2_u0_u5_n154 ) , .B1( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n164 ) );
  AOI21_X1 u2_u0_u5_U54 (.ZN( u2_u0_u5_n110 ) , .B1( u2_u0_u5_n122 ) , .B2( u2_u0_u5_n139 ) , .A( u2_u0_u5_n153 ) );
  INV_X1 u2_u0_u5_U55 (.A( u2_u0_u5_n153 ) , .ZN( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U56 (.A( u2_u0_u5_n126 ) , .ZN( u2_u0_u5_n173 ) );
  AND2_X1 u2_u0_u5_U57 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n147 ) );
  AND2_X1 u2_u0_u5_U58 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n148 ) );
  NAND2_X1 u2_u0_u5_U59 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n158 ) );
  INV_X1 u2_u0_u5_U6 (.A( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n178 ) );
  NAND2_X1 u2_u0_u5_U60 (.A2( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n139 ) );
  NAND2_X1 u2_u0_u5_U61 (.A1( u2_u0_u5_n106 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n119 ) );
  NAND2_X1 u2_u0_u5_U62 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n140 ) );
  NAND2_X1 u2_u0_u5_U63 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n155 ) );
  NAND2_X1 u2_u0_u5_U64 (.A2( u2_u0_u5_n106 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n122 ) );
  NAND2_X1 u2_u0_u5_U65 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n115 ) );
  NAND2_X1 u2_u0_u5_U66 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n103 ) , .ZN( u2_u0_u5_n161 ) );
  NAND2_X1 u2_u0_u5_U67 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n154 ) );
  INV_X1 u2_u0_u5_U68 (.A( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U69 (.A1( u2_u0_u5_n103 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n123 ) );
  OAI22_X1 u2_u0_u5_U7 (.B2( u2_u0_u5_n149 ) , .B1( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n151 ) , .A1( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n165 ) );
  NAND2_X1 u2_u0_u5_U70 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n151 ) );
  NAND2_X1 u2_u0_u5_U71 (.A2( u2_u0_u5_n107 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n120 ) );
  NAND2_X1 u2_u0_u5_U72 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n157 ) );
  AND2_X1 u2_u0_u5_U73 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n104 ) , .ZN( u2_u0_u5_n131 ) );
  INV_X1 u2_u0_u5_U74 (.A( u2_u0_u5_n102 ) , .ZN( u2_u0_u5_n195 ) );
  OAI221_X1 u2_u0_u5_U75 (.A( u2_u0_u5_n101 ) , .ZN( u2_u0_u5_n102 ) , .C2( u2_u0_u5_n115 ) , .C1( u2_u0_u5_n126 ) , .B1( u2_u0_u5_n134 ) , .B2( u2_u0_u5_n160 ) );
  OAI21_X1 u2_u0_u5_U76 (.ZN( u2_u0_u5_n101 ) , .B1( u2_u0_u5_n137 ) , .A( u2_u0_u5_n146 ) , .B2( u2_u0_u5_n147 ) );
  NOR2_X1 u2_u0_u5_U77 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n145 ) );
  NOR2_X1 u2_u0_u5_U78 (.A2( u2_u0_X_34 ) , .ZN( u2_u0_u5_n146 ) , .A1( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U79 (.A2( u2_u0_X_31 ) , .A1( u2_u0_X_32 ) , .ZN( u2_u0_u5_n103 ) );
  NOR3_X1 u2_u0_u5_U8 (.A2( u2_u0_u5_n147 ) , .A1( u2_u0_u5_n148 ) , .ZN( u2_u0_u5_n149 ) , .A3( u2_u0_u5_n194 ) );
  NOR2_X1 u2_u0_u5_U80 (.A2( u2_u0_X_36 ) , .ZN( u2_u0_u5_n105 ) , .A1( u2_u0_u5_n180 ) );
  NOR2_X1 u2_u0_u5_U81 (.A2( u2_u0_X_33 ) , .ZN( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n170 ) );
  NOR2_X1 u2_u0_u5_U82 (.A2( u2_u0_X_33 ) , .A1( u2_u0_X_36 ) , .ZN( u2_u0_u5_n107 ) );
  NOR2_X1 u2_u0_u5_U83 (.A2( u2_u0_X_31 ) , .ZN( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n181 ) );
  NAND2_X1 u2_u0_u5_U84 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n153 ) );
  NAND2_X1 u2_u0_u5_U85 (.A1( u2_u0_X_34 ) , .ZN( u2_u0_u5_n126 ) , .A2( u2_u0_u5_n171 ) );
  AND2_X1 u2_u0_u5_U86 (.A1( u2_u0_X_31 ) , .A2( u2_u0_X_32 ) , .ZN( u2_u0_u5_n106 ) );
  AND2_X1 u2_u0_u5_U87 (.A1( u2_u0_X_31 ) , .ZN( u2_u0_u5_n109 ) , .A2( u2_u0_u5_n181 ) );
  INV_X1 u2_u0_u5_U88 (.A( u2_u0_X_33 ) , .ZN( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U89 (.A( u2_u0_X_35 ) , .ZN( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U9 (.ZN( u2_u0_u5_n135 ) , .A1( u2_u0_u5_n173 ) , .A2( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U90 (.A( u2_u0_X_36 ) , .ZN( u2_u0_u5_n170 ) );
  INV_X1 u2_u0_u5_U91 (.A( u2_u0_X_32 ) , .ZN( u2_u0_u5_n181 ) );
  NAND4_X1 u2_u0_u5_U92 (.ZN( u2_out0_29 ) , .A4( u2_u0_u5_n129 ) , .A3( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n196 ) );
  AOI221_X1 u2_u0_u5_U93 (.A( u2_u0_u5_n128 ) , .ZN( u2_u0_u5_n129 ) , .C2( u2_u0_u5_n132 ) , .B2( u2_u0_u5_n159 ) , .B1( u2_u0_u5_n176 ) , .C1( u2_u0_u5_n184 ) );
  AOI222_X1 u2_u0_u5_U94 (.ZN( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n146 ) , .B1( u2_u0_u5_n147 ) , .C2( u2_u0_u5_n175 ) , .B2( u2_u0_u5_n179 ) , .A1( u2_u0_u5_n188 ) , .C1( u2_u0_u5_n194 ) );
  NAND4_X1 u2_u0_u5_U95 (.ZN( u2_out0_19 ) , .A4( u2_u0_u5_n166 ) , .A3( u2_u0_u5_n167 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n169 ) );
  AOI22_X1 u2_u0_u5_U96 (.B2( u2_u0_u5_n145 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n167 ) , .B1( u2_u0_u5_n182 ) , .A1( u2_u0_u5_n189 ) );
  NOR4_X1 u2_u0_u5_U97 (.A4( u2_u0_u5_n162 ) , .A3( u2_u0_u5_n163 ) , .A2( u2_u0_u5_n164 ) , .A1( u2_u0_u5_n165 ) , .ZN( u2_u0_u5_n166 ) );
  NAND4_X1 u2_u0_u5_U98 (.ZN( u2_out0_11 ) , .A4( u2_u0_u5_n143 ) , .A3( u2_u0_u5_n144 ) , .A2( u2_u0_u5_n169 ) , .A1( u2_u0_u5_n196 ) );
  AOI22_X1 u2_u0_u5_U99 (.A2( u2_u0_u5_n132 ) , .ZN( u2_u0_u5_n144 ) , .B2( u2_u0_u5_n145 ) , .B1( u2_u0_u5_n184 ) , .A1( u2_u0_u5_n194 ) );
  AOI22_X1 u2_u0_u6_U10 (.A2( u2_u0_u6_n151 ) , .B2( u2_u0_u6_n161 ) , .A1( u2_u0_u6_n167 ) , .B1( u2_u0_u6_n170 ) , .ZN( u2_u0_u6_n89 ) );
  AOI21_X1 u2_u0_u6_U11 (.B1( u2_u0_u6_n107 ) , .B2( u2_u0_u6_n132 ) , .A( u2_u0_u6_n158 ) , .ZN( u2_u0_u6_n88 ) );
  AOI21_X1 u2_u0_u6_U12 (.B2( u2_u0_u6_n147 ) , .B1( u2_u0_u6_n148 ) , .ZN( u2_u0_u6_n149 ) , .A( u2_u0_u6_n158 ) );
  AOI21_X1 u2_u0_u6_U13 (.ZN( u2_u0_u6_n106 ) , .A( u2_u0_u6_n142 ) , .B2( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n164 ) );
  INV_X1 u2_u0_u6_U14 (.A( u2_u0_u6_n155 ) , .ZN( u2_u0_u6_n161 ) );
  INV_X1 u2_u0_u6_U15 (.A( u2_u0_u6_n128 ) , .ZN( u2_u0_u6_n164 ) );
  NAND2_X1 u2_u0_u6_U16 (.ZN( u2_u0_u6_n110 ) , .A1( u2_u0_u6_n122 ) , .A2( u2_u0_u6_n129 ) );
  NAND2_X1 u2_u0_u6_U17 (.ZN( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n146 ) , .A1( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U18 (.A( u2_u0_u6_n132 ) , .ZN( u2_u0_u6_n171 ) );
  AND2_X1 u2_u0_u6_U19 (.A1( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n147 ) );
  INV_X1 u2_u0_u6_U20 (.A( u2_u0_u6_n127 ) , .ZN( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U21 (.A( u2_u0_u6_n121 ) , .ZN( u2_u0_u6_n167 ) );
  INV_X1 u2_u0_u6_U22 (.A( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U23 (.A( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n170 ) );
  INV_X1 u2_u0_u6_U24 (.A( u2_u0_u6_n113 ) , .ZN( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U25 (.A1( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n119 ) , .ZN( u2_u0_u6_n133 ) );
  AND2_X1 u2_u0_u6_U26 (.A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n122 ) , .ZN( u2_u0_u6_n131 ) );
  AND3_X1 u2_u0_u6_U27 (.ZN( u2_u0_u6_n120 ) , .A2( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n132 ) , .A3( u2_u0_u6_n145 ) );
  INV_X1 u2_u0_u6_U28 (.A( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n163 ) );
  AOI222_X1 u2_u0_u6_U29 (.ZN( u2_u0_u6_n114 ) , .A1( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n126 ) , .B2( u2_u0_u6_n151 ) , .C2( u2_u0_u6_n159 ) , .C1( u2_u0_u6_n168 ) , .B1( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U3 (.A( u2_u0_u6_n110 ) , .ZN( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U30 (.A1( u2_u0_u6_n162 ) , .A2( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n98 ) );
  AOI211_X1 u2_u0_u6_U31 (.B( u2_u0_u6_n134 ) , .A( u2_u0_u6_n135 ) , .C1( u2_u0_u6_n136 ) , .ZN( u2_u0_u6_n137 ) , .C2( u2_u0_u6_n151 ) );
  AOI21_X1 u2_u0_u6_U32 (.B2( u2_u0_u6_n132 ) , .B1( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n134 ) , .A( u2_u0_u6_n158 ) );
  NAND4_X1 u2_u0_u6_U33 (.A4( u2_u0_u6_n127 ) , .A3( u2_u0_u6_n128 ) , .A2( u2_u0_u6_n129 ) , .A1( u2_u0_u6_n130 ) , .ZN( u2_u0_u6_n136 ) );
  AOI21_X1 u2_u0_u6_U34 (.B1( u2_u0_u6_n131 ) , .ZN( u2_u0_u6_n135 ) , .A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n146 ) );
  NAND2_X1 u2_u0_u6_U35 (.A1( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U36 (.ZN( u2_u0_u6_n132 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n97 ) );
  AOI22_X1 u2_u0_u6_U37 (.B2( u2_u0_u6_n110 ) , .B1( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n112 ) , .ZN( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n161 ) );
  NAND4_X1 u2_u0_u6_U38 (.A3( u2_u0_u6_n109 ) , .ZN( u2_u0_u6_n112 ) , .A4( u2_u0_u6_n132 ) , .A2( u2_u0_u6_n147 ) , .A1( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U39 (.ZN( u2_u0_u6_n109 ) , .A1( u2_u0_u6_n170 ) , .A2( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U4 (.A( u2_u0_u6_n142 ) , .ZN( u2_u0_u6_n174 ) );
  NOR2_X1 u2_u0_u6_U40 (.A2( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n155 ) , .A1( u2_u0_u6_n160 ) );
  NAND2_X1 u2_u0_u6_U41 (.ZN( u2_u0_u6_n146 ) , .A2( u2_u0_u6_n94 ) , .A1( u2_u0_u6_n99 ) );
  AOI21_X1 u2_u0_u6_U42 (.A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n145 ) , .B1( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n150 ) );
  INV_X1 u2_u0_u6_U43 (.A( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U44 (.ZN( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n92 ) );
  NAND2_X1 u2_u0_u6_U45 (.ZN( u2_u0_u6_n129 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n96 ) );
  INV_X1 u2_u0_u6_U46 (.A( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n159 ) );
  NAND2_X1 u2_u0_u6_U47 (.ZN( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n97 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U48 (.ZN( u2_u0_u6_n148 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n94 ) );
  NAND2_X1 u2_u0_u6_U49 (.ZN( u2_u0_u6_n108 ) , .A2( u2_u0_u6_n139 ) , .A1( u2_u0_u6_n144 ) );
  NAND2_X1 u2_u0_u6_U5 (.A2( u2_u0_u6_n143 ) , .ZN( u2_u0_u6_n152 ) , .A1( u2_u0_u6_n166 ) );
  NAND2_X1 u2_u0_u6_U50 (.ZN( u2_u0_u6_n121 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n97 ) );
  NAND2_X1 u2_u0_u6_U51 (.ZN( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n95 ) );
  AND2_X1 u2_u0_u6_U52 (.ZN( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U53 (.ZN( u2_u0_u6_n147 ) , .A2( u2_u0_u6_n98 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U54 (.ZN( u2_u0_u6_n128 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U55 (.ZN( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U56 (.ZN( u2_u0_u6_n123 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U57 (.ZN( u2_u0_u6_n100 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U58 (.ZN( u2_u0_u6_n122 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n97 ) );
  INV_X1 u2_u0_u6_U59 (.A( u2_u0_u6_n139 ) , .ZN( u2_u0_u6_n160 ) );
  AOI22_X1 u2_u0_u6_U6 (.B2( u2_u0_u6_n101 ) , .A1( u2_u0_u6_n102 ) , .ZN( u2_u0_u6_n103 ) , .B1( u2_u0_u6_n160 ) , .A2( u2_u0_u6_n161 ) );
  NAND2_X1 u2_u0_u6_U60 (.ZN( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n96 ) , .A2( u2_u0_u6_n98 ) );
  NOR2_X1 u2_u0_u6_U61 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n126 ) );
  NOR2_X1 u2_u0_u6_U62 (.A2( u2_u0_X_39 ) , .A1( u2_u0_X_42 ) , .ZN( u2_u0_u6_n92 ) );
  NOR2_X1 u2_u0_u6_U63 (.A2( u2_u0_X_39 ) , .A1( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n97 ) );
  NOR2_X1 u2_u0_u6_U64 (.A2( u2_u0_X_38 ) , .A1( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n95 ) );
  NOR2_X1 u2_u0_u6_U65 (.A2( u2_u0_X_41 ) , .ZN( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n157 ) );
  NOR2_X1 u2_u0_u6_U66 (.A2( u2_u0_X_37 ) , .A1( u2_u0_u6_n162 ) , .ZN( u2_u0_u6_n94 ) );
  NOR2_X1 u2_u0_u6_U67 (.A2( u2_u0_X_37 ) , .A1( u2_u0_X_38 ) , .ZN( u2_u0_u6_n91 ) );
  NAND2_X1 u2_u0_u6_U68 (.A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n144 ) , .A2( u2_u0_u6_n157 ) );
  NAND2_X1 u2_u0_u6_U69 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n139 ) );
  NOR2_X1 u2_u0_u6_U7 (.A1( u2_u0_u6_n118 ) , .ZN( u2_u0_u6_n143 ) , .A2( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U70 (.A1( u2_u0_X_39 ) , .A2( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n96 ) );
  AND2_X1 u2_u0_u6_U71 (.A1( u2_u0_X_39 ) , .A2( u2_u0_X_42 ) , .ZN( u2_u0_u6_n99 ) );
  INV_X1 u2_u0_u6_U72 (.A( u2_u0_X_40 ) , .ZN( u2_u0_u6_n157 ) );
  INV_X1 u2_u0_u6_U73 (.A( u2_u0_X_37 ) , .ZN( u2_u0_u6_n165 ) );
  INV_X1 u2_u0_u6_U74 (.A( u2_u0_X_38 ) , .ZN( u2_u0_u6_n162 ) );
  INV_X1 u2_u0_u6_U75 (.A( u2_u0_X_42 ) , .ZN( u2_u0_u6_n156 ) );
  NAND4_X1 u2_u0_u6_U76 (.ZN( u2_out0_32 ) , .A4( u2_u0_u6_n103 ) , .A3( u2_u0_u6_n104 ) , .A2( u2_u0_u6_n105 ) , .A1( u2_u0_u6_n106 ) );
  AOI22_X1 u2_u0_u6_U77 (.ZN( u2_u0_u6_n105 ) , .A2( u2_u0_u6_n108 ) , .A1( u2_u0_u6_n118 ) , .B2( u2_u0_u6_n126 ) , .B1( u2_u0_u6_n171 ) );
  AOI22_X1 u2_u0_u6_U78 (.ZN( u2_u0_u6_n104 ) , .A1( u2_u0_u6_n111 ) , .B1( u2_u0_u6_n124 ) , .B2( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n93 ) );
  NAND4_X1 u2_u0_u6_U79 (.ZN( u2_out0_12 ) , .A4( u2_u0_u6_n114 ) , .A3( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n116 ) , .A1( u2_u0_u6_n117 ) );
  OAI21_X1 u2_u0_u6_U8 (.A( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n169 ) , .B2( u2_u0_u6_n173 ) , .ZN( u2_u0_u6_n90 ) );
  OAI22_X1 u2_u0_u6_U80 (.B2( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n116 ) , .B1( u2_u0_u6_n126 ) , .A2( u2_u0_u6_n164 ) , .A1( u2_u0_u6_n167 ) );
  OAI21_X1 u2_u0_u6_U81 (.A( u2_u0_u6_n108 ) , .ZN( u2_u0_u6_n117 ) , .B2( u2_u0_u6_n141 ) , .B1( u2_u0_u6_n163 ) );
  OAI211_X1 u2_u0_u6_U82 (.ZN( u2_out0_7 ) , .B( u2_u0_u6_n153 ) , .C2( u2_u0_u6_n154 ) , .C1( u2_u0_u6_n155 ) , .A( u2_u0_u6_n174 ) );
  NOR3_X1 u2_u0_u6_U83 (.A1( u2_u0_u6_n141 ) , .ZN( u2_u0_u6_n154 ) , .A3( u2_u0_u6_n164 ) , .A2( u2_u0_u6_n171 ) );
  AOI211_X1 u2_u0_u6_U84 (.B( u2_u0_u6_n149 ) , .A( u2_u0_u6_n150 ) , .C2( u2_u0_u6_n151 ) , .C1( u2_u0_u6_n152 ) , .ZN( u2_u0_u6_n153 ) );
  OAI211_X1 u2_u0_u6_U85 (.ZN( u2_out0_22 ) , .B( u2_u0_u6_n137 ) , .A( u2_u0_u6_n138 ) , .C2( u2_u0_u6_n139 ) , .C1( u2_u0_u6_n140 ) );
  AOI22_X1 u2_u0_u6_U86 (.B1( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n138 ) , .B2( u2_u0_u6_n161 ) );
  AND4_X1 u2_u0_u6_U87 (.A3( u2_u0_u6_n119 ) , .A1( u2_u0_u6_n120 ) , .A4( u2_u0_u6_n129 ) , .ZN( u2_u0_u6_n140 ) , .A2( u2_u0_u6_n143 ) );
  NAND3_X1 u2_u0_u6_U88 (.A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n130 ) , .A3( u2_u0_u6_n131 ) );
  NAND3_X1 u2_u0_u6_U89 (.A3( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n141 ) , .A1( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U9 (.ZN( u2_u0_u6_n172 ) , .A( u2_u0_u6_n88 ) );
  NAND3_X1 u2_u0_u6_U90 (.ZN( u2_u0_u6_n101 ) , .A3( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n127 ) );
  NAND3_X1 u2_u0_u6_U91 (.ZN( u2_u0_u6_n102 ) , .A3( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n145 ) , .A1( u2_u0_u6_n166 ) );
  NAND3_X1 u2_u0_u6_U92 (.A3( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n93 ) );
  NAND3_X1 u2_u0_u6_U93 (.ZN( u2_u0_u6_n142 ) , .A2( u2_u0_u6_n172 ) , .A3( u2_u0_u6_n89 ) , .A1( u2_u0_u6_n90 ) );
  INV_X1 u2_u0_u7_U10 (.A( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n176 ) );
  OAI221_X1 u2_u0_u7_U11 (.C1( u2_u0_u7_n101 ) , .C2( u2_u0_u7_n147 ) , .ZN( u2_u0_u7_n155 ) , .B2( u2_u0_u7_n162 ) , .A( u2_u0_u7_n91 ) , .B1( u2_u0_u7_n92 ) );
  AND3_X1 u2_u0_u7_U12 (.A3( u2_u0_u7_n110 ) , .A2( u2_u0_u7_n127 ) , .A1( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n92 ) );
  OAI21_X1 u2_u0_u7_U13 (.A( u2_u0_u7_n161 ) , .B1( u2_u0_u7_n168 ) , .B2( u2_u0_u7_n173 ) , .ZN( u2_u0_u7_n91 ) );
  AOI211_X1 u2_u0_u7_U14 (.A( u2_u0_u7_n117 ) , .ZN( u2_u0_u7_n118 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n177 ) , .B( u2_u0_u7_n180 ) );
  OAI22_X1 u2_u0_u7_U15 (.B1( u2_u0_u7_n115 ) , .ZN( u2_u0_u7_n117 ) , .A2( u2_u0_u7_n133 ) , .A1( u2_u0_u7_n137 ) , .B2( u2_u0_u7_n162 ) );
  INV_X1 u2_u0_u7_U16 (.A( u2_u0_u7_n116 ) , .ZN( u2_u0_u7_n180 ) );
  NOR3_X1 u2_u0_u7_U17 (.ZN( u2_u0_u7_n115 ) , .A3( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n168 ) , .A1( u2_u0_u7_n169 ) );
  NOR3_X1 u2_u0_u7_U18 (.A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n135 ) , .ZN( u2_u0_u7_n136 ) , .A3( u2_u0_u7_n171 ) );
  NOR2_X1 u2_u0_u7_U19 (.A1( u2_u0_u7_n130 ) , .A2( u2_u0_u7_n134 ) , .ZN( u2_u0_u7_n153 ) );
  INV_X1 u2_u0_u7_U20 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n165 ) );
  NOR2_X1 u2_u0_u7_U21 (.ZN( u2_u0_u7_n111 ) , .A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n169 ) );
  AOI21_X1 u2_u0_u7_U22 (.ZN( u2_u0_u7_n104 ) , .B2( u2_u0_u7_n112 ) , .B1( u2_u0_u7_n127 ) , .A( u2_u0_u7_n164 ) );
  AOI21_X1 u2_u0_u7_U23 (.ZN( u2_u0_u7_n106 ) , .B1( u2_u0_u7_n133 ) , .B2( u2_u0_u7_n146 ) , .A( u2_u0_u7_n162 ) );
  AOI21_X1 u2_u0_u7_U24 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n107 ) , .B2( u2_u0_u7_n128 ) , .B1( u2_u0_u7_n175 ) );
  INV_X1 u2_u0_u7_U25 (.A( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n171 ) );
  INV_X1 u2_u0_u7_U26 (.A( u2_u0_u7_n131 ) , .ZN( u2_u0_u7_n177 ) );
  INV_X1 u2_u0_u7_U27 (.A( u2_u0_u7_n110 ) , .ZN( u2_u0_u7_n174 ) );
  NAND2_X1 u2_u0_u7_U28 (.A1( u2_u0_u7_n129 ) , .A2( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n149 ) );
  NAND2_X1 u2_u0_u7_U29 (.A1( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n130 ) );
  OAI21_X1 u2_u0_u7_U3 (.ZN( u2_u0_u7_n159 ) , .A( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n171 ) , .B1( u2_u0_u7_n174 ) );
  INV_X1 u2_u0_u7_U30 (.A( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n173 ) );
  INV_X1 u2_u0_u7_U31 (.A( u2_u0_u7_n128 ) , .ZN( u2_u0_u7_n168 ) );
  INV_X1 u2_u0_u7_U32 (.A( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n169 ) );
  INV_X1 u2_u0_u7_U33 (.A( u2_u0_u7_n127 ) , .ZN( u2_u0_u7_n179 ) );
  NOR2_X1 u2_u0_u7_U34 (.ZN( u2_u0_u7_n101 ) , .A2( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n156 ) );
  AOI211_X1 u2_u0_u7_U35 (.B( u2_u0_u7_n139 ) , .A( u2_u0_u7_n140 ) , .C2( u2_u0_u7_n141 ) , .ZN( u2_u0_u7_n142 ) , .C1( u2_u0_u7_n156 ) );
  NAND4_X1 u2_u0_u7_U36 (.A3( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n141 ) , .A4( u2_u0_u7_n147 ) );
  AOI21_X1 u2_u0_u7_U37 (.A( u2_u0_u7_n137 ) , .B1( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n139 ) , .B2( u2_u0_u7_n146 ) );
  OAI22_X1 u2_u0_u7_U38 (.B1( u2_u0_u7_n136 ) , .ZN( u2_u0_u7_n140 ) , .A1( u2_u0_u7_n153 ) , .B2( u2_u0_u7_n162 ) , .A2( u2_u0_u7_n164 ) );
  AOI211_X1 u2_u0_u7_U39 (.B( u2_u0_u7_n154 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n156 ) , .ZN( u2_u0_u7_n157 ) , .C2( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U4 (.A( u2_u0_u7_n111 ) , .ZN( u2_u0_u7_n170 ) );
  INV_X1 u2_u0_u7_U40 (.A( u2_u0_u7_n153 ) , .ZN( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U41 (.A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n161 ) );
  NAND2_X1 u2_u0_u7_U42 (.A2( u2_u0_u7_n102 ) , .A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n133 ) );
  NAND2_X1 u2_u0_u7_U43 (.A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n99 ) );
  AOI21_X1 u2_u0_u7_U44 (.ZN( u2_u0_u7_n123 ) , .B1( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n177 ) , .A( u2_u0_u7_n97 ) );
  AOI21_X1 u2_u0_u7_U45 (.B2( u2_u0_u7_n113 ) , .B1( u2_u0_u7_n124 ) , .A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n97 ) );
  INV_X1 u2_u0_u7_U46 (.A( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n162 ) );
  AND2_X1 u2_u0_u7_U47 (.ZN( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n98 ) , .A1( u2_u0_u7_n99 ) );
  NOR2_X1 u2_u0_u7_U48 (.ZN( u2_u0_u7_n137 ) , .A1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n161 ) );
  AOI21_X1 u2_u0_u7_U49 (.ZN( u2_u0_u7_n105 ) , .B2( u2_u0_u7_n110 ) , .A( u2_u0_u7_n125 ) , .B1( u2_u0_u7_n147 ) );
  INV_X1 u2_u0_u7_U5 (.A( u2_u0_u7_n154 ) , .ZN( u2_u0_u7_n178 ) );
  NAND2_X1 u2_u0_u7_U50 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U51 (.ZN( u2_u0_u7_n146 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n98 ) );
  OR2_X1 u2_u0_u7_U52 (.ZN( u2_u0_u7_n126 ) , .A2( u2_u0_u7_n152 ) , .A1( u2_u0_u7_n156 ) );
  NAND2_X1 u2_u0_u7_U53 (.ZN( u2_u0_u7_n112 ) , .A2( u2_u0_u7_n96 ) , .A1( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U54 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U55 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U56 (.ZN( u2_u0_u7_n110 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n96 ) );
  INV_X1 u2_u0_u7_U57 (.A( u2_u0_u7_n150 ) , .ZN( u2_u0_u7_n164 ) );
  AND2_X1 u2_u0_u7_U58 (.ZN( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U59 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n131 ) , .A1( u2_u0_u7_n95 ) );
  INV_X1 u2_u0_u7_U6 (.A( u2_u0_u7_n149 ) , .ZN( u2_u0_u7_n175 ) );
  NAND2_X1 u2_u0_u7_U60 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n124 ) , .A1( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U61 (.A1( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n129 ) );
  NAND2_X1 u2_u0_u7_U62 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n138 ) , .A2( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U63 (.ZN( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U64 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n148 ) , .A2( u2_u0_u7_n95 ) );
  AOI22_X1 u2_u0_u7_U65 (.A2( u2_u0_u7_n114 ) , .ZN( u2_u0_u7_n119 ) , .B1( u2_u0_u7_n130 ) , .A1( u2_u0_u7_n156 ) , .B2( u2_u0_u7_n165 ) );
  NAND2_X1 u2_u0_u7_U66 (.A2( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n114 ) , .A1( u2_u0_u7_n175 ) );
  NOR2_X1 u2_u0_u7_U67 (.A2( u2_u0_X_47 ) , .ZN( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n163 ) );
  NOR2_X1 u2_u0_u7_U68 (.A2( u2_u0_X_48 ) , .A1( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n95 ) );
  NOR2_X1 u2_u0_u7_U69 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n99 ) );
  AOI211_X1 u2_u0_u7_U7 (.ZN( u2_u0_u7_n116 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n161 ) , .C2( u2_u0_u7_n171 ) , .B( u2_u0_u7_n94 ) );
  NOR2_X1 u2_u0_u7_U70 (.A2( u2_u0_X_44 ) , .A1( u2_u0_u7_n167 ) , .ZN( u2_u0_u7_n98 ) );
  NOR2_X1 u2_u0_u7_U71 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n152 ) );
  AND2_X1 u2_u0_u7_U72 (.A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n156 ) , .A2( u2_u0_u7_n163 ) );
  NAND2_X1 u2_u0_u7_U73 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n125 ) );
  AND2_X1 u2_u0_u7_U74 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n102 ) );
  AND2_X1 u2_u0_u7_U75 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n96 ) );
  AND2_X1 u2_u0_u7_U76 (.A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n167 ) );
  AND2_X1 u2_u0_u7_U77 (.A1( u2_u0_X_48 ) , .A2( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n93 ) );
  INV_X1 u2_u0_u7_U78 (.A( u2_u0_X_46 ) , .ZN( u2_u0_u7_n163 ) );
  INV_X1 u2_u0_u7_U79 (.A( u2_u0_X_45 ) , .ZN( u2_u0_u7_n166 ) );
  OAI222_X1 u2_u0_u7_U8 (.C2( u2_u0_u7_n101 ) , .B2( u2_u0_u7_n111 ) , .A1( u2_u0_u7_n113 ) , .C1( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n162 ) , .B1( u2_u0_u7_n164 ) , .ZN( u2_u0_u7_n94 ) );
  OAI21_X1 u2_u0_u7_U80 (.B1( u2_u0_u7_n145 ) , .ZN( u2_u0_u7_n160 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n177 ) );
  AOI22_X1 u2_u0_u7_U81 (.B2( u2_u0_u7_n149 ) , .B1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n151 ) , .A1( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n158 ) );
  NAND4_X1 u2_u0_u7_U82 (.ZN( u2_out0_27 ) , .A4( u2_u0_u7_n118 ) , .A3( u2_u0_u7_n119 ) , .A2( u2_u0_u7_n120 ) , .A1( u2_u0_u7_n121 ) );
  OAI21_X1 u2_u0_u7_U83 (.ZN( u2_u0_u7_n121 ) , .B2( u2_u0_u7_n145 ) , .A( u2_u0_u7_n150 ) , .B1( u2_u0_u7_n174 ) );
  OAI21_X1 u2_u0_u7_U84 (.ZN( u2_u0_u7_n120 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n170 ) , .B1( u2_u0_u7_n179 ) );
  NAND4_X1 u2_u0_u7_U85 (.ZN( u2_out0_15 ) , .A4( u2_u0_u7_n142 ) , .A3( u2_u0_u7_n143 ) , .A2( u2_u0_u7_n144 ) , .A1( u2_u0_u7_n178 ) );
  OR2_X1 u2_u0_u7_U86 (.A2( u2_u0_u7_n125 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n144 ) );
  AOI22_X1 u2_u0_u7_U87 (.A2( u2_u0_u7_n126 ) , .ZN( u2_u0_u7_n143 ) , .B2( u2_u0_u7_n165 ) , .B1( u2_u0_u7_n173 ) , .A1( u2_u0_u7_n174 ) );
  NAND4_X1 u2_u0_u7_U88 (.ZN( u2_out0_5 ) , .A4( u2_u0_u7_n108 ) , .A3( u2_u0_u7_n109 ) , .A1( u2_u0_u7_n116 ) , .A2( u2_u0_u7_n123 ) );
  AOI22_X1 u2_u0_u7_U89 (.ZN( u2_u0_u7_n109 ) , .A2( u2_u0_u7_n126 ) , .B2( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n156 ) , .A1( u2_u0_u7_n171 ) );
  AOI222_X1 u2_u0_u7_U9 (.ZN( u2_u0_u7_n122 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n161 ) , .A2( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n170 ) , .A1( u2_u0_u7_n176 ) );
  NOR4_X1 u2_u0_u7_U90 (.A4( u2_u0_u7_n104 ) , .A3( u2_u0_u7_n105 ) , .A2( u2_u0_u7_n106 ) , .A1( u2_u0_u7_n107 ) , .ZN( u2_u0_u7_n108 ) );
  NAND4_X1 u2_u0_u7_U91 (.ZN( u2_out0_21 ) , .A4( u2_u0_u7_n157 ) , .A3( u2_u0_u7_n158 ) , .A2( u2_u0_u7_n159 ) , .A1( u2_u0_u7_n160 ) );
  OAI211_X1 u2_u0_u7_U92 (.B( u2_u0_u7_n122 ) , .A( u2_u0_u7_n123 ) , .C2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n154 ) , .C1( u2_u0_u7_n162 ) );
  NOR2_X1 u2_u0_u7_U93 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n103 ) );
  INV_X1 u2_u0_u7_U94 (.A( u2_u0_X_43 ) , .ZN( u2_u0_u7_n167 ) );
  NAND3_X1 u2_u0_u7_U95 (.A3( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n151 ) );
  NAND3_X1 u2_u0_u7_U96 (.A3( u2_u0_u7_n131 ) , .A2( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n135 ) );
  XOR2_X1 u2_u10_U10 (.B( u2_K11_45 ) , .A( u2_R9_30 ) , .Z( u2_u10_X_45 ) );
  XOR2_X1 u2_u10_U11 (.B( u2_K11_44 ) , .A( u2_R9_29 ) , .Z( u2_u10_X_44 ) );
  XOR2_X1 u2_u10_U12 (.B( u2_K11_43 ) , .A( u2_R9_28 ) , .Z( u2_u10_X_43 ) );
  XOR2_X1 u2_u10_U13 (.B( u2_K11_42 ) , .A( u2_R9_29 ) , .Z( u2_u10_X_42 ) );
  XOR2_X1 u2_u10_U14 (.B( u2_K11_41 ) , .A( u2_R9_28 ) , .Z( u2_u10_X_41 ) );
  XOR2_X1 u2_u10_U15 (.B( u2_K11_40 ) , .A( u2_R9_27 ) , .Z( u2_u10_X_40 ) );
  XOR2_X1 u2_u10_U17 (.B( u2_K11_39 ) , .A( u2_R9_26 ) , .Z( u2_u10_X_39 ) );
  XOR2_X1 u2_u10_U18 (.B( u2_K11_38 ) , .A( u2_R9_25 ) , .Z( u2_u10_X_38 ) );
  XOR2_X1 u2_u10_U19 (.B( u2_K11_37 ) , .A( u2_R9_24 ) , .Z( u2_u10_X_37 ) );
  XOR2_X1 u2_u10_U20 (.B( u2_K11_36 ) , .A( u2_R9_25 ) , .Z( u2_u10_X_36 ) );
  XOR2_X1 u2_u10_U21 (.B( u2_K11_35 ) , .A( u2_R9_24 ) , .Z( u2_u10_X_35 ) );
  XOR2_X1 u2_u10_U22 (.B( u2_K11_34 ) , .A( u2_R9_23 ) , .Z( u2_u10_X_34 ) );
  XOR2_X1 u2_u10_U23 (.B( u2_K11_33 ) , .A( u2_R9_22 ) , .Z( u2_u10_X_33 ) );
  XOR2_X1 u2_u10_U24 (.B( u2_K11_32 ) , .A( u2_R9_21 ) , .Z( u2_u10_X_32 ) );
  XOR2_X1 u2_u10_U25 (.B( u2_K11_31 ) , .A( u2_R9_20 ) , .Z( u2_u10_X_31 ) );
  XOR2_X1 u2_u10_U40 (.B( u2_K11_18 ) , .A( u2_R9_13 ) , .Z( u2_u10_X_18 ) );
  XOR2_X1 u2_u10_U41 (.B( u2_K11_17 ) , .A( u2_R9_12 ) , .Z( u2_u10_X_17 ) );
  XOR2_X1 u2_u10_U42 (.B( u2_K11_16 ) , .A( u2_R9_11 ) , .Z( u2_u10_X_16 ) );
  XOR2_X1 u2_u10_U43 (.B( u2_K11_15 ) , .A( u2_R9_10 ) , .Z( u2_u10_X_15 ) );
  XOR2_X1 u2_u10_U44 (.B( u2_K11_14 ) , .A( u2_R9_9 ) , .Z( u2_u10_X_14 ) );
  XOR2_X1 u2_u10_U45 (.B( u2_K11_13 ) , .A( u2_R9_8 ) , .Z( u2_u10_X_13 ) );
  XOR2_X1 u2_u10_U7 (.B( u2_K11_48 ) , .A( u2_R9_1 ) , .Z( u2_u10_X_48 ) );
  XOR2_X1 u2_u10_U8 (.B( u2_K11_47 ) , .A( u2_R9_32 ) , .Z( u2_u10_X_47 ) );
  XOR2_X1 u2_u10_U9 (.B( u2_K11_46 ) , .A( u2_R9_31 ) , .Z( u2_u10_X_46 ) );
  OAI22_X1 u2_u10_u2_U10 (.ZN( u2_u10_u2_n109 ) , .A2( u2_u10_u2_n113 ) , .B2( u2_u10_u2_n133 ) , .B1( u2_u10_u2_n167 ) , .A1( u2_u10_u2_n168 ) );
  NAND3_X1 u2_u10_u2_U100 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n98 ) );
  OAI22_X1 u2_u10_u2_U11 (.B1( u2_u10_u2_n151 ) , .A2( u2_u10_u2_n152 ) , .A1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n160 ) , .B2( u2_u10_u2_n168 ) );
  NOR3_X1 u2_u10_u2_U12 (.A1( u2_u10_u2_n150 ) , .ZN( u2_u10_u2_n151 ) , .A3( u2_u10_u2_n175 ) , .A2( u2_u10_u2_n188 ) );
  AOI21_X1 u2_u10_u2_U13 (.ZN( u2_u10_u2_n144 ) , .B2( u2_u10_u2_n155 ) , .A( u2_u10_u2_n172 ) , .B1( u2_u10_u2_n185 ) );
  AOI21_X1 u2_u10_u2_U14 (.B2( u2_u10_u2_n143 ) , .ZN( u2_u10_u2_n145 ) , .B1( u2_u10_u2_n152 ) , .A( u2_u10_u2_n171 ) );
  AOI21_X1 u2_u10_u2_U15 (.B2( u2_u10_u2_n120 ) , .B1( u2_u10_u2_n121 ) , .ZN( u2_u10_u2_n126 ) , .A( u2_u10_u2_n167 ) );
  INV_X1 u2_u10_u2_U16 (.A( u2_u10_u2_n156 ) , .ZN( u2_u10_u2_n171 ) );
  INV_X1 u2_u10_u2_U17 (.A( u2_u10_u2_n120 ) , .ZN( u2_u10_u2_n188 ) );
  NAND2_X1 u2_u10_u2_U18 (.A2( u2_u10_u2_n122 ) , .ZN( u2_u10_u2_n150 ) , .A1( u2_u10_u2_n152 ) );
  INV_X1 u2_u10_u2_U19 (.A( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n170 ) );
  INV_X1 u2_u10_u2_U20 (.A( u2_u10_u2_n137 ) , .ZN( u2_u10_u2_n173 ) );
  NAND2_X1 u2_u10_u2_U21 (.A1( u2_u10_u2_n132 ) , .A2( u2_u10_u2_n139 ) , .ZN( u2_u10_u2_n157 ) );
  INV_X1 u2_u10_u2_U22 (.A( u2_u10_u2_n113 ) , .ZN( u2_u10_u2_n178 ) );
  INV_X1 u2_u10_u2_U23 (.A( u2_u10_u2_n139 ) , .ZN( u2_u10_u2_n175 ) );
  INV_X1 u2_u10_u2_U24 (.A( u2_u10_u2_n155 ) , .ZN( u2_u10_u2_n181 ) );
  INV_X1 u2_u10_u2_U25 (.A( u2_u10_u2_n119 ) , .ZN( u2_u10_u2_n177 ) );
  INV_X1 u2_u10_u2_U26 (.A( u2_u10_u2_n116 ) , .ZN( u2_u10_u2_n180 ) );
  INV_X1 u2_u10_u2_U27 (.A( u2_u10_u2_n131 ) , .ZN( u2_u10_u2_n179 ) );
  INV_X1 u2_u10_u2_U28 (.A( u2_u10_u2_n154 ) , .ZN( u2_u10_u2_n176 ) );
  NAND2_X1 u2_u10_u2_U29 (.A2( u2_u10_u2_n116 ) , .A1( u2_u10_u2_n117 ) , .ZN( u2_u10_u2_n118 ) );
  NOR2_X1 u2_u10_u2_U3 (.ZN( u2_u10_u2_n121 ) , .A2( u2_u10_u2_n177 ) , .A1( u2_u10_u2_n180 ) );
  INV_X1 u2_u10_u2_U30 (.A( u2_u10_u2_n132 ) , .ZN( u2_u10_u2_n182 ) );
  INV_X1 u2_u10_u2_U31 (.A( u2_u10_u2_n158 ) , .ZN( u2_u10_u2_n183 ) );
  OAI21_X1 u2_u10_u2_U32 (.A( u2_u10_u2_n156 ) , .B1( u2_u10_u2_n157 ) , .ZN( u2_u10_u2_n158 ) , .B2( u2_u10_u2_n179 ) );
  NOR2_X1 u2_u10_u2_U33 (.ZN( u2_u10_u2_n156 ) , .A1( u2_u10_u2_n166 ) , .A2( u2_u10_u2_n169 ) );
  NOR2_X1 u2_u10_u2_U34 (.A2( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n137 ) , .A1( u2_u10_u2_n140 ) );
  NOR2_X1 u2_u10_u2_U35 (.A2( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n153 ) , .A1( u2_u10_u2_n156 ) );
  AOI211_X1 u2_u10_u2_U36 (.ZN( u2_u10_u2_n130 ) , .C1( u2_u10_u2_n138 ) , .C2( u2_u10_u2_n179 ) , .B( u2_u10_u2_n96 ) , .A( u2_u10_u2_n97 ) );
  OAI22_X1 u2_u10_u2_U37 (.B1( u2_u10_u2_n133 ) , .A2( u2_u10_u2_n137 ) , .A1( u2_u10_u2_n152 ) , .B2( u2_u10_u2_n168 ) , .ZN( u2_u10_u2_n97 ) );
  OAI221_X1 u2_u10_u2_U38 (.B1( u2_u10_u2_n113 ) , .C1( u2_u10_u2_n132 ) , .A( u2_u10_u2_n149 ) , .B2( u2_u10_u2_n171 ) , .C2( u2_u10_u2_n172 ) , .ZN( u2_u10_u2_n96 ) );
  OAI221_X1 u2_u10_u2_U39 (.A( u2_u10_u2_n115 ) , .C2( u2_u10_u2_n123 ) , .B2( u2_u10_u2_n143 ) , .B1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n163 ) , .C1( u2_u10_u2_n168 ) );
  INV_X1 u2_u10_u2_U4 (.A( u2_u10_u2_n134 ) , .ZN( u2_u10_u2_n185 ) );
  OAI21_X1 u2_u10_u2_U40 (.A( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n115 ) , .B1( u2_u10_u2_n176 ) , .B2( u2_u10_u2_n178 ) );
  OAI221_X1 u2_u10_u2_U41 (.A( u2_u10_u2_n135 ) , .B2( u2_u10_u2_n136 ) , .B1( u2_u10_u2_n137 ) , .ZN( u2_u10_u2_n162 ) , .C2( u2_u10_u2_n167 ) , .C1( u2_u10_u2_n185 ) );
  AND3_X1 u2_u10_u2_U42 (.A3( u2_u10_u2_n131 ) , .A2( u2_u10_u2_n132 ) , .A1( u2_u10_u2_n133 ) , .ZN( u2_u10_u2_n136 ) );
  AOI22_X1 u2_u10_u2_U43 (.ZN( u2_u10_u2_n135 ) , .B1( u2_u10_u2_n140 ) , .A1( u2_u10_u2_n156 ) , .B2( u2_u10_u2_n180 ) , .A2( u2_u10_u2_n188 ) );
  AOI21_X1 u2_u10_u2_U44 (.ZN( u2_u10_u2_n149 ) , .B1( u2_u10_u2_n173 ) , .B2( u2_u10_u2_n188 ) , .A( u2_u10_u2_n95 ) );
  AND3_X1 u2_u10_u2_U45 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n156 ) , .ZN( u2_u10_u2_n95 ) );
  OAI21_X1 u2_u10_u2_U46 (.A( u2_u10_u2_n141 ) , .B2( u2_u10_u2_n142 ) , .ZN( u2_u10_u2_n146 ) , .B1( u2_u10_u2_n153 ) );
  OAI21_X1 u2_u10_u2_U47 (.A( u2_u10_u2_n140 ) , .ZN( u2_u10_u2_n141 ) , .B1( u2_u10_u2_n176 ) , .B2( u2_u10_u2_n177 ) );
  NOR3_X1 u2_u10_u2_U48 (.ZN( u2_u10_u2_n142 ) , .A3( u2_u10_u2_n175 ) , .A2( u2_u10_u2_n178 ) , .A1( u2_u10_u2_n181 ) );
  OAI21_X1 u2_u10_u2_U49 (.A( u2_u10_u2_n101 ) , .B2( u2_u10_u2_n121 ) , .B1( u2_u10_u2_n153 ) , .ZN( u2_u10_u2_n164 ) );
  INV_X1 u2_u10_u2_U5 (.A( u2_u10_u2_n150 ) , .ZN( u2_u10_u2_n184 ) );
  NAND2_X1 u2_u10_u2_U50 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n155 ) );
  NAND2_X1 u2_u10_u2_U51 (.A2( u2_u10_u2_n105 ) , .A1( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n143 ) );
  NAND2_X1 u2_u10_u2_U52 (.A1( u2_u10_u2_n104 ) , .A2( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n152 ) );
  NAND2_X1 u2_u10_u2_U53 (.A1( u2_u10_u2_n100 ) , .A2( u2_u10_u2_n105 ) , .ZN( u2_u10_u2_n132 ) );
  INV_X1 u2_u10_u2_U54 (.A( u2_u10_u2_n140 ) , .ZN( u2_u10_u2_n168 ) );
  INV_X1 u2_u10_u2_U55 (.A( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n167 ) );
  NAND2_X1 u2_u10_u2_U56 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n113 ) );
  NAND2_X1 u2_u10_u2_U57 (.A1( u2_u10_u2_n106 ) , .A2( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n131 ) );
  NAND2_X1 u2_u10_u2_U58 (.A1( u2_u10_u2_n103 ) , .A2( u2_u10_u2_n107 ) , .ZN( u2_u10_u2_n139 ) );
  NAND2_X1 u2_u10_u2_U59 (.A1( u2_u10_u2_n103 ) , .A2( u2_u10_u2_n105 ) , .ZN( u2_u10_u2_n133 ) );
  NOR4_X1 u2_u10_u2_U6 (.A4( u2_u10_u2_n124 ) , .A3( u2_u10_u2_n125 ) , .A2( u2_u10_u2_n126 ) , .A1( u2_u10_u2_n127 ) , .ZN( u2_u10_u2_n128 ) );
  NAND2_X1 u2_u10_u2_U60 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n103 ) , .ZN( u2_u10_u2_n154 ) );
  NAND2_X1 u2_u10_u2_U61 (.A2( u2_u10_u2_n103 ) , .A1( u2_u10_u2_n104 ) , .ZN( u2_u10_u2_n119 ) );
  NAND2_X1 u2_u10_u2_U62 (.A2( u2_u10_u2_n107 ) , .A1( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n123 ) );
  NAND2_X1 u2_u10_u2_U63 (.A1( u2_u10_u2_n104 ) , .A2( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n122 ) );
  INV_X1 u2_u10_u2_U64 (.A( u2_u10_u2_n114 ) , .ZN( u2_u10_u2_n172 ) );
  NAND2_X1 u2_u10_u2_U65 (.A2( u2_u10_u2_n100 ) , .A1( u2_u10_u2_n102 ) , .ZN( u2_u10_u2_n116 ) );
  NAND2_X1 u2_u10_u2_U66 (.A1( u2_u10_u2_n102 ) , .A2( u2_u10_u2_n108 ) , .ZN( u2_u10_u2_n120 ) );
  NAND2_X1 u2_u10_u2_U67 (.A2( u2_u10_u2_n105 ) , .A1( u2_u10_u2_n106 ) , .ZN( u2_u10_u2_n117 ) );
  INV_X1 u2_u10_u2_U68 (.ZN( u2_u10_u2_n187 ) , .A( u2_u10_u2_n99 ) );
  OAI21_X1 u2_u10_u2_U69 (.B1( u2_u10_u2_n137 ) , .B2( u2_u10_u2_n143 ) , .A( u2_u10_u2_n98 ) , .ZN( u2_u10_u2_n99 ) );
  AOI21_X1 u2_u10_u2_U7 (.ZN( u2_u10_u2_n124 ) , .B1( u2_u10_u2_n131 ) , .B2( u2_u10_u2_n143 ) , .A( u2_u10_u2_n172 ) );
  NOR2_X1 u2_u10_u2_U70 (.A2( u2_u10_X_16 ) , .ZN( u2_u10_u2_n140 ) , .A1( u2_u10_u2_n166 ) );
  NOR2_X1 u2_u10_u2_U71 (.A2( u2_u10_X_13 ) , .A1( u2_u10_X_14 ) , .ZN( u2_u10_u2_n100 ) );
  NOR2_X1 u2_u10_u2_U72 (.A2( u2_u10_X_16 ) , .A1( u2_u10_X_17 ) , .ZN( u2_u10_u2_n138 ) );
  NOR2_X1 u2_u10_u2_U73 (.A2( u2_u10_X_15 ) , .A1( u2_u10_X_18 ) , .ZN( u2_u10_u2_n104 ) );
  NOR2_X1 u2_u10_u2_U74 (.A2( u2_u10_X_14 ) , .ZN( u2_u10_u2_n103 ) , .A1( u2_u10_u2_n174 ) );
  NOR2_X1 u2_u10_u2_U75 (.A2( u2_u10_X_15 ) , .ZN( u2_u10_u2_n102 ) , .A1( u2_u10_u2_n165 ) );
  NOR2_X1 u2_u10_u2_U76 (.A2( u2_u10_X_17 ) , .ZN( u2_u10_u2_n114 ) , .A1( u2_u10_u2_n169 ) );
  AND2_X1 u2_u10_u2_U77 (.A1( u2_u10_X_15 ) , .ZN( u2_u10_u2_n105 ) , .A2( u2_u10_u2_n165 ) );
  AND2_X1 u2_u10_u2_U78 (.A2( u2_u10_X_15 ) , .A1( u2_u10_X_18 ) , .ZN( u2_u10_u2_n107 ) );
  AND2_X1 u2_u10_u2_U79 (.A1( u2_u10_X_14 ) , .ZN( u2_u10_u2_n106 ) , .A2( u2_u10_u2_n174 ) );
  AOI21_X1 u2_u10_u2_U8 (.B2( u2_u10_u2_n119 ) , .ZN( u2_u10_u2_n127 ) , .A( u2_u10_u2_n137 ) , .B1( u2_u10_u2_n155 ) );
  AND2_X1 u2_u10_u2_U80 (.A1( u2_u10_X_13 ) , .A2( u2_u10_X_14 ) , .ZN( u2_u10_u2_n108 ) );
  INV_X1 u2_u10_u2_U81 (.A( u2_u10_X_16 ) , .ZN( u2_u10_u2_n169 ) );
  INV_X1 u2_u10_u2_U82 (.A( u2_u10_X_17 ) , .ZN( u2_u10_u2_n166 ) );
  INV_X1 u2_u10_u2_U83 (.A( u2_u10_X_13 ) , .ZN( u2_u10_u2_n174 ) );
  INV_X1 u2_u10_u2_U84 (.A( u2_u10_X_18 ) , .ZN( u2_u10_u2_n165 ) );
  NAND4_X1 u2_u10_u2_U85 (.ZN( u2_out10_24 ) , .A4( u2_u10_u2_n111 ) , .A3( u2_u10_u2_n112 ) , .A1( u2_u10_u2_n130 ) , .A2( u2_u10_u2_n187 ) );
  AOI221_X1 u2_u10_u2_U86 (.A( u2_u10_u2_n109 ) , .B1( u2_u10_u2_n110 ) , .ZN( u2_u10_u2_n111 ) , .C1( u2_u10_u2_n134 ) , .C2( u2_u10_u2_n170 ) , .B2( u2_u10_u2_n173 ) );
  AOI21_X1 u2_u10_u2_U87 (.ZN( u2_u10_u2_n112 ) , .B2( u2_u10_u2_n156 ) , .A( u2_u10_u2_n164 ) , .B1( u2_u10_u2_n181 ) );
  NAND4_X1 u2_u10_u2_U88 (.ZN( u2_out10_16 ) , .A4( u2_u10_u2_n128 ) , .A3( u2_u10_u2_n129 ) , .A1( u2_u10_u2_n130 ) , .A2( u2_u10_u2_n186 ) );
  AOI22_X1 u2_u10_u2_U89 (.A2( u2_u10_u2_n118 ) , .ZN( u2_u10_u2_n129 ) , .A1( u2_u10_u2_n140 ) , .B1( u2_u10_u2_n157 ) , .B2( u2_u10_u2_n170 ) );
  AOI21_X1 u2_u10_u2_U9 (.B2( u2_u10_u2_n123 ) , .ZN( u2_u10_u2_n125 ) , .A( u2_u10_u2_n171 ) , .B1( u2_u10_u2_n184 ) );
  INV_X1 u2_u10_u2_U90 (.A( u2_u10_u2_n163 ) , .ZN( u2_u10_u2_n186 ) );
  NAND4_X1 u2_u10_u2_U91 (.ZN( u2_out10_30 ) , .A4( u2_u10_u2_n147 ) , .A3( u2_u10_u2_n148 ) , .A2( u2_u10_u2_n149 ) , .A1( u2_u10_u2_n187 ) );
  NOR3_X1 u2_u10_u2_U92 (.A3( u2_u10_u2_n144 ) , .A2( u2_u10_u2_n145 ) , .A1( u2_u10_u2_n146 ) , .ZN( u2_u10_u2_n147 ) );
  AOI21_X1 u2_u10_u2_U93 (.B2( u2_u10_u2_n138 ) , .ZN( u2_u10_u2_n148 ) , .A( u2_u10_u2_n162 ) , .B1( u2_u10_u2_n182 ) );
  OR4_X1 u2_u10_u2_U94 (.ZN( u2_out10_6 ) , .A4( u2_u10_u2_n161 ) , .A3( u2_u10_u2_n162 ) , .A2( u2_u10_u2_n163 ) , .A1( u2_u10_u2_n164 ) );
  OR3_X1 u2_u10_u2_U95 (.A2( u2_u10_u2_n159 ) , .A1( u2_u10_u2_n160 ) , .ZN( u2_u10_u2_n161 ) , .A3( u2_u10_u2_n183 ) );
  AOI21_X1 u2_u10_u2_U96 (.B2( u2_u10_u2_n154 ) , .B1( u2_u10_u2_n155 ) , .ZN( u2_u10_u2_n159 ) , .A( u2_u10_u2_n167 ) );
  NAND3_X1 u2_u10_u2_U97 (.A2( u2_u10_u2_n117 ) , .A1( u2_u10_u2_n122 ) , .A3( u2_u10_u2_n123 ) , .ZN( u2_u10_u2_n134 ) );
  NAND3_X1 u2_u10_u2_U98 (.ZN( u2_u10_u2_n110 ) , .A2( u2_u10_u2_n131 ) , .A3( u2_u10_u2_n139 ) , .A1( u2_u10_u2_n154 ) );
  NAND3_X1 u2_u10_u2_U99 (.A2( u2_u10_u2_n100 ) , .ZN( u2_u10_u2_n101 ) , .A1( u2_u10_u2_n104 ) , .A3( u2_u10_u2_n114 ) );
  INV_X1 u2_u10_u5_U10 (.A( u2_u10_u5_n121 ) , .ZN( u2_u10_u5_n177 ) );
  NOR3_X1 u2_u10_u5_U100 (.A3( u2_u10_u5_n141 ) , .A1( u2_u10_u5_n142 ) , .ZN( u2_u10_u5_n143 ) , .A2( u2_u10_u5_n191 ) );
  NAND4_X1 u2_u10_u5_U101 (.ZN( u2_out10_4 ) , .A4( u2_u10_u5_n112 ) , .A2( u2_u10_u5_n113 ) , .A1( u2_u10_u5_n114 ) , .A3( u2_u10_u5_n195 ) );
  AOI211_X1 u2_u10_u5_U102 (.A( u2_u10_u5_n110 ) , .C1( u2_u10_u5_n111 ) , .ZN( u2_u10_u5_n112 ) , .B( u2_u10_u5_n118 ) , .C2( u2_u10_u5_n177 ) );
  AOI222_X1 u2_u10_u5_U103 (.ZN( u2_u10_u5_n113 ) , .A1( u2_u10_u5_n131 ) , .C1( u2_u10_u5_n148 ) , .B2( u2_u10_u5_n174 ) , .C2( u2_u10_u5_n178 ) , .A2( u2_u10_u5_n179 ) , .B1( u2_u10_u5_n99 ) );
  NAND3_X1 u2_u10_u5_U104 (.A2( u2_u10_u5_n154 ) , .A3( u2_u10_u5_n158 ) , .A1( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n99 ) );
  NOR2_X1 u2_u10_u5_U11 (.ZN( u2_u10_u5_n160 ) , .A2( u2_u10_u5_n173 ) , .A1( u2_u10_u5_n177 ) );
  INV_X1 u2_u10_u5_U12 (.A( u2_u10_u5_n150 ) , .ZN( u2_u10_u5_n174 ) );
  AOI21_X1 u2_u10_u5_U13 (.A( u2_u10_u5_n160 ) , .B2( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n162 ) , .B1( u2_u10_u5_n192 ) );
  INV_X1 u2_u10_u5_U14 (.A( u2_u10_u5_n159 ) , .ZN( u2_u10_u5_n192 ) );
  AOI21_X1 u2_u10_u5_U15 (.A( u2_u10_u5_n156 ) , .B2( u2_u10_u5_n157 ) , .B1( u2_u10_u5_n158 ) , .ZN( u2_u10_u5_n163 ) );
  AOI21_X1 u2_u10_u5_U16 (.B2( u2_u10_u5_n139 ) , .B1( u2_u10_u5_n140 ) , .ZN( u2_u10_u5_n141 ) , .A( u2_u10_u5_n150 ) );
  OAI21_X1 u2_u10_u5_U17 (.A( u2_u10_u5_n133 ) , .B2( u2_u10_u5_n134 ) , .B1( u2_u10_u5_n135 ) , .ZN( u2_u10_u5_n142 ) );
  OAI21_X1 u2_u10_u5_U18 (.ZN( u2_u10_u5_n133 ) , .B2( u2_u10_u5_n147 ) , .A( u2_u10_u5_n173 ) , .B1( u2_u10_u5_n188 ) );
  NAND2_X1 u2_u10_u5_U19 (.A2( u2_u10_u5_n119 ) , .A1( u2_u10_u5_n123 ) , .ZN( u2_u10_u5_n137 ) );
  INV_X1 u2_u10_u5_U20 (.A( u2_u10_u5_n155 ) , .ZN( u2_u10_u5_n194 ) );
  NAND2_X1 u2_u10_u5_U21 (.A1( u2_u10_u5_n121 ) , .ZN( u2_u10_u5_n132 ) , .A2( u2_u10_u5_n172 ) );
  NAND2_X1 u2_u10_u5_U22 (.A2( u2_u10_u5_n122 ) , .ZN( u2_u10_u5_n136 ) , .A1( u2_u10_u5_n154 ) );
  NAND2_X1 u2_u10_u5_U23 (.A2( u2_u10_u5_n119 ) , .A1( u2_u10_u5_n120 ) , .ZN( u2_u10_u5_n159 ) );
  INV_X1 u2_u10_u5_U24 (.A( u2_u10_u5_n156 ) , .ZN( u2_u10_u5_n175 ) );
  INV_X1 u2_u10_u5_U25 (.A( u2_u10_u5_n158 ) , .ZN( u2_u10_u5_n188 ) );
  INV_X1 u2_u10_u5_U26 (.A( u2_u10_u5_n152 ) , .ZN( u2_u10_u5_n179 ) );
  INV_X1 u2_u10_u5_U27 (.A( u2_u10_u5_n140 ) , .ZN( u2_u10_u5_n182 ) );
  INV_X1 u2_u10_u5_U28 (.A( u2_u10_u5_n151 ) , .ZN( u2_u10_u5_n183 ) );
  INV_X1 u2_u10_u5_U29 (.A( u2_u10_u5_n123 ) , .ZN( u2_u10_u5_n185 ) );
  NOR2_X1 u2_u10_u5_U3 (.ZN( u2_u10_u5_n134 ) , .A1( u2_u10_u5_n183 ) , .A2( u2_u10_u5_n190 ) );
  INV_X1 u2_u10_u5_U30 (.A( u2_u10_u5_n161 ) , .ZN( u2_u10_u5_n184 ) );
  INV_X1 u2_u10_u5_U31 (.A( u2_u10_u5_n139 ) , .ZN( u2_u10_u5_n189 ) );
  INV_X1 u2_u10_u5_U32 (.A( u2_u10_u5_n157 ) , .ZN( u2_u10_u5_n190 ) );
  INV_X1 u2_u10_u5_U33 (.A( u2_u10_u5_n120 ) , .ZN( u2_u10_u5_n193 ) );
  NAND2_X1 u2_u10_u5_U34 (.ZN( u2_u10_u5_n111 ) , .A1( u2_u10_u5_n140 ) , .A2( u2_u10_u5_n155 ) );
  NOR2_X1 u2_u10_u5_U35 (.ZN( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n170 ) , .A2( u2_u10_u5_n180 ) );
  INV_X1 u2_u10_u5_U36 (.A( u2_u10_u5_n117 ) , .ZN( u2_u10_u5_n196 ) );
  OAI221_X1 u2_u10_u5_U37 (.A( u2_u10_u5_n116 ) , .ZN( u2_u10_u5_n117 ) , .B2( u2_u10_u5_n119 ) , .C1( u2_u10_u5_n153 ) , .C2( u2_u10_u5_n158 ) , .B1( u2_u10_u5_n172 ) );
  AOI222_X1 u2_u10_u5_U38 (.ZN( u2_u10_u5_n116 ) , .B2( u2_u10_u5_n145 ) , .C1( u2_u10_u5_n148 ) , .A2( u2_u10_u5_n174 ) , .C2( u2_u10_u5_n177 ) , .B1( u2_u10_u5_n187 ) , .A1( u2_u10_u5_n193 ) );
  INV_X1 u2_u10_u5_U39 (.A( u2_u10_u5_n115 ) , .ZN( u2_u10_u5_n187 ) );
  INV_X1 u2_u10_u5_U4 (.A( u2_u10_u5_n138 ) , .ZN( u2_u10_u5_n191 ) );
  AOI22_X1 u2_u10_u5_U40 (.B2( u2_u10_u5_n131 ) , .A2( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n169 ) , .B1( u2_u10_u5_n174 ) , .A1( u2_u10_u5_n185 ) );
  NOR2_X1 u2_u10_u5_U41 (.A1( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n150 ) , .A2( u2_u10_u5_n173 ) );
  AOI21_X1 u2_u10_u5_U42 (.A( u2_u10_u5_n118 ) , .B2( u2_u10_u5_n145 ) , .ZN( u2_u10_u5_n168 ) , .B1( u2_u10_u5_n186 ) );
  INV_X1 u2_u10_u5_U43 (.A( u2_u10_u5_n122 ) , .ZN( u2_u10_u5_n186 ) );
  NOR2_X1 u2_u10_u5_U44 (.A1( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n152 ) , .A2( u2_u10_u5_n176 ) );
  NOR2_X1 u2_u10_u5_U45 (.A1( u2_u10_u5_n115 ) , .ZN( u2_u10_u5_n118 ) , .A2( u2_u10_u5_n153 ) );
  NOR2_X1 u2_u10_u5_U46 (.A2( u2_u10_u5_n145 ) , .ZN( u2_u10_u5_n156 ) , .A1( u2_u10_u5_n174 ) );
  NOR2_X1 u2_u10_u5_U47 (.ZN( u2_u10_u5_n121 ) , .A2( u2_u10_u5_n145 ) , .A1( u2_u10_u5_n176 ) );
  AOI22_X1 u2_u10_u5_U48 (.ZN( u2_u10_u5_n114 ) , .A2( u2_u10_u5_n137 ) , .A1( u2_u10_u5_n145 ) , .B2( u2_u10_u5_n175 ) , .B1( u2_u10_u5_n193 ) );
  OAI211_X1 u2_u10_u5_U49 (.B( u2_u10_u5_n124 ) , .A( u2_u10_u5_n125 ) , .C2( u2_u10_u5_n126 ) , .C1( u2_u10_u5_n127 ) , .ZN( u2_u10_u5_n128 ) );
  OAI21_X1 u2_u10_u5_U5 (.B2( u2_u10_u5_n136 ) , .B1( u2_u10_u5_n137 ) , .ZN( u2_u10_u5_n138 ) , .A( u2_u10_u5_n177 ) );
  NOR3_X1 u2_u10_u5_U50 (.ZN( u2_u10_u5_n127 ) , .A1( u2_u10_u5_n136 ) , .A3( u2_u10_u5_n148 ) , .A2( u2_u10_u5_n182 ) );
  OAI21_X1 u2_u10_u5_U51 (.ZN( u2_u10_u5_n124 ) , .A( u2_u10_u5_n177 ) , .B2( u2_u10_u5_n183 ) , .B1( u2_u10_u5_n189 ) );
  OAI21_X1 u2_u10_u5_U52 (.ZN( u2_u10_u5_n125 ) , .A( u2_u10_u5_n174 ) , .B2( u2_u10_u5_n185 ) , .B1( u2_u10_u5_n190 ) );
  AOI21_X1 u2_u10_u5_U53 (.A( u2_u10_u5_n153 ) , .B2( u2_u10_u5_n154 ) , .B1( u2_u10_u5_n155 ) , .ZN( u2_u10_u5_n164 ) );
  AOI21_X1 u2_u10_u5_U54 (.ZN( u2_u10_u5_n110 ) , .B1( u2_u10_u5_n122 ) , .B2( u2_u10_u5_n139 ) , .A( u2_u10_u5_n153 ) );
  INV_X1 u2_u10_u5_U55 (.A( u2_u10_u5_n153 ) , .ZN( u2_u10_u5_n176 ) );
  INV_X1 u2_u10_u5_U56 (.A( u2_u10_u5_n126 ) , .ZN( u2_u10_u5_n173 ) );
  AND2_X1 u2_u10_u5_U57 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n147 ) );
  AND2_X1 u2_u10_u5_U58 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n148 ) );
  NAND2_X1 u2_u10_u5_U59 (.A1( u2_u10_u5_n105 ) , .A2( u2_u10_u5_n106 ) , .ZN( u2_u10_u5_n158 ) );
  INV_X1 u2_u10_u5_U6 (.A( u2_u10_u5_n135 ) , .ZN( u2_u10_u5_n178 ) );
  NAND2_X1 u2_u10_u5_U60 (.A2( u2_u10_u5_n108 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n139 ) );
  NAND2_X1 u2_u10_u5_U61 (.A1( u2_u10_u5_n106 ) , .A2( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n119 ) );
  NAND2_X1 u2_u10_u5_U62 (.A2( u2_u10_u5_n103 ) , .A1( u2_u10_u5_n105 ) , .ZN( u2_u10_u5_n140 ) );
  NAND2_X1 u2_u10_u5_U63 (.A2( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n105 ) , .ZN( u2_u10_u5_n155 ) );
  NAND2_X1 u2_u10_u5_U64 (.A2( u2_u10_u5_n106 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n122 ) );
  NAND2_X1 u2_u10_u5_U65 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n106 ) , .ZN( u2_u10_u5_n115 ) );
  NAND2_X1 u2_u10_u5_U66 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n103 ) , .ZN( u2_u10_u5_n161 ) );
  NAND2_X1 u2_u10_u5_U67 (.A1( u2_u10_u5_n105 ) , .A2( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n154 ) );
  INV_X1 u2_u10_u5_U68 (.A( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n172 ) );
  NAND2_X1 u2_u10_u5_U69 (.A1( u2_u10_u5_n103 ) , .A2( u2_u10_u5_n108 ) , .ZN( u2_u10_u5_n123 ) );
  OAI22_X1 u2_u10_u5_U7 (.B2( u2_u10_u5_n149 ) , .B1( u2_u10_u5_n150 ) , .A2( u2_u10_u5_n151 ) , .A1( u2_u10_u5_n152 ) , .ZN( u2_u10_u5_n165 ) );
  NAND2_X1 u2_u10_u5_U70 (.A2( u2_u10_u5_n103 ) , .A1( u2_u10_u5_n107 ) , .ZN( u2_u10_u5_n151 ) );
  NAND2_X1 u2_u10_u5_U71 (.A2( u2_u10_u5_n107 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n120 ) );
  NAND2_X1 u2_u10_u5_U72 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n109 ) , .ZN( u2_u10_u5_n157 ) );
  AND2_X1 u2_u10_u5_U73 (.A2( u2_u10_u5_n100 ) , .A1( u2_u10_u5_n104 ) , .ZN( u2_u10_u5_n131 ) );
  INV_X1 u2_u10_u5_U74 (.A( u2_u10_u5_n102 ) , .ZN( u2_u10_u5_n195 ) );
  OAI221_X1 u2_u10_u5_U75 (.A( u2_u10_u5_n101 ) , .ZN( u2_u10_u5_n102 ) , .C2( u2_u10_u5_n115 ) , .C1( u2_u10_u5_n126 ) , .B1( u2_u10_u5_n134 ) , .B2( u2_u10_u5_n160 ) );
  OAI21_X1 u2_u10_u5_U76 (.ZN( u2_u10_u5_n101 ) , .B1( u2_u10_u5_n137 ) , .A( u2_u10_u5_n146 ) , .B2( u2_u10_u5_n147 ) );
  NOR2_X1 u2_u10_u5_U77 (.A2( u2_u10_X_34 ) , .A1( u2_u10_X_35 ) , .ZN( u2_u10_u5_n145 ) );
  NOR2_X1 u2_u10_u5_U78 (.A2( u2_u10_X_34 ) , .ZN( u2_u10_u5_n146 ) , .A1( u2_u10_u5_n171 ) );
  NOR2_X1 u2_u10_u5_U79 (.A2( u2_u10_X_31 ) , .A1( u2_u10_X_32 ) , .ZN( u2_u10_u5_n103 ) );
  NOR3_X1 u2_u10_u5_U8 (.A2( u2_u10_u5_n147 ) , .A1( u2_u10_u5_n148 ) , .ZN( u2_u10_u5_n149 ) , .A3( u2_u10_u5_n194 ) );
  NOR2_X1 u2_u10_u5_U80 (.A2( u2_u10_X_36 ) , .ZN( u2_u10_u5_n105 ) , .A1( u2_u10_u5_n180 ) );
  NOR2_X1 u2_u10_u5_U81 (.A2( u2_u10_X_33 ) , .ZN( u2_u10_u5_n108 ) , .A1( u2_u10_u5_n170 ) );
  NOR2_X1 u2_u10_u5_U82 (.A2( u2_u10_X_33 ) , .A1( u2_u10_X_36 ) , .ZN( u2_u10_u5_n107 ) );
  NOR2_X1 u2_u10_u5_U83 (.A2( u2_u10_X_31 ) , .ZN( u2_u10_u5_n104 ) , .A1( u2_u10_u5_n181 ) );
  NAND2_X1 u2_u10_u5_U84 (.A2( u2_u10_X_34 ) , .A1( u2_u10_X_35 ) , .ZN( u2_u10_u5_n153 ) );
  NAND2_X1 u2_u10_u5_U85 (.A1( u2_u10_X_34 ) , .ZN( u2_u10_u5_n126 ) , .A2( u2_u10_u5_n171 ) );
  AND2_X1 u2_u10_u5_U86 (.A1( u2_u10_X_31 ) , .A2( u2_u10_X_32 ) , .ZN( u2_u10_u5_n106 ) );
  AND2_X1 u2_u10_u5_U87 (.A1( u2_u10_X_31 ) , .ZN( u2_u10_u5_n109 ) , .A2( u2_u10_u5_n181 ) );
  INV_X1 u2_u10_u5_U88 (.A( u2_u10_X_33 ) , .ZN( u2_u10_u5_n180 ) );
  INV_X1 u2_u10_u5_U89 (.A( u2_u10_X_35 ) , .ZN( u2_u10_u5_n171 ) );
  NOR2_X1 u2_u10_u5_U9 (.ZN( u2_u10_u5_n135 ) , .A1( u2_u10_u5_n173 ) , .A2( u2_u10_u5_n176 ) );
  INV_X1 u2_u10_u5_U90 (.A( u2_u10_X_36 ) , .ZN( u2_u10_u5_n170 ) );
  INV_X1 u2_u10_u5_U91 (.A( u2_u10_X_32 ) , .ZN( u2_u10_u5_n181 ) );
  NAND4_X1 u2_u10_u5_U92 (.ZN( u2_out10_29 ) , .A4( u2_u10_u5_n129 ) , .A3( u2_u10_u5_n130 ) , .A2( u2_u10_u5_n168 ) , .A1( u2_u10_u5_n196 ) );
  AOI221_X1 u2_u10_u5_U93 (.A( u2_u10_u5_n128 ) , .ZN( u2_u10_u5_n129 ) , .C2( u2_u10_u5_n132 ) , .B2( u2_u10_u5_n159 ) , .B1( u2_u10_u5_n176 ) , .C1( u2_u10_u5_n184 ) );
  AOI222_X1 u2_u10_u5_U94 (.ZN( u2_u10_u5_n130 ) , .A2( u2_u10_u5_n146 ) , .B1( u2_u10_u5_n147 ) , .C2( u2_u10_u5_n175 ) , .B2( u2_u10_u5_n179 ) , .A1( u2_u10_u5_n188 ) , .C1( u2_u10_u5_n194 ) );
  NAND4_X1 u2_u10_u5_U95 (.ZN( u2_out10_19 ) , .A4( u2_u10_u5_n166 ) , .A3( u2_u10_u5_n167 ) , .A2( u2_u10_u5_n168 ) , .A1( u2_u10_u5_n169 ) );
  AOI22_X1 u2_u10_u5_U96 (.B2( u2_u10_u5_n145 ) , .A2( u2_u10_u5_n146 ) , .ZN( u2_u10_u5_n167 ) , .B1( u2_u10_u5_n182 ) , .A1( u2_u10_u5_n189 ) );
  NOR4_X1 u2_u10_u5_U97 (.A4( u2_u10_u5_n162 ) , .A3( u2_u10_u5_n163 ) , .A2( u2_u10_u5_n164 ) , .A1( u2_u10_u5_n165 ) , .ZN( u2_u10_u5_n166 ) );
  NAND4_X1 u2_u10_u5_U98 (.ZN( u2_out10_11 ) , .A4( u2_u10_u5_n143 ) , .A3( u2_u10_u5_n144 ) , .A2( u2_u10_u5_n169 ) , .A1( u2_u10_u5_n196 ) );
  AOI22_X1 u2_u10_u5_U99 (.A2( u2_u10_u5_n132 ) , .ZN( u2_u10_u5_n144 ) , .B2( u2_u10_u5_n145 ) , .B1( u2_u10_u5_n184 ) , .A1( u2_u10_u5_n194 ) );
  AOI22_X1 u2_u10_u6_U10 (.A2( u2_u10_u6_n151 ) , .B2( u2_u10_u6_n161 ) , .A1( u2_u10_u6_n167 ) , .B1( u2_u10_u6_n170 ) , .ZN( u2_u10_u6_n89 ) );
  AOI21_X1 u2_u10_u6_U11 (.B1( u2_u10_u6_n107 ) , .B2( u2_u10_u6_n132 ) , .A( u2_u10_u6_n158 ) , .ZN( u2_u10_u6_n88 ) );
  AOI21_X1 u2_u10_u6_U12 (.B2( u2_u10_u6_n147 ) , .B1( u2_u10_u6_n148 ) , .ZN( u2_u10_u6_n149 ) , .A( u2_u10_u6_n158 ) );
  AOI21_X1 u2_u10_u6_U13 (.ZN( u2_u10_u6_n106 ) , .A( u2_u10_u6_n142 ) , .B2( u2_u10_u6_n159 ) , .B1( u2_u10_u6_n164 ) );
  INV_X1 u2_u10_u6_U14 (.A( u2_u10_u6_n155 ) , .ZN( u2_u10_u6_n161 ) );
  INV_X1 u2_u10_u6_U15 (.A( u2_u10_u6_n128 ) , .ZN( u2_u10_u6_n164 ) );
  NAND2_X1 u2_u10_u6_U16 (.ZN( u2_u10_u6_n110 ) , .A1( u2_u10_u6_n122 ) , .A2( u2_u10_u6_n129 ) );
  NAND2_X1 u2_u10_u6_U17 (.ZN( u2_u10_u6_n124 ) , .A2( u2_u10_u6_n146 ) , .A1( u2_u10_u6_n148 ) );
  INV_X1 u2_u10_u6_U18 (.A( u2_u10_u6_n132 ) , .ZN( u2_u10_u6_n171 ) );
  AND2_X1 u2_u10_u6_U19 (.A1( u2_u10_u6_n100 ) , .ZN( u2_u10_u6_n130 ) , .A2( u2_u10_u6_n147 ) );
  INV_X1 u2_u10_u6_U20 (.A( u2_u10_u6_n127 ) , .ZN( u2_u10_u6_n173 ) );
  INV_X1 u2_u10_u6_U21 (.A( u2_u10_u6_n121 ) , .ZN( u2_u10_u6_n167 ) );
  INV_X1 u2_u10_u6_U22 (.A( u2_u10_u6_n100 ) , .ZN( u2_u10_u6_n169 ) );
  INV_X1 u2_u10_u6_U23 (.A( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n170 ) );
  INV_X1 u2_u10_u6_U24 (.A( u2_u10_u6_n113 ) , .ZN( u2_u10_u6_n168 ) );
  AND2_X1 u2_u10_u6_U25 (.A1( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n119 ) , .ZN( u2_u10_u6_n133 ) );
  AND2_X1 u2_u10_u6_U26 (.A2( u2_u10_u6_n121 ) , .A1( u2_u10_u6_n122 ) , .ZN( u2_u10_u6_n131 ) );
  AND3_X1 u2_u10_u6_U27 (.ZN( u2_u10_u6_n120 ) , .A2( u2_u10_u6_n127 ) , .A1( u2_u10_u6_n132 ) , .A3( u2_u10_u6_n145 ) );
  INV_X1 u2_u10_u6_U28 (.A( u2_u10_u6_n146 ) , .ZN( u2_u10_u6_n163 ) );
  AOI222_X1 u2_u10_u6_U29 (.ZN( u2_u10_u6_n114 ) , .A1( u2_u10_u6_n118 ) , .A2( u2_u10_u6_n126 ) , .B2( u2_u10_u6_n151 ) , .C2( u2_u10_u6_n159 ) , .C1( u2_u10_u6_n168 ) , .B1( u2_u10_u6_n169 ) );
  INV_X1 u2_u10_u6_U3 (.A( u2_u10_u6_n110 ) , .ZN( u2_u10_u6_n166 ) );
  NOR2_X1 u2_u10_u6_U30 (.A1( u2_u10_u6_n162 ) , .A2( u2_u10_u6_n165 ) , .ZN( u2_u10_u6_n98 ) );
  AOI211_X1 u2_u10_u6_U31 (.B( u2_u10_u6_n134 ) , .A( u2_u10_u6_n135 ) , .C1( u2_u10_u6_n136 ) , .ZN( u2_u10_u6_n137 ) , .C2( u2_u10_u6_n151 ) );
  NAND4_X1 u2_u10_u6_U32 (.A4( u2_u10_u6_n127 ) , .A3( u2_u10_u6_n128 ) , .A2( u2_u10_u6_n129 ) , .A1( u2_u10_u6_n130 ) , .ZN( u2_u10_u6_n136 ) );
  AOI21_X1 u2_u10_u6_U33 (.B2( u2_u10_u6_n132 ) , .B1( u2_u10_u6_n133 ) , .ZN( u2_u10_u6_n134 ) , .A( u2_u10_u6_n158 ) );
  AOI21_X1 u2_u10_u6_U34 (.B1( u2_u10_u6_n131 ) , .ZN( u2_u10_u6_n135 ) , .A( u2_u10_u6_n144 ) , .B2( u2_u10_u6_n146 ) );
  NAND2_X1 u2_u10_u6_U35 (.A1( u2_u10_u6_n144 ) , .ZN( u2_u10_u6_n151 ) , .A2( u2_u10_u6_n158 ) );
  NAND2_X1 u2_u10_u6_U36 (.ZN( u2_u10_u6_n132 ) , .A1( u2_u10_u6_n91 ) , .A2( u2_u10_u6_n97 ) );
  AOI22_X1 u2_u10_u6_U37 (.B2( u2_u10_u6_n110 ) , .B1( u2_u10_u6_n111 ) , .A1( u2_u10_u6_n112 ) , .ZN( u2_u10_u6_n115 ) , .A2( u2_u10_u6_n161 ) );
  NAND4_X1 u2_u10_u6_U38 (.A3( u2_u10_u6_n109 ) , .ZN( u2_u10_u6_n112 ) , .A4( u2_u10_u6_n132 ) , .A2( u2_u10_u6_n147 ) , .A1( u2_u10_u6_n166 ) );
  NOR2_X1 u2_u10_u6_U39 (.ZN( u2_u10_u6_n109 ) , .A1( u2_u10_u6_n170 ) , .A2( u2_u10_u6_n173 ) );
  INV_X1 u2_u10_u6_U4 (.A( u2_u10_u6_n142 ) , .ZN( u2_u10_u6_n174 ) );
  NOR2_X1 u2_u10_u6_U40 (.A2( u2_u10_u6_n126 ) , .ZN( u2_u10_u6_n155 ) , .A1( u2_u10_u6_n160 ) );
  NAND2_X1 u2_u10_u6_U41 (.ZN( u2_u10_u6_n146 ) , .A2( u2_u10_u6_n94 ) , .A1( u2_u10_u6_n99 ) );
  AOI21_X1 u2_u10_u6_U42 (.A( u2_u10_u6_n144 ) , .B2( u2_u10_u6_n145 ) , .B1( u2_u10_u6_n146 ) , .ZN( u2_u10_u6_n150 ) );
  INV_X1 u2_u10_u6_U43 (.A( u2_u10_u6_n111 ) , .ZN( u2_u10_u6_n158 ) );
  NAND2_X1 u2_u10_u6_U44 (.ZN( u2_u10_u6_n127 ) , .A1( u2_u10_u6_n91 ) , .A2( u2_u10_u6_n92 ) );
  NAND2_X1 u2_u10_u6_U45 (.ZN( u2_u10_u6_n129 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n96 ) );
  INV_X1 u2_u10_u6_U46 (.A( u2_u10_u6_n144 ) , .ZN( u2_u10_u6_n159 ) );
  NAND2_X1 u2_u10_u6_U47 (.ZN( u2_u10_u6_n145 ) , .A2( u2_u10_u6_n97 ) , .A1( u2_u10_u6_n98 ) );
  NAND2_X1 u2_u10_u6_U48 (.ZN( u2_u10_u6_n148 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n94 ) );
  NAND2_X1 u2_u10_u6_U49 (.ZN( u2_u10_u6_n108 ) , .A2( u2_u10_u6_n139 ) , .A1( u2_u10_u6_n144 ) );
  NAND2_X1 u2_u10_u6_U5 (.A2( u2_u10_u6_n143 ) , .ZN( u2_u10_u6_n152 ) , .A1( u2_u10_u6_n166 ) );
  NAND2_X1 u2_u10_u6_U50 (.ZN( u2_u10_u6_n121 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n97 ) );
  NAND2_X1 u2_u10_u6_U51 (.ZN( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n95 ) );
  AND2_X1 u2_u10_u6_U52 (.ZN( u2_u10_u6_n118 ) , .A2( u2_u10_u6_n91 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U53 (.ZN( u2_u10_u6_n147 ) , .A2( u2_u10_u6_n98 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U54 (.ZN( u2_u10_u6_n128 ) , .A1( u2_u10_u6_n94 ) , .A2( u2_u10_u6_n96 ) );
  NAND2_X1 u2_u10_u6_U55 (.ZN( u2_u10_u6_n119 ) , .A2( u2_u10_u6_n95 ) , .A1( u2_u10_u6_n99 ) );
  NAND2_X1 u2_u10_u6_U56 (.ZN( u2_u10_u6_n123 ) , .A2( u2_u10_u6_n91 ) , .A1( u2_u10_u6_n96 ) );
  NAND2_X1 u2_u10_u6_U57 (.ZN( u2_u10_u6_n100 ) , .A2( u2_u10_u6_n92 ) , .A1( u2_u10_u6_n98 ) );
  NAND2_X1 u2_u10_u6_U58 (.ZN( u2_u10_u6_n122 ) , .A1( u2_u10_u6_n94 ) , .A2( u2_u10_u6_n97 ) );
  INV_X1 u2_u10_u6_U59 (.A( u2_u10_u6_n139 ) , .ZN( u2_u10_u6_n160 ) );
  AOI22_X1 u2_u10_u6_U6 (.B2( u2_u10_u6_n101 ) , .A1( u2_u10_u6_n102 ) , .ZN( u2_u10_u6_n103 ) , .B1( u2_u10_u6_n160 ) , .A2( u2_u10_u6_n161 ) );
  NAND2_X1 u2_u10_u6_U60 (.ZN( u2_u10_u6_n113 ) , .A1( u2_u10_u6_n96 ) , .A2( u2_u10_u6_n98 ) );
  NOR2_X1 u2_u10_u6_U61 (.A2( u2_u10_X_40 ) , .A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n126 ) );
  NOR2_X1 u2_u10_u6_U62 (.A2( u2_u10_X_39 ) , .A1( u2_u10_X_42 ) , .ZN( u2_u10_u6_n92 ) );
  NOR2_X1 u2_u10_u6_U63 (.A2( u2_u10_X_39 ) , .A1( u2_u10_u6_n156 ) , .ZN( u2_u10_u6_n97 ) );
  NOR2_X1 u2_u10_u6_U64 (.A2( u2_u10_X_38 ) , .A1( u2_u10_u6_n165 ) , .ZN( u2_u10_u6_n95 ) );
  NOR2_X1 u2_u10_u6_U65 (.A2( u2_u10_X_41 ) , .ZN( u2_u10_u6_n111 ) , .A1( u2_u10_u6_n157 ) );
  NOR2_X1 u2_u10_u6_U66 (.A2( u2_u10_X_37 ) , .A1( u2_u10_u6_n162 ) , .ZN( u2_u10_u6_n94 ) );
  NOR2_X1 u2_u10_u6_U67 (.A2( u2_u10_X_37 ) , .A1( u2_u10_X_38 ) , .ZN( u2_u10_u6_n91 ) );
  NAND2_X1 u2_u10_u6_U68 (.A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n144 ) , .A2( u2_u10_u6_n157 ) );
  NAND2_X1 u2_u10_u6_U69 (.A2( u2_u10_X_40 ) , .A1( u2_u10_X_41 ) , .ZN( u2_u10_u6_n139 ) );
  NOR2_X1 u2_u10_u6_U7 (.A1( u2_u10_u6_n118 ) , .ZN( u2_u10_u6_n143 ) , .A2( u2_u10_u6_n168 ) );
  AND2_X1 u2_u10_u6_U70 (.A1( u2_u10_X_39 ) , .A2( u2_u10_u6_n156 ) , .ZN( u2_u10_u6_n96 ) );
  AND2_X1 u2_u10_u6_U71 (.A1( u2_u10_X_39 ) , .A2( u2_u10_X_42 ) , .ZN( u2_u10_u6_n99 ) );
  INV_X1 u2_u10_u6_U72 (.A( u2_u10_X_40 ) , .ZN( u2_u10_u6_n157 ) );
  INV_X1 u2_u10_u6_U73 (.A( u2_u10_X_37 ) , .ZN( u2_u10_u6_n165 ) );
  INV_X1 u2_u10_u6_U74 (.A( u2_u10_X_38 ) , .ZN( u2_u10_u6_n162 ) );
  INV_X1 u2_u10_u6_U75 (.A( u2_u10_X_42 ) , .ZN( u2_u10_u6_n156 ) );
  NAND4_X1 u2_u10_u6_U76 (.ZN( u2_out10_12 ) , .A4( u2_u10_u6_n114 ) , .A3( u2_u10_u6_n115 ) , .A2( u2_u10_u6_n116 ) , .A1( u2_u10_u6_n117 ) );
  OAI22_X1 u2_u10_u6_U77 (.B2( u2_u10_u6_n111 ) , .ZN( u2_u10_u6_n116 ) , .B1( u2_u10_u6_n126 ) , .A2( u2_u10_u6_n164 ) , .A1( u2_u10_u6_n167 ) );
  OAI21_X1 u2_u10_u6_U78 (.A( u2_u10_u6_n108 ) , .ZN( u2_u10_u6_n117 ) , .B2( u2_u10_u6_n141 ) , .B1( u2_u10_u6_n163 ) );
  NAND4_X1 u2_u10_u6_U79 (.ZN( u2_out10_32 ) , .A4( u2_u10_u6_n103 ) , .A3( u2_u10_u6_n104 ) , .A2( u2_u10_u6_n105 ) , .A1( u2_u10_u6_n106 ) );
  INV_X1 u2_u10_u6_U8 (.ZN( u2_u10_u6_n172 ) , .A( u2_u10_u6_n88 ) );
  AOI22_X1 u2_u10_u6_U80 (.ZN( u2_u10_u6_n105 ) , .A2( u2_u10_u6_n108 ) , .A1( u2_u10_u6_n118 ) , .B2( u2_u10_u6_n126 ) , .B1( u2_u10_u6_n171 ) );
  AOI22_X1 u2_u10_u6_U81 (.ZN( u2_u10_u6_n104 ) , .A1( u2_u10_u6_n111 ) , .B1( u2_u10_u6_n124 ) , .B2( u2_u10_u6_n151 ) , .A2( u2_u10_u6_n93 ) );
  OAI211_X1 u2_u10_u6_U82 (.ZN( u2_out10_7 ) , .B( u2_u10_u6_n153 ) , .C2( u2_u10_u6_n154 ) , .C1( u2_u10_u6_n155 ) , .A( u2_u10_u6_n174 ) );
  NOR3_X1 u2_u10_u6_U83 (.A1( u2_u10_u6_n141 ) , .ZN( u2_u10_u6_n154 ) , .A3( u2_u10_u6_n164 ) , .A2( u2_u10_u6_n171 ) );
  AOI211_X1 u2_u10_u6_U84 (.B( u2_u10_u6_n149 ) , .A( u2_u10_u6_n150 ) , .C2( u2_u10_u6_n151 ) , .C1( u2_u10_u6_n152 ) , .ZN( u2_u10_u6_n153 ) );
  OAI211_X1 u2_u10_u6_U85 (.ZN( u2_out10_22 ) , .B( u2_u10_u6_n137 ) , .A( u2_u10_u6_n138 ) , .C2( u2_u10_u6_n139 ) , .C1( u2_u10_u6_n140 ) );
  AOI22_X1 u2_u10_u6_U86 (.B1( u2_u10_u6_n124 ) , .A2( u2_u10_u6_n125 ) , .A1( u2_u10_u6_n126 ) , .ZN( u2_u10_u6_n138 ) , .B2( u2_u10_u6_n161 ) );
  AND4_X1 u2_u10_u6_U87 (.A3( u2_u10_u6_n119 ) , .A1( u2_u10_u6_n120 ) , .A4( u2_u10_u6_n129 ) , .ZN( u2_u10_u6_n140 ) , .A2( u2_u10_u6_n143 ) );
  NAND3_X1 u2_u10_u6_U88 (.A2( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n125 ) , .A1( u2_u10_u6_n130 ) , .A3( u2_u10_u6_n131 ) );
  NAND3_X1 u2_u10_u6_U89 (.A3( u2_u10_u6_n133 ) , .ZN( u2_u10_u6_n141 ) , .A1( u2_u10_u6_n145 ) , .A2( u2_u10_u6_n148 ) );
  OAI21_X1 u2_u10_u6_U9 (.A( u2_u10_u6_n159 ) , .B1( u2_u10_u6_n169 ) , .B2( u2_u10_u6_n173 ) , .ZN( u2_u10_u6_n90 ) );
  NAND3_X1 u2_u10_u6_U90 (.ZN( u2_u10_u6_n101 ) , .A3( u2_u10_u6_n107 ) , .A2( u2_u10_u6_n121 ) , .A1( u2_u10_u6_n127 ) );
  NAND3_X1 u2_u10_u6_U91 (.ZN( u2_u10_u6_n102 ) , .A3( u2_u10_u6_n130 ) , .A2( u2_u10_u6_n145 ) , .A1( u2_u10_u6_n166 ) );
  NAND3_X1 u2_u10_u6_U92 (.A3( u2_u10_u6_n113 ) , .A1( u2_u10_u6_n119 ) , .A2( u2_u10_u6_n123 ) , .ZN( u2_u10_u6_n93 ) );
  NAND3_X1 u2_u10_u6_U93 (.ZN( u2_u10_u6_n142 ) , .A2( u2_u10_u6_n172 ) , .A3( u2_u10_u6_n89 ) , .A1( u2_u10_u6_n90 ) );
  AND3_X1 u2_u10_u7_U10 (.A3( u2_u10_u7_n110 ) , .A2( u2_u10_u7_n127 ) , .A1( u2_u10_u7_n132 ) , .ZN( u2_u10_u7_n92 ) );
  OAI21_X1 u2_u10_u7_U11 (.A( u2_u10_u7_n161 ) , .B1( u2_u10_u7_n168 ) , .B2( u2_u10_u7_n173 ) , .ZN( u2_u10_u7_n91 ) );
  AOI211_X1 u2_u10_u7_U12 (.A( u2_u10_u7_n117 ) , .ZN( u2_u10_u7_n118 ) , .C2( u2_u10_u7_n126 ) , .C1( u2_u10_u7_n177 ) , .B( u2_u10_u7_n180 ) );
  OAI22_X1 u2_u10_u7_U13 (.B1( u2_u10_u7_n115 ) , .ZN( u2_u10_u7_n117 ) , .A2( u2_u10_u7_n133 ) , .A1( u2_u10_u7_n137 ) , .B2( u2_u10_u7_n162 ) );
  INV_X1 u2_u10_u7_U14 (.A( u2_u10_u7_n116 ) , .ZN( u2_u10_u7_n180 ) );
  NOR3_X1 u2_u10_u7_U15 (.ZN( u2_u10_u7_n115 ) , .A3( u2_u10_u7_n145 ) , .A2( u2_u10_u7_n168 ) , .A1( u2_u10_u7_n169 ) );
  OAI211_X1 u2_u10_u7_U16 (.B( u2_u10_u7_n122 ) , .A( u2_u10_u7_n123 ) , .C2( u2_u10_u7_n124 ) , .ZN( u2_u10_u7_n154 ) , .C1( u2_u10_u7_n162 ) );
  AOI222_X1 u2_u10_u7_U17 (.ZN( u2_u10_u7_n122 ) , .C2( u2_u10_u7_n126 ) , .C1( u2_u10_u7_n145 ) , .B1( u2_u10_u7_n161 ) , .A2( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n170 ) , .A1( u2_u10_u7_n176 ) );
  INV_X1 u2_u10_u7_U18 (.A( u2_u10_u7_n133 ) , .ZN( u2_u10_u7_n176 ) );
  NOR3_X1 u2_u10_u7_U19 (.A2( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n135 ) , .ZN( u2_u10_u7_n136 ) , .A3( u2_u10_u7_n171 ) );
  NOR2_X1 u2_u10_u7_U20 (.A1( u2_u10_u7_n130 ) , .A2( u2_u10_u7_n134 ) , .ZN( u2_u10_u7_n153 ) );
  INV_X1 u2_u10_u7_U21 (.A( u2_u10_u7_n101 ) , .ZN( u2_u10_u7_n165 ) );
  NOR2_X1 u2_u10_u7_U22 (.ZN( u2_u10_u7_n111 ) , .A2( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n169 ) );
  AOI21_X1 u2_u10_u7_U23 (.ZN( u2_u10_u7_n104 ) , .B2( u2_u10_u7_n112 ) , .B1( u2_u10_u7_n127 ) , .A( u2_u10_u7_n164 ) );
  AOI21_X1 u2_u10_u7_U24 (.ZN( u2_u10_u7_n106 ) , .B1( u2_u10_u7_n133 ) , .B2( u2_u10_u7_n146 ) , .A( u2_u10_u7_n162 ) );
  AOI21_X1 u2_u10_u7_U25 (.A( u2_u10_u7_n101 ) , .ZN( u2_u10_u7_n107 ) , .B2( u2_u10_u7_n128 ) , .B1( u2_u10_u7_n175 ) );
  INV_X1 u2_u10_u7_U26 (.A( u2_u10_u7_n138 ) , .ZN( u2_u10_u7_n171 ) );
  INV_X1 u2_u10_u7_U27 (.A( u2_u10_u7_n131 ) , .ZN( u2_u10_u7_n177 ) );
  INV_X1 u2_u10_u7_U28 (.A( u2_u10_u7_n110 ) , .ZN( u2_u10_u7_n174 ) );
  NAND2_X1 u2_u10_u7_U29 (.A1( u2_u10_u7_n129 ) , .A2( u2_u10_u7_n132 ) , .ZN( u2_u10_u7_n149 ) );
  OAI21_X1 u2_u10_u7_U3 (.ZN( u2_u10_u7_n159 ) , .A( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n171 ) , .B1( u2_u10_u7_n174 ) );
  NAND2_X1 u2_u10_u7_U30 (.A1( u2_u10_u7_n113 ) , .A2( u2_u10_u7_n124 ) , .ZN( u2_u10_u7_n130 ) );
  INV_X1 u2_u10_u7_U31 (.A( u2_u10_u7_n112 ) , .ZN( u2_u10_u7_n173 ) );
  INV_X1 u2_u10_u7_U32 (.A( u2_u10_u7_n128 ) , .ZN( u2_u10_u7_n168 ) );
  INV_X1 u2_u10_u7_U33 (.A( u2_u10_u7_n148 ) , .ZN( u2_u10_u7_n169 ) );
  INV_X1 u2_u10_u7_U34 (.A( u2_u10_u7_n127 ) , .ZN( u2_u10_u7_n179 ) );
  NOR2_X1 u2_u10_u7_U35 (.ZN( u2_u10_u7_n101 ) , .A2( u2_u10_u7_n150 ) , .A1( u2_u10_u7_n156 ) );
  AOI211_X1 u2_u10_u7_U36 (.B( u2_u10_u7_n154 ) , .A( u2_u10_u7_n155 ) , .C1( u2_u10_u7_n156 ) , .ZN( u2_u10_u7_n157 ) , .C2( u2_u10_u7_n172 ) );
  INV_X1 u2_u10_u7_U37 (.A( u2_u10_u7_n153 ) , .ZN( u2_u10_u7_n172 ) );
  AOI211_X1 u2_u10_u7_U38 (.B( u2_u10_u7_n139 ) , .A( u2_u10_u7_n140 ) , .C2( u2_u10_u7_n141 ) , .ZN( u2_u10_u7_n142 ) , .C1( u2_u10_u7_n156 ) );
  NAND4_X1 u2_u10_u7_U39 (.A3( u2_u10_u7_n127 ) , .A2( u2_u10_u7_n128 ) , .A1( u2_u10_u7_n129 ) , .ZN( u2_u10_u7_n141 ) , .A4( u2_u10_u7_n147 ) );
  INV_X1 u2_u10_u7_U4 (.A( u2_u10_u7_n111 ) , .ZN( u2_u10_u7_n170 ) );
  AOI21_X1 u2_u10_u7_U40 (.A( u2_u10_u7_n137 ) , .B1( u2_u10_u7_n138 ) , .ZN( u2_u10_u7_n139 ) , .B2( u2_u10_u7_n146 ) );
  OAI22_X1 u2_u10_u7_U41 (.B1( u2_u10_u7_n136 ) , .ZN( u2_u10_u7_n140 ) , .A1( u2_u10_u7_n153 ) , .B2( u2_u10_u7_n162 ) , .A2( u2_u10_u7_n164 ) );
  AOI21_X1 u2_u10_u7_U42 (.ZN( u2_u10_u7_n123 ) , .B1( u2_u10_u7_n165 ) , .B2( u2_u10_u7_n177 ) , .A( u2_u10_u7_n97 ) );
  AOI21_X1 u2_u10_u7_U43 (.B2( u2_u10_u7_n113 ) , .B1( u2_u10_u7_n124 ) , .A( u2_u10_u7_n125 ) , .ZN( u2_u10_u7_n97 ) );
  INV_X1 u2_u10_u7_U44 (.A( u2_u10_u7_n125 ) , .ZN( u2_u10_u7_n161 ) );
  INV_X1 u2_u10_u7_U45 (.A( u2_u10_u7_n152 ) , .ZN( u2_u10_u7_n162 ) );
  AOI22_X1 u2_u10_u7_U46 (.A2( u2_u10_u7_n114 ) , .ZN( u2_u10_u7_n119 ) , .B1( u2_u10_u7_n130 ) , .A1( u2_u10_u7_n156 ) , .B2( u2_u10_u7_n165 ) );
  NAND2_X1 u2_u10_u7_U47 (.A2( u2_u10_u7_n112 ) , .ZN( u2_u10_u7_n114 ) , .A1( u2_u10_u7_n175 ) );
  AND2_X1 u2_u10_u7_U48 (.ZN( u2_u10_u7_n145 ) , .A2( u2_u10_u7_n98 ) , .A1( u2_u10_u7_n99 ) );
  NOR2_X1 u2_u10_u7_U49 (.ZN( u2_u10_u7_n137 ) , .A1( u2_u10_u7_n150 ) , .A2( u2_u10_u7_n161 ) );
  INV_X1 u2_u10_u7_U5 (.A( u2_u10_u7_n149 ) , .ZN( u2_u10_u7_n175 ) );
  AOI21_X1 u2_u10_u7_U50 (.ZN( u2_u10_u7_n105 ) , .B2( u2_u10_u7_n110 ) , .A( u2_u10_u7_n125 ) , .B1( u2_u10_u7_n147 ) );
  NAND2_X1 u2_u10_u7_U51 (.ZN( u2_u10_u7_n146 ) , .A1( u2_u10_u7_n95 ) , .A2( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U52 (.A2( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n147 ) , .A1( u2_u10_u7_n93 ) );
  NAND2_X1 u2_u10_u7_U53 (.A1( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n127 ) , .A2( u2_u10_u7_n99 ) );
  OR2_X1 u2_u10_u7_U54 (.ZN( u2_u10_u7_n126 ) , .A2( u2_u10_u7_n152 ) , .A1( u2_u10_u7_n156 ) );
  NAND2_X1 u2_u10_u7_U55 (.A2( u2_u10_u7_n102 ) , .A1( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n133 ) );
  NAND2_X1 u2_u10_u7_U56 (.ZN( u2_u10_u7_n112 ) , .A2( u2_u10_u7_n96 ) , .A1( u2_u10_u7_n99 ) );
  NAND2_X1 u2_u10_u7_U57 (.A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n128 ) , .A1( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U58 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n113 ) , .A2( u2_u10_u7_n93 ) );
  NAND2_X1 u2_u10_u7_U59 (.A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n124 ) , .A1( u2_u10_u7_n96 ) );
  INV_X1 u2_u10_u7_U6 (.A( u2_u10_u7_n154 ) , .ZN( u2_u10_u7_n178 ) );
  NAND2_X1 u2_u10_u7_U60 (.ZN( u2_u10_u7_n110 ) , .A1( u2_u10_u7_n95 ) , .A2( u2_u10_u7_n96 ) );
  INV_X1 u2_u10_u7_U61 (.A( u2_u10_u7_n150 ) , .ZN( u2_u10_u7_n164 ) );
  AND2_X1 u2_u10_u7_U62 (.ZN( u2_u10_u7_n134 ) , .A1( u2_u10_u7_n93 ) , .A2( u2_u10_u7_n98 ) );
  NAND2_X1 u2_u10_u7_U63 (.A1( u2_u10_u7_n100 ) , .A2( u2_u10_u7_n102 ) , .ZN( u2_u10_u7_n129 ) );
  NAND2_X1 u2_u10_u7_U64 (.A2( u2_u10_u7_n103 ) , .ZN( u2_u10_u7_n131 ) , .A1( u2_u10_u7_n95 ) );
  NAND2_X1 u2_u10_u7_U65 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n138 ) , .A2( u2_u10_u7_n99 ) );
  NAND2_X1 u2_u10_u7_U66 (.ZN( u2_u10_u7_n132 ) , .A1( u2_u10_u7_n93 ) , .A2( u2_u10_u7_n96 ) );
  NAND2_X1 u2_u10_u7_U67 (.A1( u2_u10_u7_n100 ) , .ZN( u2_u10_u7_n148 ) , .A2( u2_u10_u7_n95 ) );
  NOR2_X1 u2_u10_u7_U68 (.A2( u2_u10_X_47 ) , .ZN( u2_u10_u7_n150 ) , .A1( u2_u10_u7_n163 ) );
  NOR2_X1 u2_u10_u7_U69 (.A2( u2_u10_X_43 ) , .A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n103 ) );
  AOI211_X1 u2_u10_u7_U7 (.ZN( u2_u10_u7_n116 ) , .A( u2_u10_u7_n155 ) , .C1( u2_u10_u7_n161 ) , .C2( u2_u10_u7_n171 ) , .B( u2_u10_u7_n94 ) );
  NOR2_X1 u2_u10_u7_U70 (.A2( u2_u10_X_48 ) , .A1( u2_u10_u7_n166 ) , .ZN( u2_u10_u7_n95 ) );
  NOR2_X1 u2_u10_u7_U71 (.A2( u2_u10_X_45 ) , .A1( u2_u10_X_48 ) , .ZN( u2_u10_u7_n99 ) );
  NOR2_X1 u2_u10_u7_U72 (.A2( u2_u10_X_44 ) , .A1( u2_u10_u7_n167 ) , .ZN( u2_u10_u7_n98 ) );
  NOR2_X1 u2_u10_u7_U73 (.A2( u2_u10_X_46 ) , .A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n152 ) );
  AND2_X1 u2_u10_u7_U74 (.A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n156 ) , .A2( u2_u10_u7_n163 ) );
  NAND2_X1 u2_u10_u7_U75 (.A2( u2_u10_X_46 ) , .A1( u2_u10_X_47 ) , .ZN( u2_u10_u7_n125 ) );
  AND2_X1 u2_u10_u7_U76 (.A2( u2_u10_X_45 ) , .A1( u2_u10_X_48 ) , .ZN( u2_u10_u7_n102 ) );
  AND2_X1 u2_u10_u7_U77 (.A2( u2_u10_X_43 ) , .A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n96 ) );
  AND2_X1 u2_u10_u7_U78 (.A1( u2_u10_X_44 ) , .ZN( u2_u10_u7_n100 ) , .A2( u2_u10_u7_n167 ) );
  AND2_X1 u2_u10_u7_U79 (.A1( u2_u10_X_48 ) , .A2( u2_u10_u7_n166 ) , .ZN( u2_u10_u7_n93 ) );
  OAI222_X1 u2_u10_u7_U8 (.C2( u2_u10_u7_n101 ) , .B2( u2_u10_u7_n111 ) , .A1( u2_u10_u7_n113 ) , .C1( u2_u10_u7_n146 ) , .A2( u2_u10_u7_n162 ) , .B1( u2_u10_u7_n164 ) , .ZN( u2_u10_u7_n94 ) );
  INV_X1 u2_u10_u7_U80 (.A( u2_u10_X_46 ) , .ZN( u2_u10_u7_n163 ) );
  INV_X1 u2_u10_u7_U81 (.A( u2_u10_X_43 ) , .ZN( u2_u10_u7_n167 ) );
  INV_X1 u2_u10_u7_U82 (.A( u2_u10_X_45 ) , .ZN( u2_u10_u7_n166 ) );
  NAND4_X1 u2_u10_u7_U83 (.ZN( u2_out10_27 ) , .A4( u2_u10_u7_n118 ) , .A3( u2_u10_u7_n119 ) , .A2( u2_u10_u7_n120 ) , .A1( u2_u10_u7_n121 ) );
  OAI21_X1 u2_u10_u7_U84 (.ZN( u2_u10_u7_n121 ) , .B2( u2_u10_u7_n145 ) , .A( u2_u10_u7_n150 ) , .B1( u2_u10_u7_n174 ) );
  OAI21_X1 u2_u10_u7_U85 (.ZN( u2_u10_u7_n120 ) , .A( u2_u10_u7_n161 ) , .B2( u2_u10_u7_n170 ) , .B1( u2_u10_u7_n179 ) );
  NAND4_X1 u2_u10_u7_U86 (.ZN( u2_out10_21 ) , .A4( u2_u10_u7_n157 ) , .A3( u2_u10_u7_n158 ) , .A2( u2_u10_u7_n159 ) , .A1( u2_u10_u7_n160 ) );
  OAI21_X1 u2_u10_u7_U87 (.B1( u2_u10_u7_n145 ) , .ZN( u2_u10_u7_n160 ) , .A( u2_u10_u7_n161 ) , .B2( u2_u10_u7_n177 ) );
  AOI22_X1 u2_u10_u7_U88 (.B2( u2_u10_u7_n149 ) , .B1( u2_u10_u7_n150 ) , .A2( u2_u10_u7_n151 ) , .A1( u2_u10_u7_n152 ) , .ZN( u2_u10_u7_n158 ) );
  NAND4_X1 u2_u10_u7_U89 (.ZN( u2_out10_15 ) , .A4( u2_u10_u7_n142 ) , .A3( u2_u10_u7_n143 ) , .A2( u2_u10_u7_n144 ) , .A1( u2_u10_u7_n178 ) );
  OAI221_X1 u2_u10_u7_U9 (.C1( u2_u10_u7_n101 ) , .C2( u2_u10_u7_n147 ) , .ZN( u2_u10_u7_n155 ) , .B2( u2_u10_u7_n162 ) , .A( u2_u10_u7_n91 ) , .B1( u2_u10_u7_n92 ) );
  OR2_X1 u2_u10_u7_U90 (.A2( u2_u10_u7_n125 ) , .A1( u2_u10_u7_n129 ) , .ZN( u2_u10_u7_n144 ) );
  AOI22_X1 u2_u10_u7_U91 (.A2( u2_u10_u7_n126 ) , .ZN( u2_u10_u7_n143 ) , .B2( u2_u10_u7_n165 ) , .B1( u2_u10_u7_n173 ) , .A1( u2_u10_u7_n174 ) );
  NAND4_X1 u2_u10_u7_U92 (.ZN( u2_out10_5 ) , .A4( u2_u10_u7_n108 ) , .A3( u2_u10_u7_n109 ) , .A1( u2_u10_u7_n116 ) , .A2( u2_u10_u7_n123 ) );
  AOI22_X1 u2_u10_u7_U93 (.ZN( u2_u10_u7_n109 ) , .A2( u2_u10_u7_n126 ) , .B2( u2_u10_u7_n145 ) , .B1( u2_u10_u7_n156 ) , .A1( u2_u10_u7_n171 ) );
  NOR4_X1 u2_u10_u7_U94 (.A4( u2_u10_u7_n104 ) , .A3( u2_u10_u7_n105 ) , .A2( u2_u10_u7_n106 ) , .A1( u2_u10_u7_n107 ) , .ZN( u2_u10_u7_n108 ) );
  NAND3_X1 u2_u10_u7_U95 (.A3( u2_u10_u7_n146 ) , .A2( u2_u10_u7_n147 ) , .A1( u2_u10_u7_n148 ) , .ZN( u2_u10_u7_n151 ) );
  NAND3_X1 u2_u10_u7_U96 (.A3( u2_u10_u7_n131 ) , .A2( u2_u10_u7_n132 ) , .A1( u2_u10_u7_n133 ) , .ZN( u2_u10_u7_n135 ) );
  XOR2_X1 u2_u11_U10 (.B( u2_K12_45 ) , .A( u2_R10_30 ) , .Z( u2_u11_X_45 ) );
  XOR2_X1 u2_u11_U11 (.B( u2_K12_44 ) , .A( u2_R10_29 ) , .Z( u2_u11_X_44 ) );
  XOR2_X1 u2_u11_U12 (.B( u2_K12_43 ) , .A( u2_R10_28 ) , .Z( u2_u11_X_43 ) );
  XOR2_X1 u2_u11_U13 (.B( u2_K12_42 ) , .A( u2_R10_29 ) , .Z( u2_u11_X_42 ) );
  XOR2_X1 u2_u11_U14 (.B( u2_K12_41 ) , .A( u2_R10_28 ) , .Z( u2_u11_X_41 ) );
  XOR2_X1 u2_u11_U15 (.B( u2_K12_40 ) , .A( u2_R10_27 ) , .Z( u2_u11_X_40 ) );
  XOR2_X1 u2_u11_U17 (.B( u2_K12_39 ) , .A( u2_R10_26 ) , .Z( u2_u11_X_39 ) );
  XOR2_X1 u2_u11_U18 (.B( u2_K12_38 ) , .A( u2_R10_25 ) , .Z( u2_u11_X_38 ) );
  XOR2_X1 u2_u11_U19 (.B( u2_K12_37 ) , .A( u2_R10_24 ) , .Z( u2_u11_X_37 ) );
  XOR2_X1 u2_u11_U20 (.B( u2_K12_36 ) , .A( u2_R10_25 ) , .Z( u2_u11_X_36 ) );
  XOR2_X1 u2_u11_U21 (.B( u2_K12_35 ) , .A( u2_R10_24 ) , .Z( u2_u11_X_35 ) );
  XOR2_X1 u2_u11_U22 (.B( u2_K12_34 ) , .A( u2_R10_23 ) , .Z( u2_u11_X_34 ) );
  XOR2_X1 u2_u11_U23 (.B( u2_K12_33 ) , .A( u2_R10_22 ) , .Z( u2_u11_X_33 ) );
  XOR2_X1 u2_u11_U24 (.B( u2_K12_32 ) , .A( u2_R10_21 ) , .Z( u2_u11_X_32 ) );
  XOR2_X1 u2_u11_U25 (.B( u2_K12_31 ) , .A( u2_R10_20 ) , .Z( u2_u11_X_31 ) );
  XOR2_X1 u2_u11_U26 (.B( u2_K12_30 ) , .A( u2_R10_21 ) , .Z( u2_u11_X_30 ) );
  XOR2_X1 u2_u11_U28 (.B( u2_K12_29 ) , .A( u2_R10_20 ) , .Z( u2_u11_X_29 ) );
  XOR2_X1 u2_u11_U29 (.B( u2_K12_28 ) , .A( u2_R10_19 ) , .Z( u2_u11_X_28 ) );
  XOR2_X1 u2_u11_U30 (.B( u2_K12_27 ) , .A( u2_R10_18 ) , .Z( u2_u11_X_27 ) );
  XOR2_X1 u2_u11_U31 (.B( u2_K12_26 ) , .A( u2_R10_17 ) , .Z( u2_u11_X_26 ) );
  XOR2_X1 u2_u11_U32 (.B( u2_K12_25 ) , .A( u2_R10_16 ) , .Z( u2_u11_X_25 ) );
  XOR2_X1 u2_u11_U33 (.B( u2_K12_24 ) , .A( u2_R10_17 ) , .Z( u2_u11_X_24 ) );
  XOR2_X1 u2_u11_U34 (.B( u2_K12_23 ) , .A( u2_R10_16 ) , .Z( u2_u11_X_23 ) );
  XOR2_X1 u2_u11_U35 (.B( u2_K12_22 ) , .A( u2_R10_15 ) , .Z( u2_u11_X_22 ) );
  XOR2_X1 u2_u11_U36 (.B( u2_K12_21 ) , .A( u2_R10_14 ) , .Z( u2_u11_X_21 ) );
  XOR2_X1 u2_u11_U37 (.B( u2_K12_20 ) , .A( u2_R10_13 ) , .Z( u2_u11_X_20 ) );
  XOR2_X1 u2_u11_U39 (.B( u2_K12_19 ) , .A( u2_R10_12 ) , .Z( u2_u11_X_19 ) );
  XOR2_X1 u2_u11_U7 (.B( u2_K12_48 ) , .A( u2_R10_1 ) , .Z( u2_u11_X_48 ) );
  XOR2_X1 u2_u11_U8 (.B( u2_K12_47 ) , .A( u2_R10_32 ) , .Z( u2_u11_X_47 ) );
  XOR2_X1 u2_u11_U9 (.B( u2_K12_46 ) , .A( u2_R10_31 ) , .Z( u2_u11_X_46 ) );
  OAI211_X1 u2_u11_u3_U10 (.B( u2_u11_u3_n106 ) , .ZN( u2_u11_u3_n119 ) , .C2( u2_u11_u3_n128 ) , .C1( u2_u11_u3_n167 ) , .A( u2_u11_u3_n181 ) );
  INV_X1 u2_u11_u3_U11 (.ZN( u2_u11_u3_n181 ) , .A( u2_u11_u3_n98 ) );
  AOI221_X1 u2_u11_u3_U12 (.C1( u2_u11_u3_n105 ) , .ZN( u2_u11_u3_n106 ) , .A( u2_u11_u3_n131 ) , .B2( u2_u11_u3_n132 ) , .C2( u2_u11_u3_n133 ) , .B1( u2_u11_u3_n169 ) );
  OAI22_X1 u2_u11_u3_U13 (.B1( u2_u11_u3_n113 ) , .A2( u2_u11_u3_n135 ) , .A1( u2_u11_u3_n150 ) , .B2( u2_u11_u3_n164 ) , .ZN( u2_u11_u3_n98 ) );
  AOI22_X1 u2_u11_u3_U14 (.B1( u2_u11_u3_n115 ) , .A2( u2_u11_u3_n116 ) , .ZN( u2_u11_u3_n123 ) , .B2( u2_u11_u3_n133 ) , .A1( u2_u11_u3_n169 ) );
  NAND2_X1 u2_u11_u3_U15 (.ZN( u2_u11_u3_n116 ) , .A2( u2_u11_u3_n151 ) , .A1( u2_u11_u3_n182 ) );
  NOR2_X1 u2_u11_u3_U16 (.ZN( u2_u11_u3_n126 ) , .A2( u2_u11_u3_n150 ) , .A1( u2_u11_u3_n164 ) );
  AOI21_X1 u2_u11_u3_U17 (.ZN( u2_u11_u3_n112 ) , .B2( u2_u11_u3_n146 ) , .B1( u2_u11_u3_n155 ) , .A( u2_u11_u3_n167 ) );
  NAND2_X1 u2_u11_u3_U18 (.A1( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n142 ) , .A2( u2_u11_u3_n164 ) );
  NAND2_X1 u2_u11_u3_U19 (.ZN( u2_u11_u3_n132 ) , .A2( u2_u11_u3_n152 ) , .A1( u2_u11_u3_n156 ) );
  INV_X1 u2_u11_u3_U20 (.A( u2_u11_u3_n133 ) , .ZN( u2_u11_u3_n165 ) );
  AND2_X1 u2_u11_u3_U21 (.A2( u2_u11_u3_n113 ) , .A1( u2_u11_u3_n114 ) , .ZN( u2_u11_u3_n151 ) );
  INV_X1 u2_u11_u3_U22 (.A( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n170 ) );
  NAND2_X1 u2_u11_u3_U23 (.A1( u2_u11_u3_n107 ) , .A2( u2_u11_u3_n108 ) , .ZN( u2_u11_u3_n140 ) );
  NAND2_X1 u2_u11_u3_U24 (.ZN( u2_u11_u3_n117 ) , .A1( u2_u11_u3_n124 ) , .A2( u2_u11_u3_n148 ) );
  NAND2_X1 u2_u11_u3_U25 (.ZN( u2_u11_u3_n143 ) , .A1( u2_u11_u3_n165 ) , .A2( u2_u11_u3_n167 ) );
  INV_X1 u2_u11_u3_U26 (.A( u2_u11_u3_n130 ) , .ZN( u2_u11_u3_n177 ) );
  INV_X1 u2_u11_u3_U27 (.A( u2_u11_u3_n128 ) , .ZN( u2_u11_u3_n176 ) );
  NAND2_X1 u2_u11_u3_U28 (.ZN( u2_u11_u3_n105 ) , .A2( u2_u11_u3_n130 ) , .A1( u2_u11_u3_n155 ) );
  INV_X1 u2_u11_u3_U29 (.A( u2_u11_u3_n155 ) , .ZN( u2_u11_u3_n174 ) );
  INV_X1 u2_u11_u3_U3 (.A( u2_u11_u3_n140 ) , .ZN( u2_u11_u3_n182 ) );
  INV_X1 u2_u11_u3_U30 (.A( u2_u11_u3_n139 ) , .ZN( u2_u11_u3_n185 ) );
  NOR2_X1 u2_u11_u3_U31 (.ZN( u2_u11_u3_n135 ) , .A2( u2_u11_u3_n141 ) , .A1( u2_u11_u3_n169 ) );
  OAI222_X1 u2_u11_u3_U32 (.C2( u2_u11_u3_n107 ) , .A2( u2_u11_u3_n108 ) , .B1( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n138 ) , .B2( u2_u11_u3_n146 ) , .C1( u2_u11_u3_n154 ) , .A1( u2_u11_u3_n164 ) );
  NOR4_X1 u2_u11_u3_U33 (.A4( u2_u11_u3_n157 ) , .A3( u2_u11_u3_n158 ) , .A2( u2_u11_u3_n159 ) , .A1( u2_u11_u3_n160 ) , .ZN( u2_u11_u3_n161 ) );
  AOI21_X1 u2_u11_u3_U34 (.B2( u2_u11_u3_n152 ) , .B1( u2_u11_u3_n153 ) , .ZN( u2_u11_u3_n158 ) , .A( u2_u11_u3_n164 ) );
  AOI21_X1 u2_u11_u3_U35 (.A( u2_u11_u3_n154 ) , .B2( u2_u11_u3_n155 ) , .B1( u2_u11_u3_n156 ) , .ZN( u2_u11_u3_n157 ) );
  AOI21_X1 u2_u11_u3_U36 (.A( u2_u11_u3_n149 ) , .B2( u2_u11_u3_n150 ) , .B1( u2_u11_u3_n151 ) , .ZN( u2_u11_u3_n159 ) );
  AOI211_X1 u2_u11_u3_U37 (.ZN( u2_u11_u3_n109 ) , .A( u2_u11_u3_n119 ) , .C2( u2_u11_u3_n129 ) , .B( u2_u11_u3_n138 ) , .C1( u2_u11_u3_n141 ) );
  AOI211_X1 u2_u11_u3_U38 (.B( u2_u11_u3_n119 ) , .A( u2_u11_u3_n120 ) , .C2( u2_u11_u3_n121 ) , .ZN( u2_u11_u3_n122 ) , .C1( u2_u11_u3_n179 ) );
  INV_X1 u2_u11_u3_U39 (.A( u2_u11_u3_n156 ) , .ZN( u2_u11_u3_n179 ) );
  INV_X1 u2_u11_u3_U4 (.A( u2_u11_u3_n129 ) , .ZN( u2_u11_u3_n183 ) );
  OAI22_X1 u2_u11_u3_U40 (.B1( u2_u11_u3_n118 ) , .ZN( u2_u11_u3_n120 ) , .A1( u2_u11_u3_n135 ) , .B2( u2_u11_u3_n154 ) , .A2( u2_u11_u3_n178 ) );
  AND3_X1 u2_u11_u3_U41 (.ZN( u2_u11_u3_n118 ) , .A2( u2_u11_u3_n124 ) , .A1( u2_u11_u3_n144 ) , .A3( u2_u11_u3_n152 ) );
  INV_X1 u2_u11_u3_U42 (.A( u2_u11_u3_n121 ) , .ZN( u2_u11_u3_n164 ) );
  NAND2_X1 u2_u11_u3_U43 (.ZN( u2_u11_u3_n133 ) , .A1( u2_u11_u3_n154 ) , .A2( u2_u11_u3_n164 ) );
  NOR2_X1 u2_u11_u3_U44 (.A1( u2_u11_u3_n113 ) , .ZN( u2_u11_u3_n131 ) , .A2( u2_u11_u3_n154 ) );
  NAND2_X1 u2_u11_u3_U45 (.A1( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n150 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U46 (.A2( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n155 ) , .A1( u2_u11_u3_n97 ) );
  OAI211_X1 u2_u11_u3_U47 (.B( u2_u11_u3_n127 ) , .ZN( u2_u11_u3_n139 ) , .C1( u2_u11_u3_n150 ) , .C2( u2_u11_u3_n154 ) , .A( u2_u11_u3_n184 ) );
  INV_X1 u2_u11_u3_U48 (.A( u2_u11_u3_n125 ) , .ZN( u2_u11_u3_n184 ) );
  AOI221_X1 u2_u11_u3_U49 (.A( u2_u11_u3_n126 ) , .ZN( u2_u11_u3_n127 ) , .C2( u2_u11_u3_n132 ) , .C1( u2_u11_u3_n169 ) , .B2( u2_u11_u3_n170 ) , .B1( u2_u11_u3_n174 ) );
  INV_X1 u2_u11_u3_U5 (.A( u2_u11_u3_n117 ) , .ZN( u2_u11_u3_n178 ) );
  OAI22_X1 u2_u11_u3_U50 (.A1( u2_u11_u3_n124 ) , .ZN( u2_u11_u3_n125 ) , .B2( u2_u11_u3_n145 ) , .A2( u2_u11_u3_n165 ) , .B1( u2_u11_u3_n167 ) );
  INV_X1 u2_u11_u3_U51 (.A( u2_u11_u3_n141 ) , .ZN( u2_u11_u3_n167 ) );
  AOI21_X1 u2_u11_u3_U52 (.B2( u2_u11_u3_n114 ) , .B1( u2_u11_u3_n146 ) , .A( u2_u11_u3_n154 ) , .ZN( u2_u11_u3_n94 ) );
  AOI21_X1 u2_u11_u3_U53 (.ZN( u2_u11_u3_n110 ) , .B2( u2_u11_u3_n142 ) , .B1( u2_u11_u3_n186 ) , .A( u2_u11_u3_n95 ) );
  INV_X1 u2_u11_u3_U54 (.A( u2_u11_u3_n145 ) , .ZN( u2_u11_u3_n186 ) );
  AOI21_X1 u2_u11_u3_U55 (.B1( u2_u11_u3_n124 ) , .A( u2_u11_u3_n149 ) , .B2( u2_u11_u3_n155 ) , .ZN( u2_u11_u3_n95 ) );
  INV_X1 u2_u11_u3_U56 (.A( u2_u11_u3_n149 ) , .ZN( u2_u11_u3_n169 ) );
  NAND2_X1 u2_u11_u3_U57 (.ZN( u2_u11_u3_n124 ) , .A1( u2_u11_u3_n96 ) , .A2( u2_u11_u3_n97 ) );
  NAND2_X1 u2_u11_u3_U58 (.A2( u2_u11_u3_n100 ) , .ZN( u2_u11_u3_n146 ) , .A1( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U59 (.A1( u2_u11_u3_n101 ) , .ZN( u2_u11_u3_n145 ) , .A2( u2_u11_u3_n99 ) );
  AOI221_X1 u2_u11_u3_U6 (.A( u2_u11_u3_n131 ) , .C2( u2_u11_u3_n132 ) , .C1( u2_u11_u3_n133 ) , .ZN( u2_u11_u3_n134 ) , .B1( u2_u11_u3_n143 ) , .B2( u2_u11_u3_n177 ) );
  NAND2_X1 u2_u11_u3_U60 (.A1( u2_u11_u3_n100 ) , .ZN( u2_u11_u3_n156 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U61 (.A2( u2_u11_u3_n101 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n148 ) );
  NAND2_X1 u2_u11_u3_U62 (.A1( u2_u11_u3_n100 ) , .A2( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n128 ) );
  NAND2_X1 u2_u11_u3_U63 (.A2( u2_u11_u3_n101 ) , .A1( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n152 ) );
  NAND2_X1 u2_u11_u3_U64 (.A2( u2_u11_u3_n101 ) , .ZN( u2_u11_u3_n114 ) , .A1( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U65 (.ZN( u2_u11_u3_n107 ) , .A1( u2_u11_u3_n97 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U66 (.A2( u2_u11_u3_n100 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n113 ) );
  NAND2_X1 u2_u11_u3_U67 (.A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n153 ) , .A2( u2_u11_u3_n97 ) );
  NAND2_X1 u2_u11_u3_U68 (.A2( u2_u11_u3_n103 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n130 ) );
  NAND2_X1 u2_u11_u3_U69 (.A2( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n144 ) , .A1( u2_u11_u3_n96 ) );
  OAI22_X1 u2_u11_u3_U7 (.B2( u2_u11_u3_n147 ) , .A2( u2_u11_u3_n148 ) , .ZN( u2_u11_u3_n160 ) , .B1( u2_u11_u3_n165 ) , .A1( u2_u11_u3_n168 ) );
  NAND2_X1 u2_u11_u3_U70 (.A1( u2_u11_u3_n102 ) , .A2( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n108 ) );
  NOR2_X1 u2_u11_u3_U71 (.A2( u2_u11_X_19 ) , .A1( u2_u11_X_20 ) , .ZN( u2_u11_u3_n99 ) );
  NOR2_X1 u2_u11_u3_U72 (.A2( u2_u11_X_21 ) , .A1( u2_u11_X_24 ) , .ZN( u2_u11_u3_n103 ) );
  NOR2_X1 u2_u11_u3_U73 (.A2( u2_u11_X_24 ) , .A1( u2_u11_u3_n171 ) , .ZN( u2_u11_u3_n97 ) );
  NOR2_X1 u2_u11_u3_U74 (.A2( u2_u11_X_23 ) , .ZN( u2_u11_u3_n141 ) , .A1( u2_u11_u3_n166 ) );
  NOR2_X1 u2_u11_u3_U75 (.A2( u2_u11_X_19 ) , .A1( u2_u11_u3_n172 ) , .ZN( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U76 (.A1( u2_u11_X_22 ) , .A2( u2_u11_X_23 ) , .ZN( u2_u11_u3_n154 ) );
  NAND2_X1 u2_u11_u3_U77 (.A1( u2_u11_X_23 ) , .ZN( u2_u11_u3_n149 ) , .A2( u2_u11_u3_n166 ) );
  NOR2_X1 u2_u11_u3_U78 (.A2( u2_u11_X_22 ) , .A1( u2_u11_X_23 ) , .ZN( u2_u11_u3_n121 ) );
  AND2_X1 u2_u11_u3_U79 (.A1( u2_u11_X_24 ) , .ZN( u2_u11_u3_n101 ) , .A2( u2_u11_u3_n171 ) );
  AND3_X1 u2_u11_u3_U8 (.A3( u2_u11_u3_n144 ) , .A2( u2_u11_u3_n145 ) , .A1( u2_u11_u3_n146 ) , .ZN( u2_u11_u3_n147 ) );
  AND2_X1 u2_u11_u3_U80 (.A1( u2_u11_X_19 ) , .ZN( u2_u11_u3_n102 ) , .A2( u2_u11_u3_n172 ) );
  AND2_X1 u2_u11_u3_U81 (.A1( u2_u11_X_21 ) , .A2( u2_u11_X_24 ) , .ZN( u2_u11_u3_n100 ) );
  AND2_X1 u2_u11_u3_U82 (.A2( u2_u11_X_19 ) , .A1( u2_u11_X_20 ) , .ZN( u2_u11_u3_n104 ) );
  INV_X1 u2_u11_u3_U83 (.A( u2_u11_X_22 ) , .ZN( u2_u11_u3_n166 ) );
  INV_X1 u2_u11_u3_U84 (.A( u2_u11_X_21 ) , .ZN( u2_u11_u3_n171 ) );
  INV_X1 u2_u11_u3_U85 (.A( u2_u11_X_20 ) , .ZN( u2_u11_u3_n172 ) );
  NAND4_X1 u2_u11_u3_U86 (.ZN( u2_out11_26 ) , .A4( u2_u11_u3_n109 ) , .A3( u2_u11_u3_n110 ) , .A2( u2_u11_u3_n111 ) , .A1( u2_u11_u3_n173 ) );
  INV_X1 u2_u11_u3_U87 (.ZN( u2_u11_u3_n173 ) , .A( u2_u11_u3_n94 ) );
  OAI21_X1 u2_u11_u3_U88 (.ZN( u2_u11_u3_n111 ) , .B2( u2_u11_u3_n117 ) , .A( u2_u11_u3_n133 ) , .B1( u2_u11_u3_n176 ) );
  NAND4_X1 u2_u11_u3_U89 (.ZN( u2_out11_20 ) , .A4( u2_u11_u3_n122 ) , .A3( u2_u11_u3_n123 ) , .A1( u2_u11_u3_n175 ) , .A2( u2_u11_u3_n180 ) );
  INV_X1 u2_u11_u3_U9 (.A( u2_u11_u3_n143 ) , .ZN( u2_u11_u3_n168 ) );
  INV_X1 u2_u11_u3_U90 (.A( u2_u11_u3_n126 ) , .ZN( u2_u11_u3_n180 ) );
  INV_X1 u2_u11_u3_U91 (.A( u2_u11_u3_n112 ) , .ZN( u2_u11_u3_n175 ) );
  NAND4_X1 u2_u11_u3_U92 (.ZN( u2_out11_1 ) , .A4( u2_u11_u3_n161 ) , .A3( u2_u11_u3_n162 ) , .A2( u2_u11_u3_n163 ) , .A1( u2_u11_u3_n185 ) );
  NAND2_X1 u2_u11_u3_U93 (.ZN( u2_u11_u3_n163 ) , .A2( u2_u11_u3_n170 ) , .A1( u2_u11_u3_n176 ) );
  AOI22_X1 u2_u11_u3_U94 (.B2( u2_u11_u3_n140 ) , .B1( u2_u11_u3_n141 ) , .A2( u2_u11_u3_n142 ) , .ZN( u2_u11_u3_n162 ) , .A1( u2_u11_u3_n177 ) );
  OAI222_X1 u2_u11_u3_U95 (.C1( u2_u11_u3_n128 ) , .ZN( u2_u11_u3_n137 ) , .B1( u2_u11_u3_n148 ) , .A2( u2_u11_u3_n150 ) , .B2( u2_u11_u3_n154 ) , .C2( u2_u11_u3_n164 ) , .A1( u2_u11_u3_n167 ) );
  OR4_X1 u2_u11_u3_U96 (.ZN( u2_out11_10 ) , .A4( u2_u11_u3_n136 ) , .A3( u2_u11_u3_n137 ) , .A1( u2_u11_u3_n138 ) , .A2( u2_u11_u3_n139 ) );
  OAI221_X1 u2_u11_u3_U97 (.A( u2_u11_u3_n134 ) , .B2( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n136 ) , .C1( u2_u11_u3_n149 ) , .B1( u2_u11_u3_n151 ) , .C2( u2_u11_u3_n183 ) );
  NAND3_X1 u2_u11_u3_U98 (.A1( u2_u11_u3_n114 ) , .ZN( u2_u11_u3_n115 ) , .A2( u2_u11_u3_n145 ) , .A3( u2_u11_u3_n153 ) );
  NAND3_X1 u2_u11_u3_U99 (.ZN( u2_u11_u3_n129 ) , .A2( u2_u11_u3_n144 ) , .A1( u2_u11_u3_n153 ) , .A3( u2_u11_u3_n182 ) );
  OAI22_X1 u2_u11_u4_U10 (.B2( u2_u11_u4_n135 ) , .ZN( u2_u11_u4_n137 ) , .B1( u2_u11_u4_n153 ) , .A1( u2_u11_u4_n155 ) , .A2( u2_u11_u4_n171 ) );
  AND3_X1 u2_u11_u4_U11 (.A2( u2_u11_u4_n134 ) , .ZN( u2_u11_u4_n135 ) , .A3( u2_u11_u4_n145 ) , .A1( u2_u11_u4_n157 ) );
  NAND2_X1 u2_u11_u4_U12 (.ZN( u2_u11_u4_n132 ) , .A2( u2_u11_u4_n170 ) , .A1( u2_u11_u4_n173 ) );
  AOI21_X1 u2_u11_u4_U13 (.B2( u2_u11_u4_n160 ) , .B1( u2_u11_u4_n161 ) , .ZN( u2_u11_u4_n162 ) , .A( u2_u11_u4_n170 ) );
  AOI21_X1 u2_u11_u4_U14 (.ZN( u2_u11_u4_n107 ) , .B2( u2_u11_u4_n143 ) , .A( u2_u11_u4_n174 ) , .B1( u2_u11_u4_n184 ) );
  AOI21_X1 u2_u11_u4_U15 (.B2( u2_u11_u4_n158 ) , .B1( u2_u11_u4_n159 ) , .ZN( u2_u11_u4_n163 ) , .A( u2_u11_u4_n174 ) );
  AOI21_X1 u2_u11_u4_U16 (.A( u2_u11_u4_n153 ) , .B2( u2_u11_u4_n154 ) , .B1( u2_u11_u4_n155 ) , .ZN( u2_u11_u4_n165 ) );
  AOI21_X1 u2_u11_u4_U17 (.A( u2_u11_u4_n156 ) , .B2( u2_u11_u4_n157 ) , .ZN( u2_u11_u4_n164 ) , .B1( u2_u11_u4_n184 ) );
  INV_X1 u2_u11_u4_U18 (.A( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n170 ) );
  AND2_X1 u2_u11_u4_U19 (.A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n155 ) , .A1( u2_u11_u4_n160 ) );
  INV_X1 u2_u11_u4_U20 (.A( u2_u11_u4_n156 ) , .ZN( u2_u11_u4_n175 ) );
  NAND2_X1 u2_u11_u4_U21 (.A2( u2_u11_u4_n118 ) , .ZN( u2_u11_u4_n131 ) , .A1( u2_u11_u4_n147 ) );
  NAND2_X1 u2_u11_u4_U22 (.A1( u2_u11_u4_n119 ) , .A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n130 ) );
  NAND2_X1 u2_u11_u4_U23 (.ZN( u2_u11_u4_n117 ) , .A2( u2_u11_u4_n118 ) , .A1( u2_u11_u4_n148 ) );
  NAND2_X1 u2_u11_u4_U24 (.ZN( u2_u11_u4_n129 ) , .A1( u2_u11_u4_n134 ) , .A2( u2_u11_u4_n148 ) );
  AND3_X1 u2_u11_u4_U25 (.A1( u2_u11_u4_n119 ) , .A2( u2_u11_u4_n143 ) , .A3( u2_u11_u4_n154 ) , .ZN( u2_u11_u4_n161 ) );
  AND2_X1 u2_u11_u4_U26 (.A1( u2_u11_u4_n145 ) , .A2( u2_u11_u4_n147 ) , .ZN( u2_u11_u4_n159 ) );
  OR3_X1 u2_u11_u4_U27 (.A3( u2_u11_u4_n114 ) , .A2( u2_u11_u4_n115 ) , .A1( u2_u11_u4_n116 ) , .ZN( u2_u11_u4_n136 ) );
  AOI21_X1 u2_u11_u4_U28 (.A( u2_u11_u4_n113 ) , .ZN( u2_u11_u4_n116 ) , .B2( u2_u11_u4_n173 ) , .B1( u2_u11_u4_n174 ) );
  AOI21_X1 u2_u11_u4_U29 (.ZN( u2_u11_u4_n115 ) , .B2( u2_u11_u4_n145 ) , .B1( u2_u11_u4_n146 ) , .A( u2_u11_u4_n156 ) );
  NOR2_X1 u2_u11_u4_U3 (.ZN( u2_u11_u4_n121 ) , .A1( u2_u11_u4_n181 ) , .A2( u2_u11_u4_n182 ) );
  OAI22_X1 u2_u11_u4_U30 (.ZN( u2_u11_u4_n114 ) , .A2( u2_u11_u4_n121 ) , .B1( u2_u11_u4_n160 ) , .B2( u2_u11_u4_n170 ) , .A1( u2_u11_u4_n171 ) );
  INV_X1 u2_u11_u4_U31 (.A( u2_u11_u4_n158 ) , .ZN( u2_u11_u4_n182 ) );
  INV_X1 u2_u11_u4_U32 (.ZN( u2_u11_u4_n181 ) , .A( u2_u11_u4_n96 ) );
  INV_X1 u2_u11_u4_U33 (.A( u2_u11_u4_n144 ) , .ZN( u2_u11_u4_n179 ) );
  INV_X1 u2_u11_u4_U34 (.A( u2_u11_u4_n157 ) , .ZN( u2_u11_u4_n178 ) );
  NAND2_X1 u2_u11_u4_U35 (.A2( u2_u11_u4_n154 ) , .A1( u2_u11_u4_n96 ) , .ZN( u2_u11_u4_n97 ) );
  INV_X1 u2_u11_u4_U36 (.ZN( u2_u11_u4_n186 ) , .A( u2_u11_u4_n95 ) );
  OAI221_X1 u2_u11_u4_U37 (.C1( u2_u11_u4_n134 ) , .B1( u2_u11_u4_n158 ) , .B2( u2_u11_u4_n171 ) , .C2( u2_u11_u4_n173 ) , .A( u2_u11_u4_n94 ) , .ZN( u2_u11_u4_n95 ) );
  AOI222_X1 u2_u11_u4_U38 (.B2( u2_u11_u4_n132 ) , .A1( u2_u11_u4_n138 ) , .C2( u2_u11_u4_n175 ) , .A2( u2_u11_u4_n179 ) , .C1( u2_u11_u4_n181 ) , .B1( u2_u11_u4_n185 ) , .ZN( u2_u11_u4_n94 ) );
  INV_X1 u2_u11_u4_U39 (.A( u2_u11_u4_n113 ) , .ZN( u2_u11_u4_n185 ) );
  INV_X1 u2_u11_u4_U4 (.A( u2_u11_u4_n117 ) , .ZN( u2_u11_u4_n184 ) );
  INV_X1 u2_u11_u4_U40 (.A( u2_u11_u4_n143 ) , .ZN( u2_u11_u4_n183 ) );
  NOR2_X1 u2_u11_u4_U41 (.ZN( u2_u11_u4_n138 ) , .A1( u2_u11_u4_n168 ) , .A2( u2_u11_u4_n169 ) );
  NOR2_X1 u2_u11_u4_U42 (.A1( u2_u11_u4_n150 ) , .A2( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n153 ) );
  NOR2_X1 u2_u11_u4_U43 (.A2( u2_u11_u4_n128 ) , .A1( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n156 ) );
  AOI22_X1 u2_u11_u4_U44 (.B2( u2_u11_u4_n122 ) , .A1( u2_u11_u4_n123 ) , .ZN( u2_u11_u4_n124 ) , .B1( u2_u11_u4_n128 ) , .A2( u2_u11_u4_n172 ) );
  INV_X1 u2_u11_u4_U45 (.A( u2_u11_u4_n153 ) , .ZN( u2_u11_u4_n172 ) );
  NAND2_X1 u2_u11_u4_U46 (.A2( u2_u11_u4_n120 ) , .ZN( u2_u11_u4_n123 ) , .A1( u2_u11_u4_n161 ) );
  AOI22_X1 u2_u11_u4_U47 (.B2( u2_u11_u4_n132 ) , .A2( u2_u11_u4_n133 ) , .ZN( u2_u11_u4_n140 ) , .A1( u2_u11_u4_n150 ) , .B1( u2_u11_u4_n179 ) );
  NAND2_X1 u2_u11_u4_U48 (.ZN( u2_u11_u4_n133 ) , .A2( u2_u11_u4_n146 ) , .A1( u2_u11_u4_n154 ) );
  NAND2_X1 u2_u11_u4_U49 (.A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n154 ) , .A2( u2_u11_u4_n98 ) );
  NOR4_X1 u2_u11_u4_U5 (.A4( u2_u11_u4_n106 ) , .A3( u2_u11_u4_n107 ) , .A2( u2_u11_u4_n108 ) , .A1( u2_u11_u4_n109 ) , .ZN( u2_u11_u4_n110 ) );
  NAND2_X1 u2_u11_u4_U50 (.A1( u2_u11_u4_n101 ) , .ZN( u2_u11_u4_n158 ) , .A2( u2_u11_u4_n99 ) );
  AOI21_X1 u2_u11_u4_U51 (.ZN( u2_u11_u4_n127 ) , .A( u2_u11_u4_n136 ) , .B2( u2_u11_u4_n150 ) , .B1( u2_u11_u4_n180 ) );
  INV_X1 u2_u11_u4_U52 (.A( u2_u11_u4_n160 ) , .ZN( u2_u11_u4_n180 ) );
  NAND2_X1 u2_u11_u4_U53 (.A2( u2_u11_u4_n104 ) , .A1( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n146 ) );
  NAND2_X1 u2_u11_u4_U54 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n160 ) );
  NAND2_X1 u2_u11_u4_U55 (.ZN( u2_u11_u4_n134 ) , .A1( u2_u11_u4_n98 ) , .A2( u2_u11_u4_n99 ) );
  NAND2_X1 u2_u11_u4_U56 (.A1( u2_u11_u4_n103 ) , .A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n143 ) );
  NAND2_X1 u2_u11_u4_U57 (.A2( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n145 ) , .A1( u2_u11_u4_n98 ) );
  NAND2_X1 u2_u11_u4_U58 (.A1( u2_u11_u4_n100 ) , .A2( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n120 ) );
  NAND2_X1 u2_u11_u4_U59 (.A1( u2_u11_u4_n102 ) , .A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n148 ) );
  AOI21_X1 u2_u11_u4_U6 (.ZN( u2_u11_u4_n106 ) , .B2( u2_u11_u4_n146 ) , .B1( u2_u11_u4_n158 ) , .A( u2_u11_u4_n170 ) );
  NAND2_X1 u2_u11_u4_U60 (.A2( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n157 ) );
  INV_X1 u2_u11_u4_U61 (.A( u2_u11_u4_n150 ) , .ZN( u2_u11_u4_n173 ) );
  INV_X1 u2_u11_u4_U62 (.A( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n171 ) );
  NAND2_X1 u2_u11_u4_U63 (.A1( u2_u11_u4_n100 ) , .ZN( u2_u11_u4_n118 ) , .A2( u2_u11_u4_n99 ) );
  NAND2_X1 u2_u11_u4_U64 (.A2( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n144 ) );
  NAND2_X1 u2_u11_u4_U65 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n105 ) , .ZN( u2_u11_u4_n96 ) );
  INV_X1 u2_u11_u4_U66 (.A( u2_u11_u4_n128 ) , .ZN( u2_u11_u4_n174 ) );
  NAND2_X1 u2_u11_u4_U67 (.A2( u2_u11_u4_n102 ) , .ZN( u2_u11_u4_n119 ) , .A1( u2_u11_u4_n98 ) );
  NAND2_X1 u2_u11_u4_U68 (.A2( u2_u11_u4_n101 ) , .A1( u2_u11_u4_n103 ) , .ZN( u2_u11_u4_n147 ) );
  NAND2_X1 u2_u11_u4_U69 (.A2( u2_u11_u4_n104 ) , .ZN( u2_u11_u4_n113 ) , .A1( u2_u11_u4_n99 ) );
  AOI21_X1 u2_u11_u4_U7 (.ZN( u2_u11_u4_n108 ) , .B2( u2_u11_u4_n134 ) , .B1( u2_u11_u4_n155 ) , .A( u2_u11_u4_n156 ) );
  NOR2_X1 u2_u11_u4_U70 (.A2( u2_u11_X_28 ) , .ZN( u2_u11_u4_n150 ) , .A1( u2_u11_u4_n168 ) );
  NOR2_X1 u2_u11_u4_U71 (.A2( u2_u11_X_29 ) , .ZN( u2_u11_u4_n152 ) , .A1( u2_u11_u4_n169 ) );
  NOR2_X1 u2_u11_u4_U72 (.A2( u2_u11_X_26 ) , .ZN( u2_u11_u4_n100 ) , .A1( u2_u11_u4_n177 ) );
  NOR2_X1 u2_u11_u4_U73 (.A2( u2_u11_X_30 ) , .ZN( u2_u11_u4_n105 ) , .A1( u2_u11_u4_n176 ) );
  NOR2_X1 u2_u11_u4_U74 (.A2( u2_u11_X_28 ) , .A1( u2_u11_X_29 ) , .ZN( u2_u11_u4_n128 ) );
  NOR2_X1 u2_u11_u4_U75 (.A2( u2_u11_X_25 ) , .A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n98 ) );
  NOR2_X1 u2_u11_u4_U76 (.A2( u2_u11_X_27 ) , .A1( u2_u11_X_30 ) , .ZN( u2_u11_u4_n102 ) );
  AND2_X1 u2_u11_u4_U77 (.A2( u2_u11_X_25 ) , .A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n104 ) );
  AND2_X1 u2_u11_u4_U78 (.A1( u2_u11_X_30 ) , .A2( u2_u11_u4_n176 ) , .ZN( u2_u11_u4_n99 ) );
  AND2_X1 u2_u11_u4_U79 (.A1( u2_u11_X_26 ) , .ZN( u2_u11_u4_n101 ) , .A2( u2_u11_u4_n177 ) );
  AOI21_X1 u2_u11_u4_U8 (.ZN( u2_u11_u4_n109 ) , .A( u2_u11_u4_n153 ) , .B1( u2_u11_u4_n159 ) , .B2( u2_u11_u4_n184 ) );
  AND2_X1 u2_u11_u4_U80 (.A1( u2_u11_X_27 ) , .A2( u2_u11_X_30 ) , .ZN( u2_u11_u4_n103 ) );
  INV_X1 u2_u11_u4_U81 (.A( u2_u11_X_28 ) , .ZN( u2_u11_u4_n169 ) );
  INV_X1 u2_u11_u4_U82 (.A( u2_u11_X_29 ) , .ZN( u2_u11_u4_n168 ) );
  INV_X1 u2_u11_u4_U83 (.A( u2_u11_X_25 ) , .ZN( u2_u11_u4_n177 ) );
  INV_X1 u2_u11_u4_U84 (.A( u2_u11_X_27 ) , .ZN( u2_u11_u4_n176 ) );
  NAND4_X1 u2_u11_u4_U85 (.ZN( u2_out11_25 ) , .A4( u2_u11_u4_n139 ) , .A3( u2_u11_u4_n140 ) , .A2( u2_u11_u4_n141 ) , .A1( u2_u11_u4_n142 ) );
  OAI21_X1 u2_u11_u4_U86 (.A( u2_u11_u4_n128 ) , .B2( u2_u11_u4_n129 ) , .B1( u2_u11_u4_n130 ) , .ZN( u2_u11_u4_n142 ) );
  OAI21_X1 u2_u11_u4_U87 (.B2( u2_u11_u4_n131 ) , .ZN( u2_u11_u4_n141 ) , .A( u2_u11_u4_n175 ) , .B1( u2_u11_u4_n183 ) );
  NAND4_X1 u2_u11_u4_U88 (.ZN( u2_out11_14 ) , .A4( u2_u11_u4_n124 ) , .A3( u2_u11_u4_n125 ) , .A2( u2_u11_u4_n126 ) , .A1( u2_u11_u4_n127 ) );
  AOI22_X1 u2_u11_u4_U89 (.B2( u2_u11_u4_n117 ) , .ZN( u2_u11_u4_n126 ) , .A1( u2_u11_u4_n129 ) , .B1( u2_u11_u4_n152 ) , .A2( u2_u11_u4_n175 ) );
  AOI211_X1 u2_u11_u4_U9 (.B( u2_u11_u4_n136 ) , .A( u2_u11_u4_n137 ) , .C2( u2_u11_u4_n138 ) , .ZN( u2_u11_u4_n139 ) , .C1( u2_u11_u4_n182 ) );
  AOI22_X1 u2_u11_u4_U90 (.ZN( u2_u11_u4_n125 ) , .B2( u2_u11_u4_n131 ) , .A2( u2_u11_u4_n132 ) , .B1( u2_u11_u4_n138 ) , .A1( u2_u11_u4_n178 ) );
  NAND4_X1 u2_u11_u4_U91 (.ZN( u2_out11_8 ) , .A4( u2_u11_u4_n110 ) , .A3( u2_u11_u4_n111 ) , .A2( u2_u11_u4_n112 ) , .A1( u2_u11_u4_n186 ) );
  NAND2_X1 u2_u11_u4_U92 (.ZN( u2_u11_u4_n112 ) , .A2( u2_u11_u4_n130 ) , .A1( u2_u11_u4_n150 ) );
  AOI22_X1 u2_u11_u4_U93 (.ZN( u2_u11_u4_n111 ) , .B2( u2_u11_u4_n132 ) , .A1( u2_u11_u4_n152 ) , .B1( u2_u11_u4_n178 ) , .A2( u2_u11_u4_n97 ) );
  AOI22_X1 u2_u11_u4_U94 (.B2( u2_u11_u4_n149 ) , .B1( u2_u11_u4_n150 ) , .A2( u2_u11_u4_n151 ) , .A1( u2_u11_u4_n152 ) , .ZN( u2_u11_u4_n167 ) );
  NOR4_X1 u2_u11_u4_U95 (.A4( u2_u11_u4_n162 ) , .A3( u2_u11_u4_n163 ) , .A2( u2_u11_u4_n164 ) , .A1( u2_u11_u4_n165 ) , .ZN( u2_u11_u4_n166 ) );
  NAND3_X1 u2_u11_u4_U96 (.ZN( u2_out11_3 ) , .A3( u2_u11_u4_n166 ) , .A1( u2_u11_u4_n167 ) , .A2( u2_u11_u4_n186 ) );
  NAND3_X1 u2_u11_u4_U97 (.A3( u2_u11_u4_n146 ) , .A2( u2_u11_u4_n147 ) , .A1( u2_u11_u4_n148 ) , .ZN( u2_u11_u4_n149 ) );
  NAND3_X1 u2_u11_u4_U98 (.A3( u2_u11_u4_n143 ) , .A2( u2_u11_u4_n144 ) , .A1( u2_u11_u4_n145 ) , .ZN( u2_u11_u4_n151 ) );
  NAND3_X1 u2_u11_u4_U99 (.A3( u2_u11_u4_n121 ) , .ZN( u2_u11_u4_n122 ) , .A2( u2_u11_u4_n144 ) , .A1( u2_u11_u4_n154 ) );
  INV_X1 u2_u11_u5_U10 (.A( u2_u11_u5_n121 ) , .ZN( u2_u11_u5_n177 ) );
  NOR3_X1 u2_u11_u5_U100 (.A3( u2_u11_u5_n141 ) , .A1( u2_u11_u5_n142 ) , .ZN( u2_u11_u5_n143 ) , .A2( u2_u11_u5_n191 ) );
  NAND4_X1 u2_u11_u5_U101 (.ZN( u2_out11_4 ) , .A4( u2_u11_u5_n112 ) , .A2( u2_u11_u5_n113 ) , .A1( u2_u11_u5_n114 ) , .A3( u2_u11_u5_n195 ) );
  AOI211_X1 u2_u11_u5_U102 (.A( u2_u11_u5_n110 ) , .C1( u2_u11_u5_n111 ) , .ZN( u2_u11_u5_n112 ) , .B( u2_u11_u5_n118 ) , .C2( u2_u11_u5_n177 ) );
  AOI222_X1 u2_u11_u5_U103 (.ZN( u2_u11_u5_n113 ) , .A1( u2_u11_u5_n131 ) , .C1( u2_u11_u5_n148 ) , .B2( u2_u11_u5_n174 ) , .C2( u2_u11_u5_n178 ) , .A2( u2_u11_u5_n179 ) , .B1( u2_u11_u5_n99 ) );
  NAND3_X1 u2_u11_u5_U104 (.A2( u2_u11_u5_n154 ) , .A3( u2_u11_u5_n158 ) , .A1( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n99 ) );
  NOR2_X1 u2_u11_u5_U11 (.ZN( u2_u11_u5_n160 ) , .A2( u2_u11_u5_n173 ) , .A1( u2_u11_u5_n177 ) );
  INV_X1 u2_u11_u5_U12 (.A( u2_u11_u5_n150 ) , .ZN( u2_u11_u5_n174 ) );
  AOI21_X1 u2_u11_u5_U13 (.A( u2_u11_u5_n160 ) , .B2( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n162 ) , .B1( u2_u11_u5_n192 ) );
  INV_X1 u2_u11_u5_U14 (.A( u2_u11_u5_n159 ) , .ZN( u2_u11_u5_n192 ) );
  AOI21_X1 u2_u11_u5_U15 (.A( u2_u11_u5_n156 ) , .B2( u2_u11_u5_n157 ) , .B1( u2_u11_u5_n158 ) , .ZN( u2_u11_u5_n163 ) );
  AOI21_X1 u2_u11_u5_U16 (.B2( u2_u11_u5_n139 ) , .B1( u2_u11_u5_n140 ) , .ZN( u2_u11_u5_n141 ) , .A( u2_u11_u5_n150 ) );
  OAI21_X1 u2_u11_u5_U17 (.A( u2_u11_u5_n133 ) , .B2( u2_u11_u5_n134 ) , .B1( u2_u11_u5_n135 ) , .ZN( u2_u11_u5_n142 ) );
  OAI21_X1 u2_u11_u5_U18 (.ZN( u2_u11_u5_n133 ) , .B2( u2_u11_u5_n147 ) , .A( u2_u11_u5_n173 ) , .B1( u2_u11_u5_n188 ) );
  NAND2_X1 u2_u11_u5_U19 (.A2( u2_u11_u5_n119 ) , .A1( u2_u11_u5_n123 ) , .ZN( u2_u11_u5_n137 ) );
  INV_X1 u2_u11_u5_U20 (.A( u2_u11_u5_n155 ) , .ZN( u2_u11_u5_n194 ) );
  NAND2_X1 u2_u11_u5_U21 (.A1( u2_u11_u5_n121 ) , .ZN( u2_u11_u5_n132 ) , .A2( u2_u11_u5_n172 ) );
  NAND2_X1 u2_u11_u5_U22 (.A2( u2_u11_u5_n122 ) , .ZN( u2_u11_u5_n136 ) , .A1( u2_u11_u5_n154 ) );
  NAND2_X1 u2_u11_u5_U23 (.A2( u2_u11_u5_n119 ) , .A1( u2_u11_u5_n120 ) , .ZN( u2_u11_u5_n159 ) );
  INV_X1 u2_u11_u5_U24 (.A( u2_u11_u5_n156 ) , .ZN( u2_u11_u5_n175 ) );
  INV_X1 u2_u11_u5_U25 (.A( u2_u11_u5_n158 ) , .ZN( u2_u11_u5_n188 ) );
  INV_X1 u2_u11_u5_U26 (.A( u2_u11_u5_n152 ) , .ZN( u2_u11_u5_n179 ) );
  INV_X1 u2_u11_u5_U27 (.A( u2_u11_u5_n140 ) , .ZN( u2_u11_u5_n182 ) );
  INV_X1 u2_u11_u5_U28 (.A( u2_u11_u5_n151 ) , .ZN( u2_u11_u5_n183 ) );
  INV_X1 u2_u11_u5_U29 (.A( u2_u11_u5_n123 ) , .ZN( u2_u11_u5_n185 ) );
  NOR2_X1 u2_u11_u5_U3 (.ZN( u2_u11_u5_n134 ) , .A1( u2_u11_u5_n183 ) , .A2( u2_u11_u5_n190 ) );
  INV_X1 u2_u11_u5_U30 (.A( u2_u11_u5_n161 ) , .ZN( u2_u11_u5_n184 ) );
  INV_X1 u2_u11_u5_U31 (.A( u2_u11_u5_n139 ) , .ZN( u2_u11_u5_n189 ) );
  INV_X1 u2_u11_u5_U32 (.A( u2_u11_u5_n157 ) , .ZN( u2_u11_u5_n190 ) );
  INV_X1 u2_u11_u5_U33 (.A( u2_u11_u5_n120 ) , .ZN( u2_u11_u5_n193 ) );
  NAND2_X1 u2_u11_u5_U34 (.ZN( u2_u11_u5_n111 ) , .A1( u2_u11_u5_n140 ) , .A2( u2_u11_u5_n155 ) );
  NOR2_X1 u2_u11_u5_U35 (.ZN( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n170 ) , .A2( u2_u11_u5_n180 ) );
  INV_X1 u2_u11_u5_U36 (.A( u2_u11_u5_n117 ) , .ZN( u2_u11_u5_n196 ) );
  OAI221_X1 u2_u11_u5_U37 (.A( u2_u11_u5_n116 ) , .ZN( u2_u11_u5_n117 ) , .B2( u2_u11_u5_n119 ) , .C1( u2_u11_u5_n153 ) , .C2( u2_u11_u5_n158 ) , .B1( u2_u11_u5_n172 ) );
  AOI222_X1 u2_u11_u5_U38 (.ZN( u2_u11_u5_n116 ) , .B2( u2_u11_u5_n145 ) , .C1( u2_u11_u5_n148 ) , .A2( u2_u11_u5_n174 ) , .C2( u2_u11_u5_n177 ) , .B1( u2_u11_u5_n187 ) , .A1( u2_u11_u5_n193 ) );
  INV_X1 u2_u11_u5_U39 (.A( u2_u11_u5_n115 ) , .ZN( u2_u11_u5_n187 ) );
  INV_X1 u2_u11_u5_U4 (.A( u2_u11_u5_n138 ) , .ZN( u2_u11_u5_n191 ) );
  AOI22_X1 u2_u11_u5_U40 (.B2( u2_u11_u5_n131 ) , .A2( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n169 ) , .B1( u2_u11_u5_n174 ) , .A1( u2_u11_u5_n185 ) );
  NOR2_X1 u2_u11_u5_U41 (.A1( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n150 ) , .A2( u2_u11_u5_n173 ) );
  AOI21_X1 u2_u11_u5_U42 (.A( u2_u11_u5_n118 ) , .B2( u2_u11_u5_n145 ) , .ZN( u2_u11_u5_n168 ) , .B1( u2_u11_u5_n186 ) );
  INV_X1 u2_u11_u5_U43 (.A( u2_u11_u5_n122 ) , .ZN( u2_u11_u5_n186 ) );
  NOR2_X1 u2_u11_u5_U44 (.A1( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n152 ) , .A2( u2_u11_u5_n176 ) );
  NOR2_X1 u2_u11_u5_U45 (.A1( u2_u11_u5_n115 ) , .ZN( u2_u11_u5_n118 ) , .A2( u2_u11_u5_n153 ) );
  NOR2_X1 u2_u11_u5_U46 (.A2( u2_u11_u5_n145 ) , .ZN( u2_u11_u5_n156 ) , .A1( u2_u11_u5_n174 ) );
  NOR2_X1 u2_u11_u5_U47 (.ZN( u2_u11_u5_n121 ) , .A2( u2_u11_u5_n145 ) , .A1( u2_u11_u5_n176 ) );
  AOI22_X1 u2_u11_u5_U48 (.ZN( u2_u11_u5_n114 ) , .A2( u2_u11_u5_n137 ) , .A1( u2_u11_u5_n145 ) , .B2( u2_u11_u5_n175 ) , .B1( u2_u11_u5_n193 ) );
  OAI211_X1 u2_u11_u5_U49 (.B( u2_u11_u5_n124 ) , .A( u2_u11_u5_n125 ) , .C2( u2_u11_u5_n126 ) , .C1( u2_u11_u5_n127 ) , .ZN( u2_u11_u5_n128 ) );
  OAI21_X1 u2_u11_u5_U5 (.B2( u2_u11_u5_n136 ) , .B1( u2_u11_u5_n137 ) , .ZN( u2_u11_u5_n138 ) , .A( u2_u11_u5_n177 ) );
  OAI21_X1 u2_u11_u5_U50 (.ZN( u2_u11_u5_n124 ) , .A( u2_u11_u5_n177 ) , .B2( u2_u11_u5_n183 ) , .B1( u2_u11_u5_n189 ) );
  NOR3_X1 u2_u11_u5_U51 (.ZN( u2_u11_u5_n127 ) , .A1( u2_u11_u5_n136 ) , .A3( u2_u11_u5_n148 ) , .A2( u2_u11_u5_n182 ) );
  OAI21_X1 u2_u11_u5_U52 (.ZN( u2_u11_u5_n125 ) , .A( u2_u11_u5_n174 ) , .B2( u2_u11_u5_n185 ) , .B1( u2_u11_u5_n190 ) );
  AOI21_X1 u2_u11_u5_U53 (.A( u2_u11_u5_n153 ) , .B2( u2_u11_u5_n154 ) , .B1( u2_u11_u5_n155 ) , .ZN( u2_u11_u5_n164 ) );
  AOI21_X1 u2_u11_u5_U54 (.ZN( u2_u11_u5_n110 ) , .B1( u2_u11_u5_n122 ) , .B2( u2_u11_u5_n139 ) , .A( u2_u11_u5_n153 ) );
  INV_X1 u2_u11_u5_U55 (.A( u2_u11_u5_n153 ) , .ZN( u2_u11_u5_n176 ) );
  INV_X1 u2_u11_u5_U56 (.A( u2_u11_u5_n126 ) , .ZN( u2_u11_u5_n173 ) );
  AND2_X1 u2_u11_u5_U57 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n147 ) );
  AND2_X1 u2_u11_u5_U58 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n148 ) );
  NAND2_X1 u2_u11_u5_U59 (.A1( u2_u11_u5_n105 ) , .A2( u2_u11_u5_n106 ) , .ZN( u2_u11_u5_n158 ) );
  INV_X1 u2_u11_u5_U6 (.A( u2_u11_u5_n135 ) , .ZN( u2_u11_u5_n178 ) );
  NAND2_X1 u2_u11_u5_U60 (.A2( u2_u11_u5_n108 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n139 ) );
  NAND2_X1 u2_u11_u5_U61 (.A1( u2_u11_u5_n106 ) , .A2( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n119 ) );
  NAND2_X1 u2_u11_u5_U62 (.A2( u2_u11_u5_n103 ) , .A1( u2_u11_u5_n105 ) , .ZN( u2_u11_u5_n140 ) );
  NAND2_X1 u2_u11_u5_U63 (.A2( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n105 ) , .ZN( u2_u11_u5_n155 ) );
  NAND2_X1 u2_u11_u5_U64 (.A2( u2_u11_u5_n106 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n122 ) );
  NAND2_X1 u2_u11_u5_U65 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n106 ) , .ZN( u2_u11_u5_n115 ) );
  NAND2_X1 u2_u11_u5_U66 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n103 ) , .ZN( u2_u11_u5_n161 ) );
  NAND2_X1 u2_u11_u5_U67 (.A1( u2_u11_u5_n105 ) , .A2( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n154 ) );
  INV_X1 u2_u11_u5_U68 (.A( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n172 ) );
  NAND2_X1 u2_u11_u5_U69 (.A1( u2_u11_u5_n103 ) , .A2( u2_u11_u5_n108 ) , .ZN( u2_u11_u5_n123 ) );
  OAI22_X1 u2_u11_u5_U7 (.B2( u2_u11_u5_n149 ) , .B1( u2_u11_u5_n150 ) , .A2( u2_u11_u5_n151 ) , .A1( u2_u11_u5_n152 ) , .ZN( u2_u11_u5_n165 ) );
  NAND2_X1 u2_u11_u5_U70 (.A2( u2_u11_u5_n103 ) , .A1( u2_u11_u5_n107 ) , .ZN( u2_u11_u5_n151 ) );
  NAND2_X1 u2_u11_u5_U71 (.A2( u2_u11_u5_n107 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n120 ) );
  NAND2_X1 u2_u11_u5_U72 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n109 ) , .ZN( u2_u11_u5_n157 ) );
  AND2_X1 u2_u11_u5_U73 (.A2( u2_u11_u5_n100 ) , .A1( u2_u11_u5_n104 ) , .ZN( u2_u11_u5_n131 ) );
  INV_X1 u2_u11_u5_U74 (.A( u2_u11_u5_n102 ) , .ZN( u2_u11_u5_n195 ) );
  OAI221_X1 u2_u11_u5_U75 (.A( u2_u11_u5_n101 ) , .ZN( u2_u11_u5_n102 ) , .C2( u2_u11_u5_n115 ) , .C1( u2_u11_u5_n126 ) , .B1( u2_u11_u5_n134 ) , .B2( u2_u11_u5_n160 ) );
  OAI21_X1 u2_u11_u5_U76 (.ZN( u2_u11_u5_n101 ) , .B1( u2_u11_u5_n137 ) , .A( u2_u11_u5_n146 ) , .B2( u2_u11_u5_n147 ) );
  NOR2_X1 u2_u11_u5_U77 (.A2( u2_u11_X_34 ) , .A1( u2_u11_X_35 ) , .ZN( u2_u11_u5_n145 ) );
  NOR2_X1 u2_u11_u5_U78 (.A2( u2_u11_X_34 ) , .ZN( u2_u11_u5_n146 ) , .A1( u2_u11_u5_n171 ) );
  NOR2_X1 u2_u11_u5_U79 (.A2( u2_u11_X_31 ) , .A1( u2_u11_X_32 ) , .ZN( u2_u11_u5_n103 ) );
  NOR3_X1 u2_u11_u5_U8 (.A2( u2_u11_u5_n147 ) , .A1( u2_u11_u5_n148 ) , .ZN( u2_u11_u5_n149 ) , .A3( u2_u11_u5_n194 ) );
  NOR2_X1 u2_u11_u5_U80 (.A2( u2_u11_X_36 ) , .ZN( u2_u11_u5_n105 ) , .A1( u2_u11_u5_n180 ) );
  NOR2_X1 u2_u11_u5_U81 (.A2( u2_u11_X_33 ) , .ZN( u2_u11_u5_n108 ) , .A1( u2_u11_u5_n170 ) );
  NOR2_X1 u2_u11_u5_U82 (.A2( u2_u11_X_33 ) , .A1( u2_u11_X_36 ) , .ZN( u2_u11_u5_n107 ) );
  NOR2_X1 u2_u11_u5_U83 (.A2( u2_u11_X_31 ) , .ZN( u2_u11_u5_n104 ) , .A1( u2_u11_u5_n181 ) );
  NAND2_X1 u2_u11_u5_U84 (.A2( u2_u11_X_34 ) , .A1( u2_u11_X_35 ) , .ZN( u2_u11_u5_n153 ) );
  NAND2_X1 u2_u11_u5_U85 (.A1( u2_u11_X_34 ) , .ZN( u2_u11_u5_n126 ) , .A2( u2_u11_u5_n171 ) );
  AND2_X1 u2_u11_u5_U86 (.A1( u2_u11_X_31 ) , .A2( u2_u11_X_32 ) , .ZN( u2_u11_u5_n106 ) );
  AND2_X1 u2_u11_u5_U87 (.A1( u2_u11_X_31 ) , .ZN( u2_u11_u5_n109 ) , .A2( u2_u11_u5_n181 ) );
  INV_X1 u2_u11_u5_U88 (.A( u2_u11_X_33 ) , .ZN( u2_u11_u5_n180 ) );
  INV_X1 u2_u11_u5_U89 (.A( u2_u11_X_35 ) , .ZN( u2_u11_u5_n171 ) );
  NOR2_X1 u2_u11_u5_U9 (.ZN( u2_u11_u5_n135 ) , .A1( u2_u11_u5_n173 ) , .A2( u2_u11_u5_n176 ) );
  INV_X1 u2_u11_u5_U90 (.A( u2_u11_X_36 ) , .ZN( u2_u11_u5_n170 ) );
  INV_X1 u2_u11_u5_U91 (.A( u2_u11_X_32 ) , .ZN( u2_u11_u5_n181 ) );
  NAND4_X1 u2_u11_u5_U92 (.ZN( u2_out11_29 ) , .A4( u2_u11_u5_n129 ) , .A3( u2_u11_u5_n130 ) , .A2( u2_u11_u5_n168 ) , .A1( u2_u11_u5_n196 ) );
  AOI221_X1 u2_u11_u5_U93 (.A( u2_u11_u5_n128 ) , .ZN( u2_u11_u5_n129 ) , .C2( u2_u11_u5_n132 ) , .B2( u2_u11_u5_n159 ) , .B1( u2_u11_u5_n176 ) , .C1( u2_u11_u5_n184 ) );
  AOI222_X1 u2_u11_u5_U94 (.ZN( u2_u11_u5_n130 ) , .A2( u2_u11_u5_n146 ) , .B1( u2_u11_u5_n147 ) , .C2( u2_u11_u5_n175 ) , .B2( u2_u11_u5_n179 ) , .A1( u2_u11_u5_n188 ) , .C1( u2_u11_u5_n194 ) );
  NAND4_X1 u2_u11_u5_U95 (.ZN( u2_out11_19 ) , .A4( u2_u11_u5_n166 ) , .A3( u2_u11_u5_n167 ) , .A2( u2_u11_u5_n168 ) , .A1( u2_u11_u5_n169 ) );
  AOI22_X1 u2_u11_u5_U96 (.B2( u2_u11_u5_n145 ) , .A2( u2_u11_u5_n146 ) , .ZN( u2_u11_u5_n167 ) , .B1( u2_u11_u5_n182 ) , .A1( u2_u11_u5_n189 ) );
  NOR4_X1 u2_u11_u5_U97 (.A4( u2_u11_u5_n162 ) , .A3( u2_u11_u5_n163 ) , .A2( u2_u11_u5_n164 ) , .A1( u2_u11_u5_n165 ) , .ZN( u2_u11_u5_n166 ) );
  NAND4_X1 u2_u11_u5_U98 (.ZN( u2_out11_11 ) , .A4( u2_u11_u5_n143 ) , .A3( u2_u11_u5_n144 ) , .A2( u2_u11_u5_n169 ) , .A1( u2_u11_u5_n196 ) );
  AOI22_X1 u2_u11_u5_U99 (.A2( u2_u11_u5_n132 ) , .ZN( u2_u11_u5_n144 ) , .B2( u2_u11_u5_n145 ) , .B1( u2_u11_u5_n184 ) , .A1( u2_u11_u5_n194 ) );
  OAI21_X1 u2_u11_u6_U10 (.A( u2_u11_u6_n159 ) , .B1( u2_u11_u6_n169 ) , .B2( u2_u11_u6_n173 ) , .ZN( u2_u11_u6_n90 ) );
  INV_X1 u2_u11_u6_U11 (.ZN( u2_u11_u6_n172 ) , .A( u2_u11_u6_n88 ) );
  AOI22_X1 u2_u11_u6_U12 (.A2( u2_u11_u6_n151 ) , .B2( u2_u11_u6_n161 ) , .A1( u2_u11_u6_n167 ) , .B1( u2_u11_u6_n170 ) , .ZN( u2_u11_u6_n89 ) );
  AOI21_X1 u2_u11_u6_U13 (.ZN( u2_u11_u6_n106 ) , .A( u2_u11_u6_n142 ) , .B2( u2_u11_u6_n159 ) , .B1( u2_u11_u6_n164 ) );
  INV_X1 u2_u11_u6_U14 (.A( u2_u11_u6_n155 ) , .ZN( u2_u11_u6_n161 ) );
  INV_X1 u2_u11_u6_U15 (.A( u2_u11_u6_n128 ) , .ZN( u2_u11_u6_n164 ) );
  NAND2_X1 u2_u11_u6_U16 (.ZN( u2_u11_u6_n110 ) , .A1( u2_u11_u6_n122 ) , .A2( u2_u11_u6_n129 ) );
  NAND2_X1 u2_u11_u6_U17 (.ZN( u2_u11_u6_n124 ) , .A2( u2_u11_u6_n146 ) , .A1( u2_u11_u6_n148 ) );
  INV_X1 u2_u11_u6_U18 (.A( u2_u11_u6_n132 ) , .ZN( u2_u11_u6_n171 ) );
  AND2_X1 u2_u11_u6_U19 (.A1( u2_u11_u6_n100 ) , .ZN( u2_u11_u6_n130 ) , .A2( u2_u11_u6_n147 ) );
  INV_X1 u2_u11_u6_U20 (.A( u2_u11_u6_n127 ) , .ZN( u2_u11_u6_n173 ) );
  INV_X1 u2_u11_u6_U21 (.A( u2_u11_u6_n121 ) , .ZN( u2_u11_u6_n167 ) );
  INV_X1 u2_u11_u6_U22 (.A( u2_u11_u6_n100 ) , .ZN( u2_u11_u6_n169 ) );
  INV_X1 u2_u11_u6_U23 (.A( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n170 ) );
  INV_X1 u2_u11_u6_U24 (.A( u2_u11_u6_n113 ) , .ZN( u2_u11_u6_n168 ) );
  AND2_X1 u2_u11_u6_U25 (.A1( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n119 ) , .ZN( u2_u11_u6_n133 ) );
  AND2_X1 u2_u11_u6_U26 (.A2( u2_u11_u6_n121 ) , .A1( u2_u11_u6_n122 ) , .ZN( u2_u11_u6_n131 ) );
  AND3_X1 u2_u11_u6_U27 (.ZN( u2_u11_u6_n120 ) , .A2( u2_u11_u6_n127 ) , .A1( u2_u11_u6_n132 ) , .A3( u2_u11_u6_n145 ) );
  INV_X1 u2_u11_u6_U28 (.A( u2_u11_u6_n146 ) , .ZN( u2_u11_u6_n163 ) );
  AOI222_X1 u2_u11_u6_U29 (.ZN( u2_u11_u6_n114 ) , .A1( u2_u11_u6_n118 ) , .A2( u2_u11_u6_n126 ) , .B2( u2_u11_u6_n151 ) , .C2( u2_u11_u6_n159 ) , .C1( u2_u11_u6_n168 ) , .B1( u2_u11_u6_n169 ) );
  INV_X1 u2_u11_u6_U3 (.A( u2_u11_u6_n110 ) , .ZN( u2_u11_u6_n166 ) );
  NOR2_X1 u2_u11_u6_U30 (.A1( u2_u11_u6_n162 ) , .A2( u2_u11_u6_n165 ) , .ZN( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U31 (.A1( u2_u11_u6_n144 ) , .ZN( u2_u11_u6_n151 ) , .A2( u2_u11_u6_n158 ) );
  NAND2_X1 u2_u11_u6_U32 (.ZN( u2_u11_u6_n132 ) , .A1( u2_u11_u6_n91 ) , .A2( u2_u11_u6_n97 ) );
  AOI22_X1 u2_u11_u6_U33 (.B2( u2_u11_u6_n110 ) , .B1( u2_u11_u6_n111 ) , .A1( u2_u11_u6_n112 ) , .ZN( u2_u11_u6_n115 ) , .A2( u2_u11_u6_n161 ) );
  NAND4_X1 u2_u11_u6_U34 (.A3( u2_u11_u6_n109 ) , .ZN( u2_u11_u6_n112 ) , .A4( u2_u11_u6_n132 ) , .A2( u2_u11_u6_n147 ) , .A1( u2_u11_u6_n166 ) );
  NOR2_X1 u2_u11_u6_U35 (.ZN( u2_u11_u6_n109 ) , .A1( u2_u11_u6_n170 ) , .A2( u2_u11_u6_n173 ) );
  NOR2_X1 u2_u11_u6_U36 (.A2( u2_u11_u6_n126 ) , .ZN( u2_u11_u6_n155 ) , .A1( u2_u11_u6_n160 ) );
  NAND2_X1 u2_u11_u6_U37 (.ZN( u2_u11_u6_n146 ) , .A2( u2_u11_u6_n94 ) , .A1( u2_u11_u6_n99 ) );
  AOI21_X1 u2_u11_u6_U38 (.A( u2_u11_u6_n144 ) , .B2( u2_u11_u6_n145 ) , .B1( u2_u11_u6_n146 ) , .ZN( u2_u11_u6_n150 ) );
  AOI211_X1 u2_u11_u6_U39 (.B( u2_u11_u6_n134 ) , .A( u2_u11_u6_n135 ) , .C1( u2_u11_u6_n136 ) , .ZN( u2_u11_u6_n137 ) , .C2( u2_u11_u6_n151 ) );
  INV_X1 u2_u11_u6_U4 (.A( u2_u11_u6_n142 ) , .ZN( u2_u11_u6_n174 ) );
  NAND4_X1 u2_u11_u6_U40 (.A4( u2_u11_u6_n127 ) , .A3( u2_u11_u6_n128 ) , .A2( u2_u11_u6_n129 ) , .A1( u2_u11_u6_n130 ) , .ZN( u2_u11_u6_n136 ) );
  AOI21_X1 u2_u11_u6_U41 (.B2( u2_u11_u6_n132 ) , .B1( u2_u11_u6_n133 ) , .ZN( u2_u11_u6_n134 ) , .A( u2_u11_u6_n158 ) );
  AOI21_X1 u2_u11_u6_U42 (.B1( u2_u11_u6_n131 ) , .ZN( u2_u11_u6_n135 ) , .A( u2_u11_u6_n144 ) , .B2( u2_u11_u6_n146 ) );
  INV_X1 u2_u11_u6_U43 (.A( u2_u11_u6_n111 ) , .ZN( u2_u11_u6_n158 ) );
  NAND2_X1 u2_u11_u6_U44 (.ZN( u2_u11_u6_n127 ) , .A1( u2_u11_u6_n91 ) , .A2( u2_u11_u6_n92 ) );
  NAND2_X1 u2_u11_u6_U45 (.ZN( u2_u11_u6_n129 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n96 ) );
  INV_X1 u2_u11_u6_U46 (.A( u2_u11_u6_n144 ) , .ZN( u2_u11_u6_n159 ) );
  NAND2_X1 u2_u11_u6_U47 (.ZN( u2_u11_u6_n145 ) , .A2( u2_u11_u6_n97 ) , .A1( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U48 (.ZN( u2_u11_u6_n148 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n94 ) );
  NAND2_X1 u2_u11_u6_U49 (.ZN( u2_u11_u6_n108 ) , .A2( u2_u11_u6_n139 ) , .A1( u2_u11_u6_n144 ) );
  NAND2_X1 u2_u11_u6_U5 (.A2( u2_u11_u6_n143 ) , .ZN( u2_u11_u6_n152 ) , .A1( u2_u11_u6_n166 ) );
  NAND2_X1 u2_u11_u6_U50 (.ZN( u2_u11_u6_n121 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n97 ) );
  NAND2_X1 u2_u11_u6_U51 (.ZN( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n95 ) );
  AND2_X1 u2_u11_u6_U52 (.ZN( u2_u11_u6_n118 ) , .A2( u2_u11_u6_n91 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U53 (.ZN( u2_u11_u6_n147 ) , .A2( u2_u11_u6_n98 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U54 (.ZN( u2_u11_u6_n128 ) , .A1( u2_u11_u6_n94 ) , .A2( u2_u11_u6_n96 ) );
  NAND2_X1 u2_u11_u6_U55 (.ZN( u2_u11_u6_n119 ) , .A2( u2_u11_u6_n95 ) , .A1( u2_u11_u6_n99 ) );
  NAND2_X1 u2_u11_u6_U56 (.ZN( u2_u11_u6_n123 ) , .A2( u2_u11_u6_n91 ) , .A1( u2_u11_u6_n96 ) );
  NAND2_X1 u2_u11_u6_U57 (.ZN( u2_u11_u6_n100 ) , .A2( u2_u11_u6_n92 ) , .A1( u2_u11_u6_n98 ) );
  NAND2_X1 u2_u11_u6_U58 (.ZN( u2_u11_u6_n122 ) , .A1( u2_u11_u6_n94 ) , .A2( u2_u11_u6_n97 ) );
  INV_X1 u2_u11_u6_U59 (.A( u2_u11_u6_n139 ) , .ZN( u2_u11_u6_n160 ) );
  AOI22_X1 u2_u11_u6_U6 (.B2( u2_u11_u6_n101 ) , .A1( u2_u11_u6_n102 ) , .ZN( u2_u11_u6_n103 ) , .B1( u2_u11_u6_n160 ) , .A2( u2_u11_u6_n161 ) );
  NAND2_X1 u2_u11_u6_U60 (.ZN( u2_u11_u6_n113 ) , .A1( u2_u11_u6_n96 ) , .A2( u2_u11_u6_n98 ) );
  NOR2_X1 u2_u11_u6_U61 (.A2( u2_u11_X_40 ) , .A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n126 ) );
  NOR2_X1 u2_u11_u6_U62 (.A2( u2_u11_X_39 ) , .A1( u2_u11_X_42 ) , .ZN( u2_u11_u6_n92 ) );
  NOR2_X1 u2_u11_u6_U63 (.A2( u2_u11_X_39 ) , .A1( u2_u11_u6_n156 ) , .ZN( u2_u11_u6_n97 ) );
  NOR2_X1 u2_u11_u6_U64 (.A2( u2_u11_X_38 ) , .A1( u2_u11_u6_n165 ) , .ZN( u2_u11_u6_n95 ) );
  NOR2_X1 u2_u11_u6_U65 (.A2( u2_u11_X_41 ) , .ZN( u2_u11_u6_n111 ) , .A1( u2_u11_u6_n157 ) );
  NOR2_X1 u2_u11_u6_U66 (.A2( u2_u11_X_37 ) , .A1( u2_u11_u6_n162 ) , .ZN( u2_u11_u6_n94 ) );
  NOR2_X1 u2_u11_u6_U67 (.A2( u2_u11_X_37 ) , .A1( u2_u11_X_38 ) , .ZN( u2_u11_u6_n91 ) );
  NAND2_X1 u2_u11_u6_U68 (.A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n144 ) , .A2( u2_u11_u6_n157 ) );
  NAND2_X1 u2_u11_u6_U69 (.A2( u2_u11_X_40 ) , .A1( u2_u11_X_41 ) , .ZN( u2_u11_u6_n139 ) );
  NOR2_X1 u2_u11_u6_U7 (.A1( u2_u11_u6_n118 ) , .ZN( u2_u11_u6_n143 ) , .A2( u2_u11_u6_n168 ) );
  AND2_X1 u2_u11_u6_U70 (.A1( u2_u11_X_39 ) , .A2( u2_u11_u6_n156 ) , .ZN( u2_u11_u6_n96 ) );
  AND2_X1 u2_u11_u6_U71 (.A1( u2_u11_X_39 ) , .A2( u2_u11_X_42 ) , .ZN( u2_u11_u6_n99 ) );
  INV_X1 u2_u11_u6_U72 (.A( u2_u11_X_40 ) , .ZN( u2_u11_u6_n157 ) );
  INV_X1 u2_u11_u6_U73 (.A( u2_u11_X_37 ) , .ZN( u2_u11_u6_n165 ) );
  INV_X1 u2_u11_u6_U74 (.A( u2_u11_X_38 ) , .ZN( u2_u11_u6_n162 ) );
  INV_X1 u2_u11_u6_U75 (.A( u2_u11_X_42 ) , .ZN( u2_u11_u6_n156 ) );
  NAND4_X1 u2_u11_u6_U76 (.ZN( u2_out11_32 ) , .A4( u2_u11_u6_n103 ) , .A3( u2_u11_u6_n104 ) , .A2( u2_u11_u6_n105 ) , .A1( u2_u11_u6_n106 ) );
  AOI22_X1 u2_u11_u6_U77 (.ZN( u2_u11_u6_n105 ) , .A2( u2_u11_u6_n108 ) , .A1( u2_u11_u6_n118 ) , .B2( u2_u11_u6_n126 ) , .B1( u2_u11_u6_n171 ) );
  AOI22_X1 u2_u11_u6_U78 (.ZN( u2_u11_u6_n104 ) , .A1( u2_u11_u6_n111 ) , .B1( u2_u11_u6_n124 ) , .B2( u2_u11_u6_n151 ) , .A2( u2_u11_u6_n93 ) );
  NAND4_X1 u2_u11_u6_U79 (.ZN( u2_out11_12 ) , .A4( u2_u11_u6_n114 ) , .A3( u2_u11_u6_n115 ) , .A2( u2_u11_u6_n116 ) , .A1( u2_u11_u6_n117 ) );
  AOI21_X1 u2_u11_u6_U8 (.B1( u2_u11_u6_n107 ) , .B2( u2_u11_u6_n132 ) , .A( u2_u11_u6_n158 ) , .ZN( u2_u11_u6_n88 ) );
  OAI22_X1 u2_u11_u6_U80 (.B2( u2_u11_u6_n111 ) , .ZN( u2_u11_u6_n116 ) , .B1( u2_u11_u6_n126 ) , .A2( u2_u11_u6_n164 ) , .A1( u2_u11_u6_n167 ) );
  OAI21_X1 u2_u11_u6_U81 (.A( u2_u11_u6_n108 ) , .ZN( u2_u11_u6_n117 ) , .B2( u2_u11_u6_n141 ) , .B1( u2_u11_u6_n163 ) );
  OAI211_X1 u2_u11_u6_U82 (.ZN( u2_out11_7 ) , .B( u2_u11_u6_n153 ) , .C2( u2_u11_u6_n154 ) , .C1( u2_u11_u6_n155 ) , .A( u2_u11_u6_n174 ) );
  NOR3_X1 u2_u11_u6_U83 (.A1( u2_u11_u6_n141 ) , .ZN( u2_u11_u6_n154 ) , .A3( u2_u11_u6_n164 ) , .A2( u2_u11_u6_n171 ) );
  AOI211_X1 u2_u11_u6_U84 (.B( u2_u11_u6_n149 ) , .A( u2_u11_u6_n150 ) , .C2( u2_u11_u6_n151 ) , .C1( u2_u11_u6_n152 ) , .ZN( u2_u11_u6_n153 ) );
  OAI211_X1 u2_u11_u6_U85 (.ZN( u2_out11_22 ) , .B( u2_u11_u6_n137 ) , .A( u2_u11_u6_n138 ) , .C2( u2_u11_u6_n139 ) , .C1( u2_u11_u6_n140 ) );
  AOI22_X1 u2_u11_u6_U86 (.B1( u2_u11_u6_n124 ) , .A2( u2_u11_u6_n125 ) , .A1( u2_u11_u6_n126 ) , .ZN( u2_u11_u6_n138 ) , .B2( u2_u11_u6_n161 ) );
  AND4_X1 u2_u11_u6_U87 (.A3( u2_u11_u6_n119 ) , .A1( u2_u11_u6_n120 ) , .A4( u2_u11_u6_n129 ) , .ZN( u2_u11_u6_n140 ) , .A2( u2_u11_u6_n143 ) );
  NAND3_X1 u2_u11_u6_U88 (.A2( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n125 ) , .A1( u2_u11_u6_n130 ) , .A3( u2_u11_u6_n131 ) );
  NAND3_X1 u2_u11_u6_U89 (.A3( u2_u11_u6_n133 ) , .ZN( u2_u11_u6_n141 ) , .A1( u2_u11_u6_n145 ) , .A2( u2_u11_u6_n148 ) );
  AOI21_X1 u2_u11_u6_U9 (.B2( u2_u11_u6_n147 ) , .B1( u2_u11_u6_n148 ) , .ZN( u2_u11_u6_n149 ) , .A( u2_u11_u6_n158 ) );
  NAND3_X1 u2_u11_u6_U90 (.ZN( u2_u11_u6_n101 ) , .A3( u2_u11_u6_n107 ) , .A2( u2_u11_u6_n121 ) , .A1( u2_u11_u6_n127 ) );
  NAND3_X1 u2_u11_u6_U91 (.ZN( u2_u11_u6_n102 ) , .A3( u2_u11_u6_n130 ) , .A2( u2_u11_u6_n145 ) , .A1( u2_u11_u6_n166 ) );
  NAND3_X1 u2_u11_u6_U92 (.A3( u2_u11_u6_n113 ) , .A1( u2_u11_u6_n119 ) , .A2( u2_u11_u6_n123 ) , .ZN( u2_u11_u6_n93 ) );
  NAND3_X1 u2_u11_u6_U93 (.ZN( u2_u11_u6_n142 ) , .A2( u2_u11_u6_n172 ) , .A3( u2_u11_u6_n89 ) , .A1( u2_u11_u6_n90 ) );
  AND3_X1 u2_u11_u7_U10 (.A3( u2_u11_u7_n110 ) , .A2( u2_u11_u7_n127 ) , .A1( u2_u11_u7_n132 ) , .ZN( u2_u11_u7_n92 ) );
  OAI21_X1 u2_u11_u7_U11 (.A( u2_u11_u7_n161 ) , .B1( u2_u11_u7_n168 ) , .B2( u2_u11_u7_n173 ) , .ZN( u2_u11_u7_n91 ) );
  AOI211_X1 u2_u11_u7_U12 (.A( u2_u11_u7_n117 ) , .ZN( u2_u11_u7_n118 ) , .C2( u2_u11_u7_n126 ) , .C1( u2_u11_u7_n177 ) , .B( u2_u11_u7_n180 ) );
  OAI22_X1 u2_u11_u7_U13 (.B1( u2_u11_u7_n115 ) , .ZN( u2_u11_u7_n117 ) , .A2( u2_u11_u7_n133 ) , .A1( u2_u11_u7_n137 ) , .B2( u2_u11_u7_n162 ) );
  INV_X1 u2_u11_u7_U14 (.A( u2_u11_u7_n116 ) , .ZN( u2_u11_u7_n180 ) );
  NOR3_X1 u2_u11_u7_U15 (.ZN( u2_u11_u7_n115 ) , .A3( u2_u11_u7_n145 ) , .A2( u2_u11_u7_n168 ) , .A1( u2_u11_u7_n169 ) );
  OAI211_X1 u2_u11_u7_U16 (.B( u2_u11_u7_n122 ) , .A( u2_u11_u7_n123 ) , .C2( u2_u11_u7_n124 ) , .ZN( u2_u11_u7_n154 ) , .C1( u2_u11_u7_n162 ) );
  AOI222_X1 u2_u11_u7_U17 (.ZN( u2_u11_u7_n122 ) , .C2( u2_u11_u7_n126 ) , .C1( u2_u11_u7_n145 ) , .B1( u2_u11_u7_n161 ) , .A2( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n170 ) , .A1( u2_u11_u7_n176 ) );
  INV_X1 u2_u11_u7_U18 (.A( u2_u11_u7_n133 ) , .ZN( u2_u11_u7_n176 ) );
  NOR3_X1 u2_u11_u7_U19 (.A2( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n135 ) , .ZN( u2_u11_u7_n136 ) , .A3( u2_u11_u7_n171 ) );
  NOR2_X1 u2_u11_u7_U20 (.A1( u2_u11_u7_n130 ) , .A2( u2_u11_u7_n134 ) , .ZN( u2_u11_u7_n153 ) );
  INV_X1 u2_u11_u7_U21 (.A( u2_u11_u7_n101 ) , .ZN( u2_u11_u7_n165 ) );
  NOR2_X1 u2_u11_u7_U22 (.ZN( u2_u11_u7_n111 ) , .A2( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n169 ) );
  AOI21_X1 u2_u11_u7_U23 (.ZN( u2_u11_u7_n104 ) , .B2( u2_u11_u7_n112 ) , .B1( u2_u11_u7_n127 ) , .A( u2_u11_u7_n164 ) );
  AOI21_X1 u2_u11_u7_U24 (.ZN( u2_u11_u7_n106 ) , .B1( u2_u11_u7_n133 ) , .B2( u2_u11_u7_n146 ) , .A( u2_u11_u7_n162 ) );
  AOI21_X1 u2_u11_u7_U25 (.A( u2_u11_u7_n101 ) , .ZN( u2_u11_u7_n107 ) , .B2( u2_u11_u7_n128 ) , .B1( u2_u11_u7_n175 ) );
  INV_X1 u2_u11_u7_U26 (.A( u2_u11_u7_n138 ) , .ZN( u2_u11_u7_n171 ) );
  INV_X1 u2_u11_u7_U27 (.A( u2_u11_u7_n131 ) , .ZN( u2_u11_u7_n177 ) );
  INV_X1 u2_u11_u7_U28 (.A( u2_u11_u7_n110 ) , .ZN( u2_u11_u7_n174 ) );
  NAND2_X1 u2_u11_u7_U29 (.A1( u2_u11_u7_n129 ) , .A2( u2_u11_u7_n132 ) , .ZN( u2_u11_u7_n149 ) );
  OAI21_X1 u2_u11_u7_U3 (.ZN( u2_u11_u7_n159 ) , .A( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n171 ) , .B1( u2_u11_u7_n174 ) );
  NAND2_X1 u2_u11_u7_U30 (.A1( u2_u11_u7_n113 ) , .A2( u2_u11_u7_n124 ) , .ZN( u2_u11_u7_n130 ) );
  INV_X1 u2_u11_u7_U31 (.A( u2_u11_u7_n112 ) , .ZN( u2_u11_u7_n173 ) );
  INV_X1 u2_u11_u7_U32 (.A( u2_u11_u7_n128 ) , .ZN( u2_u11_u7_n168 ) );
  INV_X1 u2_u11_u7_U33 (.A( u2_u11_u7_n148 ) , .ZN( u2_u11_u7_n169 ) );
  INV_X1 u2_u11_u7_U34 (.A( u2_u11_u7_n127 ) , .ZN( u2_u11_u7_n179 ) );
  NOR2_X1 u2_u11_u7_U35 (.ZN( u2_u11_u7_n101 ) , .A2( u2_u11_u7_n150 ) , .A1( u2_u11_u7_n156 ) );
  AOI211_X1 u2_u11_u7_U36 (.B( u2_u11_u7_n154 ) , .A( u2_u11_u7_n155 ) , .C1( u2_u11_u7_n156 ) , .ZN( u2_u11_u7_n157 ) , .C2( u2_u11_u7_n172 ) );
  INV_X1 u2_u11_u7_U37 (.A( u2_u11_u7_n153 ) , .ZN( u2_u11_u7_n172 ) );
  AOI211_X1 u2_u11_u7_U38 (.B( u2_u11_u7_n139 ) , .A( u2_u11_u7_n140 ) , .C2( u2_u11_u7_n141 ) , .ZN( u2_u11_u7_n142 ) , .C1( u2_u11_u7_n156 ) );
  AOI21_X1 u2_u11_u7_U39 (.A( u2_u11_u7_n137 ) , .B1( u2_u11_u7_n138 ) , .ZN( u2_u11_u7_n139 ) , .B2( u2_u11_u7_n146 ) );
  INV_X1 u2_u11_u7_U4 (.A( u2_u11_u7_n111 ) , .ZN( u2_u11_u7_n170 ) );
  NAND4_X1 u2_u11_u7_U40 (.A3( u2_u11_u7_n127 ) , .A2( u2_u11_u7_n128 ) , .A1( u2_u11_u7_n129 ) , .ZN( u2_u11_u7_n141 ) , .A4( u2_u11_u7_n147 ) );
  OAI22_X1 u2_u11_u7_U41 (.B1( u2_u11_u7_n136 ) , .ZN( u2_u11_u7_n140 ) , .A1( u2_u11_u7_n153 ) , .B2( u2_u11_u7_n162 ) , .A2( u2_u11_u7_n164 ) );
  AOI21_X1 u2_u11_u7_U42 (.ZN( u2_u11_u7_n123 ) , .B1( u2_u11_u7_n165 ) , .B2( u2_u11_u7_n177 ) , .A( u2_u11_u7_n97 ) );
  AOI21_X1 u2_u11_u7_U43 (.B2( u2_u11_u7_n113 ) , .B1( u2_u11_u7_n124 ) , .A( u2_u11_u7_n125 ) , .ZN( u2_u11_u7_n97 ) );
  INV_X1 u2_u11_u7_U44 (.A( u2_u11_u7_n125 ) , .ZN( u2_u11_u7_n161 ) );
  INV_X1 u2_u11_u7_U45 (.A( u2_u11_u7_n152 ) , .ZN( u2_u11_u7_n162 ) );
  AOI22_X1 u2_u11_u7_U46 (.A2( u2_u11_u7_n114 ) , .ZN( u2_u11_u7_n119 ) , .B1( u2_u11_u7_n130 ) , .A1( u2_u11_u7_n156 ) , .B2( u2_u11_u7_n165 ) );
  NAND2_X1 u2_u11_u7_U47 (.A2( u2_u11_u7_n112 ) , .ZN( u2_u11_u7_n114 ) , .A1( u2_u11_u7_n175 ) );
  AND2_X1 u2_u11_u7_U48 (.ZN( u2_u11_u7_n145 ) , .A2( u2_u11_u7_n98 ) , .A1( u2_u11_u7_n99 ) );
  NOR2_X1 u2_u11_u7_U49 (.ZN( u2_u11_u7_n137 ) , .A1( u2_u11_u7_n150 ) , .A2( u2_u11_u7_n161 ) );
  INV_X1 u2_u11_u7_U5 (.A( u2_u11_u7_n149 ) , .ZN( u2_u11_u7_n175 ) );
  AOI21_X1 u2_u11_u7_U50 (.ZN( u2_u11_u7_n105 ) , .B2( u2_u11_u7_n110 ) , .A( u2_u11_u7_n125 ) , .B1( u2_u11_u7_n147 ) );
  NAND2_X1 u2_u11_u7_U51 (.ZN( u2_u11_u7_n146 ) , .A1( u2_u11_u7_n95 ) , .A2( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U52 (.A2( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n147 ) , .A1( u2_u11_u7_n93 ) );
  NAND2_X1 u2_u11_u7_U53 (.A1( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n127 ) , .A2( u2_u11_u7_n99 ) );
  OR2_X1 u2_u11_u7_U54 (.ZN( u2_u11_u7_n126 ) , .A2( u2_u11_u7_n152 ) , .A1( u2_u11_u7_n156 ) );
  NAND2_X1 u2_u11_u7_U55 (.A2( u2_u11_u7_n102 ) , .A1( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n133 ) );
  NAND2_X1 u2_u11_u7_U56 (.ZN( u2_u11_u7_n112 ) , .A2( u2_u11_u7_n96 ) , .A1( u2_u11_u7_n99 ) );
  NAND2_X1 u2_u11_u7_U57 (.A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n128 ) , .A1( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U58 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n113 ) , .A2( u2_u11_u7_n93 ) );
  NAND2_X1 u2_u11_u7_U59 (.A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n124 ) , .A1( u2_u11_u7_n96 ) );
  INV_X1 u2_u11_u7_U6 (.A( u2_u11_u7_n154 ) , .ZN( u2_u11_u7_n178 ) );
  NAND2_X1 u2_u11_u7_U60 (.ZN( u2_u11_u7_n110 ) , .A1( u2_u11_u7_n95 ) , .A2( u2_u11_u7_n96 ) );
  INV_X1 u2_u11_u7_U61 (.A( u2_u11_u7_n150 ) , .ZN( u2_u11_u7_n164 ) );
  AND2_X1 u2_u11_u7_U62 (.ZN( u2_u11_u7_n134 ) , .A1( u2_u11_u7_n93 ) , .A2( u2_u11_u7_n98 ) );
  NAND2_X1 u2_u11_u7_U63 (.A1( u2_u11_u7_n100 ) , .A2( u2_u11_u7_n102 ) , .ZN( u2_u11_u7_n129 ) );
  NAND2_X1 u2_u11_u7_U64 (.A2( u2_u11_u7_n103 ) , .ZN( u2_u11_u7_n131 ) , .A1( u2_u11_u7_n95 ) );
  NAND2_X1 u2_u11_u7_U65 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n138 ) , .A2( u2_u11_u7_n99 ) );
  NAND2_X1 u2_u11_u7_U66 (.ZN( u2_u11_u7_n132 ) , .A1( u2_u11_u7_n93 ) , .A2( u2_u11_u7_n96 ) );
  NAND2_X1 u2_u11_u7_U67 (.A1( u2_u11_u7_n100 ) , .ZN( u2_u11_u7_n148 ) , .A2( u2_u11_u7_n95 ) );
  NOR2_X1 u2_u11_u7_U68 (.A2( u2_u11_X_47 ) , .ZN( u2_u11_u7_n150 ) , .A1( u2_u11_u7_n163 ) );
  NOR2_X1 u2_u11_u7_U69 (.A2( u2_u11_X_43 ) , .A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n103 ) );
  AOI211_X1 u2_u11_u7_U7 (.ZN( u2_u11_u7_n116 ) , .A( u2_u11_u7_n155 ) , .C1( u2_u11_u7_n161 ) , .C2( u2_u11_u7_n171 ) , .B( u2_u11_u7_n94 ) );
  NOR2_X1 u2_u11_u7_U70 (.A2( u2_u11_X_48 ) , .A1( u2_u11_u7_n166 ) , .ZN( u2_u11_u7_n95 ) );
  NOR2_X1 u2_u11_u7_U71 (.A2( u2_u11_X_45 ) , .A1( u2_u11_X_48 ) , .ZN( u2_u11_u7_n99 ) );
  NOR2_X1 u2_u11_u7_U72 (.A2( u2_u11_X_44 ) , .A1( u2_u11_u7_n167 ) , .ZN( u2_u11_u7_n98 ) );
  NOR2_X1 u2_u11_u7_U73 (.A2( u2_u11_X_46 ) , .A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n152 ) );
  AND2_X1 u2_u11_u7_U74 (.A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n156 ) , .A2( u2_u11_u7_n163 ) );
  NAND2_X1 u2_u11_u7_U75 (.A2( u2_u11_X_46 ) , .A1( u2_u11_X_47 ) , .ZN( u2_u11_u7_n125 ) );
  AND2_X1 u2_u11_u7_U76 (.A2( u2_u11_X_45 ) , .A1( u2_u11_X_48 ) , .ZN( u2_u11_u7_n102 ) );
  AND2_X1 u2_u11_u7_U77 (.A2( u2_u11_X_43 ) , .A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n96 ) );
  AND2_X1 u2_u11_u7_U78 (.A1( u2_u11_X_44 ) , .ZN( u2_u11_u7_n100 ) , .A2( u2_u11_u7_n167 ) );
  AND2_X1 u2_u11_u7_U79 (.A1( u2_u11_X_48 ) , .A2( u2_u11_u7_n166 ) , .ZN( u2_u11_u7_n93 ) );
  OAI222_X1 u2_u11_u7_U8 (.C2( u2_u11_u7_n101 ) , .B2( u2_u11_u7_n111 ) , .A1( u2_u11_u7_n113 ) , .C1( u2_u11_u7_n146 ) , .A2( u2_u11_u7_n162 ) , .B1( u2_u11_u7_n164 ) , .ZN( u2_u11_u7_n94 ) );
  INV_X1 u2_u11_u7_U80 (.A( u2_u11_X_46 ) , .ZN( u2_u11_u7_n163 ) );
  INV_X1 u2_u11_u7_U81 (.A( u2_u11_X_43 ) , .ZN( u2_u11_u7_n167 ) );
  INV_X1 u2_u11_u7_U82 (.A( u2_u11_X_45 ) , .ZN( u2_u11_u7_n166 ) );
  NAND4_X1 u2_u11_u7_U83 (.ZN( u2_out11_27 ) , .A4( u2_u11_u7_n118 ) , .A3( u2_u11_u7_n119 ) , .A2( u2_u11_u7_n120 ) , .A1( u2_u11_u7_n121 ) );
  OAI21_X1 u2_u11_u7_U84 (.ZN( u2_u11_u7_n121 ) , .B2( u2_u11_u7_n145 ) , .A( u2_u11_u7_n150 ) , .B1( u2_u11_u7_n174 ) );
  OAI21_X1 u2_u11_u7_U85 (.ZN( u2_u11_u7_n120 ) , .A( u2_u11_u7_n161 ) , .B2( u2_u11_u7_n170 ) , .B1( u2_u11_u7_n179 ) );
  NAND4_X1 u2_u11_u7_U86 (.ZN( u2_out11_21 ) , .A4( u2_u11_u7_n157 ) , .A3( u2_u11_u7_n158 ) , .A2( u2_u11_u7_n159 ) , .A1( u2_u11_u7_n160 ) );
  OAI21_X1 u2_u11_u7_U87 (.B1( u2_u11_u7_n145 ) , .ZN( u2_u11_u7_n160 ) , .A( u2_u11_u7_n161 ) , .B2( u2_u11_u7_n177 ) );
  AOI22_X1 u2_u11_u7_U88 (.B2( u2_u11_u7_n149 ) , .B1( u2_u11_u7_n150 ) , .A2( u2_u11_u7_n151 ) , .A1( u2_u11_u7_n152 ) , .ZN( u2_u11_u7_n158 ) );
  NAND4_X1 u2_u11_u7_U89 (.ZN( u2_out11_15 ) , .A4( u2_u11_u7_n142 ) , .A3( u2_u11_u7_n143 ) , .A2( u2_u11_u7_n144 ) , .A1( u2_u11_u7_n178 ) );
  OAI221_X1 u2_u11_u7_U9 (.C1( u2_u11_u7_n101 ) , .C2( u2_u11_u7_n147 ) , .ZN( u2_u11_u7_n155 ) , .B2( u2_u11_u7_n162 ) , .A( u2_u11_u7_n91 ) , .B1( u2_u11_u7_n92 ) );
  OR2_X1 u2_u11_u7_U90 (.A2( u2_u11_u7_n125 ) , .A1( u2_u11_u7_n129 ) , .ZN( u2_u11_u7_n144 ) );
  AOI22_X1 u2_u11_u7_U91 (.A2( u2_u11_u7_n126 ) , .ZN( u2_u11_u7_n143 ) , .B2( u2_u11_u7_n165 ) , .B1( u2_u11_u7_n173 ) , .A1( u2_u11_u7_n174 ) );
  NAND4_X1 u2_u11_u7_U92 (.ZN( u2_out11_5 ) , .A4( u2_u11_u7_n108 ) , .A3( u2_u11_u7_n109 ) , .A1( u2_u11_u7_n116 ) , .A2( u2_u11_u7_n123 ) );
  AOI22_X1 u2_u11_u7_U93 (.ZN( u2_u11_u7_n109 ) , .A2( u2_u11_u7_n126 ) , .B2( u2_u11_u7_n145 ) , .B1( u2_u11_u7_n156 ) , .A1( u2_u11_u7_n171 ) );
  NOR4_X1 u2_u11_u7_U94 (.A4( u2_u11_u7_n104 ) , .A3( u2_u11_u7_n105 ) , .A2( u2_u11_u7_n106 ) , .A1( u2_u11_u7_n107 ) , .ZN( u2_u11_u7_n108 ) );
  NAND3_X1 u2_u11_u7_U95 (.A3( u2_u11_u7_n146 ) , .A2( u2_u11_u7_n147 ) , .A1( u2_u11_u7_n148 ) , .ZN( u2_u11_u7_n151 ) );
  NAND3_X1 u2_u11_u7_U96 (.A3( u2_u11_u7_n131 ) , .A2( u2_u11_u7_n132 ) , .A1( u2_u11_u7_n133 ) , .ZN( u2_u11_u7_n135 ) );
  XOR2_X1 u2_u12_U1 (.B( u2_K13_9 ) , .A( u2_R11_6 ) , .Z( u2_u12_X_9 ) );
  XOR2_X1 u2_u12_U16 (.B( u2_K13_3 ) , .A( u2_R11_2 ) , .Z( u2_u12_X_3 ) );
  XOR2_X1 u2_u12_U2 (.B( u2_K13_8 ) , .A( u2_R11_5 ) , .Z( u2_u12_X_8 ) );
  XOR2_X1 u2_u12_U20 (.B( u2_K13_36 ) , .A( u2_R11_25 ) , .Z( u2_u12_X_36 ) );
  XOR2_X1 u2_u12_U21 (.B( u2_K13_35 ) , .A( u2_R11_24 ) , .Z( u2_u12_X_35 ) );
  XOR2_X1 u2_u12_U22 (.B( u2_K13_34 ) , .A( u2_R11_23 ) , .Z( u2_u12_X_34 ) );
  XOR2_X1 u2_u12_U23 (.B( u2_K13_33 ) , .A( u2_R11_22 ) , .Z( u2_u12_X_33 ) );
  XOR2_X1 u2_u12_U24 (.B( u2_K13_32 ) , .A( u2_R11_21 ) , .Z( u2_u12_X_32 ) );
  XOR2_X1 u2_u12_U25 (.B( u2_K13_31 ) , .A( u2_R11_20 ) , .Z( u2_u12_X_31 ) );
  XOR2_X1 u2_u12_U26 (.B( u2_K13_30 ) , .A( u2_R11_21 ) , .Z( u2_u12_X_30 ) );
  XOR2_X1 u2_u12_U27 (.B( u2_K13_2 ) , .A( u2_R11_1 ) , .Z( u2_u12_X_2 ) );
  XOR2_X1 u2_u12_U28 (.B( u2_K13_29 ) , .A( u2_R11_20 ) , .Z( u2_u12_X_29 ) );
  XOR2_X1 u2_u12_U29 (.B( u2_K13_28 ) , .A( u2_R11_19 ) , .Z( u2_u12_X_28 ) );
  XOR2_X1 u2_u12_U3 (.B( u2_K13_7 ) , .A( u2_R11_4 ) , .Z( u2_u12_X_7 ) );
  XOR2_X1 u2_u12_U30 (.B( u2_K13_27 ) , .A( u2_R11_18 ) , .Z( u2_u12_X_27 ) );
  XOR2_X1 u2_u12_U31 (.B( u2_K13_26 ) , .A( u2_R11_17 ) , .Z( u2_u12_X_26 ) );
  XOR2_X1 u2_u12_U32 (.B( u2_K13_25 ) , .A( u2_R11_16 ) , .Z( u2_u12_X_25 ) );
  XOR2_X1 u2_u12_U33 (.B( u2_K13_24 ) , .A( u2_R11_17 ) , .Z( u2_u12_X_24 ) );
  XOR2_X1 u2_u12_U34 (.B( u2_K13_23 ) , .A( u2_R11_16 ) , .Z( u2_u12_X_23 ) );
  XOR2_X1 u2_u12_U35 (.B( u2_K13_22 ) , .A( u2_R11_15 ) , .Z( u2_u12_X_22 ) );
  XOR2_X1 u2_u12_U36 (.B( u2_K13_21 ) , .A( u2_R11_14 ) , .Z( u2_u12_X_21 ) );
  XOR2_X1 u2_u12_U37 (.B( u2_K13_20 ) , .A( u2_R11_13 ) , .Z( u2_u12_X_20 ) );
  XOR2_X1 u2_u12_U38 (.B( u2_K13_1 ) , .A( u2_R11_32 ) , .Z( u2_u12_X_1 ) );
  XOR2_X1 u2_u12_U39 (.B( u2_K13_19 ) , .A( u2_R11_12 ) , .Z( u2_u12_X_19 ) );
  XOR2_X1 u2_u12_U4 (.B( u2_K13_6 ) , .A( u2_R11_5 ) , .Z( u2_u12_X_6 ) );
  XOR2_X1 u2_u12_U40 (.B( u2_K13_18 ) , .A( u2_R11_13 ) , .Z( u2_u12_X_18 ) );
  XOR2_X1 u2_u12_U41 (.B( u2_K13_17 ) , .A( u2_R11_12 ) , .Z( u2_u12_X_17 ) );
  XOR2_X1 u2_u12_U42 (.B( u2_K13_16 ) , .A( u2_R11_11 ) , .Z( u2_u12_X_16 ) );
  XOR2_X1 u2_u12_U43 (.B( u2_K13_15 ) , .A( u2_R11_10 ) , .Z( u2_u12_X_15 ) );
  XOR2_X1 u2_u12_U44 (.B( u2_K13_14 ) , .A( u2_R11_9 ) , .Z( u2_u12_X_14 ) );
  XOR2_X1 u2_u12_U45 (.B( u2_K13_13 ) , .A( u2_R11_8 ) , .Z( u2_u12_X_13 ) );
  XOR2_X1 u2_u12_U46 (.B( u2_K13_12 ) , .A( u2_R11_9 ) , .Z( u2_u12_X_12 ) );
  XOR2_X1 u2_u12_U47 (.B( u2_K13_11 ) , .A( u2_R11_8 ) , .Z( u2_u12_X_11 ) );
  XOR2_X1 u2_u12_U48 (.B( u2_K13_10 ) , .A( u2_R11_7 ) , .Z( u2_u12_X_10 ) );
  XOR2_X1 u2_u12_U5 (.B( u2_K13_5 ) , .A( u2_R11_4 ) , .Z( u2_u12_X_5 ) );
  XOR2_X1 u2_u12_U6 (.B( u2_K13_4 ) , .A( u2_R11_3 ) , .Z( u2_u12_X_4 ) );
  AND2_X1 u2_u12_u0_U10 (.A1( u2_u12_u0_n131 ) , .ZN( u2_u12_u0_n141 ) , .A2( u2_u12_u0_n150 ) );
  AND3_X1 u2_u12_u0_U11 (.A2( u2_u12_u0_n112 ) , .ZN( u2_u12_u0_n127 ) , .A3( u2_u12_u0_n130 ) , .A1( u2_u12_u0_n148 ) );
  AND2_X1 u2_u12_u0_U12 (.ZN( u2_u12_u0_n107 ) , .A1( u2_u12_u0_n130 ) , .A2( u2_u12_u0_n140 ) );
  AND2_X1 u2_u12_u0_U13 (.A2( u2_u12_u0_n129 ) , .A1( u2_u12_u0_n130 ) , .ZN( u2_u12_u0_n151 ) );
  AND2_X1 u2_u12_u0_U14 (.A1( u2_u12_u0_n108 ) , .A2( u2_u12_u0_n125 ) , .ZN( u2_u12_u0_n145 ) );
  INV_X1 u2_u12_u0_U15 (.A( u2_u12_u0_n143 ) , .ZN( u2_u12_u0_n173 ) );
  NOR2_X1 u2_u12_u0_U16 (.A2( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n147 ) , .A1( u2_u12_u0_n160 ) );
  AOI21_X1 u2_u12_u0_U17 (.B1( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n132 ) , .A( u2_u12_u0_n165 ) , .B2( u2_u12_u0_n93 ) );
  OAI22_X1 u2_u12_u0_U18 (.B1( u2_u12_u0_n125 ) , .ZN( u2_u12_u0_n126 ) , .A1( u2_u12_u0_n138 ) , .A2( u2_u12_u0_n146 ) , .B2( u2_u12_u0_n147 ) );
  OAI22_X1 u2_u12_u0_U19 (.B1( u2_u12_u0_n131 ) , .A1( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n147 ) , .A2( u2_u12_u0_n90 ) , .ZN( u2_u12_u0_n91 ) );
  AND3_X1 u2_u12_u0_U20 (.A3( u2_u12_u0_n121 ) , .A2( u2_u12_u0_n125 ) , .A1( u2_u12_u0_n148 ) , .ZN( u2_u12_u0_n90 ) );
  NOR2_X1 u2_u12_u0_U21 (.A1( u2_u12_u0_n163 ) , .A2( u2_u12_u0_n164 ) , .ZN( u2_u12_u0_n95 ) );
  AOI22_X1 u2_u12_u0_U22 (.B2( u2_u12_u0_n109 ) , .A2( u2_u12_u0_n110 ) , .ZN( u2_u12_u0_n111 ) , .B1( u2_u12_u0_n118 ) , .A1( u2_u12_u0_n160 ) );
  NAND2_X1 u2_u12_u0_U23 (.A1( u2_u12_u0_n100 ) , .A2( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n125 ) );
  INV_X1 u2_u12_u0_U24 (.A( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n161 ) );
  INV_X1 u2_u12_u0_U25 (.A( u2_u12_u0_n118 ) , .ZN( u2_u12_u0_n158 ) );
  AOI21_X1 u2_u12_u0_U26 (.B1( u2_u12_u0_n127 ) , .B2( u2_u12_u0_n129 ) , .A( u2_u12_u0_n138 ) , .ZN( u2_u12_u0_n96 ) );
  AOI21_X1 u2_u12_u0_U27 (.ZN( u2_u12_u0_n104 ) , .B1( u2_u12_u0_n107 ) , .B2( u2_u12_u0_n141 ) , .A( u2_u12_u0_n144 ) );
  NAND2_X1 u2_u12_u0_U28 (.A2( u2_u12_u0_n102 ) , .A1( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n149 ) );
  NAND2_X1 u2_u12_u0_U29 (.A2( u2_u12_u0_n100 ) , .ZN( u2_u12_u0_n131 ) , .A1( u2_u12_u0_n92 ) );
  INV_X1 u2_u12_u0_U3 (.A( u2_u12_u0_n113 ) , .ZN( u2_u12_u0_n166 ) );
  NAND2_X1 u2_u12_u0_U30 (.A2( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n114 ) , .A1( u2_u12_u0_n92 ) );
  NOR2_X1 u2_u12_u0_U31 (.A1( u2_u12_u0_n120 ) , .ZN( u2_u12_u0_n143 ) , .A2( u2_u12_u0_n167 ) );
  OAI221_X1 u2_u12_u0_U32 (.C1( u2_u12_u0_n112 ) , .ZN( u2_u12_u0_n120 ) , .B1( u2_u12_u0_n138 ) , .B2( u2_u12_u0_n141 ) , .C2( u2_u12_u0_n147 ) , .A( u2_u12_u0_n172 ) );
  AOI211_X1 u2_u12_u0_U33 (.B( u2_u12_u0_n115 ) , .A( u2_u12_u0_n116 ) , .C2( u2_u12_u0_n117 ) , .C1( u2_u12_u0_n118 ) , .ZN( u2_u12_u0_n119 ) );
  NAND2_X1 u2_u12_u0_U34 (.A1( u2_u12_u0_n101 ) , .A2( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n150 ) );
  INV_X1 u2_u12_u0_U35 (.A( u2_u12_u0_n138 ) , .ZN( u2_u12_u0_n160 ) );
  NAND2_X1 u2_u12_u0_U36 (.A2( u2_u12_u0_n100 ) , .A1( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n139 ) );
  NAND2_X1 u2_u12_u0_U37 (.ZN( u2_u12_u0_n112 ) , .A2( u2_u12_u0_n92 ) , .A1( u2_u12_u0_n93 ) );
  INV_X1 u2_u12_u0_U38 (.ZN( u2_u12_u0_n172 ) , .A( u2_u12_u0_n88 ) );
  OAI222_X1 u2_u12_u0_U39 (.C1( u2_u12_u0_n108 ) , .A1( u2_u12_u0_n125 ) , .B2( u2_u12_u0_n128 ) , .B1( u2_u12_u0_n144 ) , .A2( u2_u12_u0_n158 ) , .C2( u2_u12_u0_n161 ) , .ZN( u2_u12_u0_n88 ) );
  AOI21_X1 u2_u12_u0_U4 (.B1( u2_u12_u0_n114 ) , .ZN( u2_u12_u0_n115 ) , .B2( u2_u12_u0_n129 ) , .A( u2_u12_u0_n161 ) );
  NAND2_X1 u2_u12_u0_U40 (.A2( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n121 ) , .A1( u2_u12_u0_n93 ) );
  OR3_X1 u2_u12_u0_U41 (.A3( u2_u12_u0_n152 ) , .A2( u2_u12_u0_n153 ) , .A1( u2_u12_u0_n154 ) , .ZN( u2_u12_u0_n155 ) );
  AOI21_X1 u2_u12_u0_U42 (.B2( u2_u12_u0_n150 ) , .B1( u2_u12_u0_n151 ) , .ZN( u2_u12_u0_n152 ) , .A( u2_u12_u0_n158 ) );
  AOI21_X1 u2_u12_u0_U43 (.A( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n145 ) , .B1( u2_u12_u0_n146 ) , .ZN( u2_u12_u0_n154 ) );
  AOI21_X1 u2_u12_u0_U44 (.A( u2_u12_u0_n147 ) , .B2( u2_u12_u0_n148 ) , .B1( u2_u12_u0_n149 ) , .ZN( u2_u12_u0_n153 ) );
  INV_X1 u2_u12_u0_U45 (.ZN( u2_u12_u0_n171 ) , .A( u2_u12_u0_n99 ) );
  OAI211_X1 u2_u12_u0_U46 (.C2( u2_u12_u0_n140 ) , .C1( u2_u12_u0_n161 ) , .A( u2_u12_u0_n169 ) , .B( u2_u12_u0_n98 ) , .ZN( u2_u12_u0_n99 ) );
  INV_X1 u2_u12_u0_U47 (.ZN( u2_u12_u0_n169 ) , .A( u2_u12_u0_n91 ) );
  AOI211_X1 u2_u12_u0_U48 (.C1( u2_u12_u0_n118 ) , .A( u2_u12_u0_n123 ) , .B( u2_u12_u0_n96 ) , .C2( u2_u12_u0_n97 ) , .ZN( u2_u12_u0_n98 ) );
  NOR2_X1 u2_u12_u0_U49 (.A2( u2_u12_X_4 ) , .A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n118 ) );
  NOR2_X1 u2_u12_u0_U5 (.A1( u2_u12_u0_n108 ) , .ZN( u2_u12_u0_n123 ) , .A2( u2_u12_u0_n158 ) );
  NOR2_X1 u2_u12_u0_U50 (.A2( u2_u12_X_1 ) , .ZN( u2_u12_u0_n101 ) , .A1( u2_u12_u0_n163 ) );
  NAND2_X1 u2_u12_u0_U51 (.A2( u2_u12_X_4 ) , .A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n144 ) );
  NOR2_X1 u2_u12_u0_U52 (.A2( u2_u12_X_5 ) , .ZN( u2_u12_u0_n136 ) , .A1( u2_u12_u0_n159 ) );
  NAND2_X1 u2_u12_u0_U53 (.A1( u2_u12_X_5 ) , .ZN( u2_u12_u0_n138 ) , .A2( u2_u12_u0_n159 ) );
  AND2_X1 u2_u12_u0_U54 (.A2( u2_u12_X_3 ) , .A1( u2_u12_X_6 ) , .ZN( u2_u12_u0_n102 ) );
  INV_X1 u2_u12_u0_U55 (.A( u2_u12_X_4 ) , .ZN( u2_u12_u0_n159 ) );
  INV_X1 u2_u12_u0_U56 (.A( u2_u12_X_1 ) , .ZN( u2_u12_u0_n164 ) );
  INV_X1 u2_u12_u0_U57 (.A( u2_u12_X_3 ) , .ZN( u2_u12_u0_n162 ) );
  INV_X1 u2_u12_u0_U58 (.A( u2_u12_u0_n126 ) , .ZN( u2_u12_u0_n168 ) );
  AOI211_X1 u2_u12_u0_U59 (.B( u2_u12_u0_n133 ) , .A( u2_u12_u0_n134 ) , .C2( u2_u12_u0_n135 ) , .C1( u2_u12_u0_n136 ) , .ZN( u2_u12_u0_n137 ) );
  AOI21_X1 u2_u12_u0_U6 (.B2( u2_u12_u0_n131 ) , .ZN( u2_u12_u0_n134 ) , .B1( u2_u12_u0_n151 ) , .A( u2_u12_u0_n158 ) );
  OR4_X1 u2_u12_u0_U60 (.ZN( u2_out12_17 ) , .A4( u2_u12_u0_n122 ) , .A2( u2_u12_u0_n123 ) , .A1( u2_u12_u0_n124 ) , .A3( u2_u12_u0_n170 ) );
  AOI21_X1 u2_u12_u0_U61 (.B2( u2_u12_u0_n107 ) , .ZN( u2_u12_u0_n124 ) , .B1( u2_u12_u0_n128 ) , .A( u2_u12_u0_n161 ) );
  INV_X1 u2_u12_u0_U62 (.A( u2_u12_u0_n111 ) , .ZN( u2_u12_u0_n170 ) );
  OR4_X1 u2_u12_u0_U63 (.ZN( u2_out12_31 ) , .A4( u2_u12_u0_n155 ) , .A2( u2_u12_u0_n156 ) , .A1( u2_u12_u0_n157 ) , .A3( u2_u12_u0_n173 ) );
  AOI21_X1 u2_u12_u0_U64 (.A( u2_u12_u0_n138 ) , .B2( u2_u12_u0_n139 ) , .B1( u2_u12_u0_n140 ) , .ZN( u2_u12_u0_n157 ) );
  INV_X1 u2_u12_u0_U65 (.ZN( u2_u12_u0_n174 ) , .A( u2_u12_u0_n89 ) );
  AOI211_X1 u2_u12_u0_U66 (.B( u2_u12_u0_n104 ) , .A( u2_u12_u0_n105 ) , .ZN( u2_u12_u0_n106 ) , .C2( u2_u12_u0_n113 ) , .C1( u2_u12_u0_n160 ) );
  AOI21_X1 u2_u12_u0_U67 (.B2( u2_u12_u0_n141 ) , .B1( u2_u12_u0_n142 ) , .ZN( u2_u12_u0_n156 ) , .A( u2_u12_u0_n161 ) );
  AOI21_X1 u2_u12_u0_U68 (.ZN( u2_u12_u0_n116 ) , .B2( u2_u12_u0_n142 ) , .A( u2_u12_u0_n144 ) , .B1( u2_u12_u0_n166 ) );
  INV_X1 u2_u12_u0_U69 (.A( u2_u12_u0_n142 ) , .ZN( u2_u12_u0_n165 ) );
  OAI21_X1 u2_u12_u0_U7 (.B1( u2_u12_u0_n150 ) , .B2( u2_u12_u0_n158 ) , .A( u2_u12_u0_n172 ) , .ZN( u2_u12_u0_n89 ) );
  NAND2_X1 u2_u12_u0_U70 (.A2( u2_u12_u0_n103 ) , .ZN( u2_u12_u0_n140 ) , .A1( u2_u12_u0_n94 ) );
  NAND2_X1 u2_u12_u0_U71 (.A1( u2_u12_u0_n101 ) , .ZN( u2_u12_u0_n130 ) , .A2( u2_u12_u0_n94 ) );
  NAND2_X1 u2_u12_u0_U72 (.ZN( u2_u12_u0_n108 ) , .A1( u2_u12_u0_n92 ) , .A2( u2_u12_u0_n94 ) );
  AND2_X1 u2_u12_u0_U73 (.A1( u2_u12_X_6 ) , .A2( u2_u12_u0_n162 ) , .ZN( u2_u12_u0_n93 ) );
  NOR2_X1 u2_u12_u0_U74 (.A2( u2_u12_X_6 ) , .ZN( u2_u12_u0_n100 ) , .A1( u2_u12_u0_n162 ) );
  NOR2_X1 u2_u12_u0_U75 (.A2( u2_u12_X_3 ) , .A1( u2_u12_X_6 ) , .ZN( u2_u12_u0_n94 ) );
  OAI221_X1 u2_u12_u0_U76 (.C1( u2_u12_u0_n121 ) , .ZN( u2_u12_u0_n122 ) , .B2( u2_u12_u0_n127 ) , .A( u2_u12_u0_n143 ) , .B1( u2_u12_u0_n144 ) , .C2( u2_u12_u0_n147 ) );
  AOI21_X1 u2_u12_u0_U77 (.B1( u2_u12_u0_n132 ) , .ZN( u2_u12_u0_n133 ) , .A( u2_u12_u0_n144 ) , .B2( u2_u12_u0_n166 ) );
  OAI22_X1 u2_u12_u0_U78 (.ZN( u2_u12_u0_n105 ) , .A2( u2_u12_u0_n132 ) , .B1( u2_u12_u0_n146 ) , .A1( u2_u12_u0_n147 ) , .B2( u2_u12_u0_n161 ) );
  NAND2_X1 u2_u12_u0_U79 (.ZN( u2_u12_u0_n110 ) , .A2( u2_u12_u0_n132 ) , .A1( u2_u12_u0_n145 ) );
  AND2_X1 u2_u12_u0_U8 (.A1( u2_u12_u0_n114 ) , .A2( u2_u12_u0_n121 ) , .ZN( u2_u12_u0_n146 ) );
  INV_X1 u2_u12_u0_U80 (.A( u2_u12_u0_n119 ) , .ZN( u2_u12_u0_n167 ) );
  NAND2_X1 u2_u12_u0_U81 (.ZN( u2_u12_u0_n148 ) , .A1( u2_u12_u0_n93 ) , .A2( u2_u12_u0_n95 ) );
  NAND2_X1 u2_u12_u0_U82 (.A1( u2_u12_u0_n100 ) , .ZN( u2_u12_u0_n129 ) , .A2( u2_u12_u0_n95 ) );
  NAND2_X1 u2_u12_u0_U83 (.A1( u2_u12_u0_n102 ) , .ZN( u2_u12_u0_n128 ) , .A2( u2_u12_u0_n95 ) );
  NOR2_X1 u2_u12_u0_U84 (.A2( u2_u12_X_1 ) , .A1( u2_u12_X_2 ) , .ZN( u2_u12_u0_n92 ) );
  NAND2_X1 u2_u12_u0_U85 (.ZN( u2_u12_u0_n142 ) , .A1( u2_u12_u0_n94 ) , .A2( u2_u12_u0_n95 ) );
  NOR2_X1 u2_u12_u0_U86 (.A2( u2_u12_X_2 ) , .ZN( u2_u12_u0_n103 ) , .A1( u2_u12_u0_n164 ) );
  INV_X1 u2_u12_u0_U87 (.A( u2_u12_X_2 ) , .ZN( u2_u12_u0_n163 ) );
  NAND3_X1 u2_u12_u0_U88 (.ZN( u2_out12_23 ) , .A3( u2_u12_u0_n137 ) , .A1( u2_u12_u0_n168 ) , .A2( u2_u12_u0_n171 ) );
  NAND3_X1 u2_u12_u0_U89 (.A3( u2_u12_u0_n127 ) , .A2( u2_u12_u0_n128 ) , .ZN( u2_u12_u0_n135 ) , .A1( u2_u12_u0_n150 ) );
  NAND2_X1 u2_u12_u0_U9 (.ZN( u2_u12_u0_n113 ) , .A1( u2_u12_u0_n139 ) , .A2( u2_u12_u0_n149 ) );
  NAND3_X1 u2_u12_u0_U90 (.ZN( u2_u12_u0_n117 ) , .A3( u2_u12_u0_n132 ) , .A2( u2_u12_u0_n139 ) , .A1( u2_u12_u0_n148 ) );
  NAND3_X1 u2_u12_u0_U91 (.ZN( u2_u12_u0_n109 ) , .A2( u2_u12_u0_n114 ) , .A3( u2_u12_u0_n140 ) , .A1( u2_u12_u0_n149 ) );
  NAND3_X1 u2_u12_u0_U92 (.ZN( u2_out12_9 ) , .A3( u2_u12_u0_n106 ) , .A2( u2_u12_u0_n171 ) , .A1( u2_u12_u0_n174 ) );
  NAND3_X1 u2_u12_u0_U93 (.A2( u2_u12_u0_n128 ) , .A1( u2_u12_u0_n132 ) , .A3( u2_u12_u0_n146 ) , .ZN( u2_u12_u0_n97 ) );
  NOR2_X1 u2_u12_u1_U10 (.A1( u2_u12_u1_n112 ) , .A2( u2_u12_u1_n116 ) , .ZN( u2_u12_u1_n118 ) );
  NAND3_X1 u2_u12_u1_U100 (.ZN( u2_u12_u1_n113 ) , .A1( u2_u12_u1_n120 ) , .A3( u2_u12_u1_n133 ) , .A2( u2_u12_u1_n155 ) );
  OAI21_X1 u2_u12_u1_U11 (.ZN( u2_u12_u1_n101 ) , .B1( u2_u12_u1_n141 ) , .A( u2_u12_u1_n146 ) , .B2( u2_u12_u1_n183 ) );
  AOI21_X1 u2_u12_u1_U12 (.B2( u2_u12_u1_n155 ) , .B1( u2_u12_u1_n156 ) , .ZN( u2_u12_u1_n157 ) , .A( u2_u12_u1_n174 ) );
  NAND2_X1 u2_u12_u1_U13 (.ZN( u2_u12_u1_n140 ) , .A2( u2_u12_u1_n150 ) , .A1( u2_u12_u1_n155 ) );
  NAND2_X1 u2_u12_u1_U14 (.A1( u2_u12_u1_n131 ) , .ZN( u2_u12_u1_n147 ) , .A2( u2_u12_u1_n153 ) );
  INV_X1 u2_u12_u1_U15 (.A( u2_u12_u1_n139 ) , .ZN( u2_u12_u1_n174 ) );
  INV_X1 u2_u12_u1_U16 (.A( u2_u12_u1_n112 ) , .ZN( u2_u12_u1_n171 ) );
  NAND2_X1 u2_u12_u1_U17 (.ZN( u2_u12_u1_n141 ) , .A1( u2_u12_u1_n153 ) , .A2( u2_u12_u1_n156 ) );
  AND2_X1 u2_u12_u1_U18 (.A1( u2_u12_u1_n123 ) , .ZN( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n161 ) );
  NAND2_X1 u2_u12_u1_U19 (.A2( u2_u12_u1_n115 ) , .A1( u2_u12_u1_n116 ) , .ZN( u2_u12_u1_n148 ) );
  NAND2_X1 u2_u12_u1_U20 (.A2( u2_u12_u1_n133 ) , .A1( u2_u12_u1_n135 ) , .ZN( u2_u12_u1_n159 ) );
  NAND2_X1 u2_u12_u1_U21 (.A2( u2_u12_u1_n115 ) , .A1( u2_u12_u1_n120 ) , .ZN( u2_u12_u1_n132 ) );
  INV_X1 u2_u12_u1_U22 (.A( u2_u12_u1_n154 ) , .ZN( u2_u12_u1_n178 ) );
  INV_X1 u2_u12_u1_U23 (.A( u2_u12_u1_n151 ) , .ZN( u2_u12_u1_n183 ) );
  AND2_X1 u2_u12_u1_U24 (.A1( u2_u12_u1_n129 ) , .A2( u2_u12_u1_n133 ) , .ZN( u2_u12_u1_n149 ) );
  INV_X1 u2_u12_u1_U25 (.A( u2_u12_u1_n131 ) , .ZN( u2_u12_u1_n180 ) );
  OR4_X1 u2_u12_u1_U26 (.A4( u2_u12_u1_n106 ) , .A3( u2_u12_u1_n107 ) , .ZN( u2_u12_u1_n108 ) , .A1( u2_u12_u1_n117 ) , .A2( u2_u12_u1_n184 ) );
  AOI21_X1 u2_u12_u1_U27 (.ZN( u2_u12_u1_n106 ) , .A( u2_u12_u1_n112 ) , .B1( u2_u12_u1_n154 ) , .B2( u2_u12_u1_n156 ) );
  AOI21_X1 u2_u12_u1_U28 (.ZN( u2_u12_u1_n107 ) , .B1( u2_u12_u1_n134 ) , .B2( u2_u12_u1_n149 ) , .A( u2_u12_u1_n174 ) );
  INV_X1 u2_u12_u1_U29 (.A( u2_u12_u1_n101 ) , .ZN( u2_u12_u1_n184 ) );
  INV_X1 u2_u12_u1_U3 (.A( u2_u12_u1_n159 ) , .ZN( u2_u12_u1_n182 ) );
  AOI221_X1 u2_u12_u1_U30 (.B1( u2_u12_u1_n140 ) , .ZN( u2_u12_u1_n167 ) , .B2( u2_u12_u1_n172 ) , .C2( u2_u12_u1_n175 ) , .C1( u2_u12_u1_n178 ) , .A( u2_u12_u1_n188 ) );
  INV_X1 u2_u12_u1_U31 (.ZN( u2_u12_u1_n188 ) , .A( u2_u12_u1_n97 ) );
  AOI211_X1 u2_u12_u1_U32 (.A( u2_u12_u1_n118 ) , .C1( u2_u12_u1_n132 ) , .C2( u2_u12_u1_n139 ) , .B( u2_u12_u1_n96 ) , .ZN( u2_u12_u1_n97 ) );
  AOI21_X1 u2_u12_u1_U33 (.B2( u2_u12_u1_n121 ) , .B1( u2_u12_u1_n135 ) , .A( u2_u12_u1_n152 ) , .ZN( u2_u12_u1_n96 ) );
  OAI221_X1 u2_u12_u1_U34 (.A( u2_u12_u1_n119 ) , .C2( u2_u12_u1_n129 ) , .ZN( u2_u12_u1_n138 ) , .B2( u2_u12_u1_n152 ) , .C1( u2_u12_u1_n174 ) , .B1( u2_u12_u1_n187 ) );
  INV_X1 u2_u12_u1_U35 (.A( u2_u12_u1_n148 ) , .ZN( u2_u12_u1_n187 ) );
  AOI211_X1 u2_u12_u1_U36 (.B( u2_u12_u1_n117 ) , .A( u2_u12_u1_n118 ) , .ZN( u2_u12_u1_n119 ) , .C2( u2_u12_u1_n146 ) , .C1( u2_u12_u1_n159 ) );
  NOR2_X1 u2_u12_u1_U37 (.A1( u2_u12_u1_n168 ) , .A2( u2_u12_u1_n176 ) , .ZN( u2_u12_u1_n98 ) );
  AOI211_X1 u2_u12_u1_U38 (.B( u2_u12_u1_n162 ) , .A( u2_u12_u1_n163 ) , .C2( u2_u12_u1_n164 ) , .ZN( u2_u12_u1_n165 ) , .C1( u2_u12_u1_n171 ) );
  AOI21_X1 u2_u12_u1_U39 (.A( u2_u12_u1_n160 ) , .B2( u2_u12_u1_n161 ) , .ZN( u2_u12_u1_n162 ) , .B1( u2_u12_u1_n182 ) );
  AOI221_X1 u2_u12_u1_U4 (.A( u2_u12_u1_n138 ) , .C2( u2_u12_u1_n139 ) , .C1( u2_u12_u1_n140 ) , .B2( u2_u12_u1_n141 ) , .ZN( u2_u12_u1_n142 ) , .B1( u2_u12_u1_n175 ) );
  OR2_X1 u2_u12_u1_U40 (.A2( u2_u12_u1_n157 ) , .A1( u2_u12_u1_n158 ) , .ZN( u2_u12_u1_n163 ) );
  NAND2_X1 u2_u12_u1_U41 (.A1( u2_u12_u1_n128 ) , .ZN( u2_u12_u1_n146 ) , .A2( u2_u12_u1_n160 ) );
  NAND2_X1 u2_u12_u1_U42 (.A2( u2_u12_u1_n112 ) , .ZN( u2_u12_u1_n139 ) , .A1( u2_u12_u1_n152 ) );
  NAND2_X1 u2_u12_u1_U43 (.A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n156 ) , .A2( u2_u12_u1_n99 ) );
  NOR2_X1 u2_u12_u1_U44 (.ZN( u2_u12_u1_n117 ) , .A1( u2_u12_u1_n121 ) , .A2( u2_u12_u1_n160 ) );
  OAI21_X1 u2_u12_u1_U45 (.B2( u2_u12_u1_n123 ) , .ZN( u2_u12_u1_n145 ) , .B1( u2_u12_u1_n160 ) , .A( u2_u12_u1_n185 ) );
  INV_X1 u2_u12_u1_U46 (.A( u2_u12_u1_n122 ) , .ZN( u2_u12_u1_n185 ) );
  AOI21_X1 u2_u12_u1_U47 (.B2( u2_u12_u1_n120 ) , .B1( u2_u12_u1_n121 ) , .ZN( u2_u12_u1_n122 ) , .A( u2_u12_u1_n128 ) );
  AOI21_X1 u2_u12_u1_U48 (.A( u2_u12_u1_n128 ) , .B2( u2_u12_u1_n129 ) , .ZN( u2_u12_u1_n130 ) , .B1( u2_u12_u1_n150 ) );
  NAND2_X1 u2_u12_u1_U49 (.ZN( u2_u12_u1_n112 ) , .A1( u2_u12_u1_n169 ) , .A2( u2_u12_u1_n170 ) );
  AOI211_X1 u2_u12_u1_U5 (.ZN( u2_u12_u1_n124 ) , .A( u2_u12_u1_n138 ) , .C2( u2_u12_u1_n139 ) , .B( u2_u12_u1_n145 ) , .C1( u2_u12_u1_n147 ) );
  NAND2_X1 u2_u12_u1_U50 (.ZN( u2_u12_u1_n129 ) , .A2( u2_u12_u1_n95 ) , .A1( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U51 (.A1( u2_u12_u1_n102 ) , .ZN( u2_u12_u1_n154 ) , .A2( u2_u12_u1_n99 ) );
  NAND2_X1 u2_u12_u1_U52 (.A2( u2_u12_u1_n100 ) , .ZN( u2_u12_u1_n135 ) , .A1( u2_u12_u1_n99 ) );
  AOI21_X1 u2_u12_u1_U53 (.A( u2_u12_u1_n152 ) , .B2( u2_u12_u1_n153 ) , .B1( u2_u12_u1_n154 ) , .ZN( u2_u12_u1_n158 ) );
  INV_X1 u2_u12_u1_U54 (.A( u2_u12_u1_n160 ) , .ZN( u2_u12_u1_n175 ) );
  NAND2_X1 u2_u12_u1_U55 (.A1( u2_u12_u1_n100 ) , .ZN( u2_u12_u1_n116 ) , .A2( u2_u12_u1_n95 ) );
  NAND2_X1 u2_u12_u1_U56 (.A1( u2_u12_u1_n102 ) , .ZN( u2_u12_u1_n131 ) , .A2( u2_u12_u1_n95 ) );
  NAND2_X1 u2_u12_u1_U57 (.A2( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n121 ) , .A1( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U58 (.A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n153 ) , .A2( u2_u12_u1_n98 ) );
  NAND2_X1 u2_u12_u1_U59 (.A2( u2_u12_u1_n104 ) , .A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n133 ) );
  AOI22_X1 u2_u12_u1_U6 (.B2( u2_u12_u1_n113 ) , .A2( u2_u12_u1_n114 ) , .ZN( u2_u12_u1_n125 ) , .A1( u2_u12_u1_n171 ) , .B1( u2_u12_u1_n173 ) );
  NAND2_X1 u2_u12_u1_U60 (.ZN( u2_u12_u1_n150 ) , .A2( u2_u12_u1_n98 ) , .A1( u2_u12_u1_n99 ) );
  NAND2_X1 u2_u12_u1_U61 (.A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n155 ) , .A2( u2_u12_u1_n95 ) );
  OAI21_X1 u2_u12_u1_U62 (.ZN( u2_u12_u1_n109 ) , .B1( u2_u12_u1_n129 ) , .B2( u2_u12_u1_n160 ) , .A( u2_u12_u1_n167 ) );
  NAND2_X1 u2_u12_u1_U63 (.A2( u2_u12_u1_n100 ) , .A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n120 ) );
  NAND2_X1 u2_u12_u1_U64 (.A1( u2_u12_u1_n102 ) , .A2( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n115 ) );
  NAND2_X1 u2_u12_u1_U65 (.A2( u2_u12_u1_n100 ) , .A1( u2_u12_u1_n104 ) , .ZN( u2_u12_u1_n151 ) );
  NAND2_X1 u2_u12_u1_U66 (.A2( u2_u12_u1_n103 ) , .A1( u2_u12_u1_n105 ) , .ZN( u2_u12_u1_n161 ) );
  INV_X1 u2_u12_u1_U67 (.A( u2_u12_u1_n152 ) , .ZN( u2_u12_u1_n173 ) );
  INV_X1 u2_u12_u1_U68 (.A( u2_u12_u1_n128 ) , .ZN( u2_u12_u1_n172 ) );
  NAND2_X1 u2_u12_u1_U69 (.A2( u2_u12_u1_n102 ) , .A1( u2_u12_u1_n103 ) , .ZN( u2_u12_u1_n123 ) );
  NAND2_X1 u2_u12_u1_U7 (.ZN( u2_u12_u1_n114 ) , .A1( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n156 ) );
  NOR2_X1 u2_u12_u1_U70 (.A2( u2_u12_X_7 ) , .A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n95 ) );
  NOR2_X1 u2_u12_u1_U71 (.A1( u2_u12_X_12 ) , .A2( u2_u12_X_9 ) , .ZN( u2_u12_u1_n100 ) );
  NOR2_X1 u2_u12_u1_U72 (.A2( u2_u12_X_8 ) , .A1( u2_u12_u1_n177 ) , .ZN( u2_u12_u1_n99 ) );
  NOR2_X1 u2_u12_u1_U73 (.A2( u2_u12_X_12 ) , .ZN( u2_u12_u1_n102 ) , .A1( u2_u12_u1_n176 ) );
  NOR2_X1 u2_u12_u1_U74 (.A2( u2_u12_X_9 ) , .ZN( u2_u12_u1_n105 ) , .A1( u2_u12_u1_n168 ) );
  NAND2_X1 u2_u12_u1_U75 (.A1( u2_u12_X_10 ) , .ZN( u2_u12_u1_n160 ) , .A2( u2_u12_u1_n169 ) );
  NAND2_X1 u2_u12_u1_U76 (.A2( u2_u12_X_10 ) , .A1( u2_u12_X_11 ) , .ZN( u2_u12_u1_n152 ) );
  NAND2_X1 u2_u12_u1_U77 (.A1( u2_u12_X_11 ) , .ZN( u2_u12_u1_n128 ) , .A2( u2_u12_u1_n170 ) );
  AND2_X1 u2_u12_u1_U78 (.A2( u2_u12_X_7 ) , .A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n104 ) );
  AND2_X1 u2_u12_u1_U79 (.A1( u2_u12_X_8 ) , .ZN( u2_u12_u1_n103 ) , .A2( u2_u12_u1_n177 ) );
  AOI22_X1 u2_u12_u1_U8 (.B2( u2_u12_u1_n136 ) , .A2( u2_u12_u1_n137 ) , .ZN( u2_u12_u1_n143 ) , .A1( u2_u12_u1_n171 ) , .B1( u2_u12_u1_n173 ) );
  INV_X1 u2_u12_u1_U80 (.A( u2_u12_X_10 ) , .ZN( u2_u12_u1_n170 ) );
  INV_X1 u2_u12_u1_U81 (.A( u2_u12_X_9 ) , .ZN( u2_u12_u1_n176 ) );
  INV_X1 u2_u12_u1_U82 (.A( u2_u12_X_11 ) , .ZN( u2_u12_u1_n169 ) );
  INV_X1 u2_u12_u1_U83 (.A( u2_u12_X_12 ) , .ZN( u2_u12_u1_n168 ) );
  INV_X1 u2_u12_u1_U84 (.A( u2_u12_X_7 ) , .ZN( u2_u12_u1_n177 ) );
  NAND4_X1 u2_u12_u1_U85 (.ZN( u2_out12_28 ) , .A4( u2_u12_u1_n124 ) , .A3( u2_u12_u1_n125 ) , .A2( u2_u12_u1_n126 ) , .A1( u2_u12_u1_n127 ) );
  OAI21_X1 u2_u12_u1_U86 (.ZN( u2_u12_u1_n127 ) , .B2( u2_u12_u1_n139 ) , .B1( u2_u12_u1_n175 ) , .A( u2_u12_u1_n183 ) );
  OAI21_X1 u2_u12_u1_U87 (.ZN( u2_u12_u1_n126 ) , .B2( u2_u12_u1_n140 ) , .A( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n178 ) );
  NAND4_X1 u2_u12_u1_U88 (.ZN( u2_out12_18 ) , .A4( u2_u12_u1_n165 ) , .A3( u2_u12_u1_n166 ) , .A1( u2_u12_u1_n167 ) , .A2( u2_u12_u1_n186 ) );
  AOI22_X1 u2_u12_u1_U89 (.B2( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n147 ) , .A2( u2_u12_u1_n148 ) , .ZN( u2_u12_u1_n166 ) , .A1( u2_u12_u1_n172 ) );
  INV_X1 u2_u12_u1_U9 (.A( u2_u12_u1_n147 ) , .ZN( u2_u12_u1_n181 ) );
  INV_X1 u2_u12_u1_U90 (.A( u2_u12_u1_n145 ) , .ZN( u2_u12_u1_n186 ) );
  NAND4_X1 u2_u12_u1_U91 (.ZN( u2_out12_2 ) , .A4( u2_u12_u1_n142 ) , .A3( u2_u12_u1_n143 ) , .A2( u2_u12_u1_n144 ) , .A1( u2_u12_u1_n179 ) );
  OAI21_X1 u2_u12_u1_U92 (.B2( u2_u12_u1_n132 ) , .ZN( u2_u12_u1_n144 ) , .A( u2_u12_u1_n146 ) , .B1( u2_u12_u1_n180 ) );
  INV_X1 u2_u12_u1_U93 (.A( u2_u12_u1_n130 ) , .ZN( u2_u12_u1_n179 ) );
  OR4_X1 u2_u12_u1_U94 (.ZN( u2_out12_13 ) , .A4( u2_u12_u1_n108 ) , .A3( u2_u12_u1_n109 ) , .A2( u2_u12_u1_n110 ) , .A1( u2_u12_u1_n111 ) );
  AOI21_X1 u2_u12_u1_U95 (.ZN( u2_u12_u1_n111 ) , .A( u2_u12_u1_n128 ) , .B2( u2_u12_u1_n131 ) , .B1( u2_u12_u1_n135 ) );
  AOI21_X1 u2_u12_u1_U96 (.ZN( u2_u12_u1_n110 ) , .A( u2_u12_u1_n116 ) , .B1( u2_u12_u1_n152 ) , .B2( u2_u12_u1_n160 ) );
  NAND3_X1 u2_u12_u1_U97 (.A3( u2_u12_u1_n149 ) , .A2( u2_u12_u1_n150 ) , .A1( u2_u12_u1_n151 ) , .ZN( u2_u12_u1_n164 ) );
  NAND3_X1 u2_u12_u1_U98 (.A3( u2_u12_u1_n134 ) , .A2( u2_u12_u1_n135 ) , .ZN( u2_u12_u1_n136 ) , .A1( u2_u12_u1_n151 ) );
  NAND3_X1 u2_u12_u1_U99 (.A1( u2_u12_u1_n133 ) , .ZN( u2_u12_u1_n137 ) , .A2( u2_u12_u1_n154 ) , .A3( u2_u12_u1_n181 ) );
  OAI22_X1 u2_u12_u2_U10 (.B1( u2_u12_u2_n151 ) , .A2( u2_u12_u2_n152 ) , .A1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n160 ) , .B2( u2_u12_u2_n168 ) );
  NAND3_X1 u2_u12_u2_U100 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n98 ) );
  NOR3_X1 u2_u12_u2_U11 (.A1( u2_u12_u2_n150 ) , .ZN( u2_u12_u2_n151 ) , .A3( u2_u12_u2_n175 ) , .A2( u2_u12_u2_n188 ) );
  AOI21_X1 u2_u12_u2_U12 (.B2( u2_u12_u2_n123 ) , .ZN( u2_u12_u2_n125 ) , .A( u2_u12_u2_n171 ) , .B1( u2_u12_u2_n184 ) );
  INV_X1 u2_u12_u2_U13 (.A( u2_u12_u2_n150 ) , .ZN( u2_u12_u2_n184 ) );
  AOI21_X1 u2_u12_u2_U14 (.ZN( u2_u12_u2_n144 ) , .B2( u2_u12_u2_n155 ) , .A( u2_u12_u2_n172 ) , .B1( u2_u12_u2_n185 ) );
  AOI21_X1 u2_u12_u2_U15 (.B2( u2_u12_u2_n143 ) , .ZN( u2_u12_u2_n145 ) , .B1( u2_u12_u2_n152 ) , .A( u2_u12_u2_n171 ) );
  INV_X1 u2_u12_u2_U16 (.A( u2_u12_u2_n156 ) , .ZN( u2_u12_u2_n171 ) );
  INV_X1 u2_u12_u2_U17 (.A( u2_u12_u2_n120 ) , .ZN( u2_u12_u2_n188 ) );
  NAND2_X1 u2_u12_u2_U18 (.A2( u2_u12_u2_n122 ) , .ZN( u2_u12_u2_n150 ) , .A1( u2_u12_u2_n152 ) );
  INV_X1 u2_u12_u2_U19 (.A( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n170 ) );
  INV_X1 u2_u12_u2_U20 (.A( u2_u12_u2_n137 ) , .ZN( u2_u12_u2_n173 ) );
  NAND2_X1 u2_u12_u2_U21 (.A1( u2_u12_u2_n132 ) , .A2( u2_u12_u2_n139 ) , .ZN( u2_u12_u2_n157 ) );
  INV_X1 u2_u12_u2_U22 (.A( u2_u12_u2_n113 ) , .ZN( u2_u12_u2_n178 ) );
  INV_X1 u2_u12_u2_U23 (.A( u2_u12_u2_n139 ) , .ZN( u2_u12_u2_n175 ) );
  INV_X1 u2_u12_u2_U24 (.A( u2_u12_u2_n155 ) , .ZN( u2_u12_u2_n181 ) );
  INV_X1 u2_u12_u2_U25 (.A( u2_u12_u2_n119 ) , .ZN( u2_u12_u2_n177 ) );
  INV_X1 u2_u12_u2_U26 (.A( u2_u12_u2_n116 ) , .ZN( u2_u12_u2_n180 ) );
  INV_X1 u2_u12_u2_U27 (.A( u2_u12_u2_n131 ) , .ZN( u2_u12_u2_n179 ) );
  INV_X1 u2_u12_u2_U28 (.A( u2_u12_u2_n154 ) , .ZN( u2_u12_u2_n176 ) );
  NAND2_X1 u2_u12_u2_U29 (.A2( u2_u12_u2_n116 ) , .A1( u2_u12_u2_n117 ) , .ZN( u2_u12_u2_n118 ) );
  NOR2_X1 u2_u12_u2_U3 (.ZN( u2_u12_u2_n121 ) , .A2( u2_u12_u2_n177 ) , .A1( u2_u12_u2_n180 ) );
  INV_X1 u2_u12_u2_U30 (.A( u2_u12_u2_n132 ) , .ZN( u2_u12_u2_n182 ) );
  INV_X1 u2_u12_u2_U31 (.A( u2_u12_u2_n158 ) , .ZN( u2_u12_u2_n183 ) );
  OAI21_X1 u2_u12_u2_U32 (.A( u2_u12_u2_n156 ) , .B1( u2_u12_u2_n157 ) , .ZN( u2_u12_u2_n158 ) , .B2( u2_u12_u2_n179 ) );
  NOR2_X1 u2_u12_u2_U33 (.ZN( u2_u12_u2_n156 ) , .A1( u2_u12_u2_n166 ) , .A2( u2_u12_u2_n169 ) );
  NOR2_X1 u2_u12_u2_U34 (.A2( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n137 ) , .A1( u2_u12_u2_n140 ) );
  NOR2_X1 u2_u12_u2_U35 (.A2( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n153 ) , .A1( u2_u12_u2_n156 ) );
  AOI211_X1 u2_u12_u2_U36 (.ZN( u2_u12_u2_n130 ) , .C1( u2_u12_u2_n138 ) , .C2( u2_u12_u2_n179 ) , .B( u2_u12_u2_n96 ) , .A( u2_u12_u2_n97 ) );
  OAI22_X1 u2_u12_u2_U37 (.B1( u2_u12_u2_n133 ) , .A2( u2_u12_u2_n137 ) , .A1( u2_u12_u2_n152 ) , .B2( u2_u12_u2_n168 ) , .ZN( u2_u12_u2_n97 ) );
  OAI221_X1 u2_u12_u2_U38 (.B1( u2_u12_u2_n113 ) , .C1( u2_u12_u2_n132 ) , .A( u2_u12_u2_n149 ) , .B2( u2_u12_u2_n171 ) , .C2( u2_u12_u2_n172 ) , .ZN( u2_u12_u2_n96 ) );
  OAI221_X1 u2_u12_u2_U39 (.A( u2_u12_u2_n115 ) , .C2( u2_u12_u2_n123 ) , .B2( u2_u12_u2_n143 ) , .B1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n163 ) , .C1( u2_u12_u2_n168 ) );
  INV_X1 u2_u12_u2_U4 (.A( u2_u12_u2_n134 ) , .ZN( u2_u12_u2_n185 ) );
  OAI21_X1 u2_u12_u2_U40 (.A( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n115 ) , .B1( u2_u12_u2_n176 ) , .B2( u2_u12_u2_n178 ) );
  OAI221_X1 u2_u12_u2_U41 (.A( u2_u12_u2_n135 ) , .B2( u2_u12_u2_n136 ) , .B1( u2_u12_u2_n137 ) , .ZN( u2_u12_u2_n162 ) , .C2( u2_u12_u2_n167 ) , .C1( u2_u12_u2_n185 ) );
  AND3_X1 u2_u12_u2_U42 (.A3( u2_u12_u2_n131 ) , .A2( u2_u12_u2_n132 ) , .A1( u2_u12_u2_n133 ) , .ZN( u2_u12_u2_n136 ) );
  AOI22_X1 u2_u12_u2_U43 (.ZN( u2_u12_u2_n135 ) , .B1( u2_u12_u2_n140 ) , .A1( u2_u12_u2_n156 ) , .B2( u2_u12_u2_n180 ) , .A2( u2_u12_u2_n188 ) );
  AOI21_X1 u2_u12_u2_U44 (.ZN( u2_u12_u2_n149 ) , .B1( u2_u12_u2_n173 ) , .B2( u2_u12_u2_n188 ) , .A( u2_u12_u2_n95 ) );
  AND3_X1 u2_u12_u2_U45 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n156 ) , .ZN( u2_u12_u2_n95 ) );
  OAI21_X1 u2_u12_u2_U46 (.A( u2_u12_u2_n101 ) , .B2( u2_u12_u2_n121 ) , .B1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n164 ) );
  NAND2_X1 u2_u12_u2_U47 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n155 ) );
  NAND2_X1 u2_u12_u2_U48 (.A2( u2_u12_u2_n105 ) , .A1( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n143 ) );
  NAND2_X1 u2_u12_u2_U49 (.A1( u2_u12_u2_n104 ) , .A2( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n152 ) );
  NOR4_X1 u2_u12_u2_U5 (.A4( u2_u12_u2_n124 ) , .A3( u2_u12_u2_n125 ) , .A2( u2_u12_u2_n126 ) , .A1( u2_u12_u2_n127 ) , .ZN( u2_u12_u2_n128 ) );
  NAND2_X1 u2_u12_u2_U50 (.A1( u2_u12_u2_n100 ) , .A2( u2_u12_u2_n105 ) , .ZN( u2_u12_u2_n132 ) );
  INV_X1 u2_u12_u2_U51 (.A( u2_u12_u2_n140 ) , .ZN( u2_u12_u2_n168 ) );
  INV_X1 u2_u12_u2_U52 (.A( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n167 ) );
  OAI21_X1 u2_u12_u2_U53 (.A( u2_u12_u2_n141 ) , .B2( u2_u12_u2_n142 ) , .ZN( u2_u12_u2_n146 ) , .B1( u2_u12_u2_n153 ) );
  OAI21_X1 u2_u12_u2_U54 (.A( u2_u12_u2_n140 ) , .ZN( u2_u12_u2_n141 ) , .B1( u2_u12_u2_n176 ) , .B2( u2_u12_u2_n177 ) );
  NOR3_X1 u2_u12_u2_U55 (.ZN( u2_u12_u2_n142 ) , .A3( u2_u12_u2_n175 ) , .A2( u2_u12_u2_n178 ) , .A1( u2_u12_u2_n181 ) );
  NAND2_X1 u2_u12_u2_U56 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n113 ) );
  NAND2_X1 u2_u12_u2_U57 (.A1( u2_u12_u2_n106 ) , .A2( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n131 ) );
  NAND2_X1 u2_u12_u2_U58 (.A1( u2_u12_u2_n103 ) , .A2( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n139 ) );
  NAND2_X1 u2_u12_u2_U59 (.A1( u2_u12_u2_n103 ) , .A2( u2_u12_u2_n105 ) , .ZN( u2_u12_u2_n133 ) );
  AOI21_X1 u2_u12_u2_U6 (.B2( u2_u12_u2_n119 ) , .ZN( u2_u12_u2_n127 ) , .A( u2_u12_u2_n137 ) , .B1( u2_u12_u2_n155 ) );
  NAND2_X1 u2_u12_u2_U60 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n103 ) , .ZN( u2_u12_u2_n154 ) );
  NAND2_X1 u2_u12_u2_U61 (.A2( u2_u12_u2_n103 ) , .A1( u2_u12_u2_n104 ) , .ZN( u2_u12_u2_n119 ) );
  NAND2_X1 u2_u12_u2_U62 (.A2( u2_u12_u2_n107 ) , .A1( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n123 ) );
  NAND2_X1 u2_u12_u2_U63 (.A1( u2_u12_u2_n104 ) , .A2( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n122 ) );
  INV_X1 u2_u12_u2_U64 (.A( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n172 ) );
  NAND2_X1 u2_u12_u2_U65 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n102 ) , .ZN( u2_u12_u2_n116 ) );
  NAND2_X1 u2_u12_u2_U66 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n120 ) );
  NAND2_X1 u2_u12_u2_U67 (.A2( u2_u12_u2_n105 ) , .A1( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n117 ) );
  INV_X1 u2_u12_u2_U68 (.ZN( u2_u12_u2_n187 ) , .A( u2_u12_u2_n99 ) );
  OAI21_X1 u2_u12_u2_U69 (.B1( u2_u12_u2_n137 ) , .B2( u2_u12_u2_n143 ) , .A( u2_u12_u2_n98 ) , .ZN( u2_u12_u2_n99 ) );
  AOI21_X1 u2_u12_u2_U7 (.ZN( u2_u12_u2_n124 ) , .B1( u2_u12_u2_n131 ) , .B2( u2_u12_u2_n143 ) , .A( u2_u12_u2_n172 ) );
  NOR2_X1 u2_u12_u2_U70 (.A2( u2_u12_X_16 ) , .ZN( u2_u12_u2_n140 ) , .A1( u2_u12_u2_n166 ) );
  NOR2_X1 u2_u12_u2_U71 (.A2( u2_u12_X_13 ) , .A1( u2_u12_X_14 ) , .ZN( u2_u12_u2_n100 ) );
  NOR2_X1 u2_u12_u2_U72 (.A2( u2_u12_X_16 ) , .A1( u2_u12_X_17 ) , .ZN( u2_u12_u2_n138 ) );
  NOR2_X1 u2_u12_u2_U73 (.A2( u2_u12_X_15 ) , .A1( u2_u12_X_18 ) , .ZN( u2_u12_u2_n104 ) );
  NOR2_X1 u2_u12_u2_U74 (.A2( u2_u12_X_14 ) , .ZN( u2_u12_u2_n103 ) , .A1( u2_u12_u2_n174 ) );
  NOR2_X1 u2_u12_u2_U75 (.A2( u2_u12_X_15 ) , .ZN( u2_u12_u2_n102 ) , .A1( u2_u12_u2_n165 ) );
  NOR2_X1 u2_u12_u2_U76 (.A2( u2_u12_X_17 ) , .ZN( u2_u12_u2_n114 ) , .A1( u2_u12_u2_n169 ) );
  AND2_X1 u2_u12_u2_U77 (.A1( u2_u12_X_15 ) , .ZN( u2_u12_u2_n105 ) , .A2( u2_u12_u2_n165 ) );
  AND2_X1 u2_u12_u2_U78 (.A2( u2_u12_X_15 ) , .A1( u2_u12_X_18 ) , .ZN( u2_u12_u2_n107 ) );
  AND2_X1 u2_u12_u2_U79 (.A1( u2_u12_X_14 ) , .ZN( u2_u12_u2_n106 ) , .A2( u2_u12_u2_n174 ) );
  AOI21_X1 u2_u12_u2_U8 (.B2( u2_u12_u2_n120 ) , .B1( u2_u12_u2_n121 ) , .ZN( u2_u12_u2_n126 ) , .A( u2_u12_u2_n167 ) );
  AND2_X1 u2_u12_u2_U80 (.A1( u2_u12_X_13 ) , .A2( u2_u12_X_14 ) , .ZN( u2_u12_u2_n108 ) );
  INV_X1 u2_u12_u2_U81 (.A( u2_u12_X_16 ) , .ZN( u2_u12_u2_n169 ) );
  INV_X1 u2_u12_u2_U82 (.A( u2_u12_X_17 ) , .ZN( u2_u12_u2_n166 ) );
  INV_X1 u2_u12_u2_U83 (.A( u2_u12_X_13 ) , .ZN( u2_u12_u2_n174 ) );
  INV_X1 u2_u12_u2_U84 (.A( u2_u12_X_18 ) , .ZN( u2_u12_u2_n165 ) );
  NAND4_X1 u2_u12_u2_U85 (.ZN( u2_out12_30 ) , .A4( u2_u12_u2_n147 ) , .A3( u2_u12_u2_n148 ) , .A2( u2_u12_u2_n149 ) , .A1( u2_u12_u2_n187 ) );
  AOI21_X1 u2_u12_u2_U86 (.B2( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n148 ) , .A( u2_u12_u2_n162 ) , .B1( u2_u12_u2_n182 ) );
  NOR3_X1 u2_u12_u2_U87 (.A3( u2_u12_u2_n144 ) , .A2( u2_u12_u2_n145 ) , .A1( u2_u12_u2_n146 ) , .ZN( u2_u12_u2_n147 ) );
  NAND4_X1 u2_u12_u2_U88 (.ZN( u2_out12_24 ) , .A4( u2_u12_u2_n111 ) , .A3( u2_u12_u2_n112 ) , .A1( u2_u12_u2_n130 ) , .A2( u2_u12_u2_n187 ) );
  AOI221_X1 u2_u12_u2_U89 (.A( u2_u12_u2_n109 ) , .B1( u2_u12_u2_n110 ) , .ZN( u2_u12_u2_n111 ) , .C1( u2_u12_u2_n134 ) , .C2( u2_u12_u2_n170 ) , .B2( u2_u12_u2_n173 ) );
  OAI22_X1 u2_u12_u2_U9 (.ZN( u2_u12_u2_n109 ) , .A2( u2_u12_u2_n113 ) , .B2( u2_u12_u2_n133 ) , .B1( u2_u12_u2_n167 ) , .A1( u2_u12_u2_n168 ) );
  AOI21_X1 u2_u12_u2_U90 (.ZN( u2_u12_u2_n112 ) , .B2( u2_u12_u2_n156 ) , .A( u2_u12_u2_n164 ) , .B1( u2_u12_u2_n181 ) );
  NAND4_X1 u2_u12_u2_U91 (.ZN( u2_out12_16 ) , .A4( u2_u12_u2_n128 ) , .A3( u2_u12_u2_n129 ) , .A1( u2_u12_u2_n130 ) , .A2( u2_u12_u2_n186 ) );
  AOI22_X1 u2_u12_u2_U92 (.A2( u2_u12_u2_n118 ) , .ZN( u2_u12_u2_n129 ) , .A1( u2_u12_u2_n140 ) , .B1( u2_u12_u2_n157 ) , .B2( u2_u12_u2_n170 ) );
  INV_X1 u2_u12_u2_U93 (.A( u2_u12_u2_n163 ) , .ZN( u2_u12_u2_n186 ) );
  OR4_X1 u2_u12_u2_U94 (.ZN( u2_out12_6 ) , .A4( u2_u12_u2_n161 ) , .A3( u2_u12_u2_n162 ) , .A2( u2_u12_u2_n163 ) , .A1( u2_u12_u2_n164 ) );
  OR3_X1 u2_u12_u2_U95 (.A2( u2_u12_u2_n159 ) , .A1( u2_u12_u2_n160 ) , .ZN( u2_u12_u2_n161 ) , .A3( u2_u12_u2_n183 ) );
  AOI21_X1 u2_u12_u2_U96 (.B2( u2_u12_u2_n154 ) , .B1( u2_u12_u2_n155 ) , .ZN( u2_u12_u2_n159 ) , .A( u2_u12_u2_n167 ) );
  NAND3_X1 u2_u12_u2_U97 (.A2( u2_u12_u2_n117 ) , .A1( u2_u12_u2_n122 ) , .A3( u2_u12_u2_n123 ) , .ZN( u2_u12_u2_n134 ) );
  NAND3_X1 u2_u12_u2_U98 (.ZN( u2_u12_u2_n110 ) , .A2( u2_u12_u2_n131 ) , .A3( u2_u12_u2_n139 ) , .A1( u2_u12_u2_n154 ) );
  NAND3_X1 u2_u12_u2_U99 (.A2( u2_u12_u2_n100 ) , .ZN( u2_u12_u2_n101 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n114 ) );
  OAI22_X1 u2_u12_u3_U10 (.B1( u2_u12_u3_n113 ) , .A2( u2_u12_u3_n135 ) , .A1( u2_u12_u3_n150 ) , .B2( u2_u12_u3_n164 ) , .ZN( u2_u12_u3_n98 ) );
  OAI211_X1 u2_u12_u3_U11 (.B( u2_u12_u3_n106 ) , .ZN( u2_u12_u3_n119 ) , .C2( u2_u12_u3_n128 ) , .C1( u2_u12_u3_n167 ) , .A( u2_u12_u3_n181 ) );
  AOI221_X1 u2_u12_u3_U12 (.C1( u2_u12_u3_n105 ) , .ZN( u2_u12_u3_n106 ) , .A( u2_u12_u3_n131 ) , .B2( u2_u12_u3_n132 ) , .C2( u2_u12_u3_n133 ) , .B1( u2_u12_u3_n169 ) );
  INV_X1 u2_u12_u3_U13 (.ZN( u2_u12_u3_n181 ) , .A( u2_u12_u3_n98 ) );
  NAND2_X1 u2_u12_u3_U14 (.ZN( u2_u12_u3_n105 ) , .A2( u2_u12_u3_n130 ) , .A1( u2_u12_u3_n155 ) );
  AOI22_X1 u2_u12_u3_U15 (.B1( u2_u12_u3_n115 ) , .A2( u2_u12_u3_n116 ) , .ZN( u2_u12_u3_n123 ) , .B2( u2_u12_u3_n133 ) , .A1( u2_u12_u3_n169 ) );
  NAND2_X1 u2_u12_u3_U16 (.ZN( u2_u12_u3_n116 ) , .A2( u2_u12_u3_n151 ) , .A1( u2_u12_u3_n182 ) );
  NOR2_X1 u2_u12_u3_U17 (.ZN( u2_u12_u3_n126 ) , .A2( u2_u12_u3_n150 ) , .A1( u2_u12_u3_n164 ) );
  AOI21_X1 u2_u12_u3_U18 (.ZN( u2_u12_u3_n112 ) , .B2( u2_u12_u3_n146 ) , .B1( u2_u12_u3_n155 ) , .A( u2_u12_u3_n167 ) );
  NAND2_X1 u2_u12_u3_U19 (.A1( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n142 ) , .A2( u2_u12_u3_n164 ) );
  NAND2_X1 u2_u12_u3_U20 (.ZN( u2_u12_u3_n132 ) , .A2( u2_u12_u3_n152 ) , .A1( u2_u12_u3_n156 ) );
  AND2_X1 u2_u12_u3_U21 (.A2( u2_u12_u3_n113 ) , .A1( u2_u12_u3_n114 ) , .ZN( u2_u12_u3_n151 ) );
  INV_X1 u2_u12_u3_U22 (.A( u2_u12_u3_n133 ) , .ZN( u2_u12_u3_n165 ) );
  INV_X1 u2_u12_u3_U23 (.A( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n170 ) );
  NAND2_X1 u2_u12_u3_U24 (.A1( u2_u12_u3_n107 ) , .A2( u2_u12_u3_n108 ) , .ZN( u2_u12_u3_n140 ) );
  NAND2_X1 u2_u12_u3_U25 (.ZN( u2_u12_u3_n117 ) , .A1( u2_u12_u3_n124 ) , .A2( u2_u12_u3_n148 ) );
  NAND2_X1 u2_u12_u3_U26 (.ZN( u2_u12_u3_n143 ) , .A1( u2_u12_u3_n165 ) , .A2( u2_u12_u3_n167 ) );
  INV_X1 u2_u12_u3_U27 (.A( u2_u12_u3_n130 ) , .ZN( u2_u12_u3_n177 ) );
  INV_X1 u2_u12_u3_U28 (.A( u2_u12_u3_n128 ) , .ZN( u2_u12_u3_n176 ) );
  INV_X1 u2_u12_u3_U29 (.A( u2_u12_u3_n155 ) , .ZN( u2_u12_u3_n174 ) );
  INV_X1 u2_u12_u3_U3 (.A( u2_u12_u3_n129 ) , .ZN( u2_u12_u3_n183 ) );
  INV_X1 u2_u12_u3_U30 (.A( u2_u12_u3_n139 ) , .ZN( u2_u12_u3_n185 ) );
  NOR2_X1 u2_u12_u3_U31 (.ZN( u2_u12_u3_n135 ) , .A2( u2_u12_u3_n141 ) , .A1( u2_u12_u3_n169 ) );
  OAI222_X1 u2_u12_u3_U32 (.C2( u2_u12_u3_n107 ) , .A2( u2_u12_u3_n108 ) , .B1( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n138 ) , .B2( u2_u12_u3_n146 ) , .C1( u2_u12_u3_n154 ) , .A1( u2_u12_u3_n164 ) );
  NOR4_X1 u2_u12_u3_U33 (.A4( u2_u12_u3_n157 ) , .A3( u2_u12_u3_n158 ) , .A2( u2_u12_u3_n159 ) , .A1( u2_u12_u3_n160 ) , .ZN( u2_u12_u3_n161 ) );
  AOI21_X1 u2_u12_u3_U34 (.B2( u2_u12_u3_n152 ) , .B1( u2_u12_u3_n153 ) , .ZN( u2_u12_u3_n158 ) , .A( u2_u12_u3_n164 ) );
  AOI21_X1 u2_u12_u3_U35 (.A( u2_u12_u3_n154 ) , .B2( u2_u12_u3_n155 ) , .B1( u2_u12_u3_n156 ) , .ZN( u2_u12_u3_n157 ) );
  AOI21_X1 u2_u12_u3_U36 (.A( u2_u12_u3_n149 ) , .B2( u2_u12_u3_n150 ) , .B1( u2_u12_u3_n151 ) , .ZN( u2_u12_u3_n159 ) );
  AOI211_X1 u2_u12_u3_U37 (.ZN( u2_u12_u3_n109 ) , .A( u2_u12_u3_n119 ) , .C2( u2_u12_u3_n129 ) , .B( u2_u12_u3_n138 ) , .C1( u2_u12_u3_n141 ) );
  AOI211_X1 u2_u12_u3_U38 (.B( u2_u12_u3_n119 ) , .A( u2_u12_u3_n120 ) , .C2( u2_u12_u3_n121 ) , .ZN( u2_u12_u3_n122 ) , .C1( u2_u12_u3_n179 ) );
  INV_X1 u2_u12_u3_U39 (.A( u2_u12_u3_n156 ) , .ZN( u2_u12_u3_n179 ) );
  INV_X1 u2_u12_u3_U4 (.A( u2_u12_u3_n140 ) , .ZN( u2_u12_u3_n182 ) );
  OAI22_X1 u2_u12_u3_U40 (.B1( u2_u12_u3_n118 ) , .ZN( u2_u12_u3_n120 ) , .A1( u2_u12_u3_n135 ) , .B2( u2_u12_u3_n154 ) , .A2( u2_u12_u3_n178 ) );
  AND3_X1 u2_u12_u3_U41 (.ZN( u2_u12_u3_n118 ) , .A2( u2_u12_u3_n124 ) , .A1( u2_u12_u3_n144 ) , .A3( u2_u12_u3_n152 ) );
  INV_X1 u2_u12_u3_U42 (.A( u2_u12_u3_n121 ) , .ZN( u2_u12_u3_n164 ) );
  NAND2_X1 u2_u12_u3_U43 (.ZN( u2_u12_u3_n133 ) , .A1( u2_u12_u3_n154 ) , .A2( u2_u12_u3_n164 ) );
  OAI211_X1 u2_u12_u3_U44 (.B( u2_u12_u3_n127 ) , .ZN( u2_u12_u3_n139 ) , .C1( u2_u12_u3_n150 ) , .C2( u2_u12_u3_n154 ) , .A( u2_u12_u3_n184 ) );
  INV_X1 u2_u12_u3_U45 (.A( u2_u12_u3_n125 ) , .ZN( u2_u12_u3_n184 ) );
  AOI221_X1 u2_u12_u3_U46 (.A( u2_u12_u3_n126 ) , .ZN( u2_u12_u3_n127 ) , .C2( u2_u12_u3_n132 ) , .C1( u2_u12_u3_n169 ) , .B2( u2_u12_u3_n170 ) , .B1( u2_u12_u3_n174 ) );
  OAI22_X1 u2_u12_u3_U47 (.A1( u2_u12_u3_n124 ) , .ZN( u2_u12_u3_n125 ) , .B2( u2_u12_u3_n145 ) , .A2( u2_u12_u3_n165 ) , .B1( u2_u12_u3_n167 ) );
  NOR2_X1 u2_u12_u3_U48 (.A1( u2_u12_u3_n113 ) , .ZN( u2_u12_u3_n131 ) , .A2( u2_u12_u3_n154 ) );
  NAND2_X1 u2_u12_u3_U49 (.A1( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n150 ) , .A2( u2_u12_u3_n99 ) );
  INV_X1 u2_u12_u3_U5 (.A( u2_u12_u3_n117 ) , .ZN( u2_u12_u3_n178 ) );
  NAND2_X1 u2_u12_u3_U50 (.A2( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n155 ) , .A1( u2_u12_u3_n97 ) );
  INV_X1 u2_u12_u3_U51 (.A( u2_u12_u3_n141 ) , .ZN( u2_u12_u3_n167 ) );
  AOI21_X1 u2_u12_u3_U52 (.B2( u2_u12_u3_n114 ) , .B1( u2_u12_u3_n146 ) , .A( u2_u12_u3_n154 ) , .ZN( u2_u12_u3_n94 ) );
  AOI21_X1 u2_u12_u3_U53 (.ZN( u2_u12_u3_n110 ) , .B2( u2_u12_u3_n142 ) , .B1( u2_u12_u3_n186 ) , .A( u2_u12_u3_n95 ) );
  INV_X1 u2_u12_u3_U54 (.A( u2_u12_u3_n145 ) , .ZN( u2_u12_u3_n186 ) );
  AOI21_X1 u2_u12_u3_U55 (.B1( u2_u12_u3_n124 ) , .A( u2_u12_u3_n149 ) , .B2( u2_u12_u3_n155 ) , .ZN( u2_u12_u3_n95 ) );
  INV_X1 u2_u12_u3_U56 (.A( u2_u12_u3_n149 ) , .ZN( u2_u12_u3_n169 ) );
  NAND2_X1 u2_u12_u3_U57 (.ZN( u2_u12_u3_n124 ) , .A1( u2_u12_u3_n96 ) , .A2( u2_u12_u3_n97 ) );
  NAND2_X1 u2_u12_u3_U58 (.A2( u2_u12_u3_n100 ) , .ZN( u2_u12_u3_n146 ) , .A1( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U59 (.A1( u2_u12_u3_n101 ) , .ZN( u2_u12_u3_n145 ) , .A2( u2_u12_u3_n99 ) );
  AOI221_X1 u2_u12_u3_U6 (.A( u2_u12_u3_n131 ) , .C2( u2_u12_u3_n132 ) , .C1( u2_u12_u3_n133 ) , .ZN( u2_u12_u3_n134 ) , .B1( u2_u12_u3_n143 ) , .B2( u2_u12_u3_n177 ) );
  NAND2_X1 u2_u12_u3_U60 (.A1( u2_u12_u3_n100 ) , .ZN( u2_u12_u3_n156 ) , .A2( u2_u12_u3_n99 ) );
  NAND2_X1 u2_u12_u3_U61 (.A2( u2_u12_u3_n101 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n148 ) );
  NAND2_X1 u2_u12_u3_U62 (.A1( u2_u12_u3_n100 ) , .A2( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n128 ) );
  NAND2_X1 u2_u12_u3_U63 (.A2( u2_u12_u3_n101 ) , .A1( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n152 ) );
  NAND2_X1 u2_u12_u3_U64 (.A2( u2_u12_u3_n101 ) , .ZN( u2_u12_u3_n114 ) , .A1( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U65 (.ZN( u2_u12_u3_n107 ) , .A1( u2_u12_u3_n97 ) , .A2( u2_u12_u3_n99 ) );
  NAND2_X1 u2_u12_u3_U66 (.A2( u2_u12_u3_n100 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n113 ) );
  NAND2_X1 u2_u12_u3_U67 (.A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n153 ) , .A2( u2_u12_u3_n97 ) );
  NAND2_X1 u2_u12_u3_U68 (.A2( u2_u12_u3_n103 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n130 ) );
  NAND2_X1 u2_u12_u3_U69 (.A2( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n144 ) , .A1( u2_u12_u3_n96 ) );
  OAI22_X1 u2_u12_u3_U7 (.B2( u2_u12_u3_n147 ) , .A2( u2_u12_u3_n148 ) , .ZN( u2_u12_u3_n160 ) , .B1( u2_u12_u3_n165 ) , .A1( u2_u12_u3_n168 ) );
  NAND2_X1 u2_u12_u3_U70 (.A1( u2_u12_u3_n102 ) , .A2( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n108 ) );
  NOR2_X1 u2_u12_u3_U71 (.A2( u2_u12_X_19 ) , .A1( u2_u12_X_20 ) , .ZN( u2_u12_u3_n99 ) );
  NOR2_X1 u2_u12_u3_U72 (.A2( u2_u12_X_21 ) , .A1( u2_u12_X_24 ) , .ZN( u2_u12_u3_n103 ) );
  NOR2_X1 u2_u12_u3_U73 (.A2( u2_u12_X_24 ) , .A1( u2_u12_u3_n171 ) , .ZN( u2_u12_u3_n97 ) );
  NOR2_X1 u2_u12_u3_U74 (.A2( u2_u12_X_23 ) , .ZN( u2_u12_u3_n141 ) , .A1( u2_u12_u3_n166 ) );
  NOR2_X1 u2_u12_u3_U75 (.A2( u2_u12_X_19 ) , .A1( u2_u12_u3_n172 ) , .ZN( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U76 (.A1( u2_u12_X_22 ) , .A2( u2_u12_X_23 ) , .ZN( u2_u12_u3_n154 ) );
  NAND2_X1 u2_u12_u3_U77 (.A1( u2_u12_X_23 ) , .ZN( u2_u12_u3_n149 ) , .A2( u2_u12_u3_n166 ) );
  NOR2_X1 u2_u12_u3_U78 (.A2( u2_u12_X_22 ) , .A1( u2_u12_X_23 ) , .ZN( u2_u12_u3_n121 ) );
  AND2_X1 u2_u12_u3_U79 (.A1( u2_u12_X_24 ) , .ZN( u2_u12_u3_n101 ) , .A2( u2_u12_u3_n171 ) );
  AND3_X1 u2_u12_u3_U8 (.A3( u2_u12_u3_n144 ) , .A2( u2_u12_u3_n145 ) , .A1( u2_u12_u3_n146 ) , .ZN( u2_u12_u3_n147 ) );
  AND2_X1 u2_u12_u3_U80 (.A1( u2_u12_X_19 ) , .ZN( u2_u12_u3_n102 ) , .A2( u2_u12_u3_n172 ) );
  AND2_X1 u2_u12_u3_U81 (.A1( u2_u12_X_21 ) , .A2( u2_u12_X_24 ) , .ZN( u2_u12_u3_n100 ) );
  AND2_X1 u2_u12_u3_U82 (.A2( u2_u12_X_19 ) , .A1( u2_u12_X_20 ) , .ZN( u2_u12_u3_n104 ) );
  INV_X1 u2_u12_u3_U83 (.A( u2_u12_X_22 ) , .ZN( u2_u12_u3_n166 ) );
  INV_X1 u2_u12_u3_U84 (.A( u2_u12_X_21 ) , .ZN( u2_u12_u3_n171 ) );
  INV_X1 u2_u12_u3_U85 (.A( u2_u12_X_20 ) , .ZN( u2_u12_u3_n172 ) );
  OR4_X1 u2_u12_u3_U86 (.ZN( u2_out12_10 ) , .A4( u2_u12_u3_n136 ) , .A3( u2_u12_u3_n137 ) , .A1( u2_u12_u3_n138 ) , .A2( u2_u12_u3_n139 ) );
  OAI222_X1 u2_u12_u3_U87 (.C1( u2_u12_u3_n128 ) , .ZN( u2_u12_u3_n137 ) , .B1( u2_u12_u3_n148 ) , .A2( u2_u12_u3_n150 ) , .B2( u2_u12_u3_n154 ) , .C2( u2_u12_u3_n164 ) , .A1( u2_u12_u3_n167 ) );
  OAI221_X1 u2_u12_u3_U88 (.A( u2_u12_u3_n134 ) , .B2( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n136 ) , .C1( u2_u12_u3_n149 ) , .B1( u2_u12_u3_n151 ) , .C2( u2_u12_u3_n183 ) );
  NAND4_X1 u2_u12_u3_U89 (.ZN( u2_out12_26 ) , .A4( u2_u12_u3_n109 ) , .A3( u2_u12_u3_n110 ) , .A2( u2_u12_u3_n111 ) , .A1( u2_u12_u3_n173 ) );
  INV_X1 u2_u12_u3_U9 (.A( u2_u12_u3_n143 ) , .ZN( u2_u12_u3_n168 ) );
  INV_X1 u2_u12_u3_U90 (.ZN( u2_u12_u3_n173 ) , .A( u2_u12_u3_n94 ) );
  OAI21_X1 u2_u12_u3_U91 (.ZN( u2_u12_u3_n111 ) , .B2( u2_u12_u3_n117 ) , .A( u2_u12_u3_n133 ) , .B1( u2_u12_u3_n176 ) );
  NAND4_X1 u2_u12_u3_U92 (.ZN( u2_out12_20 ) , .A4( u2_u12_u3_n122 ) , .A3( u2_u12_u3_n123 ) , .A1( u2_u12_u3_n175 ) , .A2( u2_u12_u3_n180 ) );
  INV_X1 u2_u12_u3_U93 (.A( u2_u12_u3_n126 ) , .ZN( u2_u12_u3_n180 ) );
  INV_X1 u2_u12_u3_U94 (.A( u2_u12_u3_n112 ) , .ZN( u2_u12_u3_n175 ) );
  NAND4_X1 u2_u12_u3_U95 (.ZN( u2_out12_1 ) , .A4( u2_u12_u3_n161 ) , .A3( u2_u12_u3_n162 ) , .A2( u2_u12_u3_n163 ) , .A1( u2_u12_u3_n185 ) );
  NAND2_X1 u2_u12_u3_U96 (.ZN( u2_u12_u3_n163 ) , .A2( u2_u12_u3_n170 ) , .A1( u2_u12_u3_n176 ) );
  AOI22_X1 u2_u12_u3_U97 (.B2( u2_u12_u3_n140 ) , .B1( u2_u12_u3_n141 ) , .A2( u2_u12_u3_n142 ) , .ZN( u2_u12_u3_n162 ) , .A1( u2_u12_u3_n177 ) );
  NAND3_X1 u2_u12_u3_U98 (.A1( u2_u12_u3_n114 ) , .ZN( u2_u12_u3_n115 ) , .A2( u2_u12_u3_n145 ) , .A3( u2_u12_u3_n153 ) );
  NAND3_X1 u2_u12_u3_U99 (.ZN( u2_u12_u3_n129 ) , .A2( u2_u12_u3_n144 ) , .A1( u2_u12_u3_n153 ) , .A3( u2_u12_u3_n182 ) );
  OAI22_X1 u2_u12_u4_U10 (.B2( u2_u12_u4_n135 ) , .ZN( u2_u12_u4_n137 ) , .B1( u2_u12_u4_n153 ) , .A1( u2_u12_u4_n155 ) , .A2( u2_u12_u4_n171 ) );
  AND3_X1 u2_u12_u4_U11 (.A2( u2_u12_u4_n134 ) , .ZN( u2_u12_u4_n135 ) , .A3( u2_u12_u4_n145 ) , .A1( u2_u12_u4_n157 ) );
  NAND2_X1 u2_u12_u4_U12 (.ZN( u2_u12_u4_n132 ) , .A2( u2_u12_u4_n170 ) , .A1( u2_u12_u4_n173 ) );
  AOI21_X1 u2_u12_u4_U13 (.B2( u2_u12_u4_n160 ) , .B1( u2_u12_u4_n161 ) , .ZN( u2_u12_u4_n162 ) , .A( u2_u12_u4_n170 ) );
  AOI21_X1 u2_u12_u4_U14 (.ZN( u2_u12_u4_n107 ) , .B2( u2_u12_u4_n143 ) , .A( u2_u12_u4_n174 ) , .B1( u2_u12_u4_n184 ) );
  AOI21_X1 u2_u12_u4_U15 (.B2( u2_u12_u4_n158 ) , .B1( u2_u12_u4_n159 ) , .ZN( u2_u12_u4_n163 ) , .A( u2_u12_u4_n174 ) );
  AOI21_X1 u2_u12_u4_U16 (.A( u2_u12_u4_n153 ) , .B2( u2_u12_u4_n154 ) , .B1( u2_u12_u4_n155 ) , .ZN( u2_u12_u4_n165 ) );
  AOI21_X1 u2_u12_u4_U17 (.A( u2_u12_u4_n156 ) , .B2( u2_u12_u4_n157 ) , .ZN( u2_u12_u4_n164 ) , .B1( u2_u12_u4_n184 ) );
  INV_X1 u2_u12_u4_U18 (.A( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n170 ) );
  AND2_X1 u2_u12_u4_U19 (.A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n155 ) , .A1( u2_u12_u4_n160 ) );
  INV_X1 u2_u12_u4_U20 (.A( u2_u12_u4_n156 ) , .ZN( u2_u12_u4_n175 ) );
  NAND2_X1 u2_u12_u4_U21 (.A2( u2_u12_u4_n118 ) , .ZN( u2_u12_u4_n131 ) , .A1( u2_u12_u4_n147 ) );
  NAND2_X1 u2_u12_u4_U22 (.A1( u2_u12_u4_n119 ) , .A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n130 ) );
  NAND2_X1 u2_u12_u4_U23 (.ZN( u2_u12_u4_n117 ) , .A2( u2_u12_u4_n118 ) , .A1( u2_u12_u4_n148 ) );
  NAND2_X1 u2_u12_u4_U24 (.ZN( u2_u12_u4_n129 ) , .A1( u2_u12_u4_n134 ) , .A2( u2_u12_u4_n148 ) );
  AND3_X1 u2_u12_u4_U25 (.A1( u2_u12_u4_n119 ) , .A2( u2_u12_u4_n143 ) , .A3( u2_u12_u4_n154 ) , .ZN( u2_u12_u4_n161 ) );
  AND2_X1 u2_u12_u4_U26 (.A1( u2_u12_u4_n145 ) , .A2( u2_u12_u4_n147 ) , .ZN( u2_u12_u4_n159 ) );
  OR3_X1 u2_u12_u4_U27 (.A3( u2_u12_u4_n114 ) , .A2( u2_u12_u4_n115 ) , .A1( u2_u12_u4_n116 ) , .ZN( u2_u12_u4_n136 ) );
  AOI21_X1 u2_u12_u4_U28 (.A( u2_u12_u4_n113 ) , .ZN( u2_u12_u4_n116 ) , .B2( u2_u12_u4_n173 ) , .B1( u2_u12_u4_n174 ) );
  AOI21_X1 u2_u12_u4_U29 (.ZN( u2_u12_u4_n115 ) , .B2( u2_u12_u4_n145 ) , .B1( u2_u12_u4_n146 ) , .A( u2_u12_u4_n156 ) );
  NOR2_X1 u2_u12_u4_U3 (.ZN( u2_u12_u4_n121 ) , .A1( u2_u12_u4_n181 ) , .A2( u2_u12_u4_n182 ) );
  OAI22_X1 u2_u12_u4_U30 (.ZN( u2_u12_u4_n114 ) , .A2( u2_u12_u4_n121 ) , .B1( u2_u12_u4_n160 ) , .B2( u2_u12_u4_n170 ) , .A1( u2_u12_u4_n171 ) );
  INV_X1 u2_u12_u4_U31 (.A( u2_u12_u4_n158 ) , .ZN( u2_u12_u4_n182 ) );
  INV_X1 u2_u12_u4_U32 (.ZN( u2_u12_u4_n181 ) , .A( u2_u12_u4_n96 ) );
  INV_X1 u2_u12_u4_U33 (.A( u2_u12_u4_n144 ) , .ZN( u2_u12_u4_n179 ) );
  INV_X1 u2_u12_u4_U34 (.A( u2_u12_u4_n157 ) , .ZN( u2_u12_u4_n178 ) );
  NAND2_X1 u2_u12_u4_U35 (.A2( u2_u12_u4_n154 ) , .A1( u2_u12_u4_n96 ) , .ZN( u2_u12_u4_n97 ) );
  INV_X1 u2_u12_u4_U36 (.ZN( u2_u12_u4_n186 ) , .A( u2_u12_u4_n95 ) );
  OAI221_X1 u2_u12_u4_U37 (.C1( u2_u12_u4_n134 ) , .B1( u2_u12_u4_n158 ) , .B2( u2_u12_u4_n171 ) , .C2( u2_u12_u4_n173 ) , .A( u2_u12_u4_n94 ) , .ZN( u2_u12_u4_n95 ) );
  AOI222_X1 u2_u12_u4_U38 (.B2( u2_u12_u4_n132 ) , .A1( u2_u12_u4_n138 ) , .C2( u2_u12_u4_n175 ) , .A2( u2_u12_u4_n179 ) , .C1( u2_u12_u4_n181 ) , .B1( u2_u12_u4_n185 ) , .ZN( u2_u12_u4_n94 ) );
  INV_X1 u2_u12_u4_U39 (.A( u2_u12_u4_n113 ) , .ZN( u2_u12_u4_n185 ) );
  INV_X1 u2_u12_u4_U4 (.A( u2_u12_u4_n117 ) , .ZN( u2_u12_u4_n184 ) );
  INV_X1 u2_u12_u4_U40 (.A( u2_u12_u4_n143 ) , .ZN( u2_u12_u4_n183 ) );
  NOR2_X1 u2_u12_u4_U41 (.ZN( u2_u12_u4_n138 ) , .A1( u2_u12_u4_n168 ) , .A2( u2_u12_u4_n169 ) );
  NOR2_X1 u2_u12_u4_U42 (.A1( u2_u12_u4_n150 ) , .A2( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n153 ) );
  NOR2_X1 u2_u12_u4_U43 (.A2( u2_u12_u4_n128 ) , .A1( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n156 ) );
  AOI22_X1 u2_u12_u4_U44 (.B2( u2_u12_u4_n122 ) , .A1( u2_u12_u4_n123 ) , .ZN( u2_u12_u4_n124 ) , .B1( u2_u12_u4_n128 ) , .A2( u2_u12_u4_n172 ) );
  INV_X1 u2_u12_u4_U45 (.A( u2_u12_u4_n153 ) , .ZN( u2_u12_u4_n172 ) );
  NAND2_X1 u2_u12_u4_U46 (.A2( u2_u12_u4_n120 ) , .ZN( u2_u12_u4_n123 ) , .A1( u2_u12_u4_n161 ) );
  AOI22_X1 u2_u12_u4_U47 (.B2( u2_u12_u4_n132 ) , .A2( u2_u12_u4_n133 ) , .ZN( u2_u12_u4_n140 ) , .A1( u2_u12_u4_n150 ) , .B1( u2_u12_u4_n179 ) );
  NAND2_X1 u2_u12_u4_U48 (.ZN( u2_u12_u4_n133 ) , .A2( u2_u12_u4_n146 ) , .A1( u2_u12_u4_n154 ) );
  NAND2_X1 u2_u12_u4_U49 (.A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n154 ) , .A2( u2_u12_u4_n98 ) );
  NOR4_X1 u2_u12_u4_U5 (.A4( u2_u12_u4_n106 ) , .A3( u2_u12_u4_n107 ) , .A2( u2_u12_u4_n108 ) , .A1( u2_u12_u4_n109 ) , .ZN( u2_u12_u4_n110 ) );
  NAND2_X1 u2_u12_u4_U50 (.A1( u2_u12_u4_n101 ) , .ZN( u2_u12_u4_n158 ) , .A2( u2_u12_u4_n99 ) );
  AOI21_X1 u2_u12_u4_U51 (.ZN( u2_u12_u4_n127 ) , .A( u2_u12_u4_n136 ) , .B2( u2_u12_u4_n150 ) , .B1( u2_u12_u4_n180 ) );
  INV_X1 u2_u12_u4_U52 (.A( u2_u12_u4_n160 ) , .ZN( u2_u12_u4_n180 ) );
  NAND2_X1 u2_u12_u4_U53 (.A2( u2_u12_u4_n104 ) , .A1( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n146 ) );
  NAND2_X1 u2_u12_u4_U54 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n160 ) );
  NAND2_X1 u2_u12_u4_U55 (.ZN( u2_u12_u4_n134 ) , .A1( u2_u12_u4_n98 ) , .A2( u2_u12_u4_n99 ) );
  NAND2_X1 u2_u12_u4_U56 (.A1( u2_u12_u4_n103 ) , .A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n143 ) );
  NAND2_X1 u2_u12_u4_U57 (.A2( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n145 ) , .A1( u2_u12_u4_n98 ) );
  NAND2_X1 u2_u12_u4_U58 (.A1( u2_u12_u4_n100 ) , .A2( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n120 ) );
  NAND2_X1 u2_u12_u4_U59 (.A1( u2_u12_u4_n102 ) , .A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n148 ) );
  AOI21_X1 u2_u12_u4_U6 (.ZN( u2_u12_u4_n106 ) , .B2( u2_u12_u4_n146 ) , .B1( u2_u12_u4_n158 ) , .A( u2_u12_u4_n170 ) );
  NAND2_X1 u2_u12_u4_U60 (.A2( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n157 ) );
  INV_X1 u2_u12_u4_U61 (.A( u2_u12_u4_n150 ) , .ZN( u2_u12_u4_n173 ) );
  INV_X1 u2_u12_u4_U62 (.A( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n171 ) );
  NAND2_X1 u2_u12_u4_U63 (.A1( u2_u12_u4_n100 ) , .ZN( u2_u12_u4_n118 ) , .A2( u2_u12_u4_n99 ) );
  NAND2_X1 u2_u12_u4_U64 (.A2( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n144 ) );
  NAND2_X1 u2_u12_u4_U65 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n105 ) , .ZN( u2_u12_u4_n96 ) );
  INV_X1 u2_u12_u4_U66 (.A( u2_u12_u4_n128 ) , .ZN( u2_u12_u4_n174 ) );
  NAND2_X1 u2_u12_u4_U67 (.A2( u2_u12_u4_n102 ) , .ZN( u2_u12_u4_n119 ) , .A1( u2_u12_u4_n98 ) );
  NAND2_X1 u2_u12_u4_U68 (.A2( u2_u12_u4_n101 ) , .A1( u2_u12_u4_n103 ) , .ZN( u2_u12_u4_n147 ) );
  NAND2_X1 u2_u12_u4_U69 (.A2( u2_u12_u4_n104 ) , .ZN( u2_u12_u4_n113 ) , .A1( u2_u12_u4_n99 ) );
  AOI21_X1 u2_u12_u4_U7 (.ZN( u2_u12_u4_n108 ) , .B2( u2_u12_u4_n134 ) , .B1( u2_u12_u4_n155 ) , .A( u2_u12_u4_n156 ) );
  NOR2_X1 u2_u12_u4_U70 (.A2( u2_u12_X_28 ) , .ZN( u2_u12_u4_n150 ) , .A1( u2_u12_u4_n168 ) );
  NOR2_X1 u2_u12_u4_U71 (.A2( u2_u12_X_29 ) , .ZN( u2_u12_u4_n152 ) , .A1( u2_u12_u4_n169 ) );
  NOR2_X1 u2_u12_u4_U72 (.A2( u2_u12_X_30 ) , .ZN( u2_u12_u4_n105 ) , .A1( u2_u12_u4_n176 ) );
  NOR2_X1 u2_u12_u4_U73 (.A2( u2_u12_X_26 ) , .ZN( u2_u12_u4_n100 ) , .A1( u2_u12_u4_n177 ) );
  NOR2_X1 u2_u12_u4_U74 (.A2( u2_u12_X_28 ) , .A1( u2_u12_X_29 ) , .ZN( u2_u12_u4_n128 ) );
  NOR2_X1 u2_u12_u4_U75 (.A2( u2_u12_X_27 ) , .A1( u2_u12_X_30 ) , .ZN( u2_u12_u4_n102 ) );
  NOR2_X1 u2_u12_u4_U76 (.A2( u2_u12_X_25 ) , .A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n98 ) );
  AND2_X1 u2_u12_u4_U77 (.A2( u2_u12_X_25 ) , .A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n104 ) );
  AND2_X1 u2_u12_u4_U78 (.A1( u2_u12_X_30 ) , .A2( u2_u12_u4_n176 ) , .ZN( u2_u12_u4_n99 ) );
  AND2_X1 u2_u12_u4_U79 (.A1( u2_u12_X_26 ) , .ZN( u2_u12_u4_n101 ) , .A2( u2_u12_u4_n177 ) );
  AOI21_X1 u2_u12_u4_U8 (.ZN( u2_u12_u4_n109 ) , .A( u2_u12_u4_n153 ) , .B1( u2_u12_u4_n159 ) , .B2( u2_u12_u4_n184 ) );
  AND2_X1 u2_u12_u4_U80 (.A1( u2_u12_X_27 ) , .A2( u2_u12_X_30 ) , .ZN( u2_u12_u4_n103 ) );
  INV_X1 u2_u12_u4_U81 (.A( u2_u12_X_28 ) , .ZN( u2_u12_u4_n169 ) );
  INV_X1 u2_u12_u4_U82 (.A( u2_u12_X_29 ) , .ZN( u2_u12_u4_n168 ) );
  INV_X1 u2_u12_u4_U83 (.A( u2_u12_X_25 ) , .ZN( u2_u12_u4_n177 ) );
  INV_X1 u2_u12_u4_U84 (.A( u2_u12_X_27 ) , .ZN( u2_u12_u4_n176 ) );
  NAND4_X1 u2_u12_u4_U85 (.ZN( u2_out12_25 ) , .A4( u2_u12_u4_n139 ) , .A3( u2_u12_u4_n140 ) , .A2( u2_u12_u4_n141 ) , .A1( u2_u12_u4_n142 ) );
  OAI21_X1 u2_u12_u4_U86 (.A( u2_u12_u4_n128 ) , .B2( u2_u12_u4_n129 ) , .B1( u2_u12_u4_n130 ) , .ZN( u2_u12_u4_n142 ) );
  OAI21_X1 u2_u12_u4_U87 (.B2( u2_u12_u4_n131 ) , .ZN( u2_u12_u4_n141 ) , .A( u2_u12_u4_n175 ) , .B1( u2_u12_u4_n183 ) );
  NAND4_X1 u2_u12_u4_U88 (.ZN( u2_out12_14 ) , .A4( u2_u12_u4_n124 ) , .A3( u2_u12_u4_n125 ) , .A2( u2_u12_u4_n126 ) , .A1( u2_u12_u4_n127 ) );
  AOI22_X1 u2_u12_u4_U89 (.B2( u2_u12_u4_n117 ) , .ZN( u2_u12_u4_n126 ) , .A1( u2_u12_u4_n129 ) , .B1( u2_u12_u4_n152 ) , .A2( u2_u12_u4_n175 ) );
  AOI211_X1 u2_u12_u4_U9 (.B( u2_u12_u4_n136 ) , .A( u2_u12_u4_n137 ) , .C2( u2_u12_u4_n138 ) , .ZN( u2_u12_u4_n139 ) , .C1( u2_u12_u4_n182 ) );
  AOI22_X1 u2_u12_u4_U90 (.ZN( u2_u12_u4_n125 ) , .B2( u2_u12_u4_n131 ) , .A2( u2_u12_u4_n132 ) , .B1( u2_u12_u4_n138 ) , .A1( u2_u12_u4_n178 ) );
  NAND4_X1 u2_u12_u4_U91 (.ZN( u2_out12_8 ) , .A4( u2_u12_u4_n110 ) , .A3( u2_u12_u4_n111 ) , .A2( u2_u12_u4_n112 ) , .A1( u2_u12_u4_n186 ) );
  NAND2_X1 u2_u12_u4_U92 (.ZN( u2_u12_u4_n112 ) , .A2( u2_u12_u4_n130 ) , .A1( u2_u12_u4_n150 ) );
  AOI22_X1 u2_u12_u4_U93 (.ZN( u2_u12_u4_n111 ) , .B2( u2_u12_u4_n132 ) , .A1( u2_u12_u4_n152 ) , .B1( u2_u12_u4_n178 ) , .A2( u2_u12_u4_n97 ) );
  AOI22_X1 u2_u12_u4_U94 (.B2( u2_u12_u4_n149 ) , .B1( u2_u12_u4_n150 ) , .A2( u2_u12_u4_n151 ) , .A1( u2_u12_u4_n152 ) , .ZN( u2_u12_u4_n167 ) );
  NOR4_X1 u2_u12_u4_U95 (.A4( u2_u12_u4_n162 ) , .A3( u2_u12_u4_n163 ) , .A2( u2_u12_u4_n164 ) , .A1( u2_u12_u4_n165 ) , .ZN( u2_u12_u4_n166 ) );
  NAND3_X1 u2_u12_u4_U96 (.ZN( u2_out12_3 ) , .A3( u2_u12_u4_n166 ) , .A1( u2_u12_u4_n167 ) , .A2( u2_u12_u4_n186 ) );
  NAND3_X1 u2_u12_u4_U97 (.A3( u2_u12_u4_n146 ) , .A2( u2_u12_u4_n147 ) , .A1( u2_u12_u4_n148 ) , .ZN( u2_u12_u4_n149 ) );
  NAND3_X1 u2_u12_u4_U98 (.A3( u2_u12_u4_n143 ) , .A2( u2_u12_u4_n144 ) , .A1( u2_u12_u4_n145 ) , .ZN( u2_u12_u4_n151 ) );
  NAND3_X1 u2_u12_u4_U99 (.A3( u2_u12_u4_n121 ) , .ZN( u2_u12_u4_n122 ) , .A2( u2_u12_u4_n144 ) , .A1( u2_u12_u4_n154 ) );
  INV_X1 u2_u12_u5_U10 (.A( u2_u12_u5_n121 ) , .ZN( u2_u12_u5_n177 ) );
  NOR3_X1 u2_u12_u5_U100 (.A3( u2_u12_u5_n141 ) , .A1( u2_u12_u5_n142 ) , .ZN( u2_u12_u5_n143 ) , .A2( u2_u12_u5_n191 ) );
  NAND4_X1 u2_u12_u5_U101 (.ZN( u2_out12_4 ) , .A4( u2_u12_u5_n112 ) , .A2( u2_u12_u5_n113 ) , .A1( u2_u12_u5_n114 ) , .A3( u2_u12_u5_n195 ) );
  AOI211_X1 u2_u12_u5_U102 (.A( u2_u12_u5_n110 ) , .C1( u2_u12_u5_n111 ) , .ZN( u2_u12_u5_n112 ) , .B( u2_u12_u5_n118 ) , .C2( u2_u12_u5_n177 ) );
  AOI222_X1 u2_u12_u5_U103 (.ZN( u2_u12_u5_n113 ) , .A1( u2_u12_u5_n131 ) , .C1( u2_u12_u5_n148 ) , .B2( u2_u12_u5_n174 ) , .C2( u2_u12_u5_n178 ) , .A2( u2_u12_u5_n179 ) , .B1( u2_u12_u5_n99 ) );
  NAND3_X1 u2_u12_u5_U104 (.A2( u2_u12_u5_n154 ) , .A3( u2_u12_u5_n158 ) , .A1( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n99 ) );
  NOR2_X1 u2_u12_u5_U11 (.ZN( u2_u12_u5_n160 ) , .A2( u2_u12_u5_n173 ) , .A1( u2_u12_u5_n177 ) );
  INV_X1 u2_u12_u5_U12 (.A( u2_u12_u5_n150 ) , .ZN( u2_u12_u5_n174 ) );
  AOI21_X1 u2_u12_u5_U13 (.A( u2_u12_u5_n160 ) , .B2( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n162 ) , .B1( u2_u12_u5_n192 ) );
  INV_X1 u2_u12_u5_U14 (.A( u2_u12_u5_n159 ) , .ZN( u2_u12_u5_n192 ) );
  AOI21_X1 u2_u12_u5_U15 (.A( u2_u12_u5_n156 ) , .B2( u2_u12_u5_n157 ) , .B1( u2_u12_u5_n158 ) , .ZN( u2_u12_u5_n163 ) );
  AOI21_X1 u2_u12_u5_U16 (.B2( u2_u12_u5_n139 ) , .B1( u2_u12_u5_n140 ) , .ZN( u2_u12_u5_n141 ) , .A( u2_u12_u5_n150 ) );
  OAI21_X1 u2_u12_u5_U17 (.A( u2_u12_u5_n133 ) , .B2( u2_u12_u5_n134 ) , .B1( u2_u12_u5_n135 ) , .ZN( u2_u12_u5_n142 ) );
  OAI21_X1 u2_u12_u5_U18 (.ZN( u2_u12_u5_n133 ) , .B2( u2_u12_u5_n147 ) , .A( u2_u12_u5_n173 ) , .B1( u2_u12_u5_n188 ) );
  NAND2_X1 u2_u12_u5_U19 (.A2( u2_u12_u5_n119 ) , .A1( u2_u12_u5_n123 ) , .ZN( u2_u12_u5_n137 ) );
  INV_X1 u2_u12_u5_U20 (.A( u2_u12_u5_n155 ) , .ZN( u2_u12_u5_n194 ) );
  NAND2_X1 u2_u12_u5_U21 (.A1( u2_u12_u5_n121 ) , .ZN( u2_u12_u5_n132 ) , .A2( u2_u12_u5_n172 ) );
  NAND2_X1 u2_u12_u5_U22 (.A2( u2_u12_u5_n122 ) , .ZN( u2_u12_u5_n136 ) , .A1( u2_u12_u5_n154 ) );
  NAND2_X1 u2_u12_u5_U23 (.A2( u2_u12_u5_n119 ) , .A1( u2_u12_u5_n120 ) , .ZN( u2_u12_u5_n159 ) );
  INV_X1 u2_u12_u5_U24 (.A( u2_u12_u5_n156 ) , .ZN( u2_u12_u5_n175 ) );
  INV_X1 u2_u12_u5_U25 (.A( u2_u12_u5_n158 ) , .ZN( u2_u12_u5_n188 ) );
  INV_X1 u2_u12_u5_U26 (.A( u2_u12_u5_n152 ) , .ZN( u2_u12_u5_n179 ) );
  INV_X1 u2_u12_u5_U27 (.A( u2_u12_u5_n140 ) , .ZN( u2_u12_u5_n182 ) );
  INV_X1 u2_u12_u5_U28 (.A( u2_u12_u5_n151 ) , .ZN( u2_u12_u5_n183 ) );
  INV_X1 u2_u12_u5_U29 (.A( u2_u12_u5_n123 ) , .ZN( u2_u12_u5_n185 ) );
  NOR2_X1 u2_u12_u5_U3 (.ZN( u2_u12_u5_n134 ) , .A1( u2_u12_u5_n183 ) , .A2( u2_u12_u5_n190 ) );
  INV_X1 u2_u12_u5_U30 (.A( u2_u12_u5_n161 ) , .ZN( u2_u12_u5_n184 ) );
  INV_X1 u2_u12_u5_U31 (.A( u2_u12_u5_n139 ) , .ZN( u2_u12_u5_n189 ) );
  INV_X1 u2_u12_u5_U32 (.A( u2_u12_u5_n157 ) , .ZN( u2_u12_u5_n190 ) );
  INV_X1 u2_u12_u5_U33 (.A( u2_u12_u5_n120 ) , .ZN( u2_u12_u5_n193 ) );
  NAND2_X1 u2_u12_u5_U34 (.ZN( u2_u12_u5_n111 ) , .A1( u2_u12_u5_n140 ) , .A2( u2_u12_u5_n155 ) );
  NOR2_X1 u2_u12_u5_U35 (.ZN( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n170 ) , .A2( u2_u12_u5_n180 ) );
  INV_X1 u2_u12_u5_U36 (.A( u2_u12_u5_n117 ) , .ZN( u2_u12_u5_n196 ) );
  OAI221_X1 u2_u12_u5_U37 (.A( u2_u12_u5_n116 ) , .ZN( u2_u12_u5_n117 ) , .B2( u2_u12_u5_n119 ) , .C1( u2_u12_u5_n153 ) , .C2( u2_u12_u5_n158 ) , .B1( u2_u12_u5_n172 ) );
  AOI222_X1 u2_u12_u5_U38 (.ZN( u2_u12_u5_n116 ) , .B2( u2_u12_u5_n145 ) , .C1( u2_u12_u5_n148 ) , .A2( u2_u12_u5_n174 ) , .C2( u2_u12_u5_n177 ) , .B1( u2_u12_u5_n187 ) , .A1( u2_u12_u5_n193 ) );
  INV_X1 u2_u12_u5_U39 (.A( u2_u12_u5_n115 ) , .ZN( u2_u12_u5_n187 ) );
  INV_X1 u2_u12_u5_U4 (.A( u2_u12_u5_n138 ) , .ZN( u2_u12_u5_n191 ) );
  AOI22_X1 u2_u12_u5_U40 (.B2( u2_u12_u5_n131 ) , .A2( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n169 ) , .B1( u2_u12_u5_n174 ) , .A1( u2_u12_u5_n185 ) );
  NOR2_X1 u2_u12_u5_U41 (.A1( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n150 ) , .A2( u2_u12_u5_n173 ) );
  AOI21_X1 u2_u12_u5_U42 (.A( u2_u12_u5_n118 ) , .B2( u2_u12_u5_n145 ) , .ZN( u2_u12_u5_n168 ) , .B1( u2_u12_u5_n186 ) );
  INV_X1 u2_u12_u5_U43 (.A( u2_u12_u5_n122 ) , .ZN( u2_u12_u5_n186 ) );
  NOR2_X1 u2_u12_u5_U44 (.A1( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n152 ) , .A2( u2_u12_u5_n176 ) );
  NOR2_X1 u2_u12_u5_U45 (.A1( u2_u12_u5_n115 ) , .ZN( u2_u12_u5_n118 ) , .A2( u2_u12_u5_n153 ) );
  NOR2_X1 u2_u12_u5_U46 (.A2( u2_u12_u5_n145 ) , .ZN( u2_u12_u5_n156 ) , .A1( u2_u12_u5_n174 ) );
  NOR2_X1 u2_u12_u5_U47 (.ZN( u2_u12_u5_n121 ) , .A2( u2_u12_u5_n145 ) , .A1( u2_u12_u5_n176 ) );
  AOI22_X1 u2_u12_u5_U48 (.ZN( u2_u12_u5_n114 ) , .A2( u2_u12_u5_n137 ) , .A1( u2_u12_u5_n145 ) , .B2( u2_u12_u5_n175 ) , .B1( u2_u12_u5_n193 ) );
  OAI211_X1 u2_u12_u5_U49 (.B( u2_u12_u5_n124 ) , .A( u2_u12_u5_n125 ) , .C2( u2_u12_u5_n126 ) , .C1( u2_u12_u5_n127 ) , .ZN( u2_u12_u5_n128 ) );
  OAI21_X1 u2_u12_u5_U5 (.B2( u2_u12_u5_n136 ) , .B1( u2_u12_u5_n137 ) , .ZN( u2_u12_u5_n138 ) , .A( u2_u12_u5_n177 ) );
  NOR3_X1 u2_u12_u5_U50 (.ZN( u2_u12_u5_n127 ) , .A1( u2_u12_u5_n136 ) , .A3( u2_u12_u5_n148 ) , .A2( u2_u12_u5_n182 ) );
  OAI21_X1 u2_u12_u5_U51 (.ZN( u2_u12_u5_n124 ) , .A( u2_u12_u5_n177 ) , .B2( u2_u12_u5_n183 ) , .B1( u2_u12_u5_n189 ) );
  OAI21_X1 u2_u12_u5_U52 (.ZN( u2_u12_u5_n125 ) , .A( u2_u12_u5_n174 ) , .B2( u2_u12_u5_n185 ) , .B1( u2_u12_u5_n190 ) );
  AOI21_X1 u2_u12_u5_U53 (.A( u2_u12_u5_n153 ) , .B2( u2_u12_u5_n154 ) , .B1( u2_u12_u5_n155 ) , .ZN( u2_u12_u5_n164 ) );
  AOI21_X1 u2_u12_u5_U54 (.ZN( u2_u12_u5_n110 ) , .B1( u2_u12_u5_n122 ) , .B2( u2_u12_u5_n139 ) , .A( u2_u12_u5_n153 ) );
  INV_X1 u2_u12_u5_U55 (.A( u2_u12_u5_n153 ) , .ZN( u2_u12_u5_n176 ) );
  INV_X1 u2_u12_u5_U56 (.A( u2_u12_u5_n126 ) , .ZN( u2_u12_u5_n173 ) );
  AND2_X1 u2_u12_u5_U57 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n147 ) );
  AND2_X1 u2_u12_u5_U58 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n148 ) );
  NAND2_X1 u2_u12_u5_U59 (.A1( u2_u12_u5_n105 ) , .A2( u2_u12_u5_n106 ) , .ZN( u2_u12_u5_n158 ) );
  INV_X1 u2_u12_u5_U6 (.A( u2_u12_u5_n135 ) , .ZN( u2_u12_u5_n178 ) );
  NAND2_X1 u2_u12_u5_U60 (.A2( u2_u12_u5_n108 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n139 ) );
  NAND2_X1 u2_u12_u5_U61 (.A1( u2_u12_u5_n106 ) , .A2( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n119 ) );
  NAND2_X1 u2_u12_u5_U62 (.A2( u2_u12_u5_n103 ) , .A1( u2_u12_u5_n105 ) , .ZN( u2_u12_u5_n140 ) );
  NAND2_X1 u2_u12_u5_U63 (.A2( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n105 ) , .ZN( u2_u12_u5_n155 ) );
  NAND2_X1 u2_u12_u5_U64 (.A2( u2_u12_u5_n106 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n122 ) );
  NAND2_X1 u2_u12_u5_U65 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n106 ) , .ZN( u2_u12_u5_n115 ) );
  NAND2_X1 u2_u12_u5_U66 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n103 ) , .ZN( u2_u12_u5_n161 ) );
  NAND2_X1 u2_u12_u5_U67 (.A1( u2_u12_u5_n105 ) , .A2( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n154 ) );
  INV_X1 u2_u12_u5_U68 (.A( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n172 ) );
  NAND2_X1 u2_u12_u5_U69 (.A1( u2_u12_u5_n103 ) , .A2( u2_u12_u5_n108 ) , .ZN( u2_u12_u5_n123 ) );
  OAI22_X1 u2_u12_u5_U7 (.B2( u2_u12_u5_n149 ) , .B1( u2_u12_u5_n150 ) , .A2( u2_u12_u5_n151 ) , .A1( u2_u12_u5_n152 ) , .ZN( u2_u12_u5_n165 ) );
  NAND2_X1 u2_u12_u5_U70 (.A2( u2_u12_u5_n103 ) , .A1( u2_u12_u5_n107 ) , .ZN( u2_u12_u5_n151 ) );
  NAND2_X1 u2_u12_u5_U71 (.A2( u2_u12_u5_n107 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n120 ) );
  NAND2_X1 u2_u12_u5_U72 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n109 ) , .ZN( u2_u12_u5_n157 ) );
  AND2_X1 u2_u12_u5_U73 (.A2( u2_u12_u5_n100 ) , .A1( u2_u12_u5_n104 ) , .ZN( u2_u12_u5_n131 ) );
  INV_X1 u2_u12_u5_U74 (.A( u2_u12_u5_n102 ) , .ZN( u2_u12_u5_n195 ) );
  OAI221_X1 u2_u12_u5_U75 (.A( u2_u12_u5_n101 ) , .ZN( u2_u12_u5_n102 ) , .C2( u2_u12_u5_n115 ) , .C1( u2_u12_u5_n126 ) , .B1( u2_u12_u5_n134 ) , .B2( u2_u12_u5_n160 ) );
  OAI21_X1 u2_u12_u5_U76 (.ZN( u2_u12_u5_n101 ) , .B1( u2_u12_u5_n137 ) , .A( u2_u12_u5_n146 ) , .B2( u2_u12_u5_n147 ) );
  NOR2_X1 u2_u12_u5_U77 (.A2( u2_u12_X_34 ) , .A1( u2_u12_X_35 ) , .ZN( u2_u12_u5_n145 ) );
  NOR2_X1 u2_u12_u5_U78 (.A2( u2_u12_X_34 ) , .ZN( u2_u12_u5_n146 ) , .A1( u2_u12_u5_n171 ) );
  NOR2_X1 u2_u12_u5_U79 (.A2( u2_u12_X_31 ) , .A1( u2_u12_X_32 ) , .ZN( u2_u12_u5_n103 ) );
  NOR3_X1 u2_u12_u5_U8 (.A2( u2_u12_u5_n147 ) , .A1( u2_u12_u5_n148 ) , .ZN( u2_u12_u5_n149 ) , .A3( u2_u12_u5_n194 ) );
  NOR2_X1 u2_u12_u5_U80 (.A2( u2_u12_X_36 ) , .ZN( u2_u12_u5_n105 ) , .A1( u2_u12_u5_n180 ) );
  NOR2_X1 u2_u12_u5_U81 (.A2( u2_u12_X_33 ) , .ZN( u2_u12_u5_n108 ) , .A1( u2_u12_u5_n170 ) );
  NOR2_X1 u2_u12_u5_U82 (.A2( u2_u12_X_33 ) , .A1( u2_u12_X_36 ) , .ZN( u2_u12_u5_n107 ) );
  NOR2_X1 u2_u12_u5_U83 (.A2( u2_u12_X_31 ) , .ZN( u2_u12_u5_n104 ) , .A1( u2_u12_u5_n181 ) );
  NAND2_X1 u2_u12_u5_U84 (.A2( u2_u12_X_34 ) , .A1( u2_u12_X_35 ) , .ZN( u2_u12_u5_n153 ) );
  NAND2_X1 u2_u12_u5_U85 (.A1( u2_u12_X_34 ) , .ZN( u2_u12_u5_n126 ) , .A2( u2_u12_u5_n171 ) );
  AND2_X1 u2_u12_u5_U86 (.A1( u2_u12_X_31 ) , .A2( u2_u12_X_32 ) , .ZN( u2_u12_u5_n106 ) );
  AND2_X1 u2_u12_u5_U87 (.A1( u2_u12_X_31 ) , .ZN( u2_u12_u5_n109 ) , .A2( u2_u12_u5_n181 ) );
  INV_X1 u2_u12_u5_U88 (.A( u2_u12_X_33 ) , .ZN( u2_u12_u5_n180 ) );
  INV_X1 u2_u12_u5_U89 (.A( u2_u12_X_35 ) , .ZN( u2_u12_u5_n171 ) );
  NOR2_X1 u2_u12_u5_U9 (.ZN( u2_u12_u5_n135 ) , .A1( u2_u12_u5_n173 ) , .A2( u2_u12_u5_n176 ) );
  INV_X1 u2_u12_u5_U90 (.A( u2_u12_X_36 ) , .ZN( u2_u12_u5_n170 ) );
  INV_X1 u2_u12_u5_U91 (.A( u2_u12_X_32 ) , .ZN( u2_u12_u5_n181 ) );
  NAND4_X1 u2_u12_u5_U92 (.ZN( u2_out12_29 ) , .A4( u2_u12_u5_n129 ) , .A3( u2_u12_u5_n130 ) , .A2( u2_u12_u5_n168 ) , .A1( u2_u12_u5_n196 ) );
  AOI221_X1 u2_u12_u5_U93 (.A( u2_u12_u5_n128 ) , .ZN( u2_u12_u5_n129 ) , .C2( u2_u12_u5_n132 ) , .B2( u2_u12_u5_n159 ) , .B1( u2_u12_u5_n176 ) , .C1( u2_u12_u5_n184 ) );
  AOI222_X1 u2_u12_u5_U94 (.ZN( u2_u12_u5_n130 ) , .A2( u2_u12_u5_n146 ) , .B1( u2_u12_u5_n147 ) , .C2( u2_u12_u5_n175 ) , .B2( u2_u12_u5_n179 ) , .A1( u2_u12_u5_n188 ) , .C1( u2_u12_u5_n194 ) );
  NAND4_X1 u2_u12_u5_U95 (.ZN( u2_out12_19 ) , .A4( u2_u12_u5_n166 ) , .A3( u2_u12_u5_n167 ) , .A2( u2_u12_u5_n168 ) , .A1( u2_u12_u5_n169 ) );
  AOI22_X1 u2_u12_u5_U96 (.B2( u2_u12_u5_n145 ) , .A2( u2_u12_u5_n146 ) , .ZN( u2_u12_u5_n167 ) , .B1( u2_u12_u5_n182 ) , .A1( u2_u12_u5_n189 ) );
  NOR4_X1 u2_u12_u5_U97 (.A4( u2_u12_u5_n162 ) , .A3( u2_u12_u5_n163 ) , .A2( u2_u12_u5_n164 ) , .A1( u2_u12_u5_n165 ) , .ZN( u2_u12_u5_n166 ) );
  NAND4_X1 u2_u12_u5_U98 (.ZN( u2_out12_11 ) , .A4( u2_u12_u5_n143 ) , .A3( u2_u12_u5_n144 ) , .A2( u2_u12_u5_n169 ) , .A1( u2_u12_u5_n196 ) );
  AOI22_X1 u2_u12_u5_U99 (.A2( u2_u12_u5_n132 ) , .ZN( u2_u12_u5_n144 ) , .B2( u2_u12_u5_n145 ) , .B1( u2_u12_u5_n184 ) , .A1( u2_u12_u5_n194 ) );
  XOR2_X1 u2_u14_U10 (.B( u2_K15_45 ) , .A( u2_R13_30 ) , .Z( u2_u14_X_45 ) );
  XOR2_X1 u2_u14_U11 (.B( u2_K15_44 ) , .A( u2_R13_29 ) , .Z( u2_u14_X_44 ) );
  XOR2_X1 u2_u14_U12 (.B( u2_K15_43 ) , .A( u2_R13_28 ) , .Z( u2_u14_X_43 ) );
  XOR2_X1 u2_u14_U33 (.B( u2_K15_24 ) , .A( u2_R13_17 ) , .Z( u2_u14_X_24 ) );
  XOR2_X1 u2_u14_U34 (.B( u2_K15_23 ) , .A( u2_R13_16 ) , .Z( u2_u14_X_23 ) );
  XOR2_X1 u2_u14_U35 (.B( u2_K15_22 ) , .A( u2_R13_15 ) , .Z( u2_u14_X_22 ) );
  XOR2_X1 u2_u14_U36 (.B( u2_K15_21 ) , .A( u2_R13_14 ) , .Z( u2_u14_X_21 ) );
  XOR2_X1 u2_u14_U37 (.B( u2_K15_20 ) , .A( u2_R13_13 ) , .Z( u2_u14_X_20 ) );
  XOR2_X1 u2_u14_U39 (.B( u2_K15_19 ) , .A( u2_R13_12 ) , .Z( u2_u14_X_19 ) );
  XOR2_X1 u2_u14_U40 (.B( u2_K15_18 ) , .A( u2_R13_13 ) , .Z( u2_u14_X_18 ) );
  XOR2_X1 u2_u14_U41 (.B( u2_K15_17 ) , .A( u2_R13_12 ) , .Z( u2_u14_X_17 ) );
  XOR2_X1 u2_u14_U42 (.B( u2_K15_16 ) , .A( u2_R13_11 ) , .Z( u2_u14_X_16 ) );
  XOR2_X1 u2_u14_U43 (.B( u2_K15_15 ) , .A( u2_R13_10 ) , .Z( u2_u14_X_15 ) );
  XOR2_X1 u2_u14_U44 (.B( u2_K15_14 ) , .A( u2_R13_9 ) , .Z( u2_u14_X_14 ) );
  XOR2_X1 u2_u14_U45 (.B( u2_K15_13 ) , .A( u2_R13_8 ) , .Z( u2_u14_X_13 ) );
  XOR2_X1 u2_u14_U7 (.B( u2_K15_48 ) , .A( u2_R13_1 ) , .Z( u2_u14_X_48 ) );
  XOR2_X1 u2_u14_U8 (.B( u2_K15_47 ) , .A( u2_R13_32 ) , .Z( u2_u14_X_47 ) );
  XOR2_X1 u2_u14_U9 (.B( u2_K15_46 ) , .A( u2_R13_31 ) , .Z( u2_u14_X_46 ) );
  OAI22_X1 u2_u14_u2_U10 (.ZN( u2_u14_u2_n109 ) , .A2( u2_u14_u2_n113 ) , .B2( u2_u14_u2_n133 ) , .B1( u2_u14_u2_n167 ) , .A1( u2_u14_u2_n168 ) );
  NAND3_X1 u2_u14_u2_U100 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n98 ) );
  OAI22_X1 u2_u14_u2_U11 (.B1( u2_u14_u2_n151 ) , .A2( u2_u14_u2_n152 ) , .A1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n160 ) , .B2( u2_u14_u2_n168 ) );
  NOR3_X1 u2_u14_u2_U12 (.A1( u2_u14_u2_n150 ) , .ZN( u2_u14_u2_n151 ) , .A3( u2_u14_u2_n175 ) , .A2( u2_u14_u2_n188 ) );
  AOI21_X1 u2_u14_u2_U13 (.ZN( u2_u14_u2_n144 ) , .B2( u2_u14_u2_n155 ) , .A( u2_u14_u2_n172 ) , .B1( u2_u14_u2_n185 ) );
  AOI21_X1 u2_u14_u2_U14 (.B2( u2_u14_u2_n143 ) , .ZN( u2_u14_u2_n145 ) , .B1( u2_u14_u2_n152 ) , .A( u2_u14_u2_n171 ) );
  AOI21_X1 u2_u14_u2_U15 (.B2( u2_u14_u2_n120 ) , .B1( u2_u14_u2_n121 ) , .ZN( u2_u14_u2_n126 ) , .A( u2_u14_u2_n167 ) );
  INV_X1 u2_u14_u2_U16 (.A( u2_u14_u2_n156 ) , .ZN( u2_u14_u2_n171 ) );
  INV_X1 u2_u14_u2_U17 (.A( u2_u14_u2_n120 ) , .ZN( u2_u14_u2_n188 ) );
  NAND2_X1 u2_u14_u2_U18 (.A2( u2_u14_u2_n122 ) , .ZN( u2_u14_u2_n150 ) , .A1( u2_u14_u2_n152 ) );
  INV_X1 u2_u14_u2_U19 (.A( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n170 ) );
  INV_X1 u2_u14_u2_U20 (.A( u2_u14_u2_n137 ) , .ZN( u2_u14_u2_n173 ) );
  NAND2_X1 u2_u14_u2_U21 (.A1( u2_u14_u2_n132 ) , .A2( u2_u14_u2_n139 ) , .ZN( u2_u14_u2_n157 ) );
  INV_X1 u2_u14_u2_U22 (.A( u2_u14_u2_n113 ) , .ZN( u2_u14_u2_n178 ) );
  INV_X1 u2_u14_u2_U23 (.A( u2_u14_u2_n139 ) , .ZN( u2_u14_u2_n175 ) );
  INV_X1 u2_u14_u2_U24 (.A( u2_u14_u2_n155 ) , .ZN( u2_u14_u2_n181 ) );
  INV_X1 u2_u14_u2_U25 (.A( u2_u14_u2_n119 ) , .ZN( u2_u14_u2_n177 ) );
  INV_X1 u2_u14_u2_U26 (.A( u2_u14_u2_n116 ) , .ZN( u2_u14_u2_n180 ) );
  INV_X1 u2_u14_u2_U27 (.A( u2_u14_u2_n131 ) , .ZN( u2_u14_u2_n179 ) );
  INV_X1 u2_u14_u2_U28 (.A( u2_u14_u2_n154 ) , .ZN( u2_u14_u2_n176 ) );
  NAND2_X1 u2_u14_u2_U29 (.A2( u2_u14_u2_n116 ) , .A1( u2_u14_u2_n117 ) , .ZN( u2_u14_u2_n118 ) );
  NOR2_X1 u2_u14_u2_U3 (.ZN( u2_u14_u2_n121 ) , .A2( u2_u14_u2_n177 ) , .A1( u2_u14_u2_n180 ) );
  INV_X1 u2_u14_u2_U30 (.A( u2_u14_u2_n132 ) , .ZN( u2_u14_u2_n182 ) );
  INV_X1 u2_u14_u2_U31 (.A( u2_u14_u2_n158 ) , .ZN( u2_u14_u2_n183 ) );
  OAI21_X1 u2_u14_u2_U32 (.A( u2_u14_u2_n156 ) , .B1( u2_u14_u2_n157 ) , .ZN( u2_u14_u2_n158 ) , .B2( u2_u14_u2_n179 ) );
  NOR2_X1 u2_u14_u2_U33 (.ZN( u2_u14_u2_n156 ) , .A1( u2_u14_u2_n166 ) , .A2( u2_u14_u2_n169 ) );
  NOR2_X1 u2_u14_u2_U34 (.A2( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n137 ) , .A1( u2_u14_u2_n140 ) );
  NOR2_X1 u2_u14_u2_U35 (.A2( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n153 ) , .A1( u2_u14_u2_n156 ) );
  AOI211_X1 u2_u14_u2_U36 (.ZN( u2_u14_u2_n130 ) , .C1( u2_u14_u2_n138 ) , .C2( u2_u14_u2_n179 ) , .B( u2_u14_u2_n96 ) , .A( u2_u14_u2_n97 ) );
  OAI22_X1 u2_u14_u2_U37 (.B1( u2_u14_u2_n133 ) , .A2( u2_u14_u2_n137 ) , .A1( u2_u14_u2_n152 ) , .B2( u2_u14_u2_n168 ) , .ZN( u2_u14_u2_n97 ) );
  OAI221_X1 u2_u14_u2_U38 (.B1( u2_u14_u2_n113 ) , .C1( u2_u14_u2_n132 ) , .A( u2_u14_u2_n149 ) , .B2( u2_u14_u2_n171 ) , .C2( u2_u14_u2_n172 ) , .ZN( u2_u14_u2_n96 ) );
  OAI221_X1 u2_u14_u2_U39 (.A( u2_u14_u2_n115 ) , .C2( u2_u14_u2_n123 ) , .B2( u2_u14_u2_n143 ) , .B1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n163 ) , .C1( u2_u14_u2_n168 ) );
  INV_X1 u2_u14_u2_U4 (.A( u2_u14_u2_n134 ) , .ZN( u2_u14_u2_n185 ) );
  OAI21_X1 u2_u14_u2_U40 (.A( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n115 ) , .B1( u2_u14_u2_n176 ) , .B2( u2_u14_u2_n178 ) );
  OAI221_X1 u2_u14_u2_U41 (.A( u2_u14_u2_n135 ) , .B2( u2_u14_u2_n136 ) , .B1( u2_u14_u2_n137 ) , .ZN( u2_u14_u2_n162 ) , .C2( u2_u14_u2_n167 ) , .C1( u2_u14_u2_n185 ) );
  AND3_X1 u2_u14_u2_U42 (.A3( u2_u14_u2_n131 ) , .A2( u2_u14_u2_n132 ) , .A1( u2_u14_u2_n133 ) , .ZN( u2_u14_u2_n136 ) );
  AOI22_X1 u2_u14_u2_U43 (.ZN( u2_u14_u2_n135 ) , .B1( u2_u14_u2_n140 ) , .A1( u2_u14_u2_n156 ) , .B2( u2_u14_u2_n180 ) , .A2( u2_u14_u2_n188 ) );
  AOI21_X1 u2_u14_u2_U44 (.ZN( u2_u14_u2_n149 ) , .B1( u2_u14_u2_n173 ) , .B2( u2_u14_u2_n188 ) , .A( u2_u14_u2_n95 ) );
  AND3_X1 u2_u14_u2_U45 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n156 ) , .ZN( u2_u14_u2_n95 ) );
  OAI21_X1 u2_u14_u2_U46 (.A( u2_u14_u2_n141 ) , .B2( u2_u14_u2_n142 ) , .ZN( u2_u14_u2_n146 ) , .B1( u2_u14_u2_n153 ) );
  OAI21_X1 u2_u14_u2_U47 (.A( u2_u14_u2_n140 ) , .ZN( u2_u14_u2_n141 ) , .B1( u2_u14_u2_n176 ) , .B2( u2_u14_u2_n177 ) );
  NOR3_X1 u2_u14_u2_U48 (.ZN( u2_u14_u2_n142 ) , .A3( u2_u14_u2_n175 ) , .A2( u2_u14_u2_n178 ) , .A1( u2_u14_u2_n181 ) );
  OAI21_X1 u2_u14_u2_U49 (.A( u2_u14_u2_n101 ) , .B2( u2_u14_u2_n121 ) , .B1( u2_u14_u2_n153 ) , .ZN( u2_u14_u2_n164 ) );
  INV_X1 u2_u14_u2_U5 (.A( u2_u14_u2_n150 ) , .ZN( u2_u14_u2_n184 ) );
  NAND2_X1 u2_u14_u2_U50 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n155 ) );
  NAND2_X1 u2_u14_u2_U51 (.A2( u2_u14_u2_n105 ) , .A1( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n143 ) );
  NAND2_X1 u2_u14_u2_U52 (.A1( u2_u14_u2_n104 ) , .A2( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n152 ) );
  NAND2_X1 u2_u14_u2_U53 (.A1( u2_u14_u2_n100 ) , .A2( u2_u14_u2_n105 ) , .ZN( u2_u14_u2_n132 ) );
  INV_X1 u2_u14_u2_U54 (.A( u2_u14_u2_n140 ) , .ZN( u2_u14_u2_n168 ) );
  INV_X1 u2_u14_u2_U55 (.A( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n167 ) );
  INV_X1 u2_u14_u2_U56 (.ZN( u2_u14_u2_n187 ) , .A( u2_u14_u2_n99 ) );
  OAI21_X1 u2_u14_u2_U57 (.B1( u2_u14_u2_n137 ) , .B2( u2_u14_u2_n143 ) , .A( u2_u14_u2_n98 ) , .ZN( u2_u14_u2_n99 ) );
  NAND2_X1 u2_u14_u2_U58 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n113 ) );
  NAND2_X1 u2_u14_u2_U59 (.A1( u2_u14_u2_n106 ) , .A2( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n131 ) );
  NOR4_X1 u2_u14_u2_U6 (.A4( u2_u14_u2_n124 ) , .A3( u2_u14_u2_n125 ) , .A2( u2_u14_u2_n126 ) , .A1( u2_u14_u2_n127 ) , .ZN( u2_u14_u2_n128 ) );
  NAND2_X1 u2_u14_u2_U60 (.A1( u2_u14_u2_n103 ) , .A2( u2_u14_u2_n107 ) , .ZN( u2_u14_u2_n139 ) );
  NAND2_X1 u2_u14_u2_U61 (.A1( u2_u14_u2_n103 ) , .A2( u2_u14_u2_n105 ) , .ZN( u2_u14_u2_n133 ) );
  NAND2_X1 u2_u14_u2_U62 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n103 ) , .ZN( u2_u14_u2_n154 ) );
  NAND2_X1 u2_u14_u2_U63 (.A2( u2_u14_u2_n103 ) , .A1( u2_u14_u2_n104 ) , .ZN( u2_u14_u2_n119 ) );
  NAND2_X1 u2_u14_u2_U64 (.A2( u2_u14_u2_n107 ) , .A1( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n123 ) );
  NAND2_X1 u2_u14_u2_U65 (.A1( u2_u14_u2_n104 ) , .A2( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n122 ) );
  INV_X1 u2_u14_u2_U66 (.A( u2_u14_u2_n114 ) , .ZN( u2_u14_u2_n172 ) );
  NAND2_X1 u2_u14_u2_U67 (.A2( u2_u14_u2_n100 ) , .A1( u2_u14_u2_n102 ) , .ZN( u2_u14_u2_n116 ) );
  NAND2_X1 u2_u14_u2_U68 (.A1( u2_u14_u2_n102 ) , .A2( u2_u14_u2_n108 ) , .ZN( u2_u14_u2_n120 ) );
  NAND2_X1 u2_u14_u2_U69 (.A2( u2_u14_u2_n105 ) , .A1( u2_u14_u2_n106 ) , .ZN( u2_u14_u2_n117 ) );
  AOI21_X1 u2_u14_u2_U7 (.B2( u2_u14_u2_n119 ) , .ZN( u2_u14_u2_n127 ) , .A( u2_u14_u2_n137 ) , .B1( u2_u14_u2_n155 ) );
  NOR2_X1 u2_u14_u2_U70 (.A2( u2_u14_X_16 ) , .ZN( u2_u14_u2_n140 ) , .A1( u2_u14_u2_n166 ) );
  NOR2_X1 u2_u14_u2_U71 (.A2( u2_u14_X_13 ) , .A1( u2_u14_X_14 ) , .ZN( u2_u14_u2_n100 ) );
  NOR2_X1 u2_u14_u2_U72 (.A2( u2_u14_X_16 ) , .A1( u2_u14_X_17 ) , .ZN( u2_u14_u2_n138 ) );
  NOR2_X1 u2_u14_u2_U73 (.A2( u2_u14_X_15 ) , .A1( u2_u14_X_18 ) , .ZN( u2_u14_u2_n104 ) );
  NOR2_X1 u2_u14_u2_U74 (.A2( u2_u14_X_14 ) , .ZN( u2_u14_u2_n103 ) , .A1( u2_u14_u2_n174 ) );
  NOR2_X1 u2_u14_u2_U75 (.A2( u2_u14_X_15 ) , .ZN( u2_u14_u2_n102 ) , .A1( u2_u14_u2_n165 ) );
  NOR2_X1 u2_u14_u2_U76 (.A2( u2_u14_X_17 ) , .ZN( u2_u14_u2_n114 ) , .A1( u2_u14_u2_n169 ) );
  AND2_X1 u2_u14_u2_U77 (.A1( u2_u14_X_15 ) , .ZN( u2_u14_u2_n105 ) , .A2( u2_u14_u2_n165 ) );
  AND2_X1 u2_u14_u2_U78 (.A2( u2_u14_X_15 ) , .A1( u2_u14_X_18 ) , .ZN( u2_u14_u2_n107 ) );
  AND2_X1 u2_u14_u2_U79 (.A1( u2_u14_X_14 ) , .ZN( u2_u14_u2_n106 ) , .A2( u2_u14_u2_n174 ) );
  AOI21_X1 u2_u14_u2_U8 (.ZN( u2_u14_u2_n124 ) , .B1( u2_u14_u2_n131 ) , .B2( u2_u14_u2_n143 ) , .A( u2_u14_u2_n172 ) );
  AND2_X1 u2_u14_u2_U80 (.A1( u2_u14_X_13 ) , .A2( u2_u14_X_14 ) , .ZN( u2_u14_u2_n108 ) );
  INV_X1 u2_u14_u2_U81 (.A( u2_u14_X_16 ) , .ZN( u2_u14_u2_n169 ) );
  INV_X1 u2_u14_u2_U82 (.A( u2_u14_X_17 ) , .ZN( u2_u14_u2_n166 ) );
  INV_X1 u2_u14_u2_U83 (.A( u2_u14_X_13 ) , .ZN( u2_u14_u2_n174 ) );
  INV_X1 u2_u14_u2_U84 (.A( u2_u14_X_18 ) , .ZN( u2_u14_u2_n165 ) );
  NAND4_X1 u2_u14_u2_U85 (.ZN( u2_out14_30 ) , .A4( u2_u14_u2_n147 ) , .A3( u2_u14_u2_n148 ) , .A2( u2_u14_u2_n149 ) , .A1( u2_u14_u2_n187 ) );
  NOR3_X1 u2_u14_u2_U86 (.A3( u2_u14_u2_n144 ) , .A2( u2_u14_u2_n145 ) , .A1( u2_u14_u2_n146 ) , .ZN( u2_u14_u2_n147 ) );
  AOI21_X1 u2_u14_u2_U87 (.B2( u2_u14_u2_n138 ) , .ZN( u2_u14_u2_n148 ) , .A( u2_u14_u2_n162 ) , .B1( u2_u14_u2_n182 ) );
  NAND4_X1 u2_u14_u2_U88 (.ZN( u2_out14_24 ) , .A4( u2_u14_u2_n111 ) , .A3( u2_u14_u2_n112 ) , .A1( u2_u14_u2_n130 ) , .A2( u2_u14_u2_n187 ) );
  AOI221_X1 u2_u14_u2_U89 (.A( u2_u14_u2_n109 ) , .B1( u2_u14_u2_n110 ) , .ZN( u2_u14_u2_n111 ) , .C1( u2_u14_u2_n134 ) , .C2( u2_u14_u2_n170 ) , .B2( u2_u14_u2_n173 ) );
  AOI21_X1 u2_u14_u2_U9 (.B2( u2_u14_u2_n123 ) , .ZN( u2_u14_u2_n125 ) , .A( u2_u14_u2_n171 ) , .B1( u2_u14_u2_n184 ) );
  AOI21_X1 u2_u14_u2_U90 (.ZN( u2_u14_u2_n112 ) , .B2( u2_u14_u2_n156 ) , .A( u2_u14_u2_n164 ) , .B1( u2_u14_u2_n181 ) );
  NAND4_X1 u2_u14_u2_U91 (.ZN( u2_out14_16 ) , .A4( u2_u14_u2_n128 ) , .A3( u2_u14_u2_n129 ) , .A1( u2_u14_u2_n130 ) , .A2( u2_u14_u2_n186 ) );
  AOI22_X1 u2_u14_u2_U92 (.A2( u2_u14_u2_n118 ) , .ZN( u2_u14_u2_n129 ) , .A1( u2_u14_u2_n140 ) , .B1( u2_u14_u2_n157 ) , .B2( u2_u14_u2_n170 ) );
  INV_X1 u2_u14_u2_U93 (.A( u2_u14_u2_n163 ) , .ZN( u2_u14_u2_n186 ) );
  OR4_X1 u2_u14_u2_U94 (.ZN( u2_out14_6 ) , .A4( u2_u14_u2_n161 ) , .A3( u2_u14_u2_n162 ) , .A2( u2_u14_u2_n163 ) , .A1( u2_u14_u2_n164 ) );
  OR3_X1 u2_u14_u2_U95 (.A2( u2_u14_u2_n159 ) , .A1( u2_u14_u2_n160 ) , .ZN( u2_u14_u2_n161 ) , .A3( u2_u14_u2_n183 ) );
  AOI21_X1 u2_u14_u2_U96 (.B2( u2_u14_u2_n154 ) , .B1( u2_u14_u2_n155 ) , .ZN( u2_u14_u2_n159 ) , .A( u2_u14_u2_n167 ) );
  NAND3_X1 u2_u14_u2_U97 (.A2( u2_u14_u2_n117 ) , .A1( u2_u14_u2_n122 ) , .A3( u2_u14_u2_n123 ) , .ZN( u2_u14_u2_n134 ) );
  NAND3_X1 u2_u14_u2_U98 (.ZN( u2_u14_u2_n110 ) , .A2( u2_u14_u2_n131 ) , .A3( u2_u14_u2_n139 ) , .A1( u2_u14_u2_n154 ) );
  NAND3_X1 u2_u14_u2_U99 (.A2( u2_u14_u2_n100 ) , .ZN( u2_u14_u2_n101 ) , .A1( u2_u14_u2_n104 ) , .A3( u2_u14_u2_n114 ) );
  OAI22_X1 u2_u14_u3_U10 (.B1( u2_u14_u3_n113 ) , .A2( u2_u14_u3_n135 ) , .A1( u2_u14_u3_n150 ) , .B2( u2_u14_u3_n164 ) , .ZN( u2_u14_u3_n98 ) );
  OAI211_X1 u2_u14_u3_U11 (.B( u2_u14_u3_n106 ) , .ZN( u2_u14_u3_n119 ) , .C2( u2_u14_u3_n128 ) , .C1( u2_u14_u3_n167 ) , .A( u2_u14_u3_n181 ) );
  AOI221_X1 u2_u14_u3_U12 (.C1( u2_u14_u3_n105 ) , .ZN( u2_u14_u3_n106 ) , .A( u2_u14_u3_n131 ) , .B2( u2_u14_u3_n132 ) , .C2( u2_u14_u3_n133 ) , .B1( u2_u14_u3_n169 ) );
  INV_X1 u2_u14_u3_U13 (.ZN( u2_u14_u3_n181 ) , .A( u2_u14_u3_n98 ) );
  NAND2_X1 u2_u14_u3_U14 (.ZN( u2_u14_u3_n105 ) , .A2( u2_u14_u3_n130 ) , .A1( u2_u14_u3_n155 ) );
  AOI22_X1 u2_u14_u3_U15 (.B1( u2_u14_u3_n115 ) , .A2( u2_u14_u3_n116 ) , .ZN( u2_u14_u3_n123 ) , .B2( u2_u14_u3_n133 ) , .A1( u2_u14_u3_n169 ) );
  NAND2_X1 u2_u14_u3_U16 (.ZN( u2_u14_u3_n116 ) , .A2( u2_u14_u3_n151 ) , .A1( u2_u14_u3_n182 ) );
  NOR2_X1 u2_u14_u3_U17 (.ZN( u2_u14_u3_n126 ) , .A2( u2_u14_u3_n150 ) , .A1( u2_u14_u3_n164 ) );
  AOI21_X1 u2_u14_u3_U18 (.ZN( u2_u14_u3_n112 ) , .B2( u2_u14_u3_n146 ) , .B1( u2_u14_u3_n155 ) , .A( u2_u14_u3_n167 ) );
  NAND2_X1 u2_u14_u3_U19 (.A1( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n142 ) , .A2( u2_u14_u3_n164 ) );
  NAND2_X1 u2_u14_u3_U20 (.ZN( u2_u14_u3_n132 ) , .A2( u2_u14_u3_n152 ) , .A1( u2_u14_u3_n156 ) );
  AND2_X1 u2_u14_u3_U21 (.A2( u2_u14_u3_n113 ) , .A1( u2_u14_u3_n114 ) , .ZN( u2_u14_u3_n151 ) );
  INV_X1 u2_u14_u3_U22 (.A( u2_u14_u3_n133 ) , .ZN( u2_u14_u3_n165 ) );
  INV_X1 u2_u14_u3_U23 (.A( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n170 ) );
  NAND2_X1 u2_u14_u3_U24 (.A1( u2_u14_u3_n107 ) , .A2( u2_u14_u3_n108 ) , .ZN( u2_u14_u3_n140 ) );
  NAND2_X1 u2_u14_u3_U25 (.ZN( u2_u14_u3_n117 ) , .A1( u2_u14_u3_n124 ) , .A2( u2_u14_u3_n148 ) );
  NAND2_X1 u2_u14_u3_U26 (.ZN( u2_u14_u3_n143 ) , .A1( u2_u14_u3_n165 ) , .A2( u2_u14_u3_n167 ) );
  INV_X1 u2_u14_u3_U27 (.A( u2_u14_u3_n130 ) , .ZN( u2_u14_u3_n177 ) );
  INV_X1 u2_u14_u3_U28 (.A( u2_u14_u3_n128 ) , .ZN( u2_u14_u3_n176 ) );
  INV_X1 u2_u14_u3_U29 (.A( u2_u14_u3_n155 ) , .ZN( u2_u14_u3_n174 ) );
  INV_X1 u2_u14_u3_U3 (.A( u2_u14_u3_n129 ) , .ZN( u2_u14_u3_n183 ) );
  INV_X1 u2_u14_u3_U30 (.A( u2_u14_u3_n139 ) , .ZN( u2_u14_u3_n185 ) );
  NOR2_X1 u2_u14_u3_U31 (.ZN( u2_u14_u3_n135 ) , .A2( u2_u14_u3_n141 ) , .A1( u2_u14_u3_n169 ) );
  OAI222_X1 u2_u14_u3_U32 (.C2( u2_u14_u3_n107 ) , .A2( u2_u14_u3_n108 ) , .B1( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n138 ) , .B2( u2_u14_u3_n146 ) , .C1( u2_u14_u3_n154 ) , .A1( u2_u14_u3_n164 ) );
  NOR4_X1 u2_u14_u3_U33 (.A4( u2_u14_u3_n157 ) , .A3( u2_u14_u3_n158 ) , .A2( u2_u14_u3_n159 ) , .A1( u2_u14_u3_n160 ) , .ZN( u2_u14_u3_n161 ) );
  AOI21_X1 u2_u14_u3_U34 (.B2( u2_u14_u3_n152 ) , .B1( u2_u14_u3_n153 ) , .ZN( u2_u14_u3_n158 ) , .A( u2_u14_u3_n164 ) );
  AOI21_X1 u2_u14_u3_U35 (.A( u2_u14_u3_n154 ) , .B2( u2_u14_u3_n155 ) , .B1( u2_u14_u3_n156 ) , .ZN( u2_u14_u3_n157 ) );
  AOI21_X1 u2_u14_u3_U36 (.A( u2_u14_u3_n149 ) , .B2( u2_u14_u3_n150 ) , .B1( u2_u14_u3_n151 ) , .ZN( u2_u14_u3_n159 ) );
  AOI211_X1 u2_u14_u3_U37 (.ZN( u2_u14_u3_n109 ) , .A( u2_u14_u3_n119 ) , .C2( u2_u14_u3_n129 ) , .B( u2_u14_u3_n138 ) , .C1( u2_u14_u3_n141 ) );
  AOI211_X1 u2_u14_u3_U38 (.B( u2_u14_u3_n119 ) , .A( u2_u14_u3_n120 ) , .C2( u2_u14_u3_n121 ) , .ZN( u2_u14_u3_n122 ) , .C1( u2_u14_u3_n179 ) );
  INV_X1 u2_u14_u3_U39 (.A( u2_u14_u3_n156 ) , .ZN( u2_u14_u3_n179 ) );
  INV_X1 u2_u14_u3_U4 (.A( u2_u14_u3_n140 ) , .ZN( u2_u14_u3_n182 ) );
  OAI22_X1 u2_u14_u3_U40 (.B1( u2_u14_u3_n118 ) , .ZN( u2_u14_u3_n120 ) , .A1( u2_u14_u3_n135 ) , .B2( u2_u14_u3_n154 ) , .A2( u2_u14_u3_n178 ) );
  AND3_X1 u2_u14_u3_U41 (.ZN( u2_u14_u3_n118 ) , .A2( u2_u14_u3_n124 ) , .A1( u2_u14_u3_n144 ) , .A3( u2_u14_u3_n152 ) );
  INV_X1 u2_u14_u3_U42 (.A( u2_u14_u3_n121 ) , .ZN( u2_u14_u3_n164 ) );
  NAND2_X1 u2_u14_u3_U43 (.ZN( u2_u14_u3_n133 ) , .A1( u2_u14_u3_n154 ) , .A2( u2_u14_u3_n164 ) );
  OAI211_X1 u2_u14_u3_U44 (.B( u2_u14_u3_n127 ) , .ZN( u2_u14_u3_n139 ) , .C1( u2_u14_u3_n150 ) , .C2( u2_u14_u3_n154 ) , .A( u2_u14_u3_n184 ) );
  INV_X1 u2_u14_u3_U45 (.A( u2_u14_u3_n125 ) , .ZN( u2_u14_u3_n184 ) );
  AOI221_X1 u2_u14_u3_U46 (.A( u2_u14_u3_n126 ) , .ZN( u2_u14_u3_n127 ) , .C2( u2_u14_u3_n132 ) , .C1( u2_u14_u3_n169 ) , .B2( u2_u14_u3_n170 ) , .B1( u2_u14_u3_n174 ) );
  OAI22_X1 u2_u14_u3_U47 (.A1( u2_u14_u3_n124 ) , .ZN( u2_u14_u3_n125 ) , .B2( u2_u14_u3_n145 ) , .A2( u2_u14_u3_n165 ) , .B1( u2_u14_u3_n167 ) );
  NOR2_X1 u2_u14_u3_U48 (.A1( u2_u14_u3_n113 ) , .ZN( u2_u14_u3_n131 ) , .A2( u2_u14_u3_n154 ) );
  NAND2_X1 u2_u14_u3_U49 (.A1( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n150 ) , .A2( u2_u14_u3_n99 ) );
  INV_X1 u2_u14_u3_U5 (.A( u2_u14_u3_n117 ) , .ZN( u2_u14_u3_n178 ) );
  NAND2_X1 u2_u14_u3_U50 (.A2( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n155 ) , .A1( u2_u14_u3_n97 ) );
  INV_X1 u2_u14_u3_U51 (.A( u2_u14_u3_n141 ) , .ZN( u2_u14_u3_n167 ) );
  AOI21_X1 u2_u14_u3_U52 (.B2( u2_u14_u3_n114 ) , .B1( u2_u14_u3_n146 ) , .A( u2_u14_u3_n154 ) , .ZN( u2_u14_u3_n94 ) );
  AOI21_X1 u2_u14_u3_U53 (.ZN( u2_u14_u3_n110 ) , .B2( u2_u14_u3_n142 ) , .B1( u2_u14_u3_n186 ) , .A( u2_u14_u3_n95 ) );
  INV_X1 u2_u14_u3_U54 (.A( u2_u14_u3_n145 ) , .ZN( u2_u14_u3_n186 ) );
  AOI21_X1 u2_u14_u3_U55 (.B1( u2_u14_u3_n124 ) , .A( u2_u14_u3_n149 ) , .B2( u2_u14_u3_n155 ) , .ZN( u2_u14_u3_n95 ) );
  INV_X1 u2_u14_u3_U56 (.A( u2_u14_u3_n149 ) , .ZN( u2_u14_u3_n169 ) );
  NAND2_X1 u2_u14_u3_U57 (.ZN( u2_u14_u3_n124 ) , .A1( u2_u14_u3_n96 ) , .A2( u2_u14_u3_n97 ) );
  NAND2_X1 u2_u14_u3_U58 (.A2( u2_u14_u3_n100 ) , .ZN( u2_u14_u3_n146 ) , .A1( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U59 (.A1( u2_u14_u3_n101 ) , .ZN( u2_u14_u3_n145 ) , .A2( u2_u14_u3_n99 ) );
  AOI221_X1 u2_u14_u3_U6 (.A( u2_u14_u3_n131 ) , .C2( u2_u14_u3_n132 ) , .C1( u2_u14_u3_n133 ) , .ZN( u2_u14_u3_n134 ) , .B1( u2_u14_u3_n143 ) , .B2( u2_u14_u3_n177 ) );
  NAND2_X1 u2_u14_u3_U60 (.A1( u2_u14_u3_n100 ) , .ZN( u2_u14_u3_n156 ) , .A2( u2_u14_u3_n99 ) );
  NAND2_X1 u2_u14_u3_U61 (.A2( u2_u14_u3_n101 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n148 ) );
  NAND2_X1 u2_u14_u3_U62 (.A1( u2_u14_u3_n100 ) , .A2( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n128 ) );
  NAND2_X1 u2_u14_u3_U63 (.A2( u2_u14_u3_n101 ) , .A1( u2_u14_u3_n102 ) , .ZN( u2_u14_u3_n152 ) );
  NAND2_X1 u2_u14_u3_U64 (.A2( u2_u14_u3_n101 ) , .ZN( u2_u14_u3_n114 ) , .A1( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U65 (.ZN( u2_u14_u3_n107 ) , .A1( u2_u14_u3_n97 ) , .A2( u2_u14_u3_n99 ) );
  NAND2_X1 u2_u14_u3_U66 (.A2( u2_u14_u3_n100 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n113 ) );
  NAND2_X1 u2_u14_u3_U67 (.A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n153 ) , .A2( u2_u14_u3_n97 ) );
  NAND2_X1 u2_u14_u3_U68 (.A2( u2_u14_u3_n103 ) , .A1( u2_u14_u3_n104 ) , .ZN( u2_u14_u3_n130 ) );
  NAND2_X1 u2_u14_u3_U69 (.A2( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n144 ) , .A1( u2_u14_u3_n96 ) );
  OAI22_X1 u2_u14_u3_U7 (.B2( u2_u14_u3_n147 ) , .A2( u2_u14_u3_n148 ) , .ZN( u2_u14_u3_n160 ) , .B1( u2_u14_u3_n165 ) , .A1( u2_u14_u3_n168 ) );
  NAND2_X1 u2_u14_u3_U70 (.A1( u2_u14_u3_n102 ) , .A2( u2_u14_u3_n103 ) , .ZN( u2_u14_u3_n108 ) );
  NOR2_X1 u2_u14_u3_U71 (.A2( u2_u14_X_19 ) , .A1( u2_u14_X_20 ) , .ZN( u2_u14_u3_n99 ) );
  NOR2_X1 u2_u14_u3_U72 (.A2( u2_u14_X_21 ) , .A1( u2_u14_X_24 ) , .ZN( u2_u14_u3_n103 ) );
  NOR2_X1 u2_u14_u3_U73 (.A2( u2_u14_X_24 ) , .A1( u2_u14_u3_n171 ) , .ZN( u2_u14_u3_n97 ) );
  NOR2_X1 u2_u14_u3_U74 (.A2( u2_u14_X_23 ) , .ZN( u2_u14_u3_n141 ) , .A1( u2_u14_u3_n166 ) );
  NOR2_X1 u2_u14_u3_U75 (.A2( u2_u14_X_19 ) , .A1( u2_u14_u3_n172 ) , .ZN( u2_u14_u3_n96 ) );
  NAND2_X1 u2_u14_u3_U76 (.A1( u2_u14_X_22 ) , .A2( u2_u14_X_23 ) , .ZN( u2_u14_u3_n154 ) );
  NAND2_X1 u2_u14_u3_U77 (.A1( u2_u14_X_23 ) , .ZN( u2_u14_u3_n149 ) , .A2( u2_u14_u3_n166 ) );
  NOR2_X1 u2_u14_u3_U78 (.A2( u2_u14_X_22 ) , .A1( u2_u14_X_23 ) , .ZN( u2_u14_u3_n121 ) );
  AND2_X1 u2_u14_u3_U79 (.A1( u2_u14_X_24 ) , .ZN( u2_u14_u3_n101 ) , .A2( u2_u14_u3_n171 ) );
  AND3_X1 u2_u14_u3_U8 (.A3( u2_u14_u3_n144 ) , .A2( u2_u14_u3_n145 ) , .A1( u2_u14_u3_n146 ) , .ZN( u2_u14_u3_n147 ) );
  AND2_X1 u2_u14_u3_U80 (.A1( u2_u14_X_19 ) , .ZN( u2_u14_u3_n102 ) , .A2( u2_u14_u3_n172 ) );
  AND2_X1 u2_u14_u3_U81 (.A1( u2_u14_X_21 ) , .A2( u2_u14_X_24 ) , .ZN( u2_u14_u3_n100 ) );
  AND2_X1 u2_u14_u3_U82 (.A2( u2_u14_X_19 ) , .A1( u2_u14_X_20 ) , .ZN( u2_u14_u3_n104 ) );
  INV_X1 u2_u14_u3_U83 (.A( u2_u14_X_22 ) , .ZN( u2_u14_u3_n166 ) );
  INV_X1 u2_u14_u3_U84 (.A( u2_u14_X_21 ) , .ZN( u2_u14_u3_n171 ) );
  INV_X1 u2_u14_u3_U85 (.A( u2_u14_X_20 ) , .ZN( u2_u14_u3_n172 ) );
  NAND4_X1 u2_u14_u3_U86 (.ZN( u2_out14_26 ) , .A4( u2_u14_u3_n109 ) , .A3( u2_u14_u3_n110 ) , .A2( u2_u14_u3_n111 ) , .A1( u2_u14_u3_n173 ) );
  INV_X1 u2_u14_u3_U87 (.ZN( u2_u14_u3_n173 ) , .A( u2_u14_u3_n94 ) );
  OAI21_X1 u2_u14_u3_U88 (.ZN( u2_u14_u3_n111 ) , .B2( u2_u14_u3_n117 ) , .A( u2_u14_u3_n133 ) , .B1( u2_u14_u3_n176 ) );
  NAND4_X1 u2_u14_u3_U89 (.ZN( u2_out14_20 ) , .A4( u2_u14_u3_n122 ) , .A3( u2_u14_u3_n123 ) , .A1( u2_u14_u3_n175 ) , .A2( u2_u14_u3_n180 ) );
  INV_X1 u2_u14_u3_U9 (.A( u2_u14_u3_n143 ) , .ZN( u2_u14_u3_n168 ) );
  INV_X1 u2_u14_u3_U90 (.A( u2_u14_u3_n126 ) , .ZN( u2_u14_u3_n180 ) );
  INV_X1 u2_u14_u3_U91 (.A( u2_u14_u3_n112 ) , .ZN( u2_u14_u3_n175 ) );
  NAND4_X1 u2_u14_u3_U92 (.ZN( u2_out14_1 ) , .A4( u2_u14_u3_n161 ) , .A3( u2_u14_u3_n162 ) , .A2( u2_u14_u3_n163 ) , .A1( u2_u14_u3_n185 ) );
  NAND2_X1 u2_u14_u3_U93 (.ZN( u2_u14_u3_n163 ) , .A2( u2_u14_u3_n170 ) , .A1( u2_u14_u3_n176 ) );
  AOI22_X1 u2_u14_u3_U94 (.B2( u2_u14_u3_n140 ) , .B1( u2_u14_u3_n141 ) , .A2( u2_u14_u3_n142 ) , .ZN( u2_u14_u3_n162 ) , .A1( u2_u14_u3_n177 ) );
  OR4_X1 u2_u14_u3_U95 (.ZN( u2_out14_10 ) , .A4( u2_u14_u3_n136 ) , .A3( u2_u14_u3_n137 ) , .A1( u2_u14_u3_n138 ) , .A2( u2_u14_u3_n139 ) );
  OAI222_X1 u2_u14_u3_U96 (.C1( u2_u14_u3_n128 ) , .ZN( u2_u14_u3_n137 ) , .B1( u2_u14_u3_n148 ) , .A2( u2_u14_u3_n150 ) , .B2( u2_u14_u3_n154 ) , .C2( u2_u14_u3_n164 ) , .A1( u2_u14_u3_n167 ) );
  OAI221_X1 u2_u14_u3_U97 (.A( u2_u14_u3_n134 ) , .B2( u2_u14_u3_n135 ) , .ZN( u2_u14_u3_n136 ) , .C1( u2_u14_u3_n149 ) , .B1( u2_u14_u3_n151 ) , .C2( u2_u14_u3_n183 ) );
  NAND3_X1 u2_u14_u3_U98 (.A1( u2_u14_u3_n114 ) , .ZN( u2_u14_u3_n115 ) , .A2( u2_u14_u3_n145 ) , .A3( u2_u14_u3_n153 ) );
  NAND3_X1 u2_u14_u3_U99 (.ZN( u2_u14_u3_n129 ) , .A2( u2_u14_u3_n144 ) , .A1( u2_u14_u3_n153 ) , .A3( u2_u14_u3_n182 ) );
  OAI21_X1 u2_u14_u7_U10 (.A( u2_u14_u7_n161 ) , .B1( u2_u14_u7_n168 ) , .B2( u2_u14_u7_n173 ) , .ZN( u2_u14_u7_n91 ) );
  AOI211_X1 u2_u14_u7_U11 (.A( u2_u14_u7_n117 ) , .ZN( u2_u14_u7_n118 ) , .C2( u2_u14_u7_n126 ) , .C1( u2_u14_u7_n177 ) , .B( u2_u14_u7_n180 ) );
  OAI22_X1 u2_u14_u7_U12 (.B1( u2_u14_u7_n115 ) , .ZN( u2_u14_u7_n117 ) , .A2( u2_u14_u7_n133 ) , .A1( u2_u14_u7_n137 ) , .B2( u2_u14_u7_n162 ) );
  INV_X1 u2_u14_u7_U13 (.A( u2_u14_u7_n116 ) , .ZN( u2_u14_u7_n180 ) );
  NOR3_X1 u2_u14_u7_U14 (.ZN( u2_u14_u7_n115 ) , .A3( u2_u14_u7_n145 ) , .A2( u2_u14_u7_n168 ) , .A1( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U15 (.A( u2_u14_u7_n133 ) , .ZN( u2_u14_u7_n176 ) );
  NOR3_X1 u2_u14_u7_U16 (.A2( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n135 ) , .ZN( u2_u14_u7_n136 ) , .A3( u2_u14_u7_n171 ) );
  NOR2_X1 u2_u14_u7_U17 (.A1( u2_u14_u7_n130 ) , .A2( u2_u14_u7_n134 ) , .ZN( u2_u14_u7_n153 ) );
  AOI21_X1 u2_u14_u7_U18 (.ZN( u2_u14_u7_n104 ) , .B2( u2_u14_u7_n112 ) , .B1( u2_u14_u7_n127 ) , .A( u2_u14_u7_n164 ) );
  AOI21_X1 u2_u14_u7_U19 (.ZN( u2_u14_u7_n106 ) , .B1( u2_u14_u7_n133 ) , .B2( u2_u14_u7_n146 ) , .A( u2_u14_u7_n162 ) );
  AOI21_X1 u2_u14_u7_U20 (.A( u2_u14_u7_n101 ) , .ZN( u2_u14_u7_n107 ) , .B2( u2_u14_u7_n128 ) , .B1( u2_u14_u7_n175 ) );
  INV_X1 u2_u14_u7_U21 (.A( u2_u14_u7_n101 ) , .ZN( u2_u14_u7_n165 ) );
  NOR2_X1 u2_u14_u7_U22 (.ZN( u2_u14_u7_n111 ) , .A2( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U23 (.A( u2_u14_u7_n138 ) , .ZN( u2_u14_u7_n171 ) );
  INV_X1 u2_u14_u7_U24 (.A( u2_u14_u7_n131 ) , .ZN( u2_u14_u7_n177 ) );
  INV_X1 u2_u14_u7_U25 (.A( u2_u14_u7_n110 ) , .ZN( u2_u14_u7_n174 ) );
  NAND2_X1 u2_u14_u7_U26 (.A1( u2_u14_u7_n129 ) , .A2( u2_u14_u7_n132 ) , .ZN( u2_u14_u7_n149 ) );
  NAND2_X1 u2_u14_u7_U27 (.A1( u2_u14_u7_n113 ) , .A2( u2_u14_u7_n124 ) , .ZN( u2_u14_u7_n130 ) );
  INV_X1 u2_u14_u7_U28 (.A( u2_u14_u7_n112 ) , .ZN( u2_u14_u7_n173 ) );
  INV_X1 u2_u14_u7_U29 (.A( u2_u14_u7_n128 ) , .ZN( u2_u14_u7_n168 ) );
  OAI21_X1 u2_u14_u7_U3 (.ZN( u2_u14_u7_n159 ) , .A( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n171 ) , .B1( u2_u14_u7_n174 ) );
  INV_X1 u2_u14_u7_U30 (.A( u2_u14_u7_n148 ) , .ZN( u2_u14_u7_n169 ) );
  INV_X1 u2_u14_u7_U31 (.A( u2_u14_u7_n127 ) , .ZN( u2_u14_u7_n179 ) );
  NOR2_X1 u2_u14_u7_U32 (.ZN( u2_u14_u7_n101 ) , .A2( u2_u14_u7_n150 ) , .A1( u2_u14_u7_n156 ) );
  AOI211_X1 u2_u14_u7_U33 (.B( u2_u14_u7_n139 ) , .A( u2_u14_u7_n140 ) , .C2( u2_u14_u7_n141 ) , .ZN( u2_u14_u7_n142 ) , .C1( u2_u14_u7_n156 ) );
  NAND4_X1 u2_u14_u7_U34 (.A3( u2_u14_u7_n127 ) , .A2( u2_u14_u7_n128 ) , .A1( u2_u14_u7_n129 ) , .ZN( u2_u14_u7_n141 ) , .A4( u2_u14_u7_n147 ) );
  AOI21_X1 u2_u14_u7_U35 (.A( u2_u14_u7_n137 ) , .B1( u2_u14_u7_n138 ) , .ZN( u2_u14_u7_n139 ) , .B2( u2_u14_u7_n146 ) );
  OAI22_X1 u2_u14_u7_U36 (.B1( u2_u14_u7_n136 ) , .ZN( u2_u14_u7_n140 ) , .A1( u2_u14_u7_n153 ) , .B2( u2_u14_u7_n162 ) , .A2( u2_u14_u7_n164 ) );
  INV_X1 u2_u14_u7_U37 (.A( u2_u14_u7_n125 ) , .ZN( u2_u14_u7_n161 ) );
  AOI21_X1 u2_u14_u7_U38 (.ZN( u2_u14_u7_n123 ) , .B1( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n177 ) , .A( u2_u14_u7_n97 ) );
  AOI21_X1 u2_u14_u7_U39 (.B2( u2_u14_u7_n113 ) , .B1( u2_u14_u7_n124 ) , .A( u2_u14_u7_n125 ) , .ZN( u2_u14_u7_n97 ) );
  INV_X1 u2_u14_u7_U4 (.A( u2_u14_u7_n149 ) , .ZN( u2_u14_u7_n175 ) );
  INV_X1 u2_u14_u7_U40 (.A( u2_u14_u7_n152 ) , .ZN( u2_u14_u7_n162 ) );
  AOI22_X1 u2_u14_u7_U41 (.A2( u2_u14_u7_n114 ) , .ZN( u2_u14_u7_n119 ) , .B1( u2_u14_u7_n130 ) , .A1( u2_u14_u7_n156 ) , .B2( u2_u14_u7_n165 ) );
  NAND2_X1 u2_u14_u7_U42 (.A2( u2_u14_u7_n112 ) , .ZN( u2_u14_u7_n114 ) , .A1( u2_u14_u7_n175 ) );
  NOR2_X1 u2_u14_u7_U43 (.ZN( u2_u14_u7_n137 ) , .A1( u2_u14_u7_n150 ) , .A2( u2_u14_u7_n161 ) );
  AND2_X1 u2_u14_u7_U44 (.ZN( u2_u14_u7_n145 ) , .A2( u2_u14_u7_n98 ) , .A1( u2_u14_u7_n99 ) );
  AOI21_X1 u2_u14_u7_U45 (.ZN( u2_u14_u7_n105 ) , .B2( u2_u14_u7_n110 ) , .A( u2_u14_u7_n125 ) , .B1( u2_u14_u7_n147 ) );
  NAND2_X1 u2_u14_u7_U46 (.ZN( u2_u14_u7_n146 ) , .A1( u2_u14_u7_n95 ) , .A2( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U47 (.A2( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n147 ) , .A1( u2_u14_u7_n93 ) );
  NAND2_X1 u2_u14_u7_U48 (.A1( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n127 ) , .A2( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U49 (.A2( u2_u14_u7_n102 ) , .A1( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n133 ) );
  INV_X1 u2_u14_u7_U5 (.A( u2_u14_u7_n154 ) , .ZN( u2_u14_u7_n178 ) );
  OR2_X1 u2_u14_u7_U50 (.ZN( u2_u14_u7_n126 ) , .A2( u2_u14_u7_n152 ) , .A1( u2_u14_u7_n156 ) );
  NAND2_X1 u2_u14_u7_U51 (.ZN( u2_u14_u7_n112 ) , .A2( u2_u14_u7_n96 ) , .A1( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U52 (.A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n128 ) , .A1( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U53 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n113 ) , .A2( u2_u14_u7_n93 ) );
  NAND2_X1 u2_u14_u7_U54 (.ZN( u2_u14_u7_n110 ) , .A1( u2_u14_u7_n95 ) , .A2( u2_u14_u7_n96 ) );
  INV_X1 u2_u14_u7_U55 (.A( u2_u14_u7_n150 ) , .ZN( u2_u14_u7_n164 ) );
  AND2_X1 u2_u14_u7_U56 (.ZN( u2_u14_u7_n134 ) , .A1( u2_u14_u7_n93 ) , .A2( u2_u14_u7_n98 ) );
  NAND2_X1 u2_u14_u7_U57 (.A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n124 ) , .A1( u2_u14_u7_n96 ) );
  NAND2_X1 u2_u14_u7_U58 (.A1( u2_u14_u7_n100 ) , .A2( u2_u14_u7_n102 ) , .ZN( u2_u14_u7_n129 ) );
  NAND2_X1 u2_u14_u7_U59 (.A2( u2_u14_u7_n103 ) , .ZN( u2_u14_u7_n131 ) , .A1( u2_u14_u7_n95 ) );
  AOI211_X1 u2_u14_u7_U6 (.ZN( u2_u14_u7_n116 ) , .A( u2_u14_u7_n155 ) , .C1( u2_u14_u7_n161 ) , .C2( u2_u14_u7_n171 ) , .B( u2_u14_u7_n94 ) );
  NAND2_X1 u2_u14_u7_U60 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n138 ) , .A2( u2_u14_u7_n99 ) );
  NAND2_X1 u2_u14_u7_U61 (.ZN( u2_u14_u7_n132 ) , .A1( u2_u14_u7_n93 ) , .A2( u2_u14_u7_n96 ) );
  NAND2_X1 u2_u14_u7_U62 (.A1( u2_u14_u7_n100 ) , .ZN( u2_u14_u7_n148 ) , .A2( u2_u14_u7_n95 ) );
  AOI211_X1 u2_u14_u7_U63 (.B( u2_u14_u7_n154 ) , .A( u2_u14_u7_n155 ) , .C1( u2_u14_u7_n156 ) , .ZN( u2_u14_u7_n157 ) , .C2( u2_u14_u7_n172 ) );
  INV_X1 u2_u14_u7_U64 (.A( u2_u14_u7_n153 ) , .ZN( u2_u14_u7_n172 ) );
  NOR2_X1 u2_u14_u7_U65 (.A2( u2_u14_X_47 ) , .ZN( u2_u14_u7_n150 ) , .A1( u2_u14_u7_n163 ) );
  NOR2_X1 u2_u14_u7_U66 (.A2( u2_u14_X_43 ) , .A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n103 ) );
  NOR2_X1 u2_u14_u7_U67 (.A2( u2_u14_X_48 ) , .A1( u2_u14_u7_n166 ) , .ZN( u2_u14_u7_n95 ) );
  NOR2_X1 u2_u14_u7_U68 (.A2( u2_u14_X_45 ) , .A1( u2_u14_X_48 ) , .ZN( u2_u14_u7_n99 ) );
  NOR2_X1 u2_u14_u7_U69 (.A2( u2_u14_X_44 ) , .A1( u2_u14_u7_n167 ) , .ZN( u2_u14_u7_n98 ) );
  OAI222_X1 u2_u14_u7_U7 (.C2( u2_u14_u7_n101 ) , .B2( u2_u14_u7_n111 ) , .A1( u2_u14_u7_n113 ) , .C1( u2_u14_u7_n146 ) , .A2( u2_u14_u7_n162 ) , .B1( u2_u14_u7_n164 ) , .ZN( u2_u14_u7_n94 ) );
  NOR2_X1 u2_u14_u7_U70 (.A2( u2_u14_X_46 ) , .A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n152 ) );
  NAND2_X1 u2_u14_u7_U71 (.A2( u2_u14_X_46 ) , .A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n125 ) );
  AND2_X1 u2_u14_u7_U72 (.A1( u2_u14_X_47 ) , .ZN( u2_u14_u7_n156 ) , .A2( u2_u14_u7_n163 ) );
  AND2_X1 u2_u14_u7_U73 (.A2( u2_u14_X_45 ) , .A1( u2_u14_X_48 ) , .ZN( u2_u14_u7_n102 ) );
  AND2_X1 u2_u14_u7_U74 (.A2( u2_u14_X_43 ) , .A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n96 ) );
  AND2_X1 u2_u14_u7_U75 (.A1( u2_u14_X_44 ) , .ZN( u2_u14_u7_n100 ) , .A2( u2_u14_u7_n167 ) );
  AND2_X1 u2_u14_u7_U76 (.A1( u2_u14_X_48 ) , .A2( u2_u14_u7_n166 ) , .ZN( u2_u14_u7_n93 ) );
  INV_X1 u2_u14_u7_U77 (.A( u2_u14_X_46 ) , .ZN( u2_u14_u7_n163 ) );
  INV_X1 u2_u14_u7_U78 (.A( u2_u14_X_45 ) , .ZN( u2_u14_u7_n166 ) );
  INV_X1 u2_u14_u7_U79 (.A( u2_u14_X_43 ) , .ZN( u2_u14_u7_n167 ) );
  OAI221_X1 u2_u14_u7_U8 (.C1( u2_u14_u7_n101 ) , .C2( u2_u14_u7_n147 ) , .ZN( u2_u14_u7_n155 ) , .B2( u2_u14_u7_n162 ) , .A( u2_u14_u7_n91 ) , .B1( u2_u14_u7_n92 ) );
  NAND4_X1 u2_u14_u7_U80 (.ZN( u2_out14_27 ) , .A4( u2_u14_u7_n118 ) , .A3( u2_u14_u7_n119 ) , .A2( u2_u14_u7_n120 ) , .A1( u2_u14_u7_n121 ) );
  OAI21_X1 u2_u14_u7_U81 (.ZN( u2_u14_u7_n121 ) , .B2( u2_u14_u7_n145 ) , .A( u2_u14_u7_n150 ) , .B1( u2_u14_u7_n174 ) );
  OAI21_X1 u2_u14_u7_U82 (.ZN( u2_u14_u7_n120 ) , .A( u2_u14_u7_n161 ) , .B2( u2_u14_u7_n170 ) , .B1( u2_u14_u7_n179 ) );
  NAND4_X1 u2_u14_u7_U83 (.ZN( u2_out14_21 ) , .A4( u2_u14_u7_n157 ) , .A3( u2_u14_u7_n158 ) , .A2( u2_u14_u7_n159 ) , .A1( u2_u14_u7_n160 ) );
  OAI21_X1 u2_u14_u7_U84 (.B1( u2_u14_u7_n145 ) , .ZN( u2_u14_u7_n160 ) , .A( u2_u14_u7_n161 ) , .B2( u2_u14_u7_n177 ) );
  AOI22_X1 u2_u14_u7_U85 (.B2( u2_u14_u7_n149 ) , .B1( u2_u14_u7_n150 ) , .A2( u2_u14_u7_n151 ) , .A1( u2_u14_u7_n152 ) , .ZN( u2_u14_u7_n158 ) );
  NAND4_X1 u2_u14_u7_U86 (.ZN( u2_out14_15 ) , .A4( u2_u14_u7_n142 ) , .A3( u2_u14_u7_n143 ) , .A2( u2_u14_u7_n144 ) , .A1( u2_u14_u7_n178 ) );
  OR2_X1 u2_u14_u7_U87 (.A2( u2_u14_u7_n125 ) , .A1( u2_u14_u7_n129 ) , .ZN( u2_u14_u7_n144 ) );
  AOI22_X1 u2_u14_u7_U88 (.A2( u2_u14_u7_n126 ) , .ZN( u2_u14_u7_n143 ) , .B2( u2_u14_u7_n165 ) , .B1( u2_u14_u7_n173 ) , .A1( u2_u14_u7_n174 ) );
  NAND4_X1 u2_u14_u7_U89 (.ZN( u2_out14_5 ) , .A4( u2_u14_u7_n108 ) , .A3( u2_u14_u7_n109 ) , .A1( u2_u14_u7_n116 ) , .A2( u2_u14_u7_n123 ) );
  AND3_X1 u2_u14_u7_U9 (.A3( u2_u14_u7_n110 ) , .A2( u2_u14_u7_n127 ) , .A1( u2_u14_u7_n132 ) , .ZN( u2_u14_u7_n92 ) );
  AOI22_X1 u2_u14_u7_U90 (.ZN( u2_u14_u7_n109 ) , .A2( u2_u14_u7_n126 ) , .B2( u2_u14_u7_n145 ) , .B1( u2_u14_u7_n156 ) , .A1( u2_u14_u7_n171 ) );
  NOR4_X1 u2_u14_u7_U91 (.A4( u2_u14_u7_n104 ) , .A3( u2_u14_u7_n105 ) , .A2( u2_u14_u7_n106 ) , .A1( u2_u14_u7_n107 ) , .ZN( u2_u14_u7_n108 ) );
  OAI211_X1 u2_u14_u7_U92 (.B( u2_u14_u7_n122 ) , .A( u2_u14_u7_n123 ) , .C2( u2_u14_u7_n124 ) , .ZN( u2_u14_u7_n154 ) , .C1( u2_u14_u7_n162 ) );
  AOI222_X1 u2_u14_u7_U93 (.ZN( u2_u14_u7_n122 ) , .C2( u2_u14_u7_n126 ) , .C1( u2_u14_u7_n145 ) , .B1( u2_u14_u7_n161 ) , .A2( u2_u14_u7_n165 ) , .B2( u2_u14_u7_n170 ) , .A1( u2_u14_u7_n176 ) );
  INV_X1 u2_u14_u7_U94 (.A( u2_u14_u7_n111 ) , .ZN( u2_u14_u7_n170 ) );
  NAND3_X1 u2_u14_u7_U95 (.A3( u2_u14_u7_n146 ) , .A2( u2_u14_u7_n147 ) , .A1( u2_u14_u7_n148 ) , .ZN( u2_u14_u7_n151 ) );
  NAND3_X1 u2_u14_u7_U96 (.A3( u2_u14_u7_n131 ) , .A2( u2_u14_u7_n132 ) , .A1( u2_u14_u7_n133 ) , .ZN( u2_u14_u7_n135 ) );
  XOR2_X1 u2_u15_U1 (.A( u2_FP_38 ) , .B( u2_K16_9 ) , .Z( u2_u15_X_9 ) );
  XOR2_X1 u2_u15_U2 (.A( u2_FP_37 ) , .B( u2_K16_8 ) , .Z( u2_u15_X_8 ) );
  XOR2_X1 u2_u15_U3 (.A( u2_FP_36 ) , .B( u2_K16_7 ) , .Z( u2_u15_X_7 ) );
  XOR2_X1 u2_u15_U33 (.A( u2_FP_49 ) , .B( u2_K16_24 ) , .Z( u2_u15_X_24 ) );
  XOR2_X1 u2_u15_U34 (.A( u2_FP_48 ) , .B( u2_K16_23 ) , .Z( u2_u15_X_23 ) );
  XOR2_X1 u2_u15_U35 (.A( u2_FP_47 ) , .B( u2_K16_22 ) , .Z( u2_u15_X_22 ) );
  XOR2_X1 u2_u15_U36 (.A( u2_FP_46 ) , .B( u2_K16_21 ) , .Z( u2_u15_X_21 ) );
  XOR2_X1 u2_u15_U37 (.A( u2_FP_45 ) , .B( u2_K16_20 ) , .Z( u2_u15_X_20 ) );
  XOR2_X1 u2_u15_U39 (.A( u2_FP_44 ) , .B( u2_K16_19 ) , .Z( u2_u15_X_19 ) );
  XOR2_X1 u2_u15_U40 (.A( u2_FP_45 ) , .B( u2_K16_18 ) , .Z( u2_u15_X_18 ) );
  XOR2_X1 u2_u15_U41 (.A( u2_FP_44 ) , .B( u2_K16_17 ) , .Z( u2_u15_X_17 ) );
  XOR2_X1 u2_u15_U42 (.A( u2_FP_43 ) , .B( u2_K16_16 ) , .Z( u2_u15_X_16 ) );
  XOR2_X1 u2_u15_U43 (.A( u2_FP_42 ) , .B( u2_K16_15 ) , .Z( u2_u15_X_15 ) );
  XOR2_X1 u2_u15_U44 (.A( u2_FP_41 ) , .B( u2_K16_14 ) , .Z( u2_u15_X_14 ) );
  XOR2_X1 u2_u15_U45 (.A( u2_FP_40 ) , .B( u2_K16_13 ) , .Z( u2_u15_X_13 ) );
  XOR2_X1 u2_u15_U46 (.A( u2_FP_41 ) , .B( u2_K16_12 ) , .Z( u2_u15_X_12 ) );
  XOR2_X1 u2_u15_U47 (.A( u2_FP_40 ) , .B( u2_K16_11 ) , .Z( u2_u15_X_11 ) );
  XOR2_X1 u2_u15_U48 (.A( u2_FP_39 ) , .B( u2_K16_10 ) , .Z( u2_u15_X_10 ) );
  NOR2_X1 u2_u15_u1_U10 (.A1( u2_u15_u1_n112 ) , .A2( u2_u15_u1_n116 ) , .ZN( u2_u15_u1_n118 ) );
  NAND3_X1 u2_u15_u1_U100 (.ZN( u2_u15_u1_n113 ) , .A1( u2_u15_u1_n120 ) , .A3( u2_u15_u1_n133 ) , .A2( u2_u15_u1_n155 ) );
  OAI21_X1 u2_u15_u1_U11 (.ZN( u2_u15_u1_n101 ) , .B1( u2_u15_u1_n141 ) , .A( u2_u15_u1_n146 ) , .B2( u2_u15_u1_n183 ) );
  AOI21_X1 u2_u15_u1_U12 (.B2( u2_u15_u1_n155 ) , .B1( u2_u15_u1_n156 ) , .ZN( u2_u15_u1_n157 ) , .A( u2_u15_u1_n174 ) );
  NAND2_X1 u2_u15_u1_U13 (.ZN( u2_u15_u1_n140 ) , .A2( u2_u15_u1_n150 ) , .A1( u2_u15_u1_n155 ) );
  NAND2_X1 u2_u15_u1_U14 (.A1( u2_u15_u1_n131 ) , .ZN( u2_u15_u1_n147 ) , .A2( u2_u15_u1_n153 ) );
  INV_X1 u2_u15_u1_U15 (.A( u2_u15_u1_n139 ) , .ZN( u2_u15_u1_n174 ) );
  OR4_X1 u2_u15_u1_U16 (.A4( u2_u15_u1_n106 ) , .A3( u2_u15_u1_n107 ) , .ZN( u2_u15_u1_n108 ) , .A1( u2_u15_u1_n117 ) , .A2( u2_u15_u1_n184 ) );
  AOI21_X1 u2_u15_u1_U17 (.ZN( u2_u15_u1_n106 ) , .A( u2_u15_u1_n112 ) , .B1( u2_u15_u1_n154 ) , .B2( u2_u15_u1_n156 ) );
  AOI21_X1 u2_u15_u1_U18 (.ZN( u2_u15_u1_n107 ) , .B1( u2_u15_u1_n134 ) , .B2( u2_u15_u1_n149 ) , .A( u2_u15_u1_n174 ) );
  INV_X1 u2_u15_u1_U19 (.A( u2_u15_u1_n101 ) , .ZN( u2_u15_u1_n184 ) );
  INV_X1 u2_u15_u1_U20 (.A( u2_u15_u1_n112 ) , .ZN( u2_u15_u1_n171 ) );
  NAND2_X1 u2_u15_u1_U21 (.ZN( u2_u15_u1_n141 ) , .A1( u2_u15_u1_n153 ) , .A2( u2_u15_u1_n156 ) );
  AND2_X1 u2_u15_u1_U22 (.A1( u2_u15_u1_n123 ) , .ZN( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n161 ) );
  NAND2_X1 u2_u15_u1_U23 (.A2( u2_u15_u1_n115 ) , .A1( u2_u15_u1_n116 ) , .ZN( u2_u15_u1_n148 ) );
  NAND2_X1 u2_u15_u1_U24 (.A2( u2_u15_u1_n133 ) , .A1( u2_u15_u1_n135 ) , .ZN( u2_u15_u1_n159 ) );
  NAND2_X1 u2_u15_u1_U25 (.A2( u2_u15_u1_n115 ) , .A1( u2_u15_u1_n120 ) , .ZN( u2_u15_u1_n132 ) );
  INV_X1 u2_u15_u1_U26 (.A( u2_u15_u1_n154 ) , .ZN( u2_u15_u1_n178 ) );
  INV_X1 u2_u15_u1_U27 (.A( u2_u15_u1_n151 ) , .ZN( u2_u15_u1_n183 ) );
  AND2_X1 u2_u15_u1_U28 (.A1( u2_u15_u1_n129 ) , .A2( u2_u15_u1_n133 ) , .ZN( u2_u15_u1_n149 ) );
  INV_X1 u2_u15_u1_U29 (.A( u2_u15_u1_n131 ) , .ZN( u2_u15_u1_n180 ) );
  INV_X1 u2_u15_u1_U3 (.A( u2_u15_u1_n159 ) , .ZN( u2_u15_u1_n182 ) );
  OAI221_X1 u2_u15_u1_U30 (.A( u2_u15_u1_n119 ) , .C2( u2_u15_u1_n129 ) , .ZN( u2_u15_u1_n138 ) , .B2( u2_u15_u1_n152 ) , .C1( u2_u15_u1_n174 ) , .B1( u2_u15_u1_n187 ) );
  INV_X1 u2_u15_u1_U31 (.A( u2_u15_u1_n148 ) , .ZN( u2_u15_u1_n187 ) );
  AOI211_X1 u2_u15_u1_U32 (.B( u2_u15_u1_n117 ) , .A( u2_u15_u1_n118 ) , .ZN( u2_u15_u1_n119 ) , .C2( u2_u15_u1_n146 ) , .C1( u2_u15_u1_n159 ) );
  NOR2_X1 u2_u15_u1_U33 (.A1( u2_u15_u1_n168 ) , .A2( u2_u15_u1_n176 ) , .ZN( u2_u15_u1_n98 ) );
  AOI211_X1 u2_u15_u1_U34 (.B( u2_u15_u1_n162 ) , .A( u2_u15_u1_n163 ) , .C2( u2_u15_u1_n164 ) , .ZN( u2_u15_u1_n165 ) , .C1( u2_u15_u1_n171 ) );
  AOI21_X1 u2_u15_u1_U35 (.A( u2_u15_u1_n160 ) , .B2( u2_u15_u1_n161 ) , .ZN( u2_u15_u1_n162 ) , .B1( u2_u15_u1_n182 ) );
  OR2_X1 u2_u15_u1_U36 (.A2( u2_u15_u1_n157 ) , .A1( u2_u15_u1_n158 ) , .ZN( u2_u15_u1_n163 ) );
  NAND2_X1 u2_u15_u1_U37 (.A1( u2_u15_u1_n128 ) , .ZN( u2_u15_u1_n146 ) , .A2( u2_u15_u1_n160 ) );
  NAND2_X1 u2_u15_u1_U38 (.A2( u2_u15_u1_n112 ) , .ZN( u2_u15_u1_n139 ) , .A1( u2_u15_u1_n152 ) );
  NAND2_X1 u2_u15_u1_U39 (.A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n156 ) , .A2( u2_u15_u1_n99 ) );
  AOI221_X1 u2_u15_u1_U4 (.A( u2_u15_u1_n138 ) , .C2( u2_u15_u1_n139 ) , .C1( u2_u15_u1_n140 ) , .B2( u2_u15_u1_n141 ) , .ZN( u2_u15_u1_n142 ) , .B1( u2_u15_u1_n175 ) );
  AOI221_X1 u2_u15_u1_U40 (.B1( u2_u15_u1_n140 ) , .ZN( u2_u15_u1_n167 ) , .B2( u2_u15_u1_n172 ) , .C2( u2_u15_u1_n175 ) , .C1( u2_u15_u1_n178 ) , .A( u2_u15_u1_n188 ) );
  INV_X1 u2_u15_u1_U41 (.ZN( u2_u15_u1_n188 ) , .A( u2_u15_u1_n97 ) );
  AOI211_X1 u2_u15_u1_U42 (.A( u2_u15_u1_n118 ) , .C1( u2_u15_u1_n132 ) , .C2( u2_u15_u1_n139 ) , .B( u2_u15_u1_n96 ) , .ZN( u2_u15_u1_n97 ) );
  AOI21_X1 u2_u15_u1_U43 (.B2( u2_u15_u1_n121 ) , .B1( u2_u15_u1_n135 ) , .A( u2_u15_u1_n152 ) , .ZN( u2_u15_u1_n96 ) );
  NOR2_X1 u2_u15_u1_U44 (.ZN( u2_u15_u1_n117 ) , .A1( u2_u15_u1_n121 ) , .A2( u2_u15_u1_n160 ) );
  AOI21_X1 u2_u15_u1_U45 (.A( u2_u15_u1_n128 ) , .B2( u2_u15_u1_n129 ) , .ZN( u2_u15_u1_n130 ) , .B1( u2_u15_u1_n150 ) );
  OAI21_X1 u2_u15_u1_U46 (.B2( u2_u15_u1_n123 ) , .ZN( u2_u15_u1_n145 ) , .B1( u2_u15_u1_n160 ) , .A( u2_u15_u1_n185 ) );
  INV_X1 u2_u15_u1_U47 (.A( u2_u15_u1_n122 ) , .ZN( u2_u15_u1_n185 ) );
  AOI21_X1 u2_u15_u1_U48 (.B2( u2_u15_u1_n120 ) , .B1( u2_u15_u1_n121 ) , .ZN( u2_u15_u1_n122 ) , .A( u2_u15_u1_n128 ) );
  NAND2_X1 u2_u15_u1_U49 (.ZN( u2_u15_u1_n112 ) , .A1( u2_u15_u1_n169 ) , .A2( u2_u15_u1_n170 ) );
  AOI211_X1 u2_u15_u1_U5 (.ZN( u2_u15_u1_n124 ) , .A( u2_u15_u1_n138 ) , .C2( u2_u15_u1_n139 ) , .B( u2_u15_u1_n145 ) , .C1( u2_u15_u1_n147 ) );
  NAND2_X1 u2_u15_u1_U50 (.ZN( u2_u15_u1_n129 ) , .A2( u2_u15_u1_n95 ) , .A1( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U51 (.A1( u2_u15_u1_n102 ) , .ZN( u2_u15_u1_n154 ) , .A2( u2_u15_u1_n99 ) );
  NAND2_X1 u2_u15_u1_U52 (.A2( u2_u15_u1_n100 ) , .ZN( u2_u15_u1_n135 ) , .A1( u2_u15_u1_n99 ) );
  AOI21_X1 u2_u15_u1_U53 (.A( u2_u15_u1_n152 ) , .B2( u2_u15_u1_n153 ) , .B1( u2_u15_u1_n154 ) , .ZN( u2_u15_u1_n158 ) );
  INV_X1 u2_u15_u1_U54 (.A( u2_u15_u1_n160 ) , .ZN( u2_u15_u1_n175 ) );
  NAND2_X1 u2_u15_u1_U55 (.A1( u2_u15_u1_n100 ) , .ZN( u2_u15_u1_n116 ) , .A2( u2_u15_u1_n95 ) );
  NAND2_X1 u2_u15_u1_U56 (.A1( u2_u15_u1_n102 ) , .ZN( u2_u15_u1_n131 ) , .A2( u2_u15_u1_n95 ) );
  NAND2_X1 u2_u15_u1_U57 (.A2( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n121 ) , .A1( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U58 (.A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n153 ) , .A2( u2_u15_u1_n98 ) );
  NAND2_X1 u2_u15_u1_U59 (.A2( u2_u15_u1_n104 ) , .A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n133 ) );
  AOI22_X1 u2_u15_u1_U6 (.B2( u2_u15_u1_n136 ) , .A2( u2_u15_u1_n137 ) , .ZN( u2_u15_u1_n143 ) , .A1( u2_u15_u1_n171 ) , .B1( u2_u15_u1_n173 ) );
  NAND2_X1 u2_u15_u1_U60 (.ZN( u2_u15_u1_n150 ) , .A2( u2_u15_u1_n98 ) , .A1( u2_u15_u1_n99 ) );
  NAND2_X1 u2_u15_u1_U61 (.A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n155 ) , .A2( u2_u15_u1_n95 ) );
  OAI21_X1 u2_u15_u1_U62 (.ZN( u2_u15_u1_n109 ) , .B1( u2_u15_u1_n129 ) , .B2( u2_u15_u1_n160 ) , .A( u2_u15_u1_n167 ) );
  NAND2_X1 u2_u15_u1_U63 (.A2( u2_u15_u1_n100 ) , .A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n120 ) );
  NAND2_X1 u2_u15_u1_U64 (.A1( u2_u15_u1_n102 ) , .A2( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n115 ) );
  NAND2_X1 u2_u15_u1_U65 (.A2( u2_u15_u1_n100 ) , .A1( u2_u15_u1_n104 ) , .ZN( u2_u15_u1_n151 ) );
  NAND2_X1 u2_u15_u1_U66 (.A2( u2_u15_u1_n103 ) , .A1( u2_u15_u1_n105 ) , .ZN( u2_u15_u1_n161 ) );
  INV_X1 u2_u15_u1_U67 (.A( u2_u15_u1_n152 ) , .ZN( u2_u15_u1_n173 ) );
  INV_X1 u2_u15_u1_U68 (.A( u2_u15_u1_n128 ) , .ZN( u2_u15_u1_n172 ) );
  NAND2_X1 u2_u15_u1_U69 (.A2( u2_u15_u1_n102 ) , .A1( u2_u15_u1_n103 ) , .ZN( u2_u15_u1_n123 ) );
  INV_X1 u2_u15_u1_U7 (.A( u2_u15_u1_n147 ) , .ZN( u2_u15_u1_n181 ) );
  NOR2_X1 u2_u15_u1_U70 (.A2( u2_u15_X_7 ) , .A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n95 ) );
  NOR2_X1 u2_u15_u1_U71 (.A1( u2_u15_X_12 ) , .A2( u2_u15_X_9 ) , .ZN( u2_u15_u1_n100 ) );
  NOR2_X1 u2_u15_u1_U72 (.A2( u2_u15_X_8 ) , .A1( u2_u15_u1_n177 ) , .ZN( u2_u15_u1_n99 ) );
  NOR2_X1 u2_u15_u1_U73 (.A2( u2_u15_X_12 ) , .ZN( u2_u15_u1_n102 ) , .A1( u2_u15_u1_n176 ) );
  NOR2_X1 u2_u15_u1_U74 (.A2( u2_u15_X_9 ) , .ZN( u2_u15_u1_n105 ) , .A1( u2_u15_u1_n168 ) );
  NAND2_X1 u2_u15_u1_U75 (.A1( u2_u15_X_10 ) , .ZN( u2_u15_u1_n160 ) , .A2( u2_u15_u1_n169 ) );
  NAND2_X1 u2_u15_u1_U76 (.A2( u2_u15_X_10 ) , .A1( u2_u15_X_11 ) , .ZN( u2_u15_u1_n152 ) );
  NAND2_X1 u2_u15_u1_U77 (.A1( u2_u15_X_11 ) , .ZN( u2_u15_u1_n128 ) , .A2( u2_u15_u1_n170 ) );
  AND2_X1 u2_u15_u1_U78 (.A2( u2_u15_X_7 ) , .A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n104 ) );
  AND2_X1 u2_u15_u1_U79 (.A1( u2_u15_X_8 ) , .ZN( u2_u15_u1_n103 ) , .A2( u2_u15_u1_n177 ) );
  AOI22_X1 u2_u15_u1_U8 (.B2( u2_u15_u1_n113 ) , .A2( u2_u15_u1_n114 ) , .ZN( u2_u15_u1_n125 ) , .A1( u2_u15_u1_n171 ) , .B1( u2_u15_u1_n173 ) );
  INV_X1 u2_u15_u1_U80 (.A( u2_u15_X_10 ) , .ZN( u2_u15_u1_n170 ) );
  INV_X1 u2_u15_u1_U81 (.A( u2_u15_X_9 ) , .ZN( u2_u15_u1_n176 ) );
  INV_X1 u2_u15_u1_U82 (.A( u2_u15_X_11 ) , .ZN( u2_u15_u1_n169 ) );
  INV_X1 u2_u15_u1_U83 (.A( u2_u15_X_12 ) , .ZN( u2_u15_u1_n168 ) );
  INV_X1 u2_u15_u1_U84 (.A( u2_u15_X_7 ) , .ZN( u2_u15_u1_n177 ) );
  NAND4_X1 u2_u15_u1_U85 (.ZN( u2_out15_18 ) , .A4( u2_u15_u1_n165 ) , .A3( u2_u15_u1_n166 ) , .A1( u2_u15_u1_n167 ) , .A2( u2_u15_u1_n186 ) );
  AOI22_X1 u2_u15_u1_U86 (.B2( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n147 ) , .A2( u2_u15_u1_n148 ) , .ZN( u2_u15_u1_n166 ) , .A1( u2_u15_u1_n172 ) );
  INV_X1 u2_u15_u1_U87 (.A( u2_u15_u1_n145 ) , .ZN( u2_u15_u1_n186 ) );
  NAND4_X1 u2_u15_u1_U88 (.ZN( u2_out15_2 ) , .A4( u2_u15_u1_n142 ) , .A3( u2_u15_u1_n143 ) , .A2( u2_u15_u1_n144 ) , .A1( u2_u15_u1_n179 ) );
  OAI21_X1 u2_u15_u1_U89 (.B2( u2_u15_u1_n132 ) , .ZN( u2_u15_u1_n144 ) , .A( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n180 ) );
  NAND2_X1 u2_u15_u1_U9 (.ZN( u2_u15_u1_n114 ) , .A1( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n156 ) );
  INV_X1 u2_u15_u1_U90 (.A( u2_u15_u1_n130 ) , .ZN( u2_u15_u1_n179 ) );
  NAND4_X1 u2_u15_u1_U91 (.ZN( u2_out15_28 ) , .A4( u2_u15_u1_n124 ) , .A3( u2_u15_u1_n125 ) , .A2( u2_u15_u1_n126 ) , .A1( u2_u15_u1_n127 ) );
  OAI21_X1 u2_u15_u1_U92 (.ZN( u2_u15_u1_n127 ) , .B2( u2_u15_u1_n139 ) , .B1( u2_u15_u1_n175 ) , .A( u2_u15_u1_n183 ) );
  OAI21_X1 u2_u15_u1_U93 (.ZN( u2_u15_u1_n126 ) , .B2( u2_u15_u1_n140 ) , .A( u2_u15_u1_n146 ) , .B1( u2_u15_u1_n178 ) );
  OR4_X1 u2_u15_u1_U94 (.ZN( u2_out15_13 ) , .A4( u2_u15_u1_n108 ) , .A3( u2_u15_u1_n109 ) , .A2( u2_u15_u1_n110 ) , .A1( u2_u15_u1_n111 ) );
  AOI21_X1 u2_u15_u1_U95 (.ZN( u2_u15_u1_n111 ) , .A( u2_u15_u1_n128 ) , .B2( u2_u15_u1_n131 ) , .B1( u2_u15_u1_n135 ) );
  AOI21_X1 u2_u15_u1_U96 (.ZN( u2_u15_u1_n110 ) , .A( u2_u15_u1_n116 ) , .B1( u2_u15_u1_n152 ) , .B2( u2_u15_u1_n160 ) );
  NAND3_X1 u2_u15_u1_U97 (.A3( u2_u15_u1_n149 ) , .A2( u2_u15_u1_n150 ) , .A1( u2_u15_u1_n151 ) , .ZN( u2_u15_u1_n164 ) );
  NAND3_X1 u2_u15_u1_U98 (.A3( u2_u15_u1_n134 ) , .A2( u2_u15_u1_n135 ) , .ZN( u2_u15_u1_n136 ) , .A1( u2_u15_u1_n151 ) );
  NAND3_X1 u2_u15_u1_U99 (.A1( u2_u15_u1_n133 ) , .ZN( u2_u15_u1_n137 ) , .A2( u2_u15_u1_n154 ) , .A3( u2_u15_u1_n181 ) );
  OAI22_X1 u2_u15_u2_U10 (.B1( u2_u15_u2_n151 ) , .A2( u2_u15_u2_n152 ) , .A1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n160 ) , .B2( u2_u15_u2_n168 ) );
  NAND3_X1 u2_u15_u2_U100 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n98 ) );
  NOR3_X1 u2_u15_u2_U11 (.A1( u2_u15_u2_n150 ) , .ZN( u2_u15_u2_n151 ) , .A3( u2_u15_u2_n175 ) , .A2( u2_u15_u2_n188 ) );
  AOI21_X1 u2_u15_u2_U12 (.B2( u2_u15_u2_n123 ) , .ZN( u2_u15_u2_n125 ) , .A( u2_u15_u2_n171 ) , .B1( u2_u15_u2_n184 ) );
  INV_X1 u2_u15_u2_U13 (.A( u2_u15_u2_n150 ) , .ZN( u2_u15_u2_n184 ) );
  AOI21_X1 u2_u15_u2_U14 (.ZN( u2_u15_u2_n144 ) , .B2( u2_u15_u2_n155 ) , .A( u2_u15_u2_n172 ) , .B1( u2_u15_u2_n185 ) );
  AOI21_X1 u2_u15_u2_U15 (.B2( u2_u15_u2_n143 ) , .ZN( u2_u15_u2_n145 ) , .B1( u2_u15_u2_n152 ) , .A( u2_u15_u2_n171 ) );
  INV_X1 u2_u15_u2_U16 (.A( u2_u15_u2_n156 ) , .ZN( u2_u15_u2_n171 ) );
  INV_X1 u2_u15_u2_U17 (.A( u2_u15_u2_n120 ) , .ZN( u2_u15_u2_n188 ) );
  NAND2_X1 u2_u15_u2_U18 (.A2( u2_u15_u2_n122 ) , .ZN( u2_u15_u2_n150 ) , .A1( u2_u15_u2_n152 ) );
  INV_X1 u2_u15_u2_U19 (.A( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n170 ) );
  INV_X1 u2_u15_u2_U20 (.A( u2_u15_u2_n137 ) , .ZN( u2_u15_u2_n173 ) );
  NAND2_X1 u2_u15_u2_U21 (.A1( u2_u15_u2_n132 ) , .A2( u2_u15_u2_n139 ) , .ZN( u2_u15_u2_n157 ) );
  INV_X1 u2_u15_u2_U22 (.A( u2_u15_u2_n113 ) , .ZN( u2_u15_u2_n178 ) );
  INV_X1 u2_u15_u2_U23 (.A( u2_u15_u2_n139 ) , .ZN( u2_u15_u2_n175 ) );
  INV_X1 u2_u15_u2_U24 (.A( u2_u15_u2_n155 ) , .ZN( u2_u15_u2_n181 ) );
  INV_X1 u2_u15_u2_U25 (.A( u2_u15_u2_n119 ) , .ZN( u2_u15_u2_n177 ) );
  INV_X1 u2_u15_u2_U26 (.A( u2_u15_u2_n116 ) , .ZN( u2_u15_u2_n180 ) );
  INV_X1 u2_u15_u2_U27 (.A( u2_u15_u2_n131 ) , .ZN( u2_u15_u2_n179 ) );
  INV_X1 u2_u15_u2_U28 (.A( u2_u15_u2_n154 ) , .ZN( u2_u15_u2_n176 ) );
  NAND2_X1 u2_u15_u2_U29 (.A2( u2_u15_u2_n116 ) , .A1( u2_u15_u2_n117 ) , .ZN( u2_u15_u2_n118 ) );
  NOR2_X1 u2_u15_u2_U3 (.ZN( u2_u15_u2_n121 ) , .A2( u2_u15_u2_n177 ) , .A1( u2_u15_u2_n180 ) );
  INV_X1 u2_u15_u2_U30 (.A( u2_u15_u2_n132 ) , .ZN( u2_u15_u2_n182 ) );
  INV_X1 u2_u15_u2_U31 (.A( u2_u15_u2_n158 ) , .ZN( u2_u15_u2_n183 ) );
  OAI21_X1 u2_u15_u2_U32 (.A( u2_u15_u2_n156 ) , .B1( u2_u15_u2_n157 ) , .ZN( u2_u15_u2_n158 ) , .B2( u2_u15_u2_n179 ) );
  NOR2_X1 u2_u15_u2_U33 (.ZN( u2_u15_u2_n156 ) , .A1( u2_u15_u2_n166 ) , .A2( u2_u15_u2_n169 ) );
  NOR2_X1 u2_u15_u2_U34 (.A2( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n137 ) , .A1( u2_u15_u2_n140 ) );
  NOR2_X1 u2_u15_u2_U35 (.A2( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n153 ) , .A1( u2_u15_u2_n156 ) );
  AOI211_X1 u2_u15_u2_U36 (.ZN( u2_u15_u2_n130 ) , .C1( u2_u15_u2_n138 ) , .C2( u2_u15_u2_n179 ) , .B( u2_u15_u2_n96 ) , .A( u2_u15_u2_n97 ) );
  OAI22_X1 u2_u15_u2_U37 (.B1( u2_u15_u2_n133 ) , .A2( u2_u15_u2_n137 ) , .A1( u2_u15_u2_n152 ) , .B2( u2_u15_u2_n168 ) , .ZN( u2_u15_u2_n97 ) );
  OAI221_X1 u2_u15_u2_U38 (.B1( u2_u15_u2_n113 ) , .C1( u2_u15_u2_n132 ) , .A( u2_u15_u2_n149 ) , .B2( u2_u15_u2_n171 ) , .C2( u2_u15_u2_n172 ) , .ZN( u2_u15_u2_n96 ) );
  OAI221_X1 u2_u15_u2_U39 (.A( u2_u15_u2_n115 ) , .C2( u2_u15_u2_n123 ) , .B2( u2_u15_u2_n143 ) , .B1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n163 ) , .C1( u2_u15_u2_n168 ) );
  INV_X1 u2_u15_u2_U4 (.A( u2_u15_u2_n134 ) , .ZN( u2_u15_u2_n185 ) );
  OAI21_X1 u2_u15_u2_U40 (.A( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n115 ) , .B1( u2_u15_u2_n176 ) , .B2( u2_u15_u2_n178 ) );
  OAI221_X1 u2_u15_u2_U41 (.A( u2_u15_u2_n135 ) , .B2( u2_u15_u2_n136 ) , .B1( u2_u15_u2_n137 ) , .ZN( u2_u15_u2_n162 ) , .C2( u2_u15_u2_n167 ) , .C1( u2_u15_u2_n185 ) );
  AND3_X1 u2_u15_u2_U42 (.A3( u2_u15_u2_n131 ) , .A2( u2_u15_u2_n132 ) , .A1( u2_u15_u2_n133 ) , .ZN( u2_u15_u2_n136 ) );
  AOI22_X1 u2_u15_u2_U43 (.ZN( u2_u15_u2_n135 ) , .B1( u2_u15_u2_n140 ) , .A1( u2_u15_u2_n156 ) , .B2( u2_u15_u2_n180 ) , .A2( u2_u15_u2_n188 ) );
  AOI21_X1 u2_u15_u2_U44 (.ZN( u2_u15_u2_n149 ) , .B1( u2_u15_u2_n173 ) , .B2( u2_u15_u2_n188 ) , .A( u2_u15_u2_n95 ) );
  AND3_X1 u2_u15_u2_U45 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n156 ) , .ZN( u2_u15_u2_n95 ) );
  OAI21_X1 u2_u15_u2_U46 (.A( u2_u15_u2_n141 ) , .B2( u2_u15_u2_n142 ) , .ZN( u2_u15_u2_n146 ) , .B1( u2_u15_u2_n153 ) );
  OAI21_X1 u2_u15_u2_U47 (.A( u2_u15_u2_n140 ) , .ZN( u2_u15_u2_n141 ) , .B1( u2_u15_u2_n176 ) , .B2( u2_u15_u2_n177 ) );
  NOR3_X1 u2_u15_u2_U48 (.ZN( u2_u15_u2_n142 ) , .A3( u2_u15_u2_n175 ) , .A2( u2_u15_u2_n178 ) , .A1( u2_u15_u2_n181 ) );
  OAI21_X1 u2_u15_u2_U49 (.A( u2_u15_u2_n101 ) , .B2( u2_u15_u2_n121 ) , .B1( u2_u15_u2_n153 ) , .ZN( u2_u15_u2_n164 ) );
  NOR4_X1 u2_u15_u2_U5 (.A4( u2_u15_u2_n124 ) , .A3( u2_u15_u2_n125 ) , .A2( u2_u15_u2_n126 ) , .A1( u2_u15_u2_n127 ) , .ZN( u2_u15_u2_n128 ) );
  NAND2_X1 u2_u15_u2_U50 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n155 ) );
  NAND2_X1 u2_u15_u2_U51 (.A2( u2_u15_u2_n105 ) , .A1( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n143 ) );
  NAND2_X1 u2_u15_u2_U52 (.A1( u2_u15_u2_n104 ) , .A2( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n152 ) );
  NAND2_X1 u2_u15_u2_U53 (.A1( u2_u15_u2_n100 ) , .A2( u2_u15_u2_n105 ) , .ZN( u2_u15_u2_n132 ) );
  INV_X1 u2_u15_u2_U54 (.A( u2_u15_u2_n140 ) , .ZN( u2_u15_u2_n168 ) );
  INV_X1 u2_u15_u2_U55 (.A( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n167 ) );
  INV_X1 u2_u15_u2_U56 (.ZN( u2_u15_u2_n187 ) , .A( u2_u15_u2_n99 ) );
  OAI21_X1 u2_u15_u2_U57 (.B1( u2_u15_u2_n137 ) , .B2( u2_u15_u2_n143 ) , .A( u2_u15_u2_n98 ) , .ZN( u2_u15_u2_n99 ) );
  NAND2_X1 u2_u15_u2_U58 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n113 ) );
  NAND2_X1 u2_u15_u2_U59 (.A1( u2_u15_u2_n106 ) , .A2( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n131 ) );
  AOI21_X1 u2_u15_u2_U6 (.B2( u2_u15_u2_n119 ) , .ZN( u2_u15_u2_n127 ) , .A( u2_u15_u2_n137 ) , .B1( u2_u15_u2_n155 ) );
  NAND2_X1 u2_u15_u2_U60 (.A1( u2_u15_u2_n103 ) , .A2( u2_u15_u2_n107 ) , .ZN( u2_u15_u2_n139 ) );
  NAND2_X1 u2_u15_u2_U61 (.A1( u2_u15_u2_n103 ) , .A2( u2_u15_u2_n105 ) , .ZN( u2_u15_u2_n133 ) );
  NAND2_X1 u2_u15_u2_U62 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n103 ) , .ZN( u2_u15_u2_n154 ) );
  NAND2_X1 u2_u15_u2_U63 (.A2( u2_u15_u2_n103 ) , .A1( u2_u15_u2_n104 ) , .ZN( u2_u15_u2_n119 ) );
  NAND2_X1 u2_u15_u2_U64 (.A2( u2_u15_u2_n107 ) , .A1( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n123 ) );
  NAND2_X1 u2_u15_u2_U65 (.A1( u2_u15_u2_n104 ) , .A2( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n122 ) );
  INV_X1 u2_u15_u2_U66 (.A( u2_u15_u2_n114 ) , .ZN( u2_u15_u2_n172 ) );
  NAND2_X1 u2_u15_u2_U67 (.A2( u2_u15_u2_n100 ) , .A1( u2_u15_u2_n102 ) , .ZN( u2_u15_u2_n116 ) );
  NAND2_X1 u2_u15_u2_U68 (.A1( u2_u15_u2_n102 ) , .A2( u2_u15_u2_n108 ) , .ZN( u2_u15_u2_n120 ) );
  NAND2_X1 u2_u15_u2_U69 (.A2( u2_u15_u2_n105 ) , .A1( u2_u15_u2_n106 ) , .ZN( u2_u15_u2_n117 ) );
  AOI21_X1 u2_u15_u2_U7 (.ZN( u2_u15_u2_n124 ) , .B1( u2_u15_u2_n131 ) , .B2( u2_u15_u2_n143 ) , .A( u2_u15_u2_n172 ) );
  NOR2_X1 u2_u15_u2_U70 (.A2( u2_u15_X_16 ) , .ZN( u2_u15_u2_n140 ) , .A1( u2_u15_u2_n166 ) );
  NOR2_X1 u2_u15_u2_U71 (.A2( u2_u15_X_13 ) , .A1( u2_u15_X_14 ) , .ZN( u2_u15_u2_n100 ) );
  NOR2_X1 u2_u15_u2_U72 (.A2( u2_u15_X_16 ) , .A1( u2_u15_X_17 ) , .ZN( u2_u15_u2_n138 ) );
  NOR2_X1 u2_u15_u2_U73 (.A2( u2_u15_X_15 ) , .A1( u2_u15_X_18 ) , .ZN( u2_u15_u2_n104 ) );
  NOR2_X1 u2_u15_u2_U74 (.A2( u2_u15_X_14 ) , .ZN( u2_u15_u2_n103 ) , .A1( u2_u15_u2_n174 ) );
  NOR2_X1 u2_u15_u2_U75 (.A2( u2_u15_X_15 ) , .ZN( u2_u15_u2_n102 ) , .A1( u2_u15_u2_n165 ) );
  NOR2_X1 u2_u15_u2_U76 (.A2( u2_u15_X_17 ) , .ZN( u2_u15_u2_n114 ) , .A1( u2_u15_u2_n169 ) );
  AND2_X1 u2_u15_u2_U77 (.A1( u2_u15_X_15 ) , .ZN( u2_u15_u2_n105 ) , .A2( u2_u15_u2_n165 ) );
  AND2_X1 u2_u15_u2_U78 (.A2( u2_u15_X_15 ) , .A1( u2_u15_X_18 ) , .ZN( u2_u15_u2_n107 ) );
  AND2_X1 u2_u15_u2_U79 (.A1( u2_u15_X_14 ) , .ZN( u2_u15_u2_n106 ) , .A2( u2_u15_u2_n174 ) );
  AOI21_X1 u2_u15_u2_U8 (.B2( u2_u15_u2_n120 ) , .B1( u2_u15_u2_n121 ) , .ZN( u2_u15_u2_n126 ) , .A( u2_u15_u2_n167 ) );
  AND2_X1 u2_u15_u2_U80 (.A1( u2_u15_X_13 ) , .A2( u2_u15_X_14 ) , .ZN( u2_u15_u2_n108 ) );
  INV_X1 u2_u15_u2_U81 (.A( u2_u15_X_16 ) , .ZN( u2_u15_u2_n169 ) );
  INV_X1 u2_u15_u2_U82 (.A( u2_u15_X_17 ) , .ZN( u2_u15_u2_n166 ) );
  INV_X1 u2_u15_u2_U83 (.A( u2_u15_X_13 ) , .ZN( u2_u15_u2_n174 ) );
  INV_X1 u2_u15_u2_U84 (.A( u2_u15_X_18 ) , .ZN( u2_u15_u2_n165 ) );
  NAND4_X1 u2_u15_u2_U85 (.ZN( u2_out15_30 ) , .A4( u2_u15_u2_n147 ) , .A3( u2_u15_u2_n148 ) , .A2( u2_u15_u2_n149 ) , .A1( u2_u15_u2_n187 ) );
  NOR3_X1 u2_u15_u2_U86 (.A3( u2_u15_u2_n144 ) , .A2( u2_u15_u2_n145 ) , .A1( u2_u15_u2_n146 ) , .ZN( u2_u15_u2_n147 ) );
  AOI21_X1 u2_u15_u2_U87 (.B2( u2_u15_u2_n138 ) , .ZN( u2_u15_u2_n148 ) , .A( u2_u15_u2_n162 ) , .B1( u2_u15_u2_n182 ) );
  NAND4_X1 u2_u15_u2_U88 (.ZN( u2_out15_24 ) , .A4( u2_u15_u2_n111 ) , .A3( u2_u15_u2_n112 ) , .A1( u2_u15_u2_n130 ) , .A2( u2_u15_u2_n187 ) );
  AOI221_X1 u2_u15_u2_U89 (.A( u2_u15_u2_n109 ) , .B1( u2_u15_u2_n110 ) , .ZN( u2_u15_u2_n111 ) , .C1( u2_u15_u2_n134 ) , .C2( u2_u15_u2_n170 ) , .B2( u2_u15_u2_n173 ) );
  OAI22_X1 u2_u15_u2_U9 (.ZN( u2_u15_u2_n109 ) , .A2( u2_u15_u2_n113 ) , .B2( u2_u15_u2_n133 ) , .B1( u2_u15_u2_n167 ) , .A1( u2_u15_u2_n168 ) );
  AOI21_X1 u2_u15_u2_U90 (.ZN( u2_u15_u2_n112 ) , .B2( u2_u15_u2_n156 ) , .A( u2_u15_u2_n164 ) , .B1( u2_u15_u2_n181 ) );
  NAND4_X1 u2_u15_u2_U91 (.ZN( u2_out15_16 ) , .A4( u2_u15_u2_n128 ) , .A3( u2_u15_u2_n129 ) , .A1( u2_u15_u2_n130 ) , .A2( u2_u15_u2_n186 ) );
  AOI22_X1 u2_u15_u2_U92 (.A2( u2_u15_u2_n118 ) , .ZN( u2_u15_u2_n129 ) , .A1( u2_u15_u2_n140 ) , .B1( u2_u15_u2_n157 ) , .B2( u2_u15_u2_n170 ) );
  INV_X1 u2_u15_u2_U93 (.A( u2_u15_u2_n163 ) , .ZN( u2_u15_u2_n186 ) );
  OR4_X1 u2_u15_u2_U94 (.ZN( u2_out15_6 ) , .A4( u2_u15_u2_n161 ) , .A3( u2_u15_u2_n162 ) , .A2( u2_u15_u2_n163 ) , .A1( u2_u15_u2_n164 ) );
  OR3_X1 u2_u15_u2_U95 (.A2( u2_u15_u2_n159 ) , .A1( u2_u15_u2_n160 ) , .ZN( u2_u15_u2_n161 ) , .A3( u2_u15_u2_n183 ) );
  AOI21_X1 u2_u15_u2_U96 (.B2( u2_u15_u2_n154 ) , .B1( u2_u15_u2_n155 ) , .ZN( u2_u15_u2_n159 ) , .A( u2_u15_u2_n167 ) );
  NAND3_X1 u2_u15_u2_U97 (.A2( u2_u15_u2_n117 ) , .A1( u2_u15_u2_n122 ) , .A3( u2_u15_u2_n123 ) , .ZN( u2_u15_u2_n134 ) );
  NAND3_X1 u2_u15_u2_U98 (.ZN( u2_u15_u2_n110 ) , .A2( u2_u15_u2_n131 ) , .A3( u2_u15_u2_n139 ) , .A1( u2_u15_u2_n154 ) );
  NAND3_X1 u2_u15_u2_U99 (.A2( u2_u15_u2_n100 ) , .ZN( u2_u15_u2_n101 ) , .A1( u2_u15_u2_n104 ) , .A3( u2_u15_u2_n114 ) );
  OAI22_X1 u2_u15_u3_U10 (.B1( u2_u15_u3_n113 ) , .A2( u2_u15_u3_n135 ) , .A1( u2_u15_u3_n150 ) , .B2( u2_u15_u3_n164 ) , .ZN( u2_u15_u3_n98 ) );
  OAI211_X1 u2_u15_u3_U11 (.B( u2_u15_u3_n106 ) , .ZN( u2_u15_u3_n119 ) , .C2( u2_u15_u3_n128 ) , .C1( u2_u15_u3_n167 ) , .A( u2_u15_u3_n181 ) );
  AOI221_X1 u2_u15_u3_U12 (.C1( u2_u15_u3_n105 ) , .ZN( u2_u15_u3_n106 ) , .A( u2_u15_u3_n131 ) , .B2( u2_u15_u3_n132 ) , .C2( u2_u15_u3_n133 ) , .B1( u2_u15_u3_n169 ) );
  INV_X1 u2_u15_u3_U13 (.ZN( u2_u15_u3_n181 ) , .A( u2_u15_u3_n98 ) );
  NAND2_X1 u2_u15_u3_U14 (.ZN( u2_u15_u3_n105 ) , .A2( u2_u15_u3_n130 ) , .A1( u2_u15_u3_n155 ) );
  AOI22_X1 u2_u15_u3_U15 (.B1( u2_u15_u3_n115 ) , .A2( u2_u15_u3_n116 ) , .ZN( u2_u15_u3_n123 ) , .B2( u2_u15_u3_n133 ) , .A1( u2_u15_u3_n169 ) );
  NAND2_X1 u2_u15_u3_U16 (.ZN( u2_u15_u3_n116 ) , .A2( u2_u15_u3_n151 ) , .A1( u2_u15_u3_n182 ) );
  NOR2_X1 u2_u15_u3_U17 (.ZN( u2_u15_u3_n126 ) , .A2( u2_u15_u3_n150 ) , .A1( u2_u15_u3_n164 ) );
  AOI21_X1 u2_u15_u3_U18 (.ZN( u2_u15_u3_n112 ) , .B2( u2_u15_u3_n146 ) , .B1( u2_u15_u3_n155 ) , .A( u2_u15_u3_n167 ) );
  NAND2_X1 u2_u15_u3_U19 (.A1( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n142 ) , .A2( u2_u15_u3_n164 ) );
  NAND2_X1 u2_u15_u3_U20 (.ZN( u2_u15_u3_n132 ) , .A2( u2_u15_u3_n152 ) , .A1( u2_u15_u3_n156 ) );
  AND2_X1 u2_u15_u3_U21 (.A2( u2_u15_u3_n113 ) , .A1( u2_u15_u3_n114 ) , .ZN( u2_u15_u3_n151 ) );
  INV_X1 u2_u15_u3_U22 (.A( u2_u15_u3_n133 ) , .ZN( u2_u15_u3_n165 ) );
  INV_X1 u2_u15_u3_U23 (.A( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n170 ) );
  NAND2_X1 u2_u15_u3_U24 (.A1( u2_u15_u3_n107 ) , .A2( u2_u15_u3_n108 ) , .ZN( u2_u15_u3_n140 ) );
  NAND2_X1 u2_u15_u3_U25 (.ZN( u2_u15_u3_n117 ) , .A1( u2_u15_u3_n124 ) , .A2( u2_u15_u3_n148 ) );
  NAND2_X1 u2_u15_u3_U26 (.ZN( u2_u15_u3_n143 ) , .A1( u2_u15_u3_n165 ) , .A2( u2_u15_u3_n167 ) );
  INV_X1 u2_u15_u3_U27 (.A( u2_u15_u3_n130 ) , .ZN( u2_u15_u3_n177 ) );
  INV_X1 u2_u15_u3_U28 (.A( u2_u15_u3_n128 ) , .ZN( u2_u15_u3_n176 ) );
  INV_X1 u2_u15_u3_U29 (.A( u2_u15_u3_n155 ) , .ZN( u2_u15_u3_n174 ) );
  INV_X1 u2_u15_u3_U3 (.A( u2_u15_u3_n129 ) , .ZN( u2_u15_u3_n183 ) );
  INV_X1 u2_u15_u3_U30 (.A( u2_u15_u3_n139 ) , .ZN( u2_u15_u3_n185 ) );
  NOR2_X1 u2_u15_u3_U31 (.ZN( u2_u15_u3_n135 ) , .A2( u2_u15_u3_n141 ) , .A1( u2_u15_u3_n169 ) );
  OAI222_X1 u2_u15_u3_U32 (.C2( u2_u15_u3_n107 ) , .A2( u2_u15_u3_n108 ) , .B1( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n138 ) , .B2( u2_u15_u3_n146 ) , .C1( u2_u15_u3_n154 ) , .A1( u2_u15_u3_n164 ) );
  NOR4_X1 u2_u15_u3_U33 (.A4( u2_u15_u3_n157 ) , .A3( u2_u15_u3_n158 ) , .A2( u2_u15_u3_n159 ) , .A1( u2_u15_u3_n160 ) , .ZN( u2_u15_u3_n161 ) );
  AOI21_X1 u2_u15_u3_U34 (.B2( u2_u15_u3_n152 ) , .B1( u2_u15_u3_n153 ) , .ZN( u2_u15_u3_n158 ) , .A( u2_u15_u3_n164 ) );
  AOI21_X1 u2_u15_u3_U35 (.A( u2_u15_u3_n154 ) , .B2( u2_u15_u3_n155 ) , .B1( u2_u15_u3_n156 ) , .ZN( u2_u15_u3_n157 ) );
  AOI21_X1 u2_u15_u3_U36 (.A( u2_u15_u3_n149 ) , .B2( u2_u15_u3_n150 ) , .B1( u2_u15_u3_n151 ) , .ZN( u2_u15_u3_n159 ) );
  AOI211_X1 u2_u15_u3_U37 (.ZN( u2_u15_u3_n109 ) , .A( u2_u15_u3_n119 ) , .C2( u2_u15_u3_n129 ) , .B( u2_u15_u3_n138 ) , .C1( u2_u15_u3_n141 ) );
  AOI211_X1 u2_u15_u3_U38 (.B( u2_u15_u3_n119 ) , .A( u2_u15_u3_n120 ) , .C2( u2_u15_u3_n121 ) , .ZN( u2_u15_u3_n122 ) , .C1( u2_u15_u3_n179 ) );
  INV_X1 u2_u15_u3_U39 (.A( u2_u15_u3_n156 ) , .ZN( u2_u15_u3_n179 ) );
  INV_X1 u2_u15_u3_U4 (.A( u2_u15_u3_n140 ) , .ZN( u2_u15_u3_n182 ) );
  OAI22_X1 u2_u15_u3_U40 (.B1( u2_u15_u3_n118 ) , .ZN( u2_u15_u3_n120 ) , .A1( u2_u15_u3_n135 ) , .B2( u2_u15_u3_n154 ) , .A2( u2_u15_u3_n178 ) );
  AND3_X1 u2_u15_u3_U41 (.ZN( u2_u15_u3_n118 ) , .A2( u2_u15_u3_n124 ) , .A1( u2_u15_u3_n144 ) , .A3( u2_u15_u3_n152 ) );
  INV_X1 u2_u15_u3_U42 (.A( u2_u15_u3_n121 ) , .ZN( u2_u15_u3_n164 ) );
  NAND2_X1 u2_u15_u3_U43 (.ZN( u2_u15_u3_n133 ) , .A1( u2_u15_u3_n154 ) , .A2( u2_u15_u3_n164 ) );
  OAI211_X1 u2_u15_u3_U44 (.B( u2_u15_u3_n127 ) , .ZN( u2_u15_u3_n139 ) , .C1( u2_u15_u3_n150 ) , .C2( u2_u15_u3_n154 ) , .A( u2_u15_u3_n184 ) );
  INV_X1 u2_u15_u3_U45 (.A( u2_u15_u3_n125 ) , .ZN( u2_u15_u3_n184 ) );
  AOI221_X1 u2_u15_u3_U46 (.A( u2_u15_u3_n126 ) , .ZN( u2_u15_u3_n127 ) , .C2( u2_u15_u3_n132 ) , .C1( u2_u15_u3_n169 ) , .B2( u2_u15_u3_n170 ) , .B1( u2_u15_u3_n174 ) );
  OAI22_X1 u2_u15_u3_U47 (.A1( u2_u15_u3_n124 ) , .ZN( u2_u15_u3_n125 ) , .B2( u2_u15_u3_n145 ) , .A2( u2_u15_u3_n165 ) , .B1( u2_u15_u3_n167 ) );
  NOR2_X1 u2_u15_u3_U48 (.A1( u2_u15_u3_n113 ) , .ZN( u2_u15_u3_n131 ) , .A2( u2_u15_u3_n154 ) );
  NAND2_X1 u2_u15_u3_U49 (.A1( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n150 ) , .A2( u2_u15_u3_n99 ) );
  INV_X1 u2_u15_u3_U5 (.A( u2_u15_u3_n117 ) , .ZN( u2_u15_u3_n178 ) );
  NAND2_X1 u2_u15_u3_U50 (.A2( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n155 ) , .A1( u2_u15_u3_n97 ) );
  INV_X1 u2_u15_u3_U51 (.A( u2_u15_u3_n141 ) , .ZN( u2_u15_u3_n167 ) );
  AOI21_X1 u2_u15_u3_U52 (.B2( u2_u15_u3_n114 ) , .B1( u2_u15_u3_n146 ) , .A( u2_u15_u3_n154 ) , .ZN( u2_u15_u3_n94 ) );
  AOI21_X1 u2_u15_u3_U53 (.ZN( u2_u15_u3_n110 ) , .B2( u2_u15_u3_n142 ) , .B1( u2_u15_u3_n186 ) , .A( u2_u15_u3_n95 ) );
  INV_X1 u2_u15_u3_U54 (.A( u2_u15_u3_n145 ) , .ZN( u2_u15_u3_n186 ) );
  AOI21_X1 u2_u15_u3_U55 (.B1( u2_u15_u3_n124 ) , .A( u2_u15_u3_n149 ) , .B2( u2_u15_u3_n155 ) , .ZN( u2_u15_u3_n95 ) );
  INV_X1 u2_u15_u3_U56 (.A( u2_u15_u3_n149 ) , .ZN( u2_u15_u3_n169 ) );
  NAND2_X1 u2_u15_u3_U57 (.ZN( u2_u15_u3_n124 ) , .A1( u2_u15_u3_n96 ) , .A2( u2_u15_u3_n97 ) );
  NAND2_X1 u2_u15_u3_U58 (.A2( u2_u15_u3_n100 ) , .ZN( u2_u15_u3_n146 ) , .A1( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U59 (.A1( u2_u15_u3_n101 ) , .ZN( u2_u15_u3_n145 ) , .A2( u2_u15_u3_n99 ) );
  AOI221_X1 u2_u15_u3_U6 (.A( u2_u15_u3_n131 ) , .C2( u2_u15_u3_n132 ) , .C1( u2_u15_u3_n133 ) , .ZN( u2_u15_u3_n134 ) , .B1( u2_u15_u3_n143 ) , .B2( u2_u15_u3_n177 ) );
  NAND2_X1 u2_u15_u3_U60 (.A1( u2_u15_u3_n100 ) , .ZN( u2_u15_u3_n156 ) , .A2( u2_u15_u3_n99 ) );
  NAND2_X1 u2_u15_u3_U61 (.A2( u2_u15_u3_n101 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n148 ) );
  NAND2_X1 u2_u15_u3_U62 (.A1( u2_u15_u3_n100 ) , .A2( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n128 ) );
  NAND2_X1 u2_u15_u3_U63 (.A2( u2_u15_u3_n101 ) , .A1( u2_u15_u3_n102 ) , .ZN( u2_u15_u3_n152 ) );
  NAND2_X1 u2_u15_u3_U64 (.A2( u2_u15_u3_n101 ) , .ZN( u2_u15_u3_n114 ) , .A1( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U65 (.ZN( u2_u15_u3_n107 ) , .A1( u2_u15_u3_n97 ) , .A2( u2_u15_u3_n99 ) );
  NAND2_X1 u2_u15_u3_U66 (.A2( u2_u15_u3_n100 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n113 ) );
  NAND2_X1 u2_u15_u3_U67 (.A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n153 ) , .A2( u2_u15_u3_n97 ) );
  NAND2_X1 u2_u15_u3_U68 (.A2( u2_u15_u3_n103 ) , .A1( u2_u15_u3_n104 ) , .ZN( u2_u15_u3_n130 ) );
  NAND2_X1 u2_u15_u3_U69 (.A2( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n144 ) , .A1( u2_u15_u3_n96 ) );
  OAI22_X1 u2_u15_u3_U7 (.B2( u2_u15_u3_n147 ) , .A2( u2_u15_u3_n148 ) , .ZN( u2_u15_u3_n160 ) , .B1( u2_u15_u3_n165 ) , .A1( u2_u15_u3_n168 ) );
  NAND2_X1 u2_u15_u3_U70 (.A1( u2_u15_u3_n102 ) , .A2( u2_u15_u3_n103 ) , .ZN( u2_u15_u3_n108 ) );
  NOR2_X1 u2_u15_u3_U71 (.A2( u2_u15_X_19 ) , .A1( u2_u15_X_20 ) , .ZN( u2_u15_u3_n99 ) );
  NOR2_X1 u2_u15_u3_U72 (.A2( u2_u15_X_21 ) , .A1( u2_u15_X_24 ) , .ZN( u2_u15_u3_n103 ) );
  NOR2_X1 u2_u15_u3_U73 (.A2( u2_u15_X_24 ) , .A1( u2_u15_u3_n171 ) , .ZN( u2_u15_u3_n97 ) );
  NOR2_X1 u2_u15_u3_U74 (.A2( u2_u15_X_23 ) , .ZN( u2_u15_u3_n141 ) , .A1( u2_u15_u3_n166 ) );
  NOR2_X1 u2_u15_u3_U75 (.A2( u2_u15_X_19 ) , .A1( u2_u15_u3_n172 ) , .ZN( u2_u15_u3_n96 ) );
  NAND2_X1 u2_u15_u3_U76 (.A1( u2_u15_X_22 ) , .A2( u2_u15_X_23 ) , .ZN( u2_u15_u3_n154 ) );
  NAND2_X1 u2_u15_u3_U77 (.A1( u2_u15_X_23 ) , .ZN( u2_u15_u3_n149 ) , .A2( u2_u15_u3_n166 ) );
  NOR2_X1 u2_u15_u3_U78 (.A2( u2_u15_X_22 ) , .A1( u2_u15_X_23 ) , .ZN( u2_u15_u3_n121 ) );
  AND2_X1 u2_u15_u3_U79 (.A1( u2_u15_X_24 ) , .ZN( u2_u15_u3_n101 ) , .A2( u2_u15_u3_n171 ) );
  AND3_X1 u2_u15_u3_U8 (.A3( u2_u15_u3_n144 ) , .A2( u2_u15_u3_n145 ) , .A1( u2_u15_u3_n146 ) , .ZN( u2_u15_u3_n147 ) );
  AND2_X1 u2_u15_u3_U80 (.A1( u2_u15_X_19 ) , .ZN( u2_u15_u3_n102 ) , .A2( u2_u15_u3_n172 ) );
  AND2_X1 u2_u15_u3_U81 (.A1( u2_u15_X_21 ) , .A2( u2_u15_X_24 ) , .ZN( u2_u15_u3_n100 ) );
  AND2_X1 u2_u15_u3_U82 (.A2( u2_u15_X_19 ) , .A1( u2_u15_X_20 ) , .ZN( u2_u15_u3_n104 ) );
  INV_X1 u2_u15_u3_U83 (.A( u2_u15_X_22 ) , .ZN( u2_u15_u3_n166 ) );
  INV_X1 u2_u15_u3_U84 (.A( u2_u15_X_21 ) , .ZN( u2_u15_u3_n171 ) );
  INV_X1 u2_u15_u3_U85 (.A( u2_u15_X_20 ) , .ZN( u2_u15_u3_n172 ) );
  OR4_X1 u2_u15_u3_U86 (.ZN( u2_out15_10 ) , .A4( u2_u15_u3_n136 ) , .A3( u2_u15_u3_n137 ) , .A1( u2_u15_u3_n138 ) , .A2( u2_u15_u3_n139 ) );
  OAI222_X1 u2_u15_u3_U87 (.C1( u2_u15_u3_n128 ) , .ZN( u2_u15_u3_n137 ) , .B1( u2_u15_u3_n148 ) , .A2( u2_u15_u3_n150 ) , .B2( u2_u15_u3_n154 ) , .C2( u2_u15_u3_n164 ) , .A1( u2_u15_u3_n167 ) );
  OAI221_X1 u2_u15_u3_U88 (.A( u2_u15_u3_n134 ) , .B2( u2_u15_u3_n135 ) , .ZN( u2_u15_u3_n136 ) , .C1( u2_u15_u3_n149 ) , .B1( u2_u15_u3_n151 ) , .C2( u2_u15_u3_n183 ) );
  NAND4_X1 u2_u15_u3_U89 (.ZN( u2_out15_1 ) , .A4( u2_u15_u3_n161 ) , .A3( u2_u15_u3_n162 ) , .A2( u2_u15_u3_n163 ) , .A1( u2_u15_u3_n185 ) );
  INV_X1 u2_u15_u3_U9 (.A( u2_u15_u3_n143 ) , .ZN( u2_u15_u3_n168 ) );
  NAND2_X1 u2_u15_u3_U90 (.ZN( u2_u15_u3_n163 ) , .A2( u2_u15_u3_n170 ) , .A1( u2_u15_u3_n176 ) );
  AOI22_X1 u2_u15_u3_U91 (.B2( u2_u15_u3_n140 ) , .B1( u2_u15_u3_n141 ) , .A2( u2_u15_u3_n142 ) , .ZN( u2_u15_u3_n162 ) , .A1( u2_u15_u3_n177 ) );
  NAND4_X1 u2_u15_u3_U92 (.ZN( u2_out15_26 ) , .A4( u2_u15_u3_n109 ) , .A3( u2_u15_u3_n110 ) , .A2( u2_u15_u3_n111 ) , .A1( u2_u15_u3_n173 ) );
  INV_X1 u2_u15_u3_U93 (.ZN( u2_u15_u3_n173 ) , .A( u2_u15_u3_n94 ) );
  OAI21_X1 u2_u15_u3_U94 (.ZN( u2_u15_u3_n111 ) , .B2( u2_u15_u3_n117 ) , .A( u2_u15_u3_n133 ) , .B1( u2_u15_u3_n176 ) );
  NAND4_X1 u2_u15_u3_U95 (.ZN( u2_out15_20 ) , .A4( u2_u15_u3_n122 ) , .A3( u2_u15_u3_n123 ) , .A1( u2_u15_u3_n175 ) , .A2( u2_u15_u3_n180 ) );
  INV_X1 u2_u15_u3_U96 (.A( u2_u15_u3_n126 ) , .ZN( u2_u15_u3_n180 ) );
  INV_X1 u2_u15_u3_U97 (.A( u2_u15_u3_n112 ) , .ZN( u2_u15_u3_n175 ) );
  NAND3_X1 u2_u15_u3_U98 (.A1( u2_u15_u3_n114 ) , .ZN( u2_u15_u3_n115 ) , .A2( u2_u15_u3_n145 ) , .A3( u2_u15_u3_n153 ) );
  NAND3_X1 u2_u15_u3_U99 (.ZN( u2_u15_u3_n129 ) , .A2( u2_u15_u3_n144 ) , .A1( u2_u15_u3_n153 ) , .A3( u2_u15_u3_n182 ) );
  XOR2_X1 u2_u1_U1 (.B( u2_K2_9 ) , .A( u2_R0_6 ) , .Z( u2_u1_X_9 ) );
  XOR2_X1 u2_u1_U2 (.B( u2_K2_8 ) , .A( u2_R0_5 ) , .Z( u2_u1_X_8 ) );
  XOR2_X1 u2_u1_U3 (.B( u2_K2_7 ) , .A( u2_R0_4 ) , .Z( u2_u1_X_7 ) );
  XOR2_X1 u2_u1_U33 (.B( u2_K2_24 ) , .A( u2_R0_17 ) , .Z( u2_u1_X_24 ) );
  XOR2_X1 u2_u1_U34 (.B( u2_K2_23 ) , .A( u2_R0_16 ) , .Z( u2_u1_X_23 ) );
  XOR2_X1 u2_u1_U35 (.B( u2_K2_22 ) , .A( u2_R0_15 ) , .Z( u2_u1_X_22 ) );
  XOR2_X1 u2_u1_U36 (.B( u2_K2_21 ) , .A( u2_R0_14 ) , .Z( u2_u1_X_21 ) );
  XOR2_X1 u2_u1_U37 (.B( u2_K2_20 ) , .A( u2_R0_13 ) , .Z( u2_u1_X_20 ) );
  XOR2_X1 u2_u1_U39 (.B( u2_K2_19 ) , .A( u2_R0_12 ) , .Z( u2_u1_X_19 ) );
  XOR2_X1 u2_u1_U40 (.B( u2_K2_18 ) , .A( u2_R0_13 ) , .Z( u2_u1_X_18 ) );
  XOR2_X1 u2_u1_U41 (.B( u2_K2_17 ) , .A( u2_R0_12 ) , .Z( u2_u1_X_17 ) );
  XOR2_X1 u2_u1_U42 (.B( u2_K2_16 ) , .A( u2_R0_11 ) , .Z( u2_u1_X_16 ) );
  XOR2_X1 u2_u1_U43 (.B( u2_K2_15 ) , .A( u2_R0_10 ) , .Z( u2_u1_X_15 ) );
  XOR2_X1 u2_u1_U44 (.B( u2_K2_14 ) , .A( u2_R0_9 ) , .Z( u2_u1_X_14 ) );
  XOR2_X1 u2_u1_U45 (.B( u2_K2_13 ) , .A( u2_R0_8 ) , .Z( u2_u1_X_13 ) );
  XOR2_X1 u2_u1_U46 (.B( u2_K2_12 ) , .A( u2_R0_9 ) , .Z( u2_u1_X_12 ) );
  XOR2_X1 u2_u1_U47 (.B( u2_K2_11 ) , .A( u2_R0_8 ) , .Z( u2_u1_X_11 ) );
  XOR2_X1 u2_u1_U48 (.B( u2_K2_10 ) , .A( u2_R0_7 ) , .Z( u2_u1_X_10 ) );
  NOR2_X1 u2_u1_u1_U10 (.A1( u2_u1_u1_n112 ) , .A2( u2_u1_u1_n116 ) , .ZN( u2_u1_u1_n118 ) );
  NAND3_X1 u2_u1_u1_U100 (.ZN( u2_u1_u1_n113 ) , .A1( u2_u1_u1_n120 ) , .A3( u2_u1_u1_n133 ) , .A2( u2_u1_u1_n155 ) );
  OAI21_X1 u2_u1_u1_U11 (.ZN( u2_u1_u1_n101 ) , .B1( u2_u1_u1_n141 ) , .A( u2_u1_u1_n146 ) , .B2( u2_u1_u1_n183 ) );
  AOI21_X1 u2_u1_u1_U12 (.B2( u2_u1_u1_n155 ) , .B1( u2_u1_u1_n156 ) , .ZN( u2_u1_u1_n157 ) , .A( u2_u1_u1_n174 ) );
  OR4_X1 u2_u1_u1_U13 (.A4( u2_u1_u1_n106 ) , .A3( u2_u1_u1_n107 ) , .ZN( u2_u1_u1_n108 ) , .A1( u2_u1_u1_n117 ) , .A2( u2_u1_u1_n184 ) );
  AOI21_X1 u2_u1_u1_U14 (.ZN( u2_u1_u1_n106 ) , .A( u2_u1_u1_n112 ) , .B1( u2_u1_u1_n154 ) , .B2( u2_u1_u1_n156 ) );
  INV_X1 u2_u1_u1_U15 (.A( u2_u1_u1_n101 ) , .ZN( u2_u1_u1_n184 ) );
  AOI21_X1 u2_u1_u1_U16 (.ZN( u2_u1_u1_n107 ) , .B1( u2_u1_u1_n134 ) , .B2( u2_u1_u1_n149 ) , .A( u2_u1_u1_n174 ) );
  NAND2_X1 u2_u1_u1_U17 (.ZN( u2_u1_u1_n140 ) , .A2( u2_u1_u1_n150 ) , .A1( u2_u1_u1_n155 ) );
  NAND2_X1 u2_u1_u1_U18 (.A1( u2_u1_u1_n131 ) , .ZN( u2_u1_u1_n147 ) , .A2( u2_u1_u1_n153 ) );
  INV_X1 u2_u1_u1_U19 (.A( u2_u1_u1_n139 ) , .ZN( u2_u1_u1_n174 ) );
  INV_X1 u2_u1_u1_U20 (.A( u2_u1_u1_n112 ) , .ZN( u2_u1_u1_n171 ) );
  NAND2_X1 u2_u1_u1_U21 (.ZN( u2_u1_u1_n141 ) , .A1( u2_u1_u1_n153 ) , .A2( u2_u1_u1_n156 ) );
  AND2_X1 u2_u1_u1_U22 (.A1( u2_u1_u1_n123 ) , .ZN( u2_u1_u1_n134 ) , .A2( u2_u1_u1_n161 ) );
  NAND2_X1 u2_u1_u1_U23 (.A2( u2_u1_u1_n115 ) , .A1( u2_u1_u1_n116 ) , .ZN( u2_u1_u1_n148 ) );
  NAND2_X1 u2_u1_u1_U24 (.A2( u2_u1_u1_n133 ) , .A1( u2_u1_u1_n135 ) , .ZN( u2_u1_u1_n159 ) );
  NAND2_X1 u2_u1_u1_U25 (.A2( u2_u1_u1_n115 ) , .A1( u2_u1_u1_n120 ) , .ZN( u2_u1_u1_n132 ) );
  INV_X1 u2_u1_u1_U26 (.A( u2_u1_u1_n154 ) , .ZN( u2_u1_u1_n178 ) );
  INV_X1 u2_u1_u1_U27 (.A( u2_u1_u1_n151 ) , .ZN( u2_u1_u1_n183 ) );
  AND2_X1 u2_u1_u1_U28 (.A1( u2_u1_u1_n129 ) , .A2( u2_u1_u1_n133 ) , .ZN( u2_u1_u1_n149 ) );
  INV_X1 u2_u1_u1_U29 (.A( u2_u1_u1_n131 ) , .ZN( u2_u1_u1_n180 ) );
  INV_X1 u2_u1_u1_U3 (.A( u2_u1_u1_n159 ) , .ZN( u2_u1_u1_n182 ) );
  AOI221_X1 u2_u1_u1_U30 (.B1( u2_u1_u1_n140 ) , .ZN( u2_u1_u1_n167 ) , .B2( u2_u1_u1_n172 ) , .C2( u2_u1_u1_n175 ) , .C1( u2_u1_u1_n178 ) , .A( u2_u1_u1_n188 ) );
  INV_X1 u2_u1_u1_U31 (.ZN( u2_u1_u1_n188 ) , .A( u2_u1_u1_n97 ) );
  AOI211_X1 u2_u1_u1_U32 (.A( u2_u1_u1_n118 ) , .C1( u2_u1_u1_n132 ) , .C2( u2_u1_u1_n139 ) , .B( u2_u1_u1_n96 ) , .ZN( u2_u1_u1_n97 ) );
  AOI21_X1 u2_u1_u1_U33 (.B2( u2_u1_u1_n121 ) , .B1( u2_u1_u1_n135 ) , .A( u2_u1_u1_n152 ) , .ZN( u2_u1_u1_n96 ) );
  OAI221_X1 u2_u1_u1_U34 (.A( u2_u1_u1_n119 ) , .C2( u2_u1_u1_n129 ) , .ZN( u2_u1_u1_n138 ) , .B2( u2_u1_u1_n152 ) , .C1( u2_u1_u1_n174 ) , .B1( u2_u1_u1_n187 ) );
  INV_X1 u2_u1_u1_U35 (.A( u2_u1_u1_n148 ) , .ZN( u2_u1_u1_n187 ) );
  AOI211_X1 u2_u1_u1_U36 (.B( u2_u1_u1_n117 ) , .A( u2_u1_u1_n118 ) , .ZN( u2_u1_u1_n119 ) , .C2( u2_u1_u1_n146 ) , .C1( u2_u1_u1_n159 ) );
  NOR2_X1 u2_u1_u1_U37 (.A1( u2_u1_u1_n168 ) , .A2( u2_u1_u1_n176 ) , .ZN( u2_u1_u1_n98 ) );
  AOI211_X1 u2_u1_u1_U38 (.B( u2_u1_u1_n162 ) , .A( u2_u1_u1_n163 ) , .C2( u2_u1_u1_n164 ) , .ZN( u2_u1_u1_n165 ) , .C1( u2_u1_u1_n171 ) );
  AOI21_X1 u2_u1_u1_U39 (.A( u2_u1_u1_n160 ) , .B2( u2_u1_u1_n161 ) , .ZN( u2_u1_u1_n162 ) , .B1( u2_u1_u1_n182 ) );
  AOI221_X1 u2_u1_u1_U4 (.A( u2_u1_u1_n138 ) , .C2( u2_u1_u1_n139 ) , .C1( u2_u1_u1_n140 ) , .B2( u2_u1_u1_n141 ) , .ZN( u2_u1_u1_n142 ) , .B1( u2_u1_u1_n175 ) );
  OR2_X1 u2_u1_u1_U40 (.A2( u2_u1_u1_n157 ) , .A1( u2_u1_u1_n158 ) , .ZN( u2_u1_u1_n163 ) );
  OAI21_X1 u2_u1_u1_U41 (.B2( u2_u1_u1_n123 ) , .ZN( u2_u1_u1_n145 ) , .B1( u2_u1_u1_n160 ) , .A( u2_u1_u1_n185 ) );
  INV_X1 u2_u1_u1_U42 (.A( u2_u1_u1_n122 ) , .ZN( u2_u1_u1_n185 ) );
  AOI21_X1 u2_u1_u1_U43 (.B2( u2_u1_u1_n120 ) , .B1( u2_u1_u1_n121 ) , .ZN( u2_u1_u1_n122 ) , .A( u2_u1_u1_n128 ) );
  NAND2_X1 u2_u1_u1_U44 (.A1( u2_u1_u1_n128 ) , .ZN( u2_u1_u1_n146 ) , .A2( u2_u1_u1_n160 ) );
  NAND2_X1 u2_u1_u1_U45 (.A2( u2_u1_u1_n112 ) , .ZN( u2_u1_u1_n139 ) , .A1( u2_u1_u1_n152 ) );
  NAND2_X1 u2_u1_u1_U46 (.A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n156 ) , .A2( u2_u1_u1_n99 ) );
  NOR2_X1 u2_u1_u1_U47 (.ZN( u2_u1_u1_n117 ) , .A1( u2_u1_u1_n121 ) , .A2( u2_u1_u1_n160 ) );
  AOI21_X1 u2_u1_u1_U48 (.A( u2_u1_u1_n128 ) , .B2( u2_u1_u1_n129 ) , .ZN( u2_u1_u1_n130 ) , .B1( u2_u1_u1_n150 ) );
  NAND2_X1 u2_u1_u1_U49 (.ZN( u2_u1_u1_n112 ) , .A1( u2_u1_u1_n169 ) , .A2( u2_u1_u1_n170 ) );
  AOI211_X1 u2_u1_u1_U5 (.ZN( u2_u1_u1_n124 ) , .A( u2_u1_u1_n138 ) , .C2( u2_u1_u1_n139 ) , .B( u2_u1_u1_n145 ) , .C1( u2_u1_u1_n147 ) );
  NAND2_X1 u2_u1_u1_U50 (.ZN( u2_u1_u1_n129 ) , .A2( u2_u1_u1_n95 ) , .A1( u2_u1_u1_n98 ) );
  NAND2_X1 u2_u1_u1_U51 (.A1( u2_u1_u1_n102 ) , .ZN( u2_u1_u1_n154 ) , .A2( u2_u1_u1_n99 ) );
  NAND2_X1 u2_u1_u1_U52 (.A2( u2_u1_u1_n100 ) , .ZN( u2_u1_u1_n135 ) , .A1( u2_u1_u1_n99 ) );
  AOI21_X1 u2_u1_u1_U53 (.A( u2_u1_u1_n152 ) , .B2( u2_u1_u1_n153 ) , .B1( u2_u1_u1_n154 ) , .ZN( u2_u1_u1_n158 ) );
  INV_X1 u2_u1_u1_U54 (.A( u2_u1_u1_n160 ) , .ZN( u2_u1_u1_n175 ) );
  NAND2_X1 u2_u1_u1_U55 (.A1( u2_u1_u1_n100 ) , .ZN( u2_u1_u1_n116 ) , .A2( u2_u1_u1_n95 ) );
  NAND2_X1 u2_u1_u1_U56 (.A1( u2_u1_u1_n102 ) , .ZN( u2_u1_u1_n131 ) , .A2( u2_u1_u1_n95 ) );
  NAND2_X1 u2_u1_u1_U57 (.A2( u2_u1_u1_n104 ) , .ZN( u2_u1_u1_n121 ) , .A1( u2_u1_u1_n98 ) );
  NAND2_X1 u2_u1_u1_U58 (.A1( u2_u1_u1_n103 ) , .ZN( u2_u1_u1_n153 ) , .A2( u2_u1_u1_n98 ) );
  NAND2_X1 u2_u1_u1_U59 (.A2( u2_u1_u1_n104 ) , .A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n133 ) );
  AOI22_X1 u2_u1_u1_U6 (.B2( u2_u1_u1_n113 ) , .A2( u2_u1_u1_n114 ) , .ZN( u2_u1_u1_n125 ) , .A1( u2_u1_u1_n171 ) , .B1( u2_u1_u1_n173 ) );
  NAND2_X1 u2_u1_u1_U60 (.ZN( u2_u1_u1_n150 ) , .A2( u2_u1_u1_n98 ) , .A1( u2_u1_u1_n99 ) );
  NAND2_X1 u2_u1_u1_U61 (.A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n155 ) , .A2( u2_u1_u1_n95 ) );
  OAI21_X1 u2_u1_u1_U62 (.ZN( u2_u1_u1_n109 ) , .B1( u2_u1_u1_n129 ) , .B2( u2_u1_u1_n160 ) , .A( u2_u1_u1_n167 ) );
  NAND2_X1 u2_u1_u1_U63 (.A2( u2_u1_u1_n100 ) , .A1( u2_u1_u1_n103 ) , .ZN( u2_u1_u1_n120 ) );
  NAND2_X1 u2_u1_u1_U64 (.A1( u2_u1_u1_n102 ) , .A2( u2_u1_u1_n104 ) , .ZN( u2_u1_u1_n115 ) );
  NAND2_X1 u2_u1_u1_U65 (.A2( u2_u1_u1_n100 ) , .A1( u2_u1_u1_n104 ) , .ZN( u2_u1_u1_n151 ) );
  NAND2_X1 u2_u1_u1_U66 (.A2( u2_u1_u1_n103 ) , .A1( u2_u1_u1_n105 ) , .ZN( u2_u1_u1_n161 ) );
  INV_X1 u2_u1_u1_U67 (.A( u2_u1_u1_n152 ) , .ZN( u2_u1_u1_n173 ) );
  INV_X1 u2_u1_u1_U68 (.A( u2_u1_u1_n128 ) , .ZN( u2_u1_u1_n172 ) );
  NAND2_X1 u2_u1_u1_U69 (.A2( u2_u1_u1_n102 ) , .A1( u2_u1_u1_n103 ) , .ZN( u2_u1_u1_n123 ) );
  NAND2_X1 u2_u1_u1_U7 (.ZN( u2_u1_u1_n114 ) , .A1( u2_u1_u1_n134 ) , .A2( u2_u1_u1_n156 ) );
  NOR2_X1 u2_u1_u1_U70 (.A2( u2_u1_X_7 ) , .A1( u2_u1_X_8 ) , .ZN( u2_u1_u1_n95 ) );
  NOR2_X1 u2_u1_u1_U71 (.A1( u2_u1_X_12 ) , .A2( u2_u1_X_9 ) , .ZN( u2_u1_u1_n100 ) );
  NOR2_X1 u2_u1_u1_U72 (.A2( u2_u1_X_8 ) , .A1( u2_u1_u1_n177 ) , .ZN( u2_u1_u1_n99 ) );
  NOR2_X1 u2_u1_u1_U73 (.A2( u2_u1_X_12 ) , .ZN( u2_u1_u1_n102 ) , .A1( u2_u1_u1_n176 ) );
  NOR2_X1 u2_u1_u1_U74 (.A2( u2_u1_X_9 ) , .ZN( u2_u1_u1_n105 ) , .A1( u2_u1_u1_n168 ) );
  NAND2_X1 u2_u1_u1_U75 (.A1( u2_u1_X_10 ) , .ZN( u2_u1_u1_n160 ) , .A2( u2_u1_u1_n169 ) );
  NAND2_X1 u2_u1_u1_U76 (.A2( u2_u1_X_10 ) , .A1( u2_u1_X_11 ) , .ZN( u2_u1_u1_n152 ) );
  NAND2_X1 u2_u1_u1_U77 (.A1( u2_u1_X_11 ) , .ZN( u2_u1_u1_n128 ) , .A2( u2_u1_u1_n170 ) );
  AND2_X1 u2_u1_u1_U78 (.A2( u2_u1_X_7 ) , .A1( u2_u1_X_8 ) , .ZN( u2_u1_u1_n104 ) );
  AND2_X1 u2_u1_u1_U79 (.A1( u2_u1_X_8 ) , .ZN( u2_u1_u1_n103 ) , .A2( u2_u1_u1_n177 ) );
  AOI22_X1 u2_u1_u1_U8 (.B2( u2_u1_u1_n136 ) , .A2( u2_u1_u1_n137 ) , .ZN( u2_u1_u1_n143 ) , .A1( u2_u1_u1_n171 ) , .B1( u2_u1_u1_n173 ) );
  INV_X1 u2_u1_u1_U80 (.A( u2_u1_X_10 ) , .ZN( u2_u1_u1_n170 ) );
  INV_X1 u2_u1_u1_U81 (.A( u2_u1_X_9 ) , .ZN( u2_u1_u1_n176 ) );
  INV_X1 u2_u1_u1_U82 (.A( u2_u1_X_11 ) , .ZN( u2_u1_u1_n169 ) );
  INV_X1 u2_u1_u1_U83 (.A( u2_u1_X_12 ) , .ZN( u2_u1_u1_n168 ) );
  INV_X1 u2_u1_u1_U84 (.A( u2_u1_X_7 ) , .ZN( u2_u1_u1_n177 ) );
  NAND4_X1 u2_u1_u1_U85 (.ZN( u2_out1_18 ) , .A4( u2_u1_u1_n165 ) , .A3( u2_u1_u1_n166 ) , .A1( u2_u1_u1_n167 ) , .A2( u2_u1_u1_n186 ) );
  AOI22_X1 u2_u1_u1_U86 (.B2( u2_u1_u1_n146 ) , .B1( u2_u1_u1_n147 ) , .A2( u2_u1_u1_n148 ) , .ZN( u2_u1_u1_n166 ) , .A1( u2_u1_u1_n172 ) );
  INV_X1 u2_u1_u1_U87 (.A( u2_u1_u1_n145 ) , .ZN( u2_u1_u1_n186 ) );
  NAND4_X1 u2_u1_u1_U88 (.ZN( u2_out1_2 ) , .A4( u2_u1_u1_n142 ) , .A3( u2_u1_u1_n143 ) , .A2( u2_u1_u1_n144 ) , .A1( u2_u1_u1_n179 ) );
  INV_X1 u2_u1_u1_U89 (.A( u2_u1_u1_n130 ) , .ZN( u2_u1_u1_n179 ) );
  INV_X1 u2_u1_u1_U9 (.A( u2_u1_u1_n147 ) , .ZN( u2_u1_u1_n181 ) );
  OAI21_X1 u2_u1_u1_U90 (.B2( u2_u1_u1_n132 ) , .ZN( u2_u1_u1_n144 ) , .A( u2_u1_u1_n146 ) , .B1( u2_u1_u1_n180 ) );
  NAND4_X1 u2_u1_u1_U91 (.ZN( u2_out1_28 ) , .A4( u2_u1_u1_n124 ) , .A3( u2_u1_u1_n125 ) , .A2( u2_u1_u1_n126 ) , .A1( u2_u1_u1_n127 ) );
  OAI21_X1 u2_u1_u1_U92 (.ZN( u2_u1_u1_n127 ) , .B2( u2_u1_u1_n139 ) , .B1( u2_u1_u1_n175 ) , .A( u2_u1_u1_n183 ) );
  OAI21_X1 u2_u1_u1_U93 (.ZN( u2_u1_u1_n126 ) , .B2( u2_u1_u1_n140 ) , .A( u2_u1_u1_n146 ) , .B1( u2_u1_u1_n178 ) );
  OR4_X1 u2_u1_u1_U94 (.ZN( u2_out1_13 ) , .A4( u2_u1_u1_n108 ) , .A3( u2_u1_u1_n109 ) , .A2( u2_u1_u1_n110 ) , .A1( u2_u1_u1_n111 ) );
  AOI21_X1 u2_u1_u1_U95 (.ZN( u2_u1_u1_n111 ) , .A( u2_u1_u1_n128 ) , .B2( u2_u1_u1_n131 ) , .B1( u2_u1_u1_n135 ) );
  AOI21_X1 u2_u1_u1_U96 (.ZN( u2_u1_u1_n110 ) , .A( u2_u1_u1_n116 ) , .B1( u2_u1_u1_n152 ) , .B2( u2_u1_u1_n160 ) );
  NAND3_X1 u2_u1_u1_U97 (.A3( u2_u1_u1_n149 ) , .A2( u2_u1_u1_n150 ) , .A1( u2_u1_u1_n151 ) , .ZN( u2_u1_u1_n164 ) );
  NAND3_X1 u2_u1_u1_U98 (.A3( u2_u1_u1_n134 ) , .A2( u2_u1_u1_n135 ) , .ZN( u2_u1_u1_n136 ) , .A1( u2_u1_u1_n151 ) );
  NAND3_X1 u2_u1_u1_U99 (.A1( u2_u1_u1_n133 ) , .ZN( u2_u1_u1_n137 ) , .A2( u2_u1_u1_n154 ) , .A3( u2_u1_u1_n181 ) );
  OAI22_X1 u2_u1_u2_U10 (.ZN( u2_u1_u2_n109 ) , .A2( u2_u1_u2_n113 ) , .B2( u2_u1_u2_n133 ) , .B1( u2_u1_u2_n167 ) , .A1( u2_u1_u2_n168 ) );
  NAND3_X1 u2_u1_u2_U100 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n104 ) , .A3( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n98 ) );
  OAI22_X1 u2_u1_u2_U11 (.B1( u2_u1_u2_n151 ) , .A2( u2_u1_u2_n152 ) , .A1( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n160 ) , .B2( u2_u1_u2_n168 ) );
  NOR3_X1 u2_u1_u2_U12 (.A1( u2_u1_u2_n150 ) , .ZN( u2_u1_u2_n151 ) , .A3( u2_u1_u2_n175 ) , .A2( u2_u1_u2_n188 ) );
  AOI21_X1 u2_u1_u2_U13 (.ZN( u2_u1_u2_n144 ) , .B2( u2_u1_u2_n155 ) , .A( u2_u1_u2_n172 ) , .B1( u2_u1_u2_n185 ) );
  AOI21_X1 u2_u1_u2_U14 (.B2( u2_u1_u2_n143 ) , .ZN( u2_u1_u2_n145 ) , .B1( u2_u1_u2_n152 ) , .A( u2_u1_u2_n171 ) );
  AOI21_X1 u2_u1_u2_U15 (.B2( u2_u1_u2_n120 ) , .B1( u2_u1_u2_n121 ) , .ZN( u2_u1_u2_n126 ) , .A( u2_u1_u2_n167 ) );
  INV_X1 u2_u1_u2_U16 (.A( u2_u1_u2_n156 ) , .ZN( u2_u1_u2_n171 ) );
  INV_X1 u2_u1_u2_U17 (.A( u2_u1_u2_n120 ) , .ZN( u2_u1_u2_n188 ) );
  NAND2_X1 u2_u1_u2_U18 (.A2( u2_u1_u2_n122 ) , .ZN( u2_u1_u2_n150 ) , .A1( u2_u1_u2_n152 ) );
  INV_X1 u2_u1_u2_U19 (.A( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n170 ) );
  INV_X1 u2_u1_u2_U20 (.A( u2_u1_u2_n137 ) , .ZN( u2_u1_u2_n173 ) );
  NAND2_X1 u2_u1_u2_U21 (.A1( u2_u1_u2_n132 ) , .A2( u2_u1_u2_n139 ) , .ZN( u2_u1_u2_n157 ) );
  INV_X1 u2_u1_u2_U22 (.A( u2_u1_u2_n113 ) , .ZN( u2_u1_u2_n178 ) );
  INV_X1 u2_u1_u2_U23 (.A( u2_u1_u2_n139 ) , .ZN( u2_u1_u2_n175 ) );
  INV_X1 u2_u1_u2_U24 (.A( u2_u1_u2_n155 ) , .ZN( u2_u1_u2_n181 ) );
  INV_X1 u2_u1_u2_U25 (.A( u2_u1_u2_n119 ) , .ZN( u2_u1_u2_n177 ) );
  INV_X1 u2_u1_u2_U26 (.A( u2_u1_u2_n116 ) , .ZN( u2_u1_u2_n180 ) );
  INV_X1 u2_u1_u2_U27 (.A( u2_u1_u2_n131 ) , .ZN( u2_u1_u2_n179 ) );
  INV_X1 u2_u1_u2_U28 (.A( u2_u1_u2_n154 ) , .ZN( u2_u1_u2_n176 ) );
  NAND2_X1 u2_u1_u2_U29 (.A2( u2_u1_u2_n116 ) , .A1( u2_u1_u2_n117 ) , .ZN( u2_u1_u2_n118 ) );
  NOR2_X1 u2_u1_u2_U3 (.ZN( u2_u1_u2_n121 ) , .A2( u2_u1_u2_n177 ) , .A1( u2_u1_u2_n180 ) );
  INV_X1 u2_u1_u2_U30 (.A( u2_u1_u2_n132 ) , .ZN( u2_u1_u2_n182 ) );
  INV_X1 u2_u1_u2_U31 (.A( u2_u1_u2_n158 ) , .ZN( u2_u1_u2_n183 ) );
  OAI21_X1 u2_u1_u2_U32 (.A( u2_u1_u2_n156 ) , .B1( u2_u1_u2_n157 ) , .ZN( u2_u1_u2_n158 ) , .B2( u2_u1_u2_n179 ) );
  NOR2_X1 u2_u1_u2_U33 (.ZN( u2_u1_u2_n156 ) , .A1( u2_u1_u2_n166 ) , .A2( u2_u1_u2_n169 ) );
  NOR2_X1 u2_u1_u2_U34 (.A2( u2_u1_u2_n114 ) , .ZN( u2_u1_u2_n137 ) , .A1( u2_u1_u2_n140 ) );
  NOR2_X1 u2_u1_u2_U35 (.A2( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n153 ) , .A1( u2_u1_u2_n156 ) );
  AOI211_X1 u2_u1_u2_U36 (.ZN( u2_u1_u2_n130 ) , .C1( u2_u1_u2_n138 ) , .C2( u2_u1_u2_n179 ) , .B( u2_u1_u2_n96 ) , .A( u2_u1_u2_n97 ) );
  OAI22_X1 u2_u1_u2_U37 (.B1( u2_u1_u2_n133 ) , .A2( u2_u1_u2_n137 ) , .A1( u2_u1_u2_n152 ) , .B2( u2_u1_u2_n168 ) , .ZN( u2_u1_u2_n97 ) );
  OAI221_X1 u2_u1_u2_U38 (.B1( u2_u1_u2_n113 ) , .C1( u2_u1_u2_n132 ) , .A( u2_u1_u2_n149 ) , .B2( u2_u1_u2_n171 ) , .C2( u2_u1_u2_n172 ) , .ZN( u2_u1_u2_n96 ) );
  OAI221_X1 u2_u1_u2_U39 (.A( u2_u1_u2_n115 ) , .C2( u2_u1_u2_n123 ) , .B2( u2_u1_u2_n143 ) , .B1( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n163 ) , .C1( u2_u1_u2_n168 ) );
  INV_X1 u2_u1_u2_U4 (.A( u2_u1_u2_n134 ) , .ZN( u2_u1_u2_n185 ) );
  OAI21_X1 u2_u1_u2_U40 (.A( u2_u1_u2_n114 ) , .ZN( u2_u1_u2_n115 ) , .B1( u2_u1_u2_n176 ) , .B2( u2_u1_u2_n178 ) );
  OAI221_X1 u2_u1_u2_U41 (.A( u2_u1_u2_n135 ) , .B2( u2_u1_u2_n136 ) , .B1( u2_u1_u2_n137 ) , .ZN( u2_u1_u2_n162 ) , .C2( u2_u1_u2_n167 ) , .C1( u2_u1_u2_n185 ) );
  AND3_X1 u2_u1_u2_U42 (.A3( u2_u1_u2_n131 ) , .A2( u2_u1_u2_n132 ) , .A1( u2_u1_u2_n133 ) , .ZN( u2_u1_u2_n136 ) );
  AOI22_X1 u2_u1_u2_U43 (.ZN( u2_u1_u2_n135 ) , .B1( u2_u1_u2_n140 ) , .A1( u2_u1_u2_n156 ) , .B2( u2_u1_u2_n180 ) , .A2( u2_u1_u2_n188 ) );
  AOI21_X1 u2_u1_u2_U44 (.ZN( u2_u1_u2_n149 ) , .B1( u2_u1_u2_n173 ) , .B2( u2_u1_u2_n188 ) , .A( u2_u1_u2_n95 ) );
  AND3_X1 u2_u1_u2_U45 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n104 ) , .A3( u2_u1_u2_n156 ) , .ZN( u2_u1_u2_n95 ) );
  OAI21_X1 u2_u1_u2_U46 (.A( u2_u1_u2_n101 ) , .B2( u2_u1_u2_n121 ) , .B1( u2_u1_u2_n153 ) , .ZN( u2_u1_u2_n164 ) );
  NAND2_X1 u2_u1_u2_U47 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n107 ) , .ZN( u2_u1_u2_n155 ) );
  NAND2_X1 u2_u1_u2_U48 (.A2( u2_u1_u2_n105 ) , .A1( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n143 ) );
  NAND2_X1 u2_u1_u2_U49 (.A1( u2_u1_u2_n104 ) , .A2( u2_u1_u2_n106 ) , .ZN( u2_u1_u2_n152 ) );
  INV_X1 u2_u1_u2_U5 (.A( u2_u1_u2_n150 ) , .ZN( u2_u1_u2_n184 ) );
  NAND2_X1 u2_u1_u2_U50 (.A1( u2_u1_u2_n100 ) , .A2( u2_u1_u2_n105 ) , .ZN( u2_u1_u2_n132 ) );
  INV_X1 u2_u1_u2_U51 (.A( u2_u1_u2_n140 ) , .ZN( u2_u1_u2_n168 ) );
  INV_X1 u2_u1_u2_U52 (.A( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n167 ) );
  OAI21_X1 u2_u1_u2_U53 (.A( u2_u1_u2_n141 ) , .B2( u2_u1_u2_n142 ) , .ZN( u2_u1_u2_n146 ) , .B1( u2_u1_u2_n153 ) );
  OAI21_X1 u2_u1_u2_U54 (.A( u2_u1_u2_n140 ) , .ZN( u2_u1_u2_n141 ) , .B1( u2_u1_u2_n176 ) , .B2( u2_u1_u2_n177 ) );
  NOR3_X1 u2_u1_u2_U55 (.ZN( u2_u1_u2_n142 ) , .A3( u2_u1_u2_n175 ) , .A2( u2_u1_u2_n178 ) , .A1( u2_u1_u2_n181 ) );
  NAND2_X1 u2_u1_u2_U56 (.A1( u2_u1_u2_n102 ) , .A2( u2_u1_u2_n106 ) , .ZN( u2_u1_u2_n113 ) );
  NAND2_X1 u2_u1_u2_U57 (.A1( u2_u1_u2_n106 ) , .A2( u2_u1_u2_n107 ) , .ZN( u2_u1_u2_n131 ) );
  NAND2_X1 u2_u1_u2_U58 (.A1( u2_u1_u2_n103 ) , .A2( u2_u1_u2_n107 ) , .ZN( u2_u1_u2_n139 ) );
  NAND2_X1 u2_u1_u2_U59 (.A1( u2_u1_u2_n103 ) , .A2( u2_u1_u2_n105 ) , .ZN( u2_u1_u2_n133 ) );
  NOR4_X1 u2_u1_u2_U6 (.A4( u2_u1_u2_n124 ) , .A3( u2_u1_u2_n125 ) , .A2( u2_u1_u2_n126 ) , .A1( u2_u1_u2_n127 ) , .ZN( u2_u1_u2_n128 ) );
  NAND2_X1 u2_u1_u2_U60 (.A1( u2_u1_u2_n102 ) , .A2( u2_u1_u2_n103 ) , .ZN( u2_u1_u2_n154 ) );
  NAND2_X1 u2_u1_u2_U61 (.A2( u2_u1_u2_n103 ) , .A1( u2_u1_u2_n104 ) , .ZN( u2_u1_u2_n119 ) );
  NAND2_X1 u2_u1_u2_U62 (.A2( u2_u1_u2_n107 ) , .A1( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n123 ) );
  NAND2_X1 u2_u1_u2_U63 (.A1( u2_u1_u2_n104 ) , .A2( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n122 ) );
  INV_X1 u2_u1_u2_U64 (.A( u2_u1_u2_n114 ) , .ZN( u2_u1_u2_n172 ) );
  NAND2_X1 u2_u1_u2_U65 (.A2( u2_u1_u2_n100 ) , .A1( u2_u1_u2_n102 ) , .ZN( u2_u1_u2_n116 ) );
  NAND2_X1 u2_u1_u2_U66 (.A1( u2_u1_u2_n102 ) , .A2( u2_u1_u2_n108 ) , .ZN( u2_u1_u2_n120 ) );
  NAND2_X1 u2_u1_u2_U67 (.A2( u2_u1_u2_n105 ) , .A1( u2_u1_u2_n106 ) , .ZN( u2_u1_u2_n117 ) );
  INV_X1 u2_u1_u2_U68 (.ZN( u2_u1_u2_n187 ) , .A( u2_u1_u2_n99 ) );
  OAI21_X1 u2_u1_u2_U69 (.B1( u2_u1_u2_n137 ) , .B2( u2_u1_u2_n143 ) , .A( u2_u1_u2_n98 ) , .ZN( u2_u1_u2_n99 ) );
  AOI21_X1 u2_u1_u2_U7 (.B2( u2_u1_u2_n119 ) , .ZN( u2_u1_u2_n127 ) , .A( u2_u1_u2_n137 ) , .B1( u2_u1_u2_n155 ) );
  NOR2_X1 u2_u1_u2_U70 (.A2( u2_u1_X_16 ) , .ZN( u2_u1_u2_n140 ) , .A1( u2_u1_u2_n166 ) );
  NOR2_X1 u2_u1_u2_U71 (.A2( u2_u1_X_13 ) , .A1( u2_u1_X_14 ) , .ZN( u2_u1_u2_n100 ) );
  NOR2_X1 u2_u1_u2_U72 (.A2( u2_u1_X_16 ) , .A1( u2_u1_X_17 ) , .ZN( u2_u1_u2_n138 ) );
  NOR2_X1 u2_u1_u2_U73 (.A2( u2_u1_X_15 ) , .A1( u2_u1_X_18 ) , .ZN( u2_u1_u2_n104 ) );
  NOR2_X1 u2_u1_u2_U74 (.A2( u2_u1_X_14 ) , .ZN( u2_u1_u2_n103 ) , .A1( u2_u1_u2_n174 ) );
  NOR2_X1 u2_u1_u2_U75 (.A2( u2_u1_X_15 ) , .ZN( u2_u1_u2_n102 ) , .A1( u2_u1_u2_n165 ) );
  NOR2_X1 u2_u1_u2_U76 (.A2( u2_u1_X_17 ) , .ZN( u2_u1_u2_n114 ) , .A1( u2_u1_u2_n169 ) );
  AND2_X1 u2_u1_u2_U77 (.A1( u2_u1_X_15 ) , .ZN( u2_u1_u2_n105 ) , .A2( u2_u1_u2_n165 ) );
  AND2_X1 u2_u1_u2_U78 (.A2( u2_u1_X_15 ) , .A1( u2_u1_X_18 ) , .ZN( u2_u1_u2_n107 ) );
  AND2_X1 u2_u1_u2_U79 (.A1( u2_u1_X_14 ) , .ZN( u2_u1_u2_n106 ) , .A2( u2_u1_u2_n174 ) );
  AOI21_X1 u2_u1_u2_U8 (.ZN( u2_u1_u2_n124 ) , .B1( u2_u1_u2_n131 ) , .B2( u2_u1_u2_n143 ) , .A( u2_u1_u2_n172 ) );
  AND2_X1 u2_u1_u2_U80 (.A1( u2_u1_X_13 ) , .A2( u2_u1_X_14 ) , .ZN( u2_u1_u2_n108 ) );
  INV_X1 u2_u1_u2_U81 (.A( u2_u1_X_16 ) , .ZN( u2_u1_u2_n169 ) );
  INV_X1 u2_u1_u2_U82 (.A( u2_u1_X_17 ) , .ZN( u2_u1_u2_n166 ) );
  INV_X1 u2_u1_u2_U83 (.A( u2_u1_X_13 ) , .ZN( u2_u1_u2_n174 ) );
  INV_X1 u2_u1_u2_U84 (.A( u2_u1_X_18 ) , .ZN( u2_u1_u2_n165 ) );
  NAND4_X1 u2_u1_u2_U85 (.ZN( u2_out1_30 ) , .A4( u2_u1_u2_n147 ) , .A3( u2_u1_u2_n148 ) , .A2( u2_u1_u2_n149 ) , .A1( u2_u1_u2_n187 ) );
  NOR3_X1 u2_u1_u2_U86 (.A3( u2_u1_u2_n144 ) , .A2( u2_u1_u2_n145 ) , .A1( u2_u1_u2_n146 ) , .ZN( u2_u1_u2_n147 ) );
  AOI21_X1 u2_u1_u2_U87 (.B2( u2_u1_u2_n138 ) , .ZN( u2_u1_u2_n148 ) , .A( u2_u1_u2_n162 ) , .B1( u2_u1_u2_n182 ) );
  NAND4_X1 u2_u1_u2_U88 (.ZN( u2_out1_24 ) , .A4( u2_u1_u2_n111 ) , .A3( u2_u1_u2_n112 ) , .A1( u2_u1_u2_n130 ) , .A2( u2_u1_u2_n187 ) );
  AOI221_X1 u2_u1_u2_U89 (.A( u2_u1_u2_n109 ) , .B1( u2_u1_u2_n110 ) , .ZN( u2_u1_u2_n111 ) , .C1( u2_u1_u2_n134 ) , .C2( u2_u1_u2_n170 ) , .B2( u2_u1_u2_n173 ) );
  AOI21_X1 u2_u1_u2_U9 (.B2( u2_u1_u2_n123 ) , .ZN( u2_u1_u2_n125 ) , .A( u2_u1_u2_n171 ) , .B1( u2_u1_u2_n184 ) );
  AOI21_X1 u2_u1_u2_U90 (.ZN( u2_u1_u2_n112 ) , .B2( u2_u1_u2_n156 ) , .A( u2_u1_u2_n164 ) , .B1( u2_u1_u2_n181 ) );
  NAND4_X1 u2_u1_u2_U91 (.ZN( u2_out1_16 ) , .A4( u2_u1_u2_n128 ) , .A3( u2_u1_u2_n129 ) , .A1( u2_u1_u2_n130 ) , .A2( u2_u1_u2_n186 ) );
  AOI22_X1 u2_u1_u2_U92 (.A2( u2_u1_u2_n118 ) , .ZN( u2_u1_u2_n129 ) , .A1( u2_u1_u2_n140 ) , .B1( u2_u1_u2_n157 ) , .B2( u2_u1_u2_n170 ) );
  INV_X1 u2_u1_u2_U93 (.A( u2_u1_u2_n163 ) , .ZN( u2_u1_u2_n186 ) );
  OR4_X1 u2_u1_u2_U94 (.ZN( u2_out1_6 ) , .A4( u2_u1_u2_n161 ) , .A3( u2_u1_u2_n162 ) , .A2( u2_u1_u2_n163 ) , .A1( u2_u1_u2_n164 ) );
  OR3_X1 u2_u1_u2_U95 (.A2( u2_u1_u2_n159 ) , .A1( u2_u1_u2_n160 ) , .ZN( u2_u1_u2_n161 ) , .A3( u2_u1_u2_n183 ) );
  AOI21_X1 u2_u1_u2_U96 (.B2( u2_u1_u2_n154 ) , .B1( u2_u1_u2_n155 ) , .ZN( u2_u1_u2_n159 ) , .A( u2_u1_u2_n167 ) );
  NAND3_X1 u2_u1_u2_U97 (.A2( u2_u1_u2_n117 ) , .A1( u2_u1_u2_n122 ) , .A3( u2_u1_u2_n123 ) , .ZN( u2_u1_u2_n134 ) );
  NAND3_X1 u2_u1_u2_U98 (.ZN( u2_u1_u2_n110 ) , .A2( u2_u1_u2_n131 ) , .A3( u2_u1_u2_n139 ) , .A1( u2_u1_u2_n154 ) );
  NAND3_X1 u2_u1_u2_U99 (.A2( u2_u1_u2_n100 ) , .ZN( u2_u1_u2_n101 ) , .A1( u2_u1_u2_n104 ) , .A3( u2_u1_u2_n114 ) );
  OAI22_X1 u2_u1_u3_U10 (.B1( u2_u1_u3_n113 ) , .A2( u2_u1_u3_n135 ) , .A1( u2_u1_u3_n150 ) , .B2( u2_u1_u3_n164 ) , .ZN( u2_u1_u3_n98 ) );
  OAI211_X1 u2_u1_u3_U11 (.B( u2_u1_u3_n106 ) , .ZN( u2_u1_u3_n119 ) , .C2( u2_u1_u3_n128 ) , .C1( u2_u1_u3_n167 ) , .A( u2_u1_u3_n181 ) );
  AOI221_X1 u2_u1_u3_U12 (.C1( u2_u1_u3_n105 ) , .ZN( u2_u1_u3_n106 ) , .A( u2_u1_u3_n131 ) , .B2( u2_u1_u3_n132 ) , .C2( u2_u1_u3_n133 ) , .B1( u2_u1_u3_n169 ) );
  INV_X1 u2_u1_u3_U13 (.ZN( u2_u1_u3_n181 ) , .A( u2_u1_u3_n98 ) );
  NAND2_X1 u2_u1_u3_U14 (.ZN( u2_u1_u3_n105 ) , .A2( u2_u1_u3_n130 ) , .A1( u2_u1_u3_n155 ) );
  AOI22_X1 u2_u1_u3_U15 (.B1( u2_u1_u3_n115 ) , .A2( u2_u1_u3_n116 ) , .ZN( u2_u1_u3_n123 ) , .B2( u2_u1_u3_n133 ) , .A1( u2_u1_u3_n169 ) );
  NAND2_X1 u2_u1_u3_U16 (.ZN( u2_u1_u3_n116 ) , .A2( u2_u1_u3_n151 ) , .A1( u2_u1_u3_n182 ) );
  NOR2_X1 u2_u1_u3_U17 (.ZN( u2_u1_u3_n126 ) , .A2( u2_u1_u3_n150 ) , .A1( u2_u1_u3_n164 ) );
  AOI21_X1 u2_u1_u3_U18 (.ZN( u2_u1_u3_n112 ) , .B2( u2_u1_u3_n146 ) , .B1( u2_u1_u3_n155 ) , .A( u2_u1_u3_n167 ) );
  NAND2_X1 u2_u1_u3_U19 (.A1( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n142 ) , .A2( u2_u1_u3_n164 ) );
  NAND2_X1 u2_u1_u3_U20 (.ZN( u2_u1_u3_n132 ) , .A2( u2_u1_u3_n152 ) , .A1( u2_u1_u3_n156 ) );
  AND2_X1 u2_u1_u3_U21 (.A2( u2_u1_u3_n113 ) , .A1( u2_u1_u3_n114 ) , .ZN( u2_u1_u3_n151 ) );
  INV_X1 u2_u1_u3_U22 (.A( u2_u1_u3_n133 ) , .ZN( u2_u1_u3_n165 ) );
  INV_X1 u2_u1_u3_U23 (.A( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n170 ) );
  NAND2_X1 u2_u1_u3_U24 (.A1( u2_u1_u3_n107 ) , .A2( u2_u1_u3_n108 ) , .ZN( u2_u1_u3_n140 ) );
  NAND2_X1 u2_u1_u3_U25 (.ZN( u2_u1_u3_n117 ) , .A1( u2_u1_u3_n124 ) , .A2( u2_u1_u3_n148 ) );
  NAND2_X1 u2_u1_u3_U26 (.ZN( u2_u1_u3_n143 ) , .A1( u2_u1_u3_n165 ) , .A2( u2_u1_u3_n167 ) );
  INV_X1 u2_u1_u3_U27 (.A( u2_u1_u3_n130 ) , .ZN( u2_u1_u3_n177 ) );
  INV_X1 u2_u1_u3_U28 (.A( u2_u1_u3_n128 ) , .ZN( u2_u1_u3_n176 ) );
  INV_X1 u2_u1_u3_U29 (.A( u2_u1_u3_n155 ) , .ZN( u2_u1_u3_n174 ) );
  INV_X1 u2_u1_u3_U3 (.A( u2_u1_u3_n129 ) , .ZN( u2_u1_u3_n183 ) );
  INV_X1 u2_u1_u3_U30 (.A( u2_u1_u3_n139 ) , .ZN( u2_u1_u3_n185 ) );
  NOR2_X1 u2_u1_u3_U31 (.ZN( u2_u1_u3_n135 ) , .A2( u2_u1_u3_n141 ) , .A1( u2_u1_u3_n169 ) );
  OAI222_X1 u2_u1_u3_U32 (.C2( u2_u1_u3_n107 ) , .A2( u2_u1_u3_n108 ) , .B1( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n138 ) , .B2( u2_u1_u3_n146 ) , .C1( u2_u1_u3_n154 ) , .A1( u2_u1_u3_n164 ) );
  NOR4_X1 u2_u1_u3_U33 (.A4( u2_u1_u3_n157 ) , .A3( u2_u1_u3_n158 ) , .A2( u2_u1_u3_n159 ) , .A1( u2_u1_u3_n160 ) , .ZN( u2_u1_u3_n161 ) );
  AOI21_X1 u2_u1_u3_U34 (.B2( u2_u1_u3_n152 ) , .B1( u2_u1_u3_n153 ) , .ZN( u2_u1_u3_n158 ) , .A( u2_u1_u3_n164 ) );
  AOI21_X1 u2_u1_u3_U35 (.A( u2_u1_u3_n154 ) , .B2( u2_u1_u3_n155 ) , .B1( u2_u1_u3_n156 ) , .ZN( u2_u1_u3_n157 ) );
  AOI21_X1 u2_u1_u3_U36 (.A( u2_u1_u3_n149 ) , .B2( u2_u1_u3_n150 ) , .B1( u2_u1_u3_n151 ) , .ZN( u2_u1_u3_n159 ) );
  AOI211_X1 u2_u1_u3_U37 (.ZN( u2_u1_u3_n109 ) , .A( u2_u1_u3_n119 ) , .C2( u2_u1_u3_n129 ) , .B( u2_u1_u3_n138 ) , .C1( u2_u1_u3_n141 ) );
  AOI211_X1 u2_u1_u3_U38 (.B( u2_u1_u3_n119 ) , .A( u2_u1_u3_n120 ) , .C2( u2_u1_u3_n121 ) , .ZN( u2_u1_u3_n122 ) , .C1( u2_u1_u3_n179 ) );
  INV_X1 u2_u1_u3_U39 (.A( u2_u1_u3_n156 ) , .ZN( u2_u1_u3_n179 ) );
  INV_X1 u2_u1_u3_U4 (.A( u2_u1_u3_n140 ) , .ZN( u2_u1_u3_n182 ) );
  OAI22_X1 u2_u1_u3_U40 (.B1( u2_u1_u3_n118 ) , .ZN( u2_u1_u3_n120 ) , .A1( u2_u1_u3_n135 ) , .B2( u2_u1_u3_n154 ) , .A2( u2_u1_u3_n178 ) );
  AND3_X1 u2_u1_u3_U41 (.ZN( u2_u1_u3_n118 ) , .A2( u2_u1_u3_n124 ) , .A1( u2_u1_u3_n144 ) , .A3( u2_u1_u3_n152 ) );
  INV_X1 u2_u1_u3_U42 (.A( u2_u1_u3_n121 ) , .ZN( u2_u1_u3_n164 ) );
  NAND2_X1 u2_u1_u3_U43 (.ZN( u2_u1_u3_n133 ) , .A1( u2_u1_u3_n154 ) , .A2( u2_u1_u3_n164 ) );
  OAI211_X1 u2_u1_u3_U44 (.B( u2_u1_u3_n127 ) , .ZN( u2_u1_u3_n139 ) , .C1( u2_u1_u3_n150 ) , .C2( u2_u1_u3_n154 ) , .A( u2_u1_u3_n184 ) );
  INV_X1 u2_u1_u3_U45 (.A( u2_u1_u3_n125 ) , .ZN( u2_u1_u3_n184 ) );
  AOI221_X1 u2_u1_u3_U46 (.A( u2_u1_u3_n126 ) , .ZN( u2_u1_u3_n127 ) , .C2( u2_u1_u3_n132 ) , .C1( u2_u1_u3_n169 ) , .B2( u2_u1_u3_n170 ) , .B1( u2_u1_u3_n174 ) );
  OAI22_X1 u2_u1_u3_U47 (.A1( u2_u1_u3_n124 ) , .ZN( u2_u1_u3_n125 ) , .B2( u2_u1_u3_n145 ) , .A2( u2_u1_u3_n165 ) , .B1( u2_u1_u3_n167 ) );
  NOR2_X1 u2_u1_u3_U48 (.A1( u2_u1_u3_n113 ) , .ZN( u2_u1_u3_n131 ) , .A2( u2_u1_u3_n154 ) );
  NAND2_X1 u2_u1_u3_U49 (.A1( u2_u1_u3_n103 ) , .ZN( u2_u1_u3_n150 ) , .A2( u2_u1_u3_n99 ) );
  INV_X1 u2_u1_u3_U5 (.A( u2_u1_u3_n117 ) , .ZN( u2_u1_u3_n178 ) );
  NAND2_X1 u2_u1_u3_U50 (.A2( u2_u1_u3_n102 ) , .ZN( u2_u1_u3_n155 ) , .A1( u2_u1_u3_n97 ) );
  INV_X1 u2_u1_u3_U51 (.A( u2_u1_u3_n141 ) , .ZN( u2_u1_u3_n167 ) );
  AOI21_X1 u2_u1_u3_U52 (.B2( u2_u1_u3_n114 ) , .B1( u2_u1_u3_n146 ) , .A( u2_u1_u3_n154 ) , .ZN( u2_u1_u3_n94 ) );
  AOI21_X1 u2_u1_u3_U53 (.ZN( u2_u1_u3_n110 ) , .B2( u2_u1_u3_n142 ) , .B1( u2_u1_u3_n186 ) , .A( u2_u1_u3_n95 ) );
  INV_X1 u2_u1_u3_U54 (.A( u2_u1_u3_n145 ) , .ZN( u2_u1_u3_n186 ) );
  AOI21_X1 u2_u1_u3_U55 (.B1( u2_u1_u3_n124 ) , .A( u2_u1_u3_n149 ) , .B2( u2_u1_u3_n155 ) , .ZN( u2_u1_u3_n95 ) );
  INV_X1 u2_u1_u3_U56 (.A( u2_u1_u3_n149 ) , .ZN( u2_u1_u3_n169 ) );
  NAND2_X1 u2_u1_u3_U57 (.ZN( u2_u1_u3_n124 ) , .A1( u2_u1_u3_n96 ) , .A2( u2_u1_u3_n97 ) );
  NAND2_X1 u2_u1_u3_U58 (.A2( u2_u1_u3_n100 ) , .ZN( u2_u1_u3_n146 ) , .A1( u2_u1_u3_n96 ) );
  NAND2_X1 u2_u1_u3_U59 (.A1( u2_u1_u3_n101 ) , .ZN( u2_u1_u3_n145 ) , .A2( u2_u1_u3_n99 ) );
  AOI221_X1 u2_u1_u3_U6 (.A( u2_u1_u3_n131 ) , .C2( u2_u1_u3_n132 ) , .C1( u2_u1_u3_n133 ) , .ZN( u2_u1_u3_n134 ) , .B1( u2_u1_u3_n143 ) , .B2( u2_u1_u3_n177 ) );
  NAND2_X1 u2_u1_u3_U60 (.A1( u2_u1_u3_n100 ) , .ZN( u2_u1_u3_n156 ) , .A2( u2_u1_u3_n99 ) );
  NAND2_X1 u2_u1_u3_U61 (.A2( u2_u1_u3_n101 ) , .A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n148 ) );
  NAND2_X1 u2_u1_u3_U62 (.A1( u2_u1_u3_n100 ) , .A2( u2_u1_u3_n102 ) , .ZN( u2_u1_u3_n128 ) );
  NAND2_X1 u2_u1_u3_U63 (.A2( u2_u1_u3_n101 ) , .A1( u2_u1_u3_n102 ) , .ZN( u2_u1_u3_n152 ) );
  NAND2_X1 u2_u1_u3_U64 (.A2( u2_u1_u3_n101 ) , .ZN( u2_u1_u3_n114 ) , .A1( u2_u1_u3_n96 ) );
  NAND2_X1 u2_u1_u3_U65 (.ZN( u2_u1_u3_n107 ) , .A1( u2_u1_u3_n97 ) , .A2( u2_u1_u3_n99 ) );
  NAND2_X1 u2_u1_u3_U66 (.A2( u2_u1_u3_n100 ) , .A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n113 ) );
  NAND2_X1 u2_u1_u3_U67 (.A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n153 ) , .A2( u2_u1_u3_n97 ) );
  NAND2_X1 u2_u1_u3_U68 (.A2( u2_u1_u3_n103 ) , .A1( u2_u1_u3_n104 ) , .ZN( u2_u1_u3_n130 ) );
  NAND2_X1 u2_u1_u3_U69 (.A2( u2_u1_u3_n103 ) , .ZN( u2_u1_u3_n144 ) , .A1( u2_u1_u3_n96 ) );
  OAI22_X1 u2_u1_u3_U7 (.B2( u2_u1_u3_n147 ) , .A2( u2_u1_u3_n148 ) , .ZN( u2_u1_u3_n160 ) , .B1( u2_u1_u3_n165 ) , .A1( u2_u1_u3_n168 ) );
  NAND2_X1 u2_u1_u3_U70 (.A1( u2_u1_u3_n102 ) , .A2( u2_u1_u3_n103 ) , .ZN( u2_u1_u3_n108 ) );
  NOR2_X1 u2_u1_u3_U71 (.A2( u2_u1_X_19 ) , .A1( u2_u1_X_20 ) , .ZN( u2_u1_u3_n99 ) );
  NOR2_X1 u2_u1_u3_U72 (.A2( u2_u1_X_21 ) , .A1( u2_u1_X_24 ) , .ZN( u2_u1_u3_n103 ) );
  NOR2_X1 u2_u1_u3_U73 (.A2( u2_u1_X_24 ) , .A1( u2_u1_u3_n171 ) , .ZN( u2_u1_u3_n97 ) );
  NOR2_X1 u2_u1_u3_U74 (.A2( u2_u1_X_23 ) , .ZN( u2_u1_u3_n141 ) , .A1( u2_u1_u3_n166 ) );
  NOR2_X1 u2_u1_u3_U75 (.A2( u2_u1_X_19 ) , .A1( u2_u1_u3_n172 ) , .ZN( u2_u1_u3_n96 ) );
  NAND2_X1 u2_u1_u3_U76 (.A1( u2_u1_X_22 ) , .A2( u2_u1_X_23 ) , .ZN( u2_u1_u3_n154 ) );
  NAND2_X1 u2_u1_u3_U77 (.A1( u2_u1_X_23 ) , .ZN( u2_u1_u3_n149 ) , .A2( u2_u1_u3_n166 ) );
  NOR2_X1 u2_u1_u3_U78 (.A2( u2_u1_X_22 ) , .A1( u2_u1_X_23 ) , .ZN( u2_u1_u3_n121 ) );
  AND2_X1 u2_u1_u3_U79 (.A1( u2_u1_X_24 ) , .ZN( u2_u1_u3_n101 ) , .A2( u2_u1_u3_n171 ) );
  AND3_X1 u2_u1_u3_U8 (.A3( u2_u1_u3_n144 ) , .A2( u2_u1_u3_n145 ) , .A1( u2_u1_u3_n146 ) , .ZN( u2_u1_u3_n147 ) );
  AND2_X1 u2_u1_u3_U80 (.A1( u2_u1_X_19 ) , .ZN( u2_u1_u3_n102 ) , .A2( u2_u1_u3_n172 ) );
  AND2_X1 u2_u1_u3_U81 (.A1( u2_u1_X_21 ) , .A2( u2_u1_X_24 ) , .ZN( u2_u1_u3_n100 ) );
  AND2_X1 u2_u1_u3_U82 (.A2( u2_u1_X_19 ) , .A1( u2_u1_X_20 ) , .ZN( u2_u1_u3_n104 ) );
  INV_X1 u2_u1_u3_U83 (.A( u2_u1_X_22 ) , .ZN( u2_u1_u3_n166 ) );
  INV_X1 u2_u1_u3_U84 (.A( u2_u1_X_21 ) , .ZN( u2_u1_u3_n171 ) );
  INV_X1 u2_u1_u3_U85 (.A( u2_u1_X_20 ) , .ZN( u2_u1_u3_n172 ) );
  OR4_X1 u2_u1_u3_U86 (.ZN( u2_out1_10 ) , .A4( u2_u1_u3_n136 ) , .A3( u2_u1_u3_n137 ) , .A1( u2_u1_u3_n138 ) , .A2( u2_u1_u3_n139 ) );
  OAI222_X1 u2_u1_u3_U87 (.C1( u2_u1_u3_n128 ) , .ZN( u2_u1_u3_n137 ) , .B1( u2_u1_u3_n148 ) , .A2( u2_u1_u3_n150 ) , .B2( u2_u1_u3_n154 ) , .C2( u2_u1_u3_n164 ) , .A1( u2_u1_u3_n167 ) );
  OAI221_X1 u2_u1_u3_U88 (.A( u2_u1_u3_n134 ) , .B2( u2_u1_u3_n135 ) , .ZN( u2_u1_u3_n136 ) , .C1( u2_u1_u3_n149 ) , .B1( u2_u1_u3_n151 ) , .C2( u2_u1_u3_n183 ) );
  NAND4_X1 u2_u1_u3_U89 (.ZN( u2_out1_26 ) , .A4( u2_u1_u3_n109 ) , .A3( u2_u1_u3_n110 ) , .A2( u2_u1_u3_n111 ) , .A1( u2_u1_u3_n173 ) );
  INV_X1 u2_u1_u3_U9 (.A( u2_u1_u3_n143 ) , .ZN( u2_u1_u3_n168 ) );
  INV_X1 u2_u1_u3_U90 (.ZN( u2_u1_u3_n173 ) , .A( u2_u1_u3_n94 ) );
  OAI21_X1 u2_u1_u3_U91 (.ZN( u2_u1_u3_n111 ) , .B2( u2_u1_u3_n117 ) , .A( u2_u1_u3_n133 ) , .B1( u2_u1_u3_n176 ) );
  NAND4_X1 u2_u1_u3_U92 (.ZN( u2_out1_20 ) , .A4( u2_u1_u3_n122 ) , .A3( u2_u1_u3_n123 ) , .A1( u2_u1_u3_n175 ) , .A2( u2_u1_u3_n180 ) );
  INV_X1 u2_u1_u3_U93 (.A( u2_u1_u3_n112 ) , .ZN( u2_u1_u3_n175 ) );
  INV_X1 u2_u1_u3_U94 (.A( u2_u1_u3_n126 ) , .ZN( u2_u1_u3_n180 ) );
  NAND4_X1 u2_u1_u3_U95 (.ZN( u2_out1_1 ) , .A4( u2_u1_u3_n161 ) , .A3( u2_u1_u3_n162 ) , .A2( u2_u1_u3_n163 ) , .A1( u2_u1_u3_n185 ) );
  NAND2_X1 u2_u1_u3_U96 (.ZN( u2_u1_u3_n163 ) , .A2( u2_u1_u3_n170 ) , .A1( u2_u1_u3_n176 ) );
  AOI22_X1 u2_u1_u3_U97 (.B2( u2_u1_u3_n140 ) , .B1( u2_u1_u3_n141 ) , .A2( u2_u1_u3_n142 ) , .ZN( u2_u1_u3_n162 ) , .A1( u2_u1_u3_n177 ) );
  NAND3_X1 u2_u1_u3_U98 (.A1( u2_u1_u3_n114 ) , .ZN( u2_u1_u3_n115 ) , .A2( u2_u1_u3_n145 ) , .A3( u2_u1_u3_n153 ) );
  NAND3_X1 u2_u1_u3_U99 (.ZN( u2_u1_u3_n129 ) , .A2( u2_u1_u3_n144 ) , .A1( u2_u1_u3_n153 ) , .A3( u2_u1_u3_n182 ) );
  XOR2_X1 u2_u2_U26 (.B( u2_K3_30 ) , .A( u2_R1_21 ) , .Z( u2_u2_X_30 ) );
  XOR2_X1 u2_u2_U28 (.B( u2_K3_29 ) , .A( u2_R1_20 ) , .Z( u2_u2_X_29 ) );
  XOR2_X1 u2_u2_U29 (.B( u2_K3_28 ) , .A( u2_R1_19 ) , .Z( u2_u2_X_28 ) );
  XOR2_X1 u2_u2_U30 (.B( u2_K3_27 ) , .A( u2_R1_18 ) , .Z( u2_u2_X_27 ) );
  XOR2_X1 u2_u2_U31 (.B( u2_K3_26 ) , .A( u2_R1_17 ) , .Z( u2_u2_X_26 ) );
  XOR2_X1 u2_u2_U32 (.B( u2_K3_25 ) , .A( u2_R1_16 ) , .Z( u2_u2_X_25 ) );
  OAI22_X1 u2_u2_u4_U10 (.B2( u2_u2_u4_n135 ) , .ZN( u2_u2_u4_n137 ) , .B1( u2_u2_u4_n153 ) , .A1( u2_u2_u4_n155 ) , .A2( u2_u2_u4_n171 ) );
  AND3_X1 u2_u2_u4_U11 (.A2( u2_u2_u4_n134 ) , .ZN( u2_u2_u4_n135 ) , .A3( u2_u2_u4_n145 ) , .A1( u2_u2_u4_n157 ) );
  NAND2_X1 u2_u2_u4_U12 (.ZN( u2_u2_u4_n132 ) , .A2( u2_u2_u4_n170 ) , .A1( u2_u2_u4_n173 ) );
  AOI21_X1 u2_u2_u4_U13 (.B2( u2_u2_u4_n160 ) , .B1( u2_u2_u4_n161 ) , .ZN( u2_u2_u4_n162 ) , .A( u2_u2_u4_n170 ) );
  AOI21_X1 u2_u2_u4_U14 (.ZN( u2_u2_u4_n107 ) , .B2( u2_u2_u4_n143 ) , .A( u2_u2_u4_n174 ) , .B1( u2_u2_u4_n184 ) );
  AOI21_X1 u2_u2_u4_U15 (.B2( u2_u2_u4_n158 ) , .B1( u2_u2_u4_n159 ) , .ZN( u2_u2_u4_n163 ) , .A( u2_u2_u4_n174 ) );
  AOI21_X1 u2_u2_u4_U16 (.A( u2_u2_u4_n153 ) , .B2( u2_u2_u4_n154 ) , .B1( u2_u2_u4_n155 ) , .ZN( u2_u2_u4_n165 ) );
  AOI21_X1 u2_u2_u4_U17 (.A( u2_u2_u4_n156 ) , .B2( u2_u2_u4_n157 ) , .ZN( u2_u2_u4_n164 ) , .B1( u2_u2_u4_n184 ) );
  INV_X1 u2_u2_u4_U18 (.A( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n170 ) );
  AND2_X1 u2_u2_u4_U19 (.A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n155 ) , .A1( u2_u2_u4_n160 ) );
  INV_X1 u2_u2_u4_U20 (.A( u2_u2_u4_n156 ) , .ZN( u2_u2_u4_n175 ) );
  NAND2_X1 u2_u2_u4_U21 (.A2( u2_u2_u4_n118 ) , .ZN( u2_u2_u4_n131 ) , .A1( u2_u2_u4_n147 ) );
  NAND2_X1 u2_u2_u4_U22 (.A1( u2_u2_u4_n119 ) , .A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n130 ) );
  NAND2_X1 u2_u2_u4_U23 (.ZN( u2_u2_u4_n117 ) , .A2( u2_u2_u4_n118 ) , .A1( u2_u2_u4_n148 ) );
  NAND2_X1 u2_u2_u4_U24 (.ZN( u2_u2_u4_n129 ) , .A1( u2_u2_u4_n134 ) , .A2( u2_u2_u4_n148 ) );
  AND3_X1 u2_u2_u4_U25 (.A1( u2_u2_u4_n119 ) , .A2( u2_u2_u4_n143 ) , .A3( u2_u2_u4_n154 ) , .ZN( u2_u2_u4_n161 ) );
  AND2_X1 u2_u2_u4_U26 (.A1( u2_u2_u4_n145 ) , .A2( u2_u2_u4_n147 ) , .ZN( u2_u2_u4_n159 ) );
  OR3_X1 u2_u2_u4_U27 (.A3( u2_u2_u4_n114 ) , .A2( u2_u2_u4_n115 ) , .A1( u2_u2_u4_n116 ) , .ZN( u2_u2_u4_n136 ) );
  AOI21_X1 u2_u2_u4_U28 (.A( u2_u2_u4_n113 ) , .ZN( u2_u2_u4_n116 ) , .B2( u2_u2_u4_n173 ) , .B1( u2_u2_u4_n174 ) );
  AOI21_X1 u2_u2_u4_U29 (.ZN( u2_u2_u4_n115 ) , .B2( u2_u2_u4_n145 ) , .B1( u2_u2_u4_n146 ) , .A( u2_u2_u4_n156 ) );
  NOR2_X1 u2_u2_u4_U3 (.ZN( u2_u2_u4_n121 ) , .A1( u2_u2_u4_n181 ) , .A2( u2_u2_u4_n182 ) );
  OAI22_X1 u2_u2_u4_U30 (.ZN( u2_u2_u4_n114 ) , .A2( u2_u2_u4_n121 ) , .B1( u2_u2_u4_n160 ) , .B2( u2_u2_u4_n170 ) , .A1( u2_u2_u4_n171 ) );
  INV_X1 u2_u2_u4_U31 (.A( u2_u2_u4_n158 ) , .ZN( u2_u2_u4_n182 ) );
  INV_X1 u2_u2_u4_U32 (.ZN( u2_u2_u4_n181 ) , .A( u2_u2_u4_n96 ) );
  INV_X1 u2_u2_u4_U33 (.A( u2_u2_u4_n144 ) , .ZN( u2_u2_u4_n179 ) );
  INV_X1 u2_u2_u4_U34 (.A( u2_u2_u4_n157 ) , .ZN( u2_u2_u4_n178 ) );
  NAND2_X1 u2_u2_u4_U35 (.A2( u2_u2_u4_n154 ) , .A1( u2_u2_u4_n96 ) , .ZN( u2_u2_u4_n97 ) );
  INV_X1 u2_u2_u4_U36 (.ZN( u2_u2_u4_n186 ) , .A( u2_u2_u4_n95 ) );
  OAI221_X1 u2_u2_u4_U37 (.C1( u2_u2_u4_n134 ) , .B1( u2_u2_u4_n158 ) , .B2( u2_u2_u4_n171 ) , .C2( u2_u2_u4_n173 ) , .A( u2_u2_u4_n94 ) , .ZN( u2_u2_u4_n95 ) );
  AOI222_X1 u2_u2_u4_U38 (.B2( u2_u2_u4_n132 ) , .A1( u2_u2_u4_n138 ) , .C2( u2_u2_u4_n175 ) , .A2( u2_u2_u4_n179 ) , .C1( u2_u2_u4_n181 ) , .B1( u2_u2_u4_n185 ) , .ZN( u2_u2_u4_n94 ) );
  INV_X1 u2_u2_u4_U39 (.A( u2_u2_u4_n113 ) , .ZN( u2_u2_u4_n185 ) );
  INV_X1 u2_u2_u4_U4 (.A( u2_u2_u4_n117 ) , .ZN( u2_u2_u4_n184 ) );
  INV_X1 u2_u2_u4_U40 (.A( u2_u2_u4_n143 ) , .ZN( u2_u2_u4_n183 ) );
  NOR2_X1 u2_u2_u4_U41 (.ZN( u2_u2_u4_n138 ) , .A1( u2_u2_u4_n168 ) , .A2( u2_u2_u4_n169 ) );
  NOR2_X1 u2_u2_u4_U42 (.A1( u2_u2_u4_n150 ) , .A2( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n153 ) );
  NOR2_X1 u2_u2_u4_U43 (.A2( u2_u2_u4_n128 ) , .A1( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n156 ) );
  AOI22_X1 u2_u2_u4_U44 (.B2( u2_u2_u4_n122 ) , .A1( u2_u2_u4_n123 ) , .ZN( u2_u2_u4_n124 ) , .B1( u2_u2_u4_n128 ) , .A2( u2_u2_u4_n172 ) );
  INV_X1 u2_u2_u4_U45 (.A( u2_u2_u4_n153 ) , .ZN( u2_u2_u4_n172 ) );
  NAND2_X1 u2_u2_u4_U46 (.A2( u2_u2_u4_n120 ) , .ZN( u2_u2_u4_n123 ) , .A1( u2_u2_u4_n161 ) );
  AOI22_X1 u2_u2_u4_U47 (.B2( u2_u2_u4_n132 ) , .A2( u2_u2_u4_n133 ) , .ZN( u2_u2_u4_n140 ) , .A1( u2_u2_u4_n150 ) , .B1( u2_u2_u4_n179 ) );
  NAND2_X1 u2_u2_u4_U48 (.ZN( u2_u2_u4_n133 ) , .A2( u2_u2_u4_n146 ) , .A1( u2_u2_u4_n154 ) );
  NAND2_X1 u2_u2_u4_U49 (.A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n154 ) , .A2( u2_u2_u4_n98 ) );
  NOR4_X1 u2_u2_u4_U5 (.A4( u2_u2_u4_n106 ) , .A3( u2_u2_u4_n107 ) , .A2( u2_u2_u4_n108 ) , .A1( u2_u2_u4_n109 ) , .ZN( u2_u2_u4_n110 ) );
  NAND2_X1 u2_u2_u4_U50 (.A1( u2_u2_u4_n101 ) , .ZN( u2_u2_u4_n158 ) , .A2( u2_u2_u4_n99 ) );
  AOI21_X1 u2_u2_u4_U51 (.ZN( u2_u2_u4_n127 ) , .A( u2_u2_u4_n136 ) , .B2( u2_u2_u4_n150 ) , .B1( u2_u2_u4_n180 ) );
  INV_X1 u2_u2_u4_U52 (.A( u2_u2_u4_n160 ) , .ZN( u2_u2_u4_n180 ) );
  NAND2_X1 u2_u2_u4_U53 (.A2( u2_u2_u4_n104 ) , .A1( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n146 ) );
  NAND2_X1 u2_u2_u4_U54 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n160 ) );
  NAND2_X1 u2_u2_u4_U55 (.ZN( u2_u2_u4_n134 ) , .A1( u2_u2_u4_n98 ) , .A2( u2_u2_u4_n99 ) );
  NAND2_X1 u2_u2_u4_U56 (.A1( u2_u2_u4_n103 ) , .A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n143 ) );
  NAND2_X1 u2_u2_u4_U57 (.A2( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n145 ) , .A1( u2_u2_u4_n98 ) );
  NAND2_X1 u2_u2_u4_U58 (.A1( u2_u2_u4_n100 ) , .A2( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n120 ) );
  NAND2_X1 u2_u2_u4_U59 (.A1( u2_u2_u4_n102 ) , .A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n148 ) );
  AOI21_X1 u2_u2_u4_U6 (.ZN( u2_u2_u4_n106 ) , .B2( u2_u2_u4_n146 ) , .B1( u2_u2_u4_n158 ) , .A( u2_u2_u4_n170 ) );
  NAND2_X1 u2_u2_u4_U60 (.A2( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n157 ) );
  INV_X1 u2_u2_u4_U61 (.A( u2_u2_u4_n150 ) , .ZN( u2_u2_u4_n173 ) );
  INV_X1 u2_u2_u4_U62 (.A( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n171 ) );
  NAND2_X1 u2_u2_u4_U63 (.A1( u2_u2_u4_n100 ) , .ZN( u2_u2_u4_n118 ) , .A2( u2_u2_u4_n99 ) );
  NAND2_X1 u2_u2_u4_U64 (.A2( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n144 ) );
  NAND2_X1 u2_u2_u4_U65 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n105 ) , .ZN( u2_u2_u4_n96 ) );
  INV_X1 u2_u2_u4_U66 (.A( u2_u2_u4_n128 ) , .ZN( u2_u2_u4_n174 ) );
  NAND2_X1 u2_u2_u4_U67 (.A2( u2_u2_u4_n102 ) , .ZN( u2_u2_u4_n119 ) , .A1( u2_u2_u4_n98 ) );
  NAND2_X1 u2_u2_u4_U68 (.A2( u2_u2_u4_n101 ) , .A1( u2_u2_u4_n103 ) , .ZN( u2_u2_u4_n147 ) );
  NAND2_X1 u2_u2_u4_U69 (.A2( u2_u2_u4_n104 ) , .ZN( u2_u2_u4_n113 ) , .A1( u2_u2_u4_n99 ) );
  AOI21_X1 u2_u2_u4_U7 (.ZN( u2_u2_u4_n108 ) , .B2( u2_u2_u4_n134 ) , .B1( u2_u2_u4_n155 ) , .A( u2_u2_u4_n156 ) );
  NOR2_X1 u2_u2_u4_U70 (.A2( u2_u2_X_28 ) , .ZN( u2_u2_u4_n150 ) , .A1( u2_u2_u4_n168 ) );
  NOR2_X1 u2_u2_u4_U71 (.A2( u2_u2_X_29 ) , .ZN( u2_u2_u4_n152 ) , .A1( u2_u2_u4_n169 ) );
  NOR2_X1 u2_u2_u4_U72 (.A2( u2_u2_X_30 ) , .ZN( u2_u2_u4_n105 ) , .A1( u2_u2_u4_n176 ) );
  NOR2_X1 u2_u2_u4_U73 (.A2( u2_u2_X_26 ) , .ZN( u2_u2_u4_n100 ) , .A1( u2_u2_u4_n177 ) );
  NOR2_X1 u2_u2_u4_U74 (.A2( u2_u2_X_28 ) , .A1( u2_u2_X_29 ) , .ZN( u2_u2_u4_n128 ) );
  NOR2_X1 u2_u2_u4_U75 (.A2( u2_u2_X_27 ) , .A1( u2_u2_X_30 ) , .ZN( u2_u2_u4_n102 ) );
  NOR2_X1 u2_u2_u4_U76 (.A2( u2_u2_X_25 ) , .A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n98 ) );
  AND2_X1 u2_u2_u4_U77 (.A2( u2_u2_X_25 ) , .A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n104 ) );
  AND2_X1 u2_u2_u4_U78 (.A1( u2_u2_X_30 ) , .A2( u2_u2_u4_n176 ) , .ZN( u2_u2_u4_n99 ) );
  AND2_X1 u2_u2_u4_U79 (.A1( u2_u2_X_26 ) , .ZN( u2_u2_u4_n101 ) , .A2( u2_u2_u4_n177 ) );
  AOI21_X1 u2_u2_u4_U8 (.ZN( u2_u2_u4_n109 ) , .A( u2_u2_u4_n153 ) , .B1( u2_u2_u4_n159 ) , .B2( u2_u2_u4_n184 ) );
  AND2_X1 u2_u2_u4_U80 (.A1( u2_u2_X_27 ) , .A2( u2_u2_X_30 ) , .ZN( u2_u2_u4_n103 ) );
  INV_X1 u2_u2_u4_U81 (.A( u2_u2_X_28 ) , .ZN( u2_u2_u4_n169 ) );
  INV_X1 u2_u2_u4_U82 (.A( u2_u2_X_29 ) , .ZN( u2_u2_u4_n168 ) );
  INV_X1 u2_u2_u4_U83 (.A( u2_u2_X_25 ) , .ZN( u2_u2_u4_n177 ) );
  INV_X1 u2_u2_u4_U84 (.A( u2_u2_X_27 ) , .ZN( u2_u2_u4_n176 ) );
  NAND4_X1 u2_u2_u4_U85 (.ZN( u2_out2_25 ) , .A4( u2_u2_u4_n139 ) , .A3( u2_u2_u4_n140 ) , .A2( u2_u2_u4_n141 ) , .A1( u2_u2_u4_n142 ) );
  OAI21_X1 u2_u2_u4_U86 (.A( u2_u2_u4_n128 ) , .B2( u2_u2_u4_n129 ) , .B1( u2_u2_u4_n130 ) , .ZN( u2_u2_u4_n142 ) );
  OAI21_X1 u2_u2_u4_U87 (.B2( u2_u2_u4_n131 ) , .ZN( u2_u2_u4_n141 ) , .A( u2_u2_u4_n175 ) , .B1( u2_u2_u4_n183 ) );
  NAND4_X1 u2_u2_u4_U88 (.ZN( u2_out2_14 ) , .A4( u2_u2_u4_n124 ) , .A3( u2_u2_u4_n125 ) , .A2( u2_u2_u4_n126 ) , .A1( u2_u2_u4_n127 ) );
  AOI22_X1 u2_u2_u4_U89 (.B2( u2_u2_u4_n117 ) , .ZN( u2_u2_u4_n126 ) , .A1( u2_u2_u4_n129 ) , .B1( u2_u2_u4_n152 ) , .A2( u2_u2_u4_n175 ) );
  AOI211_X1 u2_u2_u4_U9 (.B( u2_u2_u4_n136 ) , .A( u2_u2_u4_n137 ) , .C2( u2_u2_u4_n138 ) , .ZN( u2_u2_u4_n139 ) , .C1( u2_u2_u4_n182 ) );
  AOI22_X1 u2_u2_u4_U90 (.ZN( u2_u2_u4_n125 ) , .B2( u2_u2_u4_n131 ) , .A2( u2_u2_u4_n132 ) , .B1( u2_u2_u4_n138 ) , .A1( u2_u2_u4_n178 ) );
  NAND4_X1 u2_u2_u4_U91 (.ZN( u2_out2_8 ) , .A4( u2_u2_u4_n110 ) , .A3( u2_u2_u4_n111 ) , .A2( u2_u2_u4_n112 ) , .A1( u2_u2_u4_n186 ) );
  NAND2_X1 u2_u2_u4_U92 (.ZN( u2_u2_u4_n112 ) , .A2( u2_u2_u4_n130 ) , .A1( u2_u2_u4_n150 ) );
  AOI22_X1 u2_u2_u4_U93 (.ZN( u2_u2_u4_n111 ) , .B2( u2_u2_u4_n132 ) , .A1( u2_u2_u4_n152 ) , .B1( u2_u2_u4_n178 ) , .A2( u2_u2_u4_n97 ) );
  AOI22_X1 u2_u2_u4_U94 (.B2( u2_u2_u4_n149 ) , .B1( u2_u2_u4_n150 ) , .A2( u2_u2_u4_n151 ) , .A1( u2_u2_u4_n152 ) , .ZN( u2_u2_u4_n167 ) );
  NOR4_X1 u2_u2_u4_U95 (.A4( u2_u2_u4_n162 ) , .A3( u2_u2_u4_n163 ) , .A2( u2_u2_u4_n164 ) , .A1( u2_u2_u4_n165 ) , .ZN( u2_u2_u4_n166 ) );
  NAND3_X1 u2_u2_u4_U96 (.ZN( u2_out2_3 ) , .A3( u2_u2_u4_n166 ) , .A1( u2_u2_u4_n167 ) , .A2( u2_u2_u4_n186 ) );
  NAND3_X1 u2_u2_u4_U97 (.A3( u2_u2_u4_n146 ) , .A2( u2_u2_u4_n147 ) , .A1( u2_u2_u4_n148 ) , .ZN( u2_u2_u4_n149 ) );
  NAND3_X1 u2_u2_u4_U98 (.A3( u2_u2_u4_n143 ) , .A2( u2_u2_u4_n144 ) , .A1( u2_u2_u4_n145 ) , .ZN( u2_u2_u4_n151 ) );
  NAND3_X1 u2_u2_u4_U99 (.A3( u2_u2_u4_n121 ) , .ZN( u2_u2_u4_n122 ) , .A2( u2_u2_u4_n144 ) , .A1( u2_u2_u4_n154 ) );
  XOR2_X1 u2_u3_U1 (.B( u2_K4_9 ) , .A( u2_R2_6 ) , .Z( u2_u3_X_9 ) );
  XOR2_X1 u2_u3_U10 (.B( u2_K4_45 ) , .A( u2_R2_30 ) , .Z( u2_u3_X_45 ) );
  XOR2_X1 u2_u3_U11 (.B( u2_K4_44 ) , .A( u2_R2_29 ) , .Z( u2_u3_X_44 ) );
  XOR2_X1 u2_u3_U12 (.B( u2_K4_43 ) , .A( u2_R2_28 ) , .Z( u2_u3_X_43 ) );
  XOR2_X1 u2_u3_U13 (.B( u2_K4_42 ) , .A( u2_R2_29 ) , .Z( u2_u3_X_42 ) );
  XOR2_X1 u2_u3_U14 (.B( u2_K4_41 ) , .A( u2_R2_28 ) , .Z( u2_u3_X_41 ) );
  XOR2_X1 u2_u3_U15 (.B( u2_K4_40 ) , .A( u2_R2_27 ) , .Z( u2_u3_X_40 ) );
  XOR2_X1 u2_u3_U16 (.B( u2_K4_3 ) , .A( u2_R2_2 ) , .Z( u2_u3_X_3 ) );
  XOR2_X1 u2_u3_U17 (.B( u2_K4_39 ) , .A( u2_R2_26 ) , .Z( u2_u3_X_39 ) );
  XOR2_X1 u2_u3_U18 (.B( u2_K4_38 ) , .A( u2_R2_25 ) , .Z( u2_u3_X_38 ) );
  XOR2_X1 u2_u3_U19 (.B( u2_K4_37 ) , .A( u2_R2_24 ) , .Z( u2_u3_X_37 ) );
  XOR2_X1 u2_u3_U2 (.B( u2_K4_8 ) , .A( u2_R2_5 ) , .Z( u2_u3_X_8 ) );
  XOR2_X1 u2_u3_U27 (.B( u2_K4_2 ) , .A( u2_R2_1 ) , .Z( u2_u3_X_2 ) );
  XOR2_X1 u2_u3_U3 (.B( u2_K4_7 ) , .A( u2_R2_4 ) , .Z( u2_u3_X_7 ) );
  XOR2_X1 u2_u3_U38 (.B( u2_K4_1 ) , .A( u2_R2_32 ) , .Z( u2_u3_X_1 ) );
  XOR2_X1 u2_u3_U4 (.B( u2_K4_6 ) , .A( u2_R2_5 ) , .Z( u2_u3_X_6 ) );
  XOR2_X1 u2_u3_U46 (.B( u2_K4_12 ) , .A( u2_R2_9 ) , .Z( u2_u3_X_12 ) );
  XOR2_X1 u2_u3_U47 (.B( u2_K4_11 ) , .A( u2_R2_8 ) , .Z( u2_u3_X_11 ) );
  XOR2_X1 u2_u3_U48 (.B( u2_K4_10 ) , .A( u2_R2_7 ) , .Z( u2_u3_X_10 ) );
  XOR2_X1 u2_u3_U5 (.B( u2_K4_5 ) , .A( u2_R2_4 ) , .Z( u2_u3_X_5 ) );
  XOR2_X1 u2_u3_U6 (.B( u2_K4_4 ) , .A( u2_R2_3 ) , .Z( u2_u3_X_4 ) );
  XOR2_X1 u2_u3_U7 (.B( u2_K4_48 ) , .A( u2_R2_1 ) , .Z( u2_u3_X_48 ) );
  XOR2_X1 u2_u3_U8 (.B( u2_K4_47 ) , .A( u2_R2_32 ) , .Z( u2_u3_X_47 ) );
  XOR2_X1 u2_u3_U9 (.B( u2_K4_46 ) , .A( u2_R2_31 ) , .Z( u2_u3_X_46 ) );
  AND3_X1 u2_u3_u0_U10 (.A2( u2_u3_u0_n112 ) , .ZN( u2_u3_u0_n127 ) , .A3( u2_u3_u0_n130 ) , .A1( u2_u3_u0_n148 ) );
  NAND2_X1 u2_u3_u0_U11 (.ZN( u2_u3_u0_n113 ) , .A1( u2_u3_u0_n139 ) , .A2( u2_u3_u0_n149 ) );
  AND2_X1 u2_u3_u0_U12 (.ZN( u2_u3_u0_n107 ) , .A1( u2_u3_u0_n130 ) , .A2( u2_u3_u0_n140 ) );
  AND2_X1 u2_u3_u0_U13 (.A2( u2_u3_u0_n129 ) , .A1( u2_u3_u0_n130 ) , .ZN( u2_u3_u0_n151 ) );
  AND2_X1 u2_u3_u0_U14 (.A1( u2_u3_u0_n108 ) , .A2( u2_u3_u0_n125 ) , .ZN( u2_u3_u0_n145 ) );
  INV_X1 u2_u3_u0_U15 (.A( u2_u3_u0_n143 ) , .ZN( u2_u3_u0_n173 ) );
  NOR2_X1 u2_u3_u0_U16 (.A2( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n147 ) , .A1( u2_u3_u0_n160 ) );
  INV_X1 u2_u3_u0_U17 (.ZN( u2_u3_u0_n172 ) , .A( u2_u3_u0_n88 ) );
  OAI222_X1 u2_u3_u0_U18 (.C1( u2_u3_u0_n108 ) , .A1( u2_u3_u0_n125 ) , .B2( u2_u3_u0_n128 ) , .B1( u2_u3_u0_n144 ) , .A2( u2_u3_u0_n158 ) , .C2( u2_u3_u0_n161 ) , .ZN( u2_u3_u0_n88 ) );
  AOI21_X1 u2_u3_u0_U19 (.B1( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n132 ) , .A( u2_u3_u0_n165 ) , .B2( u2_u3_u0_n93 ) );
  INV_X1 u2_u3_u0_U20 (.A( u2_u3_u0_n142 ) , .ZN( u2_u3_u0_n165 ) );
  OAI22_X1 u2_u3_u0_U21 (.B1( u2_u3_u0_n125 ) , .ZN( u2_u3_u0_n126 ) , .A1( u2_u3_u0_n138 ) , .A2( u2_u3_u0_n146 ) , .B2( u2_u3_u0_n147 ) );
  OAI22_X1 u2_u3_u0_U22 (.B1( u2_u3_u0_n131 ) , .A1( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n147 ) , .A2( u2_u3_u0_n90 ) , .ZN( u2_u3_u0_n91 ) );
  AND3_X1 u2_u3_u0_U23 (.A3( u2_u3_u0_n121 ) , .A2( u2_u3_u0_n125 ) , .A1( u2_u3_u0_n148 ) , .ZN( u2_u3_u0_n90 ) );
  INV_X1 u2_u3_u0_U24 (.A( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n161 ) );
  AOI22_X1 u2_u3_u0_U25 (.B2( u2_u3_u0_n109 ) , .A2( u2_u3_u0_n110 ) , .ZN( u2_u3_u0_n111 ) , .B1( u2_u3_u0_n118 ) , .A1( u2_u3_u0_n160 ) );
  NAND2_X1 u2_u3_u0_U26 (.A2( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n140 ) , .A1( u2_u3_u0_n94 ) );
  INV_X1 u2_u3_u0_U27 (.A( u2_u3_u0_n118 ) , .ZN( u2_u3_u0_n158 ) );
  AOI21_X1 u2_u3_u0_U28 (.ZN( u2_u3_u0_n104 ) , .B1( u2_u3_u0_n107 ) , .B2( u2_u3_u0_n141 ) , .A( u2_u3_u0_n144 ) );
  AOI21_X1 u2_u3_u0_U29 (.B1( u2_u3_u0_n127 ) , .B2( u2_u3_u0_n129 ) , .A( u2_u3_u0_n138 ) , .ZN( u2_u3_u0_n96 ) );
  INV_X1 u2_u3_u0_U3 (.A( u2_u3_u0_n113 ) , .ZN( u2_u3_u0_n166 ) );
  NOR2_X1 u2_u3_u0_U30 (.A1( u2_u3_u0_n120 ) , .ZN( u2_u3_u0_n143 ) , .A2( u2_u3_u0_n167 ) );
  OAI221_X1 u2_u3_u0_U31 (.C1( u2_u3_u0_n112 ) , .ZN( u2_u3_u0_n120 ) , .B1( u2_u3_u0_n138 ) , .B2( u2_u3_u0_n141 ) , .C2( u2_u3_u0_n147 ) , .A( u2_u3_u0_n172 ) );
  AOI21_X1 u2_u3_u0_U32 (.ZN( u2_u3_u0_n116 ) , .B2( u2_u3_u0_n142 ) , .A( u2_u3_u0_n144 ) , .B1( u2_u3_u0_n166 ) );
  NAND2_X1 u2_u3_u0_U33 (.A1( u2_u3_u0_n101 ) , .A2( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n150 ) );
  INV_X1 u2_u3_u0_U34 (.A( u2_u3_u0_n138 ) , .ZN( u2_u3_u0_n160 ) );
  NAND2_X1 u2_u3_u0_U35 (.ZN( u2_u3_u0_n108 ) , .A1( u2_u3_u0_n92 ) , .A2( u2_u3_u0_n94 ) );
  NAND2_X1 u2_u3_u0_U36 (.A2( u2_u3_u0_n102 ) , .A1( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n149 ) );
  NAND2_X1 u2_u3_u0_U37 (.A1( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n130 ) , .A2( u2_u3_u0_n94 ) );
  NAND2_X1 u2_u3_u0_U38 (.A2( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n114 ) , .A1( u2_u3_u0_n92 ) );
  NAND2_X1 u2_u3_u0_U39 (.A2( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n121 ) , .A1( u2_u3_u0_n93 ) );
  AOI21_X1 u2_u3_u0_U4 (.B2( u2_u3_u0_n131 ) , .ZN( u2_u3_u0_n134 ) , .B1( u2_u3_u0_n151 ) , .A( u2_u3_u0_n158 ) );
  NAND2_X1 u2_u3_u0_U40 (.ZN( u2_u3_u0_n112 ) , .A2( u2_u3_u0_n92 ) , .A1( u2_u3_u0_n93 ) );
  OR3_X1 u2_u3_u0_U41 (.A3( u2_u3_u0_n152 ) , .A2( u2_u3_u0_n153 ) , .A1( u2_u3_u0_n154 ) , .ZN( u2_u3_u0_n155 ) );
  AOI21_X1 u2_u3_u0_U42 (.A( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n145 ) , .B1( u2_u3_u0_n146 ) , .ZN( u2_u3_u0_n154 ) );
  AOI21_X1 u2_u3_u0_U43 (.B2( u2_u3_u0_n150 ) , .B1( u2_u3_u0_n151 ) , .ZN( u2_u3_u0_n152 ) , .A( u2_u3_u0_n158 ) );
  AOI21_X1 u2_u3_u0_U44 (.A( u2_u3_u0_n147 ) , .B2( u2_u3_u0_n148 ) , .B1( u2_u3_u0_n149 ) , .ZN( u2_u3_u0_n153 ) );
  INV_X1 u2_u3_u0_U45 (.ZN( u2_u3_u0_n171 ) , .A( u2_u3_u0_n99 ) );
  OAI211_X1 u2_u3_u0_U46 (.C2( u2_u3_u0_n140 ) , .C1( u2_u3_u0_n161 ) , .A( u2_u3_u0_n169 ) , .B( u2_u3_u0_n98 ) , .ZN( u2_u3_u0_n99 ) );
  AOI211_X1 u2_u3_u0_U47 (.C1( u2_u3_u0_n118 ) , .A( u2_u3_u0_n123 ) , .B( u2_u3_u0_n96 ) , .C2( u2_u3_u0_n97 ) , .ZN( u2_u3_u0_n98 ) );
  INV_X1 u2_u3_u0_U48 (.ZN( u2_u3_u0_n169 ) , .A( u2_u3_u0_n91 ) );
  NOR2_X1 u2_u3_u0_U49 (.A2( u2_u3_X_2 ) , .ZN( u2_u3_u0_n103 ) , .A1( u2_u3_u0_n164 ) );
  NOR2_X1 u2_u3_u0_U5 (.A1( u2_u3_u0_n108 ) , .ZN( u2_u3_u0_n123 ) , .A2( u2_u3_u0_n158 ) );
  NOR2_X1 u2_u3_u0_U50 (.A2( u2_u3_X_1 ) , .A1( u2_u3_X_2 ) , .ZN( u2_u3_u0_n92 ) );
  NOR2_X1 u2_u3_u0_U51 (.A2( u2_u3_X_4 ) , .A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n118 ) );
  NOR2_X1 u2_u3_u0_U52 (.A2( u2_u3_X_1 ) , .ZN( u2_u3_u0_n101 ) , .A1( u2_u3_u0_n163 ) );
  NAND2_X1 u2_u3_u0_U53 (.A2( u2_u3_X_4 ) , .A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n144 ) );
  NOR2_X1 u2_u3_u0_U54 (.A2( u2_u3_X_5 ) , .ZN( u2_u3_u0_n136 ) , .A1( u2_u3_u0_n159 ) );
  NAND2_X1 u2_u3_u0_U55 (.A1( u2_u3_X_5 ) , .ZN( u2_u3_u0_n138 ) , .A2( u2_u3_u0_n159 ) );
  NOR2_X1 u2_u3_u0_U56 (.A2( u2_u3_X_6 ) , .ZN( u2_u3_u0_n100 ) , .A1( u2_u3_u0_n162 ) );
  AND2_X1 u2_u3_u0_U57 (.A2( u2_u3_X_3 ) , .A1( u2_u3_X_6 ) , .ZN( u2_u3_u0_n102 ) );
  AND2_X1 u2_u3_u0_U58 (.A1( u2_u3_X_6 ) , .A2( u2_u3_u0_n162 ) , .ZN( u2_u3_u0_n93 ) );
  INV_X1 u2_u3_u0_U59 (.A( u2_u3_X_4 ) , .ZN( u2_u3_u0_n159 ) );
  OAI21_X1 u2_u3_u0_U6 (.B1( u2_u3_u0_n150 ) , .B2( u2_u3_u0_n158 ) , .A( u2_u3_u0_n172 ) , .ZN( u2_u3_u0_n89 ) );
  INV_X1 u2_u3_u0_U60 (.A( u2_u3_X_1 ) , .ZN( u2_u3_u0_n164 ) );
  INV_X1 u2_u3_u0_U61 (.A( u2_u3_X_2 ) , .ZN( u2_u3_u0_n163 ) );
  INV_X1 u2_u3_u0_U62 (.A( u2_u3_u0_n126 ) , .ZN( u2_u3_u0_n168 ) );
  AOI211_X1 u2_u3_u0_U63 (.B( u2_u3_u0_n133 ) , .A( u2_u3_u0_n134 ) , .C2( u2_u3_u0_n135 ) , .C1( u2_u3_u0_n136 ) , .ZN( u2_u3_u0_n137 ) );
  OR4_X1 u2_u3_u0_U64 (.ZN( u2_out3_17 ) , .A4( u2_u3_u0_n122 ) , .A2( u2_u3_u0_n123 ) , .A1( u2_u3_u0_n124 ) , .A3( u2_u3_u0_n170 ) );
  AOI21_X1 u2_u3_u0_U65 (.B2( u2_u3_u0_n107 ) , .ZN( u2_u3_u0_n124 ) , .B1( u2_u3_u0_n128 ) , .A( u2_u3_u0_n161 ) );
  INV_X1 u2_u3_u0_U66 (.A( u2_u3_u0_n111 ) , .ZN( u2_u3_u0_n170 ) );
  OR4_X1 u2_u3_u0_U67 (.ZN( u2_out3_31 ) , .A4( u2_u3_u0_n155 ) , .A2( u2_u3_u0_n156 ) , .A1( u2_u3_u0_n157 ) , .A3( u2_u3_u0_n173 ) );
  AOI21_X1 u2_u3_u0_U68 (.A( u2_u3_u0_n138 ) , .B2( u2_u3_u0_n139 ) , .B1( u2_u3_u0_n140 ) , .ZN( u2_u3_u0_n157 ) );
  AOI21_X1 u2_u3_u0_U69 (.B2( u2_u3_u0_n141 ) , .B1( u2_u3_u0_n142 ) , .ZN( u2_u3_u0_n156 ) , .A( u2_u3_u0_n161 ) );
  AOI21_X1 u2_u3_u0_U7 (.B1( u2_u3_u0_n114 ) , .ZN( u2_u3_u0_n115 ) , .B2( u2_u3_u0_n129 ) , .A( u2_u3_u0_n161 ) );
  INV_X1 u2_u3_u0_U70 (.ZN( u2_u3_u0_n174 ) , .A( u2_u3_u0_n89 ) );
  AOI211_X1 u2_u3_u0_U71 (.B( u2_u3_u0_n104 ) , .A( u2_u3_u0_n105 ) , .ZN( u2_u3_u0_n106 ) , .C2( u2_u3_u0_n113 ) , .C1( u2_u3_u0_n160 ) );
  AOI211_X1 u2_u3_u0_U72 (.B( u2_u3_u0_n115 ) , .A( u2_u3_u0_n116 ) , .C2( u2_u3_u0_n117 ) , .C1( u2_u3_u0_n118 ) , .ZN( u2_u3_u0_n119 ) );
  NAND2_X1 u2_u3_u0_U73 (.A2( u2_u3_u0_n100 ) , .ZN( u2_u3_u0_n131 ) , .A1( u2_u3_u0_n92 ) );
  NAND2_X1 u2_u3_u0_U74 (.A1( u2_u3_u0_n100 ) , .A2( u2_u3_u0_n103 ) , .ZN( u2_u3_u0_n125 ) );
  NAND2_X1 u2_u3_u0_U75 (.A2( u2_u3_u0_n100 ) , .A1( u2_u3_u0_n101 ) , .ZN( u2_u3_u0_n139 ) );
  NOR2_X1 u2_u3_u0_U76 (.A2( u2_u3_X_3 ) , .A1( u2_u3_X_6 ) , .ZN( u2_u3_u0_n94 ) );
  INV_X1 u2_u3_u0_U77 (.A( u2_u3_X_3 ) , .ZN( u2_u3_u0_n162 ) );
  NOR2_X1 u2_u3_u0_U78 (.A1( u2_u3_u0_n163 ) , .A2( u2_u3_u0_n164 ) , .ZN( u2_u3_u0_n95 ) );
  OAI221_X1 u2_u3_u0_U79 (.C1( u2_u3_u0_n121 ) , .ZN( u2_u3_u0_n122 ) , .B2( u2_u3_u0_n127 ) , .A( u2_u3_u0_n143 ) , .B1( u2_u3_u0_n144 ) , .C2( u2_u3_u0_n147 ) );
  AND2_X1 u2_u3_u0_U8 (.A1( u2_u3_u0_n114 ) , .A2( u2_u3_u0_n121 ) , .ZN( u2_u3_u0_n146 ) );
  AOI21_X1 u2_u3_u0_U80 (.B1( u2_u3_u0_n132 ) , .ZN( u2_u3_u0_n133 ) , .A( u2_u3_u0_n144 ) , .B2( u2_u3_u0_n166 ) );
  OAI22_X1 u2_u3_u0_U81 (.ZN( u2_u3_u0_n105 ) , .A2( u2_u3_u0_n132 ) , .B1( u2_u3_u0_n146 ) , .A1( u2_u3_u0_n147 ) , .B2( u2_u3_u0_n161 ) );
  NAND2_X1 u2_u3_u0_U82 (.ZN( u2_u3_u0_n110 ) , .A2( u2_u3_u0_n132 ) , .A1( u2_u3_u0_n145 ) );
  INV_X1 u2_u3_u0_U83 (.A( u2_u3_u0_n119 ) , .ZN( u2_u3_u0_n167 ) );
  NAND2_X1 u2_u3_u0_U84 (.ZN( u2_u3_u0_n148 ) , .A1( u2_u3_u0_n93 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U85 (.A1( u2_u3_u0_n100 ) , .ZN( u2_u3_u0_n129 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U86 (.A1( u2_u3_u0_n102 ) , .ZN( u2_u3_u0_n128 ) , .A2( u2_u3_u0_n95 ) );
  NAND2_X1 u2_u3_u0_U87 (.ZN( u2_u3_u0_n142 ) , .A1( u2_u3_u0_n94 ) , .A2( u2_u3_u0_n95 ) );
  NAND3_X1 u2_u3_u0_U88 (.ZN( u2_out3_23 ) , .A3( u2_u3_u0_n137 ) , .A1( u2_u3_u0_n168 ) , .A2( u2_u3_u0_n171 ) );
  NAND3_X1 u2_u3_u0_U89 (.A3( u2_u3_u0_n127 ) , .A2( u2_u3_u0_n128 ) , .ZN( u2_u3_u0_n135 ) , .A1( u2_u3_u0_n150 ) );
  AND2_X1 u2_u3_u0_U9 (.A1( u2_u3_u0_n131 ) , .ZN( u2_u3_u0_n141 ) , .A2( u2_u3_u0_n150 ) );
  NAND3_X1 u2_u3_u0_U90 (.ZN( u2_u3_u0_n117 ) , .A3( u2_u3_u0_n132 ) , .A2( u2_u3_u0_n139 ) , .A1( u2_u3_u0_n148 ) );
  NAND3_X1 u2_u3_u0_U91 (.ZN( u2_u3_u0_n109 ) , .A2( u2_u3_u0_n114 ) , .A3( u2_u3_u0_n140 ) , .A1( u2_u3_u0_n149 ) );
  NAND3_X1 u2_u3_u0_U92 (.ZN( u2_out3_9 ) , .A3( u2_u3_u0_n106 ) , .A2( u2_u3_u0_n171 ) , .A1( u2_u3_u0_n174 ) );
  NAND3_X1 u2_u3_u0_U93 (.A2( u2_u3_u0_n128 ) , .A1( u2_u3_u0_n132 ) , .A3( u2_u3_u0_n146 ) , .ZN( u2_u3_u0_n97 ) );
  NOR2_X1 u2_u3_u1_U10 (.A1( u2_u3_u1_n112 ) , .A2( u2_u3_u1_n116 ) , .ZN( u2_u3_u1_n118 ) );
  NAND3_X1 u2_u3_u1_U100 (.ZN( u2_u3_u1_n113 ) , .A1( u2_u3_u1_n120 ) , .A3( u2_u3_u1_n133 ) , .A2( u2_u3_u1_n155 ) );
  OAI21_X1 u2_u3_u1_U11 (.ZN( u2_u3_u1_n101 ) , .B1( u2_u3_u1_n141 ) , .A( u2_u3_u1_n146 ) , .B2( u2_u3_u1_n183 ) );
  AOI21_X1 u2_u3_u1_U12 (.B2( u2_u3_u1_n155 ) , .B1( u2_u3_u1_n156 ) , .ZN( u2_u3_u1_n157 ) , .A( u2_u3_u1_n174 ) );
  NAND2_X1 u2_u3_u1_U13 (.ZN( u2_u3_u1_n140 ) , .A2( u2_u3_u1_n150 ) , .A1( u2_u3_u1_n155 ) );
  NAND2_X1 u2_u3_u1_U14 (.A1( u2_u3_u1_n131 ) , .ZN( u2_u3_u1_n147 ) , .A2( u2_u3_u1_n153 ) );
  INV_X1 u2_u3_u1_U15 (.A( u2_u3_u1_n139 ) , .ZN( u2_u3_u1_n174 ) );
  OR4_X1 u2_u3_u1_U16 (.A4( u2_u3_u1_n106 ) , .A3( u2_u3_u1_n107 ) , .ZN( u2_u3_u1_n108 ) , .A1( u2_u3_u1_n117 ) , .A2( u2_u3_u1_n184 ) );
  AOI21_X1 u2_u3_u1_U17 (.ZN( u2_u3_u1_n106 ) , .A( u2_u3_u1_n112 ) , .B1( u2_u3_u1_n154 ) , .B2( u2_u3_u1_n156 ) );
  INV_X1 u2_u3_u1_U18 (.A( u2_u3_u1_n101 ) , .ZN( u2_u3_u1_n184 ) );
  AOI21_X1 u2_u3_u1_U19 (.ZN( u2_u3_u1_n107 ) , .B1( u2_u3_u1_n134 ) , .B2( u2_u3_u1_n149 ) , .A( u2_u3_u1_n174 ) );
  INV_X1 u2_u3_u1_U20 (.A( u2_u3_u1_n112 ) , .ZN( u2_u3_u1_n171 ) );
  NAND2_X1 u2_u3_u1_U21 (.ZN( u2_u3_u1_n141 ) , .A1( u2_u3_u1_n153 ) , .A2( u2_u3_u1_n156 ) );
  AND2_X1 u2_u3_u1_U22 (.A1( u2_u3_u1_n123 ) , .ZN( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n161 ) );
  NAND2_X1 u2_u3_u1_U23 (.A2( u2_u3_u1_n115 ) , .A1( u2_u3_u1_n116 ) , .ZN( u2_u3_u1_n148 ) );
  NAND2_X1 u2_u3_u1_U24 (.A2( u2_u3_u1_n133 ) , .A1( u2_u3_u1_n135 ) , .ZN( u2_u3_u1_n159 ) );
  NAND2_X1 u2_u3_u1_U25 (.A2( u2_u3_u1_n115 ) , .A1( u2_u3_u1_n120 ) , .ZN( u2_u3_u1_n132 ) );
  INV_X1 u2_u3_u1_U26 (.A( u2_u3_u1_n154 ) , .ZN( u2_u3_u1_n178 ) );
  INV_X1 u2_u3_u1_U27 (.A( u2_u3_u1_n151 ) , .ZN( u2_u3_u1_n183 ) );
  AND2_X1 u2_u3_u1_U28 (.A1( u2_u3_u1_n129 ) , .A2( u2_u3_u1_n133 ) , .ZN( u2_u3_u1_n149 ) );
  INV_X1 u2_u3_u1_U29 (.A( u2_u3_u1_n131 ) , .ZN( u2_u3_u1_n180 ) );
  INV_X1 u2_u3_u1_U3 (.A( u2_u3_u1_n159 ) , .ZN( u2_u3_u1_n182 ) );
  AOI221_X1 u2_u3_u1_U30 (.B1( u2_u3_u1_n140 ) , .ZN( u2_u3_u1_n167 ) , .B2( u2_u3_u1_n172 ) , .C2( u2_u3_u1_n175 ) , .C1( u2_u3_u1_n178 ) , .A( u2_u3_u1_n188 ) );
  INV_X1 u2_u3_u1_U31 (.ZN( u2_u3_u1_n188 ) , .A( u2_u3_u1_n97 ) );
  AOI211_X1 u2_u3_u1_U32 (.A( u2_u3_u1_n118 ) , .C1( u2_u3_u1_n132 ) , .C2( u2_u3_u1_n139 ) , .B( u2_u3_u1_n96 ) , .ZN( u2_u3_u1_n97 ) );
  AOI21_X1 u2_u3_u1_U33 (.B2( u2_u3_u1_n121 ) , .B1( u2_u3_u1_n135 ) , .A( u2_u3_u1_n152 ) , .ZN( u2_u3_u1_n96 ) );
  OAI221_X1 u2_u3_u1_U34 (.A( u2_u3_u1_n119 ) , .C2( u2_u3_u1_n129 ) , .ZN( u2_u3_u1_n138 ) , .B2( u2_u3_u1_n152 ) , .C1( u2_u3_u1_n174 ) , .B1( u2_u3_u1_n187 ) );
  INV_X1 u2_u3_u1_U35 (.A( u2_u3_u1_n148 ) , .ZN( u2_u3_u1_n187 ) );
  AOI211_X1 u2_u3_u1_U36 (.B( u2_u3_u1_n117 ) , .A( u2_u3_u1_n118 ) , .ZN( u2_u3_u1_n119 ) , .C2( u2_u3_u1_n146 ) , .C1( u2_u3_u1_n159 ) );
  NOR2_X1 u2_u3_u1_U37 (.A1( u2_u3_u1_n168 ) , .A2( u2_u3_u1_n176 ) , .ZN( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U38 (.A1( u2_u3_u1_n128 ) , .ZN( u2_u3_u1_n146 ) , .A2( u2_u3_u1_n160 ) );
  NAND2_X1 u2_u3_u1_U39 (.A2( u2_u3_u1_n112 ) , .ZN( u2_u3_u1_n139 ) , .A1( u2_u3_u1_n152 ) );
  AOI221_X1 u2_u3_u1_U4 (.A( u2_u3_u1_n138 ) , .C2( u2_u3_u1_n139 ) , .C1( u2_u3_u1_n140 ) , .B2( u2_u3_u1_n141 ) , .ZN( u2_u3_u1_n142 ) , .B1( u2_u3_u1_n175 ) );
  NAND2_X1 u2_u3_u1_U40 (.A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n156 ) , .A2( u2_u3_u1_n99 ) );
  NOR2_X1 u2_u3_u1_U41 (.ZN( u2_u3_u1_n117 ) , .A1( u2_u3_u1_n121 ) , .A2( u2_u3_u1_n160 ) );
  OAI21_X1 u2_u3_u1_U42 (.B2( u2_u3_u1_n123 ) , .ZN( u2_u3_u1_n145 ) , .B1( u2_u3_u1_n160 ) , .A( u2_u3_u1_n185 ) );
  INV_X1 u2_u3_u1_U43 (.A( u2_u3_u1_n122 ) , .ZN( u2_u3_u1_n185 ) );
  AOI21_X1 u2_u3_u1_U44 (.B2( u2_u3_u1_n120 ) , .B1( u2_u3_u1_n121 ) , .ZN( u2_u3_u1_n122 ) , .A( u2_u3_u1_n128 ) );
  AOI21_X1 u2_u3_u1_U45 (.A( u2_u3_u1_n128 ) , .B2( u2_u3_u1_n129 ) , .ZN( u2_u3_u1_n130 ) , .B1( u2_u3_u1_n150 ) );
  NAND2_X1 u2_u3_u1_U46 (.ZN( u2_u3_u1_n112 ) , .A1( u2_u3_u1_n169 ) , .A2( u2_u3_u1_n170 ) );
  NAND2_X1 u2_u3_u1_U47 (.ZN( u2_u3_u1_n129 ) , .A2( u2_u3_u1_n95 ) , .A1( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U48 (.A1( u2_u3_u1_n102 ) , .ZN( u2_u3_u1_n154 ) , .A2( u2_u3_u1_n99 ) );
  NAND2_X1 u2_u3_u1_U49 (.A2( u2_u3_u1_n100 ) , .ZN( u2_u3_u1_n135 ) , .A1( u2_u3_u1_n99 ) );
  AOI211_X1 u2_u3_u1_U5 (.ZN( u2_u3_u1_n124 ) , .A( u2_u3_u1_n138 ) , .C2( u2_u3_u1_n139 ) , .B( u2_u3_u1_n145 ) , .C1( u2_u3_u1_n147 ) );
  AOI21_X1 u2_u3_u1_U50 (.A( u2_u3_u1_n152 ) , .B2( u2_u3_u1_n153 ) , .B1( u2_u3_u1_n154 ) , .ZN( u2_u3_u1_n158 ) );
  INV_X1 u2_u3_u1_U51 (.A( u2_u3_u1_n160 ) , .ZN( u2_u3_u1_n175 ) );
  NAND2_X1 u2_u3_u1_U52 (.A1( u2_u3_u1_n100 ) , .ZN( u2_u3_u1_n116 ) , .A2( u2_u3_u1_n95 ) );
  NAND2_X1 u2_u3_u1_U53 (.A1( u2_u3_u1_n102 ) , .ZN( u2_u3_u1_n131 ) , .A2( u2_u3_u1_n95 ) );
  NAND2_X1 u2_u3_u1_U54 (.A2( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n121 ) , .A1( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U55 (.A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n153 ) , .A2( u2_u3_u1_n98 ) );
  NAND2_X1 u2_u3_u1_U56 (.A2( u2_u3_u1_n104 ) , .A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n133 ) );
  NAND2_X1 u2_u3_u1_U57 (.ZN( u2_u3_u1_n150 ) , .A2( u2_u3_u1_n98 ) , .A1( u2_u3_u1_n99 ) );
  NAND2_X1 u2_u3_u1_U58 (.A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n155 ) , .A2( u2_u3_u1_n95 ) );
  OAI21_X1 u2_u3_u1_U59 (.ZN( u2_u3_u1_n109 ) , .B1( u2_u3_u1_n129 ) , .B2( u2_u3_u1_n160 ) , .A( u2_u3_u1_n167 ) );
  AOI22_X1 u2_u3_u1_U6 (.B2( u2_u3_u1_n113 ) , .A2( u2_u3_u1_n114 ) , .ZN( u2_u3_u1_n125 ) , .A1( u2_u3_u1_n171 ) , .B1( u2_u3_u1_n173 ) );
  NAND2_X1 u2_u3_u1_U60 (.A2( u2_u3_u1_n100 ) , .A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n120 ) );
  NAND2_X1 u2_u3_u1_U61 (.A1( u2_u3_u1_n102 ) , .A2( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n115 ) );
  NAND2_X1 u2_u3_u1_U62 (.A2( u2_u3_u1_n100 ) , .A1( u2_u3_u1_n104 ) , .ZN( u2_u3_u1_n151 ) );
  NAND2_X1 u2_u3_u1_U63 (.A2( u2_u3_u1_n103 ) , .A1( u2_u3_u1_n105 ) , .ZN( u2_u3_u1_n161 ) );
  INV_X1 u2_u3_u1_U64 (.A( u2_u3_u1_n152 ) , .ZN( u2_u3_u1_n173 ) );
  INV_X1 u2_u3_u1_U65 (.A( u2_u3_u1_n128 ) , .ZN( u2_u3_u1_n172 ) );
  NAND2_X1 u2_u3_u1_U66 (.A2( u2_u3_u1_n102 ) , .A1( u2_u3_u1_n103 ) , .ZN( u2_u3_u1_n123 ) );
  AOI211_X1 u2_u3_u1_U67 (.B( u2_u3_u1_n162 ) , .A( u2_u3_u1_n163 ) , .C2( u2_u3_u1_n164 ) , .ZN( u2_u3_u1_n165 ) , .C1( u2_u3_u1_n171 ) );
  AOI21_X1 u2_u3_u1_U68 (.A( u2_u3_u1_n160 ) , .B2( u2_u3_u1_n161 ) , .ZN( u2_u3_u1_n162 ) , .B1( u2_u3_u1_n182 ) );
  OR2_X1 u2_u3_u1_U69 (.A2( u2_u3_u1_n157 ) , .A1( u2_u3_u1_n158 ) , .ZN( u2_u3_u1_n163 ) );
  NAND2_X1 u2_u3_u1_U7 (.ZN( u2_u3_u1_n114 ) , .A1( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n156 ) );
  NOR2_X1 u2_u3_u1_U70 (.A2( u2_u3_X_7 ) , .A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n95 ) );
  NOR2_X1 u2_u3_u1_U71 (.A1( u2_u3_X_12 ) , .A2( u2_u3_X_9 ) , .ZN( u2_u3_u1_n100 ) );
  NOR2_X1 u2_u3_u1_U72 (.A2( u2_u3_X_8 ) , .A1( u2_u3_u1_n177 ) , .ZN( u2_u3_u1_n99 ) );
  NOR2_X1 u2_u3_u1_U73 (.A2( u2_u3_X_12 ) , .ZN( u2_u3_u1_n102 ) , .A1( u2_u3_u1_n176 ) );
  NOR2_X1 u2_u3_u1_U74 (.A2( u2_u3_X_9 ) , .ZN( u2_u3_u1_n105 ) , .A1( u2_u3_u1_n168 ) );
  NAND2_X1 u2_u3_u1_U75 (.A1( u2_u3_X_10 ) , .ZN( u2_u3_u1_n160 ) , .A2( u2_u3_u1_n169 ) );
  NAND2_X1 u2_u3_u1_U76 (.A2( u2_u3_X_10 ) , .A1( u2_u3_X_11 ) , .ZN( u2_u3_u1_n152 ) );
  NAND2_X1 u2_u3_u1_U77 (.A1( u2_u3_X_11 ) , .ZN( u2_u3_u1_n128 ) , .A2( u2_u3_u1_n170 ) );
  AND2_X1 u2_u3_u1_U78 (.A2( u2_u3_X_7 ) , .A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n104 ) );
  AND2_X1 u2_u3_u1_U79 (.A1( u2_u3_X_8 ) , .ZN( u2_u3_u1_n103 ) , .A2( u2_u3_u1_n177 ) );
  AOI22_X1 u2_u3_u1_U8 (.B2( u2_u3_u1_n136 ) , .A2( u2_u3_u1_n137 ) , .ZN( u2_u3_u1_n143 ) , .A1( u2_u3_u1_n171 ) , .B1( u2_u3_u1_n173 ) );
  INV_X1 u2_u3_u1_U80 (.A( u2_u3_X_10 ) , .ZN( u2_u3_u1_n170 ) );
  INV_X1 u2_u3_u1_U81 (.A( u2_u3_X_9 ) , .ZN( u2_u3_u1_n176 ) );
  INV_X1 u2_u3_u1_U82 (.A( u2_u3_X_11 ) , .ZN( u2_u3_u1_n169 ) );
  INV_X1 u2_u3_u1_U83 (.A( u2_u3_X_12 ) , .ZN( u2_u3_u1_n168 ) );
  INV_X1 u2_u3_u1_U84 (.A( u2_u3_X_7 ) , .ZN( u2_u3_u1_n177 ) );
  NAND4_X1 u2_u3_u1_U85 (.ZN( u2_out3_28 ) , .A4( u2_u3_u1_n124 ) , .A3( u2_u3_u1_n125 ) , .A2( u2_u3_u1_n126 ) , .A1( u2_u3_u1_n127 ) );
  OAI21_X1 u2_u3_u1_U86 (.ZN( u2_u3_u1_n127 ) , .B2( u2_u3_u1_n139 ) , .B1( u2_u3_u1_n175 ) , .A( u2_u3_u1_n183 ) );
  OAI21_X1 u2_u3_u1_U87 (.ZN( u2_u3_u1_n126 ) , .B2( u2_u3_u1_n140 ) , .A( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n178 ) );
  NAND4_X1 u2_u3_u1_U88 (.ZN( u2_out3_18 ) , .A4( u2_u3_u1_n165 ) , .A3( u2_u3_u1_n166 ) , .A1( u2_u3_u1_n167 ) , .A2( u2_u3_u1_n186 ) );
  AOI22_X1 u2_u3_u1_U89 (.B2( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n147 ) , .A2( u2_u3_u1_n148 ) , .ZN( u2_u3_u1_n166 ) , .A1( u2_u3_u1_n172 ) );
  INV_X1 u2_u3_u1_U9 (.A( u2_u3_u1_n147 ) , .ZN( u2_u3_u1_n181 ) );
  INV_X1 u2_u3_u1_U90 (.A( u2_u3_u1_n145 ) , .ZN( u2_u3_u1_n186 ) );
  NAND4_X1 u2_u3_u1_U91 (.ZN( u2_out3_2 ) , .A4( u2_u3_u1_n142 ) , .A3( u2_u3_u1_n143 ) , .A2( u2_u3_u1_n144 ) , .A1( u2_u3_u1_n179 ) );
  OAI21_X1 u2_u3_u1_U92 (.B2( u2_u3_u1_n132 ) , .ZN( u2_u3_u1_n144 ) , .A( u2_u3_u1_n146 ) , .B1( u2_u3_u1_n180 ) );
  INV_X1 u2_u3_u1_U93 (.A( u2_u3_u1_n130 ) , .ZN( u2_u3_u1_n179 ) );
  OR4_X1 u2_u3_u1_U94 (.ZN( u2_out3_13 ) , .A4( u2_u3_u1_n108 ) , .A3( u2_u3_u1_n109 ) , .A2( u2_u3_u1_n110 ) , .A1( u2_u3_u1_n111 ) );
  AOI21_X1 u2_u3_u1_U95 (.ZN( u2_u3_u1_n111 ) , .A( u2_u3_u1_n128 ) , .B2( u2_u3_u1_n131 ) , .B1( u2_u3_u1_n135 ) );
  AOI21_X1 u2_u3_u1_U96 (.ZN( u2_u3_u1_n110 ) , .A( u2_u3_u1_n116 ) , .B1( u2_u3_u1_n152 ) , .B2( u2_u3_u1_n160 ) );
  NAND3_X1 u2_u3_u1_U97 (.A3( u2_u3_u1_n149 ) , .A2( u2_u3_u1_n150 ) , .A1( u2_u3_u1_n151 ) , .ZN( u2_u3_u1_n164 ) );
  NAND3_X1 u2_u3_u1_U98 (.A3( u2_u3_u1_n134 ) , .A2( u2_u3_u1_n135 ) , .ZN( u2_u3_u1_n136 ) , .A1( u2_u3_u1_n151 ) );
  NAND3_X1 u2_u3_u1_U99 (.A1( u2_u3_u1_n133 ) , .ZN( u2_u3_u1_n137 ) , .A2( u2_u3_u1_n154 ) , .A3( u2_u3_u1_n181 ) );
  INV_X1 u2_u3_u6_U10 (.ZN( u2_u3_u6_n172 ) , .A( u2_u3_u6_n88 ) );
  OAI21_X1 u2_u3_u6_U11 (.A( u2_u3_u6_n159 ) , .B1( u2_u3_u6_n169 ) , .B2( u2_u3_u6_n173 ) , .ZN( u2_u3_u6_n90 ) );
  AOI22_X1 u2_u3_u6_U12 (.A2( u2_u3_u6_n151 ) , .B2( u2_u3_u6_n161 ) , .A1( u2_u3_u6_n167 ) , .B1( u2_u3_u6_n170 ) , .ZN( u2_u3_u6_n89 ) );
  AOI21_X1 u2_u3_u6_U13 (.ZN( u2_u3_u6_n106 ) , .A( u2_u3_u6_n142 ) , .B2( u2_u3_u6_n159 ) , .B1( u2_u3_u6_n164 ) );
  INV_X1 u2_u3_u6_U14 (.A( u2_u3_u6_n155 ) , .ZN( u2_u3_u6_n161 ) );
  INV_X1 u2_u3_u6_U15 (.A( u2_u3_u6_n128 ) , .ZN( u2_u3_u6_n164 ) );
  NAND2_X1 u2_u3_u6_U16 (.ZN( u2_u3_u6_n110 ) , .A1( u2_u3_u6_n122 ) , .A2( u2_u3_u6_n129 ) );
  NAND2_X1 u2_u3_u6_U17 (.ZN( u2_u3_u6_n124 ) , .A2( u2_u3_u6_n146 ) , .A1( u2_u3_u6_n148 ) );
  INV_X1 u2_u3_u6_U18 (.A( u2_u3_u6_n132 ) , .ZN( u2_u3_u6_n171 ) );
  AND2_X1 u2_u3_u6_U19 (.A1( u2_u3_u6_n100 ) , .ZN( u2_u3_u6_n130 ) , .A2( u2_u3_u6_n147 ) );
  INV_X1 u2_u3_u6_U20 (.A( u2_u3_u6_n127 ) , .ZN( u2_u3_u6_n173 ) );
  INV_X1 u2_u3_u6_U21 (.A( u2_u3_u6_n121 ) , .ZN( u2_u3_u6_n167 ) );
  INV_X1 u2_u3_u6_U22 (.A( u2_u3_u6_n100 ) , .ZN( u2_u3_u6_n169 ) );
  INV_X1 u2_u3_u6_U23 (.A( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n170 ) );
  INV_X1 u2_u3_u6_U24 (.A( u2_u3_u6_n113 ) , .ZN( u2_u3_u6_n168 ) );
  AND2_X1 u2_u3_u6_U25 (.A1( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n119 ) , .ZN( u2_u3_u6_n133 ) );
  AND2_X1 u2_u3_u6_U26 (.A2( u2_u3_u6_n121 ) , .A1( u2_u3_u6_n122 ) , .ZN( u2_u3_u6_n131 ) );
  AND3_X1 u2_u3_u6_U27 (.ZN( u2_u3_u6_n120 ) , .A2( u2_u3_u6_n127 ) , .A1( u2_u3_u6_n132 ) , .A3( u2_u3_u6_n145 ) );
  INV_X1 u2_u3_u6_U28 (.A( u2_u3_u6_n146 ) , .ZN( u2_u3_u6_n163 ) );
  AOI222_X1 u2_u3_u6_U29 (.ZN( u2_u3_u6_n114 ) , .A1( u2_u3_u6_n118 ) , .A2( u2_u3_u6_n126 ) , .B2( u2_u3_u6_n151 ) , .C2( u2_u3_u6_n159 ) , .C1( u2_u3_u6_n168 ) , .B1( u2_u3_u6_n169 ) );
  INV_X1 u2_u3_u6_U3 (.A( u2_u3_u6_n110 ) , .ZN( u2_u3_u6_n166 ) );
  NOR2_X1 u2_u3_u6_U30 (.A1( u2_u3_u6_n162 ) , .A2( u2_u3_u6_n165 ) , .ZN( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U31 (.A1( u2_u3_u6_n144 ) , .ZN( u2_u3_u6_n151 ) , .A2( u2_u3_u6_n158 ) );
  NAND2_X1 u2_u3_u6_U32 (.ZN( u2_u3_u6_n132 ) , .A1( u2_u3_u6_n91 ) , .A2( u2_u3_u6_n97 ) );
  AOI22_X1 u2_u3_u6_U33 (.B2( u2_u3_u6_n110 ) , .B1( u2_u3_u6_n111 ) , .A1( u2_u3_u6_n112 ) , .ZN( u2_u3_u6_n115 ) , .A2( u2_u3_u6_n161 ) );
  NAND4_X1 u2_u3_u6_U34 (.A3( u2_u3_u6_n109 ) , .ZN( u2_u3_u6_n112 ) , .A4( u2_u3_u6_n132 ) , .A2( u2_u3_u6_n147 ) , .A1( u2_u3_u6_n166 ) );
  NOR2_X1 u2_u3_u6_U35 (.ZN( u2_u3_u6_n109 ) , .A1( u2_u3_u6_n170 ) , .A2( u2_u3_u6_n173 ) );
  NOR2_X1 u2_u3_u6_U36 (.A2( u2_u3_u6_n126 ) , .ZN( u2_u3_u6_n155 ) , .A1( u2_u3_u6_n160 ) );
  NAND2_X1 u2_u3_u6_U37 (.ZN( u2_u3_u6_n146 ) , .A2( u2_u3_u6_n94 ) , .A1( u2_u3_u6_n99 ) );
  AOI21_X1 u2_u3_u6_U38 (.A( u2_u3_u6_n144 ) , .B2( u2_u3_u6_n145 ) , .B1( u2_u3_u6_n146 ) , .ZN( u2_u3_u6_n150 ) );
  AOI211_X1 u2_u3_u6_U39 (.B( u2_u3_u6_n134 ) , .A( u2_u3_u6_n135 ) , .C1( u2_u3_u6_n136 ) , .ZN( u2_u3_u6_n137 ) , .C2( u2_u3_u6_n151 ) );
  INV_X1 u2_u3_u6_U4 (.A( u2_u3_u6_n142 ) , .ZN( u2_u3_u6_n174 ) );
  AOI21_X1 u2_u3_u6_U40 (.B2( u2_u3_u6_n132 ) , .B1( u2_u3_u6_n133 ) , .ZN( u2_u3_u6_n134 ) , .A( u2_u3_u6_n158 ) );
  NAND4_X1 u2_u3_u6_U41 (.A4( u2_u3_u6_n127 ) , .A3( u2_u3_u6_n128 ) , .A2( u2_u3_u6_n129 ) , .A1( u2_u3_u6_n130 ) , .ZN( u2_u3_u6_n136 ) );
  AOI21_X1 u2_u3_u6_U42 (.B1( u2_u3_u6_n131 ) , .ZN( u2_u3_u6_n135 ) , .A( u2_u3_u6_n144 ) , .B2( u2_u3_u6_n146 ) );
  INV_X1 u2_u3_u6_U43 (.A( u2_u3_u6_n111 ) , .ZN( u2_u3_u6_n158 ) );
  NAND2_X1 u2_u3_u6_U44 (.ZN( u2_u3_u6_n127 ) , .A1( u2_u3_u6_n91 ) , .A2( u2_u3_u6_n92 ) );
  NAND2_X1 u2_u3_u6_U45 (.ZN( u2_u3_u6_n129 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n96 ) );
  INV_X1 u2_u3_u6_U46 (.A( u2_u3_u6_n144 ) , .ZN( u2_u3_u6_n159 ) );
  NAND2_X1 u2_u3_u6_U47 (.ZN( u2_u3_u6_n145 ) , .A2( u2_u3_u6_n97 ) , .A1( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U48 (.ZN( u2_u3_u6_n148 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n94 ) );
  NAND2_X1 u2_u3_u6_U49 (.ZN( u2_u3_u6_n108 ) , .A2( u2_u3_u6_n139 ) , .A1( u2_u3_u6_n144 ) );
  NAND2_X1 u2_u3_u6_U5 (.A2( u2_u3_u6_n143 ) , .ZN( u2_u3_u6_n152 ) , .A1( u2_u3_u6_n166 ) );
  NAND2_X1 u2_u3_u6_U50 (.ZN( u2_u3_u6_n121 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n97 ) );
  NAND2_X1 u2_u3_u6_U51 (.ZN( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n95 ) );
  AND2_X1 u2_u3_u6_U52 (.ZN( u2_u3_u6_n118 ) , .A2( u2_u3_u6_n91 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U53 (.ZN( u2_u3_u6_n147 ) , .A2( u2_u3_u6_n98 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U54 (.ZN( u2_u3_u6_n128 ) , .A1( u2_u3_u6_n94 ) , .A2( u2_u3_u6_n96 ) );
  NAND2_X1 u2_u3_u6_U55 (.ZN( u2_u3_u6_n119 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U56 (.ZN( u2_u3_u6_n123 ) , .A2( u2_u3_u6_n91 ) , .A1( u2_u3_u6_n96 ) );
  NAND2_X1 u2_u3_u6_U57 (.ZN( u2_u3_u6_n100 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U58 (.ZN( u2_u3_u6_n122 ) , .A1( u2_u3_u6_n94 ) , .A2( u2_u3_u6_n97 ) );
  INV_X1 u2_u3_u6_U59 (.A( u2_u3_u6_n139 ) , .ZN( u2_u3_u6_n160 ) );
  AOI22_X1 u2_u3_u6_U6 (.B2( u2_u3_u6_n101 ) , .A1( u2_u3_u6_n102 ) , .ZN( u2_u3_u6_n103 ) , .B1( u2_u3_u6_n160 ) , .A2( u2_u3_u6_n161 ) );
  NAND2_X1 u2_u3_u6_U60 (.ZN( u2_u3_u6_n113 ) , .A1( u2_u3_u6_n96 ) , .A2( u2_u3_u6_n98 ) );
  NOR2_X1 u2_u3_u6_U61 (.A2( u2_u3_X_40 ) , .A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n126 ) );
  NOR2_X1 u2_u3_u6_U62 (.A2( u2_u3_X_39 ) , .A1( u2_u3_X_42 ) , .ZN( u2_u3_u6_n92 ) );
  NOR2_X1 u2_u3_u6_U63 (.A2( u2_u3_X_39 ) , .A1( u2_u3_u6_n156 ) , .ZN( u2_u3_u6_n97 ) );
  NOR2_X1 u2_u3_u6_U64 (.A2( u2_u3_X_38 ) , .A1( u2_u3_u6_n165 ) , .ZN( u2_u3_u6_n95 ) );
  NOR2_X1 u2_u3_u6_U65 (.A2( u2_u3_X_41 ) , .ZN( u2_u3_u6_n111 ) , .A1( u2_u3_u6_n157 ) );
  NOR2_X1 u2_u3_u6_U66 (.A2( u2_u3_X_37 ) , .A1( u2_u3_u6_n162 ) , .ZN( u2_u3_u6_n94 ) );
  NOR2_X1 u2_u3_u6_U67 (.A2( u2_u3_X_37 ) , .A1( u2_u3_X_38 ) , .ZN( u2_u3_u6_n91 ) );
  NAND2_X1 u2_u3_u6_U68 (.A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n144 ) , .A2( u2_u3_u6_n157 ) );
  NAND2_X1 u2_u3_u6_U69 (.A2( u2_u3_X_40 ) , .A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n139 ) );
  NOR2_X1 u2_u3_u6_U7 (.A1( u2_u3_u6_n118 ) , .ZN( u2_u3_u6_n143 ) , .A2( u2_u3_u6_n168 ) );
  AND2_X1 u2_u3_u6_U70 (.A1( u2_u3_X_39 ) , .A2( u2_u3_u6_n156 ) , .ZN( u2_u3_u6_n96 ) );
  AND2_X1 u2_u3_u6_U71 (.A1( u2_u3_X_39 ) , .A2( u2_u3_X_42 ) , .ZN( u2_u3_u6_n99 ) );
  INV_X1 u2_u3_u6_U72 (.A( u2_u3_X_40 ) , .ZN( u2_u3_u6_n157 ) );
  INV_X1 u2_u3_u6_U73 (.A( u2_u3_X_37 ) , .ZN( u2_u3_u6_n165 ) );
  INV_X1 u2_u3_u6_U74 (.A( u2_u3_X_38 ) , .ZN( u2_u3_u6_n162 ) );
  INV_X1 u2_u3_u6_U75 (.A( u2_u3_X_42 ) , .ZN( u2_u3_u6_n156 ) );
  NAND4_X1 u2_u3_u6_U76 (.ZN( u2_out3_32 ) , .A4( u2_u3_u6_n103 ) , .A3( u2_u3_u6_n104 ) , .A2( u2_u3_u6_n105 ) , .A1( u2_u3_u6_n106 ) );
  AOI22_X1 u2_u3_u6_U77 (.ZN( u2_u3_u6_n105 ) , .A2( u2_u3_u6_n108 ) , .A1( u2_u3_u6_n118 ) , .B2( u2_u3_u6_n126 ) , .B1( u2_u3_u6_n171 ) );
  AOI22_X1 u2_u3_u6_U78 (.ZN( u2_u3_u6_n104 ) , .A1( u2_u3_u6_n111 ) , .B1( u2_u3_u6_n124 ) , .B2( u2_u3_u6_n151 ) , .A2( u2_u3_u6_n93 ) );
  NAND4_X1 u2_u3_u6_U79 (.ZN( u2_out3_12 ) , .A4( u2_u3_u6_n114 ) , .A3( u2_u3_u6_n115 ) , .A2( u2_u3_u6_n116 ) , .A1( u2_u3_u6_n117 ) );
  AOI21_X1 u2_u3_u6_U8 (.B1( u2_u3_u6_n107 ) , .B2( u2_u3_u6_n132 ) , .A( u2_u3_u6_n158 ) , .ZN( u2_u3_u6_n88 ) );
  OAI22_X1 u2_u3_u6_U80 (.B2( u2_u3_u6_n111 ) , .ZN( u2_u3_u6_n116 ) , .B1( u2_u3_u6_n126 ) , .A2( u2_u3_u6_n164 ) , .A1( u2_u3_u6_n167 ) );
  OAI21_X1 u2_u3_u6_U81 (.A( u2_u3_u6_n108 ) , .ZN( u2_u3_u6_n117 ) , .B2( u2_u3_u6_n141 ) , .B1( u2_u3_u6_n163 ) );
  OAI211_X1 u2_u3_u6_U82 (.ZN( u2_out3_22 ) , .B( u2_u3_u6_n137 ) , .A( u2_u3_u6_n138 ) , .C2( u2_u3_u6_n139 ) , .C1( u2_u3_u6_n140 ) );
  AOI22_X1 u2_u3_u6_U83 (.B1( u2_u3_u6_n124 ) , .A2( u2_u3_u6_n125 ) , .A1( u2_u3_u6_n126 ) , .ZN( u2_u3_u6_n138 ) , .B2( u2_u3_u6_n161 ) );
  AND4_X1 u2_u3_u6_U84 (.A3( u2_u3_u6_n119 ) , .A1( u2_u3_u6_n120 ) , .A4( u2_u3_u6_n129 ) , .ZN( u2_u3_u6_n140 ) , .A2( u2_u3_u6_n143 ) );
  OAI211_X1 u2_u3_u6_U85 (.ZN( u2_out3_7 ) , .B( u2_u3_u6_n153 ) , .C2( u2_u3_u6_n154 ) , .C1( u2_u3_u6_n155 ) , .A( u2_u3_u6_n174 ) );
  NOR3_X1 u2_u3_u6_U86 (.A1( u2_u3_u6_n141 ) , .ZN( u2_u3_u6_n154 ) , .A3( u2_u3_u6_n164 ) , .A2( u2_u3_u6_n171 ) );
  AOI211_X1 u2_u3_u6_U87 (.B( u2_u3_u6_n149 ) , .A( u2_u3_u6_n150 ) , .C2( u2_u3_u6_n151 ) , .C1( u2_u3_u6_n152 ) , .ZN( u2_u3_u6_n153 ) );
  NAND3_X1 u2_u3_u6_U88 (.A2( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n125 ) , .A1( u2_u3_u6_n130 ) , .A3( u2_u3_u6_n131 ) );
  NAND3_X1 u2_u3_u6_U89 (.A3( u2_u3_u6_n133 ) , .ZN( u2_u3_u6_n141 ) , .A1( u2_u3_u6_n145 ) , .A2( u2_u3_u6_n148 ) );
  AOI21_X1 u2_u3_u6_U9 (.B2( u2_u3_u6_n147 ) , .B1( u2_u3_u6_n148 ) , .ZN( u2_u3_u6_n149 ) , .A( u2_u3_u6_n158 ) );
  NAND3_X1 u2_u3_u6_U90 (.ZN( u2_u3_u6_n101 ) , .A3( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n121 ) , .A1( u2_u3_u6_n127 ) );
  NAND3_X1 u2_u3_u6_U91 (.ZN( u2_u3_u6_n102 ) , .A3( u2_u3_u6_n130 ) , .A2( u2_u3_u6_n145 ) , .A1( u2_u3_u6_n166 ) );
  NAND3_X1 u2_u3_u6_U92 (.A3( u2_u3_u6_n113 ) , .A1( u2_u3_u6_n119 ) , .A2( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n93 ) );
  NAND3_X1 u2_u3_u6_U93 (.ZN( u2_u3_u6_n142 ) , .A2( u2_u3_u6_n172 ) , .A3( u2_u3_u6_n89 ) , .A1( u2_u3_u6_n90 ) );
  AND3_X1 u2_u3_u7_U10 (.A3( u2_u3_u7_n110 ) , .A2( u2_u3_u7_n127 ) , .A1( u2_u3_u7_n132 ) , .ZN( u2_u3_u7_n92 ) );
  OAI21_X1 u2_u3_u7_U11 (.A( u2_u3_u7_n161 ) , .B1( u2_u3_u7_n168 ) , .B2( u2_u3_u7_n173 ) , .ZN( u2_u3_u7_n91 ) );
  AOI211_X1 u2_u3_u7_U12 (.A( u2_u3_u7_n117 ) , .ZN( u2_u3_u7_n118 ) , .C2( u2_u3_u7_n126 ) , .C1( u2_u3_u7_n177 ) , .B( u2_u3_u7_n180 ) );
  OAI22_X1 u2_u3_u7_U13 (.B1( u2_u3_u7_n115 ) , .ZN( u2_u3_u7_n117 ) , .A2( u2_u3_u7_n133 ) , .A1( u2_u3_u7_n137 ) , .B2( u2_u3_u7_n162 ) );
  INV_X1 u2_u3_u7_U14 (.A( u2_u3_u7_n116 ) , .ZN( u2_u3_u7_n180 ) );
  NOR3_X1 u2_u3_u7_U15 (.ZN( u2_u3_u7_n115 ) , .A3( u2_u3_u7_n145 ) , .A2( u2_u3_u7_n168 ) , .A1( u2_u3_u7_n169 ) );
  OAI211_X1 u2_u3_u7_U16 (.B( u2_u3_u7_n122 ) , .A( u2_u3_u7_n123 ) , .C2( u2_u3_u7_n124 ) , .ZN( u2_u3_u7_n154 ) , .C1( u2_u3_u7_n162 ) );
  AOI222_X1 u2_u3_u7_U17 (.ZN( u2_u3_u7_n122 ) , .C2( u2_u3_u7_n126 ) , .C1( u2_u3_u7_n145 ) , .B1( u2_u3_u7_n161 ) , .A2( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n170 ) , .A1( u2_u3_u7_n176 ) );
  INV_X1 u2_u3_u7_U18 (.A( u2_u3_u7_n133 ) , .ZN( u2_u3_u7_n176 ) );
  NOR3_X1 u2_u3_u7_U19 (.A2( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n135 ) , .ZN( u2_u3_u7_n136 ) , .A3( u2_u3_u7_n171 ) );
  NOR2_X1 u2_u3_u7_U20 (.A1( u2_u3_u7_n130 ) , .A2( u2_u3_u7_n134 ) , .ZN( u2_u3_u7_n153 ) );
  INV_X1 u2_u3_u7_U21 (.A( u2_u3_u7_n101 ) , .ZN( u2_u3_u7_n165 ) );
  NOR2_X1 u2_u3_u7_U22 (.ZN( u2_u3_u7_n111 ) , .A2( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n169 ) );
  AOI21_X1 u2_u3_u7_U23 (.ZN( u2_u3_u7_n104 ) , .B2( u2_u3_u7_n112 ) , .B1( u2_u3_u7_n127 ) , .A( u2_u3_u7_n164 ) );
  AOI21_X1 u2_u3_u7_U24 (.ZN( u2_u3_u7_n106 ) , .B1( u2_u3_u7_n133 ) , .B2( u2_u3_u7_n146 ) , .A( u2_u3_u7_n162 ) );
  AOI21_X1 u2_u3_u7_U25 (.A( u2_u3_u7_n101 ) , .ZN( u2_u3_u7_n107 ) , .B2( u2_u3_u7_n128 ) , .B1( u2_u3_u7_n175 ) );
  INV_X1 u2_u3_u7_U26 (.A( u2_u3_u7_n138 ) , .ZN( u2_u3_u7_n171 ) );
  INV_X1 u2_u3_u7_U27 (.A( u2_u3_u7_n131 ) , .ZN( u2_u3_u7_n177 ) );
  INV_X1 u2_u3_u7_U28 (.A( u2_u3_u7_n110 ) , .ZN( u2_u3_u7_n174 ) );
  NAND2_X1 u2_u3_u7_U29 (.A1( u2_u3_u7_n129 ) , .A2( u2_u3_u7_n132 ) , .ZN( u2_u3_u7_n149 ) );
  OAI21_X1 u2_u3_u7_U3 (.ZN( u2_u3_u7_n159 ) , .A( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n171 ) , .B1( u2_u3_u7_n174 ) );
  NAND2_X1 u2_u3_u7_U30 (.A1( u2_u3_u7_n113 ) , .A2( u2_u3_u7_n124 ) , .ZN( u2_u3_u7_n130 ) );
  INV_X1 u2_u3_u7_U31 (.A( u2_u3_u7_n112 ) , .ZN( u2_u3_u7_n173 ) );
  INV_X1 u2_u3_u7_U32 (.A( u2_u3_u7_n128 ) , .ZN( u2_u3_u7_n168 ) );
  INV_X1 u2_u3_u7_U33 (.A( u2_u3_u7_n148 ) , .ZN( u2_u3_u7_n169 ) );
  INV_X1 u2_u3_u7_U34 (.A( u2_u3_u7_n127 ) , .ZN( u2_u3_u7_n179 ) );
  NOR2_X1 u2_u3_u7_U35 (.ZN( u2_u3_u7_n101 ) , .A2( u2_u3_u7_n150 ) , .A1( u2_u3_u7_n156 ) );
  AOI211_X1 u2_u3_u7_U36 (.B( u2_u3_u7_n154 ) , .A( u2_u3_u7_n155 ) , .C1( u2_u3_u7_n156 ) , .ZN( u2_u3_u7_n157 ) , .C2( u2_u3_u7_n172 ) );
  INV_X1 u2_u3_u7_U37 (.A( u2_u3_u7_n153 ) , .ZN( u2_u3_u7_n172 ) );
  AOI211_X1 u2_u3_u7_U38 (.B( u2_u3_u7_n139 ) , .A( u2_u3_u7_n140 ) , .C2( u2_u3_u7_n141 ) , .ZN( u2_u3_u7_n142 ) , .C1( u2_u3_u7_n156 ) );
  NAND4_X1 u2_u3_u7_U39 (.A3( u2_u3_u7_n127 ) , .A2( u2_u3_u7_n128 ) , .A1( u2_u3_u7_n129 ) , .ZN( u2_u3_u7_n141 ) , .A4( u2_u3_u7_n147 ) );
  INV_X1 u2_u3_u7_U4 (.A( u2_u3_u7_n111 ) , .ZN( u2_u3_u7_n170 ) );
  AOI21_X1 u2_u3_u7_U40 (.A( u2_u3_u7_n137 ) , .B1( u2_u3_u7_n138 ) , .ZN( u2_u3_u7_n139 ) , .B2( u2_u3_u7_n146 ) );
  OAI22_X1 u2_u3_u7_U41 (.B1( u2_u3_u7_n136 ) , .ZN( u2_u3_u7_n140 ) , .A1( u2_u3_u7_n153 ) , .B2( u2_u3_u7_n162 ) , .A2( u2_u3_u7_n164 ) );
  AOI21_X1 u2_u3_u7_U42 (.ZN( u2_u3_u7_n123 ) , .B1( u2_u3_u7_n165 ) , .B2( u2_u3_u7_n177 ) , .A( u2_u3_u7_n97 ) );
  AOI21_X1 u2_u3_u7_U43 (.B2( u2_u3_u7_n113 ) , .B1( u2_u3_u7_n124 ) , .A( u2_u3_u7_n125 ) , .ZN( u2_u3_u7_n97 ) );
  INV_X1 u2_u3_u7_U44 (.A( u2_u3_u7_n125 ) , .ZN( u2_u3_u7_n161 ) );
  INV_X1 u2_u3_u7_U45 (.A( u2_u3_u7_n152 ) , .ZN( u2_u3_u7_n162 ) );
  AOI22_X1 u2_u3_u7_U46 (.A2( u2_u3_u7_n114 ) , .ZN( u2_u3_u7_n119 ) , .B1( u2_u3_u7_n130 ) , .A1( u2_u3_u7_n156 ) , .B2( u2_u3_u7_n165 ) );
  NAND2_X1 u2_u3_u7_U47 (.A2( u2_u3_u7_n112 ) , .ZN( u2_u3_u7_n114 ) , .A1( u2_u3_u7_n175 ) );
  AND2_X1 u2_u3_u7_U48 (.ZN( u2_u3_u7_n145 ) , .A2( u2_u3_u7_n98 ) , .A1( u2_u3_u7_n99 ) );
  NOR2_X1 u2_u3_u7_U49 (.ZN( u2_u3_u7_n137 ) , .A1( u2_u3_u7_n150 ) , .A2( u2_u3_u7_n161 ) );
  INV_X1 u2_u3_u7_U5 (.A( u2_u3_u7_n149 ) , .ZN( u2_u3_u7_n175 ) );
  AOI21_X1 u2_u3_u7_U50 (.ZN( u2_u3_u7_n105 ) , .B2( u2_u3_u7_n110 ) , .A( u2_u3_u7_n125 ) , .B1( u2_u3_u7_n147 ) );
  NAND2_X1 u2_u3_u7_U51 (.ZN( u2_u3_u7_n146 ) , .A1( u2_u3_u7_n95 ) , .A2( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U52 (.A2( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n147 ) , .A1( u2_u3_u7_n93 ) );
  NAND2_X1 u2_u3_u7_U53 (.A1( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n127 ) , .A2( u2_u3_u7_n99 ) );
  OR2_X1 u2_u3_u7_U54 (.ZN( u2_u3_u7_n126 ) , .A2( u2_u3_u7_n152 ) , .A1( u2_u3_u7_n156 ) );
  NAND2_X1 u2_u3_u7_U55 (.A2( u2_u3_u7_n102 ) , .A1( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n133 ) );
  NAND2_X1 u2_u3_u7_U56 (.ZN( u2_u3_u7_n112 ) , .A2( u2_u3_u7_n96 ) , .A1( u2_u3_u7_n99 ) );
  NAND2_X1 u2_u3_u7_U57 (.A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n128 ) , .A1( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U58 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n113 ) , .A2( u2_u3_u7_n93 ) );
  NAND2_X1 u2_u3_u7_U59 (.A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n124 ) , .A1( u2_u3_u7_n96 ) );
  INV_X1 u2_u3_u7_U6 (.A( u2_u3_u7_n154 ) , .ZN( u2_u3_u7_n178 ) );
  NAND2_X1 u2_u3_u7_U60 (.ZN( u2_u3_u7_n110 ) , .A1( u2_u3_u7_n95 ) , .A2( u2_u3_u7_n96 ) );
  INV_X1 u2_u3_u7_U61 (.A( u2_u3_u7_n150 ) , .ZN( u2_u3_u7_n164 ) );
  AND2_X1 u2_u3_u7_U62 (.ZN( u2_u3_u7_n134 ) , .A1( u2_u3_u7_n93 ) , .A2( u2_u3_u7_n98 ) );
  NAND2_X1 u2_u3_u7_U63 (.A1( u2_u3_u7_n100 ) , .A2( u2_u3_u7_n102 ) , .ZN( u2_u3_u7_n129 ) );
  NAND2_X1 u2_u3_u7_U64 (.A2( u2_u3_u7_n103 ) , .ZN( u2_u3_u7_n131 ) , .A1( u2_u3_u7_n95 ) );
  NAND2_X1 u2_u3_u7_U65 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n138 ) , .A2( u2_u3_u7_n99 ) );
  NAND2_X1 u2_u3_u7_U66 (.ZN( u2_u3_u7_n132 ) , .A1( u2_u3_u7_n93 ) , .A2( u2_u3_u7_n96 ) );
  NAND2_X1 u2_u3_u7_U67 (.A1( u2_u3_u7_n100 ) , .ZN( u2_u3_u7_n148 ) , .A2( u2_u3_u7_n95 ) );
  NOR2_X1 u2_u3_u7_U68 (.A2( u2_u3_X_47 ) , .ZN( u2_u3_u7_n150 ) , .A1( u2_u3_u7_n163 ) );
  NOR2_X1 u2_u3_u7_U69 (.A2( u2_u3_X_43 ) , .A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n103 ) );
  AOI211_X1 u2_u3_u7_U7 (.ZN( u2_u3_u7_n116 ) , .A( u2_u3_u7_n155 ) , .C1( u2_u3_u7_n161 ) , .C2( u2_u3_u7_n171 ) , .B( u2_u3_u7_n94 ) );
  NOR2_X1 u2_u3_u7_U70 (.A2( u2_u3_X_48 ) , .A1( u2_u3_u7_n166 ) , .ZN( u2_u3_u7_n95 ) );
  NOR2_X1 u2_u3_u7_U71 (.A2( u2_u3_X_45 ) , .A1( u2_u3_X_48 ) , .ZN( u2_u3_u7_n99 ) );
  NOR2_X1 u2_u3_u7_U72 (.A2( u2_u3_X_44 ) , .A1( u2_u3_u7_n167 ) , .ZN( u2_u3_u7_n98 ) );
  NOR2_X1 u2_u3_u7_U73 (.A2( u2_u3_X_46 ) , .A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n152 ) );
  AND2_X1 u2_u3_u7_U74 (.A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n156 ) , .A2( u2_u3_u7_n163 ) );
  NAND2_X1 u2_u3_u7_U75 (.A2( u2_u3_X_46 ) , .A1( u2_u3_X_47 ) , .ZN( u2_u3_u7_n125 ) );
  AND2_X1 u2_u3_u7_U76 (.A2( u2_u3_X_45 ) , .A1( u2_u3_X_48 ) , .ZN( u2_u3_u7_n102 ) );
  AND2_X1 u2_u3_u7_U77 (.A2( u2_u3_X_43 ) , .A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n96 ) );
  AND2_X1 u2_u3_u7_U78 (.A1( u2_u3_X_44 ) , .ZN( u2_u3_u7_n100 ) , .A2( u2_u3_u7_n167 ) );
  AND2_X1 u2_u3_u7_U79 (.A1( u2_u3_X_48 ) , .A2( u2_u3_u7_n166 ) , .ZN( u2_u3_u7_n93 ) );
  OAI222_X1 u2_u3_u7_U8 (.C2( u2_u3_u7_n101 ) , .B2( u2_u3_u7_n111 ) , .A1( u2_u3_u7_n113 ) , .C1( u2_u3_u7_n146 ) , .A2( u2_u3_u7_n162 ) , .B1( u2_u3_u7_n164 ) , .ZN( u2_u3_u7_n94 ) );
  INV_X1 u2_u3_u7_U80 (.A( u2_u3_X_46 ) , .ZN( u2_u3_u7_n163 ) );
  INV_X1 u2_u3_u7_U81 (.A( u2_u3_X_43 ) , .ZN( u2_u3_u7_n167 ) );
  INV_X1 u2_u3_u7_U82 (.A( u2_u3_X_45 ) , .ZN( u2_u3_u7_n166 ) );
  NAND4_X1 u2_u3_u7_U83 (.ZN( u2_out3_5 ) , .A4( u2_u3_u7_n108 ) , .A3( u2_u3_u7_n109 ) , .A1( u2_u3_u7_n116 ) , .A2( u2_u3_u7_n123 ) );
  AOI22_X1 u2_u3_u7_U84 (.ZN( u2_u3_u7_n109 ) , .A2( u2_u3_u7_n126 ) , .B2( u2_u3_u7_n145 ) , .B1( u2_u3_u7_n156 ) , .A1( u2_u3_u7_n171 ) );
  NOR4_X1 u2_u3_u7_U85 (.A4( u2_u3_u7_n104 ) , .A3( u2_u3_u7_n105 ) , .A2( u2_u3_u7_n106 ) , .A1( u2_u3_u7_n107 ) , .ZN( u2_u3_u7_n108 ) );
  NAND4_X1 u2_u3_u7_U86 (.ZN( u2_out3_27 ) , .A4( u2_u3_u7_n118 ) , .A3( u2_u3_u7_n119 ) , .A2( u2_u3_u7_n120 ) , .A1( u2_u3_u7_n121 ) );
  OAI21_X1 u2_u3_u7_U87 (.ZN( u2_u3_u7_n121 ) , .B2( u2_u3_u7_n145 ) , .A( u2_u3_u7_n150 ) , .B1( u2_u3_u7_n174 ) );
  OAI21_X1 u2_u3_u7_U88 (.ZN( u2_u3_u7_n120 ) , .A( u2_u3_u7_n161 ) , .B2( u2_u3_u7_n170 ) , .B1( u2_u3_u7_n179 ) );
  NAND4_X1 u2_u3_u7_U89 (.ZN( u2_out3_21 ) , .A4( u2_u3_u7_n157 ) , .A3( u2_u3_u7_n158 ) , .A2( u2_u3_u7_n159 ) , .A1( u2_u3_u7_n160 ) );
  OAI221_X1 u2_u3_u7_U9 (.C1( u2_u3_u7_n101 ) , .C2( u2_u3_u7_n147 ) , .ZN( u2_u3_u7_n155 ) , .B2( u2_u3_u7_n162 ) , .A( u2_u3_u7_n91 ) , .B1( u2_u3_u7_n92 ) );
  OAI21_X1 u2_u3_u7_U90 (.B1( u2_u3_u7_n145 ) , .ZN( u2_u3_u7_n160 ) , .A( u2_u3_u7_n161 ) , .B2( u2_u3_u7_n177 ) );
  AOI22_X1 u2_u3_u7_U91 (.B2( u2_u3_u7_n149 ) , .B1( u2_u3_u7_n150 ) , .A2( u2_u3_u7_n151 ) , .A1( u2_u3_u7_n152 ) , .ZN( u2_u3_u7_n158 ) );
  NAND4_X1 u2_u3_u7_U92 (.ZN( u2_out3_15 ) , .A4( u2_u3_u7_n142 ) , .A3( u2_u3_u7_n143 ) , .A2( u2_u3_u7_n144 ) , .A1( u2_u3_u7_n178 ) );
  OR2_X1 u2_u3_u7_U93 (.A2( u2_u3_u7_n125 ) , .A1( u2_u3_u7_n129 ) , .ZN( u2_u3_u7_n144 ) );
  AOI22_X1 u2_u3_u7_U94 (.A2( u2_u3_u7_n126 ) , .ZN( u2_u3_u7_n143 ) , .B2( u2_u3_u7_n165 ) , .B1( u2_u3_u7_n173 ) , .A1( u2_u3_u7_n174 ) );
  NAND3_X1 u2_u3_u7_U95 (.A3( u2_u3_u7_n146 ) , .A2( u2_u3_u7_n147 ) , .A1( u2_u3_u7_n148 ) , .ZN( u2_u3_u7_n151 ) );
  NAND3_X1 u2_u3_u7_U96 (.A3( u2_u3_u7_n131 ) , .A2( u2_u3_u7_n132 ) , .A1( u2_u3_u7_n133 ) , .ZN( u2_u3_u7_n135 ) );
  XOR2_X1 u2_u4_U13 (.B( u2_K5_42 ) , .A( u2_R3_29 ) , .Z( u2_u4_X_42 ) );
  XOR2_X1 u2_u4_U14 (.B( u2_K5_41 ) , .A( u2_R3_28 ) , .Z( u2_u4_X_41 ) );
  XOR2_X1 u2_u4_U15 (.B( u2_K5_40 ) , .A( u2_R3_27 ) , .Z( u2_u4_X_40 ) );
  XOR2_X1 u2_u4_U17 (.B( u2_K5_39 ) , .A( u2_R3_26 ) , .Z( u2_u4_X_39 ) );
  XOR2_X1 u2_u4_U18 (.B( u2_K5_38 ) , .A( u2_R3_25 ) , .Z( u2_u4_X_38 ) );
  XOR2_X1 u2_u4_U19 (.B( u2_K5_37 ) , .A( u2_R3_24 ) , .Z( u2_u4_X_37 ) );
  XOR2_X1 u2_u4_U20 (.B( u2_K5_36 ) , .A( u2_R3_25 ) , .Z( u2_u4_X_36 ) );
  XOR2_X1 u2_u4_U21 (.B( u2_K5_35 ) , .A( u2_R3_24 ) , .Z( u2_u4_X_35 ) );
  XOR2_X1 u2_u4_U22 (.B( u2_K5_34 ) , .A( u2_R3_23 ) , .Z( u2_u4_X_34 ) );
  XOR2_X1 u2_u4_U23 (.B( u2_K5_33 ) , .A( u2_R3_22 ) , .Z( u2_u4_X_33 ) );
  XOR2_X1 u2_u4_U24 (.B( u2_K5_32 ) , .A( u2_R3_21 ) , .Z( u2_u4_X_32 ) );
  XOR2_X1 u2_u4_U25 (.B( u2_K5_31 ) , .A( u2_R3_20 ) , .Z( u2_u4_X_31 ) );
  XOR2_X1 u2_u4_U26 (.B( u2_K5_30 ) , .A( u2_R3_21 ) , .Z( u2_u4_X_30 ) );
  XOR2_X1 u2_u4_U28 (.B( u2_K5_29 ) , .A( u2_R3_20 ) , .Z( u2_u4_X_29 ) );
  XOR2_X1 u2_u4_U29 (.B( u2_K5_28 ) , .A( u2_R3_19 ) , .Z( u2_u4_X_28 ) );
  XOR2_X1 u2_u4_U30 (.B( u2_K5_27 ) , .A( u2_R3_18 ) , .Z( u2_u4_X_27 ) );
  XOR2_X1 u2_u4_U31 (.B( u2_K5_26 ) , .A( u2_R3_17 ) , .Z( u2_u4_X_26 ) );
  XOR2_X1 u2_u4_U32 (.B( u2_K5_25 ) , .A( u2_R3_16 ) , .Z( u2_u4_X_25 ) );
  OAI22_X1 u2_u4_u4_U10 (.B2( u2_u4_u4_n135 ) , .ZN( u2_u4_u4_n137 ) , .B1( u2_u4_u4_n153 ) , .A1( u2_u4_u4_n155 ) , .A2( u2_u4_u4_n171 ) );
  AND3_X1 u2_u4_u4_U11 (.A2( u2_u4_u4_n134 ) , .ZN( u2_u4_u4_n135 ) , .A3( u2_u4_u4_n145 ) , .A1( u2_u4_u4_n157 ) );
  NAND2_X1 u2_u4_u4_U12 (.ZN( u2_u4_u4_n132 ) , .A2( u2_u4_u4_n170 ) , .A1( u2_u4_u4_n173 ) );
  AOI21_X1 u2_u4_u4_U13 (.B2( u2_u4_u4_n160 ) , .B1( u2_u4_u4_n161 ) , .ZN( u2_u4_u4_n162 ) , .A( u2_u4_u4_n170 ) );
  AOI21_X1 u2_u4_u4_U14 (.ZN( u2_u4_u4_n107 ) , .B2( u2_u4_u4_n143 ) , .A( u2_u4_u4_n174 ) , .B1( u2_u4_u4_n184 ) );
  AOI21_X1 u2_u4_u4_U15 (.B2( u2_u4_u4_n158 ) , .B1( u2_u4_u4_n159 ) , .ZN( u2_u4_u4_n163 ) , .A( u2_u4_u4_n174 ) );
  AOI21_X1 u2_u4_u4_U16 (.A( u2_u4_u4_n153 ) , .B2( u2_u4_u4_n154 ) , .B1( u2_u4_u4_n155 ) , .ZN( u2_u4_u4_n165 ) );
  AOI21_X1 u2_u4_u4_U17 (.A( u2_u4_u4_n156 ) , .B2( u2_u4_u4_n157 ) , .ZN( u2_u4_u4_n164 ) , .B1( u2_u4_u4_n184 ) );
  INV_X1 u2_u4_u4_U18 (.A( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n170 ) );
  AND2_X1 u2_u4_u4_U19 (.A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n155 ) , .A1( u2_u4_u4_n160 ) );
  INV_X1 u2_u4_u4_U20 (.A( u2_u4_u4_n156 ) , .ZN( u2_u4_u4_n175 ) );
  NAND2_X1 u2_u4_u4_U21 (.A2( u2_u4_u4_n118 ) , .ZN( u2_u4_u4_n131 ) , .A1( u2_u4_u4_n147 ) );
  NAND2_X1 u2_u4_u4_U22 (.A1( u2_u4_u4_n119 ) , .A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n130 ) );
  NAND2_X1 u2_u4_u4_U23 (.ZN( u2_u4_u4_n117 ) , .A2( u2_u4_u4_n118 ) , .A1( u2_u4_u4_n148 ) );
  NAND2_X1 u2_u4_u4_U24 (.ZN( u2_u4_u4_n129 ) , .A1( u2_u4_u4_n134 ) , .A2( u2_u4_u4_n148 ) );
  AND3_X1 u2_u4_u4_U25 (.A1( u2_u4_u4_n119 ) , .A2( u2_u4_u4_n143 ) , .A3( u2_u4_u4_n154 ) , .ZN( u2_u4_u4_n161 ) );
  AND2_X1 u2_u4_u4_U26 (.A1( u2_u4_u4_n145 ) , .A2( u2_u4_u4_n147 ) , .ZN( u2_u4_u4_n159 ) );
  OR3_X1 u2_u4_u4_U27 (.A3( u2_u4_u4_n114 ) , .A2( u2_u4_u4_n115 ) , .A1( u2_u4_u4_n116 ) , .ZN( u2_u4_u4_n136 ) );
  AOI21_X1 u2_u4_u4_U28 (.A( u2_u4_u4_n113 ) , .ZN( u2_u4_u4_n116 ) , .B2( u2_u4_u4_n173 ) , .B1( u2_u4_u4_n174 ) );
  AOI21_X1 u2_u4_u4_U29 (.ZN( u2_u4_u4_n115 ) , .B2( u2_u4_u4_n145 ) , .B1( u2_u4_u4_n146 ) , .A( u2_u4_u4_n156 ) );
  NOR2_X1 u2_u4_u4_U3 (.ZN( u2_u4_u4_n121 ) , .A1( u2_u4_u4_n181 ) , .A2( u2_u4_u4_n182 ) );
  OAI22_X1 u2_u4_u4_U30 (.ZN( u2_u4_u4_n114 ) , .A2( u2_u4_u4_n121 ) , .B1( u2_u4_u4_n160 ) , .B2( u2_u4_u4_n170 ) , .A1( u2_u4_u4_n171 ) );
  INV_X1 u2_u4_u4_U31 (.A( u2_u4_u4_n158 ) , .ZN( u2_u4_u4_n182 ) );
  INV_X1 u2_u4_u4_U32 (.ZN( u2_u4_u4_n181 ) , .A( u2_u4_u4_n96 ) );
  INV_X1 u2_u4_u4_U33 (.A( u2_u4_u4_n144 ) , .ZN( u2_u4_u4_n179 ) );
  INV_X1 u2_u4_u4_U34 (.A( u2_u4_u4_n157 ) , .ZN( u2_u4_u4_n178 ) );
  NAND2_X1 u2_u4_u4_U35 (.A2( u2_u4_u4_n154 ) , .A1( u2_u4_u4_n96 ) , .ZN( u2_u4_u4_n97 ) );
  INV_X1 u2_u4_u4_U36 (.ZN( u2_u4_u4_n186 ) , .A( u2_u4_u4_n95 ) );
  OAI221_X1 u2_u4_u4_U37 (.C1( u2_u4_u4_n134 ) , .B1( u2_u4_u4_n158 ) , .B2( u2_u4_u4_n171 ) , .C2( u2_u4_u4_n173 ) , .A( u2_u4_u4_n94 ) , .ZN( u2_u4_u4_n95 ) );
  AOI222_X1 u2_u4_u4_U38 (.B2( u2_u4_u4_n132 ) , .A1( u2_u4_u4_n138 ) , .C2( u2_u4_u4_n175 ) , .A2( u2_u4_u4_n179 ) , .C1( u2_u4_u4_n181 ) , .B1( u2_u4_u4_n185 ) , .ZN( u2_u4_u4_n94 ) );
  INV_X1 u2_u4_u4_U39 (.A( u2_u4_u4_n113 ) , .ZN( u2_u4_u4_n185 ) );
  INV_X1 u2_u4_u4_U4 (.A( u2_u4_u4_n117 ) , .ZN( u2_u4_u4_n184 ) );
  INV_X1 u2_u4_u4_U40 (.A( u2_u4_u4_n143 ) , .ZN( u2_u4_u4_n183 ) );
  NOR2_X1 u2_u4_u4_U41 (.ZN( u2_u4_u4_n138 ) , .A1( u2_u4_u4_n168 ) , .A2( u2_u4_u4_n169 ) );
  NOR2_X1 u2_u4_u4_U42 (.A1( u2_u4_u4_n150 ) , .A2( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n153 ) );
  NOR2_X1 u2_u4_u4_U43 (.A2( u2_u4_u4_n128 ) , .A1( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n156 ) );
  AOI22_X1 u2_u4_u4_U44 (.B2( u2_u4_u4_n122 ) , .A1( u2_u4_u4_n123 ) , .ZN( u2_u4_u4_n124 ) , .B1( u2_u4_u4_n128 ) , .A2( u2_u4_u4_n172 ) );
  INV_X1 u2_u4_u4_U45 (.A( u2_u4_u4_n153 ) , .ZN( u2_u4_u4_n172 ) );
  NAND2_X1 u2_u4_u4_U46 (.A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n123 ) , .A1( u2_u4_u4_n161 ) );
  AOI22_X1 u2_u4_u4_U47 (.B2( u2_u4_u4_n132 ) , .A2( u2_u4_u4_n133 ) , .ZN( u2_u4_u4_n140 ) , .A1( u2_u4_u4_n150 ) , .B1( u2_u4_u4_n179 ) );
  NAND2_X1 u2_u4_u4_U48 (.ZN( u2_u4_u4_n133 ) , .A2( u2_u4_u4_n146 ) , .A1( u2_u4_u4_n154 ) );
  NAND2_X1 u2_u4_u4_U49 (.A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n154 ) , .A2( u2_u4_u4_n98 ) );
  NOR4_X1 u2_u4_u4_U5 (.A4( u2_u4_u4_n106 ) , .A3( u2_u4_u4_n107 ) , .A2( u2_u4_u4_n108 ) , .A1( u2_u4_u4_n109 ) , .ZN( u2_u4_u4_n110 ) );
  NAND2_X1 u2_u4_u4_U50 (.A1( u2_u4_u4_n101 ) , .ZN( u2_u4_u4_n158 ) , .A2( u2_u4_u4_n99 ) );
  AOI21_X1 u2_u4_u4_U51 (.ZN( u2_u4_u4_n127 ) , .A( u2_u4_u4_n136 ) , .B2( u2_u4_u4_n150 ) , .B1( u2_u4_u4_n180 ) );
  INV_X1 u2_u4_u4_U52 (.A( u2_u4_u4_n160 ) , .ZN( u2_u4_u4_n180 ) );
  NAND2_X1 u2_u4_u4_U53 (.A2( u2_u4_u4_n104 ) , .A1( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n146 ) );
  NAND2_X1 u2_u4_u4_U54 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n160 ) );
  NAND2_X1 u2_u4_u4_U55 (.ZN( u2_u4_u4_n134 ) , .A1( u2_u4_u4_n98 ) , .A2( u2_u4_u4_n99 ) );
  NAND2_X1 u2_u4_u4_U56 (.A1( u2_u4_u4_n103 ) , .A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n143 ) );
  NAND2_X1 u2_u4_u4_U57 (.A2( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n145 ) , .A1( u2_u4_u4_n98 ) );
  NAND2_X1 u2_u4_u4_U58 (.A1( u2_u4_u4_n100 ) , .A2( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n120 ) );
  NAND2_X1 u2_u4_u4_U59 (.A1( u2_u4_u4_n102 ) , .A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n148 ) );
  AOI21_X1 u2_u4_u4_U6 (.ZN( u2_u4_u4_n106 ) , .B2( u2_u4_u4_n146 ) , .B1( u2_u4_u4_n158 ) , .A( u2_u4_u4_n170 ) );
  NAND2_X1 u2_u4_u4_U60 (.A2( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n157 ) );
  INV_X1 u2_u4_u4_U61 (.A( u2_u4_u4_n150 ) , .ZN( u2_u4_u4_n173 ) );
  INV_X1 u2_u4_u4_U62 (.A( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n171 ) );
  NAND2_X1 u2_u4_u4_U63 (.A1( u2_u4_u4_n100 ) , .ZN( u2_u4_u4_n118 ) , .A2( u2_u4_u4_n99 ) );
  NAND2_X1 u2_u4_u4_U64 (.A2( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n144 ) );
  NAND2_X1 u2_u4_u4_U65 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n96 ) );
  INV_X1 u2_u4_u4_U66 (.A( u2_u4_u4_n128 ) , .ZN( u2_u4_u4_n174 ) );
  NAND2_X1 u2_u4_u4_U67 (.A2( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n119 ) , .A1( u2_u4_u4_n98 ) );
  NAND2_X1 u2_u4_u4_U68 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n147 ) );
  NAND2_X1 u2_u4_u4_U69 (.A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n113 ) , .A1( u2_u4_u4_n99 ) );
  AOI21_X1 u2_u4_u4_U7 (.ZN( u2_u4_u4_n108 ) , .B2( u2_u4_u4_n134 ) , .B1( u2_u4_u4_n155 ) , .A( u2_u4_u4_n156 ) );
  NOR2_X1 u2_u4_u4_U70 (.A2( u2_u4_X_28 ) , .ZN( u2_u4_u4_n150 ) , .A1( u2_u4_u4_n168 ) );
  NOR2_X1 u2_u4_u4_U71 (.A2( u2_u4_X_29 ) , .ZN( u2_u4_u4_n152 ) , .A1( u2_u4_u4_n169 ) );
  NOR2_X1 u2_u4_u4_U72 (.A2( u2_u4_X_30 ) , .ZN( u2_u4_u4_n105 ) , .A1( u2_u4_u4_n176 ) );
  NOR2_X1 u2_u4_u4_U73 (.A2( u2_u4_X_26 ) , .ZN( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n177 ) );
  NOR2_X1 u2_u4_u4_U74 (.A2( u2_u4_X_28 ) , .A1( u2_u4_X_29 ) , .ZN( u2_u4_u4_n128 ) );
  NOR2_X1 u2_u4_u4_U75 (.A2( u2_u4_X_27 ) , .A1( u2_u4_X_30 ) , .ZN( u2_u4_u4_n102 ) );
  NOR2_X1 u2_u4_u4_U76 (.A2( u2_u4_X_25 ) , .A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n98 ) );
  AND2_X1 u2_u4_u4_U77 (.A2( u2_u4_X_25 ) , .A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n104 ) );
  AND2_X1 u2_u4_u4_U78 (.A1( u2_u4_X_30 ) , .A2( u2_u4_u4_n176 ) , .ZN( u2_u4_u4_n99 ) );
  AND2_X1 u2_u4_u4_U79 (.A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n101 ) , .A2( u2_u4_u4_n177 ) );
  AOI21_X1 u2_u4_u4_U8 (.ZN( u2_u4_u4_n109 ) , .A( u2_u4_u4_n153 ) , .B1( u2_u4_u4_n159 ) , .B2( u2_u4_u4_n184 ) );
  AND2_X1 u2_u4_u4_U80 (.A1( u2_u4_X_27 ) , .A2( u2_u4_X_30 ) , .ZN( u2_u4_u4_n103 ) );
  INV_X1 u2_u4_u4_U81 (.A( u2_u4_X_28 ) , .ZN( u2_u4_u4_n169 ) );
  INV_X1 u2_u4_u4_U82 (.A( u2_u4_X_29 ) , .ZN( u2_u4_u4_n168 ) );
  INV_X1 u2_u4_u4_U83 (.A( u2_u4_X_25 ) , .ZN( u2_u4_u4_n177 ) );
  INV_X1 u2_u4_u4_U84 (.A( u2_u4_X_27 ) , .ZN( u2_u4_u4_n176 ) );
  NAND4_X1 u2_u4_u4_U85 (.ZN( u2_out4_25 ) , .A4( u2_u4_u4_n139 ) , .A3( u2_u4_u4_n140 ) , .A2( u2_u4_u4_n141 ) , .A1( u2_u4_u4_n142 ) );
  OAI21_X1 u2_u4_u4_U86 (.B2( u2_u4_u4_n131 ) , .ZN( u2_u4_u4_n141 ) , .A( u2_u4_u4_n175 ) , .B1( u2_u4_u4_n183 ) );
  OAI21_X1 u2_u4_u4_U87 (.A( u2_u4_u4_n128 ) , .B2( u2_u4_u4_n129 ) , .B1( u2_u4_u4_n130 ) , .ZN( u2_u4_u4_n142 ) );
  NAND4_X1 u2_u4_u4_U88 (.ZN( u2_out4_14 ) , .A4( u2_u4_u4_n124 ) , .A3( u2_u4_u4_n125 ) , .A2( u2_u4_u4_n126 ) , .A1( u2_u4_u4_n127 ) );
  AOI22_X1 u2_u4_u4_U89 (.B2( u2_u4_u4_n117 ) , .ZN( u2_u4_u4_n126 ) , .A1( u2_u4_u4_n129 ) , .B1( u2_u4_u4_n152 ) , .A2( u2_u4_u4_n175 ) );
  AOI211_X1 u2_u4_u4_U9 (.B( u2_u4_u4_n136 ) , .A( u2_u4_u4_n137 ) , .C2( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n139 ) , .C1( u2_u4_u4_n182 ) );
  AOI22_X1 u2_u4_u4_U90 (.ZN( u2_u4_u4_n125 ) , .B2( u2_u4_u4_n131 ) , .A2( u2_u4_u4_n132 ) , .B1( u2_u4_u4_n138 ) , .A1( u2_u4_u4_n178 ) );
  NAND4_X1 u2_u4_u4_U91 (.ZN( u2_out4_8 ) , .A4( u2_u4_u4_n110 ) , .A3( u2_u4_u4_n111 ) , .A2( u2_u4_u4_n112 ) , .A1( u2_u4_u4_n186 ) );
  NAND2_X1 u2_u4_u4_U92 (.ZN( u2_u4_u4_n112 ) , .A2( u2_u4_u4_n130 ) , .A1( u2_u4_u4_n150 ) );
  AOI22_X1 u2_u4_u4_U93 (.ZN( u2_u4_u4_n111 ) , .B2( u2_u4_u4_n132 ) , .A1( u2_u4_u4_n152 ) , .B1( u2_u4_u4_n178 ) , .A2( u2_u4_u4_n97 ) );
  AOI22_X1 u2_u4_u4_U94 (.B2( u2_u4_u4_n149 ) , .B1( u2_u4_u4_n150 ) , .A2( u2_u4_u4_n151 ) , .A1( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n167 ) );
  NOR4_X1 u2_u4_u4_U95 (.A4( u2_u4_u4_n162 ) , .A3( u2_u4_u4_n163 ) , .A2( u2_u4_u4_n164 ) , .A1( u2_u4_u4_n165 ) , .ZN( u2_u4_u4_n166 ) );
  NAND3_X1 u2_u4_u4_U96 (.ZN( u2_out4_3 ) , .A3( u2_u4_u4_n166 ) , .A1( u2_u4_u4_n167 ) , .A2( u2_u4_u4_n186 ) );
  NAND3_X1 u2_u4_u4_U97 (.A3( u2_u4_u4_n146 ) , .A2( u2_u4_u4_n147 ) , .A1( u2_u4_u4_n148 ) , .ZN( u2_u4_u4_n149 ) );
  NAND3_X1 u2_u4_u4_U98 (.A3( u2_u4_u4_n143 ) , .A2( u2_u4_u4_n144 ) , .A1( u2_u4_u4_n145 ) , .ZN( u2_u4_u4_n151 ) );
  NAND3_X1 u2_u4_u4_U99 (.A3( u2_u4_u4_n121 ) , .ZN( u2_u4_u4_n122 ) , .A2( u2_u4_u4_n144 ) , .A1( u2_u4_u4_n154 ) );
  NOR2_X1 u2_u4_u5_U10 (.ZN( u2_u4_u5_n135 ) , .A1( u2_u4_u5_n173 ) , .A2( u2_u4_u5_n176 ) );
  NOR3_X1 u2_u4_u5_U100 (.A3( u2_u4_u5_n141 ) , .A1( u2_u4_u5_n142 ) , .ZN( u2_u4_u5_n143 ) , .A2( u2_u4_u5_n191 ) );
  NAND4_X1 u2_u4_u5_U101 (.ZN( u2_out4_4 ) , .A4( u2_u4_u5_n112 ) , .A2( u2_u4_u5_n113 ) , .A1( u2_u4_u5_n114 ) , .A3( u2_u4_u5_n195 ) );
  AOI211_X1 u2_u4_u5_U102 (.A( u2_u4_u5_n110 ) , .C1( u2_u4_u5_n111 ) , .ZN( u2_u4_u5_n112 ) , .B( u2_u4_u5_n118 ) , .C2( u2_u4_u5_n177 ) );
  INV_X1 u2_u4_u5_U103 (.A( u2_u4_u5_n102 ) , .ZN( u2_u4_u5_n195 ) );
  NAND3_X1 u2_u4_u5_U104 (.A2( u2_u4_u5_n154 ) , .A3( u2_u4_u5_n158 ) , .A1( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n99 ) );
  INV_X1 u2_u4_u5_U11 (.A( u2_u4_u5_n121 ) , .ZN( u2_u4_u5_n177 ) );
  NOR2_X1 u2_u4_u5_U12 (.ZN( u2_u4_u5_n160 ) , .A2( u2_u4_u5_n173 ) , .A1( u2_u4_u5_n177 ) );
  INV_X1 u2_u4_u5_U13 (.A( u2_u4_u5_n150 ) , .ZN( u2_u4_u5_n174 ) );
  AOI21_X1 u2_u4_u5_U14 (.A( u2_u4_u5_n160 ) , .B2( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n162 ) , .B1( u2_u4_u5_n192 ) );
  INV_X1 u2_u4_u5_U15 (.A( u2_u4_u5_n159 ) , .ZN( u2_u4_u5_n192 ) );
  AOI21_X1 u2_u4_u5_U16 (.A( u2_u4_u5_n156 ) , .B2( u2_u4_u5_n157 ) , .B1( u2_u4_u5_n158 ) , .ZN( u2_u4_u5_n163 ) );
  AOI21_X1 u2_u4_u5_U17 (.B2( u2_u4_u5_n139 ) , .B1( u2_u4_u5_n140 ) , .ZN( u2_u4_u5_n141 ) , .A( u2_u4_u5_n150 ) );
  OAI21_X1 u2_u4_u5_U18 (.A( u2_u4_u5_n133 ) , .B2( u2_u4_u5_n134 ) , .B1( u2_u4_u5_n135 ) , .ZN( u2_u4_u5_n142 ) );
  OAI21_X1 u2_u4_u5_U19 (.ZN( u2_u4_u5_n133 ) , .B2( u2_u4_u5_n147 ) , .A( u2_u4_u5_n173 ) , .B1( u2_u4_u5_n188 ) );
  NAND2_X1 u2_u4_u5_U20 (.A2( u2_u4_u5_n119 ) , .A1( u2_u4_u5_n123 ) , .ZN( u2_u4_u5_n137 ) );
  INV_X1 u2_u4_u5_U21 (.A( u2_u4_u5_n155 ) , .ZN( u2_u4_u5_n194 ) );
  NAND2_X1 u2_u4_u5_U22 (.A1( u2_u4_u5_n121 ) , .ZN( u2_u4_u5_n132 ) , .A2( u2_u4_u5_n172 ) );
  NAND2_X1 u2_u4_u5_U23 (.A2( u2_u4_u5_n122 ) , .ZN( u2_u4_u5_n136 ) , .A1( u2_u4_u5_n154 ) );
  NAND2_X1 u2_u4_u5_U24 (.A2( u2_u4_u5_n119 ) , .A1( u2_u4_u5_n120 ) , .ZN( u2_u4_u5_n159 ) );
  INV_X1 u2_u4_u5_U25 (.A( u2_u4_u5_n156 ) , .ZN( u2_u4_u5_n175 ) );
  INV_X1 u2_u4_u5_U26 (.A( u2_u4_u5_n158 ) , .ZN( u2_u4_u5_n188 ) );
  INV_X1 u2_u4_u5_U27 (.A( u2_u4_u5_n152 ) , .ZN( u2_u4_u5_n179 ) );
  INV_X1 u2_u4_u5_U28 (.A( u2_u4_u5_n140 ) , .ZN( u2_u4_u5_n182 ) );
  INV_X1 u2_u4_u5_U29 (.A( u2_u4_u5_n151 ) , .ZN( u2_u4_u5_n183 ) );
  NOR2_X1 u2_u4_u5_U3 (.ZN( u2_u4_u5_n134 ) , .A1( u2_u4_u5_n183 ) , .A2( u2_u4_u5_n190 ) );
  INV_X1 u2_u4_u5_U30 (.A( u2_u4_u5_n123 ) , .ZN( u2_u4_u5_n185 ) );
  INV_X1 u2_u4_u5_U31 (.A( u2_u4_u5_n161 ) , .ZN( u2_u4_u5_n184 ) );
  INV_X1 u2_u4_u5_U32 (.A( u2_u4_u5_n139 ) , .ZN( u2_u4_u5_n189 ) );
  INV_X1 u2_u4_u5_U33 (.A( u2_u4_u5_n157 ) , .ZN( u2_u4_u5_n190 ) );
  INV_X1 u2_u4_u5_U34 (.A( u2_u4_u5_n120 ) , .ZN( u2_u4_u5_n193 ) );
  NAND2_X1 u2_u4_u5_U35 (.ZN( u2_u4_u5_n111 ) , .A1( u2_u4_u5_n140 ) , .A2( u2_u4_u5_n155 ) );
  INV_X1 u2_u4_u5_U36 (.A( u2_u4_u5_n117 ) , .ZN( u2_u4_u5_n196 ) );
  OAI221_X1 u2_u4_u5_U37 (.A( u2_u4_u5_n116 ) , .ZN( u2_u4_u5_n117 ) , .B2( u2_u4_u5_n119 ) , .C1( u2_u4_u5_n153 ) , .C2( u2_u4_u5_n158 ) , .B1( u2_u4_u5_n172 ) );
  AOI222_X1 u2_u4_u5_U38 (.ZN( u2_u4_u5_n116 ) , .B2( u2_u4_u5_n145 ) , .C1( u2_u4_u5_n148 ) , .A2( u2_u4_u5_n174 ) , .C2( u2_u4_u5_n177 ) , .B1( u2_u4_u5_n187 ) , .A1( u2_u4_u5_n193 ) );
  INV_X1 u2_u4_u5_U39 (.A( u2_u4_u5_n115 ) , .ZN( u2_u4_u5_n187 ) );
  INV_X1 u2_u4_u5_U4 (.A( u2_u4_u5_n138 ) , .ZN( u2_u4_u5_n191 ) );
  NOR2_X1 u2_u4_u5_U40 (.ZN( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n170 ) , .A2( u2_u4_u5_n180 ) );
  OAI221_X1 u2_u4_u5_U41 (.A( u2_u4_u5_n101 ) , .ZN( u2_u4_u5_n102 ) , .C2( u2_u4_u5_n115 ) , .C1( u2_u4_u5_n126 ) , .B1( u2_u4_u5_n134 ) , .B2( u2_u4_u5_n160 ) );
  OAI21_X1 u2_u4_u5_U42 (.ZN( u2_u4_u5_n101 ) , .B1( u2_u4_u5_n137 ) , .A( u2_u4_u5_n146 ) , .B2( u2_u4_u5_n147 ) );
  AOI22_X1 u2_u4_u5_U43 (.B2( u2_u4_u5_n131 ) , .A2( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n169 ) , .B1( u2_u4_u5_n174 ) , .A1( u2_u4_u5_n185 ) );
  NOR2_X1 u2_u4_u5_U44 (.A1( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n150 ) , .A2( u2_u4_u5_n173 ) );
  AOI21_X1 u2_u4_u5_U45 (.A( u2_u4_u5_n118 ) , .B2( u2_u4_u5_n145 ) , .ZN( u2_u4_u5_n168 ) , .B1( u2_u4_u5_n186 ) );
  INV_X1 u2_u4_u5_U46 (.A( u2_u4_u5_n122 ) , .ZN( u2_u4_u5_n186 ) );
  NOR2_X1 u2_u4_u5_U47 (.A1( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n152 ) , .A2( u2_u4_u5_n176 ) );
  NOR2_X1 u2_u4_u5_U48 (.A1( u2_u4_u5_n115 ) , .ZN( u2_u4_u5_n118 ) , .A2( u2_u4_u5_n153 ) );
  NOR2_X1 u2_u4_u5_U49 (.A2( u2_u4_u5_n145 ) , .ZN( u2_u4_u5_n156 ) , .A1( u2_u4_u5_n174 ) );
  OAI21_X1 u2_u4_u5_U5 (.B2( u2_u4_u5_n136 ) , .B1( u2_u4_u5_n137 ) , .ZN( u2_u4_u5_n138 ) , .A( u2_u4_u5_n177 ) );
  NOR2_X1 u2_u4_u5_U50 (.ZN( u2_u4_u5_n121 ) , .A2( u2_u4_u5_n145 ) , .A1( u2_u4_u5_n176 ) );
  AOI22_X1 u2_u4_u5_U51 (.ZN( u2_u4_u5_n114 ) , .A2( u2_u4_u5_n137 ) , .A1( u2_u4_u5_n145 ) , .B2( u2_u4_u5_n175 ) , .B1( u2_u4_u5_n193 ) );
  OAI211_X1 u2_u4_u5_U52 (.B( u2_u4_u5_n124 ) , .A( u2_u4_u5_n125 ) , .C2( u2_u4_u5_n126 ) , .C1( u2_u4_u5_n127 ) , .ZN( u2_u4_u5_n128 ) );
  NOR3_X1 u2_u4_u5_U53 (.ZN( u2_u4_u5_n127 ) , .A1( u2_u4_u5_n136 ) , .A3( u2_u4_u5_n148 ) , .A2( u2_u4_u5_n182 ) );
  OAI21_X1 u2_u4_u5_U54 (.ZN( u2_u4_u5_n124 ) , .A( u2_u4_u5_n177 ) , .B2( u2_u4_u5_n183 ) , .B1( u2_u4_u5_n189 ) );
  OAI21_X1 u2_u4_u5_U55 (.ZN( u2_u4_u5_n125 ) , .A( u2_u4_u5_n174 ) , .B2( u2_u4_u5_n185 ) , .B1( u2_u4_u5_n190 ) );
  AOI21_X1 u2_u4_u5_U56 (.A( u2_u4_u5_n153 ) , .B2( u2_u4_u5_n154 ) , .B1( u2_u4_u5_n155 ) , .ZN( u2_u4_u5_n164 ) );
  AOI21_X1 u2_u4_u5_U57 (.ZN( u2_u4_u5_n110 ) , .B1( u2_u4_u5_n122 ) , .B2( u2_u4_u5_n139 ) , .A( u2_u4_u5_n153 ) );
  INV_X1 u2_u4_u5_U58 (.A( u2_u4_u5_n153 ) , .ZN( u2_u4_u5_n176 ) );
  INV_X1 u2_u4_u5_U59 (.A( u2_u4_u5_n126 ) , .ZN( u2_u4_u5_n173 ) );
  AOI222_X1 u2_u4_u5_U6 (.ZN( u2_u4_u5_n113 ) , .A1( u2_u4_u5_n131 ) , .C1( u2_u4_u5_n148 ) , .B2( u2_u4_u5_n174 ) , .C2( u2_u4_u5_n178 ) , .A2( u2_u4_u5_n179 ) , .B1( u2_u4_u5_n99 ) );
  AND2_X1 u2_u4_u5_U60 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n147 ) );
  AND2_X1 u2_u4_u5_U61 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n148 ) );
  NAND2_X1 u2_u4_u5_U62 (.A1( u2_u4_u5_n105 ) , .A2( u2_u4_u5_n106 ) , .ZN( u2_u4_u5_n158 ) );
  NAND2_X1 u2_u4_u5_U63 (.A2( u2_u4_u5_n108 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n139 ) );
  NAND2_X1 u2_u4_u5_U64 (.A1( u2_u4_u5_n106 ) , .A2( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n119 ) );
  NAND2_X1 u2_u4_u5_U65 (.A2( u2_u4_u5_n103 ) , .A1( u2_u4_u5_n105 ) , .ZN( u2_u4_u5_n140 ) );
  NAND2_X1 u2_u4_u5_U66 (.A2( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n105 ) , .ZN( u2_u4_u5_n155 ) );
  NAND2_X1 u2_u4_u5_U67 (.A2( u2_u4_u5_n106 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n122 ) );
  NAND2_X1 u2_u4_u5_U68 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n106 ) , .ZN( u2_u4_u5_n115 ) );
  NAND2_X1 u2_u4_u5_U69 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n103 ) , .ZN( u2_u4_u5_n161 ) );
  INV_X1 u2_u4_u5_U7 (.A( u2_u4_u5_n135 ) , .ZN( u2_u4_u5_n178 ) );
  NAND2_X1 u2_u4_u5_U70 (.A1( u2_u4_u5_n105 ) , .A2( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n154 ) );
  INV_X1 u2_u4_u5_U71 (.A( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n172 ) );
  NAND2_X1 u2_u4_u5_U72 (.A1( u2_u4_u5_n103 ) , .A2( u2_u4_u5_n108 ) , .ZN( u2_u4_u5_n123 ) );
  NAND2_X1 u2_u4_u5_U73 (.A2( u2_u4_u5_n103 ) , .A1( u2_u4_u5_n107 ) , .ZN( u2_u4_u5_n151 ) );
  NAND2_X1 u2_u4_u5_U74 (.A2( u2_u4_u5_n107 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n120 ) );
  NAND2_X1 u2_u4_u5_U75 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n109 ) , .ZN( u2_u4_u5_n157 ) );
  AND2_X1 u2_u4_u5_U76 (.A2( u2_u4_u5_n100 ) , .A1( u2_u4_u5_n104 ) , .ZN( u2_u4_u5_n131 ) );
  NOR2_X1 u2_u4_u5_U77 (.A2( u2_u4_X_34 ) , .A1( u2_u4_X_35 ) , .ZN( u2_u4_u5_n145 ) );
  NOR2_X1 u2_u4_u5_U78 (.A2( u2_u4_X_34 ) , .ZN( u2_u4_u5_n146 ) , .A1( u2_u4_u5_n171 ) );
  NOR2_X1 u2_u4_u5_U79 (.A2( u2_u4_X_31 ) , .A1( u2_u4_X_32 ) , .ZN( u2_u4_u5_n103 ) );
  OAI22_X1 u2_u4_u5_U8 (.B2( u2_u4_u5_n149 ) , .B1( u2_u4_u5_n150 ) , .A2( u2_u4_u5_n151 ) , .A1( u2_u4_u5_n152 ) , .ZN( u2_u4_u5_n165 ) );
  NOR2_X1 u2_u4_u5_U80 (.A2( u2_u4_X_36 ) , .ZN( u2_u4_u5_n105 ) , .A1( u2_u4_u5_n180 ) );
  NOR2_X1 u2_u4_u5_U81 (.A2( u2_u4_X_33 ) , .ZN( u2_u4_u5_n108 ) , .A1( u2_u4_u5_n170 ) );
  NOR2_X1 u2_u4_u5_U82 (.A2( u2_u4_X_33 ) , .A1( u2_u4_X_36 ) , .ZN( u2_u4_u5_n107 ) );
  NOR2_X1 u2_u4_u5_U83 (.A2( u2_u4_X_31 ) , .ZN( u2_u4_u5_n104 ) , .A1( u2_u4_u5_n181 ) );
  NAND2_X1 u2_u4_u5_U84 (.A2( u2_u4_X_34 ) , .A1( u2_u4_X_35 ) , .ZN( u2_u4_u5_n153 ) );
  NAND2_X1 u2_u4_u5_U85 (.A1( u2_u4_X_34 ) , .ZN( u2_u4_u5_n126 ) , .A2( u2_u4_u5_n171 ) );
  AND2_X1 u2_u4_u5_U86 (.A1( u2_u4_X_31 ) , .A2( u2_u4_X_32 ) , .ZN( u2_u4_u5_n106 ) );
  AND2_X1 u2_u4_u5_U87 (.A1( u2_u4_X_31 ) , .ZN( u2_u4_u5_n109 ) , .A2( u2_u4_u5_n181 ) );
  INV_X1 u2_u4_u5_U88 (.A( u2_u4_X_33 ) , .ZN( u2_u4_u5_n180 ) );
  INV_X1 u2_u4_u5_U89 (.A( u2_u4_X_35 ) , .ZN( u2_u4_u5_n171 ) );
  NOR3_X1 u2_u4_u5_U9 (.A2( u2_u4_u5_n147 ) , .A1( u2_u4_u5_n148 ) , .ZN( u2_u4_u5_n149 ) , .A3( u2_u4_u5_n194 ) );
  INV_X1 u2_u4_u5_U90 (.A( u2_u4_X_36 ) , .ZN( u2_u4_u5_n170 ) );
  INV_X1 u2_u4_u5_U91 (.A( u2_u4_X_32 ) , .ZN( u2_u4_u5_n181 ) );
  NAND4_X1 u2_u4_u5_U92 (.ZN( u2_out4_29 ) , .A4( u2_u4_u5_n129 ) , .A3( u2_u4_u5_n130 ) , .A2( u2_u4_u5_n168 ) , .A1( u2_u4_u5_n196 ) );
  AOI221_X1 u2_u4_u5_U93 (.A( u2_u4_u5_n128 ) , .ZN( u2_u4_u5_n129 ) , .C2( u2_u4_u5_n132 ) , .B2( u2_u4_u5_n159 ) , .B1( u2_u4_u5_n176 ) , .C1( u2_u4_u5_n184 ) );
  AOI222_X1 u2_u4_u5_U94 (.ZN( u2_u4_u5_n130 ) , .A2( u2_u4_u5_n146 ) , .B1( u2_u4_u5_n147 ) , .C2( u2_u4_u5_n175 ) , .B2( u2_u4_u5_n179 ) , .A1( u2_u4_u5_n188 ) , .C1( u2_u4_u5_n194 ) );
  NAND4_X1 u2_u4_u5_U95 (.ZN( u2_out4_19 ) , .A4( u2_u4_u5_n166 ) , .A3( u2_u4_u5_n167 ) , .A2( u2_u4_u5_n168 ) , .A1( u2_u4_u5_n169 ) );
  AOI22_X1 u2_u4_u5_U96 (.B2( u2_u4_u5_n145 ) , .A2( u2_u4_u5_n146 ) , .ZN( u2_u4_u5_n167 ) , .B1( u2_u4_u5_n182 ) , .A1( u2_u4_u5_n189 ) );
  NOR4_X1 u2_u4_u5_U97 (.A4( u2_u4_u5_n162 ) , .A3( u2_u4_u5_n163 ) , .A2( u2_u4_u5_n164 ) , .A1( u2_u4_u5_n165 ) , .ZN( u2_u4_u5_n166 ) );
  NAND4_X1 u2_u4_u5_U98 (.ZN( u2_out4_11 ) , .A4( u2_u4_u5_n143 ) , .A3( u2_u4_u5_n144 ) , .A2( u2_u4_u5_n169 ) , .A1( u2_u4_u5_n196 ) );
  AOI22_X1 u2_u4_u5_U99 (.A2( u2_u4_u5_n132 ) , .ZN( u2_u4_u5_n144 ) , .B2( u2_u4_u5_n145 ) , .B1( u2_u4_u5_n184 ) , .A1( u2_u4_u5_n194 ) );
  AOI22_X1 u2_u4_u6_U10 (.A2( u2_u4_u6_n151 ) , .B2( u2_u4_u6_n161 ) , .A1( u2_u4_u6_n167 ) , .B1( u2_u4_u6_n170 ) , .ZN( u2_u4_u6_n89 ) );
  AOI21_X1 u2_u4_u6_U11 (.B1( u2_u4_u6_n107 ) , .B2( u2_u4_u6_n132 ) , .A( u2_u4_u6_n158 ) , .ZN( u2_u4_u6_n88 ) );
  AOI21_X1 u2_u4_u6_U12 (.B2( u2_u4_u6_n147 ) , .B1( u2_u4_u6_n148 ) , .ZN( u2_u4_u6_n149 ) , .A( u2_u4_u6_n158 ) );
  AOI21_X1 u2_u4_u6_U13 (.ZN( u2_u4_u6_n106 ) , .A( u2_u4_u6_n142 ) , .B2( u2_u4_u6_n159 ) , .B1( u2_u4_u6_n164 ) );
  INV_X1 u2_u4_u6_U14 (.A( u2_u4_u6_n155 ) , .ZN( u2_u4_u6_n161 ) );
  INV_X1 u2_u4_u6_U15 (.A( u2_u4_u6_n128 ) , .ZN( u2_u4_u6_n164 ) );
  NAND2_X1 u2_u4_u6_U16 (.ZN( u2_u4_u6_n110 ) , .A1( u2_u4_u6_n122 ) , .A2( u2_u4_u6_n129 ) );
  NAND2_X1 u2_u4_u6_U17 (.ZN( u2_u4_u6_n124 ) , .A2( u2_u4_u6_n146 ) , .A1( u2_u4_u6_n148 ) );
  INV_X1 u2_u4_u6_U18 (.A( u2_u4_u6_n132 ) , .ZN( u2_u4_u6_n171 ) );
  AND2_X1 u2_u4_u6_U19 (.A1( u2_u4_u6_n100 ) , .ZN( u2_u4_u6_n130 ) , .A2( u2_u4_u6_n147 ) );
  INV_X1 u2_u4_u6_U20 (.A( u2_u4_u6_n127 ) , .ZN( u2_u4_u6_n173 ) );
  INV_X1 u2_u4_u6_U21 (.A( u2_u4_u6_n121 ) , .ZN( u2_u4_u6_n167 ) );
  INV_X1 u2_u4_u6_U22 (.A( u2_u4_u6_n100 ) , .ZN( u2_u4_u6_n169 ) );
  INV_X1 u2_u4_u6_U23 (.A( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n170 ) );
  INV_X1 u2_u4_u6_U24 (.A( u2_u4_u6_n113 ) , .ZN( u2_u4_u6_n168 ) );
  AND2_X1 u2_u4_u6_U25 (.A1( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n119 ) , .ZN( u2_u4_u6_n133 ) );
  AND2_X1 u2_u4_u6_U26 (.A2( u2_u4_u6_n121 ) , .A1( u2_u4_u6_n122 ) , .ZN( u2_u4_u6_n131 ) );
  AND3_X1 u2_u4_u6_U27 (.ZN( u2_u4_u6_n120 ) , .A2( u2_u4_u6_n127 ) , .A1( u2_u4_u6_n132 ) , .A3( u2_u4_u6_n145 ) );
  INV_X1 u2_u4_u6_U28 (.A( u2_u4_u6_n146 ) , .ZN( u2_u4_u6_n163 ) );
  AOI222_X1 u2_u4_u6_U29 (.ZN( u2_u4_u6_n114 ) , .A1( u2_u4_u6_n118 ) , .A2( u2_u4_u6_n126 ) , .B2( u2_u4_u6_n151 ) , .C2( u2_u4_u6_n159 ) , .C1( u2_u4_u6_n168 ) , .B1( u2_u4_u6_n169 ) );
  INV_X1 u2_u4_u6_U3 (.A( u2_u4_u6_n110 ) , .ZN( u2_u4_u6_n166 ) );
  NOR2_X1 u2_u4_u6_U30 (.A1( u2_u4_u6_n162 ) , .A2( u2_u4_u6_n165 ) , .ZN( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U31 (.A1( u2_u4_u6_n144 ) , .ZN( u2_u4_u6_n151 ) , .A2( u2_u4_u6_n158 ) );
  NAND2_X1 u2_u4_u6_U32 (.ZN( u2_u4_u6_n132 ) , .A1( u2_u4_u6_n91 ) , .A2( u2_u4_u6_n97 ) );
  AOI22_X1 u2_u4_u6_U33 (.B2( u2_u4_u6_n110 ) , .B1( u2_u4_u6_n111 ) , .A1( u2_u4_u6_n112 ) , .ZN( u2_u4_u6_n115 ) , .A2( u2_u4_u6_n161 ) );
  NAND4_X1 u2_u4_u6_U34 (.A3( u2_u4_u6_n109 ) , .ZN( u2_u4_u6_n112 ) , .A4( u2_u4_u6_n132 ) , .A2( u2_u4_u6_n147 ) , .A1( u2_u4_u6_n166 ) );
  NOR2_X1 u2_u4_u6_U35 (.ZN( u2_u4_u6_n109 ) , .A1( u2_u4_u6_n170 ) , .A2( u2_u4_u6_n173 ) );
  NOR2_X1 u2_u4_u6_U36 (.A2( u2_u4_u6_n126 ) , .ZN( u2_u4_u6_n155 ) , .A1( u2_u4_u6_n160 ) );
  NAND2_X1 u2_u4_u6_U37 (.ZN( u2_u4_u6_n146 ) , .A2( u2_u4_u6_n94 ) , .A1( u2_u4_u6_n99 ) );
  AOI21_X1 u2_u4_u6_U38 (.A( u2_u4_u6_n144 ) , .B2( u2_u4_u6_n145 ) , .B1( u2_u4_u6_n146 ) , .ZN( u2_u4_u6_n150 ) );
  AOI211_X1 u2_u4_u6_U39 (.B( u2_u4_u6_n134 ) , .A( u2_u4_u6_n135 ) , .C1( u2_u4_u6_n136 ) , .ZN( u2_u4_u6_n137 ) , .C2( u2_u4_u6_n151 ) );
  INV_X1 u2_u4_u6_U4 (.A( u2_u4_u6_n142 ) , .ZN( u2_u4_u6_n174 ) );
  NAND4_X1 u2_u4_u6_U40 (.A4( u2_u4_u6_n127 ) , .A3( u2_u4_u6_n128 ) , .A2( u2_u4_u6_n129 ) , .A1( u2_u4_u6_n130 ) , .ZN( u2_u4_u6_n136 ) );
  AOI21_X1 u2_u4_u6_U41 (.B2( u2_u4_u6_n132 ) , .B1( u2_u4_u6_n133 ) , .ZN( u2_u4_u6_n134 ) , .A( u2_u4_u6_n158 ) );
  AOI21_X1 u2_u4_u6_U42 (.B1( u2_u4_u6_n131 ) , .ZN( u2_u4_u6_n135 ) , .A( u2_u4_u6_n144 ) , .B2( u2_u4_u6_n146 ) );
  INV_X1 u2_u4_u6_U43 (.A( u2_u4_u6_n111 ) , .ZN( u2_u4_u6_n158 ) );
  NAND2_X1 u2_u4_u6_U44 (.ZN( u2_u4_u6_n127 ) , .A1( u2_u4_u6_n91 ) , .A2( u2_u4_u6_n92 ) );
  NAND2_X1 u2_u4_u6_U45 (.ZN( u2_u4_u6_n129 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n96 ) );
  INV_X1 u2_u4_u6_U46 (.A( u2_u4_u6_n144 ) , .ZN( u2_u4_u6_n159 ) );
  NAND2_X1 u2_u4_u6_U47 (.ZN( u2_u4_u6_n145 ) , .A2( u2_u4_u6_n97 ) , .A1( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U48 (.ZN( u2_u4_u6_n148 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n94 ) );
  NAND2_X1 u2_u4_u6_U49 (.ZN( u2_u4_u6_n108 ) , .A2( u2_u4_u6_n139 ) , .A1( u2_u4_u6_n144 ) );
  NAND2_X1 u2_u4_u6_U5 (.A2( u2_u4_u6_n143 ) , .ZN( u2_u4_u6_n152 ) , .A1( u2_u4_u6_n166 ) );
  NAND2_X1 u2_u4_u6_U50 (.ZN( u2_u4_u6_n121 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n97 ) );
  NAND2_X1 u2_u4_u6_U51 (.ZN( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n95 ) );
  AND2_X1 u2_u4_u6_U52 (.ZN( u2_u4_u6_n118 ) , .A2( u2_u4_u6_n91 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U53 (.ZN( u2_u4_u6_n147 ) , .A2( u2_u4_u6_n98 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U54 (.ZN( u2_u4_u6_n128 ) , .A1( u2_u4_u6_n94 ) , .A2( u2_u4_u6_n96 ) );
  NAND2_X1 u2_u4_u6_U55 (.ZN( u2_u4_u6_n119 ) , .A2( u2_u4_u6_n95 ) , .A1( u2_u4_u6_n99 ) );
  NAND2_X1 u2_u4_u6_U56 (.ZN( u2_u4_u6_n123 ) , .A2( u2_u4_u6_n91 ) , .A1( u2_u4_u6_n96 ) );
  NAND2_X1 u2_u4_u6_U57 (.ZN( u2_u4_u6_n100 ) , .A2( u2_u4_u6_n92 ) , .A1( u2_u4_u6_n98 ) );
  NAND2_X1 u2_u4_u6_U58 (.ZN( u2_u4_u6_n122 ) , .A1( u2_u4_u6_n94 ) , .A2( u2_u4_u6_n97 ) );
  INV_X1 u2_u4_u6_U59 (.A( u2_u4_u6_n139 ) , .ZN( u2_u4_u6_n160 ) );
  AOI22_X1 u2_u4_u6_U6 (.B2( u2_u4_u6_n101 ) , .A1( u2_u4_u6_n102 ) , .ZN( u2_u4_u6_n103 ) , .B1( u2_u4_u6_n160 ) , .A2( u2_u4_u6_n161 ) );
  NAND2_X1 u2_u4_u6_U60 (.ZN( u2_u4_u6_n113 ) , .A1( u2_u4_u6_n96 ) , .A2( u2_u4_u6_n98 ) );
  NOR2_X1 u2_u4_u6_U61 (.A2( u2_u4_X_40 ) , .A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n126 ) );
  NOR2_X1 u2_u4_u6_U62 (.A2( u2_u4_X_39 ) , .A1( u2_u4_X_42 ) , .ZN( u2_u4_u6_n92 ) );
  NOR2_X1 u2_u4_u6_U63 (.A2( u2_u4_X_39 ) , .A1( u2_u4_u6_n156 ) , .ZN( u2_u4_u6_n97 ) );
  NOR2_X1 u2_u4_u6_U64 (.A2( u2_u4_X_38 ) , .A1( u2_u4_u6_n165 ) , .ZN( u2_u4_u6_n95 ) );
  NOR2_X1 u2_u4_u6_U65 (.A2( u2_u4_X_41 ) , .ZN( u2_u4_u6_n111 ) , .A1( u2_u4_u6_n157 ) );
  NOR2_X1 u2_u4_u6_U66 (.A2( u2_u4_X_37 ) , .A1( u2_u4_u6_n162 ) , .ZN( u2_u4_u6_n94 ) );
  NOR2_X1 u2_u4_u6_U67 (.A2( u2_u4_X_37 ) , .A1( u2_u4_X_38 ) , .ZN( u2_u4_u6_n91 ) );
  NAND2_X1 u2_u4_u6_U68 (.A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n144 ) , .A2( u2_u4_u6_n157 ) );
  NAND2_X1 u2_u4_u6_U69 (.A2( u2_u4_X_40 ) , .A1( u2_u4_X_41 ) , .ZN( u2_u4_u6_n139 ) );
  NOR2_X1 u2_u4_u6_U7 (.A1( u2_u4_u6_n118 ) , .ZN( u2_u4_u6_n143 ) , .A2( u2_u4_u6_n168 ) );
  AND2_X1 u2_u4_u6_U70 (.A1( u2_u4_X_39 ) , .A2( u2_u4_u6_n156 ) , .ZN( u2_u4_u6_n96 ) );
  AND2_X1 u2_u4_u6_U71 (.A1( u2_u4_X_39 ) , .A2( u2_u4_X_42 ) , .ZN( u2_u4_u6_n99 ) );
  INV_X1 u2_u4_u6_U72 (.A( u2_u4_X_40 ) , .ZN( u2_u4_u6_n157 ) );
  INV_X1 u2_u4_u6_U73 (.A( u2_u4_X_37 ) , .ZN( u2_u4_u6_n165 ) );
  INV_X1 u2_u4_u6_U74 (.A( u2_u4_X_38 ) , .ZN( u2_u4_u6_n162 ) );
  INV_X1 u2_u4_u6_U75 (.A( u2_u4_X_42 ) , .ZN( u2_u4_u6_n156 ) );
  NAND4_X1 u2_u4_u6_U76 (.ZN( u2_out4_32 ) , .A4( u2_u4_u6_n103 ) , .A3( u2_u4_u6_n104 ) , .A2( u2_u4_u6_n105 ) , .A1( u2_u4_u6_n106 ) );
  AOI22_X1 u2_u4_u6_U77 (.ZN( u2_u4_u6_n105 ) , .A2( u2_u4_u6_n108 ) , .A1( u2_u4_u6_n118 ) , .B2( u2_u4_u6_n126 ) , .B1( u2_u4_u6_n171 ) );
  AOI22_X1 u2_u4_u6_U78 (.ZN( u2_u4_u6_n104 ) , .A1( u2_u4_u6_n111 ) , .B1( u2_u4_u6_n124 ) , .B2( u2_u4_u6_n151 ) , .A2( u2_u4_u6_n93 ) );
  NAND4_X1 u2_u4_u6_U79 (.ZN( u2_out4_12 ) , .A4( u2_u4_u6_n114 ) , .A3( u2_u4_u6_n115 ) , .A2( u2_u4_u6_n116 ) , .A1( u2_u4_u6_n117 ) );
  INV_X1 u2_u4_u6_U8 (.ZN( u2_u4_u6_n172 ) , .A( u2_u4_u6_n88 ) );
  OAI22_X1 u2_u4_u6_U80 (.B2( u2_u4_u6_n111 ) , .ZN( u2_u4_u6_n116 ) , .B1( u2_u4_u6_n126 ) , .A2( u2_u4_u6_n164 ) , .A1( u2_u4_u6_n167 ) );
  OAI21_X1 u2_u4_u6_U81 (.A( u2_u4_u6_n108 ) , .ZN( u2_u4_u6_n117 ) , .B2( u2_u4_u6_n141 ) , .B1( u2_u4_u6_n163 ) );
  OAI211_X1 u2_u4_u6_U82 (.ZN( u2_out4_22 ) , .B( u2_u4_u6_n137 ) , .A( u2_u4_u6_n138 ) , .C2( u2_u4_u6_n139 ) , .C1( u2_u4_u6_n140 ) );
  AOI22_X1 u2_u4_u6_U83 (.B1( u2_u4_u6_n124 ) , .A2( u2_u4_u6_n125 ) , .A1( u2_u4_u6_n126 ) , .ZN( u2_u4_u6_n138 ) , .B2( u2_u4_u6_n161 ) );
  AND4_X1 u2_u4_u6_U84 (.A3( u2_u4_u6_n119 ) , .A1( u2_u4_u6_n120 ) , .A4( u2_u4_u6_n129 ) , .ZN( u2_u4_u6_n140 ) , .A2( u2_u4_u6_n143 ) );
  OAI211_X1 u2_u4_u6_U85 (.ZN( u2_out4_7 ) , .B( u2_u4_u6_n153 ) , .C2( u2_u4_u6_n154 ) , .C1( u2_u4_u6_n155 ) , .A( u2_u4_u6_n174 ) );
  NOR3_X1 u2_u4_u6_U86 (.A1( u2_u4_u6_n141 ) , .ZN( u2_u4_u6_n154 ) , .A3( u2_u4_u6_n164 ) , .A2( u2_u4_u6_n171 ) );
  AOI211_X1 u2_u4_u6_U87 (.B( u2_u4_u6_n149 ) , .A( u2_u4_u6_n150 ) , .C2( u2_u4_u6_n151 ) , .C1( u2_u4_u6_n152 ) , .ZN( u2_u4_u6_n153 ) );
  NAND3_X1 u2_u4_u6_U88 (.A2( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n125 ) , .A1( u2_u4_u6_n130 ) , .A3( u2_u4_u6_n131 ) );
  NAND3_X1 u2_u4_u6_U89 (.A3( u2_u4_u6_n133 ) , .ZN( u2_u4_u6_n141 ) , .A1( u2_u4_u6_n145 ) , .A2( u2_u4_u6_n148 ) );
  OAI21_X1 u2_u4_u6_U9 (.A( u2_u4_u6_n159 ) , .B1( u2_u4_u6_n169 ) , .B2( u2_u4_u6_n173 ) , .ZN( u2_u4_u6_n90 ) );
  NAND3_X1 u2_u4_u6_U90 (.ZN( u2_u4_u6_n101 ) , .A3( u2_u4_u6_n107 ) , .A2( u2_u4_u6_n121 ) , .A1( u2_u4_u6_n127 ) );
  NAND3_X1 u2_u4_u6_U91 (.ZN( u2_u4_u6_n102 ) , .A3( u2_u4_u6_n130 ) , .A2( u2_u4_u6_n145 ) , .A1( u2_u4_u6_n166 ) );
  NAND3_X1 u2_u4_u6_U92 (.A3( u2_u4_u6_n113 ) , .A1( u2_u4_u6_n119 ) , .A2( u2_u4_u6_n123 ) , .ZN( u2_u4_u6_n93 ) );
  NAND3_X1 u2_u4_u6_U93 (.ZN( u2_u4_u6_n142 ) , .A2( u2_u4_u6_n172 ) , .A3( u2_u4_u6_n89 ) , .A1( u2_u4_u6_n90 ) );
  XOR2_X1 u2_u5_U1 (.B( u2_K6_9 ) , .A( u2_R4_6 ) , .Z( u2_u5_X_9 ) );
  XOR2_X1 u2_u5_U10 (.B( u2_K6_45 ) , .A( u2_R4_30 ) , .Z( u2_u5_X_45 ) );
  XOR2_X1 u2_u5_U11 (.B( u2_K6_44 ) , .A( u2_R4_29 ) , .Z( u2_u5_X_44 ) );
  XOR2_X1 u2_u5_U12 (.B( u2_K6_43 ) , .A( u2_R4_28 ) , .Z( u2_u5_X_43 ) );
  XOR2_X1 u2_u5_U13 (.B( u2_K6_42 ) , .A( u2_R4_29 ) , .Z( u2_u5_X_42 ) );
  XOR2_X1 u2_u5_U14 (.B( u2_K6_41 ) , .A( u2_R4_28 ) , .Z( u2_u5_X_41 ) );
  XOR2_X1 u2_u5_U15 (.B( u2_K6_40 ) , .A( u2_R4_27 ) , .Z( u2_u5_X_40 ) );
  XOR2_X1 u2_u5_U16 (.B( u2_K6_3 ) , .A( u2_R4_2 ) , .Z( u2_u5_X_3 ) );
  XOR2_X1 u2_u5_U17 (.B( u2_K6_39 ) , .A( u2_R4_26 ) , .Z( u2_u5_X_39 ) );
  XOR2_X1 u2_u5_U18 (.B( u2_K6_38 ) , .A( u2_R4_25 ) , .Z( u2_u5_X_38 ) );
  XOR2_X1 u2_u5_U19 (.B( u2_K6_37 ) , .A( u2_R4_24 ) , .Z( u2_u5_X_37 ) );
  XOR2_X1 u2_u5_U2 (.B( u2_K6_8 ) , .A( u2_R4_5 ) , .Z( u2_u5_X_8 ) );
  XOR2_X1 u2_u5_U20 (.B( u2_K6_36 ) , .A( u2_R4_25 ) , .Z( u2_u5_X_36 ) );
  XOR2_X1 u2_u5_U21 (.B( u2_K6_35 ) , .A( u2_R4_24 ) , .Z( u2_u5_X_35 ) );
  XOR2_X1 u2_u5_U22 (.B( u2_K6_34 ) , .A( u2_R4_23 ) , .Z( u2_u5_X_34 ) );
  XOR2_X1 u2_u5_U23 (.B( u2_K6_33 ) , .A( u2_R4_22 ) , .Z( u2_u5_X_33 ) );
  XOR2_X1 u2_u5_U24 (.B( u2_K6_32 ) , .A( u2_R4_21 ) , .Z( u2_u5_X_32 ) );
  XOR2_X1 u2_u5_U25 (.B( u2_K6_31 ) , .A( u2_R4_20 ) , .Z( u2_u5_X_31 ) );
  XOR2_X1 u2_u5_U27 (.B( u2_K6_2 ) , .A( u2_R4_1 ) , .Z( u2_u5_X_2 ) );
  XOR2_X1 u2_u5_U3 (.B( u2_K6_7 ) , .A( u2_R4_4 ) , .Z( u2_u5_X_7 ) );
  XOR2_X1 u2_u5_U38 (.B( u2_K6_1 ) , .A( u2_R4_32 ) , .Z( u2_u5_X_1 ) );
  XOR2_X1 u2_u5_U4 (.B( u2_K6_6 ) , .A( u2_R4_5 ) , .Z( u2_u5_X_6 ) );
  XOR2_X1 u2_u5_U46 (.B( u2_K6_12 ) , .A( u2_R4_9 ) , .Z( u2_u5_X_12 ) );
  XOR2_X1 u2_u5_U47 (.B( u2_K6_11 ) , .A( u2_R4_8 ) , .Z( u2_u5_X_11 ) );
  XOR2_X1 u2_u5_U48 (.B( u2_K6_10 ) , .A( u2_R4_7 ) , .Z( u2_u5_X_10 ) );
  XOR2_X1 u2_u5_U5 (.B( u2_K6_5 ) , .A( u2_R4_4 ) , .Z( u2_u5_X_5 ) );
  XOR2_X1 u2_u5_U6 (.B( u2_K6_4 ) , .A( u2_R4_3 ) , .Z( u2_u5_X_4 ) );
  XOR2_X1 u2_u5_U7 (.B( u2_K6_48 ) , .A( u2_R4_1 ) , .Z( u2_u5_X_48 ) );
  XOR2_X1 u2_u5_U8 (.B( u2_K6_47 ) , .A( u2_R4_32 ) , .Z( u2_u5_X_47 ) );
  XOR2_X1 u2_u5_U9 (.B( u2_K6_46 ) , .A( u2_R4_31 ) , .Z( u2_u5_X_46 ) );
  AND3_X1 u2_u5_u0_U10 (.A2( u2_u5_u0_n112 ) , .ZN( u2_u5_u0_n127 ) , .A3( u2_u5_u0_n130 ) , .A1( u2_u5_u0_n148 ) );
  NAND2_X1 u2_u5_u0_U11 (.ZN( u2_u5_u0_n113 ) , .A1( u2_u5_u0_n139 ) , .A2( u2_u5_u0_n149 ) );
  AND2_X1 u2_u5_u0_U12 (.ZN( u2_u5_u0_n107 ) , .A1( u2_u5_u0_n130 ) , .A2( u2_u5_u0_n140 ) );
  AND2_X1 u2_u5_u0_U13 (.A2( u2_u5_u0_n129 ) , .A1( u2_u5_u0_n130 ) , .ZN( u2_u5_u0_n151 ) );
  AND2_X1 u2_u5_u0_U14 (.A1( u2_u5_u0_n108 ) , .A2( u2_u5_u0_n125 ) , .ZN( u2_u5_u0_n145 ) );
  INV_X1 u2_u5_u0_U15 (.A( u2_u5_u0_n143 ) , .ZN( u2_u5_u0_n173 ) );
  NOR2_X1 u2_u5_u0_U16 (.A2( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n147 ) , .A1( u2_u5_u0_n160 ) );
  AOI21_X1 u2_u5_u0_U17 (.B1( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n132 ) , .A( u2_u5_u0_n165 ) , .B2( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U18 (.A( u2_u5_u0_n142 ) , .ZN( u2_u5_u0_n165 ) );
  OAI22_X1 u2_u5_u0_U19 (.B1( u2_u5_u0_n125 ) , .ZN( u2_u5_u0_n126 ) , .A1( u2_u5_u0_n138 ) , .A2( u2_u5_u0_n146 ) , .B2( u2_u5_u0_n147 ) );
  OAI22_X1 u2_u5_u0_U20 (.B1( u2_u5_u0_n131 ) , .A1( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n147 ) , .A2( u2_u5_u0_n90 ) , .ZN( u2_u5_u0_n91 ) );
  AND3_X1 u2_u5_u0_U21 (.A3( u2_u5_u0_n121 ) , .A2( u2_u5_u0_n125 ) , .A1( u2_u5_u0_n148 ) , .ZN( u2_u5_u0_n90 ) );
  INV_X1 u2_u5_u0_U22 (.A( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n161 ) );
  AOI22_X1 u2_u5_u0_U23 (.B2( u2_u5_u0_n109 ) , .A2( u2_u5_u0_n110 ) , .ZN( u2_u5_u0_n111 ) , .B1( u2_u5_u0_n118 ) , .A1( u2_u5_u0_n160 ) );
  INV_X1 u2_u5_u0_U24 (.A( u2_u5_u0_n118 ) , .ZN( u2_u5_u0_n158 ) );
  AOI21_X1 u2_u5_u0_U25 (.ZN( u2_u5_u0_n104 ) , .B1( u2_u5_u0_n107 ) , .B2( u2_u5_u0_n141 ) , .A( u2_u5_u0_n144 ) );
  AOI21_X1 u2_u5_u0_U26 (.B1( u2_u5_u0_n127 ) , .B2( u2_u5_u0_n129 ) , .A( u2_u5_u0_n138 ) , .ZN( u2_u5_u0_n96 ) );
  AOI21_X1 u2_u5_u0_U27 (.ZN( u2_u5_u0_n116 ) , .B2( u2_u5_u0_n142 ) , .A( u2_u5_u0_n144 ) , .B1( u2_u5_u0_n166 ) );
  NOR2_X1 u2_u5_u0_U28 (.A1( u2_u5_u0_n120 ) , .ZN( u2_u5_u0_n143 ) , .A2( u2_u5_u0_n167 ) );
  OAI221_X1 u2_u5_u0_U29 (.C1( u2_u5_u0_n112 ) , .ZN( u2_u5_u0_n120 ) , .B1( u2_u5_u0_n138 ) , .B2( u2_u5_u0_n141 ) , .C2( u2_u5_u0_n147 ) , .A( u2_u5_u0_n172 ) );
  INV_X1 u2_u5_u0_U3 (.A( u2_u5_u0_n113 ) , .ZN( u2_u5_u0_n166 ) );
  AOI211_X1 u2_u5_u0_U30 (.B( u2_u5_u0_n115 ) , .A( u2_u5_u0_n116 ) , .C2( u2_u5_u0_n117 ) , .C1( u2_u5_u0_n118 ) , .ZN( u2_u5_u0_n119 ) );
  NAND2_X1 u2_u5_u0_U31 (.A1( u2_u5_u0_n100 ) , .A2( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n125 ) );
  NAND2_X1 u2_u5_u0_U32 (.A2( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n140 ) , .A1( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U33 (.A1( u2_u5_u0_n101 ) , .A2( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n150 ) );
  INV_X1 u2_u5_u0_U34 (.A( u2_u5_u0_n138 ) , .ZN( u2_u5_u0_n160 ) );
  NAND2_X1 u2_u5_u0_U35 (.A2( u2_u5_u0_n102 ) , .A1( u2_u5_u0_n103 ) , .ZN( u2_u5_u0_n149 ) );
  NAND2_X1 u2_u5_u0_U36 (.A2( u2_u5_u0_n100 ) , .A1( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n139 ) );
  NAND2_X1 u2_u5_u0_U37 (.A2( u2_u5_u0_n100 ) , .ZN( u2_u5_u0_n131 ) , .A1( u2_u5_u0_n92 ) );
  NAND2_X1 u2_u5_u0_U38 (.ZN( u2_u5_u0_n108 ) , .A1( u2_u5_u0_n92 ) , .A2( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U39 (.A2( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n114 ) , .A1( u2_u5_u0_n92 ) );
  AOI21_X1 u2_u5_u0_U4 (.B1( u2_u5_u0_n114 ) , .ZN( u2_u5_u0_n115 ) , .B2( u2_u5_u0_n129 ) , .A( u2_u5_u0_n161 ) );
  NAND2_X1 u2_u5_u0_U40 (.A1( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n130 ) , .A2( u2_u5_u0_n94 ) );
  NAND2_X1 u2_u5_u0_U41 (.A2( u2_u5_u0_n101 ) , .ZN( u2_u5_u0_n121 ) , .A1( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U42 (.ZN( u2_u5_u0_n172 ) , .A( u2_u5_u0_n88 ) );
  OAI222_X1 u2_u5_u0_U43 (.C1( u2_u5_u0_n108 ) , .A1( u2_u5_u0_n125 ) , .B2( u2_u5_u0_n128 ) , .B1( u2_u5_u0_n144 ) , .A2( u2_u5_u0_n158 ) , .C2( u2_u5_u0_n161 ) , .ZN( u2_u5_u0_n88 ) );
  NAND2_X1 u2_u5_u0_U44 (.ZN( u2_u5_u0_n112 ) , .A2( u2_u5_u0_n92 ) , .A1( u2_u5_u0_n93 ) );
  OR3_X1 u2_u5_u0_U45 (.A3( u2_u5_u0_n152 ) , .A2( u2_u5_u0_n153 ) , .A1( u2_u5_u0_n154 ) , .ZN( u2_u5_u0_n155 ) );
  AOI21_X1 u2_u5_u0_U46 (.A( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n145 ) , .B1( u2_u5_u0_n146 ) , .ZN( u2_u5_u0_n154 ) );
  AOI21_X1 u2_u5_u0_U47 (.B2( u2_u5_u0_n150 ) , .B1( u2_u5_u0_n151 ) , .ZN( u2_u5_u0_n152 ) , .A( u2_u5_u0_n158 ) );
  AOI21_X1 u2_u5_u0_U48 (.A( u2_u5_u0_n147 ) , .B2( u2_u5_u0_n148 ) , .B1( u2_u5_u0_n149 ) , .ZN( u2_u5_u0_n153 ) );
  INV_X1 u2_u5_u0_U49 (.ZN( u2_u5_u0_n171 ) , .A( u2_u5_u0_n99 ) );
  AOI21_X1 u2_u5_u0_U5 (.B2( u2_u5_u0_n131 ) , .ZN( u2_u5_u0_n134 ) , .B1( u2_u5_u0_n151 ) , .A( u2_u5_u0_n158 ) );
  OAI211_X1 u2_u5_u0_U50 (.C2( u2_u5_u0_n140 ) , .C1( u2_u5_u0_n161 ) , .A( u2_u5_u0_n169 ) , .B( u2_u5_u0_n98 ) , .ZN( u2_u5_u0_n99 ) );
  AOI211_X1 u2_u5_u0_U51 (.C1( u2_u5_u0_n118 ) , .A( u2_u5_u0_n123 ) , .B( u2_u5_u0_n96 ) , .C2( u2_u5_u0_n97 ) , .ZN( u2_u5_u0_n98 ) );
  INV_X1 u2_u5_u0_U52 (.ZN( u2_u5_u0_n169 ) , .A( u2_u5_u0_n91 ) );
  NOR2_X1 u2_u5_u0_U53 (.A2( u2_u5_X_2 ) , .ZN( u2_u5_u0_n103 ) , .A1( u2_u5_u0_n164 ) );
  NOR2_X1 u2_u5_u0_U54 (.A2( u2_u5_X_4 ) , .A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n118 ) );
  NOR2_X1 u2_u5_u0_U55 (.A2( u2_u5_X_1 ) , .A1( u2_u5_X_2 ) , .ZN( u2_u5_u0_n92 ) );
  NOR2_X1 u2_u5_u0_U56 (.A2( u2_u5_X_1 ) , .ZN( u2_u5_u0_n101 ) , .A1( u2_u5_u0_n163 ) );
  NOR2_X1 u2_u5_u0_U57 (.A2( u2_u5_X_3 ) , .A1( u2_u5_X_6 ) , .ZN( u2_u5_u0_n94 ) );
  NOR2_X1 u2_u5_u0_U58 (.A2( u2_u5_X_6 ) , .ZN( u2_u5_u0_n100 ) , .A1( u2_u5_u0_n162 ) );
  NAND2_X1 u2_u5_u0_U59 (.A2( u2_u5_X_4 ) , .A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n144 ) );
  NOR2_X1 u2_u5_u0_U6 (.A1( u2_u5_u0_n108 ) , .ZN( u2_u5_u0_n123 ) , .A2( u2_u5_u0_n158 ) );
  NOR2_X1 u2_u5_u0_U60 (.A2( u2_u5_X_5 ) , .ZN( u2_u5_u0_n136 ) , .A1( u2_u5_u0_n159 ) );
  NAND2_X1 u2_u5_u0_U61 (.A1( u2_u5_X_5 ) , .ZN( u2_u5_u0_n138 ) , .A2( u2_u5_u0_n159 ) );
  AND2_X1 u2_u5_u0_U62 (.A2( u2_u5_X_3 ) , .A1( u2_u5_X_6 ) , .ZN( u2_u5_u0_n102 ) );
  AND2_X1 u2_u5_u0_U63 (.A1( u2_u5_X_6 ) , .A2( u2_u5_u0_n162 ) , .ZN( u2_u5_u0_n93 ) );
  INV_X1 u2_u5_u0_U64 (.A( u2_u5_X_4 ) , .ZN( u2_u5_u0_n159 ) );
  INV_X1 u2_u5_u0_U65 (.A( u2_u5_X_1 ) , .ZN( u2_u5_u0_n164 ) );
  INV_X1 u2_u5_u0_U66 (.A( u2_u5_X_2 ) , .ZN( u2_u5_u0_n163 ) );
  INV_X1 u2_u5_u0_U67 (.A( u2_u5_X_3 ) , .ZN( u2_u5_u0_n162 ) );
  INV_X1 u2_u5_u0_U68 (.A( u2_u5_u0_n126 ) , .ZN( u2_u5_u0_n168 ) );
  AOI211_X1 u2_u5_u0_U69 (.B( u2_u5_u0_n133 ) , .A( u2_u5_u0_n134 ) , .C2( u2_u5_u0_n135 ) , .C1( u2_u5_u0_n136 ) , .ZN( u2_u5_u0_n137 ) );
  OAI21_X1 u2_u5_u0_U7 (.B1( u2_u5_u0_n150 ) , .B2( u2_u5_u0_n158 ) , .A( u2_u5_u0_n172 ) , .ZN( u2_u5_u0_n89 ) );
  OR4_X1 u2_u5_u0_U70 (.ZN( u2_out5_17 ) , .A4( u2_u5_u0_n122 ) , .A2( u2_u5_u0_n123 ) , .A1( u2_u5_u0_n124 ) , .A3( u2_u5_u0_n170 ) );
  AOI21_X1 u2_u5_u0_U71 (.B2( u2_u5_u0_n107 ) , .ZN( u2_u5_u0_n124 ) , .B1( u2_u5_u0_n128 ) , .A( u2_u5_u0_n161 ) );
  INV_X1 u2_u5_u0_U72 (.A( u2_u5_u0_n111 ) , .ZN( u2_u5_u0_n170 ) );
  OR4_X1 u2_u5_u0_U73 (.ZN( u2_out5_31 ) , .A4( u2_u5_u0_n155 ) , .A2( u2_u5_u0_n156 ) , .A1( u2_u5_u0_n157 ) , .A3( u2_u5_u0_n173 ) );
  AOI21_X1 u2_u5_u0_U74 (.A( u2_u5_u0_n138 ) , .B2( u2_u5_u0_n139 ) , .B1( u2_u5_u0_n140 ) , .ZN( u2_u5_u0_n157 ) );
  AOI21_X1 u2_u5_u0_U75 (.B2( u2_u5_u0_n141 ) , .B1( u2_u5_u0_n142 ) , .ZN( u2_u5_u0_n156 ) , .A( u2_u5_u0_n161 ) );
  INV_X1 u2_u5_u0_U76 (.ZN( u2_u5_u0_n174 ) , .A( u2_u5_u0_n89 ) );
  AOI211_X1 u2_u5_u0_U77 (.B( u2_u5_u0_n104 ) , .A( u2_u5_u0_n105 ) , .ZN( u2_u5_u0_n106 ) , .C2( u2_u5_u0_n113 ) , .C1( u2_u5_u0_n160 ) );
  NOR2_X1 u2_u5_u0_U78 (.A1( u2_u5_u0_n163 ) , .A2( u2_u5_u0_n164 ) , .ZN( u2_u5_u0_n95 ) );
  OAI221_X1 u2_u5_u0_U79 (.C1( u2_u5_u0_n121 ) , .ZN( u2_u5_u0_n122 ) , .B2( u2_u5_u0_n127 ) , .A( u2_u5_u0_n143 ) , .B1( u2_u5_u0_n144 ) , .C2( u2_u5_u0_n147 ) );
  AND2_X1 u2_u5_u0_U8 (.A1( u2_u5_u0_n114 ) , .A2( u2_u5_u0_n121 ) , .ZN( u2_u5_u0_n146 ) );
  AOI21_X1 u2_u5_u0_U80 (.B1( u2_u5_u0_n132 ) , .ZN( u2_u5_u0_n133 ) , .A( u2_u5_u0_n144 ) , .B2( u2_u5_u0_n166 ) );
  OAI22_X1 u2_u5_u0_U81 (.ZN( u2_u5_u0_n105 ) , .A2( u2_u5_u0_n132 ) , .B1( u2_u5_u0_n146 ) , .A1( u2_u5_u0_n147 ) , .B2( u2_u5_u0_n161 ) );
  NAND2_X1 u2_u5_u0_U82 (.ZN( u2_u5_u0_n110 ) , .A2( u2_u5_u0_n132 ) , .A1( u2_u5_u0_n145 ) );
  INV_X1 u2_u5_u0_U83 (.A( u2_u5_u0_n119 ) , .ZN( u2_u5_u0_n167 ) );
  NAND2_X1 u2_u5_u0_U84 (.ZN( u2_u5_u0_n148 ) , .A1( u2_u5_u0_n93 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U85 (.A1( u2_u5_u0_n100 ) , .ZN( u2_u5_u0_n129 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U86 (.A1( u2_u5_u0_n102 ) , .ZN( u2_u5_u0_n128 ) , .A2( u2_u5_u0_n95 ) );
  NAND2_X1 u2_u5_u0_U87 (.ZN( u2_u5_u0_n142 ) , .A1( u2_u5_u0_n94 ) , .A2( u2_u5_u0_n95 ) );
  NAND3_X1 u2_u5_u0_U88 (.ZN( u2_out5_23 ) , .A3( u2_u5_u0_n137 ) , .A1( u2_u5_u0_n168 ) , .A2( u2_u5_u0_n171 ) );
  NAND3_X1 u2_u5_u0_U89 (.A3( u2_u5_u0_n127 ) , .A2( u2_u5_u0_n128 ) , .ZN( u2_u5_u0_n135 ) , .A1( u2_u5_u0_n150 ) );
  AND2_X1 u2_u5_u0_U9 (.A1( u2_u5_u0_n131 ) , .ZN( u2_u5_u0_n141 ) , .A2( u2_u5_u0_n150 ) );
  NAND3_X1 u2_u5_u0_U90 (.ZN( u2_u5_u0_n117 ) , .A3( u2_u5_u0_n132 ) , .A2( u2_u5_u0_n139 ) , .A1( u2_u5_u0_n148 ) );
  NAND3_X1 u2_u5_u0_U91 (.ZN( u2_u5_u0_n109 ) , .A2( u2_u5_u0_n114 ) , .A3( u2_u5_u0_n140 ) , .A1( u2_u5_u0_n149 ) );
  NAND3_X1 u2_u5_u0_U92 (.ZN( u2_out5_9 ) , .A3( u2_u5_u0_n106 ) , .A2( u2_u5_u0_n171 ) , .A1( u2_u5_u0_n174 ) );
  NAND3_X1 u2_u5_u0_U93 (.A2( u2_u5_u0_n128 ) , .A1( u2_u5_u0_n132 ) , .A3( u2_u5_u0_n146 ) , .ZN( u2_u5_u0_n97 ) );
  NOR2_X1 u2_u5_u1_U10 (.A1( u2_u5_u1_n112 ) , .A2( u2_u5_u1_n116 ) , .ZN( u2_u5_u1_n118 ) );
  NAND3_X1 u2_u5_u1_U100 (.ZN( u2_u5_u1_n113 ) , .A1( u2_u5_u1_n120 ) , .A3( u2_u5_u1_n133 ) , .A2( u2_u5_u1_n155 ) );
  OAI21_X1 u2_u5_u1_U11 (.ZN( u2_u5_u1_n101 ) , .B1( u2_u5_u1_n141 ) , .A( u2_u5_u1_n146 ) , .B2( u2_u5_u1_n183 ) );
  AOI21_X1 u2_u5_u1_U12 (.B2( u2_u5_u1_n155 ) , .B1( u2_u5_u1_n156 ) , .ZN( u2_u5_u1_n157 ) , .A( u2_u5_u1_n174 ) );
  NAND2_X1 u2_u5_u1_U13 (.ZN( u2_u5_u1_n140 ) , .A2( u2_u5_u1_n150 ) , .A1( u2_u5_u1_n155 ) );
  NAND2_X1 u2_u5_u1_U14 (.A1( u2_u5_u1_n131 ) , .ZN( u2_u5_u1_n147 ) , .A2( u2_u5_u1_n153 ) );
  INV_X1 u2_u5_u1_U15 (.A( u2_u5_u1_n139 ) , .ZN( u2_u5_u1_n174 ) );
  OR4_X1 u2_u5_u1_U16 (.A4( u2_u5_u1_n106 ) , .A3( u2_u5_u1_n107 ) , .ZN( u2_u5_u1_n108 ) , .A1( u2_u5_u1_n117 ) , .A2( u2_u5_u1_n184 ) );
  AOI21_X1 u2_u5_u1_U17 (.ZN( u2_u5_u1_n106 ) , .A( u2_u5_u1_n112 ) , .B1( u2_u5_u1_n154 ) , .B2( u2_u5_u1_n156 ) );
  INV_X1 u2_u5_u1_U18 (.A( u2_u5_u1_n101 ) , .ZN( u2_u5_u1_n184 ) );
  AOI21_X1 u2_u5_u1_U19 (.ZN( u2_u5_u1_n107 ) , .B1( u2_u5_u1_n134 ) , .B2( u2_u5_u1_n149 ) , .A( u2_u5_u1_n174 ) );
  INV_X1 u2_u5_u1_U20 (.A( u2_u5_u1_n112 ) , .ZN( u2_u5_u1_n171 ) );
  NAND2_X1 u2_u5_u1_U21 (.ZN( u2_u5_u1_n141 ) , .A1( u2_u5_u1_n153 ) , .A2( u2_u5_u1_n156 ) );
  AND2_X1 u2_u5_u1_U22 (.A1( u2_u5_u1_n123 ) , .ZN( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n161 ) );
  NAND2_X1 u2_u5_u1_U23 (.A2( u2_u5_u1_n115 ) , .A1( u2_u5_u1_n116 ) , .ZN( u2_u5_u1_n148 ) );
  NAND2_X1 u2_u5_u1_U24 (.A2( u2_u5_u1_n133 ) , .A1( u2_u5_u1_n135 ) , .ZN( u2_u5_u1_n159 ) );
  NAND2_X1 u2_u5_u1_U25 (.A2( u2_u5_u1_n115 ) , .A1( u2_u5_u1_n120 ) , .ZN( u2_u5_u1_n132 ) );
  INV_X1 u2_u5_u1_U26 (.A( u2_u5_u1_n154 ) , .ZN( u2_u5_u1_n178 ) );
  INV_X1 u2_u5_u1_U27 (.A( u2_u5_u1_n151 ) , .ZN( u2_u5_u1_n183 ) );
  AND2_X1 u2_u5_u1_U28 (.A1( u2_u5_u1_n129 ) , .A2( u2_u5_u1_n133 ) , .ZN( u2_u5_u1_n149 ) );
  INV_X1 u2_u5_u1_U29 (.A( u2_u5_u1_n131 ) , .ZN( u2_u5_u1_n180 ) );
  INV_X1 u2_u5_u1_U3 (.A( u2_u5_u1_n159 ) , .ZN( u2_u5_u1_n182 ) );
  OAI221_X1 u2_u5_u1_U30 (.A( u2_u5_u1_n119 ) , .C2( u2_u5_u1_n129 ) , .ZN( u2_u5_u1_n138 ) , .B2( u2_u5_u1_n152 ) , .C1( u2_u5_u1_n174 ) , .B1( u2_u5_u1_n187 ) );
  INV_X1 u2_u5_u1_U31 (.A( u2_u5_u1_n148 ) , .ZN( u2_u5_u1_n187 ) );
  AOI211_X1 u2_u5_u1_U32 (.B( u2_u5_u1_n117 ) , .A( u2_u5_u1_n118 ) , .ZN( u2_u5_u1_n119 ) , .C2( u2_u5_u1_n146 ) , .C1( u2_u5_u1_n159 ) );
  NOR2_X1 u2_u5_u1_U33 (.A1( u2_u5_u1_n168 ) , .A2( u2_u5_u1_n176 ) , .ZN( u2_u5_u1_n98 ) );
  OAI21_X1 u2_u5_u1_U34 (.B2( u2_u5_u1_n123 ) , .ZN( u2_u5_u1_n145 ) , .B1( u2_u5_u1_n160 ) , .A( u2_u5_u1_n185 ) );
  INV_X1 u2_u5_u1_U35 (.A( u2_u5_u1_n122 ) , .ZN( u2_u5_u1_n185 ) );
  AOI21_X1 u2_u5_u1_U36 (.B2( u2_u5_u1_n120 ) , .B1( u2_u5_u1_n121 ) , .ZN( u2_u5_u1_n122 ) , .A( u2_u5_u1_n128 ) );
  NAND2_X1 u2_u5_u1_U37 (.A1( u2_u5_u1_n128 ) , .ZN( u2_u5_u1_n146 ) , .A2( u2_u5_u1_n160 ) );
  NAND2_X1 u2_u5_u1_U38 (.A2( u2_u5_u1_n112 ) , .ZN( u2_u5_u1_n139 ) , .A1( u2_u5_u1_n152 ) );
  NAND2_X1 u2_u5_u1_U39 (.A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n156 ) , .A2( u2_u5_u1_n99 ) );
  AOI221_X1 u2_u5_u1_U4 (.A( u2_u5_u1_n138 ) , .C2( u2_u5_u1_n139 ) , .C1( u2_u5_u1_n140 ) , .B2( u2_u5_u1_n141 ) , .ZN( u2_u5_u1_n142 ) , .B1( u2_u5_u1_n175 ) );
  AOI221_X1 u2_u5_u1_U40 (.B1( u2_u5_u1_n140 ) , .ZN( u2_u5_u1_n167 ) , .B2( u2_u5_u1_n172 ) , .C2( u2_u5_u1_n175 ) , .C1( u2_u5_u1_n178 ) , .A( u2_u5_u1_n188 ) );
  INV_X1 u2_u5_u1_U41 (.ZN( u2_u5_u1_n188 ) , .A( u2_u5_u1_n97 ) );
  AOI211_X1 u2_u5_u1_U42 (.A( u2_u5_u1_n118 ) , .C1( u2_u5_u1_n132 ) , .C2( u2_u5_u1_n139 ) , .B( u2_u5_u1_n96 ) , .ZN( u2_u5_u1_n97 ) );
  AOI21_X1 u2_u5_u1_U43 (.B2( u2_u5_u1_n121 ) , .B1( u2_u5_u1_n135 ) , .A( u2_u5_u1_n152 ) , .ZN( u2_u5_u1_n96 ) );
  NOR2_X1 u2_u5_u1_U44 (.ZN( u2_u5_u1_n117 ) , .A1( u2_u5_u1_n121 ) , .A2( u2_u5_u1_n160 ) );
  AOI21_X1 u2_u5_u1_U45 (.A( u2_u5_u1_n128 ) , .B2( u2_u5_u1_n129 ) , .ZN( u2_u5_u1_n130 ) , .B1( u2_u5_u1_n150 ) );
  NAND2_X1 u2_u5_u1_U46 (.ZN( u2_u5_u1_n112 ) , .A1( u2_u5_u1_n169 ) , .A2( u2_u5_u1_n170 ) );
  NAND2_X1 u2_u5_u1_U47 (.ZN( u2_u5_u1_n129 ) , .A2( u2_u5_u1_n95 ) , .A1( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U48 (.A1( u2_u5_u1_n102 ) , .ZN( u2_u5_u1_n154 ) , .A2( u2_u5_u1_n99 ) );
  NAND2_X1 u2_u5_u1_U49 (.A2( u2_u5_u1_n100 ) , .ZN( u2_u5_u1_n135 ) , .A1( u2_u5_u1_n99 ) );
  AOI211_X1 u2_u5_u1_U5 (.ZN( u2_u5_u1_n124 ) , .A( u2_u5_u1_n138 ) , .C2( u2_u5_u1_n139 ) , .B( u2_u5_u1_n145 ) , .C1( u2_u5_u1_n147 ) );
  AOI21_X1 u2_u5_u1_U50 (.A( u2_u5_u1_n152 ) , .B2( u2_u5_u1_n153 ) , .B1( u2_u5_u1_n154 ) , .ZN( u2_u5_u1_n158 ) );
  INV_X1 u2_u5_u1_U51 (.A( u2_u5_u1_n160 ) , .ZN( u2_u5_u1_n175 ) );
  NAND2_X1 u2_u5_u1_U52 (.A1( u2_u5_u1_n100 ) , .ZN( u2_u5_u1_n116 ) , .A2( u2_u5_u1_n95 ) );
  NAND2_X1 u2_u5_u1_U53 (.A1( u2_u5_u1_n102 ) , .ZN( u2_u5_u1_n131 ) , .A2( u2_u5_u1_n95 ) );
  NAND2_X1 u2_u5_u1_U54 (.A2( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n121 ) , .A1( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U55 (.A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n153 ) , .A2( u2_u5_u1_n98 ) );
  NAND2_X1 u2_u5_u1_U56 (.A2( u2_u5_u1_n104 ) , .A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n133 ) );
  NAND2_X1 u2_u5_u1_U57 (.ZN( u2_u5_u1_n150 ) , .A2( u2_u5_u1_n98 ) , .A1( u2_u5_u1_n99 ) );
  NAND2_X1 u2_u5_u1_U58 (.A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n155 ) , .A2( u2_u5_u1_n95 ) );
  OAI21_X1 u2_u5_u1_U59 (.ZN( u2_u5_u1_n109 ) , .B1( u2_u5_u1_n129 ) , .B2( u2_u5_u1_n160 ) , .A( u2_u5_u1_n167 ) );
  AOI22_X1 u2_u5_u1_U6 (.B2( u2_u5_u1_n136 ) , .A2( u2_u5_u1_n137 ) , .ZN( u2_u5_u1_n143 ) , .A1( u2_u5_u1_n171 ) , .B1( u2_u5_u1_n173 ) );
  NAND2_X1 u2_u5_u1_U60 (.A2( u2_u5_u1_n100 ) , .A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n120 ) );
  NAND2_X1 u2_u5_u1_U61 (.A1( u2_u5_u1_n102 ) , .A2( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n115 ) );
  NAND2_X1 u2_u5_u1_U62 (.A2( u2_u5_u1_n100 ) , .A1( u2_u5_u1_n104 ) , .ZN( u2_u5_u1_n151 ) );
  NAND2_X1 u2_u5_u1_U63 (.A2( u2_u5_u1_n103 ) , .A1( u2_u5_u1_n105 ) , .ZN( u2_u5_u1_n161 ) );
  INV_X1 u2_u5_u1_U64 (.A( u2_u5_u1_n152 ) , .ZN( u2_u5_u1_n173 ) );
  INV_X1 u2_u5_u1_U65 (.A( u2_u5_u1_n128 ) , .ZN( u2_u5_u1_n172 ) );
  NAND2_X1 u2_u5_u1_U66 (.A2( u2_u5_u1_n102 ) , .A1( u2_u5_u1_n103 ) , .ZN( u2_u5_u1_n123 ) );
  AOI211_X1 u2_u5_u1_U67 (.B( u2_u5_u1_n162 ) , .A( u2_u5_u1_n163 ) , .C2( u2_u5_u1_n164 ) , .ZN( u2_u5_u1_n165 ) , .C1( u2_u5_u1_n171 ) );
  AOI21_X1 u2_u5_u1_U68 (.A( u2_u5_u1_n160 ) , .B2( u2_u5_u1_n161 ) , .ZN( u2_u5_u1_n162 ) , .B1( u2_u5_u1_n182 ) );
  OR2_X1 u2_u5_u1_U69 (.A2( u2_u5_u1_n157 ) , .A1( u2_u5_u1_n158 ) , .ZN( u2_u5_u1_n163 ) );
  INV_X1 u2_u5_u1_U7 (.A( u2_u5_u1_n147 ) , .ZN( u2_u5_u1_n181 ) );
  NOR2_X1 u2_u5_u1_U70 (.A2( u2_u5_X_7 ) , .A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n95 ) );
  NOR2_X1 u2_u5_u1_U71 (.A1( u2_u5_X_12 ) , .A2( u2_u5_X_9 ) , .ZN( u2_u5_u1_n100 ) );
  NOR2_X1 u2_u5_u1_U72 (.A2( u2_u5_X_8 ) , .A1( u2_u5_u1_n177 ) , .ZN( u2_u5_u1_n99 ) );
  NOR2_X1 u2_u5_u1_U73 (.A2( u2_u5_X_12 ) , .ZN( u2_u5_u1_n102 ) , .A1( u2_u5_u1_n176 ) );
  NOR2_X1 u2_u5_u1_U74 (.A2( u2_u5_X_9 ) , .ZN( u2_u5_u1_n105 ) , .A1( u2_u5_u1_n168 ) );
  NAND2_X1 u2_u5_u1_U75 (.A1( u2_u5_X_10 ) , .ZN( u2_u5_u1_n160 ) , .A2( u2_u5_u1_n169 ) );
  NAND2_X1 u2_u5_u1_U76 (.A2( u2_u5_X_10 ) , .A1( u2_u5_X_11 ) , .ZN( u2_u5_u1_n152 ) );
  NAND2_X1 u2_u5_u1_U77 (.A1( u2_u5_X_11 ) , .ZN( u2_u5_u1_n128 ) , .A2( u2_u5_u1_n170 ) );
  AND2_X1 u2_u5_u1_U78 (.A2( u2_u5_X_7 ) , .A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n104 ) );
  AND2_X1 u2_u5_u1_U79 (.A1( u2_u5_X_8 ) , .ZN( u2_u5_u1_n103 ) , .A2( u2_u5_u1_n177 ) );
  AOI22_X1 u2_u5_u1_U8 (.B2( u2_u5_u1_n113 ) , .A2( u2_u5_u1_n114 ) , .ZN( u2_u5_u1_n125 ) , .A1( u2_u5_u1_n171 ) , .B1( u2_u5_u1_n173 ) );
  INV_X1 u2_u5_u1_U80 (.A( u2_u5_X_10 ) , .ZN( u2_u5_u1_n170 ) );
  INV_X1 u2_u5_u1_U81 (.A( u2_u5_X_9 ) , .ZN( u2_u5_u1_n176 ) );
  INV_X1 u2_u5_u1_U82 (.A( u2_u5_X_11 ) , .ZN( u2_u5_u1_n169 ) );
  INV_X1 u2_u5_u1_U83 (.A( u2_u5_X_12 ) , .ZN( u2_u5_u1_n168 ) );
  INV_X1 u2_u5_u1_U84 (.A( u2_u5_X_7 ) , .ZN( u2_u5_u1_n177 ) );
  NAND4_X1 u2_u5_u1_U85 (.ZN( u2_out5_28 ) , .A4( u2_u5_u1_n124 ) , .A3( u2_u5_u1_n125 ) , .A2( u2_u5_u1_n126 ) , .A1( u2_u5_u1_n127 ) );
  OAI21_X1 u2_u5_u1_U86 (.ZN( u2_u5_u1_n127 ) , .B2( u2_u5_u1_n139 ) , .B1( u2_u5_u1_n175 ) , .A( u2_u5_u1_n183 ) );
  OAI21_X1 u2_u5_u1_U87 (.ZN( u2_u5_u1_n126 ) , .B2( u2_u5_u1_n140 ) , .A( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n178 ) );
  NAND4_X1 u2_u5_u1_U88 (.ZN( u2_out5_18 ) , .A4( u2_u5_u1_n165 ) , .A3( u2_u5_u1_n166 ) , .A1( u2_u5_u1_n167 ) , .A2( u2_u5_u1_n186 ) );
  AOI22_X1 u2_u5_u1_U89 (.B2( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n147 ) , .A2( u2_u5_u1_n148 ) , .ZN( u2_u5_u1_n166 ) , .A1( u2_u5_u1_n172 ) );
  NAND2_X1 u2_u5_u1_U9 (.ZN( u2_u5_u1_n114 ) , .A1( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n156 ) );
  INV_X1 u2_u5_u1_U90 (.A( u2_u5_u1_n145 ) , .ZN( u2_u5_u1_n186 ) );
  NAND4_X1 u2_u5_u1_U91 (.ZN( u2_out5_2 ) , .A4( u2_u5_u1_n142 ) , .A3( u2_u5_u1_n143 ) , .A2( u2_u5_u1_n144 ) , .A1( u2_u5_u1_n179 ) );
  OAI21_X1 u2_u5_u1_U92 (.B2( u2_u5_u1_n132 ) , .ZN( u2_u5_u1_n144 ) , .A( u2_u5_u1_n146 ) , .B1( u2_u5_u1_n180 ) );
  INV_X1 u2_u5_u1_U93 (.A( u2_u5_u1_n130 ) , .ZN( u2_u5_u1_n179 ) );
  OR4_X1 u2_u5_u1_U94 (.ZN( u2_out5_13 ) , .A4( u2_u5_u1_n108 ) , .A3( u2_u5_u1_n109 ) , .A2( u2_u5_u1_n110 ) , .A1( u2_u5_u1_n111 ) );
  AOI21_X1 u2_u5_u1_U95 (.ZN( u2_u5_u1_n110 ) , .A( u2_u5_u1_n116 ) , .B1( u2_u5_u1_n152 ) , .B2( u2_u5_u1_n160 ) );
  AOI21_X1 u2_u5_u1_U96 (.ZN( u2_u5_u1_n111 ) , .A( u2_u5_u1_n128 ) , .B2( u2_u5_u1_n131 ) , .B1( u2_u5_u1_n135 ) );
  NAND3_X1 u2_u5_u1_U97 (.A3( u2_u5_u1_n149 ) , .A2( u2_u5_u1_n150 ) , .A1( u2_u5_u1_n151 ) , .ZN( u2_u5_u1_n164 ) );
  NAND3_X1 u2_u5_u1_U98 (.A3( u2_u5_u1_n134 ) , .A2( u2_u5_u1_n135 ) , .ZN( u2_u5_u1_n136 ) , .A1( u2_u5_u1_n151 ) );
  NAND3_X1 u2_u5_u1_U99 (.A1( u2_u5_u1_n133 ) , .ZN( u2_u5_u1_n137 ) , .A2( u2_u5_u1_n154 ) , .A3( u2_u5_u1_n181 ) );
  INV_X1 u2_u5_u5_U10 (.A( u2_u5_u5_n121 ) , .ZN( u2_u5_u5_n177 ) );
  NOR3_X1 u2_u5_u5_U100 (.A3( u2_u5_u5_n141 ) , .A1( u2_u5_u5_n142 ) , .ZN( u2_u5_u5_n143 ) , .A2( u2_u5_u5_n191 ) );
  NAND4_X1 u2_u5_u5_U101 (.ZN( u2_out5_4 ) , .A4( u2_u5_u5_n112 ) , .A2( u2_u5_u5_n113 ) , .A1( u2_u5_u5_n114 ) , .A3( u2_u5_u5_n195 ) );
  AOI211_X1 u2_u5_u5_U102 (.A( u2_u5_u5_n110 ) , .C1( u2_u5_u5_n111 ) , .ZN( u2_u5_u5_n112 ) , .B( u2_u5_u5_n118 ) , .C2( u2_u5_u5_n177 ) );
  AOI222_X1 u2_u5_u5_U103 (.ZN( u2_u5_u5_n113 ) , .A1( u2_u5_u5_n131 ) , .C1( u2_u5_u5_n148 ) , .B2( u2_u5_u5_n174 ) , .C2( u2_u5_u5_n178 ) , .A2( u2_u5_u5_n179 ) , .B1( u2_u5_u5_n99 ) );
  NAND3_X1 u2_u5_u5_U104 (.A2( u2_u5_u5_n154 ) , .A3( u2_u5_u5_n158 ) , .A1( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n99 ) );
  NOR2_X1 u2_u5_u5_U11 (.ZN( u2_u5_u5_n160 ) , .A2( u2_u5_u5_n173 ) , .A1( u2_u5_u5_n177 ) );
  INV_X1 u2_u5_u5_U12 (.A( u2_u5_u5_n150 ) , .ZN( u2_u5_u5_n174 ) );
  AOI21_X1 u2_u5_u5_U13 (.A( u2_u5_u5_n160 ) , .B2( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n162 ) , .B1( u2_u5_u5_n192 ) );
  INV_X1 u2_u5_u5_U14 (.A( u2_u5_u5_n159 ) , .ZN( u2_u5_u5_n192 ) );
  AOI21_X1 u2_u5_u5_U15 (.A( u2_u5_u5_n156 ) , .B2( u2_u5_u5_n157 ) , .B1( u2_u5_u5_n158 ) , .ZN( u2_u5_u5_n163 ) );
  AOI21_X1 u2_u5_u5_U16 (.B2( u2_u5_u5_n139 ) , .B1( u2_u5_u5_n140 ) , .ZN( u2_u5_u5_n141 ) , .A( u2_u5_u5_n150 ) );
  OAI21_X1 u2_u5_u5_U17 (.A( u2_u5_u5_n133 ) , .B2( u2_u5_u5_n134 ) , .B1( u2_u5_u5_n135 ) , .ZN( u2_u5_u5_n142 ) );
  OAI21_X1 u2_u5_u5_U18 (.ZN( u2_u5_u5_n133 ) , .B2( u2_u5_u5_n147 ) , .A( u2_u5_u5_n173 ) , .B1( u2_u5_u5_n188 ) );
  NAND2_X1 u2_u5_u5_U19 (.A2( u2_u5_u5_n119 ) , .A1( u2_u5_u5_n123 ) , .ZN( u2_u5_u5_n137 ) );
  INV_X1 u2_u5_u5_U20 (.A( u2_u5_u5_n155 ) , .ZN( u2_u5_u5_n194 ) );
  NAND2_X1 u2_u5_u5_U21 (.A1( u2_u5_u5_n121 ) , .ZN( u2_u5_u5_n132 ) , .A2( u2_u5_u5_n172 ) );
  NAND2_X1 u2_u5_u5_U22 (.A2( u2_u5_u5_n122 ) , .ZN( u2_u5_u5_n136 ) , .A1( u2_u5_u5_n154 ) );
  NAND2_X1 u2_u5_u5_U23 (.A2( u2_u5_u5_n119 ) , .A1( u2_u5_u5_n120 ) , .ZN( u2_u5_u5_n159 ) );
  INV_X1 u2_u5_u5_U24 (.A( u2_u5_u5_n156 ) , .ZN( u2_u5_u5_n175 ) );
  INV_X1 u2_u5_u5_U25 (.A( u2_u5_u5_n158 ) , .ZN( u2_u5_u5_n188 ) );
  INV_X1 u2_u5_u5_U26 (.A( u2_u5_u5_n152 ) , .ZN( u2_u5_u5_n179 ) );
  INV_X1 u2_u5_u5_U27 (.A( u2_u5_u5_n140 ) , .ZN( u2_u5_u5_n182 ) );
  INV_X1 u2_u5_u5_U28 (.A( u2_u5_u5_n151 ) , .ZN( u2_u5_u5_n183 ) );
  INV_X1 u2_u5_u5_U29 (.A( u2_u5_u5_n123 ) , .ZN( u2_u5_u5_n185 ) );
  NOR2_X1 u2_u5_u5_U3 (.ZN( u2_u5_u5_n134 ) , .A1( u2_u5_u5_n183 ) , .A2( u2_u5_u5_n190 ) );
  INV_X1 u2_u5_u5_U30 (.A( u2_u5_u5_n161 ) , .ZN( u2_u5_u5_n184 ) );
  INV_X1 u2_u5_u5_U31 (.A( u2_u5_u5_n139 ) , .ZN( u2_u5_u5_n189 ) );
  INV_X1 u2_u5_u5_U32 (.A( u2_u5_u5_n157 ) , .ZN( u2_u5_u5_n190 ) );
  INV_X1 u2_u5_u5_U33 (.A( u2_u5_u5_n120 ) , .ZN( u2_u5_u5_n193 ) );
  NAND2_X1 u2_u5_u5_U34 (.ZN( u2_u5_u5_n111 ) , .A1( u2_u5_u5_n140 ) , .A2( u2_u5_u5_n155 ) );
  NOR2_X1 u2_u5_u5_U35 (.ZN( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n170 ) , .A2( u2_u5_u5_n180 ) );
  INV_X1 u2_u5_u5_U36 (.A( u2_u5_u5_n117 ) , .ZN( u2_u5_u5_n196 ) );
  OAI221_X1 u2_u5_u5_U37 (.A( u2_u5_u5_n116 ) , .ZN( u2_u5_u5_n117 ) , .B2( u2_u5_u5_n119 ) , .C1( u2_u5_u5_n153 ) , .C2( u2_u5_u5_n158 ) , .B1( u2_u5_u5_n172 ) );
  AOI222_X1 u2_u5_u5_U38 (.ZN( u2_u5_u5_n116 ) , .B2( u2_u5_u5_n145 ) , .C1( u2_u5_u5_n148 ) , .A2( u2_u5_u5_n174 ) , .C2( u2_u5_u5_n177 ) , .B1( u2_u5_u5_n187 ) , .A1( u2_u5_u5_n193 ) );
  INV_X1 u2_u5_u5_U39 (.A( u2_u5_u5_n115 ) , .ZN( u2_u5_u5_n187 ) );
  INV_X1 u2_u5_u5_U4 (.A( u2_u5_u5_n138 ) , .ZN( u2_u5_u5_n191 ) );
  AOI22_X1 u2_u5_u5_U40 (.B2( u2_u5_u5_n131 ) , .A2( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n169 ) , .B1( u2_u5_u5_n174 ) , .A1( u2_u5_u5_n185 ) );
  NOR2_X1 u2_u5_u5_U41 (.A1( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n150 ) , .A2( u2_u5_u5_n173 ) );
  AOI21_X1 u2_u5_u5_U42 (.A( u2_u5_u5_n118 ) , .B2( u2_u5_u5_n145 ) , .ZN( u2_u5_u5_n168 ) , .B1( u2_u5_u5_n186 ) );
  INV_X1 u2_u5_u5_U43 (.A( u2_u5_u5_n122 ) , .ZN( u2_u5_u5_n186 ) );
  NOR2_X1 u2_u5_u5_U44 (.A1( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n152 ) , .A2( u2_u5_u5_n176 ) );
  NOR2_X1 u2_u5_u5_U45 (.A1( u2_u5_u5_n115 ) , .ZN( u2_u5_u5_n118 ) , .A2( u2_u5_u5_n153 ) );
  NOR2_X1 u2_u5_u5_U46 (.A2( u2_u5_u5_n145 ) , .ZN( u2_u5_u5_n156 ) , .A1( u2_u5_u5_n174 ) );
  NOR2_X1 u2_u5_u5_U47 (.ZN( u2_u5_u5_n121 ) , .A2( u2_u5_u5_n145 ) , .A1( u2_u5_u5_n176 ) );
  AOI22_X1 u2_u5_u5_U48 (.ZN( u2_u5_u5_n114 ) , .A2( u2_u5_u5_n137 ) , .A1( u2_u5_u5_n145 ) , .B2( u2_u5_u5_n175 ) , .B1( u2_u5_u5_n193 ) );
  OAI211_X1 u2_u5_u5_U49 (.B( u2_u5_u5_n124 ) , .A( u2_u5_u5_n125 ) , .C2( u2_u5_u5_n126 ) , .C1( u2_u5_u5_n127 ) , .ZN( u2_u5_u5_n128 ) );
  OAI21_X1 u2_u5_u5_U5 (.B2( u2_u5_u5_n136 ) , .B1( u2_u5_u5_n137 ) , .ZN( u2_u5_u5_n138 ) , .A( u2_u5_u5_n177 ) );
  NOR3_X1 u2_u5_u5_U50 (.ZN( u2_u5_u5_n127 ) , .A1( u2_u5_u5_n136 ) , .A3( u2_u5_u5_n148 ) , .A2( u2_u5_u5_n182 ) );
  OAI21_X1 u2_u5_u5_U51 (.ZN( u2_u5_u5_n124 ) , .A( u2_u5_u5_n177 ) , .B2( u2_u5_u5_n183 ) , .B1( u2_u5_u5_n189 ) );
  OAI21_X1 u2_u5_u5_U52 (.ZN( u2_u5_u5_n125 ) , .A( u2_u5_u5_n174 ) , .B2( u2_u5_u5_n185 ) , .B1( u2_u5_u5_n190 ) );
  AOI21_X1 u2_u5_u5_U53 (.A( u2_u5_u5_n153 ) , .B2( u2_u5_u5_n154 ) , .B1( u2_u5_u5_n155 ) , .ZN( u2_u5_u5_n164 ) );
  AOI21_X1 u2_u5_u5_U54 (.ZN( u2_u5_u5_n110 ) , .B1( u2_u5_u5_n122 ) , .B2( u2_u5_u5_n139 ) , .A( u2_u5_u5_n153 ) );
  INV_X1 u2_u5_u5_U55 (.A( u2_u5_u5_n153 ) , .ZN( u2_u5_u5_n176 ) );
  INV_X1 u2_u5_u5_U56 (.A( u2_u5_u5_n126 ) , .ZN( u2_u5_u5_n173 ) );
  AND2_X1 u2_u5_u5_U57 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n147 ) );
  AND2_X1 u2_u5_u5_U58 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n148 ) );
  NAND2_X1 u2_u5_u5_U59 (.A1( u2_u5_u5_n105 ) , .A2( u2_u5_u5_n106 ) , .ZN( u2_u5_u5_n158 ) );
  INV_X1 u2_u5_u5_U6 (.A( u2_u5_u5_n135 ) , .ZN( u2_u5_u5_n178 ) );
  NAND2_X1 u2_u5_u5_U60 (.A2( u2_u5_u5_n108 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n139 ) );
  NAND2_X1 u2_u5_u5_U61 (.A1( u2_u5_u5_n106 ) , .A2( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n119 ) );
  NAND2_X1 u2_u5_u5_U62 (.A2( u2_u5_u5_n103 ) , .A1( u2_u5_u5_n105 ) , .ZN( u2_u5_u5_n140 ) );
  NAND2_X1 u2_u5_u5_U63 (.A2( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n105 ) , .ZN( u2_u5_u5_n155 ) );
  NAND2_X1 u2_u5_u5_U64 (.A2( u2_u5_u5_n106 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n122 ) );
  NAND2_X1 u2_u5_u5_U65 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n106 ) , .ZN( u2_u5_u5_n115 ) );
  NAND2_X1 u2_u5_u5_U66 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n103 ) , .ZN( u2_u5_u5_n161 ) );
  NAND2_X1 u2_u5_u5_U67 (.A1( u2_u5_u5_n105 ) , .A2( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n154 ) );
  INV_X1 u2_u5_u5_U68 (.A( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n172 ) );
  NAND2_X1 u2_u5_u5_U69 (.A1( u2_u5_u5_n103 ) , .A2( u2_u5_u5_n108 ) , .ZN( u2_u5_u5_n123 ) );
  OAI22_X1 u2_u5_u5_U7 (.B2( u2_u5_u5_n149 ) , .B1( u2_u5_u5_n150 ) , .A2( u2_u5_u5_n151 ) , .A1( u2_u5_u5_n152 ) , .ZN( u2_u5_u5_n165 ) );
  NAND2_X1 u2_u5_u5_U70 (.A2( u2_u5_u5_n103 ) , .A1( u2_u5_u5_n107 ) , .ZN( u2_u5_u5_n151 ) );
  NAND2_X1 u2_u5_u5_U71 (.A2( u2_u5_u5_n107 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n120 ) );
  NAND2_X1 u2_u5_u5_U72 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n109 ) , .ZN( u2_u5_u5_n157 ) );
  AND2_X1 u2_u5_u5_U73 (.A2( u2_u5_u5_n100 ) , .A1( u2_u5_u5_n104 ) , .ZN( u2_u5_u5_n131 ) );
  INV_X1 u2_u5_u5_U74 (.A( u2_u5_u5_n102 ) , .ZN( u2_u5_u5_n195 ) );
  OAI221_X1 u2_u5_u5_U75 (.A( u2_u5_u5_n101 ) , .ZN( u2_u5_u5_n102 ) , .C2( u2_u5_u5_n115 ) , .C1( u2_u5_u5_n126 ) , .B1( u2_u5_u5_n134 ) , .B2( u2_u5_u5_n160 ) );
  OAI21_X1 u2_u5_u5_U76 (.ZN( u2_u5_u5_n101 ) , .B1( u2_u5_u5_n137 ) , .A( u2_u5_u5_n146 ) , .B2( u2_u5_u5_n147 ) );
  NOR2_X1 u2_u5_u5_U77 (.A2( u2_u5_X_34 ) , .A1( u2_u5_X_35 ) , .ZN( u2_u5_u5_n145 ) );
  NOR2_X1 u2_u5_u5_U78 (.A2( u2_u5_X_34 ) , .ZN( u2_u5_u5_n146 ) , .A1( u2_u5_u5_n171 ) );
  NOR2_X1 u2_u5_u5_U79 (.A2( u2_u5_X_31 ) , .A1( u2_u5_X_32 ) , .ZN( u2_u5_u5_n103 ) );
  NOR3_X1 u2_u5_u5_U8 (.A2( u2_u5_u5_n147 ) , .A1( u2_u5_u5_n148 ) , .ZN( u2_u5_u5_n149 ) , .A3( u2_u5_u5_n194 ) );
  NOR2_X1 u2_u5_u5_U80 (.A2( u2_u5_X_36 ) , .ZN( u2_u5_u5_n105 ) , .A1( u2_u5_u5_n180 ) );
  NOR2_X1 u2_u5_u5_U81 (.A2( u2_u5_X_33 ) , .ZN( u2_u5_u5_n108 ) , .A1( u2_u5_u5_n170 ) );
  NOR2_X1 u2_u5_u5_U82 (.A2( u2_u5_X_33 ) , .A1( u2_u5_X_36 ) , .ZN( u2_u5_u5_n107 ) );
  NOR2_X1 u2_u5_u5_U83 (.A2( u2_u5_X_31 ) , .ZN( u2_u5_u5_n104 ) , .A1( u2_u5_u5_n181 ) );
  NAND2_X1 u2_u5_u5_U84 (.A2( u2_u5_X_34 ) , .A1( u2_u5_X_35 ) , .ZN( u2_u5_u5_n153 ) );
  NAND2_X1 u2_u5_u5_U85 (.A1( u2_u5_X_34 ) , .ZN( u2_u5_u5_n126 ) , .A2( u2_u5_u5_n171 ) );
  AND2_X1 u2_u5_u5_U86 (.A1( u2_u5_X_31 ) , .A2( u2_u5_X_32 ) , .ZN( u2_u5_u5_n106 ) );
  AND2_X1 u2_u5_u5_U87 (.A1( u2_u5_X_31 ) , .ZN( u2_u5_u5_n109 ) , .A2( u2_u5_u5_n181 ) );
  INV_X1 u2_u5_u5_U88 (.A( u2_u5_X_33 ) , .ZN( u2_u5_u5_n180 ) );
  INV_X1 u2_u5_u5_U89 (.A( u2_u5_X_35 ) , .ZN( u2_u5_u5_n171 ) );
  NOR2_X1 u2_u5_u5_U9 (.ZN( u2_u5_u5_n135 ) , .A1( u2_u5_u5_n173 ) , .A2( u2_u5_u5_n176 ) );
  INV_X1 u2_u5_u5_U90 (.A( u2_u5_X_36 ) , .ZN( u2_u5_u5_n170 ) );
  INV_X1 u2_u5_u5_U91 (.A( u2_u5_X_32 ) , .ZN( u2_u5_u5_n181 ) );
  NAND4_X1 u2_u5_u5_U92 (.ZN( u2_out5_29 ) , .A4( u2_u5_u5_n129 ) , .A3( u2_u5_u5_n130 ) , .A2( u2_u5_u5_n168 ) , .A1( u2_u5_u5_n196 ) );
  AOI221_X1 u2_u5_u5_U93 (.A( u2_u5_u5_n128 ) , .ZN( u2_u5_u5_n129 ) , .C2( u2_u5_u5_n132 ) , .B2( u2_u5_u5_n159 ) , .B1( u2_u5_u5_n176 ) , .C1( u2_u5_u5_n184 ) );
  AOI222_X1 u2_u5_u5_U94 (.ZN( u2_u5_u5_n130 ) , .A2( u2_u5_u5_n146 ) , .B1( u2_u5_u5_n147 ) , .C2( u2_u5_u5_n175 ) , .B2( u2_u5_u5_n179 ) , .A1( u2_u5_u5_n188 ) , .C1( u2_u5_u5_n194 ) );
  NAND4_X1 u2_u5_u5_U95 (.ZN( u2_out5_19 ) , .A4( u2_u5_u5_n166 ) , .A3( u2_u5_u5_n167 ) , .A2( u2_u5_u5_n168 ) , .A1( u2_u5_u5_n169 ) );
  AOI22_X1 u2_u5_u5_U96 (.B2( u2_u5_u5_n145 ) , .A2( u2_u5_u5_n146 ) , .ZN( u2_u5_u5_n167 ) , .B1( u2_u5_u5_n182 ) , .A1( u2_u5_u5_n189 ) );
  NOR4_X1 u2_u5_u5_U97 (.A4( u2_u5_u5_n162 ) , .A3( u2_u5_u5_n163 ) , .A2( u2_u5_u5_n164 ) , .A1( u2_u5_u5_n165 ) , .ZN( u2_u5_u5_n166 ) );
  NAND4_X1 u2_u5_u5_U98 (.ZN( u2_out5_11 ) , .A4( u2_u5_u5_n143 ) , .A3( u2_u5_u5_n144 ) , .A2( u2_u5_u5_n169 ) , .A1( u2_u5_u5_n196 ) );
  AOI22_X1 u2_u5_u5_U99 (.A2( u2_u5_u5_n132 ) , .ZN( u2_u5_u5_n144 ) , .B2( u2_u5_u5_n145 ) , .B1( u2_u5_u5_n184 ) , .A1( u2_u5_u5_n194 ) );
  OAI21_X1 u2_u5_u6_U10 (.A( u2_u5_u6_n159 ) , .B1( u2_u5_u6_n169 ) , .B2( u2_u5_u6_n173 ) , .ZN( u2_u5_u6_n90 ) );
  INV_X1 u2_u5_u6_U11 (.ZN( u2_u5_u6_n172 ) , .A( u2_u5_u6_n88 ) );
  AOI22_X1 u2_u5_u6_U12 (.A2( u2_u5_u6_n151 ) , .B2( u2_u5_u6_n161 ) , .A1( u2_u5_u6_n167 ) , .B1( u2_u5_u6_n170 ) , .ZN( u2_u5_u6_n89 ) );
  AOI21_X1 u2_u5_u6_U13 (.ZN( u2_u5_u6_n106 ) , .A( u2_u5_u6_n142 ) , .B2( u2_u5_u6_n159 ) , .B1( u2_u5_u6_n164 ) );
  INV_X1 u2_u5_u6_U14 (.A( u2_u5_u6_n155 ) , .ZN( u2_u5_u6_n161 ) );
  INV_X1 u2_u5_u6_U15 (.A( u2_u5_u6_n128 ) , .ZN( u2_u5_u6_n164 ) );
  NAND2_X1 u2_u5_u6_U16 (.ZN( u2_u5_u6_n110 ) , .A1( u2_u5_u6_n122 ) , .A2( u2_u5_u6_n129 ) );
  NAND2_X1 u2_u5_u6_U17 (.ZN( u2_u5_u6_n124 ) , .A2( u2_u5_u6_n146 ) , .A1( u2_u5_u6_n148 ) );
  INV_X1 u2_u5_u6_U18 (.A( u2_u5_u6_n132 ) , .ZN( u2_u5_u6_n171 ) );
  AND2_X1 u2_u5_u6_U19 (.A1( u2_u5_u6_n100 ) , .ZN( u2_u5_u6_n130 ) , .A2( u2_u5_u6_n147 ) );
  INV_X1 u2_u5_u6_U20 (.A( u2_u5_u6_n127 ) , .ZN( u2_u5_u6_n173 ) );
  INV_X1 u2_u5_u6_U21 (.A( u2_u5_u6_n121 ) , .ZN( u2_u5_u6_n167 ) );
  INV_X1 u2_u5_u6_U22 (.A( u2_u5_u6_n100 ) , .ZN( u2_u5_u6_n169 ) );
  INV_X1 u2_u5_u6_U23 (.A( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n170 ) );
  INV_X1 u2_u5_u6_U24 (.A( u2_u5_u6_n113 ) , .ZN( u2_u5_u6_n168 ) );
  AND2_X1 u2_u5_u6_U25 (.A1( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n119 ) , .ZN( u2_u5_u6_n133 ) );
  AND2_X1 u2_u5_u6_U26 (.A2( u2_u5_u6_n121 ) , .A1( u2_u5_u6_n122 ) , .ZN( u2_u5_u6_n131 ) );
  AND3_X1 u2_u5_u6_U27 (.ZN( u2_u5_u6_n120 ) , .A2( u2_u5_u6_n127 ) , .A1( u2_u5_u6_n132 ) , .A3( u2_u5_u6_n145 ) );
  INV_X1 u2_u5_u6_U28 (.A( u2_u5_u6_n146 ) , .ZN( u2_u5_u6_n163 ) );
  AOI222_X1 u2_u5_u6_U29 (.ZN( u2_u5_u6_n114 ) , .A1( u2_u5_u6_n118 ) , .A2( u2_u5_u6_n126 ) , .B2( u2_u5_u6_n151 ) , .C2( u2_u5_u6_n159 ) , .C1( u2_u5_u6_n168 ) , .B1( u2_u5_u6_n169 ) );
  INV_X1 u2_u5_u6_U3 (.A( u2_u5_u6_n110 ) , .ZN( u2_u5_u6_n166 ) );
  NOR2_X1 u2_u5_u6_U30 (.A1( u2_u5_u6_n162 ) , .A2( u2_u5_u6_n165 ) , .ZN( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U31 (.A1( u2_u5_u6_n144 ) , .ZN( u2_u5_u6_n151 ) , .A2( u2_u5_u6_n158 ) );
  NAND2_X1 u2_u5_u6_U32 (.ZN( u2_u5_u6_n132 ) , .A1( u2_u5_u6_n91 ) , .A2( u2_u5_u6_n97 ) );
  NOR2_X1 u2_u5_u6_U33 (.A2( u2_u5_u6_n126 ) , .ZN( u2_u5_u6_n155 ) , .A1( u2_u5_u6_n160 ) );
  NAND2_X1 u2_u5_u6_U34 (.ZN( u2_u5_u6_n146 ) , .A2( u2_u5_u6_n94 ) , .A1( u2_u5_u6_n99 ) );
  AOI21_X1 u2_u5_u6_U35 (.A( u2_u5_u6_n144 ) , .B2( u2_u5_u6_n145 ) , .B1( u2_u5_u6_n146 ) , .ZN( u2_u5_u6_n150 ) );
  INV_X1 u2_u5_u6_U36 (.A( u2_u5_u6_n111 ) , .ZN( u2_u5_u6_n158 ) );
  NAND2_X1 u2_u5_u6_U37 (.ZN( u2_u5_u6_n127 ) , .A1( u2_u5_u6_n91 ) , .A2( u2_u5_u6_n92 ) );
  NAND2_X1 u2_u5_u6_U38 (.ZN( u2_u5_u6_n129 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n96 ) );
  INV_X1 u2_u5_u6_U39 (.A( u2_u5_u6_n144 ) , .ZN( u2_u5_u6_n159 ) );
  INV_X1 u2_u5_u6_U4 (.A( u2_u5_u6_n142 ) , .ZN( u2_u5_u6_n174 ) );
  NAND2_X1 u2_u5_u6_U40 (.ZN( u2_u5_u6_n145 ) , .A2( u2_u5_u6_n97 ) , .A1( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U41 (.ZN( u2_u5_u6_n148 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n94 ) );
  NAND2_X1 u2_u5_u6_U42 (.ZN( u2_u5_u6_n108 ) , .A2( u2_u5_u6_n139 ) , .A1( u2_u5_u6_n144 ) );
  NAND2_X1 u2_u5_u6_U43 (.ZN( u2_u5_u6_n121 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n97 ) );
  NAND2_X1 u2_u5_u6_U44 (.ZN( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n95 ) );
  AND2_X1 u2_u5_u6_U45 (.ZN( u2_u5_u6_n118 ) , .A2( u2_u5_u6_n91 ) , .A1( u2_u5_u6_n99 ) );
  AOI22_X1 u2_u5_u6_U46 (.B2( u2_u5_u6_n110 ) , .B1( u2_u5_u6_n111 ) , .A1( u2_u5_u6_n112 ) , .ZN( u2_u5_u6_n115 ) , .A2( u2_u5_u6_n161 ) );
  NAND4_X1 u2_u5_u6_U47 (.A3( u2_u5_u6_n109 ) , .ZN( u2_u5_u6_n112 ) , .A4( u2_u5_u6_n132 ) , .A2( u2_u5_u6_n147 ) , .A1( u2_u5_u6_n166 ) );
  NOR2_X1 u2_u5_u6_U48 (.ZN( u2_u5_u6_n109 ) , .A1( u2_u5_u6_n170 ) , .A2( u2_u5_u6_n173 ) );
  NAND2_X1 u2_u5_u6_U49 (.ZN( u2_u5_u6_n147 ) , .A2( u2_u5_u6_n98 ) , .A1( u2_u5_u6_n99 ) );
  NAND2_X1 u2_u5_u6_U5 (.A2( u2_u5_u6_n143 ) , .ZN( u2_u5_u6_n152 ) , .A1( u2_u5_u6_n166 ) );
  NAND2_X1 u2_u5_u6_U50 (.ZN( u2_u5_u6_n128 ) , .A1( u2_u5_u6_n94 ) , .A2( u2_u5_u6_n96 ) );
  AOI211_X1 u2_u5_u6_U51 (.B( u2_u5_u6_n134 ) , .A( u2_u5_u6_n135 ) , .C1( u2_u5_u6_n136 ) , .ZN( u2_u5_u6_n137 ) , .C2( u2_u5_u6_n151 ) );
  AOI21_X1 u2_u5_u6_U52 (.B2( u2_u5_u6_n132 ) , .B1( u2_u5_u6_n133 ) , .ZN( u2_u5_u6_n134 ) , .A( u2_u5_u6_n158 ) );
  AOI21_X1 u2_u5_u6_U53 (.B1( u2_u5_u6_n131 ) , .ZN( u2_u5_u6_n135 ) , .A( u2_u5_u6_n144 ) , .B2( u2_u5_u6_n146 ) );
  NAND4_X1 u2_u5_u6_U54 (.A4( u2_u5_u6_n127 ) , .A3( u2_u5_u6_n128 ) , .A2( u2_u5_u6_n129 ) , .A1( u2_u5_u6_n130 ) , .ZN( u2_u5_u6_n136 ) );
  NAND2_X1 u2_u5_u6_U55 (.ZN( u2_u5_u6_n119 ) , .A2( u2_u5_u6_n95 ) , .A1( u2_u5_u6_n99 ) );
  NAND2_X1 u2_u5_u6_U56 (.ZN( u2_u5_u6_n123 ) , .A2( u2_u5_u6_n91 ) , .A1( u2_u5_u6_n96 ) );
  NAND2_X1 u2_u5_u6_U57 (.ZN( u2_u5_u6_n100 ) , .A2( u2_u5_u6_n92 ) , .A1( u2_u5_u6_n98 ) );
  NAND2_X1 u2_u5_u6_U58 (.ZN( u2_u5_u6_n122 ) , .A1( u2_u5_u6_n94 ) , .A2( u2_u5_u6_n97 ) );
  INV_X1 u2_u5_u6_U59 (.A( u2_u5_u6_n139 ) , .ZN( u2_u5_u6_n160 ) );
  AOI22_X1 u2_u5_u6_U6 (.B2( u2_u5_u6_n101 ) , .A1( u2_u5_u6_n102 ) , .ZN( u2_u5_u6_n103 ) , .B1( u2_u5_u6_n160 ) , .A2( u2_u5_u6_n161 ) );
  NAND2_X1 u2_u5_u6_U60 (.ZN( u2_u5_u6_n113 ) , .A1( u2_u5_u6_n96 ) , .A2( u2_u5_u6_n98 ) );
  NOR2_X1 u2_u5_u6_U61 (.A2( u2_u5_X_40 ) , .A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n126 ) );
  NOR2_X1 u2_u5_u6_U62 (.A2( u2_u5_X_39 ) , .A1( u2_u5_X_42 ) , .ZN( u2_u5_u6_n92 ) );
  NOR2_X1 u2_u5_u6_U63 (.A2( u2_u5_X_39 ) , .A1( u2_u5_u6_n156 ) , .ZN( u2_u5_u6_n97 ) );
  NOR2_X1 u2_u5_u6_U64 (.A2( u2_u5_X_38 ) , .A1( u2_u5_u6_n165 ) , .ZN( u2_u5_u6_n95 ) );
  NOR2_X1 u2_u5_u6_U65 (.A2( u2_u5_X_41 ) , .ZN( u2_u5_u6_n111 ) , .A1( u2_u5_u6_n157 ) );
  NOR2_X1 u2_u5_u6_U66 (.A2( u2_u5_X_37 ) , .A1( u2_u5_u6_n162 ) , .ZN( u2_u5_u6_n94 ) );
  NOR2_X1 u2_u5_u6_U67 (.A2( u2_u5_X_37 ) , .A1( u2_u5_X_38 ) , .ZN( u2_u5_u6_n91 ) );
  NAND2_X1 u2_u5_u6_U68 (.A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n144 ) , .A2( u2_u5_u6_n157 ) );
  NAND2_X1 u2_u5_u6_U69 (.A2( u2_u5_X_40 ) , .A1( u2_u5_X_41 ) , .ZN( u2_u5_u6_n139 ) );
  NOR2_X1 u2_u5_u6_U7 (.A1( u2_u5_u6_n118 ) , .ZN( u2_u5_u6_n143 ) , .A2( u2_u5_u6_n168 ) );
  AND2_X1 u2_u5_u6_U70 (.A1( u2_u5_X_39 ) , .A2( u2_u5_u6_n156 ) , .ZN( u2_u5_u6_n96 ) );
  AND2_X1 u2_u5_u6_U71 (.A1( u2_u5_X_39 ) , .A2( u2_u5_X_42 ) , .ZN( u2_u5_u6_n99 ) );
  INV_X1 u2_u5_u6_U72 (.A( u2_u5_X_40 ) , .ZN( u2_u5_u6_n157 ) );
  INV_X1 u2_u5_u6_U73 (.A( u2_u5_X_37 ) , .ZN( u2_u5_u6_n165 ) );
  INV_X1 u2_u5_u6_U74 (.A( u2_u5_X_38 ) , .ZN( u2_u5_u6_n162 ) );
  INV_X1 u2_u5_u6_U75 (.A( u2_u5_X_42 ) , .ZN( u2_u5_u6_n156 ) );
  NAND4_X1 u2_u5_u6_U76 (.ZN( u2_out5_32 ) , .A4( u2_u5_u6_n103 ) , .A3( u2_u5_u6_n104 ) , .A2( u2_u5_u6_n105 ) , .A1( u2_u5_u6_n106 ) );
  AOI22_X1 u2_u5_u6_U77 (.ZN( u2_u5_u6_n105 ) , .A2( u2_u5_u6_n108 ) , .A1( u2_u5_u6_n118 ) , .B2( u2_u5_u6_n126 ) , .B1( u2_u5_u6_n171 ) );
  AOI22_X1 u2_u5_u6_U78 (.ZN( u2_u5_u6_n104 ) , .A1( u2_u5_u6_n111 ) , .B1( u2_u5_u6_n124 ) , .B2( u2_u5_u6_n151 ) , .A2( u2_u5_u6_n93 ) );
  NAND4_X1 u2_u5_u6_U79 (.ZN( u2_out5_12 ) , .A4( u2_u5_u6_n114 ) , .A3( u2_u5_u6_n115 ) , .A2( u2_u5_u6_n116 ) , .A1( u2_u5_u6_n117 ) );
  AOI21_X1 u2_u5_u6_U8 (.B1( u2_u5_u6_n107 ) , .B2( u2_u5_u6_n132 ) , .A( u2_u5_u6_n158 ) , .ZN( u2_u5_u6_n88 ) );
  OAI22_X1 u2_u5_u6_U80 (.B2( u2_u5_u6_n111 ) , .ZN( u2_u5_u6_n116 ) , .B1( u2_u5_u6_n126 ) , .A2( u2_u5_u6_n164 ) , .A1( u2_u5_u6_n167 ) );
  OAI21_X1 u2_u5_u6_U81 (.A( u2_u5_u6_n108 ) , .ZN( u2_u5_u6_n117 ) , .B2( u2_u5_u6_n141 ) , .B1( u2_u5_u6_n163 ) );
  OAI211_X1 u2_u5_u6_U82 (.ZN( u2_out5_22 ) , .B( u2_u5_u6_n137 ) , .A( u2_u5_u6_n138 ) , .C2( u2_u5_u6_n139 ) , .C1( u2_u5_u6_n140 ) );
  AOI22_X1 u2_u5_u6_U83 (.B1( u2_u5_u6_n124 ) , .A2( u2_u5_u6_n125 ) , .A1( u2_u5_u6_n126 ) , .ZN( u2_u5_u6_n138 ) , .B2( u2_u5_u6_n161 ) );
  AND4_X1 u2_u5_u6_U84 (.A3( u2_u5_u6_n119 ) , .A1( u2_u5_u6_n120 ) , .A4( u2_u5_u6_n129 ) , .ZN( u2_u5_u6_n140 ) , .A2( u2_u5_u6_n143 ) );
  OAI211_X1 u2_u5_u6_U85 (.ZN( u2_out5_7 ) , .B( u2_u5_u6_n153 ) , .C2( u2_u5_u6_n154 ) , .C1( u2_u5_u6_n155 ) , .A( u2_u5_u6_n174 ) );
  NOR3_X1 u2_u5_u6_U86 (.A1( u2_u5_u6_n141 ) , .ZN( u2_u5_u6_n154 ) , .A3( u2_u5_u6_n164 ) , .A2( u2_u5_u6_n171 ) );
  AOI211_X1 u2_u5_u6_U87 (.B( u2_u5_u6_n149 ) , .A( u2_u5_u6_n150 ) , .C2( u2_u5_u6_n151 ) , .C1( u2_u5_u6_n152 ) , .ZN( u2_u5_u6_n153 ) );
  NAND3_X1 u2_u5_u6_U88 (.A2( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n125 ) , .A1( u2_u5_u6_n130 ) , .A3( u2_u5_u6_n131 ) );
  NAND3_X1 u2_u5_u6_U89 (.A3( u2_u5_u6_n133 ) , .ZN( u2_u5_u6_n141 ) , .A1( u2_u5_u6_n145 ) , .A2( u2_u5_u6_n148 ) );
  AOI21_X1 u2_u5_u6_U9 (.B2( u2_u5_u6_n147 ) , .B1( u2_u5_u6_n148 ) , .ZN( u2_u5_u6_n149 ) , .A( u2_u5_u6_n158 ) );
  NAND3_X1 u2_u5_u6_U90 (.ZN( u2_u5_u6_n101 ) , .A3( u2_u5_u6_n107 ) , .A2( u2_u5_u6_n121 ) , .A1( u2_u5_u6_n127 ) );
  NAND3_X1 u2_u5_u6_U91 (.ZN( u2_u5_u6_n102 ) , .A3( u2_u5_u6_n130 ) , .A2( u2_u5_u6_n145 ) , .A1( u2_u5_u6_n166 ) );
  NAND3_X1 u2_u5_u6_U92 (.A3( u2_u5_u6_n113 ) , .A1( u2_u5_u6_n119 ) , .A2( u2_u5_u6_n123 ) , .ZN( u2_u5_u6_n93 ) );
  NAND3_X1 u2_u5_u6_U93 (.ZN( u2_u5_u6_n142 ) , .A2( u2_u5_u6_n172 ) , .A3( u2_u5_u6_n89 ) , .A1( u2_u5_u6_n90 ) );
  AND3_X1 u2_u5_u7_U10 (.A3( u2_u5_u7_n110 ) , .A2( u2_u5_u7_n127 ) , .A1( u2_u5_u7_n132 ) , .ZN( u2_u5_u7_n92 ) );
  OAI21_X1 u2_u5_u7_U11 (.A( u2_u5_u7_n161 ) , .B1( u2_u5_u7_n168 ) , .B2( u2_u5_u7_n173 ) , .ZN( u2_u5_u7_n91 ) );
  AOI211_X1 u2_u5_u7_U12 (.A( u2_u5_u7_n117 ) , .ZN( u2_u5_u7_n118 ) , .C2( u2_u5_u7_n126 ) , .C1( u2_u5_u7_n177 ) , .B( u2_u5_u7_n180 ) );
  OAI22_X1 u2_u5_u7_U13 (.B1( u2_u5_u7_n115 ) , .ZN( u2_u5_u7_n117 ) , .A2( u2_u5_u7_n133 ) , .A1( u2_u5_u7_n137 ) , .B2( u2_u5_u7_n162 ) );
  INV_X1 u2_u5_u7_U14 (.A( u2_u5_u7_n116 ) , .ZN( u2_u5_u7_n180 ) );
  NOR3_X1 u2_u5_u7_U15 (.ZN( u2_u5_u7_n115 ) , .A3( u2_u5_u7_n145 ) , .A2( u2_u5_u7_n168 ) , .A1( u2_u5_u7_n169 ) );
  OAI211_X1 u2_u5_u7_U16 (.B( u2_u5_u7_n122 ) , .A( u2_u5_u7_n123 ) , .C2( u2_u5_u7_n124 ) , .ZN( u2_u5_u7_n154 ) , .C1( u2_u5_u7_n162 ) );
  AOI222_X1 u2_u5_u7_U17 (.ZN( u2_u5_u7_n122 ) , .C2( u2_u5_u7_n126 ) , .C1( u2_u5_u7_n145 ) , .B1( u2_u5_u7_n161 ) , .A2( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n170 ) , .A1( u2_u5_u7_n176 ) );
  INV_X1 u2_u5_u7_U18 (.A( u2_u5_u7_n133 ) , .ZN( u2_u5_u7_n176 ) );
  NOR3_X1 u2_u5_u7_U19 (.A2( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n135 ) , .ZN( u2_u5_u7_n136 ) , .A3( u2_u5_u7_n171 ) );
  NOR2_X1 u2_u5_u7_U20 (.A1( u2_u5_u7_n130 ) , .A2( u2_u5_u7_n134 ) , .ZN( u2_u5_u7_n153 ) );
  INV_X1 u2_u5_u7_U21 (.A( u2_u5_u7_n101 ) , .ZN( u2_u5_u7_n165 ) );
  NOR2_X1 u2_u5_u7_U22 (.ZN( u2_u5_u7_n111 ) , .A2( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n169 ) );
  AOI21_X1 u2_u5_u7_U23 (.ZN( u2_u5_u7_n104 ) , .B2( u2_u5_u7_n112 ) , .B1( u2_u5_u7_n127 ) , .A( u2_u5_u7_n164 ) );
  AOI21_X1 u2_u5_u7_U24 (.ZN( u2_u5_u7_n106 ) , .B1( u2_u5_u7_n133 ) , .B2( u2_u5_u7_n146 ) , .A( u2_u5_u7_n162 ) );
  AOI21_X1 u2_u5_u7_U25 (.A( u2_u5_u7_n101 ) , .ZN( u2_u5_u7_n107 ) , .B2( u2_u5_u7_n128 ) , .B1( u2_u5_u7_n175 ) );
  INV_X1 u2_u5_u7_U26 (.A( u2_u5_u7_n138 ) , .ZN( u2_u5_u7_n171 ) );
  INV_X1 u2_u5_u7_U27 (.A( u2_u5_u7_n131 ) , .ZN( u2_u5_u7_n177 ) );
  INV_X1 u2_u5_u7_U28 (.A( u2_u5_u7_n110 ) , .ZN( u2_u5_u7_n174 ) );
  NAND2_X1 u2_u5_u7_U29 (.A1( u2_u5_u7_n129 ) , .A2( u2_u5_u7_n132 ) , .ZN( u2_u5_u7_n149 ) );
  OAI21_X1 u2_u5_u7_U3 (.ZN( u2_u5_u7_n159 ) , .A( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n171 ) , .B1( u2_u5_u7_n174 ) );
  NAND2_X1 u2_u5_u7_U30 (.A1( u2_u5_u7_n113 ) , .A2( u2_u5_u7_n124 ) , .ZN( u2_u5_u7_n130 ) );
  INV_X1 u2_u5_u7_U31 (.A( u2_u5_u7_n112 ) , .ZN( u2_u5_u7_n173 ) );
  INV_X1 u2_u5_u7_U32 (.A( u2_u5_u7_n128 ) , .ZN( u2_u5_u7_n168 ) );
  INV_X1 u2_u5_u7_U33 (.A( u2_u5_u7_n148 ) , .ZN( u2_u5_u7_n169 ) );
  INV_X1 u2_u5_u7_U34 (.A( u2_u5_u7_n127 ) , .ZN( u2_u5_u7_n179 ) );
  NOR2_X1 u2_u5_u7_U35 (.ZN( u2_u5_u7_n101 ) , .A2( u2_u5_u7_n150 ) , .A1( u2_u5_u7_n156 ) );
  AOI211_X1 u2_u5_u7_U36 (.B( u2_u5_u7_n154 ) , .A( u2_u5_u7_n155 ) , .C1( u2_u5_u7_n156 ) , .ZN( u2_u5_u7_n157 ) , .C2( u2_u5_u7_n172 ) );
  INV_X1 u2_u5_u7_U37 (.A( u2_u5_u7_n153 ) , .ZN( u2_u5_u7_n172 ) );
  AOI211_X1 u2_u5_u7_U38 (.B( u2_u5_u7_n139 ) , .A( u2_u5_u7_n140 ) , .C2( u2_u5_u7_n141 ) , .ZN( u2_u5_u7_n142 ) , .C1( u2_u5_u7_n156 ) );
  NAND4_X1 u2_u5_u7_U39 (.A3( u2_u5_u7_n127 ) , .A2( u2_u5_u7_n128 ) , .A1( u2_u5_u7_n129 ) , .ZN( u2_u5_u7_n141 ) , .A4( u2_u5_u7_n147 ) );
  INV_X1 u2_u5_u7_U4 (.A( u2_u5_u7_n111 ) , .ZN( u2_u5_u7_n170 ) );
  AOI21_X1 u2_u5_u7_U40 (.A( u2_u5_u7_n137 ) , .B1( u2_u5_u7_n138 ) , .ZN( u2_u5_u7_n139 ) , .B2( u2_u5_u7_n146 ) );
  OAI22_X1 u2_u5_u7_U41 (.B1( u2_u5_u7_n136 ) , .ZN( u2_u5_u7_n140 ) , .A1( u2_u5_u7_n153 ) , .B2( u2_u5_u7_n162 ) , .A2( u2_u5_u7_n164 ) );
  AOI21_X1 u2_u5_u7_U42 (.ZN( u2_u5_u7_n123 ) , .B1( u2_u5_u7_n165 ) , .B2( u2_u5_u7_n177 ) , .A( u2_u5_u7_n97 ) );
  AOI21_X1 u2_u5_u7_U43 (.B2( u2_u5_u7_n113 ) , .B1( u2_u5_u7_n124 ) , .A( u2_u5_u7_n125 ) , .ZN( u2_u5_u7_n97 ) );
  INV_X1 u2_u5_u7_U44 (.A( u2_u5_u7_n125 ) , .ZN( u2_u5_u7_n161 ) );
  INV_X1 u2_u5_u7_U45 (.A( u2_u5_u7_n152 ) , .ZN( u2_u5_u7_n162 ) );
  AOI22_X1 u2_u5_u7_U46 (.A2( u2_u5_u7_n114 ) , .ZN( u2_u5_u7_n119 ) , .B1( u2_u5_u7_n130 ) , .A1( u2_u5_u7_n156 ) , .B2( u2_u5_u7_n165 ) );
  NAND2_X1 u2_u5_u7_U47 (.A2( u2_u5_u7_n112 ) , .ZN( u2_u5_u7_n114 ) , .A1( u2_u5_u7_n175 ) );
  AND2_X1 u2_u5_u7_U48 (.ZN( u2_u5_u7_n145 ) , .A2( u2_u5_u7_n98 ) , .A1( u2_u5_u7_n99 ) );
  NOR2_X1 u2_u5_u7_U49 (.ZN( u2_u5_u7_n137 ) , .A1( u2_u5_u7_n150 ) , .A2( u2_u5_u7_n161 ) );
  INV_X1 u2_u5_u7_U5 (.A( u2_u5_u7_n149 ) , .ZN( u2_u5_u7_n175 ) );
  AOI21_X1 u2_u5_u7_U50 (.ZN( u2_u5_u7_n105 ) , .B2( u2_u5_u7_n110 ) , .A( u2_u5_u7_n125 ) , .B1( u2_u5_u7_n147 ) );
  NAND2_X1 u2_u5_u7_U51 (.ZN( u2_u5_u7_n146 ) , .A1( u2_u5_u7_n95 ) , .A2( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U52 (.A2( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n147 ) , .A1( u2_u5_u7_n93 ) );
  NAND2_X1 u2_u5_u7_U53 (.A1( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n127 ) , .A2( u2_u5_u7_n99 ) );
  OR2_X1 u2_u5_u7_U54 (.ZN( u2_u5_u7_n126 ) , .A2( u2_u5_u7_n152 ) , .A1( u2_u5_u7_n156 ) );
  NAND2_X1 u2_u5_u7_U55 (.A2( u2_u5_u7_n102 ) , .A1( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n133 ) );
  NAND2_X1 u2_u5_u7_U56 (.ZN( u2_u5_u7_n112 ) , .A2( u2_u5_u7_n96 ) , .A1( u2_u5_u7_n99 ) );
  NAND2_X1 u2_u5_u7_U57 (.A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n128 ) , .A1( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U58 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n113 ) , .A2( u2_u5_u7_n93 ) );
  NAND2_X1 u2_u5_u7_U59 (.A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n124 ) , .A1( u2_u5_u7_n96 ) );
  INV_X1 u2_u5_u7_U6 (.A( u2_u5_u7_n154 ) , .ZN( u2_u5_u7_n178 ) );
  NAND2_X1 u2_u5_u7_U60 (.ZN( u2_u5_u7_n110 ) , .A1( u2_u5_u7_n95 ) , .A2( u2_u5_u7_n96 ) );
  INV_X1 u2_u5_u7_U61 (.A( u2_u5_u7_n150 ) , .ZN( u2_u5_u7_n164 ) );
  AND2_X1 u2_u5_u7_U62 (.ZN( u2_u5_u7_n134 ) , .A1( u2_u5_u7_n93 ) , .A2( u2_u5_u7_n98 ) );
  NAND2_X1 u2_u5_u7_U63 (.A1( u2_u5_u7_n100 ) , .A2( u2_u5_u7_n102 ) , .ZN( u2_u5_u7_n129 ) );
  NAND2_X1 u2_u5_u7_U64 (.A2( u2_u5_u7_n103 ) , .ZN( u2_u5_u7_n131 ) , .A1( u2_u5_u7_n95 ) );
  NAND2_X1 u2_u5_u7_U65 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n138 ) , .A2( u2_u5_u7_n99 ) );
  NAND2_X1 u2_u5_u7_U66 (.ZN( u2_u5_u7_n132 ) , .A1( u2_u5_u7_n93 ) , .A2( u2_u5_u7_n96 ) );
  NAND2_X1 u2_u5_u7_U67 (.A1( u2_u5_u7_n100 ) , .ZN( u2_u5_u7_n148 ) , .A2( u2_u5_u7_n95 ) );
  NOR2_X1 u2_u5_u7_U68 (.A2( u2_u5_X_47 ) , .ZN( u2_u5_u7_n150 ) , .A1( u2_u5_u7_n163 ) );
  NOR2_X1 u2_u5_u7_U69 (.A2( u2_u5_X_43 ) , .A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n103 ) );
  AOI211_X1 u2_u5_u7_U7 (.ZN( u2_u5_u7_n116 ) , .A( u2_u5_u7_n155 ) , .C1( u2_u5_u7_n161 ) , .C2( u2_u5_u7_n171 ) , .B( u2_u5_u7_n94 ) );
  NOR2_X1 u2_u5_u7_U70 (.A2( u2_u5_X_48 ) , .A1( u2_u5_u7_n166 ) , .ZN( u2_u5_u7_n95 ) );
  NOR2_X1 u2_u5_u7_U71 (.A2( u2_u5_X_45 ) , .A1( u2_u5_X_48 ) , .ZN( u2_u5_u7_n99 ) );
  NOR2_X1 u2_u5_u7_U72 (.A2( u2_u5_X_44 ) , .A1( u2_u5_u7_n167 ) , .ZN( u2_u5_u7_n98 ) );
  NOR2_X1 u2_u5_u7_U73 (.A2( u2_u5_X_46 ) , .A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n152 ) );
  AND2_X1 u2_u5_u7_U74 (.A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n156 ) , .A2( u2_u5_u7_n163 ) );
  NAND2_X1 u2_u5_u7_U75 (.A2( u2_u5_X_46 ) , .A1( u2_u5_X_47 ) , .ZN( u2_u5_u7_n125 ) );
  AND2_X1 u2_u5_u7_U76 (.A2( u2_u5_X_45 ) , .A1( u2_u5_X_48 ) , .ZN( u2_u5_u7_n102 ) );
  AND2_X1 u2_u5_u7_U77 (.A2( u2_u5_X_43 ) , .A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n96 ) );
  AND2_X1 u2_u5_u7_U78 (.A1( u2_u5_X_44 ) , .ZN( u2_u5_u7_n100 ) , .A2( u2_u5_u7_n167 ) );
  AND2_X1 u2_u5_u7_U79 (.A1( u2_u5_X_48 ) , .A2( u2_u5_u7_n166 ) , .ZN( u2_u5_u7_n93 ) );
  OAI222_X1 u2_u5_u7_U8 (.C2( u2_u5_u7_n101 ) , .B2( u2_u5_u7_n111 ) , .A1( u2_u5_u7_n113 ) , .C1( u2_u5_u7_n146 ) , .A2( u2_u5_u7_n162 ) , .B1( u2_u5_u7_n164 ) , .ZN( u2_u5_u7_n94 ) );
  INV_X1 u2_u5_u7_U80 (.A( u2_u5_X_46 ) , .ZN( u2_u5_u7_n163 ) );
  INV_X1 u2_u5_u7_U81 (.A( u2_u5_X_43 ) , .ZN( u2_u5_u7_n167 ) );
  INV_X1 u2_u5_u7_U82 (.A( u2_u5_X_45 ) , .ZN( u2_u5_u7_n166 ) );
  NAND4_X1 u2_u5_u7_U83 (.ZN( u2_out5_27 ) , .A4( u2_u5_u7_n118 ) , .A3( u2_u5_u7_n119 ) , .A2( u2_u5_u7_n120 ) , .A1( u2_u5_u7_n121 ) );
  OAI21_X1 u2_u5_u7_U84 (.ZN( u2_u5_u7_n121 ) , .B2( u2_u5_u7_n145 ) , .A( u2_u5_u7_n150 ) , .B1( u2_u5_u7_n174 ) );
  OAI21_X1 u2_u5_u7_U85 (.ZN( u2_u5_u7_n120 ) , .A( u2_u5_u7_n161 ) , .B2( u2_u5_u7_n170 ) , .B1( u2_u5_u7_n179 ) );
  NAND4_X1 u2_u5_u7_U86 (.ZN( u2_out5_21 ) , .A4( u2_u5_u7_n157 ) , .A3( u2_u5_u7_n158 ) , .A2( u2_u5_u7_n159 ) , .A1( u2_u5_u7_n160 ) );
  OAI21_X1 u2_u5_u7_U87 (.B1( u2_u5_u7_n145 ) , .ZN( u2_u5_u7_n160 ) , .A( u2_u5_u7_n161 ) , .B2( u2_u5_u7_n177 ) );
  AOI22_X1 u2_u5_u7_U88 (.B2( u2_u5_u7_n149 ) , .B1( u2_u5_u7_n150 ) , .A2( u2_u5_u7_n151 ) , .A1( u2_u5_u7_n152 ) , .ZN( u2_u5_u7_n158 ) );
  NAND4_X1 u2_u5_u7_U89 (.ZN( u2_out5_15 ) , .A4( u2_u5_u7_n142 ) , .A3( u2_u5_u7_n143 ) , .A2( u2_u5_u7_n144 ) , .A1( u2_u5_u7_n178 ) );
  OAI221_X1 u2_u5_u7_U9 (.C1( u2_u5_u7_n101 ) , .C2( u2_u5_u7_n147 ) , .ZN( u2_u5_u7_n155 ) , .B2( u2_u5_u7_n162 ) , .A( u2_u5_u7_n91 ) , .B1( u2_u5_u7_n92 ) );
  OR2_X1 u2_u5_u7_U90 (.A2( u2_u5_u7_n125 ) , .A1( u2_u5_u7_n129 ) , .ZN( u2_u5_u7_n144 ) );
  AOI22_X1 u2_u5_u7_U91 (.A2( u2_u5_u7_n126 ) , .ZN( u2_u5_u7_n143 ) , .B2( u2_u5_u7_n165 ) , .B1( u2_u5_u7_n173 ) , .A1( u2_u5_u7_n174 ) );
  NAND4_X1 u2_u5_u7_U92 (.ZN( u2_out5_5 ) , .A4( u2_u5_u7_n108 ) , .A3( u2_u5_u7_n109 ) , .A1( u2_u5_u7_n116 ) , .A2( u2_u5_u7_n123 ) );
  AOI22_X1 u2_u5_u7_U93 (.ZN( u2_u5_u7_n109 ) , .A2( u2_u5_u7_n126 ) , .B2( u2_u5_u7_n145 ) , .B1( u2_u5_u7_n156 ) , .A1( u2_u5_u7_n171 ) );
  NOR4_X1 u2_u5_u7_U94 (.A4( u2_u5_u7_n104 ) , .A3( u2_u5_u7_n105 ) , .A2( u2_u5_u7_n106 ) , .A1( u2_u5_u7_n107 ) , .ZN( u2_u5_u7_n108 ) );
  NAND3_X1 u2_u5_u7_U95 (.A3( u2_u5_u7_n146 ) , .A2( u2_u5_u7_n147 ) , .A1( u2_u5_u7_n148 ) , .ZN( u2_u5_u7_n151 ) );
  NAND3_X1 u2_u5_u7_U96 (.A3( u2_u5_u7_n131 ) , .A2( u2_u5_u7_n132 ) , .A1( u2_u5_u7_n133 ) , .ZN( u2_u5_u7_n135 ) );
  XOR2_X1 u2_u6_U20 (.B( u2_K7_36 ) , .A( u2_R5_25 ) , .Z( u2_u6_X_36 ) );
  XOR2_X1 u2_u6_U21 (.B( u2_K7_35 ) , .A( u2_R5_24 ) , .Z( u2_u6_X_35 ) );
  XOR2_X1 u2_u6_U22 (.B( u2_K7_34 ) , .A( u2_R5_23 ) , .Z( u2_u6_X_34 ) );
  XOR2_X1 u2_u6_U23 (.B( u2_K7_33 ) , .A( u2_R5_22 ) , .Z( u2_u6_X_33 ) );
  XOR2_X1 u2_u6_U24 (.B( u2_K7_32 ) , .A( u2_R5_21 ) , .Z( u2_u6_X_32 ) );
  XOR2_X1 u2_u6_U25 (.B( u2_K7_31 ) , .A( u2_R5_20 ) , .Z( u2_u6_X_31 ) );
  INV_X1 u2_u6_u5_U10 (.A( u2_u6_u5_n121 ) , .ZN( u2_u6_u5_n177 ) );
  NOR3_X1 u2_u6_u5_U100 (.A3( u2_u6_u5_n141 ) , .A1( u2_u6_u5_n142 ) , .ZN( u2_u6_u5_n143 ) , .A2( u2_u6_u5_n191 ) );
  NAND4_X1 u2_u6_u5_U101 (.ZN( u2_out6_4 ) , .A4( u2_u6_u5_n112 ) , .A2( u2_u6_u5_n113 ) , .A1( u2_u6_u5_n114 ) , .A3( u2_u6_u5_n195 ) );
  AOI211_X1 u2_u6_u5_U102 (.A( u2_u6_u5_n110 ) , .C1( u2_u6_u5_n111 ) , .ZN( u2_u6_u5_n112 ) , .B( u2_u6_u5_n118 ) , .C2( u2_u6_u5_n177 ) );
  AOI222_X1 u2_u6_u5_U103 (.ZN( u2_u6_u5_n113 ) , .A1( u2_u6_u5_n131 ) , .C1( u2_u6_u5_n148 ) , .B2( u2_u6_u5_n174 ) , .C2( u2_u6_u5_n178 ) , .A2( u2_u6_u5_n179 ) , .B1( u2_u6_u5_n99 ) );
  NAND3_X1 u2_u6_u5_U104 (.A2( u2_u6_u5_n154 ) , .A3( u2_u6_u5_n158 ) , .A1( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n99 ) );
  NOR2_X1 u2_u6_u5_U11 (.ZN( u2_u6_u5_n160 ) , .A2( u2_u6_u5_n173 ) , .A1( u2_u6_u5_n177 ) );
  INV_X1 u2_u6_u5_U12 (.A( u2_u6_u5_n150 ) , .ZN( u2_u6_u5_n174 ) );
  AOI21_X1 u2_u6_u5_U13 (.A( u2_u6_u5_n160 ) , .B2( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n162 ) , .B1( u2_u6_u5_n192 ) );
  INV_X1 u2_u6_u5_U14 (.A( u2_u6_u5_n159 ) , .ZN( u2_u6_u5_n192 ) );
  AOI21_X1 u2_u6_u5_U15 (.A( u2_u6_u5_n156 ) , .B2( u2_u6_u5_n157 ) , .B1( u2_u6_u5_n158 ) , .ZN( u2_u6_u5_n163 ) );
  AOI21_X1 u2_u6_u5_U16 (.B2( u2_u6_u5_n139 ) , .B1( u2_u6_u5_n140 ) , .ZN( u2_u6_u5_n141 ) , .A( u2_u6_u5_n150 ) );
  OAI21_X1 u2_u6_u5_U17 (.A( u2_u6_u5_n133 ) , .B2( u2_u6_u5_n134 ) , .B1( u2_u6_u5_n135 ) , .ZN( u2_u6_u5_n142 ) );
  OAI21_X1 u2_u6_u5_U18 (.ZN( u2_u6_u5_n133 ) , .B2( u2_u6_u5_n147 ) , .A( u2_u6_u5_n173 ) , .B1( u2_u6_u5_n188 ) );
  NAND2_X1 u2_u6_u5_U19 (.A2( u2_u6_u5_n119 ) , .A1( u2_u6_u5_n123 ) , .ZN( u2_u6_u5_n137 ) );
  INV_X1 u2_u6_u5_U20 (.A( u2_u6_u5_n155 ) , .ZN( u2_u6_u5_n194 ) );
  NAND2_X1 u2_u6_u5_U21 (.A1( u2_u6_u5_n121 ) , .ZN( u2_u6_u5_n132 ) , .A2( u2_u6_u5_n172 ) );
  NAND2_X1 u2_u6_u5_U22 (.A2( u2_u6_u5_n122 ) , .ZN( u2_u6_u5_n136 ) , .A1( u2_u6_u5_n154 ) );
  NAND2_X1 u2_u6_u5_U23 (.A2( u2_u6_u5_n119 ) , .A1( u2_u6_u5_n120 ) , .ZN( u2_u6_u5_n159 ) );
  INV_X1 u2_u6_u5_U24 (.A( u2_u6_u5_n156 ) , .ZN( u2_u6_u5_n175 ) );
  INV_X1 u2_u6_u5_U25 (.A( u2_u6_u5_n158 ) , .ZN( u2_u6_u5_n188 ) );
  INV_X1 u2_u6_u5_U26 (.A( u2_u6_u5_n152 ) , .ZN( u2_u6_u5_n179 ) );
  INV_X1 u2_u6_u5_U27 (.A( u2_u6_u5_n140 ) , .ZN( u2_u6_u5_n182 ) );
  INV_X1 u2_u6_u5_U28 (.A( u2_u6_u5_n151 ) , .ZN( u2_u6_u5_n183 ) );
  INV_X1 u2_u6_u5_U29 (.A( u2_u6_u5_n123 ) , .ZN( u2_u6_u5_n185 ) );
  NOR2_X1 u2_u6_u5_U3 (.ZN( u2_u6_u5_n134 ) , .A1( u2_u6_u5_n183 ) , .A2( u2_u6_u5_n190 ) );
  INV_X1 u2_u6_u5_U30 (.A( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n184 ) );
  INV_X1 u2_u6_u5_U31 (.A( u2_u6_u5_n139 ) , .ZN( u2_u6_u5_n189 ) );
  INV_X1 u2_u6_u5_U32 (.A( u2_u6_u5_n157 ) , .ZN( u2_u6_u5_n190 ) );
  INV_X1 u2_u6_u5_U33 (.A( u2_u6_u5_n120 ) , .ZN( u2_u6_u5_n193 ) );
  NAND2_X1 u2_u6_u5_U34 (.ZN( u2_u6_u5_n111 ) , .A1( u2_u6_u5_n140 ) , .A2( u2_u6_u5_n155 ) );
  INV_X1 u2_u6_u5_U35 (.A( u2_u6_u5_n117 ) , .ZN( u2_u6_u5_n196 ) );
  OAI221_X1 u2_u6_u5_U36 (.A( u2_u6_u5_n116 ) , .ZN( u2_u6_u5_n117 ) , .B2( u2_u6_u5_n119 ) , .C1( u2_u6_u5_n153 ) , .C2( u2_u6_u5_n158 ) , .B1( u2_u6_u5_n172 ) );
  AOI222_X1 u2_u6_u5_U37 (.ZN( u2_u6_u5_n116 ) , .B2( u2_u6_u5_n145 ) , .C1( u2_u6_u5_n148 ) , .A2( u2_u6_u5_n174 ) , .C2( u2_u6_u5_n177 ) , .B1( u2_u6_u5_n187 ) , .A1( u2_u6_u5_n193 ) );
  INV_X1 u2_u6_u5_U38 (.A( u2_u6_u5_n115 ) , .ZN( u2_u6_u5_n187 ) );
  NOR2_X1 u2_u6_u5_U39 (.ZN( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n170 ) , .A2( u2_u6_u5_n180 ) );
  INV_X1 u2_u6_u5_U4 (.A( u2_u6_u5_n138 ) , .ZN( u2_u6_u5_n191 ) );
  AOI22_X1 u2_u6_u5_U40 (.B2( u2_u6_u5_n131 ) , .A2( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n169 ) , .B1( u2_u6_u5_n174 ) , .A1( u2_u6_u5_n185 ) );
  NOR2_X1 u2_u6_u5_U41 (.A1( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n150 ) , .A2( u2_u6_u5_n173 ) );
  AOI21_X1 u2_u6_u5_U42 (.A( u2_u6_u5_n118 ) , .B2( u2_u6_u5_n145 ) , .ZN( u2_u6_u5_n168 ) , .B1( u2_u6_u5_n186 ) );
  INV_X1 u2_u6_u5_U43 (.A( u2_u6_u5_n122 ) , .ZN( u2_u6_u5_n186 ) );
  NOR2_X1 u2_u6_u5_U44 (.A1( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n152 ) , .A2( u2_u6_u5_n176 ) );
  NOR2_X1 u2_u6_u5_U45 (.A1( u2_u6_u5_n115 ) , .ZN( u2_u6_u5_n118 ) , .A2( u2_u6_u5_n153 ) );
  NOR2_X1 u2_u6_u5_U46 (.A2( u2_u6_u5_n145 ) , .ZN( u2_u6_u5_n156 ) , .A1( u2_u6_u5_n174 ) );
  NOR2_X1 u2_u6_u5_U47 (.ZN( u2_u6_u5_n121 ) , .A2( u2_u6_u5_n145 ) , .A1( u2_u6_u5_n176 ) );
  AOI22_X1 u2_u6_u5_U48 (.ZN( u2_u6_u5_n114 ) , .A2( u2_u6_u5_n137 ) , .A1( u2_u6_u5_n145 ) , .B2( u2_u6_u5_n175 ) , .B1( u2_u6_u5_n193 ) );
  OAI211_X1 u2_u6_u5_U49 (.B( u2_u6_u5_n124 ) , .A( u2_u6_u5_n125 ) , .C2( u2_u6_u5_n126 ) , .C1( u2_u6_u5_n127 ) , .ZN( u2_u6_u5_n128 ) );
  OAI21_X1 u2_u6_u5_U5 (.B2( u2_u6_u5_n136 ) , .B1( u2_u6_u5_n137 ) , .ZN( u2_u6_u5_n138 ) , .A( u2_u6_u5_n177 ) );
  NOR3_X1 u2_u6_u5_U50 (.ZN( u2_u6_u5_n127 ) , .A1( u2_u6_u5_n136 ) , .A3( u2_u6_u5_n148 ) , .A2( u2_u6_u5_n182 ) );
  OAI21_X1 u2_u6_u5_U51 (.ZN( u2_u6_u5_n124 ) , .A( u2_u6_u5_n177 ) , .B2( u2_u6_u5_n183 ) , .B1( u2_u6_u5_n189 ) );
  OAI21_X1 u2_u6_u5_U52 (.ZN( u2_u6_u5_n125 ) , .A( u2_u6_u5_n174 ) , .B2( u2_u6_u5_n185 ) , .B1( u2_u6_u5_n190 ) );
  AOI21_X1 u2_u6_u5_U53 (.A( u2_u6_u5_n153 ) , .B2( u2_u6_u5_n154 ) , .B1( u2_u6_u5_n155 ) , .ZN( u2_u6_u5_n164 ) );
  AOI21_X1 u2_u6_u5_U54 (.ZN( u2_u6_u5_n110 ) , .B1( u2_u6_u5_n122 ) , .B2( u2_u6_u5_n139 ) , .A( u2_u6_u5_n153 ) );
  INV_X1 u2_u6_u5_U55 (.A( u2_u6_u5_n153 ) , .ZN( u2_u6_u5_n176 ) );
  INV_X1 u2_u6_u5_U56 (.A( u2_u6_u5_n126 ) , .ZN( u2_u6_u5_n173 ) );
  AND2_X1 u2_u6_u5_U57 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n147 ) );
  AND2_X1 u2_u6_u5_U58 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n148 ) );
  NAND2_X1 u2_u6_u5_U59 (.A1( u2_u6_u5_n105 ) , .A2( u2_u6_u5_n106 ) , .ZN( u2_u6_u5_n158 ) );
  INV_X1 u2_u6_u5_U6 (.A( u2_u6_u5_n135 ) , .ZN( u2_u6_u5_n178 ) );
  NAND2_X1 u2_u6_u5_U60 (.A2( u2_u6_u5_n108 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n139 ) );
  NAND2_X1 u2_u6_u5_U61 (.A1( u2_u6_u5_n106 ) , .A2( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n119 ) );
  NAND2_X1 u2_u6_u5_U62 (.A2( u2_u6_u5_n103 ) , .A1( u2_u6_u5_n105 ) , .ZN( u2_u6_u5_n140 ) );
  NAND2_X1 u2_u6_u5_U63 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n105 ) , .ZN( u2_u6_u5_n155 ) );
  NAND2_X1 u2_u6_u5_U64 (.A2( u2_u6_u5_n106 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n122 ) );
  NAND2_X1 u2_u6_u5_U65 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n106 ) , .ZN( u2_u6_u5_n115 ) );
  NAND2_X1 u2_u6_u5_U66 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n103 ) , .ZN( u2_u6_u5_n161 ) );
  NAND2_X1 u2_u6_u5_U67 (.A1( u2_u6_u5_n105 ) , .A2( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n154 ) );
  INV_X1 u2_u6_u5_U68 (.A( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n172 ) );
  NAND2_X1 u2_u6_u5_U69 (.A1( u2_u6_u5_n103 ) , .A2( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n123 ) );
  OAI22_X1 u2_u6_u5_U7 (.B2( u2_u6_u5_n149 ) , .B1( u2_u6_u5_n150 ) , .A2( u2_u6_u5_n151 ) , .A1( u2_u6_u5_n152 ) , .ZN( u2_u6_u5_n165 ) );
  NAND2_X1 u2_u6_u5_U70 (.A2( u2_u6_u5_n103 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n151 ) );
  NAND2_X1 u2_u6_u5_U71 (.A2( u2_u6_u5_n107 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n120 ) );
  NAND2_X1 u2_u6_u5_U72 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n157 ) );
  AND2_X1 u2_u6_u5_U73 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n104 ) , .ZN( u2_u6_u5_n131 ) );
  INV_X1 u2_u6_u5_U74 (.A( u2_u6_u5_n102 ) , .ZN( u2_u6_u5_n195 ) );
  OAI221_X1 u2_u6_u5_U75 (.A( u2_u6_u5_n101 ) , .ZN( u2_u6_u5_n102 ) , .C2( u2_u6_u5_n115 ) , .C1( u2_u6_u5_n126 ) , .B1( u2_u6_u5_n134 ) , .B2( u2_u6_u5_n160 ) );
  OAI21_X1 u2_u6_u5_U76 (.ZN( u2_u6_u5_n101 ) , .B1( u2_u6_u5_n137 ) , .A( u2_u6_u5_n146 ) , .B2( u2_u6_u5_n147 ) );
  NOR2_X1 u2_u6_u5_U77 (.A2( u2_u6_X_34 ) , .A1( u2_u6_X_35 ) , .ZN( u2_u6_u5_n145 ) );
  NOR2_X1 u2_u6_u5_U78 (.A2( u2_u6_X_34 ) , .ZN( u2_u6_u5_n146 ) , .A1( u2_u6_u5_n171 ) );
  NOR2_X1 u2_u6_u5_U79 (.A2( u2_u6_X_31 ) , .A1( u2_u6_X_32 ) , .ZN( u2_u6_u5_n103 ) );
  NOR3_X1 u2_u6_u5_U8 (.A2( u2_u6_u5_n147 ) , .A1( u2_u6_u5_n148 ) , .ZN( u2_u6_u5_n149 ) , .A3( u2_u6_u5_n194 ) );
  NOR2_X1 u2_u6_u5_U80 (.A2( u2_u6_X_36 ) , .ZN( u2_u6_u5_n105 ) , .A1( u2_u6_u5_n180 ) );
  NOR2_X1 u2_u6_u5_U81 (.A2( u2_u6_X_33 ) , .ZN( u2_u6_u5_n108 ) , .A1( u2_u6_u5_n170 ) );
  NOR2_X1 u2_u6_u5_U82 (.A2( u2_u6_X_33 ) , .A1( u2_u6_X_36 ) , .ZN( u2_u6_u5_n107 ) );
  NOR2_X1 u2_u6_u5_U83 (.A2( u2_u6_X_31 ) , .ZN( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n181 ) );
  NAND2_X1 u2_u6_u5_U84 (.A2( u2_u6_X_34 ) , .A1( u2_u6_X_35 ) , .ZN( u2_u6_u5_n153 ) );
  NAND2_X1 u2_u6_u5_U85 (.A1( u2_u6_X_34 ) , .ZN( u2_u6_u5_n126 ) , .A2( u2_u6_u5_n171 ) );
  AND2_X1 u2_u6_u5_U86 (.A1( u2_u6_X_31 ) , .A2( u2_u6_X_32 ) , .ZN( u2_u6_u5_n106 ) );
  AND2_X1 u2_u6_u5_U87 (.A1( u2_u6_X_31 ) , .ZN( u2_u6_u5_n109 ) , .A2( u2_u6_u5_n181 ) );
  INV_X1 u2_u6_u5_U88 (.A( u2_u6_X_33 ) , .ZN( u2_u6_u5_n180 ) );
  INV_X1 u2_u6_u5_U89 (.A( u2_u6_X_35 ) , .ZN( u2_u6_u5_n171 ) );
  NOR2_X1 u2_u6_u5_U9 (.ZN( u2_u6_u5_n135 ) , .A1( u2_u6_u5_n173 ) , .A2( u2_u6_u5_n176 ) );
  INV_X1 u2_u6_u5_U90 (.A( u2_u6_X_36 ) , .ZN( u2_u6_u5_n170 ) );
  INV_X1 u2_u6_u5_U91 (.A( u2_u6_X_32 ) , .ZN( u2_u6_u5_n181 ) );
  NAND4_X1 u2_u6_u5_U92 (.ZN( u2_out6_29 ) , .A4( u2_u6_u5_n129 ) , .A3( u2_u6_u5_n130 ) , .A2( u2_u6_u5_n168 ) , .A1( u2_u6_u5_n196 ) );
  AOI221_X1 u2_u6_u5_U93 (.A( u2_u6_u5_n128 ) , .ZN( u2_u6_u5_n129 ) , .C2( u2_u6_u5_n132 ) , .B2( u2_u6_u5_n159 ) , .B1( u2_u6_u5_n176 ) , .C1( u2_u6_u5_n184 ) );
  AOI222_X1 u2_u6_u5_U94 (.ZN( u2_u6_u5_n130 ) , .A2( u2_u6_u5_n146 ) , .B1( u2_u6_u5_n147 ) , .C2( u2_u6_u5_n175 ) , .B2( u2_u6_u5_n179 ) , .A1( u2_u6_u5_n188 ) , .C1( u2_u6_u5_n194 ) );
  NAND4_X1 u2_u6_u5_U95 (.ZN( u2_out6_19 ) , .A4( u2_u6_u5_n166 ) , .A3( u2_u6_u5_n167 ) , .A2( u2_u6_u5_n168 ) , .A1( u2_u6_u5_n169 ) );
  AOI22_X1 u2_u6_u5_U96 (.B2( u2_u6_u5_n145 ) , .A2( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n167 ) , .B1( u2_u6_u5_n182 ) , .A1( u2_u6_u5_n189 ) );
  NOR4_X1 u2_u6_u5_U97 (.A4( u2_u6_u5_n162 ) , .A3( u2_u6_u5_n163 ) , .A2( u2_u6_u5_n164 ) , .A1( u2_u6_u5_n165 ) , .ZN( u2_u6_u5_n166 ) );
  NAND4_X1 u2_u6_u5_U98 (.ZN( u2_out6_11 ) , .A4( u2_u6_u5_n143 ) , .A3( u2_u6_u5_n144 ) , .A2( u2_u6_u5_n169 ) , .A1( u2_u6_u5_n196 ) );
  AOI22_X1 u2_u6_u5_U99 (.A2( u2_u6_u5_n132 ) , .ZN( u2_u6_u5_n144 ) , .B2( u2_u6_u5_n145 ) , .B1( u2_u6_u5_n184 ) , .A1( u2_u6_u5_n194 ) );
  XOR2_X1 u2_u7_U20 (.B( u2_K8_36 ) , .A( u2_R6_25 ) , .Z( u2_u7_X_36 ) );
  XOR2_X1 u2_u7_U21 (.B( u2_K8_35 ) , .A( u2_R6_24 ) , .Z( u2_u7_X_35 ) );
  XOR2_X1 u2_u7_U22 (.B( u2_K8_34 ) , .A( u2_R6_23 ) , .Z( u2_u7_X_34 ) );
  XOR2_X1 u2_u7_U23 (.B( u2_K8_33 ) , .A( u2_R6_22 ) , .Z( u2_u7_X_33 ) );
  XOR2_X1 u2_u7_U24 (.B( u2_K8_32 ) , .A( u2_R6_21 ) , .Z( u2_u7_X_32 ) );
  XOR2_X1 u2_u7_U25 (.B( u2_K8_31 ) , .A( u2_R6_20 ) , .Z( u2_u7_X_31 ) );
  XOR2_X1 u2_u7_U26 (.B( u2_K8_30 ) , .A( u2_R6_21 ) , .Z( u2_u7_X_30 ) );
  XOR2_X1 u2_u7_U28 (.B( u2_K8_29 ) , .A( u2_R6_20 ) , .Z( u2_u7_X_29 ) );
  XOR2_X1 u2_u7_U29 (.B( u2_K8_28 ) , .A( u2_R6_19 ) , .Z( u2_u7_X_28 ) );
  XOR2_X1 u2_u7_U30 (.B( u2_K8_27 ) , .A( u2_R6_18 ) , .Z( u2_u7_X_27 ) );
  XOR2_X1 u2_u7_U31 (.B( u2_K8_26 ) , .A( u2_R6_17 ) , .Z( u2_u7_X_26 ) );
  XOR2_X1 u2_u7_U32 (.B( u2_K8_25 ) , .A( u2_R6_16 ) , .Z( u2_u7_X_25 ) );
  OAI22_X1 u2_u7_u4_U10 (.B2( u2_u7_u4_n135 ) , .ZN( u2_u7_u4_n137 ) , .B1( u2_u7_u4_n153 ) , .A1( u2_u7_u4_n155 ) , .A2( u2_u7_u4_n171 ) );
  AND3_X1 u2_u7_u4_U11 (.A2( u2_u7_u4_n134 ) , .ZN( u2_u7_u4_n135 ) , .A3( u2_u7_u4_n145 ) , .A1( u2_u7_u4_n157 ) );
  OR3_X1 u2_u7_u4_U12 (.A3( u2_u7_u4_n114 ) , .A2( u2_u7_u4_n115 ) , .A1( u2_u7_u4_n116 ) , .ZN( u2_u7_u4_n136 ) );
  AOI21_X1 u2_u7_u4_U13 (.A( u2_u7_u4_n113 ) , .ZN( u2_u7_u4_n116 ) , .B2( u2_u7_u4_n173 ) , .B1( u2_u7_u4_n174 ) );
  AOI21_X1 u2_u7_u4_U14 (.ZN( u2_u7_u4_n115 ) , .B2( u2_u7_u4_n145 ) , .B1( u2_u7_u4_n146 ) , .A( u2_u7_u4_n156 ) );
  OAI22_X1 u2_u7_u4_U15 (.ZN( u2_u7_u4_n114 ) , .A2( u2_u7_u4_n121 ) , .B1( u2_u7_u4_n160 ) , .B2( u2_u7_u4_n170 ) , .A1( u2_u7_u4_n171 ) );
  NAND2_X1 u2_u7_u4_U16 (.ZN( u2_u7_u4_n132 ) , .A2( u2_u7_u4_n170 ) , .A1( u2_u7_u4_n173 ) );
  AOI21_X1 u2_u7_u4_U17 (.B2( u2_u7_u4_n160 ) , .B1( u2_u7_u4_n161 ) , .ZN( u2_u7_u4_n162 ) , .A( u2_u7_u4_n170 ) );
  AOI21_X1 u2_u7_u4_U18 (.ZN( u2_u7_u4_n107 ) , .B2( u2_u7_u4_n143 ) , .A( u2_u7_u4_n174 ) , .B1( u2_u7_u4_n184 ) );
  AOI21_X1 u2_u7_u4_U19 (.B2( u2_u7_u4_n158 ) , .B1( u2_u7_u4_n159 ) , .ZN( u2_u7_u4_n163 ) , .A( u2_u7_u4_n174 ) );
  AOI21_X1 u2_u7_u4_U20 (.A( u2_u7_u4_n153 ) , .B2( u2_u7_u4_n154 ) , .B1( u2_u7_u4_n155 ) , .ZN( u2_u7_u4_n165 ) );
  AOI21_X1 u2_u7_u4_U21 (.A( u2_u7_u4_n156 ) , .B2( u2_u7_u4_n157 ) , .ZN( u2_u7_u4_n164 ) , .B1( u2_u7_u4_n184 ) );
  INV_X1 u2_u7_u4_U22 (.A( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n170 ) );
  AND2_X1 u2_u7_u4_U23 (.A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n155 ) , .A1( u2_u7_u4_n160 ) );
  INV_X1 u2_u7_u4_U24 (.A( u2_u7_u4_n156 ) , .ZN( u2_u7_u4_n175 ) );
  NAND2_X1 u2_u7_u4_U25 (.A2( u2_u7_u4_n118 ) , .ZN( u2_u7_u4_n131 ) , .A1( u2_u7_u4_n147 ) );
  NAND2_X1 u2_u7_u4_U26 (.A1( u2_u7_u4_n119 ) , .A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n130 ) );
  NAND2_X1 u2_u7_u4_U27 (.ZN( u2_u7_u4_n117 ) , .A2( u2_u7_u4_n118 ) , .A1( u2_u7_u4_n148 ) );
  NAND2_X1 u2_u7_u4_U28 (.ZN( u2_u7_u4_n129 ) , .A1( u2_u7_u4_n134 ) , .A2( u2_u7_u4_n148 ) );
  AND3_X1 u2_u7_u4_U29 (.A1( u2_u7_u4_n119 ) , .A2( u2_u7_u4_n143 ) , .A3( u2_u7_u4_n154 ) , .ZN( u2_u7_u4_n161 ) );
  NOR2_X1 u2_u7_u4_U3 (.ZN( u2_u7_u4_n121 ) , .A1( u2_u7_u4_n181 ) , .A2( u2_u7_u4_n182 ) );
  AND2_X1 u2_u7_u4_U30 (.A1( u2_u7_u4_n145 ) , .A2( u2_u7_u4_n147 ) , .ZN( u2_u7_u4_n159 ) );
  INV_X1 u2_u7_u4_U31 (.A( u2_u7_u4_n158 ) , .ZN( u2_u7_u4_n182 ) );
  INV_X1 u2_u7_u4_U32 (.ZN( u2_u7_u4_n181 ) , .A( u2_u7_u4_n96 ) );
  INV_X1 u2_u7_u4_U33 (.A( u2_u7_u4_n144 ) , .ZN( u2_u7_u4_n179 ) );
  INV_X1 u2_u7_u4_U34 (.A( u2_u7_u4_n157 ) , .ZN( u2_u7_u4_n178 ) );
  NAND2_X1 u2_u7_u4_U35 (.A2( u2_u7_u4_n154 ) , .A1( u2_u7_u4_n96 ) , .ZN( u2_u7_u4_n97 ) );
  INV_X1 u2_u7_u4_U36 (.ZN( u2_u7_u4_n186 ) , .A( u2_u7_u4_n95 ) );
  OAI221_X1 u2_u7_u4_U37 (.C1( u2_u7_u4_n134 ) , .B1( u2_u7_u4_n158 ) , .B2( u2_u7_u4_n171 ) , .C2( u2_u7_u4_n173 ) , .A( u2_u7_u4_n94 ) , .ZN( u2_u7_u4_n95 ) );
  AOI222_X1 u2_u7_u4_U38 (.B2( u2_u7_u4_n132 ) , .A1( u2_u7_u4_n138 ) , .C2( u2_u7_u4_n175 ) , .A2( u2_u7_u4_n179 ) , .C1( u2_u7_u4_n181 ) , .B1( u2_u7_u4_n185 ) , .ZN( u2_u7_u4_n94 ) );
  INV_X1 u2_u7_u4_U39 (.A( u2_u7_u4_n113 ) , .ZN( u2_u7_u4_n185 ) );
  INV_X1 u2_u7_u4_U4 (.A( u2_u7_u4_n117 ) , .ZN( u2_u7_u4_n184 ) );
  INV_X1 u2_u7_u4_U40 (.A( u2_u7_u4_n143 ) , .ZN( u2_u7_u4_n183 ) );
  NOR2_X1 u2_u7_u4_U41 (.ZN( u2_u7_u4_n138 ) , .A1( u2_u7_u4_n168 ) , .A2( u2_u7_u4_n169 ) );
  NOR2_X1 u2_u7_u4_U42 (.A1( u2_u7_u4_n150 ) , .A2( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n153 ) );
  NOR2_X1 u2_u7_u4_U43 (.A2( u2_u7_u4_n128 ) , .A1( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n156 ) );
  AOI22_X1 u2_u7_u4_U44 (.B2( u2_u7_u4_n122 ) , .A1( u2_u7_u4_n123 ) , .ZN( u2_u7_u4_n124 ) , .B1( u2_u7_u4_n128 ) , .A2( u2_u7_u4_n172 ) );
  NAND2_X1 u2_u7_u4_U45 (.A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n123 ) , .A1( u2_u7_u4_n161 ) );
  INV_X1 u2_u7_u4_U46 (.A( u2_u7_u4_n153 ) , .ZN( u2_u7_u4_n172 ) );
  AOI22_X1 u2_u7_u4_U47 (.B2( u2_u7_u4_n132 ) , .A2( u2_u7_u4_n133 ) , .ZN( u2_u7_u4_n140 ) , .A1( u2_u7_u4_n150 ) , .B1( u2_u7_u4_n179 ) );
  NAND2_X1 u2_u7_u4_U48 (.ZN( u2_u7_u4_n133 ) , .A2( u2_u7_u4_n146 ) , .A1( u2_u7_u4_n154 ) );
  NAND2_X1 u2_u7_u4_U49 (.A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n154 ) , .A2( u2_u7_u4_n98 ) );
  NOR4_X1 u2_u7_u4_U5 (.A4( u2_u7_u4_n106 ) , .A3( u2_u7_u4_n107 ) , .A2( u2_u7_u4_n108 ) , .A1( u2_u7_u4_n109 ) , .ZN( u2_u7_u4_n110 ) );
  NAND2_X1 u2_u7_u4_U50 (.A1( u2_u7_u4_n101 ) , .ZN( u2_u7_u4_n158 ) , .A2( u2_u7_u4_n99 ) );
  AOI21_X1 u2_u7_u4_U51 (.ZN( u2_u7_u4_n127 ) , .A( u2_u7_u4_n136 ) , .B2( u2_u7_u4_n150 ) , .B1( u2_u7_u4_n180 ) );
  INV_X1 u2_u7_u4_U52 (.A( u2_u7_u4_n160 ) , .ZN( u2_u7_u4_n180 ) );
  NAND2_X1 u2_u7_u4_U53 (.A2( u2_u7_u4_n104 ) , .A1( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n146 ) );
  NAND2_X1 u2_u7_u4_U54 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n160 ) );
  NAND2_X1 u2_u7_u4_U55 (.ZN( u2_u7_u4_n134 ) , .A1( u2_u7_u4_n98 ) , .A2( u2_u7_u4_n99 ) );
  NAND2_X1 u2_u7_u4_U56 (.A1( u2_u7_u4_n103 ) , .A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n143 ) );
  NAND2_X1 u2_u7_u4_U57 (.A2( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n145 ) , .A1( u2_u7_u4_n98 ) );
  NAND2_X1 u2_u7_u4_U58 (.A1( u2_u7_u4_n100 ) , .A2( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n120 ) );
  NAND2_X1 u2_u7_u4_U59 (.A1( u2_u7_u4_n102 ) , .A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n148 ) );
  AOI21_X1 u2_u7_u4_U6 (.ZN( u2_u7_u4_n106 ) , .B2( u2_u7_u4_n146 ) , .B1( u2_u7_u4_n158 ) , .A( u2_u7_u4_n170 ) );
  NAND2_X1 u2_u7_u4_U60 (.A2( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n157 ) );
  INV_X1 u2_u7_u4_U61 (.A( u2_u7_u4_n150 ) , .ZN( u2_u7_u4_n173 ) );
  INV_X1 u2_u7_u4_U62 (.A( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n171 ) );
  NAND2_X1 u2_u7_u4_U63 (.A1( u2_u7_u4_n100 ) , .ZN( u2_u7_u4_n118 ) , .A2( u2_u7_u4_n99 ) );
  NAND2_X1 u2_u7_u4_U64 (.A2( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n144 ) );
  NAND2_X1 u2_u7_u4_U65 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n96 ) );
  INV_X1 u2_u7_u4_U66 (.A( u2_u7_u4_n128 ) , .ZN( u2_u7_u4_n174 ) );
  NAND2_X1 u2_u7_u4_U67 (.A2( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n119 ) , .A1( u2_u7_u4_n98 ) );
  NAND2_X1 u2_u7_u4_U68 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n147 ) );
  NAND2_X1 u2_u7_u4_U69 (.A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n113 ) , .A1( u2_u7_u4_n99 ) );
  AOI21_X1 u2_u7_u4_U7 (.ZN( u2_u7_u4_n108 ) , .B2( u2_u7_u4_n134 ) , .B1( u2_u7_u4_n155 ) , .A( u2_u7_u4_n156 ) );
  NOR2_X1 u2_u7_u4_U70 (.A2( u2_u7_X_28 ) , .ZN( u2_u7_u4_n150 ) , .A1( u2_u7_u4_n168 ) );
  NOR2_X1 u2_u7_u4_U71 (.A2( u2_u7_X_29 ) , .ZN( u2_u7_u4_n152 ) , .A1( u2_u7_u4_n169 ) );
  NOR2_X1 u2_u7_u4_U72 (.A2( u2_u7_X_26 ) , .ZN( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n177 ) );
  NOR2_X1 u2_u7_u4_U73 (.A2( u2_u7_X_30 ) , .ZN( u2_u7_u4_n105 ) , .A1( u2_u7_u4_n176 ) );
  NOR2_X1 u2_u7_u4_U74 (.A2( u2_u7_X_28 ) , .A1( u2_u7_X_29 ) , .ZN( u2_u7_u4_n128 ) );
  NOR2_X1 u2_u7_u4_U75 (.A2( u2_u7_X_25 ) , .A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n98 ) );
  NOR2_X1 u2_u7_u4_U76 (.A2( u2_u7_X_27 ) , .A1( u2_u7_X_30 ) , .ZN( u2_u7_u4_n102 ) );
  AND2_X1 u2_u7_u4_U77 (.A2( u2_u7_X_25 ) , .A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n104 ) );
  AND2_X1 u2_u7_u4_U78 (.A1( u2_u7_X_30 ) , .A2( u2_u7_u4_n176 ) , .ZN( u2_u7_u4_n99 ) );
  AND2_X1 u2_u7_u4_U79 (.A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n101 ) , .A2( u2_u7_u4_n177 ) );
  AOI21_X1 u2_u7_u4_U8 (.ZN( u2_u7_u4_n109 ) , .A( u2_u7_u4_n153 ) , .B1( u2_u7_u4_n159 ) , .B2( u2_u7_u4_n184 ) );
  AND2_X1 u2_u7_u4_U80 (.A1( u2_u7_X_27 ) , .A2( u2_u7_X_30 ) , .ZN( u2_u7_u4_n103 ) );
  INV_X1 u2_u7_u4_U81 (.A( u2_u7_X_28 ) , .ZN( u2_u7_u4_n169 ) );
  INV_X1 u2_u7_u4_U82 (.A( u2_u7_X_29 ) , .ZN( u2_u7_u4_n168 ) );
  INV_X1 u2_u7_u4_U83 (.A( u2_u7_X_25 ) , .ZN( u2_u7_u4_n177 ) );
  INV_X1 u2_u7_u4_U84 (.A( u2_u7_X_27 ) , .ZN( u2_u7_u4_n176 ) );
  NAND4_X1 u2_u7_u4_U85 (.ZN( u2_out7_25 ) , .A4( u2_u7_u4_n139 ) , .A3( u2_u7_u4_n140 ) , .A2( u2_u7_u4_n141 ) , .A1( u2_u7_u4_n142 ) );
  OAI21_X1 u2_u7_u4_U86 (.A( u2_u7_u4_n128 ) , .B2( u2_u7_u4_n129 ) , .B1( u2_u7_u4_n130 ) , .ZN( u2_u7_u4_n142 ) );
  OAI21_X1 u2_u7_u4_U87 (.B2( u2_u7_u4_n131 ) , .ZN( u2_u7_u4_n141 ) , .A( u2_u7_u4_n175 ) , .B1( u2_u7_u4_n183 ) );
  NAND4_X1 u2_u7_u4_U88 (.ZN( u2_out7_14 ) , .A4( u2_u7_u4_n124 ) , .A3( u2_u7_u4_n125 ) , .A2( u2_u7_u4_n126 ) , .A1( u2_u7_u4_n127 ) );
  AOI22_X1 u2_u7_u4_U89 (.B2( u2_u7_u4_n117 ) , .ZN( u2_u7_u4_n126 ) , .A1( u2_u7_u4_n129 ) , .B1( u2_u7_u4_n152 ) , .A2( u2_u7_u4_n175 ) );
  AOI211_X1 u2_u7_u4_U9 (.B( u2_u7_u4_n136 ) , .A( u2_u7_u4_n137 ) , .C2( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n139 ) , .C1( u2_u7_u4_n182 ) );
  AOI22_X1 u2_u7_u4_U90 (.ZN( u2_u7_u4_n125 ) , .B2( u2_u7_u4_n131 ) , .A2( u2_u7_u4_n132 ) , .B1( u2_u7_u4_n138 ) , .A1( u2_u7_u4_n178 ) );
  NAND4_X1 u2_u7_u4_U91 (.ZN( u2_out7_8 ) , .A4( u2_u7_u4_n110 ) , .A3( u2_u7_u4_n111 ) , .A2( u2_u7_u4_n112 ) , .A1( u2_u7_u4_n186 ) );
  NAND2_X1 u2_u7_u4_U92 (.ZN( u2_u7_u4_n112 ) , .A2( u2_u7_u4_n130 ) , .A1( u2_u7_u4_n150 ) );
  AOI22_X1 u2_u7_u4_U93 (.ZN( u2_u7_u4_n111 ) , .B2( u2_u7_u4_n132 ) , .A1( u2_u7_u4_n152 ) , .B1( u2_u7_u4_n178 ) , .A2( u2_u7_u4_n97 ) );
  AOI22_X1 u2_u7_u4_U94 (.B2( u2_u7_u4_n149 ) , .B1( u2_u7_u4_n150 ) , .A2( u2_u7_u4_n151 ) , .A1( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n167 ) );
  NOR4_X1 u2_u7_u4_U95 (.A4( u2_u7_u4_n162 ) , .A3( u2_u7_u4_n163 ) , .A2( u2_u7_u4_n164 ) , .A1( u2_u7_u4_n165 ) , .ZN( u2_u7_u4_n166 ) );
  NAND3_X1 u2_u7_u4_U96 (.ZN( u2_out7_3 ) , .A3( u2_u7_u4_n166 ) , .A1( u2_u7_u4_n167 ) , .A2( u2_u7_u4_n186 ) );
  NAND3_X1 u2_u7_u4_U97 (.A3( u2_u7_u4_n146 ) , .A2( u2_u7_u4_n147 ) , .A1( u2_u7_u4_n148 ) , .ZN( u2_u7_u4_n149 ) );
  NAND3_X1 u2_u7_u4_U98 (.A3( u2_u7_u4_n143 ) , .A2( u2_u7_u4_n144 ) , .A1( u2_u7_u4_n145 ) , .ZN( u2_u7_u4_n151 ) );
  NAND3_X1 u2_u7_u4_U99 (.A3( u2_u7_u4_n121 ) , .ZN( u2_u7_u4_n122 ) , .A2( u2_u7_u4_n144 ) , .A1( u2_u7_u4_n154 ) );
  INV_X1 u2_u7_u5_U10 (.A( u2_u7_u5_n121 ) , .ZN( u2_u7_u5_n177 ) );
  NOR3_X1 u2_u7_u5_U100 (.A3( u2_u7_u5_n141 ) , .A1( u2_u7_u5_n142 ) , .ZN( u2_u7_u5_n143 ) , .A2( u2_u7_u5_n191 ) );
  NAND4_X1 u2_u7_u5_U101 (.ZN( u2_out7_4 ) , .A4( u2_u7_u5_n112 ) , .A2( u2_u7_u5_n113 ) , .A1( u2_u7_u5_n114 ) , .A3( u2_u7_u5_n195 ) );
  AOI211_X1 u2_u7_u5_U102 (.A( u2_u7_u5_n110 ) , .C1( u2_u7_u5_n111 ) , .ZN( u2_u7_u5_n112 ) , .B( u2_u7_u5_n118 ) , .C2( u2_u7_u5_n177 ) );
  AOI222_X1 u2_u7_u5_U103 (.ZN( u2_u7_u5_n113 ) , .A1( u2_u7_u5_n131 ) , .C1( u2_u7_u5_n148 ) , .B2( u2_u7_u5_n174 ) , .C2( u2_u7_u5_n178 ) , .A2( u2_u7_u5_n179 ) , .B1( u2_u7_u5_n99 ) );
  NAND3_X1 u2_u7_u5_U104 (.A2( u2_u7_u5_n154 ) , .A3( u2_u7_u5_n158 ) , .A1( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n99 ) );
  NOR2_X1 u2_u7_u5_U11 (.ZN( u2_u7_u5_n160 ) , .A2( u2_u7_u5_n173 ) , .A1( u2_u7_u5_n177 ) );
  INV_X1 u2_u7_u5_U12 (.A( u2_u7_u5_n150 ) , .ZN( u2_u7_u5_n174 ) );
  AOI21_X1 u2_u7_u5_U13 (.A( u2_u7_u5_n160 ) , .B2( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n162 ) , .B1( u2_u7_u5_n192 ) );
  INV_X1 u2_u7_u5_U14 (.A( u2_u7_u5_n159 ) , .ZN( u2_u7_u5_n192 ) );
  AOI21_X1 u2_u7_u5_U15 (.A( u2_u7_u5_n156 ) , .B2( u2_u7_u5_n157 ) , .B1( u2_u7_u5_n158 ) , .ZN( u2_u7_u5_n163 ) );
  AOI21_X1 u2_u7_u5_U16 (.B2( u2_u7_u5_n139 ) , .B1( u2_u7_u5_n140 ) , .ZN( u2_u7_u5_n141 ) , .A( u2_u7_u5_n150 ) );
  OAI21_X1 u2_u7_u5_U17 (.A( u2_u7_u5_n133 ) , .B2( u2_u7_u5_n134 ) , .B1( u2_u7_u5_n135 ) , .ZN( u2_u7_u5_n142 ) );
  OAI21_X1 u2_u7_u5_U18 (.ZN( u2_u7_u5_n133 ) , .B2( u2_u7_u5_n147 ) , .A( u2_u7_u5_n173 ) , .B1( u2_u7_u5_n188 ) );
  NAND2_X1 u2_u7_u5_U19 (.A2( u2_u7_u5_n119 ) , .A1( u2_u7_u5_n123 ) , .ZN( u2_u7_u5_n137 ) );
  INV_X1 u2_u7_u5_U20 (.A( u2_u7_u5_n155 ) , .ZN( u2_u7_u5_n194 ) );
  NAND2_X1 u2_u7_u5_U21 (.A1( u2_u7_u5_n121 ) , .ZN( u2_u7_u5_n132 ) , .A2( u2_u7_u5_n172 ) );
  NAND2_X1 u2_u7_u5_U22 (.A2( u2_u7_u5_n122 ) , .ZN( u2_u7_u5_n136 ) , .A1( u2_u7_u5_n154 ) );
  NAND2_X1 u2_u7_u5_U23 (.A2( u2_u7_u5_n119 ) , .A1( u2_u7_u5_n120 ) , .ZN( u2_u7_u5_n159 ) );
  INV_X1 u2_u7_u5_U24 (.A( u2_u7_u5_n156 ) , .ZN( u2_u7_u5_n175 ) );
  INV_X1 u2_u7_u5_U25 (.A( u2_u7_u5_n158 ) , .ZN( u2_u7_u5_n188 ) );
  INV_X1 u2_u7_u5_U26 (.A( u2_u7_u5_n152 ) , .ZN( u2_u7_u5_n179 ) );
  INV_X1 u2_u7_u5_U27 (.A( u2_u7_u5_n140 ) , .ZN( u2_u7_u5_n182 ) );
  INV_X1 u2_u7_u5_U28 (.A( u2_u7_u5_n151 ) , .ZN( u2_u7_u5_n183 ) );
  INV_X1 u2_u7_u5_U29 (.A( u2_u7_u5_n123 ) , .ZN( u2_u7_u5_n185 ) );
  NOR2_X1 u2_u7_u5_U3 (.ZN( u2_u7_u5_n134 ) , .A1( u2_u7_u5_n183 ) , .A2( u2_u7_u5_n190 ) );
  INV_X1 u2_u7_u5_U30 (.A( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n184 ) );
  INV_X1 u2_u7_u5_U31 (.A( u2_u7_u5_n139 ) , .ZN( u2_u7_u5_n189 ) );
  INV_X1 u2_u7_u5_U32 (.A( u2_u7_u5_n157 ) , .ZN( u2_u7_u5_n190 ) );
  INV_X1 u2_u7_u5_U33 (.A( u2_u7_u5_n120 ) , .ZN( u2_u7_u5_n193 ) );
  NAND2_X1 u2_u7_u5_U34 (.ZN( u2_u7_u5_n111 ) , .A1( u2_u7_u5_n140 ) , .A2( u2_u7_u5_n155 ) );
  NOR2_X1 u2_u7_u5_U35 (.ZN( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n170 ) , .A2( u2_u7_u5_n180 ) );
  INV_X1 u2_u7_u5_U36 (.A( u2_u7_u5_n117 ) , .ZN( u2_u7_u5_n196 ) );
  OAI221_X1 u2_u7_u5_U37 (.A( u2_u7_u5_n116 ) , .ZN( u2_u7_u5_n117 ) , .B2( u2_u7_u5_n119 ) , .C1( u2_u7_u5_n153 ) , .C2( u2_u7_u5_n158 ) , .B1( u2_u7_u5_n172 ) );
  AOI222_X1 u2_u7_u5_U38 (.ZN( u2_u7_u5_n116 ) , .B2( u2_u7_u5_n145 ) , .C1( u2_u7_u5_n148 ) , .A2( u2_u7_u5_n174 ) , .C2( u2_u7_u5_n177 ) , .B1( u2_u7_u5_n187 ) , .A1( u2_u7_u5_n193 ) );
  INV_X1 u2_u7_u5_U39 (.A( u2_u7_u5_n115 ) , .ZN( u2_u7_u5_n187 ) );
  INV_X1 u2_u7_u5_U4 (.A( u2_u7_u5_n138 ) , .ZN( u2_u7_u5_n191 ) );
  AOI22_X1 u2_u7_u5_U40 (.B2( u2_u7_u5_n131 ) , .A2( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n169 ) , .B1( u2_u7_u5_n174 ) , .A1( u2_u7_u5_n185 ) );
  NOR2_X1 u2_u7_u5_U41 (.A1( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n150 ) , .A2( u2_u7_u5_n173 ) );
  AOI21_X1 u2_u7_u5_U42 (.A( u2_u7_u5_n118 ) , .B2( u2_u7_u5_n145 ) , .ZN( u2_u7_u5_n168 ) , .B1( u2_u7_u5_n186 ) );
  INV_X1 u2_u7_u5_U43 (.A( u2_u7_u5_n122 ) , .ZN( u2_u7_u5_n186 ) );
  NOR2_X1 u2_u7_u5_U44 (.A1( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n152 ) , .A2( u2_u7_u5_n176 ) );
  NOR2_X1 u2_u7_u5_U45 (.A1( u2_u7_u5_n115 ) , .ZN( u2_u7_u5_n118 ) , .A2( u2_u7_u5_n153 ) );
  NOR2_X1 u2_u7_u5_U46 (.A2( u2_u7_u5_n145 ) , .ZN( u2_u7_u5_n156 ) , .A1( u2_u7_u5_n174 ) );
  NOR2_X1 u2_u7_u5_U47 (.ZN( u2_u7_u5_n121 ) , .A2( u2_u7_u5_n145 ) , .A1( u2_u7_u5_n176 ) );
  AOI22_X1 u2_u7_u5_U48 (.ZN( u2_u7_u5_n114 ) , .A2( u2_u7_u5_n137 ) , .A1( u2_u7_u5_n145 ) , .B2( u2_u7_u5_n175 ) , .B1( u2_u7_u5_n193 ) );
  OAI211_X1 u2_u7_u5_U49 (.B( u2_u7_u5_n124 ) , .A( u2_u7_u5_n125 ) , .C2( u2_u7_u5_n126 ) , .C1( u2_u7_u5_n127 ) , .ZN( u2_u7_u5_n128 ) );
  OAI21_X1 u2_u7_u5_U5 (.B2( u2_u7_u5_n136 ) , .B1( u2_u7_u5_n137 ) , .ZN( u2_u7_u5_n138 ) , .A( u2_u7_u5_n177 ) );
  NOR3_X1 u2_u7_u5_U50 (.ZN( u2_u7_u5_n127 ) , .A1( u2_u7_u5_n136 ) , .A3( u2_u7_u5_n148 ) , .A2( u2_u7_u5_n182 ) );
  OAI21_X1 u2_u7_u5_U51 (.ZN( u2_u7_u5_n124 ) , .A( u2_u7_u5_n177 ) , .B2( u2_u7_u5_n183 ) , .B1( u2_u7_u5_n189 ) );
  OAI21_X1 u2_u7_u5_U52 (.ZN( u2_u7_u5_n125 ) , .A( u2_u7_u5_n174 ) , .B2( u2_u7_u5_n185 ) , .B1( u2_u7_u5_n190 ) );
  AOI21_X1 u2_u7_u5_U53 (.A( u2_u7_u5_n153 ) , .B2( u2_u7_u5_n154 ) , .B1( u2_u7_u5_n155 ) , .ZN( u2_u7_u5_n164 ) );
  AOI21_X1 u2_u7_u5_U54 (.ZN( u2_u7_u5_n110 ) , .B1( u2_u7_u5_n122 ) , .B2( u2_u7_u5_n139 ) , .A( u2_u7_u5_n153 ) );
  INV_X1 u2_u7_u5_U55 (.A( u2_u7_u5_n153 ) , .ZN( u2_u7_u5_n176 ) );
  INV_X1 u2_u7_u5_U56 (.A( u2_u7_u5_n126 ) , .ZN( u2_u7_u5_n173 ) );
  AND2_X1 u2_u7_u5_U57 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n147 ) );
  AND2_X1 u2_u7_u5_U58 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n148 ) );
  NAND2_X1 u2_u7_u5_U59 (.A1( u2_u7_u5_n105 ) , .A2( u2_u7_u5_n106 ) , .ZN( u2_u7_u5_n158 ) );
  INV_X1 u2_u7_u5_U6 (.A( u2_u7_u5_n135 ) , .ZN( u2_u7_u5_n178 ) );
  NAND2_X1 u2_u7_u5_U60 (.A2( u2_u7_u5_n108 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n139 ) );
  NAND2_X1 u2_u7_u5_U61 (.A1( u2_u7_u5_n106 ) , .A2( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n119 ) );
  NAND2_X1 u2_u7_u5_U62 (.A2( u2_u7_u5_n103 ) , .A1( u2_u7_u5_n105 ) , .ZN( u2_u7_u5_n140 ) );
  NAND2_X1 u2_u7_u5_U63 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n105 ) , .ZN( u2_u7_u5_n155 ) );
  NAND2_X1 u2_u7_u5_U64 (.A2( u2_u7_u5_n106 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n122 ) );
  NAND2_X1 u2_u7_u5_U65 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n106 ) , .ZN( u2_u7_u5_n115 ) );
  NAND2_X1 u2_u7_u5_U66 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n103 ) , .ZN( u2_u7_u5_n161 ) );
  NAND2_X1 u2_u7_u5_U67 (.A1( u2_u7_u5_n105 ) , .A2( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n154 ) );
  INV_X1 u2_u7_u5_U68 (.A( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n172 ) );
  NAND2_X1 u2_u7_u5_U69 (.A1( u2_u7_u5_n103 ) , .A2( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n123 ) );
  OAI22_X1 u2_u7_u5_U7 (.B2( u2_u7_u5_n149 ) , .B1( u2_u7_u5_n150 ) , .A2( u2_u7_u5_n151 ) , .A1( u2_u7_u5_n152 ) , .ZN( u2_u7_u5_n165 ) );
  NAND2_X1 u2_u7_u5_U70 (.A2( u2_u7_u5_n103 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n151 ) );
  NAND2_X1 u2_u7_u5_U71 (.A2( u2_u7_u5_n107 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n120 ) );
  NAND2_X1 u2_u7_u5_U72 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n157 ) );
  AND2_X1 u2_u7_u5_U73 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n104 ) , .ZN( u2_u7_u5_n131 ) );
  INV_X1 u2_u7_u5_U74 (.A( u2_u7_u5_n102 ) , .ZN( u2_u7_u5_n195 ) );
  OAI221_X1 u2_u7_u5_U75 (.A( u2_u7_u5_n101 ) , .ZN( u2_u7_u5_n102 ) , .C2( u2_u7_u5_n115 ) , .C1( u2_u7_u5_n126 ) , .B1( u2_u7_u5_n134 ) , .B2( u2_u7_u5_n160 ) );
  OAI21_X1 u2_u7_u5_U76 (.ZN( u2_u7_u5_n101 ) , .B1( u2_u7_u5_n137 ) , .A( u2_u7_u5_n146 ) , .B2( u2_u7_u5_n147 ) );
  NOR2_X1 u2_u7_u5_U77 (.A2( u2_u7_X_34 ) , .A1( u2_u7_X_35 ) , .ZN( u2_u7_u5_n145 ) );
  NOR2_X1 u2_u7_u5_U78 (.A2( u2_u7_X_34 ) , .ZN( u2_u7_u5_n146 ) , .A1( u2_u7_u5_n171 ) );
  NOR2_X1 u2_u7_u5_U79 (.A2( u2_u7_X_31 ) , .A1( u2_u7_X_32 ) , .ZN( u2_u7_u5_n103 ) );
  NOR3_X1 u2_u7_u5_U8 (.A2( u2_u7_u5_n147 ) , .A1( u2_u7_u5_n148 ) , .ZN( u2_u7_u5_n149 ) , .A3( u2_u7_u5_n194 ) );
  NOR2_X1 u2_u7_u5_U80 (.A2( u2_u7_X_36 ) , .ZN( u2_u7_u5_n105 ) , .A1( u2_u7_u5_n180 ) );
  NOR2_X1 u2_u7_u5_U81 (.A2( u2_u7_X_33 ) , .ZN( u2_u7_u5_n108 ) , .A1( u2_u7_u5_n170 ) );
  NOR2_X1 u2_u7_u5_U82 (.A2( u2_u7_X_33 ) , .A1( u2_u7_X_36 ) , .ZN( u2_u7_u5_n107 ) );
  NOR2_X1 u2_u7_u5_U83 (.A2( u2_u7_X_31 ) , .ZN( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n181 ) );
  NAND2_X1 u2_u7_u5_U84 (.A2( u2_u7_X_34 ) , .A1( u2_u7_X_35 ) , .ZN( u2_u7_u5_n153 ) );
  NAND2_X1 u2_u7_u5_U85 (.A1( u2_u7_X_34 ) , .ZN( u2_u7_u5_n126 ) , .A2( u2_u7_u5_n171 ) );
  AND2_X1 u2_u7_u5_U86 (.A1( u2_u7_X_31 ) , .A2( u2_u7_X_32 ) , .ZN( u2_u7_u5_n106 ) );
  AND2_X1 u2_u7_u5_U87 (.A1( u2_u7_X_31 ) , .ZN( u2_u7_u5_n109 ) , .A2( u2_u7_u5_n181 ) );
  INV_X1 u2_u7_u5_U88 (.A( u2_u7_X_33 ) , .ZN( u2_u7_u5_n180 ) );
  INV_X1 u2_u7_u5_U89 (.A( u2_u7_X_35 ) , .ZN( u2_u7_u5_n171 ) );
  NOR2_X1 u2_u7_u5_U9 (.ZN( u2_u7_u5_n135 ) , .A1( u2_u7_u5_n173 ) , .A2( u2_u7_u5_n176 ) );
  INV_X1 u2_u7_u5_U90 (.A( u2_u7_X_36 ) , .ZN( u2_u7_u5_n170 ) );
  INV_X1 u2_u7_u5_U91 (.A( u2_u7_X_32 ) , .ZN( u2_u7_u5_n181 ) );
  NAND4_X1 u2_u7_u5_U92 (.ZN( u2_out7_29 ) , .A4( u2_u7_u5_n129 ) , .A3( u2_u7_u5_n130 ) , .A2( u2_u7_u5_n168 ) , .A1( u2_u7_u5_n196 ) );
  AOI221_X1 u2_u7_u5_U93 (.A( u2_u7_u5_n128 ) , .ZN( u2_u7_u5_n129 ) , .C2( u2_u7_u5_n132 ) , .B2( u2_u7_u5_n159 ) , .B1( u2_u7_u5_n176 ) , .C1( u2_u7_u5_n184 ) );
  AOI222_X1 u2_u7_u5_U94 (.ZN( u2_u7_u5_n130 ) , .A2( u2_u7_u5_n146 ) , .B1( u2_u7_u5_n147 ) , .C2( u2_u7_u5_n175 ) , .B2( u2_u7_u5_n179 ) , .A1( u2_u7_u5_n188 ) , .C1( u2_u7_u5_n194 ) );
  NAND4_X1 u2_u7_u5_U95 (.ZN( u2_out7_19 ) , .A4( u2_u7_u5_n166 ) , .A3( u2_u7_u5_n167 ) , .A2( u2_u7_u5_n168 ) , .A1( u2_u7_u5_n169 ) );
  AOI22_X1 u2_u7_u5_U96 (.B2( u2_u7_u5_n145 ) , .A2( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n167 ) , .B1( u2_u7_u5_n182 ) , .A1( u2_u7_u5_n189 ) );
  NOR4_X1 u2_u7_u5_U97 (.A4( u2_u7_u5_n162 ) , .A3( u2_u7_u5_n163 ) , .A2( u2_u7_u5_n164 ) , .A1( u2_u7_u5_n165 ) , .ZN( u2_u7_u5_n166 ) );
  NAND4_X1 u2_u7_u5_U98 (.ZN( u2_out7_11 ) , .A4( u2_u7_u5_n143 ) , .A3( u2_u7_u5_n144 ) , .A2( u2_u7_u5_n169 ) , .A1( u2_u7_u5_n196 ) );
  AOI22_X1 u2_u7_u5_U99 (.A2( u2_u7_u5_n132 ) , .ZN( u2_u7_u5_n144 ) , .B2( u2_u7_u5_n145 ) , .B1( u2_u7_u5_n184 ) , .A1( u2_u7_u5_n194 ) );
  XOR2_X1 u2_u8_U1 (.B( u2_K9_9 ) , .A( u2_R7_6 ) , .Z( u2_u8_X_9 ) );
  XOR2_X1 u2_u8_U10 (.B( u2_K9_45 ) , .A( u2_R7_30 ) , .Z( u2_u8_X_45 ) );
  XOR2_X1 u2_u8_U11 (.B( u2_K9_44 ) , .A( u2_R7_29 ) , .Z( u2_u8_X_44 ) );
  XOR2_X1 u2_u8_U12 (.B( u2_K9_43 ) , .A( u2_R7_28 ) , .Z( u2_u8_X_43 ) );
  XOR2_X1 u2_u8_U13 (.B( u2_K9_42 ) , .A( u2_R7_29 ) , .Z( u2_u8_X_42 ) );
  XOR2_X1 u2_u8_U14 (.B( u2_K9_41 ) , .A( u2_R7_28 ) , .Z( u2_u8_X_41 ) );
  XOR2_X1 u2_u8_U15 (.B( u2_K9_40 ) , .A( u2_R7_27 ) , .Z( u2_u8_X_40 ) );
  XOR2_X1 u2_u8_U16 (.B( u2_K9_3 ) , .A( u2_R7_2 ) , .Z( u2_u8_X_3 ) );
  XOR2_X1 u2_u8_U17 (.B( u2_K9_39 ) , .A( u2_R7_26 ) , .Z( u2_u8_X_39 ) );
  XOR2_X1 u2_u8_U18 (.B( u2_K9_38 ) , .A( u2_R7_25 ) , .Z( u2_u8_X_38 ) );
  XOR2_X1 u2_u8_U19 (.B( u2_K9_37 ) , .A( u2_R7_24 ) , .Z( u2_u8_X_37 ) );
  XOR2_X1 u2_u8_U2 (.B( u2_K9_8 ) , .A( u2_R7_5 ) , .Z( u2_u8_X_8 ) );
  XOR2_X1 u2_u8_U26 (.B( u2_K9_30 ) , .A( u2_R7_21 ) , .Z( u2_u8_X_30 ) );
  XOR2_X1 u2_u8_U27 (.B( u2_K9_2 ) , .A( u2_R7_1 ) , .Z( u2_u8_X_2 ) );
  XOR2_X1 u2_u8_U28 (.B( u2_K9_29 ) , .A( u2_R7_20 ) , .Z( u2_u8_X_29 ) );
  XOR2_X1 u2_u8_U29 (.B( u2_K9_28 ) , .A( u2_R7_19 ) , .Z( u2_u8_X_28 ) );
  XOR2_X1 u2_u8_U3 (.B( u2_K9_7 ) , .A( u2_R7_4 ) , .Z( u2_u8_X_7 ) );
  XOR2_X1 u2_u8_U30 (.B( u2_K9_27 ) , .A( u2_R7_18 ) , .Z( u2_u8_X_27 ) );
  XOR2_X1 u2_u8_U31 (.B( u2_K9_26 ) , .A( u2_R7_17 ) , .Z( u2_u8_X_26 ) );
  XOR2_X1 u2_u8_U32 (.B( u2_K9_25 ) , .A( u2_R7_16 ) , .Z( u2_u8_X_25 ) );
  XOR2_X1 u2_u8_U33 (.B( u2_K9_24 ) , .A( u2_R7_17 ) , .Z( u2_u8_X_24 ) );
  XOR2_X1 u2_u8_U34 (.B( u2_K9_23 ) , .A( u2_R7_16 ) , .Z( u2_u8_X_23 ) );
  XOR2_X1 u2_u8_U35 (.B( u2_K9_22 ) , .A( u2_R7_15 ) , .Z( u2_u8_X_22 ) );
  XOR2_X1 u2_u8_U36 (.B( u2_K9_21 ) , .A( u2_R7_14 ) , .Z( u2_u8_X_21 ) );
  XOR2_X1 u2_u8_U37 (.B( u2_K9_20 ) , .A( u2_R7_13 ) , .Z( u2_u8_X_20 ) );
  XOR2_X1 u2_u8_U38 (.B( u2_K9_1 ) , .A( u2_R7_32 ) , .Z( u2_u8_X_1 ) );
  XOR2_X1 u2_u8_U39 (.B( u2_K9_19 ) , .A( u2_R7_12 ) , .Z( u2_u8_X_19 ) );
  XOR2_X1 u2_u8_U4 (.B( u2_K9_6 ) , .A( u2_R7_5 ) , .Z( u2_u8_X_6 ) );
  XOR2_X1 u2_u8_U40 (.B( u2_K9_18 ) , .A( u2_R7_13 ) , .Z( u2_u8_X_18 ) );
  XOR2_X1 u2_u8_U41 (.B( u2_K9_17 ) , .A( u2_R7_12 ) , .Z( u2_u8_X_17 ) );
  XOR2_X1 u2_u8_U42 (.B( u2_K9_16 ) , .A( u2_R7_11 ) , .Z( u2_u8_X_16 ) );
  XOR2_X1 u2_u8_U43 (.B( u2_K9_15 ) , .A( u2_R7_10 ) , .Z( u2_u8_X_15 ) );
  XOR2_X1 u2_u8_U44 (.B( u2_K9_14 ) , .A( u2_R7_9 ) , .Z( u2_u8_X_14 ) );
  XOR2_X1 u2_u8_U45 (.B( u2_K9_13 ) , .A( u2_R7_8 ) , .Z( u2_u8_X_13 ) );
  XOR2_X1 u2_u8_U46 (.B( u2_K9_12 ) , .A( u2_R7_9 ) , .Z( u2_u8_X_12 ) );
  XOR2_X1 u2_u8_U47 (.B( u2_K9_11 ) , .A( u2_R7_8 ) , .Z( u2_u8_X_11 ) );
  XOR2_X1 u2_u8_U48 (.B( u2_K9_10 ) , .A( u2_R7_7 ) , .Z( u2_u8_X_10 ) );
  XOR2_X1 u2_u8_U5 (.B( u2_K9_5 ) , .A( u2_R7_4 ) , .Z( u2_u8_X_5 ) );
  XOR2_X1 u2_u8_U6 (.B( u2_K9_4 ) , .A( u2_R7_3 ) , .Z( u2_u8_X_4 ) );
  XOR2_X1 u2_u8_U7 (.B( u2_K9_48 ) , .A( u2_R7_1 ) , .Z( u2_u8_X_48 ) );
  XOR2_X1 u2_u8_U8 (.B( u2_K9_47 ) , .A( u2_R7_32 ) , .Z( u2_u8_X_47 ) );
  XOR2_X1 u2_u8_U9 (.B( u2_K9_46 ) , .A( u2_R7_31 ) , .Z( u2_u8_X_46 ) );
  AND2_X1 u2_u8_u0_U10 (.A1( u2_u8_u0_n131 ) , .ZN( u2_u8_u0_n141 ) , .A2( u2_u8_u0_n150 ) );
  AND3_X1 u2_u8_u0_U11 (.A2( u2_u8_u0_n112 ) , .ZN( u2_u8_u0_n127 ) , .A3( u2_u8_u0_n130 ) , .A1( u2_u8_u0_n148 ) );
  AND2_X1 u2_u8_u0_U12 (.ZN( u2_u8_u0_n107 ) , .A1( u2_u8_u0_n130 ) , .A2( u2_u8_u0_n140 ) );
  AND2_X1 u2_u8_u0_U13 (.A2( u2_u8_u0_n129 ) , .A1( u2_u8_u0_n130 ) , .ZN( u2_u8_u0_n151 ) );
  AND2_X1 u2_u8_u0_U14 (.A1( u2_u8_u0_n108 ) , .A2( u2_u8_u0_n125 ) , .ZN( u2_u8_u0_n145 ) );
  INV_X1 u2_u8_u0_U15 (.A( u2_u8_u0_n143 ) , .ZN( u2_u8_u0_n173 ) );
  NOR2_X1 u2_u8_u0_U16 (.A2( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n147 ) , .A1( u2_u8_u0_n160 ) );
  AOI21_X1 u2_u8_u0_U17 (.B1( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n132 ) , .A( u2_u8_u0_n165 ) , .B2( u2_u8_u0_n93 ) );
  OAI22_X1 u2_u8_u0_U18 (.B1( u2_u8_u0_n131 ) , .A1( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n147 ) , .A2( u2_u8_u0_n90 ) , .ZN( u2_u8_u0_n91 ) );
  AND3_X1 u2_u8_u0_U19 (.A3( u2_u8_u0_n121 ) , .A2( u2_u8_u0_n125 ) , .A1( u2_u8_u0_n148 ) , .ZN( u2_u8_u0_n90 ) );
  OAI22_X1 u2_u8_u0_U20 (.B1( u2_u8_u0_n125 ) , .ZN( u2_u8_u0_n126 ) , .A1( u2_u8_u0_n138 ) , .A2( u2_u8_u0_n146 ) , .B2( u2_u8_u0_n147 ) );
  NOR2_X1 u2_u8_u0_U21 (.A1( u2_u8_u0_n163 ) , .A2( u2_u8_u0_n164 ) , .ZN( u2_u8_u0_n95 ) );
  AOI22_X1 u2_u8_u0_U22 (.B2( u2_u8_u0_n109 ) , .A2( u2_u8_u0_n110 ) , .ZN( u2_u8_u0_n111 ) , .B1( u2_u8_u0_n118 ) , .A1( u2_u8_u0_n160 ) );
  NAND2_X1 u2_u8_u0_U23 (.A2( u2_u8_u0_n102 ) , .A1( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n149 ) );
  INV_X1 u2_u8_u0_U24 (.A( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n161 ) );
  INV_X1 u2_u8_u0_U25 (.A( u2_u8_u0_n118 ) , .ZN( u2_u8_u0_n158 ) );
  NAND2_X1 u2_u8_u0_U26 (.A2( u2_u8_u0_n100 ) , .ZN( u2_u8_u0_n131 ) , .A1( u2_u8_u0_n92 ) );
  NAND2_X1 u2_u8_u0_U27 (.ZN( u2_u8_u0_n108 ) , .A1( u2_u8_u0_n92 ) , .A2( u2_u8_u0_n94 ) );
  AOI21_X1 u2_u8_u0_U28 (.ZN( u2_u8_u0_n104 ) , .B1( u2_u8_u0_n107 ) , .B2( u2_u8_u0_n141 ) , .A( u2_u8_u0_n144 ) );
  AOI21_X1 u2_u8_u0_U29 (.B1( u2_u8_u0_n127 ) , .B2( u2_u8_u0_n129 ) , .A( u2_u8_u0_n138 ) , .ZN( u2_u8_u0_n96 ) );
  INV_X1 u2_u8_u0_U3 (.A( u2_u8_u0_n113 ) , .ZN( u2_u8_u0_n166 ) );
  NAND2_X1 u2_u8_u0_U30 (.A2( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n114 ) , .A1( u2_u8_u0_n92 ) );
  NOR2_X1 u2_u8_u0_U31 (.A1( u2_u8_u0_n120 ) , .ZN( u2_u8_u0_n143 ) , .A2( u2_u8_u0_n167 ) );
  OAI221_X1 u2_u8_u0_U32 (.C1( u2_u8_u0_n112 ) , .ZN( u2_u8_u0_n120 ) , .B1( u2_u8_u0_n138 ) , .B2( u2_u8_u0_n141 ) , .C2( u2_u8_u0_n147 ) , .A( u2_u8_u0_n172 ) );
  AOI211_X1 u2_u8_u0_U33 (.B( u2_u8_u0_n115 ) , .A( u2_u8_u0_n116 ) , .C2( u2_u8_u0_n117 ) , .C1( u2_u8_u0_n118 ) , .ZN( u2_u8_u0_n119 ) );
  NAND2_X1 u2_u8_u0_U34 (.A2( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n140 ) , .A1( u2_u8_u0_n94 ) );
  NAND2_X1 u2_u8_u0_U35 (.A1( u2_u8_u0_n100 ) , .A2( u2_u8_u0_n103 ) , .ZN( u2_u8_u0_n125 ) );
  NAND2_X1 u2_u8_u0_U36 (.A1( u2_u8_u0_n101 ) , .A2( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n150 ) );
  INV_X1 u2_u8_u0_U37 (.A( u2_u8_u0_n138 ) , .ZN( u2_u8_u0_n160 ) );
  NAND2_X1 u2_u8_u0_U38 (.A2( u2_u8_u0_n100 ) , .A1( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n139 ) );
  NAND2_X1 u2_u8_u0_U39 (.ZN( u2_u8_u0_n112 ) , .A2( u2_u8_u0_n92 ) , .A1( u2_u8_u0_n93 ) );
  AOI21_X1 u2_u8_u0_U4 (.B1( u2_u8_u0_n114 ) , .ZN( u2_u8_u0_n115 ) , .B2( u2_u8_u0_n129 ) , .A( u2_u8_u0_n161 ) );
  NAND2_X1 u2_u8_u0_U40 (.A1( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n130 ) , .A2( u2_u8_u0_n94 ) );
  INV_X1 u2_u8_u0_U41 (.ZN( u2_u8_u0_n172 ) , .A( u2_u8_u0_n88 ) );
  OAI222_X1 u2_u8_u0_U42 (.C1( u2_u8_u0_n108 ) , .A1( u2_u8_u0_n125 ) , .B2( u2_u8_u0_n128 ) , .B1( u2_u8_u0_n144 ) , .A2( u2_u8_u0_n158 ) , .C2( u2_u8_u0_n161 ) , .ZN( u2_u8_u0_n88 ) );
  NAND2_X1 u2_u8_u0_U43 (.A2( u2_u8_u0_n101 ) , .ZN( u2_u8_u0_n121 ) , .A1( u2_u8_u0_n93 ) );
  OR3_X1 u2_u8_u0_U44 (.A3( u2_u8_u0_n152 ) , .A2( u2_u8_u0_n153 ) , .A1( u2_u8_u0_n154 ) , .ZN( u2_u8_u0_n155 ) );
  AOI21_X1 u2_u8_u0_U45 (.A( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n145 ) , .B1( u2_u8_u0_n146 ) , .ZN( u2_u8_u0_n154 ) );
  AOI21_X1 u2_u8_u0_U46 (.B2( u2_u8_u0_n150 ) , .B1( u2_u8_u0_n151 ) , .ZN( u2_u8_u0_n152 ) , .A( u2_u8_u0_n158 ) );
  AOI21_X1 u2_u8_u0_U47 (.A( u2_u8_u0_n147 ) , .B2( u2_u8_u0_n148 ) , .B1( u2_u8_u0_n149 ) , .ZN( u2_u8_u0_n153 ) );
  INV_X1 u2_u8_u0_U48 (.ZN( u2_u8_u0_n171 ) , .A( u2_u8_u0_n99 ) );
  OAI211_X1 u2_u8_u0_U49 (.C2( u2_u8_u0_n140 ) , .C1( u2_u8_u0_n161 ) , .A( u2_u8_u0_n169 ) , .B( u2_u8_u0_n98 ) , .ZN( u2_u8_u0_n99 ) );
  AOI21_X1 u2_u8_u0_U5 (.B2( u2_u8_u0_n131 ) , .ZN( u2_u8_u0_n134 ) , .B1( u2_u8_u0_n151 ) , .A( u2_u8_u0_n158 ) );
  INV_X1 u2_u8_u0_U50 (.ZN( u2_u8_u0_n169 ) , .A( u2_u8_u0_n91 ) );
  AOI211_X1 u2_u8_u0_U51 (.C1( u2_u8_u0_n118 ) , .A( u2_u8_u0_n123 ) , .B( u2_u8_u0_n96 ) , .C2( u2_u8_u0_n97 ) , .ZN( u2_u8_u0_n98 ) );
  NOR2_X1 u2_u8_u0_U52 (.A2( u2_u8_X_4 ) , .A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n118 ) );
  NOR2_X1 u2_u8_u0_U53 (.A2( u2_u8_X_1 ) , .ZN( u2_u8_u0_n101 ) , .A1( u2_u8_u0_n163 ) );
  NOR2_X1 u2_u8_u0_U54 (.A2( u2_u8_X_3 ) , .A1( u2_u8_X_6 ) , .ZN( u2_u8_u0_n94 ) );
  NOR2_X1 u2_u8_u0_U55 (.A2( u2_u8_X_6 ) , .ZN( u2_u8_u0_n100 ) , .A1( u2_u8_u0_n162 ) );
  NAND2_X1 u2_u8_u0_U56 (.A2( u2_u8_X_4 ) , .A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n144 ) );
  NOR2_X1 u2_u8_u0_U57 (.A2( u2_u8_X_5 ) , .ZN( u2_u8_u0_n136 ) , .A1( u2_u8_u0_n159 ) );
  NAND2_X1 u2_u8_u0_U58 (.A1( u2_u8_X_5 ) , .ZN( u2_u8_u0_n138 ) , .A2( u2_u8_u0_n159 ) );
  AND2_X1 u2_u8_u0_U59 (.A2( u2_u8_X_3 ) , .A1( u2_u8_X_6 ) , .ZN( u2_u8_u0_n102 ) );
  NOR2_X1 u2_u8_u0_U6 (.A1( u2_u8_u0_n108 ) , .ZN( u2_u8_u0_n123 ) , .A2( u2_u8_u0_n158 ) );
  AND2_X1 u2_u8_u0_U60 (.A1( u2_u8_X_6 ) , .A2( u2_u8_u0_n162 ) , .ZN( u2_u8_u0_n93 ) );
  INV_X1 u2_u8_u0_U61 (.A( u2_u8_X_4 ) , .ZN( u2_u8_u0_n159 ) );
  INV_X1 u2_u8_u0_U62 (.A( u2_u8_X_1 ) , .ZN( u2_u8_u0_n164 ) );
  INV_X1 u2_u8_u0_U63 (.A( u2_u8_X_3 ) , .ZN( u2_u8_u0_n162 ) );
  INV_X1 u2_u8_u0_U64 (.A( u2_u8_u0_n126 ) , .ZN( u2_u8_u0_n168 ) );
  AOI211_X1 u2_u8_u0_U65 (.B( u2_u8_u0_n133 ) , .A( u2_u8_u0_n134 ) , .C2( u2_u8_u0_n135 ) , .C1( u2_u8_u0_n136 ) , .ZN( u2_u8_u0_n137 ) );
  OR4_X1 u2_u8_u0_U66 (.ZN( u2_out8_17 ) , .A4( u2_u8_u0_n122 ) , .A2( u2_u8_u0_n123 ) , .A1( u2_u8_u0_n124 ) , .A3( u2_u8_u0_n170 ) );
  AOI21_X1 u2_u8_u0_U67 (.B2( u2_u8_u0_n107 ) , .ZN( u2_u8_u0_n124 ) , .B1( u2_u8_u0_n128 ) , .A( u2_u8_u0_n161 ) );
  INV_X1 u2_u8_u0_U68 (.A( u2_u8_u0_n111 ) , .ZN( u2_u8_u0_n170 ) );
  OR4_X1 u2_u8_u0_U69 (.ZN( u2_out8_31 ) , .A4( u2_u8_u0_n155 ) , .A2( u2_u8_u0_n156 ) , .A1( u2_u8_u0_n157 ) , .A3( u2_u8_u0_n173 ) );
  OAI21_X1 u2_u8_u0_U7 (.B1( u2_u8_u0_n150 ) , .B2( u2_u8_u0_n158 ) , .A( u2_u8_u0_n172 ) , .ZN( u2_u8_u0_n89 ) );
  AOI21_X1 u2_u8_u0_U70 (.A( u2_u8_u0_n138 ) , .B2( u2_u8_u0_n139 ) , .B1( u2_u8_u0_n140 ) , .ZN( u2_u8_u0_n157 ) );
  AOI211_X1 u2_u8_u0_U71 (.B( u2_u8_u0_n104 ) , .A( u2_u8_u0_n105 ) , .ZN( u2_u8_u0_n106 ) , .C2( u2_u8_u0_n113 ) , .C1( u2_u8_u0_n160 ) );
  INV_X1 u2_u8_u0_U72 (.ZN( u2_u8_u0_n174 ) , .A( u2_u8_u0_n89 ) );
  INV_X1 u2_u8_u0_U73 (.A( u2_u8_u0_n142 ) , .ZN( u2_u8_u0_n165 ) );
  AOI21_X1 u2_u8_u0_U74 (.ZN( u2_u8_u0_n116 ) , .B2( u2_u8_u0_n142 ) , .A( u2_u8_u0_n144 ) , .B1( u2_u8_u0_n166 ) );
  AOI21_X1 u2_u8_u0_U75 (.B2( u2_u8_u0_n141 ) , .B1( u2_u8_u0_n142 ) , .ZN( u2_u8_u0_n156 ) , .A( u2_u8_u0_n161 ) );
  OAI221_X1 u2_u8_u0_U76 (.C1( u2_u8_u0_n121 ) , .ZN( u2_u8_u0_n122 ) , .B2( u2_u8_u0_n127 ) , .A( u2_u8_u0_n143 ) , .B1( u2_u8_u0_n144 ) , .C2( u2_u8_u0_n147 ) );
  AOI21_X1 u2_u8_u0_U77 (.B1( u2_u8_u0_n132 ) , .ZN( u2_u8_u0_n133 ) , .A( u2_u8_u0_n144 ) , .B2( u2_u8_u0_n166 ) );
  OAI22_X1 u2_u8_u0_U78 (.ZN( u2_u8_u0_n105 ) , .A2( u2_u8_u0_n132 ) , .B1( u2_u8_u0_n146 ) , .A1( u2_u8_u0_n147 ) , .B2( u2_u8_u0_n161 ) );
  NAND2_X1 u2_u8_u0_U79 (.ZN( u2_u8_u0_n110 ) , .A2( u2_u8_u0_n132 ) , .A1( u2_u8_u0_n145 ) );
  AND2_X1 u2_u8_u0_U8 (.A1( u2_u8_u0_n114 ) , .A2( u2_u8_u0_n121 ) , .ZN( u2_u8_u0_n146 ) );
  INV_X1 u2_u8_u0_U80 (.A( u2_u8_u0_n119 ) , .ZN( u2_u8_u0_n167 ) );
  NAND2_X1 u2_u8_u0_U81 (.ZN( u2_u8_u0_n148 ) , .A1( u2_u8_u0_n93 ) , .A2( u2_u8_u0_n95 ) );
  NAND2_X1 u2_u8_u0_U82 (.A1( u2_u8_u0_n100 ) , .ZN( u2_u8_u0_n129 ) , .A2( u2_u8_u0_n95 ) );
  NAND2_X1 u2_u8_u0_U83 (.A1( u2_u8_u0_n102 ) , .ZN( u2_u8_u0_n128 ) , .A2( u2_u8_u0_n95 ) );
  NOR2_X1 u2_u8_u0_U84 (.A2( u2_u8_X_1 ) , .A1( u2_u8_X_2 ) , .ZN( u2_u8_u0_n92 ) );
  NAND2_X1 u2_u8_u0_U85 (.ZN( u2_u8_u0_n142 ) , .A1( u2_u8_u0_n94 ) , .A2( u2_u8_u0_n95 ) );
  NOR2_X1 u2_u8_u0_U86 (.A2( u2_u8_X_2 ) , .ZN( u2_u8_u0_n103 ) , .A1( u2_u8_u0_n164 ) );
  INV_X1 u2_u8_u0_U87 (.A( u2_u8_X_2 ) , .ZN( u2_u8_u0_n163 ) );
  NAND3_X1 u2_u8_u0_U88 (.ZN( u2_out8_23 ) , .A3( u2_u8_u0_n137 ) , .A1( u2_u8_u0_n168 ) , .A2( u2_u8_u0_n171 ) );
  NAND3_X1 u2_u8_u0_U89 (.A3( u2_u8_u0_n127 ) , .A2( u2_u8_u0_n128 ) , .ZN( u2_u8_u0_n135 ) , .A1( u2_u8_u0_n150 ) );
  NAND2_X1 u2_u8_u0_U9 (.ZN( u2_u8_u0_n113 ) , .A1( u2_u8_u0_n139 ) , .A2( u2_u8_u0_n149 ) );
  NAND3_X1 u2_u8_u0_U90 (.ZN( u2_u8_u0_n117 ) , .A3( u2_u8_u0_n132 ) , .A2( u2_u8_u0_n139 ) , .A1( u2_u8_u0_n148 ) );
  NAND3_X1 u2_u8_u0_U91 (.ZN( u2_u8_u0_n109 ) , .A2( u2_u8_u0_n114 ) , .A3( u2_u8_u0_n140 ) , .A1( u2_u8_u0_n149 ) );
  NAND3_X1 u2_u8_u0_U92 (.ZN( u2_out8_9 ) , .A3( u2_u8_u0_n106 ) , .A2( u2_u8_u0_n171 ) , .A1( u2_u8_u0_n174 ) );
  NAND3_X1 u2_u8_u0_U93 (.A2( u2_u8_u0_n128 ) , .A1( u2_u8_u0_n132 ) , .A3( u2_u8_u0_n146 ) , .ZN( u2_u8_u0_n97 ) );
  AOI21_X1 u2_u8_u1_U10 (.B2( u2_u8_u1_n155 ) , .B1( u2_u8_u1_n156 ) , .ZN( u2_u8_u1_n157 ) , .A( u2_u8_u1_n174 ) );
  NAND3_X1 u2_u8_u1_U100 (.ZN( u2_u8_u1_n113 ) , .A1( u2_u8_u1_n120 ) , .A3( u2_u8_u1_n133 ) , .A2( u2_u8_u1_n155 ) );
  NAND2_X1 u2_u8_u1_U11 (.ZN( u2_u8_u1_n140 ) , .A2( u2_u8_u1_n150 ) , .A1( u2_u8_u1_n155 ) );
  NAND2_X1 u2_u8_u1_U12 (.A1( u2_u8_u1_n131 ) , .ZN( u2_u8_u1_n147 ) , .A2( u2_u8_u1_n153 ) );
  AOI22_X1 u2_u8_u1_U13 (.B2( u2_u8_u1_n136 ) , .A2( u2_u8_u1_n137 ) , .ZN( u2_u8_u1_n143 ) , .A1( u2_u8_u1_n171 ) , .B1( u2_u8_u1_n173 ) );
  INV_X1 u2_u8_u1_U14 (.A( u2_u8_u1_n147 ) , .ZN( u2_u8_u1_n181 ) );
  INV_X1 u2_u8_u1_U15 (.A( u2_u8_u1_n139 ) , .ZN( u2_u8_u1_n174 ) );
  OR4_X1 u2_u8_u1_U16 (.A4( u2_u8_u1_n106 ) , .A3( u2_u8_u1_n107 ) , .ZN( u2_u8_u1_n108 ) , .A1( u2_u8_u1_n117 ) , .A2( u2_u8_u1_n184 ) );
  AOI21_X1 u2_u8_u1_U17 (.ZN( u2_u8_u1_n106 ) , .A( u2_u8_u1_n112 ) , .B1( u2_u8_u1_n154 ) , .B2( u2_u8_u1_n156 ) );
  AOI21_X1 u2_u8_u1_U18 (.ZN( u2_u8_u1_n107 ) , .B1( u2_u8_u1_n134 ) , .B2( u2_u8_u1_n149 ) , .A( u2_u8_u1_n174 ) );
  INV_X1 u2_u8_u1_U19 (.A( u2_u8_u1_n101 ) , .ZN( u2_u8_u1_n184 ) );
  INV_X1 u2_u8_u1_U20 (.A( u2_u8_u1_n112 ) , .ZN( u2_u8_u1_n171 ) );
  NAND2_X1 u2_u8_u1_U21 (.ZN( u2_u8_u1_n141 ) , .A1( u2_u8_u1_n153 ) , .A2( u2_u8_u1_n156 ) );
  AND2_X1 u2_u8_u1_U22 (.A1( u2_u8_u1_n123 ) , .ZN( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n161 ) );
  NAND2_X1 u2_u8_u1_U23 (.A2( u2_u8_u1_n115 ) , .A1( u2_u8_u1_n116 ) , .ZN( u2_u8_u1_n148 ) );
  NAND2_X1 u2_u8_u1_U24 (.A2( u2_u8_u1_n133 ) , .A1( u2_u8_u1_n135 ) , .ZN( u2_u8_u1_n159 ) );
  NAND2_X1 u2_u8_u1_U25 (.A2( u2_u8_u1_n115 ) , .A1( u2_u8_u1_n120 ) , .ZN( u2_u8_u1_n132 ) );
  INV_X1 u2_u8_u1_U26 (.A( u2_u8_u1_n154 ) , .ZN( u2_u8_u1_n178 ) );
  INV_X1 u2_u8_u1_U27 (.A( u2_u8_u1_n151 ) , .ZN( u2_u8_u1_n183 ) );
  AND2_X1 u2_u8_u1_U28 (.A1( u2_u8_u1_n129 ) , .A2( u2_u8_u1_n133 ) , .ZN( u2_u8_u1_n149 ) );
  INV_X1 u2_u8_u1_U29 (.A( u2_u8_u1_n131 ) , .ZN( u2_u8_u1_n180 ) );
  INV_X1 u2_u8_u1_U3 (.A( u2_u8_u1_n159 ) , .ZN( u2_u8_u1_n182 ) );
  AOI221_X1 u2_u8_u1_U30 (.B1( u2_u8_u1_n140 ) , .ZN( u2_u8_u1_n167 ) , .B2( u2_u8_u1_n172 ) , .C2( u2_u8_u1_n175 ) , .C1( u2_u8_u1_n178 ) , .A( u2_u8_u1_n188 ) );
  INV_X1 u2_u8_u1_U31 (.ZN( u2_u8_u1_n188 ) , .A( u2_u8_u1_n97 ) );
  AOI211_X1 u2_u8_u1_U32 (.A( u2_u8_u1_n118 ) , .C1( u2_u8_u1_n132 ) , .C2( u2_u8_u1_n139 ) , .B( u2_u8_u1_n96 ) , .ZN( u2_u8_u1_n97 ) );
  AOI21_X1 u2_u8_u1_U33 (.B2( u2_u8_u1_n121 ) , .B1( u2_u8_u1_n135 ) , .A( u2_u8_u1_n152 ) , .ZN( u2_u8_u1_n96 ) );
  OAI221_X1 u2_u8_u1_U34 (.A( u2_u8_u1_n119 ) , .C2( u2_u8_u1_n129 ) , .ZN( u2_u8_u1_n138 ) , .B2( u2_u8_u1_n152 ) , .C1( u2_u8_u1_n174 ) , .B1( u2_u8_u1_n187 ) );
  INV_X1 u2_u8_u1_U35 (.A( u2_u8_u1_n148 ) , .ZN( u2_u8_u1_n187 ) );
  AOI211_X1 u2_u8_u1_U36 (.B( u2_u8_u1_n117 ) , .A( u2_u8_u1_n118 ) , .ZN( u2_u8_u1_n119 ) , .C2( u2_u8_u1_n146 ) , .C1( u2_u8_u1_n159 ) );
  NOR2_X1 u2_u8_u1_U37 (.A1( u2_u8_u1_n168 ) , .A2( u2_u8_u1_n176 ) , .ZN( u2_u8_u1_n98 ) );
  AOI211_X1 u2_u8_u1_U38 (.B( u2_u8_u1_n162 ) , .A( u2_u8_u1_n163 ) , .C2( u2_u8_u1_n164 ) , .ZN( u2_u8_u1_n165 ) , .C1( u2_u8_u1_n171 ) );
  AOI21_X1 u2_u8_u1_U39 (.A( u2_u8_u1_n160 ) , .B2( u2_u8_u1_n161 ) , .ZN( u2_u8_u1_n162 ) , .B1( u2_u8_u1_n182 ) );
  AOI221_X1 u2_u8_u1_U4 (.A( u2_u8_u1_n138 ) , .C2( u2_u8_u1_n139 ) , .C1( u2_u8_u1_n140 ) , .B2( u2_u8_u1_n141 ) , .ZN( u2_u8_u1_n142 ) , .B1( u2_u8_u1_n175 ) );
  OR2_X1 u2_u8_u1_U40 (.A2( u2_u8_u1_n157 ) , .A1( u2_u8_u1_n158 ) , .ZN( u2_u8_u1_n163 ) );
  NAND2_X1 u2_u8_u1_U41 (.A1( u2_u8_u1_n128 ) , .ZN( u2_u8_u1_n146 ) , .A2( u2_u8_u1_n160 ) );
  NAND2_X1 u2_u8_u1_U42 (.A2( u2_u8_u1_n112 ) , .ZN( u2_u8_u1_n139 ) , .A1( u2_u8_u1_n152 ) );
  NAND2_X1 u2_u8_u1_U43 (.A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n156 ) , .A2( u2_u8_u1_n99 ) );
  NOR2_X1 u2_u8_u1_U44 (.ZN( u2_u8_u1_n117 ) , .A1( u2_u8_u1_n121 ) , .A2( u2_u8_u1_n160 ) );
  OAI21_X1 u2_u8_u1_U45 (.B2( u2_u8_u1_n123 ) , .ZN( u2_u8_u1_n145 ) , .B1( u2_u8_u1_n160 ) , .A( u2_u8_u1_n185 ) );
  INV_X1 u2_u8_u1_U46 (.A( u2_u8_u1_n122 ) , .ZN( u2_u8_u1_n185 ) );
  AOI21_X1 u2_u8_u1_U47 (.B2( u2_u8_u1_n120 ) , .B1( u2_u8_u1_n121 ) , .ZN( u2_u8_u1_n122 ) , .A( u2_u8_u1_n128 ) );
  AOI21_X1 u2_u8_u1_U48 (.A( u2_u8_u1_n128 ) , .B2( u2_u8_u1_n129 ) , .ZN( u2_u8_u1_n130 ) , .B1( u2_u8_u1_n150 ) );
  NAND2_X1 u2_u8_u1_U49 (.ZN( u2_u8_u1_n112 ) , .A1( u2_u8_u1_n169 ) , .A2( u2_u8_u1_n170 ) );
  AOI211_X1 u2_u8_u1_U5 (.ZN( u2_u8_u1_n124 ) , .A( u2_u8_u1_n138 ) , .C2( u2_u8_u1_n139 ) , .B( u2_u8_u1_n145 ) , .C1( u2_u8_u1_n147 ) );
  NAND2_X1 u2_u8_u1_U50 (.ZN( u2_u8_u1_n129 ) , .A2( u2_u8_u1_n95 ) , .A1( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U51 (.A1( u2_u8_u1_n102 ) , .ZN( u2_u8_u1_n154 ) , .A2( u2_u8_u1_n99 ) );
  NAND2_X1 u2_u8_u1_U52 (.A2( u2_u8_u1_n100 ) , .ZN( u2_u8_u1_n135 ) , .A1( u2_u8_u1_n99 ) );
  AOI21_X1 u2_u8_u1_U53 (.A( u2_u8_u1_n152 ) , .B2( u2_u8_u1_n153 ) , .B1( u2_u8_u1_n154 ) , .ZN( u2_u8_u1_n158 ) );
  INV_X1 u2_u8_u1_U54 (.A( u2_u8_u1_n160 ) , .ZN( u2_u8_u1_n175 ) );
  NAND2_X1 u2_u8_u1_U55 (.A1( u2_u8_u1_n100 ) , .ZN( u2_u8_u1_n116 ) , .A2( u2_u8_u1_n95 ) );
  NAND2_X1 u2_u8_u1_U56 (.A1( u2_u8_u1_n102 ) , .ZN( u2_u8_u1_n131 ) , .A2( u2_u8_u1_n95 ) );
  NAND2_X1 u2_u8_u1_U57 (.A2( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n121 ) , .A1( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U58 (.A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n153 ) , .A2( u2_u8_u1_n98 ) );
  NAND2_X1 u2_u8_u1_U59 (.A2( u2_u8_u1_n104 ) , .A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n133 ) );
  AOI22_X1 u2_u8_u1_U6 (.B2( u2_u8_u1_n113 ) , .A2( u2_u8_u1_n114 ) , .ZN( u2_u8_u1_n125 ) , .A1( u2_u8_u1_n171 ) , .B1( u2_u8_u1_n173 ) );
  NAND2_X1 u2_u8_u1_U60 (.ZN( u2_u8_u1_n150 ) , .A2( u2_u8_u1_n98 ) , .A1( u2_u8_u1_n99 ) );
  NAND2_X1 u2_u8_u1_U61 (.A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n155 ) , .A2( u2_u8_u1_n95 ) );
  OAI21_X1 u2_u8_u1_U62 (.ZN( u2_u8_u1_n109 ) , .B1( u2_u8_u1_n129 ) , .B2( u2_u8_u1_n160 ) , .A( u2_u8_u1_n167 ) );
  NAND2_X1 u2_u8_u1_U63 (.A2( u2_u8_u1_n100 ) , .A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n120 ) );
  NAND2_X1 u2_u8_u1_U64 (.A1( u2_u8_u1_n102 ) , .A2( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n115 ) );
  NAND2_X1 u2_u8_u1_U65 (.A2( u2_u8_u1_n100 ) , .A1( u2_u8_u1_n104 ) , .ZN( u2_u8_u1_n151 ) );
  NAND2_X1 u2_u8_u1_U66 (.A2( u2_u8_u1_n103 ) , .A1( u2_u8_u1_n105 ) , .ZN( u2_u8_u1_n161 ) );
  INV_X1 u2_u8_u1_U67 (.A( u2_u8_u1_n152 ) , .ZN( u2_u8_u1_n173 ) );
  INV_X1 u2_u8_u1_U68 (.A( u2_u8_u1_n128 ) , .ZN( u2_u8_u1_n172 ) );
  NAND2_X1 u2_u8_u1_U69 (.A2( u2_u8_u1_n102 ) , .A1( u2_u8_u1_n103 ) , .ZN( u2_u8_u1_n123 ) );
  NAND2_X1 u2_u8_u1_U7 (.ZN( u2_u8_u1_n114 ) , .A1( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n156 ) );
  NOR2_X1 u2_u8_u1_U70 (.A2( u2_u8_X_7 ) , .A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n95 ) );
  NOR2_X1 u2_u8_u1_U71 (.A1( u2_u8_X_12 ) , .A2( u2_u8_X_9 ) , .ZN( u2_u8_u1_n100 ) );
  NOR2_X1 u2_u8_u1_U72 (.A2( u2_u8_X_8 ) , .A1( u2_u8_u1_n177 ) , .ZN( u2_u8_u1_n99 ) );
  NOR2_X1 u2_u8_u1_U73 (.A2( u2_u8_X_12 ) , .ZN( u2_u8_u1_n102 ) , .A1( u2_u8_u1_n176 ) );
  NOR2_X1 u2_u8_u1_U74 (.A2( u2_u8_X_9 ) , .ZN( u2_u8_u1_n105 ) , .A1( u2_u8_u1_n168 ) );
  NAND2_X1 u2_u8_u1_U75 (.A1( u2_u8_X_10 ) , .ZN( u2_u8_u1_n160 ) , .A2( u2_u8_u1_n169 ) );
  NAND2_X1 u2_u8_u1_U76 (.A2( u2_u8_X_10 ) , .A1( u2_u8_X_11 ) , .ZN( u2_u8_u1_n152 ) );
  NAND2_X1 u2_u8_u1_U77 (.A1( u2_u8_X_11 ) , .ZN( u2_u8_u1_n128 ) , .A2( u2_u8_u1_n170 ) );
  AND2_X1 u2_u8_u1_U78 (.A2( u2_u8_X_7 ) , .A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n104 ) );
  AND2_X1 u2_u8_u1_U79 (.A1( u2_u8_X_8 ) , .ZN( u2_u8_u1_n103 ) , .A2( u2_u8_u1_n177 ) );
  NOR2_X1 u2_u8_u1_U8 (.A1( u2_u8_u1_n112 ) , .A2( u2_u8_u1_n116 ) , .ZN( u2_u8_u1_n118 ) );
  INV_X1 u2_u8_u1_U80 (.A( u2_u8_X_10 ) , .ZN( u2_u8_u1_n170 ) );
  INV_X1 u2_u8_u1_U81 (.A( u2_u8_X_9 ) , .ZN( u2_u8_u1_n176 ) );
  INV_X1 u2_u8_u1_U82 (.A( u2_u8_X_11 ) , .ZN( u2_u8_u1_n169 ) );
  INV_X1 u2_u8_u1_U83 (.A( u2_u8_X_12 ) , .ZN( u2_u8_u1_n168 ) );
  INV_X1 u2_u8_u1_U84 (.A( u2_u8_X_7 ) , .ZN( u2_u8_u1_n177 ) );
  NAND4_X1 u2_u8_u1_U85 (.ZN( u2_out8_28 ) , .A4( u2_u8_u1_n124 ) , .A3( u2_u8_u1_n125 ) , .A2( u2_u8_u1_n126 ) , .A1( u2_u8_u1_n127 ) );
  OAI21_X1 u2_u8_u1_U86 (.ZN( u2_u8_u1_n127 ) , .B2( u2_u8_u1_n139 ) , .B1( u2_u8_u1_n175 ) , .A( u2_u8_u1_n183 ) );
  OAI21_X1 u2_u8_u1_U87 (.ZN( u2_u8_u1_n126 ) , .B2( u2_u8_u1_n140 ) , .A( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n178 ) );
  NAND4_X1 u2_u8_u1_U88 (.ZN( u2_out8_18 ) , .A4( u2_u8_u1_n165 ) , .A3( u2_u8_u1_n166 ) , .A1( u2_u8_u1_n167 ) , .A2( u2_u8_u1_n186 ) );
  AOI22_X1 u2_u8_u1_U89 (.B2( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n147 ) , .A2( u2_u8_u1_n148 ) , .ZN( u2_u8_u1_n166 ) , .A1( u2_u8_u1_n172 ) );
  OAI21_X1 u2_u8_u1_U9 (.ZN( u2_u8_u1_n101 ) , .B1( u2_u8_u1_n141 ) , .A( u2_u8_u1_n146 ) , .B2( u2_u8_u1_n183 ) );
  INV_X1 u2_u8_u1_U90 (.A( u2_u8_u1_n145 ) , .ZN( u2_u8_u1_n186 ) );
  NAND4_X1 u2_u8_u1_U91 (.ZN( u2_out8_2 ) , .A4( u2_u8_u1_n142 ) , .A3( u2_u8_u1_n143 ) , .A2( u2_u8_u1_n144 ) , .A1( u2_u8_u1_n179 ) );
  OAI21_X1 u2_u8_u1_U92 (.B2( u2_u8_u1_n132 ) , .ZN( u2_u8_u1_n144 ) , .A( u2_u8_u1_n146 ) , .B1( u2_u8_u1_n180 ) );
  INV_X1 u2_u8_u1_U93 (.A( u2_u8_u1_n130 ) , .ZN( u2_u8_u1_n179 ) );
  OR4_X1 u2_u8_u1_U94 (.ZN( u2_out8_13 ) , .A4( u2_u8_u1_n108 ) , .A3( u2_u8_u1_n109 ) , .A2( u2_u8_u1_n110 ) , .A1( u2_u8_u1_n111 ) );
  AOI21_X1 u2_u8_u1_U95 (.ZN( u2_u8_u1_n111 ) , .A( u2_u8_u1_n128 ) , .B2( u2_u8_u1_n131 ) , .B1( u2_u8_u1_n135 ) );
  AOI21_X1 u2_u8_u1_U96 (.ZN( u2_u8_u1_n110 ) , .A( u2_u8_u1_n116 ) , .B1( u2_u8_u1_n152 ) , .B2( u2_u8_u1_n160 ) );
  NAND3_X1 u2_u8_u1_U97 (.A3( u2_u8_u1_n149 ) , .A2( u2_u8_u1_n150 ) , .A1( u2_u8_u1_n151 ) , .ZN( u2_u8_u1_n164 ) );
  NAND3_X1 u2_u8_u1_U98 (.A3( u2_u8_u1_n134 ) , .A2( u2_u8_u1_n135 ) , .ZN( u2_u8_u1_n136 ) , .A1( u2_u8_u1_n151 ) );
  NAND3_X1 u2_u8_u1_U99 (.A1( u2_u8_u1_n133 ) , .ZN( u2_u8_u1_n137 ) , .A2( u2_u8_u1_n154 ) , .A3( u2_u8_u1_n181 ) );
  OAI22_X1 u2_u8_u2_U10 (.B1( u2_u8_u2_n151 ) , .A2( u2_u8_u2_n152 ) , .A1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n160 ) , .B2( u2_u8_u2_n168 ) );
  NAND3_X1 u2_u8_u2_U100 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n98 ) );
  NOR3_X1 u2_u8_u2_U11 (.A1( u2_u8_u2_n150 ) , .ZN( u2_u8_u2_n151 ) , .A3( u2_u8_u2_n175 ) , .A2( u2_u8_u2_n188 ) );
  AOI21_X1 u2_u8_u2_U12 (.B2( u2_u8_u2_n123 ) , .ZN( u2_u8_u2_n125 ) , .A( u2_u8_u2_n171 ) , .B1( u2_u8_u2_n184 ) );
  INV_X1 u2_u8_u2_U13 (.A( u2_u8_u2_n150 ) , .ZN( u2_u8_u2_n184 ) );
  AOI21_X1 u2_u8_u2_U14 (.ZN( u2_u8_u2_n144 ) , .B2( u2_u8_u2_n155 ) , .A( u2_u8_u2_n172 ) , .B1( u2_u8_u2_n185 ) );
  AOI21_X1 u2_u8_u2_U15 (.B2( u2_u8_u2_n143 ) , .ZN( u2_u8_u2_n145 ) , .B1( u2_u8_u2_n152 ) , .A( u2_u8_u2_n171 ) );
  INV_X1 u2_u8_u2_U16 (.A( u2_u8_u2_n156 ) , .ZN( u2_u8_u2_n171 ) );
  INV_X1 u2_u8_u2_U17 (.A( u2_u8_u2_n120 ) , .ZN( u2_u8_u2_n188 ) );
  NAND2_X1 u2_u8_u2_U18 (.A2( u2_u8_u2_n122 ) , .ZN( u2_u8_u2_n150 ) , .A1( u2_u8_u2_n152 ) );
  INV_X1 u2_u8_u2_U19 (.A( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n170 ) );
  INV_X1 u2_u8_u2_U20 (.A( u2_u8_u2_n137 ) , .ZN( u2_u8_u2_n173 ) );
  NAND2_X1 u2_u8_u2_U21 (.A1( u2_u8_u2_n132 ) , .A2( u2_u8_u2_n139 ) , .ZN( u2_u8_u2_n157 ) );
  INV_X1 u2_u8_u2_U22 (.A( u2_u8_u2_n113 ) , .ZN( u2_u8_u2_n178 ) );
  INV_X1 u2_u8_u2_U23 (.A( u2_u8_u2_n139 ) , .ZN( u2_u8_u2_n175 ) );
  INV_X1 u2_u8_u2_U24 (.A( u2_u8_u2_n155 ) , .ZN( u2_u8_u2_n181 ) );
  INV_X1 u2_u8_u2_U25 (.A( u2_u8_u2_n119 ) , .ZN( u2_u8_u2_n177 ) );
  INV_X1 u2_u8_u2_U26 (.A( u2_u8_u2_n116 ) , .ZN( u2_u8_u2_n180 ) );
  INV_X1 u2_u8_u2_U27 (.A( u2_u8_u2_n131 ) , .ZN( u2_u8_u2_n179 ) );
  INV_X1 u2_u8_u2_U28 (.A( u2_u8_u2_n154 ) , .ZN( u2_u8_u2_n176 ) );
  NAND2_X1 u2_u8_u2_U29 (.A2( u2_u8_u2_n116 ) , .A1( u2_u8_u2_n117 ) , .ZN( u2_u8_u2_n118 ) );
  NOR2_X1 u2_u8_u2_U3 (.ZN( u2_u8_u2_n121 ) , .A2( u2_u8_u2_n177 ) , .A1( u2_u8_u2_n180 ) );
  INV_X1 u2_u8_u2_U30 (.A( u2_u8_u2_n132 ) , .ZN( u2_u8_u2_n182 ) );
  INV_X1 u2_u8_u2_U31 (.A( u2_u8_u2_n158 ) , .ZN( u2_u8_u2_n183 ) );
  OAI21_X1 u2_u8_u2_U32 (.A( u2_u8_u2_n156 ) , .B1( u2_u8_u2_n157 ) , .ZN( u2_u8_u2_n158 ) , .B2( u2_u8_u2_n179 ) );
  NOR2_X1 u2_u8_u2_U33 (.ZN( u2_u8_u2_n156 ) , .A1( u2_u8_u2_n166 ) , .A2( u2_u8_u2_n169 ) );
  NOR2_X1 u2_u8_u2_U34 (.A2( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n137 ) , .A1( u2_u8_u2_n140 ) );
  NOR2_X1 u2_u8_u2_U35 (.A2( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n153 ) , .A1( u2_u8_u2_n156 ) );
  AOI211_X1 u2_u8_u2_U36 (.ZN( u2_u8_u2_n130 ) , .C1( u2_u8_u2_n138 ) , .C2( u2_u8_u2_n179 ) , .B( u2_u8_u2_n96 ) , .A( u2_u8_u2_n97 ) );
  OAI22_X1 u2_u8_u2_U37 (.B1( u2_u8_u2_n133 ) , .A2( u2_u8_u2_n137 ) , .A1( u2_u8_u2_n152 ) , .B2( u2_u8_u2_n168 ) , .ZN( u2_u8_u2_n97 ) );
  OAI221_X1 u2_u8_u2_U38 (.B1( u2_u8_u2_n113 ) , .C1( u2_u8_u2_n132 ) , .A( u2_u8_u2_n149 ) , .B2( u2_u8_u2_n171 ) , .C2( u2_u8_u2_n172 ) , .ZN( u2_u8_u2_n96 ) );
  OAI221_X1 u2_u8_u2_U39 (.A( u2_u8_u2_n115 ) , .C2( u2_u8_u2_n123 ) , .B2( u2_u8_u2_n143 ) , .B1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n163 ) , .C1( u2_u8_u2_n168 ) );
  INV_X1 u2_u8_u2_U4 (.A( u2_u8_u2_n134 ) , .ZN( u2_u8_u2_n185 ) );
  OAI21_X1 u2_u8_u2_U40 (.A( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n115 ) , .B1( u2_u8_u2_n176 ) , .B2( u2_u8_u2_n178 ) );
  OAI221_X1 u2_u8_u2_U41 (.A( u2_u8_u2_n135 ) , .B2( u2_u8_u2_n136 ) , .B1( u2_u8_u2_n137 ) , .ZN( u2_u8_u2_n162 ) , .C2( u2_u8_u2_n167 ) , .C1( u2_u8_u2_n185 ) );
  AND3_X1 u2_u8_u2_U42 (.A3( u2_u8_u2_n131 ) , .A2( u2_u8_u2_n132 ) , .A1( u2_u8_u2_n133 ) , .ZN( u2_u8_u2_n136 ) );
  AOI22_X1 u2_u8_u2_U43 (.ZN( u2_u8_u2_n135 ) , .B1( u2_u8_u2_n140 ) , .A1( u2_u8_u2_n156 ) , .B2( u2_u8_u2_n180 ) , .A2( u2_u8_u2_n188 ) );
  AOI21_X1 u2_u8_u2_U44 (.ZN( u2_u8_u2_n149 ) , .B1( u2_u8_u2_n173 ) , .B2( u2_u8_u2_n188 ) , .A( u2_u8_u2_n95 ) );
  AND3_X1 u2_u8_u2_U45 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n156 ) , .ZN( u2_u8_u2_n95 ) );
  OAI21_X1 u2_u8_u2_U46 (.A( u2_u8_u2_n141 ) , .B2( u2_u8_u2_n142 ) , .ZN( u2_u8_u2_n146 ) , .B1( u2_u8_u2_n153 ) );
  OAI21_X1 u2_u8_u2_U47 (.A( u2_u8_u2_n140 ) , .ZN( u2_u8_u2_n141 ) , .B1( u2_u8_u2_n176 ) , .B2( u2_u8_u2_n177 ) );
  NOR3_X1 u2_u8_u2_U48 (.ZN( u2_u8_u2_n142 ) , .A3( u2_u8_u2_n175 ) , .A2( u2_u8_u2_n178 ) , .A1( u2_u8_u2_n181 ) );
  OAI21_X1 u2_u8_u2_U49 (.A( u2_u8_u2_n101 ) , .B2( u2_u8_u2_n121 ) , .B1( u2_u8_u2_n153 ) , .ZN( u2_u8_u2_n164 ) );
  NOR4_X1 u2_u8_u2_U5 (.A4( u2_u8_u2_n124 ) , .A3( u2_u8_u2_n125 ) , .A2( u2_u8_u2_n126 ) , .A1( u2_u8_u2_n127 ) , .ZN( u2_u8_u2_n128 ) );
  NAND2_X1 u2_u8_u2_U50 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n155 ) );
  NAND2_X1 u2_u8_u2_U51 (.A2( u2_u8_u2_n105 ) , .A1( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n143 ) );
  NAND2_X1 u2_u8_u2_U52 (.A1( u2_u8_u2_n104 ) , .A2( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n152 ) );
  NAND2_X1 u2_u8_u2_U53 (.A1( u2_u8_u2_n100 ) , .A2( u2_u8_u2_n105 ) , .ZN( u2_u8_u2_n132 ) );
  INV_X1 u2_u8_u2_U54 (.A( u2_u8_u2_n140 ) , .ZN( u2_u8_u2_n168 ) );
  INV_X1 u2_u8_u2_U55 (.A( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n167 ) );
  NAND2_X1 u2_u8_u2_U56 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n113 ) );
  NAND2_X1 u2_u8_u2_U57 (.A1( u2_u8_u2_n106 ) , .A2( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n131 ) );
  NAND2_X1 u2_u8_u2_U58 (.A1( u2_u8_u2_n103 ) , .A2( u2_u8_u2_n107 ) , .ZN( u2_u8_u2_n139 ) );
  NAND2_X1 u2_u8_u2_U59 (.A1( u2_u8_u2_n103 ) , .A2( u2_u8_u2_n105 ) , .ZN( u2_u8_u2_n133 ) );
  AOI21_X1 u2_u8_u2_U6 (.B2( u2_u8_u2_n119 ) , .ZN( u2_u8_u2_n127 ) , .A( u2_u8_u2_n137 ) , .B1( u2_u8_u2_n155 ) );
  NAND2_X1 u2_u8_u2_U60 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n103 ) , .ZN( u2_u8_u2_n154 ) );
  NAND2_X1 u2_u8_u2_U61 (.A2( u2_u8_u2_n103 ) , .A1( u2_u8_u2_n104 ) , .ZN( u2_u8_u2_n119 ) );
  NAND2_X1 u2_u8_u2_U62 (.A2( u2_u8_u2_n107 ) , .A1( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n123 ) );
  NAND2_X1 u2_u8_u2_U63 (.A1( u2_u8_u2_n104 ) , .A2( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n122 ) );
  INV_X1 u2_u8_u2_U64 (.A( u2_u8_u2_n114 ) , .ZN( u2_u8_u2_n172 ) );
  NAND2_X1 u2_u8_u2_U65 (.A2( u2_u8_u2_n100 ) , .A1( u2_u8_u2_n102 ) , .ZN( u2_u8_u2_n116 ) );
  NAND2_X1 u2_u8_u2_U66 (.A1( u2_u8_u2_n102 ) , .A2( u2_u8_u2_n108 ) , .ZN( u2_u8_u2_n120 ) );
  NAND2_X1 u2_u8_u2_U67 (.A2( u2_u8_u2_n105 ) , .A1( u2_u8_u2_n106 ) , .ZN( u2_u8_u2_n117 ) );
  INV_X1 u2_u8_u2_U68 (.ZN( u2_u8_u2_n187 ) , .A( u2_u8_u2_n99 ) );
  OAI21_X1 u2_u8_u2_U69 (.B1( u2_u8_u2_n137 ) , .B2( u2_u8_u2_n143 ) , .A( u2_u8_u2_n98 ) , .ZN( u2_u8_u2_n99 ) );
  AOI21_X1 u2_u8_u2_U7 (.ZN( u2_u8_u2_n124 ) , .B1( u2_u8_u2_n131 ) , .B2( u2_u8_u2_n143 ) , .A( u2_u8_u2_n172 ) );
  NOR2_X1 u2_u8_u2_U70 (.A2( u2_u8_X_16 ) , .ZN( u2_u8_u2_n140 ) , .A1( u2_u8_u2_n166 ) );
  NOR2_X1 u2_u8_u2_U71 (.A2( u2_u8_X_13 ) , .A1( u2_u8_X_14 ) , .ZN( u2_u8_u2_n100 ) );
  NOR2_X1 u2_u8_u2_U72 (.A2( u2_u8_X_16 ) , .A1( u2_u8_X_17 ) , .ZN( u2_u8_u2_n138 ) );
  NOR2_X1 u2_u8_u2_U73 (.A2( u2_u8_X_15 ) , .A1( u2_u8_X_18 ) , .ZN( u2_u8_u2_n104 ) );
  NOR2_X1 u2_u8_u2_U74 (.A2( u2_u8_X_14 ) , .ZN( u2_u8_u2_n103 ) , .A1( u2_u8_u2_n174 ) );
  NOR2_X1 u2_u8_u2_U75 (.A2( u2_u8_X_15 ) , .ZN( u2_u8_u2_n102 ) , .A1( u2_u8_u2_n165 ) );
  NOR2_X1 u2_u8_u2_U76 (.A2( u2_u8_X_17 ) , .ZN( u2_u8_u2_n114 ) , .A1( u2_u8_u2_n169 ) );
  AND2_X1 u2_u8_u2_U77 (.A1( u2_u8_X_15 ) , .ZN( u2_u8_u2_n105 ) , .A2( u2_u8_u2_n165 ) );
  AND2_X1 u2_u8_u2_U78 (.A2( u2_u8_X_15 ) , .A1( u2_u8_X_18 ) , .ZN( u2_u8_u2_n107 ) );
  AND2_X1 u2_u8_u2_U79 (.A1( u2_u8_X_14 ) , .ZN( u2_u8_u2_n106 ) , .A2( u2_u8_u2_n174 ) );
  AOI21_X1 u2_u8_u2_U8 (.B2( u2_u8_u2_n120 ) , .B1( u2_u8_u2_n121 ) , .ZN( u2_u8_u2_n126 ) , .A( u2_u8_u2_n167 ) );
  AND2_X1 u2_u8_u2_U80 (.A1( u2_u8_X_13 ) , .A2( u2_u8_X_14 ) , .ZN( u2_u8_u2_n108 ) );
  INV_X1 u2_u8_u2_U81 (.A( u2_u8_X_16 ) , .ZN( u2_u8_u2_n169 ) );
  INV_X1 u2_u8_u2_U82 (.A( u2_u8_X_17 ) , .ZN( u2_u8_u2_n166 ) );
  INV_X1 u2_u8_u2_U83 (.A( u2_u8_X_13 ) , .ZN( u2_u8_u2_n174 ) );
  INV_X1 u2_u8_u2_U84 (.A( u2_u8_X_18 ) , .ZN( u2_u8_u2_n165 ) );
  NAND4_X1 u2_u8_u2_U85 (.ZN( u2_out8_30 ) , .A4( u2_u8_u2_n147 ) , .A3( u2_u8_u2_n148 ) , .A2( u2_u8_u2_n149 ) , .A1( u2_u8_u2_n187 ) );
  NOR3_X1 u2_u8_u2_U86 (.A3( u2_u8_u2_n144 ) , .A2( u2_u8_u2_n145 ) , .A1( u2_u8_u2_n146 ) , .ZN( u2_u8_u2_n147 ) );
  AOI21_X1 u2_u8_u2_U87 (.B2( u2_u8_u2_n138 ) , .ZN( u2_u8_u2_n148 ) , .A( u2_u8_u2_n162 ) , .B1( u2_u8_u2_n182 ) );
  NAND4_X1 u2_u8_u2_U88 (.ZN( u2_out8_24 ) , .A4( u2_u8_u2_n111 ) , .A3( u2_u8_u2_n112 ) , .A1( u2_u8_u2_n130 ) , .A2( u2_u8_u2_n187 ) );
  AOI221_X1 u2_u8_u2_U89 (.A( u2_u8_u2_n109 ) , .B1( u2_u8_u2_n110 ) , .ZN( u2_u8_u2_n111 ) , .C1( u2_u8_u2_n134 ) , .C2( u2_u8_u2_n170 ) , .B2( u2_u8_u2_n173 ) );
  OAI22_X1 u2_u8_u2_U9 (.ZN( u2_u8_u2_n109 ) , .A2( u2_u8_u2_n113 ) , .B2( u2_u8_u2_n133 ) , .B1( u2_u8_u2_n167 ) , .A1( u2_u8_u2_n168 ) );
  AOI21_X1 u2_u8_u2_U90 (.ZN( u2_u8_u2_n112 ) , .B2( u2_u8_u2_n156 ) , .A( u2_u8_u2_n164 ) , .B1( u2_u8_u2_n181 ) );
  NAND4_X1 u2_u8_u2_U91 (.ZN( u2_out8_16 ) , .A4( u2_u8_u2_n128 ) , .A3( u2_u8_u2_n129 ) , .A1( u2_u8_u2_n130 ) , .A2( u2_u8_u2_n186 ) );
  AOI22_X1 u2_u8_u2_U92 (.A2( u2_u8_u2_n118 ) , .ZN( u2_u8_u2_n129 ) , .A1( u2_u8_u2_n140 ) , .B1( u2_u8_u2_n157 ) , .B2( u2_u8_u2_n170 ) );
  INV_X1 u2_u8_u2_U93 (.A( u2_u8_u2_n163 ) , .ZN( u2_u8_u2_n186 ) );
  OR4_X1 u2_u8_u2_U94 (.ZN( u2_out8_6 ) , .A4( u2_u8_u2_n161 ) , .A3( u2_u8_u2_n162 ) , .A2( u2_u8_u2_n163 ) , .A1( u2_u8_u2_n164 ) );
  OR3_X1 u2_u8_u2_U95 (.A2( u2_u8_u2_n159 ) , .A1( u2_u8_u2_n160 ) , .ZN( u2_u8_u2_n161 ) , .A3( u2_u8_u2_n183 ) );
  AOI21_X1 u2_u8_u2_U96 (.B2( u2_u8_u2_n154 ) , .B1( u2_u8_u2_n155 ) , .ZN( u2_u8_u2_n159 ) , .A( u2_u8_u2_n167 ) );
  NAND3_X1 u2_u8_u2_U97 (.A2( u2_u8_u2_n117 ) , .A1( u2_u8_u2_n122 ) , .A3( u2_u8_u2_n123 ) , .ZN( u2_u8_u2_n134 ) );
  NAND3_X1 u2_u8_u2_U98 (.ZN( u2_u8_u2_n110 ) , .A2( u2_u8_u2_n131 ) , .A3( u2_u8_u2_n139 ) , .A1( u2_u8_u2_n154 ) );
  NAND3_X1 u2_u8_u2_U99 (.A2( u2_u8_u2_n100 ) , .ZN( u2_u8_u2_n101 ) , .A1( u2_u8_u2_n104 ) , .A3( u2_u8_u2_n114 ) );
  OAI22_X1 u2_u8_u3_U10 (.B1( u2_u8_u3_n113 ) , .A2( u2_u8_u3_n135 ) , .A1( u2_u8_u3_n150 ) , .B2( u2_u8_u3_n164 ) , .ZN( u2_u8_u3_n98 ) );
  OAI211_X1 u2_u8_u3_U11 (.B( u2_u8_u3_n106 ) , .ZN( u2_u8_u3_n119 ) , .C2( u2_u8_u3_n128 ) , .C1( u2_u8_u3_n167 ) , .A( u2_u8_u3_n181 ) );
  AOI221_X1 u2_u8_u3_U12 (.C1( u2_u8_u3_n105 ) , .ZN( u2_u8_u3_n106 ) , .A( u2_u8_u3_n131 ) , .B2( u2_u8_u3_n132 ) , .C2( u2_u8_u3_n133 ) , .B1( u2_u8_u3_n169 ) );
  INV_X1 u2_u8_u3_U13 (.ZN( u2_u8_u3_n181 ) , .A( u2_u8_u3_n98 ) );
  NAND2_X1 u2_u8_u3_U14 (.ZN( u2_u8_u3_n105 ) , .A2( u2_u8_u3_n130 ) , .A1( u2_u8_u3_n155 ) );
  AOI22_X1 u2_u8_u3_U15 (.B1( u2_u8_u3_n115 ) , .A2( u2_u8_u3_n116 ) , .ZN( u2_u8_u3_n123 ) , .B2( u2_u8_u3_n133 ) , .A1( u2_u8_u3_n169 ) );
  NAND2_X1 u2_u8_u3_U16 (.ZN( u2_u8_u3_n116 ) , .A2( u2_u8_u3_n151 ) , .A1( u2_u8_u3_n182 ) );
  NOR2_X1 u2_u8_u3_U17 (.ZN( u2_u8_u3_n126 ) , .A2( u2_u8_u3_n150 ) , .A1( u2_u8_u3_n164 ) );
  AOI21_X1 u2_u8_u3_U18 (.ZN( u2_u8_u3_n112 ) , .B2( u2_u8_u3_n146 ) , .B1( u2_u8_u3_n155 ) , .A( u2_u8_u3_n167 ) );
  NAND2_X1 u2_u8_u3_U19 (.A1( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n142 ) , .A2( u2_u8_u3_n164 ) );
  NAND2_X1 u2_u8_u3_U20 (.ZN( u2_u8_u3_n132 ) , .A2( u2_u8_u3_n152 ) , .A1( u2_u8_u3_n156 ) );
  AND2_X1 u2_u8_u3_U21 (.A2( u2_u8_u3_n113 ) , .A1( u2_u8_u3_n114 ) , .ZN( u2_u8_u3_n151 ) );
  INV_X1 u2_u8_u3_U22 (.A( u2_u8_u3_n133 ) , .ZN( u2_u8_u3_n165 ) );
  INV_X1 u2_u8_u3_U23 (.A( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n170 ) );
  NAND2_X1 u2_u8_u3_U24 (.A1( u2_u8_u3_n107 ) , .A2( u2_u8_u3_n108 ) , .ZN( u2_u8_u3_n140 ) );
  NAND2_X1 u2_u8_u3_U25 (.ZN( u2_u8_u3_n117 ) , .A1( u2_u8_u3_n124 ) , .A2( u2_u8_u3_n148 ) );
  NAND2_X1 u2_u8_u3_U26 (.ZN( u2_u8_u3_n143 ) , .A1( u2_u8_u3_n165 ) , .A2( u2_u8_u3_n167 ) );
  INV_X1 u2_u8_u3_U27 (.A( u2_u8_u3_n130 ) , .ZN( u2_u8_u3_n177 ) );
  INV_X1 u2_u8_u3_U28 (.A( u2_u8_u3_n128 ) , .ZN( u2_u8_u3_n176 ) );
  INV_X1 u2_u8_u3_U29 (.A( u2_u8_u3_n155 ) , .ZN( u2_u8_u3_n174 ) );
  INV_X1 u2_u8_u3_U3 (.A( u2_u8_u3_n129 ) , .ZN( u2_u8_u3_n183 ) );
  INV_X1 u2_u8_u3_U30 (.A( u2_u8_u3_n139 ) , .ZN( u2_u8_u3_n185 ) );
  NOR2_X1 u2_u8_u3_U31 (.ZN( u2_u8_u3_n135 ) , .A2( u2_u8_u3_n141 ) , .A1( u2_u8_u3_n169 ) );
  OAI222_X1 u2_u8_u3_U32 (.C2( u2_u8_u3_n107 ) , .A2( u2_u8_u3_n108 ) , .B1( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n138 ) , .B2( u2_u8_u3_n146 ) , .C1( u2_u8_u3_n154 ) , .A1( u2_u8_u3_n164 ) );
  NOR4_X1 u2_u8_u3_U33 (.A4( u2_u8_u3_n157 ) , .A3( u2_u8_u3_n158 ) , .A2( u2_u8_u3_n159 ) , .A1( u2_u8_u3_n160 ) , .ZN( u2_u8_u3_n161 ) );
  AOI21_X1 u2_u8_u3_U34 (.B2( u2_u8_u3_n152 ) , .B1( u2_u8_u3_n153 ) , .ZN( u2_u8_u3_n158 ) , .A( u2_u8_u3_n164 ) );
  AOI21_X1 u2_u8_u3_U35 (.A( u2_u8_u3_n149 ) , .B2( u2_u8_u3_n150 ) , .B1( u2_u8_u3_n151 ) , .ZN( u2_u8_u3_n159 ) );
  AOI21_X1 u2_u8_u3_U36 (.A( u2_u8_u3_n154 ) , .B2( u2_u8_u3_n155 ) , .B1( u2_u8_u3_n156 ) , .ZN( u2_u8_u3_n157 ) );
  AOI211_X1 u2_u8_u3_U37 (.ZN( u2_u8_u3_n109 ) , .A( u2_u8_u3_n119 ) , .C2( u2_u8_u3_n129 ) , .B( u2_u8_u3_n138 ) , .C1( u2_u8_u3_n141 ) );
  AOI211_X1 u2_u8_u3_U38 (.B( u2_u8_u3_n119 ) , .A( u2_u8_u3_n120 ) , .C2( u2_u8_u3_n121 ) , .ZN( u2_u8_u3_n122 ) , .C1( u2_u8_u3_n179 ) );
  INV_X1 u2_u8_u3_U39 (.A( u2_u8_u3_n156 ) , .ZN( u2_u8_u3_n179 ) );
  INV_X1 u2_u8_u3_U4 (.A( u2_u8_u3_n140 ) , .ZN( u2_u8_u3_n182 ) );
  OAI22_X1 u2_u8_u3_U40 (.B1( u2_u8_u3_n118 ) , .ZN( u2_u8_u3_n120 ) , .A1( u2_u8_u3_n135 ) , .B2( u2_u8_u3_n154 ) , .A2( u2_u8_u3_n178 ) );
  AND3_X1 u2_u8_u3_U41 (.ZN( u2_u8_u3_n118 ) , .A2( u2_u8_u3_n124 ) , .A1( u2_u8_u3_n144 ) , .A3( u2_u8_u3_n152 ) );
  INV_X1 u2_u8_u3_U42 (.A( u2_u8_u3_n121 ) , .ZN( u2_u8_u3_n164 ) );
  NAND2_X1 u2_u8_u3_U43 (.ZN( u2_u8_u3_n133 ) , .A1( u2_u8_u3_n154 ) , .A2( u2_u8_u3_n164 ) );
  OAI211_X1 u2_u8_u3_U44 (.B( u2_u8_u3_n127 ) , .ZN( u2_u8_u3_n139 ) , .C1( u2_u8_u3_n150 ) , .C2( u2_u8_u3_n154 ) , .A( u2_u8_u3_n184 ) );
  INV_X1 u2_u8_u3_U45 (.A( u2_u8_u3_n125 ) , .ZN( u2_u8_u3_n184 ) );
  AOI221_X1 u2_u8_u3_U46 (.A( u2_u8_u3_n126 ) , .ZN( u2_u8_u3_n127 ) , .C2( u2_u8_u3_n132 ) , .C1( u2_u8_u3_n169 ) , .B2( u2_u8_u3_n170 ) , .B1( u2_u8_u3_n174 ) );
  OAI22_X1 u2_u8_u3_U47 (.A1( u2_u8_u3_n124 ) , .ZN( u2_u8_u3_n125 ) , .B2( u2_u8_u3_n145 ) , .A2( u2_u8_u3_n165 ) , .B1( u2_u8_u3_n167 ) );
  NOR2_X1 u2_u8_u3_U48 (.A1( u2_u8_u3_n113 ) , .ZN( u2_u8_u3_n131 ) , .A2( u2_u8_u3_n154 ) );
  NAND2_X1 u2_u8_u3_U49 (.A1( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n150 ) , .A2( u2_u8_u3_n99 ) );
  INV_X1 u2_u8_u3_U5 (.A( u2_u8_u3_n117 ) , .ZN( u2_u8_u3_n178 ) );
  NAND2_X1 u2_u8_u3_U50 (.A2( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n155 ) , .A1( u2_u8_u3_n97 ) );
  INV_X1 u2_u8_u3_U51 (.A( u2_u8_u3_n141 ) , .ZN( u2_u8_u3_n167 ) );
  AOI21_X1 u2_u8_u3_U52 (.B2( u2_u8_u3_n114 ) , .B1( u2_u8_u3_n146 ) , .A( u2_u8_u3_n154 ) , .ZN( u2_u8_u3_n94 ) );
  AOI21_X1 u2_u8_u3_U53 (.ZN( u2_u8_u3_n110 ) , .B2( u2_u8_u3_n142 ) , .B1( u2_u8_u3_n186 ) , .A( u2_u8_u3_n95 ) );
  INV_X1 u2_u8_u3_U54 (.A( u2_u8_u3_n145 ) , .ZN( u2_u8_u3_n186 ) );
  AOI21_X1 u2_u8_u3_U55 (.B1( u2_u8_u3_n124 ) , .A( u2_u8_u3_n149 ) , .B2( u2_u8_u3_n155 ) , .ZN( u2_u8_u3_n95 ) );
  INV_X1 u2_u8_u3_U56 (.A( u2_u8_u3_n149 ) , .ZN( u2_u8_u3_n169 ) );
  NAND2_X1 u2_u8_u3_U57 (.ZN( u2_u8_u3_n124 ) , .A1( u2_u8_u3_n96 ) , .A2( u2_u8_u3_n97 ) );
  NAND2_X1 u2_u8_u3_U58 (.A2( u2_u8_u3_n100 ) , .ZN( u2_u8_u3_n146 ) , .A1( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U59 (.A1( u2_u8_u3_n101 ) , .ZN( u2_u8_u3_n145 ) , .A2( u2_u8_u3_n99 ) );
  AOI221_X1 u2_u8_u3_U6 (.A( u2_u8_u3_n131 ) , .C2( u2_u8_u3_n132 ) , .C1( u2_u8_u3_n133 ) , .ZN( u2_u8_u3_n134 ) , .B1( u2_u8_u3_n143 ) , .B2( u2_u8_u3_n177 ) );
  NAND2_X1 u2_u8_u3_U60 (.A1( u2_u8_u3_n100 ) , .ZN( u2_u8_u3_n156 ) , .A2( u2_u8_u3_n99 ) );
  NAND2_X1 u2_u8_u3_U61 (.A2( u2_u8_u3_n101 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n148 ) );
  NAND2_X1 u2_u8_u3_U62 (.A1( u2_u8_u3_n100 ) , .A2( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n128 ) );
  NAND2_X1 u2_u8_u3_U63 (.A2( u2_u8_u3_n101 ) , .A1( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n152 ) );
  NAND2_X1 u2_u8_u3_U64 (.A2( u2_u8_u3_n101 ) , .ZN( u2_u8_u3_n114 ) , .A1( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U65 (.ZN( u2_u8_u3_n107 ) , .A1( u2_u8_u3_n97 ) , .A2( u2_u8_u3_n99 ) );
  NAND2_X1 u2_u8_u3_U66 (.A2( u2_u8_u3_n100 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n113 ) );
  NAND2_X1 u2_u8_u3_U67 (.A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n153 ) , .A2( u2_u8_u3_n97 ) );
  NAND2_X1 u2_u8_u3_U68 (.A2( u2_u8_u3_n103 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n130 ) );
  NAND2_X1 u2_u8_u3_U69 (.A2( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n144 ) , .A1( u2_u8_u3_n96 ) );
  OAI22_X1 u2_u8_u3_U7 (.B2( u2_u8_u3_n147 ) , .A2( u2_u8_u3_n148 ) , .ZN( u2_u8_u3_n160 ) , .B1( u2_u8_u3_n165 ) , .A1( u2_u8_u3_n168 ) );
  NAND2_X1 u2_u8_u3_U70 (.A1( u2_u8_u3_n102 ) , .A2( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n108 ) );
  NOR2_X1 u2_u8_u3_U71 (.A2( u2_u8_X_19 ) , .A1( u2_u8_X_20 ) , .ZN( u2_u8_u3_n99 ) );
  NOR2_X1 u2_u8_u3_U72 (.A2( u2_u8_X_21 ) , .A1( u2_u8_X_24 ) , .ZN( u2_u8_u3_n103 ) );
  NOR2_X1 u2_u8_u3_U73 (.A2( u2_u8_X_24 ) , .A1( u2_u8_u3_n171 ) , .ZN( u2_u8_u3_n97 ) );
  NOR2_X1 u2_u8_u3_U74 (.A2( u2_u8_X_23 ) , .ZN( u2_u8_u3_n141 ) , .A1( u2_u8_u3_n166 ) );
  NOR2_X1 u2_u8_u3_U75 (.A2( u2_u8_X_19 ) , .A1( u2_u8_u3_n172 ) , .ZN( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U76 (.A1( u2_u8_X_22 ) , .A2( u2_u8_X_23 ) , .ZN( u2_u8_u3_n154 ) );
  NAND2_X1 u2_u8_u3_U77 (.A1( u2_u8_X_23 ) , .ZN( u2_u8_u3_n149 ) , .A2( u2_u8_u3_n166 ) );
  NOR2_X1 u2_u8_u3_U78 (.A2( u2_u8_X_22 ) , .A1( u2_u8_X_23 ) , .ZN( u2_u8_u3_n121 ) );
  AND2_X1 u2_u8_u3_U79 (.A1( u2_u8_X_24 ) , .ZN( u2_u8_u3_n101 ) , .A2( u2_u8_u3_n171 ) );
  AND3_X1 u2_u8_u3_U8 (.A3( u2_u8_u3_n144 ) , .A2( u2_u8_u3_n145 ) , .A1( u2_u8_u3_n146 ) , .ZN( u2_u8_u3_n147 ) );
  AND2_X1 u2_u8_u3_U80 (.A1( u2_u8_X_19 ) , .ZN( u2_u8_u3_n102 ) , .A2( u2_u8_u3_n172 ) );
  AND2_X1 u2_u8_u3_U81 (.A1( u2_u8_X_21 ) , .A2( u2_u8_X_24 ) , .ZN( u2_u8_u3_n100 ) );
  AND2_X1 u2_u8_u3_U82 (.A2( u2_u8_X_19 ) , .A1( u2_u8_X_20 ) , .ZN( u2_u8_u3_n104 ) );
  INV_X1 u2_u8_u3_U83 (.A( u2_u8_X_22 ) , .ZN( u2_u8_u3_n166 ) );
  INV_X1 u2_u8_u3_U84 (.A( u2_u8_X_21 ) , .ZN( u2_u8_u3_n171 ) );
  INV_X1 u2_u8_u3_U85 (.A( u2_u8_X_20 ) , .ZN( u2_u8_u3_n172 ) );
  OR4_X1 u2_u8_u3_U86 (.ZN( u2_out8_10 ) , .A4( u2_u8_u3_n136 ) , .A3( u2_u8_u3_n137 ) , .A1( u2_u8_u3_n138 ) , .A2( u2_u8_u3_n139 ) );
  OAI222_X1 u2_u8_u3_U87 (.C1( u2_u8_u3_n128 ) , .ZN( u2_u8_u3_n137 ) , .B1( u2_u8_u3_n148 ) , .A2( u2_u8_u3_n150 ) , .B2( u2_u8_u3_n154 ) , .C2( u2_u8_u3_n164 ) , .A1( u2_u8_u3_n167 ) );
  OAI221_X1 u2_u8_u3_U88 (.A( u2_u8_u3_n134 ) , .B2( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n136 ) , .C1( u2_u8_u3_n149 ) , .B1( u2_u8_u3_n151 ) , .C2( u2_u8_u3_n183 ) );
  NAND4_X1 u2_u8_u3_U89 (.ZN( u2_out8_26 ) , .A4( u2_u8_u3_n109 ) , .A3( u2_u8_u3_n110 ) , .A2( u2_u8_u3_n111 ) , .A1( u2_u8_u3_n173 ) );
  INV_X1 u2_u8_u3_U9 (.A( u2_u8_u3_n143 ) , .ZN( u2_u8_u3_n168 ) );
  INV_X1 u2_u8_u3_U90 (.ZN( u2_u8_u3_n173 ) , .A( u2_u8_u3_n94 ) );
  OAI21_X1 u2_u8_u3_U91 (.ZN( u2_u8_u3_n111 ) , .B2( u2_u8_u3_n117 ) , .A( u2_u8_u3_n133 ) , .B1( u2_u8_u3_n176 ) );
  NAND4_X1 u2_u8_u3_U92 (.ZN( u2_out8_20 ) , .A4( u2_u8_u3_n122 ) , .A3( u2_u8_u3_n123 ) , .A1( u2_u8_u3_n175 ) , .A2( u2_u8_u3_n180 ) );
  INV_X1 u2_u8_u3_U93 (.A( u2_u8_u3_n126 ) , .ZN( u2_u8_u3_n180 ) );
  INV_X1 u2_u8_u3_U94 (.A( u2_u8_u3_n112 ) , .ZN( u2_u8_u3_n175 ) );
  NAND4_X1 u2_u8_u3_U95 (.ZN( u2_out8_1 ) , .A4( u2_u8_u3_n161 ) , .A3( u2_u8_u3_n162 ) , .A2( u2_u8_u3_n163 ) , .A1( u2_u8_u3_n185 ) );
  NAND2_X1 u2_u8_u3_U96 (.ZN( u2_u8_u3_n163 ) , .A2( u2_u8_u3_n170 ) , .A1( u2_u8_u3_n176 ) );
  AOI22_X1 u2_u8_u3_U97 (.B2( u2_u8_u3_n140 ) , .B1( u2_u8_u3_n141 ) , .A2( u2_u8_u3_n142 ) , .ZN( u2_u8_u3_n162 ) , .A1( u2_u8_u3_n177 ) );
  NAND3_X1 u2_u8_u3_U98 (.A1( u2_u8_u3_n114 ) , .ZN( u2_u8_u3_n115 ) , .A2( u2_u8_u3_n145 ) , .A3( u2_u8_u3_n153 ) );
  NAND3_X1 u2_u8_u3_U99 (.ZN( u2_u8_u3_n129 ) , .A2( u2_u8_u3_n144 ) , .A1( u2_u8_u3_n153 ) , .A3( u2_u8_u3_n182 ) );
  OAI22_X1 u2_u8_u4_U10 (.B2( u2_u8_u4_n135 ) , .ZN( u2_u8_u4_n137 ) , .B1( u2_u8_u4_n153 ) , .A1( u2_u8_u4_n155 ) , .A2( u2_u8_u4_n171 ) );
  AND3_X1 u2_u8_u4_U11 (.A2( u2_u8_u4_n134 ) , .ZN( u2_u8_u4_n135 ) , .A3( u2_u8_u4_n145 ) , .A1( u2_u8_u4_n157 ) );
  NAND2_X1 u2_u8_u4_U12 (.ZN( u2_u8_u4_n132 ) , .A2( u2_u8_u4_n170 ) , .A1( u2_u8_u4_n173 ) );
  AOI21_X1 u2_u8_u4_U13 (.B2( u2_u8_u4_n160 ) , .B1( u2_u8_u4_n161 ) , .ZN( u2_u8_u4_n162 ) , .A( u2_u8_u4_n170 ) );
  AOI21_X1 u2_u8_u4_U14 (.ZN( u2_u8_u4_n107 ) , .B2( u2_u8_u4_n143 ) , .A( u2_u8_u4_n174 ) , .B1( u2_u8_u4_n184 ) );
  AOI21_X1 u2_u8_u4_U15 (.B2( u2_u8_u4_n158 ) , .B1( u2_u8_u4_n159 ) , .ZN( u2_u8_u4_n163 ) , .A( u2_u8_u4_n174 ) );
  AOI21_X1 u2_u8_u4_U16 (.A( u2_u8_u4_n153 ) , .B2( u2_u8_u4_n154 ) , .B1( u2_u8_u4_n155 ) , .ZN( u2_u8_u4_n165 ) );
  AOI21_X1 u2_u8_u4_U17 (.A( u2_u8_u4_n156 ) , .B2( u2_u8_u4_n157 ) , .ZN( u2_u8_u4_n164 ) , .B1( u2_u8_u4_n184 ) );
  INV_X1 u2_u8_u4_U18 (.A( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n170 ) );
  AND2_X1 u2_u8_u4_U19 (.A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n155 ) , .A1( u2_u8_u4_n160 ) );
  INV_X1 u2_u8_u4_U20 (.A( u2_u8_u4_n156 ) , .ZN( u2_u8_u4_n175 ) );
  NAND2_X1 u2_u8_u4_U21 (.A2( u2_u8_u4_n118 ) , .ZN( u2_u8_u4_n131 ) , .A1( u2_u8_u4_n147 ) );
  NAND2_X1 u2_u8_u4_U22 (.A1( u2_u8_u4_n119 ) , .A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n130 ) );
  NAND2_X1 u2_u8_u4_U23 (.ZN( u2_u8_u4_n117 ) , .A2( u2_u8_u4_n118 ) , .A1( u2_u8_u4_n148 ) );
  NAND2_X1 u2_u8_u4_U24 (.ZN( u2_u8_u4_n129 ) , .A1( u2_u8_u4_n134 ) , .A2( u2_u8_u4_n148 ) );
  AND3_X1 u2_u8_u4_U25 (.A1( u2_u8_u4_n119 ) , .A2( u2_u8_u4_n143 ) , .A3( u2_u8_u4_n154 ) , .ZN( u2_u8_u4_n161 ) );
  AND2_X1 u2_u8_u4_U26 (.A1( u2_u8_u4_n145 ) , .A2( u2_u8_u4_n147 ) , .ZN( u2_u8_u4_n159 ) );
  OR3_X1 u2_u8_u4_U27 (.A3( u2_u8_u4_n114 ) , .A2( u2_u8_u4_n115 ) , .A1( u2_u8_u4_n116 ) , .ZN( u2_u8_u4_n136 ) );
  AOI21_X1 u2_u8_u4_U28 (.A( u2_u8_u4_n113 ) , .ZN( u2_u8_u4_n116 ) , .B2( u2_u8_u4_n173 ) , .B1( u2_u8_u4_n174 ) );
  AOI21_X1 u2_u8_u4_U29 (.ZN( u2_u8_u4_n115 ) , .B2( u2_u8_u4_n145 ) , .B1( u2_u8_u4_n146 ) , .A( u2_u8_u4_n156 ) );
  NOR2_X1 u2_u8_u4_U3 (.ZN( u2_u8_u4_n121 ) , .A1( u2_u8_u4_n181 ) , .A2( u2_u8_u4_n182 ) );
  OAI22_X1 u2_u8_u4_U30 (.ZN( u2_u8_u4_n114 ) , .A2( u2_u8_u4_n121 ) , .B1( u2_u8_u4_n160 ) , .B2( u2_u8_u4_n170 ) , .A1( u2_u8_u4_n171 ) );
  INV_X1 u2_u8_u4_U31 (.A( u2_u8_u4_n158 ) , .ZN( u2_u8_u4_n182 ) );
  INV_X1 u2_u8_u4_U32 (.ZN( u2_u8_u4_n181 ) , .A( u2_u8_u4_n96 ) );
  INV_X1 u2_u8_u4_U33 (.A( u2_u8_u4_n144 ) , .ZN( u2_u8_u4_n179 ) );
  INV_X1 u2_u8_u4_U34 (.A( u2_u8_u4_n157 ) , .ZN( u2_u8_u4_n178 ) );
  NAND2_X1 u2_u8_u4_U35 (.A2( u2_u8_u4_n154 ) , .A1( u2_u8_u4_n96 ) , .ZN( u2_u8_u4_n97 ) );
  INV_X1 u2_u8_u4_U36 (.ZN( u2_u8_u4_n186 ) , .A( u2_u8_u4_n95 ) );
  OAI221_X1 u2_u8_u4_U37 (.C1( u2_u8_u4_n134 ) , .B1( u2_u8_u4_n158 ) , .B2( u2_u8_u4_n171 ) , .C2( u2_u8_u4_n173 ) , .A( u2_u8_u4_n94 ) , .ZN( u2_u8_u4_n95 ) );
  AOI222_X1 u2_u8_u4_U38 (.B2( u2_u8_u4_n132 ) , .A1( u2_u8_u4_n138 ) , .C2( u2_u8_u4_n175 ) , .A2( u2_u8_u4_n179 ) , .C1( u2_u8_u4_n181 ) , .B1( u2_u8_u4_n185 ) , .ZN( u2_u8_u4_n94 ) );
  INV_X1 u2_u8_u4_U39 (.A( u2_u8_u4_n113 ) , .ZN( u2_u8_u4_n185 ) );
  INV_X1 u2_u8_u4_U4 (.A( u2_u8_u4_n117 ) , .ZN( u2_u8_u4_n184 ) );
  INV_X1 u2_u8_u4_U40 (.A( u2_u8_u4_n143 ) , .ZN( u2_u8_u4_n183 ) );
  NOR2_X1 u2_u8_u4_U41 (.ZN( u2_u8_u4_n138 ) , .A1( u2_u8_u4_n168 ) , .A2( u2_u8_u4_n169 ) );
  NOR2_X1 u2_u8_u4_U42 (.A1( u2_u8_u4_n150 ) , .A2( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n153 ) );
  NOR2_X1 u2_u8_u4_U43 (.A2( u2_u8_u4_n128 ) , .A1( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n156 ) );
  AOI22_X1 u2_u8_u4_U44 (.B2( u2_u8_u4_n122 ) , .A1( u2_u8_u4_n123 ) , .ZN( u2_u8_u4_n124 ) , .B1( u2_u8_u4_n128 ) , .A2( u2_u8_u4_n172 ) );
  INV_X1 u2_u8_u4_U45 (.A( u2_u8_u4_n153 ) , .ZN( u2_u8_u4_n172 ) );
  NAND2_X1 u2_u8_u4_U46 (.A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n123 ) , .A1( u2_u8_u4_n161 ) );
  AOI22_X1 u2_u8_u4_U47 (.B2( u2_u8_u4_n132 ) , .A2( u2_u8_u4_n133 ) , .ZN( u2_u8_u4_n140 ) , .A1( u2_u8_u4_n150 ) , .B1( u2_u8_u4_n179 ) );
  NAND2_X1 u2_u8_u4_U48 (.ZN( u2_u8_u4_n133 ) , .A2( u2_u8_u4_n146 ) , .A1( u2_u8_u4_n154 ) );
  NAND2_X1 u2_u8_u4_U49 (.A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n154 ) , .A2( u2_u8_u4_n98 ) );
  NOR4_X1 u2_u8_u4_U5 (.A4( u2_u8_u4_n106 ) , .A3( u2_u8_u4_n107 ) , .A2( u2_u8_u4_n108 ) , .A1( u2_u8_u4_n109 ) , .ZN( u2_u8_u4_n110 ) );
  NAND2_X1 u2_u8_u4_U50 (.A1( u2_u8_u4_n101 ) , .ZN( u2_u8_u4_n158 ) , .A2( u2_u8_u4_n99 ) );
  AOI21_X1 u2_u8_u4_U51 (.ZN( u2_u8_u4_n127 ) , .A( u2_u8_u4_n136 ) , .B2( u2_u8_u4_n150 ) , .B1( u2_u8_u4_n180 ) );
  INV_X1 u2_u8_u4_U52 (.A( u2_u8_u4_n160 ) , .ZN( u2_u8_u4_n180 ) );
  NAND2_X1 u2_u8_u4_U53 (.A2( u2_u8_u4_n104 ) , .A1( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n146 ) );
  NAND2_X1 u2_u8_u4_U54 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n160 ) );
  NAND2_X1 u2_u8_u4_U55 (.ZN( u2_u8_u4_n134 ) , .A1( u2_u8_u4_n98 ) , .A2( u2_u8_u4_n99 ) );
  NAND2_X1 u2_u8_u4_U56 (.A1( u2_u8_u4_n103 ) , .A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n143 ) );
  NAND2_X1 u2_u8_u4_U57 (.A2( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n145 ) , .A1( u2_u8_u4_n98 ) );
  NAND2_X1 u2_u8_u4_U58 (.A1( u2_u8_u4_n100 ) , .A2( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n120 ) );
  NAND2_X1 u2_u8_u4_U59 (.A1( u2_u8_u4_n102 ) , .A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n148 ) );
  AOI21_X1 u2_u8_u4_U6 (.ZN( u2_u8_u4_n106 ) , .B2( u2_u8_u4_n146 ) , .B1( u2_u8_u4_n158 ) , .A( u2_u8_u4_n170 ) );
  NAND2_X1 u2_u8_u4_U60 (.A2( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n157 ) );
  INV_X1 u2_u8_u4_U61 (.A( u2_u8_u4_n150 ) , .ZN( u2_u8_u4_n173 ) );
  INV_X1 u2_u8_u4_U62 (.A( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n171 ) );
  NAND2_X1 u2_u8_u4_U63 (.A1( u2_u8_u4_n100 ) , .ZN( u2_u8_u4_n118 ) , .A2( u2_u8_u4_n99 ) );
  NAND2_X1 u2_u8_u4_U64 (.A2( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n144 ) );
  NAND2_X1 u2_u8_u4_U65 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n96 ) );
  INV_X1 u2_u8_u4_U66 (.A( u2_u8_u4_n128 ) , .ZN( u2_u8_u4_n174 ) );
  NAND2_X1 u2_u8_u4_U67 (.A2( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n119 ) , .A1( u2_u8_u4_n98 ) );
  NAND2_X1 u2_u8_u4_U68 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n147 ) );
  NAND2_X1 u2_u8_u4_U69 (.A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n113 ) , .A1( u2_u8_u4_n99 ) );
  AOI21_X1 u2_u8_u4_U7 (.ZN( u2_u8_u4_n108 ) , .B2( u2_u8_u4_n134 ) , .B1( u2_u8_u4_n155 ) , .A( u2_u8_u4_n156 ) );
  NOR2_X1 u2_u8_u4_U70 (.A2( u2_u8_X_28 ) , .ZN( u2_u8_u4_n150 ) , .A1( u2_u8_u4_n168 ) );
  NOR2_X1 u2_u8_u4_U71 (.A2( u2_u8_X_29 ) , .ZN( u2_u8_u4_n152 ) , .A1( u2_u8_u4_n169 ) );
  NOR2_X1 u2_u8_u4_U72 (.A2( u2_u8_X_30 ) , .ZN( u2_u8_u4_n105 ) , .A1( u2_u8_u4_n176 ) );
  NOR2_X1 u2_u8_u4_U73 (.A2( u2_u8_X_26 ) , .ZN( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n177 ) );
  NOR2_X1 u2_u8_u4_U74 (.A2( u2_u8_X_28 ) , .A1( u2_u8_X_29 ) , .ZN( u2_u8_u4_n128 ) );
  NOR2_X1 u2_u8_u4_U75 (.A2( u2_u8_X_27 ) , .A1( u2_u8_X_30 ) , .ZN( u2_u8_u4_n102 ) );
  NOR2_X1 u2_u8_u4_U76 (.A2( u2_u8_X_25 ) , .A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n98 ) );
  AND2_X1 u2_u8_u4_U77 (.A2( u2_u8_X_25 ) , .A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n104 ) );
  AND2_X1 u2_u8_u4_U78 (.A1( u2_u8_X_30 ) , .A2( u2_u8_u4_n176 ) , .ZN( u2_u8_u4_n99 ) );
  AND2_X1 u2_u8_u4_U79 (.A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n101 ) , .A2( u2_u8_u4_n177 ) );
  AOI21_X1 u2_u8_u4_U8 (.ZN( u2_u8_u4_n109 ) , .A( u2_u8_u4_n153 ) , .B1( u2_u8_u4_n159 ) , .B2( u2_u8_u4_n184 ) );
  AND2_X1 u2_u8_u4_U80 (.A1( u2_u8_X_27 ) , .A2( u2_u8_X_30 ) , .ZN( u2_u8_u4_n103 ) );
  INV_X1 u2_u8_u4_U81 (.A( u2_u8_X_28 ) , .ZN( u2_u8_u4_n169 ) );
  INV_X1 u2_u8_u4_U82 (.A( u2_u8_X_29 ) , .ZN( u2_u8_u4_n168 ) );
  INV_X1 u2_u8_u4_U83 (.A( u2_u8_X_25 ) , .ZN( u2_u8_u4_n177 ) );
  INV_X1 u2_u8_u4_U84 (.A( u2_u8_X_27 ) , .ZN( u2_u8_u4_n176 ) );
  NAND4_X1 u2_u8_u4_U85 (.ZN( u2_out8_25 ) , .A4( u2_u8_u4_n139 ) , .A3( u2_u8_u4_n140 ) , .A2( u2_u8_u4_n141 ) , .A1( u2_u8_u4_n142 ) );
  OAI21_X1 u2_u8_u4_U86 (.B2( u2_u8_u4_n131 ) , .ZN( u2_u8_u4_n141 ) , .A( u2_u8_u4_n175 ) , .B1( u2_u8_u4_n183 ) );
  OAI21_X1 u2_u8_u4_U87 (.A( u2_u8_u4_n128 ) , .B2( u2_u8_u4_n129 ) , .B1( u2_u8_u4_n130 ) , .ZN( u2_u8_u4_n142 ) );
  NAND4_X1 u2_u8_u4_U88 (.ZN( u2_out8_14 ) , .A4( u2_u8_u4_n124 ) , .A3( u2_u8_u4_n125 ) , .A2( u2_u8_u4_n126 ) , .A1( u2_u8_u4_n127 ) );
  AOI22_X1 u2_u8_u4_U89 (.B2( u2_u8_u4_n117 ) , .ZN( u2_u8_u4_n126 ) , .A1( u2_u8_u4_n129 ) , .B1( u2_u8_u4_n152 ) , .A2( u2_u8_u4_n175 ) );
  AOI211_X1 u2_u8_u4_U9 (.B( u2_u8_u4_n136 ) , .A( u2_u8_u4_n137 ) , .C2( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n139 ) , .C1( u2_u8_u4_n182 ) );
  AOI22_X1 u2_u8_u4_U90 (.ZN( u2_u8_u4_n125 ) , .B2( u2_u8_u4_n131 ) , .A2( u2_u8_u4_n132 ) , .B1( u2_u8_u4_n138 ) , .A1( u2_u8_u4_n178 ) );
  NAND4_X1 u2_u8_u4_U91 (.ZN( u2_out8_8 ) , .A4( u2_u8_u4_n110 ) , .A3( u2_u8_u4_n111 ) , .A2( u2_u8_u4_n112 ) , .A1( u2_u8_u4_n186 ) );
  NAND2_X1 u2_u8_u4_U92 (.ZN( u2_u8_u4_n112 ) , .A2( u2_u8_u4_n130 ) , .A1( u2_u8_u4_n150 ) );
  AOI22_X1 u2_u8_u4_U93 (.ZN( u2_u8_u4_n111 ) , .B2( u2_u8_u4_n132 ) , .A1( u2_u8_u4_n152 ) , .B1( u2_u8_u4_n178 ) , .A2( u2_u8_u4_n97 ) );
  AOI22_X1 u2_u8_u4_U94 (.B2( u2_u8_u4_n149 ) , .B1( u2_u8_u4_n150 ) , .A2( u2_u8_u4_n151 ) , .A1( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n167 ) );
  NOR4_X1 u2_u8_u4_U95 (.A4( u2_u8_u4_n162 ) , .A3( u2_u8_u4_n163 ) , .A2( u2_u8_u4_n164 ) , .A1( u2_u8_u4_n165 ) , .ZN( u2_u8_u4_n166 ) );
  NAND3_X1 u2_u8_u4_U96 (.ZN( u2_out8_3 ) , .A3( u2_u8_u4_n166 ) , .A1( u2_u8_u4_n167 ) , .A2( u2_u8_u4_n186 ) );
  NAND3_X1 u2_u8_u4_U97 (.A3( u2_u8_u4_n146 ) , .A2( u2_u8_u4_n147 ) , .A1( u2_u8_u4_n148 ) , .ZN( u2_u8_u4_n149 ) );
  NAND3_X1 u2_u8_u4_U98 (.A3( u2_u8_u4_n143 ) , .A2( u2_u8_u4_n144 ) , .A1( u2_u8_u4_n145 ) , .ZN( u2_u8_u4_n151 ) );
  NAND3_X1 u2_u8_u4_U99 (.A3( u2_u8_u4_n121 ) , .ZN( u2_u8_u4_n122 ) , .A2( u2_u8_u4_n144 ) , .A1( u2_u8_u4_n154 ) );
  AOI22_X1 u2_u8_u6_U10 (.A2( u2_u8_u6_n151 ) , .B2( u2_u8_u6_n161 ) , .A1( u2_u8_u6_n167 ) , .B1( u2_u8_u6_n170 ) , .ZN( u2_u8_u6_n89 ) );
  AOI21_X1 u2_u8_u6_U11 (.B1( u2_u8_u6_n107 ) , .B2( u2_u8_u6_n132 ) , .A( u2_u8_u6_n158 ) , .ZN( u2_u8_u6_n88 ) );
  AOI21_X1 u2_u8_u6_U12 (.B2( u2_u8_u6_n147 ) , .B1( u2_u8_u6_n148 ) , .ZN( u2_u8_u6_n149 ) , .A( u2_u8_u6_n158 ) );
  AOI21_X1 u2_u8_u6_U13 (.ZN( u2_u8_u6_n106 ) , .A( u2_u8_u6_n142 ) , .B2( u2_u8_u6_n159 ) , .B1( u2_u8_u6_n164 ) );
  INV_X1 u2_u8_u6_U14 (.A( u2_u8_u6_n155 ) , .ZN( u2_u8_u6_n161 ) );
  INV_X1 u2_u8_u6_U15 (.A( u2_u8_u6_n128 ) , .ZN( u2_u8_u6_n164 ) );
  NAND2_X1 u2_u8_u6_U16 (.ZN( u2_u8_u6_n110 ) , .A1( u2_u8_u6_n122 ) , .A2( u2_u8_u6_n129 ) );
  NAND2_X1 u2_u8_u6_U17 (.ZN( u2_u8_u6_n124 ) , .A2( u2_u8_u6_n146 ) , .A1( u2_u8_u6_n148 ) );
  INV_X1 u2_u8_u6_U18 (.A( u2_u8_u6_n132 ) , .ZN( u2_u8_u6_n171 ) );
  AND2_X1 u2_u8_u6_U19 (.A1( u2_u8_u6_n100 ) , .ZN( u2_u8_u6_n130 ) , .A2( u2_u8_u6_n147 ) );
  INV_X1 u2_u8_u6_U20 (.A( u2_u8_u6_n127 ) , .ZN( u2_u8_u6_n173 ) );
  INV_X1 u2_u8_u6_U21 (.A( u2_u8_u6_n121 ) , .ZN( u2_u8_u6_n167 ) );
  INV_X1 u2_u8_u6_U22 (.A( u2_u8_u6_n100 ) , .ZN( u2_u8_u6_n169 ) );
  INV_X1 u2_u8_u6_U23 (.A( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n170 ) );
  INV_X1 u2_u8_u6_U24 (.A( u2_u8_u6_n113 ) , .ZN( u2_u8_u6_n168 ) );
  AND2_X1 u2_u8_u6_U25 (.A1( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n119 ) , .ZN( u2_u8_u6_n133 ) );
  AND2_X1 u2_u8_u6_U26 (.A2( u2_u8_u6_n121 ) , .A1( u2_u8_u6_n122 ) , .ZN( u2_u8_u6_n131 ) );
  AND3_X1 u2_u8_u6_U27 (.ZN( u2_u8_u6_n120 ) , .A2( u2_u8_u6_n127 ) , .A1( u2_u8_u6_n132 ) , .A3( u2_u8_u6_n145 ) );
  INV_X1 u2_u8_u6_U28 (.A( u2_u8_u6_n146 ) , .ZN( u2_u8_u6_n163 ) );
  AOI222_X1 u2_u8_u6_U29 (.ZN( u2_u8_u6_n114 ) , .A1( u2_u8_u6_n118 ) , .A2( u2_u8_u6_n126 ) , .B2( u2_u8_u6_n151 ) , .C2( u2_u8_u6_n159 ) , .C1( u2_u8_u6_n168 ) , .B1( u2_u8_u6_n169 ) );
  INV_X1 u2_u8_u6_U3 (.A( u2_u8_u6_n110 ) , .ZN( u2_u8_u6_n166 ) );
  NOR2_X1 u2_u8_u6_U30 (.A1( u2_u8_u6_n162 ) , .A2( u2_u8_u6_n165 ) , .ZN( u2_u8_u6_n98 ) );
  AOI211_X1 u2_u8_u6_U31 (.B( u2_u8_u6_n134 ) , .A( u2_u8_u6_n135 ) , .C1( u2_u8_u6_n136 ) , .ZN( u2_u8_u6_n137 ) , .C2( u2_u8_u6_n151 ) );
  AOI21_X1 u2_u8_u6_U32 (.B2( u2_u8_u6_n132 ) , .B1( u2_u8_u6_n133 ) , .ZN( u2_u8_u6_n134 ) , .A( u2_u8_u6_n158 ) );
  NAND4_X1 u2_u8_u6_U33 (.A4( u2_u8_u6_n127 ) , .A3( u2_u8_u6_n128 ) , .A2( u2_u8_u6_n129 ) , .A1( u2_u8_u6_n130 ) , .ZN( u2_u8_u6_n136 ) );
  AOI21_X1 u2_u8_u6_U34 (.B1( u2_u8_u6_n131 ) , .ZN( u2_u8_u6_n135 ) , .A( u2_u8_u6_n144 ) , .B2( u2_u8_u6_n146 ) );
  NAND2_X1 u2_u8_u6_U35 (.A1( u2_u8_u6_n144 ) , .ZN( u2_u8_u6_n151 ) , .A2( u2_u8_u6_n158 ) );
  NAND2_X1 u2_u8_u6_U36 (.ZN( u2_u8_u6_n132 ) , .A1( u2_u8_u6_n91 ) , .A2( u2_u8_u6_n97 ) );
  AOI22_X1 u2_u8_u6_U37 (.B2( u2_u8_u6_n110 ) , .B1( u2_u8_u6_n111 ) , .A1( u2_u8_u6_n112 ) , .ZN( u2_u8_u6_n115 ) , .A2( u2_u8_u6_n161 ) );
  NAND4_X1 u2_u8_u6_U38 (.A3( u2_u8_u6_n109 ) , .ZN( u2_u8_u6_n112 ) , .A4( u2_u8_u6_n132 ) , .A2( u2_u8_u6_n147 ) , .A1( u2_u8_u6_n166 ) );
  NOR2_X1 u2_u8_u6_U39 (.ZN( u2_u8_u6_n109 ) , .A1( u2_u8_u6_n170 ) , .A2( u2_u8_u6_n173 ) );
  INV_X1 u2_u8_u6_U4 (.A( u2_u8_u6_n142 ) , .ZN( u2_u8_u6_n174 ) );
  NOR2_X1 u2_u8_u6_U40 (.A2( u2_u8_u6_n126 ) , .ZN( u2_u8_u6_n155 ) , .A1( u2_u8_u6_n160 ) );
  NAND2_X1 u2_u8_u6_U41 (.ZN( u2_u8_u6_n146 ) , .A2( u2_u8_u6_n94 ) , .A1( u2_u8_u6_n99 ) );
  AOI21_X1 u2_u8_u6_U42 (.A( u2_u8_u6_n144 ) , .B2( u2_u8_u6_n145 ) , .B1( u2_u8_u6_n146 ) , .ZN( u2_u8_u6_n150 ) );
  INV_X1 u2_u8_u6_U43 (.A( u2_u8_u6_n111 ) , .ZN( u2_u8_u6_n158 ) );
  NAND2_X1 u2_u8_u6_U44 (.ZN( u2_u8_u6_n127 ) , .A1( u2_u8_u6_n91 ) , .A2( u2_u8_u6_n92 ) );
  NAND2_X1 u2_u8_u6_U45 (.ZN( u2_u8_u6_n129 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n96 ) );
  INV_X1 u2_u8_u6_U46 (.A( u2_u8_u6_n144 ) , .ZN( u2_u8_u6_n159 ) );
  NAND2_X1 u2_u8_u6_U47 (.ZN( u2_u8_u6_n145 ) , .A2( u2_u8_u6_n97 ) , .A1( u2_u8_u6_n98 ) );
  NAND2_X1 u2_u8_u6_U48 (.ZN( u2_u8_u6_n148 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n94 ) );
  NAND2_X1 u2_u8_u6_U49 (.ZN( u2_u8_u6_n108 ) , .A2( u2_u8_u6_n139 ) , .A1( u2_u8_u6_n144 ) );
  NAND2_X1 u2_u8_u6_U5 (.A2( u2_u8_u6_n143 ) , .ZN( u2_u8_u6_n152 ) , .A1( u2_u8_u6_n166 ) );
  NAND2_X1 u2_u8_u6_U50 (.ZN( u2_u8_u6_n121 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n97 ) );
  NAND2_X1 u2_u8_u6_U51 (.ZN( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n95 ) );
  AND2_X1 u2_u8_u6_U52 (.ZN( u2_u8_u6_n118 ) , .A2( u2_u8_u6_n91 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U53 (.ZN( u2_u8_u6_n147 ) , .A2( u2_u8_u6_n98 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U54 (.ZN( u2_u8_u6_n128 ) , .A1( u2_u8_u6_n94 ) , .A2( u2_u8_u6_n96 ) );
  NAND2_X1 u2_u8_u6_U55 (.ZN( u2_u8_u6_n119 ) , .A2( u2_u8_u6_n95 ) , .A1( u2_u8_u6_n99 ) );
  NAND2_X1 u2_u8_u6_U56 (.ZN( u2_u8_u6_n123 ) , .A2( u2_u8_u6_n91 ) , .A1( u2_u8_u6_n96 ) );
  NAND2_X1 u2_u8_u6_U57 (.ZN( u2_u8_u6_n100 ) , .A2( u2_u8_u6_n92 ) , .A1( u2_u8_u6_n98 ) );
  NAND2_X1 u2_u8_u6_U58 (.ZN( u2_u8_u6_n122 ) , .A1( u2_u8_u6_n94 ) , .A2( u2_u8_u6_n97 ) );
  INV_X1 u2_u8_u6_U59 (.A( u2_u8_u6_n139 ) , .ZN( u2_u8_u6_n160 ) );
  AOI22_X1 u2_u8_u6_U6 (.B2( u2_u8_u6_n101 ) , .A1( u2_u8_u6_n102 ) , .ZN( u2_u8_u6_n103 ) , .B1( u2_u8_u6_n160 ) , .A2( u2_u8_u6_n161 ) );
  NAND2_X1 u2_u8_u6_U60 (.ZN( u2_u8_u6_n113 ) , .A1( u2_u8_u6_n96 ) , .A2( u2_u8_u6_n98 ) );
  NOR2_X1 u2_u8_u6_U61 (.A2( u2_u8_X_40 ) , .A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n126 ) );
  NOR2_X1 u2_u8_u6_U62 (.A2( u2_u8_X_39 ) , .A1( u2_u8_X_42 ) , .ZN( u2_u8_u6_n92 ) );
  NOR2_X1 u2_u8_u6_U63 (.A2( u2_u8_X_39 ) , .A1( u2_u8_u6_n156 ) , .ZN( u2_u8_u6_n97 ) );
  NOR2_X1 u2_u8_u6_U64 (.A2( u2_u8_X_38 ) , .A1( u2_u8_u6_n165 ) , .ZN( u2_u8_u6_n95 ) );
  NOR2_X1 u2_u8_u6_U65 (.A2( u2_u8_X_41 ) , .ZN( u2_u8_u6_n111 ) , .A1( u2_u8_u6_n157 ) );
  NOR2_X1 u2_u8_u6_U66 (.A2( u2_u8_X_37 ) , .A1( u2_u8_u6_n162 ) , .ZN( u2_u8_u6_n94 ) );
  NOR2_X1 u2_u8_u6_U67 (.A2( u2_u8_X_37 ) , .A1( u2_u8_X_38 ) , .ZN( u2_u8_u6_n91 ) );
  NAND2_X1 u2_u8_u6_U68 (.A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n144 ) , .A2( u2_u8_u6_n157 ) );
  NAND2_X1 u2_u8_u6_U69 (.A2( u2_u8_X_40 ) , .A1( u2_u8_X_41 ) , .ZN( u2_u8_u6_n139 ) );
  NOR2_X1 u2_u8_u6_U7 (.A1( u2_u8_u6_n118 ) , .ZN( u2_u8_u6_n143 ) , .A2( u2_u8_u6_n168 ) );
  AND2_X1 u2_u8_u6_U70 (.A1( u2_u8_X_39 ) , .A2( u2_u8_u6_n156 ) , .ZN( u2_u8_u6_n96 ) );
  AND2_X1 u2_u8_u6_U71 (.A1( u2_u8_X_39 ) , .A2( u2_u8_X_42 ) , .ZN( u2_u8_u6_n99 ) );
  INV_X1 u2_u8_u6_U72 (.A( u2_u8_X_40 ) , .ZN( u2_u8_u6_n157 ) );
  INV_X1 u2_u8_u6_U73 (.A( u2_u8_X_37 ) , .ZN( u2_u8_u6_n165 ) );
  INV_X1 u2_u8_u6_U74 (.A( u2_u8_X_38 ) , .ZN( u2_u8_u6_n162 ) );
  INV_X1 u2_u8_u6_U75 (.A( u2_u8_X_42 ) , .ZN( u2_u8_u6_n156 ) );
  NAND4_X1 u2_u8_u6_U76 (.ZN( u2_out8_32 ) , .A4( u2_u8_u6_n103 ) , .A3( u2_u8_u6_n104 ) , .A2( u2_u8_u6_n105 ) , .A1( u2_u8_u6_n106 ) );
  AOI22_X1 u2_u8_u6_U77 (.ZN( u2_u8_u6_n105 ) , .A2( u2_u8_u6_n108 ) , .A1( u2_u8_u6_n118 ) , .B2( u2_u8_u6_n126 ) , .B1( u2_u8_u6_n171 ) );
  AOI22_X1 u2_u8_u6_U78 (.ZN( u2_u8_u6_n104 ) , .A1( u2_u8_u6_n111 ) , .B1( u2_u8_u6_n124 ) , .B2( u2_u8_u6_n151 ) , .A2( u2_u8_u6_n93 ) );
  NAND4_X1 u2_u8_u6_U79 (.ZN( u2_out8_12 ) , .A4( u2_u8_u6_n114 ) , .A3( u2_u8_u6_n115 ) , .A2( u2_u8_u6_n116 ) , .A1( u2_u8_u6_n117 ) );
  OAI21_X1 u2_u8_u6_U8 (.A( u2_u8_u6_n159 ) , .B1( u2_u8_u6_n169 ) , .B2( u2_u8_u6_n173 ) , .ZN( u2_u8_u6_n90 ) );
  OAI22_X1 u2_u8_u6_U80 (.B2( u2_u8_u6_n111 ) , .ZN( u2_u8_u6_n116 ) , .B1( u2_u8_u6_n126 ) , .A2( u2_u8_u6_n164 ) , .A1( u2_u8_u6_n167 ) );
  OAI21_X1 u2_u8_u6_U81 (.A( u2_u8_u6_n108 ) , .ZN( u2_u8_u6_n117 ) , .B2( u2_u8_u6_n141 ) , .B1( u2_u8_u6_n163 ) );
  OAI211_X1 u2_u8_u6_U82 (.ZN( u2_out8_7 ) , .B( u2_u8_u6_n153 ) , .C2( u2_u8_u6_n154 ) , .C1( u2_u8_u6_n155 ) , .A( u2_u8_u6_n174 ) );
  NOR3_X1 u2_u8_u6_U83 (.A1( u2_u8_u6_n141 ) , .ZN( u2_u8_u6_n154 ) , .A3( u2_u8_u6_n164 ) , .A2( u2_u8_u6_n171 ) );
  AOI211_X1 u2_u8_u6_U84 (.B( u2_u8_u6_n149 ) , .A( u2_u8_u6_n150 ) , .C2( u2_u8_u6_n151 ) , .C1( u2_u8_u6_n152 ) , .ZN( u2_u8_u6_n153 ) );
  OAI211_X1 u2_u8_u6_U85 (.ZN( u2_out8_22 ) , .B( u2_u8_u6_n137 ) , .A( u2_u8_u6_n138 ) , .C2( u2_u8_u6_n139 ) , .C1( u2_u8_u6_n140 ) );
  AOI22_X1 u2_u8_u6_U86 (.B1( u2_u8_u6_n124 ) , .A2( u2_u8_u6_n125 ) , .A1( u2_u8_u6_n126 ) , .ZN( u2_u8_u6_n138 ) , .B2( u2_u8_u6_n161 ) );
  AND4_X1 u2_u8_u6_U87 (.A3( u2_u8_u6_n119 ) , .A1( u2_u8_u6_n120 ) , .A4( u2_u8_u6_n129 ) , .ZN( u2_u8_u6_n140 ) , .A2( u2_u8_u6_n143 ) );
  NAND3_X1 u2_u8_u6_U88 (.A2( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n125 ) , .A1( u2_u8_u6_n130 ) , .A3( u2_u8_u6_n131 ) );
  NAND3_X1 u2_u8_u6_U89 (.A3( u2_u8_u6_n133 ) , .ZN( u2_u8_u6_n141 ) , .A1( u2_u8_u6_n145 ) , .A2( u2_u8_u6_n148 ) );
  INV_X1 u2_u8_u6_U9 (.ZN( u2_u8_u6_n172 ) , .A( u2_u8_u6_n88 ) );
  NAND3_X1 u2_u8_u6_U90 (.ZN( u2_u8_u6_n101 ) , .A3( u2_u8_u6_n107 ) , .A2( u2_u8_u6_n121 ) , .A1( u2_u8_u6_n127 ) );
  NAND3_X1 u2_u8_u6_U91 (.ZN( u2_u8_u6_n102 ) , .A3( u2_u8_u6_n130 ) , .A2( u2_u8_u6_n145 ) , .A1( u2_u8_u6_n166 ) );
  NAND3_X1 u2_u8_u6_U92 (.A3( u2_u8_u6_n113 ) , .A1( u2_u8_u6_n119 ) , .A2( u2_u8_u6_n123 ) , .ZN( u2_u8_u6_n93 ) );
  NAND3_X1 u2_u8_u6_U93 (.ZN( u2_u8_u6_n142 ) , .A2( u2_u8_u6_n172 ) , .A3( u2_u8_u6_n89 ) , .A1( u2_u8_u6_n90 ) );
  AND3_X1 u2_u8_u7_U10 (.A3( u2_u8_u7_n110 ) , .A2( u2_u8_u7_n127 ) , .A1( u2_u8_u7_n132 ) , .ZN( u2_u8_u7_n92 ) );
  OAI21_X1 u2_u8_u7_U11 (.A( u2_u8_u7_n161 ) , .B1( u2_u8_u7_n168 ) , .B2( u2_u8_u7_n173 ) , .ZN( u2_u8_u7_n91 ) );
  AOI211_X1 u2_u8_u7_U12 (.A( u2_u8_u7_n117 ) , .ZN( u2_u8_u7_n118 ) , .C2( u2_u8_u7_n126 ) , .C1( u2_u8_u7_n177 ) , .B( u2_u8_u7_n180 ) );
  OAI22_X1 u2_u8_u7_U13 (.B1( u2_u8_u7_n115 ) , .ZN( u2_u8_u7_n117 ) , .A2( u2_u8_u7_n133 ) , .A1( u2_u8_u7_n137 ) , .B2( u2_u8_u7_n162 ) );
  INV_X1 u2_u8_u7_U14 (.A( u2_u8_u7_n116 ) , .ZN( u2_u8_u7_n180 ) );
  NOR3_X1 u2_u8_u7_U15 (.ZN( u2_u8_u7_n115 ) , .A3( u2_u8_u7_n145 ) , .A2( u2_u8_u7_n168 ) , .A1( u2_u8_u7_n169 ) );
  OAI211_X1 u2_u8_u7_U16 (.B( u2_u8_u7_n122 ) , .A( u2_u8_u7_n123 ) , .C2( u2_u8_u7_n124 ) , .ZN( u2_u8_u7_n154 ) , .C1( u2_u8_u7_n162 ) );
  AOI222_X1 u2_u8_u7_U17 (.ZN( u2_u8_u7_n122 ) , .C2( u2_u8_u7_n126 ) , .C1( u2_u8_u7_n145 ) , .B1( u2_u8_u7_n161 ) , .A2( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n170 ) , .A1( u2_u8_u7_n176 ) );
  INV_X1 u2_u8_u7_U18 (.A( u2_u8_u7_n133 ) , .ZN( u2_u8_u7_n176 ) );
  NOR3_X1 u2_u8_u7_U19 (.A2( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n135 ) , .ZN( u2_u8_u7_n136 ) , .A3( u2_u8_u7_n171 ) );
  NOR2_X1 u2_u8_u7_U20 (.A1( u2_u8_u7_n130 ) , .A2( u2_u8_u7_n134 ) , .ZN( u2_u8_u7_n153 ) );
  INV_X1 u2_u8_u7_U21 (.A( u2_u8_u7_n101 ) , .ZN( u2_u8_u7_n165 ) );
  NOR2_X1 u2_u8_u7_U22 (.ZN( u2_u8_u7_n111 ) , .A2( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n169 ) );
  AOI21_X1 u2_u8_u7_U23 (.ZN( u2_u8_u7_n104 ) , .B2( u2_u8_u7_n112 ) , .B1( u2_u8_u7_n127 ) , .A( u2_u8_u7_n164 ) );
  AOI21_X1 u2_u8_u7_U24 (.ZN( u2_u8_u7_n106 ) , .B1( u2_u8_u7_n133 ) , .B2( u2_u8_u7_n146 ) , .A( u2_u8_u7_n162 ) );
  AOI21_X1 u2_u8_u7_U25 (.A( u2_u8_u7_n101 ) , .ZN( u2_u8_u7_n107 ) , .B2( u2_u8_u7_n128 ) , .B1( u2_u8_u7_n175 ) );
  INV_X1 u2_u8_u7_U26 (.A( u2_u8_u7_n138 ) , .ZN( u2_u8_u7_n171 ) );
  INV_X1 u2_u8_u7_U27 (.A( u2_u8_u7_n131 ) , .ZN( u2_u8_u7_n177 ) );
  INV_X1 u2_u8_u7_U28 (.A( u2_u8_u7_n110 ) , .ZN( u2_u8_u7_n174 ) );
  NAND2_X1 u2_u8_u7_U29 (.A1( u2_u8_u7_n129 ) , .A2( u2_u8_u7_n132 ) , .ZN( u2_u8_u7_n149 ) );
  OAI21_X1 u2_u8_u7_U3 (.ZN( u2_u8_u7_n159 ) , .A( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n171 ) , .B1( u2_u8_u7_n174 ) );
  NAND2_X1 u2_u8_u7_U30 (.A1( u2_u8_u7_n113 ) , .A2( u2_u8_u7_n124 ) , .ZN( u2_u8_u7_n130 ) );
  INV_X1 u2_u8_u7_U31 (.A( u2_u8_u7_n112 ) , .ZN( u2_u8_u7_n173 ) );
  INV_X1 u2_u8_u7_U32 (.A( u2_u8_u7_n128 ) , .ZN( u2_u8_u7_n168 ) );
  INV_X1 u2_u8_u7_U33 (.A( u2_u8_u7_n148 ) , .ZN( u2_u8_u7_n169 ) );
  INV_X1 u2_u8_u7_U34 (.A( u2_u8_u7_n127 ) , .ZN( u2_u8_u7_n179 ) );
  NOR2_X1 u2_u8_u7_U35 (.ZN( u2_u8_u7_n101 ) , .A2( u2_u8_u7_n150 ) , .A1( u2_u8_u7_n156 ) );
  AOI211_X1 u2_u8_u7_U36 (.B( u2_u8_u7_n154 ) , .A( u2_u8_u7_n155 ) , .C1( u2_u8_u7_n156 ) , .ZN( u2_u8_u7_n157 ) , .C2( u2_u8_u7_n172 ) );
  INV_X1 u2_u8_u7_U37 (.A( u2_u8_u7_n153 ) , .ZN( u2_u8_u7_n172 ) );
  AOI211_X1 u2_u8_u7_U38 (.B( u2_u8_u7_n139 ) , .A( u2_u8_u7_n140 ) , .C2( u2_u8_u7_n141 ) , .ZN( u2_u8_u7_n142 ) , .C1( u2_u8_u7_n156 ) );
  NAND4_X1 u2_u8_u7_U39 (.A3( u2_u8_u7_n127 ) , .A2( u2_u8_u7_n128 ) , .A1( u2_u8_u7_n129 ) , .ZN( u2_u8_u7_n141 ) , .A4( u2_u8_u7_n147 ) );
  INV_X1 u2_u8_u7_U4 (.A( u2_u8_u7_n111 ) , .ZN( u2_u8_u7_n170 ) );
  AOI21_X1 u2_u8_u7_U40 (.A( u2_u8_u7_n137 ) , .B1( u2_u8_u7_n138 ) , .ZN( u2_u8_u7_n139 ) , .B2( u2_u8_u7_n146 ) );
  OAI22_X1 u2_u8_u7_U41 (.B1( u2_u8_u7_n136 ) , .ZN( u2_u8_u7_n140 ) , .A1( u2_u8_u7_n153 ) , .B2( u2_u8_u7_n162 ) , .A2( u2_u8_u7_n164 ) );
  AOI21_X1 u2_u8_u7_U42 (.ZN( u2_u8_u7_n123 ) , .B1( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n177 ) , .A( u2_u8_u7_n97 ) );
  AOI21_X1 u2_u8_u7_U43 (.B2( u2_u8_u7_n113 ) , .B1( u2_u8_u7_n124 ) , .A( u2_u8_u7_n125 ) , .ZN( u2_u8_u7_n97 ) );
  INV_X1 u2_u8_u7_U44 (.A( u2_u8_u7_n125 ) , .ZN( u2_u8_u7_n161 ) );
  INV_X1 u2_u8_u7_U45 (.A( u2_u8_u7_n152 ) , .ZN( u2_u8_u7_n162 ) );
  AOI22_X1 u2_u8_u7_U46 (.A2( u2_u8_u7_n114 ) , .ZN( u2_u8_u7_n119 ) , .B1( u2_u8_u7_n130 ) , .A1( u2_u8_u7_n156 ) , .B2( u2_u8_u7_n165 ) );
  NAND2_X1 u2_u8_u7_U47 (.A2( u2_u8_u7_n112 ) , .ZN( u2_u8_u7_n114 ) , .A1( u2_u8_u7_n175 ) );
  AND2_X1 u2_u8_u7_U48 (.ZN( u2_u8_u7_n145 ) , .A2( u2_u8_u7_n98 ) , .A1( u2_u8_u7_n99 ) );
  NOR2_X1 u2_u8_u7_U49 (.ZN( u2_u8_u7_n137 ) , .A1( u2_u8_u7_n150 ) , .A2( u2_u8_u7_n161 ) );
  INV_X1 u2_u8_u7_U5 (.A( u2_u8_u7_n149 ) , .ZN( u2_u8_u7_n175 ) );
  AOI21_X1 u2_u8_u7_U50 (.ZN( u2_u8_u7_n105 ) , .B2( u2_u8_u7_n110 ) , .A( u2_u8_u7_n125 ) , .B1( u2_u8_u7_n147 ) );
  NAND2_X1 u2_u8_u7_U51 (.ZN( u2_u8_u7_n146 ) , .A1( u2_u8_u7_n95 ) , .A2( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U52 (.A2( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n147 ) , .A1( u2_u8_u7_n93 ) );
  NAND2_X1 u2_u8_u7_U53 (.A1( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n127 ) , .A2( u2_u8_u7_n99 ) );
  OR2_X1 u2_u8_u7_U54 (.ZN( u2_u8_u7_n126 ) , .A2( u2_u8_u7_n152 ) , .A1( u2_u8_u7_n156 ) );
  NAND2_X1 u2_u8_u7_U55 (.A2( u2_u8_u7_n102 ) , .A1( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n133 ) );
  NAND2_X1 u2_u8_u7_U56 (.ZN( u2_u8_u7_n112 ) , .A2( u2_u8_u7_n96 ) , .A1( u2_u8_u7_n99 ) );
  NAND2_X1 u2_u8_u7_U57 (.A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n128 ) , .A1( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U58 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n113 ) , .A2( u2_u8_u7_n93 ) );
  NAND2_X1 u2_u8_u7_U59 (.A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n124 ) , .A1( u2_u8_u7_n96 ) );
  INV_X1 u2_u8_u7_U6 (.A( u2_u8_u7_n154 ) , .ZN( u2_u8_u7_n178 ) );
  NAND2_X1 u2_u8_u7_U60 (.ZN( u2_u8_u7_n110 ) , .A1( u2_u8_u7_n95 ) , .A2( u2_u8_u7_n96 ) );
  INV_X1 u2_u8_u7_U61 (.A( u2_u8_u7_n150 ) , .ZN( u2_u8_u7_n164 ) );
  AND2_X1 u2_u8_u7_U62 (.ZN( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n93 ) , .A2( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U63 (.A1( u2_u8_u7_n100 ) , .A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n129 ) );
  NAND2_X1 u2_u8_u7_U64 (.A2( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n131 ) , .A1( u2_u8_u7_n95 ) );
  NAND2_X1 u2_u8_u7_U65 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n138 ) , .A2( u2_u8_u7_n99 ) );
  NAND2_X1 u2_u8_u7_U66 (.ZN( u2_u8_u7_n132 ) , .A1( u2_u8_u7_n93 ) , .A2( u2_u8_u7_n96 ) );
  NAND2_X1 u2_u8_u7_U67 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n148 ) , .A2( u2_u8_u7_n95 ) );
  NOR2_X1 u2_u8_u7_U68 (.A2( u2_u8_X_47 ) , .ZN( u2_u8_u7_n150 ) , .A1( u2_u8_u7_n163 ) );
  NOR2_X1 u2_u8_u7_U69 (.A2( u2_u8_X_43 ) , .A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n103 ) );
  AOI211_X1 u2_u8_u7_U7 (.ZN( u2_u8_u7_n116 ) , .A( u2_u8_u7_n155 ) , .C1( u2_u8_u7_n161 ) , .C2( u2_u8_u7_n171 ) , .B( u2_u8_u7_n94 ) );
  NOR2_X1 u2_u8_u7_U70 (.A2( u2_u8_X_48 ) , .A1( u2_u8_u7_n166 ) , .ZN( u2_u8_u7_n95 ) );
  NOR2_X1 u2_u8_u7_U71 (.A2( u2_u8_X_45 ) , .A1( u2_u8_X_48 ) , .ZN( u2_u8_u7_n99 ) );
  NOR2_X1 u2_u8_u7_U72 (.A2( u2_u8_X_44 ) , .A1( u2_u8_u7_n167 ) , .ZN( u2_u8_u7_n98 ) );
  NOR2_X1 u2_u8_u7_U73 (.A2( u2_u8_X_46 ) , .A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n152 ) );
  AND2_X1 u2_u8_u7_U74 (.A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n156 ) , .A2( u2_u8_u7_n163 ) );
  NAND2_X1 u2_u8_u7_U75 (.A2( u2_u8_X_46 ) , .A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n125 ) );
  AND2_X1 u2_u8_u7_U76 (.A2( u2_u8_X_45 ) , .A1( u2_u8_X_48 ) , .ZN( u2_u8_u7_n102 ) );
  AND2_X1 u2_u8_u7_U77 (.A2( u2_u8_X_43 ) , .A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n96 ) );
  AND2_X1 u2_u8_u7_U78 (.A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n100 ) , .A2( u2_u8_u7_n167 ) );
  AND2_X1 u2_u8_u7_U79 (.A1( u2_u8_X_48 ) , .A2( u2_u8_u7_n166 ) , .ZN( u2_u8_u7_n93 ) );
  OAI222_X1 u2_u8_u7_U8 (.C2( u2_u8_u7_n101 ) , .B2( u2_u8_u7_n111 ) , .A1( u2_u8_u7_n113 ) , .C1( u2_u8_u7_n146 ) , .A2( u2_u8_u7_n162 ) , .B1( u2_u8_u7_n164 ) , .ZN( u2_u8_u7_n94 ) );
  INV_X1 u2_u8_u7_U80 (.A( u2_u8_X_46 ) , .ZN( u2_u8_u7_n163 ) );
  INV_X1 u2_u8_u7_U81 (.A( u2_u8_X_43 ) , .ZN( u2_u8_u7_n167 ) );
  INV_X1 u2_u8_u7_U82 (.A( u2_u8_X_45 ) , .ZN( u2_u8_u7_n166 ) );
  NAND4_X1 u2_u8_u7_U83 (.ZN( u2_out8_27 ) , .A4( u2_u8_u7_n118 ) , .A3( u2_u8_u7_n119 ) , .A2( u2_u8_u7_n120 ) , .A1( u2_u8_u7_n121 ) );
  OAI21_X1 u2_u8_u7_U84 (.ZN( u2_u8_u7_n121 ) , .B2( u2_u8_u7_n145 ) , .A( u2_u8_u7_n150 ) , .B1( u2_u8_u7_n174 ) );
  OAI21_X1 u2_u8_u7_U85 (.ZN( u2_u8_u7_n120 ) , .A( u2_u8_u7_n161 ) , .B2( u2_u8_u7_n170 ) , .B1( u2_u8_u7_n179 ) );
  NAND4_X1 u2_u8_u7_U86 (.ZN( u2_out8_21 ) , .A4( u2_u8_u7_n157 ) , .A3( u2_u8_u7_n158 ) , .A2( u2_u8_u7_n159 ) , .A1( u2_u8_u7_n160 ) );
  OAI21_X1 u2_u8_u7_U87 (.B1( u2_u8_u7_n145 ) , .ZN( u2_u8_u7_n160 ) , .A( u2_u8_u7_n161 ) , .B2( u2_u8_u7_n177 ) );
  AOI22_X1 u2_u8_u7_U88 (.B2( u2_u8_u7_n149 ) , .B1( u2_u8_u7_n150 ) , .A2( u2_u8_u7_n151 ) , .A1( u2_u8_u7_n152 ) , .ZN( u2_u8_u7_n158 ) );
  NAND4_X1 u2_u8_u7_U89 (.ZN( u2_out8_15 ) , .A4( u2_u8_u7_n142 ) , .A3( u2_u8_u7_n143 ) , .A2( u2_u8_u7_n144 ) , .A1( u2_u8_u7_n178 ) );
  OAI221_X1 u2_u8_u7_U9 (.C1( u2_u8_u7_n101 ) , .C2( u2_u8_u7_n147 ) , .ZN( u2_u8_u7_n155 ) , .B2( u2_u8_u7_n162 ) , .A( u2_u8_u7_n91 ) , .B1( u2_u8_u7_n92 ) );
  OR2_X1 u2_u8_u7_U90 (.A2( u2_u8_u7_n125 ) , .A1( u2_u8_u7_n129 ) , .ZN( u2_u8_u7_n144 ) );
  AOI22_X1 u2_u8_u7_U91 (.A2( u2_u8_u7_n126 ) , .ZN( u2_u8_u7_n143 ) , .B2( u2_u8_u7_n165 ) , .B1( u2_u8_u7_n173 ) , .A1( u2_u8_u7_n174 ) );
  NAND4_X1 u2_u8_u7_U92 (.ZN( u2_out8_5 ) , .A4( u2_u8_u7_n108 ) , .A3( u2_u8_u7_n109 ) , .A1( u2_u8_u7_n116 ) , .A2( u2_u8_u7_n123 ) );
  AOI22_X1 u2_u8_u7_U93 (.ZN( u2_u8_u7_n109 ) , .A2( u2_u8_u7_n126 ) , .B2( u2_u8_u7_n145 ) , .B1( u2_u8_u7_n156 ) , .A1( u2_u8_u7_n171 ) );
  NOR4_X1 u2_u8_u7_U94 (.A4( u2_u8_u7_n104 ) , .A3( u2_u8_u7_n105 ) , .A2( u2_u8_u7_n106 ) , .A1( u2_u8_u7_n107 ) , .ZN( u2_u8_u7_n108 ) );
  NAND3_X1 u2_u8_u7_U95 (.A3( u2_u8_u7_n146 ) , .A2( u2_u8_u7_n147 ) , .A1( u2_u8_u7_n148 ) , .ZN( u2_u8_u7_n151 ) );
  NAND3_X1 u2_u8_u7_U96 (.A3( u2_u8_u7_n131 ) , .A2( u2_u8_u7_n132 ) , .A1( u2_u8_u7_n133 ) , .ZN( u2_u8_u7_n135 ) );
  XOR2_X1 u2_u9_U13 (.B( u2_K10_42 ) , .A( u2_R8_29 ) , .Z( u2_u9_X_42 ) );
  XOR2_X1 u2_u9_U14 (.B( u2_K10_41 ) , .A( u2_R8_28 ) , .Z( u2_u9_X_41 ) );
  XOR2_X1 u2_u9_U15 (.B( u2_K10_40 ) , .A( u2_R8_27 ) , .Z( u2_u9_X_40 ) );
  XOR2_X1 u2_u9_U17 (.B( u2_K10_39 ) , .A( u2_R8_26 ) , .Z( u2_u9_X_39 ) );
  XOR2_X1 u2_u9_U18 (.B( u2_K10_38 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_38 ) );
  XOR2_X1 u2_u9_U19 (.B( u2_K10_37 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_37 ) );
  XOR2_X1 u2_u9_U20 (.B( u2_K10_36 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_36 ) );
  XOR2_X1 u2_u9_U21 (.B( u2_K10_35 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_35 ) );
  XOR2_X1 u2_u9_U22 (.B( u2_K10_34 ) , .A( u2_R8_23 ) , .Z( u2_u9_X_34 ) );
  XOR2_X1 u2_u9_U23 (.B( u2_K10_33 ) , .A( u2_R8_22 ) , .Z( u2_u9_X_33 ) );
  XOR2_X1 u2_u9_U24 (.B( u2_K10_32 ) , .A( u2_R8_21 ) , .Z( u2_u9_X_32 ) );
  XOR2_X1 u2_u9_U25 (.B( u2_K10_31 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_31 ) );
  XOR2_X1 u2_u9_U26 (.B( u2_K10_30 ) , .A( u2_R8_21 ) , .Z( u2_u9_X_30 ) );
  XOR2_X1 u2_u9_U28 (.B( u2_K10_29 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_29 ) );
  XOR2_X1 u2_u9_U29 (.B( u2_K10_28 ) , .A( u2_R8_19 ) , .Z( u2_u9_X_28 ) );
  XOR2_X1 u2_u9_U30 (.B( u2_K10_27 ) , .A( u2_R8_18 ) , .Z( u2_u9_X_27 ) );
  XOR2_X1 u2_u9_U31 (.B( u2_K10_26 ) , .A( u2_R8_17 ) , .Z( u2_u9_X_26 ) );
  XOR2_X1 u2_u9_U32 (.B( u2_K10_25 ) , .A( u2_R8_16 ) , .Z( u2_u9_X_25 ) );
  XOR2_X1 u2_u9_U33 (.B( u2_K10_24 ) , .A( u2_R8_17 ) , .Z( u2_u9_X_24 ) );
  XOR2_X1 u2_u9_U34 (.B( u2_K10_23 ) , .A( u2_R8_16 ) , .Z( u2_u9_X_23 ) );
  XOR2_X1 u2_u9_U35 (.B( u2_K10_22 ) , .A( u2_R8_15 ) , .Z( u2_u9_X_22 ) );
  XOR2_X1 u2_u9_U36 (.B( u2_K10_21 ) , .A( u2_R8_14 ) , .Z( u2_u9_X_21 ) );
  XOR2_X1 u2_u9_U37 (.B( u2_K10_20 ) , .A( u2_R8_13 ) , .Z( u2_u9_X_20 ) );
  XOR2_X1 u2_u9_U39 (.B( u2_K10_19 ) , .A( u2_R8_12 ) , .Z( u2_u9_X_19 ) );
  OAI22_X1 u2_u9_u3_U10 (.B1( u2_u9_u3_n113 ) , .A2( u2_u9_u3_n135 ) , .A1( u2_u9_u3_n150 ) , .B2( u2_u9_u3_n164 ) , .ZN( u2_u9_u3_n98 ) );
  OAI211_X1 u2_u9_u3_U11 (.B( u2_u9_u3_n106 ) , .ZN( u2_u9_u3_n119 ) , .C2( u2_u9_u3_n128 ) , .C1( u2_u9_u3_n167 ) , .A( u2_u9_u3_n181 ) );
  AOI221_X1 u2_u9_u3_U12 (.C1( u2_u9_u3_n105 ) , .ZN( u2_u9_u3_n106 ) , .A( u2_u9_u3_n131 ) , .B2( u2_u9_u3_n132 ) , .C2( u2_u9_u3_n133 ) , .B1( u2_u9_u3_n169 ) );
  INV_X1 u2_u9_u3_U13 (.ZN( u2_u9_u3_n181 ) , .A( u2_u9_u3_n98 ) );
  NAND2_X1 u2_u9_u3_U14 (.ZN( u2_u9_u3_n105 ) , .A2( u2_u9_u3_n130 ) , .A1( u2_u9_u3_n155 ) );
  AOI22_X1 u2_u9_u3_U15 (.B1( u2_u9_u3_n115 ) , .A2( u2_u9_u3_n116 ) , .ZN( u2_u9_u3_n123 ) , .B2( u2_u9_u3_n133 ) , .A1( u2_u9_u3_n169 ) );
  NAND2_X1 u2_u9_u3_U16 (.ZN( u2_u9_u3_n116 ) , .A2( u2_u9_u3_n151 ) , .A1( u2_u9_u3_n182 ) );
  NOR2_X1 u2_u9_u3_U17 (.ZN( u2_u9_u3_n126 ) , .A2( u2_u9_u3_n150 ) , .A1( u2_u9_u3_n164 ) );
  AOI21_X1 u2_u9_u3_U18 (.ZN( u2_u9_u3_n112 ) , .B2( u2_u9_u3_n146 ) , .B1( u2_u9_u3_n155 ) , .A( u2_u9_u3_n167 ) );
  NAND2_X1 u2_u9_u3_U19 (.A1( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n142 ) , .A2( u2_u9_u3_n164 ) );
  NAND2_X1 u2_u9_u3_U20 (.ZN( u2_u9_u3_n132 ) , .A2( u2_u9_u3_n152 ) , .A1( u2_u9_u3_n156 ) );
  AND2_X1 u2_u9_u3_U21 (.A2( u2_u9_u3_n113 ) , .A1( u2_u9_u3_n114 ) , .ZN( u2_u9_u3_n151 ) );
  INV_X1 u2_u9_u3_U22 (.A( u2_u9_u3_n133 ) , .ZN( u2_u9_u3_n165 ) );
  INV_X1 u2_u9_u3_U23 (.A( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n170 ) );
  NAND2_X1 u2_u9_u3_U24 (.A1( u2_u9_u3_n107 ) , .A2( u2_u9_u3_n108 ) , .ZN( u2_u9_u3_n140 ) );
  NAND2_X1 u2_u9_u3_U25 (.ZN( u2_u9_u3_n117 ) , .A1( u2_u9_u3_n124 ) , .A2( u2_u9_u3_n148 ) );
  NAND2_X1 u2_u9_u3_U26 (.ZN( u2_u9_u3_n143 ) , .A1( u2_u9_u3_n165 ) , .A2( u2_u9_u3_n167 ) );
  INV_X1 u2_u9_u3_U27 (.A( u2_u9_u3_n130 ) , .ZN( u2_u9_u3_n177 ) );
  INV_X1 u2_u9_u3_U28 (.A( u2_u9_u3_n128 ) , .ZN( u2_u9_u3_n176 ) );
  INV_X1 u2_u9_u3_U29 (.A( u2_u9_u3_n155 ) , .ZN( u2_u9_u3_n174 ) );
  INV_X1 u2_u9_u3_U3 (.A( u2_u9_u3_n129 ) , .ZN( u2_u9_u3_n183 ) );
  INV_X1 u2_u9_u3_U30 (.A( u2_u9_u3_n139 ) , .ZN( u2_u9_u3_n185 ) );
  NOR2_X1 u2_u9_u3_U31 (.ZN( u2_u9_u3_n135 ) , .A2( u2_u9_u3_n141 ) , .A1( u2_u9_u3_n169 ) );
  OAI222_X1 u2_u9_u3_U32 (.C2( u2_u9_u3_n107 ) , .A2( u2_u9_u3_n108 ) , .B1( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n138 ) , .B2( u2_u9_u3_n146 ) , .C1( u2_u9_u3_n154 ) , .A1( u2_u9_u3_n164 ) );
  NOR4_X1 u2_u9_u3_U33 (.A4( u2_u9_u3_n157 ) , .A3( u2_u9_u3_n158 ) , .A2( u2_u9_u3_n159 ) , .A1( u2_u9_u3_n160 ) , .ZN( u2_u9_u3_n161 ) );
  AOI21_X1 u2_u9_u3_U34 (.B2( u2_u9_u3_n152 ) , .B1( u2_u9_u3_n153 ) , .ZN( u2_u9_u3_n158 ) , .A( u2_u9_u3_n164 ) );
  AOI21_X1 u2_u9_u3_U35 (.A( u2_u9_u3_n154 ) , .B2( u2_u9_u3_n155 ) , .B1( u2_u9_u3_n156 ) , .ZN( u2_u9_u3_n157 ) );
  AOI21_X1 u2_u9_u3_U36 (.A( u2_u9_u3_n149 ) , .B2( u2_u9_u3_n150 ) , .B1( u2_u9_u3_n151 ) , .ZN( u2_u9_u3_n159 ) );
  AOI211_X1 u2_u9_u3_U37 (.ZN( u2_u9_u3_n109 ) , .A( u2_u9_u3_n119 ) , .C2( u2_u9_u3_n129 ) , .B( u2_u9_u3_n138 ) , .C1( u2_u9_u3_n141 ) );
  AOI211_X1 u2_u9_u3_U38 (.B( u2_u9_u3_n119 ) , .A( u2_u9_u3_n120 ) , .C2( u2_u9_u3_n121 ) , .ZN( u2_u9_u3_n122 ) , .C1( u2_u9_u3_n179 ) );
  INV_X1 u2_u9_u3_U39 (.A( u2_u9_u3_n156 ) , .ZN( u2_u9_u3_n179 ) );
  INV_X1 u2_u9_u3_U4 (.A( u2_u9_u3_n140 ) , .ZN( u2_u9_u3_n182 ) );
  OAI22_X1 u2_u9_u3_U40 (.B1( u2_u9_u3_n118 ) , .ZN( u2_u9_u3_n120 ) , .A1( u2_u9_u3_n135 ) , .B2( u2_u9_u3_n154 ) , .A2( u2_u9_u3_n178 ) );
  AND3_X1 u2_u9_u3_U41 (.ZN( u2_u9_u3_n118 ) , .A2( u2_u9_u3_n124 ) , .A1( u2_u9_u3_n144 ) , .A3( u2_u9_u3_n152 ) );
  INV_X1 u2_u9_u3_U42 (.A( u2_u9_u3_n121 ) , .ZN( u2_u9_u3_n164 ) );
  NAND2_X1 u2_u9_u3_U43 (.ZN( u2_u9_u3_n133 ) , .A1( u2_u9_u3_n154 ) , .A2( u2_u9_u3_n164 ) );
  OAI211_X1 u2_u9_u3_U44 (.B( u2_u9_u3_n127 ) , .ZN( u2_u9_u3_n139 ) , .C1( u2_u9_u3_n150 ) , .C2( u2_u9_u3_n154 ) , .A( u2_u9_u3_n184 ) );
  INV_X1 u2_u9_u3_U45 (.A( u2_u9_u3_n125 ) , .ZN( u2_u9_u3_n184 ) );
  AOI221_X1 u2_u9_u3_U46 (.A( u2_u9_u3_n126 ) , .ZN( u2_u9_u3_n127 ) , .C2( u2_u9_u3_n132 ) , .C1( u2_u9_u3_n169 ) , .B2( u2_u9_u3_n170 ) , .B1( u2_u9_u3_n174 ) );
  OAI22_X1 u2_u9_u3_U47 (.A1( u2_u9_u3_n124 ) , .ZN( u2_u9_u3_n125 ) , .B2( u2_u9_u3_n145 ) , .A2( u2_u9_u3_n165 ) , .B1( u2_u9_u3_n167 ) );
  NOR2_X1 u2_u9_u3_U48 (.A1( u2_u9_u3_n113 ) , .ZN( u2_u9_u3_n131 ) , .A2( u2_u9_u3_n154 ) );
  NAND2_X1 u2_u9_u3_U49 (.A1( u2_u9_u3_n103 ) , .ZN( u2_u9_u3_n150 ) , .A2( u2_u9_u3_n99 ) );
  INV_X1 u2_u9_u3_U5 (.A( u2_u9_u3_n117 ) , .ZN( u2_u9_u3_n178 ) );
  NAND2_X1 u2_u9_u3_U50 (.A2( u2_u9_u3_n102 ) , .ZN( u2_u9_u3_n155 ) , .A1( u2_u9_u3_n97 ) );
  INV_X1 u2_u9_u3_U51 (.A( u2_u9_u3_n141 ) , .ZN( u2_u9_u3_n167 ) );
  AOI21_X1 u2_u9_u3_U52 (.B2( u2_u9_u3_n114 ) , .B1( u2_u9_u3_n146 ) , .A( u2_u9_u3_n154 ) , .ZN( u2_u9_u3_n94 ) );
  AOI21_X1 u2_u9_u3_U53 (.ZN( u2_u9_u3_n110 ) , .B2( u2_u9_u3_n142 ) , .B1( u2_u9_u3_n186 ) , .A( u2_u9_u3_n95 ) );
  INV_X1 u2_u9_u3_U54 (.A( u2_u9_u3_n145 ) , .ZN( u2_u9_u3_n186 ) );
  AOI21_X1 u2_u9_u3_U55 (.B1( u2_u9_u3_n124 ) , .A( u2_u9_u3_n149 ) , .B2( u2_u9_u3_n155 ) , .ZN( u2_u9_u3_n95 ) );
  INV_X1 u2_u9_u3_U56 (.A( u2_u9_u3_n149 ) , .ZN( u2_u9_u3_n169 ) );
  NAND2_X1 u2_u9_u3_U57 (.ZN( u2_u9_u3_n124 ) , .A1( u2_u9_u3_n96 ) , .A2( u2_u9_u3_n97 ) );
  NAND2_X1 u2_u9_u3_U58 (.A2( u2_u9_u3_n100 ) , .ZN( u2_u9_u3_n146 ) , .A1( u2_u9_u3_n96 ) );
  NAND2_X1 u2_u9_u3_U59 (.A1( u2_u9_u3_n101 ) , .ZN( u2_u9_u3_n145 ) , .A2( u2_u9_u3_n99 ) );
  AOI221_X1 u2_u9_u3_U6 (.A( u2_u9_u3_n131 ) , .C2( u2_u9_u3_n132 ) , .C1( u2_u9_u3_n133 ) , .ZN( u2_u9_u3_n134 ) , .B1( u2_u9_u3_n143 ) , .B2( u2_u9_u3_n177 ) );
  NAND2_X1 u2_u9_u3_U60 (.A1( u2_u9_u3_n100 ) , .ZN( u2_u9_u3_n156 ) , .A2( u2_u9_u3_n99 ) );
  NAND2_X1 u2_u9_u3_U61 (.A2( u2_u9_u3_n101 ) , .A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n148 ) );
  NAND2_X1 u2_u9_u3_U62 (.A1( u2_u9_u3_n100 ) , .A2( u2_u9_u3_n102 ) , .ZN( u2_u9_u3_n128 ) );
  NAND2_X1 u2_u9_u3_U63 (.A2( u2_u9_u3_n101 ) , .A1( u2_u9_u3_n102 ) , .ZN( u2_u9_u3_n152 ) );
  NAND2_X1 u2_u9_u3_U64 (.A2( u2_u9_u3_n101 ) , .ZN( u2_u9_u3_n114 ) , .A1( u2_u9_u3_n96 ) );
  NAND2_X1 u2_u9_u3_U65 (.ZN( u2_u9_u3_n107 ) , .A1( u2_u9_u3_n97 ) , .A2( u2_u9_u3_n99 ) );
  NAND2_X1 u2_u9_u3_U66 (.A2( u2_u9_u3_n100 ) , .A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n113 ) );
  NAND2_X1 u2_u9_u3_U67 (.A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n153 ) , .A2( u2_u9_u3_n97 ) );
  NAND2_X1 u2_u9_u3_U68 (.A2( u2_u9_u3_n103 ) , .A1( u2_u9_u3_n104 ) , .ZN( u2_u9_u3_n130 ) );
  NAND2_X1 u2_u9_u3_U69 (.A2( u2_u9_u3_n103 ) , .ZN( u2_u9_u3_n144 ) , .A1( u2_u9_u3_n96 ) );
  OAI22_X1 u2_u9_u3_U7 (.B2( u2_u9_u3_n147 ) , .A2( u2_u9_u3_n148 ) , .ZN( u2_u9_u3_n160 ) , .B1( u2_u9_u3_n165 ) , .A1( u2_u9_u3_n168 ) );
  NAND2_X1 u2_u9_u3_U70 (.A1( u2_u9_u3_n102 ) , .A2( u2_u9_u3_n103 ) , .ZN( u2_u9_u3_n108 ) );
  NOR2_X1 u2_u9_u3_U71 (.A2( u2_u9_X_19 ) , .A1( u2_u9_X_20 ) , .ZN( u2_u9_u3_n99 ) );
  NOR2_X1 u2_u9_u3_U72 (.A2( u2_u9_X_21 ) , .A1( u2_u9_X_24 ) , .ZN( u2_u9_u3_n103 ) );
  NOR2_X1 u2_u9_u3_U73 (.A2( u2_u9_X_24 ) , .A1( u2_u9_u3_n171 ) , .ZN( u2_u9_u3_n97 ) );
  NOR2_X1 u2_u9_u3_U74 (.A2( u2_u9_X_23 ) , .ZN( u2_u9_u3_n141 ) , .A1( u2_u9_u3_n166 ) );
  NOR2_X1 u2_u9_u3_U75 (.A2( u2_u9_X_19 ) , .A1( u2_u9_u3_n172 ) , .ZN( u2_u9_u3_n96 ) );
  NAND2_X1 u2_u9_u3_U76 (.A1( u2_u9_X_22 ) , .A2( u2_u9_X_23 ) , .ZN( u2_u9_u3_n154 ) );
  NAND2_X1 u2_u9_u3_U77 (.A1( u2_u9_X_23 ) , .ZN( u2_u9_u3_n149 ) , .A2( u2_u9_u3_n166 ) );
  NOR2_X1 u2_u9_u3_U78 (.A2( u2_u9_X_22 ) , .A1( u2_u9_X_23 ) , .ZN( u2_u9_u3_n121 ) );
  AND2_X1 u2_u9_u3_U79 (.A1( u2_u9_X_24 ) , .ZN( u2_u9_u3_n101 ) , .A2( u2_u9_u3_n171 ) );
  AND3_X1 u2_u9_u3_U8 (.A3( u2_u9_u3_n144 ) , .A2( u2_u9_u3_n145 ) , .A1( u2_u9_u3_n146 ) , .ZN( u2_u9_u3_n147 ) );
  AND2_X1 u2_u9_u3_U80 (.A1( u2_u9_X_19 ) , .ZN( u2_u9_u3_n102 ) , .A2( u2_u9_u3_n172 ) );
  AND2_X1 u2_u9_u3_U81 (.A1( u2_u9_X_21 ) , .A2( u2_u9_X_24 ) , .ZN( u2_u9_u3_n100 ) );
  AND2_X1 u2_u9_u3_U82 (.A2( u2_u9_X_19 ) , .A1( u2_u9_X_20 ) , .ZN( u2_u9_u3_n104 ) );
  INV_X1 u2_u9_u3_U83 (.A( u2_u9_X_22 ) , .ZN( u2_u9_u3_n166 ) );
  INV_X1 u2_u9_u3_U84 (.A( u2_u9_X_21 ) , .ZN( u2_u9_u3_n171 ) );
  INV_X1 u2_u9_u3_U85 (.A( u2_u9_X_20 ) , .ZN( u2_u9_u3_n172 ) );
  OR4_X1 u2_u9_u3_U86 (.ZN( u2_out9_10 ) , .A4( u2_u9_u3_n136 ) , .A3( u2_u9_u3_n137 ) , .A1( u2_u9_u3_n138 ) , .A2( u2_u9_u3_n139 ) );
  OAI222_X1 u2_u9_u3_U87 (.C1( u2_u9_u3_n128 ) , .ZN( u2_u9_u3_n137 ) , .B1( u2_u9_u3_n148 ) , .A2( u2_u9_u3_n150 ) , .B2( u2_u9_u3_n154 ) , .C2( u2_u9_u3_n164 ) , .A1( u2_u9_u3_n167 ) );
  OAI221_X1 u2_u9_u3_U88 (.A( u2_u9_u3_n134 ) , .B2( u2_u9_u3_n135 ) , .ZN( u2_u9_u3_n136 ) , .C1( u2_u9_u3_n149 ) , .B1( u2_u9_u3_n151 ) , .C2( u2_u9_u3_n183 ) );
  NAND4_X1 u2_u9_u3_U89 (.ZN( u2_out9_26 ) , .A4( u2_u9_u3_n109 ) , .A3( u2_u9_u3_n110 ) , .A2( u2_u9_u3_n111 ) , .A1( u2_u9_u3_n173 ) );
  INV_X1 u2_u9_u3_U9 (.A( u2_u9_u3_n143 ) , .ZN( u2_u9_u3_n168 ) );
  INV_X1 u2_u9_u3_U90 (.ZN( u2_u9_u3_n173 ) , .A( u2_u9_u3_n94 ) );
  OAI21_X1 u2_u9_u3_U91 (.ZN( u2_u9_u3_n111 ) , .B2( u2_u9_u3_n117 ) , .A( u2_u9_u3_n133 ) , .B1( u2_u9_u3_n176 ) );
  NAND4_X1 u2_u9_u3_U92 (.ZN( u2_out9_20 ) , .A4( u2_u9_u3_n122 ) , .A3( u2_u9_u3_n123 ) , .A1( u2_u9_u3_n175 ) , .A2( u2_u9_u3_n180 ) );
  INV_X1 u2_u9_u3_U93 (.A( u2_u9_u3_n126 ) , .ZN( u2_u9_u3_n180 ) );
  INV_X1 u2_u9_u3_U94 (.A( u2_u9_u3_n112 ) , .ZN( u2_u9_u3_n175 ) );
  NAND4_X1 u2_u9_u3_U95 (.ZN( u2_out9_1 ) , .A4( u2_u9_u3_n161 ) , .A3( u2_u9_u3_n162 ) , .A2( u2_u9_u3_n163 ) , .A1( u2_u9_u3_n185 ) );
  NAND2_X1 u2_u9_u3_U96 (.ZN( u2_u9_u3_n163 ) , .A2( u2_u9_u3_n170 ) , .A1( u2_u9_u3_n176 ) );
  AOI22_X1 u2_u9_u3_U97 (.B2( u2_u9_u3_n140 ) , .B1( u2_u9_u3_n141 ) , .A2( u2_u9_u3_n142 ) , .ZN( u2_u9_u3_n162 ) , .A1( u2_u9_u3_n177 ) );
  NAND3_X1 u2_u9_u3_U98 (.A1( u2_u9_u3_n114 ) , .ZN( u2_u9_u3_n115 ) , .A2( u2_u9_u3_n145 ) , .A3( u2_u9_u3_n153 ) );
  NAND3_X1 u2_u9_u3_U99 (.ZN( u2_u9_u3_n129 ) , .A2( u2_u9_u3_n144 ) , .A1( u2_u9_u3_n153 ) , .A3( u2_u9_u3_n182 ) );
  OAI22_X1 u2_u9_u4_U10 (.B2( u2_u9_u4_n135 ) , .ZN( u2_u9_u4_n137 ) , .B1( u2_u9_u4_n153 ) , .A1( u2_u9_u4_n155 ) , .A2( u2_u9_u4_n171 ) );
  AND3_X1 u2_u9_u4_U11 (.A2( u2_u9_u4_n134 ) , .ZN( u2_u9_u4_n135 ) , .A3( u2_u9_u4_n145 ) , .A1( u2_u9_u4_n157 ) );
  NAND2_X1 u2_u9_u4_U12 (.ZN( u2_u9_u4_n132 ) , .A2( u2_u9_u4_n170 ) , .A1( u2_u9_u4_n173 ) );
  AOI21_X1 u2_u9_u4_U13 (.B2( u2_u9_u4_n160 ) , .B1( u2_u9_u4_n161 ) , .ZN( u2_u9_u4_n162 ) , .A( u2_u9_u4_n170 ) );
  AOI21_X1 u2_u9_u4_U14 (.ZN( u2_u9_u4_n107 ) , .B2( u2_u9_u4_n143 ) , .A( u2_u9_u4_n174 ) , .B1( u2_u9_u4_n184 ) );
  AOI21_X1 u2_u9_u4_U15 (.B2( u2_u9_u4_n158 ) , .B1( u2_u9_u4_n159 ) , .ZN( u2_u9_u4_n163 ) , .A( u2_u9_u4_n174 ) );
  AOI21_X1 u2_u9_u4_U16 (.A( u2_u9_u4_n153 ) , .B2( u2_u9_u4_n154 ) , .B1( u2_u9_u4_n155 ) , .ZN( u2_u9_u4_n165 ) );
  AOI21_X1 u2_u9_u4_U17 (.A( u2_u9_u4_n156 ) , .B2( u2_u9_u4_n157 ) , .ZN( u2_u9_u4_n164 ) , .B1( u2_u9_u4_n184 ) );
  INV_X1 u2_u9_u4_U18 (.A( u2_u9_u4_n138 ) , .ZN( u2_u9_u4_n170 ) );
  AND2_X1 u2_u9_u4_U19 (.A2( u2_u9_u4_n120 ) , .ZN( u2_u9_u4_n155 ) , .A1( u2_u9_u4_n160 ) );
  INV_X1 u2_u9_u4_U20 (.A( u2_u9_u4_n156 ) , .ZN( u2_u9_u4_n175 ) );
  NAND2_X1 u2_u9_u4_U21 (.A2( u2_u9_u4_n118 ) , .ZN( u2_u9_u4_n131 ) , .A1( u2_u9_u4_n147 ) );
  NAND2_X1 u2_u9_u4_U22 (.A1( u2_u9_u4_n119 ) , .A2( u2_u9_u4_n120 ) , .ZN( u2_u9_u4_n130 ) );
  NAND2_X1 u2_u9_u4_U23 (.ZN( u2_u9_u4_n117 ) , .A2( u2_u9_u4_n118 ) , .A1( u2_u9_u4_n148 ) );
  NAND2_X1 u2_u9_u4_U24 (.ZN( u2_u9_u4_n129 ) , .A1( u2_u9_u4_n134 ) , .A2( u2_u9_u4_n148 ) );
  AND3_X1 u2_u9_u4_U25 (.A1( u2_u9_u4_n119 ) , .A2( u2_u9_u4_n143 ) , .A3( u2_u9_u4_n154 ) , .ZN( u2_u9_u4_n161 ) );
  AND2_X1 u2_u9_u4_U26 (.A1( u2_u9_u4_n145 ) , .A2( u2_u9_u4_n147 ) , .ZN( u2_u9_u4_n159 ) );
  OR3_X1 u2_u9_u4_U27 (.A3( u2_u9_u4_n114 ) , .A2( u2_u9_u4_n115 ) , .A1( u2_u9_u4_n116 ) , .ZN( u2_u9_u4_n136 ) );
  AOI21_X1 u2_u9_u4_U28 (.A( u2_u9_u4_n113 ) , .ZN( u2_u9_u4_n116 ) , .B2( u2_u9_u4_n173 ) , .B1( u2_u9_u4_n174 ) );
  AOI21_X1 u2_u9_u4_U29 (.ZN( u2_u9_u4_n115 ) , .B2( u2_u9_u4_n145 ) , .B1( u2_u9_u4_n146 ) , .A( u2_u9_u4_n156 ) );
  NOR2_X1 u2_u9_u4_U3 (.ZN( u2_u9_u4_n121 ) , .A1( u2_u9_u4_n181 ) , .A2( u2_u9_u4_n182 ) );
  OAI22_X1 u2_u9_u4_U30 (.ZN( u2_u9_u4_n114 ) , .A2( u2_u9_u4_n121 ) , .B1( u2_u9_u4_n160 ) , .B2( u2_u9_u4_n170 ) , .A1( u2_u9_u4_n171 ) );
  INV_X1 u2_u9_u4_U31 (.A( u2_u9_u4_n158 ) , .ZN( u2_u9_u4_n182 ) );
  INV_X1 u2_u9_u4_U32 (.ZN( u2_u9_u4_n181 ) , .A( u2_u9_u4_n96 ) );
  INV_X1 u2_u9_u4_U33 (.A( u2_u9_u4_n144 ) , .ZN( u2_u9_u4_n179 ) );
  INV_X1 u2_u9_u4_U34 (.A( u2_u9_u4_n157 ) , .ZN( u2_u9_u4_n178 ) );
  NAND2_X1 u2_u9_u4_U35 (.A2( u2_u9_u4_n154 ) , .A1( u2_u9_u4_n96 ) , .ZN( u2_u9_u4_n97 ) );
  INV_X1 u2_u9_u4_U36 (.ZN( u2_u9_u4_n186 ) , .A( u2_u9_u4_n95 ) );
  OAI221_X1 u2_u9_u4_U37 (.C1( u2_u9_u4_n134 ) , .B1( u2_u9_u4_n158 ) , .B2( u2_u9_u4_n171 ) , .C2( u2_u9_u4_n173 ) , .A( u2_u9_u4_n94 ) , .ZN( u2_u9_u4_n95 ) );
  AOI222_X1 u2_u9_u4_U38 (.B2( u2_u9_u4_n132 ) , .A1( u2_u9_u4_n138 ) , .C2( u2_u9_u4_n175 ) , .A2( u2_u9_u4_n179 ) , .C1( u2_u9_u4_n181 ) , .B1( u2_u9_u4_n185 ) , .ZN( u2_u9_u4_n94 ) );
  INV_X1 u2_u9_u4_U39 (.A( u2_u9_u4_n113 ) , .ZN( u2_u9_u4_n185 ) );
  INV_X1 u2_u9_u4_U4 (.A( u2_u9_u4_n117 ) , .ZN( u2_u9_u4_n184 ) );
  INV_X1 u2_u9_u4_U40 (.A( u2_u9_u4_n143 ) , .ZN( u2_u9_u4_n183 ) );
  NOR2_X1 u2_u9_u4_U41 (.ZN( u2_u9_u4_n138 ) , .A1( u2_u9_u4_n168 ) , .A2( u2_u9_u4_n169 ) );
  NOR2_X1 u2_u9_u4_U42 (.A1( u2_u9_u4_n150 ) , .A2( u2_u9_u4_n152 ) , .ZN( u2_u9_u4_n153 ) );
  NOR2_X1 u2_u9_u4_U43 (.A2( u2_u9_u4_n128 ) , .A1( u2_u9_u4_n138 ) , .ZN( u2_u9_u4_n156 ) );
  AOI22_X1 u2_u9_u4_U44 (.B2( u2_u9_u4_n122 ) , .A1( u2_u9_u4_n123 ) , .ZN( u2_u9_u4_n124 ) , .B1( u2_u9_u4_n128 ) , .A2( u2_u9_u4_n172 ) );
  INV_X1 u2_u9_u4_U45 (.A( u2_u9_u4_n153 ) , .ZN( u2_u9_u4_n172 ) );
  NAND2_X1 u2_u9_u4_U46 (.A2( u2_u9_u4_n120 ) , .ZN( u2_u9_u4_n123 ) , .A1( u2_u9_u4_n161 ) );
  AOI22_X1 u2_u9_u4_U47 (.B2( u2_u9_u4_n132 ) , .A2( u2_u9_u4_n133 ) , .ZN( u2_u9_u4_n140 ) , .A1( u2_u9_u4_n150 ) , .B1( u2_u9_u4_n179 ) );
  NAND2_X1 u2_u9_u4_U48 (.ZN( u2_u9_u4_n133 ) , .A2( u2_u9_u4_n146 ) , .A1( u2_u9_u4_n154 ) );
  NAND2_X1 u2_u9_u4_U49 (.A1( u2_u9_u4_n103 ) , .ZN( u2_u9_u4_n154 ) , .A2( u2_u9_u4_n98 ) );
  NOR4_X1 u2_u9_u4_U5 (.A4( u2_u9_u4_n106 ) , .A3( u2_u9_u4_n107 ) , .A2( u2_u9_u4_n108 ) , .A1( u2_u9_u4_n109 ) , .ZN( u2_u9_u4_n110 ) );
  NAND2_X1 u2_u9_u4_U50 (.A1( u2_u9_u4_n101 ) , .ZN( u2_u9_u4_n158 ) , .A2( u2_u9_u4_n99 ) );
  AOI21_X1 u2_u9_u4_U51 (.ZN( u2_u9_u4_n127 ) , .A( u2_u9_u4_n136 ) , .B2( u2_u9_u4_n150 ) , .B1( u2_u9_u4_n180 ) );
  INV_X1 u2_u9_u4_U52 (.A( u2_u9_u4_n160 ) , .ZN( u2_u9_u4_n180 ) );
  NAND2_X1 u2_u9_u4_U53 (.A2( u2_u9_u4_n104 ) , .A1( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n146 ) );
  NAND2_X1 u2_u9_u4_U54 (.A2( u2_u9_u4_n101 ) , .A1( u2_u9_u4_n102 ) , .ZN( u2_u9_u4_n160 ) );
  NAND2_X1 u2_u9_u4_U55 (.ZN( u2_u9_u4_n134 ) , .A1( u2_u9_u4_n98 ) , .A2( u2_u9_u4_n99 ) );
  NAND2_X1 u2_u9_u4_U56 (.A1( u2_u9_u4_n103 ) , .A2( u2_u9_u4_n104 ) , .ZN( u2_u9_u4_n143 ) );
  NAND2_X1 u2_u9_u4_U57 (.A2( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n145 ) , .A1( u2_u9_u4_n98 ) );
  NAND2_X1 u2_u9_u4_U58 (.A1( u2_u9_u4_n100 ) , .A2( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n120 ) );
  NAND2_X1 u2_u9_u4_U59 (.A1( u2_u9_u4_n102 ) , .A2( u2_u9_u4_n104 ) , .ZN( u2_u9_u4_n148 ) );
  AOI21_X1 u2_u9_u4_U6 (.ZN( u2_u9_u4_n106 ) , .B2( u2_u9_u4_n146 ) , .B1( u2_u9_u4_n158 ) , .A( u2_u9_u4_n170 ) );
  NAND2_X1 u2_u9_u4_U60 (.A2( u2_u9_u4_n100 ) , .A1( u2_u9_u4_n103 ) , .ZN( u2_u9_u4_n157 ) );
  INV_X1 u2_u9_u4_U61 (.A( u2_u9_u4_n150 ) , .ZN( u2_u9_u4_n173 ) );
  INV_X1 u2_u9_u4_U62 (.A( u2_u9_u4_n152 ) , .ZN( u2_u9_u4_n171 ) );
  NAND2_X1 u2_u9_u4_U63 (.A1( u2_u9_u4_n100 ) , .ZN( u2_u9_u4_n118 ) , .A2( u2_u9_u4_n99 ) );
  NAND2_X1 u2_u9_u4_U64 (.A2( u2_u9_u4_n100 ) , .A1( u2_u9_u4_n102 ) , .ZN( u2_u9_u4_n144 ) );
  NAND2_X1 u2_u9_u4_U65 (.A2( u2_u9_u4_n101 ) , .A1( u2_u9_u4_n105 ) , .ZN( u2_u9_u4_n96 ) );
  INV_X1 u2_u9_u4_U66 (.A( u2_u9_u4_n128 ) , .ZN( u2_u9_u4_n174 ) );
  NAND2_X1 u2_u9_u4_U67 (.A2( u2_u9_u4_n102 ) , .ZN( u2_u9_u4_n119 ) , .A1( u2_u9_u4_n98 ) );
  NAND2_X1 u2_u9_u4_U68 (.A2( u2_u9_u4_n101 ) , .A1( u2_u9_u4_n103 ) , .ZN( u2_u9_u4_n147 ) );
  NAND2_X1 u2_u9_u4_U69 (.A2( u2_u9_u4_n104 ) , .ZN( u2_u9_u4_n113 ) , .A1( u2_u9_u4_n99 ) );
  AOI21_X1 u2_u9_u4_U7 (.ZN( u2_u9_u4_n108 ) , .B2( u2_u9_u4_n134 ) , .B1( u2_u9_u4_n155 ) , .A( u2_u9_u4_n156 ) );
  NOR2_X1 u2_u9_u4_U70 (.A2( u2_u9_X_28 ) , .ZN( u2_u9_u4_n150 ) , .A1( u2_u9_u4_n168 ) );
  NOR2_X1 u2_u9_u4_U71 (.A2( u2_u9_X_29 ) , .ZN( u2_u9_u4_n152 ) , .A1( u2_u9_u4_n169 ) );
  NOR2_X1 u2_u9_u4_U72 (.A2( u2_u9_X_30 ) , .ZN( u2_u9_u4_n105 ) , .A1( u2_u9_u4_n176 ) );
  NOR2_X1 u2_u9_u4_U73 (.A2( u2_u9_X_26 ) , .ZN( u2_u9_u4_n100 ) , .A1( u2_u9_u4_n177 ) );
  NOR2_X1 u2_u9_u4_U74 (.A2( u2_u9_X_28 ) , .A1( u2_u9_X_29 ) , .ZN( u2_u9_u4_n128 ) );
  NOR2_X1 u2_u9_u4_U75 (.A2( u2_u9_X_27 ) , .A1( u2_u9_X_30 ) , .ZN( u2_u9_u4_n102 ) );
  NOR2_X1 u2_u9_u4_U76 (.A2( u2_u9_X_25 ) , .A1( u2_u9_X_26 ) , .ZN( u2_u9_u4_n98 ) );
  AND2_X1 u2_u9_u4_U77 (.A2( u2_u9_X_25 ) , .A1( u2_u9_X_26 ) , .ZN( u2_u9_u4_n104 ) );
  AND2_X1 u2_u9_u4_U78 (.A1( u2_u9_X_30 ) , .A2( u2_u9_u4_n176 ) , .ZN( u2_u9_u4_n99 ) );
  AND2_X1 u2_u9_u4_U79 (.A1( u2_u9_X_26 ) , .ZN( u2_u9_u4_n101 ) , .A2( u2_u9_u4_n177 ) );
  AOI21_X1 u2_u9_u4_U8 (.ZN( u2_u9_u4_n109 ) , .A( u2_u9_u4_n153 ) , .B1( u2_u9_u4_n159 ) , .B2( u2_u9_u4_n184 ) );
  AND2_X1 u2_u9_u4_U80 (.A1( u2_u9_X_27 ) , .A2( u2_u9_X_30 ) , .ZN( u2_u9_u4_n103 ) );
  INV_X1 u2_u9_u4_U81 (.A( u2_u9_X_28 ) , .ZN( u2_u9_u4_n169 ) );
  INV_X1 u2_u9_u4_U82 (.A( u2_u9_X_29 ) , .ZN( u2_u9_u4_n168 ) );
  INV_X1 u2_u9_u4_U83 (.A( u2_u9_X_25 ) , .ZN( u2_u9_u4_n177 ) );
  INV_X1 u2_u9_u4_U84 (.A( u2_u9_X_27 ) , .ZN( u2_u9_u4_n176 ) );
  NAND4_X1 u2_u9_u4_U85 (.ZN( u2_out9_25 ) , .A4( u2_u9_u4_n139 ) , .A3( u2_u9_u4_n140 ) , .A2( u2_u9_u4_n141 ) , .A1( u2_u9_u4_n142 ) );
  OAI21_X1 u2_u9_u4_U86 (.A( u2_u9_u4_n128 ) , .B2( u2_u9_u4_n129 ) , .B1( u2_u9_u4_n130 ) , .ZN( u2_u9_u4_n142 ) );
  OAI21_X1 u2_u9_u4_U87 (.B2( u2_u9_u4_n131 ) , .ZN( u2_u9_u4_n141 ) , .A( u2_u9_u4_n175 ) , .B1( u2_u9_u4_n183 ) );
  NAND4_X1 u2_u9_u4_U88 (.ZN( u2_out9_14 ) , .A4( u2_u9_u4_n124 ) , .A3( u2_u9_u4_n125 ) , .A2( u2_u9_u4_n126 ) , .A1( u2_u9_u4_n127 ) );
  AOI22_X1 u2_u9_u4_U89 (.B2( u2_u9_u4_n117 ) , .ZN( u2_u9_u4_n126 ) , .A1( u2_u9_u4_n129 ) , .B1( u2_u9_u4_n152 ) , .A2( u2_u9_u4_n175 ) );
  AOI211_X1 u2_u9_u4_U9 (.B( u2_u9_u4_n136 ) , .A( u2_u9_u4_n137 ) , .C2( u2_u9_u4_n138 ) , .ZN( u2_u9_u4_n139 ) , .C1( u2_u9_u4_n182 ) );
  AOI22_X1 u2_u9_u4_U90 (.ZN( u2_u9_u4_n125 ) , .B2( u2_u9_u4_n131 ) , .A2( u2_u9_u4_n132 ) , .B1( u2_u9_u4_n138 ) , .A1( u2_u9_u4_n178 ) );
  NAND4_X1 u2_u9_u4_U91 (.ZN( u2_out9_8 ) , .A4( u2_u9_u4_n110 ) , .A3( u2_u9_u4_n111 ) , .A2( u2_u9_u4_n112 ) , .A1( u2_u9_u4_n186 ) );
  NAND2_X1 u2_u9_u4_U92 (.ZN( u2_u9_u4_n112 ) , .A2( u2_u9_u4_n130 ) , .A1( u2_u9_u4_n150 ) );
  AOI22_X1 u2_u9_u4_U93 (.ZN( u2_u9_u4_n111 ) , .B2( u2_u9_u4_n132 ) , .A1( u2_u9_u4_n152 ) , .B1( u2_u9_u4_n178 ) , .A2( u2_u9_u4_n97 ) );
  AOI22_X1 u2_u9_u4_U94 (.B2( u2_u9_u4_n149 ) , .B1( u2_u9_u4_n150 ) , .A2( u2_u9_u4_n151 ) , .A1( u2_u9_u4_n152 ) , .ZN( u2_u9_u4_n167 ) );
  NOR4_X1 u2_u9_u4_U95 (.A4( u2_u9_u4_n162 ) , .A3( u2_u9_u4_n163 ) , .A2( u2_u9_u4_n164 ) , .A1( u2_u9_u4_n165 ) , .ZN( u2_u9_u4_n166 ) );
  NAND3_X1 u2_u9_u4_U96 (.ZN( u2_out9_3 ) , .A3( u2_u9_u4_n166 ) , .A1( u2_u9_u4_n167 ) , .A2( u2_u9_u4_n186 ) );
  NAND3_X1 u2_u9_u4_U97 (.A3( u2_u9_u4_n146 ) , .A2( u2_u9_u4_n147 ) , .A1( u2_u9_u4_n148 ) , .ZN( u2_u9_u4_n149 ) );
  NAND3_X1 u2_u9_u4_U98 (.A3( u2_u9_u4_n143 ) , .A2( u2_u9_u4_n144 ) , .A1( u2_u9_u4_n145 ) , .ZN( u2_u9_u4_n151 ) );
  NAND3_X1 u2_u9_u4_U99 (.A3( u2_u9_u4_n121 ) , .ZN( u2_u9_u4_n122 ) , .A2( u2_u9_u4_n144 ) , .A1( u2_u9_u4_n154 ) );
  NOR2_X1 u2_u9_u5_U10 (.ZN( u2_u9_u5_n135 ) , .A1( u2_u9_u5_n173 ) , .A2( u2_u9_u5_n176 ) );
  NOR3_X1 u2_u9_u5_U100 (.A3( u2_u9_u5_n141 ) , .A1( u2_u9_u5_n142 ) , .ZN( u2_u9_u5_n143 ) , .A2( u2_u9_u5_n191 ) );
  NAND4_X1 u2_u9_u5_U101 (.ZN( u2_out9_4 ) , .A4( u2_u9_u5_n112 ) , .A2( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n114 ) , .A3( u2_u9_u5_n195 ) );
  AOI211_X1 u2_u9_u5_U102 (.A( u2_u9_u5_n110 ) , .C1( u2_u9_u5_n111 ) , .ZN( u2_u9_u5_n112 ) , .B( u2_u9_u5_n118 ) , .C2( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U103 (.A( u2_u9_u5_n102 ) , .ZN( u2_u9_u5_n195 ) );
  NAND3_X1 u2_u9_u5_U104 (.A2( u2_u9_u5_n154 ) , .A3( u2_u9_u5_n158 ) , .A1( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n99 ) );
  INV_X1 u2_u9_u5_U11 (.A( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U12 (.ZN( u2_u9_u5_n160 ) , .A2( u2_u9_u5_n173 ) , .A1( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U13 (.A( u2_u9_u5_n150 ) , .ZN( u2_u9_u5_n174 ) );
  AOI21_X1 u2_u9_u5_U14 (.A( u2_u9_u5_n160 ) , .B2( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n162 ) , .B1( u2_u9_u5_n192 ) );
  INV_X1 u2_u9_u5_U15 (.A( u2_u9_u5_n159 ) , .ZN( u2_u9_u5_n192 ) );
  AOI21_X1 u2_u9_u5_U16 (.A( u2_u9_u5_n156 ) , .B2( u2_u9_u5_n157 ) , .B1( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n163 ) );
  AOI21_X1 u2_u9_u5_U17 (.B2( u2_u9_u5_n139 ) , .B1( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n141 ) , .A( u2_u9_u5_n150 ) );
  OAI21_X1 u2_u9_u5_U18 (.A( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n134 ) , .B1( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n142 ) );
  OAI21_X1 u2_u9_u5_U19 (.ZN( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n147 ) , .A( u2_u9_u5_n173 ) , .B1( u2_u9_u5_n188 ) );
  NAND2_X1 u2_u9_u5_U20 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n137 ) );
  INV_X1 u2_u9_u5_U21 (.A( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n194 ) );
  NAND2_X1 u2_u9_u5_U22 (.A1( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n132 ) , .A2( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U23 (.A2( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n136 ) , .A1( u2_u9_u5_n154 ) );
  NAND2_X1 u2_u9_u5_U24 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n159 ) );
  INV_X1 u2_u9_u5_U25 (.A( u2_u9_u5_n156 ) , .ZN( u2_u9_u5_n175 ) );
  INV_X1 u2_u9_u5_U26 (.A( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n188 ) );
  INV_X1 u2_u9_u5_U27 (.A( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n179 ) );
  INV_X1 u2_u9_u5_U28 (.A( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n182 ) );
  INV_X1 u2_u9_u5_U29 (.A( u2_u9_u5_n151 ) , .ZN( u2_u9_u5_n183 ) );
  NOR2_X1 u2_u9_u5_U3 (.ZN( u2_u9_u5_n134 ) , .A1( u2_u9_u5_n183 ) , .A2( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U30 (.A( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n185 ) );
  INV_X1 u2_u9_u5_U31 (.A( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n184 ) );
  INV_X1 u2_u9_u5_U32 (.A( u2_u9_u5_n139 ) , .ZN( u2_u9_u5_n189 ) );
  INV_X1 u2_u9_u5_U33 (.A( u2_u9_u5_n157 ) , .ZN( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U34 (.A( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n193 ) );
  NAND2_X1 u2_u9_u5_U35 (.ZN( u2_u9_u5_n111 ) , .A1( u2_u9_u5_n140 ) , .A2( u2_u9_u5_n155 ) );
  NOR2_X1 u2_u9_u5_U36 (.ZN( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n170 ) , .A2( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U37 (.A( u2_u9_u5_n117 ) , .ZN( u2_u9_u5_n196 ) );
  OAI221_X1 u2_u9_u5_U38 (.A( u2_u9_u5_n116 ) , .ZN( u2_u9_u5_n117 ) , .B2( u2_u9_u5_n119 ) , .C1( u2_u9_u5_n153 ) , .C2( u2_u9_u5_n158 ) , .B1( u2_u9_u5_n172 ) );
  AOI222_X1 u2_u9_u5_U39 (.ZN( u2_u9_u5_n116 ) , .B2( u2_u9_u5_n145 ) , .C1( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n177 ) , .B1( u2_u9_u5_n187 ) , .A1( u2_u9_u5_n193 ) );
  INV_X1 u2_u9_u5_U4 (.A( u2_u9_u5_n138 ) , .ZN( u2_u9_u5_n191 ) );
  INV_X1 u2_u9_u5_U40 (.A( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n187 ) );
  OAI221_X1 u2_u9_u5_U41 (.A( u2_u9_u5_n101 ) , .ZN( u2_u9_u5_n102 ) , .C2( u2_u9_u5_n115 ) , .C1( u2_u9_u5_n126 ) , .B1( u2_u9_u5_n134 ) , .B2( u2_u9_u5_n160 ) );
  OAI21_X1 u2_u9_u5_U42 (.ZN( u2_u9_u5_n101 ) , .B1( u2_u9_u5_n137 ) , .A( u2_u9_u5_n146 ) , .B2( u2_u9_u5_n147 ) );
  AOI22_X1 u2_u9_u5_U43 (.B2( u2_u9_u5_n131 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n169 ) , .B1( u2_u9_u5_n174 ) , .A1( u2_u9_u5_n185 ) );
  NOR2_X1 u2_u9_u5_U44 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n173 ) );
  AOI21_X1 u2_u9_u5_U45 (.A( u2_u9_u5_n118 ) , .B2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n168 ) , .B1( u2_u9_u5_n186 ) );
  INV_X1 u2_u9_u5_U46 (.A( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n186 ) );
  NOR2_X1 u2_u9_u5_U47 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n152 ) , .A2( u2_u9_u5_n176 ) );
  NOR2_X1 u2_u9_u5_U48 (.A1( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n118 ) , .A2( u2_u9_u5_n153 ) );
  NOR2_X1 u2_u9_u5_U49 (.A2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n156 ) , .A1( u2_u9_u5_n174 ) );
  OAI21_X1 u2_u9_u5_U5 (.B2( u2_u9_u5_n136 ) , .B1( u2_u9_u5_n137 ) , .ZN( u2_u9_u5_n138 ) , .A( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U50 (.ZN( u2_u9_u5_n121 ) , .A2( u2_u9_u5_n145 ) , .A1( u2_u9_u5_n176 ) );
  AOI22_X1 u2_u9_u5_U51 (.ZN( u2_u9_u5_n114 ) , .A2( u2_u9_u5_n137 ) , .A1( u2_u9_u5_n145 ) , .B2( u2_u9_u5_n175 ) , .B1( u2_u9_u5_n193 ) );
  OAI211_X1 u2_u9_u5_U52 (.B( u2_u9_u5_n124 ) , .A( u2_u9_u5_n125 ) , .C2( u2_u9_u5_n126 ) , .C1( u2_u9_u5_n127 ) , .ZN( u2_u9_u5_n128 ) );
  NOR3_X1 u2_u9_u5_U53 (.ZN( u2_u9_u5_n127 ) , .A1( u2_u9_u5_n136 ) , .A3( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n182 ) );
  OAI21_X1 u2_u9_u5_U54 (.ZN( u2_u9_u5_n124 ) , .A( u2_u9_u5_n177 ) , .B2( u2_u9_u5_n183 ) , .B1( u2_u9_u5_n189 ) );
  OAI21_X1 u2_u9_u5_U55 (.ZN( u2_u9_u5_n125 ) , .A( u2_u9_u5_n174 ) , .B2( u2_u9_u5_n185 ) , .B1( u2_u9_u5_n190 ) );
  AOI21_X1 u2_u9_u5_U56 (.A( u2_u9_u5_n153 ) , .B2( u2_u9_u5_n154 ) , .B1( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n164 ) );
  AOI21_X1 u2_u9_u5_U57 (.ZN( u2_u9_u5_n110 ) , .B1( u2_u9_u5_n122 ) , .B2( u2_u9_u5_n139 ) , .A( u2_u9_u5_n153 ) );
  INV_X1 u2_u9_u5_U58 (.A( u2_u9_u5_n153 ) , .ZN( u2_u9_u5_n176 ) );
  INV_X1 u2_u9_u5_U59 (.A( u2_u9_u5_n126 ) , .ZN( u2_u9_u5_n173 ) );
  AOI222_X1 u2_u9_u5_U6 (.ZN( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n131 ) , .C1( u2_u9_u5_n148 ) , .B2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n178 ) , .A2( u2_u9_u5_n179 ) , .B1( u2_u9_u5_n99 ) );
  AND2_X1 u2_u9_u5_U60 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n147 ) );
  AND2_X1 u2_u9_u5_U61 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n148 ) );
  NAND2_X1 u2_u9_u5_U62 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n158 ) );
  NAND2_X1 u2_u9_u5_U63 (.A2( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n139 ) );
  NAND2_X1 u2_u9_u5_U64 (.A1( u2_u9_u5_n106 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n119 ) );
  NAND2_X1 u2_u9_u5_U65 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n140 ) );
  NAND2_X1 u2_u9_u5_U66 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n155 ) );
  NAND2_X1 u2_u9_u5_U67 (.A2( u2_u9_u5_n106 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n122 ) );
  NAND2_X1 u2_u9_u5_U68 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n115 ) );
  NAND2_X1 u2_u9_u5_U69 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n103 ) , .ZN( u2_u9_u5_n161 ) );
  INV_X1 u2_u9_u5_U7 (.A( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n178 ) );
  NAND2_X1 u2_u9_u5_U70 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n154 ) );
  INV_X1 u2_u9_u5_U71 (.A( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U72 (.A1( u2_u9_u5_n103 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n123 ) );
  NAND2_X1 u2_u9_u5_U73 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n151 ) );
  NAND2_X1 u2_u9_u5_U74 (.A2( u2_u9_u5_n107 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n120 ) );
  NAND2_X1 u2_u9_u5_U75 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n157 ) );
  AND2_X1 u2_u9_u5_U76 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n104 ) , .ZN( u2_u9_u5_n131 ) );
  NOR2_X1 u2_u9_u5_U77 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n145 ) );
  NOR2_X1 u2_u9_u5_U78 (.A2( u2_u9_X_34 ) , .ZN( u2_u9_u5_n146 ) , .A1( u2_u9_u5_n171 ) );
  NOR2_X1 u2_u9_u5_U79 (.A2( u2_u9_X_31 ) , .A1( u2_u9_X_32 ) , .ZN( u2_u9_u5_n103 ) );
  OAI22_X1 u2_u9_u5_U8 (.B2( u2_u9_u5_n149 ) , .B1( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n151 ) , .A1( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n165 ) );
  NOR2_X1 u2_u9_u5_U80 (.A2( u2_u9_X_36 ) , .ZN( u2_u9_u5_n105 ) , .A1( u2_u9_u5_n180 ) );
  NOR2_X1 u2_u9_u5_U81 (.A2( u2_u9_X_33 ) , .ZN( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n170 ) );
  NOR2_X1 u2_u9_u5_U82 (.A2( u2_u9_X_33 ) , .A1( u2_u9_X_36 ) , .ZN( u2_u9_u5_n107 ) );
  NOR2_X1 u2_u9_u5_U83 (.A2( u2_u9_X_31 ) , .ZN( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n181 ) );
  NAND2_X1 u2_u9_u5_U84 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n153 ) );
  NAND2_X1 u2_u9_u5_U85 (.A1( u2_u9_X_34 ) , .ZN( u2_u9_u5_n126 ) , .A2( u2_u9_u5_n171 ) );
  AND2_X1 u2_u9_u5_U86 (.A1( u2_u9_X_31 ) , .A2( u2_u9_X_32 ) , .ZN( u2_u9_u5_n106 ) );
  AND2_X1 u2_u9_u5_U87 (.A1( u2_u9_X_31 ) , .ZN( u2_u9_u5_n109 ) , .A2( u2_u9_u5_n181 ) );
  INV_X1 u2_u9_u5_U88 (.A( u2_u9_X_33 ) , .ZN( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U89 (.A( u2_u9_X_35 ) , .ZN( u2_u9_u5_n171 ) );
  NOR3_X1 u2_u9_u5_U9 (.A2( u2_u9_u5_n147 ) , .A1( u2_u9_u5_n148 ) , .ZN( u2_u9_u5_n149 ) , .A3( u2_u9_u5_n194 ) );
  INV_X1 u2_u9_u5_U90 (.A( u2_u9_X_36 ) , .ZN( u2_u9_u5_n170 ) );
  INV_X1 u2_u9_u5_U91 (.A( u2_u9_X_32 ) , .ZN( u2_u9_u5_n181 ) );
  NAND4_X1 u2_u9_u5_U92 (.ZN( u2_out9_29 ) , .A4( u2_u9_u5_n129 ) , .A3( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n196 ) );
  AOI221_X1 u2_u9_u5_U93 (.A( u2_u9_u5_n128 ) , .ZN( u2_u9_u5_n129 ) , .C2( u2_u9_u5_n132 ) , .B2( u2_u9_u5_n159 ) , .B1( u2_u9_u5_n176 ) , .C1( u2_u9_u5_n184 ) );
  AOI222_X1 u2_u9_u5_U94 (.ZN( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n146 ) , .B1( u2_u9_u5_n147 ) , .C2( u2_u9_u5_n175 ) , .B2( u2_u9_u5_n179 ) , .A1( u2_u9_u5_n188 ) , .C1( u2_u9_u5_n194 ) );
  NAND4_X1 u2_u9_u5_U95 (.ZN( u2_out9_19 ) , .A4( u2_u9_u5_n166 ) , .A3( u2_u9_u5_n167 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n169 ) );
  AOI22_X1 u2_u9_u5_U96 (.B2( u2_u9_u5_n145 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n167 ) , .B1( u2_u9_u5_n182 ) , .A1( u2_u9_u5_n189 ) );
  NOR4_X1 u2_u9_u5_U97 (.A4( u2_u9_u5_n162 ) , .A3( u2_u9_u5_n163 ) , .A2( u2_u9_u5_n164 ) , .A1( u2_u9_u5_n165 ) , .ZN( u2_u9_u5_n166 ) );
  NAND4_X1 u2_u9_u5_U98 (.ZN( u2_out9_11 ) , .A4( u2_u9_u5_n143 ) , .A3( u2_u9_u5_n144 ) , .A2( u2_u9_u5_n169 ) , .A1( u2_u9_u5_n196 ) );
  AOI22_X1 u2_u9_u5_U99 (.A2( u2_u9_u5_n132 ) , .ZN( u2_u9_u5_n144 ) , .B2( u2_u9_u5_n145 ) , .B1( u2_u9_u5_n184 ) , .A1( u2_u9_u5_n194 ) );
  AOI22_X1 u2_u9_u6_U10 (.A2( u2_u9_u6_n151 ) , .B2( u2_u9_u6_n161 ) , .A1( u2_u9_u6_n167 ) , .B1( u2_u9_u6_n170 ) , .ZN( u2_u9_u6_n89 ) );
  AOI21_X1 u2_u9_u6_U11 (.B1( u2_u9_u6_n107 ) , .B2( u2_u9_u6_n132 ) , .A( u2_u9_u6_n158 ) , .ZN( u2_u9_u6_n88 ) );
  AOI21_X1 u2_u9_u6_U12 (.B2( u2_u9_u6_n147 ) , .B1( u2_u9_u6_n148 ) , .ZN( u2_u9_u6_n149 ) , .A( u2_u9_u6_n158 ) );
  AOI21_X1 u2_u9_u6_U13 (.ZN( u2_u9_u6_n106 ) , .A( u2_u9_u6_n142 ) , .B2( u2_u9_u6_n159 ) , .B1( u2_u9_u6_n164 ) );
  INV_X1 u2_u9_u6_U14 (.A( u2_u9_u6_n155 ) , .ZN( u2_u9_u6_n161 ) );
  INV_X1 u2_u9_u6_U15 (.A( u2_u9_u6_n128 ) , .ZN( u2_u9_u6_n164 ) );
  NAND2_X1 u2_u9_u6_U16 (.ZN( u2_u9_u6_n110 ) , .A1( u2_u9_u6_n122 ) , .A2( u2_u9_u6_n129 ) );
  NAND2_X1 u2_u9_u6_U17 (.ZN( u2_u9_u6_n124 ) , .A2( u2_u9_u6_n146 ) , .A1( u2_u9_u6_n148 ) );
  INV_X1 u2_u9_u6_U18 (.A( u2_u9_u6_n132 ) , .ZN( u2_u9_u6_n171 ) );
  AND2_X1 u2_u9_u6_U19 (.A1( u2_u9_u6_n100 ) , .ZN( u2_u9_u6_n130 ) , .A2( u2_u9_u6_n147 ) );
  INV_X1 u2_u9_u6_U20 (.A( u2_u9_u6_n127 ) , .ZN( u2_u9_u6_n173 ) );
  INV_X1 u2_u9_u6_U21 (.A( u2_u9_u6_n121 ) , .ZN( u2_u9_u6_n167 ) );
  INV_X1 u2_u9_u6_U22 (.A( u2_u9_u6_n100 ) , .ZN( u2_u9_u6_n169 ) );
  INV_X1 u2_u9_u6_U23 (.A( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n170 ) );
  INV_X1 u2_u9_u6_U24 (.A( u2_u9_u6_n113 ) , .ZN( u2_u9_u6_n168 ) );
  AND2_X1 u2_u9_u6_U25 (.A1( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n119 ) , .ZN( u2_u9_u6_n133 ) );
  AND2_X1 u2_u9_u6_U26 (.A2( u2_u9_u6_n121 ) , .A1( u2_u9_u6_n122 ) , .ZN( u2_u9_u6_n131 ) );
  AND3_X1 u2_u9_u6_U27 (.ZN( u2_u9_u6_n120 ) , .A2( u2_u9_u6_n127 ) , .A1( u2_u9_u6_n132 ) , .A3( u2_u9_u6_n145 ) );
  INV_X1 u2_u9_u6_U28 (.A( u2_u9_u6_n146 ) , .ZN( u2_u9_u6_n163 ) );
  AOI222_X1 u2_u9_u6_U29 (.ZN( u2_u9_u6_n114 ) , .A1( u2_u9_u6_n118 ) , .A2( u2_u9_u6_n126 ) , .B2( u2_u9_u6_n151 ) , .C2( u2_u9_u6_n159 ) , .C1( u2_u9_u6_n168 ) , .B1( u2_u9_u6_n169 ) );
  INV_X1 u2_u9_u6_U3 (.A( u2_u9_u6_n110 ) , .ZN( u2_u9_u6_n166 ) );
  NOR2_X1 u2_u9_u6_U30 (.A1( u2_u9_u6_n162 ) , .A2( u2_u9_u6_n165 ) , .ZN( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U31 (.A1( u2_u9_u6_n144 ) , .ZN( u2_u9_u6_n151 ) , .A2( u2_u9_u6_n158 ) );
  NAND2_X1 u2_u9_u6_U32 (.ZN( u2_u9_u6_n132 ) , .A1( u2_u9_u6_n91 ) , .A2( u2_u9_u6_n97 ) );
  AOI22_X1 u2_u9_u6_U33 (.B2( u2_u9_u6_n110 ) , .B1( u2_u9_u6_n111 ) , .A1( u2_u9_u6_n112 ) , .ZN( u2_u9_u6_n115 ) , .A2( u2_u9_u6_n161 ) );
  NAND4_X1 u2_u9_u6_U34 (.A3( u2_u9_u6_n109 ) , .ZN( u2_u9_u6_n112 ) , .A4( u2_u9_u6_n132 ) , .A2( u2_u9_u6_n147 ) , .A1( u2_u9_u6_n166 ) );
  NOR2_X1 u2_u9_u6_U35 (.ZN( u2_u9_u6_n109 ) , .A1( u2_u9_u6_n170 ) , .A2( u2_u9_u6_n173 ) );
  NOR2_X1 u2_u9_u6_U36 (.A2( u2_u9_u6_n126 ) , .ZN( u2_u9_u6_n155 ) , .A1( u2_u9_u6_n160 ) );
  NAND2_X1 u2_u9_u6_U37 (.ZN( u2_u9_u6_n146 ) , .A2( u2_u9_u6_n94 ) , .A1( u2_u9_u6_n99 ) );
  AOI21_X1 u2_u9_u6_U38 (.A( u2_u9_u6_n144 ) , .B2( u2_u9_u6_n145 ) , .B1( u2_u9_u6_n146 ) , .ZN( u2_u9_u6_n150 ) );
  AOI211_X1 u2_u9_u6_U39 (.B( u2_u9_u6_n134 ) , .A( u2_u9_u6_n135 ) , .C1( u2_u9_u6_n136 ) , .ZN( u2_u9_u6_n137 ) , .C2( u2_u9_u6_n151 ) );
  INV_X1 u2_u9_u6_U4 (.A( u2_u9_u6_n142 ) , .ZN( u2_u9_u6_n174 ) );
  NAND4_X1 u2_u9_u6_U40 (.A4( u2_u9_u6_n127 ) , .A3( u2_u9_u6_n128 ) , .A2( u2_u9_u6_n129 ) , .A1( u2_u9_u6_n130 ) , .ZN( u2_u9_u6_n136 ) );
  AOI21_X1 u2_u9_u6_U41 (.B2( u2_u9_u6_n132 ) , .B1( u2_u9_u6_n133 ) , .ZN( u2_u9_u6_n134 ) , .A( u2_u9_u6_n158 ) );
  AOI21_X1 u2_u9_u6_U42 (.B1( u2_u9_u6_n131 ) , .ZN( u2_u9_u6_n135 ) , .A( u2_u9_u6_n144 ) , .B2( u2_u9_u6_n146 ) );
  INV_X1 u2_u9_u6_U43 (.A( u2_u9_u6_n111 ) , .ZN( u2_u9_u6_n158 ) );
  NAND2_X1 u2_u9_u6_U44 (.ZN( u2_u9_u6_n127 ) , .A1( u2_u9_u6_n91 ) , .A2( u2_u9_u6_n92 ) );
  NAND2_X1 u2_u9_u6_U45 (.ZN( u2_u9_u6_n129 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n96 ) );
  INV_X1 u2_u9_u6_U46 (.A( u2_u9_u6_n144 ) , .ZN( u2_u9_u6_n159 ) );
  NAND2_X1 u2_u9_u6_U47 (.ZN( u2_u9_u6_n145 ) , .A2( u2_u9_u6_n97 ) , .A1( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U48 (.ZN( u2_u9_u6_n148 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n94 ) );
  NAND2_X1 u2_u9_u6_U49 (.ZN( u2_u9_u6_n108 ) , .A2( u2_u9_u6_n139 ) , .A1( u2_u9_u6_n144 ) );
  NAND2_X1 u2_u9_u6_U5 (.A2( u2_u9_u6_n143 ) , .ZN( u2_u9_u6_n152 ) , .A1( u2_u9_u6_n166 ) );
  NAND2_X1 u2_u9_u6_U50 (.ZN( u2_u9_u6_n121 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n97 ) );
  NAND2_X1 u2_u9_u6_U51 (.ZN( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n95 ) );
  AND2_X1 u2_u9_u6_U52 (.ZN( u2_u9_u6_n118 ) , .A2( u2_u9_u6_n91 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U53 (.ZN( u2_u9_u6_n147 ) , .A2( u2_u9_u6_n98 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U54 (.ZN( u2_u9_u6_n128 ) , .A1( u2_u9_u6_n94 ) , .A2( u2_u9_u6_n96 ) );
  NAND2_X1 u2_u9_u6_U55 (.ZN( u2_u9_u6_n119 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U56 (.ZN( u2_u9_u6_n123 ) , .A2( u2_u9_u6_n91 ) , .A1( u2_u9_u6_n96 ) );
  NAND2_X1 u2_u9_u6_U57 (.ZN( u2_u9_u6_n100 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U58 (.ZN( u2_u9_u6_n122 ) , .A1( u2_u9_u6_n94 ) , .A2( u2_u9_u6_n97 ) );
  INV_X1 u2_u9_u6_U59 (.A( u2_u9_u6_n139 ) , .ZN( u2_u9_u6_n160 ) );
  AOI22_X1 u2_u9_u6_U6 (.B2( u2_u9_u6_n101 ) , .A1( u2_u9_u6_n102 ) , .ZN( u2_u9_u6_n103 ) , .B1( u2_u9_u6_n160 ) , .A2( u2_u9_u6_n161 ) );
  NAND2_X1 u2_u9_u6_U60 (.ZN( u2_u9_u6_n113 ) , .A1( u2_u9_u6_n96 ) , .A2( u2_u9_u6_n98 ) );
  NOR2_X1 u2_u9_u6_U61 (.A2( u2_u9_X_40 ) , .A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n126 ) );
  NOR2_X1 u2_u9_u6_U62 (.A2( u2_u9_X_39 ) , .A1( u2_u9_X_42 ) , .ZN( u2_u9_u6_n92 ) );
  NOR2_X1 u2_u9_u6_U63 (.A2( u2_u9_X_39 ) , .A1( u2_u9_u6_n156 ) , .ZN( u2_u9_u6_n97 ) );
  NOR2_X1 u2_u9_u6_U64 (.A2( u2_u9_X_38 ) , .A1( u2_u9_u6_n165 ) , .ZN( u2_u9_u6_n95 ) );
  NOR2_X1 u2_u9_u6_U65 (.A2( u2_u9_X_41 ) , .ZN( u2_u9_u6_n111 ) , .A1( u2_u9_u6_n157 ) );
  NOR2_X1 u2_u9_u6_U66 (.A2( u2_u9_X_37 ) , .A1( u2_u9_u6_n162 ) , .ZN( u2_u9_u6_n94 ) );
  NOR2_X1 u2_u9_u6_U67 (.A2( u2_u9_X_37 ) , .A1( u2_u9_X_38 ) , .ZN( u2_u9_u6_n91 ) );
  NAND2_X1 u2_u9_u6_U68 (.A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n144 ) , .A2( u2_u9_u6_n157 ) );
  NAND2_X1 u2_u9_u6_U69 (.A2( u2_u9_X_40 ) , .A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n139 ) );
  NOR2_X1 u2_u9_u6_U7 (.A1( u2_u9_u6_n118 ) , .ZN( u2_u9_u6_n143 ) , .A2( u2_u9_u6_n168 ) );
  AND2_X1 u2_u9_u6_U70 (.A1( u2_u9_X_39 ) , .A2( u2_u9_u6_n156 ) , .ZN( u2_u9_u6_n96 ) );
  AND2_X1 u2_u9_u6_U71 (.A1( u2_u9_X_39 ) , .A2( u2_u9_X_42 ) , .ZN( u2_u9_u6_n99 ) );
  INV_X1 u2_u9_u6_U72 (.A( u2_u9_X_40 ) , .ZN( u2_u9_u6_n157 ) );
  INV_X1 u2_u9_u6_U73 (.A( u2_u9_X_37 ) , .ZN( u2_u9_u6_n165 ) );
  INV_X1 u2_u9_u6_U74 (.A( u2_u9_X_38 ) , .ZN( u2_u9_u6_n162 ) );
  INV_X1 u2_u9_u6_U75 (.A( u2_u9_X_42 ) , .ZN( u2_u9_u6_n156 ) );
  NAND4_X1 u2_u9_u6_U76 (.ZN( u2_out9_32 ) , .A4( u2_u9_u6_n103 ) , .A3( u2_u9_u6_n104 ) , .A2( u2_u9_u6_n105 ) , .A1( u2_u9_u6_n106 ) );
  AOI22_X1 u2_u9_u6_U77 (.ZN( u2_u9_u6_n105 ) , .A2( u2_u9_u6_n108 ) , .A1( u2_u9_u6_n118 ) , .B2( u2_u9_u6_n126 ) , .B1( u2_u9_u6_n171 ) );
  AOI22_X1 u2_u9_u6_U78 (.ZN( u2_u9_u6_n104 ) , .A1( u2_u9_u6_n111 ) , .B1( u2_u9_u6_n124 ) , .B2( u2_u9_u6_n151 ) , .A2( u2_u9_u6_n93 ) );
  NAND4_X1 u2_u9_u6_U79 (.ZN( u2_out9_12 ) , .A4( u2_u9_u6_n114 ) , .A3( u2_u9_u6_n115 ) , .A2( u2_u9_u6_n116 ) , .A1( u2_u9_u6_n117 ) );
  OAI21_X1 u2_u9_u6_U8 (.A( u2_u9_u6_n159 ) , .B1( u2_u9_u6_n169 ) , .B2( u2_u9_u6_n173 ) , .ZN( u2_u9_u6_n90 ) );
  OAI22_X1 u2_u9_u6_U80 (.B2( u2_u9_u6_n111 ) , .ZN( u2_u9_u6_n116 ) , .B1( u2_u9_u6_n126 ) , .A2( u2_u9_u6_n164 ) , .A1( u2_u9_u6_n167 ) );
  OAI21_X1 u2_u9_u6_U81 (.A( u2_u9_u6_n108 ) , .ZN( u2_u9_u6_n117 ) , .B2( u2_u9_u6_n141 ) , .B1( u2_u9_u6_n163 ) );
  OAI211_X1 u2_u9_u6_U82 (.ZN( u2_out9_7 ) , .B( u2_u9_u6_n153 ) , .C2( u2_u9_u6_n154 ) , .C1( u2_u9_u6_n155 ) , .A( u2_u9_u6_n174 ) );
  NOR3_X1 u2_u9_u6_U83 (.A1( u2_u9_u6_n141 ) , .ZN( u2_u9_u6_n154 ) , .A3( u2_u9_u6_n164 ) , .A2( u2_u9_u6_n171 ) );
  AOI211_X1 u2_u9_u6_U84 (.B( u2_u9_u6_n149 ) , .A( u2_u9_u6_n150 ) , .C2( u2_u9_u6_n151 ) , .C1( u2_u9_u6_n152 ) , .ZN( u2_u9_u6_n153 ) );
  OAI211_X1 u2_u9_u6_U85 (.ZN( u2_out9_22 ) , .B( u2_u9_u6_n137 ) , .A( u2_u9_u6_n138 ) , .C2( u2_u9_u6_n139 ) , .C1( u2_u9_u6_n140 ) );
  AOI22_X1 u2_u9_u6_U86 (.B1( u2_u9_u6_n124 ) , .A2( u2_u9_u6_n125 ) , .A1( u2_u9_u6_n126 ) , .ZN( u2_u9_u6_n138 ) , .B2( u2_u9_u6_n161 ) );
  AND4_X1 u2_u9_u6_U87 (.A3( u2_u9_u6_n119 ) , .A1( u2_u9_u6_n120 ) , .A4( u2_u9_u6_n129 ) , .ZN( u2_u9_u6_n140 ) , .A2( u2_u9_u6_n143 ) );
  NAND3_X1 u2_u9_u6_U88 (.A2( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n125 ) , .A1( u2_u9_u6_n130 ) , .A3( u2_u9_u6_n131 ) );
  NAND3_X1 u2_u9_u6_U89 (.A3( u2_u9_u6_n133 ) , .ZN( u2_u9_u6_n141 ) , .A1( u2_u9_u6_n145 ) , .A2( u2_u9_u6_n148 ) );
  INV_X1 u2_u9_u6_U9 (.ZN( u2_u9_u6_n172 ) , .A( u2_u9_u6_n88 ) );
  NAND3_X1 u2_u9_u6_U90 (.ZN( u2_u9_u6_n101 ) , .A3( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n121 ) , .A1( u2_u9_u6_n127 ) );
  NAND3_X1 u2_u9_u6_U91 (.ZN( u2_u9_u6_n102 ) , .A3( u2_u9_u6_n130 ) , .A2( u2_u9_u6_n145 ) , .A1( u2_u9_u6_n166 ) );
  NAND3_X1 u2_u9_u6_U92 (.A3( u2_u9_u6_n113 ) , .A1( u2_u9_u6_n119 ) , .A2( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n93 ) );
  NAND3_X1 u2_u9_u6_U93 (.ZN( u2_u9_u6_n142 ) , .A2( u2_u9_u6_n172 ) , .A3( u2_u9_u6_n89 ) , .A1( u2_u9_u6_n90 ) );
  INV_X1 u2_uk_U10 (.A( u2_uk_n188 ) , .ZN( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U1005 (.ZN( u2_K10_21 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1630 ) , .A( u2_uk_n252 ) );
  NAND2_X1 u2_uk_U1006 (.A1( u2_uk_K_r8_19 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n252 ) );
  OAI21_X1 u2_uk_U1009 (.ZN( u2_K9_39 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1135 ) , .B2( u2_uk_n1571 ) );
  NAND2_X1 u2_uk_U1010 (.A1( u2_uk_K_r7_31 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n1135 ) );
  OAI21_X1 u2_uk_U1013 (.ZN( u2_K9_44 ) , .A( u2_uk_n1138 ) , .B2( u2_uk_n1585 ) , .B1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U1014 (.A1( u2_uk_K_r7_0 ) , .ZN( u2_uk_n1138 ) , .A2( u2_uk_n155 ) );
  OAI21_X1 u2_uk_U1019 (.ZN( u2_K12_36 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1698 ) , .A( u2_uk_n472 ) );
  OAI21_X1 u2_uk_U1021 (.ZN( u2_K6_41 ) , .A( u2_uk_n1069 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1445 ) );
  OAI21_X1 u2_uk_U1023 (.ZN( u2_K8_28 ) , .A( u2_uk_n1103 ) , .B2( u2_uk_n1532 ) , .B1( u2_uk_n27 ) );
  NAND2_X1 u2_uk_U1024 (.A1( u2_uk_K_r6_51 ) , .ZN( u2_uk_n1103 ) , .A2( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U1029 (.ZN( u2_K12_40 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1699 ) , .A( u2_uk_n501 ) );
  NAND2_X1 u2_uk_U1030 (.A1( u2_uk_K_r10_49 ) , .A2( u2_uk_n102 ) , .ZN( u2_uk_n501 ) );
  OAI21_X1 u2_uk_U1031 (.ZN( u2_K15_14 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1821 ) , .A( u2_uk_n936 ) );
  NAND2_X1 u2_uk_U1032 (.A1( u2_uk_K_r13_32 ) , .A2( u2_uk_n83 ) , .ZN( u2_uk_n936 ) );
  OAI21_X1 u2_uk_U1037 (.ZN( u2_K5_42 ) , .A( u2_uk_n1052 ) , .B2( u2_uk_n1382 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U1038 (.A1( u2_uk_K_r3_9 ) , .ZN( u2_uk_n1052 ) , .A2( u2_uk_n60 ) );
  NAND2_X1 u2_uk_U1040 (.A1( u2_uk_K_r2_50 ) , .A2( u2_uk_n102 ) , .ZN( u2_uk_n1034 ) );
  INV_X1 u2_uk_U1043 (.A( u2_key_r_9 ) , .ZN( u2_uk_n1149 ) );
  INV_X1 u2_uk_U1044 (.A( u2_key_r_7 ) , .ZN( u2_uk_n1147 ) );
  INV_X1 u2_uk_U1047 (.A( u2_key_r_23 ) , .ZN( u2_uk_n1158 ) );
  INV_X1 u2_uk_U1049 (.A( u2_key_r_30 ) , .ZN( u2_uk_n1165 ) );
  INV_X1 u2_uk_U1055 (.A( u2_key_r_37 ) , .ZN( u2_uk_n1171 ) );
  INV_X1 u2_uk_U1056 (.A( u2_key_r_52 ) , .ZN( u2_uk_n1183 ) );
  INV_X1 u2_uk_U1057 (.A( u2_key_r_0 ) , .ZN( u2_uk_n1142 ) );
  INV_X1 u2_uk_U1058 (.A( u2_key_r_16 ) , .ZN( u2_uk_n1152 ) );
  OAI22_X1 u2_uk_U106 (.ZN( u2_K10_41 ) , .A2( u2_uk_n1594 ) , .B2( u2_uk_n1622 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n231 ) );
  INV_X1 u2_uk_U1061 (.A( u2_key_r_2 ) , .ZN( u2_uk_n1144 ) );
  OAI21_X1 u2_uk_U1066 (.ZN( u2_K13_28 ) , .B2( u2_uk_n1753 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n662 ) );
  NAND2_X1 u2_uk_U1067 (.A1( u2_uk_K_r11_21 ) , .A2( u2_uk_n238 ) , .ZN( u2_uk_n662 ) );
  OAI21_X1 u2_uk_U1070 (.ZN( u2_K16_14 ) , .B2( u2_uk_n1205 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n951 ) );
  NAND2_X1 u2_uk_U1071 (.A1( u2_uk_K_r14_18 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n951 ) );
  OAI21_X1 u2_uk_U1078 (.ZN( u2_K5_39 ) , .A( u2_uk_n1051 ) , .B2( u2_uk_n1376 ) , .B1( u2_uk_n162 ) );
  NAND2_X1 u2_uk_U1079 (.A1( u2_uk_K_r3_16 ) , .ZN( u2_uk_n1051 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1081 (.ZN( u2_K13_10 ) , .A( u2_uk_n524 ) );
  INV_X1 u2_uk_U1082 (.ZN( u2_K2_10 ) , .A( u2_uk_n991 ) );
  AOI22_X1 u2_uk_U1083 (.B2( u2_uk_K_r0_34 ) , .A2( u2_uk_K_r0_55 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n147 ) , .ZN( u2_uk_n991 ) );
  INV_X1 u2_uk_U1092 (.ZN( u2_K1_41 ) , .A( u2_uk_n985 ) );
  AOI22_X1 u2_uk_U1093 (.B2( u2_key_r_35 ) , .A2( u2_key_r_42 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) , .ZN( u2_uk_n985 ) );
  INV_X1 u2_uk_U11 (.A( u2_uk_n163 ) , .ZN( u2_uk_n60 ) );
  INV_X1 u2_uk_U1104 (.ZN( u2_K4_3 ) , .A( u2_uk_n1035 ) );
  INV_X1 u2_uk_U1106 (.ZN( u2_K12_23 ) , .A( u2_uk_n454 ) );
  AOI22_X1 u2_uk_U1107 (.B2( u2_uk_K_r10_32 ) , .A2( u2_uk_K_r10_41 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n454 ) );
  INV_X1 u2_uk_U1108 (.ZN( u2_K2_7 ) , .A( u2_uk_n1004 ) );
  AOI22_X1 u2_uk_U1109 (.B2( u2_uk_K_r0_13 ) , .A2( u2_uk_K_r0_34 ) , .ZN( u2_uk_n1004 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U1110 (.ZN( u2_K12_32 ) , .A( u2_uk_n467 ) );
  INV_X1 u2_uk_U1112 (.ZN( u2_K9_20 ) , .A( u2_uk_n1126 ) );
  AOI22_X1 u2_uk_U1113 (.B2( u2_uk_K_r7_32 ) , .A2( u2_uk_K_r7_39 ) , .ZN( u2_uk_n1126 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1118 (.ZN( u2_K1_32 ) , .A( u2_uk_n980 ) );
  AOI22_X1 u2_uk_U1119 (.B2( u2_key_r_22 ) , .A2( u2_key_r_29 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n980 ) );
  INV_X1 u2_uk_U1120 (.ZN( u2_K7_32 ) , .A( u2_uk_n1088 ) );
  AOI22_X1 u2_uk_U1121 (.B2( u2_uk_K_r5_0 ) , .A2( u2_uk_K_r5_51 ) , .ZN( u2_uk_n1088 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n231 ) );
  INV_X1 u2_uk_U1124 (.ZN( u2_K4_4 ) , .A( u2_uk_n1037 ) );
  AOI22_X1 u2_uk_U1125 (.B2( u2_uk_K_r2_13 ) , .A2( u2_uk_K_r2_18 ) , .ZN( u2_uk_n1037 ) , .B1( u2_uk_n147 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U1126 (.ZN( u2_K5_35 ) , .A( u2_uk_n1049 ) );
  INV_X1 u2_uk_U1128 (.ZN( u2_K6_4 ) , .A( u2_uk_n1071 ) );
  AOI22_X1 u2_uk_U1129 (.B2( u2_uk_K_r4_41 ) , .A2( u2_uk_K_r4_47 ) , .ZN( u2_uk_n1071 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n60 ) );
  INV_X1 u2_uk_U113 (.ZN( u2_K11_47 ) , .A( u2_uk_n386 ) );
  INV_X1 u2_uk_U1130 (.ZN( u2_K4_10 ) , .A( u2_uk_n1020 ) );
  AOI22_X1 u2_uk_U1131 (.B2( u2_uk_K_r2_26 ) , .A2( u2_uk_K_r2_6 ) , .ZN( u2_uk_n1020 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n60 ) );
  INV_X1 u2_uk_U1134 (.ZN( u2_K13_12 ) , .A( u2_uk_n551 ) );
  AOI22_X1 u2_uk_U114 (.B2( u2_uk_K_r9_15 ) , .A2( u2_uk_K_r9_23 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n223 ) , .ZN( u2_uk_n386 ) );
  INV_X1 u2_uk_U1143 (.ZN( u2_K15_43 ) , .A( u2_uk_n944 ) );
  INV_X1 u2_uk_U1146 (.ZN( u2_K13_2 ) , .A( u2_uk_n665 ) );
  AOI22_X1 u2_uk_U1147 (.B2( u2_uk_K_r11_26 ) , .A2( u2_uk_K_r11_6 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n524 ) );
  INV_X1 u2_uk_U1149 (.ZN( u2_K13_6 ) , .A( u2_uk_n681 ) );
  INV_X1 u2_uk_U1153 (.ZN( u2_K9_2 ) , .A( u2_uk_n1130 ) );
  AOI22_X1 u2_uk_U1154 (.B2( u2_uk_K_r4_17 ) , .A2( u2_uk_K_r4_55 ) , .ZN( u2_uk_n1066 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1155 (.ZN( u2_K6_2 ) , .A( u2_uk_n1066 ) );
  INV_X1 u2_uk_U1157 (.ZN( u2_K4_2 ) , .A( u2_uk_n1031 ) );
  OAI21_X1 u2_uk_U118 (.ZN( u2_K6_47 ) , .A( u2_uk_n1070 ) , .B2( u2_uk_n1419 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U121 (.ZN( u2_K4_47 ) , .B2( u2_uk_n1350 ) , .A2( u2_uk_n1359 ) , .A1( u2_uk_n187 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U128 (.ZN( u2_K13_15 ) , .A( u2_uk_n586 ) );
  INV_X1 u2_uk_U134 (.ZN( u2_K13_19 ) , .A( u2_uk_n601 ) );
  AOI22_X1 u2_uk_U135 (.B2( u2_uk_K_r11_19 ) , .A2( u2_uk_K_r11_39 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n601 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U136 (.ZN( u2_K11_15 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1646 ) , .A2( u2_uk_n1661 ) , .B1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U139 (.ZN( u2_K2_15 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1261 ) , .A( u2_uk_n994 ) );
  OAI22_X1 u2_uk_U142 (.ZN( u2_K16_15 ) , .B2( u2_uk_n1206 ) , .A2( u2_uk_n1213 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U144 (.ZN( u2_K15_15 ) , .B2( u2_uk_n1843 ) , .B1( u2_uk_n188 ) , .A( u2_uk_n937 ) );
  NAND2_X1 u2_uk_U145 (.A1( u2_uk_K_r13_19 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n937 ) );
  INV_X1 u2_uk_U151 (.ZN( u2_K9_19 ) , .A( u2_uk_n1124 ) );
  AOI22_X1 u2_uk_U152 (.B1( u2_uk_K_r7_13 ) , .A2( u2_uk_K_r7_20 ) , .B2( u2_uk_n10 ) , .ZN( u2_uk_n1124 ) , .A1( u2_uk_n162 ) );
  INV_X1 u2_uk_U156 (.ZN( u2_K2_19 ) , .A( u2_uk_n995 ) );
  AOI22_X1 u2_uk_U157 (.B2( u2_uk_K_r0_11 ) , .A2( u2_uk_K_r0_47 ) , .A1( u2_uk_n128 ) , .B1( u2_uk_n231 ) , .ZN( u2_uk_n995 ) );
  OAI22_X1 u2_uk_U158 (.ZN( u2_K16_19 ) , .B2( u2_uk_n1190 ) , .A2( u2_uk_n1228 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U16 (.A( u2_uk_n146 ) , .ZN( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U160 (.ZN( u2_K10_19 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1603 ) , .A2( u2_uk_n1613 ) , .B1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U161 (.ZN( u2_K5_30 ) , .B2( u2_uk_n1378 ) , .A2( u2_uk_n1395 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U164 (.ZN( u2_K12_30 ) , .A( u2_uk_n456 ) );
  INV_X1 u2_uk_U17 (.ZN( u2_uk_n109 ) , .A( u2_uk_n146 ) );
  OAI21_X1 u2_uk_U171 (.ZN( u2_K8_30 ) , .A( u2_uk_n1106 ) , .B2( u2_uk_n1525 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U172 (.A1( u2_uk_K_r6_29 ) , .ZN( u2_uk_n1106 ) , .A2( u2_uk_n191 ) );
  INV_X1 u2_uk_U177 (.ZN( u2_K11_14 ) , .A( u2_uk_n319 ) );
  OAI21_X1 u2_uk_U179 (.ZN( u2_K10_24 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1599 ) , .A( u2_uk_n277 ) );
  INV_X1 u2_uk_U18 (.ZN( u2_uk_n110 ) , .A( u2_uk_n209 ) );
  NAND2_X1 u2_uk_U180 (.A1( u2_uk_K_r8_40 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n277 ) );
  OAI21_X1 u2_uk_U181 (.ZN( u2_K9_14 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1121 ) , .B2( u2_uk_n1574 ) );
  INV_X1 u2_uk_U184 (.ZN( u2_K2_14 ) , .A( u2_uk_n993 ) );
  AOI22_X1 u2_uk_U185 (.B2( u2_uk_K_r0_11 ) , .A2( u2_uk_K_r0_32 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n993 ) );
  OAI21_X1 u2_uk_U190 (.ZN( u2_K13_30 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1746 ) , .A( u2_uk_n671 ) );
  NAND2_X1 u2_uk_U191 (.A1( u2_uk_K_r11_28 ) , .A2( u2_uk_n17 ) , .ZN( u2_uk_n671 ) );
  OAI22_X1 u2_uk_U199 (.ZN( u2_K15_24 ) , .A2( u2_uk_n1816 ) , .B2( u2_uk_n1834 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U20 (.ZN( u2_uk_n102 ) , .A( u2_uk_n146 ) );
  OAI21_X1 u2_uk_U200 (.ZN( u2_K1_30 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1183 ) , .A( u2_uk_n979 ) );
  OAI21_X1 u2_uk_U202 (.ZN( u2_K9_30 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1131 ) , .B2( u2_uk_n1570 ) );
  INV_X1 u2_uk_U21 (.ZN( u2_uk_n128 ) , .A( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U211 (.ZN( u2_K1_31 ) , .A2( u2_uk_n1147 ) , .B2( u2_uk_n1151 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U212 (.A( u2_key_r_14 ) , .ZN( u2_uk_n1151 ) );
  OAI21_X1 u2_uk_U215 (.ZN( u2_K12_31 ) , .B2( u2_uk_n1685 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n460 ) );
  NAND2_X1 u2_uk_U216 (.A1( u2_uk_K_r10_44 ) , .A2( u2_uk_n217 ) , .ZN( u2_uk_n460 ) );
  INV_X1 u2_uk_U217 (.ZN( u2_K11_31 ) , .A( u2_uk_n373 ) );
  INV_X1 u2_uk_U220 (.ZN( u2_K11_39 ) , .A( u2_uk_n379 ) );
  INV_X1 u2_uk_U222 (.ZN( u2_K10_39 ) , .A( u2_uk_n305 ) );
  AOI22_X1 u2_uk_U223 (.B2( u2_uk_K_r8_44 ) , .A2( u2_uk_K_r8_52 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n305 ) );
  OAI21_X1 u2_uk_U225 (.ZN( u2_K10_31 ) , .B2( u2_uk_n1615 ) , .B1( u2_uk_n164 ) , .A( u2_uk_n291 ) );
  NAND2_X1 u2_uk_U226 (.A1( u2_uk_K_r8_16 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n291 ) );
  OAI22_X1 u2_uk_U227 (.ZN( u2_K6_31 ) , .B2( u2_uk_n1425 ) , .A2( u2_uk_n1430 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n60 ) );
  BUF_X1 u2_uk_U23 (.Z( u2_uk_n155 ) , .A( u2_uk_n214 ) );
  OAI21_X1 u2_uk_U232 (.ZN( u2_K1_39 ) , .B2( u2_uk_n1157 ) , .B1( u2_uk_n63 ) , .A( u2_uk_n984 ) );
  INV_X1 u2_uk_U234 (.A( u2_key_r_22 ) , .ZN( u2_uk_n1157 ) );
  BUF_X1 u2_uk_U24 (.Z( u2_uk_n145 ) , .A( u2_uk_n222 ) );
  OAI21_X1 u2_uk_U240 (.ZN( u2_K12_39 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1690 ) , .A( u2_uk_n496 ) );
  NAND2_X1 u2_uk_U241 (.A1( u2_uk_K_r10_16 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n496 ) );
  INV_X1 u2_uk_U247 (.ZN( u2_K1_48 ) , .A( u2_uk_n989 ) );
  AOI22_X1 u2_uk_U248 (.B2( u2_key_r_21 ) , .A2( u2_key_r_28 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n217 ) , .ZN( u2_uk_n989 ) );
  OAI22_X1 u2_uk_U249 (.ZN( u2_K15_44 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1836 ) , .A2( u2_uk_n1854 ) , .A1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U250 (.ZN( u2_K15_48 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1824 ) , .A( u2_uk_n945 ) );
  INV_X1 u2_uk_U256 (.ZN( u2_K12_44 ) , .A( u2_uk_n504 ) );
  OAI22_X1 u2_uk_U258 (.ZN( u2_K12_48 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1691 ) , .A2( u2_uk_n1700 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U259 (.ZN( u2_K11_44 ) , .A1( u2_uk_n142 ) , .B2( u2_uk_n1653 ) , .A2( u2_uk_n1673 ) , .B1( u2_uk_n63 ) );
  BUF_X1 u2_uk_U26 (.Z( u2_uk_n148 ) , .A( u2_uk_n217 ) );
  INV_X1 u2_uk_U262 (.ZN( u2_K9_48 ) , .A( u2_uk_n1140 ) );
  OAI22_X1 u2_uk_U269 (.ZN( u2_K6_44 ) , .B2( u2_uk_n1428 ) , .A2( u2_uk_n1446 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U270 (.ZN( u2_K6_48 ) , .B2( u2_uk_n1433 ) , .A2( u2_uk_n1440 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U271 (.ZN( u2_K4_44 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1320 ) , .A2( u2_uk_n1337 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U280 (.ZN( u2_K6_6 ) , .B2( u2_uk_n1444 ) , .A2( u2_uk_n1448 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U281 (.ZN( u2_K6_8 ) , .A( u2_uk_n1073 ) , .B2( u2_uk_n1416 ) , .B1( u2_uk_n31 ) );
  BUF_X1 u2_uk_U29 (.Z( u2_uk_n147 ) , .A( u2_uk_n217 ) );
  INV_X1 u2_uk_U292 (.ZN( u2_K4_8 ) , .A( u2_uk_n1040 ) );
  OAI21_X1 u2_uk_U295 (.ZN( u2_K2_8 ) , .A( u2_uk_n1005 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1240 ) );
  NAND2_X1 u2_uk_U296 (.A1( u2_uk_K_r0_17 ) , .ZN( u2_uk_n1005 ) , .A2( u2_uk_n93 ) );
  INV_X1 u2_uk_U298 (.ZN( u2_K1_26 ) , .A( u2_uk_n976 ) );
  AOI22_X1 u2_uk_U299 (.B2( u2_key_r_31 ) , .A2( u2_key_r_51 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n976 ) );
  INV_X1 u2_uk_U301 (.ZN( u2_K9_26 ) , .A( u2_uk_n1128 ) );
  BUF_X1 u2_uk_U31 (.Z( u2_uk_n163 ) , .A( u2_uk_n209 ) );
  BUF_X1 u2_uk_U32 (.Z( u2_uk_n162 ) , .A( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U320 (.ZN( u2_K3_26 ) , .B2( u2_uk_n1299 ) , .A2( u2_uk_n1315 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U322 (.ZN( u2_K15_46 ) , .B1( u2_uk_n17 ) , .A2( u2_uk_n1818 ) , .B2( u2_uk_n1845 ) , .A1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U325 (.ZN( u2_K4_46 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1330 ) , .A2( u2_uk_n1344 ) , .B1( u2_uk_n155 ) );
  INV_X1 u2_uk_U334 (.ZN( u2_K11_46 ) , .A( u2_uk_n385 ) );
  OAI21_X1 u2_uk_U336 (.ZN( u2_K9_46 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1139 ) , .B2( u2_uk_n1577 ) );
  NAND2_X1 u2_uk_U337 (.A1( u2_uk_K_r7_37 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n1139 ) );
  INV_X1 u2_uk_U350 (.ZN( u2_K10_40 ) , .A( u2_uk_n306 ) );
  AOI22_X1 u2_uk_U351 (.A2( u2_uk_K_r8_2 ) , .B2( u2_uk_K_r8_22 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n306 ) );
  OAI22_X1 u2_uk_U357 (.ZN( u2_K11_40 ) , .A1( u2_uk_n161 ) , .A2( u2_uk_n1634 ) , .B2( u2_uk_n1642 ) , .B1( u2_uk_n63 ) );
  BUF_X1 u2_uk_U36 (.Z( u2_uk_n188 ) , .A( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U360 (.ZN( u2_K4_40 ) , .B2( u2_uk_n1342 ) , .A2( u2_uk_n1352 ) , .A1( u2_uk_n146 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U373 (.ZN( u2_K3_28 ) , .B2( u2_uk_n1298 ) , .A2( u2_uk_n1303 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U374 (.ZN( u2_K5_33 ) , .A( u2_uk_n1048 ) , .B2( u2_uk_n1401 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U375 (.A1( u2_uk_K_r3_14 ) , .ZN( u2_uk_n1048 ) , .A2( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U377 (.ZN( u2_K12_28 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1680 ) , .A2( u2_uk_n1684 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U378 (.ZN( u2_K10_28 ) , .B2( u2_uk_n1610 ) , .A2( u2_uk_n1617 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U388 (.ZN( u2_K4_1 ) , .A( u2_uk_n1023 ) , .B2( u2_uk_n1323 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U389 (.A1( u2_uk_K_r2_25 ) , .ZN( u2_uk_n1023 ) , .A2( u2_uk_n214 ) );
  BUF_X1 u2_uk_U39 (.Z( u2_uk_n214 ) , .A( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U395 (.ZN( u2_K13_16 ) , .B2( u2_uk_n1731 ) , .A2( u2_uk_n1736 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U398 (.ZN( u2_K9_16 ) , .B2( u2_uk_n1548 ) , .A2( u2_uk_n1555 ) , .B1( u2_uk_n220 ) , .A1( u2_uk_n99 ) );
  BUF_X1 u2_uk_U40 (.Z( u2_uk_n209 ) , .A( u2_uk_n231 ) );
  BUF_X1 u2_uk_U41 (.Z( u2_uk_n203 ) , .A( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U411 (.ZN( u2_K13_9 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1731 ) , .A2( u2_uk_n1743 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U415 (.ZN( u2_K4_9 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1329 ) , .A2( u2_uk_n1339 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U416 (.ZN( u2_K10_37 ) , .A( u2_uk_n299 ) );
  INV_X1 u2_uk_U422 (.ZN( u2_K9_9 ) , .A( u2_uk_n1141 ) );
  INV_X1 u2_uk_U424 (.ZN( u2_K6_9 ) , .A( u2_uk_n1074 ) );
  OAI22_X1 u2_uk_U430 (.ZN( u2_K2_9 ) , .A2( u2_uk_n1232 ) , .B2( u2_uk_n1261 ) , .B1( u2_uk_n145 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U434 (.ZN( u2_K16_16 ) , .B2( u2_uk_n1207 ) , .A2( u2_uk_n1214 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U438 (.ZN( u2_K4_37 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1331 ) , .A2( u2_uk_n1345 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U446 (.ZN( u2_K10_33 ) , .A( u2_uk_n294 ) );
  AOI22_X1 u2_uk_U447 (.B2( u2_uk_K_r8_22 ) , .A2( u2_uk_K_r8_42 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n294 ) );
  INV_X1 u2_uk_U448 (.ZN( u2_K1_33 ) , .A( u2_uk_n981 ) );
  AOI22_X1 u2_uk_U449 (.B2( u2_key_r_44 ) , .A2( u2_key_r_51 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n981 ) );
  BUF_X1 u2_uk_U45 (.A( u2_uk_n203 ) , .Z( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U450 (.ZN( u2_K12_33 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1718 ) , .A( u2_uk_n468 ) );
  OAI22_X1 u2_uk_U454 (.ZN( u2_K13_33 ) , .B2( u2_uk_n1723 ) , .A2( u2_uk_n1728 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U455 (.ZN( u2_K11_33 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1653 ) , .A2( u2_uk_n1659 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U456 (.ZN( u2_K8_33 ) , .B2( u2_uk_n1498 ) , .A2( u2_uk_n1503 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U457 (.ZN( u2_K6_33 ) , .B2( u2_uk_n1428 ) , .A2( u2_uk_n1433 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n60 ) );
  BUF_X1 u2_uk_U46 (.A( u2_uk_n155 ) , .Z( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U464 (.ZN( u2_K11_37 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1664 ) , .A( u2_uk_n377 ) );
  OAI21_X1 u2_uk_U466 (.ZN( u2_K9_37 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1134 ) , .B2( u2_uk_n1551 ) );
  OAI21_X1 u2_uk_U468 (.ZN( u2_K6_37 ) , .A( u2_uk_n1068 ) , .B2( u2_uk_n1438 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U469 (.A1( u2_uk_K_r4_38 ) , .ZN( u2_uk_n1068 ) , .A2( u2_uk_n217 ) );
  BUF_X1 u2_uk_U47 (.Z( u2_uk_n223 ) , .A( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U470 (.ZN( u2_K5_37 ) , .B2( u2_uk_n1365 ) , .A2( u2_uk_n1403 ) , .B1( u2_uk_n147 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U472 (.ZN( u2_K1_29 ) , .B2( u2_uk_n1152 ) , .A2( u2_uk_n1158 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U477 (.ZN( u2_K13_29 ) , .B2( u2_uk_n1742 ) , .A2( u2_uk_n1745 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  BUF_X1 u2_uk_U48 (.Z( u2_uk_n191 ) , .A( u2_uk_n217 ) );
  OAI21_X1 u2_uk_U485 (.ZN( u2_K3_29 ) , .A( u2_uk_n1010 ) , .B2( u2_uk_n1313 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U486 (.A1( u2_uk_K_r1_44 ) , .ZN( u2_uk_n1010 ) , .A2( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U489 (.ZN( u2_K10_29 ) , .B2( u2_uk_n1597 ) , .A2( u2_uk_n1625 ) , .B1( u2_uk_n202 ) , .A1( u2_uk_n92 ) );
  BUF_X1 u2_uk_U49 (.Z( u2_uk_n231 ) , .A( u2_uk_n238 ) );
  INV_X1 u2_uk_U491 (.ZN( u2_K8_29 ) , .A( u2_uk_n1104 ) );
  OAI22_X1 u2_uk_U494 (.ZN( u2_K5_29 ) , .B2( u2_uk_n1377 ) , .A2( u2_uk_n1396 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n92 ) );
  BUF_X1 u2_uk_U50 (.Z( u2_uk_n230 ) , .A( u2_uk_n238 ) );
  OAI21_X1 u2_uk_U505 (.ZN( u2_K9_12 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1119 ) , .B2( u2_uk_n1543 ) );
  OAI21_X1 u2_uk_U509 (.ZN( u2_K13_17 ) , .B2( u2_uk_n1743 ) , .A( u2_uk_n587 ) , .B1( u2_uk_n60 ) );
  NAND2_X1 u2_uk_U510 (.A1( u2_uk_K_r11_27 ) , .ZN( u2_uk_n587 ) , .A2( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U512 (.ZN( u2_K9_17 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1122 ) , .B2( u2_uk_n1568 ) );
  NAND2_X1 u2_uk_U513 (.A1( u2_uk_K_r7_26 ) , .ZN( u2_uk_n1122 ) , .A2( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U529 (.ZN( u2_K4_12 ) , .A1( u2_uk_n109 ) , .B2( u2_uk_n1341 ) , .A2( u2_uk_n1361 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U531 (.ZN( u2_K2_12 ) , .A2( u2_uk_n1233 ) , .B2( u2_uk_n1248 ) , .A1( u2_uk_n141 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U533 (.ZN( u2_K1_36 ) , .B2( u2_uk_n1158 ) , .A2( u2_uk_n1165 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U534 (.ZN( u2_K16_12 ) , .B2( u2_uk_n1198 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n949 ) );
  NAND2_X1 u2_uk_U535 (.A1( u2_uk_K_r14_12 ) , .A2( u2_uk_n145 ) , .ZN( u2_uk_n949 ) );
  OAI21_X1 u2_uk_U536 (.ZN( u2_K16_17 ) , .B2( u2_uk_n1197 ) , .B1( u2_uk_n188 ) , .A( u2_uk_n952 ) );
  NAND2_X1 u2_uk_U537 (.A1( u2_uk_K_r14_10 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n952 ) );
  OAI22_X1 u2_uk_U539 (.ZN( u2_K15_17 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1814 ) , .B2( u2_uk_n1832 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U54 (.ZN( u2_K11_34 ) , .A( u2_uk_n375 ) );
  INV_X1 u2_uk_U544 (.ZN( u2_K11_17 ) , .A( u2_uk_n335 ) );
  AOI22_X1 u2_uk_U545 (.B2( u2_uk_K_r9_4 ) , .A2( u2_uk_K_r9_55 ) , .A1( u2_uk_n109 ) , .B1( u2_uk_n231 ) , .ZN( u2_uk_n335 ) );
  AOI22_X1 u2_uk_U55 (.B2( u2_uk_K_r9_45 ) , .A2( u2_uk_K_r9_49 ) , .B1( u2_uk_n10 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n375 ) );
  OAI22_X1 u2_uk_U550 (.ZN( u2_K13_36 ) , .B2( u2_uk_n1747 ) , .A2( u2_uk_n1753 ) , .B1( u2_uk_n202 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U553 (.ZN( u2_K1_38 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1165 ) , .A2( u2_uk_n1171 ) , .B1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U554 (.ZN( u2_K12_38 ) , .A1( u2_uk_n10 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1678 ) , .A2( u2_uk_n1705 ) );
  INV_X1 u2_uk_U557 (.ZN( u2_K7_36 ) , .A( u2_uk_n1091 ) );
  AOI22_X1 u2_uk_U558 (.B2( u2_uk_K_r5_1 ) , .A2( u2_uk_K_r5_21 ) , .ZN( u2_uk_n1091 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n202 ) );
  INV_X1 u2_uk_U559 (.ZN( u2_K11_36 ) , .A( u2_uk_n376 ) );
  INV_X1 u2_uk_U56 (.ZN( u2_K8_34 ) , .A( u2_uk_n1107 ) );
  INV_X1 u2_uk_U561 (.ZN( u2_K5_36 ) , .A( u2_uk_n1050 ) );
  AOI22_X1 u2_uk_U562 (.B2( u2_uk_K_r3_29 ) , .A2( u2_uk_K_r3_52 ) , .ZN( u2_uk_n1050 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n191 ) );
  INV_X1 u2_uk_U566 (.ZN( u2_K10_38 ) , .A( u2_uk_n301 ) );
  AOI22_X1 u2_uk_U567 (.B2( u2_uk_K_r8_28 ) , .A2( u2_uk_K_r8_8 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n301 ) );
  OAI22_X1 u2_uk_U568 (.ZN( u2_K8_36 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1524 ) , .A2( u2_uk_n1530 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U569 (.ZN( u2_K6_38 ) , .B2( u2_uk_n1418 ) , .A2( u2_uk_n1425 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U578 (.ZN( u2_K16_10 ) , .B2( u2_uk_n1219 ) , .A2( u2_uk_n1222 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n217 ) );
  INV_X1 u2_uk_U579 (.ZN( u2_K9_10 ) , .A( u2_uk_n1117 ) );
  INV_X1 u2_uk_U58 (.ZN( u2_K7_34 ) , .A( u2_uk_n1089 ) );
  AOI22_X1 u2_uk_U580 (.B2( u2_uk_K_r7_25 ) , .A2( u2_uk_K_r7_32 ) , .B1( u2_uk_n110 ) , .ZN( u2_uk_n1117 ) , .A1( u2_uk_n163 ) );
  INV_X1 u2_uk_U582 (.ZN( u2_K6_10 ) , .A( u2_uk_n1058 ) );
  AOI22_X1 u2_uk_U583 (.B2( u2_uk_K_r4_3 ) , .A2( u2_uk_K_r4_54 ) , .ZN( u2_uk_n1058 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U588 (.ZN( u2_K16_22 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1205 ) , .A2( u2_uk_n1212 ) , .A1( u2_uk_n213 ) );
  INV_X1 u2_uk_U589 (.ZN( u2_K13_22 ) , .A( u2_uk_n634 ) );
  AOI22_X1 u2_uk_U590 (.B2( u2_uk_K_r11_10 ) , .A2( u2_uk_K_r11_47 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n634 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U593 (.ZN( u2_K10_22 ) , .A( u2_uk_n257 ) );
  INV_X1 u2_uk_U595 (.ZN( u2_K9_22 ) , .A( u2_uk_n1127 ) );
  AOI22_X1 u2_uk_U596 (.B2( u2_uk_K_r7_41 ) , .A2( u2_uk_K_r7_48 ) , .B1( u2_uk_n109 ) , .ZN( u2_uk_n1127 ) , .A1( u2_uk_n213 ) );
  INV_X1 u2_uk_U6 (.A( u2_uk_n146 ) , .ZN( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U605 (.ZN( u2_K11_35 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1665 ) , .A2( u2_uk_n1673 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U606 (.ZN( u2_K8_35 ) , .B2( u2_uk_n1511 ) , .A2( u2_uk_n1517 ) , .A1( u2_uk_n203 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U610 (.ZN( u2_K13_35 ) , .B2( u2_uk_n1734 ) , .A2( u2_uk_n1763 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U611 (.ZN( u2_K12_35 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1698 ) , .A2( u2_uk_n1707 ) , .B1( u2_uk_n230 ) );
  INV_X1 u2_uk_U614 (.ZN( u2_K10_35 ) , .A( u2_uk_n297 ) );
  AOI22_X1 u2_uk_U615 (.B2( u2_uk_K_r8_2 ) , .A2( u2_uk_K_r8_37 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n297 ) );
  OAI22_X1 u2_uk_U618 (.ZN( u2_K6_35 ) , .B2( u2_uk_n1439 ) , .A2( u2_uk_n1446 ) , .A1( u2_uk_n217 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U621 (.ZN( u2_K1_35 ) , .A( u2_uk_n982 ) );
  AOI22_X1 u2_uk_U622 (.B2( u2_key_r_28 ) , .A2( u2_key_r_35 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n982 ) );
  OAI21_X1 u2_uk_U623 (.ZN( u2_K16_11 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1212 ) , .A( u2_uk_n948 ) );
  INV_X1 u2_uk_U630 (.ZN( u2_K13_11 ) , .A( u2_uk_n526 ) );
  INV_X1 u2_uk_U635 (.ZN( u2_K9_11 ) , .A( u2_uk_n1118 ) );
  AOI22_X1 u2_uk_U636 (.B2( u2_uk_K_r7_48 ) , .A2( u2_uk_K_r7_55 ) , .B1( u2_uk_n100 ) , .ZN( u2_uk_n1118 ) , .A1( u2_uk_n223 ) );
  OAI21_X1 u2_uk_U640 (.ZN( u2_K2_11 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1267 ) , .A( u2_uk_n992 ) );
  NAND2_X1 u2_uk_U641 (.A1( u2_uk_K_r0_25 ) , .A2( u2_uk_n100 ) , .ZN( u2_uk_n992 ) );
  NAND2_X1 u2_uk_U643 (.A1( u2_uk_K_r2_24 ) , .ZN( u2_uk_n1039 ) , .A2( u2_uk_n60 ) );
  INV_X1 u2_uk_U644 (.ZN( u2_K1_44 ) , .A( u2_uk_n987 ) );
  AOI22_X1 u2_uk_U645 (.B2( u2_key_r_36 ) , .A2( u2_key_r_43 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n182 ) , .ZN( u2_uk_n987 ) );
  INV_X1 u2_uk_U650 (.A( u2_key_r_44 ) , .ZN( u2_uk_n1178 ) );
  OAI22_X1 u2_uk_U652 (.ZN( u2_K9_43 ) , .A1( u2_uk_n102 ) , .B2( u2_uk_n1558 ) , .A2( u2_uk_n1565 ) , .B1( u2_uk_n214 ) );
  OAI21_X1 u2_uk_U653 (.ZN( u2_K4_43 ) , .A( u2_uk_n1036 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1359 ) );
  OAI21_X1 u2_uk_U669 (.ZN( u2_K12_45 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1684 ) , .A( u2_uk_n509 ) );
  NAND2_X1 u2_uk_U670 (.A1( u2_uk_K_r10_43 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n509 ) );
  OAI22_X1 u2_uk_U671 (.ZN( u2_K11_43 ) , .A1( u2_uk_n161 ) , .B2( u2_uk_n1632 ) , .A2( u2_uk_n1674 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U680 (.ZN( u2_K6_7 ) , .A( u2_uk_n1072 ) , .B2( u2_uk_n1435 ) , .B1( u2_uk_n238 ) );
  NAND2_X1 u2_uk_U681 (.A1( u2_uk_K_r4_33 ) , .ZN( u2_uk_n1072 ) , .A2( u2_uk_n217 ) );
  NAND2_X1 u2_uk_U686 (.A1( u2_uk_K_r9_33 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n395 ) );
  OAI22_X1 u2_uk_U687 (.ZN( u2_K16_7 ) , .B2( u2_uk_n1199 ) , .A2( u2_uk_n1207 ) , .A1( u2_uk_n141 ) , .B1( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U689 (.ZN( u2_K13_25 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1735 ) , .A2( u2_uk_n1760 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U696 (.ZN( u2_K8_25 ) , .B2( u2_uk_n1533 ) , .A2( u2_uk_n1538 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n27 ) );
  INV_X1 u2_uk_U697 (.ZN( u2_K13_7 ) , .A( u2_uk_n682 ) );
  OAI22_X1 u2_uk_U70 (.ZN( u2_K16_23 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1213 ) , .A2( u2_uk_n1218 ) , .A1( u2_uk_n164 ) );
  INV_X1 u2_uk_U703 (.ZN( u2_K1_25 ) , .A( u2_uk_n975 ) );
  AOI22_X1 u2_uk_U704 (.B2( u2_key_r_29 ) , .A2( u2_key_r_36 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n975 ) );
  OAI22_X1 u2_uk_U715 (.ZN( u2_K8_32 ) , .B2( u2_uk_n1526 ) , .A2( u2_uk_n1533 ) , .A1( u2_uk_n238 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U716 (.ZN( u2_K11_32 ) , .B2( u2_uk_n1640 ) , .A2( u2_uk_n1660 ) , .A1( u2_uk_n203 ) , .B1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U73 (.ZN( u2_K10_23 ) , .B2( u2_uk_n1590 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n271 ) );
  INV_X1 u2_uk_U739 (.ZN( u2_K1_42 ) , .A( u2_uk_n986 ) );
  NAND2_X1 u2_uk_U74 (.A1( u2_uk_K_r8_13 ) , .A2( u2_uk_n129 ) , .ZN( u2_uk_n271 ) );
  OAI21_X1 u2_uk_U744 (.ZN( u2_K10_27 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1602 ) , .A( u2_uk_n279 ) );
  NAND2_X1 u2_uk_U745 (.A1( u2_uk_K_r8_43 ) , .ZN( u2_uk_n279 ) , .A2( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U746 (.ZN( u2_K8_27 ) , .B2( u2_uk_n1499 ) , .A2( u2_uk_n1504 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U752 (.ZN( u2_K2_13 ) , .A2( u2_uk_n1231 ) , .B2( u2_uk_n1260 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U754 (.ZN( u2_K9_13 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1120 ) , .B2( u2_uk_n1549 ) );
  OAI22_X1 u2_uk_U757 (.ZN( u2_K13_27 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1724 ) , .A2( u2_uk_n1747 ) , .B1( u2_uk_n222 ) );
  NAND2_X1 u2_uk_U760 (.A1( u2_uk_K_r9_5 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n346 ) );
  OAI22_X1 u2_uk_U761 (.ZN( u2_K9_21 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1568 ) , .A2( u2_uk_n1573 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U764 (.ZN( u2_K2_21 ) , .A2( u2_uk_n1234 ) , .B2( u2_uk_n1238 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U770 (.ZN( u2_K12_21 ) , .A( u2_uk_n443 ) );
  OAI21_X1 u2_uk_U772 (.ZN( u2_K3_27 ) , .A( u2_uk_n1009 ) , .B2( u2_uk_n1315 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U773 (.A1( u2_uk_K_r1_42 ) , .ZN( u2_uk_n1009 ) , .A2( u2_uk_n188 ) );
  INV_X1 u2_uk_U776 (.ZN( u2_K13_21 ) , .A( u2_uk_n608 ) );
  OAI21_X1 u2_uk_U780 (.ZN( u2_K16_13 ) , .B2( u2_uk_n1227 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n950 ) );
  NAND2_X1 u2_uk_U781 (.A1( u2_uk_K_r14_46 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n950 ) );
  INV_X1 u2_uk_U785 (.ZN( u2_K5_27 ) , .A( u2_uk_n1046 ) );
  INV_X1 u2_uk_U787 (.ZN( u2_K13_13 ) , .A( u2_uk_n582 ) );
  AOI22_X1 u2_uk_U788 (.B2( u2_uk_K_r11_11 ) , .A2( u2_uk_K_r11_6 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n582 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U79 (.ZN( u2_K2_23 ) , .B2( u2_uk_n1248 ) , .A2( u2_uk_n1269 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U791 (.ZN( u2_K1_27 ) , .A( u2_uk_n977 ) );
  AOI22_X1 u2_uk_U792 (.B2( u2_key_r_14 ) , .A2( u2_key_r_21 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n977 ) );
  INV_X1 u2_uk_U793 (.ZN( u2_K9_27 ) , .A( u2_uk_n1129 ) );
  AOI22_X1 u2_uk_U794 (.B2( u2_uk_K_r7_2 ) , .A2( u2_uk_K_r7_9 ) , .B1( u2_uk_n109 ) , .ZN( u2_uk_n1129 ) , .A1( u2_uk_n163 ) );
  OAI21_X1 u2_uk_U795 (.ZN( u2_K13_1 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1727 ) , .A( u2_uk_n603 ) );
  NAND2_X1 u2_uk_U796 (.A1( u2_uk_K_r11_25 ) , .ZN( u2_uk_n603 ) , .A2( u2_uk_n93 ) );
  INV_X1 u2_uk_U797 (.ZN( u2_K9_1 ) , .A( u2_uk_n1125 ) );
  INV_X1 u2_uk_U8 (.A( u2_uk_n145 ) , .ZN( u2_uk_n63 ) );
  NAND2_X1 u2_uk_U804 (.A1( u2_uk_K_r11_33 ) , .ZN( u2_uk_n605 ) , .A2( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U808 (.ZN( u2_K16_18 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1229 ) , .A( u2_uk_n953 ) );
  NAND2_X1 u2_uk_U809 (.A1( u2_uk_K_r14_5 ) , .A2( u2_uk_n109 ) , .ZN( u2_uk_n953 ) );
  OAI21_X1 u2_uk_U812 (.ZN( u2_K13_18 ) , .B2( u2_uk_n1750 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n590 ) );
  NAND2_X1 u2_uk_U813 (.A1( u2_uk_K_r11_20 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n590 ) );
  OAI22_X1 u2_uk_U817 (.ZN( u2_K16_20 ) , .B2( u2_uk_n1222 ) , .A2( u2_uk_n1229 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n209 ) );
  OAI21_X1 u2_uk_U82 (.ZN( u2_K11_41 ) , .B2( u2_uk_n1672 ) , .B1( u2_uk_n214 ) , .A( u2_uk_n382 ) );
  INV_X1 u2_uk_U820 (.ZN( u2_K9_18 ) , .A( u2_uk_n1123 ) );
  AOI22_X1 u2_uk_U821 (.B2( u2_uk_K_r7_39 ) , .A2( u2_uk_K_r7_46 ) , .B1( u2_uk_n110 ) , .ZN( u2_uk_n1123 ) , .A1( u2_uk_n163 ) );
  NAND2_X1 u2_uk_U83 (.A1( u2_uk_K_r9_31 ) , .A2( u2_uk_n203 ) , .ZN( u2_uk_n382 ) );
  NAND2_X1 u2_uk_U834 (.A1( u2_uk_K_r11_4 ) , .A2( u2_uk_n128 ) , .ZN( u2_uk_n672 ) );
  NAND2_X1 u2_uk_U841 (.A1( u2_uk_K_r3_10 ) , .ZN( u2_uk_n1056 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U849 (.ZN( u2_K15_22 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1828 ) , .A2( u2_uk_n1842 ) );
  OAI22_X1 u2_uk_U858 (.ZN( u2_K6_5 ) , .B2( u2_uk_n1422 ) , .A2( u2_uk_n1426 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U862 (.ZN( u2_K4_11 ) , .B2( u2_uk_n1333 ) , .A2( u2_uk_n1361 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U864 (.ZN( u2_K15_45 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1837 ) , .A2( u2_uk_n1855 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U866 (.ZN( u2_K12_43 ) , .B2( u2_uk_n1687 ) , .A2( u2_uk_n1707 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U867 (.ZN( u2_K6_45 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1424 ) , .A2( u2_uk_n1429 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U873 (.ZN( u2_K9_7 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1544 ) , .B2( u2_uk_n1548 ) );
  OAI22_X1 u2_uk_U874 (.ZN( u2_K6_12 ) , .A2( u2_uk_n1410 ) , .B2( u2_uk_n1426 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U877 (.ZN( u2_K13_24 ) , .B2( u2_uk_n1726 ) , .A2( u2_uk_n1767 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U881 (.ZN( u2_K9_24 ) , .B1( u2_uk_n128 ) , .B2( u2_uk_n1544 ) , .A2( u2_uk_n1586 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U884 (.ZN( u2_K2_24 ) , .A2( u2_uk_n1234 ) , .B2( u2_uk_n1249 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U885 (.ZN( u2_K16_21 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1197 ) , .A2( u2_uk_n1204 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U887 (.ZN( u2_K16_24 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1194 ) , .A2( u2_uk_n1199 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U894 (.ZN( u2_K2_17 ) , .A2( u2_uk_n1231 ) , .B2( u2_uk_n1247 ) , .A1( u2_uk_n145 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U896 (.ZN( u2_K3_25 ) , .B1( u2_uk_n117 ) , .B2( u2_uk_n1279 ) , .A2( u2_uk_n1283 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U900 (.ZN( u2_K6_42 ) , .B2( u2_uk_n1438 ) , .A2( u2_uk_n1445 ) , .A1( u2_uk_n163 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U901 (.ZN( u2_K6_39 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1411 ) , .B2( u2_uk_n1430 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U907 (.ZN( u2_K13_23 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1737 ) , .A2( u2_uk_n1767 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U909 (.ZN( u2_K9_47 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1576 ) , .A2( u2_uk_n1583 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U91 (.ZN( u2_K4_41 ) , .B2( u2_uk_n1319 ) , .A2( u2_uk_n1336 ) , .B1( u2_uk_n162 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U913 (.ZN( u2_K9_6 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1555 ) , .A2( u2_uk_n1563 ) , .B1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U914 (.ZN( u2_K9_8 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1573 ) , .A2( u2_uk_n1580 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U923 (.ZN( u2_K15_47 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1824 ) , .A2( u2_uk_n1856 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U928 (.ZN( u2_K6_46 ) , .A2( u2_uk_n1413 ) , .B2( u2_uk_n1441 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U929 (.ZN( u2_K13_4 ) , .B2( u2_uk_n1732 ) , .A2( u2_uk_n1737 ) , .B1( u2_uk_n187 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U930 (.ZN( u2_K9_4 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1549 ) , .A2( u2_uk_n1556 ) , .B1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U931 (.ZN( u2_K4_48 ) , .A1( u2_uk_n109 ) , .A2( u2_uk_n1325 ) , .B2( u2_uk_n1353 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U938 (.ZN( u2_K12_19 ) , .A1( u2_uk_n128 ) , .A2( u2_uk_n1682 ) , .B2( u2_uk_n1720 ) , .B1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U939 (.ZN( u2_K15_19 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1821 ) , .A2( u2_uk_n1851 ) , .B1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U940 (.ZN( u2_K10_20 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1599 ) , .A2( u2_uk_n1629 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U949 (.ZN( u2_K5_40 ) , .B2( u2_uk_n1383 ) , .A2( u2_uk_n1400 ) , .B1( u2_uk_n146 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U950 (.ZN( u2_K2_22 ) , .B2( u2_uk_n1243 ) , .A2( u2_uk_n1260 ) , .B1( u2_uk_n230 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U954 (.ZN( u2_K6_43 ) , .B2( u2_uk_n1408 ) , .A2( u2_uk_n1447 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U955 (.ZN( u2_K4_45 ) , .A1( u2_uk_n102 ) , .B2( u2_uk_n1321 ) , .A2( u2_uk_n1360 ) , .B1( u2_uk_n155 ) );
  INV_X1 u2_uk_U96 (.ZN( u2_K13_5 ) , .A( u2_uk_n678 ) );
  OAI22_X1 u2_uk_U965 (.ZN( u2_K1_34 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1144 ) , .A2( u2_uk_n1149 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U966 (.ZN( u2_K1_47 ) , .B2( u2_uk_n1142 ) , .A2( u2_uk_n1147 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U968 (.ZN( u2_K9_41 ) , .A( u2_uk_n1136 ) );
  AOI22_X1 u2_uk_U97 (.B2( u2_uk_K_r11_48 ) , .A2( u2_uk_K_r11_53 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n678 ) );
  INV_X1 u2_uk_U970 (.ZN( u2_K12_42 ) , .A( u2_uk_n503 ) );
  INV_X1 u2_uk_U972 (.ZN( u2_K9_42 ) , .A( u2_uk_n1137 ) );
  AOI22_X1 u2_uk_U974 (.B2( u2_uk_K_r11_19 ) , .A2( u2_uk_K_r11_24 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n681 ) );
  OAI21_X1 u2_uk_U985 (.ZN( u2_K4_5 ) , .A( u2_uk_n1038 ) , .B2( u2_uk_n1356 ) , .B1( u2_uk_n27 ) );
endmodule

