module des_des_die_0 ( clk, decrypt, desIn, key1, key2, key3, desOut, u0_out0_1, u0_out0_10, 
       u0_out0_11, u0_out0_12, u0_out0_13, u0_out0_14, u0_out0_15, u0_out0_16, u0_out0_17, u0_out0_18, u0_out0_19, 
       u0_out0_2, u0_out0_20, u0_out0_21, u0_out0_22, u0_out0_23, u0_out0_24, u0_out0_25, u0_out0_26, u0_out0_27, 
       u0_out0_28, u0_out0_29, u0_out0_3, u0_out0_30, u0_out0_31, u0_out0_32, u0_out0_4, u0_out0_5, u0_out0_6, 
       u0_out0_7, u0_out0_8, u0_out0_9, u0_out10_1, u0_out10_10, u0_out10_11, u0_out10_12, u0_out10_13, u0_out10_14, 
       u0_out10_15, u0_out10_16, u0_out10_17, u0_out10_18, u0_out10_19, u0_out10_2, u0_out10_20, u0_out10_21, u0_out10_22, 
       u0_out10_23, u0_out10_24, u0_out10_25, u0_out10_26, u0_out10_27, u0_out10_28, u0_out10_29, u0_out10_3, u0_out10_30, 
       u0_out10_31, u0_out10_32, u0_out10_4, u0_out10_5, u0_out10_6, u0_out10_7, u0_out10_8, u0_out10_9, u0_out11_1, 
       u0_out11_10, u0_out11_11, u0_out11_12, u0_out11_13, u0_out11_14, u0_out11_15, u0_out11_16, u0_out11_17, u0_out11_18, 
       u0_out11_19, u0_out11_2, u0_out11_20, u0_out11_21, u0_out11_22, u0_out11_23, u0_out11_24, u0_out11_25, u0_out11_26, 
       u0_out11_27, u0_out11_28, u0_out11_29, u0_out11_3, u0_out11_30, u0_out11_31, u0_out11_32, u0_out11_4, u0_out11_5, 
       u0_out11_6, u0_out11_7, u0_out11_8, u0_out11_9, u0_out12_1, u0_out12_10, u0_out12_11, u0_out12_12, u0_out12_13, 
       u0_out12_14, u0_out12_15, u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_19, u0_out12_2, u0_out12_20, u0_out12_21, 
       u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_25, u0_out12_26, u0_out12_27, u0_out12_28, u0_out12_29, u0_out12_3, 
       u0_out12_30, u0_out12_31, u0_out12_32, u0_out12_4, u0_out12_5, u0_out12_6, u0_out12_7, u0_out12_8, u0_out12_9, 
       u0_out13_1, u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_13, u0_out13_14, u0_out13_15, u0_out13_17, u0_out13_18, 
       u0_out13_19, u0_out13_2, u0_out13_20, u0_out13_21, u0_out13_22, u0_out13_23, u0_out13_25, u0_out13_26, u0_out13_27, 
       u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_31, u0_out13_32, u0_out13_4, u0_out13_5, u0_out13_7, u0_out13_8, 
       u0_out13_9, u0_out14_1, u0_out14_10, u0_out14_11, u0_out14_12, u0_out14_13, u0_out14_14, u0_out14_15, u0_out14_16, 
       u0_out14_18, u0_out14_19, u0_out14_2, u0_out14_20, u0_out14_21, u0_out14_22, u0_out14_24, u0_out14_25, u0_out14_26, 
       u0_out14_27, u0_out14_28, u0_out14_29, u0_out14_3, u0_out14_30, u0_out14_32, u0_out14_4, u0_out14_5, u0_out14_6, 
       u0_out14_7, u0_out14_8, u0_out15_1, u0_out15_10, u0_out15_11, u0_out15_12, u0_out15_13, u0_out15_14, u0_out15_15, 
       u0_out15_16, u0_out15_17, u0_out15_18, u0_out15_19, u0_out15_2, u0_out15_20, u0_out15_21, u0_out15_22, u0_out15_23, 
       u0_out15_24, u0_out15_25, u0_out15_26, u0_out15_27, u0_out15_28, u0_out15_29, u0_out15_3, u0_out15_30, u0_out15_31, 
       u0_out15_32, u0_out15_4, u0_out15_5, u0_out15_6, u0_out15_7, u0_out15_8, u0_out15_9, u0_out1_1, u0_out1_10, 
       u0_out1_11, u0_out1_12, u0_out1_13, u0_out1_14, u0_out1_16, u0_out1_17, u0_out1_18, u0_out1_19, u0_out1_2, 
       u0_out1_20, u0_out1_22, u0_out1_23, u0_out1_24, u0_out1_25, u0_out1_26, u0_out1_28, u0_out1_29, u0_out1_3, 
       u0_out1_30, u0_out1_31, u0_out1_32, u0_out1_4, u0_out1_6, u0_out1_7, u0_out1_8, u0_out1_9, u0_out2_1, 
       u0_out2_10, u0_out2_11, u0_out2_12, u0_out2_13, u0_out2_14, u0_out2_15, u0_out2_16, u0_out2_17, u0_out2_18, 
       u0_out2_19, u0_out2_2, u0_out2_20, u0_out2_21, u0_out2_22, u0_out2_23, u0_out2_24, u0_out2_25, u0_out2_26, 
       u0_out2_27, u0_out2_28, u0_out2_29, u0_out2_3, u0_out2_30, u0_out2_31, u0_out2_32, u0_out2_4, u0_out2_5, 
       u0_out2_6, u0_out2_7, u0_out2_8, u0_out2_9, u0_out3_1, u0_out3_10, u0_out3_11, u0_out3_12, u0_out3_13, 
       u0_out3_14, u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, u0_out3_20, u0_out3_21, 
       u0_out3_22, u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, u0_out3_29, u0_out3_3, 
       u0_out3_30, u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, u0_out3_8, u0_out3_9, 
       u0_out4_1, u0_out4_10, u0_out4_11, u0_out4_13, u0_out4_14, u0_out4_15, u0_out4_16, u0_out4_17, u0_out4_18, 
       u0_out4_19, u0_out4_2, u0_out4_20, u0_out4_21, u0_out4_23, u0_out4_24, u0_out4_25, u0_out4_26, u0_out4_27, 
       u0_out4_28, u0_out4_29, u0_out4_3, u0_out4_30, u0_out4_31, u0_out4_4, u0_out4_5, u0_out4_6, u0_out4_8, 
       u0_out4_9, u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, u0_out5_13, u0_out5_14, u0_out5_15, u0_out5_16, 
       u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, u0_out5_21, u0_out5_22, u0_out5_23, u0_out5_24, 
       u0_out5_25, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_3, u0_out5_30, u0_out5_31, u0_out5_32, 
       u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, u0_out5_9, u0_out6_1, u0_out6_10, u0_out6_11, 
       u0_out6_13, u0_out6_16, u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, u0_out6_23, u0_out6_24, 
       u0_out6_26, u0_out6_28, u0_out6_29, u0_out6_30, u0_out6_31, u0_out6_4, u0_out6_6, u0_out6_9, u0_out7_1, 
       u0_out7_10, u0_out7_11, u0_out7_12, u0_out7_13, u0_out7_14, u0_out7_15, u0_out7_16, u0_out7_17, u0_out7_18, 
       u0_out7_19, u0_out7_2, u0_out7_20, u0_out7_21, u0_out7_22, u0_out7_23, u0_out7_24, u0_out7_25, u0_out7_26, 
       u0_out7_27, u0_out7_28, u0_out7_29, u0_out7_3, u0_out7_30, u0_out7_31, u0_out7_32, u0_out7_4, u0_out7_5, 
       u0_out7_6, u0_out7_7, u0_out7_8, u0_out7_9, u0_out8_1, u0_out8_10, u0_out8_11, u0_out8_12, u0_out8_13, 
       u0_out8_14, u0_out8_15, u0_out8_16, u0_out8_17, u0_out8_18, u0_out8_19, u0_out8_2, u0_out8_20, u0_out8_21, 
       u0_out8_22, u0_out8_23, u0_out8_24, u0_out8_25, u0_out8_26, u0_out8_27, u0_out8_28, u0_out8_29, u0_out8_3, 
       u0_out8_30, u0_out8_31, u0_out8_32, u0_out8_4, u0_out8_5, u0_out8_6, u0_out8_7, u0_out8_8, u0_out8_9, 
       u0_out9_1, u0_out9_10, u0_out9_11, u0_out9_12, u0_out9_13, u0_out9_14, u0_out9_15, u0_out9_16, u0_out9_17, 
       u0_out9_18, u0_out9_19, u0_out9_2, u0_out9_20, u0_out9_21, u0_out9_22, u0_out9_23, u0_out9_24, u0_out9_25, 
       u0_out9_26, u0_out9_27, u0_out9_28, u0_out9_29, u0_out9_3, u0_out9_30, u0_out9_31, u0_out9_32, u0_out9_4, 
       u0_out9_5, u0_out9_6, u0_out9_7, u0_out9_8, u0_out9_9, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n109, 
       u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n129, u0_uk_n141, u0_uk_n142, u0_uk_n145, 
       u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, 
       u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n203, u0_uk_n207, u0_uk_n208, u0_uk_n209, 
       u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n230, u0_uk_n231, u0_uk_n238, 
       u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n27, u0_uk_n31, u0_uk_n60, u0_uk_n63, 
       u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_out0_1, u1_out0_10, u1_out0_11, u1_out0_12, 
       u1_out0_13, u1_out0_14, u1_out0_15, u1_out0_16, u1_out0_17, u1_out0_18, u1_out0_19, u1_out0_2, u1_out0_20, 
       u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_24, u1_out0_25, u1_out0_26, u1_out0_27, u1_out0_28, u1_out0_29, 
       u1_out0_3, u1_out0_30, u1_out0_31, u1_out0_32, u1_out0_4, u1_out0_5, u1_out0_6, u1_out0_7, u1_out0_8, 
       u1_out0_9, u1_out10_1, u1_out10_10, u1_out10_11, u1_out10_12, u1_out10_13, u1_out10_14, u1_out10_15, u1_out10_16, 
       u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_20, u1_out10_21, u1_out10_22, u1_out10_23, u1_out10_24, 
       u1_out10_25, u1_out10_26, u1_out10_27, u1_out10_28, u1_out10_29, u1_out10_3, u1_out10_30, u1_out10_31, u1_out10_32, 
       u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_8, u1_out10_9, u1_out11_1, u1_out11_10, u1_out11_11, 
       u1_out11_12, u1_out11_13, u1_out11_14, u1_out11_15, u1_out11_16, u1_out11_17, u1_out11_18, u1_out11_19, u1_out11_2, 
       u1_out11_20, u1_out11_21, u1_out11_22, u1_out11_23, u1_out11_24, u1_out11_25, u1_out11_26, u1_out11_27, u1_out11_28, 
       u1_out11_29, u1_out11_3, u1_out11_30, u1_out11_31, u1_out11_32, u1_out11_4, u1_out11_5, u1_out11_6, u1_out11_7, 
       u1_out11_8, u1_out11_9, u1_out12_1, u1_out12_10, u1_out12_11, u1_out12_12, u1_out12_13, u1_out12_14, u1_out12_15, 
       u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_19, u1_out12_2, u1_out12_20, u1_out12_21, u1_out12_22, u1_out12_23, 
       u1_out12_24, u1_out12_25, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_29, u1_out12_3, u1_out12_30, u1_out12_31, 
       u1_out12_32, u1_out12_4, u1_out12_5, u1_out12_6, u1_out12_7, u1_out12_8, u1_out12_9, u1_out13_1, u1_out13_10, 
       u1_out13_11, u1_out13_12, u1_out13_13, u1_out13_14, u1_out13_15, u1_out13_16, u1_out13_17, u1_out13_18, u1_out13_19, 
       u1_out13_2, u1_out13_20, u1_out13_21, u1_out13_22, u1_out13_23, u1_out13_24, u1_out13_25, u1_out13_26, u1_out13_27, 
       u1_out13_28, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_31, u1_out13_32, u1_out13_4, u1_out13_5, u1_out13_6, 
       u1_out13_7, u1_out13_8, u1_out13_9, u1_out14_1, u1_out14_10, u1_out14_11, u1_out14_12, u1_out14_13, u1_out14_14, 
       u1_out14_15, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_20, u1_out14_21, u1_out14_22, 
       u1_out14_23, u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_27, u1_out14_28, u1_out14_29, u1_out14_3, u1_out14_30, 
       u1_out14_31, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, u1_out14_8, u1_out14_9, u1_out15_1, 
       u1_out15_10, u1_out15_11, u1_out15_12, u1_out15_13, u1_out15_14, u1_out15_15, u1_out15_16, u1_out15_17, u1_out15_18, 
       u1_out15_19, u1_out15_2, u1_out15_20, u1_out15_21, u1_out15_22, u1_out15_23, u1_out15_24, u1_out15_25, u1_out15_26, 
       u1_out15_27, u1_out15_28, u1_out15_29, u1_out15_3, u1_out15_30, u1_out15_31, u1_out15_32, u1_out15_4, u1_out15_5, 
       u1_out15_6, u1_out15_7, u1_out15_8, u1_out15_9, u1_out1_1, u1_out1_10, u1_out1_11, u1_out1_12, u1_out1_13, 
       u1_out1_14, u1_out1_15, u1_out1_16, u1_out1_17, u1_out1_18, u1_out1_19, u1_out1_2, u1_out1_20, u1_out1_21, 
       u1_out1_22, u1_out1_23, u1_out1_24, u1_out1_25, u1_out1_26, u1_out1_27, u1_out1_28, u1_out1_29, u1_out1_3, 
       u1_out1_30, u1_out1_31, u1_out1_32, u1_out1_4, u1_out1_5, u1_out1_6, u1_out1_7, u1_out1_8, u1_out1_9, 
       u1_out2_1, u1_out2_10, u1_out2_11, u1_out2_12, u1_out2_13, u1_out2_14, u1_out2_15, u1_out2_16, u1_out2_17, 
       u1_out2_18, u1_out2_19, u1_out2_2, u1_out2_20, u1_out2_21, u1_out2_22, u1_out2_23, u1_out2_24, u1_out2_25, 
       u1_out2_26, u1_out2_27, u1_out2_28, u1_out2_29, u1_out2_3, u1_out2_30, u1_out2_31, u1_out2_32, u1_out2_4, 
       u1_out2_5, u1_out2_6, u1_out2_7, u1_out2_8, u1_out2_9, u1_out3_1, u1_out3_10, u1_out3_11, u1_out3_12, 
       u1_out3_13, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_17, u1_out3_18, u1_out3_19, u1_out3_2, u1_out3_20, 
       u1_out3_21, u1_out3_22, u1_out3_23, u1_out3_24, u1_out3_25, u1_out3_26, u1_out3_27, u1_out3_28, u1_out3_29, 
       u1_out3_3, u1_out3_30, u1_out3_31, u1_out3_32, u1_out3_4, u1_out3_5, u1_out3_6, u1_out3_7, u1_out3_8, 
       u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_11, u1_out4_12, u1_out4_13, u1_out4_14, u1_out4_15, u1_out4_16, 
       u1_out4_17, u1_out4_18, u1_out4_19, u1_out4_2, u1_out4_20, u1_out4_21, u1_out4_22, u1_out4_23, u1_out4_24, 
       u1_out4_25, u1_out4_26, u1_out4_27, u1_out4_28, u1_out4_29, u1_out4_3, u1_out4_30, u1_out4_31, u1_out4_32, 
       u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out4_9, u1_out5_1, u1_out5_10, u1_out5_11, 
       u1_out5_12, u1_out5_13, u1_out5_14, u1_out5_15, u1_out5_16, u1_out5_17, u1_out5_18, u1_out5_19, u1_out5_2, 
       u1_out5_20, u1_out5_21, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_25, u1_out5_26, u1_out5_27, u1_out5_28, 
       u1_out5_29, u1_out5_3, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_5, u1_out5_6, u1_out5_7, 
       u1_out5_8, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_11, u1_out6_12, u1_out6_13, u1_out6_14, u1_out6_15, 
       u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_19, u1_out6_2, u1_out6_20, u1_out6_21, u1_out6_22, u1_out6_23, 
       u1_out6_24, u1_out6_25, u1_out6_26, u1_out6_27, u1_out6_28, u1_out6_29, u1_out6_3, u1_out6_30, u1_out6_31, 
       u1_out6_32, u1_out6_4, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_8, u1_out6_9, u1_out7_1, u1_out7_10, 
       u1_out7_11, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_15, u1_out7_16, u1_out7_17, u1_out7_18, u1_out7_19, 
       u1_out7_2, u1_out7_20, u1_out7_21, u1_out7_22, u1_out7_23, u1_out7_24, u1_out7_25, u1_out7_26, u1_out7_27, 
       u1_out7_28, u1_out7_29, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, u1_out7_4, u1_out7_5, u1_out7_6, 
       u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_11, u1_out8_12, u1_out8_13, u1_out8_14, 
       u1_out8_15, u1_out8_16, u1_out8_17, u1_out8_18, u1_out8_19, u1_out8_2, u1_out8_20, u1_out8_21, u1_out8_22, 
       u1_out8_23, u1_out8_24, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_28, u1_out8_29, u1_out8_3, u1_out8_30, 
       u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_5, u1_out8_6, u1_out8_7, u1_out8_8, u1_out8_9, u1_out9_1, 
       u1_out9_10, u1_out9_11, u1_out9_12, u1_out9_13, u1_out9_14, u1_out9_15, u1_out9_16, u1_out9_17, u1_out9_18, 
       u1_out9_19, u1_out9_2, u1_out9_20, u1_out9_21, u1_out9_22, u1_out9_23, u1_out9_24, u1_out9_25, u1_out9_26, 
       u1_out9_27, u1_out9_28, u1_out9_29, u1_out9_3, u1_out9_30, u1_out9_31, u1_out9_32, u1_out9_4, u1_out9_5, 
       u1_out9_6, u1_out9_7, u1_out9_8, u1_out9_9, u2_out0_11, u2_out0_12, u2_out0_13, u2_out0_14, u2_out0_15, 
       u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, u2_out0_28, u2_out0_29, 
       u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, u2_out10_1, u2_out10_10, u2_out10_11, 
       u2_out10_12, u2_out10_13, u2_out10_14, u2_out10_15, u2_out10_16, u2_out10_18, u2_out10_19, u2_out10_2, u2_out10_20, 
       u2_out10_21, u2_out10_22, u2_out10_24, u2_out10_25, u2_out10_26, u2_out10_27, u2_out10_28, u2_out10_29, u2_out10_3, 
       u2_out10_30, u2_out10_32, u2_out10_4, u2_out10_5, u2_out10_6, u2_out10_7, u2_out10_8, u2_out11_1, u2_out11_10, 
       u2_out11_11, u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, u2_out11_16, u2_out11_17, u2_out11_18, u2_out11_19, 
       u2_out11_2, u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, u2_out11_24, u2_out11_25, u2_out11_26, u2_out11_27, 
       u2_out11_28, u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, u2_out11_32, u2_out11_4, u2_out11_5, u2_out11_6, 
       u2_out11_7, u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, u2_out12_13, u2_out12_14, u2_out12_15, u2_out12_17, 
       u2_out12_18, u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, u2_out12_23, u2_out12_25, u2_out12_27, u2_out12_28, 
       u2_out12_29, u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, u2_out12_5, u2_out12_7, u2_out12_8, u2_out12_9, 
       u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, u2_out13_21, u2_out13_22, u2_out13_25, u2_out13_27, 
       u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, u2_out13_7, u2_out13_8, u2_out14_1, u2_out14_10, 
       u2_out14_11, u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, u2_out14_16, u2_out14_17, u2_out14_18, u2_out14_19, 
       u2_out14_2, u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, u2_out14_24, u2_out14_25, u2_out14_26, u2_out14_27, 
       u2_out14_28, u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, u2_out14_32, u2_out14_4, u2_out14_5, u2_out14_6, 
       u2_out14_7, u2_out14_8, u2_out14_9, u2_out15_1, u2_out15_10, u2_out15_11, u2_out15_12, u2_out15_13, u2_out15_14, 
       u2_out15_15, u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_19, u2_out15_2, u2_out15_20, u2_out15_21, u2_out15_22, 
       u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_27, u2_out15_28, u2_out15_29, u2_out15_3, u2_out15_30, 
       u2_out15_31, u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_6, u2_out15_7, u2_out15_8, u2_out15_9, u2_out1_1, 
       u2_out1_10, u2_out1_11, u2_out1_12, u2_out1_13, u2_out1_14, u2_out1_15, u2_out1_16, u2_out1_17, u2_out1_18, 
       u2_out1_19, u2_out1_2, u2_out1_20, u2_out1_21, u2_out1_22, u2_out1_23, u2_out1_24, u2_out1_25, u2_out1_26, 
       u2_out1_27, u2_out1_28, u2_out1_29, u2_out1_3, u2_out1_30, u2_out1_31, u2_out1_32, u2_out1_4, u2_out1_5, 
       u2_out1_6, u2_out1_7, u2_out1_8, u2_out1_9, u2_out2_1, u2_out2_10, u2_out2_11, u2_out2_12, u2_out2_13, 
       u2_out2_14, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, u2_out2_20, u2_out2_21, 
       u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, u2_out2_29, u2_out2_3, 
       u2_out2_30, u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, u2_out2_8, u2_out2_9, 
       u2_out3_1, u2_out3_10, u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, u2_out3_16, u2_out3_17, u2_out3_18, 
       u2_out3_19, u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, u2_out3_25, u2_out3_26, u2_out3_27, 
       u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, u2_out3_5, u2_out3_6, u2_out3_8, 
       u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, u2_out4_15, u2_out4_16, 
       u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, u2_out4_23, u2_out4_24, 
       u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, u2_out4_31, u2_out4_32, 
       u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, u2_out5_10, u2_out5_11, 
       u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, u2_out5_19, u2_out5_2, 
       u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, u2_out5_27, u2_out5_28, 
       u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, u2_out5_6, u2_out5_7, 
       u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, u2_out6_14, u2_out6_15, 
       u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, u2_out6_22, u2_out6_23, 
       u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, u2_out6_30, u2_out6_31, 
       u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, u2_out7_1, u2_out7_10, 
       u2_out7_13, u2_out7_15, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, u2_out7_21, u2_out7_23, 
       u2_out7_24, u2_out7_26, u2_out7_27, u2_out7_28, u2_out7_30, u2_out7_31, u2_out7_5, u2_out7_6, u2_out7_9, 
       u2_out8_1, u2_out8_10, u2_out8_11, u2_out8_12, u2_out8_13, u2_out8_14, u2_out8_15, u2_out8_16, u2_out8_17, 
       u2_out8_18, u2_out8_19, u2_out8_2, u2_out8_20, u2_out8_21, u2_out8_22, u2_out8_23, u2_out8_24, u2_out8_25, 
       u2_out8_26, u2_out8_27, u2_out8_28, u2_out8_29, u2_out8_3, u2_out8_30, u2_out8_31, u2_out8_32, u2_out8_4, 
       u2_out8_5, u2_out8_6, u2_out8_7, u2_out8_8, u2_out8_9, u2_out9_1, u2_out9_10, u2_out9_11, u2_out9_12, 
       u2_out9_13, u2_out9_14, u2_out9_15, u2_out9_16, u2_out9_17, u2_out9_18, u2_out9_19, u2_out9_2, u2_out9_20, 
       u2_out9_21, u2_out9_22, u2_out9_23, u2_out9_24, u2_out9_25, u2_out9_26, u2_out9_27, u2_out9_28, u2_out9_29, 
       u2_out9_3, u2_out9_30, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_6, u2_out9_7, u2_out9_8, 
       u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n117, u2_uk_n118, 
       u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
       u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n182, u2_uk_n187, u2_uk_n188, u2_uk_n191, 
       u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, 
       u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, u2_uk_n31, u2_uk_n60, u2_uk_n63, u2_uk_n83, 
       u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99, u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_39, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, 
        u0_FP_45, u0_FP_46, u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_55, 
        u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_63, u0_FP_64, u0_K10_1, u0_K10_14, 
        u0_K10_17, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_32, u0_K11_37, u0_K11_42, u0_K11_48, u0_K12_19, 
        u0_K12_25, u0_K12_35, u0_K12_36, u0_K12_48, u0_K12_5, u0_K12_7, u0_K12_8, u0_K13_41, u0_K14_23, 
        u0_K14_24, u0_K14_25, u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K15_13, u0_K16_18, u0_K16_19, 
        u0_K16_24, u0_K16_26, u0_K16_36, u0_K16_38, u0_K16_5, u0_K16_8, u0_K1_13, u0_K1_14, u0_K1_17, 
        u0_K1_30, u0_K1_31, u0_K2_11, u0_K2_12, u0_K2_18, u0_K2_20, u0_K2_29, u0_K2_30, u0_K2_31, 
        u0_K2_5, u0_K3_12, u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_5, 
        u0_K3_6, u0_K4_36, u0_K4_43, u0_K4_48, u0_K4_6, u0_K5_1, u0_K5_18, u0_K5_24, u0_K5_26, 
        u0_K5_29, u0_K5_31, u0_K5_47, u0_K5_8, u0_K6_11, u0_K6_13, u0_K6_19, u0_K6_20, u0_K6_23, 
        u0_K6_24, u0_K6_41, u0_K8_11, u0_K8_13, u0_K8_19, u0_K9_12, u0_K9_13, u0_K9_14, u0_K9_30, 
        u0_K9_32, u0_K9_44, u0_K9_6, u0_R0_1, u0_R0_13, u0_R0_15, u0_R0_18, u0_R0_19, u0_R0_20, 
        u0_R0_21, u0_R0_28, u0_R0_32, u0_R0_4, u0_R0_7, u0_R0_8, u0_R0_9, u0_R10_1, u0_R10_12, 
        u0_R10_14, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_24, 
        u0_R10_25, u0_R10_28, u0_R10_29, u0_R10_3, u0_R10_4, u0_R10_5, u0_R11_10, u0_R11_11, u0_R11_12, 
        u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_2, u0_R11_20, u0_R11_28, u0_R11_3, u0_R11_32, 
        u0_R11_5, u0_R11_6, u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, u0_R12_23, u0_R12_24, 
        u0_R12_30, u0_R12_4, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, 
        u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, u0_R13_8, 
        u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, u0_R1_19, u0_R1_20, u0_R1_21, 
        u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_30, 
        u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, 
        u0_R2_13, u0_R2_14, u0_R2_16, u0_R2_2, u0_R2_21, u0_R2_22, u0_R2_25, u0_R2_28, u0_R2_3, 
        u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_13, u0_R3_15, 
        u0_R3_17, u0_R3_18, u0_R3_20, u0_R3_22, u0_R3_24, u0_R3_25, u0_R3_32, u0_R3_5, u0_R4_1, 
        u0_R4_12, u0_R4_13, u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_24, 
        u0_R4_25, u0_R4_26, u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, u0_R4_4, 
        u0_R4_5, u0_R4_8, u0_R4_9, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, u0_R5_32, 
        u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, 
        u0_R6_14, u0_R6_17, u0_R6_24, u0_R6_26, u0_R6_28, u0_R6_29, u0_R6_4, u0_R6_5, u0_R6_7, 
        u0_R6_8, u0_R6_9, u0_R7_1, u0_R7_12, u0_R7_14, u0_R7_17, u0_R7_20, u0_R7_21, u0_R7_22, 
        u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_28, u0_R7_29, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_8, 
        u0_R7_9, u0_R8_1, u0_R8_12, u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, 
        u0_R8_27, u0_R8_29, u0_R8_30, u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_R9_1, u0_R9_10, 
        u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, 
        u0_R9_21, u0_R9_22, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_29, u0_R9_3, u0_R9_30, 
        u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_1, 
        u0_desIn_r_11, u0_desIn_r_15, u0_desIn_r_17, u0_desIn_r_23, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, 
        u0_desIn_r_35, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_51, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_59, 
        u0_desIn_r_63, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_14, u0_key_r_16, 
        u0_key_r_19, u0_key_r_2, u0_key_r_20, u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, 
        u0_key_r_35, u0_key_r_4, u0_key_r_41, u0_key_r_42, u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_50, u0_key_r_54, 
        u0_key_r_55, u0_key_r_6, u0_key_r_9, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, u0_u0_X_25, 
        u0_u0_X_28, u0_u0_X_33, u0_u0_X_42, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u10_X_22, u0_u10_X_34, 
        u0_u10_X_41, u0_u10_X_43, u0_u11_X_1, u0_u11_X_10, u0_u11_X_11, u0_u11_X_12, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, 
        u0_u11_X_16, u0_u11_X_18, u0_u11_X_20, u0_u11_X_22, u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u11_X_45, 
        u0_u11_X_46, u0_u11_X_47, u0_u11_X_9, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, u0_u12_X_2, 
        u0_u12_X_24, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, 
        u0_u12_X_36, u0_u12_X_37, u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, 
        u0_u12_X_48, u0_u12_X_5, u0_u12_X_7, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, u0_u13_X_2, 
        u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, u0_u13_X_38, 
        u0_u13_X_39, u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, 
        u0_u13_X_48, u0_u13_X_6, u0_u13_X_8, u0_u13_X_9, u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, 
        u0_u14_X_17, u0_u14_X_18, u0_u14_X_19, u0_u14_X_20, u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_25, 
        u0_u14_X_47, u0_u14_X_48, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_11, u0_u15_X_13, u0_u15_X_22, u0_u15_X_33, 
        u0_u15_X_4, u0_u15_X_42, u0_u15_X_44, u0_u15_X_45, u0_u15_X_9, u0_u1_X_15, u0_u1_X_16, u0_u1_X_17, u0_u1_X_19, 
        u0_u1_X_21, u0_u1_X_23, u0_u1_X_24, u0_u1_X_25, u0_u1_X_26, u0_u1_X_3, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, 
        u0_u1_X_36, u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_4, u0_u1_X_40, u0_u1_X_42, u0_u1_X_6, u0_u1_X_8, 
        u0_u1_X_9, u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_24, u0_u2_X_26, u0_u2_X_27, u0_u2_X_3, u0_u2_X_34, 
        u0_u2_X_46, u0_u2_X_9, u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, u0_u3_X_31, 
        u0_u3_X_34, u0_u3_X_35, u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, u0_u3_X_46, 
        u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, u0_u4_X_19, 
        u0_u4_X_2, u0_u4_X_21, u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, u0_u4_X_34, 
        u0_u4_X_4, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, u0_u4_X_9, 
        u0_u5_X_10, u0_u5_X_15, u0_u5_X_16, u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, 
        u0_u5_X_9, u0_u6_X_15, u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, 
        u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, 
        u0_u7_X_25, u0_u7_X_27, u0_u7_X_28, u0_u7_X_29, u0_u7_X_3, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, 
        u0_u7_X_34, u0_u7_X_36, u0_u7_X_38, u0_u7_X_4, u0_u7_X_40, u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, 
        u0_u7_X_9, u0_u8_X_10, u0_u8_X_15, u0_u8_X_16, u0_u8_X_18, u0_u8_X_20, u0_u8_X_22, u0_u8_X_23, u0_u8_X_25, 
        u0_u8_X_27, u0_u8_X_28, u0_u8_X_3, u0_u8_X_39, u0_u8_X_4, u0_u8_X_40, u0_u8_X_45, u0_u8_X_46, u0_u8_X_9, 
        u0_u9_X_10, u0_u9_X_11, u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, 
        u0_u9_X_27, u0_u9_X_3, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, 
        u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r0_15, u0_uk_K_r0_28, u0_uk_K_r0_36, u0_uk_K_r0_49, 
        u0_uk_K_r0_7, u0_uk_K_r10_10, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_37, u0_uk_K_r10_41, 
        u0_uk_K_r10_42, u0_uk_K_r10_44, u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, 
        u0_uk_K_r11_33, u0_uk_K_r11_39, u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_0, u0_uk_K_r13_25, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r14_10, 
        u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_50, u0_uk_K_r14_8, 
        u0_uk_K_r14_9, u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, 
        u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, 
        u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, u0_uk_K_r4_35, u0_uk_K_r4_38, 
        u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_0, u0_uk_K_r6_22, u0_uk_K_r6_26, 
        u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r7_26, u0_uk_K_r8_16, u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r9_0, u0_uk_K_r9_1, 
        u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_6, 
        u0_uk_K_r9_7, u0_uk_K_r9_9, u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1005, u0_uk_n1006, u0_uk_n101, 
        u0_uk_n1012, u0_uk_n1024, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n12, 
        u0_uk_n121, u0_uk_n122, u0_uk_n123, u0_uk_n126, u0_uk_n127, u0_uk_n13, u0_uk_n131, u0_uk_n139, u0_uk_n143, 
        u0_uk_n144, u0_uk_n151, u0_uk_n153, u0_uk_n156, u0_uk_n167, u0_uk_n168, u0_uk_n171, u0_uk_n172, u0_uk_n173, 
        u0_uk_n174, u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, u0_uk_n181, u0_uk_n183, u0_uk_n184, 
        u0_uk_n185, u0_uk_n189, u0_uk_n190, u0_uk_n192, u0_uk_n193, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, 
        u0_uk_n199, u0_uk_n200, u0_uk_n201, u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n21, u0_uk_n210, u0_uk_n211, 
        u0_uk_n212, u0_uk_n215, u0_uk_n216, u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n221, u0_uk_n224, u0_uk_n225, 
        u0_uk_n23, u0_uk_n232, u0_uk_n233, u0_uk_n239, u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, 
        u0_uk_n253, u0_uk_n257, u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, 
        u0_uk_n272, u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n289, 
        u0_uk_n290, u0_uk_n293, u0_uk_n3, u0_uk_n300, u0_uk_n307, u0_uk_n310, u0_uk_n314, u0_uk_n316, u0_uk_n318, 
        u0_uk_n32, u0_uk_n320, u0_uk_n324, u0_uk_n329, u0_uk_n33, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n336, 
        u0_uk_n337, u0_uk_n339, u0_uk_n341, u0_uk_n344, u0_uk_n347, u0_uk_n348, u0_uk_n352, u0_uk_n355, u0_uk_n358, 
        u0_uk_n361, u0_uk_n370, u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n396, 
        u0_uk_n4, u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n410, u0_uk_n411, u0_uk_n412, 
        u0_uk_n413, u0_uk_n414, u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, 
        u0_uk_n428, u0_uk_n429, u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, u0_uk_n439, 
        u0_uk_n440, u0_uk_n442, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n45, u0_uk_n450, u0_uk_n457, 
        u0_uk_n471, u0_uk_n497, u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, u0_uk_n511, 
        u0_uk_n513, u0_uk_n517, u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, 
        u0_uk_n532, u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n542, u0_uk_n544, u0_uk_n545, u0_uk_n546, 
        u0_uk_n547, u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, u0_uk_n555, u0_uk_n557, 
        u0_uk_n558, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, u0_uk_n567, u0_uk_n568, u0_uk_n570, 
        u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n577, u0_uk_n578, u0_uk_n579, u0_uk_n58, u0_uk_n580, u0_uk_n581, 
        u0_uk_n583, u0_uk_n598, u0_uk_n604, u0_uk_n61, u0_uk_n615, u0_uk_n627, u0_uk_n629, u0_uk_n632, u0_uk_n635, 
        u0_uk_n636, u0_uk_n637, u0_uk_n639, u0_uk_n640, u0_uk_n642, u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n649, 
        u0_uk_n650, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n654, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n660, 
        u0_uk_n661, u0_uk_n663, u0_uk_n666, u0_uk_n668, u0_uk_n669, u0_uk_n67, u0_uk_n670, u0_uk_n674, u0_uk_n675, 
        u0_uk_n684, u0_uk_n687, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, u0_uk_n711, u0_uk_n719, u0_uk_n722, 
        u0_uk_n723, u0_uk_n725, u0_uk_n726, u0_uk_n727, u0_uk_n729, u0_uk_n73, u0_uk_n731, u0_uk_n734, u0_uk_n735, 
        u0_uk_n741, u0_uk_n746, u0_uk_n748, u0_uk_n751, u0_uk_n759, u0_uk_n761, u0_uk_n763, u0_uk_n768, u0_uk_n780, 
        u0_uk_n783, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n8, u0_uk_n800, u0_uk_n809, u0_uk_n810, u0_uk_n813, 
        u0_uk_n815, u0_uk_n816, u0_uk_n832, u0_uk_n839, u0_uk_n855, u0_uk_n866, u0_uk_n868, u0_uk_n869, u0_uk_n875, 
        u0_uk_n883, u0_uk_n892, u0_uk_n898, u0_uk_n9, u0_uk_n904, u0_uk_n91, u0_uk_n915, u0_uk_n916, u0_uk_n917, 
        u0_uk_n918, u0_uk_n933, u0_uk_n934, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n963, u0_uk_n976, 
        u0_uk_n98, u0_uk_n982, u0_uk_n985, u0_uk_n990, u0_uk_n999, u1_FP_33, u1_FP_37, u1_FP_40, u1_FP_41, 
        u1_FP_44, u1_FP_45, u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, u1_FP_60, u1_FP_61, u1_K10_1, 
        u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_18, u1_K10_2, u1_K10_20, u1_K10_23, u1_K10_24, u1_K10_25, 
        u1_K10_26, u1_K10_29, u1_K10_30, u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, 
        u1_K10_44, u1_K10_47, u1_K10_48, u1_K10_5, u1_K10_6, u1_K10_7, u1_K10_8, u1_K11_11, u1_K11_13, 
        u1_K11_2, u1_K11_23, u1_K11_25, u1_K11_29, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, 
        u1_K11_7, u1_K12_18, u1_K12_19, u1_K12_2, u1_K12_20, u1_K12_24, u1_K12_25, u1_K12_26, u1_K12_35, 
        u1_K12_36, u1_K12_37, u1_K12_38, u1_K12_41, u1_K12_43, u1_K12_47, u1_K12_48, u1_K12_6, u1_K12_8, 
        u1_K13_14, u1_K13_17, u1_K13_18, u1_K13_20, u1_K13_29, u1_K13_30, u1_K13_31, u1_K13_32, u1_K13_35, 
        u1_K13_37, u1_K13_48, u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_29, u1_K14_30, u1_K14_31, u1_K14_32, 
        u1_K14_42, u1_K14_44, u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, 
        u1_K15_2, u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, 
        u1_K15_36, u1_K15_37, u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, 
        u1_K16_11, u1_K16_12, u1_K16_13, u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_2, u1_K16_20, 
        u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_35, u1_K16_41, u1_K16_42, u1_K16_44, u1_K16_48, u1_K16_6, 
        u1_K16_8, u1_K1_1, u1_K1_17, u1_K1_19, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_1, 
        u1_K2_11, u1_K2_12, u1_K2_13, u1_K2_17, u1_K2_18, u1_K2_2, u1_K2_20, u1_K2_23, u1_K2_24, 
        u1_K2_25, u1_K2_26, u1_K2_29, u1_K2_30, u1_K2_31, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, 
        u1_K2_48, u1_K2_5, u1_K2_6, u1_K2_8, u1_K3_1, u1_K3_12, u1_K3_14, u1_K3_17, u1_K3_18, 
        u1_K3_19, u1_K3_2, u1_K3_20, u1_K3_23, u1_K3_25, u1_K3_26, u1_K3_29, u1_K3_31, u1_K3_35, 
        u1_K3_36, u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, 
        u1_K3_5, u1_K3_6, u1_K3_7, u1_K3_8, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_13, u1_K4_14, 
        u1_K4_17, u1_K4_18, u1_K4_19, u1_K4_24, u1_K4_30, u1_K4_32, u1_K4_35, u1_K4_36, u1_K4_37, 
        u1_K4_38, u1_K4_41, u1_K4_42, u1_K4_43, u1_K4_44, u1_K4_47, u1_K4_48, u1_K4_6, u1_K5_1, 
        u1_K5_11, u1_K5_12, u1_K5_13, u1_K5_14, u1_K5_17, u1_K5_18, u1_K5_19, u1_K5_2, u1_K5_23, 
        u1_K5_24, u1_K5_25, u1_K5_26, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_37, u1_K5_38, 
        u1_K5_41, u1_K5_42, u1_K5_44, u1_K5_47, u1_K5_48, u1_K5_5, u1_K5_6, u1_K5_7, u1_K5_8, 
        u1_K6_1, u1_K6_11, u1_K6_12, u1_K6_13, u1_K6_14, u1_K6_20, u1_K6_23, u1_K6_24, u1_K6_25, 
        u1_K6_26, u1_K6_29, u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, 
        u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_47, u1_K6_48, u1_K6_5, u1_K6_6, u1_K6_7, 
        u1_K6_8, u1_K7_1, u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_19, u1_K7_2, u1_K7_23, 
        u1_K7_26, u1_K7_29, u1_K7_30, u1_K7_31, u1_K7_35, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, 
        u1_K7_44, u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_7, u1_K8_1, u1_K8_11, u1_K8_13, u1_K8_14, 
        u1_K8_18, u1_K8_2, u1_K8_20, u1_K8_23, u1_K8_24, u1_K8_25, u1_K8_26, u1_K8_30, u1_K8_31, 
        u1_K8_32, u1_K8_35, u1_K8_36, u1_K8_38, u1_K8_41, u1_K8_42, u1_K8_44, u1_K8_47, u1_K8_48, 
        u1_K8_5, u1_K8_7, u1_K9_12, u1_K9_13, u1_K9_14, u1_K9_17, u1_K9_23, u1_K9_24, u1_K9_25, 
        u1_K9_29, u1_K9_31, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, 
        u1_K9_6, u1_K9_7, u1_K9_8, u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, 
        u1_R0_21, u1_R0_28, u1_R0_29, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_7, u1_R0_8, u1_R0_9, 
        u1_R10_1, u1_R10_10, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_16, u1_R10_17, u1_R10_24, u1_R10_25, 
        u1_R10_28, u1_R10_29, u1_R10_32, u1_R10_5, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_20, 
        u1_R11_21, u1_R11_24, u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_20, u1_R12_21, 
        u1_R12_23, u1_R12_29, u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, 
        u1_R13_24, u1_R13_25, u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, 
        u1_R1_12, u1_R1_13, u1_R1_16, u1_R1_17, u1_R1_20, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, 
        u1_R1_32, u1_R1_4, u1_R1_5, u1_R1_9, u1_R2_1, u1_R2_12, u1_R2_13, u1_R2_16, u1_R2_17, 
        u1_R2_2, u1_R2_20, u1_R2_21, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_32, u1_R2_5, 
        u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, u1_R3_17, 
        u1_R3_18, u1_R3_20, u1_R3_21, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_32, u1_R3_4, 
        u1_R3_5, u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_13, u1_R4_14, u1_R4_16, u1_R4_17, u1_R4_20, 
        u1_R4_21, u1_R4_24, u1_R4_25, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, 
        u1_R4_6, u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_12, u1_R5_13, u1_R5_16, u1_R5_17, 
        u1_R5_18, u1_R5_20, u1_R5_21, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, 
        u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_8, u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_13, u1_R6_16, 
        u1_R6_17, u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_28, u1_R6_29, u1_R6_32, 
        u1_R6_4, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, 
        u1_R7_18, u1_R7_20, u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, 
        u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_13, u1_R8_15, u1_R8_16, u1_R8_17, 
        u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R8_4, 
        u1_R8_5, u1_R8_6, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_12, u1_R9_15, u1_R9_16, u1_R9_20, 
        u1_R9_21, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, u1_desIn_r_25, u1_desIn_r_29, 
        u1_desIn_r_37, u1_desIn_r_39, u1_desIn_r_57, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_13, u1_u0_X_14, u1_u0_X_15, 
        u1_u0_X_16, u1_u0_X_2, u1_u0_X_21, u1_u0_X_22, u1_u0_X_23, u1_u0_X_24, u1_u0_X_25, u1_u0_X_26, u1_u0_X_27, 
        u1_u0_X_28, u1_u0_X_29, u1_u0_X_3, u1_u0_X_30, u1_u0_X_31, u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, 
        u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, 
        u1_u0_X_46, u1_u0_X_48, u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, 
        u1_u10_X_18, u1_u10_X_20, u1_u10_X_21, u1_u10_X_24, u1_u10_X_26, u1_u10_X_27, u1_u10_X_28, u1_u10_X_3, u1_u10_X_33, 
        u1_u10_X_39, u1_u10_X_4, u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, 
        u1_u10_X_47, u1_u10_X_6, u1_u10_X_8, u1_u10_X_9, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, u1_u11_X_14, 
        u1_u11_X_16, u1_u11_X_22, u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_3, u1_u11_X_30, u1_u11_X_31, u1_u11_X_32, 
        u1_u11_X_33, u1_u11_X_34, u1_u11_X_39, u1_u11_X_4, u1_u11_X_40, u1_u11_X_45, u1_u11_X_46, u1_u11_X_5, u1_u11_X_7, 
        u1_u11_X_9, u1_u12_X_1, u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, u1_u12_X_25, 
        u1_u12_X_26, u1_u12_X_27, u1_u12_X_28, u1_u12_X_3, u1_u12_X_33, u1_u12_X_34, u1_u12_X_36, u1_u12_X_38, u1_u12_X_39, 
        u1_u12_X_4, u1_u12_X_40, u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, 
        u1_u12_X_9, u1_u13_X_10, u1_u13_X_11, u1_u13_X_12, u1_u13_X_13, u1_u13_X_14, u1_u13_X_15, u1_u13_X_16, u1_u13_X_17, 
        u1_u13_X_18, u1_u13_X_19, u1_u13_X_20, u1_u13_X_21, u1_u13_X_22, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, 
        u1_u13_X_27, u1_u13_X_28, u1_u13_X_3, u1_u13_X_33, u1_u13_X_35, u1_u13_X_36, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, 
        u1_u13_X_4, u1_u13_X_40, u1_u13_X_41, u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, 
        u1_u13_X_8, u1_u13_X_9, u1_u14_X_1, u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, 
        u1_u14_X_22, u1_u14_X_27, u1_u14_X_28, u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, 
        u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, u1_u14_X_9, u1_u15_X_1, u1_u15_X_10, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, 
        u1_u15_X_22, u1_u15_X_23, u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, u1_u15_X_27, u1_u15_X_28, u1_u15_X_3, u1_u15_X_33, 
        u1_u15_X_36, u1_u15_X_38, u1_u15_X_39, u1_u15_X_4, u1_u15_X_40, u1_u15_X_45, u1_u15_X_46, u1_u15_X_47, u1_u15_X_5, 
        u1_u15_X_7, u1_u15_X_9, u1_u1_X_15, u1_u1_X_16, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_3, 
        u1_u1_X_33, u1_u1_X_34, u1_u1_X_35, u1_u1_X_36, u1_u1_X_37, u1_u1_X_38, u1_u1_X_39, u1_u1_X_4, u1_u1_X_40, 
        u1_u1_X_45, u1_u1_X_46, u1_u1_X_9, u1_u2_X_10, u1_u2_X_11, u1_u2_X_13, u1_u2_X_15, u1_u2_X_16, u1_u2_X_21, 
        u1_u2_X_22, u1_u2_X_27, u1_u2_X_28, u1_u2_X_3, u1_u2_X_30, u1_u2_X_32, u1_u2_X_33, u1_u2_X_34, u1_u2_X_39, 
        u1_u2_X_4, u1_u2_X_40, u1_u2_X_45, u1_u2_X_46, u1_u2_X_9, u1_u3_X_15, u1_u3_X_16, u1_u3_X_21, u1_u3_X_22, 
        u1_u3_X_27, u1_u3_X_28, u1_u3_X_33, u1_u3_X_34, u1_u3_X_39, u1_u3_X_4, u1_u3_X_40, u1_u3_X_45, u1_u3_X_46, 
        u1_u3_X_5, u1_u3_X_7, u1_u3_X_9, u1_u4_X_10, u1_u4_X_15, u1_u4_X_16, u1_u4_X_21, u1_u4_X_28, u1_u4_X_3, 
        u1_u4_X_33, u1_u4_X_34, u1_u4_X_39, u1_u4_X_4, u1_u4_X_40, u1_u4_X_45, u1_u4_X_46, u1_u4_X_9, u1_u5_X_15, 
        u1_u5_X_16, u1_u5_X_17, u1_u5_X_19, u1_u5_X_22, u1_u5_X_27, u1_u5_X_28, u1_u5_X_3, u1_u5_X_33, u1_u5_X_34, 
        u1_u5_X_39, u1_u5_X_40, u1_u5_X_45, u1_u5_X_46, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_21, u1_u6_X_22, 
        u1_u6_X_28, u1_u6_X_3, u1_u6_X_33, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, u1_u6_X_45, u1_u6_X_9, u1_u7_X_10, 
        u1_u7_X_16, u1_u7_X_17, u1_u7_X_19, u1_u7_X_21, u1_u7_X_22, u1_u7_X_27, u1_u7_X_28, u1_u7_X_33, u1_u7_X_34, 
        u1_u7_X_39, u1_u7_X_4, u1_u7_X_40, u1_u7_X_45, u1_u7_X_46, u1_u7_X_6, u1_u7_X_8, u1_u7_X_9, u1_u8_X_15, 
        u1_u8_X_16, u1_u8_X_21, u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, u1_u8_X_39, 
        u1_u8_X_4, u1_u8_X_40, u1_u8_X_45, u1_u8_X_46, u1_u9_X_10, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_19, 
        u1_u9_X_21, u1_u9_X_27, u1_u9_X_28, u1_u9_X_3, u1_u9_X_34, u1_u9_X_39, u1_u9_X_4, u1_u9_X_40, u1_u9_X_45, 
        u1_u9_X_46, u1_uk_n1002, u1_uk_n1003, u1_uk_n1015, u1_uk_n1021, u1_uk_n1023, u1_uk_n1025, u1_uk_n1029, u1_uk_n1031, 
        u1_uk_n1034, u1_uk_n1038, u1_uk_n1050, u1_uk_n1054, u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1060, u1_uk_n1061, 
        u1_uk_n1063, u1_uk_n1065, u1_uk_n1070, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, 
        u1_uk_n1088, u1_uk_n1090, u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, 
        u1_uk_n1113, u1_uk_n1114, u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1121, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, 
        u1_uk_n1126, u1_uk_n1128, u1_uk_n1130, u1_uk_n1134, u1_uk_n1138, u1_uk_n1140, u1_uk_n1143, u1_uk_n1147, u1_uk_n1148, 
        u1_uk_n1153, u1_uk_n1154, u1_uk_n1155, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, 
        u1_uk_n1166, u1_uk_n1167, u1_uk_n1170, u1_uk_n1171, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, u1_uk_n366, 
        u1_uk_n369, u1_uk_n376, u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n386, u1_uk_n407, u1_uk_n421, u1_uk_n437, 
        u1_uk_n443, u1_uk_n454, u1_uk_n496, u1_uk_n504, u1_uk_n509, u1_uk_n515, u1_uk_n520, u1_uk_n524, u1_uk_n605, 
        u1_uk_n608, u1_uk_n672, u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, u1_uk_n949, 
        u1_uk_n950, u1_uk_n955, u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, 
        u1_uk_n989, u1_uk_n993, u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, 
        u2_FP_48, u2_FP_49, u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, 
        u2_FP_64, u2_K10_1, u2_K10_11, u2_K10_13, u2_K10_14, u2_K10_17, u2_K10_18, u2_K10_19, u2_K10_20, 
        u2_K10_23, u2_K10_24, u2_K10_25, u2_K10_26, u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, 
        u2_K10_5, u2_K10_7, u2_K10_8, u2_K11_11, u2_K11_13, u2_K11_24, u2_K11_26, u2_K11_29, u2_K12_2, 
        u2_K12_20, u2_K12_25, u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, u2_K13_37, 
        u2_K13_48, u2_K14_38, u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, u2_K15_31, 
        u2_K15_35, u2_K15_44, u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, 
        u2_K16_19, u2_K16_2, u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, 
        u2_K16_32, u2_K16_35, u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, 
        u2_K16_5, u2_K16_6, u2_K16_7, u2_K16_8, u2_K1_43, u2_K2_1, u2_K2_11, u2_K2_12, u2_K2_13, 
        u2_K2_17, u2_K2_18, u2_K2_2, u2_K2_20, u2_K2_23, u2_K2_24, u2_K2_25, u2_K2_26, u2_K2_29, 
        u2_K2_30, u2_K2_31, u2_K2_35, u2_K2_36, u2_K2_37, u2_K2_38, u2_K2_42, u2_K2_44, u2_K2_47, 
        u2_K2_48, u2_K2_5, u2_K2_6, u2_K2_8, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, 
        u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, 
        u2_K4_6, u2_K4_7, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, 
        u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, 
        u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, 
        u2_K6_13, u2_K6_14, u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, 
        u2_K7_26, u2_K7_30, u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, 
        u2_K7_7, u2_K8_1, u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, u2_K8_19, u2_K8_2, 
        u2_K8_20, u2_K8_47, u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, u2_K9_12, u2_K9_14, 
        u2_K9_23, u2_K9_25, u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_K9_5, u2_R0_1, u2_R0_12, 
        u2_R0_13, u2_R0_16, u2_R0_17, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_29, 
        u2_R0_32, u2_R0_4, u2_R0_5, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_12, u2_R10_13, 
        u2_R10_16, u2_R10_21, u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, 
        u2_R10_9, u2_R11_1, u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, 
        u2_R13_1, u2_R13_12, u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, 
        u2_R13_29, u2_R13_32, u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, 
        u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, 
        u2_R1_31, u2_R1_32, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, 
        u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, 
        u2_R2_25, u2_R2_3, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, 
        u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, 
        u2_R3_24, u2_R3_25, u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, 
        u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, 
        u2_R4_29, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, 
        u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, 
        u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, 
        u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, u2_R6_32, u2_R6_4, 
        u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, 
        u2_R7_16, u2_R7_17, u2_R7_22, u2_R7_24, u2_R7_25, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_4, 
        u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, 
        u2_R8_16, u2_R8_17, u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, 
        u2_R8_29, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_R9_12, u2_R9_13, 
        u2_R9_17, u2_R9_20, u2_R9_32, u2_R9_8, u2_R9_9, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_33, 
        u2_desIn_r_57, u2_key_r_14, u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, u2_u0_X_25, 
        u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, u2_u0_X_37, 
        u2_u0_X_39, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, u2_u10_X_10, 
        u2_u10_X_15, u2_u10_X_16, u2_u10_X_18, u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, 
        u2_u10_X_30, u2_u10_X_32, u2_u10_X_33, u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, 
        u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u10_X_7, 
        u2_u10_X_8, u2_u10_X_9, u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, u2_u11_X_22, u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, 
        u2_u11_X_28, u2_u11_X_29, u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, 
        u2_u11_X_40, u2_u11_X_41, u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, u2_u11_X_6, u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, 
        u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, 
        u2_u12_X_31, u2_u12_X_33, u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, u2_u12_X_39, u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, 
        u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, 
        u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, u2_u13_X_35, u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, 
        u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, 
        u2_u14_X_11, u2_u14_X_13, u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, u2_u14_X_20, u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, 
        u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, 
        u2_u14_X_45, u2_u14_X_46, u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, 
        u2_u15_X_22, u2_u15_X_27, u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, 
        u2_u15_X_46, u2_u15_X_9, u2_u1_X_15, u2_u1_X_16, u2_u1_X_21, u2_u1_X_22, u2_u1_X_27, u2_u1_X_3, u2_u1_X_33, 
        u2_u1_X_34, u2_u1_X_39, u2_u1_X_4, u2_u1_X_40, u2_u1_X_41, u2_u1_X_43, u2_u1_X_45, u2_u1_X_46, u2_u1_X_9, 
        u2_u2_X_15, u2_u2_X_16, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, 
        u2_u2_X_34, u2_u2_X_35, u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, 
        u2_u3_X_33, u2_u3_X_34, u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, 
        u2_u4_X_15, u2_u4_X_16, u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, 
        u2_u4_X_40, u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, 
        u2_u5_X_25, u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, 
        u2_u5_X_39, u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, 
        u2_u6_X_33, u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, 
        u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, u2_u7_X_44, u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, 
        u2_u8_X_1, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u8_X_31, u2_u8_X_32, 
        u2_u8_X_34, u2_u8_X_39, u2_u8_X_40, u2_u8_X_45, u2_u8_X_46, u2_u8_X_47, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, 
        u2_u9_X_21, u2_u9_X_27, u2_u9_X_28, u2_u9_X_29, u2_u9_X_3, u2_u9_X_30, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, 
        u2_u9_X_45, u2_u9_X_46, u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, 
        u2_uk_K_r1_16, u2_uk_K_r1_18, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, 
        u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, 
        u2_uk_K_r3_43, u2_uk_K_r3_9, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, 
        u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_0, u2_uk_K_r7_25, 
        u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, 
        u2_uk_K_r8_37, u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r9_10, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_n1004, u2_uk_n1008, u2_uk_n1020, 
        u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, 
        u2_uk_n1049, u2_uk_n1050, u2_uk_n1053, u2_uk_n1069, u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, 
        u2_uk_n1083, u2_uk_n1084, u2_uk_n1088, u2_uk_n1089, u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1098, u2_uk_n1110, 
        u2_uk_n1113, u2_uk_n1120, u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1132, u2_uk_n1133, u2_uk_n1136, 
        u2_uk_n1137, u2_uk_n1140, u2_uk_n1141, u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, 
        u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, 
        u2_uk_n1293, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, 
        u2_uk_n1310, u2_uk_n1311, u2_uk_n1314, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, 
        u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, 
        u2_uk_n1356, u2_uk_n1359, u2_uk_n1361, u2_uk_n1370, u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, 
        u2_uk_n1410, u2_uk_n1413, u2_uk_n1422, u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, 
        u2_uk_n1440, u2_uk_n1441, u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, 
        u2_uk_n1459, u2_uk_n1462, u2_uk_n1465, u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1488, 
        u2_uk_n1490, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, 
        u2_uk_n1556, u2_uk_n1563, u2_uk_n1568, u2_uk_n1573, u2_uk_n1580, u2_uk_n1585, u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, 
        u2_uk_n1609, u2_uk_n1615, u2_uk_n1622, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n1708, 
        u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1746, u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, 
        u2_uk_n1803, u2_uk_n1807, u2_uk_n1808, u2_uk_n1816, u2_uk_n1817, u2_uk_n1819, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, 
        u2_uk_n1834, u2_uk_n1840, u2_uk_n1846, u2_uk_n1849, u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, 
        u2_uk_n240, u2_uk_n257, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n308, u2_uk_n313, u2_uk_n319, u2_uk_n335, 
        u2_uk_n373, u2_uk_n386, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, 
        u2_uk_n504, u2_uk_n515, u2_uk_n520, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n939, u2_uk_n942, u2_uk_n943, 
        u2_uk_n945, u2_uk_n946, u2_uk_n955, u2_uk_n958, u2_uk_n959, u2_uk_n963, u2_uk_n985, u2_uk_n986, u2_uk_n987, 
        u2_uk_n991, u2_uk_n993, u2_uk_n995, u2_uk_n998, u2_uk_n999 );
  input clk;
  input decrypt;
  input [63:0] desIn;
  input [55:0] key1;
  input [55:0] key2;
  input [55:0] key3;
  output [63:0] desOut;
  input u0_out0_1, u0_out0_10, u0_out0_11, u0_out0_12, u0_out0_13, u0_out0_14, u0_out0_15, u0_out0_16, u0_out0_17, 
        u0_out0_18, u0_out0_19, u0_out0_2, u0_out0_20, u0_out0_21, u0_out0_22, u0_out0_23, u0_out0_24, u0_out0_25, 
        u0_out0_26, u0_out0_27, u0_out0_28, u0_out0_29, u0_out0_3, u0_out0_30, u0_out0_31, u0_out0_32, u0_out0_4, 
        u0_out0_5, u0_out0_6, u0_out0_7, u0_out0_8, u0_out0_9, u0_out10_1, u0_out10_10, u0_out10_11, u0_out10_12, 
        u0_out10_13, u0_out10_14, u0_out10_15, u0_out10_16, u0_out10_17, u0_out10_18, u0_out10_19, u0_out10_2, u0_out10_20, 
        u0_out10_21, u0_out10_22, u0_out10_23, u0_out10_24, u0_out10_25, u0_out10_26, u0_out10_27, u0_out10_28, u0_out10_29, 
        u0_out10_3, u0_out10_30, u0_out10_31, u0_out10_32, u0_out10_4, u0_out10_5, u0_out10_6, u0_out10_7, u0_out10_8, 
        u0_out10_9, u0_out11_1, u0_out11_10, u0_out11_11, u0_out11_12, u0_out11_13, u0_out11_14, u0_out11_15, u0_out11_16, 
        u0_out11_17, u0_out11_18, u0_out11_19, u0_out11_2, u0_out11_20, u0_out11_21, u0_out11_22, u0_out11_23, u0_out11_24, 
        u0_out11_25, u0_out11_26, u0_out11_27, u0_out11_28, u0_out11_29, u0_out11_3, u0_out11_30, u0_out11_31, u0_out11_32, 
        u0_out11_4, u0_out11_5, u0_out11_6, u0_out11_7, u0_out11_8, u0_out11_9, u0_out12_1, u0_out12_10, u0_out12_11, 
        u0_out12_12, u0_out12_13, u0_out12_14, u0_out12_15, u0_out12_16, u0_out12_17, u0_out12_18, u0_out12_19, u0_out12_2, 
        u0_out12_20, u0_out12_21, u0_out12_22, u0_out12_23, u0_out12_24, u0_out12_25, u0_out12_26, u0_out12_27, u0_out12_28, 
        u0_out12_29, u0_out12_3, u0_out12_30, u0_out12_31, u0_out12_32, u0_out12_4, u0_out12_5, u0_out12_6, u0_out12_7, 
        u0_out12_8, u0_out12_9, u0_out13_1, u0_out13_10, u0_out13_11, u0_out13_12, u0_out13_13, u0_out13_14, u0_out13_15, 
        u0_out13_17, u0_out13_18, u0_out13_19, u0_out13_2, u0_out13_20, u0_out13_21, u0_out13_22, u0_out13_23, u0_out13_25, 
        u0_out13_26, u0_out13_27, u0_out13_28, u0_out13_29, u0_out13_3, u0_out13_31, u0_out13_32, u0_out13_4, u0_out13_5, 
        u0_out13_7, u0_out13_8, u0_out13_9, u0_out14_1, u0_out14_10, u0_out14_11, u0_out14_12, u0_out14_13, u0_out14_14, 
        u0_out14_15, u0_out14_16, u0_out14_18, u0_out14_19, u0_out14_2, u0_out14_20, u0_out14_21, u0_out14_22, u0_out14_24, 
        u0_out14_25, u0_out14_26, u0_out14_27, u0_out14_28, u0_out14_29, u0_out14_3, u0_out14_30, u0_out14_32, u0_out14_4, 
        u0_out14_5, u0_out14_6, u0_out14_7, u0_out14_8, u0_out15_1, u0_out15_10, u0_out15_11, u0_out15_12, u0_out15_13, 
        u0_out15_14, u0_out15_15, u0_out15_16, u0_out15_17, u0_out15_18, u0_out15_19, u0_out15_2, u0_out15_20, u0_out15_21, 
        u0_out15_22, u0_out15_23, u0_out15_24, u0_out15_25, u0_out15_26, u0_out15_27, u0_out15_28, u0_out15_29, u0_out15_3, 
        u0_out15_30, u0_out15_31, u0_out15_32, u0_out15_4, u0_out15_5, u0_out15_6, u0_out15_7, u0_out15_8, u0_out15_9, 
        u0_out1_1, u0_out1_10, u0_out1_11, u0_out1_12, u0_out1_13, u0_out1_14, u0_out1_16, u0_out1_17, u0_out1_18, 
        u0_out1_19, u0_out1_2, u0_out1_20, u0_out1_22, u0_out1_23, u0_out1_24, u0_out1_25, u0_out1_26, u0_out1_28, 
        u0_out1_29, u0_out1_3, u0_out1_30, u0_out1_31, u0_out1_32, u0_out1_4, u0_out1_6, u0_out1_7, u0_out1_8, 
        u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_11, u0_out2_12, u0_out2_13, u0_out2_14, u0_out2_15, u0_out2_16, 
        u0_out2_17, u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, u0_out2_21, u0_out2_22, u0_out2_23, u0_out2_24, 
        u0_out2_25, u0_out2_26, u0_out2_27, u0_out2_28, u0_out2_29, u0_out2_3, u0_out2_30, u0_out2_31, u0_out2_32, 
        u0_out2_4, u0_out2_5, u0_out2_6, u0_out2_7, u0_out2_8, u0_out2_9, u0_out3_1, u0_out3_10, u0_out3_11, 
        u0_out3_12, u0_out3_13, u0_out3_14, u0_out3_15, u0_out3_16, u0_out3_17, u0_out3_18, u0_out3_19, u0_out3_2, 
        u0_out3_20, u0_out3_21, u0_out3_22, u0_out3_23, u0_out3_24, u0_out3_25, u0_out3_26, u0_out3_27, u0_out3_28, 
        u0_out3_29, u0_out3_3, u0_out3_30, u0_out3_31, u0_out3_32, u0_out3_4, u0_out3_5, u0_out3_6, u0_out3_7, 
        u0_out3_8, u0_out3_9, u0_out4_1, u0_out4_10, u0_out4_11, u0_out4_13, u0_out4_14, u0_out4_15, u0_out4_16, 
        u0_out4_17, u0_out4_18, u0_out4_19, u0_out4_2, u0_out4_20, u0_out4_21, u0_out4_23, u0_out4_24, u0_out4_25, 
        u0_out4_26, u0_out4_27, u0_out4_28, u0_out4_29, u0_out4_3, u0_out4_30, u0_out4_31, u0_out4_4, u0_out4_5, 
        u0_out4_6, u0_out4_8, u0_out4_9, u0_out5_1, u0_out5_10, u0_out5_11, u0_out5_12, u0_out5_13, u0_out5_14, 
        u0_out5_15, u0_out5_16, u0_out5_17, u0_out5_18, u0_out5_19, u0_out5_2, u0_out5_20, u0_out5_21, u0_out5_22, 
        u0_out5_23, u0_out5_24, u0_out5_25, u0_out5_26, u0_out5_27, u0_out5_28, u0_out5_29, u0_out5_3, u0_out5_30, 
        u0_out5_31, u0_out5_32, u0_out5_4, u0_out5_5, u0_out5_6, u0_out5_7, u0_out5_8, u0_out5_9, u0_out6_1, 
        u0_out6_10, u0_out6_11, u0_out6_13, u0_out6_16, u0_out6_17, u0_out6_18, u0_out6_19, u0_out6_2, u0_out6_20, 
        u0_out6_23, u0_out6_24, u0_out6_26, u0_out6_28, u0_out6_29, u0_out6_30, u0_out6_31, u0_out6_4, u0_out6_6, 
        u0_out6_9, u0_out7_1, u0_out7_10, u0_out7_11, u0_out7_12, u0_out7_13, u0_out7_14, u0_out7_15, u0_out7_16, 
        u0_out7_17, u0_out7_18, u0_out7_19, u0_out7_2, u0_out7_20, u0_out7_21, u0_out7_22, u0_out7_23, u0_out7_24, 
        u0_out7_25, u0_out7_26, u0_out7_27, u0_out7_28, u0_out7_29, u0_out7_3, u0_out7_30, u0_out7_31, u0_out7_32, 
        u0_out7_4, u0_out7_5, u0_out7_6, u0_out7_7, u0_out7_8, u0_out7_9, u0_out8_1, u0_out8_10, u0_out8_11, 
        u0_out8_12, u0_out8_13, u0_out8_14, u0_out8_15, u0_out8_16, u0_out8_17, u0_out8_18, u0_out8_19, u0_out8_2, 
        u0_out8_20, u0_out8_21, u0_out8_22, u0_out8_23, u0_out8_24, u0_out8_25, u0_out8_26, u0_out8_27, u0_out8_28, 
        u0_out8_29, u0_out8_3, u0_out8_30, u0_out8_31, u0_out8_32, u0_out8_4, u0_out8_5, u0_out8_6, u0_out8_7, 
        u0_out8_8, u0_out8_9, u0_out9_1, u0_out9_10, u0_out9_11, u0_out9_12, u0_out9_13, u0_out9_14, u0_out9_15, 
        u0_out9_16, u0_out9_17, u0_out9_18, u0_out9_19, u0_out9_2, u0_out9_20, u0_out9_21, u0_out9_22, u0_out9_23, 
        u0_out9_24, u0_out9_25, u0_out9_26, u0_out9_27, u0_out9_28, u0_out9_29, u0_out9_3, u0_out9_30, u0_out9_31, 
        u0_out9_32, u0_out9_4, u0_out9_5, u0_out9_6, u0_out9_7, u0_out9_8, u0_out9_9, u0_uk_n10, u0_uk_n100, 
        u0_uk_n102, u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n129, u0_uk_n141, 
        u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n162, u0_uk_n163, 
        u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, u0_uk_n191, u0_uk_n202, u0_uk_n203, u0_uk_n207, 
        u0_uk_n208, u0_uk_n209, u0_uk_n213, u0_uk_n214, u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n223, u0_uk_n230, 
        u0_uk_n231, u0_uk_n238, u0_uk_n240, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n27, u0_uk_n31, 
        u0_uk_n60, u0_uk_n63, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u1_out0_1, u1_out0_10, 
        u1_out0_11, u1_out0_12, u1_out0_13, u1_out0_14, u1_out0_15, u1_out0_16, u1_out0_17, u1_out0_18, u1_out0_19, 
        u1_out0_2, u1_out0_20, u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_24, u1_out0_25, u1_out0_26, u1_out0_27, 
        u1_out0_28, u1_out0_29, u1_out0_3, u1_out0_30, u1_out0_31, u1_out0_32, u1_out0_4, u1_out0_5, u1_out0_6, 
        u1_out0_7, u1_out0_8, u1_out0_9, u1_out10_1, u1_out10_10, u1_out10_11, u1_out10_12, u1_out10_13, u1_out10_14, 
        u1_out10_15, u1_out10_16, u1_out10_17, u1_out10_18, u1_out10_19, u1_out10_2, u1_out10_20, u1_out10_21, u1_out10_22, 
        u1_out10_23, u1_out10_24, u1_out10_25, u1_out10_26, u1_out10_27, u1_out10_28, u1_out10_29, u1_out10_3, u1_out10_30, 
        u1_out10_31, u1_out10_32, u1_out10_4, u1_out10_5, u1_out10_6, u1_out10_7, u1_out10_8, u1_out10_9, u1_out11_1, 
        u1_out11_10, u1_out11_11, u1_out11_12, u1_out11_13, u1_out11_14, u1_out11_15, u1_out11_16, u1_out11_17, u1_out11_18, 
        u1_out11_19, u1_out11_2, u1_out11_20, u1_out11_21, u1_out11_22, u1_out11_23, u1_out11_24, u1_out11_25, u1_out11_26, 
        u1_out11_27, u1_out11_28, u1_out11_29, u1_out11_3, u1_out11_30, u1_out11_31, u1_out11_32, u1_out11_4, u1_out11_5, 
        u1_out11_6, u1_out11_7, u1_out11_8, u1_out11_9, u1_out12_1, u1_out12_10, u1_out12_11, u1_out12_12, u1_out12_13, 
        u1_out12_14, u1_out12_15, u1_out12_16, u1_out12_17, u1_out12_18, u1_out12_19, u1_out12_2, u1_out12_20, u1_out12_21, 
        u1_out12_22, u1_out12_23, u1_out12_24, u1_out12_25, u1_out12_26, u1_out12_27, u1_out12_28, u1_out12_29, u1_out12_3, 
        u1_out12_30, u1_out12_31, u1_out12_32, u1_out12_4, u1_out12_5, u1_out12_6, u1_out12_7, u1_out12_8, u1_out12_9, 
        u1_out13_1, u1_out13_10, u1_out13_11, u1_out13_12, u1_out13_13, u1_out13_14, u1_out13_15, u1_out13_16, u1_out13_17, 
        u1_out13_18, u1_out13_19, u1_out13_2, u1_out13_20, u1_out13_21, u1_out13_22, u1_out13_23, u1_out13_24, u1_out13_25, 
        u1_out13_26, u1_out13_27, u1_out13_28, u1_out13_29, u1_out13_3, u1_out13_30, u1_out13_31, u1_out13_32, u1_out13_4, 
        u1_out13_5, u1_out13_6, u1_out13_7, u1_out13_8, u1_out13_9, u1_out14_1, u1_out14_10, u1_out14_11, u1_out14_12, 
        u1_out14_13, u1_out14_14, u1_out14_15, u1_out14_16, u1_out14_17, u1_out14_18, u1_out14_19, u1_out14_2, u1_out14_20, 
        u1_out14_21, u1_out14_22, u1_out14_23, u1_out14_24, u1_out14_25, u1_out14_26, u1_out14_27, u1_out14_28, u1_out14_29, 
        u1_out14_3, u1_out14_30, u1_out14_31, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, u1_out14_8, 
        u1_out14_9, u1_out15_1, u1_out15_10, u1_out15_11, u1_out15_12, u1_out15_13, u1_out15_14, u1_out15_15, u1_out15_16, 
        u1_out15_17, u1_out15_18, u1_out15_19, u1_out15_2, u1_out15_20, u1_out15_21, u1_out15_22, u1_out15_23, u1_out15_24, 
        u1_out15_25, u1_out15_26, u1_out15_27, u1_out15_28, u1_out15_29, u1_out15_3, u1_out15_30, u1_out15_31, u1_out15_32, 
        u1_out15_4, u1_out15_5, u1_out15_6, u1_out15_7, u1_out15_8, u1_out15_9, u1_out1_1, u1_out1_10, u1_out1_11, 
        u1_out1_12, u1_out1_13, u1_out1_14, u1_out1_15, u1_out1_16, u1_out1_17, u1_out1_18, u1_out1_19, u1_out1_2, 
        u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_23, u1_out1_24, u1_out1_25, u1_out1_26, u1_out1_27, u1_out1_28, 
        u1_out1_29, u1_out1_3, u1_out1_30, u1_out1_31, u1_out1_32, u1_out1_4, u1_out1_5, u1_out1_6, u1_out1_7, 
        u1_out1_8, u1_out1_9, u1_out2_1, u1_out2_10, u1_out2_11, u1_out2_12, u1_out2_13, u1_out2_14, u1_out2_15, 
        u1_out2_16, u1_out2_17, u1_out2_18, u1_out2_19, u1_out2_2, u1_out2_20, u1_out2_21, u1_out2_22, u1_out2_23, 
        u1_out2_24, u1_out2_25, u1_out2_26, u1_out2_27, u1_out2_28, u1_out2_29, u1_out2_3, u1_out2_30, u1_out2_31, 
        u1_out2_32, u1_out2_4, u1_out2_5, u1_out2_6, u1_out2_7, u1_out2_8, u1_out2_9, u1_out3_1, u1_out3_10, 
        u1_out3_11, u1_out3_12, u1_out3_13, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_17, u1_out3_18, u1_out3_19, 
        u1_out3_2, u1_out3_20, u1_out3_21, u1_out3_22, u1_out3_23, u1_out3_24, u1_out3_25, u1_out3_26, u1_out3_27, 
        u1_out3_28, u1_out3_29, u1_out3_3, u1_out3_30, u1_out3_31, u1_out3_32, u1_out3_4, u1_out3_5, u1_out3_6, 
        u1_out3_7, u1_out3_8, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_11, u1_out4_12, u1_out4_13, u1_out4_14, 
        u1_out4_15, u1_out4_16, u1_out4_17, u1_out4_18, u1_out4_19, u1_out4_2, u1_out4_20, u1_out4_21, u1_out4_22, 
        u1_out4_23, u1_out4_24, u1_out4_25, u1_out4_26, u1_out4_27, u1_out4_28, u1_out4_29, u1_out4_3, u1_out4_30, 
        u1_out4_31, u1_out4_32, u1_out4_4, u1_out4_5, u1_out4_6, u1_out4_7, u1_out4_8, u1_out4_9, u1_out5_1, 
        u1_out5_10, u1_out5_11, u1_out5_12, u1_out5_13, u1_out5_14, u1_out5_15, u1_out5_16, u1_out5_17, u1_out5_18, 
        u1_out5_19, u1_out5_2, u1_out5_20, u1_out5_21, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_25, u1_out5_26, 
        u1_out5_27, u1_out5_28, u1_out5_29, u1_out5_3, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_4, u1_out5_5, 
        u1_out5_6, u1_out5_7, u1_out5_8, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_11, u1_out6_12, u1_out6_13, 
        u1_out6_14, u1_out6_15, u1_out6_16, u1_out6_17, u1_out6_18, u1_out6_19, u1_out6_2, u1_out6_20, u1_out6_21, 
        u1_out6_22, u1_out6_23, u1_out6_24, u1_out6_25, u1_out6_26, u1_out6_27, u1_out6_28, u1_out6_29, u1_out6_3, 
        u1_out6_30, u1_out6_31, u1_out6_32, u1_out6_4, u1_out6_5, u1_out6_6, u1_out6_7, u1_out6_8, u1_out6_9, 
        u1_out7_1, u1_out7_10, u1_out7_11, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_15, u1_out7_16, u1_out7_17, 
        u1_out7_18, u1_out7_19, u1_out7_2, u1_out7_20, u1_out7_21, u1_out7_22, u1_out7_23, u1_out7_24, u1_out7_25, 
        u1_out7_26, u1_out7_27, u1_out7_28, u1_out7_29, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, u1_out7_4, 
        u1_out7_5, u1_out7_6, u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_11, u1_out8_12, 
        u1_out8_13, u1_out8_14, u1_out8_15, u1_out8_16, u1_out8_17, u1_out8_18, u1_out8_19, u1_out8_2, u1_out8_20, 
        u1_out8_21, u1_out8_22, u1_out8_23, u1_out8_24, u1_out8_25, u1_out8_26, u1_out8_27, u1_out8_28, u1_out8_29, 
        u1_out8_3, u1_out8_30, u1_out8_31, u1_out8_32, u1_out8_4, u1_out8_5, u1_out8_6, u1_out8_7, u1_out8_8, 
        u1_out8_9, u1_out9_1, u1_out9_10, u1_out9_11, u1_out9_12, u1_out9_13, u1_out9_14, u1_out9_15, u1_out9_16, 
        u1_out9_17, u1_out9_18, u1_out9_19, u1_out9_2, u1_out9_20, u1_out9_21, u1_out9_22, u1_out9_23, u1_out9_24, 
        u1_out9_25, u1_out9_26, u1_out9_27, u1_out9_28, u1_out9_29, u1_out9_3, u1_out9_30, u1_out9_31, u1_out9_32, 
        u1_out9_4, u1_out9_5, u1_out9_6, u1_out9_7, u1_out9_8, u1_out9_9, u2_out0_11, u2_out0_12, u2_out0_13, 
        u2_out0_14, u2_out0_15, u2_out0_18, u2_out0_19, u2_out0_2, u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_27, 
        u2_out0_28, u2_out0_29, u2_out0_3, u2_out0_32, u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, u2_out10_1, 
        u2_out10_10, u2_out10_11, u2_out10_12, u2_out10_13, u2_out10_14, u2_out10_15, u2_out10_16, u2_out10_18, u2_out10_19, 
        u2_out10_2, u2_out10_20, u2_out10_21, u2_out10_22, u2_out10_24, u2_out10_25, u2_out10_26, u2_out10_27, u2_out10_28, 
        u2_out10_29, u2_out10_3, u2_out10_30, u2_out10_32, u2_out10_4, u2_out10_5, u2_out10_6, u2_out10_7, u2_out10_8, 
        u2_out11_1, u2_out11_10, u2_out11_11, u2_out11_12, u2_out11_13, u2_out11_14, u2_out11_15, u2_out11_16, u2_out11_17, 
        u2_out11_18, u2_out11_19, u2_out11_2, u2_out11_20, u2_out11_21, u2_out11_22, u2_out11_23, u2_out11_24, u2_out11_25, 
        u2_out11_26, u2_out11_27, u2_out11_28, u2_out11_29, u2_out11_3, u2_out11_30, u2_out11_31, u2_out11_32, u2_out11_4, 
        u2_out11_5, u2_out11_6, u2_out11_7, u2_out11_8, u2_out11_9, u2_out12_11, u2_out12_12, u2_out12_13, u2_out12_14, 
        u2_out12_15, u2_out12_17, u2_out12_18, u2_out12_19, u2_out12_2, u2_out12_21, u2_out12_22, u2_out12_23, u2_out12_25, 
        u2_out12_27, u2_out12_28, u2_out12_29, u2_out12_3, u2_out12_31, u2_out12_32, u2_out12_4, u2_out12_5, u2_out12_7, 
        u2_out12_8, u2_out12_9, u2_out13_11, u2_out13_12, u2_out13_14, u2_out13_15, u2_out13_19, u2_out13_21, u2_out13_22, 
        u2_out13_25, u2_out13_27, u2_out13_29, u2_out13_3, u2_out13_32, u2_out13_4, u2_out13_5, u2_out13_7, u2_out13_8, 
        u2_out14_1, u2_out14_10, u2_out14_11, u2_out14_12, u2_out14_13, u2_out14_14, u2_out14_15, u2_out14_16, u2_out14_17, 
        u2_out14_18, u2_out14_19, u2_out14_2, u2_out14_20, u2_out14_21, u2_out14_22, u2_out14_23, u2_out14_24, u2_out14_25, 
        u2_out14_26, u2_out14_27, u2_out14_28, u2_out14_29, u2_out14_3, u2_out14_30, u2_out14_31, u2_out14_32, u2_out14_4, 
        u2_out14_5, u2_out14_6, u2_out14_7, u2_out14_8, u2_out14_9, u2_out15_1, u2_out15_10, u2_out15_11, u2_out15_12, 
        u2_out15_13, u2_out15_14, u2_out15_15, u2_out15_16, u2_out15_17, u2_out15_18, u2_out15_19, u2_out15_2, u2_out15_20, 
        u2_out15_21, u2_out15_22, u2_out15_23, u2_out15_24, u2_out15_25, u2_out15_26, u2_out15_27, u2_out15_28, u2_out15_29, 
        u2_out15_3, u2_out15_30, u2_out15_31, u2_out15_32, u2_out15_4, u2_out15_5, u2_out15_6, u2_out15_7, u2_out15_8, 
        u2_out15_9, u2_out1_1, u2_out1_10, u2_out1_11, u2_out1_12, u2_out1_13, u2_out1_14, u2_out1_15, u2_out1_16, 
        u2_out1_17, u2_out1_18, u2_out1_19, u2_out1_2, u2_out1_20, u2_out1_21, u2_out1_22, u2_out1_23, u2_out1_24, 
        u2_out1_25, u2_out1_26, u2_out1_27, u2_out1_28, u2_out1_29, u2_out1_3, u2_out1_30, u2_out1_31, u2_out1_32, 
        u2_out1_4, u2_out1_5, u2_out1_6, u2_out1_7, u2_out1_8, u2_out1_9, u2_out2_1, u2_out2_10, u2_out2_11, 
        u2_out2_12, u2_out2_13, u2_out2_14, u2_out2_15, u2_out2_16, u2_out2_17, u2_out2_18, u2_out2_19, u2_out2_2, 
        u2_out2_20, u2_out2_21, u2_out2_22, u2_out2_23, u2_out2_24, u2_out2_25, u2_out2_26, u2_out2_27, u2_out2_28, 
        u2_out2_29, u2_out2_3, u2_out2_30, u2_out2_31, u2_out2_32, u2_out2_4, u2_out2_5, u2_out2_6, u2_out2_7, 
        u2_out2_8, u2_out2_9, u2_out3_1, u2_out3_10, u2_out3_11, u2_out3_13, u2_out3_14, u2_out3_15, u2_out3_16, 
        u2_out3_17, u2_out3_18, u2_out3_19, u2_out3_2, u2_out3_20, u2_out3_21, u2_out3_23, u2_out3_24, u2_out3_25, 
        u2_out3_26, u2_out3_27, u2_out3_28, u2_out3_29, u2_out3_3, u2_out3_30, u2_out3_31, u2_out3_4, u2_out3_5, 
        u2_out3_6, u2_out3_8, u2_out3_9, u2_out4_1, u2_out4_10, u2_out4_11, u2_out4_12, u2_out4_13, u2_out4_14, 
        u2_out4_15, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_19, u2_out4_2, u2_out4_20, u2_out4_21, u2_out4_22, 
        u2_out4_23, u2_out4_24, u2_out4_25, u2_out4_26, u2_out4_27, u2_out4_28, u2_out4_29, u2_out4_3, u2_out4_30, 
        u2_out4_31, u2_out4_32, u2_out4_4, u2_out4_5, u2_out4_6, u2_out4_7, u2_out4_8, u2_out4_9, u2_out5_1, 
        u2_out5_10, u2_out5_11, u2_out5_12, u2_out5_13, u2_out5_14, u2_out5_15, u2_out5_16, u2_out5_17, u2_out5_18, 
        u2_out5_19, u2_out5_2, u2_out5_20, u2_out5_21, u2_out5_22, u2_out5_23, u2_out5_24, u2_out5_25, u2_out5_26, 
        u2_out5_27, u2_out5_28, u2_out5_29, u2_out5_3, u2_out5_30, u2_out5_31, u2_out5_32, u2_out5_4, u2_out5_5, 
        u2_out5_6, u2_out5_7, u2_out5_8, u2_out5_9, u2_out6_1, u2_out6_10, u2_out6_11, u2_out6_12, u2_out6_13, 
        u2_out6_14, u2_out6_15, u2_out6_16, u2_out6_17, u2_out6_18, u2_out6_19, u2_out6_2, u2_out6_20, u2_out6_21, 
        u2_out6_22, u2_out6_23, u2_out6_24, u2_out6_25, u2_out6_26, u2_out6_27, u2_out6_28, u2_out6_29, u2_out6_3, 
        u2_out6_30, u2_out6_31, u2_out6_32, u2_out6_4, u2_out6_5, u2_out6_6, u2_out6_7, u2_out6_8, u2_out6_9, 
        u2_out7_1, u2_out7_10, u2_out7_13, u2_out7_15, u2_out7_16, u2_out7_17, u2_out7_18, u2_out7_2, u2_out7_20, 
        u2_out7_21, u2_out7_23, u2_out7_24, u2_out7_26, u2_out7_27, u2_out7_28, u2_out7_30, u2_out7_31, u2_out7_5, 
        u2_out7_6, u2_out7_9, u2_out8_1, u2_out8_10, u2_out8_11, u2_out8_12, u2_out8_13, u2_out8_14, u2_out8_15, 
        u2_out8_16, u2_out8_17, u2_out8_18, u2_out8_19, u2_out8_2, u2_out8_20, u2_out8_21, u2_out8_22, u2_out8_23, 
        u2_out8_24, u2_out8_25, u2_out8_26, u2_out8_27, u2_out8_28, u2_out8_29, u2_out8_3, u2_out8_30, u2_out8_31, 
        u2_out8_32, u2_out8_4, u2_out8_5, u2_out8_6, u2_out8_7, u2_out8_8, u2_out8_9, u2_out9_1, u2_out9_10, 
        u2_out9_11, u2_out9_12, u2_out9_13, u2_out9_14, u2_out9_15, u2_out9_16, u2_out9_17, u2_out9_18, u2_out9_19, 
        u2_out9_2, u2_out9_20, u2_out9_21, u2_out9_22, u2_out9_23, u2_out9_24, u2_out9_25, u2_out9_26, u2_out9_27, 
        u2_out9_28, u2_out9_29, u2_out9_3, u2_out9_30, u2_out9_31, u2_out9_32, u2_out9_4, u2_out9_5, u2_out9_6, 
        u2_out9_7, u2_out9_8, u2_out9_9, u2_uk_n10, u2_uk_n100, u2_uk_n102, u2_uk_n109, u2_uk_n11, u2_uk_n110, 
        u2_uk_n117, u2_uk_n118, u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, 
        u2_uk_n148, u2_uk_n155, u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n164, u2_uk_n17, u2_uk_n182, u2_uk_n187, 
        u2_uk_n188, u2_uk_n191, u2_uk_n202, u2_uk_n203, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, 
        u2_uk_n217, u2_uk_n220, u2_uk_n222, u2_uk_n223, u2_uk_n230, u2_uk_n231, u2_uk_n27, u2_uk_n31, u2_uk_n60, 
        u2_uk_n63, u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n94, u2_uk_n99;
  output u0_FP_33, u0_FP_34, u0_FP_36, u0_FP_37, u0_FP_39, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, 
        u0_FP_45, u0_FP_46, u0_FP_48, u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_FP_55, 
        u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, u0_FP_60, u0_FP_63, u0_FP_64, u0_K10_1, u0_K10_14, 
        u0_K10_17, u0_K10_18, u0_K10_19, u0_K10_20, u0_K10_32, u0_K11_37, u0_K11_42, u0_K11_48, u0_K12_19, 
        u0_K12_25, u0_K12_35, u0_K12_36, u0_K12_48, u0_K12_5, u0_K12_7, u0_K12_8, u0_K13_41, u0_K14_23, 
        u0_K14_24, u0_K14_25, u0_K14_26, u0_K14_29, u0_K14_5, u0_K14_7, u0_K15_13, u0_K16_18, u0_K16_19, 
        u0_K16_24, u0_K16_26, u0_K16_36, u0_K16_38, u0_K16_5, u0_K16_8, u0_K1_13, u0_K1_14, u0_K1_17, 
        u0_K1_30, u0_K1_31, u0_K2_11, u0_K2_12, u0_K2_18, u0_K2_20, u0_K2_29, u0_K2_30, u0_K2_31, 
        u0_K2_5, u0_K3_12, u0_K3_13, u0_K3_14, u0_K3_17, u0_K3_18, u0_K3_19, u0_K3_23, u0_K3_5, 
        u0_K3_6, u0_K4_36, u0_K4_43, u0_K4_48, u0_K4_6, u0_K5_1, u0_K5_18, u0_K5_24, u0_K5_26, 
        u0_K5_29, u0_K5_31, u0_K5_47, u0_K5_8, u0_K6_11, u0_K6_13, u0_K6_19, u0_K6_20, u0_K6_23, 
        u0_K6_24, u0_K6_41, u0_K8_11, u0_K8_13, u0_K8_19, u0_K9_12, u0_K9_13, u0_K9_14, u0_K9_30, 
        u0_K9_32, u0_K9_44, u0_K9_6, u0_R0_1, u0_R0_13, u0_R0_15, u0_R0_18, u0_R0_19, u0_R0_20, 
        u0_R0_21, u0_R0_28, u0_R0_32, u0_R0_4, u0_R0_7, u0_R0_8, u0_R0_9, u0_R10_1, u0_R10_12, 
        u0_R10_14, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_2, u0_R10_20, u0_R10_21, u0_R10_24, 
        u0_R10_25, u0_R10_28, u0_R10_29, u0_R10_3, u0_R10_4, u0_R10_5, u0_R11_10, u0_R11_11, u0_R11_12, 
        u0_R11_13, u0_R11_14, u0_R11_15, u0_R11_16, u0_R11_2, u0_R11_20, u0_R11_28, u0_R11_3, u0_R11_32, 
        u0_R11_5, u0_R11_6, u0_R12_16, u0_R12_17, u0_R12_19, u0_R12_20, u0_R12_22, u0_R12_23, u0_R12_24, 
        u0_R12_30, u0_R12_4, u0_R13_17, u0_R13_18, u0_R13_19, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, 
        u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, u0_R13_28, u0_R13_29, u0_R13_30, u0_R13_31, u0_R13_8, 
        u0_R1_1, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, u0_R1_19, u0_R1_20, u0_R1_21, 
        u0_R1_22, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_3, u0_R1_30, 
        u0_R1_32, u0_R1_4, u0_R1_5, u0_R1_8, u0_R1_9, u0_R2_1, u0_R2_10, u0_R2_11, u0_R2_12, 
        u0_R2_13, u0_R2_14, u0_R2_16, u0_R2_2, u0_R2_21, u0_R2_22, u0_R2_25, u0_R2_28, u0_R2_3, 
        u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_13, u0_R3_15, 
        u0_R3_17, u0_R3_18, u0_R3_20, u0_R3_22, u0_R3_24, u0_R3_25, u0_R3_32, u0_R3_5, u0_R4_1, 
        u0_R4_12, u0_R4_13, u0_R4_16, u0_R4_17, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_22, u0_R4_24, 
        u0_R4_25, u0_R4_26, u0_R4_27, u0_R4_28, u0_R4_29, u0_R4_3, u0_R4_30, u0_R4_32, u0_R4_4, 
        u0_R4_5, u0_R4_8, u0_R4_9, u0_R5_12, u0_R5_13, u0_R5_2, u0_R5_25, u0_R5_3, u0_R5_32, 
        u0_R5_4, u0_R5_5, u0_R5_7, u0_R5_8, u0_R5_9, u0_R6_10, u0_R6_11, u0_R6_12, u0_R6_13, 
        u0_R6_14, u0_R6_17, u0_R6_24, u0_R6_26, u0_R6_28, u0_R6_29, u0_R6_4, u0_R6_5, u0_R6_7, 
        u0_R6_8, u0_R6_9, u0_R7_1, u0_R7_12, u0_R7_14, u0_R7_17, u0_R7_20, u0_R7_21, u0_R7_22, 
        u0_R7_23, u0_R7_24, u0_R7_25, u0_R7_28, u0_R7_29, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_8, 
        u0_R7_9, u0_R8_1, u0_R8_12, u0_R8_13, u0_R8_17, u0_R8_19, u0_R8_20, u0_R8_21, u0_R8_22, 
        u0_R8_27, u0_R8_29, u0_R8_30, u0_R8_32, u0_R8_5, u0_R8_6, u0_R8_9, u0_R9_1, u0_R9_10, 
        u0_R9_11, u0_R9_12, u0_R9_13, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_2, u0_R9_20, 
        u0_R9_21, u0_R9_22, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_29, u0_R9_3, u0_R9_30, 
        u0_R9_31, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_desIn_r_1, 
        u0_desIn_r_11, u0_desIn_r_15, u0_desIn_r_17, u0_desIn_r_23, u0_desIn_r_25, u0_desIn_r_27, u0_desIn_r_29, u0_desIn_r_3, u0_desIn_r_31, 
        u0_desIn_r_35, u0_desIn_r_37, u0_desIn_r_39, u0_desIn_r_47, u0_desIn_r_5, u0_desIn_r_51, u0_desIn_r_55, u0_desIn_r_57, u0_desIn_r_59, 
        u0_desIn_r_63, u0_desIn_r_7, u0_desIn_r_9, u0_key_r_0, u0_key_r_11, u0_key_r_12, u0_key_r_13, u0_key_r_14, u0_key_r_16, 
        u0_key_r_19, u0_key_r_2, u0_key_r_20, u0_key_r_21, u0_key_r_22, u0_key_r_23, u0_key_r_28, u0_key_r_29, u0_key_r_30, 
        u0_key_r_35, u0_key_r_4, u0_key_r_41, u0_key_r_42, u0_key_r_47, u0_key_r_48, u0_key_r_5, u0_key_r_50, u0_key_r_54, 
        u0_key_r_55, u0_key_r_6, u0_key_r_9, u0_u0_X_15, u0_u0_X_16, u0_u0_X_21, u0_u0_X_22, u0_u0_X_23, u0_u0_X_25, 
        u0_u0_X_28, u0_u0_X_33, u0_u0_X_42, u0_u0_X_44, u0_u0_X_45, u0_u0_X_46, u0_u10_X_21, u0_u10_X_22, u0_u10_X_34, 
        u0_u10_X_41, u0_u10_X_43, u0_u11_X_1, u0_u11_X_10, u0_u11_X_11, u0_u11_X_12, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, 
        u0_u11_X_16, u0_u11_X_18, u0_u11_X_20, u0_u11_X_22, u0_u11_X_33, u0_u11_X_34, u0_u11_X_39, u0_u11_X_40, u0_u11_X_45, 
        u0_u11_X_46, u0_u11_X_47, u0_u11_X_9, u0_u12_X_10, u0_u12_X_11, u0_u12_X_12, u0_u12_X_13, u0_u12_X_14, u0_u12_X_2, 
        u0_u12_X_24, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_30, u0_u12_X_32, u0_u12_X_33, u0_u12_X_34, u0_u12_X_35, 
        u0_u12_X_36, u0_u12_X_37, u0_u12_X_38, u0_u12_X_39, u0_u12_X_40, u0_u12_X_42, u0_u12_X_44, u0_u12_X_45, u0_u12_X_46, 
        u0_u12_X_48, u0_u12_X_5, u0_u12_X_7, u0_u13_X_1, u0_u13_X_10, u0_u13_X_11, u0_u13_X_12, u0_u13_X_19, u0_u13_X_2, 
        u0_u13_X_20, u0_u13_X_21, u0_u13_X_22, u0_u13_X_27, u0_u13_X_3, u0_u13_X_30, u0_u13_X_32, u0_u13_X_36, u0_u13_X_38, 
        u0_u13_X_39, u0_u13_X_4, u0_u13_X_40, u0_u13_X_41, u0_u13_X_42, u0_u13_X_43, u0_u13_X_44, u0_u13_X_46, u0_u13_X_47, 
        u0_u13_X_48, u0_u13_X_6, u0_u13_X_8, u0_u13_X_9, u0_u14_X_10, u0_u14_X_12, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, 
        u0_u14_X_17, u0_u14_X_18, u0_u14_X_19, u0_u14_X_20, u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_25, 
        u0_u14_X_47, u0_u14_X_48, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u15_X_11, u0_u15_X_13, u0_u15_X_22, u0_u15_X_33, 
        u0_u15_X_4, u0_u15_X_42, u0_u15_X_44, u0_u15_X_45, u0_u15_X_9, u0_u1_X_15, u0_u1_X_16, u0_u1_X_17, u0_u1_X_19, 
        u0_u1_X_21, u0_u1_X_23, u0_u1_X_24, u0_u1_X_25, u0_u1_X_26, u0_u1_X_3, u0_u1_X_33, u0_u1_X_34, u0_u1_X_35, 
        u0_u1_X_36, u0_u1_X_37, u0_u1_X_38, u0_u1_X_39, u0_u1_X_4, u0_u1_X_40, u0_u1_X_42, u0_u1_X_6, u0_u1_X_8, 
        u0_u1_X_9, u0_u2_X_10, u0_u2_X_15, u0_u2_X_16, u0_u2_X_24, u0_u2_X_26, u0_u2_X_27, u0_u2_X_3, u0_u2_X_34, 
        u0_u2_X_46, u0_u2_X_9, u0_u3_X_22, u0_u3_X_24, u0_u3_X_26, u0_u3_X_27, u0_u3_X_28, u0_u3_X_29, u0_u3_X_31, 
        u0_u3_X_34, u0_u3_X_35, u0_u3_X_37, u0_u3_X_39, u0_u3_X_40, u0_u3_X_42, u0_u3_X_44, u0_u3_X_45, u0_u3_X_46, 
        u0_u4_X_10, u0_u4_X_11, u0_u4_X_12, u0_u4_X_13, u0_u4_X_14, u0_u4_X_15, u0_u4_X_16, u0_u4_X_17, u0_u4_X_19, 
        u0_u4_X_2, u0_u4_X_21, u0_u4_X_23, u0_u4_X_25, u0_u4_X_28, u0_u4_X_3, u0_u4_X_30, u0_u4_X_32, u0_u4_X_34, 
        u0_u4_X_4, u0_u4_X_43, u0_u4_X_44, u0_u4_X_45, u0_u4_X_46, u0_u4_X_48, u0_u4_X_5, u0_u4_X_7, u0_u4_X_9, 
        u0_u5_X_10, u0_u5_X_15, u0_u5_X_16, u0_u5_X_21, u0_u5_X_22, u0_u5_X_27, u0_u5_X_3, u0_u5_X_34, u0_u5_X_46, 
        u0_u5_X_9, u0_u6_X_15, u0_u6_X_16, u0_u6_X_2, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, u0_u6_X_31, 
        u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, u0_u6_X_9, u0_u7_X_1, u0_u7_X_2, u0_u7_X_22, u0_u7_X_23, 
        u0_u7_X_25, u0_u7_X_27, u0_u7_X_28, u0_u7_X_29, u0_u7_X_3, u0_u7_X_30, u0_u7_X_31, u0_u7_X_32, u0_u7_X_33, 
        u0_u7_X_34, u0_u7_X_36, u0_u7_X_38, u0_u7_X_4, u0_u7_X_40, u0_u7_X_45, u0_u7_X_46, u0_u7_X_47, u0_u7_X_48, 
        u0_u7_X_9, u0_u8_X_10, u0_u8_X_15, u0_u8_X_16, u0_u8_X_18, u0_u8_X_20, u0_u8_X_22, u0_u8_X_23, u0_u8_X_25, 
        u0_u8_X_27, u0_u8_X_28, u0_u8_X_3, u0_u8_X_39, u0_u8_X_4, u0_u8_X_40, u0_u8_X_45, u0_u8_X_46, u0_u8_X_9, 
        u0_u9_X_10, u0_u9_X_11, u0_u9_X_13, u0_u9_X_15, u0_u9_X_16, u0_u9_X_21, u0_u9_X_22, u0_u9_X_23, u0_u9_X_25, 
        u0_u9_X_27, u0_u9_X_3, u0_u9_X_34, u0_u9_X_35, u0_u9_X_36, u0_u9_X_37, u0_u9_X_38, u0_u9_X_39, u0_u9_X_4, 
        u0_u9_X_41, u0_u9_X_43, u0_u9_X_46, u0_u9_X_5, u0_u9_X_7, u0_uk_K_r0_15, u0_uk_K_r0_28, u0_uk_K_r0_36, u0_uk_K_r0_49, 
        u0_uk_K_r0_7, u0_uk_K_r10_10, u0_uk_K_r10_18, u0_uk_K_r10_23, u0_uk_K_r10_27, u0_uk_K_r10_28, u0_uk_K_r10_32, u0_uk_K_r10_37, u0_uk_K_r10_41, 
        u0_uk_K_r10_42, u0_uk_K_r10_44, u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_20, u0_uk_K_r11_24, u0_uk_K_r11_25, u0_uk_K_r11_27, u0_uk_K_r11_29, 
        u0_uk_K_r11_33, u0_uk_K_r11_39, u0_uk_K_r11_4, u0_uk_K_r12_16, u0_uk_K_r13_0, u0_uk_K_r13_25, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r14_10, 
        u0_uk_K_r14_11, u0_uk_K_r14_12, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_18, u0_uk_K_r14_2, u0_uk_K_r14_45, u0_uk_K_r14_50, u0_uk_K_r14_8, 
        u0_uk_K_r14_9, u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_44, u0_uk_K_r1_7, u0_uk_K_r2_13, u0_uk_K_r2_18, u0_uk_K_r2_20, 
        u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_28, u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, u0_uk_K_r2_50, 
        u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_10, u0_uk_K_r3_14, u0_uk_K_r4_0, u0_uk_K_r4_23, u0_uk_K_r4_33, u0_uk_K_r4_35, u0_uk_K_r4_38, 
        u0_uk_K_r4_41, u0_uk_K_r4_47, u0_uk_K_r5_10, u0_uk_K_r5_17, u0_uk_K_r5_39, u0_uk_K_r5_4, u0_uk_K_r6_0, u0_uk_K_r6_22, u0_uk_K_r6_26, 
        u0_uk_K_r6_31, u0_uk_K_r6_34, u0_uk_K_r6_46, u0_uk_K_r7_26, u0_uk_K_r8_16, u0_uk_K_r8_40, u0_uk_K_r8_41, u0_uk_K_r9_0, u0_uk_K_r9_1, 
        u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_25, u0_uk_K_r9_27, u0_uk_K_r9_30, u0_uk_K_r9_33, u0_uk_K_r9_35, u0_uk_K_r9_45, u0_uk_K_r9_6, 
        u0_uk_K_r9_7, u0_uk_K_r9_9, u0_uk_n1000, u0_uk_n1001, u0_uk_n1002, u0_uk_n1004, u0_uk_n1005, u0_uk_n1006, u0_uk_n101, 
        u0_uk_n1012, u0_uk_n1024, u0_uk_n106, u0_uk_n107, u0_uk_n108, u0_uk_n113, u0_uk_n115, u0_uk_n116, u0_uk_n12, 
        u0_uk_n121, u0_uk_n122, u0_uk_n123, u0_uk_n126, u0_uk_n127, u0_uk_n13, u0_uk_n131, u0_uk_n139, u0_uk_n143, 
        u0_uk_n144, u0_uk_n151, u0_uk_n153, u0_uk_n156, u0_uk_n167, u0_uk_n168, u0_uk_n171, u0_uk_n172, u0_uk_n173, 
        u0_uk_n174, u0_uk_n177, u0_uk_n178, u0_uk_n179, u0_uk_n18, u0_uk_n180, u0_uk_n181, u0_uk_n183, u0_uk_n184, 
        u0_uk_n185, u0_uk_n189, u0_uk_n190, u0_uk_n192, u0_uk_n193, u0_uk_n195, u0_uk_n196, u0_uk_n197, u0_uk_n198, 
        u0_uk_n199, u0_uk_n200, u0_uk_n201, u0_uk_n204, u0_uk_n205, u0_uk_n206, u0_uk_n21, u0_uk_n210, u0_uk_n211, 
        u0_uk_n212, u0_uk_n215, u0_uk_n216, u0_uk_n218, u0_uk_n219, u0_uk_n22, u0_uk_n221, u0_uk_n224, u0_uk_n225, 
        u0_uk_n23, u0_uk_n232, u0_uk_n233, u0_uk_n239, u0_uk_n241, u0_uk_n243, u0_uk_n244, u0_uk_n248, u0_uk_n249, 
        u0_uk_n253, u0_uk_n257, u0_uk_n259, u0_uk_n260, u0_uk_n261, u0_uk_n264, u0_uk_n266, u0_uk_n267, u0_uk_n269, 
        u0_uk_n272, u0_uk_n275, u0_uk_n276, u0_uk_n278, u0_uk_n28, u0_uk_n282, u0_uk_n283, u0_uk_n285, u0_uk_n289, 
        u0_uk_n290, u0_uk_n293, u0_uk_n3, u0_uk_n300, u0_uk_n307, u0_uk_n310, u0_uk_n314, u0_uk_n316, u0_uk_n318, 
        u0_uk_n32, u0_uk_n320, u0_uk_n324, u0_uk_n329, u0_uk_n33, u0_uk_n330, u0_uk_n331, u0_uk_n332, u0_uk_n336, 
        u0_uk_n337, u0_uk_n339, u0_uk_n341, u0_uk_n344, u0_uk_n347, u0_uk_n348, u0_uk_n352, u0_uk_n355, u0_uk_n358, 
        u0_uk_n361, u0_uk_n370, u0_uk_n371, u0_uk_n383, u0_uk_n384, u0_uk_n39, u0_uk_n392, u0_uk_n393, u0_uk_n396, 
        u0_uk_n4, u0_uk_n40, u0_uk_n400, u0_uk_n401, u0_uk_n405, u0_uk_n41, u0_uk_n410, u0_uk_n411, u0_uk_n412, 
        u0_uk_n413, u0_uk_n414, u0_uk_n418, u0_uk_n419, u0_uk_n420, u0_uk_n423, u0_uk_n424, u0_uk_n425, u0_uk_n426, 
        u0_uk_n428, u0_uk_n429, u0_uk_n430, u0_uk_n432, u0_uk_n433, u0_uk_n434, u0_uk_n436, u0_uk_n438, u0_uk_n439, 
        u0_uk_n440, u0_uk_n442, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n448, u0_uk_n45, u0_uk_n450, u0_uk_n457, 
        u0_uk_n471, u0_uk_n497, u0_uk_n499, u0_uk_n5, u0_uk_n502, u0_uk_n505, u0_uk_n508, u0_uk_n510, u0_uk_n511, 
        u0_uk_n513, u0_uk_n517, u0_uk_n519, u0_uk_n522, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, 
        u0_uk_n532, u0_uk_n534, u0_uk_n535, u0_uk_n536, u0_uk_n539, u0_uk_n542, u0_uk_n544, u0_uk_n545, u0_uk_n546, 
        u0_uk_n547, u0_uk_n549, u0_uk_n55, u0_uk_n550, u0_uk_n552, u0_uk_n553, u0_uk_n554, u0_uk_n555, u0_uk_n557, 
        u0_uk_n558, u0_uk_n560, u0_uk_n561, u0_uk_n562, u0_uk_n565, u0_uk_n566, u0_uk_n567, u0_uk_n568, u0_uk_n570, 
        u0_uk_n573, u0_uk_n574, u0_uk_n575, u0_uk_n577, u0_uk_n578, u0_uk_n579, u0_uk_n58, u0_uk_n580, u0_uk_n581, 
        u0_uk_n583, u0_uk_n598, u0_uk_n604, u0_uk_n61, u0_uk_n615, u0_uk_n627, u0_uk_n629, u0_uk_n632, u0_uk_n635, 
        u0_uk_n636, u0_uk_n637, u0_uk_n639, u0_uk_n640, u0_uk_n642, u0_uk_n643, u0_uk_n644, u0_uk_n645, u0_uk_n649, 
        u0_uk_n650, u0_uk_n651, u0_uk_n652, u0_uk_n653, u0_uk_n654, u0_uk_n657, u0_uk_n658, u0_uk_n659, u0_uk_n660, 
        u0_uk_n661, u0_uk_n663, u0_uk_n666, u0_uk_n668, u0_uk_n669, u0_uk_n67, u0_uk_n670, u0_uk_n674, u0_uk_n675, 
        u0_uk_n684, u0_uk_n687, u0_uk_n690, u0_uk_n696, u0_uk_n697, u0_uk_n699, u0_uk_n711, u0_uk_n719, u0_uk_n722, 
        u0_uk_n723, u0_uk_n725, u0_uk_n726, u0_uk_n727, u0_uk_n729, u0_uk_n73, u0_uk_n731, u0_uk_n734, u0_uk_n735, 
        u0_uk_n741, u0_uk_n746, u0_uk_n748, u0_uk_n751, u0_uk_n759, u0_uk_n761, u0_uk_n763, u0_uk_n768, u0_uk_n780, 
        u0_uk_n783, u0_uk_n786, u0_uk_n793, u0_uk_n799, u0_uk_n8, u0_uk_n800, u0_uk_n809, u0_uk_n810, u0_uk_n813, 
        u0_uk_n815, u0_uk_n816, u0_uk_n832, u0_uk_n839, u0_uk_n855, u0_uk_n866, u0_uk_n868, u0_uk_n869, u0_uk_n875, 
        u0_uk_n883, u0_uk_n892, u0_uk_n898, u0_uk_n9, u0_uk_n904, u0_uk_n91, u0_uk_n915, u0_uk_n916, u0_uk_n917, 
        u0_uk_n918, u0_uk_n933, u0_uk_n934, u0_uk_n949, u0_uk_n950, u0_uk_n956, u0_uk_n96, u0_uk_n963, u0_uk_n976, 
        u0_uk_n98, u0_uk_n982, u0_uk_n985, u0_uk_n990, u0_uk_n999, u1_FP_33, u1_FP_37, u1_FP_40, u1_FP_41, 
        u1_FP_44, u1_FP_45, u1_FP_52, u1_FP_53, u1_FP_55, u1_FP_56, u1_FP_60, u1_FP_61, u1_K10_1, 
        u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_18, u1_K10_2, u1_K10_20, u1_K10_23, u1_K10_24, u1_K10_25, 
        u1_K10_26, u1_K10_29, u1_K10_30, u1_K10_31, u1_K10_32, u1_K10_36, u1_K10_41, u1_K10_42, u1_K10_43, 
        u1_K10_44, u1_K10_47, u1_K10_48, u1_K10_5, u1_K10_6, u1_K10_7, u1_K10_8, u1_K11_11, u1_K11_13, 
        u1_K11_2, u1_K11_23, u1_K11_25, u1_K11_29, u1_K11_32, u1_K11_35, u1_K11_37, u1_K11_38, u1_K11_48, 
        u1_K11_7, u1_K12_18, u1_K12_19, u1_K12_2, u1_K12_20, u1_K12_24, u1_K12_25, u1_K12_26, u1_K12_35, 
        u1_K12_36, u1_K12_37, u1_K12_38, u1_K12_41, u1_K12_43, u1_K12_47, u1_K12_48, u1_K12_6, u1_K12_8, 
        u1_K13_14, u1_K13_17, u1_K13_18, u1_K13_20, u1_K13_29, u1_K13_30, u1_K13_31, u1_K13_32, u1_K13_35, 
        u1_K13_37, u1_K13_48, u1_K13_8, u1_K14_1, u1_K14_2, u1_K14_29, u1_K14_30, u1_K14_31, u1_K14_32, 
        u1_K14_42, u1_K14_44, u1_K14_47, u1_K14_48, u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_18, 
        u1_K15_2, u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_29, u1_K15_31, u1_K15_32, u1_K15_35, 
        u1_K15_36, u1_K15_37, u1_K15_41, u1_K15_42, u1_K15_44, u1_K15_48, u1_K15_5, u1_K15_6, u1_K15_7, 
        u1_K16_11, u1_K16_12, u1_K16_13, u1_K16_14, u1_K16_17, u1_K16_18, u1_K16_19, u1_K16_2, u1_K16_20, 
        u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_35, u1_K16_41, u1_K16_42, u1_K16_44, u1_K16_48, u1_K16_6, 
        u1_K16_8, u1_K1_1, u1_K1_17, u1_K1_19, u1_K1_43, u1_K1_47, u1_K1_6, u1_K1_8, u1_K2_1, 
        u1_K2_11, u1_K2_12, u1_K2_13, u1_K2_17, u1_K2_18, u1_K2_2, u1_K2_20, u1_K2_23, u1_K2_24, 
        u1_K2_25, u1_K2_26, u1_K2_29, u1_K2_30, u1_K2_31, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_47, 
        u1_K2_48, u1_K2_5, u1_K2_6, u1_K2_8, u1_K3_1, u1_K3_12, u1_K3_14, u1_K3_17, u1_K3_18, 
        u1_K3_19, u1_K3_2, u1_K3_20, u1_K3_23, u1_K3_25, u1_K3_26, u1_K3_29, u1_K3_31, u1_K3_35, 
        u1_K3_36, u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_47, u1_K3_48, 
        u1_K3_5, u1_K3_6, u1_K3_7, u1_K3_8, u1_K4_1, u1_K4_11, u1_K4_12, u1_K4_13, u1_K4_14, 
        u1_K4_17, u1_K4_18, u1_K4_19, u1_K4_24, u1_K4_30, u1_K4_32, u1_K4_35, u1_K4_36, u1_K4_37, 
        u1_K4_38, u1_K4_41, u1_K4_42, u1_K4_43, u1_K4_44, u1_K4_47, u1_K4_48, u1_K4_6, u1_K5_1, 
        u1_K5_11, u1_K5_12, u1_K5_13, u1_K5_14, u1_K5_17, u1_K5_18, u1_K5_19, u1_K5_2, u1_K5_23, 
        u1_K5_24, u1_K5_25, u1_K5_26, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, u1_K5_37, u1_K5_38, 
        u1_K5_41, u1_K5_42, u1_K5_44, u1_K5_47, u1_K5_48, u1_K5_5, u1_K5_6, u1_K5_7, u1_K5_8, 
        u1_K6_1, u1_K6_11, u1_K6_12, u1_K6_13, u1_K6_14, u1_K6_20, u1_K6_23, u1_K6_24, u1_K6_25, 
        u1_K6_26, u1_K6_29, u1_K6_30, u1_K6_31, u1_K6_32, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, 
        u1_K6_41, u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_47, u1_K6_48, u1_K6_5, u1_K6_6, u1_K6_7, 
        u1_K6_8, u1_K7_1, u1_K7_11, u1_K7_14, u1_K7_17, u1_K7_18, u1_K7_19, u1_K7_2, u1_K7_23, 
        u1_K7_26, u1_K7_29, u1_K7_30, u1_K7_31, u1_K7_35, u1_K7_37, u1_K7_38, u1_K7_41, u1_K7_43, 
        u1_K7_44, u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_7, u1_K8_1, u1_K8_11, u1_K8_13, u1_K8_14, 
        u1_K8_18, u1_K8_2, u1_K8_20, u1_K8_23, u1_K8_24, u1_K8_25, u1_K8_26, u1_K8_30, u1_K8_31, 
        u1_K8_32, u1_K8_35, u1_K8_36, u1_K8_38, u1_K8_41, u1_K8_42, u1_K8_44, u1_K8_47, u1_K8_48, 
        u1_K8_5, u1_K8_7, u1_K9_12, u1_K9_13, u1_K9_14, u1_K9_17, u1_K9_23, u1_K9_24, u1_K9_25, 
        u1_K9_29, u1_K9_31, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_43, u1_K9_44, u1_K9_47, u1_K9_5, 
        u1_K9_6, u1_K9_7, u1_K9_8, u1_R0_1, u1_R0_12, u1_R0_13, u1_R0_16, u1_R0_17, u1_R0_20, 
        u1_R0_21, u1_R0_28, u1_R0_29, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_7, u1_R0_8, u1_R0_9, 
        u1_R10_1, u1_R10_10, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_16, u1_R10_17, u1_R10_24, u1_R10_25, 
        u1_R10_28, u1_R10_29, u1_R10_32, u1_R10_5, u1_R11_1, u1_R11_10, u1_R11_12, u1_R11_13, u1_R11_20, 
        u1_R11_21, u1_R11_24, u1_R11_4, u1_R11_5, u1_R11_8, u1_R11_9, u1_R12_1, u1_R12_20, u1_R12_21, 
        u1_R12_23, u1_R12_29, u1_R12_32, u1_R13_1, u1_R13_13, u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, 
        u1_R13_24, u1_R13_25, u1_R13_28, u1_R13_29, u1_R13_4, u1_R13_5, u1_R13_8, u1_R13_9, u1_R1_1, 
        u1_R1_12, u1_R1_13, u1_R1_16, u1_R1_17, u1_R1_20, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, 
        u1_R1_32, u1_R1_4, u1_R1_5, u1_R1_9, u1_R2_1, u1_R2_12, u1_R2_13, u1_R2_16, u1_R2_17, 
        u1_R2_2, u1_R2_20, u1_R2_21, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_32, u1_R2_5, 
        u1_R2_7, u1_R2_8, u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_15, u1_R3_16, u1_R3_17, 
        u1_R3_18, u1_R3_20, u1_R3_21, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_32, u1_R3_4, 
        u1_R3_5, u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_13, u1_R4_14, u1_R4_16, u1_R4_17, u1_R4_20, 
        u1_R4_21, u1_R4_24, u1_R4_25, u1_R4_28, u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, 
        u1_R4_6, u1_R4_7, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_12, u1_R5_13, u1_R5_16, u1_R5_17, 
        u1_R5_18, u1_R5_20, u1_R5_21, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_31, 
        u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_8, u1_R5_9, u1_R6_1, u1_R6_10, u1_R6_13, u1_R6_16, 
        u1_R6_17, u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_28, u1_R6_29, u1_R6_32, 
        u1_R6_4, u1_R6_8, u1_R6_9, u1_R7_1, u1_R7_12, u1_R7_13, u1_R7_15, u1_R7_16, u1_R7_17, 
        u1_R7_18, u1_R7_20, u1_R7_24, u1_R7_25, u1_R7_28, u1_R7_29, u1_R7_32, u1_R7_4, u1_R7_5, 
        u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_13, u1_R8_15, u1_R8_16, u1_R8_17, 
        u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_24, u1_R8_25, u1_R8_28, u1_R8_29, u1_R8_32, u1_R8_4, 
        u1_R8_5, u1_R8_6, u1_R8_8, u1_R8_9, u1_R9_1, u1_R9_12, u1_R9_15, u1_R9_16, u1_R9_20, 
        u1_R9_21, u1_R9_23, u1_R9_24, u1_R9_25, u1_R9_4, u1_R9_8, u1_R9_9, u1_desIn_r_25, u1_desIn_r_29, 
        u1_desIn_r_37, u1_desIn_r_39, u1_desIn_r_57, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_13, u1_u0_X_14, u1_u0_X_15, 
        u1_u0_X_16, u1_u0_X_2, u1_u0_X_21, u1_u0_X_22, u1_u0_X_23, u1_u0_X_24, u1_u0_X_25, u1_u0_X_26, u1_u0_X_27, 
        u1_u0_X_28, u1_u0_X_29, u1_u0_X_3, u1_u0_X_30, u1_u0_X_31, u1_u0_X_32, u1_u0_X_33, u1_u0_X_34, u1_u0_X_35, 
        u1_u0_X_36, u1_u0_X_37, u1_u0_X_38, u1_u0_X_39, u1_u0_X_4, u1_u0_X_40, u1_u0_X_42, u1_u0_X_44, u1_u0_X_45, 
        u1_u0_X_46, u1_u0_X_48, u1_u0_X_5, u1_u0_X_7, u1_u0_X_9, u1_u10_X_1, u1_u10_X_10, u1_u10_X_15, u1_u10_X_16, 
        u1_u10_X_18, u1_u10_X_20, u1_u10_X_21, u1_u10_X_24, u1_u10_X_26, u1_u10_X_27, u1_u10_X_28, u1_u10_X_3, u1_u10_X_33, 
        u1_u10_X_39, u1_u10_X_4, u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_X_43, u1_u10_X_44, u1_u10_X_45, u1_u10_X_46, 
        u1_u10_X_47, u1_u10_X_6, u1_u10_X_8, u1_u10_X_9, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, u1_u11_X_14, 
        u1_u11_X_16, u1_u11_X_22, u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_3, u1_u11_X_30, u1_u11_X_31, u1_u11_X_32, 
        u1_u11_X_33, u1_u11_X_34, u1_u11_X_39, u1_u11_X_4, u1_u11_X_40, u1_u11_X_45, u1_u11_X_46, u1_u11_X_5, u1_u11_X_7, 
        u1_u11_X_9, u1_u12_X_1, u1_u12_X_10, u1_u12_X_16, u1_u12_X_21, u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, u1_u12_X_25, 
        u1_u12_X_26, u1_u12_X_27, u1_u12_X_28, u1_u12_X_3, u1_u12_X_33, u1_u12_X_34, u1_u12_X_36, u1_u12_X_38, u1_u12_X_39, 
        u1_u12_X_4, u1_u12_X_40, u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, 
        u1_u12_X_9, u1_u13_X_10, u1_u13_X_11, u1_u13_X_12, u1_u13_X_13, u1_u13_X_14, u1_u13_X_15, u1_u13_X_16, u1_u13_X_17, 
        u1_u13_X_18, u1_u13_X_19, u1_u13_X_20, u1_u13_X_21, u1_u13_X_22, u1_u13_X_23, u1_u13_X_24, u1_u13_X_25, u1_u13_X_26, 
        u1_u13_X_27, u1_u13_X_28, u1_u13_X_3, u1_u13_X_33, u1_u13_X_35, u1_u13_X_36, u1_u13_X_37, u1_u13_X_38, u1_u13_X_39, 
        u1_u13_X_4, u1_u13_X_40, u1_u13_X_41, u1_u13_X_43, u1_u13_X_45, u1_u13_X_46, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, 
        u1_u13_X_8, u1_u13_X_9, u1_u14_X_1, u1_u14_X_10, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_19, u1_u14_X_21, 
        u1_u14_X_22, u1_u14_X_27, u1_u14_X_28, u1_u14_X_3, u1_u14_X_33, u1_u14_X_34, u1_u14_X_39, u1_u14_X_4, u1_u14_X_40, 
        u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, u1_u14_X_9, u1_u15_X_1, u1_u15_X_10, u1_u15_X_15, u1_u15_X_16, u1_u15_X_21, 
        u1_u15_X_22, u1_u15_X_23, u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, u1_u15_X_27, u1_u15_X_28, u1_u15_X_3, u1_u15_X_33, 
        u1_u15_X_36, u1_u15_X_38, u1_u15_X_39, u1_u15_X_4, u1_u15_X_40, u1_u15_X_45, u1_u15_X_46, u1_u15_X_47, u1_u15_X_5, 
        u1_u15_X_7, u1_u15_X_9, u1_u1_X_15, u1_u1_X_16, u1_u1_X_21, u1_u1_X_22, u1_u1_X_27, u1_u1_X_28, u1_u1_X_3, 
        u1_u1_X_33, u1_u1_X_34, u1_u1_X_35, u1_u1_X_36, u1_u1_X_37, u1_u1_X_38, u1_u1_X_39, u1_u1_X_4, u1_u1_X_40, 
        u1_u1_X_45, u1_u1_X_46, u1_u1_X_9, u1_u2_X_10, u1_u2_X_11, u1_u2_X_13, u1_u2_X_15, u1_u2_X_16, u1_u2_X_21, 
        u1_u2_X_22, u1_u2_X_27, u1_u2_X_28, u1_u2_X_3, u1_u2_X_30, u1_u2_X_32, u1_u2_X_33, u1_u2_X_34, u1_u2_X_39, 
        u1_u2_X_4, u1_u2_X_40, u1_u2_X_45, u1_u2_X_46, u1_u2_X_9, u1_u3_X_15, u1_u3_X_16, u1_u3_X_21, u1_u3_X_22, 
        u1_u3_X_27, u1_u3_X_28, u1_u3_X_33, u1_u3_X_34, u1_u3_X_39, u1_u3_X_4, u1_u3_X_40, u1_u3_X_45, u1_u3_X_46, 
        u1_u3_X_5, u1_u3_X_7, u1_u3_X_9, u1_u4_X_10, u1_u4_X_15, u1_u4_X_16, u1_u4_X_21, u1_u4_X_28, u1_u4_X_3, 
        u1_u4_X_33, u1_u4_X_34, u1_u4_X_39, u1_u4_X_4, u1_u4_X_40, u1_u4_X_45, u1_u4_X_46, u1_u4_X_9, u1_u5_X_15, 
        u1_u5_X_16, u1_u5_X_17, u1_u5_X_19, u1_u5_X_22, u1_u5_X_27, u1_u5_X_28, u1_u5_X_3, u1_u5_X_33, u1_u5_X_34, 
        u1_u5_X_39, u1_u5_X_40, u1_u5_X_45, u1_u5_X_46, u1_u6_X_10, u1_u6_X_15, u1_u6_X_16, u1_u6_X_21, u1_u6_X_22, 
        u1_u6_X_28, u1_u6_X_3, u1_u6_X_33, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, u1_u6_X_45, u1_u6_X_9, u1_u7_X_10, 
        u1_u7_X_16, u1_u7_X_17, u1_u7_X_19, u1_u7_X_21, u1_u7_X_22, u1_u7_X_27, u1_u7_X_28, u1_u7_X_33, u1_u7_X_34, 
        u1_u7_X_39, u1_u7_X_4, u1_u7_X_40, u1_u7_X_45, u1_u7_X_46, u1_u7_X_6, u1_u7_X_8, u1_u7_X_9, u1_u8_X_15, 
        u1_u8_X_16, u1_u8_X_21, u1_u8_X_28, u1_u8_X_3, u1_u8_X_30, u1_u8_X_32, u1_u8_X_33, u1_u8_X_34, u1_u8_X_39, 
        u1_u8_X_4, u1_u8_X_40, u1_u8_X_45, u1_u8_X_46, u1_u9_X_10, u1_u9_X_15, u1_u9_X_16, u1_u9_X_17, u1_u9_X_19, 
        u1_u9_X_21, u1_u9_X_27, u1_u9_X_28, u1_u9_X_3, u1_u9_X_34, u1_u9_X_39, u1_u9_X_4, u1_u9_X_40, u1_u9_X_45, 
        u1_u9_X_46, u1_uk_n1002, u1_uk_n1003, u1_uk_n1015, u1_uk_n1021, u1_uk_n1023, u1_uk_n1025, u1_uk_n1029, u1_uk_n1031, 
        u1_uk_n1034, u1_uk_n1038, u1_uk_n1050, u1_uk_n1054, u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1060, u1_uk_n1061, 
        u1_uk_n1063, u1_uk_n1065, u1_uk_n1070, u1_uk_n1073, u1_uk_n1074, u1_uk_n1076, u1_uk_n1079, u1_uk_n1080, u1_uk_n1083, 
        u1_uk_n1088, u1_uk_n1090, u1_uk_n1092, u1_uk_n1096, u1_uk_n1101, u1_uk_n1104, u1_uk_n1105, u1_uk_n1106, u1_uk_n1109, 
        u1_uk_n1113, u1_uk_n1114, u1_uk_n1115, u1_uk_n1118, u1_uk_n1119, u1_uk_n1121, u1_uk_n1123, u1_uk_n1124, u1_uk_n1125, 
        u1_uk_n1126, u1_uk_n1128, u1_uk_n1130, u1_uk_n1134, u1_uk_n1138, u1_uk_n1140, u1_uk_n1143, u1_uk_n1147, u1_uk_n1148, 
        u1_uk_n1153, u1_uk_n1154, u1_uk_n1155, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1159, u1_uk_n1160, u1_uk_n1163, 
        u1_uk_n1166, u1_uk_n1167, u1_uk_n1170, u1_uk_n1171, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, u1_uk_n366, 
        u1_uk_n369, u1_uk_n376, u1_uk_n379, u1_uk_n382, u1_uk_n385, u1_uk_n386, u1_uk_n407, u1_uk_n421, u1_uk_n437, 
        u1_uk_n443, u1_uk_n454, u1_uk_n496, u1_uk_n504, u1_uk_n509, u1_uk_n515, u1_uk_n520, u1_uk_n524, u1_uk_n605, 
        u1_uk_n608, u1_uk_n672, u1_uk_n676, u1_uk_n677, u1_uk_n678, u1_uk_n685, u1_uk_n702, u1_uk_n948, u1_uk_n949, 
        u1_uk_n950, u1_uk_n955, u1_uk_n969, u1_uk_n970, u1_uk_n973, u1_uk_n974, u1_uk_n976, u1_uk_n985, u1_uk_n988, 
        u1_uk_n989, u1_uk_n993, u2_FP_33, u2_FP_36, u2_FP_37, u2_FP_40, u2_FP_41, u2_FP_44, u2_FP_45, 
        u2_FP_48, u2_FP_49, u2_FP_52, u2_FP_53, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_60, u2_FP_61, 
        u2_FP_64, u2_K10_1, u2_K10_11, u2_K10_13, u2_K10_14, u2_K10_17, u2_K10_18, u2_K10_19, u2_K10_20, 
        u2_K10_23, u2_K10_24, u2_K10_25, u2_K10_26, u2_K10_36, u2_K10_42, u2_K10_43, u2_K10_44, u2_K10_48, 
        u2_K10_5, u2_K10_7, u2_K10_8, u2_K11_11, u2_K11_13, u2_K11_24, u2_K11_26, u2_K11_29, u2_K12_2, 
        u2_K12_20, u2_K12_25, u2_K12_36, u2_K12_38, u2_K12_47, u2_K12_48, u2_K13_32, u2_K13_35, u2_K13_37, 
        u2_K13_48, u2_K14_38, u2_K15_1, u2_K15_12, u2_K15_17, u2_K15_2, u2_K15_23, u2_K15_29, u2_K15_31, 
        u2_K15_35, u2_K15_44, u2_K16_1, u2_K16_11, u2_K16_12, u2_K16_13, u2_K16_14, u2_K16_17, u2_K16_18, 
        u2_K16_19, u2_K16_2, u2_K16_20, u2_K16_23, u2_K16_24, u2_K16_25, u2_K16_26, u2_K16_30, u2_K16_31, 
        u2_K16_32, u2_K16_35, u2_K16_36, u2_K16_38, u2_K16_41, u2_K16_42, u2_K16_44, u2_K16_47, u2_K16_48, 
        u2_K16_5, u2_K16_6, u2_K16_7, u2_K16_8, u2_K1_43, u2_K2_1, u2_K2_11, u2_K2_12, u2_K2_13, 
        u2_K2_17, u2_K2_18, u2_K2_2, u2_K2_20, u2_K2_23, u2_K2_24, u2_K2_25, u2_K2_26, u2_K2_29, 
        u2_K2_30, u2_K2_31, u2_K2_35, u2_K2_36, u2_K2_37, u2_K2_38, u2_K2_42, u2_K2_44, u2_K2_47, 
        u2_K2_48, u2_K2_5, u2_K2_6, u2_K2_8, u2_K3_13, u2_K3_19, u2_K3_20, u2_K3_23, u2_K3_26, 
        u2_K3_42, u2_K3_43, u2_K3_47, u2_K3_48, u2_K4_14, u2_K4_18, u2_K4_19, u2_K4_24, u2_K4_48, 
        u2_K4_6, u2_K4_7, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_17, u2_K5_18, u2_K5_19, u2_K5_2, 
        u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_29, u2_K5_30, u2_K5_31, u2_K5_32, u2_K5_37, 
        u2_K5_38, u2_K5_41, u2_K5_44, u2_K5_48, u2_K5_5, u2_K5_6, u2_K5_8, u2_K6_1, u2_K6_11, 
        u2_K6_13, u2_K6_14, u2_K6_19, u2_K6_20, u2_K6_24, u2_K6_32, u2_K6_47, u2_K6_6, u2_K6_8, 
        u2_K7_26, u2_K7_30, u2_K7_31, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_48, u2_K7_5, 
        u2_K7_7, u2_K8_1, u2_K8_11, u2_K8_13, u2_K8_14, u2_K8_17, u2_K8_18, u2_K8_19, u2_K8_2, 
        u2_K8_20, u2_K8_47, u2_K8_48, u2_K8_5, u2_K8_6, u2_K8_7, u2_K8_8, u2_K9_12, u2_K9_14, 
        u2_K9_23, u2_K9_25, u2_K9_36, u2_K9_37, u2_K9_38, u2_K9_43, u2_K9_5, u2_R0_1, u2_R0_12, 
        u2_R0_13, u2_R0_16, u2_R0_17, u2_R0_19, u2_R0_20, u2_R0_21, u2_R0_24, u2_R0_25, u2_R0_29, 
        u2_R0_32, u2_R0_4, u2_R0_5, u2_R0_7, u2_R0_8, u2_R0_9, u2_R10_1, u2_R10_12, u2_R10_13, 
        u2_R10_16, u2_R10_21, u2_R10_25, u2_R10_29, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_7, u2_R10_8, 
        u2_R10_9, u2_R11_1, u2_R11_21, u2_R11_24, u2_R11_4, u2_R12_20, u2_R12_21, u2_R12_22, u2_R12_25, 
        u2_R13_1, u2_R13_12, u2_R13_16, u2_R13_17, u2_R13_20, u2_R13_22, u2_R13_24, u2_R13_25, u2_R13_27, 
        u2_R13_29, u2_R13_32, u2_R13_5, u2_R13_9, u2_R1_1, u2_R1_12, u2_R1_13, u2_R1_14, u2_R1_15, 
        u2_R1_16, u2_R1_17, u2_R1_2, u2_R1_25, u2_R1_27, u2_R1_28, u2_R1_29, u2_R1_3, u2_R1_30, 
        u2_R1_31, u2_R1_32, u2_R1_5, u2_R1_6, u2_R1_7, u2_R1_8, u2_R1_9, u2_R2_1, u2_R2_10, 
        u2_R2_11, u2_R2_12, u2_R2_13, u2_R2_16, u2_R2_17, u2_R2_19, u2_R2_2, u2_R2_20, u2_R2_21, 
        u2_R2_25, u2_R2_3, u2_R2_32, u2_R2_4, u2_R2_5, u2_R2_6, u2_R2_7, u2_R2_8, u2_R2_9, 
        u2_R3_1, u2_R3_12, u2_R3_13, u2_R3_16, u2_R3_17, u2_R3_18, u2_R3_20, u2_R3_21, u2_R3_22, 
        u2_R3_24, u2_R3_25, u2_R3_28, u2_R3_29, u2_R3_30, u2_R3_4, u2_R3_5, u2_R3_8, u2_R3_9, 
        u2_R4_1, u2_R4_12, u2_R4_13, u2_R4_14, u2_R4_17, u2_R4_21, u2_R4_22, u2_R4_24, u2_R4_28, 
        u2_R4_29, u2_R4_31, u2_R4_32, u2_R4_4, u2_R4_5, u2_R4_6, u2_R4_8, u2_R4_9, u2_R5_1, 
        u2_R5_10, u2_R5_11, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_16, u2_R5_17, u2_R5_20, u2_R5_21, 
        u2_R5_23, u2_R5_24, u2_R5_25, u2_R5_26, u2_R5_28, u2_R5_29, u2_R5_32, u2_R5_4, u2_R5_5, 
        u2_R5_8, u2_R5_9, u2_R6_1, u2_R6_12, u2_R6_13, u2_R6_2, u2_R6_28, u2_R6_32, u2_R6_4, 
        u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_1, u2_R7_11, u2_R7_12, u2_R7_13, u2_R7_14, u2_R7_15, 
        u2_R7_16, u2_R7_17, u2_R7_22, u2_R7_24, u2_R7_25, u2_R7_28, u2_R7_29, u2_R7_3, u2_R7_4, 
        u2_R7_5, u2_R7_6, u2_R7_7, u2_R7_8, u2_R7_9, u2_R8_1, u2_R8_12, u2_R8_13, u2_R8_15, 
        u2_R8_16, u2_R8_17, u2_R8_20, u2_R8_22, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, 
        u2_R8_29, u2_R8_32, u2_R8_4, u2_R8_5, u2_R8_6, u2_R8_8, u2_R8_9, u2_R9_12, u2_R9_13, 
        u2_R9_17, u2_R9_20, u2_R9_32, u2_R9_8, u2_R9_9, u2_desIn_r_1, u2_desIn_r_25, u2_desIn_r_27, u2_desIn_r_33, 
        u2_desIn_r_57, u2_key_r_14, u2_key_r_23, u2_key_r_30, u2_key_r_7, u2_u0_X_10, u2_u0_X_11, u2_u0_X_12, u2_u0_X_25, 
        u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_30, u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, u2_u0_X_37, 
        u2_u0_X_39, u2_u0_X_40, u2_u0_X_45, u2_u0_X_46, u2_u0_X_48, u2_u0_X_7, u2_u0_X_8, u2_u0_X_9, u2_u10_X_10, 
        u2_u10_X_15, u2_u10_X_16, u2_u10_X_18, u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_25, u2_u10_X_27, u2_u10_X_28, 
        u2_u10_X_30, u2_u10_X_32, u2_u10_X_33, u2_u10_X_34, u2_u10_X_35, u2_u10_X_36, u2_u10_X_37, u2_u10_X_38, u2_u10_X_39, 
        u2_u10_X_40, u2_u10_X_41, u2_u10_X_42, u2_u10_X_43, u2_u10_X_44, u2_u10_X_45, u2_u10_X_46, u2_u10_X_48, u2_u10_X_7, 
        u2_u10_X_8, u2_u10_X_9, u2_u11_X_15, u2_u11_X_16, u2_u11_X_21, u2_u11_X_22, u2_u11_X_24, u2_u11_X_26, u2_u11_X_27, 
        u2_u11_X_28, u2_u11_X_29, u2_u11_X_3, u2_u11_X_31, u2_u11_X_33, u2_u11_X_34, u2_u11_X_35, u2_u11_X_37, u2_u11_X_39, 
        u2_u11_X_40, u2_u11_X_41, u2_u11_X_43, u2_u11_X_45, u2_u11_X_46, u2_u11_X_6, u2_u11_X_8, u2_u11_X_9, u2_u12_X_1, 
        u2_u12_X_10, u2_u12_X_11, u2_u12_X_12, u2_u12_X_25, u2_u12_X_26, u2_u12_X_27, u2_u12_X_28, u2_u12_X_29, u2_u12_X_3, 
        u2_u12_X_31, u2_u12_X_33, u2_u12_X_34, u2_u12_X_36, u2_u12_X_38, u2_u12_X_39, u2_u12_X_4, u2_u12_X_40, u2_u12_X_41, 
        u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, u2_u12_X_46, u2_u12_X_47, u2_u12_X_6, u2_u12_X_8, u2_u12_X_9, 
        u2_u13_X_25, u2_u13_X_26, u2_u13_X_27, u2_u13_X_28, u2_u13_X_34, u2_u13_X_35, u2_u13_X_37, u2_u13_X_39, u2_u13_X_40, 
        u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, u2_u13_X_47, u2_u13_X_48, u2_u14_X_10, 
        u2_u14_X_11, u2_u14_X_13, u2_u14_X_15, u2_u14_X_16, u2_u14_X_18, u2_u14_X_20, u2_u14_X_21, u2_u14_X_22, u2_u14_X_27, 
        u2_u14_X_28, u2_u14_X_3, u2_u14_X_30, u2_u14_X_32, u2_u14_X_34, u2_u14_X_39, u2_u14_X_4, u2_u14_X_41, u2_u14_X_43, 
        u2_u14_X_45, u2_u14_X_46, u2_u14_X_5, u2_u14_X_7, u2_u14_X_9, u2_u15_X_10, u2_u15_X_15, u2_u15_X_16, u2_u15_X_21, 
        u2_u15_X_22, u2_u15_X_27, u2_u15_X_28, u2_u15_X_3, u2_u15_X_33, u2_u15_X_39, u2_u15_X_4, u2_u15_X_40, u2_u15_X_45, 
        u2_u15_X_46, u2_u15_X_9, u2_u1_X_15, u2_u1_X_16, u2_u1_X_21, u2_u1_X_22, u2_u1_X_27, u2_u1_X_3, u2_u1_X_33, 
        u2_u1_X_34, u2_u1_X_39, u2_u1_X_4, u2_u1_X_40, u2_u1_X_41, u2_u1_X_43, u2_u1_X_45, u2_u1_X_46, u2_u1_X_9, 
        u2_u2_X_15, u2_u2_X_16, u2_u2_X_27, u2_u2_X_28, u2_u2_X_29, u2_u2_X_30, u2_u2_X_31, u2_u2_X_32, u2_u2_X_33, 
        u2_u2_X_34, u2_u2_X_35, u2_u2_X_37, u2_u2_X_39, u2_u2_X_5, u2_u2_X_7, u2_u3_X_21, u2_u3_X_22, u2_u3_X_27, 
        u2_u3_X_33, u2_u3_X_34, u2_u3_X_35, u2_u3_X_43, u2_u3_X_44, u2_u3_X_45, u2_u3_X_46, u2_u4_X_1, u2_u4_X_10, 
        u2_u4_X_15, u2_u4_X_16, u2_u4_X_21, u2_u4_X_22, u2_u4_X_28, u2_u4_X_3, u2_u4_X_34, u2_u4_X_39, u2_u4_X_4, 
        u2_u4_X_40, u2_u4_X_46, u2_u4_X_47, u2_u4_X_9, u2_u5_X_10, u2_u5_X_15, u2_u5_X_16, u2_u5_X_22, u2_u5_X_23, 
        u2_u5_X_25, u2_u5_X_27, u2_u5_X_28, u2_u5_X_29, u2_u5_X_3, u2_u5_X_31, u2_u5_X_34, u2_u5_X_36, u2_u5_X_38, 
        u2_u5_X_39, u2_u5_X_4, u2_u5_X_40, u2_u5_X_45, u2_u6_X_10, u2_u6_X_22, u2_u6_X_27, u2_u6_X_28, u2_u6_X_3, 
        u2_u6_X_33, u2_u6_X_4, u2_u6_X_40, u2_u6_X_45, u2_u6_X_46, u2_u6_X_9, u2_u7_X_10, u2_u7_X_15, u2_u7_X_16, 
        u2_u7_X_21, u2_u7_X_22, u2_u7_X_23, u2_u7_X_24, u2_u7_X_4, u2_u7_X_44, u2_u7_X_45, u2_u7_X_46, u2_u7_X_9, 
        u2_u8_X_1, u2_u8_X_15, u2_u8_X_27, u2_u8_X_28, u2_u8_X_29, u2_u8_X_3, u2_u8_X_30, u2_u8_X_31, u2_u8_X_32, 
        u2_u8_X_34, u2_u8_X_39, u2_u8_X_40, u2_u8_X_45, u2_u8_X_46, u2_u8_X_47, u2_u9_X_10, u2_u9_X_15, u2_u9_X_16, 
        u2_u9_X_21, u2_u9_X_27, u2_u9_X_28, u2_u9_X_29, u2_u9_X_3, u2_u9_X_30, u2_u9_X_32, u2_u9_X_34, u2_u9_X_4, 
        u2_u9_X_45, u2_u9_X_46, u2_u9_X_6, u2_uk_K_r11_28, u2_uk_K_r11_48, u2_uk_K_r11_53, u2_uk_K_r13_22, u2_uk_K_r13_32, u2_uk_K_r1_15, 
        u2_uk_K_r1_16, u2_uk_K_r1_18, u2_uk_K_r1_21, u2_uk_K_r1_22, u2_uk_K_r1_47, u2_uk_K_r2_13, u2_uk_K_r2_18, u2_uk_K_r2_21, u2_uk_K_r2_25, 
        u2_uk_K_r2_27, u2_uk_K_r2_28, u2_uk_K_r2_31, u2_uk_K_r2_36, u2_uk_K_r2_49, u2_uk_K_r2_55, u2_uk_K_r3_11, u2_uk_K_r3_14, u2_uk_K_r3_19, 
        u2_uk_K_r3_43, u2_uk_K_r3_9, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_33, u2_uk_K_r4_35, u2_uk_K_r4_38, u2_uk_K_r4_4, u2_uk_K_r4_5, 
        u2_uk_K_r4_55, u2_uk_K_r5_10, u2_uk_K_r5_17, u2_uk_K_r5_19, u2_uk_K_r5_39, u2_uk_K_r5_4, u2_uk_K_r5_41, u2_uk_K_r7_0, u2_uk_K_r7_25, 
        u2_uk_K_r7_26, u2_uk_K_r7_32, u2_uk_K_r7_39, u2_uk_K_r7_41, u2_uk_K_r7_48, u2_uk_K_r7_55, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, 
        u2_uk_K_r8_37, u2_uk_K_r8_41, u2_uk_K_r8_42, u2_uk_K_r9_10, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_n1004, u2_uk_n1008, u2_uk_n1020, 
        u2_uk_n1024, u2_uk_n1027, u2_uk_n1028, u2_uk_n1031, u2_uk_n1035, u2_uk_n1038, u2_uk_n1040, u2_uk_n1043, u2_uk_n1046, 
        u2_uk_n1049, u2_uk_n1050, u2_uk_n1053, u2_uk_n1069, u2_uk_n1074, u2_uk_n1076, u2_uk_n1077, u2_uk_n1079, u2_uk_n1082, 
        u2_uk_n1083, u2_uk_n1084, u2_uk_n1088, u2_uk_n1089, u2_uk_n1091, u2_uk_n1093, u2_uk_n1096, u2_uk_n1098, u2_uk_n1110, 
        u2_uk_n1113, u2_uk_n1120, u2_uk_n1123, u2_uk_n1124, u2_uk_n1128, u2_uk_n1130, u2_uk_n1132, u2_uk_n1133, u2_uk_n1136, 
        u2_uk_n1137, u2_uk_n1140, u2_uk_n1141, u2_uk_n1142, u2_uk_n1152, u2_uk_n1171, u2_uk_n1279, u2_uk_n1280, u2_uk_n1281, 
        u2_uk_n1282, u2_uk_n1283, u2_uk_n1284, u2_uk_n1285, u2_uk_n1286, u2_uk_n1287, u2_uk_n1288, u2_uk_n1290, u2_uk_n1291, 
        u2_uk_n1293, u2_uk_n1295, u2_uk_n1296, u2_uk_n1297, u2_uk_n1300, u2_uk_n1301, u2_uk_n1302, u2_uk_n1305, u2_uk_n1306, 
        u2_uk_n1310, u2_uk_n1311, u2_uk_n1314, u2_uk_n1316, u2_uk_n1317, u2_uk_n1318, u2_uk_n1323, u2_uk_n1324, u2_uk_n1326, 
        u2_uk_n1328, u2_uk_n1329, u2_uk_n1333, u2_uk_n1339, u2_uk_n1341, u2_uk_n1345, u2_uk_n1346, u2_uk_n1350, u2_uk_n1351, 
        u2_uk_n1356, u2_uk_n1359, u2_uk_n1361, u2_uk_n1370, u2_uk_n1375, u2_uk_n1382, u2_uk_n1401, u2_uk_n1405, u2_uk_n1408, 
        u2_uk_n1410, u2_uk_n1413, u2_uk_n1422, u2_uk_n1426, u2_uk_n1428, u2_uk_n1433, u2_uk_n1435, u2_uk_n1438, u2_uk_n1439, 
        u2_uk_n1440, u2_uk_n1441, u2_uk_n1445, u2_uk_n1446, u2_uk_n1447, u2_uk_n1453, u2_uk_n1454, u2_uk_n1456, u2_uk_n1458, 
        u2_uk_n1459, u2_uk_n1462, u2_uk_n1465, u2_uk_n1466, u2_uk_n1470, u2_uk_n1475, u2_uk_n1480, u2_uk_n1486, u2_uk_n1488, 
        u2_uk_n1490, u2_uk_n1493, u2_uk_n1494, u2_uk_n1496, u2_uk_n1497, u2_uk_n1544, u2_uk_n1548, u2_uk_n1549, u2_uk_n1555, 
        u2_uk_n1556, u2_uk_n1563, u2_uk_n1568, u2_uk_n1573, u2_uk_n1580, u2_uk_n1585, u2_uk_n1586, u2_uk_n1592, u2_uk_n1594, 
        u2_uk_n1609, u2_uk_n1615, u2_uk_n1622, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n1693, u2_uk_n1708, 
        u2_uk_n1709, u2_uk_n1720, u2_uk_n1721, u2_uk_n1746, u2_uk_n1769, u2_uk_n1770, u2_uk_n1781, u2_uk_n1785, u2_uk_n1797, 
        u2_uk_n1803, u2_uk_n1807, u2_uk_n1808, u2_uk_n1816, u2_uk_n1817, u2_uk_n1819, u2_uk_n1821, u2_uk_n1824, u2_uk_n1826, 
        u2_uk_n1834, u2_uk_n1840, u2_uk_n1846, u2_uk_n1849, u2_uk_n1851, u2_uk_n1852, u2_uk_n1855, u2_uk_n1856, u2_uk_n238, 
        u2_uk_n240, u2_uk_n257, u2_uk_n299, u2_uk_n301, u2_uk_n305, u2_uk_n308, u2_uk_n313, u2_uk_n319, u2_uk_n335, 
        u2_uk_n373, u2_uk_n386, u2_uk_n408, u2_uk_n415, u2_uk_n421, u2_uk_n454, u2_uk_n456, u2_uk_n467, u2_uk_n503, 
        u2_uk_n504, u2_uk_n515, u2_uk_n520, u2_uk_n665, u2_uk_n682, u2_uk_n689, u2_uk_n939, u2_uk_n942, u2_uk_n943, 
        u2_uk_n945, u2_uk_n946, u2_uk_n955, u2_uk_n958, u2_uk_n959, u2_uk_n963, u2_uk_n985, u2_uk_n986, u2_uk_n987, 
        u2_uk_n991, u2_uk_n993, u2_uk_n995, u2_uk_n998, u2_uk_n999;
  wire key_a_0, key_a_1, key_a_10, key_a_11, key_a_12, key_a_13, key_a_14, key_a_15, key_a_16, 
       key_a_17, key_a_18, key_a_19, key_a_2, key_a_20, key_a_21, key_a_22, key_a_23, key_a_24, 
       key_a_25, key_a_26, key_a_27, key_a_28, key_a_29, key_a_3, key_a_30, key_a_31, key_a_32, 
       key_a_33, key_a_34, key_a_35, key_a_36, key_a_37, key_a_38, key_a_39, key_a_4, key_a_40, 
       key_a_41, key_a_42, key_a_43, key_a_44, key_a_45, key_a_46, key_a_47, key_a_48, key_a_49, 
       key_a_5, key_a_50, key_a_51, key_a_52, key_a_53, key_a_54, key_a_55, key_a_6, key_a_7, 
       key_a_8, key_a_9, key_b_r_0_0, key_b_r_0_1, key_b_r_0_10, key_b_r_0_11, key_b_r_0_12, key_b_r_0_13, key_b_r_0_14, 
       key_b_r_0_15, key_b_r_0_16, key_b_r_0_17, key_b_r_0_18, key_b_r_0_19, key_b_r_0_2, key_b_r_0_20, key_b_r_0_21, key_b_r_0_22, 
       key_b_r_0_23, key_b_r_0_24, key_b_r_0_25, key_b_r_0_26, key_b_r_0_27, key_b_r_0_28, key_b_r_0_29, key_b_r_0_3, key_b_r_0_30, 
       key_b_r_0_31, key_b_r_0_32, key_b_r_0_33, key_b_r_0_34, key_b_r_0_35, key_b_r_0_36, key_b_r_0_37, key_b_r_0_38, key_b_r_0_39, 
       key_b_r_0_4, key_b_r_0_40, key_b_r_0_41, key_b_r_0_42, key_b_r_0_43, key_b_r_0_44, key_b_r_0_45, key_b_r_0_46, key_b_r_0_47, 
       key_b_r_0_48, key_b_r_0_49, key_b_r_0_5, key_b_r_0_50, key_b_r_0_51, key_b_r_0_52, key_b_r_0_53, key_b_r_0_54, key_b_r_0_55, 
       key_b_r_0_6, key_b_r_0_7, key_b_r_0_8, key_b_r_0_9, key_b_r_10_0, key_b_r_10_1, key_b_r_10_10, key_b_r_10_11, key_b_r_10_12, 
       key_b_r_10_13, key_b_r_10_14, key_b_r_10_15, key_b_r_10_16, key_b_r_10_17, key_b_r_10_18, key_b_r_10_19, key_b_r_10_2, key_b_r_10_20, 
       key_b_r_10_21, key_b_r_10_22, key_b_r_10_23, key_b_r_10_24, key_b_r_10_25, key_b_r_10_26, key_b_r_10_27, key_b_r_10_28, key_b_r_10_29, 
       key_b_r_10_3, key_b_r_10_30, key_b_r_10_31, key_b_r_10_32, key_b_r_10_33, key_b_r_10_34, key_b_r_10_35, key_b_r_10_36, key_b_r_10_37, 
       key_b_r_10_38, key_b_r_10_39, key_b_r_10_4, key_b_r_10_40, key_b_r_10_41, key_b_r_10_42, key_b_r_10_43, key_b_r_10_44, key_b_r_10_45, 
       key_b_r_10_46, key_b_r_10_47, key_b_r_10_48, key_b_r_10_49, key_b_r_10_5, key_b_r_10_50, key_b_r_10_51, key_b_r_10_52, key_b_r_10_53, 
       key_b_r_10_54, key_b_r_10_55, key_b_r_10_6, key_b_r_10_7, key_b_r_10_8, key_b_r_10_9, key_b_r_11_0, key_b_r_11_1, key_b_r_11_10, 
       key_b_r_11_11, key_b_r_11_12, key_b_r_11_13, key_b_r_11_14, key_b_r_11_15, key_b_r_11_16, key_b_r_11_17, key_b_r_11_18, key_b_r_11_19, 
       key_b_r_11_2, key_b_r_11_20, key_b_r_11_21, key_b_r_11_22, key_b_r_11_23, key_b_r_11_24, key_b_r_11_25, key_b_r_11_26, key_b_r_11_27, 
       key_b_r_11_28, key_b_r_11_29, key_b_r_11_3, key_b_r_11_30, key_b_r_11_31, key_b_r_11_32, key_b_r_11_33, key_b_r_11_34, key_b_r_11_35, 
       key_b_r_11_36, key_b_r_11_37, key_b_r_11_38, key_b_r_11_39, key_b_r_11_4, key_b_r_11_40, key_b_r_11_41, key_b_r_11_42, key_b_r_11_43, 
       key_b_r_11_44, key_b_r_11_45, key_b_r_11_46, key_b_r_11_47, key_b_r_11_48, key_b_r_11_49, key_b_r_11_5, key_b_r_11_50, key_b_r_11_51, 
       key_b_r_11_52, key_b_r_11_53, key_b_r_11_54, key_b_r_11_55, key_b_r_11_6, key_b_r_11_7, key_b_r_11_8, key_b_r_11_9, key_b_r_12_0, 
       key_b_r_12_1, key_b_r_12_10, key_b_r_12_11, key_b_r_12_12, key_b_r_12_13, key_b_r_12_14, key_b_r_12_15, key_b_r_12_16, key_b_r_12_17, 
       key_b_r_12_18, key_b_r_12_19, key_b_r_12_2, key_b_r_12_20, key_b_r_12_21, key_b_r_12_22, key_b_r_12_23, key_b_r_12_24, key_b_r_12_25, 
       key_b_r_12_26, key_b_r_12_27, key_b_r_12_28, key_b_r_12_29, key_b_r_12_3, key_b_r_12_30, key_b_r_12_31, key_b_r_12_32, key_b_r_12_33, 
       key_b_r_12_34, key_b_r_12_35, key_b_r_12_36, key_b_r_12_37, key_b_r_12_38, key_b_r_12_39, key_b_r_12_4, key_b_r_12_40, key_b_r_12_41, 
       key_b_r_12_42, key_b_r_12_43, key_b_r_12_44, key_b_r_12_45, key_b_r_12_46, key_b_r_12_47, key_b_r_12_48, key_b_r_12_49, key_b_r_12_5, 
       key_b_r_12_50, key_b_r_12_51, key_b_r_12_52, key_b_r_12_53, key_b_r_12_54, key_b_r_12_55, key_b_r_12_6, key_b_r_12_7, key_b_r_12_8, 
       key_b_r_12_9, key_b_r_13_0, key_b_r_13_1, key_b_r_13_10, key_b_r_13_11, key_b_r_13_12, key_b_r_13_13, key_b_r_13_14, key_b_r_13_15, 
       key_b_r_13_16, key_b_r_13_17, key_b_r_13_18, key_b_r_13_19, key_b_r_13_2, key_b_r_13_20, key_b_r_13_21, key_b_r_13_22, key_b_r_13_23, 
       key_b_r_13_24, key_b_r_13_25, key_b_r_13_26, key_b_r_13_27, key_b_r_13_28, key_b_r_13_29, key_b_r_13_3, key_b_r_13_30, key_b_r_13_31, 
       key_b_r_13_32, key_b_r_13_33, key_b_r_13_34, key_b_r_13_35, key_b_r_13_36, key_b_r_13_37, key_b_r_13_38, key_b_r_13_39, key_b_r_13_4, 
       key_b_r_13_40, key_b_r_13_41, key_b_r_13_42, key_b_r_13_43, key_b_r_13_44, key_b_r_13_45, key_b_r_13_46, key_b_r_13_47, key_b_r_13_48, 
       key_b_r_13_49, key_b_r_13_5, key_b_r_13_50, key_b_r_13_51, key_b_r_13_52, key_b_r_13_53, key_b_r_13_54, key_b_r_13_55, key_b_r_13_6, 
       key_b_r_13_7, key_b_r_13_8, key_b_r_13_9, key_b_r_14_0, key_b_r_14_1, key_b_r_14_10, key_b_r_14_11, key_b_r_14_12, key_b_r_14_13, 
       key_b_r_14_14, key_b_r_14_15, key_b_r_14_16, key_b_r_14_17, key_b_r_14_18, key_b_r_14_19, key_b_r_14_2, key_b_r_14_20, key_b_r_14_21, 
       key_b_r_14_22, key_b_r_14_23, key_b_r_14_24, key_b_r_14_25, key_b_r_14_26, key_b_r_14_27, key_b_r_14_28, key_b_r_14_29, key_b_r_14_3, 
       key_b_r_14_30, key_b_r_14_31, key_b_r_14_32, key_b_r_14_33, key_b_r_14_34, key_b_r_14_35, key_b_r_14_36, key_b_r_14_37, key_b_r_14_38, 
       key_b_r_14_39, key_b_r_14_4, key_b_r_14_40, key_b_r_14_41, key_b_r_14_42, key_b_r_14_43, key_b_r_14_44, key_b_r_14_45, key_b_r_14_46, 
       key_b_r_14_47, key_b_r_14_48, key_b_r_14_49, key_b_r_14_5, key_b_r_14_50, key_b_r_14_51, key_b_r_14_52, key_b_r_14_53, key_b_r_14_54, 
       key_b_r_14_55, key_b_r_14_6, key_b_r_14_7, key_b_r_14_8, key_b_r_14_9, key_b_r_15_0, key_b_r_15_1, key_b_r_15_10, key_b_r_15_11, 
       key_b_r_15_12, key_b_r_15_13, key_b_r_15_14, key_b_r_15_15, key_b_r_15_16, key_b_r_15_17, key_b_r_15_18, key_b_r_15_19, key_b_r_15_2, 
       key_b_r_15_20, key_b_r_15_21, key_b_r_15_22, key_b_r_15_23, key_b_r_15_24, key_b_r_15_25, key_b_r_15_26, key_b_r_15_27, key_b_r_15_28, 
       key_b_r_15_29, key_b_r_15_3, key_b_r_15_30, key_b_r_15_31, key_b_r_15_32, key_b_r_15_33, key_b_r_15_34, key_b_r_15_35, key_b_r_15_36, 
       key_b_r_15_37, key_b_r_15_38, key_b_r_15_39, key_b_r_15_4, key_b_r_15_40, key_b_r_15_41, key_b_r_15_42, key_b_r_15_43, key_b_r_15_44, 
       key_b_r_15_45, key_b_r_15_46, key_b_r_15_47, key_b_r_15_48, key_b_r_15_49, key_b_r_15_5, key_b_r_15_50, key_b_r_15_51, key_b_r_15_52, 
       key_b_r_15_53, key_b_r_15_54, key_b_r_15_55, key_b_r_15_6, key_b_r_15_7, key_b_r_15_8, key_b_r_15_9, key_b_r_16_0, key_b_r_16_1, 
       key_b_r_16_10, key_b_r_16_11, key_b_r_16_12, key_b_r_16_13, key_b_r_16_14, key_b_r_16_15, key_b_r_16_16, key_b_r_16_17, key_b_r_16_18, 
       key_b_r_16_19, key_b_r_16_2, key_b_r_16_20, key_b_r_16_21, key_b_r_16_22, key_b_r_16_23, key_b_r_16_24, key_b_r_16_25, key_b_r_16_26, 
       key_b_r_16_27, key_b_r_16_28, key_b_r_16_29, key_b_r_16_3, key_b_r_16_30, key_b_r_16_31, key_b_r_16_32, key_b_r_16_33, key_b_r_16_34, 
       key_b_r_16_35, key_b_r_16_36, key_b_r_16_37, key_b_r_16_38, key_b_r_16_39, key_b_r_16_4, key_b_r_16_40, key_b_r_16_41, key_b_r_16_42, 
       key_b_r_16_43, key_b_r_16_44, key_b_r_16_45, key_b_r_16_46, key_b_r_16_47, key_b_r_16_48, key_b_r_16_49, key_b_r_16_5, key_b_r_16_50, 
       key_b_r_16_51, key_b_r_16_52, key_b_r_16_53, key_b_r_16_54, key_b_r_16_55, key_b_r_16_6, key_b_r_16_7, key_b_r_16_8, key_b_r_16_9, 
       key_b_r_1_0, key_b_r_1_1, key_b_r_1_10, key_b_r_1_11, key_b_r_1_12, key_b_r_1_13, key_b_r_1_14, key_b_r_1_15, key_b_r_1_16, 
       key_b_r_1_17, key_b_r_1_18, key_b_r_1_19, key_b_r_1_2, key_b_r_1_20, key_b_r_1_21, key_b_r_1_22, key_b_r_1_23, key_b_r_1_24, 
       key_b_r_1_25, key_b_r_1_26, key_b_r_1_27, key_b_r_1_28, key_b_r_1_29, key_b_r_1_3, key_b_r_1_30, key_b_r_1_31, key_b_r_1_32, 
       key_b_r_1_33, key_b_r_1_34, key_b_r_1_35, key_b_r_1_36, key_b_r_1_37, key_b_r_1_38, key_b_r_1_39, key_b_r_1_4, key_b_r_1_40, 
       key_b_r_1_41, key_b_r_1_42, key_b_r_1_43, key_b_r_1_44, key_b_r_1_45, key_b_r_1_46, key_b_r_1_47, key_b_r_1_48, key_b_r_1_49, 
       key_b_r_1_5, key_b_r_1_50, key_b_r_1_51, key_b_r_1_52, key_b_r_1_53, key_b_r_1_54, key_b_r_1_55, key_b_r_1_6, key_b_r_1_7, 
       key_b_r_1_8, key_b_r_1_9, key_b_r_2_0, key_b_r_2_1, key_b_r_2_10, key_b_r_2_11, key_b_r_2_12, key_b_r_2_13, key_b_r_2_14, 
       key_b_r_2_15, key_b_r_2_16, key_b_r_2_17, key_b_r_2_18, key_b_r_2_19, key_b_r_2_2, key_b_r_2_20, key_b_r_2_21, key_b_r_2_22, 
       key_b_r_2_23, key_b_r_2_24, key_b_r_2_25, key_b_r_2_26, key_b_r_2_27, key_b_r_2_28, key_b_r_2_29, key_b_r_2_3, key_b_r_2_30, 
       key_b_r_2_31, key_b_r_2_32, key_b_r_2_33, key_b_r_2_34, key_b_r_2_35, key_b_r_2_36, key_b_r_2_37, key_b_r_2_38, key_b_r_2_39, 
       key_b_r_2_4, key_b_r_2_40, key_b_r_2_41, key_b_r_2_42, key_b_r_2_43, key_b_r_2_44, key_b_r_2_45, key_b_r_2_46, key_b_r_2_47, 
       key_b_r_2_48, key_b_r_2_49, key_b_r_2_5, key_b_r_2_50, key_b_r_2_51, key_b_r_2_52, key_b_r_2_53, key_b_r_2_54, key_b_r_2_55, 
       key_b_r_2_6, key_b_r_2_7, key_b_r_2_8, key_b_r_2_9, key_b_r_3_0, key_b_r_3_1, key_b_r_3_10, key_b_r_3_11, key_b_r_3_12, 
       key_b_r_3_13, key_b_r_3_14, key_b_r_3_15, key_b_r_3_16, key_b_r_3_17, key_b_r_3_18, key_b_r_3_19, key_b_r_3_2, key_b_r_3_20, 
       key_b_r_3_21, key_b_r_3_22, key_b_r_3_23, key_b_r_3_24, key_b_r_3_25, key_b_r_3_26, key_b_r_3_27, key_b_r_3_28, key_b_r_3_29, 
       key_b_r_3_3, key_b_r_3_30, key_b_r_3_31, key_b_r_3_32, key_b_r_3_33, key_b_r_3_34, key_b_r_3_35, key_b_r_3_36, key_b_r_3_37, 
       key_b_r_3_38, key_b_r_3_39, key_b_r_3_4, key_b_r_3_40, key_b_r_3_41, key_b_r_3_42, key_b_r_3_43, key_b_r_3_44, key_b_r_3_45, 
       key_b_r_3_46, key_b_r_3_47, key_b_r_3_48, key_b_r_3_49, key_b_r_3_5, key_b_r_3_50, key_b_r_3_51, key_b_r_3_52, key_b_r_3_53, 
       key_b_r_3_54, key_b_r_3_55, key_b_r_3_6, key_b_r_3_7, key_b_r_3_8, key_b_r_3_9, key_b_r_4_0, key_b_r_4_1, key_b_r_4_10, 
       key_b_r_4_11, key_b_r_4_12, key_b_r_4_13, key_b_r_4_14, key_b_r_4_15, key_b_r_4_16, key_b_r_4_17, key_b_r_4_18, key_b_r_4_19, 
       key_b_r_4_2, key_b_r_4_20, key_b_r_4_21, key_b_r_4_22, key_b_r_4_23, key_b_r_4_24, key_b_r_4_25, key_b_r_4_26, key_b_r_4_27, 
       key_b_r_4_28, key_b_r_4_29, key_b_r_4_3, key_b_r_4_30, key_b_r_4_31, key_b_r_4_32, key_b_r_4_33, key_b_r_4_34, key_b_r_4_35, 
       key_b_r_4_36, key_b_r_4_37, key_b_r_4_38, key_b_r_4_39, key_b_r_4_4, key_b_r_4_40, key_b_r_4_41, key_b_r_4_42, key_b_r_4_43, 
       key_b_r_4_44, key_b_r_4_45, key_b_r_4_46, key_b_r_4_47, key_b_r_4_48, key_b_r_4_49, key_b_r_4_5, key_b_r_4_50, key_b_r_4_51, 
       key_b_r_4_52, key_b_r_4_53, key_b_r_4_54, key_b_r_4_55, key_b_r_4_6, key_b_r_4_7, key_b_r_4_8, key_b_r_4_9, key_b_r_5_0, 
       key_b_r_5_1, key_b_r_5_10, key_b_r_5_11, key_b_r_5_12, key_b_r_5_13, key_b_r_5_14, key_b_r_5_15, key_b_r_5_16, key_b_r_5_17, 
       key_b_r_5_18, key_b_r_5_19, key_b_r_5_2, key_b_r_5_20, key_b_r_5_21, key_b_r_5_22, key_b_r_5_23, key_b_r_5_24, key_b_r_5_25, 
       key_b_r_5_26, key_b_r_5_27, key_b_r_5_28, key_b_r_5_29, key_b_r_5_3, key_b_r_5_30, key_b_r_5_31, key_b_r_5_32, key_b_r_5_33, 
       key_b_r_5_34, key_b_r_5_35, key_b_r_5_36, key_b_r_5_37, key_b_r_5_38, key_b_r_5_39, key_b_r_5_4, key_b_r_5_40, key_b_r_5_41, 
       key_b_r_5_42, key_b_r_5_43, key_b_r_5_44, key_b_r_5_45, key_b_r_5_46, key_b_r_5_47, key_b_r_5_48, key_b_r_5_49, key_b_r_5_5, 
       key_b_r_5_50, key_b_r_5_51, key_b_r_5_52, key_b_r_5_53, key_b_r_5_54, key_b_r_5_55, key_b_r_5_6, key_b_r_5_7, key_b_r_5_8, 
       key_b_r_5_9, key_b_r_6_0, key_b_r_6_1, key_b_r_6_10, key_b_r_6_11, key_b_r_6_12, key_b_r_6_13, key_b_r_6_14, key_b_r_6_15, 
       key_b_r_6_16, key_b_r_6_17, key_b_r_6_18, key_b_r_6_19, key_b_r_6_2, key_b_r_6_20, key_b_r_6_21, key_b_r_6_22, key_b_r_6_23, 
       key_b_r_6_24, key_b_r_6_25, key_b_r_6_26, key_b_r_6_27, key_b_r_6_28, key_b_r_6_29, key_b_r_6_3, key_b_r_6_30, key_b_r_6_31, 
       key_b_r_6_32, key_b_r_6_33, key_b_r_6_34, key_b_r_6_35, key_b_r_6_36, key_b_r_6_37, key_b_r_6_38, key_b_r_6_39, key_b_r_6_4, 
       key_b_r_6_40, key_b_r_6_41, key_b_r_6_42, key_b_r_6_43, key_b_r_6_44, key_b_r_6_45, key_b_r_6_46, key_b_r_6_47, key_b_r_6_48, 
       key_b_r_6_49, key_b_r_6_5, key_b_r_6_50, key_b_r_6_51, key_b_r_6_52, key_b_r_6_53, key_b_r_6_54, key_b_r_6_55, key_b_r_6_6, 
       key_b_r_6_7, key_b_r_6_8, key_b_r_6_9, key_b_r_7_0, key_b_r_7_1, key_b_r_7_10, key_b_r_7_11, key_b_r_7_12, key_b_r_7_13, 
       key_b_r_7_14, key_b_r_7_15, key_b_r_7_16, key_b_r_7_17, key_b_r_7_18, key_b_r_7_19, key_b_r_7_2, key_b_r_7_20, key_b_r_7_21, 
       key_b_r_7_22, key_b_r_7_23, key_b_r_7_24, key_b_r_7_25, key_b_r_7_26, key_b_r_7_27, key_b_r_7_28, key_b_r_7_29, key_b_r_7_3, 
       key_b_r_7_30, key_b_r_7_31, key_b_r_7_32, key_b_r_7_33, key_b_r_7_34, key_b_r_7_35, key_b_r_7_36, key_b_r_7_37, key_b_r_7_38, 
       key_b_r_7_39, key_b_r_7_4, key_b_r_7_40, key_b_r_7_41, key_b_r_7_42, key_b_r_7_43, key_b_r_7_44, key_b_r_7_45, key_b_r_7_46, 
       key_b_r_7_47, key_b_r_7_48, key_b_r_7_49, key_b_r_7_5, key_b_r_7_50, key_b_r_7_51, key_b_r_7_52, key_b_r_7_53, key_b_r_7_54, 
       key_b_r_7_55, key_b_r_7_6, key_b_r_7_7, key_b_r_7_8, key_b_r_7_9, key_b_r_8_0, key_b_r_8_1, key_b_r_8_10, key_b_r_8_11, 
       key_b_r_8_12, key_b_r_8_13, key_b_r_8_14, key_b_r_8_15, key_b_r_8_16, key_b_r_8_17, key_b_r_8_18, key_b_r_8_19, key_b_r_8_2, 
       key_b_r_8_20, key_b_r_8_21, key_b_r_8_22, key_b_r_8_23, key_b_r_8_24, key_b_r_8_25, key_b_r_8_26, key_b_r_8_27, key_b_r_8_28, 
       key_b_r_8_29, key_b_r_8_3, key_b_r_8_30, key_b_r_8_31, key_b_r_8_32, key_b_r_8_33, key_b_r_8_34, key_b_r_8_35, key_b_r_8_36, 
       key_b_r_8_37, key_b_r_8_38, key_b_r_8_39, key_b_r_8_4, key_b_r_8_40, key_b_r_8_41, key_b_r_8_42, key_b_r_8_43, key_b_r_8_44, 
       key_b_r_8_45, key_b_r_8_46, key_b_r_8_47, key_b_r_8_48, key_b_r_8_49, key_b_r_8_5, key_b_r_8_50, key_b_r_8_51, key_b_r_8_52, 
       key_b_r_8_53, key_b_r_8_54, key_b_r_8_55, key_b_r_8_6, key_b_r_8_7, key_b_r_8_8, key_b_r_8_9, key_b_r_9_0, key_b_r_9_1, 
       key_b_r_9_10, key_b_r_9_11, key_b_r_9_12, key_b_r_9_13, key_b_r_9_14, key_b_r_9_15, key_b_r_9_16, key_b_r_9_17, key_b_r_9_18, 
       key_b_r_9_19, key_b_r_9_2, key_b_r_9_20, key_b_r_9_21, key_b_r_9_22, key_b_r_9_23, key_b_r_9_24, key_b_r_9_25, key_b_r_9_26, 
       key_b_r_9_27, key_b_r_9_28, key_b_r_9_29, key_b_r_9_3, key_b_r_9_30, key_b_r_9_31, key_b_r_9_32, key_b_r_9_33, key_b_r_9_34, 
       key_b_r_9_35, key_b_r_9_36, key_b_r_9_37, key_b_r_9_38, key_b_r_9_39, key_b_r_9_4, key_b_r_9_40, key_b_r_9_41, key_b_r_9_42, 
       key_b_r_9_43, key_b_r_9_44, key_b_r_9_45, key_b_r_9_46, key_b_r_9_47, key_b_r_9_48, key_b_r_9_49, key_b_r_9_5, key_b_r_9_50, 
       key_b_r_9_51, key_b_r_9_52, key_b_r_9_53, key_b_r_9_54, key_b_r_9_55, key_b_r_9_6, key_b_r_9_7, key_b_r_9_8, key_b_r_9_9, 
       key_c_r_0_0, key_c_r_0_1, key_c_r_0_10, key_c_r_0_11, key_c_r_0_12, key_c_r_0_13, key_c_r_0_14, key_c_r_0_15, key_c_r_0_16, 
       key_c_r_0_17, key_c_r_0_18, key_c_r_0_19, key_c_r_0_2, key_c_r_0_20, key_c_r_0_21, key_c_r_0_22, key_c_r_0_23, key_c_r_0_24, 
       key_c_r_0_25, key_c_r_0_26, key_c_r_0_27, key_c_r_0_28, key_c_r_0_29, key_c_r_0_3, key_c_r_0_30, key_c_r_0_31, key_c_r_0_32, 
       key_c_r_0_33, key_c_r_0_34, key_c_r_0_35, key_c_r_0_36, key_c_r_0_37, key_c_r_0_38, key_c_r_0_39, key_c_r_0_4, key_c_r_0_40, 
       key_c_r_0_41, key_c_r_0_42, key_c_r_0_43, key_c_r_0_44, key_c_r_0_45, key_c_r_0_46, key_c_r_0_47, key_c_r_0_48, key_c_r_0_49, 
       key_c_r_0_5, key_c_r_0_50, key_c_r_0_51, key_c_r_0_52, key_c_r_0_53, key_c_r_0_54, key_c_r_0_55, key_c_r_0_6, key_c_r_0_7, 
       key_c_r_0_8, key_c_r_0_9, key_c_r_10_0, key_c_r_10_1, key_c_r_10_10, key_c_r_10_11, key_c_r_10_12, key_c_r_10_13, key_c_r_10_14, 
       key_c_r_10_15, key_c_r_10_16, key_c_r_10_17, key_c_r_10_18, key_c_r_10_19, key_c_r_10_2, key_c_r_10_20, key_c_r_10_21, key_c_r_10_22, 
       key_c_r_10_23, key_c_r_10_24, key_c_r_10_25, key_c_r_10_26, key_c_r_10_27, key_c_r_10_28, key_c_r_10_29, key_c_r_10_3, key_c_r_10_30, 
       key_c_r_10_31, key_c_r_10_32, key_c_r_10_33, key_c_r_10_34, key_c_r_10_35, key_c_r_10_36, key_c_r_10_37, key_c_r_10_38, key_c_r_10_39, 
       key_c_r_10_4, key_c_r_10_40, key_c_r_10_41, key_c_r_10_42, key_c_r_10_43, key_c_r_10_44, key_c_r_10_45, key_c_r_10_46, key_c_r_10_47, 
       key_c_r_10_48, key_c_r_10_49, key_c_r_10_5, key_c_r_10_50, key_c_r_10_51, key_c_r_10_52, key_c_r_10_53, key_c_r_10_54, key_c_r_10_55, 
       key_c_r_10_6, key_c_r_10_7, key_c_r_10_8, key_c_r_10_9, key_c_r_11_0, key_c_r_11_1, key_c_r_11_10, key_c_r_11_11, key_c_r_11_12, 
       key_c_r_11_13, key_c_r_11_14, key_c_r_11_15, key_c_r_11_16, key_c_r_11_17, key_c_r_11_18, key_c_r_11_19, key_c_r_11_2, key_c_r_11_20, 
       key_c_r_11_21, key_c_r_11_22, key_c_r_11_23, key_c_r_11_24, key_c_r_11_25, key_c_r_11_26, key_c_r_11_27, key_c_r_11_28, key_c_r_11_29, 
       key_c_r_11_3, key_c_r_11_30, key_c_r_11_31, key_c_r_11_32, key_c_r_11_33, key_c_r_11_34, key_c_r_11_35, key_c_r_11_36, key_c_r_11_37, 
       key_c_r_11_38, key_c_r_11_39, key_c_r_11_4, key_c_r_11_40, key_c_r_11_41, key_c_r_11_42, key_c_r_11_43, key_c_r_11_44, key_c_r_11_45, 
       key_c_r_11_46, key_c_r_11_47, key_c_r_11_48, key_c_r_11_49, key_c_r_11_5, key_c_r_11_50, key_c_r_11_51, key_c_r_11_52, key_c_r_11_53, 
       key_c_r_11_54, key_c_r_11_55, key_c_r_11_6, key_c_r_11_7, key_c_r_11_8, key_c_r_11_9, key_c_r_12_0, key_c_r_12_1, key_c_r_12_10, 
       key_c_r_12_11, key_c_r_12_12, key_c_r_12_13, key_c_r_12_14, key_c_r_12_15, key_c_r_12_16, key_c_r_12_17, key_c_r_12_18, key_c_r_12_19, 
       key_c_r_12_2, key_c_r_12_20, key_c_r_12_21, key_c_r_12_22, key_c_r_12_23, key_c_r_12_24, key_c_r_12_25, key_c_r_12_26, key_c_r_12_27, 
       key_c_r_12_28, key_c_r_12_29, key_c_r_12_3, key_c_r_12_30, key_c_r_12_31, key_c_r_12_32, key_c_r_12_33, key_c_r_12_34, key_c_r_12_35, 
       key_c_r_12_36, key_c_r_12_37, key_c_r_12_38, key_c_r_12_39, key_c_r_12_4, key_c_r_12_40, key_c_r_12_41, key_c_r_12_42, key_c_r_12_43, 
       key_c_r_12_44, key_c_r_12_45, key_c_r_12_46, key_c_r_12_47, key_c_r_12_48, key_c_r_12_49, key_c_r_12_5, key_c_r_12_50, key_c_r_12_51, 
       key_c_r_12_52, key_c_r_12_53, key_c_r_12_54, key_c_r_12_55, key_c_r_12_6, key_c_r_12_7, key_c_r_12_8, key_c_r_12_9, key_c_r_13_0, 
       key_c_r_13_1, key_c_r_13_10, key_c_r_13_11, key_c_r_13_12, key_c_r_13_13, key_c_r_13_14, key_c_r_13_15, key_c_r_13_16, key_c_r_13_17, 
       key_c_r_13_18, key_c_r_13_19, key_c_r_13_2, key_c_r_13_20, key_c_r_13_21, key_c_r_13_22, key_c_r_13_23, key_c_r_13_24, key_c_r_13_25, 
       key_c_r_13_26, key_c_r_13_27, key_c_r_13_28, key_c_r_13_29, key_c_r_13_3, key_c_r_13_30, key_c_r_13_31, key_c_r_13_32, key_c_r_13_33, 
       key_c_r_13_34, key_c_r_13_35, key_c_r_13_36, key_c_r_13_37, key_c_r_13_38, key_c_r_13_39, key_c_r_13_4, key_c_r_13_40, key_c_r_13_41, 
       key_c_r_13_42, key_c_r_13_43, key_c_r_13_44, key_c_r_13_45, key_c_r_13_46, key_c_r_13_47, key_c_r_13_48, key_c_r_13_49, key_c_r_13_5, 
       key_c_r_13_50, key_c_r_13_51, key_c_r_13_52, key_c_r_13_53, key_c_r_13_54, key_c_r_13_55, key_c_r_13_6, key_c_r_13_7, key_c_r_13_8, 
       key_c_r_13_9, key_c_r_14_0, key_c_r_14_1, key_c_r_14_10, key_c_r_14_11, key_c_r_14_12, key_c_r_14_13, key_c_r_14_14, key_c_r_14_15, 
       key_c_r_14_16, key_c_r_14_17, key_c_r_14_18, key_c_r_14_19, key_c_r_14_2, key_c_r_14_20, key_c_r_14_21, key_c_r_14_22, key_c_r_14_23, 
       key_c_r_14_24, key_c_r_14_25, key_c_r_14_26, key_c_r_14_27, key_c_r_14_28, key_c_r_14_29, key_c_r_14_3, key_c_r_14_30, key_c_r_14_31, 
       key_c_r_14_32, key_c_r_14_33, key_c_r_14_34, key_c_r_14_35, key_c_r_14_36, key_c_r_14_37, key_c_r_14_38, key_c_r_14_39, key_c_r_14_4, 
       key_c_r_14_40, key_c_r_14_41, key_c_r_14_42, key_c_r_14_43, key_c_r_14_44, key_c_r_14_45, key_c_r_14_46, key_c_r_14_47, key_c_r_14_48, 
       key_c_r_14_49, key_c_r_14_5, key_c_r_14_50, key_c_r_14_51, key_c_r_14_52, key_c_r_14_53, key_c_r_14_54, key_c_r_14_55, key_c_r_14_6, 
       key_c_r_14_7, key_c_r_14_8, key_c_r_14_9, key_c_r_15_0, key_c_r_15_1, key_c_r_15_10, key_c_r_15_11, key_c_r_15_12, key_c_r_15_13, 
       key_c_r_15_14, key_c_r_15_15, key_c_r_15_16, key_c_r_15_17, key_c_r_15_18, key_c_r_15_19, key_c_r_15_2, key_c_r_15_20, key_c_r_15_21, 
       key_c_r_15_22, key_c_r_15_23, key_c_r_15_24, key_c_r_15_25, key_c_r_15_26, key_c_r_15_27, key_c_r_15_28, key_c_r_15_29, key_c_r_15_3, 
       key_c_r_15_30, key_c_r_15_31, key_c_r_15_32, key_c_r_15_33, key_c_r_15_34, key_c_r_15_35, key_c_r_15_36, key_c_r_15_37, key_c_r_15_38, 
       key_c_r_15_39, key_c_r_15_4, key_c_r_15_40, key_c_r_15_41, key_c_r_15_42, key_c_r_15_43, key_c_r_15_44, key_c_r_15_45, key_c_r_15_46, 
       key_c_r_15_47, key_c_r_15_48, key_c_r_15_49, key_c_r_15_5, key_c_r_15_50, key_c_r_15_51, key_c_r_15_52, key_c_r_15_53, key_c_r_15_54, 
       key_c_r_15_55, key_c_r_15_6, key_c_r_15_7, key_c_r_15_8, key_c_r_15_9, key_c_r_16_0, key_c_r_16_1, key_c_r_16_10, key_c_r_16_11, 
       key_c_r_16_12, key_c_r_16_13, key_c_r_16_14, key_c_r_16_15, key_c_r_16_16, key_c_r_16_17, key_c_r_16_18, key_c_r_16_19, key_c_r_16_2, 
       key_c_r_16_20, key_c_r_16_21, key_c_r_16_22, key_c_r_16_23, key_c_r_16_24, key_c_r_16_25, key_c_r_16_26, key_c_r_16_27, key_c_r_16_28, 
       key_c_r_16_29, key_c_r_16_3, key_c_r_16_30, key_c_r_16_31, key_c_r_16_32, key_c_r_16_33, key_c_r_16_34, key_c_r_16_35, key_c_r_16_36, 
       key_c_r_16_37, key_c_r_16_38, key_c_r_16_39, key_c_r_16_4, key_c_r_16_40, key_c_r_16_41, key_c_r_16_42, key_c_r_16_43, key_c_r_16_44, 
       key_c_r_16_45, key_c_r_16_46, key_c_r_16_47, key_c_r_16_48, key_c_r_16_49, key_c_r_16_5, key_c_r_16_50, key_c_r_16_51, key_c_r_16_52, 
       key_c_r_16_53, key_c_r_16_54, key_c_r_16_55, key_c_r_16_6, key_c_r_16_7, key_c_r_16_8, key_c_r_16_9, key_c_r_17_0, key_c_r_17_1, 
       key_c_r_17_10, key_c_r_17_11, key_c_r_17_12, key_c_r_17_13, key_c_r_17_14, key_c_r_17_15, key_c_r_17_16, key_c_r_17_17, key_c_r_17_18, 
       key_c_r_17_19, key_c_r_17_2, key_c_r_17_20, key_c_r_17_21, key_c_r_17_22, key_c_r_17_23, key_c_r_17_24, key_c_r_17_25, key_c_r_17_26, 
       key_c_r_17_27, key_c_r_17_28, key_c_r_17_29, key_c_r_17_3, key_c_r_17_30, key_c_r_17_31, key_c_r_17_32, key_c_r_17_33, key_c_r_17_34, 
       key_c_r_17_35, key_c_r_17_36, key_c_r_17_37, key_c_r_17_38, key_c_r_17_39, key_c_r_17_4, key_c_r_17_40, key_c_r_17_41, key_c_r_17_42, 
       key_c_r_17_43, key_c_r_17_44, key_c_r_17_45, key_c_r_17_46, key_c_r_17_47, key_c_r_17_48, key_c_r_17_49, key_c_r_17_5, key_c_r_17_50, 
       key_c_r_17_51, key_c_r_17_52, key_c_r_17_53, key_c_r_17_54, key_c_r_17_55, key_c_r_17_6, key_c_r_17_7, key_c_r_17_8, key_c_r_17_9, 
       key_c_r_18_0, key_c_r_18_1, key_c_r_18_10, key_c_r_18_11, key_c_r_18_12, key_c_r_18_13, key_c_r_18_14, key_c_r_18_15, key_c_r_18_16, 
       key_c_r_18_17, key_c_r_18_18, key_c_r_18_19, key_c_r_18_2, key_c_r_18_20, key_c_r_18_21, key_c_r_18_22, key_c_r_18_23, key_c_r_18_24, 
       key_c_r_18_25, key_c_r_18_26, key_c_r_18_27, key_c_r_18_28, key_c_r_18_29, key_c_r_18_3, key_c_r_18_30, key_c_r_18_31, key_c_r_18_32, 
       key_c_r_18_33, key_c_r_18_34, key_c_r_18_35, key_c_r_18_36, key_c_r_18_37, key_c_r_18_38, key_c_r_18_39, key_c_r_18_4, key_c_r_18_40, 
       key_c_r_18_41, key_c_r_18_42, key_c_r_18_43, key_c_r_18_44, key_c_r_18_45, key_c_r_18_46, key_c_r_18_47, key_c_r_18_48, key_c_r_18_49, 
       key_c_r_18_5, key_c_r_18_50, key_c_r_18_51, key_c_r_18_52, key_c_r_18_53, key_c_r_18_54, key_c_r_18_55, key_c_r_18_6, key_c_r_18_7, 
       key_c_r_18_8, key_c_r_18_9, key_c_r_19_0, key_c_r_19_1, key_c_r_19_10, key_c_r_19_11, key_c_r_19_12, key_c_r_19_13, key_c_r_19_14, 
       key_c_r_19_15, key_c_r_19_16, key_c_r_19_17, key_c_r_19_18, key_c_r_19_19, key_c_r_19_2, key_c_r_19_20, key_c_r_19_21, key_c_r_19_22, 
       key_c_r_19_23, key_c_r_19_24, key_c_r_19_25, key_c_r_19_26, key_c_r_19_27, key_c_r_19_28, key_c_r_19_29, key_c_r_19_3, key_c_r_19_30, 
       key_c_r_19_31, key_c_r_19_32, key_c_r_19_33, key_c_r_19_34, key_c_r_19_35, key_c_r_19_36, key_c_r_19_37, key_c_r_19_38, key_c_r_19_39, 
       key_c_r_19_4, key_c_r_19_40, key_c_r_19_41, key_c_r_19_42, key_c_r_19_43, key_c_r_19_44, key_c_r_19_45, key_c_r_19_46, key_c_r_19_47, 
       key_c_r_19_48, key_c_r_19_49, key_c_r_19_5, key_c_r_19_50, key_c_r_19_51, key_c_r_19_52, key_c_r_19_53, key_c_r_19_54, key_c_r_19_55, 
       key_c_r_19_6, key_c_r_19_7, key_c_r_19_8, key_c_r_19_9, key_c_r_1_0, key_c_r_1_1, key_c_r_1_10, key_c_r_1_11, key_c_r_1_12, 
       key_c_r_1_13, key_c_r_1_14, key_c_r_1_15, key_c_r_1_16, key_c_r_1_17, key_c_r_1_18, key_c_r_1_19, key_c_r_1_2, key_c_r_1_20, 
       key_c_r_1_21, key_c_r_1_22, key_c_r_1_23, key_c_r_1_24, key_c_r_1_25, key_c_r_1_26, key_c_r_1_27, key_c_r_1_28, key_c_r_1_29, 
       key_c_r_1_3, key_c_r_1_30, key_c_r_1_31, key_c_r_1_32, key_c_r_1_33, key_c_r_1_34, key_c_r_1_35, key_c_r_1_36, key_c_r_1_37, 
       key_c_r_1_38, key_c_r_1_39, key_c_r_1_4, key_c_r_1_40, key_c_r_1_41, key_c_r_1_42, key_c_r_1_43, key_c_r_1_44, key_c_r_1_45, 
       key_c_r_1_46, key_c_r_1_47, key_c_r_1_48, key_c_r_1_49, key_c_r_1_5, key_c_r_1_50, key_c_r_1_51, key_c_r_1_52, key_c_r_1_53, 
       key_c_r_1_54, key_c_r_1_55, key_c_r_1_6, key_c_r_1_7, key_c_r_1_8, key_c_r_1_9, key_c_r_20_0, key_c_r_20_1, key_c_r_20_10, 
       key_c_r_20_11, key_c_r_20_12, key_c_r_20_13, key_c_r_20_14, key_c_r_20_15, key_c_r_20_16, key_c_r_20_17, key_c_r_20_18, key_c_r_20_19, 
       key_c_r_20_2, key_c_r_20_20, key_c_r_20_21, key_c_r_20_22, key_c_r_20_23, key_c_r_20_24, key_c_r_20_25, key_c_r_20_26, key_c_r_20_27, 
       key_c_r_20_28, key_c_r_20_29, key_c_r_20_3, key_c_r_20_30, key_c_r_20_31, key_c_r_20_32, key_c_r_20_33, key_c_r_20_34, key_c_r_20_35, 
       key_c_r_20_36, key_c_r_20_37, key_c_r_20_38, key_c_r_20_39, key_c_r_20_4, key_c_r_20_40, key_c_r_20_41, key_c_r_20_42, key_c_r_20_43, 
       key_c_r_20_44, key_c_r_20_45, key_c_r_20_46, key_c_r_20_47, key_c_r_20_48, key_c_r_20_49, key_c_r_20_5, key_c_r_20_50, key_c_r_20_51, 
       key_c_r_20_52, key_c_r_20_53, key_c_r_20_54, key_c_r_20_55, key_c_r_20_6, key_c_r_20_7, key_c_r_20_8, key_c_r_20_9, key_c_r_21_0, 
       key_c_r_21_1, key_c_r_21_10, key_c_r_21_11, key_c_r_21_12, key_c_r_21_13, key_c_r_21_14, key_c_r_21_15, key_c_r_21_16, key_c_r_21_17, 
       key_c_r_21_18, key_c_r_21_19, key_c_r_21_2, key_c_r_21_20, key_c_r_21_21, key_c_r_21_22, key_c_r_21_23, key_c_r_21_24, key_c_r_21_25, 
       key_c_r_21_26, key_c_r_21_27, key_c_r_21_28, key_c_r_21_29, key_c_r_21_3, key_c_r_21_30, key_c_r_21_31, key_c_r_21_32, key_c_r_21_33, 
       key_c_r_21_34, key_c_r_21_35, key_c_r_21_36, key_c_r_21_37, key_c_r_21_38, key_c_r_21_39, key_c_r_21_4, key_c_r_21_40, key_c_r_21_41, 
       key_c_r_21_42, key_c_r_21_43, key_c_r_21_44, key_c_r_21_45, key_c_r_21_46, key_c_r_21_47, key_c_r_21_48, key_c_r_21_49, key_c_r_21_5, 
       key_c_r_21_50, key_c_r_21_51, key_c_r_21_52, key_c_r_21_53, key_c_r_21_54, key_c_r_21_55, key_c_r_21_6, key_c_r_21_7, key_c_r_21_8, 
       key_c_r_21_9, key_c_r_22_0, key_c_r_22_1, key_c_r_22_10, key_c_r_22_11, key_c_r_22_12, key_c_r_22_13, key_c_r_22_14, key_c_r_22_15, 
       key_c_r_22_16, key_c_r_22_17, key_c_r_22_18, key_c_r_22_19, key_c_r_22_2, key_c_r_22_20, key_c_r_22_21, key_c_r_22_22, key_c_r_22_23, 
       key_c_r_22_24, key_c_r_22_25, key_c_r_22_26, key_c_r_22_27, key_c_r_22_28, key_c_r_22_29, key_c_r_22_3, key_c_r_22_30, key_c_r_22_31, 
       key_c_r_22_32, key_c_r_22_33, key_c_r_22_34, key_c_r_22_35, key_c_r_22_36, key_c_r_22_37, key_c_r_22_38, key_c_r_22_39, key_c_r_22_4, 
       key_c_r_22_40, key_c_r_22_41, key_c_r_22_42, key_c_r_22_43, key_c_r_22_44, key_c_r_22_45, key_c_r_22_46, key_c_r_22_47, key_c_r_22_48, 
       key_c_r_22_49, key_c_r_22_5, key_c_r_22_50, key_c_r_22_51, key_c_r_22_52, key_c_r_22_53, key_c_r_22_54, key_c_r_22_55, key_c_r_22_6, 
       key_c_r_22_7, key_c_r_22_8, key_c_r_22_9, key_c_r_23_0, key_c_r_23_1, key_c_r_23_10, key_c_r_23_11, key_c_r_23_12, key_c_r_23_13, 
       key_c_r_23_14, key_c_r_23_15, key_c_r_23_16, key_c_r_23_17, key_c_r_23_18, key_c_r_23_19, key_c_r_23_2, key_c_r_23_20, key_c_r_23_21, 
       key_c_r_23_22, key_c_r_23_23, key_c_r_23_24, key_c_r_23_25, key_c_r_23_26, key_c_r_23_27, key_c_r_23_28, key_c_r_23_29, key_c_r_23_3, 
       key_c_r_23_30, key_c_r_23_31, key_c_r_23_32, key_c_r_23_33, key_c_r_23_34, key_c_r_23_35, key_c_r_23_36, key_c_r_23_37, key_c_r_23_38, 
       key_c_r_23_39, key_c_r_23_4, key_c_r_23_40, key_c_r_23_41, key_c_r_23_42, key_c_r_23_43, key_c_r_23_44, key_c_r_23_45, key_c_r_23_46, 
       key_c_r_23_47, key_c_r_23_48, key_c_r_23_49, key_c_r_23_5, key_c_r_23_50, key_c_r_23_51, key_c_r_23_52, key_c_r_23_53, key_c_r_23_54, 
       key_c_r_23_55, key_c_r_23_6, key_c_r_23_7, key_c_r_23_8, key_c_r_23_9, key_c_r_24_0, key_c_r_24_1, key_c_r_24_10, key_c_r_24_11, 
       key_c_r_24_12, key_c_r_24_13, key_c_r_24_14, key_c_r_24_15, key_c_r_24_16, key_c_r_24_17, key_c_r_24_18, key_c_r_24_19, key_c_r_24_2, 
       key_c_r_24_20, key_c_r_24_21, key_c_r_24_22, key_c_r_24_23, key_c_r_24_24, key_c_r_24_25, key_c_r_24_26, key_c_r_24_27, key_c_r_24_28, 
       key_c_r_24_29, key_c_r_24_3, key_c_r_24_30, key_c_r_24_31, key_c_r_24_32, key_c_r_24_33, key_c_r_24_34, key_c_r_24_35, key_c_r_24_36, 
       key_c_r_24_37, key_c_r_24_38, key_c_r_24_39, key_c_r_24_4, key_c_r_24_40, key_c_r_24_41, key_c_r_24_42, key_c_r_24_43, key_c_r_24_44, 
       key_c_r_24_45, key_c_r_24_46, key_c_r_24_47, key_c_r_24_48, key_c_r_24_49, key_c_r_24_5, key_c_r_24_50, key_c_r_24_51, key_c_r_24_52, 
       key_c_r_24_53, key_c_r_24_54, key_c_r_24_55, key_c_r_24_6, key_c_r_24_7, key_c_r_24_8, key_c_r_24_9, key_c_r_25_0, key_c_r_25_1, 
       key_c_r_25_10, key_c_r_25_11, key_c_r_25_12, key_c_r_25_13, key_c_r_25_14, key_c_r_25_15, key_c_r_25_16, key_c_r_25_17, key_c_r_25_18, 
       key_c_r_25_19, key_c_r_25_2, key_c_r_25_20, key_c_r_25_21, key_c_r_25_22, key_c_r_25_23, key_c_r_25_24, key_c_r_25_25, key_c_r_25_26, 
       key_c_r_25_27, key_c_r_25_28, key_c_r_25_29, key_c_r_25_3, key_c_r_25_30, key_c_r_25_31, key_c_r_25_32, key_c_r_25_33, key_c_r_25_34, 
       key_c_r_25_35, key_c_r_25_36, key_c_r_25_37, key_c_r_25_38, key_c_r_25_39, key_c_r_25_4, key_c_r_25_40, key_c_r_25_41, key_c_r_25_42, 
       key_c_r_25_43, key_c_r_25_44, key_c_r_25_45, key_c_r_25_46, key_c_r_25_47, key_c_r_25_48, key_c_r_25_49, key_c_r_25_5, key_c_r_25_50, 
       key_c_r_25_51, key_c_r_25_52, key_c_r_25_53, key_c_r_25_54, key_c_r_25_55, key_c_r_25_6, key_c_r_25_7, key_c_r_25_8, key_c_r_25_9, 
       key_c_r_26_0, key_c_r_26_1, key_c_r_26_10, key_c_r_26_11, key_c_r_26_12, key_c_r_26_13, key_c_r_26_14, key_c_r_26_15, key_c_r_26_16, 
       key_c_r_26_17, key_c_r_26_18, key_c_r_26_19, key_c_r_26_2, key_c_r_26_20, key_c_r_26_21, key_c_r_26_22, key_c_r_26_23, key_c_r_26_24, 
       key_c_r_26_25, key_c_r_26_26, key_c_r_26_27, key_c_r_26_28, key_c_r_26_29, key_c_r_26_3, key_c_r_26_30, key_c_r_26_31, key_c_r_26_32, 
       key_c_r_26_33, key_c_r_26_34, key_c_r_26_35, key_c_r_26_36, key_c_r_26_37, key_c_r_26_38, key_c_r_26_39, key_c_r_26_4, key_c_r_26_40, 
       key_c_r_26_41, key_c_r_26_42, key_c_r_26_43, key_c_r_26_44, key_c_r_26_45, key_c_r_26_46, key_c_r_26_47, key_c_r_26_48, key_c_r_26_49, 
       key_c_r_26_5, key_c_r_26_50, key_c_r_26_51, key_c_r_26_52, key_c_r_26_53, key_c_r_26_54, key_c_r_26_55, key_c_r_26_6, key_c_r_26_7, 
       key_c_r_26_8, key_c_r_26_9, key_c_r_27_0, key_c_r_27_1, key_c_r_27_10, key_c_r_27_11, key_c_r_27_12, key_c_r_27_13, key_c_r_27_14, 
       key_c_r_27_15, key_c_r_27_16, key_c_r_27_17, key_c_r_27_18, key_c_r_27_19, key_c_r_27_2, key_c_r_27_20, key_c_r_27_21, key_c_r_27_22, 
       key_c_r_27_23, key_c_r_27_24, key_c_r_27_25, key_c_r_27_26, key_c_r_27_27, key_c_r_27_28, key_c_r_27_29, key_c_r_27_3, key_c_r_27_30, 
       key_c_r_27_31, key_c_r_27_32, key_c_r_27_33, key_c_r_27_34, key_c_r_27_35, key_c_r_27_36, key_c_r_27_37, key_c_r_27_38, key_c_r_27_39, 
       key_c_r_27_4, key_c_r_27_40, key_c_r_27_41, key_c_r_27_42, key_c_r_27_43, key_c_r_27_44, key_c_r_27_45, key_c_r_27_46, key_c_r_27_47, 
       key_c_r_27_48, key_c_r_27_49, key_c_r_27_5, key_c_r_27_50, key_c_r_27_51, key_c_r_27_52, key_c_r_27_53, key_c_r_27_54, key_c_r_27_55, 
       key_c_r_27_6, key_c_r_27_7, key_c_r_27_8, key_c_r_27_9, key_c_r_28_0, key_c_r_28_1, key_c_r_28_10, key_c_r_28_11, key_c_r_28_12, 
       key_c_r_28_13, key_c_r_28_14, key_c_r_28_15, key_c_r_28_16, key_c_r_28_17, key_c_r_28_18, key_c_r_28_19, key_c_r_28_2, key_c_r_28_20, 
       key_c_r_28_21, key_c_r_28_22, key_c_r_28_23, key_c_r_28_24, key_c_r_28_25, key_c_r_28_26, key_c_r_28_27, key_c_r_28_28, key_c_r_28_29, 
       key_c_r_28_3, key_c_r_28_30, key_c_r_28_31, key_c_r_28_32, key_c_r_28_33, key_c_r_28_34, key_c_r_28_35, key_c_r_28_36, key_c_r_28_37, 
       key_c_r_28_38, key_c_r_28_39, key_c_r_28_4, key_c_r_28_40, key_c_r_28_41, key_c_r_28_42, key_c_r_28_43, key_c_r_28_44, key_c_r_28_45, 
       key_c_r_28_46, key_c_r_28_47, key_c_r_28_48, key_c_r_28_49, key_c_r_28_5, key_c_r_28_50, key_c_r_28_51, key_c_r_28_52, key_c_r_28_53, 
       key_c_r_28_54, key_c_r_28_55, key_c_r_28_6, key_c_r_28_7, key_c_r_28_8, key_c_r_28_9, key_c_r_29_0, key_c_r_29_1, key_c_r_29_10, 
       key_c_r_29_11, key_c_r_29_12, key_c_r_29_13, key_c_r_29_14, key_c_r_29_15, key_c_r_29_16, key_c_r_29_17, key_c_r_29_18, key_c_r_29_19, 
       key_c_r_29_2, key_c_r_29_20, key_c_r_29_21, key_c_r_29_22, key_c_r_29_23, key_c_r_29_24, key_c_r_29_25, key_c_r_29_26, key_c_r_29_27, 
       key_c_r_29_28, key_c_r_29_29, key_c_r_29_3, key_c_r_29_30, key_c_r_29_31, key_c_r_29_32, key_c_r_29_33, key_c_r_29_34, key_c_r_29_35, 
       key_c_r_29_36, key_c_r_29_37, key_c_r_29_38, key_c_r_29_39, key_c_r_29_4, key_c_r_29_40, key_c_r_29_41, key_c_r_29_42, key_c_r_29_43, 
       key_c_r_29_44, key_c_r_29_45, key_c_r_29_46, key_c_r_29_47, key_c_r_29_48, key_c_r_29_49, key_c_r_29_5, key_c_r_29_50, key_c_r_29_51, 
       key_c_r_29_52, key_c_r_29_53, key_c_r_29_54, key_c_r_29_55, key_c_r_29_6, key_c_r_29_7, key_c_r_29_8, key_c_r_29_9, key_c_r_2_0, 
       key_c_r_2_1, key_c_r_2_10, key_c_r_2_11, key_c_r_2_12, key_c_r_2_13, key_c_r_2_14, key_c_r_2_15, key_c_r_2_16, key_c_r_2_17, 
       key_c_r_2_18, key_c_r_2_19, key_c_r_2_2, key_c_r_2_20, key_c_r_2_21, key_c_r_2_22, key_c_r_2_23, key_c_r_2_24, key_c_r_2_25, 
       key_c_r_2_26, key_c_r_2_27, key_c_r_2_28, key_c_r_2_29, key_c_r_2_3, key_c_r_2_30, key_c_r_2_31, key_c_r_2_32, key_c_r_2_33, 
       key_c_r_2_34, key_c_r_2_35, key_c_r_2_36, key_c_r_2_37, key_c_r_2_38, key_c_r_2_39, key_c_r_2_4, key_c_r_2_40, key_c_r_2_41, 
       key_c_r_2_42, key_c_r_2_43, key_c_r_2_44, key_c_r_2_45, key_c_r_2_46, key_c_r_2_47, key_c_r_2_48, key_c_r_2_49, key_c_r_2_5, 
       key_c_r_2_50, key_c_r_2_51, key_c_r_2_52, key_c_r_2_53, key_c_r_2_54, key_c_r_2_55, key_c_r_2_6, key_c_r_2_7, key_c_r_2_8, 
       key_c_r_2_9, key_c_r_30_0, key_c_r_30_1, key_c_r_30_10, key_c_r_30_11, key_c_r_30_12, key_c_r_30_13, key_c_r_30_14, key_c_r_30_15, 
       key_c_r_30_16, key_c_r_30_17, key_c_r_30_18, key_c_r_30_19, key_c_r_30_2, key_c_r_30_20, key_c_r_30_21, key_c_r_30_22, key_c_r_30_23, 
       key_c_r_30_24, key_c_r_30_25, key_c_r_30_26, key_c_r_30_27, key_c_r_30_28, key_c_r_30_29, key_c_r_30_3, key_c_r_30_30, key_c_r_30_31, 
       key_c_r_30_32, key_c_r_30_33, key_c_r_30_34, key_c_r_30_35, key_c_r_30_36, key_c_r_30_37, key_c_r_30_38, key_c_r_30_39, key_c_r_30_4, 
       key_c_r_30_40, key_c_r_30_41, key_c_r_30_42, key_c_r_30_43, key_c_r_30_44, key_c_r_30_45, key_c_r_30_46, key_c_r_30_47, key_c_r_30_48, 
       key_c_r_30_49, key_c_r_30_5, key_c_r_30_50, key_c_r_30_51, key_c_r_30_52, key_c_r_30_53, key_c_r_30_54, key_c_r_30_55, key_c_r_30_6, 
       key_c_r_30_7, key_c_r_30_8, key_c_r_30_9, key_c_r_31_0, key_c_r_31_1, key_c_r_31_10, key_c_r_31_11, key_c_r_31_12, key_c_r_31_13, 
       key_c_r_31_14, key_c_r_31_15, key_c_r_31_16, key_c_r_31_17, key_c_r_31_18, key_c_r_31_19, key_c_r_31_2, key_c_r_31_20, key_c_r_31_21, 
       key_c_r_31_22, key_c_r_31_23, key_c_r_31_24, key_c_r_31_25, key_c_r_31_26, key_c_r_31_27, key_c_r_31_28, key_c_r_31_29, key_c_r_31_3, 
       key_c_r_31_30, key_c_r_31_31, key_c_r_31_32, key_c_r_31_33, key_c_r_31_34, key_c_r_31_35, key_c_r_31_36, key_c_r_31_37, key_c_r_31_38, 
       key_c_r_31_39, key_c_r_31_4, key_c_r_31_40, key_c_r_31_41, key_c_r_31_42, key_c_r_31_43, key_c_r_31_44, key_c_r_31_45, key_c_r_31_46, 
       key_c_r_31_47, key_c_r_31_48, key_c_r_31_49, key_c_r_31_5, key_c_r_31_50, key_c_r_31_51, key_c_r_31_52, key_c_r_31_53, key_c_r_31_54, 
       key_c_r_31_55, key_c_r_31_6, key_c_r_31_7, key_c_r_31_8, key_c_r_31_9, key_c_r_32_0, key_c_r_32_1, key_c_r_32_10, key_c_r_32_11, 
       key_c_r_32_12, key_c_r_32_13, key_c_r_32_14, key_c_r_32_15, key_c_r_32_16, key_c_r_32_17, key_c_r_32_18, key_c_r_32_19, key_c_r_32_2, 
       key_c_r_32_20, key_c_r_32_21, key_c_r_32_22, key_c_r_32_23, key_c_r_32_24, key_c_r_32_25, key_c_r_32_26, key_c_r_32_27, key_c_r_32_28, 
       key_c_r_32_29, key_c_r_32_3, key_c_r_32_30, key_c_r_32_31, key_c_r_32_32, key_c_r_32_33, key_c_r_32_34, key_c_r_32_35, key_c_r_32_36, 
       key_c_r_32_37, key_c_r_32_38, key_c_r_32_39, key_c_r_32_4, key_c_r_32_40, key_c_r_32_41, key_c_r_32_42, key_c_r_32_43, key_c_r_32_44, 
       key_c_r_32_45, key_c_r_32_46, key_c_r_32_47, key_c_r_32_48, key_c_r_32_49, key_c_r_32_5, key_c_r_32_50, key_c_r_32_51, key_c_r_32_52, 
       key_c_r_32_53, key_c_r_32_54, key_c_r_32_55, key_c_r_32_6, key_c_r_32_7, key_c_r_32_8, key_c_r_32_9, key_c_r_33_0, key_c_r_33_1, 
       key_c_r_33_10, key_c_r_33_11, key_c_r_33_12, key_c_r_33_13, key_c_r_33_14, key_c_r_33_15, key_c_r_33_16, key_c_r_33_17, key_c_r_33_18, 
       key_c_r_33_19, key_c_r_33_2, key_c_r_33_20, key_c_r_33_21, key_c_r_33_22, key_c_r_33_23, key_c_r_33_24, key_c_r_33_25, key_c_r_33_26, 
       key_c_r_33_27, key_c_r_33_28, key_c_r_33_29, key_c_r_33_3, key_c_r_33_30, key_c_r_33_31, key_c_r_33_32, key_c_r_33_33, key_c_r_33_34, 
       key_c_r_33_35, key_c_r_33_36, key_c_r_33_37, key_c_r_33_38, key_c_r_33_39, key_c_r_33_4, key_c_r_33_40, key_c_r_33_41, key_c_r_33_42, 
       key_c_r_33_43, key_c_r_33_44, key_c_r_33_45, key_c_r_33_46, key_c_r_33_47, key_c_r_33_48, key_c_r_33_49, key_c_r_33_5, key_c_r_33_50, 
       key_c_r_33_51, key_c_r_33_52, key_c_r_33_53, key_c_r_33_54, key_c_r_33_55, key_c_r_33_6, key_c_r_33_7, key_c_r_33_8, key_c_r_33_9, 
       key_c_r_3_0, key_c_r_3_1, key_c_r_3_10, key_c_r_3_11, key_c_r_3_12, key_c_r_3_13, key_c_r_3_14, key_c_r_3_15, key_c_r_3_16, 
       key_c_r_3_17, key_c_r_3_18, key_c_r_3_19, key_c_r_3_2, key_c_r_3_20, key_c_r_3_21, key_c_r_3_22, key_c_r_3_23, key_c_r_3_24, 
       key_c_r_3_25, key_c_r_3_26, key_c_r_3_27, key_c_r_3_28, key_c_r_3_29, key_c_r_3_3, key_c_r_3_30, key_c_r_3_31, key_c_r_3_32, 
       key_c_r_3_33, key_c_r_3_34, key_c_r_3_35, key_c_r_3_36, key_c_r_3_37, key_c_r_3_38, key_c_r_3_39, key_c_r_3_4, key_c_r_3_40, 
       key_c_r_3_41, key_c_r_3_42, key_c_r_3_43, key_c_r_3_44, key_c_r_3_45, key_c_r_3_46, key_c_r_3_47, key_c_r_3_48, key_c_r_3_49, 
       key_c_r_3_5, key_c_r_3_50, key_c_r_3_51, key_c_r_3_52, key_c_r_3_53, key_c_r_3_54, key_c_r_3_55, key_c_r_3_6, key_c_r_3_7, 
       key_c_r_3_8, key_c_r_3_9, key_c_r_4_0, key_c_r_4_1, key_c_r_4_10, key_c_r_4_11, key_c_r_4_12, key_c_r_4_13, key_c_r_4_14, 
       key_c_r_4_15, key_c_r_4_16, key_c_r_4_17, key_c_r_4_18, key_c_r_4_19, key_c_r_4_2, key_c_r_4_20, key_c_r_4_21, key_c_r_4_22, 
       key_c_r_4_23, key_c_r_4_24, key_c_r_4_25, key_c_r_4_26, key_c_r_4_27, key_c_r_4_28, key_c_r_4_29, key_c_r_4_3, key_c_r_4_30, 
       key_c_r_4_31, key_c_r_4_32, key_c_r_4_33, key_c_r_4_34, key_c_r_4_35, key_c_r_4_36, key_c_r_4_37, key_c_r_4_38, key_c_r_4_39, 
       key_c_r_4_4, key_c_r_4_40, key_c_r_4_41, key_c_r_4_42, key_c_r_4_43, key_c_r_4_44, key_c_r_4_45, key_c_r_4_46, key_c_r_4_47, 
       key_c_r_4_48, key_c_r_4_49, key_c_r_4_5, key_c_r_4_50, key_c_r_4_51, key_c_r_4_52, key_c_r_4_53, key_c_r_4_54, key_c_r_4_55, 
       key_c_r_4_6, key_c_r_4_7, key_c_r_4_8, key_c_r_4_9, key_c_r_5_0, key_c_r_5_1, key_c_r_5_10, key_c_r_5_11, key_c_r_5_12, 
       key_c_r_5_13, key_c_r_5_14, key_c_r_5_15, key_c_r_5_16, key_c_r_5_17, key_c_r_5_18, key_c_r_5_19, key_c_r_5_2, key_c_r_5_20, 
       key_c_r_5_21, key_c_r_5_22, key_c_r_5_23, key_c_r_5_24, key_c_r_5_25, key_c_r_5_26, key_c_r_5_27, key_c_r_5_28, key_c_r_5_29, 
       key_c_r_5_3, key_c_r_5_30, key_c_r_5_31, key_c_r_5_32, key_c_r_5_33, key_c_r_5_34, key_c_r_5_35, key_c_r_5_36, key_c_r_5_37, 
       key_c_r_5_38, key_c_r_5_39, key_c_r_5_4, key_c_r_5_40, key_c_r_5_41, key_c_r_5_42, key_c_r_5_43, key_c_r_5_44, key_c_r_5_45, 
       key_c_r_5_46, key_c_r_5_47, key_c_r_5_48, key_c_r_5_49, key_c_r_5_5, key_c_r_5_50, key_c_r_5_51, key_c_r_5_52, key_c_r_5_53, 
       key_c_r_5_54, key_c_r_5_55, key_c_r_5_6, key_c_r_5_7, key_c_r_5_8, key_c_r_5_9, key_c_r_6_0, key_c_r_6_1, key_c_r_6_10, 
       key_c_r_6_11, key_c_r_6_12, key_c_r_6_13, key_c_r_6_14, key_c_r_6_15, key_c_r_6_16, key_c_r_6_17, key_c_r_6_18, key_c_r_6_19, 
       key_c_r_6_2, key_c_r_6_20, key_c_r_6_21, key_c_r_6_22, key_c_r_6_23, key_c_r_6_24, key_c_r_6_25, key_c_r_6_26, key_c_r_6_27, 
       key_c_r_6_28, key_c_r_6_29, key_c_r_6_3, key_c_r_6_30, key_c_r_6_31, key_c_r_6_32, key_c_r_6_33, key_c_r_6_34, key_c_r_6_35, 
       key_c_r_6_36, key_c_r_6_37, key_c_r_6_38, key_c_r_6_39, key_c_r_6_4, key_c_r_6_40, key_c_r_6_41, key_c_r_6_42, key_c_r_6_43, 
       key_c_r_6_44, key_c_r_6_45, key_c_r_6_46, key_c_r_6_47, key_c_r_6_48, key_c_r_6_49, key_c_r_6_5, key_c_r_6_50, key_c_r_6_51, 
       key_c_r_6_52, key_c_r_6_53, key_c_r_6_54, key_c_r_6_55, key_c_r_6_6, key_c_r_6_7, key_c_r_6_8, key_c_r_6_9, key_c_r_7_0, 
       key_c_r_7_1, key_c_r_7_10, key_c_r_7_11, key_c_r_7_12, key_c_r_7_13, key_c_r_7_14, key_c_r_7_15, key_c_r_7_16, key_c_r_7_17, 
       key_c_r_7_18, key_c_r_7_19, key_c_r_7_2, key_c_r_7_20, key_c_r_7_21, key_c_r_7_22, key_c_r_7_23, key_c_r_7_24, key_c_r_7_25, 
       key_c_r_7_26, key_c_r_7_27, key_c_r_7_28, key_c_r_7_29, key_c_r_7_3, key_c_r_7_30, key_c_r_7_31, key_c_r_7_32, key_c_r_7_33, 
       key_c_r_7_34, key_c_r_7_35, key_c_r_7_36, key_c_r_7_37, key_c_r_7_38, key_c_r_7_39, key_c_r_7_4, key_c_r_7_40, key_c_r_7_41, 
       key_c_r_7_42, key_c_r_7_43, key_c_r_7_44, key_c_r_7_45, key_c_r_7_46, key_c_r_7_47, key_c_r_7_48, key_c_r_7_49, key_c_r_7_5, 
       key_c_r_7_50, key_c_r_7_51, key_c_r_7_52, key_c_r_7_53, key_c_r_7_54, key_c_r_7_55, key_c_r_7_6, key_c_r_7_7, key_c_r_7_8, 
       key_c_r_7_9, key_c_r_8_0, key_c_r_8_1, key_c_r_8_10, key_c_r_8_11, key_c_r_8_12, key_c_r_8_13, key_c_r_8_14, key_c_r_8_15, 
       key_c_r_8_16, key_c_r_8_17, key_c_r_8_18, key_c_r_8_19, key_c_r_8_2, key_c_r_8_20, key_c_r_8_21, key_c_r_8_22, key_c_r_8_23, 
       key_c_r_8_24, key_c_r_8_25, key_c_r_8_26, key_c_r_8_27, key_c_r_8_28, key_c_r_8_29, key_c_r_8_3, key_c_r_8_30, key_c_r_8_31, 
       key_c_r_8_32, key_c_r_8_33, key_c_r_8_34, key_c_r_8_35, key_c_r_8_36, key_c_r_8_37, key_c_r_8_38, key_c_r_8_39, key_c_r_8_4, 
       key_c_r_8_40, key_c_r_8_41, key_c_r_8_42, key_c_r_8_43, key_c_r_8_44, key_c_r_8_45, key_c_r_8_46, key_c_r_8_47, key_c_r_8_48, 
       key_c_r_8_49, key_c_r_8_5, key_c_r_8_50, key_c_r_8_51, key_c_r_8_52, key_c_r_8_53, key_c_r_8_54, key_c_r_8_55, key_c_r_8_6, 
       key_c_r_8_7, key_c_r_8_8, key_c_r_8_9, key_c_r_9_0, key_c_r_9_1, key_c_r_9_10, key_c_r_9_11, key_c_r_9_12, key_c_r_9_13, 
       key_c_r_9_14, key_c_r_9_15, key_c_r_9_16, key_c_r_9_17, key_c_r_9_18, key_c_r_9_19, key_c_r_9_2, key_c_r_9_20, key_c_r_9_21, 
       key_c_r_9_22, key_c_r_9_23, key_c_r_9_24, key_c_r_9_25, key_c_r_9_26, key_c_r_9_27, key_c_r_9_28, key_c_r_9_29, key_c_r_9_3, 
       key_c_r_9_30, key_c_r_9_31, key_c_r_9_32, key_c_r_9_33, key_c_r_9_34, key_c_r_9_35, key_c_r_9_36, key_c_r_9_37, key_c_r_9_38, 
       key_c_r_9_39, key_c_r_9_4, key_c_r_9_40, key_c_r_9_41, key_c_r_9_42, key_c_r_9_43, key_c_r_9_44, key_c_r_9_45, key_c_r_9_46, 
       key_c_r_9_47, key_c_r_9_48, key_c_r_9_49, key_c_r_9_5, key_c_r_9_50, key_c_r_9_51, key_c_r_9_52, key_c_r_9_53, key_c_r_9_54, 
       key_c_r_9_55, key_c_r_9_6, key_c_r_9_7, key_c_r_9_8, key_c_r_9_9, n1, n10, n100, n101, 
       n102, n103, n104, n105, n106, n107, n108, n109, n11, 
       n110, n111, n112, n114, n115, n116, n12, n13, n14, 
       n15, n16, n17, n18, n19, n2, n20, n21, n22, 
       n23, n24, n25, n26, n27, n28, n29, n3, n30, 
       n31, n32, n33, n34, n35, n36, n37, n38, n39, 
       n4, n40, n41, n42, n43, n44, n45, n46, n47, 
       n48, n49, n5, n50, n51, n52, n53, n54, n55, 
       n56, n57, n58, n59, n6, n60, n61, n62, n63, 
       n64, n65, n66, n67, n68, n69, n7, n70, n71, 
       n72, n73, n74, n75, n76, n77, n78, n79, n8, 
       n80, n81, n82, n83, n84, n85, n86, n87, n88, 
       n89, n9, n90, n91, n92, n93, n94, n95, n96, 
       n97, n98, n99, stage1_out_0, stage1_out_1, stage1_out_10, stage1_out_11, stage1_out_12, stage1_out_13, 
       stage1_out_14, stage1_out_15, stage1_out_16, stage1_out_17, stage1_out_18, stage1_out_19, stage1_out_2, stage1_out_20, stage1_out_21, 
       stage1_out_22, stage1_out_23, stage1_out_24, stage1_out_25, stage1_out_26, stage1_out_27, stage1_out_28, stage1_out_29, stage1_out_3, 
       stage1_out_30, stage1_out_31, stage1_out_32, stage1_out_33, stage1_out_34, stage1_out_35, stage1_out_36, stage1_out_37, stage1_out_38, 
       stage1_out_39, stage1_out_4, stage1_out_40, stage1_out_41, stage1_out_42, stage1_out_43, stage1_out_44, stage1_out_45, stage1_out_46, 
       stage1_out_47, stage1_out_48, stage1_out_49, stage1_out_5, stage1_out_50, stage1_out_51, stage1_out_52, stage1_out_53, stage1_out_54, 
       stage1_out_55, stage1_out_56, stage1_out_57, stage1_out_58, stage1_out_59, stage1_out_6, stage1_out_60, stage1_out_61, stage1_out_62, 
       stage1_out_63, stage1_out_7, stage1_out_8, stage1_out_9, stage2_out_0, stage2_out_1, stage2_out_10, stage2_out_11, stage2_out_12, 
       stage2_out_13, stage2_out_14, stage2_out_15, stage2_out_16, stage2_out_17, stage2_out_18, stage2_out_19, stage2_out_2, stage2_out_20, 
       stage2_out_21, stage2_out_22, stage2_out_23, stage2_out_24, stage2_out_25, stage2_out_26, stage2_out_27, stage2_out_28, stage2_out_29, 
       stage2_out_3, stage2_out_30, stage2_out_31, stage2_out_32, stage2_out_33, stage2_out_34, stage2_out_35, stage2_out_36, stage2_out_37, 
       stage2_out_38, stage2_out_39, stage2_out_4, stage2_out_40, stage2_out_41, stage2_out_42, stage2_out_43, stage2_out_44, stage2_out_45, 
       stage2_out_46, stage2_out_47, stage2_out_48, stage2_out_49, stage2_out_5, stage2_out_50, stage2_out_51, stage2_out_52, stage2_out_53, 
       stage2_out_54, stage2_out_55, stage2_out_56, stage2_out_57, stage2_out_58, stage2_out_59, stage2_out_6, stage2_out_60, stage2_out_61, 
       stage2_out_62, stage2_out_63, stage2_out_7, stage2_out_8, stage2_out_9, u0_FP_1, u0_FP_10, u0_FP_11, u0_FP_12, 
       u0_FP_13, u0_FP_14, u0_FP_15, u0_FP_16, u0_FP_17, u0_FP_18, u0_FP_19, u0_FP_2, u0_FP_20, 
       u0_FP_21, u0_FP_22, u0_FP_23, u0_FP_24, u0_FP_25, u0_FP_26, u0_FP_27, u0_FP_28, u0_FP_29, 
       u0_FP_3, u0_FP_30, u0_FP_31, u0_FP_32, u0_FP_35, u0_FP_38, u0_FP_4, u0_FP_40, u0_FP_47, 
       u0_FP_5, u0_FP_54, u0_FP_6, u0_FP_61, u0_FP_62, u0_FP_7, u0_FP_8, u0_FP_9, u0_K10_10, 
       u0_K10_11, u0_K10_13, u0_K10_15, u0_K10_16, u0_K10_21, u0_K10_22, u0_K10_23, u0_K10_25, u0_K10_27, 
       u0_K10_3, u0_K10_34, u0_K10_35, u0_K10_36, u0_K10_37, u0_K10_38, u0_K10_39, u0_K10_4, u0_K10_41, 
       u0_K10_43, u0_K10_46, u0_K10_5, u0_K10_7, u0_K11_21, u0_K11_22, u0_K11_34, u0_K11_41, u0_K11_43, 
       u0_K12_1, u0_K12_10, u0_K12_11, u0_K12_12, u0_K12_13, u0_K12_14, u0_K12_15, u0_K12_16, u0_K12_18, 
       u0_K12_20, u0_K12_22, u0_K12_33, u0_K12_34, u0_K12_39, u0_K12_40, u0_K12_45, u0_K12_46, u0_K12_47, 
       u0_K12_9, u0_K13_10, u0_K13_11, u0_K13_12, u0_K13_13, u0_K13_14, u0_K13_2, u0_K13_24, u0_K13_26, 
       u0_K13_27, u0_K13_28, u0_K13_30, u0_K13_32, u0_K13_33, u0_K13_34, u0_K13_35, u0_K13_36, u0_K13_37, 
       u0_K13_38, u0_K13_39, u0_K13_40, u0_K13_42, u0_K13_44, u0_K13_45, u0_K13_46, u0_K13_48, u0_K13_5, 
       u0_K13_7, u0_K14_1, u0_K14_10, u0_K14_11, u0_K14_12, u0_K14_13, u0_K14_14, u0_K14_15, u0_K14_16, 
       u0_K14_17, u0_K14_18, u0_K14_19, u0_K14_2, u0_K14_20, u0_K14_21, u0_K14_22, u0_K14_27, u0_K14_3, 
       u0_K14_30, u0_K14_32, u0_K14_36, u0_K14_38, u0_K14_39, u0_K14_4, u0_K14_40, u0_K14_41, u0_K14_42, 
       u0_K14_43, u0_K14_44, u0_K14_46, u0_K14_47, u0_K14_48, u0_K14_6, u0_K14_8, u0_K14_9, u0_K15_1, 
       u0_K15_10, u0_K15_12, u0_K15_14, u0_K15_15, u0_K15_16, u0_K15_17, u0_K15_18, u0_K15_19, u0_K15_2, 
       u0_K15_20, u0_K15_21, u0_K15_22, u0_K15_23, u0_K15_24, u0_K15_25, u0_K15_3, u0_K15_4, u0_K15_47, 
       u0_K15_48, u0_K15_5, u0_K15_6, u0_K15_7, u0_K15_8, u0_K15_9, u0_K16_11, u0_K16_13, u0_K16_22, 
       u0_K16_33, u0_K16_4, u0_K16_42, u0_K16_44, u0_K16_45, u0_K16_9, u0_K1_15, u0_K1_16, u0_K1_21, 
       u0_K1_22, u0_K1_23, u0_K1_25, u0_K1_28, u0_K1_33, u0_K1_42, u0_K1_44, u0_K1_45, u0_K1_46, 
       u0_K2_15, u0_K2_16, u0_K2_17, u0_K2_19, u0_K2_21, u0_K2_23, u0_K2_24, u0_K2_25, u0_K2_26, 
       u0_K2_3, u0_K2_33, u0_K2_34, u0_K2_35, u0_K2_36, u0_K2_37, u0_K2_38, u0_K2_39, u0_K2_4, 
       u0_K2_40, u0_K2_42, u0_K2_43, u0_K2_44, u0_K2_45, u0_K2_46, u0_K2_47, u0_K2_48, u0_K2_6, 
       u0_K2_8, u0_K2_9, u0_K3_10, u0_K3_15, u0_K3_16, u0_K3_24, u0_K3_26, u0_K3_27, u0_K3_3, 
       u0_K3_34, u0_K3_46, u0_K3_9, u0_K4_22, u0_K4_24, u0_K4_26, u0_K4_27, u0_K4_28, u0_K4_29, 
       u0_K4_31, u0_K4_34, u0_K4_35, u0_K4_37, u0_K4_39, u0_K4_40, u0_K4_42, u0_K4_44, u0_K4_45, 
       u0_K4_46, u0_K5_10, u0_K5_11, u0_K5_12, u0_K5_13, u0_K5_14, u0_K5_15, u0_K5_16, u0_K5_17, 
       u0_K5_19, u0_K5_2, u0_K5_21, u0_K5_23, u0_K5_25, u0_K5_28, u0_K5_3, u0_K5_30, u0_K5_32, 
       u0_K5_34, u0_K5_37, u0_K5_38, u0_K5_39, u0_K5_4, u0_K5_40, u0_K5_41, u0_K5_42, u0_K5_43, 
       u0_K5_44, u0_K5_45, u0_K5_46, u0_K5_48, u0_K5_5, u0_K5_7, u0_K5_9, u0_K6_10, u0_K6_15, 
       u0_K6_16, u0_K6_21, u0_K6_22, u0_K6_27, u0_K6_3, u0_K6_34, u0_K6_46, u0_K6_9, u0_K7_15, 
       u0_K7_16, u0_K7_2, u0_K7_21, u0_K7_22, u0_K7_23, u0_K7_24, u0_K7_25, u0_K7_26, u0_K7_27, 
       u0_K7_28, u0_K7_29, u0_K7_30, u0_K7_31, u0_K7_32, u0_K7_33, u0_K7_34, u0_K7_35, u0_K7_37, 
       u0_K7_38, u0_K7_39, u0_K7_40, u0_K7_41, u0_K7_42, u0_K7_43, u0_K7_44, u0_K7_45, u0_K7_46, 
       u0_K7_47, u0_K7_48, u0_K7_9, u0_K8_1, u0_K8_2, u0_K8_22, u0_K8_23, u0_K8_25, u0_K8_27, 
       u0_K8_28, u0_K8_29, u0_K8_3, u0_K8_30, u0_K8_31, u0_K8_32, u0_K8_33, u0_K8_34, u0_K8_36, 
       u0_K8_38, u0_K8_4, u0_K8_40, u0_K8_45, u0_K8_46, u0_K8_47, u0_K8_48, u0_K8_9, u0_K9_10, 
       u0_K9_15, u0_K9_16, u0_K9_18, u0_K9_20, u0_K9_22, u0_K9_23, u0_K9_25, u0_K9_27, u0_K9_28, 
       u0_K9_3, u0_K9_39, u0_K9_4, u0_K9_40, u0_K9_45, u0_K9_46, u0_K9_9, u0_L0_1, u0_L0_10, 
       u0_L0_11, u0_L0_12, u0_L0_13, u0_L0_14, u0_L0_15, u0_L0_16, u0_L0_17, u0_L0_18, u0_L0_19, 
       u0_L0_2, u0_L0_20, u0_L0_21, u0_L0_22, u0_L0_23, u0_L0_24, u0_L0_25, u0_L0_26, u0_L0_27, 
       u0_L0_28, u0_L0_29, u0_L0_3, u0_L0_30, u0_L0_31, u0_L0_32, u0_L0_4, u0_L0_5, u0_L0_6, 
       u0_L0_7, u0_L0_8, u0_L0_9, u0_L10_1, u0_L10_10, u0_L10_11, u0_L10_12, u0_L10_13, u0_L10_14, 
       u0_L10_15, u0_L10_16, u0_L10_17, u0_L10_18, u0_L10_19, u0_L10_2, u0_L10_20, u0_L10_21, u0_L10_22, 
       u0_L10_23, u0_L10_24, u0_L10_25, u0_L10_26, u0_L10_27, u0_L10_28, u0_L10_29, u0_L10_3, u0_L10_30, 
       u0_L10_31, u0_L10_32, u0_L10_4, u0_L10_5, u0_L10_6, u0_L10_7, u0_L10_8, u0_L10_9, u0_L11_1, 
       u0_L11_10, u0_L11_11, u0_L11_12, u0_L11_13, u0_L11_14, u0_L11_15, u0_L11_16, u0_L11_17, u0_L11_18, 
       u0_L11_19, u0_L11_2, u0_L11_20, u0_L11_21, u0_L11_22, u0_L11_23, u0_L11_24, u0_L11_25, u0_L11_26, 
       u0_L11_27, u0_L11_28, u0_L11_29, u0_L11_3, u0_L11_30, u0_L11_31, u0_L11_32, u0_L11_4, u0_L11_5, 
       u0_L11_6, u0_L11_7, u0_L11_8, u0_L11_9, u0_L12_1, u0_L12_10, u0_L12_11, u0_L12_12, u0_L12_13, 
       u0_L12_14, u0_L12_15, u0_L12_16, u0_L12_17, u0_L12_18, u0_L12_19, u0_L12_2, u0_L12_20, u0_L12_21, 
       u0_L12_22, u0_L12_23, u0_L12_24, u0_L12_25, u0_L12_26, u0_L12_27, u0_L12_28, u0_L12_29, u0_L12_3, 
       u0_L12_30, u0_L12_31, u0_L12_32, u0_L12_4, u0_L12_5, u0_L12_6, u0_L12_7, u0_L12_8, u0_L12_9, 
       u0_L13_1, u0_L13_10, u0_L13_11, u0_L13_12, u0_L13_13, u0_L13_14, u0_L13_15, u0_L13_16, u0_L13_17, 
       u0_L13_18, u0_L13_19, u0_L13_2, u0_L13_20, u0_L13_21, u0_L13_22, u0_L13_23, u0_L13_24, u0_L13_25, 
       u0_L13_26, u0_L13_27, u0_L13_28, u0_L13_29, u0_L13_3, u0_L13_30, u0_L13_31, u0_L13_32, u0_L13_4, 
       u0_L13_5, u0_L13_6, u0_L13_7, u0_L13_8, u0_L13_9, u0_L14_1, u0_L14_10, u0_L14_11, u0_L14_12, 
       u0_L14_13, u0_L14_14, u0_L14_15, u0_L14_16, u0_L14_17, u0_L14_18, u0_L14_19, u0_L14_2, u0_L14_20, 
       u0_L14_21, u0_L14_22, u0_L14_23, u0_L14_24, u0_L14_25, u0_L14_26, u0_L14_27, u0_L14_28, u0_L14_29, 
       u0_L14_3, u0_L14_30, u0_L14_31, u0_L14_32, u0_L14_4, u0_L14_5, u0_L14_6, u0_L14_7, u0_L14_8, 
       u0_L14_9, u0_L1_1, u0_L1_10, u0_L1_11, u0_L1_12, u0_L1_13, u0_L1_14, u0_L1_15, u0_L1_16, 
       u0_L1_17, u0_L1_18, u0_L1_19, u0_L1_2, u0_L1_20, u0_L1_21, u0_L1_22, u0_L1_23, u0_L1_24, 
       u0_L1_25, u0_L1_26, u0_L1_27, u0_L1_28, u0_L1_29, u0_L1_3, u0_L1_30, u0_L1_31, u0_L1_32, 
       u0_L1_4, u0_L1_5, u0_L1_6, u0_L1_7, u0_L1_8, u0_L1_9, u0_L2_1, u0_L2_10, u0_L2_11, 
       u0_L2_12, u0_L2_13, u0_L2_14, u0_L2_15, u0_L2_16, u0_L2_17, u0_L2_18, u0_L2_19, u0_L2_2, 
       u0_L2_20, u0_L2_21, u0_L2_22, u0_L2_23, u0_L2_24, u0_L2_25, u0_L2_26, u0_L2_27, u0_L2_28, 
       u0_L2_29, u0_L2_3, u0_L2_30, u0_L2_31, u0_L2_32, u0_L2_4, u0_L2_5, u0_L2_6, u0_L2_7, 
       u0_L2_8, u0_L2_9, u0_L3_1, u0_L3_10, u0_L3_11, u0_L3_12, u0_L3_13, u0_L3_14, u0_L3_15, 
       u0_L3_16, u0_L3_17, u0_L3_18, u0_L3_19, u0_L3_2, u0_L3_20, u0_L3_21, u0_L3_22, u0_L3_23, 
       u0_L3_24, u0_L3_25, u0_L3_26, u0_L3_27, u0_L3_28, u0_L3_29, u0_L3_3, u0_L3_30, u0_L3_31, 
       u0_L3_32, u0_L3_4, u0_L3_5, u0_L3_6, u0_L3_7, u0_L3_8, u0_L3_9, u0_L4_1, u0_L4_10, 
       u0_L4_11, u0_L4_12, u0_L4_13, u0_L4_14, u0_L4_15, u0_L4_16, u0_L4_17, u0_L4_18, u0_L4_19, 
       u0_L4_2, u0_L4_20, u0_L4_21, u0_L4_22, u0_L4_23, u0_L4_24, u0_L4_25, u0_L4_26, u0_L4_27, 
       u0_L4_28, u0_L4_29, u0_L4_3, u0_L4_30, u0_L4_31, u0_L4_32, u0_L4_4, u0_L4_5, u0_L4_6, 
       u0_L4_7, u0_L4_8, u0_L4_9, u0_L5_1, u0_L5_10, u0_L5_11, u0_L5_12, u0_L5_13, u0_L5_14, 
       u0_L5_15, u0_L5_16, u0_L5_17, u0_L5_18, u0_L5_19, u0_L5_2, u0_L5_20, u0_L5_21, u0_L5_22, 
       u0_L5_23, u0_L5_24, u0_L5_25, u0_L5_26, u0_L5_27, u0_L5_28, u0_L5_29, u0_L5_3, u0_L5_30, 
       u0_L5_31, u0_L5_32, u0_L5_4, u0_L5_5, u0_L5_6, u0_L5_7, u0_L5_8, u0_L5_9, u0_L6_1, 
       u0_L6_10, u0_L6_11, u0_L6_12, u0_L6_13, u0_L6_14, u0_L6_15, u0_L6_16, u0_L6_17, u0_L6_18, 
       u0_L6_19, u0_L6_2, u0_L6_20, u0_L6_21, u0_L6_22, u0_L6_23, u0_L6_24, u0_L6_25, u0_L6_26, 
       u0_L6_27, u0_L6_28, u0_L6_29, u0_L6_3, u0_L6_30, u0_L6_31, u0_L6_32, u0_L6_4, u0_L6_5, 
       u0_L6_6, u0_L6_7, u0_L6_8, u0_L6_9, u0_L7_1, u0_L7_10, u0_L7_11, u0_L7_12, u0_L7_13, 
       u0_L7_14, u0_L7_15, u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_19, u0_L7_2, u0_L7_20, u0_L7_21, 
       u0_L7_22, u0_L7_23, u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_28, u0_L7_29, u0_L7_3, 
       u0_L7_30, u0_L7_31, u0_L7_32, u0_L7_4, u0_L7_5, u0_L7_6, u0_L7_7, u0_L7_8, u0_L7_9, 
       u0_L8_1, u0_L8_10, u0_L8_11, u0_L8_12, u0_L8_13, u0_L8_14, u0_L8_15, u0_L8_16, u0_L8_17, 
       u0_L8_18, u0_L8_19, u0_L8_2, u0_L8_20, u0_L8_21, u0_L8_22, u0_L8_23, u0_L8_24, u0_L8_25, 
       u0_L8_26, u0_L8_27, u0_L8_28, u0_L8_29, u0_L8_3, u0_L8_30, u0_L8_31, u0_L8_32, u0_L8_4, 
       u0_L8_5, u0_L8_6, u0_L8_7, u0_L8_8, u0_L8_9, u0_L9_1, u0_L9_10, u0_L9_11, u0_L9_12, 
       u0_L9_13, u0_L9_14, u0_L9_15, u0_L9_16, u0_L9_17, u0_L9_18, u0_L9_19, u0_L9_2, u0_L9_20, 
       u0_L9_21, u0_L9_22, u0_L9_23, u0_L9_24, u0_L9_25, u0_L9_26, u0_L9_27, u0_L9_28, u0_L9_29, 
       u0_L9_3, u0_L9_30, u0_L9_31, u0_L9_32, u0_L9_4, u0_L9_5, u0_L9_6, u0_L9_7, u0_L9_8, 
       u0_L9_9, u0_N0, u0_N1, u0_N10, u0_N100, u0_N101, u0_N102, u0_N103, u0_N104, 
       u0_N105, u0_N106, u0_N107, u0_N108, u0_N109, u0_N11, u0_N110, u0_N111, u0_N112, 
       u0_N113, u0_N114, u0_N115, u0_N116, u0_N117, u0_N118, u0_N119, u0_N12, u0_N120, 
       u0_N121, u0_N122, u0_N123, u0_N124, u0_N125, u0_N126, u0_N127, u0_N128, u0_N129, 
       u0_N13, u0_N130, u0_N131, u0_N132, u0_N133, u0_N134, u0_N135, u0_N136, u0_N137, 
       u0_N138, u0_N139, u0_N14, u0_N140, u0_N141, u0_N142, u0_N143, u0_N144, u0_N145, 
       u0_N146, u0_N147, u0_N148, u0_N149, u0_N15, u0_N150, u0_N151, u0_N152, u0_N153, 
       u0_N154, u0_N155, u0_N156, u0_N157, u0_N158, u0_N159, u0_N16, u0_N160, u0_N161, 
       u0_N162, u0_N163, u0_N164, u0_N165, u0_N166, u0_N167, u0_N168, u0_N169, u0_N17, 
       u0_N170, u0_N171, u0_N172, u0_N173, u0_N174, u0_N175, u0_N176, u0_N177, u0_N178, 
       u0_N179, u0_N18, u0_N180, u0_N181, u0_N182, u0_N183, u0_N184, u0_N185, u0_N186, 
       u0_N187, u0_N188, u0_N189, u0_N19, u0_N190, u0_N191, u0_N192, u0_N193, u0_N194, 
       u0_N195, u0_N196, u0_N197, u0_N198, u0_N199, u0_N2, u0_N20, u0_N200, u0_N201, 
       u0_N202, u0_N203, u0_N204, u0_N205, u0_N206, u0_N207, u0_N208, u0_N209, u0_N21, 
       u0_N210, u0_N211, u0_N212, u0_N213, u0_N214, u0_N215, u0_N216, u0_N217, u0_N218, 
       u0_N219, u0_N22, u0_N220, u0_N221, u0_N222, u0_N223, u0_N224, u0_N225, u0_N226, 
       u0_N227, u0_N228, u0_N229, u0_N23, u0_N230, u0_N231, u0_N232, u0_N233, u0_N234, 
       u0_N235, u0_N236, u0_N237, u0_N238, u0_N239, u0_N24, u0_N240, u0_N241, u0_N242, 
       u0_N243, u0_N244, u0_N245, u0_N246, u0_N247, u0_N248, u0_N249, u0_N25, u0_N250, 
       u0_N251, u0_N252, u0_N253, u0_N254, u0_N255, u0_N256, u0_N257, u0_N258, u0_N259, 
       u0_N26, u0_N260, u0_N261, u0_N262, u0_N263, u0_N264, u0_N265, u0_N266, u0_N267, 
       u0_N268, u0_N269, u0_N27, u0_N270, u0_N271, u0_N272, u0_N273, u0_N274, u0_N275, 
       u0_N276, u0_N277, u0_N278, u0_N279, u0_N28, u0_N280, u0_N281, u0_N282, u0_N283, 
       u0_N284, u0_N285, u0_N286, u0_N287, u0_N288, u0_N289, u0_N29, u0_N290, u0_N291, 
       u0_N292, u0_N293, u0_N294, u0_N295, u0_N296, u0_N297, u0_N298, u0_N299, u0_N3, 
       u0_N30, u0_N300, u0_N301, u0_N302, u0_N303, u0_N304, u0_N305, u0_N306, u0_N307, 
       u0_N308, u0_N309, u0_N31, u0_N310, u0_N311, u0_N312, u0_N313, u0_N314, u0_N315, 
       u0_N316, u0_N317, u0_N318, u0_N319, u0_N32, u0_N320, u0_N321, u0_N322, u0_N323, 
       u0_N324, u0_N325, u0_N326, u0_N327, u0_N328, u0_N329, u0_N33, u0_N330, u0_N331, 
       u0_N332, u0_N333, u0_N334, u0_N335, u0_N336, u0_N337, u0_N338, u0_N339, u0_N34, 
       u0_N340, u0_N341, u0_N342, u0_N343, u0_N344, u0_N345, u0_N346, u0_N347, u0_N348, 
       u0_N349, u0_N35, u0_N350, u0_N351, u0_N352, u0_N353, u0_N354, u0_N355, u0_N356, 
       u0_N357, u0_N358, u0_N359, u0_N36, u0_N360, u0_N361, u0_N362, u0_N363, u0_N364, 
       u0_N365, u0_N366, u0_N367, u0_N368, u0_N369, u0_N37, u0_N370, u0_N371, u0_N372, 
       u0_N373, u0_N374, u0_N375, u0_N376, u0_N377, u0_N378, u0_N379, u0_N38, u0_N380, 
       u0_N381, u0_N382, u0_N383, u0_N384, u0_N385, u0_N386, u0_N387, u0_N388, u0_N389, 
       u0_N39, u0_N390, u0_N391, u0_N392, u0_N393, u0_N394, u0_N395, u0_N396, u0_N397, 
       u0_N398, u0_N399, u0_N4, u0_N40, u0_N400, u0_N401, u0_N402, u0_N403, u0_N404, 
       u0_N405, u0_N406, u0_N407, u0_N408, u0_N409, u0_N41, u0_N410, u0_N411, u0_N412, 
       u0_N413, u0_N414, u0_N415, u0_N416, u0_N417, u0_N418, u0_N419, u0_N42, u0_N420, 
       u0_N421, u0_N422, u0_N423, u0_N424, u0_N425, u0_N426, u0_N427, u0_N428, u0_N429, 
       u0_N43, u0_N430, u0_N431, u0_N432, u0_N433, u0_N434, u0_N435, u0_N436, u0_N437, 
       u0_N438, u0_N439, u0_N44, u0_N440, u0_N441, u0_N442, u0_N443, u0_N444, u0_N445, 
       u0_N446, u0_N447, u0_N448, u0_N449, u0_N45, u0_N450, u0_N451, u0_N452, u0_N453, 
       u0_N454, u0_N455, u0_N456, u0_N457, u0_N458, u0_N459, u0_N46, u0_N460, u0_N461, 
       u0_N462, u0_N463, u0_N464, u0_N465, u0_N466, u0_N467, u0_N468, u0_N469, u0_N47, 
       u0_N470, u0_N471, u0_N472, u0_N473, u0_N474, u0_N475, u0_N476, u0_N477, u0_N478, 
       u0_N479, u0_N48, u0_N49, u0_N5, u0_N50, u0_N51, u0_N52, u0_N53, u0_N54, 
       u0_N55, u0_N56, u0_N57, u0_N58, u0_N59, u0_N6, u0_N60, u0_N61, u0_N62, 
       u0_N63, u0_N64, u0_N65, u0_N66, u0_N67, u0_N68, u0_N69, u0_N7, u0_N70, 
       u0_N71, u0_N72, u0_N73, u0_N74, u0_N75, u0_N76, u0_N77, u0_N78, u0_N79, 
       u0_N8, u0_N80, u0_N81, u0_N82, u0_N83, u0_N84, u0_N85, u0_N86, u0_N87, 
       u0_N88, u0_N89, u0_N9, u0_N90, u0_N91, u0_N92, u0_N93, u0_N94, u0_N95, 
       u0_N96, u0_N97, u0_N98, u0_N99, u0_R0_10, u0_R0_11, u0_R0_12, u0_R0_14, u0_R0_16, 
       u0_R0_17, u0_R0_2, u0_R0_22, u0_R0_23, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, u0_R0_29, 
       u0_R0_3, u0_R0_30, u0_R0_31, u0_R0_5, u0_R0_6, u0_R10_10, u0_R10_11, u0_R10_13, u0_R10_15, 
       u0_R10_22, u0_R10_23, u0_R10_26, u0_R10_27, u0_R10_30, u0_R10_31, u0_R10_32, u0_R10_6, u0_R10_7, 
       u0_R10_8, u0_R10_9, u0_R11_1, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_21, u0_R11_22, u0_R11_23, 
       u0_R11_24, u0_R11_25, u0_R11_26, u0_R11_27, u0_R11_29, u0_R11_30, u0_R11_31, u0_R11_4, u0_R11_7, 
       u0_R11_8, u0_R11_9, u0_R12_1, u0_R12_10, u0_R12_11, u0_R12_12, u0_R12_13, u0_R12_14, u0_R12_15, 
       u0_R12_18, u0_R12_2, u0_R12_21, u0_R12_25, u0_R12_26, u0_R12_27, u0_R12_28, u0_R12_29, u0_R12_3, 
       u0_R12_31, u0_R12_32, u0_R12_5, u0_R12_6, u0_R12_7, u0_R12_8, u0_R12_9, u0_R13_1, u0_R13_10, 
       u0_R13_11, u0_R13_12, u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_2, u0_R13_3, u0_R13_32, 
       u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_9, u0_R1_10, u0_R1_11, u0_R1_17, u0_R1_18, 
       u0_R1_2, u0_R1_23, u0_R1_31, u0_R1_6, u0_R1_7, u0_R2_15, u0_R2_17, u0_R2_18, u0_R2_19, 
       u0_R2_20, u0_R2_23, u0_R2_24, u0_R2_26, u0_R2_27, u0_R2_29, u0_R2_30, u0_R2_31, u0_R3_1, 
       u0_R3_10, u0_R3_11, u0_R3_12, u0_R3_14, u0_R3_16, u0_R3_19, u0_R3_2, u0_R3_21, u0_R3_23, 
       u0_R3_26, u0_R3_27, u0_R3_28, u0_R3_29, u0_R3_3, u0_R3_30, u0_R3_31, u0_R3_4, u0_R3_6, 
       u0_R3_7, u0_R3_8, u0_R3_9, u0_R4_10, u0_R4_11, u0_R4_14, u0_R4_15, u0_R4_18, u0_R4_2, 
       u0_R4_23, u0_R4_31, u0_R4_6, u0_R4_7, u0_R5_1, u0_R5_10, u0_R5_11, u0_R5_14, u0_R5_15, 
       u0_R5_16, u0_R5_17, u0_R5_18, u0_R5_19, u0_R5_20, u0_R5_21, u0_R5_22, u0_R5_23, u0_R5_24, 
       u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R5_30, u0_R5_31, u0_R5_6, u0_R6_1, u0_R6_15, 
       u0_R6_16, u0_R6_18, u0_R6_19, u0_R6_2, u0_R6_20, u0_R6_21, u0_R6_22, u0_R6_23, u0_R6_25, 
       u0_R6_27, u0_R6_3, u0_R6_30, u0_R6_31, u0_R6_32, u0_R6_6, u0_R7_10, u0_R7_11, u0_R7_13, 
       u0_R7_15, u0_R7_16, u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_26, u0_R7_27, u0_R7_3, u0_R7_30, 
       u0_R7_31, u0_R7_6, u0_R7_7, u0_R8_10, u0_R8_11, u0_R8_14, u0_R8_15, u0_R8_16, u0_R8_18, 
       u0_R8_2, u0_R8_23, u0_R8_24, u0_R8_25, u0_R8_26, u0_R8_28, u0_R8_3, u0_R8_31, u0_R8_4, 
       u0_R8_7, u0_R8_8, u0_R9_14, u0_R9_15, u0_R9_23, u0_R9_28, u0_desIn_r_0, u0_desIn_r_10, u0_desIn_r_12, 
       u0_desIn_r_13, u0_desIn_r_14, u0_desIn_r_16, u0_desIn_r_18, u0_desIn_r_19, u0_desIn_r_2, u0_desIn_r_20, u0_desIn_r_21, u0_desIn_r_22, 
       u0_desIn_r_24, u0_desIn_r_26, u0_desIn_r_28, u0_desIn_r_30, u0_desIn_r_32, u0_desIn_r_33, u0_desIn_r_34, u0_desIn_r_36, u0_desIn_r_38, 
       u0_desIn_r_4, u0_desIn_r_40, u0_desIn_r_41, u0_desIn_r_42, u0_desIn_r_43, u0_desIn_r_44, u0_desIn_r_45, u0_desIn_r_46, u0_desIn_r_48, 
       u0_desIn_r_49, u0_desIn_r_50, u0_desIn_r_52, u0_desIn_r_53, u0_desIn_r_54, u0_desIn_r_56, u0_desIn_r_58, u0_desIn_r_6, u0_desIn_r_60, 
       u0_desIn_r_61, u0_desIn_r_62, u0_desIn_r_8, u0_key_r_1, u0_key_r_10, u0_key_r_15, u0_key_r_17, u0_key_r_18, u0_key_r_24, 
       u0_key_r_25, u0_key_r_26, u0_key_r_27, u0_key_r_3, u0_key_r_31, u0_key_r_32, u0_key_r_33, u0_key_r_34, u0_key_r_36, 
       u0_key_r_37, u0_key_r_38, u0_key_r_39, u0_key_r_40, u0_key_r_43, u0_key_r_44, u0_key_r_45, u0_key_r_46, u0_key_r_49, 
       u0_key_r_51, u0_key_r_52, u0_key_r_53, u0_key_r_7, u0_key_r_8, u0_out13_16, u0_out13_24, u0_out13_30, u0_out13_6, 
       u0_out14_17, u0_out14_23, u0_out14_31, u0_out14_9, u0_out1_15, u0_out1_21, u0_out1_27, u0_out1_5, u0_out4_12, 
       u0_out4_22, u0_out4_32, u0_out4_7, u0_out6_12, u0_out6_14, u0_out6_15, u0_out6_21, u0_out6_22, u0_out6_25, 
       u0_out6_27, u0_out6_3, u0_out6_32, u0_out6_5, u0_out6_7, u0_out6_8, u0_u13_X_13, u0_u13_X_14, u0_u13_X_15, 
       u0_u13_X_16, u0_u13_X_17, u0_u13_X_18, u0_u13_u2_n100, u0_u13_u2_n101, u0_u13_u2_n102, u0_u13_u2_n103, u0_u13_u2_n104, u0_u13_u2_n105, 
       u0_u13_u2_n106, u0_u13_u2_n107, u0_u13_u2_n108, u0_u13_u2_n109, u0_u13_u2_n110, u0_u13_u2_n111, u0_u13_u2_n112, u0_u13_u2_n113, u0_u13_u2_n114, 
       u0_u13_u2_n115, u0_u13_u2_n116, u0_u13_u2_n117, u0_u13_u2_n118, u0_u13_u2_n119, u0_u13_u2_n120, u0_u13_u2_n121, u0_u13_u2_n122, u0_u13_u2_n123, 
       u0_u13_u2_n124, u0_u13_u2_n125, u0_u13_u2_n126, u0_u13_u2_n127, u0_u13_u2_n128, u0_u13_u2_n129, u0_u13_u2_n130, u0_u13_u2_n131, u0_u13_u2_n132, 
       u0_u13_u2_n133, u0_u13_u2_n134, u0_u13_u2_n135, u0_u13_u2_n136, u0_u13_u2_n137, u0_u13_u2_n138, u0_u13_u2_n139, u0_u13_u2_n140, u0_u13_u2_n141, 
       u0_u13_u2_n142, u0_u13_u2_n143, u0_u13_u2_n144, u0_u13_u2_n145, u0_u13_u2_n146, u0_u13_u2_n147, u0_u13_u2_n148, u0_u13_u2_n149, u0_u13_u2_n150, 
       u0_u13_u2_n151, u0_u13_u2_n152, u0_u13_u2_n153, u0_u13_u2_n154, u0_u13_u2_n155, u0_u13_u2_n156, u0_u13_u2_n157, u0_u13_u2_n158, u0_u13_u2_n159, 
       u0_u13_u2_n160, u0_u13_u2_n161, u0_u13_u2_n162, u0_u13_u2_n163, u0_u13_u2_n164, u0_u13_u2_n165, u0_u13_u2_n166, u0_u13_u2_n167, u0_u13_u2_n168, 
       u0_u13_u2_n169, u0_u13_u2_n170, u0_u13_u2_n171, u0_u13_u2_n172, u0_u13_u2_n173, u0_u13_u2_n174, u0_u13_u2_n175, u0_u13_u2_n176, u0_u13_u2_n177, 
       u0_u13_u2_n178, u0_u13_u2_n179, u0_u13_u2_n180, u0_u13_u2_n181, u0_u13_u2_n182, u0_u13_u2_n183, u0_u13_u2_n184, u0_u13_u2_n185, u0_u13_u2_n186, 
       u0_u13_u2_n187, u0_u13_u2_n188, u0_u13_u2_n95, u0_u13_u2_n96, u0_u13_u2_n97, u0_u13_u2_n98, u0_u13_u2_n99, u0_u14_X_1, u0_u14_X_2, 
       u0_u14_X_3, u0_u14_X_4, u0_u14_X_5, u0_u14_X_6, u0_u14_u0_n100, u0_u14_u0_n101, u0_u14_u0_n102, u0_u14_u0_n103, u0_u14_u0_n104, 
       u0_u14_u0_n105, u0_u14_u0_n106, u0_u14_u0_n107, u0_u14_u0_n108, u0_u14_u0_n109, u0_u14_u0_n110, u0_u14_u0_n111, u0_u14_u0_n112, u0_u14_u0_n113, 
       u0_u14_u0_n114, u0_u14_u0_n115, u0_u14_u0_n116, u0_u14_u0_n117, u0_u14_u0_n118, u0_u14_u0_n119, u0_u14_u0_n120, u0_u14_u0_n121, u0_u14_u0_n122, 
       u0_u14_u0_n123, u0_u14_u0_n124, u0_u14_u0_n125, u0_u14_u0_n126, u0_u14_u0_n127, u0_u14_u0_n128, u0_u14_u0_n129, u0_u14_u0_n130, u0_u14_u0_n131, 
       u0_u14_u0_n132, u0_u14_u0_n133, u0_u14_u0_n134, u0_u14_u0_n135, u0_u14_u0_n136, u0_u14_u0_n137, u0_u14_u0_n138, u0_u14_u0_n139, u0_u14_u0_n140, 
       u0_u14_u0_n141, u0_u14_u0_n142, u0_u14_u0_n143, u0_u14_u0_n144, u0_u14_u0_n145, u0_u14_u0_n146, u0_u14_u0_n147, u0_u14_u0_n148, u0_u14_u0_n149, 
       u0_u14_u0_n150, u0_u14_u0_n151, u0_u14_u0_n152, u0_u14_u0_n153, u0_u14_u0_n154, u0_u14_u0_n155, u0_u14_u0_n156, u0_u14_u0_n157, u0_u14_u0_n158, 
       u0_u14_u0_n159, u0_u14_u0_n160, u0_u14_u0_n161, u0_u14_u0_n162, u0_u14_u0_n163, u0_u14_u0_n164, u0_u14_u0_n165, u0_u14_u0_n166, u0_u14_u0_n167, 
       u0_u14_u0_n168, u0_u14_u0_n169, u0_u14_u0_n170, u0_u14_u0_n171, u0_u14_u0_n172, u0_u14_u0_n173, u0_u14_u0_n174, u0_u14_u0_n88, u0_u14_u0_n89, 
       u0_u14_u0_n90, u0_u14_u0_n91, u0_u14_u0_n92, u0_u14_u0_n93, u0_u14_u0_n94, u0_u14_u0_n95, u0_u14_u0_n96, u0_u14_u0_n97, u0_u14_u0_n98, 
       u0_u14_u0_n99, u0_u1_X_43, u0_u1_X_44, u0_u1_X_45, u0_u1_X_46, u0_u1_X_47, u0_u1_X_48, u0_u1_u7_n100, u0_u1_u7_n101, 
       u0_u1_u7_n102, u0_u1_u7_n103, u0_u1_u7_n104, u0_u1_u7_n105, u0_u1_u7_n106, u0_u1_u7_n107, u0_u1_u7_n108, u0_u1_u7_n109, u0_u1_u7_n110, 
       u0_u1_u7_n111, u0_u1_u7_n112, u0_u1_u7_n113, u0_u1_u7_n114, u0_u1_u7_n115, u0_u1_u7_n116, u0_u1_u7_n117, u0_u1_u7_n118, u0_u1_u7_n119, 
       u0_u1_u7_n120, u0_u1_u7_n121, u0_u1_u7_n122, u0_u1_u7_n123, u0_u1_u7_n124, u0_u1_u7_n125, u0_u1_u7_n126, u0_u1_u7_n127, u0_u1_u7_n128, 
       u0_u1_u7_n129, u0_u1_u7_n130, u0_u1_u7_n131, u0_u1_u7_n132, u0_u1_u7_n133, u0_u1_u7_n134, u0_u1_u7_n135, u0_u1_u7_n136, u0_u1_u7_n137, 
       u0_u1_u7_n138, u0_u1_u7_n139, u0_u1_u7_n140, u0_u1_u7_n141, u0_u1_u7_n142, u0_u1_u7_n143, u0_u1_u7_n144, u0_u1_u7_n145, u0_u1_u7_n146, 
       u0_u1_u7_n147, u0_u1_u7_n148, u0_u1_u7_n149, u0_u1_u7_n150, u0_u1_u7_n151, u0_u1_u7_n152, u0_u1_u7_n153, u0_u1_u7_n154, u0_u1_u7_n155, 
       u0_u1_u7_n156, u0_u1_u7_n157, u0_u1_u7_n158, u0_u1_u7_n159, u0_u1_u7_n160, u0_u1_u7_n161, u0_u1_u7_n162, u0_u1_u7_n163, u0_u1_u7_n164, 
       u0_u1_u7_n165, u0_u1_u7_n166, u0_u1_u7_n167, u0_u1_u7_n168, u0_u1_u7_n169, u0_u1_u7_n170, u0_u1_u7_n171, u0_u1_u7_n172, u0_u1_u7_n173, 
       u0_u1_u7_n174, u0_u1_u7_n175, u0_u1_u7_n176, u0_u1_u7_n177, u0_u1_u7_n178, u0_u1_u7_n179, u0_u1_u7_n180, u0_u1_u7_n91, u0_u1_u7_n92, 
       u0_u1_u7_n93, u0_u1_u7_n94, u0_u1_u7_n95, u0_u1_u7_n96, u0_u1_u7_n97, u0_u1_u7_n98, u0_u1_u7_n99, u0_u4_X_37, u0_u4_X_38, 
       u0_u4_X_39, u0_u4_X_40, u0_u4_X_41, u0_u4_X_42, u0_u4_u6_n100, u0_u4_u6_n101, u0_u4_u6_n102, u0_u4_u6_n103, u0_u4_u6_n104, 
       u0_u4_u6_n105, u0_u4_u6_n106, u0_u4_u6_n107, u0_u4_u6_n108, u0_u4_u6_n109, u0_u4_u6_n110, u0_u4_u6_n111, u0_u4_u6_n112, u0_u4_u6_n113, 
       u0_u4_u6_n114, u0_u4_u6_n115, u0_u4_u6_n116, u0_u4_u6_n117, u0_u4_u6_n118, u0_u4_u6_n119, u0_u4_u6_n120, u0_u4_u6_n121, u0_u4_u6_n122, 
       u0_u4_u6_n123, u0_u4_u6_n124, u0_u4_u6_n125, u0_u4_u6_n126, u0_u4_u6_n127, u0_u4_u6_n128, u0_u4_u6_n129, u0_u4_u6_n130, u0_u4_u6_n131, 
       u0_u4_u6_n132, u0_u4_u6_n133, u0_u4_u6_n134, u0_u4_u6_n135, u0_u4_u6_n136, u0_u4_u6_n137, u0_u4_u6_n138, u0_u4_u6_n139, u0_u4_u6_n140, 
       u0_u4_u6_n141, u0_u4_u6_n142, u0_u4_u6_n143, u0_u4_u6_n144, u0_u4_u6_n145, u0_u4_u6_n146, u0_u4_u6_n147, u0_u4_u6_n148, u0_u4_u6_n149, 
       u0_u4_u6_n150, u0_u4_u6_n151, u0_u4_u6_n152, u0_u4_u6_n153, u0_u4_u6_n154, u0_u4_u6_n155, u0_u4_u6_n156, u0_u4_u6_n157, u0_u4_u6_n158, 
       u0_u4_u6_n159, u0_u4_u6_n160, u0_u4_u6_n161, u0_u4_u6_n162, u0_u4_u6_n163, u0_u4_u6_n164, u0_u4_u6_n165, u0_u4_u6_n166, u0_u4_u6_n167, 
       u0_u4_u6_n168, u0_u4_u6_n169, u0_u4_u6_n170, u0_u4_u6_n171, u0_u4_u6_n172, u0_u4_u6_n173, u0_u4_u6_n174, u0_u4_u6_n88, u0_u4_u6_n89, 
       u0_u4_u6_n90, u0_u4_u6_n91, u0_u4_u6_n92, u0_u4_u6_n93, u0_u4_u6_n94, u0_u4_u6_n95, u0_u4_u6_n96, u0_u4_u6_n97, u0_u4_u6_n98, 
       u0_u4_u6_n99, u0_u6_X_25, u0_u6_X_26, u0_u6_X_27, u0_u6_X_28, u0_u6_X_29, u0_u6_X_30, u0_u6_X_37, u0_u6_X_38, 
       u0_u6_X_39, u0_u6_X_40, u0_u6_X_41, u0_u6_X_42, u0_u6_X_43, u0_u6_X_44, u0_u6_X_45, u0_u6_X_46, u0_u6_X_47, 
       u0_u6_X_48, u0_u6_u4_n100, u0_u6_u4_n101, u0_u6_u4_n102, u0_u6_u4_n103, u0_u6_u4_n104, u0_u6_u4_n105, u0_u6_u4_n106, u0_u6_u4_n107, 
       u0_u6_u4_n108, u0_u6_u4_n109, u0_u6_u4_n110, u0_u6_u4_n111, u0_u6_u4_n112, u0_u6_u4_n113, u0_u6_u4_n114, u0_u6_u4_n115, u0_u6_u4_n116, 
       u0_u6_u4_n117, u0_u6_u4_n118, u0_u6_u4_n119, u0_u6_u4_n120, u0_u6_u4_n121, u0_u6_u4_n122, u0_u6_u4_n123, u0_u6_u4_n124, u0_u6_u4_n125, 
       u0_u6_u4_n126, u0_u6_u4_n127, u0_u6_u4_n128, u0_u6_u4_n129, u0_u6_u4_n130, u0_u6_u4_n131, u0_u6_u4_n132, u0_u6_u4_n133, u0_u6_u4_n134, 
       u0_u6_u4_n135, u0_u6_u4_n136, u0_u6_u4_n137, u0_u6_u4_n138, u0_u6_u4_n139, u0_u6_u4_n140, u0_u6_u4_n141, u0_u6_u4_n142, u0_u6_u4_n143, 
       u0_u6_u4_n144, u0_u6_u4_n145, u0_u6_u4_n146, u0_u6_u4_n147, u0_u6_u4_n148, u0_u6_u4_n149, u0_u6_u4_n150, u0_u6_u4_n151, u0_u6_u4_n152, 
       u0_u6_u4_n153, u0_u6_u4_n154, u0_u6_u4_n155, u0_u6_u4_n156, u0_u6_u4_n157, u0_u6_u4_n158, u0_u6_u4_n159, u0_u6_u4_n160, u0_u6_u4_n161, 
       u0_u6_u4_n162, u0_u6_u4_n163, u0_u6_u4_n164, u0_u6_u4_n165, u0_u6_u4_n166, u0_u6_u4_n167, u0_u6_u4_n168, u0_u6_u4_n169, u0_u6_u4_n170, 
       u0_u6_u4_n171, u0_u6_u4_n172, u0_u6_u4_n173, u0_u6_u4_n174, u0_u6_u4_n175, u0_u6_u4_n176, u0_u6_u4_n177, u0_u6_u4_n178, u0_u6_u4_n179, 
       u0_u6_u4_n180, u0_u6_u4_n181, u0_u6_u4_n182, u0_u6_u4_n183, u0_u6_u4_n184, u0_u6_u4_n185, u0_u6_u4_n186, u0_u6_u4_n94, u0_u6_u4_n95, 
       u0_u6_u4_n96, u0_u6_u4_n97, u0_u6_u4_n98, u0_u6_u4_n99, u0_u6_u6_n100, u0_u6_u6_n101, u0_u6_u6_n102, u0_u6_u6_n103, u0_u6_u6_n104, 
       u0_u6_u6_n105, u0_u6_u6_n106, u0_u6_u6_n107, u0_u6_u6_n108, u0_u6_u6_n109, u0_u6_u6_n110, u0_u6_u6_n111, u0_u6_u6_n112, u0_u6_u6_n113, 
       u0_u6_u6_n114, u0_u6_u6_n115, u0_u6_u6_n116, u0_u6_u6_n117, u0_u6_u6_n118, u0_u6_u6_n119, u0_u6_u6_n120, u0_u6_u6_n121, u0_u6_u6_n122, 
       u0_u6_u6_n123, u0_u6_u6_n124, u0_u6_u6_n125, u0_u6_u6_n126, u0_u6_u6_n127, u0_u6_u6_n128, u0_u6_u6_n129, u0_u6_u6_n130, u0_u6_u6_n131, 
       u0_u6_u6_n132, u0_u6_u6_n133, u0_u6_u6_n134, u0_u6_u6_n135, u0_u6_u6_n136, u0_u6_u6_n137, u0_u6_u6_n138, u0_u6_u6_n139, u0_u6_u6_n140, 
       u0_u6_u6_n141, u0_u6_u6_n142, u0_u6_u6_n143, u0_u6_u6_n144, u0_u6_u6_n145, u0_u6_u6_n146, u0_u6_u6_n147, u0_u6_u6_n148, u0_u6_u6_n149, 
       u0_u6_u6_n150, u0_u6_u6_n151, u0_u6_u6_n152, u0_u6_u6_n153, u0_u6_u6_n154, u0_u6_u6_n155, u0_u6_u6_n156, u0_u6_u6_n157, u0_u6_u6_n158, 
       u0_u6_u6_n159, u0_u6_u6_n160, u0_u6_u6_n161, u0_u6_u6_n162, u0_u6_u6_n163, u0_u6_u6_n164, u0_u6_u6_n165, u0_u6_u6_n166, u0_u6_u6_n167, 
       u0_u6_u6_n168, u0_u6_u6_n169, u0_u6_u6_n170, u0_u6_u6_n171, u0_u6_u6_n172, u0_u6_u6_n173, u0_u6_u6_n174, u0_u6_u6_n88, u0_u6_u6_n89, 
       u0_u6_u6_n90, u0_u6_u6_n91, u0_u6_u6_n92, u0_u6_u6_n93, u0_u6_u6_n94, u0_u6_u6_n95, u0_u6_u6_n96, u0_u6_u6_n97, u0_u6_u6_n98, 
       u0_u6_u6_n99, u0_u6_u7_n100, u0_u6_u7_n101, u0_u6_u7_n102, u0_u6_u7_n103, u0_u6_u7_n104, u0_u6_u7_n105, u0_u6_u7_n106, u0_u6_u7_n107, 
       u0_u6_u7_n108, u0_u6_u7_n109, u0_u6_u7_n110, u0_u6_u7_n111, u0_u6_u7_n112, u0_u6_u7_n113, u0_u6_u7_n114, u0_u6_u7_n115, u0_u6_u7_n116, 
       u0_u6_u7_n117, u0_u6_u7_n118, u0_u6_u7_n119, u0_u6_u7_n120, u0_u6_u7_n121, u0_u6_u7_n122, u0_u6_u7_n123, u0_u6_u7_n124, u0_u6_u7_n125, 
       u0_u6_u7_n126, u0_u6_u7_n127, u0_u6_u7_n128, u0_u6_u7_n129, u0_u6_u7_n130, u0_u6_u7_n131, u0_u6_u7_n132, u0_u6_u7_n133, u0_u6_u7_n134, 
       u0_u6_u7_n135, u0_u6_u7_n136, u0_u6_u7_n137, u0_u6_u7_n138, u0_u6_u7_n139, u0_u6_u7_n140, u0_u6_u7_n141, u0_u6_u7_n142, u0_u6_u7_n143, 
       u0_u6_u7_n144, u0_u6_u7_n145, u0_u6_u7_n146, u0_u6_u7_n147, u0_u6_u7_n148, u0_u6_u7_n149, u0_u6_u7_n150, u0_u6_u7_n151, u0_u6_u7_n152, 
       u0_u6_u7_n153, u0_u6_u7_n154, u0_u6_u7_n155, u0_u6_u7_n156, u0_u6_u7_n157, u0_u6_u7_n158, u0_u6_u7_n159, u0_u6_u7_n160, u0_u6_u7_n161, 
       u0_u6_u7_n162, u0_u6_u7_n163, u0_u6_u7_n164, u0_u6_u7_n165, u0_u6_u7_n166, u0_u6_u7_n167, u0_u6_u7_n168, u0_u6_u7_n169, u0_u6_u7_n170, 
       u0_u6_u7_n171, u0_u6_u7_n172, u0_u6_u7_n173, u0_u6_u7_n174, u0_u6_u7_n175, u0_u6_u7_n176, u0_u6_u7_n177, u0_u6_u7_n178, u0_u6_u7_n179, 
       u0_u6_u7_n180, u0_u6_u7_n91, u0_u6_u7_n92, u0_u6_u7_n93, u0_u6_u7_n94, u0_u6_u7_n95, u0_u6_u7_n96, u0_u6_u7_n97, u0_u6_u7_n98, 
       u0_u6_u7_n99, u0_uk_K_r0_0, u0_uk_K_r0_1, u0_uk_K_r0_10, u0_uk_K_r0_11, u0_uk_K_r0_12, u0_uk_K_r0_13, u0_uk_K_r0_14, u0_uk_K_r0_16, 
       u0_uk_K_r0_17, u0_uk_K_r0_18, u0_uk_K_r0_19, u0_uk_K_r0_2, u0_uk_K_r0_20, u0_uk_K_r0_21, u0_uk_K_r0_22, u0_uk_K_r0_23, u0_uk_K_r0_24, 
       u0_uk_K_r0_25, u0_uk_K_r0_26, u0_uk_K_r0_27, u0_uk_K_r0_29, u0_uk_K_r0_3, u0_uk_K_r0_30, u0_uk_K_r0_31, u0_uk_K_r0_32, u0_uk_K_r0_33, 
       u0_uk_K_r0_34, u0_uk_K_r0_35, u0_uk_K_r0_37, u0_uk_K_r0_38, u0_uk_K_r0_39, u0_uk_K_r0_4, u0_uk_K_r0_40, u0_uk_K_r0_41, u0_uk_K_r0_42, 
       u0_uk_K_r0_43, u0_uk_K_r0_44, u0_uk_K_r0_45, u0_uk_K_r0_46, u0_uk_K_r0_47, u0_uk_K_r0_48, u0_uk_K_r0_5, u0_uk_K_r0_50, u0_uk_K_r0_51, 
       u0_uk_K_r0_52, u0_uk_K_r0_53, u0_uk_K_r0_54, u0_uk_K_r0_55, u0_uk_K_r0_6, u0_uk_K_r0_8, u0_uk_K_r0_9, u0_uk_K_r10_0, u0_uk_K_r10_1, 
       u0_uk_K_r10_11, u0_uk_K_r10_12, u0_uk_K_r10_13, u0_uk_K_r10_14, u0_uk_K_r10_15, u0_uk_K_r10_16, u0_uk_K_r10_17, u0_uk_K_r10_19, u0_uk_K_r10_2, 
       u0_uk_K_r10_20, u0_uk_K_r10_21, u0_uk_K_r10_22, u0_uk_K_r10_24, u0_uk_K_r10_25, u0_uk_K_r10_26, u0_uk_K_r10_29, u0_uk_K_r10_3, u0_uk_K_r10_30, 
       u0_uk_K_r10_31, u0_uk_K_r10_33, u0_uk_K_r10_34, u0_uk_K_r10_35, u0_uk_K_r10_36, u0_uk_K_r10_38, u0_uk_K_r10_39, u0_uk_K_r10_4, u0_uk_K_r10_40, 
       u0_uk_K_r10_43, u0_uk_K_r10_45, u0_uk_K_r10_46, u0_uk_K_r10_47, u0_uk_K_r10_48, u0_uk_K_r10_49, u0_uk_K_r10_5, u0_uk_K_r10_50, u0_uk_K_r10_51, 
       u0_uk_K_r10_52, u0_uk_K_r10_53, u0_uk_K_r10_54, u0_uk_K_r10_55, u0_uk_K_r10_6, u0_uk_K_r10_7, u0_uk_K_r10_8, u0_uk_K_r11_0, u0_uk_K_r11_1, 
       u0_uk_K_r11_10, u0_uk_K_r11_11, u0_uk_K_r11_12, u0_uk_K_r11_13, u0_uk_K_r11_14, u0_uk_K_r11_15, u0_uk_K_r11_16, u0_uk_K_r11_17, u0_uk_K_r11_18, 
       u0_uk_K_r11_2, u0_uk_K_r11_21, u0_uk_K_r11_22, u0_uk_K_r11_23, u0_uk_K_r11_26, u0_uk_K_r11_28, u0_uk_K_r11_3, u0_uk_K_r11_30, u0_uk_K_r11_31, 
       u0_uk_K_r11_32, u0_uk_K_r11_34, u0_uk_K_r11_35, u0_uk_K_r11_36, u0_uk_K_r11_37, u0_uk_K_r11_38, u0_uk_K_r11_40, u0_uk_K_r11_41, u0_uk_K_r11_42, 
       u0_uk_K_r11_43, u0_uk_K_r11_44, u0_uk_K_r11_45, u0_uk_K_r11_46, u0_uk_K_r11_47, u0_uk_K_r11_48, u0_uk_K_r11_49, u0_uk_K_r11_5, u0_uk_K_r11_50, 
       u0_uk_K_r11_51, u0_uk_K_r11_52, u0_uk_K_r11_53, u0_uk_K_r11_54, u0_uk_K_r11_55, u0_uk_K_r11_6, u0_uk_K_r11_7, u0_uk_K_r11_8, u0_uk_K_r11_9, 
       u0_uk_K_r12_0, u0_uk_K_r12_1, u0_uk_K_r12_10, u0_uk_K_r12_11, u0_uk_K_r12_12, u0_uk_K_r12_13, u0_uk_K_r12_14, u0_uk_K_r12_15, u0_uk_K_r12_17, 
       u0_uk_K_r12_18, u0_uk_K_r12_19, u0_uk_K_r12_2, u0_uk_K_r12_20, u0_uk_K_r12_21, u0_uk_K_r12_22, u0_uk_K_r12_23, u0_uk_K_r12_24, u0_uk_K_r12_25, 
       u0_uk_K_r12_26, u0_uk_K_r12_27, u0_uk_K_r12_28, u0_uk_K_r12_29, u0_uk_K_r12_3, u0_uk_K_r12_30, u0_uk_K_r12_31, u0_uk_K_r12_32, u0_uk_K_r12_33, 
       u0_uk_K_r12_34, u0_uk_K_r12_35, u0_uk_K_r12_36, u0_uk_K_r12_37, u0_uk_K_r12_38, u0_uk_K_r12_39, u0_uk_K_r12_4, u0_uk_K_r12_40, u0_uk_K_r12_41, 
       u0_uk_K_r12_42, u0_uk_K_r12_43, u0_uk_K_r12_44, u0_uk_K_r12_45, u0_uk_K_r12_46, u0_uk_K_r12_47, u0_uk_K_r12_48, u0_uk_K_r12_49, u0_uk_K_r12_5, 
       u0_uk_K_r12_50, u0_uk_K_r12_51, u0_uk_K_r12_52, u0_uk_K_r12_53, u0_uk_K_r12_54, u0_uk_K_r12_55, u0_uk_K_r12_6, u0_uk_K_r12_7, u0_uk_K_r12_8, 
       u0_uk_K_r12_9, u0_uk_K_r13_1, u0_uk_K_r13_10, u0_uk_K_r13_11, u0_uk_K_r13_12, u0_uk_K_r13_13, u0_uk_K_r13_14, u0_uk_K_r13_15, u0_uk_K_r13_16, 
       u0_uk_K_r13_17, u0_uk_K_r13_18, u0_uk_K_r13_19, u0_uk_K_r13_2, u0_uk_K_r13_20, u0_uk_K_r13_21, u0_uk_K_r13_22, u0_uk_K_r13_23, u0_uk_K_r13_24, 
       u0_uk_K_r13_26, u0_uk_K_r13_27, u0_uk_K_r13_28, u0_uk_K_r13_29, u0_uk_K_r13_3, u0_uk_K_r13_30, u0_uk_K_r13_31, u0_uk_K_r13_32, u0_uk_K_r13_33, 
       u0_uk_K_r13_34, u0_uk_K_r13_35, u0_uk_K_r13_36, u0_uk_K_r13_37, u0_uk_K_r13_39, u0_uk_K_r13_4, u0_uk_K_r13_40, u0_uk_K_r13_41, u0_uk_K_r13_42, 
       u0_uk_K_r13_43, u0_uk_K_r13_45, u0_uk_K_r13_46, u0_uk_K_r13_47, u0_uk_K_r13_48, u0_uk_K_r13_49, u0_uk_K_r13_5, u0_uk_K_r13_50, u0_uk_K_r13_51, 
       u0_uk_K_r13_52, u0_uk_K_r13_53, u0_uk_K_r13_54, u0_uk_K_r13_55, u0_uk_K_r13_6, u0_uk_K_r13_7, u0_uk_K_r13_8, u0_uk_K_r13_9, u0_uk_K_r14_23, 
       u0_uk_K_r14_3, u0_uk_K_r14_38, u0_uk_K_r14_39, u0_uk_K_r14_42, u0_uk_K_r14_43, u0_uk_K_r14_46, u0_uk_K_r14_5, u0_uk_K_r1_0, u0_uk_K_r1_1, 
       u0_uk_K_r1_10, u0_uk_K_r1_11, u0_uk_K_r1_12, u0_uk_K_r1_13, u0_uk_K_r1_14, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_19, u0_uk_K_r1_2, 
       u0_uk_K_r1_20, u0_uk_K_r1_22, u0_uk_K_r1_23, u0_uk_K_r1_24, u0_uk_K_r1_25, u0_uk_K_r1_26, u0_uk_K_r1_27, u0_uk_K_r1_28, u0_uk_K_r1_29, 
       u0_uk_K_r1_3, u0_uk_K_r1_30, u0_uk_K_r1_31, u0_uk_K_r1_32, u0_uk_K_r1_33, u0_uk_K_r1_34, u0_uk_K_r1_35, u0_uk_K_r1_36, u0_uk_K_r1_37, 
       u0_uk_K_r1_38, u0_uk_K_r1_39, u0_uk_K_r1_4, u0_uk_K_r1_40, u0_uk_K_r1_41, u0_uk_K_r1_42, u0_uk_K_r1_43, u0_uk_K_r1_45, u0_uk_K_r1_46, 
       u0_uk_K_r1_47, u0_uk_K_r1_48, u0_uk_K_r1_49, u0_uk_K_r1_5, u0_uk_K_r1_50, u0_uk_K_r1_51, u0_uk_K_r1_52, u0_uk_K_r1_53, u0_uk_K_r1_54, 
       u0_uk_K_r1_55, u0_uk_K_r1_6, u0_uk_K_r1_8, u0_uk_K_r1_9, u0_uk_K_r2_0, u0_uk_K_r2_1, u0_uk_K_r2_10, u0_uk_K_r2_11, u0_uk_K_r2_12, 
       u0_uk_K_r2_14, u0_uk_K_r2_15, u0_uk_K_r2_16, u0_uk_K_r2_17, u0_uk_K_r2_19, u0_uk_K_r2_2, u0_uk_K_r2_21, u0_uk_K_r2_22, u0_uk_K_r2_23, 
       u0_uk_K_r2_24, u0_uk_K_r2_29, u0_uk_K_r2_3, u0_uk_K_r2_30, u0_uk_K_r2_31, u0_uk_K_r2_32, u0_uk_K_r2_34, u0_uk_K_r2_35, u0_uk_K_r2_36, 
       u0_uk_K_r2_37, u0_uk_K_r2_38, u0_uk_K_r2_39, u0_uk_K_r2_40, u0_uk_K_r2_42, u0_uk_K_r2_43, u0_uk_K_r2_44, u0_uk_K_r2_45, u0_uk_K_r2_47, 
       u0_uk_K_r2_48, u0_uk_K_r2_49, u0_uk_K_r2_5, u0_uk_K_r2_51, u0_uk_K_r2_52, u0_uk_K_r2_54, u0_uk_K_r2_6, u0_uk_K_r2_7, u0_uk_K_r2_8, 
       u0_uk_K_r2_9, u0_uk_K_r3_0, u0_uk_K_r3_1, u0_uk_K_r3_11, u0_uk_K_r3_12, u0_uk_K_r3_13, u0_uk_K_r3_15, u0_uk_K_r3_16, u0_uk_K_r3_17, 
       u0_uk_K_r3_18, u0_uk_K_r3_19, u0_uk_K_r3_2, u0_uk_K_r3_20, u0_uk_K_r3_21, u0_uk_K_r3_22, u0_uk_K_r3_23, u0_uk_K_r3_24, u0_uk_K_r3_25, 
       u0_uk_K_r3_26, u0_uk_K_r3_27, u0_uk_K_r3_28, u0_uk_K_r3_29, u0_uk_K_r3_3, u0_uk_K_r3_30, u0_uk_K_r3_31, u0_uk_K_r3_32, u0_uk_K_r3_33, 
       u0_uk_K_r3_34, u0_uk_K_r3_35, u0_uk_K_r3_36, u0_uk_K_r3_37, u0_uk_K_r3_38, u0_uk_K_r3_39, u0_uk_K_r3_4, u0_uk_K_r3_40, u0_uk_K_r3_41, 
       u0_uk_K_r3_42, u0_uk_K_r3_43, u0_uk_K_r3_44, u0_uk_K_r3_45, u0_uk_K_r3_46, u0_uk_K_r3_47, u0_uk_K_r3_48, u0_uk_K_r3_49, u0_uk_K_r3_5, 
       u0_uk_K_r3_50, u0_uk_K_r3_51, u0_uk_K_r3_52, u0_uk_K_r3_53, u0_uk_K_r3_54, u0_uk_K_r3_55, u0_uk_K_r3_6, u0_uk_K_r3_7, u0_uk_K_r3_8, 
       u0_uk_K_r3_9, u0_uk_K_r4_1, u0_uk_K_r4_10, u0_uk_K_r4_11, u0_uk_K_r4_12, u0_uk_K_r4_13, u0_uk_K_r4_14, u0_uk_K_r4_15, u0_uk_K_r4_16, 
       u0_uk_K_r4_17, u0_uk_K_r4_18, u0_uk_K_r4_19, u0_uk_K_r4_2, u0_uk_K_r4_20, u0_uk_K_r4_21, u0_uk_K_r4_22, u0_uk_K_r4_24, u0_uk_K_r4_25, 
       u0_uk_K_r4_26, u0_uk_K_r4_27, u0_uk_K_r4_28, u0_uk_K_r4_29, u0_uk_K_r4_3, u0_uk_K_r4_30, u0_uk_K_r4_31, u0_uk_K_r4_32, u0_uk_K_r4_34, 
       u0_uk_K_r4_36, u0_uk_K_r4_37, u0_uk_K_r4_39, u0_uk_K_r4_4, u0_uk_K_r4_40, u0_uk_K_r4_42, u0_uk_K_r4_43, u0_uk_K_r4_44, u0_uk_K_r4_45, 
       u0_uk_K_r4_46, u0_uk_K_r4_48, u0_uk_K_r4_49, u0_uk_K_r4_5, u0_uk_K_r4_50, u0_uk_K_r4_51, u0_uk_K_r4_52, u0_uk_K_r4_53, u0_uk_K_r4_54, 
       u0_uk_K_r4_55, u0_uk_K_r4_6, u0_uk_K_r4_7, u0_uk_K_r4_8, u0_uk_K_r4_9, u0_uk_K_r5_0, u0_uk_K_r5_1, u0_uk_K_r5_11, u0_uk_K_r5_12, 
       u0_uk_K_r5_13, u0_uk_K_r5_14, u0_uk_K_r5_15, u0_uk_K_r5_16, u0_uk_K_r5_18, u0_uk_K_r5_19, u0_uk_K_r5_2, u0_uk_K_r5_20, u0_uk_K_r5_21, 
       u0_uk_K_r5_22, u0_uk_K_r5_23, u0_uk_K_r5_24, u0_uk_K_r5_25, u0_uk_K_r5_26, u0_uk_K_r5_27, u0_uk_K_r5_28, u0_uk_K_r5_29, u0_uk_K_r5_3, 
       u0_uk_K_r5_30, u0_uk_K_r5_31, u0_uk_K_r5_32, u0_uk_K_r5_33, u0_uk_K_r5_34, u0_uk_K_r5_35, u0_uk_K_r5_36, u0_uk_K_r5_37, u0_uk_K_r5_38, 
       u0_uk_K_r5_40, u0_uk_K_r5_41, u0_uk_K_r5_42, u0_uk_K_r5_43, u0_uk_K_r5_44, u0_uk_K_r5_45, u0_uk_K_r5_46, u0_uk_K_r5_47, u0_uk_K_r5_48, 
       u0_uk_K_r5_49, u0_uk_K_r5_5, u0_uk_K_r5_50, u0_uk_K_r5_51, u0_uk_K_r5_52, u0_uk_K_r5_53, u0_uk_K_r5_54, u0_uk_K_r5_55, u0_uk_K_r5_6, 
       u0_uk_K_r5_7, u0_uk_K_r5_8, u0_uk_K_r5_9, u0_uk_K_r6_1, u0_uk_K_r6_10, u0_uk_K_r6_11, u0_uk_K_r6_12, u0_uk_K_r6_13, u0_uk_K_r6_14, 
       u0_uk_K_r6_15, u0_uk_K_r6_16, u0_uk_K_r6_17, u0_uk_K_r6_18, u0_uk_K_r6_19, u0_uk_K_r6_2, u0_uk_K_r6_20, u0_uk_K_r6_21, u0_uk_K_r6_23, 
       u0_uk_K_r6_24, u0_uk_K_r6_25, u0_uk_K_r6_27, u0_uk_K_r6_28, u0_uk_K_r6_29, u0_uk_K_r6_3, u0_uk_K_r6_30, u0_uk_K_r6_32, u0_uk_K_r6_33, 
       u0_uk_K_r6_35, u0_uk_K_r6_36, u0_uk_K_r6_37, u0_uk_K_r6_38, u0_uk_K_r6_39, u0_uk_K_r6_4, u0_uk_K_r6_40, u0_uk_K_r6_41, u0_uk_K_r6_42, 
       u0_uk_K_r6_43, u0_uk_K_r6_44, u0_uk_K_r6_45, u0_uk_K_r6_47, u0_uk_K_r6_48, u0_uk_K_r6_49, u0_uk_K_r6_5, u0_uk_K_r6_50, u0_uk_K_r6_51, 
       u0_uk_K_r6_52, u0_uk_K_r6_53, u0_uk_K_r6_54, u0_uk_K_r6_55, u0_uk_K_r6_6, u0_uk_K_r6_7, u0_uk_K_r6_8, u0_uk_K_r6_9, u0_uk_K_r7_0, 
       u0_uk_K_r7_1, u0_uk_K_r7_10, u0_uk_K_r7_11, u0_uk_K_r7_12, u0_uk_K_r7_13, u0_uk_K_r7_14, u0_uk_K_r7_15, u0_uk_K_r7_16, u0_uk_K_r7_17, 
       u0_uk_K_r7_18, u0_uk_K_r7_19, u0_uk_K_r7_2, u0_uk_K_r7_20, u0_uk_K_r7_21, u0_uk_K_r7_22, u0_uk_K_r7_23, u0_uk_K_r7_24, u0_uk_K_r7_25, 
       u0_uk_K_r7_27, u0_uk_K_r7_28, u0_uk_K_r7_29, u0_uk_K_r7_3, u0_uk_K_r7_30, u0_uk_K_r7_31, u0_uk_K_r7_32, u0_uk_K_r7_33, u0_uk_K_r7_34, 
       u0_uk_K_r7_35, u0_uk_K_r7_36, u0_uk_K_r7_37, u0_uk_K_r7_38, u0_uk_K_r7_39, u0_uk_K_r7_4, u0_uk_K_r7_40, u0_uk_K_r7_41, u0_uk_K_r7_42, 
       u0_uk_K_r7_43, u0_uk_K_r7_44, u0_uk_K_r7_45, u0_uk_K_r7_46, u0_uk_K_r7_47, u0_uk_K_r7_48, u0_uk_K_r7_49, u0_uk_K_r7_5, u0_uk_K_r7_50, 
       u0_uk_K_r7_51, u0_uk_K_r7_52, u0_uk_K_r7_53, u0_uk_K_r7_54, u0_uk_K_r7_55, u0_uk_K_r7_6, u0_uk_K_r7_7, u0_uk_K_r7_8, u0_uk_K_r7_9, 
       u0_uk_K_r8_0, u0_uk_K_r8_1, u0_uk_K_r8_10, u0_uk_K_r8_11, u0_uk_K_r8_12, u0_uk_K_r8_13, u0_uk_K_r8_14, u0_uk_K_r8_15, u0_uk_K_r8_17, 
       u0_uk_K_r8_18, u0_uk_K_r8_19, u0_uk_K_r8_2, u0_uk_K_r8_20, u0_uk_K_r8_21, u0_uk_K_r8_22, u0_uk_K_r8_23, u0_uk_K_r8_24, u0_uk_K_r8_25, 
       u0_uk_K_r8_26, u0_uk_K_r8_27, u0_uk_K_r8_28, u0_uk_K_r8_29, u0_uk_K_r8_3, u0_uk_K_r8_30, u0_uk_K_r8_31, u0_uk_K_r8_32, u0_uk_K_r8_33, 
       u0_uk_K_r8_34, u0_uk_K_r8_35, u0_uk_K_r8_36, u0_uk_K_r8_37, u0_uk_K_r8_38, u0_uk_K_r8_39, u0_uk_K_r8_4, u0_uk_K_r8_42, u0_uk_K_r8_43, 
       u0_uk_K_r8_44, u0_uk_K_r8_45, u0_uk_K_r8_46, u0_uk_K_r8_47, u0_uk_K_r8_48, u0_uk_K_r8_49, u0_uk_K_r8_5, u0_uk_K_r8_50, u0_uk_K_r8_51, 
       u0_uk_K_r8_52, u0_uk_K_r8_53, u0_uk_K_r8_54, u0_uk_K_r8_55, u0_uk_K_r8_6, u0_uk_K_r8_7, u0_uk_K_r8_8, u0_uk_K_r8_9, u0_uk_K_r9_10, 
       u0_uk_K_r9_11, u0_uk_K_r9_12, u0_uk_K_r9_13, u0_uk_K_r9_14, u0_uk_K_r9_15, u0_uk_K_r9_16, u0_uk_K_r9_17, u0_uk_K_r9_18, u0_uk_K_r9_2, 
       u0_uk_K_r9_20, u0_uk_K_r9_21, u0_uk_K_r9_23, u0_uk_K_r9_24, u0_uk_K_r9_26, u0_uk_K_r9_28, u0_uk_K_r9_29, u0_uk_K_r9_3, u0_uk_K_r9_31, 
       u0_uk_K_r9_32, u0_uk_K_r9_34, u0_uk_K_r9_36, u0_uk_K_r9_37, u0_uk_K_r9_38, u0_uk_K_r9_39, u0_uk_K_r9_4, u0_uk_K_r9_40, u0_uk_K_r9_41, 
       u0_uk_K_r9_42, u0_uk_K_r9_43, u0_uk_K_r9_44, u0_uk_K_r9_46, u0_uk_K_r9_47, u0_uk_K_r9_48, u0_uk_K_r9_49, u0_uk_K_r9_5, u0_uk_K_r9_50, 
       u0_uk_K_r9_51, u0_uk_K_r9_52, u0_uk_K_r9_53, u0_uk_K_r9_54, u0_uk_K_r9_55, u0_uk_K_r9_8, u0_uk_n1, u0_uk_n1007, u0_uk_n1008, 
       u0_uk_n1009, u0_uk_n1010, u0_uk_n1011, u0_uk_n1013, u0_uk_n1016, u0_uk_n1018, u0_uk_n1019, u0_uk_n1020, u0_uk_n1021, 
       u0_uk_n1022, u0_uk_n1023, u0_uk_n103, u0_uk_n104, u0_uk_n105, u0_uk_n111, u0_uk_n112, u0_uk_n114, u0_uk_n119, 
       u0_uk_n120, u0_uk_n124, u0_uk_n125, u0_uk_n130, u0_uk_n132, u0_uk_n133, u0_uk_n134, u0_uk_n135, u0_uk_n136, 
       u0_uk_n137, u0_uk_n138, u0_uk_n14, u0_uk_n140, u0_uk_n149, u0_uk_n15, u0_uk_n150, u0_uk_n152, u0_uk_n154, 
       u0_uk_n157, u0_uk_n158, u0_uk_n159, u0_uk_n16, u0_uk_n160, u0_uk_n165, u0_uk_n166, u0_uk_n169, u0_uk_n170, 
       u0_uk_n175, u0_uk_n176, u0_uk_n186, u0_uk_n19, u0_uk_n194, u0_uk_n2, u0_uk_n20, u0_uk_n226, u0_uk_n227, 
       u0_uk_n228, u0_uk_n229, u0_uk_n234, u0_uk_n235, u0_uk_n236, u0_uk_n237, u0_uk_n24, u0_uk_n245, u0_uk_n246, 
       u0_uk_n247, u0_uk_n25, u0_uk_n254, u0_uk_n255, u0_uk_n256, u0_uk_n258, u0_uk_n26, u0_uk_n262, u0_uk_n263, 
       u0_uk_n265, u0_uk_n268, u0_uk_n270, u0_uk_n273, u0_uk_n274, u0_uk_n280, u0_uk_n281, u0_uk_n284, u0_uk_n287, 
       u0_uk_n288, u0_uk_n29, u0_uk_n295, u0_uk_n296, u0_uk_n30, u0_uk_n302, u0_uk_n303, u0_uk_n304, u0_uk_n309, 
       u0_uk_n311, u0_uk_n315, u0_uk_n317, u0_uk_n321, u0_uk_n322, u0_uk_n323, u0_uk_n325, u0_uk_n326, u0_uk_n327, 
       u0_uk_n328, u0_uk_n333, u0_uk_n334, u0_uk_n34, u0_uk_n340, u0_uk_n343, u0_uk_n345, u0_uk_n35, u0_uk_n350, 
       u0_uk_n351, u0_uk_n354, u0_uk_n356, u0_uk_n357, u0_uk_n359, u0_uk_n36, u0_uk_n360, u0_uk_n362, u0_uk_n364, 
       u0_uk_n365, u0_uk_n367, u0_uk_n368, u0_uk_n37, u0_uk_n372, u0_uk_n374, u0_uk_n378, u0_uk_n38, u0_uk_n380, 
       u0_uk_n381, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n390, u0_uk_n394, u0_uk_n397, u0_uk_n398, u0_uk_n399, 
       u0_uk_n402, u0_uk_n403, u0_uk_n404, u0_uk_n406, u0_uk_n416, u0_uk_n417, u0_uk_n42, u0_uk_n422, u0_uk_n427, 
       u0_uk_n43, u0_uk_n431, u0_uk_n435, u0_uk_n44, u0_uk_n441, u0_uk_n444, u0_uk_n449, u0_uk_n451, u0_uk_n452, 
       u0_uk_n453, u0_uk_n455, u0_uk_n458, u0_uk_n459, u0_uk_n46, u0_uk_n461, u0_uk_n462, u0_uk_n463, u0_uk_n464, 
       u0_uk_n465, u0_uk_n466, u0_uk_n469, u0_uk_n47, u0_uk_n470, u0_uk_n473, u0_uk_n474, u0_uk_n475, u0_uk_n476, 
       u0_uk_n477, u0_uk_n478, u0_uk_n479, u0_uk_n48, u0_uk_n480, u0_uk_n481, u0_uk_n482, u0_uk_n483, u0_uk_n484, 
       u0_uk_n485, u0_uk_n486, u0_uk_n487, u0_uk_n488, u0_uk_n489, u0_uk_n49, u0_uk_n490, u0_uk_n491, u0_uk_n492, 
       u0_uk_n493, u0_uk_n494, u0_uk_n495, u0_uk_n498, u0_uk_n50, u0_uk_n506, u0_uk_n507, u0_uk_n51, u0_uk_n512, 
       u0_uk_n514, u0_uk_n516, u0_uk_n52, u0_uk_n521, u0_uk_n527, u0_uk_n528, u0_uk_n53, u0_uk_n533, u0_uk_n537, 
       u0_uk_n538, u0_uk_n54, u0_uk_n540, u0_uk_n541, u0_uk_n543, u0_uk_n548, u0_uk_n556, u0_uk_n559, u0_uk_n56, 
       u0_uk_n563, u0_uk_n564, u0_uk_n569, u0_uk_n57, u0_uk_n571, u0_uk_n572, u0_uk_n576, u0_uk_n584, u0_uk_n585, 
       u0_uk_n588, u0_uk_n589, u0_uk_n59, u0_uk_n591, u0_uk_n592, u0_uk_n593, u0_uk_n594, u0_uk_n595, u0_uk_n596, 
       u0_uk_n597, u0_uk_n599, u0_uk_n6, u0_uk_n600, u0_uk_n602, u0_uk_n606, u0_uk_n607, u0_uk_n609, u0_uk_n610, 
       u0_uk_n611, u0_uk_n612, u0_uk_n613, u0_uk_n614, u0_uk_n616, u0_uk_n617, u0_uk_n618, u0_uk_n619, u0_uk_n62, 
       u0_uk_n620, u0_uk_n621, u0_uk_n622, u0_uk_n623, u0_uk_n624, u0_uk_n625, u0_uk_n626, u0_uk_n628, u0_uk_n630, 
       u0_uk_n631, u0_uk_n633, u0_uk_n638, u0_uk_n64, u0_uk_n641, u0_uk_n646, u0_uk_n647, u0_uk_n648, u0_uk_n65, 
       u0_uk_n655, u0_uk_n66, u0_uk_n664, u0_uk_n667, u0_uk_n68, u0_uk_n680, u0_uk_n69, u0_uk_n691, u0_uk_n698, 
       u0_uk_n7, u0_uk_n70, u0_uk_n705, u0_uk_n707, u0_uk_n71, u0_uk_n710, u0_uk_n715, u0_uk_n718, u0_uk_n72, 
       u0_uk_n720, u0_uk_n721, u0_uk_n724, u0_uk_n728, u0_uk_n730, u0_uk_n732, u0_uk_n733, u0_uk_n736, u0_uk_n738, 
       u0_uk_n739, u0_uk_n74, u0_uk_n740, u0_uk_n742, u0_uk_n743, u0_uk_n744, u0_uk_n749, u0_uk_n75, u0_uk_n752, 
       u0_uk_n753, u0_uk_n754, u0_uk_n755, u0_uk_n756, u0_uk_n76, u0_uk_n762, u0_uk_n765, u0_uk_n766, u0_uk_n767, 
       u0_uk_n769, u0_uk_n77, u0_uk_n770, u0_uk_n771, u0_uk_n772, u0_uk_n773, u0_uk_n774, u0_uk_n775, u0_uk_n776, 
       u0_uk_n777, u0_uk_n778, u0_uk_n779, u0_uk_n78, u0_uk_n782, u0_uk_n785, u0_uk_n79, u0_uk_n790, u0_uk_n792, 
       u0_uk_n796, u0_uk_n797, u0_uk_n798, u0_uk_n80, u0_uk_n801, u0_uk_n802, u0_uk_n804, u0_uk_n805, u0_uk_n806, 
       u0_uk_n807, u0_uk_n808, u0_uk_n81, u0_uk_n812, u0_uk_n814, u0_uk_n817, u0_uk_n818, u0_uk_n82, u0_uk_n820, 
       u0_uk_n823, u0_uk_n826, u0_uk_n829, u0_uk_n830, u0_uk_n831, u0_uk_n834, u0_uk_n84, u0_uk_n840, u0_uk_n841, 
       u0_uk_n842, u0_uk_n846, u0_uk_n848, u0_uk_n85, u0_uk_n850, u0_uk_n851, u0_uk_n852, u0_uk_n853, u0_uk_n854, 
       u0_uk_n856, u0_uk_n857, u0_uk_n859, u0_uk_n86, u0_uk_n863, u0_uk_n864, u0_uk_n865, u0_uk_n867, u0_uk_n87, 
       u0_uk_n871, u0_uk_n872, u0_uk_n873, u0_uk_n878, u0_uk_n88, u0_uk_n880, u0_uk_n884, u0_uk_n885, u0_uk_n888, 
       u0_uk_n889, u0_uk_n89, u0_uk_n890, u0_uk_n894, u0_uk_n895, u0_uk_n897, u0_uk_n90, u0_uk_n906, u0_uk_n909, 
       u0_uk_n911, u0_uk_n912, u0_uk_n913, u0_uk_n914, u0_uk_n921, u0_uk_n922, u0_uk_n923, u0_uk_n925, u0_uk_n926, 
       u0_uk_n927, u0_uk_n928, u0_uk_n930, u0_uk_n931, u0_uk_n932, u0_uk_n935, u0_uk_n936, u0_uk_n937, u0_uk_n938, 
       u0_uk_n939, u0_uk_n941, u0_uk_n942, u0_uk_n945, u0_uk_n946, u0_uk_n947, u0_uk_n948, u0_uk_n95, u0_uk_n957, 
       u0_uk_n958, u0_uk_n959, u0_uk_n960, u0_uk_n961, u0_uk_n964, u0_uk_n967, u0_uk_n969, u0_uk_n97, u0_uk_n970, 
       u0_uk_n971, u0_uk_n977, u0_uk_n978, u0_uk_n980, u0_uk_n981, u0_uk_n987, u0_uk_n989, u0_uk_n991, u0_uk_n997, 
       u0_uk_n998, u1_FP_1, u1_FP_10, u1_FP_11, u1_FP_12, u1_FP_13, u1_FP_14, u1_FP_15, u1_FP_16, 
       u1_FP_17, u1_FP_18, u1_FP_19, u1_FP_2, u1_FP_20, u1_FP_21, u1_FP_22, u1_FP_23, u1_FP_24, 
       u1_FP_25, u1_FP_26, u1_FP_27, u1_FP_28, u1_FP_29, u1_FP_3, u1_FP_30, u1_FP_31, u1_FP_32, 
       u1_FP_34, u1_FP_35, u1_FP_36, u1_FP_38, u1_FP_39, u1_FP_4, u1_FP_42, u1_FP_43, u1_FP_46, 
       u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_5, u1_FP_50, u1_FP_51, u1_FP_54, u1_FP_57, u1_FP_58, 
       u1_FP_59, u1_FP_6, u1_FP_62, u1_FP_63, u1_FP_64, u1_FP_7, u1_FP_8, u1_FP_9, u1_K10_10, 
       u1_K10_15, u1_K10_16, u1_K10_17, u1_K10_19, u1_K10_21, u1_K10_27, u1_K10_28, u1_K10_3, u1_K10_34, 
       u1_K10_39, u1_K10_4, u1_K10_40, u1_K10_45, u1_K10_46, u1_K11_1, u1_K11_10, u1_K11_15, u1_K11_16, 
       u1_K11_18, u1_K11_20, u1_K11_21, u1_K11_24, u1_K11_26, u1_K11_27, u1_K11_28, u1_K11_3, u1_K11_33, 
       u1_K11_39, u1_K11_4, u1_K11_40, u1_K11_41, u1_K11_42, u1_K11_43, u1_K11_44, u1_K11_45, u1_K11_46, 
       u1_K11_47, u1_K11_6, u1_K11_8, u1_K11_9, u1_K12_10, u1_K12_11, u1_K12_12, u1_K12_13, u1_K12_14, 
       u1_K12_16, u1_K12_22, u1_K12_27, u1_K12_28, u1_K12_29, u1_K12_3, u1_K12_30, u1_K12_31, u1_K12_32, 
       u1_K12_33, u1_K12_34, u1_K12_39, u1_K12_4, u1_K12_40, u1_K12_45, u1_K12_46, u1_K12_5, u1_K12_7, 
       u1_K12_9, u1_K13_1, u1_K13_10, u1_K13_16, u1_K13_21, u1_K13_22, u1_K13_23, u1_K13_24, u1_K13_25, 
       u1_K13_26, u1_K13_27, u1_K13_28, u1_K13_3, u1_K13_33, u1_K13_34, u1_K13_36, u1_K13_38, u1_K13_39, 
       u1_K13_4, u1_K13_40, u1_K13_41, u1_K13_42, u1_K13_43, u1_K13_44, u1_K13_45, u1_K13_46, u1_K13_47, 
       u1_K13_9, u1_K14_10, u1_K14_11, u1_K14_12, u1_K14_13, u1_K14_14, u1_K14_15, u1_K14_16, u1_K14_17, 
       u1_K14_18, u1_K14_19, u1_K14_20, u1_K14_21, u1_K14_22, u1_K14_23, u1_K14_24, u1_K14_25, u1_K14_26, 
       u1_K14_27, u1_K14_28, u1_K14_3, u1_K14_33, u1_K14_35, u1_K14_36, u1_K14_37, u1_K14_38, u1_K14_39, 
       u1_K14_4, u1_K14_40, u1_K14_41, u1_K14_43, u1_K14_45, u1_K14_46, u1_K14_5, u1_K14_6, u1_K14_7, 
       u1_K14_8, u1_K14_9, u1_K15_1, u1_K15_10, u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_19, u1_K15_21, 
       u1_K15_22, u1_K15_27, u1_K15_28, u1_K15_3, u1_K15_33, u1_K15_34, u1_K15_39, u1_K15_4, u1_K15_40, 
       u1_K15_45, u1_K15_46, u1_K15_47, u1_K15_9, u1_K16_1, u1_K16_10, u1_K16_15, u1_K16_16, u1_K16_21, 
       u1_K16_22, u1_K16_23, u1_K16_24, u1_K16_25, u1_K16_26, u1_K16_27, u1_K16_28, u1_K16_3, u1_K16_33, 
       u1_K16_36, u1_K16_38, u1_K16_39, u1_K16_4, u1_K16_40, u1_K16_45, u1_K16_46, u1_K16_47, u1_K16_5, 
       u1_K16_7, u1_K16_9, u1_K1_10, u1_K1_11, u1_K1_12, u1_K1_13, u1_K1_14, u1_K1_15, u1_K1_16, 
       u1_K1_2, u1_K1_21, u1_K1_22, u1_K1_23, u1_K1_24, u1_K1_25, u1_K1_26, u1_K1_27, u1_K1_28, 
       u1_K1_29, u1_K1_3, u1_K1_30, u1_K1_31, u1_K1_32, u1_K1_33, u1_K1_34, u1_K1_35, u1_K1_36, 
       u1_K1_37, u1_K1_38, u1_K1_39, u1_K1_4, u1_K1_40, u1_K1_42, u1_K1_44, u1_K1_45, u1_K1_46, 
       u1_K1_48, u1_K1_5, u1_K1_7, u1_K1_9, u1_K2_15, u1_K2_16, u1_K2_21, u1_K2_22, u1_K2_27, 
       u1_K2_28, u1_K2_3, u1_K2_33, u1_K2_34, u1_K2_35, u1_K2_36, u1_K2_37, u1_K2_38, u1_K2_39, 
       u1_K2_4, u1_K2_40, u1_K2_45, u1_K2_46, u1_K2_9, u1_K3_10, u1_K3_11, u1_K3_13, u1_K3_15, 
       u1_K3_16, u1_K3_21, u1_K3_22, u1_K3_27, u1_K3_28, u1_K3_3, u1_K3_30, u1_K3_32, u1_K3_33, 
       u1_K3_34, u1_K3_39, u1_K3_4, u1_K3_40, u1_K3_45, u1_K3_46, u1_K3_9, u1_K4_15, u1_K4_16, 
       u1_K4_21, u1_K4_22, u1_K4_27, u1_K4_28, u1_K4_33, u1_K4_34, u1_K4_39, u1_K4_4, u1_K4_40, 
       u1_K4_45, u1_K4_46, u1_K4_5, u1_K4_7, u1_K4_9, u1_K5_10, u1_K5_15, u1_K5_16, u1_K5_21, 
       u1_K5_28, u1_K5_3, u1_K5_33, u1_K5_34, u1_K5_39, u1_K5_4, u1_K5_40, u1_K5_45, u1_K5_46, 
       u1_K5_9, u1_K6_15, u1_K6_16, u1_K6_17, u1_K6_19, u1_K6_22, u1_K6_27, u1_K6_28, u1_K6_3, 
       u1_K6_33, u1_K6_34, u1_K6_39, u1_K6_40, u1_K6_45, u1_K6_46, u1_K7_10, u1_K7_15, u1_K7_16, 
       u1_K7_21, u1_K7_22, u1_K7_28, u1_K7_3, u1_K7_33, u1_K7_39, u1_K7_4, u1_K7_40, u1_K7_45, 
       u1_K7_9, u1_K8_10, u1_K8_16, u1_K8_17, u1_K8_19, u1_K8_21, u1_K8_22, u1_K8_27, u1_K8_28, 
       u1_K8_33, u1_K8_34, u1_K8_39, u1_K8_4, u1_K8_40, u1_K8_45, u1_K8_46, u1_K8_6, u1_K8_8, 
       u1_K8_9, u1_K9_15, u1_K9_16, u1_K9_21, u1_K9_28, u1_K9_3, u1_K9_30, u1_K9_32, u1_K9_33, 
       u1_K9_34, u1_K9_39, u1_K9_4, u1_K9_40, u1_K9_45, u1_K9_46, u1_L0_1, u1_L0_10, u1_L0_11, 
       u1_L0_12, u1_L0_13, u1_L0_14, u1_L0_15, u1_L0_16, u1_L0_17, u1_L0_18, u1_L0_19, u1_L0_2, 
       u1_L0_20, u1_L0_21, u1_L0_22, u1_L0_23, u1_L0_24, u1_L0_25, u1_L0_26, u1_L0_27, u1_L0_28, 
       u1_L0_29, u1_L0_3, u1_L0_30, u1_L0_31, u1_L0_32, u1_L0_4, u1_L0_5, u1_L0_6, u1_L0_7, 
       u1_L0_8, u1_L0_9, u1_L10_1, u1_L10_10, u1_L10_11, u1_L10_12, u1_L10_13, u1_L10_14, u1_L10_15, 
       u1_L10_16, u1_L10_17, u1_L10_18, u1_L10_19, u1_L10_2, u1_L10_20, u1_L10_21, u1_L10_22, u1_L10_23, 
       u1_L10_24, u1_L10_25, u1_L10_26, u1_L10_27, u1_L10_28, u1_L10_29, u1_L10_3, u1_L10_30, u1_L10_31, 
       u1_L10_32, u1_L10_4, u1_L10_5, u1_L10_6, u1_L10_7, u1_L10_8, u1_L10_9, u1_L11_1, u1_L11_10, 
       u1_L11_11, u1_L11_12, u1_L11_13, u1_L11_14, u1_L11_15, u1_L11_16, u1_L11_17, u1_L11_18, u1_L11_19, 
       u1_L11_2, u1_L11_20, u1_L11_21, u1_L11_22, u1_L11_23, u1_L11_24, u1_L11_25, u1_L11_26, u1_L11_27, 
       u1_L11_28, u1_L11_29, u1_L11_3, u1_L11_30, u1_L11_31, u1_L11_32, u1_L11_4, u1_L11_5, u1_L11_6, 
       u1_L11_7, u1_L11_8, u1_L11_9, u1_L12_1, u1_L12_10, u1_L12_11, u1_L12_12, u1_L12_13, u1_L12_14, 
       u1_L12_15, u1_L12_16, u1_L12_17, u1_L12_18, u1_L12_19, u1_L12_2, u1_L12_20, u1_L12_21, u1_L12_22, 
       u1_L12_23, u1_L12_24, u1_L12_25, u1_L12_26, u1_L12_27, u1_L12_28, u1_L12_29, u1_L12_3, u1_L12_30, 
       u1_L12_31, u1_L12_32, u1_L12_4, u1_L12_5, u1_L12_6, u1_L12_7, u1_L12_8, u1_L12_9, u1_L13_1, 
       u1_L13_10, u1_L13_11, u1_L13_12, u1_L13_13, u1_L13_14, u1_L13_15, u1_L13_16, u1_L13_17, u1_L13_18, 
       u1_L13_19, u1_L13_2, u1_L13_20, u1_L13_21, u1_L13_22, u1_L13_23, u1_L13_24, u1_L13_25, u1_L13_26, 
       u1_L13_27, u1_L13_28, u1_L13_29, u1_L13_3, u1_L13_30, u1_L13_31, u1_L13_32, u1_L13_4, u1_L13_5, 
       u1_L13_6, u1_L13_7, u1_L13_8, u1_L13_9, u1_L14_1, u1_L14_10, u1_L14_11, u1_L14_12, u1_L14_13, 
       u1_L14_14, u1_L14_15, u1_L14_16, u1_L14_17, u1_L14_18, u1_L14_19, u1_L14_2, u1_L14_20, u1_L14_21, 
       u1_L14_22, u1_L14_23, u1_L14_24, u1_L14_25, u1_L14_26, u1_L14_27, u1_L14_28, u1_L14_29, u1_L14_3, 
       u1_L14_30, u1_L14_31, u1_L14_32, u1_L14_4, u1_L14_5, u1_L14_6, u1_L14_7, u1_L14_8, u1_L14_9, 
       u1_L1_1, u1_L1_10, u1_L1_11, u1_L1_12, u1_L1_13, u1_L1_14, u1_L1_15, u1_L1_16, u1_L1_17, 
       u1_L1_18, u1_L1_19, u1_L1_2, u1_L1_20, u1_L1_21, u1_L1_22, u1_L1_23, u1_L1_24, u1_L1_25, 
       u1_L1_26, u1_L1_27, u1_L1_28, u1_L1_29, u1_L1_3, u1_L1_30, u1_L1_31, u1_L1_32, u1_L1_4, 
       u1_L1_5, u1_L1_6, u1_L1_7, u1_L1_8, u1_L1_9, u1_L2_1, u1_L2_10, u1_L2_11, u1_L2_12, 
       u1_L2_13, u1_L2_14, u1_L2_15, u1_L2_16, u1_L2_17, u1_L2_18, u1_L2_19, u1_L2_2, u1_L2_20, 
       u1_L2_21, u1_L2_22, u1_L2_23, u1_L2_24, u1_L2_25, u1_L2_26, u1_L2_27, u1_L2_28, u1_L2_29, 
       u1_L2_3, u1_L2_30, u1_L2_31, u1_L2_32, u1_L2_4, u1_L2_5, u1_L2_6, u1_L2_7, u1_L2_8, 
       u1_L2_9, u1_L3_1, u1_L3_10, u1_L3_11, u1_L3_12, u1_L3_13, u1_L3_14, u1_L3_15, u1_L3_16, 
       u1_L3_17, u1_L3_18, u1_L3_19, u1_L3_2, u1_L3_20, u1_L3_21, u1_L3_22, u1_L3_23, u1_L3_24, 
       u1_L3_25, u1_L3_26, u1_L3_27, u1_L3_28, u1_L3_29, u1_L3_3, u1_L3_30, u1_L3_31, u1_L3_32, 
       u1_L3_4, u1_L3_5, u1_L3_6, u1_L3_7, u1_L3_8, u1_L3_9, u1_L4_1, u1_L4_10, u1_L4_11, 
       u1_L4_12, u1_L4_13, u1_L4_14, u1_L4_15, u1_L4_16, u1_L4_17, u1_L4_18, u1_L4_19, u1_L4_2, 
       u1_L4_20, u1_L4_21, u1_L4_22, u1_L4_23, u1_L4_24, u1_L4_25, u1_L4_26, u1_L4_27, u1_L4_28, 
       u1_L4_29, u1_L4_3, u1_L4_30, u1_L4_31, u1_L4_32, u1_L4_4, u1_L4_5, u1_L4_6, u1_L4_7, 
       u1_L4_8, u1_L4_9, u1_L5_1, u1_L5_10, u1_L5_11, u1_L5_12, u1_L5_13, u1_L5_14, u1_L5_15, 
       u1_L5_16, u1_L5_17, u1_L5_18, u1_L5_19, u1_L5_2, u1_L5_20, u1_L5_21, u1_L5_22, u1_L5_23, 
       u1_L5_24, u1_L5_25, u1_L5_26, u1_L5_27, u1_L5_28, u1_L5_29, u1_L5_3, u1_L5_30, u1_L5_31, 
       u1_L5_32, u1_L5_4, u1_L5_5, u1_L5_6, u1_L5_7, u1_L5_8, u1_L5_9, u1_L6_1, u1_L6_10, 
       u1_L6_11, u1_L6_12, u1_L6_13, u1_L6_14, u1_L6_15, u1_L6_16, u1_L6_17, u1_L6_18, u1_L6_19, 
       u1_L6_2, u1_L6_20, u1_L6_21, u1_L6_22, u1_L6_23, u1_L6_24, u1_L6_25, u1_L6_26, u1_L6_27, 
       u1_L6_28, u1_L6_29, u1_L6_3, u1_L6_30, u1_L6_31, u1_L6_32, u1_L6_4, u1_L6_5, u1_L6_6, 
       u1_L6_7, u1_L6_8, u1_L6_9, u1_L7_1, u1_L7_10, u1_L7_11, u1_L7_12, u1_L7_13, u1_L7_14, 
       u1_L7_15, u1_L7_16, u1_L7_17, u1_L7_18, u1_L7_19, u1_L7_2, u1_L7_20, u1_L7_21, u1_L7_22, 
       u1_L7_23, u1_L7_24, u1_L7_25, u1_L7_26, u1_L7_27, u1_L7_28, u1_L7_29, u1_L7_3, u1_L7_30, 
       u1_L7_31, u1_L7_32, u1_L7_4, u1_L7_5, u1_L7_6, u1_L7_7, u1_L7_8, u1_L7_9, u1_L8_1, 
       u1_L8_10, u1_L8_11, u1_L8_12, u1_L8_13, u1_L8_14, u1_L8_15, u1_L8_16, u1_L8_17, u1_L8_18, 
       u1_L8_19, u1_L8_2, u1_L8_20, u1_L8_21, u1_L8_22, u1_L8_23, u1_L8_24, u1_L8_25, u1_L8_26, 
       u1_L8_27, u1_L8_28, u1_L8_29, u1_L8_3, u1_L8_30, u1_L8_31, u1_L8_32, u1_L8_4, u1_L8_5, 
       u1_L8_6, u1_L8_7, u1_L8_8, u1_L8_9, u1_L9_1, u1_L9_10, u1_L9_11, u1_L9_12, u1_L9_13, 
       u1_L9_14, u1_L9_15, u1_L9_16, u1_L9_17, u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_20, u1_L9_21, 
       u1_L9_22, u1_L9_23, u1_L9_24, u1_L9_25, u1_L9_26, u1_L9_27, u1_L9_28, u1_L9_29, u1_L9_3, 
       u1_L9_30, u1_L9_31, u1_L9_32, u1_L9_4, u1_L9_5, u1_L9_6, u1_L9_7, u1_L9_8, u1_L9_9, 
       u1_N0, u1_N1, u1_N10, u1_N100, u1_N101, u1_N102, u1_N103, u1_N104, u1_N105, 
       u1_N106, u1_N107, u1_N108, u1_N109, u1_N11, u1_N110, u1_N111, u1_N112, u1_N113, 
       u1_N114, u1_N115, u1_N116, u1_N117, u1_N118, u1_N119, u1_N12, u1_N120, u1_N121, 
       u1_N122, u1_N123, u1_N124, u1_N125, u1_N126, u1_N127, u1_N128, u1_N129, u1_N13, 
       u1_N130, u1_N131, u1_N132, u1_N133, u1_N134, u1_N135, u1_N136, u1_N137, u1_N138, 
       u1_N139, u1_N14, u1_N140, u1_N141, u1_N142, u1_N143, u1_N144, u1_N145, u1_N146, 
       u1_N147, u1_N148, u1_N149, u1_N15, u1_N150, u1_N151, u1_N152, u1_N153, u1_N154, 
       u1_N155, u1_N156, u1_N157, u1_N158, u1_N159, u1_N16, u1_N160, u1_N161, u1_N162, 
       u1_N163, u1_N164, u1_N165, u1_N166, u1_N167, u1_N168, u1_N169, u1_N17, u1_N170, 
       u1_N171, u1_N172, u1_N173, u1_N174, u1_N175, u1_N176, u1_N177, u1_N178, u1_N179, 
       u1_N18, u1_N180, u1_N181, u1_N182, u1_N183, u1_N184, u1_N185, u1_N186, u1_N187, 
       u1_N188, u1_N189, u1_N19, u1_N190, u1_N191, u1_N192, u1_N193, u1_N194, u1_N195, 
       u1_N196, u1_N197, u1_N198, u1_N199, u1_N2, u1_N20, u1_N200, u1_N201, u1_N202, 
       u1_N203, u1_N204, u1_N205, u1_N206, u1_N207, u1_N208, u1_N209, u1_N21, u1_N210, 
       u1_N211, u1_N212, u1_N213, u1_N214, u1_N215, u1_N216, u1_N217, u1_N218, u1_N219, 
       u1_N22, u1_N220, u1_N221, u1_N222, u1_N223, u1_N224, u1_N225, u1_N226, u1_N227, 
       u1_N228, u1_N229, u1_N23, u1_N230, u1_N231, u1_N232, u1_N233, u1_N234, u1_N235, 
       u1_N236, u1_N237, u1_N238, u1_N239, u1_N24, u1_N240, u1_N241, u1_N242, u1_N243, 
       u1_N244, u1_N245, u1_N246, u1_N247, u1_N248, u1_N249, u1_N25, u1_N250, u1_N251, 
       u1_N252, u1_N253, u1_N254, u1_N255, u1_N256, u1_N257, u1_N258, u1_N259, u1_N26, 
       u1_N260, u1_N261, u1_N262, u1_N263, u1_N264, u1_N265, u1_N266, u1_N267, u1_N268, 
       u1_N269, u1_N27, u1_N270, u1_N271, u1_N272, u1_N273, u1_N274, u1_N275, u1_N276, 
       u1_N277, u1_N278, u1_N279, u1_N28, u1_N280, u1_N281, u1_N282, u1_N283, u1_N284, 
       u1_N285, u1_N286, u1_N287, u1_N288, u1_N289, u1_N29, u1_N290, u1_N291, u1_N292, 
       u1_N293, u1_N294, u1_N295, u1_N296, u1_N297, u1_N298, u1_N299, u1_N3, u1_N30, 
       u1_N300, u1_N301, u1_N302, u1_N303, u1_N304, u1_N305, u1_N306, u1_N307, u1_N308, 
       u1_N309, u1_N31, u1_N310, u1_N311, u1_N312, u1_N313, u1_N314, u1_N315, u1_N316, 
       u1_N317, u1_N318, u1_N319, u1_N32, u1_N320, u1_N321, u1_N322, u1_N323, u1_N324, 
       u1_N325, u1_N326, u1_N327, u1_N328, u1_N329, u1_N33, u1_N330, u1_N331, u1_N332, 
       u1_N333, u1_N334, u1_N335, u1_N336, u1_N337, u1_N338, u1_N339, u1_N34, u1_N340, 
       u1_N341, u1_N342, u1_N343, u1_N344, u1_N345, u1_N346, u1_N347, u1_N348, u1_N349, 
       u1_N35, u1_N350, u1_N351, u1_N352, u1_N353, u1_N354, u1_N355, u1_N356, u1_N357, 
       u1_N358, u1_N359, u1_N36, u1_N360, u1_N361, u1_N362, u1_N363, u1_N364, u1_N365, 
       u1_N366, u1_N367, u1_N368, u1_N369, u1_N37, u1_N370, u1_N371, u1_N372, u1_N373, 
       u1_N374, u1_N375, u1_N376, u1_N377, u1_N378, u1_N379, u1_N38, u1_N380, u1_N381, 
       u1_N382, u1_N383, u1_N384, u1_N385, u1_N386, u1_N387, u1_N388, u1_N389, u1_N39, 
       u1_N390, u1_N391, u1_N392, u1_N393, u1_N394, u1_N395, u1_N396, u1_N397, u1_N398, 
       u1_N399, u1_N4, u1_N40, u1_N400, u1_N401, u1_N402, u1_N403, u1_N404, u1_N405, 
       u1_N406, u1_N407, u1_N408, u1_N409, u1_N41, u1_N410, u1_N411, u1_N412, u1_N413, 
       u1_N414, u1_N415, u1_N416, u1_N417, u1_N418, u1_N419, u1_N42, u1_N420, u1_N421, 
       u1_N422, u1_N423, u1_N424, u1_N425, u1_N426, u1_N427, u1_N428, u1_N429, u1_N43, 
       u1_N430, u1_N431, u1_N432, u1_N433, u1_N434, u1_N435, u1_N436, u1_N437, u1_N438, 
       u1_N439, u1_N44, u1_N440, u1_N441, u1_N442, u1_N443, u1_N444, u1_N445, u1_N446, 
       u1_N447, u1_N448, u1_N449, u1_N45, u1_N450, u1_N451, u1_N452, u1_N453, u1_N454, 
       u1_N455, u1_N456, u1_N457, u1_N458, u1_N459, u1_N46, u1_N460, u1_N461, u1_N462, 
       u1_N463, u1_N464, u1_N465, u1_N466, u1_N467, u1_N468, u1_N469, u1_N47, u1_N470, 
       u1_N471, u1_N472, u1_N473, u1_N474, u1_N475, u1_N476, u1_N477, u1_N478, u1_N479, 
       u1_N48, u1_N49, u1_N5, u1_N50, u1_N51, u1_N52, u1_N53, u1_N54, u1_N55, 
       u1_N56, u1_N57, u1_N58, u1_N59, u1_N6, u1_N60, u1_N61, u1_N62, u1_N63, 
       u1_N64, u1_N65, u1_N66, u1_N67, u1_N68, u1_N69, u1_N7, u1_N70, u1_N71, 
       u1_N72, u1_N73, u1_N74, u1_N75, u1_N76, u1_N77, u1_N78, u1_N79, u1_N8, 
       u1_N80, u1_N81, u1_N82, u1_N83, u1_N84, u1_N85, u1_N86, u1_N87, u1_N88, 
       u1_N89, u1_N9, u1_N90, u1_N91, u1_N92, u1_N93, u1_N94, u1_N95, u1_N96, 
       u1_N97, u1_N98, u1_N99, u1_R0_10, u1_R0_11, u1_R0_14, u1_R0_15, u1_R0_18, u1_R0_19, 
       u1_R0_2, u1_R0_22, u1_R0_23, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_3, u1_R0_30, 
       u1_R0_31, u1_R0_6, u1_R10_11, u1_R10_15, u1_R10_18, u1_R10_19, u1_R10_2, u1_R10_20, u1_R10_21, 
       u1_R10_22, u1_R10_23, u1_R10_26, u1_R10_27, u1_R10_3, u1_R10_30, u1_R10_31, u1_R10_4, u1_R10_6, 
       u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_11, u1_R11_14, u1_R11_15, u1_R11_16, u1_R11_17, u1_R11_18, 
       u1_R11_19, u1_R11_2, u1_R11_22, u1_R11_23, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, u1_R11_29, 
       u1_R11_3, u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_6, u1_R11_7, u1_R12_10, u1_R12_11, u1_R12_12, 
       u1_R12_13, u1_R12_14, u1_R12_15, u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, u1_R12_2, u1_R12_22, 
       u1_R12_24, u1_R12_25, u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_3, u1_R12_30, u1_R12_31, u1_R12_4, 
       u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_14, 
       u1_R13_15, u1_R13_18, u1_R13_19, u1_R13_2, u1_R13_22, u1_R13_23, u1_R13_26, u1_R13_27, u1_R13_3, 
       u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_6, u1_R13_7, u1_R1_10, u1_R1_11, u1_R1_14, u1_R1_15, 
       u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_21, u1_R1_22, u1_R1_23, u1_R1_26, u1_R1_27, u1_R1_3, 
       u1_R1_30, u1_R1_31, u1_R1_6, u1_R1_7, u1_R1_8, u1_R2_10, u1_R2_11, u1_R2_14, u1_R2_15, 
       u1_R2_18, u1_R2_19, u1_R2_22, u1_R2_23, u1_R2_26, u1_R2_27, u1_R2_3, u1_R2_30, u1_R2_31, 
       u1_R2_4, u1_R2_6, u1_R3_10, u1_R3_11, u1_R3_14, u1_R3_19, u1_R3_2, u1_R3_22, u1_R3_23, 
       u1_R3_26, u1_R3_27, u1_R3_3, u1_R3_30, u1_R3_31, u1_R3_6, u1_R3_7, u1_R4_10, u1_R4_11, 
       u1_R4_12, u1_R4_15, u1_R4_18, u1_R4_19, u1_R4_2, u1_R4_22, u1_R4_23, u1_R4_26, u1_R4_27, 
       u1_R4_30, u1_R4_31, u1_R5_10, u1_R5_11, u1_R5_14, u1_R5_15, u1_R5_19, u1_R5_2, u1_R5_22, 
       u1_R5_26, u1_R5_27, u1_R5_3, u1_R5_30, u1_R5_6, u1_R5_7, u1_R6_11, u1_R6_12, u1_R6_14, 
       u1_R6_15, u1_R6_18, u1_R6_19, u1_R6_22, u1_R6_23, u1_R6_26, u1_R6_27, u1_R6_3, u1_R6_30, 
       u1_R6_31, u1_R6_5, u1_R6_6, u1_R6_7, u1_R7_10, u1_R7_11, u1_R7_14, u1_R7_19, u1_R7_2, 
       u1_R7_21, u1_R7_22, u1_R7_23, u1_R7_26, u1_R7_27, u1_R7_3, u1_R7_30, u1_R7_31, u1_R8_10, 
       u1_R8_11, u1_R8_12, u1_R8_14, u1_R8_18, u1_R8_19, u1_R8_2, u1_R8_23, u1_R8_26, u1_R8_27, 
       u1_R8_3, u1_R8_30, u1_R8_31, u1_R8_7, u1_R9_10, u1_R9_11, u1_R9_13, u1_R9_14, u1_R9_17, 
       u1_R9_18, u1_R9_19, u1_R9_2, u1_R9_22, u1_R9_26, u1_R9_27, u1_R9_28, u1_R9_29, u1_R9_3, 
       u1_R9_30, u1_R9_31, u1_R9_32, u1_R9_5, u1_R9_6, u1_R9_7, u1_desIn_r_0, u1_desIn_r_1, u1_desIn_r_10, 
       u1_desIn_r_11, u1_desIn_r_12, u1_desIn_r_13, u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_16, u1_desIn_r_17, u1_desIn_r_18, u1_desIn_r_19, 
       u1_desIn_r_2, u1_desIn_r_20, u1_desIn_r_21, u1_desIn_r_22, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_26, u1_desIn_r_27, u1_desIn_r_28, 
       u1_desIn_r_3, u1_desIn_r_30, u1_desIn_r_31, u1_desIn_r_32, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_36, u1_desIn_r_38, 
       u1_desIn_r_4, u1_desIn_r_40, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_43, u1_desIn_r_44, u1_desIn_r_45, u1_desIn_r_46, u1_desIn_r_47, 
       u1_desIn_r_48, u1_desIn_r_49, u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_51, u1_desIn_r_52, u1_desIn_r_53, u1_desIn_r_54, u1_desIn_r_55, 
       u1_desIn_r_56, u1_desIn_r_58, u1_desIn_r_59, u1_desIn_r_6, u1_desIn_r_60, u1_desIn_r_61, u1_desIn_r_62, u1_desIn_r_63, u1_desIn_r_7, 
       u1_desIn_r_8, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_14, 
       u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, u1_key_r_2, u1_key_r_20, u1_key_r_21, u1_key_r_22, 
       u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, u1_key_r_28, u1_key_r_29, u1_key_r_3, u1_key_r_30, 
       u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, u1_key_r_36, u1_key_r_37, u1_key_r_38, u1_key_r_39, 
       u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, u1_key_r_44, u1_key_r_45, u1_key_r_46, u1_key_r_47, 
       u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, u1_key_r_52, u1_key_r_53, u1_key_r_54, u1_key_r_55, 
       u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_0, u1_uk_K_r0_1, u1_uk_K_r0_10, u1_uk_K_r0_11, u1_uk_K_r0_12, 
       u1_uk_K_r0_13, u1_uk_K_r0_14, u1_uk_K_r0_15, u1_uk_K_r0_16, u1_uk_K_r0_17, u1_uk_K_r0_18, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_20, 
       u1_uk_K_r0_21, u1_uk_K_r0_22, u1_uk_K_r0_23, u1_uk_K_r0_24, u1_uk_K_r0_25, u1_uk_K_r0_26, u1_uk_K_r0_27, u1_uk_K_r0_28, u1_uk_K_r0_29, 
       u1_uk_K_r0_3, u1_uk_K_r0_30, u1_uk_K_r0_31, u1_uk_K_r0_32, u1_uk_K_r0_33, u1_uk_K_r0_34, u1_uk_K_r0_35, u1_uk_K_r0_36, u1_uk_K_r0_37, 
       u1_uk_K_r0_38, u1_uk_K_r0_39, u1_uk_K_r0_4, u1_uk_K_r0_40, u1_uk_K_r0_41, u1_uk_K_r0_42, u1_uk_K_r0_43, u1_uk_K_r0_44, u1_uk_K_r0_45, 
       u1_uk_K_r0_46, u1_uk_K_r0_47, u1_uk_K_r0_48, u1_uk_K_r0_49, u1_uk_K_r0_5, u1_uk_K_r0_50, u1_uk_K_r0_51, u1_uk_K_r0_52, u1_uk_K_r0_53, 
       u1_uk_K_r0_54, u1_uk_K_r0_55, u1_uk_K_r0_6, u1_uk_K_r0_7, u1_uk_K_r0_8, u1_uk_K_r0_9, u1_uk_K_r10_0, u1_uk_K_r10_1, u1_uk_K_r10_10, 
       u1_uk_K_r10_11, u1_uk_K_r10_12, u1_uk_K_r10_13, u1_uk_K_r10_14, u1_uk_K_r10_15, u1_uk_K_r10_16, u1_uk_K_r10_17, u1_uk_K_r10_18, u1_uk_K_r10_19, 
       u1_uk_K_r10_2, u1_uk_K_r10_20, u1_uk_K_r10_21, u1_uk_K_r10_22, u1_uk_K_r10_23, u1_uk_K_r10_24, u1_uk_K_r10_25, u1_uk_K_r10_26, u1_uk_K_r10_27, 
       u1_uk_K_r10_28, u1_uk_K_r10_29, u1_uk_K_r10_3, u1_uk_K_r10_30, u1_uk_K_r10_31, u1_uk_K_r10_32, u1_uk_K_r10_33, u1_uk_K_r10_34, u1_uk_K_r10_35, 
       u1_uk_K_r10_36, u1_uk_K_r10_37, u1_uk_K_r10_38, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_40, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, 
       u1_uk_K_r10_44, u1_uk_K_r10_45, u1_uk_K_r10_46, u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r10_49, u1_uk_K_r10_5, u1_uk_K_r10_50, u1_uk_K_r10_51, 
       u1_uk_K_r10_52, u1_uk_K_r10_53, u1_uk_K_r10_54, u1_uk_K_r10_55, u1_uk_K_r10_6, u1_uk_K_r10_7, u1_uk_K_r10_8, u1_uk_K_r10_9, u1_uk_K_r11_0, 
       u1_uk_K_r11_1, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_12, u1_uk_K_r11_13, u1_uk_K_r11_14, u1_uk_K_r11_15, u1_uk_K_r11_16, u1_uk_K_r11_17, 
       u1_uk_K_r11_18, u1_uk_K_r11_19, u1_uk_K_r11_2, u1_uk_K_r11_20, u1_uk_K_r11_21, u1_uk_K_r11_22, u1_uk_K_r11_23, u1_uk_K_r11_24, u1_uk_K_r11_25, 
       u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_3, u1_uk_K_r11_30, u1_uk_K_r11_31, u1_uk_K_r11_32, u1_uk_K_r11_33, 
       u1_uk_K_r11_34, u1_uk_K_r11_35, u1_uk_K_r11_36, u1_uk_K_r11_37, u1_uk_K_r11_38, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_40, u1_uk_K_r11_41, 
       u1_uk_K_r11_42, u1_uk_K_r11_43, u1_uk_K_r11_44, u1_uk_K_r11_45, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_49, u1_uk_K_r11_5, 
       u1_uk_K_r11_50, u1_uk_K_r11_51, u1_uk_K_r11_52, u1_uk_K_r11_53, u1_uk_K_r11_54, u1_uk_K_r11_55, u1_uk_K_r11_6, u1_uk_K_r11_7, u1_uk_K_r11_8, 
       u1_uk_K_r11_9, u1_uk_K_r12_0, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_11, u1_uk_K_r12_12, u1_uk_K_r12_13, u1_uk_K_r12_14, u1_uk_K_r12_15, 
       u1_uk_K_r12_16, u1_uk_K_r12_17, u1_uk_K_r12_18, u1_uk_K_r12_19, u1_uk_K_r12_2, u1_uk_K_r12_20, u1_uk_K_r12_21, u1_uk_K_r12_22, u1_uk_K_r12_23, 
       u1_uk_K_r12_24, u1_uk_K_r12_25, u1_uk_K_r12_26, u1_uk_K_r12_27, u1_uk_K_r12_28, u1_uk_K_r12_29, u1_uk_K_r12_3, u1_uk_K_r12_30, u1_uk_K_r12_31, 
       u1_uk_K_r12_32, u1_uk_K_r12_33, u1_uk_K_r12_34, u1_uk_K_r12_35, u1_uk_K_r12_36, u1_uk_K_r12_37, u1_uk_K_r12_38, u1_uk_K_r12_39, u1_uk_K_r12_4, 
       u1_uk_K_r12_40, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_43, u1_uk_K_r12_44, u1_uk_K_r12_45, u1_uk_K_r12_46, u1_uk_K_r12_47, u1_uk_K_r12_48, 
       u1_uk_K_r12_49, u1_uk_K_r12_5, u1_uk_K_r12_50, u1_uk_K_r12_51, u1_uk_K_r12_52, u1_uk_K_r12_53, u1_uk_K_r12_54, u1_uk_K_r12_55, u1_uk_K_r12_6, 
       u1_uk_K_r12_7, u1_uk_K_r12_8, u1_uk_K_r12_9, u1_uk_K_r13_0, u1_uk_K_r13_1, u1_uk_K_r13_10, u1_uk_K_r13_11, u1_uk_K_r13_12, u1_uk_K_r13_13, 
       u1_uk_K_r13_14, u1_uk_K_r13_15, u1_uk_K_r13_16, u1_uk_K_r13_17, u1_uk_K_r13_18, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_20, u1_uk_K_r13_21, 
       u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_24, u1_uk_K_r13_25, u1_uk_K_r13_26, u1_uk_K_r13_27, u1_uk_K_r13_28, u1_uk_K_r13_29, u1_uk_K_r13_3, 
       u1_uk_K_r13_30, u1_uk_K_r13_31, u1_uk_K_r13_32, u1_uk_K_r13_33, u1_uk_K_r13_34, u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_37, u1_uk_K_r13_38, 
       u1_uk_K_r13_39, u1_uk_K_r13_4, u1_uk_K_r13_40, u1_uk_K_r13_41, u1_uk_K_r13_42, u1_uk_K_r13_43, u1_uk_K_r13_44, u1_uk_K_r13_45, u1_uk_K_r13_46, 
       u1_uk_K_r13_47, u1_uk_K_r13_48, u1_uk_K_r13_49, u1_uk_K_r13_5, u1_uk_K_r13_50, u1_uk_K_r13_51, u1_uk_K_r13_52, u1_uk_K_r13_53, u1_uk_K_r13_54, 
       u1_uk_K_r13_55, u1_uk_K_r13_6, u1_uk_K_r13_7, u1_uk_K_r13_8, u1_uk_K_r13_9, u1_uk_K_r14_10, u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_15, 
       u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, u1_uk_K_r14_39, u1_uk_K_r14_42, u1_uk_K_r14_43, 
       u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, u1_uk_K_r1_0, u1_uk_K_r1_1, u1_uk_K_r1_10, 
       u1_uk_K_r1_11, u1_uk_K_r1_12, u1_uk_K_r1_13, u1_uk_K_r1_14, u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_19, 
       u1_uk_K_r1_2, u1_uk_K_r1_20, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_23, u1_uk_K_r1_24, u1_uk_K_r1_25, u1_uk_K_r1_26, u1_uk_K_r1_27, 
       u1_uk_K_r1_28, u1_uk_K_r1_29, u1_uk_K_r1_3, u1_uk_K_r1_30, u1_uk_K_r1_31, u1_uk_K_r1_32, u1_uk_K_r1_33, u1_uk_K_r1_34, u1_uk_K_r1_35, 
       u1_uk_K_r1_36, u1_uk_K_r1_37, u1_uk_K_r1_38, u1_uk_K_r1_39, u1_uk_K_r1_4, u1_uk_K_r1_40, u1_uk_K_r1_41, u1_uk_K_r1_42, u1_uk_K_r1_43, 
       u1_uk_K_r1_44, u1_uk_K_r1_45, u1_uk_K_r1_46, u1_uk_K_r1_47, u1_uk_K_r1_48, u1_uk_K_r1_49, u1_uk_K_r1_5, u1_uk_K_r1_50, u1_uk_K_r1_51, 
       u1_uk_K_r1_52, u1_uk_K_r1_53, u1_uk_K_r1_54, u1_uk_K_r1_55, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r1_8, u1_uk_K_r1_9, u1_uk_K_r2_0, 
       u1_uk_K_r2_1, u1_uk_K_r2_10, u1_uk_K_r2_11, u1_uk_K_r2_12, u1_uk_K_r2_13, u1_uk_K_r2_14, u1_uk_K_r2_15, u1_uk_K_r2_16, u1_uk_K_r2_17, 
       u1_uk_K_r2_18, u1_uk_K_r2_19, u1_uk_K_r2_2, u1_uk_K_r2_20, u1_uk_K_r2_21, u1_uk_K_r2_22, u1_uk_K_r2_23, u1_uk_K_r2_24, u1_uk_K_r2_25, 
       u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_3, u1_uk_K_r2_30, u1_uk_K_r2_31, u1_uk_K_r2_32, u1_uk_K_r2_33, 
       u1_uk_K_r2_34, u1_uk_K_r2_35, u1_uk_K_r2_36, u1_uk_K_r2_37, u1_uk_K_r2_38, u1_uk_K_r2_39, u1_uk_K_r2_4, u1_uk_K_r2_40, u1_uk_K_r2_41, 
       u1_uk_K_r2_42, u1_uk_K_r2_43, u1_uk_K_r2_44, u1_uk_K_r2_45, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_48, u1_uk_K_r2_49, u1_uk_K_r2_5, 
       u1_uk_K_r2_50, u1_uk_K_r2_51, u1_uk_K_r2_52, u1_uk_K_r2_53, u1_uk_K_r2_54, u1_uk_K_r2_55, u1_uk_K_r2_6, u1_uk_K_r2_7, u1_uk_K_r2_8, 
       u1_uk_K_r2_9, u1_uk_K_r3_0, u1_uk_K_r3_1, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_12, u1_uk_K_r3_13, u1_uk_K_r3_14, u1_uk_K_r3_15, 
       u1_uk_K_r3_16, u1_uk_K_r3_17, u1_uk_K_r3_18, u1_uk_K_r3_19, u1_uk_K_r3_2, u1_uk_K_r3_20, u1_uk_K_r3_21, u1_uk_K_r3_22, u1_uk_K_r3_23, 
       u1_uk_K_r3_24, u1_uk_K_r3_25, u1_uk_K_r3_26, u1_uk_K_r3_27, u1_uk_K_r3_28, u1_uk_K_r3_29, u1_uk_K_r3_3, u1_uk_K_r3_30, u1_uk_K_r3_31, 
       u1_uk_K_r3_32, u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_36, u1_uk_K_r3_37, u1_uk_K_r3_38, u1_uk_K_r3_39, u1_uk_K_r3_4, 
       u1_uk_K_r3_40, u1_uk_K_r3_41, u1_uk_K_r3_42, u1_uk_K_r3_43, u1_uk_K_r3_44, u1_uk_K_r3_45, u1_uk_K_r3_46, u1_uk_K_r3_47, u1_uk_K_r3_48, 
       u1_uk_K_r3_49, u1_uk_K_r3_5, u1_uk_K_r3_50, u1_uk_K_r3_51, u1_uk_K_r3_52, u1_uk_K_r3_53, u1_uk_K_r3_54, u1_uk_K_r3_55, u1_uk_K_r3_6, 
       u1_uk_K_r3_7, u1_uk_K_r3_8, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_1, u1_uk_K_r4_10, u1_uk_K_r4_11, u1_uk_K_r4_12, u1_uk_K_r4_13, 
       u1_uk_K_r4_14, u1_uk_K_r4_15, u1_uk_K_r4_16, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_19, u1_uk_K_r4_2, u1_uk_K_r4_20, u1_uk_K_r4_21, 
       u1_uk_K_r4_22, u1_uk_K_r4_23, u1_uk_K_r4_24, u1_uk_K_r4_25, u1_uk_K_r4_26, u1_uk_K_r4_27, u1_uk_K_r4_28, u1_uk_K_r4_29, u1_uk_K_r4_3, 
       u1_uk_K_r4_30, u1_uk_K_r4_31, u1_uk_K_r4_32, u1_uk_K_r4_33, u1_uk_K_r4_34, u1_uk_K_r4_35, u1_uk_K_r4_36, u1_uk_K_r4_37, u1_uk_K_r4_38, 
       u1_uk_K_r4_39, u1_uk_K_r4_4, u1_uk_K_r4_40, u1_uk_K_r4_41, u1_uk_K_r4_42, u1_uk_K_r4_43, u1_uk_K_r4_44, u1_uk_K_r4_45, u1_uk_K_r4_46, 
       u1_uk_K_r4_47, u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_50, u1_uk_K_r4_51, u1_uk_K_r4_52, u1_uk_K_r4_53, u1_uk_K_r4_54, 
       u1_uk_K_r4_55, u1_uk_K_r4_6, u1_uk_K_r4_7, u1_uk_K_r4_8, u1_uk_K_r4_9, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_11, 
       u1_uk_K_r5_12, u1_uk_K_r5_13, u1_uk_K_r5_14, u1_uk_K_r5_15, u1_uk_K_r5_16, u1_uk_K_r5_17, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_2, 
       u1_uk_K_r5_20, u1_uk_K_r5_21, u1_uk_K_r5_22, u1_uk_K_r5_23, u1_uk_K_r5_24, u1_uk_K_r5_25, u1_uk_K_r5_26, u1_uk_K_r5_27, u1_uk_K_r5_28, 
       u1_uk_K_r5_29, u1_uk_K_r5_3, u1_uk_K_r5_30, u1_uk_K_r5_31, u1_uk_K_r5_32, u1_uk_K_r5_33, u1_uk_K_r5_34, u1_uk_K_r5_35, u1_uk_K_r5_36, 
       u1_uk_K_r5_37, u1_uk_K_r5_38, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_42, u1_uk_K_r5_43, u1_uk_K_r5_44, 
       u1_uk_K_r5_45, u1_uk_K_r5_46, u1_uk_K_r5_47, u1_uk_K_r5_48, u1_uk_K_r5_49, u1_uk_K_r5_5, u1_uk_K_r5_50, u1_uk_K_r5_51, u1_uk_K_r5_52, 
       u1_uk_K_r5_53, u1_uk_K_r5_54, u1_uk_K_r5_55, u1_uk_K_r5_6, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r5_9, u1_uk_K_r6_0, u1_uk_K_r6_1, 
       u1_uk_K_r6_10, u1_uk_K_r6_11, u1_uk_K_r6_12, u1_uk_K_r6_13, u1_uk_K_r6_14, u1_uk_K_r6_15, u1_uk_K_r6_16, u1_uk_K_r6_17, u1_uk_K_r6_18, 
       u1_uk_K_r6_19, u1_uk_K_r6_2, u1_uk_K_r6_20, u1_uk_K_r6_21, u1_uk_K_r6_22, u1_uk_K_r6_23, u1_uk_K_r6_24, u1_uk_K_r6_25, u1_uk_K_r6_26, 
       u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, u1_uk_K_r6_31, u1_uk_K_r6_32, u1_uk_K_r6_33, u1_uk_K_r6_34, 
       u1_uk_K_r6_35, u1_uk_K_r6_36, u1_uk_K_r6_37, u1_uk_K_r6_38, u1_uk_K_r6_39, u1_uk_K_r6_4, u1_uk_K_r6_40, u1_uk_K_r6_41, u1_uk_K_r6_42, 
       u1_uk_K_r6_43, u1_uk_K_r6_44, u1_uk_K_r6_45, u1_uk_K_r6_46, u1_uk_K_r6_47, u1_uk_K_r6_48, u1_uk_K_r6_49, u1_uk_K_r6_5, u1_uk_K_r6_50, 
       u1_uk_K_r6_51, u1_uk_K_r6_52, u1_uk_K_r6_53, u1_uk_K_r6_54, u1_uk_K_r6_55, u1_uk_K_r6_6, u1_uk_K_r6_7, u1_uk_K_r6_8, u1_uk_K_r6_9, 
       u1_uk_K_r7_0, u1_uk_K_r7_1, u1_uk_K_r7_10, u1_uk_K_r7_11, u1_uk_K_r7_12, u1_uk_K_r7_13, u1_uk_K_r7_14, u1_uk_K_r7_15, u1_uk_K_r7_16, 
       u1_uk_K_r7_17, u1_uk_K_r7_18, u1_uk_K_r7_19, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_21, u1_uk_K_r7_22, u1_uk_K_r7_23, u1_uk_K_r7_24, 
       u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_28, u1_uk_K_r7_29, u1_uk_K_r7_3, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, 
       u1_uk_K_r7_33, u1_uk_K_r7_34, u1_uk_K_r7_35, u1_uk_K_r7_36, u1_uk_K_r7_37, u1_uk_K_r7_38, u1_uk_K_r7_39, u1_uk_K_r7_4, u1_uk_K_r7_40, 
       u1_uk_K_r7_41, u1_uk_K_r7_42, u1_uk_K_r7_43, u1_uk_K_r7_44, u1_uk_K_r7_45, u1_uk_K_r7_46, u1_uk_K_r7_47, u1_uk_K_r7_48, u1_uk_K_r7_49, 
       u1_uk_K_r7_5, u1_uk_K_r7_50, u1_uk_K_r7_51, u1_uk_K_r7_52, u1_uk_K_r7_53, u1_uk_K_r7_54, u1_uk_K_r7_55, u1_uk_K_r7_6, u1_uk_K_r7_7, 
       u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_0, u1_uk_K_r8_1, u1_uk_K_r8_10, u1_uk_K_r8_11, u1_uk_K_r8_12, u1_uk_K_r8_13, u1_uk_K_r8_14, 
       u1_uk_K_r8_15, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_18, u1_uk_K_r8_19, u1_uk_K_r8_2, u1_uk_K_r8_20, u1_uk_K_r8_21, u1_uk_K_r8_22, 
       u1_uk_K_r8_23, u1_uk_K_r8_24, u1_uk_K_r8_25, u1_uk_K_r8_26, u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_29, u1_uk_K_r8_3, u1_uk_K_r8_30, 
       u1_uk_K_r8_31, u1_uk_K_r8_32, u1_uk_K_r8_33, u1_uk_K_r8_34, u1_uk_K_r8_35, u1_uk_K_r8_36, u1_uk_K_r8_37, u1_uk_K_r8_38, u1_uk_K_r8_39, 
       u1_uk_K_r8_4, u1_uk_K_r8_40, u1_uk_K_r8_41, u1_uk_K_r8_42, u1_uk_K_r8_43, u1_uk_K_r8_44, u1_uk_K_r8_45, u1_uk_K_r8_46, u1_uk_K_r8_47, 
       u1_uk_K_r8_48, u1_uk_K_r8_49, u1_uk_K_r8_5, u1_uk_K_r8_50, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_53, u1_uk_K_r8_54, u1_uk_K_r8_55, 
       u1_uk_K_r8_6, u1_uk_K_r8_7, u1_uk_K_r8_8, u1_uk_K_r8_9, u1_uk_K_r9_0, u1_uk_K_r9_1, u1_uk_K_r9_10, u1_uk_K_r9_11, u1_uk_K_r9_12, 
       u1_uk_K_r9_13, u1_uk_K_r9_14, u1_uk_K_r9_15, u1_uk_K_r9_16, u1_uk_K_r9_17, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_2, u1_uk_K_r9_20, 
       u1_uk_K_r9_21, u1_uk_K_r9_22, u1_uk_K_r9_23, u1_uk_K_r9_24, u1_uk_K_r9_25, u1_uk_K_r9_26, u1_uk_K_r9_27, u1_uk_K_r9_28, u1_uk_K_r9_29, 
       u1_uk_K_r9_3, u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_32, u1_uk_K_r9_33, u1_uk_K_r9_34, u1_uk_K_r9_35, u1_uk_K_r9_36, u1_uk_K_r9_37, 
       u1_uk_K_r9_38, u1_uk_K_r9_39, u1_uk_K_r9_4, u1_uk_K_r9_40, u1_uk_K_r9_41, u1_uk_K_r9_42, u1_uk_K_r9_43, u1_uk_K_r9_44, u1_uk_K_r9_45, 
       u1_uk_K_r9_46, u1_uk_K_r9_47, u1_uk_K_r9_48, u1_uk_K_r9_49, u1_uk_K_r9_5, u1_uk_K_r9_50, u1_uk_K_r9_51, u1_uk_K_r9_52, u1_uk_K_r9_53, 
       u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_8, u1_uk_K_r9_9, u1_uk_n10, u1_uk_n100, u1_uk_n1000, 
       u1_uk_n1001, u1_uk_n1004, u1_uk_n1005, u1_uk_n1006, u1_uk_n1007, u1_uk_n1008, u1_uk_n1009, u1_uk_n1010, u1_uk_n1011, 
       u1_uk_n1012, u1_uk_n1013, u1_uk_n1014, u1_uk_n1016, u1_uk_n1017, u1_uk_n1018, u1_uk_n1019, u1_uk_n102, u1_uk_n1020, 
       u1_uk_n1022, u1_uk_n1024, u1_uk_n1026, u1_uk_n1027, u1_uk_n1028, u1_uk_n1030, u1_uk_n1032, u1_uk_n1033, u1_uk_n1035, 
       u1_uk_n1036, u1_uk_n1037, u1_uk_n1039, u1_uk_n1040, u1_uk_n1041, u1_uk_n1042, u1_uk_n1043, u1_uk_n1044, u1_uk_n1045, 
       u1_uk_n1046, u1_uk_n1047, u1_uk_n1048, u1_uk_n1049, u1_uk_n1051, u1_uk_n1052, u1_uk_n1053, u1_uk_n1055, u1_uk_n1059, 
       u1_uk_n1062, u1_uk_n1064, u1_uk_n1066, u1_uk_n1067, u1_uk_n1068, u1_uk_n1069, u1_uk_n1071, u1_uk_n1072, u1_uk_n1075, 
       u1_uk_n1077, u1_uk_n1078, u1_uk_n1081, u1_uk_n1082, u1_uk_n1084, u1_uk_n1085, u1_uk_n1086, u1_uk_n1087, u1_uk_n1089, 
       u1_uk_n109, u1_uk_n1091, u1_uk_n1093, u1_uk_n1094, u1_uk_n1095, u1_uk_n1097, u1_uk_n1098, u1_uk_n1099, u1_uk_n11, 
       u1_uk_n110, u1_uk_n1100, u1_uk_n1102, u1_uk_n1103, u1_uk_n1107, u1_uk_n1108, u1_uk_n1110, u1_uk_n1111, u1_uk_n1112, 
       u1_uk_n1116, u1_uk_n1117, u1_uk_n1120, u1_uk_n1122, u1_uk_n1127, u1_uk_n1129, u1_uk_n1131, u1_uk_n1132, u1_uk_n1133, 
       u1_uk_n1135, u1_uk_n1136, u1_uk_n1137, u1_uk_n1139, u1_uk_n1141, u1_uk_n1142, u1_uk_n1144, u1_uk_n1145, u1_uk_n1146, 
       u1_uk_n1149, u1_uk_n1150, u1_uk_n1151, u1_uk_n1152, u1_uk_n1161, u1_uk_n1162, u1_uk_n1164, u1_uk_n1165, u1_uk_n1168, 
       u1_uk_n1169, u1_uk_n117, u1_uk_n1172, u1_uk_n1173, u1_uk_n1174, u1_uk_n1175, u1_uk_n1176, u1_uk_n1177, u1_uk_n1178, 
       u1_uk_n1179, u1_uk_n118, u1_uk_n1180, u1_uk_n1181, u1_uk_n1182, u1_uk_n1183, u1_uk_n1184, u1_uk_n1185, u1_uk_n1187, 
       u1_uk_n1188, u1_uk_n1189, u1_uk_n1190, u1_uk_n1191, u1_uk_n1192, u1_uk_n1195, u1_uk_n1197, u1_uk_n1198, u1_uk_n1201, 
       u1_uk_n1204, u1_uk_n1205, u1_uk_n1208, u1_uk_n1209, u1_uk_n1213, u1_uk_n1214, u1_uk_n1215, u1_uk_n1218, u1_uk_n1219, 
       u1_uk_n1220, u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1230, 
       u1_uk_n1231, u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, u1_uk_n1240, 
       u1_uk_n1241, u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, u1_uk_n1249, 
       u1_uk_n1250, u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, 
       u1_uk_n1260, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1268, 
       u1_uk_n1269, u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, u1_uk_n1277, 
       u1_uk_n1278, u1_uk_n1279, u1_uk_n128, u1_uk_n1281, u1_uk_n1282, u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, 
       u1_uk_n129, u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, 
       u1_uk_n1299, u1_uk_n1300, u1_uk_n1303, u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, 
       u1_uk_n1311, u1_uk_n1312, u1_uk_n1313, u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, 
       u1_uk_n1320, u1_uk_n1321, u1_uk_n1322, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, 
       u1_uk_n1329, u1_uk_n1330, u1_uk_n1331, u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, 
       u1_uk_n1339, u1_uk_n1340, u1_uk_n1341, u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, 
       u1_uk_n1348, u1_uk_n1349, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, 
       u1_uk_n1357, u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, 
       u1_uk_n1369, u1_uk_n1371, u1_uk_n1372, u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, 
       u1_uk_n1381, u1_uk_n1382, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, 
       u1_uk_n1395, u1_uk_n1396, u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, 
       u1_uk_n1404, u1_uk_n1405, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, u1_uk_n141, u1_uk_n1410, u1_uk_n1411, 
       u1_uk_n1412, u1_uk_n1413, u1_uk_n1414, u1_uk_n1415, u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, u1_uk_n142, u1_uk_n1422, 
       u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, u1_uk_n1426, u1_uk_n1427, u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, u1_uk_n1433, 
       u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, 
       u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, u1_uk_n1448, u1_uk_n1449, u1_uk_n145, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, 
       u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n146, u1_uk_n1460, u1_uk_n1461, 
       u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, u1_uk_n1468, u1_uk_n1469, u1_uk_n147, u1_uk_n1470, 
       u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, u1_uk_n1478, u1_uk_n148, u1_uk_n1482, 
       u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, u1_uk_n1490, u1_uk_n1491, 
       u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, u1_uk_n1501, u1_uk_n1504, 
       u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, u1_uk_n1518, u1_uk_n1520, 
       u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1530, u1_uk_n1531, 
       u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, u1_uk_n1541, u1_uk_n1543, 
       u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, u1_uk_n1548, u1_uk_n1549, u1_uk_n155, u1_uk_n1551, u1_uk_n1552, u1_uk_n1554, 
       u1_uk_n1555, u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, u1_uk_n1563, 
       u1_uk_n1564, u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, u1_uk_n1573, 
       u1_uk_n1574, u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, u1_uk_n1588, 
       u1_uk_n1592, u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, u1_uk_n1604, 
       u1_uk_n1605, u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, u1_uk_n161, u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, 
       u1_uk_n1615, u1_uk_n1616, u1_uk_n1618, u1_uk_n1619, u1_uk_n162, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, 
       u1_uk_n1624, u1_uk_n1625, u1_uk_n1626, u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, u1_uk_n163, u1_uk_n1630, u1_uk_n1632, 
       u1_uk_n1633, u1_uk_n1634, u1_uk_n1635, u1_uk_n1639, u1_uk_n164, u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, u1_uk_n1643, 
       u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, u1_uk_n1649, u1_uk_n1651, u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, u1_uk_n1655, 
       u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, u1_uk_n1661, u1_uk_n1662, u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, u1_uk_n1669, 
       u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, u1_uk_n1676, u1_uk_n1677, u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, 
       u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, u1_uk_n1690, u1_uk_n1691, u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, u1_uk_n1695, 
       u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, u1_uk_n17, u1_uk_n1702, u1_uk_n1703, u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, 
       u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, 
       u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, u1_uk_n1721, u1_uk_n1722, u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, 
       u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, 
       u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, u1_uk_n1750, u1_uk_n1751, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, 
       u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, u1_uk_n1761, u1_uk_n1762, u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, 
       u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, u1_uk_n1772, u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, 
       u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, u1_uk_n1783, u1_uk_n1784, u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, 
       u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, u1_uk_n1798, u1_uk_n1799, u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, 
       u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, 
       u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n182, u1_uk_n1820, 
       u1_uk_n1821, u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, u1_uk_n1827, u1_uk_n1829, u1_uk_n1830, u1_uk_n1831, 
       u1_uk_n1832, u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n1840, 
       u1_uk_n1841, u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, u1_uk_n1846, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, 
       u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, u1_uk_n1855, u1_uk_n1856, u1_uk_n1858, u1_uk_n1859, 
       u1_uk_n1860, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, u1_uk_n1866, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, 
       u1_uk_n187, u1_uk_n1870, u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, u1_uk_n1876, u1_uk_n1879, u1_uk_n188, 
       u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, u1_uk_n1887, u1_uk_n191, 
       u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, u1_uk_n209, u1_uk_n213, u1_uk_n214, u1_uk_n217, u1_uk_n220, 
       u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n231, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, 
       u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n291, u1_uk_n292, 
       u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n301, u1_uk_n305, u1_uk_n306, u1_uk_n308, u1_uk_n31, u1_uk_n313, 
       u1_uk_n319, u1_uk_n335, u1_uk_n338, u1_uk_n342, u1_uk_n346, u1_uk_n363, u1_uk_n373, u1_uk_n375, u1_uk_n377, 
       u1_uk_n391, u1_uk_n395, u1_uk_n408, u1_uk_n409, u1_uk_n415, u1_uk_n456, u1_uk_n460, u1_uk_n467, u1_uk_n468, 
       u1_uk_n472, u1_uk_n500, u1_uk_n501, u1_uk_n503, u1_uk_n518, u1_uk_n526, u1_uk_n551, u1_uk_n582, u1_uk_n586, 
       u1_uk_n587, u1_uk_n590, u1_uk_n60, u1_uk_n601, u1_uk_n603, u1_uk_n63, u1_uk_n634, u1_uk_n656, u1_uk_n662, 
       u1_uk_n665, u1_uk_n671, u1_uk_n681, u1_uk_n682, u1_uk_n686, u1_uk_n688, u1_uk_n689, u1_uk_n692, u1_uk_n694, 
       u1_uk_n695, u1_uk_n717, u1_uk_n83, u1_uk_n92, u1_uk_n93, u1_uk_n94, u1_uk_n945, u1_uk_n946, u1_uk_n947, 
       u1_uk_n951, u1_uk_n952, u1_uk_n953, u1_uk_n954, u1_uk_n956, u1_uk_n957, u1_uk_n958, u1_uk_n959, u1_uk_n960, 
       u1_uk_n961, u1_uk_n962, u1_uk_n963, u1_uk_n964, u1_uk_n965, u1_uk_n966, u1_uk_n967, u1_uk_n968, u1_uk_n971, 
       u1_uk_n972, u1_uk_n975, u1_uk_n977, u1_uk_n978, u1_uk_n979, u1_uk_n980, u1_uk_n981, u1_uk_n982, u1_uk_n983, 
       u1_uk_n984, u1_uk_n986, u1_uk_n987, u1_uk_n99, u1_uk_n990, u1_uk_n991, u1_uk_n992, u1_uk_n994, u1_uk_n995, 
       u1_uk_n996, u1_uk_n997, u1_uk_n998, u1_uk_n999, u2_FP_1, u2_FP_10, u2_FP_11, u2_FP_12, u2_FP_13, 
       u2_FP_14, u2_FP_15, u2_FP_16, u2_FP_17, u2_FP_18, u2_FP_19, u2_FP_2, u2_FP_20, u2_FP_21, 
       u2_FP_22, u2_FP_23, u2_FP_24, u2_FP_25, u2_FP_26, u2_FP_27, u2_FP_28, u2_FP_29, u2_FP_3, 
       u2_FP_30, u2_FP_31, u2_FP_32, u2_FP_34, u2_FP_35, u2_FP_38, u2_FP_39, u2_FP_4, u2_FP_42, 
       u2_FP_43, u2_FP_46, u2_FP_47, u2_FP_5, u2_FP_50, u2_FP_51, u2_FP_54, u2_FP_58, u2_FP_59, 
       u2_FP_6, u2_FP_62, u2_FP_63, u2_FP_7, u2_FP_8, u2_FP_9, u2_K10_10, u2_K10_15, u2_K10_16, 
       u2_K10_21, u2_K10_27, u2_K10_28, u2_K10_29, u2_K10_3, u2_K10_30, u2_K10_32, u2_K10_34, u2_K10_4, 
       u2_K10_45, u2_K10_46, u2_K10_6, u2_K11_1, u2_K11_10, u2_K11_15, u2_K11_16, u2_K11_18, u2_K11_2, 
       u2_K11_21, u2_K11_22, u2_K11_23, u2_K11_25, u2_K11_27, u2_K11_28, u2_K11_3, u2_K11_30, u2_K11_32, 
       u2_K11_33, u2_K11_34, u2_K11_35, u2_K11_36, u2_K11_37, u2_K11_38, u2_K11_39, u2_K11_4, u2_K11_40, 
       u2_K11_41, u2_K11_42, u2_K11_43, u2_K11_44, u2_K11_45, u2_K11_46, u2_K11_48, u2_K11_5, u2_K11_6, 
       u2_K11_7, u2_K11_8, u2_K11_9, u2_K12_15, u2_K12_16, u2_K12_21, u2_K12_22, u2_K12_24, u2_K12_26, 
       u2_K12_27, u2_K12_28, u2_K12_29, u2_K12_3, u2_K12_31, u2_K12_33, u2_K12_34, u2_K12_35, u2_K12_37, 
       u2_K12_39, u2_K12_40, u2_K12_41, u2_K12_43, u2_K12_45, u2_K12_46, u2_K12_6, u2_K12_8, u2_K12_9, 
       u2_K13_1, u2_K13_10, u2_K13_11, u2_K13_12, u2_K13_13, u2_K13_14, u2_K13_15, u2_K13_16, u2_K13_17, 
       u2_K13_18, u2_K13_19, u2_K13_20, u2_K13_21, u2_K13_22, u2_K13_23, u2_K13_24, u2_K13_25, u2_K13_26, 
       u2_K13_27, u2_K13_28, u2_K13_29, u2_K13_3, u2_K13_31, u2_K13_33, u2_K13_34, u2_K13_36, u2_K13_38, 
       u2_K13_39, u2_K13_4, u2_K13_40, u2_K13_41, u2_K13_42, u2_K13_43, u2_K13_44, u2_K13_45, u2_K13_46, 
       u2_K13_47, u2_K13_6, u2_K13_8, u2_K13_9, u2_K14_1, u2_K14_10, u2_K14_11, u2_K14_12, u2_K14_13, 
       u2_K14_14, u2_K14_15, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_19, u2_K14_2, u2_K14_20, u2_K14_21, 
       u2_K14_22, u2_K14_23, u2_K14_24, u2_K14_25, u2_K14_26, u2_K14_27, u2_K14_28, u2_K14_3, u2_K14_34, 
       u2_K14_35, u2_K14_37, u2_K14_39, u2_K14_4, u2_K14_40, u2_K14_41, u2_K14_42, u2_K14_43, u2_K14_44, 
       u2_K14_45, u2_K14_46, u2_K14_47, u2_K14_48, u2_K14_5, u2_K14_6, u2_K14_7, u2_K14_8, u2_K14_9, 
       u2_K15_10, u2_K15_11, u2_K15_13, u2_K15_15, u2_K15_16, u2_K15_18, u2_K15_20, u2_K15_21, u2_K15_22, 
       u2_K15_27, u2_K15_28, u2_K15_3, u2_K15_30, u2_K15_32, u2_K15_34, u2_K15_39, u2_K15_4, u2_K15_41, 
       u2_K15_43, u2_K15_45, u2_K15_46, u2_K15_5, u2_K15_7, u2_K15_9, u2_K16_10, u2_K16_15, u2_K16_16, 
       u2_K16_21, u2_K16_22, u2_K16_27, u2_K16_28, u2_K16_3, u2_K16_33, u2_K16_39, u2_K16_4, u2_K16_40, 
       u2_K16_45, u2_K16_46, u2_K16_9, u2_K1_1, u2_K1_10, u2_K1_11, u2_K1_12, u2_K1_13, u2_K1_14, 
       u2_K1_15, u2_K1_16, u2_K1_17, u2_K1_18, u2_K1_19, u2_K1_2, u2_K1_20, u2_K1_21, u2_K1_22, 
       u2_K1_23, u2_K1_24, u2_K1_25, u2_K1_26, u2_K1_27, u2_K1_28, u2_K1_3, u2_K1_30, u2_K1_32, 
       u2_K1_33, u2_K1_34, u2_K1_35, u2_K1_37, u2_K1_39, u2_K1_4, u2_K1_40, u2_K1_45, u2_K1_46, 
       u2_K1_48, u2_K1_5, u2_K1_6, u2_K1_7, u2_K1_8, u2_K1_9, u2_K2_15, u2_K2_16, u2_K2_21, 
       u2_K2_22, u2_K2_27, u2_K2_3, u2_K2_33, u2_K2_34, u2_K2_39, u2_K2_4, u2_K2_40, u2_K2_41, 
       u2_K2_43, u2_K2_45, u2_K2_46, u2_K2_9, u2_K3_15, u2_K3_16, u2_K3_27, u2_K3_28, u2_K3_29, 
       u2_K3_30, u2_K3_31, u2_K3_32, u2_K3_33, u2_K3_34, u2_K3_35, u2_K3_37, u2_K3_39, u2_K3_5, 
       u2_K3_7, u2_K4_21, u2_K4_22, u2_K4_27, u2_K4_33, u2_K4_34, u2_K4_35, u2_K4_37, u2_K4_38, 
       u2_K4_39, u2_K4_40, u2_K4_41, u2_K4_42, u2_K4_43, u2_K4_44, u2_K4_45, u2_K4_46, u2_K5_1, 
       u2_K5_10, u2_K5_15, u2_K5_16, u2_K5_21, u2_K5_22, u2_K5_28, u2_K5_3, u2_K5_34, u2_K5_39, 
       u2_K5_4, u2_K5_40, u2_K5_46, u2_K5_47, u2_K5_9, u2_K6_10, u2_K6_15, u2_K6_16, u2_K6_22, 
       u2_K6_23, u2_K6_25, u2_K6_27, u2_K6_28, u2_K6_29, u2_K6_3, u2_K6_31, u2_K6_34, u2_K6_36, 
       u2_K6_38, u2_K6_39, u2_K6_4, u2_K6_40, u2_K6_45, u2_K7_10, u2_K7_22, u2_K7_27, u2_K7_28, 
       u2_K7_3, u2_K7_33, u2_K7_4, u2_K7_40, u2_K7_45, u2_K7_46, u2_K7_9, u2_K8_10, u2_K8_15, 
       u2_K8_16, u2_K8_21, u2_K8_22, u2_K8_23, u2_K8_24, u2_K8_25, u2_K8_26, u2_K8_27, u2_K8_28, 
       u2_K8_29, u2_K8_30, u2_K8_31, u2_K8_32, u2_K8_33, u2_K8_34, u2_K8_35, u2_K8_36, u2_K8_37, 
       u2_K8_38, u2_K8_39, u2_K8_4, u2_K8_40, u2_K8_41, u2_K8_42, u2_K8_44, u2_K8_45, u2_K8_46, 
       u2_K8_9, u2_K9_1, u2_K9_15, u2_K9_27, u2_K9_28, u2_K9_29, u2_K9_3, u2_K9_30, u2_K9_31, 
       u2_K9_32, u2_K9_34, u2_K9_39, u2_K9_40, u2_K9_45, u2_K9_46, u2_K9_47, u2_L0_1, u2_L0_10, 
       u2_L0_11, u2_L0_12, u2_L0_13, u2_L0_14, u2_L0_15, u2_L0_16, u2_L0_17, u2_L0_18, u2_L0_19, 
       u2_L0_2, u2_L0_20, u2_L0_21, u2_L0_22, u2_L0_23, u2_L0_24, u2_L0_25, u2_L0_26, u2_L0_27, 
       u2_L0_28, u2_L0_29, u2_L0_3, u2_L0_30, u2_L0_31, u2_L0_32, u2_L0_4, u2_L0_5, u2_L0_6, 
       u2_L0_7, u2_L0_8, u2_L0_9, u2_L10_1, u2_L10_10, u2_L10_11, u2_L10_12, u2_L10_13, u2_L10_14, 
       u2_L10_15, u2_L10_16, u2_L10_17, u2_L10_18, u2_L10_19, u2_L10_2, u2_L10_20, u2_L10_21, u2_L10_22, 
       u2_L10_23, u2_L10_24, u2_L10_25, u2_L10_26, u2_L10_27, u2_L10_28, u2_L10_29, u2_L10_3, u2_L10_30, 
       u2_L10_31, u2_L10_32, u2_L10_4, u2_L10_5, u2_L10_6, u2_L10_7, u2_L10_8, u2_L10_9, u2_L11_1, 
       u2_L11_10, u2_L11_11, u2_L11_12, u2_L11_13, u2_L11_14, u2_L11_15, u2_L11_16, u2_L11_17, u2_L11_18, 
       u2_L11_19, u2_L11_2, u2_L11_20, u2_L11_21, u2_L11_22, u2_L11_23, u2_L11_24, u2_L11_25, u2_L11_26, 
       u2_L11_27, u2_L11_28, u2_L11_29, u2_L11_3, u2_L11_30, u2_L11_31, u2_L11_32, u2_L11_4, u2_L11_5, 
       u2_L11_6, u2_L11_7, u2_L11_8, u2_L11_9, u2_L12_1, u2_L12_10, u2_L12_11, u2_L12_12, u2_L12_13, 
       u2_L12_14, u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_19, u2_L12_2, u2_L12_20, u2_L12_21, 
       u2_L12_22, u2_L12_23, u2_L12_24, u2_L12_25, u2_L12_26, u2_L12_27, u2_L12_28, u2_L12_29, u2_L12_3, 
       u2_L12_30, u2_L12_31, u2_L12_32, u2_L12_4, u2_L12_5, u2_L12_6, u2_L12_7, u2_L12_8, u2_L12_9, 
       u2_L13_1, u2_L13_10, u2_L13_11, u2_L13_12, u2_L13_13, u2_L13_14, u2_L13_15, u2_L13_16, u2_L13_17, 
       u2_L13_18, u2_L13_19, u2_L13_2, u2_L13_20, u2_L13_21, u2_L13_22, u2_L13_23, u2_L13_24, u2_L13_25, 
       u2_L13_26, u2_L13_27, u2_L13_28, u2_L13_29, u2_L13_3, u2_L13_30, u2_L13_31, u2_L13_32, u2_L13_4, 
       u2_L13_5, u2_L13_6, u2_L13_7, u2_L13_8, u2_L13_9, u2_L14_1, u2_L14_10, u2_L14_11, u2_L14_12, 
       u2_L14_13, u2_L14_14, u2_L14_15, u2_L14_16, u2_L14_17, u2_L14_18, u2_L14_19, u2_L14_2, u2_L14_20, 
       u2_L14_21, u2_L14_22, u2_L14_23, u2_L14_24, u2_L14_25, u2_L14_26, u2_L14_27, u2_L14_28, u2_L14_29, 
       u2_L14_3, u2_L14_30, u2_L14_31, u2_L14_32, u2_L14_4, u2_L14_5, u2_L14_6, u2_L14_7, u2_L14_8, 
       u2_L14_9, u2_L1_1, u2_L1_10, u2_L1_11, u2_L1_12, u2_L1_13, u2_L1_14, u2_L1_15, u2_L1_16, 
       u2_L1_17, u2_L1_18, u2_L1_19, u2_L1_2, u2_L1_20, u2_L1_21, u2_L1_22, u2_L1_23, u2_L1_24, 
       u2_L1_25, u2_L1_26, u2_L1_27, u2_L1_28, u2_L1_29, u2_L1_3, u2_L1_30, u2_L1_31, u2_L1_32, 
       u2_L1_4, u2_L1_5, u2_L1_6, u2_L1_7, u2_L1_8, u2_L1_9, u2_L2_1, u2_L2_10, u2_L2_11, 
       u2_L2_12, u2_L2_13, u2_L2_14, u2_L2_15, u2_L2_16, u2_L2_17, u2_L2_18, u2_L2_19, u2_L2_2, 
       u2_L2_20, u2_L2_21, u2_L2_22, u2_L2_23, u2_L2_24, u2_L2_25, u2_L2_26, u2_L2_27, u2_L2_28, 
       u2_L2_29, u2_L2_3, u2_L2_30, u2_L2_31, u2_L2_32, u2_L2_4, u2_L2_5, u2_L2_6, u2_L2_7, 
       u2_L2_8, u2_L2_9, u2_L3_1, u2_L3_10, u2_L3_11, u2_L3_12, u2_L3_13, u2_L3_14, u2_L3_15, 
       u2_L3_16, u2_L3_17, u2_L3_18, u2_L3_19, u2_L3_2, u2_L3_20, u2_L3_21, u2_L3_22, u2_L3_23, 
       u2_L3_24, u2_L3_25, u2_L3_26, u2_L3_27, u2_L3_28, u2_L3_29, u2_L3_3, u2_L3_30, u2_L3_31, 
       u2_L3_32, u2_L3_4, u2_L3_5, u2_L3_6, u2_L3_7, u2_L3_8, u2_L3_9, u2_L4_1, u2_L4_10, 
       u2_L4_11, u2_L4_12, u2_L4_13, u2_L4_14, u2_L4_15, u2_L4_16, u2_L4_17, u2_L4_18, u2_L4_19, 
       u2_L4_2, u2_L4_20, u2_L4_21, u2_L4_22, u2_L4_23, u2_L4_24, u2_L4_25, u2_L4_26, u2_L4_27, 
       u2_L4_28, u2_L4_29, u2_L4_3, u2_L4_30, u2_L4_31, u2_L4_32, u2_L4_4, u2_L4_5, u2_L4_6, 
       u2_L4_7, u2_L4_8, u2_L4_9, u2_L5_1, u2_L5_10, u2_L5_11, u2_L5_12, u2_L5_13, u2_L5_14, 
       u2_L5_15, u2_L5_16, u2_L5_17, u2_L5_18, u2_L5_19, u2_L5_2, u2_L5_20, u2_L5_21, u2_L5_22, 
       u2_L5_23, u2_L5_24, u2_L5_25, u2_L5_26, u2_L5_27, u2_L5_28, u2_L5_29, u2_L5_3, u2_L5_30, 
       u2_L5_31, u2_L5_32, u2_L5_4, u2_L5_5, u2_L5_6, u2_L5_7, u2_L5_8, u2_L5_9, u2_L6_1, 
       u2_L6_10, u2_L6_11, u2_L6_12, u2_L6_13, u2_L6_14, u2_L6_15, u2_L6_16, u2_L6_17, u2_L6_18, 
       u2_L6_19, u2_L6_2, u2_L6_20, u2_L6_21, u2_L6_22, u2_L6_23, u2_L6_24, u2_L6_25, u2_L6_26, 
       u2_L6_27, u2_L6_28, u2_L6_29, u2_L6_3, u2_L6_30, u2_L6_31, u2_L6_32, u2_L6_4, u2_L6_5, 
       u2_L6_6, u2_L6_7, u2_L6_8, u2_L6_9, u2_L7_1, u2_L7_10, u2_L7_11, u2_L7_12, u2_L7_13, 
       u2_L7_14, u2_L7_15, u2_L7_16, u2_L7_17, u2_L7_18, u2_L7_19, u2_L7_2, u2_L7_20, u2_L7_21, 
       u2_L7_22, u2_L7_23, u2_L7_24, u2_L7_25, u2_L7_26, u2_L7_27, u2_L7_28, u2_L7_29, u2_L7_3, 
       u2_L7_30, u2_L7_31, u2_L7_32, u2_L7_4, u2_L7_5, u2_L7_6, u2_L7_7, u2_L7_8, u2_L7_9, 
       u2_L8_1, u2_L8_10, u2_L8_11, u2_L8_12, u2_L8_13, u2_L8_14, u2_L8_15, u2_L8_16, u2_L8_17, 
       u2_L8_18, u2_L8_19, u2_L8_2, u2_L8_20, u2_L8_21, u2_L8_22, u2_L8_23, u2_L8_24, u2_L8_25, 
       u2_L8_26, u2_L8_27, u2_L8_28, u2_L8_29, u2_L8_3, u2_L8_30, u2_L8_31, u2_L8_32, u2_L8_4, 
       u2_L8_5, u2_L8_6, u2_L8_7, u2_L8_8, u2_L8_9, u2_L9_1, u2_L9_10, u2_L9_11, u2_L9_12, 
       u2_L9_13, u2_L9_14, u2_L9_15, u2_L9_16, u2_L9_17, u2_L9_18, u2_L9_19, u2_L9_2, u2_L9_20, 
       u2_L9_21, u2_L9_22, u2_L9_23, u2_L9_24, u2_L9_25, u2_L9_26, u2_L9_27, u2_L9_28, u2_L9_29, 
       u2_L9_3, u2_L9_30, u2_L9_31, u2_L9_32, u2_L9_4, u2_L9_5, u2_L9_6, u2_L9_7, u2_L9_8, 
       u2_L9_9, u2_N0, u2_N1, u2_N10, u2_N100, u2_N101, u2_N102, u2_N103, u2_N104, 
       u2_N105, u2_N106, u2_N107, u2_N108, u2_N109, u2_N11, u2_N110, u2_N111, u2_N112, 
       u2_N113, u2_N114, u2_N115, u2_N116, u2_N117, u2_N118, u2_N119, u2_N12, u2_N120, 
       u2_N121, u2_N122, u2_N123, u2_N124, u2_N125, u2_N126, u2_N127, u2_N128, u2_N129, 
       u2_N13, u2_N130, u2_N131, u2_N132, u2_N133, u2_N134, u2_N135, u2_N136, u2_N137, 
       u2_N138, u2_N139, u2_N14, u2_N140, u2_N141, u2_N142, u2_N143, u2_N144, u2_N145, 
       u2_N146, u2_N147, u2_N148, u2_N149, u2_N15, u2_N150, u2_N151, u2_N152, u2_N153, 
       u2_N154, u2_N155, u2_N156, u2_N157, u2_N158, u2_N159, u2_N16, u2_N160, u2_N161, 
       u2_N162, u2_N163, u2_N164, u2_N165, u2_N166, u2_N167, u2_N168, u2_N169, u2_N17, 
       u2_N170, u2_N171, u2_N172, u2_N173, u2_N174, u2_N175, u2_N176, u2_N177, u2_N178, 
       u2_N179, u2_N18, u2_N180, u2_N181, u2_N182, u2_N183, u2_N184, u2_N185, u2_N186, 
       u2_N187, u2_N188, u2_N189, u2_N19, u2_N190, u2_N191, u2_N192, u2_N193, u2_N194, 
       u2_N195, u2_N196, u2_N197, u2_N198, u2_N199, u2_N2, u2_N20, u2_N200, u2_N201, 
       u2_N202, u2_N203, u2_N204, u2_N205, u2_N206, u2_N207, u2_N208, u2_N209, u2_N21, 
       u2_N210, u2_N211, u2_N212, u2_N213, u2_N214, u2_N215, u2_N216, u2_N217, u2_N218, 
       u2_N219, u2_N22, u2_N220, u2_N221, u2_N222, u2_N223, u2_N224, u2_N225, u2_N226, 
       u2_N227, u2_N228, u2_N229, u2_N23, u2_N230, u2_N231, u2_N232, u2_N233, u2_N234, 
       u2_N235, u2_N236, u2_N237, u2_N238, u2_N239, u2_N24, u2_N240, u2_N241, u2_N242, 
       u2_N243, u2_N244, u2_N245, u2_N246, u2_N247, u2_N248, u2_N249, u2_N25, u2_N250, 
       u2_N251, u2_N252, u2_N253, u2_N254, u2_N255, u2_N256, u2_N257, u2_N258, u2_N259, 
       u2_N26, u2_N260, u2_N261, u2_N262, u2_N263, u2_N264, u2_N265, u2_N266, u2_N267, 
       u2_N268, u2_N269, u2_N27, u2_N270, u2_N271, u2_N272, u2_N273, u2_N274, u2_N275, 
       u2_N276, u2_N277, u2_N278, u2_N279, u2_N28, u2_N280, u2_N281, u2_N282, u2_N283, 
       u2_N284, u2_N285, u2_N286, u2_N287, u2_N288, u2_N289, u2_N29, u2_N290, u2_N291, 
       u2_N292, u2_N293, u2_N294, u2_N295, u2_N296, u2_N297, u2_N298, u2_N299, u2_N3, 
       u2_N30, u2_N300, u2_N301, u2_N302, u2_N303, u2_N304, u2_N305, u2_N306, u2_N307, 
       u2_N308, u2_N309, u2_N31, u2_N310, u2_N311, u2_N312, u2_N313, u2_N314, u2_N315, 
       u2_N316, u2_N317, u2_N318, u2_N319, u2_N32, u2_N320, u2_N321, u2_N322, u2_N323, 
       u2_N324, u2_N325, u2_N326, u2_N327, u2_N328, u2_N329, u2_N33, u2_N330, u2_N331, 
       u2_N332, u2_N333, u2_N334, u2_N335, u2_N336, u2_N337, u2_N338, u2_N339, u2_N34, 
       u2_N340, u2_N341, u2_N342, u2_N343, u2_N344, u2_N345, u2_N346, u2_N347, u2_N348, 
       u2_N349, u2_N35, u2_N350, u2_N351, u2_N352, u2_N353, u2_N354, u2_N355, u2_N356, 
       u2_N357, u2_N358, u2_N359, u2_N36, u2_N360, u2_N361, u2_N362, u2_N363, u2_N364, 
       u2_N365, u2_N366, u2_N367, u2_N368, u2_N369, u2_N37, u2_N370, u2_N371, u2_N372, 
       u2_N373, u2_N374, u2_N375, u2_N376, u2_N377, u2_N378, u2_N379, u2_N38, u2_N380, 
       u2_N381, u2_N382, u2_N383, u2_N384, u2_N385, u2_N386, u2_N387, u2_N388, u2_N389, 
       u2_N39, u2_N390, u2_N391, u2_N392, u2_N393, u2_N394, u2_N395, u2_N396, u2_N397, 
       u2_N398, u2_N399, u2_N4, u2_N40, u2_N400, u2_N401, u2_N402, u2_N403, u2_N404, 
       u2_N405, u2_N406, u2_N407, u2_N408, u2_N409, u2_N41, u2_N410, u2_N411, u2_N412, 
       u2_N413, u2_N414, u2_N415, u2_N416, u2_N417, u2_N418, u2_N419, u2_N42, u2_N420, 
       u2_N421, u2_N422, u2_N423, u2_N424, u2_N425, u2_N426, u2_N427, u2_N428, u2_N429, 
       u2_N43, u2_N430, u2_N431, u2_N432, u2_N433, u2_N434, u2_N435, u2_N436, u2_N437, 
       u2_N438, u2_N439, u2_N44, u2_N440, u2_N441, u2_N442, u2_N443, u2_N444, u2_N445, 
       u2_N446, u2_N447, u2_N448, u2_N449, u2_N45, u2_N450, u2_N451, u2_N452, u2_N453, 
       u2_N454, u2_N455, u2_N456, u2_N457, u2_N458, u2_N459, u2_N46, u2_N460, u2_N461, 
       u2_N462, u2_N463, u2_N464, u2_N465, u2_N466, u2_N467, u2_N468, u2_N469, u2_N47, 
       u2_N470, u2_N471, u2_N472, u2_N473, u2_N474, u2_N475, u2_N476, u2_N477, u2_N478, 
       u2_N479, u2_N48, u2_N49, u2_N5, u2_N50, u2_N51, u2_N52, u2_N53, u2_N54, 
       u2_N55, u2_N56, u2_N57, u2_N58, u2_N59, u2_N6, u2_N60, u2_N61, u2_N62, 
       u2_N63, u2_N64, u2_N65, u2_N66, u2_N67, u2_N68, u2_N69, u2_N7, u2_N70, 
       u2_N71, u2_N72, u2_N73, u2_N74, u2_N75, u2_N76, u2_N77, u2_N78, u2_N79, 
       u2_N8, u2_N80, u2_N81, u2_N82, u2_N83, u2_N84, u2_N85, u2_N86, u2_N87, 
       u2_N88, u2_N89, u2_N9, u2_N90, u2_N91, u2_N92, u2_N93, u2_N94, u2_N95, 
       u2_N96, u2_N97, u2_N98, u2_N99, u2_R0_10, u2_R0_11, u2_R0_14, u2_R0_15, u2_R0_18, 
       u2_R0_2, u2_R0_22, u2_R0_23, u2_R0_26, u2_R0_27, u2_R0_28, u2_R0_3, u2_R0_30, u2_R0_31, 
       u2_R0_6, u2_R10_10, u2_R10_11, u2_R10_14, u2_R10_15, u2_R10_17, u2_R10_18, u2_R10_19, u2_R10_2, 
       u2_R10_20, u2_R10_22, u2_R10_23, u2_R10_24, u2_R10_26, u2_R10_27, u2_R10_28, u2_R10_30, u2_R10_31, 
       u2_R10_5, u2_R10_6, u2_R11_10, u2_R11_11, u2_R11_12, u2_R11_13, u2_R11_14, u2_R11_15, u2_R11_16, 
       u2_R11_17, u2_R11_18, u2_R11_19, u2_R11_2, u2_R11_20, u2_R11_22, u2_R11_23, u2_R11_25, u2_R11_26, 
       u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_3, u2_R11_30, u2_R11_31, u2_R11_32, u2_R11_5, u2_R11_6, 
       u2_R11_7, u2_R11_8, u2_R11_9, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_14, 
       u2_R12_15, u2_R12_16, u2_R12_17, u2_R12_18, u2_R12_19, u2_R12_2, u2_R12_23, u2_R12_24, u2_R12_26, 
       u2_R12_27, u2_R12_28, u2_R12_29, u2_R12_3, u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, 
       u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, u2_R13_10, u2_R13_11, u2_R13_13, u2_R13_14, u2_R13_15, 
       u2_R13_18, u2_R13_19, u2_R13_2, u2_R13_21, u2_R13_23, u2_R13_26, u2_R13_28, u2_R13_3, u2_R13_30, 
       u2_R13_31, u2_R13_4, u2_R13_6, u2_R13_7, u2_R13_8, u2_R1_10, u2_R1_11, u2_R1_18, u2_R1_19, 
       u2_R1_20, u2_R1_21, u2_R1_22, u2_R1_23, u2_R1_24, u2_R1_26, u2_R1_4, u2_R2_14, u2_R2_15, 
       u2_R2_18, u2_R2_22, u2_R2_23, u2_R2_24, u2_R2_26, u2_R2_27, u2_R2_28, u2_R2_29, u2_R2_30, 
       u2_R2_31, u2_R3_10, u2_R3_11, u2_R3_14, u2_R3_15, u2_R3_19, u2_R3_2, u2_R3_23, u2_R3_26, 
       u2_R3_27, u2_R3_3, u2_R3_31, u2_R3_32, u2_R3_6, u2_R3_7, u2_R4_10, u2_R4_11, u2_R4_15, 
       u2_R4_16, u2_R4_18, u2_R4_19, u2_R4_2, u2_R4_20, u2_R4_23, u2_R4_25, u2_R4_26, u2_R4_27, 
       u2_R4_3, u2_R4_30, u2_R4_7, u2_R5_15, u2_R5_18, u2_R5_19, u2_R5_2, u2_R5_22, u2_R5_27, 
       u2_R5_3, u2_R5_30, u2_R5_31, u2_R5_6, u2_R5_7, u2_R6_10, u2_R6_11, u2_R6_14, u2_R6_15, 
       u2_R6_16, u2_R6_17, u2_R6_18, u2_R6_19, u2_R6_20, u2_R6_21, u2_R6_22, u2_R6_23, u2_R6_24, 
       u2_R6_25, u2_R6_26, u2_R6_27, u2_R6_29, u2_R6_3, u2_R6_30, u2_R6_31, u2_R6_6, u2_R6_7, 
       u2_R7_10, u2_R7_18, u2_R7_19, u2_R7_2, u2_R7_20, u2_R7_21, u2_R7_23, u2_R7_26, u2_R7_27, 
       u2_R7_30, u2_R7_31, u2_R7_32, u2_R8_10, u2_R8_11, u2_R8_14, u2_R8_18, u2_R8_19, u2_R8_2, 
       u2_R8_21, u2_R8_23, u2_R8_3, u2_R8_30, u2_R8_31, u2_R8_7, u2_R9_1, u2_R9_10, u2_R9_11, 
       u2_R9_14, u2_R9_15, u2_R9_16, u2_R9_18, u2_R9_19, u2_R9_2, u2_R9_21, u2_R9_22, u2_R9_23, 
       u2_R9_24, u2_R9_25, u2_R9_26, u2_R9_27, u2_R9_28, u2_R9_29, u2_R9_3, u2_R9_30, u2_R9_31, 
       u2_R9_4, u2_R9_5, u2_R9_6, u2_R9_7, u2_desIn_r_0, u2_desIn_r_10, u2_desIn_r_11, u2_desIn_r_12, u2_desIn_r_13, 
       u2_desIn_r_14, u2_desIn_r_15, u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, u2_desIn_r_19, u2_desIn_r_2, u2_desIn_r_20, u2_desIn_r_21, 
       u2_desIn_r_22, u2_desIn_r_23, u2_desIn_r_24, u2_desIn_r_26, u2_desIn_r_28, u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_31, 
       u2_desIn_r_32, u2_desIn_r_34, u2_desIn_r_35, u2_desIn_r_36, u2_desIn_r_37, u2_desIn_r_38, u2_desIn_r_39, u2_desIn_r_4, u2_desIn_r_40, 
       u2_desIn_r_41, u2_desIn_r_42, u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_45, u2_desIn_r_46, u2_desIn_r_47, u2_desIn_r_48, u2_desIn_r_49, 
       u2_desIn_r_5, u2_desIn_r_50, u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_53, u2_desIn_r_54, u2_desIn_r_55, u2_desIn_r_56, u2_desIn_r_58, 
       u2_desIn_r_59, u2_desIn_r_6, u2_desIn_r_60, u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_63, u2_desIn_r_7, u2_desIn_r_8, u2_desIn_r_9, 
       u2_key_r_0, u2_key_r_1, u2_key_r_10, u2_key_r_11, u2_key_r_12, u2_key_r_13, u2_key_r_15, u2_key_r_16, u2_key_r_17, 
       u2_key_r_18, u2_key_r_19, u2_key_r_2, u2_key_r_20, u2_key_r_21, u2_key_r_22, u2_key_r_24, u2_key_r_25, u2_key_r_26, 
       u2_key_r_27, u2_key_r_28, u2_key_r_29, u2_key_r_3, u2_key_r_31, u2_key_r_32, u2_key_r_33, u2_key_r_34, u2_key_r_35, 
       u2_key_r_36, u2_key_r_37, u2_key_r_38, u2_key_r_39, u2_key_r_4, u2_key_r_40, u2_key_r_41, u2_key_r_42, u2_key_r_43, 
       u2_key_r_44, u2_key_r_45, u2_key_r_46, u2_key_r_47, u2_key_r_48, u2_key_r_49, u2_key_r_5, u2_key_r_50, u2_key_r_51, 
       u2_key_r_52, u2_key_r_53, u2_key_r_54, u2_key_r_55, u2_key_r_6, u2_key_r_8, u2_key_r_9, u2_out0_1, u2_out0_10, 
       u2_out0_16, u2_out0_17, u2_out0_20, u2_out0_23, u2_out0_24, u2_out0_26, u2_out0_30, u2_out0_31, u2_out0_6, 
       u2_out0_9, u2_out10_17, u2_out10_23, u2_out10_31, u2_out10_9, u2_out12_1, u2_out12_10, u2_out12_16, u2_out12_20, 
       u2_out12_24, u2_out12_26, u2_out12_30, u2_out12_6, u2_out13_1, u2_out13_10, u2_out13_13, u2_out13_16, u2_out13_17, 
       u2_out13_18, u2_out13_2, u2_out13_20, u2_out13_23, u2_out13_24, u2_out13_26, u2_out13_28, u2_out13_30, u2_out13_31, 
       u2_out13_6, u2_out13_9, u2_out3_12, u2_out3_22, u2_out3_32, u2_out3_7, u2_out7_11, u2_out7_12, u2_out7_14, 
       u2_out7_19, u2_out7_22, u2_out7_25, u2_out7_29, u2_out7_3, u2_out7_32, u2_out7_4, u2_out7_7, u2_out7_8, 
       u2_u0_X_1, u2_u0_X_13, u2_u0_X_14, u2_u0_X_15, u2_u0_X_16, u2_u0_X_17, u2_u0_X_18, u2_u0_X_19, u2_u0_X_2, 
       u2_u0_X_20, u2_u0_X_21, u2_u0_X_22, u2_u0_X_23, u2_u0_X_24, u2_u0_X_3, u2_u0_X_4, u2_u0_X_5, u2_u0_X_6, 
       u2_u0_u0_n100, u2_u0_u0_n101, u2_u0_u0_n102, u2_u0_u0_n103, u2_u0_u0_n104, u2_u0_u0_n105, u2_u0_u0_n106, u2_u0_u0_n107, u2_u0_u0_n108, 
       u2_u0_u0_n109, u2_u0_u0_n110, u2_u0_u0_n111, u2_u0_u0_n112, u2_u0_u0_n113, u2_u0_u0_n114, u2_u0_u0_n115, u2_u0_u0_n116, u2_u0_u0_n117, 
       u2_u0_u0_n118, u2_u0_u0_n119, u2_u0_u0_n120, u2_u0_u0_n121, u2_u0_u0_n122, u2_u0_u0_n123, u2_u0_u0_n124, u2_u0_u0_n125, u2_u0_u0_n126, 
       u2_u0_u0_n127, u2_u0_u0_n128, u2_u0_u0_n129, u2_u0_u0_n130, u2_u0_u0_n131, u2_u0_u0_n132, u2_u0_u0_n133, u2_u0_u0_n134, u2_u0_u0_n135, 
       u2_u0_u0_n136, u2_u0_u0_n137, u2_u0_u0_n138, u2_u0_u0_n139, u2_u0_u0_n140, u2_u0_u0_n141, u2_u0_u0_n142, u2_u0_u0_n143, u2_u0_u0_n144, 
       u2_u0_u0_n145, u2_u0_u0_n146, u2_u0_u0_n147, u2_u0_u0_n148, u2_u0_u0_n149, u2_u0_u0_n150, u2_u0_u0_n151, u2_u0_u0_n152, u2_u0_u0_n153, 
       u2_u0_u0_n154, u2_u0_u0_n155, u2_u0_u0_n156, u2_u0_u0_n157, u2_u0_u0_n158, u2_u0_u0_n159, u2_u0_u0_n160, u2_u0_u0_n161, u2_u0_u0_n162, 
       u2_u0_u0_n163, u2_u0_u0_n164, u2_u0_u0_n165, u2_u0_u0_n166, u2_u0_u0_n167, u2_u0_u0_n168, u2_u0_u0_n169, u2_u0_u0_n170, u2_u0_u0_n171, 
       u2_u0_u0_n172, u2_u0_u0_n173, u2_u0_u0_n174, u2_u0_u0_n88, u2_u0_u0_n89, u2_u0_u0_n90, u2_u0_u0_n91, u2_u0_u0_n92, u2_u0_u0_n93, 
       u2_u0_u0_n94, u2_u0_u0_n95, u2_u0_u0_n96, u2_u0_u0_n97, u2_u0_u0_n98, u2_u0_u0_n99, u2_u0_u2_n100, u2_u0_u2_n101, u2_u0_u2_n102, 
       u2_u0_u2_n103, u2_u0_u2_n104, u2_u0_u2_n105, u2_u0_u2_n106, u2_u0_u2_n107, u2_u0_u2_n108, u2_u0_u2_n109, u2_u0_u2_n110, u2_u0_u2_n111, 
       u2_u0_u2_n112, u2_u0_u2_n113, u2_u0_u2_n114, u2_u0_u2_n115, u2_u0_u2_n116, u2_u0_u2_n117, u2_u0_u2_n118, u2_u0_u2_n119, u2_u0_u2_n120, 
       u2_u0_u2_n121, u2_u0_u2_n122, u2_u0_u2_n123, u2_u0_u2_n124, u2_u0_u2_n125, u2_u0_u2_n126, u2_u0_u2_n127, u2_u0_u2_n128, u2_u0_u2_n129, 
       u2_u0_u2_n130, u2_u0_u2_n131, u2_u0_u2_n132, u2_u0_u2_n133, u2_u0_u2_n134, u2_u0_u2_n135, u2_u0_u2_n136, u2_u0_u2_n137, u2_u0_u2_n138, 
       u2_u0_u2_n139, u2_u0_u2_n140, u2_u0_u2_n141, u2_u0_u2_n142, u2_u0_u2_n143, u2_u0_u2_n144, u2_u0_u2_n145, u2_u0_u2_n146, u2_u0_u2_n147, 
       u2_u0_u2_n148, u2_u0_u2_n149, u2_u0_u2_n150, u2_u0_u2_n151, u2_u0_u2_n152, u2_u0_u2_n153, u2_u0_u2_n154, u2_u0_u2_n155, u2_u0_u2_n156, 
       u2_u0_u2_n157, u2_u0_u2_n158, u2_u0_u2_n159, u2_u0_u2_n160, u2_u0_u2_n161, u2_u0_u2_n162, u2_u0_u2_n163, u2_u0_u2_n164, u2_u0_u2_n165, 
       u2_u0_u2_n166, u2_u0_u2_n167, u2_u0_u2_n168, u2_u0_u2_n169, u2_u0_u2_n170, u2_u0_u2_n171, u2_u0_u2_n172, u2_u0_u2_n173, u2_u0_u2_n174, 
       u2_u0_u2_n175, u2_u0_u2_n176, u2_u0_u2_n177, u2_u0_u2_n178, u2_u0_u2_n179, u2_u0_u2_n180, u2_u0_u2_n181, u2_u0_u2_n182, u2_u0_u2_n183, 
       u2_u0_u2_n184, u2_u0_u2_n185, u2_u0_u2_n186, u2_u0_u2_n187, u2_u0_u2_n188, u2_u0_u2_n95, u2_u0_u2_n96, u2_u0_u2_n97, u2_u0_u2_n98, 
       u2_u0_u2_n99, u2_u0_u3_n100, u2_u0_u3_n101, u2_u0_u3_n102, u2_u0_u3_n103, u2_u0_u3_n104, u2_u0_u3_n105, u2_u0_u3_n106, u2_u0_u3_n107, 
       u2_u0_u3_n108, u2_u0_u3_n109, u2_u0_u3_n110, u2_u0_u3_n111, u2_u0_u3_n112, u2_u0_u3_n113, u2_u0_u3_n114, u2_u0_u3_n115, u2_u0_u3_n116, 
       u2_u0_u3_n117, u2_u0_u3_n118, u2_u0_u3_n119, u2_u0_u3_n120, u2_u0_u3_n121, u2_u0_u3_n122, u2_u0_u3_n123, u2_u0_u3_n124, u2_u0_u3_n125, 
       u2_u0_u3_n126, u2_u0_u3_n127, u2_u0_u3_n128, u2_u0_u3_n129, u2_u0_u3_n130, u2_u0_u3_n131, u2_u0_u3_n132, u2_u0_u3_n133, u2_u0_u3_n134, 
       u2_u0_u3_n135, u2_u0_u3_n136, u2_u0_u3_n137, u2_u0_u3_n138, u2_u0_u3_n139, u2_u0_u3_n140, u2_u0_u3_n141, u2_u0_u3_n142, u2_u0_u3_n143, 
       u2_u0_u3_n144, u2_u0_u3_n145, u2_u0_u3_n146, u2_u0_u3_n147, u2_u0_u3_n148, u2_u0_u3_n149, u2_u0_u3_n150, u2_u0_u3_n151, u2_u0_u3_n152, 
       u2_u0_u3_n153, u2_u0_u3_n154, u2_u0_u3_n155, u2_u0_u3_n156, u2_u0_u3_n157, u2_u0_u3_n158, u2_u0_u3_n159, u2_u0_u3_n160, u2_u0_u3_n161, 
       u2_u0_u3_n162, u2_u0_u3_n163, u2_u0_u3_n164, u2_u0_u3_n165, u2_u0_u3_n166, u2_u0_u3_n167, u2_u0_u3_n168, u2_u0_u3_n169, u2_u0_u3_n170, 
       u2_u0_u3_n171, u2_u0_u3_n172, u2_u0_u3_n173, u2_u0_u3_n174, u2_u0_u3_n175, u2_u0_u3_n176, u2_u0_u3_n177, u2_u0_u3_n178, u2_u0_u3_n179, 
       u2_u0_u3_n180, u2_u0_u3_n181, u2_u0_u3_n182, u2_u0_u3_n183, u2_u0_u3_n184, u2_u0_u3_n185, u2_u0_u3_n186, u2_u0_u3_n94, u2_u0_u3_n95, 
       u2_u0_u3_n96, u2_u0_u3_n97, u2_u0_u3_n98, u2_u0_u3_n99, u2_u10_X_1, u2_u10_X_2, u2_u10_X_3, u2_u10_X_4, u2_u10_X_5, 
       u2_u10_X_6, u2_u10_u0_n100, u2_u10_u0_n101, u2_u10_u0_n102, u2_u10_u0_n103, u2_u10_u0_n104, u2_u10_u0_n105, u2_u10_u0_n106, u2_u10_u0_n107, 
       u2_u10_u0_n108, u2_u10_u0_n109, u2_u10_u0_n110, u2_u10_u0_n111, u2_u10_u0_n112, u2_u10_u0_n113, u2_u10_u0_n114, u2_u10_u0_n115, u2_u10_u0_n116, 
       u2_u10_u0_n117, u2_u10_u0_n118, u2_u10_u0_n119, u2_u10_u0_n120, u2_u10_u0_n121, u2_u10_u0_n122, u2_u10_u0_n123, u2_u10_u0_n124, u2_u10_u0_n125, 
       u2_u10_u0_n126, u2_u10_u0_n127, u2_u10_u0_n128, u2_u10_u0_n129, u2_u10_u0_n130, u2_u10_u0_n131, u2_u10_u0_n132, u2_u10_u0_n133, u2_u10_u0_n134, 
       u2_u10_u0_n135, u2_u10_u0_n136, u2_u10_u0_n137, u2_u10_u0_n138, u2_u10_u0_n139, u2_u10_u0_n140, u2_u10_u0_n141, u2_u10_u0_n142, u2_u10_u0_n143, 
       u2_u10_u0_n144, u2_u10_u0_n145, u2_u10_u0_n146, u2_u10_u0_n147, u2_u10_u0_n148, u2_u10_u0_n149, u2_u10_u0_n150, u2_u10_u0_n151, u2_u10_u0_n152, 
       u2_u10_u0_n153, u2_u10_u0_n154, u2_u10_u0_n155, u2_u10_u0_n156, u2_u10_u0_n157, u2_u10_u0_n158, u2_u10_u0_n159, u2_u10_u0_n160, u2_u10_u0_n161, 
       u2_u10_u0_n162, u2_u10_u0_n163, u2_u10_u0_n164, u2_u10_u0_n165, u2_u10_u0_n166, u2_u10_u0_n167, u2_u10_u0_n168, u2_u10_u0_n169, u2_u10_u0_n170, 
       u2_u10_u0_n171, u2_u10_u0_n172, u2_u10_u0_n173, u2_u10_u0_n174, u2_u10_u0_n88, u2_u10_u0_n89, u2_u10_u0_n90, u2_u10_u0_n91, u2_u10_u0_n92, 
       u2_u10_u0_n93, u2_u10_u0_n94, u2_u10_u0_n95, u2_u10_u0_n96, u2_u10_u0_n97, u2_u10_u0_n98, u2_u10_u0_n99, u2_u12_X_13, u2_u12_X_14, 
       u2_u12_X_15, u2_u12_X_16, u2_u12_X_17, u2_u12_X_18, u2_u12_X_19, u2_u12_X_20, u2_u12_X_21, u2_u12_X_22, u2_u12_X_23, 
       u2_u12_X_24, u2_u12_u2_n100, u2_u12_u2_n101, u2_u12_u2_n102, u2_u12_u2_n103, u2_u12_u2_n104, u2_u12_u2_n105, u2_u12_u2_n106, u2_u12_u2_n107, 
       u2_u12_u2_n108, u2_u12_u2_n109, u2_u12_u2_n110, u2_u12_u2_n111, u2_u12_u2_n112, u2_u12_u2_n113, u2_u12_u2_n114, u2_u12_u2_n115, u2_u12_u2_n116, 
       u2_u12_u2_n117, u2_u12_u2_n118, u2_u12_u2_n119, u2_u12_u2_n120, u2_u12_u2_n121, u2_u12_u2_n122, u2_u12_u2_n123, u2_u12_u2_n124, u2_u12_u2_n125, 
       u2_u12_u2_n126, u2_u12_u2_n127, u2_u12_u2_n128, u2_u12_u2_n129, u2_u12_u2_n130, u2_u12_u2_n131, u2_u12_u2_n132, u2_u12_u2_n133, u2_u12_u2_n134, 
       u2_u12_u2_n135, u2_u12_u2_n136, u2_u12_u2_n137, u2_u12_u2_n138, u2_u12_u2_n139, u2_u12_u2_n140, u2_u12_u2_n141, u2_u12_u2_n142, u2_u12_u2_n143, 
       u2_u12_u2_n144, u2_u12_u2_n145, u2_u12_u2_n146, u2_u12_u2_n147, u2_u12_u2_n148, u2_u12_u2_n149, u2_u12_u2_n150, u2_u12_u2_n151, u2_u12_u2_n152, 
       u2_u12_u2_n153, u2_u12_u2_n154, u2_u12_u2_n155, u2_u12_u2_n156, u2_u12_u2_n157, u2_u12_u2_n158, u2_u12_u2_n159, u2_u12_u2_n160, u2_u12_u2_n161, 
       u2_u12_u2_n162, u2_u12_u2_n163, u2_u12_u2_n164, u2_u12_u2_n165, u2_u12_u2_n166, u2_u12_u2_n167, u2_u12_u2_n168, u2_u12_u2_n169, u2_u12_u2_n170, 
       u2_u12_u2_n171, u2_u12_u2_n172, u2_u12_u2_n173, u2_u12_u2_n174, u2_u12_u2_n175, u2_u12_u2_n176, u2_u12_u2_n177, u2_u12_u2_n178, u2_u12_u2_n179, 
       u2_u12_u2_n180, u2_u12_u2_n181, u2_u12_u2_n182, u2_u12_u2_n183, u2_u12_u2_n184, u2_u12_u2_n185, u2_u12_u2_n186, u2_u12_u2_n187, u2_u12_u2_n188, 
       u2_u12_u2_n95, u2_u12_u2_n96, u2_u12_u2_n97, u2_u12_u2_n98, u2_u12_u2_n99, u2_u12_u3_n100, u2_u12_u3_n101, u2_u12_u3_n102, u2_u12_u3_n103, 
       u2_u12_u3_n104, u2_u12_u3_n105, u2_u12_u3_n106, u2_u12_u3_n107, u2_u12_u3_n108, u2_u12_u3_n109, u2_u12_u3_n110, u2_u12_u3_n111, u2_u12_u3_n112, 
       u2_u12_u3_n113, u2_u12_u3_n114, u2_u12_u3_n115, u2_u12_u3_n116, u2_u12_u3_n117, u2_u12_u3_n118, u2_u12_u3_n119, u2_u12_u3_n120, u2_u12_u3_n121, 
       u2_u12_u3_n122, u2_u12_u3_n123, u2_u12_u3_n124, u2_u12_u3_n125, u2_u12_u3_n126, u2_u12_u3_n127, u2_u12_u3_n128, u2_u12_u3_n129, u2_u12_u3_n130, 
       u2_u12_u3_n131, u2_u12_u3_n132, u2_u12_u3_n133, u2_u12_u3_n134, u2_u12_u3_n135, u2_u12_u3_n136, u2_u12_u3_n137, u2_u12_u3_n138, u2_u12_u3_n139, 
       u2_u12_u3_n140, u2_u12_u3_n141, u2_u12_u3_n142, u2_u12_u3_n143, u2_u12_u3_n144, u2_u12_u3_n145, u2_u12_u3_n146, u2_u12_u3_n147, u2_u12_u3_n148, 
       u2_u12_u3_n149, u2_u12_u3_n150, u2_u12_u3_n151, u2_u12_u3_n152, u2_u12_u3_n153, u2_u12_u3_n154, u2_u12_u3_n155, u2_u12_u3_n156, u2_u12_u3_n157, 
       u2_u12_u3_n158, u2_u12_u3_n159, u2_u12_u3_n160, u2_u12_u3_n161, u2_u12_u3_n162, u2_u12_u3_n163, u2_u12_u3_n164, u2_u12_u3_n165, u2_u12_u3_n166, 
       u2_u12_u3_n167, u2_u12_u3_n168, u2_u12_u3_n169, u2_u12_u3_n170, u2_u12_u3_n171, u2_u12_u3_n172, u2_u12_u3_n173, u2_u12_u3_n174, u2_u12_u3_n175, 
       u2_u12_u3_n176, u2_u12_u3_n177, u2_u12_u3_n178, u2_u12_u3_n179, u2_u12_u3_n180, u2_u12_u3_n181, u2_u12_u3_n182, u2_u12_u3_n183, u2_u12_u3_n184, 
       u2_u12_u3_n185, u2_u12_u3_n186, u2_u12_u3_n94, u2_u12_u3_n95, u2_u12_u3_n96, u2_u12_u3_n97, u2_u12_u3_n98, u2_u12_u3_n99, u2_u13_X_1, 
       u2_u13_X_10, u2_u13_X_11, u2_u13_X_12, u2_u13_X_13, u2_u13_X_14, u2_u13_X_15, u2_u13_X_16, u2_u13_X_17, u2_u13_X_18, 
       u2_u13_X_19, u2_u13_X_2, u2_u13_X_20, u2_u13_X_21, u2_u13_X_22, u2_u13_X_23, u2_u13_X_24, u2_u13_X_3, u2_u13_X_4, 
       u2_u13_X_5, u2_u13_X_6, u2_u13_X_7, u2_u13_X_8, u2_u13_X_9, u2_u13_u0_n100, u2_u13_u0_n101, u2_u13_u0_n102, u2_u13_u0_n103, 
       u2_u13_u0_n104, u2_u13_u0_n105, u2_u13_u0_n106, u2_u13_u0_n107, u2_u13_u0_n108, u2_u13_u0_n109, u2_u13_u0_n110, u2_u13_u0_n111, u2_u13_u0_n112, 
       u2_u13_u0_n113, u2_u13_u0_n114, u2_u13_u0_n115, u2_u13_u0_n116, u2_u13_u0_n117, u2_u13_u0_n118, u2_u13_u0_n119, u2_u13_u0_n120, u2_u13_u0_n121, 
       u2_u13_u0_n122, u2_u13_u0_n123, u2_u13_u0_n124, u2_u13_u0_n125, u2_u13_u0_n126, u2_u13_u0_n127, u2_u13_u0_n128, u2_u13_u0_n129, u2_u13_u0_n130, 
       u2_u13_u0_n131, u2_u13_u0_n132, u2_u13_u0_n133, u2_u13_u0_n134, u2_u13_u0_n135, u2_u13_u0_n136, u2_u13_u0_n137, u2_u13_u0_n138, u2_u13_u0_n139, 
       u2_u13_u0_n140, u2_u13_u0_n141, u2_u13_u0_n142, u2_u13_u0_n143, u2_u13_u0_n144, u2_u13_u0_n145, u2_u13_u0_n146, u2_u13_u0_n147, u2_u13_u0_n148, 
       u2_u13_u0_n149, u2_u13_u0_n150, u2_u13_u0_n151, u2_u13_u0_n152, u2_u13_u0_n153, u2_u13_u0_n154, u2_u13_u0_n155, u2_u13_u0_n156, u2_u13_u0_n157, 
       u2_u13_u0_n158, u2_u13_u0_n159, u2_u13_u0_n160, u2_u13_u0_n161, u2_u13_u0_n162, u2_u13_u0_n163, u2_u13_u0_n164, u2_u13_u0_n165, u2_u13_u0_n166, 
       u2_u13_u0_n167, u2_u13_u0_n168, u2_u13_u0_n169, u2_u13_u0_n170, u2_u13_u0_n171, u2_u13_u0_n172, u2_u13_u0_n173, u2_u13_u0_n174, u2_u13_u0_n88, 
       u2_u13_u0_n89, u2_u13_u0_n90, u2_u13_u0_n91, u2_u13_u0_n92, u2_u13_u0_n93, u2_u13_u0_n94, u2_u13_u0_n95, u2_u13_u0_n96, u2_u13_u0_n97, 
       u2_u13_u0_n98, u2_u13_u0_n99, u2_u13_u1_n100, u2_u13_u1_n101, u2_u13_u1_n102, u2_u13_u1_n103, u2_u13_u1_n104, u2_u13_u1_n105, u2_u13_u1_n106, 
       u2_u13_u1_n107, u2_u13_u1_n108, u2_u13_u1_n109, u2_u13_u1_n110, u2_u13_u1_n111, u2_u13_u1_n112, u2_u13_u1_n113, u2_u13_u1_n114, u2_u13_u1_n115, 
       u2_u13_u1_n116, u2_u13_u1_n117, u2_u13_u1_n118, u2_u13_u1_n119, u2_u13_u1_n120, u2_u13_u1_n121, u2_u13_u1_n122, u2_u13_u1_n123, u2_u13_u1_n124, 
       u2_u13_u1_n125, u2_u13_u1_n126, u2_u13_u1_n127, u2_u13_u1_n128, u2_u13_u1_n129, u2_u13_u1_n130, u2_u13_u1_n131, u2_u13_u1_n132, u2_u13_u1_n133, 
       u2_u13_u1_n134, u2_u13_u1_n135, u2_u13_u1_n136, u2_u13_u1_n137, u2_u13_u1_n138, u2_u13_u1_n139, u2_u13_u1_n140, u2_u13_u1_n141, u2_u13_u1_n142, 
       u2_u13_u1_n143, u2_u13_u1_n144, u2_u13_u1_n145, u2_u13_u1_n146, u2_u13_u1_n147, u2_u13_u1_n148, u2_u13_u1_n149, u2_u13_u1_n150, u2_u13_u1_n151, 
       u2_u13_u1_n152, u2_u13_u1_n153, u2_u13_u1_n154, u2_u13_u1_n155, u2_u13_u1_n156, u2_u13_u1_n157, u2_u13_u1_n158, u2_u13_u1_n159, u2_u13_u1_n160, 
       u2_u13_u1_n161, u2_u13_u1_n162, u2_u13_u1_n163, u2_u13_u1_n164, u2_u13_u1_n165, u2_u13_u1_n166, u2_u13_u1_n167, u2_u13_u1_n168, u2_u13_u1_n169, 
       u2_u13_u1_n170, u2_u13_u1_n171, u2_u13_u1_n172, u2_u13_u1_n173, u2_u13_u1_n174, u2_u13_u1_n175, u2_u13_u1_n176, u2_u13_u1_n177, u2_u13_u1_n178, 
       u2_u13_u1_n179, u2_u13_u1_n180, u2_u13_u1_n181, u2_u13_u1_n182, u2_u13_u1_n183, u2_u13_u1_n184, u2_u13_u1_n185, u2_u13_u1_n186, u2_u13_u1_n187, 
       u2_u13_u1_n188, u2_u13_u1_n95, u2_u13_u1_n96, u2_u13_u1_n97, u2_u13_u1_n98, u2_u13_u1_n99, u2_u13_u2_n100, u2_u13_u2_n101, u2_u13_u2_n102, 
       u2_u13_u2_n103, u2_u13_u2_n104, u2_u13_u2_n105, u2_u13_u2_n106, u2_u13_u2_n107, u2_u13_u2_n108, u2_u13_u2_n109, u2_u13_u2_n110, u2_u13_u2_n111, 
       u2_u13_u2_n112, u2_u13_u2_n113, u2_u13_u2_n114, u2_u13_u2_n115, u2_u13_u2_n116, u2_u13_u2_n117, u2_u13_u2_n118, u2_u13_u2_n119, u2_u13_u2_n120, 
       u2_u13_u2_n121, u2_u13_u2_n122, u2_u13_u2_n123, u2_u13_u2_n124, u2_u13_u2_n125, u2_u13_u2_n126, u2_u13_u2_n127, u2_u13_u2_n128, u2_u13_u2_n129, 
       u2_u13_u2_n130, u2_u13_u2_n131, u2_u13_u2_n132, u2_u13_u2_n133, u2_u13_u2_n134, u2_u13_u2_n135, u2_u13_u2_n136, u2_u13_u2_n137, u2_u13_u2_n138, 
       u2_u13_u2_n139, u2_u13_u2_n140, u2_u13_u2_n141, u2_u13_u2_n142, u2_u13_u2_n143, u2_u13_u2_n144, u2_u13_u2_n145, u2_u13_u2_n146, u2_u13_u2_n147, 
       u2_u13_u2_n148, u2_u13_u2_n149, u2_u13_u2_n150, u2_u13_u2_n151, u2_u13_u2_n152, u2_u13_u2_n153, u2_u13_u2_n154, u2_u13_u2_n155, u2_u13_u2_n156, 
       u2_u13_u2_n157, u2_u13_u2_n158, u2_u13_u2_n159, u2_u13_u2_n160, u2_u13_u2_n161, u2_u13_u2_n162, u2_u13_u2_n163, u2_u13_u2_n164, u2_u13_u2_n165, 
       u2_u13_u2_n166, u2_u13_u2_n167, u2_u13_u2_n168, u2_u13_u2_n169, u2_u13_u2_n170, u2_u13_u2_n171, u2_u13_u2_n172, u2_u13_u2_n173, u2_u13_u2_n174, 
       u2_u13_u2_n175, u2_u13_u2_n176, u2_u13_u2_n177, u2_u13_u2_n178, u2_u13_u2_n179, u2_u13_u2_n180, u2_u13_u2_n181, u2_u13_u2_n182, u2_u13_u2_n183, 
       u2_u13_u2_n184, u2_u13_u2_n185, u2_u13_u2_n186, u2_u13_u2_n187, u2_u13_u2_n188, u2_u13_u2_n95, u2_u13_u2_n96, u2_u13_u2_n97, u2_u13_u2_n98, 
       u2_u13_u2_n99, u2_u13_u3_n100, u2_u13_u3_n101, u2_u13_u3_n102, u2_u13_u3_n103, u2_u13_u3_n104, u2_u13_u3_n105, u2_u13_u3_n106, u2_u13_u3_n107, 
       u2_u13_u3_n108, u2_u13_u3_n109, u2_u13_u3_n110, u2_u13_u3_n111, u2_u13_u3_n112, u2_u13_u3_n113, u2_u13_u3_n114, u2_u13_u3_n115, u2_u13_u3_n116, 
       u2_u13_u3_n117, u2_u13_u3_n118, u2_u13_u3_n119, u2_u13_u3_n120, u2_u13_u3_n121, u2_u13_u3_n122, u2_u13_u3_n123, u2_u13_u3_n124, u2_u13_u3_n125, 
       u2_u13_u3_n126, u2_u13_u3_n127, u2_u13_u3_n128, u2_u13_u3_n129, u2_u13_u3_n130, u2_u13_u3_n131, u2_u13_u3_n132, u2_u13_u3_n133, u2_u13_u3_n134, 
       u2_u13_u3_n135, u2_u13_u3_n136, u2_u13_u3_n137, u2_u13_u3_n138, u2_u13_u3_n139, u2_u13_u3_n140, u2_u13_u3_n141, u2_u13_u3_n142, u2_u13_u3_n143, 
       u2_u13_u3_n144, u2_u13_u3_n145, u2_u13_u3_n146, u2_u13_u3_n147, u2_u13_u3_n148, u2_u13_u3_n149, u2_u13_u3_n150, u2_u13_u3_n151, u2_u13_u3_n152, 
       u2_u13_u3_n153, u2_u13_u3_n154, u2_u13_u3_n155, u2_u13_u3_n156, u2_u13_u3_n157, u2_u13_u3_n158, u2_u13_u3_n159, u2_u13_u3_n160, u2_u13_u3_n161, 
       u2_u13_u3_n162, u2_u13_u3_n163, u2_u13_u3_n164, u2_u13_u3_n165, u2_u13_u3_n166, u2_u13_u3_n167, u2_u13_u3_n168, u2_u13_u3_n169, u2_u13_u3_n170, 
       u2_u13_u3_n171, u2_u13_u3_n172, u2_u13_u3_n173, u2_u13_u3_n174, u2_u13_u3_n175, u2_u13_u3_n176, u2_u13_u3_n177, u2_u13_u3_n178, u2_u13_u3_n179, 
       u2_u13_u3_n180, u2_u13_u3_n181, u2_u13_u3_n182, u2_u13_u3_n183, u2_u13_u3_n184, u2_u13_u3_n185, u2_u13_u3_n186, u2_u13_u3_n94, u2_u13_u3_n95, 
       u2_u13_u3_n96, u2_u13_u3_n97, u2_u13_u3_n98, u2_u13_u3_n99, u2_u3_X_37, u2_u3_X_38, u2_u3_X_39, u2_u3_X_40, u2_u3_X_41, 
       u2_u3_X_42, u2_u3_u6_n100, u2_u3_u6_n101, u2_u3_u6_n102, u2_u3_u6_n103, u2_u3_u6_n104, u2_u3_u6_n105, u2_u3_u6_n106, u2_u3_u6_n107, 
       u2_u3_u6_n108, u2_u3_u6_n109, u2_u3_u6_n110, u2_u3_u6_n111, u2_u3_u6_n112, u2_u3_u6_n113, u2_u3_u6_n114, u2_u3_u6_n115, u2_u3_u6_n116, 
       u2_u3_u6_n117, u2_u3_u6_n118, u2_u3_u6_n119, u2_u3_u6_n120, u2_u3_u6_n121, u2_u3_u6_n122, u2_u3_u6_n123, u2_u3_u6_n124, u2_u3_u6_n125, 
       u2_u3_u6_n126, u2_u3_u6_n127, u2_u3_u6_n128, u2_u3_u6_n129, u2_u3_u6_n130, u2_u3_u6_n131, u2_u3_u6_n132, u2_u3_u6_n133, u2_u3_u6_n134, 
       u2_u3_u6_n135, u2_u3_u6_n136, u2_u3_u6_n137, u2_u3_u6_n138, u2_u3_u6_n139, u2_u3_u6_n140, u2_u3_u6_n141, u2_u3_u6_n142, u2_u3_u6_n143, 
       u2_u3_u6_n144, u2_u3_u6_n145, u2_u3_u6_n146, u2_u3_u6_n147, u2_u3_u6_n148, u2_u3_u6_n149, u2_u3_u6_n150, u2_u3_u6_n151, u2_u3_u6_n152, 
       u2_u3_u6_n153, u2_u3_u6_n154, u2_u3_u6_n155, u2_u3_u6_n156, u2_u3_u6_n157, u2_u3_u6_n158, u2_u3_u6_n159, u2_u3_u6_n160, u2_u3_u6_n161, 
       u2_u3_u6_n162, u2_u3_u6_n163, u2_u3_u6_n164, u2_u3_u6_n165, u2_u3_u6_n166, u2_u3_u6_n167, u2_u3_u6_n168, u2_u3_u6_n169, u2_u3_u6_n170, 
       u2_u3_u6_n171, u2_u3_u6_n172, u2_u3_u6_n173, u2_u3_u6_n174, u2_u3_u6_n88, u2_u3_u6_n89, u2_u3_u6_n90, u2_u3_u6_n91, u2_u3_u6_n92, 
       u2_u3_u6_n93, u2_u3_u6_n94, u2_u3_u6_n95, u2_u3_u6_n96, u2_u3_u6_n97, u2_u3_u6_n98, u2_u3_u6_n99, u2_u7_X_25, u2_u7_X_26, 
       u2_u7_X_27, u2_u7_X_28, u2_u7_X_29, u2_u7_X_30, u2_u7_X_31, u2_u7_X_32, u2_u7_X_33, u2_u7_X_34, u2_u7_X_35, 
       u2_u7_X_36, u2_u7_X_37, u2_u7_X_38, u2_u7_X_39, u2_u7_X_40, u2_u7_X_41, u2_u7_X_42, u2_u7_u4_n100, u2_u7_u4_n101, 
       u2_u7_u4_n102, u2_u7_u4_n103, u2_u7_u4_n104, u2_u7_u4_n105, u2_u7_u4_n106, u2_u7_u4_n107, u2_u7_u4_n108, u2_u7_u4_n109, u2_u7_u4_n110, 
       u2_u7_u4_n111, u2_u7_u4_n112, u2_u7_u4_n113, u2_u7_u4_n114, u2_u7_u4_n115, u2_u7_u4_n116, u2_u7_u4_n117, u2_u7_u4_n118, u2_u7_u4_n119, 
       u2_u7_u4_n120, u2_u7_u4_n121, u2_u7_u4_n122, u2_u7_u4_n123, u2_u7_u4_n124, u2_u7_u4_n125, u2_u7_u4_n126, u2_u7_u4_n127, u2_u7_u4_n128, 
       u2_u7_u4_n129, u2_u7_u4_n130, u2_u7_u4_n131, u2_u7_u4_n132, u2_u7_u4_n133, u2_u7_u4_n134, u2_u7_u4_n135, u2_u7_u4_n136, u2_u7_u4_n137, 
       u2_u7_u4_n138, u2_u7_u4_n139, u2_u7_u4_n140, u2_u7_u4_n141, u2_u7_u4_n142, u2_u7_u4_n143, u2_u7_u4_n144, u2_u7_u4_n145, u2_u7_u4_n146, 
       u2_u7_u4_n147, u2_u7_u4_n148, u2_u7_u4_n149, u2_u7_u4_n150, u2_u7_u4_n151, u2_u7_u4_n152, u2_u7_u4_n153, u2_u7_u4_n154, u2_u7_u4_n155, 
       u2_u7_u4_n156, u2_u7_u4_n157, u2_u7_u4_n158, u2_u7_u4_n159, u2_u7_u4_n160, u2_u7_u4_n161, u2_u7_u4_n162, u2_u7_u4_n163, u2_u7_u4_n164, 
       u2_u7_u4_n165, u2_u7_u4_n166, u2_u7_u4_n167, u2_u7_u4_n168, u2_u7_u4_n169, u2_u7_u4_n170, u2_u7_u4_n171, u2_u7_u4_n172, u2_u7_u4_n173, 
       u2_u7_u4_n174, u2_u7_u4_n175, u2_u7_u4_n176, u2_u7_u4_n177, u2_u7_u4_n178, u2_u7_u4_n179, u2_u7_u4_n180, u2_u7_u4_n181, u2_u7_u4_n182, 
       u2_u7_u4_n183, u2_u7_u4_n184, u2_u7_u4_n185, u2_u7_u4_n186, u2_u7_u4_n94, u2_u7_u4_n95, u2_u7_u4_n96, u2_u7_u4_n97, u2_u7_u4_n98, 
       u2_u7_u4_n99, u2_u7_u5_n100, u2_u7_u5_n101, u2_u7_u5_n102, u2_u7_u5_n103, u2_u7_u5_n104, u2_u7_u5_n105, u2_u7_u5_n106, u2_u7_u5_n107, 
       u2_u7_u5_n108, u2_u7_u5_n109, u2_u7_u5_n110, u2_u7_u5_n111, u2_u7_u5_n112, u2_u7_u5_n113, u2_u7_u5_n114, u2_u7_u5_n115, u2_u7_u5_n116, 
       u2_u7_u5_n117, u2_u7_u5_n118, u2_u7_u5_n119, u2_u7_u5_n120, u2_u7_u5_n121, u2_u7_u5_n122, u2_u7_u5_n123, u2_u7_u5_n124, u2_u7_u5_n125, 
       u2_u7_u5_n126, u2_u7_u5_n127, u2_u7_u5_n128, u2_u7_u5_n129, u2_u7_u5_n130, u2_u7_u5_n131, u2_u7_u5_n132, u2_u7_u5_n133, u2_u7_u5_n134, 
       u2_u7_u5_n135, u2_u7_u5_n136, u2_u7_u5_n137, u2_u7_u5_n138, u2_u7_u5_n139, u2_u7_u5_n140, u2_u7_u5_n141, u2_u7_u5_n142, u2_u7_u5_n143, 
       u2_u7_u5_n144, u2_u7_u5_n145, u2_u7_u5_n146, u2_u7_u5_n147, u2_u7_u5_n148, u2_u7_u5_n149, u2_u7_u5_n150, u2_u7_u5_n151, u2_u7_u5_n152, 
       u2_u7_u5_n153, u2_u7_u5_n154, u2_u7_u5_n155, u2_u7_u5_n156, u2_u7_u5_n157, u2_u7_u5_n158, u2_u7_u5_n159, u2_u7_u5_n160, u2_u7_u5_n161, 
       u2_u7_u5_n162, u2_u7_u5_n163, u2_u7_u5_n164, u2_u7_u5_n165, u2_u7_u5_n166, u2_u7_u5_n167, u2_u7_u5_n168, u2_u7_u5_n169, u2_u7_u5_n170, 
       u2_u7_u5_n171, u2_u7_u5_n172, u2_u7_u5_n173, u2_u7_u5_n174, u2_u7_u5_n175, u2_u7_u5_n176, u2_u7_u5_n177, u2_u7_u5_n178, u2_u7_u5_n179, 
       u2_u7_u5_n180, u2_u7_u5_n181, u2_u7_u5_n182, u2_u7_u5_n183, u2_u7_u5_n184, u2_u7_u5_n185, u2_u7_u5_n186, u2_u7_u5_n187, u2_u7_u5_n188, 
       u2_u7_u5_n189, u2_u7_u5_n190, u2_u7_u5_n191, u2_u7_u5_n192, u2_u7_u5_n193, u2_u7_u5_n194, u2_u7_u5_n195, u2_u7_u5_n196, u2_u7_u5_n99, 
       u2_u7_u6_n100, u2_u7_u6_n101, u2_u7_u6_n102, u2_u7_u6_n103, u2_u7_u6_n104, u2_u7_u6_n105, u2_u7_u6_n106, u2_u7_u6_n107, u2_u7_u6_n108, 
       u2_u7_u6_n109, u2_u7_u6_n110, u2_u7_u6_n111, u2_u7_u6_n112, u2_u7_u6_n113, u2_u7_u6_n114, u2_u7_u6_n115, u2_u7_u6_n116, u2_u7_u6_n117, 
       u2_u7_u6_n118, u2_u7_u6_n119, u2_u7_u6_n120, u2_u7_u6_n121, u2_u7_u6_n122, u2_u7_u6_n123, u2_u7_u6_n124, u2_u7_u6_n125, u2_u7_u6_n126, 
       u2_u7_u6_n127, u2_u7_u6_n128, u2_u7_u6_n129, u2_u7_u6_n130, u2_u7_u6_n131, u2_u7_u6_n132, u2_u7_u6_n133, u2_u7_u6_n134, u2_u7_u6_n135, 
       u2_u7_u6_n136, u2_u7_u6_n137, u2_u7_u6_n138, u2_u7_u6_n139, u2_u7_u6_n140, u2_u7_u6_n141, u2_u7_u6_n142, u2_u7_u6_n143, u2_u7_u6_n144, 
       u2_u7_u6_n145, u2_u7_u6_n146, u2_u7_u6_n147, u2_u7_u6_n148, u2_u7_u6_n149, u2_u7_u6_n150, u2_u7_u6_n151, u2_u7_u6_n152, u2_u7_u6_n153, 
       u2_u7_u6_n154, u2_u7_u6_n155, u2_u7_u6_n156, u2_u7_u6_n157, u2_u7_u6_n158, u2_u7_u6_n159, u2_u7_u6_n160, u2_u7_u6_n161, u2_u7_u6_n162, 
       u2_u7_u6_n163, u2_u7_u6_n164, u2_u7_u6_n165, u2_u7_u6_n166, u2_u7_u6_n167, u2_u7_u6_n168, u2_u7_u6_n169, u2_u7_u6_n170, u2_u7_u6_n171, 
       u2_u7_u6_n172, u2_u7_u6_n173, u2_u7_u6_n174, u2_u7_u6_n88, u2_u7_u6_n89, u2_u7_u6_n90, u2_u7_u6_n91, u2_u7_u6_n92, u2_u7_u6_n93, 
       u2_u7_u6_n94, u2_u7_u6_n95, u2_u7_u6_n96, u2_u7_u6_n97, u2_u7_u6_n98, u2_u7_u6_n99, u2_uk_K_r0_0, u2_uk_K_r0_1, u2_uk_K_r0_10, 
       u2_uk_K_r0_11, u2_uk_K_r0_12, u2_uk_K_r0_13, u2_uk_K_r0_14, u2_uk_K_r0_15, u2_uk_K_r0_16, u2_uk_K_r0_17, u2_uk_K_r0_18, u2_uk_K_r0_19, 
       u2_uk_K_r0_2, u2_uk_K_r0_20, u2_uk_K_r0_21, u2_uk_K_r0_22, u2_uk_K_r0_23, u2_uk_K_r0_24, u2_uk_K_r0_25, u2_uk_K_r0_26, u2_uk_K_r0_27, 
       u2_uk_K_r0_28, u2_uk_K_r0_29, u2_uk_K_r0_3, u2_uk_K_r0_30, u2_uk_K_r0_31, u2_uk_K_r0_32, u2_uk_K_r0_33, u2_uk_K_r0_34, u2_uk_K_r0_35, 
       u2_uk_K_r0_36, u2_uk_K_r0_37, u2_uk_K_r0_38, u2_uk_K_r0_39, u2_uk_K_r0_4, u2_uk_K_r0_40, u2_uk_K_r0_41, u2_uk_K_r0_42, u2_uk_K_r0_43, 
       u2_uk_K_r0_44, u2_uk_K_r0_45, u2_uk_K_r0_46, u2_uk_K_r0_47, u2_uk_K_r0_48, u2_uk_K_r0_49, u2_uk_K_r0_5, u2_uk_K_r0_50, u2_uk_K_r0_51, 
       u2_uk_K_r0_52, u2_uk_K_r0_53, u2_uk_K_r0_54, u2_uk_K_r0_55, u2_uk_K_r0_6, u2_uk_K_r0_7, u2_uk_K_r0_8, u2_uk_K_r0_9, u2_uk_K_r10_0, 
       u2_uk_K_r10_1, u2_uk_K_r10_10, u2_uk_K_r10_11, u2_uk_K_r10_12, u2_uk_K_r10_13, u2_uk_K_r10_14, u2_uk_K_r10_15, u2_uk_K_r10_16, u2_uk_K_r10_17, 
       u2_uk_K_r10_18, u2_uk_K_r10_19, u2_uk_K_r10_2, u2_uk_K_r10_20, u2_uk_K_r10_21, u2_uk_K_r10_22, u2_uk_K_r10_23, u2_uk_K_r10_24, u2_uk_K_r10_25, 
       u2_uk_K_r10_26, u2_uk_K_r10_27, u2_uk_K_r10_28, u2_uk_K_r10_29, u2_uk_K_r10_3, u2_uk_K_r10_30, u2_uk_K_r10_31, u2_uk_K_r10_32, u2_uk_K_r10_33, 
       u2_uk_K_r10_34, u2_uk_K_r10_35, u2_uk_K_r10_36, u2_uk_K_r10_37, u2_uk_K_r10_38, u2_uk_K_r10_39, u2_uk_K_r10_4, u2_uk_K_r10_40, u2_uk_K_r10_41, 
       u2_uk_K_r10_42, u2_uk_K_r10_43, u2_uk_K_r10_44, u2_uk_K_r10_45, u2_uk_K_r10_46, u2_uk_K_r10_47, u2_uk_K_r10_48, u2_uk_K_r10_49, u2_uk_K_r10_5, 
       u2_uk_K_r10_50, u2_uk_K_r10_51, u2_uk_K_r10_52, u2_uk_K_r10_53, u2_uk_K_r10_54, u2_uk_K_r10_55, u2_uk_K_r10_6, u2_uk_K_r10_7, u2_uk_K_r10_8, 
       u2_uk_K_r10_9, u2_uk_K_r11_0, u2_uk_K_r11_1, u2_uk_K_r11_10, u2_uk_K_r11_11, u2_uk_K_r11_12, u2_uk_K_r11_13, u2_uk_K_r11_14, u2_uk_K_r11_15, 
       u2_uk_K_r11_16, u2_uk_K_r11_17, u2_uk_K_r11_18, u2_uk_K_r11_19, u2_uk_K_r11_2, u2_uk_K_r11_20, u2_uk_K_r11_21, u2_uk_K_r11_22, u2_uk_K_r11_23, 
       u2_uk_K_r11_24, u2_uk_K_r11_25, u2_uk_K_r11_26, u2_uk_K_r11_27, u2_uk_K_r11_29, u2_uk_K_r11_3, u2_uk_K_r11_30, u2_uk_K_r11_31, u2_uk_K_r11_32, 
       u2_uk_K_r11_33, u2_uk_K_r11_34, u2_uk_K_r11_35, u2_uk_K_r11_36, u2_uk_K_r11_37, u2_uk_K_r11_38, u2_uk_K_r11_39, u2_uk_K_r11_4, u2_uk_K_r11_40, 
       u2_uk_K_r11_41, u2_uk_K_r11_42, u2_uk_K_r11_43, u2_uk_K_r11_44, u2_uk_K_r11_45, u2_uk_K_r11_46, u2_uk_K_r11_47, u2_uk_K_r11_49, u2_uk_K_r11_5, 
       u2_uk_K_r11_50, u2_uk_K_r11_51, u2_uk_K_r11_52, u2_uk_K_r11_54, u2_uk_K_r11_55, u2_uk_K_r11_6, u2_uk_K_r11_7, u2_uk_K_r11_8, u2_uk_K_r11_9, 
       u2_uk_K_r12_0, u2_uk_K_r12_1, u2_uk_K_r12_10, u2_uk_K_r12_11, u2_uk_K_r12_12, u2_uk_K_r12_13, u2_uk_K_r12_14, u2_uk_K_r12_15, u2_uk_K_r12_16, 
       u2_uk_K_r12_17, u2_uk_K_r12_18, u2_uk_K_r12_19, u2_uk_K_r12_2, u2_uk_K_r12_20, u2_uk_K_r12_21, u2_uk_K_r12_22, u2_uk_K_r12_23, u2_uk_K_r12_24, 
       u2_uk_K_r12_25, u2_uk_K_r12_26, u2_uk_K_r12_27, u2_uk_K_r12_28, u2_uk_K_r12_29, u2_uk_K_r12_3, u2_uk_K_r12_30, u2_uk_K_r12_31, u2_uk_K_r12_32, 
       u2_uk_K_r12_33, u2_uk_K_r12_34, u2_uk_K_r12_35, u2_uk_K_r12_36, u2_uk_K_r12_37, u2_uk_K_r12_38, u2_uk_K_r12_39, u2_uk_K_r12_4, u2_uk_K_r12_40, 
       u2_uk_K_r12_41, u2_uk_K_r12_42, u2_uk_K_r12_43, u2_uk_K_r12_44, u2_uk_K_r12_45, u2_uk_K_r12_46, u2_uk_K_r12_47, u2_uk_K_r12_48, u2_uk_K_r12_49, 
       u2_uk_K_r12_5, u2_uk_K_r12_50, u2_uk_K_r12_51, u2_uk_K_r12_52, u2_uk_K_r12_53, u2_uk_K_r12_54, u2_uk_K_r12_55, u2_uk_K_r12_6, u2_uk_K_r12_7, 
       u2_uk_K_r12_8, u2_uk_K_r12_9, u2_uk_K_r13_0, u2_uk_K_r13_1, u2_uk_K_r13_10, u2_uk_K_r13_11, u2_uk_K_r13_12, u2_uk_K_r13_13, u2_uk_K_r13_14, 
       u2_uk_K_r13_15, u2_uk_K_r13_16, u2_uk_K_r13_17, u2_uk_K_r13_18, u2_uk_K_r13_19, u2_uk_K_r13_2, u2_uk_K_r13_20, u2_uk_K_r13_21, u2_uk_K_r13_23, 
       u2_uk_K_r13_24, u2_uk_K_r13_25, u2_uk_K_r13_26, u2_uk_K_r13_27, u2_uk_K_r13_28, u2_uk_K_r13_29, u2_uk_K_r13_3, u2_uk_K_r13_30, u2_uk_K_r13_31, 
       u2_uk_K_r13_33, u2_uk_K_r13_34, u2_uk_K_r13_35, u2_uk_K_r13_36, u2_uk_K_r13_37, u2_uk_K_r13_38, u2_uk_K_r13_39, u2_uk_K_r13_4, u2_uk_K_r13_40, 
       u2_uk_K_r13_41, u2_uk_K_r13_42, u2_uk_K_r13_43, u2_uk_K_r13_44, u2_uk_K_r13_45, u2_uk_K_r13_46, u2_uk_K_r13_47, u2_uk_K_r13_48, u2_uk_K_r13_49, 
       u2_uk_K_r13_5, u2_uk_K_r13_50, u2_uk_K_r13_51, u2_uk_K_r13_52, u2_uk_K_r13_53, u2_uk_K_r13_54, u2_uk_K_r13_55, u2_uk_K_r13_6, u2_uk_K_r13_7, 
       u2_uk_K_r13_8, u2_uk_K_r13_9, u2_uk_K_r14_10, u2_uk_K_r14_11, u2_uk_K_r14_12, u2_uk_K_r14_15, u2_uk_K_r14_16, u2_uk_K_r14_18, u2_uk_K_r14_2, 
       u2_uk_K_r14_23, u2_uk_K_r14_3, u2_uk_K_r14_38, u2_uk_K_r14_39, u2_uk_K_r14_42, u2_uk_K_r14_43, u2_uk_K_r14_45, u2_uk_K_r14_46, u2_uk_K_r14_5, 
       u2_uk_K_r14_50, u2_uk_K_r14_8, u2_uk_K_r14_9, u2_uk_K_r1_0, u2_uk_K_r1_1, u2_uk_K_r1_10, u2_uk_K_r1_11, u2_uk_K_r1_12, u2_uk_K_r1_13, 
       u2_uk_K_r1_14, u2_uk_K_r1_17, u2_uk_K_r1_19, u2_uk_K_r1_2, u2_uk_K_r1_20, u2_uk_K_r1_23, u2_uk_K_r1_24, u2_uk_K_r1_25, u2_uk_K_r1_26, 
       u2_uk_K_r1_27, u2_uk_K_r1_28, u2_uk_K_r1_29, u2_uk_K_r1_3, u2_uk_K_r1_30, u2_uk_K_r1_31, u2_uk_K_r1_32, u2_uk_K_r1_33, u2_uk_K_r1_34, 
       u2_uk_K_r1_35, u2_uk_K_r1_36, u2_uk_K_r1_37, u2_uk_K_r1_38, u2_uk_K_r1_39, u2_uk_K_r1_4, u2_uk_K_r1_40, u2_uk_K_r1_41, u2_uk_K_r1_42, 
       u2_uk_K_r1_43, u2_uk_K_r1_44, u2_uk_K_r1_45, u2_uk_K_r1_46, u2_uk_K_r1_48, u2_uk_K_r1_49, u2_uk_K_r1_5, u2_uk_K_r1_50, u2_uk_K_r1_51, 
       u2_uk_K_r1_52, u2_uk_K_r1_53, u2_uk_K_r1_54, u2_uk_K_r1_55, u2_uk_K_r1_6, u2_uk_K_r1_7, u2_uk_K_r1_8, u2_uk_K_r1_9, u2_uk_K_r2_0, 
       u2_uk_K_r2_1, u2_uk_K_r2_10, u2_uk_K_r2_11, u2_uk_K_r2_12, u2_uk_K_r2_14, u2_uk_K_r2_15, u2_uk_K_r2_16, u2_uk_K_r2_17, u2_uk_K_r2_19, 
       u2_uk_K_r2_2, u2_uk_K_r2_20, u2_uk_K_r2_22, u2_uk_K_r2_23, u2_uk_K_r2_24, u2_uk_K_r2_26, u2_uk_K_r2_29, u2_uk_K_r2_3, u2_uk_K_r2_30, 
       u2_uk_K_r2_32, u2_uk_K_r2_33, u2_uk_K_r2_34, u2_uk_K_r2_35, u2_uk_K_r2_37, u2_uk_K_r2_38, u2_uk_K_r2_39, u2_uk_K_r2_4, u2_uk_K_r2_40, 
       u2_uk_K_r2_41, u2_uk_K_r2_42, u2_uk_K_r2_43, u2_uk_K_r2_44, u2_uk_K_r2_45, u2_uk_K_r2_46, u2_uk_K_r2_47, u2_uk_K_r2_48, u2_uk_K_r2_5, 
       u2_uk_K_r2_50, u2_uk_K_r2_51, u2_uk_K_r2_52, u2_uk_K_r2_53, u2_uk_K_r2_54, u2_uk_K_r2_6, u2_uk_K_r2_7, u2_uk_K_r2_8, u2_uk_K_r2_9, 
       u2_uk_K_r3_0, u2_uk_K_r3_1, u2_uk_K_r3_10, u2_uk_K_r3_12, u2_uk_K_r3_13, u2_uk_K_r3_15, u2_uk_K_r3_16, u2_uk_K_r3_17, u2_uk_K_r3_18, 
       u2_uk_K_r3_2, u2_uk_K_r3_20, u2_uk_K_r3_21, u2_uk_K_r3_22, u2_uk_K_r3_23, u2_uk_K_r3_24, u2_uk_K_r3_25, u2_uk_K_r3_26, u2_uk_K_r3_27, 
       u2_uk_K_r3_28, u2_uk_K_r3_29, u2_uk_K_r3_3, u2_uk_K_r3_30, u2_uk_K_r3_31, u2_uk_K_r3_32, u2_uk_K_r3_33, u2_uk_K_r3_34, u2_uk_K_r3_35, 
       u2_uk_K_r3_36, u2_uk_K_r3_37, u2_uk_K_r3_38, u2_uk_K_r3_39, u2_uk_K_r3_4, u2_uk_K_r3_40, u2_uk_K_r3_41, u2_uk_K_r3_42, u2_uk_K_r3_44, 
       u2_uk_K_r3_45, u2_uk_K_r3_46, u2_uk_K_r3_47, u2_uk_K_r3_48, u2_uk_K_r3_49, u2_uk_K_r3_5, u2_uk_K_r3_50, u2_uk_K_r3_51, u2_uk_K_r3_52, 
       u2_uk_K_r3_53, u2_uk_K_r3_54, u2_uk_K_r3_55, u2_uk_K_r3_6, u2_uk_K_r3_7, u2_uk_K_r3_8, u2_uk_K_r4_0, u2_uk_K_r4_1, u2_uk_K_r4_10, 
       u2_uk_K_r4_12, u2_uk_K_r4_13, u2_uk_K_r4_14, u2_uk_K_r4_15, u2_uk_K_r4_16, u2_uk_K_r4_18, u2_uk_K_r4_19, u2_uk_K_r4_2, u2_uk_K_r4_20, 
       u2_uk_K_r4_21, u2_uk_K_r4_22, u2_uk_K_r4_23, u2_uk_K_r4_24, u2_uk_K_r4_25, u2_uk_K_r4_26, u2_uk_K_r4_27, u2_uk_K_r4_28, u2_uk_K_r4_29, 
       u2_uk_K_r4_3, u2_uk_K_r4_30, u2_uk_K_r4_31, u2_uk_K_r4_32, u2_uk_K_r4_34, u2_uk_K_r4_36, u2_uk_K_r4_37, u2_uk_K_r4_39, u2_uk_K_r4_40, 
       u2_uk_K_r4_41, u2_uk_K_r4_42, u2_uk_K_r4_43, u2_uk_K_r4_44, u2_uk_K_r4_45, u2_uk_K_r4_46, u2_uk_K_r4_47, u2_uk_K_r4_48, u2_uk_K_r4_49, 
       u2_uk_K_r4_50, u2_uk_K_r4_51, u2_uk_K_r4_52, u2_uk_K_r4_53, u2_uk_K_r4_54, u2_uk_K_r4_6, u2_uk_K_r4_7, u2_uk_K_r4_8, u2_uk_K_r4_9, 
       u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_11, u2_uk_K_r5_12, u2_uk_K_r5_13, u2_uk_K_r5_14, u2_uk_K_r5_15, u2_uk_K_r5_16, u2_uk_K_r5_18, 
       u2_uk_K_r5_2, u2_uk_K_r5_20, u2_uk_K_r5_21, u2_uk_K_r5_22, u2_uk_K_r5_23, u2_uk_K_r5_24, u2_uk_K_r5_25, u2_uk_K_r5_26, u2_uk_K_r5_27, 
       u2_uk_K_r5_28, u2_uk_K_r5_29, u2_uk_K_r5_3, u2_uk_K_r5_30, u2_uk_K_r5_31, u2_uk_K_r5_32, u2_uk_K_r5_33, u2_uk_K_r5_34, u2_uk_K_r5_35, 
       u2_uk_K_r5_36, u2_uk_K_r5_37, u2_uk_K_r5_38, u2_uk_K_r5_40, u2_uk_K_r5_42, u2_uk_K_r5_43, u2_uk_K_r5_44, u2_uk_K_r5_45, u2_uk_K_r5_46, 
       u2_uk_K_r5_47, u2_uk_K_r5_48, u2_uk_K_r5_49, u2_uk_K_r5_5, u2_uk_K_r5_50, u2_uk_K_r5_51, u2_uk_K_r5_52, u2_uk_K_r5_53, u2_uk_K_r5_54, 
       u2_uk_K_r5_55, u2_uk_K_r5_6, u2_uk_K_r5_7, u2_uk_K_r5_8, u2_uk_K_r5_9, u2_uk_K_r6_0, u2_uk_K_r6_1, u2_uk_K_r6_10, u2_uk_K_r6_11, 
       u2_uk_K_r6_12, u2_uk_K_r6_13, u2_uk_K_r6_14, u2_uk_K_r6_15, u2_uk_K_r6_16, u2_uk_K_r6_17, u2_uk_K_r6_18, u2_uk_K_r6_19, u2_uk_K_r6_2, 
       u2_uk_K_r6_20, u2_uk_K_r6_21, u2_uk_K_r6_22, u2_uk_K_r6_23, u2_uk_K_r6_24, u2_uk_K_r6_25, u2_uk_K_r6_26, u2_uk_K_r6_27, u2_uk_K_r6_28, 
       u2_uk_K_r6_29, u2_uk_K_r6_3, u2_uk_K_r6_30, u2_uk_K_r6_31, u2_uk_K_r6_32, u2_uk_K_r6_33, u2_uk_K_r6_34, u2_uk_K_r6_35, u2_uk_K_r6_36, 
       u2_uk_K_r6_37, u2_uk_K_r6_38, u2_uk_K_r6_39, u2_uk_K_r6_4, u2_uk_K_r6_40, u2_uk_K_r6_41, u2_uk_K_r6_42, u2_uk_K_r6_43, u2_uk_K_r6_44, 
       u2_uk_K_r6_45, u2_uk_K_r6_46, u2_uk_K_r6_47, u2_uk_K_r6_48, u2_uk_K_r6_49, u2_uk_K_r6_5, u2_uk_K_r6_50, u2_uk_K_r6_51, u2_uk_K_r6_52, 
       u2_uk_K_r6_53, u2_uk_K_r6_54, u2_uk_K_r6_55, u2_uk_K_r6_6, u2_uk_K_r6_7, u2_uk_K_r6_8, u2_uk_K_r6_9, u2_uk_K_r7_1, u2_uk_K_r7_10, 
       u2_uk_K_r7_11, u2_uk_K_r7_12, u2_uk_K_r7_13, u2_uk_K_r7_14, u2_uk_K_r7_15, u2_uk_K_r7_16, u2_uk_K_r7_17, u2_uk_K_r7_18, u2_uk_K_r7_19, 
       u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_21, u2_uk_K_r7_22, u2_uk_K_r7_23, u2_uk_K_r7_24, u2_uk_K_r7_27, u2_uk_K_r7_28, u2_uk_K_r7_29, 
       u2_uk_K_r7_3, u2_uk_K_r7_30, u2_uk_K_r7_31, u2_uk_K_r7_33, u2_uk_K_r7_34, u2_uk_K_r7_35, u2_uk_K_r7_36, u2_uk_K_r7_37, u2_uk_K_r7_38, 
       u2_uk_K_r7_4, u2_uk_K_r7_40, u2_uk_K_r7_42, u2_uk_K_r7_43, u2_uk_K_r7_44, u2_uk_K_r7_45, u2_uk_K_r7_46, u2_uk_K_r7_47, u2_uk_K_r7_49, 
       u2_uk_K_r7_5, u2_uk_K_r7_50, u2_uk_K_r7_51, u2_uk_K_r7_52, u2_uk_K_r7_53, u2_uk_K_r7_54, u2_uk_K_r7_6, u2_uk_K_r7_7, u2_uk_K_r7_8, 
       u2_uk_K_r7_9, u2_uk_K_r8_0, u2_uk_K_r8_1, u2_uk_K_r8_10, u2_uk_K_r8_11, u2_uk_K_r8_12, u2_uk_K_r8_13, u2_uk_K_r8_14, u2_uk_K_r8_15, 
       u2_uk_K_r8_17, u2_uk_K_r8_18, u2_uk_K_r8_19, u2_uk_K_r8_20, u2_uk_K_r8_21, u2_uk_K_r8_23, u2_uk_K_r8_24, u2_uk_K_r8_25, u2_uk_K_r8_26, 
       u2_uk_K_r8_27, u2_uk_K_r8_28, u2_uk_K_r8_29, u2_uk_K_r8_3, u2_uk_K_r8_30, u2_uk_K_r8_31, u2_uk_K_r8_32, u2_uk_K_r8_33, u2_uk_K_r8_34, 
       u2_uk_K_r8_35, u2_uk_K_r8_36, u2_uk_K_r8_38, u2_uk_K_r8_39, u2_uk_K_r8_4, u2_uk_K_r8_40, u2_uk_K_r8_43, u2_uk_K_r8_44, u2_uk_K_r8_45, 
       u2_uk_K_r8_46, u2_uk_K_r8_47, u2_uk_K_r8_48, u2_uk_K_r8_49, u2_uk_K_r8_5, u2_uk_K_r8_50, u2_uk_K_r8_51, u2_uk_K_r8_52, u2_uk_K_r8_53, 
       u2_uk_K_r8_54, u2_uk_K_r8_55, u2_uk_K_r8_6, u2_uk_K_r8_7, u2_uk_K_r8_8, u2_uk_K_r8_9, u2_uk_K_r9_0, u2_uk_K_r9_1, u2_uk_K_r9_11, 
       u2_uk_K_r9_12, u2_uk_K_r9_13, u2_uk_K_r9_14, u2_uk_K_r9_15, u2_uk_K_r9_16, u2_uk_K_r9_17, u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_2, 
       u2_uk_K_r9_20, u2_uk_K_r9_21, u2_uk_K_r9_22, u2_uk_K_r9_23, u2_uk_K_r9_24, u2_uk_K_r9_25, u2_uk_K_r9_26, u2_uk_K_r9_27, u2_uk_K_r9_28, 
       u2_uk_K_r9_29, u2_uk_K_r9_3, u2_uk_K_r9_30, u2_uk_K_r9_31, u2_uk_K_r9_32, u2_uk_K_r9_33, u2_uk_K_r9_34, u2_uk_K_r9_35, u2_uk_K_r9_36, 
       u2_uk_K_r9_37, u2_uk_K_r9_38, u2_uk_K_r9_39, u2_uk_K_r9_40, u2_uk_K_r9_41, u2_uk_K_r9_42, u2_uk_K_r9_43, u2_uk_K_r9_44, u2_uk_K_r9_45, 
       u2_uk_K_r9_46, u2_uk_K_r9_47, u2_uk_K_r9_49, u2_uk_K_r9_5, u2_uk_K_r9_50, u2_uk_K_r9_51, u2_uk_K_r9_52, u2_uk_K_r9_53, u2_uk_K_r9_54, 
       u2_uk_K_r9_55, u2_uk_K_r9_6, u2_uk_K_r9_7, u2_uk_K_r9_8, u2_uk_K_r9_9, u2_uk_n1000, u2_uk_n1001, u2_uk_n1002, u2_uk_n1003, 
       u2_uk_n1005, u2_uk_n1006, u2_uk_n1007, u2_uk_n1009, u2_uk_n1010, u2_uk_n1011, u2_uk_n1012, u2_uk_n1018, u2_uk_n1022, 
       u2_uk_n1025, u2_uk_n1034, u2_uk_n1036, u2_uk_n1039, u2_uk_n1042, u2_uk_n1044, u2_uk_n1045, u2_uk_n1047, u2_uk_n1051, 
       u2_uk_n1055, u2_uk_n1056, u2_uk_n1058, u2_uk_n1061, u2_uk_n1063, u2_uk_n1065, u2_uk_n1067, u2_uk_n1070, u2_uk_n1071, 
       u2_uk_n1073, u2_uk_n1081, u2_uk_n1085, u2_uk_n1087, u2_uk_n1090, u2_uk_n1092, u2_uk_n1094, u2_uk_n1097, u2_uk_n1099, 
       u2_uk_n1100, u2_uk_n1101, u2_uk_n1102, u2_uk_n1103, u2_uk_n1104, u2_uk_n1105, u2_uk_n1106, u2_uk_n1107, u2_uk_n1108, 
       u2_uk_n1109, u2_uk_n1111, u2_uk_n1112, u2_uk_n1114, u2_uk_n1115, u2_uk_n1116, u2_uk_n1119, u2_uk_n1121, u2_uk_n1125, 
       u2_uk_n1129, u2_uk_n1131, u2_uk_n1134, u2_uk_n1135, u2_uk_n1139, u2_uk_n1143, u2_uk_n1144, u2_uk_n1145, u2_uk_n1146, 
       u2_uk_n1148, u2_uk_n1149, u2_uk_n1150, u2_uk_n1153, u2_uk_n1154, u2_uk_n1155, u2_uk_n1157, u2_uk_n1159, u2_uk_n1160, 
       u2_uk_n1161, u2_uk_n1162, u2_uk_n1167, u2_uk_n1168, u2_uk_n1174, u2_uk_n1175, u2_uk_n1178, u2_uk_n1179, u2_uk_n1183, 
       u2_uk_n1184, u2_uk_n1185, u2_uk_n1188, u2_uk_n1189, u2_uk_n1190, u2_uk_n1191, u2_uk_n1192, u2_uk_n1194, u2_uk_n1195, 
       u2_uk_n1197, u2_uk_n1198, u2_uk_n1199, u2_uk_n1200, u2_uk_n1201, u2_uk_n1203, u2_uk_n1204, u2_uk_n1205, u2_uk_n1206, 
       u2_uk_n1207, u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1211, u2_uk_n1212, u2_uk_n1213, u2_uk_n1214, u2_uk_n1215, 
       u2_uk_n1216, u2_uk_n1217, u2_uk_n1218, u2_uk_n1219, u2_uk_n1220, u2_uk_n1221, u2_uk_n1222, u2_uk_n1223, u2_uk_n1225, 
       u2_uk_n1226, u2_uk_n1227, u2_uk_n1228, u2_uk_n1229, u2_uk_n1230, u2_uk_n1231, u2_uk_n1232, u2_uk_n1233, u2_uk_n1234, 
       u2_uk_n1235, u2_uk_n1236, u2_uk_n1237, u2_uk_n1238, u2_uk_n1239, u2_uk_n1240, u2_uk_n1241, u2_uk_n1242, u2_uk_n1243, 
       u2_uk_n1244, u2_uk_n1245, u2_uk_n1246, u2_uk_n1247, u2_uk_n1248, u2_uk_n1249, u2_uk_n1251, u2_uk_n1252, u2_uk_n1254, 
       u2_uk_n1256, u2_uk_n1258, u2_uk_n1259, u2_uk_n1260, u2_uk_n1261, u2_uk_n1262, u2_uk_n1263, u2_uk_n1264, u2_uk_n1265, 
       u2_uk_n1266, u2_uk_n1267, u2_uk_n1269, u2_uk_n1270, u2_uk_n1273, u2_uk_n1274, u2_uk_n1275, u2_uk_n1277, u2_uk_n1278, 
       u2_uk_n1289, u2_uk_n1292, u2_uk_n1294, u2_uk_n1298, u2_uk_n1299, u2_uk_n1303, u2_uk_n1304, u2_uk_n1308, u2_uk_n1309, 
       u2_uk_n1312, u2_uk_n1313, u2_uk_n1315, u2_uk_n1319, u2_uk_n1320, u2_uk_n1321, u2_uk_n1322, u2_uk_n1325, u2_uk_n1327, 
       u2_uk_n1330, u2_uk_n1331, u2_uk_n1335, u2_uk_n1336, u2_uk_n1337, u2_uk_n1342, u2_uk_n1344, u2_uk_n1347, u2_uk_n1348, 
       u2_uk_n1352, u2_uk_n1353, u2_uk_n1360, u2_uk_n1363, u2_uk_n1364, u2_uk_n1365, u2_uk_n1366, u2_uk_n1367, u2_uk_n1368, 
       u2_uk_n1369, u2_uk_n1371, u2_uk_n1372, u2_uk_n1373, u2_uk_n1374, u2_uk_n1376, u2_uk_n1377, u2_uk_n1378, u2_uk_n1379, 
       u2_uk_n1380, u2_uk_n1381, u2_uk_n1383, u2_uk_n1384, u2_uk_n1385, u2_uk_n1387, u2_uk_n1388, u2_uk_n1389, u2_uk_n1392, 
       u2_uk_n1393, u2_uk_n1394, u2_uk_n1395, u2_uk_n1396, u2_uk_n1397, u2_uk_n1399, u2_uk_n1400, u2_uk_n1403, u2_uk_n1406, 
       u2_uk_n1407, u2_uk_n1409, u2_uk_n1411, u2_uk_n1412, u2_uk_n1414, u2_uk_n1416, u2_uk_n1417, u2_uk_n1418, u2_uk_n1419, 
       u2_uk_n1420, u2_uk_n1423, u2_uk_n1424, u2_uk_n1425, u2_uk_n1427, u2_uk_n1429, u2_uk_n1430, u2_uk_n1431, u2_uk_n1432, 
       u2_uk_n1434, u2_uk_n1436, u2_uk_n1442, u2_uk_n1444, u2_uk_n1448, u2_uk_n1452, u2_uk_n1455, u2_uk_n1457, u2_uk_n1460, 
       u2_uk_n1461, u2_uk_n1464, u2_uk_n1468, u2_uk_n1469, u2_uk_n1471, u2_uk_n1474, u2_uk_n1477, u2_uk_n1478, u2_uk_n1484, 
       u2_uk_n1487, u2_uk_n1491, u2_uk_n1498, u2_uk_n1499, u2_uk_n1500, u2_uk_n1501, u2_uk_n1502, u2_uk_n1503, u2_uk_n1504, 
       u2_uk_n1506, u2_uk_n1507, u2_uk_n1508, u2_uk_n1510, u2_uk_n1511, u2_uk_n1513, u2_uk_n1514, u2_uk_n1515, u2_uk_n1517, 
       u2_uk_n1518, u2_uk_n1519, u2_uk_n1521, u2_uk_n1522, u2_uk_n1524, u2_uk_n1525, u2_uk_n1526, u2_uk_n1527, u2_uk_n1528, 
       u2_uk_n1529, u2_uk_n1530, u2_uk_n1531, u2_uk_n1532, u2_uk_n1533, u2_uk_n1534, u2_uk_n1535, u2_uk_n1536, u2_uk_n1537, 
       u2_uk_n1538, u2_uk_n1540, u2_uk_n1541, u2_uk_n1542, u2_uk_n1543, u2_uk_n1547, u2_uk_n1551, u2_uk_n1554, u2_uk_n1558, 
       u2_uk_n1562, u2_uk_n1565, u2_uk_n1569, u2_uk_n1570, u2_uk_n1571, u2_uk_n1574, u2_uk_n1575, u2_uk_n1576, u2_uk_n1577, 
       u2_uk_n1578, u2_uk_n1582, u2_uk_n1583, u2_uk_n1584, u2_uk_n1588, u2_uk_n1589, u2_uk_n1590, u2_uk_n1591, u2_uk_n1593, 
       u2_uk_n1595, u2_uk_n1596, u2_uk_n1597, u2_uk_n1598, u2_uk_n1599, u2_uk_n1600, u2_uk_n1602, u2_uk_n1603, u2_uk_n1604, 
       u2_uk_n1605, u2_uk_n1610, u2_uk_n1611, u2_uk_n1612, u2_uk_n1613, u2_uk_n1614, u2_uk_n1617, u2_uk_n1619, u2_uk_n1621, 
       u2_uk_n1623, u2_uk_n1624, u2_uk_n1625, u2_uk_n1626, u2_uk_n1629, u2_uk_n1630, u2_uk_n1631, u2_uk_n1632, u2_uk_n1633, 
       u2_uk_n1634, u2_uk_n1637, u2_uk_n1639, u2_uk_n1640, u2_uk_n1642, u2_uk_n1643, u2_uk_n1646, u2_uk_n1647, u2_uk_n1648, 
       u2_uk_n1652, u2_uk_n1653, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, u2_uk_n1659, u2_uk_n1660, u2_uk_n1661, u2_uk_n1662, 
       u2_uk_n1663, u2_uk_n1664, u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1669, u2_uk_n1672, u2_uk_n1673, u2_uk_n1674, 
       u2_uk_n1675, u2_uk_n1677, u2_uk_n1678, u2_uk_n1679, u2_uk_n1680, u2_uk_n1681, u2_uk_n1684, u2_uk_n1685, u2_uk_n1686, 
       u2_uk_n1687, u2_uk_n1690, u2_uk_n1691, u2_uk_n1692, u2_uk_n1698, u2_uk_n1699, u2_uk_n1700, u2_uk_n1701, u2_uk_n1702, 
       u2_uk_n1704, u2_uk_n1705, u2_uk_n1706, u2_uk_n1707, u2_uk_n1714, u2_uk_n1715, u2_uk_n1718, u2_uk_n1719, u2_uk_n1722, 
       u2_uk_n1723, u2_uk_n1724, u2_uk_n1725, u2_uk_n1726, u2_uk_n1727, u2_uk_n1728, u2_uk_n1731, u2_uk_n1732, u2_uk_n1733, 
       u2_uk_n1734, u2_uk_n1735, u2_uk_n1736, u2_uk_n1737, u2_uk_n1738, u2_uk_n1739, u2_uk_n1742, u2_uk_n1743, u2_uk_n1744, 
       u2_uk_n1745, u2_uk_n1747, u2_uk_n1750, u2_uk_n1751, u2_uk_n1752, u2_uk_n1753, u2_uk_n1754, u2_uk_n1755, u2_uk_n1757, 
       u2_uk_n1760, u2_uk_n1761, u2_uk_n1762, u2_uk_n1763, u2_uk_n1767, u2_uk_n1768, u2_uk_n1771, u2_uk_n1772, u2_uk_n1773, 
       u2_uk_n1774, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1779, u2_uk_n1780, u2_uk_n1782, u2_uk_n1783, u2_uk_n1784, 
       u2_uk_n1786, u2_uk_n1787, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, u2_uk_n1791, u2_uk_n1792, u2_uk_n1793, u2_uk_n1794, 
       u2_uk_n1796, u2_uk_n1799, u2_uk_n1800, u2_uk_n1801, u2_uk_n1802, u2_uk_n1804, u2_uk_n1805, u2_uk_n1806, u2_uk_n1809, 
       u2_uk_n1810, u2_uk_n1811, u2_uk_n1812, u2_uk_n1813, u2_uk_n1814, u2_uk_n1815, u2_uk_n1818, u2_uk_n1820, u2_uk_n1822, 
       u2_uk_n1823, u2_uk_n1825, u2_uk_n1828, u2_uk_n1829, u2_uk_n1830, u2_uk_n1832, u2_uk_n1833, u2_uk_n1835, u2_uk_n1836, 
       u2_uk_n1837, u2_uk_n1838, u2_uk_n1839, u2_uk_n1842, u2_uk_n1843, u2_uk_n1844, u2_uk_n1845, u2_uk_n1850, u2_uk_n1853, 
       u2_uk_n1854, u2_uk_n1857, u2_uk_n242, u2_uk_n250, u2_uk_n251, u2_uk_n252, u2_uk_n271, u2_uk_n277, u2_uk_n279, 
       u2_uk_n292, u2_uk_n298, u2_uk_n312, u2_uk_n346, u2_uk_n349, u2_uk_n353, u2_uk_n363, u2_uk_n366, u2_uk_n369, 
       u2_uk_n375, u2_uk_n376, u2_uk_n377, u2_uk_n379, u2_uk_n382, u2_uk_n385, u2_uk_n391, u2_uk_n395, u2_uk_n407, 
       u2_uk_n409, u2_uk_n437, u2_uk_n443, u2_uk_n460, u2_uk_n468, u2_uk_n472, u2_uk_n496, u2_uk_n500, u2_uk_n501, 
       u2_uk_n509, u2_uk_n518, u2_uk_n524, u2_uk_n526, u2_uk_n551, u2_uk_n582, u2_uk_n586, u2_uk_n587, u2_uk_n590, 
       u2_uk_n601, u2_uk_n603, u2_uk_n605, u2_uk_n608, u2_uk_n634, u2_uk_n656, u2_uk_n662, u2_uk_n672, u2_uk_n676, 
       u2_uk_n677, u2_uk_n681, u2_uk_n685, u2_uk_n686, u2_uk_n688, u2_uk_n692, u2_uk_n694, u2_uk_n695, u2_uk_n702, 
       u2_uk_n717, u2_uk_n930, u2_uk_n931, u2_uk_n932, u2_uk_n933, u2_uk_n934, u2_uk_n935, u2_uk_n937, u2_uk_n940, 
       u2_uk_n941, u2_uk_n944, u2_uk_n947, u2_uk_n948, u2_uk_n949, u2_uk_n950, u2_uk_n951, u2_uk_n952, u2_uk_n953, 
       u2_uk_n954, u2_uk_n956, u2_uk_n957, u2_uk_n960, u2_uk_n961, u2_uk_n962, u2_uk_n964, u2_uk_n965, u2_uk_n966, 
       u2_uk_n967, u2_uk_n968, u2_uk_n969, u2_uk_n970, u2_uk_n971, u2_uk_n972, u2_uk_n973, u2_uk_n974, u2_uk_n975, 
       u2_uk_n976, u2_uk_n977, u2_uk_n978, u2_uk_n979, u2_uk_n980, u2_uk_n981, u2_uk_n982, u2_uk_n983, u2_uk_n984, 
       u2_uk_n988, u2_uk_n989, u2_uk_n990, u2_uk_n992, u2_uk_n994, u2_uk_n996,  u2_uk_n997;
  OAI22_X1 U172 (.B1( decrypt ) , .ZN( key_a_0 ) , .A2( n112 ) , .A1( n115 ) , .B2( n56 ) );
  INV_X1 U173 (.A( key1[0] ) , .ZN( n56 ) );
  INV_X1 U174 (.A( key3[0] ) , .ZN( n112 ) );
  OAI22_X1 U175 (.B1( decrypt ) , .ZN( key_a_10 ) , .A2( n102 ) , .A1( n114 ) , .B2( n46 ) );
  INV_X1 U176 (.A( key1[10] ) , .ZN( n46 ) );
  INV_X1 U177 (.A( key3[10] ) , .ZN( n102 ) );
  OAI22_X1 U178 (.B1( decrypt ) , .ZN( key_a_11 ) , .A2( n101 ) , .A1( n116 ) , .B2( n45 ) );
  INV_X1 U179 (.A( key1[11] ) , .ZN( n45 ) );
  INV_X1 U180 (.A( key3[11] ) , .ZN( n101 ) );
  OAI22_X1 U181 (.B1( decrypt ) , .ZN( key_a_12 ) , .A2( n100 ) , .A1( n116 ) , .B2( n44 ) );
  INV_X1 U182 (.A( key1[12] ) , .ZN( n44 ) );
  INV_X1 U183 (.A( key3[12] ) , .ZN( n100 ) );
  OAI22_X1 U184 (.B1( decrypt ) , .ZN( key_a_13 ) , .A1( n116 ) , .B2( n43 ) , .A2( n99 ) );
  INV_X1 U185 (.A( key1[13] ) , .ZN( n43 ) );
  INV_X1 U186 (.A( key3[13] ) , .ZN( n99 ) );
  OAI22_X1 U187 (.B1( decrypt ) , .ZN( key_a_14 ) , .A1( n116 ) , .B2( n42 ) , .A2( n98 ) );
  INV_X1 U188 (.A( key1[14] ) , .ZN( n42 ) );
  INV_X1 U189 (.A( key3[14] ) , .ZN( n98 ) );
  OAI22_X1 U190 (.B1( decrypt ) , .ZN( key_a_1 ) , .A2( n111 ) , .A1( n116 ) , .B2( n55 ) );
  INV_X1 U191 (.A( key1[1] ) , .ZN( n55 ) );
  INV_X1 U192 (.A( key3[1] ) , .ZN( n111 ) );
  OAI22_X1 U193 (.B1( decrypt ) , .ZN( key_a_2 ) , .A2( n110 ) , .A1( n115 ) , .B2( n54 ) );
  INV_X1 U194 (.A( key1[2] ) , .ZN( n54 ) );
  INV_X1 U195 (.A( key3[2] ) , .ZN( n110 ) );
  OAI22_X1 U196 (.B1( decrypt ) , .ZN( key_a_3 ) , .A2( n109 ) , .A1( n114 ) , .B2( n53 ) );
  INV_X1 U197 (.A( key1[3] ) , .ZN( n53 ) );
  INV_X1 U198 (.A( key3[3] ) , .ZN( n109 ) );
  OAI22_X1 U199 (.B1( decrypt ) , .ZN( key_a_4 ) , .A2( n108 ) , .A1( n114 ) , .B2( n52 ) );
  INV_X1 U200 (.A( key1[4] ) , .ZN( n52 ) );
  INV_X1 U201 (.A( key3[4] ) , .ZN( n108 ) );
  OAI22_X1 U202 (.B1( decrypt ) , .ZN( key_a_9 ) , .A2( n103 ) , .A1( n115 ) , .B2( n47 ) );
  INV_X1 U203 (.A( key1[9] ) , .ZN( n47 ) );
  INV_X1 U204 (.A( key3[9] ) , .ZN( n103 ) );
  OAI22_X1 U205 (.B1( decrypt ) , .ZN( key_a_15 ) , .A1( n116 ) , .B2( n41 ) , .A2( n97 ) );
  INV_X1 U206 (.A( key1[15] ) , .ZN( n41 ) );
  INV_X1 U207 (.A( key3[15] ) , .ZN( n97 ) );
  OAI22_X1 U208 (.B1( decrypt ) , .ZN( key_a_16 ) , .A1( n116 ) , .B2( n40 ) , .A2( n96 ) );
  INV_X1 U209 (.A( key1[16] ) , .ZN( n40 ) );
  INV_X1 U210 (.A( key3[16] ) , .ZN( n96 ) );
  OAI22_X1 U211 (.B1( decrypt ) , .ZN( key_a_17 ) , .A1( n116 ) , .B2( n39 ) , .A2( n95 ) );
  INV_X1 U212 (.A( key1[17] ) , .ZN( n39 ) );
  INV_X1 U213 (.A( key3[17] ) , .ZN( n95 ) );
  OAI22_X1 U214 (.B1( decrypt ) , .ZN( key_a_18 ) , .A1( n116 ) , .B2( n38 ) , .A2( n94 ) );
  INV_X1 U215 (.A( key1[18] ) , .ZN( n38 ) );
  INV_X1 U216 (.A( key3[18] ) , .ZN( n94 ) );
  OAI22_X1 U217 (.B1( decrypt ) , .ZN( key_a_19 ) , .A1( n116 ) , .B2( n37 ) , .A2( n93 ) );
  INV_X1 U218 (.A( key1[19] ) , .ZN( n37 ) );
  INV_X1 U219 (.A( key3[19] ) , .ZN( n93 ) );
  OAI22_X1 U220 (.B1( decrypt ) , .ZN( key_a_20 ) , .A1( n116 ) , .B2( n36 ) , .A2( n92 ) );
  INV_X1 U221 (.A( key1[20] ) , .ZN( n36 ) );
  INV_X1 U222 (.A( key3[20] ) , .ZN( n92 ) );
  OAI22_X1 U223 (.B1( decrypt ) , .ZN( key_a_21 ) , .A1( n116 ) , .B2( n35 ) , .A2( n91 ) );
  INV_X1 U224 (.A( key1[21] ) , .ZN( n35 ) );
  INV_X1 U225 (.A( key3[21] ) , .ZN( n91 ) );
  OAI22_X1 U226 (.B1( decrypt ) , .ZN( key_a_22 ) , .A1( n116 ) , .B2( n34 ) , .A2( n90 ) );
  INV_X1 U227 (.A( key1[22] ) , .ZN( n34 ) );
  INV_X1 U228 (.A( key3[22] ) , .ZN( n90 ) );
  OAI22_X1 U229 (.B1( decrypt ) , .ZN( key_a_23 ) , .A1( n116 ) , .B2( n33 ) , .A2( n89 ) );
  INV_X1 U230 (.A( key1[23] ) , .ZN( n33 ) );
  INV_X1 U231 (.A( key3[23] ) , .ZN( n89 ) );
  OAI22_X1 U232 (.B1( decrypt ) , .ZN( key_a_24 ) , .A1( n116 ) , .B2( n32 ) , .A2( n88 ) );
  INV_X1 U233 (.A( key1[24] ) , .ZN( n32 ) );
  INV_X1 U234 (.A( key3[24] ) , .ZN( n88 ) );
  OAI22_X1 U235 (.B1( decrypt ) , .ZN( key_a_25 ) , .A1( n116 ) , .B2( n31 ) , .A2( n87 ) );
  INV_X1 U236 (.A( key1[25] ) , .ZN( n31 ) );
  INV_X1 U237 (.A( key3[25] ) , .ZN( n87 ) );
  OAI22_X1 U238 (.B1( decrypt ) , .ZN( key_a_26 ) , .A1( n115 ) , .B2( n30 ) , .A2( n86 ) );
  INV_X1 U239 (.A( key1[26] ) , .ZN( n30 ) );
  INV_X1 U240 (.A( key3[26] ) , .ZN( n86 ) );
  OAI22_X1 U241 (.B1( decrypt ) , .ZN( key_a_27 ) , .A1( n115 ) , .B2( n29 ) , .A2( n85 ) );
  INV_X1 U242 (.A( key1[27] ) , .ZN( n29 ) );
  INV_X1 U243 (.A( key3[27] ) , .ZN( n85 ) );
  OAI22_X1 U244 (.B1( decrypt ) , .ZN( key_a_28 ) , .A1( n115 ) , .B2( n28 ) , .A2( n84 ) );
  INV_X1 U245 (.A( key1[28] ) , .ZN( n28 ) );
  INV_X1 U246 (.A( key3[28] ) , .ZN( n84 ) );
  OAI22_X1 U247 (.B1( decrypt ) , .ZN( key_a_29 ) , .A1( n115 ) , .B2( n27 ) , .A2( n83 ) );
  INV_X1 U248 (.A( key1[29] ) , .ZN( n27 ) );
  INV_X1 U249 (.A( key3[29] ) , .ZN( n83 ) );
  OAI22_X1 U250 (.B1( decrypt ) , .ZN( key_a_30 ) , .A1( n115 ) , .B2( n26 ) , .A2( n82 ) );
  INV_X1 U251 (.A( key1[30] ) , .ZN( n26 ) );
  INV_X1 U252 (.A( key3[30] ) , .ZN( n82 ) );
  OAI22_X1 U253 (.B1( decrypt ) , .ZN( key_a_31 ) , .A1( n115 ) , .B2( n25 ) , .A2( n81 ) );
  INV_X1 U254 (.A( key1[31] ) , .ZN( n25 ) );
  INV_X1 U255 (.A( key3[31] ) , .ZN( n81 ) );
  OAI22_X1 U256 (.B1( decrypt ) , .ZN( key_a_32 ) , .A1( n115 ) , .B2( n24 ) , .A2( n80 ) );
  INV_X1 U257 (.A( key1[32] ) , .ZN( n24 ) );
  INV_X1 U258 (.A( key3[32] ) , .ZN( n80 ) );
  OAI22_X1 U259 (.B1( decrypt ) , .ZN( key_a_33 ) , .A1( n115 ) , .B2( n23 ) , .A2( n79 ) );
  INV_X1 U260 (.A( key1[33] ) , .ZN( n23 ) );
  INV_X1 U261 (.A( key3[33] ) , .ZN( n79 ) );
  OAI22_X1 U262 (.B1( decrypt ) , .ZN( key_a_34 ) , .A1( n115 ) , .B2( n22 ) , .A2( n78 ) );
  INV_X1 U263 (.A( key1[34] ) , .ZN( n22 ) );
  INV_X1 U264 (.A( key3[34] ) , .ZN( n78 ) );
  OAI22_X1 U265 (.B1( decrypt ) , .ZN( key_a_35 ) , .A1( n115 ) , .B2( n21 ) , .A2( n77 ) );
  INV_X1 U266 (.A( key1[35] ) , .ZN( n21 ) );
  INV_X1 U267 (.A( key3[35] ) , .ZN( n77 ) );
  OAI22_X1 U268 (.B1( decrypt ) , .ZN( key_a_36 ) , .A1( n115 ) , .B2( n20 ) , .A2( n76 ) );
  INV_X1 U269 (.A( key1[36] ) , .ZN( n20 ) );
  INV_X1 U270 (.A( key3[36] ) , .ZN( n76 ) );
  OAI22_X1 U271 (.B1( decrypt ) , .ZN( key_a_37 ) , .A1( n115 ) , .B2( n19 ) , .A2( n75 ) );
  INV_X1 U272 (.A( key1[37] ) , .ZN( n19 ) );
  INV_X1 U273 (.A( key3[37] ) , .ZN( n75 ) );
  OAI22_X1 U274 (.B1( decrypt ) , .ZN( key_a_38 ) , .A1( n115 ) , .B2( n18 ) , .A2( n74 ) );
  INV_X1 U275 (.A( key1[38] ) , .ZN( n18 ) );
  INV_X1 U276 (.A( key3[38] ) , .ZN( n74 ) );
  OAI22_X1 U277 (.B1( decrypt ) , .ZN( key_a_39 ) , .A1( n115 ) , .B2( n17 ) , .A2( n73 ) );
  INV_X1 U278 (.A( key1[39] ) , .ZN( n17 ) );
  INV_X1 U279 (.A( key3[39] ) , .ZN( n73 ) );
  OAI22_X1 U280 (.B1( decrypt ) , .ZN( key_a_40 ) , .A1( n114 ) , .B2( n16 ) , .A2( n72 ) );
  INV_X1 U281 (.A( key1[40] ) , .ZN( n16 ) );
  INV_X1 U282 (.A( key3[40] ) , .ZN( n72 ) );
  OAI22_X1 U283 (.B1( decrypt ) , .ZN( key_a_41 ) , .A1( n114 ) , .B2( n15 ) , .A2( n71 ) );
  INV_X1 U284 (.A( key1[41] ) , .ZN( n15 ) );
  INV_X1 U285 (.A( key3[41] ) , .ZN( n71 ) );
  OAI22_X1 U286 (.B1( decrypt ) , .ZN( key_a_42 ) , .A1( n114 ) , .B2( n14 ) , .A2( n70 ) );
  INV_X1 U287 (.A( key1[42] ) , .ZN( n14 ) );
  INV_X1 U288 (.A( key3[42] ) , .ZN( n70 ) );
  OAI22_X1 U289 (.B1( decrypt ) , .ZN( key_a_43 ) , .A1( n114 ) , .B2( n13 ) , .A2( n69 ) );
  INV_X1 U290 (.A( key1[43] ) , .ZN( n13 ) );
  INV_X1 U291 (.A( key3[43] ) , .ZN( n69 ) );
  OAI22_X1 U292 (.B1( decrypt ) , .ZN( key_a_44 ) , .A1( n114 ) , .B2( n12 ) , .A2( n68 ) );
  INV_X1 U293 (.A( key1[44] ) , .ZN( n12 ) );
  INV_X1 U294 (.A( key3[44] ) , .ZN( n68 ) );
  OAI22_X1 U295 (.B1( decrypt ) , .ZN( key_a_45 ) , .B2( n11 ) , .A1( n114 ) , .A2( n67 ) );
  INV_X1 U296 (.A( key1[45] ) , .ZN( n11 ) );
  INV_X1 U297 (.A( key3[45] ) , .ZN( n67 ) );
  OAI22_X1 U298 (.B1( decrypt ) , .ZN( key_a_46 ) , .B2( n10 ) , .A1( n114 ) , .A2( n66 ) );
  INV_X1 U299 (.A( key1[46] ) , .ZN( n10 ) );
  INV_X1 U300 (.A( key3[46] ) , .ZN( n66 ) );
  OAI22_X1 U301 (.B1( decrypt ) , .ZN( key_a_47 ) , .A1( n114 ) , .A2( n65 ) , .B2( n9 ) );
  INV_X1 U302 (.A( key1[47] ) , .ZN( n9 ) );
  INV_X1 U303 (.A( key3[47] ) , .ZN( n65 ) );
  OAI22_X1 U304 (.B1( decrypt ) , .ZN( key_a_48 ) , .A1( n114 ) , .A2( n64 ) , .B2( n8 ) );
  INV_X1 U305 (.A( key1[48] ) , .ZN( n8 ) );
  INV_X1 U306 (.A( key3[48] ) , .ZN( n64 ) );
  OAI22_X1 U307 (.B1( decrypt ) , .ZN( key_a_49 ) , .A1( n114 ) , .A2( n63 ) , .B2( n7 ) );
  INV_X1 U308 (.A( key1[49] ) , .ZN( n7 ) );
  INV_X1 U309 (.A( key3[49] ) , .ZN( n63 ) );
  OAI22_X1 U310 (.B1( decrypt ) , .ZN( key_a_50 ) , .A1( n114 ) , .B2( n6 ) , .A2( n62 ) );
  INV_X1 U311 (.A( key1[50] ) , .ZN( n6 ) );
  INV_X1 U312 (.A( key3[50] ) , .ZN( n62 ) );
  OAI22_X1 U313 (.B1( decrypt ) , .ZN( key_a_51 ) , .A1( n114 ) , .B2( n5 ) , .A2( n61 ) );
  INV_X1 U314 (.A( key1[51] ) , .ZN( n5 ) );
  INV_X1 U315 (.A( key3[51] ) , .ZN( n61 ) );
  OAI22_X1 U316 (.B1( decrypt ) , .ZN( key_a_5 ) , .A2( n107 ) , .A1( n114 ) , .B2( n51 ) );
  INV_X1 U317 (.A( key1[5] ) , .ZN( n51 ) );
  INV_X1 U318 (.A( key3[5] ) , .ZN( n107 ) );
  OAI22_X1 U319 (.B1( decrypt ) , .ZN( key_a_6 ) , .A2( n106 ) , .A1( n114 ) , .B2( n50 ) );
  INV_X1 U320 (.A( key1[6] ) , .ZN( n50 ) );
  INV_X1 U321 (.A( key3[6] ) , .ZN( n106 ) );
  OAI22_X1 U322 (.B1( decrypt ) , .ZN( key_a_7 ) , .A2( n105 ) , .A1( n116 ) , .B2( n49 ) );
  INV_X1 U323 (.A( key1[7] ) , .ZN( n49 ) );
  INV_X1 U324 (.A( key3[7] ) , .ZN( n105 ) );
  OAI22_X1 U325 (.B1( decrypt ) , .ZN( key_a_8 ) , .A2( n104 ) , .A1( n115 ) , .B2( n48 ) );
  INV_X1 U326 (.A( key1[8] ) , .ZN( n48 ) );
  INV_X1 U327 (.A( key3[8] ) , .ZN( n104 ) );
  OAI22_X1 U328 (.B1( decrypt ) , .ZN( key_a_52 ) , .A1( n114 ) , .B2( n4 ) , .A2( n60 ) );
  INV_X1 U329 (.A( key1[52] ) , .ZN( n4 ) );
  INV_X1 U330 (.A( key3[52] ) , .ZN( n60 ) );
  OAI22_X1 U331 (.B1( decrypt ) , .ZN( key_a_53 ) , .A1( n114 ) , .B2( n3 ) , .A2( n59 ) );
  INV_X1 U332 (.A( key1[53] ) , .ZN( n3 ) );
  INV_X1 U333 (.A( key3[53] ) , .ZN( n59 ) );
  OAI22_X1 U334 (.B1( decrypt ) , .ZN( key_a_54 ) , .A1( n114 ) , .B2( n2 ) , .A2( n58 ) );
  INV_X1 U335 (.A( key1[54] ) , .ZN( n2 ) );
  INV_X1 U336 (.A( key3[54] ) , .ZN( n58 ) );
  OAI22_X1 U337 (.B1( decrypt ) , .ZN( key_a_55 ) , .B2( n1 ) , .A1( n116 ) , .A2( n57 ) );
  INV_X1 U338 (.A( key1[55] ) , .ZN( n1 ) );
  INV_X1 U339 (.A( key3[55] ) , .ZN( n57 ) );
  INV_X1 U340 (.A( decrypt ) , .ZN( n116 ) );
  INV_X1 U341 (.A( decrypt ) , .ZN( n115 ) );
  INV_X1 U342 (.A( decrypt ) , .ZN( n114 ) );
  DFF_X1 key_b_r_reg_0_0 (.CK( clk ) , .D( key2[0] ) , .Q( key_b_r_0_0 ) );
  DFF_X1 key_b_r_reg_0_1 (.CK( clk ) , .D( key2[1] ) , .Q( key_b_r_0_1 ) );
  DFF_X1 key_b_r_reg_0_10 (.CK( clk ) , .D( key2[10] ) , .Q( key_b_r_0_10 ) );
  DFF_X1 key_b_r_reg_0_11 (.CK( clk ) , .D( key2[11] ) , .Q( key_b_r_0_11 ) );
  DFF_X1 key_b_r_reg_0_12 (.CK( clk ) , .D( key2[12] ) , .Q( key_b_r_0_12 ) );
  DFF_X1 key_b_r_reg_0_13 (.CK( clk ) , .D( key2[13] ) , .Q( key_b_r_0_13 ) );
  DFF_X1 key_b_r_reg_0_14 (.CK( clk ) , .D( key2[14] ) , .Q( key_b_r_0_14 ) );
  DFF_X1 key_b_r_reg_0_15 (.CK( clk ) , .D( key2[15] ) , .Q( key_b_r_0_15 ) );
  DFF_X1 key_b_r_reg_0_16 (.CK( clk ) , .D( key2[16] ) , .Q( key_b_r_0_16 ) );
  DFF_X1 key_b_r_reg_0_17 (.CK( clk ) , .D( key2[17] ) , .Q( key_b_r_0_17 ) );
  DFF_X1 key_b_r_reg_0_18 (.CK( clk ) , .D( key2[18] ) , .Q( key_b_r_0_18 ) );
  DFF_X1 key_b_r_reg_0_19 (.CK( clk ) , .D( key2[19] ) , .Q( key_b_r_0_19 ) );
  DFF_X1 key_b_r_reg_0_2 (.CK( clk ) , .D( key2[2] ) , .Q( key_b_r_0_2 ) );
  DFF_X1 key_b_r_reg_0_20 (.CK( clk ) , .D( key2[20] ) , .Q( key_b_r_0_20 ) );
  DFF_X1 key_b_r_reg_0_21 (.CK( clk ) , .D( key2[21] ) , .Q( key_b_r_0_21 ) );
  DFF_X1 key_b_r_reg_0_22 (.CK( clk ) , .D( key2[22] ) , .Q( key_b_r_0_22 ) );
  DFF_X1 key_b_r_reg_0_23 (.CK( clk ) , .D( key2[23] ) , .Q( key_b_r_0_23 ) );
  DFF_X1 key_b_r_reg_0_24 (.CK( clk ) , .D( key2[24] ) , .Q( key_b_r_0_24 ) );
  DFF_X1 key_b_r_reg_0_25 (.CK( clk ) , .D( key2[25] ) , .Q( key_b_r_0_25 ) );
  DFF_X1 key_b_r_reg_0_26 (.CK( clk ) , .D( key2[26] ) , .Q( key_b_r_0_26 ) );
  DFF_X1 key_b_r_reg_0_27 (.CK( clk ) , .D( key2[27] ) , .Q( key_b_r_0_27 ) );
  DFF_X1 key_b_r_reg_0_28 (.CK( clk ) , .D( key2[28] ) , .Q( key_b_r_0_28 ) );
  DFF_X1 key_b_r_reg_0_29 (.CK( clk ) , .D( key2[29] ) , .Q( key_b_r_0_29 ) );
  DFF_X1 key_b_r_reg_0_3 (.CK( clk ) , .D( key2[3] ) , .Q( key_b_r_0_3 ) );
  DFF_X1 key_b_r_reg_0_30 (.CK( clk ) , .D( key2[30] ) , .Q( key_b_r_0_30 ) );
  DFF_X1 key_b_r_reg_0_31 (.CK( clk ) , .D( key2[31] ) , .Q( key_b_r_0_31 ) );
  DFF_X1 key_b_r_reg_0_32 (.CK( clk ) , .D( key2[32] ) , .Q( key_b_r_0_32 ) );
  DFF_X1 key_b_r_reg_0_33 (.CK( clk ) , .D( key2[33] ) , .Q( key_b_r_0_33 ) );
  DFF_X1 key_b_r_reg_0_34 (.CK( clk ) , .D( key2[34] ) , .Q( key_b_r_0_34 ) );
  DFF_X1 key_b_r_reg_0_35 (.CK( clk ) , .D( key2[35] ) , .Q( key_b_r_0_35 ) );
  DFF_X1 key_b_r_reg_0_36 (.CK( clk ) , .D( key2[36] ) , .Q( key_b_r_0_36 ) );
  DFF_X1 key_b_r_reg_0_37 (.CK( clk ) , .D( key2[37] ) , .Q( key_b_r_0_37 ) );
  DFF_X1 key_b_r_reg_0_38 (.CK( clk ) , .D( key2[38] ) , .Q( key_b_r_0_38 ) );
  DFF_X1 key_b_r_reg_0_39 (.CK( clk ) , .D( key2[39] ) , .Q( key_b_r_0_39 ) );
  DFF_X1 key_b_r_reg_0_4 (.CK( clk ) , .D( key2[4] ) , .Q( key_b_r_0_4 ) );
  DFF_X1 key_b_r_reg_0_40 (.CK( clk ) , .D( key2[40] ) , .Q( key_b_r_0_40 ) );
  DFF_X1 key_b_r_reg_0_41 (.CK( clk ) , .D( key2[41] ) , .Q( key_b_r_0_41 ) );
  DFF_X1 key_b_r_reg_0_42 (.CK( clk ) , .D( key2[42] ) , .Q( key_b_r_0_42 ) );
  DFF_X1 key_b_r_reg_0_43 (.CK( clk ) , .D( key2[43] ) , .Q( key_b_r_0_43 ) );
  DFF_X1 key_b_r_reg_0_44 (.CK( clk ) , .D( key2[44] ) , .Q( key_b_r_0_44 ) );
  DFF_X1 key_b_r_reg_0_45 (.CK( clk ) , .D( key2[45] ) , .Q( key_b_r_0_45 ) );
  DFF_X1 key_b_r_reg_0_46 (.CK( clk ) , .D( key2[46] ) , .Q( key_b_r_0_46 ) );
  DFF_X1 key_b_r_reg_0_47 (.CK( clk ) , .D( key2[47] ) , .Q( key_b_r_0_47 ) );
  DFF_X1 key_b_r_reg_0_48 (.CK( clk ) , .D( key2[48] ) , .Q( key_b_r_0_48 ) );
  DFF_X1 key_b_r_reg_0_49 (.CK( clk ) , .D( key2[49] ) , .Q( key_b_r_0_49 ) );
  DFF_X1 key_b_r_reg_0_5 (.CK( clk ) , .D( key2[5] ) , .Q( key_b_r_0_5 ) );
  DFF_X1 key_b_r_reg_0_50 (.CK( clk ) , .D( key2[50] ) , .Q( key_b_r_0_50 ) );
  DFF_X1 key_b_r_reg_0_51 (.CK( clk ) , .D( key2[51] ) , .Q( key_b_r_0_51 ) );
  DFF_X1 key_b_r_reg_0_52 (.CK( clk ) , .D( key2[52] ) , .Q( key_b_r_0_52 ) );
  DFF_X1 key_b_r_reg_0_53 (.CK( clk ) , .D( key2[53] ) , .Q( key_b_r_0_53 ) );
  DFF_X1 key_b_r_reg_0_54 (.CK( clk ) , .D( key2[54] ) , .Q( key_b_r_0_54 ) );
  DFF_X1 key_b_r_reg_0_55 (.CK( clk ) , .D( key2[55] ) , .Q( key_b_r_0_55 ) );
  DFF_X1 key_b_r_reg_0_6 (.CK( clk ) , .D( key2[6] ) , .Q( key_b_r_0_6 ) );
  DFF_X1 key_b_r_reg_0_7 (.CK( clk ) , .D( key2[7] ) , .Q( key_b_r_0_7 ) );
  DFF_X1 key_b_r_reg_0_8 (.CK( clk ) , .D( key2[8] ) , .Q( key_b_r_0_8 ) );
  DFF_X1 key_b_r_reg_0_9 (.CK( clk ) , .D( key2[9] ) , .Q( key_b_r_0_9 ) );
  DFF_X1 key_b_r_reg_10_0 (.CK( clk ) , .Q( key_b_r_10_0 ) , .D( key_b_r_9_0 ) );
  DFF_X1 key_b_r_reg_10_1 (.CK( clk ) , .Q( key_b_r_10_1 ) , .D( key_b_r_9_1 ) );
  DFF_X1 key_b_r_reg_10_10 (.CK( clk ) , .Q( key_b_r_10_10 ) , .D( key_b_r_9_10 ) );
  DFF_X1 key_b_r_reg_10_11 (.CK( clk ) , .Q( key_b_r_10_11 ) , .D( key_b_r_9_11 ) );
  DFF_X1 key_b_r_reg_10_12 (.CK( clk ) , .Q( key_b_r_10_12 ) , .D( key_b_r_9_12 ) );
  DFF_X1 key_b_r_reg_10_13 (.CK( clk ) , .Q( key_b_r_10_13 ) , .D( key_b_r_9_13 ) );
  DFF_X1 key_b_r_reg_10_14 (.CK( clk ) , .Q( key_b_r_10_14 ) , .D( key_b_r_9_14 ) );
  DFF_X1 key_b_r_reg_10_15 (.CK( clk ) , .Q( key_b_r_10_15 ) , .D( key_b_r_9_15 ) );
  DFF_X1 key_b_r_reg_10_16 (.CK( clk ) , .Q( key_b_r_10_16 ) , .D( key_b_r_9_16 ) );
  DFF_X1 key_b_r_reg_10_17 (.CK( clk ) , .Q( key_b_r_10_17 ) , .D( key_b_r_9_17 ) );
  DFF_X1 key_b_r_reg_10_18 (.CK( clk ) , .Q( key_b_r_10_18 ) , .D( key_b_r_9_18 ) );
  DFF_X1 key_b_r_reg_10_19 (.CK( clk ) , .Q( key_b_r_10_19 ) , .D( key_b_r_9_19 ) );
  DFF_X1 key_b_r_reg_10_2 (.CK( clk ) , .Q( key_b_r_10_2 ) , .D( key_b_r_9_2 ) );
  DFF_X1 key_b_r_reg_10_20 (.CK( clk ) , .Q( key_b_r_10_20 ) , .D( key_b_r_9_20 ) );
  DFF_X1 key_b_r_reg_10_21 (.CK( clk ) , .Q( key_b_r_10_21 ) , .D( key_b_r_9_21 ) );
  DFF_X1 key_b_r_reg_10_22 (.CK( clk ) , .Q( key_b_r_10_22 ) , .D( key_b_r_9_22 ) );
  DFF_X1 key_b_r_reg_10_23 (.CK( clk ) , .Q( key_b_r_10_23 ) , .D( key_b_r_9_23 ) );
  DFF_X1 key_b_r_reg_10_24 (.CK( clk ) , .Q( key_b_r_10_24 ) , .D( key_b_r_9_24 ) );
  DFF_X1 key_b_r_reg_10_25 (.CK( clk ) , .Q( key_b_r_10_25 ) , .D( key_b_r_9_25 ) );
  DFF_X1 key_b_r_reg_10_26 (.CK( clk ) , .Q( key_b_r_10_26 ) , .D( key_b_r_9_26 ) );
  DFF_X1 key_b_r_reg_10_27 (.CK( clk ) , .Q( key_b_r_10_27 ) , .D( key_b_r_9_27 ) );
  DFF_X1 key_b_r_reg_10_28 (.CK( clk ) , .Q( key_b_r_10_28 ) , .D( key_b_r_9_28 ) );
  DFF_X1 key_b_r_reg_10_29 (.CK( clk ) , .Q( key_b_r_10_29 ) , .D( key_b_r_9_29 ) );
  DFF_X1 key_b_r_reg_10_3 (.CK( clk ) , .Q( key_b_r_10_3 ) , .D( key_b_r_9_3 ) );
  DFF_X1 key_b_r_reg_10_30 (.CK( clk ) , .Q( key_b_r_10_30 ) , .D( key_b_r_9_30 ) );
  DFF_X1 key_b_r_reg_10_31 (.CK( clk ) , .Q( key_b_r_10_31 ) , .D( key_b_r_9_31 ) );
  DFF_X1 key_b_r_reg_10_32 (.CK( clk ) , .Q( key_b_r_10_32 ) , .D( key_b_r_9_32 ) );
  DFF_X1 key_b_r_reg_10_33 (.CK( clk ) , .Q( key_b_r_10_33 ) , .D( key_b_r_9_33 ) );
  DFF_X1 key_b_r_reg_10_34 (.CK( clk ) , .Q( key_b_r_10_34 ) , .D( key_b_r_9_34 ) );
  DFF_X1 key_b_r_reg_10_35 (.CK( clk ) , .Q( key_b_r_10_35 ) , .D( key_b_r_9_35 ) );
  DFF_X1 key_b_r_reg_10_36 (.CK( clk ) , .Q( key_b_r_10_36 ) , .D( key_b_r_9_36 ) );
  DFF_X1 key_b_r_reg_10_37 (.CK( clk ) , .Q( key_b_r_10_37 ) , .D( key_b_r_9_37 ) );
  DFF_X1 key_b_r_reg_10_38 (.CK( clk ) , .Q( key_b_r_10_38 ) , .D( key_b_r_9_38 ) );
  DFF_X1 key_b_r_reg_10_39 (.CK( clk ) , .Q( key_b_r_10_39 ) , .D( key_b_r_9_39 ) );
  DFF_X1 key_b_r_reg_10_4 (.CK( clk ) , .Q( key_b_r_10_4 ) , .D( key_b_r_9_4 ) );
  DFF_X1 key_b_r_reg_10_40 (.CK( clk ) , .Q( key_b_r_10_40 ) , .D( key_b_r_9_40 ) );
  DFF_X1 key_b_r_reg_10_41 (.CK( clk ) , .Q( key_b_r_10_41 ) , .D( key_b_r_9_41 ) );
  DFF_X1 key_b_r_reg_10_42 (.CK( clk ) , .Q( key_b_r_10_42 ) , .D( key_b_r_9_42 ) );
  DFF_X1 key_b_r_reg_10_43 (.CK( clk ) , .Q( key_b_r_10_43 ) , .D( key_b_r_9_43 ) );
  DFF_X1 key_b_r_reg_10_44 (.CK( clk ) , .Q( key_b_r_10_44 ) , .D( key_b_r_9_44 ) );
  DFF_X1 key_b_r_reg_10_45 (.CK( clk ) , .Q( key_b_r_10_45 ) , .D( key_b_r_9_45 ) );
  DFF_X1 key_b_r_reg_10_46 (.CK( clk ) , .Q( key_b_r_10_46 ) , .D( key_b_r_9_46 ) );
  DFF_X1 key_b_r_reg_10_47 (.CK( clk ) , .Q( key_b_r_10_47 ) , .D( key_b_r_9_47 ) );
  DFF_X1 key_b_r_reg_10_48 (.CK( clk ) , .Q( key_b_r_10_48 ) , .D( key_b_r_9_48 ) );
  DFF_X1 key_b_r_reg_10_49 (.CK( clk ) , .Q( key_b_r_10_49 ) , .D( key_b_r_9_49 ) );
  DFF_X1 key_b_r_reg_10_5 (.CK( clk ) , .Q( key_b_r_10_5 ) , .D( key_b_r_9_5 ) );
  DFF_X1 key_b_r_reg_10_50 (.CK( clk ) , .Q( key_b_r_10_50 ) , .D( key_b_r_9_50 ) );
  DFF_X1 key_b_r_reg_10_51 (.CK( clk ) , .Q( key_b_r_10_51 ) , .D( key_b_r_9_51 ) );
  DFF_X1 key_b_r_reg_10_52 (.CK( clk ) , .Q( key_b_r_10_52 ) , .D( key_b_r_9_52 ) );
  DFF_X1 key_b_r_reg_10_53 (.CK( clk ) , .Q( key_b_r_10_53 ) , .D( key_b_r_9_53 ) );
  DFF_X1 key_b_r_reg_10_54 (.CK( clk ) , .Q( key_b_r_10_54 ) , .D( key_b_r_9_54 ) );
  DFF_X1 key_b_r_reg_10_55 (.CK( clk ) , .Q( key_b_r_10_55 ) , .D( key_b_r_9_55 ) );
  DFF_X1 key_b_r_reg_10_6 (.CK( clk ) , .Q( key_b_r_10_6 ) , .D( key_b_r_9_6 ) );
  DFF_X1 key_b_r_reg_10_7 (.CK( clk ) , .Q( key_b_r_10_7 ) , .D( key_b_r_9_7 ) );
  DFF_X1 key_b_r_reg_10_8 (.CK( clk ) , .Q( key_b_r_10_8 ) , .D( key_b_r_9_8 ) );
  DFF_X1 key_b_r_reg_10_9 (.CK( clk ) , .Q( key_b_r_10_9 ) , .D( key_b_r_9_9 ) );
  DFF_X1 key_b_r_reg_11_0 (.CK( clk ) , .D( key_b_r_10_0 ) , .Q( key_b_r_11_0 ) );
  DFF_X1 key_b_r_reg_11_1 (.CK( clk ) , .D( key_b_r_10_1 ) , .Q( key_b_r_11_1 ) );
  DFF_X1 key_b_r_reg_11_10 (.CK( clk ) , .D( key_b_r_10_10 ) , .Q( key_b_r_11_10 ) );
  DFF_X1 key_b_r_reg_11_11 (.CK( clk ) , .D( key_b_r_10_11 ) , .Q( key_b_r_11_11 ) );
  DFF_X1 key_b_r_reg_11_12 (.CK( clk ) , .D( key_b_r_10_12 ) , .Q( key_b_r_11_12 ) );
  DFF_X1 key_b_r_reg_11_13 (.CK( clk ) , .D( key_b_r_10_13 ) , .Q( key_b_r_11_13 ) );
  DFF_X1 key_b_r_reg_11_14 (.CK( clk ) , .D( key_b_r_10_14 ) , .Q( key_b_r_11_14 ) );
  DFF_X1 key_b_r_reg_11_15 (.CK( clk ) , .D( key_b_r_10_15 ) , .Q( key_b_r_11_15 ) );
  DFF_X1 key_b_r_reg_11_16 (.CK( clk ) , .D( key_b_r_10_16 ) , .Q( key_b_r_11_16 ) );
  DFF_X1 key_b_r_reg_11_17 (.CK( clk ) , .D( key_b_r_10_17 ) , .Q( key_b_r_11_17 ) );
  DFF_X1 key_b_r_reg_11_18 (.CK( clk ) , .D( key_b_r_10_18 ) , .Q( key_b_r_11_18 ) );
  DFF_X1 key_b_r_reg_11_19 (.CK( clk ) , .D( key_b_r_10_19 ) , .Q( key_b_r_11_19 ) );
  DFF_X1 key_b_r_reg_11_2 (.CK( clk ) , .D( key_b_r_10_2 ) , .Q( key_b_r_11_2 ) );
  DFF_X1 key_b_r_reg_11_20 (.CK( clk ) , .D( key_b_r_10_20 ) , .Q( key_b_r_11_20 ) );
  DFF_X1 key_b_r_reg_11_21 (.CK( clk ) , .D( key_b_r_10_21 ) , .Q( key_b_r_11_21 ) );
  DFF_X1 key_b_r_reg_11_22 (.CK( clk ) , .D( key_b_r_10_22 ) , .Q( key_b_r_11_22 ) );
  DFF_X1 key_b_r_reg_11_23 (.CK( clk ) , .D( key_b_r_10_23 ) , .Q( key_b_r_11_23 ) );
  DFF_X1 key_b_r_reg_11_24 (.CK( clk ) , .D( key_b_r_10_24 ) , .Q( key_b_r_11_24 ) );
  DFF_X1 key_b_r_reg_11_25 (.CK( clk ) , .D( key_b_r_10_25 ) , .Q( key_b_r_11_25 ) );
  DFF_X1 key_b_r_reg_11_26 (.CK( clk ) , .D( key_b_r_10_26 ) , .Q( key_b_r_11_26 ) );
  DFF_X1 key_b_r_reg_11_27 (.CK( clk ) , .D( key_b_r_10_27 ) , .Q( key_b_r_11_27 ) );
  DFF_X1 key_b_r_reg_11_28 (.CK( clk ) , .D( key_b_r_10_28 ) , .Q( key_b_r_11_28 ) );
  DFF_X1 key_b_r_reg_11_29 (.CK( clk ) , .D( key_b_r_10_29 ) , .Q( key_b_r_11_29 ) );
  DFF_X1 key_b_r_reg_11_3 (.CK( clk ) , .D( key_b_r_10_3 ) , .Q( key_b_r_11_3 ) );
  DFF_X1 key_b_r_reg_11_30 (.CK( clk ) , .D( key_b_r_10_30 ) , .Q( key_b_r_11_30 ) );
  DFF_X1 key_b_r_reg_11_31 (.CK( clk ) , .D( key_b_r_10_31 ) , .Q( key_b_r_11_31 ) );
  DFF_X1 key_b_r_reg_11_32 (.CK( clk ) , .D( key_b_r_10_32 ) , .Q( key_b_r_11_32 ) );
  DFF_X1 key_b_r_reg_11_33 (.CK( clk ) , .D( key_b_r_10_33 ) , .Q( key_b_r_11_33 ) );
  DFF_X1 key_b_r_reg_11_34 (.CK( clk ) , .D( key_b_r_10_34 ) , .Q( key_b_r_11_34 ) );
  DFF_X1 key_b_r_reg_11_35 (.CK( clk ) , .D( key_b_r_10_35 ) , .Q( key_b_r_11_35 ) );
  DFF_X1 key_b_r_reg_11_36 (.CK( clk ) , .D( key_b_r_10_36 ) , .Q( key_b_r_11_36 ) );
  DFF_X1 key_b_r_reg_11_37 (.CK( clk ) , .D( key_b_r_10_37 ) , .Q( key_b_r_11_37 ) );
  DFF_X1 key_b_r_reg_11_38 (.CK( clk ) , .D( key_b_r_10_38 ) , .Q( key_b_r_11_38 ) );
  DFF_X1 key_b_r_reg_11_39 (.CK( clk ) , .D( key_b_r_10_39 ) , .Q( key_b_r_11_39 ) );
  DFF_X1 key_b_r_reg_11_4 (.CK( clk ) , .D( key_b_r_10_4 ) , .Q( key_b_r_11_4 ) );
  DFF_X1 key_b_r_reg_11_40 (.CK( clk ) , .D( key_b_r_10_40 ) , .Q( key_b_r_11_40 ) );
  DFF_X1 key_b_r_reg_11_41 (.CK( clk ) , .D( key_b_r_10_41 ) , .Q( key_b_r_11_41 ) );
  DFF_X1 key_b_r_reg_11_42 (.CK( clk ) , .D( key_b_r_10_42 ) , .Q( key_b_r_11_42 ) );
  DFF_X1 key_b_r_reg_11_43 (.CK( clk ) , .D( key_b_r_10_43 ) , .Q( key_b_r_11_43 ) );
  DFF_X1 key_b_r_reg_11_44 (.CK( clk ) , .D( key_b_r_10_44 ) , .Q( key_b_r_11_44 ) );
  DFF_X1 key_b_r_reg_11_45 (.CK( clk ) , .D( key_b_r_10_45 ) , .Q( key_b_r_11_45 ) );
  DFF_X1 key_b_r_reg_11_46 (.CK( clk ) , .D( key_b_r_10_46 ) , .Q( key_b_r_11_46 ) );
  DFF_X1 key_b_r_reg_11_47 (.CK( clk ) , .D( key_b_r_10_47 ) , .Q( key_b_r_11_47 ) );
  DFF_X1 key_b_r_reg_11_48 (.CK( clk ) , .D( key_b_r_10_48 ) , .Q( key_b_r_11_48 ) );
  DFF_X1 key_b_r_reg_11_49 (.CK( clk ) , .D( key_b_r_10_49 ) , .Q( key_b_r_11_49 ) );
  DFF_X1 key_b_r_reg_11_5 (.CK( clk ) , .D( key_b_r_10_5 ) , .Q( key_b_r_11_5 ) );
  DFF_X1 key_b_r_reg_11_50 (.CK( clk ) , .D( key_b_r_10_50 ) , .Q( key_b_r_11_50 ) );
  DFF_X1 key_b_r_reg_11_51 (.CK( clk ) , .D( key_b_r_10_51 ) , .Q( key_b_r_11_51 ) );
  DFF_X1 key_b_r_reg_11_52 (.CK( clk ) , .D( key_b_r_10_52 ) , .Q( key_b_r_11_52 ) );
  DFF_X1 key_b_r_reg_11_53 (.CK( clk ) , .D( key_b_r_10_53 ) , .Q( key_b_r_11_53 ) );
  DFF_X1 key_b_r_reg_11_54 (.CK( clk ) , .D( key_b_r_10_54 ) , .Q( key_b_r_11_54 ) );
  DFF_X1 key_b_r_reg_11_55 (.CK( clk ) , .D( key_b_r_10_55 ) , .Q( key_b_r_11_55 ) );
  DFF_X1 key_b_r_reg_11_6 (.CK( clk ) , .D( key_b_r_10_6 ) , .Q( key_b_r_11_6 ) );
  DFF_X1 key_b_r_reg_11_7 (.CK( clk ) , .D( key_b_r_10_7 ) , .Q( key_b_r_11_7 ) );
  DFF_X1 key_b_r_reg_11_8 (.CK( clk ) , .D( key_b_r_10_8 ) , .Q( key_b_r_11_8 ) );
  DFF_X1 key_b_r_reg_11_9 (.CK( clk ) , .D( key_b_r_10_9 ) , .Q( key_b_r_11_9 ) );
  DFF_X1 key_b_r_reg_12_0 (.CK( clk ) , .D( key_b_r_11_0 ) , .Q( key_b_r_12_0 ) );
  DFF_X1 key_b_r_reg_12_1 (.CK( clk ) , .D( key_b_r_11_1 ) , .Q( key_b_r_12_1 ) );
  DFF_X1 key_b_r_reg_12_10 (.CK( clk ) , .D( key_b_r_11_10 ) , .Q( key_b_r_12_10 ) );
  DFF_X1 key_b_r_reg_12_11 (.CK( clk ) , .D( key_b_r_11_11 ) , .Q( key_b_r_12_11 ) );
  DFF_X1 key_b_r_reg_12_12 (.CK( clk ) , .D( key_b_r_11_12 ) , .Q( key_b_r_12_12 ) );
  DFF_X1 key_b_r_reg_12_13 (.CK( clk ) , .D( key_b_r_11_13 ) , .Q( key_b_r_12_13 ) );
  DFF_X1 key_b_r_reg_12_14 (.CK( clk ) , .D( key_b_r_11_14 ) , .Q( key_b_r_12_14 ) );
  DFF_X1 key_b_r_reg_12_15 (.CK( clk ) , .D( key_b_r_11_15 ) , .Q( key_b_r_12_15 ) );
  DFF_X1 key_b_r_reg_12_16 (.CK( clk ) , .D( key_b_r_11_16 ) , .Q( key_b_r_12_16 ) );
  DFF_X1 key_b_r_reg_12_17 (.CK( clk ) , .D( key_b_r_11_17 ) , .Q( key_b_r_12_17 ) );
  DFF_X1 key_b_r_reg_12_18 (.CK( clk ) , .D( key_b_r_11_18 ) , .Q( key_b_r_12_18 ) );
  DFF_X1 key_b_r_reg_12_19 (.CK( clk ) , .D( key_b_r_11_19 ) , .Q( key_b_r_12_19 ) );
  DFF_X1 key_b_r_reg_12_2 (.CK( clk ) , .D( key_b_r_11_2 ) , .Q( key_b_r_12_2 ) );
  DFF_X1 key_b_r_reg_12_20 (.CK( clk ) , .D( key_b_r_11_20 ) , .Q( key_b_r_12_20 ) );
  DFF_X1 key_b_r_reg_12_21 (.CK( clk ) , .D( key_b_r_11_21 ) , .Q( key_b_r_12_21 ) );
  DFF_X1 key_b_r_reg_12_22 (.CK( clk ) , .D( key_b_r_11_22 ) , .Q( key_b_r_12_22 ) );
  DFF_X1 key_b_r_reg_12_23 (.CK( clk ) , .D( key_b_r_11_23 ) , .Q( key_b_r_12_23 ) );
  DFF_X1 key_b_r_reg_12_24 (.CK( clk ) , .D( key_b_r_11_24 ) , .Q( key_b_r_12_24 ) );
  DFF_X1 key_b_r_reg_12_25 (.CK( clk ) , .D( key_b_r_11_25 ) , .Q( key_b_r_12_25 ) );
  DFF_X1 key_b_r_reg_12_26 (.CK( clk ) , .D( key_b_r_11_26 ) , .Q( key_b_r_12_26 ) );
  DFF_X1 key_b_r_reg_12_27 (.CK( clk ) , .D( key_b_r_11_27 ) , .Q( key_b_r_12_27 ) );
  DFF_X1 key_b_r_reg_12_28 (.CK( clk ) , .D( key_b_r_11_28 ) , .Q( key_b_r_12_28 ) );
  DFF_X1 key_b_r_reg_12_29 (.CK( clk ) , .D( key_b_r_11_29 ) , .Q( key_b_r_12_29 ) );
  DFF_X1 key_b_r_reg_12_3 (.CK( clk ) , .D( key_b_r_11_3 ) , .Q( key_b_r_12_3 ) );
  DFF_X1 key_b_r_reg_12_30 (.CK( clk ) , .D( key_b_r_11_30 ) , .Q( key_b_r_12_30 ) );
  DFF_X1 key_b_r_reg_12_31 (.CK( clk ) , .D( key_b_r_11_31 ) , .Q( key_b_r_12_31 ) );
  DFF_X1 key_b_r_reg_12_32 (.CK( clk ) , .D( key_b_r_11_32 ) , .Q( key_b_r_12_32 ) );
  DFF_X1 key_b_r_reg_12_33 (.CK( clk ) , .D( key_b_r_11_33 ) , .Q( key_b_r_12_33 ) );
  DFF_X1 key_b_r_reg_12_34 (.CK( clk ) , .D( key_b_r_11_34 ) , .Q( key_b_r_12_34 ) );
  DFF_X1 key_b_r_reg_12_35 (.CK( clk ) , .D( key_b_r_11_35 ) , .Q( key_b_r_12_35 ) );
  DFF_X1 key_b_r_reg_12_36 (.CK( clk ) , .D( key_b_r_11_36 ) , .Q( key_b_r_12_36 ) );
  DFF_X1 key_b_r_reg_12_37 (.CK( clk ) , .D( key_b_r_11_37 ) , .Q( key_b_r_12_37 ) );
  DFF_X1 key_b_r_reg_12_38 (.CK( clk ) , .D( key_b_r_11_38 ) , .Q( key_b_r_12_38 ) );
  DFF_X1 key_b_r_reg_12_39 (.CK( clk ) , .D( key_b_r_11_39 ) , .Q( key_b_r_12_39 ) );
  DFF_X1 key_b_r_reg_12_4 (.CK( clk ) , .D( key_b_r_11_4 ) , .Q( key_b_r_12_4 ) );
  DFF_X1 key_b_r_reg_12_40 (.CK( clk ) , .D( key_b_r_11_40 ) , .Q( key_b_r_12_40 ) );
  DFF_X1 key_b_r_reg_12_41 (.CK( clk ) , .D( key_b_r_11_41 ) , .Q( key_b_r_12_41 ) );
  DFF_X1 key_b_r_reg_12_42 (.CK( clk ) , .D( key_b_r_11_42 ) , .Q( key_b_r_12_42 ) );
  DFF_X1 key_b_r_reg_12_43 (.CK( clk ) , .D( key_b_r_11_43 ) , .Q( key_b_r_12_43 ) );
  DFF_X1 key_b_r_reg_12_44 (.CK( clk ) , .D( key_b_r_11_44 ) , .Q( key_b_r_12_44 ) );
  DFF_X1 key_b_r_reg_12_45 (.CK( clk ) , .D( key_b_r_11_45 ) , .Q( key_b_r_12_45 ) );
  DFF_X1 key_b_r_reg_12_46 (.CK( clk ) , .D( key_b_r_11_46 ) , .Q( key_b_r_12_46 ) );
  DFF_X1 key_b_r_reg_12_47 (.CK( clk ) , .D( key_b_r_11_47 ) , .Q( key_b_r_12_47 ) );
  DFF_X1 key_b_r_reg_12_48 (.CK( clk ) , .D( key_b_r_11_48 ) , .Q( key_b_r_12_48 ) );
  DFF_X1 key_b_r_reg_12_49 (.CK( clk ) , .D( key_b_r_11_49 ) , .Q( key_b_r_12_49 ) );
  DFF_X1 key_b_r_reg_12_5 (.CK( clk ) , .D( key_b_r_11_5 ) , .Q( key_b_r_12_5 ) );
  DFF_X1 key_b_r_reg_12_50 (.CK( clk ) , .D( key_b_r_11_50 ) , .Q( key_b_r_12_50 ) );
  DFF_X1 key_b_r_reg_12_51 (.CK( clk ) , .D( key_b_r_11_51 ) , .Q( key_b_r_12_51 ) );
  DFF_X1 key_b_r_reg_12_52 (.CK( clk ) , .D( key_b_r_11_52 ) , .Q( key_b_r_12_52 ) );
  DFF_X1 key_b_r_reg_12_53 (.CK( clk ) , .D( key_b_r_11_53 ) , .Q( key_b_r_12_53 ) );
  DFF_X1 key_b_r_reg_12_54 (.CK( clk ) , .D( key_b_r_11_54 ) , .Q( key_b_r_12_54 ) );
  DFF_X1 key_b_r_reg_12_55 (.CK( clk ) , .D( key_b_r_11_55 ) , .Q( key_b_r_12_55 ) );
  DFF_X1 key_b_r_reg_12_6 (.CK( clk ) , .D( key_b_r_11_6 ) , .Q( key_b_r_12_6 ) );
  DFF_X1 key_b_r_reg_12_7 (.CK( clk ) , .D( key_b_r_11_7 ) , .Q( key_b_r_12_7 ) );
  DFF_X1 key_b_r_reg_12_8 (.CK( clk ) , .D( key_b_r_11_8 ) , .Q( key_b_r_12_8 ) );
  DFF_X1 key_b_r_reg_12_9 (.CK( clk ) , .D( key_b_r_11_9 ) , .Q( key_b_r_12_9 ) );
  DFF_X1 key_b_r_reg_13_0 (.CK( clk ) , .D( key_b_r_12_0 ) , .Q( key_b_r_13_0 ) );
  DFF_X1 key_b_r_reg_13_1 (.CK( clk ) , .D( key_b_r_12_1 ) , .Q( key_b_r_13_1 ) );
  DFF_X1 key_b_r_reg_13_10 (.CK( clk ) , .D( key_b_r_12_10 ) , .Q( key_b_r_13_10 ) );
  DFF_X1 key_b_r_reg_13_11 (.CK( clk ) , .D( key_b_r_12_11 ) , .Q( key_b_r_13_11 ) );
  DFF_X1 key_b_r_reg_13_12 (.CK( clk ) , .D( key_b_r_12_12 ) , .Q( key_b_r_13_12 ) );
  DFF_X1 key_b_r_reg_13_13 (.CK( clk ) , .D( key_b_r_12_13 ) , .Q( key_b_r_13_13 ) );
  DFF_X1 key_b_r_reg_13_14 (.CK( clk ) , .D( key_b_r_12_14 ) , .Q( key_b_r_13_14 ) );
  DFF_X1 key_b_r_reg_13_15 (.CK( clk ) , .D( key_b_r_12_15 ) , .Q( key_b_r_13_15 ) );
  DFF_X1 key_b_r_reg_13_16 (.CK( clk ) , .D( key_b_r_12_16 ) , .Q( key_b_r_13_16 ) );
  DFF_X1 key_b_r_reg_13_17 (.CK( clk ) , .D( key_b_r_12_17 ) , .Q( key_b_r_13_17 ) );
  DFF_X1 key_b_r_reg_13_18 (.CK( clk ) , .D( key_b_r_12_18 ) , .Q( key_b_r_13_18 ) );
  DFF_X1 key_b_r_reg_13_19 (.CK( clk ) , .D( key_b_r_12_19 ) , .Q( key_b_r_13_19 ) );
  DFF_X1 key_b_r_reg_13_2 (.CK( clk ) , .D( key_b_r_12_2 ) , .Q( key_b_r_13_2 ) );
  DFF_X1 key_b_r_reg_13_20 (.CK( clk ) , .D( key_b_r_12_20 ) , .Q( key_b_r_13_20 ) );
  DFF_X1 key_b_r_reg_13_21 (.CK( clk ) , .D( key_b_r_12_21 ) , .Q( key_b_r_13_21 ) );
  DFF_X1 key_b_r_reg_13_22 (.CK( clk ) , .D( key_b_r_12_22 ) , .Q( key_b_r_13_22 ) );
  DFF_X1 key_b_r_reg_13_23 (.CK( clk ) , .D( key_b_r_12_23 ) , .Q( key_b_r_13_23 ) );
  DFF_X1 key_b_r_reg_13_24 (.CK( clk ) , .D( key_b_r_12_24 ) , .Q( key_b_r_13_24 ) );
  DFF_X1 key_b_r_reg_13_25 (.CK( clk ) , .D( key_b_r_12_25 ) , .Q( key_b_r_13_25 ) );
  DFF_X1 key_b_r_reg_13_26 (.CK( clk ) , .D( key_b_r_12_26 ) , .Q( key_b_r_13_26 ) );
  DFF_X1 key_b_r_reg_13_27 (.CK( clk ) , .D( key_b_r_12_27 ) , .Q( key_b_r_13_27 ) );
  DFF_X1 key_b_r_reg_13_28 (.CK( clk ) , .D( key_b_r_12_28 ) , .Q( key_b_r_13_28 ) );
  DFF_X1 key_b_r_reg_13_29 (.CK( clk ) , .D( key_b_r_12_29 ) , .Q( key_b_r_13_29 ) );
  DFF_X1 key_b_r_reg_13_3 (.CK( clk ) , .D( key_b_r_12_3 ) , .Q( key_b_r_13_3 ) );
  DFF_X1 key_b_r_reg_13_30 (.CK( clk ) , .D( key_b_r_12_30 ) , .Q( key_b_r_13_30 ) );
  DFF_X1 key_b_r_reg_13_31 (.CK( clk ) , .D( key_b_r_12_31 ) , .Q( key_b_r_13_31 ) );
  DFF_X1 key_b_r_reg_13_32 (.CK( clk ) , .D( key_b_r_12_32 ) , .Q( key_b_r_13_32 ) );
  DFF_X1 key_b_r_reg_13_33 (.CK( clk ) , .D( key_b_r_12_33 ) , .Q( key_b_r_13_33 ) );
  DFF_X1 key_b_r_reg_13_34 (.CK( clk ) , .D( key_b_r_12_34 ) , .Q( key_b_r_13_34 ) );
  DFF_X1 key_b_r_reg_13_35 (.CK( clk ) , .D( key_b_r_12_35 ) , .Q( key_b_r_13_35 ) );
  DFF_X1 key_b_r_reg_13_36 (.CK( clk ) , .D( key_b_r_12_36 ) , .Q( key_b_r_13_36 ) );
  DFF_X1 key_b_r_reg_13_37 (.CK( clk ) , .D( key_b_r_12_37 ) , .Q( key_b_r_13_37 ) );
  DFF_X1 key_b_r_reg_13_38 (.CK( clk ) , .D( key_b_r_12_38 ) , .Q( key_b_r_13_38 ) );
  DFF_X1 key_b_r_reg_13_39 (.CK( clk ) , .D( key_b_r_12_39 ) , .Q( key_b_r_13_39 ) );
  DFF_X1 key_b_r_reg_13_4 (.CK( clk ) , .D( key_b_r_12_4 ) , .Q( key_b_r_13_4 ) );
  DFF_X1 key_b_r_reg_13_40 (.CK( clk ) , .D( key_b_r_12_40 ) , .Q( key_b_r_13_40 ) );
  DFF_X1 key_b_r_reg_13_41 (.CK( clk ) , .D( key_b_r_12_41 ) , .Q( key_b_r_13_41 ) );
  DFF_X1 key_b_r_reg_13_42 (.CK( clk ) , .D( key_b_r_12_42 ) , .Q( key_b_r_13_42 ) );
  DFF_X1 key_b_r_reg_13_43 (.CK( clk ) , .D( key_b_r_12_43 ) , .Q( key_b_r_13_43 ) );
  DFF_X1 key_b_r_reg_13_44 (.CK( clk ) , .D( key_b_r_12_44 ) , .Q( key_b_r_13_44 ) );
  DFF_X1 key_b_r_reg_13_45 (.CK( clk ) , .D( key_b_r_12_45 ) , .Q( key_b_r_13_45 ) );
  DFF_X1 key_b_r_reg_13_46 (.CK( clk ) , .D( key_b_r_12_46 ) , .Q( key_b_r_13_46 ) );
  DFF_X1 key_b_r_reg_13_47 (.CK( clk ) , .D( key_b_r_12_47 ) , .Q( key_b_r_13_47 ) );
  DFF_X1 key_b_r_reg_13_48 (.CK( clk ) , .D( key_b_r_12_48 ) , .Q( key_b_r_13_48 ) );
  DFF_X1 key_b_r_reg_13_49 (.CK( clk ) , .D( key_b_r_12_49 ) , .Q( key_b_r_13_49 ) );
  DFF_X1 key_b_r_reg_13_5 (.CK( clk ) , .D( key_b_r_12_5 ) , .Q( key_b_r_13_5 ) );
  DFF_X1 key_b_r_reg_13_50 (.CK( clk ) , .D( key_b_r_12_50 ) , .Q( key_b_r_13_50 ) );
  DFF_X1 key_b_r_reg_13_51 (.CK( clk ) , .D( key_b_r_12_51 ) , .Q( key_b_r_13_51 ) );
  DFF_X1 key_b_r_reg_13_52 (.CK( clk ) , .D( key_b_r_12_52 ) , .Q( key_b_r_13_52 ) );
  DFF_X1 key_b_r_reg_13_53 (.CK( clk ) , .D( key_b_r_12_53 ) , .Q( key_b_r_13_53 ) );
  DFF_X1 key_b_r_reg_13_54 (.CK( clk ) , .D( key_b_r_12_54 ) , .Q( key_b_r_13_54 ) );
  DFF_X1 key_b_r_reg_13_55 (.CK( clk ) , .D( key_b_r_12_55 ) , .Q( key_b_r_13_55 ) );
  DFF_X1 key_b_r_reg_13_6 (.CK( clk ) , .D( key_b_r_12_6 ) , .Q( key_b_r_13_6 ) );
  DFF_X1 key_b_r_reg_13_7 (.CK( clk ) , .D( key_b_r_12_7 ) , .Q( key_b_r_13_7 ) );
  DFF_X1 key_b_r_reg_13_8 (.CK( clk ) , .D( key_b_r_12_8 ) , .Q( key_b_r_13_8 ) );
  DFF_X1 key_b_r_reg_13_9 (.CK( clk ) , .D( key_b_r_12_9 ) , .Q( key_b_r_13_9 ) );
  DFF_X1 key_b_r_reg_14_0 (.CK( clk ) , .D( key_b_r_13_0 ) , .Q( key_b_r_14_0 ) );
  DFF_X1 key_b_r_reg_14_1 (.CK( clk ) , .D( key_b_r_13_1 ) , .Q( key_b_r_14_1 ) );
  DFF_X1 key_b_r_reg_14_10 (.CK( clk ) , .D( key_b_r_13_10 ) , .Q( key_b_r_14_10 ) );
  DFF_X1 key_b_r_reg_14_11 (.CK( clk ) , .D( key_b_r_13_11 ) , .Q( key_b_r_14_11 ) );
  DFF_X1 key_b_r_reg_14_12 (.CK( clk ) , .D( key_b_r_13_12 ) , .Q( key_b_r_14_12 ) );
  DFF_X1 key_b_r_reg_14_13 (.CK( clk ) , .D( key_b_r_13_13 ) , .Q( key_b_r_14_13 ) );
  DFF_X1 key_b_r_reg_14_14 (.CK( clk ) , .D( key_b_r_13_14 ) , .Q( key_b_r_14_14 ) );
  DFF_X1 key_b_r_reg_14_15 (.CK( clk ) , .D( key_b_r_13_15 ) , .Q( key_b_r_14_15 ) );
  DFF_X1 key_b_r_reg_14_16 (.CK( clk ) , .D( key_b_r_13_16 ) , .Q( key_b_r_14_16 ) );
  DFF_X1 key_b_r_reg_14_17 (.CK( clk ) , .D( key_b_r_13_17 ) , .Q( key_b_r_14_17 ) );
  DFF_X1 key_b_r_reg_14_18 (.CK( clk ) , .D( key_b_r_13_18 ) , .Q( key_b_r_14_18 ) );
  DFF_X1 key_b_r_reg_14_19 (.CK( clk ) , .D( key_b_r_13_19 ) , .Q( key_b_r_14_19 ) );
  DFF_X1 key_b_r_reg_14_2 (.CK( clk ) , .D( key_b_r_13_2 ) , .Q( key_b_r_14_2 ) );
  DFF_X1 key_b_r_reg_14_20 (.CK( clk ) , .D( key_b_r_13_20 ) , .Q( key_b_r_14_20 ) );
  DFF_X1 key_b_r_reg_14_21 (.CK( clk ) , .D( key_b_r_13_21 ) , .Q( key_b_r_14_21 ) );
  DFF_X1 key_b_r_reg_14_22 (.CK( clk ) , .D( key_b_r_13_22 ) , .Q( key_b_r_14_22 ) );
  DFF_X1 key_b_r_reg_14_23 (.CK( clk ) , .D( key_b_r_13_23 ) , .Q( key_b_r_14_23 ) );
  DFF_X1 key_b_r_reg_14_24 (.CK( clk ) , .D( key_b_r_13_24 ) , .Q( key_b_r_14_24 ) );
  DFF_X1 key_b_r_reg_14_25 (.CK( clk ) , .D( key_b_r_13_25 ) , .Q( key_b_r_14_25 ) );
  DFF_X1 key_b_r_reg_14_26 (.CK( clk ) , .D( key_b_r_13_26 ) , .Q( key_b_r_14_26 ) );
  DFF_X1 key_b_r_reg_14_27 (.CK( clk ) , .D( key_b_r_13_27 ) , .Q( key_b_r_14_27 ) );
  DFF_X1 key_b_r_reg_14_28 (.CK( clk ) , .D( key_b_r_13_28 ) , .Q( key_b_r_14_28 ) );
  DFF_X1 key_b_r_reg_14_29 (.CK( clk ) , .D( key_b_r_13_29 ) , .Q( key_b_r_14_29 ) );
  DFF_X1 key_b_r_reg_14_3 (.CK( clk ) , .D( key_b_r_13_3 ) , .Q( key_b_r_14_3 ) );
  DFF_X1 key_b_r_reg_14_30 (.CK( clk ) , .D( key_b_r_13_30 ) , .Q( key_b_r_14_30 ) );
  DFF_X1 key_b_r_reg_14_31 (.CK( clk ) , .D( key_b_r_13_31 ) , .Q( key_b_r_14_31 ) );
  DFF_X1 key_b_r_reg_14_32 (.CK( clk ) , .D( key_b_r_13_32 ) , .Q( key_b_r_14_32 ) );
  DFF_X1 key_b_r_reg_14_33 (.CK( clk ) , .D( key_b_r_13_33 ) , .Q( key_b_r_14_33 ) );
  DFF_X1 key_b_r_reg_14_34 (.CK( clk ) , .D( key_b_r_13_34 ) , .Q( key_b_r_14_34 ) );
  DFF_X1 key_b_r_reg_14_35 (.CK( clk ) , .D( key_b_r_13_35 ) , .Q( key_b_r_14_35 ) );
  DFF_X1 key_b_r_reg_14_36 (.CK( clk ) , .D( key_b_r_13_36 ) , .Q( key_b_r_14_36 ) );
  DFF_X1 key_b_r_reg_14_37 (.CK( clk ) , .D( key_b_r_13_37 ) , .Q( key_b_r_14_37 ) );
  DFF_X1 key_b_r_reg_14_38 (.CK( clk ) , .D( key_b_r_13_38 ) , .Q( key_b_r_14_38 ) );
  DFF_X1 key_b_r_reg_14_39 (.CK( clk ) , .D( key_b_r_13_39 ) , .Q( key_b_r_14_39 ) );
  DFF_X1 key_b_r_reg_14_4 (.CK( clk ) , .D( key_b_r_13_4 ) , .Q( key_b_r_14_4 ) );
  DFF_X1 key_b_r_reg_14_40 (.CK( clk ) , .D( key_b_r_13_40 ) , .Q( key_b_r_14_40 ) );
  DFF_X1 key_b_r_reg_14_41 (.CK( clk ) , .D( key_b_r_13_41 ) , .Q( key_b_r_14_41 ) );
  DFF_X1 key_b_r_reg_14_42 (.CK( clk ) , .D( key_b_r_13_42 ) , .Q( key_b_r_14_42 ) );
  DFF_X1 key_b_r_reg_14_43 (.CK( clk ) , .D( key_b_r_13_43 ) , .Q( key_b_r_14_43 ) );
  DFF_X1 key_b_r_reg_14_44 (.CK( clk ) , .D( key_b_r_13_44 ) , .Q( key_b_r_14_44 ) );
  DFF_X1 key_b_r_reg_14_45 (.CK( clk ) , .D( key_b_r_13_45 ) , .Q( key_b_r_14_45 ) );
  DFF_X1 key_b_r_reg_14_46 (.CK( clk ) , .D( key_b_r_13_46 ) , .Q( key_b_r_14_46 ) );
  DFF_X1 key_b_r_reg_14_47 (.CK( clk ) , .D( key_b_r_13_47 ) , .Q( key_b_r_14_47 ) );
  DFF_X1 key_b_r_reg_14_48 (.CK( clk ) , .D( key_b_r_13_48 ) , .Q( key_b_r_14_48 ) );
  DFF_X1 key_b_r_reg_14_49 (.CK( clk ) , .D( key_b_r_13_49 ) , .Q( key_b_r_14_49 ) );
  DFF_X1 key_b_r_reg_14_5 (.CK( clk ) , .D( key_b_r_13_5 ) , .Q( key_b_r_14_5 ) );
  DFF_X1 key_b_r_reg_14_50 (.CK( clk ) , .D( key_b_r_13_50 ) , .Q( key_b_r_14_50 ) );
  DFF_X1 key_b_r_reg_14_51 (.CK( clk ) , .D( key_b_r_13_51 ) , .Q( key_b_r_14_51 ) );
  DFF_X1 key_b_r_reg_14_52 (.CK( clk ) , .D( key_b_r_13_52 ) , .Q( key_b_r_14_52 ) );
  DFF_X1 key_b_r_reg_14_53 (.CK( clk ) , .D( key_b_r_13_53 ) , .Q( key_b_r_14_53 ) );
  DFF_X1 key_b_r_reg_14_54 (.CK( clk ) , .D( key_b_r_13_54 ) , .Q( key_b_r_14_54 ) );
  DFF_X1 key_b_r_reg_14_55 (.CK( clk ) , .D( key_b_r_13_55 ) , .Q( key_b_r_14_55 ) );
  DFF_X1 key_b_r_reg_14_6 (.CK( clk ) , .D( key_b_r_13_6 ) , .Q( key_b_r_14_6 ) );
  DFF_X1 key_b_r_reg_14_7 (.CK( clk ) , .D( key_b_r_13_7 ) , .Q( key_b_r_14_7 ) );
  DFF_X1 key_b_r_reg_14_8 (.CK( clk ) , .D( key_b_r_13_8 ) , .Q( key_b_r_14_8 ) );
  DFF_X1 key_b_r_reg_14_9 (.CK( clk ) , .D( key_b_r_13_9 ) , .Q( key_b_r_14_9 ) );
  DFF_X1 key_b_r_reg_15_0 (.CK( clk ) , .D( key_b_r_14_0 ) , .Q( key_b_r_15_0 ) );
  DFF_X1 key_b_r_reg_15_1 (.CK( clk ) , .D( key_b_r_14_1 ) , .Q( key_b_r_15_1 ) );
  DFF_X1 key_b_r_reg_15_10 (.CK( clk ) , .D( key_b_r_14_10 ) , .Q( key_b_r_15_10 ) );
  DFF_X1 key_b_r_reg_15_11 (.CK( clk ) , .D( key_b_r_14_11 ) , .Q( key_b_r_15_11 ) );
  DFF_X1 key_b_r_reg_15_12 (.CK( clk ) , .D( key_b_r_14_12 ) , .Q( key_b_r_15_12 ) );
  DFF_X1 key_b_r_reg_15_13 (.CK( clk ) , .D( key_b_r_14_13 ) , .Q( key_b_r_15_13 ) );
  DFF_X1 key_b_r_reg_15_14 (.CK( clk ) , .D( key_b_r_14_14 ) , .Q( key_b_r_15_14 ) );
  DFF_X1 key_b_r_reg_15_15 (.CK( clk ) , .D( key_b_r_14_15 ) , .Q( key_b_r_15_15 ) );
  DFF_X1 key_b_r_reg_15_16 (.CK( clk ) , .D( key_b_r_14_16 ) , .Q( key_b_r_15_16 ) );
  DFF_X1 key_b_r_reg_15_17 (.CK( clk ) , .D( key_b_r_14_17 ) , .Q( key_b_r_15_17 ) );
  DFF_X1 key_b_r_reg_15_18 (.CK( clk ) , .D( key_b_r_14_18 ) , .Q( key_b_r_15_18 ) );
  DFF_X1 key_b_r_reg_15_19 (.CK( clk ) , .D( key_b_r_14_19 ) , .Q( key_b_r_15_19 ) );
  DFF_X1 key_b_r_reg_15_2 (.CK( clk ) , .D( key_b_r_14_2 ) , .Q( key_b_r_15_2 ) );
  DFF_X1 key_b_r_reg_15_20 (.CK( clk ) , .D( key_b_r_14_20 ) , .Q( key_b_r_15_20 ) );
  DFF_X1 key_b_r_reg_15_21 (.CK( clk ) , .D( key_b_r_14_21 ) , .Q( key_b_r_15_21 ) );
  DFF_X1 key_b_r_reg_15_22 (.CK( clk ) , .D( key_b_r_14_22 ) , .Q( key_b_r_15_22 ) );
  DFF_X1 key_b_r_reg_15_23 (.CK( clk ) , .D( key_b_r_14_23 ) , .Q( key_b_r_15_23 ) );
  DFF_X1 key_b_r_reg_15_24 (.CK( clk ) , .D( key_b_r_14_24 ) , .Q( key_b_r_15_24 ) );
  DFF_X1 key_b_r_reg_15_25 (.CK( clk ) , .D( key_b_r_14_25 ) , .Q( key_b_r_15_25 ) );
  DFF_X1 key_b_r_reg_15_26 (.CK( clk ) , .D( key_b_r_14_26 ) , .Q( key_b_r_15_26 ) );
  DFF_X1 key_b_r_reg_15_27 (.CK( clk ) , .D( key_b_r_14_27 ) , .Q( key_b_r_15_27 ) );
  DFF_X1 key_b_r_reg_15_28 (.CK( clk ) , .D( key_b_r_14_28 ) , .Q( key_b_r_15_28 ) );
  DFF_X1 key_b_r_reg_15_29 (.CK( clk ) , .D( key_b_r_14_29 ) , .Q( key_b_r_15_29 ) );
  DFF_X1 key_b_r_reg_15_3 (.CK( clk ) , .D( key_b_r_14_3 ) , .Q( key_b_r_15_3 ) );
  DFF_X1 key_b_r_reg_15_30 (.CK( clk ) , .D( key_b_r_14_30 ) , .Q( key_b_r_15_30 ) );
  DFF_X1 key_b_r_reg_15_31 (.CK( clk ) , .D( key_b_r_14_31 ) , .Q( key_b_r_15_31 ) );
  DFF_X1 key_b_r_reg_15_32 (.CK( clk ) , .D( key_b_r_14_32 ) , .Q( key_b_r_15_32 ) );
  DFF_X1 key_b_r_reg_15_33 (.CK( clk ) , .D( key_b_r_14_33 ) , .Q( key_b_r_15_33 ) );
  DFF_X1 key_b_r_reg_15_34 (.CK( clk ) , .D( key_b_r_14_34 ) , .Q( key_b_r_15_34 ) );
  DFF_X1 key_b_r_reg_15_35 (.CK( clk ) , .D( key_b_r_14_35 ) , .Q( key_b_r_15_35 ) );
  DFF_X1 key_b_r_reg_15_36 (.CK( clk ) , .D( key_b_r_14_36 ) , .Q( key_b_r_15_36 ) );
  DFF_X1 key_b_r_reg_15_37 (.CK( clk ) , .D( key_b_r_14_37 ) , .Q( key_b_r_15_37 ) );
  DFF_X1 key_b_r_reg_15_38 (.CK( clk ) , .D( key_b_r_14_38 ) , .Q( key_b_r_15_38 ) );
  DFF_X1 key_b_r_reg_15_39 (.CK( clk ) , .D( key_b_r_14_39 ) , .Q( key_b_r_15_39 ) );
  DFF_X1 key_b_r_reg_15_4 (.CK( clk ) , .D( key_b_r_14_4 ) , .Q( key_b_r_15_4 ) );
  DFF_X1 key_b_r_reg_15_40 (.CK( clk ) , .D( key_b_r_14_40 ) , .Q( key_b_r_15_40 ) );
  DFF_X1 key_b_r_reg_15_41 (.CK( clk ) , .D( key_b_r_14_41 ) , .Q( key_b_r_15_41 ) );
  DFF_X1 key_b_r_reg_15_42 (.CK( clk ) , .D( key_b_r_14_42 ) , .Q( key_b_r_15_42 ) );
  DFF_X1 key_b_r_reg_15_43 (.CK( clk ) , .D( key_b_r_14_43 ) , .Q( key_b_r_15_43 ) );
  DFF_X1 key_b_r_reg_15_44 (.CK( clk ) , .D( key_b_r_14_44 ) , .Q( key_b_r_15_44 ) );
  DFF_X1 key_b_r_reg_15_45 (.CK( clk ) , .D( key_b_r_14_45 ) , .Q( key_b_r_15_45 ) );
  DFF_X1 key_b_r_reg_15_46 (.CK( clk ) , .D( key_b_r_14_46 ) , .Q( key_b_r_15_46 ) );
  DFF_X1 key_b_r_reg_15_47 (.CK( clk ) , .D( key_b_r_14_47 ) , .Q( key_b_r_15_47 ) );
  DFF_X1 key_b_r_reg_15_48 (.CK( clk ) , .D( key_b_r_14_48 ) , .Q( key_b_r_15_48 ) );
  DFF_X1 key_b_r_reg_15_49 (.CK( clk ) , .D( key_b_r_14_49 ) , .Q( key_b_r_15_49 ) );
  DFF_X1 key_b_r_reg_15_5 (.CK( clk ) , .D( key_b_r_14_5 ) , .Q( key_b_r_15_5 ) );
  DFF_X1 key_b_r_reg_15_50 (.CK( clk ) , .D( key_b_r_14_50 ) , .Q( key_b_r_15_50 ) );
  DFF_X1 key_b_r_reg_15_51 (.CK( clk ) , .D( key_b_r_14_51 ) , .Q( key_b_r_15_51 ) );
  DFF_X1 key_b_r_reg_15_52 (.CK( clk ) , .D( key_b_r_14_52 ) , .Q( key_b_r_15_52 ) );
  DFF_X1 key_b_r_reg_15_53 (.CK( clk ) , .D( key_b_r_14_53 ) , .Q( key_b_r_15_53 ) );
  DFF_X1 key_b_r_reg_15_54 (.CK( clk ) , .D( key_b_r_14_54 ) , .Q( key_b_r_15_54 ) );
  DFF_X1 key_b_r_reg_15_55 (.CK( clk ) , .D( key_b_r_14_55 ) , .Q( key_b_r_15_55 ) );
  DFF_X1 key_b_r_reg_15_6 (.CK( clk ) , .D( key_b_r_14_6 ) , .Q( key_b_r_15_6 ) );
  DFF_X1 key_b_r_reg_15_7 (.CK( clk ) , .D( key_b_r_14_7 ) , .Q( key_b_r_15_7 ) );
  DFF_X1 key_b_r_reg_15_8 (.CK( clk ) , .D( key_b_r_14_8 ) , .Q( key_b_r_15_8 ) );
  DFF_X1 key_b_r_reg_15_9 (.CK( clk ) , .D( key_b_r_14_9 ) , .Q( key_b_r_15_9 ) );
  DFF_X1 key_b_r_reg_16_0 (.CK( clk ) , .D( key_b_r_15_0 ) , .Q( key_b_r_16_0 ) );
  DFF_X1 key_b_r_reg_16_1 (.CK( clk ) , .D( key_b_r_15_1 ) , .Q( key_b_r_16_1 ) );
  DFF_X1 key_b_r_reg_16_10 (.CK( clk ) , .D( key_b_r_15_10 ) , .Q( key_b_r_16_10 ) );
  DFF_X1 key_b_r_reg_16_11 (.CK( clk ) , .D( key_b_r_15_11 ) , .Q( key_b_r_16_11 ) );
  DFF_X1 key_b_r_reg_16_12 (.CK( clk ) , .D( key_b_r_15_12 ) , .Q( key_b_r_16_12 ) );
  DFF_X1 key_b_r_reg_16_13 (.CK( clk ) , .D( key_b_r_15_13 ) , .Q( key_b_r_16_13 ) );
  DFF_X1 key_b_r_reg_16_14 (.CK( clk ) , .D( key_b_r_15_14 ) , .Q( key_b_r_16_14 ) );
  DFF_X1 key_b_r_reg_16_15 (.CK( clk ) , .D( key_b_r_15_15 ) , .Q( key_b_r_16_15 ) );
  DFF_X1 key_b_r_reg_16_16 (.CK( clk ) , .D( key_b_r_15_16 ) , .Q( key_b_r_16_16 ) );
  DFF_X1 key_b_r_reg_16_17 (.CK( clk ) , .D( key_b_r_15_17 ) , .Q( key_b_r_16_17 ) );
  DFF_X1 key_b_r_reg_16_18 (.CK( clk ) , .D( key_b_r_15_18 ) , .Q( key_b_r_16_18 ) );
  DFF_X1 key_b_r_reg_16_19 (.CK( clk ) , .D( key_b_r_15_19 ) , .Q( key_b_r_16_19 ) );
  DFF_X1 key_b_r_reg_16_2 (.CK( clk ) , .D( key_b_r_15_2 ) , .Q( key_b_r_16_2 ) );
  DFF_X1 key_b_r_reg_16_20 (.CK( clk ) , .D( key_b_r_15_20 ) , .Q( key_b_r_16_20 ) );
  DFF_X1 key_b_r_reg_16_21 (.CK( clk ) , .D( key_b_r_15_21 ) , .Q( key_b_r_16_21 ) );
  DFF_X1 key_b_r_reg_16_22 (.CK( clk ) , .D( key_b_r_15_22 ) , .Q( key_b_r_16_22 ) );
  DFF_X1 key_b_r_reg_16_23 (.CK( clk ) , .D( key_b_r_15_23 ) , .Q( key_b_r_16_23 ) );
  DFF_X1 key_b_r_reg_16_24 (.CK( clk ) , .D( key_b_r_15_24 ) , .Q( key_b_r_16_24 ) );
  DFF_X1 key_b_r_reg_16_25 (.CK( clk ) , .D( key_b_r_15_25 ) , .Q( key_b_r_16_25 ) );
  DFF_X1 key_b_r_reg_16_26 (.CK( clk ) , .D( key_b_r_15_26 ) , .Q( key_b_r_16_26 ) );
  DFF_X1 key_b_r_reg_16_27 (.CK( clk ) , .D( key_b_r_15_27 ) , .Q( key_b_r_16_27 ) );
  DFF_X1 key_b_r_reg_16_28 (.CK( clk ) , .D( key_b_r_15_28 ) , .Q( key_b_r_16_28 ) );
  DFF_X1 key_b_r_reg_16_29 (.CK( clk ) , .D( key_b_r_15_29 ) , .Q( key_b_r_16_29 ) );
  DFF_X1 key_b_r_reg_16_3 (.CK( clk ) , .D( key_b_r_15_3 ) , .Q( key_b_r_16_3 ) );
  DFF_X1 key_b_r_reg_16_30 (.CK( clk ) , .D( key_b_r_15_30 ) , .Q( key_b_r_16_30 ) );
  DFF_X1 key_b_r_reg_16_31 (.CK( clk ) , .D( key_b_r_15_31 ) , .Q( key_b_r_16_31 ) );
  DFF_X1 key_b_r_reg_16_32 (.CK( clk ) , .D( key_b_r_15_32 ) , .Q( key_b_r_16_32 ) );
  DFF_X1 key_b_r_reg_16_33 (.CK( clk ) , .D( key_b_r_15_33 ) , .Q( key_b_r_16_33 ) );
  DFF_X1 key_b_r_reg_16_34 (.CK( clk ) , .D( key_b_r_15_34 ) , .Q( key_b_r_16_34 ) );
  DFF_X1 key_b_r_reg_16_35 (.CK( clk ) , .D( key_b_r_15_35 ) , .Q( key_b_r_16_35 ) );
  DFF_X1 key_b_r_reg_16_36 (.CK( clk ) , .D( key_b_r_15_36 ) , .Q( key_b_r_16_36 ) );
  DFF_X1 key_b_r_reg_16_37 (.CK( clk ) , .D( key_b_r_15_37 ) , .Q( key_b_r_16_37 ) );
  DFF_X1 key_b_r_reg_16_38 (.CK( clk ) , .D( key_b_r_15_38 ) , .Q( key_b_r_16_38 ) );
  DFF_X1 key_b_r_reg_16_39 (.CK( clk ) , .D( key_b_r_15_39 ) , .Q( key_b_r_16_39 ) );
  DFF_X1 key_b_r_reg_16_4 (.CK( clk ) , .D( key_b_r_15_4 ) , .Q( key_b_r_16_4 ) );
  DFF_X1 key_b_r_reg_16_40 (.CK( clk ) , .D( key_b_r_15_40 ) , .Q( key_b_r_16_40 ) );
  DFF_X1 key_b_r_reg_16_41 (.CK( clk ) , .D( key_b_r_15_41 ) , .Q( key_b_r_16_41 ) );
  DFF_X1 key_b_r_reg_16_42 (.CK( clk ) , .D( key_b_r_15_42 ) , .Q( key_b_r_16_42 ) );
  DFF_X1 key_b_r_reg_16_43 (.CK( clk ) , .D( key_b_r_15_43 ) , .Q( key_b_r_16_43 ) );
  DFF_X1 key_b_r_reg_16_44 (.CK( clk ) , .D( key_b_r_15_44 ) , .Q( key_b_r_16_44 ) );
  DFF_X1 key_b_r_reg_16_45 (.CK( clk ) , .D( key_b_r_15_45 ) , .Q( key_b_r_16_45 ) );
  DFF_X1 key_b_r_reg_16_46 (.CK( clk ) , .D( key_b_r_15_46 ) , .Q( key_b_r_16_46 ) );
  DFF_X1 key_b_r_reg_16_47 (.CK( clk ) , .D( key_b_r_15_47 ) , .Q( key_b_r_16_47 ) );
  DFF_X1 key_b_r_reg_16_48 (.CK( clk ) , .D( key_b_r_15_48 ) , .Q( key_b_r_16_48 ) );
  DFF_X1 key_b_r_reg_16_49 (.CK( clk ) , .D( key_b_r_15_49 ) , .Q( key_b_r_16_49 ) );
  DFF_X1 key_b_r_reg_16_5 (.CK( clk ) , .D( key_b_r_15_5 ) , .Q( key_b_r_16_5 ) );
  DFF_X1 key_b_r_reg_16_50 (.CK( clk ) , .D( key_b_r_15_50 ) , .Q( key_b_r_16_50 ) );
  DFF_X1 key_b_r_reg_16_51 (.CK( clk ) , .D( key_b_r_15_51 ) , .Q( key_b_r_16_51 ) );
  DFF_X1 key_b_r_reg_16_52 (.CK( clk ) , .D( key_b_r_15_52 ) , .Q( key_b_r_16_52 ) );
  DFF_X1 key_b_r_reg_16_53 (.CK( clk ) , .D( key_b_r_15_53 ) , .Q( key_b_r_16_53 ) );
  DFF_X1 key_b_r_reg_16_54 (.CK( clk ) , .D( key_b_r_15_54 ) , .Q( key_b_r_16_54 ) );
  DFF_X1 key_b_r_reg_16_55 (.CK( clk ) , .D( key_b_r_15_55 ) , .Q( key_b_r_16_55 ) );
  DFF_X1 key_b_r_reg_16_6 (.CK( clk ) , .D( key_b_r_15_6 ) , .Q( key_b_r_16_6 ) );
  DFF_X1 key_b_r_reg_16_7 (.CK( clk ) , .D( key_b_r_15_7 ) , .Q( key_b_r_16_7 ) );
  DFF_X1 key_b_r_reg_16_8 (.CK( clk ) , .D( key_b_r_15_8 ) , .Q( key_b_r_16_8 ) );
  DFF_X1 key_b_r_reg_16_9 (.CK( clk ) , .D( key_b_r_15_9 ) , .Q( key_b_r_16_9 ) );
  DFF_X1 key_b_r_reg_1_0 (.CK( clk ) , .D( key_b_r_0_0 ) , .Q( key_b_r_1_0 ) );
  DFF_X1 key_b_r_reg_1_1 (.CK( clk ) , .D( key_b_r_0_1 ) , .Q( key_b_r_1_1 ) );
  DFF_X1 key_b_r_reg_1_10 (.CK( clk ) , .D( key_b_r_0_10 ) , .Q( key_b_r_1_10 ) );
  DFF_X1 key_b_r_reg_1_11 (.CK( clk ) , .D( key_b_r_0_11 ) , .Q( key_b_r_1_11 ) );
  DFF_X1 key_b_r_reg_1_12 (.CK( clk ) , .D( key_b_r_0_12 ) , .Q( key_b_r_1_12 ) );
  DFF_X1 key_b_r_reg_1_13 (.CK( clk ) , .D( key_b_r_0_13 ) , .Q( key_b_r_1_13 ) );
  DFF_X1 key_b_r_reg_1_14 (.CK( clk ) , .D( key_b_r_0_14 ) , .Q( key_b_r_1_14 ) );
  DFF_X1 key_b_r_reg_1_15 (.CK( clk ) , .D( key_b_r_0_15 ) , .Q( key_b_r_1_15 ) );
  DFF_X1 key_b_r_reg_1_16 (.CK( clk ) , .D( key_b_r_0_16 ) , .Q( key_b_r_1_16 ) );
  DFF_X1 key_b_r_reg_1_17 (.CK( clk ) , .D( key_b_r_0_17 ) , .Q( key_b_r_1_17 ) );
  DFF_X1 key_b_r_reg_1_18 (.CK( clk ) , .D( key_b_r_0_18 ) , .Q( key_b_r_1_18 ) );
  DFF_X1 key_b_r_reg_1_19 (.CK( clk ) , .D( key_b_r_0_19 ) , .Q( key_b_r_1_19 ) );
  DFF_X1 key_b_r_reg_1_2 (.CK( clk ) , .D( key_b_r_0_2 ) , .Q( key_b_r_1_2 ) );
  DFF_X1 key_b_r_reg_1_20 (.CK( clk ) , .D( key_b_r_0_20 ) , .Q( key_b_r_1_20 ) );
  DFF_X1 key_b_r_reg_1_21 (.CK( clk ) , .D( key_b_r_0_21 ) , .Q( key_b_r_1_21 ) );
  DFF_X1 key_b_r_reg_1_22 (.CK( clk ) , .D( key_b_r_0_22 ) , .Q( key_b_r_1_22 ) );
  DFF_X1 key_b_r_reg_1_23 (.CK( clk ) , .D( key_b_r_0_23 ) , .Q( key_b_r_1_23 ) );
  DFF_X1 key_b_r_reg_1_24 (.CK( clk ) , .D( key_b_r_0_24 ) , .Q( key_b_r_1_24 ) );
  DFF_X1 key_b_r_reg_1_25 (.CK( clk ) , .D( key_b_r_0_25 ) , .Q( key_b_r_1_25 ) );
  DFF_X1 key_b_r_reg_1_26 (.CK( clk ) , .D( key_b_r_0_26 ) , .Q( key_b_r_1_26 ) );
  DFF_X1 key_b_r_reg_1_27 (.CK( clk ) , .D( key_b_r_0_27 ) , .Q( key_b_r_1_27 ) );
  DFF_X1 key_b_r_reg_1_28 (.CK( clk ) , .D( key_b_r_0_28 ) , .Q( key_b_r_1_28 ) );
  DFF_X1 key_b_r_reg_1_29 (.CK( clk ) , .D( key_b_r_0_29 ) , .Q( key_b_r_1_29 ) );
  DFF_X1 key_b_r_reg_1_3 (.CK( clk ) , .D( key_b_r_0_3 ) , .Q( key_b_r_1_3 ) );
  DFF_X1 key_b_r_reg_1_30 (.CK( clk ) , .D( key_b_r_0_30 ) , .Q( key_b_r_1_30 ) );
  DFF_X1 key_b_r_reg_1_31 (.CK( clk ) , .D( key_b_r_0_31 ) , .Q( key_b_r_1_31 ) );
  DFF_X1 key_b_r_reg_1_32 (.CK( clk ) , .D( key_b_r_0_32 ) , .Q( key_b_r_1_32 ) );
  DFF_X1 key_b_r_reg_1_33 (.CK( clk ) , .D( key_b_r_0_33 ) , .Q( key_b_r_1_33 ) );
  DFF_X1 key_b_r_reg_1_34 (.CK( clk ) , .D( key_b_r_0_34 ) , .Q( key_b_r_1_34 ) );
  DFF_X1 key_b_r_reg_1_35 (.CK( clk ) , .D( key_b_r_0_35 ) , .Q( key_b_r_1_35 ) );
  DFF_X1 key_b_r_reg_1_36 (.CK( clk ) , .D( key_b_r_0_36 ) , .Q( key_b_r_1_36 ) );
  DFF_X1 key_b_r_reg_1_37 (.CK( clk ) , .D( key_b_r_0_37 ) , .Q( key_b_r_1_37 ) );
  DFF_X1 key_b_r_reg_1_38 (.CK( clk ) , .D( key_b_r_0_38 ) , .Q( key_b_r_1_38 ) );
  DFF_X1 key_b_r_reg_1_39 (.CK( clk ) , .D( key_b_r_0_39 ) , .Q( key_b_r_1_39 ) );
  DFF_X1 key_b_r_reg_1_4 (.CK( clk ) , .D( key_b_r_0_4 ) , .Q( key_b_r_1_4 ) );
  DFF_X1 key_b_r_reg_1_40 (.CK( clk ) , .D( key_b_r_0_40 ) , .Q( key_b_r_1_40 ) );
  DFF_X1 key_b_r_reg_1_41 (.CK( clk ) , .D( key_b_r_0_41 ) , .Q( key_b_r_1_41 ) );
  DFF_X1 key_b_r_reg_1_42 (.CK( clk ) , .D( key_b_r_0_42 ) , .Q( key_b_r_1_42 ) );
  DFF_X1 key_b_r_reg_1_43 (.CK( clk ) , .D( key_b_r_0_43 ) , .Q( key_b_r_1_43 ) );
  DFF_X1 key_b_r_reg_1_44 (.CK( clk ) , .D( key_b_r_0_44 ) , .Q( key_b_r_1_44 ) );
  DFF_X1 key_b_r_reg_1_45 (.CK( clk ) , .D( key_b_r_0_45 ) , .Q( key_b_r_1_45 ) );
  DFF_X1 key_b_r_reg_1_46 (.CK( clk ) , .D( key_b_r_0_46 ) , .Q( key_b_r_1_46 ) );
  DFF_X1 key_b_r_reg_1_47 (.CK( clk ) , .D( key_b_r_0_47 ) , .Q( key_b_r_1_47 ) );
  DFF_X1 key_b_r_reg_1_48 (.CK( clk ) , .D( key_b_r_0_48 ) , .Q( key_b_r_1_48 ) );
  DFF_X1 key_b_r_reg_1_49 (.CK( clk ) , .D( key_b_r_0_49 ) , .Q( key_b_r_1_49 ) );
  DFF_X1 key_b_r_reg_1_5 (.CK( clk ) , .D( key_b_r_0_5 ) , .Q( key_b_r_1_5 ) );
  DFF_X1 key_b_r_reg_1_50 (.CK( clk ) , .D( key_b_r_0_50 ) , .Q( key_b_r_1_50 ) );
  DFF_X1 key_b_r_reg_1_51 (.CK( clk ) , .D( key_b_r_0_51 ) , .Q( key_b_r_1_51 ) );
  DFF_X1 key_b_r_reg_1_52 (.CK( clk ) , .D( key_b_r_0_52 ) , .Q( key_b_r_1_52 ) );
  DFF_X1 key_b_r_reg_1_53 (.CK( clk ) , .D( key_b_r_0_53 ) , .Q( key_b_r_1_53 ) );
  DFF_X1 key_b_r_reg_1_54 (.CK( clk ) , .D( key_b_r_0_54 ) , .Q( key_b_r_1_54 ) );
  DFF_X1 key_b_r_reg_1_55 (.CK( clk ) , .D( key_b_r_0_55 ) , .Q( key_b_r_1_55 ) );
  DFF_X1 key_b_r_reg_1_6 (.CK( clk ) , .D( key_b_r_0_6 ) , .Q( key_b_r_1_6 ) );
  DFF_X1 key_b_r_reg_1_7 (.CK( clk ) , .D( key_b_r_0_7 ) , .Q( key_b_r_1_7 ) );
  DFF_X1 key_b_r_reg_1_8 (.CK( clk ) , .D( key_b_r_0_8 ) , .Q( key_b_r_1_8 ) );
  DFF_X1 key_b_r_reg_1_9 (.CK( clk ) , .D( key_b_r_0_9 ) , .Q( key_b_r_1_9 ) );
  DFF_X1 key_b_r_reg_2_0 (.CK( clk ) , .D( key_b_r_1_0 ) , .Q( key_b_r_2_0 ) );
  DFF_X1 key_b_r_reg_2_1 (.CK( clk ) , .D( key_b_r_1_1 ) , .Q( key_b_r_2_1 ) );
  DFF_X1 key_b_r_reg_2_10 (.CK( clk ) , .D( key_b_r_1_10 ) , .Q( key_b_r_2_10 ) );
  DFF_X1 key_b_r_reg_2_11 (.CK( clk ) , .D( key_b_r_1_11 ) , .Q( key_b_r_2_11 ) );
  DFF_X1 key_b_r_reg_2_12 (.CK( clk ) , .D( key_b_r_1_12 ) , .Q( key_b_r_2_12 ) );
  DFF_X1 key_b_r_reg_2_13 (.CK( clk ) , .D( key_b_r_1_13 ) , .Q( key_b_r_2_13 ) );
  DFF_X1 key_b_r_reg_2_14 (.CK( clk ) , .D( key_b_r_1_14 ) , .Q( key_b_r_2_14 ) );
  DFF_X1 key_b_r_reg_2_15 (.CK( clk ) , .D( key_b_r_1_15 ) , .Q( key_b_r_2_15 ) );
  DFF_X1 key_b_r_reg_2_16 (.CK( clk ) , .D( key_b_r_1_16 ) , .Q( key_b_r_2_16 ) );
  DFF_X1 key_b_r_reg_2_17 (.CK( clk ) , .D( key_b_r_1_17 ) , .Q( key_b_r_2_17 ) );
  DFF_X1 key_b_r_reg_2_18 (.CK( clk ) , .D( key_b_r_1_18 ) , .Q( key_b_r_2_18 ) );
  DFF_X1 key_b_r_reg_2_19 (.CK( clk ) , .D( key_b_r_1_19 ) , .Q( key_b_r_2_19 ) );
  DFF_X1 key_b_r_reg_2_2 (.CK( clk ) , .D( key_b_r_1_2 ) , .Q( key_b_r_2_2 ) );
  DFF_X1 key_b_r_reg_2_20 (.CK( clk ) , .D( key_b_r_1_20 ) , .Q( key_b_r_2_20 ) );
  DFF_X1 key_b_r_reg_2_21 (.CK( clk ) , .D( key_b_r_1_21 ) , .Q( key_b_r_2_21 ) );
  DFF_X1 key_b_r_reg_2_22 (.CK( clk ) , .D( key_b_r_1_22 ) , .Q( key_b_r_2_22 ) );
  DFF_X1 key_b_r_reg_2_23 (.CK( clk ) , .D( key_b_r_1_23 ) , .Q( key_b_r_2_23 ) );
  DFF_X1 key_b_r_reg_2_24 (.CK( clk ) , .D( key_b_r_1_24 ) , .Q( key_b_r_2_24 ) );
  DFF_X1 key_b_r_reg_2_25 (.CK( clk ) , .D( key_b_r_1_25 ) , .Q( key_b_r_2_25 ) );
  DFF_X1 key_b_r_reg_2_26 (.CK( clk ) , .D( key_b_r_1_26 ) , .Q( key_b_r_2_26 ) );
  DFF_X1 key_b_r_reg_2_27 (.CK( clk ) , .D( key_b_r_1_27 ) , .Q( key_b_r_2_27 ) );
  DFF_X1 key_b_r_reg_2_28 (.CK( clk ) , .D( key_b_r_1_28 ) , .Q( key_b_r_2_28 ) );
  DFF_X1 key_b_r_reg_2_29 (.CK( clk ) , .D( key_b_r_1_29 ) , .Q( key_b_r_2_29 ) );
  DFF_X1 key_b_r_reg_2_3 (.CK( clk ) , .D( key_b_r_1_3 ) , .Q( key_b_r_2_3 ) );
  DFF_X1 key_b_r_reg_2_30 (.CK( clk ) , .D( key_b_r_1_30 ) , .Q( key_b_r_2_30 ) );
  DFF_X1 key_b_r_reg_2_31 (.CK( clk ) , .D( key_b_r_1_31 ) , .Q( key_b_r_2_31 ) );
  DFF_X1 key_b_r_reg_2_32 (.CK( clk ) , .D( key_b_r_1_32 ) , .Q( key_b_r_2_32 ) );
  DFF_X1 key_b_r_reg_2_33 (.CK( clk ) , .D( key_b_r_1_33 ) , .Q( key_b_r_2_33 ) );
  DFF_X1 key_b_r_reg_2_34 (.CK( clk ) , .D( key_b_r_1_34 ) , .Q( key_b_r_2_34 ) );
  DFF_X1 key_b_r_reg_2_35 (.CK( clk ) , .D( key_b_r_1_35 ) , .Q( key_b_r_2_35 ) );
  DFF_X1 key_b_r_reg_2_36 (.CK( clk ) , .D( key_b_r_1_36 ) , .Q( key_b_r_2_36 ) );
  DFF_X1 key_b_r_reg_2_37 (.CK( clk ) , .D( key_b_r_1_37 ) , .Q( key_b_r_2_37 ) );
  DFF_X1 key_b_r_reg_2_38 (.CK( clk ) , .D( key_b_r_1_38 ) , .Q( key_b_r_2_38 ) );
  DFF_X1 key_b_r_reg_2_39 (.CK( clk ) , .D( key_b_r_1_39 ) , .Q( key_b_r_2_39 ) );
  DFF_X1 key_b_r_reg_2_4 (.CK( clk ) , .D( key_b_r_1_4 ) , .Q( key_b_r_2_4 ) );
  DFF_X1 key_b_r_reg_2_40 (.CK( clk ) , .D( key_b_r_1_40 ) , .Q( key_b_r_2_40 ) );
  DFF_X1 key_b_r_reg_2_41 (.CK( clk ) , .D( key_b_r_1_41 ) , .Q( key_b_r_2_41 ) );
  DFF_X1 key_b_r_reg_2_42 (.CK( clk ) , .D( key_b_r_1_42 ) , .Q( key_b_r_2_42 ) );
  DFF_X1 key_b_r_reg_2_43 (.CK( clk ) , .D( key_b_r_1_43 ) , .Q( key_b_r_2_43 ) );
  DFF_X1 key_b_r_reg_2_44 (.CK( clk ) , .D( key_b_r_1_44 ) , .Q( key_b_r_2_44 ) );
  DFF_X1 key_b_r_reg_2_45 (.CK( clk ) , .D( key_b_r_1_45 ) , .Q( key_b_r_2_45 ) );
  DFF_X1 key_b_r_reg_2_46 (.CK( clk ) , .D( key_b_r_1_46 ) , .Q( key_b_r_2_46 ) );
  DFF_X1 key_b_r_reg_2_47 (.CK( clk ) , .D( key_b_r_1_47 ) , .Q( key_b_r_2_47 ) );
  DFF_X1 key_b_r_reg_2_48 (.CK( clk ) , .D( key_b_r_1_48 ) , .Q( key_b_r_2_48 ) );
  DFF_X1 key_b_r_reg_2_49 (.CK( clk ) , .D( key_b_r_1_49 ) , .Q( key_b_r_2_49 ) );
  DFF_X1 key_b_r_reg_2_5 (.CK( clk ) , .D( key_b_r_1_5 ) , .Q( key_b_r_2_5 ) );
  DFF_X1 key_b_r_reg_2_50 (.CK( clk ) , .D( key_b_r_1_50 ) , .Q( key_b_r_2_50 ) );
  DFF_X1 key_b_r_reg_2_51 (.CK( clk ) , .D( key_b_r_1_51 ) , .Q( key_b_r_2_51 ) );
  DFF_X1 key_b_r_reg_2_52 (.CK( clk ) , .D( key_b_r_1_52 ) , .Q( key_b_r_2_52 ) );
  DFF_X1 key_b_r_reg_2_53 (.CK( clk ) , .D( key_b_r_1_53 ) , .Q( key_b_r_2_53 ) );
  DFF_X1 key_b_r_reg_2_54 (.CK( clk ) , .D( key_b_r_1_54 ) , .Q( key_b_r_2_54 ) );
  DFF_X1 key_b_r_reg_2_55 (.CK( clk ) , .D( key_b_r_1_55 ) , .Q( key_b_r_2_55 ) );
  DFF_X1 key_b_r_reg_2_6 (.CK( clk ) , .D( key_b_r_1_6 ) , .Q( key_b_r_2_6 ) );
  DFF_X1 key_b_r_reg_2_7 (.CK( clk ) , .D( key_b_r_1_7 ) , .Q( key_b_r_2_7 ) );
  DFF_X1 key_b_r_reg_2_8 (.CK( clk ) , .D( key_b_r_1_8 ) , .Q( key_b_r_2_8 ) );
  DFF_X1 key_b_r_reg_2_9 (.CK( clk ) , .D( key_b_r_1_9 ) , .Q( key_b_r_2_9 ) );
  DFF_X1 key_b_r_reg_3_0 (.CK( clk ) , .D( key_b_r_2_0 ) , .Q( key_b_r_3_0 ) );
  DFF_X1 key_b_r_reg_3_1 (.CK( clk ) , .D( key_b_r_2_1 ) , .Q( key_b_r_3_1 ) );
  DFF_X1 key_b_r_reg_3_10 (.CK( clk ) , .D( key_b_r_2_10 ) , .Q( key_b_r_3_10 ) );
  DFF_X1 key_b_r_reg_3_11 (.CK( clk ) , .D( key_b_r_2_11 ) , .Q( key_b_r_3_11 ) );
  DFF_X1 key_b_r_reg_3_12 (.CK( clk ) , .D( key_b_r_2_12 ) , .Q( key_b_r_3_12 ) );
  DFF_X1 key_b_r_reg_3_13 (.CK( clk ) , .D( key_b_r_2_13 ) , .Q( key_b_r_3_13 ) );
  DFF_X1 key_b_r_reg_3_14 (.CK( clk ) , .D( key_b_r_2_14 ) , .Q( key_b_r_3_14 ) );
  DFF_X1 key_b_r_reg_3_15 (.CK( clk ) , .D( key_b_r_2_15 ) , .Q( key_b_r_3_15 ) );
  DFF_X1 key_b_r_reg_3_16 (.CK( clk ) , .D( key_b_r_2_16 ) , .Q( key_b_r_3_16 ) );
  DFF_X1 key_b_r_reg_3_17 (.CK( clk ) , .D( key_b_r_2_17 ) , .Q( key_b_r_3_17 ) );
  DFF_X1 key_b_r_reg_3_18 (.CK( clk ) , .D( key_b_r_2_18 ) , .Q( key_b_r_3_18 ) );
  DFF_X1 key_b_r_reg_3_19 (.CK( clk ) , .D( key_b_r_2_19 ) , .Q( key_b_r_3_19 ) );
  DFF_X1 key_b_r_reg_3_2 (.CK( clk ) , .D( key_b_r_2_2 ) , .Q( key_b_r_3_2 ) );
  DFF_X1 key_b_r_reg_3_20 (.CK( clk ) , .D( key_b_r_2_20 ) , .Q( key_b_r_3_20 ) );
  DFF_X1 key_b_r_reg_3_21 (.CK( clk ) , .D( key_b_r_2_21 ) , .Q( key_b_r_3_21 ) );
  DFF_X1 key_b_r_reg_3_22 (.CK( clk ) , .D( key_b_r_2_22 ) , .Q( key_b_r_3_22 ) );
  DFF_X1 key_b_r_reg_3_23 (.CK( clk ) , .D( key_b_r_2_23 ) , .Q( key_b_r_3_23 ) );
  DFF_X1 key_b_r_reg_3_24 (.CK( clk ) , .D( key_b_r_2_24 ) , .Q( key_b_r_3_24 ) );
  DFF_X1 key_b_r_reg_3_25 (.CK( clk ) , .D( key_b_r_2_25 ) , .Q( key_b_r_3_25 ) );
  DFF_X1 key_b_r_reg_3_26 (.CK( clk ) , .D( key_b_r_2_26 ) , .Q( key_b_r_3_26 ) );
  DFF_X1 key_b_r_reg_3_27 (.CK( clk ) , .D( key_b_r_2_27 ) , .Q( key_b_r_3_27 ) );
  DFF_X1 key_b_r_reg_3_28 (.CK( clk ) , .D( key_b_r_2_28 ) , .Q( key_b_r_3_28 ) );
  DFF_X1 key_b_r_reg_3_29 (.CK( clk ) , .D( key_b_r_2_29 ) , .Q( key_b_r_3_29 ) );
  DFF_X1 key_b_r_reg_3_3 (.CK( clk ) , .D( key_b_r_2_3 ) , .Q( key_b_r_3_3 ) );
  DFF_X1 key_b_r_reg_3_30 (.CK( clk ) , .D( key_b_r_2_30 ) , .Q( key_b_r_3_30 ) );
  DFF_X1 key_b_r_reg_3_31 (.CK( clk ) , .D( key_b_r_2_31 ) , .Q( key_b_r_3_31 ) );
  DFF_X1 key_b_r_reg_3_32 (.CK( clk ) , .D( key_b_r_2_32 ) , .Q( key_b_r_3_32 ) );
  DFF_X1 key_b_r_reg_3_33 (.CK( clk ) , .D( key_b_r_2_33 ) , .Q( key_b_r_3_33 ) );
  DFF_X1 key_b_r_reg_3_34 (.CK( clk ) , .D( key_b_r_2_34 ) , .Q( key_b_r_3_34 ) );
  DFF_X1 key_b_r_reg_3_35 (.CK( clk ) , .D( key_b_r_2_35 ) , .Q( key_b_r_3_35 ) );
  DFF_X1 key_b_r_reg_3_36 (.CK( clk ) , .D( key_b_r_2_36 ) , .Q( key_b_r_3_36 ) );
  DFF_X1 key_b_r_reg_3_37 (.CK( clk ) , .D( key_b_r_2_37 ) , .Q( key_b_r_3_37 ) );
  DFF_X1 key_b_r_reg_3_38 (.CK( clk ) , .D( key_b_r_2_38 ) , .Q( key_b_r_3_38 ) );
  DFF_X1 key_b_r_reg_3_39 (.CK( clk ) , .D( key_b_r_2_39 ) , .Q( key_b_r_3_39 ) );
  DFF_X1 key_b_r_reg_3_4 (.CK( clk ) , .D( key_b_r_2_4 ) , .Q( key_b_r_3_4 ) );
  DFF_X1 key_b_r_reg_3_40 (.CK( clk ) , .D( key_b_r_2_40 ) , .Q( key_b_r_3_40 ) );
  DFF_X1 key_b_r_reg_3_41 (.CK( clk ) , .D( key_b_r_2_41 ) , .Q( key_b_r_3_41 ) );
  DFF_X1 key_b_r_reg_3_42 (.CK( clk ) , .D( key_b_r_2_42 ) , .Q( key_b_r_3_42 ) );
  DFF_X1 key_b_r_reg_3_43 (.CK( clk ) , .D( key_b_r_2_43 ) , .Q( key_b_r_3_43 ) );
  DFF_X1 key_b_r_reg_3_44 (.CK( clk ) , .D( key_b_r_2_44 ) , .Q( key_b_r_3_44 ) );
  DFF_X1 key_b_r_reg_3_45 (.CK( clk ) , .D( key_b_r_2_45 ) , .Q( key_b_r_3_45 ) );
  DFF_X1 key_b_r_reg_3_46 (.CK( clk ) , .D( key_b_r_2_46 ) , .Q( key_b_r_3_46 ) );
  DFF_X1 key_b_r_reg_3_47 (.CK( clk ) , .D( key_b_r_2_47 ) , .Q( key_b_r_3_47 ) );
  DFF_X1 key_b_r_reg_3_48 (.CK( clk ) , .D( key_b_r_2_48 ) , .Q( key_b_r_3_48 ) );
  DFF_X1 key_b_r_reg_3_49 (.CK( clk ) , .D( key_b_r_2_49 ) , .Q( key_b_r_3_49 ) );
  DFF_X1 key_b_r_reg_3_5 (.CK( clk ) , .D( key_b_r_2_5 ) , .Q( key_b_r_3_5 ) );
  DFF_X1 key_b_r_reg_3_50 (.CK( clk ) , .D( key_b_r_2_50 ) , .Q( key_b_r_3_50 ) );
  DFF_X1 key_b_r_reg_3_51 (.CK( clk ) , .D( key_b_r_2_51 ) , .Q( key_b_r_3_51 ) );
  DFF_X1 key_b_r_reg_3_52 (.CK( clk ) , .D( key_b_r_2_52 ) , .Q( key_b_r_3_52 ) );
  DFF_X1 key_b_r_reg_3_53 (.CK( clk ) , .D( key_b_r_2_53 ) , .Q( key_b_r_3_53 ) );
  DFF_X1 key_b_r_reg_3_54 (.CK( clk ) , .D( key_b_r_2_54 ) , .Q( key_b_r_3_54 ) );
  DFF_X1 key_b_r_reg_3_55 (.CK( clk ) , .D( key_b_r_2_55 ) , .Q( key_b_r_3_55 ) );
  DFF_X1 key_b_r_reg_3_6 (.CK( clk ) , .D( key_b_r_2_6 ) , .Q( key_b_r_3_6 ) );
  DFF_X1 key_b_r_reg_3_7 (.CK( clk ) , .D( key_b_r_2_7 ) , .Q( key_b_r_3_7 ) );
  DFF_X1 key_b_r_reg_3_8 (.CK( clk ) , .D( key_b_r_2_8 ) , .Q( key_b_r_3_8 ) );
  DFF_X1 key_b_r_reg_3_9 (.CK( clk ) , .D( key_b_r_2_9 ) , .Q( key_b_r_3_9 ) );
  DFF_X1 key_b_r_reg_4_0 (.CK( clk ) , .D( key_b_r_3_0 ) , .Q( key_b_r_4_0 ) );
  DFF_X1 key_b_r_reg_4_1 (.CK( clk ) , .D( key_b_r_3_1 ) , .Q( key_b_r_4_1 ) );
  DFF_X1 key_b_r_reg_4_10 (.CK( clk ) , .D( key_b_r_3_10 ) , .Q( key_b_r_4_10 ) );
  DFF_X1 key_b_r_reg_4_11 (.CK( clk ) , .D( key_b_r_3_11 ) , .Q( key_b_r_4_11 ) );
  DFF_X1 key_b_r_reg_4_12 (.CK( clk ) , .D( key_b_r_3_12 ) , .Q( key_b_r_4_12 ) );
  DFF_X1 key_b_r_reg_4_13 (.CK( clk ) , .D( key_b_r_3_13 ) , .Q( key_b_r_4_13 ) );
  DFF_X1 key_b_r_reg_4_14 (.CK( clk ) , .D( key_b_r_3_14 ) , .Q( key_b_r_4_14 ) );
  DFF_X1 key_b_r_reg_4_15 (.CK( clk ) , .D( key_b_r_3_15 ) , .Q( key_b_r_4_15 ) );
  DFF_X1 key_b_r_reg_4_16 (.CK( clk ) , .D( key_b_r_3_16 ) , .Q( key_b_r_4_16 ) );
  DFF_X1 key_b_r_reg_4_17 (.CK( clk ) , .D( key_b_r_3_17 ) , .Q( key_b_r_4_17 ) );
  DFF_X1 key_b_r_reg_4_18 (.CK( clk ) , .D( key_b_r_3_18 ) , .Q( key_b_r_4_18 ) );
  DFF_X1 key_b_r_reg_4_19 (.CK( clk ) , .D( key_b_r_3_19 ) , .Q( key_b_r_4_19 ) );
  DFF_X1 key_b_r_reg_4_2 (.CK( clk ) , .D( key_b_r_3_2 ) , .Q( key_b_r_4_2 ) );
  DFF_X1 key_b_r_reg_4_20 (.CK( clk ) , .D( key_b_r_3_20 ) , .Q( key_b_r_4_20 ) );
  DFF_X1 key_b_r_reg_4_21 (.CK( clk ) , .D( key_b_r_3_21 ) , .Q( key_b_r_4_21 ) );
  DFF_X1 key_b_r_reg_4_22 (.CK( clk ) , .D( key_b_r_3_22 ) , .Q( key_b_r_4_22 ) );
  DFF_X1 key_b_r_reg_4_23 (.CK( clk ) , .D( key_b_r_3_23 ) , .Q( key_b_r_4_23 ) );
  DFF_X1 key_b_r_reg_4_24 (.CK( clk ) , .D( key_b_r_3_24 ) , .Q( key_b_r_4_24 ) );
  DFF_X1 key_b_r_reg_4_25 (.CK( clk ) , .D( key_b_r_3_25 ) , .Q( key_b_r_4_25 ) );
  DFF_X1 key_b_r_reg_4_26 (.CK( clk ) , .D( key_b_r_3_26 ) , .Q( key_b_r_4_26 ) );
  DFF_X1 key_b_r_reg_4_27 (.CK( clk ) , .D( key_b_r_3_27 ) , .Q( key_b_r_4_27 ) );
  DFF_X1 key_b_r_reg_4_28 (.CK( clk ) , .D( key_b_r_3_28 ) , .Q( key_b_r_4_28 ) );
  DFF_X1 key_b_r_reg_4_29 (.CK( clk ) , .D( key_b_r_3_29 ) , .Q( key_b_r_4_29 ) );
  DFF_X1 key_b_r_reg_4_3 (.CK( clk ) , .D( key_b_r_3_3 ) , .Q( key_b_r_4_3 ) );
  DFF_X1 key_b_r_reg_4_30 (.CK( clk ) , .D( key_b_r_3_30 ) , .Q( key_b_r_4_30 ) );
  DFF_X1 key_b_r_reg_4_31 (.CK( clk ) , .D( key_b_r_3_31 ) , .Q( key_b_r_4_31 ) );
  DFF_X1 key_b_r_reg_4_32 (.CK( clk ) , .D( key_b_r_3_32 ) , .Q( key_b_r_4_32 ) );
  DFF_X1 key_b_r_reg_4_33 (.CK( clk ) , .D( key_b_r_3_33 ) , .Q( key_b_r_4_33 ) );
  DFF_X1 key_b_r_reg_4_34 (.CK( clk ) , .D( key_b_r_3_34 ) , .Q( key_b_r_4_34 ) );
  DFF_X1 key_b_r_reg_4_35 (.CK( clk ) , .D( key_b_r_3_35 ) , .Q( key_b_r_4_35 ) );
  DFF_X1 key_b_r_reg_4_36 (.CK( clk ) , .D( key_b_r_3_36 ) , .Q( key_b_r_4_36 ) );
  DFF_X1 key_b_r_reg_4_37 (.CK( clk ) , .D( key_b_r_3_37 ) , .Q( key_b_r_4_37 ) );
  DFF_X1 key_b_r_reg_4_38 (.CK( clk ) , .D( key_b_r_3_38 ) , .Q( key_b_r_4_38 ) );
  DFF_X1 key_b_r_reg_4_39 (.CK( clk ) , .D( key_b_r_3_39 ) , .Q( key_b_r_4_39 ) );
  DFF_X1 key_b_r_reg_4_4 (.CK( clk ) , .D( key_b_r_3_4 ) , .Q( key_b_r_4_4 ) );
  DFF_X1 key_b_r_reg_4_40 (.CK( clk ) , .D( key_b_r_3_40 ) , .Q( key_b_r_4_40 ) );
  DFF_X1 key_b_r_reg_4_41 (.CK( clk ) , .D( key_b_r_3_41 ) , .Q( key_b_r_4_41 ) );
  DFF_X1 key_b_r_reg_4_42 (.CK( clk ) , .D( key_b_r_3_42 ) , .Q( key_b_r_4_42 ) );
  DFF_X1 key_b_r_reg_4_43 (.CK( clk ) , .D( key_b_r_3_43 ) , .Q( key_b_r_4_43 ) );
  DFF_X1 key_b_r_reg_4_44 (.CK( clk ) , .D( key_b_r_3_44 ) , .Q( key_b_r_4_44 ) );
  DFF_X1 key_b_r_reg_4_45 (.CK( clk ) , .D( key_b_r_3_45 ) , .Q( key_b_r_4_45 ) );
  DFF_X1 key_b_r_reg_4_46 (.CK( clk ) , .D( key_b_r_3_46 ) , .Q( key_b_r_4_46 ) );
  DFF_X1 key_b_r_reg_4_47 (.CK( clk ) , .D( key_b_r_3_47 ) , .Q( key_b_r_4_47 ) );
  DFF_X1 key_b_r_reg_4_48 (.CK( clk ) , .D( key_b_r_3_48 ) , .Q( key_b_r_4_48 ) );
  DFF_X1 key_b_r_reg_4_49 (.CK( clk ) , .D( key_b_r_3_49 ) , .Q( key_b_r_4_49 ) );
  DFF_X1 key_b_r_reg_4_5 (.CK( clk ) , .D( key_b_r_3_5 ) , .Q( key_b_r_4_5 ) );
  DFF_X1 key_b_r_reg_4_50 (.CK( clk ) , .D( key_b_r_3_50 ) , .Q( key_b_r_4_50 ) );
  DFF_X1 key_b_r_reg_4_51 (.CK( clk ) , .D( key_b_r_3_51 ) , .Q( key_b_r_4_51 ) );
  DFF_X1 key_b_r_reg_4_52 (.CK( clk ) , .D( key_b_r_3_52 ) , .Q( key_b_r_4_52 ) );
  DFF_X1 key_b_r_reg_4_53 (.CK( clk ) , .D( key_b_r_3_53 ) , .Q( key_b_r_4_53 ) );
  DFF_X1 key_b_r_reg_4_54 (.CK( clk ) , .D( key_b_r_3_54 ) , .Q( key_b_r_4_54 ) );
  DFF_X1 key_b_r_reg_4_55 (.CK( clk ) , .D( key_b_r_3_55 ) , .Q( key_b_r_4_55 ) );
  DFF_X1 key_b_r_reg_4_6 (.CK( clk ) , .D( key_b_r_3_6 ) , .Q( key_b_r_4_6 ) );
  DFF_X1 key_b_r_reg_4_7 (.CK( clk ) , .D( key_b_r_3_7 ) , .Q( key_b_r_4_7 ) );
  DFF_X1 key_b_r_reg_4_8 (.CK( clk ) , .D( key_b_r_3_8 ) , .Q( key_b_r_4_8 ) );
  DFF_X1 key_b_r_reg_4_9 (.CK( clk ) , .D( key_b_r_3_9 ) , .Q( key_b_r_4_9 ) );
  DFF_X1 key_b_r_reg_5_0 (.CK( clk ) , .D( key_b_r_4_0 ) , .Q( key_b_r_5_0 ) );
  DFF_X1 key_b_r_reg_5_1 (.CK( clk ) , .D( key_b_r_4_1 ) , .Q( key_b_r_5_1 ) );
  DFF_X1 key_b_r_reg_5_10 (.CK( clk ) , .D( key_b_r_4_10 ) , .Q( key_b_r_5_10 ) );
  DFF_X1 key_b_r_reg_5_11 (.CK( clk ) , .D( key_b_r_4_11 ) , .Q( key_b_r_5_11 ) );
  DFF_X1 key_b_r_reg_5_12 (.CK( clk ) , .D( key_b_r_4_12 ) , .Q( key_b_r_5_12 ) );
  DFF_X1 key_b_r_reg_5_13 (.CK( clk ) , .D( key_b_r_4_13 ) , .Q( key_b_r_5_13 ) );
  DFF_X1 key_b_r_reg_5_14 (.CK( clk ) , .D( key_b_r_4_14 ) , .Q( key_b_r_5_14 ) );
  DFF_X1 key_b_r_reg_5_15 (.CK( clk ) , .D( key_b_r_4_15 ) , .Q( key_b_r_5_15 ) );
  DFF_X1 key_b_r_reg_5_16 (.CK( clk ) , .D( key_b_r_4_16 ) , .Q( key_b_r_5_16 ) );
  DFF_X1 key_b_r_reg_5_17 (.CK( clk ) , .D( key_b_r_4_17 ) , .Q( key_b_r_5_17 ) );
  DFF_X1 key_b_r_reg_5_18 (.CK( clk ) , .D( key_b_r_4_18 ) , .Q( key_b_r_5_18 ) );
  DFF_X1 key_b_r_reg_5_19 (.CK( clk ) , .D( key_b_r_4_19 ) , .Q( key_b_r_5_19 ) );
  DFF_X1 key_b_r_reg_5_2 (.CK( clk ) , .D( key_b_r_4_2 ) , .Q( key_b_r_5_2 ) );
  DFF_X1 key_b_r_reg_5_20 (.CK( clk ) , .D( key_b_r_4_20 ) , .Q( key_b_r_5_20 ) );
  DFF_X1 key_b_r_reg_5_21 (.CK( clk ) , .D( key_b_r_4_21 ) , .Q( key_b_r_5_21 ) );
  DFF_X1 key_b_r_reg_5_22 (.CK( clk ) , .D( key_b_r_4_22 ) , .Q( key_b_r_5_22 ) );
  DFF_X1 key_b_r_reg_5_23 (.CK( clk ) , .D( key_b_r_4_23 ) , .Q( key_b_r_5_23 ) );
  DFF_X1 key_b_r_reg_5_24 (.CK( clk ) , .D( key_b_r_4_24 ) , .Q( key_b_r_5_24 ) );
  DFF_X1 key_b_r_reg_5_25 (.CK( clk ) , .D( key_b_r_4_25 ) , .Q( key_b_r_5_25 ) );
  DFF_X1 key_b_r_reg_5_26 (.CK( clk ) , .D( key_b_r_4_26 ) , .Q( key_b_r_5_26 ) );
  DFF_X1 key_b_r_reg_5_27 (.CK( clk ) , .D( key_b_r_4_27 ) , .Q( key_b_r_5_27 ) );
  DFF_X1 key_b_r_reg_5_28 (.CK( clk ) , .D( key_b_r_4_28 ) , .Q( key_b_r_5_28 ) );
  DFF_X1 key_b_r_reg_5_29 (.CK( clk ) , .D( key_b_r_4_29 ) , .Q( key_b_r_5_29 ) );
  DFF_X1 key_b_r_reg_5_3 (.CK( clk ) , .D( key_b_r_4_3 ) , .Q( key_b_r_5_3 ) );
  DFF_X1 key_b_r_reg_5_30 (.CK( clk ) , .D( key_b_r_4_30 ) , .Q( key_b_r_5_30 ) );
  DFF_X1 key_b_r_reg_5_31 (.CK( clk ) , .D( key_b_r_4_31 ) , .Q( key_b_r_5_31 ) );
  DFF_X1 key_b_r_reg_5_32 (.CK( clk ) , .D( key_b_r_4_32 ) , .Q( key_b_r_5_32 ) );
  DFF_X1 key_b_r_reg_5_33 (.CK( clk ) , .D( key_b_r_4_33 ) , .Q( key_b_r_5_33 ) );
  DFF_X1 key_b_r_reg_5_34 (.CK( clk ) , .D( key_b_r_4_34 ) , .Q( key_b_r_5_34 ) );
  DFF_X1 key_b_r_reg_5_35 (.CK( clk ) , .D( key_b_r_4_35 ) , .Q( key_b_r_5_35 ) );
  DFF_X1 key_b_r_reg_5_36 (.CK( clk ) , .D( key_b_r_4_36 ) , .Q( key_b_r_5_36 ) );
  DFF_X1 key_b_r_reg_5_37 (.CK( clk ) , .D( key_b_r_4_37 ) , .Q( key_b_r_5_37 ) );
  DFF_X1 key_b_r_reg_5_38 (.CK( clk ) , .D( key_b_r_4_38 ) , .Q( key_b_r_5_38 ) );
  DFF_X1 key_b_r_reg_5_39 (.CK( clk ) , .D( key_b_r_4_39 ) , .Q( key_b_r_5_39 ) );
  DFF_X1 key_b_r_reg_5_4 (.CK( clk ) , .D( key_b_r_4_4 ) , .Q( key_b_r_5_4 ) );
  DFF_X1 key_b_r_reg_5_40 (.CK( clk ) , .D( key_b_r_4_40 ) , .Q( key_b_r_5_40 ) );
  DFF_X1 key_b_r_reg_5_41 (.CK( clk ) , .D( key_b_r_4_41 ) , .Q( key_b_r_5_41 ) );
  DFF_X1 key_b_r_reg_5_42 (.CK( clk ) , .D( key_b_r_4_42 ) , .Q( key_b_r_5_42 ) );
  DFF_X1 key_b_r_reg_5_43 (.CK( clk ) , .D( key_b_r_4_43 ) , .Q( key_b_r_5_43 ) );
  DFF_X1 key_b_r_reg_5_44 (.CK( clk ) , .D( key_b_r_4_44 ) , .Q( key_b_r_5_44 ) );
  DFF_X1 key_b_r_reg_5_45 (.CK( clk ) , .D( key_b_r_4_45 ) , .Q( key_b_r_5_45 ) );
  DFF_X1 key_b_r_reg_5_46 (.CK( clk ) , .D( key_b_r_4_46 ) , .Q( key_b_r_5_46 ) );
  DFF_X1 key_b_r_reg_5_47 (.CK( clk ) , .D( key_b_r_4_47 ) , .Q( key_b_r_5_47 ) );
  DFF_X1 key_b_r_reg_5_48 (.CK( clk ) , .D( key_b_r_4_48 ) , .Q( key_b_r_5_48 ) );
  DFF_X1 key_b_r_reg_5_49 (.CK( clk ) , .D( key_b_r_4_49 ) , .Q( key_b_r_5_49 ) );
  DFF_X1 key_b_r_reg_5_5 (.CK( clk ) , .D( key_b_r_4_5 ) , .Q( key_b_r_5_5 ) );
  DFF_X1 key_b_r_reg_5_50 (.CK( clk ) , .D( key_b_r_4_50 ) , .Q( key_b_r_5_50 ) );
  DFF_X1 key_b_r_reg_5_51 (.CK( clk ) , .D( key_b_r_4_51 ) , .Q( key_b_r_5_51 ) );
  DFF_X1 key_b_r_reg_5_52 (.CK( clk ) , .D( key_b_r_4_52 ) , .Q( key_b_r_5_52 ) );
  DFF_X1 key_b_r_reg_5_53 (.CK( clk ) , .D( key_b_r_4_53 ) , .Q( key_b_r_5_53 ) );
  DFF_X1 key_b_r_reg_5_54 (.CK( clk ) , .D( key_b_r_4_54 ) , .Q( key_b_r_5_54 ) );
  DFF_X1 key_b_r_reg_5_55 (.CK( clk ) , .D( key_b_r_4_55 ) , .Q( key_b_r_5_55 ) );
  DFF_X1 key_b_r_reg_5_6 (.CK( clk ) , .D( key_b_r_4_6 ) , .Q( key_b_r_5_6 ) );
  DFF_X1 key_b_r_reg_5_7 (.CK( clk ) , .D( key_b_r_4_7 ) , .Q( key_b_r_5_7 ) );
  DFF_X1 key_b_r_reg_5_8 (.CK( clk ) , .D( key_b_r_4_8 ) , .Q( key_b_r_5_8 ) );
  DFF_X1 key_b_r_reg_5_9 (.CK( clk ) , .D( key_b_r_4_9 ) , .Q( key_b_r_5_9 ) );
  DFF_X1 key_b_r_reg_6_0 (.CK( clk ) , .D( key_b_r_5_0 ) , .Q( key_b_r_6_0 ) );
  DFF_X1 key_b_r_reg_6_1 (.CK( clk ) , .D( key_b_r_5_1 ) , .Q( key_b_r_6_1 ) );
  DFF_X1 key_b_r_reg_6_10 (.CK( clk ) , .D( key_b_r_5_10 ) , .Q( key_b_r_6_10 ) );
  DFF_X1 key_b_r_reg_6_11 (.CK( clk ) , .D( key_b_r_5_11 ) , .Q( key_b_r_6_11 ) );
  DFF_X1 key_b_r_reg_6_12 (.CK( clk ) , .D( key_b_r_5_12 ) , .Q( key_b_r_6_12 ) );
  DFF_X1 key_b_r_reg_6_13 (.CK( clk ) , .D( key_b_r_5_13 ) , .Q( key_b_r_6_13 ) );
  DFF_X1 key_b_r_reg_6_14 (.CK( clk ) , .D( key_b_r_5_14 ) , .Q( key_b_r_6_14 ) );
  DFF_X1 key_b_r_reg_6_15 (.CK( clk ) , .D( key_b_r_5_15 ) , .Q( key_b_r_6_15 ) );
  DFF_X1 key_b_r_reg_6_16 (.CK( clk ) , .D( key_b_r_5_16 ) , .Q( key_b_r_6_16 ) );
  DFF_X1 key_b_r_reg_6_17 (.CK( clk ) , .D( key_b_r_5_17 ) , .Q( key_b_r_6_17 ) );
  DFF_X1 key_b_r_reg_6_18 (.CK( clk ) , .D( key_b_r_5_18 ) , .Q( key_b_r_6_18 ) );
  DFF_X1 key_b_r_reg_6_19 (.CK( clk ) , .D( key_b_r_5_19 ) , .Q( key_b_r_6_19 ) );
  DFF_X1 key_b_r_reg_6_2 (.CK( clk ) , .D( key_b_r_5_2 ) , .Q( key_b_r_6_2 ) );
  DFF_X1 key_b_r_reg_6_20 (.CK( clk ) , .D( key_b_r_5_20 ) , .Q( key_b_r_6_20 ) );
  DFF_X1 key_b_r_reg_6_21 (.CK( clk ) , .D( key_b_r_5_21 ) , .Q( key_b_r_6_21 ) );
  DFF_X1 key_b_r_reg_6_22 (.CK( clk ) , .D( key_b_r_5_22 ) , .Q( key_b_r_6_22 ) );
  DFF_X1 key_b_r_reg_6_23 (.CK( clk ) , .D( key_b_r_5_23 ) , .Q( key_b_r_6_23 ) );
  DFF_X1 key_b_r_reg_6_24 (.CK( clk ) , .D( key_b_r_5_24 ) , .Q( key_b_r_6_24 ) );
  DFF_X1 key_b_r_reg_6_25 (.CK( clk ) , .D( key_b_r_5_25 ) , .Q( key_b_r_6_25 ) );
  DFF_X1 key_b_r_reg_6_26 (.CK( clk ) , .D( key_b_r_5_26 ) , .Q( key_b_r_6_26 ) );
  DFF_X1 key_b_r_reg_6_27 (.CK( clk ) , .D( key_b_r_5_27 ) , .Q( key_b_r_6_27 ) );
  DFF_X1 key_b_r_reg_6_28 (.CK( clk ) , .D( key_b_r_5_28 ) , .Q( key_b_r_6_28 ) );
  DFF_X1 key_b_r_reg_6_29 (.CK( clk ) , .D( key_b_r_5_29 ) , .Q( key_b_r_6_29 ) );
  DFF_X1 key_b_r_reg_6_3 (.CK( clk ) , .D( key_b_r_5_3 ) , .Q( key_b_r_6_3 ) );
  DFF_X1 key_b_r_reg_6_30 (.CK( clk ) , .D( key_b_r_5_30 ) , .Q( key_b_r_6_30 ) );
  DFF_X1 key_b_r_reg_6_31 (.CK( clk ) , .D( key_b_r_5_31 ) , .Q( key_b_r_6_31 ) );
  DFF_X1 key_b_r_reg_6_32 (.CK( clk ) , .D( key_b_r_5_32 ) , .Q( key_b_r_6_32 ) );
  DFF_X1 key_b_r_reg_6_33 (.CK( clk ) , .D( key_b_r_5_33 ) , .Q( key_b_r_6_33 ) );
  DFF_X1 key_b_r_reg_6_34 (.CK( clk ) , .D( key_b_r_5_34 ) , .Q( key_b_r_6_34 ) );
  DFF_X1 key_b_r_reg_6_35 (.CK( clk ) , .D( key_b_r_5_35 ) , .Q( key_b_r_6_35 ) );
  DFF_X1 key_b_r_reg_6_36 (.CK( clk ) , .D( key_b_r_5_36 ) , .Q( key_b_r_6_36 ) );
  DFF_X1 key_b_r_reg_6_37 (.CK( clk ) , .D( key_b_r_5_37 ) , .Q( key_b_r_6_37 ) );
  DFF_X1 key_b_r_reg_6_38 (.CK( clk ) , .D( key_b_r_5_38 ) , .Q( key_b_r_6_38 ) );
  DFF_X1 key_b_r_reg_6_39 (.CK( clk ) , .D( key_b_r_5_39 ) , .Q( key_b_r_6_39 ) );
  DFF_X1 key_b_r_reg_6_4 (.CK( clk ) , .D( key_b_r_5_4 ) , .Q( key_b_r_6_4 ) );
  DFF_X1 key_b_r_reg_6_40 (.CK( clk ) , .D( key_b_r_5_40 ) , .Q( key_b_r_6_40 ) );
  DFF_X1 key_b_r_reg_6_41 (.CK( clk ) , .D( key_b_r_5_41 ) , .Q( key_b_r_6_41 ) );
  DFF_X1 key_b_r_reg_6_42 (.CK( clk ) , .D( key_b_r_5_42 ) , .Q( key_b_r_6_42 ) );
  DFF_X1 key_b_r_reg_6_43 (.CK( clk ) , .D( key_b_r_5_43 ) , .Q( key_b_r_6_43 ) );
  DFF_X1 key_b_r_reg_6_44 (.CK( clk ) , .D( key_b_r_5_44 ) , .Q( key_b_r_6_44 ) );
  DFF_X1 key_b_r_reg_6_45 (.CK( clk ) , .D( key_b_r_5_45 ) , .Q( key_b_r_6_45 ) );
  DFF_X1 key_b_r_reg_6_46 (.CK( clk ) , .D( key_b_r_5_46 ) , .Q( key_b_r_6_46 ) );
  DFF_X1 key_b_r_reg_6_47 (.CK( clk ) , .D( key_b_r_5_47 ) , .Q( key_b_r_6_47 ) );
  DFF_X1 key_b_r_reg_6_48 (.CK( clk ) , .D( key_b_r_5_48 ) , .Q( key_b_r_6_48 ) );
  DFF_X1 key_b_r_reg_6_49 (.CK( clk ) , .D( key_b_r_5_49 ) , .Q( key_b_r_6_49 ) );
  DFF_X1 key_b_r_reg_6_5 (.CK( clk ) , .D( key_b_r_5_5 ) , .Q( key_b_r_6_5 ) );
  DFF_X1 key_b_r_reg_6_50 (.CK( clk ) , .D( key_b_r_5_50 ) , .Q( key_b_r_6_50 ) );
  DFF_X1 key_b_r_reg_6_51 (.CK( clk ) , .D( key_b_r_5_51 ) , .Q( key_b_r_6_51 ) );
  DFF_X1 key_b_r_reg_6_52 (.CK( clk ) , .D( key_b_r_5_52 ) , .Q( key_b_r_6_52 ) );
  DFF_X1 key_b_r_reg_6_53 (.CK( clk ) , .D( key_b_r_5_53 ) , .Q( key_b_r_6_53 ) );
  DFF_X1 key_b_r_reg_6_54 (.CK( clk ) , .D( key_b_r_5_54 ) , .Q( key_b_r_6_54 ) );
  DFF_X1 key_b_r_reg_6_55 (.CK( clk ) , .D( key_b_r_5_55 ) , .Q( key_b_r_6_55 ) );
  DFF_X1 key_b_r_reg_6_6 (.CK( clk ) , .D( key_b_r_5_6 ) , .Q( key_b_r_6_6 ) );
  DFF_X1 key_b_r_reg_6_7 (.CK( clk ) , .D( key_b_r_5_7 ) , .Q( key_b_r_6_7 ) );
  DFF_X1 key_b_r_reg_6_8 (.CK( clk ) , .D( key_b_r_5_8 ) , .Q( key_b_r_6_8 ) );
  DFF_X1 key_b_r_reg_6_9 (.CK( clk ) , .D( key_b_r_5_9 ) , .Q( key_b_r_6_9 ) );
  DFF_X1 key_b_r_reg_7_0 (.CK( clk ) , .D( key_b_r_6_0 ) , .Q( key_b_r_7_0 ) );
  DFF_X1 key_b_r_reg_7_1 (.CK( clk ) , .D( key_b_r_6_1 ) , .Q( key_b_r_7_1 ) );
  DFF_X1 key_b_r_reg_7_10 (.CK( clk ) , .D( key_b_r_6_10 ) , .Q( key_b_r_7_10 ) );
  DFF_X1 key_b_r_reg_7_11 (.CK( clk ) , .D( key_b_r_6_11 ) , .Q( key_b_r_7_11 ) );
  DFF_X1 key_b_r_reg_7_12 (.CK( clk ) , .D( key_b_r_6_12 ) , .Q( key_b_r_7_12 ) );
  DFF_X1 key_b_r_reg_7_13 (.CK( clk ) , .D( key_b_r_6_13 ) , .Q( key_b_r_7_13 ) );
  DFF_X1 key_b_r_reg_7_14 (.CK( clk ) , .D( key_b_r_6_14 ) , .Q( key_b_r_7_14 ) );
  DFF_X1 key_b_r_reg_7_15 (.CK( clk ) , .D( key_b_r_6_15 ) , .Q( key_b_r_7_15 ) );
  DFF_X1 key_b_r_reg_7_16 (.CK( clk ) , .D( key_b_r_6_16 ) , .Q( key_b_r_7_16 ) );
  DFF_X1 key_b_r_reg_7_17 (.CK( clk ) , .D( key_b_r_6_17 ) , .Q( key_b_r_7_17 ) );
  DFF_X1 key_b_r_reg_7_18 (.CK( clk ) , .D( key_b_r_6_18 ) , .Q( key_b_r_7_18 ) );
  DFF_X1 key_b_r_reg_7_19 (.CK( clk ) , .D( key_b_r_6_19 ) , .Q( key_b_r_7_19 ) );
  DFF_X1 key_b_r_reg_7_2 (.CK( clk ) , .D( key_b_r_6_2 ) , .Q( key_b_r_7_2 ) );
  DFF_X1 key_b_r_reg_7_20 (.CK( clk ) , .D( key_b_r_6_20 ) , .Q( key_b_r_7_20 ) );
  DFF_X1 key_b_r_reg_7_21 (.CK( clk ) , .D( key_b_r_6_21 ) , .Q( key_b_r_7_21 ) );
  DFF_X1 key_b_r_reg_7_22 (.CK( clk ) , .D( key_b_r_6_22 ) , .Q( key_b_r_7_22 ) );
  DFF_X1 key_b_r_reg_7_23 (.CK( clk ) , .D( key_b_r_6_23 ) , .Q( key_b_r_7_23 ) );
  DFF_X1 key_b_r_reg_7_24 (.CK( clk ) , .D( key_b_r_6_24 ) , .Q( key_b_r_7_24 ) );
  DFF_X1 key_b_r_reg_7_25 (.CK( clk ) , .D( key_b_r_6_25 ) , .Q( key_b_r_7_25 ) );
  DFF_X1 key_b_r_reg_7_26 (.CK( clk ) , .D( key_b_r_6_26 ) , .Q( key_b_r_7_26 ) );
  DFF_X1 key_b_r_reg_7_27 (.CK( clk ) , .D( key_b_r_6_27 ) , .Q( key_b_r_7_27 ) );
  DFF_X1 key_b_r_reg_7_28 (.CK( clk ) , .D( key_b_r_6_28 ) , .Q( key_b_r_7_28 ) );
  DFF_X1 key_b_r_reg_7_29 (.CK( clk ) , .D( key_b_r_6_29 ) , .Q( key_b_r_7_29 ) );
  DFF_X1 key_b_r_reg_7_3 (.CK( clk ) , .D( key_b_r_6_3 ) , .Q( key_b_r_7_3 ) );
  DFF_X1 key_b_r_reg_7_30 (.CK( clk ) , .D( key_b_r_6_30 ) , .Q( key_b_r_7_30 ) );
  DFF_X1 key_b_r_reg_7_31 (.CK( clk ) , .D( key_b_r_6_31 ) , .Q( key_b_r_7_31 ) );
  DFF_X1 key_b_r_reg_7_32 (.CK( clk ) , .D( key_b_r_6_32 ) , .Q( key_b_r_7_32 ) );
  DFF_X1 key_b_r_reg_7_33 (.CK( clk ) , .D( key_b_r_6_33 ) , .Q( key_b_r_7_33 ) );
  DFF_X1 key_b_r_reg_7_34 (.CK( clk ) , .D( key_b_r_6_34 ) , .Q( key_b_r_7_34 ) );
  DFF_X1 key_b_r_reg_7_35 (.CK( clk ) , .D( key_b_r_6_35 ) , .Q( key_b_r_7_35 ) );
  DFF_X1 key_b_r_reg_7_36 (.CK( clk ) , .D( key_b_r_6_36 ) , .Q( key_b_r_7_36 ) );
  DFF_X1 key_b_r_reg_7_37 (.CK( clk ) , .D( key_b_r_6_37 ) , .Q( key_b_r_7_37 ) );
  DFF_X1 key_b_r_reg_7_38 (.CK( clk ) , .D( key_b_r_6_38 ) , .Q( key_b_r_7_38 ) );
  DFF_X1 key_b_r_reg_7_39 (.CK( clk ) , .D( key_b_r_6_39 ) , .Q( key_b_r_7_39 ) );
  DFF_X1 key_b_r_reg_7_4 (.CK( clk ) , .D( key_b_r_6_4 ) , .Q( key_b_r_7_4 ) );
  DFF_X1 key_b_r_reg_7_40 (.CK( clk ) , .D( key_b_r_6_40 ) , .Q( key_b_r_7_40 ) );
  DFF_X1 key_b_r_reg_7_41 (.CK( clk ) , .D( key_b_r_6_41 ) , .Q( key_b_r_7_41 ) );
  DFF_X1 key_b_r_reg_7_42 (.CK( clk ) , .D( key_b_r_6_42 ) , .Q( key_b_r_7_42 ) );
  DFF_X1 key_b_r_reg_7_43 (.CK( clk ) , .D( key_b_r_6_43 ) , .Q( key_b_r_7_43 ) );
  DFF_X1 key_b_r_reg_7_44 (.CK( clk ) , .D( key_b_r_6_44 ) , .Q( key_b_r_7_44 ) );
  DFF_X1 key_b_r_reg_7_45 (.CK( clk ) , .D( key_b_r_6_45 ) , .Q( key_b_r_7_45 ) );
  DFF_X1 key_b_r_reg_7_46 (.CK( clk ) , .D( key_b_r_6_46 ) , .Q( key_b_r_7_46 ) );
  DFF_X1 key_b_r_reg_7_47 (.CK( clk ) , .D( key_b_r_6_47 ) , .Q( key_b_r_7_47 ) );
  DFF_X1 key_b_r_reg_7_48 (.CK( clk ) , .D( key_b_r_6_48 ) , .Q( key_b_r_7_48 ) );
  DFF_X1 key_b_r_reg_7_49 (.CK( clk ) , .D( key_b_r_6_49 ) , .Q( key_b_r_7_49 ) );
  DFF_X1 key_b_r_reg_7_5 (.CK( clk ) , .D( key_b_r_6_5 ) , .Q( key_b_r_7_5 ) );
  DFF_X1 key_b_r_reg_7_50 (.CK( clk ) , .D( key_b_r_6_50 ) , .Q( key_b_r_7_50 ) );
  DFF_X1 key_b_r_reg_7_51 (.CK( clk ) , .D( key_b_r_6_51 ) , .Q( key_b_r_7_51 ) );
  DFF_X1 key_b_r_reg_7_52 (.CK( clk ) , .D( key_b_r_6_52 ) , .Q( key_b_r_7_52 ) );
  DFF_X1 key_b_r_reg_7_53 (.CK( clk ) , .D( key_b_r_6_53 ) , .Q( key_b_r_7_53 ) );
  DFF_X1 key_b_r_reg_7_54 (.CK( clk ) , .D( key_b_r_6_54 ) , .Q( key_b_r_7_54 ) );
  DFF_X1 key_b_r_reg_7_55 (.CK( clk ) , .D( key_b_r_6_55 ) , .Q( key_b_r_7_55 ) );
  DFF_X1 key_b_r_reg_7_6 (.CK( clk ) , .D( key_b_r_6_6 ) , .Q( key_b_r_7_6 ) );
  DFF_X1 key_b_r_reg_7_7 (.CK( clk ) , .D( key_b_r_6_7 ) , .Q( key_b_r_7_7 ) );
  DFF_X1 key_b_r_reg_7_8 (.CK( clk ) , .D( key_b_r_6_8 ) , .Q( key_b_r_7_8 ) );
  DFF_X1 key_b_r_reg_7_9 (.CK( clk ) , .D( key_b_r_6_9 ) , .Q( key_b_r_7_9 ) );
  DFF_X1 key_b_r_reg_8_0 (.CK( clk ) , .D( key_b_r_7_0 ) , .Q( key_b_r_8_0 ) );
  DFF_X1 key_b_r_reg_8_1 (.CK( clk ) , .D( key_b_r_7_1 ) , .Q( key_b_r_8_1 ) );
  DFF_X1 key_b_r_reg_8_10 (.CK( clk ) , .D( key_b_r_7_10 ) , .Q( key_b_r_8_10 ) );
  DFF_X1 key_b_r_reg_8_11 (.CK( clk ) , .D( key_b_r_7_11 ) , .Q( key_b_r_8_11 ) );
  DFF_X1 key_b_r_reg_8_12 (.CK( clk ) , .D( key_b_r_7_12 ) , .Q( key_b_r_8_12 ) );
  DFF_X1 key_b_r_reg_8_13 (.CK( clk ) , .D( key_b_r_7_13 ) , .Q( key_b_r_8_13 ) );
  DFF_X1 key_b_r_reg_8_14 (.CK( clk ) , .D( key_b_r_7_14 ) , .Q( key_b_r_8_14 ) );
  DFF_X1 key_b_r_reg_8_15 (.CK( clk ) , .D( key_b_r_7_15 ) , .Q( key_b_r_8_15 ) );
  DFF_X1 key_b_r_reg_8_16 (.CK( clk ) , .D( key_b_r_7_16 ) , .Q( key_b_r_8_16 ) );
  DFF_X1 key_b_r_reg_8_17 (.CK( clk ) , .D( key_b_r_7_17 ) , .Q( key_b_r_8_17 ) );
  DFF_X1 key_b_r_reg_8_18 (.CK( clk ) , .D( key_b_r_7_18 ) , .Q( key_b_r_8_18 ) );
  DFF_X1 key_b_r_reg_8_19 (.CK( clk ) , .D( key_b_r_7_19 ) , .Q( key_b_r_8_19 ) );
  DFF_X1 key_b_r_reg_8_2 (.CK( clk ) , .D( key_b_r_7_2 ) , .Q( key_b_r_8_2 ) );
  DFF_X1 key_b_r_reg_8_20 (.CK( clk ) , .D( key_b_r_7_20 ) , .Q( key_b_r_8_20 ) );
  DFF_X1 key_b_r_reg_8_21 (.CK( clk ) , .D( key_b_r_7_21 ) , .Q( key_b_r_8_21 ) );
  DFF_X1 key_b_r_reg_8_22 (.CK( clk ) , .D( key_b_r_7_22 ) , .Q( key_b_r_8_22 ) );
  DFF_X1 key_b_r_reg_8_23 (.CK( clk ) , .D( key_b_r_7_23 ) , .Q( key_b_r_8_23 ) );
  DFF_X1 key_b_r_reg_8_24 (.CK( clk ) , .D( key_b_r_7_24 ) , .Q( key_b_r_8_24 ) );
  DFF_X1 key_b_r_reg_8_25 (.CK( clk ) , .D( key_b_r_7_25 ) , .Q( key_b_r_8_25 ) );
  DFF_X1 key_b_r_reg_8_26 (.CK( clk ) , .D( key_b_r_7_26 ) , .Q( key_b_r_8_26 ) );
  DFF_X1 key_b_r_reg_8_27 (.CK( clk ) , .D( key_b_r_7_27 ) , .Q( key_b_r_8_27 ) );
  DFF_X1 key_b_r_reg_8_28 (.CK( clk ) , .D( key_b_r_7_28 ) , .Q( key_b_r_8_28 ) );
  DFF_X1 key_b_r_reg_8_29 (.CK( clk ) , .D( key_b_r_7_29 ) , .Q( key_b_r_8_29 ) );
  DFF_X1 key_b_r_reg_8_3 (.CK( clk ) , .D( key_b_r_7_3 ) , .Q( key_b_r_8_3 ) );
  DFF_X1 key_b_r_reg_8_30 (.CK( clk ) , .D( key_b_r_7_30 ) , .Q( key_b_r_8_30 ) );
  DFF_X1 key_b_r_reg_8_31 (.CK( clk ) , .D( key_b_r_7_31 ) , .Q( key_b_r_8_31 ) );
  DFF_X1 key_b_r_reg_8_32 (.CK( clk ) , .D( key_b_r_7_32 ) , .Q( key_b_r_8_32 ) );
  DFF_X1 key_b_r_reg_8_33 (.CK( clk ) , .D( key_b_r_7_33 ) , .Q( key_b_r_8_33 ) );
  DFF_X1 key_b_r_reg_8_34 (.CK( clk ) , .D( key_b_r_7_34 ) , .Q( key_b_r_8_34 ) );
  DFF_X1 key_b_r_reg_8_35 (.CK( clk ) , .D( key_b_r_7_35 ) , .Q( key_b_r_8_35 ) );
  DFF_X1 key_b_r_reg_8_36 (.CK( clk ) , .D( key_b_r_7_36 ) , .Q( key_b_r_8_36 ) );
  DFF_X1 key_b_r_reg_8_37 (.CK( clk ) , .D( key_b_r_7_37 ) , .Q( key_b_r_8_37 ) );
  DFF_X1 key_b_r_reg_8_38 (.CK( clk ) , .D( key_b_r_7_38 ) , .Q( key_b_r_8_38 ) );
  DFF_X1 key_b_r_reg_8_39 (.CK( clk ) , .D( key_b_r_7_39 ) , .Q( key_b_r_8_39 ) );
  DFF_X1 key_b_r_reg_8_4 (.CK( clk ) , .D( key_b_r_7_4 ) , .Q( key_b_r_8_4 ) );
  DFF_X1 key_b_r_reg_8_40 (.CK( clk ) , .D( key_b_r_7_40 ) , .Q( key_b_r_8_40 ) );
  DFF_X1 key_b_r_reg_8_41 (.CK( clk ) , .D( key_b_r_7_41 ) , .Q( key_b_r_8_41 ) );
  DFF_X1 key_b_r_reg_8_42 (.CK( clk ) , .D( key_b_r_7_42 ) , .Q( key_b_r_8_42 ) );
  DFF_X1 key_b_r_reg_8_43 (.CK( clk ) , .D( key_b_r_7_43 ) , .Q( key_b_r_8_43 ) );
  DFF_X1 key_b_r_reg_8_44 (.CK( clk ) , .D( key_b_r_7_44 ) , .Q( key_b_r_8_44 ) );
  DFF_X1 key_b_r_reg_8_45 (.CK( clk ) , .D( key_b_r_7_45 ) , .Q( key_b_r_8_45 ) );
  DFF_X1 key_b_r_reg_8_46 (.CK( clk ) , .D( key_b_r_7_46 ) , .Q( key_b_r_8_46 ) );
  DFF_X1 key_b_r_reg_8_47 (.CK( clk ) , .D( key_b_r_7_47 ) , .Q( key_b_r_8_47 ) );
  DFF_X1 key_b_r_reg_8_48 (.CK( clk ) , .D( key_b_r_7_48 ) , .Q( key_b_r_8_48 ) );
  DFF_X1 key_b_r_reg_8_49 (.CK( clk ) , .D( key_b_r_7_49 ) , .Q( key_b_r_8_49 ) );
  DFF_X1 key_b_r_reg_8_5 (.CK( clk ) , .D( key_b_r_7_5 ) , .Q( key_b_r_8_5 ) );
  DFF_X1 key_b_r_reg_8_50 (.CK( clk ) , .D( key_b_r_7_50 ) , .Q( key_b_r_8_50 ) );
  DFF_X1 key_b_r_reg_8_51 (.CK( clk ) , .D( key_b_r_7_51 ) , .Q( key_b_r_8_51 ) );
  DFF_X1 key_b_r_reg_8_52 (.CK( clk ) , .D( key_b_r_7_52 ) , .Q( key_b_r_8_52 ) );
  DFF_X1 key_b_r_reg_8_53 (.CK( clk ) , .D( key_b_r_7_53 ) , .Q( key_b_r_8_53 ) );
  DFF_X1 key_b_r_reg_8_54 (.CK( clk ) , .D( key_b_r_7_54 ) , .Q( key_b_r_8_54 ) );
  DFF_X1 key_b_r_reg_8_55 (.CK( clk ) , .D( key_b_r_7_55 ) , .Q( key_b_r_8_55 ) );
  DFF_X1 key_b_r_reg_8_6 (.CK( clk ) , .D( key_b_r_7_6 ) , .Q( key_b_r_8_6 ) );
  DFF_X1 key_b_r_reg_8_7 (.CK( clk ) , .D( key_b_r_7_7 ) , .Q( key_b_r_8_7 ) );
  DFF_X1 key_b_r_reg_8_8 (.CK( clk ) , .D( key_b_r_7_8 ) , .Q( key_b_r_8_8 ) );
  DFF_X1 key_b_r_reg_8_9 (.CK( clk ) , .D( key_b_r_7_9 ) , .Q( key_b_r_8_9 ) );
  DFF_X1 key_b_r_reg_9_0 (.CK( clk ) , .D( key_b_r_8_0 ) , .Q( key_b_r_9_0 ) );
  DFF_X1 key_b_r_reg_9_1 (.CK( clk ) , .D( key_b_r_8_1 ) , .Q( key_b_r_9_1 ) );
  DFF_X1 key_b_r_reg_9_10 (.CK( clk ) , .D( key_b_r_8_10 ) , .Q( key_b_r_9_10 ) );
  DFF_X1 key_b_r_reg_9_11 (.CK( clk ) , .D( key_b_r_8_11 ) , .Q( key_b_r_9_11 ) );
  DFF_X1 key_b_r_reg_9_12 (.CK( clk ) , .D( key_b_r_8_12 ) , .Q( key_b_r_9_12 ) );
  DFF_X1 key_b_r_reg_9_13 (.CK( clk ) , .D( key_b_r_8_13 ) , .Q( key_b_r_9_13 ) );
  DFF_X1 key_b_r_reg_9_14 (.CK( clk ) , .D( key_b_r_8_14 ) , .Q( key_b_r_9_14 ) );
  DFF_X1 key_b_r_reg_9_15 (.CK( clk ) , .D( key_b_r_8_15 ) , .Q( key_b_r_9_15 ) );
  DFF_X1 key_b_r_reg_9_16 (.CK( clk ) , .D( key_b_r_8_16 ) , .Q( key_b_r_9_16 ) );
  DFF_X1 key_b_r_reg_9_17 (.CK( clk ) , .D( key_b_r_8_17 ) , .Q( key_b_r_9_17 ) );
  DFF_X1 key_b_r_reg_9_18 (.CK( clk ) , .D( key_b_r_8_18 ) , .Q( key_b_r_9_18 ) );
  DFF_X1 key_b_r_reg_9_19 (.CK( clk ) , .D( key_b_r_8_19 ) , .Q( key_b_r_9_19 ) );
  DFF_X1 key_b_r_reg_9_2 (.CK( clk ) , .D( key_b_r_8_2 ) , .Q( key_b_r_9_2 ) );
  DFF_X1 key_b_r_reg_9_20 (.CK( clk ) , .D( key_b_r_8_20 ) , .Q( key_b_r_9_20 ) );
  DFF_X1 key_b_r_reg_9_21 (.CK( clk ) , .D( key_b_r_8_21 ) , .Q( key_b_r_9_21 ) );
  DFF_X1 key_b_r_reg_9_22 (.CK( clk ) , .D( key_b_r_8_22 ) , .Q( key_b_r_9_22 ) );
  DFF_X1 key_b_r_reg_9_23 (.CK( clk ) , .D( key_b_r_8_23 ) , .Q( key_b_r_9_23 ) );
  DFF_X1 key_b_r_reg_9_24 (.CK( clk ) , .D( key_b_r_8_24 ) , .Q( key_b_r_9_24 ) );
  DFF_X1 key_b_r_reg_9_25 (.CK( clk ) , .D( key_b_r_8_25 ) , .Q( key_b_r_9_25 ) );
  DFF_X1 key_b_r_reg_9_26 (.CK( clk ) , .D( key_b_r_8_26 ) , .Q( key_b_r_9_26 ) );
  DFF_X1 key_b_r_reg_9_27 (.CK( clk ) , .D( key_b_r_8_27 ) , .Q( key_b_r_9_27 ) );
  DFF_X1 key_b_r_reg_9_28 (.CK( clk ) , .D( key_b_r_8_28 ) , .Q( key_b_r_9_28 ) );
  DFF_X1 key_b_r_reg_9_29 (.CK( clk ) , .D( key_b_r_8_29 ) , .Q( key_b_r_9_29 ) );
  DFF_X1 key_b_r_reg_9_3 (.CK( clk ) , .D( key_b_r_8_3 ) , .Q( key_b_r_9_3 ) );
  DFF_X1 key_b_r_reg_9_30 (.CK( clk ) , .D( key_b_r_8_30 ) , .Q( key_b_r_9_30 ) );
  DFF_X1 key_b_r_reg_9_31 (.CK( clk ) , .D( key_b_r_8_31 ) , .Q( key_b_r_9_31 ) );
  DFF_X1 key_b_r_reg_9_32 (.CK( clk ) , .D( key_b_r_8_32 ) , .Q( key_b_r_9_32 ) );
  DFF_X1 key_b_r_reg_9_33 (.CK( clk ) , .D( key_b_r_8_33 ) , .Q( key_b_r_9_33 ) );
  DFF_X1 key_b_r_reg_9_34 (.CK( clk ) , .D( key_b_r_8_34 ) , .Q( key_b_r_9_34 ) );
  DFF_X1 key_b_r_reg_9_35 (.CK( clk ) , .D( key_b_r_8_35 ) , .Q( key_b_r_9_35 ) );
  DFF_X1 key_b_r_reg_9_36 (.CK( clk ) , .D( key_b_r_8_36 ) , .Q( key_b_r_9_36 ) );
  DFF_X1 key_b_r_reg_9_37 (.CK( clk ) , .D( key_b_r_8_37 ) , .Q( key_b_r_9_37 ) );
  DFF_X1 key_b_r_reg_9_38 (.CK( clk ) , .D( key_b_r_8_38 ) , .Q( key_b_r_9_38 ) );
  DFF_X1 key_b_r_reg_9_39 (.CK( clk ) , .D( key_b_r_8_39 ) , .Q( key_b_r_9_39 ) );
  DFF_X1 key_b_r_reg_9_4 (.CK( clk ) , .D( key_b_r_8_4 ) , .Q( key_b_r_9_4 ) );
  DFF_X1 key_b_r_reg_9_40 (.CK( clk ) , .D( key_b_r_8_40 ) , .Q( key_b_r_9_40 ) );
  DFF_X1 key_b_r_reg_9_41 (.CK( clk ) , .D( key_b_r_8_41 ) , .Q( key_b_r_9_41 ) );
  DFF_X1 key_b_r_reg_9_42 (.CK( clk ) , .D( key_b_r_8_42 ) , .Q( key_b_r_9_42 ) );
  DFF_X1 key_b_r_reg_9_43 (.CK( clk ) , .D( key_b_r_8_43 ) , .Q( key_b_r_9_43 ) );
  DFF_X1 key_b_r_reg_9_44 (.CK( clk ) , .D( key_b_r_8_44 ) , .Q( key_b_r_9_44 ) );
  DFF_X1 key_b_r_reg_9_45 (.CK( clk ) , .D( key_b_r_8_45 ) , .Q( key_b_r_9_45 ) );
  DFF_X1 key_b_r_reg_9_46 (.CK( clk ) , .D( key_b_r_8_46 ) , .Q( key_b_r_9_46 ) );
  DFF_X1 key_b_r_reg_9_47 (.CK( clk ) , .D( key_b_r_8_47 ) , .Q( key_b_r_9_47 ) );
  DFF_X1 key_b_r_reg_9_48 (.CK( clk ) , .D( key_b_r_8_48 ) , .Q( key_b_r_9_48 ) );
  DFF_X1 key_b_r_reg_9_49 (.CK( clk ) , .D( key_b_r_8_49 ) , .Q( key_b_r_9_49 ) );
  DFF_X1 key_b_r_reg_9_5 (.CK( clk ) , .D( key_b_r_8_5 ) , .Q( key_b_r_9_5 ) );
  DFF_X1 key_b_r_reg_9_50 (.CK( clk ) , .D( key_b_r_8_50 ) , .Q( key_b_r_9_50 ) );
  DFF_X1 key_b_r_reg_9_51 (.CK( clk ) , .D( key_b_r_8_51 ) , .Q( key_b_r_9_51 ) );
  DFF_X1 key_b_r_reg_9_52 (.CK( clk ) , .D( key_b_r_8_52 ) , .Q( key_b_r_9_52 ) );
  DFF_X1 key_b_r_reg_9_53 (.CK( clk ) , .D( key_b_r_8_53 ) , .Q( key_b_r_9_53 ) );
  DFF_X1 key_b_r_reg_9_54 (.CK( clk ) , .D( key_b_r_8_54 ) , .Q( key_b_r_9_54 ) );
  DFF_X1 key_b_r_reg_9_55 (.CK( clk ) , .D( key_b_r_8_55 ) , .Q( key_b_r_9_55 ) );
  DFF_X1 key_b_r_reg_9_6 (.CK( clk ) , .D( key_b_r_8_6 ) , .Q( key_b_r_9_6 ) );
  DFF_X1 key_b_r_reg_9_7 (.CK( clk ) , .D( key_b_r_8_7 ) , .Q( key_b_r_9_7 ) );
  DFF_X1 key_b_r_reg_9_8 (.CK( clk ) , .D( key_b_r_8_8 ) , .Q( key_b_r_9_8 ) );
  DFF_X1 key_b_r_reg_9_9 (.CK( clk ) , .D( key_b_r_8_9 ) , .Q( key_b_r_9_9 ) );
  SDFF_X1 key_c_r_reg_0_0 (.CK( clk ) , .SE( decrypt ) , .SI( key1[0] ) , .D( key3[0] ) , .Q( key_c_r_0_0 ) );
  SDFF_X1 key_c_r_reg_0_1 (.CK( clk ) , .SE( decrypt ) , .SI( key1[1] ) , .D( key3[1] ) , .Q( key_c_r_0_1 ) );
  SDFF_X1 key_c_r_reg_0_10 (.CK( clk ) , .SE( decrypt ) , .SI( key1[10] ) , .D( key3[10] ) , .Q( key_c_r_0_10 ) );
  SDFF_X1 key_c_r_reg_0_11 (.CK( clk ) , .SE( decrypt ) , .SI( key1[11] ) , .D( key3[11] ) , .Q( key_c_r_0_11 ) );
  SDFF_X1 key_c_r_reg_0_12 (.CK( clk ) , .SE( decrypt ) , .SI( key1[12] ) , .D( key3[12] ) , .Q( key_c_r_0_12 ) );
  SDFF_X1 key_c_r_reg_0_13 (.CK( clk ) , .SE( decrypt ) , .SI( key1[13] ) , .D( key3[13] ) , .Q( key_c_r_0_13 ) );
  SDFF_X1 key_c_r_reg_0_14 (.CK( clk ) , .SE( decrypt ) , .SI( key1[14] ) , .D( key3[14] ) , .Q( key_c_r_0_14 ) );
  SDFF_X1 key_c_r_reg_0_15 (.CK( clk ) , .SE( decrypt ) , .SI( key1[15] ) , .D( key3[15] ) , .Q( key_c_r_0_15 ) );
  SDFF_X1 key_c_r_reg_0_16 (.CK( clk ) , .SE( decrypt ) , .SI( key1[16] ) , .D( key3[16] ) , .Q( key_c_r_0_16 ) );
  SDFF_X1 key_c_r_reg_0_17 (.CK( clk ) , .SE( decrypt ) , .SI( key1[17] ) , .D( key3[17] ) , .Q( key_c_r_0_17 ) );
  SDFF_X1 key_c_r_reg_0_18 (.CK( clk ) , .SE( decrypt ) , .SI( key1[18] ) , .D( key3[18] ) , .Q( key_c_r_0_18 ) );
  SDFF_X1 key_c_r_reg_0_19 (.CK( clk ) , .SE( decrypt ) , .SI( key1[19] ) , .D( key3[19] ) , .Q( key_c_r_0_19 ) );
  SDFF_X1 key_c_r_reg_0_2 (.CK( clk ) , .SE( decrypt ) , .SI( key1[2] ) , .D( key3[2] ) , .Q( key_c_r_0_2 ) );
  SDFF_X1 key_c_r_reg_0_20 (.CK( clk ) , .SE( decrypt ) , .SI( key1[20] ) , .D( key3[20] ) , .Q( key_c_r_0_20 ) );
  SDFF_X1 key_c_r_reg_0_21 (.CK( clk ) , .SE( decrypt ) , .SI( key1[21] ) , .D( key3[21] ) , .Q( key_c_r_0_21 ) );
  SDFF_X1 key_c_r_reg_0_22 (.CK( clk ) , .SE( decrypt ) , .SI( key1[22] ) , .D( key3[22] ) , .Q( key_c_r_0_22 ) );
  SDFF_X1 key_c_r_reg_0_23 (.CK( clk ) , .SE( decrypt ) , .SI( key1[23] ) , .D( key3[23] ) , .Q( key_c_r_0_23 ) );
  SDFF_X1 key_c_r_reg_0_24 (.CK( clk ) , .SE( decrypt ) , .SI( key1[24] ) , .D( key3[24] ) , .Q( key_c_r_0_24 ) );
  SDFF_X1 key_c_r_reg_0_25 (.CK( clk ) , .SE( decrypt ) , .SI( key1[25] ) , .D( key3[25] ) , .Q( key_c_r_0_25 ) );
  SDFF_X1 key_c_r_reg_0_26 (.CK( clk ) , .SE( decrypt ) , .SI( key1[26] ) , .D( key3[26] ) , .Q( key_c_r_0_26 ) );
  SDFF_X1 key_c_r_reg_0_27 (.CK( clk ) , .SE( decrypt ) , .SI( key1[27] ) , .D( key3[27] ) , .Q( key_c_r_0_27 ) );
  SDFF_X1 key_c_r_reg_0_28 (.CK( clk ) , .SE( decrypt ) , .SI( key1[28] ) , .D( key3[28] ) , .Q( key_c_r_0_28 ) );
  SDFF_X1 key_c_r_reg_0_29 (.CK( clk ) , .SE( decrypt ) , .SI( key1[29] ) , .D( key3[29] ) , .Q( key_c_r_0_29 ) );
  SDFF_X1 key_c_r_reg_0_3 (.CK( clk ) , .SE( decrypt ) , .SI( key1[3] ) , .D( key3[3] ) , .Q( key_c_r_0_3 ) );
  SDFF_X1 key_c_r_reg_0_30 (.CK( clk ) , .SE( decrypt ) , .SI( key1[30] ) , .D( key3[30] ) , .Q( key_c_r_0_30 ) );
  SDFF_X1 key_c_r_reg_0_31 (.CK( clk ) , .SE( decrypt ) , .SI( key1[31] ) , .D( key3[31] ) , .Q( key_c_r_0_31 ) );
  SDFF_X1 key_c_r_reg_0_32 (.CK( clk ) , .SE( decrypt ) , .SI( key1[32] ) , .D( key3[32] ) , .Q( key_c_r_0_32 ) );
  SDFF_X1 key_c_r_reg_0_33 (.CK( clk ) , .SE( decrypt ) , .SI( key1[33] ) , .D( key3[33] ) , .Q( key_c_r_0_33 ) );
  SDFF_X1 key_c_r_reg_0_34 (.CK( clk ) , .SE( decrypt ) , .SI( key1[34] ) , .D( key3[34] ) , .Q( key_c_r_0_34 ) );
  SDFF_X1 key_c_r_reg_0_35 (.CK( clk ) , .SE( decrypt ) , .SI( key1[35] ) , .D( key3[35] ) , .Q( key_c_r_0_35 ) );
  SDFF_X1 key_c_r_reg_0_36 (.CK( clk ) , .SE( decrypt ) , .SI( key1[36] ) , .D( key3[36] ) , .Q( key_c_r_0_36 ) );
  SDFF_X1 key_c_r_reg_0_37 (.CK( clk ) , .SE( decrypt ) , .SI( key1[37] ) , .D( key3[37] ) , .Q( key_c_r_0_37 ) );
  SDFF_X1 key_c_r_reg_0_38 (.CK( clk ) , .SE( decrypt ) , .SI( key1[38] ) , .D( key3[38] ) , .Q( key_c_r_0_38 ) );
  SDFF_X1 key_c_r_reg_0_39 (.CK( clk ) , .SE( decrypt ) , .SI( key1[39] ) , .D( key3[39] ) , .Q( key_c_r_0_39 ) );
  SDFF_X1 key_c_r_reg_0_4 (.CK( clk ) , .SE( decrypt ) , .SI( key1[4] ) , .D( key3[4] ) , .Q( key_c_r_0_4 ) );
  SDFF_X1 key_c_r_reg_0_40 (.CK( clk ) , .SE( decrypt ) , .SI( key1[40] ) , .D( key3[40] ) , .Q( key_c_r_0_40 ) );
  SDFF_X1 key_c_r_reg_0_41 (.CK( clk ) , .SE( decrypt ) , .SI( key1[41] ) , .D( key3[41] ) , .Q( key_c_r_0_41 ) );
  SDFF_X1 key_c_r_reg_0_42 (.CK( clk ) , .SE( decrypt ) , .SI( key1[42] ) , .D( key3[42] ) , .Q( key_c_r_0_42 ) );
  SDFF_X1 key_c_r_reg_0_43 (.CK( clk ) , .SE( decrypt ) , .SI( key1[43] ) , .D( key3[43] ) , .Q( key_c_r_0_43 ) );
  SDFF_X1 key_c_r_reg_0_44 (.CK( clk ) , .SE( decrypt ) , .SI( key1[44] ) , .D( key3[44] ) , .Q( key_c_r_0_44 ) );
  SDFF_X1 key_c_r_reg_0_45 (.CK( clk ) , .SE( decrypt ) , .SI( key1[45] ) , .D( key3[45] ) , .Q( key_c_r_0_45 ) );
  SDFF_X1 key_c_r_reg_0_46 (.CK( clk ) , .SE( decrypt ) , .SI( key1[46] ) , .D( key3[46] ) , .Q( key_c_r_0_46 ) );
  SDFF_X1 key_c_r_reg_0_47 (.CK( clk ) , .SE( decrypt ) , .SI( key1[47] ) , .D( key3[47] ) , .Q( key_c_r_0_47 ) );
  SDFF_X1 key_c_r_reg_0_48 (.CK( clk ) , .SE( decrypt ) , .SI( key1[48] ) , .D( key3[48] ) , .Q( key_c_r_0_48 ) );
  SDFF_X1 key_c_r_reg_0_49 (.CK( clk ) , .SE( decrypt ) , .SI( key1[49] ) , .D( key3[49] ) , .Q( key_c_r_0_49 ) );
  SDFF_X1 key_c_r_reg_0_5 (.CK( clk ) , .SE( decrypt ) , .SI( key1[5] ) , .D( key3[5] ) , .Q( key_c_r_0_5 ) );
  SDFF_X1 key_c_r_reg_0_50 (.CK( clk ) , .SE( decrypt ) , .SI( key1[50] ) , .D( key3[50] ) , .Q( key_c_r_0_50 ) );
  SDFF_X1 key_c_r_reg_0_51 (.CK( clk ) , .SE( decrypt ) , .SI( key1[51] ) , .D( key3[51] ) , .Q( key_c_r_0_51 ) );
  SDFF_X1 key_c_r_reg_0_52 (.CK( clk ) , .SE( decrypt ) , .SI( key1[52] ) , .D( key3[52] ) , .Q( key_c_r_0_52 ) );
  SDFF_X1 key_c_r_reg_0_53 (.CK( clk ) , .SE( decrypt ) , .SI( key1[53] ) , .D( key3[53] ) , .Q( key_c_r_0_53 ) );
  SDFF_X1 key_c_r_reg_0_54 (.CK( clk ) , .SE( decrypt ) , .SI( key1[54] ) , .D( key3[54] ) , .Q( key_c_r_0_54 ) );
  SDFF_X1 key_c_r_reg_0_55 (.CK( clk ) , .SE( decrypt ) , .SI( key1[55] ) , .D( key3[55] ) , .Q( key_c_r_0_55 ) );
  SDFF_X1 key_c_r_reg_0_6 (.CK( clk ) , .SE( decrypt ) , .SI( key1[6] ) , .D( key3[6] ) , .Q( key_c_r_0_6 ) );
  SDFF_X1 key_c_r_reg_0_7 (.CK( clk ) , .SE( decrypt ) , .SI( key1[7] ) , .D( key3[7] ) , .Q( key_c_r_0_7 ) );
  SDFF_X1 key_c_r_reg_0_8 (.CK( clk ) , .SE( decrypt ) , .SI( key1[8] ) , .D( key3[8] ) , .Q( key_c_r_0_8 ) );
  SDFF_X1 key_c_r_reg_0_9 (.CK( clk ) , .SE( decrypt ) , .SI( key1[9] ) , .D( key3[9] ) , .Q( key_c_r_0_9 ) );
  DFF_X1 key_c_r_reg_10_0 (.CK( clk ) , .Q( key_c_r_10_0 ) , .D( key_c_r_9_0 ) );
  DFF_X1 key_c_r_reg_10_1 (.CK( clk ) , .Q( key_c_r_10_1 ) , .D( key_c_r_9_1 ) );
  DFF_X1 key_c_r_reg_10_10 (.CK( clk ) , .Q( key_c_r_10_10 ) , .D( key_c_r_9_10 ) );
  DFF_X1 key_c_r_reg_10_11 (.CK( clk ) , .Q( key_c_r_10_11 ) , .D( key_c_r_9_11 ) );
  DFF_X1 key_c_r_reg_10_12 (.CK( clk ) , .Q( key_c_r_10_12 ) , .D( key_c_r_9_12 ) );
  DFF_X1 key_c_r_reg_10_13 (.CK( clk ) , .Q( key_c_r_10_13 ) , .D( key_c_r_9_13 ) );
  DFF_X1 key_c_r_reg_10_14 (.CK( clk ) , .Q( key_c_r_10_14 ) , .D( key_c_r_9_14 ) );
  DFF_X1 key_c_r_reg_10_15 (.CK( clk ) , .Q( key_c_r_10_15 ) , .D( key_c_r_9_15 ) );
  DFF_X1 key_c_r_reg_10_16 (.CK( clk ) , .Q( key_c_r_10_16 ) , .D( key_c_r_9_16 ) );
  DFF_X1 key_c_r_reg_10_17 (.CK( clk ) , .Q( key_c_r_10_17 ) , .D( key_c_r_9_17 ) );
  DFF_X1 key_c_r_reg_10_18 (.CK( clk ) , .Q( key_c_r_10_18 ) , .D( key_c_r_9_18 ) );
  DFF_X1 key_c_r_reg_10_19 (.CK( clk ) , .Q( key_c_r_10_19 ) , .D( key_c_r_9_19 ) );
  DFF_X1 key_c_r_reg_10_2 (.CK( clk ) , .Q( key_c_r_10_2 ) , .D( key_c_r_9_2 ) );
  DFF_X1 key_c_r_reg_10_20 (.CK( clk ) , .Q( key_c_r_10_20 ) , .D( key_c_r_9_20 ) );
  DFF_X1 key_c_r_reg_10_21 (.CK( clk ) , .Q( key_c_r_10_21 ) , .D( key_c_r_9_21 ) );
  DFF_X1 key_c_r_reg_10_22 (.CK( clk ) , .Q( key_c_r_10_22 ) , .D( key_c_r_9_22 ) );
  DFF_X1 key_c_r_reg_10_23 (.CK( clk ) , .Q( key_c_r_10_23 ) , .D( key_c_r_9_23 ) );
  DFF_X1 key_c_r_reg_10_24 (.CK( clk ) , .Q( key_c_r_10_24 ) , .D( key_c_r_9_24 ) );
  DFF_X1 key_c_r_reg_10_25 (.CK( clk ) , .Q( key_c_r_10_25 ) , .D( key_c_r_9_25 ) );
  DFF_X1 key_c_r_reg_10_26 (.CK( clk ) , .Q( key_c_r_10_26 ) , .D( key_c_r_9_26 ) );
  DFF_X1 key_c_r_reg_10_27 (.CK( clk ) , .Q( key_c_r_10_27 ) , .D( key_c_r_9_27 ) );
  DFF_X1 key_c_r_reg_10_28 (.CK( clk ) , .Q( key_c_r_10_28 ) , .D( key_c_r_9_28 ) );
  DFF_X1 key_c_r_reg_10_29 (.CK( clk ) , .Q( key_c_r_10_29 ) , .D( key_c_r_9_29 ) );
  DFF_X1 key_c_r_reg_10_3 (.CK( clk ) , .Q( key_c_r_10_3 ) , .D( key_c_r_9_3 ) );
  DFF_X1 key_c_r_reg_10_30 (.CK( clk ) , .Q( key_c_r_10_30 ) , .D( key_c_r_9_30 ) );
  DFF_X1 key_c_r_reg_10_31 (.CK( clk ) , .Q( key_c_r_10_31 ) , .D( key_c_r_9_31 ) );
  DFF_X1 key_c_r_reg_10_32 (.CK( clk ) , .Q( key_c_r_10_32 ) , .D( key_c_r_9_32 ) );
  DFF_X1 key_c_r_reg_10_33 (.CK( clk ) , .Q( key_c_r_10_33 ) , .D( key_c_r_9_33 ) );
  DFF_X1 key_c_r_reg_10_34 (.CK( clk ) , .Q( key_c_r_10_34 ) , .D( key_c_r_9_34 ) );
  DFF_X1 key_c_r_reg_10_35 (.CK( clk ) , .Q( key_c_r_10_35 ) , .D( key_c_r_9_35 ) );
  DFF_X1 key_c_r_reg_10_36 (.CK( clk ) , .Q( key_c_r_10_36 ) , .D( key_c_r_9_36 ) );
  DFF_X1 key_c_r_reg_10_37 (.CK( clk ) , .Q( key_c_r_10_37 ) , .D( key_c_r_9_37 ) );
  DFF_X1 key_c_r_reg_10_38 (.CK( clk ) , .Q( key_c_r_10_38 ) , .D( key_c_r_9_38 ) );
  DFF_X1 key_c_r_reg_10_39 (.CK( clk ) , .Q( key_c_r_10_39 ) , .D( key_c_r_9_39 ) );
  DFF_X1 key_c_r_reg_10_4 (.CK( clk ) , .Q( key_c_r_10_4 ) , .D( key_c_r_9_4 ) );
  DFF_X1 key_c_r_reg_10_40 (.CK( clk ) , .Q( key_c_r_10_40 ) , .D( key_c_r_9_40 ) );
  DFF_X1 key_c_r_reg_10_41 (.CK( clk ) , .Q( key_c_r_10_41 ) , .D( key_c_r_9_41 ) );
  DFF_X1 key_c_r_reg_10_42 (.CK( clk ) , .Q( key_c_r_10_42 ) , .D( key_c_r_9_42 ) );
  DFF_X1 key_c_r_reg_10_43 (.CK( clk ) , .Q( key_c_r_10_43 ) , .D( key_c_r_9_43 ) );
  DFF_X1 key_c_r_reg_10_44 (.CK( clk ) , .Q( key_c_r_10_44 ) , .D( key_c_r_9_44 ) );
  DFF_X1 key_c_r_reg_10_45 (.CK( clk ) , .Q( key_c_r_10_45 ) , .D( key_c_r_9_45 ) );
  DFF_X1 key_c_r_reg_10_46 (.CK( clk ) , .Q( key_c_r_10_46 ) , .D( key_c_r_9_46 ) );
  DFF_X1 key_c_r_reg_10_47 (.CK( clk ) , .Q( key_c_r_10_47 ) , .D( key_c_r_9_47 ) );
  DFF_X1 key_c_r_reg_10_48 (.CK( clk ) , .Q( key_c_r_10_48 ) , .D( key_c_r_9_48 ) );
  DFF_X1 key_c_r_reg_10_49 (.CK( clk ) , .Q( key_c_r_10_49 ) , .D( key_c_r_9_49 ) );
  DFF_X1 key_c_r_reg_10_5 (.CK( clk ) , .Q( key_c_r_10_5 ) , .D( key_c_r_9_5 ) );
  DFF_X1 key_c_r_reg_10_50 (.CK( clk ) , .Q( key_c_r_10_50 ) , .D( key_c_r_9_50 ) );
  DFF_X1 key_c_r_reg_10_51 (.CK( clk ) , .Q( key_c_r_10_51 ) , .D( key_c_r_9_51 ) );
  DFF_X1 key_c_r_reg_10_52 (.CK( clk ) , .Q( key_c_r_10_52 ) , .D( key_c_r_9_52 ) );
  DFF_X1 key_c_r_reg_10_53 (.CK( clk ) , .Q( key_c_r_10_53 ) , .D( key_c_r_9_53 ) );
  DFF_X1 key_c_r_reg_10_54 (.CK( clk ) , .Q( key_c_r_10_54 ) , .D( key_c_r_9_54 ) );
  DFF_X1 key_c_r_reg_10_55 (.CK( clk ) , .Q( key_c_r_10_55 ) , .D( key_c_r_9_55 ) );
  DFF_X1 key_c_r_reg_10_6 (.CK( clk ) , .Q( key_c_r_10_6 ) , .D( key_c_r_9_6 ) );
  DFF_X1 key_c_r_reg_10_7 (.CK( clk ) , .Q( key_c_r_10_7 ) , .D( key_c_r_9_7 ) );
  DFF_X1 key_c_r_reg_10_8 (.CK( clk ) , .Q( key_c_r_10_8 ) , .D( key_c_r_9_8 ) );
  DFF_X1 key_c_r_reg_10_9 (.CK( clk ) , .Q( key_c_r_10_9 ) , .D( key_c_r_9_9 ) );
  DFF_X1 key_c_r_reg_11_0 (.CK( clk ) , .D( key_c_r_10_0 ) , .Q( key_c_r_11_0 ) );
  DFF_X1 key_c_r_reg_11_1 (.CK( clk ) , .D( key_c_r_10_1 ) , .Q( key_c_r_11_1 ) );
  DFF_X1 key_c_r_reg_11_10 (.CK( clk ) , .D( key_c_r_10_10 ) , .Q( key_c_r_11_10 ) );
  DFF_X1 key_c_r_reg_11_11 (.CK( clk ) , .D( key_c_r_10_11 ) , .Q( key_c_r_11_11 ) );
  DFF_X1 key_c_r_reg_11_12 (.CK( clk ) , .D( key_c_r_10_12 ) , .Q( key_c_r_11_12 ) );
  DFF_X1 key_c_r_reg_11_13 (.CK( clk ) , .D( key_c_r_10_13 ) , .Q( key_c_r_11_13 ) );
  DFF_X1 key_c_r_reg_11_14 (.CK( clk ) , .D( key_c_r_10_14 ) , .Q( key_c_r_11_14 ) );
  DFF_X1 key_c_r_reg_11_15 (.CK( clk ) , .D( key_c_r_10_15 ) , .Q( key_c_r_11_15 ) );
  DFF_X1 key_c_r_reg_11_16 (.CK( clk ) , .D( key_c_r_10_16 ) , .Q( key_c_r_11_16 ) );
  DFF_X1 key_c_r_reg_11_17 (.CK( clk ) , .D( key_c_r_10_17 ) , .Q( key_c_r_11_17 ) );
  DFF_X1 key_c_r_reg_11_18 (.CK( clk ) , .D( key_c_r_10_18 ) , .Q( key_c_r_11_18 ) );
  DFF_X1 key_c_r_reg_11_19 (.CK( clk ) , .D( key_c_r_10_19 ) , .Q( key_c_r_11_19 ) );
  DFF_X1 key_c_r_reg_11_2 (.CK( clk ) , .D( key_c_r_10_2 ) , .Q( key_c_r_11_2 ) );
  DFF_X1 key_c_r_reg_11_20 (.CK( clk ) , .D( key_c_r_10_20 ) , .Q( key_c_r_11_20 ) );
  DFF_X1 key_c_r_reg_11_21 (.CK( clk ) , .D( key_c_r_10_21 ) , .Q( key_c_r_11_21 ) );
  DFF_X1 key_c_r_reg_11_22 (.CK( clk ) , .D( key_c_r_10_22 ) , .Q( key_c_r_11_22 ) );
  DFF_X1 key_c_r_reg_11_23 (.CK( clk ) , .D( key_c_r_10_23 ) , .Q( key_c_r_11_23 ) );
  DFF_X1 key_c_r_reg_11_24 (.CK( clk ) , .D( key_c_r_10_24 ) , .Q( key_c_r_11_24 ) );
  DFF_X1 key_c_r_reg_11_25 (.CK( clk ) , .D( key_c_r_10_25 ) , .Q( key_c_r_11_25 ) );
  DFF_X1 key_c_r_reg_11_26 (.CK( clk ) , .D( key_c_r_10_26 ) , .Q( key_c_r_11_26 ) );
  DFF_X1 key_c_r_reg_11_27 (.CK( clk ) , .D( key_c_r_10_27 ) , .Q( key_c_r_11_27 ) );
  DFF_X1 key_c_r_reg_11_28 (.CK( clk ) , .D( key_c_r_10_28 ) , .Q( key_c_r_11_28 ) );
  DFF_X1 key_c_r_reg_11_29 (.CK( clk ) , .D( key_c_r_10_29 ) , .Q( key_c_r_11_29 ) );
  DFF_X1 key_c_r_reg_11_3 (.CK( clk ) , .D( key_c_r_10_3 ) , .Q( key_c_r_11_3 ) );
  DFF_X1 key_c_r_reg_11_30 (.CK( clk ) , .D( key_c_r_10_30 ) , .Q( key_c_r_11_30 ) );
  DFF_X1 key_c_r_reg_11_31 (.CK( clk ) , .D( key_c_r_10_31 ) , .Q( key_c_r_11_31 ) );
  DFF_X1 key_c_r_reg_11_32 (.CK( clk ) , .D( key_c_r_10_32 ) , .Q( key_c_r_11_32 ) );
  DFF_X1 key_c_r_reg_11_33 (.CK( clk ) , .D( key_c_r_10_33 ) , .Q( key_c_r_11_33 ) );
  DFF_X1 key_c_r_reg_11_34 (.CK( clk ) , .D( key_c_r_10_34 ) , .Q( key_c_r_11_34 ) );
  DFF_X1 key_c_r_reg_11_35 (.CK( clk ) , .D( key_c_r_10_35 ) , .Q( key_c_r_11_35 ) );
  DFF_X1 key_c_r_reg_11_36 (.CK( clk ) , .D( key_c_r_10_36 ) , .Q( key_c_r_11_36 ) );
  DFF_X1 key_c_r_reg_11_37 (.CK( clk ) , .D( key_c_r_10_37 ) , .Q( key_c_r_11_37 ) );
  DFF_X1 key_c_r_reg_11_38 (.CK( clk ) , .D( key_c_r_10_38 ) , .Q( key_c_r_11_38 ) );
  DFF_X1 key_c_r_reg_11_39 (.CK( clk ) , .D( key_c_r_10_39 ) , .Q( key_c_r_11_39 ) );
  DFF_X1 key_c_r_reg_11_4 (.CK( clk ) , .D( key_c_r_10_4 ) , .Q( key_c_r_11_4 ) );
  DFF_X1 key_c_r_reg_11_40 (.CK( clk ) , .D( key_c_r_10_40 ) , .Q( key_c_r_11_40 ) );
  DFF_X1 key_c_r_reg_11_41 (.CK( clk ) , .D( key_c_r_10_41 ) , .Q( key_c_r_11_41 ) );
  DFF_X1 key_c_r_reg_11_42 (.CK( clk ) , .D( key_c_r_10_42 ) , .Q( key_c_r_11_42 ) );
  DFF_X1 key_c_r_reg_11_43 (.CK( clk ) , .D( key_c_r_10_43 ) , .Q( key_c_r_11_43 ) );
  DFF_X1 key_c_r_reg_11_44 (.CK( clk ) , .D( key_c_r_10_44 ) , .Q( key_c_r_11_44 ) );
  DFF_X1 key_c_r_reg_11_45 (.CK( clk ) , .D( key_c_r_10_45 ) , .Q( key_c_r_11_45 ) );
  DFF_X1 key_c_r_reg_11_46 (.CK( clk ) , .D( key_c_r_10_46 ) , .Q( key_c_r_11_46 ) );
  DFF_X1 key_c_r_reg_11_47 (.CK( clk ) , .D( key_c_r_10_47 ) , .Q( key_c_r_11_47 ) );
  DFF_X1 key_c_r_reg_11_48 (.CK( clk ) , .D( key_c_r_10_48 ) , .Q( key_c_r_11_48 ) );
  DFF_X1 key_c_r_reg_11_49 (.CK( clk ) , .D( key_c_r_10_49 ) , .Q( key_c_r_11_49 ) );
  DFF_X1 key_c_r_reg_11_5 (.CK( clk ) , .D( key_c_r_10_5 ) , .Q( key_c_r_11_5 ) );
  DFF_X1 key_c_r_reg_11_50 (.CK( clk ) , .D( key_c_r_10_50 ) , .Q( key_c_r_11_50 ) );
  DFF_X1 key_c_r_reg_11_51 (.CK( clk ) , .D( key_c_r_10_51 ) , .Q( key_c_r_11_51 ) );
  DFF_X1 key_c_r_reg_11_52 (.CK( clk ) , .D( key_c_r_10_52 ) , .Q( key_c_r_11_52 ) );
  DFF_X1 key_c_r_reg_11_53 (.CK( clk ) , .D( key_c_r_10_53 ) , .Q( key_c_r_11_53 ) );
  DFF_X1 key_c_r_reg_11_54 (.CK( clk ) , .D( key_c_r_10_54 ) , .Q( key_c_r_11_54 ) );
  DFF_X1 key_c_r_reg_11_55 (.CK( clk ) , .D( key_c_r_10_55 ) , .Q( key_c_r_11_55 ) );
  DFF_X1 key_c_r_reg_11_6 (.CK( clk ) , .D( key_c_r_10_6 ) , .Q( key_c_r_11_6 ) );
  DFF_X1 key_c_r_reg_11_7 (.CK( clk ) , .D( key_c_r_10_7 ) , .Q( key_c_r_11_7 ) );
  DFF_X1 key_c_r_reg_11_8 (.CK( clk ) , .D( key_c_r_10_8 ) , .Q( key_c_r_11_8 ) );
  DFF_X1 key_c_r_reg_11_9 (.CK( clk ) , .D( key_c_r_10_9 ) , .Q( key_c_r_11_9 ) );
  DFF_X1 key_c_r_reg_12_0 (.CK( clk ) , .D( key_c_r_11_0 ) , .Q( key_c_r_12_0 ) );
  DFF_X1 key_c_r_reg_12_1 (.CK( clk ) , .D( key_c_r_11_1 ) , .Q( key_c_r_12_1 ) );
  DFF_X1 key_c_r_reg_12_10 (.CK( clk ) , .D( key_c_r_11_10 ) , .Q( key_c_r_12_10 ) );
  DFF_X1 key_c_r_reg_12_11 (.CK( clk ) , .D( key_c_r_11_11 ) , .Q( key_c_r_12_11 ) );
  DFF_X1 key_c_r_reg_12_12 (.CK( clk ) , .D( key_c_r_11_12 ) , .Q( key_c_r_12_12 ) );
  DFF_X1 key_c_r_reg_12_13 (.CK( clk ) , .D( key_c_r_11_13 ) , .Q( key_c_r_12_13 ) );
  DFF_X1 key_c_r_reg_12_14 (.CK( clk ) , .D( key_c_r_11_14 ) , .Q( key_c_r_12_14 ) );
  DFF_X1 key_c_r_reg_12_15 (.CK( clk ) , .D( key_c_r_11_15 ) , .Q( key_c_r_12_15 ) );
  DFF_X1 key_c_r_reg_12_16 (.CK( clk ) , .D( key_c_r_11_16 ) , .Q( key_c_r_12_16 ) );
  DFF_X1 key_c_r_reg_12_17 (.CK( clk ) , .D( key_c_r_11_17 ) , .Q( key_c_r_12_17 ) );
  DFF_X1 key_c_r_reg_12_18 (.CK( clk ) , .D( key_c_r_11_18 ) , .Q( key_c_r_12_18 ) );
  DFF_X1 key_c_r_reg_12_19 (.CK( clk ) , .D( key_c_r_11_19 ) , .Q( key_c_r_12_19 ) );
  DFF_X1 key_c_r_reg_12_2 (.CK( clk ) , .D( key_c_r_11_2 ) , .Q( key_c_r_12_2 ) );
  DFF_X1 key_c_r_reg_12_20 (.CK( clk ) , .D( key_c_r_11_20 ) , .Q( key_c_r_12_20 ) );
  DFF_X1 key_c_r_reg_12_21 (.CK( clk ) , .D( key_c_r_11_21 ) , .Q( key_c_r_12_21 ) );
  DFF_X1 key_c_r_reg_12_22 (.CK( clk ) , .D( key_c_r_11_22 ) , .Q( key_c_r_12_22 ) );
  DFF_X1 key_c_r_reg_12_23 (.CK( clk ) , .D( key_c_r_11_23 ) , .Q( key_c_r_12_23 ) );
  DFF_X1 key_c_r_reg_12_24 (.CK( clk ) , .D( key_c_r_11_24 ) , .Q( key_c_r_12_24 ) );
  DFF_X1 key_c_r_reg_12_25 (.CK( clk ) , .D( key_c_r_11_25 ) , .Q( key_c_r_12_25 ) );
  DFF_X1 key_c_r_reg_12_26 (.CK( clk ) , .D( key_c_r_11_26 ) , .Q( key_c_r_12_26 ) );
  DFF_X1 key_c_r_reg_12_27 (.CK( clk ) , .D( key_c_r_11_27 ) , .Q( key_c_r_12_27 ) );
  DFF_X1 key_c_r_reg_12_28 (.CK( clk ) , .D( key_c_r_11_28 ) , .Q( key_c_r_12_28 ) );
  DFF_X1 key_c_r_reg_12_29 (.CK( clk ) , .D( key_c_r_11_29 ) , .Q( key_c_r_12_29 ) );
  DFF_X1 key_c_r_reg_12_3 (.CK( clk ) , .D( key_c_r_11_3 ) , .Q( key_c_r_12_3 ) );
  DFF_X1 key_c_r_reg_12_30 (.CK( clk ) , .D( key_c_r_11_30 ) , .Q( key_c_r_12_30 ) );
  DFF_X1 key_c_r_reg_12_31 (.CK( clk ) , .D( key_c_r_11_31 ) , .Q( key_c_r_12_31 ) );
  DFF_X1 key_c_r_reg_12_32 (.CK( clk ) , .D( key_c_r_11_32 ) , .Q( key_c_r_12_32 ) );
  DFF_X1 key_c_r_reg_12_33 (.CK( clk ) , .D( key_c_r_11_33 ) , .Q( key_c_r_12_33 ) );
  DFF_X1 key_c_r_reg_12_34 (.CK( clk ) , .D( key_c_r_11_34 ) , .Q( key_c_r_12_34 ) );
  DFF_X1 key_c_r_reg_12_35 (.CK( clk ) , .D( key_c_r_11_35 ) , .Q( key_c_r_12_35 ) );
  DFF_X1 key_c_r_reg_12_36 (.CK( clk ) , .D( key_c_r_11_36 ) , .Q( key_c_r_12_36 ) );
  DFF_X1 key_c_r_reg_12_37 (.CK( clk ) , .D( key_c_r_11_37 ) , .Q( key_c_r_12_37 ) );
  DFF_X1 key_c_r_reg_12_38 (.CK( clk ) , .D( key_c_r_11_38 ) , .Q( key_c_r_12_38 ) );
  DFF_X1 key_c_r_reg_12_39 (.CK( clk ) , .D( key_c_r_11_39 ) , .Q( key_c_r_12_39 ) );
  DFF_X1 key_c_r_reg_12_4 (.CK( clk ) , .D( key_c_r_11_4 ) , .Q( key_c_r_12_4 ) );
  DFF_X1 key_c_r_reg_12_40 (.CK( clk ) , .D( key_c_r_11_40 ) , .Q( key_c_r_12_40 ) );
  DFF_X1 key_c_r_reg_12_41 (.CK( clk ) , .D( key_c_r_11_41 ) , .Q( key_c_r_12_41 ) );
  DFF_X1 key_c_r_reg_12_42 (.CK( clk ) , .D( key_c_r_11_42 ) , .Q( key_c_r_12_42 ) );
  DFF_X1 key_c_r_reg_12_43 (.CK( clk ) , .D( key_c_r_11_43 ) , .Q( key_c_r_12_43 ) );
  DFF_X1 key_c_r_reg_12_44 (.CK( clk ) , .D( key_c_r_11_44 ) , .Q( key_c_r_12_44 ) );
  DFF_X1 key_c_r_reg_12_45 (.CK( clk ) , .D( key_c_r_11_45 ) , .Q( key_c_r_12_45 ) );
  DFF_X1 key_c_r_reg_12_46 (.CK( clk ) , .D( key_c_r_11_46 ) , .Q( key_c_r_12_46 ) );
  DFF_X1 key_c_r_reg_12_47 (.CK( clk ) , .D( key_c_r_11_47 ) , .Q( key_c_r_12_47 ) );
  DFF_X1 key_c_r_reg_12_48 (.CK( clk ) , .D( key_c_r_11_48 ) , .Q( key_c_r_12_48 ) );
  DFF_X1 key_c_r_reg_12_49 (.CK( clk ) , .D( key_c_r_11_49 ) , .Q( key_c_r_12_49 ) );
  DFF_X1 key_c_r_reg_12_5 (.CK( clk ) , .D( key_c_r_11_5 ) , .Q( key_c_r_12_5 ) );
  DFF_X1 key_c_r_reg_12_50 (.CK( clk ) , .D( key_c_r_11_50 ) , .Q( key_c_r_12_50 ) );
  DFF_X1 key_c_r_reg_12_51 (.CK( clk ) , .D( key_c_r_11_51 ) , .Q( key_c_r_12_51 ) );
  DFF_X1 key_c_r_reg_12_52 (.CK( clk ) , .D( key_c_r_11_52 ) , .Q( key_c_r_12_52 ) );
  DFF_X1 key_c_r_reg_12_53 (.CK( clk ) , .D( key_c_r_11_53 ) , .Q( key_c_r_12_53 ) );
  DFF_X1 key_c_r_reg_12_54 (.CK( clk ) , .D( key_c_r_11_54 ) , .Q( key_c_r_12_54 ) );
  DFF_X1 key_c_r_reg_12_55 (.CK( clk ) , .D( key_c_r_11_55 ) , .Q( key_c_r_12_55 ) );
  DFF_X1 key_c_r_reg_12_6 (.CK( clk ) , .D( key_c_r_11_6 ) , .Q( key_c_r_12_6 ) );
  DFF_X1 key_c_r_reg_12_7 (.CK( clk ) , .D( key_c_r_11_7 ) , .Q( key_c_r_12_7 ) );
  DFF_X1 key_c_r_reg_12_8 (.CK( clk ) , .D( key_c_r_11_8 ) , .Q( key_c_r_12_8 ) );
  DFF_X1 key_c_r_reg_12_9 (.CK( clk ) , .D( key_c_r_11_9 ) , .Q( key_c_r_12_9 ) );
  DFF_X1 key_c_r_reg_13_0 (.CK( clk ) , .D( key_c_r_12_0 ) , .Q( key_c_r_13_0 ) );
  DFF_X1 key_c_r_reg_13_1 (.CK( clk ) , .D( key_c_r_12_1 ) , .Q( key_c_r_13_1 ) );
  DFF_X1 key_c_r_reg_13_10 (.CK( clk ) , .D( key_c_r_12_10 ) , .Q( key_c_r_13_10 ) );
  DFF_X1 key_c_r_reg_13_11 (.CK( clk ) , .D( key_c_r_12_11 ) , .Q( key_c_r_13_11 ) );
  DFF_X1 key_c_r_reg_13_12 (.CK( clk ) , .D( key_c_r_12_12 ) , .Q( key_c_r_13_12 ) );
  DFF_X1 key_c_r_reg_13_13 (.CK( clk ) , .D( key_c_r_12_13 ) , .Q( key_c_r_13_13 ) );
  DFF_X1 key_c_r_reg_13_14 (.CK( clk ) , .D( key_c_r_12_14 ) , .Q( key_c_r_13_14 ) );
  DFF_X1 key_c_r_reg_13_15 (.CK( clk ) , .D( key_c_r_12_15 ) , .Q( key_c_r_13_15 ) );
  DFF_X1 key_c_r_reg_13_16 (.CK( clk ) , .D( key_c_r_12_16 ) , .Q( key_c_r_13_16 ) );
  DFF_X1 key_c_r_reg_13_17 (.CK( clk ) , .D( key_c_r_12_17 ) , .Q( key_c_r_13_17 ) );
  DFF_X1 key_c_r_reg_13_18 (.CK( clk ) , .D( key_c_r_12_18 ) , .Q( key_c_r_13_18 ) );
  DFF_X1 key_c_r_reg_13_19 (.CK( clk ) , .D( key_c_r_12_19 ) , .Q( key_c_r_13_19 ) );
  DFF_X1 key_c_r_reg_13_2 (.CK( clk ) , .D( key_c_r_12_2 ) , .Q( key_c_r_13_2 ) );
  DFF_X1 key_c_r_reg_13_20 (.CK( clk ) , .D( key_c_r_12_20 ) , .Q( key_c_r_13_20 ) );
  DFF_X1 key_c_r_reg_13_21 (.CK( clk ) , .D( key_c_r_12_21 ) , .Q( key_c_r_13_21 ) );
  DFF_X1 key_c_r_reg_13_22 (.CK( clk ) , .D( key_c_r_12_22 ) , .Q( key_c_r_13_22 ) );
  DFF_X1 key_c_r_reg_13_23 (.CK( clk ) , .D( key_c_r_12_23 ) , .Q( key_c_r_13_23 ) );
  DFF_X1 key_c_r_reg_13_24 (.CK( clk ) , .D( key_c_r_12_24 ) , .Q( key_c_r_13_24 ) );
  DFF_X1 key_c_r_reg_13_25 (.CK( clk ) , .D( key_c_r_12_25 ) , .Q( key_c_r_13_25 ) );
  DFF_X1 key_c_r_reg_13_26 (.CK( clk ) , .D( key_c_r_12_26 ) , .Q( key_c_r_13_26 ) );
  DFF_X1 key_c_r_reg_13_27 (.CK( clk ) , .D( key_c_r_12_27 ) , .Q( key_c_r_13_27 ) );
  DFF_X1 key_c_r_reg_13_28 (.CK( clk ) , .D( key_c_r_12_28 ) , .Q( key_c_r_13_28 ) );
  DFF_X1 key_c_r_reg_13_29 (.CK( clk ) , .D( key_c_r_12_29 ) , .Q( key_c_r_13_29 ) );
  DFF_X1 key_c_r_reg_13_3 (.CK( clk ) , .D( key_c_r_12_3 ) , .Q( key_c_r_13_3 ) );
  DFF_X1 key_c_r_reg_13_30 (.CK( clk ) , .D( key_c_r_12_30 ) , .Q( key_c_r_13_30 ) );
  DFF_X1 key_c_r_reg_13_31 (.CK( clk ) , .D( key_c_r_12_31 ) , .Q( key_c_r_13_31 ) );
  DFF_X1 key_c_r_reg_13_32 (.CK( clk ) , .D( key_c_r_12_32 ) , .Q( key_c_r_13_32 ) );
  DFF_X1 key_c_r_reg_13_33 (.CK( clk ) , .D( key_c_r_12_33 ) , .Q( key_c_r_13_33 ) );
  DFF_X1 key_c_r_reg_13_34 (.CK( clk ) , .D( key_c_r_12_34 ) , .Q( key_c_r_13_34 ) );
  DFF_X1 key_c_r_reg_13_35 (.CK( clk ) , .D( key_c_r_12_35 ) , .Q( key_c_r_13_35 ) );
  DFF_X1 key_c_r_reg_13_36 (.CK( clk ) , .D( key_c_r_12_36 ) , .Q( key_c_r_13_36 ) );
  DFF_X1 key_c_r_reg_13_37 (.CK( clk ) , .D( key_c_r_12_37 ) , .Q( key_c_r_13_37 ) );
  DFF_X1 key_c_r_reg_13_38 (.CK( clk ) , .D( key_c_r_12_38 ) , .Q( key_c_r_13_38 ) );
  DFF_X1 key_c_r_reg_13_39 (.CK( clk ) , .D( key_c_r_12_39 ) , .Q( key_c_r_13_39 ) );
  DFF_X1 key_c_r_reg_13_4 (.CK( clk ) , .D( key_c_r_12_4 ) , .Q( key_c_r_13_4 ) );
  DFF_X1 key_c_r_reg_13_40 (.CK( clk ) , .D( key_c_r_12_40 ) , .Q( key_c_r_13_40 ) );
  DFF_X1 key_c_r_reg_13_41 (.CK( clk ) , .D( key_c_r_12_41 ) , .Q( key_c_r_13_41 ) );
  DFF_X1 key_c_r_reg_13_42 (.CK( clk ) , .D( key_c_r_12_42 ) , .Q( key_c_r_13_42 ) );
  DFF_X1 key_c_r_reg_13_43 (.CK( clk ) , .D( key_c_r_12_43 ) , .Q( key_c_r_13_43 ) );
  DFF_X1 key_c_r_reg_13_44 (.CK( clk ) , .D( key_c_r_12_44 ) , .Q( key_c_r_13_44 ) );
  DFF_X1 key_c_r_reg_13_45 (.CK( clk ) , .D( key_c_r_12_45 ) , .Q( key_c_r_13_45 ) );
  DFF_X1 key_c_r_reg_13_46 (.CK( clk ) , .D( key_c_r_12_46 ) , .Q( key_c_r_13_46 ) );
  DFF_X1 key_c_r_reg_13_47 (.CK( clk ) , .D( key_c_r_12_47 ) , .Q( key_c_r_13_47 ) );
  DFF_X1 key_c_r_reg_13_48 (.CK( clk ) , .D( key_c_r_12_48 ) , .Q( key_c_r_13_48 ) );
  DFF_X1 key_c_r_reg_13_49 (.CK( clk ) , .D( key_c_r_12_49 ) , .Q( key_c_r_13_49 ) );
  DFF_X1 key_c_r_reg_13_5 (.CK( clk ) , .D( key_c_r_12_5 ) , .Q( key_c_r_13_5 ) );
  DFF_X1 key_c_r_reg_13_50 (.CK( clk ) , .D( key_c_r_12_50 ) , .Q( key_c_r_13_50 ) );
  DFF_X1 key_c_r_reg_13_51 (.CK( clk ) , .D( key_c_r_12_51 ) , .Q( key_c_r_13_51 ) );
  DFF_X1 key_c_r_reg_13_52 (.CK( clk ) , .D( key_c_r_12_52 ) , .Q( key_c_r_13_52 ) );
  DFF_X1 key_c_r_reg_13_53 (.CK( clk ) , .D( key_c_r_12_53 ) , .Q( key_c_r_13_53 ) );
  DFF_X1 key_c_r_reg_13_54 (.CK( clk ) , .D( key_c_r_12_54 ) , .Q( key_c_r_13_54 ) );
  DFF_X1 key_c_r_reg_13_55 (.CK( clk ) , .D( key_c_r_12_55 ) , .Q( key_c_r_13_55 ) );
  DFF_X1 key_c_r_reg_13_6 (.CK( clk ) , .D( key_c_r_12_6 ) , .Q( key_c_r_13_6 ) );
  DFF_X1 key_c_r_reg_13_7 (.CK( clk ) , .D( key_c_r_12_7 ) , .Q( key_c_r_13_7 ) );
  DFF_X1 key_c_r_reg_13_8 (.CK( clk ) , .D( key_c_r_12_8 ) , .Q( key_c_r_13_8 ) );
  DFF_X1 key_c_r_reg_13_9 (.CK( clk ) , .D( key_c_r_12_9 ) , .Q( key_c_r_13_9 ) );
  DFF_X1 key_c_r_reg_14_0 (.CK( clk ) , .D( key_c_r_13_0 ) , .Q( key_c_r_14_0 ) );
  DFF_X1 key_c_r_reg_14_1 (.CK( clk ) , .D( key_c_r_13_1 ) , .Q( key_c_r_14_1 ) );
  DFF_X1 key_c_r_reg_14_10 (.CK( clk ) , .D( key_c_r_13_10 ) , .Q( key_c_r_14_10 ) );
  DFF_X1 key_c_r_reg_14_11 (.CK( clk ) , .D( key_c_r_13_11 ) , .Q( key_c_r_14_11 ) );
  DFF_X1 key_c_r_reg_14_12 (.CK( clk ) , .D( key_c_r_13_12 ) , .Q( key_c_r_14_12 ) );
  DFF_X1 key_c_r_reg_14_13 (.CK( clk ) , .D( key_c_r_13_13 ) , .Q( key_c_r_14_13 ) );
  DFF_X1 key_c_r_reg_14_14 (.CK( clk ) , .D( key_c_r_13_14 ) , .Q( key_c_r_14_14 ) );
  DFF_X1 key_c_r_reg_14_15 (.CK( clk ) , .D( key_c_r_13_15 ) , .Q( key_c_r_14_15 ) );
  DFF_X1 key_c_r_reg_14_16 (.CK( clk ) , .D( key_c_r_13_16 ) , .Q( key_c_r_14_16 ) );
  DFF_X1 key_c_r_reg_14_17 (.CK( clk ) , .D( key_c_r_13_17 ) , .Q( key_c_r_14_17 ) );
  DFF_X1 key_c_r_reg_14_18 (.CK( clk ) , .D( key_c_r_13_18 ) , .Q( key_c_r_14_18 ) );
  DFF_X1 key_c_r_reg_14_19 (.CK( clk ) , .D( key_c_r_13_19 ) , .Q( key_c_r_14_19 ) );
  DFF_X1 key_c_r_reg_14_2 (.CK( clk ) , .D( key_c_r_13_2 ) , .Q( key_c_r_14_2 ) );
  DFF_X1 key_c_r_reg_14_20 (.CK( clk ) , .D( key_c_r_13_20 ) , .Q( key_c_r_14_20 ) );
  DFF_X1 key_c_r_reg_14_21 (.CK( clk ) , .D( key_c_r_13_21 ) , .Q( key_c_r_14_21 ) );
  DFF_X1 key_c_r_reg_14_22 (.CK( clk ) , .D( key_c_r_13_22 ) , .Q( key_c_r_14_22 ) );
  DFF_X1 key_c_r_reg_14_23 (.CK( clk ) , .D( key_c_r_13_23 ) , .Q( key_c_r_14_23 ) );
  DFF_X1 key_c_r_reg_14_24 (.CK( clk ) , .D( key_c_r_13_24 ) , .Q( key_c_r_14_24 ) );
  DFF_X1 key_c_r_reg_14_25 (.CK( clk ) , .D( key_c_r_13_25 ) , .Q( key_c_r_14_25 ) );
  DFF_X1 key_c_r_reg_14_26 (.CK( clk ) , .D( key_c_r_13_26 ) , .Q( key_c_r_14_26 ) );
  DFF_X1 key_c_r_reg_14_27 (.CK( clk ) , .D( key_c_r_13_27 ) , .Q( key_c_r_14_27 ) );
  DFF_X1 key_c_r_reg_14_28 (.CK( clk ) , .D( key_c_r_13_28 ) , .Q( key_c_r_14_28 ) );
  DFF_X1 key_c_r_reg_14_29 (.CK( clk ) , .D( key_c_r_13_29 ) , .Q( key_c_r_14_29 ) );
  DFF_X1 key_c_r_reg_14_3 (.CK( clk ) , .D( key_c_r_13_3 ) , .Q( key_c_r_14_3 ) );
  DFF_X1 key_c_r_reg_14_30 (.CK( clk ) , .D( key_c_r_13_30 ) , .Q( key_c_r_14_30 ) );
  DFF_X1 key_c_r_reg_14_31 (.CK( clk ) , .D( key_c_r_13_31 ) , .Q( key_c_r_14_31 ) );
  DFF_X1 key_c_r_reg_14_32 (.CK( clk ) , .D( key_c_r_13_32 ) , .Q( key_c_r_14_32 ) );
  DFF_X1 key_c_r_reg_14_33 (.CK( clk ) , .D( key_c_r_13_33 ) , .Q( key_c_r_14_33 ) );
  DFF_X1 key_c_r_reg_14_34 (.CK( clk ) , .D( key_c_r_13_34 ) , .Q( key_c_r_14_34 ) );
  DFF_X1 key_c_r_reg_14_35 (.CK( clk ) , .D( key_c_r_13_35 ) , .Q( key_c_r_14_35 ) );
  DFF_X1 key_c_r_reg_14_36 (.CK( clk ) , .D( key_c_r_13_36 ) , .Q( key_c_r_14_36 ) );
  DFF_X1 key_c_r_reg_14_37 (.CK( clk ) , .D( key_c_r_13_37 ) , .Q( key_c_r_14_37 ) );
  DFF_X1 key_c_r_reg_14_38 (.CK( clk ) , .D( key_c_r_13_38 ) , .Q( key_c_r_14_38 ) );
  DFF_X1 key_c_r_reg_14_39 (.CK( clk ) , .D( key_c_r_13_39 ) , .Q( key_c_r_14_39 ) );
  DFF_X1 key_c_r_reg_14_4 (.CK( clk ) , .D( key_c_r_13_4 ) , .Q( key_c_r_14_4 ) );
  DFF_X1 key_c_r_reg_14_40 (.CK( clk ) , .D( key_c_r_13_40 ) , .Q( key_c_r_14_40 ) );
  DFF_X1 key_c_r_reg_14_41 (.CK( clk ) , .D( key_c_r_13_41 ) , .Q( key_c_r_14_41 ) );
  DFF_X1 key_c_r_reg_14_42 (.CK( clk ) , .D( key_c_r_13_42 ) , .Q( key_c_r_14_42 ) );
  DFF_X1 key_c_r_reg_14_43 (.CK( clk ) , .D( key_c_r_13_43 ) , .Q( key_c_r_14_43 ) );
  DFF_X1 key_c_r_reg_14_44 (.CK( clk ) , .D( key_c_r_13_44 ) , .Q( key_c_r_14_44 ) );
  DFF_X1 key_c_r_reg_14_45 (.CK( clk ) , .D( key_c_r_13_45 ) , .Q( key_c_r_14_45 ) );
  DFF_X1 key_c_r_reg_14_46 (.CK( clk ) , .D( key_c_r_13_46 ) , .Q( key_c_r_14_46 ) );
  DFF_X1 key_c_r_reg_14_47 (.CK( clk ) , .D( key_c_r_13_47 ) , .Q( key_c_r_14_47 ) );
  DFF_X1 key_c_r_reg_14_48 (.CK( clk ) , .D( key_c_r_13_48 ) , .Q( key_c_r_14_48 ) );
  DFF_X1 key_c_r_reg_14_49 (.CK( clk ) , .D( key_c_r_13_49 ) , .Q( key_c_r_14_49 ) );
  DFF_X1 key_c_r_reg_14_5 (.CK( clk ) , .D( key_c_r_13_5 ) , .Q( key_c_r_14_5 ) );
  DFF_X1 key_c_r_reg_14_50 (.CK( clk ) , .D( key_c_r_13_50 ) , .Q( key_c_r_14_50 ) );
  DFF_X1 key_c_r_reg_14_51 (.CK( clk ) , .D( key_c_r_13_51 ) , .Q( key_c_r_14_51 ) );
  DFF_X1 key_c_r_reg_14_52 (.CK( clk ) , .D( key_c_r_13_52 ) , .Q( key_c_r_14_52 ) );
  DFF_X1 key_c_r_reg_14_53 (.CK( clk ) , .D( key_c_r_13_53 ) , .Q( key_c_r_14_53 ) );
  DFF_X1 key_c_r_reg_14_54 (.CK( clk ) , .D( key_c_r_13_54 ) , .Q( key_c_r_14_54 ) );
  DFF_X1 key_c_r_reg_14_55 (.CK( clk ) , .D( key_c_r_13_55 ) , .Q( key_c_r_14_55 ) );
  DFF_X1 key_c_r_reg_14_6 (.CK( clk ) , .D( key_c_r_13_6 ) , .Q( key_c_r_14_6 ) );
  DFF_X1 key_c_r_reg_14_7 (.CK( clk ) , .D( key_c_r_13_7 ) , .Q( key_c_r_14_7 ) );
  DFF_X1 key_c_r_reg_14_8 (.CK( clk ) , .D( key_c_r_13_8 ) , .Q( key_c_r_14_8 ) );
  DFF_X1 key_c_r_reg_14_9 (.CK( clk ) , .D( key_c_r_13_9 ) , .Q( key_c_r_14_9 ) );
  DFF_X1 key_c_r_reg_15_0 (.CK( clk ) , .D( key_c_r_14_0 ) , .Q( key_c_r_15_0 ) );
  DFF_X1 key_c_r_reg_15_1 (.CK( clk ) , .D( key_c_r_14_1 ) , .Q( key_c_r_15_1 ) );
  DFF_X1 key_c_r_reg_15_10 (.CK( clk ) , .D( key_c_r_14_10 ) , .Q( key_c_r_15_10 ) );
  DFF_X1 key_c_r_reg_15_11 (.CK( clk ) , .D( key_c_r_14_11 ) , .Q( key_c_r_15_11 ) );
  DFF_X1 key_c_r_reg_15_12 (.CK( clk ) , .D( key_c_r_14_12 ) , .Q( key_c_r_15_12 ) );
  DFF_X1 key_c_r_reg_15_13 (.CK( clk ) , .D( key_c_r_14_13 ) , .Q( key_c_r_15_13 ) );
  DFF_X1 key_c_r_reg_15_14 (.CK( clk ) , .D( key_c_r_14_14 ) , .Q( key_c_r_15_14 ) );
  DFF_X1 key_c_r_reg_15_15 (.CK( clk ) , .D( key_c_r_14_15 ) , .Q( key_c_r_15_15 ) );
  DFF_X1 key_c_r_reg_15_16 (.CK( clk ) , .D( key_c_r_14_16 ) , .Q( key_c_r_15_16 ) );
  DFF_X1 key_c_r_reg_15_17 (.CK( clk ) , .D( key_c_r_14_17 ) , .Q( key_c_r_15_17 ) );
  DFF_X1 key_c_r_reg_15_18 (.CK( clk ) , .D( key_c_r_14_18 ) , .Q( key_c_r_15_18 ) );
  DFF_X1 key_c_r_reg_15_19 (.CK( clk ) , .D( key_c_r_14_19 ) , .Q( key_c_r_15_19 ) );
  DFF_X1 key_c_r_reg_15_2 (.CK( clk ) , .D( key_c_r_14_2 ) , .Q( key_c_r_15_2 ) );
  DFF_X1 key_c_r_reg_15_20 (.CK( clk ) , .D( key_c_r_14_20 ) , .Q( key_c_r_15_20 ) );
  DFF_X1 key_c_r_reg_15_21 (.CK( clk ) , .D( key_c_r_14_21 ) , .Q( key_c_r_15_21 ) );
  DFF_X1 key_c_r_reg_15_22 (.CK( clk ) , .D( key_c_r_14_22 ) , .Q( key_c_r_15_22 ) );
  DFF_X1 key_c_r_reg_15_23 (.CK( clk ) , .D( key_c_r_14_23 ) , .Q( key_c_r_15_23 ) );
  DFF_X1 key_c_r_reg_15_24 (.CK( clk ) , .D( key_c_r_14_24 ) , .Q( key_c_r_15_24 ) );
  DFF_X1 key_c_r_reg_15_25 (.CK( clk ) , .D( key_c_r_14_25 ) , .Q( key_c_r_15_25 ) );
  DFF_X1 key_c_r_reg_15_26 (.CK( clk ) , .D( key_c_r_14_26 ) , .Q( key_c_r_15_26 ) );
  DFF_X1 key_c_r_reg_15_27 (.CK( clk ) , .D( key_c_r_14_27 ) , .Q( key_c_r_15_27 ) );
  DFF_X1 key_c_r_reg_15_28 (.CK( clk ) , .D( key_c_r_14_28 ) , .Q( key_c_r_15_28 ) );
  DFF_X1 key_c_r_reg_15_29 (.CK( clk ) , .D( key_c_r_14_29 ) , .Q( key_c_r_15_29 ) );
  DFF_X1 key_c_r_reg_15_3 (.CK( clk ) , .D( key_c_r_14_3 ) , .Q( key_c_r_15_3 ) );
  DFF_X1 key_c_r_reg_15_30 (.CK( clk ) , .D( key_c_r_14_30 ) , .Q( key_c_r_15_30 ) );
  DFF_X1 key_c_r_reg_15_31 (.CK( clk ) , .D( key_c_r_14_31 ) , .Q( key_c_r_15_31 ) );
  DFF_X1 key_c_r_reg_15_32 (.CK( clk ) , .D( key_c_r_14_32 ) , .Q( key_c_r_15_32 ) );
  DFF_X1 key_c_r_reg_15_33 (.CK( clk ) , .D( key_c_r_14_33 ) , .Q( key_c_r_15_33 ) );
  DFF_X1 key_c_r_reg_15_34 (.CK( clk ) , .D( key_c_r_14_34 ) , .Q( key_c_r_15_34 ) );
  DFF_X1 key_c_r_reg_15_35 (.CK( clk ) , .D( key_c_r_14_35 ) , .Q( key_c_r_15_35 ) );
  DFF_X1 key_c_r_reg_15_36 (.CK( clk ) , .D( key_c_r_14_36 ) , .Q( key_c_r_15_36 ) );
  DFF_X1 key_c_r_reg_15_37 (.CK( clk ) , .D( key_c_r_14_37 ) , .Q( key_c_r_15_37 ) );
  DFF_X1 key_c_r_reg_15_38 (.CK( clk ) , .D( key_c_r_14_38 ) , .Q( key_c_r_15_38 ) );
  DFF_X1 key_c_r_reg_15_39 (.CK( clk ) , .D( key_c_r_14_39 ) , .Q( key_c_r_15_39 ) );
  DFF_X1 key_c_r_reg_15_4 (.CK( clk ) , .D( key_c_r_14_4 ) , .Q( key_c_r_15_4 ) );
  DFF_X1 key_c_r_reg_15_40 (.CK( clk ) , .D( key_c_r_14_40 ) , .Q( key_c_r_15_40 ) );
  DFF_X1 key_c_r_reg_15_41 (.CK( clk ) , .D( key_c_r_14_41 ) , .Q( key_c_r_15_41 ) );
  DFF_X1 key_c_r_reg_15_42 (.CK( clk ) , .D( key_c_r_14_42 ) , .Q( key_c_r_15_42 ) );
  DFF_X1 key_c_r_reg_15_43 (.CK( clk ) , .D( key_c_r_14_43 ) , .Q( key_c_r_15_43 ) );
  DFF_X1 key_c_r_reg_15_44 (.CK( clk ) , .D( key_c_r_14_44 ) , .Q( key_c_r_15_44 ) );
  DFF_X1 key_c_r_reg_15_45 (.CK( clk ) , .D( key_c_r_14_45 ) , .Q( key_c_r_15_45 ) );
  DFF_X1 key_c_r_reg_15_46 (.CK( clk ) , .D( key_c_r_14_46 ) , .Q( key_c_r_15_46 ) );
  DFF_X1 key_c_r_reg_15_47 (.CK( clk ) , .D( key_c_r_14_47 ) , .Q( key_c_r_15_47 ) );
  DFF_X1 key_c_r_reg_15_48 (.CK( clk ) , .D( key_c_r_14_48 ) , .Q( key_c_r_15_48 ) );
  DFF_X1 key_c_r_reg_15_49 (.CK( clk ) , .D( key_c_r_14_49 ) , .Q( key_c_r_15_49 ) );
  DFF_X1 key_c_r_reg_15_5 (.CK( clk ) , .D( key_c_r_14_5 ) , .Q( key_c_r_15_5 ) );
  DFF_X1 key_c_r_reg_15_50 (.CK( clk ) , .D( key_c_r_14_50 ) , .Q( key_c_r_15_50 ) );
  DFF_X1 key_c_r_reg_15_51 (.CK( clk ) , .D( key_c_r_14_51 ) , .Q( key_c_r_15_51 ) );
  DFF_X1 key_c_r_reg_15_52 (.CK( clk ) , .D( key_c_r_14_52 ) , .Q( key_c_r_15_52 ) );
  DFF_X1 key_c_r_reg_15_53 (.CK( clk ) , .D( key_c_r_14_53 ) , .Q( key_c_r_15_53 ) );
  DFF_X1 key_c_r_reg_15_54 (.CK( clk ) , .D( key_c_r_14_54 ) , .Q( key_c_r_15_54 ) );
  DFF_X1 key_c_r_reg_15_55 (.CK( clk ) , .D( key_c_r_14_55 ) , .Q( key_c_r_15_55 ) );
  DFF_X1 key_c_r_reg_15_6 (.CK( clk ) , .D( key_c_r_14_6 ) , .Q( key_c_r_15_6 ) );
  DFF_X1 key_c_r_reg_15_7 (.CK( clk ) , .D( key_c_r_14_7 ) , .Q( key_c_r_15_7 ) );
  DFF_X1 key_c_r_reg_15_8 (.CK( clk ) , .D( key_c_r_14_8 ) , .Q( key_c_r_15_8 ) );
  DFF_X1 key_c_r_reg_15_9 (.CK( clk ) , .D( key_c_r_14_9 ) , .Q( key_c_r_15_9 ) );
  DFF_X1 key_c_r_reg_16_0 (.CK( clk ) , .D( key_c_r_15_0 ) , .Q( key_c_r_16_0 ) );
  DFF_X1 key_c_r_reg_16_1 (.CK( clk ) , .D( key_c_r_15_1 ) , .Q( key_c_r_16_1 ) );
  DFF_X1 key_c_r_reg_16_10 (.CK( clk ) , .D( key_c_r_15_10 ) , .Q( key_c_r_16_10 ) );
  DFF_X1 key_c_r_reg_16_11 (.CK( clk ) , .D( key_c_r_15_11 ) , .Q( key_c_r_16_11 ) );
  DFF_X1 key_c_r_reg_16_12 (.CK( clk ) , .D( key_c_r_15_12 ) , .Q( key_c_r_16_12 ) );
  DFF_X1 key_c_r_reg_16_13 (.CK( clk ) , .D( key_c_r_15_13 ) , .Q( key_c_r_16_13 ) );
  DFF_X1 key_c_r_reg_16_14 (.CK( clk ) , .D( key_c_r_15_14 ) , .Q( key_c_r_16_14 ) );
  DFF_X1 key_c_r_reg_16_15 (.CK( clk ) , .D( key_c_r_15_15 ) , .Q( key_c_r_16_15 ) );
  DFF_X1 key_c_r_reg_16_16 (.CK( clk ) , .D( key_c_r_15_16 ) , .Q( key_c_r_16_16 ) );
  DFF_X1 key_c_r_reg_16_17 (.CK( clk ) , .D( key_c_r_15_17 ) , .Q( key_c_r_16_17 ) );
  DFF_X1 key_c_r_reg_16_18 (.CK( clk ) , .D( key_c_r_15_18 ) , .Q( key_c_r_16_18 ) );
  DFF_X1 key_c_r_reg_16_19 (.CK( clk ) , .D( key_c_r_15_19 ) , .Q( key_c_r_16_19 ) );
  DFF_X1 key_c_r_reg_16_2 (.CK( clk ) , .D( key_c_r_15_2 ) , .Q( key_c_r_16_2 ) );
  DFF_X1 key_c_r_reg_16_20 (.CK( clk ) , .D( key_c_r_15_20 ) , .Q( key_c_r_16_20 ) );
  DFF_X1 key_c_r_reg_16_21 (.CK( clk ) , .D( key_c_r_15_21 ) , .Q( key_c_r_16_21 ) );
  DFF_X1 key_c_r_reg_16_22 (.CK( clk ) , .D( key_c_r_15_22 ) , .Q( key_c_r_16_22 ) );
  DFF_X1 key_c_r_reg_16_23 (.CK( clk ) , .D( key_c_r_15_23 ) , .Q( key_c_r_16_23 ) );
  DFF_X1 key_c_r_reg_16_24 (.CK( clk ) , .D( key_c_r_15_24 ) , .Q( key_c_r_16_24 ) );
  DFF_X1 key_c_r_reg_16_25 (.CK( clk ) , .D( key_c_r_15_25 ) , .Q( key_c_r_16_25 ) );
  DFF_X1 key_c_r_reg_16_26 (.CK( clk ) , .D( key_c_r_15_26 ) , .Q( key_c_r_16_26 ) );
  DFF_X1 key_c_r_reg_16_27 (.CK( clk ) , .D( key_c_r_15_27 ) , .Q( key_c_r_16_27 ) );
  DFF_X1 key_c_r_reg_16_28 (.CK( clk ) , .D( key_c_r_15_28 ) , .Q( key_c_r_16_28 ) );
  DFF_X1 key_c_r_reg_16_29 (.CK( clk ) , .D( key_c_r_15_29 ) , .Q( key_c_r_16_29 ) );
  DFF_X1 key_c_r_reg_16_3 (.CK( clk ) , .D( key_c_r_15_3 ) , .Q( key_c_r_16_3 ) );
  DFF_X1 key_c_r_reg_16_30 (.CK( clk ) , .D( key_c_r_15_30 ) , .Q( key_c_r_16_30 ) );
  DFF_X1 key_c_r_reg_16_31 (.CK( clk ) , .D( key_c_r_15_31 ) , .Q( key_c_r_16_31 ) );
  DFF_X1 key_c_r_reg_16_32 (.CK( clk ) , .D( key_c_r_15_32 ) , .Q( key_c_r_16_32 ) );
  DFF_X1 key_c_r_reg_16_33 (.CK( clk ) , .D( key_c_r_15_33 ) , .Q( key_c_r_16_33 ) );
  DFF_X1 key_c_r_reg_16_34 (.CK( clk ) , .D( key_c_r_15_34 ) , .Q( key_c_r_16_34 ) );
  DFF_X1 key_c_r_reg_16_35 (.CK( clk ) , .D( key_c_r_15_35 ) , .Q( key_c_r_16_35 ) );
  DFF_X1 key_c_r_reg_16_36 (.CK( clk ) , .D( key_c_r_15_36 ) , .Q( key_c_r_16_36 ) );
  DFF_X1 key_c_r_reg_16_37 (.CK( clk ) , .D( key_c_r_15_37 ) , .Q( key_c_r_16_37 ) );
  DFF_X1 key_c_r_reg_16_38 (.CK( clk ) , .D( key_c_r_15_38 ) , .Q( key_c_r_16_38 ) );
  DFF_X1 key_c_r_reg_16_39 (.CK( clk ) , .D( key_c_r_15_39 ) , .Q( key_c_r_16_39 ) );
  DFF_X1 key_c_r_reg_16_4 (.CK( clk ) , .D( key_c_r_15_4 ) , .Q( key_c_r_16_4 ) );
  DFF_X1 key_c_r_reg_16_40 (.CK( clk ) , .D( key_c_r_15_40 ) , .Q( key_c_r_16_40 ) );
  DFF_X1 key_c_r_reg_16_41 (.CK( clk ) , .D( key_c_r_15_41 ) , .Q( key_c_r_16_41 ) );
  DFF_X1 key_c_r_reg_16_42 (.CK( clk ) , .D( key_c_r_15_42 ) , .Q( key_c_r_16_42 ) );
  DFF_X1 key_c_r_reg_16_43 (.CK( clk ) , .D( key_c_r_15_43 ) , .Q( key_c_r_16_43 ) );
  DFF_X1 key_c_r_reg_16_44 (.CK( clk ) , .D( key_c_r_15_44 ) , .Q( key_c_r_16_44 ) );
  DFF_X1 key_c_r_reg_16_45 (.CK( clk ) , .D( key_c_r_15_45 ) , .Q( key_c_r_16_45 ) );
  DFF_X1 key_c_r_reg_16_46 (.CK( clk ) , .D( key_c_r_15_46 ) , .Q( key_c_r_16_46 ) );
  DFF_X1 key_c_r_reg_16_47 (.CK( clk ) , .D( key_c_r_15_47 ) , .Q( key_c_r_16_47 ) );
  DFF_X1 key_c_r_reg_16_48 (.CK( clk ) , .D( key_c_r_15_48 ) , .Q( key_c_r_16_48 ) );
  DFF_X1 key_c_r_reg_16_49 (.CK( clk ) , .D( key_c_r_15_49 ) , .Q( key_c_r_16_49 ) );
  DFF_X1 key_c_r_reg_16_5 (.CK( clk ) , .D( key_c_r_15_5 ) , .Q( key_c_r_16_5 ) );
  DFF_X1 key_c_r_reg_16_50 (.CK( clk ) , .D( key_c_r_15_50 ) , .Q( key_c_r_16_50 ) );
  DFF_X1 key_c_r_reg_16_51 (.CK( clk ) , .D( key_c_r_15_51 ) , .Q( key_c_r_16_51 ) );
  DFF_X1 key_c_r_reg_16_52 (.CK( clk ) , .D( key_c_r_15_52 ) , .Q( key_c_r_16_52 ) );
  DFF_X1 key_c_r_reg_16_53 (.CK( clk ) , .D( key_c_r_15_53 ) , .Q( key_c_r_16_53 ) );
  DFF_X1 key_c_r_reg_16_54 (.CK( clk ) , .D( key_c_r_15_54 ) , .Q( key_c_r_16_54 ) );
  DFF_X1 key_c_r_reg_16_55 (.CK( clk ) , .D( key_c_r_15_55 ) , .Q( key_c_r_16_55 ) );
  DFF_X1 key_c_r_reg_16_6 (.CK( clk ) , .D( key_c_r_15_6 ) , .Q( key_c_r_16_6 ) );
  DFF_X1 key_c_r_reg_16_7 (.CK( clk ) , .D( key_c_r_15_7 ) , .Q( key_c_r_16_7 ) );
  DFF_X1 key_c_r_reg_16_8 (.CK( clk ) , .D( key_c_r_15_8 ) , .Q( key_c_r_16_8 ) );
  DFF_X1 key_c_r_reg_16_9 (.CK( clk ) , .D( key_c_r_15_9 ) , .Q( key_c_r_16_9 ) );
  DFF_X1 key_c_r_reg_17_0 (.CK( clk ) , .D( key_c_r_16_0 ) , .Q( key_c_r_17_0 ) );
  DFF_X1 key_c_r_reg_17_1 (.CK( clk ) , .D( key_c_r_16_1 ) , .Q( key_c_r_17_1 ) );
  DFF_X1 key_c_r_reg_17_10 (.CK( clk ) , .D( key_c_r_16_10 ) , .Q( key_c_r_17_10 ) );
  DFF_X1 key_c_r_reg_17_11 (.CK( clk ) , .D( key_c_r_16_11 ) , .Q( key_c_r_17_11 ) );
  DFF_X1 key_c_r_reg_17_12 (.CK( clk ) , .D( key_c_r_16_12 ) , .Q( key_c_r_17_12 ) );
  DFF_X1 key_c_r_reg_17_13 (.CK( clk ) , .D( key_c_r_16_13 ) , .Q( key_c_r_17_13 ) );
  DFF_X1 key_c_r_reg_17_14 (.CK( clk ) , .D( key_c_r_16_14 ) , .Q( key_c_r_17_14 ) );
  DFF_X1 key_c_r_reg_17_15 (.CK( clk ) , .D( key_c_r_16_15 ) , .Q( key_c_r_17_15 ) );
  DFF_X1 key_c_r_reg_17_16 (.CK( clk ) , .D( key_c_r_16_16 ) , .Q( key_c_r_17_16 ) );
  DFF_X1 key_c_r_reg_17_17 (.CK( clk ) , .D( key_c_r_16_17 ) , .Q( key_c_r_17_17 ) );
  DFF_X1 key_c_r_reg_17_18 (.CK( clk ) , .D( key_c_r_16_18 ) , .Q( key_c_r_17_18 ) );
  DFF_X1 key_c_r_reg_17_19 (.CK( clk ) , .D( key_c_r_16_19 ) , .Q( key_c_r_17_19 ) );
  DFF_X1 key_c_r_reg_17_2 (.CK( clk ) , .D( key_c_r_16_2 ) , .Q( key_c_r_17_2 ) );
  DFF_X1 key_c_r_reg_17_20 (.CK( clk ) , .D( key_c_r_16_20 ) , .Q( key_c_r_17_20 ) );
  DFF_X1 key_c_r_reg_17_21 (.CK( clk ) , .D( key_c_r_16_21 ) , .Q( key_c_r_17_21 ) );
  DFF_X1 key_c_r_reg_17_22 (.CK( clk ) , .D( key_c_r_16_22 ) , .Q( key_c_r_17_22 ) );
  DFF_X1 key_c_r_reg_17_23 (.CK( clk ) , .D( key_c_r_16_23 ) , .Q( key_c_r_17_23 ) );
  DFF_X1 key_c_r_reg_17_24 (.CK( clk ) , .D( key_c_r_16_24 ) , .Q( key_c_r_17_24 ) );
  DFF_X1 key_c_r_reg_17_25 (.CK( clk ) , .D( key_c_r_16_25 ) , .Q( key_c_r_17_25 ) );
  DFF_X1 key_c_r_reg_17_26 (.CK( clk ) , .D( key_c_r_16_26 ) , .Q( key_c_r_17_26 ) );
  DFF_X1 key_c_r_reg_17_27 (.CK( clk ) , .D( key_c_r_16_27 ) , .Q( key_c_r_17_27 ) );
  DFF_X1 key_c_r_reg_17_28 (.CK( clk ) , .D( key_c_r_16_28 ) , .Q( key_c_r_17_28 ) );
  DFF_X1 key_c_r_reg_17_29 (.CK( clk ) , .D( key_c_r_16_29 ) , .Q( key_c_r_17_29 ) );
  DFF_X1 key_c_r_reg_17_3 (.CK( clk ) , .D( key_c_r_16_3 ) , .Q( key_c_r_17_3 ) );
  DFF_X1 key_c_r_reg_17_30 (.CK( clk ) , .D( key_c_r_16_30 ) , .Q( key_c_r_17_30 ) );
  DFF_X1 key_c_r_reg_17_31 (.CK( clk ) , .D( key_c_r_16_31 ) , .Q( key_c_r_17_31 ) );
  DFF_X1 key_c_r_reg_17_32 (.CK( clk ) , .D( key_c_r_16_32 ) , .Q( key_c_r_17_32 ) );
  DFF_X1 key_c_r_reg_17_33 (.CK( clk ) , .D( key_c_r_16_33 ) , .Q( key_c_r_17_33 ) );
  DFF_X1 key_c_r_reg_17_34 (.CK( clk ) , .D( key_c_r_16_34 ) , .Q( key_c_r_17_34 ) );
  DFF_X1 key_c_r_reg_17_35 (.CK( clk ) , .D( key_c_r_16_35 ) , .Q( key_c_r_17_35 ) );
  DFF_X1 key_c_r_reg_17_36 (.CK( clk ) , .D( key_c_r_16_36 ) , .Q( key_c_r_17_36 ) );
  DFF_X1 key_c_r_reg_17_37 (.CK( clk ) , .D( key_c_r_16_37 ) , .Q( key_c_r_17_37 ) );
  DFF_X1 key_c_r_reg_17_38 (.CK( clk ) , .D( key_c_r_16_38 ) , .Q( key_c_r_17_38 ) );
  DFF_X1 key_c_r_reg_17_39 (.CK( clk ) , .D( key_c_r_16_39 ) , .Q( key_c_r_17_39 ) );
  DFF_X1 key_c_r_reg_17_4 (.CK( clk ) , .D( key_c_r_16_4 ) , .Q( key_c_r_17_4 ) );
  DFF_X1 key_c_r_reg_17_40 (.CK( clk ) , .D( key_c_r_16_40 ) , .Q( key_c_r_17_40 ) );
  DFF_X1 key_c_r_reg_17_41 (.CK( clk ) , .D( key_c_r_16_41 ) , .Q( key_c_r_17_41 ) );
  DFF_X1 key_c_r_reg_17_42 (.CK( clk ) , .D( key_c_r_16_42 ) , .Q( key_c_r_17_42 ) );
  DFF_X1 key_c_r_reg_17_43 (.CK( clk ) , .D( key_c_r_16_43 ) , .Q( key_c_r_17_43 ) );
  DFF_X1 key_c_r_reg_17_44 (.CK( clk ) , .D( key_c_r_16_44 ) , .Q( key_c_r_17_44 ) );
  DFF_X1 key_c_r_reg_17_45 (.CK( clk ) , .D( key_c_r_16_45 ) , .Q( key_c_r_17_45 ) );
  DFF_X1 key_c_r_reg_17_46 (.CK( clk ) , .D( key_c_r_16_46 ) , .Q( key_c_r_17_46 ) );
  DFF_X1 key_c_r_reg_17_47 (.CK( clk ) , .D( key_c_r_16_47 ) , .Q( key_c_r_17_47 ) );
  DFF_X1 key_c_r_reg_17_48 (.CK( clk ) , .D( key_c_r_16_48 ) , .Q( key_c_r_17_48 ) );
  DFF_X1 key_c_r_reg_17_49 (.CK( clk ) , .D( key_c_r_16_49 ) , .Q( key_c_r_17_49 ) );
  DFF_X1 key_c_r_reg_17_5 (.CK( clk ) , .D( key_c_r_16_5 ) , .Q( key_c_r_17_5 ) );
  DFF_X1 key_c_r_reg_17_50 (.CK( clk ) , .D( key_c_r_16_50 ) , .Q( key_c_r_17_50 ) );
  DFF_X1 key_c_r_reg_17_51 (.CK( clk ) , .D( key_c_r_16_51 ) , .Q( key_c_r_17_51 ) );
  DFF_X1 key_c_r_reg_17_52 (.CK( clk ) , .D( key_c_r_16_52 ) , .Q( key_c_r_17_52 ) );
  DFF_X1 key_c_r_reg_17_53 (.CK( clk ) , .D( key_c_r_16_53 ) , .Q( key_c_r_17_53 ) );
  DFF_X1 key_c_r_reg_17_54 (.CK( clk ) , .D( key_c_r_16_54 ) , .Q( key_c_r_17_54 ) );
  DFF_X1 key_c_r_reg_17_55 (.CK( clk ) , .D( key_c_r_16_55 ) , .Q( key_c_r_17_55 ) );
  DFF_X1 key_c_r_reg_17_6 (.CK( clk ) , .D( key_c_r_16_6 ) , .Q( key_c_r_17_6 ) );
  DFF_X1 key_c_r_reg_17_7 (.CK( clk ) , .D( key_c_r_16_7 ) , .Q( key_c_r_17_7 ) );
  DFF_X1 key_c_r_reg_17_8 (.CK( clk ) , .D( key_c_r_16_8 ) , .Q( key_c_r_17_8 ) );
  DFF_X1 key_c_r_reg_17_9 (.CK( clk ) , .D( key_c_r_16_9 ) , .Q( key_c_r_17_9 ) );
  DFF_X1 key_c_r_reg_18_0 (.CK( clk ) , .D( key_c_r_17_0 ) , .Q( key_c_r_18_0 ) );
  DFF_X1 key_c_r_reg_18_1 (.CK( clk ) , .D( key_c_r_17_1 ) , .Q( key_c_r_18_1 ) );
  DFF_X1 key_c_r_reg_18_10 (.CK( clk ) , .D( key_c_r_17_10 ) , .Q( key_c_r_18_10 ) );
  DFF_X1 key_c_r_reg_18_11 (.CK( clk ) , .D( key_c_r_17_11 ) , .Q( key_c_r_18_11 ) );
  DFF_X1 key_c_r_reg_18_12 (.CK( clk ) , .D( key_c_r_17_12 ) , .Q( key_c_r_18_12 ) );
  DFF_X1 key_c_r_reg_18_13 (.CK( clk ) , .D( key_c_r_17_13 ) , .Q( key_c_r_18_13 ) );
  DFF_X1 key_c_r_reg_18_14 (.CK( clk ) , .D( key_c_r_17_14 ) , .Q( key_c_r_18_14 ) );
  DFF_X1 key_c_r_reg_18_15 (.CK( clk ) , .D( key_c_r_17_15 ) , .Q( key_c_r_18_15 ) );
  DFF_X1 key_c_r_reg_18_16 (.CK( clk ) , .D( key_c_r_17_16 ) , .Q( key_c_r_18_16 ) );
  DFF_X1 key_c_r_reg_18_17 (.CK( clk ) , .D( key_c_r_17_17 ) , .Q( key_c_r_18_17 ) );
  DFF_X1 key_c_r_reg_18_18 (.CK( clk ) , .D( key_c_r_17_18 ) , .Q( key_c_r_18_18 ) );
  DFF_X1 key_c_r_reg_18_19 (.CK( clk ) , .D( key_c_r_17_19 ) , .Q( key_c_r_18_19 ) );
  DFF_X1 key_c_r_reg_18_2 (.CK( clk ) , .D( key_c_r_17_2 ) , .Q( key_c_r_18_2 ) );
  DFF_X1 key_c_r_reg_18_20 (.CK( clk ) , .D( key_c_r_17_20 ) , .Q( key_c_r_18_20 ) );
  DFF_X1 key_c_r_reg_18_21 (.CK( clk ) , .D( key_c_r_17_21 ) , .Q( key_c_r_18_21 ) );
  DFF_X1 key_c_r_reg_18_22 (.CK( clk ) , .D( key_c_r_17_22 ) , .Q( key_c_r_18_22 ) );
  DFF_X1 key_c_r_reg_18_23 (.CK( clk ) , .D( key_c_r_17_23 ) , .Q( key_c_r_18_23 ) );
  DFF_X1 key_c_r_reg_18_24 (.CK( clk ) , .D( key_c_r_17_24 ) , .Q( key_c_r_18_24 ) );
  DFF_X1 key_c_r_reg_18_25 (.CK( clk ) , .D( key_c_r_17_25 ) , .Q( key_c_r_18_25 ) );
  DFF_X1 key_c_r_reg_18_26 (.CK( clk ) , .D( key_c_r_17_26 ) , .Q( key_c_r_18_26 ) );
  DFF_X1 key_c_r_reg_18_27 (.CK( clk ) , .D( key_c_r_17_27 ) , .Q( key_c_r_18_27 ) );
  DFF_X1 key_c_r_reg_18_28 (.CK( clk ) , .D( key_c_r_17_28 ) , .Q( key_c_r_18_28 ) );
  DFF_X1 key_c_r_reg_18_29 (.CK( clk ) , .D( key_c_r_17_29 ) , .Q( key_c_r_18_29 ) );
  DFF_X1 key_c_r_reg_18_3 (.CK( clk ) , .D( key_c_r_17_3 ) , .Q( key_c_r_18_3 ) );
  DFF_X1 key_c_r_reg_18_30 (.CK( clk ) , .D( key_c_r_17_30 ) , .Q( key_c_r_18_30 ) );
  DFF_X1 key_c_r_reg_18_31 (.CK( clk ) , .D( key_c_r_17_31 ) , .Q( key_c_r_18_31 ) );
  DFF_X1 key_c_r_reg_18_32 (.CK( clk ) , .D( key_c_r_17_32 ) , .Q( key_c_r_18_32 ) );
  DFF_X1 key_c_r_reg_18_33 (.CK( clk ) , .D( key_c_r_17_33 ) , .Q( key_c_r_18_33 ) );
  DFF_X1 key_c_r_reg_18_34 (.CK( clk ) , .D( key_c_r_17_34 ) , .Q( key_c_r_18_34 ) );
  DFF_X1 key_c_r_reg_18_35 (.CK( clk ) , .D( key_c_r_17_35 ) , .Q( key_c_r_18_35 ) );
  DFF_X1 key_c_r_reg_18_36 (.CK( clk ) , .D( key_c_r_17_36 ) , .Q( key_c_r_18_36 ) );
  DFF_X1 key_c_r_reg_18_37 (.CK( clk ) , .D( key_c_r_17_37 ) , .Q( key_c_r_18_37 ) );
  DFF_X1 key_c_r_reg_18_38 (.CK( clk ) , .D( key_c_r_17_38 ) , .Q( key_c_r_18_38 ) );
  DFF_X1 key_c_r_reg_18_39 (.CK( clk ) , .D( key_c_r_17_39 ) , .Q( key_c_r_18_39 ) );
  DFF_X1 key_c_r_reg_18_4 (.CK( clk ) , .D( key_c_r_17_4 ) , .Q( key_c_r_18_4 ) );
  DFF_X1 key_c_r_reg_18_40 (.CK( clk ) , .D( key_c_r_17_40 ) , .Q( key_c_r_18_40 ) );
  DFF_X1 key_c_r_reg_18_41 (.CK( clk ) , .D( key_c_r_17_41 ) , .Q( key_c_r_18_41 ) );
  DFF_X1 key_c_r_reg_18_42 (.CK( clk ) , .D( key_c_r_17_42 ) , .Q( key_c_r_18_42 ) );
  DFF_X1 key_c_r_reg_18_43 (.CK( clk ) , .D( key_c_r_17_43 ) , .Q( key_c_r_18_43 ) );
  DFF_X1 key_c_r_reg_18_44 (.CK( clk ) , .D( key_c_r_17_44 ) , .Q( key_c_r_18_44 ) );
  DFF_X1 key_c_r_reg_18_45 (.CK( clk ) , .D( key_c_r_17_45 ) , .Q( key_c_r_18_45 ) );
  DFF_X1 key_c_r_reg_18_46 (.CK( clk ) , .D( key_c_r_17_46 ) , .Q( key_c_r_18_46 ) );
  DFF_X1 key_c_r_reg_18_47 (.CK( clk ) , .D( key_c_r_17_47 ) , .Q( key_c_r_18_47 ) );
  DFF_X1 key_c_r_reg_18_48 (.CK( clk ) , .D( key_c_r_17_48 ) , .Q( key_c_r_18_48 ) );
  DFF_X1 key_c_r_reg_18_49 (.CK( clk ) , .D( key_c_r_17_49 ) , .Q( key_c_r_18_49 ) );
  DFF_X1 key_c_r_reg_18_5 (.CK( clk ) , .D( key_c_r_17_5 ) , .Q( key_c_r_18_5 ) );
  DFF_X1 key_c_r_reg_18_50 (.CK( clk ) , .D( key_c_r_17_50 ) , .Q( key_c_r_18_50 ) );
  DFF_X1 key_c_r_reg_18_51 (.CK( clk ) , .D( key_c_r_17_51 ) , .Q( key_c_r_18_51 ) );
  DFF_X1 key_c_r_reg_18_52 (.CK( clk ) , .D( key_c_r_17_52 ) , .Q( key_c_r_18_52 ) );
  DFF_X1 key_c_r_reg_18_53 (.CK( clk ) , .D( key_c_r_17_53 ) , .Q( key_c_r_18_53 ) );
  DFF_X1 key_c_r_reg_18_54 (.CK( clk ) , .D( key_c_r_17_54 ) , .Q( key_c_r_18_54 ) );
  DFF_X1 key_c_r_reg_18_55 (.CK( clk ) , .D( key_c_r_17_55 ) , .Q( key_c_r_18_55 ) );
  DFF_X1 key_c_r_reg_18_6 (.CK( clk ) , .D( key_c_r_17_6 ) , .Q( key_c_r_18_6 ) );
  DFF_X1 key_c_r_reg_18_7 (.CK( clk ) , .D( key_c_r_17_7 ) , .Q( key_c_r_18_7 ) );
  DFF_X1 key_c_r_reg_18_8 (.CK( clk ) , .D( key_c_r_17_8 ) , .Q( key_c_r_18_8 ) );
  DFF_X1 key_c_r_reg_18_9 (.CK( clk ) , .D( key_c_r_17_9 ) , .Q( key_c_r_18_9 ) );
  DFF_X1 key_c_r_reg_19_0 (.CK( clk ) , .D( key_c_r_18_0 ) , .Q( key_c_r_19_0 ) );
  DFF_X1 key_c_r_reg_19_1 (.CK( clk ) , .D( key_c_r_18_1 ) , .Q( key_c_r_19_1 ) );
  DFF_X1 key_c_r_reg_19_10 (.CK( clk ) , .D( key_c_r_18_10 ) , .Q( key_c_r_19_10 ) );
  DFF_X1 key_c_r_reg_19_11 (.CK( clk ) , .D( key_c_r_18_11 ) , .Q( key_c_r_19_11 ) );
  DFF_X1 key_c_r_reg_19_12 (.CK( clk ) , .D( key_c_r_18_12 ) , .Q( key_c_r_19_12 ) );
  DFF_X1 key_c_r_reg_19_13 (.CK( clk ) , .D( key_c_r_18_13 ) , .Q( key_c_r_19_13 ) );
  DFF_X1 key_c_r_reg_19_14 (.CK( clk ) , .D( key_c_r_18_14 ) , .Q( key_c_r_19_14 ) );
  DFF_X1 key_c_r_reg_19_15 (.CK( clk ) , .D( key_c_r_18_15 ) , .Q( key_c_r_19_15 ) );
  DFF_X1 key_c_r_reg_19_16 (.CK( clk ) , .D( key_c_r_18_16 ) , .Q( key_c_r_19_16 ) );
  DFF_X1 key_c_r_reg_19_17 (.CK( clk ) , .D( key_c_r_18_17 ) , .Q( key_c_r_19_17 ) );
  DFF_X1 key_c_r_reg_19_18 (.CK( clk ) , .D( key_c_r_18_18 ) , .Q( key_c_r_19_18 ) );
  DFF_X1 key_c_r_reg_19_19 (.CK( clk ) , .D( key_c_r_18_19 ) , .Q( key_c_r_19_19 ) );
  DFF_X1 key_c_r_reg_19_2 (.CK( clk ) , .D( key_c_r_18_2 ) , .Q( key_c_r_19_2 ) );
  DFF_X1 key_c_r_reg_19_20 (.CK( clk ) , .D( key_c_r_18_20 ) , .Q( key_c_r_19_20 ) );
  DFF_X1 key_c_r_reg_19_21 (.CK( clk ) , .D( key_c_r_18_21 ) , .Q( key_c_r_19_21 ) );
  DFF_X1 key_c_r_reg_19_22 (.CK( clk ) , .D( key_c_r_18_22 ) , .Q( key_c_r_19_22 ) );
  DFF_X1 key_c_r_reg_19_23 (.CK( clk ) , .D( key_c_r_18_23 ) , .Q( key_c_r_19_23 ) );
  DFF_X1 key_c_r_reg_19_24 (.CK( clk ) , .D( key_c_r_18_24 ) , .Q( key_c_r_19_24 ) );
  DFF_X1 key_c_r_reg_19_25 (.CK( clk ) , .D( key_c_r_18_25 ) , .Q( key_c_r_19_25 ) );
  DFF_X1 key_c_r_reg_19_26 (.CK( clk ) , .D( key_c_r_18_26 ) , .Q( key_c_r_19_26 ) );
  DFF_X1 key_c_r_reg_19_27 (.CK( clk ) , .D( key_c_r_18_27 ) , .Q( key_c_r_19_27 ) );
  DFF_X1 key_c_r_reg_19_28 (.CK( clk ) , .D( key_c_r_18_28 ) , .Q( key_c_r_19_28 ) );
  DFF_X1 key_c_r_reg_19_29 (.CK( clk ) , .D( key_c_r_18_29 ) , .Q( key_c_r_19_29 ) );
  DFF_X1 key_c_r_reg_19_3 (.CK( clk ) , .D( key_c_r_18_3 ) , .Q( key_c_r_19_3 ) );
  DFF_X1 key_c_r_reg_19_30 (.CK( clk ) , .D( key_c_r_18_30 ) , .Q( key_c_r_19_30 ) );
  DFF_X1 key_c_r_reg_19_31 (.CK( clk ) , .D( key_c_r_18_31 ) , .Q( key_c_r_19_31 ) );
  DFF_X1 key_c_r_reg_19_32 (.CK( clk ) , .D( key_c_r_18_32 ) , .Q( key_c_r_19_32 ) );
  DFF_X1 key_c_r_reg_19_33 (.CK( clk ) , .D( key_c_r_18_33 ) , .Q( key_c_r_19_33 ) );
  DFF_X1 key_c_r_reg_19_34 (.CK( clk ) , .D( key_c_r_18_34 ) , .Q( key_c_r_19_34 ) );
  DFF_X1 key_c_r_reg_19_35 (.CK( clk ) , .D( key_c_r_18_35 ) , .Q( key_c_r_19_35 ) );
  DFF_X1 key_c_r_reg_19_36 (.CK( clk ) , .D( key_c_r_18_36 ) , .Q( key_c_r_19_36 ) );
  DFF_X1 key_c_r_reg_19_37 (.CK( clk ) , .D( key_c_r_18_37 ) , .Q( key_c_r_19_37 ) );
  DFF_X1 key_c_r_reg_19_38 (.CK( clk ) , .D( key_c_r_18_38 ) , .Q( key_c_r_19_38 ) );
  DFF_X1 key_c_r_reg_19_39 (.CK( clk ) , .D( key_c_r_18_39 ) , .Q( key_c_r_19_39 ) );
  DFF_X1 key_c_r_reg_19_4 (.CK( clk ) , .D( key_c_r_18_4 ) , .Q( key_c_r_19_4 ) );
  DFF_X1 key_c_r_reg_19_40 (.CK( clk ) , .D( key_c_r_18_40 ) , .Q( key_c_r_19_40 ) );
  DFF_X1 key_c_r_reg_19_41 (.CK( clk ) , .D( key_c_r_18_41 ) , .Q( key_c_r_19_41 ) );
  DFF_X1 key_c_r_reg_19_42 (.CK( clk ) , .D( key_c_r_18_42 ) , .Q( key_c_r_19_42 ) );
  DFF_X1 key_c_r_reg_19_43 (.CK( clk ) , .D( key_c_r_18_43 ) , .Q( key_c_r_19_43 ) );
  DFF_X1 key_c_r_reg_19_44 (.CK( clk ) , .D( key_c_r_18_44 ) , .Q( key_c_r_19_44 ) );
  DFF_X1 key_c_r_reg_19_45 (.CK( clk ) , .D( key_c_r_18_45 ) , .Q( key_c_r_19_45 ) );
  DFF_X1 key_c_r_reg_19_46 (.CK( clk ) , .D( key_c_r_18_46 ) , .Q( key_c_r_19_46 ) );
  DFF_X1 key_c_r_reg_19_47 (.CK( clk ) , .D( key_c_r_18_47 ) , .Q( key_c_r_19_47 ) );
  DFF_X1 key_c_r_reg_19_48 (.CK( clk ) , .D( key_c_r_18_48 ) , .Q( key_c_r_19_48 ) );
  DFF_X1 key_c_r_reg_19_49 (.CK( clk ) , .D( key_c_r_18_49 ) , .Q( key_c_r_19_49 ) );
  DFF_X1 key_c_r_reg_19_5 (.CK( clk ) , .D( key_c_r_18_5 ) , .Q( key_c_r_19_5 ) );
  DFF_X1 key_c_r_reg_19_50 (.CK( clk ) , .D( key_c_r_18_50 ) , .Q( key_c_r_19_50 ) );
  DFF_X1 key_c_r_reg_19_51 (.CK( clk ) , .D( key_c_r_18_51 ) , .Q( key_c_r_19_51 ) );
  DFF_X1 key_c_r_reg_19_52 (.CK( clk ) , .D( key_c_r_18_52 ) , .Q( key_c_r_19_52 ) );
  DFF_X1 key_c_r_reg_19_53 (.CK( clk ) , .D( key_c_r_18_53 ) , .Q( key_c_r_19_53 ) );
  DFF_X1 key_c_r_reg_19_54 (.CK( clk ) , .D( key_c_r_18_54 ) , .Q( key_c_r_19_54 ) );
  DFF_X1 key_c_r_reg_19_55 (.CK( clk ) , .D( key_c_r_18_55 ) , .Q( key_c_r_19_55 ) );
  DFF_X1 key_c_r_reg_19_6 (.CK( clk ) , .D( key_c_r_18_6 ) , .Q( key_c_r_19_6 ) );
  DFF_X1 key_c_r_reg_19_7 (.CK( clk ) , .D( key_c_r_18_7 ) , .Q( key_c_r_19_7 ) );
  DFF_X1 key_c_r_reg_19_8 (.CK( clk ) , .D( key_c_r_18_8 ) , .Q( key_c_r_19_8 ) );
  DFF_X1 key_c_r_reg_19_9 (.CK( clk ) , .D( key_c_r_18_9 ) , .Q( key_c_r_19_9 ) );
  DFF_X1 key_c_r_reg_1_0 (.CK( clk ) , .D( key_c_r_0_0 ) , .Q( key_c_r_1_0 ) );
  DFF_X1 key_c_r_reg_1_1 (.CK( clk ) , .D( key_c_r_0_1 ) , .Q( key_c_r_1_1 ) );
  DFF_X1 key_c_r_reg_1_10 (.CK( clk ) , .D( key_c_r_0_10 ) , .Q( key_c_r_1_10 ) );
  DFF_X1 key_c_r_reg_1_11 (.CK( clk ) , .D( key_c_r_0_11 ) , .Q( key_c_r_1_11 ) );
  DFF_X1 key_c_r_reg_1_12 (.CK( clk ) , .D( key_c_r_0_12 ) , .Q( key_c_r_1_12 ) );
  DFF_X1 key_c_r_reg_1_13 (.CK( clk ) , .D( key_c_r_0_13 ) , .Q( key_c_r_1_13 ) );
  DFF_X1 key_c_r_reg_1_14 (.CK( clk ) , .D( key_c_r_0_14 ) , .Q( key_c_r_1_14 ) );
  DFF_X1 key_c_r_reg_1_15 (.CK( clk ) , .D( key_c_r_0_15 ) , .Q( key_c_r_1_15 ) );
  DFF_X1 key_c_r_reg_1_16 (.CK( clk ) , .D( key_c_r_0_16 ) , .Q( key_c_r_1_16 ) );
  DFF_X1 key_c_r_reg_1_17 (.CK( clk ) , .D( key_c_r_0_17 ) , .Q( key_c_r_1_17 ) );
  DFF_X1 key_c_r_reg_1_18 (.CK( clk ) , .D( key_c_r_0_18 ) , .Q( key_c_r_1_18 ) );
  DFF_X1 key_c_r_reg_1_19 (.CK( clk ) , .D( key_c_r_0_19 ) , .Q( key_c_r_1_19 ) );
  DFF_X1 key_c_r_reg_1_2 (.CK( clk ) , .D( key_c_r_0_2 ) , .Q( key_c_r_1_2 ) );
  DFF_X1 key_c_r_reg_1_20 (.CK( clk ) , .D( key_c_r_0_20 ) , .Q( key_c_r_1_20 ) );
  DFF_X1 key_c_r_reg_1_21 (.CK( clk ) , .D( key_c_r_0_21 ) , .Q( key_c_r_1_21 ) );
  DFF_X1 key_c_r_reg_1_22 (.CK( clk ) , .D( key_c_r_0_22 ) , .Q( key_c_r_1_22 ) );
  DFF_X1 key_c_r_reg_1_23 (.CK( clk ) , .D( key_c_r_0_23 ) , .Q( key_c_r_1_23 ) );
  DFF_X1 key_c_r_reg_1_24 (.CK( clk ) , .D( key_c_r_0_24 ) , .Q( key_c_r_1_24 ) );
  DFF_X1 key_c_r_reg_1_25 (.CK( clk ) , .D( key_c_r_0_25 ) , .Q( key_c_r_1_25 ) );
  DFF_X1 key_c_r_reg_1_26 (.CK( clk ) , .D( key_c_r_0_26 ) , .Q( key_c_r_1_26 ) );
  DFF_X1 key_c_r_reg_1_27 (.CK( clk ) , .D( key_c_r_0_27 ) , .Q( key_c_r_1_27 ) );
  DFF_X1 key_c_r_reg_1_28 (.CK( clk ) , .D( key_c_r_0_28 ) , .Q( key_c_r_1_28 ) );
  DFF_X1 key_c_r_reg_1_29 (.CK( clk ) , .D( key_c_r_0_29 ) , .Q( key_c_r_1_29 ) );
  DFF_X1 key_c_r_reg_1_3 (.CK( clk ) , .D( key_c_r_0_3 ) , .Q( key_c_r_1_3 ) );
  DFF_X1 key_c_r_reg_1_30 (.CK( clk ) , .D( key_c_r_0_30 ) , .Q( key_c_r_1_30 ) );
  DFF_X1 key_c_r_reg_1_31 (.CK( clk ) , .D( key_c_r_0_31 ) , .Q( key_c_r_1_31 ) );
  DFF_X1 key_c_r_reg_1_32 (.CK( clk ) , .D( key_c_r_0_32 ) , .Q( key_c_r_1_32 ) );
  DFF_X1 key_c_r_reg_1_33 (.CK( clk ) , .D( key_c_r_0_33 ) , .Q( key_c_r_1_33 ) );
  DFF_X1 key_c_r_reg_1_34 (.CK( clk ) , .D( key_c_r_0_34 ) , .Q( key_c_r_1_34 ) );
  DFF_X1 key_c_r_reg_1_35 (.CK( clk ) , .D( key_c_r_0_35 ) , .Q( key_c_r_1_35 ) );
  DFF_X1 key_c_r_reg_1_36 (.CK( clk ) , .D( key_c_r_0_36 ) , .Q( key_c_r_1_36 ) );
  DFF_X1 key_c_r_reg_1_37 (.CK( clk ) , .D( key_c_r_0_37 ) , .Q( key_c_r_1_37 ) );
  DFF_X1 key_c_r_reg_1_38 (.CK( clk ) , .D( key_c_r_0_38 ) , .Q( key_c_r_1_38 ) );
  DFF_X1 key_c_r_reg_1_39 (.CK( clk ) , .D( key_c_r_0_39 ) , .Q( key_c_r_1_39 ) );
  DFF_X1 key_c_r_reg_1_4 (.CK( clk ) , .D( key_c_r_0_4 ) , .Q( key_c_r_1_4 ) );
  DFF_X1 key_c_r_reg_1_40 (.CK( clk ) , .D( key_c_r_0_40 ) , .Q( key_c_r_1_40 ) );
  DFF_X1 key_c_r_reg_1_41 (.CK( clk ) , .D( key_c_r_0_41 ) , .Q( key_c_r_1_41 ) );
  DFF_X1 key_c_r_reg_1_42 (.CK( clk ) , .D( key_c_r_0_42 ) , .Q( key_c_r_1_42 ) );
  DFF_X1 key_c_r_reg_1_43 (.CK( clk ) , .D( key_c_r_0_43 ) , .Q( key_c_r_1_43 ) );
  DFF_X1 key_c_r_reg_1_44 (.CK( clk ) , .D( key_c_r_0_44 ) , .Q( key_c_r_1_44 ) );
  DFF_X1 key_c_r_reg_1_45 (.CK( clk ) , .D( key_c_r_0_45 ) , .Q( key_c_r_1_45 ) );
  DFF_X1 key_c_r_reg_1_46 (.CK( clk ) , .D( key_c_r_0_46 ) , .Q( key_c_r_1_46 ) );
  DFF_X1 key_c_r_reg_1_47 (.CK( clk ) , .D( key_c_r_0_47 ) , .Q( key_c_r_1_47 ) );
  DFF_X1 key_c_r_reg_1_48 (.CK( clk ) , .D( key_c_r_0_48 ) , .Q( key_c_r_1_48 ) );
  DFF_X1 key_c_r_reg_1_49 (.CK( clk ) , .D( key_c_r_0_49 ) , .Q( key_c_r_1_49 ) );
  DFF_X1 key_c_r_reg_1_5 (.CK( clk ) , .D( key_c_r_0_5 ) , .Q( key_c_r_1_5 ) );
  DFF_X1 key_c_r_reg_1_50 (.CK( clk ) , .D( key_c_r_0_50 ) , .Q( key_c_r_1_50 ) );
  DFF_X1 key_c_r_reg_1_51 (.CK( clk ) , .D( key_c_r_0_51 ) , .Q( key_c_r_1_51 ) );
  DFF_X1 key_c_r_reg_1_52 (.CK( clk ) , .D( key_c_r_0_52 ) , .Q( key_c_r_1_52 ) );
  DFF_X1 key_c_r_reg_1_53 (.CK( clk ) , .D( key_c_r_0_53 ) , .Q( key_c_r_1_53 ) );
  DFF_X1 key_c_r_reg_1_54 (.CK( clk ) , .D( key_c_r_0_54 ) , .Q( key_c_r_1_54 ) );
  DFF_X1 key_c_r_reg_1_55 (.CK( clk ) , .D( key_c_r_0_55 ) , .Q( key_c_r_1_55 ) );
  DFF_X1 key_c_r_reg_1_6 (.CK( clk ) , .D( key_c_r_0_6 ) , .Q( key_c_r_1_6 ) );
  DFF_X1 key_c_r_reg_1_7 (.CK( clk ) , .D( key_c_r_0_7 ) , .Q( key_c_r_1_7 ) );
  DFF_X1 key_c_r_reg_1_8 (.CK( clk ) , .D( key_c_r_0_8 ) , .Q( key_c_r_1_8 ) );
  DFF_X1 key_c_r_reg_1_9 (.CK( clk ) , .D( key_c_r_0_9 ) , .Q( key_c_r_1_9 ) );
  DFF_X1 key_c_r_reg_20_0 (.CK( clk ) , .D( key_c_r_19_0 ) , .Q( key_c_r_20_0 ) );
  DFF_X1 key_c_r_reg_20_1 (.CK( clk ) , .D( key_c_r_19_1 ) , .Q( key_c_r_20_1 ) );
  DFF_X1 key_c_r_reg_20_10 (.CK( clk ) , .D( key_c_r_19_10 ) , .Q( key_c_r_20_10 ) );
  DFF_X1 key_c_r_reg_20_11 (.CK( clk ) , .D( key_c_r_19_11 ) , .Q( key_c_r_20_11 ) );
  DFF_X1 key_c_r_reg_20_12 (.CK( clk ) , .D( key_c_r_19_12 ) , .Q( key_c_r_20_12 ) );
  DFF_X1 key_c_r_reg_20_13 (.CK( clk ) , .D( key_c_r_19_13 ) , .Q( key_c_r_20_13 ) );
  DFF_X1 key_c_r_reg_20_14 (.CK( clk ) , .D( key_c_r_19_14 ) , .Q( key_c_r_20_14 ) );
  DFF_X1 key_c_r_reg_20_15 (.CK( clk ) , .D( key_c_r_19_15 ) , .Q( key_c_r_20_15 ) );
  DFF_X1 key_c_r_reg_20_16 (.CK( clk ) , .D( key_c_r_19_16 ) , .Q( key_c_r_20_16 ) );
  DFF_X1 key_c_r_reg_20_17 (.CK( clk ) , .D( key_c_r_19_17 ) , .Q( key_c_r_20_17 ) );
  DFF_X1 key_c_r_reg_20_18 (.CK( clk ) , .D( key_c_r_19_18 ) , .Q( key_c_r_20_18 ) );
  DFF_X1 key_c_r_reg_20_19 (.CK( clk ) , .D( key_c_r_19_19 ) , .Q( key_c_r_20_19 ) );
  DFF_X1 key_c_r_reg_20_2 (.CK( clk ) , .D( key_c_r_19_2 ) , .Q( key_c_r_20_2 ) );
  DFF_X1 key_c_r_reg_20_20 (.CK( clk ) , .D( key_c_r_19_20 ) , .Q( key_c_r_20_20 ) );
  DFF_X1 key_c_r_reg_20_21 (.CK( clk ) , .D( key_c_r_19_21 ) , .Q( key_c_r_20_21 ) );
  DFF_X1 key_c_r_reg_20_22 (.CK( clk ) , .D( key_c_r_19_22 ) , .Q( key_c_r_20_22 ) );
  DFF_X1 key_c_r_reg_20_23 (.CK( clk ) , .D( key_c_r_19_23 ) , .Q( key_c_r_20_23 ) );
  DFF_X1 key_c_r_reg_20_24 (.CK( clk ) , .D( key_c_r_19_24 ) , .Q( key_c_r_20_24 ) );
  DFF_X1 key_c_r_reg_20_25 (.CK( clk ) , .D( key_c_r_19_25 ) , .Q( key_c_r_20_25 ) );
  DFF_X1 key_c_r_reg_20_26 (.CK( clk ) , .D( key_c_r_19_26 ) , .Q( key_c_r_20_26 ) );
  DFF_X1 key_c_r_reg_20_27 (.CK( clk ) , .D( key_c_r_19_27 ) , .Q( key_c_r_20_27 ) );
  DFF_X1 key_c_r_reg_20_28 (.CK( clk ) , .D( key_c_r_19_28 ) , .Q( key_c_r_20_28 ) );
  DFF_X1 key_c_r_reg_20_29 (.CK( clk ) , .D( key_c_r_19_29 ) , .Q( key_c_r_20_29 ) );
  DFF_X1 key_c_r_reg_20_3 (.CK( clk ) , .D( key_c_r_19_3 ) , .Q( key_c_r_20_3 ) );
  DFF_X1 key_c_r_reg_20_30 (.CK( clk ) , .D( key_c_r_19_30 ) , .Q( key_c_r_20_30 ) );
  DFF_X1 key_c_r_reg_20_31 (.CK( clk ) , .D( key_c_r_19_31 ) , .Q( key_c_r_20_31 ) );
  DFF_X1 key_c_r_reg_20_32 (.CK( clk ) , .D( key_c_r_19_32 ) , .Q( key_c_r_20_32 ) );
  DFF_X1 key_c_r_reg_20_33 (.CK( clk ) , .D( key_c_r_19_33 ) , .Q( key_c_r_20_33 ) );
  DFF_X1 key_c_r_reg_20_34 (.CK( clk ) , .D( key_c_r_19_34 ) , .Q( key_c_r_20_34 ) );
  DFF_X1 key_c_r_reg_20_35 (.CK( clk ) , .D( key_c_r_19_35 ) , .Q( key_c_r_20_35 ) );
  DFF_X1 key_c_r_reg_20_36 (.CK( clk ) , .D( key_c_r_19_36 ) , .Q( key_c_r_20_36 ) );
  DFF_X1 key_c_r_reg_20_37 (.CK( clk ) , .D( key_c_r_19_37 ) , .Q( key_c_r_20_37 ) );
  DFF_X1 key_c_r_reg_20_38 (.CK( clk ) , .D( key_c_r_19_38 ) , .Q( key_c_r_20_38 ) );
  DFF_X1 key_c_r_reg_20_39 (.CK( clk ) , .D( key_c_r_19_39 ) , .Q( key_c_r_20_39 ) );
  DFF_X1 key_c_r_reg_20_4 (.CK( clk ) , .D( key_c_r_19_4 ) , .Q( key_c_r_20_4 ) );
  DFF_X1 key_c_r_reg_20_40 (.CK( clk ) , .D( key_c_r_19_40 ) , .Q( key_c_r_20_40 ) );
  DFF_X1 key_c_r_reg_20_41 (.CK( clk ) , .D( key_c_r_19_41 ) , .Q( key_c_r_20_41 ) );
  DFF_X1 key_c_r_reg_20_42 (.CK( clk ) , .D( key_c_r_19_42 ) , .Q( key_c_r_20_42 ) );
  DFF_X1 key_c_r_reg_20_43 (.CK( clk ) , .D( key_c_r_19_43 ) , .Q( key_c_r_20_43 ) );
  DFF_X1 key_c_r_reg_20_44 (.CK( clk ) , .D( key_c_r_19_44 ) , .Q( key_c_r_20_44 ) );
  DFF_X1 key_c_r_reg_20_45 (.CK( clk ) , .D( key_c_r_19_45 ) , .Q( key_c_r_20_45 ) );
  DFF_X1 key_c_r_reg_20_46 (.CK( clk ) , .D( key_c_r_19_46 ) , .Q( key_c_r_20_46 ) );
  DFF_X1 key_c_r_reg_20_47 (.CK( clk ) , .D( key_c_r_19_47 ) , .Q( key_c_r_20_47 ) );
  DFF_X1 key_c_r_reg_20_48 (.CK( clk ) , .D( key_c_r_19_48 ) , .Q( key_c_r_20_48 ) );
  DFF_X1 key_c_r_reg_20_49 (.CK( clk ) , .D( key_c_r_19_49 ) , .Q( key_c_r_20_49 ) );
  DFF_X1 key_c_r_reg_20_5 (.CK( clk ) , .D( key_c_r_19_5 ) , .Q( key_c_r_20_5 ) );
  DFF_X1 key_c_r_reg_20_50 (.CK( clk ) , .D( key_c_r_19_50 ) , .Q( key_c_r_20_50 ) );
  DFF_X1 key_c_r_reg_20_51 (.CK( clk ) , .D( key_c_r_19_51 ) , .Q( key_c_r_20_51 ) );
  DFF_X1 key_c_r_reg_20_52 (.CK( clk ) , .D( key_c_r_19_52 ) , .Q( key_c_r_20_52 ) );
  DFF_X1 key_c_r_reg_20_53 (.CK( clk ) , .D( key_c_r_19_53 ) , .Q( key_c_r_20_53 ) );
  DFF_X1 key_c_r_reg_20_54 (.CK( clk ) , .D( key_c_r_19_54 ) , .Q( key_c_r_20_54 ) );
  DFF_X1 key_c_r_reg_20_55 (.CK( clk ) , .D( key_c_r_19_55 ) , .Q( key_c_r_20_55 ) );
  DFF_X1 key_c_r_reg_20_6 (.CK( clk ) , .D( key_c_r_19_6 ) , .Q( key_c_r_20_6 ) );
  DFF_X1 key_c_r_reg_20_7 (.CK( clk ) , .D( key_c_r_19_7 ) , .Q( key_c_r_20_7 ) );
  DFF_X1 key_c_r_reg_20_8 (.CK( clk ) , .D( key_c_r_19_8 ) , .Q( key_c_r_20_8 ) );
  DFF_X1 key_c_r_reg_20_9 (.CK( clk ) , .D( key_c_r_19_9 ) , .Q( key_c_r_20_9 ) );
  DFF_X1 key_c_r_reg_21_0 (.CK( clk ) , .D( key_c_r_20_0 ) , .Q( key_c_r_21_0 ) );
  DFF_X1 key_c_r_reg_21_1 (.CK( clk ) , .D( key_c_r_20_1 ) , .Q( key_c_r_21_1 ) );
  DFF_X1 key_c_r_reg_21_10 (.CK( clk ) , .D( key_c_r_20_10 ) , .Q( key_c_r_21_10 ) );
  DFF_X1 key_c_r_reg_21_11 (.CK( clk ) , .D( key_c_r_20_11 ) , .Q( key_c_r_21_11 ) );
  DFF_X1 key_c_r_reg_21_12 (.CK( clk ) , .D( key_c_r_20_12 ) , .Q( key_c_r_21_12 ) );
  DFF_X1 key_c_r_reg_21_13 (.CK( clk ) , .D( key_c_r_20_13 ) , .Q( key_c_r_21_13 ) );
  DFF_X1 key_c_r_reg_21_14 (.CK( clk ) , .D( key_c_r_20_14 ) , .Q( key_c_r_21_14 ) );
  DFF_X1 key_c_r_reg_21_15 (.CK( clk ) , .D( key_c_r_20_15 ) , .Q( key_c_r_21_15 ) );
  DFF_X1 key_c_r_reg_21_16 (.CK( clk ) , .D( key_c_r_20_16 ) , .Q( key_c_r_21_16 ) );
  DFF_X1 key_c_r_reg_21_17 (.CK( clk ) , .D( key_c_r_20_17 ) , .Q( key_c_r_21_17 ) );
  DFF_X1 key_c_r_reg_21_18 (.CK( clk ) , .D( key_c_r_20_18 ) , .Q( key_c_r_21_18 ) );
  DFF_X1 key_c_r_reg_21_19 (.CK( clk ) , .D( key_c_r_20_19 ) , .Q( key_c_r_21_19 ) );
  DFF_X1 key_c_r_reg_21_2 (.CK( clk ) , .D( key_c_r_20_2 ) , .Q( key_c_r_21_2 ) );
  DFF_X1 key_c_r_reg_21_20 (.CK( clk ) , .D( key_c_r_20_20 ) , .Q( key_c_r_21_20 ) );
  DFF_X1 key_c_r_reg_21_21 (.CK( clk ) , .D( key_c_r_20_21 ) , .Q( key_c_r_21_21 ) );
  DFF_X1 key_c_r_reg_21_22 (.CK( clk ) , .D( key_c_r_20_22 ) , .Q( key_c_r_21_22 ) );
  DFF_X1 key_c_r_reg_21_23 (.CK( clk ) , .D( key_c_r_20_23 ) , .Q( key_c_r_21_23 ) );
  DFF_X1 key_c_r_reg_21_24 (.CK( clk ) , .D( key_c_r_20_24 ) , .Q( key_c_r_21_24 ) );
  DFF_X1 key_c_r_reg_21_25 (.CK( clk ) , .D( key_c_r_20_25 ) , .Q( key_c_r_21_25 ) );
  DFF_X1 key_c_r_reg_21_26 (.CK( clk ) , .D( key_c_r_20_26 ) , .Q( key_c_r_21_26 ) );
  DFF_X1 key_c_r_reg_21_27 (.CK( clk ) , .D( key_c_r_20_27 ) , .Q( key_c_r_21_27 ) );
  DFF_X1 key_c_r_reg_21_28 (.CK( clk ) , .D( key_c_r_20_28 ) , .Q( key_c_r_21_28 ) );
  DFF_X1 key_c_r_reg_21_29 (.CK( clk ) , .D( key_c_r_20_29 ) , .Q( key_c_r_21_29 ) );
  DFF_X1 key_c_r_reg_21_3 (.CK( clk ) , .D( key_c_r_20_3 ) , .Q( key_c_r_21_3 ) );
  DFF_X1 key_c_r_reg_21_30 (.CK( clk ) , .D( key_c_r_20_30 ) , .Q( key_c_r_21_30 ) );
  DFF_X1 key_c_r_reg_21_31 (.CK( clk ) , .D( key_c_r_20_31 ) , .Q( key_c_r_21_31 ) );
  DFF_X1 key_c_r_reg_21_32 (.CK( clk ) , .D( key_c_r_20_32 ) , .Q( key_c_r_21_32 ) );
  DFF_X1 key_c_r_reg_21_33 (.CK( clk ) , .D( key_c_r_20_33 ) , .Q( key_c_r_21_33 ) );
  DFF_X1 key_c_r_reg_21_34 (.CK( clk ) , .D( key_c_r_20_34 ) , .Q( key_c_r_21_34 ) );
  DFF_X1 key_c_r_reg_21_35 (.CK( clk ) , .D( key_c_r_20_35 ) , .Q( key_c_r_21_35 ) );
  DFF_X1 key_c_r_reg_21_36 (.CK( clk ) , .D( key_c_r_20_36 ) , .Q( key_c_r_21_36 ) );
  DFF_X1 key_c_r_reg_21_37 (.CK( clk ) , .D( key_c_r_20_37 ) , .Q( key_c_r_21_37 ) );
  DFF_X1 key_c_r_reg_21_38 (.CK( clk ) , .D( key_c_r_20_38 ) , .Q( key_c_r_21_38 ) );
  DFF_X1 key_c_r_reg_21_39 (.CK( clk ) , .D( key_c_r_20_39 ) , .Q( key_c_r_21_39 ) );
  DFF_X1 key_c_r_reg_21_4 (.CK( clk ) , .D( key_c_r_20_4 ) , .Q( key_c_r_21_4 ) );
  DFF_X1 key_c_r_reg_21_40 (.CK( clk ) , .D( key_c_r_20_40 ) , .Q( key_c_r_21_40 ) );
  DFF_X1 key_c_r_reg_21_41 (.CK( clk ) , .D( key_c_r_20_41 ) , .Q( key_c_r_21_41 ) );
  DFF_X1 key_c_r_reg_21_42 (.CK( clk ) , .D( key_c_r_20_42 ) , .Q( key_c_r_21_42 ) );
  DFF_X1 key_c_r_reg_21_43 (.CK( clk ) , .D( key_c_r_20_43 ) , .Q( key_c_r_21_43 ) );
  DFF_X1 key_c_r_reg_21_44 (.CK( clk ) , .D( key_c_r_20_44 ) , .Q( key_c_r_21_44 ) );
  DFF_X1 key_c_r_reg_21_45 (.CK( clk ) , .D( key_c_r_20_45 ) , .Q( key_c_r_21_45 ) );
  DFF_X1 key_c_r_reg_21_46 (.CK( clk ) , .D( key_c_r_20_46 ) , .Q( key_c_r_21_46 ) );
  DFF_X1 key_c_r_reg_21_47 (.CK( clk ) , .D( key_c_r_20_47 ) , .Q( key_c_r_21_47 ) );
  DFF_X1 key_c_r_reg_21_48 (.CK( clk ) , .D( key_c_r_20_48 ) , .Q( key_c_r_21_48 ) );
  DFF_X1 key_c_r_reg_21_49 (.CK( clk ) , .D( key_c_r_20_49 ) , .Q( key_c_r_21_49 ) );
  DFF_X1 key_c_r_reg_21_5 (.CK( clk ) , .D( key_c_r_20_5 ) , .Q( key_c_r_21_5 ) );
  DFF_X1 key_c_r_reg_21_50 (.CK( clk ) , .D( key_c_r_20_50 ) , .Q( key_c_r_21_50 ) );
  DFF_X1 key_c_r_reg_21_51 (.CK( clk ) , .D( key_c_r_20_51 ) , .Q( key_c_r_21_51 ) );
  DFF_X1 key_c_r_reg_21_52 (.CK( clk ) , .D( key_c_r_20_52 ) , .Q( key_c_r_21_52 ) );
  DFF_X1 key_c_r_reg_21_53 (.CK( clk ) , .D( key_c_r_20_53 ) , .Q( key_c_r_21_53 ) );
  DFF_X1 key_c_r_reg_21_54 (.CK( clk ) , .D( key_c_r_20_54 ) , .Q( key_c_r_21_54 ) );
  DFF_X1 key_c_r_reg_21_55 (.CK( clk ) , .D( key_c_r_20_55 ) , .Q( key_c_r_21_55 ) );
  DFF_X1 key_c_r_reg_21_6 (.CK( clk ) , .D( key_c_r_20_6 ) , .Q( key_c_r_21_6 ) );
  DFF_X1 key_c_r_reg_21_7 (.CK( clk ) , .D( key_c_r_20_7 ) , .Q( key_c_r_21_7 ) );
  DFF_X1 key_c_r_reg_21_8 (.CK( clk ) , .D( key_c_r_20_8 ) , .Q( key_c_r_21_8 ) );
  DFF_X1 key_c_r_reg_21_9 (.CK( clk ) , .D( key_c_r_20_9 ) , .Q( key_c_r_21_9 ) );
  DFF_X1 key_c_r_reg_22_0 (.CK( clk ) , .D( key_c_r_21_0 ) , .Q( key_c_r_22_0 ) );
  DFF_X1 key_c_r_reg_22_1 (.CK( clk ) , .D( key_c_r_21_1 ) , .Q( key_c_r_22_1 ) );
  DFF_X1 key_c_r_reg_22_10 (.CK( clk ) , .D( key_c_r_21_10 ) , .Q( key_c_r_22_10 ) );
  DFF_X1 key_c_r_reg_22_11 (.CK( clk ) , .D( key_c_r_21_11 ) , .Q( key_c_r_22_11 ) );
  DFF_X1 key_c_r_reg_22_12 (.CK( clk ) , .D( key_c_r_21_12 ) , .Q( key_c_r_22_12 ) );
  DFF_X1 key_c_r_reg_22_13 (.CK( clk ) , .D( key_c_r_21_13 ) , .Q( key_c_r_22_13 ) );
  DFF_X1 key_c_r_reg_22_14 (.CK( clk ) , .D( key_c_r_21_14 ) , .Q( key_c_r_22_14 ) );
  DFF_X1 key_c_r_reg_22_15 (.CK( clk ) , .D( key_c_r_21_15 ) , .Q( key_c_r_22_15 ) );
  DFF_X1 key_c_r_reg_22_16 (.CK( clk ) , .D( key_c_r_21_16 ) , .Q( key_c_r_22_16 ) );
  DFF_X1 key_c_r_reg_22_17 (.CK( clk ) , .D( key_c_r_21_17 ) , .Q( key_c_r_22_17 ) );
  DFF_X1 key_c_r_reg_22_18 (.CK( clk ) , .D( key_c_r_21_18 ) , .Q( key_c_r_22_18 ) );
  DFF_X1 key_c_r_reg_22_19 (.CK( clk ) , .D( key_c_r_21_19 ) , .Q( key_c_r_22_19 ) );
  DFF_X1 key_c_r_reg_22_2 (.CK( clk ) , .D( key_c_r_21_2 ) , .Q( key_c_r_22_2 ) );
  DFF_X1 key_c_r_reg_22_20 (.CK( clk ) , .D( key_c_r_21_20 ) , .Q( key_c_r_22_20 ) );
  DFF_X1 key_c_r_reg_22_21 (.CK( clk ) , .D( key_c_r_21_21 ) , .Q( key_c_r_22_21 ) );
  DFF_X1 key_c_r_reg_22_22 (.CK( clk ) , .D( key_c_r_21_22 ) , .Q( key_c_r_22_22 ) );
  DFF_X1 key_c_r_reg_22_23 (.CK( clk ) , .D( key_c_r_21_23 ) , .Q( key_c_r_22_23 ) );
  DFF_X1 key_c_r_reg_22_24 (.CK( clk ) , .D( key_c_r_21_24 ) , .Q( key_c_r_22_24 ) );
  DFF_X1 key_c_r_reg_22_25 (.CK( clk ) , .D( key_c_r_21_25 ) , .Q( key_c_r_22_25 ) );
  DFF_X1 key_c_r_reg_22_26 (.CK( clk ) , .D( key_c_r_21_26 ) , .Q( key_c_r_22_26 ) );
  DFF_X1 key_c_r_reg_22_27 (.CK( clk ) , .D( key_c_r_21_27 ) , .Q( key_c_r_22_27 ) );
  DFF_X1 key_c_r_reg_22_28 (.CK( clk ) , .D( key_c_r_21_28 ) , .Q( key_c_r_22_28 ) );
  DFF_X1 key_c_r_reg_22_29 (.CK( clk ) , .D( key_c_r_21_29 ) , .Q( key_c_r_22_29 ) );
  DFF_X1 key_c_r_reg_22_3 (.CK( clk ) , .D( key_c_r_21_3 ) , .Q( key_c_r_22_3 ) );
  DFF_X1 key_c_r_reg_22_30 (.CK( clk ) , .D( key_c_r_21_30 ) , .Q( key_c_r_22_30 ) );
  DFF_X1 key_c_r_reg_22_31 (.CK( clk ) , .D( key_c_r_21_31 ) , .Q( key_c_r_22_31 ) );
  DFF_X1 key_c_r_reg_22_32 (.CK( clk ) , .D( key_c_r_21_32 ) , .Q( key_c_r_22_32 ) );
  DFF_X1 key_c_r_reg_22_33 (.CK( clk ) , .D( key_c_r_21_33 ) , .Q( key_c_r_22_33 ) );
  DFF_X1 key_c_r_reg_22_34 (.CK( clk ) , .D( key_c_r_21_34 ) , .Q( key_c_r_22_34 ) );
  DFF_X1 key_c_r_reg_22_35 (.CK( clk ) , .D( key_c_r_21_35 ) , .Q( key_c_r_22_35 ) );
  DFF_X1 key_c_r_reg_22_36 (.CK( clk ) , .D( key_c_r_21_36 ) , .Q( key_c_r_22_36 ) );
  DFF_X1 key_c_r_reg_22_37 (.CK( clk ) , .D( key_c_r_21_37 ) , .Q( key_c_r_22_37 ) );
  DFF_X1 key_c_r_reg_22_38 (.CK( clk ) , .D( key_c_r_21_38 ) , .Q( key_c_r_22_38 ) );
  DFF_X1 key_c_r_reg_22_39 (.CK( clk ) , .D( key_c_r_21_39 ) , .Q( key_c_r_22_39 ) );
  DFF_X1 key_c_r_reg_22_4 (.CK( clk ) , .D( key_c_r_21_4 ) , .Q( key_c_r_22_4 ) );
  DFF_X1 key_c_r_reg_22_40 (.CK( clk ) , .D( key_c_r_21_40 ) , .Q( key_c_r_22_40 ) );
  DFF_X1 key_c_r_reg_22_41 (.CK( clk ) , .D( key_c_r_21_41 ) , .Q( key_c_r_22_41 ) );
  DFF_X1 key_c_r_reg_22_42 (.CK( clk ) , .D( key_c_r_21_42 ) , .Q( key_c_r_22_42 ) );
  DFF_X1 key_c_r_reg_22_43 (.CK( clk ) , .D( key_c_r_21_43 ) , .Q( key_c_r_22_43 ) );
  DFF_X1 key_c_r_reg_22_44 (.CK( clk ) , .D( key_c_r_21_44 ) , .Q( key_c_r_22_44 ) );
  DFF_X1 key_c_r_reg_22_45 (.CK( clk ) , .D( key_c_r_21_45 ) , .Q( key_c_r_22_45 ) );
  DFF_X1 key_c_r_reg_22_46 (.CK( clk ) , .D( key_c_r_21_46 ) , .Q( key_c_r_22_46 ) );
  DFF_X1 key_c_r_reg_22_47 (.CK( clk ) , .D( key_c_r_21_47 ) , .Q( key_c_r_22_47 ) );
  DFF_X1 key_c_r_reg_22_48 (.CK( clk ) , .D( key_c_r_21_48 ) , .Q( key_c_r_22_48 ) );
  DFF_X1 key_c_r_reg_22_49 (.CK( clk ) , .D( key_c_r_21_49 ) , .Q( key_c_r_22_49 ) );
  DFF_X1 key_c_r_reg_22_5 (.CK( clk ) , .D( key_c_r_21_5 ) , .Q( key_c_r_22_5 ) );
  DFF_X1 key_c_r_reg_22_50 (.CK( clk ) , .D( key_c_r_21_50 ) , .Q( key_c_r_22_50 ) );
  DFF_X1 key_c_r_reg_22_51 (.CK( clk ) , .D( key_c_r_21_51 ) , .Q( key_c_r_22_51 ) );
  DFF_X1 key_c_r_reg_22_52 (.CK( clk ) , .D( key_c_r_21_52 ) , .Q( key_c_r_22_52 ) );
  DFF_X1 key_c_r_reg_22_53 (.CK( clk ) , .D( key_c_r_21_53 ) , .Q( key_c_r_22_53 ) );
  DFF_X1 key_c_r_reg_22_54 (.CK( clk ) , .D( key_c_r_21_54 ) , .Q( key_c_r_22_54 ) );
  DFF_X1 key_c_r_reg_22_55 (.CK( clk ) , .D( key_c_r_21_55 ) , .Q( key_c_r_22_55 ) );
  DFF_X1 key_c_r_reg_22_6 (.CK( clk ) , .D( key_c_r_21_6 ) , .Q( key_c_r_22_6 ) );
  DFF_X1 key_c_r_reg_22_7 (.CK( clk ) , .D( key_c_r_21_7 ) , .Q( key_c_r_22_7 ) );
  DFF_X1 key_c_r_reg_22_8 (.CK( clk ) , .D( key_c_r_21_8 ) , .Q( key_c_r_22_8 ) );
  DFF_X1 key_c_r_reg_22_9 (.CK( clk ) , .D( key_c_r_21_9 ) , .Q( key_c_r_22_9 ) );
  DFF_X1 key_c_r_reg_23_0 (.CK( clk ) , .D( key_c_r_22_0 ) , .Q( key_c_r_23_0 ) );
  DFF_X1 key_c_r_reg_23_1 (.CK( clk ) , .D( key_c_r_22_1 ) , .Q( key_c_r_23_1 ) );
  DFF_X1 key_c_r_reg_23_10 (.CK( clk ) , .D( key_c_r_22_10 ) , .Q( key_c_r_23_10 ) );
  DFF_X1 key_c_r_reg_23_11 (.CK( clk ) , .D( key_c_r_22_11 ) , .Q( key_c_r_23_11 ) );
  DFF_X1 key_c_r_reg_23_12 (.CK( clk ) , .D( key_c_r_22_12 ) , .Q( key_c_r_23_12 ) );
  DFF_X1 key_c_r_reg_23_13 (.CK( clk ) , .D( key_c_r_22_13 ) , .Q( key_c_r_23_13 ) );
  DFF_X1 key_c_r_reg_23_14 (.CK( clk ) , .D( key_c_r_22_14 ) , .Q( key_c_r_23_14 ) );
  DFF_X1 key_c_r_reg_23_15 (.CK( clk ) , .D( key_c_r_22_15 ) , .Q( key_c_r_23_15 ) );
  DFF_X1 key_c_r_reg_23_16 (.CK( clk ) , .D( key_c_r_22_16 ) , .Q( key_c_r_23_16 ) );
  DFF_X1 key_c_r_reg_23_17 (.CK( clk ) , .D( key_c_r_22_17 ) , .Q( key_c_r_23_17 ) );
  DFF_X1 key_c_r_reg_23_18 (.CK( clk ) , .D( key_c_r_22_18 ) , .Q( key_c_r_23_18 ) );
  DFF_X1 key_c_r_reg_23_19 (.CK( clk ) , .D( key_c_r_22_19 ) , .Q( key_c_r_23_19 ) );
  DFF_X1 key_c_r_reg_23_2 (.CK( clk ) , .D( key_c_r_22_2 ) , .Q( key_c_r_23_2 ) );
  DFF_X1 key_c_r_reg_23_20 (.CK( clk ) , .D( key_c_r_22_20 ) , .Q( key_c_r_23_20 ) );
  DFF_X1 key_c_r_reg_23_21 (.CK( clk ) , .D( key_c_r_22_21 ) , .Q( key_c_r_23_21 ) );
  DFF_X1 key_c_r_reg_23_22 (.CK( clk ) , .D( key_c_r_22_22 ) , .Q( key_c_r_23_22 ) );
  DFF_X1 key_c_r_reg_23_23 (.CK( clk ) , .D( key_c_r_22_23 ) , .Q( key_c_r_23_23 ) );
  DFF_X1 key_c_r_reg_23_24 (.CK( clk ) , .D( key_c_r_22_24 ) , .Q( key_c_r_23_24 ) );
  DFF_X1 key_c_r_reg_23_25 (.CK( clk ) , .D( key_c_r_22_25 ) , .Q( key_c_r_23_25 ) );
  DFF_X1 key_c_r_reg_23_26 (.CK( clk ) , .D( key_c_r_22_26 ) , .Q( key_c_r_23_26 ) );
  DFF_X1 key_c_r_reg_23_27 (.CK( clk ) , .D( key_c_r_22_27 ) , .Q( key_c_r_23_27 ) );
  DFF_X1 key_c_r_reg_23_28 (.CK( clk ) , .D( key_c_r_22_28 ) , .Q( key_c_r_23_28 ) );
  DFF_X1 key_c_r_reg_23_29 (.CK( clk ) , .D( key_c_r_22_29 ) , .Q( key_c_r_23_29 ) );
  DFF_X1 key_c_r_reg_23_3 (.CK( clk ) , .D( key_c_r_22_3 ) , .Q( key_c_r_23_3 ) );
  DFF_X1 key_c_r_reg_23_30 (.CK( clk ) , .D( key_c_r_22_30 ) , .Q( key_c_r_23_30 ) );
  DFF_X1 key_c_r_reg_23_31 (.CK( clk ) , .D( key_c_r_22_31 ) , .Q( key_c_r_23_31 ) );
  DFF_X1 key_c_r_reg_23_32 (.CK( clk ) , .D( key_c_r_22_32 ) , .Q( key_c_r_23_32 ) );
  DFF_X1 key_c_r_reg_23_33 (.CK( clk ) , .D( key_c_r_22_33 ) , .Q( key_c_r_23_33 ) );
  DFF_X1 key_c_r_reg_23_34 (.CK( clk ) , .D( key_c_r_22_34 ) , .Q( key_c_r_23_34 ) );
  DFF_X1 key_c_r_reg_23_35 (.CK( clk ) , .D( key_c_r_22_35 ) , .Q( key_c_r_23_35 ) );
  DFF_X1 key_c_r_reg_23_36 (.CK( clk ) , .D( key_c_r_22_36 ) , .Q( key_c_r_23_36 ) );
  DFF_X1 key_c_r_reg_23_37 (.CK( clk ) , .D( key_c_r_22_37 ) , .Q( key_c_r_23_37 ) );
  DFF_X1 key_c_r_reg_23_38 (.CK( clk ) , .D( key_c_r_22_38 ) , .Q( key_c_r_23_38 ) );
  DFF_X1 key_c_r_reg_23_39 (.CK( clk ) , .D( key_c_r_22_39 ) , .Q( key_c_r_23_39 ) );
  DFF_X1 key_c_r_reg_23_4 (.CK( clk ) , .D( key_c_r_22_4 ) , .Q( key_c_r_23_4 ) );
  DFF_X1 key_c_r_reg_23_40 (.CK( clk ) , .D( key_c_r_22_40 ) , .Q( key_c_r_23_40 ) );
  DFF_X1 key_c_r_reg_23_41 (.CK( clk ) , .D( key_c_r_22_41 ) , .Q( key_c_r_23_41 ) );
  DFF_X1 key_c_r_reg_23_42 (.CK( clk ) , .D( key_c_r_22_42 ) , .Q( key_c_r_23_42 ) );
  DFF_X1 key_c_r_reg_23_43 (.CK( clk ) , .D( key_c_r_22_43 ) , .Q( key_c_r_23_43 ) );
  DFF_X1 key_c_r_reg_23_44 (.CK( clk ) , .D( key_c_r_22_44 ) , .Q( key_c_r_23_44 ) );
  DFF_X1 key_c_r_reg_23_45 (.CK( clk ) , .D( key_c_r_22_45 ) , .Q( key_c_r_23_45 ) );
  DFF_X1 key_c_r_reg_23_46 (.CK( clk ) , .D( key_c_r_22_46 ) , .Q( key_c_r_23_46 ) );
  DFF_X1 key_c_r_reg_23_47 (.CK( clk ) , .D( key_c_r_22_47 ) , .Q( key_c_r_23_47 ) );
  DFF_X1 key_c_r_reg_23_48 (.CK( clk ) , .D( key_c_r_22_48 ) , .Q( key_c_r_23_48 ) );
  DFF_X1 key_c_r_reg_23_49 (.CK( clk ) , .D( key_c_r_22_49 ) , .Q( key_c_r_23_49 ) );
  DFF_X1 key_c_r_reg_23_5 (.CK( clk ) , .D( key_c_r_22_5 ) , .Q( key_c_r_23_5 ) );
  DFF_X1 key_c_r_reg_23_50 (.CK( clk ) , .D( key_c_r_22_50 ) , .Q( key_c_r_23_50 ) );
  DFF_X1 key_c_r_reg_23_51 (.CK( clk ) , .D( key_c_r_22_51 ) , .Q( key_c_r_23_51 ) );
  DFF_X1 key_c_r_reg_23_52 (.CK( clk ) , .D( key_c_r_22_52 ) , .Q( key_c_r_23_52 ) );
  DFF_X1 key_c_r_reg_23_53 (.CK( clk ) , .D( key_c_r_22_53 ) , .Q( key_c_r_23_53 ) );
  DFF_X1 key_c_r_reg_23_54 (.CK( clk ) , .D( key_c_r_22_54 ) , .Q( key_c_r_23_54 ) );
  DFF_X1 key_c_r_reg_23_55 (.CK( clk ) , .D( key_c_r_22_55 ) , .Q( key_c_r_23_55 ) );
  DFF_X1 key_c_r_reg_23_6 (.CK( clk ) , .D( key_c_r_22_6 ) , .Q( key_c_r_23_6 ) );
  DFF_X1 key_c_r_reg_23_7 (.CK( clk ) , .D( key_c_r_22_7 ) , .Q( key_c_r_23_7 ) );
  DFF_X1 key_c_r_reg_23_8 (.CK( clk ) , .D( key_c_r_22_8 ) , .Q( key_c_r_23_8 ) );
  DFF_X1 key_c_r_reg_23_9 (.CK( clk ) , .D( key_c_r_22_9 ) , .Q( key_c_r_23_9 ) );
  DFF_X1 key_c_r_reg_24_0 (.CK( clk ) , .D( key_c_r_23_0 ) , .Q( key_c_r_24_0 ) );
  DFF_X1 key_c_r_reg_24_1 (.CK( clk ) , .D( key_c_r_23_1 ) , .Q( key_c_r_24_1 ) );
  DFF_X1 key_c_r_reg_24_10 (.CK( clk ) , .D( key_c_r_23_10 ) , .Q( key_c_r_24_10 ) );
  DFF_X1 key_c_r_reg_24_11 (.CK( clk ) , .D( key_c_r_23_11 ) , .Q( key_c_r_24_11 ) );
  DFF_X1 key_c_r_reg_24_12 (.CK( clk ) , .D( key_c_r_23_12 ) , .Q( key_c_r_24_12 ) );
  DFF_X1 key_c_r_reg_24_13 (.CK( clk ) , .D( key_c_r_23_13 ) , .Q( key_c_r_24_13 ) );
  DFF_X1 key_c_r_reg_24_14 (.CK( clk ) , .D( key_c_r_23_14 ) , .Q( key_c_r_24_14 ) );
  DFF_X1 key_c_r_reg_24_15 (.CK( clk ) , .D( key_c_r_23_15 ) , .Q( key_c_r_24_15 ) );
  DFF_X1 key_c_r_reg_24_16 (.CK( clk ) , .D( key_c_r_23_16 ) , .Q( key_c_r_24_16 ) );
  DFF_X1 key_c_r_reg_24_17 (.CK( clk ) , .D( key_c_r_23_17 ) , .Q( key_c_r_24_17 ) );
  DFF_X1 key_c_r_reg_24_18 (.CK( clk ) , .D( key_c_r_23_18 ) , .Q( key_c_r_24_18 ) );
  DFF_X1 key_c_r_reg_24_19 (.CK( clk ) , .D( key_c_r_23_19 ) , .Q( key_c_r_24_19 ) );
  DFF_X1 key_c_r_reg_24_2 (.CK( clk ) , .D( key_c_r_23_2 ) , .Q( key_c_r_24_2 ) );
  DFF_X1 key_c_r_reg_24_20 (.CK( clk ) , .D( key_c_r_23_20 ) , .Q( key_c_r_24_20 ) );
  DFF_X1 key_c_r_reg_24_21 (.CK( clk ) , .D( key_c_r_23_21 ) , .Q( key_c_r_24_21 ) );
  DFF_X1 key_c_r_reg_24_22 (.CK( clk ) , .D( key_c_r_23_22 ) , .Q( key_c_r_24_22 ) );
  DFF_X1 key_c_r_reg_24_23 (.CK( clk ) , .D( key_c_r_23_23 ) , .Q( key_c_r_24_23 ) );
  DFF_X1 key_c_r_reg_24_24 (.CK( clk ) , .D( key_c_r_23_24 ) , .Q( key_c_r_24_24 ) );
  DFF_X1 key_c_r_reg_24_25 (.CK( clk ) , .D( key_c_r_23_25 ) , .Q( key_c_r_24_25 ) );
  DFF_X1 key_c_r_reg_24_26 (.CK( clk ) , .D( key_c_r_23_26 ) , .Q( key_c_r_24_26 ) );
  DFF_X1 key_c_r_reg_24_27 (.CK( clk ) , .D( key_c_r_23_27 ) , .Q( key_c_r_24_27 ) );
  DFF_X1 key_c_r_reg_24_28 (.CK( clk ) , .D( key_c_r_23_28 ) , .Q( key_c_r_24_28 ) );
  DFF_X1 key_c_r_reg_24_29 (.CK( clk ) , .D( key_c_r_23_29 ) , .Q( key_c_r_24_29 ) );
  DFF_X1 key_c_r_reg_24_3 (.CK( clk ) , .D( key_c_r_23_3 ) , .Q( key_c_r_24_3 ) );
  DFF_X1 key_c_r_reg_24_30 (.CK( clk ) , .D( key_c_r_23_30 ) , .Q( key_c_r_24_30 ) );
  DFF_X1 key_c_r_reg_24_31 (.CK( clk ) , .D( key_c_r_23_31 ) , .Q( key_c_r_24_31 ) );
  DFF_X1 key_c_r_reg_24_32 (.CK( clk ) , .D( key_c_r_23_32 ) , .Q( key_c_r_24_32 ) );
  DFF_X1 key_c_r_reg_24_33 (.CK( clk ) , .D( key_c_r_23_33 ) , .Q( key_c_r_24_33 ) );
  DFF_X1 key_c_r_reg_24_34 (.CK( clk ) , .D( key_c_r_23_34 ) , .Q( key_c_r_24_34 ) );
  DFF_X1 key_c_r_reg_24_35 (.CK( clk ) , .D( key_c_r_23_35 ) , .Q( key_c_r_24_35 ) );
  DFF_X1 key_c_r_reg_24_36 (.CK( clk ) , .D( key_c_r_23_36 ) , .Q( key_c_r_24_36 ) );
  DFF_X1 key_c_r_reg_24_37 (.CK( clk ) , .D( key_c_r_23_37 ) , .Q( key_c_r_24_37 ) );
  DFF_X1 key_c_r_reg_24_38 (.CK( clk ) , .D( key_c_r_23_38 ) , .Q( key_c_r_24_38 ) );
  DFF_X1 key_c_r_reg_24_39 (.CK( clk ) , .D( key_c_r_23_39 ) , .Q( key_c_r_24_39 ) );
  DFF_X1 key_c_r_reg_24_4 (.CK( clk ) , .D( key_c_r_23_4 ) , .Q( key_c_r_24_4 ) );
  DFF_X1 key_c_r_reg_24_40 (.CK( clk ) , .D( key_c_r_23_40 ) , .Q( key_c_r_24_40 ) );
  DFF_X1 key_c_r_reg_24_41 (.CK( clk ) , .D( key_c_r_23_41 ) , .Q( key_c_r_24_41 ) );
  DFF_X1 key_c_r_reg_24_42 (.CK( clk ) , .D( key_c_r_23_42 ) , .Q( key_c_r_24_42 ) );
  DFF_X1 key_c_r_reg_24_43 (.CK( clk ) , .D( key_c_r_23_43 ) , .Q( key_c_r_24_43 ) );
  DFF_X1 key_c_r_reg_24_44 (.CK( clk ) , .D( key_c_r_23_44 ) , .Q( key_c_r_24_44 ) );
  DFF_X1 key_c_r_reg_24_45 (.CK( clk ) , .D( key_c_r_23_45 ) , .Q( key_c_r_24_45 ) );
  DFF_X1 key_c_r_reg_24_46 (.CK( clk ) , .D( key_c_r_23_46 ) , .Q( key_c_r_24_46 ) );
  DFF_X1 key_c_r_reg_24_47 (.CK( clk ) , .D( key_c_r_23_47 ) , .Q( key_c_r_24_47 ) );
  DFF_X1 key_c_r_reg_24_48 (.CK( clk ) , .D( key_c_r_23_48 ) , .Q( key_c_r_24_48 ) );
  DFF_X1 key_c_r_reg_24_49 (.CK( clk ) , .D( key_c_r_23_49 ) , .Q( key_c_r_24_49 ) );
  DFF_X1 key_c_r_reg_24_5 (.CK( clk ) , .D( key_c_r_23_5 ) , .Q( key_c_r_24_5 ) );
  DFF_X1 key_c_r_reg_24_50 (.CK( clk ) , .D( key_c_r_23_50 ) , .Q( key_c_r_24_50 ) );
  DFF_X1 key_c_r_reg_24_51 (.CK( clk ) , .D( key_c_r_23_51 ) , .Q( key_c_r_24_51 ) );
  DFF_X1 key_c_r_reg_24_52 (.CK( clk ) , .D( key_c_r_23_52 ) , .Q( key_c_r_24_52 ) );
  DFF_X1 key_c_r_reg_24_53 (.CK( clk ) , .D( key_c_r_23_53 ) , .Q( key_c_r_24_53 ) );
  DFF_X1 key_c_r_reg_24_54 (.CK( clk ) , .D( key_c_r_23_54 ) , .Q( key_c_r_24_54 ) );
  DFF_X1 key_c_r_reg_24_55 (.CK( clk ) , .D( key_c_r_23_55 ) , .Q( key_c_r_24_55 ) );
  DFF_X1 key_c_r_reg_24_6 (.CK( clk ) , .D( key_c_r_23_6 ) , .Q( key_c_r_24_6 ) );
  DFF_X1 key_c_r_reg_24_7 (.CK( clk ) , .D( key_c_r_23_7 ) , .Q( key_c_r_24_7 ) );
  DFF_X1 key_c_r_reg_24_8 (.CK( clk ) , .D( key_c_r_23_8 ) , .Q( key_c_r_24_8 ) );
  DFF_X1 key_c_r_reg_24_9 (.CK( clk ) , .D( key_c_r_23_9 ) , .Q( key_c_r_24_9 ) );
  DFF_X1 key_c_r_reg_25_0 (.CK( clk ) , .D( key_c_r_24_0 ) , .Q( key_c_r_25_0 ) );
  DFF_X1 key_c_r_reg_25_1 (.CK( clk ) , .D( key_c_r_24_1 ) , .Q( key_c_r_25_1 ) );
  DFF_X1 key_c_r_reg_25_10 (.CK( clk ) , .D( key_c_r_24_10 ) , .Q( key_c_r_25_10 ) );
  DFF_X1 key_c_r_reg_25_11 (.CK( clk ) , .D( key_c_r_24_11 ) , .Q( key_c_r_25_11 ) );
  DFF_X1 key_c_r_reg_25_12 (.CK( clk ) , .D( key_c_r_24_12 ) , .Q( key_c_r_25_12 ) );
  DFF_X1 key_c_r_reg_25_13 (.CK( clk ) , .D( key_c_r_24_13 ) , .Q( key_c_r_25_13 ) );
  DFF_X1 key_c_r_reg_25_14 (.CK( clk ) , .D( key_c_r_24_14 ) , .Q( key_c_r_25_14 ) );
  DFF_X1 key_c_r_reg_25_15 (.CK( clk ) , .D( key_c_r_24_15 ) , .Q( key_c_r_25_15 ) );
  DFF_X1 key_c_r_reg_25_16 (.CK( clk ) , .D( key_c_r_24_16 ) , .Q( key_c_r_25_16 ) );
  DFF_X1 key_c_r_reg_25_17 (.CK( clk ) , .D( key_c_r_24_17 ) , .Q( key_c_r_25_17 ) );
  DFF_X1 key_c_r_reg_25_18 (.CK( clk ) , .D( key_c_r_24_18 ) , .Q( key_c_r_25_18 ) );
  DFF_X1 key_c_r_reg_25_19 (.CK( clk ) , .D( key_c_r_24_19 ) , .Q( key_c_r_25_19 ) );
  DFF_X1 key_c_r_reg_25_2 (.CK( clk ) , .D( key_c_r_24_2 ) , .Q( key_c_r_25_2 ) );
  DFF_X1 key_c_r_reg_25_20 (.CK( clk ) , .D( key_c_r_24_20 ) , .Q( key_c_r_25_20 ) );
  DFF_X1 key_c_r_reg_25_21 (.CK( clk ) , .D( key_c_r_24_21 ) , .Q( key_c_r_25_21 ) );
  DFF_X1 key_c_r_reg_25_22 (.CK( clk ) , .D( key_c_r_24_22 ) , .Q( key_c_r_25_22 ) );
  DFF_X1 key_c_r_reg_25_23 (.CK( clk ) , .D( key_c_r_24_23 ) , .Q( key_c_r_25_23 ) );
  DFF_X1 key_c_r_reg_25_24 (.CK( clk ) , .D( key_c_r_24_24 ) , .Q( key_c_r_25_24 ) );
  DFF_X1 key_c_r_reg_25_25 (.CK( clk ) , .D( key_c_r_24_25 ) , .Q( key_c_r_25_25 ) );
  DFF_X1 key_c_r_reg_25_26 (.CK( clk ) , .D( key_c_r_24_26 ) , .Q( key_c_r_25_26 ) );
  DFF_X1 key_c_r_reg_25_27 (.CK( clk ) , .D( key_c_r_24_27 ) , .Q( key_c_r_25_27 ) );
  DFF_X1 key_c_r_reg_25_28 (.CK( clk ) , .D( key_c_r_24_28 ) , .Q( key_c_r_25_28 ) );
  DFF_X1 key_c_r_reg_25_29 (.CK( clk ) , .D( key_c_r_24_29 ) , .Q( key_c_r_25_29 ) );
  DFF_X1 key_c_r_reg_25_3 (.CK( clk ) , .D( key_c_r_24_3 ) , .Q( key_c_r_25_3 ) );
  DFF_X1 key_c_r_reg_25_30 (.CK( clk ) , .D( key_c_r_24_30 ) , .Q( key_c_r_25_30 ) );
  DFF_X1 key_c_r_reg_25_31 (.CK( clk ) , .D( key_c_r_24_31 ) , .Q( key_c_r_25_31 ) );
  DFF_X1 key_c_r_reg_25_32 (.CK( clk ) , .D( key_c_r_24_32 ) , .Q( key_c_r_25_32 ) );
  DFF_X1 key_c_r_reg_25_33 (.CK( clk ) , .D( key_c_r_24_33 ) , .Q( key_c_r_25_33 ) );
  DFF_X1 key_c_r_reg_25_34 (.CK( clk ) , .D( key_c_r_24_34 ) , .Q( key_c_r_25_34 ) );
  DFF_X1 key_c_r_reg_25_35 (.CK( clk ) , .D( key_c_r_24_35 ) , .Q( key_c_r_25_35 ) );
  DFF_X1 key_c_r_reg_25_36 (.CK( clk ) , .D( key_c_r_24_36 ) , .Q( key_c_r_25_36 ) );
  DFF_X1 key_c_r_reg_25_37 (.CK( clk ) , .D( key_c_r_24_37 ) , .Q( key_c_r_25_37 ) );
  DFF_X1 key_c_r_reg_25_38 (.CK( clk ) , .D( key_c_r_24_38 ) , .Q( key_c_r_25_38 ) );
  DFF_X1 key_c_r_reg_25_39 (.CK( clk ) , .D( key_c_r_24_39 ) , .Q( key_c_r_25_39 ) );
  DFF_X1 key_c_r_reg_25_4 (.CK( clk ) , .D( key_c_r_24_4 ) , .Q( key_c_r_25_4 ) );
  DFF_X1 key_c_r_reg_25_40 (.CK( clk ) , .D( key_c_r_24_40 ) , .Q( key_c_r_25_40 ) );
  DFF_X1 key_c_r_reg_25_41 (.CK( clk ) , .D( key_c_r_24_41 ) , .Q( key_c_r_25_41 ) );
  DFF_X1 key_c_r_reg_25_42 (.CK( clk ) , .D( key_c_r_24_42 ) , .Q( key_c_r_25_42 ) );
  DFF_X1 key_c_r_reg_25_43 (.CK( clk ) , .D( key_c_r_24_43 ) , .Q( key_c_r_25_43 ) );
  DFF_X1 key_c_r_reg_25_44 (.CK( clk ) , .D( key_c_r_24_44 ) , .Q( key_c_r_25_44 ) );
  DFF_X1 key_c_r_reg_25_45 (.CK( clk ) , .D( key_c_r_24_45 ) , .Q( key_c_r_25_45 ) );
  DFF_X1 key_c_r_reg_25_46 (.CK( clk ) , .D( key_c_r_24_46 ) , .Q( key_c_r_25_46 ) );
  DFF_X1 key_c_r_reg_25_47 (.CK( clk ) , .D( key_c_r_24_47 ) , .Q( key_c_r_25_47 ) );
  DFF_X1 key_c_r_reg_25_48 (.CK( clk ) , .D( key_c_r_24_48 ) , .Q( key_c_r_25_48 ) );
  DFF_X1 key_c_r_reg_25_49 (.CK( clk ) , .D( key_c_r_24_49 ) , .Q( key_c_r_25_49 ) );
  DFF_X1 key_c_r_reg_25_5 (.CK( clk ) , .D( key_c_r_24_5 ) , .Q( key_c_r_25_5 ) );
  DFF_X1 key_c_r_reg_25_50 (.CK( clk ) , .D( key_c_r_24_50 ) , .Q( key_c_r_25_50 ) );
  DFF_X1 key_c_r_reg_25_51 (.CK( clk ) , .D( key_c_r_24_51 ) , .Q( key_c_r_25_51 ) );
  DFF_X1 key_c_r_reg_25_52 (.CK( clk ) , .D( key_c_r_24_52 ) , .Q( key_c_r_25_52 ) );
  DFF_X1 key_c_r_reg_25_53 (.CK( clk ) , .D( key_c_r_24_53 ) , .Q( key_c_r_25_53 ) );
  DFF_X1 key_c_r_reg_25_54 (.CK( clk ) , .D( key_c_r_24_54 ) , .Q( key_c_r_25_54 ) );
  DFF_X1 key_c_r_reg_25_55 (.CK( clk ) , .D( key_c_r_24_55 ) , .Q( key_c_r_25_55 ) );
  DFF_X1 key_c_r_reg_25_6 (.CK( clk ) , .D( key_c_r_24_6 ) , .Q( key_c_r_25_6 ) );
  DFF_X1 key_c_r_reg_25_7 (.CK( clk ) , .D( key_c_r_24_7 ) , .Q( key_c_r_25_7 ) );
  DFF_X1 key_c_r_reg_25_8 (.CK( clk ) , .D( key_c_r_24_8 ) , .Q( key_c_r_25_8 ) );
  DFF_X1 key_c_r_reg_25_9 (.CK( clk ) , .D( key_c_r_24_9 ) , .Q( key_c_r_25_9 ) );
  DFF_X1 key_c_r_reg_26_0 (.CK( clk ) , .D( key_c_r_25_0 ) , .Q( key_c_r_26_0 ) );
  DFF_X1 key_c_r_reg_26_1 (.CK( clk ) , .D( key_c_r_25_1 ) , .Q( key_c_r_26_1 ) );
  DFF_X1 key_c_r_reg_26_10 (.CK( clk ) , .D( key_c_r_25_10 ) , .Q( key_c_r_26_10 ) );
  DFF_X1 key_c_r_reg_26_11 (.CK( clk ) , .D( key_c_r_25_11 ) , .Q( key_c_r_26_11 ) );
  DFF_X1 key_c_r_reg_26_12 (.CK( clk ) , .D( key_c_r_25_12 ) , .Q( key_c_r_26_12 ) );
  DFF_X1 key_c_r_reg_26_13 (.CK( clk ) , .D( key_c_r_25_13 ) , .Q( key_c_r_26_13 ) );
  DFF_X1 key_c_r_reg_26_14 (.CK( clk ) , .D( key_c_r_25_14 ) , .Q( key_c_r_26_14 ) );
  DFF_X1 key_c_r_reg_26_15 (.CK( clk ) , .D( key_c_r_25_15 ) , .Q( key_c_r_26_15 ) );
  DFF_X1 key_c_r_reg_26_16 (.CK( clk ) , .D( key_c_r_25_16 ) , .Q( key_c_r_26_16 ) );
  DFF_X1 key_c_r_reg_26_17 (.CK( clk ) , .D( key_c_r_25_17 ) , .Q( key_c_r_26_17 ) );
  DFF_X1 key_c_r_reg_26_18 (.CK( clk ) , .D( key_c_r_25_18 ) , .Q( key_c_r_26_18 ) );
  DFF_X1 key_c_r_reg_26_19 (.CK( clk ) , .D( key_c_r_25_19 ) , .Q( key_c_r_26_19 ) );
  DFF_X1 key_c_r_reg_26_2 (.CK( clk ) , .D( key_c_r_25_2 ) , .Q( key_c_r_26_2 ) );
  DFF_X1 key_c_r_reg_26_20 (.CK( clk ) , .D( key_c_r_25_20 ) , .Q( key_c_r_26_20 ) );
  DFF_X1 key_c_r_reg_26_21 (.CK( clk ) , .D( key_c_r_25_21 ) , .Q( key_c_r_26_21 ) );
  DFF_X1 key_c_r_reg_26_22 (.CK( clk ) , .D( key_c_r_25_22 ) , .Q( key_c_r_26_22 ) );
  DFF_X1 key_c_r_reg_26_23 (.CK( clk ) , .D( key_c_r_25_23 ) , .Q( key_c_r_26_23 ) );
  DFF_X1 key_c_r_reg_26_24 (.CK( clk ) , .D( key_c_r_25_24 ) , .Q( key_c_r_26_24 ) );
  DFF_X1 key_c_r_reg_26_25 (.CK( clk ) , .D( key_c_r_25_25 ) , .Q( key_c_r_26_25 ) );
  DFF_X1 key_c_r_reg_26_26 (.CK( clk ) , .D( key_c_r_25_26 ) , .Q( key_c_r_26_26 ) );
  DFF_X1 key_c_r_reg_26_27 (.CK( clk ) , .D( key_c_r_25_27 ) , .Q( key_c_r_26_27 ) );
  DFF_X1 key_c_r_reg_26_28 (.CK( clk ) , .D( key_c_r_25_28 ) , .Q( key_c_r_26_28 ) );
  DFF_X1 key_c_r_reg_26_29 (.CK( clk ) , .D( key_c_r_25_29 ) , .Q( key_c_r_26_29 ) );
  DFF_X1 key_c_r_reg_26_3 (.CK( clk ) , .D( key_c_r_25_3 ) , .Q( key_c_r_26_3 ) );
  DFF_X1 key_c_r_reg_26_30 (.CK( clk ) , .D( key_c_r_25_30 ) , .Q( key_c_r_26_30 ) );
  DFF_X1 key_c_r_reg_26_31 (.CK( clk ) , .D( key_c_r_25_31 ) , .Q( key_c_r_26_31 ) );
  DFF_X1 key_c_r_reg_26_32 (.CK( clk ) , .D( key_c_r_25_32 ) , .Q( key_c_r_26_32 ) );
  DFF_X1 key_c_r_reg_26_33 (.CK( clk ) , .D( key_c_r_25_33 ) , .Q( key_c_r_26_33 ) );
  DFF_X1 key_c_r_reg_26_34 (.CK( clk ) , .D( key_c_r_25_34 ) , .Q( key_c_r_26_34 ) );
  DFF_X1 key_c_r_reg_26_35 (.CK( clk ) , .D( key_c_r_25_35 ) , .Q( key_c_r_26_35 ) );
  DFF_X1 key_c_r_reg_26_36 (.CK( clk ) , .D( key_c_r_25_36 ) , .Q( key_c_r_26_36 ) );
  DFF_X1 key_c_r_reg_26_37 (.CK( clk ) , .D( key_c_r_25_37 ) , .Q( key_c_r_26_37 ) );
  DFF_X1 key_c_r_reg_26_38 (.CK( clk ) , .D( key_c_r_25_38 ) , .Q( key_c_r_26_38 ) );
  DFF_X1 key_c_r_reg_26_39 (.CK( clk ) , .D( key_c_r_25_39 ) , .Q( key_c_r_26_39 ) );
  DFF_X1 key_c_r_reg_26_4 (.CK( clk ) , .D( key_c_r_25_4 ) , .Q( key_c_r_26_4 ) );
  DFF_X1 key_c_r_reg_26_40 (.CK( clk ) , .D( key_c_r_25_40 ) , .Q( key_c_r_26_40 ) );
  DFF_X1 key_c_r_reg_26_41 (.CK( clk ) , .D( key_c_r_25_41 ) , .Q( key_c_r_26_41 ) );
  DFF_X1 key_c_r_reg_26_42 (.CK( clk ) , .D( key_c_r_25_42 ) , .Q( key_c_r_26_42 ) );
  DFF_X1 key_c_r_reg_26_43 (.CK( clk ) , .D( key_c_r_25_43 ) , .Q( key_c_r_26_43 ) );
  DFF_X1 key_c_r_reg_26_44 (.CK( clk ) , .D( key_c_r_25_44 ) , .Q( key_c_r_26_44 ) );
  DFF_X1 key_c_r_reg_26_45 (.CK( clk ) , .D( key_c_r_25_45 ) , .Q( key_c_r_26_45 ) );
  DFF_X1 key_c_r_reg_26_46 (.CK( clk ) , .D( key_c_r_25_46 ) , .Q( key_c_r_26_46 ) );
  DFF_X1 key_c_r_reg_26_47 (.CK( clk ) , .D( key_c_r_25_47 ) , .Q( key_c_r_26_47 ) );
  DFF_X1 key_c_r_reg_26_48 (.CK( clk ) , .D( key_c_r_25_48 ) , .Q( key_c_r_26_48 ) );
  DFF_X1 key_c_r_reg_26_49 (.CK( clk ) , .D( key_c_r_25_49 ) , .Q( key_c_r_26_49 ) );
  DFF_X1 key_c_r_reg_26_5 (.CK( clk ) , .D( key_c_r_25_5 ) , .Q( key_c_r_26_5 ) );
  DFF_X1 key_c_r_reg_26_50 (.CK( clk ) , .D( key_c_r_25_50 ) , .Q( key_c_r_26_50 ) );
  DFF_X1 key_c_r_reg_26_51 (.CK( clk ) , .D( key_c_r_25_51 ) , .Q( key_c_r_26_51 ) );
  DFF_X1 key_c_r_reg_26_52 (.CK( clk ) , .D( key_c_r_25_52 ) , .Q( key_c_r_26_52 ) );
  DFF_X1 key_c_r_reg_26_53 (.CK( clk ) , .D( key_c_r_25_53 ) , .Q( key_c_r_26_53 ) );
  DFF_X1 key_c_r_reg_26_54 (.CK( clk ) , .D( key_c_r_25_54 ) , .Q( key_c_r_26_54 ) );
  DFF_X1 key_c_r_reg_26_55 (.CK( clk ) , .D( key_c_r_25_55 ) , .Q( key_c_r_26_55 ) );
  DFF_X1 key_c_r_reg_26_6 (.CK( clk ) , .D( key_c_r_25_6 ) , .Q( key_c_r_26_6 ) );
  DFF_X1 key_c_r_reg_26_7 (.CK( clk ) , .D( key_c_r_25_7 ) , .Q( key_c_r_26_7 ) );
  DFF_X1 key_c_r_reg_26_8 (.CK( clk ) , .D( key_c_r_25_8 ) , .Q( key_c_r_26_8 ) );
  DFF_X1 key_c_r_reg_26_9 (.CK( clk ) , .D( key_c_r_25_9 ) , .Q( key_c_r_26_9 ) );
  DFF_X1 key_c_r_reg_27_0 (.CK( clk ) , .D( key_c_r_26_0 ) , .Q( key_c_r_27_0 ) );
  DFF_X1 key_c_r_reg_27_1 (.CK( clk ) , .D( key_c_r_26_1 ) , .Q( key_c_r_27_1 ) );
  DFF_X1 key_c_r_reg_27_10 (.CK( clk ) , .D( key_c_r_26_10 ) , .Q( key_c_r_27_10 ) );
  DFF_X1 key_c_r_reg_27_11 (.CK( clk ) , .D( key_c_r_26_11 ) , .Q( key_c_r_27_11 ) );
  DFF_X1 key_c_r_reg_27_12 (.CK( clk ) , .D( key_c_r_26_12 ) , .Q( key_c_r_27_12 ) );
  DFF_X1 key_c_r_reg_27_13 (.CK( clk ) , .D( key_c_r_26_13 ) , .Q( key_c_r_27_13 ) );
  DFF_X1 key_c_r_reg_27_14 (.CK( clk ) , .D( key_c_r_26_14 ) , .Q( key_c_r_27_14 ) );
  DFF_X1 key_c_r_reg_27_15 (.CK( clk ) , .D( key_c_r_26_15 ) , .Q( key_c_r_27_15 ) );
  DFF_X1 key_c_r_reg_27_16 (.CK( clk ) , .D( key_c_r_26_16 ) , .Q( key_c_r_27_16 ) );
  DFF_X1 key_c_r_reg_27_17 (.CK( clk ) , .D( key_c_r_26_17 ) , .Q( key_c_r_27_17 ) );
  DFF_X1 key_c_r_reg_27_18 (.CK( clk ) , .D( key_c_r_26_18 ) , .Q( key_c_r_27_18 ) );
  DFF_X1 key_c_r_reg_27_19 (.CK( clk ) , .D( key_c_r_26_19 ) , .Q( key_c_r_27_19 ) );
  DFF_X1 key_c_r_reg_27_2 (.CK( clk ) , .D( key_c_r_26_2 ) , .Q( key_c_r_27_2 ) );
  DFF_X1 key_c_r_reg_27_20 (.CK( clk ) , .D( key_c_r_26_20 ) , .Q( key_c_r_27_20 ) );
  DFF_X1 key_c_r_reg_27_21 (.CK( clk ) , .D( key_c_r_26_21 ) , .Q( key_c_r_27_21 ) );
  DFF_X1 key_c_r_reg_27_22 (.CK( clk ) , .D( key_c_r_26_22 ) , .Q( key_c_r_27_22 ) );
  DFF_X1 key_c_r_reg_27_23 (.CK( clk ) , .D( key_c_r_26_23 ) , .Q( key_c_r_27_23 ) );
  DFF_X1 key_c_r_reg_27_24 (.CK( clk ) , .D( key_c_r_26_24 ) , .Q( key_c_r_27_24 ) );
  DFF_X1 key_c_r_reg_27_25 (.CK( clk ) , .D( key_c_r_26_25 ) , .Q( key_c_r_27_25 ) );
  DFF_X1 key_c_r_reg_27_26 (.CK( clk ) , .D( key_c_r_26_26 ) , .Q( key_c_r_27_26 ) );
  DFF_X1 key_c_r_reg_27_27 (.CK( clk ) , .D( key_c_r_26_27 ) , .Q( key_c_r_27_27 ) );
  DFF_X1 key_c_r_reg_27_28 (.CK( clk ) , .D( key_c_r_26_28 ) , .Q( key_c_r_27_28 ) );
  DFF_X1 key_c_r_reg_27_29 (.CK( clk ) , .D( key_c_r_26_29 ) , .Q( key_c_r_27_29 ) );
  DFF_X1 key_c_r_reg_27_3 (.CK( clk ) , .D( key_c_r_26_3 ) , .Q( key_c_r_27_3 ) );
  DFF_X1 key_c_r_reg_27_30 (.CK( clk ) , .D( key_c_r_26_30 ) , .Q( key_c_r_27_30 ) );
  DFF_X1 key_c_r_reg_27_31 (.CK( clk ) , .D( key_c_r_26_31 ) , .Q( key_c_r_27_31 ) );
  DFF_X1 key_c_r_reg_27_32 (.CK( clk ) , .D( key_c_r_26_32 ) , .Q( key_c_r_27_32 ) );
  DFF_X1 key_c_r_reg_27_33 (.CK( clk ) , .D( key_c_r_26_33 ) , .Q( key_c_r_27_33 ) );
  DFF_X1 key_c_r_reg_27_34 (.CK( clk ) , .D( key_c_r_26_34 ) , .Q( key_c_r_27_34 ) );
  DFF_X1 key_c_r_reg_27_35 (.CK( clk ) , .D( key_c_r_26_35 ) , .Q( key_c_r_27_35 ) );
  DFF_X1 key_c_r_reg_27_36 (.CK( clk ) , .D( key_c_r_26_36 ) , .Q( key_c_r_27_36 ) );
  DFF_X1 key_c_r_reg_27_37 (.CK( clk ) , .D( key_c_r_26_37 ) , .Q( key_c_r_27_37 ) );
  DFF_X1 key_c_r_reg_27_38 (.CK( clk ) , .D( key_c_r_26_38 ) , .Q( key_c_r_27_38 ) );
  DFF_X1 key_c_r_reg_27_39 (.CK( clk ) , .D( key_c_r_26_39 ) , .Q( key_c_r_27_39 ) );
  DFF_X1 key_c_r_reg_27_4 (.CK( clk ) , .D( key_c_r_26_4 ) , .Q( key_c_r_27_4 ) );
  DFF_X1 key_c_r_reg_27_40 (.CK( clk ) , .D( key_c_r_26_40 ) , .Q( key_c_r_27_40 ) );
  DFF_X1 key_c_r_reg_27_41 (.CK( clk ) , .D( key_c_r_26_41 ) , .Q( key_c_r_27_41 ) );
  DFF_X1 key_c_r_reg_27_42 (.CK( clk ) , .D( key_c_r_26_42 ) , .Q( key_c_r_27_42 ) );
  DFF_X1 key_c_r_reg_27_43 (.CK( clk ) , .D( key_c_r_26_43 ) , .Q( key_c_r_27_43 ) );
  DFF_X1 key_c_r_reg_27_44 (.CK( clk ) , .D( key_c_r_26_44 ) , .Q( key_c_r_27_44 ) );
  DFF_X1 key_c_r_reg_27_45 (.CK( clk ) , .D( key_c_r_26_45 ) , .Q( key_c_r_27_45 ) );
  DFF_X1 key_c_r_reg_27_46 (.CK( clk ) , .D( key_c_r_26_46 ) , .Q( key_c_r_27_46 ) );
  DFF_X1 key_c_r_reg_27_47 (.CK( clk ) , .D( key_c_r_26_47 ) , .Q( key_c_r_27_47 ) );
  DFF_X1 key_c_r_reg_27_48 (.CK( clk ) , .D( key_c_r_26_48 ) , .Q( key_c_r_27_48 ) );
  DFF_X1 key_c_r_reg_27_49 (.CK( clk ) , .D( key_c_r_26_49 ) , .Q( key_c_r_27_49 ) );
  DFF_X1 key_c_r_reg_27_5 (.CK( clk ) , .D( key_c_r_26_5 ) , .Q( key_c_r_27_5 ) );
  DFF_X1 key_c_r_reg_27_50 (.CK( clk ) , .D( key_c_r_26_50 ) , .Q( key_c_r_27_50 ) );
  DFF_X1 key_c_r_reg_27_51 (.CK( clk ) , .D( key_c_r_26_51 ) , .Q( key_c_r_27_51 ) );
  DFF_X1 key_c_r_reg_27_52 (.CK( clk ) , .D( key_c_r_26_52 ) , .Q( key_c_r_27_52 ) );
  DFF_X1 key_c_r_reg_27_53 (.CK( clk ) , .D( key_c_r_26_53 ) , .Q( key_c_r_27_53 ) );
  DFF_X1 key_c_r_reg_27_54 (.CK( clk ) , .D( key_c_r_26_54 ) , .Q( key_c_r_27_54 ) );
  DFF_X1 key_c_r_reg_27_55 (.CK( clk ) , .D( key_c_r_26_55 ) , .Q( key_c_r_27_55 ) );
  DFF_X1 key_c_r_reg_27_6 (.CK( clk ) , .D( key_c_r_26_6 ) , .Q( key_c_r_27_6 ) );
  DFF_X1 key_c_r_reg_27_7 (.CK( clk ) , .D( key_c_r_26_7 ) , .Q( key_c_r_27_7 ) );
  DFF_X1 key_c_r_reg_27_8 (.CK( clk ) , .D( key_c_r_26_8 ) , .Q( key_c_r_27_8 ) );
  DFF_X1 key_c_r_reg_27_9 (.CK( clk ) , .D( key_c_r_26_9 ) , .Q( key_c_r_27_9 ) );
  DFF_X1 key_c_r_reg_28_0 (.CK( clk ) , .D( key_c_r_27_0 ) , .Q( key_c_r_28_0 ) );
  DFF_X1 key_c_r_reg_28_1 (.CK( clk ) , .D( key_c_r_27_1 ) , .Q( key_c_r_28_1 ) );
  DFF_X1 key_c_r_reg_28_10 (.CK( clk ) , .D( key_c_r_27_10 ) , .Q( key_c_r_28_10 ) );
  DFF_X1 key_c_r_reg_28_11 (.CK( clk ) , .D( key_c_r_27_11 ) , .Q( key_c_r_28_11 ) );
  DFF_X1 key_c_r_reg_28_12 (.CK( clk ) , .D( key_c_r_27_12 ) , .Q( key_c_r_28_12 ) );
  DFF_X1 key_c_r_reg_28_13 (.CK( clk ) , .D( key_c_r_27_13 ) , .Q( key_c_r_28_13 ) );
  DFF_X1 key_c_r_reg_28_14 (.CK( clk ) , .D( key_c_r_27_14 ) , .Q( key_c_r_28_14 ) );
  DFF_X1 key_c_r_reg_28_15 (.CK( clk ) , .D( key_c_r_27_15 ) , .Q( key_c_r_28_15 ) );
  DFF_X1 key_c_r_reg_28_16 (.CK( clk ) , .D( key_c_r_27_16 ) , .Q( key_c_r_28_16 ) );
  DFF_X1 key_c_r_reg_28_17 (.CK( clk ) , .D( key_c_r_27_17 ) , .Q( key_c_r_28_17 ) );
  DFF_X1 key_c_r_reg_28_18 (.CK( clk ) , .D( key_c_r_27_18 ) , .Q( key_c_r_28_18 ) );
  DFF_X1 key_c_r_reg_28_19 (.CK( clk ) , .D( key_c_r_27_19 ) , .Q( key_c_r_28_19 ) );
  DFF_X1 key_c_r_reg_28_2 (.CK( clk ) , .D( key_c_r_27_2 ) , .Q( key_c_r_28_2 ) );
  DFF_X1 key_c_r_reg_28_20 (.CK( clk ) , .D( key_c_r_27_20 ) , .Q( key_c_r_28_20 ) );
  DFF_X1 key_c_r_reg_28_21 (.CK( clk ) , .D( key_c_r_27_21 ) , .Q( key_c_r_28_21 ) );
  DFF_X1 key_c_r_reg_28_22 (.CK( clk ) , .D( key_c_r_27_22 ) , .Q( key_c_r_28_22 ) );
  DFF_X1 key_c_r_reg_28_23 (.CK( clk ) , .D( key_c_r_27_23 ) , .Q( key_c_r_28_23 ) );
  DFF_X1 key_c_r_reg_28_24 (.CK( clk ) , .D( key_c_r_27_24 ) , .Q( key_c_r_28_24 ) );
  DFF_X1 key_c_r_reg_28_25 (.CK( clk ) , .D( key_c_r_27_25 ) , .Q( key_c_r_28_25 ) );
  DFF_X1 key_c_r_reg_28_26 (.CK( clk ) , .D( key_c_r_27_26 ) , .Q( key_c_r_28_26 ) );
  DFF_X1 key_c_r_reg_28_27 (.CK( clk ) , .D( key_c_r_27_27 ) , .Q( key_c_r_28_27 ) );
  DFF_X1 key_c_r_reg_28_28 (.CK( clk ) , .D( key_c_r_27_28 ) , .Q( key_c_r_28_28 ) );
  DFF_X1 key_c_r_reg_28_29 (.CK( clk ) , .D( key_c_r_27_29 ) , .Q( key_c_r_28_29 ) );
  DFF_X1 key_c_r_reg_28_3 (.CK( clk ) , .D( key_c_r_27_3 ) , .Q( key_c_r_28_3 ) );
  DFF_X1 key_c_r_reg_28_30 (.CK( clk ) , .D( key_c_r_27_30 ) , .Q( key_c_r_28_30 ) );
  DFF_X1 key_c_r_reg_28_31 (.CK( clk ) , .D( key_c_r_27_31 ) , .Q( key_c_r_28_31 ) );
  DFF_X1 key_c_r_reg_28_32 (.CK( clk ) , .D( key_c_r_27_32 ) , .Q( key_c_r_28_32 ) );
  DFF_X1 key_c_r_reg_28_33 (.CK( clk ) , .D( key_c_r_27_33 ) , .Q( key_c_r_28_33 ) );
  DFF_X1 key_c_r_reg_28_34 (.CK( clk ) , .D( key_c_r_27_34 ) , .Q( key_c_r_28_34 ) );
  DFF_X1 key_c_r_reg_28_35 (.CK( clk ) , .D( key_c_r_27_35 ) , .Q( key_c_r_28_35 ) );
  DFF_X1 key_c_r_reg_28_36 (.CK( clk ) , .D( key_c_r_27_36 ) , .Q( key_c_r_28_36 ) );
  DFF_X1 key_c_r_reg_28_37 (.CK( clk ) , .D( key_c_r_27_37 ) , .Q( key_c_r_28_37 ) );
  DFF_X1 key_c_r_reg_28_38 (.CK( clk ) , .D( key_c_r_27_38 ) , .Q( key_c_r_28_38 ) );
  DFF_X1 key_c_r_reg_28_39 (.CK( clk ) , .D( key_c_r_27_39 ) , .Q( key_c_r_28_39 ) );
  DFF_X1 key_c_r_reg_28_4 (.CK( clk ) , .D( key_c_r_27_4 ) , .Q( key_c_r_28_4 ) );
  DFF_X1 key_c_r_reg_28_40 (.CK( clk ) , .D( key_c_r_27_40 ) , .Q( key_c_r_28_40 ) );
  DFF_X1 key_c_r_reg_28_41 (.CK( clk ) , .D( key_c_r_27_41 ) , .Q( key_c_r_28_41 ) );
  DFF_X1 key_c_r_reg_28_42 (.CK( clk ) , .D( key_c_r_27_42 ) , .Q( key_c_r_28_42 ) );
  DFF_X1 key_c_r_reg_28_43 (.CK( clk ) , .D( key_c_r_27_43 ) , .Q( key_c_r_28_43 ) );
  DFF_X1 key_c_r_reg_28_44 (.CK( clk ) , .D( key_c_r_27_44 ) , .Q( key_c_r_28_44 ) );
  DFF_X1 key_c_r_reg_28_45 (.CK( clk ) , .D( key_c_r_27_45 ) , .Q( key_c_r_28_45 ) );
  DFF_X1 key_c_r_reg_28_46 (.CK( clk ) , .D( key_c_r_27_46 ) , .Q( key_c_r_28_46 ) );
  DFF_X1 key_c_r_reg_28_47 (.CK( clk ) , .D( key_c_r_27_47 ) , .Q( key_c_r_28_47 ) );
  DFF_X1 key_c_r_reg_28_48 (.CK( clk ) , .D( key_c_r_27_48 ) , .Q( key_c_r_28_48 ) );
  DFF_X1 key_c_r_reg_28_49 (.CK( clk ) , .D( key_c_r_27_49 ) , .Q( key_c_r_28_49 ) );
  DFF_X1 key_c_r_reg_28_5 (.CK( clk ) , .D( key_c_r_27_5 ) , .Q( key_c_r_28_5 ) );
  DFF_X1 key_c_r_reg_28_50 (.CK( clk ) , .D( key_c_r_27_50 ) , .Q( key_c_r_28_50 ) );
  DFF_X1 key_c_r_reg_28_51 (.CK( clk ) , .D( key_c_r_27_51 ) , .Q( key_c_r_28_51 ) );
  DFF_X1 key_c_r_reg_28_52 (.CK( clk ) , .D( key_c_r_27_52 ) , .Q( key_c_r_28_52 ) );
  DFF_X1 key_c_r_reg_28_53 (.CK( clk ) , .D( key_c_r_27_53 ) , .Q( key_c_r_28_53 ) );
  DFF_X1 key_c_r_reg_28_54 (.CK( clk ) , .D( key_c_r_27_54 ) , .Q( key_c_r_28_54 ) );
  DFF_X1 key_c_r_reg_28_55 (.CK( clk ) , .D( key_c_r_27_55 ) , .Q( key_c_r_28_55 ) );
  DFF_X1 key_c_r_reg_28_6 (.CK( clk ) , .D( key_c_r_27_6 ) , .Q( key_c_r_28_6 ) );
  DFF_X1 key_c_r_reg_28_7 (.CK( clk ) , .D( key_c_r_27_7 ) , .Q( key_c_r_28_7 ) );
  DFF_X1 key_c_r_reg_28_8 (.CK( clk ) , .D( key_c_r_27_8 ) , .Q( key_c_r_28_8 ) );
  DFF_X1 key_c_r_reg_28_9 (.CK( clk ) , .D( key_c_r_27_9 ) , .Q( key_c_r_28_9 ) );
  DFF_X1 key_c_r_reg_29_0 (.CK( clk ) , .D( key_c_r_28_0 ) , .Q( key_c_r_29_0 ) );
  DFF_X1 key_c_r_reg_29_1 (.CK( clk ) , .D( key_c_r_28_1 ) , .Q( key_c_r_29_1 ) );
  DFF_X1 key_c_r_reg_29_10 (.CK( clk ) , .D( key_c_r_28_10 ) , .Q( key_c_r_29_10 ) );
  DFF_X1 key_c_r_reg_29_11 (.CK( clk ) , .D( key_c_r_28_11 ) , .Q( key_c_r_29_11 ) );
  DFF_X1 key_c_r_reg_29_12 (.CK( clk ) , .D( key_c_r_28_12 ) , .Q( key_c_r_29_12 ) );
  DFF_X1 key_c_r_reg_29_13 (.CK( clk ) , .D( key_c_r_28_13 ) , .Q( key_c_r_29_13 ) );
  DFF_X1 key_c_r_reg_29_14 (.CK( clk ) , .D( key_c_r_28_14 ) , .Q( key_c_r_29_14 ) );
  DFF_X1 key_c_r_reg_29_15 (.CK( clk ) , .D( key_c_r_28_15 ) , .Q( key_c_r_29_15 ) );
  DFF_X1 key_c_r_reg_29_16 (.CK( clk ) , .D( key_c_r_28_16 ) , .Q( key_c_r_29_16 ) );
  DFF_X1 key_c_r_reg_29_17 (.CK( clk ) , .D( key_c_r_28_17 ) , .Q( key_c_r_29_17 ) );
  DFF_X1 key_c_r_reg_29_18 (.CK( clk ) , .D( key_c_r_28_18 ) , .Q( key_c_r_29_18 ) );
  DFF_X1 key_c_r_reg_29_19 (.CK( clk ) , .D( key_c_r_28_19 ) , .Q( key_c_r_29_19 ) );
  DFF_X1 key_c_r_reg_29_2 (.CK( clk ) , .D( key_c_r_28_2 ) , .Q( key_c_r_29_2 ) );
  DFF_X1 key_c_r_reg_29_20 (.CK( clk ) , .D( key_c_r_28_20 ) , .Q( key_c_r_29_20 ) );
  DFF_X1 key_c_r_reg_29_21 (.CK( clk ) , .D( key_c_r_28_21 ) , .Q( key_c_r_29_21 ) );
  DFF_X1 key_c_r_reg_29_22 (.CK( clk ) , .D( key_c_r_28_22 ) , .Q( key_c_r_29_22 ) );
  DFF_X1 key_c_r_reg_29_23 (.CK( clk ) , .D( key_c_r_28_23 ) , .Q( key_c_r_29_23 ) );
  DFF_X1 key_c_r_reg_29_24 (.CK( clk ) , .D( key_c_r_28_24 ) , .Q( key_c_r_29_24 ) );
  DFF_X1 key_c_r_reg_29_25 (.CK( clk ) , .D( key_c_r_28_25 ) , .Q( key_c_r_29_25 ) );
  DFF_X1 key_c_r_reg_29_26 (.CK( clk ) , .D( key_c_r_28_26 ) , .Q( key_c_r_29_26 ) );
  DFF_X1 key_c_r_reg_29_27 (.CK( clk ) , .D( key_c_r_28_27 ) , .Q( key_c_r_29_27 ) );
  DFF_X1 key_c_r_reg_29_28 (.CK( clk ) , .D( key_c_r_28_28 ) , .Q( key_c_r_29_28 ) );
  DFF_X1 key_c_r_reg_29_29 (.CK( clk ) , .D( key_c_r_28_29 ) , .Q( key_c_r_29_29 ) );
  DFF_X1 key_c_r_reg_29_3 (.CK( clk ) , .D( key_c_r_28_3 ) , .Q( key_c_r_29_3 ) );
  DFF_X1 key_c_r_reg_29_30 (.CK( clk ) , .D( key_c_r_28_30 ) , .Q( key_c_r_29_30 ) );
  DFF_X1 key_c_r_reg_29_31 (.CK( clk ) , .D( key_c_r_28_31 ) , .Q( key_c_r_29_31 ) );
  DFF_X1 key_c_r_reg_29_32 (.CK( clk ) , .D( key_c_r_28_32 ) , .Q( key_c_r_29_32 ) );
  DFF_X1 key_c_r_reg_29_33 (.CK( clk ) , .D( key_c_r_28_33 ) , .Q( key_c_r_29_33 ) );
  DFF_X1 key_c_r_reg_29_34 (.CK( clk ) , .D( key_c_r_28_34 ) , .Q( key_c_r_29_34 ) );
  DFF_X1 key_c_r_reg_29_35 (.CK( clk ) , .D( key_c_r_28_35 ) , .Q( key_c_r_29_35 ) );
  DFF_X1 key_c_r_reg_29_36 (.CK( clk ) , .D( key_c_r_28_36 ) , .Q( key_c_r_29_36 ) );
  DFF_X1 key_c_r_reg_29_37 (.CK( clk ) , .D( key_c_r_28_37 ) , .Q( key_c_r_29_37 ) );
  DFF_X1 key_c_r_reg_29_38 (.CK( clk ) , .D( key_c_r_28_38 ) , .Q( key_c_r_29_38 ) );
  DFF_X1 key_c_r_reg_29_39 (.CK( clk ) , .D( key_c_r_28_39 ) , .Q( key_c_r_29_39 ) );
  DFF_X1 key_c_r_reg_29_4 (.CK( clk ) , .D( key_c_r_28_4 ) , .Q( key_c_r_29_4 ) );
  DFF_X1 key_c_r_reg_29_40 (.CK( clk ) , .D( key_c_r_28_40 ) , .Q( key_c_r_29_40 ) );
  DFF_X1 key_c_r_reg_29_41 (.CK( clk ) , .D( key_c_r_28_41 ) , .Q( key_c_r_29_41 ) );
  DFF_X1 key_c_r_reg_29_42 (.CK( clk ) , .D( key_c_r_28_42 ) , .Q( key_c_r_29_42 ) );
  DFF_X1 key_c_r_reg_29_43 (.CK( clk ) , .D( key_c_r_28_43 ) , .Q( key_c_r_29_43 ) );
  DFF_X1 key_c_r_reg_29_44 (.CK( clk ) , .D( key_c_r_28_44 ) , .Q( key_c_r_29_44 ) );
  DFF_X1 key_c_r_reg_29_45 (.CK( clk ) , .D( key_c_r_28_45 ) , .Q( key_c_r_29_45 ) );
  DFF_X1 key_c_r_reg_29_46 (.CK( clk ) , .D( key_c_r_28_46 ) , .Q( key_c_r_29_46 ) );
  DFF_X1 key_c_r_reg_29_47 (.CK( clk ) , .D( key_c_r_28_47 ) , .Q( key_c_r_29_47 ) );
  DFF_X1 key_c_r_reg_29_48 (.CK( clk ) , .D( key_c_r_28_48 ) , .Q( key_c_r_29_48 ) );
  DFF_X1 key_c_r_reg_29_49 (.CK( clk ) , .D( key_c_r_28_49 ) , .Q( key_c_r_29_49 ) );
  DFF_X1 key_c_r_reg_29_5 (.CK( clk ) , .D( key_c_r_28_5 ) , .Q( key_c_r_29_5 ) );
  DFF_X1 key_c_r_reg_29_50 (.CK( clk ) , .D( key_c_r_28_50 ) , .Q( key_c_r_29_50 ) );
  DFF_X1 key_c_r_reg_29_51 (.CK( clk ) , .D( key_c_r_28_51 ) , .Q( key_c_r_29_51 ) );
  DFF_X1 key_c_r_reg_29_52 (.CK( clk ) , .D( key_c_r_28_52 ) , .Q( key_c_r_29_52 ) );
  DFF_X1 key_c_r_reg_29_53 (.CK( clk ) , .D( key_c_r_28_53 ) , .Q( key_c_r_29_53 ) );
  DFF_X1 key_c_r_reg_29_54 (.CK( clk ) , .D( key_c_r_28_54 ) , .Q( key_c_r_29_54 ) );
  DFF_X1 key_c_r_reg_29_55 (.CK( clk ) , .D( key_c_r_28_55 ) , .Q( key_c_r_29_55 ) );
  DFF_X1 key_c_r_reg_29_6 (.CK( clk ) , .D( key_c_r_28_6 ) , .Q( key_c_r_29_6 ) );
  DFF_X1 key_c_r_reg_29_7 (.CK( clk ) , .D( key_c_r_28_7 ) , .Q( key_c_r_29_7 ) );
  DFF_X1 key_c_r_reg_29_8 (.CK( clk ) , .D( key_c_r_28_8 ) , .Q( key_c_r_29_8 ) );
  DFF_X1 key_c_r_reg_29_9 (.CK( clk ) , .D( key_c_r_28_9 ) , .Q( key_c_r_29_9 ) );
  DFF_X1 key_c_r_reg_2_0 (.CK( clk ) , .D( key_c_r_1_0 ) , .Q( key_c_r_2_0 ) );
  DFF_X1 key_c_r_reg_2_1 (.CK( clk ) , .D( key_c_r_1_1 ) , .Q( key_c_r_2_1 ) );
  DFF_X1 key_c_r_reg_2_10 (.CK( clk ) , .D( key_c_r_1_10 ) , .Q( key_c_r_2_10 ) );
  DFF_X1 key_c_r_reg_2_11 (.CK( clk ) , .D( key_c_r_1_11 ) , .Q( key_c_r_2_11 ) );
  DFF_X1 key_c_r_reg_2_12 (.CK( clk ) , .D( key_c_r_1_12 ) , .Q( key_c_r_2_12 ) );
  DFF_X1 key_c_r_reg_2_13 (.CK( clk ) , .D( key_c_r_1_13 ) , .Q( key_c_r_2_13 ) );
  DFF_X1 key_c_r_reg_2_14 (.CK( clk ) , .D( key_c_r_1_14 ) , .Q( key_c_r_2_14 ) );
  DFF_X1 key_c_r_reg_2_15 (.CK( clk ) , .D( key_c_r_1_15 ) , .Q( key_c_r_2_15 ) );
  DFF_X1 key_c_r_reg_2_16 (.CK( clk ) , .D( key_c_r_1_16 ) , .Q( key_c_r_2_16 ) );
  DFF_X1 key_c_r_reg_2_17 (.CK( clk ) , .D( key_c_r_1_17 ) , .Q( key_c_r_2_17 ) );
  DFF_X1 key_c_r_reg_2_18 (.CK( clk ) , .D( key_c_r_1_18 ) , .Q( key_c_r_2_18 ) );
  DFF_X1 key_c_r_reg_2_19 (.CK( clk ) , .D( key_c_r_1_19 ) , .Q( key_c_r_2_19 ) );
  DFF_X1 key_c_r_reg_2_2 (.CK( clk ) , .D( key_c_r_1_2 ) , .Q( key_c_r_2_2 ) );
  DFF_X1 key_c_r_reg_2_20 (.CK( clk ) , .D( key_c_r_1_20 ) , .Q( key_c_r_2_20 ) );
  DFF_X1 key_c_r_reg_2_21 (.CK( clk ) , .D( key_c_r_1_21 ) , .Q( key_c_r_2_21 ) );
  DFF_X1 key_c_r_reg_2_22 (.CK( clk ) , .D( key_c_r_1_22 ) , .Q( key_c_r_2_22 ) );
  DFF_X1 key_c_r_reg_2_23 (.CK( clk ) , .D( key_c_r_1_23 ) , .Q( key_c_r_2_23 ) );
  DFF_X1 key_c_r_reg_2_24 (.CK( clk ) , .D( key_c_r_1_24 ) , .Q( key_c_r_2_24 ) );
  DFF_X1 key_c_r_reg_2_25 (.CK( clk ) , .D( key_c_r_1_25 ) , .Q( key_c_r_2_25 ) );
  DFF_X1 key_c_r_reg_2_26 (.CK( clk ) , .D( key_c_r_1_26 ) , .Q( key_c_r_2_26 ) );
  DFF_X1 key_c_r_reg_2_27 (.CK( clk ) , .D( key_c_r_1_27 ) , .Q( key_c_r_2_27 ) );
  DFF_X1 key_c_r_reg_2_28 (.CK( clk ) , .D( key_c_r_1_28 ) , .Q( key_c_r_2_28 ) );
  DFF_X1 key_c_r_reg_2_29 (.CK( clk ) , .D( key_c_r_1_29 ) , .Q( key_c_r_2_29 ) );
  DFF_X1 key_c_r_reg_2_3 (.CK( clk ) , .D( key_c_r_1_3 ) , .Q( key_c_r_2_3 ) );
  DFF_X1 key_c_r_reg_2_30 (.CK( clk ) , .D( key_c_r_1_30 ) , .Q( key_c_r_2_30 ) );
  DFF_X1 key_c_r_reg_2_31 (.CK( clk ) , .D( key_c_r_1_31 ) , .Q( key_c_r_2_31 ) );
  DFF_X1 key_c_r_reg_2_32 (.CK( clk ) , .D( key_c_r_1_32 ) , .Q( key_c_r_2_32 ) );
  DFF_X1 key_c_r_reg_2_33 (.CK( clk ) , .D( key_c_r_1_33 ) , .Q( key_c_r_2_33 ) );
  DFF_X1 key_c_r_reg_2_34 (.CK( clk ) , .D( key_c_r_1_34 ) , .Q( key_c_r_2_34 ) );
  DFF_X1 key_c_r_reg_2_35 (.CK( clk ) , .D( key_c_r_1_35 ) , .Q( key_c_r_2_35 ) );
  DFF_X1 key_c_r_reg_2_36 (.CK( clk ) , .D( key_c_r_1_36 ) , .Q( key_c_r_2_36 ) );
  DFF_X1 key_c_r_reg_2_37 (.CK( clk ) , .D( key_c_r_1_37 ) , .Q( key_c_r_2_37 ) );
  DFF_X1 key_c_r_reg_2_38 (.CK( clk ) , .D( key_c_r_1_38 ) , .Q( key_c_r_2_38 ) );
  DFF_X1 key_c_r_reg_2_39 (.CK( clk ) , .D( key_c_r_1_39 ) , .Q( key_c_r_2_39 ) );
  DFF_X1 key_c_r_reg_2_4 (.CK( clk ) , .D( key_c_r_1_4 ) , .Q( key_c_r_2_4 ) );
  DFF_X1 key_c_r_reg_2_40 (.CK( clk ) , .D( key_c_r_1_40 ) , .Q( key_c_r_2_40 ) );
  DFF_X1 key_c_r_reg_2_41 (.CK( clk ) , .D( key_c_r_1_41 ) , .Q( key_c_r_2_41 ) );
  DFF_X1 key_c_r_reg_2_42 (.CK( clk ) , .D( key_c_r_1_42 ) , .Q( key_c_r_2_42 ) );
  DFF_X1 key_c_r_reg_2_43 (.CK( clk ) , .D( key_c_r_1_43 ) , .Q( key_c_r_2_43 ) );
  DFF_X1 key_c_r_reg_2_44 (.CK( clk ) , .D( key_c_r_1_44 ) , .Q( key_c_r_2_44 ) );
  DFF_X1 key_c_r_reg_2_45 (.CK( clk ) , .D( key_c_r_1_45 ) , .Q( key_c_r_2_45 ) );
  DFF_X1 key_c_r_reg_2_46 (.CK( clk ) , .D( key_c_r_1_46 ) , .Q( key_c_r_2_46 ) );
  DFF_X1 key_c_r_reg_2_47 (.CK( clk ) , .D( key_c_r_1_47 ) , .Q( key_c_r_2_47 ) );
  DFF_X1 key_c_r_reg_2_48 (.CK( clk ) , .D( key_c_r_1_48 ) , .Q( key_c_r_2_48 ) );
  DFF_X1 key_c_r_reg_2_49 (.CK( clk ) , .D( key_c_r_1_49 ) , .Q( key_c_r_2_49 ) );
  DFF_X1 key_c_r_reg_2_5 (.CK( clk ) , .D( key_c_r_1_5 ) , .Q( key_c_r_2_5 ) );
  DFF_X1 key_c_r_reg_2_50 (.CK( clk ) , .D( key_c_r_1_50 ) , .Q( key_c_r_2_50 ) );
  DFF_X1 key_c_r_reg_2_51 (.CK( clk ) , .D( key_c_r_1_51 ) , .Q( key_c_r_2_51 ) );
  DFF_X1 key_c_r_reg_2_52 (.CK( clk ) , .D( key_c_r_1_52 ) , .Q( key_c_r_2_52 ) );
  DFF_X1 key_c_r_reg_2_53 (.CK( clk ) , .D( key_c_r_1_53 ) , .Q( key_c_r_2_53 ) );
  DFF_X1 key_c_r_reg_2_54 (.CK( clk ) , .D( key_c_r_1_54 ) , .Q( key_c_r_2_54 ) );
  DFF_X1 key_c_r_reg_2_55 (.CK( clk ) , .D( key_c_r_1_55 ) , .Q( key_c_r_2_55 ) );
  DFF_X1 key_c_r_reg_2_6 (.CK( clk ) , .D( key_c_r_1_6 ) , .Q( key_c_r_2_6 ) );
  DFF_X1 key_c_r_reg_2_7 (.CK( clk ) , .D( key_c_r_1_7 ) , .Q( key_c_r_2_7 ) );
  DFF_X1 key_c_r_reg_2_8 (.CK( clk ) , .D( key_c_r_1_8 ) , .Q( key_c_r_2_8 ) );
  DFF_X1 key_c_r_reg_2_9 (.CK( clk ) , .D( key_c_r_1_9 ) , .Q( key_c_r_2_9 ) );
  DFF_X1 key_c_r_reg_30_0 (.CK( clk ) , .D( key_c_r_29_0 ) , .Q( key_c_r_30_0 ) );
  DFF_X1 key_c_r_reg_30_1 (.CK( clk ) , .D( key_c_r_29_1 ) , .Q( key_c_r_30_1 ) );
  DFF_X1 key_c_r_reg_30_10 (.CK( clk ) , .D( key_c_r_29_10 ) , .Q( key_c_r_30_10 ) );
  DFF_X1 key_c_r_reg_30_11 (.CK( clk ) , .D( key_c_r_29_11 ) , .Q( key_c_r_30_11 ) );
  DFF_X1 key_c_r_reg_30_12 (.CK( clk ) , .D( key_c_r_29_12 ) , .Q( key_c_r_30_12 ) );
  DFF_X1 key_c_r_reg_30_13 (.CK( clk ) , .D( key_c_r_29_13 ) , .Q( key_c_r_30_13 ) );
  DFF_X1 key_c_r_reg_30_14 (.CK( clk ) , .D( key_c_r_29_14 ) , .Q( key_c_r_30_14 ) );
  DFF_X1 key_c_r_reg_30_15 (.CK( clk ) , .D( key_c_r_29_15 ) , .Q( key_c_r_30_15 ) );
  DFF_X1 key_c_r_reg_30_16 (.CK( clk ) , .D( key_c_r_29_16 ) , .Q( key_c_r_30_16 ) );
  DFF_X1 key_c_r_reg_30_17 (.CK( clk ) , .D( key_c_r_29_17 ) , .Q( key_c_r_30_17 ) );
  DFF_X1 key_c_r_reg_30_18 (.CK( clk ) , .D( key_c_r_29_18 ) , .Q( key_c_r_30_18 ) );
  DFF_X1 key_c_r_reg_30_19 (.CK( clk ) , .D( key_c_r_29_19 ) , .Q( key_c_r_30_19 ) );
  DFF_X1 key_c_r_reg_30_2 (.CK( clk ) , .D( key_c_r_29_2 ) , .Q( key_c_r_30_2 ) );
  DFF_X1 key_c_r_reg_30_20 (.CK( clk ) , .D( key_c_r_29_20 ) , .Q( key_c_r_30_20 ) );
  DFF_X1 key_c_r_reg_30_21 (.CK( clk ) , .D( key_c_r_29_21 ) , .Q( key_c_r_30_21 ) );
  DFF_X1 key_c_r_reg_30_22 (.CK( clk ) , .D( key_c_r_29_22 ) , .Q( key_c_r_30_22 ) );
  DFF_X1 key_c_r_reg_30_23 (.CK( clk ) , .D( key_c_r_29_23 ) , .Q( key_c_r_30_23 ) );
  DFF_X1 key_c_r_reg_30_24 (.CK( clk ) , .D( key_c_r_29_24 ) , .Q( key_c_r_30_24 ) );
  DFF_X1 key_c_r_reg_30_25 (.CK( clk ) , .D( key_c_r_29_25 ) , .Q( key_c_r_30_25 ) );
  DFF_X1 key_c_r_reg_30_26 (.CK( clk ) , .D( key_c_r_29_26 ) , .Q( key_c_r_30_26 ) );
  DFF_X1 key_c_r_reg_30_27 (.CK( clk ) , .D( key_c_r_29_27 ) , .Q( key_c_r_30_27 ) );
  DFF_X1 key_c_r_reg_30_28 (.CK( clk ) , .D( key_c_r_29_28 ) , .Q( key_c_r_30_28 ) );
  DFF_X1 key_c_r_reg_30_29 (.CK( clk ) , .D( key_c_r_29_29 ) , .Q( key_c_r_30_29 ) );
  DFF_X1 key_c_r_reg_30_3 (.CK( clk ) , .D( key_c_r_29_3 ) , .Q( key_c_r_30_3 ) );
  DFF_X1 key_c_r_reg_30_30 (.CK( clk ) , .D( key_c_r_29_30 ) , .Q( key_c_r_30_30 ) );
  DFF_X1 key_c_r_reg_30_31 (.CK( clk ) , .D( key_c_r_29_31 ) , .Q( key_c_r_30_31 ) );
  DFF_X1 key_c_r_reg_30_32 (.CK( clk ) , .D( key_c_r_29_32 ) , .Q( key_c_r_30_32 ) );
  DFF_X1 key_c_r_reg_30_33 (.CK( clk ) , .D( key_c_r_29_33 ) , .Q( key_c_r_30_33 ) );
  DFF_X1 key_c_r_reg_30_34 (.CK( clk ) , .D( key_c_r_29_34 ) , .Q( key_c_r_30_34 ) );
  DFF_X1 key_c_r_reg_30_35 (.CK( clk ) , .D( key_c_r_29_35 ) , .Q( key_c_r_30_35 ) );
  DFF_X1 key_c_r_reg_30_36 (.CK( clk ) , .D( key_c_r_29_36 ) , .Q( key_c_r_30_36 ) );
  DFF_X1 key_c_r_reg_30_37 (.CK( clk ) , .D( key_c_r_29_37 ) , .Q( key_c_r_30_37 ) );
  DFF_X1 key_c_r_reg_30_38 (.CK( clk ) , .D( key_c_r_29_38 ) , .Q( key_c_r_30_38 ) );
  DFF_X1 key_c_r_reg_30_39 (.CK( clk ) , .D( key_c_r_29_39 ) , .Q( key_c_r_30_39 ) );
  DFF_X1 key_c_r_reg_30_4 (.CK( clk ) , .D( key_c_r_29_4 ) , .Q( key_c_r_30_4 ) );
  DFF_X1 key_c_r_reg_30_40 (.CK( clk ) , .D( key_c_r_29_40 ) , .Q( key_c_r_30_40 ) );
  DFF_X1 key_c_r_reg_30_41 (.CK( clk ) , .D( key_c_r_29_41 ) , .Q( key_c_r_30_41 ) );
  DFF_X1 key_c_r_reg_30_42 (.CK( clk ) , .D( key_c_r_29_42 ) , .Q( key_c_r_30_42 ) );
  DFF_X1 key_c_r_reg_30_43 (.CK( clk ) , .D( key_c_r_29_43 ) , .Q( key_c_r_30_43 ) );
  DFF_X1 key_c_r_reg_30_44 (.CK( clk ) , .D( key_c_r_29_44 ) , .Q( key_c_r_30_44 ) );
  DFF_X1 key_c_r_reg_30_45 (.CK( clk ) , .D( key_c_r_29_45 ) , .Q( key_c_r_30_45 ) );
  DFF_X1 key_c_r_reg_30_46 (.CK( clk ) , .D( key_c_r_29_46 ) , .Q( key_c_r_30_46 ) );
  DFF_X1 key_c_r_reg_30_47 (.CK( clk ) , .D( key_c_r_29_47 ) , .Q( key_c_r_30_47 ) );
  DFF_X1 key_c_r_reg_30_48 (.CK( clk ) , .D( key_c_r_29_48 ) , .Q( key_c_r_30_48 ) );
  DFF_X1 key_c_r_reg_30_49 (.CK( clk ) , .D( key_c_r_29_49 ) , .Q( key_c_r_30_49 ) );
  DFF_X1 key_c_r_reg_30_5 (.CK( clk ) , .D( key_c_r_29_5 ) , .Q( key_c_r_30_5 ) );
  DFF_X1 key_c_r_reg_30_50 (.CK( clk ) , .D( key_c_r_29_50 ) , .Q( key_c_r_30_50 ) );
  DFF_X1 key_c_r_reg_30_51 (.CK( clk ) , .D( key_c_r_29_51 ) , .Q( key_c_r_30_51 ) );
  DFF_X1 key_c_r_reg_30_52 (.CK( clk ) , .D( key_c_r_29_52 ) , .Q( key_c_r_30_52 ) );
  DFF_X1 key_c_r_reg_30_53 (.CK( clk ) , .D( key_c_r_29_53 ) , .Q( key_c_r_30_53 ) );
  DFF_X1 key_c_r_reg_30_54 (.CK( clk ) , .D( key_c_r_29_54 ) , .Q( key_c_r_30_54 ) );
  DFF_X1 key_c_r_reg_30_55 (.CK( clk ) , .D( key_c_r_29_55 ) , .Q( key_c_r_30_55 ) );
  DFF_X1 key_c_r_reg_30_6 (.CK( clk ) , .D( key_c_r_29_6 ) , .Q( key_c_r_30_6 ) );
  DFF_X1 key_c_r_reg_30_7 (.CK( clk ) , .D( key_c_r_29_7 ) , .Q( key_c_r_30_7 ) );
  DFF_X1 key_c_r_reg_30_8 (.CK( clk ) , .D( key_c_r_29_8 ) , .Q( key_c_r_30_8 ) );
  DFF_X1 key_c_r_reg_30_9 (.CK( clk ) , .D( key_c_r_29_9 ) , .Q( key_c_r_30_9 ) );
  DFF_X1 key_c_r_reg_31_0 (.CK( clk ) , .D( key_c_r_30_0 ) , .Q( key_c_r_31_0 ) );
  DFF_X1 key_c_r_reg_31_1 (.CK( clk ) , .D( key_c_r_30_1 ) , .Q( key_c_r_31_1 ) );
  DFF_X1 key_c_r_reg_31_10 (.CK( clk ) , .D( key_c_r_30_10 ) , .Q( key_c_r_31_10 ) );
  DFF_X1 key_c_r_reg_31_11 (.CK( clk ) , .D( key_c_r_30_11 ) , .Q( key_c_r_31_11 ) );
  DFF_X1 key_c_r_reg_31_12 (.CK( clk ) , .D( key_c_r_30_12 ) , .Q( key_c_r_31_12 ) );
  DFF_X1 key_c_r_reg_31_13 (.CK( clk ) , .D( key_c_r_30_13 ) , .Q( key_c_r_31_13 ) );
  DFF_X1 key_c_r_reg_31_14 (.CK( clk ) , .D( key_c_r_30_14 ) , .Q( key_c_r_31_14 ) );
  DFF_X1 key_c_r_reg_31_15 (.CK( clk ) , .D( key_c_r_30_15 ) , .Q( key_c_r_31_15 ) );
  DFF_X1 key_c_r_reg_31_16 (.CK( clk ) , .D( key_c_r_30_16 ) , .Q( key_c_r_31_16 ) );
  DFF_X1 key_c_r_reg_31_17 (.CK( clk ) , .D( key_c_r_30_17 ) , .Q( key_c_r_31_17 ) );
  DFF_X1 key_c_r_reg_31_18 (.CK( clk ) , .D( key_c_r_30_18 ) , .Q( key_c_r_31_18 ) );
  DFF_X1 key_c_r_reg_31_19 (.CK( clk ) , .D( key_c_r_30_19 ) , .Q( key_c_r_31_19 ) );
  DFF_X1 key_c_r_reg_31_2 (.CK( clk ) , .D( key_c_r_30_2 ) , .Q( key_c_r_31_2 ) );
  DFF_X1 key_c_r_reg_31_20 (.CK( clk ) , .D( key_c_r_30_20 ) , .Q( key_c_r_31_20 ) );
  DFF_X1 key_c_r_reg_31_21 (.CK( clk ) , .D( key_c_r_30_21 ) , .Q( key_c_r_31_21 ) );
  DFF_X1 key_c_r_reg_31_22 (.CK( clk ) , .D( key_c_r_30_22 ) , .Q( key_c_r_31_22 ) );
  DFF_X1 key_c_r_reg_31_23 (.CK( clk ) , .D( key_c_r_30_23 ) , .Q( key_c_r_31_23 ) );
  DFF_X1 key_c_r_reg_31_24 (.CK( clk ) , .D( key_c_r_30_24 ) , .Q( key_c_r_31_24 ) );
  DFF_X1 key_c_r_reg_31_25 (.CK( clk ) , .D( key_c_r_30_25 ) , .Q( key_c_r_31_25 ) );
  DFF_X1 key_c_r_reg_31_26 (.CK( clk ) , .D( key_c_r_30_26 ) , .Q( key_c_r_31_26 ) );
  DFF_X1 key_c_r_reg_31_27 (.CK( clk ) , .D( key_c_r_30_27 ) , .Q( key_c_r_31_27 ) );
  DFF_X1 key_c_r_reg_31_28 (.CK( clk ) , .D( key_c_r_30_28 ) , .Q( key_c_r_31_28 ) );
  DFF_X1 key_c_r_reg_31_29 (.CK( clk ) , .D( key_c_r_30_29 ) , .Q( key_c_r_31_29 ) );
  DFF_X1 key_c_r_reg_31_3 (.CK( clk ) , .D( key_c_r_30_3 ) , .Q( key_c_r_31_3 ) );
  DFF_X1 key_c_r_reg_31_30 (.CK( clk ) , .D( key_c_r_30_30 ) , .Q( key_c_r_31_30 ) );
  DFF_X1 key_c_r_reg_31_31 (.CK( clk ) , .D( key_c_r_30_31 ) , .Q( key_c_r_31_31 ) );
  DFF_X1 key_c_r_reg_31_32 (.CK( clk ) , .D( key_c_r_30_32 ) , .Q( key_c_r_31_32 ) );
  DFF_X1 key_c_r_reg_31_33 (.CK( clk ) , .D( key_c_r_30_33 ) , .Q( key_c_r_31_33 ) );
  DFF_X1 key_c_r_reg_31_34 (.CK( clk ) , .D( key_c_r_30_34 ) , .Q( key_c_r_31_34 ) );
  DFF_X1 key_c_r_reg_31_35 (.CK( clk ) , .D( key_c_r_30_35 ) , .Q( key_c_r_31_35 ) );
  DFF_X1 key_c_r_reg_31_36 (.CK( clk ) , .D( key_c_r_30_36 ) , .Q( key_c_r_31_36 ) );
  DFF_X1 key_c_r_reg_31_37 (.CK( clk ) , .D( key_c_r_30_37 ) , .Q( key_c_r_31_37 ) );
  DFF_X1 key_c_r_reg_31_38 (.CK( clk ) , .D( key_c_r_30_38 ) , .Q( key_c_r_31_38 ) );
  DFF_X1 key_c_r_reg_31_39 (.CK( clk ) , .D( key_c_r_30_39 ) , .Q( key_c_r_31_39 ) );
  DFF_X1 key_c_r_reg_31_4 (.CK( clk ) , .D( key_c_r_30_4 ) , .Q( key_c_r_31_4 ) );
  DFF_X1 key_c_r_reg_31_40 (.CK( clk ) , .D( key_c_r_30_40 ) , .Q( key_c_r_31_40 ) );
  DFF_X1 key_c_r_reg_31_41 (.CK( clk ) , .D( key_c_r_30_41 ) , .Q( key_c_r_31_41 ) );
  DFF_X1 key_c_r_reg_31_42 (.CK( clk ) , .D( key_c_r_30_42 ) , .Q( key_c_r_31_42 ) );
  DFF_X1 key_c_r_reg_31_43 (.CK( clk ) , .D( key_c_r_30_43 ) , .Q( key_c_r_31_43 ) );
  DFF_X1 key_c_r_reg_31_44 (.CK( clk ) , .D( key_c_r_30_44 ) , .Q( key_c_r_31_44 ) );
  DFF_X1 key_c_r_reg_31_45 (.CK( clk ) , .D( key_c_r_30_45 ) , .Q( key_c_r_31_45 ) );
  DFF_X1 key_c_r_reg_31_46 (.CK( clk ) , .D( key_c_r_30_46 ) , .Q( key_c_r_31_46 ) );
  DFF_X1 key_c_r_reg_31_47 (.CK( clk ) , .D( key_c_r_30_47 ) , .Q( key_c_r_31_47 ) );
  DFF_X1 key_c_r_reg_31_48 (.CK( clk ) , .D( key_c_r_30_48 ) , .Q( key_c_r_31_48 ) );
  DFF_X1 key_c_r_reg_31_49 (.CK( clk ) , .D( key_c_r_30_49 ) , .Q( key_c_r_31_49 ) );
  DFF_X1 key_c_r_reg_31_5 (.CK( clk ) , .D( key_c_r_30_5 ) , .Q( key_c_r_31_5 ) );
  DFF_X1 key_c_r_reg_31_50 (.CK( clk ) , .D( key_c_r_30_50 ) , .Q( key_c_r_31_50 ) );
  DFF_X1 key_c_r_reg_31_51 (.CK( clk ) , .D( key_c_r_30_51 ) , .Q( key_c_r_31_51 ) );
  DFF_X1 key_c_r_reg_31_52 (.CK( clk ) , .D( key_c_r_30_52 ) , .Q( key_c_r_31_52 ) );
  DFF_X1 key_c_r_reg_31_53 (.CK( clk ) , .D( key_c_r_30_53 ) , .Q( key_c_r_31_53 ) );
  DFF_X1 key_c_r_reg_31_54 (.CK( clk ) , .D( key_c_r_30_54 ) , .Q( key_c_r_31_54 ) );
  DFF_X1 key_c_r_reg_31_55 (.CK( clk ) , .D( key_c_r_30_55 ) , .Q( key_c_r_31_55 ) );
  DFF_X1 key_c_r_reg_31_6 (.CK( clk ) , .D( key_c_r_30_6 ) , .Q( key_c_r_31_6 ) );
  DFF_X1 key_c_r_reg_31_7 (.CK( clk ) , .D( key_c_r_30_7 ) , .Q( key_c_r_31_7 ) );
  DFF_X1 key_c_r_reg_31_8 (.CK( clk ) , .D( key_c_r_30_8 ) , .Q( key_c_r_31_8 ) );
  DFF_X1 key_c_r_reg_31_9 (.CK( clk ) , .D( key_c_r_30_9 ) , .Q( key_c_r_31_9 ) );
  DFF_X1 key_c_r_reg_32_0 (.CK( clk ) , .D( key_c_r_31_0 ) , .Q( key_c_r_32_0 ) );
  DFF_X1 key_c_r_reg_32_1 (.CK( clk ) , .D( key_c_r_31_1 ) , .Q( key_c_r_32_1 ) );
  DFF_X1 key_c_r_reg_32_10 (.CK( clk ) , .D( key_c_r_31_10 ) , .Q( key_c_r_32_10 ) );
  DFF_X1 key_c_r_reg_32_11 (.CK( clk ) , .D( key_c_r_31_11 ) , .Q( key_c_r_32_11 ) );
  DFF_X1 key_c_r_reg_32_12 (.CK( clk ) , .D( key_c_r_31_12 ) , .Q( key_c_r_32_12 ) );
  DFF_X1 key_c_r_reg_32_13 (.CK( clk ) , .D( key_c_r_31_13 ) , .Q( key_c_r_32_13 ) );
  DFF_X1 key_c_r_reg_32_14 (.CK( clk ) , .D( key_c_r_31_14 ) , .Q( key_c_r_32_14 ) );
  DFF_X1 key_c_r_reg_32_15 (.CK( clk ) , .D( key_c_r_31_15 ) , .Q( key_c_r_32_15 ) );
  DFF_X1 key_c_r_reg_32_16 (.CK( clk ) , .D( key_c_r_31_16 ) , .Q( key_c_r_32_16 ) );
  DFF_X1 key_c_r_reg_32_17 (.CK( clk ) , .D( key_c_r_31_17 ) , .Q( key_c_r_32_17 ) );
  DFF_X1 key_c_r_reg_32_18 (.CK( clk ) , .D( key_c_r_31_18 ) , .Q( key_c_r_32_18 ) );
  DFF_X1 key_c_r_reg_32_19 (.CK( clk ) , .D( key_c_r_31_19 ) , .Q( key_c_r_32_19 ) );
  DFF_X1 key_c_r_reg_32_2 (.CK( clk ) , .D( key_c_r_31_2 ) , .Q( key_c_r_32_2 ) );
  DFF_X1 key_c_r_reg_32_20 (.CK( clk ) , .D( key_c_r_31_20 ) , .Q( key_c_r_32_20 ) );
  DFF_X1 key_c_r_reg_32_21 (.CK( clk ) , .D( key_c_r_31_21 ) , .Q( key_c_r_32_21 ) );
  DFF_X1 key_c_r_reg_32_22 (.CK( clk ) , .D( key_c_r_31_22 ) , .Q( key_c_r_32_22 ) );
  DFF_X1 key_c_r_reg_32_23 (.CK( clk ) , .D( key_c_r_31_23 ) , .Q( key_c_r_32_23 ) );
  DFF_X1 key_c_r_reg_32_24 (.CK( clk ) , .D( key_c_r_31_24 ) , .Q( key_c_r_32_24 ) );
  DFF_X1 key_c_r_reg_32_25 (.CK( clk ) , .D( key_c_r_31_25 ) , .Q( key_c_r_32_25 ) );
  DFF_X1 key_c_r_reg_32_26 (.CK( clk ) , .D( key_c_r_31_26 ) , .Q( key_c_r_32_26 ) );
  DFF_X1 key_c_r_reg_32_27 (.CK( clk ) , .D( key_c_r_31_27 ) , .Q( key_c_r_32_27 ) );
  DFF_X1 key_c_r_reg_32_28 (.CK( clk ) , .D( key_c_r_31_28 ) , .Q( key_c_r_32_28 ) );
  DFF_X1 key_c_r_reg_32_29 (.CK( clk ) , .D( key_c_r_31_29 ) , .Q( key_c_r_32_29 ) );
  DFF_X1 key_c_r_reg_32_3 (.CK( clk ) , .D( key_c_r_31_3 ) , .Q( key_c_r_32_3 ) );
  DFF_X1 key_c_r_reg_32_30 (.CK( clk ) , .D( key_c_r_31_30 ) , .Q( key_c_r_32_30 ) );
  DFF_X1 key_c_r_reg_32_31 (.CK( clk ) , .D( key_c_r_31_31 ) , .Q( key_c_r_32_31 ) );
  DFF_X1 key_c_r_reg_32_32 (.CK( clk ) , .D( key_c_r_31_32 ) , .Q( key_c_r_32_32 ) );
  DFF_X1 key_c_r_reg_32_33 (.CK( clk ) , .D( key_c_r_31_33 ) , .Q( key_c_r_32_33 ) );
  DFF_X1 key_c_r_reg_32_34 (.CK( clk ) , .D( key_c_r_31_34 ) , .Q( key_c_r_32_34 ) );
  DFF_X1 key_c_r_reg_32_35 (.CK( clk ) , .D( key_c_r_31_35 ) , .Q( key_c_r_32_35 ) );
  DFF_X1 key_c_r_reg_32_36 (.CK( clk ) , .D( key_c_r_31_36 ) , .Q( key_c_r_32_36 ) );
  DFF_X1 key_c_r_reg_32_37 (.CK( clk ) , .D( key_c_r_31_37 ) , .Q( key_c_r_32_37 ) );
  DFF_X1 key_c_r_reg_32_38 (.CK( clk ) , .D( key_c_r_31_38 ) , .Q( key_c_r_32_38 ) );
  DFF_X1 key_c_r_reg_32_39 (.CK( clk ) , .D( key_c_r_31_39 ) , .Q( key_c_r_32_39 ) );
  DFF_X1 key_c_r_reg_32_4 (.CK( clk ) , .D( key_c_r_31_4 ) , .Q( key_c_r_32_4 ) );
  DFF_X1 key_c_r_reg_32_40 (.CK( clk ) , .D( key_c_r_31_40 ) , .Q( key_c_r_32_40 ) );
  DFF_X1 key_c_r_reg_32_41 (.CK( clk ) , .D( key_c_r_31_41 ) , .Q( key_c_r_32_41 ) );
  DFF_X1 key_c_r_reg_32_42 (.CK( clk ) , .D( key_c_r_31_42 ) , .Q( key_c_r_32_42 ) );
  DFF_X1 key_c_r_reg_32_43 (.CK( clk ) , .D( key_c_r_31_43 ) , .Q( key_c_r_32_43 ) );
  DFF_X1 key_c_r_reg_32_44 (.CK( clk ) , .D( key_c_r_31_44 ) , .Q( key_c_r_32_44 ) );
  DFF_X1 key_c_r_reg_32_45 (.CK( clk ) , .D( key_c_r_31_45 ) , .Q( key_c_r_32_45 ) );
  DFF_X1 key_c_r_reg_32_46 (.CK( clk ) , .D( key_c_r_31_46 ) , .Q( key_c_r_32_46 ) );
  DFF_X1 key_c_r_reg_32_47 (.CK( clk ) , .D( key_c_r_31_47 ) , .Q( key_c_r_32_47 ) );
  DFF_X1 key_c_r_reg_32_48 (.CK( clk ) , .D( key_c_r_31_48 ) , .Q( key_c_r_32_48 ) );
  DFF_X1 key_c_r_reg_32_49 (.CK( clk ) , .D( key_c_r_31_49 ) , .Q( key_c_r_32_49 ) );
  DFF_X1 key_c_r_reg_32_5 (.CK( clk ) , .D( key_c_r_31_5 ) , .Q( key_c_r_32_5 ) );
  DFF_X1 key_c_r_reg_32_50 (.CK( clk ) , .D( key_c_r_31_50 ) , .Q( key_c_r_32_50 ) );
  DFF_X1 key_c_r_reg_32_51 (.CK( clk ) , .D( key_c_r_31_51 ) , .Q( key_c_r_32_51 ) );
  DFF_X1 key_c_r_reg_32_52 (.CK( clk ) , .D( key_c_r_31_52 ) , .Q( key_c_r_32_52 ) );
  DFF_X1 key_c_r_reg_32_53 (.CK( clk ) , .D( key_c_r_31_53 ) , .Q( key_c_r_32_53 ) );
  DFF_X1 key_c_r_reg_32_54 (.CK( clk ) , .D( key_c_r_31_54 ) , .Q( key_c_r_32_54 ) );
  DFF_X1 key_c_r_reg_32_55 (.CK( clk ) , .D( key_c_r_31_55 ) , .Q( key_c_r_32_55 ) );
  DFF_X1 key_c_r_reg_32_6 (.CK( clk ) , .D( key_c_r_31_6 ) , .Q( key_c_r_32_6 ) );
  DFF_X1 key_c_r_reg_32_7 (.CK( clk ) , .D( key_c_r_31_7 ) , .Q( key_c_r_32_7 ) );
  DFF_X1 key_c_r_reg_32_8 (.CK( clk ) , .D( key_c_r_31_8 ) , .Q( key_c_r_32_8 ) );
  DFF_X1 key_c_r_reg_32_9 (.CK( clk ) , .D( key_c_r_31_9 ) , .Q( key_c_r_32_9 ) );
  DFF_X1 key_c_r_reg_33_0 (.CK( clk ) , .D( key_c_r_32_0 ) , .Q( key_c_r_33_0 ) );
  DFF_X1 key_c_r_reg_33_1 (.CK( clk ) , .D( key_c_r_32_1 ) , .Q( key_c_r_33_1 ) );
  DFF_X1 key_c_r_reg_33_10 (.CK( clk ) , .D( key_c_r_32_10 ) , .Q( key_c_r_33_10 ) );
  DFF_X1 key_c_r_reg_33_11 (.CK( clk ) , .D( key_c_r_32_11 ) , .Q( key_c_r_33_11 ) );
  DFF_X1 key_c_r_reg_33_12 (.CK( clk ) , .D( key_c_r_32_12 ) , .Q( key_c_r_33_12 ) );
  DFF_X1 key_c_r_reg_33_13 (.CK( clk ) , .D( key_c_r_32_13 ) , .Q( key_c_r_33_13 ) );
  DFF_X1 key_c_r_reg_33_14 (.CK( clk ) , .D( key_c_r_32_14 ) , .Q( key_c_r_33_14 ) );
  DFF_X1 key_c_r_reg_33_15 (.CK( clk ) , .D( key_c_r_32_15 ) , .Q( key_c_r_33_15 ) );
  DFF_X1 key_c_r_reg_33_16 (.CK( clk ) , .D( key_c_r_32_16 ) , .Q( key_c_r_33_16 ) );
  DFF_X1 key_c_r_reg_33_17 (.CK( clk ) , .D( key_c_r_32_17 ) , .Q( key_c_r_33_17 ) );
  DFF_X1 key_c_r_reg_33_18 (.CK( clk ) , .D( key_c_r_32_18 ) , .Q( key_c_r_33_18 ) );
  DFF_X1 key_c_r_reg_33_19 (.CK( clk ) , .D( key_c_r_32_19 ) , .Q( key_c_r_33_19 ) );
  DFF_X1 key_c_r_reg_33_2 (.CK( clk ) , .D( key_c_r_32_2 ) , .Q( key_c_r_33_2 ) );
  DFF_X1 key_c_r_reg_33_20 (.CK( clk ) , .D( key_c_r_32_20 ) , .Q( key_c_r_33_20 ) );
  DFF_X1 key_c_r_reg_33_21 (.CK( clk ) , .D( key_c_r_32_21 ) , .Q( key_c_r_33_21 ) );
  DFF_X1 key_c_r_reg_33_22 (.CK( clk ) , .D( key_c_r_32_22 ) , .Q( key_c_r_33_22 ) );
  DFF_X1 key_c_r_reg_33_23 (.CK( clk ) , .D( key_c_r_32_23 ) , .Q( key_c_r_33_23 ) );
  DFF_X1 key_c_r_reg_33_24 (.CK( clk ) , .D( key_c_r_32_24 ) , .Q( key_c_r_33_24 ) );
  DFF_X1 key_c_r_reg_33_25 (.CK( clk ) , .D( key_c_r_32_25 ) , .Q( key_c_r_33_25 ) );
  DFF_X1 key_c_r_reg_33_26 (.CK( clk ) , .D( key_c_r_32_26 ) , .Q( key_c_r_33_26 ) );
  DFF_X1 key_c_r_reg_33_27 (.CK( clk ) , .D( key_c_r_32_27 ) , .Q( key_c_r_33_27 ) );
  DFF_X1 key_c_r_reg_33_28 (.CK( clk ) , .D( key_c_r_32_28 ) , .Q( key_c_r_33_28 ) );
  DFF_X1 key_c_r_reg_33_29 (.CK( clk ) , .D( key_c_r_32_29 ) , .Q( key_c_r_33_29 ) );
  DFF_X1 key_c_r_reg_33_3 (.CK( clk ) , .D( key_c_r_32_3 ) , .Q( key_c_r_33_3 ) );
  DFF_X1 key_c_r_reg_33_30 (.CK( clk ) , .D( key_c_r_32_30 ) , .Q( key_c_r_33_30 ) );
  DFF_X1 key_c_r_reg_33_31 (.CK( clk ) , .D( key_c_r_32_31 ) , .Q( key_c_r_33_31 ) );
  DFF_X1 key_c_r_reg_33_32 (.CK( clk ) , .D( key_c_r_32_32 ) , .Q( key_c_r_33_32 ) );
  DFF_X1 key_c_r_reg_33_33 (.CK( clk ) , .D( key_c_r_32_33 ) , .Q( key_c_r_33_33 ) );
  DFF_X1 key_c_r_reg_33_34 (.CK( clk ) , .D( key_c_r_32_34 ) , .Q( key_c_r_33_34 ) );
  DFF_X1 key_c_r_reg_33_35 (.CK( clk ) , .D( key_c_r_32_35 ) , .Q( key_c_r_33_35 ) );
  DFF_X1 key_c_r_reg_33_36 (.CK( clk ) , .D( key_c_r_32_36 ) , .Q( key_c_r_33_36 ) );
  DFF_X1 key_c_r_reg_33_37 (.CK( clk ) , .D( key_c_r_32_37 ) , .Q( key_c_r_33_37 ) );
  DFF_X1 key_c_r_reg_33_38 (.CK( clk ) , .D( key_c_r_32_38 ) , .Q( key_c_r_33_38 ) );
  DFF_X1 key_c_r_reg_33_39 (.CK( clk ) , .D( key_c_r_32_39 ) , .Q( key_c_r_33_39 ) );
  DFF_X1 key_c_r_reg_33_4 (.CK( clk ) , .D( key_c_r_32_4 ) , .Q( key_c_r_33_4 ) );
  DFF_X1 key_c_r_reg_33_40 (.CK( clk ) , .D( key_c_r_32_40 ) , .Q( key_c_r_33_40 ) );
  DFF_X1 key_c_r_reg_33_41 (.CK( clk ) , .D( key_c_r_32_41 ) , .Q( key_c_r_33_41 ) );
  DFF_X1 key_c_r_reg_33_42 (.CK( clk ) , .D( key_c_r_32_42 ) , .Q( key_c_r_33_42 ) );
  DFF_X1 key_c_r_reg_33_43 (.CK( clk ) , .D( key_c_r_32_43 ) , .Q( key_c_r_33_43 ) );
  DFF_X1 key_c_r_reg_33_44 (.CK( clk ) , .D( key_c_r_32_44 ) , .Q( key_c_r_33_44 ) );
  DFF_X1 key_c_r_reg_33_45 (.CK( clk ) , .D( key_c_r_32_45 ) , .Q( key_c_r_33_45 ) );
  DFF_X1 key_c_r_reg_33_46 (.CK( clk ) , .D( key_c_r_32_46 ) , .Q( key_c_r_33_46 ) );
  DFF_X1 key_c_r_reg_33_47 (.CK( clk ) , .D( key_c_r_32_47 ) , .Q( key_c_r_33_47 ) );
  DFF_X1 key_c_r_reg_33_48 (.CK( clk ) , .D( key_c_r_32_48 ) , .Q( key_c_r_33_48 ) );
  DFF_X1 key_c_r_reg_33_49 (.CK( clk ) , .D( key_c_r_32_49 ) , .Q( key_c_r_33_49 ) );
  DFF_X1 key_c_r_reg_33_5 (.CK( clk ) , .D( key_c_r_32_5 ) , .Q( key_c_r_33_5 ) );
  DFF_X1 key_c_r_reg_33_50 (.CK( clk ) , .D( key_c_r_32_50 ) , .Q( key_c_r_33_50 ) );
  DFF_X1 key_c_r_reg_33_51 (.CK( clk ) , .D( key_c_r_32_51 ) , .Q( key_c_r_33_51 ) );
  DFF_X1 key_c_r_reg_33_52 (.CK( clk ) , .D( key_c_r_32_52 ) , .Q( key_c_r_33_52 ) );
  DFF_X1 key_c_r_reg_33_53 (.CK( clk ) , .D( key_c_r_32_53 ) , .Q( key_c_r_33_53 ) );
  DFF_X1 key_c_r_reg_33_54 (.CK( clk ) , .D( key_c_r_32_54 ) , .Q( key_c_r_33_54 ) );
  DFF_X1 key_c_r_reg_33_55 (.CK( clk ) , .D( key_c_r_32_55 ) , .Q( key_c_r_33_55 ) );
  DFF_X1 key_c_r_reg_33_6 (.CK( clk ) , .D( key_c_r_32_6 ) , .Q( key_c_r_33_6 ) );
  DFF_X1 key_c_r_reg_33_7 (.CK( clk ) , .D( key_c_r_32_7 ) , .Q( key_c_r_33_7 ) );
  DFF_X1 key_c_r_reg_33_8 (.CK( clk ) , .D( key_c_r_32_8 ) , .Q( key_c_r_33_8 ) );
  DFF_X1 key_c_r_reg_33_9 (.CK( clk ) , .D( key_c_r_32_9 ) , .Q( key_c_r_33_9 ) );
  DFF_X1 key_c_r_reg_3_0 (.CK( clk ) , .D( key_c_r_2_0 ) , .Q( key_c_r_3_0 ) );
  DFF_X1 key_c_r_reg_3_1 (.CK( clk ) , .D( key_c_r_2_1 ) , .Q( key_c_r_3_1 ) );
  DFF_X1 key_c_r_reg_3_10 (.CK( clk ) , .D( key_c_r_2_10 ) , .Q( key_c_r_3_10 ) );
  DFF_X1 key_c_r_reg_3_11 (.CK( clk ) , .D( key_c_r_2_11 ) , .Q( key_c_r_3_11 ) );
  DFF_X1 key_c_r_reg_3_12 (.CK( clk ) , .D( key_c_r_2_12 ) , .Q( key_c_r_3_12 ) );
  DFF_X1 key_c_r_reg_3_13 (.CK( clk ) , .D( key_c_r_2_13 ) , .Q( key_c_r_3_13 ) );
  DFF_X1 key_c_r_reg_3_14 (.CK( clk ) , .D( key_c_r_2_14 ) , .Q( key_c_r_3_14 ) );
  DFF_X1 key_c_r_reg_3_15 (.CK( clk ) , .D( key_c_r_2_15 ) , .Q( key_c_r_3_15 ) );
  DFF_X1 key_c_r_reg_3_16 (.CK( clk ) , .D( key_c_r_2_16 ) , .Q( key_c_r_3_16 ) );
  DFF_X1 key_c_r_reg_3_17 (.CK( clk ) , .D( key_c_r_2_17 ) , .Q( key_c_r_3_17 ) );
  DFF_X1 key_c_r_reg_3_18 (.CK( clk ) , .D( key_c_r_2_18 ) , .Q( key_c_r_3_18 ) );
  DFF_X1 key_c_r_reg_3_19 (.CK( clk ) , .D( key_c_r_2_19 ) , .Q( key_c_r_3_19 ) );
  DFF_X1 key_c_r_reg_3_2 (.CK( clk ) , .D( key_c_r_2_2 ) , .Q( key_c_r_3_2 ) );
  DFF_X1 key_c_r_reg_3_20 (.CK( clk ) , .D( key_c_r_2_20 ) , .Q( key_c_r_3_20 ) );
  DFF_X1 key_c_r_reg_3_21 (.CK( clk ) , .D( key_c_r_2_21 ) , .Q( key_c_r_3_21 ) );
  DFF_X1 key_c_r_reg_3_22 (.CK( clk ) , .D( key_c_r_2_22 ) , .Q( key_c_r_3_22 ) );
  DFF_X1 key_c_r_reg_3_23 (.CK( clk ) , .D( key_c_r_2_23 ) , .Q( key_c_r_3_23 ) );
  DFF_X1 key_c_r_reg_3_24 (.CK( clk ) , .D( key_c_r_2_24 ) , .Q( key_c_r_3_24 ) );
  DFF_X1 key_c_r_reg_3_25 (.CK( clk ) , .D( key_c_r_2_25 ) , .Q( key_c_r_3_25 ) );
  DFF_X1 key_c_r_reg_3_26 (.CK( clk ) , .D( key_c_r_2_26 ) , .Q( key_c_r_3_26 ) );
  DFF_X1 key_c_r_reg_3_27 (.CK( clk ) , .D( key_c_r_2_27 ) , .Q( key_c_r_3_27 ) );
  DFF_X1 key_c_r_reg_3_28 (.CK( clk ) , .D( key_c_r_2_28 ) , .Q( key_c_r_3_28 ) );
  DFF_X1 key_c_r_reg_3_29 (.CK( clk ) , .D( key_c_r_2_29 ) , .Q( key_c_r_3_29 ) );
  DFF_X1 key_c_r_reg_3_3 (.CK( clk ) , .D( key_c_r_2_3 ) , .Q( key_c_r_3_3 ) );
  DFF_X1 key_c_r_reg_3_30 (.CK( clk ) , .D( key_c_r_2_30 ) , .Q( key_c_r_3_30 ) );
  DFF_X1 key_c_r_reg_3_31 (.CK( clk ) , .D( key_c_r_2_31 ) , .Q( key_c_r_3_31 ) );
  DFF_X1 key_c_r_reg_3_32 (.CK( clk ) , .D( key_c_r_2_32 ) , .Q( key_c_r_3_32 ) );
  DFF_X1 key_c_r_reg_3_33 (.CK( clk ) , .D( key_c_r_2_33 ) , .Q( key_c_r_3_33 ) );
  DFF_X1 key_c_r_reg_3_34 (.CK( clk ) , .D( key_c_r_2_34 ) , .Q( key_c_r_3_34 ) );
  DFF_X1 key_c_r_reg_3_35 (.CK( clk ) , .D( key_c_r_2_35 ) , .Q( key_c_r_3_35 ) );
  DFF_X1 key_c_r_reg_3_36 (.CK( clk ) , .D( key_c_r_2_36 ) , .Q( key_c_r_3_36 ) );
  DFF_X1 key_c_r_reg_3_37 (.CK( clk ) , .D( key_c_r_2_37 ) , .Q( key_c_r_3_37 ) );
  DFF_X1 key_c_r_reg_3_38 (.CK( clk ) , .D( key_c_r_2_38 ) , .Q( key_c_r_3_38 ) );
  DFF_X1 key_c_r_reg_3_39 (.CK( clk ) , .D( key_c_r_2_39 ) , .Q( key_c_r_3_39 ) );
  DFF_X1 key_c_r_reg_3_4 (.CK( clk ) , .D( key_c_r_2_4 ) , .Q( key_c_r_3_4 ) );
  DFF_X1 key_c_r_reg_3_40 (.CK( clk ) , .D( key_c_r_2_40 ) , .Q( key_c_r_3_40 ) );
  DFF_X1 key_c_r_reg_3_41 (.CK( clk ) , .D( key_c_r_2_41 ) , .Q( key_c_r_3_41 ) );
  DFF_X1 key_c_r_reg_3_42 (.CK( clk ) , .D( key_c_r_2_42 ) , .Q( key_c_r_3_42 ) );
  DFF_X1 key_c_r_reg_3_43 (.CK( clk ) , .D( key_c_r_2_43 ) , .Q( key_c_r_3_43 ) );
  DFF_X1 key_c_r_reg_3_44 (.CK( clk ) , .D( key_c_r_2_44 ) , .Q( key_c_r_3_44 ) );
  DFF_X1 key_c_r_reg_3_45 (.CK( clk ) , .D( key_c_r_2_45 ) , .Q( key_c_r_3_45 ) );
  DFF_X1 key_c_r_reg_3_46 (.CK( clk ) , .D( key_c_r_2_46 ) , .Q( key_c_r_3_46 ) );
  DFF_X1 key_c_r_reg_3_47 (.CK( clk ) , .D( key_c_r_2_47 ) , .Q( key_c_r_3_47 ) );
  DFF_X1 key_c_r_reg_3_48 (.CK( clk ) , .D( key_c_r_2_48 ) , .Q( key_c_r_3_48 ) );
  DFF_X1 key_c_r_reg_3_49 (.CK( clk ) , .D( key_c_r_2_49 ) , .Q( key_c_r_3_49 ) );
  DFF_X1 key_c_r_reg_3_5 (.CK( clk ) , .D( key_c_r_2_5 ) , .Q( key_c_r_3_5 ) );
  DFF_X1 key_c_r_reg_3_50 (.CK( clk ) , .D( key_c_r_2_50 ) , .Q( key_c_r_3_50 ) );
  DFF_X1 key_c_r_reg_3_51 (.CK( clk ) , .D( key_c_r_2_51 ) , .Q( key_c_r_3_51 ) );
  DFF_X1 key_c_r_reg_3_52 (.CK( clk ) , .D( key_c_r_2_52 ) , .Q( key_c_r_3_52 ) );
  DFF_X1 key_c_r_reg_3_53 (.CK( clk ) , .D( key_c_r_2_53 ) , .Q( key_c_r_3_53 ) );
  DFF_X1 key_c_r_reg_3_54 (.CK( clk ) , .D( key_c_r_2_54 ) , .Q( key_c_r_3_54 ) );
  DFF_X1 key_c_r_reg_3_55 (.CK( clk ) , .D( key_c_r_2_55 ) , .Q( key_c_r_3_55 ) );
  DFF_X1 key_c_r_reg_3_6 (.CK( clk ) , .D( key_c_r_2_6 ) , .Q( key_c_r_3_6 ) );
  DFF_X1 key_c_r_reg_3_7 (.CK( clk ) , .D( key_c_r_2_7 ) , .Q( key_c_r_3_7 ) );
  DFF_X1 key_c_r_reg_3_8 (.CK( clk ) , .D( key_c_r_2_8 ) , .Q( key_c_r_3_8 ) );
  DFF_X1 key_c_r_reg_3_9 (.CK( clk ) , .D( key_c_r_2_9 ) , .Q( key_c_r_3_9 ) );
  DFF_X1 key_c_r_reg_4_0 (.CK( clk ) , .D( key_c_r_3_0 ) , .Q( key_c_r_4_0 ) );
  DFF_X1 key_c_r_reg_4_1 (.CK( clk ) , .D( key_c_r_3_1 ) , .Q( key_c_r_4_1 ) );
  DFF_X1 key_c_r_reg_4_10 (.CK( clk ) , .D( key_c_r_3_10 ) , .Q( key_c_r_4_10 ) );
  DFF_X1 key_c_r_reg_4_11 (.CK( clk ) , .D( key_c_r_3_11 ) , .Q( key_c_r_4_11 ) );
  DFF_X1 key_c_r_reg_4_12 (.CK( clk ) , .D( key_c_r_3_12 ) , .Q( key_c_r_4_12 ) );
  DFF_X1 key_c_r_reg_4_13 (.CK( clk ) , .D( key_c_r_3_13 ) , .Q( key_c_r_4_13 ) );
  DFF_X1 key_c_r_reg_4_14 (.CK( clk ) , .D( key_c_r_3_14 ) , .Q( key_c_r_4_14 ) );
  DFF_X1 key_c_r_reg_4_15 (.CK( clk ) , .D( key_c_r_3_15 ) , .Q( key_c_r_4_15 ) );
  DFF_X1 key_c_r_reg_4_16 (.CK( clk ) , .D( key_c_r_3_16 ) , .Q( key_c_r_4_16 ) );
  DFF_X1 key_c_r_reg_4_17 (.CK( clk ) , .D( key_c_r_3_17 ) , .Q( key_c_r_4_17 ) );
  DFF_X1 key_c_r_reg_4_18 (.CK( clk ) , .D( key_c_r_3_18 ) , .Q( key_c_r_4_18 ) );
  DFF_X1 key_c_r_reg_4_19 (.CK( clk ) , .D( key_c_r_3_19 ) , .Q( key_c_r_4_19 ) );
  DFF_X1 key_c_r_reg_4_2 (.CK( clk ) , .D( key_c_r_3_2 ) , .Q( key_c_r_4_2 ) );
  DFF_X1 key_c_r_reg_4_20 (.CK( clk ) , .D( key_c_r_3_20 ) , .Q( key_c_r_4_20 ) );
  DFF_X1 key_c_r_reg_4_21 (.CK( clk ) , .D( key_c_r_3_21 ) , .Q( key_c_r_4_21 ) );
  DFF_X1 key_c_r_reg_4_22 (.CK( clk ) , .D( key_c_r_3_22 ) , .Q( key_c_r_4_22 ) );
  DFF_X1 key_c_r_reg_4_23 (.CK( clk ) , .D( key_c_r_3_23 ) , .Q( key_c_r_4_23 ) );
  DFF_X1 key_c_r_reg_4_24 (.CK( clk ) , .D( key_c_r_3_24 ) , .Q( key_c_r_4_24 ) );
  DFF_X1 key_c_r_reg_4_25 (.CK( clk ) , .D( key_c_r_3_25 ) , .Q( key_c_r_4_25 ) );
  DFF_X1 key_c_r_reg_4_26 (.CK( clk ) , .D( key_c_r_3_26 ) , .Q( key_c_r_4_26 ) );
  DFF_X1 key_c_r_reg_4_27 (.CK( clk ) , .D( key_c_r_3_27 ) , .Q( key_c_r_4_27 ) );
  DFF_X1 key_c_r_reg_4_28 (.CK( clk ) , .D( key_c_r_3_28 ) , .Q( key_c_r_4_28 ) );
  DFF_X1 key_c_r_reg_4_29 (.CK( clk ) , .D( key_c_r_3_29 ) , .Q( key_c_r_4_29 ) );
  DFF_X1 key_c_r_reg_4_3 (.CK( clk ) , .D( key_c_r_3_3 ) , .Q( key_c_r_4_3 ) );
  DFF_X1 key_c_r_reg_4_30 (.CK( clk ) , .D( key_c_r_3_30 ) , .Q( key_c_r_4_30 ) );
  DFF_X1 key_c_r_reg_4_31 (.CK( clk ) , .D( key_c_r_3_31 ) , .Q( key_c_r_4_31 ) );
  DFF_X1 key_c_r_reg_4_32 (.CK( clk ) , .D( key_c_r_3_32 ) , .Q( key_c_r_4_32 ) );
  DFF_X1 key_c_r_reg_4_33 (.CK( clk ) , .D( key_c_r_3_33 ) , .Q( key_c_r_4_33 ) );
  DFF_X1 key_c_r_reg_4_34 (.CK( clk ) , .D( key_c_r_3_34 ) , .Q( key_c_r_4_34 ) );
  DFF_X1 key_c_r_reg_4_35 (.CK( clk ) , .D( key_c_r_3_35 ) , .Q( key_c_r_4_35 ) );
  DFF_X1 key_c_r_reg_4_36 (.CK( clk ) , .D( key_c_r_3_36 ) , .Q( key_c_r_4_36 ) );
  DFF_X1 key_c_r_reg_4_37 (.CK( clk ) , .D( key_c_r_3_37 ) , .Q( key_c_r_4_37 ) );
  DFF_X1 key_c_r_reg_4_38 (.CK( clk ) , .D( key_c_r_3_38 ) , .Q( key_c_r_4_38 ) );
  DFF_X1 key_c_r_reg_4_39 (.CK( clk ) , .D( key_c_r_3_39 ) , .Q( key_c_r_4_39 ) );
  DFF_X1 key_c_r_reg_4_4 (.CK( clk ) , .D( key_c_r_3_4 ) , .Q( key_c_r_4_4 ) );
  DFF_X1 key_c_r_reg_4_40 (.CK( clk ) , .D( key_c_r_3_40 ) , .Q( key_c_r_4_40 ) );
  DFF_X1 key_c_r_reg_4_41 (.CK( clk ) , .D( key_c_r_3_41 ) , .Q( key_c_r_4_41 ) );
  DFF_X1 key_c_r_reg_4_42 (.CK( clk ) , .D( key_c_r_3_42 ) , .Q( key_c_r_4_42 ) );
  DFF_X1 key_c_r_reg_4_43 (.CK( clk ) , .D( key_c_r_3_43 ) , .Q( key_c_r_4_43 ) );
  DFF_X1 key_c_r_reg_4_44 (.CK( clk ) , .D( key_c_r_3_44 ) , .Q( key_c_r_4_44 ) );
  DFF_X1 key_c_r_reg_4_45 (.CK( clk ) , .D( key_c_r_3_45 ) , .Q( key_c_r_4_45 ) );
  DFF_X1 key_c_r_reg_4_46 (.CK( clk ) , .D( key_c_r_3_46 ) , .Q( key_c_r_4_46 ) );
  DFF_X1 key_c_r_reg_4_47 (.CK( clk ) , .D( key_c_r_3_47 ) , .Q( key_c_r_4_47 ) );
  DFF_X1 key_c_r_reg_4_48 (.CK( clk ) , .D( key_c_r_3_48 ) , .Q( key_c_r_4_48 ) );
  DFF_X1 key_c_r_reg_4_49 (.CK( clk ) , .D( key_c_r_3_49 ) , .Q( key_c_r_4_49 ) );
  DFF_X1 key_c_r_reg_4_5 (.CK( clk ) , .D( key_c_r_3_5 ) , .Q( key_c_r_4_5 ) );
  DFF_X1 key_c_r_reg_4_50 (.CK( clk ) , .D( key_c_r_3_50 ) , .Q( key_c_r_4_50 ) );
  DFF_X1 key_c_r_reg_4_51 (.CK( clk ) , .D( key_c_r_3_51 ) , .Q( key_c_r_4_51 ) );
  DFF_X1 key_c_r_reg_4_52 (.CK( clk ) , .D( key_c_r_3_52 ) , .Q( key_c_r_4_52 ) );
  DFF_X1 key_c_r_reg_4_53 (.CK( clk ) , .D( key_c_r_3_53 ) , .Q( key_c_r_4_53 ) );
  DFF_X1 key_c_r_reg_4_54 (.CK( clk ) , .D( key_c_r_3_54 ) , .Q( key_c_r_4_54 ) );
  DFF_X1 key_c_r_reg_4_55 (.CK( clk ) , .D( key_c_r_3_55 ) , .Q( key_c_r_4_55 ) );
  DFF_X1 key_c_r_reg_4_6 (.CK( clk ) , .D( key_c_r_3_6 ) , .Q( key_c_r_4_6 ) );
  DFF_X1 key_c_r_reg_4_7 (.CK( clk ) , .D( key_c_r_3_7 ) , .Q( key_c_r_4_7 ) );
  DFF_X1 key_c_r_reg_4_8 (.CK( clk ) , .D( key_c_r_3_8 ) , .Q( key_c_r_4_8 ) );
  DFF_X1 key_c_r_reg_4_9 (.CK( clk ) , .D( key_c_r_3_9 ) , .Q( key_c_r_4_9 ) );
  DFF_X1 key_c_r_reg_5_0 (.CK( clk ) , .D( key_c_r_4_0 ) , .Q( key_c_r_5_0 ) );
  DFF_X1 key_c_r_reg_5_1 (.CK( clk ) , .D( key_c_r_4_1 ) , .Q( key_c_r_5_1 ) );
  DFF_X1 key_c_r_reg_5_10 (.CK( clk ) , .D( key_c_r_4_10 ) , .Q( key_c_r_5_10 ) );
  DFF_X1 key_c_r_reg_5_11 (.CK( clk ) , .D( key_c_r_4_11 ) , .Q( key_c_r_5_11 ) );
  DFF_X1 key_c_r_reg_5_12 (.CK( clk ) , .D( key_c_r_4_12 ) , .Q( key_c_r_5_12 ) );
  DFF_X1 key_c_r_reg_5_13 (.CK( clk ) , .D( key_c_r_4_13 ) , .Q( key_c_r_5_13 ) );
  DFF_X1 key_c_r_reg_5_14 (.CK( clk ) , .D( key_c_r_4_14 ) , .Q( key_c_r_5_14 ) );
  DFF_X1 key_c_r_reg_5_15 (.CK( clk ) , .D( key_c_r_4_15 ) , .Q( key_c_r_5_15 ) );
  DFF_X1 key_c_r_reg_5_16 (.CK( clk ) , .D( key_c_r_4_16 ) , .Q( key_c_r_5_16 ) );
  DFF_X1 key_c_r_reg_5_17 (.CK( clk ) , .D( key_c_r_4_17 ) , .Q( key_c_r_5_17 ) );
  DFF_X1 key_c_r_reg_5_18 (.CK( clk ) , .D( key_c_r_4_18 ) , .Q( key_c_r_5_18 ) );
  DFF_X1 key_c_r_reg_5_19 (.CK( clk ) , .D( key_c_r_4_19 ) , .Q( key_c_r_5_19 ) );
  DFF_X1 key_c_r_reg_5_2 (.CK( clk ) , .D( key_c_r_4_2 ) , .Q( key_c_r_5_2 ) );
  DFF_X1 key_c_r_reg_5_20 (.CK( clk ) , .D( key_c_r_4_20 ) , .Q( key_c_r_5_20 ) );
  DFF_X1 key_c_r_reg_5_21 (.CK( clk ) , .D( key_c_r_4_21 ) , .Q( key_c_r_5_21 ) );
  DFF_X1 key_c_r_reg_5_22 (.CK( clk ) , .D( key_c_r_4_22 ) , .Q( key_c_r_5_22 ) );
  DFF_X1 key_c_r_reg_5_23 (.CK( clk ) , .D( key_c_r_4_23 ) , .Q( key_c_r_5_23 ) );
  DFF_X1 key_c_r_reg_5_24 (.CK( clk ) , .D( key_c_r_4_24 ) , .Q( key_c_r_5_24 ) );
  DFF_X1 key_c_r_reg_5_25 (.CK( clk ) , .D( key_c_r_4_25 ) , .Q( key_c_r_5_25 ) );
  DFF_X1 key_c_r_reg_5_26 (.CK( clk ) , .D( key_c_r_4_26 ) , .Q( key_c_r_5_26 ) );
  DFF_X1 key_c_r_reg_5_27 (.CK( clk ) , .D( key_c_r_4_27 ) , .Q( key_c_r_5_27 ) );
  DFF_X1 key_c_r_reg_5_28 (.CK( clk ) , .D( key_c_r_4_28 ) , .Q( key_c_r_5_28 ) );
  DFF_X1 key_c_r_reg_5_29 (.CK( clk ) , .D( key_c_r_4_29 ) , .Q( key_c_r_5_29 ) );
  DFF_X1 key_c_r_reg_5_3 (.CK( clk ) , .D( key_c_r_4_3 ) , .Q( key_c_r_5_3 ) );
  DFF_X1 key_c_r_reg_5_30 (.CK( clk ) , .D( key_c_r_4_30 ) , .Q( key_c_r_5_30 ) );
  DFF_X1 key_c_r_reg_5_31 (.CK( clk ) , .D( key_c_r_4_31 ) , .Q( key_c_r_5_31 ) );
  DFF_X1 key_c_r_reg_5_32 (.CK( clk ) , .D( key_c_r_4_32 ) , .Q( key_c_r_5_32 ) );
  DFF_X1 key_c_r_reg_5_33 (.CK( clk ) , .D( key_c_r_4_33 ) , .Q( key_c_r_5_33 ) );
  DFF_X1 key_c_r_reg_5_34 (.CK( clk ) , .D( key_c_r_4_34 ) , .Q( key_c_r_5_34 ) );
  DFF_X1 key_c_r_reg_5_35 (.CK( clk ) , .D( key_c_r_4_35 ) , .Q( key_c_r_5_35 ) );
  DFF_X1 key_c_r_reg_5_36 (.CK( clk ) , .D( key_c_r_4_36 ) , .Q( key_c_r_5_36 ) );
  DFF_X1 key_c_r_reg_5_37 (.CK( clk ) , .D( key_c_r_4_37 ) , .Q( key_c_r_5_37 ) );
  DFF_X1 key_c_r_reg_5_38 (.CK( clk ) , .D( key_c_r_4_38 ) , .Q( key_c_r_5_38 ) );
  DFF_X1 key_c_r_reg_5_39 (.CK( clk ) , .D( key_c_r_4_39 ) , .Q( key_c_r_5_39 ) );
  DFF_X1 key_c_r_reg_5_4 (.CK( clk ) , .D( key_c_r_4_4 ) , .Q( key_c_r_5_4 ) );
  DFF_X1 key_c_r_reg_5_40 (.CK( clk ) , .D( key_c_r_4_40 ) , .Q( key_c_r_5_40 ) );
  DFF_X1 key_c_r_reg_5_41 (.CK( clk ) , .D( key_c_r_4_41 ) , .Q( key_c_r_5_41 ) );
  DFF_X1 key_c_r_reg_5_42 (.CK( clk ) , .D( key_c_r_4_42 ) , .Q( key_c_r_5_42 ) );
  DFF_X1 key_c_r_reg_5_43 (.CK( clk ) , .D( key_c_r_4_43 ) , .Q( key_c_r_5_43 ) );
  DFF_X1 key_c_r_reg_5_44 (.CK( clk ) , .D( key_c_r_4_44 ) , .Q( key_c_r_5_44 ) );
  DFF_X1 key_c_r_reg_5_45 (.CK( clk ) , .D( key_c_r_4_45 ) , .Q( key_c_r_5_45 ) );
  DFF_X1 key_c_r_reg_5_46 (.CK( clk ) , .D( key_c_r_4_46 ) , .Q( key_c_r_5_46 ) );
  DFF_X1 key_c_r_reg_5_47 (.CK( clk ) , .D( key_c_r_4_47 ) , .Q( key_c_r_5_47 ) );
  DFF_X1 key_c_r_reg_5_48 (.CK( clk ) , .D( key_c_r_4_48 ) , .Q( key_c_r_5_48 ) );
  DFF_X1 key_c_r_reg_5_49 (.CK( clk ) , .D( key_c_r_4_49 ) , .Q( key_c_r_5_49 ) );
  DFF_X1 key_c_r_reg_5_5 (.CK( clk ) , .D( key_c_r_4_5 ) , .Q( key_c_r_5_5 ) );
  DFF_X1 key_c_r_reg_5_50 (.CK( clk ) , .D( key_c_r_4_50 ) , .Q( key_c_r_5_50 ) );
  DFF_X1 key_c_r_reg_5_51 (.CK( clk ) , .D( key_c_r_4_51 ) , .Q( key_c_r_5_51 ) );
  DFF_X1 key_c_r_reg_5_52 (.CK( clk ) , .D( key_c_r_4_52 ) , .Q( key_c_r_5_52 ) );
  DFF_X1 key_c_r_reg_5_53 (.CK( clk ) , .D( key_c_r_4_53 ) , .Q( key_c_r_5_53 ) );
  DFF_X1 key_c_r_reg_5_54 (.CK( clk ) , .D( key_c_r_4_54 ) , .Q( key_c_r_5_54 ) );
  DFF_X1 key_c_r_reg_5_55 (.CK( clk ) , .D( key_c_r_4_55 ) , .Q( key_c_r_5_55 ) );
  DFF_X1 key_c_r_reg_5_6 (.CK( clk ) , .D( key_c_r_4_6 ) , .Q( key_c_r_5_6 ) );
  DFF_X1 key_c_r_reg_5_7 (.CK( clk ) , .D( key_c_r_4_7 ) , .Q( key_c_r_5_7 ) );
  DFF_X1 key_c_r_reg_5_8 (.CK( clk ) , .D( key_c_r_4_8 ) , .Q( key_c_r_5_8 ) );
  DFF_X1 key_c_r_reg_5_9 (.CK( clk ) , .D( key_c_r_4_9 ) , .Q( key_c_r_5_9 ) );
  DFF_X1 key_c_r_reg_6_0 (.CK( clk ) , .D( key_c_r_5_0 ) , .Q( key_c_r_6_0 ) );
  DFF_X1 key_c_r_reg_6_1 (.CK( clk ) , .D( key_c_r_5_1 ) , .Q( key_c_r_6_1 ) );
  DFF_X1 key_c_r_reg_6_10 (.CK( clk ) , .D( key_c_r_5_10 ) , .Q( key_c_r_6_10 ) );
  DFF_X1 key_c_r_reg_6_11 (.CK( clk ) , .D( key_c_r_5_11 ) , .Q( key_c_r_6_11 ) );
  DFF_X1 key_c_r_reg_6_12 (.CK( clk ) , .D( key_c_r_5_12 ) , .Q( key_c_r_6_12 ) );
  DFF_X1 key_c_r_reg_6_13 (.CK( clk ) , .D( key_c_r_5_13 ) , .Q( key_c_r_6_13 ) );
  DFF_X1 key_c_r_reg_6_14 (.CK( clk ) , .D( key_c_r_5_14 ) , .Q( key_c_r_6_14 ) );
  DFF_X1 key_c_r_reg_6_15 (.CK( clk ) , .D( key_c_r_5_15 ) , .Q( key_c_r_6_15 ) );
  DFF_X1 key_c_r_reg_6_16 (.CK( clk ) , .D( key_c_r_5_16 ) , .Q( key_c_r_6_16 ) );
  DFF_X1 key_c_r_reg_6_17 (.CK( clk ) , .D( key_c_r_5_17 ) , .Q( key_c_r_6_17 ) );
  DFF_X1 key_c_r_reg_6_18 (.CK( clk ) , .D( key_c_r_5_18 ) , .Q( key_c_r_6_18 ) );
  DFF_X1 key_c_r_reg_6_19 (.CK( clk ) , .D( key_c_r_5_19 ) , .Q( key_c_r_6_19 ) );
  DFF_X1 key_c_r_reg_6_2 (.CK( clk ) , .D( key_c_r_5_2 ) , .Q( key_c_r_6_2 ) );
  DFF_X1 key_c_r_reg_6_20 (.CK( clk ) , .D( key_c_r_5_20 ) , .Q( key_c_r_6_20 ) );
  DFF_X1 key_c_r_reg_6_21 (.CK( clk ) , .D( key_c_r_5_21 ) , .Q( key_c_r_6_21 ) );
  DFF_X1 key_c_r_reg_6_22 (.CK( clk ) , .D( key_c_r_5_22 ) , .Q( key_c_r_6_22 ) );
  DFF_X1 key_c_r_reg_6_23 (.CK( clk ) , .D( key_c_r_5_23 ) , .Q( key_c_r_6_23 ) );
  DFF_X1 key_c_r_reg_6_24 (.CK( clk ) , .D( key_c_r_5_24 ) , .Q( key_c_r_6_24 ) );
  DFF_X1 key_c_r_reg_6_25 (.CK( clk ) , .D( key_c_r_5_25 ) , .Q( key_c_r_6_25 ) );
  DFF_X1 key_c_r_reg_6_26 (.CK( clk ) , .D( key_c_r_5_26 ) , .Q( key_c_r_6_26 ) );
  DFF_X1 key_c_r_reg_6_27 (.CK( clk ) , .D( key_c_r_5_27 ) , .Q( key_c_r_6_27 ) );
  DFF_X1 key_c_r_reg_6_28 (.CK( clk ) , .D( key_c_r_5_28 ) , .Q( key_c_r_6_28 ) );
  DFF_X1 key_c_r_reg_6_29 (.CK( clk ) , .D( key_c_r_5_29 ) , .Q( key_c_r_6_29 ) );
  DFF_X1 key_c_r_reg_6_3 (.CK( clk ) , .D( key_c_r_5_3 ) , .Q( key_c_r_6_3 ) );
  DFF_X1 key_c_r_reg_6_30 (.CK( clk ) , .D( key_c_r_5_30 ) , .Q( key_c_r_6_30 ) );
  DFF_X1 key_c_r_reg_6_31 (.CK( clk ) , .D( key_c_r_5_31 ) , .Q( key_c_r_6_31 ) );
  DFF_X1 key_c_r_reg_6_32 (.CK( clk ) , .D( key_c_r_5_32 ) , .Q( key_c_r_6_32 ) );
  DFF_X1 key_c_r_reg_6_33 (.CK( clk ) , .D( key_c_r_5_33 ) , .Q( key_c_r_6_33 ) );
  DFF_X1 key_c_r_reg_6_34 (.CK( clk ) , .D( key_c_r_5_34 ) , .Q( key_c_r_6_34 ) );
  DFF_X1 key_c_r_reg_6_35 (.CK( clk ) , .D( key_c_r_5_35 ) , .Q( key_c_r_6_35 ) );
  DFF_X1 key_c_r_reg_6_36 (.CK( clk ) , .D( key_c_r_5_36 ) , .Q( key_c_r_6_36 ) );
  DFF_X1 key_c_r_reg_6_37 (.CK( clk ) , .D( key_c_r_5_37 ) , .Q( key_c_r_6_37 ) );
  DFF_X1 key_c_r_reg_6_38 (.CK( clk ) , .D( key_c_r_5_38 ) , .Q( key_c_r_6_38 ) );
  DFF_X1 key_c_r_reg_6_39 (.CK( clk ) , .D( key_c_r_5_39 ) , .Q( key_c_r_6_39 ) );
  DFF_X1 key_c_r_reg_6_4 (.CK( clk ) , .D( key_c_r_5_4 ) , .Q( key_c_r_6_4 ) );
  DFF_X1 key_c_r_reg_6_40 (.CK( clk ) , .D( key_c_r_5_40 ) , .Q( key_c_r_6_40 ) );
  DFF_X1 key_c_r_reg_6_41 (.CK( clk ) , .D( key_c_r_5_41 ) , .Q( key_c_r_6_41 ) );
  DFF_X1 key_c_r_reg_6_42 (.CK( clk ) , .D( key_c_r_5_42 ) , .Q( key_c_r_6_42 ) );
  DFF_X1 key_c_r_reg_6_43 (.CK( clk ) , .D( key_c_r_5_43 ) , .Q( key_c_r_6_43 ) );
  DFF_X1 key_c_r_reg_6_44 (.CK( clk ) , .D( key_c_r_5_44 ) , .Q( key_c_r_6_44 ) );
  DFF_X1 key_c_r_reg_6_45 (.CK( clk ) , .D( key_c_r_5_45 ) , .Q( key_c_r_6_45 ) );
  DFF_X1 key_c_r_reg_6_46 (.CK( clk ) , .D( key_c_r_5_46 ) , .Q( key_c_r_6_46 ) );
  DFF_X1 key_c_r_reg_6_47 (.CK( clk ) , .D( key_c_r_5_47 ) , .Q( key_c_r_6_47 ) );
  DFF_X1 key_c_r_reg_6_48 (.CK( clk ) , .D( key_c_r_5_48 ) , .Q( key_c_r_6_48 ) );
  DFF_X1 key_c_r_reg_6_49 (.CK( clk ) , .D( key_c_r_5_49 ) , .Q( key_c_r_6_49 ) );
  DFF_X1 key_c_r_reg_6_5 (.CK( clk ) , .D( key_c_r_5_5 ) , .Q( key_c_r_6_5 ) );
  DFF_X1 key_c_r_reg_6_50 (.CK( clk ) , .D( key_c_r_5_50 ) , .Q( key_c_r_6_50 ) );
  DFF_X1 key_c_r_reg_6_51 (.CK( clk ) , .D( key_c_r_5_51 ) , .Q( key_c_r_6_51 ) );
  DFF_X1 key_c_r_reg_6_52 (.CK( clk ) , .D( key_c_r_5_52 ) , .Q( key_c_r_6_52 ) );
  DFF_X1 key_c_r_reg_6_53 (.CK( clk ) , .D( key_c_r_5_53 ) , .Q( key_c_r_6_53 ) );
  DFF_X1 key_c_r_reg_6_54 (.CK( clk ) , .D( key_c_r_5_54 ) , .Q( key_c_r_6_54 ) );
  DFF_X1 key_c_r_reg_6_55 (.CK( clk ) , .D( key_c_r_5_55 ) , .Q( key_c_r_6_55 ) );
  DFF_X1 key_c_r_reg_6_6 (.CK( clk ) , .D( key_c_r_5_6 ) , .Q( key_c_r_6_6 ) );
  DFF_X1 key_c_r_reg_6_7 (.CK( clk ) , .D( key_c_r_5_7 ) , .Q( key_c_r_6_7 ) );
  DFF_X1 key_c_r_reg_6_8 (.CK( clk ) , .D( key_c_r_5_8 ) , .Q( key_c_r_6_8 ) );
  DFF_X1 key_c_r_reg_6_9 (.CK( clk ) , .D( key_c_r_5_9 ) , .Q( key_c_r_6_9 ) );
  DFF_X1 key_c_r_reg_7_0 (.CK( clk ) , .D( key_c_r_6_0 ) , .Q( key_c_r_7_0 ) );
  DFF_X1 key_c_r_reg_7_1 (.CK( clk ) , .D( key_c_r_6_1 ) , .Q( key_c_r_7_1 ) );
  DFF_X1 key_c_r_reg_7_10 (.CK( clk ) , .D( key_c_r_6_10 ) , .Q( key_c_r_7_10 ) );
  DFF_X1 key_c_r_reg_7_11 (.CK( clk ) , .D( key_c_r_6_11 ) , .Q( key_c_r_7_11 ) );
  DFF_X1 key_c_r_reg_7_12 (.CK( clk ) , .D( key_c_r_6_12 ) , .Q( key_c_r_7_12 ) );
  DFF_X1 key_c_r_reg_7_13 (.CK( clk ) , .D( key_c_r_6_13 ) , .Q( key_c_r_7_13 ) );
  DFF_X1 key_c_r_reg_7_14 (.CK( clk ) , .D( key_c_r_6_14 ) , .Q( key_c_r_7_14 ) );
  DFF_X1 key_c_r_reg_7_15 (.CK( clk ) , .D( key_c_r_6_15 ) , .Q( key_c_r_7_15 ) );
  DFF_X1 key_c_r_reg_7_16 (.CK( clk ) , .D( key_c_r_6_16 ) , .Q( key_c_r_7_16 ) );
  DFF_X1 key_c_r_reg_7_17 (.CK( clk ) , .D( key_c_r_6_17 ) , .Q( key_c_r_7_17 ) );
  DFF_X1 key_c_r_reg_7_18 (.CK( clk ) , .D( key_c_r_6_18 ) , .Q( key_c_r_7_18 ) );
  DFF_X1 key_c_r_reg_7_19 (.CK( clk ) , .D( key_c_r_6_19 ) , .Q( key_c_r_7_19 ) );
  DFF_X1 key_c_r_reg_7_2 (.CK( clk ) , .D( key_c_r_6_2 ) , .Q( key_c_r_7_2 ) );
  DFF_X1 key_c_r_reg_7_20 (.CK( clk ) , .D( key_c_r_6_20 ) , .Q( key_c_r_7_20 ) );
  DFF_X1 key_c_r_reg_7_21 (.CK( clk ) , .D( key_c_r_6_21 ) , .Q( key_c_r_7_21 ) );
  DFF_X1 key_c_r_reg_7_22 (.CK( clk ) , .D( key_c_r_6_22 ) , .Q( key_c_r_7_22 ) );
  DFF_X1 key_c_r_reg_7_23 (.CK( clk ) , .D( key_c_r_6_23 ) , .Q( key_c_r_7_23 ) );
  DFF_X1 key_c_r_reg_7_24 (.CK( clk ) , .D( key_c_r_6_24 ) , .Q( key_c_r_7_24 ) );
  DFF_X1 key_c_r_reg_7_25 (.CK( clk ) , .D( key_c_r_6_25 ) , .Q( key_c_r_7_25 ) );
  DFF_X1 key_c_r_reg_7_26 (.CK( clk ) , .D( key_c_r_6_26 ) , .Q( key_c_r_7_26 ) );
  DFF_X1 key_c_r_reg_7_27 (.CK( clk ) , .D( key_c_r_6_27 ) , .Q( key_c_r_7_27 ) );
  DFF_X1 key_c_r_reg_7_28 (.CK( clk ) , .D( key_c_r_6_28 ) , .Q( key_c_r_7_28 ) );
  DFF_X1 key_c_r_reg_7_29 (.CK( clk ) , .D( key_c_r_6_29 ) , .Q( key_c_r_7_29 ) );
  DFF_X1 key_c_r_reg_7_3 (.CK( clk ) , .D( key_c_r_6_3 ) , .Q( key_c_r_7_3 ) );
  DFF_X1 key_c_r_reg_7_30 (.CK( clk ) , .D( key_c_r_6_30 ) , .Q( key_c_r_7_30 ) );
  DFF_X1 key_c_r_reg_7_31 (.CK( clk ) , .D( key_c_r_6_31 ) , .Q( key_c_r_7_31 ) );
  DFF_X1 key_c_r_reg_7_32 (.CK( clk ) , .D( key_c_r_6_32 ) , .Q( key_c_r_7_32 ) );
  DFF_X1 key_c_r_reg_7_33 (.CK( clk ) , .D( key_c_r_6_33 ) , .Q( key_c_r_7_33 ) );
  DFF_X1 key_c_r_reg_7_34 (.CK( clk ) , .D( key_c_r_6_34 ) , .Q( key_c_r_7_34 ) );
  DFF_X1 key_c_r_reg_7_35 (.CK( clk ) , .D( key_c_r_6_35 ) , .Q( key_c_r_7_35 ) );
  DFF_X1 key_c_r_reg_7_36 (.CK( clk ) , .D( key_c_r_6_36 ) , .Q( key_c_r_7_36 ) );
  DFF_X1 key_c_r_reg_7_37 (.CK( clk ) , .D( key_c_r_6_37 ) , .Q( key_c_r_7_37 ) );
  DFF_X1 key_c_r_reg_7_38 (.CK( clk ) , .D( key_c_r_6_38 ) , .Q( key_c_r_7_38 ) );
  DFF_X1 key_c_r_reg_7_39 (.CK( clk ) , .D( key_c_r_6_39 ) , .Q( key_c_r_7_39 ) );
  DFF_X1 key_c_r_reg_7_4 (.CK( clk ) , .D( key_c_r_6_4 ) , .Q( key_c_r_7_4 ) );
  DFF_X1 key_c_r_reg_7_40 (.CK( clk ) , .D( key_c_r_6_40 ) , .Q( key_c_r_7_40 ) );
  DFF_X1 key_c_r_reg_7_41 (.CK( clk ) , .D( key_c_r_6_41 ) , .Q( key_c_r_7_41 ) );
  DFF_X1 key_c_r_reg_7_42 (.CK( clk ) , .D( key_c_r_6_42 ) , .Q( key_c_r_7_42 ) );
  DFF_X1 key_c_r_reg_7_43 (.CK( clk ) , .D( key_c_r_6_43 ) , .Q( key_c_r_7_43 ) );
  DFF_X1 key_c_r_reg_7_44 (.CK( clk ) , .D( key_c_r_6_44 ) , .Q( key_c_r_7_44 ) );
  DFF_X1 key_c_r_reg_7_45 (.CK( clk ) , .D( key_c_r_6_45 ) , .Q( key_c_r_7_45 ) );
  DFF_X1 key_c_r_reg_7_46 (.CK( clk ) , .D( key_c_r_6_46 ) , .Q( key_c_r_7_46 ) );
  DFF_X1 key_c_r_reg_7_47 (.CK( clk ) , .D( key_c_r_6_47 ) , .Q( key_c_r_7_47 ) );
  DFF_X1 key_c_r_reg_7_48 (.CK( clk ) , .D( key_c_r_6_48 ) , .Q( key_c_r_7_48 ) );
  DFF_X1 key_c_r_reg_7_49 (.CK( clk ) , .D( key_c_r_6_49 ) , .Q( key_c_r_7_49 ) );
  DFF_X1 key_c_r_reg_7_5 (.CK( clk ) , .D( key_c_r_6_5 ) , .Q( key_c_r_7_5 ) );
  DFF_X1 key_c_r_reg_7_50 (.CK( clk ) , .D( key_c_r_6_50 ) , .Q( key_c_r_7_50 ) );
  DFF_X1 key_c_r_reg_7_51 (.CK( clk ) , .D( key_c_r_6_51 ) , .Q( key_c_r_7_51 ) );
  DFF_X1 key_c_r_reg_7_52 (.CK( clk ) , .D( key_c_r_6_52 ) , .Q( key_c_r_7_52 ) );
  DFF_X1 key_c_r_reg_7_53 (.CK( clk ) , .D( key_c_r_6_53 ) , .Q( key_c_r_7_53 ) );
  DFF_X1 key_c_r_reg_7_54 (.CK( clk ) , .D( key_c_r_6_54 ) , .Q( key_c_r_7_54 ) );
  DFF_X1 key_c_r_reg_7_55 (.CK( clk ) , .D( key_c_r_6_55 ) , .Q( key_c_r_7_55 ) );
  DFF_X1 key_c_r_reg_7_6 (.CK( clk ) , .D( key_c_r_6_6 ) , .Q( key_c_r_7_6 ) );
  DFF_X1 key_c_r_reg_7_7 (.CK( clk ) , .D( key_c_r_6_7 ) , .Q( key_c_r_7_7 ) );
  DFF_X1 key_c_r_reg_7_8 (.CK( clk ) , .D( key_c_r_6_8 ) , .Q( key_c_r_7_8 ) );
  DFF_X1 key_c_r_reg_7_9 (.CK( clk ) , .D( key_c_r_6_9 ) , .Q( key_c_r_7_9 ) );
  DFF_X1 key_c_r_reg_8_0 (.CK( clk ) , .D( key_c_r_7_0 ) , .Q( key_c_r_8_0 ) );
  DFF_X1 key_c_r_reg_8_1 (.CK( clk ) , .D( key_c_r_7_1 ) , .Q( key_c_r_8_1 ) );
  DFF_X1 key_c_r_reg_8_10 (.CK( clk ) , .D( key_c_r_7_10 ) , .Q( key_c_r_8_10 ) );
  DFF_X1 key_c_r_reg_8_11 (.CK( clk ) , .D( key_c_r_7_11 ) , .Q( key_c_r_8_11 ) );
  DFF_X1 key_c_r_reg_8_12 (.CK( clk ) , .D( key_c_r_7_12 ) , .Q( key_c_r_8_12 ) );
  DFF_X1 key_c_r_reg_8_13 (.CK( clk ) , .D( key_c_r_7_13 ) , .Q( key_c_r_8_13 ) );
  DFF_X1 key_c_r_reg_8_14 (.CK( clk ) , .D( key_c_r_7_14 ) , .Q( key_c_r_8_14 ) );
  DFF_X1 key_c_r_reg_8_15 (.CK( clk ) , .D( key_c_r_7_15 ) , .Q( key_c_r_8_15 ) );
  DFF_X1 key_c_r_reg_8_16 (.CK( clk ) , .D( key_c_r_7_16 ) , .Q( key_c_r_8_16 ) );
  DFF_X1 key_c_r_reg_8_17 (.CK( clk ) , .D( key_c_r_7_17 ) , .Q( key_c_r_8_17 ) );
  DFF_X1 key_c_r_reg_8_18 (.CK( clk ) , .D( key_c_r_7_18 ) , .Q( key_c_r_8_18 ) );
  DFF_X1 key_c_r_reg_8_19 (.CK( clk ) , .D( key_c_r_7_19 ) , .Q( key_c_r_8_19 ) );
  DFF_X1 key_c_r_reg_8_2 (.CK( clk ) , .D( key_c_r_7_2 ) , .Q( key_c_r_8_2 ) );
  DFF_X1 key_c_r_reg_8_20 (.CK( clk ) , .D( key_c_r_7_20 ) , .Q( key_c_r_8_20 ) );
  DFF_X1 key_c_r_reg_8_21 (.CK( clk ) , .D( key_c_r_7_21 ) , .Q( key_c_r_8_21 ) );
  DFF_X1 key_c_r_reg_8_22 (.CK( clk ) , .D( key_c_r_7_22 ) , .Q( key_c_r_8_22 ) );
  DFF_X1 key_c_r_reg_8_23 (.CK( clk ) , .D( key_c_r_7_23 ) , .Q( key_c_r_8_23 ) );
  DFF_X1 key_c_r_reg_8_24 (.CK( clk ) , .D( key_c_r_7_24 ) , .Q( key_c_r_8_24 ) );
  DFF_X1 key_c_r_reg_8_25 (.CK( clk ) , .D( key_c_r_7_25 ) , .Q( key_c_r_8_25 ) );
  DFF_X1 key_c_r_reg_8_26 (.CK( clk ) , .D( key_c_r_7_26 ) , .Q( key_c_r_8_26 ) );
  DFF_X1 key_c_r_reg_8_27 (.CK( clk ) , .D( key_c_r_7_27 ) , .Q( key_c_r_8_27 ) );
  DFF_X1 key_c_r_reg_8_28 (.CK( clk ) , .D( key_c_r_7_28 ) , .Q( key_c_r_8_28 ) );
  DFF_X1 key_c_r_reg_8_29 (.CK( clk ) , .D( key_c_r_7_29 ) , .Q( key_c_r_8_29 ) );
  DFF_X1 key_c_r_reg_8_3 (.CK( clk ) , .D( key_c_r_7_3 ) , .Q( key_c_r_8_3 ) );
  DFF_X1 key_c_r_reg_8_30 (.CK( clk ) , .D( key_c_r_7_30 ) , .Q( key_c_r_8_30 ) );
  DFF_X1 key_c_r_reg_8_31 (.CK( clk ) , .D( key_c_r_7_31 ) , .Q( key_c_r_8_31 ) );
  DFF_X1 key_c_r_reg_8_32 (.CK( clk ) , .D( key_c_r_7_32 ) , .Q( key_c_r_8_32 ) );
  DFF_X1 key_c_r_reg_8_33 (.CK( clk ) , .D( key_c_r_7_33 ) , .Q( key_c_r_8_33 ) );
  DFF_X1 key_c_r_reg_8_34 (.CK( clk ) , .D( key_c_r_7_34 ) , .Q( key_c_r_8_34 ) );
  DFF_X1 key_c_r_reg_8_35 (.CK( clk ) , .D( key_c_r_7_35 ) , .Q( key_c_r_8_35 ) );
  DFF_X1 key_c_r_reg_8_36 (.CK( clk ) , .D( key_c_r_7_36 ) , .Q( key_c_r_8_36 ) );
  DFF_X1 key_c_r_reg_8_37 (.CK( clk ) , .D( key_c_r_7_37 ) , .Q( key_c_r_8_37 ) );
  DFF_X1 key_c_r_reg_8_38 (.CK( clk ) , .D( key_c_r_7_38 ) , .Q( key_c_r_8_38 ) );
  DFF_X1 key_c_r_reg_8_39 (.CK( clk ) , .D( key_c_r_7_39 ) , .Q( key_c_r_8_39 ) );
  DFF_X1 key_c_r_reg_8_4 (.CK( clk ) , .D( key_c_r_7_4 ) , .Q( key_c_r_8_4 ) );
  DFF_X1 key_c_r_reg_8_40 (.CK( clk ) , .D( key_c_r_7_40 ) , .Q( key_c_r_8_40 ) );
  DFF_X1 key_c_r_reg_8_41 (.CK( clk ) , .D( key_c_r_7_41 ) , .Q( key_c_r_8_41 ) );
  DFF_X1 key_c_r_reg_8_42 (.CK( clk ) , .D( key_c_r_7_42 ) , .Q( key_c_r_8_42 ) );
  DFF_X1 key_c_r_reg_8_43 (.CK( clk ) , .D( key_c_r_7_43 ) , .Q( key_c_r_8_43 ) );
  DFF_X1 key_c_r_reg_8_44 (.CK( clk ) , .D( key_c_r_7_44 ) , .Q( key_c_r_8_44 ) );
  DFF_X1 key_c_r_reg_8_45 (.CK( clk ) , .D( key_c_r_7_45 ) , .Q( key_c_r_8_45 ) );
  DFF_X1 key_c_r_reg_8_46 (.CK( clk ) , .D( key_c_r_7_46 ) , .Q( key_c_r_8_46 ) );
  DFF_X1 key_c_r_reg_8_47 (.CK( clk ) , .D( key_c_r_7_47 ) , .Q( key_c_r_8_47 ) );
  DFF_X1 key_c_r_reg_8_48 (.CK( clk ) , .D( key_c_r_7_48 ) , .Q( key_c_r_8_48 ) );
  DFF_X1 key_c_r_reg_8_49 (.CK( clk ) , .D( key_c_r_7_49 ) , .Q( key_c_r_8_49 ) );
  DFF_X1 key_c_r_reg_8_5 (.CK( clk ) , .D( key_c_r_7_5 ) , .Q( key_c_r_8_5 ) );
  DFF_X1 key_c_r_reg_8_50 (.CK( clk ) , .D( key_c_r_7_50 ) , .Q( key_c_r_8_50 ) );
  DFF_X1 key_c_r_reg_8_51 (.CK( clk ) , .D( key_c_r_7_51 ) , .Q( key_c_r_8_51 ) );
  DFF_X1 key_c_r_reg_8_52 (.CK( clk ) , .D( key_c_r_7_52 ) , .Q( key_c_r_8_52 ) );
  DFF_X1 key_c_r_reg_8_53 (.CK( clk ) , .D( key_c_r_7_53 ) , .Q( key_c_r_8_53 ) );
  DFF_X1 key_c_r_reg_8_54 (.CK( clk ) , .D( key_c_r_7_54 ) , .Q( key_c_r_8_54 ) );
  DFF_X1 key_c_r_reg_8_55 (.CK( clk ) , .D( key_c_r_7_55 ) , .Q( key_c_r_8_55 ) );
  DFF_X1 key_c_r_reg_8_6 (.CK( clk ) , .D( key_c_r_7_6 ) , .Q( key_c_r_8_6 ) );
  DFF_X1 key_c_r_reg_8_7 (.CK( clk ) , .D( key_c_r_7_7 ) , .Q( key_c_r_8_7 ) );
  DFF_X1 key_c_r_reg_8_8 (.CK( clk ) , .D( key_c_r_7_8 ) , .Q( key_c_r_8_8 ) );
  DFF_X1 key_c_r_reg_8_9 (.CK( clk ) , .D( key_c_r_7_9 ) , .Q( key_c_r_8_9 ) );
  DFF_X1 key_c_r_reg_9_0 (.CK( clk ) , .D( key_c_r_8_0 ) , .Q( key_c_r_9_0 ) );
  DFF_X1 key_c_r_reg_9_1 (.CK( clk ) , .D( key_c_r_8_1 ) , .Q( key_c_r_9_1 ) );
  DFF_X1 key_c_r_reg_9_10 (.CK( clk ) , .D( key_c_r_8_10 ) , .Q( key_c_r_9_10 ) );
  DFF_X1 key_c_r_reg_9_11 (.CK( clk ) , .D( key_c_r_8_11 ) , .Q( key_c_r_9_11 ) );
  DFF_X1 key_c_r_reg_9_12 (.CK( clk ) , .D( key_c_r_8_12 ) , .Q( key_c_r_9_12 ) );
  DFF_X1 key_c_r_reg_9_13 (.CK( clk ) , .D( key_c_r_8_13 ) , .Q( key_c_r_9_13 ) );
  DFF_X1 key_c_r_reg_9_14 (.CK( clk ) , .D( key_c_r_8_14 ) , .Q( key_c_r_9_14 ) );
  DFF_X1 key_c_r_reg_9_15 (.CK( clk ) , .D( key_c_r_8_15 ) , .Q( key_c_r_9_15 ) );
  DFF_X1 key_c_r_reg_9_16 (.CK( clk ) , .D( key_c_r_8_16 ) , .Q( key_c_r_9_16 ) );
  DFF_X1 key_c_r_reg_9_17 (.CK( clk ) , .D( key_c_r_8_17 ) , .Q( key_c_r_9_17 ) );
  DFF_X1 key_c_r_reg_9_18 (.CK( clk ) , .D( key_c_r_8_18 ) , .Q( key_c_r_9_18 ) );
  DFF_X1 key_c_r_reg_9_19 (.CK( clk ) , .D( key_c_r_8_19 ) , .Q( key_c_r_9_19 ) );
  DFF_X1 key_c_r_reg_9_2 (.CK( clk ) , .D( key_c_r_8_2 ) , .Q( key_c_r_9_2 ) );
  DFF_X1 key_c_r_reg_9_20 (.CK( clk ) , .D( key_c_r_8_20 ) , .Q( key_c_r_9_20 ) );
  DFF_X1 key_c_r_reg_9_21 (.CK( clk ) , .D( key_c_r_8_21 ) , .Q( key_c_r_9_21 ) );
  DFF_X1 key_c_r_reg_9_22 (.CK( clk ) , .D( key_c_r_8_22 ) , .Q( key_c_r_9_22 ) );
  DFF_X1 key_c_r_reg_9_23 (.CK( clk ) , .D( key_c_r_8_23 ) , .Q( key_c_r_9_23 ) );
  DFF_X1 key_c_r_reg_9_24 (.CK( clk ) , .D( key_c_r_8_24 ) , .Q( key_c_r_9_24 ) );
  DFF_X1 key_c_r_reg_9_25 (.CK( clk ) , .D( key_c_r_8_25 ) , .Q( key_c_r_9_25 ) );
  DFF_X1 key_c_r_reg_9_26 (.CK( clk ) , .D( key_c_r_8_26 ) , .Q( key_c_r_9_26 ) );
  DFF_X1 key_c_r_reg_9_27 (.CK( clk ) , .D( key_c_r_8_27 ) , .Q( key_c_r_9_27 ) );
  DFF_X1 key_c_r_reg_9_28 (.CK( clk ) , .D( key_c_r_8_28 ) , .Q( key_c_r_9_28 ) );
  DFF_X1 key_c_r_reg_9_29 (.CK( clk ) , .D( key_c_r_8_29 ) , .Q( key_c_r_9_29 ) );
  DFF_X1 key_c_r_reg_9_3 (.CK( clk ) , .D( key_c_r_8_3 ) , .Q( key_c_r_9_3 ) );
  DFF_X1 key_c_r_reg_9_30 (.CK( clk ) , .D( key_c_r_8_30 ) , .Q( key_c_r_9_30 ) );
  DFF_X1 key_c_r_reg_9_31 (.CK( clk ) , .D( key_c_r_8_31 ) , .Q( key_c_r_9_31 ) );
  DFF_X1 key_c_r_reg_9_32 (.CK( clk ) , .D( key_c_r_8_32 ) , .Q( key_c_r_9_32 ) );
  DFF_X1 key_c_r_reg_9_33 (.CK( clk ) , .D( key_c_r_8_33 ) , .Q( key_c_r_9_33 ) );
  DFF_X1 key_c_r_reg_9_34 (.CK( clk ) , .D( key_c_r_8_34 ) , .Q( key_c_r_9_34 ) );
  DFF_X1 key_c_r_reg_9_35 (.CK( clk ) , .D( key_c_r_8_35 ) , .Q( key_c_r_9_35 ) );
  DFF_X1 key_c_r_reg_9_36 (.CK( clk ) , .D( key_c_r_8_36 ) , .Q( key_c_r_9_36 ) );
  DFF_X1 key_c_r_reg_9_37 (.CK( clk ) , .D( key_c_r_8_37 ) , .Q( key_c_r_9_37 ) );
  DFF_X1 key_c_r_reg_9_38 (.CK( clk ) , .D( key_c_r_8_38 ) , .Q( key_c_r_9_38 ) );
  DFF_X1 key_c_r_reg_9_39 (.CK( clk ) , .D( key_c_r_8_39 ) , .Q( key_c_r_9_39 ) );
  DFF_X1 key_c_r_reg_9_4 (.CK( clk ) , .D( key_c_r_8_4 ) , .Q( key_c_r_9_4 ) );
  DFF_X1 key_c_r_reg_9_40 (.CK( clk ) , .D( key_c_r_8_40 ) , .Q( key_c_r_9_40 ) );
  DFF_X1 key_c_r_reg_9_41 (.CK( clk ) , .D( key_c_r_8_41 ) , .Q( key_c_r_9_41 ) );
  DFF_X1 key_c_r_reg_9_42 (.CK( clk ) , .D( key_c_r_8_42 ) , .Q( key_c_r_9_42 ) );
  DFF_X1 key_c_r_reg_9_43 (.CK( clk ) , .D( key_c_r_8_43 ) , .Q( key_c_r_9_43 ) );
  DFF_X1 key_c_r_reg_9_44 (.CK( clk ) , .D( key_c_r_8_44 ) , .Q( key_c_r_9_44 ) );
  DFF_X1 key_c_r_reg_9_45 (.CK( clk ) , .D( key_c_r_8_45 ) , .Q( key_c_r_9_45 ) );
  DFF_X1 key_c_r_reg_9_46 (.CK( clk ) , .D( key_c_r_8_46 ) , .Q( key_c_r_9_46 ) );
  DFF_X1 key_c_r_reg_9_47 (.CK( clk ) , .D( key_c_r_8_47 ) , .Q( key_c_r_9_47 ) );
  DFF_X1 key_c_r_reg_9_48 (.CK( clk ) , .D( key_c_r_8_48 ) , .Q( key_c_r_9_48 ) );
  DFF_X1 key_c_r_reg_9_49 (.CK( clk ) , .D( key_c_r_8_49 ) , .Q( key_c_r_9_49 ) );
  DFF_X1 key_c_r_reg_9_5 (.CK( clk ) , .D( key_c_r_8_5 ) , .Q( key_c_r_9_5 ) );
  DFF_X1 key_c_r_reg_9_50 (.CK( clk ) , .D( key_c_r_8_50 ) , .Q( key_c_r_9_50 ) );
  DFF_X1 key_c_r_reg_9_51 (.CK( clk ) , .D( key_c_r_8_51 ) , .Q( key_c_r_9_51 ) );
  DFF_X1 key_c_r_reg_9_52 (.CK( clk ) , .D( key_c_r_8_52 ) , .Q( key_c_r_9_52 ) );
  DFF_X1 key_c_r_reg_9_53 (.CK( clk ) , .D( key_c_r_8_53 ) , .Q( key_c_r_9_53 ) );
  DFF_X1 key_c_r_reg_9_54 (.CK( clk ) , .D( key_c_r_8_54 ) , .Q( key_c_r_9_54 ) );
  DFF_X1 key_c_r_reg_9_55 (.CK( clk ) , .D( key_c_r_8_55 ) , .Q( key_c_r_9_55 ) );
  DFF_X1 key_c_r_reg_9_6 (.CK( clk ) , .D( key_c_r_8_6 ) , .Q( key_c_r_9_6 ) );
  DFF_X1 key_c_r_reg_9_7 (.CK( clk ) , .D( key_c_r_8_7 ) , .Q( key_c_r_9_7 ) );
  DFF_X1 key_c_r_reg_9_8 (.CK( clk ) , .D( key_c_r_8_8 ) , .Q( key_c_r_9_8 ) );
  DFF_X1 key_c_r_reg_9_9 (.CK( clk ) , .D( key_c_r_8_9 ) , .Q( key_c_r_9_9 ) );
  DFF_X1 u0_L0_reg_1 (.CK( clk ) , .Q( u0_L0_1 ) , .D( u0_desIn_r_7 ) );
  DFF_X1 u0_L0_reg_10 (.CK( clk ) , .Q( u0_L0_10 ) , .D( u0_desIn_r_13 ) );
  DFF_X1 u0_L0_reg_11 (.CK( clk ) , .Q( u0_L0_11 ) , .D( u0_desIn_r_21 ) );
  DFF_X1 u0_L0_reg_12 (.CK( clk ) , .Q( u0_L0_12 ) , .D( u0_desIn_r_29 ) );
  DFF_X1 u0_L0_reg_13 (.CK( clk ) , .Q( u0_L0_13 ) , .D( u0_desIn_r_37 ) );
  DFF_X1 u0_L0_reg_14 (.CK( clk ) , .Q( u0_L0_14 ) , .D( u0_desIn_r_45 ) );
  DFF_X1 u0_L0_reg_15 (.CK( clk ) , .Q( u0_L0_15 ) , .D( u0_desIn_r_53 ) );
  DFF_X1 u0_L0_reg_16 (.CK( clk ) , .Q( u0_L0_16 ) , .D( u0_desIn_r_61 ) );
  DFF_X1 u0_L0_reg_17 (.CK( clk ) , .Q( u0_L0_17 ) , .D( u0_desIn_r_3 ) );
  DFF_X1 u0_L0_reg_18 (.CK( clk ) , .Q( u0_L0_18 ) , .D( u0_desIn_r_11 ) );
  DFF_X1 u0_L0_reg_19 (.CK( clk ) , .Q( u0_L0_19 ) , .D( u0_desIn_r_19 ) );
  DFF_X1 u0_L0_reg_2 (.CK( clk ) , .Q( u0_L0_2 ) , .D( u0_desIn_r_15 ) );
  DFF_X1 u0_L0_reg_20 (.CK( clk ) , .Q( u0_L0_20 ) , .D( u0_desIn_r_27 ) );
  DFF_X1 u0_L0_reg_21 (.CK( clk ) , .Q( u0_L0_21 ) , .D( u0_desIn_r_35 ) );
  DFF_X1 u0_L0_reg_22 (.CK( clk ) , .Q( u0_L0_22 ) , .D( u0_desIn_r_43 ) );
  DFF_X1 u0_L0_reg_23 (.CK( clk ) , .Q( u0_L0_23 ) , .D( u0_desIn_r_51 ) );
  DFF_X1 u0_L0_reg_24 (.CK( clk ) , .Q( u0_L0_24 ) , .D( u0_desIn_r_59 ) );
  DFF_X1 u0_L0_reg_25 (.CK( clk ) , .Q( u0_L0_25 ) , .D( u0_desIn_r_1 ) );
  DFF_X1 u0_L0_reg_26 (.CK( clk ) , .Q( u0_L0_26 ) , .D( u0_desIn_r_9 ) );
  DFF_X1 u0_L0_reg_27 (.CK( clk ) , .Q( u0_L0_27 ) , .D( u0_desIn_r_17 ) );
  DFF_X1 u0_L0_reg_28 (.CK( clk ) , .Q( u0_L0_28 ) , .D( u0_desIn_r_25 ) );
  DFF_X1 u0_L0_reg_29 (.CK( clk ) , .Q( u0_L0_29 ) , .D( u0_desIn_r_33 ) );
  DFF_X1 u0_L0_reg_3 (.CK( clk ) , .Q( u0_L0_3 ) , .D( u0_desIn_r_23 ) );
  DFF_X1 u0_L0_reg_30 (.CK( clk ) , .Q( u0_L0_30 ) , .D( u0_desIn_r_41 ) );
  DFF_X1 u0_L0_reg_31 (.CK( clk ) , .Q( u0_L0_31 ) , .D( u0_desIn_r_49 ) );
  DFF_X1 u0_L0_reg_32 (.CK( clk ) , .Q( u0_L0_32 ) , .D( u0_desIn_r_57 ) );
  DFF_X1 u0_L0_reg_4 (.CK( clk ) , .Q( u0_L0_4 ) , .D( u0_desIn_r_31 ) );
  DFF_X1 u0_L0_reg_5 (.CK( clk ) , .Q( u0_L0_5 ) , .D( u0_desIn_r_39 ) );
  DFF_X1 u0_L0_reg_6 (.CK( clk ) , .Q( u0_L0_6 ) , .D( u0_desIn_r_47 ) );
  DFF_X1 u0_L0_reg_7 (.CK( clk ) , .Q( u0_L0_7 ) , .D( u0_desIn_r_55 ) );
  DFF_X1 u0_L0_reg_8 (.CK( clk ) , .Q( u0_L0_8 ) , .D( u0_desIn_r_63 ) );
  DFF_X1 u0_L0_reg_9 (.CK( clk ) , .Q( u0_L0_9 ) , .D( u0_desIn_r_5 ) );
  DFF_X1 u0_L10_reg_1 (.CK( clk ) , .Q( u0_L10_1 ) , .D( u0_R9_1 ) );
  DFF_X1 u0_L10_reg_10 (.CK( clk ) , .Q( u0_L10_10 ) , .D( u0_R9_10 ) );
  DFF_X1 u0_L10_reg_11 (.CK( clk ) , .Q( u0_L10_11 ) , .D( u0_R9_11 ) );
  DFF_X1 u0_L10_reg_12 (.CK( clk ) , .Q( u0_L10_12 ) , .D( u0_R9_12 ) );
  DFF_X1 u0_L10_reg_13 (.CK( clk ) , .Q( u0_L10_13 ) , .D( u0_R9_13 ) );
  DFF_X1 u0_L10_reg_14 (.CK( clk ) , .Q( u0_L10_14 ) , .D( u0_R9_14 ) );
  DFF_X1 u0_L10_reg_15 (.CK( clk ) , .Q( u0_L10_15 ) , .D( u0_R9_15 ) );
  DFF_X1 u0_L10_reg_16 (.CK( clk ) , .Q( u0_L10_16 ) , .D( u0_R9_16 ) );
  DFF_X1 u0_L10_reg_17 (.CK( clk ) , .Q( u0_L10_17 ) , .D( u0_R9_17 ) );
  DFF_X1 u0_L10_reg_18 (.CK( clk ) , .Q( u0_L10_18 ) , .D( u0_R9_18 ) );
  DFF_X1 u0_L10_reg_19 (.CK( clk ) , .Q( u0_L10_19 ) , .D( u0_R9_19 ) );
  DFF_X1 u0_L10_reg_2 (.CK( clk ) , .Q( u0_L10_2 ) , .D( u0_R9_2 ) );
  DFF_X1 u0_L10_reg_20 (.CK( clk ) , .Q( u0_L10_20 ) , .D( u0_R9_20 ) );
  DFF_X1 u0_L10_reg_21 (.CK( clk ) , .Q( u0_L10_21 ) , .D( u0_R9_21 ) );
  DFF_X1 u0_L10_reg_22 (.CK( clk ) , .Q( u0_L10_22 ) , .D( u0_R9_22 ) );
  DFF_X1 u0_L10_reg_23 (.CK( clk ) , .Q( u0_L10_23 ) , .D( u0_R9_23 ) );
  DFF_X1 u0_L10_reg_24 (.CK( clk ) , .Q( u0_L10_24 ) , .D( u0_R9_24 ) );
  DFF_X1 u0_L10_reg_25 (.CK( clk ) , .Q( u0_L10_25 ) , .D( u0_R9_25 ) );
  DFF_X1 u0_L10_reg_26 (.CK( clk ) , .Q( u0_L10_26 ) , .D( u0_R9_26 ) );
  DFF_X1 u0_L10_reg_27 (.CK( clk ) , .Q( u0_L10_27 ) , .D( u0_R9_27 ) );
  DFF_X1 u0_L10_reg_28 (.CK( clk ) , .Q( u0_L10_28 ) , .D( u0_R9_28 ) );
  DFF_X1 u0_L10_reg_29 (.CK( clk ) , .Q( u0_L10_29 ) , .D( u0_R9_29 ) );
  DFF_X1 u0_L10_reg_3 (.CK( clk ) , .Q( u0_L10_3 ) , .D( u0_R9_3 ) );
  DFF_X1 u0_L10_reg_30 (.CK( clk ) , .Q( u0_L10_30 ) , .D( u0_R9_30 ) );
  DFF_X1 u0_L10_reg_31 (.CK( clk ) , .Q( u0_L10_31 ) , .D( u0_R9_31 ) );
  DFF_X1 u0_L10_reg_32 (.CK( clk ) , .Q( u0_L10_32 ) , .D( u0_R9_32 ) );
  DFF_X1 u0_L10_reg_4 (.CK( clk ) , .Q( u0_L10_4 ) , .D( u0_R9_4 ) );
  DFF_X1 u0_L10_reg_5 (.CK( clk ) , .Q( u0_L10_5 ) , .D( u0_R9_5 ) );
  DFF_X1 u0_L10_reg_6 (.CK( clk ) , .Q( u0_L10_6 ) , .D( u0_R9_6 ) );
  DFF_X1 u0_L10_reg_7 (.CK( clk ) , .Q( u0_L10_7 ) , .D( u0_R9_7 ) );
  DFF_X1 u0_L10_reg_8 (.CK( clk ) , .Q( u0_L10_8 ) , .D( u0_R9_8 ) );
  DFF_X1 u0_L10_reg_9 (.CK( clk ) , .Q( u0_L10_9 ) , .D( u0_R9_9 ) );
  DFF_X1 u0_L11_reg_1 (.CK( clk ) , .Q( u0_L11_1 ) , .D( u0_R10_1 ) );
  DFF_X1 u0_L11_reg_10 (.CK( clk ) , .Q( u0_L11_10 ) , .D( u0_R10_10 ) );
  DFF_X1 u0_L11_reg_11 (.CK( clk ) , .Q( u0_L11_11 ) , .D( u0_R10_11 ) );
  DFF_X1 u0_L11_reg_12 (.CK( clk ) , .Q( u0_L11_12 ) , .D( u0_R10_12 ) );
  DFF_X1 u0_L11_reg_13 (.CK( clk ) , .Q( u0_L11_13 ) , .D( u0_R10_13 ) );
  DFF_X1 u0_L11_reg_14 (.CK( clk ) , .Q( u0_L11_14 ) , .D( u0_R10_14 ) );
  DFF_X1 u0_L11_reg_15 (.CK( clk ) , .Q( u0_L11_15 ) , .D( u0_R10_15 ) );
  DFF_X1 u0_L11_reg_16 (.CK( clk ) , .Q( u0_L11_16 ) , .D( u0_R10_16 ) );
  DFF_X1 u0_L11_reg_17 (.CK( clk ) , .Q( u0_L11_17 ) , .D( u0_R10_17 ) );
  DFF_X1 u0_L11_reg_18 (.CK( clk ) , .Q( u0_L11_18 ) , .D( u0_R10_18 ) );
  DFF_X1 u0_L11_reg_19 (.CK( clk ) , .Q( u0_L11_19 ) , .D( u0_R10_19 ) );
  DFF_X1 u0_L11_reg_2 (.CK( clk ) , .Q( u0_L11_2 ) , .D( u0_R10_2 ) );
  DFF_X1 u0_L11_reg_20 (.CK( clk ) , .Q( u0_L11_20 ) , .D( u0_R10_20 ) );
  DFF_X1 u0_L11_reg_21 (.CK( clk ) , .Q( u0_L11_21 ) , .D( u0_R10_21 ) );
  DFF_X1 u0_L11_reg_22 (.CK( clk ) , .Q( u0_L11_22 ) , .D( u0_R10_22 ) );
  DFF_X1 u0_L11_reg_23 (.CK( clk ) , .Q( u0_L11_23 ) , .D( u0_R10_23 ) );
  DFF_X1 u0_L11_reg_24 (.CK( clk ) , .Q( u0_L11_24 ) , .D( u0_R10_24 ) );
  DFF_X1 u0_L11_reg_25 (.CK( clk ) , .Q( u0_L11_25 ) , .D( u0_R10_25 ) );
  DFF_X1 u0_L11_reg_26 (.CK( clk ) , .Q( u0_L11_26 ) , .D( u0_R10_26 ) );
  DFF_X1 u0_L11_reg_27 (.CK( clk ) , .Q( u0_L11_27 ) , .D( u0_R10_27 ) );
  DFF_X1 u0_L11_reg_28 (.CK( clk ) , .Q( u0_L11_28 ) , .D( u0_R10_28 ) );
  DFF_X1 u0_L11_reg_29 (.CK( clk ) , .Q( u0_L11_29 ) , .D( u0_R10_29 ) );
  DFF_X1 u0_L11_reg_3 (.CK( clk ) , .Q( u0_L11_3 ) , .D( u0_R10_3 ) );
  DFF_X1 u0_L11_reg_30 (.CK( clk ) , .Q( u0_L11_30 ) , .D( u0_R10_30 ) );
  DFF_X1 u0_L11_reg_31 (.CK( clk ) , .Q( u0_L11_31 ) , .D( u0_R10_31 ) );
  DFF_X1 u0_L11_reg_32 (.CK( clk ) , .Q( u0_L11_32 ) , .D( u0_R10_32 ) );
  DFF_X1 u0_L11_reg_4 (.CK( clk ) , .Q( u0_L11_4 ) , .D( u0_R10_4 ) );
  DFF_X1 u0_L11_reg_5 (.CK( clk ) , .Q( u0_L11_5 ) , .D( u0_R10_5 ) );
  DFF_X1 u0_L11_reg_6 (.CK( clk ) , .Q( u0_L11_6 ) , .D( u0_R10_6 ) );
  DFF_X1 u0_L11_reg_7 (.CK( clk ) , .Q( u0_L11_7 ) , .D( u0_R10_7 ) );
  DFF_X1 u0_L11_reg_8 (.CK( clk ) , .Q( u0_L11_8 ) , .D( u0_R10_8 ) );
  DFF_X1 u0_L11_reg_9 (.CK( clk ) , .Q( u0_L11_9 ) , .D( u0_R10_9 ) );
  DFF_X1 u0_L12_reg_1 (.CK( clk ) , .Q( u0_L12_1 ) , .D( u0_R11_1 ) );
  DFF_X1 u0_L12_reg_10 (.CK( clk ) , .Q( u0_L12_10 ) , .D( u0_R11_10 ) );
  DFF_X1 u0_L12_reg_11 (.CK( clk ) , .Q( u0_L12_11 ) , .D( u0_R11_11 ) );
  DFF_X1 u0_L12_reg_12 (.CK( clk ) , .Q( u0_L12_12 ) , .D( u0_R11_12 ) );
  DFF_X1 u0_L12_reg_13 (.CK( clk ) , .Q( u0_L12_13 ) , .D( u0_R11_13 ) );
  DFF_X1 u0_L12_reg_14 (.CK( clk ) , .Q( u0_L12_14 ) , .D( u0_R11_14 ) );
  DFF_X1 u0_L12_reg_15 (.CK( clk ) , .Q( u0_L12_15 ) , .D( u0_R11_15 ) );
  DFF_X1 u0_L12_reg_16 (.CK( clk ) , .Q( u0_L12_16 ) , .D( u0_R11_16 ) );
  DFF_X1 u0_L12_reg_17 (.CK( clk ) , .Q( u0_L12_17 ) , .D( u0_R11_17 ) );
  DFF_X1 u0_L12_reg_18 (.CK( clk ) , .Q( u0_L12_18 ) , .D( u0_R11_18 ) );
  DFF_X1 u0_L12_reg_19 (.CK( clk ) , .Q( u0_L12_19 ) , .D( u0_R11_19 ) );
  DFF_X1 u0_L12_reg_2 (.CK( clk ) , .Q( u0_L12_2 ) , .D( u0_R11_2 ) );
  DFF_X1 u0_L12_reg_20 (.CK( clk ) , .Q( u0_L12_20 ) , .D( u0_R11_20 ) );
  DFF_X1 u0_L12_reg_21 (.CK( clk ) , .Q( u0_L12_21 ) , .D( u0_R11_21 ) );
  DFF_X1 u0_L12_reg_22 (.CK( clk ) , .Q( u0_L12_22 ) , .D( u0_R11_22 ) );
  DFF_X1 u0_L12_reg_23 (.CK( clk ) , .Q( u0_L12_23 ) , .D( u0_R11_23 ) );
  DFF_X1 u0_L12_reg_24 (.CK( clk ) , .Q( u0_L12_24 ) , .D( u0_R11_24 ) );
  DFF_X1 u0_L12_reg_25 (.CK( clk ) , .Q( u0_L12_25 ) , .D( u0_R11_25 ) );
  DFF_X1 u0_L12_reg_26 (.CK( clk ) , .Q( u0_L12_26 ) , .D( u0_R11_26 ) );
  DFF_X1 u0_L12_reg_27 (.CK( clk ) , .Q( u0_L12_27 ) , .D( u0_R11_27 ) );
  DFF_X1 u0_L12_reg_28 (.CK( clk ) , .Q( u0_L12_28 ) , .D( u0_R11_28 ) );
  DFF_X1 u0_L12_reg_29 (.CK( clk ) , .Q( u0_L12_29 ) , .D( u0_R11_29 ) );
  DFF_X1 u0_L12_reg_3 (.CK( clk ) , .Q( u0_L12_3 ) , .D( u0_R11_3 ) );
  DFF_X1 u0_L12_reg_30 (.CK( clk ) , .Q( u0_L12_30 ) , .D( u0_R11_30 ) );
  DFF_X1 u0_L12_reg_31 (.CK( clk ) , .Q( u0_L12_31 ) , .D( u0_R11_31 ) );
  DFF_X1 u0_L12_reg_32 (.CK( clk ) , .Q( u0_L12_32 ) , .D( u0_R11_32 ) );
  DFF_X1 u0_L12_reg_4 (.CK( clk ) , .Q( u0_L12_4 ) , .D( u0_R11_4 ) );
  DFF_X1 u0_L12_reg_5 (.CK( clk ) , .Q( u0_L12_5 ) , .D( u0_R11_5 ) );
  DFF_X1 u0_L12_reg_6 (.CK( clk ) , .Q( u0_L12_6 ) , .D( u0_R11_6 ) );
  DFF_X1 u0_L12_reg_7 (.CK( clk ) , .Q( u0_L12_7 ) , .D( u0_R11_7 ) );
  DFF_X1 u0_L12_reg_8 (.CK( clk ) , .Q( u0_L12_8 ) , .D( u0_R11_8 ) );
  DFF_X1 u0_L12_reg_9 (.CK( clk ) , .Q( u0_L12_9 ) , .D( u0_R11_9 ) );
  DFF_X1 u0_L13_reg_1 (.CK( clk ) , .Q( u0_L13_1 ) , .D( u0_R12_1 ) );
  DFF_X1 u0_L13_reg_10 (.CK( clk ) , .Q( u0_L13_10 ) , .D( u0_R12_10 ) );
  DFF_X1 u0_L13_reg_11 (.CK( clk ) , .Q( u0_L13_11 ) , .D( u0_R12_11 ) );
  DFF_X1 u0_L13_reg_12 (.CK( clk ) , .Q( u0_L13_12 ) , .D( u0_R12_12 ) );
  DFF_X1 u0_L13_reg_13 (.CK( clk ) , .Q( u0_L13_13 ) , .D( u0_R12_13 ) );
  DFF_X1 u0_L13_reg_14 (.CK( clk ) , .Q( u0_L13_14 ) , .D( u0_R12_14 ) );
  DFF_X1 u0_L13_reg_15 (.CK( clk ) , .Q( u0_L13_15 ) , .D( u0_R12_15 ) );
  DFF_X1 u0_L13_reg_16 (.CK( clk ) , .Q( u0_L13_16 ) , .D( u0_R12_16 ) );
  DFF_X1 u0_L13_reg_17 (.CK( clk ) , .Q( u0_L13_17 ) , .D( u0_R12_17 ) );
  DFF_X1 u0_L13_reg_18 (.CK( clk ) , .Q( u0_L13_18 ) , .D( u0_R12_18 ) );
  DFF_X1 u0_L13_reg_19 (.CK( clk ) , .Q( u0_L13_19 ) , .D( u0_R12_19 ) );
  DFF_X1 u0_L13_reg_2 (.CK( clk ) , .Q( u0_L13_2 ) , .D( u0_R12_2 ) );
  DFF_X1 u0_L13_reg_20 (.CK( clk ) , .Q( u0_L13_20 ) , .D( u0_R12_20 ) );
  DFF_X1 u0_L13_reg_21 (.CK( clk ) , .Q( u0_L13_21 ) , .D( u0_R12_21 ) );
  DFF_X1 u0_L13_reg_22 (.CK( clk ) , .Q( u0_L13_22 ) , .D( u0_R12_22 ) );
  DFF_X1 u0_L13_reg_23 (.CK( clk ) , .Q( u0_L13_23 ) , .D( u0_R12_23 ) );
  DFF_X1 u0_L13_reg_24 (.CK( clk ) , .Q( u0_L13_24 ) , .D( u0_R12_24 ) );
  DFF_X1 u0_L13_reg_25 (.CK( clk ) , .Q( u0_L13_25 ) , .D( u0_R12_25 ) );
  DFF_X1 u0_L13_reg_26 (.CK( clk ) , .Q( u0_L13_26 ) , .D( u0_R12_26 ) );
  DFF_X1 u0_L13_reg_27 (.CK( clk ) , .Q( u0_L13_27 ) , .D( u0_R12_27 ) );
  DFF_X1 u0_L13_reg_28 (.CK( clk ) , .Q( u0_L13_28 ) , .D( u0_R12_28 ) );
  DFF_X1 u0_L13_reg_29 (.CK( clk ) , .Q( u0_L13_29 ) , .D( u0_R12_29 ) );
  DFF_X1 u0_L13_reg_3 (.CK( clk ) , .Q( u0_L13_3 ) , .D( u0_R12_3 ) );
  DFF_X1 u0_L13_reg_30 (.CK( clk ) , .Q( u0_L13_30 ) , .D( u0_R12_30 ) );
  DFF_X1 u0_L13_reg_31 (.CK( clk ) , .Q( u0_L13_31 ) , .D( u0_R12_31 ) );
  DFF_X1 u0_L13_reg_32 (.CK( clk ) , .Q( u0_L13_32 ) , .D( u0_R12_32 ) );
  DFF_X1 u0_L13_reg_4 (.CK( clk ) , .Q( u0_L13_4 ) , .D( u0_R12_4 ) );
  DFF_X1 u0_L13_reg_5 (.CK( clk ) , .Q( u0_L13_5 ) , .D( u0_R12_5 ) );
  DFF_X1 u0_L13_reg_6 (.CK( clk ) , .Q( u0_L13_6 ) , .D( u0_R12_6 ) );
  DFF_X1 u0_L13_reg_7 (.CK( clk ) , .Q( u0_L13_7 ) , .D( u0_R12_7 ) );
  DFF_X1 u0_L13_reg_8 (.CK( clk ) , .Q( u0_L13_8 ) , .D( u0_R12_8 ) );
  DFF_X1 u0_L13_reg_9 (.CK( clk ) , .Q( u0_L13_9 ) , .D( u0_R12_9 ) );
  DFF_X1 u0_L14_reg_1 (.CK( clk ) , .Q( u0_L14_1 ) , .D( u0_R13_1 ) );
  DFF_X1 u0_L14_reg_10 (.CK( clk ) , .Q( u0_L14_10 ) , .D( u0_R13_10 ) );
  DFF_X1 u0_L14_reg_11 (.CK( clk ) , .Q( u0_L14_11 ) , .D( u0_R13_11 ) );
  DFF_X1 u0_L14_reg_12 (.CK( clk ) , .Q( u0_L14_12 ) , .D( u0_R13_12 ) );
  DFF_X1 u0_L14_reg_13 (.CK( clk ) , .Q( u0_L14_13 ) , .D( u0_R13_13 ) );
  DFF_X1 u0_L14_reg_14 (.CK( clk ) , .Q( u0_L14_14 ) , .D( u0_R13_14 ) );
  DFF_X1 u0_L14_reg_15 (.CK( clk ) , .Q( u0_L14_15 ) , .D( u0_R13_15 ) );
  DFF_X1 u0_L14_reg_16 (.CK( clk ) , .Q( u0_L14_16 ) , .D( u0_R13_16 ) );
  DFF_X1 u0_L14_reg_17 (.CK( clk ) , .Q( u0_L14_17 ) , .D( u0_R13_17 ) );
  DFF_X1 u0_L14_reg_18 (.CK( clk ) , .Q( u0_L14_18 ) , .D( u0_R13_18 ) );
  DFF_X1 u0_L14_reg_19 (.CK( clk ) , .Q( u0_L14_19 ) , .D( u0_R13_19 ) );
  DFF_X1 u0_L14_reg_2 (.CK( clk ) , .Q( u0_L14_2 ) , .D( u0_R13_2 ) );
  DFF_X1 u0_L14_reg_20 (.CK( clk ) , .Q( u0_L14_20 ) , .D( u0_R13_20 ) );
  DFF_X1 u0_L14_reg_21 (.CK( clk ) , .Q( u0_L14_21 ) , .D( u0_R13_21 ) );
  DFF_X1 u0_L14_reg_22 (.CK( clk ) , .Q( u0_L14_22 ) , .D( u0_R13_22 ) );
  DFF_X1 u0_L14_reg_23 (.CK( clk ) , .Q( u0_L14_23 ) , .D( u0_R13_23 ) );
  DFF_X1 u0_L14_reg_24 (.CK( clk ) , .Q( u0_L14_24 ) , .D( u0_R13_24 ) );
  DFF_X1 u0_L14_reg_25 (.CK( clk ) , .Q( u0_L14_25 ) , .D( u0_R13_25 ) );
  DFF_X1 u0_L14_reg_26 (.CK( clk ) , .Q( u0_L14_26 ) , .D( u0_R13_26 ) );
  DFF_X1 u0_L14_reg_27 (.CK( clk ) , .Q( u0_L14_27 ) , .D( u0_R13_27 ) );
  DFF_X1 u0_L14_reg_28 (.CK( clk ) , .Q( u0_L14_28 ) , .D( u0_R13_28 ) );
  DFF_X1 u0_L14_reg_29 (.CK( clk ) , .Q( u0_L14_29 ) , .D( u0_R13_29 ) );
  DFF_X1 u0_L14_reg_3 (.CK( clk ) , .Q( u0_L14_3 ) , .D( u0_R13_3 ) );
  DFF_X1 u0_L14_reg_30 (.CK( clk ) , .Q( u0_L14_30 ) , .D( u0_R13_30 ) );
  DFF_X1 u0_L14_reg_31 (.CK( clk ) , .Q( u0_L14_31 ) , .D( u0_R13_31 ) );
  DFF_X1 u0_L14_reg_32 (.CK( clk ) , .Q( u0_L14_32 ) , .D( u0_R13_32 ) );
  DFF_X1 u0_L14_reg_4 (.CK( clk ) , .Q( u0_L14_4 ) , .D( u0_R13_4 ) );
  DFF_X1 u0_L14_reg_5 (.CK( clk ) , .Q( u0_L14_5 ) , .D( u0_R13_5 ) );
  DFF_X1 u0_L14_reg_6 (.CK( clk ) , .Q( u0_L14_6 ) , .D( u0_R13_6 ) );
  DFF_X1 u0_L14_reg_7 (.CK( clk ) , .Q( u0_L14_7 ) , .D( u0_R13_7 ) );
  DFF_X1 u0_L14_reg_8 (.CK( clk ) , .Q( u0_L14_8 ) , .D( u0_R13_8 ) );
  DFF_X1 u0_L14_reg_9 (.CK( clk ) , .Q( u0_L14_9 ) , .D( u0_R13_9 ) );
  DFF_X1 u0_L1_reg_1 (.CK( clk ) , .Q( u0_L1_1 ) , .D( u0_R0_1 ) );
  DFF_X1 u0_L1_reg_10 (.CK( clk ) , .Q( u0_L1_10 ) , .D( u0_R0_10 ) );
  DFF_X1 u0_L1_reg_11 (.CK( clk ) , .Q( u0_L1_11 ) , .D( u0_R0_11 ) );
  DFF_X1 u0_L1_reg_12 (.CK( clk ) , .Q( u0_L1_12 ) , .D( u0_R0_12 ) );
  DFF_X1 u0_L1_reg_13 (.CK( clk ) , .Q( u0_L1_13 ) , .D( u0_R0_13 ) );
  DFF_X1 u0_L1_reg_14 (.CK( clk ) , .Q( u0_L1_14 ) , .D( u0_R0_14 ) );
  DFF_X1 u0_L1_reg_15 (.CK( clk ) , .Q( u0_L1_15 ) , .D( u0_R0_15 ) );
  DFF_X1 u0_L1_reg_16 (.CK( clk ) , .Q( u0_L1_16 ) , .D( u0_R0_16 ) );
  DFF_X1 u0_L1_reg_17 (.CK( clk ) , .Q( u0_L1_17 ) , .D( u0_R0_17 ) );
  DFF_X1 u0_L1_reg_18 (.CK( clk ) , .Q( u0_L1_18 ) , .D( u0_R0_18 ) );
  DFF_X1 u0_L1_reg_19 (.CK( clk ) , .Q( u0_L1_19 ) , .D( u0_R0_19 ) );
  DFF_X1 u0_L1_reg_2 (.CK( clk ) , .Q( u0_L1_2 ) , .D( u0_R0_2 ) );
  DFF_X1 u0_L1_reg_20 (.CK( clk ) , .Q( u0_L1_20 ) , .D( u0_R0_20 ) );
  DFF_X1 u0_L1_reg_21 (.CK( clk ) , .Q( u0_L1_21 ) , .D( u0_R0_21 ) );
  DFF_X1 u0_L1_reg_22 (.CK( clk ) , .Q( u0_L1_22 ) , .D( u0_R0_22 ) );
  DFF_X1 u0_L1_reg_23 (.CK( clk ) , .Q( u0_L1_23 ) , .D( u0_R0_23 ) );
  DFF_X1 u0_L1_reg_24 (.CK( clk ) , .Q( u0_L1_24 ) , .D( u0_R0_24 ) );
  DFF_X1 u0_L1_reg_25 (.CK( clk ) , .Q( u0_L1_25 ) , .D( u0_R0_25 ) );
  DFF_X1 u0_L1_reg_26 (.CK( clk ) , .Q( u0_L1_26 ) , .D( u0_R0_26 ) );
  DFF_X1 u0_L1_reg_27 (.CK( clk ) , .Q( u0_L1_27 ) , .D( u0_R0_27 ) );
  DFF_X1 u0_L1_reg_28 (.CK( clk ) , .Q( u0_L1_28 ) , .D( u0_R0_28 ) );
  DFF_X1 u0_L1_reg_29 (.CK( clk ) , .Q( u0_L1_29 ) , .D( u0_R0_29 ) );
  DFF_X1 u0_L1_reg_3 (.CK( clk ) , .Q( u0_L1_3 ) , .D( u0_R0_3 ) );
  DFF_X1 u0_L1_reg_30 (.CK( clk ) , .Q( u0_L1_30 ) , .D( u0_R0_30 ) );
  DFF_X1 u0_L1_reg_31 (.CK( clk ) , .Q( u0_L1_31 ) , .D( u0_R0_31 ) );
  DFF_X1 u0_L1_reg_32 (.CK( clk ) , .Q( u0_L1_32 ) , .D( u0_R0_32 ) );
  DFF_X1 u0_L1_reg_4 (.CK( clk ) , .Q( u0_L1_4 ) , .D( u0_R0_4 ) );
  DFF_X1 u0_L1_reg_5 (.CK( clk ) , .Q( u0_L1_5 ) , .D( u0_R0_5 ) );
  DFF_X1 u0_L1_reg_6 (.CK( clk ) , .Q( u0_L1_6 ) , .D( u0_R0_6 ) );
  DFF_X1 u0_L1_reg_7 (.CK( clk ) , .Q( u0_L1_7 ) , .D( u0_R0_7 ) );
  DFF_X1 u0_L1_reg_8 (.CK( clk ) , .Q( u0_L1_8 ) , .D( u0_R0_8 ) );
  DFF_X1 u0_L1_reg_9 (.CK( clk ) , .Q( u0_L1_9 ) , .D( u0_R0_9 ) );
  DFF_X1 u0_L2_reg_1 (.CK( clk ) , .Q( u0_L2_1 ) , .D( u0_R1_1 ) );
  DFF_X1 u0_L2_reg_10 (.CK( clk ) , .Q( u0_L2_10 ) , .D( u0_R1_10 ) );
  DFF_X1 u0_L2_reg_11 (.CK( clk ) , .Q( u0_L2_11 ) , .D( u0_R1_11 ) );
  DFF_X1 u0_L2_reg_12 (.CK( clk ) , .Q( u0_L2_12 ) , .D( u0_R1_12 ) );
  DFF_X1 u0_L2_reg_13 (.CK( clk ) , .Q( u0_L2_13 ) , .D( u0_R1_13 ) );
  DFF_X1 u0_L2_reg_14 (.CK( clk ) , .Q( u0_L2_14 ) , .D( u0_R1_14 ) );
  DFF_X1 u0_L2_reg_15 (.CK( clk ) , .Q( u0_L2_15 ) , .D( u0_R1_15 ) );
  DFF_X1 u0_L2_reg_16 (.CK( clk ) , .Q( u0_L2_16 ) , .D( u0_R1_16 ) );
  DFF_X1 u0_L2_reg_17 (.CK( clk ) , .Q( u0_L2_17 ) , .D( u0_R1_17 ) );
  DFF_X1 u0_L2_reg_18 (.CK( clk ) , .Q( u0_L2_18 ) , .D( u0_R1_18 ) );
  DFF_X1 u0_L2_reg_19 (.CK( clk ) , .Q( u0_L2_19 ) , .D( u0_R1_19 ) );
  DFF_X1 u0_L2_reg_2 (.CK( clk ) , .Q( u0_L2_2 ) , .D( u0_R1_2 ) );
  DFF_X1 u0_L2_reg_20 (.CK( clk ) , .Q( u0_L2_20 ) , .D( u0_R1_20 ) );
  DFF_X1 u0_L2_reg_21 (.CK( clk ) , .Q( u0_L2_21 ) , .D( u0_R1_21 ) );
  DFF_X1 u0_L2_reg_22 (.CK( clk ) , .Q( u0_L2_22 ) , .D( u0_R1_22 ) );
  DFF_X1 u0_L2_reg_23 (.CK( clk ) , .Q( u0_L2_23 ) , .D( u0_R1_23 ) );
  DFF_X1 u0_L2_reg_24 (.CK( clk ) , .Q( u0_L2_24 ) , .D( u0_R1_24 ) );
  DFF_X1 u0_L2_reg_25 (.CK( clk ) , .Q( u0_L2_25 ) , .D( u0_R1_25 ) );
  DFF_X1 u0_L2_reg_26 (.CK( clk ) , .Q( u0_L2_26 ) , .D( u0_R1_26 ) );
  DFF_X1 u0_L2_reg_27 (.CK( clk ) , .Q( u0_L2_27 ) , .D( u0_R1_27 ) );
  DFF_X1 u0_L2_reg_28 (.CK( clk ) , .Q( u0_L2_28 ) , .D( u0_R1_28 ) );
  DFF_X1 u0_L2_reg_29 (.CK( clk ) , .Q( u0_L2_29 ) , .D( u0_R1_29 ) );
  DFF_X1 u0_L2_reg_3 (.CK( clk ) , .Q( u0_L2_3 ) , .D( u0_R1_3 ) );
  DFF_X1 u0_L2_reg_30 (.CK( clk ) , .Q( u0_L2_30 ) , .D( u0_R1_30 ) );
  DFF_X1 u0_L2_reg_31 (.CK( clk ) , .Q( u0_L2_31 ) , .D( u0_R1_31 ) );
  DFF_X1 u0_L2_reg_32 (.CK( clk ) , .Q( u0_L2_32 ) , .D( u0_R1_32 ) );
  DFF_X1 u0_L2_reg_4 (.CK( clk ) , .Q( u0_L2_4 ) , .D( u0_R1_4 ) );
  DFF_X1 u0_L2_reg_5 (.CK( clk ) , .Q( u0_L2_5 ) , .D( u0_R1_5 ) );
  DFF_X1 u0_L2_reg_6 (.CK( clk ) , .Q( u0_L2_6 ) , .D( u0_R1_6 ) );
  DFF_X1 u0_L2_reg_7 (.CK( clk ) , .Q( u0_L2_7 ) , .D( u0_R1_7 ) );
  DFF_X1 u0_L2_reg_8 (.CK( clk ) , .Q( u0_L2_8 ) , .D( u0_R1_8 ) );
  DFF_X1 u0_L2_reg_9 (.CK( clk ) , .Q( u0_L2_9 ) , .D( u0_R1_9 ) );
  DFF_X1 u0_L3_reg_1 (.CK( clk ) , .Q( u0_L3_1 ) , .D( u0_R2_1 ) );
  DFF_X1 u0_L3_reg_10 (.CK( clk ) , .Q( u0_L3_10 ) , .D( u0_R2_10 ) );
  DFF_X1 u0_L3_reg_11 (.CK( clk ) , .Q( u0_L3_11 ) , .D( u0_R2_11 ) );
  DFF_X1 u0_L3_reg_12 (.CK( clk ) , .Q( u0_L3_12 ) , .D( u0_R2_12 ) );
  DFF_X1 u0_L3_reg_13 (.CK( clk ) , .Q( u0_L3_13 ) , .D( u0_R2_13 ) );
  DFF_X1 u0_L3_reg_14 (.CK( clk ) , .Q( u0_L3_14 ) , .D( u0_R2_14 ) );
  DFF_X1 u0_L3_reg_15 (.CK( clk ) , .Q( u0_L3_15 ) , .D( u0_R2_15 ) );
  DFF_X1 u0_L3_reg_16 (.CK( clk ) , .Q( u0_L3_16 ) , .D( u0_R2_16 ) );
  DFF_X1 u0_L3_reg_17 (.CK( clk ) , .Q( u0_L3_17 ) , .D( u0_R2_17 ) );
  DFF_X1 u0_L3_reg_18 (.CK( clk ) , .Q( u0_L3_18 ) , .D( u0_R2_18 ) );
  DFF_X1 u0_L3_reg_19 (.CK( clk ) , .Q( u0_L3_19 ) , .D( u0_R2_19 ) );
  DFF_X1 u0_L3_reg_2 (.CK( clk ) , .Q( u0_L3_2 ) , .D( u0_R2_2 ) );
  DFF_X1 u0_L3_reg_20 (.CK( clk ) , .Q( u0_L3_20 ) , .D( u0_R2_20 ) );
  DFF_X1 u0_L3_reg_21 (.CK( clk ) , .Q( u0_L3_21 ) , .D( u0_R2_21 ) );
  DFF_X1 u0_L3_reg_22 (.CK( clk ) , .Q( u0_L3_22 ) , .D( u0_R2_22 ) );
  DFF_X1 u0_L3_reg_23 (.CK( clk ) , .Q( u0_L3_23 ) , .D( u0_R2_23 ) );
  DFF_X1 u0_L3_reg_24 (.CK( clk ) , .Q( u0_L3_24 ) , .D( u0_R2_24 ) );
  DFF_X1 u0_L3_reg_25 (.CK( clk ) , .Q( u0_L3_25 ) , .D( u0_R2_25 ) );
  DFF_X1 u0_L3_reg_26 (.CK( clk ) , .Q( u0_L3_26 ) , .D( u0_R2_26 ) );
  DFF_X1 u0_L3_reg_27 (.CK( clk ) , .Q( u0_L3_27 ) , .D( u0_R2_27 ) );
  DFF_X1 u0_L3_reg_28 (.CK( clk ) , .Q( u0_L3_28 ) , .D( u0_R2_28 ) );
  DFF_X1 u0_L3_reg_29 (.CK( clk ) , .Q( u0_L3_29 ) , .D( u0_R2_29 ) );
  DFF_X1 u0_L3_reg_3 (.CK( clk ) , .Q( u0_L3_3 ) , .D( u0_R2_3 ) );
  DFF_X1 u0_L3_reg_30 (.CK( clk ) , .Q( u0_L3_30 ) , .D( u0_R2_30 ) );
  DFF_X1 u0_L3_reg_31 (.CK( clk ) , .Q( u0_L3_31 ) , .D( u0_R2_31 ) );
  DFF_X1 u0_L3_reg_32 (.CK( clk ) , .Q( u0_L3_32 ) , .D( u0_R2_32 ) );
  DFF_X1 u0_L3_reg_4 (.CK( clk ) , .Q( u0_L3_4 ) , .D( u0_R2_4 ) );
  DFF_X1 u0_L3_reg_5 (.CK( clk ) , .Q( u0_L3_5 ) , .D( u0_R2_5 ) );
  DFF_X1 u0_L3_reg_6 (.CK( clk ) , .Q( u0_L3_6 ) , .D( u0_R2_6 ) );
  DFF_X1 u0_L3_reg_7 (.CK( clk ) , .Q( u0_L3_7 ) , .D( u0_R2_7 ) );
  DFF_X1 u0_L3_reg_8 (.CK( clk ) , .Q( u0_L3_8 ) , .D( u0_R2_8 ) );
  DFF_X1 u0_L3_reg_9 (.CK( clk ) , .Q( u0_L3_9 ) , .D( u0_R2_9 ) );
  DFF_X1 u0_L4_reg_1 (.CK( clk ) , .Q( u0_L4_1 ) , .D( u0_R3_1 ) );
  DFF_X1 u0_L4_reg_10 (.CK( clk ) , .Q( u0_L4_10 ) , .D( u0_R3_10 ) );
  DFF_X1 u0_L4_reg_11 (.CK( clk ) , .Q( u0_L4_11 ) , .D( u0_R3_11 ) );
  DFF_X1 u0_L4_reg_12 (.CK( clk ) , .Q( u0_L4_12 ) , .D( u0_R3_12 ) );
  DFF_X1 u0_L4_reg_13 (.CK( clk ) , .Q( u0_L4_13 ) , .D( u0_R3_13 ) );
  DFF_X1 u0_L4_reg_14 (.CK( clk ) , .Q( u0_L4_14 ) , .D( u0_R3_14 ) );
  DFF_X1 u0_L4_reg_15 (.CK( clk ) , .Q( u0_L4_15 ) , .D( u0_R3_15 ) );
  DFF_X1 u0_L4_reg_16 (.CK( clk ) , .Q( u0_L4_16 ) , .D( u0_R3_16 ) );
  DFF_X1 u0_L4_reg_17 (.CK( clk ) , .Q( u0_L4_17 ) , .D( u0_R3_17 ) );
  DFF_X1 u0_L4_reg_18 (.CK( clk ) , .Q( u0_L4_18 ) , .D( u0_R3_18 ) );
  DFF_X1 u0_L4_reg_19 (.CK( clk ) , .Q( u0_L4_19 ) , .D( u0_R3_19 ) );
  DFF_X1 u0_L4_reg_2 (.CK( clk ) , .Q( u0_L4_2 ) , .D( u0_R3_2 ) );
  DFF_X1 u0_L4_reg_20 (.CK( clk ) , .Q( u0_L4_20 ) , .D( u0_R3_20 ) );
  DFF_X1 u0_L4_reg_21 (.CK( clk ) , .Q( u0_L4_21 ) , .D( u0_R3_21 ) );
  DFF_X1 u0_L4_reg_22 (.CK( clk ) , .Q( u0_L4_22 ) , .D( u0_R3_22 ) );
  DFF_X1 u0_L4_reg_23 (.CK( clk ) , .Q( u0_L4_23 ) , .D( u0_R3_23 ) );
  DFF_X1 u0_L4_reg_24 (.CK( clk ) , .Q( u0_L4_24 ) , .D( u0_R3_24 ) );
  DFF_X1 u0_L4_reg_25 (.CK( clk ) , .Q( u0_L4_25 ) , .D( u0_R3_25 ) );
  DFF_X1 u0_L4_reg_26 (.CK( clk ) , .Q( u0_L4_26 ) , .D( u0_R3_26 ) );
  DFF_X1 u0_L4_reg_27 (.CK( clk ) , .Q( u0_L4_27 ) , .D( u0_R3_27 ) );
  DFF_X1 u0_L4_reg_28 (.CK( clk ) , .Q( u0_L4_28 ) , .D( u0_R3_28 ) );
  DFF_X1 u0_L4_reg_29 (.CK( clk ) , .Q( u0_L4_29 ) , .D( u0_R3_29 ) );
  DFF_X1 u0_L4_reg_3 (.CK( clk ) , .Q( u0_L4_3 ) , .D( u0_R3_3 ) );
  DFF_X1 u0_L4_reg_30 (.CK( clk ) , .Q( u0_L4_30 ) , .D( u0_R3_30 ) );
  DFF_X1 u0_L4_reg_31 (.CK( clk ) , .Q( u0_L4_31 ) , .D( u0_R3_31 ) );
  DFF_X1 u0_L4_reg_32 (.CK( clk ) , .Q( u0_L4_32 ) , .D( u0_R3_32 ) );
  DFF_X1 u0_L4_reg_4 (.CK( clk ) , .Q( u0_L4_4 ) , .D( u0_R3_4 ) );
  DFF_X1 u0_L4_reg_5 (.CK( clk ) , .Q( u0_L4_5 ) , .D( u0_R3_5 ) );
  DFF_X1 u0_L4_reg_6 (.CK( clk ) , .Q( u0_L4_6 ) , .D( u0_R3_6 ) );
  DFF_X1 u0_L4_reg_7 (.CK( clk ) , .Q( u0_L4_7 ) , .D( u0_R3_7 ) );
  DFF_X1 u0_L4_reg_8 (.CK( clk ) , .Q( u0_L4_8 ) , .D( u0_R3_8 ) );
  DFF_X1 u0_L4_reg_9 (.CK( clk ) , .Q( u0_L4_9 ) , .D( u0_R3_9 ) );
  DFF_X1 u0_L5_reg_1 (.CK( clk ) , .Q( u0_L5_1 ) , .D( u0_R4_1 ) );
  DFF_X1 u0_L5_reg_10 (.CK( clk ) , .Q( u0_L5_10 ) , .D( u0_R4_10 ) );
  DFF_X1 u0_L5_reg_11 (.CK( clk ) , .Q( u0_L5_11 ) , .D( u0_R4_11 ) );
  DFF_X1 u0_L5_reg_12 (.CK( clk ) , .Q( u0_L5_12 ) , .D( u0_R4_12 ) );
  DFF_X1 u0_L5_reg_13 (.CK( clk ) , .Q( u0_L5_13 ) , .D( u0_R4_13 ) );
  DFF_X1 u0_L5_reg_14 (.CK( clk ) , .Q( u0_L5_14 ) , .D( u0_R4_14 ) );
  DFF_X1 u0_L5_reg_15 (.CK( clk ) , .Q( u0_L5_15 ) , .D( u0_R4_15 ) );
  DFF_X1 u0_L5_reg_16 (.CK( clk ) , .Q( u0_L5_16 ) , .D( u0_R4_16 ) );
  DFF_X1 u0_L5_reg_17 (.CK( clk ) , .Q( u0_L5_17 ) , .D( u0_R4_17 ) );
  DFF_X1 u0_L5_reg_18 (.CK( clk ) , .Q( u0_L5_18 ) , .D( u0_R4_18 ) );
  DFF_X1 u0_L5_reg_19 (.CK( clk ) , .Q( u0_L5_19 ) , .D( u0_R4_19 ) );
  DFF_X1 u0_L5_reg_2 (.CK( clk ) , .Q( u0_L5_2 ) , .D( u0_R4_2 ) );
  DFF_X1 u0_L5_reg_20 (.CK( clk ) , .Q( u0_L5_20 ) , .D( u0_R4_20 ) );
  DFF_X1 u0_L5_reg_21 (.CK( clk ) , .Q( u0_L5_21 ) , .D( u0_R4_21 ) );
  DFF_X1 u0_L5_reg_22 (.CK( clk ) , .Q( u0_L5_22 ) , .D( u0_R4_22 ) );
  DFF_X1 u0_L5_reg_23 (.CK( clk ) , .Q( u0_L5_23 ) , .D( u0_R4_23 ) );
  DFF_X1 u0_L5_reg_24 (.CK( clk ) , .Q( u0_L5_24 ) , .D( u0_R4_24 ) );
  DFF_X1 u0_L5_reg_25 (.CK( clk ) , .Q( u0_L5_25 ) , .D( u0_R4_25 ) );
  DFF_X1 u0_L5_reg_26 (.CK( clk ) , .Q( u0_L5_26 ) , .D( u0_R4_26 ) );
  DFF_X1 u0_L5_reg_27 (.CK( clk ) , .Q( u0_L5_27 ) , .D( u0_R4_27 ) );
  DFF_X1 u0_L5_reg_28 (.CK( clk ) , .Q( u0_L5_28 ) , .D( u0_R4_28 ) );
  DFF_X1 u0_L5_reg_29 (.CK( clk ) , .Q( u0_L5_29 ) , .D( u0_R4_29 ) );
  DFF_X1 u0_L5_reg_3 (.CK( clk ) , .Q( u0_L5_3 ) , .D( u0_R4_3 ) );
  DFF_X1 u0_L5_reg_30 (.CK( clk ) , .Q( u0_L5_30 ) , .D( u0_R4_30 ) );
  DFF_X1 u0_L5_reg_31 (.CK( clk ) , .Q( u0_L5_31 ) , .D( u0_R4_31 ) );
  DFF_X1 u0_L5_reg_32 (.CK( clk ) , .Q( u0_L5_32 ) , .D( u0_R4_32 ) );
  DFF_X1 u0_L5_reg_4 (.CK( clk ) , .Q( u0_L5_4 ) , .D( u0_R4_4 ) );
  DFF_X1 u0_L5_reg_5 (.CK( clk ) , .Q( u0_L5_5 ) , .D( u0_R4_5 ) );
  DFF_X1 u0_L5_reg_6 (.CK( clk ) , .Q( u0_L5_6 ) , .D( u0_R4_6 ) );
  DFF_X1 u0_L5_reg_7 (.CK( clk ) , .Q( u0_L5_7 ) , .D( u0_R4_7 ) );
  DFF_X1 u0_L5_reg_8 (.CK( clk ) , .Q( u0_L5_8 ) , .D( u0_R4_8 ) );
  DFF_X1 u0_L5_reg_9 (.CK( clk ) , .Q( u0_L5_9 ) , .D( u0_R4_9 ) );
  DFF_X1 u0_L6_reg_1 (.CK( clk ) , .Q( u0_L6_1 ) , .D( u0_R5_1 ) );
  DFF_X1 u0_L6_reg_10 (.CK( clk ) , .Q( u0_L6_10 ) , .D( u0_R5_10 ) );
  DFF_X1 u0_L6_reg_11 (.CK( clk ) , .Q( u0_L6_11 ) , .D( u0_R5_11 ) );
  DFF_X1 u0_L6_reg_12 (.CK( clk ) , .Q( u0_L6_12 ) , .D( u0_R5_12 ) );
  DFF_X1 u0_L6_reg_13 (.CK( clk ) , .Q( u0_L6_13 ) , .D( u0_R5_13 ) );
  DFF_X1 u0_L6_reg_14 (.CK( clk ) , .Q( u0_L6_14 ) , .D( u0_R5_14 ) );
  DFF_X1 u0_L6_reg_15 (.CK( clk ) , .Q( u0_L6_15 ) , .D( u0_R5_15 ) );
  DFF_X1 u0_L6_reg_16 (.CK( clk ) , .Q( u0_L6_16 ) , .D( u0_R5_16 ) );
  DFF_X1 u0_L6_reg_17 (.CK( clk ) , .Q( u0_L6_17 ) , .D( u0_R5_17 ) );
  DFF_X1 u0_L6_reg_18 (.CK( clk ) , .Q( u0_L6_18 ) , .D( u0_R5_18 ) );
  DFF_X1 u0_L6_reg_19 (.CK( clk ) , .Q( u0_L6_19 ) , .D( u0_R5_19 ) );
  DFF_X1 u0_L6_reg_2 (.CK( clk ) , .Q( u0_L6_2 ) , .D( u0_R5_2 ) );
  DFF_X1 u0_L6_reg_20 (.CK( clk ) , .Q( u0_L6_20 ) , .D( u0_R5_20 ) );
  DFF_X1 u0_L6_reg_21 (.CK( clk ) , .Q( u0_L6_21 ) , .D( u0_R5_21 ) );
  DFF_X1 u0_L6_reg_22 (.CK( clk ) , .Q( u0_L6_22 ) , .D( u0_R5_22 ) );
  DFF_X1 u0_L6_reg_23 (.CK( clk ) , .Q( u0_L6_23 ) , .D( u0_R5_23 ) );
  DFF_X1 u0_L6_reg_24 (.CK( clk ) , .Q( u0_L6_24 ) , .D( u0_R5_24 ) );
  DFF_X1 u0_L6_reg_25 (.CK( clk ) , .Q( u0_L6_25 ) , .D( u0_R5_25 ) );
  DFF_X1 u0_L6_reg_26 (.CK( clk ) , .Q( u0_L6_26 ) , .D( u0_R5_26 ) );
  DFF_X1 u0_L6_reg_27 (.CK( clk ) , .Q( u0_L6_27 ) , .D( u0_R5_27 ) );
  DFF_X1 u0_L6_reg_28 (.CK( clk ) , .Q( u0_L6_28 ) , .D( u0_R5_28 ) );
  DFF_X1 u0_L6_reg_29 (.CK( clk ) , .Q( u0_L6_29 ) , .D( u0_R5_29 ) );
  DFF_X1 u0_L6_reg_3 (.CK( clk ) , .Q( u0_L6_3 ) , .D( u0_R5_3 ) );
  DFF_X1 u0_L6_reg_30 (.CK( clk ) , .Q( u0_L6_30 ) , .D( u0_R5_30 ) );
  DFF_X1 u0_L6_reg_31 (.CK( clk ) , .Q( u0_L6_31 ) , .D( u0_R5_31 ) );
  DFF_X1 u0_L6_reg_32 (.CK( clk ) , .Q( u0_L6_32 ) , .D( u0_R5_32 ) );
  DFF_X1 u0_L6_reg_4 (.CK( clk ) , .Q( u0_L6_4 ) , .D( u0_R5_4 ) );
  DFF_X1 u0_L6_reg_5 (.CK( clk ) , .Q( u0_L6_5 ) , .D( u0_R5_5 ) );
  DFF_X1 u0_L6_reg_6 (.CK( clk ) , .Q( u0_L6_6 ) , .D( u0_R5_6 ) );
  DFF_X1 u0_L6_reg_7 (.CK( clk ) , .Q( u0_L6_7 ) , .D( u0_R5_7 ) );
  DFF_X1 u0_L6_reg_8 (.CK( clk ) , .Q( u0_L6_8 ) , .D( u0_R5_8 ) );
  DFF_X1 u0_L6_reg_9 (.CK( clk ) , .Q( u0_L6_9 ) , .D( u0_R5_9 ) );
  DFF_X1 u0_L7_reg_1 (.CK( clk ) , .Q( u0_L7_1 ) , .D( u0_R6_1 ) );
  DFF_X1 u0_L7_reg_10 (.CK( clk ) , .Q( u0_L7_10 ) , .D( u0_R6_10 ) );
  DFF_X1 u0_L7_reg_11 (.CK( clk ) , .Q( u0_L7_11 ) , .D( u0_R6_11 ) );
  DFF_X1 u0_L7_reg_12 (.CK( clk ) , .Q( u0_L7_12 ) , .D( u0_R6_12 ) );
  DFF_X1 u0_L7_reg_13 (.CK( clk ) , .Q( u0_L7_13 ) , .D( u0_R6_13 ) );
  DFF_X1 u0_L7_reg_14 (.CK( clk ) , .Q( u0_L7_14 ) , .D( u0_R6_14 ) );
  DFF_X1 u0_L7_reg_15 (.CK( clk ) , .Q( u0_L7_15 ) , .D( u0_R6_15 ) );
  DFF_X1 u0_L7_reg_16 (.CK( clk ) , .Q( u0_L7_16 ) , .D( u0_R6_16 ) );
  DFF_X1 u0_L7_reg_17 (.CK( clk ) , .Q( u0_L7_17 ) , .D( u0_R6_17 ) );
  DFF_X1 u0_L7_reg_18 (.CK( clk ) , .Q( u0_L7_18 ) , .D( u0_R6_18 ) );
  DFF_X1 u0_L7_reg_19 (.CK( clk ) , .Q( u0_L7_19 ) , .D( u0_R6_19 ) );
  DFF_X1 u0_L7_reg_2 (.CK( clk ) , .Q( u0_L7_2 ) , .D( u0_R6_2 ) );
  DFF_X1 u0_L7_reg_20 (.CK( clk ) , .Q( u0_L7_20 ) , .D( u0_R6_20 ) );
  DFF_X1 u0_L7_reg_21 (.CK( clk ) , .Q( u0_L7_21 ) , .D( u0_R6_21 ) );
  DFF_X1 u0_L7_reg_22 (.CK( clk ) , .Q( u0_L7_22 ) , .D( u0_R6_22 ) );
  DFF_X1 u0_L7_reg_23 (.CK( clk ) , .Q( u0_L7_23 ) , .D( u0_R6_23 ) );
  DFF_X1 u0_L7_reg_24 (.CK( clk ) , .Q( u0_L7_24 ) , .D( u0_R6_24 ) );
  DFF_X1 u0_L7_reg_25 (.CK( clk ) , .Q( u0_L7_25 ) , .D( u0_R6_25 ) );
  DFF_X1 u0_L7_reg_26 (.CK( clk ) , .Q( u0_L7_26 ) , .D( u0_R6_26 ) );
  DFF_X1 u0_L7_reg_27 (.CK( clk ) , .Q( u0_L7_27 ) , .D( u0_R6_27 ) );
  DFF_X1 u0_L7_reg_28 (.CK( clk ) , .Q( u0_L7_28 ) , .D( u0_R6_28 ) );
  DFF_X1 u0_L7_reg_29 (.CK( clk ) , .Q( u0_L7_29 ) , .D( u0_R6_29 ) );
  DFF_X1 u0_L7_reg_3 (.CK( clk ) , .Q( u0_L7_3 ) , .D( u0_R6_3 ) );
  DFF_X1 u0_L7_reg_30 (.CK( clk ) , .Q( u0_L7_30 ) , .D( u0_R6_30 ) );
  DFF_X1 u0_L7_reg_31 (.CK( clk ) , .Q( u0_L7_31 ) , .D( u0_R6_31 ) );
  DFF_X1 u0_L7_reg_32 (.CK( clk ) , .Q( u0_L7_32 ) , .D( u0_R6_32 ) );
  DFF_X1 u0_L7_reg_4 (.CK( clk ) , .Q( u0_L7_4 ) , .D( u0_R6_4 ) );
  DFF_X1 u0_L7_reg_5 (.CK( clk ) , .Q( u0_L7_5 ) , .D( u0_R6_5 ) );
  DFF_X1 u0_L7_reg_6 (.CK( clk ) , .Q( u0_L7_6 ) , .D( u0_R6_6 ) );
  DFF_X1 u0_L7_reg_7 (.CK( clk ) , .Q( u0_L7_7 ) , .D( u0_R6_7 ) );
  DFF_X1 u0_L7_reg_8 (.CK( clk ) , .Q( u0_L7_8 ) , .D( u0_R6_8 ) );
  DFF_X1 u0_L7_reg_9 (.CK( clk ) , .Q( u0_L7_9 ) , .D( u0_R6_9 ) );
  DFF_X1 u0_L8_reg_1 (.CK( clk ) , .Q( u0_L8_1 ) , .D( u0_R7_1 ) );
  DFF_X1 u0_L8_reg_10 (.CK( clk ) , .Q( u0_L8_10 ) , .D( u0_R7_10 ) );
  DFF_X1 u0_L8_reg_11 (.CK( clk ) , .Q( u0_L8_11 ) , .D( u0_R7_11 ) );
  DFF_X1 u0_L8_reg_12 (.CK( clk ) , .Q( u0_L8_12 ) , .D( u0_R7_12 ) );
  DFF_X1 u0_L8_reg_13 (.CK( clk ) , .Q( u0_L8_13 ) , .D( u0_R7_13 ) );
  DFF_X1 u0_L8_reg_14 (.CK( clk ) , .Q( u0_L8_14 ) , .D( u0_R7_14 ) );
  DFF_X1 u0_L8_reg_15 (.CK( clk ) , .Q( u0_L8_15 ) , .D( u0_R7_15 ) );
  DFF_X1 u0_L8_reg_16 (.CK( clk ) , .Q( u0_L8_16 ) , .D( u0_R7_16 ) );
  DFF_X1 u0_L8_reg_17 (.CK( clk ) , .Q( u0_L8_17 ) , .D( u0_R7_17 ) );
  DFF_X1 u0_L8_reg_18 (.CK( clk ) , .Q( u0_L8_18 ) , .D( u0_R7_18 ) );
  DFF_X1 u0_L8_reg_19 (.CK( clk ) , .Q( u0_L8_19 ) , .D( u0_R7_19 ) );
  DFF_X1 u0_L8_reg_2 (.CK( clk ) , .Q( u0_L8_2 ) , .D( u0_R7_2 ) );
  DFF_X1 u0_L8_reg_20 (.CK( clk ) , .Q( u0_L8_20 ) , .D( u0_R7_20 ) );
  DFF_X1 u0_L8_reg_21 (.CK( clk ) , .Q( u0_L8_21 ) , .D( u0_R7_21 ) );
  DFF_X1 u0_L8_reg_22 (.CK( clk ) , .Q( u0_L8_22 ) , .D( u0_R7_22 ) );
  DFF_X1 u0_L8_reg_23 (.CK( clk ) , .Q( u0_L8_23 ) , .D( u0_R7_23 ) );
  DFF_X1 u0_L8_reg_24 (.CK( clk ) , .Q( u0_L8_24 ) , .D( u0_R7_24 ) );
  DFF_X1 u0_L8_reg_25 (.CK( clk ) , .Q( u0_L8_25 ) , .D( u0_R7_25 ) );
  DFF_X1 u0_L8_reg_26 (.CK( clk ) , .Q( u0_L8_26 ) , .D( u0_R7_26 ) );
  DFF_X1 u0_L8_reg_27 (.CK( clk ) , .Q( u0_L8_27 ) , .D( u0_R7_27 ) );
  DFF_X1 u0_L8_reg_28 (.CK( clk ) , .Q( u0_L8_28 ) , .D( u0_R7_28 ) );
  DFF_X1 u0_L8_reg_29 (.CK( clk ) , .Q( u0_L8_29 ) , .D( u0_R7_29 ) );
  DFF_X1 u0_L8_reg_3 (.CK( clk ) , .Q( u0_L8_3 ) , .D( u0_R7_3 ) );
  DFF_X1 u0_L8_reg_30 (.CK( clk ) , .Q( u0_L8_30 ) , .D( u0_R7_30 ) );
  DFF_X1 u0_L8_reg_31 (.CK( clk ) , .Q( u0_L8_31 ) , .D( u0_R7_31 ) );
  DFF_X1 u0_L8_reg_32 (.CK( clk ) , .Q( u0_L8_32 ) , .D( u0_R7_32 ) );
  DFF_X1 u0_L8_reg_4 (.CK( clk ) , .Q( u0_L8_4 ) , .D( u0_R7_4 ) );
  DFF_X1 u0_L8_reg_5 (.CK( clk ) , .Q( u0_L8_5 ) , .D( u0_R7_5 ) );
  DFF_X1 u0_L8_reg_6 (.CK( clk ) , .Q( u0_L8_6 ) , .D( u0_R7_6 ) );
  DFF_X1 u0_L8_reg_7 (.CK( clk ) , .Q( u0_L8_7 ) , .D( u0_R7_7 ) );
  DFF_X1 u0_L8_reg_8 (.CK( clk ) , .Q( u0_L8_8 ) , .D( u0_R7_8 ) );
  DFF_X1 u0_L8_reg_9 (.CK( clk ) , .Q( u0_L8_9 ) , .D( u0_R7_9 ) );
  DFF_X1 u0_L9_reg_1 (.CK( clk ) , .Q( u0_L9_1 ) , .D( u0_R8_1 ) );
  DFF_X1 u0_L9_reg_10 (.CK( clk ) , .Q( u0_L9_10 ) , .D( u0_R8_10 ) );
  DFF_X1 u0_L9_reg_11 (.CK( clk ) , .Q( u0_L9_11 ) , .D( u0_R8_11 ) );
  DFF_X1 u0_L9_reg_12 (.CK( clk ) , .Q( u0_L9_12 ) , .D( u0_R8_12 ) );
  DFF_X1 u0_L9_reg_13 (.CK( clk ) , .Q( u0_L9_13 ) , .D( u0_R8_13 ) );
  DFF_X1 u0_L9_reg_14 (.CK( clk ) , .Q( u0_L9_14 ) , .D( u0_R8_14 ) );
  DFF_X1 u0_L9_reg_15 (.CK( clk ) , .Q( u0_L9_15 ) , .D( u0_R8_15 ) );
  DFF_X1 u0_L9_reg_16 (.CK( clk ) , .Q( u0_L9_16 ) , .D( u0_R8_16 ) );
  DFF_X1 u0_L9_reg_17 (.CK( clk ) , .Q( u0_L9_17 ) , .D( u0_R8_17 ) );
  DFF_X1 u0_L9_reg_18 (.CK( clk ) , .Q( u0_L9_18 ) , .D( u0_R8_18 ) );
  DFF_X1 u0_L9_reg_19 (.CK( clk ) , .Q( u0_L9_19 ) , .D( u0_R8_19 ) );
  DFF_X1 u0_L9_reg_2 (.CK( clk ) , .Q( u0_L9_2 ) , .D( u0_R8_2 ) );
  DFF_X1 u0_L9_reg_20 (.CK( clk ) , .Q( u0_L9_20 ) , .D( u0_R8_20 ) );
  DFF_X1 u0_L9_reg_21 (.CK( clk ) , .Q( u0_L9_21 ) , .D( u0_R8_21 ) );
  DFF_X1 u0_L9_reg_22 (.CK( clk ) , .Q( u0_L9_22 ) , .D( u0_R8_22 ) );
  DFF_X1 u0_L9_reg_23 (.CK( clk ) , .Q( u0_L9_23 ) , .D( u0_R8_23 ) );
  DFF_X1 u0_L9_reg_24 (.CK( clk ) , .Q( u0_L9_24 ) , .D( u0_R8_24 ) );
  DFF_X1 u0_L9_reg_25 (.CK( clk ) , .Q( u0_L9_25 ) , .D( u0_R8_25 ) );
  DFF_X1 u0_L9_reg_26 (.CK( clk ) , .Q( u0_L9_26 ) , .D( u0_R8_26 ) );
  DFF_X1 u0_L9_reg_27 (.CK( clk ) , .Q( u0_L9_27 ) , .D( u0_R8_27 ) );
  DFF_X1 u0_L9_reg_28 (.CK( clk ) , .Q( u0_L9_28 ) , .D( u0_R8_28 ) );
  DFF_X1 u0_L9_reg_29 (.CK( clk ) , .Q( u0_L9_29 ) , .D( u0_R8_29 ) );
  DFF_X1 u0_L9_reg_3 (.CK( clk ) , .Q( u0_L9_3 ) , .D( u0_R8_3 ) );
  DFF_X1 u0_L9_reg_30 (.CK( clk ) , .Q( u0_L9_30 ) , .D( u0_R8_30 ) );
  DFF_X1 u0_L9_reg_31 (.CK( clk ) , .Q( u0_L9_31 ) , .D( u0_R8_31 ) );
  DFF_X1 u0_L9_reg_32 (.CK( clk ) , .Q( u0_L9_32 ) , .D( u0_R8_32 ) );
  DFF_X1 u0_L9_reg_4 (.CK( clk ) , .Q( u0_L9_4 ) , .D( u0_R8_4 ) );
  DFF_X1 u0_L9_reg_5 (.CK( clk ) , .Q( u0_L9_5 ) , .D( u0_R8_5 ) );
  DFF_X1 u0_L9_reg_6 (.CK( clk ) , .Q( u0_L9_6 ) , .D( u0_R8_6 ) );
  DFF_X1 u0_L9_reg_7 (.CK( clk ) , .Q( u0_L9_7 ) , .D( u0_R8_7 ) );
  DFF_X1 u0_L9_reg_8 (.CK( clk ) , .Q( u0_L9_8 ) , .D( u0_R8_8 ) );
  DFF_X1 u0_L9_reg_9 (.CK( clk ) , .Q( u0_L9_9 ) , .D( u0_R8_9 ) );
  DFF_X1 u0_R0_reg_1 (.CK( clk ) , .D( u0_N0 ) , .Q( u0_R0_1 ) );
  DFF_X1 u0_R0_reg_10 (.CK( clk ) , .D( u0_N9 ) , .Q( u0_R0_10 ) );
  DFF_X1 u0_R0_reg_11 (.CK( clk ) , .D( u0_N10 ) , .Q( u0_R0_11 ) );
  DFF_X1 u0_R0_reg_12 (.CK( clk ) , .D( u0_N11 ) , .Q( u0_R0_12 ) );
  DFF_X1 u0_R0_reg_13 (.CK( clk ) , .D( u0_N12 ) , .Q( u0_R0_13 ) );
  DFF_X1 u0_R0_reg_14 (.CK( clk ) , .D( u0_N13 ) , .Q( u0_R0_14 ) );
  DFF_X1 u0_R0_reg_15 (.CK( clk ) , .D( u0_N14 ) , .Q( u0_R0_15 ) );
  DFF_X1 u0_R0_reg_16 (.CK( clk ) , .D( u0_N15 ) , .Q( u0_R0_16 ) );
  DFF_X1 u0_R0_reg_17 (.CK( clk ) , .D( u0_N16 ) , .Q( u0_R0_17 ) );
  DFF_X1 u0_R0_reg_18 (.CK( clk ) , .D( u0_N17 ) , .Q( u0_R0_18 ) );
  DFF_X1 u0_R0_reg_19 (.CK( clk ) , .D( u0_N18 ) , .Q( u0_R0_19 ) );
  DFF_X1 u0_R0_reg_2 (.CK( clk ) , .D( u0_N1 ) , .Q( u0_R0_2 ) );
  DFF_X1 u0_R0_reg_20 (.CK( clk ) , .D( u0_N19 ) , .Q( u0_R0_20 ) );
  DFF_X1 u0_R0_reg_21 (.CK( clk ) , .D( u0_N20 ) , .Q( u0_R0_21 ) );
  DFF_X1 u0_R0_reg_22 (.CK( clk ) , .D( u0_N21 ) , .Q( u0_R0_22 ) );
  DFF_X1 u0_R0_reg_23 (.CK( clk ) , .D( u0_N22 ) , .Q( u0_R0_23 ) );
  DFF_X1 u0_R0_reg_24 (.CK( clk ) , .D( u0_N23 ) , .Q( u0_R0_24 ) );
  DFF_X1 u0_R0_reg_25 (.CK( clk ) , .D( u0_N24 ) , .Q( u0_R0_25 ) );
  DFF_X1 u0_R0_reg_26 (.CK( clk ) , .D( u0_N25 ) , .Q( u0_R0_26 ) );
  DFF_X1 u0_R0_reg_27 (.CK( clk ) , .D( u0_N26 ) , .Q( u0_R0_27 ) );
  DFF_X1 u0_R0_reg_28 (.CK( clk ) , .D( u0_N27 ) , .Q( u0_R0_28 ) );
  DFF_X1 u0_R0_reg_29 (.CK( clk ) , .D( u0_N28 ) , .Q( u0_R0_29 ) );
  DFF_X1 u0_R0_reg_3 (.CK( clk ) , .D( u0_N2 ) , .Q( u0_R0_3 ) );
  DFF_X1 u0_R0_reg_30 (.CK( clk ) , .D( u0_N29 ) , .Q( u0_R0_30 ) );
  DFF_X1 u0_R0_reg_31 (.CK( clk ) , .D( u0_N30 ) , .Q( u0_R0_31 ) );
  DFF_X1 u0_R0_reg_32 (.CK( clk ) , .D( u0_N31 ) , .Q( u0_R0_32 ) );
  DFF_X1 u0_R0_reg_4 (.CK( clk ) , .D( u0_N3 ) , .Q( u0_R0_4 ) );
  DFF_X1 u0_R0_reg_5 (.CK( clk ) , .D( u0_N4 ) , .Q( u0_R0_5 ) );
  DFF_X1 u0_R0_reg_6 (.CK( clk ) , .D( u0_N5 ) , .Q( u0_R0_6 ) );
  DFF_X1 u0_R0_reg_7 (.CK( clk ) , .D( u0_N6 ) , .Q( u0_R0_7 ) );
  DFF_X1 u0_R0_reg_8 (.CK( clk ) , .D( u0_N7 ) , .Q( u0_R0_8 ) );
  DFF_X1 u0_R0_reg_9 (.CK( clk ) , .D( u0_N8 ) , .Q( u0_R0_9 ) );
  DFF_X1 u0_R10_reg_1 (.CK( clk ) , .D( u0_N320 ) , .Q( u0_R10_1 ) );
  DFF_X1 u0_R10_reg_10 (.CK( clk ) , .D( u0_N329 ) , .Q( u0_R10_10 ) );
  DFF_X1 u0_R10_reg_11 (.CK( clk ) , .D( u0_N330 ) , .Q( u0_R10_11 ) );
  DFF_X1 u0_R10_reg_12 (.CK( clk ) , .D( u0_N331 ) , .Q( u0_R10_12 ) );
  DFF_X1 u0_R10_reg_13 (.CK( clk ) , .D( u0_N332 ) , .Q( u0_R10_13 ) );
  DFF_X1 u0_R10_reg_14 (.CK( clk ) , .D( u0_N333 ) , .Q( u0_R10_14 ) );
  DFF_X1 u0_R10_reg_15 (.CK( clk ) , .D( u0_N334 ) , .Q( u0_R10_15 ) );
  DFF_X1 u0_R10_reg_16 (.CK( clk ) , .D( u0_N335 ) , .Q( u0_R10_16 ) );
  DFF_X1 u0_R10_reg_17 (.CK( clk ) , .D( u0_N336 ) , .Q( u0_R10_17 ) );
  DFF_X1 u0_R10_reg_18 (.CK( clk ) , .D( u0_N337 ) , .Q( u0_R10_18 ) );
  DFF_X1 u0_R10_reg_19 (.CK( clk ) , .D( u0_N338 ) , .Q( u0_R10_19 ) );
  DFF_X1 u0_R10_reg_2 (.CK( clk ) , .D( u0_N321 ) , .Q( u0_R10_2 ) );
  DFF_X1 u0_R10_reg_20 (.CK( clk ) , .D( u0_N339 ) , .Q( u0_R10_20 ) );
  DFF_X1 u0_R10_reg_21 (.CK( clk ) , .D( u0_N340 ) , .Q( u0_R10_21 ) );
  DFF_X1 u0_R10_reg_22 (.CK( clk ) , .D( u0_N341 ) , .Q( u0_R10_22 ) );
  DFF_X1 u0_R10_reg_23 (.CK( clk ) , .D( u0_N342 ) , .Q( u0_R10_23 ) );
  DFF_X1 u0_R10_reg_24 (.CK( clk ) , .D( u0_N343 ) , .Q( u0_R10_24 ) );
  DFF_X1 u0_R10_reg_25 (.CK( clk ) , .D( u0_N344 ) , .Q( u0_R10_25 ) );
  DFF_X1 u0_R10_reg_26 (.CK( clk ) , .D( u0_N345 ) , .Q( u0_R10_26 ) );
  DFF_X1 u0_R10_reg_27 (.CK( clk ) , .D( u0_N346 ) , .Q( u0_R10_27 ) );
  DFF_X1 u0_R10_reg_28 (.CK( clk ) , .D( u0_N347 ) , .Q( u0_R10_28 ) );
  DFF_X1 u0_R10_reg_29 (.CK( clk ) , .D( u0_N348 ) , .Q( u0_R10_29 ) );
  DFF_X1 u0_R10_reg_3 (.CK( clk ) , .D( u0_N322 ) , .Q( u0_R10_3 ) );
  DFF_X1 u0_R10_reg_30 (.CK( clk ) , .D( u0_N349 ) , .Q( u0_R10_30 ) );
  DFF_X1 u0_R10_reg_31 (.CK( clk ) , .D( u0_N350 ) , .Q( u0_R10_31 ) );
  DFF_X1 u0_R10_reg_32 (.CK( clk ) , .D( u0_N351 ) , .Q( u0_R10_32 ) );
  DFF_X1 u0_R10_reg_4 (.CK( clk ) , .D( u0_N323 ) , .Q( u0_R10_4 ) );
  DFF_X1 u0_R10_reg_5 (.CK( clk ) , .D( u0_N324 ) , .Q( u0_R10_5 ) );
  DFF_X1 u0_R10_reg_6 (.CK( clk ) , .D( u0_N325 ) , .Q( u0_R10_6 ) );
  DFF_X1 u0_R10_reg_7 (.CK( clk ) , .D( u0_N326 ) , .Q( u0_R10_7 ) );
  DFF_X1 u0_R10_reg_8 (.CK( clk ) , .D( u0_N327 ) , .Q( u0_R10_8 ) );
  DFF_X1 u0_R10_reg_9 (.CK( clk ) , .D( u0_N328 ) , .Q( u0_R10_9 ) );
  DFF_X1 u0_R11_reg_1 (.CK( clk ) , .D( u0_N352 ) , .Q( u0_R11_1 ) );
  DFF_X1 u0_R11_reg_10 (.CK( clk ) , .D( u0_N361 ) , .Q( u0_R11_10 ) );
  DFF_X1 u0_R11_reg_11 (.CK( clk ) , .D( u0_N362 ) , .Q( u0_R11_11 ) );
  DFF_X1 u0_R11_reg_12 (.CK( clk ) , .D( u0_N363 ) , .Q( u0_R11_12 ) );
  DFF_X1 u0_R11_reg_13 (.CK( clk ) , .D( u0_N364 ) , .Q( u0_R11_13 ) );
  DFF_X1 u0_R11_reg_14 (.CK( clk ) , .D( u0_N365 ) , .Q( u0_R11_14 ) );
  DFF_X1 u0_R11_reg_15 (.CK( clk ) , .D( u0_N366 ) , .Q( u0_R11_15 ) );
  DFF_X1 u0_R11_reg_16 (.CK( clk ) , .D( u0_N367 ) , .Q( u0_R11_16 ) );
  DFF_X1 u0_R11_reg_17 (.CK( clk ) , .D( u0_N368 ) , .Q( u0_R11_17 ) );
  DFF_X1 u0_R11_reg_18 (.CK( clk ) , .D( u0_N369 ) , .Q( u0_R11_18 ) );
  DFF_X1 u0_R11_reg_19 (.CK( clk ) , .D( u0_N370 ) , .Q( u0_R11_19 ) );
  DFF_X1 u0_R11_reg_2 (.CK( clk ) , .D( u0_N353 ) , .Q( u0_R11_2 ) );
  DFF_X1 u0_R11_reg_20 (.CK( clk ) , .D( u0_N371 ) , .Q( u0_R11_20 ) );
  DFF_X1 u0_R11_reg_21 (.CK( clk ) , .D( u0_N372 ) , .Q( u0_R11_21 ) );
  DFF_X1 u0_R11_reg_22 (.CK( clk ) , .D( u0_N373 ) , .Q( u0_R11_22 ) );
  DFF_X1 u0_R11_reg_23 (.CK( clk ) , .D( u0_N374 ) , .Q( u0_R11_23 ) );
  DFF_X1 u0_R11_reg_24 (.CK( clk ) , .D( u0_N375 ) , .Q( u0_R11_24 ) );
  DFF_X1 u0_R11_reg_25 (.CK( clk ) , .D( u0_N376 ) , .Q( u0_R11_25 ) );
  DFF_X1 u0_R11_reg_26 (.CK( clk ) , .D( u0_N377 ) , .Q( u0_R11_26 ) );
  DFF_X1 u0_R11_reg_27 (.CK( clk ) , .D( u0_N378 ) , .Q( u0_R11_27 ) );
  DFF_X1 u0_R11_reg_28 (.CK( clk ) , .D( u0_N379 ) , .Q( u0_R11_28 ) );
  DFF_X1 u0_R11_reg_29 (.CK( clk ) , .D( u0_N380 ) , .Q( u0_R11_29 ) );
  DFF_X1 u0_R11_reg_3 (.CK( clk ) , .D( u0_N354 ) , .Q( u0_R11_3 ) );
  DFF_X1 u0_R11_reg_30 (.CK( clk ) , .D( u0_N381 ) , .Q( u0_R11_30 ) );
  DFF_X1 u0_R11_reg_31 (.CK( clk ) , .D( u0_N382 ) , .Q( u0_R11_31 ) );
  DFF_X1 u0_R11_reg_32 (.CK( clk ) , .D( u0_N383 ) , .Q( u0_R11_32 ) );
  DFF_X1 u0_R11_reg_4 (.CK( clk ) , .D( u0_N355 ) , .Q( u0_R11_4 ) );
  DFF_X1 u0_R11_reg_5 (.CK( clk ) , .D( u0_N356 ) , .Q( u0_R11_5 ) );
  DFF_X1 u0_R11_reg_6 (.CK( clk ) , .D( u0_N357 ) , .Q( u0_R11_6 ) );
  DFF_X1 u0_R11_reg_7 (.CK( clk ) , .D( u0_N358 ) , .Q( u0_R11_7 ) );
  DFF_X1 u0_R11_reg_8 (.CK( clk ) , .D( u0_N359 ) , .Q( u0_R11_8 ) );
  DFF_X1 u0_R11_reg_9 (.CK( clk ) , .D( u0_N360 ) , .Q( u0_R11_9 ) );
  DFF_X1 u0_R12_reg_1 (.CK( clk ) , .D( u0_N384 ) , .Q( u0_R12_1 ) );
  DFF_X1 u0_R12_reg_10 (.CK( clk ) , .D( u0_N393 ) , .Q( u0_R12_10 ) );
  DFF_X1 u0_R12_reg_11 (.CK( clk ) , .D( u0_N394 ) , .Q( u0_R12_11 ) );
  DFF_X1 u0_R12_reg_12 (.CK( clk ) , .D( u0_N395 ) , .Q( u0_R12_12 ) );
  DFF_X1 u0_R12_reg_13 (.CK( clk ) , .D( u0_N396 ) , .Q( u0_R12_13 ) );
  DFF_X1 u0_R12_reg_14 (.CK( clk ) , .D( u0_N397 ) , .Q( u0_R12_14 ) );
  DFF_X1 u0_R12_reg_15 (.CK( clk ) , .D( u0_N398 ) , .Q( u0_R12_15 ) );
  DFF_X1 u0_R12_reg_16 (.CK( clk ) , .D( u0_N399 ) , .Q( u0_R12_16 ) );
  DFF_X1 u0_R12_reg_17 (.CK( clk ) , .D( u0_N400 ) , .Q( u0_R12_17 ) );
  DFF_X1 u0_R12_reg_18 (.CK( clk ) , .D( u0_N401 ) , .Q( u0_R12_18 ) );
  DFF_X1 u0_R12_reg_19 (.CK( clk ) , .D( u0_N402 ) , .Q( u0_R12_19 ) );
  DFF_X1 u0_R12_reg_2 (.CK( clk ) , .D( u0_N385 ) , .Q( u0_R12_2 ) );
  DFF_X1 u0_R12_reg_20 (.CK( clk ) , .D( u0_N403 ) , .Q( u0_R12_20 ) );
  DFF_X1 u0_R12_reg_21 (.CK( clk ) , .D( u0_N404 ) , .Q( u0_R12_21 ) );
  DFF_X1 u0_R12_reg_22 (.CK( clk ) , .D( u0_N405 ) , .Q( u0_R12_22 ) );
  DFF_X1 u0_R12_reg_23 (.CK( clk ) , .D( u0_N406 ) , .Q( u0_R12_23 ) );
  DFF_X1 u0_R12_reg_24 (.CK( clk ) , .D( u0_N407 ) , .Q( u0_R12_24 ) );
  DFF_X1 u0_R12_reg_25 (.CK( clk ) , .D( u0_N408 ) , .Q( u0_R12_25 ) );
  DFF_X1 u0_R12_reg_26 (.CK( clk ) , .D( u0_N409 ) , .Q( u0_R12_26 ) );
  DFF_X1 u0_R12_reg_27 (.CK( clk ) , .D( u0_N410 ) , .Q( u0_R12_27 ) );
  DFF_X1 u0_R12_reg_28 (.CK( clk ) , .D( u0_N411 ) , .Q( u0_R12_28 ) );
  DFF_X1 u0_R12_reg_29 (.CK( clk ) , .D( u0_N412 ) , .Q( u0_R12_29 ) );
  DFF_X1 u0_R12_reg_3 (.CK( clk ) , .D( u0_N386 ) , .Q( u0_R12_3 ) );
  DFF_X1 u0_R12_reg_30 (.CK( clk ) , .D( u0_N413 ) , .Q( u0_R12_30 ) );
  DFF_X1 u0_R12_reg_31 (.CK( clk ) , .D( u0_N414 ) , .Q( u0_R12_31 ) );
  DFF_X1 u0_R12_reg_32 (.CK( clk ) , .D( u0_N415 ) , .Q( u0_R12_32 ) );
  DFF_X1 u0_R12_reg_4 (.CK( clk ) , .D( u0_N387 ) , .Q( u0_R12_4 ) );
  DFF_X1 u0_R12_reg_5 (.CK( clk ) , .D( u0_N388 ) , .Q( u0_R12_5 ) );
  DFF_X1 u0_R12_reg_6 (.CK( clk ) , .D( u0_N389 ) , .Q( u0_R12_6 ) );
  DFF_X1 u0_R12_reg_7 (.CK( clk ) , .D( u0_N390 ) , .Q( u0_R12_7 ) );
  DFF_X1 u0_R12_reg_8 (.CK( clk ) , .D( u0_N391 ) , .Q( u0_R12_8 ) );
  DFF_X1 u0_R12_reg_9 (.CK( clk ) , .D( u0_N392 ) , .Q( u0_R12_9 ) );
  DFF_X1 u0_R13_reg_1 (.CK( clk ) , .D( u0_N416 ) , .Q( u0_R13_1 ) );
  DFF_X1 u0_R13_reg_10 (.CK( clk ) , .D( u0_N425 ) , .Q( u0_R13_10 ) );
  DFF_X1 u0_R13_reg_11 (.CK( clk ) , .D( u0_N426 ) , .Q( u0_R13_11 ) );
  DFF_X1 u0_R13_reg_12 (.CK( clk ) , .D( u0_N427 ) , .Q( u0_R13_12 ) );
  DFF_X1 u0_R13_reg_13 (.CK( clk ) , .D( u0_N428 ) , .Q( u0_R13_13 ) );
  DFF_X1 u0_R13_reg_14 (.CK( clk ) , .D( u0_N429 ) , .Q( u0_R13_14 ) );
  DFF_X1 u0_R13_reg_15 (.CK( clk ) , .D( u0_N430 ) , .Q( u0_R13_15 ) );
  DFF_X1 u0_R13_reg_16 (.CK( clk ) , .D( u0_N431 ) , .Q( u0_R13_16 ) );
  DFF_X1 u0_R13_reg_17 (.CK( clk ) , .D( u0_N432 ) , .Q( u0_R13_17 ) );
  DFF_X1 u0_R13_reg_18 (.CK( clk ) , .D( u0_N433 ) , .Q( u0_R13_18 ) );
  DFF_X1 u0_R13_reg_19 (.CK( clk ) , .D( u0_N434 ) , .Q( u0_R13_19 ) );
  DFF_X1 u0_R13_reg_2 (.CK( clk ) , .D( u0_N417 ) , .Q( u0_R13_2 ) );
  DFF_X1 u0_R13_reg_20 (.CK( clk ) , .D( u0_N435 ) , .Q( u0_R13_20 ) );
  DFF_X1 u0_R13_reg_21 (.CK( clk ) , .D( u0_N436 ) , .Q( u0_R13_21 ) );
  DFF_X1 u0_R13_reg_22 (.CK( clk ) , .D( u0_N437 ) , .Q( u0_R13_22 ) );
  DFF_X1 u0_R13_reg_23 (.CK( clk ) , .D( u0_N438 ) , .Q( u0_R13_23 ) );
  DFF_X1 u0_R13_reg_24 (.CK( clk ) , .D( u0_N439 ) , .Q( u0_R13_24 ) );
  DFF_X1 u0_R13_reg_25 (.CK( clk ) , .D( u0_N440 ) , .Q( u0_R13_25 ) );
  DFF_X1 u0_R13_reg_26 (.CK( clk ) , .D( u0_N441 ) , .Q( u0_R13_26 ) );
  DFF_X1 u0_R13_reg_27 (.CK( clk ) , .D( u0_N442 ) , .Q( u0_R13_27 ) );
  DFF_X1 u0_R13_reg_28 (.CK( clk ) , .D( u0_N443 ) , .Q( u0_R13_28 ) );
  DFF_X1 u0_R13_reg_29 (.CK( clk ) , .D( u0_N444 ) , .Q( u0_R13_29 ) );
  DFF_X1 u0_R13_reg_3 (.CK( clk ) , .D( u0_N418 ) , .Q( u0_R13_3 ) );
  DFF_X1 u0_R13_reg_30 (.CK( clk ) , .D( u0_N445 ) , .Q( u0_R13_30 ) );
  DFF_X1 u0_R13_reg_31 (.CK( clk ) , .D( u0_N446 ) , .Q( u0_R13_31 ) );
  DFF_X1 u0_R13_reg_32 (.CK( clk ) , .D( u0_N447 ) , .Q( u0_R13_32 ) );
  DFF_X1 u0_R13_reg_4 (.CK( clk ) , .D( u0_N419 ) , .Q( u0_R13_4 ) );
  DFF_X1 u0_R13_reg_5 (.CK( clk ) , .D( u0_N420 ) , .Q( u0_R13_5 ) );
  DFF_X1 u0_R13_reg_6 (.CK( clk ) , .D( u0_N421 ) , .Q( u0_R13_6 ) );
  DFF_X1 u0_R13_reg_7 (.CK( clk ) , .D( u0_N422 ) , .Q( u0_R13_7 ) );
  DFF_X1 u0_R13_reg_8 (.CK( clk ) , .D( u0_N423 ) , .Q( u0_R13_8 ) );
  DFF_X1 u0_R13_reg_9 (.CK( clk ) , .D( u0_N424 ) , .Q( u0_R13_9 ) );
  DFF_X1 u0_R14_reg_1 (.CK( clk ) , .Q( u0_FP_33 ) , .D( u0_N448 ) );
  DFF_X1 u0_R14_reg_10 (.CK( clk ) , .Q( u0_FP_42 ) , .D( u0_N457 ) );
  DFF_X1 u0_R14_reg_11 (.CK( clk ) , .Q( u0_FP_43 ) , .D( u0_N458 ) );
  DFF_X1 u0_R14_reg_12 (.CK( clk ) , .Q( u0_FP_44 ) , .D( u0_N459 ) );
  DFF_X1 u0_R14_reg_13 (.CK( clk ) , .Q( u0_FP_45 ) , .D( u0_N460 ) );
  DFF_X1 u0_R14_reg_14 (.CK( clk ) , .Q( u0_FP_46 ) , .D( u0_N461 ) );
  DFF_X1 u0_R14_reg_15 (.CK( clk ) , .Q( u0_FP_47 ) , .D( u0_N462 ) );
  DFF_X1 u0_R14_reg_16 (.CK( clk ) , .Q( u0_FP_48 ) , .D( u0_N463 ) );
  DFF_X1 u0_R14_reg_17 (.CK( clk ) , .Q( u0_FP_49 ) , .D( u0_N464 ) );
  DFF_X1 u0_R14_reg_18 (.CK( clk ) , .Q( u0_FP_50 ) , .D( u0_N465 ) );
  DFF_X1 u0_R14_reg_19 (.CK( clk ) , .Q( u0_FP_51 ) , .D( u0_N466 ) );
  DFF_X1 u0_R14_reg_2 (.CK( clk ) , .Q( u0_FP_34 ) , .D( u0_N449 ) );
  DFF_X1 u0_R14_reg_20 (.CK( clk ) , .Q( u0_FP_52 ) , .D( u0_N467 ) );
  DFF_X1 u0_R14_reg_21 (.CK( clk ) , .Q( u0_FP_53 ) , .D( u0_N468 ) );
  DFF_X1 u0_R14_reg_22 (.CK( clk ) , .Q( u0_FP_54 ) , .D( u0_N469 ) );
  DFF_X1 u0_R14_reg_23 (.CK( clk ) , .Q( u0_FP_55 ) , .D( u0_N470 ) );
  DFF_X1 u0_R14_reg_24 (.CK( clk ) , .Q( u0_FP_56 ) , .D( u0_N471 ) );
  DFF_X1 u0_R14_reg_25 (.CK( clk ) , .Q( u0_FP_57 ) , .D( u0_N472 ) );
  DFF_X1 u0_R14_reg_26 (.CK( clk ) , .Q( u0_FP_58 ) , .D( u0_N473 ) );
  DFF_X1 u0_R14_reg_27 (.CK( clk ) , .Q( u0_FP_59 ) , .D( u0_N474 ) );
  DFF_X1 u0_R14_reg_28 (.CK( clk ) , .Q( u0_FP_60 ) , .D( u0_N475 ) );
  DFF_X1 u0_R14_reg_29 (.CK( clk ) , .Q( u0_FP_61 ) , .D( u0_N476 ) );
  DFF_X1 u0_R14_reg_3 (.CK( clk ) , .Q( u0_FP_35 ) , .D( u0_N450 ) );
  DFF_X1 u0_R14_reg_30 (.CK( clk ) , .Q( u0_FP_62 ) , .D( u0_N477 ) );
  DFF_X1 u0_R14_reg_31 (.CK( clk ) , .Q( u0_FP_63 ) , .D( u0_N478 ) );
  DFF_X1 u0_R14_reg_32 (.CK( clk ) , .Q( u0_FP_64 ) , .D( u0_N479 ) );
  DFF_X1 u0_R14_reg_4 (.CK( clk ) , .Q( u0_FP_36 ) , .D( u0_N451 ) );
  DFF_X1 u0_R14_reg_5 (.CK( clk ) , .Q( u0_FP_37 ) , .D( u0_N452 ) );
  DFF_X1 u0_R14_reg_6 (.CK( clk ) , .Q( u0_FP_38 ) , .D( u0_N453 ) );
  DFF_X1 u0_R14_reg_7 (.CK( clk ) , .Q( u0_FP_39 ) , .D( u0_N454 ) );
  DFF_X1 u0_R14_reg_8 (.CK( clk ) , .Q( u0_FP_40 ) , .D( u0_N455 ) );
  DFF_X1 u0_R14_reg_9 (.CK( clk ) , .Q( u0_FP_41 ) , .D( u0_N456 ) );
  DFF_X1 u0_R1_reg_1 (.CK( clk ) , .D( u0_N32 ) , .Q( u0_R1_1 ) );
  DFF_X1 u0_R1_reg_10 (.CK( clk ) , .D( u0_N41 ) , .Q( u0_R1_10 ) );
  DFF_X1 u0_R1_reg_11 (.CK( clk ) , .D( u0_N42 ) , .Q( u0_R1_11 ) );
  DFF_X1 u0_R1_reg_12 (.CK( clk ) , .D( u0_N43 ) , .Q( u0_R1_12 ) );
  DFF_X1 u0_R1_reg_13 (.CK( clk ) , .D( u0_N44 ) , .Q( u0_R1_13 ) );
  DFF_X1 u0_R1_reg_14 (.CK( clk ) , .D( u0_N45 ) , .Q( u0_R1_14 ) );
  DFF_X1 u0_R1_reg_15 (.CK( clk ) , .D( u0_N46 ) , .Q( u0_R1_15 ) );
  DFF_X1 u0_R1_reg_16 (.CK( clk ) , .D( u0_N47 ) , .Q( u0_R1_16 ) );
  DFF_X1 u0_R1_reg_17 (.CK( clk ) , .D( u0_N48 ) , .Q( u0_R1_17 ) );
  DFF_X1 u0_R1_reg_18 (.CK( clk ) , .D( u0_N49 ) , .Q( u0_R1_18 ) );
  DFF_X1 u0_R1_reg_19 (.CK( clk ) , .D( u0_N50 ) , .Q( u0_R1_19 ) );
  DFF_X1 u0_R1_reg_2 (.CK( clk ) , .D( u0_N33 ) , .Q( u0_R1_2 ) );
  DFF_X1 u0_R1_reg_20 (.CK( clk ) , .D( u0_N51 ) , .Q( u0_R1_20 ) );
  DFF_X1 u0_R1_reg_21 (.CK( clk ) , .D( u0_N52 ) , .Q( u0_R1_21 ) );
  DFF_X1 u0_R1_reg_22 (.CK( clk ) , .D( u0_N53 ) , .Q( u0_R1_22 ) );
  DFF_X1 u0_R1_reg_23 (.CK( clk ) , .D( u0_N54 ) , .Q( u0_R1_23 ) );
  DFF_X1 u0_R1_reg_24 (.CK( clk ) , .D( u0_N55 ) , .Q( u0_R1_24 ) );
  DFF_X1 u0_R1_reg_25 (.CK( clk ) , .D( u0_N56 ) , .Q( u0_R1_25 ) );
  DFF_X1 u0_R1_reg_26 (.CK( clk ) , .D( u0_N57 ) , .Q( u0_R1_26 ) );
  DFF_X1 u0_R1_reg_27 (.CK( clk ) , .D( u0_N58 ) , .Q( u0_R1_27 ) );
  DFF_X1 u0_R1_reg_28 (.CK( clk ) , .D( u0_N59 ) , .Q( u0_R1_28 ) );
  DFF_X1 u0_R1_reg_29 (.CK( clk ) , .D( u0_N60 ) , .Q( u0_R1_29 ) );
  DFF_X1 u0_R1_reg_3 (.CK( clk ) , .D( u0_N34 ) , .Q( u0_R1_3 ) );
  DFF_X1 u0_R1_reg_30 (.CK( clk ) , .D( u0_N61 ) , .Q( u0_R1_30 ) );
  DFF_X1 u0_R1_reg_31 (.CK( clk ) , .D( u0_N62 ) , .Q( u0_R1_31 ) );
  DFF_X1 u0_R1_reg_32 (.CK( clk ) , .D( u0_N63 ) , .Q( u0_R1_32 ) );
  DFF_X1 u0_R1_reg_4 (.CK( clk ) , .D( u0_N35 ) , .Q( u0_R1_4 ) );
  DFF_X1 u0_R1_reg_5 (.CK( clk ) , .D( u0_N36 ) , .Q( u0_R1_5 ) );
  DFF_X1 u0_R1_reg_6 (.CK( clk ) , .D( u0_N37 ) , .Q( u0_R1_6 ) );
  DFF_X1 u0_R1_reg_7 (.CK( clk ) , .D( u0_N38 ) , .Q( u0_R1_7 ) );
  DFF_X1 u0_R1_reg_8 (.CK( clk ) , .D( u0_N39 ) , .Q( u0_R1_8 ) );
  DFF_X1 u0_R1_reg_9 (.CK( clk ) , .D( u0_N40 ) , .Q( u0_R1_9 ) );
  DFF_X1 u0_R2_reg_1 (.CK( clk ) , .D( u0_N64 ) , .Q( u0_R2_1 ) );
  DFF_X1 u0_R2_reg_10 (.CK( clk ) , .D( u0_N73 ) , .Q( u0_R2_10 ) );
  DFF_X1 u0_R2_reg_11 (.CK( clk ) , .D( u0_N74 ) , .Q( u0_R2_11 ) );
  DFF_X1 u0_R2_reg_12 (.CK( clk ) , .D( u0_N75 ) , .Q( u0_R2_12 ) );
  DFF_X1 u0_R2_reg_13 (.CK( clk ) , .D( u0_N76 ) , .Q( u0_R2_13 ) );
  DFF_X1 u0_R2_reg_14 (.CK( clk ) , .D( u0_N77 ) , .Q( u0_R2_14 ) );
  DFF_X1 u0_R2_reg_15 (.CK( clk ) , .D( u0_N78 ) , .Q( u0_R2_15 ) );
  DFF_X1 u0_R2_reg_16 (.CK( clk ) , .D( u0_N79 ) , .Q( u0_R2_16 ) );
  DFF_X1 u0_R2_reg_17 (.CK( clk ) , .D( u0_N80 ) , .Q( u0_R2_17 ) );
  DFF_X1 u0_R2_reg_18 (.CK( clk ) , .D( u0_N81 ) , .Q( u0_R2_18 ) );
  DFF_X1 u0_R2_reg_19 (.CK( clk ) , .D( u0_N82 ) , .Q( u0_R2_19 ) );
  DFF_X1 u0_R2_reg_2 (.CK( clk ) , .D( u0_N65 ) , .Q( u0_R2_2 ) );
  DFF_X1 u0_R2_reg_20 (.CK( clk ) , .D( u0_N83 ) , .Q( u0_R2_20 ) );
  DFF_X1 u0_R2_reg_21 (.CK( clk ) , .D( u0_N84 ) , .Q( u0_R2_21 ) );
  DFF_X1 u0_R2_reg_22 (.CK( clk ) , .D( u0_N85 ) , .Q( u0_R2_22 ) );
  DFF_X1 u0_R2_reg_23 (.CK( clk ) , .D( u0_N86 ) , .Q( u0_R2_23 ) );
  DFF_X1 u0_R2_reg_24 (.CK( clk ) , .D( u0_N87 ) , .Q( u0_R2_24 ) );
  DFF_X1 u0_R2_reg_25 (.CK( clk ) , .D( u0_N88 ) , .Q( u0_R2_25 ) );
  DFF_X1 u0_R2_reg_26 (.CK( clk ) , .D( u0_N89 ) , .Q( u0_R2_26 ) );
  DFF_X1 u0_R2_reg_27 (.CK( clk ) , .D( u0_N90 ) , .Q( u0_R2_27 ) );
  DFF_X1 u0_R2_reg_28 (.CK( clk ) , .D( u0_N91 ) , .Q( u0_R2_28 ) );
  DFF_X1 u0_R2_reg_29 (.CK( clk ) , .D( u0_N92 ) , .Q( u0_R2_29 ) );
  DFF_X1 u0_R2_reg_3 (.CK( clk ) , .D( u0_N66 ) , .Q( u0_R2_3 ) );
  DFF_X1 u0_R2_reg_30 (.CK( clk ) , .D( u0_N93 ) , .Q( u0_R2_30 ) );
  DFF_X1 u0_R2_reg_31 (.CK( clk ) , .D( u0_N94 ) , .Q( u0_R2_31 ) );
  DFF_X1 u0_R2_reg_32 (.CK( clk ) , .D( u0_N95 ) , .Q( u0_R2_32 ) );
  DFF_X1 u0_R2_reg_4 (.CK( clk ) , .D( u0_N67 ) , .Q( u0_R2_4 ) );
  DFF_X1 u0_R2_reg_5 (.CK( clk ) , .D( u0_N68 ) , .Q( u0_R2_5 ) );
  DFF_X1 u0_R2_reg_6 (.CK( clk ) , .D( u0_N69 ) , .Q( u0_R2_6 ) );
  DFF_X1 u0_R2_reg_7 (.CK( clk ) , .D( u0_N70 ) , .Q( u0_R2_7 ) );
  DFF_X1 u0_R2_reg_8 (.CK( clk ) , .D( u0_N71 ) , .Q( u0_R2_8 ) );
  DFF_X1 u0_R2_reg_9 (.CK( clk ) , .D( u0_N72 ) , .Q( u0_R2_9 ) );
  DFF_X1 u0_R3_reg_1 (.CK( clk ) , .D( u0_N96 ) , .Q( u0_R3_1 ) );
  DFF_X1 u0_R3_reg_10 (.CK( clk ) , .D( u0_N105 ) , .Q( u0_R3_10 ) );
  DFF_X1 u0_R3_reg_11 (.CK( clk ) , .D( u0_N106 ) , .Q( u0_R3_11 ) );
  DFF_X1 u0_R3_reg_12 (.CK( clk ) , .D( u0_N107 ) , .Q( u0_R3_12 ) );
  DFF_X1 u0_R3_reg_13 (.CK( clk ) , .D( u0_N108 ) , .Q( u0_R3_13 ) );
  DFF_X1 u0_R3_reg_14 (.CK( clk ) , .D( u0_N109 ) , .Q( u0_R3_14 ) );
  DFF_X1 u0_R3_reg_15 (.CK( clk ) , .D( u0_N110 ) , .Q( u0_R3_15 ) );
  DFF_X1 u0_R3_reg_16 (.CK( clk ) , .D( u0_N111 ) , .Q( u0_R3_16 ) );
  DFF_X1 u0_R3_reg_17 (.CK( clk ) , .D( u0_N112 ) , .Q( u0_R3_17 ) );
  DFF_X1 u0_R3_reg_18 (.CK( clk ) , .D( u0_N113 ) , .Q( u0_R3_18 ) );
  DFF_X1 u0_R3_reg_19 (.CK( clk ) , .D( u0_N114 ) , .Q( u0_R3_19 ) );
  DFF_X1 u0_R3_reg_2 (.CK( clk ) , .D( u0_N97 ) , .Q( u0_R3_2 ) );
  DFF_X1 u0_R3_reg_20 (.CK( clk ) , .D( u0_N115 ) , .Q( u0_R3_20 ) );
  DFF_X1 u0_R3_reg_21 (.CK( clk ) , .D( u0_N116 ) , .Q( u0_R3_21 ) );
  DFF_X1 u0_R3_reg_22 (.CK( clk ) , .D( u0_N117 ) , .Q( u0_R3_22 ) );
  DFF_X1 u0_R3_reg_23 (.CK( clk ) , .D( u0_N118 ) , .Q( u0_R3_23 ) );
  DFF_X1 u0_R3_reg_24 (.CK( clk ) , .D( u0_N119 ) , .Q( u0_R3_24 ) );
  DFF_X1 u0_R3_reg_25 (.CK( clk ) , .D( u0_N120 ) , .Q( u0_R3_25 ) );
  DFF_X1 u0_R3_reg_26 (.CK( clk ) , .D( u0_N121 ) , .Q( u0_R3_26 ) );
  DFF_X1 u0_R3_reg_27 (.CK( clk ) , .D( u0_N122 ) , .Q( u0_R3_27 ) );
  DFF_X1 u0_R3_reg_28 (.CK( clk ) , .D( u0_N123 ) , .Q( u0_R3_28 ) );
  DFF_X1 u0_R3_reg_29 (.CK( clk ) , .D( u0_N124 ) , .Q( u0_R3_29 ) );
  DFF_X1 u0_R3_reg_3 (.CK( clk ) , .D( u0_N98 ) , .Q( u0_R3_3 ) );
  DFF_X1 u0_R3_reg_30 (.CK( clk ) , .D( u0_N125 ) , .Q( u0_R3_30 ) );
  DFF_X1 u0_R3_reg_31 (.CK( clk ) , .D( u0_N126 ) , .Q( u0_R3_31 ) );
  DFF_X1 u0_R3_reg_32 (.CK( clk ) , .D( u0_N127 ) , .Q( u0_R3_32 ) );
  DFF_X1 u0_R3_reg_4 (.CK( clk ) , .D( u0_N99 ) , .Q( u0_R3_4 ) );
  DFF_X1 u0_R3_reg_5 (.CK( clk ) , .D( u0_N100 ) , .Q( u0_R3_5 ) );
  DFF_X1 u0_R3_reg_6 (.CK( clk ) , .D( u0_N101 ) , .Q( u0_R3_6 ) );
  DFF_X1 u0_R3_reg_7 (.CK( clk ) , .D( u0_N102 ) , .Q( u0_R3_7 ) );
  DFF_X1 u0_R3_reg_8 (.CK( clk ) , .D( u0_N103 ) , .Q( u0_R3_8 ) );
  DFF_X1 u0_R3_reg_9 (.CK( clk ) , .D( u0_N104 ) , .Q( u0_R3_9 ) );
  DFF_X1 u0_R4_reg_1 (.CK( clk ) , .D( u0_N128 ) , .Q( u0_R4_1 ) );
  DFF_X1 u0_R4_reg_10 (.CK( clk ) , .D( u0_N137 ) , .Q( u0_R4_10 ) );
  DFF_X1 u0_R4_reg_11 (.CK( clk ) , .D( u0_N138 ) , .Q( u0_R4_11 ) );
  DFF_X1 u0_R4_reg_12 (.CK( clk ) , .D( u0_N139 ) , .Q( u0_R4_12 ) );
  DFF_X1 u0_R4_reg_13 (.CK( clk ) , .D( u0_N140 ) , .Q( u0_R4_13 ) );
  DFF_X1 u0_R4_reg_14 (.CK( clk ) , .D( u0_N141 ) , .Q( u0_R4_14 ) );
  DFF_X1 u0_R4_reg_15 (.CK( clk ) , .D( u0_N142 ) , .Q( u0_R4_15 ) );
  DFF_X1 u0_R4_reg_16 (.CK( clk ) , .D( u0_N143 ) , .Q( u0_R4_16 ) );
  DFF_X1 u0_R4_reg_17 (.CK( clk ) , .D( u0_N144 ) , .Q( u0_R4_17 ) );
  DFF_X1 u0_R4_reg_18 (.CK( clk ) , .D( u0_N145 ) , .Q( u0_R4_18 ) );
  DFF_X1 u0_R4_reg_19 (.CK( clk ) , .D( u0_N146 ) , .Q( u0_R4_19 ) );
  DFF_X1 u0_R4_reg_2 (.CK( clk ) , .D( u0_N129 ) , .Q( u0_R4_2 ) );
  DFF_X1 u0_R4_reg_20 (.CK( clk ) , .D( u0_N147 ) , .Q( u0_R4_20 ) );
  DFF_X1 u0_R4_reg_21 (.CK( clk ) , .D( u0_N148 ) , .Q( u0_R4_21 ) );
  DFF_X1 u0_R4_reg_22 (.CK( clk ) , .D( u0_N149 ) , .Q( u0_R4_22 ) );
  DFF_X1 u0_R4_reg_23 (.CK( clk ) , .D( u0_N150 ) , .Q( u0_R4_23 ) );
  DFF_X1 u0_R4_reg_24 (.CK( clk ) , .D( u0_N151 ) , .Q( u0_R4_24 ) );
  DFF_X1 u0_R4_reg_25 (.CK( clk ) , .D( u0_N152 ) , .Q( u0_R4_25 ) );
  DFF_X1 u0_R4_reg_26 (.CK( clk ) , .D( u0_N153 ) , .Q( u0_R4_26 ) );
  DFF_X1 u0_R4_reg_27 (.CK( clk ) , .D( u0_N154 ) , .Q( u0_R4_27 ) );
  DFF_X1 u0_R4_reg_28 (.CK( clk ) , .D( u0_N155 ) , .Q( u0_R4_28 ) );
  DFF_X1 u0_R4_reg_29 (.CK( clk ) , .D( u0_N156 ) , .Q( u0_R4_29 ) );
  DFF_X1 u0_R4_reg_3 (.CK( clk ) , .D( u0_N130 ) , .Q( u0_R4_3 ) );
  DFF_X1 u0_R4_reg_30 (.CK( clk ) , .D( u0_N157 ) , .Q( u0_R4_30 ) );
  DFF_X1 u0_R4_reg_31 (.CK( clk ) , .D( u0_N158 ) , .Q( u0_R4_31 ) );
  DFF_X1 u0_R4_reg_32 (.CK( clk ) , .D( u0_N159 ) , .Q( u0_R4_32 ) );
  DFF_X1 u0_R4_reg_4 (.CK( clk ) , .D( u0_N131 ) , .Q( u0_R4_4 ) );
  DFF_X1 u0_R4_reg_5 (.CK( clk ) , .D( u0_N132 ) , .Q( u0_R4_5 ) );
  DFF_X1 u0_R4_reg_6 (.CK( clk ) , .D( u0_N133 ) , .Q( u0_R4_6 ) );
  DFF_X1 u0_R4_reg_7 (.CK( clk ) , .D( u0_N134 ) , .Q( u0_R4_7 ) );
  DFF_X1 u0_R4_reg_8 (.CK( clk ) , .D( u0_N135 ) , .Q( u0_R4_8 ) );
  DFF_X1 u0_R4_reg_9 (.CK( clk ) , .D( u0_N136 ) , .Q( u0_R4_9 ) );
  DFF_X1 u0_R5_reg_1 (.CK( clk ) , .D( u0_N160 ) , .Q( u0_R5_1 ) );
  DFF_X1 u0_R5_reg_10 (.CK( clk ) , .D( u0_N169 ) , .Q( u0_R5_10 ) );
  DFF_X1 u0_R5_reg_11 (.CK( clk ) , .D( u0_N170 ) , .Q( u0_R5_11 ) );
  DFF_X1 u0_R5_reg_12 (.CK( clk ) , .D( u0_N171 ) , .Q( u0_R5_12 ) );
  DFF_X1 u0_R5_reg_13 (.CK( clk ) , .D( u0_N172 ) , .Q( u0_R5_13 ) );
  DFF_X1 u0_R5_reg_14 (.CK( clk ) , .D( u0_N173 ) , .Q( u0_R5_14 ) );
  DFF_X1 u0_R5_reg_15 (.CK( clk ) , .D( u0_N174 ) , .Q( u0_R5_15 ) );
  DFF_X1 u0_R5_reg_16 (.CK( clk ) , .D( u0_N175 ) , .Q( u0_R5_16 ) );
  DFF_X1 u0_R5_reg_17 (.CK( clk ) , .D( u0_N176 ) , .Q( u0_R5_17 ) );
  DFF_X1 u0_R5_reg_18 (.CK( clk ) , .D( u0_N177 ) , .Q( u0_R5_18 ) );
  DFF_X1 u0_R5_reg_19 (.CK( clk ) , .D( u0_N178 ) , .Q( u0_R5_19 ) );
  DFF_X1 u0_R5_reg_2 (.CK( clk ) , .D( u0_N161 ) , .Q( u0_R5_2 ) );
  DFF_X1 u0_R5_reg_20 (.CK( clk ) , .D( u0_N179 ) , .Q( u0_R5_20 ) );
  DFF_X1 u0_R5_reg_21 (.CK( clk ) , .D( u0_N180 ) , .Q( u0_R5_21 ) );
  DFF_X1 u0_R5_reg_22 (.CK( clk ) , .D( u0_N181 ) , .Q( u0_R5_22 ) );
  DFF_X1 u0_R5_reg_23 (.CK( clk ) , .D( u0_N182 ) , .Q( u0_R5_23 ) );
  DFF_X1 u0_R5_reg_24 (.CK( clk ) , .D( u0_N183 ) , .Q( u0_R5_24 ) );
  DFF_X1 u0_R5_reg_25 (.CK( clk ) , .D( u0_N184 ) , .Q( u0_R5_25 ) );
  DFF_X1 u0_R5_reg_26 (.CK( clk ) , .D( u0_N185 ) , .Q( u0_R5_26 ) );
  DFF_X1 u0_R5_reg_27 (.CK( clk ) , .D( u0_N186 ) , .Q( u0_R5_27 ) );
  DFF_X1 u0_R5_reg_28 (.CK( clk ) , .D( u0_N187 ) , .Q( u0_R5_28 ) );
  DFF_X1 u0_R5_reg_29 (.CK( clk ) , .D( u0_N188 ) , .Q( u0_R5_29 ) );
  DFF_X1 u0_R5_reg_3 (.CK( clk ) , .D( u0_N162 ) , .Q( u0_R5_3 ) );
  DFF_X1 u0_R5_reg_30 (.CK( clk ) , .D( u0_N189 ) , .Q( u0_R5_30 ) );
  DFF_X1 u0_R5_reg_31 (.CK( clk ) , .D( u0_N190 ) , .Q( u0_R5_31 ) );
  DFF_X1 u0_R5_reg_32 (.CK( clk ) , .D( u0_N191 ) , .Q( u0_R5_32 ) );
  DFF_X1 u0_R5_reg_4 (.CK( clk ) , .D( u0_N163 ) , .Q( u0_R5_4 ) );
  DFF_X1 u0_R5_reg_5 (.CK( clk ) , .D( u0_N164 ) , .Q( u0_R5_5 ) );
  DFF_X1 u0_R5_reg_6 (.CK( clk ) , .D( u0_N165 ) , .Q( u0_R5_6 ) );
  DFF_X1 u0_R5_reg_7 (.CK( clk ) , .D( u0_N166 ) , .Q( u0_R5_7 ) );
  DFF_X1 u0_R5_reg_8 (.CK( clk ) , .D( u0_N167 ) , .Q( u0_R5_8 ) );
  DFF_X1 u0_R5_reg_9 (.CK( clk ) , .D( u0_N168 ) , .Q( u0_R5_9 ) );
  DFF_X1 u0_R6_reg_1 (.CK( clk ) , .D( u0_N192 ) , .Q( u0_R6_1 ) );
  DFF_X1 u0_R6_reg_10 (.CK( clk ) , .D( u0_N201 ) , .Q( u0_R6_10 ) );
  DFF_X1 u0_R6_reg_11 (.CK( clk ) , .D( u0_N202 ) , .Q( u0_R6_11 ) );
  DFF_X1 u0_R6_reg_12 (.CK( clk ) , .D( u0_N203 ) , .Q( u0_R6_12 ) );
  DFF_X1 u0_R6_reg_13 (.CK( clk ) , .D( u0_N204 ) , .Q( u0_R6_13 ) );
  DFF_X1 u0_R6_reg_14 (.CK( clk ) , .D( u0_N205 ) , .Q( u0_R6_14 ) );
  DFF_X1 u0_R6_reg_15 (.CK( clk ) , .D( u0_N206 ) , .Q( u0_R6_15 ) );
  DFF_X1 u0_R6_reg_16 (.CK( clk ) , .D( u0_N207 ) , .Q( u0_R6_16 ) );
  DFF_X1 u0_R6_reg_17 (.CK( clk ) , .D( u0_N208 ) , .Q( u0_R6_17 ) );
  DFF_X1 u0_R6_reg_18 (.CK( clk ) , .D( u0_N209 ) , .Q( u0_R6_18 ) );
  DFF_X1 u0_R6_reg_19 (.CK( clk ) , .D( u0_N210 ) , .Q( u0_R6_19 ) );
  DFF_X1 u0_R6_reg_2 (.CK( clk ) , .D( u0_N193 ) , .Q( u0_R6_2 ) );
  DFF_X1 u0_R6_reg_20 (.CK( clk ) , .D( u0_N211 ) , .Q( u0_R6_20 ) );
  DFF_X1 u0_R6_reg_21 (.CK( clk ) , .D( u0_N212 ) , .Q( u0_R6_21 ) );
  DFF_X1 u0_R6_reg_22 (.CK( clk ) , .D( u0_N213 ) , .Q( u0_R6_22 ) );
  DFF_X1 u0_R6_reg_23 (.CK( clk ) , .D( u0_N214 ) , .Q( u0_R6_23 ) );
  DFF_X1 u0_R6_reg_24 (.CK( clk ) , .D( u0_N215 ) , .Q( u0_R6_24 ) );
  DFF_X1 u0_R6_reg_25 (.CK( clk ) , .D( u0_N216 ) , .Q( u0_R6_25 ) );
  DFF_X1 u0_R6_reg_26 (.CK( clk ) , .D( u0_N217 ) , .Q( u0_R6_26 ) );
  DFF_X1 u0_R6_reg_27 (.CK( clk ) , .D( u0_N218 ) , .Q( u0_R6_27 ) );
  DFF_X1 u0_R6_reg_28 (.CK( clk ) , .D( u0_N219 ) , .Q( u0_R6_28 ) );
  DFF_X1 u0_R6_reg_29 (.CK( clk ) , .D( u0_N220 ) , .Q( u0_R6_29 ) );
  DFF_X1 u0_R6_reg_3 (.CK( clk ) , .D( u0_N194 ) , .Q( u0_R6_3 ) );
  DFF_X1 u0_R6_reg_30 (.CK( clk ) , .D( u0_N221 ) , .Q( u0_R6_30 ) );
  DFF_X1 u0_R6_reg_31 (.CK( clk ) , .D( u0_N222 ) , .Q( u0_R6_31 ) );
  DFF_X1 u0_R6_reg_32 (.CK( clk ) , .D( u0_N223 ) , .Q( u0_R6_32 ) );
  DFF_X1 u0_R6_reg_4 (.CK( clk ) , .D( u0_N195 ) , .Q( u0_R6_4 ) );
  DFF_X1 u0_R6_reg_5 (.CK( clk ) , .D( u0_N196 ) , .Q( u0_R6_5 ) );
  DFF_X1 u0_R6_reg_6 (.CK( clk ) , .D( u0_N197 ) , .Q( u0_R6_6 ) );
  DFF_X1 u0_R6_reg_7 (.CK( clk ) , .D( u0_N198 ) , .Q( u0_R6_7 ) );
  DFF_X1 u0_R6_reg_8 (.CK( clk ) , .D( u0_N199 ) , .Q( u0_R6_8 ) );
  DFF_X1 u0_R6_reg_9 (.CK( clk ) , .D( u0_N200 ) , .Q( u0_R6_9 ) );
  DFF_X1 u0_R7_reg_1 (.CK( clk ) , .D( u0_N224 ) , .Q( u0_R7_1 ) );
  DFF_X1 u0_R7_reg_10 (.CK( clk ) , .D( u0_N233 ) , .Q( u0_R7_10 ) );
  DFF_X1 u0_R7_reg_11 (.CK( clk ) , .D( u0_N234 ) , .Q( u0_R7_11 ) );
  DFF_X1 u0_R7_reg_12 (.CK( clk ) , .D( u0_N235 ) , .Q( u0_R7_12 ) );
  DFF_X1 u0_R7_reg_13 (.CK( clk ) , .D( u0_N236 ) , .Q( u0_R7_13 ) );
  DFF_X1 u0_R7_reg_14 (.CK( clk ) , .D( u0_N237 ) , .Q( u0_R7_14 ) );
  DFF_X1 u0_R7_reg_15 (.CK( clk ) , .D( u0_N238 ) , .Q( u0_R7_15 ) );
  DFF_X1 u0_R7_reg_16 (.CK( clk ) , .D( u0_N239 ) , .Q( u0_R7_16 ) );
  DFF_X1 u0_R7_reg_17 (.CK( clk ) , .D( u0_N240 ) , .Q( u0_R7_17 ) );
  DFF_X1 u0_R7_reg_18 (.CK( clk ) , .D( u0_N241 ) , .Q( u0_R7_18 ) );
  DFF_X1 u0_R7_reg_19 (.CK( clk ) , .D( u0_N242 ) , .Q( u0_R7_19 ) );
  DFF_X1 u0_R7_reg_2 (.CK( clk ) , .D( u0_N225 ) , .Q( u0_R7_2 ) );
  DFF_X1 u0_R7_reg_20 (.CK( clk ) , .D( u0_N243 ) , .Q( u0_R7_20 ) );
  DFF_X1 u0_R7_reg_21 (.CK( clk ) , .D( u0_N244 ) , .Q( u0_R7_21 ) );
  DFF_X1 u0_R7_reg_22 (.CK( clk ) , .D( u0_N245 ) , .Q( u0_R7_22 ) );
  DFF_X1 u0_R7_reg_23 (.CK( clk ) , .D( u0_N246 ) , .Q( u0_R7_23 ) );
  DFF_X1 u0_R7_reg_24 (.CK( clk ) , .D( u0_N247 ) , .Q( u0_R7_24 ) );
  DFF_X1 u0_R7_reg_25 (.CK( clk ) , .D( u0_N248 ) , .Q( u0_R7_25 ) );
  DFF_X1 u0_R7_reg_26 (.CK( clk ) , .D( u0_N249 ) , .Q( u0_R7_26 ) );
  DFF_X1 u0_R7_reg_27 (.CK( clk ) , .D( u0_N250 ) , .Q( u0_R7_27 ) );
  DFF_X1 u0_R7_reg_28 (.CK( clk ) , .D( u0_N251 ) , .Q( u0_R7_28 ) );
  DFF_X1 u0_R7_reg_29 (.CK( clk ) , .D( u0_N252 ) , .Q( u0_R7_29 ) );
  DFF_X1 u0_R7_reg_3 (.CK( clk ) , .D( u0_N226 ) , .Q( u0_R7_3 ) );
  DFF_X1 u0_R7_reg_30 (.CK( clk ) , .D( u0_N253 ) , .Q( u0_R7_30 ) );
  DFF_X1 u0_R7_reg_31 (.CK( clk ) , .D( u0_N254 ) , .Q( u0_R7_31 ) );
  DFF_X1 u0_R7_reg_32 (.CK( clk ) , .D( u0_N255 ) , .Q( u0_R7_32 ) );
  DFF_X1 u0_R7_reg_4 (.CK( clk ) , .D( u0_N227 ) , .Q( u0_R7_4 ) );
  DFF_X1 u0_R7_reg_5 (.CK( clk ) , .D( u0_N228 ) , .Q( u0_R7_5 ) );
  DFF_X1 u0_R7_reg_6 (.CK( clk ) , .D( u0_N229 ) , .Q( u0_R7_6 ) );
  DFF_X1 u0_R7_reg_7 (.CK( clk ) , .D( u0_N230 ) , .Q( u0_R7_7 ) );
  DFF_X1 u0_R7_reg_8 (.CK( clk ) , .D( u0_N231 ) , .Q( u0_R7_8 ) );
  DFF_X1 u0_R7_reg_9 (.CK( clk ) , .D( u0_N232 ) , .Q( u0_R7_9 ) );
  DFF_X1 u0_R8_reg_1 (.CK( clk ) , .D( u0_N256 ) , .Q( u0_R8_1 ) );
  DFF_X1 u0_R8_reg_10 (.CK( clk ) , .D( u0_N265 ) , .Q( u0_R8_10 ) );
  DFF_X1 u0_R8_reg_11 (.CK( clk ) , .D( u0_N266 ) , .Q( u0_R8_11 ) );
  DFF_X1 u0_R8_reg_12 (.CK( clk ) , .D( u0_N267 ) , .Q( u0_R8_12 ) );
  DFF_X1 u0_R8_reg_13 (.CK( clk ) , .D( u0_N268 ) , .Q( u0_R8_13 ) );
  DFF_X1 u0_R8_reg_14 (.CK( clk ) , .D( u0_N269 ) , .Q( u0_R8_14 ) );
  DFF_X1 u0_R8_reg_15 (.CK( clk ) , .D( u0_N270 ) , .Q( u0_R8_15 ) );
  DFF_X1 u0_R8_reg_16 (.CK( clk ) , .D( u0_N271 ) , .Q( u0_R8_16 ) );
  DFF_X1 u0_R8_reg_17 (.CK( clk ) , .D( u0_N272 ) , .Q( u0_R8_17 ) );
  DFF_X1 u0_R8_reg_18 (.CK( clk ) , .D( u0_N273 ) , .Q( u0_R8_18 ) );
  DFF_X1 u0_R8_reg_19 (.CK( clk ) , .D( u0_N274 ) , .Q( u0_R8_19 ) );
  DFF_X1 u0_R8_reg_2 (.CK( clk ) , .D( u0_N257 ) , .Q( u0_R8_2 ) );
  DFF_X1 u0_R8_reg_20 (.CK( clk ) , .D( u0_N275 ) , .Q( u0_R8_20 ) );
  DFF_X1 u0_R8_reg_21 (.CK( clk ) , .D( u0_N276 ) , .Q( u0_R8_21 ) );
  DFF_X1 u0_R8_reg_22 (.CK( clk ) , .D( u0_N277 ) , .Q( u0_R8_22 ) );
  DFF_X1 u0_R8_reg_23 (.CK( clk ) , .D( u0_N278 ) , .Q( u0_R8_23 ) );
  DFF_X1 u0_R8_reg_24 (.CK( clk ) , .D( u0_N279 ) , .Q( u0_R8_24 ) );
  DFF_X1 u0_R8_reg_25 (.CK( clk ) , .D( u0_N280 ) , .Q( u0_R8_25 ) );
  DFF_X1 u0_R8_reg_26 (.CK( clk ) , .D( u0_N281 ) , .Q( u0_R8_26 ) );
  DFF_X1 u0_R8_reg_27 (.CK( clk ) , .D( u0_N282 ) , .Q( u0_R8_27 ) );
  DFF_X1 u0_R8_reg_28 (.CK( clk ) , .D( u0_N283 ) , .Q( u0_R8_28 ) );
  DFF_X1 u0_R8_reg_29 (.CK( clk ) , .D( u0_N284 ) , .Q( u0_R8_29 ) );
  DFF_X1 u0_R8_reg_3 (.CK( clk ) , .D( u0_N258 ) , .Q( u0_R8_3 ) );
  DFF_X1 u0_R8_reg_30 (.CK( clk ) , .D( u0_N285 ) , .Q( u0_R8_30 ) );
  DFF_X1 u0_R8_reg_31 (.CK( clk ) , .D( u0_N286 ) , .Q( u0_R8_31 ) );
  DFF_X1 u0_R8_reg_32 (.CK( clk ) , .D( u0_N287 ) , .Q( u0_R8_32 ) );
  DFF_X1 u0_R8_reg_4 (.CK( clk ) , .D( u0_N259 ) , .Q( u0_R8_4 ) );
  DFF_X1 u0_R8_reg_5 (.CK( clk ) , .D( u0_N260 ) , .Q( u0_R8_5 ) );
  DFF_X1 u0_R8_reg_6 (.CK( clk ) , .D( u0_N261 ) , .Q( u0_R8_6 ) );
  DFF_X1 u0_R8_reg_7 (.CK( clk ) , .D( u0_N262 ) , .Q( u0_R8_7 ) );
  DFF_X1 u0_R8_reg_8 (.CK( clk ) , .D( u0_N263 ) , .Q( u0_R8_8 ) );
  DFF_X1 u0_R8_reg_9 (.CK( clk ) , .D( u0_N264 ) , .Q( u0_R8_9 ) );
  DFF_X1 u0_R9_reg_1 (.CK( clk ) , .D( u0_N288 ) , .Q( u0_R9_1 ) );
  DFF_X1 u0_R9_reg_10 (.CK( clk ) , .D( u0_N297 ) , .Q( u0_R9_10 ) );
  DFF_X1 u0_R9_reg_11 (.CK( clk ) , .D( u0_N298 ) , .Q( u0_R9_11 ) );
  DFF_X1 u0_R9_reg_12 (.CK( clk ) , .D( u0_N299 ) , .Q( u0_R9_12 ) );
  DFF_X1 u0_R9_reg_13 (.CK( clk ) , .D( u0_N300 ) , .Q( u0_R9_13 ) );
  DFF_X1 u0_R9_reg_14 (.CK( clk ) , .D( u0_N301 ) , .Q( u0_R9_14 ) );
  DFF_X1 u0_R9_reg_15 (.CK( clk ) , .D( u0_N302 ) , .Q( u0_R9_15 ) );
  DFF_X1 u0_R9_reg_16 (.CK( clk ) , .D( u0_N303 ) , .Q( u0_R9_16 ) );
  DFF_X1 u0_R9_reg_17 (.CK( clk ) , .D( u0_N304 ) , .Q( u0_R9_17 ) );
  DFF_X1 u0_R9_reg_18 (.CK( clk ) , .D( u0_N305 ) , .Q( u0_R9_18 ) );
  DFF_X1 u0_R9_reg_19 (.CK( clk ) , .D( u0_N306 ) , .Q( u0_R9_19 ) );
  DFF_X1 u0_R9_reg_2 (.CK( clk ) , .D( u0_N289 ) , .Q( u0_R9_2 ) );
  DFF_X1 u0_R9_reg_20 (.CK( clk ) , .D( u0_N307 ) , .Q( u0_R9_20 ) );
  DFF_X1 u0_R9_reg_21 (.CK( clk ) , .D( u0_N308 ) , .Q( u0_R9_21 ) );
  DFF_X1 u0_R9_reg_22 (.CK( clk ) , .D( u0_N309 ) , .Q( u0_R9_22 ) );
  DFF_X1 u0_R9_reg_23 (.CK( clk ) , .D( u0_N310 ) , .Q( u0_R9_23 ) );
  DFF_X1 u0_R9_reg_24 (.CK( clk ) , .D( u0_N311 ) , .Q( u0_R9_24 ) );
  DFF_X1 u0_R9_reg_25 (.CK( clk ) , .D( u0_N312 ) , .Q( u0_R9_25 ) );
  DFF_X1 u0_R9_reg_26 (.CK( clk ) , .D( u0_N313 ) , .Q( u0_R9_26 ) );
  DFF_X1 u0_R9_reg_27 (.CK( clk ) , .D( u0_N314 ) , .Q( u0_R9_27 ) );
  DFF_X1 u0_R9_reg_28 (.CK( clk ) , .D( u0_N315 ) , .Q( u0_R9_28 ) );
  DFF_X1 u0_R9_reg_29 (.CK( clk ) , .D( u0_N316 ) , .Q( u0_R9_29 ) );
  DFF_X1 u0_R9_reg_3 (.CK( clk ) , .D( u0_N290 ) , .Q( u0_R9_3 ) );
  DFF_X1 u0_R9_reg_30 (.CK( clk ) , .D( u0_N317 ) , .Q( u0_R9_30 ) );
  DFF_X1 u0_R9_reg_31 (.CK( clk ) , .D( u0_N318 ) , .Q( u0_R9_31 ) );
  DFF_X1 u0_R9_reg_32 (.CK( clk ) , .D( u0_N319 ) , .Q( u0_R9_32 ) );
  DFF_X1 u0_R9_reg_4 (.CK( clk ) , .D( u0_N291 ) , .Q( u0_R9_4 ) );
  DFF_X1 u0_R9_reg_5 (.CK( clk ) , .D( u0_N292 ) , .Q( u0_R9_5 ) );
  DFF_X1 u0_R9_reg_6 (.CK( clk ) , .D( u0_N293 ) , .Q( u0_R9_6 ) );
  DFF_X1 u0_R9_reg_7 (.CK( clk ) , .D( u0_N294 ) , .Q( u0_R9_7 ) );
  DFF_X1 u0_R9_reg_8 (.CK( clk ) , .D( u0_N295 ) , .Q( u0_R9_8 ) );
  DFF_X1 u0_R9_reg_9 (.CK( clk ) , .D( u0_N296 ) , .Q( u0_R9_9 ) );
  XOR2_X1 u0_U10 (.B( u0_L1_29 ) , .Z( u0_N92 ) , .A( u0_out2_29 ) );
  XOR2_X1 u0_U100 (.B( u0_L12_27 ) , .Z( u0_N442 ) , .A( u0_out13_27 ) );
  XOR2_X1 u0_U101 (.B( u0_L12_26 ) , .Z( u0_N441 ) , .A( u0_out13_26 ) );
  XOR2_X1 u0_U102 (.B( u0_L12_25 ) , .Z( u0_N440 ) , .A( u0_out13_25 ) );
  XOR2_X1 u0_U103 (.B( u0_L0_13 ) , .Z( u0_N44 ) , .A( u0_out1_13 ) );
  XOR2_X1 u0_U104 (.B( u0_L12_24 ) , .Z( u0_N439 ) , .A( u0_out13_24 ) );
  XOR2_X1 u0_U105 (.B( u0_L12_23 ) , .Z( u0_N438 ) , .A( u0_out13_23 ) );
  XOR2_X1 u0_U106 (.B( u0_L12_22 ) , .Z( u0_N437 ) , .A( u0_out13_22 ) );
  XOR2_X1 u0_U107 (.B( u0_L12_21 ) , .Z( u0_N436 ) , .A( u0_out13_21 ) );
  XOR2_X1 u0_U108 (.B( u0_L12_20 ) , .Z( u0_N435 ) , .A( u0_out13_20 ) );
  XOR2_X1 u0_U109 (.B( u0_L12_19 ) , .Z( u0_N434 ) , .A( u0_out13_19 ) );
  XOR2_X1 u0_U11 (.B( u0_L1_28 ) , .Z( u0_N91 ) , .A( u0_out2_28 ) );
  XOR2_X1 u0_U110 (.B( u0_L12_18 ) , .Z( u0_N433 ) , .A( u0_out13_18 ) );
  XOR2_X1 u0_U111 (.B( u0_L12_17 ) , .Z( u0_N432 ) , .A( u0_out13_17 ) );
  XOR2_X1 u0_U112 (.B( u0_L12_16 ) , .Z( u0_N431 ) , .A( u0_out13_16 ) );
  XOR2_X1 u0_U113 (.B( u0_L12_15 ) , .Z( u0_N430 ) , .A( u0_out13_15 ) );
  XOR2_X1 u0_U114 (.B( u0_L0_12 ) , .Z( u0_N43 ) , .A( u0_out1_12 ) );
  XOR2_X1 u0_U115 (.B( u0_L12_14 ) , .Z( u0_N429 ) , .A( u0_out13_14 ) );
  XOR2_X1 u0_U116 (.B( u0_L12_13 ) , .Z( u0_N428 ) , .A( u0_out13_13 ) );
  XOR2_X1 u0_U117 (.B( u0_L12_12 ) , .Z( u0_N427 ) , .A( u0_out13_12 ) );
  XOR2_X1 u0_U118 (.B( u0_L12_11 ) , .Z( u0_N426 ) , .A( u0_out13_11 ) );
  XOR2_X1 u0_U119 (.B( u0_L12_10 ) , .Z( u0_N425 ) , .A( u0_out13_10 ) );
  XOR2_X1 u0_U12 (.B( u0_L1_27 ) , .Z( u0_N90 ) , .A( u0_out2_27 ) );
  XOR2_X1 u0_U120 (.B( u0_L12_9 ) , .Z( u0_N424 ) , .A( u0_out13_9 ) );
  XOR2_X1 u0_U121 (.B( u0_L12_8 ) , .Z( u0_N423 ) , .A( u0_out13_8 ) );
  XOR2_X1 u0_U122 (.B( u0_L12_7 ) , .Z( u0_N422 ) , .A( u0_out13_7 ) );
  XOR2_X1 u0_U123 (.B( u0_L12_6 ) , .Z( u0_N421 ) , .A( u0_out13_6 ) );
  XOR2_X1 u0_U124 (.B( u0_L12_5 ) , .Z( u0_N420 ) , .A( u0_out13_5 ) );
  XOR2_X1 u0_U125 (.B( u0_L0_11 ) , .Z( u0_N42 ) , .A( u0_out1_11 ) );
  XOR2_X1 u0_U126 (.B( u0_L12_4 ) , .Z( u0_N419 ) , .A( u0_out13_4 ) );
  XOR2_X1 u0_U127 (.B( u0_L12_3 ) , .Z( u0_N418 ) , .A( u0_out13_3 ) );
  XOR2_X1 u0_U128 (.B( u0_L12_2 ) , .Z( u0_N417 ) , .A( u0_out13_2 ) );
  XOR2_X1 u0_U129 (.B( u0_L12_1 ) , .Z( u0_N416 ) , .A( u0_out13_1 ) );
  XOR2_X1 u0_U13 (.Z( u0_N9 ) , .B( u0_desIn_r_12 ) , .A( u0_out0_10 ) );
  XOR2_X1 u0_U130 (.B( u0_L11_32 ) , .Z( u0_N415 ) , .A( u0_out12_32 ) );
  XOR2_X1 u0_U131 (.B( u0_L11_31 ) , .Z( u0_N414 ) , .A( u0_out12_31 ) );
  XOR2_X1 u0_U132 (.B( u0_L11_30 ) , .Z( u0_N413 ) , .A( u0_out12_30 ) );
  XOR2_X1 u0_U133 (.B( u0_L11_29 ) , .Z( u0_N412 ) , .A( u0_out12_29 ) );
  XOR2_X1 u0_U134 (.B( u0_L11_28 ) , .Z( u0_N411 ) , .A( u0_out12_28 ) );
  XOR2_X1 u0_U135 (.B( u0_L11_27 ) , .Z( u0_N410 ) , .A( u0_out12_27 ) );
  XOR2_X1 u0_U136 (.B( u0_L0_10 ) , .Z( u0_N41 ) , .A( u0_out1_10 ) );
  XOR2_X1 u0_U137 (.B( u0_L11_26 ) , .Z( u0_N409 ) , .A( u0_out12_26 ) );
  XOR2_X1 u0_U138 (.B( u0_L11_25 ) , .Z( u0_N408 ) , .A( u0_out12_25 ) );
  XOR2_X1 u0_U139 (.B( u0_L11_24 ) , .Z( u0_N407 ) , .A( u0_out12_24 ) );
  XOR2_X1 u0_U14 (.B( u0_L1_26 ) , .Z( u0_N89 ) , .A( u0_out2_26 ) );
  XOR2_X1 u0_U140 (.B( u0_L11_23 ) , .Z( u0_N406 ) , .A( u0_out12_23 ) );
  XOR2_X1 u0_U141 (.B( u0_L11_22 ) , .Z( u0_N405 ) , .A( u0_out12_22 ) );
  XOR2_X1 u0_U142 (.B( u0_L11_21 ) , .Z( u0_N404 ) , .A( u0_out12_21 ) );
  XOR2_X1 u0_U143 (.B( u0_L11_20 ) , .Z( u0_N403 ) , .A( u0_out12_20 ) );
  XOR2_X1 u0_U144 (.B( u0_L11_19 ) , .Z( u0_N402 ) , .A( u0_out12_19 ) );
  XOR2_X1 u0_U145 (.B( u0_L11_18 ) , .Z( u0_N401 ) , .A( u0_out12_18 ) );
  XOR2_X1 u0_U146 (.B( u0_L11_17 ) , .Z( u0_N400 ) , .A( u0_out12_17 ) );
  XOR2_X1 u0_U147 (.B( u0_L0_9 ) , .Z( u0_N40 ) , .A( u0_out1_9 ) );
  XOR2_X1 u0_U148 (.Z( u0_N4 ) , .B( u0_desIn_r_38 ) , .A( u0_out0_5 ) );
  XOR2_X1 u0_U149 (.B( u0_L11_16 ) , .Z( u0_N399 ) , .A( u0_out12_16 ) );
  XOR2_X1 u0_U15 (.B( u0_L1_25 ) , .Z( u0_N88 ) , .A( u0_out2_25 ) );
  XOR2_X1 u0_U150 (.B( u0_L11_15 ) , .Z( u0_N398 ) , .A( u0_out12_15 ) );
  XOR2_X1 u0_U151 (.B( u0_L11_14 ) , .Z( u0_N397 ) , .A( u0_out12_14 ) );
  XOR2_X1 u0_U152 (.B( u0_L11_13 ) , .Z( u0_N396 ) , .A( u0_out12_13 ) );
  XOR2_X1 u0_U153 (.B( u0_L11_12 ) , .Z( u0_N395 ) , .A( u0_out12_12 ) );
  XOR2_X1 u0_U154 (.B( u0_L11_11 ) , .Z( u0_N394 ) , .A( u0_out12_11 ) );
  XOR2_X1 u0_U155 (.B( u0_L11_10 ) , .Z( u0_N393 ) , .A( u0_out12_10 ) );
  XOR2_X1 u0_U156 (.B( u0_L11_9 ) , .Z( u0_N392 ) , .A( u0_out12_9 ) );
  XOR2_X1 u0_U157 (.B( u0_L11_8 ) , .Z( u0_N391 ) , .A( u0_out12_8 ) );
  XOR2_X1 u0_U158 (.B( u0_L11_7 ) , .Z( u0_N390 ) , .A( u0_out12_7 ) );
  XOR2_X1 u0_U159 (.B( u0_L0_8 ) , .Z( u0_N39 ) , .A( u0_out1_8 ) );
  XOR2_X1 u0_U16 (.B( u0_L1_24 ) , .Z( u0_N87 ) , .A( u0_out2_24 ) );
  XOR2_X1 u0_U160 (.B( u0_L11_6 ) , .Z( u0_N389 ) , .A( u0_out12_6 ) );
  XOR2_X1 u0_U161 (.B( u0_L11_5 ) , .Z( u0_N388 ) , .A( u0_out12_5 ) );
  XOR2_X1 u0_U162 (.B( u0_L11_4 ) , .Z( u0_N387 ) , .A( u0_out12_4 ) );
  XOR2_X1 u0_U163 (.B( u0_L11_3 ) , .Z( u0_N386 ) , .A( u0_out12_3 ) );
  XOR2_X1 u0_U164 (.B( u0_L11_2 ) , .Z( u0_N385 ) , .A( u0_out12_2 ) );
  XOR2_X1 u0_U165 (.B( u0_L11_1 ) , .Z( u0_N384 ) , .A( u0_out12_1 ) );
  XOR2_X1 u0_U166 (.B( u0_L10_32 ) , .Z( u0_N383 ) , .A( u0_out11_32 ) );
  XOR2_X1 u0_U167 (.B( u0_L10_31 ) , .Z( u0_N382 ) , .A( u0_out11_31 ) );
  XOR2_X1 u0_U168 (.B( u0_L10_30 ) , .Z( u0_N381 ) , .A( u0_out11_30 ) );
  XOR2_X1 u0_U169 (.B( u0_L10_29 ) , .Z( u0_N380 ) , .A( u0_out11_29 ) );
  XOR2_X1 u0_U17 (.B( u0_L1_23 ) , .Z( u0_N86 ) , .A( u0_out2_23 ) );
  XOR2_X1 u0_U170 (.B( u0_L0_7 ) , .Z( u0_N38 ) , .A( u0_out1_7 ) );
  XOR2_X1 u0_U171 (.B( u0_L10_28 ) , .Z( u0_N379 ) , .A( u0_out11_28 ) );
  XOR2_X1 u0_U172 (.B( u0_L10_27 ) , .Z( u0_N378 ) , .A( u0_out11_27 ) );
  XOR2_X1 u0_U173 (.B( u0_L10_26 ) , .Z( u0_N377 ) , .A( u0_out11_26 ) );
  XOR2_X1 u0_U174 (.B( u0_L10_25 ) , .Z( u0_N376 ) , .A( u0_out11_25 ) );
  XOR2_X1 u0_U175 (.B( u0_L10_24 ) , .Z( u0_N375 ) , .A( u0_out11_24 ) );
  XOR2_X1 u0_U176 (.B( u0_L10_23 ) , .Z( u0_N374 ) , .A( u0_out11_23 ) );
  XOR2_X1 u0_U177 (.B( u0_L10_22 ) , .Z( u0_N373 ) , .A( u0_out11_22 ) );
  XOR2_X1 u0_U178 (.B( u0_L10_21 ) , .Z( u0_N372 ) , .A( u0_out11_21 ) );
  XOR2_X1 u0_U179 (.B( u0_L10_20 ) , .Z( u0_N371 ) , .A( u0_out11_20 ) );
  XOR2_X1 u0_U18 (.B( u0_L1_22 ) , .Z( u0_N85 ) , .A( u0_out2_22 ) );
  XOR2_X1 u0_U180 (.B( u0_L10_19 ) , .Z( u0_N370 ) , .A( u0_out11_19 ) );
  XOR2_X1 u0_U181 (.B( u0_L0_6 ) , .Z( u0_N37 ) , .A( u0_out1_6 ) );
  XOR2_X1 u0_U182 (.B( u0_L10_18 ) , .Z( u0_N369 ) , .A( u0_out11_18 ) );
  XOR2_X1 u0_U183 (.B( u0_L10_17 ) , .Z( u0_N368 ) , .A( u0_out11_17 ) );
  XOR2_X1 u0_U184 (.B( u0_L10_16 ) , .Z( u0_N367 ) , .A( u0_out11_16 ) );
  XOR2_X1 u0_U185 (.B( u0_L10_15 ) , .Z( u0_N366 ) , .A( u0_out11_15 ) );
  XOR2_X1 u0_U186 (.B( u0_L10_14 ) , .Z( u0_N365 ) , .A( u0_out11_14 ) );
  XOR2_X1 u0_U187 (.B( u0_L10_13 ) , .Z( u0_N364 ) , .A( u0_out11_13 ) );
  XOR2_X1 u0_U188 (.B( u0_L10_12 ) , .Z( u0_N363 ) , .A( u0_out11_12 ) );
  XOR2_X1 u0_U189 (.B( u0_L10_11 ) , .Z( u0_N362 ) , .A( u0_out11_11 ) );
  XOR2_X1 u0_U19 (.B( u0_L1_21 ) , .Z( u0_N84 ) , .A( u0_out2_21 ) );
  XOR2_X1 u0_U190 (.B( u0_L10_10 ) , .Z( u0_N361 ) , .A( u0_out11_10 ) );
  XOR2_X1 u0_U191 (.B( u0_L10_9 ) , .Z( u0_N360 ) , .A( u0_out11_9 ) );
  XOR2_X1 u0_U192 (.B( u0_L0_5 ) , .Z( u0_N36 ) , .A( u0_out1_5 ) );
  XOR2_X1 u0_U193 (.B( u0_L10_8 ) , .Z( u0_N359 ) , .A( u0_out11_8 ) );
  XOR2_X1 u0_U194 (.B( u0_L10_7 ) , .Z( u0_N358 ) , .A( u0_out11_7 ) );
  XOR2_X1 u0_U195 (.B( u0_L10_6 ) , .Z( u0_N357 ) , .A( u0_out11_6 ) );
  XOR2_X1 u0_U196 (.B( u0_L10_5 ) , .Z( u0_N356 ) , .A( u0_out11_5 ) );
  XOR2_X1 u0_U197 (.B( u0_L10_4 ) , .Z( u0_N355 ) , .A( u0_out11_4 ) );
  XOR2_X1 u0_U198 (.B( u0_L10_3 ) , .Z( u0_N354 ) , .A( u0_out11_3 ) );
  XOR2_X1 u0_U199 (.B( u0_L10_2 ) , .Z( u0_N353 ) , .A( u0_out11_2 ) );
  XOR2_X1 u0_U20 (.B( u0_L1_20 ) , .Z( u0_N83 ) , .A( u0_out2_20 ) );
  XOR2_X1 u0_U200 (.B( u0_L10_1 ) , .Z( u0_N352 ) , .A( u0_out11_1 ) );
  XOR2_X1 u0_U201 (.B( u0_L9_32 ) , .Z( u0_N351 ) , .A( u0_out10_32 ) );
  XOR2_X1 u0_U202 (.B( u0_L9_31 ) , .Z( u0_N350 ) , .A( u0_out10_31 ) );
  XOR2_X1 u0_U203 (.B( u0_L0_4 ) , .Z( u0_N35 ) , .A( u0_out1_4 ) );
  XOR2_X1 u0_U204 (.B( u0_L9_30 ) , .Z( u0_N349 ) , .A( u0_out10_30 ) );
  XOR2_X1 u0_U205 (.B( u0_L9_29 ) , .Z( u0_N348 ) , .A( u0_out10_29 ) );
  XOR2_X1 u0_U206 (.B( u0_L9_28 ) , .Z( u0_N347 ) , .A( u0_out10_28 ) );
  XOR2_X1 u0_U207 (.B( u0_L9_27 ) , .Z( u0_N346 ) , .A( u0_out10_27 ) );
  XOR2_X1 u0_U208 (.B( u0_L9_26 ) , .Z( u0_N345 ) , .A( u0_out10_26 ) );
  XOR2_X1 u0_U209 (.B( u0_L9_25 ) , .Z( u0_N344 ) , .A( u0_out10_25 ) );
  XOR2_X1 u0_U21 (.B( u0_L1_19 ) , .Z( u0_N82 ) , .A( u0_out2_19 ) );
  XOR2_X1 u0_U210 (.B( u0_L9_24 ) , .Z( u0_N343 ) , .A( u0_out10_24 ) );
  XOR2_X1 u0_U211 (.B( u0_L9_23 ) , .Z( u0_N342 ) , .A( u0_out10_23 ) );
  XOR2_X1 u0_U212 (.B( u0_L9_22 ) , .Z( u0_N341 ) , .A( u0_out10_22 ) );
  XOR2_X1 u0_U213 (.B( u0_L9_21 ) , .Z( u0_N340 ) , .A( u0_out10_21 ) );
  XOR2_X1 u0_U214 (.B( u0_L0_3 ) , .Z( u0_N34 ) , .A( u0_out1_3 ) );
  XOR2_X1 u0_U215 (.B( u0_L9_20 ) , .Z( u0_N339 ) , .A( u0_out10_20 ) );
  XOR2_X1 u0_U216 (.B( u0_L9_19 ) , .Z( u0_N338 ) , .A( u0_out10_19 ) );
  XOR2_X1 u0_U217 (.B( u0_L9_18 ) , .Z( u0_N337 ) , .A( u0_out10_18 ) );
  XOR2_X1 u0_U218 (.B( u0_L9_17 ) , .Z( u0_N336 ) , .A( u0_out10_17 ) );
  XOR2_X1 u0_U219 (.B( u0_L9_16 ) , .Z( u0_N335 ) , .A( u0_out10_16 ) );
  XOR2_X1 u0_U22 (.B( u0_L1_18 ) , .Z( u0_N81 ) , .A( u0_out2_18 ) );
  XOR2_X1 u0_U220 (.B( u0_L9_15 ) , .Z( u0_N334 ) , .A( u0_out10_15 ) );
  XOR2_X1 u0_U221 (.B( u0_L9_14 ) , .Z( u0_N333 ) , .A( u0_out10_14 ) );
  XOR2_X1 u0_U222 (.B( u0_L9_13 ) , .Z( u0_N332 ) , .A( u0_out10_13 ) );
  XOR2_X1 u0_U223 (.B( u0_L9_12 ) , .Z( u0_N331 ) , .A( u0_out10_12 ) );
  XOR2_X1 u0_U224 (.B( u0_L9_11 ) , .Z( u0_N330 ) , .A( u0_out10_11 ) );
  XOR2_X1 u0_U225 (.B( u0_L0_2 ) , .Z( u0_N33 ) , .A( u0_out1_2 ) );
  XOR2_X1 u0_U226 (.B( u0_L9_10 ) , .Z( u0_N329 ) , .A( u0_out10_10 ) );
  XOR2_X1 u0_U227 (.B( u0_L9_9 ) , .Z( u0_N328 ) , .A( u0_out10_9 ) );
  XOR2_X1 u0_U228 (.B( u0_L9_8 ) , .Z( u0_N327 ) , .A( u0_out10_8 ) );
  XOR2_X1 u0_U229 (.B( u0_L9_7 ) , .Z( u0_N326 ) , .A( u0_out10_7 ) );
  XOR2_X1 u0_U23 (.B( u0_L1_17 ) , .Z( u0_N80 ) , .A( u0_out2_17 ) );
  XOR2_X1 u0_U230 (.B( u0_L9_6 ) , .Z( u0_N325 ) , .A( u0_out10_6 ) );
  XOR2_X1 u0_U231 (.B( u0_L9_5 ) , .Z( u0_N324 ) , .A( u0_out10_5 ) );
  XOR2_X1 u0_U232 (.B( u0_L9_4 ) , .Z( u0_N323 ) , .A( u0_out10_4 ) );
  XOR2_X1 u0_U233 (.B( u0_L9_3 ) , .Z( u0_N322 ) , .A( u0_out10_3 ) );
  XOR2_X1 u0_U234 (.B( u0_L9_2 ) , .Z( u0_N321 ) , .A( u0_out10_2 ) );
  XOR2_X1 u0_U235 (.B( u0_L9_1 ) , .Z( u0_N320 ) , .A( u0_out10_1 ) );
  XOR2_X1 u0_U236 (.B( u0_L0_1 ) , .Z( u0_N32 ) , .A( u0_out1_1 ) );
  XOR2_X1 u0_U237 (.B( u0_L8_32 ) , .Z( u0_N319 ) , .A( u0_out9_32 ) );
  XOR2_X1 u0_U238 (.B( u0_L8_31 ) , .Z( u0_N318 ) , .A( u0_out9_31 ) );
  XOR2_X1 u0_U239 (.B( u0_L8_30 ) , .Z( u0_N317 ) , .A( u0_out9_30 ) );
  XOR2_X1 u0_U24 (.Z( u0_N8 ) , .B( u0_desIn_r_4 ) , .A( u0_out0_9 ) );
  XOR2_X1 u0_U240 (.B( u0_L8_29 ) , .Z( u0_N316 ) , .A( u0_out9_29 ) );
  XOR2_X1 u0_U241 (.B( u0_L8_28 ) , .Z( u0_N315 ) , .A( u0_out9_28 ) );
  XOR2_X1 u0_U242 (.B( u0_L8_27 ) , .Z( u0_N314 ) , .A( u0_out9_27 ) );
  XOR2_X1 u0_U243 (.B( u0_L8_26 ) , .Z( u0_N313 ) , .A( u0_out9_26 ) );
  XOR2_X1 u0_U244 (.B( u0_L8_25 ) , .Z( u0_N312 ) , .A( u0_out9_25 ) );
  XOR2_X1 u0_U245 (.B( u0_L8_24 ) , .Z( u0_N311 ) , .A( u0_out9_24 ) );
  XOR2_X1 u0_U246 (.B( u0_L8_23 ) , .Z( u0_N310 ) , .A( u0_out9_23 ) );
  XOR2_X1 u0_U247 (.Z( u0_N31 ) , .B( u0_desIn_r_56 ) , .A( u0_out0_32 ) );
  XOR2_X1 u0_U248 (.B( u0_L8_22 ) , .Z( u0_N309 ) , .A( u0_out9_22 ) );
  XOR2_X1 u0_U249 (.B( u0_L8_21 ) , .Z( u0_N308 ) , .A( u0_out9_21 ) );
  XOR2_X1 u0_U25 (.B( u0_L1_16 ) , .Z( u0_N79 ) , .A( u0_out2_16 ) );
  XOR2_X1 u0_U250 (.B( u0_L8_20 ) , .Z( u0_N307 ) , .A( u0_out9_20 ) );
  XOR2_X1 u0_U251 (.B( u0_L8_19 ) , .Z( u0_N306 ) , .A( u0_out9_19 ) );
  XOR2_X1 u0_U252 (.B( u0_L8_18 ) , .Z( u0_N305 ) , .A( u0_out9_18 ) );
  XOR2_X1 u0_U253 (.B( u0_L8_17 ) , .Z( u0_N304 ) , .A( u0_out9_17 ) );
  XOR2_X1 u0_U254 (.B( u0_L8_16 ) , .Z( u0_N303 ) , .A( u0_out9_16 ) );
  XOR2_X1 u0_U255 (.B( u0_L8_15 ) , .Z( u0_N302 ) , .A( u0_out9_15 ) );
  XOR2_X1 u0_U256 (.B( u0_L8_14 ) , .Z( u0_N301 ) , .A( u0_out9_14 ) );
  XOR2_X1 u0_U257 (.B( u0_L8_13 ) , .Z( u0_N300 ) , .A( u0_out9_13 ) );
  XOR2_X1 u0_U258 (.Z( u0_N30 ) , .B( u0_desIn_r_48 ) , .A( u0_out0_31 ) );
  XOR2_X1 u0_U259 (.Z( u0_N3 ) , .B( u0_desIn_r_30 ) , .A( u0_out0_4 ) );
  XOR2_X1 u0_U26 (.B( u0_L1_15 ) , .Z( u0_N78 ) , .A( u0_out2_15 ) );
  XOR2_X1 u0_U260 (.B( u0_L8_12 ) , .Z( u0_N299 ) , .A( u0_out9_12 ) );
  XOR2_X1 u0_U261 (.B( u0_L8_11 ) , .Z( u0_N298 ) , .A( u0_out9_11 ) );
  XOR2_X1 u0_U262 (.B( u0_L8_10 ) , .Z( u0_N297 ) , .A( u0_out9_10 ) );
  XOR2_X1 u0_U263 (.B( u0_L8_9 ) , .Z( u0_N296 ) , .A( u0_out9_9 ) );
  XOR2_X1 u0_U264 (.B( u0_L8_8 ) , .Z( u0_N295 ) , .A( u0_out9_8 ) );
  XOR2_X1 u0_U265 (.B( u0_L8_7 ) , .Z( u0_N294 ) , .A( u0_out9_7 ) );
  XOR2_X1 u0_U266 (.B( u0_L8_6 ) , .Z( u0_N293 ) , .A( u0_out9_6 ) );
  XOR2_X1 u0_U267 (.B( u0_L8_5 ) , .Z( u0_N292 ) , .A( u0_out9_5 ) );
  XOR2_X1 u0_U268 (.B( u0_L8_4 ) , .Z( u0_N291 ) , .A( u0_out9_4 ) );
  XOR2_X1 u0_U269 (.B( u0_L8_3 ) , .Z( u0_N290 ) , .A( u0_out9_3 ) );
  XOR2_X1 u0_U27 (.B( u0_L1_14 ) , .Z( u0_N77 ) , .A( u0_out2_14 ) );
  XOR2_X1 u0_U270 (.Z( u0_N29 ) , .B( u0_desIn_r_40 ) , .A( u0_out0_30 ) );
  XOR2_X1 u0_U271 (.B( u0_L8_2 ) , .Z( u0_N289 ) , .A( u0_out9_2 ) );
  XOR2_X1 u0_U272 (.B( u0_L8_1 ) , .Z( u0_N288 ) , .A( u0_out9_1 ) );
  XOR2_X1 u0_U273 (.B( u0_L7_32 ) , .Z( u0_N287 ) , .A( u0_out8_32 ) );
  XOR2_X1 u0_U274 (.B( u0_L7_31 ) , .Z( u0_N286 ) , .A( u0_out8_31 ) );
  XOR2_X1 u0_U275 (.B( u0_L7_30 ) , .Z( u0_N285 ) , .A( u0_out8_30 ) );
  XOR2_X1 u0_U276 (.B( u0_L7_29 ) , .Z( u0_N284 ) , .A( u0_out8_29 ) );
  XOR2_X1 u0_U277 (.B( u0_L7_28 ) , .Z( u0_N283 ) , .A( u0_out8_28 ) );
  XOR2_X1 u0_U278 (.B( u0_L7_27 ) , .Z( u0_N282 ) , .A( u0_out8_27 ) );
  XOR2_X1 u0_U279 (.B( u0_L7_26 ) , .Z( u0_N281 ) , .A( u0_out8_26 ) );
  XOR2_X1 u0_U28 (.B( u0_L1_13 ) , .Z( u0_N76 ) , .A( u0_out2_13 ) );
  XOR2_X1 u0_U280 (.B( u0_L7_25 ) , .Z( u0_N280 ) , .A( u0_out8_25 ) );
  XOR2_X1 u0_U281 (.Z( u0_N28 ) , .B( u0_desIn_r_32 ) , .A( u0_out0_29 ) );
  XOR2_X1 u0_U282 (.B( u0_L7_24 ) , .Z( u0_N279 ) , .A( u0_out8_24 ) );
  XOR2_X1 u0_U283 (.B( u0_L7_23 ) , .Z( u0_N278 ) , .A( u0_out8_23 ) );
  XOR2_X1 u0_U284 (.B( u0_L7_22 ) , .Z( u0_N277 ) , .A( u0_out8_22 ) );
  XOR2_X1 u0_U285 (.B( u0_L7_21 ) , .Z( u0_N276 ) , .A( u0_out8_21 ) );
  XOR2_X1 u0_U286 (.B( u0_L7_20 ) , .Z( u0_N275 ) , .A( u0_out8_20 ) );
  XOR2_X1 u0_U287 (.B( u0_L7_19 ) , .Z( u0_N274 ) , .A( u0_out8_19 ) );
  XOR2_X1 u0_U288 (.B( u0_L7_18 ) , .Z( u0_N273 ) , .A( u0_out8_18 ) );
  XOR2_X1 u0_U289 (.B( u0_L7_17 ) , .Z( u0_N272 ) , .A( u0_out8_17 ) );
  XOR2_X1 u0_U29 (.B( u0_L1_12 ) , .Z( u0_N75 ) , .A( u0_out2_12 ) );
  XOR2_X1 u0_U290 (.B( u0_L7_16 ) , .Z( u0_N271 ) , .A( u0_out8_16 ) );
  XOR2_X1 u0_U291 (.B( u0_L7_15 ) , .Z( u0_N270 ) , .A( u0_out8_15 ) );
  XOR2_X1 u0_U292 (.Z( u0_N27 ) , .B( u0_desIn_r_24 ) , .A( u0_out0_28 ) );
  XOR2_X1 u0_U293 (.B( u0_L7_14 ) , .Z( u0_N269 ) , .A( u0_out8_14 ) );
  XOR2_X1 u0_U294 (.B( u0_L7_13 ) , .Z( u0_N268 ) , .A( u0_out8_13 ) );
  XOR2_X1 u0_U295 (.B( u0_L7_12 ) , .Z( u0_N267 ) , .A( u0_out8_12 ) );
  XOR2_X1 u0_U296 (.B( u0_L7_11 ) , .Z( u0_N266 ) , .A( u0_out8_11 ) );
  XOR2_X1 u0_U297 (.B( u0_L7_10 ) , .Z( u0_N265 ) , .A( u0_out8_10 ) );
  XOR2_X1 u0_U298 (.B( u0_L7_9 ) , .Z( u0_N264 ) , .A( u0_out8_9 ) );
  XOR2_X1 u0_U299 (.B( u0_L7_8 ) , .Z( u0_N263 ) , .A( u0_out8_8 ) );
  XOR2_X1 u0_U3 (.B( u0_L2_4 ) , .Z( u0_N99 ) , .A( u0_out3_4 ) );
  XOR2_X1 u0_U30 (.B( u0_L1_11 ) , .Z( u0_N74 ) , .A( u0_out2_11 ) );
  XOR2_X1 u0_U300 (.B( u0_L7_7 ) , .Z( u0_N262 ) , .A( u0_out8_7 ) );
  XOR2_X1 u0_U301 (.B( u0_L7_6 ) , .Z( u0_N261 ) , .A( u0_out8_6 ) );
  XOR2_X1 u0_U302 (.B( u0_L7_5 ) , .Z( u0_N260 ) , .A( u0_out8_5 ) );
  XOR2_X1 u0_U303 (.Z( u0_N26 ) , .B( u0_desIn_r_16 ) , .A( u0_out0_27 ) );
  XOR2_X1 u0_U304 (.B( u0_L7_4 ) , .Z( u0_N259 ) , .A( u0_out8_4 ) );
  XOR2_X1 u0_U305 (.B( u0_L7_3 ) , .Z( u0_N258 ) , .A( u0_out8_3 ) );
  XOR2_X1 u0_U306 (.B( u0_L7_2 ) , .Z( u0_N257 ) , .A( u0_out8_2 ) );
  XOR2_X1 u0_U307 (.B( u0_L7_1 ) , .Z( u0_N256 ) , .A( u0_out8_1 ) );
  XOR2_X1 u0_U308 (.B( u0_L6_32 ) , .Z( u0_N255 ) , .A( u0_out7_32 ) );
  XOR2_X1 u0_U309 (.B( u0_L6_31 ) , .Z( u0_N254 ) , .A( u0_out7_31 ) );
  XOR2_X1 u0_U31 (.B( u0_L1_10 ) , .Z( u0_N73 ) , .A( u0_out2_10 ) );
  XOR2_X1 u0_U310 (.B( u0_L6_30 ) , .Z( u0_N253 ) , .A( u0_out7_30 ) );
  XOR2_X1 u0_U311 (.B( u0_L6_29 ) , .Z( u0_N252 ) , .A( u0_out7_29 ) );
  XOR2_X1 u0_U312 (.B( u0_L6_28 ) , .Z( u0_N251 ) , .A( u0_out7_28 ) );
  XOR2_X1 u0_U313 (.B( u0_L6_27 ) , .Z( u0_N250 ) , .A( u0_out7_27 ) );
  XOR2_X1 u0_U314 (.Z( u0_N25 ) , .B( u0_desIn_r_8 ) , .A( u0_out0_26 ) );
  XOR2_X1 u0_U315 (.B( u0_L6_26 ) , .Z( u0_N249 ) , .A( u0_out7_26 ) );
  XOR2_X1 u0_U316 (.B( u0_L6_25 ) , .Z( u0_N248 ) , .A( u0_out7_25 ) );
  XOR2_X1 u0_U317 (.B( u0_L6_24 ) , .Z( u0_N247 ) , .A( u0_out7_24 ) );
  XOR2_X1 u0_U318 (.B( u0_L6_23 ) , .Z( u0_N246 ) , .A( u0_out7_23 ) );
  XOR2_X1 u0_U319 (.B( u0_L6_22 ) , .Z( u0_N245 ) , .A( u0_out7_22 ) );
  XOR2_X1 u0_U32 (.B( u0_L1_9 ) , .Z( u0_N72 ) , .A( u0_out2_9 ) );
  XOR2_X1 u0_U320 (.B( u0_L6_21 ) , .Z( u0_N244 ) , .A( u0_out7_21 ) );
  XOR2_X1 u0_U321 (.B( u0_L6_20 ) , .Z( u0_N243 ) , .A( u0_out7_20 ) );
  XOR2_X1 u0_U322 (.B( u0_L6_19 ) , .Z( u0_N242 ) , .A( u0_out7_19 ) );
  XOR2_X1 u0_U323 (.B( u0_L6_18 ) , .Z( u0_N241 ) , .A( u0_out7_18 ) );
  XOR2_X1 u0_U324 (.B( u0_L6_17 ) , .Z( u0_N240 ) , .A( u0_out7_17 ) );
  XOR2_X1 u0_U325 (.Z( u0_N24 ) , .B( u0_desIn_r_0 ) , .A( u0_out0_25 ) );
  XOR2_X1 u0_U326 (.B( u0_L6_16 ) , .Z( u0_N239 ) , .A( u0_out7_16 ) );
  XOR2_X1 u0_U327 (.B( u0_L6_15 ) , .Z( u0_N238 ) , .A( u0_out7_15 ) );
  XOR2_X1 u0_U328 (.B( u0_L6_14 ) , .Z( u0_N237 ) , .A( u0_out7_14 ) );
  XOR2_X1 u0_U329 (.B( u0_L6_13 ) , .Z( u0_N236 ) , .A( u0_out7_13 ) );
  XOR2_X1 u0_U33 (.B( u0_L1_8 ) , .Z( u0_N71 ) , .A( u0_out2_8 ) );
  XOR2_X1 u0_U330 (.B( u0_L6_12 ) , .Z( u0_N235 ) , .A( u0_out7_12 ) );
  XOR2_X1 u0_U331 (.B( u0_L6_11 ) , .Z( u0_N234 ) , .A( u0_out7_11 ) );
  XOR2_X1 u0_U332 (.B( u0_L6_10 ) , .Z( u0_N233 ) , .A( u0_out7_10 ) );
  XOR2_X1 u0_U333 (.B( u0_L6_9 ) , .Z( u0_N232 ) , .A( u0_out7_9 ) );
  XOR2_X1 u0_U334 (.B( u0_L6_8 ) , .Z( u0_N231 ) , .A( u0_out7_8 ) );
  XOR2_X1 u0_U335 (.B( u0_L6_7 ) , .Z( u0_N230 ) , .A( u0_out7_7 ) );
  XOR2_X1 u0_U336 (.Z( u0_N23 ) , .B( u0_desIn_r_58 ) , .A( u0_out0_24 ) );
  XOR2_X1 u0_U337 (.B( u0_L6_6 ) , .Z( u0_N229 ) , .A( u0_out7_6 ) );
  XOR2_X1 u0_U338 (.B( u0_L6_5 ) , .Z( u0_N228 ) , .A( u0_out7_5 ) );
  XOR2_X1 u0_U339 (.B( u0_L6_4 ) , .Z( u0_N227 ) , .A( u0_out7_4 ) );
  XOR2_X1 u0_U34 (.B( u0_L1_7 ) , .Z( u0_N70 ) , .A( u0_out2_7 ) );
  XOR2_X1 u0_U340 (.B( u0_L6_3 ) , .Z( u0_N226 ) , .A( u0_out7_3 ) );
  XOR2_X1 u0_U341 (.B( u0_L6_2 ) , .Z( u0_N225 ) , .A( u0_out7_2 ) );
  XOR2_X1 u0_U342 (.B( u0_L6_1 ) , .Z( u0_N224 ) , .A( u0_out7_1 ) );
  XOR2_X1 u0_U343 (.B( u0_L5_32 ) , .Z( u0_N223 ) , .A( u0_out6_32 ) );
  XOR2_X1 u0_U344 (.B( u0_L5_31 ) , .Z( u0_N222 ) , .A( u0_out6_31 ) );
  XOR2_X1 u0_U345 (.B( u0_L5_30 ) , .Z( u0_N221 ) , .A( u0_out6_30 ) );
  XOR2_X1 u0_U346 (.B( u0_L5_29 ) , .Z( u0_N220 ) , .A( u0_out6_29 ) );
  XOR2_X1 u0_U347 (.Z( u0_N22 ) , .B( u0_desIn_r_50 ) , .A( u0_out0_23 ) );
  XOR2_X1 u0_U348 (.B( u0_L5_28 ) , .Z( u0_N219 ) , .A( u0_out6_28 ) );
  XOR2_X1 u0_U349 (.B( u0_L5_27 ) , .Z( u0_N218 ) , .A( u0_out6_27 ) );
  XOR2_X1 u0_U35 (.Z( u0_N7 ) , .B( u0_desIn_r_62 ) , .A( u0_out0_8 ) );
  XOR2_X1 u0_U350 (.B( u0_L5_26 ) , .Z( u0_N217 ) , .A( u0_out6_26 ) );
  XOR2_X1 u0_U351 (.B( u0_L5_25 ) , .Z( u0_N216 ) , .A( u0_out6_25 ) );
  XOR2_X1 u0_U352 (.B( u0_L5_24 ) , .Z( u0_N215 ) , .A( u0_out6_24 ) );
  XOR2_X1 u0_U353 (.B( u0_L5_23 ) , .Z( u0_N214 ) , .A( u0_out6_23 ) );
  XOR2_X1 u0_U354 (.B( u0_L5_22 ) , .Z( u0_N213 ) , .A( u0_out6_22 ) );
  XOR2_X1 u0_U355 (.B( u0_L5_21 ) , .Z( u0_N212 ) , .A( u0_out6_21 ) );
  XOR2_X1 u0_U356 (.B( u0_L5_20 ) , .Z( u0_N211 ) , .A( u0_out6_20 ) );
  XOR2_X1 u0_U357 (.B( u0_L5_19 ) , .Z( u0_N210 ) , .A( u0_out6_19 ) );
  XOR2_X1 u0_U358 (.Z( u0_N21 ) , .B( u0_desIn_r_42 ) , .A( u0_out0_22 ) );
  XOR2_X1 u0_U359 (.B( u0_L5_18 ) , .Z( u0_N209 ) , .A( u0_out6_18 ) );
  XOR2_X1 u0_U36 (.B( u0_L1_6 ) , .Z( u0_N69 ) , .A( u0_out2_6 ) );
  XOR2_X1 u0_U360 (.B( u0_L5_17 ) , .Z( u0_N208 ) , .A( u0_out6_17 ) );
  XOR2_X1 u0_U361 (.B( u0_L5_16 ) , .Z( u0_N207 ) , .A( u0_out6_16 ) );
  XOR2_X1 u0_U362 (.B( u0_L5_15 ) , .Z( u0_N206 ) , .A( u0_out6_15 ) );
  XOR2_X1 u0_U363 (.B( u0_L5_14 ) , .Z( u0_N205 ) , .A( u0_out6_14 ) );
  XOR2_X1 u0_U364 (.B( u0_L5_13 ) , .Z( u0_N204 ) , .A( u0_out6_13 ) );
  XOR2_X1 u0_U365 (.B( u0_L5_12 ) , .Z( u0_N203 ) , .A( u0_out6_12 ) );
  XOR2_X1 u0_U366 (.B( u0_L5_11 ) , .Z( u0_N202 ) , .A( u0_out6_11 ) );
  XOR2_X1 u0_U367 (.B( u0_L5_10 ) , .Z( u0_N201 ) , .A( u0_out6_10 ) );
  XOR2_X1 u0_U368 (.B( u0_L5_9 ) , .Z( u0_N200 ) , .A( u0_out6_9 ) );
  XOR2_X1 u0_U369 (.Z( u0_N20 ) , .B( u0_desIn_r_34 ) , .A( u0_out0_21 ) );
  XOR2_X1 u0_U37 (.B( u0_L1_5 ) , .Z( u0_N68 ) , .A( u0_out2_5 ) );
  XOR2_X1 u0_U370 (.Z( u0_N2 ) , .B( u0_desIn_r_22 ) , .A( u0_out0_3 ) );
  XOR2_X1 u0_U371 (.B( u0_L5_8 ) , .Z( u0_N199 ) , .A( u0_out6_8 ) );
  XOR2_X1 u0_U372 (.B( u0_L5_7 ) , .Z( u0_N198 ) , .A( u0_out6_7 ) );
  XOR2_X1 u0_U373 (.B( u0_L5_6 ) , .Z( u0_N197 ) , .A( u0_out6_6 ) );
  XOR2_X1 u0_U374 (.B( u0_L5_5 ) , .Z( u0_N196 ) , .A( u0_out6_5 ) );
  XOR2_X1 u0_U375 (.B( u0_L5_4 ) , .Z( u0_N195 ) , .A( u0_out6_4 ) );
  XOR2_X1 u0_U376 (.B( u0_L5_3 ) , .Z( u0_N194 ) , .A( u0_out6_3 ) );
  XOR2_X1 u0_U377 (.B( u0_L5_2 ) , .Z( u0_N193 ) , .A( u0_out6_2 ) );
  XOR2_X1 u0_U378 (.B( u0_L5_1 ) , .Z( u0_N192 ) , .A( u0_out6_1 ) );
  XOR2_X1 u0_U379 (.B( u0_L4_32 ) , .Z( u0_N191 ) , .A( u0_out5_32 ) );
  XOR2_X1 u0_U38 (.B( u0_L1_4 ) , .Z( u0_N67 ) , .A( u0_out2_4 ) );
  XOR2_X1 u0_U380 (.B( u0_L4_31 ) , .Z( u0_N190 ) , .A( u0_out5_31 ) );
  XOR2_X1 u0_U381 (.Z( u0_N19 ) , .B( u0_desIn_r_26 ) , .A( u0_out0_20 ) );
  XOR2_X1 u0_U382 (.B( u0_L4_30 ) , .Z( u0_N189 ) , .A( u0_out5_30 ) );
  XOR2_X1 u0_U383 (.B( u0_L4_29 ) , .Z( u0_N188 ) , .A( u0_out5_29 ) );
  XOR2_X1 u0_U384 (.B( u0_L4_28 ) , .Z( u0_N187 ) , .A( u0_out5_28 ) );
  XOR2_X1 u0_U385 (.B( u0_L4_27 ) , .Z( u0_N186 ) , .A( u0_out5_27 ) );
  XOR2_X1 u0_U386 (.B( u0_L4_26 ) , .Z( u0_N185 ) , .A( u0_out5_26 ) );
  XOR2_X1 u0_U387 (.B( u0_L4_25 ) , .Z( u0_N184 ) , .A( u0_out5_25 ) );
  XOR2_X1 u0_U388 (.B( u0_L4_24 ) , .Z( u0_N183 ) , .A( u0_out5_24 ) );
  XOR2_X1 u0_U389 (.B( u0_L4_23 ) , .Z( u0_N182 ) , .A( u0_out5_23 ) );
  XOR2_X1 u0_U39 (.B( u0_L1_3 ) , .Z( u0_N66 ) , .A( u0_out2_3 ) );
  XOR2_X1 u0_U390 (.B( u0_L4_22 ) , .Z( u0_N181 ) , .A( u0_out5_22 ) );
  XOR2_X1 u0_U391 (.B( u0_L4_21 ) , .Z( u0_N180 ) , .A( u0_out5_21 ) );
  XOR2_X1 u0_U392 (.Z( u0_N18 ) , .B( u0_desIn_r_18 ) , .A( u0_out0_19 ) );
  XOR2_X1 u0_U393 (.B( u0_L4_20 ) , .Z( u0_N179 ) , .A( u0_out5_20 ) );
  XOR2_X1 u0_U394 (.B( u0_L4_19 ) , .Z( u0_N178 ) , .A( u0_out5_19 ) );
  XOR2_X1 u0_U395 (.B( u0_L4_18 ) , .Z( u0_N177 ) , .A( u0_out5_18 ) );
  XOR2_X1 u0_U396 (.B( u0_L4_17 ) , .Z( u0_N176 ) , .A( u0_out5_17 ) );
  XOR2_X1 u0_U397 (.B( u0_L4_16 ) , .Z( u0_N175 ) , .A( u0_out5_16 ) );
  XOR2_X1 u0_U398 (.B( u0_L4_15 ) , .Z( u0_N174 ) , .A( u0_out5_15 ) );
  XOR2_X1 u0_U399 (.B( u0_L4_14 ) , .Z( u0_N173 ) , .A( u0_out5_14 ) );
  XOR2_X1 u0_U4 (.B( u0_L2_3 ) , .Z( u0_N98 ) , .A( u0_out3_3 ) );
  XOR2_X1 u0_U40 (.B( u0_L1_2 ) , .Z( u0_N65 ) , .A( u0_out2_2 ) );
  XOR2_X1 u0_U400 (.B( u0_L4_13 ) , .Z( u0_N172 ) , .A( u0_out5_13 ) );
  XOR2_X1 u0_U401 (.B( u0_L4_12 ) , .Z( u0_N171 ) , .A( u0_out5_12 ) );
  XOR2_X1 u0_U402 (.B( u0_L4_11 ) , .Z( u0_N170 ) , .A( u0_out5_11 ) );
  XOR2_X1 u0_U403 (.Z( u0_N17 ) , .B( u0_desIn_r_10 ) , .A( u0_out0_18 ) );
  XOR2_X1 u0_U404 (.B( u0_L4_10 ) , .Z( u0_N169 ) , .A( u0_out5_10 ) );
  XOR2_X1 u0_U405 (.B( u0_L4_9 ) , .Z( u0_N168 ) , .A( u0_out5_9 ) );
  XOR2_X1 u0_U406 (.B( u0_L4_8 ) , .Z( u0_N167 ) , .A( u0_out5_8 ) );
  XOR2_X1 u0_U407 (.B( u0_L4_7 ) , .Z( u0_N166 ) , .A( u0_out5_7 ) );
  XOR2_X1 u0_U408 (.B( u0_L4_6 ) , .Z( u0_N165 ) , .A( u0_out5_6 ) );
  XOR2_X1 u0_U409 (.B( u0_L4_5 ) , .Z( u0_N164 ) , .A( u0_out5_5 ) );
  XOR2_X1 u0_U41 (.B( u0_L1_1 ) , .Z( u0_N64 ) , .A( u0_out2_1 ) );
  XOR2_X1 u0_U410 (.B( u0_L4_4 ) , .Z( u0_N163 ) , .A( u0_out5_4 ) );
  XOR2_X1 u0_U411 (.B( u0_L4_3 ) , .Z( u0_N162 ) , .A( u0_out5_3 ) );
  XOR2_X1 u0_U412 (.B( u0_L4_2 ) , .Z( u0_N161 ) , .A( u0_out5_2 ) );
  XOR2_X1 u0_U413 (.B( u0_L4_1 ) , .Z( u0_N160 ) , .A( u0_out5_1 ) );
  XOR2_X1 u0_U414 (.Z( u0_N16 ) , .B( u0_desIn_r_2 ) , .A( u0_out0_17 ) );
  XOR2_X1 u0_U415 (.B( u0_L3_32 ) , .Z( u0_N159 ) , .A( u0_out4_32 ) );
  XOR2_X1 u0_U416 (.B( u0_L3_31 ) , .Z( u0_N158 ) , .A( u0_out4_31 ) );
  XOR2_X1 u0_U417 (.B( u0_L3_30 ) , .Z( u0_N157 ) , .A( u0_out4_30 ) );
  XOR2_X1 u0_U418 (.B( u0_L3_29 ) , .Z( u0_N156 ) , .A( u0_out4_29 ) );
  XOR2_X1 u0_U419 (.B( u0_L3_28 ) , .Z( u0_N155 ) , .A( u0_out4_28 ) );
  XOR2_X1 u0_U42 (.B( u0_L0_32 ) , .Z( u0_N63 ) , .A( u0_out1_32 ) );
  XOR2_X1 u0_U420 (.B( u0_L3_27 ) , .Z( u0_N154 ) , .A( u0_out4_27 ) );
  XOR2_X1 u0_U421 (.B( u0_L3_26 ) , .Z( u0_N153 ) , .A( u0_out4_26 ) );
  XOR2_X1 u0_U422 (.B( u0_L3_25 ) , .Z( u0_N152 ) , .A( u0_out4_25 ) );
  XOR2_X1 u0_U423 (.B( u0_L3_24 ) , .Z( u0_N151 ) , .A( u0_out4_24 ) );
  XOR2_X1 u0_U424 (.B( u0_L3_23 ) , .Z( u0_N150 ) , .A( u0_out4_23 ) );
  XOR2_X1 u0_U425 (.Z( u0_N15 ) , .B( u0_desIn_r_60 ) , .A( u0_out0_16 ) );
  XOR2_X1 u0_U426 (.B( u0_L3_22 ) , .Z( u0_N149 ) , .A( u0_out4_22 ) );
  XOR2_X1 u0_U427 (.B( u0_L3_21 ) , .Z( u0_N148 ) , .A( u0_out4_21 ) );
  XOR2_X1 u0_U428 (.B( u0_L3_20 ) , .Z( u0_N147 ) , .A( u0_out4_20 ) );
  XOR2_X1 u0_U429 (.B( u0_L3_19 ) , .Z( u0_N146 ) , .A( u0_out4_19 ) );
  XOR2_X1 u0_U43 (.B( u0_L0_31 ) , .Z( u0_N62 ) , .A( u0_out1_31 ) );
  XOR2_X1 u0_U430 (.B( u0_L3_18 ) , .Z( u0_N145 ) , .A( u0_out4_18 ) );
  XOR2_X1 u0_U431 (.B( u0_L3_17 ) , .Z( u0_N144 ) , .A( u0_out4_17 ) );
  XOR2_X1 u0_U432 (.B( u0_L3_16 ) , .Z( u0_N143 ) , .A( u0_out4_16 ) );
  XOR2_X1 u0_U433 (.B( u0_L3_15 ) , .Z( u0_N142 ) , .A( u0_out4_15 ) );
  XOR2_X1 u0_U434 (.B( u0_L3_14 ) , .Z( u0_N141 ) , .A( u0_out4_14 ) );
  XOR2_X1 u0_U435 (.B( u0_L3_13 ) , .Z( u0_N140 ) , .A( u0_out4_13 ) );
  XOR2_X1 u0_U436 (.Z( u0_N14 ) , .B( u0_desIn_r_52 ) , .A( u0_out0_15 ) );
  XOR2_X1 u0_U437 (.B( u0_L3_12 ) , .Z( u0_N139 ) , .A( u0_out4_12 ) );
  XOR2_X1 u0_U438 (.B( u0_L3_11 ) , .Z( u0_N138 ) , .A( u0_out4_11 ) );
  XOR2_X1 u0_U439 (.B( u0_L3_10 ) , .Z( u0_N137 ) , .A( u0_out4_10 ) );
  XOR2_X1 u0_U44 (.B( u0_L0_30 ) , .Z( u0_N61 ) , .A( u0_out1_30 ) );
  XOR2_X1 u0_U440 (.B( u0_L3_9 ) , .Z( u0_N136 ) , .A( u0_out4_9 ) );
  XOR2_X1 u0_U441 (.B( u0_L3_8 ) , .Z( u0_N135 ) , .A( u0_out4_8 ) );
  XOR2_X1 u0_U442 (.B( u0_L3_7 ) , .Z( u0_N134 ) , .A( u0_out4_7 ) );
  XOR2_X1 u0_U443 (.B( u0_L3_6 ) , .Z( u0_N133 ) , .A( u0_out4_6 ) );
  XOR2_X1 u0_U444 (.B( u0_L3_5 ) , .Z( u0_N132 ) , .A( u0_out4_5 ) );
  XOR2_X1 u0_U445 (.B( u0_L3_4 ) , .Z( u0_N131 ) , .A( u0_out4_4 ) );
  XOR2_X1 u0_U446 (.B( u0_L3_3 ) , .Z( u0_N130 ) , .A( u0_out4_3 ) );
  XOR2_X1 u0_U447 (.Z( u0_N13 ) , .B( u0_desIn_r_44 ) , .A( u0_out0_14 ) );
  XOR2_X1 u0_U448 (.B( u0_L3_2 ) , .Z( u0_N129 ) , .A( u0_out4_2 ) );
  XOR2_X1 u0_U449 (.B( u0_L3_1 ) , .Z( u0_N128 ) , .A( u0_out4_1 ) );
  XOR2_X1 u0_U45 (.B( u0_L0_29 ) , .Z( u0_N60 ) , .A( u0_out1_29 ) );
  XOR2_X1 u0_U450 (.B( u0_L2_32 ) , .Z( u0_N127 ) , .A( u0_out3_32 ) );
  XOR2_X1 u0_U451 (.B( u0_L2_31 ) , .Z( u0_N126 ) , .A( u0_out3_31 ) );
  XOR2_X1 u0_U452 (.B( u0_L2_30 ) , .Z( u0_N125 ) , .A( u0_out3_30 ) );
  XOR2_X1 u0_U453 (.B( u0_L2_29 ) , .Z( u0_N124 ) , .A( u0_out3_29 ) );
  XOR2_X1 u0_U454 (.B( u0_L2_28 ) , .Z( u0_N123 ) , .A( u0_out3_28 ) );
  XOR2_X1 u0_U455 (.B( u0_L2_27 ) , .Z( u0_N122 ) , .A( u0_out3_27 ) );
  XOR2_X1 u0_U456 (.B( u0_L2_26 ) , .Z( u0_N121 ) , .A( u0_out3_26 ) );
  XOR2_X1 u0_U457 (.B( u0_L2_25 ) , .Z( u0_N120 ) , .A( u0_out3_25 ) );
  XOR2_X1 u0_U458 (.Z( u0_N12 ) , .B( u0_desIn_r_36 ) , .A( u0_out0_13 ) );
  XOR2_X1 u0_U459 (.B( u0_L2_24 ) , .Z( u0_N119 ) , .A( u0_out3_24 ) );
  XOR2_X1 u0_U46 (.Z( u0_N6 ) , .B( u0_desIn_r_54 ) , .A( u0_out0_7 ) );
  XOR2_X1 u0_U460 (.B( u0_L2_23 ) , .Z( u0_N118 ) , .A( u0_out3_23 ) );
  XOR2_X1 u0_U461 (.B( u0_L2_22 ) , .Z( u0_N117 ) , .A( u0_out3_22 ) );
  XOR2_X1 u0_U462 (.B( u0_L2_21 ) , .Z( u0_N116 ) , .A( u0_out3_21 ) );
  XOR2_X1 u0_U463 (.B( u0_L2_20 ) , .Z( u0_N115 ) , .A( u0_out3_20 ) );
  XOR2_X1 u0_U464 (.B( u0_L2_19 ) , .Z( u0_N114 ) , .A( u0_out3_19 ) );
  XOR2_X1 u0_U465 (.B( u0_L2_18 ) , .Z( u0_N113 ) , .A( u0_out3_18 ) );
  XOR2_X1 u0_U466 (.B( u0_L2_17 ) , .Z( u0_N112 ) , .A( u0_out3_17 ) );
  XOR2_X1 u0_U467 (.B( u0_L2_16 ) , .Z( u0_N111 ) , .A( u0_out3_16 ) );
  XOR2_X1 u0_U468 (.B( u0_L2_15 ) , .Z( u0_N110 ) , .A( u0_out3_15 ) );
  XOR2_X1 u0_U469 (.Z( u0_N11 ) , .B( u0_desIn_r_28 ) , .A( u0_out0_12 ) );
  XOR2_X1 u0_U47 (.B( u0_L0_28 ) , .Z( u0_N59 ) , .A( u0_out1_28 ) );
  XOR2_X1 u0_U470 (.B( u0_L2_14 ) , .Z( u0_N109 ) , .A( u0_out3_14 ) );
  XOR2_X1 u0_U471 (.B( u0_L2_13 ) , .Z( u0_N108 ) , .A( u0_out3_13 ) );
  XOR2_X1 u0_U472 (.B( u0_L2_12 ) , .Z( u0_N107 ) , .A( u0_out3_12 ) );
  XOR2_X1 u0_U473 (.B( u0_L2_11 ) , .Z( u0_N106 ) , .A( u0_out3_11 ) );
  XOR2_X1 u0_U474 (.B( u0_L2_10 ) , .Z( u0_N105 ) , .A( u0_out3_10 ) );
  XOR2_X1 u0_U475 (.B( u0_L2_9 ) , .Z( u0_N104 ) , .A( u0_out3_9 ) );
  XOR2_X1 u0_U476 (.B( u0_L2_8 ) , .Z( u0_N103 ) , .A( u0_out3_8 ) );
  XOR2_X1 u0_U477 (.B( u0_L2_7 ) , .Z( u0_N102 ) , .A( u0_out3_7 ) );
  XOR2_X1 u0_U478 (.B( u0_L2_6 ) , .Z( u0_N101 ) , .A( u0_out3_6 ) );
  XOR2_X1 u0_U479 (.B( u0_L2_5 ) , .Z( u0_N100 ) , .A( u0_out3_5 ) );
  XOR2_X1 u0_U48 (.B( u0_L0_27 ) , .Z( u0_N58 ) , .A( u0_out1_27 ) );
  XOR2_X1 u0_U480 (.Z( u0_N10 ) , .B( u0_desIn_r_20 ) , .A( u0_out0_11 ) );
  XOR2_X1 u0_U481 (.Z( u0_N1 ) , .B( u0_desIn_r_14 ) , .A( u0_out0_2 ) );
  XOR2_X1 u0_U482 (.Z( u0_N0 ) , .B( u0_desIn_r_6 ) , .A( u0_out0_1 ) );
  XOR2_X1 u0_U483 (.Z( u0_FP_9 ) , .B( u0_L14_9 ) , .A( u0_out15_9 ) );
  XOR2_X1 u0_U484 (.Z( u0_FP_8 ) , .B( u0_L14_8 ) , .A( u0_out15_8 ) );
  XOR2_X1 u0_U485 (.Z( u0_FP_7 ) , .B( u0_L14_7 ) , .A( u0_out15_7 ) );
  XOR2_X1 u0_U486 (.Z( u0_FP_6 ) , .B( u0_L14_6 ) , .A( u0_out15_6 ) );
  XOR2_X1 u0_U487 (.Z( u0_FP_5 ) , .B( u0_L14_5 ) , .A( u0_out15_5 ) );
  XOR2_X1 u0_U488 (.Z( u0_FP_4 ) , .B( u0_L14_4 ) , .A( u0_out15_4 ) );
  XOR2_X1 u0_U489 (.Z( u0_FP_3 ) , .B( u0_L14_3 ) , .A( u0_out15_3 ) );
  XOR2_X1 u0_U49 (.B( u0_L0_26 ) , .Z( u0_N57 ) , .A( u0_out1_26 ) );
  XOR2_X1 u0_U490 (.Z( u0_FP_32 ) , .B( u0_L14_32 ) , .A( u0_out15_32 ) );
  XOR2_X1 u0_U491 (.Z( u0_FP_31 ) , .B( u0_L14_31 ) , .A( u0_out15_31 ) );
  XOR2_X1 u0_U492 (.Z( u0_FP_30 ) , .B( u0_L14_30 ) , .A( u0_out15_30 ) );
  XOR2_X1 u0_U493 (.Z( u0_FP_2 ) , .B( u0_L14_2 ) , .A( u0_out15_2 ) );
  XOR2_X1 u0_U494 (.Z( u0_FP_29 ) , .B( u0_L14_29 ) , .A( u0_out15_29 ) );
  XOR2_X1 u0_U495 (.Z( u0_FP_28 ) , .B( u0_L14_28 ) , .A( u0_out15_28 ) );
  XOR2_X1 u0_U496 (.Z( u0_FP_27 ) , .B( u0_L14_27 ) , .A( u0_out15_27 ) );
  XOR2_X1 u0_U497 (.Z( u0_FP_26 ) , .B( u0_L14_26 ) , .A( u0_out15_26 ) );
  XOR2_X1 u0_U498 (.Z( u0_FP_25 ) , .B( u0_L14_25 ) , .A( u0_out15_25 ) );
  XOR2_X1 u0_U499 (.Z( u0_FP_24 ) , .B( u0_L14_24 ) , .A( u0_out15_24 ) );
  XOR2_X1 u0_U5 (.B( u0_L2_2 ) , .Z( u0_N97 ) , .A( u0_out3_2 ) );
  XOR2_X1 u0_U50 (.B( u0_L0_25 ) , .Z( u0_N56 ) , .A( u0_out1_25 ) );
  XOR2_X1 u0_U500 (.Z( u0_FP_23 ) , .B( u0_L14_23 ) , .A( u0_out15_23 ) );
  XOR2_X1 u0_U501 (.Z( u0_FP_22 ) , .B( u0_L14_22 ) , .A( u0_out15_22 ) );
  XOR2_X1 u0_U502 (.Z( u0_FP_21 ) , .B( u0_L14_21 ) , .A( u0_out15_21 ) );
  XOR2_X1 u0_U503 (.Z( u0_FP_20 ) , .B( u0_L14_20 ) , .A( u0_out15_20 ) );
  XOR2_X1 u0_U504 (.Z( u0_FP_1 ) , .B( u0_L14_1 ) , .A( u0_out15_1 ) );
  XOR2_X1 u0_U505 (.Z( u0_FP_19 ) , .B( u0_L14_19 ) , .A( u0_out15_19 ) );
  XOR2_X1 u0_U506 (.Z( u0_FP_18 ) , .B( u0_L14_18 ) , .A( u0_out15_18 ) );
  XOR2_X1 u0_U507 (.Z( u0_FP_17 ) , .B( u0_L14_17 ) , .A( u0_out15_17 ) );
  XOR2_X1 u0_U508 (.Z( u0_FP_16 ) , .B( u0_L14_16 ) , .A( u0_out15_16 ) );
  XOR2_X1 u0_U509 (.Z( u0_FP_15 ) , .B( u0_L14_15 ) , .A( u0_out15_15 ) );
  XOR2_X1 u0_U51 (.B( u0_L0_24 ) , .Z( u0_N55 ) , .A( u0_out1_24 ) );
  XOR2_X1 u0_U510 (.Z( u0_FP_14 ) , .B( u0_L14_14 ) , .A( u0_out15_14 ) );
  XOR2_X1 u0_U511 (.Z( u0_FP_13 ) , .B( u0_L14_13 ) , .A( u0_out15_13 ) );
  XOR2_X1 u0_U512 (.Z( u0_FP_12 ) , .B( u0_L14_12 ) , .A( u0_out15_12 ) );
  XOR2_X1 u0_U513 (.Z( u0_FP_11 ) , .B( u0_L14_11 ) , .A( u0_out15_11 ) );
  XOR2_X1 u0_U514 (.Z( u0_FP_10 ) , .B( u0_L14_10 ) , .A( u0_out15_10 ) );
  XOR2_X1 u0_U52 (.B( u0_L0_23 ) , .Z( u0_N54 ) , .A( u0_out1_23 ) );
  XOR2_X1 u0_U53 (.B( u0_L0_22 ) , .Z( u0_N53 ) , .A( u0_out1_22 ) );
  XOR2_X1 u0_U54 (.B( u0_L0_21 ) , .Z( u0_N52 ) , .A( u0_out1_21 ) );
  XOR2_X1 u0_U55 (.B( u0_L0_20 ) , .Z( u0_N51 ) , .A( u0_out1_20 ) );
  XOR2_X1 u0_U56 (.B( u0_L0_19 ) , .Z( u0_N50 ) , .A( u0_out1_19 ) );
  XOR2_X1 u0_U57 (.Z( u0_N5 ) , .B( u0_desIn_r_46 ) , .A( u0_out0_6 ) );
  XOR2_X1 u0_U58 (.B( u0_L0_18 ) , .Z( u0_N49 ) , .A( u0_out1_18 ) );
  XOR2_X1 u0_U59 (.B( u0_L0_17 ) , .Z( u0_N48 ) , .A( u0_out1_17 ) );
  XOR2_X1 u0_U6 (.B( u0_L2_1 ) , .Z( u0_N96 ) , .A( u0_out3_1 ) );
  XOR2_X1 u0_U60 (.B( u0_L13_32 ) , .Z( u0_N479 ) , .A( u0_out14_32 ) );
  XOR2_X1 u0_U61 (.B( u0_L13_31 ) , .Z( u0_N478 ) , .A( u0_out14_31 ) );
  XOR2_X1 u0_U62 (.B( u0_L13_30 ) , .Z( u0_N477 ) , .A( u0_out14_30 ) );
  XOR2_X1 u0_U63 (.B( u0_L13_29 ) , .Z( u0_N476 ) , .A( u0_out14_29 ) );
  XOR2_X1 u0_U64 (.B( u0_L13_28 ) , .Z( u0_N475 ) , .A( u0_out14_28 ) );
  XOR2_X1 u0_U65 (.B( u0_L13_27 ) , .Z( u0_N474 ) , .A( u0_out14_27 ) );
  XOR2_X1 u0_U66 (.B( u0_L13_26 ) , .Z( u0_N473 ) , .A( u0_out14_26 ) );
  XOR2_X1 u0_U67 (.B( u0_L13_25 ) , .Z( u0_N472 ) , .A( u0_out14_25 ) );
  XOR2_X1 u0_U68 (.B( u0_L13_24 ) , .Z( u0_N471 ) , .A( u0_out14_24 ) );
  XOR2_X1 u0_U69 (.B( u0_L13_23 ) , .Z( u0_N470 ) , .A( u0_out14_23 ) );
  XOR2_X1 u0_U7 (.B( u0_L1_32 ) , .Z( u0_N95 ) , .A( u0_out2_32 ) );
  XOR2_X1 u0_U70 (.B( u0_L0_16 ) , .Z( u0_N47 ) , .A( u0_out1_16 ) );
  XOR2_X1 u0_U71 (.B( u0_L13_22 ) , .Z( u0_N469 ) , .A( u0_out14_22 ) );
  XOR2_X1 u0_U72 (.B( u0_L13_21 ) , .Z( u0_N468 ) , .A( u0_out14_21 ) );
  XOR2_X1 u0_U73 (.B( u0_L13_20 ) , .Z( u0_N467 ) , .A( u0_out14_20 ) );
  XOR2_X1 u0_U74 (.B( u0_L13_19 ) , .Z( u0_N466 ) , .A( u0_out14_19 ) );
  XOR2_X1 u0_U75 (.B( u0_L13_18 ) , .Z( u0_N465 ) , .A( u0_out14_18 ) );
  XOR2_X1 u0_U76 (.B( u0_L13_17 ) , .Z( u0_N464 ) , .A( u0_out14_17 ) );
  XOR2_X1 u0_U77 (.B( u0_L13_16 ) , .Z( u0_N463 ) , .A( u0_out14_16 ) );
  XOR2_X1 u0_U78 (.B( u0_L13_15 ) , .Z( u0_N462 ) , .A( u0_out14_15 ) );
  XOR2_X1 u0_U79 (.B( u0_L13_14 ) , .Z( u0_N461 ) , .A( u0_out14_14 ) );
  XOR2_X1 u0_U8 (.B( u0_L1_31 ) , .Z( u0_N94 ) , .A( u0_out2_31 ) );
  XOR2_X1 u0_U80 (.B( u0_L13_13 ) , .Z( u0_N460 ) , .A( u0_out14_13 ) );
  XOR2_X1 u0_U81 (.B( u0_L0_15 ) , .Z( u0_N46 ) , .A( u0_out1_15 ) );
  XOR2_X1 u0_U82 (.B( u0_L13_12 ) , .Z( u0_N459 ) , .A( u0_out14_12 ) );
  XOR2_X1 u0_U83 (.B( u0_L13_11 ) , .Z( u0_N458 ) , .A( u0_out14_11 ) );
  XOR2_X1 u0_U84 (.B( u0_L13_10 ) , .Z( u0_N457 ) , .A( u0_out14_10 ) );
  XOR2_X1 u0_U85 (.B( u0_L13_9 ) , .Z( u0_N456 ) , .A( u0_out14_9 ) );
  XOR2_X1 u0_U86 (.B( u0_L13_8 ) , .Z( u0_N455 ) , .A( u0_out14_8 ) );
  XOR2_X1 u0_U87 (.B( u0_L13_7 ) , .Z( u0_N454 ) , .A( u0_out14_7 ) );
  XOR2_X1 u0_U88 (.B( u0_L13_6 ) , .Z( u0_N453 ) , .A( u0_out14_6 ) );
  XOR2_X1 u0_U89 (.B( u0_L13_5 ) , .Z( u0_N452 ) , .A( u0_out14_5 ) );
  XOR2_X1 u0_U9 (.B( u0_L1_30 ) , .Z( u0_N93 ) , .A( u0_out2_30 ) );
  XOR2_X1 u0_U90 (.B( u0_L13_4 ) , .Z( u0_N451 ) , .A( u0_out14_4 ) );
  XOR2_X1 u0_U91 (.B( u0_L13_3 ) , .Z( u0_N450 ) , .A( u0_out14_3 ) );
  XOR2_X1 u0_U92 (.B( u0_L0_14 ) , .Z( u0_N45 ) , .A( u0_out1_14 ) );
  XOR2_X1 u0_U93 (.B( u0_L13_2 ) , .Z( u0_N449 ) , .A( u0_out14_2 ) );
  XOR2_X1 u0_U94 (.B( u0_L13_1 ) , .Z( u0_N448 ) , .A( u0_out14_1 ) );
  XOR2_X1 u0_U95 (.B( u0_L12_32 ) , .Z( u0_N447 ) , .A( u0_out13_32 ) );
  XOR2_X1 u0_U96 (.B( u0_L12_31 ) , .Z( u0_N446 ) , .A( u0_out13_31 ) );
  XOR2_X1 u0_U97 (.B( u0_L12_30 ) , .Z( u0_N445 ) , .A( u0_out13_30 ) );
  XOR2_X1 u0_U98 (.B( u0_L12_29 ) , .Z( u0_N444 ) , .A( u0_out13_29 ) );
  XOR2_X1 u0_U99 (.B( u0_L12_28 ) , .Z( u0_N443 ) , .A( u0_out13_28 ) );
  DFF_X1 u0_desIn_r_reg_0 (.CK( clk ) , .D( desIn[0] ) , .Q( u0_desIn_r_0 ) );
  DFF_X1 u0_desIn_r_reg_1 (.CK( clk ) , .D( desIn[1] ) , .Q( u0_desIn_r_1 ) );
  DFF_X1 u0_desIn_r_reg_10 (.CK( clk ) , .D( desIn[10] ) , .Q( u0_desIn_r_10 ) );
  DFF_X1 u0_desIn_r_reg_11 (.CK( clk ) , .D( desIn[11] ) , .Q( u0_desIn_r_11 ) );
  DFF_X1 u0_desIn_r_reg_12 (.CK( clk ) , .D( desIn[12] ) , .Q( u0_desIn_r_12 ) );
  DFF_X1 u0_desIn_r_reg_13 (.CK( clk ) , .D( desIn[13] ) , .Q( u0_desIn_r_13 ) );
  DFF_X1 u0_desIn_r_reg_14 (.CK( clk ) , .D( desIn[14] ) , .Q( u0_desIn_r_14 ) );
  DFF_X1 u0_desIn_r_reg_15 (.CK( clk ) , .D( desIn[15] ) , .Q( u0_desIn_r_15 ) );
  DFF_X1 u0_desIn_r_reg_16 (.CK( clk ) , .D( desIn[16] ) , .Q( u0_desIn_r_16 ) );
  DFF_X1 u0_desIn_r_reg_17 (.CK( clk ) , .D( desIn[17] ) , .Q( u0_desIn_r_17 ) );
  DFF_X1 u0_desIn_r_reg_18 (.CK( clk ) , .D( desIn[18] ) , .Q( u0_desIn_r_18 ) );
  DFF_X1 u0_desIn_r_reg_19 (.CK( clk ) , .D( desIn[19] ) , .Q( u0_desIn_r_19 ) );
  DFF_X1 u0_desIn_r_reg_2 (.CK( clk ) , .D( desIn[2] ) , .Q( u0_desIn_r_2 ) );
  DFF_X1 u0_desIn_r_reg_20 (.CK( clk ) , .D( desIn[20] ) , .Q( u0_desIn_r_20 ) );
  DFF_X1 u0_desIn_r_reg_21 (.CK( clk ) , .D( desIn[21] ) , .Q( u0_desIn_r_21 ) );
  DFF_X1 u0_desIn_r_reg_22 (.CK( clk ) , .D( desIn[22] ) , .Q( u0_desIn_r_22 ) );
  DFF_X1 u0_desIn_r_reg_23 (.CK( clk ) , .D( desIn[23] ) , .Q( u0_desIn_r_23 ) );
  DFF_X1 u0_desIn_r_reg_24 (.CK( clk ) , .D( desIn[24] ) , .Q( u0_desIn_r_24 ) );
  DFF_X1 u0_desIn_r_reg_25 (.CK( clk ) , .D( desIn[25] ) , .Q( u0_desIn_r_25 ) );
  DFF_X1 u0_desIn_r_reg_26 (.CK( clk ) , .D( desIn[26] ) , .Q( u0_desIn_r_26 ) );
  DFF_X1 u0_desIn_r_reg_27 (.CK( clk ) , .D( desIn[27] ) , .Q( u0_desIn_r_27 ) );
  DFF_X1 u0_desIn_r_reg_28 (.CK( clk ) , .D( desIn[28] ) , .Q( u0_desIn_r_28 ) );
  DFF_X1 u0_desIn_r_reg_29 (.CK( clk ) , .D( desIn[29] ) , .Q( u0_desIn_r_29 ) );
  DFF_X1 u0_desIn_r_reg_3 (.CK( clk ) , .D( desIn[3] ) , .Q( u0_desIn_r_3 ) );
  DFF_X1 u0_desIn_r_reg_30 (.CK( clk ) , .D( desIn[30] ) , .Q( u0_desIn_r_30 ) );
  DFF_X1 u0_desIn_r_reg_31 (.CK( clk ) , .D( desIn[31] ) , .Q( u0_desIn_r_31 ) );
  DFF_X1 u0_desIn_r_reg_32 (.CK( clk ) , .D( desIn[32] ) , .Q( u0_desIn_r_32 ) );
  DFF_X1 u0_desIn_r_reg_33 (.CK( clk ) , .D( desIn[33] ) , .Q( u0_desIn_r_33 ) );
  DFF_X1 u0_desIn_r_reg_34 (.CK( clk ) , .D( desIn[34] ) , .Q( u0_desIn_r_34 ) );
  DFF_X1 u0_desIn_r_reg_35 (.CK( clk ) , .D( desIn[35] ) , .Q( u0_desIn_r_35 ) );
  DFF_X1 u0_desIn_r_reg_36 (.CK( clk ) , .D( desIn[36] ) , .Q( u0_desIn_r_36 ) );
  DFF_X1 u0_desIn_r_reg_37 (.CK( clk ) , .D( desIn[37] ) , .Q( u0_desIn_r_37 ) );
  DFF_X1 u0_desIn_r_reg_38 (.CK( clk ) , .D( desIn[38] ) , .Q( u0_desIn_r_38 ) );
  DFF_X1 u0_desIn_r_reg_39 (.CK( clk ) , .D( desIn[39] ) , .Q( u0_desIn_r_39 ) );
  DFF_X1 u0_desIn_r_reg_4 (.CK( clk ) , .D( desIn[4] ) , .Q( u0_desIn_r_4 ) );
  DFF_X1 u0_desIn_r_reg_40 (.CK( clk ) , .D( desIn[40] ) , .Q( u0_desIn_r_40 ) );
  DFF_X1 u0_desIn_r_reg_41 (.CK( clk ) , .D( desIn[41] ) , .Q( u0_desIn_r_41 ) );
  DFF_X1 u0_desIn_r_reg_42 (.CK( clk ) , .D( desIn[42] ) , .Q( u0_desIn_r_42 ) );
  DFF_X1 u0_desIn_r_reg_43 (.CK( clk ) , .D( desIn[43] ) , .Q( u0_desIn_r_43 ) );
  DFF_X1 u0_desIn_r_reg_44 (.CK( clk ) , .D( desIn[44] ) , .Q( u0_desIn_r_44 ) );
  DFF_X1 u0_desIn_r_reg_45 (.CK( clk ) , .D( desIn[45] ) , .Q( u0_desIn_r_45 ) );
  DFF_X1 u0_desIn_r_reg_46 (.CK( clk ) , .D( desIn[46] ) , .Q( u0_desIn_r_46 ) );
  DFF_X1 u0_desIn_r_reg_47 (.CK( clk ) , .D( desIn[47] ) , .Q( u0_desIn_r_47 ) );
  DFF_X1 u0_desIn_r_reg_48 (.CK( clk ) , .D( desIn[48] ) , .Q( u0_desIn_r_48 ) );
  DFF_X1 u0_desIn_r_reg_49 (.CK( clk ) , .D( desIn[49] ) , .Q( u0_desIn_r_49 ) );
  DFF_X1 u0_desIn_r_reg_5 (.CK( clk ) , .D( desIn[5] ) , .Q( u0_desIn_r_5 ) );
  DFF_X1 u0_desIn_r_reg_50 (.CK( clk ) , .D( desIn[50] ) , .Q( u0_desIn_r_50 ) );
  DFF_X1 u0_desIn_r_reg_51 (.CK( clk ) , .D( desIn[51] ) , .Q( u0_desIn_r_51 ) );
  DFF_X1 u0_desIn_r_reg_52 (.CK( clk ) , .D( desIn[52] ) , .Q( u0_desIn_r_52 ) );
  DFF_X1 u0_desIn_r_reg_53 (.CK( clk ) , .D( desIn[53] ) , .Q( u0_desIn_r_53 ) );
  DFF_X1 u0_desIn_r_reg_54 (.CK( clk ) , .D( desIn[54] ) , .Q( u0_desIn_r_54 ) );
  DFF_X1 u0_desIn_r_reg_55 (.CK( clk ) , .D( desIn[55] ) , .Q( u0_desIn_r_55 ) );
  DFF_X1 u0_desIn_r_reg_56 (.CK( clk ) , .D( desIn[56] ) , .Q( u0_desIn_r_56 ) );
  DFF_X1 u0_desIn_r_reg_57 (.CK( clk ) , .D( desIn[57] ) , .Q( u0_desIn_r_57 ) );
  DFF_X1 u0_desIn_r_reg_58 (.CK( clk ) , .D( desIn[58] ) , .Q( u0_desIn_r_58 ) );
  DFF_X1 u0_desIn_r_reg_59 (.CK( clk ) , .D( desIn[59] ) , .Q( u0_desIn_r_59 ) );
  DFF_X1 u0_desIn_r_reg_6 (.CK( clk ) , .D( desIn[6] ) , .Q( u0_desIn_r_6 ) );
  DFF_X1 u0_desIn_r_reg_60 (.CK( clk ) , .D( desIn[60] ) , .Q( u0_desIn_r_60 ) );
  DFF_X1 u0_desIn_r_reg_61 (.CK( clk ) , .D( desIn[61] ) , .Q( u0_desIn_r_61 ) );
  DFF_X1 u0_desIn_r_reg_62 (.CK( clk ) , .D( desIn[62] ) , .Q( u0_desIn_r_62 ) );
  DFF_X1 u0_desIn_r_reg_63 (.CK( clk ) , .D( desIn[63] ) , .Q( u0_desIn_r_63 ) );
  DFF_X1 u0_desIn_r_reg_7 (.CK( clk ) , .D( desIn[7] ) , .Q( u0_desIn_r_7 ) );
  DFF_X1 u0_desIn_r_reg_8 (.CK( clk ) , .D( desIn[8] ) , .Q( u0_desIn_r_8 ) );
  DFF_X1 u0_desIn_r_reg_9 (.CK( clk ) , .D( desIn[9] ) , .Q( u0_desIn_r_9 ) );
  DFF_X1 u0_desOut_reg_0 (.CK( clk ) , .Q( stage1_out_0 ) , .D( u0_FP_25 ) );
  DFF_X1 u0_desOut_reg_1 (.CK( clk ) , .Q( stage1_out_1 ) , .D( u0_FP_57 ) );
  DFF_X1 u0_desOut_reg_10 (.CK( clk ) , .Q( stage1_out_10 ) , .D( u0_FP_18 ) );
  DFF_X1 u0_desOut_reg_11 (.CK( clk ) , .Q( stage1_out_11 ) , .D( u0_FP_50 ) );
  DFF_X1 u0_desOut_reg_12 (.CK( clk ) , .Q( stage1_out_12 ) , .D( u0_FP_10 ) );
  DFF_X1 u0_desOut_reg_13 (.CK( clk ) , .Q( stage1_out_13 ) , .D( u0_FP_42 ) );
  DFF_X1 u0_desOut_reg_14 (.CK( clk ) , .Q( stage1_out_14 ) , .D( u0_FP_2 ) );
  DFF_X1 u0_desOut_reg_15 (.CK( clk ) , .Q( stage1_out_15 ) , .D( u0_FP_34 ) );
  DFF_X1 u0_desOut_reg_16 (.CK( clk ) , .Q( stage1_out_16 ) , .D( u0_FP_27 ) );
  DFF_X1 u0_desOut_reg_17 (.CK( clk ) , .Q( stage1_out_17 ) , .D( u0_FP_59 ) );
  DFF_X1 u0_desOut_reg_18 (.CK( clk ) , .Q( stage1_out_18 ) , .D( u0_FP_19 ) );
  DFF_X1 u0_desOut_reg_19 (.CK( clk ) , .Q( stage1_out_19 ) , .D( u0_FP_51 ) );
  DFF_X1 u0_desOut_reg_2 (.CK( clk ) , .Q( stage1_out_2 ) , .D( u0_FP_17 ) );
  DFF_X1 u0_desOut_reg_20 (.CK( clk ) , .Q( stage1_out_20 ) , .D( u0_FP_11 ) );
  DFF_X1 u0_desOut_reg_21 (.CK( clk ) , .Q( stage1_out_21 ) , .D( u0_FP_43 ) );
  DFF_X1 u0_desOut_reg_22 (.CK( clk ) , .Q( stage1_out_22 ) , .D( u0_FP_3 ) );
  DFF_X1 u0_desOut_reg_23 (.CK( clk ) , .Q( stage1_out_23 ) , .D( u0_FP_35 ) );
  DFF_X1 u0_desOut_reg_24 (.CK( clk ) , .Q( stage1_out_24 ) , .D( u0_FP_28 ) );
  DFF_X1 u0_desOut_reg_25 (.CK( clk ) , .Q( stage1_out_25 ) , .D( u0_FP_60 ) );
  DFF_X1 u0_desOut_reg_26 (.CK( clk ) , .Q( stage1_out_26 ) , .D( u0_FP_20 ) );
  DFF_X1 u0_desOut_reg_27 (.CK( clk ) , .Q( stage1_out_27 ) , .D( u0_FP_52 ) );
  DFF_X1 u0_desOut_reg_28 (.CK( clk ) , .Q( stage1_out_28 ) , .D( u0_FP_12 ) );
  DFF_X1 u0_desOut_reg_29 (.CK( clk ) , .Q( stage1_out_29 ) , .D( u0_FP_44 ) );
  DFF_X1 u0_desOut_reg_3 (.CK( clk ) , .Q( stage1_out_3 ) , .D( u0_FP_49 ) );
  DFF_X1 u0_desOut_reg_30 (.CK( clk ) , .Q( stage1_out_30 ) , .D( u0_FP_4 ) );
  DFF_X1 u0_desOut_reg_31 (.CK( clk ) , .Q( stage1_out_31 ) , .D( u0_FP_36 ) );
  DFF_X1 u0_desOut_reg_32 (.CK( clk ) , .Q( stage1_out_32 ) , .D( u0_FP_29 ) );
  DFF_X1 u0_desOut_reg_33 (.CK( clk ) , .Q( stage1_out_33 ) , .D( u0_FP_61 ) );
  DFF_X1 u0_desOut_reg_34 (.CK( clk ) , .Q( stage1_out_34 ) , .D( u0_FP_21 ) );
  DFF_X1 u0_desOut_reg_35 (.CK( clk ) , .Q( stage1_out_35 ) , .D( u0_FP_53 ) );
  DFF_X1 u0_desOut_reg_36 (.CK( clk ) , .Q( stage1_out_36 ) , .D( u0_FP_13 ) );
  DFF_X1 u0_desOut_reg_37 (.CK( clk ) , .Q( stage1_out_37 ) , .D( u0_FP_45 ) );
  DFF_X1 u0_desOut_reg_38 (.CK( clk ) , .Q( stage1_out_38 ) , .D( u0_FP_5 ) );
  DFF_X1 u0_desOut_reg_39 (.CK( clk ) , .Q( stage1_out_39 ) , .D( u0_FP_37 ) );
  DFF_X1 u0_desOut_reg_4 (.CK( clk ) , .Q( stage1_out_4 ) , .D( u0_FP_9 ) );
  DFF_X1 u0_desOut_reg_40 (.CK( clk ) , .Q( stage1_out_40 ) , .D( u0_FP_30 ) );
  DFF_X1 u0_desOut_reg_41 (.CK( clk ) , .Q( stage1_out_41 ) , .D( u0_FP_62 ) );
  DFF_X1 u0_desOut_reg_42 (.CK( clk ) , .Q( stage1_out_42 ) , .D( u0_FP_22 ) );
  DFF_X1 u0_desOut_reg_43 (.CK( clk ) , .Q( stage1_out_43 ) , .D( u0_FP_54 ) );
  DFF_X1 u0_desOut_reg_44 (.CK( clk ) , .Q( stage1_out_44 ) , .D( u0_FP_14 ) );
  DFF_X1 u0_desOut_reg_45 (.CK( clk ) , .Q( stage1_out_45 ) , .D( u0_FP_46 ) );
  DFF_X1 u0_desOut_reg_46 (.CK( clk ) , .Q( stage1_out_46 ) , .D( u0_FP_6 ) );
  DFF_X1 u0_desOut_reg_47 (.CK( clk ) , .Q( stage1_out_47 ) , .D( u0_FP_38 ) );
  DFF_X1 u0_desOut_reg_48 (.CK( clk ) , .Q( stage1_out_48 ) , .D( u0_FP_31 ) );
  DFF_X1 u0_desOut_reg_49 (.CK( clk ) , .Q( stage1_out_49 ) , .D( u0_FP_63 ) );
  DFF_X1 u0_desOut_reg_5 (.CK( clk ) , .Q( stage1_out_5 ) , .D( u0_FP_41 ) );
  DFF_X1 u0_desOut_reg_50 (.CK( clk ) , .Q( stage1_out_50 ) , .D( u0_FP_23 ) );
  DFF_X1 u0_desOut_reg_51 (.CK( clk ) , .Q( stage1_out_51 ) , .D( u0_FP_55 ) );
  DFF_X1 u0_desOut_reg_52 (.CK( clk ) , .Q( stage1_out_52 ) , .D( u0_FP_15 ) );
  DFF_X1 u0_desOut_reg_53 (.CK( clk ) , .Q( stage1_out_53 ) , .D( u0_FP_47 ) );
  DFF_X1 u0_desOut_reg_54 (.CK( clk ) , .Q( stage1_out_54 ) , .D( u0_FP_7 ) );
  DFF_X1 u0_desOut_reg_55 (.CK( clk ) , .Q( stage1_out_55 ) , .D( u0_FP_39 ) );
  DFF_X1 u0_desOut_reg_56 (.CK( clk ) , .Q( stage1_out_56 ) , .D( u0_FP_32 ) );
  DFF_X1 u0_desOut_reg_57 (.CK( clk ) , .Q( stage1_out_57 ) , .D( u0_FP_64 ) );
  DFF_X1 u0_desOut_reg_58 (.CK( clk ) , .Q( stage1_out_58 ) , .D( u0_FP_24 ) );
  DFF_X1 u0_desOut_reg_59 (.CK( clk ) , .Q( stage1_out_59 ) , .D( u0_FP_56 ) );
  DFF_X1 u0_desOut_reg_6 (.CK( clk ) , .Q( stage1_out_6 ) , .D( u0_FP_1 ) );
  DFF_X1 u0_desOut_reg_60 (.CK( clk ) , .Q( stage1_out_60 ) , .D( u0_FP_16 ) );
  DFF_X1 u0_desOut_reg_61 (.CK( clk ) , .Q( stage1_out_61 ) , .D( u0_FP_48 ) );
  DFF_X1 u0_desOut_reg_62 (.CK( clk ) , .Q( stage1_out_62 ) , .D( u0_FP_8 ) );
  DFF_X1 u0_desOut_reg_63 (.CK( clk ) , .Q( stage1_out_63 ) , .D( u0_FP_40 ) );
  DFF_X1 u0_desOut_reg_7 (.CK( clk ) , .Q( stage1_out_7 ) , .D( u0_FP_33 ) );
  DFF_X1 u0_desOut_reg_8 (.CK( clk ) , .Q( stage1_out_8 ) , .D( u0_FP_26 ) );
  DFF_X1 u0_desOut_reg_9 (.CK( clk ) , .Q( stage1_out_9 ) , .D( u0_FP_58 ) );
  DFF_X1 u0_key_r_reg_0 (.CK( clk ) , .D( key_a_0 ) , .Q( u0_key_r_0 ) );
  DFF_X1 u0_key_r_reg_1 (.CK( clk ) , .D( key_a_1 ) , .Q( u0_key_r_1 ) );
  DFF_X1 u0_key_r_reg_10 (.CK( clk ) , .D( key_a_10 ) , .Q( u0_key_r_10 ) );
  DFF_X1 u0_key_r_reg_11 (.CK( clk ) , .D( key_a_11 ) , .Q( u0_key_r_11 ) );
  DFF_X1 u0_key_r_reg_12 (.CK( clk ) , .D( key_a_12 ) , .Q( u0_key_r_12 ) );
  DFF_X1 u0_key_r_reg_13 (.CK( clk ) , .D( key_a_13 ) , .Q( u0_key_r_13 ) );
  DFF_X1 u0_key_r_reg_14 (.CK( clk ) , .D( key_a_14 ) , .Q( u0_key_r_14 ) );
  DFF_X1 u0_key_r_reg_15 (.CK( clk ) , .D( key_a_15 ) , .Q( u0_key_r_15 ) );
  DFF_X1 u0_key_r_reg_16 (.CK( clk ) , .D( key_a_16 ) , .Q( u0_key_r_16 ) );
  DFF_X1 u0_key_r_reg_17 (.CK( clk ) , .D( key_a_17 ) , .Q( u0_key_r_17 ) );
  DFF_X1 u0_key_r_reg_18 (.CK( clk ) , .D( key_a_18 ) , .Q( u0_key_r_18 ) );
  DFF_X1 u0_key_r_reg_19 (.CK( clk ) , .D( key_a_19 ) , .Q( u0_key_r_19 ) );
  DFF_X1 u0_key_r_reg_2 (.CK( clk ) , .D( key_a_2 ) , .Q( u0_key_r_2 ) );
  DFF_X1 u0_key_r_reg_20 (.CK( clk ) , .D( key_a_20 ) , .Q( u0_key_r_20 ) );
  DFF_X1 u0_key_r_reg_21 (.CK( clk ) , .D( key_a_21 ) , .Q( u0_key_r_21 ) );
  DFF_X1 u0_key_r_reg_22 (.CK( clk ) , .D( key_a_22 ) , .Q( u0_key_r_22 ) );
  DFF_X1 u0_key_r_reg_23 (.CK( clk ) , .D( key_a_23 ) , .Q( u0_key_r_23 ) );
  DFF_X1 u0_key_r_reg_24 (.CK( clk ) , .D( key_a_24 ) , .Q( u0_key_r_24 ) );
  DFF_X1 u0_key_r_reg_25 (.CK( clk ) , .D( key_a_25 ) , .Q( u0_key_r_25 ) );
  DFF_X1 u0_key_r_reg_26 (.CK( clk ) , .D( key_a_26 ) , .Q( u0_key_r_26 ) );
  DFF_X1 u0_key_r_reg_27 (.CK( clk ) , .D( key_a_27 ) , .Q( u0_key_r_27 ) );
  DFF_X1 u0_key_r_reg_28 (.CK( clk ) , .D( key_a_28 ) , .Q( u0_key_r_28 ) );
  DFF_X1 u0_key_r_reg_29 (.CK( clk ) , .D( key_a_29 ) , .Q( u0_key_r_29 ) );
  DFF_X1 u0_key_r_reg_3 (.CK( clk ) , .D( key_a_3 ) , .Q( u0_key_r_3 ) );
  DFF_X1 u0_key_r_reg_30 (.CK( clk ) , .D( key_a_30 ) , .Q( u0_key_r_30 ) );
  DFF_X1 u0_key_r_reg_31 (.CK( clk ) , .D( key_a_31 ) , .Q( u0_key_r_31 ) );
  DFF_X1 u0_key_r_reg_32 (.CK( clk ) , .D( key_a_32 ) , .Q( u0_key_r_32 ) );
  DFF_X1 u0_key_r_reg_33 (.CK( clk ) , .D( key_a_33 ) , .Q( u0_key_r_33 ) );
  DFF_X1 u0_key_r_reg_34 (.CK( clk ) , .D( key_a_34 ) , .Q( u0_key_r_34 ) );
  DFF_X1 u0_key_r_reg_35 (.CK( clk ) , .D( key_a_35 ) , .Q( u0_key_r_35 ) );
  DFF_X1 u0_key_r_reg_36 (.CK( clk ) , .D( key_a_36 ) , .Q( u0_key_r_36 ) );
  DFF_X1 u0_key_r_reg_37 (.CK( clk ) , .D( key_a_37 ) , .Q( u0_key_r_37 ) );
  DFF_X1 u0_key_r_reg_38 (.CK( clk ) , .D( key_a_38 ) , .Q( u0_key_r_38 ) );
  DFF_X1 u0_key_r_reg_39 (.CK( clk ) , .D( key_a_39 ) , .Q( u0_key_r_39 ) );
  DFF_X1 u0_key_r_reg_4 (.CK( clk ) , .D( key_a_4 ) , .Q( u0_key_r_4 ) );
  DFF_X1 u0_key_r_reg_40 (.CK( clk ) , .D( key_a_40 ) , .Q( u0_key_r_40 ) );
  DFF_X1 u0_key_r_reg_41 (.CK( clk ) , .D( key_a_41 ) , .Q( u0_key_r_41 ) );
  DFF_X1 u0_key_r_reg_42 (.CK( clk ) , .D( key_a_42 ) , .Q( u0_key_r_42 ) );
  DFF_X1 u0_key_r_reg_43 (.CK( clk ) , .D( key_a_43 ) , .Q( u0_key_r_43 ) );
  DFF_X1 u0_key_r_reg_44 (.CK( clk ) , .D( key_a_44 ) , .Q( u0_key_r_44 ) );
  DFF_X1 u0_key_r_reg_45 (.CK( clk ) , .D( key_a_45 ) , .Q( u0_key_r_45 ) );
  DFF_X1 u0_key_r_reg_46 (.CK( clk ) , .D( key_a_46 ) , .Q( u0_key_r_46 ) );
  DFF_X1 u0_key_r_reg_47 (.CK( clk ) , .D( key_a_47 ) , .Q( u0_key_r_47 ) );
  DFF_X1 u0_key_r_reg_48 (.CK( clk ) , .D( key_a_48 ) , .Q( u0_key_r_48 ) );
  DFF_X1 u0_key_r_reg_49 (.CK( clk ) , .D( key_a_49 ) , .Q( u0_key_r_49 ) );
  DFF_X1 u0_key_r_reg_5 (.CK( clk ) , .D( key_a_5 ) , .Q( u0_key_r_5 ) );
  DFF_X1 u0_key_r_reg_50 (.CK( clk ) , .D( key_a_50 ) , .Q( u0_key_r_50 ) );
  DFF_X1 u0_key_r_reg_51 (.CK( clk ) , .D( key_a_51 ) , .Q( u0_key_r_51 ) );
  DFF_X1 u0_key_r_reg_52 (.CK( clk ) , .D( key_a_52 ) , .Q( u0_key_r_52 ) );
  DFF_X1 u0_key_r_reg_53 (.CK( clk ) , .D( key_a_53 ) , .Q( u0_key_r_53 ) );
  DFF_X1 u0_key_r_reg_54 (.CK( clk ) , .D( key_a_54 ) , .Q( u0_key_r_54 ) );
  DFF_X1 u0_key_r_reg_55 (.CK( clk ) , .D( key_a_55 ) , .Q( u0_key_r_55 ) );
  DFF_X1 u0_key_r_reg_6 (.CK( clk ) , .D( key_a_6 ) , .Q( u0_key_r_6 ) );
  DFF_X1 u0_key_r_reg_7 (.CK( clk ) , .D( key_a_7 ) , .Q( u0_key_r_7 ) );
  DFF_X1 u0_key_r_reg_8 (.CK( clk ) , .D( key_a_8 ) , .Q( u0_key_r_8 ) );
  DFF_X1 u0_key_r_reg_9 (.CK( clk ) , .D( key_a_9 ) , .Q( u0_key_r_9 ) );
  XOR2_X1 u0_u0_U10 (.B( u0_K1_45 ) , .A( u0_desIn_r_41 ) , .Z( u0_u0_X_45 ) );
  XOR2_X1 u0_u0_U11 (.B( u0_K1_44 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_44 ) );
  XOR2_X1 u0_u0_U13 (.B( u0_K1_42 ) , .A( u0_desIn_r_33 ) , .Z( u0_u0_X_42 ) );
  XOR2_X1 u0_u0_U23 (.B( u0_K1_33 ) , .A( u0_desIn_r_43 ) , .Z( u0_u0_X_33 ) );
  XOR2_X1 u0_u0_U29 (.B( u0_K1_28 ) , .A( u0_desIn_r_19 ) , .Z( u0_u0_X_28 ) );
  XOR2_X1 u0_u0_U32 (.B( u0_K1_25 ) , .A( u0_desIn_r_61 ) , .Z( u0_u0_X_25 ) );
  XOR2_X1 u0_u0_U34 (.B( u0_K1_23 ) , .A( u0_desIn_r_61 ) , .Z( u0_u0_X_23 ) );
  XOR2_X1 u0_u0_U35 (.B( u0_K1_22 ) , .A( u0_desIn_r_53 ) , .Z( u0_u0_X_22 ) );
  XOR2_X1 u0_u0_U36 (.B( u0_K1_21 ) , .A( u0_desIn_r_45 ) , .Z( u0_u0_X_21 ) );
  XOR2_X1 u0_u0_U42 (.B( u0_K1_16 ) , .A( u0_desIn_r_21 ) , .Z( u0_u0_X_16 ) );
  XOR2_X1 u0_u0_U43 (.B( u0_K1_15 ) , .A( u0_desIn_r_13 ) , .Z( u0_u0_X_15 ) );
  XOR2_X1 u0_u0_U9 (.B( u0_K1_46 ) , .A( u0_desIn_r_49 ) , .Z( u0_u0_X_46 ) );
  XOR2_X1 u0_u10_U12 (.B( u0_K11_43 ) , .A( u0_R9_28 ) , .Z( u0_u10_X_43 ) );
  XOR2_X1 u0_u10_U14 (.B( u0_K11_41 ) , .A( u0_R9_28 ) , .Z( u0_u10_X_41 ) );
  XOR2_X1 u0_u10_U22 (.B( u0_K11_34 ) , .A( u0_R9_23 ) , .Z( u0_u10_X_34 ) );
  XOR2_X1 u0_u10_U35 (.B( u0_K11_22 ) , .A( u0_R9_15 ) , .Z( u0_u10_X_22 ) );
  XOR2_X1 u0_u10_U36 (.B( u0_K11_21 ) , .A( u0_R9_14 ) , .Z( u0_u10_X_21 ) );
  XOR2_X1 u0_u11_U1 (.B( u0_K12_9 ) , .A( u0_R10_6 ) , .Z( u0_u11_X_9 ) );
  XOR2_X1 u0_u11_U10 (.B( u0_K12_45 ) , .A( u0_R10_30 ) , .Z( u0_u11_X_45 ) );
  XOR2_X1 u0_u11_U15 (.B( u0_K12_40 ) , .A( u0_R10_27 ) , .Z( u0_u11_X_40 ) );
  XOR2_X1 u0_u11_U17 (.B( u0_K12_39 ) , .A( u0_R10_26 ) , .Z( u0_u11_X_39 ) );
  XOR2_X1 u0_u11_U22 (.B( u0_K12_34 ) , .A( u0_R10_23 ) , .Z( u0_u11_X_34 ) );
  XOR2_X1 u0_u11_U23 (.B( u0_K12_33 ) , .A( u0_R10_22 ) , .Z( u0_u11_X_33 ) );
  XOR2_X1 u0_u11_U35 (.B( u0_K12_22 ) , .A( u0_R10_15 ) , .Z( u0_u11_X_22 ) );
  XOR2_X1 u0_u11_U37 (.B( u0_K12_20 ) , .A( u0_R10_13 ) , .Z( u0_u11_X_20 ) );
  XOR2_X1 u0_u11_U38 (.B( u0_K12_1 ) , .A( u0_R10_32 ) , .Z( u0_u11_X_1 ) );
  XOR2_X1 u0_u11_U40 (.B( u0_K12_18 ) , .A( u0_R10_13 ) , .Z( u0_u11_X_18 ) );
  XOR2_X1 u0_u11_U42 (.B( u0_K12_16 ) , .A( u0_R10_11 ) , .Z( u0_u11_X_16 ) );
  XOR2_X1 u0_u11_U43 (.B( u0_K12_15 ) , .A( u0_R10_10 ) , .Z( u0_u11_X_15 ) );
  XOR2_X1 u0_u11_U44 (.B( u0_K12_14 ) , .A( u0_R10_9 ) , .Z( u0_u11_X_14 ) );
  XOR2_X1 u0_u11_U45 (.B( u0_K12_13 ) , .A( u0_R10_8 ) , .Z( u0_u11_X_13 ) );
  XOR2_X1 u0_u11_U46 (.B( u0_K12_12 ) , .A( u0_R10_9 ) , .Z( u0_u11_X_12 ) );
  XOR2_X1 u0_u11_U47 (.B( u0_K12_11 ) , .A( u0_R10_8 ) , .Z( u0_u11_X_11 ) );
  XOR2_X1 u0_u11_U48 (.B( u0_K12_10 ) , .A( u0_R10_7 ) , .Z( u0_u11_X_10 ) );
  XOR2_X1 u0_u11_U8 (.B( u0_K12_47 ) , .A( u0_R10_32 ) , .Z( u0_u11_X_47 ) );
  XOR2_X1 u0_u11_U9 (.B( u0_K12_46 ) , .A( u0_R10_31 ) , .Z( u0_u11_X_46 ) );
  XOR2_X1 u0_u12_U10 (.B( u0_K13_45 ) , .A( u0_R11_30 ) , .Z( u0_u12_X_45 ) );
  XOR2_X1 u0_u12_U11 (.B( u0_K13_44 ) , .A( u0_R11_29 ) , .Z( u0_u12_X_44 ) );
  XOR2_X1 u0_u12_U13 (.B( u0_K13_42 ) , .A( u0_R11_29 ) , .Z( u0_u12_X_42 ) );
  XOR2_X1 u0_u12_U15 (.B( u0_K13_40 ) , .A( u0_R11_27 ) , .Z( u0_u12_X_40 ) );
  XOR2_X1 u0_u12_U17 (.B( u0_K13_39 ) , .A( u0_R11_26 ) , .Z( u0_u12_X_39 ) );
  XOR2_X1 u0_u12_U18 (.B( u0_K13_38 ) , .A( u0_R11_25 ) , .Z( u0_u12_X_38 ) );
  XOR2_X1 u0_u12_U19 (.B( u0_K13_37 ) , .A( u0_R11_24 ) , .Z( u0_u12_X_37 ) );
  XOR2_X1 u0_u12_U20 (.B( u0_K13_36 ) , .A( u0_R11_25 ) , .Z( u0_u12_X_36 ) );
  XOR2_X1 u0_u12_U21 (.B( u0_K13_35 ) , .A( u0_R11_24 ) , .Z( u0_u12_X_35 ) );
  XOR2_X1 u0_u12_U22 (.B( u0_K13_34 ) , .A( u0_R11_23 ) , .Z( u0_u12_X_34 ) );
  XOR2_X1 u0_u12_U23 (.B( u0_K13_33 ) , .A( u0_R11_22 ) , .Z( u0_u12_X_33 ) );
  XOR2_X1 u0_u12_U24 (.B( u0_K13_32 ) , .A( u0_R11_21 ) , .Z( u0_u12_X_32 ) );
  XOR2_X1 u0_u12_U26 (.B( u0_K13_30 ) , .A( u0_R11_21 ) , .Z( u0_u12_X_30 ) );
  XOR2_X1 u0_u12_U27 (.B( u0_K13_2 ) , .A( u0_R11_1 ) , .Z( u0_u12_X_2 ) );
  XOR2_X1 u0_u12_U29 (.B( u0_K13_28 ) , .A( u0_R11_19 ) , .Z( u0_u12_X_28 ) );
  XOR2_X1 u0_u12_U3 (.B( u0_K13_7 ) , .A( u0_R11_4 ) , .Z( u0_u12_X_7 ) );
  XOR2_X1 u0_u12_U30 (.B( u0_K13_27 ) , .A( u0_R11_18 ) , .Z( u0_u12_X_27 ) );
  XOR2_X1 u0_u12_U31 (.B( u0_K13_26 ) , .A( u0_R11_17 ) , .Z( u0_u12_X_26 ) );
  XOR2_X1 u0_u12_U33 (.B( u0_K13_24 ) , .A( u0_R11_17 ) , .Z( u0_u12_X_24 ) );
  XOR2_X1 u0_u12_U44 (.B( u0_K13_14 ) , .A( u0_R11_9 ) , .Z( u0_u12_X_14 ) );
  XOR2_X1 u0_u12_U45 (.B( u0_K13_13 ) , .A( u0_R11_8 ) , .Z( u0_u12_X_13 ) );
  XOR2_X1 u0_u12_U46 (.B( u0_K13_12 ) , .A( u0_R11_9 ) , .Z( u0_u12_X_12 ) );
  XOR2_X1 u0_u12_U47 (.B( u0_K13_11 ) , .A( u0_R11_8 ) , .Z( u0_u12_X_11 ) );
  XOR2_X1 u0_u12_U48 (.B( u0_K13_10 ) , .A( u0_R11_7 ) , .Z( u0_u12_X_10 ) );
  XOR2_X1 u0_u12_U5 (.B( u0_K13_5 ) , .A( u0_R11_4 ) , .Z( u0_u12_X_5 ) );
  XOR2_X1 u0_u12_U7 (.B( u0_K13_48 ) , .A( u0_R11_1 ) , .Z( u0_u12_X_48 ) );
  XOR2_X1 u0_u12_U9 (.B( u0_K13_46 ) , .A( u0_R11_31 ) , .Z( u0_u12_X_46 ) );
  XOR2_X1 u0_u13_U1 (.B( u0_K14_9 ) , .A( u0_R12_6 ) , .Z( u0_u13_X_9 ) );
  XOR2_X1 u0_u13_U11 (.B( u0_K14_44 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_44 ) );
  XOR2_X1 u0_u13_U12 (.B( u0_K14_43 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_43 ) );
  XOR2_X1 u0_u13_U13 (.B( u0_K14_42 ) , .A( u0_R12_29 ) , .Z( u0_u13_X_42 ) );
  XOR2_X1 u0_u13_U14 (.B( u0_K14_41 ) , .A( u0_R12_28 ) , .Z( u0_u13_X_41 ) );
  XOR2_X1 u0_u13_U15 (.B( u0_K14_40 ) , .A( u0_R12_27 ) , .Z( u0_u13_X_40 ) );
  XOR2_X1 u0_u13_U16 (.B( u0_K14_3 ) , .A( u0_R12_2 ) , .Z( u0_u13_X_3 ) );
  XOR2_X1 u0_u13_U17 (.B( u0_K14_39 ) , .A( u0_R12_26 ) , .Z( u0_u13_X_39 ) );
  XOR2_X1 u0_u13_U18 (.B( u0_K14_38 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_38 ) );
  XOR2_X1 u0_u13_U2 (.B( u0_K14_8 ) , .A( u0_R12_5 ) , .Z( u0_u13_X_8 ) );
  XOR2_X1 u0_u13_U20 (.B( u0_K14_36 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_36 ) );
  XOR2_X1 u0_u13_U24 (.B( u0_K14_32 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_32 ) );
  XOR2_X1 u0_u13_U26 (.B( u0_K14_30 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_30 ) );
  XOR2_X1 u0_u13_U27 (.B( u0_K14_2 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_2 ) );
  XOR2_X1 u0_u13_U30 (.B( u0_K14_27 ) , .A( u0_R12_18 ) , .Z( u0_u13_X_27 ) );
  XOR2_X1 u0_u13_U35 (.B( u0_K14_22 ) , .A( u0_R12_15 ) , .Z( u0_u13_X_22 ) );
  XOR2_X1 u0_u13_U36 (.B( u0_K14_21 ) , .A( u0_R12_14 ) , .Z( u0_u13_X_21 ) );
  XOR2_X1 u0_u13_U37 (.B( u0_K14_20 ) , .A( u0_R12_13 ) , .Z( u0_u13_X_20 ) );
  XOR2_X1 u0_u13_U38 (.B( u0_K14_1 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_1 ) );
  XOR2_X1 u0_u13_U39 (.B( u0_K14_19 ) , .A( u0_R12_12 ) , .Z( u0_u13_X_19 ) );
  XOR2_X1 u0_u13_U4 (.B( u0_K14_6 ) , .A( u0_R12_5 ) , .Z( u0_u13_X_6 ) );
  XOR2_X1 u0_u13_U40 (.B( u0_K14_18 ) , .A( u0_R12_13 ) , .Z( u0_u13_X_18 ) );
  XOR2_X1 u0_u13_U41 (.B( u0_K14_17 ) , .A( u0_R12_12 ) , .Z( u0_u13_X_17 ) );
  XOR2_X1 u0_u13_U42 (.B( u0_K14_16 ) , .A( u0_R12_11 ) , .Z( u0_u13_X_16 ) );
  XOR2_X1 u0_u13_U43 (.B( u0_K14_15 ) , .A( u0_R12_10 ) , .Z( u0_u13_X_15 ) );
  XOR2_X1 u0_u13_U44 (.B( u0_K14_14 ) , .A( u0_R12_9 ) , .Z( u0_u13_X_14 ) );
  XOR2_X1 u0_u13_U45 (.B( u0_K14_13 ) , .A( u0_R12_8 ) , .Z( u0_u13_X_13 ) );
  XOR2_X1 u0_u13_U46 (.B( u0_K14_12 ) , .A( u0_R12_9 ) , .Z( u0_u13_X_12 ) );
  XOR2_X1 u0_u13_U47 (.B( u0_K14_11 ) , .A( u0_R12_8 ) , .Z( u0_u13_X_11 ) );
  XOR2_X1 u0_u13_U48 (.B( u0_K14_10 ) , .A( u0_R12_7 ) , .Z( u0_u13_X_10 ) );
  XOR2_X1 u0_u13_U6 (.B( u0_K14_4 ) , .A( u0_R12_3 ) , .Z( u0_u13_X_4 ) );
  XOR2_X1 u0_u13_U7 (.B( u0_K14_48 ) , .A( u0_R12_1 ) , .Z( u0_u13_X_48 ) );
  XOR2_X1 u0_u13_U8 (.B( u0_K14_47 ) , .A( u0_R12_32 ) , .Z( u0_u13_X_47 ) );
  XOR2_X1 u0_u13_U9 (.B( u0_K14_46 ) , .A( u0_R12_31 ) , .Z( u0_u13_X_46 ) );
  OAI22_X1 u0_u13_u2_U10 (.B1( u0_u13_u2_n151 ) , .A2( u0_u13_u2_n152 ) , .A1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n160 ) , .B2( u0_u13_u2_n168 ) );
  NAND3_X1 u0_u13_u2_U100 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n98 ) );
  NOR3_X1 u0_u13_u2_U11 (.A1( u0_u13_u2_n150 ) , .ZN( u0_u13_u2_n151 ) , .A3( u0_u13_u2_n175 ) , .A2( u0_u13_u2_n188 ) );
  AOI21_X1 u0_u13_u2_U12 (.B2( u0_u13_u2_n123 ) , .ZN( u0_u13_u2_n125 ) , .A( u0_u13_u2_n171 ) , .B1( u0_u13_u2_n184 ) );
  INV_X1 u0_u13_u2_U13 (.A( u0_u13_u2_n150 ) , .ZN( u0_u13_u2_n184 ) );
  AOI21_X1 u0_u13_u2_U14 (.ZN( u0_u13_u2_n144 ) , .B2( u0_u13_u2_n155 ) , .A( u0_u13_u2_n172 ) , .B1( u0_u13_u2_n185 ) );
  AOI21_X1 u0_u13_u2_U15 (.B2( u0_u13_u2_n143 ) , .ZN( u0_u13_u2_n145 ) , .B1( u0_u13_u2_n152 ) , .A( u0_u13_u2_n171 ) );
  INV_X1 u0_u13_u2_U16 (.A( u0_u13_u2_n156 ) , .ZN( u0_u13_u2_n171 ) );
  INV_X1 u0_u13_u2_U17 (.A( u0_u13_u2_n120 ) , .ZN( u0_u13_u2_n188 ) );
  NAND2_X1 u0_u13_u2_U18 (.A2( u0_u13_u2_n122 ) , .ZN( u0_u13_u2_n150 ) , .A1( u0_u13_u2_n152 ) );
  INV_X1 u0_u13_u2_U19 (.A( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n170 ) );
  INV_X1 u0_u13_u2_U20 (.A( u0_u13_u2_n137 ) , .ZN( u0_u13_u2_n173 ) );
  NAND2_X1 u0_u13_u2_U21 (.A1( u0_u13_u2_n132 ) , .A2( u0_u13_u2_n139 ) , .ZN( u0_u13_u2_n157 ) );
  INV_X1 u0_u13_u2_U22 (.A( u0_u13_u2_n113 ) , .ZN( u0_u13_u2_n178 ) );
  INV_X1 u0_u13_u2_U23 (.A( u0_u13_u2_n139 ) , .ZN( u0_u13_u2_n175 ) );
  INV_X1 u0_u13_u2_U24 (.A( u0_u13_u2_n155 ) , .ZN( u0_u13_u2_n181 ) );
  INV_X1 u0_u13_u2_U25 (.A( u0_u13_u2_n119 ) , .ZN( u0_u13_u2_n177 ) );
  INV_X1 u0_u13_u2_U26 (.A( u0_u13_u2_n116 ) , .ZN( u0_u13_u2_n180 ) );
  INV_X1 u0_u13_u2_U27 (.A( u0_u13_u2_n131 ) , .ZN( u0_u13_u2_n179 ) );
  INV_X1 u0_u13_u2_U28 (.A( u0_u13_u2_n154 ) , .ZN( u0_u13_u2_n176 ) );
  NAND2_X1 u0_u13_u2_U29 (.A2( u0_u13_u2_n116 ) , .A1( u0_u13_u2_n117 ) , .ZN( u0_u13_u2_n118 ) );
  NOR2_X1 u0_u13_u2_U3 (.ZN( u0_u13_u2_n121 ) , .A2( u0_u13_u2_n177 ) , .A1( u0_u13_u2_n180 ) );
  INV_X1 u0_u13_u2_U30 (.A( u0_u13_u2_n132 ) , .ZN( u0_u13_u2_n182 ) );
  INV_X1 u0_u13_u2_U31 (.A( u0_u13_u2_n158 ) , .ZN( u0_u13_u2_n183 ) );
  OAI21_X1 u0_u13_u2_U32 (.A( u0_u13_u2_n156 ) , .B1( u0_u13_u2_n157 ) , .ZN( u0_u13_u2_n158 ) , .B2( u0_u13_u2_n179 ) );
  NOR2_X1 u0_u13_u2_U33 (.ZN( u0_u13_u2_n156 ) , .A1( u0_u13_u2_n166 ) , .A2( u0_u13_u2_n169 ) );
  NOR2_X1 u0_u13_u2_U34 (.A2( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n137 ) , .A1( u0_u13_u2_n140 ) );
  NOR2_X1 u0_u13_u2_U35 (.A2( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n153 ) , .A1( u0_u13_u2_n156 ) );
  AOI211_X1 u0_u13_u2_U36 (.ZN( u0_u13_u2_n130 ) , .C1( u0_u13_u2_n138 ) , .C2( u0_u13_u2_n179 ) , .B( u0_u13_u2_n96 ) , .A( u0_u13_u2_n97 ) );
  OAI22_X1 u0_u13_u2_U37 (.B1( u0_u13_u2_n133 ) , .A2( u0_u13_u2_n137 ) , .A1( u0_u13_u2_n152 ) , .B2( u0_u13_u2_n168 ) , .ZN( u0_u13_u2_n97 ) );
  OAI221_X1 u0_u13_u2_U38 (.B1( u0_u13_u2_n113 ) , .C1( u0_u13_u2_n132 ) , .A( u0_u13_u2_n149 ) , .B2( u0_u13_u2_n171 ) , .C2( u0_u13_u2_n172 ) , .ZN( u0_u13_u2_n96 ) );
  OAI221_X1 u0_u13_u2_U39 (.A( u0_u13_u2_n115 ) , .C2( u0_u13_u2_n123 ) , .B2( u0_u13_u2_n143 ) , .B1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n163 ) , .C1( u0_u13_u2_n168 ) );
  INV_X1 u0_u13_u2_U4 (.A( u0_u13_u2_n134 ) , .ZN( u0_u13_u2_n185 ) );
  OAI21_X1 u0_u13_u2_U40 (.A( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n115 ) , .B1( u0_u13_u2_n176 ) , .B2( u0_u13_u2_n178 ) );
  OAI221_X1 u0_u13_u2_U41 (.A( u0_u13_u2_n135 ) , .B2( u0_u13_u2_n136 ) , .B1( u0_u13_u2_n137 ) , .ZN( u0_u13_u2_n162 ) , .C2( u0_u13_u2_n167 ) , .C1( u0_u13_u2_n185 ) );
  AND3_X1 u0_u13_u2_U42 (.A3( u0_u13_u2_n131 ) , .A2( u0_u13_u2_n132 ) , .A1( u0_u13_u2_n133 ) , .ZN( u0_u13_u2_n136 ) );
  AOI22_X1 u0_u13_u2_U43 (.ZN( u0_u13_u2_n135 ) , .B1( u0_u13_u2_n140 ) , .A1( u0_u13_u2_n156 ) , .B2( u0_u13_u2_n180 ) , .A2( u0_u13_u2_n188 ) );
  AOI21_X1 u0_u13_u2_U44 (.ZN( u0_u13_u2_n149 ) , .B1( u0_u13_u2_n173 ) , .B2( u0_u13_u2_n188 ) , .A( u0_u13_u2_n95 ) );
  AND3_X1 u0_u13_u2_U45 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n156 ) , .ZN( u0_u13_u2_n95 ) );
  OAI21_X1 u0_u13_u2_U46 (.A( u0_u13_u2_n141 ) , .B2( u0_u13_u2_n142 ) , .ZN( u0_u13_u2_n146 ) , .B1( u0_u13_u2_n153 ) );
  OAI21_X1 u0_u13_u2_U47 (.A( u0_u13_u2_n140 ) , .ZN( u0_u13_u2_n141 ) , .B1( u0_u13_u2_n176 ) , .B2( u0_u13_u2_n177 ) );
  NOR3_X1 u0_u13_u2_U48 (.ZN( u0_u13_u2_n142 ) , .A3( u0_u13_u2_n175 ) , .A2( u0_u13_u2_n178 ) , .A1( u0_u13_u2_n181 ) );
  OAI21_X1 u0_u13_u2_U49 (.A( u0_u13_u2_n101 ) , .B2( u0_u13_u2_n121 ) , .B1( u0_u13_u2_n153 ) , .ZN( u0_u13_u2_n164 ) );
  NOR4_X1 u0_u13_u2_U5 (.A4( u0_u13_u2_n124 ) , .A3( u0_u13_u2_n125 ) , .A2( u0_u13_u2_n126 ) , .A1( u0_u13_u2_n127 ) , .ZN( u0_u13_u2_n128 ) );
  NAND2_X1 u0_u13_u2_U50 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n155 ) );
  NAND2_X1 u0_u13_u2_U51 (.A2( u0_u13_u2_n105 ) , .A1( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n143 ) );
  NAND2_X1 u0_u13_u2_U52 (.A1( u0_u13_u2_n104 ) , .A2( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n152 ) );
  NAND2_X1 u0_u13_u2_U53 (.A1( u0_u13_u2_n100 ) , .A2( u0_u13_u2_n105 ) , .ZN( u0_u13_u2_n132 ) );
  INV_X1 u0_u13_u2_U54 (.A( u0_u13_u2_n140 ) , .ZN( u0_u13_u2_n168 ) );
  INV_X1 u0_u13_u2_U55 (.A( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n167 ) );
  NAND2_X1 u0_u13_u2_U56 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n113 ) );
  NAND2_X1 u0_u13_u2_U57 (.A1( u0_u13_u2_n106 ) , .A2( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n131 ) );
  NAND2_X1 u0_u13_u2_U58 (.A1( u0_u13_u2_n103 ) , .A2( u0_u13_u2_n107 ) , .ZN( u0_u13_u2_n139 ) );
  NAND2_X1 u0_u13_u2_U59 (.A1( u0_u13_u2_n103 ) , .A2( u0_u13_u2_n105 ) , .ZN( u0_u13_u2_n133 ) );
  AOI21_X1 u0_u13_u2_U6 (.B2( u0_u13_u2_n119 ) , .ZN( u0_u13_u2_n127 ) , .A( u0_u13_u2_n137 ) , .B1( u0_u13_u2_n155 ) );
  NAND2_X1 u0_u13_u2_U60 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n103 ) , .ZN( u0_u13_u2_n154 ) );
  NAND2_X1 u0_u13_u2_U61 (.A2( u0_u13_u2_n103 ) , .A1( u0_u13_u2_n104 ) , .ZN( u0_u13_u2_n119 ) );
  NAND2_X1 u0_u13_u2_U62 (.A2( u0_u13_u2_n107 ) , .A1( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n123 ) );
  NAND2_X1 u0_u13_u2_U63 (.A1( u0_u13_u2_n104 ) , .A2( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n122 ) );
  INV_X1 u0_u13_u2_U64 (.A( u0_u13_u2_n114 ) , .ZN( u0_u13_u2_n172 ) );
  NAND2_X1 u0_u13_u2_U65 (.A2( u0_u13_u2_n100 ) , .A1( u0_u13_u2_n102 ) , .ZN( u0_u13_u2_n116 ) );
  NAND2_X1 u0_u13_u2_U66 (.A1( u0_u13_u2_n102 ) , .A2( u0_u13_u2_n108 ) , .ZN( u0_u13_u2_n120 ) );
  NAND2_X1 u0_u13_u2_U67 (.A2( u0_u13_u2_n105 ) , .A1( u0_u13_u2_n106 ) , .ZN( u0_u13_u2_n117 ) );
  INV_X1 u0_u13_u2_U68 (.ZN( u0_u13_u2_n187 ) , .A( u0_u13_u2_n99 ) );
  OAI21_X1 u0_u13_u2_U69 (.B1( u0_u13_u2_n137 ) , .B2( u0_u13_u2_n143 ) , .A( u0_u13_u2_n98 ) , .ZN( u0_u13_u2_n99 ) );
  AOI21_X1 u0_u13_u2_U7 (.ZN( u0_u13_u2_n124 ) , .B1( u0_u13_u2_n131 ) , .B2( u0_u13_u2_n143 ) , .A( u0_u13_u2_n172 ) );
  NOR2_X1 u0_u13_u2_U70 (.A2( u0_u13_X_16 ) , .ZN( u0_u13_u2_n140 ) , .A1( u0_u13_u2_n166 ) );
  NOR2_X1 u0_u13_u2_U71 (.A2( u0_u13_X_13 ) , .A1( u0_u13_X_14 ) , .ZN( u0_u13_u2_n100 ) );
  NOR2_X1 u0_u13_u2_U72 (.A2( u0_u13_X_16 ) , .A1( u0_u13_X_17 ) , .ZN( u0_u13_u2_n138 ) );
  NOR2_X1 u0_u13_u2_U73 (.A2( u0_u13_X_15 ) , .A1( u0_u13_X_18 ) , .ZN( u0_u13_u2_n104 ) );
  NOR2_X1 u0_u13_u2_U74 (.A2( u0_u13_X_14 ) , .ZN( u0_u13_u2_n103 ) , .A1( u0_u13_u2_n174 ) );
  NOR2_X1 u0_u13_u2_U75 (.A2( u0_u13_X_15 ) , .ZN( u0_u13_u2_n102 ) , .A1( u0_u13_u2_n165 ) );
  NOR2_X1 u0_u13_u2_U76 (.A2( u0_u13_X_17 ) , .ZN( u0_u13_u2_n114 ) , .A1( u0_u13_u2_n169 ) );
  AND2_X1 u0_u13_u2_U77 (.A1( u0_u13_X_15 ) , .ZN( u0_u13_u2_n105 ) , .A2( u0_u13_u2_n165 ) );
  AND2_X1 u0_u13_u2_U78 (.A2( u0_u13_X_15 ) , .A1( u0_u13_X_18 ) , .ZN( u0_u13_u2_n107 ) );
  AND2_X1 u0_u13_u2_U79 (.A1( u0_u13_X_14 ) , .ZN( u0_u13_u2_n106 ) , .A2( u0_u13_u2_n174 ) );
  AOI21_X1 u0_u13_u2_U8 (.B2( u0_u13_u2_n120 ) , .B1( u0_u13_u2_n121 ) , .ZN( u0_u13_u2_n126 ) , .A( u0_u13_u2_n167 ) );
  AND2_X1 u0_u13_u2_U80 (.A1( u0_u13_X_13 ) , .A2( u0_u13_X_14 ) , .ZN( u0_u13_u2_n108 ) );
  INV_X1 u0_u13_u2_U81 (.A( u0_u13_X_16 ) , .ZN( u0_u13_u2_n169 ) );
  INV_X1 u0_u13_u2_U82 (.A( u0_u13_X_17 ) , .ZN( u0_u13_u2_n166 ) );
  INV_X1 u0_u13_u2_U83 (.A( u0_u13_X_13 ) , .ZN( u0_u13_u2_n174 ) );
  INV_X1 u0_u13_u2_U84 (.A( u0_u13_X_18 ) , .ZN( u0_u13_u2_n165 ) );
  NAND4_X1 u0_u13_u2_U85 (.ZN( u0_out13_30 ) , .A4( u0_u13_u2_n147 ) , .A3( u0_u13_u2_n148 ) , .A2( u0_u13_u2_n149 ) , .A1( u0_u13_u2_n187 ) );
  NOR3_X1 u0_u13_u2_U86 (.A3( u0_u13_u2_n144 ) , .A2( u0_u13_u2_n145 ) , .A1( u0_u13_u2_n146 ) , .ZN( u0_u13_u2_n147 ) );
  AOI21_X1 u0_u13_u2_U87 (.B2( u0_u13_u2_n138 ) , .ZN( u0_u13_u2_n148 ) , .A( u0_u13_u2_n162 ) , .B1( u0_u13_u2_n182 ) );
  NAND4_X1 u0_u13_u2_U88 (.ZN( u0_out13_24 ) , .A4( u0_u13_u2_n111 ) , .A3( u0_u13_u2_n112 ) , .A1( u0_u13_u2_n130 ) , .A2( u0_u13_u2_n187 ) );
  AOI221_X1 u0_u13_u2_U89 (.A( u0_u13_u2_n109 ) , .B1( u0_u13_u2_n110 ) , .ZN( u0_u13_u2_n111 ) , .C1( u0_u13_u2_n134 ) , .C2( u0_u13_u2_n170 ) , .B2( u0_u13_u2_n173 ) );
  OAI22_X1 u0_u13_u2_U9 (.ZN( u0_u13_u2_n109 ) , .A2( u0_u13_u2_n113 ) , .B2( u0_u13_u2_n133 ) , .B1( u0_u13_u2_n167 ) , .A1( u0_u13_u2_n168 ) );
  AOI21_X1 u0_u13_u2_U90 (.ZN( u0_u13_u2_n112 ) , .B2( u0_u13_u2_n156 ) , .A( u0_u13_u2_n164 ) , .B1( u0_u13_u2_n181 ) );
  NAND4_X1 u0_u13_u2_U91 (.ZN( u0_out13_16 ) , .A4( u0_u13_u2_n128 ) , .A3( u0_u13_u2_n129 ) , .A1( u0_u13_u2_n130 ) , .A2( u0_u13_u2_n186 ) );
  AOI22_X1 u0_u13_u2_U92 (.A2( u0_u13_u2_n118 ) , .ZN( u0_u13_u2_n129 ) , .A1( u0_u13_u2_n140 ) , .B1( u0_u13_u2_n157 ) , .B2( u0_u13_u2_n170 ) );
  INV_X1 u0_u13_u2_U93 (.A( u0_u13_u2_n163 ) , .ZN( u0_u13_u2_n186 ) );
  OR4_X1 u0_u13_u2_U94 (.ZN( u0_out13_6 ) , .A4( u0_u13_u2_n161 ) , .A3( u0_u13_u2_n162 ) , .A2( u0_u13_u2_n163 ) , .A1( u0_u13_u2_n164 ) );
  OR3_X1 u0_u13_u2_U95 (.A2( u0_u13_u2_n159 ) , .A1( u0_u13_u2_n160 ) , .ZN( u0_u13_u2_n161 ) , .A3( u0_u13_u2_n183 ) );
  AOI21_X1 u0_u13_u2_U96 (.B2( u0_u13_u2_n154 ) , .B1( u0_u13_u2_n155 ) , .ZN( u0_u13_u2_n159 ) , .A( u0_u13_u2_n167 ) );
  NAND3_X1 u0_u13_u2_U97 (.A2( u0_u13_u2_n117 ) , .A1( u0_u13_u2_n122 ) , .A3( u0_u13_u2_n123 ) , .ZN( u0_u13_u2_n134 ) );
  NAND3_X1 u0_u13_u2_U98 (.ZN( u0_u13_u2_n110 ) , .A2( u0_u13_u2_n131 ) , .A3( u0_u13_u2_n139 ) , .A1( u0_u13_u2_n154 ) );
  NAND3_X1 u0_u13_u2_U99 (.A2( u0_u13_u2_n100 ) , .ZN( u0_u13_u2_n101 ) , .A1( u0_u13_u2_n104 ) , .A3( u0_u13_u2_n114 ) );
  XOR2_X1 u0_u14_U1 (.B( u0_K15_9 ) , .A( u0_R13_6 ) , .Z( u0_u14_X_9 ) );
  XOR2_X1 u0_u14_U16 (.B( u0_K15_3 ) , .A( u0_R13_2 ) , .Z( u0_u14_X_3 ) );
  XOR2_X1 u0_u14_U2 (.B( u0_K15_8 ) , .A( u0_R13_5 ) , .Z( u0_u14_X_8 ) );
  XOR2_X1 u0_u14_U27 (.B( u0_K15_2 ) , .A( u0_R13_1 ) , .Z( u0_u14_X_2 ) );
  XOR2_X1 u0_u14_U3 (.B( u0_K15_7 ) , .A( u0_R13_4 ) , .Z( u0_u14_X_7 ) );
  XOR2_X1 u0_u14_U32 (.B( u0_K15_25 ) , .A( u0_R13_16 ) , .Z( u0_u14_X_25 ) );
  XOR2_X1 u0_u14_U33 (.B( u0_K15_24 ) , .A( u0_R13_17 ) , .Z( u0_u14_X_24 ) );
  XOR2_X1 u0_u14_U34 (.B( u0_K15_23 ) , .A( u0_R13_16 ) , .Z( u0_u14_X_23 ) );
  XOR2_X1 u0_u14_U35 (.B( u0_K15_22 ) , .A( u0_R13_15 ) , .Z( u0_u14_X_22 ) );
  XOR2_X1 u0_u14_U36 (.B( u0_K15_21 ) , .A( u0_R13_14 ) , .Z( u0_u14_X_21 ) );
  XOR2_X1 u0_u14_U37 (.B( u0_K15_20 ) , .A( u0_R13_13 ) , .Z( u0_u14_X_20 ) );
  XOR2_X1 u0_u14_U38 (.B( u0_K15_1 ) , .A( u0_R13_32 ) , .Z( u0_u14_X_1 ) );
  XOR2_X1 u0_u14_U39 (.B( u0_K15_19 ) , .A( u0_R13_12 ) , .Z( u0_u14_X_19 ) );
  XOR2_X1 u0_u14_U4 (.B( u0_K15_6 ) , .A( u0_R13_5 ) , .Z( u0_u14_X_6 ) );
  XOR2_X1 u0_u14_U40 (.B( u0_K15_18 ) , .A( u0_R13_13 ) , .Z( u0_u14_X_18 ) );
  XOR2_X1 u0_u14_U41 (.B( u0_K15_17 ) , .A( u0_R13_12 ) , .Z( u0_u14_X_17 ) );
  XOR2_X1 u0_u14_U42 (.B( u0_K15_16 ) , .A( u0_R13_11 ) , .Z( u0_u14_X_16 ) );
  XOR2_X1 u0_u14_U43 (.B( u0_K15_15 ) , .A( u0_R13_10 ) , .Z( u0_u14_X_15 ) );
  XOR2_X1 u0_u14_U44 (.B( u0_K15_14 ) , .A( u0_R13_9 ) , .Z( u0_u14_X_14 ) );
  XOR2_X1 u0_u14_U46 (.B( u0_K15_12 ) , .A( u0_R13_9 ) , .Z( u0_u14_X_12 ) );
  XOR2_X1 u0_u14_U48 (.B( u0_K15_10 ) , .A( u0_R13_7 ) , .Z( u0_u14_X_10 ) );
  XOR2_X1 u0_u14_U5 (.B( u0_K15_5 ) , .A( u0_R13_4 ) , .Z( u0_u14_X_5 ) );
  XOR2_X1 u0_u14_U6 (.B( u0_K15_4 ) , .A( u0_R13_3 ) , .Z( u0_u14_X_4 ) );
  XOR2_X1 u0_u14_U7 (.B( u0_K15_48 ) , .A( u0_R13_1 ) , .Z( u0_u14_X_48 ) );
  XOR2_X1 u0_u14_U8 (.B( u0_K15_47 ) , .A( u0_R13_32 ) , .Z( u0_u14_X_47 ) );
  AND3_X1 u0_u14_u0_U10 (.A2( u0_u14_u0_n112 ) , .ZN( u0_u14_u0_n127 ) , .A3( u0_u14_u0_n130 ) , .A1( u0_u14_u0_n148 ) );
  NAND2_X1 u0_u14_u0_U11 (.ZN( u0_u14_u0_n113 ) , .A1( u0_u14_u0_n139 ) , .A2( u0_u14_u0_n149 ) );
  AND2_X1 u0_u14_u0_U12 (.ZN( u0_u14_u0_n107 ) , .A1( u0_u14_u0_n130 ) , .A2( u0_u14_u0_n140 ) );
  AND2_X1 u0_u14_u0_U13 (.A2( u0_u14_u0_n129 ) , .A1( u0_u14_u0_n130 ) , .ZN( u0_u14_u0_n151 ) );
  AND2_X1 u0_u14_u0_U14 (.A1( u0_u14_u0_n108 ) , .A2( u0_u14_u0_n125 ) , .ZN( u0_u14_u0_n145 ) );
  INV_X1 u0_u14_u0_U15 (.A( u0_u14_u0_n143 ) , .ZN( u0_u14_u0_n173 ) );
  NOR2_X1 u0_u14_u0_U16 (.A2( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n147 ) , .A1( u0_u14_u0_n160 ) );
  NOR2_X1 u0_u14_u0_U17 (.A1( u0_u14_u0_n163 ) , .A2( u0_u14_u0_n164 ) , .ZN( u0_u14_u0_n95 ) );
  AOI21_X1 u0_u14_u0_U18 (.B1( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n132 ) , .A( u0_u14_u0_n165 ) , .B2( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U19 (.A( u0_u14_u0_n142 ) , .ZN( u0_u14_u0_n165 ) );
  OAI221_X1 u0_u14_u0_U20 (.C1( u0_u14_u0_n121 ) , .ZN( u0_u14_u0_n122 ) , .B2( u0_u14_u0_n127 ) , .A( u0_u14_u0_n143 ) , .B1( u0_u14_u0_n144 ) , .C2( u0_u14_u0_n147 ) );
  OAI22_X1 u0_u14_u0_U21 (.B1( u0_u14_u0_n125 ) , .ZN( u0_u14_u0_n126 ) , .A1( u0_u14_u0_n138 ) , .A2( u0_u14_u0_n146 ) , .B2( u0_u14_u0_n147 ) );
  OAI22_X1 u0_u14_u0_U22 (.B1( u0_u14_u0_n131 ) , .A1( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n147 ) , .A2( u0_u14_u0_n90 ) , .ZN( u0_u14_u0_n91 ) );
  AND3_X1 u0_u14_u0_U23 (.A3( u0_u14_u0_n121 ) , .A2( u0_u14_u0_n125 ) , .A1( u0_u14_u0_n148 ) , .ZN( u0_u14_u0_n90 ) );
  NAND2_X1 u0_u14_u0_U24 (.A1( u0_u14_u0_n100 ) , .A2( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n125 ) );
  INV_X1 u0_u14_u0_U25 (.A( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n161 ) );
  NOR2_X1 u0_u14_u0_U26 (.A1( u0_u14_u0_n120 ) , .ZN( u0_u14_u0_n143 ) , .A2( u0_u14_u0_n167 ) );
  OAI221_X1 u0_u14_u0_U27 (.C1( u0_u14_u0_n112 ) , .ZN( u0_u14_u0_n120 ) , .B1( u0_u14_u0_n138 ) , .B2( u0_u14_u0_n141 ) , .C2( u0_u14_u0_n147 ) , .A( u0_u14_u0_n172 ) );
  AOI211_X1 u0_u14_u0_U28 (.B( u0_u14_u0_n115 ) , .A( u0_u14_u0_n116 ) , .C2( u0_u14_u0_n117 ) , .C1( u0_u14_u0_n118 ) , .ZN( u0_u14_u0_n119 ) );
  AOI22_X1 u0_u14_u0_U29 (.B2( u0_u14_u0_n109 ) , .A2( u0_u14_u0_n110 ) , .ZN( u0_u14_u0_n111 ) , .B1( u0_u14_u0_n118 ) , .A1( u0_u14_u0_n160 ) );
  INV_X1 u0_u14_u0_U3 (.A( u0_u14_u0_n113 ) , .ZN( u0_u14_u0_n166 ) );
  NAND2_X1 u0_u14_u0_U30 (.A1( u0_u14_u0_n100 ) , .ZN( u0_u14_u0_n129 ) , .A2( u0_u14_u0_n95 ) );
  INV_X1 u0_u14_u0_U31 (.A( u0_u14_u0_n118 ) , .ZN( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U32 (.ZN( u0_u14_u0_n104 ) , .B1( u0_u14_u0_n107 ) , .B2( u0_u14_u0_n141 ) , .A( u0_u14_u0_n144 ) );
  AOI21_X1 u0_u14_u0_U33 (.B1( u0_u14_u0_n127 ) , .B2( u0_u14_u0_n129 ) , .A( u0_u14_u0_n138 ) , .ZN( u0_u14_u0_n96 ) );
  AOI21_X1 u0_u14_u0_U34 (.ZN( u0_u14_u0_n116 ) , .B2( u0_u14_u0_n142 ) , .A( u0_u14_u0_n144 ) , .B1( u0_u14_u0_n166 ) );
  NAND2_X1 u0_u14_u0_U35 (.A2( u0_u14_u0_n100 ) , .A1( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n139 ) );
  NAND2_X1 u0_u14_u0_U36 (.A2( u0_u14_u0_n100 ) , .ZN( u0_u14_u0_n131 ) , .A1( u0_u14_u0_n92 ) );
  NAND2_X1 u0_u14_u0_U37 (.A1( u0_u14_u0_n101 ) , .A2( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n150 ) );
  INV_X1 u0_u14_u0_U38 (.A( u0_u14_u0_n138 ) , .ZN( u0_u14_u0_n160 ) );
  NAND2_X1 u0_u14_u0_U39 (.A1( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n128 ) , .A2( u0_u14_u0_n95 ) );
  AOI21_X1 u0_u14_u0_U4 (.B1( u0_u14_u0_n114 ) , .ZN( u0_u14_u0_n115 ) , .B2( u0_u14_u0_n129 ) , .A( u0_u14_u0_n161 ) );
  NAND2_X1 u0_u14_u0_U40 (.ZN( u0_u14_u0_n148 ) , .A1( u0_u14_u0_n93 ) , .A2( u0_u14_u0_n95 ) );
  NAND2_X1 u0_u14_u0_U41 (.A2( u0_u14_u0_n102 ) , .A1( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n149 ) );
  NAND2_X1 u0_u14_u0_U42 (.A2( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n114 ) , .A1( u0_u14_u0_n92 ) );
  NAND2_X1 u0_u14_u0_U43 (.A2( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n121 ) , .A1( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U44 (.ZN( u0_u14_u0_n172 ) , .A( u0_u14_u0_n88 ) );
  OAI222_X1 u0_u14_u0_U45 (.C1( u0_u14_u0_n108 ) , .A1( u0_u14_u0_n125 ) , .B2( u0_u14_u0_n128 ) , .B1( u0_u14_u0_n144 ) , .A2( u0_u14_u0_n158 ) , .C2( u0_u14_u0_n161 ) , .ZN( u0_u14_u0_n88 ) );
  NAND2_X1 u0_u14_u0_U46 (.ZN( u0_u14_u0_n112 ) , .A2( u0_u14_u0_n92 ) , .A1( u0_u14_u0_n93 ) );
  OR3_X1 u0_u14_u0_U47 (.A3( u0_u14_u0_n152 ) , .A2( u0_u14_u0_n153 ) , .A1( u0_u14_u0_n154 ) , .ZN( u0_u14_u0_n155 ) );
  AOI21_X1 u0_u14_u0_U48 (.B2( u0_u14_u0_n150 ) , .B1( u0_u14_u0_n151 ) , .ZN( u0_u14_u0_n152 ) , .A( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U49 (.A( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n145 ) , .B1( u0_u14_u0_n146 ) , .ZN( u0_u14_u0_n154 ) );
  AOI21_X1 u0_u14_u0_U5 (.B2( u0_u14_u0_n131 ) , .ZN( u0_u14_u0_n134 ) , .B1( u0_u14_u0_n151 ) , .A( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U50 (.A( u0_u14_u0_n147 ) , .B2( u0_u14_u0_n148 ) , .B1( u0_u14_u0_n149 ) , .ZN( u0_u14_u0_n153 ) );
  INV_X1 u0_u14_u0_U51 (.ZN( u0_u14_u0_n171 ) , .A( u0_u14_u0_n99 ) );
  OAI211_X1 u0_u14_u0_U52 (.C2( u0_u14_u0_n140 ) , .C1( u0_u14_u0_n161 ) , .A( u0_u14_u0_n169 ) , .B( u0_u14_u0_n98 ) , .ZN( u0_u14_u0_n99 ) );
  AOI211_X1 u0_u14_u0_U53 (.C1( u0_u14_u0_n118 ) , .A( u0_u14_u0_n123 ) , .B( u0_u14_u0_n96 ) , .C2( u0_u14_u0_n97 ) , .ZN( u0_u14_u0_n98 ) );
  INV_X1 u0_u14_u0_U54 (.ZN( u0_u14_u0_n169 ) , .A( u0_u14_u0_n91 ) );
  NOR2_X1 u0_u14_u0_U55 (.A2( u0_u14_X_4 ) , .A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n118 ) );
  NOR2_X1 u0_u14_u0_U56 (.A2( u0_u14_X_2 ) , .ZN( u0_u14_u0_n103 ) , .A1( u0_u14_u0_n164 ) );
  NOR2_X1 u0_u14_u0_U57 (.A2( u0_u14_X_1 ) , .A1( u0_u14_X_2 ) , .ZN( u0_u14_u0_n92 ) );
  NOR2_X1 u0_u14_u0_U58 (.A2( u0_u14_X_1 ) , .ZN( u0_u14_u0_n101 ) , .A1( u0_u14_u0_n163 ) );
  NAND2_X1 u0_u14_u0_U59 (.A2( u0_u14_X_4 ) , .A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n144 ) );
  NOR2_X1 u0_u14_u0_U6 (.A1( u0_u14_u0_n108 ) , .ZN( u0_u14_u0_n123 ) , .A2( u0_u14_u0_n158 ) );
  NOR2_X1 u0_u14_u0_U60 (.A2( u0_u14_X_5 ) , .ZN( u0_u14_u0_n136 ) , .A1( u0_u14_u0_n159 ) );
  NAND2_X1 u0_u14_u0_U61 (.A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n138 ) , .A2( u0_u14_u0_n159 ) );
  AND2_X1 u0_u14_u0_U62 (.A2( u0_u14_X_3 ) , .A1( u0_u14_X_6 ) , .ZN( u0_u14_u0_n102 ) );
  AND2_X1 u0_u14_u0_U63 (.A1( u0_u14_X_6 ) , .A2( u0_u14_u0_n162 ) , .ZN( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U64 (.A( u0_u14_X_4 ) , .ZN( u0_u14_u0_n159 ) );
  INV_X1 u0_u14_u0_U65 (.A( u0_u14_X_1 ) , .ZN( u0_u14_u0_n164 ) );
  INV_X1 u0_u14_u0_U66 (.A( u0_u14_X_2 ) , .ZN( u0_u14_u0_n163 ) );
  INV_X1 u0_u14_u0_U67 (.A( u0_u14_X_3 ) , .ZN( u0_u14_u0_n162 ) );
  INV_X1 u0_u14_u0_U68 (.A( u0_u14_u0_n126 ) , .ZN( u0_u14_u0_n168 ) );
  AOI211_X1 u0_u14_u0_U69 (.B( u0_u14_u0_n133 ) , .A( u0_u14_u0_n134 ) , .C2( u0_u14_u0_n135 ) , .C1( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n137 ) );
  OAI21_X1 u0_u14_u0_U7 (.B1( u0_u14_u0_n150 ) , .B2( u0_u14_u0_n158 ) , .A( u0_u14_u0_n172 ) , .ZN( u0_u14_u0_n89 ) );
  INV_X1 u0_u14_u0_U70 (.ZN( u0_u14_u0_n174 ) , .A( u0_u14_u0_n89 ) );
  AOI211_X1 u0_u14_u0_U71 (.B( u0_u14_u0_n104 ) , .A( u0_u14_u0_n105 ) , .ZN( u0_u14_u0_n106 ) , .C2( u0_u14_u0_n113 ) , .C1( u0_u14_u0_n160 ) );
  OR4_X1 u0_u14_u0_U72 (.ZN( u0_out14_31 ) , .A4( u0_u14_u0_n155 ) , .A2( u0_u14_u0_n156 ) , .A1( u0_u14_u0_n157 ) , .A3( u0_u14_u0_n173 ) );
  AOI21_X1 u0_u14_u0_U73 (.A( u0_u14_u0_n138 ) , .B2( u0_u14_u0_n139 ) , .B1( u0_u14_u0_n140 ) , .ZN( u0_u14_u0_n157 ) );
  AOI21_X1 u0_u14_u0_U74 (.B2( u0_u14_u0_n141 ) , .B1( u0_u14_u0_n142 ) , .ZN( u0_u14_u0_n156 ) , .A( u0_u14_u0_n161 ) );
  OR4_X1 u0_u14_u0_U75 (.ZN( u0_out14_17 ) , .A4( u0_u14_u0_n122 ) , .A2( u0_u14_u0_n123 ) , .A1( u0_u14_u0_n124 ) , .A3( u0_u14_u0_n170 ) );
  AOI21_X1 u0_u14_u0_U76 (.B2( u0_u14_u0_n107 ) , .ZN( u0_u14_u0_n124 ) , .B1( u0_u14_u0_n128 ) , .A( u0_u14_u0_n161 ) );
  INV_X1 u0_u14_u0_U77 (.A( u0_u14_u0_n111 ) , .ZN( u0_u14_u0_n170 ) );
  AOI21_X1 u0_u14_u0_U78 (.B1( u0_u14_u0_n132 ) , .ZN( u0_u14_u0_n133 ) , .A( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n166 ) );
  OAI22_X1 u0_u14_u0_U79 (.ZN( u0_u14_u0_n105 ) , .A2( u0_u14_u0_n132 ) , .B1( u0_u14_u0_n146 ) , .A1( u0_u14_u0_n147 ) , .B2( u0_u14_u0_n161 ) );
  AND2_X1 u0_u14_u0_U8 (.A1( u0_u14_u0_n114 ) , .A2( u0_u14_u0_n121 ) , .ZN( u0_u14_u0_n146 ) );
  NAND2_X1 u0_u14_u0_U80 (.ZN( u0_u14_u0_n110 ) , .A2( u0_u14_u0_n132 ) , .A1( u0_u14_u0_n145 ) );
  INV_X1 u0_u14_u0_U81 (.A( u0_u14_u0_n119 ) , .ZN( u0_u14_u0_n167 ) );
  NAND2_X1 u0_u14_u0_U82 (.A2( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n140 ) , .A1( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U83 (.A1( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n130 ) , .A2( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U84 (.ZN( u0_u14_u0_n108 ) , .A1( u0_u14_u0_n92 ) , .A2( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U85 (.ZN( u0_u14_u0_n142 ) , .A1( u0_u14_u0_n94 ) , .A2( u0_u14_u0_n95 ) );
  NOR2_X1 u0_u14_u0_U86 (.A2( u0_u14_X_6 ) , .ZN( u0_u14_u0_n100 ) , .A1( u0_u14_u0_n162 ) );
  NOR2_X1 u0_u14_u0_U87 (.A2( u0_u14_X_3 ) , .A1( u0_u14_X_6 ) , .ZN( u0_u14_u0_n94 ) );
  NAND3_X1 u0_u14_u0_U88 (.ZN( u0_out14_23 ) , .A3( u0_u14_u0_n137 ) , .A1( u0_u14_u0_n168 ) , .A2( u0_u14_u0_n171 ) );
  NAND3_X1 u0_u14_u0_U89 (.A3( u0_u14_u0_n127 ) , .A2( u0_u14_u0_n128 ) , .ZN( u0_u14_u0_n135 ) , .A1( u0_u14_u0_n150 ) );
  AND2_X1 u0_u14_u0_U9 (.A1( u0_u14_u0_n131 ) , .ZN( u0_u14_u0_n141 ) , .A2( u0_u14_u0_n150 ) );
  NAND3_X1 u0_u14_u0_U90 (.ZN( u0_u14_u0_n117 ) , .A3( u0_u14_u0_n132 ) , .A2( u0_u14_u0_n139 ) , .A1( u0_u14_u0_n148 ) );
  NAND3_X1 u0_u14_u0_U91 (.ZN( u0_u14_u0_n109 ) , .A2( u0_u14_u0_n114 ) , .A3( u0_u14_u0_n140 ) , .A1( u0_u14_u0_n149 ) );
  NAND3_X1 u0_u14_u0_U92 (.ZN( u0_out14_9 ) , .A3( u0_u14_u0_n106 ) , .A2( u0_u14_u0_n171 ) , .A1( u0_u14_u0_n174 ) );
  NAND3_X1 u0_u14_u0_U93 (.A2( u0_u14_u0_n128 ) , .A1( u0_u14_u0_n132 ) , .A3( u0_u14_u0_n146 ) , .ZN( u0_u14_u0_n97 ) );
  XOR2_X1 u0_u15_U1 (.A( u0_FP_38 ) , .B( u0_K16_9 ) , .Z( u0_u15_X_9 ) );
  XOR2_X1 u0_u15_U10 (.A( u0_FP_62 ) , .B( u0_K16_45 ) , .Z( u0_u15_X_45 ) );
  XOR2_X1 u0_u15_U11 (.A( u0_FP_61 ) , .B( u0_K16_44 ) , .Z( u0_u15_X_44 ) );
  XOR2_X1 u0_u15_U13 (.A( u0_FP_61 ) , .B( u0_K16_42 ) , .Z( u0_u15_X_42 ) );
  XOR2_X1 u0_u15_U23 (.A( u0_FP_54 ) , .B( u0_K16_33 ) , .Z( u0_u15_X_33 ) );
  XOR2_X1 u0_u15_U35 (.A( u0_FP_47 ) , .B( u0_K16_22 ) , .Z( u0_u15_X_22 ) );
  XOR2_X1 u0_u15_U45 (.A( u0_FP_40 ) , .B( u0_K16_13 ) , .Z( u0_u15_X_13 ) );
  XOR2_X1 u0_u15_U47 (.A( u0_FP_40 ) , .B( u0_K16_11 ) , .Z( u0_u15_X_11 ) );
  XOR2_X1 u0_u15_U6 (.A( u0_FP_35 ) , .B( u0_K16_4 ) , .Z( u0_u15_X_4 ) );
  XOR2_X1 u0_u1_U1 (.B( u0_K2_9 ) , .A( u0_R0_6 ) , .Z( u0_u1_X_9 ) );
  XOR2_X1 u0_u1_U10 (.B( u0_K2_45 ) , .A( u0_R0_30 ) , .Z( u0_u1_X_45 ) );
  XOR2_X1 u0_u1_U11 (.B( u0_K2_44 ) , .A( u0_R0_29 ) , .Z( u0_u1_X_44 ) );
  XOR2_X1 u0_u1_U12 (.B( u0_K2_43 ) , .A( u0_R0_28 ) , .Z( u0_u1_X_43 ) );
  XOR2_X1 u0_u1_U13 (.B( u0_K2_42 ) , .A( u0_R0_29 ) , .Z( u0_u1_X_42 ) );
  XOR2_X1 u0_u1_U15 (.B( u0_K2_40 ) , .A( u0_R0_27 ) , .Z( u0_u1_X_40 ) );
  XOR2_X1 u0_u1_U16 (.B( u0_K2_3 ) , .A( u0_R0_2 ) , .Z( u0_u1_X_3 ) );
  XOR2_X1 u0_u1_U17 (.B( u0_K2_39 ) , .A( u0_R0_26 ) , .Z( u0_u1_X_39 ) );
  XOR2_X1 u0_u1_U18 (.B( u0_K2_38 ) , .A( u0_R0_25 ) , .Z( u0_u1_X_38 ) );
  XOR2_X1 u0_u1_U19 (.B( u0_K2_37 ) , .A( u0_R0_24 ) , .Z( u0_u1_X_37 ) );
  XOR2_X1 u0_u1_U2 (.B( u0_K2_8 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_8 ) );
  XOR2_X1 u0_u1_U20 (.B( u0_K2_36 ) , .A( u0_R0_25 ) , .Z( u0_u1_X_36 ) );
  XOR2_X1 u0_u1_U21 (.B( u0_K2_35 ) , .A( u0_R0_24 ) , .Z( u0_u1_X_35 ) );
  XOR2_X1 u0_u1_U22 (.B( u0_K2_34 ) , .A( u0_R0_23 ) , .Z( u0_u1_X_34 ) );
  XOR2_X1 u0_u1_U23 (.B( u0_K2_33 ) , .A( u0_R0_22 ) , .Z( u0_u1_X_33 ) );
  XOR2_X1 u0_u1_U31 (.B( u0_K2_26 ) , .A( u0_R0_17 ) , .Z( u0_u1_X_26 ) );
  XOR2_X1 u0_u1_U32 (.B( u0_K2_25 ) , .A( u0_R0_16 ) , .Z( u0_u1_X_25 ) );
  XOR2_X1 u0_u1_U33 (.B( u0_K2_24 ) , .A( u0_R0_17 ) , .Z( u0_u1_X_24 ) );
  XOR2_X1 u0_u1_U34 (.B( u0_K2_23 ) , .A( u0_R0_16 ) , .Z( u0_u1_X_23 ) );
  XOR2_X1 u0_u1_U36 (.B( u0_K2_21 ) , .A( u0_R0_14 ) , .Z( u0_u1_X_21 ) );
  XOR2_X1 u0_u1_U39 (.B( u0_K2_19 ) , .A( u0_R0_12 ) , .Z( u0_u1_X_19 ) );
  XOR2_X1 u0_u1_U4 (.B( u0_K2_6 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_6 ) );
  XOR2_X1 u0_u1_U41 (.B( u0_K2_17 ) , .A( u0_R0_12 ) , .Z( u0_u1_X_17 ) );
  XOR2_X1 u0_u1_U42 (.B( u0_K2_16 ) , .A( u0_R0_11 ) , .Z( u0_u1_X_16 ) );
  XOR2_X1 u0_u1_U43 (.B( u0_K2_15 ) , .A( u0_R0_10 ) , .Z( u0_u1_X_15 ) );
  XOR2_X1 u0_u1_U6 (.B( u0_K2_4 ) , .A( u0_R0_3 ) , .Z( u0_u1_X_4 ) );
  XOR2_X1 u0_u1_U7 (.B( u0_K2_48 ) , .A( u0_R0_1 ) , .Z( u0_u1_X_48 ) );
  XOR2_X1 u0_u1_U8 (.B( u0_K2_47 ) , .A( u0_R0_32 ) , .Z( u0_u1_X_47 ) );
  XOR2_X1 u0_u1_U9 (.B( u0_K2_46 ) , .A( u0_R0_31 ) , .Z( u0_u1_X_46 ) );
  AND3_X1 u0_u1_u7_U10 (.A3( u0_u1_u7_n110 ) , .A2( u0_u1_u7_n127 ) , .A1( u0_u1_u7_n132 ) , .ZN( u0_u1_u7_n92 ) );
  OAI21_X1 u0_u1_u7_U11 (.A( u0_u1_u7_n161 ) , .B1( u0_u1_u7_n168 ) , .B2( u0_u1_u7_n173 ) , .ZN( u0_u1_u7_n91 ) );
  AOI211_X1 u0_u1_u7_U12 (.A( u0_u1_u7_n117 ) , .ZN( u0_u1_u7_n118 ) , .C2( u0_u1_u7_n126 ) , .C1( u0_u1_u7_n177 ) , .B( u0_u1_u7_n180 ) );
  OAI22_X1 u0_u1_u7_U13 (.B1( u0_u1_u7_n115 ) , .ZN( u0_u1_u7_n117 ) , .A2( u0_u1_u7_n133 ) , .A1( u0_u1_u7_n137 ) , .B2( u0_u1_u7_n162 ) );
  INV_X1 u0_u1_u7_U14 (.A( u0_u1_u7_n116 ) , .ZN( u0_u1_u7_n180 ) );
  NOR3_X1 u0_u1_u7_U15 (.ZN( u0_u1_u7_n115 ) , .A3( u0_u1_u7_n145 ) , .A2( u0_u1_u7_n168 ) , .A1( u0_u1_u7_n169 ) );
  OAI211_X1 u0_u1_u7_U16 (.B( u0_u1_u7_n122 ) , .A( u0_u1_u7_n123 ) , .C2( u0_u1_u7_n124 ) , .ZN( u0_u1_u7_n154 ) , .C1( u0_u1_u7_n162 ) );
  AOI222_X1 u0_u1_u7_U17 (.ZN( u0_u1_u7_n122 ) , .C2( u0_u1_u7_n126 ) , .C1( u0_u1_u7_n145 ) , .B1( u0_u1_u7_n161 ) , .A2( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n170 ) , .A1( u0_u1_u7_n176 ) );
  INV_X1 u0_u1_u7_U18 (.A( u0_u1_u7_n133 ) , .ZN( u0_u1_u7_n176 ) );
  NOR3_X1 u0_u1_u7_U19 (.A2( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n135 ) , .ZN( u0_u1_u7_n136 ) , .A3( u0_u1_u7_n171 ) );
  NOR2_X1 u0_u1_u7_U20 (.A1( u0_u1_u7_n130 ) , .A2( u0_u1_u7_n134 ) , .ZN( u0_u1_u7_n153 ) );
  INV_X1 u0_u1_u7_U21 (.A( u0_u1_u7_n101 ) , .ZN( u0_u1_u7_n165 ) );
  NOR2_X1 u0_u1_u7_U22 (.ZN( u0_u1_u7_n111 ) , .A2( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n169 ) );
  AOI21_X1 u0_u1_u7_U23 (.ZN( u0_u1_u7_n104 ) , .B2( u0_u1_u7_n112 ) , .B1( u0_u1_u7_n127 ) , .A( u0_u1_u7_n164 ) );
  AOI21_X1 u0_u1_u7_U24 (.ZN( u0_u1_u7_n106 ) , .B1( u0_u1_u7_n133 ) , .B2( u0_u1_u7_n146 ) , .A( u0_u1_u7_n162 ) );
  AOI21_X1 u0_u1_u7_U25 (.A( u0_u1_u7_n101 ) , .ZN( u0_u1_u7_n107 ) , .B2( u0_u1_u7_n128 ) , .B1( u0_u1_u7_n175 ) );
  INV_X1 u0_u1_u7_U26 (.A( u0_u1_u7_n138 ) , .ZN( u0_u1_u7_n171 ) );
  INV_X1 u0_u1_u7_U27 (.A( u0_u1_u7_n131 ) , .ZN( u0_u1_u7_n177 ) );
  INV_X1 u0_u1_u7_U28 (.A( u0_u1_u7_n110 ) , .ZN( u0_u1_u7_n174 ) );
  NAND2_X1 u0_u1_u7_U29 (.A1( u0_u1_u7_n129 ) , .A2( u0_u1_u7_n132 ) , .ZN( u0_u1_u7_n149 ) );
  OAI21_X1 u0_u1_u7_U3 (.ZN( u0_u1_u7_n159 ) , .A( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n171 ) , .B1( u0_u1_u7_n174 ) );
  NAND2_X1 u0_u1_u7_U30 (.A1( u0_u1_u7_n113 ) , .A2( u0_u1_u7_n124 ) , .ZN( u0_u1_u7_n130 ) );
  INV_X1 u0_u1_u7_U31 (.A( u0_u1_u7_n112 ) , .ZN( u0_u1_u7_n173 ) );
  INV_X1 u0_u1_u7_U32 (.A( u0_u1_u7_n128 ) , .ZN( u0_u1_u7_n168 ) );
  INV_X1 u0_u1_u7_U33 (.A( u0_u1_u7_n148 ) , .ZN( u0_u1_u7_n169 ) );
  INV_X1 u0_u1_u7_U34 (.A( u0_u1_u7_n127 ) , .ZN( u0_u1_u7_n179 ) );
  NOR2_X1 u0_u1_u7_U35 (.ZN( u0_u1_u7_n101 ) , .A2( u0_u1_u7_n150 ) , .A1( u0_u1_u7_n156 ) );
  AOI211_X1 u0_u1_u7_U36 (.B( u0_u1_u7_n154 ) , .A( u0_u1_u7_n155 ) , .C1( u0_u1_u7_n156 ) , .ZN( u0_u1_u7_n157 ) , .C2( u0_u1_u7_n172 ) );
  INV_X1 u0_u1_u7_U37 (.A( u0_u1_u7_n153 ) , .ZN( u0_u1_u7_n172 ) );
  AOI211_X1 u0_u1_u7_U38 (.B( u0_u1_u7_n139 ) , .A( u0_u1_u7_n140 ) , .C2( u0_u1_u7_n141 ) , .ZN( u0_u1_u7_n142 ) , .C1( u0_u1_u7_n156 ) );
  NAND4_X1 u0_u1_u7_U39 (.A3( u0_u1_u7_n127 ) , .A2( u0_u1_u7_n128 ) , .A1( u0_u1_u7_n129 ) , .ZN( u0_u1_u7_n141 ) , .A4( u0_u1_u7_n147 ) );
  INV_X1 u0_u1_u7_U4 (.A( u0_u1_u7_n111 ) , .ZN( u0_u1_u7_n170 ) );
  AOI21_X1 u0_u1_u7_U40 (.A( u0_u1_u7_n137 ) , .B1( u0_u1_u7_n138 ) , .ZN( u0_u1_u7_n139 ) , .B2( u0_u1_u7_n146 ) );
  OAI22_X1 u0_u1_u7_U41 (.B1( u0_u1_u7_n136 ) , .ZN( u0_u1_u7_n140 ) , .A1( u0_u1_u7_n153 ) , .B2( u0_u1_u7_n162 ) , .A2( u0_u1_u7_n164 ) );
  AOI21_X1 u0_u1_u7_U42 (.ZN( u0_u1_u7_n123 ) , .B1( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n177 ) , .A( u0_u1_u7_n97 ) );
  AOI21_X1 u0_u1_u7_U43 (.B2( u0_u1_u7_n113 ) , .B1( u0_u1_u7_n124 ) , .A( u0_u1_u7_n125 ) , .ZN( u0_u1_u7_n97 ) );
  INV_X1 u0_u1_u7_U44 (.A( u0_u1_u7_n125 ) , .ZN( u0_u1_u7_n161 ) );
  INV_X1 u0_u1_u7_U45 (.A( u0_u1_u7_n152 ) , .ZN( u0_u1_u7_n162 ) );
  AOI22_X1 u0_u1_u7_U46 (.A2( u0_u1_u7_n114 ) , .ZN( u0_u1_u7_n119 ) , .B1( u0_u1_u7_n130 ) , .A1( u0_u1_u7_n156 ) , .B2( u0_u1_u7_n165 ) );
  NAND2_X1 u0_u1_u7_U47 (.A2( u0_u1_u7_n112 ) , .ZN( u0_u1_u7_n114 ) , .A1( u0_u1_u7_n175 ) );
  AND2_X1 u0_u1_u7_U48 (.ZN( u0_u1_u7_n145 ) , .A2( u0_u1_u7_n98 ) , .A1( u0_u1_u7_n99 ) );
  NOR2_X1 u0_u1_u7_U49 (.ZN( u0_u1_u7_n137 ) , .A1( u0_u1_u7_n150 ) , .A2( u0_u1_u7_n161 ) );
  INV_X1 u0_u1_u7_U5 (.A( u0_u1_u7_n149 ) , .ZN( u0_u1_u7_n175 ) );
  AOI21_X1 u0_u1_u7_U50 (.ZN( u0_u1_u7_n105 ) , .B2( u0_u1_u7_n110 ) , .A( u0_u1_u7_n125 ) , .B1( u0_u1_u7_n147 ) );
  NAND2_X1 u0_u1_u7_U51 (.ZN( u0_u1_u7_n146 ) , .A1( u0_u1_u7_n95 ) , .A2( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U52 (.A2( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n147 ) , .A1( u0_u1_u7_n93 ) );
  NAND2_X1 u0_u1_u7_U53 (.A1( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n127 ) , .A2( u0_u1_u7_n99 ) );
  OR2_X1 u0_u1_u7_U54 (.ZN( u0_u1_u7_n126 ) , .A2( u0_u1_u7_n152 ) , .A1( u0_u1_u7_n156 ) );
  NAND2_X1 u0_u1_u7_U55 (.A2( u0_u1_u7_n102 ) , .A1( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n133 ) );
  NAND2_X1 u0_u1_u7_U56 (.ZN( u0_u1_u7_n112 ) , .A2( u0_u1_u7_n96 ) , .A1( u0_u1_u7_n99 ) );
  NAND2_X1 u0_u1_u7_U57 (.A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n128 ) , .A1( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U58 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n113 ) , .A2( u0_u1_u7_n93 ) );
  NAND2_X1 u0_u1_u7_U59 (.A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n124 ) , .A1( u0_u1_u7_n96 ) );
  INV_X1 u0_u1_u7_U6 (.A( u0_u1_u7_n154 ) , .ZN( u0_u1_u7_n178 ) );
  NAND2_X1 u0_u1_u7_U60 (.ZN( u0_u1_u7_n110 ) , .A1( u0_u1_u7_n95 ) , .A2( u0_u1_u7_n96 ) );
  INV_X1 u0_u1_u7_U61 (.A( u0_u1_u7_n150 ) , .ZN( u0_u1_u7_n164 ) );
  AND2_X1 u0_u1_u7_U62 (.ZN( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n93 ) , .A2( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U63 (.A1( u0_u1_u7_n100 ) , .A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n129 ) );
  NAND2_X1 u0_u1_u7_U64 (.A2( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n131 ) , .A1( u0_u1_u7_n95 ) );
  NAND2_X1 u0_u1_u7_U65 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n138 ) , .A2( u0_u1_u7_n99 ) );
  NAND2_X1 u0_u1_u7_U66 (.ZN( u0_u1_u7_n132 ) , .A1( u0_u1_u7_n93 ) , .A2( u0_u1_u7_n96 ) );
  NAND2_X1 u0_u1_u7_U67 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n148 ) , .A2( u0_u1_u7_n95 ) );
  NOR2_X1 u0_u1_u7_U68 (.A2( u0_u1_X_47 ) , .ZN( u0_u1_u7_n150 ) , .A1( u0_u1_u7_n163 ) );
  NOR2_X1 u0_u1_u7_U69 (.A2( u0_u1_X_43 ) , .A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n103 ) );
  AOI211_X1 u0_u1_u7_U7 (.ZN( u0_u1_u7_n116 ) , .A( u0_u1_u7_n155 ) , .C1( u0_u1_u7_n161 ) , .C2( u0_u1_u7_n171 ) , .B( u0_u1_u7_n94 ) );
  NOR2_X1 u0_u1_u7_U70 (.A2( u0_u1_X_48 ) , .A1( u0_u1_u7_n166 ) , .ZN( u0_u1_u7_n95 ) );
  NOR2_X1 u0_u1_u7_U71 (.A2( u0_u1_X_45 ) , .A1( u0_u1_X_48 ) , .ZN( u0_u1_u7_n99 ) );
  NOR2_X1 u0_u1_u7_U72 (.A2( u0_u1_X_44 ) , .A1( u0_u1_u7_n167 ) , .ZN( u0_u1_u7_n98 ) );
  NOR2_X1 u0_u1_u7_U73 (.A2( u0_u1_X_46 ) , .A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n152 ) );
  AND2_X1 u0_u1_u7_U74 (.A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n156 ) , .A2( u0_u1_u7_n163 ) );
  NAND2_X1 u0_u1_u7_U75 (.A2( u0_u1_X_46 ) , .A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n125 ) );
  AND2_X1 u0_u1_u7_U76 (.A2( u0_u1_X_45 ) , .A1( u0_u1_X_48 ) , .ZN( u0_u1_u7_n102 ) );
  AND2_X1 u0_u1_u7_U77 (.A2( u0_u1_X_43 ) , .A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n96 ) );
  AND2_X1 u0_u1_u7_U78 (.A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n100 ) , .A2( u0_u1_u7_n167 ) );
  AND2_X1 u0_u1_u7_U79 (.A1( u0_u1_X_48 ) , .A2( u0_u1_u7_n166 ) , .ZN( u0_u1_u7_n93 ) );
  OAI222_X1 u0_u1_u7_U8 (.C2( u0_u1_u7_n101 ) , .B2( u0_u1_u7_n111 ) , .A1( u0_u1_u7_n113 ) , .C1( u0_u1_u7_n146 ) , .A2( u0_u1_u7_n162 ) , .B1( u0_u1_u7_n164 ) , .ZN( u0_u1_u7_n94 ) );
  INV_X1 u0_u1_u7_U80 (.A( u0_u1_X_46 ) , .ZN( u0_u1_u7_n163 ) );
  INV_X1 u0_u1_u7_U81 (.A( u0_u1_X_43 ) , .ZN( u0_u1_u7_n167 ) );
  INV_X1 u0_u1_u7_U82 (.A( u0_u1_X_45 ) , .ZN( u0_u1_u7_n166 ) );
  NAND4_X1 u0_u1_u7_U83 (.ZN( u0_out1_27 ) , .A4( u0_u1_u7_n118 ) , .A3( u0_u1_u7_n119 ) , .A2( u0_u1_u7_n120 ) , .A1( u0_u1_u7_n121 ) );
  OAI21_X1 u0_u1_u7_U84 (.ZN( u0_u1_u7_n121 ) , .B2( u0_u1_u7_n145 ) , .A( u0_u1_u7_n150 ) , .B1( u0_u1_u7_n174 ) );
  OAI21_X1 u0_u1_u7_U85 (.ZN( u0_u1_u7_n120 ) , .A( u0_u1_u7_n161 ) , .B2( u0_u1_u7_n170 ) , .B1( u0_u1_u7_n179 ) );
  NAND4_X1 u0_u1_u7_U86 (.ZN( u0_out1_15 ) , .A4( u0_u1_u7_n142 ) , .A3( u0_u1_u7_n143 ) , .A2( u0_u1_u7_n144 ) , .A1( u0_u1_u7_n178 ) );
  OR2_X1 u0_u1_u7_U87 (.A2( u0_u1_u7_n125 ) , .A1( u0_u1_u7_n129 ) , .ZN( u0_u1_u7_n144 ) );
  AOI22_X1 u0_u1_u7_U88 (.A2( u0_u1_u7_n126 ) , .ZN( u0_u1_u7_n143 ) , .B2( u0_u1_u7_n165 ) , .B1( u0_u1_u7_n173 ) , .A1( u0_u1_u7_n174 ) );
  NAND4_X1 u0_u1_u7_U89 (.ZN( u0_out1_5 ) , .A4( u0_u1_u7_n108 ) , .A3( u0_u1_u7_n109 ) , .A1( u0_u1_u7_n116 ) , .A2( u0_u1_u7_n123 ) );
  OAI221_X1 u0_u1_u7_U9 (.C1( u0_u1_u7_n101 ) , .C2( u0_u1_u7_n147 ) , .ZN( u0_u1_u7_n155 ) , .B2( u0_u1_u7_n162 ) , .A( u0_u1_u7_n91 ) , .B1( u0_u1_u7_n92 ) );
  AOI22_X1 u0_u1_u7_U90 (.ZN( u0_u1_u7_n109 ) , .A2( u0_u1_u7_n126 ) , .B2( u0_u1_u7_n145 ) , .B1( u0_u1_u7_n156 ) , .A1( u0_u1_u7_n171 ) );
  NOR4_X1 u0_u1_u7_U91 (.A4( u0_u1_u7_n104 ) , .A3( u0_u1_u7_n105 ) , .A2( u0_u1_u7_n106 ) , .A1( u0_u1_u7_n107 ) , .ZN( u0_u1_u7_n108 ) );
  NAND4_X1 u0_u1_u7_U92 (.ZN( u0_out1_21 ) , .A4( u0_u1_u7_n157 ) , .A3( u0_u1_u7_n158 ) , .A2( u0_u1_u7_n159 ) , .A1( u0_u1_u7_n160 ) );
  OAI21_X1 u0_u1_u7_U93 (.B1( u0_u1_u7_n145 ) , .ZN( u0_u1_u7_n160 ) , .A( u0_u1_u7_n161 ) , .B2( u0_u1_u7_n177 ) );
  AOI22_X1 u0_u1_u7_U94 (.B2( u0_u1_u7_n149 ) , .B1( u0_u1_u7_n150 ) , .A2( u0_u1_u7_n151 ) , .A1( u0_u1_u7_n152 ) , .ZN( u0_u1_u7_n158 ) );
  NAND3_X1 u0_u1_u7_U95 (.A3( u0_u1_u7_n146 ) , .A2( u0_u1_u7_n147 ) , .A1( u0_u1_u7_n148 ) , .ZN( u0_u1_u7_n151 ) );
  NAND3_X1 u0_u1_u7_U96 (.A3( u0_u1_u7_n131 ) , .A2( u0_u1_u7_n132 ) , .A1( u0_u1_u7_n133 ) , .ZN( u0_u1_u7_n135 ) );
  XOR2_X1 u0_u2_U1 (.B( u0_K3_9 ) , .A( u0_R1_6 ) , .Z( u0_u2_X_9 ) );
  XOR2_X1 u0_u2_U16 (.B( u0_K3_3 ) , .A( u0_R1_2 ) , .Z( u0_u2_X_3 ) );
  XOR2_X1 u0_u2_U22 (.B( u0_K3_34 ) , .A( u0_R1_23 ) , .Z( u0_u2_X_34 ) );
  XOR2_X1 u0_u2_U30 (.B( u0_K3_27 ) , .A( u0_R1_18 ) , .Z( u0_u2_X_27 ) );
  XOR2_X1 u0_u2_U31 (.B( u0_K3_26 ) , .A( u0_R1_17 ) , .Z( u0_u2_X_26 ) );
  XOR2_X1 u0_u2_U33 (.B( u0_K3_24 ) , .A( u0_R1_17 ) , .Z( u0_u2_X_24 ) );
  XOR2_X1 u0_u2_U42 (.B( u0_K3_16 ) , .A( u0_R1_11 ) , .Z( u0_u2_X_16 ) );
  XOR2_X1 u0_u2_U43 (.B( u0_K3_15 ) , .A( u0_R1_10 ) , .Z( u0_u2_X_15 ) );
  XOR2_X1 u0_u2_U48 (.B( u0_K3_10 ) , .A( u0_R1_7 ) , .Z( u0_u2_X_10 ) );
  XOR2_X1 u0_u2_U9 (.B( u0_K3_46 ) , .A( u0_R1_31 ) , .Z( u0_u2_X_46 ) );
  XOR2_X1 u0_u3_U10 (.B( u0_K4_45 ) , .A( u0_R2_30 ) , .Z( u0_u3_X_45 ) );
  XOR2_X1 u0_u3_U11 (.B( u0_K4_44 ) , .A( u0_R2_29 ) , .Z( u0_u3_X_44 ) );
  XOR2_X1 u0_u3_U13 (.B( u0_K4_42 ) , .A( u0_R2_29 ) , .Z( u0_u3_X_42 ) );
  XOR2_X1 u0_u3_U15 (.B( u0_K4_40 ) , .A( u0_R2_27 ) , .Z( u0_u3_X_40 ) );
  XOR2_X1 u0_u3_U17 (.B( u0_K4_39 ) , .A( u0_R2_26 ) , .Z( u0_u3_X_39 ) );
  XOR2_X1 u0_u3_U19 (.B( u0_K4_37 ) , .A( u0_R2_24 ) , .Z( u0_u3_X_37 ) );
  XOR2_X1 u0_u3_U21 (.B( u0_K4_35 ) , .A( u0_R2_24 ) , .Z( u0_u3_X_35 ) );
  XOR2_X1 u0_u3_U22 (.B( u0_K4_34 ) , .A( u0_R2_23 ) , .Z( u0_u3_X_34 ) );
  XOR2_X1 u0_u3_U25 (.B( u0_K4_31 ) , .A( u0_R2_20 ) , .Z( u0_u3_X_31 ) );
  XOR2_X1 u0_u3_U28 (.B( u0_K4_29 ) , .A( u0_R2_20 ) , .Z( u0_u3_X_29 ) );
  XOR2_X1 u0_u3_U29 (.B( u0_K4_28 ) , .A( u0_R2_19 ) , .Z( u0_u3_X_28 ) );
  XOR2_X1 u0_u3_U30 (.B( u0_K4_27 ) , .A( u0_R2_18 ) , .Z( u0_u3_X_27 ) );
  XOR2_X1 u0_u3_U31 (.B( u0_K4_26 ) , .A( u0_R2_17 ) , .Z( u0_u3_X_26 ) );
  XOR2_X1 u0_u3_U33 (.B( u0_K4_24 ) , .A( u0_R2_17 ) , .Z( u0_u3_X_24 ) );
  XOR2_X1 u0_u3_U35 (.B( u0_K4_22 ) , .A( u0_R2_15 ) , .Z( u0_u3_X_22 ) );
  XOR2_X1 u0_u3_U9 (.B( u0_K4_46 ) , .A( u0_R2_31 ) , .Z( u0_u3_X_46 ) );
  XOR2_X1 u0_u4_U1 (.B( u0_K5_9 ) , .A( u0_R3_6 ) , .Z( u0_u4_X_9 ) );
  XOR2_X1 u0_u4_U10 (.B( u0_K5_45 ) , .A( u0_R3_30 ) , .Z( u0_u4_X_45 ) );
  XOR2_X1 u0_u4_U11 (.B( u0_K5_44 ) , .A( u0_R3_29 ) , .Z( u0_u4_X_44 ) );
  XOR2_X1 u0_u4_U12 (.B( u0_K5_43 ) , .A( u0_R3_28 ) , .Z( u0_u4_X_43 ) );
  XOR2_X1 u0_u4_U13 (.B( u0_K5_42 ) , .A( u0_R3_29 ) , .Z( u0_u4_X_42 ) );
  XOR2_X1 u0_u4_U14 (.B( u0_K5_41 ) , .A( u0_R3_28 ) , .Z( u0_u4_X_41 ) );
  XOR2_X1 u0_u4_U15 (.B( u0_K5_40 ) , .A( u0_R3_27 ) , .Z( u0_u4_X_40 ) );
  XOR2_X1 u0_u4_U16 (.B( u0_K5_3 ) , .A( u0_R3_2 ) , .Z( u0_u4_X_3 ) );
  XOR2_X1 u0_u4_U17 (.B( u0_K5_39 ) , .A( u0_R3_26 ) , .Z( u0_u4_X_39 ) );
  XOR2_X1 u0_u4_U18 (.B( u0_K5_38 ) , .A( u0_R3_25 ) , .Z( u0_u4_X_38 ) );
  XOR2_X1 u0_u4_U19 (.B( u0_K5_37 ) , .A( u0_R3_24 ) , .Z( u0_u4_X_37 ) );
  XOR2_X1 u0_u4_U22 (.B( u0_K5_34 ) , .A( u0_R3_23 ) , .Z( u0_u4_X_34 ) );
  XOR2_X1 u0_u4_U24 (.B( u0_K5_32 ) , .A( u0_R3_21 ) , .Z( u0_u4_X_32 ) );
  XOR2_X1 u0_u4_U26 (.B( u0_K5_30 ) , .A( u0_R3_21 ) , .Z( u0_u4_X_30 ) );
  XOR2_X1 u0_u4_U27 (.B( u0_K5_2 ) , .A( u0_R3_1 ) , .Z( u0_u4_X_2 ) );
  XOR2_X1 u0_u4_U29 (.B( u0_K5_28 ) , .A( u0_R3_19 ) , .Z( u0_u4_X_28 ) );
  XOR2_X1 u0_u4_U3 (.B( u0_K5_7 ) , .A( u0_R3_4 ) , .Z( u0_u4_X_7 ) );
  XOR2_X1 u0_u4_U32 (.B( u0_K5_25 ) , .A( u0_R3_16 ) , .Z( u0_u4_X_25 ) );
  XOR2_X1 u0_u4_U34 (.B( u0_K5_23 ) , .A( u0_R3_16 ) , .Z( u0_u4_X_23 ) );
  XOR2_X1 u0_u4_U36 (.B( u0_K5_21 ) , .A( u0_R3_14 ) , .Z( u0_u4_X_21 ) );
  XOR2_X1 u0_u4_U39 (.B( u0_K5_19 ) , .A( u0_R3_12 ) , .Z( u0_u4_X_19 ) );
  XOR2_X1 u0_u4_U41 (.B( u0_K5_17 ) , .A( u0_R3_12 ) , .Z( u0_u4_X_17 ) );
  XOR2_X1 u0_u4_U42 (.B( u0_K5_16 ) , .A( u0_R3_11 ) , .Z( u0_u4_X_16 ) );
  XOR2_X1 u0_u4_U43 (.B( u0_K5_15 ) , .A( u0_R3_10 ) , .Z( u0_u4_X_15 ) );
  XOR2_X1 u0_u4_U44 (.B( u0_K5_14 ) , .A( u0_R3_9 ) , .Z( u0_u4_X_14 ) );
  XOR2_X1 u0_u4_U45 (.B( u0_K5_13 ) , .A( u0_R3_8 ) , .Z( u0_u4_X_13 ) );
  XOR2_X1 u0_u4_U46 (.B( u0_K5_12 ) , .A( u0_R3_9 ) , .Z( u0_u4_X_12 ) );
  XOR2_X1 u0_u4_U47 (.B( u0_K5_11 ) , .A( u0_R3_8 ) , .Z( u0_u4_X_11 ) );
  XOR2_X1 u0_u4_U48 (.B( u0_K5_10 ) , .A( u0_R3_7 ) , .Z( u0_u4_X_10 ) );
  XOR2_X1 u0_u4_U5 (.B( u0_K5_5 ) , .A( u0_R3_4 ) , .Z( u0_u4_X_5 ) );
  XOR2_X1 u0_u4_U6 (.B( u0_K5_4 ) , .A( u0_R3_3 ) , .Z( u0_u4_X_4 ) );
  XOR2_X1 u0_u4_U7 (.B( u0_K5_48 ) , .A( u0_R3_1 ) , .Z( u0_u4_X_48 ) );
  XOR2_X1 u0_u4_U9 (.B( u0_K5_46 ) , .A( u0_R3_31 ) , .Z( u0_u4_X_46 ) );
  AOI22_X1 u0_u4_u6_U10 (.A2( u0_u4_u6_n151 ) , .B2( u0_u4_u6_n161 ) , .A1( u0_u4_u6_n167 ) , .B1( u0_u4_u6_n170 ) , .ZN( u0_u4_u6_n89 ) );
  AOI21_X1 u0_u4_u6_U11 (.B1( u0_u4_u6_n107 ) , .B2( u0_u4_u6_n132 ) , .A( u0_u4_u6_n158 ) , .ZN( u0_u4_u6_n88 ) );
  AOI21_X1 u0_u4_u6_U12 (.B2( u0_u4_u6_n147 ) , .B1( u0_u4_u6_n148 ) , .ZN( u0_u4_u6_n149 ) , .A( u0_u4_u6_n158 ) );
  AOI21_X1 u0_u4_u6_U13 (.ZN( u0_u4_u6_n106 ) , .A( u0_u4_u6_n142 ) , .B2( u0_u4_u6_n159 ) , .B1( u0_u4_u6_n164 ) );
  INV_X1 u0_u4_u6_U14 (.A( u0_u4_u6_n155 ) , .ZN( u0_u4_u6_n161 ) );
  INV_X1 u0_u4_u6_U15 (.A( u0_u4_u6_n128 ) , .ZN( u0_u4_u6_n164 ) );
  NAND2_X1 u0_u4_u6_U16 (.ZN( u0_u4_u6_n110 ) , .A1( u0_u4_u6_n122 ) , .A2( u0_u4_u6_n129 ) );
  NAND2_X1 u0_u4_u6_U17 (.ZN( u0_u4_u6_n124 ) , .A2( u0_u4_u6_n146 ) , .A1( u0_u4_u6_n148 ) );
  INV_X1 u0_u4_u6_U18 (.A( u0_u4_u6_n132 ) , .ZN( u0_u4_u6_n171 ) );
  AND2_X1 u0_u4_u6_U19 (.A1( u0_u4_u6_n100 ) , .ZN( u0_u4_u6_n130 ) , .A2( u0_u4_u6_n147 ) );
  INV_X1 u0_u4_u6_U20 (.A( u0_u4_u6_n127 ) , .ZN( u0_u4_u6_n173 ) );
  INV_X1 u0_u4_u6_U21 (.A( u0_u4_u6_n121 ) , .ZN( u0_u4_u6_n167 ) );
  INV_X1 u0_u4_u6_U22 (.A( u0_u4_u6_n100 ) , .ZN( u0_u4_u6_n169 ) );
  INV_X1 u0_u4_u6_U23 (.A( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n170 ) );
  INV_X1 u0_u4_u6_U24 (.A( u0_u4_u6_n113 ) , .ZN( u0_u4_u6_n168 ) );
  AND2_X1 u0_u4_u6_U25 (.A1( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n119 ) , .ZN( u0_u4_u6_n133 ) );
  AND2_X1 u0_u4_u6_U26 (.A2( u0_u4_u6_n121 ) , .A1( u0_u4_u6_n122 ) , .ZN( u0_u4_u6_n131 ) );
  AND3_X1 u0_u4_u6_U27 (.ZN( u0_u4_u6_n120 ) , .A2( u0_u4_u6_n127 ) , .A1( u0_u4_u6_n132 ) , .A3( u0_u4_u6_n145 ) );
  INV_X1 u0_u4_u6_U28 (.A( u0_u4_u6_n146 ) , .ZN( u0_u4_u6_n163 ) );
  AOI222_X1 u0_u4_u6_U29 (.ZN( u0_u4_u6_n114 ) , .A1( u0_u4_u6_n118 ) , .A2( u0_u4_u6_n126 ) , .B2( u0_u4_u6_n151 ) , .C2( u0_u4_u6_n159 ) , .C1( u0_u4_u6_n168 ) , .B1( u0_u4_u6_n169 ) );
  INV_X1 u0_u4_u6_U3 (.A( u0_u4_u6_n110 ) , .ZN( u0_u4_u6_n166 ) );
  NOR2_X1 u0_u4_u6_U30 (.A1( u0_u4_u6_n162 ) , .A2( u0_u4_u6_n165 ) , .ZN( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U31 (.A1( u0_u4_u6_n144 ) , .ZN( u0_u4_u6_n151 ) , .A2( u0_u4_u6_n158 ) );
  NAND2_X1 u0_u4_u6_U32 (.ZN( u0_u4_u6_n132 ) , .A1( u0_u4_u6_n91 ) , .A2( u0_u4_u6_n97 ) );
  AOI22_X1 u0_u4_u6_U33 (.B2( u0_u4_u6_n110 ) , .B1( u0_u4_u6_n111 ) , .A1( u0_u4_u6_n112 ) , .ZN( u0_u4_u6_n115 ) , .A2( u0_u4_u6_n161 ) );
  NAND4_X1 u0_u4_u6_U34 (.A3( u0_u4_u6_n109 ) , .ZN( u0_u4_u6_n112 ) , .A4( u0_u4_u6_n132 ) , .A2( u0_u4_u6_n147 ) , .A1( u0_u4_u6_n166 ) );
  NOR2_X1 u0_u4_u6_U35 (.ZN( u0_u4_u6_n109 ) , .A1( u0_u4_u6_n170 ) , .A2( u0_u4_u6_n173 ) );
  NOR2_X1 u0_u4_u6_U36 (.A2( u0_u4_u6_n126 ) , .ZN( u0_u4_u6_n155 ) , .A1( u0_u4_u6_n160 ) );
  NAND2_X1 u0_u4_u6_U37 (.ZN( u0_u4_u6_n146 ) , .A2( u0_u4_u6_n94 ) , .A1( u0_u4_u6_n99 ) );
  AOI21_X1 u0_u4_u6_U38 (.A( u0_u4_u6_n144 ) , .B2( u0_u4_u6_n145 ) , .B1( u0_u4_u6_n146 ) , .ZN( u0_u4_u6_n150 ) );
  AOI211_X1 u0_u4_u6_U39 (.B( u0_u4_u6_n134 ) , .A( u0_u4_u6_n135 ) , .C1( u0_u4_u6_n136 ) , .ZN( u0_u4_u6_n137 ) , .C2( u0_u4_u6_n151 ) );
  INV_X1 u0_u4_u6_U4 (.A( u0_u4_u6_n142 ) , .ZN( u0_u4_u6_n174 ) );
  NAND4_X1 u0_u4_u6_U40 (.A4( u0_u4_u6_n127 ) , .A3( u0_u4_u6_n128 ) , .A2( u0_u4_u6_n129 ) , .A1( u0_u4_u6_n130 ) , .ZN( u0_u4_u6_n136 ) );
  AOI21_X1 u0_u4_u6_U41 (.B2( u0_u4_u6_n132 ) , .B1( u0_u4_u6_n133 ) , .ZN( u0_u4_u6_n134 ) , .A( u0_u4_u6_n158 ) );
  AOI21_X1 u0_u4_u6_U42 (.B1( u0_u4_u6_n131 ) , .ZN( u0_u4_u6_n135 ) , .A( u0_u4_u6_n144 ) , .B2( u0_u4_u6_n146 ) );
  INV_X1 u0_u4_u6_U43 (.A( u0_u4_u6_n111 ) , .ZN( u0_u4_u6_n158 ) );
  NAND2_X1 u0_u4_u6_U44 (.ZN( u0_u4_u6_n127 ) , .A1( u0_u4_u6_n91 ) , .A2( u0_u4_u6_n92 ) );
  NAND2_X1 u0_u4_u6_U45 (.ZN( u0_u4_u6_n129 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n96 ) );
  INV_X1 u0_u4_u6_U46 (.A( u0_u4_u6_n144 ) , .ZN( u0_u4_u6_n159 ) );
  NAND2_X1 u0_u4_u6_U47 (.ZN( u0_u4_u6_n145 ) , .A2( u0_u4_u6_n97 ) , .A1( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U48 (.ZN( u0_u4_u6_n148 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n94 ) );
  NAND2_X1 u0_u4_u6_U49 (.ZN( u0_u4_u6_n108 ) , .A2( u0_u4_u6_n139 ) , .A1( u0_u4_u6_n144 ) );
  NAND2_X1 u0_u4_u6_U5 (.A2( u0_u4_u6_n143 ) , .ZN( u0_u4_u6_n152 ) , .A1( u0_u4_u6_n166 ) );
  NAND2_X1 u0_u4_u6_U50 (.ZN( u0_u4_u6_n121 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n97 ) );
  NAND2_X1 u0_u4_u6_U51 (.ZN( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n95 ) );
  AND2_X1 u0_u4_u6_U52 (.ZN( u0_u4_u6_n118 ) , .A2( u0_u4_u6_n91 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U53 (.ZN( u0_u4_u6_n147 ) , .A2( u0_u4_u6_n98 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U54 (.ZN( u0_u4_u6_n128 ) , .A1( u0_u4_u6_n94 ) , .A2( u0_u4_u6_n96 ) );
  NAND2_X1 u0_u4_u6_U55 (.ZN( u0_u4_u6_n119 ) , .A2( u0_u4_u6_n95 ) , .A1( u0_u4_u6_n99 ) );
  NAND2_X1 u0_u4_u6_U56 (.ZN( u0_u4_u6_n123 ) , .A2( u0_u4_u6_n91 ) , .A1( u0_u4_u6_n96 ) );
  NAND2_X1 u0_u4_u6_U57 (.ZN( u0_u4_u6_n100 ) , .A2( u0_u4_u6_n92 ) , .A1( u0_u4_u6_n98 ) );
  NAND2_X1 u0_u4_u6_U58 (.ZN( u0_u4_u6_n122 ) , .A1( u0_u4_u6_n94 ) , .A2( u0_u4_u6_n97 ) );
  INV_X1 u0_u4_u6_U59 (.A( u0_u4_u6_n139 ) , .ZN( u0_u4_u6_n160 ) );
  AOI22_X1 u0_u4_u6_U6 (.B2( u0_u4_u6_n101 ) , .A1( u0_u4_u6_n102 ) , .ZN( u0_u4_u6_n103 ) , .B1( u0_u4_u6_n160 ) , .A2( u0_u4_u6_n161 ) );
  NAND2_X1 u0_u4_u6_U60 (.ZN( u0_u4_u6_n113 ) , .A1( u0_u4_u6_n96 ) , .A2( u0_u4_u6_n98 ) );
  NOR2_X1 u0_u4_u6_U61 (.A2( u0_u4_X_40 ) , .A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n126 ) );
  NOR2_X1 u0_u4_u6_U62 (.A2( u0_u4_X_39 ) , .A1( u0_u4_X_42 ) , .ZN( u0_u4_u6_n92 ) );
  NOR2_X1 u0_u4_u6_U63 (.A2( u0_u4_X_39 ) , .A1( u0_u4_u6_n156 ) , .ZN( u0_u4_u6_n97 ) );
  NOR2_X1 u0_u4_u6_U64 (.A2( u0_u4_X_38 ) , .A1( u0_u4_u6_n165 ) , .ZN( u0_u4_u6_n95 ) );
  NOR2_X1 u0_u4_u6_U65 (.A2( u0_u4_X_41 ) , .ZN( u0_u4_u6_n111 ) , .A1( u0_u4_u6_n157 ) );
  NOR2_X1 u0_u4_u6_U66 (.A2( u0_u4_X_37 ) , .A1( u0_u4_u6_n162 ) , .ZN( u0_u4_u6_n94 ) );
  NOR2_X1 u0_u4_u6_U67 (.A2( u0_u4_X_37 ) , .A1( u0_u4_X_38 ) , .ZN( u0_u4_u6_n91 ) );
  NAND2_X1 u0_u4_u6_U68 (.A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n144 ) , .A2( u0_u4_u6_n157 ) );
  NAND2_X1 u0_u4_u6_U69 (.A2( u0_u4_X_40 ) , .A1( u0_u4_X_41 ) , .ZN( u0_u4_u6_n139 ) );
  NOR2_X1 u0_u4_u6_U7 (.A1( u0_u4_u6_n118 ) , .ZN( u0_u4_u6_n143 ) , .A2( u0_u4_u6_n168 ) );
  AND2_X1 u0_u4_u6_U70 (.A1( u0_u4_X_39 ) , .A2( u0_u4_u6_n156 ) , .ZN( u0_u4_u6_n96 ) );
  AND2_X1 u0_u4_u6_U71 (.A1( u0_u4_X_39 ) , .A2( u0_u4_X_42 ) , .ZN( u0_u4_u6_n99 ) );
  INV_X1 u0_u4_u6_U72 (.A( u0_u4_X_40 ) , .ZN( u0_u4_u6_n157 ) );
  INV_X1 u0_u4_u6_U73 (.A( u0_u4_X_37 ) , .ZN( u0_u4_u6_n165 ) );
  INV_X1 u0_u4_u6_U74 (.A( u0_u4_X_38 ) , .ZN( u0_u4_u6_n162 ) );
  INV_X1 u0_u4_u6_U75 (.A( u0_u4_X_42 ) , .ZN( u0_u4_u6_n156 ) );
  NAND4_X1 u0_u4_u6_U76 (.ZN( u0_out4_32 ) , .A4( u0_u4_u6_n103 ) , .A3( u0_u4_u6_n104 ) , .A2( u0_u4_u6_n105 ) , .A1( u0_u4_u6_n106 ) );
  AOI22_X1 u0_u4_u6_U77 (.ZN( u0_u4_u6_n105 ) , .A2( u0_u4_u6_n108 ) , .A1( u0_u4_u6_n118 ) , .B2( u0_u4_u6_n126 ) , .B1( u0_u4_u6_n171 ) );
  AOI22_X1 u0_u4_u6_U78 (.ZN( u0_u4_u6_n104 ) , .A1( u0_u4_u6_n111 ) , .B1( u0_u4_u6_n124 ) , .B2( u0_u4_u6_n151 ) , .A2( u0_u4_u6_n93 ) );
  NAND4_X1 u0_u4_u6_U79 (.ZN( u0_out4_12 ) , .A4( u0_u4_u6_n114 ) , .A3( u0_u4_u6_n115 ) , .A2( u0_u4_u6_n116 ) , .A1( u0_u4_u6_n117 ) );
  INV_X1 u0_u4_u6_U8 (.ZN( u0_u4_u6_n172 ) , .A( u0_u4_u6_n88 ) );
  OAI22_X1 u0_u4_u6_U80 (.B2( u0_u4_u6_n111 ) , .ZN( u0_u4_u6_n116 ) , .B1( u0_u4_u6_n126 ) , .A2( u0_u4_u6_n164 ) , .A1( u0_u4_u6_n167 ) );
  OAI21_X1 u0_u4_u6_U81 (.A( u0_u4_u6_n108 ) , .ZN( u0_u4_u6_n117 ) , .B2( u0_u4_u6_n141 ) , .B1( u0_u4_u6_n163 ) );
  OAI211_X1 u0_u4_u6_U82 (.ZN( u0_out4_22 ) , .B( u0_u4_u6_n137 ) , .A( u0_u4_u6_n138 ) , .C2( u0_u4_u6_n139 ) , .C1( u0_u4_u6_n140 ) );
  AOI22_X1 u0_u4_u6_U83 (.B1( u0_u4_u6_n124 ) , .A2( u0_u4_u6_n125 ) , .A1( u0_u4_u6_n126 ) , .ZN( u0_u4_u6_n138 ) , .B2( u0_u4_u6_n161 ) );
  AND4_X1 u0_u4_u6_U84 (.A3( u0_u4_u6_n119 ) , .A1( u0_u4_u6_n120 ) , .A4( u0_u4_u6_n129 ) , .ZN( u0_u4_u6_n140 ) , .A2( u0_u4_u6_n143 ) );
  OAI211_X1 u0_u4_u6_U85 (.ZN( u0_out4_7 ) , .B( u0_u4_u6_n153 ) , .C2( u0_u4_u6_n154 ) , .C1( u0_u4_u6_n155 ) , .A( u0_u4_u6_n174 ) );
  NOR3_X1 u0_u4_u6_U86 (.A1( u0_u4_u6_n141 ) , .ZN( u0_u4_u6_n154 ) , .A3( u0_u4_u6_n164 ) , .A2( u0_u4_u6_n171 ) );
  AOI211_X1 u0_u4_u6_U87 (.B( u0_u4_u6_n149 ) , .A( u0_u4_u6_n150 ) , .C2( u0_u4_u6_n151 ) , .C1( u0_u4_u6_n152 ) , .ZN( u0_u4_u6_n153 ) );
  NAND3_X1 u0_u4_u6_U88 (.A2( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n125 ) , .A1( u0_u4_u6_n130 ) , .A3( u0_u4_u6_n131 ) );
  NAND3_X1 u0_u4_u6_U89 (.A3( u0_u4_u6_n133 ) , .ZN( u0_u4_u6_n141 ) , .A1( u0_u4_u6_n145 ) , .A2( u0_u4_u6_n148 ) );
  OAI21_X1 u0_u4_u6_U9 (.A( u0_u4_u6_n159 ) , .B1( u0_u4_u6_n169 ) , .B2( u0_u4_u6_n173 ) , .ZN( u0_u4_u6_n90 ) );
  NAND3_X1 u0_u4_u6_U90 (.ZN( u0_u4_u6_n101 ) , .A3( u0_u4_u6_n107 ) , .A2( u0_u4_u6_n121 ) , .A1( u0_u4_u6_n127 ) );
  NAND3_X1 u0_u4_u6_U91 (.ZN( u0_u4_u6_n102 ) , .A3( u0_u4_u6_n130 ) , .A2( u0_u4_u6_n145 ) , .A1( u0_u4_u6_n166 ) );
  NAND3_X1 u0_u4_u6_U92 (.A3( u0_u4_u6_n113 ) , .A1( u0_u4_u6_n119 ) , .A2( u0_u4_u6_n123 ) , .ZN( u0_u4_u6_n93 ) );
  NAND3_X1 u0_u4_u6_U93 (.ZN( u0_u4_u6_n142 ) , .A2( u0_u4_u6_n172 ) , .A3( u0_u4_u6_n89 ) , .A1( u0_u4_u6_n90 ) );
  XOR2_X1 u0_u5_U1 (.B( u0_K6_9 ) , .A( u0_R4_6 ) , .Z( u0_u5_X_9 ) );
  XOR2_X1 u0_u5_U16 (.B( u0_K6_3 ) , .A( u0_R4_2 ) , .Z( u0_u5_X_3 ) );
  XOR2_X1 u0_u5_U22 (.B( u0_K6_34 ) , .A( u0_R4_23 ) , .Z( u0_u5_X_34 ) );
  XOR2_X1 u0_u5_U30 (.B( u0_K6_27 ) , .A( u0_R4_18 ) , .Z( u0_u5_X_27 ) );
  XOR2_X1 u0_u5_U35 (.B( u0_K6_22 ) , .A( u0_R4_15 ) , .Z( u0_u5_X_22 ) );
  XOR2_X1 u0_u5_U36 (.B( u0_K6_21 ) , .A( u0_R4_14 ) , .Z( u0_u5_X_21 ) );
  XOR2_X1 u0_u5_U42 (.B( u0_K6_16 ) , .A( u0_R4_11 ) , .Z( u0_u5_X_16 ) );
  XOR2_X1 u0_u5_U43 (.B( u0_K6_15 ) , .A( u0_R4_10 ) , .Z( u0_u5_X_15 ) );
  XOR2_X1 u0_u5_U48 (.B( u0_K6_10 ) , .A( u0_R4_7 ) , .Z( u0_u5_X_10 ) );
  XOR2_X1 u0_u5_U9 (.B( u0_K6_46 ) , .A( u0_R4_31 ) , .Z( u0_u5_X_46 ) );
  XOR2_X1 u0_u6_U1 (.B( u0_K7_9 ) , .A( u0_R5_6 ) , .Z( u0_u6_X_9 ) );
  XOR2_X1 u0_u6_U10 (.B( u0_K7_45 ) , .A( u0_R5_30 ) , .Z( u0_u6_X_45 ) );
  XOR2_X1 u0_u6_U11 (.B( u0_K7_44 ) , .A( u0_R5_29 ) , .Z( u0_u6_X_44 ) );
  XOR2_X1 u0_u6_U12 (.B( u0_K7_43 ) , .A( u0_R5_28 ) , .Z( u0_u6_X_43 ) );
  XOR2_X1 u0_u6_U13 (.B( u0_K7_42 ) , .A( u0_R5_29 ) , .Z( u0_u6_X_42 ) );
  XOR2_X1 u0_u6_U14 (.B( u0_K7_41 ) , .A( u0_R5_28 ) , .Z( u0_u6_X_41 ) );
  XOR2_X1 u0_u6_U15 (.B( u0_K7_40 ) , .A( u0_R5_27 ) , .Z( u0_u6_X_40 ) );
  XOR2_X1 u0_u6_U17 (.B( u0_K7_39 ) , .A( u0_R5_26 ) , .Z( u0_u6_X_39 ) );
  XOR2_X1 u0_u6_U18 (.B( u0_K7_38 ) , .A( u0_R5_25 ) , .Z( u0_u6_X_38 ) );
  XOR2_X1 u0_u6_U19 (.B( u0_K7_37 ) , .A( u0_R5_24 ) , .Z( u0_u6_X_37 ) );
  XOR2_X1 u0_u6_U21 (.B( u0_K7_35 ) , .A( u0_R5_24 ) , .Z( u0_u6_X_35 ) );
  XOR2_X1 u0_u6_U22 (.B( u0_K7_34 ) , .A( u0_R5_23 ) , .Z( u0_u6_X_34 ) );
  XOR2_X1 u0_u6_U23 (.B( u0_K7_33 ) , .A( u0_R5_22 ) , .Z( u0_u6_X_33 ) );
  XOR2_X1 u0_u6_U24 (.B( u0_K7_32 ) , .A( u0_R5_21 ) , .Z( u0_u6_X_32 ) );
  XOR2_X1 u0_u6_U25 (.B( u0_K7_31 ) , .A( u0_R5_20 ) , .Z( u0_u6_X_31 ) );
  XOR2_X1 u0_u6_U26 (.B( u0_K7_30 ) , .A( u0_R5_21 ) , .Z( u0_u6_X_30 ) );
  XOR2_X1 u0_u6_U27 (.B( u0_K7_2 ) , .A( u0_R5_1 ) , .Z( u0_u6_X_2 ) );
  XOR2_X1 u0_u6_U28 (.B( u0_K7_29 ) , .A( u0_R5_20 ) , .Z( u0_u6_X_29 ) );
  XOR2_X1 u0_u6_U29 (.B( u0_K7_28 ) , .A( u0_R5_19 ) , .Z( u0_u6_X_28 ) );
  XOR2_X1 u0_u6_U30 (.B( u0_K7_27 ) , .A( u0_R5_18 ) , .Z( u0_u6_X_27 ) );
  XOR2_X1 u0_u6_U31 (.B( u0_K7_26 ) , .A( u0_R5_17 ) , .Z( u0_u6_X_26 ) );
  XOR2_X1 u0_u6_U32 (.B( u0_K7_25 ) , .A( u0_R5_16 ) , .Z( u0_u6_X_25 ) );
  XOR2_X1 u0_u6_U33 (.B( u0_K7_24 ) , .A( u0_R5_17 ) , .Z( u0_u6_X_24 ) );
  XOR2_X1 u0_u6_U34 (.B( u0_K7_23 ) , .A( u0_R5_16 ) , .Z( u0_u6_X_23 ) );
  XOR2_X1 u0_u6_U35 (.B( u0_K7_22 ) , .A( u0_R5_15 ) , .Z( u0_u6_X_22 ) );
  XOR2_X1 u0_u6_U36 (.B( u0_K7_21 ) , .A( u0_R5_14 ) , .Z( u0_u6_X_21 ) );
  XOR2_X1 u0_u6_U42 (.B( u0_K7_16 ) , .A( u0_R5_11 ) , .Z( u0_u6_X_16 ) );
  XOR2_X1 u0_u6_U43 (.B( u0_K7_15 ) , .A( u0_R5_10 ) , .Z( u0_u6_X_15 ) );
  XOR2_X1 u0_u6_U7 (.B( u0_K7_48 ) , .A( u0_R5_1 ) , .Z( u0_u6_X_48 ) );
  XOR2_X1 u0_u6_U8 (.B( u0_K7_47 ) , .A( u0_R5_32 ) , .Z( u0_u6_X_47 ) );
  XOR2_X1 u0_u6_U9 (.B( u0_K7_46 ) , .A( u0_R5_31 ) , .Z( u0_u6_X_46 ) );
  OAI22_X1 u0_u6_u4_U10 (.B2( u0_u6_u4_n135 ) , .ZN( u0_u6_u4_n137 ) , .B1( u0_u6_u4_n153 ) , .A1( u0_u6_u4_n155 ) , .A2( u0_u6_u4_n171 ) );
  AND3_X1 u0_u6_u4_U11 (.A2( u0_u6_u4_n134 ) , .ZN( u0_u6_u4_n135 ) , .A3( u0_u6_u4_n145 ) , .A1( u0_u6_u4_n157 ) );
  NAND2_X1 u0_u6_u4_U12 (.ZN( u0_u6_u4_n132 ) , .A2( u0_u6_u4_n170 ) , .A1( u0_u6_u4_n173 ) );
  AOI21_X1 u0_u6_u4_U13 (.B2( u0_u6_u4_n160 ) , .B1( u0_u6_u4_n161 ) , .ZN( u0_u6_u4_n162 ) , .A( u0_u6_u4_n170 ) );
  AOI21_X1 u0_u6_u4_U14 (.ZN( u0_u6_u4_n107 ) , .B2( u0_u6_u4_n143 ) , .A( u0_u6_u4_n174 ) , .B1( u0_u6_u4_n184 ) );
  AOI21_X1 u0_u6_u4_U15 (.B2( u0_u6_u4_n158 ) , .B1( u0_u6_u4_n159 ) , .ZN( u0_u6_u4_n163 ) , .A( u0_u6_u4_n174 ) );
  AOI21_X1 u0_u6_u4_U16 (.A( u0_u6_u4_n153 ) , .B2( u0_u6_u4_n154 ) , .B1( u0_u6_u4_n155 ) , .ZN( u0_u6_u4_n165 ) );
  AOI21_X1 u0_u6_u4_U17 (.A( u0_u6_u4_n156 ) , .B2( u0_u6_u4_n157 ) , .ZN( u0_u6_u4_n164 ) , .B1( u0_u6_u4_n184 ) );
  INV_X1 u0_u6_u4_U18 (.A( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n170 ) );
  AND2_X1 u0_u6_u4_U19 (.A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n155 ) , .A1( u0_u6_u4_n160 ) );
  INV_X1 u0_u6_u4_U20 (.A( u0_u6_u4_n156 ) , .ZN( u0_u6_u4_n175 ) );
  NAND2_X1 u0_u6_u4_U21 (.A2( u0_u6_u4_n118 ) , .ZN( u0_u6_u4_n131 ) , .A1( u0_u6_u4_n147 ) );
  NAND2_X1 u0_u6_u4_U22 (.A1( u0_u6_u4_n119 ) , .A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n130 ) );
  NAND2_X1 u0_u6_u4_U23 (.ZN( u0_u6_u4_n117 ) , .A2( u0_u6_u4_n118 ) , .A1( u0_u6_u4_n148 ) );
  NAND2_X1 u0_u6_u4_U24 (.ZN( u0_u6_u4_n129 ) , .A1( u0_u6_u4_n134 ) , .A2( u0_u6_u4_n148 ) );
  AND3_X1 u0_u6_u4_U25 (.A1( u0_u6_u4_n119 ) , .A2( u0_u6_u4_n143 ) , .A3( u0_u6_u4_n154 ) , .ZN( u0_u6_u4_n161 ) );
  AND2_X1 u0_u6_u4_U26 (.A1( u0_u6_u4_n145 ) , .A2( u0_u6_u4_n147 ) , .ZN( u0_u6_u4_n159 ) );
  OR3_X1 u0_u6_u4_U27 (.A3( u0_u6_u4_n114 ) , .A2( u0_u6_u4_n115 ) , .A1( u0_u6_u4_n116 ) , .ZN( u0_u6_u4_n136 ) );
  AOI21_X1 u0_u6_u4_U28 (.A( u0_u6_u4_n113 ) , .ZN( u0_u6_u4_n116 ) , .B2( u0_u6_u4_n173 ) , .B1( u0_u6_u4_n174 ) );
  AOI21_X1 u0_u6_u4_U29 (.ZN( u0_u6_u4_n115 ) , .B2( u0_u6_u4_n145 ) , .B1( u0_u6_u4_n146 ) , .A( u0_u6_u4_n156 ) );
  NOR2_X1 u0_u6_u4_U3 (.ZN( u0_u6_u4_n121 ) , .A1( u0_u6_u4_n181 ) , .A2( u0_u6_u4_n182 ) );
  OAI22_X1 u0_u6_u4_U30 (.ZN( u0_u6_u4_n114 ) , .A2( u0_u6_u4_n121 ) , .B1( u0_u6_u4_n160 ) , .B2( u0_u6_u4_n170 ) , .A1( u0_u6_u4_n171 ) );
  INV_X1 u0_u6_u4_U31 (.A( u0_u6_u4_n158 ) , .ZN( u0_u6_u4_n182 ) );
  INV_X1 u0_u6_u4_U32 (.ZN( u0_u6_u4_n181 ) , .A( u0_u6_u4_n96 ) );
  INV_X1 u0_u6_u4_U33 (.A( u0_u6_u4_n144 ) , .ZN( u0_u6_u4_n179 ) );
  INV_X1 u0_u6_u4_U34 (.A( u0_u6_u4_n157 ) , .ZN( u0_u6_u4_n178 ) );
  NAND2_X1 u0_u6_u4_U35 (.A2( u0_u6_u4_n154 ) , .A1( u0_u6_u4_n96 ) , .ZN( u0_u6_u4_n97 ) );
  INV_X1 u0_u6_u4_U36 (.ZN( u0_u6_u4_n186 ) , .A( u0_u6_u4_n95 ) );
  OAI221_X1 u0_u6_u4_U37 (.C1( u0_u6_u4_n134 ) , .B1( u0_u6_u4_n158 ) , .B2( u0_u6_u4_n171 ) , .C2( u0_u6_u4_n173 ) , .A( u0_u6_u4_n94 ) , .ZN( u0_u6_u4_n95 ) );
  AOI222_X1 u0_u6_u4_U38 (.B2( u0_u6_u4_n132 ) , .A1( u0_u6_u4_n138 ) , .C2( u0_u6_u4_n175 ) , .A2( u0_u6_u4_n179 ) , .C1( u0_u6_u4_n181 ) , .B1( u0_u6_u4_n185 ) , .ZN( u0_u6_u4_n94 ) );
  INV_X1 u0_u6_u4_U39 (.A( u0_u6_u4_n113 ) , .ZN( u0_u6_u4_n185 ) );
  INV_X1 u0_u6_u4_U4 (.A( u0_u6_u4_n117 ) , .ZN( u0_u6_u4_n184 ) );
  INV_X1 u0_u6_u4_U40 (.A( u0_u6_u4_n143 ) , .ZN( u0_u6_u4_n183 ) );
  NOR2_X1 u0_u6_u4_U41 (.ZN( u0_u6_u4_n138 ) , .A1( u0_u6_u4_n168 ) , .A2( u0_u6_u4_n169 ) );
  NOR2_X1 u0_u6_u4_U42 (.A1( u0_u6_u4_n150 ) , .A2( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n153 ) );
  NOR2_X1 u0_u6_u4_U43 (.A2( u0_u6_u4_n128 ) , .A1( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n156 ) );
  AOI22_X1 u0_u6_u4_U44 (.B2( u0_u6_u4_n122 ) , .A1( u0_u6_u4_n123 ) , .ZN( u0_u6_u4_n124 ) , .B1( u0_u6_u4_n128 ) , .A2( u0_u6_u4_n172 ) );
  INV_X1 u0_u6_u4_U45 (.A( u0_u6_u4_n153 ) , .ZN( u0_u6_u4_n172 ) );
  NAND2_X1 u0_u6_u4_U46 (.A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n123 ) , .A1( u0_u6_u4_n161 ) );
  AOI22_X1 u0_u6_u4_U47 (.B2( u0_u6_u4_n132 ) , .A2( u0_u6_u4_n133 ) , .ZN( u0_u6_u4_n140 ) , .A1( u0_u6_u4_n150 ) , .B1( u0_u6_u4_n179 ) );
  NAND2_X1 u0_u6_u4_U48 (.ZN( u0_u6_u4_n133 ) , .A2( u0_u6_u4_n146 ) , .A1( u0_u6_u4_n154 ) );
  NAND2_X1 u0_u6_u4_U49 (.A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n154 ) , .A2( u0_u6_u4_n98 ) );
  NOR4_X1 u0_u6_u4_U5 (.A4( u0_u6_u4_n106 ) , .A3( u0_u6_u4_n107 ) , .A2( u0_u6_u4_n108 ) , .A1( u0_u6_u4_n109 ) , .ZN( u0_u6_u4_n110 ) );
  NAND2_X1 u0_u6_u4_U50 (.A1( u0_u6_u4_n101 ) , .ZN( u0_u6_u4_n158 ) , .A2( u0_u6_u4_n99 ) );
  AOI21_X1 u0_u6_u4_U51 (.ZN( u0_u6_u4_n127 ) , .A( u0_u6_u4_n136 ) , .B2( u0_u6_u4_n150 ) , .B1( u0_u6_u4_n180 ) );
  INV_X1 u0_u6_u4_U52 (.A( u0_u6_u4_n160 ) , .ZN( u0_u6_u4_n180 ) );
  NAND2_X1 u0_u6_u4_U53 (.A2( u0_u6_u4_n104 ) , .A1( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n146 ) );
  NAND2_X1 u0_u6_u4_U54 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n160 ) );
  NAND2_X1 u0_u6_u4_U55 (.ZN( u0_u6_u4_n134 ) , .A1( u0_u6_u4_n98 ) , .A2( u0_u6_u4_n99 ) );
  NAND2_X1 u0_u6_u4_U56 (.A1( u0_u6_u4_n103 ) , .A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n143 ) );
  NAND2_X1 u0_u6_u4_U57 (.A2( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n145 ) , .A1( u0_u6_u4_n98 ) );
  NAND2_X1 u0_u6_u4_U58 (.A1( u0_u6_u4_n100 ) , .A2( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n120 ) );
  NAND2_X1 u0_u6_u4_U59 (.A1( u0_u6_u4_n102 ) , .A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n148 ) );
  AOI21_X1 u0_u6_u4_U6 (.ZN( u0_u6_u4_n106 ) , .B2( u0_u6_u4_n146 ) , .B1( u0_u6_u4_n158 ) , .A( u0_u6_u4_n170 ) );
  NAND2_X1 u0_u6_u4_U60 (.A2( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n157 ) );
  INV_X1 u0_u6_u4_U61 (.A( u0_u6_u4_n150 ) , .ZN( u0_u6_u4_n173 ) );
  INV_X1 u0_u6_u4_U62 (.A( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n171 ) );
  NAND2_X1 u0_u6_u4_U63 (.A1( u0_u6_u4_n100 ) , .ZN( u0_u6_u4_n118 ) , .A2( u0_u6_u4_n99 ) );
  NAND2_X1 u0_u6_u4_U64 (.A2( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n144 ) );
  NAND2_X1 u0_u6_u4_U65 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n96 ) );
  INV_X1 u0_u6_u4_U66 (.A( u0_u6_u4_n128 ) , .ZN( u0_u6_u4_n174 ) );
  NAND2_X1 u0_u6_u4_U67 (.A2( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n119 ) , .A1( u0_u6_u4_n98 ) );
  NAND2_X1 u0_u6_u4_U68 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n147 ) );
  NAND2_X1 u0_u6_u4_U69 (.A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n113 ) , .A1( u0_u6_u4_n99 ) );
  AOI21_X1 u0_u6_u4_U7 (.ZN( u0_u6_u4_n108 ) , .B2( u0_u6_u4_n134 ) , .B1( u0_u6_u4_n155 ) , .A( u0_u6_u4_n156 ) );
  NOR2_X1 u0_u6_u4_U70 (.A2( u0_u6_X_28 ) , .ZN( u0_u6_u4_n150 ) , .A1( u0_u6_u4_n168 ) );
  NOR2_X1 u0_u6_u4_U71 (.A2( u0_u6_X_29 ) , .ZN( u0_u6_u4_n152 ) , .A1( u0_u6_u4_n169 ) );
  NOR2_X1 u0_u6_u4_U72 (.A2( u0_u6_X_30 ) , .ZN( u0_u6_u4_n105 ) , .A1( u0_u6_u4_n176 ) );
  NOR2_X1 u0_u6_u4_U73 (.A2( u0_u6_X_26 ) , .ZN( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n177 ) );
  NOR2_X1 u0_u6_u4_U74 (.A2( u0_u6_X_28 ) , .A1( u0_u6_X_29 ) , .ZN( u0_u6_u4_n128 ) );
  NOR2_X1 u0_u6_u4_U75 (.A2( u0_u6_X_27 ) , .A1( u0_u6_X_30 ) , .ZN( u0_u6_u4_n102 ) );
  NOR2_X1 u0_u6_u4_U76 (.A2( u0_u6_X_25 ) , .A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n98 ) );
  AND2_X1 u0_u6_u4_U77 (.A2( u0_u6_X_25 ) , .A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n104 ) );
  AND2_X1 u0_u6_u4_U78 (.A1( u0_u6_X_30 ) , .A2( u0_u6_u4_n176 ) , .ZN( u0_u6_u4_n99 ) );
  AND2_X1 u0_u6_u4_U79 (.A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n101 ) , .A2( u0_u6_u4_n177 ) );
  AOI21_X1 u0_u6_u4_U8 (.ZN( u0_u6_u4_n109 ) , .A( u0_u6_u4_n153 ) , .B1( u0_u6_u4_n159 ) , .B2( u0_u6_u4_n184 ) );
  AND2_X1 u0_u6_u4_U80 (.A1( u0_u6_X_27 ) , .A2( u0_u6_X_30 ) , .ZN( u0_u6_u4_n103 ) );
  INV_X1 u0_u6_u4_U81 (.A( u0_u6_X_28 ) , .ZN( u0_u6_u4_n169 ) );
  INV_X1 u0_u6_u4_U82 (.A( u0_u6_X_29 ) , .ZN( u0_u6_u4_n168 ) );
  INV_X1 u0_u6_u4_U83 (.A( u0_u6_X_25 ) , .ZN( u0_u6_u4_n177 ) );
  INV_X1 u0_u6_u4_U84 (.A( u0_u6_X_27 ) , .ZN( u0_u6_u4_n176 ) );
  NAND4_X1 u0_u6_u4_U85 (.ZN( u0_out6_25 ) , .A4( u0_u6_u4_n139 ) , .A3( u0_u6_u4_n140 ) , .A2( u0_u6_u4_n141 ) , .A1( u0_u6_u4_n142 ) );
  OAI21_X1 u0_u6_u4_U86 (.B2( u0_u6_u4_n131 ) , .ZN( u0_u6_u4_n141 ) , .A( u0_u6_u4_n175 ) , .B1( u0_u6_u4_n183 ) );
  OAI21_X1 u0_u6_u4_U87 (.A( u0_u6_u4_n128 ) , .B2( u0_u6_u4_n129 ) , .B1( u0_u6_u4_n130 ) , .ZN( u0_u6_u4_n142 ) );
  NAND4_X1 u0_u6_u4_U88 (.ZN( u0_out6_14 ) , .A4( u0_u6_u4_n124 ) , .A3( u0_u6_u4_n125 ) , .A2( u0_u6_u4_n126 ) , .A1( u0_u6_u4_n127 ) );
  AOI22_X1 u0_u6_u4_U89 (.B2( u0_u6_u4_n117 ) , .ZN( u0_u6_u4_n126 ) , .A1( u0_u6_u4_n129 ) , .B1( u0_u6_u4_n152 ) , .A2( u0_u6_u4_n175 ) );
  AOI211_X1 u0_u6_u4_U9 (.B( u0_u6_u4_n136 ) , .A( u0_u6_u4_n137 ) , .C2( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n139 ) , .C1( u0_u6_u4_n182 ) );
  AOI22_X1 u0_u6_u4_U90 (.ZN( u0_u6_u4_n125 ) , .B2( u0_u6_u4_n131 ) , .A2( u0_u6_u4_n132 ) , .B1( u0_u6_u4_n138 ) , .A1( u0_u6_u4_n178 ) );
  NAND4_X1 u0_u6_u4_U91 (.ZN( u0_out6_8 ) , .A4( u0_u6_u4_n110 ) , .A3( u0_u6_u4_n111 ) , .A2( u0_u6_u4_n112 ) , .A1( u0_u6_u4_n186 ) );
  NAND2_X1 u0_u6_u4_U92 (.ZN( u0_u6_u4_n112 ) , .A2( u0_u6_u4_n130 ) , .A1( u0_u6_u4_n150 ) );
  AOI22_X1 u0_u6_u4_U93 (.ZN( u0_u6_u4_n111 ) , .B2( u0_u6_u4_n132 ) , .A1( u0_u6_u4_n152 ) , .B1( u0_u6_u4_n178 ) , .A2( u0_u6_u4_n97 ) );
  AOI22_X1 u0_u6_u4_U94 (.B2( u0_u6_u4_n149 ) , .B1( u0_u6_u4_n150 ) , .A2( u0_u6_u4_n151 ) , .A1( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n167 ) );
  NOR4_X1 u0_u6_u4_U95 (.A4( u0_u6_u4_n162 ) , .A3( u0_u6_u4_n163 ) , .A2( u0_u6_u4_n164 ) , .A1( u0_u6_u4_n165 ) , .ZN( u0_u6_u4_n166 ) );
  NAND3_X1 u0_u6_u4_U96 (.ZN( u0_out6_3 ) , .A3( u0_u6_u4_n166 ) , .A1( u0_u6_u4_n167 ) , .A2( u0_u6_u4_n186 ) );
  NAND3_X1 u0_u6_u4_U97 (.A3( u0_u6_u4_n146 ) , .A2( u0_u6_u4_n147 ) , .A1( u0_u6_u4_n148 ) , .ZN( u0_u6_u4_n149 ) );
  NAND3_X1 u0_u6_u4_U98 (.A3( u0_u6_u4_n143 ) , .A2( u0_u6_u4_n144 ) , .A1( u0_u6_u4_n145 ) , .ZN( u0_u6_u4_n151 ) );
  NAND3_X1 u0_u6_u4_U99 (.A3( u0_u6_u4_n121 ) , .ZN( u0_u6_u4_n122 ) , .A2( u0_u6_u4_n144 ) , .A1( u0_u6_u4_n154 ) );
  AOI21_X1 u0_u6_u6_U10 (.ZN( u0_u6_u6_n106 ) , .A( u0_u6_u6_n142 ) , .B2( u0_u6_u6_n159 ) , .B1( u0_u6_u6_n164 ) );
  INV_X1 u0_u6_u6_U11 (.A( u0_u6_u6_n155 ) , .ZN( u0_u6_u6_n161 ) );
  INV_X1 u0_u6_u6_U12 (.A( u0_u6_u6_n128 ) , .ZN( u0_u6_u6_n164 ) );
  NAND2_X1 u0_u6_u6_U13 (.ZN( u0_u6_u6_n110 ) , .A1( u0_u6_u6_n122 ) , .A2( u0_u6_u6_n129 ) );
  NAND2_X1 u0_u6_u6_U14 (.ZN( u0_u6_u6_n124 ) , .A2( u0_u6_u6_n146 ) , .A1( u0_u6_u6_n148 ) );
  INV_X1 u0_u6_u6_U15 (.A( u0_u6_u6_n132 ) , .ZN( u0_u6_u6_n171 ) );
  AND2_X1 u0_u6_u6_U16 (.A1( u0_u6_u6_n100 ) , .ZN( u0_u6_u6_n130 ) , .A2( u0_u6_u6_n147 ) );
  INV_X1 u0_u6_u6_U17 (.A( u0_u6_u6_n127 ) , .ZN( u0_u6_u6_n173 ) );
  INV_X1 u0_u6_u6_U18 (.A( u0_u6_u6_n121 ) , .ZN( u0_u6_u6_n167 ) );
  INV_X1 u0_u6_u6_U19 (.A( u0_u6_u6_n100 ) , .ZN( u0_u6_u6_n169 ) );
  INV_X1 u0_u6_u6_U20 (.A( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n170 ) );
  INV_X1 u0_u6_u6_U21 (.A( u0_u6_u6_n113 ) , .ZN( u0_u6_u6_n168 ) );
  AND2_X1 u0_u6_u6_U22 (.A1( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n119 ) , .ZN( u0_u6_u6_n133 ) );
  AND2_X1 u0_u6_u6_U23 (.A2( u0_u6_u6_n121 ) , .A1( u0_u6_u6_n122 ) , .ZN( u0_u6_u6_n131 ) );
  AND3_X1 u0_u6_u6_U24 (.ZN( u0_u6_u6_n120 ) , .A2( u0_u6_u6_n127 ) , .A1( u0_u6_u6_n132 ) , .A3( u0_u6_u6_n145 ) );
  INV_X1 u0_u6_u6_U25 (.A( u0_u6_u6_n146 ) , .ZN( u0_u6_u6_n163 ) );
  AOI222_X1 u0_u6_u6_U26 (.ZN( u0_u6_u6_n114 ) , .A1( u0_u6_u6_n118 ) , .A2( u0_u6_u6_n126 ) , .B2( u0_u6_u6_n151 ) , .C2( u0_u6_u6_n159 ) , .C1( u0_u6_u6_n168 ) , .B1( u0_u6_u6_n169 ) );
  NOR2_X1 u0_u6_u6_U27 (.A1( u0_u6_u6_n162 ) , .A2( u0_u6_u6_n165 ) , .ZN( u0_u6_u6_n98 ) );
  AOI211_X1 u0_u6_u6_U28 (.B( u0_u6_u6_n149 ) , .A( u0_u6_u6_n150 ) , .C2( u0_u6_u6_n151 ) , .C1( u0_u6_u6_n152 ) , .ZN( u0_u6_u6_n153 ) );
  AOI21_X1 u0_u6_u6_U29 (.B2( u0_u6_u6_n147 ) , .B1( u0_u6_u6_n148 ) , .ZN( u0_u6_u6_n149 ) , .A( u0_u6_u6_n158 ) );
  INV_X1 u0_u6_u6_U3 (.A( u0_u6_u6_n110 ) , .ZN( u0_u6_u6_n166 ) );
  AOI21_X1 u0_u6_u6_U30 (.A( u0_u6_u6_n144 ) , .B2( u0_u6_u6_n145 ) , .B1( u0_u6_u6_n146 ) , .ZN( u0_u6_u6_n150 ) );
  NAND2_X1 u0_u6_u6_U31 (.A2( u0_u6_u6_n143 ) , .ZN( u0_u6_u6_n152 ) , .A1( u0_u6_u6_n166 ) );
  NAND2_X1 u0_u6_u6_U32 (.A1( u0_u6_u6_n144 ) , .ZN( u0_u6_u6_n151 ) , .A2( u0_u6_u6_n158 ) );
  NAND2_X1 u0_u6_u6_U33 (.ZN( u0_u6_u6_n132 ) , .A1( u0_u6_u6_n91 ) , .A2( u0_u6_u6_n97 ) );
  AOI22_X1 u0_u6_u6_U34 (.B2( u0_u6_u6_n110 ) , .B1( u0_u6_u6_n111 ) , .A1( u0_u6_u6_n112 ) , .ZN( u0_u6_u6_n115 ) , .A2( u0_u6_u6_n161 ) );
  NAND4_X1 u0_u6_u6_U35 (.A3( u0_u6_u6_n109 ) , .ZN( u0_u6_u6_n112 ) , .A4( u0_u6_u6_n132 ) , .A2( u0_u6_u6_n147 ) , .A1( u0_u6_u6_n166 ) );
  NOR2_X1 u0_u6_u6_U36 (.ZN( u0_u6_u6_n109 ) , .A1( u0_u6_u6_n170 ) , .A2( u0_u6_u6_n173 ) );
  NOR2_X1 u0_u6_u6_U37 (.A2( u0_u6_u6_n126 ) , .ZN( u0_u6_u6_n155 ) , .A1( u0_u6_u6_n160 ) );
  NAND2_X1 u0_u6_u6_U38 (.ZN( u0_u6_u6_n146 ) , .A2( u0_u6_u6_n94 ) , .A1( u0_u6_u6_n99 ) );
  AOI211_X1 u0_u6_u6_U39 (.B( u0_u6_u6_n134 ) , .A( u0_u6_u6_n135 ) , .C1( u0_u6_u6_n136 ) , .ZN( u0_u6_u6_n137 ) , .C2( u0_u6_u6_n151 ) );
  AOI22_X1 u0_u6_u6_U4 (.B2( u0_u6_u6_n101 ) , .A1( u0_u6_u6_n102 ) , .ZN( u0_u6_u6_n103 ) , .B1( u0_u6_u6_n160 ) , .A2( u0_u6_u6_n161 ) );
  NAND4_X1 u0_u6_u6_U40 (.A4( u0_u6_u6_n127 ) , .A3( u0_u6_u6_n128 ) , .A2( u0_u6_u6_n129 ) , .A1( u0_u6_u6_n130 ) , .ZN( u0_u6_u6_n136 ) );
  AOI21_X1 u0_u6_u6_U41 (.B2( u0_u6_u6_n132 ) , .B1( u0_u6_u6_n133 ) , .ZN( u0_u6_u6_n134 ) , .A( u0_u6_u6_n158 ) );
  AOI21_X1 u0_u6_u6_U42 (.B1( u0_u6_u6_n131 ) , .ZN( u0_u6_u6_n135 ) , .A( u0_u6_u6_n144 ) , .B2( u0_u6_u6_n146 ) );
  INV_X1 u0_u6_u6_U43 (.A( u0_u6_u6_n111 ) , .ZN( u0_u6_u6_n158 ) );
  NAND2_X1 u0_u6_u6_U44 (.ZN( u0_u6_u6_n127 ) , .A1( u0_u6_u6_n91 ) , .A2( u0_u6_u6_n92 ) );
  NAND2_X1 u0_u6_u6_U45 (.ZN( u0_u6_u6_n129 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n96 ) );
  INV_X1 u0_u6_u6_U46 (.A( u0_u6_u6_n144 ) , .ZN( u0_u6_u6_n159 ) );
  NAND2_X1 u0_u6_u6_U47 (.ZN( u0_u6_u6_n145 ) , .A2( u0_u6_u6_n97 ) , .A1( u0_u6_u6_n98 ) );
  NAND2_X1 u0_u6_u6_U48 (.ZN( u0_u6_u6_n148 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n94 ) );
  NAND2_X1 u0_u6_u6_U49 (.ZN( u0_u6_u6_n108 ) , .A2( u0_u6_u6_n139 ) , .A1( u0_u6_u6_n144 ) );
  NOR2_X1 u0_u6_u6_U5 (.A1( u0_u6_u6_n118 ) , .ZN( u0_u6_u6_n143 ) , .A2( u0_u6_u6_n168 ) );
  NAND2_X1 u0_u6_u6_U50 (.ZN( u0_u6_u6_n121 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n97 ) );
  NAND2_X1 u0_u6_u6_U51 (.ZN( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n95 ) );
  AND2_X1 u0_u6_u6_U52 (.ZN( u0_u6_u6_n118 ) , .A2( u0_u6_u6_n91 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U53 (.ZN( u0_u6_u6_n147 ) , .A2( u0_u6_u6_n98 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U54 (.ZN( u0_u6_u6_n128 ) , .A1( u0_u6_u6_n94 ) , .A2( u0_u6_u6_n96 ) );
  NAND2_X1 u0_u6_u6_U55 (.ZN( u0_u6_u6_n119 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U56 (.ZN( u0_u6_u6_n123 ) , .A2( u0_u6_u6_n91 ) , .A1( u0_u6_u6_n96 ) );
  NAND2_X1 u0_u6_u6_U57 (.ZN( u0_u6_u6_n100 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n98 ) );
  NAND2_X1 u0_u6_u6_U58 (.ZN( u0_u6_u6_n122 ) , .A1( u0_u6_u6_n94 ) , .A2( u0_u6_u6_n97 ) );
  INV_X1 u0_u6_u6_U59 (.A( u0_u6_u6_n139 ) , .ZN( u0_u6_u6_n160 ) );
  AOI21_X1 u0_u6_u6_U6 (.B1( u0_u6_u6_n107 ) , .B2( u0_u6_u6_n132 ) , .A( u0_u6_u6_n158 ) , .ZN( u0_u6_u6_n88 ) );
  NAND2_X1 u0_u6_u6_U60 (.ZN( u0_u6_u6_n113 ) , .A1( u0_u6_u6_n96 ) , .A2( u0_u6_u6_n98 ) );
  NOR2_X1 u0_u6_u6_U61 (.A2( u0_u6_X_40 ) , .A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n126 ) );
  NOR2_X1 u0_u6_u6_U62 (.A2( u0_u6_X_39 ) , .A1( u0_u6_X_42 ) , .ZN( u0_u6_u6_n92 ) );
  NOR2_X1 u0_u6_u6_U63 (.A2( u0_u6_X_39 ) , .A1( u0_u6_u6_n156 ) , .ZN( u0_u6_u6_n97 ) );
  NOR2_X1 u0_u6_u6_U64 (.A2( u0_u6_X_38 ) , .A1( u0_u6_u6_n165 ) , .ZN( u0_u6_u6_n95 ) );
  NOR2_X1 u0_u6_u6_U65 (.A2( u0_u6_X_41 ) , .ZN( u0_u6_u6_n111 ) , .A1( u0_u6_u6_n157 ) );
  NOR2_X1 u0_u6_u6_U66 (.A2( u0_u6_X_37 ) , .A1( u0_u6_u6_n162 ) , .ZN( u0_u6_u6_n94 ) );
  NOR2_X1 u0_u6_u6_U67 (.A2( u0_u6_X_37 ) , .A1( u0_u6_X_38 ) , .ZN( u0_u6_u6_n91 ) );
  NAND2_X1 u0_u6_u6_U68 (.A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n144 ) , .A2( u0_u6_u6_n157 ) );
  NAND2_X1 u0_u6_u6_U69 (.A2( u0_u6_X_40 ) , .A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n139 ) );
  OAI21_X1 u0_u6_u6_U7 (.A( u0_u6_u6_n159 ) , .B1( u0_u6_u6_n169 ) , .B2( u0_u6_u6_n173 ) , .ZN( u0_u6_u6_n90 ) );
  AND2_X1 u0_u6_u6_U70 (.A1( u0_u6_X_39 ) , .A2( u0_u6_u6_n156 ) , .ZN( u0_u6_u6_n96 ) );
  AND2_X1 u0_u6_u6_U71 (.A1( u0_u6_X_39 ) , .A2( u0_u6_X_42 ) , .ZN( u0_u6_u6_n99 ) );
  INV_X1 u0_u6_u6_U72 (.A( u0_u6_X_40 ) , .ZN( u0_u6_u6_n157 ) );
  INV_X1 u0_u6_u6_U73 (.A( u0_u6_X_37 ) , .ZN( u0_u6_u6_n165 ) );
  INV_X1 u0_u6_u6_U74 (.A( u0_u6_X_38 ) , .ZN( u0_u6_u6_n162 ) );
  INV_X1 u0_u6_u6_U75 (.A( u0_u6_X_42 ) , .ZN( u0_u6_u6_n156 ) );
  NAND4_X1 u0_u6_u6_U76 (.ZN( u0_out6_32 ) , .A4( u0_u6_u6_n103 ) , .A3( u0_u6_u6_n104 ) , .A2( u0_u6_u6_n105 ) , .A1( u0_u6_u6_n106 ) );
  AOI22_X1 u0_u6_u6_U77 (.ZN( u0_u6_u6_n104 ) , .A1( u0_u6_u6_n111 ) , .B1( u0_u6_u6_n124 ) , .B2( u0_u6_u6_n151 ) , .A2( u0_u6_u6_n93 ) );
  AOI22_X1 u0_u6_u6_U78 (.ZN( u0_u6_u6_n105 ) , .A2( u0_u6_u6_n108 ) , .A1( u0_u6_u6_n118 ) , .B2( u0_u6_u6_n126 ) , .B1( u0_u6_u6_n171 ) );
  NAND4_X1 u0_u6_u6_U79 (.ZN( u0_out6_12 ) , .A4( u0_u6_u6_n114 ) , .A3( u0_u6_u6_n115 ) , .A2( u0_u6_u6_n116 ) , .A1( u0_u6_u6_n117 ) );
  INV_X1 u0_u6_u6_U8 (.ZN( u0_u6_u6_n172 ) , .A( u0_u6_u6_n88 ) );
  OAI22_X1 u0_u6_u6_U80 (.B2( u0_u6_u6_n111 ) , .ZN( u0_u6_u6_n116 ) , .B1( u0_u6_u6_n126 ) , .A2( u0_u6_u6_n164 ) , .A1( u0_u6_u6_n167 ) );
  OAI21_X1 u0_u6_u6_U81 (.A( u0_u6_u6_n108 ) , .ZN( u0_u6_u6_n117 ) , .B2( u0_u6_u6_n141 ) , .B1( u0_u6_u6_n163 ) );
  OAI211_X1 u0_u6_u6_U82 (.ZN( u0_out6_22 ) , .B( u0_u6_u6_n137 ) , .A( u0_u6_u6_n138 ) , .C2( u0_u6_u6_n139 ) , .C1( u0_u6_u6_n140 ) );
  AOI22_X1 u0_u6_u6_U83 (.B1( u0_u6_u6_n124 ) , .A2( u0_u6_u6_n125 ) , .A1( u0_u6_u6_n126 ) , .ZN( u0_u6_u6_n138 ) , .B2( u0_u6_u6_n161 ) );
  AND4_X1 u0_u6_u6_U84 (.A3( u0_u6_u6_n119 ) , .A1( u0_u6_u6_n120 ) , .A4( u0_u6_u6_n129 ) , .ZN( u0_u6_u6_n140 ) , .A2( u0_u6_u6_n143 ) );
  OAI211_X1 u0_u6_u6_U85 (.ZN( u0_out6_7 ) , .B( u0_u6_u6_n153 ) , .C2( u0_u6_u6_n154 ) , .C1( u0_u6_u6_n155 ) , .A( u0_u6_u6_n174 ) );
  NOR3_X1 u0_u6_u6_U86 (.A1( u0_u6_u6_n141 ) , .ZN( u0_u6_u6_n154 ) , .A3( u0_u6_u6_n164 ) , .A2( u0_u6_u6_n171 ) );
  INV_X1 u0_u6_u6_U87 (.A( u0_u6_u6_n142 ) , .ZN( u0_u6_u6_n174 ) );
  NAND3_X1 u0_u6_u6_U88 (.A2( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n125 ) , .A1( u0_u6_u6_n130 ) , .A3( u0_u6_u6_n131 ) );
  NAND3_X1 u0_u6_u6_U89 (.A3( u0_u6_u6_n133 ) , .ZN( u0_u6_u6_n141 ) , .A1( u0_u6_u6_n145 ) , .A2( u0_u6_u6_n148 ) );
  AOI22_X1 u0_u6_u6_U9 (.A2( u0_u6_u6_n151 ) , .B2( u0_u6_u6_n161 ) , .A1( u0_u6_u6_n167 ) , .B1( u0_u6_u6_n170 ) , .ZN( u0_u6_u6_n89 ) );
  NAND3_X1 u0_u6_u6_U90 (.ZN( u0_u6_u6_n101 ) , .A3( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n121 ) , .A1( u0_u6_u6_n127 ) );
  NAND3_X1 u0_u6_u6_U91 (.ZN( u0_u6_u6_n102 ) , .A3( u0_u6_u6_n130 ) , .A2( u0_u6_u6_n145 ) , .A1( u0_u6_u6_n166 ) );
  NAND3_X1 u0_u6_u6_U92 (.A3( u0_u6_u6_n113 ) , .A1( u0_u6_u6_n119 ) , .A2( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n93 ) );
  NAND3_X1 u0_u6_u6_U93 (.ZN( u0_u6_u6_n142 ) , .A2( u0_u6_u6_n172 ) , .A3( u0_u6_u6_n89 ) , .A1( u0_u6_u6_n90 ) );
  AND3_X1 u0_u6_u7_U10 (.A3( u0_u6_u7_n110 ) , .A2( u0_u6_u7_n127 ) , .A1( u0_u6_u7_n132 ) , .ZN( u0_u6_u7_n92 ) );
  OAI21_X1 u0_u6_u7_U11 (.A( u0_u6_u7_n161 ) , .B1( u0_u6_u7_n168 ) , .B2( u0_u6_u7_n173 ) , .ZN( u0_u6_u7_n91 ) );
  AOI211_X1 u0_u6_u7_U12 (.A( u0_u6_u7_n117 ) , .ZN( u0_u6_u7_n118 ) , .C2( u0_u6_u7_n126 ) , .C1( u0_u6_u7_n177 ) , .B( u0_u6_u7_n180 ) );
  OAI22_X1 u0_u6_u7_U13 (.B1( u0_u6_u7_n115 ) , .ZN( u0_u6_u7_n117 ) , .A2( u0_u6_u7_n133 ) , .A1( u0_u6_u7_n137 ) , .B2( u0_u6_u7_n162 ) );
  INV_X1 u0_u6_u7_U14 (.A( u0_u6_u7_n116 ) , .ZN( u0_u6_u7_n180 ) );
  NOR3_X1 u0_u6_u7_U15 (.ZN( u0_u6_u7_n115 ) , .A3( u0_u6_u7_n145 ) , .A2( u0_u6_u7_n168 ) , .A1( u0_u6_u7_n169 ) );
  OAI211_X1 u0_u6_u7_U16 (.B( u0_u6_u7_n122 ) , .A( u0_u6_u7_n123 ) , .C2( u0_u6_u7_n124 ) , .ZN( u0_u6_u7_n154 ) , .C1( u0_u6_u7_n162 ) );
  AOI222_X1 u0_u6_u7_U17 (.ZN( u0_u6_u7_n122 ) , .C2( u0_u6_u7_n126 ) , .C1( u0_u6_u7_n145 ) , .B1( u0_u6_u7_n161 ) , .A2( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n170 ) , .A1( u0_u6_u7_n176 ) );
  INV_X1 u0_u6_u7_U18 (.A( u0_u6_u7_n133 ) , .ZN( u0_u6_u7_n176 ) );
  NOR3_X1 u0_u6_u7_U19 (.A2( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n135 ) , .ZN( u0_u6_u7_n136 ) , .A3( u0_u6_u7_n171 ) );
  NOR2_X1 u0_u6_u7_U20 (.A1( u0_u6_u7_n130 ) , .A2( u0_u6_u7_n134 ) , .ZN( u0_u6_u7_n153 ) );
  INV_X1 u0_u6_u7_U21 (.A( u0_u6_u7_n101 ) , .ZN( u0_u6_u7_n165 ) );
  NOR2_X1 u0_u6_u7_U22 (.ZN( u0_u6_u7_n111 ) , .A2( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n169 ) );
  AOI21_X1 u0_u6_u7_U23 (.ZN( u0_u6_u7_n104 ) , .B2( u0_u6_u7_n112 ) , .B1( u0_u6_u7_n127 ) , .A( u0_u6_u7_n164 ) );
  AOI21_X1 u0_u6_u7_U24 (.ZN( u0_u6_u7_n106 ) , .B1( u0_u6_u7_n133 ) , .B2( u0_u6_u7_n146 ) , .A( u0_u6_u7_n162 ) );
  AOI21_X1 u0_u6_u7_U25 (.A( u0_u6_u7_n101 ) , .ZN( u0_u6_u7_n107 ) , .B2( u0_u6_u7_n128 ) , .B1( u0_u6_u7_n175 ) );
  INV_X1 u0_u6_u7_U26 (.A( u0_u6_u7_n138 ) , .ZN( u0_u6_u7_n171 ) );
  INV_X1 u0_u6_u7_U27 (.A( u0_u6_u7_n131 ) , .ZN( u0_u6_u7_n177 ) );
  INV_X1 u0_u6_u7_U28 (.A( u0_u6_u7_n110 ) , .ZN( u0_u6_u7_n174 ) );
  NAND2_X1 u0_u6_u7_U29 (.A1( u0_u6_u7_n129 ) , .A2( u0_u6_u7_n132 ) , .ZN( u0_u6_u7_n149 ) );
  OAI21_X1 u0_u6_u7_U3 (.ZN( u0_u6_u7_n159 ) , .A( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n171 ) , .B1( u0_u6_u7_n174 ) );
  NAND2_X1 u0_u6_u7_U30 (.A1( u0_u6_u7_n113 ) , .A2( u0_u6_u7_n124 ) , .ZN( u0_u6_u7_n130 ) );
  INV_X1 u0_u6_u7_U31 (.A( u0_u6_u7_n112 ) , .ZN( u0_u6_u7_n173 ) );
  INV_X1 u0_u6_u7_U32 (.A( u0_u6_u7_n128 ) , .ZN( u0_u6_u7_n168 ) );
  INV_X1 u0_u6_u7_U33 (.A( u0_u6_u7_n148 ) , .ZN( u0_u6_u7_n169 ) );
  INV_X1 u0_u6_u7_U34 (.A( u0_u6_u7_n127 ) , .ZN( u0_u6_u7_n179 ) );
  NOR2_X1 u0_u6_u7_U35 (.ZN( u0_u6_u7_n101 ) , .A2( u0_u6_u7_n150 ) , .A1( u0_u6_u7_n156 ) );
  AOI211_X1 u0_u6_u7_U36 (.B( u0_u6_u7_n154 ) , .A( u0_u6_u7_n155 ) , .C1( u0_u6_u7_n156 ) , .ZN( u0_u6_u7_n157 ) , .C2( u0_u6_u7_n172 ) );
  INV_X1 u0_u6_u7_U37 (.A( u0_u6_u7_n153 ) , .ZN( u0_u6_u7_n172 ) );
  AOI211_X1 u0_u6_u7_U38 (.B( u0_u6_u7_n139 ) , .A( u0_u6_u7_n140 ) , .C2( u0_u6_u7_n141 ) , .ZN( u0_u6_u7_n142 ) , .C1( u0_u6_u7_n156 ) );
  NAND4_X1 u0_u6_u7_U39 (.A3( u0_u6_u7_n127 ) , .A2( u0_u6_u7_n128 ) , .A1( u0_u6_u7_n129 ) , .ZN( u0_u6_u7_n141 ) , .A4( u0_u6_u7_n147 ) );
  INV_X1 u0_u6_u7_U4 (.A( u0_u6_u7_n111 ) , .ZN( u0_u6_u7_n170 ) );
  AOI21_X1 u0_u6_u7_U40 (.A( u0_u6_u7_n137 ) , .B1( u0_u6_u7_n138 ) , .ZN( u0_u6_u7_n139 ) , .B2( u0_u6_u7_n146 ) );
  OAI22_X1 u0_u6_u7_U41 (.B1( u0_u6_u7_n136 ) , .ZN( u0_u6_u7_n140 ) , .A1( u0_u6_u7_n153 ) , .B2( u0_u6_u7_n162 ) , .A2( u0_u6_u7_n164 ) );
  AOI21_X1 u0_u6_u7_U42 (.ZN( u0_u6_u7_n123 ) , .B1( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n177 ) , .A( u0_u6_u7_n97 ) );
  AOI21_X1 u0_u6_u7_U43 (.B2( u0_u6_u7_n113 ) , .B1( u0_u6_u7_n124 ) , .A( u0_u6_u7_n125 ) , .ZN( u0_u6_u7_n97 ) );
  INV_X1 u0_u6_u7_U44 (.A( u0_u6_u7_n125 ) , .ZN( u0_u6_u7_n161 ) );
  INV_X1 u0_u6_u7_U45 (.A( u0_u6_u7_n152 ) , .ZN( u0_u6_u7_n162 ) );
  AOI22_X1 u0_u6_u7_U46 (.A2( u0_u6_u7_n114 ) , .ZN( u0_u6_u7_n119 ) , .B1( u0_u6_u7_n130 ) , .A1( u0_u6_u7_n156 ) , .B2( u0_u6_u7_n165 ) );
  NAND2_X1 u0_u6_u7_U47 (.A2( u0_u6_u7_n112 ) , .ZN( u0_u6_u7_n114 ) , .A1( u0_u6_u7_n175 ) );
  AND2_X1 u0_u6_u7_U48 (.ZN( u0_u6_u7_n145 ) , .A2( u0_u6_u7_n98 ) , .A1( u0_u6_u7_n99 ) );
  NOR2_X1 u0_u6_u7_U49 (.ZN( u0_u6_u7_n137 ) , .A1( u0_u6_u7_n150 ) , .A2( u0_u6_u7_n161 ) );
  INV_X1 u0_u6_u7_U5 (.A( u0_u6_u7_n149 ) , .ZN( u0_u6_u7_n175 ) );
  AOI21_X1 u0_u6_u7_U50 (.ZN( u0_u6_u7_n105 ) , .B2( u0_u6_u7_n110 ) , .A( u0_u6_u7_n125 ) , .B1( u0_u6_u7_n147 ) );
  NAND2_X1 u0_u6_u7_U51 (.ZN( u0_u6_u7_n146 ) , .A1( u0_u6_u7_n95 ) , .A2( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U52 (.A2( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n147 ) , .A1( u0_u6_u7_n93 ) );
  NAND2_X1 u0_u6_u7_U53 (.A1( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n127 ) , .A2( u0_u6_u7_n99 ) );
  OR2_X1 u0_u6_u7_U54 (.ZN( u0_u6_u7_n126 ) , .A2( u0_u6_u7_n152 ) , .A1( u0_u6_u7_n156 ) );
  NAND2_X1 u0_u6_u7_U55 (.A2( u0_u6_u7_n102 ) , .A1( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n133 ) );
  NAND2_X1 u0_u6_u7_U56 (.ZN( u0_u6_u7_n112 ) , .A2( u0_u6_u7_n96 ) , .A1( u0_u6_u7_n99 ) );
  NAND2_X1 u0_u6_u7_U57 (.A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n128 ) , .A1( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U58 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n113 ) , .A2( u0_u6_u7_n93 ) );
  NAND2_X1 u0_u6_u7_U59 (.A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n124 ) , .A1( u0_u6_u7_n96 ) );
  INV_X1 u0_u6_u7_U6 (.A( u0_u6_u7_n154 ) , .ZN( u0_u6_u7_n178 ) );
  NAND2_X1 u0_u6_u7_U60 (.ZN( u0_u6_u7_n110 ) , .A1( u0_u6_u7_n95 ) , .A2( u0_u6_u7_n96 ) );
  INV_X1 u0_u6_u7_U61 (.A( u0_u6_u7_n150 ) , .ZN( u0_u6_u7_n164 ) );
  AND2_X1 u0_u6_u7_U62 (.ZN( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n93 ) , .A2( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U63 (.A1( u0_u6_u7_n100 ) , .A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n129 ) );
  NAND2_X1 u0_u6_u7_U64 (.A2( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n131 ) , .A1( u0_u6_u7_n95 ) );
  NAND2_X1 u0_u6_u7_U65 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n138 ) , .A2( u0_u6_u7_n99 ) );
  NAND2_X1 u0_u6_u7_U66 (.ZN( u0_u6_u7_n132 ) , .A1( u0_u6_u7_n93 ) , .A2( u0_u6_u7_n96 ) );
  NAND2_X1 u0_u6_u7_U67 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n148 ) , .A2( u0_u6_u7_n95 ) );
  NOR2_X1 u0_u6_u7_U68 (.A2( u0_u6_X_47 ) , .ZN( u0_u6_u7_n150 ) , .A1( u0_u6_u7_n163 ) );
  NOR2_X1 u0_u6_u7_U69 (.A2( u0_u6_X_43 ) , .A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n103 ) );
  AOI211_X1 u0_u6_u7_U7 (.ZN( u0_u6_u7_n116 ) , .A( u0_u6_u7_n155 ) , .C1( u0_u6_u7_n161 ) , .C2( u0_u6_u7_n171 ) , .B( u0_u6_u7_n94 ) );
  NOR2_X1 u0_u6_u7_U70 (.A2( u0_u6_X_48 ) , .A1( u0_u6_u7_n166 ) , .ZN( u0_u6_u7_n95 ) );
  NOR2_X1 u0_u6_u7_U71 (.A2( u0_u6_X_45 ) , .A1( u0_u6_X_48 ) , .ZN( u0_u6_u7_n99 ) );
  NOR2_X1 u0_u6_u7_U72 (.A2( u0_u6_X_44 ) , .A1( u0_u6_u7_n167 ) , .ZN( u0_u6_u7_n98 ) );
  NOR2_X1 u0_u6_u7_U73 (.A2( u0_u6_X_46 ) , .A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n152 ) );
  AND2_X1 u0_u6_u7_U74 (.A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n156 ) , .A2( u0_u6_u7_n163 ) );
  NAND2_X1 u0_u6_u7_U75 (.A2( u0_u6_X_46 ) , .A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n125 ) );
  AND2_X1 u0_u6_u7_U76 (.A2( u0_u6_X_45 ) , .A1( u0_u6_X_48 ) , .ZN( u0_u6_u7_n102 ) );
  AND2_X1 u0_u6_u7_U77 (.A2( u0_u6_X_43 ) , .A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n96 ) );
  AND2_X1 u0_u6_u7_U78 (.A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n100 ) , .A2( u0_u6_u7_n167 ) );
  AND2_X1 u0_u6_u7_U79 (.A1( u0_u6_X_48 ) , .A2( u0_u6_u7_n166 ) , .ZN( u0_u6_u7_n93 ) );
  OAI222_X1 u0_u6_u7_U8 (.C2( u0_u6_u7_n101 ) , .B2( u0_u6_u7_n111 ) , .A1( u0_u6_u7_n113 ) , .C1( u0_u6_u7_n146 ) , .A2( u0_u6_u7_n162 ) , .B1( u0_u6_u7_n164 ) , .ZN( u0_u6_u7_n94 ) );
  INV_X1 u0_u6_u7_U80 (.A( u0_u6_X_46 ) , .ZN( u0_u6_u7_n163 ) );
  INV_X1 u0_u6_u7_U81 (.A( u0_u6_X_43 ) , .ZN( u0_u6_u7_n167 ) );
  INV_X1 u0_u6_u7_U82 (.A( u0_u6_X_45 ) , .ZN( u0_u6_u7_n166 ) );
  NAND4_X1 u0_u6_u7_U83 (.ZN( u0_out6_5 ) , .A4( u0_u6_u7_n108 ) , .A3( u0_u6_u7_n109 ) , .A1( u0_u6_u7_n116 ) , .A2( u0_u6_u7_n123 ) );
  AOI22_X1 u0_u6_u7_U84 (.ZN( u0_u6_u7_n109 ) , .A2( u0_u6_u7_n126 ) , .B2( u0_u6_u7_n145 ) , .B1( u0_u6_u7_n156 ) , .A1( u0_u6_u7_n171 ) );
  NOR4_X1 u0_u6_u7_U85 (.A4( u0_u6_u7_n104 ) , .A3( u0_u6_u7_n105 ) , .A2( u0_u6_u7_n106 ) , .A1( u0_u6_u7_n107 ) , .ZN( u0_u6_u7_n108 ) );
  NAND4_X1 u0_u6_u7_U86 (.ZN( u0_out6_27 ) , .A4( u0_u6_u7_n118 ) , .A3( u0_u6_u7_n119 ) , .A2( u0_u6_u7_n120 ) , .A1( u0_u6_u7_n121 ) );
  OAI21_X1 u0_u6_u7_U87 (.ZN( u0_u6_u7_n121 ) , .B2( u0_u6_u7_n145 ) , .A( u0_u6_u7_n150 ) , .B1( u0_u6_u7_n174 ) );
  OAI21_X1 u0_u6_u7_U88 (.ZN( u0_u6_u7_n120 ) , .A( u0_u6_u7_n161 ) , .B2( u0_u6_u7_n170 ) , .B1( u0_u6_u7_n179 ) );
  NAND4_X1 u0_u6_u7_U89 (.ZN( u0_out6_21 ) , .A4( u0_u6_u7_n157 ) , .A3( u0_u6_u7_n158 ) , .A2( u0_u6_u7_n159 ) , .A1( u0_u6_u7_n160 ) );
  OAI221_X1 u0_u6_u7_U9 (.C1( u0_u6_u7_n101 ) , .C2( u0_u6_u7_n147 ) , .ZN( u0_u6_u7_n155 ) , .B2( u0_u6_u7_n162 ) , .A( u0_u6_u7_n91 ) , .B1( u0_u6_u7_n92 ) );
  OAI21_X1 u0_u6_u7_U90 (.B1( u0_u6_u7_n145 ) , .ZN( u0_u6_u7_n160 ) , .A( u0_u6_u7_n161 ) , .B2( u0_u6_u7_n177 ) );
  AOI22_X1 u0_u6_u7_U91 (.B2( u0_u6_u7_n149 ) , .B1( u0_u6_u7_n150 ) , .A2( u0_u6_u7_n151 ) , .A1( u0_u6_u7_n152 ) , .ZN( u0_u6_u7_n158 ) );
  NAND4_X1 u0_u6_u7_U92 (.ZN( u0_out6_15 ) , .A4( u0_u6_u7_n142 ) , .A3( u0_u6_u7_n143 ) , .A2( u0_u6_u7_n144 ) , .A1( u0_u6_u7_n178 ) );
  OR2_X1 u0_u6_u7_U93 (.A2( u0_u6_u7_n125 ) , .A1( u0_u6_u7_n129 ) , .ZN( u0_u6_u7_n144 ) );
  AOI22_X1 u0_u6_u7_U94 (.A2( u0_u6_u7_n126 ) , .ZN( u0_u6_u7_n143 ) , .B2( u0_u6_u7_n165 ) , .B1( u0_u6_u7_n173 ) , .A1( u0_u6_u7_n174 ) );
  NAND3_X1 u0_u6_u7_U95 (.A3( u0_u6_u7_n146 ) , .A2( u0_u6_u7_n147 ) , .A1( u0_u6_u7_n148 ) , .ZN( u0_u6_u7_n151 ) );
  NAND3_X1 u0_u6_u7_U96 (.A3( u0_u6_u7_n131 ) , .A2( u0_u6_u7_n132 ) , .A1( u0_u6_u7_n133 ) , .ZN( u0_u6_u7_n135 ) );
  XOR2_X1 u0_u7_U1 (.B( u0_K8_9 ) , .A( u0_R6_6 ) , .Z( u0_u7_X_9 ) );
  XOR2_X1 u0_u7_U10 (.B( u0_K8_45 ) , .A( u0_R6_30 ) , .Z( u0_u7_X_45 ) );
  XOR2_X1 u0_u7_U15 (.B( u0_K8_40 ) , .A( u0_R6_27 ) , .Z( u0_u7_X_40 ) );
  XOR2_X1 u0_u7_U16 (.B( u0_K8_3 ) , .A( u0_R6_2 ) , .Z( u0_u7_X_3 ) );
  XOR2_X1 u0_u7_U18 (.B( u0_K8_38 ) , .A( u0_R6_25 ) , .Z( u0_u7_X_38 ) );
  XOR2_X1 u0_u7_U20 (.B( u0_K8_36 ) , .A( u0_R6_25 ) , .Z( u0_u7_X_36 ) );
  XOR2_X1 u0_u7_U22 (.B( u0_K8_34 ) , .A( u0_R6_23 ) , .Z( u0_u7_X_34 ) );
  XOR2_X1 u0_u7_U23 (.B( u0_K8_33 ) , .A( u0_R6_22 ) , .Z( u0_u7_X_33 ) );
  XOR2_X1 u0_u7_U24 (.B( u0_K8_32 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_32 ) );
  XOR2_X1 u0_u7_U25 (.B( u0_K8_31 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_31 ) );
  XOR2_X1 u0_u7_U26 (.B( u0_K8_30 ) , .A( u0_R6_21 ) , .Z( u0_u7_X_30 ) );
  XOR2_X1 u0_u7_U27 (.B( u0_K8_2 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_2 ) );
  XOR2_X1 u0_u7_U28 (.B( u0_K8_29 ) , .A( u0_R6_20 ) , .Z( u0_u7_X_29 ) );
  XOR2_X1 u0_u7_U29 (.B( u0_K8_28 ) , .A( u0_R6_19 ) , .Z( u0_u7_X_28 ) );
  XOR2_X1 u0_u7_U30 (.B( u0_K8_27 ) , .A( u0_R6_18 ) , .Z( u0_u7_X_27 ) );
  XOR2_X1 u0_u7_U32 (.B( u0_K8_25 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_25 ) );
  XOR2_X1 u0_u7_U34 (.B( u0_K8_23 ) , .A( u0_R6_16 ) , .Z( u0_u7_X_23 ) );
  XOR2_X1 u0_u7_U35 (.B( u0_K8_22 ) , .A( u0_R6_15 ) , .Z( u0_u7_X_22 ) );
  XOR2_X1 u0_u7_U38 (.B( u0_K8_1 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_1 ) );
  XOR2_X1 u0_u7_U6 (.B( u0_K8_4 ) , .A( u0_R6_3 ) , .Z( u0_u7_X_4 ) );
  XOR2_X1 u0_u7_U7 (.B( u0_K8_48 ) , .A( u0_R6_1 ) , .Z( u0_u7_X_48 ) );
  XOR2_X1 u0_u7_U8 (.B( u0_K8_47 ) , .A( u0_R6_32 ) , .Z( u0_u7_X_47 ) );
  XOR2_X1 u0_u7_U9 (.B( u0_K8_46 ) , .A( u0_R6_31 ) , .Z( u0_u7_X_46 ) );
  XOR2_X1 u0_u8_U1 (.B( u0_K9_9 ) , .A( u0_R7_6 ) , .Z( u0_u8_X_9 ) );
  XOR2_X1 u0_u8_U10 (.B( u0_K9_45 ) , .A( u0_R7_30 ) , .Z( u0_u8_X_45 ) );
  XOR2_X1 u0_u8_U15 (.B( u0_K9_40 ) , .A( u0_R7_27 ) , .Z( u0_u8_X_40 ) );
  XOR2_X1 u0_u8_U16 (.B( u0_K9_3 ) , .A( u0_R7_2 ) , .Z( u0_u8_X_3 ) );
  XOR2_X1 u0_u8_U17 (.B( u0_K9_39 ) , .A( u0_R7_26 ) , .Z( u0_u8_X_39 ) );
  XOR2_X1 u0_u8_U29 (.B( u0_K9_28 ) , .A( u0_R7_19 ) , .Z( u0_u8_X_28 ) );
  XOR2_X1 u0_u8_U30 (.B( u0_K9_27 ) , .A( u0_R7_18 ) , .Z( u0_u8_X_27 ) );
  XOR2_X1 u0_u8_U32 (.B( u0_K9_25 ) , .A( u0_R7_16 ) , .Z( u0_u8_X_25 ) );
  XOR2_X1 u0_u8_U34 (.B( u0_K9_23 ) , .A( u0_R7_16 ) , .Z( u0_u8_X_23 ) );
  XOR2_X1 u0_u8_U35 (.B( u0_K9_22 ) , .A( u0_R7_15 ) , .Z( u0_u8_X_22 ) );
  XOR2_X1 u0_u8_U37 (.B( u0_K9_20 ) , .A( u0_R7_13 ) , .Z( u0_u8_X_20 ) );
  XOR2_X1 u0_u8_U40 (.B( u0_K9_18 ) , .A( u0_R7_13 ) , .Z( u0_u8_X_18 ) );
  XOR2_X1 u0_u8_U42 (.B( u0_K9_16 ) , .A( u0_R7_11 ) , .Z( u0_u8_X_16 ) );
  XOR2_X1 u0_u8_U43 (.B( u0_K9_15 ) , .A( u0_R7_10 ) , .Z( u0_u8_X_15 ) );
  XOR2_X1 u0_u8_U48 (.B( u0_K9_10 ) , .A( u0_R7_7 ) , .Z( u0_u8_X_10 ) );
  XOR2_X1 u0_u8_U6 (.B( u0_K9_4 ) , .A( u0_R7_3 ) , .Z( u0_u8_X_4 ) );
  XOR2_X1 u0_u8_U9 (.B( u0_K9_46 ) , .A( u0_R7_31 ) , .Z( u0_u8_X_46 ) );
  XOR2_X1 u0_u9_U12 (.B( u0_K10_43 ) , .A( u0_R8_28 ) , .Z( u0_u9_X_43 ) );
  XOR2_X1 u0_u9_U14 (.B( u0_K10_41 ) , .A( u0_R8_28 ) , .Z( u0_u9_X_41 ) );
  XOR2_X1 u0_u9_U16 (.B( u0_K10_3 ) , .A( u0_R8_2 ) , .Z( u0_u9_X_3 ) );
  XOR2_X1 u0_u9_U17 (.B( u0_K10_39 ) , .A( u0_R8_26 ) , .Z( u0_u9_X_39 ) );
  XOR2_X1 u0_u9_U18 (.B( u0_K10_38 ) , .A( u0_R8_25 ) , .Z( u0_u9_X_38 ) );
  XOR2_X1 u0_u9_U19 (.B( u0_K10_37 ) , .A( u0_R8_24 ) , .Z( u0_u9_X_37 ) );
  XOR2_X1 u0_u9_U20 (.B( u0_K10_36 ) , .A( u0_R8_25 ) , .Z( u0_u9_X_36 ) );
  XOR2_X1 u0_u9_U21 (.B( u0_K10_35 ) , .A( u0_R8_24 ) , .Z( u0_u9_X_35 ) );
  XOR2_X1 u0_u9_U22 (.B( u0_K10_34 ) , .A( u0_R8_23 ) , .Z( u0_u9_X_34 ) );
  XOR2_X1 u0_u9_U3 (.B( u0_K10_7 ) , .A( u0_R8_4 ) , .Z( u0_u9_X_7 ) );
  XOR2_X1 u0_u9_U30 (.B( u0_K10_27 ) , .A( u0_R8_18 ) , .Z( u0_u9_X_27 ) );
  XOR2_X1 u0_u9_U32 (.B( u0_K10_25 ) , .A( u0_R8_16 ) , .Z( u0_u9_X_25 ) );
  XOR2_X1 u0_u9_U34 (.B( u0_K10_23 ) , .A( u0_R8_16 ) , .Z( u0_u9_X_23 ) );
  XOR2_X1 u0_u9_U35 (.B( u0_K10_22 ) , .A( u0_R8_15 ) , .Z( u0_u9_X_22 ) );
  XOR2_X1 u0_u9_U36 (.B( u0_K10_21 ) , .A( u0_R8_14 ) , .Z( u0_u9_X_21 ) );
  XOR2_X1 u0_u9_U42 (.B( u0_K10_16 ) , .A( u0_R8_11 ) , .Z( u0_u9_X_16 ) );
  XOR2_X1 u0_u9_U43 (.B( u0_K10_15 ) , .A( u0_R8_10 ) , .Z( u0_u9_X_15 ) );
  XOR2_X1 u0_u9_U45 (.B( u0_K10_13 ) , .A( u0_R8_8 ) , .Z( u0_u9_X_13 ) );
  XOR2_X1 u0_u9_U47 (.B( u0_K10_11 ) , .A( u0_R8_8 ) , .Z( u0_u9_X_11 ) );
  XOR2_X1 u0_u9_U48 (.B( u0_K10_10 ) , .A( u0_R8_7 ) , .Z( u0_u9_X_10 ) );
  XOR2_X1 u0_u9_U5 (.B( u0_K10_5 ) , .A( u0_R8_4 ) , .Z( u0_u9_X_5 ) );
  XOR2_X1 u0_u9_U6 (.B( u0_K10_4 ) , .A( u0_R8_3 ) , .Z( u0_u9_X_4 ) );
  XOR2_X1 u0_u9_U9 (.B( u0_K10_46 ) , .A( u0_R8_31 ) , .Z( u0_u9_X_46 ) );
  DFF_X1 u0_uk_K_r0_reg_0 (.CK( clk ) , .D( u0_key_r_0 ) , .Q( u0_uk_K_r0_0 ) , .QN( u0_uk_n628 ) );
  DFF_X1 u0_uk_K_r0_reg_1 (.CK( clk ) , .D( u0_key_r_1 ) , .Q( u0_uk_K_r0_1 ) );
  DFF_X1 u0_uk_K_r0_reg_10 (.CK( clk ) , .D( u0_key_r_10 ) , .Q( u0_uk_K_r0_10 ) , .QN( u0_uk_n620 ) );
  DFF_X1 u0_uk_K_r0_reg_11 (.CK( clk ) , .D( u0_key_r_11 ) , .Q( u0_uk_K_r0_11 ) );
  DFF_X1 u0_uk_K_r0_reg_12 (.CK( clk ) , .D( u0_key_r_12 ) , .Q( u0_uk_K_r0_12 ) , .QN( u0_uk_n619 ) );
  DFF_X1 u0_uk_K_r0_reg_13 (.CK( clk ) , .D( u0_key_r_13 ) , .Q( u0_uk_K_r0_13 ) , .QN( u0_uk_n618 ) );
  DFF_X1 u0_uk_K_r0_reg_14 (.CK( clk ) , .D( u0_key_r_14 ) , .Q( u0_uk_K_r0_14 ) , .QN( u0_uk_n617 ) );
  DFF_X1 u0_uk_K_r0_reg_15 (.CK( clk ) , .D( u0_key_r_15 ) , .Q( u0_uk_K_r0_15 ) );
  DFF_X1 u0_uk_K_r0_reg_16 (.CK( clk ) , .D( u0_key_r_16 ) , .Q( u0_uk_K_r0_16 ) , .QN( u0_uk_n616 ) );
  DFF_X1 u0_uk_K_r0_reg_17 (.CK( clk ) , .D( u0_key_r_17 ) , .Q( u0_uk_K_r0_17 ) );
  DFF_X1 u0_uk_K_r0_reg_18 (.CK( clk ) , .D( u0_key_r_18 ) , .Q( u0_uk_K_r0_18 ) , .QN( u0_uk_n615 ) );
  DFF_X1 u0_uk_K_r0_reg_19 (.CK( clk ) , .D( u0_key_r_19 ) , .Q( u0_uk_K_r0_19 ) );
  DFF_X1 u0_uk_K_r0_reg_2 (.CK( clk ) , .D( u0_key_r_2 ) , .Q( u0_uk_K_r0_2 ) );
  DFF_X1 u0_uk_K_r0_reg_20 (.CK( clk ) , .D( u0_key_r_20 ) , .Q( u0_uk_K_r0_20 ) , .QN( u0_uk_n614 ) );
  DFF_X1 u0_uk_K_r0_reg_21 (.CK( clk ) , .D( u0_key_r_21 ) , .Q( u0_uk_K_r0_21 ) , .QN( u0_uk_n613 ) );
  DFF_X1 u0_uk_K_r0_reg_22 (.CK( clk ) , .D( u0_key_r_22 ) , .Q( u0_uk_K_r0_22 ) );
  DFF_X1 u0_uk_K_r0_reg_23 (.CK( clk ) , .D( u0_key_r_23 ) , .Q( u0_uk_K_r0_23 ) , .QN( u0_uk_n612 ) );
  DFF_X1 u0_uk_K_r0_reg_24 (.CK( clk ) , .D( u0_key_r_24 ) , .Q( u0_uk_K_r0_24 ) , .QN( u0_uk_n611 ) );
  DFF_X1 u0_uk_K_r0_reg_25 (.CK( clk ) , .D( u0_key_r_25 ) , .Q( u0_uk_K_r0_25 ) );
  DFF_X1 u0_uk_K_r0_reg_26 (.CK( clk ) , .D( u0_key_r_26 ) , .Q( u0_uk_K_r0_26 ) , .QN( u0_uk_n610 ) );
  DFF_X1 u0_uk_K_r0_reg_27 (.CK( clk ) , .D( u0_key_r_27 ) , .Q( u0_uk_K_r0_27 ) , .QN( u0_uk_n609 ) );
  DFF_X1 u0_uk_K_r0_reg_28 (.CK( clk ) , .D( u0_key_r_28 ) , .Q( u0_uk_K_r0_28 ) );
  DFF_X1 u0_uk_K_r0_reg_29 (.CK( clk ) , .D( u0_key_r_29 ) , .Q( u0_uk_K_r0_29 ) , .QN( u0_uk_n607 ) );
  DFF_X1 u0_uk_K_r0_reg_3 (.CK( clk ) , .D( u0_key_r_3 ) , .Q( u0_uk_K_r0_3 ) , .QN( u0_uk_n627 ) );
  DFF_X1 u0_uk_K_r0_reg_30 (.CK( clk ) , .D( u0_key_r_30 ) , .Q( u0_uk_K_r0_30 ) , .QN( u0_uk_n606 ) );
  DFF_X1 u0_uk_K_r0_reg_31 (.CK( clk ) , .D( u0_key_r_31 ) , .Q( u0_uk_K_r0_31 ) );
  DFF_X1 u0_uk_K_r0_reg_32 (.CK( clk ) , .D( u0_key_r_32 ) , .Q( u0_uk_K_r0_32 ) );
  DFF_X1 u0_uk_K_r0_reg_33 (.CK( clk ) , .D( u0_key_r_33 ) , .Q( u0_uk_K_r0_33 ) , .QN( u0_uk_n604 ) );
  DFF_X1 u0_uk_K_r0_reg_34 (.CK( clk ) , .D( u0_key_r_34 ) , .Q( u0_uk_K_r0_34 ) );
  DFF_X1 u0_uk_K_r0_reg_35 (.CK( clk ) , .D( u0_key_r_35 ) , .Q( u0_uk_K_r0_35 ) , .QN( u0_uk_n602 ) );
  DFF_X1 u0_uk_K_r0_reg_36 (.CK( clk ) , .D( u0_key_r_36 ) , .Q( u0_uk_K_r0_36 ) );
  DFF_X1 u0_uk_K_r0_reg_37 (.CK( clk ) , .D( u0_key_r_37 ) , .Q( u0_uk_K_r0_37 ) , .QN( u0_uk_n600 ) );
  DFF_X1 u0_uk_K_r0_reg_38 (.CK( clk ) , .D( u0_key_r_38 ) , .Q( u0_uk_K_r0_38 ) , .QN( u0_uk_n599 ) );
  DFF_X1 u0_uk_K_r0_reg_39 (.CK( clk ) , .D( u0_key_r_39 ) , .Q( u0_uk_K_r0_39 ) , .QN( u0_uk_n598 ) );
  DFF_X1 u0_uk_K_r0_reg_4 (.CK( clk ) , .D( u0_key_r_4 ) , .Q( u0_uk_K_r0_4 ) , .QN( u0_uk_n626 ) );
  DFF_X1 u0_uk_K_r0_reg_40 (.CK( clk ) , .D( u0_key_r_40 ) , .Q( u0_uk_K_r0_40 ) , .QN( u0_uk_n597 ) );
  DFF_X1 u0_uk_K_r0_reg_41 (.CK( clk ) , .D( u0_key_r_41 ) , .Q( u0_uk_K_r0_41 ) , .QN( u0_uk_n596 ) );
  DFF_X1 u0_uk_K_r0_reg_42 (.CK( clk ) , .D( u0_key_r_42 ) , .Q( u0_uk_K_r0_42 ) , .QN( u0_uk_n595 ) );
  DFF_X1 u0_uk_K_r0_reg_43 (.CK( clk ) , .D( u0_key_r_43 ) , .Q( u0_uk_K_r0_43 ) , .QN( u0_uk_n594 ) );
  DFF_X1 u0_uk_K_r0_reg_44 (.CK( clk ) , .D( u0_key_r_44 ) , .Q( u0_uk_K_r0_44 ) , .QN( u0_uk_n593 ) );
  DFF_X1 u0_uk_K_r0_reg_45 (.CK( clk ) , .D( u0_key_r_45 ) , .Q( u0_uk_K_r0_45 ) , .QN( u0_uk_n592 ) );
  DFF_X1 u0_uk_K_r0_reg_46 (.CK( clk ) , .D( u0_key_r_46 ) , .Q( u0_uk_K_r0_46 ) , .QN( u0_uk_n591 ) );
  DFF_X1 u0_uk_K_r0_reg_47 (.CK( clk ) , .D( u0_key_r_47 ) , .Q( u0_uk_K_r0_47 ) , .QN( u0_uk_n589 ) );
  DFF_X1 u0_uk_K_r0_reg_48 (.CK( clk ) , .D( u0_key_r_48 ) , .Q( u0_uk_K_r0_48 ) , .QN( u0_uk_n588 ) );
  DFF_X1 u0_uk_K_r0_reg_49 (.CK( clk ) , .D( u0_key_r_49 ) , .Q( u0_uk_K_r0_49 ) );
  DFF_X1 u0_uk_K_r0_reg_5 (.CK( clk ) , .D( u0_key_r_5 ) , .Q( u0_uk_K_r0_5 ) , .QN( u0_uk_n625 ) );
  DFF_X1 u0_uk_K_r0_reg_50 (.CK( clk ) , .D( u0_key_r_50 ) , .Q( u0_uk_K_r0_50 ) , .QN( u0_uk_n585 ) );
  DFF_X1 u0_uk_K_r0_reg_51 (.CK( clk ) , .D( u0_key_r_51 ) , .Q( u0_uk_K_r0_51 ) , .QN( u0_uk_n584 ) );
  DFF_X1 u0_uk_K_r0_reg_52 (.CK( clk ) , .D( u0_key_r_52 ) , .Q( u0_uk_K_r0_52 ) );
  DFF_X1 u0_uk_K_r0_reg_53 (.CK( clk ) , .D( u0_key_r_53 ) , .Q( u0_uk_K_r0_53 ) );
  DFF_X1 u0_uk_K_r0_reg_54 (.CK( clk ) , .D( u0_key_r_54 ) , .Q( u0_uk_K_r0_54 ) , .QN( u0_uk_n583 ) );
  DFF_X1 u0_uk_K_r0_reg_55 (.CK( clk ) , .D( u0_key_r_55 ) , .Q( u0_uk_K_r0_55 ) );
  DFF_X1 u0_uk_K_r0_reg_6 (.CK( clk ) , .D( u0_key_r_6 ) , .Q( u0_uk_K_r0_6 ) , .QN( u0_uk_n624 ) );
  DFF_X1 u0_uk_K_r0_reg_7 (.CK( clk ) , .D( u0_key_r_7 ) , .Q( u0_uk_K_r0_7 ) , .QN( u0_uk_n623 ) );
  DFF_X1 u0_uk_K_r0_reg_8 (.CK( clk ) , .D( u0_key_r_8 ) , .Q( u0_uk_K_r0_8 ) , .QN( u0_uk_n622 ) );
  DFF_X1 u0_uk_K_r0_reg_9 (.CK( clk ) , .D( u0_key_r_9 ) , .Q( u0_uk_K_r0_9 ) , .QN( u0_uk_n621 ) );
  DFF_X1 u0_uk_K_r10_reg_0 (.CK( clk ) , .Q( u0_uk_K_r10_0 ) , .D( u0_uk_K_r9_0 ) , .QN( u0_uk_n180 ) );
  DFF_X1 u0_uk_K_r10_reg_1 (.CK( clk ) , .Q( u0_uk_K_r10_1 ) , .D( u0_uk_K_r9_1 ) , .QN( u0_uk_n179 ) );
  DFF_X1 u0_uk_K_r10_reg_10 (.CK( clk ) , .Q( u0_uk_K_r10_10 ) , .D( u0_uk_K_r9_10 ) );
  DFF_X1 u0_uk_K_r10_reg_11 (.CK( clk ) , .Q( u0_uk_K_r10_11 ) , .D( u0_uk_K_r9_11 ) );
  DFF_X1 u0_uk_K_r10_reg_12 (.CK( clk ) , .Q( u0_uk_K_r10_12 ) , .D( u0_uk_K_r9_12 ) , .QN( u0_uk_n172 ) );
  DFF_X1 u0_uk_K_r10_reg_13 (.CK( clk ) , .Q( u0_uk_K_r10_13 ) , .D( u0_uk_K_r9_13 ) );
  DFF_X1 u0_uk_K_r10_reg_14 (.CK( clk ) , .Q( u0_uk_K_r10_14 ) , .D( u0_uk_K_r9_14 ) );
  DFF_X1 u0_uk_K_r10_reg_15 (.CK( clk ) , .Q( u0_uk_K_r10_15 ) , .D( u0_uk_K_r9_15 ) , .QN( u0_uk_n171 ) );
  DFF_X1 u0_uk_K_r10_reg_16 (.CK( clk ) , .Q( u0_uk_K_r10_16 ) , .D( u0_uk_K_r9_16 ) );
  DFF_X1 u0_uk_K_r10_reg_17 (.CK( clk ) , .Q( u0_uk_K_r10_17 ) , .D( u0_uk_K_r9_17 ) , .QN( u0_uk_n170 ) );
  DFF_X1 u0_uk_K_r10_reg_18 (.CK( clk ) , .Q( u0_uk_K_r10_18 ) , .D( u0_uk_K_r9_18 ) );
  DFF_X1 u0_uk_K_r10_reg_19 (.CK( clk ) , .Q( u0_uk_K_r10_19 ) , .D( u0_uk_K_r9_19 ) );
  DFF_X1 u0_uk_K_r10_reg_2 (.CK( clk ) , .Q( u0_uk_K_r10_2 ) , .D( u0_uk_K_r9_2 ) , .QN( u0_uk_n178 ) );
  DFF_X1 u0_uk_K_r10_reg_20 (.CK( clk ) , .Q( u0_uk_K_r10_20 ) , .D( u0_uk_K_r9_20 ) , .QN( u0_uk_n169 ) );
  DFF_X1 u0_uk_K_r10_reg_21 (.CK( clk ) , .Q( u0_uk_K_r10_21 ) , .D( u0_uk_K_r9_21 ) , .QN( u0_uk_n168 ) );
  DFF_X1 u0_uk_K_r10_reg_22 (.CK( clk ) , .Q( u0_uk_K_r10_22 ) , .D( u0_uk_K_r9_22 ) , .QN( u0_uk_n167 ) );
  DFF_X1 u0_uk_K_r10_reg_23 (.CK( clk ) , .Q( u0_uk_K_r10_23 ) , .D( u0_uk_K_r9_23 ) );
  DFF_X1 u0_uk_K_r10_reg_24 (.CK( clk ) , .Q( u0_uk_K_r10_24 ) , .D( u0_uk_K_r9_24 ) , .QN( u0_uk_n166 ) );
  DFF_X1 u0_uk_K_r10_reg_25 (.CK( clk ) , .Q( u0_uk_K_r10_25 ) , .D( u0_uk_K_r9_25 ) );
  DFF_X1 u0_uk_K_r10_reg_26 (.CK( clk ) , .Q( u0_uk_K_r10_26 ) , .D( u0_uk_K_r9_26 ) , .QN( u0_uk_n165 ) );
  DFF_X1 u0_uk_K_r10_reg_27 (.CK( clk ) , .Q( u0_uk_K_r10_27 ) , .D( u0_uk_K_r9_27 ) );
  DFF_X1 u0_uk_K_r10_reg_28 (.CK( clk ) , .Q( u0_uk_K_r10_28 ) , .D( u0_uk_K_r9_28 ) );
  DFF_X1 u0_uk_K_r10_reg_29 (.CK( clk ) , .Q( u0_uk_K_r10_29 ) , .D( u0_uk_K_r9_29 ) , .QN( u0_uk_n160 ) );
  DFF_X1 u0_uk_K_r10_reg_3 (.CK( clk ) , .Q( u0_uk_K_r10_3 ) , .D( u0_uk_K_r9_3 ) , .QN( u0_uk_n177 ) );
  DFF_X1 u0_uk_K_r10_reg_30 (.CK( clk ) , .Q( u0_uk_K_r10_30 ) , .D( u0_uk_K_r9_30 ) , .QN( u0_uk_n159 ) );
  DFF_X1 u0_uk_K_r10_reg_31 (.CK( clk ) , .Q( u0_uk_K_r10_31 ) , .D( u0_uk_K_r9_31 ) , .QN( u0_uk_n158 ) );
  DFF_X1 u0_uk_K_r10_reg_32 (.CK( clk ) , .Q( u0_uk_K_r10_32 ) , .D( u0_uk_K_r9_32 ) , .QN( u0_uk_n157 ) );
  DFF_X1 u0_uk_K_r10_reg_33 (.CK( clk ) , .Q( u0_uk_K_r10_33 ) , .D( u0_uk_K_r9_33 ) , .QN( u0_uk_n156 ) );
  DFF_X1 u0_uk_K_r10_reg_34 (.CK( clk ) , .Q( u0_uk_K_r10_34 ) , .D( u0_uk_K_r9_34 ) );
  DFF_X1 u0_uk_K_r10_reg_35 (.CK( clk ) , .Q( u0_uk_K_r10_35 ) , .D( u0_uk_K_r9_35 ) , .QN( u0_uk_n154 ) );
  DFF_X1 u0_uk_K_r10_reg_36 (.CK( clk ) , .Q( u0_uk_K_r10_36 ) , .D( u0_uk_K_r9_36 ) , .QN( u0_uk_n153 ) );
  DFF_X1 u0_uk_K_r10_reg_37 (.CK( clk ) , .Q( u0_uk_K_r10_37 ) , .D( u0_uk_K_r9_37 ) , .QN( u0_uk_n152 ) );
  DFF_X1 u0_uk_K_r10_reg_38 (.CK( clk ) , .Q( u0_uk_K_r10_38 ) , .D( u0_uk_K_r9_38 ) , .QN( u0_uk_n151 ) );
  DFF_X1 u0_uk_K_r10_reg_39 (.CK( clk ) , .Q( u0_uk_K_r10_39 ) , .D( u0_uk_K_r9_39 ) , .QN( u0_uk_n150 ) );
  DFF_X1 u0_uk_K_r10_reg_4 (.CK( clk ) , .Q( u0_uk_K_r10_4 ) , .D( u0_uk_K_r9_4 ) );
  DFF_X1 u0_uk_K_r10_reg_40 (.CK( clk ) , .Q( u0_uk_K_r10_40 ) , .D( u0_uk_K_r9_40 ) , .QN( u0_uk_n149 ) );
  DFF_X1 u0_uk_K_r10_reg_41 (.CK( clk ) , .Q( u0_uk_K_r10_41 ) , .D( u0_uk_K_r9_41 ) );
  DFF_X1 u0_uk_K_r10_reg_42 (.CK( clk ) , .Q( u0_uk_K_r10_42 ) , .D( u0_uk_K_r9_42 ) );
  DFF_X1 u0_uk_K_r10_reg_43 (.CK( clk ) , .Q( u0_uk_K_r10_43 ) , .D( u0_uk_K_r9_43 ) );
  DFF_X1 u0_uk_K_r10_reg_44 (.CK( clk ) , .Q( u0_uk_K_r10_44 ) , .D( u0_uk_K_r9_44 ) );
  DFF_X1 u0_uk_K_r10_reg_45 (.CK( clk ) , .Q( u0_uk_K_r10_45 ) , .D( u0_uk_K_r9_45 ) , .QN( u0_uk_n144 ) );
  DFF_X1 u0_uk_K_r10_reg_46 (.CK( clk ) , .Q( u0_uk_K_r10_46 ) , .D( u0_uk_K_r9_46 ) , .QN( u0_uk_n143 ) );
  DFF_X1 u0_uk_K_r10_reg_47 (.CK( clk ) , .Q( u0_uk_K_r10_47 ) , .D( u0_uk_K_r9_47 ) );
  DFF_X1 u0_uk_K_r10_reg_48 (.CK( clk ) , .Q( u0_uk_K_r10_48 ) , .D( u0_uk_K_r9_48 ) );
  DFF_X1 u0_uk_K_r10_reg_49 (.CK( clk ) , .Q( u0_uk_K_r10_49 ) , .D( u0_uk_K_r9_49 ) );
  DFF_X1 u0_uk_K_r10_reg_5 (.CK( clk ) , .Q( u0_uk_K_r10_5 ) , .D( u0_uk_K_r9_5 ) , .QN( u0_uk_n176 ) );
  DFF_X1 u0_uk_K_r10_reg_50 (.CK( clk ) , .Q( u0_uk_K_r10_50 ) , .D( u0_uk_K_r9_50 ) , .QN( u0_uk_n140 ) );
  DFF_X1 u0_uk_K_r10_reg_51 (.CK( clk ) , .Q( u0_uk_K_r10_51 ) , .D( u0_uk_K_r9_51 ) , .QN( u0_uk_n139 ) );
  DFF_X1 u0_uk_K_r10_reg_52 (.CK( clk ) , .Q( u0_uk_K_r10_52 ) , .D( u0_uk_K_r9_52 ) );
  DFF_X1 u0_uk_K_r10_reg_53 (.CK( clk ) , .Q( u0_uk_K_r10_53 ) , .D( u0_uk_K_r9_53 ) , .QN( u0_uk_n138 ) );
  DFF_X1 u0_uk_K_r10_reg_54 (.CK( clk ) , .Q( u0_uk_K_r10_54 ) , .D( u0_uk_K_r9_54 ) , .QN( u0_uk_n137 ) );
  DFF_X1 u0_uk_K_r10_reg_55 (.CK( clk ) , .Q( u0_uk_K_r10_55 ) , .D( u0_uk_K_r9_55 ) , .QN( u0_uk_n136 ) );
  DFF_X1 u0_uk_K_r10_reg_6 (.CK( clk ) , .Q( u0_uk_K_r10_6 ) , .D( u0_uk_K_r9_6 ) , .QN( u0_uk_n175 ) );
  DFF_X1 u0_uk_K_r10_reg_7 (.CK( clk ) , .Q( u0_uk_K_r10_7 ) , .D( u0_uk_K_r9_7 ) , .QN( u0_uk_n174 ) );
  DFF_X1 u0_uk_K_r10_reg_8 (.CK( clk ) , .Q( u0_uk_K_r10_8 ) , .D( u0_uk_K_r9_8 ) , .QN( u0_uk_n173 ) );
  DFF_X1 u0_uk_K_r10_reg_9 (.CK( clk ) , .Q( u0_uk_K_r10_9 ) , .D( u0_uk_K_r9_9 ) );
  DFF_X1 u0_uk_K_r11_reg_0 (.CK( clk ) , .D( u0_uk_K_r10_0 ) , .Q( u0_uk_K_r11_0 ) , .QN( u0_uk_n135 ) );
  DFF_X1 u0_uk_K_r11_reg_1 (.CK( clk ) , .D( u0_uk_K_r10_1 ) , .Q( u0_uk_K_r11_1 ) , .QN( u0_uk_n134 ) );
  DFF_X1 u0_uk_K_r11_reg_10 (.CK( clk ) , .D( u0_uk_K_r10_10 ) , .Q( u0_uk_K_r11_10 ) );
  DFF_X1 u0_uk_K_r11_reg_11 (.CK( clk ) , .D( u0_uk_K_r10_11 ) , .Q( u0_uk_K_r11_11 ) );
  DFF_X1 u0_uk_K_r11_reg_12 (.CK( clk ) , .D( u0_uk_K_r10_12 ) , .Q( u0_uk_K_r11_12 ) , .QN( u0_uk_n127 ) );
  DFF_X1 u0_uk_K_r11_reg_13 (.CK( clk ) , .D( u0_uk_K_r10_13 ) , .Q( u0_uk_K_r11_13 ) , .QN( u0_uk_n126 ) );
  DFF_X1 u0_uk_K_r11_reg_14 (.CK( clk ) , .D( u0_uk_K_r10_14 ) , .Q( u0_uk_K_r11_14 ) , .QN( u0_uk_n125 ) );
  DFF_X1 u0_uk_K_r11_reg_15 (.CK( clk ) , .D( u0_uk_K_r10_15 ) , .Q( u0_uk_K_r11_15 ) , .QN( u0_uk_n124 ) );
  DFF_X1 u0_uk_K_r11_reg_16 (.CK( clk ) , .D( u0_uk_K_r10_16 ) , .Q( u0_uk_K_r11_16 ) , .QN( u0_uk_n123 ) );
  DFF_X1 u0_uk_K_r11_reg_17 (.CK( clk ) , .D( u0_uk_K_r10_17 ) , .Q( u0_uk_K_r11_17 ) , .QN( u0_uk_n122 ) );
  DFF_X1 u0_uk_K_r11_reg_18 (.CK( clk ) , .D( u0_uk_K_r10_18 ) , .Q( u0_uk_K_r11_18 ) , .QN( u0_uk_n121 ) );
  DFF_X1 u0_uk_K_r11_reg_19 (.CK( clk ) , .D( u0_uk_K_r10_19 ) , .Q( u0_uk_K_r11_19 ) );
  DFF_X1 u0_uk_K_r11_reg_2 (.CK( clk ) , .D( u0_uk_K_r10_2 ) , .Q( u0_uk_K_r11_2 ) , .QN( u0_uk_n133 ) );
  DFF_X1 u0_uk_K_r11_reg_20 (.CK( clk ) , .D( u0_uk_K_r10_20 ) , .Q( u0_uk_K_r11_20 ) );
  DFF_X1 u0_uk_K_r11_reg_21 (.CK( clk ) , .D( u0_uk_K_r10_21 ) , .Q( u0_uk_K_r11_21 ) );
  DFF_X1 u0_uk_K_r11_reg_22 (.CK( clk ) , .D( u0_uk_K_r10_22 ) , .Q( u0_uk_K_r11_22 ) , .QN( u0_uk_n120 ) );
  DFF_X1 u0_uk_K_r11_reg_23 (.CK( clk ) , .D( u0_uk_K_r10_23 ) , .Q( u0_uk_K_r11_23 ) , .QN( u0_uk_n119 ) );
  DFF_X1 u0_uk_K_r11_reg_24 (.CK( clk ) , .D( u0_uk_K_r10_24 ) , .Q( u0_uk_K_r11_24 ) );
  DFF_X1 u0_uk_K_r11_reg_25 (.CK( clk ) , .D( u0_uk_K_r10_25 ) , .Q( u0_uk_K_r11_25 ) );
  DFF_X1 u0_uk_K_r11_reg_26 (.CK( clk ) , .D( u0_uk_K_r10_26 ) , .Q( u0_uk_K_r11_26 ) );
  DFF_X1 u0_uk_K_r11_reg_27 (.CK( clk ) , .D( u0_uk_K_r10_27 ) , .Q( u0_uk_K_r11_27 ) );
  DFF_X1 u0_uk_K_r11_reg_28 (.CK( clk ) , .D( u0_uk_K_r10_28 ) , .Q( u0_uk_K_r11_28 ) );
  DFF_X1 u0_uk_K_r11_reg_29 (.CK( clk ) , .D( u0_uk_K_r10_29 ) , .Q( u0_uk_K_r11_29 ) );
  DFF_X1 u0_uk_K_r11_reg_3 (.CK( clk ) , .D( u0_uk_K_r10_3 ) , .Q( u0_uk_K_r11_3 ) , .QN( u0_uk_n132 ) );
  DFF_X1 u0_uk_K_r11_reg_30 (.CK( clk ) , .D( u0_uk_K_r10_30 ) , .Q( u0_uk_K_r11_30 ) );
  DFF_X1 u0_uk_K_r11_reg_31 (.CK( clk ) , .D( u0_uk_K_r10_31 ) , .Q( u0_uk_K_r11_31 ) , .QN( u0_uk_n116 ) );
  DFF_X1 u0_uk_K_r11_reg_32 (.CK( clk ) , .D( u0_uk_K_r10_32 ) , .Q( u0_uk_K_r11_32 ) , .QN( u0_uk_n115 ) );
  DFF_X1 u0_uk_K_r11_reg_33 (.CK( clk ) , .D( u0_uk_K_r10_33 ) , .Q( u0_uk_K_r11_33 ) );
  DFF_X1 u0_uk_K_r11_reg_34 (.CK( clk ) , .D( u0_uk_K_r10_34 ) , .Q( u0_uk_K_r11_34 ) );
  DFF_X1 u0_uk_K_r11_reg_35 (.CK( clk ) , .D( u0_uk_K_r10_35 ) , .Q( u0_uk_K_r11_35 ) , .QN( u0_uk_n114 ) );
  DFF_X1 u0_uk_K_r11_reg_36 (.CK( clk ) , .D( u0_uk_K_r10_36 ) , .Q( u0_uk_K_r11_36 ) , .QN( u0_uk_n113 ) );
  DFF_X1 u0_uk_K_r11_reg_37 (.CK( clk ) , .D( u0_uk_K_r10_37 ) , .Q( u0_uk_K_r11_37 ) , .QN( u0_uk_n112 ) );
  DFF_X1 u0_uk_K_r11_reg_38 (.CK( clk ) , .D( u0_uk_K_r10_38 ) , .Q( u0_uk_K_r11_38 ) , .QN( u0_uk_n111 ) );
  DFF_X1 u0_uk_K_r11_reg_39 (.CK( clk ) , .D( u0_uk_K_r10_39 ) , .Q( u0_uk_K_r11_39 ) );
  DFF_X1 u0_uk_K_r11_reg_4 (.CK( clk ) , .D( u0_uk_K_r10_4 ) , .Q( u0_uk_K_r11_4 ) );
  DFF_X1 u0_uk_K_r11_reg_40 (.CK( clk ) , .D( u0_uk_K_r10_40 ) , .Q( u0_uk_K_r11_40 ) , .QN( u0_uk_n108 ) );
  DFF_X1 u0_uk_K_r11_reg_41 (.CK( clk ) , .D( u0_uk_K_r10_41 ) , .Q( u0_uk_K_r11_41 ) , .QN( u0_uk_n107 ) );
  DFF_X1 u0_uk_K_r11_reg_42 (.CK( clk ) , .D( u0_uk_K_r10_42 ) , .Q( u0_uk_K_r11_42 ) , .QN( u0_uk_n106 ) );
  DFF_X1 u0_uk_K_r11_reg_43 (.CK( clk ) , .D( u0_uk_K_r10_43 ) , .Q( u0_uk_K_r11_43 ) , .QN( u0_uk_n105 ) );
  DFF_X1 u0_uk_K_r11_reg_44 (.CK( clk ) , .D( u0_uk_K_r10_44 ) , .Q( u0_uk_K_r11_44 ) , .QN( u0_uk_n104 ) );
  DFF_X1 u0_uk_K_r11_reg_45 (.CK( clk ) , .D( u0_uk_K_r10_45 ) , .Q( u0_uk_K_r11_45 ) , .QN( u0_uk_n103 ) );
  DFF_X1 u0_uk_K_r11_reg_46 (.CK( clk ) , .D( u0_uk_K_r10_46 ) , .Q( u0_uk_K_r11_46 ) , .QN( u0_uk_n101 ) );
  DFF_X1 u0_uk_K_r11_reg_47 (.CK( clk ) , .D( u0_uk_K_r10_47 ) , .Q( u0_uk_K_r11_47 ) );
  DFF_X1 u0_uk_K_r11_reg_48 (.CK( clk ) , .D( u0_uk_K_r10_48 ) , .Q( u0_uk_K_r11_48 ) );
  DFF_X1 u0_uk_K_r11_reg_49 (.CK( clk ) , .D( u0_uk_K_r10_49 ) , .Q( u0_uk_K_r11_49 ) , .QN( u0_uk_n98 ) );
  DFF_X1 u0_uk_K_r11_reg_5 (.CK( clk ) , .D( u0_uk_K_r10_5 ) , .Q( u0_uk_K_r11_5 ) , .QN( u0_uk_n131 ) );
  DFF_X1 u0_uk_K_r11_reg_50 (.CK( clk ) , .D( u0_uk_K_r10_50 ) , .Q( u0_uk_K_r11_50 ) , .QN( u0_uk_n97 ) );
  DFF_X1 u0_uk_K_r11_reg_51 (.CK( clk ) , .D( u0_uk_K_r10_51 ) , .Q( u0_uk_K_r11_51 ) , .QN( u0_uk_n96 ) );
  DFF_X1 u0_uk_K_r11_reg_52 (.CK( clk ) , .D( u0_uk_K_r10_52 ) , .Q( u0_uk_K_r11_52 ) , .QN( u0_uk_n95 ) );
  DFF_X1 u0_uk_K_r11_reg_53 (.CK( clk ) , .D( u0_uk_K_r10_53 ) , .Q( u0_uk_K_r11_53 ) );
  DFF_X1 u0_uk_K_r11_reg_54 (.CK( clk ) , .D( u0_uk_K_r10_54 ) , .Q( u0_uk_K_r11_54 ) );
  DFF_X1 u0_uk_K_r11_reg_55 (.CK( clk ) , .D( u0_uk_K_r10_55 ) , .Q( u0_uk_K_r11_55 ) , .QN( u0_uk_n91 ) );
  DFF_X1 u0_uk_K_r11_reg_6 (.CK( clk ) , .D( u0_uk_K_r10_6 ) , .Q( u0_uk_K_r11_6 ) );
  DFF_X1 u0_uk_K_r11_reg_7 (.CK( clk ) , .D( u0_uk_K_r10_7 ) , .Q( u0_uk_K_r11_7 ) );
  DFF_X1 u0_uk_K_r11_reg_8 (.CK( clk ) , .D( u0_uk_K_r10_8 ) , .Q( u0_uk_K_r11_8 ) );
  DFF_X1 u0_uk_K_r11_reg_9 (.CK( clk ) , .D( u0_uk_K_r10_9 ) , .Q( u0_uk_K_r11_9 ) , .QN( u0_uk_n130 ) );
  DFF_X1 u0_uk_K_r12_reg_0 (.CK( clk ) , .D( u0_uk_K_r11_0 ) , .Q( u0_uk_K_r12_0 ) , .QN( u0_uk_n90 ) );
  DFF_X1 u0_uk_K_r12_reg_1 (.CK( clk ) , .D( u0_uk_K_r11_1 ) , .Q( u0_uk_K_r12_1 ) , .QN( u0_uk_n89 ) );
  DFF_X1 u0_uk_K_r12_reg_10 (.CK( clk ) , .D( u0_uk_K_r11_10 ) , .Q( u0_uk_K_r12_10 ) );
  DFF_X1 u0_uk_K_r12_reg_11 (.CK( clk ) , .D( u0_uk_K_r11_11 ) , .Q( u0_uk_K_r12_11 ) , .QN( u0_uk_n80 ) );
  DFF_X1 u0_uk_K_r12_reg_12 (.CK( clk ) , .D( u0_uk_K_r11_12 ) , .Q( u0_uk_K_r12_12 ) , .QN( u0_uk_n79 ) );
  DFF_X1 u0_uk_K_r12_reg_13 (.CK( clk ) , .D( u0_uk_K_r11_13 ) , .Q( u0_uk_K_r12_13 ) , .QN( u0_uk_n78 ) );
  DFF_X1 u0_uk_K_r12_reg_14 (.CK( clk ) , .D( u0_uk_K_r11_14 ) , .Q( u0_uk_K_r12_14 ) , .QN( u0_uk_n77 ) );
  DFF_X1 u0_uk_K_r12_reg_15 (.CK( clk ) , .D( u0_uk_K_r11_15 ) , .Q( u0_uk_K_r12_15 ) );
  DFF_X1 u0_uk_K_r12_reg_16 (.CK( clk ) , .D( u0_uk_K_r11_16 ) , .Q( u0_uk_K_r12_16 ) );
  DFF_X1 u0_uk_K_r12_reg_17 (.CK( clk ) , .D( u0_uk_K_r11_17 ) , .Q( u0_uk_K_r12_17 ) , .QN( u0_uk_n76 ) );
  DFF_X1 u0_uk_K_r12_reg_18 (.CK( clk ) , .D( u0_uk_K_r11_18 ) , .Q( u0_uk_K_r12_18 ) );
  DFF_X1 u0_uk_K_r12_reg_19 (.CK( clk ) , .D( u0_uk_K_r11_19 ) , .Q( u0_uk_K_r12_19 ) , .QN( u0_uk_n75 ) );
  DFF_X1 u0_uk_K_r12_reg_2 (.CK( clk ) , .D( u0_uk_K_r11_2 ) , .Q( u0_uk_K_r12_2 ) , .QN( u0_uk_n88 ) );
  DFF_X1 u0_uk_K_r12_reg_20 (.CK( clk ) , .D( u0_uk_K_r11_20 ) , .Q( u0_uk_K_r12_20 ) , .QN( u0_uk_n74 ) );
  DFF_X1 u0_uk_K_r12_reg_21 (.CK( clk ) , .D( u0_uk_K_r11_21 ) , .Q( u0_uk_K_r12_21 ) );
  DFF_X1 u0_uk_K_r12_reg_22 (.CK( clk ) , .D( u0_uk_K_r11_22 ) , .Q( u0_uk_K_r12_22 ) );
  DFF_X1 u0_uk_K_r12_reg_23 (.CK( clk ) , .D( u0_uk_K_r11_23 ) , .Q( u0_uk_K_r12_23 ) , .QN( u0_uk_n73 ) );
  DFF_X1 u0_uk_K_r12_reg_24 (.CK( clk ) , .D( u0_uk_K_r11_24 ) , .Q( u0_uk_K_r12_24 ) , .QN( u0_uk_n72 ) );
  DFF_X1 u0_uk_K_r12_reg_25 (.CK( clk ) , .D( u0_uk_K_r11_25 ) , .Q( u0_uk_K_r12_25 ) , .QN( u0_uk_n71 ) );
  DFF_X1 u0_uk_K_r12_reg_26 (.CK( clk ) , .D( u0_uk_K_r11_26 ) , .Q( u0_uk_K_r12_26 ) , .QN( u0_uk_n70 ) );
  DFF_X1 u0_uk_K_r12_reg_27 (.CK( clk ) , .D( u0_uk_K_r11_27 ) , .Q( u0_uk_K_r12_27 ) , .QN( u0_uk_n69 ) );
  DFF_X1 u0_uk_K_r12_reg_28 (.CK( clk ) , .D( u0_uk_K_r11_28 ) , .Q( u0_uk_K_r12_28 ) , .QN( u0_uk_n68 ) );
  DFF_X1 u0_uk_K_r12_reg_29 (.CK( clk ) , .D( u0_uk_K_r11_29 ) , .Q( u0_uk_K_r12_29 ) , .QN( u0_uk_n67 ) );
  DFF_X1 u0_uk_K_r12_reg_3 (.CK( clk ) , .D( u0_uk_K_r11_3 ) , .Q( u0_uk_K_r12_3 ) , .QN( u0_uk_n87 ) );
  DFF_X1 u0_uk_K_r12_reg_30 (.CK( clk ) , .D( u0_uk_K_r11_30 ) , .Q( u0_uk_K_r12_30 ) , .QN( u0_uk_n66 ) );
  DFF_X1 u0_uk_K_r12_reg_31 (.CK( clk ) , .D( u0_uk_K_r11_31 ) , .Q( u0_uk_K_r12_31 ) , .QN( u0_uk_n65 ) );
  DFF_X1 u0_uk_K_r12_reg_32 (.CK( clk ) , .D( u0_uk_K_r11_32 ) , .Q( u0_uk_K_r12_32 ) , .QN( u0_uk_n64 ) );
  DFF_X1 u0_uk_K_r12_reg_33 (.CK( clk ) , .D( u0_uk_K_r11_33 ) , .Q( u0_uk_K_r12_33 ) );
  DFF_X1 u0_uk_K_r12_reg_34 (.CK( clk ) , .D( u0_uk_K_r11_34 ) , .Q( u0_uk_K_r12_34 ) , .QN( u0_uk_n62 ) );
  DFF_X1 u0_uk_K_r12_reg_35 (.CK( clk ) , .D( u0_uk_K_r11_35 ) , .Q( u0_uk_K_r12_35 ) , .QN( u0_uk_n61 ) );
  DFF_X1 u0_uk_K_r12_reg_36 (.CK( clk ) , .D( u0_uk_K_r11_36 ) , .Q( u0_uk_K_r12_36 ) );
  DFF_X1 u0_uk_K_r12_reg_37 (.CK( clk ) , .D( u0_uk_K_r11_37 ) , .Q( u0_uk_K_r12_37 ) , .QN( u0_uk_n59 ) );
  DFF_X1 u0_uk_K_r12_reg_38 (.CK( clk ) , .D( u0_uk_K_r11_38 ) , .Q( u0_uk_K_r12_38 ) , .QN( u0_uk_n58 ) );
  DFF_X1 u0_uk_K_r12_reg_39 (.CK( clk ) , .D( u0_uk_K_r11_39 ) , .Q( u0_uk_K_r12_39 ) );
  DFF_X1 u0_uk_K_r12_reg_4 (.CK( clk ) , .D( u0_uk_K_r11_4 ) , .Q( u0_uk_K_r12_4 ) , .QN( u0_uk_n86 ) );
  DFF_X1 u0_uk_K_r12_reg_40 (.CK( clk ) , .D( u0_uk_K_r11_40 ) , .Q( u0_uk_K_r12_40 ) , .QN( u0_uk_n57 ) );
  DFF_X1 u0_uk_K_r12_reg_41 (.CK( clk ) , .D( u0_uk_K_r11_41 ) , .Q( u0_uk_K_r12_41 ) );
  DFF_X1 u0_uk_K_r12_reg_42 (.CK( clk ) , .D( u0_uk_K_r11_42 ) , .Q( u0_uk_K_r12_42 ) );
  DFF_X1 u0_uk_K_r12_reg_43 (.CK( clk ) , .D( u0_uk_K_r11_43 ) , .Q( u0_uk_K_r12_43 ) , .QN( u0_uk_n56 ) );
  DFF_X1 u0_uk_K_r12_reg_44 (.CK( clk ) , .D( u0_uk_K_r11_44 ) , .Q( u0_uk_K_r12_44 ) );
  DFF_X1 u0_uk_K_r12_reg_45 (.CK( clk ) , .D( u0_uk_K_r11_45 ) , .Q( u0_uk_K_r12_45 ) , .QN( u0_uk_n55 ) );
  DFF_X1 u0_uk_K_r12_reg_46 (.CK( clk ) , .D( u0_uk_K_r11_46 ) , .Q( u0_uk_K_r12_46 ) , .QN( u0_uk_n54 ) );
  DFF_X1 u0_uk_K_r12_reg_47 (.CK( clk ) , .D( u0_uk_K_r11_47 ) , .Q( u0_uk_K_r12_47 ) );
  DFF_X1 u0_uk_K_r12_reg_48 (.CK( clk ) , .D( u0_uk_K_r11_48 ) , .Q( u0_uk_K_r12_48 ) , .QN( u0_uk_n53 ) );
  DFF_X1 u0_uk_K_r12_reg_49 (.CK( clk ) , .D( u0_uk_K_r11_49 ) , .Q( u0_uk_K_r12_49 ) , .QN( u0_uk_n52 ) );
  DFF_X1 u0_uk_K_r12_reg_5 (.CK( clk ) , .D( u0_uk_K_r11_5 ) , .Q( u0_uk_K_r12_5 ) , .QN( u0_uk_n85 ) );
  DFF_X1 u0_uk_K_r12_reg_50 (.CK( clk ) , .D( u0_uk_K_r11_50 ) , .Q( u0_uk_K_r12_50 ) , .QN( u0_uk_n51 ) );
  DFF_X1 u0_uk_K_r12_reg_51 (.CK( clk ) , .D( u0_uk_K_r11_51 ) , .Q( u0_uk_K_r12_51 ) , .QN( u0_uk_n50 ) );
  DFF_X1 u0_uk_K_r12_reg_52 (.CK( clk ) , .D( u0_uk_K_r11_52 ) , .Q( u0_uk_K_r12_52 ) , .QN( u0_uk_n49 ) );
  DFF_X1 u0_uk_K_r12_reg_53 (.CK( clk ) , .D( u0_uk_K_r11_53 ) , .Q( u0_uk_K_r12_53 ) , .QN( u0_uk_n48 ) );
  DFF_X1 u0_uk_K_r12_reg_54 (.CK( clk ) , .D( u0_uk_K_r11_54 ) , .Q( u0_uk_K_r12_54 ) , .QN( u0_uk_n47 ) );
  DFF_X1 u0_uk_K_r12_reg_55 (.CK( clk ) , .D( u0_uk_K_r11_55 ) , .Q( u0_uk_K_r12_55 ) , .QN( u0_uk_n46 ) );
  DFF_X1 u0_uk_K_r12_reg_6 (.CK( clk ) , .D( u0_uk_K_r11_6 ) , .Q( u0_uk_K_r12_6 ) , .QN( u0_uk_n84 ) );
  DFF_X1 u0_uk_K_r12_reg_7 (.CK( clk ) , .D( u0_uk_K_r11_7 ) , .Q( u0_uk_K_r12_7 ) );
  DFF_X1 u0_uk_K_r12_reg_8 (.CK( clk ) , .D( u0_uk_K_r11_8 ) , .Q( u0_uk_K_r12_8 ) , .QN( u0_uk_n82 ) );
  DFF_X1 u0_uk_K_r12_reg_9 (.CK( clk ) , .D( u0_uk_K_r11_9 ) , .Q( u0_uk_K_r12_9 ) , .QN( u0_uk_n81 ) );
  DFF_X1 u0_uk_K_r13_reg_0 (.CK( clk ) , .D( u0_uk_K_r12_0 ) , .Q( u0_uk_K_r13_0 ) , .QN( u0_uk_n45 ) );
  DFF_X1 u0_uk_K_r13_reg_1 (.CK( clk ) , .D( u0_uk_K_r12_1 ) , .Q( u0_uk_K_r13_1 ) );
  DFF_X1 u0_uk_K_r13_reg_10 (.CK( clk ) , .D( u0_uk_K_r12_10 ) , .Q( u0_uk_K_r13_10 ) , .QN( u0_uk_n38 ) );
  DFF_X1 u0_uk_K_r13_reg_11 (.CK( clk ) , .D( u0_uk_K_r12_11 ) , .Q( u0_uk_K_r13_11 ) , .QN( u0_uk_n37 ) );
  DFF_X1 u0_uk_K_r13_reg_12 (.CK( clk ) , .D( u0_uk_K_r12_12 ) , .Q( u0_uk_K_r13_12 ) , .QN( u0_uk_n36 ) );
  DFF_X1 u0_uk_K_r13_reg_13 (.CK( clk ) , .D( u0_uk_K_r12_13 ) , .Q( u0_uk_K_r13_13 ) , .QN( u0_uk_n35 ) );
  DFF_X1 u0_uk_K_r13_reg_14 (.CK( clk ) , .D( u0_uk_K_r12_14 ) , .Q( u0_uk_K_r13_14 ) , .QN( u0_uk_n34 ) );
  DFF_X1 u0_uk_K_r13_reg_15 (.CK( clk ) , .D( u0_uk_K_r12_15 ) , .Q( u0_uk_K_r13_15 ) , .QN( u0_uk_n33 ) );
  DFF_X1 u0_uk_K_r13_reg_16 (.CK( clk ) , .D( u0_uk_K_r12_16 ) , .Q( u0_uk_K_r13_16 ) , .QN( u0_uk_n32 ) );
  DFF_X1 u0_uk_K_r13_reg_17 (.CK( clk ) , .D( u0_uk_K_r12_17 ) , .Q( u0_uk_K_r13_17 ) );
  DFF_X1 u0_uk_K_r13_reg_18 (.CK( clk ) , .D( u0_uk_K_r12_18 ) , .Q( u0_uk_K_r13_18 ) , .QN( u0_uk_n30 ) );
  DFF_X1 u0_uk_K_r13_reg_19 (.CK( clk ) , .D( u0_uk_K_r12_19 ) , .Q( u0_uk_K_r13_19 ) );
  DFF_X1 u0_uk_K_r13_reg_2 (.CK( clk ) , .D( u0_uk_K_r12_2 ) , .Q( u0_uk_K_r13_2 ) );
  DFF_X1 u0_uk_K_r13_reg_20 (.CK( clk ) , .D( u0_uk_K_r12_20 ) , .Q( u0_uk_K_r13_20 ) , .QN( u0_uk_n29 ) );
  DFF_X1 u0_uk_K_r13_reg_21 (.CK( clk ) , .D( u0_uk_K_r12_21 ) , .Q( u0_uk_K_r13_21 ) , .QN( u0_uk_n28 ) );
  DFF_X1 u0_uk_K_r13_reg_22 (.CK( clk ) , .D( u0_uk_K_r12_22 ) , .Q( u0_uk_K_r13_22 ) );
  DFF_X1 u0_uk_K_r13_reg_23 (.CK( clk ) , .D( u0_uk_K_r12_23 ) , .Q( u0_uk_K_r13_23 ) );
  DFF_X1 u0_uk_K_r13_reg_24 (.CK( clk ) , .D( u0_uk_K_r12_24 ) , .Q( u0_uk_K_r13_24 ) , .QN( u0_uk_n26 ) );
  DFF_X1 u0_uk_K_r13_reg_25 (.CK( clk ) , .D( u0_uk_K_r12_25 ) , .Q( u0_uk_K_r13_25 ) );
  DFF_X1 u0_uk_K_r13_reg_26 (.CK( clk ) , .D( u0_uk_K_r12_26 ) , .Q( u0_uk_K_r13_26 ) , .QN( u0_uk_n25 ) );
  DFF_X1 u0_uk_K_r13_reg_27 (.CK( clk ) , .D( u0_uk_K_r12_27 ) , .Q( u0_uk_K_r13_27 ) , .QN( u0_uk_n24 ) );
  DFF_X1 u0_uk_K_r13_reg_28 (.CK( clk ) , .D( u0_uk_K_r12_28 ) , .Q( u0_uk_K_r13_28 ) , .QN( u0_uk_n23 ) );
  DFF_X1 u0_uk_K_r13_reg_29 (.CK( clk ) , .D( u0_uk_K_r12_29 ) , .Q( u0_uk_K_r13_29 ) , .QN( u0_uk_n22 ) );
  DFF_X1 u0_uk_K_r13_reg_3 (.CK( clk ) , .D( u0_uk_K_r12_3 ) , .Q( u0_uk_K_r13_3 ) , .QN( u0_uk_n44 ) );
  DFF_X1 u0_uk_K_r13_reg_30 (.CK( clk ) , .D( u0_uk_K_r12_30 ) , .Q( u0_uk_K_r13_30 ) , .QN( u0_uk_n21 ) );
  DFF_X1 u0_uk_K_r13_reg_31 (.CK( clk ) , .D( u0_uk_K_r12_31 ) , .Q( u0_uk_K_r13_31 ) );
  DFF_X1 u0_uk_K_r13_reg_32 (.CK( clk ) , .D( u0_uk_K_r12_32 ) , .Q( u0_uk_K_r13_32 ) );
  DFF_X1 u0_uk_K_r13_reg_33 (.CK( clk ) , .D( u0_uk_K_r12_33 ) , .Q( u0_uk_K_r13_33 ) , .QN( u0_uk_n20 ) );
  DFF_X1 u0_uk_K_r13_reg_34 (.CK( clk ) , .D( u0_uk_K_r12_34 ) , .Q( u0_uk_K_r13_34 ) , .QN( u0_uk_n19 ) );
  DFF_X1 u0_uk_K_r13_reg_35 (.CK( clk ) , .D( u0_uk_K_r12_35 ) , .Q( u0_uk_K_r13_35 ) );
  DFF_X1 u0_uk_K_r13_reg_36 (.CK( clk ) , .D( u0_uk_K_r12_36 ) , .Q( u0_uk_K_r13_36 ) );
  DFF_X1 u0_uk_K_r13_reg_37 (.CK( clk ) , .D( u0_uk_K_r12_37 ) , .Q( u0_uk_K_r13_37 ) , .QN( u0_uk_n18 ) );
  DFF_X1 u0_uk_K_r13_reg_38 (.CK( clk ) , .D( u0_uk_K_r12_38 ) , .Q( u0_uk_K_r13_38 ) );
  DFF_X1 u0_uk_K_r13_reg_39 (.CK( clk ) , .D( u0_uk_K_r12_39 ) , .Q( u0_uk_K_r13_39 ) , .QN( u0_uk_n16 ) );
  DFF_X1 u0_uk_K_r13_reg_4 (.CK( clk ) , .D( u0_uk_K_r12_4 ) , .Q( u0_uk_K_r13_4 ) );
  DFF_X1 u0_uk_K_r13_reg_40 (.CK( clk ) , .D( u0_uk_K_r12_40 ) , .Q( u0_uk_K_r13_40 ) , .QN( u0_uk_n15 ) );
  DFF_X1 u0_uk_K_r13_reg_41 (.CK( clk ) , .D( u0_uk_K_r12_41 ) , .Q( u0_uk_K_r13_41 ) , .QN( u0_uk_n14 ) );
  DFF_X1 u0_uk_K_r13_reg_42 (.CK( clk ) , .D( u0_uk_K_r12_42 ) , .Q( u0_uk_K_r13_42 ) , .QN( u0_uk_n13 ) );
  DFF_X1 u0_uk_K_r13_reg_43 (.CK( clk ) , .D( u0_uk_K_r12_43 ) , .Q( u0_uk_K_r13_43 ) , .QN( u0_uk_n12 ) );
  DFF_X1 u0_uk_K_r13_reg_44 (.CK( clk ) , .D( u0_uk_K_r12_44 ) , .Q( u0_uk_K_r13_44 ) );
  DFF_X1 u0_uk_K_r13_reg_45 (.CK( clk ) , .D( u0_uk_K_r12_45 ) , .Q( u0_uk_K_r13_45 ) , .QN( u0_uk_n9 ) );
  DFF_X1 u0_uk_K_r13_reg_46 (.CK( clk ) , .D( u0_uk_K_r12_46 ) , .Q( u0_uk_K_r13_46 ) , .QN( u0_uk_n8 ) );
  DFF_X1 u0_uk_K_r13_reg_47 (.CK( clk ) , .D( u0_uk_K_r12_47 ) , .Q( u0_uk_K_r13_47 ) , .QN( u0_uk_n7 ) );
  DFF_X1 u0_uk_K_r13_reg_48 (.CK( clk ) , .D( u0_uk_K_r12_48 ) , .Q( u0_uk_K_r13_48 ) , .QN( u0_uk_n6 ) );
  DFF_X1 u0_uk_K_r13_reg_49 (.CK( clk ) , .D( u0_uk_K_r12_49 ) , .Q( u0_uk_K_r13_49 ) , .QN( u0_uk_n5 ) );
  DFF_X1 u0_uk_K_r13_reg_5 (.CK( clk ) , .D( u0_uk_K_r12_5 ) , .Q( u0_uk_K_r13_5 ) , .QN( u0_uk_n43 ) );
  DFF_X1 u0_uk_K_r13_reg_50 (.CK( clk ) , .D( u0_uk_K_r12_50 ) , .Q( u0_uk_K_r13_50 ) , .QN( u0_uk_n4 ) );
  DFF_X1 u0_uk_K_r13_reg_51 (.CK( clk ) , .D( u0_uk_K_r12_51 ) , .Q( u0_uk_K_r13_51 ) , .QN( u0_uk_n3 ) );
  DFF_X1 u0_uk_K_r13_reg_52 (.CK( clk ) , .D( u0_uk_K_r12_52 ) , .Q( u0_uk_K_r13_52 ) , .QN( u0_uk_n2 ) );
  DFF_X1 u0_uk_K_r13_reg_53 (.CK( clk ) , .D( u0_uk_K_r12_53 ) , .Q( u0_uk_K_r13_53 ) );
  DFF_X1 u0_uk_K_r13_reg_54 (.CK( clk ) , .D( u0_uk_K_r12_54 ) , .Q( u0_uk_K_r13_54 ) , .QN( u0_uk_n1 ) );
  DFF_X1 u0_uk_K_r13_reg_55 (.CK( clk ) , .D( u0_uk_K_r12_55 ) , .Q( u0_uk_K_r13_55 ) );
  DFF_X1 u0_uk_K_r13_reg_6 (.CK( clk ) , .D( u0_uk_K_r12_6 ) , .Q( u0_uk_K_r13_6 ) , .QN( u0_uk_n42 ) );
  DFF_X1 u0_uk_K_r13_reg_7 (.CK( clk ) , .D( u0_uk_K_r12_7 ) , .Q( u0_uk_K_r13_7 ) , .QN( u0_uk_n41 ) );
  DFF_X1 u0_uk_K_r13_reg_8 (.CK( clk ) , .D( u0_uk_K_r12_8 ) , .Q( u0_uk_K_r13_8 ) , .QN( u0_uk_n40 ) );
  DFF_X1 u0_uk_K_r13_reg_9 (.CK( clk ) , .D( u0_uk_K_r12_9 ) , .Q( u0_uk_K_r13_9 ) , .QN( u0_uk_n39 ) );
  DFF_X1 u0_uk_K_r14_reg_0 (.CK( clk ) , .D( u0_uk_K_r13_0 ) , .QN( u0_uk_n670 ) );
  DFF_X1 u0_uk_K_r14_reg_1 (.CK( clk ) , .D( u0_uk_K_r13_1 ) , .QN( u0_uk_n669 ) );
  DFF_X1 u0_uk_K_r14_reg_10 (.CK( clk ) , .D( u0_uk_K_r13_10 ) , .Q( u0_uk_K_r14_10 ) );
  DFF_X1 u0_uk_K_r14_reg_11 (.CK( clk ) , .D( u0_uk_K_r13_11 ) , .Q( u0_uk_K_r14_11 ) );
  DFF_X1 u0_uk_K_r14_reg_12 (.CK( clk ) , .D( u0_uk_K_r13_12 ) , .Q( u0_uk_K_r14_12 ) );
  DFF_X1 u0_uk_K_r14_reg_13 (.CK( clk ) , .D( u0_uk_K_r13_13 ) , .QN( u0_uk_n664 ) );
  DFF_X1 u0_uk_K_r14_reg_14 (.CK( clk ) , .D( u0_uk_K_r13_14 ) , .QN( u0_uk_n663 ) );
  DFF_X1 u0_uk_K_r14_reg_15 (.CK( clk ) , .D( u0_uk_K_r13_15 ) , .Q( u0_uk_K_r14_15 ) );
  DFF_X1 u0_uk_K_r14_reg_16 (.CK( clk ) , .D( u0_uk_K_r13_16 ) , .Q( u0_uk_K_r14_16 ) );
  DFF_X1 u0_uk_K_r14_reg_17 (.CK( clk ) , .D( u0_uk_K_r13_17 ) , .QN( u0_uk_n661 ) );
  DFF_X1 u0_uk_K_r14_reg_18 (.CK( clk ) , .D( u0_uk_K_r13_18 ) , .Q( u0_uk_K_r14_18 ) );
  DFF_X1 u0_uk_K_r14_reg_19 (.CK( clk ) , .D( u0_uk_K_r13_19 ) , .QN( u0_uk_n660 ) );
  DFF_X1 u0_uk_K_r14_reg_2 (.CK( clk ) , .D( u0_uk_K_r13_2 ) , .Q( u0_uk_K_r14_2 ) );
  DFF_X1 u0_uk_K_r14_reg_20 (.CK( clk ) , .D( u0_uk_K_r13_20 ) , .QN( u0_uk_n659 ) );
  DFF_X1 u0_uk_K_r14_reg_21 (.CK( clk ) , .D( u0_uk_K_r13_21 ) , .QN( u0_uk_n658 ) );
  DFF_X1 u0_uk_K_r14_reg_22 (.CK( clk ) , .D( u0_uk_K_r13_22 ) , .QN( u0_uk_n657 ) );
  DFF_X1 u0_uk_K_r14_reg_23 (.CK( clk ) , .D( u0_uk_K_r13_23 ) , .Q( u0_uk_K_r14_23 ) , .QN( u0_uk_n655 ) );
  DFF_X1 u0_uk_K_r14_reg_24 (.CK( clk ) , .D( u0_uk_K_r13_24 ) , .QN( u0_uk_n654 ) );
  DFF_X1 u0_uk_K_r14_reg_25 (.CK( clk ) , .D( u0_uk_K_r13_25 ) , .QN( u0_uk_n653 ) );
  DFF_X1 u0_uk_K_r14_reg_26 (.CK( clk ) , .D( u0_uk_K_r13_26 ) , .QN( u0_uk_n652 ) );
  DFF_X1 u0_uk_K_r14_reg_27 (.CK( clk ) , .D( u0_uk_K_r13_27 ) , .QN( u0_uk_n651 ) );
  DFF_X1 u0_uk_K_r14_reg_28 (.CK( clk ) , .D( u0_uk_K_r13_28 ) , .QN( u0_uk_n650 ) );
  DFF_X1 u0_uk_K_r14_reg_29 (.CK( clk ) , .D( u0_uk_K_r13_29 ) , .QN( u0_uk_n649 ) );
  DFF_X1 u0_uk_K_r14_reg_3 (.CK( clk ) , .D( u0_uk_K_r13_3 ) , .Q( u0_uk_K_r14_3 ) );
  DFF_X1 u0_uk_K_r14_reg_30 (.CK( clk ) , .D( u0_uk_K_r13_30 ) , .QN( u0_uk_n648 ) );
  DFF_X1 u0_uk_K_r14_reg_31 (.CK( clk ) , .D( u0_uk_K_r13_31 ) , .QN( u0_uk_n647 ) );
  DFF_X1 u0_uk_K_r14_reg_32 (.CK( clk ) , .D( u0_uk_K_r13_32 ) , .QN( u0_uk_n646 ) );
  DFF_X1 u0_uk_K_r14_reg_33 (.CK( clk ) , .D( u0_uk_K_r13_33 ) , .QN( u0_uk_n645 ) );
  DFF_X1 u0_uk_K_r14_reg_34 (.CK( clk ) , .D( u0_uk_K_r13_34 ) , .QN( u0_uk_n644 ) );
  DFF_X1 u0_uk_K_r14_reg_35 (.CK( clk ) , .D( u0_uk_K_r13_35 ) , .QN( u0_uk_n643 ) );
  DFF_X1 u0_uk_K_r14_reg_36 (.CK( clk ) , .D( u0_uk_K_r13_36 ) , .QN( u0_uk_n642 ) );
  DFF_X1 u0_uk_K_r14_reg_37 (.CK( clk ) , .D( u0_uk_K_r13_37 ) , .QN( u0_uk_n641 ) );
  DFF_X1 u0_uk_K_r14_reg_38 (.CK( clk ) , .D( u0_uk_K_r13_38 ) , .Q( u0_uk_K_r14_38 ) );
  DFF_X1 u0_uk_K_r14_reg_39 (.CK( clk ) , .D( u0_uk_K_r13_39 ) , .Q( u0_uk_K_r14_39 ) );
  DFF_X1 u0_uk_K_r14_reg_4 (.CK( clk ) , .D( u0_uk_K_r13_4 ) , .QN( u0_uk_n668 ) );
  DFF_X1 u0_uk_K_r14_reg_40 (.CK( clk ) , .D( u0_uk_K_r13_40 ) , .QN( u0_uk_n640 ) );
  DFF_X1 u0_uk_K_r14_reg_41 (.CK( clk ) , .D( u0_uk_K_r13_41 ) , .QN( u0_uk_n639 ) );
  DFF_X1 u0_uk_K_r14_reg_42 (.CK( clk ) , .D( u0_uk_K_r13_42 ) , .Q( u0_uk_K_r14_42 ) );
  DFF_X1 u0_uk_K_r14_reg_43 (.CK( clk ) , .D( u0_uk_K_r13_43 ) , .Q( u0_uk_K_r14_43 ) );
  DFF_X1 u0_uk_K_r14_reg_44 (.CK( clk ) , .D( u0_uk_K_r13_44 ) , .QN( u0_uk_n638 ) );
  DFF_X1 u0_uk_K_r14_reg_45 (.CK( clk ) , .D( u0_uk_K_r13_45 ) , .Q( u0_uk_K_r14_45 ) );
  DFF_X1 u0_uk_K_r14_reg_46 (.CK( clk ) , .D( u0_uk_K_r13_46 ) , .Q( u0_uk_K_r14_46 ) );
  DFF_X1 u0_uk_K_r14_reg_47 (.CK( clk ) , .D( u0_uk_K_r13_47 ) , .QN( u0_uk_n637 ) );
  DFF_X1 u0_uk_K_r14_reg_48 (.CK( clk ) , .D( u0_uk_K_r13_48 ) , .QN( u0_uk_n636 ) );
  DFF_X1 u0_uk_K_r14_reg_49 (.CK( clk ) , .D( u0_uk_K_r13_49 ) , .QN( u0_uk_n635 ) );
  DFF_X1 u0_uk_K_r14_reg_5 (.CK( clk ) , .D( u0_uk_K_r13_5 ) , .Q( u0_uk_K_r14_5 ) );
  DFF_X1 u0_uk_K_r14_reg_50 (.CK( clk ) , .D( u0_uk_K_r13_50 ) , .Q( u0_uk_K_r14_50 ) );
  DFF_X1 u0_uk_K_r14_reg_51 (.CK( clk ) , .D( u0_uk_K_r13_51 ) , .QN( u0_uk_n633 ) );
  DFF_X1 u0_uk_K_r14_reg_52 (.CK( clk ) , .D( u0_uk_K_r13_52 ) , .QN( u0_uk_n632 ) );
  DFF_X1 u0_uk_K_r14_reg_53 (.CK( clk ) , .D( u0_uk_K_r13_53 ) , .QN( u0_uk_n631 ) );
  DFF_X1 u0_uk_K_r14_reg_54 (.CK( clk ) , .D( u0_uk_K_r13_54 ) , .QN( u0_uk_n630 ) );
  DFF_X1 u0_uk_K_r14_reg_55 (.CK( clk ) , .D( u0_uk_K_r13_55 ) , .QN( u0_uk_n629 ) );
  DFF_X1 u0_uk_K_r14_reg_6 (.CK( clk ) , .D( u0_uk_K_r13_6 ) , .QN( u0_uk_n667 ) );
  DFF_X1 u0_uk_K_r14_reg_7 (.CK( clk ) , .D( u0_uk_K_r13_7 ) , .QN( u0_uk_n666 ) );
  DFF_X1 u0_uk_K_r14_reg_8 (.CK( clk ) , .D( u0_uk_K_r13_8 ) , .Q( u0_uk_K_r14_8 ) );
  DFF_X1 u0_uk_K_r14_reg_9 (.CK( clk ) , .D( u0_uk_K_r13_9 ) , .Q( u0_uk_K_r14_9 ) );
  DFF_X1 u0_uk_K_r1_reg_0 (.CK( clk ) , .D( u0_uk_K_r0_0 ) , .Q( u0_uk_K_r1_0 ) , .QN( u0_uk_n581 ) );
  DFF_X1 u0_uk_K_r1_reg_1 (.CK( clk ) , .D( u0_uk_K_r0_1 ) , .Q( u0_uk_K_r1_1 ) , .QN( u0_uk_n580 ) );
  DFF_X1 u0_uk_K_r1_reg_10 (.CK( clk ) , .D( u0_uk_K_r0_10 ) , .Q( u0_uk_K_r1_10 ) );
  DFF_X1 u0_uk_K_r1_reg_11 (.CK( clk ) , .D( u0_uk_K_r0_11 ) , .Q( u0_uk_K_r1_11 ) , .QN( u0_uk_n573 ) );
  DFF_X1 u0_uk_K_r1_reg_12 (.CK( clk ) , .D( u0_uk_K_r0_12 ) , .Q( u0_uk_K_r1_12 ) , .QN( u0_uk_n572 ) );
  DFF_X1 u0_uk_K_r1_reg_13 (.CK( clk ) , .D( u0_uk_K_r0_13 ) , .Q( u0_uk_K_r1_13 ) , .QN( u0_uk_n571 ) );
  DFF_X1 u0_uk_K_r1_reg_14 (.CK( clk ) , .D( u0_uk_K_r0_14 ) , .Q( u0_uk_K_r1_14 ) , .QN( u0_uk_n570 ) );
  DFF_X1 u0_uk_K_r1_reg_15 (.CK( clk ) , .D( u0_uk_K_r0_15 ) , .Q( u0_uk_K_r1_15 ) );
  DFF_X1 u0_uk_K_r1_reg_16 (.CK( clk ) , .D( u0_uk_K_r0_16 ) , .Q( u0_uk_K_r1_16 ) );
  DFF_X1 u0_uk_K_r1_reg_17 (.CK( clk ) , .D( u0_uk_K_r0_17 ) , .Q( u0_uk_K_r1_17 ) , .QN( u0_uk_n569 ) );
  DFF_X1 u0_uk_K_r1_reg_18 (.CK( clk ) , .D( u0_uk_K_r0_18 ) , .Q( u0_uk_K_r1_18 ) );
  DFF_X1 u0_uk_K_r1_reg_19 (.CK( clk ) , .D( u0_uk_K_r0_19 ) , .Q( u0_uk_K_r1_19 ) , .QN( u0_uk_n568 ) );
  DFF_X1 u0_uk_K_r1_reg_2 (.CK( clk ) , .D( u0_uk_K_r0_2 ) , .Q( u0_uk_K_r1_2 ) , .QN( u0_uk_n579 ) );
  DFF_X1 u0_uk_K_r1_reg_20 (.CK( clk ) , .D( u0_uk_K_r0_20 ) , .Q( u0_uk_K_r1_20 ) , .QN( u0_uk_n567 ) );
  DFF_X1 u0_uk_K_r1_reg_21 (.CK( clk ) , .D( u0_uk_K_r0_21 ) , .Q( u0_uk_K_r1_21 ) );
  DFF_X1 u0_uk_K_r1_reg_22 (.CK( clk ) , .D( u0_uk_K_r0_22 ) , .Q( u0_uk_K_r1_22 ) );
  DFF_X1 u0_uk_K_r1_reg_23 (.CK( clk ) , .D( u0_uk_K_r0_23 ) , .Q( u0_uk_K_r1_23 ) , .QN( u0_uk_n566 ) );
  DFF_X1 u0_uk_K_r1_reg_24 (.CK( clk ) , .D( u0_uk_K_r0_24 ) , .Q( u0_uk_K_r1_24 ) , .QN( u0_uk_n565 ) );
  DFF_X1 u0_uk_K_r1_reg_25 (.CK( clk ) , .D( u0_uk_K_r0_25 ) , .Q( u0_uk_K_r1_25 ) , .QN( u0_uk_n564 ) );
  DFF_X1 u0_uk_K_r1_reg_26 (.CK( clk ) , .D( u0_uk_K_r0_26 ) , .Q( u0_uk_K_r1_26 ) , .QN( u0_uk_n563 ) );
  DFF_X1 u0_uk_K_r1_reg_27 (.CK( clk ) , .D( u0_uk_K_r0_27 ) , .Q( u0_uk_K_r1_27 ) , .QN( u0_uk_n562 ) );
  DFF_X1 u0_uk_K_r1_reg_28 (.CK( clk ) , .D( u0_uk_K_r0_28 ) , .Q( u0_uk_K_r1_28 ) , .QN( u0_uk_n561 ) );
  DFF_X1 u0_uk_K_r1_reg_29 (.CK( clk ) , .D( u0_uk_K_r0_29 ) , .Q( u0_uk_K_r1_29 ) , .QN( u0_uk_n560 ) );
  DFF_X1 u0_uk_K_r1_reg_3 (.CK( clk ) , .D( u0_uk_K_r0_3 ) , .Q( u0_uk_K_r1_3 ) , .QN( u0_uk_n578 ) );
  DFF_X1 u0_uk_K_r1_reg_30 (.CK( clk ) , .D( u0_uk_K_r0_30 ) , .Q( u0_uk_K_r1_30 ) , .QN( u0_uk_n559 ) );
  DFF_X1 u0_uk_K_r1_reg_31 (.CK( clk ) , .D( u0_uk_K_r0_31 ) , .Q( u0_uk_K_r1_31 ) , .QN( u0_uk_n558 ) );
  DFF_X1 u0_uk_K_r1_reg_32 (.CK( clk ) , .D( u0_uk_K_r0_32 ) , .Q( u0_uk_K_r1_32 ) , .QN( u0_uk_n557 ) );
  DFF_X1 u0_uk_K_r1_reg_33 (.CK( clk ) , .D( u0_uk_K_r0_33 ) , .Q( u0_uk_K_r1_33 ) );
  DFF_X1 u0_uk_K_r1_reg_34 (.CK( clk ) , .D( u0_uk_K_r0_34 ) , .Q( u0_uk_K_r1_34 ) , .QN( u0_uk_n556 ) );
  DFF_X1 u0_uk_K_r1_reg_35 (.CK( clk ) , .D( u0_uk_K_r0_35 ) , .Q( u0_uk_K_r1_35 ) , .QN( u0_uk_n555 ) );
  DFF_X1 u0_uk_K_r1_reg_36 (.CK( clk ) , .D( u0_uk_K_r0_36 ) , .Q( u0_uk_K_r1_36 ) );
  DFF_X1 u0_uk_K_r1_reg_37 (.CK( clk ) , .D( u0_uk_K_r0_37 ) , .Q( u0_uk_K_r1_37 ) , .QN( u0_uk_n554 ) );
  DFF_X1 u0_uk_K_r1_reg_38 (.CK( clk ) , .D( u0_uk_K_r0_38 ) , .Q( u0_uk_K_r1_38 ) , .QN( u0_uk_n553 ) );
  DFF_X1 u0_uk_K_r1_reg_39 (.CK( clk ) , .D( u0_uk_K_r0_39 ) , .Q( u0_uk_K_r1_39 ) );
  DFF_X1 u0_uk_K_r1_reg_4 (.CK( clk ) , .D( u0_uk_K_r0_4 ) , .Q( u0_uk_K_r1_4 ) , .QN( u0_uk_n577 ) );
  DFF_X1 u0_uk_K_r1_reg_40 (.CK( clk ) , .D( u0_uk_K_r0_40 ) , .Q( u0_uk_K_r1_40 ) , .QN( u0_uk_n552 ) );
  DFF_X1 u0_uk_K_r1_reg_41 (.CK( clk ) , .D( u0_uk_K_r0_41 ) , .Q( u0_uk_K_r1_41 ) );
  DFF_X1 u0_uk_K_r1_reg_42 (.CK( clk ) , .D( u0_uk_K_r0_42 ) , .Q( u0_uk_K_r1_42 ) );
  DFF_X1 u0_uk_K_r1_reg_43 (.CK( clk ) , .D( u0_uk_K_r0_43 ) , .Q( u0_uk_K_r1_43 ) , .QN( u0_uk_n550 ) );
  DFF_X1 u0_uk_K_r1_reg_44 (.CK( clk ) , .D( u0_uk_K_r0_44 ) , .Q( u0_uk_K_r1_44 ) );
  DFF_X1 u0_uk_K_r1_reg_45 (.CK( clk ) , .D( u0_uk_K_r0_45 ) , .Q( u0_uk_K_r1_45 ) , .QN( u0_uk_n549 ) );
  DFF_X1 u0_uk_K_r1_reg_46 (.CK( clk ) , .D( u0_uk_K_r0_46 ) , .Q( u0_uk_K_r1_46 ) , .QN( u0_uk_n548 ) );
  DFF_X1 u0_uk_K_r1_reg_47 (.CK( clk ) , .D( u0_uk_K_r0_47 ) , .Q( u0_uk_K_r1_47 ) );
  DFF_X1 u0_uk_K_r1_reg_48 (.CK( clk ) , .D( u0_uk_K_r0_48 ) , .Q( u0_uk_K_r1_48 ) , .QN( u0_uk_n547 ) );
  DFF_X1 u0_uk_K_r1_reg_49 (.CK( clk ) , .D( u0_uk_K_r0_49 ) , .Q( u0_uk_K_r1_49 ) , .QN( u0_uk_n546 ) );
  DFF_X1 u0_uk_K_r1_reg_5 (.CK( clk ) , .D( u0_uk_K_r0_5 ) , .Q( u0_uk_K_r1_5 ) , .QN( u0_uk_n576 ) );
  DFF_X1 u0_uk_K_r1_reg_50 (.CK( clk ) , .D( u0_uk_K_r0_50 ) , .Q( u0_uk_K_r1_50 ) , .QN( u0_uk_n545 ) );
  DFF_X1 u0_uk_K_r1_reg_51 (.CK( clk ) , .D( u0_uk_K_r0_51 ) , .Q( u0_uk_K_r1_51 ) , .QN( u0_uk_n544 ) );
  DFF_X1 u0_uk_K_r1_reg_52 (.CK( clk ) , .D( u0_uk_K_r0_52 ) , .Q( u0_uk_K_r1_52 ) , .QN( u0_uk_n543 ) );
  DFF_X1 u0_uk_K_r1_reg_53 (.CK( clk ) , .D( u0_uk_K_r0_53 ) , .Q( u0_uk_K_r1_53 ) , .QN( u0_uk_n542 ) );
  DFF_X1 u0_uk_K_r1_reg_54 (.CK( clk ) , .D( u0_uk_K_r0_54 ) , .Q( u0_uk_K_r1_54 ) , .QN( u0_uk_n541 ) );
  DFF_X1 u0_uk_K_r1_reg_55 (.CK( clk ) , .D( u0_uk_K_r0_55 ) , .Q( u0_uk_K_r1_55 ) , .QN( u0_uk_n540 ) );
  DFF_X1 u0_uk_K_r1_reg_6 (.CK( clk ) , .D( u0_uk_K_r0_6 ) , .Q( u0_uk_K_r1_6 ) );
  DFF_X1 u0_uk_K_r1_reg_7 (.CK( clk ) , .D( u0_uk_K_r0_7 ) , .Q( u0_uk_K_r1_7 ) );
  DFF_X1 u0_uk_K_r1_reg_8 (.CK( clk ) , .D( u0_uk_K_r0_8 ) , .Q( u0_uk_K_r1_8 ) , .QN( u0_uk_n575 ) );
  DFF_X1 u0_uk_K_r1_reg_9 (.CK( clk ) , .D( u0_uk_K_r0_9 ) , .Q( u0_uk_K_r1_9 ) , .QN( u0_uk_n574 ) );
  DFF_X1 u0_uk_K_r2_reg_0 (.CK( clk ) , .D( u0_uk_K_r1_0 ) , .Q( u0_uk_K_r2_0 ) , .QN( u0_uk_n539 ) );
  DFF_X1 u0_uk_K_r2_reg_1 (.CK( clk ) , .D( u0_uk_K_r1_1 ) , .Q( u0_uk_K_r2_1 ) , .QN( u0_uk_n538 ) );
  DFF_X1 u0_uk_K_r2_reg_10 (.CK( clk ) , .D( u0_uk_K_r1_10 ) , .Q( u0_uk_K_r2_10 ) , .QN( u0_uk_n531 ) );
  DFF_X1 u0_uk_K_r2_reg_11 (.CK( clk ) , .D( u0_uk_K_r1_11 ) , .Q( u0_uk_K_r2_11 ) , .QN( u0_uk_n530 ) );
  DFF_X1 u0_uk_K_r2_reg_12 (.CK( clk ) , .D( u0_uk_K_r1_12 ) , .Q( u0_uk_K_r2_12 ) , .QN( u0_uk_n529 ) );
  DFF_X1 u0_uk_K_r2_reg_13 (.CK( clk ) , .D( u0_uk_K_r1_13 ) , .Q( u0_uk_K_r2_13 ) );
  DFF_X1 u0_uk_K_r2_reg_14 (.CK( clk ) , .D( u0_uk_K_r1_14 ) , .Q( u0_uk_K_r2_14 ) , .QN( u0_uk_n528 ) );
  DFF_X1 u0_uk_K_r2_reg_15 (.CK( clk ) , .D( u0_uk_K_r1_15 ) , .Q( u0_uk_K_r2_15 ) , .QN( u0_uk_n527 ) );
  DFF_X1 u0_uk_K_r2_reg_16 (.CK( clk ) , .D( u0_uk_K_r1_16 ) , .Q( u0_uk_K_r2_16 ) );
  DFF_X1 u0_uk_K_r2_reg_17 (.CK( clk ) , .D( u0_uk_K_r1_17 ) , .Q( u0_uk_K_r2_17 ) , .QN( u0_uk_n525 ) );
  DFF_X1 u0_uk_K_r2_reg_18 (.CK( clk ) , .D( u0_uk_K_r1_18 ) , .Q( u0_uk_K_r2_18 ) );
  DFF_X1 u0_uk_K_r2_reg_19 (.CK( clk ) , .D( u0_uk_K_r1_19 ) , .Q( u0_uk_K_r2_19 ) , .QN( u0_uk_n523 ) );
  DFF_X1 u0_uk_K_r2_reg_2 (.CK( clk ) , .D( u0_uk_K_r1_2 ) , .Q( u0_uk_K_r2_2 ) , .QN( u0_uk_n537 ) );
  DFF_X1 u0_uk_K_r2_reg_20 (.CK( clk ) , .D( u0_uk_K_r1_20 ) , .Q( u0_uk_K_r2_20 ) );
  DFF_X1 u0_uk_K_r2_reg_21 (.CK( clk ) , .D( u0_uk_K_r1_21 ) , .Q( u0_uk_K_r2_21 ) );
  DFF_X1 u0_uk_K_r2_reg_22 (.CK( clk ) , .D( u0_uk_K_r1_22 ) , .Q( u0_uk_K_r2_22 ) , .QN( u0_uk_n522 ) );
  DFF_X1 u0_uk_K_r2_reg_23 (.CK( clk ) , .D( u0_uk_K_r1_23 ) , .Q( u0_uk_K_r2_23 ) , .QN( u0_uk_n521 ) );
  DFF_X1 u0_uk_K_r2_reg_24 (.CK( clk ) , .D( u0_uk_K_r1_24 ) , .Q( u0_uk_K_r2_24 ) );
  DFF_X1 u0_uk_K_r2_reg_25 (.CK( clk ) , .D( u0_uk_K_r1_25 ) , .Q( u0_uk_K_r2_25 ) );
  DFF_X1 u0_uk_K_r2_reg_26 (.CK( clk ) , .D( u0_uk_K_r1_26 ) , .Q( u0_uk_K_r2_26 ) );
  DFF_X1 u0_uk_K_r2_reg_27 (.CK( clk ) , .D( u0_uk_K_r1_27 ) , .Q( u0_uk_K_r2_27 ) );
  DFF_X1 u0_uk_K_r2_reg_28 (.CK( clk ) , .D( u0_uk_K_r1_28 ) , .Q( u0_uk_K_r2_28 ) );
  DFF_X1 u0_uk_K_r2_reg_29 (.CK( clk ) , .D( u0_uk_K_r1_29 ) , .Q( u0_uk_K_r2_29 ) );
  DFF_X1 u0_uk_K_r2_reg_3 (.CK( clk ) , .D( u0_uk_K_r1_3 ) , .Q( u0_uk_K_r2_3 ) , .QN( u0_uk_n536 ) );
  DFF_X1 u0_uk_K_r2_reg_30 (.CK( clk ) , .D( u0_uk_K_r1_30 ) , .Q( u0_uk_K_r2_30 ) );
  DFF_X1 u0_uk_K_r2_reg_31 (.CK( clk ) , .D( u0_uk_K_r1_31 ) , .Q( u0_uk_K_r2_31 ) );
  DFF_X1 u0_uk_K_r2_reg_32 (.CK( clk ) , .D( u0_uk_K_r1_32 ) , .Q( u0_uk_K_r2_32 ) , .QN( u0_uk_n519 ) );
  DFF_X1 u0_uk_K_r2_reg_33 (.CK( clk ) , .D( u0_uk_K_r1_33 ) , .Q( u0_uk_K_r2_33 ) );
  DFF_X1 u0_uk_K_r2_reg_34 (.CK( clk ) , .D( u0_uk_K_r1_34 ) , .Q( u0_uk_K_r2_34 ) , .QN( u0_uk_n517 ) );
  DFF_X1 u0_uk_K_r2_reg_35 (.CK( clk ) , .D( u0_uk_K_r1_35 ) , .Q( u0_uk_K_r2_35 ) , .QN( u0_uk_n516 ) );
  DFF_X1 u0_uk_K_r2_reg_36 (.CK( clk ) , .D( u0_uk_K_r1_36 ) , .Q( u0_uk_K_r2_36 ) , .QN( u0_uk_n514 ) );
  DFF_X1 u0_uk_K_r2_reg_37 (.CK( clk ) , .D( u0_uk_K_r1_37 ) , .Q( u0_uk_K_r2_37 ) , .QN( u0_uk_n513 ) );
  DFF_X1 u0_uk_K_r2_reg_38 (.CK( clk ) , .D( u0_uk_K_r1_38 ) , .Q( u0_uk_K_r2_38 ) , .QN( u0_uk_n512 ) );
  DFF_X1 u0_uk_K_r2_reg_39 (.CK( clk ) , .D( u0_uk_K_r1_39 ) , .Q( u0_uk_K_r2_39 ) , .QN( u0_uk_n511 ) );
  DFF_X1 u0_uk_K_r2_reg_4 (.CK( clk ) , .D( u0_uk_K_r1_4 ) , .Q( u0_uk_K_r2_4 ) );
  DFF_X1 u0_uk_K_r2_reg_40 (.CK( clk ) , .D( u0_uk_K_r1_40 ) , .Q( u0_uk_K_r2_40 ) , .QN( u0_uk_n510 ) );
  DFF_X1 u0_uk_K_r2_reg_41 (.CK( clk ) , .D( u0_uk_K_r1_41 ) , .Q( u0_uk_K_r2_41 ) );
  DFF_X1 u0_uk_K_r2_reg_42 (.CK( clk ) , .D( u0_uk_K_r1_42 ) , .Q( u0_uk_K_r2_42 ) , .QN( u0_uk_n508 ) );
  DFF_X1 u0_uk_K_r2_reg_43 (.CK( clk ) , .D( u0_uk_K_r1_43 ) , .Q( u0_uk_K_r2_43 ) , .QN( u0_uk_n507 ) );
  DFF_X1 u0_uk_K_r2_reg_44 (.CK( clk ) , .D( u0_uk_K_r1_44 ) , .Q( u0_uk_K_r2_44 ) , .QN( u0_uk_n506 ) );
  DFF_X1 u0_uk_K_r2_reg_45 (.CK( clk ) , .D( u0_uk_K_r1_45 ) , .Q( u0_uk_K_r2_45 ) , .QN( u0_uk_n505 ) );
  DFF_X1 u0_uk_K_r2_reg_46 (.CK( clk ) , .D( u0_uk_K_r1_46 ) , .Q( u0_uk_K_r2_46 ) );
  DFF_X1 u0_uk_K_r2_reg_47 (.CK( clk ) , .D( u0_uk_K_r1_47 ) , .Q( u0_uk_K_r2_47 ) );
  DFF_X1 u0_uk_K_r2_reg_48 (.CK( clk ) , .D( u0_uk_K_r1_48 ) , .Q( u0_uk_K_r2_48 ) , .QN( u0_uk_n502 ) );
  DFF_X1 u0_uk_K_r2_reg_49 (.CK( clk ) , .D( u0_uk_K_r1_49 ) , .Q( u0_uk_K_r2_49 ) );
  DFF_X1 u0_uk_K_r2_reg_5 (.CK( clk ) , .D( u0_uk_K_r1_5 ) , .Q( u0_uk_K_r2_5 ) , .QN( u0_uk_n535 ) );
  DFF_X1 u0_uk_K_r2_reg_50 (.CK( clk ) , .D( u0_uk_K_r1_50 ) , .Q( u0_uk_K_r2_50 ) );
  DFF_X1 u0_uk_K_r2_reg_51 (.CK( clk ) , .D( u0_uk_K_r1_51 ) , .Q( u0_uk_K_r2_51 ) , .QN( u0_uk_n499 ) );
  DFF_X1 u0_uk_K_r2_reg_52 (.CK( clk ) , .D( u0_uk_K_r1_52 ) , .Q( u0_uk_K_r2_52 ) , .QN( u0_uk_n498 ) );
  DFF_X1 u0_uk_K_r2_reg_53 (.CK( clk ) , .D( u0_uk_K_r1_53 ) , .Q( u0_uk_K_r2_53 ) );
  DFF_X1 u0_uk_K_r2_reg_54 (.CK( clk ) , .D( u0_uk_K_r1_54 ) , .Q( u0_uk_K_r2_54 ) , .QN( u0_uk_n497 ) );
  DFF_X1 u0_uk_K_r2_reg_55 (.CK( clk ) , .D( u0_uk_K_r1_55 ) , .Q( u0_uk_K_r2_55 ) , .QN( u0_uk_n495 ) );
  DFF_X1 u0_uk_K_r2_reg_6 (.CK( clk ) , .D( u0_uk_K_r1_6 ) , .Q( u0_uk_K_r2_6 ) , .QN( u0_uk_n534 ) );
  DFF_X1 u0_uk_K_r2_reg_7 (.CK( clk ) , .D( u0_uk_K_r1_7 ) , .Q( u0_uk_K_r2_7 ) );
  DFF_X1 u0_uk_K_r2_reg_8 (.CK( clk ) , .D( u0_uk_K_r1_8 ) , .Q( u0_uk_K_r2_8 ) , .QN( u0_uk_n533 ) );
  DFF_X1 u0_uk_K_r2_reg_9 (.CK( clk ) , .D( u0_uk_K_r1_9 ) , .Q( u0_uk_K_r2_9 ) , .QN( u0_uk_n532 ) );
  DFF_X1 u0_uk_K_r3_reg_0 (.CK( clk ) , .D( u0_uk_K_r2_0 ) , .Q( u0_uk_K_r3_0 ) , .QN( u0_uk_n494 ) );
  DFF_X1 u0_uk_K_r3_reg_1 (.CK( clk ) , .D( u0_uk_K_r2_1 ) , .Q( u0_uk_K_r3_1 ) , .QN( u0_uk_n493 ) );
  DFF_X1 u0_uk_K_r3_reg_10 (.CK( clk ) , .D( u0_uk_K_r2_10 ) , .Q( u0_uk_K_r3_10 ) );
  DFF_X1 u0_uk_K_r3_reg_11 (.CK( clk ) , .D( u0_uk_K_r2_11 ) , .Q( u0_uk_K_r3_11 ) );
  DFF_X1 u0_uk_K_r3_reg_12 (.CK( clk ) , .D( u0_uk_K_r2_12 ) , .Q( u0_uk_K_r3_12 ) , .QN( u0_uk_n486 ) );
  DFF_X1 u0_uk_K_r3_reg_13 (.CK( clk ) , .D( u0_uk_K_r2_13 ) , .Q( u0_uk_K_r3_13 ) );
  DFF_X1 u0_uk_K_r3_reg_14 (.CK( clk ) , .D( u0_uk_K_r2_14 ) , .Q( u0_uk_K_r3_14 ) );
  DFF_X1 u0_uk_K_r3_reg_15 (.CK( clk ) , .D( u0_uk_K_r2_15 ) , .Q( u0_uk_K_r3_15 ) );
  DFF_X1 u0_uk_K_r3_reg_16 (.CK( clk ) , .D( u0_uk_K_r2_16 ) , .Q( u0_uk_K_r3_16 ) );
  DFF_X1 u0_uk_K_r3_reg_17 (.CK( clk ) , .D( u0_uk_K_r2_17 ) , .Q( u0_uk_K_r3_17 ) , .QN( u0_uk_n485 ) );
  DFF_X1 u0_uk_K_r3_reg_18 (.CK( clk ) , .D( u0_uk_K_r2_18 ) , .Q( u0_uk_K_r3_18 ) , .QN( u0_uk_n484 ) );
  DFF_X1 u0_uk_K_r3_reg_19 (.CK( clk ) , .D( u0_uk_K_r2_19 ) , .Q( u0_uk_K_r3_19 ) );
  DFF_X1 u0_uk_K_r3_reg_2 (.CK( clk ) , .D( u0_uk_K_r2_2 ) , .Q( u0_uk_K_r3_2 ) , .QN( u0_uk_n492 ) );
  DFF_X1 u0_uk_K_r3_reg_20 (.CK( clk ) , .D( u0_uk_K_r2_20 ) , .Q( u0_uk_K_r3_20 ) , .QN( u0_uk_n483 ) );
  DFF_X1 u0_uk_K_r3_reg_21 (.CK( clk ) , .D( u0_uk_K_r2_21 ) , .Q( u0_uk_K_r3_21 ) , .QN( u0_uk_n482 ) );
  DFF_X1 u0_uk_K_r3_reg_22 (.CK( clk ) , .D( u0_uk_K_r2_22 ) , .Q( u0_uk_K_r3_22 ) , .QN( u0_uk_n481 ) );
  DFF_X1 u0_uk_K_r3_reg_23 (.CK( clk ) , .D( u0_uk_K_r2_23 ) , .Q( u0_uk_K_r3_23 ) , .QN( u0_uk_n480 ) );
  DFF_X1 u0_uk_K_r3_reg_24 (.CK( clk ) , .D( u0_uk_K_r2_24 ) , .Q( u0_uk_K_r3_24 ) );
  DFF_X1 u0_uk_K_r3_reg_25 (.CK( clk ) , .D( u0_uk_K_r2_25 ) , .Q( u0_uk_K_r3_25 ) , .QN( u0_uk_n479 ) );
  DFF_X1 u0_uk_K_r3_reg_26 (.CK( clk ) , .D( u0_uk_K_r2_26 ) , .Q( u0_uk_K_r3_26 ) , .QN( u0_uk_n478 ) );
  DFF_X1 u0_uk_K_r3_reg_27 (.CK( clk ) , .D( u0_uk_K_r2_27 ) , .Q( u0_uk_K_r3_27 ) , .QN( u0_uk_n477 ) );
  DFF_X1 u0_uk_K_r3_reg_28 (.CK( clk ) , .D( u0_uk_K_r2_28 ) , .Q( u0_uk_K_r3_28 ) , .QN( u0_uk_n476 ) );
  DFF_X1 u0_uk_K_r3_reg_29 (.CK( clk ) , .D( u0_uk_K_r2_29 ) , .Q( u0_uk_K_r3_29 ) );
  DFF_X1 u0_uk_K_r3_reg_3 (.CK( clk ) , .D( u0_uk_K_r2_3 ) , .Q( u0_uk_K_r3_3 ) , .QN( u0_uk_n491 ) );
  DFF_X1 u0_uk_K_r3_reg_30 (.CK( clk ) , .D( u0_uk_K_r2_30 ) , .Q( u0_uk_K_r3_30 ) , .QN( u0_uk_n475 ) );
  DFF_X1 u0_uk_K_r3_reg_31 (.CK( clk ) , .D( u0_uk_K_r2_31 ) , .Q( u0_uk_K_r3_31 ) , .QN( u0_uk_n474 ) );
  DFF_X1 u0_uk_K_r3_reg_32 (.CK( clk ) , .D( u0_uk_K_r2_32 ) , .Q( u0_uk_K_r3_32 ) , .QN( u0_uk_n473 ) );
  DFF_X1 u0_uk_K_r3_reg_33 (.CK( clk ) , .D( u0_uk_K_r2_33 ) , .Q( u0_uk_K_r3_33 ) , .QN( u0_uk_n471 ) );
  DFF_X1 u0_uk_K_r3_reg_34 (.CK( clk ) , .D( u0_uk_K_r2_34 ) , .Q( u0_uk_K_r3_34 ) );
  DFF_X1 u0_uk_K_r3_reg_35 (.CK( clk ) , .D( u0_uk_K_r2_35 ) , .Q( u0_uk_K_r3_35 ) );
  DFF_X1 u0_uk_K_r3_reg_36 (.CK( clk ) , .D( u0_uk_K_r2_36 ) , .Q( u0_uk_K_r3_36 ) , .QN( u0_uk_n470 ) );
  DFF_X1 u0_uk_K_r3_reg_37 (.CK( clk ) , .D( u0_uk_K_r2_37 ) , .Q( u0_uk_K_r3_37 ) , .QN( u0_uk_n469 ) );
  DFF_X1 u0_uk_K_r3_reg_38 (.CK( clk ) , .D( u0_uk_K_r2_38 ) , .Q( u0_uk_K_r3_38 ) );
  DFF_X1 u0_uk_K_r3_reg_39 (.CK( clk ) , .D( u0_uk_K_r2_39 ) , .Q( u0_uk_K_r3_39 ) , .QN( u0_uk_n466 ) );
  DFF_X1 u0_uk_K_r3_reg_4 (.CK( clk ) , .D( u0_uk_K_r2_4 ) , .Q( u0_uk_K_r3_4 ) );
  DFF_X1 u0_uk_K_r3_reg_40 (.CK( clk ) , .D( u0_uk_K_r2_40 ) , .Q( u0_uk_K_r3_40 ) , .QN( u0_uk_n465 ) );
  DFF_X1 u0_uk_K_r3_reg_41 (.CK( clk ) , .D( u0_uk_K_r2_41 ) , .Q( u0_uk_K_r3_41 ) , .QN( u0_uk_n464 ) );
  DFF_X1 u0_uk_K_r3_reg_42 (.CK( clk ) , .D( u0_uk_K_r2_42 ) , .Q( u0_uk_K_r3_42 ) , .QN( u0_uk_n463 ) );
  DFF_X1 u0_uk_K_r3_reg_43 (.CK( clk ) , .D( u0_uk_K_r2_43 ) , .Q( u0_uk_K_r3_43 ) );
  DFF_X1 u0_uk_K_r3_reg_44 (.CK( clk ) , .D( u0_uk_K_r2_44 ) , .Q( u0_uk_K_r3_44 ) );
  DFF_X1 u0_uk_K_r3_reg_45 (.CK( clk ) , .D( u0_uk_K_r2_45 ) , .Q( u0_uk_K_r3_45 ) , .QN( u0_uk_n462 ) );
  DFF_X1 u0_uk_K_r3_reg_46 (.CK( clk ) , .D( u0_uk_K_r2_46 ) , .Q( u0_uk_K_r3_46 ) , .QN( u0_uk_n461 ) );
  DFF_X1 u0_uk_K_r3_reg_47 (.CK( clk ) , .D( u0_uk_K_r2_47 ) , .Q( u0_uk_K_r3_47 ) );
  DFF_X1 u0_uk_K_r3_reg_48 (.CK( clk ) , .D( u0_uk_K_r2_48 ) , .Q( u0_uk_K_r3_48 ) , .QN( u0_uk_n459 ) );
  DFF_X1 u0_uk_K_r3_reg_49 (.CK( clk ) , .D( u0_uk_K_r2_49 ) , .Q( u0_uk_K_r3_49 ) , .QN( u0_uk_n458 ) );
  DFF_X1 u0_uk_K_r3_reg_5 (.CK( clk ) , .D( u0_uk_K_r2_5 ) , .Q( u0_uk_K_r3_5 ) , .QN( u0_uk_n490 ) );
  DFF_X1 u0_uk_K_r3_reg_50 (.CK( clk ) , .D( u0_uk_K_r2_50 ) , .Q( u0_uk_K_r3_50 ) , .QN( u0_uk_n457 ) );
  DFF_X1 u0_uk_K_r3_reg_51 (.CK( clk ) , .D( u0_uk_K_r2_51 ) , .Q( u0_uk_K_r3_51 ) , .QN( u0_uk_n455 ) );
  DFF_X1 u0_uk_K_r3_reg_52 (.CK( clk ) , .D( u0_uk_K_r2_52 ) , .Q( u0_uk_K_r3_52 ) );
  DFF_X1 u0_uk_K_r3_reg_53 (.CK( clk ) , .D( u0_uk_K_r2_53 ) , .Q( u0_uk_K_r3_53 ) , .QN( u0_uk_n453 ) );
  DFF_X1 u0_uk_K_r3_reg_54 (.CK( clk ) , .D( u0_uk_K_r2_54 ) , .Q( u0_uk_K_r3_54 ) , .QN( u0_uk_n452 ) );
  DFF_X1 u0_uk_K_r3_reg_55 (.CK( clk ) , .D( u0_uk_K_r2_55 ) , .Q( u0_uk_K_r3_55 ) , .QN( u0_uk_n451 ) );
  DFF_X1 u0_uk_K_r3_reg_6 (.CK( clk ) , .D( u0_uk_K_r2_6 ) , .Q( u0_uk_K_r3_6 ) , .QN( u0_uk_n489 ) );
  DFF_X1 u0_uk_K_r3_reg_7 (.CK( clk ) , .D( u0_uk_K_r2_7 ) , .Q( u0_uk_K_r3_7 ) , .QN( u0_uk_n488 ) );
  DFF_X1 u0_uk_K_r3_reg_8 (.CK( clk ) , .D( u0_uk_K_r2_8 ) , .Q( u0_uk_K_r3_8 ) , .QN( u0_uk_n487 ) );
  DFF_X1 u0_uk_K_r3_reg_9 (.CK( clk ) , .D( u0_uk_K_r2_9 ) , .Q( u0_uk_K_r3_9 ) );
  DFF_X1 u0_uk_K_r4_reg_0 (.CK( clk ) , .D( u0_uk_K_r3_0 ) , .Q( u0_uk_K_r4_0 ) );
  DFF_X1 u0_uk_K_r4_reg_1 (.CK( clk ) , .D( u0_uk_K_r3_1 ) , .Q( u0_uk_K_r4_1 ) , .QN( u0_uk_n450 ) );
  DFF_X1 u0_uk_K_r4_reg_10 (.CK( clk ) , .D( u0_uk_K_r3_10 ) , .Q( u0_uk_K_r4_10 ) , .QN( u0_uk_n444 ) );
  DFF_X1 u0_uk_K_r4_reg_11 (.CK( clk ) , .D( u0_uk_K_r3_11 ) , .Q( u0_uk_K_r4_11 ) );
  DFF_X1 u0_uk_K_r4_reg_12 (.CK( clk ) , .D( u0_uk_K_r3_12 ) , .Q( u0_uk_K_r4_12 ) , .QN( u0_uk_n442 ) );
  DFF_X1 u0_uk_K_r4_reg_13 (.CK( clk ) , .D( u0_uk_K_r3_13 ) , .Q( u0_uk_K_r4_13 ) , .QN( u0_uk_n441 ) );
  DFF_X1 u0_uk_K_r4_reg_14 (.CK( clk ) , .D( u0_uk_K_r3_14 ) , .Q( u0_uk_K_r4_14 ) , .QN( u0_uk_n440 ) );
  DFF_X1 u0_uk_K_r4_reg_15 (.CK( clk ) , .D( u0_uk_K_r3_15 ) , .Q( u0_uk_K_r4_15 ) , .QN( u0_uk_n439 ) );
  DFF_X1 u0_uk_K_r4_reg_16 (.CK( clk ) , .D( u0_uk_K_r3_16 ) , .Q( u0_uk_K_r4_16 ) , .QN( u0_uk_n438 ) );
  DFF_X1 u0_uk_K_r4_reg_17 (.CK( clk ) , .D( u0_uk_K_r3_17 ) , .Q( u0_uk_K_r4_17 ) );
  DFF_X1 u0_uk_K_r4_reg_18 (.CK( clk ) , .D( u0_uk_K_r3_18 ) , .Q( u0_uk_K_r4_18 ) );
  DFF_X1 u0_uk_K_r4_reg_19 (.CK( clk ) , .D( u0_uk_K_r3_19 ) , .Q( u0_uk_K_r4_19 ) , .QN( u0_uk_n436 ) );
  DFF_X1 u0_uk_K_r4_reg_2 (.CK( clk ) , .D( u0_uk_K_r3_2 ) , .Q( u0_uk_K_r4_2 ) );
  DFF_X1 u0_uk_K_r4_reg_20 (.CK( clk ) , .D( u0_uk_K_r3_20 ) , .Q( u0_uk_K_r4_20 ) , .QN( u0_uk_n435 ) );
  DFF_X1 u0_uk_K_r4_reg_21 (.CK( clk ) , .D( u0_uk_K_r3_21 ) , .Q( u0_uk_K_r4_21 ) , .QN( u0_uk_n434 ) );
  DFF_X1 u0_uk_K_r4_reg_22 (.CK( clk ) , .D( u0_uk_K_r3_22 ) , .Q( u0_uk_K_r4_22 ) , .QN( u0_uk_n433 ) );
  DFF_X1 u0_uk_K_r4_reg_23 (.CK( clk ) , .D( u0_uk_K_r3_23 ) , .Q( u0_uk_K_r4_23 ) );
  DFF_X1 u0_uk_K_r4_reg_24 (.CK( clk ) , .D( u0_uk_K_r3_24 ) , .Q( u0_uk_K_r4_24 ) );
  DFF_X1 u0_uk_K_r4_reg_25 (.CK( clk ) , .D( u0_uk_K_r3_25 ) , .Q( u0_uk_K_r4_25 ) , .QN( u0_uk_n432 ) );
  DFF_X1 u0_uk_K_r4_reg_26 (.CK( clk ) , .D( u0_uk_K_r3_26 ) , .Q( u0_uk_K_r4_26 ) , .QN( u0_uk_n431 ) );
  DFF_X1 u0_uk_K_r4_reg_27 (.CK( clk ) , .D( u0_uk_K_r3_27 ) , .Q( u0_uk_K_r4_27 ) );
  DFF_X1 u0_uk_K_r4_reg_28 (.CK( clk ) , .D( u0_uk_K_r3_28 ) , .Q( u0_uk_K_r4_28 ) , .QN( u0_uk_n430 ) );
  DFF_X1 u0_uk_K_r4_reg_29 (.CK( clk ) , .D( u0_uk_K_r3_29 ) , .Q( u0_uk_K_r4_29 ) , .QN( u0_uk_n429 ) );
  DFF_X1 u0_uk_K_r4_reg_3 (.CK( clk ) , .D( u0_uk_K_r3_3 ) , .Q( u0_uk_K_r4_3 ) );
  DFF_X1 u0_uk_K_r4_reg_30 (.CK( clk ) , .D( u0_uk_K_r3_30 ) , .Q( u0_uk_K_r4_30 ) , .QN( u0_uk_n428 ) );
  DFF_X1 u0_uk_K_r4_reg_31 (.CK( clk ) , .D( u0_uk_K_r3_31 ) , .Q( u0_uk_K_r4_31 ) );
  DFF_X1 u0_uk_K_r4_reg_32 (.CK( clk ) , .D( u0_uk_K_r3_32 ) , .Q( u0_uk_K_r4_32 ) , .QN( u0_uk_n427 ) );
  DFF_X1 u0_uk_K_r4_reg_33 (.CK( clk ) , .D( u0_uk_K_r3_33 ) , .Q( u0_uk_K_r4_33 ) );
  DFF_X1 u0_uk_K_r4_reg_34 (.CK( clk ) , .D( u0_uk_K_r3_34 ) , .Q( u0_uk_K_r4_34 ) , .QN( u0_uk_n426 ) );
  DFF_X1 u0_uk_K_r4_reg_35 (.CK( clk ) , .D( u0_uk_K_r3_35 ) , .Q( u0_uk_K_r4_35 ) );
  DFF_X1 u0_uk_K_r4_reg_36 (.CK( clk ) , .D( u0_uk_K_r3_36 ) , .Q( u0_uk_K_r4_36 ) , .QN( u0_uk_n425 ) );
  DFF_X1 u0_uk_K_r4_reg_37 (.CK( clk ) , .D( u0_uk_K_r3_37 ) , .Q( u0_uk_K_r4_37 ) , .QN( u0_uk_n424 ) );
  DFF_X1 u0_uk_K_r4_reg_38 (.CK( clk ) , .D( u0_uk_K_r3_38 ) , .Q( u0_uk_K_r4_38 ) );
  DFF_X1 u0_uk_K_r4_reg_39 (.CK( clk ) , .D( u0_uk_K_r3_39 ) , .Q( u0_uk_K_r4_39 ) , .QN( u0_uk_n423 ) );
  DFF_X1 u0_uk_K_r4_reg_4 (.CK( clk ) , .D( u0_uk_K_r3_4 ) , .Q( u0_uk_K_r4_4 ) , .QN( u0_uk_n449 ) );
  DFF_X1 u0_uk_K_r4_reg_40 (.CK( clk ) , .D( u0_uk_K_r3_40 ) , .Q( u0_uk_K_r4_40 ) , .QN( u0_uk_n422 ) );
  DFF_X1 u0_uk_K_r4_reg_41 (.CK( clk ) , .D( u0_uk_K_r3_41 ) , .Q( u0_uk_K_r4_41 ) );
  DFF_X1 u0_uk_K_r4_reg_42 (.CK( clk ) , .D( u0_uk_K_r3_42 ) , .Q( u0_uk_K_r4_42 ) , .QN( u0_uk_n420 ) );
  DFF_X1 u0_uk_K_r4_reg_43 (.CK( clk ) , .D( u0_uk_K_r3_43 ) , .Q( u0_uk_K_r4_43 ) , .QN( u0_uk_n419 ) );
  DFF_X1 u0_uk_K_r4_reg_44 (.CK( clk ) , .D( u0_uk_K_r3_44 ) , .Q( u0_uk_K_r4_44 ) , .QN( u0_uk_n418 ) );
  DFF_X1 u0_uk_K_r4_reg_45 (.CK( clk ) , .D( u0_uk_K_r3_45 ) , .Q( u0_uk_K_r4_45 ) , .QN( u0_uk_n417 ) );
  DFF_X1 u0_uk_K_r4_reg_46 (.CK( clk ) , .D( u0_uk_K_r3_46 ) , .Q( u0_uk_K_r4_46 ) , .QN( u0_uk_n416 ) );
  DFF_X1 u0_uk_K_r4_reg_47 (.CK( clk ) , .D( u0_uk_K_r3_47 ) , .Q( u0_uk_K_r4_47 ) , .QN( u0_uk_n414 ) );
  DFF_X1 u0_uk_K_r4_reg_48 (.CK( clk ) , .D( u0_uk_K_r3_48 ) , .Q( u0_uk_K_r4_48 ) );
  DFF_X1 u0_uk_K_r4_reg_49 (.CK( clk ) , .D( u0_uk_K_r3_49 ) , .Q( u0_uk_K_r4_49 ) );
  DFF_X1 u0_uk_K_r4_reg_5 (.CK( clk ) , .D( u0_uk_K_r3_5 ) , .Q( u0_uk_K_r4_5 ) );
  DFF_X1 u0_uk_K_r4_reg_50 (.CK( clk ) , .D( u0_uk_K_r3_50 ) , .Q( u0_uk_K_r4_50 ) , .QN( u0_uk_n413 ) );
  DFF_X1 u0_uk_K_r4_reg_51 (.CK( clk ) , .D( u0_uk_K_r3_51 ) , .Q( u0_uk_K_r4_51 ) , .QN( u0_uk_n412 ) );
  DFF_X1 u0_uk_K_r4_reg_52 (.CK( clk ) , .D( u0_uk_K_r3_52 ) , .Q( u0_uk_K_r4_52 ) , .QN( u0_uk_n411 ) );
  DFF_X1 u0_uk_K_r4_reg_53 (.CK( clk ) , .D( u0_uk_K_r3_53 ) , .Q( u0_uk_K_r4_53 ) , .QN( u0_uk_n410 ) );
  DFF_X1 u0_uk_K_r4_reg_54 (.CK( clk ) , .D( u0_uk_K_r3_54 ) , .Q( u0_uk_K_r4_54 ) );
  DFF_X1 u0_uk_K_r4_reg_55 (.CK( clk ) , .D( u0_uk_K_r3_55 ) , .Q( u0_uk_K_r4_55 ) );
  DFF_X1 u0_uk_K_r4_reg_6 (.CK( clk ) , .D( u0_uk_K_r3_6 ) , .Q( u0_uk_K_r4_6 ) , .QN( u0_uk_n448 ) );
  DFF_X1 u0_uk_K_r4_reg_7 (.CK( clk ) , .D( u0_uk_K_r3_7 ) , .Q( u0_uk_K_r4_7 ) , .QN( u0_uk_n447 ) );
  DFF_X1 u0_uk_K_r4_reg_8 (.CK( clk ) , .D( u0_uk_K_r3_8 ) , .Q( u0_uk_K_r4_8 ) , .QN( u0_uk_n446 ) );
  DFF_X1 u0_uk_K_r4_reg_9 (.CK( clk ) , .D( u0_uk_K_r3_9 ) , .Q( u0_uk_K_r4_9 ) , .QN( u0_uk_n445 ) );
  DFF_X1 u0_uk_K_r5_reg_0 (.CK( clk ) , .D( u0_uk_K_r4_0 ) , .Q( u0_uk_K_r5_0 ) );
  DFF_X1 u0_uk_K_r5_reg_1 (.CK( clk ) , .D( u0_uk_K_r4_1 ) , .Q( u0_uk_K_r5_1 ) );
  DFF_X1 u0_uk_K_r5_reg_10 (.CK( clk ) , .D( u0_uk_K_r4_10 ) , .Q( u0_uk_K_r5_10 ) );
  DFF_X1 u0_uk_K_r5_reg_11 (.CK( clk ) , .D( u0_uk_K_r4_11 ) , .Q( u0_uk_K_r5_11 ) , .QN( u0_uk_n401 ) );
  DFF_X1 u0_uk_K_r5_reg_12 (.CK( clk ) , .D( u0_uk_K_r4_12 ) , .Q( u0_uk_K_r5_12 ) , .QN( u0_uk_n400 ) );
  DFF_X1 u0_uk_K_r5_reg_13 (.CK( clk ) , .D( u0_uk_K_r4_13 ) , .Q( u0_uk_K_r5_13 ) );
  DFF_X1 u0_uk_K_r5_reg_14 (.CK( clk ) , .D( u0_uk_K_r4_14 ) , .Q( u0_uk_K_r5_14 ) , .QN( u0_uk_n399 ) );
  DFF_X1 u0_uk_K_r5_reg_15 (.CK( clk ) , .D( u0_uk_K_r4_15 ) , .Q( u0_uk_K_r5_15 ) , .QN( u0_uk_n398 ) );
  DFF_X1 u0_uk_K_r5_reg_16 (.CK( clk ) , .D( u0_uk_K_r4_16 ) , .Q( u0_uk_K_r5_16 ) );
  DFF_X1 u0_uk_K_r5_reg_17 (.CK( clk ) , .D( u0_uk_K_r4_17 ) , .Q( u0_uk_K_r5_17 ) , .QN( u0_uk_n397 ) );
  DFF_X1 u0_uk_K_r5_reg_18 (.CK( clk ) , .D( u0_uk_K_r4_18 ) , .Q( u0_uk_K_r5_18 ) );
  DFF_X1 u0_uk_K_r5_reg_19 (.CK( clk ) , .D( u0_uk_K_r4_19 ) , .Q( u0_uk_K_r5_19 ) );
  DFF_X1 u0_uk_K_r5_reg_2 (.CK( clk ) , .D( u0_uk_K_r4_2 ) , .Q( u0_uk_K_r5_2 ) , .QN( u0_uk_n406 ) );
  DFF_X1 u0_uk_K_r5_reg_20 (.CK( clk ) , .D( u0_uk_K_r4_20 ) , .Q( u0_uk_K_r5_20 ) , .QN( u0_uk_n396 ) );
  DFF_X1 u0_uk_K_r5_reg_21 (.CK( clk ) , .D( u0_uk_K_r4_21 ) , .Q( u0_uk_K_r5_21 ) );
  DFF_X1 u0_uk_K_r5_reg_22 (.CK( clk ) , .D( u0_uk_K_r4_22 ) , .Q( u0_uk_K_r5_22 ) , .QN( u0_uk_n394 ) );
  DFF_X1 u0_uk_K_r5_reg_23 (.CK( clk ) , .D( u0_uk_K_r4_23 ) , .Q( u0_uk_K_r5_23 ) );
  DFF_X1 u0_uk_K_r5_reg_24 (.CK( clk ) , .D( u0_uk_K_r4_24 ) , .Q( u0_uk_K_r5_24 ) , .QN( u0_uk_n393 ) );
  DFF_X1 u0_uk_K_r5_reg_25 (.CK( clk ) , .D( u0_uk_K_r4_25 ) , .Q( u0_uk_K_r5_25 ) , .QN( u0_uk_n392 ) );
  DFF_X1 u0_uk_K_r5_reg_26 (.CK( clk ) , .D( u0_uk_K_r4_26 ) , .Q( u0_uk_K_r5_26 ) );
  DFF_X1 u0_uk_K_r5_reg_27 (.CK( clk ) , .D( u0_uk_K_r4_27 ) , .Q( u0_uk_K_r5_27 ) , .QN( u0_uk_n390 ) );
  DFF_X1 u0_uk_K_r5_reg_28 (.CK( clk ) , .D( u0_uk_K_r4_28 ) , .Q( u0_uk_K_r5_28 ) , .QN( u0_uk_n389 ) );
  DFF_X1 u0_uk_K_r5_reg_29 (.CK( clk ) , .D( u0_uk_K_r4_29 ) , .Q( u0_uk_K_r5_29 ) , .QN( u0_uk_n388 ) );
  DFF_X1 u0_uk_K_r5_reg_3 (.CK( clk ) , .D( u0_uk_K_r4_3 ) , .Q( u0_uk_K_r5_3 ) , .QN( u0_uk_n405 ) );
  DFF_X1 u0_uk_K_r5_reg_30 (.CK( clk ) , .D( u0_uk_K_r4_30 ) , .Q( u0_uk_K_r5_30 ) , .QN( u0_uk_n387 ) );
  DFF_X1 u0_uk_K_r5_reg_31 (.CK( clk ) , .D( u0_uk_K_r4_31 ) , .Q( u0_uk_K_r5_31 ) );
  DFF_X1 u0_uk_K_r5_reg_32 (.CK( clk ) , .D( u0_uk_K_r4_32 ) , .Q( u0_uk_K_r5_32 ) );
  DFF_X1 u0_uk_K_r5_reg_33 (.CK( clk ) , .D( u0_uk_K_r4_33 ) , .Q( u0_uk_K_r5_33 ) , .QN( u0_uk_n384 ) );
  DFF_X1 u0_uk_K_r5_reg_34 (.CK( clk ) , .D( u0_uk_K_r4_34 ) , .Q( u0_uk_K_r5_34 ) , .QN( u0_uk_n383 ) );
  DFF_X1 u0_uk_K_r5_reg_35 (.CK( clk ) , .D( u0_uk_K_r4_35 ) , .Q( u0_uk_K_r5_35 ) , .QN( u0_uk_n381 ) );
  DFF_X1 u0_uk_K_r5_reg_36 (.CK( clk ) , .D( u0_uk_K_r4_36 ) , .Q( u0_uk_K_r5_36 ) , .QN( u0_uk_n380 ) );
  DFF_X1 u0_uk_K_r5_reg_37 (.CK( clk ) , .D( u0_uk_K_r4_37 ) , .Q( u0_uk_K_r5_37 ) );
  DFF_X1 u0_uk_K_r5_reg_38 (.CK( clk ) , .D( u0_uk_K_r4_38 ) , .Q( u0_uk_K_r5_38 ) , .QN( u0_uk_n378 ) );
  DFF_X1 u0_uk_K_r5_reg_39 (.CK( clk ) , .D( u0_uk_K_r4_39 ) , .Q( u0_uk_K_r5_39 ) );
  DFF_X1 u0_uk_K_r5_reg_4 (.CK( clk ) , .D( u0_uk_K_r4_4 ) , .Q( u0_uk_K_r5_4 ) );
  DFF_X1 u0_uk_K_r5_reg_40 (.CK( clk ) , .D( u0_uk_K_r4_40 ) , .Q( u0_uk_K_r5_40 ) );
  DFF_X1 u0_uk_K_r5_reg_41 (.CK( clk ) , .D( u0_uk_K_r4_41 ) , .Q( u0_uk_K_r5_41 ) );
  DFF_X1 u0_uk_K_r5_reg_42 (.CK( clk ) , .D( u0_uk_K_r4_42 ) , .Q( u0_uk_K_r5_42 ) , .QN( u0_uk_n374 ) );
  DFF_X1 u0_uk_K_r5_reg_43 (.CK( clk ) , .D( u0_uk_K_r4_43 ) , .Q( u0_uk_K_r5_43 ) );
  DFF_X1 u0_uk_K_r5_reg_44 (.CK( clk ) , .D( u0_uk_K_r4_44 ) , .Q( u0_uk_K_r5_44 ) , .QN( u0_uk_n372 ) );
  DFF_X1 u0_uk_K_r5_reg_45 (.CK( clk ) , .D( u0_uk_K_r4_45 ) , .Q( u0_uk_K_r5_45 ) );
  DFF_X1 u0_uk_K_r5_reg_46 (.CK( clk ) , .D( u0_uk_K_r4_46 ) , .Q( u0_uk_K_r5_46 ) , .QN( u0_uk_n371 ) );
  DFF_X1 u0_uk_K_r5_reg_47 (.CK( clk ) , .D( u0_uk_K_r4_47 ) , .Q( u0_uk_K_r5_47 ) , .QN( u0_uk_n370 ) );
  DFF_X1 u0_uk_K_r5_reg_48 (.CK( clk ) , .D( u0_uk_K_r4_48 ) , .Q( u0_uk_K_r5_48 ) );
  DFF_X1 u0_uk_K_r5_reg_49 (.CK( clk ) , .D( u0_uk_K_r4_49 ) , .Q( u0_uk_K_r5_49 ) , .QN( u0_uk_n368 ) );
  DFF_X1 u0_uk_K_r5_reg_5 (.CK( clk ) , .D( u0_uk_K_r4_5 ) , .Q( u0_uk_K_r5_5 ) );
  DFF_X1 u0_uk_K_r5_reg_50 (.CK( clk ) , .D( u0_uk_K_r4_50 ) , .Q( u0_uk_K_r5_50 ) , .QN( u0_uk_n367 ) );
  DFF_X1 u0_uk_K_r5_reg_51 (.CK( clk ) , .D( u0_uk_K_r4_51 ) , .Q( u0_uk_K_r5_51 ) );
  DFF_X1 u0_uk_K_r5_reg_52 (.CK( clk ) , .D( u0_uk_K_r4_52 ) , .Q( u0_uk_K_r5_52 ) , .QN( u0_uk_n365 ) );
  DFF_X1 u0_uk_K_r5_reg_53 (.CK( clk ) , .D( u0_uk_K_r4_53 ) , .Q( u0_uk_K_r5_53 ) , .QN( u0_uk_n364 ) );
  DFF_X1 u0_uk_K_r5_reg_54 (.CK( clk ) , .D( u0_uk_K_r4_54 ) , .Q( u0_uk_K_r5_54 ) , .QN( u0_uk_n362 ) );
  DFF_X1 u0_uk_K_r5_reg_55 (.CK( clk ) , .D( u0_uk_K_r4_55 ) , .Q( u0_uk_K_r5_55 ) , .QN( u0_uk_n361 ) );
  DFF_X1 u0_uk_K_r5_reg_6 (.CK( clk ) , .D( u0_uk_K_r4_6 ) , .Q( u0_uk_K_r5_6 ) , .QN( u0_uk_n404 ) );
  DFF_X1 u0_uk_K_r5_reg_7 (.CK( clk ) , .D( u0_uk_K_r4_7 ) , .Q( u0_uk_K_r5_7 ) , .QN( u0_uk_n403 ) );
  DFF_X1 u0_uk_K_r5_reg_8 (.CK( clk ) , .D( u0_uk_K_r4_8 ) , .Q( u0_uk_K_r5_8 ) );
  DFF_X1 u0_uk_K_r5_reg_9 (.CK( clk ) , .D( u0_uk_K_r4_9 ) , .Q( u0_uk_K_r5_9 ) , .QN( u0_uk_n402 ) );
  DFF_X1 u0_uk_K_r6_reg_0 (.CK( clk ) , .D( u0_uk_K_r5_0 ) , .Q( u0_uk_K_r6_0 ) );
  DFF_X1 u0_uk_K_r6_reg_1 (.CK( clk ) , .D( u0_uk_K_r5_1 ) , .Q( u0_uk_K_r6_1 ) , .QN( u0_uk_n360 ) );
  DFF_X1 u0_uk_K_r6_reg_10 (.CK( clk ) , .D( u0_uk_K_r5_10 ) , .Q( u0_uk_K_r6_10 ) );
  DFF_X1 u0_uk_K_r6_reg_11 (.CK( clk ) , .D( u0_uk_K_r5_11 ) , .Q( u0_uk_K_r6_11 ) , .QN( u0_uk_n352 ) );
  DFF_X1 u0_uk_K_r6_reg_12 (.CK( clk ) , .D( u0_uk_K_r5_12 ) , .Q( u0_uk_K_r6_12 ) , .QN( u0_uk_n351 ) );
  DFF_X1 u0_uk_K_r6_reg_13 (.CK( clk ) , .D( u0_uk_K_r5_13 ) , .Q( u0_uk_K_r6_13 ) , .QN( u0_uk_n350 ) );
  DFF_X1 u0_uk_K_r6_reg_14 (.CK( clk ) , .D( u0_uk_K_r5_14 ) , .Q( u0_uk_K_r6_14 ) );
  DFF_X1 u0_uk_K_r6_reg_15 (.CK( clk ) , .D( u0_uk_K_r5_15 ) , .Q( u0_uk_K_r6_15 ) , .QN( u0_uk_n348 ) );
  DFF_X1 u0_uk_K_r6_reg_16 (.CK( clk ) , .D( u0_uk_K_r5_16 ) , .Q( u0_uk_K_r6_16 ) , .QN( u0_uk_n347 ) );
  DFF_X1 u0_uk_K_r6_reg_17 (.CK( clk ) , .D( u0_uk_K_r5_17 ) , .Q( u0_uk_K_r6_17 ) , .QN( u0_uk_n345 ) );
  DFF_X1 u0_uk_K_r6_reg_18 (.CK( clk ) , .D( u0_uk_K_r5_18 ) , .Q( u0_uk_K_r6_18 ) , .QN( u0_uk_n344 ) );
  DFF_X1 u0_uk_K_r6_reg_19 (.CK( clk ) , .D( u0_uk_K_r5_19 ) , .Q( u0_uk_K_r6_19 ) );
  DFF_X1 u0_uk_K_r6_reg_2 (.CK( clk ) , .D( u0_uk_K_r5_2 ) , .Q( u0_uk_K_r6_2 ) , .QN( u0_uk_n359 ) );
  DFF_X1 u0_uk_K_r6_reg_20 (.CK( clk ) , .D( u0_uk_K_r5_20 ) , .Q( u0_uk_K_r6_20 ) , .QN( u0_uk_n343 ) );
  DFF_X1 u0_uk_K_r6_reg_21 (.CK( clk ) , .D( u0_uk_K_r5_21 ) , .Q( u0_uk_K_r6_21 ) );
  DFF_X1 u0_uk_K_r6_reg_22 (.CK( clk ) , .D( u0_uk_K_r5_22 ) , .Q( u0_uk_K_r6_22 ) );
  DFF_X1 u0_uk_K_r6_reg_23 (.CK( clk ) , .D( u0_uk_K_r5_23 ) , .Q( u0_uk_K_r6_23 ) , .QN( u0_uk_n341 ) );
  DFF_X1 u0_uk_K_r6_reg_24 (.CK( clk ) , .D( u0_uk_K_r5_24 ) , .Q( u0_uk_K_r6_24 ) , .QN( u0_uk_n340 ) );
  DFF_X1 u0_uk_K_r6_reg_25 (.CK( clk ) , .D( u0_uk_K_r5_25 ) , .Q( u0_uk_K_r6_25 ) , .QN( u0_uk_n339 ) );
  DFF_X1 u0_uk_K_r6_reg_26 (.CK( clk ) , .D( u0_uk_K_r5_26 ) , .Q( u0_uk_K_r6_26 ) );
  DFF_X1 u0_uk_K_r6_reg_27 (.CK( clk ) , .D( u0_uk_K_r5_27 ) , .Q( u0_uk_K_r6_27 ) );
  DFF_X1 u0_uk_K_r6_reg_28 (.CK( clk ) , .D( u0_uk_K_r5_28 ) , .Q( u0_uk_K_r6_28 ) );
  DFF_X1 u0_uk_K_r6_reg_29 (.CK( clk ) , .D( u0_uk_K_r5_29 ) , .Q( u0_uk_K_r6_29 ) );
  DFF_X1 u0_uk_K_r6_reg_3 (.CK( clk ) , .D( u0_uk_K_r5_3 ) , .Q( u0_uk_K_r6_3 ) );
  DFF_X1 u0_uk_K_r6_reg_30 (.CK( clk ) , .D( u0_uk_K_r5_30 ) , .Q( u0_uk_K_r6_30 ) );
  DFF_X1 u0_uk_K_r6_reg_31 (.CK( clk ) , .D( u0_uk_K_r5_31 ) , .Q( u0_uk_K_r6_31 ) );
  DFF_X1 u0_uk_K_r6_reg_32 (.CK( clk ) , .D( u0_uk_K_r5_32 ) , .Q( u0_uk_K_r6_32 ) , .QN( u0_uk_n337 ) );
  DFF_X1 u0_uk_K_r6_reg_33 (.CK( clk ) , .D( u0_uk_K_r5_33 ) , .Q( u0_uk_K_r6_33 ) , .QN( u0_uk_n336 ) );
  DFF_X1 u0_uk_K_r6_reg_34 (.CK( clk ) , .D( u0_uk_K_r5_34 ) , .Q( u0_uk_K_r6_34 ) );
  DFF_X1 u0_uk_K_r6_reg_35 (.CK( clk ) , .D( u0_uk_K_r5_35 ) , .Q( u0_uk_K_r6_35 ) , .QN( u0_uk_n334 ) );
  DFF_X1 u0_uk_K_r6_reg_36 (.CK( clk ) , .D( u0_uk_K_r5_36 ) , .Q( u0_uk_K_r6_36 ) , .QN( u0_uk_n333 ) );
  DFF_X1 u0_uk_K_r6_reg_37 (.CK( clk ) , .D( u0_uk_K_r5_37 ) , .Q( u0_uk_K_r6_37 ) );
  DFF_X1 u0_uk_K_r6_reg_38 (.CK( clk ) , .D( u0_uk_K_r5_38 ) , .Q( u0_uk_K_r6_38 ) , .QN( u0_uk_n332 ) );
  DFF_X1 u0_uk_K_r6_reg_39 (.CK( clk ) , .D( u0_uk_K_r5_39 ) , .Q( u0_uk_K_r6_39 ) , .QN( u0_uk_n331 ) );
  DFF_X1 u0_uk_K_r6_reg_4 (.CK( clk ) , .D( u0_uk_K_r5_4 ) , .Q( u0_uk_K_r6_4 ) , .QN( u0_uk_n358 ) );
  DFF_X1 u0_uk_K_r6_reg_40 (.CK( clk ) , .D( u0_uk_K_r5_40 ) , .Q( u0_uk_K_r6_40 ) , .QN( u0_uk_n330 ) );
  DFF_X1 u0_uk_K_r6_reg_41 (.CK( clk ) , .D( u0_uk_K_r5_41 ) , .Q( u0_uk_K_r6_41 ) , .QN( u0_uk_n329 ) );
  DFF_X1 u0_uk_K_r6_reg_42 (.CK( clk ) , .D( u0_uk_K_r5_42 ) , .Q( u0_uk_K_r6_42 ) , .QN( u0_uk_n328 ) );
  DFF_X1 u0_uk_K_r6_reg_43 (.CK( clk ) , .D( u0_uk_K_r5_43 ) , .Q( u0_uk_K_r6_43 ) , .QN( u0_uk_n327 ) );
  DFF_X1 u0_uk_K_r6_reg_44 (.CK( clk ) , .D( u0_uk_K_r5_44 ) , .Q( u0_uk_K_r6_44 ) , .QN( u0_uk_n326 ) );
  DFF_X1 u0_uk_K_r6_reg_45 (.CK( clk ) , .D( u0_uk_K_r5_45 ) , .Q( u0_uk_K_r6_45 ) , .QN( u0_uk_n325 ) );
  DFF_X1 u0_uk_K_r6_reg_46 (.CK( clk ) , .D( u0_uk_K_r5_46 ) , .Q( u0_uk_K_r6_46 ) );
  DFF_X1 u0_uk_K_r6_reg_47 (.CK( clk ) , .D( u0_uk_K_r5_47 ) , .Q( u0_uk_K_r6_47 ) , .QN( u0_uk_n324 ) );
  DFF_X1 u0_uk_K_r6_reg_48 (.CK( clk ) , .D( u0_uk_K_r5_48 ) , .Q( u0_uk_K_r6_48 ) , .QN( u0_uk_n323 ) );
  DFF_X1 u0_uk_K_r6_reg_49 (.CK( clk ) , .D( u0_uk_K_r5_49 ) , .Q( u0_uk_K_r6_49 ) , .QN( u0_uk_n322 ) );
  DFF_X1 u0_uk_K_r6_reg_5 (.CK( clk ) , .D( u0_uk_K_r5_5 ) , .Q( u0_uk_K_r6_5 ) , .QN( u0_uk_n357 ) );
  DFF_X1 u0_uk_K_r6_reg_50 (.CK( clk ) , .D( u0_uk_K_r5_50 ) , .Q( u0_uk_K_r6_50 ) , .QN( u0_uk_n321 ) );
  DFF_X1 u0_uk_K_r6_reg_51 (.CK( clk ) , .D( u0_uk_K_r5_51 ) , .Q( u0_uk_K_r6_51 ) );
  DFF_X1 u0_uk_K_r6_reg_52 (.CK( clk ) , .D( u0_uk_K_r5_52 ) , .Q( u0_uk_K_r6_52 ) , .QN( u0_uk_n320 ) );
  DFF_X1 u0_uk_K_r6_reg_53 (.CK( clk ) , .D( u0_uk_K_r5_53 ) , .Q( u0_uk_K_r6_53 ) );
  DFF_X1 u0_uk_K_r6_reg_54 (.CK( clk ) , .D( u0_uk_K_r5_54 ) , .Q( u0_uk_K_r6_54 ) , .QN( u0_uk_n318 ) );
  DFF_X1 u0_uk_K_r6_reg_55 (.CK( clk ) , .D( u0_uk_K_r5_55 ) , .Q( u0_uk_K_r6_55 ) );
  DFF_X1 u0_uk_K_r6_reg_6 (.CK( clk ) , .D( u0_uk_K_r5_6 ) , .Q( u0_uk_K_r6_6 ) , .QN( u0_uk_n356 ) );
  DFF_X1 u0_uk_K_r6_reg_7 (.CK( clk ) , .D( u0_uk_K_r5_7 ) , .Q( u0_uk_K_r6_7 ) );
  DFF_X1 u0_uk_K_r6_reg_8 (.CK( clk ) , .D( u0_uk_K_r5_8 ) , .Q( u0_uk_K_r6_8 ) , .QN( u0_uk_n355 ) );
  DFF_X1 u0_uk_K_r6_reg_9 (.CK( clk ) , .D( u0_uk_K_r5_9 ) , .Q( u0_uk_K_r6_9 ) , .QN( u0_uk_n354 ) );
  DFF_X1 u0_uk_K_r7_reg_0 (.CK( clk ) , .D( u0_uk_K_r6_0 ) , .Q( u0_uk_K_r7_0 ) );
  DFF_X1 u0_uk_K_r7_reg_1 (.CK( clk ) , .D( u0_uk_K_r6_1 ) , .Q( u0_uk_K_r7_1 ) , .QN( u0_uk_n317 ) );
  DFF_X1 u0_uk_K_r7_reg_10 (.CK( clk ) , .D( u0_uk_K_r6_10 ) , .Q( u0_uk_K_r7_10 ) , .QN( u0_uk_n311 ) );
  DFF_X1 u0_uk_K_r7_reg_11 (.CK( clk ) , .D( u0_uk_K_r6_11 ) , .Q( u0_uk_K_r7_11 ) , .QN( u0_uk_n310 ) );
  DFF_X1 u0_uk_K_r7_reg_12 (.CK( clk ) , .D( u0_uk_K_r6_12 ) , .Q( u0_uk_K_r7_12 ) , .QN( u0_uk_n309 ) );
  DFF_X1 u0_uk_K_r7_reg_13 (.CK( clk ) , .D( u0_uk_K_r6_13 ) , .Q( u0_uk_K_r7_13 ) );
  DFF_X1 u0_uk_K_r7_reg_14 (.CK( clk ) , .D( u0_uk_K_r6_14 ) , .Q( u0_uk_K_r7_14 ) , .QN( u0_uk_n307 ) );
  DFF_X1 u0_uk_K_r7_reg_15 (.CK( clk ) , .D( u0_uk_K_r6_15 ) , .Q( u0_uk_K_r7_15 ) );
  DFF_X1 u0_uk_K_r7_reg_16 (.CK( clk ) , .D( u0_uk_K_r6_16 ) , .Q( u0_uk_K_r7_16 ) );
  DFF_X1 u0_uk_K_r7_reg_17 (.CK( clk ) , .D( u0_uk_K_r6_17 ) , .Q( u0_uk_K_r7_17 ) , .QN( u0_uk_n304 ) );
  DFF_X1 u0_uk_K_r7_reg_18 (.CK( clk ) , .D( u0_uk_K_r6_18 ) , .Q( u0_uk_K_r7_18 ) , .QN( u0_uk_n303 ) );
  DFF_X1 u0_uk_K_r7_reg_19 (.CK( clk ) , .D( u0_uk_K_r6_19 ) , .Q( u0_uk_K_r7_19 ) , .QN( u0_uk_n302 ) );
  DFF_X1 u0_uk_K_r7_reg_2 (.CK( clk ) , .D( u0_uk_K_r6_2 ) , .Q( u0_uk_K_r7_2 ) , .QN( u0_uk_n316 ) );
  DFF_X1 u0_uk_K_r7_reg_20 (.CK( clk ) , .D( u0_uk_K_r6_20 ) , .Q( u0_uk_K_r7_20 ) );
  DFF_X1 u0_uk_K_r7_reg_21 (.CK( clk ) , .D( u0_uk_K_r6_21 ) , .Q( u0_uk_K_r7_21 ) , .QN( u0_uk_n300 ) );
  DFF_X1 u0_uk_K_r7_reg_22 (.CK( clk ) , .D( u0_uk_K_r6_22 ) , .Q( u0_uk_K_r7_22 ) );
  DFF_X1 u0_uk_K_r7_reg_23 (.CK( clk ) , .D( u0_uk_K_r6_23 ) , .Q( u0_uk_K_r7_23 ) );
  DFF_X1 u0_uk_K_r7_reg_24 (.CK( clk ) , .D( u0_uk_K_r6_24 ) , .Q( u0_uk_K_r7_24 ) , .QN( u0_uk_n296 ) );
  DFF_X1 u0_uk_K_r7_reg_25 (.CK( clk ) , .D( u0_uk_K_r6_25 ) , .Q( u0_uk_K_r7_25 ) , .QN( u0_uk_n295 ) );
  DFF_X1 u0_uk_K_r7_reg_26 (.CK( clk ) , .D( u0_uk_K_r6_26 ) , .Q( u0_uk_K_r7_26 ) );
  DFF_X1 u0_uk_K_r7_reg_27 (.CK( clk ) , .D( u0_uk_K_r6_27 ) , .Q( u0_uk_K_r7_27 ) );
  DFF_X1 u0_uk_K_r7_reg_28 (.CK( clk ) , .D( u0_uk_K_r6_28 ) , .Q( u0_uk_K_r7_28 ) , .QN( u0_uk_n293 ) );
  DFF_X1 u0_uk_K_r7_reg_29 (.CK( clk ) , .D( u0_uk_K_r6_29 ) , .Q( u0_uk_K_r7_29 ) );
  DFF_X1 u0_uk_K_r7_reg_3 (.CK( clk ) , .D( u0_uk_K_r6_3 ) , .Q( u0_uk_K_r7_3 ) , .QN( u0_uk_n315 ) );
  DFF_X1 u0_uk_K_r7_reg_30 (.CK( clk ) , .D( u0_uk_K_r6_30 ) , .Q( u0_uk_K_r7_30 ) );
  DFF_X1 u0_uk_K_r7_reg_31 (.CK( clk ) , .D( u0_uk_K_r6_31 ) , .Q( u0_uk_K_r7_31 ) );
  DFF_X1 u0_uk_K_r7_reg_32 (.CK( clk ) , .D( u0_uk_K_r6_32 ) , .Q( u0_uk_K_r7_32 ) );
  DFF_X1 u0_uk_K_r7_reg_33 (.CK( clk ) , .D( u0_uk_K_r6_33 ) , .Q( u0_uk_K_r7_33 ) , .QN( u0_uk_n290 ) );
  DFF_X1 u0_uk_K_r7_reg_34 (.CK( clk ) , .D( u0_uk_K_r6_34 ) , .Q( u0_uk_K_r7_34 ) );
  DFF_X1 u0_uk_K_r7_reg_35 (.CK( clk ) , .D( u0_uk_K_r6_35 ) , .Q( u0_uk_K_r7_35 ) , .QN( u0_uk_n289 ) );
  DFF_X1 u0_uk_K_r7_reg_36 (.CK( clk ) , .D( u0_uk_K_r6_36 ) , .Q( u0_uk_K_r7_36 ) , .QN( u0_uk_n288 ) );
  DFF_X1 u0_uk_K_r7_reg_37 (.CK( clk ) , .D( u0_uk_K_r6_37 ) , .Q( u0_uk_K_r7_37 ) );
  DFF_X1 u0_uk_K_r7_reg_38 (.CK( clk ) , .D( u0_uk_K_r6_38 ) , .Q( u0_uk_K_r7_38 ) , .QN( u0_uk_n287 ) );
  DFF_X1 u0_uk_K_r7_reg_39 (.CK( clk ) , .D( u0_uk_K_r6_39 ) , .Q( u0_uk_K_r7_39 ) );
  DFF_X1 u0_uk_K_r7_reg_4 (.CK( clk ) , .D( u0_uk_K_r6_4 ) , .Q( u0_uk_K_r7_4 ) , .QN( u0_uk_n314 ) );
  DFF_X1 u0_uk_K_r7_reg_40 (.CK( clk ) , .D( u0_uk_K_r6_40 ) , .Q( u0_uk_K_r7_40 ) , .QN( u0_uk_n285 ) );
  DFF_X1 u0_uk_K_r7_reg_41 (.CK( clk ) , .D( u0_uk_K_r6_41 ) , .Q( u0_uk_K_r7_41 ) , .QN( u0_uk_n284 ) );
  DFF_X1 u0_uk_K_r7_reg_42 (.CK( clk ) , .D( u0_uk_K_r6_42 ) , .Q( u0_uk_K_r7_42 ) , .QN( u0_uk_n283 ) );
  DFF_X1 u0_uk_K_r7_reg_43 (.CK( clk ) , .D( u0_uk_K_r6_43 ) , .Q( u0_uk_K_r7_43 ) , .QN( u0_uk_n282 ) );
  DFF_X1 u0_uk_K_r7_reg_44 (.CK( clk ) , .D( u0_uk_K_r6_44 ) , .Q( u0_uk_K_r7_44 ) , .QN( u0_uk_n281 ) );
  DFF_X1 u0_uk_K_r7_reg_45 (.CK( clk ) , .D( u0_uk_K_r6_45 ) , .Q( u0_uk_K_r7_45 ) , .QN( u0_uk_n280 ) );
  DFF_X1 u0_uk_K_r7_reg_46 (.CK( clk ) , .D( u0_uk_K_r6_46 ) , .Q( u0_uk_K_r7_46 ) );
  DFF_X1 u0_uk_K_r7_reg_47 (.CK( clk ) , .D( u0_uk_K_r6_47 ) , .Q( u0_uk_K_r7_47 ) , .QN( u0_uk_n278 ) );
  DFF_X1 u0_uk_K_r7_reg_48 (.CK( clk ) , .D( u0_uk_K_r6_48 ) , .Q( u0_uk_K_r7_48 ) );
  DFF_X1 u0_uk_K_r7_reg_49 (.CK( clk ) , .D( u0_uk_K_r6_49 ) , .Q( u0_uk_K_r7_49 ) , .QN( u0_uk_n276 ) );
  DFF_X1 u0_uk_K_r7_reg_5 (.CK( clk ) , .D( u0_uk_K_r6_5 ) , .Q( u0_uk_K_r7_5 ) );
  DFF_X1 u0_uk_K_r7_reg_50 (.CK( clk ) , .D( u0_uk_K_r6_50 ) , .Q( u0_uk_K_r7_50 ) , .QN( u0_uk_n275 ) );
  DFF_X1 u0_uk_K_r7_reg_51 (.CK( clk ) , .D( u0_uk_K_r6_51 ) , .Q( u0_uk_K_r7_51 ) , .QN( u0_uk_n274 ) );
  DFF_X1 u0_uk_K_r7_reg_52 (.CK( clk ) , .D( u0_uk_K_r6_52 ) , .Q( u0_uk_K_r7_52 ) , .QN( u0_uk_n273 ) );
  DFF_X1 u0_uk_K_r7_reg_53 (.CK( clk ) , .D( u0_uk_K_r6_53 ) , .Q( u0_uk_K_r7_53 ) );
  DFF_X1 u0_uk_K_r7_reg_54 (.CK( clk ) , .D( u0_uk_K_r6_54 ) , .Q( u0_uk_K_r7_54 ) , .QN( u0_uk_n272 ) );
  DFF_X1 u0_uk_K_r7_reg_55 (.CK( clk ) , .D( u0_uk_K_r6_55 ) , .Q( u0_uk_K_r7_55 ) );
  DFF_X1 u0_uk_K_r7_reg_6 (.CK( clk ) , .D( u0_uk_K_r6_6 ) , .Q( u0_uk_K_r7_6 ) );
  DFF_X1 u0_uk_K_r7_reg_7 (.CK( clk ) , .D( u0_uk_K_r6_7 ) , .Q( u0_uk_K_r7_7 ) );
  DFF_X1 u0_uk_K_r7_reg_8 (.CK( clk ) , .D( u0_uk_K_r6_8 ) , .Q( u0_uk_K_r7_8 ) );
  DFF_X1 u0_uk_K_r7_reg_9 (.CK( clk ) , .D( u0_uk_K_r6_9 ) , .Q( u0_uk_K_r7_9 ) );
  DFF_X1 u0_uk_K_r8_reg_0 (.CK( clk ) , .D( u0_uk_K_r7_0 ) , .Q( u0_uk_K_r8_0 ) , .QN( u0_uk_n270 ) );
  DFF_X1 u0_uk_K_r8_reg_1 (.CK( clk ) , .D( u0_uk_K_r7_1 ) , .Q( u0_uk_K_r8_1 ) , .QN( u0_uk_n269 ) );
  DFF_X1 u0_uk_K_r8_reg_10 (.CK( clk ) , .D( u0_uk_K_r7_10 ) , .Q( u0_uk_K_r8_10 ) );
  DFF_X1 u0_uk_K_r8_reg_11 (.CK( clk ) , .D( u0_uk_K_r7_11 ) , .Q( u0_uk_K_r8_11 ) , .QN( u0_uk_n263 ) );
  DFF_X1 u0_uk_K_r8_reg_12 (.CK( clk ) , .D( u0_uk_K_r7_12 ) , .Q( u0_uk_K_r8_12 ) , .QN( u0_uk_n262 ) );
  DFF_X1 u0_uk_K_r8_reg_13 (.CK( clk ) , .D( u0_uk_K_r7_13 ) , .Q( u0_uk_K_r8_13 ) );
  DFF_X1 u0_uk_K_r8_reg_14 (.CK( clk ) , .D( u0_uk_K_r7_14 ) , .Q( u0_uk_K_r8_14 ) , .QN( u0_uk_n261 ) );
  DFF_X1 u0_uk_K_r8_reg_15 (.CK( clk ) , .D( u0_uk_K_r7_15 ) , .Q( u0_uk_K_r8_15 ) , .QN( u0_uk_n260 ) );
  DFF_X1 u0_uk_K_r8_reg_16 (.CK( clk ) , .D( u0_uk_K_r7_16 ) , .Q( u0_uk_K_r8_16 ) );
  DFF_X1 u0_uk_K_r8_reg_17 (.CK( clk ) , .D( u0_uk_K_r7_17 ) , .Q( u0_uk_K_r8_17 ) );
  DFF_X1 u0_uk_K_r8_reg_18 (.CK( clk ) , .D( u0_uk_K_r7_18 ) , .Q( u0_uk_K_r8_18 ) , .QN( u0_uk_n259 ) );
  DFF_X1 u0_uk_K_r8_reg_19 (.CK( clk ) , .D( u0_uk_K_r7_19 ) , .Q( u0_uk_K_r8_19 ) );
  DFF_X1 u0_uk_K_r8_reg_2 (.CK( clk ) , .D( u0_uk_K_r7_2 ) , .Q( u0_uk_K_r8_2 ) );
  DFF_X1 u0_uk_K_r8_reg_20 (.CK( clk ) , .D( u0_uk_K_r7_20 ) , .Q( u0_uk_K_r8_20 ) , .QN( u0_uk_n258 ) );
  DFF_X1 u0_uk_K_r8_reg_21 (.CK( clk ) , .D( u0_uk_K_r7_21 ) , .Q( u0_uk_K_r8_21 ) );
  DFF_X1 u0_uk_K_r8_reg_22 (.CK( clk ) , .D( u0_uk_K_r7_22 ) , .Q( u0_uk_K_r8_22 ) );
  DFF_X1 u0_uk_K_r8_reg_23 (.CK( clk ) , .D( u0_uk_K_r7_23 ) , .Q( u0_uk_K_r8_23 ) , .QN( u0_uk_n256 ) );
  DFF_X1 u0_uk_K_r8_reg_24 (.CK( clk ) , .D( u0_uk_K_r7_24 ) , .Q( u0_uk_K_r8_24 ) , .QN( u0_uk_n255 ) );
  DFF_X1 u0_uk_K_r8_reg_25 (.CK( clk ) , .D( u0_uk_K_r7_25 ) , .Q( u0_uk_K_r8_25 ) , .QN( u0_uk_n254 ) );
  DFF_X1 u0_uk_K_r8_reg_26 (.CK( clk ) , .D( u0_uk_K_r7_26 ) , .Q( u0_uk_K_r8_26 ) , .QN( u0_uk_n253 ) );
  DFF_X1 u0_uk_K_r8_reg_27 (.CK( clk ) , .D( u0_uk_K_r7_27 ) , .Q( u0_uk_K_r8_27 ) );
  DFF_X1 u0_uk_K_r8_reg_28 (.CK( clk ) , .D( u0_uk_K_r7_28 ) , .Q( u0_uk_K_r8_28 ) );
  DFF_X1 u0_uk_K_r8_reg_29 (.CK( clk ) , .D( u0_uk_K_r7_29 ) , .Q( u0_uk_K_r8_29 ) , .QN( u0_uk_n249 ) );
  DFF_X1 u0_uk_K_r8_reg_3 (.CK( clk ) , .D( u0_uk_K_r7_3 ) , .Q( u0_uk_K_r8_3 ) , .QN( u0_uk_n268 ) );
  DFF_X1 u0_uk_K_r8_reg_30 (.CK( clk ) , .D( u0_uk_K_r7_30 ) , .Q( u0_uk_K_r8_30 ) , .QN( u0_uk_n248 ) );
  DFF_X1 u0_uk_K_r8_reg_31 (.CK( clk ) , .D( u0_uk_K_r7_31 ) , .Q( u0_uk_K_r8_31 ) , .QN( u0_uk_n247 ) );
  DFF_X1 u0_uk_K_r8_reg_32 (.CK( clk ) , .D( u0_uk_K_r7_32 ) , .Q( u0_uk_K_r8_32 ) );
  DFF_X1 u0_uk_K_r8_reg_33 (.CK( clk ) , .D( u0_uk_K_r7_33 ) , .Q( u0_uk_K_r8_33 ) , .QN( u0_uk_n246 ) );
  DFF_X1 u0_uk_K_r8_reg_34 (.CK( clk ) , .D( u0_uk_K_r7_34 ) , .Q( u0_uk_K_r8_34 ) , .QN( u0_uk_n245 ) );
  DFF_X1 u0_uk_K_r8_reg_35 (.CK( clk ) , .D( u0_uk_K_r7_35 ) , .Q( u0_uk_K_r8_35 ) , .QN( u0_uk_n244 ) );
  DFF_X1 u0_uk_K_r8_reg_36 (.CK( clk ) , .D( u0_uk_K_r7_36 ) , .Q( u0_uk_K_r8_36 ) , .QN( u0_uk_n243 ) );
  DFF_X1 u0_uk_K_r8_reg_37 (.CK( clk ) , .D( u0_uk_K_r7_37 ) , .Q( u0_uk_K_r8_37 ) );
  DFF_X1 u0_uk_K_r8_reg_38 (.CK( clk ) , .D( u0_uk_K_r7_38 ) , .Q( u0_uk_K_r8_38 ) , .QN( u0_uk_n241 ) );
  DFF_X1 u0_uk_K_r8_reg_39 (.CK( clk ) , .D( u0_uk_K_r7_39 ) , .Q( u0_uk_K_r8_39 ) , .QN( u0_uk_n239 ) );
  DFF_X1 u0_uk_K_r8_reg_4 (.CK( clk ) , .D( u0_uk_K_r7_4 ) , .Q( u0_uk_K_r8_4 ) , .QN( u0_uk_n267 ) );
  DFF_X1 u0_uk_K_r8_reg_40 (.CK( clk ) , .D( u0_uk_K_r7_40 ) , .Q( u0_uk_K_r8_40 ) );
  DFF_X1 u0_uk_K_r8_reg_41 (.CK( clk ) , .D( u0_uk_K_r7_41 ) , .Q( u0_uk_K_r8_41 ) );
  DFF_X1 u0_uk_K_r8_reg_42 (.CK( clk ) , .D( u0_uk_K_r7_42 ) , .Q( u0_uk_K_r8_42 ) , .QN( u0_uk_n237 ) );
  DFF_X1 u0_uk_K_r8_reg_43 (.CK( clk ) , .D( u0_uk_K_r7_43 ) , .Q( u0_uk_K_r8_43 ) );
  DFF_X1 u0_uk_K_r8_reg_44 (.CK( clk ) , .D( u0_uk_K_r7_44 ) , .Q( u0_uk_K_r8_44 ) , .QN( u0_uk_n236 ) );
  DFF_X1 u0_uk_K_r8_reg_45 (.CK( clk ) , .D( u0_uk_K_r7_45 ) , .Q( u0_uk_K_r8_45 ) );
  DFF_X1 u0_uk_K_r8_reg_46 (.CK( clk ) , .D( u0_uk_K_r7_46 ) , .Q( u0_uk_K_r8_46 ) , .QN( u0_uk_n235 ) );
  DFF_X1 u0_uk_K_r8_reg_47 (.CK( clk ) , .D( u0_uk_K_r7_47 ) , .Q( u0_uk_K_r8_47 ) , .QN( u0_uk_n234 ) );
  DFF_X1 u0_uk_K_r8_reg_48 (.CK( clk ) , .D( u0_uk_K_r7_48 ) , .Q( u0_uk_K_r8_48 ) );
  DFF_X1 u0_uk_K_r8_reg_49 (.CK( clk ) , .D( u0_uk_K_r7_49 ) , .Q( u0_uk_K_r8_49 ) , .QN( u0_uk_n233 ) );
  DFF_X1 u0_uk_K_r8_reg_5 (.CK( clk ) , .D( u0_uk_K_r7_5 ) , .Q( u0_uk_K_r8_5 ) );
  DFF_X1 u0_uk_K_r8_reg_50 (.CK( clk ) , .D( u0_uk_K_r7_50 ) , .Q( u0_uk_K_r8_50 ) , .QN( u0_uk_n232 ) );
  DFF_X1 u0_uk_K_r8_reg_51 (.CK( clk ) , .D( u0_uk_K_r7_51 ) , .Q( u0_uk_K_r8_51 ) );
  DFF_X1 u0_uk_K_r8_reg_52 (.CK( clk ) , .D( u0_uk_K_r7_52 ) , .Q( u0_uk_K_r8_52 ) );
  DFF_X1 u0_uk_K_r8_reg_53 (.CK( clk ) , .D( u0_uk_K_r7_53 ) , .Q( u0_uk_K_r8_53 ) , .QN( u0_uk_n229 ) );
  DFF_X1 u0_uk_K_r8_reg_54 (.CK( clk ) , .D( u0_uk_K_r7_54 ) , .Q( u0_uk_K_r8_54 ) , .QN( u0_uk_n228 ) );
  DFF_X1 u0_uk_K_r8_reg_55 (.CK( clk ) , .D( u0_uk_K_r7_55 ) , .Q( u0_uk_K_r8_55 ) , .QN( u0_uk_n227 ) );
  DFF_X1 u0_uk_K_r8_reg_6 (.CK( clk ) , .D( u0_uk_K_r7_6 ) , .Q( u0_uk_K_r8_6 ) , .QN( u0_uk_n266 ) );
  DFF_X1 u0_uk_K_r8_reg_7 (.CK( clk ) , .D( u0_uk_K_r7_7 ) , .Q( u0_uk_K_r8_7 ) , .QN( u0_uk_n265 ) );
  DFF_X1 u0_uk_K_r8_reg_8 (.CK( clk ) , .D( u0_uk_K_r7_8 ) , .Q( u0_uk_K_r8_8 ) );
  DFF_X1 u0_uk_K_r8_reg_9 (.CK( clk ) , .D( u0_uk_K_r7_9 ) , .Q( u0_uk_K_r8_9 ) , .QN( u0_uk_n264 ) );
  DFF_X1 u0_uk_K_r9_reg_0 (.CK( clk ) , .D( u0_uk_K_r8_0 ) , .Q( u0_uk_K_r9_0 ) );
  DFF_X1 u0_uk_K_r9_reg_1 (.CK( clk ) , .D( u0_uk_K_r8_1 ) , .Q( u0_uk_K_r9_1 ) , .QN( u0_uk_n226 ) );
  DFF_X1 u0_uk_K_r9_reg_10 (.CK( clk ) , .D( u0_uk_K_r8_10 ) , .Q( u0_uk_K_r9_10 ) );
  DFF_X1 u0_uk_K_r9_reg_11 (.CK( clk ) , .D( u0_uk_K_r8_11 ) , .Q( u0_uk_K_r9_11 ) , .QN( u0_uk_n221 ) );
  DFF_X1 u0_uk_K_r9_reg_12 (.CK( clk ) , .D( u0_uk_K_r8_12 ) , .Q( u0_uk_K_r9_12 ) );
  DFF_X1 u0_uk_K_r9_reg_13 (.CK( clk ) , .D( u0_uk_K_r8_13 ) , .Q( u0_uk_K_r9_13 ) , .QN( u0_uk_n219 ) );
  DFF_X1 u0_uk_K_r9_reg_14 (.CK( clk ) , .D( u0_uk_K_r8_14 ) , .Q( u0_uk_K_r9_14 ) , .QN( u0_uk_n218 ) );
  DFF_X1 u0_uk_K_r9_reg_15 (.CK( clk ) , .D( u0_uk_K_r8_15 ) , .Q( u0_uk_K_r9_15 ) );
  DFF_X1 u0_uk_K_r9_reg_16 (.CK( clk ) , .D( u0_uk_K_r8_16 ) , .Q( u0_uk_K_r9_16 ) , .QN( u0_uk_n216 ) );
  DFF_X1 u0_uk_K_r9_reg_17 (.CK( clk ) , .D( u0_uk_K_r8_17 ) , .Q( u0_uk_K_r9_17 ) , .QN( u0_uk_n215 ) );
  DFF_X1 u0_uk_K_r9_reg_18 (.CK( clk ) , .D( u0_uk_K_r8_18 ) , .Q( u0_uk_K_r9_18 ) );
  DFF_X1 u0_uk_K_r9_reg_19 (.CK( clk ) , .D( u0_uk_K_r8_19 ) , .Q( u0_uk_K_r9_19 ) );
  DFF_X1 u0_uk_K_r9_reg_2 (.CK( clk ) , .D( u0_uk_K_r8_2 ) , .Q( u0_uk_K_r9_2 ) );
  DFF_X1 u0_uk_K_r9_reg_20 (.CK( clk ) , .D( u0_uk_K_r8_20 ) , .Q( u0_uk_K_r9_20 ) , .QN( u0_uk_n212 ) );
  DFF_X1 u0_uk_K_r9_reg_21 (.CK( clk ) , .D( u0_uk_K_r8_21 ) , .Q( u0_uk_K_r9_21 ) , .QN( u0_uk_n211 ) );
  DFF_X1 u0_uk_K_r9_reg_22 (.CK( clk ) , .D( u0_uk_K_r8_22 ) , .Q( u0_uk_K_r9_22 ) , .QN( u0_uk_n210 ) );
  DFF_X1 u0_uk_K_r9_reg_23 (.CK( clk ) , .D( u0_uk_K_r8_23 ) , .Q( u0_uk_K_r9_23 ) );
  DFF_X1 u0_uk_K_r9_reg_24 (.CK( clk ) , .D( u0_uk_K_r8_24 ) , .Q( u0_uk_K_r9_24 ) );
  DFF_X1 u0_uk_K_r9_reg_25 (.CK( clk ) , .D( u0_uk_K_r8_25 ) , .Q( u0_uk_K_r9_25 ) );
  DFF_X1 u0_uk_K_r9_reg_26 (.CK( clk ) , .D( u0_uk_K_r8_26 ) , .Q( u0_uk_K_r9_26 ) , .QN( u0_uk_n206 ) );
  DFF_X1 u0_uk_K_r9_reg_27 (.CK( clk ) , .D( u0_uk_K_r8_27 ) , .Q( u0_uk_K_r9_27 ) );
  DFF_X1 u0_uk_K_r9_reg_28 (.CK( clk ) , .D( u0_uk_K_r8_28 ) , .Q( u0_uk_K_r9_28 ) , .QN( u0_uk_n205 ) );
  DFF_X1 u0_uk_K_r9_reg_29 (.CK( clk ) , .D( u0_uk_K_r8_29 ) , .Q( u0_uk_K_r9_29 ) , .QN( u0_uk_n204 ) );
  DFF_X1 u0_uk_K_r9_reg_3 (.CK( clk ) , .D( u0_uk_K_r8_3 ) , .Q( u0_uk_K_r9_3 ) , .QN( u0_uk_n225 ) );
  DFF_X1 u0_uk_K_r9_reg_30 (.CK( clk ) , .D( u0_uk_K_r8_30 ) , .Q( u0_uk_K_r9_30 ) );
  DFF_X1 u0_uk_K_r9_reg_31 (.CK( clk ) , .D( u0_uk_K_r8_31 ) , .Q( u0_uk_K_r9_31 ) );
  DFF_X1 u0_uk_K_r9_reg_32 (.CK( clk ) , .D( u0_uk_K_r8_32 ) , .Q( u0_uk_K_r9_32 ) , .QN( u0_uk_n201 ) );
  DFF_X1 u0_uk_K_r9_reg_33 (.CK( clk ) , .D( u0_uk_K_r8_33 ) , .Q( u0_uk_K_r9_33 ) );
  DFF_X1 u0_uk_K_r9_reg_34 (.CK( clk ) , .D( u0_uk_K_r8_34 ) , .Q( u0_uk_K_r9_34 ) , .QN( u0_uk_n200 ) );
  DFF_X1 u0_uk_K_r9_reg_35 (.CK( clk ) , .D( u0_uk_K_r8_35 ) , .Q( u0_uk_K_r9_35 ) );
  DFF_X1 u0_uk_K_r9_reg_36 (.CK( clk ) , .D( u0_uk_K_r8_36 ) , .Q( u0_uk_K_r9_36 ) , .QN( u0_uk_n199 ) );
  DFF_X1 u0_uk_K_r9_reg_37 (.CK( clk ) , .D( u0_uk_K_r8_37 ) , .Q( u0_uk_K_r9_37 ) , .QN( u0_uk_n198 ) );
  DFF_X1 u0_uk_K_r9_reg_38 (.CK( clk ) , .D( u0_uk_K_r8_38 ) , .Q( u0_uk_K_r9_38 ) );
  DFF_X1 u0_uk_K_r9_reg_39 (.CK( clk ) , .D( u0_uk_K_r8_39 ) , .Q( u0_uk_K_r9_39 ) , .QN( u0_uk_n197 ) );
  DFF_X1 u0_uk_K_r9_reg_4 (.CK( clk ) , .D( u0_uk_K_r8_4 ) , .Q( u0_uk_K_r9_4 ) );
  DFF_X1 u0_uk_K_r9_reg_40 (.CK( clk ) , .D( u0_uk_K_r8_40 ) , .Q( u0_uk_K_r9_40 ) , .QN( u0_uk_n196 ) );
  DFF_X1 u0_uk_K_r9_reg_41 (.CK( clk ) , .D( u0_uk_K_r8_41 ) , .Q( u0_uk_K_r9_41 ) , .QN( u0_uk_n195 ) );
  DFF_X1 u0_uk_K_r9_reg_42 (.CK( clk ) , .D( u0_uk_K_r8_42 ) , .Q( u0_uk_K_r9_42 ) , .QN( u0_uk_n194 ) );
  DFF_X1 u0_uk_K_r9_reg_43 (.CK( clk ) , .D( u0_uk_K_r8_43 ) , .Q( u0_uk_K_r9_43 ) , .QN( u0_uk_n193 ) );
  DFF_X1 u0_uk_K_r9_reg_44 (.CK( clk ) , .D( u0_uk_K_r8_44 ) , .Q( u0_uk_K_r9_44 ) , .QN( u0_uk_n192 ) );
  DFF_X1 u0_uk_K_r9_reg_45 (.CK( clk ) , .D( u0_uk_K_r8_45 ) , .Q( u0_uk_K_r9_45 ) );
  DFF_X1 u0_uk_K_r9_reg_46 (.CK( clk ) , .D( u0_uk_K_r8_46 ) , .Q( u0_uk_K_r9_46 ) , .QN( u0_uk_n190 ) );
  DFF_X1 u0_uk_K_r9_reg_47 (.CK( clk ) , .D( u0_uk_K_r8_47 ) , .Q( u0_uk_K_r9_47 ) , .QN( u0_uk_n189 ) );
  DFF_X1 u0_uk_K_r9_reg_48 (.CK( clk ) , .D( u0_uk_K_r8_48 ) , .Q( u0_uk_K_r9_48 ) );
  DFF_X1 u0_uk_K_r9_reg_49 (.CK( clk ) , .D( u0_uk_K_r8_49 ) , .Q( u0_uk_K_r9_49 ) );
  DFF_X1 u0_uk_K_r9_reg_5 (.CK( clk ) , .D( u0_uk_K_r8_5 ) , .Q( u0_uk_K_r9_5 ) );
  DFF_X1 u0_uk_K_r9_reg_50 (.CK( clk ) , .D( u0_uk_K_r8_50 ) , .Q( u0_uk_K_r9_50 ) , .QN( u0_uk_n186 ) );
  DFF_X1 u0_uk_K_r9_reg_51 (.CK( clk ) , .D( u0_uk_K_r8_51 ) , .Q( u0_uk_K_r9_51 ) , .QN( u0_uk_n185 ) );
  DFF_X1 u0_uk_K_r9_reg_52 (.CK( clk ) , .D( u0_uk_K_r8_52 ) , .Q( u0_uk_K_r9_52 ) , .QN( u0_uk_n184 ) );
  DFF_X1 u0_uk_K_r9_reg_53 (.CK( clk ) , .D( u0_uk_K_r8_53 ) , .Q( u0_uk_K_r9_53 ) , .QN( u0_uk_n183 ) );
  DFF_X1 u0_uk_K_r9_reg_54 (.CK( clk ) , .D( u0_uk_K_r8_54 ) , .Q( u0_uk_K_r9_54 ) );
  DFF_X1 u0_uk_K_r9_reg_55 (.CK( clk ) , .D( u0_uk_K_r8_55 ) , .Q( u0_uk_K_r9_55 ) , .QN( u0_uk_n181 ) );
  DFF_X1 u0_uk_K_r9_reg_6 (.CK( clk ) , .D( u0_uk_K_r8_6 ) , .Q( u0_uk_K_r9_6 ) );
  DFF_X1 u0_uk_K_r9_reg_7 (.CK( clk ) , .D( u0_uk_K_r8_7 ) , .Q( u0_uk_K_r9_7 ) );
  DFF_X1 u0_uk_K_r9_reg_8 (.CK( clk ) , .D( u0_uk_K_r8_8 ) , .Q( u0_uk_K_r9_8 ) , .QN( u0_uk_n224 ) );
  DFF_X1 u0_uk_K_r9_reg_9 (.CK( clk ) , .D( u0_uk_K_r8_9 ) , .Q( u0_uk_K_r9_9 ) );
  OAI22_X1 u0_uk_U100 (.ZN( u0_K12_5 ) , .B2( u0_uk_n150 ) , .A2( u0_uk_n176 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U1000 (.B1( decrypt ) , .ZN( u0_K14_46 ) , .B2( u0_uk_n68 ) , .A( u0_uk_n928 ) );
  NAND2_X1 u0_uk_U1001 (.A2( decrypt ) , .A1( u0_uk_K_r12_22 ) , .ZN( u0_uk_n928 ) );
  OAI21_X1 u0_uk_U1002 (.ZN( u0_K8_4 ) , .B2( u0_uk_n351 ) , .A( u0_uk_n743 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U1003 (.A1( u0_uk_K_r6_19 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n743 ) );
  OAI21_X1 u0_uk_U1004 (.B1( decrypt ) , .ZN( u0_K3_5 ) , .B2( u0_uk_n556 ) , .A( u0_uk_n841 ) );
  NAND2_X1 u0_uk_U1005 (.A1( u0_uk_K_r1_10 ) , .A2( u0_uk_n100 ) , .ZN( u0_uk_n841 ) );
  OAI21_X1 u0_uk_U1008 (.B1( decrypt ) , .ZN( u0_K1_13 ) , .B2( u0_uk_n674 ) , .A( u0_uk_n890 ) );
  NAND2_X1 u0_uk_U1009 (.A1( u0_key_r_46 ) , .A2( u0_uk_n60 ) , .ZN( u0_uk_n890 ) );
  OAI21_X1 u0_uk_U1010 (.B1( decrypt ) , .ZN( u0_K1_17 ) , .B2( u0_uk_n705 ) , .A( u0_uk_n888 ) );
  NAND2_X1 u0_uk_U1011 (.A1( u0_key_r_10 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n888 ) );
  OAI21_X1 u0_uk_U1012 (.ZN( u0_K10_21 ) , .A( u0_uk_n1020 ) , .B2( u0_uk_n228 ) , .B1( u0_uk_n31 ) );
  NAND2_X1 u0_uk_U1013 (.A2( decrypt ) , .A1( u0_uk_K_r8_19 ) , .ZN( u0_uk_n1020 ) );
  OAI21_X1 u0_uk_U1016 (.B1( decrypt ) , .ZN( u0_K9_39 ) , .B2( u0_uk_n287 ) , .A( u0_uk_n724 ) );
  NAND2_X1 u0_uk_U1017 (.A2( decrypt ) , .A1( u0_uk_K_r7_31 ) , .ZN( u0_uk_n724 ) );
  OAI21_X1 u0_uk_U1018 (.B1( decrypt ) , .ZN( u0_K4_6 ) , .B2( u0_uk_n523 ) , .A( u0_uk_n820 ) );
  NAND2_X1 u0_uk_U1019 (.A2( decrypt ) , .A1( u0_uk_K_r2_24 ) , .ZN( u0_uk_n820 ) );
  OAI21_X1 u0_uk_U1020 (.ZN( u0_K14_44 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n81 ) , .A( u0_uk_n930 ) );
  NAND2_X1 u0_uk_U1021 (.A1( u0_uk_K_r12_15 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n930 ) );
  OAI21_X1 u0_uk_U1022 (.ZN( u0_K9_44 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n273 ) , .A( u0_uk_n721 ) );
  NAND2_X1 u0_uk_U1023 (.A1( u0_uk_K_r7_0 ) , .A2( u0_uk_n217 ) , .ZN( u0_uk_n721 ) );
  OAI21_X1 u0_uk_U1024 (.ZN( u0_K8_46 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n326 ) , .A( u0_uk_n744 ) );
  NAND2_X1 u0_uk_U1025 (.A1( u0_uk_K_r6_37 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n744 ) );
  OAI21_X1 u0_uk_U1026 (.B1( decrypt ) , .ZN( u0_K10_13 ) , .A( u0_uk_n1023 ) , .B2( u0_uk_n253 ) );
  NAND2_X1 u0_uk_U1027 (.A2( decrypt ) , .A1( u0_uk_K_r8_48 ) , .ZN( u0_uk_n1023 ) );
  OAI21_X1 u0_uk_U1028 (.B1( decrypt ) , .ZN( u0_K12_36 ) , .B2( u0_uk_n160 ) , .A( u0_uk_n970 ) );
  NAND2_X1 u0_uk_U1029 (.A2( decrypt ) , .A1( u0_uk_K_r10_52 ) , .ZN( u0_uk_n970 ) );
  OAI22_X1 u0_uk_U103 (.ZN( u0_K5_5 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n466 ) , .A2( u0_uk_n490 ) );
  NAND2_X1 u0_uk_U1031 (.A2( decrypt ) , .A1( u0_uk_K_r14_42 ) , .ZN( u0_uk_n898 ) );
  NAND2_X1 u0_uk_U1033 (.A2( decrypt ) , .A1( u0_uk_K_r6_30 ) , .ZN( u0_uk_n748 ) );
  OAI21_X1 u0_uk_U1034 (.B1( decrypt ) , .ZN( u0_K6_41 ) , .B2( u0_uk_n413 ) , .A( u0_uk_n790 ) );
  NAND2_X1 u0_uk_U1035 (.A1( u0_uk_K_r4_31 ) , .ZN( u0_uk_n790 ) , .A2( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U1038 (.B1( decrypt ) , .ZN( u0_K8_28 ) , .B2( u0_uk_n326 ) , .A( u0_uk_n756 ) );
  NAND2_X1 u0_uk_U1039 (.A1( u0_uk_K_r6_51 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n756 ) );
  OAI21_X1 u0_uk_U1040 (.ZN( u0_K7_31 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n380 ) , .A( u0_uk_n772 ) );
  NAND2_X1 u0_uk_U1041 (.A1( u0_uk_K_r5_16 ) , .A2( u0_uk_n102 ) , .ZN( u0_uk_n772 ) );
  OAI21_X1 u0_uk_U1042 (.ZN( u0_K14_40 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n65 ) , .A( u0_uk_n931 ) );
  NAND2_X1 u0_uk_U1043 (.A1( u0_uk_K_r12_21 ) , .A2( u0_uk_n110 ) , .ZN( u0_uk_n931 ) );
  OAI21_X1 u0_uk_U1044 (.ZN( u0_K15_14 ) , .B2( u0_uk_n37 ) , .B1( u0_uk_n92 ) , .A( u0_uk_n923 ) );
  NAND2_X1 u0_uk_U1045 (.A1( u0_uk_K_r13_32 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n923 ) );
  OAI21_X1 u0_uk_U1046 (.B1( decrypt ) , .ZN( u0_K10_32 ) , .A( u0_uk_n1013 ) , .B2( u0_uk_n270 ) );
  NAND2_X1 u0_uk_U1047 (.A2( decrypt ) , .A1( u0_uk_K_r8_51 ) , .ZN( u0_uk_n1013 ) );
  OAI21_X1 u0_uk_U1048 (.B1( decrypt ) , .ZN( u0_K5_31 ) , .B2( u0_uk_n487 ) , .A( u0_uk_n812 ) );
  NAND2_X1 u0_uk_U1049 (.A2( decrypt ) , .A1( u0_uk_K_r3_44 ) , .ZN( u0_uk_n812 ) );
  NAND2_X1 u0_uk_U1051 (.A2( decrypt ) , .A1( u0_uk_K_r13_36 ) , .ZN( u0_uk_n918 ) );
  OAI21_X1 u0_uk_U1052 (.ZN( u0_K16_42 ) , .B2( u0_uk_n647 ) , .A( u0_uk_n897 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U1053 (.A2( decrypt ) , .A1( u0_uk_K_r14_38 ) , .ZN( u0_uk_n897 ) );
  OAI21_X1 u0_uk_U1056 (.ZN( u0_K7_38 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n389 ) , .A( u0_uk_n767 ) );
  NAND2_X1 u0_uk_U1057 (.A1( u0_uk_K_r5_8 ) , .A2( u0_uk_n117 ) , .ZN( u0_uk_n767 ) );
  OAI22_X1 u0_uk_U106 (.B1( decrypt ) , .ZN( u0_K2_5 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n611 ) , .B2( u0_uk_n614 ) );
  OAI21_X1 u0_uk_U1060 (.B1( decrypt ) , .ZN( u0_K14_24 ) , .B2( u0_uk_n76 ) , .A( u0_uk_n937 ) );
  NAND2_X1 u0_uk_U1061 (.A2( decrypt ) , .A1( u0_uk_K_r12_41 ) , .ZN( u0_uk_n937 ) );
  INV_X1 u0_uk_U1063 (.A( u0_key_r_7 ) , .ZN( u0_uk_n711 ) );
  INV_X1 u0_uk_U1066 (.A( u0_key_r_33 ) , .ZN( u0_uk_n691 ) );
  INV_X1 u0_uk_U1068 (.A( u0_key_r_26 ) , .ZN( u0_uk_n697 ) );
  INV_X1 u0_uk_U1070 (.A( u0_key_r_34 ) , .ZN( u0_uk_n690 ) );
  INV_X1 u0_uk_U1071 (.A( u0_key_r_27 ) , .ZN( u0_uk_n696 ) );
  INV_X1 u0_uk_U1072 (.A( u0_key_r_24 ) , .ZN( u0_uk_n699 ) );
  INV_X1 u0_uk_U1074 (.A( u0_key_r_37 ) , .ZN( u0_uk_n687 ) );
  INV_X1 u0_uk_U1075 (.A( u0_key_r_52 ) , .ZN( u0_uk_n675 ) );
  INV_X1 u0_uk_U1079 (.A( u0_key_r_1 ) , .ZN( u0_uk_n715 ) );
  OAI22_X1 u0_uk_U108 (.B1( decrypt ) , .ZN( u0_K10_41 ) , .A1( u0_uk_n163 ) , .B2( u0_uk_n236 ) , .A2( u0_uk_n264 ) );
  INV_X1 u0_uk_U1083 (.A( u0_key_r_17 ) , .ZN( u0_uk_n705 ) );
  INV_X1 u0_uk_U1084 (.A( u0_key_r_53 ) , .ZN( u0_uk_n674 ) );
  OAI21_X1 u0_uk_U1085 (.ZN( u0_K13_28 ) , .B2( u0_uk_n105 ) , .B1( u0_uk_n252 ) , .A( u0_uk_n947 ) );
  NAND2_X1 u0_uk_U1086 (.A1( u0_uk_K_r11_21 ) , .A2( u0_uk_n214 ) , .ZN( u0_uk_n947 ) );
  OAI22_X1 u0_uk_U109 (.ZN( u0_K14_41 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n77 ) , .A2( u0_uk_n82 ) , .B1( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U1097 (.ZN( u0_K5_39 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n482 ) , .A( u0_uk_n808 ) );
  NAND2_X1 u0_uk_U1098 (.A1( u0_uk_K_r3_16 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n808 ) );
  INV_X1 u0_uk_U1099 (.A( u0_key_r_40 ) , .ZN( u0_uk_n684 ) );
  AOI22_X1 u0_uk_U1102 (.B2( u0_uk_K_r0_34 ) , .A2( u0_uk_K_r0_55 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n868 ) );
  AOI22_X1 u0_uk_U1104 (.B2( u0_key_r_32 ) , .A2( u0_key_r_39 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n892 ) );
  AOI22_X1 u0_uk_U1110 (.B2( u0_uk_K_r9_12 ) , .A2( u0_uk_K_r9_18 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n982 ) );
  AOI22_X1 u0_uk_U1114 (.B2( u0_uk_K_r6_3 ) , .A2( u0_uk_K_r6_53 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n761 ) );
  AOI22_X1 u0_uk_U1118 (.B1( decrypt ) , .B2( u0_uk_K_r10_27 ) , .A2( u0_uk_K_r10_4 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n963 ) );
  AOI22_X1 u0_uk_U1120 (.B1( decrypt ) , .B2( u0_uk_K_r0_13 ) , .A2( u0_uk_K_r0_34 ) , .A1( u0_uk_n222 ) , .ZN( u0_uk_n855 ) );
  AOI22_X1 u0_uk_U1122 (.B2( u0_uk_K_r3_24 ) , .A2( u0_uk_K_r3_47 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n816 ) );
  AOI22_X1 u0_uk_U1124 (.B2( u0_uk_K_r5_26 ) , .A2( u0_uk_K_r5_48 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n188 ) , .ZN( u0_uk_n783 ) );
  INV_X1 u0_uk_U1127 (.ZN( u0_K7_32 ) , .A( u0_uk_n771 ) );
  AOI22_X1 u0_uk_U1128 (.B2( u0_uk_K_r5_0 ) , .A2( u0_uk_K_r5_51 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n771 ) );
  AOI22_X1 u0_uk_U1130 (.B2( u0_uk_K_r7_23 ) , .A2( u0_uk_K_r7_30 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n148 ) , .ZN( u0_uk_n723 ) );
  AOI22_X1 u0_uk_U1134 (.B2( u0_uk_K_r7_15 ) , .A2( u0_uk_K_r7_22 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n722 ) );
  INV_X1 u0_uk_U1139 (.ZN( u0_K7_34 ) , .A( u0_uk_n770 ) );
  OAI22_X1 u0_uk_U114 (.ZN( u0_K12_47 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n152 ) , .B2( u0_uk_n179 ) );
  AOI22_X1 u0_uk_U1140 (.A1( decrypt ) , .B2( u0_uk_K_r5_0 ) , .A2( u0_uk_K_r5_35 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n770 ) );
  AOI22_X1 u0_uk_U1142 (.A1( decrypt ) , .B2( u0_uk_K_r8_17 ) , .A2( u0_uk_K_r8_39 ) , .ZN( u0_uk_n1024 ) , .B1( u0_uk_n203 ) );
  INV_X1 u0_uk_U1143 (.ZN( u0_K13_12 ) , .A( u0_uk_n958 ) );
  AOI22_X1 u0_uk_U1144 (.B2( u0_uk_K_r11_34 ) , .A2( u0_uk_K_r11_54 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n958 ) );
  AOI22_X1 u0_uk_U1146 (.A1( decrypt ) , .B2( u0_uk_K_r6_10 ) , .A2( u0_uk_K_r6_17 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n759 ) );
  AOI22_X1 u0_uk_U1148 (.A1( decrypt ) , .B2( u0_uk_K_r3_29 ) , .A2( u0_uk_K_r3_38 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n810 ) );
  AOI22_X1 u0_uk_U1149 (.B2( u0_uk_K_r3_15 ) , .A2( u0_uk_K_r3_38 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n230 ) , .ZN( u0_uk_n806 ) );
  INV_X1 u0_uk_U1150 (.ZN( u0_K5_43 ) , .A( u0_uk_n806 ) );
  AOI22_X1 u0_uk_U1153 (.B2( u0_uk_K_r7_24 ) , .A2( u0_uk_K_r7_6 ) , .B1( u0_uk_n10 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n734 ) );
  AOI22_X1 u0_uk_U1155 (.A1( decrypt ) , .B2( u0_uk_K_r4_17 ) , .A2( u0_uk_K_r4_55 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n793 ) );
  INV_X1 u0_uk_U1158 (.ZN( u0_K8_3 ) , .A( u0_uk_n749 ) );
  AOI22_X1 u0_uk_U116 (.B2( u0_uk_K_r9_15 ) , .A2( u0_uk_K_r9_23 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n985 ) );
  AOI22_X1 u0_uk_U1160 (.B2( u0_uk_K_r10_39 ) , .A2( u0_uk_K_r10_48 ) , .B1( u0_uk_n11 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n978 ) );
  INV_X1 u0_uk_U1161 (.ZN( u0_K12_1 ) , .A( u0_uk_n978 ) );
  AOI22_X1 u0_uk_U1162 (.B2( u0_uk_K_r7_20 ) , .A2( u0_uk_K_r7_27 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n729 ) );
  OAI22_X1 u0_uk_U118 (.ZN( u0_K8_47 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n327 ) );
  OAI22_X1 u0_uk_U119 (.ZN( u0_K7_47 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n388 ) , .A2( u0_uk_n402 ) );
  OAI22_X1 u0_uk_U122 (.B1( decrypt ) , .ZN( u0_K5_47 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n469 ) , .B2( u0_uk_n493 ) );
  OAI21_X1 u0_uk_U124 (.B1( decrypt ) , .ZN( u0_K2_47 ) , .B2( u0_uk_n617 ) , .A( u0_uk_n856 ) );
  NAND2_X1 u0_uk_U125 (.A1( u0_uk_K_r0_52 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n856 ) );
  OAI22_X1 u0_uk_U126 (.A1( decrypt ) , .ZN( u0_K1_15 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n691 ) , .B2( u0_uk_n697 ) );
  OAI21_X1 u0_uk_U128 (.B1( decrypt ) , .ZN( u0_K5_15 ) , .B2( u0_uk_n479 ) , .A( u0_uk_n817 ) );
  NAND2_X1 u0_uk_U129 (.A2( decrypt ) , .A1( u0_uk_K_r3_34 ) , .ZN( u0_uk_n817 ) );
  AOI22_X1 u0_uk_U131 (.B2( u0_uk_K_r11_11 ) , .A2( u0_uk_K_r11_48 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n956 ) );
  OAI22_X1 u0_uk_U132 (.ZN( u0_K7_15 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n364 ) , .A2( u0_uk_n404 ) );
  INV_X1 u0_uk_U133 (.ZN( u0_K12_15 ) , .A( u0_uk_n980 ) );
  AOI22_X1 u0_uk_U134 (.B2( u0_uk_K_r10_25 ) , .A2( u0_uk_K_r10_34 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n980 ) );
  OAI22_X1 u0_uk_U135 (.B1( decrypt ) , .ZN( u0_K3_15 ) , .A1( u0_uk_n191 ) , .B2( u0_uk_n541 ) , .A2( u0_uk_n576 ) );
  OAI22_X1 u0_uk_U138 (.A1( decrypt ) , .ZN( u0_K12_19 ) , .B2( u0_uk_n138 ) , .A2( u0_uk_n176 ) , .B1( u0_uk_n217 ) );
  OAI21_X1 u0_uk_U140 (.B1( decrypt ) , .ZN( u0_K6_19 ) , .B2( u0_uk_n444 ) , .A( u0_uk_n798 ) );
  NAND2_X1 u0_uk_U141 (.A1( u0_uk_K_r4_48 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n798 ) );
  OAI21_X1 u0_uk_U142 (.ZN( u0_K2_15 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n597 ) , .A( u0_uk_n865 ) );
  NAND2_X1 u0_uk_U143 (.A1( u0_uk_K_r0_19 ) , .A2( u0_uk_n102 ) , .ZN( u0_uk_n865 ) );
  OAI22_X1 u0_uk_U146 (.ZN( u0_K10_15 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n229 ) , .A2( u0_uk_n266 ) , .A1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U147 (.ZN( u0_K15_15 ) , .B2( u0_uk_n15 ) , .B1( u0_uk_n163 ) , .A( u0_uk_n922 ) );
  NAND2_X1 u0_uk_U148 (.A1( u0_uk_K_r13_19 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n922 ) );
  INV_X1 u0_uk_U149 (.ZN( u0_K14_19 ) , .A( u0_uk_n938 ) );
  AOI22_X1 u0_uk_U150 (.B2( u0_uk_K_r12_25 ) , .A2( u0_uk_K_r12_33 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n207 ) , .ZN( u0_uk_n938 ) );
  AOI22_X1 u0_uk_U152 (.B2( u0_uk_K_r9_10 ) , .A2( u0_uk_K_r9_48 ) , .ZN( u0_uk_n1000 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n220 ) );
  AOI22_X1 u0_uk_U154 (.B2( decrypt ) , .B1( u0_uk_K_r7_13 ) , .A2( u0_uk_K_r7_20 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n735 ) );
  OAI21_X1 u0_uk_U157 (.B1( decrypt ) , .ZN( u0_K3_19 ) , .B2( u0_uk_n564 ) , .A( u0_uk_n852 ) );
  NAND2_X1 u0_uk_U158 (.A2( decrypt ) , .A1( u0_uk_K_r1_33 ) , .ZN( u0_uk_n852 ) );
  INV_X1 u0_uk_U159 (.ZN( u0_K2_19 ) , .A( u0_uk_n864 ) );
  AOI22_X1 u0_uk_U160 (.B2( u0_uk_K_r0_11 ) , .A2( u0_uk_K_r0_47 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n864 ) );
  OAI22_X1 u0_uk_U161 (.A1( decrypt ) , .ZN( u0_K14_15 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n47 ) , .A2( u0_uk_n85 ) );
  OAI22_X1 u0_uk_U162 (.B1( decrypt ) , .ZN( u0_K8_19 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n343 ) , .B2( u0_uk_n350 ) );
  OAI22_X1 u0_uk_U163 (.A1( decrypt ) , .ZN( u0_K10_19 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n245 ) , .B2( u0_uk_n255 ) );
  OAI22_X1 u0_uk_U164 (.ZN( u0_K5_30 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n463 ) , .B2( u0_uk_n480 ) );
  OAI22_X1 u0_uk_U165 (.B1( decrypt ) , .ZN( u0_K2_30 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n599 ) , .B2( u0_uk_n628 ) );
  OAI22_X1 u0_uk_U166 (.ZN( u0_K14_30 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n250 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n77 ) );
  OAI21_X1 u0_uk_U170 (.B1( decrypt ) , .ZN( u0_K1_14 ) , .B2( u0_uk_n698 ) , .A( u0_uk_n889 ) );
  NAND2_X1 u0_uk_U171 (.A1( u0_key_r_18 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n889 ) );
  INV_X1 u0_uk_U172 (.A( u0_key_r_25 ) , .ZN( u0_uk_n698 ) );
  OAI21_X1 u0_uk_U173 (.ZN( u0_K8_30 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n333 ) , .A( u0_uk_n753 ) );
  NAND2_X1 u0_uk_U174 (.A1( u0_uk_K_r6_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n753 ) );
  OAI22_X1 u0_uk_U177 (.ZN( u0_K13_14 ) , .A2( u0_uk_n108 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n132 ) , .B1( u0_uk_n242 ) );
  OAI22_X1 u0_uk_U178 (.ZN( u0_K12_14 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n165 ) , .B2( u0_uk_n170 ) , .B1( u0_uk_n202 ) );
  AOI22_X1 u0_uk_U181 (.A1( decrypt ) , .B2( u0_uk_K_r9_12 ) , .A2( u0_uk_K_r9_6 ) , .ZN( u0_uk_n1002 ) , .B1( u0_uk_n163 ) );
  OAI21_X1 u0_uk_U184 (.B1( decrypt ) , .ZN( u0_K9_14 ) , .B2( u0_uk_n284 ) , .A( u0_uk_n738 ) );
  NAND2_X1 u0_uk_U185 (.A2( decrypt ) , .A1( u0_uk_K_r7_34 ) , .ZN( u0_uk_n738 ) );
  AOI22_X1 u0_uk_U188 (.B2( u0_uk_K_r0_11 ) , .A2( u0_uk_K_r0_32 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n866 ) );
  OAI22_X1 u0_uk_U192 (.A1( decrypt ) , .ZN( u0_K10_14 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n227 ) , .B2( u0_uk_n258 ) );
  OAI21_X1 u0_uk_U193 (.B1( decrypt ) , .ZN( u0_K13_30 ) , .B2( u0_uk_n112 ) , .A( u0_uk_n945 ) );
  NAND2_X1 u0_uk_U194 (.A1( u0_uk_K_r11_28 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n945 ) );
  INV_X1 u0_uk_U195 (.ZN( u0_K7_24 ) , .A( u0_uk_n776 ) );
  AOI22_X1 u0_uk_U196 (.B2( u0_uk_K_r5_18 ) , .A2( u0_uk_K_r5_40 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n776 ) );
  OAI22_X1 u0_uk_U197 (.A1( decrypt ) , .ZN( u0_K4_24 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n495 ) , .B2( u0_uk_n536 ) );
  INV_X1 u0_uk_U198 (.ZN( u0_K3_24 ) , .A( u0_uk_n851 ) );
  AOI22_X1 u0_uk_U199 (.B2( u0_uk_K_r1_17 ) , .A2( u0_uk_K_r1_41 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n851 ) );
  OAI22_X1 u0_uk_U200 (.ZN( u0_K15_24 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n24 ) , .A2( u0_uk_n42 ) );
  OAI21_X1 u0_uk_U201 (.B1( decrypt ) , .ZN( u0_K1_30 ) , .B2( u0_uk_n675 ) , .A( u0_uk_n880 ) );
  NAND2_X1 u0_uk_U202 (.A1( u0_key_r_45 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n880 ) );
  OAI21_X1 u0_uk_U203 (.ZN( u0_K9_30 ) , .B2( u0_uk_n288 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n728 ) );
  NAND2_X1 u0_uk_U204 (.A2( decrypt ) , .A1( u0_uk_K_r7_29 ) , .ZN( u0_uk_n728 ) );
  OAI22_X1 u0_uk_U209 (.B1( decrypt ) , .ZN( u0_K3_14 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n541 ) , .B2( u0_uk_n548 ) );
  INV_X1 u0_uk_U210 (.ZN( u0_K4_31 ) , .A( u0_uk_n826 ) );
  AOI22_X1 u0_uk_U211 (.B1( decrypt ) , .B2( u0_uk_K_r2_31 ) , .A2( u0_uk_K_r2_49 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n826 ) );
  OAI22_X1 u0_uk_U212 (.B1( decrypt ) , .ZN( u0_K1_31 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n707 ) , .A2( u0_uk_n711 ) );
  INV_X1 u0_uk_U213 (.A( u0_key_r_14 ) , .ZN( u0_uk_n707 ) );
  OAI22_X1 u0_uk_U215 (.ZN( u0_K8_31 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n321 ) , .B2( u0_uk_n359 ) );
  OAI22_X1 u0_uk_U220 (.ZN( u0_K2_31 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n613 ) , .B2( u0_uk_n628 ) );
  INV_X1 u0_uk_U223 (.ZN( u0_K10_39 ) , .A( u0_uk_n1007 ) );
  AOI22_X1 u0_uk_U224 (.B2( u0_uk_K_r8_44 ) , .A2( u0_uk_K_r8_52 ) , .ZN( u0_uk_n1007 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n217 ) );
  NAND2_X1 u0_uk_U232 (.A2( decrypt ) , .A1( u0_key_r_15 ) , .ZN( u0_uk_n875 ) );
  OAI22_X1 u0_uk_U237 (.ZN( u0_K14_39 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n56 ) );
  OAI22_X1 u0_uk_U238 (.A1( decrypt ) , .ZN( u0_K13_39 ) , .A2( u0_uk_n114 ) , .B2( u0_uk_n133 ) , .B1( u0_uk_n250 ) );
  OAI21_X1 u0_uk_U239 (.B1( decrypt ) , .ZN( u0_K12_39 ) , .B2( u0_uk_n168 ) , .A( u0_uk_n969 ) );
  NAND2_X1 u0_uk_U240 (.A1( u0_uk_K_r10_16 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n969 ) );
  OAI21_X1 u0_uk_U242 (.ZN( u0_K16_44 ) , .B1( u0_uk_n110 ) , .B2( u0_uk_n642 ) , .A( u0_uk_n895 ) );
  NAND2_X1 u0_uk_U243 (.A1( u0_uk_K_r14_43 ) , .ZN( u0_uk_n895 ) , .A2( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U245 (.ZN( u0_K15_48 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n34 ) , .A( u0_uk_n914 ) );
  NAND2_X1 u0_uk_U246 (.A1( u0_uk_K_r13_35 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n914 ) );
  OAI22_X1 u0_uk_U249 (.ZN( u0_K8_48 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n223 ) , .B2( u0_uk_n347 ) , .A2( u0_uk_n354 ) );
  INV_X1 u0_uk_U252 (.ZN( u0_K1_44 ) , .A( u0_uk_n872 ) );
  AOI22_X1 u0_uk_U253 (.B2( u0_key_r_36 ) , .A2( u0_key_r_43 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n872 ) );
  OAI22_X1 u0_uk_U254 (.ZN( u0_K14_48 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n52 ) , .B2( u0_uk_n90 ) );
  OAI22_X1 u0_uk_U255 (.ZN( u0_K13_44 ) , .B1( u0_uk_n110 ) , .A2( u0_uk_n119 ) , .B2( u0_uk_n134 ) , .A1( u0_uk_n191 ) );
  OAI21_X1 u0_uk_U256 (.B1( decrypt ) , .ZN( u0_K13_48 ) , .B2( u0_uk_n103 ) , .A( u0_uk_n942 ) );
  NAND2_X1 u0_uk_U257 (.A1( u0_uk_K_r11_8 ) , .A2( u0_uk_n141 ) , .ZN( u0_uk_n942 ) );
  OAI22_X1 u0_uk_U260 (.A1( decrypt ) , .ZN( u0_K12_48 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n158 ) , .B2( u0_uk_n167 ) );
  AOI22_X1 u0_uk_U265 (.A1( decrypt ) , .B2( u0_uk_K_r7_16 ) , .A2( u0_uk_K_r7_9 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n719 ) );
  OAI22_X1 u0_uk_U266 (.ZN( u0_K7_44 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n378 ) , .B2( u0_uk_n399 ) );
  OAI22_X1 u0_uk_U267 (.ZN( u0_K7_48 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n257 ) , .A2( u0_uk_n367 ) , .B2( u0_uk_n387 ) );
  OAI22_X1 u0_uk_U270 (.B1( decrypt ) , .ZN( u0_K5_44 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n463 ) , .B2( u0_uk_n469 ) );
  OAI22_X1 u0_uk_U271 (.B1( decrypt ) , .ZN( u0_K5_48 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n474 ) , .B2( u0_uk_n481 ) );
  OAI22_X1 u0_uk_U272 (.ZN( u0_K4_44 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .A2( u0_uk_n521 ) , .B2( u0_uk_n538 ) );
  OAI22_X1 u0_uk_U276 (.A1( decrypt ) , .ZN( u0_K2_44 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n585 ) , .B2( u0_uk_n607 ) );
  NAND2_X1 u0_uk_U281 (.A2( decrypt ) , .A1( u0_uk_K_r4_18 ) , .ZN( u0_uk_n786 ) );
  OAI22_X1 u0_uk_U282 (.A1( decrypt ) , .ZN( u0_K2_6 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n588 ) , .B2( u0_uk_n609 ) );
  INV_X1 u0_uk_U284 (.ZN( u0_K15_8 ) , .A( u0_uk_n913 ) );
  AOI22_X1 u0_uk_U285 (.B2( u0_uk_K_r13_13 ) , .A2( u0_uk_K_r13_17 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n230 ) , .ZN( u0_uk_n913 ) );
  OAI22_X1 u0_uk_U286 (.ZN( u0_K12_8 ) , .A2( u0_uk_n136 ) , .B2( u0_uk_n157 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n83 ) );
  AOI22_X1 u0_uk_U289 (.A1( decrypt ) , .B2( u0_uk_K_r5_26 ) , .A2( u0_uk_K_r5_4 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n763 ) );
  OAI22_X1 u0_uk_U290 (.ZN( u0_K5_8 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n451 ) , .B2( u0_uk_n473 ) );
  OAI21_X1 u0_uk_U294 (.B1( decrypt ) , .ZN( u0_K2_8 ) , .B2( u0_uk_n618 ) , .A( u0_uk_n854 ) );
  NAND2_X1 u0_uk_U295 (.A2( decrypt ) , .A1( u0_uk_K_r0_17 ) , .ZN( u0_uk_n854 ) );
  OAI22_X1 u0_uk_U296 (.ZN( u0_K7_26 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n368 ) , .B2( u0_uk_n388 ) );
  AOI22_X1 u0_uk_U298 (.B2( u0_key_r_31 ) , .A2( u0_key_r_51 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n883 ) );
  OAI22_X1 u0_uk_U299 (.B1( decrypt ) , .ZN( u0_K16_8 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n654 ) , .A2( u0_uk_n667 ) );
  AOI22_X1 u0_uk_U301 (.A1( decrypt ) , .B2( u0_uk_K_r7_15 ) , .A2( u0_uk_K_r7_8 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n731 ) );
  INV_X1 u0_uk_U302 (.ZN( u0_K4_26 ) , .A( u0_uk_n831 ) );
  AOI22_X1 u0_uk_U303 (.B2( u0_uk_K_r2_16 ) , .A2( u0_uk_K_r2_7 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n831 ) );
  OAI21_X1 u0_uk_U310 (.ZN( u0_K13_26 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n123 ) , .A( u0_uk_n948 ) );
  NAND2_X1 u0_uk_U311 (.A2( decrypt ) , .A1( u0_uk_K_r11_7 ) , .ZN( u0_uk_n948 ) );
  OAI22_X1 u0_uk_U312 (.B1( decrypt ) , .ZN( u0_K5_26 ) , .A1( u0_uk_n242 ) , .B2( u0_uk_n482 ) , .A2( u0_uk_n492 ) );
  OAI22_X1 u0_uk_U313 (.ZN( u0_K2_26 ) , .A1( u0_uk_n164 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n593 ) , .B2( u0_uk_n599 ) );
  OAI22_X1 u0_uk_U314 (.A1( decrypt ) , .ZN( u0_K16_26 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n633 ) , .B2( u0_uk_n647 ) );
  OAI22_X1 u0_uk_U315 (.ZN( u0_K14_26 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n49 ) , .B2( u0_uk_n66 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U319 (.ZN( u0_K3_26 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n242 ) , .A2( u0_uk_n543 ) , .B2( u0_uk_n559 ) );
  OAI22_X1 u0_uk_U321 (.B1( decrypt ) , .ZN( u0_K13_46 ) , .A2( u0_uk_n113 ) , .B2( u0_uk_n125 ) , .A1( u0_uk_n230 ) );
  OAI22_X1 u0_uk_U322 (.ZN( u0_K12_46 ) , .A2( u0_uk_n140 ) , .B2( u0_uk_n180 ) , .A1( u0_uk_n252 ) , .B1( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U323 (.ZN( u0_K9_46 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n281 ) , .A( u0_uk_n720 ) );
  NAND2_X1 u0_uk_U324 (.A2( decrypt ) , .A1( u0_uk_K_r7_37 ) , .ZN( u0_uk_n720 ) );
  OAI22_X1 u0_uk_U325 (.ZN( u0_K5_46 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n457 ) , .B2( u0_uk_n494 ) );
  OAI22_X1 u0_uk_U326 (.ZN( u0_K4_46 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n514 ) , .B2( u0_uk_n528 ) );
  OAI21_X1 u0_uk_U327 (.ZN( u0_K3_46 ) , .B1( u0_uk_n209 ) , .B2( u0_uk_n561 ) , .A( u0_uk_n842 ) );
  NAND2_X1 u0_uk_U328 (.A1( u0_uk_K_r1_22 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n842 ) );
  OAI22_X1 u0_uk_U329 (.A1( decrypt ) , .ZN( u0_K2_46 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n595 ) , .A2( u0_uk_n622 ) );
  OAI21_X1 u0_uk_U330 (.B1( decrypt ) , .ZN( u0_K1_46 ) , .B2( u0_uk_n715 ) , .A( u0_uk_n871 ) );
  NAND2_X1 u0_uk_U331 (.A1( u0_key_r_49 ) , .A2( u0_uk_n117 ) , .ZN( u0_uk_n871 ) );
  INV_X1 u0_uk_U333 (.ZN( u0_K7_46 ) , .A( u0_uk_n765 ) );
  AOI22_X1 u0_uk_U334 (.A1( decrypt ) , .B2( u0_uk_K_r5_23 ) , .A2( u0_uk_K_r5_31 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n765 ) );
  OAI21_X1 u0_uk_U335 (.B1( decrypt ) , .ZN( u0_K16_4 ) , .B2( u0_uk_n631 ) , .A( u0_uk_n894 ) );
  NAND2_X1 u0_uk_U336 (.A1( u0_uk_K_r14_3 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n894 ) );
  OAI22_X1 u0_uk_U337 (.ZN( u0_K15_4 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n38 ) , .A2( u0_uk_n8 ) );
  OAI22_X1 u0_uk_U338 (.A1( decrypt ) , .ZN( u0_K14_4 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n64 ) , .B2( u0_uk_n72 ) );
  OAI22_X1 u0_uk_U339 (.ZN( u0_K10_4 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n227 ) , .B2( u0_uk_n246 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U343 (.B1( decrypt ) , .ZN( u0_K5_4 ) , .B2( u0_uk_n477 ) , .A( u0_uk_n804 ) );
  NAND2_X1 u0_uk_U344 (.A1( u0_uk_K_r3_4 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n804 ) );
  OAI22_X1 u0_uk_U348 (.B1( decrypt ) , .ZN( u0_K2_4 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n591 ) , .B2( u0_uk_n620 ) );
  NAND2_X1 u0_uk_U350 (.A1( u0_key_r_3 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n869 ) );
  AOI22_X1 u0_uk_U356 (.A2( u0_uk_K_r8_2 ) , .B2( u0_uk_K_r8_22 ) , .ZN( u0_uk_n1006 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n217 ) );
  OAI21_X1 u0_uk_U358 (.B1( decrypt ) , .ZN( u0_K12_40 ) , .B2( u0_uk_n159 ) , .A( u0_uk_n967 ) );
  NAND2_X1 u0_uk_U359 (.A2( decrypt ) , .A1( u0_uk_K_r10_49 ) , .ZN( u0_uk_n967 ) );
  OAI22_X1 u0_uk_U361 (.A1( decrypt ) , .ZN( u0_K13_40 ) , .A2( u0_uk_n104 ) , .B2( u0_uk_n114 ) , .B1( u0_uk_n147 ) );
  OAI22_X1 u0_uk_U363 (.ZN( u0_K8_40 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n327 ) , .B2( u0_uk_n333 ) );
  OAI22_X1 u0_uk_U364 (.ZN( u0_K7_40 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n394 ) , .A2( u0_uk_n406 ) );
  OAI22_X1 u0_uk_U365 (.ZN( u0_K4_40 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n506 ) , .B2( u0_uk_n516 ) );
  OAI22_X1 u0_uk_U366 (.ZN( u0_K2_40 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n592 ) , .A2( u0_uk_n623 ) );
  NAND2_X1 u0_uk_U368 (.A2( decrypt ) , .A1( u0_uk_K_r13_31 ) , .ZN( u0_uk_n917 ) );
  OAI21_X1 u0_uk_U369 (.ZN( u0_K2_33 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n600 ) , .A( u0_uk_n859 ) );
  NAND2_X1 u0_uk_U370 (.A1( u0_uk_K_r0_31 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n859 ) );
  OAI22_X1 u0_uk_U371 (.ZN( u0_K1_28 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n710 ) , .B2( u0_uk_n715 ) );
  INV_X1 u0_uk_U372 (.A( u0_key_r_8 ) , .ZN( u0_uk_n710 ) );
  OAI21_X1 u0_uk_U376 (.B1( decrypt ) , .ZN( u0_K4_28 ) , .B2( u0_uk_n507 ) , .A( u0_uk_n830 ) );
  NAND2_X1 u0_uk_U377 (.A2( decrypt ) , .A1( u0_uk_K_r2_21 ) , .ZN( u0_uk_n830 ) );
  OAI22_X1 u0_uk_U384 (.ZN( u0_K9_28 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n274 ) , .B2( u0_uk_n281 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U385 (.ZN( u0_K7_28 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n378 ) , .B2( u0_uk_n387 ) );
  OAI22_X1 u0_uk_U386 (.B1( decrypt ) , .ZN( u0_K5_28 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n488 ) , .B2( u0_uk_n492 ) );
  OAI22_X1 u0_uk_U387 (.ZN( u0_K14_1 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n75 ) , .B2( u0_uk_n80 ) );
  OAI21_X1 u0_uk_U393 (.ZN( u0_K10_16 ) , .A( u0_uk_n1022 ) , .B2( u0_uk_n228 ) , .B1( u0_uk_n250 ) );
  NAND2_X1 u0_uk_U394 (.A1( u0_uk_K_r8_32 ) , .ZN( u0_uk_n1022 ) , .A2( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U395 (.ZN( u0_K9_16 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n303 ) , .B2( u0_uk_n310 ) );
  OAI22_X1 u0_uk_U397 (.B1( decrypt ) , .ZN( u0_K6_16 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n416 ) , .B2( u0_uk_n422 ) );
  OAI21_X1 u0_uk_U398 (.ZN( u0_K3_16 ) , .B1( u0_uk_n102 ) , .B2( u0_uk_n540 ) , .A( u0_uk_n853 ) );
  NAND2_X1 u0_uk_U399 (.A2( decrypt ) , .A1( u0_uk_K_r1_6 ) , .ZN( u0_uk_n853 ) );
  OAI22_X1 u0_uk_U400 (.A1( decrypt ) , .ZN( u0_K1_16 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n690 ) , .B2( u0_uk_n696 ) );
  OAI21_X1 u0_uk_U402 (.ZN( u0_K15_9 ) , .B2( u0_uk_n15 ) , .A( u0_uk_n912 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U403 (.A1( u0_uk_K_r13_4 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n912 ) );
  OAI21_X1 u0_uk_U404 (.B1( decrypt ) , .ZN( u0_K14_9 ) , .B2( u0_uk_n70 ) , .A( u0_uk_n926 ) );
  NAND2_X1 u0_uk_U405 (.A1( u0_uk_K_r12_18 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n926 ) );
  OAI22_X1 u0_uk_U407 (.A1( decrypt ) , .ZN( u0_K12_9 ) , .A2( u0_uk_n136 ) , .B2( u0_uk_n143 ) , .B1( u0_uk_n148 ) );
  OAI22_X1 u0_uk_U409 (.ZN( u0_K8_9 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n162 ) , .B2( u0_uk_n350 ) , .A2( u0_uk_n356 ) );
  INV_X1 u0_uk_U412 (.ZN( u0_K10_37 ) , .A( u0_uk_n1009 ) );
  AOI22_X1 u0_uk_U413 (.A1( decrypt ) , .B2( u0_uk_K_r8_28 ) , .A2( u0_uk_K_r8_52 ) , .ZN( u0_uk_n1009 ) , .B1( u0_uk_n207 ) );
  AOI22_X1 u0_uk_U415 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_7 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n751 ) );
  AOI22_X1 u0_uk_U417 (.B2( u0_uk_K_r8_17 ) , .A2( u0_uk_K_r8_27 ) , .ZN( u0_uk_n1005 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) );
  INV_X1 u0_uk_U418 (.ZN( u0_K9_9 ) , .A( u0_uk_n718 ) );
  AOI22_X1 u0_uk_U419 (.B2( u0_uk_K_r7_13 ) , .A1( u0_uk_K_r7_6 ) , .A2( u0_uk_n128 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n718 ) );
  OAI22_X1 u0_uk_U420 (.ZN( u0_K7_9 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n390 ) , .B2( u0_uk_n397 ) );
  OAI21_X1 u0_uk_U422 (.ZN( u0_K3_9 ) , .B1( u0_uk_n209 ) , .B2( u0_uk_n563 ) , .A( u0_uk_n840 ) );
  NAND2_X1 u0_uk_U423 (.A1( u0_uk_K_r1_18 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n840 ) );
  OAI22_X1 u0_uk_U424 (.ZN( u0_K2_9 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n597 ) , .A2( u0_uk_n626 ) );
  OAI22_X1 u0_uk_U425 (.ZN( u0_K15_1 ) , .A2( u0_uk_n1 ) , .B2( u0_uk_n20 ) , .A1( u0_uk_n230 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U426 (.ZN( u0_K1_33 ) , .A( u0_uk_n878 ) );
  AOI22_X1 u0_uk_U427 (.B1( decrypt ) , .B2( u0_key_r_44 ) , .A2( u0_key_r_51 ) , .A1( u0_uk_n222 ) , .ZN( u0_uk_n878 ) );
  OAI22_X1 u0_uk_U428 (.B1( decrypt ) , .ZN( u0_K5_1 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n459 ) , .B2( u0_uk_n466 ) );
  OAI22_X1 u0_uk_U429 (.ZN( u0_K16_9 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n630 ) , .B2( u0_uk_n637 ) );
  OAI22_X1 u0_uk_U431 (.ZN( u0_K2_16 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n596 ) , .B2( u0_uk_n614 ) , .A1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U432 (.ZN( u0_K7_16 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n362 ) , .A( u0_uk_n782 ) );
  NAND2_X1 u0_uk_U433 (.A1( u0_uk_K_r5_32 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n782 ) );
  OAI22_X1 u0_uk_U434 (.ZN( u0_K15_16 ) , .A2( u0_uk_n14 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n29 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U435 (.B1( decrypt ) , .ZN( u0_K5_16 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n478 ) , .A2( u0_uk_n491 ) );
  AOI22_X1 u0_uk_U438 (.B2( u0_uk_K_r7_1 ) , .A2( u0_uk_K_r7_8 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n727 ) );
  AOI22_X1 u0_uk_U440 (.A1( decrypt ) , .B2( u0_uk_K_r8_22 ) , .A2( u0_uk_K_r8_42 ) , .ZN( u0_uk_n1012 ) , .B1( u0_uk_n207 ) );
  OAI21_X1 u0_uk_U441 (.ZN( u0_K12_33 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n140 ) , .A( u0_uk_n971 ) );
  NAND2_X1 u0_uk_U442 (.A1( u0_uk_K_r10_14 ) , .A2( u0_uk_n118 ) , .ZN( u0_uk_n971 ) );
  OAI22_X1 u0_uk_U443 (.ZN( u0_K16_33 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n633 ) , .B2( u0_uk_n638 ) );
  OAI22_X1 u0_uk_U445 (.ZN( u0_K13_33 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n130 ) , .B2( u0_uk_n135 ) , .B1( u0_uk_n238 ) );
  OAI22_X1 u0_uk_U446 (.B1( decrypt ) , .ZN( u0_K8_33 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n355 ) , .B2( u0_uk_n360 ) );
  OAI22_X1 u0_uk_U447 (.ZN( u0_K7_33 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n374 ) , .B2( u0_uk_n394 ) );
  OAI22_X1 u0_uk_U455 (.ZN( u0_K13_37 ) , .A2( u0_uk_n112 ) , .B2( u0_uk_n124 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U457 (.B1( decrypt ) , .ZN( u0_K11_37 ) , .B2( u0_uk_n194 ) , .A( u0_uk_n989 ) );
  NAND2_X1 u0_uk_U458 (.A1( u0_uk_K_r9_38 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n989 ) );
  NAND2_X1 u0_uk_U460 (.A2( decrypt ) , .A1( u0_uk_K_r7_7 ) , .ZN( u0_uk_n725 ) );
  OAI22_X1 u0_uk_U463 (.ZN( u0_K4_37 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n251 ) , .A2( u0_uk_n513 ) , .B2( u0_uk_n527 ) );
  INV_X1 u0_uk_U464 (.ZN( u0_K6_9 ) , .A( u0_uk_n785 ) );
  AOI22_X1 u0_uk_U465 (.A1( decrypt ) , .B2( u0_uk_K_r4_3 ) , .A2( u0_uk_K_r4_41 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n785 ) );
  OAI22_X1 u0_uk_U466 (.B1( decrypt ) , .ZN( u0_K5_9 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n451 ) , .B2( u0_uk_n461 ) );
  OAI22_X1 u0_uk_U467 (.ZN( u0_K5_37 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n455 ) , .B2( u0_uk_n493 ) );
  OAI21_X1 u0_uk_U470 (.B1( decrypt ) , .ZN( u0_K10_36 ) , .A( u0_uk_n1010 ) , .B2( u0_uk_n269 ) );
  NAND2_X1 u0_uk_U471 (.A1( u0_uk_K_r8_21 ) , .ZN( u0_uk_n1010 ) , .A2( u0_uk_n11 ) );
  OAI21_X1 u0_uk_U472 (.ZN( u0_K14_29 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n51 ) , .A( u0_uk_n935 ) );
  NAND2_X1 u0_uk_U473 (.A1( u0_uk_K_r12_44 ) , .A2( u0_uk_n145 ) , .ZN( u0_uk_n935 ) );
  OAI22_X1 u0_uk_U481 (.ZN( u0_K2_29 ) , .A1( u0_uk_n188 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n606 ) , .A2( u0_uk_n621 ) );
  OAI22_X1 u0_uk_U486 (.ZN( u0_K7_29 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n368 ) , .B2( u0_uk_n399 ) );
  OAI22_X1 u0_uk_U487 (.ZN( u0_K5_29 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n462 ) , .B2( u0_uk_n481 ) );
  OAI22_X1 u0_uk_U488 (.ZN( u0_K14_2 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n57 ) , .B2( u0_uk_n64 ) );
  OAI21_X1 u0_uk_U493 (.ZN( u0_K8_2 ) , .B2( u0_uk_n343 ) , .A( u0_uk_n754 ) , .B1( u0_uk_n83 ) );
  NAND2_X1 u0_uk_U494 (.A1( u0_uk_K_r6_27 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n754 ) );
  OAI21_X1 u0_uk_U497 (.ZN( u0_K9_12 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n315 ) , .A( u0_uk_n740 ) );
  NAND2_X1 u0_uk_U498 (.A2( decrypt ) , .A1( u0_uk_K_r7_53 ) , .ZN( u0_uk_n740 ) );
  OAI22_X1 u0_uk_U503 (.ZN( u0_K10_17 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n234 ) , .B2( u0_uk_n262 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U506 (.ZN( u0_K8_29 ) , .A( u0_uk_n755 ) );
  AOI22_X1 u0_uk_U507 (.A1( decrypt ) , .B2( u0_uk_K_r6_28 ) , .A2( u0_uk_K_r6_35 ) , .B1( u0_uk_n208 ) , .ZN( u0_uk_n755 ) );
  AOI22_X1 u0_uk_U509 (.A1( decrypt ) , .B2( u0_uk_K_r9_4 ) , .A2( u0_uk_K_r9_55 ) , .ZN( u0_uk_n1001 ) , .B1( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U515 (.B1( decrypt ) , .ZN( u0_K3_17 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n548 ) , .B2( u0_uk_n571 ) );
  INV_X1 u0_uk_U516 (.ZN( u0_K4_29 ) , .A( u0_uk_n829 ) );
  AOI22_X1 u0_uk_U517 (.B2( u0_uk_K_r2_31 ) , .A2( u0_uk_K_r2_36 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n829 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U518 (.ZN( u0_K15_12 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n25 ) , .A2( u0_uk_n43 ) );
  OAI22_X1 u0_uk_U519 (.A1( decrypt ) , .ZN( u0_K14_12 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n53 ) , .B2( u0_uk_n57 ) );
  OAI21_X1 u0_uk_U520 (.ZN( u0_K12_12 ) , .B1( u0_uk_n109 ) , .B2( u0_uk_n169 ) , .A( u0_uk_n981 ) );
  NAND2_X1 u0_uk_U521 (.A2( decrypt ) , .A1( u0_uk_K_r10_11 ) , .ZN( u0_uk_n981 ) );
  OAI21_X1 u0_uk_U524 (.ZN( u0_K5_12 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n483 ) , .A( u0_uk_n818 ) );
  NAND2_X1 u0_uk_U525 (.A1( u0_uk_K_r3_11 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n818 ) );
  OAI22_X1 u0_uk_U527 (.B1( decrypt ) , .ZN( u0_K3_12 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n547 ) , .B2( u0_uk_n552 ) );
  OAI22_X1 u0_uk_U528 (.B1( decrypt ) , .ZN( u0_K2_12 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n610 ) , .A2( u0_uk_n625 ) );
  OAI22_X1 u0_uk_U529 (.ZN( u0_K15_2 ) , .A2( u0_uk_n1 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n30 ) );
  OAI22_X1 u0_uk_U530 (.ZN( u0_K5_2 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n486 ) , .A2( u0_uk_n491 ) );
  OAI22_X1 u0_uk_U537 (.ZN( u0_K15_17 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n220 ) , .B2( u0_uk_n26 ) , .A2( u0_uk_n44 ) );
  OAI22_X1 u0_uk_U538 (.ZN( u0_K14_17 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n54 ) , .B2( u0_uk_n78 ) );
  OAI22_X1 u0_uk_U539 (.ZN( u0_K5_17 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n464 ) , .B2( u0_uk_n484 ) , .A1( u0_uk_n99 ) );
  AOI22_X1 u0_uk_U543 (.B2( u0_uk_K_r4_4 ) , .A2( u0_uk_K_r4_55 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n800 ) );
  OAI22_X1 u0_uk_U545 (.ZN( u0_K14_36 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n88 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U546 (.A1( decrypt ) , .ZN( u0_K13_36 ) , .A2( u0_uk_n105 ) , .B2( u0_uk_n111 ) , .B1( u0_uk_n147 ) );
  OAI22_X1 u0_uk_U548 (.ZN( u0_K2_36 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n250 ) , .A2( u0_uk_n600 ) , .B2( u0_uk_n616 ) );
  AOI22_X1 u0_uk_U551 (.B2( u0_uk_K_r3_29 ) , .A2( u0_uk_K_r3_52 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n809 ) );
  AOI22_X1 u0_uk_U553 (.A1( decrypt ) , .B2( u0_uk_K_r14_16 ) , .A2( u0_uk_K_r14_23 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n904 ) );
  OAI22_X1 u0_uk_U554 (.ZN( u0_K16_36 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n63 ) , .A2( u0_uk_n648 ) , .B2( u0_uk_n655 ) );
  AOI22_X1 u0_uk_U559 (.B2( u0_uk_K_r5_1 ) , .A2( u0_uk_K_r5_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n768 ) );
  AOI22_X1 u0_uk_U561 (.A1( decrypt ) , .B2( u0_uk_K_r9_15 ) , .A2( u0_uk_K_r9_7 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n990 ) );
  AOI22_X1 u0_uk_U563 (.A1( decrypt ) , .B2( u0_uk_K_r13_23 ) , .A2( u0_uk_K_r13_44 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n916 ) );
  INV_X1 u0_uk_U564 (.ZN( u0_K10_38 ) , .A( u0_uk_n1008 ) );
  AOI22_X1 u0_uk_U565 (.B2( u0_uk_K_r8_28 ) , .A2( u0_uk_K_r8_8 ) , .ZN( u0_uk_n1008 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U566 (.B1( decrypt ) , .ZN( u0_K8_36 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n328 ) , .B2( u0_uk_n334 ) );
  OAI22_X1 u0_uk_U568 (.B1( decrypt ) , .ZN( u0_K5_38 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n470 ) , .B2( u0_uk_n494 ) );
  OAI22_X1 u0_uk_U569 (.A1( decrypt ) , .ZN( u0_K10_10 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n235 ) , .B2( u0_uk_n263 ) );
  INV_X1 u0_uk_U57 (.A( decrypt ) , .ZN( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U570 (.ZN( u0_K5_10 ) , .B1( u0_uk_n208 ) , .A2( u0_uk_n465 ) , .B2( u0_uk_n485 ) , .A1( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U572 (.ZN( u0_K15_10 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n19 ) , .A( u0_uk_n925 ) );
  NAND2_X1 u0_uk_U573 (.A1( u0_uk_K_r13_55 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n925 ) );
  OAI22_X1 u0_uk_U574 (.A1( decrypt ) , .ZN( u0_K14_10 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n74 ) , .B2( u0_uk_n79 ) );
  NAND2_X1 u0_uk_U576 (.A2( decrypt ) , .A1( u0_uk_K_r9_54 ) , .ZN( u0_uk_n1004 ) );
  INV_X1 u0_uk_U577 (.ZN( u0_K13_10 ) , .A( u0_uk_n960 ) );
  AOI22_X1 u0_uk_U578 (.B1( decrypt ) , .B2( u0_uk_K_r11_26 ) , .A2( u0_uk_K_r11_6 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n960 ) );
  INV_X1 u0_uk_U579 (.ZN( u0_K9_10 ) , .A( u0_uk_n742 ) );
  AOI22_X1 u0_uk_U580 (.B2( u0_uk_K_r7_25 ) , .A2( u0_uk_K_r7_32 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n742 ) );
  INV_X1 u0_uk_U582 (.ZN( u0_K6_10 ) , .A( u0_uk_n801 ) );
  AOI22_X1 u0_uk_U583 (.B2( u0_uk_K_r4_3 ) , .A2( u0_uk_K_r4_54 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n801 ) );
  AOI22_X1 u0_uk_U585 (.A1( decrypt ) , .B2( u0_uk_K_r2_26 ) , .A2( u0_uk_K_r2_6 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n839 ) );
  OAI22_X1 u0_uk_U589 (.B1( decrypt ) , .ZN( u0_K16_22 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n646 ) , .B2( u0_uk_n653 ) );
  AOI22_X1 u0_uk_U591 (.B2( u0_uk_K_r11_10 ) , .A2( u0_uk_K_r11_47 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n949 ) );
  INV_X1 u0_uk_U592 (.ZN( u0_K11_22 ) , .A( u0_uk_n997 ) );
  AOI22_X1 u0_uk_U593 (.B2( u0_uk_K_r9_13 ) , .A2( u0_uk_K_r9_19 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n997 ) );
  INV_X1 u0_uk_U594 (.ZN( u0_K10_22 ) , .A( u0_uk_n1019 ) );
  AOI22_X1 u0_uk_U595 (.B1( decrypt ) , .B2( u0_uk_K_r8_27 ) , .A2( u0_uk_K_r8_5 ) , .ZN( u0_uk_n1019 ) , .A1( u0_uk_n162 ) );
  INV_X1 u0_uk_U596 (.ZN( u0_K9_22 ) , .A( u0_uk_n732 ) );
  AOI22_X1 u0_uk_U597 (.B1( decrypt ) , .B2( u0_uk_K_r7_41 ) , .A2( u0_uk_K_r7_48 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n732 ) );
  OAI22_X1 u0_uk_U598 (.ZN( u0_K8_22 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n323 ) , .B2( u0_uk_n329 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U60 (.ZN( u0_K11_34 ) , .A( u0_uk_n991 ) );
  AOI22_X1 u0_uk_U600 (.A1( decrypt ) , .B2( u0_uk_K_r3_24 ) , .A2( u0_uk_K_r3_33 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n815 ) );
  INV_X1 u0_uk_U601 (.ZN( u0_K1_22 ) , .A( u0_uk_n885 ) );
  AOI22_X1 u0_uk_U602 (.B2( u0_key_r_25 ) , .A2( u0_key_r_32 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n885 ) );
  OAI21_X1 u0_uk_U606 (.ZN( u0_K7_35 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n406 ) , .A( u0_uk_n769 ) );
  NAND2_X1 u0_uk_U607 (.A1( u0_uk_K_r5_37 ) , .ZN( u0_uk_n769 ) , .A2( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U608 (.A1( decrypt ) , .ZN( u0_K2_35 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n595 ) , .B2( u0_uk_n613 ) );
  OAI22_X1 u0_uk_U609 (.ZN( u0_K13_35 ) , .B2( u0_uk_n124 ) , .B1( u0_uk_n214 ) , .A1( u0_uk_n27 ) , .A2( u0_uk_n95 ) );
  AOI22_X1 u0_uk_U61 (.B2( u0_uk_K_r9_45 ) , .A2( u0_uk_K_r9_49 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n991 ) );
  OAI22_X1 u0_uk_U610 (.A1( decrypt ) , .ZN( u0_K12_35 ) , .A2( u0_uk_n151 ) , .B2( u0_uk_n160 ) , .B1( u0_uk_n238 ) );
  AOI22_X1 u0_uk_U613 (.B2( u0_uk_K_r12_1 ) , .A2( u0_uk_K_r12_7 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n933 ) );
  INV_X1 u0_uk_U614 (.ZN( u0_K10_35 ) , .A( u0_uk_n1011 ) );
  AOI22_X1 u0_uk_U615 (.B2( u0_uk_K_r8_2 ) , .A2( u0_uk_K_r8_37 ) , .ZN( u0_uk_n1011 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n222 ) );
  AOI22_X1 u0_uk_U617 (.B1( decrypt ) , .B2( u0_uk_K_r7_16 ) , .A2( u0_uk_K_r7_23 ) , .A1( u0_uk_n191 ) , .ZN( u0_uk_n726 ) );
  OAI22_X1 u0_uk_U619 (.B1( decrypt ) , .ZN( u0_K4_35 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n498 ) , .B2( u0_uk_n527 ) );
  INV_X1 u0_uk_U62 (.ZN( u0_K8_34 ) , .A( u0_uk_n752 ) );
  OAI21_X1 u0_uk_U622 (.ZN( u0_K16_11 ) , .B1( u0_uk_n146 ) , .B2( u0_uk_n646 ) , .A( u0_uk_n911 ) );
  NAND2_X1 u0_uk_U623 (.A1( u0_uk_K_r14_39 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n911 ) );
  OAI22_X1 u0_uk_U626 (.ZN( u0_K14_11 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n80 ) , .B1( u0_uk_n83 ) , .A2( u0_uk_n87 ) );
  INV_X1 u0_uk_U628 (.ZN( u0_K13_11 ) , .A( u0_uk_n959 ) );
  AOI22_X1 u0_uk_U629 (.B2( u0_uk_K_r11_17 ) , .A2( u0_uk_K_r11_54 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n959 ) );
  AOI22_X1 u0_uk_U63 (.B2( u0_uk_K_r6_14 ) , .A2( u0_uk_K_r6_21 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n752 ) );
  OAI22_X1 u0_uk_U630 (.ZN( u0_K10_11 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n245 ) , .B2( u0_uk_n262 ) , .B1( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U631 (.B1( decrypt ) , .ZN( u0_K8_11 ) , .B2( u0_uk_n323 ) , .A( u0_uk_n762 ) );
  NAND2_X1 u0_uk_U632 (.A1( u0_uk_K_r6_55 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n762 ) );
  OAI21_X1 u0_uk_U635 (.B1( decrypt ) , .ZN( u0_K2_11 ) , .B2( u0_uk_n591 ) , .A( u0_uk_n867 ) );
  NAND2_X1 u0_uk_U636 (.A1( u0_uk_K_r0_25 ) , .A2( u0_uk_n109 ) , .ZN( u0_uk_n867 ) );
  AOI22_X1 u0_uk_U638 (.B2( u0_uk_K_r7_48 ) , .A2( u0_uk_K_r7_55 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n741 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U639 (.B1( decrypt ) , .ZN( u0_K6_11 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n431 ) , .B2( u0_uk_n435 ) );
  OAI22_X1 u0_uk_U640 (.ZN( u0_K5_11 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n465 ) , .A2( u0_uk_n489 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U647 (.ZN( u0_K16_45 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n638 ) , .B2( u0_uk_n641 ) );
  OAI22_X1 u0_uk_U648 (.A1( decrypt ) , .ZN( u0_K1_45 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n680 ) , .B2( u0_uk_n687 ) );
  INV_X1 u0_uk_U649 (.A( u0_key_r_44 ) , .ZN( u0_uk_n680 ) );
  OAI22_X1 u0_uk_U650 (.ZN( u0_K14_43 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n56 ) , .B2( u0_uk_n59 ) , .A1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U651 (.ZN( u0_K7_43 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n374 ) , .A2( u0_uk_n403 ) );
  OAI21_X1 u0_uk_U653 (.ZN( u0_K2_43 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n612 ) , .A( u0_uk_n857 ) );
  NAND2_X1 u0_uk_U654 (.A1( u0_uk_K_r0_2 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n857 ) );
  OAI22_X1 u0_uk_U657 (.ZN( u0_K9_25 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n273 ) , .B2( u0_uk_n280 ) , .A1( u0_uk_n99 ) );
  AOI22_X1 u0_uk_U66 (.B2( u0_uk_K_r12_30 ) , .A2( u0_uk_K_r12_36 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n934 ) );
  AOI22_X1 u0_uk_U661 (.A2( u0_uk_K_r13_2 ) , .B2( u0_uk_K_r13_23 ) , .A1( u0_uk_n163 ) , .ZN( u0_uk_n915 ) , .B1( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U666 (.ZN( u0_K12_45 ) , .B2( u0_uk_n174 ) , .B1( u0_uk_n191 ) , .A( u0_uk_n964 ) );
  NAND2_X1 u0_uk_U667 (.A1( u0_uk_K_r10_43 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n964 ) );
  OAI22_X1 u0_uk_U668 (.ZN( u0_K11_43 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n184 ) , .B2( u0_uk_n226 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U669 (.ZN( u0_K10_43 ) , .A1( u0_uk_n214 ) , .B2( u0_uk_n237 ) , .A2( u0_uk_n265 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U67 (.A1( decrypt ) , .ZN( u0_K12_34 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n158 ) , .A2( u0_uk_n173 ) );
  OAI22_X1 u0_uk_U672 (.B1( decrypt ) , .ZN( u0_K9_45 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n276 ) , .B2( u0_uk_n317 ) );
  OAI21_X1 u0_uk_U673 (.ZN( u0_K5_45 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n488 ) , .A( u0_uk_n805 ) );
  NAND2_X1 u0_uk_U674 (.A2( decrypt ) , .A1( u0_uk_K_r3_43 ) , .ZN( u0_uk_n805 ) );
  OAI21_X1 u0_uk_U675 (.B1( decrypt ) , .ZN( u0_K4_43 ) , .B2( u0_uk_n499 ) , .A( u0_uk_n823 ) );
  NAND2_X1 u0_uk_U676 (.A1( u0_uk_K_r2_29 ) , .A2( u0_uk_n100 ) , .ZN( u0_uk_n823 ) );
  OAI22_X1 u0_uk_U678 (.ZN( u0_K10_7 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n234 ) , .B2( u0_uk_n254 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U679 (.ZN( u0_K15_7 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n19 ) , .B2( u0_uk_n35 ) );
  OAI21_X1 u0_uk_U68 (.ZN( u0_K6_34 ) , .B1( u0_uk_n118 ) , .B2( u0_uk_n417 ) , .A( u0_uk_n792 ) );
  OAI21_X1 u0_uk_U680 (.B1( decrypt ) , .ZN( u0_K12_7 ) , .B2( u0_uk_n138 ) , .A( u0_uk_n961 ) );
  NAND2_X1 u0_uk_U681 (.A1( u0_uk_K_r10_19 ) , .A2( u0_uk_n27 ) , .ZN( u0_uk_n961 ) );
  OAI21_X1 u0_uk_U686 (.ZN( u0_K15_25 ) , .B2( u0_uk_n12 ) , .B1( u0_uk_n147 ) , .A( u0_uk_n921 ) );
  NAND2_X1 u0_uk_U687 (.A1( u0_uk_K_r13_22 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n921 ) );
  NAND2_X1 u0_uk_U69 (.A1( u0_uk_K_r4_49 ) , .ZN( u0_uk_n792 ) , .A2( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U690 (.ZN( u0_K5_25 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n475 ) , .A( u0_uk_n814 ) );
  NAND2_X1 u0_uk_U691 (.A1( u0_uk_K_r3_35 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n814 ) );
  OAI21_X1 u0_uk_U692 (.B1( decrypt ) , .ZN( u0_K2_25 ) , .B2( u0_uk_n594 ) , .A( u0_uk_n863 ) );
  NAND2_X1 u0_uk_U693 (.A1( u0_uk_K_r0_22 ) , .ZN( u0_uk_n863 ) , .A2( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U695 (.ZN( u0_K12_25 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n154 ) , .B2( u0_uk_n159 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U696 (.A1( decrypt ) , .ZN( u0_K10_25 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n247 ) , .A2( u0_uk_n265 ) );
  AOI22_X1 u0_uk_U698 (.A1( decrypt ) , .B2( u0_uk_K_r6_21 ) , .A2( u0_uk_K_r6_28 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n746 ) );
  OAI22_X1 u0_uk_U70 (.ZN( u0_K4_34 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n208 ) , .A2( u0_uk_n506 ) , .B2( u0_uk_n522 ) );
  OAI22_X1 u0_uk_U701 (.ZN( u0_K8_25 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n320 ) , .B2( u0_uk_n325 ) , .B1( u0_uk_n60 ) );
  INV_X1 u0_uk_U704 (.ZN( u0_K13_7 ) , .A( u0_uk_n939 ) );
  AOI22_X1 u0_uk_U705 (.A1( decrypt ) , .B2( u0_uk_K_r11_10 ) , .A2( u0_uk_K_r11_5 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n939 ) );
  OAI21_X1 u0_uk_U706 (.ZN( u0_K5_7 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n453 ) , .A( u0_uk_n802 ) );
  NAND2_X1 u0_uk_U707 (.A1( u0_uk_K_r3_19 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n802 ) );
  INV_X1 u0_uk_U708 (.ZN( u0_K7_25 ) , .A( u0_uk_n775 ) );
  AOI22_X1 u0_uk_U709 (.A1( decrypt ) , .B2( u0_uk_K_r5_31 ) , .A2( u0_uk_K_r5_7 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n775 ) );
  OAI21_X1 u0_uk_U71 (.B1( decrypt ) , .ZN( u0_K3_34 ) , .B2( u0_uk_n559 ) , .A( u0_uk_n848 ) );
  INV_X1 u0_uk_U710 (.ZN( u0_K1_25 ) , .A( u0_uk_n884 ) );
  AOI22_X1 u0_uk_U711 (.B2( u0_key_r_29 ) , .A2( u0_key_r_36 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n884 ) );
  AOI22_X1 u0_uk_U713 (.A1( decrypt ) , .B2( u0_uk_K_r2_16 ) , .A2( u0_uk_K_r2_49 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n832 ) );
  OAI22_X1 u0_uk_U718 (.ZN( u0_K8_32 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n325 ) , .B2( u0_uk_n332 ) );
  NAND2_X1 u0_uk_U72 (.A1( u0_uk_K_r1_36 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n848 ) );
  OAI22_X1 u0_uk_U720 (.ZN( u0_K13_32 ) , .B2( u0_uk_n106 ) , .A2( u0_uk_n130 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U723 (.B1( decrypt ) , .ZN( u0_K5_32 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n476 ) , .B2( u0_uk_n480 ) );
  OAI22_X1 u0_uk_U724 (.ZN( u0_K14_32 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n51 ) , .B2( u0_uk_n89 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U725 (.A1( decrypt ) , .ZN( u0_K9_32 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n280 ) , .B2( u0_uk_n287 ) );
  OAI22_X1 u0_uk_U727 (.A1( decrypt ) , .ZN( u0_K14_42 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n59 ) , .B2( u0_uk_n90 ) );
  OAI22_X1 u0_uk_U728 (.A1( decrypt ) , .ZN( u0_K13_42 ) , .A2( u0_uk_n119 ) , .B2( u0_uk_n125 ) , .B1( u0_uk_n147 ) );
  OAI22_X1 u0_uk_U729 (.ZN( u0_K11_42 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n186 ) , .B2( u0_uk_n194 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U73 (.B1( decrypt ) , .ZN( u0_K2_34 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n585 ) , .B2( u0_uk_n616 ) );
  OAI21_X1 u0_uk_U731 (.ZN( u0_K5_42 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n476 ) , .A( u0_uk_n807 ) );
  NAND2_X1 u0_uk_U732 (.A1( u0_uk_K_r3_9 ) , .ZN( u0_uk_n807 ) , .A2( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U733 (.ZN( u0_K4_42 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n521 ) , .B2( u0_uk_n528 ) );
  OAI22_X1 u0_uk_U735 (.ZN( u0_K2_42 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n584 ) , .B2( u0_uk_n592 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U736 (.ZN( u0_K7_42 ) , .A( u0_uk_n766 ) );
  AOI22_X1 u0_uk_U737 (.A1( decrypt ) , .B2( u0_uk_K_r5_1 ) , .A2( u0_uk_K_r5_36 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n766 ) );
  INV_X1 u0_uk_U742 (.ZN( u0_K1_42 ) , .A( u0_uk_n873 ) );
  AOI22_X1 u0_uk_U743 (.B2( u0_key_r_31 ) , .A2( u0_key_r_38 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n873 ) );
  OAI21_X1 u0_uk_U744 (.B1( decrypt ) , .ZN( u0_K14_27 ) , .B2( u0_uk_n49 ) , .A( u0_uk_n936 ) );
  NAND2_X1 u0_uk_U745 (.A1( u0_uk_K_r12_42 ) , .A2( u0_uk_n129 ) , .ZN( u0_uk_n936 ) );
  OAI21_X1 u0_uk_U747 (.B1( decrypt ) , .ZN( u0_K10_27 ) , .A( u0_uk_n1016 ) , .B2( u0_uk_n256 ) );
  NAND2_X1 u0_uk_U748 (.A1( u0_uk_K_r8_43 ) , .ZN( u0_uk_n1016 ) , .A2( u0_uk_n11 ) );
  OAI22_X1 u0_uk_U749 (.ZN( u0_K8_27 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n354 ) , .B2( u0_uk_n359 ) );
  OAI22_X1 u0_uk_U751 (.ZN( u0_K12_13 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n137 ) , .B2( u0_uk_n169 ) , .B1( u0_uk_n238 ) );
  OAI22_X1 u0_uk_U753 (.ZN( u0_K8_13 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n257 ) , .B2( u0_uk_n351 ) , .A2( u0_uk_n357 ) );
  OAI22_X1 u0_uk_U754 (.B1( decrypt ) , .ZN( u0_K6_13 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n422 ) , .B2( u0_uk_n426 ) );
  OAI22_X1 u0_uk_U756 (.ZN( u0_K1_21 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n699 ) , .B2( u0_uk_n705 ) );
  OAI21_X1 u0_uk_U757 (.ZN( u0_K9_13 ) , .B2( u0_uk_n309 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n739 ) );
  NAND2_X1 u0_uk_U758 (.A2( decrypt ) , .A1( u0_uk_K_r7_5 ) , .ZN( u0_uk_n739 ) );
  OAI22_X1 u0_uk_U760 (.ZN( u0_K13_27 ) , .A2( u0_uk_n111 ) , .B2( u0_uk_n134 ) , .B1( u0_uk_n238 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U761 (.A1( decrypt ) , .ZN( u0_K14_21 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n48 ) , .B2( u0_uk_n74 ) );
  OAI21_X1 u0_uk_U762 (.B1( decrypt ) , .ZN( u0_K11_21 ) , .B2( u0_uk_n221 ) , .A( u0_uk_n998 ) );
  NAND2_X1 u0_uk_U763 (.A1( u0_uk_K_r9_5 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n998 ) );
  OAI22_X1 u0_uk_U765 (.ZN( u0_K5_21 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n459 ) , .B2( u0_uk_n479 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U767 (.ZN( u0_K2_21 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n620 ) , .A2( u0_uk_n624 ) );
  OAI22_X1 u0_uk_U768 (.ZN( u0_K15_21 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n38 ) , .A2( u0_uk_n42 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U769 (.A1( decrypt ) , .ZN( u0_K14_13 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n71 ) , .B2( u0_uk_n76 ) );
  OAI21_X1 u0_uk_U77 (.ZN( u0_K10_23 ) , .A( u0_uk_n1018 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n268 ) );
  OAI22_X1 u0_uk_U770 (.B1( decrypt ) , .ZN( u0_K4_27 ) , .A1( u0_uk_n202 ) , .A2( u0_uk_n512 ) , .B2( u0_uk_n538 ) );
  OAI22_X1 u0_uk_U773 (.B1( decrypt ) , .ZN( u0_K6_27 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n424 ) , .B2( u0_uk_n429 ) );
  AOI22_X1 u0_uk_U775 (.A1( decrypt ) , .B2( u0_uk_K_r3_15 ) , .A2( u0_uk_K_r3_51 ) , .B1( u0_uk_n217 ) , .ZN( u0_uk_n813 ) );
  OAI21_X1 u0_uk_U778 (.ZN( u0_K3_27 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n543 ) , .A( u0_uk_n850 ) );
  NAND2_X1 u0_uk_U779 (.A1( u0_uk_K_r1_42 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n850 ) );
  NAND2_X1 u0_uk_U78 (.A1( u0_uk_K_r8_13 ) , .ZN( u0_uk_n1018 ) , .A2( u0_uk_n252 ) );
  INV_X1 u0_uk_U780 (.ZN( u0_K13_13 ) , .A( u0_uk_n957 ) );
  AOI22_X1 u0_uk_U781 (.B2( u0_uk_K_r11_11 ) , .A2( u0_uk_K_r11_6 ) , .B1( u0_uk_n207 ) , .A1( u0_uk_n94 ) , .ZN( u0_uk_n957 ) );
  AOI22_X1 u0_uk_U783 (.B1( decrypt ) , .B2( u0_uk_K_r11_34 ) , .A2( u0_uk_K_r11_39 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n950 ) );
  AOI22_X1 u0_uk_U785 (.B2( u0_uk_K_r10_25 ) , .A2( u0_uk_K_r10_48 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n976 ) );
  INV_X1 u0_uk_U786 (.ZN( u0_K6_21 ) , .A( u0_uk_n797 ) );
  AOI22_X1 u0_uk_U787 (.B2( u0_uk_K_r4_11 ) , .A2( u0_uk_K_r4_5 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n797 ) );
  OAI21_X1 u0_uk_U788 (.ZN( u0_K16_13 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n631 ) , .A( u0_uk_n909 ) );
  NAND2_X1 u0_uk_U789 (.A1( u0_uk_K_r14_46 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n909 ) );
  OAI22_X1 u0_uk_U79 (.ZN( u0_K8_23 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n340 ) , .B2( u0_uk_n345 ) , .B1( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U790 (.ZN( u0_K7_21 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n362 ) , .A( u0_uk_n779 ) );
  NAND2_X1 u0_uk_U791 (.A1( u0_uk_K_r5_19 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n779 ) );
  INV_X1 u0_uk_U792 (.ZN( u0_K7_27 ) , .A( u0_uk_n774 ) );
  AOI22_X1 u0_uk_U793 (.B2( u0_uk_K_r5_23 ) , .A2( u0_uk_K_r5_43 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n774 ) );
  INV_X1 u0_uk_U796 (.ZN( u0_K9_27 ) , .A( u0_uk_n730 ) );
  AOI22_X1 u0_uk_U797 (.B2( u0_uk_K_r7_2 ) , .A2( u0_uk_K_r7_9 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n730 ) , .B1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U80 (.B1( decrypt ) , .ZN( u0_K6_23 ) , .B2( u0_uk_n416 ) , .A( u0_uk_n796 ) );
  OAI22_X1 u0_uk_U806 (.B1( decrypt ) , .ZN( u0_K5_18 ) , .A1( u0_uk_n251 ) , .B2( u0_uk_n452 ) , .A2( u0_uk_n489 ) );
  NAND2_X1 u0_uk_U81 (.A2( decrypt ) , .A1( u0_uk_K_r4_27 ) , .ZN( u0_uk_n796 ) );
  OAI21_X1 u0_uk_U810 (.ZN( u0_K12_20 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n166 ) , .A( u0_uk_n977 ) );
  NAND2_X1 u0_uk_U811 (.A1( u0_uk_K_r10_47 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n977 ) );
  OAI22_X1 u0_uk_U814 (.ZN( u0_K2_18 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n588 ) , .B2( u0_uk_n619 ) , .B1( u0_uk_n63 ) );
  OAI21_X1 u0_uk_U815 (.B1( decrypt ) , .ZN( u0_K16_18 ) , .B2( u0_uk_n629 ) , .A( u0_uk_n906 ) );
  NAND2_X1 u0_uk_U816 (.A1( u0_uk_K_r14_5 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n906 ) );
  OAI22_X1 u0_uk_U817 (.A1( decrypt ) , .ZN( u0_K10_18 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n254 ) , .A2( u0_uk_n268 ) );
  OAI22_X1 u0_uk_U818 (.A1( decrypt ) , .ZN( u0_K15_18 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n36 ) , .A2( u0_uk_n6 ) );
  OAI22_X1 u0_uk_U82 (.A1( decrypt ) , .ZN( u0_K3_23 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n572 ) , .A2( u0_uk_n577 ) );
  OAI22_X1 u0_uk_U823 (.ZN( u0_K15_20 ) , .B2( u0_uk_n14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n43 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U825 (.ZN( u0_K9_18 ) , .A( u0_uk_n736 ) );
  AOI22_X1 u0_uk_U826 (.B1( decrypt ) , .B2( u0_uk_K_r7_39 ) , .A2( u0_uk_K_r7_46 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n736 ) );
  AOI22_X1 u0_uk_U828 (.A1( decrypt ) , .B2( u0_uk_K_r4_11 ) , .A2( u0_uk_K_r4_17 ) , .B1( u0_uk_n208 ) , .ZN( u0_uk_n799 ) );
  OAI22_X1 u0_uk_U83 (.ZN( u0_K2_23 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n589 ) , .B2( u0_uk_n610 ) );
  AOI22_X1 u0_uk_U830 (.A1( decrypt ) , .B2( u0_uk_K_r9_10 ) , .A2( u0_uk_K_r9_4 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n999 ) );
  INV_X1 u0_uk_U831 (.ZN( u0_K9_20 ) , .A( u0_uk_n733 ) );
  AOI22_X1 u0_uk_U832 (.B2( u0_uk_K_r7_32 ) , .A2( u0_uk_K_r7_39 ) , .B1( u0_uk_n10 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n733 ) );
  AOI22_X1 u0_uk_U834 (.A1( decrypt ) , .B2( u0_uk_K_r5_18 ) , .A2( u0_uk_K_r5_53 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n780 ) );
  OAI22_X1 u0_uk_U837 (.A1( decrypt ) , .ZN( u0_K12_22 ) , .A2( u0_uk_n156 ) , .B2( u0_uk_n166 ) , .B1( u0_uk_n222 ) );
  OAI21_X1 u0_uk_U838 (.ZN( u0_K4_22 ) , .B2( u0_uk_n531 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n834 ) );
  NAND2_X1 u0_uk_U839 (.A2( decrypt ) , .A1( u0_uk_K_r2_47 ) , .ZN( u0_uk_n834 ) );
  OAI21_X1 u0_uk_U84 (.ZN( u0_K11_41 ) , .B2( u0_uk_n186 ) , .B1( u0_uk_n203 ) , .A( u0_uk_n987 ) );
  OAI22_X1 u0_uk_U842 (.ZN( u0_K15_6 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n24 ) , .A2( u0_uk_n6 ) );
  AOI22_X1 u0_uk_U846 (.B2( u0_uk_K_r6_10 ) , .A2( u0_uk_K_r6_3 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n749 ) );
  NAND2_X1 u0_uk_U85 (.A1( u0_uk_K_r9_31 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n987 ) );
  OAI22_X1 u0_uk_U850 (.ZN( u0_K15_3 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n20 ) , .B2( u0_uk_n36 ) );
  OAI22_X1 u0_uk_U851 (.B1( decrypt ) , .ZN( u0_K5_3 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n477 ) , .B2( u0_uk_n484 ) );
  INV_X1 u0_uk_U852 (.ZN( u0_K13_2 ) , .A( u0_uk_n946 ) );
  AOI22_X1 u0_uk_U853 (.B2( u0_uk_K_r11_26 ) , .A2( u0_uk_K_r11_46 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n946 ) );
  OAI21_X1 u0_uk_U856 (.ZN( u0_K14_3 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n46 ) , .A( u0_uk_n932 ) );
  NAND2_X1 u0_uk_U857 (.A1( u0_uk_K_r12_47 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n932 ) );
  OAI21_X1 u0_uk_U858 (.ZN( u0_K3_3 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n540 ) , .A( u0_uk_n846 ) );
  NAND2_X1 u0_uk_U859 (.A1( u0_uk_K_r1_47 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n846 ) );
  OAI21_X1 u0_uk_U862 (.B1( decrypt ) , .ZN( u0_K7_2 ) , .B2( u0_uk_n404 ) , .A( u0_uk_n773 ) );
  NAND2_X1 u0_uk_U863 (.A1( u0_uk_K_r5_41 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n773 ) );
  OAI21_X1 u0_uk_U864 (.ZN( u0_K10_1 ) , .A( u0_uk_n1021 ) , .B2( u0_uk_n258 ) , .B1( u0_uk_n63 ) );
  NAND2_X1 u0_uk_U865 (.A2( decrypt ) , .A1( u0_uk_K_r8_10 ) , .ZN( u0_uk_n1021 ) );
  OAI22_X1 u0_uk_U867 (.B1( decrypt ) , .ZN( u0_K3_18 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n556 ) , .B2( u0_uk_n563 ) );
  OAI22_X1 u0_uk_U868 (.ZN( u0_K14_22 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n48 ) , .B2( u0_uk_n86 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U869 (.ZN( u0_K10_5 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n246 ) , .B2( u0_uk_n263 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U870 (.B1( decrypt ) , .ZN( u0_K5_41 ) , .A1( u0_uk_n220 ) , .A2( u0_uk_n462 ) , .B2( u0_uk_n470 ) );
  OAI22_X1 u0_uk_U871 (.ZN( u0_K15_22 ) , .A2( u0_uk_n16 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n30 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U872 (.B1( decrypt ) , .ZN( u0_K6_22 ) , .A1( u0_uk_n257 ) , .A2( u0_uk_n436 ) , .B2( u0_uk_n441 ) );
  OAI22_X1 u0_uk_U873 (.ZN( u0_K15_23 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n25 ) , .A2( u0_uk_n7 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U874 (.ZN( u0_K14_23 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n79 ) , .A2( u0_uk_n86 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U875 (.B1( decrypt ) , .ZN( u0_K5_23 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n464 ) , .B2( u0_uk_n473 ) );
  OAI22_X1 u0_uk_U876 (.ZN( u0_K13_34 ) , .A2( u0_uk_n104 ) , .B2( u0_uk_n120 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U877 (.B1( decrypt ) , .ZN( u0_K5_34 ) , .A1( u0_uk_n240 ) , .B2( u0_uk_n474 ) , .A2( u0_uk_n487 ) );
  OAI22_X1 u0_uk_U881 (.ZN( u0_K12_10 ) , .B1( u0_uk_n142 ) , .A2( u0_uk_n149 ) , .B2( u0_uk_n170 ) , .A1( u0_uk_n191 ) );
  OAI22_X1 u0_uk_U882 (.ZN( u0_K12_11 ) , .B2( u0_uk_n149 ) , .A2( u0_uk_n175 ) , .A1( u0_uk_n182 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U885 (.B1( decrypt ) , .ZN( u0_K3_10 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n567 ) , .B2( u0_uk_n572 ) );
  OAI22_X1 u0_uk_U887 (.B1( decrypt ) , .ZN( u0_K13_45 ) , .B2( u0_uk_n133 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n95 ) );
  OAI22_X1 u0_uk_U89 (.ZN( u0_K13_41 ) , .A2( u0_uk_n120 ) , .B2( u0_uk_n135 ) , .A1( u0_uk_n209 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U892 (.B1( decrypt ) , .ZN( u0_K8_1 ) , .A1( u0_uk_n257 ) , .B2( u0_uk_n340 ) , .A2( u0_uk_n356 ) );
  OAI22_X1 u0_uk_U893 (.ZN( u0_K14_6 ) , .A1( u0_uk_n230 ) , .B2( u0_uk_n78 ) , .A2( u0_uk_n85 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U894 (.ZN( u0_K10_3 ) , .A2( u0_uk_n235 ) , .A1( u0_uk_n238 ) , .B2( u0_uk_n255 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U895 (.ZN( u0_K9_3 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n311 ) , .A2( u0_uk_n315 ) );
  OAI22_X1 u0_uk_U899 (.ZN( u0_K14_7 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n53 ) , .B2( u0_uk_n72 ) );
  OAI22_X1 u0_uk_U90 (.ZN( u0_K7_41 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n372 ) , .A2( u0_uk_n402 ) );
  OAI22_X1 u0_uk_U900 (.ZN( u0_K13_24 ) , .B2( u0_uk_n132 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n83 ) , .A2( u0_uk_n91 ) );
  OAI22_X1 u0_uk_U901 (.B1( decrypt ) , .ZN( u0_K6_24 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n427 ) , .B2( u0_uk_n431 ) );
  OAI22_X1 u0_uk_U902 (.ZN( u0_K15_13 ) , .B2( u0_uk_n16 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n44 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U905 (.B1( decrypt ) , .ZN( u0_K5_19 ) , .A1( u0_uk_n161 ) , .B2( u0_uk_n453 ) , .A2( u0_uk_n490 ) );
  OAI22_X1 u0_uk_U906 (.B1( decrypt ) , .ZN( u0_K5_24 ) , .A1( u0_uk_n202 ) , .A2( u0_uk_n461 ) , .B2( u0_uk_n486 ) );
  OAI22_X1 u0_uk_U907 (.ZN( u0_K2_24 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n609 ) , .A2( u0_uk_n624 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U910 (.B1( decrypt ) , .ZN( u0_K16_24 ) , .A1( u0_uk_n162 ) , .A2( u0_uk_n659 ) , .B2( u0_uk_n664 ) );
  OAI22_X1 u0_uk_U911 (.ZN( u0_K7_30 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n367 ) , .B2( u0_uk_n398 ) );
  OAI22_X1 u0_uk_U912 (.B1( decrypt ) , .ZN( u0_K5_13 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n452 ) , .B2( u0_uk_n483 ) );
  OAI22_X1 u0_uk_U913 (.B1( decrypt ) , .ZN( u0_K5_14 ) , .A1( u0_uk_n222 ) , .A2( u0_uk_n478 ) , .B2( u0_uk_n485 ) );
  OAI22_X1 u0_uk_U915 (.ZN( u0_K3_13 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n564 ) , .B2( u0_uk_n569 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U916 (.ZN( u0_K4_36 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n208 ) , .A2( u0_uk_n507 ) , .B2( u0_uk_n512 ) );
  OAI22_X1 u0_uk_U917 (.ZN( u0_K2_17 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n611 ) , .A2( u0_uk_n627 ) );
  OAI22_X1 u0_uk_U920 (.B1( decrypt ) , .ZN( u0_K16_38 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n641 ) , .B2( u0_uk_n648 ) );
  OAI22_X1 u0_uk_U921 (.ZN( u0_K8_38 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n322 ) , .B2( u0_uk_n328 ) );
  OAI22_X1 u0_uk_U922 (.ZN( u0_K7_39 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n365 ) , .B2( u0_uk_n372 ) );
  OAI22_X1 u0_uk_U925 (.ZN( u0_K4_39 ) , .A1( u0_uk_n182 ) , .A2( u0_uk_n516 ) , .B2( u0_uk_n537 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U928 (.ZN( u0_K2_39 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n607 ) , .A2( u0_uk_n622 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U930 (.ZN( u0_K9_23 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n296 ) , .B2( u0_uk_n304 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U932 (.ZN( u0_K12_16 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n165 ) , .A2( u0_uk_n177 ) );
  OAI22_X1 u0_uk_U934 (.A1( decrypt ) , .ZN( u0_K11_48 ) , .A2( u0_uk_n192 ) , .B2( u0_uk_n199 ) , .B1( u0_uk_n202 ) );
  OAI22_X1 u0_uk_U936 (.A1( decrypt ) , .ZN( u0_K9_6 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n295 ) , .B2( u0_uk_n303 ) );
  OAI22_X1 u0_uk_U938 (.ZN( u0_K14_8 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n69 ) , .A2( u0_uk_n87 ) );
  OAI22_X1 u0_uk_U939 (.ZN( u0_K12_18 ) , .A1( u0_uk_n100 ) , .B2( u0_uk_n137 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n175 ) );
  OAI22_X1 u0_uk_U94 (.ZN( u0_K16_5 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n187 ) , .B2( u0_uk_n664 ) , .A2( u0_uk_n667 ) );
  OAI22_X1 u0_uk_U940 (.ZN( u0_K14_20 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n69 ) , .B2( u0_uk_n75 ) , .A1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U941 (.ZN( u0_K2_20 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n238 ) , .B2( u0_uk_n596 ) , .A2( u0_uk_n625 ) );
  OAI22_X1 u0_uk_U943 (.A1( decrypt ) , .ZN( u0_K14_14 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n47 ) , .B2( u0_uk_n54 ) );
  OAI22_X1 u0_uk_U946 (.A1( decrypt ) , .ZN( u0_K15_47 ) , .A2( u0_uk_n2 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n34 ) );
  OAI22_X1 u0_uk_U947 (.ZN( u0_K14_47 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n58 ) , .B2( u0_uk_n68 ) );
  OAI22_X1 u0_uk_U948 (.ZN( u0_K10_46 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n247 ) , .B2( u0_uk_n256 ) );
  OAI22_X1 u0_uk_U949 (.A1( decrypt ) , .ZN( u0_K10_34 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n244 ) , .B2( u0_uk_n270 ) );
  OAI22_X1 u0_uk_U95 (.ZN( u0_K15_5 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n26 ) , .B2( u0_uk_n29 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U951 (.ZN( u0_K6_46 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n417 ) , .A2( u0_uk_n445 ) );
  OAI22_X1 u0_uk_U953 (.A1( decrypt ) , .ZN( u0_K9_4 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n302 ) , .B2( u0_uk_n309 ) );
  OAI22_X1 u0_uk_U954 (.A1( decrypt ) , .ZN( u0_K4_48 ) , .B1( u0_uk_n208 ) , .B2( u0_uk_n505 ) , .A2( u0_uk_n533 ) );
  OAI22_X1 u0_uk_U955 (.A1( decrypt ) , .ZN( u0_K2_48 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n602 ) , .B2( u0_uk_n617 ) );
  OAI22_X1 u0_uk_U958 (.A1( decrypt ) , .ZN( u0_K6_20 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n444 ) , .A2( u0_uk_n449 ) );
  OAI21_X1 u0_uk_U96 (.ZN( u0_K14_5 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n62 ) , .A( u0_uk_n927 ) );
  OAI22_X1 u0_uk_U960 (.A1( decrypt ) , .ZN( u0_K14_18 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n62 ) , .B2( u0_uk_n70 ) );
  OAI22_X1 u0_uk_U961 (.A1( decrypt ) , .ZN( u0_K16_19 ) , .B1( u0_uk_n187 ) , .A2( u0_uk_n630 ) , .B2( u0_uk_n668 ) );
  OAI22_X1 u0_uk_U962 (.ZN( u0_K15_19 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n37 ) , .A2( u0_uk_n7 ) );
  OAI22_X1 u0_uk_U963 (.A1( decrypt ) , .ZN( u0_K10_20 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n229 ) , .B2( u0_uk_n259 ) );
  OAI22_X1 u0_uk_U964 (.ZN( u0_K14_16 ) , .A1( u0_uk_n17 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n46 ) , .A2( u0_uk_n84 ) );
  OAI22_X1 u0_uk_U966 (.ZN( u0_K14_38 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n65 ) , .A2( u0_uk_n81 ) );
  OAI22_X1 u0_uk_U967 (.ZN( u0_K13_38 ) , .B2( u0_uk_n103 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n97 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U968 (.ZN( u0_K2_38 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n593 ) , .B2( u0_uk_n612 ) );
  OAI22_X1 u0_uk_U969 (.ZN( u0_K7_37 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n365 ) , .B2( u0_uk_n389 ) );
  NAND2_X1 u0_uk_U97 (.A1( u0_uk_K_r12_10 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n927 ) );
  OAI22_X1 u0_uk_U970 (.ZN( u0_K2_37 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n594 ) , .A2( u0_uk_n621 ) );
  OAI22_X1 u0_uk_U971 (.A1( decrypt ) , .ZN( u0_K9_40 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n282 ) , .B2( u0_uk_n288 ) );
  OAI22_X1 u0_uk_U972 (.ZN( u0_K5_40 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n458 ) , .B2( u0_uk_n475 ) );
  OAI22_X1 u0_uk_U974 (.A1( decrypt ) , .ZN( u0_K8_45 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n322 ) , .B2( u0_uk_n360 ) );
  OAI22_X1 u0_uk_U976 (.ZN( u0_K7_45 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n381 ) , .B2( u0_uk_n398 ) );
  OAI22_X1 u0_uk_U978 (.ZN( u0_K4_45 ) , .B1( u0_uk_n163 ) , .A1( u0_uk_n27 ) , .A2( u0_uk_n498 ) , .B2( u0_uk_n537 ) );
  OAI22_X1 u0_uk_U979 (.A1( decrypt ) , .ZN( u0_K2_45 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n584 ) , .B2( u0_uk_n606 ) );
  INV_X1 u0_uk_U98 (.ZN( u0_K13_5 ) , .A( u0_uk_n941 ) );
  OAI22_X1 u0_uk_U980 (.ZN( u0_K2_3 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n604 ) , .B2( u0_uk_n619 ) );
  OAI22_X1 u0_uk_U981 (.ZN( u0_K6_3 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n427 ) , .B2( u0_uk_n441 ) );
  OAI22_X1 u0_uk_U982 (.ZN( u0_K3_6 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n571 ) , .A2( u0_uk_n576 ) );
  OAI22_X1 u0_uk_U986 (.A1( decrypt ) , .ZN( u0_K9_15 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n304 ) , .B2( u0_uk_n311 ) );
  OAI22_X1 u0_uk_U987 (.ZN( u0_K6_15 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n423 ) , .B2( u0_uk_n435 ) );
  OAI22_X1 u0_uk_U989 (.ZN( u0_K14_25 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n82 ) , .B2( u0_uk_n88 ) );
  AOI22_X1 u0_uk_U99 (.B2( u0_uk_K_r11_48 ) , .A2( u0_uk_K_r11_53 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n941 ) );
  OAI22_X1 u0_uk_U990 (.A1( decrypt ) , .ZN( u0_K1_23 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n684 ) , .B2( u0_uk_n691 ) );
  OAI21_X1 u0_uk_U994 (.B1( decrypt ) , .ZN( u0_K7_22 ) , .B2( u0_uk_n390 ) , .A( u0_uk_n778 ) );
  NAND2_X1 u0_uk_U995 (.A1( u0_uk_K_r5_5 ) , .ZN( u0_uk_n778 ) , .A2( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U996 (.B1( decrypt ) , .ZN( u0_K7_23 ) , .B2( u0_uk_n405 ) , .A( u0_uk_n777 ) );
  NAND2_X1 u0_uk_U997 (.A1( u0_uk_K_r5_13 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n777 ) );
  DFF_X1 u1_L0_reg_1 (.CK( clk ) , .Q( u1_L0_1 ) , .D( u1_desIn_r_7 ) );
  DFF_X1 u1_L0_reg_10 (.CK( clk ) , .Q( u1_L0_10 ) , .D( u1_desIn_r_13 ) );
  DFF_X1 u1_L0_reg_11 (.CK( clk ) , .Q( u1_L0_11 ) , .D( u1_desIn_r_21 ) );
  DFF_X1 u1_L0_reg_12 (.CK( clk ) , .Q( u1_L0_12 ) , .D( u1_desIn_r_29 ) );
  DFF_X1 u1_L0_reg_13 (.CK( clk ) , .Q( u1_L0_13 ) , .D( u1_desIn_r_37 ) );
  DFF_X1 u1_L0_reg_14 (.CK( clk ) , .Q( u1_L0_14 ) , .D( u1_desIn_r_45 ) );
  DFF_X1 u1_L0_reg_15 (.CK( clk ) , .Q( u1_L0_15 ) , .D( u1_desIn_r_53 ) );
  DFF_X1 u1_L0_reg_16 (.CK( clk ) , .Q( u1_L0_16 ) , .D( u1_desIn_r_61 ) );
  DFF_X1 u1_L0_reg_17 (.CK( clk ) , .Q( u1_L0_17 ) , .D( u1_desIn_r_3 ) );
  DFF_X1 u1_L0_reg_18 (.CK( clk ) , .Q( u1_L0_18 ) , .D( u1_desIn_r_11 ) );
  DFF_X1 u1_L0_reg_19 (.CK( clk ) , .Q( u1_L0_19 ) , .D( u1_desIn_r_19 ) );
  DFF_X1 u1_L0_reg_2 (.CK( clk ) , .Q( u1_L0_2 ) , .D( u1_desIn_r_15 ) );
  DFF_X1 u1_L0_reg_20 (.CK( clk ) , .Q( u1_L0_20 ) , .D( u1_desIn_r_27 ) );
  DFF_X1 u1_L0_reg_21 (.CK( clk ) , .Q( u1_L0_21 ) , .D( u1_desIn_r_35 ) );
  DFF_X1 u1_L0_reg_22 (.CK( clk ) , .Q( u1_L0_22 ) , .D( u1_desIn_r_43 ) );
  DFF_X1 u1_L0_reg_23 (.CK( clk ) , .Q( u1_L0_23 ) , .D( u1_desIn_r_51 ) );
  DFF_X1 u1_L0_reg_24 (.CK( clk ) , .Q( u1_L0_24 ) , .D( u1_desIn_r_59 ) );
  DFF_X1 u1_L0_reg_25 (.CK( clk ) , .Q( u1_L0_25 ) , .D( u1_desIn_r_1 ) );
  DFF_X1 u1_L0_reg_26 (.CK( clk ) , .Q( u1_L0_26 ) , .D( u1_desIn_r_9 ) );
  DFF_X1 u1_L0_reg_27 (.CK( clk ) , .Q( u1_L0_27 ) , .D( u1_desIn_r_17 ) );
  DFF_X1 u1_L0_reg_28 (.CK( clk ) , .Q( u1_L0_28 ) , .D( u1_desIn_r_25 ) );
  DFF_X1 u1_L0_reg_29 (.CK( clk ) , .Q( u1_L0_29 ) , .D( u1_desIn_r_33 ) );
  DFF_X1 u1_L0_reg_3 (.CK( clk ) , .Q( u1_L0_3 ) , .D( u1_desIn_r_23 ) );
  DFF_X1 u1_L0_reg_30 (.CK( clk ) , .Q( u1_L0_30 ) , .D( u1_desIn_r_41 ) );
  DFF_X1 u1_L0_reg_31 (.CK( clk ) , .Q( u1_L0_31 ) , .D( u1_desIn_r_49 ) );
  DFF_X1 u1_L0_reg_32 (.CK( clk ) , .Q( u1_L0_32 ) , .D( u1_desIn_r_57 ) );
  DFF_X1 u1_L0_reg_4 (.CK( clk ) , .Q( u1_L0_4 ) , .D( u1_desIn_r_31 ) );
  DFF_X1 u1_L0_reg_5 (.CK( clk ) , .Q( u1_L0_5 ) , .D( u1_desIn_r_39 ) );
  DFF_X1 u1_L0_reg_6 (.CK( clk ) , .Q( u1_L0_6 ) , .D( u1_desIn_r_47 ) );
  DFF_X1 u1_L0_reg_7 (.CK( clk ) , .Q( u1_L0_7 ) , .D( u1_desIn_r_55 ) );
  DFF_X1 u1_L0_reg_8 (.CK( clk ) , .Q( u1_L0_8 ) , .D( u1_desIn_r_63 ) );
  DFF_X1 u1_L0_reg_9 (.CK( clk ) , .Q( u1_L0_9 ) , .D( u1_desIn_r_5 ) );
  DFF_X1 u1_L10_reg_1 (.CK( clk ) , .Q( u1_L10_1 ) , .D( u1_R9_1 ) );
  DFF_X1 u1_L10_reg_10 (.CK( clk ) , .Q( u1_L10_10 ) , .D( u1_R9_10 ) );
  DFF_X1 u1_L10_reg_11 (.CK( clk ) , .Q( u1_L10_11 ) , .D( u1_R9_11 ) );
  DFF_X1 u1_L10_reg_12 (.CK( clk ) , .Q( u1_L10_12 ) , .D( u1_R9_12 ) );
  DFF_X1 u1_L10_reg_13 (.CK( clk ) , .Q( u1_L10_13 ) , .D( u1_R9_13 ) );
  DFF_X1 u1_L10_reg_14 (.CK( clk ) , .Q( u1_L10_14 ) , .D( u1_R9_14 ) );
  DFF_X1 u1_L10_reg_15 (.CK( clk ) , .Q( u1_L10_15 ) , .D( u1_R9_15 ) );
  DFF_X1 u1_L10_reg_16 (.CK( clk ) , .Q( u1_L10_16 ) , .D( u1_R9_16 ) );
  DFF_X1 u1_L10_reg_17 (.CK( clk ) , .Q( u1_L10_17 ) , .D( u1_R9_17 ) );
  DFF_X1 u1_L10_reg_18 (.CK( clk ) , .Q( u1_L10_18 ) , .D( u1_R9_18 ) );
  DFF_X1 u1_L10_reg_19 (.CK( clk ) , .Q( u1_L10_19 ) , .D( u1_R9_19 ) );
  DFF_X1 u1_L10_reg_2 (.CK( clk ) , .Q( u1_L10_2 ) , .D( u1_R9_2 ) );
  DFF_X1 u1_L10_reg_20 (.CK( clk ) , .Q( u1_L10_20 ) , .D( u1_R9_20 ) );
  DFF_X1 u1_L10_reg_21 (.CK( clk ) , .Q( u1_L10_21 ) , .D( u1_R9_21 ) );
  DFF_X1 u1_L10_reg_22 (.CK( clk ) , .Q( u1_L10_22 ) , .D( u1_R9_22 ) );
  DFF_X1 u1_L10_reg_23 (.CK( clk ) , .Q( u1_L10_23 ) , .D( u1_R9_23 ) );
  DFF_X1 u1_L10_reg_24 (.CK( clk ) , .Q( u1_L10_24 ) , .D( u1_R9_24 ) );
  DFF_X1 u1_L10_reg_25 (.CK( clk ) , .Q( u1_L10_25 ) , .D( u1_R9_25 ) );
  DFF_X1 u1_L10_reg_26 (.CK( clk ) , .Q( u1_L10_26 ) , .D( u1_R9_26 ) );
  DFF_X1 u1_L10_reg_27 (.CK( clk ) , .Q( u1_L10_27 ) , .D( u1_R9_27 ) );
  DFF_X1 u1_L10_reg_28 (.CK( clk ) , .Q( u1_L10_28 ) , .D( u1_R9_28 ) );
  DFF_X1 u1_L10_reg_29 (.CK( clk ) , .Q( u1_L10_29 ) , .D( u1_R9_29 ) );
  DFF_X1 u1_L10_reg_3 (.CK( clk ) , .Q( u1_L10_3 ) , .D( u1_R9_3 ) );
  DFF_X1 u1_L10_reg_30 (.CK( clk ) , .Q( u1_L10_30 ) , .D( u1_R9_30 ) );
  DFF_X1 u1_L10_reg_31 (.CK( clk ) , .Q( u1_L10_31 ) , .D( u1_R9_31 ) );
  DFF_X1 u1_L10_reg_32 (.CK( clk ) , .Q( u1_L10_32 ) , .D( u1_R9_32 ) );
  DFF_X1 u1_L10_reg_4 (.CK( clk ) , .Q( u1_L10_4 ) , .D( u1_R9_4 ) );
  DFF_X1 u1_L10_reg_5 (.CK( clk ) , .Q( u1_L10_5 ) , .D( u1_R9_5 ) );
  DFF_X1 u1_L10_reg_6 (.CK( clk ) , .Q( u1_L10_6 ) , .D( u1_R9_6 ) );
  DFF_X1 u1_L10_reg_7 (.CK( clk ) , .Q( u1_L10_7 ) , .D( u1_R9_7 ) );
  DFF_X1 u1_L10_reg_8 (.CK( clk ) , .Q( u1_L10_8 ) , .D( u1_R9_8 ) );
  DFF_X1 u1_L10_reg_9 (.CK( clk ) , .Q( u1_L10_9 ) , .D( u1_R9_9 ) );
  DFF_X1 u1_L11_reg_1 (.CK( clk ) , .Q( u1_L11_1 ) , .D( u1_R10_1 ) );
  DFF_X1 u1_L11_reg_10 (.CK( clk ) , .Q( u1_L11_10 ) , .D( u1_R10_10 ) );
  DFF_X1 u1_L11_reg_11 (.CK( clk ) , .Q( u1_L11_11 ) , .D( u1_R10_11 ) );
  DFF_X1 u1_L11_reg_12 (.CK( clk ) , .Q( u1_L11_12 ) , .D( u1_R10_12 ) );
  DFF_X1 u1_L11_reg_13 (.CK( clk ) , .Q( u1_L11_13 ) , .D( u1_R10_13 ) );
  DFF_X1 u1_L11_reg_14 (.CK( clk ) , .Q( u1_L11_14 ) , .D( u1_R10_14 ) );
  DFF_X1 u1_L11_reg_15 (.CK( clk ) , .Q( u1_L11_15 ) , .D( u1_R10_15 ) );
  DFF_X1 u1_L11_reg_16 (.CK( clk ) , .Q( u1_L11_16 ) , .D( u1_R10_16 ) );
  DFF_X1 u1_L11_reg_17 (.CK( clk ) , .Q( u1_L11_17 ) , .D( u1_R10_17 ) );
  DFF_X1 u1_L11_reg_18 (.CK( clk ) , .Q( u1_L11_18 ) , .D( u1_R10_18 ) );
  DFF_X1 u1_L11_reg_19 (.CK( clk ) , .Q( u1_L11_19 ) , .D( u1_R10_19 ) );
  DFF_X1 u1_L11_reg_2 (.CK( clk ) , .Q( u1_L11_2 ) , .D( u1_R10_2 ) );
  DFF_X1 u1_L11_reg_20 (.CK( clk ) , .Q( u1_L11_20 ) , .D( u1_R10_20 ) );
  DFF_X1 u1_L11_reg_21 (.CK( clk ) , .Q( u1_L11_21 ) , .D( u1_R10_21 ) );
  DFF_X1 u1_L11_reg_22 (.CK( clk ) , .Q( u1_L11_22 ) , .D( u1_R10_22 ) );
  DFF_X1 u1_L11_reg_23 (.CK( clk ) , .Q( u1_L11_23 ) , .D( u1_R10_23 ) );
  DFF_X1 u1_L11_reg_24 (.CK( clk ) , .Q( u1_L11_24 ) , .D( u1_R10_24 ) );
  DFF_X1 u1_L11_reg_25 (.CK( clk ) , .Q( u1_L11_25 ) , .D( u1_R10_25 ) );
  DFF_X1 u1_L11_reg_26 (.CK( clk ) , .Q( u1_L11_26 ) , .D( u1_R10_26 ) );
  DFF_X1 u1_L11_reg_27 (.CK( clk ) , .Q( u1_L11_27 ) , .D( u1_R10_27 ) );
  DFF_X1 u1_L11_reg_28 (.CK( clk ) , .Q( u1_L11_28 ) , .D( u1_R10_28 ) );
  DFF_X1 u1_L11_reg_29 (.CK( clk ) , .Q( u1_L11_29 ) , .D( u1_R10_29 ) );
  DFF_X1 u1_L11_reg_3 (.CK( clk ) , .Q( u1_L11_3 ) , .D( u1_R10_3 ) );
  DFF_X1 u1_L11_reg_30 (.CK( clk ) , .Q( u1_L11_30 ) , .D( u1_R10_30 ) );
  DFF_X1 u1_L11_reg_31 (.CK( clk ) , .Q( u1_L11_31 ) , .D( u1_R10_31 ) );
  DFF_X1 u1_L11_reg_32 (.CK( clk ) , .Q( u1_L11_32 ) , .D( u1_R10_32 ) );
  DFF_X1 u1_L11_reg_4 (.CK( clk ) , .Q( u1_L11_4 ) , .D( u1_R10_4 ) );
  DFF_X1 u1_L11_reg_5 (.CK( clk ) , .Q( u1_L11_5 ) , .D( u1_R10_5 ) );
  DFF_X1 u1_L11_reg_6 (.CK( clk ) , .Q( u1_L11_6 ) , .D( u1_R10_6 ) );
  DFF_X1 u1_L11_reg_7 (.CK( clk ) , .Q( u1_L11_7 ) , .D( u1_R10_7 ) );
  DFF_X1 u1_L11_reg_8 (.CK( clk ) , .Q( u1_L11_8 ) , .D( u1_R10_8 ) );
  DFF_X1 u1_L11_reg_9 (.CK( clk ) , .Q( u1_L11_9 ) , .D( u1_R10_9 ) );
  DFF_X1 u1_L12_reg_1 (.CK( clk ) , .Q( u1_L12_1 ) , .D( u1_R11_1 ) );
  DFF_X1 u1_L12_reg_10 (.CK( clk ) , .Q( u1_L12_10 ) , .D( u1_R11_10 ) );
  DFF_X1 u1_L12_reg_11 (.CK( clk ) , .Q( u1_L12_11 ) , .D( u1_R11_11 ) );
  DFF_X1 u1_L12_reg_12 (.CK( clk ) , .Q( u1_L12_12 ) , .D( u1_R11_12 ) );
  DFF_X1 u1_L12_reg_13 (.CK( clk ) , .Q( u1_L12_13 ) , .D( u1_R11_13 ) );
  DFF_X1 u1_L12_reg_14 (.CK( clk ) , .Q( u1_L12_14 ) , .D( u1_R11_14 ) );
  DFF_X1 u1_L12_reg_15 (.CK( clk ) , .Q( u1_L12_15 ) , .D( u1_R11_15 ) );
  DFF_X1 u1_L12_reg_16 (.CK( clk ) , .Q( u1_L12_16 ) , .D( u1_R11_16 ) );
  DFF_X1 u1_L12_reg_17 (.CK( clk ) , .Q( u1_L12_17 ) , .D( u1_R11_17 ) );
  DFF_X1 u1_L12_reg_18 (.CK( clk ) , .Q( u1_L12_18 ) , .D( u1_R11_18 ) );
  DFF_X1 u1_L12_reg_19 (.CK( clk ) , .Q( u1_L12_19 ) , .D( u1_R11_19 ) );
  DFF_X1 u1_L12_reg_2 (.CK( clk ) , .Q( u1_L12_2 ) , .D( u1_R11_2 ) );
  DFF_X1 u1_L12_reg_20 (.CK( clk ) , .Q( u1_L12_20 ) , .D( u1_R11_20 ) );
  DFF_X1 u1_L12_reg_21 (.CK( clk ) , .Q( u1_L12_21 ) , .D( u1_R11_21 ) );
  DFF_X1 u1_L12_reg_22 (.CK( clk ) , .Q( u1_L12_22 ) , .D( u1_R11_22 ) );
  DFF_X1 u1_L12_reg_23 (.CK( clk ) , .Q( u1_L12_23 ) , .D( u1_R11_23 ) );
  DFF_X1 u1_L12_reg_24 (.CK( clk ) , .Q( u1_L12_24 ) , .D( u1_R11_24 ) );
  DFF_X1 u1_L12_reg_25 (.CK( clk ) , .Q( u1_L12_25 ) , .D( u1_R11_25 ) );
  DFF_X1 u1_L12_reg_26 (.CK( clk ) , .Q( u1_L12_26 ) , .D( u1_R11_26 ) );
  DFF_X1 u1_L12_reg_27 (.CK( clk ) , .Q( u1_L12_27 ) , .D( u1_R11_27 ) );
  DFF_X1 u1_L12_reg_28 (.CK( clk ) , .Q( u1_L12_28 ) , .D( u1_R11_28 ) );
  DFF_X1 u1_L12_reg_29 (.CK( clk ) , .Q( u1_L12_29 ) , .D( u1_R11_29 ) );
  DFF_X1 u1_L12_reg_3 (.CK( clk ) , .Q( u1_L12_3 ) , .D( u1_R11_3 ) );
  DFF_X1 u1_L12_reg_30 (.CK( clk ) , .Q( u1_L12_30 ) , .D( u1_R11_30 ) );
  DFF_X1 u1_L12_reg_31 (.CK( clk ) , .Q( u1_L12_31 ) , .D( u1_R11_31 ) );
  DFF_X1 u1_L12_reg_32 (.CK( clk ) , .Q( u1_L12_32 ) , .D( u1_R11_32 ) );
  DFF_X1 u1_L12_reg_4 (.CK( clk ) , .Q( u1_L12_4 ) , .D( u1_R11_4 ) );
  DFF_X1 u1_L12_reg_5 (.CK( clk ) , .Q( u1_L12_5 ) , .D( u1_R11_5 ) );
  DFF_X1 u1_L12_reg_6 (.CK( clk ) , .Q( u1_L12_6 ) , .D( u1_R11_6 ) );
  DFF_X1 u1_L12_reg_7 (.CK( clk ) , .Q( u1_L12_7 ) , .D( u1_R11_7 ) );
  DFF_X1 u1_L12_reg_8 (.CK( clk ) , .Q( u1_L12_8 ) , .D( u1_R11_8 ) );
  DFF_X1 u1_L12_reg_9 (.CK( clk ) , .Q( u1_L12_9 ) , .D( u1_R11_9 ) );
  DFF_X1 u1_L13_reg_1 (.CK( clk ) , .Q( u1_L13_1 ) , .D( u1_R12_1 ) );
  DFF_X1 u1_L13_reg_10 (.CK( clk ) , .Q( u1_L13_10 ) , .D( u1_R12_10 ) );
  DFF_X1 u1_L13_reg_11 (.CK( clk ) , .Q( u1_L13_11 ) , .D( u1_R12_11 ) );
  DFF_X1 u1_L13_reg_12 (.CK( clk ) , .Q( u1_L13_12 ) , .D( u1_R12_12 ) );
  DFF_X1 u1_L13_reg_13 (.CK( clk ) , .Q( u1_L13_13 ) , .D( u1_R12_13 ) );
  DFF_X1 u1_L13_reg_14 (.CK( clk ) , .Q( u1_L13_14 ) , .D( u1_R12_14 ) );
  DFF_X1 u1_L13_reg_15 (.CK( clk ) , .Q( u1_L13_15 ) , .D( u1_R12_15 ) );
  DFF_X1 u1_L13_reg_16 (.CK( clk ) , .Q( u1_L13_16 ) , .D( u1_R12_16 ) );
  DFF_X1 u1_L13_reg_17 (.CK( clk ) , .Q( u1_L13_17 ) , .D( u1_R12_17 ) );
  DFF_X1 u1_L13_reg_18 (.CK( clk ) , .Q( u1_L13_18 ) , .D( u1_R12_18 ) );
  DFF_X1 u1_L13_reg_19 (.CK( clk ) , .Q( u1_L13_19 ) , .D( u1_R12_19 ) );
  DFF_X1 u1_L13_reg_2 (.CK( clk ) , .Q( u1_L13_2 ) , .D( u1_R12_2 ) );
  DFF_X1 u1_L13_reg_20 (.CK( clk ) , .Q( u1_L13_20 ) , .D( u1_R12_20 ) );
  DFF_X1 u1_L13_reg_21 (.CK( clk ) , .Q( u1_L13_21 ) , .D( u1_R12_21 ) );
  DFF_X1 u1_L13_reg_22 (.CK( clk ) , .Q( u1_L13_22 ) , .D( u1_R12_22 ) );
  DFF_X1 u1_L13_reg_23 (.CK( clk ) , .Q( u1_L13_23 ) , .D( u1_R12_23 ) );
  DFF_X1 u1_L13_reg_24 (.CK( clk ) , .Q( u1_L13_24 ) , .D( u1_R12_24 ) );
  DFF_X1 u1_L13_reg_25 (.CK( clk ) , .Q( u1_L13_25 ) , .D( u1_R12_25 ) );
  DFF_X1 u1_L13_reg_26 (.CK( clk ) , .Q( u1_L13_26 ) , .D( u1_R12_26 ) );
  DFF_X1 u1_L13_reg_27 (.CK( clk ) , .Q( u1_L13_27 ) , .D( u1_R12_27 ) );
  DFF_X1 u1_L13_reg_28 (.CK( clk ) , .Q( u1_L13_28 ) , .D( u1_R12_28 ) );
  DFF_X1 u1_L13_reg_29 (.CK( clk ) , .Q( u1_L13_29 ) , .D( u1_R12_29 ) );
  DFF_X1 u1_L13_reg_3 (.CK( clk ) , .Q( u1_L13_3 ) , .D( u1_R12_3 ) );
  DFF_X1 u1_L13_reg_30 (.CK( clk ) , .Q( u1_L13_30 ) , .D( u1_R12_30 ) );
  DFF_X1 u1_L13_reg_31 (.CK( clk ) , .Q( u1_L13_31 ) , .D( u1_R12_31 ) );
  DFF_X1 u1_L13_reg_32 (.CK( clk ) , .Q( u1_L13_32 ) , .D( u1_R12_32 ) );
  DFF_X1 u1_L13_reg_4 (.CK( clk ) , .Q( u1_L13_4 ) , .D( u1_R12_4 ) );
  DFF_X1 u1_L13_reg_5 (.CK( clk ) , .Q( u1_L13_5 ) , .D( u1_R12_5 ) );
  DFF_X1 u1_L13_reg_6 (.CK( clk ) , .Q( u1_L13_6 ) , .D( u1_R12_6 ) );
  DFF_X1 u1_L13_reg_7 (.CK( clk ) , .Q( u1_L13_7 ) , .D( u1_R12_7 ) );
  DFF_X1 u1_L13_reg_8 (.CK( clk ) , .Q( u1_L13_8 ) , .D( u1_R12_8 ) );
  DFF_X1 u1_L13_reg_9 (.CK( clk ) , .Q( u1_L13_9 ) , .D( u1_R12_9 ) );
  DFF_X1 u1_L14_reg_1 (.CK( clk ) , .Q( u1_L14_1 ) , .D( u1_R13_1 ) );
  DFF_X1 u1_L14_reg_10 (.CK( clk ) , .Q( u1_L14_10 ) , .D( u1_R13_10 ) );
  DFF_X1 u1_L14_reg_11 (.CK( clk ) , .Q( u1_L14_11 ) , .D( u1_R13_11 ) );
  DFF_X1 u1_L14_reg_12 (.CK( clk ) , .Q( u1_L14_12 ) , .D( u1_R13_12 ) );
  DFF_X1 u1_L14_reg_13 (.CK( clk ) , .Q( u1_L14_13 ) , .D( u1_R13_13 ) );
  DFF_X1 u1_L14_reg_14 (.CK( clk ) , .Q( u1_L14_14 ) , .D( u1_R13_14 ) );
  DFF_X1 u1_L14_reg_15 (.CK( clk ) , .Q( u1_L14_15 ) , .D( u1_R13_15 ) );
  DFF_X1 u1_L14_reg_16 (.CK( clk ) , .Q( u1_L14_16 ) , .D( u1_R13_16 ) );
  DFF_X1 u1_L14_reg_17 (.CK( clk ) , .Q( u1_L14_17 ) , .D( u1_R13_17 ) );
  DFF_X1 u1_L14_reg_18 (.CK( clk ) , .Q( u1_L14_18 ) , .D( u1_R13_18 ) );
  DFF_X1 u1_L14_reg_19 (.CK( clk ) , .Q( u1_L14_19 ) , .D( u1_R13_19 ) );
  DFF_X1 u1_L14_reg_2 (.CK( clk ) , .Q( u1_L14_2 ) , .D( u1_R13_2 ) );
  DFF_X1 u1_L14_reg_20 (.CK( clk ) , .Q( u1_L14_20 ) , .D( u1_R13_20 ) );
  DFF_X1 u1_L14_reg_21 (.CK( clk ) , .Q( u1_L14_21 ) , .D( u1_R13_21 ) );
  DFF_X1 u1_L14_reg_22 (.CK( clk ) , .Q( u1_L14_22 ) , .D( u1_R13_22 ) );
  DFF_X1 u1_L14_reg_23 (.CK( clk ) , .Q( u1_L14_23 ) , .D( u1_R13_23 ) );
  DFF_X1 u1_L14_reg_24 (.CK( clk ) , .Q( u1_L14_24 ) , .D( u1_R13_24 ) );
  DFF_X1 u1_L14_reg_25 (.CK( clk ) , .Q( u1_L14_25 ) , .D( u1_R13_25 ) );
  DFF_X1 u1_L14_reg_26 (.CK( clk ) , .Q( u1_L14_26 ) , .D( u1_R13_26 ) );
  DFF_X1 u1_L14_reg_27 (.CK( clk ) , .Q( u1_L14_27 ) , .D( u1_R13_27 ) );
  DFF_X1 u1_L14_reg_28 (.CK( clk ) , .Q( u1_L14_28 ) , .D( u1_R13_28 ) );
  DFF_X1 u1_L14_reg_29 (.CK( clk ) , .Q( u1_L14_29 ) , .D( u1_R13_29 ) );
  DFF_X1 u1_L14_reg_3 (.CK( clk ) , .Q( u1_L14_3 ) , .D( u1_R13_3 ) );
  DFF_X1 u1_L14_reg_30 (.CK( clk ) , .Q( u1_L14_30 ) , .D( u1_R13_30 ) );
  DFF_X1 u1_L14_reg_31 (.CK( clk ) , .Q( u1_L14_31 ) , .D( u1_R13_31 ) );
  DFF_X1 u1_L14_reg_32 (.CK( clk ) , .Q( u1_L14_32 ) , .D( u1_R13_32 ) );
  DFF_X1 u1_L14_reg_4 (.CK( clk ) , .Q( u1_L14_4 ) , .D( u1_R13_4 ) );
  DFF_X1 u1_L14_reg_5 (.CK( clk ) , .Q( u1_L14_5 ) , .D( u1_R13_5 ) );
  DFF_X1 u1_L14_reg_6 (.CK( clk ) , .Q( u1_L14_6 ) , .D( u1_R13_6 ) );
  DFF_X1 u1_L14_reg_7 (.CK( clk ) , .Q( u1_L14_7 ) , .D( u1_R13_7 ) );
  DFF_X1 u1_L14_reg_8 (.CK( clk ) , .Q( u1_L14_8 ) , .D( u1_R13_8 ) );
  DFF_X1 u1_L14_reg_9 (.CK( clk ) , .Q( u1_L14_9 ) , .D( u1_R13_9 ) );
  DFF_X1 u1_L1_reg_1 (.CK( clk ) , .Q( u1_L1_1 ) , .D( u1_R0_1 ) );
  DFF_X1 u1_L1_reg_10 (.CK( clk ) , .Q( u1_L1_10 ) , .D( u1_R0_10 ) );
  DFF_X1 u1_L1_reg_11 (.CK( clk ) , .Q( u1_L1_11 ) , .D( u1_R0_11 ) );
  DFF_X1 u1_L1_reg_12 (.CK( clk ) , .Q( u1_L1_12 ) , .D( u1_R0_12 ) );
  DFF_X1 u1_L1_reg_13 (.CK( clk ) , .Q( u1_L1_13 ) , .D( u1_R0_13 ) );
  DFF_X1 u1_L1_reg_14 (.CK( clk ) , .Q( u1_L1_14 ) , .D( u1_R0_14 ) );
  DFF_X1 u1_L1_reg_15 (.CK( clk ) , .Q( u1_L1_15 ) , .D( u1_R0_15 ) );
  DFF_X1 u1_L1_reg_16 (.CK( clk ) , .Q( u1_L1_16 ) , .D( u1_R0_16 ) );
  DFF_X1 u1_L1_reg_17 (.CK( clk ) , .Q( u1_L1_17 ) , .D( u1_R0_17 ) );
  DFF_X1 u1_L1_reg_18 (.CK( clk ) , .Q( u1_L1_18 ) , .D( u1_R0_18 ) );
  DFF_X1 u1_L1_reg_19 (.CK( clk ) , .Q( u1_L1_19 ) , .D( u1_R0_19 ) );
  DFF_X1 u1_L1_reg_2 (.CK( clk ) , .Q( u1_L1_2 ) , .D( u1_R0_2 ) );
  DFF_X1 u1_L1_reg_20 (.CK( clk ) , .Q( u1_L1_20 ) , .D( u1_R0_20 ) );
  DFF_X1 u1_L1_reg_21 (.CK( clk ) , .Q( u1_L1_21 ) , .D( u1_R0_21 ) );
  DFF_X1 u1_L1_reg_22 (.CK( clk ) , .Q( u1_L1_22 ) , .D( u1_R0_22 ) );
  DFF_X1 u1_L1_reg_23 (.CK( clk ) , .Q( u1_L1_23 ) , .D( u1_R0_23 ) );
  DFF_X1 u1_L1_reg_24 (.CK( clk ) , .Q( u1_L1_24 ) , .D( u1_R0_24 ) );
  DFF_X1 u1_L1_reg_25 (.CK( clk ) , .Q( u1_L1_25 ) , .D( u1_R0_25 ) );
  DFF_X1 u1_L1_reg_26 (.CK( clk ) , .Q( u1_L1_26 ) , .D( u1_R0_26 ) );
  DFF_X1 u1_L1_reg_27 (.CK( clk ) , .Q( u1_L1_27 ) , .D( u1_R0_27 ) );
  DFF_X1 u1_L1_reg_28 (.CK( clk ) , .Q( u1_L1_28 ) , .D( u1_R0_28 ) );
  DFF_X1 u1_L1_reg_29 (.CK( clk ) , .Q( u1_L1_29 ) , .D( u1_R0_29 ) );
  DFF_X1 u1_L1_reg_3 (.CK( clk ) , .Q( u1_L1_3 ) , .D( u1_R0_3 ) );
  DFF_X1 u1_L1_reg_30 (.CK( clk ) , .Q( u1_L1_30 ) , .D( u1_R0_30 ) );
  DFF_X1 u1_L1_reg_31 (.CK( clk ) , .Q( u1_L1_31 ) , .D( u1_R0_31 ) );
  DFF_X1 u1_L1_reg_32 (.CK( clk ) , .Q( u1_L1_32 ) , .D( u1_R0_32 ) );
  DFF_X1 u1_L1_reg_4 (.CK( clk ) , .Q( u1_L1_4 ) , .D( u1_R0_4 ) );
  DFF_X1 u1_L1_reg_5 (.CK( clk ) , .Q( u1_L1_5 ) , .D( u1_R0_5 ) );
  DFF_X1 u1_L1_reg_6 (.CK( clk ) , .Q( u1_L1_6 ) , .D( u1_R0_6 ) );
  DFF_X1 u1_L1_reg_7 (.CK( clk ) , .Q( u1_L1_7 ) , .D( u1_R0_7 ) );
  DFF_X1 u1_L1_reg_8 (.CK( clk ) , .Q( u1_L1_8 ) , .D( u1_R0_8 ) );
  DFF_X1 u1_L1_reg_9 (.CK( clk ) , .Q( u1_L1_9 ) , .D( u1_R0_9 ) );
  DFF_X1 u1_L2_reg_1 (.CK( clk ) , .Q( u1_L2_1 ) , .D( u1_R1_1 ) );
  DFF_X1 u1_L2_reg_10 (.CK( clk ) , .Q( u1_L2_10 ) , .D( u1_R1_10 ) );
  DFF_X1 u1_L2_reg_11 (.CK( clk ) , .Q( u1_L2_11 ) , .D( u1_R1_11 ) );
  DFF_X1 u1_L2_reg_12 (.CK( clk ) , .Q( u1_L2_12 ) , .D( u1_R1_12 ) );
  DFF_X1 u1_L2_reg_13 (.CK( clk ) , .Q( u1_L2_13 ) , .D( u1_R1_13 ) );
  DFF_X1 u1_L2_reg_14 (.CK( clk ) , .Q( u1_L2_14 ) , .D( u1_R1_14 ) );
  DFF_X1 u1_L2_reg_15 (.CK( clk ) , .Q( u1_L2_15 ) , .D( u1_R1_15 ) );
  DFF_X1 u1_L2_reg_16 (.CK( clk ) , .Q( u1_L2_16 ) , .D( u1_R1_16 ) );
  DFF_X1 u1_L2_reg_17 (.CK( clk ) , .Q( u1_L2_17 ) , .D( u1_R1_17 ) );
  DFF_X1 u1_L2_reg_18 (.CK( clk ) , .Q( u1_L2_18 ) , .D( u1_R1_18 ) );
  DFF_X1 u1_L2_reg_19 (.CK( clk ) , .Q( u1_L2_19 ) , .D( u1_R1_19 ) );
  DFF_X1 u1_L2_reg_2 (.CK( clk ) , .Q( u1_L2_2 ) , .D( u1_R1_2 ) );
  DFF_X1 u1_L2_reg_20 (.CK( clk ) , .Q( u1_L2_20 ) , .D( u1_R1_20 ) );
  DFF_X1 u1_L2_reg_21 (.CK( clk ) , .Q( u1_L2_21 ) , .D( u1_R1_21 ) );
  DFF_X1 u1_L2_reg_22 (.CK( clk ) , .Q( u1_L2_22 ) , .D( u1_R1_22 ) );
  DFF_X1 u1_L2_reg_23 (.CK( clk ) , .Q( u1_L2_23 ) , .D( u1_R1_23 ) );
  DFF_X1 u1_L2_reg_24 (.CK( clk ) , .Q( u1_L2_24 ) , .D( u1_R1_24 ) );
  DFF_X1 u1_L2_reg_25 (.CK( clk ) , .Q( u1_L2_25 ) , .D( u1_R1_25 ) );
  DFF_X1 u1_L2_reg_26 (.CK( clk ) , .Q( u1_L2_26 ) , .D( u1_R1_26 ) );
  DFF_X1 u1_L2_reg_27 (.CK( clk ) , .Q( u1_L2_27 ) , .D( u1_R1_27 ) );
  DFF_X1 u1_L2_reg_28 (.CK( clk ) , .Q( u1_L2_28 ) , .D( u1_R1_28 ) );
  DFF_X1 u1_L2_reg_29 (.CK( clk ) , .Q( u1_L2_29 ) , .D( u1_R1_29 ) );
  DFF_X1 u1_L2_reg_3 (.CK( clk ) , .Q( u1_L2_3 ) , .D( u1_R1_3 ) );
  DFF_X1 u1_L2_reg_30 (.CK( clk ) , .Q( u1_L2_30 ) , .D( u1_R1_30 ) );
  DFF_X1 u1_L2_reg_31 (.CK( clk ) , .Q( u1_L2_31 ) , .D( u1_R1_31 ) );
  DFF_X1 u1_L2_reg_32 (.CK( clk ) , .Q( u1_L2_32 ) , .D( u1_R1_32 ) );
  DFF_X1 u1_L2_reg_4 (.CK( clk ) , .Q( u1_L2_4 ) , .D( u1_R1_4 ) );
  DFF_X1 u1_L2_reg_5 (.CK( clk ) , .Q( u1_L2_5 ) , .D( u1_R1_5 ) );
  DFF_X1 u1_L2_reg_6 (.CK( clk ) , .Q( u1_L2_6 ) , .D( u1_R1_6 ) );
  DFF_X1 u1_L2_reg_7 (.CK( clk ) , .Q( u1_L2_7 ) , .D( u1_R1_7 ) );
  DFF_X1 u1_L2_reg_8 (.CK( clk ) , .Q( u1_L2_8 ) , .D( u1_R1_8 ) );
  DFF_X1 u1_L2_reg_9 (.CK( clk ) , .Q( u1_L2_9 ) , .D( u1_R1_9 ) );
  DFF_X1 u1_L3_reg_1 (.CK( clk ) , .Q( u1_L3_1 ) , .D( u1_R2_1 ) );
  DFF_X1 u1_L3_reg_10 (.CK( clk ) , .Q( u1_L3_10 ) , .D( u1_R2_10 ) );
  DFF_X1 u1_L3_reg_11 (.CK( clk ) , .Q( u1_L3_11 ) , .D( u1_R2_11 ) );
  DFF_X1 u1_L3_reg_12 (.CK( clk ) , .Q( u1_L3_12 ) , .D( u1_R2_12 ) );
  DFF_X1 u1_L3_reg_13 (.CK( clk ) , .Q( u1_L3_13 ) , .D( u1_R2_13 ) );
  DFF_X1 u1_L3_reg_14 (.CK( clk ) , .Q( u1_L3_14 ) , .D( u1_R2_14 ) );
  DFF_X1 u1_L3_reg_15 (.CK( clk ) , .Q( u1_L3_15 ) , .D( u1_R2_15 ) );
  DFF_X1 u1_L3_reg_16 (.CK( clk ) , .Q( u1_L3_16 ) , .D( u1_R2_16 ) );
  DFF_X1 u1_L3_reg_17 (.CK( clk ) , .Q( u1_L3_17 ) , .D( u1_R2_17 ) );
  DFF_X1 u1_L3_reg_18 (.CK( clk ) , .Q( u1_L3_18 ) , .D( u1_R2_18 ) );
  DFF_X1 u1_L3_reg_19 (.CK( clk ) , .Q( u1_L3_19 ) , .D( u1_R2_19 ) );
  DFF_X1 u1_L3_reg_2 (.CK( clk ) , .Q( u1_L3_2 ) , .D( u1_R2_2 ) );
  DFF_X1 u1_L3_reg_20 (.CK( clk ) , .Q( u1_L3_20 ) , .D( u1_R2_20 ) );
  DFF_X1 u1_L3_reg_21 (.CK( clk ) , .Q( u1_L3_21 ) , .D( u1_R2_21 ) );
  DFF_X1 u1_L3_reg_22 (.CK( clk ) , .Q( u1_L3_22 ) , .D( u1_R2_22 ) );
  DFF_X1 u1_L3_reg_23 (.CK( clk ) , .Q( u1_L3_23 ) , .D( u1_R2_23 ) );
  DFF_X1 u1_L3_reg_24 (.CK( clk ) , .Q( u1_L3_24 ) , .D( u1_R2_24 ) );
  DFF_X1 u1_L3_reg_25 (.CK( clk ) , .Q( u1_L3_25 ) , .D( u1_R2_25 ) );
  DFF_X1 u1_L3_reg_26 (.CK( clk ) , .Q( u1_L3_26 ) , .D( u1_R2_26 ) );
  DFF_X1 u1_L3_reg_27 (.CK( clk ) , .Q( u1_L3_27 ) , .D( u1_R2_27 ) );
  DFF_X1 u1_L3_reg_28 (.CK( clk ) , .Q( u1_L3_28 ) , .D( u1_R2_28 ) );
  DFF_X1 u1_L3_reg_29 (.CK( clk ) , .Q( u1_L3_29 ) , .D( u1_R2_29 ) );
  DFF_X1 u1_L3_reg_3 (.CK( clk ) , .Q( u1_L3_3 ) , .D( u1_R2_3 ) );
  DFF_X1 u1_L3_reg_30 (.CK( clk ) , .Q( u1_L3_30 ) , .D( u1_R2_30 ) );
  DFF_X1 u1_L3_reg_31 (.CK( clk ) , .Q( u1_L3_31 ) , .D( u1_R2_31 ) );
  DFF_X1 u1_L3_reg_32 (.CK( clk ) , .Q( u1_L3_32 ) , .D( u1_R2_32 ) );
  DFF_X1 u1_L3_reg_4 (.CK( clk ) , .Q( u1_L3_4 ) , .D( u1_R2_4 ) );
  DFF_X1 u1_L3_reg_5 (.CK( clk ) , .Q( u1_L3_5 ) , .D( u1_R2_5 ) );
  DFF_X1 u1_L3_reg_6 (.CK( clk ) , .Q( u1_L3_6 ) , .D( u1_R2_6 ) );
  DFF_X1 u1_L3_reg_7 (.CK( clk ) , .Q( u1_L3_7 ) , .D( u1_R2_7 ) );
  DFF_X1 u1_L3_reg_8 (.CK( clk ) , .Q( u1_L3_8 ) , .D( u1_R2_8 ) );
  DFF_X1 u1_L3_reg_9 (.CK( clk ) , .Q( u1_L3_9 ) , .D( u1_R2_9 ) );
  DFF_X1 u1_L4_reg_1 (.CK( clk ) , .Q( u1_L4_1 ) , .D( u1_R3_1 ) );
  DFF_X1 u1_L4_reg_10 (.CK( clk ) , .Q( u1_L4_10 ) , .D( u1_R3_10 ) );
  DFF_X1 u1_L4_reg_11 (.CK( clk ) , .Q( u1_L4_11 ) , .D( u1_R3_11 ) );
  DFF_X1 u1_L4_reg_12 (.CK( clk ) , .Q( u1_L4_12 ) , .D( u1_R3_12 ) );
  DFF_X1 u1_L4_reg_13 (.CK( clk ) , .Q( u1_L4_13 ) , .D( u1_R3_13 ) );
  DFF_X1 u1_L4_reg_14 (.CK( clk ) , .Q( u1_L4_14 ) , .D( u1_R3_14 ) );
  DFF_X1 u1_L4_reg_15 (.CK( clk ) , .Q( u1_L4_15 ) , .D( u1_R3_15 ) );
  DFF_X1 u1_L4_reg_16 (.CK( clk ) , .Q( u1_L4_16 ) , .D( u1_R3_16 ) );
  DFF_X1 u1_L4_reg_17 (.CK( clk ) , .Q( u1_L4_17 ) , .D( u1_R3_17 ) );
  DFF_X1 u1_L4_reg_18 (.CK( clk ) , .Q( u1_L4_18 ) , .D( u1_R3_18 ) );
  DFF_X1 u1_L4_reg_19 (.CK( clk ) , .Q( u1_L4_19 ) , .D( u1_R3_19 ) );
  DFF_X1 u1_L4_reg_2 (.CK( clk ) , .Q( u1_L4_2 ) , .D( u1_R3_2 ) );
  DFF_X1 u1_L4_reg_20 (.CK( clk ) , .Q( u1_L4_20 ) , .D( u1_R3_20 ) );
  DFF_X1 u1_L4_reg_21 (.CK( clk ) , .Q( u1_L4_21 ) , .D( u1_R3_21 ) );
  DFF_X1 u1_L4_reg_22 (.CK( clk ) , .Q( u1_L4_22 ) , .D( u1_R3_22 ) );
  DFF_X1 u1_L4_reg_23 (.CK( clk ) , .Q( u1_L4_23 ) , .D( u1_R3_23 ) );
  DFF_X1 u1_L4_reg_24 (.CK( clk ) , .Q( u1_L4_24 ) , .D( u1_R3_24 ) );
  DFF_X1 u1_L4_reg_25 (.CK( clk ) , .Q( u1_L4_25 ) , .D( u1_R3_25 ) );
  DFF_X1 u1_L4_reg_26 (.CK( clk ) , .Q( u1_L4_26 ) , .D( u1_R3_26 ) );
  DFF_X1 u1_L4_reg_27 (.CK( clk ) , .Q( u1_L4_27 ) , .D( u1_R3_27 ) );
  DFF_X1 u1_L4_reg_28 (.CK( clk ) , .Q( u1_L4_28 ) , .D( u1_R3_28 ) );
  DFF_X1 u1_L4_reg_29 (.CK( clk ) , .Q( u1_L4_29 ) , .D( u1_R3_29 ) );
  DFF_X1 u1_L4_reg_3 (.CK( clk ) , .Q( u1_L4_3 ) , .D( u1_R3_3 ) );
  DFF_X1 u1_L4_reg_30 (.CK( clk ) , .Q( u1_L4_30 ) , .D( u1_R3_30 ) );
  DFF_X1 u1_L4_reg_31 (.CK( clk ) , .Q( u1_L4_31 ) , .D( u1_R3_31 ) );
  DFF_X1 u1_L4_reg_32 (.CK( clk ) , .Q( u1_L4_32 ) , .D( u1_R3_32 ) );
  DFF_X1 u1_L4_reg_4 (.CK( clk ) , .Q( u1_L4_4 ) , .D( u1_R3_4 ) );
  DFF_X1 u1_L4_reg_5 (.CK( clk ) , .Q( u1_L4_5 ) , .D( u1_R3_5 ) );
  DFF_X1 u1_L4_reg_6 (.CK( clk ) , .Q( u1_L4_6 ) , .D( u1_R3_6 ) );
  DFF_X1 u1_L4_reg_7 (.CK( clk ) , .Q( u1_L4_7 ) , .D( u1_R3_7 ) );
  DFF_X1 u1_L4_reg_8 (.CK( clk ) , .Q( u1_L4_8 ) , .D( u1_R3_8 ) );
  DFF_X1 u1_L4_reg_9 (.CK( clk ) , .Q( u1_L4_9 ) , .D( u1_R3_9 ) );
  DFF_X1 u1_L5_reg_1 (.CK( clk ) , .Q( u1_L5_1 ) , .D( u1_R4_1 ) );
  DFF_X1 u1_L5_reg_10 (.CK( clk ) , .Q( u1_L5_10 ) , .D( u1_R4_10 ) );
  DFF_X1 u1_L5_reg_11 (.CK( clk ) , .Q( u1_L5_11 ) , .D( u1_R4_11 ) );
  DFF_X1 u1_L5_reg_12 (.CK( clk ) , .Q( u1_L5_12 ) , .D( u1_R4_12 ) );
  DFF_X1 u1_L5_reg_13 (.CK( clk ) , .Q( u1_L5_13 ) , .D( u1_R4_13 ) );
  DFF_X1 u1_L5_reg_14 (.CK( clk ) , .Q( u1_L5_14 ) , .D( u1_R4_14 ) );
  DFF_X1 u1_L5_reg_15 (.CK( clk ) , .Q( u1_L5_15 ) , .D( u1_R4_15 ) );
  DFF_X1 u1_L5_reg_16 (.CK( clk ) , .Q( u1_L5_16 ) , .D( u1_R4_16 ) );
  DFF_X1 u1_L5_reg_17 (.CK( clk ) , .Q( u1_L5_17 ) , .D( u1_R4_17 ) );
  DFF_X1 u1_L5_reg_18 (.CK( clk ) , .Q( u1_L5_18 ) , .D( u1_R4_18 ) );
  DFF_X1 u1_L5_reg_19 (.CK( clk ) , .Q( u1_L5_19 ) , .D( u1_R4_19 ) );
  DFF_X1 u1_L5_reg_2 (.CK( clk ) , .Q( u1_L5_2 ) , .D( u1_R4_2 ) );
  DFF_X1 u1_L5_reg_20 (.CK( clk ) , .Q( u1_L5_20 ) , .D( u1_R4_20 ) );
  DFF_X1 u1_L5_reg_21 (.CK( clk ) , .Q( u1_L5_21 ) , .D( u1_R4_21 ) );
  DFF_X1 u1_L5_reg_22 (.CK( clk ) , .Q( u1_L5_22 ) , .D( u1_R4_22 ) );
  DFF_X1 u1_L5_reg_23 (.CK( clk ) , .Q( u1_L5_23 ) , .D( u1_R4_23 ) );
  DFF_X1 u1_L5_reg_24 (.CK( clk ) , .Q( u1_L5_24 ) , .D( u1_R4_24 ) );
  DFF_X1 u1_L5_reg_25 (.CK( clk ) , .Q( u1_L5_25 ) , .D( u1_R4_25 ) );
  DFF_X1 u1_L5_reg_26 (.CK( clk ) , .Q( u1_L5_26 ) , .D( u1_R4_26 ) );
  DFF_X1 u1_L5_reg_27 (.CK( clk ) , .Q( u1_L5_27 ) , .D( u1_R4_27 ) );
  DFF_X1 u1_L5_reg_28 (.CK( clk ) , .Q( u1_L5_28 ) , .D( u1_R4_28 ) );
  DFF_X1 u1_L5_reg_29 (.CK( clk ) , .Q( u1_L5_29 ) , .D( u1_R4_29 ) );
  DFF_X1 u1_L5_reg_3 (.CK( clk ) , .Q( u1_L5_3 ) , .D( u1_R4_3 ) );
  DFF_X1 u1_L5_reg_30 (.CK( clk ) , .Q( u1_L5_30 ) , .D( u1_R4_30 ) );
  DFF_X1 u1_L5_reg_31 (.CK( clk ) , .Q( u1_L5_31 ) , .D( u1_R4_31 ) );
  DFF_X1 u1_L5_reg_32 (.CK( clk ) , .Q( u1_L5_32 ) , .D( u1_R4_32 ) );
  DFF_X1 u1_L5_reg_4 (.CK( clk ) , .Q( u1_L5_4 ) , .D( u1_R4_4 ) );
  DFF_X1 u1_L5_reg_5 (.CK( clk ) , .Q( u1_L5_5 ) , .D( u1_R4_5 ) );
  DFF_X1 u1_L5_reg_6 (.CK( clk ) , .Q( u1_L5_6 ) , .D( u1_R4_6 ) );
  DFF_X1 u1_L5_reg_7 (.CK( clk ) , .Q( u1_L5_7 ) , .D( u1_R4_7 ) );
  DFF_X1 u1_L5_reg_8 (.CK( clk ) , .Q( u1_L5_8 ) , .D( u1_R4_8 ) );
  DFF_X1 u1_L5_reg_9 (.CK( clk ) , .Q( u1_L5_9 ) , .D( u1_R4_9 ) );
  DFF_X1 u1_L6_reg_1 (.CK( clk ) , .Q( u1_L6_1 ) , .D( u1_R5_1 ) );
  DFF_X1 u1_L6_reg_10 (.CK( clk ) , .Q( u1_L6_10 ) , .D( u1_R5_10 ) );
  DFF_X1 u1_L6_reg_11 (.CK( clk ) , .Q( u1_L6_11 ) , .D( u1_R5_11 ) );
  DFF_X1 u1_L6_reg_12 (.CK( clk ) , .Q( u1_L6_12 ) , .D( u1_R5_12 ) );
  DFF_X1 u1_L6_reg_13 (.CK( clk ) , .Q( u1_L6_13 ) , .D( u1_R5_13 ) );
  DFF_X1 u1_L6_reg_14 (.CK( clk ) , .Q( u1_L6_14 ) , .D( u1_R5_14 ) );
  DFF_X1 u1_L6_reg_15 (.CK( clk ) , .Q( u1_L6_15 ) , .D( u1_R5_15 ) );
  DFF_X1 u1_L6_reg_16 (.CK( clk ) , .Q( u1_L6_16 ) , .D( u1_R5_16 ) );
  DFF_X1 u1_L6_reg_17 (.CK( clk ) , .Q( u1_L6_17 ) , .D( u1_R5_17 ) );
  DFF_X1 u1_L6_reg_18 (.CK( clk ) , .Q( u1_L6_18 ) , .D( u1_R5_18 ) );
  DFF_X1 u1_L6_reg_19 (.CK( clk ) , .Q( u1_L6_19 ) , .D( u1_R5_19 ) );
  DFF_X1 u1_L6_reg_2 (.CK( clk ) , .Q( u1_L6_2 ) , .D( u1_R5_2 ) );
  DFF_X1 u1_L6_reg_20 (.CK( clk ) , .Q( u1_L6_20 ) , .D( u1_R5_20 ) );
  DFF_X1 u1_L6_reg_21 (.CK( clk ) , .Q( u1_L6_21 ) , .D( u1_R5_21 ) );
  DFF_X1 u1_L6_reg_22 (.CK( clk ) , .Q( u1_L6_22 ) , .D( u1_R5_22 ) );
  DFF_X1 u1_L6_reg_23 (.CK( clk ) , .Q( u1_L6_23 ) , .D( u1_R5_23 ) );
  DFF_X1 u1_L6_reg_24 (.CK( clk ) , .Q( u1_L6_24 ) , .D( u1_R5_24 ) );
  DFF_X1 u1_L6_reg_25 (.CK( clk ) , .Q( u1_L6_25 ) , .D( u1_R5_25 ) );
  DFF_X1 u1_L6_reg_26 (.CK( clk ) , .Q( u1_L6_26 ) , .D( u1_R5_26 ) );
  DFF_X1 u1_L6_reg_27 (.CK( clk ) , .Q( u1_L6_27 ) , .D( u1_R5_27 ) );
  DFF_X1 u1_L6_reg_28 (.CK( clk ) , .Q( u1_L6_28 ) , .D( u1_R5_28 ) );
  DFF_X1 u1_L6_reg_29 (.CK( clk ) , .Q( u1_L6_29 ) , .D( u1_R5_29 ) );
  DFF_X1 u1_L6_reg_3 (.CK( clk ) , .Q( u1_L6_3 ) , .D( u1_R5_3 ) );
  DFF_X1 u1_L6_reg_30 (.CK( clk ) , .Q( u1_L6_30 ) , .D( u1_R5_30 ) );
  DFF_X1 u1_L6_reg_31 (.CK( clk ) , .Q( u1_L6_31 ) , .D( u1_R5_31 ) );
  DFF_X1 u1_L6_reg_32 (.CK( clk ) , .Q( u1_L6_32 ) , .D( u1_R5_32 ) );
  DFF_X1 u1_L6_reg_4 (.CK( clk ) , .Q( u1_L6_4 ) , .D( u1_R5_4 ) );
  DFF_X1 u1_L6_reg_5 (.CK( clk ) , .Q( u1_L6_5 ) , .D( u1_R5_5 ) );
  DFF_X1 u1_L6_reg_6 (.CK( clk ) , .Q( u1_L6_6 ) , .D( u1_R5_6 ) );
  DFF_X1 u1_L6_reg_7 (.CK( clk ) , .Q( u1_L6_7 ) , .D( u1_R5_7 ) );
  DFF_X1 u1_L6_reg_8 (.CK( clk ) , .Q( u1_L6_8 ) , .D( u1_R5_8 ) );
  DFF_X1 u1_L6_reg_9 (.CK( clk ) , .Q( u1_L6_9 ) , .D( u1_R5_9 ) );
  DFF_X1 u1_L7_reg_1 (.CK( clk ) , .Q( u1_L7_1 ) , .D( u1_R6_1 ) );
  DFF_X1 u1_L7_reg_10 (.CK( clk ) , .Q( u1_L7_10 ) , .D( u1_R6_10 ) );
  DFF_X1 u1_L7_reg_11 (.CK( clk ) , .Q( u1_L7_11 ) , .D( u1_R6_11 ) );
  DFF_X1 u1_L7_reg_12 (.CK( clk ) , .Q( u1_L7_12 ) , .D( u1_R6_12 ) );
  DFF_X1 u1_L7_reg_13 (.CK( clk ) , .Q( u1_L7_13 ) , .D( u1_R6_13 ) );
  DFF_X1 u1_L7_reg_14 (.CK( clk ) , .Q( u1_L7_14 ) , .D( u1_R6_14 ) );
  DFF_X1 u1_L7_reg_15 (.CK( clk ) , .Q( u1_L7_15 ) , .D( u1_R6_15 ) );
  DFF_X1 u1_L7_reg_16 (.CK( clk ) , .Q( u1_L7_16 ) , .D( u1_R6_16 ) );
  DFF_X1 u1_L7_reg_17 (.CK( clk ) , .Q( u1_L7_17 ) , .D( u1_R6_17 ) );
  DFF_X1 u1_L7_reg_18 (.CK( clk ) , .Q( u1_L7_18 ) , .D( u1_R6_18 ) );
  DFF_X1 u1_L7_reg_19 (.CK( clk ) , .Q( u1_L7_19 ) , .D( u1_R6_19 ) );
  DFF_X1 u1_L7_reg_2 (.CK( clk ) , .Q( u1_L7_2 ) , .D( u1_R6_2 ) );
  DFF_X1 u1_L7_reg_20 (.CK( clk ) , .Q( u1_L7_20 ) , .D( u1_R6_20 ) );
  DFF_X1 u1_L7_reg_21 (.CK( clk ) , .Q( u1_L7_21 ) , .D( u1_R6_21 ) );
  DFF_X1 u1_L7_reg_22 (.CK( clk ) , .Q( u1_L7_22 ) , .D( u1_R6_22 ) );
  DFF_X1 u1_L7_reg_23 (.CK( clk ) , .Q( u1_L7_23 ) , .D( u1_R6_23 ) );
  DFF_X1 u1_L7_reg_24 (.CK( clk ) , .Q( u1_L7_24 ) , .D( u1_R6_24 ) );
  DFF_X1 u1_L7_reg_25 (.CK( clk ) , .Q( u1_L7_25 ) , .D( u1_R6_25 ) );
  DFF_X1 u1_L7_reg_26 (.CK( clk ) , .Q( u1_L7_26 ) , .D( u1_R6_26 ) );
  DFF_X1 u1_L7_reg_27 (.CK( clk ) , .Q( u1_L7_27 ) , .D( u1_R6_27 ) );
  DFF_X1 u1_L7_reg_28 (.CK( clk ) , .Q( u1_L7_28 ) , .D( u1_R6_28 ) );
  DFF_X1 u1_L7_reg_29 (.CK( clk ) , .Q( u1_L7_29 ) , .D( u1_R6_29 ) );
  DFF_X1 u1_L7_reg_3 (.CK( clk ) , .Q( u1_L7_3 ) , .D( u1_R6_3 ) );
  DFF_X1 u1_L7_reg_30 (.CK( clk ) , .Q( u1_L7_30 ) , .D( u1_R6_30 ) );
  DFF_X1 u1_L7_reg_31 (.CK( clk ) , .Q( u1_L7_31 ) , .D( u1_R6_31 ) );
  DFF_X1 u1_L7_reg_32 (.CK( clk ) , .Q( u1_L7_32 ) , .D( u1_R6_32 ) );
  DFF_X1 u1_L7_reg_4 (.CK( clk ) , .Q( u1_L7_4 ) , .D( u1_R6_4 ) );
  DFF_X1 u1_L7_reg_5 (.CK( clk ) , .Q( u1_L7_5 ) , .D( u1_R6_5 ) );
  DFF_X1 u1_L7_reg_6 (.CK( clk ) , .Q( u1_L7_6 ) , .D( u1_R6_6 ) );
  DFF_X1 u1_L7_reg_7 (.CK( clk ) , .Q( u1_L7_7 ) , .D( u1_R6_7 ) );
  DFF_X1 u1_L7_reg_8 (.CK( clk ) , .Q( u1_L7_8 ) , .D( u1_R6_8 ) );
  DFF_X1 u1_L7_reg_9 (.CK( clk ) , .Q( u1_L7_9 ) , .D( u1_R6_9 ) );
  DFF_X1 u1_L8_reg_1 (.CK( clk ) , .Q( u1_L8_1 ) , .D( u1_R7_1 ) );
  DFF_X1 u1_L8_reg_10 (.CK( clk ) , .Q( u1_L8_10 ) , .D( u1_R7_10 ) );
  DFF_X1 u1_L8_reg_11 (.CK( clk ) , .Q( u1_L8_11 ) , .D( u1_R7_11 ) );
  DFF_X1 u1_L8_reg_12 (.CK( clk ) , .Q( u1_L8_12 ) , .D( u1_R7_12 ) );
  DFF_X1 u1_L8_reg_13 (.CK( clk ) , .Q( u1_L8_13 ) , .D( u1_R7_13 ) );
  DFF_X1 u1_L8_reg_14 (.CK( clk ) , .Q( u1_L8_14 ) , .D( u1_R7_14 ) );
  DFF_X1 u1_L8_reg_15 (.CK( clk ) , .Q( u1_L8_15 ) , .D( u1_R7_15 ) );
  DFF_X1 u1_L8_reg_16 (.CK( clk ) , .Q( u1_L8_16 ) , .D( u1_R7_16 ) );
  DFF_X1 u1_L8_reg_17 (.CK( clk ) , .Q( u1_L8_17 ) , .D( u1_R7_17 ) );
  DFF_X1 u1_L8_reg_18 (.CK( clk ) , .Q( u1_L8_18 ) , .D( u1_R7_18 ) );
  DFF_X1 u1_L8_reg_19 (.CK( clk ) , .Q( u1_L8_19 ) , .D( u1_R7_19 ) );
  DFF_X1 u1_L8_reg_2 (.CK( clk ) , .Q( u1_L8_2 ) , .D( u1_R7_2 ) );
  DFF_X1 u1_L8_reg_20 (.CK( clk ) , .Q( u1_L8_20 ) , .D( u1_R7_20 ) );
  DFF_X1 u1_L8_reg_21 (.CK( clk ) , .Q( u1_L8_21 ) , .D( u1_R7_21 ) );
  DFF_X1 u1_L8_reg_22 (.CK( clk ) , .Q( u1_L8_22 ) , .D( u1_R7_22 ) );
  DFF_X1 u1_L8_reg_23 (.CK( clk ) , .Q( u1_L8_23 ) , .D( u1_R7_23 ) );
  DFF_X1 u1_L8_reg_24 (.CK( clk ) , .Q( u1_L8_24 ) , .D( u1_R7_24 ) );
  DFF_X1 u1_L8_reg_25 (.CK( clk ) , .Q( u1_L8_25 ) , .D( u1_R7_25 ) );
  DFF_X1 u1_L8_reg_26 (.CK( clk ) , .Q( u1_L8_26 ) , .D( u1_R7_26 ) );
  DFF_X1 u1_L8_reg_27 (.CK( clk ) , .Q( u1_L8_27 ) , .D( u1_R7_27 ) );
  DFF_X1 u1_L8_reg_28 (.CK( clk ) , .Q( u1_L8_28 ) , .D( u1_R7_28 ) );
  DFF_X1 u1_L8_reg_29 (.CK( clk ) , .Q( u1_L8_29 ) , .D( u1_R7_29 ) );
  DFF_X1 u1_L8_reg_3 (.CK( clk ) , .Q( u1_L8_3 ) , .D( u1_R7_3 ) );
  DFF_X1 u1_L8_reg_30 (.CK( clk ) , .Q( u1_L8_30 ) , .D( u1_R7_30 ) );
  DFF_X1 u1_L8_reg_31 (.CK( clk ) , .Q( u1_L8_31 ) , .D( u1_R7_31 ) );
  DFF_X1 u1_L8_reg_32 (.CK( clk ) , .Q( u1_L8_32 ) , .D( u1_R7_32 ) );
  DFF_X1 u1_L8_reg_4 (.CK( clk ) , .Q( u1_L8_4 ) , .D( u1_R7_4 ) );
  DFF_X1 u1_L8_reg_5 (.CK( clk ) , .Q( u1_L8_5 ) , .D( u1_R7_5 ) );
  DFF_X1 u1_L8_reg_6 (.CK( clk ) , .Q( u1_L8_6 ) , .D( u1_R7_6 ) );
  DFF_X1 u1_L8_reg_7 (.CK( clk ) , .Q( u1_L8_7 ) , .D( u1_R7_7 ) );
  DFF_X1 u1_L8_reg_8 (.CK( clk ) , .Q( u1_L8_8 ) , .D( u1_R7_8 ) );
  DFF_X1 u1_L8_reg_9 (.CK( clk ) , .Q( u1_L8_9 ) , .D( u1_R7_9 ) );
  DFF_X1 u1_L9_reg_1 (.CK( clk ) , .Q( u1_L9_1 ) , .D( u1_R8_1 ) );
  DFF_X1 u1_L9_reg_10 (.CK( clk ) , .Q( u1_L9_10 ) , .D( u1_R8_10 ) );
  DFF_X1 u1_L9_reg_11 (.CK( clk ) , .Q( u1_L9_11 ) , .D( u1_R8_11 ) );
  DFF_X1 u1_L9_reg_12 (.CK( clk ) , .Q( u1_L9_12 ) , .D( u1_R8_12 ) );
  DFF_X1 u1_L9_reg_13 (.CK( clk ) , .Q( u1_L9_13 ) , .D( u1_R8_13 ) );
  DFF_X1 u1_L9_reg_14 (.CK( clk ) , .Q( u1_L9_14 ) , .D( u1_R8_14 ) );
  DFF_X1 u1_L9_reg_15 (.CK( clk ) , .Q( u1_L9_15 ) , .D( u1_R8_15 ) );
  DFF_X1 u1_L9_reg_16 (.CK( clk ) , .Q( u1_L9_16 ) , .D( u1_R8_16 ) );
  DFF_X1 u1_L9_reg_17 (.CK( clk ) , .Q( u1_L9_17 ) , .D( u1_R8_17 ) );
  DFF_X1 u1_L9_reg_18 (.CK( clk ) , .Q( u1_L9_18 ) , .D( u1_R8_18 ) );
  DFF_X1 u1_L9_reg_19 (.CK( clk ) , .Q( u1_L9_19 ) , .D( u1_R8_19 ) );
  DFF_X1 u1_L9_reg_2 (.CK( clk ) , .Q( u1_L9_2 ) , .D( u1_R8_2 ) );
  DFF_X1 u1_L9_reg_20 (.CK( clk ) , .Q( u1_L9_20 ) , .D( u1_R8_20 ) );
  DFF_X1 u1_L9_reg_21 (.CK( clk ) , .Q( u1_L9_21 ) , .D( u1_R8_21 ) );
  DFF_X1 u1_L9_reg_22 (.CK( clk ) , .Q( u1_L9_22 ) , .D( u1_R8_22 ) );
  DFF_X1 u1_L9_reg_23 (.CK( clk ) , .Q( u1_L9_23 ) , .D( u1_R8_23 ) );
  DFF_X1 u1_L9_reg_24 (.CK( clk ) , .Q( u1_L9_24 ) , .D( u1_R8_24 ) );
  DFF_X1 u1_L9_reg_25 (.CK( clk ) , .Q( u1_L9_25 ) , .D( u1_R8_25 ) );
  DFF_X1 u1_L9_reg_26 (.CK( clk ) , .Q( u1_L9_26 ) , .D( u1_R8_26 ) );
  DFF_X1 u1_L9_reg_27 (.CK( clk ) , .Q( u1_L9_27 ) , .D( u1_R8_27 ) );
  DFF_X1 u1_L9_reg_28 (.CK( clk ) , .Q( u1_L9_28 ) , .D( u1_R8_28 ) );
  DFF_X1 u1_L9_reg_29 (.CK( clk ) , .Q( u1_L9_29 ) , .D( u1_R8_29 ) );
  DFF_X1 u1_L9_reg_3 (.CK( clk ) , .Q( u1_L9_3 ) , .D( u1_R8_3 ) );
  DFF_X1 u1_L9_reg_30 (.CK( clk ) , .Q( u1_L9_30 ) , .D( u1_R8_30 ) );
  DFF_X1 u1_L9_reg_31 (.CK( clk ) , .Q( u1_L9_31 ) , .D( u1_R8_31 ) );
  DFF_X1 u1_L9_reg_32 (.CK( clk ) , .Q( u1_L9_32 ) , .D( u1_R8_32 ) );
  DFF_X1 u1_L9_reg_4 (.CK( clk ) , .Q( u1_L9_4 ) , .D( u1_R8_4 ) );
  DFF_X1 u1_L9_reg_5 (.CK( clk ) , .Q( u1_L9_5 ) , .D( u1_R8_5 ) );
  DFF_X1 u1_L9_reg_6 (.CK( clk ) , .Q( u1_L9_6 ) , .D( u1_R8_6 ) );
  DFF_X1 u1_L9_reg_7 (.CK( clk ) , .Q( u1_L9_7 ) , .D( u1_R8_7 ) );
  DFF_X1 u1_L9_reg_8 (.CK( clk ) , .Q( u1_L9_8 ) , .D( u1_R8_8 ) );
  DFF_X1 u1_L9_reg_9 (.CK( clk ) , .Q( u1_L9_9 ) , .D( u1_R8_9 ) );
  DFF_X1 u1_R0_reg_1 (.CK( clk ) , .D( u1_N0 ) , .Q( u1_R0_1 ) );
  DFF_X1 u1_R0_reg_10 (.CK( clk ) , .D( u1_N9 ) , .Q( u1_R0_10 ) );
  DFF_X1 u1_R0_reg_11 (.CK( clk ) , .D( u1_N10 ) , .Q( u1_R0_11 ) );
  DFF_X1 u1_R0_reg_12 (.CK( clk ) , .D( u1_N11 ) , .Q( u1_R0_12 ) );
  DFF_X1 u1_R0_reg_13 (.CK( clk ) , .D( u1_N12 ) , .Q( u1_R0_13 ) );
  DFF_X1 u1_R0_reg_14 (.CK( clk ) , .D( u1_N13 ) , .Q( u1_R0_14 ) );
  DFF_X1 u1_R0_reg_15 (.CK( clk ) , .D( u1_N14 ) , .Q( u1_R0_15 ) );
  DFF_X1 u1_R0_reg_16 (.CK( clk ) , .D( u1_N15 ) , .Q( u1_R0_16 ) );
  DFF_X1 u1_R0_reg_17 (.CK( clk ) , .D( u1_N16 ) , .Q( u1_R0_17 ) );
  DFF_X1 u1_R0_reg_18 (.CK( clk ) , .D( u1_N17 ) , .Q( u1_R0_18 ) );
  DFF_X1 u1_R0_reg_19 (.CK( clk ) , .D( u1_N18 ) , .Q( u1_R0_19 ) );
  DFF_X1 u1_R0_reg_2 (.CK( clk ) , .D( u1_N1 ) , .Q( u1_R0_2 ) );
  DFF_X1 u1_R0_reg_20 (.CK( clk ) , .D( u1_N19 ) , .Q( u1_R0_20 ) );
  DFF_X1 u1_R0_reg_21 (.CK( clk ) , .D( u1_N20 ) , .Q( u1_R0_21 ) );
  DFF_X1 u1_R0_reg_22 (.CK( clk ) , .D( u1_N21 ) , .Q( u1_R0_22 ) );
  DFF_X1 u1_R0_reg_23 (.CK( clk ) , .D( u1_N22 ) , .Q( u1_R0_23 ) );
  DFF_X1 u1_R0_reg_24 (.CK( clk ) , .D( u1_N23 ) , .Q( u1_R0_24 ) );
  DFF_X1 u1_R0_reg_25 (.CK( clk ) , .D( u1_N24 ) , .Q( u1_R0_25 ) );
  DFF_X1 u1_R0_reg_26 (.CK( clk ) , .D( u1_N25 ) , .Q( u1_R0_26 ) );
  DFF_X1 u1_R0_reg_27 (.CK( clk ) , .D( u1_N26 ) , .Q( u1_R0_27 ) );
  DFF_X1 u1_R0_reg_28 (.CK( clk ) , .D( u1_N27 ) , .Q( u1_R0_28 ) );
  DFF_X1 u1_R0_reg_29 (.CK( clk ) , .D( u1_N28 ) , .Q( u1_R0_29 ) );
  DFF_X1 u1_R0_reg_3 (.CK( clk ) , .D( u1_N2 ) , .Q( u1_R0_3 ) );
  DFF_X1 u1_R0_reg_30 (.CK( clk ) , .D( u1_N29 ) , .Q( u1_R0_30 ) );
  DFF_X1 u1_R0_reg_31 (.CK( clk ) , .D( u1_N30 ) , .Q( u1_R0_31 ) );
  DFF_X1 u1_R0_reg_32 (.CK( clk ) , .D( u1_N31 ) , .Q( u1_R0_32 ) );
  DFF_X1 u1_R0_reg_4 (.CK( clk ) , .D( u1_N3 ) , .Q( u1_R0_4 ) );
  DFF_X1 u1_R0_reg_5 (.CK( clk ) , .D( u1_N4 ) , .Q( u1_R0_5 ) );
  DFF_X1 u1_R0_reg_6 (.CK( clk ) , .D( u1_N5 ) , .Q( u1_R0_6 ) );
  DFF_X1 u1_R0_reg_7 (.CK( clk ) , .D( u1_N6 ) , .Q( u1_R0_7 ) );
  DFF_X1 u1_R0_reg_8 (.CK( clk ) , .D( u1_N7 ) , .Q( u1_R0_8 ) );
  DFF_X1 u1_R0_reg_9 (.CK( clk ) , .D( u1_N8 ) , .Q( u1_R0_9 ) );
  DFF_X1 u1_R10_reg_1 (.CK( clk ) , .D( u1_N320 ) , .Q( u1_R10_1 ) );
  DFF_X1 u1_R10_reg_10 (.CK( clk ) , .D( u1_N329 ) , .Q( u1_R10_10 ) );
  DFF_X1 u1_R10_reg_11 (.CK( clk ) , .D( u1_N330 ) , .Q( u1_R10_11 ) );
  DFF_X1 u1_R10_reg_12 (.CK( clk ) , .D( u1_N331 ) , .Q( u1_R10_12 ) );
  DFF_X1 u1_R10_reg_13 (.CK( clk ) , .D( u1_N332 ) , .Q( u1_R10_13 ) );
  DFF_X1 u1_R10_reg_14 (.CK( clk ) , .D( u1_N333 ) , .Q( u1_R10_14 ) );
  DFF_X1 u1_R10_reg_15 (.CK( clk ) , .D( u1_N334 ) , .Q( u1_R10_15 ) );
  DFF_X1 u1_R10_reg_16 (.CK( clk ) , .D( u1_N335 ) , .Q( u1_R10_16 ) );
  DFF_X1 u1_R10_reg_17 (.CK( clk ) , .D( u1_N336 ) , .Q( u1_R10_17 ) );
  DFF_X1 u1_R10_reg_18 (.CK( clk ) , .D( u1_N337 ) , .Q( u1_R10_18 ) );
  DFF_X1 u1_R10_reg_19 (.CK( clk ) , .D( u1_N338 ) , .Q( u1_R10_19 ) );
  DFF_X1 u1_R10_reg_2 (.CK( clk ) , .D( u1_N321 ) , .Q( u1_R10_2 ) );
  DFF_X1 u1_R10_reg_20 (.CK( clk ) , .D( u1_N339 ) , .Q( u1_R10_20 ) );
  DFF_X1 u1_R10_reg_21 (.CK( clk ) , .D( u1_N340 ) , .Q( u1_R10_21 ) );
  DFF_X1 u1_R10_reg_22 (.CK( clk ) , .D( u1_N341 ) , .Q( u1_R10_22 ) );
  DFF_X1 u1_R10_reg_23 (.CK( clk ) , .D( u1_N342 ) , .Q( u1_R10_23 ) );
  DFF_X1 u1_R10_reg_24 (.CK( clk ) , .D( u1_N343 ) , .Q( u1_R10_24 ) );
  DFF_X1 u1_R10_reg_25 (.CK( clk ) , .D( u1_N344 ) , .Q( u1_R10_25 ) );
  DFF_X1 u1_R10_reg_26 (.CK( clk ) , .D( u1_N345 ) , .Q( u1_R10_26 ) );
  DFF_X1 u1_R10_reg_27 (.CK( clk ) , .D( u1_N346 ) , .Q( u1_R10_27 ) );
  DFF_X1 u1_R10_reg_28 (.CK( clk ) , .D( u1_N347 ) , .Q( u1_R10_28 ) );
  DFF_X1 u1_R10_reg_29 (.CK( clk ) , .D( u1_N348 ) , .Q( u1_R10_29 ) );
  DFF_X1 u1_R10_reg_3 (.CK( clk ) , .D( u1_N322 ) , .Q( u1_R10_3 ) );
  DFF_X1 u1_R10_reg_30 (.CK( clk ) , .D( u1_N349 ) , .Q( u1_R10_30 ) );
  DFF_X1 u1_R10_reg_31 (.CK( clk ) , .D( u1_N350 ) , .Q( u1_R10_31 ) );
  DFF_X1 u1_R10_reg_32 (.CK( clk ) , .D( u1_N351 ) , .Q( u1_R10_32 ) );
  DFF_X1 u1_R10_reg_4 (.CK( clk ) , .D( u1_N323 ) , .Q( u1_R10_4 ) );
  DFF_X1 u1_R10_reg_5 (.CK( clk ) , .D( u1_N324 ) , .Q( u1_R10_5 ) );
  DFF_X1 u1_R10_reg_6 (.CK( clk ) , .D( u1_N325 ) , .Q( u1_R10_6 ) );
  DFF_X1 u1_R10_reg_7 (.CK( clk ) , .D( u1_N326 ) , .Q( u1_R10_7 ) );
  DFF_X1 u1_R10_reg_8 (.CK( clk ) , .D( u1_N327 ) , .Q( u1_R10_8 ) );
  DFF_X1 u1_R10_reg_9 (.CK( clk ) , .D( u1_N328 ) , .Q( u1_R10_9 ) );
  DFF_X1 u1_R11_reg_1 (.CK( clk ) , .D( u1_N352 ) , .Q( u1_R11_1 ) );
  DFF_X1 u1_R11_reg_10 (.CK( clk ) , .D( u1_N361 ) , .Q( u1_R11_10 ) );
  DFF_X1 u1_R11_reg_11 (.CK( clk ) , .D( u1_N362 ) , .Q( u1_R11_11 ) );
  DFF_X1 u1_R11_reg_12 (.CK( clk ) , .D( u1_N363 ) , .Q( u1_R11_12 ) );
  DFF_X1 u1_R11_reg_13 (.CK( clk ) , .D( u1_N364 ) , .Q( u1_R11_13 ) );
  DFF_X1 u1_R11_reg_14 (.CK( clk ) , .D( u1_N365 ) , .Q( u1_R11_14 ) );
  DFF_X1 u1_R11_reg_15 (.CK( clk ) , .D( u1_N366 ) , .Q( u1_R11_15 ) );
  DFF_X1 u1_R11_reg_16 (.CK( clk ) , .D( u1_N367 ) , .Q( u1_R11_16 ) );
  DFF_X1 u1_R11_reg_17 (.CK( clk ) , .D( u1_N368 ) , .Q( u1_R11_17 ) );
  DFF_X1 u1_R11_reg_18 (.CK( clk ) , .D( u1_N369 ) , .Q( u1_R11_18 ) );
  DFF_X1 u1_R11_reg_19 (.CK( clk ) , .D( u1_N370 ) , .Q( u1_R11_19 ) );
  DFF_X1 u1_R11_reg_2 (.CK( clk ) , .D( u1_N353 ) , .Q( u1_R11_2 ) );
  DFF_X1 u1_R11_reg_20 (.CK( clk ) , .D( u1_N371 ) , .Q( u1_R11_20 ) );
  DFF_X1 u1_R11_reg_21 (.CK( clk ) , .D( u1_N372 ) , .Q( u1_R11_21 ) );
  DFF_X1 u1_R11_reg_22 (.CK( clk ) , .D( u1_N373 ) , .Q( u1_R11_22 ) );
  DFF_X1 u1_R11_reg_23 (.CK( clk ) , .D( u1_N374 ) , .Q( u1_R11_23 ) );
  DFF_X1 u1_R11_reg_24 (.CK( clk ) , .D( u1_N375 ) , .Q( u1_R11_24 ) );
  DFF_X1 u1_R11_reg_25 (.CK( clk ) , .D( u1_N376 ) , .Q( u1_R11_25 ) );
  DFF_X1 u1_R11_reg_26 (.CK( clk ) , .D( u1_N377 ) , .Q( u1_R11_26 ) );
  DFF_X1 u1_R11_reg_27 (.CK( clk ) , .D( u1_N378 ) , .Q( u1_R11_27 ) );
  DFF_X1 u1_R11_reg_28 (.CK( clk ) , .D( u1_N379 ) , .Q( u1_R11_28 ) );
  DFF_X1 u1_R11_reg_29 (.CK( clk ) , .D( u1_N380 ) , .Q( u1_R11_29 ) );
  DFF_X1 u1_R11_reg_3 (.CK( clk ) , .D( u1_N354 ) , .Q( u1_R11_3 ) );
  DFF_X1 u1_R11_reg_30 (.CK( clk ) , .D( u1_N381 ) , .Q( u1_R11_30 ) );
  DFF_X1 u1_R11_reg_31 (.CK( clk ) , .D( u1_N382 ) , .Q( u1_R11_31 ) );
  DFF_X1 u1_R11_reg_32 (.CK( clk ) , .D( u1_N383 ) , .Q( u1_R11_32 ) );
  DFF_X1 u1_R11_reg_4 (.CK( clk ) , .D( u1_N355 ) , .Q( u1_R11_4 ) );
  DFF_X1 u1_R11_reg_5 (.CK( clk ) , .D( u1_N356 ) , .Q( u1_R11_5 ) );
  DFF_X1 u1_R11_reg_6 (.CK( clk ) , .D( u1_N357 ) , .Q( u1_R11_6 ) );
  DFF_X1 u1_R11_reg_7 (.CK( clk ) , .D( u1_N358 ) , .Q( u1_R11_7 ) );
  DFF_X1 u1_R11_reg_8 (.CK( clk ) , .D( u1_N359 ) , .Q( u1_R11_8 ) );
  DFF_X1 u1_R11_reg_9 (.CK( clk ) , .D( u1_N360 ) , .Q( u1_R11_9 ) );
  DFF_X1 u1_R12_reg_1 (.CK( clk ) , .D( u1_N384 ) , .Q( u1_R12_1 ) );
  DFF_X1 u1_R12_reg_10 (.CK( clk ) , .D( u1_N393 ) , .Q( u1_R12_10 ) );
  DFF_X1 u1_R12_reg_11 (.CK( clk ) , .D( u1_N394 ) , .Q( u1_R12_11 ) );
  DFF_X1 u1_R12_reg_12 (.CK( clk ) , .D( u1_N395 ) , .Q( u1_R12_12 ) );
  DFF_X1 u1_R12_reg_13 (.CK( clk ) , .D( u1_N396 ) , .Q( u1_R12_13 ) );
  DFF_X1 u1_R12_reg_14 (.CK( clk ) , .D( u1_N397 ) , .Q( u1_R12_14 ) );
  DFF_X1 u1_R12_reg_15 (.CK( clk ) , .D( u1_N398 ) , .Q( u1_R12_15 ) );
  DFF_X1 u1_R12_reg_16 (.CK( clk ) , .D( u1_N399 ) , .Q( u1_R12_16 ) );
  DFF_X1 u1_R12_reg_17 (.CK( clk ) , .D( u1_N400 ) , .Q( u1_R12_17 ) );
  DFF_X1 u1_R12_reg_18 (.CK( clk ) , .D( u1_N401 ) , .Q( u1_R12_18 ) );
  DFF_X1 u1_R12_reg_19 (.CK( clk ) , .D( u1_N402 ) , .Q( u1_R12_19 ) );
  DFF_X1 u1_R12_reg_2 (.CK( clk ) , .D( u1_N385 ) , .Q( u1_R12_2 ) );
  DFF_X1 u1_R12_reg_20 (.CK( clk ) , .D( u1_N403 ) , .Q( u1_R12_20 ) );
  DFF_X1 u1_R12_reg_21 (.CK( clk ) , .D( u1_N404 ) , .Q( u1_R12_21 ) );
  DFF_X1 u1_R12_reg_22 (.CK( clk ) , .D( u1_N405 ) , .Q( u1_R12_22 ) );
  DFF_X1 u1_R12_reg_23 (.CK( clk ) , .D( u1_N406 ) , .Q( u1_R12_23 ) );
  DFF_X1 u1_R12_reg_24 (.CK( clk ) , .D( u1_N407 ) , .Q( u1_R12_24 ) );
  DFF_X1 u1_R12_reg_25 (.CK( clk ) , .D( u1_N408 ) , .Q( u1_R12_25 ) );
  DFF_X1 u1_R12_reg_26 (.CK( clk ) , .D( u1_N409 ) , .Q( u1_R12_26 ) );
  DFF_X1 u1_R12_reg_27 (.CK( clk ) , .D( u1_N410 ) , .Q( u1_R12_27 ) );
  DFF_X1 u1_R12_reg_28 (.CK( clk ) , .D( u1_N411 ) , .Q( u1_R12_28 ) );
  DFF_X1 u1_R12_reg_29 (.CK( clk ) , .D( u1_N412 ) , .Q( u1_R12_29 ) );
  DFF_X1 u1_R12_reg_3 (.CK( clk ) , .D( u1_N386 ) , .Q( u1_R12_3 ) );
  DFF_X1 u1_R12_reg_30 (.CK( clk ) , .D( u1_N413 ) , .Q( u1_R12_30 ) );
  DFF_X1 u1_R12_reg_31 (.CK( clk ) , .D( u1_N414 ) , .Q( u1_R12_31 ) );
  DFF_X1 u1_R12_reg_32 (.CK( clk ) , .D( u1_N415 ) , .Q( u1_R12_32 ) );
  DFF_X1 u1_R12_reg_4 (.CK( clk ) , .D( u1_N387 ) , .Q( u1_R12_4 ) );
  DFF_X1 u1_R12_reg_5 (.CK( clk ) , .D( u1_N388 ) , .Q( u1_R12_5 ) );
  DFF_X1 u1_R12_reg_6 (.CK( clk ) , .D( u1_N389 ) , .Q( u1_R12_6 ) );
  DFF_X1 u1_R12_reg_7 (.CK( clk ) , .D( u1_N390 ) , .Q( u1_R12_7 ) );
  DFF_X1 u1_R12_reg_8 (.CK( clk ) , .D( u1_N391 ) , .Q( u1_R12_8 ) );
  DFF_X1 u1_R12_reg_9 (.CK( clk ) , .D( u1_N392 ) , .Q( u1_R12_9 ) );
  DFF_X1 u1_R13_reg_1 (.CK( clk ) , .D( u1_N416 ) , .Q( u1_R13_1 ) );
  DFF_X1 u1_R13_reg_10 (.CK( clk ) , .D( u1_N425 ) , .Q( u1_R13_10 ) );
  DFF_X1 u1_R13_reg_11 (.CK( clk ) , .D( u1_N426 ) , .Q( u1_R13_11 ) );
  DFF_X1 u1_R13_reg_12 (.CK( clk ) , .D( u1_N427 ) , .Q( u1_R13_12 ) );
  DFF_X1 u1_R13_reg_13 (.CK( clk ) , .D( u1_N428 ) , .Q( u1_R13_13 ) );
  DFF_X1 u1_R13_reg_14 (.CK( clk ) , .D( u1_N429 ) , .Q( u1_R13_14 ) );
  DFF_X1 u1_R13_reg_15 (.CK( clk ) , .D( u1_N430 ) , .Q( u1_R13_15 ) );
  DFF_X1 u1_R13_reg_16 (.CK( clk ) , .D( u1_N431 ) , .Q( u1_R13_16 ) );
  DFF_X1 u1_R13_reg_17 (.CK( clk ) , .D( u1_N432 ) , .Q( u1_R13_17 ) );
  DFF_X1 u1_R13_reg_18 (.CK( clk ) , .D( u1_N433 ) , .Q( u1_R13_18 ) );
  DFF_X1 u1_R13_reg_19 (.CK( clk ) , .D( u1_N434 ) , .Q( u1_R13_19 ) );
  DFF_X1 u1_R13_reg_2 (.CK( clk ) , .D( u1_N417 ) , .Q( u1_R13_2 ) );
  DFF_X1 u1_R13_reg_20 (.CK( clk ) , .D( u1_N435 ) , .Q( u1_R13_20 ) );
  DFF_X1 u1_R13_reg_21 (.CK( clk ) , .D( u1_N436 ) , .Q( u1_R13_21 ) );
  DFF_X1 u1_R13_reg_22 (.CK( clk ) , .D( u1_N437 ) , .Q( u1_R13_22 ) );
  DFF_X1 u1_R13_reg_23 (.CK( clk ) , .D( u1_N438 ) , .Q( u1_R13_23 ) );
  DFF_X1 u1_R13_reg_24 (.CK( clk ) , .D( u1_N439 ) , .Q( u1_R13_24 ) );
  DFF_X1 u1_R13_reg_25 (.CK( clk ) , .D( u1_N440 ) , .Q( u1_R13_25 ) );
  DFF_X1 u1_R13_reg_26 (.CK( clk ) , .D( u1_N441 ) , .Q( u1_R13_26 ) );
  DFF_X1 u1_R13_reg_27 (.CK( clk ) , .D( u1_N442 ) , .Q( u1_R13_27 ) );
  DFF_X1 u1_R13_reg_28 (.CK( clk ) , .D( u1_N443 ) , .Q( u1_R13_28 ) );
  DFF_X1 u1_R13_reg_29 (.CK( clk ) , .D( u1_N444 ) , .Q( u1_R13_29 ) );
  DFF_X1 u1_R13_reg_3 (.CK( clk ) , .D( u1_N418 ) , .Q( u1_R13_3 ) );
  DFF_X1 u1_R13_reg_30 (.CK( clk ) , .D( u1_N445 ) , .Q( u1_R13_30 ) );
  DFF_X1 u1_R13_reg_31 (.CK( clk ) , .D( u1_N446 ) , .Q( u1_R13_31 ) );
  DFF_X1 u1_R13_reg_32 (.CK( clk ) , .D( u1_N447 ) , .Q( u1_R13_32 ) );
  DFF_X1 u1_R13_reg_4 (.CK( clk ) , .D( u1_N419 ) , .Q( u1_R13_4 ) );
  DFF_X1 u1_R13_reg_5 (.CK( clk ) , .D( u1_N420 ) , .Q( u1_R13_5 ) );
  DFF_X1 u1_R13_reg_6 (.CK( clk ) , .D( u1_N421 ) , .Q( u1_R13_6 ) );
  DFF_X1 u1_R13_reg_7 (.CK( clk ) , .D( u1_N422 ) , .Q( u1_R13_7 ) );
  DFF_X1 u1_R13_reg_8 (.CK( clk ) , .D( u1_N423 ) , .Q( u1_R13_8 ) );
  DFF_X1 u1_R13_reg_9 (.CK( clk ) , .D( u1_N424 ) , .Q( u1_R13_9 ) );
  DFF_X1 u1_R14_reg_1 (.CK( clk ) , .Q( u1_FP_33 ) , .D( u1_N448 ) );
  DFF_X1 u1_R14_reg_10 (.CK( clk ) , .Q( u1_FP_42 ) , .D( u1_N457 ) );
  DFF_X1 u1_R14_reg_11 (.CK( clk ) , .Q( u1_FP_43 ) , .D( u1_N458 ) );
  DFF_X1 u1_R14_reg_12 (.CK( clk ) , .Q( u1_FP_44 ) , .D( u1_N459 ) );
  DFF_X1 u1_R14_reg_13 (.CK( clk ) , .Q( u1_FP_45 ) , .D( u1_N460 ) );
  DFF_X1 u1_R14_reg_14 (.CK( clk ) , .Q( u1_FP_46 ) , .D( u1_N461 ) );
  DFF_X1 u1_R14_reg_15 (.CK( clk ) , .Q( u1_FP_47 ) , .D( u1_N462 ) );
  DFF_X1 u1_R14_reg_16 (.CK( clk ) , .Q( u1_FP_48 ) , .D( u1_N463 ) );
  DFF_X1 u1_R14_reg_17 (.CK( clk ) , .Q( u1_FP_49 ) , .D( u1_N464 ) );
  DFF_X1 u1_R14_reg_18 (.CK( clk ) , .Q( u1_FP_50 ) , .D( u1_N465 ) );
  DFF_X1 u1_R14_reg_19 (.CK( clk ) , .Q( u1_FP_51 ) , .D( u1_N466 ) );
  DFF_X1 u1_R14_reg_2 (.CK( clk ) , .Q( u1_FP_34 ) , .D( u1_N449 ) );
  DFF_X1 u1_R14_reg_20 (.CK( clk ) , .Q( u1_FP_52 ) , .D( u1_N467 ) );
  DFF_X1 u1_R14_reg_21 (.CK( clk ) , .Q( u1_FP_53 ) , .D( u1_N468 ) );
  DFF_X1 u1_R14_reg_22 (.CK( clk ) , .Q( u1_FP_54 ) , .D( u1_N469 ) );
  DFF_X1 u1_R14_reg_23 (.CK( clk ) , .Q( u1_FP_55 ) , .D( u1_N470 ) );
  DFF_X1 u1_R14_reg_24 (.CK( clk ) , .Q( u1_FP_56 ) , .D( u1_N471 ) );
  DFF_X1 u1_R14_reg_25 (.CK( clk ) , .Q( u1_FP_57 ) , .D( u1_N472 ) );
  DFF_X1 u1_R14_reg_26 (.CK( clk ) , .Q( u1_FP_58 ) , .D( u1_N473 ) );
  DFF_X1 u1_R14_reg_27 (.CK( clk ) , .Q( u1_FP_59 ) , .D( u1_N474 ) );
  DFF_X1 u1_R14_reg_28 (.CK( clk ) , .Q( u1_FP_60 ) , .D( u1_N475 ) );
  DFF_X1 u1_R14_reg_29 (.CK( clk ) , .Q( u1_FP_61 ) , .D( u1_N476 ) );
  DFF_X1 u1_R14_reg_3 (.CK( clk ) , .Q( u1_FP_35 ) , .D( u1_N450 ) );
  DFF_X1 u1_R14_reg_30 (.CK( clk ) , .Q( u1_FP_62 ) , .D( u1_N477 ) );
  DFF_X1 u1_R14_reg_31 (.CK( clk ) , .Q( u1_FP_63 ) , .D( u1_N478 ) );
  DFF_X1 u1_R14_reg_32 (.CK( clk ) , .Q( u1_FP_64 ) , .D( u1_N479 ) );
  DFF_X1 u1_R14_reg_4 (.CK( clk ) , .Q( u1_FP_36 ) , .D( u1_N451 ) );
  DFF_X1 u1_R14_reg_5 (.CK( clk ) , .Q( u1_FP_37 ) , .D( u1_N452 ) );
  DFF_X1 u1_R14_reg_6 (.CK( clk ) , .Q( u1_FP_38 ) , .D( u1_N453 ) );
  DFF_X1 u1_R14_reg_7 (.CK( clk ) , .Q( u1_FP_39 ) , .D( u1_N454 ) );
  DFF_X1 u1_R14_reg_8 (.CK( clk ) , .Q( u1_FP_40 ) , .D( u1_N455 ) );
  DFF_X1 u1_R14_reg_9 (.CK( clk ) , .Q( u1_FP_41 ) , .D( u1_N456 ) );
  DFF_X1 u1_R1_reg_1 (.CK( clk ) , .D( u1_N32 ) , .Q( u1_R1_1 ) );
  DFF_X1 u1_R1_reg_10 (.CK( clk ) , .D( u1_N41 ) , .Q( u1_R1_10 ) );
  DFF_X1 u1_R1_reg_11 (.CK( clk ) , .D( u1_N42 ) , .Q( u1_R1_11 ) );
  DFF_X1 u1_R1_reg_12 (.CK( clk ) , .D( u1_N43 ) , .Q( u1_R1_12 ) );
  DFF_X1 u1_R1_reg_13 (.CK( clk ) , .D( u1_N44 ) , .Q( u1_R1_13 ) );
  DFF_X1 u1_R1_reg_14 (.CK( clk ) , .D( u1_N45 ) , .Q( u1_R1_14 ) );
  DFF_X1 u1_R1_reg_15 (.CK( clk ) , .D( u1_N46 ) , .Q( u1_R1_15 ) );
  DFF_X1 u1_R1_reg_16 (.CK( clk ) , .D( u1_N47 ) , .Q( u1_R1_16 ) );
  DFF_X1 u1_R1_reg_17 (.CK( clk ) , .D( u1_N48 ) , .Q( u1_R1_17 ) );
  DFF_X1 u1_R1_reg_18 (.CK( clk ) , .D( u1_N49 ) , .Q( u1_R1_18 ) );
  DFF_X1 u1_R1_reg_19 (.CK( clk ) , .D( u1_N50 ) , .Q( u1_R1_19 ) );
  DFF_X1 u1_R1_reg_2 (.CK( clk ) , .D( u1_N33 ) , .Q( u1_R1_2 ) );
  DFF_X1 u1_R1_reg_20 (.CK( clk ) , .D( u1_N51 ) , .Q( u1_R1_20 ) );
  DFF_X1 u1_R1_reg_21 (.CK( clk ) , .D( u1_N52 ) , .Q( u1_R1_21 ) );
  DFF_X1 u1_R1_reg_22 (.CK( clk ) , .D( u1_N53 ) , .Q( u1_R1_22 ) );
  DFF_X1 u1_R1_reg_23 (.CK( clk ) , .D( u1_N54 ) , .Q( u1_R1_23 ) );
  DFF_X1 u1_R1_reg_24 (.CK( clk ) , .D( u1_N55 ) , .Q( u1_R1_24 ) );
  DFF_X1 u1_R1_reg_25 (.CK( clk ) , .D( u1_N56 ) , .Q( u1_R1_25 ) );
  DFF_X1 u1_R1_reg_26 (.CK( clk ) , .D( u1_N57 ) , .Q( u1_R1_26 ) );
  DFF_X1 u1_R1_reg_27 (.CK( clk ) , .D( u1_N58 ) , .Q( u1_R1_27 ) );
  DFF_X1 u1_R1_reg_28 (.CK( clk ) , .D( u1_N59 ) , .Q( u1_R1_28 ) );
  DFF_X1 u1_R1_reg_29 (.CK( clk ) , .D( u1_N60 ) , .Q( u1_R1_29 ) );
  DFF_X1 u1_R1_reg_3 (.CK( clk ) , .D( u1_N34 ) , .Q( u1_R1_3 ) );
  DFF_X1 u1_R1_reg_30 (.CK( clk ) , .D( u1_N61 ) , .Q( u1_R1_30 ) );
  DFF_X1 u1_R1_reg_31 (.CK( clk ) , .D( u1_N62 ) , .Q( u1_R1_31 ) );
  DFF_X1 u1_R1_reg_32 (.CK( clk ) , .D( u1_N63 ) , .Q( u1_R1_32 ) );
  DFF_X1 u1_R1_reg_4 (.CK( clk ) , .D( u1_N35 ) , .Q( u1_R1_4 ) );
  DFF_X1 u1_R1_reg_5 (.CK( clk ) , .D( u1_N36 ) , .Q( u1_R1_5 ) );
  DFF_X1 u1_R1_reg_6 (.CK( clk ) , .D( u1_N37 ) , .Q( u1_R1_6 ) );
  DFF_X1 u1_R1_reg_7 (.CK( clk ) , .D( u1_N38 ) , .Q( u1_R1_7 ) );
  DFF_X1 u1_R1_reg_8 (.CK( clk ) , .D( u1_N39 ) , .Q( u1_R1_8 ) );
  DFF_X1 u1_R1_reg_9 (.CK( clk ) , .D( u1_N40 ) , .Q( u1_R1_9 ) );
  DFF_X1 u1_R2_reg_1 (.CK( clk ) , .D( u1_N64 ) , .Q( u1_R2_1 ) );
  DFF_X1 u1_R2_reg_10 (.CK( clk ) , .D( u1_N73 ) , .Q( u1_R2_10 ) );
  DFF_X1 u1_R2_reg_11 (.CK( clk ) , .D( u1_N74 ) , .Q( u1_R2_11 ) );
  DFF_X1 u1_R2_reg_12 (.CK( clk ) , .D( u1_N75 ) , .Q( u1_R2_12 ) );
  DFF_X1 u1_R2_reg_13 (.CK( clk ) , .D( u1_N76 ) , .Q( u1_R2_13 ) );
  DFF_X1 u1_R2_reg_14 (.CK( clk ) , .D( u1_N77 ) , .Q( u1_R2_14 ) );
  DFF_X1 u1_R2_reg_15 (.CK( clk ) , .D( u1_N78 ) , .Q( u1_R2_15 ) );
  DFF_X1 u1_R2_reg_16 (.CK( clk ) , .D( u1_N79 ) , .Q( u1_R2_16 ) );
  DFF_X1 u1_R2_reg_17 (.CK( clk ) , .D( u1_N80 ) , .Q( u1_R2_17 ) );
  DFF_X1 u1_R2_reg_18 (.CK( clk ) , .D( u1_N81 ) , .Q( u1_R2_18 ) );
  DFF_X1 u1_R2_reg_19 (.CK( clk ) , .D( u1_N82 ) , .Q( u1_R2_19 ) );
  DFF_X1 u1_R2_reg_2 (.CK( clk ) , .D( u1_N65 ) , .Q( u1_R2_2 ) );
  DFF_X1 u1_R2_reg_20 (.CK( clk ) , .D( u1_N83 ) , .Q( u1_R2_20 ) );
  DFF_X1 u1_R2_reg_21 (.CK( clk ) , .D( u1_N84 ) , .Q( u1_R2_21 ) );
  DFF_X1 u1_R2_reg_22 (.CK( clk ) , .D( u1_N85 ) , .Q( u1_R2_22 ) );
  DFF_X1 u1_R2_reg_23 (.CK( clk ) , .D( u1_N86 ) , .Q( u1_R2_23 ) );
  DFF_X1 u1_R2_reg_24 (.CK( clk ) , .D( u1_N87 ) , .Q( u1_R2_24 ) );
  DFF_X1 u1_R2_reg_25 (.CK( clk ) , .D( u1_N88 ) , .Q( u1_R2_25 ) );
  DFF_X1 u1_R2_reg_26 (.CK( clk ) , .D( u1_N89 ) , .Q( u1_R2_26 ) );
  DFF_X1 u1_R2_reg_27 (.CK( clk ) , .D( u1_N90 ) , .Q( u1_R2_27 ) );
  DFF_X1 u1_R2_reg_28 (.CK( clk ) , .D( u1_N91 ) , .Q( u1_R2_28 ) );
  DFF_X1 u1_R2_reg_29 (.CK( clk ) , .D( u1_N92 ) , .Q( u1_R2_29 ) );
  DFF_X1 u1_R2_reg_3 (.CK( clk ) , .D( u1_N66 ) , .Q( u1_R2_3 ) );
  DFF_X1 u1_R2_reg_30 (.CK( clk ) , .D( u1_N93 ) , .Q( u1_R2_30 ) );
  DFF_X1 u1_R2_reg_31 (.CK( clk ) , .D( u1_N94 ) , .Q( u1_R2_31 ) );
  DFF_X1 u1_R2_reg_32 (.CK( clk ) , .D( u1_N95 ) , .Q( u1_R2_32 ) );
  DFF_X1 u1_R2_reg_4 (.CK( clk ) , .D( u1_N67 ) , .Q( u1_R2_4 ) );
  DFF_X1 u1_R2_reg_5 (.CK( clk ) , .D( u1_N68 ) , .Q( u1_R2_5 ) );
  DFF_X1 u1_R2_reg_6 (.CK( clk ) , .D( u1_N69 ) , .Q( u1_R2_6 ) );
  DFF_X1 u1_R2_reg_7 (.CK( clk ) , .D( u1_N70 ) , .Q( u1_R2_7 ) );
  DFF_X1 u1_R2_reg_8 (.CK( clk ) , .D( u1_N71 ) , .Q( u1_R2_8 ) );
  DFF_X1 u1_R2_reg_9 (.CK( clk ) , .D( u1_N72 ) , .Q( u1_R2_9 ) );
  DFF_X1 u1_R3_reg_1 (.CK( clk ) , .D( u1_N96 ) , .Q( u1_R3_1 ) );
  DFF_X1 u1_R3_reg_10 (.CK( clk ) , .D( u1_N105 ) , .Q( u1_R3_10 ) );
  DFF_X1 u1_R3_reg_11 (.CK( clk ) , .D( u1_N106 ) , .Q( u1_R3_11 ) );
  DFF_X1 u1_R3_reg_12 (.CK( clk ) , .D( u1_N107 ) , .Q( u1_R3_12 ) );
  DFF_X1 u1_R3_reg_13 (.CK( clk ) , .D( u1_N108 ) , .Q( u1_R3_13 ) );
  DFF_X1 u1_R3_reg_14 (.CK( clk ) , .D( u1_N109 ) , .Q( u1_R3_14 ) );
  DFF_X1 u1_R3_reg_15 (.CK( clk ) , .D( u1_N110 ) , .Q( u1_R3_15 ) );
  DFF_X1 u1_R3_reg_16 (.CK( clk ) , .D( u1_N111 ) , .Q( u1_R3_16 ) );
  DFF_X1 u1_R3_reg_17 (.CK( clk ) , .D( u1_N112 ) , .Q( u1_R3_17 ) );
  DFF_X1 u1_R3_reg_18 (.CK( clk ) , .D( u1_N113 ) , .Q( u1_R3_18 ) );
  DFF_X1 u1_R3_reg_19 (.CK( clk ) , .D( u1_N114 ) , .Q( u1_R3_19 ) );
  DFF_X1 u1_R3_reg_2 (.CK( clk ) , .D( u1_N97 ) , .Q( u1_R3_2 ) );
  DFF_X1 u1_R3_reg_20 (.CK( clk ) , .D( u1_N115 ) , .Q( u1_R3_20 ) );
  DFF_X1 u1_R3_reg_21 (.CK( clk ) , .D( u1_N116 ) , .Q( u1_R3_21 ) );
  DFF_X1 u1_R3_reg_22 (.CK( clk ) , .D( u1_N117 ) , .Q( u1_R3_22 ) );
  DFF_X1 u1_R3_reg_23 (.CK( clk ) , .D( u1_N118 ) , .Q( u1_R3_23 ) );
  DFF_X1 u1_R3_reg_24 (.CK( clk ) , .D( u1_N119 ) , .Q( u1_R3_24 ) );
  DFF_X1 u1_R3_reg_25 (.CK( clk ) , .D( u1_N120 ) , .Q( u1_R3_25 ) );
  DFF_X1 u1_R3_reg_26 (.CK( clk ) , .D( u1_N121 ) , .Q( u1_R3_26 ) );
  DFF_X1 u1_R3_reg_27 (.CK( clk ) , .D( u1_N122 ) , .Q( u1_R3_27 ) );
  DFF_X1 u1_R3_reg_28 (.CK( clk ) , .D( u1_N123 ) , .Q( u1_R3_28 ) );
  DFF_X1 u1_R3_reg_29 (.CK( clk ) , .D( u1_N124 ) , .Q( u1_R3_29 ) );
  DFF_X1 u1_R3_reg_3 (.CK( clk ) , .D( u1_N98 ) , .Q( u1_R3_3 ) );
  DFF_X1 u1_R3_reg_30 (.CK( clk ) , .D( u1_N125 ) , .Q( u1_R3_30 ) );
  DFF_X1 u1_R3_reg_31 (.CK( clk ) , .D( u1_N126 ) , .Q( u1_R3_31 ) );
  DFF_X1 u1_R3_reg_32 (.CK( clk ) , .D( u1_N127 ) , .Q( u1_R3_32 ) );
  DFF_X1 u1_R3_reg_4 (.CK( clk ) , .D( u1_N99 ) , .Q( u1_R3_4 ) );
  DFF_X1 u1_R3_reg_5 (.CK( clk ) , .D( u1_N100 ) , .Q( u1_R3_5 ) );
  DFF_X1 u1_R3_reg_6 (.CK( clk ) , .D( u1_N101 ) , .Q( u1_R3_6 ) );
  DFF_X1 u1_R3_reg_7 (.CK( clk ) , .D( u1_N102 ) , .Q( u1_R3_7 ) );
  DFF_X1 u1_R3_reg_8 (.CK( clk ) , .D( u1_N103 ) , .Q( u1_R3_8 ) );
  DFF_X1 u1_R3_reg_9 (.CK( clk ) , .D( u1_N104 ) , .Q( u1_R3_9 ) );
  DFF_X1 u1_R4_reg_1 (.CK( clk ) , .D( u1_N128 ) , .Q( u1_R4_1 ) );
  DFF_X1 u1_R4_reg_10 (.CK( clk ) , .D( u1_N137 ) , .Q( u1_R4_10 ) );
  DFF_X1 u1_R4_reg_11 (.CK( clk ) , .D( u1_N138 ) , .Q( u1_R4_11 ) );
  DFF_X1 u1_R4_reg_12 (.CK( clk ) , .D( u1_N139 ) , .Q( u1_R4_12 ) );
  DFF_X1 u1_R4_reg_13 (.CK( clk ) , .D( u1_N140 ) , .Q( u1_R4_13 ) );
  DFF_X1 u1_R4_reg_14 (.CK( clk ) , .D( u1_N141 ) , .Q( u1_R4_14 ) );
  DFF_X1 u1_R4_reg_15 (.CK( clk ) , .D( u1_N142 ) , .Q( u1_R4_15 ) );
  DFF_X1 u1_R4_reg_16 (.CK( clk ) , .D( u1_N143 ) , .Q( u1_R4_16 ) );
  DFF_X1 u1_R4_reg_17 (.CK( clk ) , .D( u1_N144 ) , .Q( u1_R4_17 ) );
  DFF_X1 u1_R4_reg_18 (.CK( clk ) , .D( u1_N145 ) , .Q( u1_R4_18 ) );
  DFF_X1 u1_R4_reg_19 (.CK( clk ) , .D( u1_N146 ) , .Q( u1_R4_19 ) );
  DFF_X1 u1_R4_reg_2 (.CK( clk ) , .D( u1_N129 ) , .Q( u1_R4_2 ) );
  DFF_X1 u1_R4_reg_20 (.CK( clk ) , .D( u1_N147 ) , .Q( u1_R4_20 ) );
  DFF_X1 u1_R4_reg_21 (.CK( clk ) , .D( u1_N148 ) , .Q( u1_R4_21 ) );
  DFF_X1 u1_R4_reg_22 (.CK( clk ) , .D( u1_N149 ) , .Q( u1_R4_22 ) );
  DFF_X1 u1_R4_reg_23 (.CK( clk ) , .D( u1_N150 ) , .Q( u1_R4_23 ) );
  DFF_X1 u1_R4_reg_24 (.CK( clk ) , .D( u1_N151 ) , .Q( u1_R4_24 ) );
  DFF_X1 u1_R4_reg_25 (.CK( clk ) , .D( u1_N152 ) , .Q( u1_R4_25 ) );
  DFF_X1 u1_R4_reg_26 (.CK( clk ) , .D( u1_N153 ) , .Q( u1_R4_26 ) );
  DFF_X1 u1_R4_reg_27 (.CK( clk ) , .D( u1_N154 ) , .Q( u1_R4_27 ) );
  DFF_X1 u1_R4_reg_28 (.CK( clk ) , .D( u1_N155 ) , .Q( u1_R4_28 ) );
  DFF_X1 u1_R4_reg_29 (.CK( clk ) , .D( u1_N156 ) , .Q( u1_R4_29 ) );
  DFF_X1 u1_R4_reg_3 (.CK( clk ) , .D( u1_N130 ) , .Q( u1_R4_3 ) );
  DFF_X1 u1_R4_reg_30 (.CK( clk ) , .D( u1_N157 ) , .Q( u1_R4_30 ) );
  DFF_X1 u1_R4_reg_31 (.CK( clk ) , .D( u1_N158 ) , .Q( u1_R4_31 ) );
  DFF_X1 u1_R4_reg_32 (.CK( clk ) , .D( u1_N159 ) , .Q( u1_R4_32 ) );
  DFF_X1 u1_R4_reg_4 (.CK( clk ) , .D( u1_N131 ) , .Q( u1_R4_4 ) );
  DFF_X1 u1_R4_reg_5 (.CK( clk ) , .D( u1_N132 ) , .Q( u1_R4_5 ) );
  DFF_X1 u1_R4_reg_6 (.CK( clk ) , .D( u1_N133 ) , .Q( u1_R4_6 ) );
  DFF_X1 u1_R4_reg_7 (.CK( clk ) , .D( u1_N134 ) , .Q( u1_R4_7 ) );
  DFF_X1 u1_R4_reg_8 (.CK( clk ) , .D( u1_N135 ) , .Q( u1_R4_8 ) );
  DFF_X1 u1_R4_reg_9 (.CK( clk ) , .D( u1_N136 ) , .Q( u1_R4_9 ) );
  DFF_X1 u1_R5_reg_1 (.CK( clk ) , .D( u1_N160 ) , .Q( u1_R5_1 ) );
  DFF_X1 u1_R5_reg_10 (.CK( clk ) , .D( u1_N169 ) , .Q( u1_R5_10 ) );
  DFF_X1 u1_R5_reg_11 (.CK( clk ) , .D( u1_N170 ) , .Q( u1_R5_11 ) );
  DFF_X1 u1_R5_reg_12 (.CK( clk ) , .D( u1_N171 ) , .Q( u1_R5_12 ) );
  DFF_X1 u1_R5_reg_13 (.CK( clk ) , .D( u1_N172 ) , .Q( u1_R5_13 ) );
  DFF_X1 u1_R5_reg_14 (.CK( clk ) , .D( u1_N173 ) , .Q( u1_R5_14 ) );
  DFF_X1 u1_R5_reg_15 (.CK( clk ) , .D( u1_N174 ) , .Q( u1_R5_15 ) );
  DFF_X1 u1_R5_reg_16 (.CK( clk ) , .D( u1_N175 ) , .Q( u1_R5_16 ) );
  DFF_X1 u1_R5_reg_17 (.CK( clk ) , .D( u1_N176 ) , .Q( u1_R5_17 ) );
  DFF_X1 u1_R5_reg_18 (.CK( clk ) , .D( u1_N177 ) , .Q( u1_R5_18 ) );
  DFF_X1 u1_R5_reg_19 (.CK( clk ) , .D( u1_N178 ) , .Q( u1_R5_19 ) );
  DFF_X1 u1_R5_reg_2 (.CK( clk ) , .D( u1_N161 ) , .Q( u1_R5_2 ) );
  DFF_X1 u1_R5_reg_20 (.CK( clk ) , .D( u1_N179 ) , .Q( u1_R5_20 ) );
  DFF_X1 u1_R5_reg_21 (.CK( clk ) , .D( u1_N180 ) , .Q( u1_R5_21 ) );
  DFF_X1 u1_R5_reg_22 (.CK( clk ) , .D( u1_N181 ) , .Q( u1_R5_22 ) );
  DFF_X1 u1_R5_reg_23 (.CK( clk ) , .D( u1_N182 ) , .Q( u1_R5_23 ) );
  DFF_X1 u1_R5_reg_24 (.CK( clk ) , .D( u1_N183 ) , .Q( u1_R5_24 ) );
  DFF_X1 u1_R5_reg_25 (.CK( clk ) , .D( u1_N184 ) , .Q( u1_R5_25 ) );
  DFF_X1 u1_R5_reg_26 (.CK( clk ) , .D( u1_N185 ) , .Q( u1_R5_26 ) );
  DFF_X1 u1_R5_reg_27 (.CK( clk ) , .D( u1_N186 ) , .Q( u1_R5_27 ) );
  DFF_X1 u1_R5_reg_28 (.CK( clk ) , .D( u1_N187 ) , .Q( u1_R5_28 ) );
  DFF_X1 u1_R5_reg_29 (.CK( clk ) , .D( u1_N188 ) , .Q( u1_R5_29 ) );
  DFF_X1 u1_R5_reg_3 (.CK( clk ) , .D( u1_N162 ) , .Q( u1_R5_3 ) );
  DFF_X1 u1_R5_reg_30 (.CK( clk ) , .D( u1_N189 ) , .Q( u1_R5_30 ) );
  DFF_X1 u1_R5_reg_31 (.CK( clk ) , .D( u1_N190 ) , .Q( u1_R5_31 ) );
  DFF_X1 u1_R5_reg_32 (.CK( clk ) , .D( u1_N191 ) , .Q( u1_R5_32 ) );
  DFF_X1 u1_R5_reg_4 (.CK( clk ) , .D( u1_N163 ) , .Q( u1_R5_4 ) );
  DFF_X1 u1_R5_reg_5 (.CK( clk ) , .D( u1_N164 ) , .Q( u1_R5_5 ) );
  DFF_X1 u1_R5_reg_6 (.CK( clk ) , .D( u1_N165 ) , .Q( u1_R5_6 ) );
  DFF_X1 u1_R5_reg_7 (.CK( clk ) , .D( u1_N166 ) , .Q( u1_R5_7 ) );
  DFF_X1 u1_R5_reg_8 (.CK( clk ) , .D( u1_N167 ) , .Q( u1_R5_8 ) );
  DFF_X1 u1_R5_reg_9 (.CK( clk ) , .D( u1_N168 ) , .Q( u1_R5_9 ) );
  DFF_X1 u1_R6_reg_1 (.CK( clk ) , .D( u1_N192 ) , .Q( u1_R6_1 ) );
  DFF_X1 u1_R6_reg_10 (.CK( clk ) , .D( u1_N201 ) , .Q( u1_R6_10 ) );
  DFF_X1 u1_R6_reg_11 (.CK( clk ) , .D( u1_N202 ) , .Q( u1_R6_11 ) );
  DFF_X1 u1_R6_reg_12 (.CK( clk ) , .D( u1_N203 ) , .Q( u1_R6_12 ) );
  DFF_X1 u1_R6_reg_13 (.CK( clk ) , .D( u1_N204 ) , .Q( u1_R6_13 ) );
  DFF_X1 u1_R6_reg_14 (.CK( clk ) , .D( u1_N205 ) , .Q( u1_R6_14 ) );
  DFF_X1 u1_R6_reg_15 (.CK( clk ) , .D( u1_N206 ) , .Q( u1_R6_15 ) );
  DFF_X1 u1_R6_reg_16 (.CK( clk ) , .D( u1_N207 ) , .Q( u1_R6_16 ) );
  DFF_X1 u1_R6_reg_17 (.CK( clk ) , .D( u1_N208 ) , .Q( u1_R6_17 ) );
  DFF_X1 u1_R6_reg_18 (.CK( clk ) , .D( u1_N209 ) , .Q( u1_R6_18 ) );
  DFF_X1 u1_R6_reg_19 (.CK( clk ) , .D( u1_N210 ) , .Q( u1_R6_19 ) );
  DFF_X1 u1_R6_reg_2 (.CK( clk ) , .D( u1_N193 ) , .Q( u1_R6_2 ) );
  DFF_X1 u1_R6_reg_20 (.CK( clk ) , .D( u1_N211 ) , .Q( u1_R6_20 ) );
  DFF_X1 u1_R6_reg_21 (.CK( clk ) , .D( u1_N212 ) , .Q( u1_R6_21 ) );
  DFF_X1 u1_R6_reg_22 (.CK( clk ) , .D( u1_N213 ) , .Q( u1_R6_22 ) );
  DFF_X1 u1_R6_reg_23 (.CK( clk ) , .D( u1_N214 ) , .Q( u1_R6_23 ) );
  DFF_X1 u1_R6_reg_24 (.CK( clk ) , .D( u1_N215 ) , .Q( u1_R6_24 ) );
  DFF_X1 u1_R6_reg_25 (.CK( clk ) , .D( u1_N216 ) , .Q( u1_R6_25 ) );
  DFF_X1 u1_R6_reg_26 (.CK( clk ) , .D( u1_N217 ) , .Q( u1_R6_26 ) );
  DFF_X1 u1_R6_reg_27 (.CK( clk ) , .D( u1_N218 ) , .Q( u1_R6_27 ) );
  DFF_X1 u1_R6_reg_28 (.CK( clk ) , .D( u1_N219 ) , .Q( u1_R6_28 ) );
  DFF_X1 u1_R6_reg_29 (.CK( clk ) , .D( u1_N220 ) , .Q( u1_R6_29 ) );
  DFF_X1 u1_R6_reg_3 (.CK( clk ) , .D( u1_N194 ) , .Q( u1_R6_3 ) );
  DFF_X1 u1_R6_reg_30 (.CK( clk ) , .D( u1_N221 ) , .Q( u1_R6_30 ) );
  DFF_X1 u1_R6_reg_31 (.CK( clk ) , .D( u1_N222 ) , .Q( u1_R6_31 ) );
  DFF_X1 u1_R6_reg_32 (.CK( clk ) , .D( u1_N223 ) , .Q( u1_R6_32 ) );
  DFF_X1 u1_R6_reg_4 (.CK( clk ) , .D( u1_N195 ) , .Q( u1_R6_4 ) );
  DFF_X1 u1_R6_reg_5 (.CK( clk ) , .D( u1_N196 ) , .Q( u1_R6_5 ) );
  DFF_X1 u1_R6_reg_6 (.CK( clk ) , .D( u1_N197 ) , .Q( u1_R6_6 ) );
  DFF_X1 u1_R6_reg_7 (.CK( clk ) , .D( u1_N198 ) , .Q( u1_R6_7 ) );
  DFF_X1 u1_R6_reg_8 (.CK( clk ) , .D( u1_N199 ) , .Q( u1_R6_8 ) );
  DFF_X1 u1_R6_reg_9 (.CK( clk ) , .D( u1_N200 ) , .Q( u1_R6_9 ) );
  DFF_X1 u1_R7_reg_1 (.CK( clk ) , .D( u1_N224 ) , .Q( u1_R7_1 ) );
  DFF_X1 u1_R7_reg_10 (.CK( clk ) , .D( u1_N233 ) , .Q( u1_R7_10 ) );
  DFF_X1 u1_R7_reg_11 (.CK( clk ) , .D( u1_N234 ) , .Q( u1_R7_11 ) );
  DFF_X1 u1_R7_reg_12 (.CK( clk ) , .D( u1_N235 ) , .Q( u1_R7_12 ) );
  DFF_X1 u1_R7_reg_13 (.CK( clk ) , .D( u1_N236 ) , .Q( u1_R7_13 ) );
  DFF_X1 u1_R7_reg_14 (.CK( clk ) , .D( u1_N237 ) , .Q( u1_R7_14 ) );
  DFF_X1 u1_R7_reg_15 (.CK( clk ) , .D( u1_N238 ) , .Q( u1_R7_15 ) );
  DFF_X1 u1_R7_reg_16 (.CK( clk ) , .D( u1_N239 ) , .Q( u1_R7_16 ) );
  DFF_X1 u1_R7_reg_17 (.CK( clk ) , .D( u1_N240 ) , .Q( u1_R7_17 ) );
  DFF_X1 u1_R7_reg_18 (.CK( clk ) , .D( u1_N241 ) , .Q( u1_R7_18 ) );
  DFF_X1 u1_R7_reg_19 (.CK( clk ) , .D( u1_N242 ) , .Q( u1_R7_19 ) );
  DFF_X1 u1_R7_reg_2 (.CK( clk ) , .D( u1_N225 ) , .Q( u1_R7_2 ) );
  DFF_X1 u1_R7_reg_20 (.CK( clk ) , .D( u1_N243 ) , .Q( u1_R7_20 ) );
  DFF_X1 u1_R7_reg_21 (.CK( clk ) , .D( u1_N244 ) , .Q( u1_R7_21 ) );
  DFF_X1 u1_R7_reg_22 (.CK( clk ) , .D( u1_N245 ) , .Q( u1_R7_22 ) );
  DFF_X1 u1_R7_reg_23 (.CK( clk ) , .D( u1_N246 ) , .Q( u1_R7_23 ) );
  DFF_X1 u1_R7_reg_24 (.CK( clk ) , .D( u1_N247 ) , .Q( u1_R7_24 ) );
  DFF_X1 u1_R7_reg_25 (.CK( clk ) , .D( u1_N248 ) , .Q( u1_R7_25 ) );
  DFF_X1 u1_R7_reg_26 (.CK( clk ) , .D( u1_N249 ) , .Q( u1_R7_26 ) );
  DFF_X1 u1_R7_reg_27 (.CK( clk ) , .D( u1_N250 ) , .Q( u1_R7_27 ) );
  DFF_X1 u1_R7_reg_28 (.CK( clk ) , .D( u1_N251 ) , .Q( u1_R7_28 ) );
  DFF_X1 u1_R7_reg_29 (.CK( clk ) , .D( u1_N252 ) , .Q( u1_R7_29 ) );
  DFF_X1 u1_R7_reg_3 (.CK( clk ) , .D( u1_N226 ) , .Q( u1_R7_3 ) );
  DFF_X1 u1_R7_reg_30 (.CK( clk ) , .D( u1_N253 ) , .Q( u1_R7_30 ) );
  DFF_X1 u1_R7_reg_31 (.CK( clk ) , .D( u1_N254 ) , .Q( u1_R7_31 ) );
  DFF_X1 u1_R7_reg_32 (.CK( clk ) , .D( u1_N255 ) , .Q( u1_R7_32 ) );
  DFF_X1 u1_R7_reg_4 (.CK( clk ) , .D( u1_N227 ) , .Q( u1_R7_4 ) );
  DFF_X1 u1_R7_reg_5 (.CK( clk ) , .D( u1_N228 ) , .Q( u1_R7_5 ) );
  DFF_X1 u1_R7_reg_6 (.CK( clk ) , .D( u1_N229 ) , .Q( u1_R7_6 ) );
  DFF_X1 u1_R7_reg_7 (.CK( clk ) , .D( u1_N230 ) , .Q( u1_R7_7 ) );
  DFF_X1 u1_R7_reg_8 (.CK( clk ) , .D( u1_N231 ) , .Q( u1_R7_8 ) );
  DFF_X1 u1_R7_reg_9 (.CK( clk ) , .D( u1_N232 ) , .Q( u1_R7_9 ) );
  DFF_X1 u1_R8_reg_1 (.CK( clk ) , .D( u1_N256 ) , .Q( u1_R8_1 ) );
  DFF_X1 u1_R8_reg_10 (.CK( clk ) , .D( u1_N265 ) , .Q( u1_R8_10 ) );
  DFF_X1 u1_R8_reg_11 (.CK( clk ) , .D( u1_N266 ) , .Q( u1_R8_11 ) );
  DFF_X1 u1_R8_reg_12 (.CK( clk ) , .D( u1_N267 ) , .Q( u1_R8_12 ) );
  DFF_X1 u1_R8_reg_13 (.CK( clk ) , .D( u1_N268 ) , .Q( u1_R8_13 ) );
  DFF_X1 u1_R8_reg_14 (.CK( clk ) , .D( u1_N269 ) , .Q( u1_R8_14 ) );
  DFF_X1 u1_R8_reg_15 (.CK( clk ) , .D( u1_N270 ) , .Q( u1_R8_15 ) );
  DFF_X1 u1_R8_reg_16 (.CK( clk ) , .D( u1_N271 ) , .Q( u1_R8_16 ) );
  DFF_X1 u1_R8_reg_17 (.CK( clk ) , .D( u1_N272 ) , .Q( u1_R8_17 ) );
  DFF_X1 u1_R8_reg_18 (.CK( clk ) , .D( u1_N273 ) , .Q( u1_R8_18 ) );
  DFF_X1 u1_R8_reg_19 (.CK( clk ) , .D( u1_N274 ) , .Q( u1_R8_19 ) );
  DFF_X1 u1_R8_reg_2 (.CK( clk ) , .D( u1_N257 ) , .Q( u1_R8_2 ) );
  DFF_X1 u1_R8_reg_20 (.CK( clk ) , .D( u1_N275 ) , .Q( u1_R8_20 ) );
  DFF_X1 u1_R8_reg_21 (.CK( clk ) , .D( u1_N276 ) , .Q( u1_R8_21 ) );
  DFF_X1 u1_R8_reg_22 (.CK( clk ) , .D( u1_N277 ) , .Q( u1_R8_22 ) );
  DFF_X1 u1_R8_reg_23 (.CK( clk ) , .D( u1_N278 ) , .Q( u1_R8_23 ) );
  DFF_X1 u1_R8_reg_24 (.CK( clk ) , .D( u1_N279 ) , .Q( u1_R8_24 ) );
  DFF_X1 u1_R8_reg_25 (.CK( clk ) , .D( u1_N280 ) , .Q( u1_R8_25 ) );
  DFF_X1 u1_R8_reg_26 (.CK( clk ) , .D( u1_N281 ) , .Q( u1_R8_26 ) );
  DFF_X1 u1_R8_reg_27 (.CK( clk ) , .D( u1_N282 ) , .Q( u1_R8_27 ) );
  DFF_X1 u1_R8_reg_28 (.CK( clk ) , .D( u1_N283 ) , .Q( u1_R8_28 ) );
  DFF_X1 u1_R8_reg_29 (.CK( clk ) , .D( u1_N284 ) , .Q( u1_R8_29 ) );
  DFF_X1 u1_R8_reg_3 (.CK( clk ) , .D( u1_N258 ) , .Q( u1_R8_3 ) );
  DFF_X1 u1_R8_reg_30 (.CK( clk ) , .D( u1_N285 ) , .Q( u1_R8_30 ) );
  DFF_X1 u1_R8_reg_31 (.CK( clk ) , .D( u1_N286 ) , .Q( u1_R8_31 ) );
  DFF_X1 u1_R8_reg_32 (.CK( clk ) , .D( u1_N287 ) , .Q( u1_R8_32 ) );
  DFF_X1 u1_R8_reg_4 (.CK( clk ) , .D( u1_N259 ) , .Q( u1_R8_4 ) );
  DFF_X1 u1_R8_reg_5 (.CK( clk ) , .D( u1_N260 ) , .Q( u1_R8_5 ) );
  DFF_X1 u1_R8_reg_6 (.CK( clk ) , .D( u1_N261 ) , .Q( u1_R8_6 ) );
  DFF_X1 u1_R8_reg_7 (.CK( clk ) , .D( u1_N262 ) , .Q( u1_R8_7 ) );
  DFF_X1 u1_R8_reg_8 (.CK( clk ) , .D( u1_N263 ) , .Q( u1_R8_8 ) );
  DFF_X1 u1_R8_reg_9 (.CK( clk ) , .D( u1_N264 ) , .Q( u1_R8_9 ) );
  DFF_X1 u1_R9_reg_1 (.CK( clk ) , .D( u1_N288 ) , .Q( u1_R9_1 ) );
  DFF_X1 u1_R9_reg_10 (.CK( clk ) , .D( u1_N297 ) , .Q( u1_R9_10 ) );
  DFF_X1 u1_R9_reg_11 (.CK( clk ) , .D( u1_N298 ) , .Q( u1_R9_11 ) );
  DFF_X1 u1_R9_reg_12 (.CK( clk ) , .D( u1_N299 ) , .Q( u1_R9_12 ) );
  DFF_X1 u1_R9_reg_13 (.CK( clk ) , .D( u1_N300 ) , .Q( u1_R9_13 ) );
  DFF_X1 u1_R9_reg_14 (.CK( clk ) , .D( u1_N301 ) , .Q( u1_R9_14 ) );
  DFF_X1 u1_R9_reg_15 (.CK( clk ) , .D( u1_N302 ) , .Q( u1_R9_15 ) );
  DFF_X1 u1_R9_reg_16 (.CK( clk ) , .D( u1_N303 ) , .Q( u1_R9_16 ) );
  DFF_X1 u1_R9_reg_17 (.CK( clk ) , .D( u1_N304 ) , .Q( u1_R9_17 ) );
  DFF_X1 u1_R9_reg_18 (.CK( clk ) , .D( u1_N305 ) , .Q( u1_R9_18 ) );
  DFF_X1 u1_R9_reg_19 (.CK( clk ) , .D( u1_N306 ) , .Q( u1_R9_19 ) );
  DFF_X1 u1_R9_reg_2 (.CK( clk ) , .D( u1_N289 ) , .Q( u1_R9_2 ) );
  DFF_X1 u1_R9_reg_20 (.CK( clk ) , .D( u1_N307 ) , .Q( u1_R9_20 ) );
  DFF_X1 u1_R9_reg_21 (.CK( clk ) , .D( u1_N308 ) , .Q( u1_R9_21 ) );
  DFF_X1 u1_R9_reg_22 (.CK( clk ) , .D( u1_N309 ) , .Q( u1_R9_22 ) );
  DFF_X1 u1_R9_reg_23 (.CK( clk ) , .D( u1_N310 ) , .Q( u1_R9_23 ) );
  DFF_X1 u1_R9_reg_24 (.CK( clk ) , .D( u1_N311 ) , .Q( u1_R9_24 ) );
  DFF_X1 u1_R9_reg_25 (.CK( clk ) , .D( u1_N312 ) , .Q( u1_R9_25 ) );
  DFF_X1 u1_R9_reg_26 (.CK( clk ) , .D( u1_N313 ) , .Q( u1_R9_26 ) );
  DFF_X1 u1_R9_reg_27 (.CK( clk ) , .D( u1_N314 ) , .Q( u1_R9_27 ) );
  DFF_X1 u1_R9_reg_28 (.CK( clk ) , .D( u1_N315 ) , .Q( u1_R9_28 ) );
  DFF_X1 u1_R9_reg_29 (.CK( clk ) , .D( u1_N316 ) , .Q( u1_R9_29 ) );
  DFF_X1 u1_R9_reg_3 (.CK( clk ) , .D( u1_N290 ) , .Q( u1_R9_3 ) );
  DFF_X1 u1_R9_reg_30 (.CK( clk ) , .D( u1_N317 ) , .Q( u1_R9_30 ) );
  DFF_X1 u1_R9_reg_31 (.CK( clk ) , .D( u1_N318 ) , .Q( u1_R9_31 ) );
  DFF_X1 u1_R9_reg_32 (.CK( clk ) , .D( u1_N319 ) , .Q( u1_R9_32 ) );
  DFF_X1 u1_R9_reg_4 (.CK( clk ) , .D( u1_N291 ) , .Q( u1_R9_4 ) );
  DFF_X1 u1_R9_reg_5 (.CK( clk ) , .D( u1_N292 ) , .Q( u1_R9_5 ) );
  DFF_X1 u1_R9_reg_6 (.CK( clk ) , .D( u1_N293 ) , .Q( u1_R9_6 ) );
  DFF_X1 u1_R9_reg_7 (.CK( clk ) , .D( u1_N294 ) , .Q( u1_R9_7 ) );
  DFF_X1 u1_R9_reg_8 (.CK( clk ) , .D( u1_N295 ) , .Q( u1_R9_8 ) );
  DFF_X1 u1_R9_reg_9 (.CK( clk ) , .D( u1_N296 ) , .Q( u1_R9_9 ) );
  XOR2_X1 u1_U10 (.B( u1_L1_29 ) , .Z( u1_N92 ) , .A( u1_out2_29 ) );
  XOR2_X1 u1_U100 (.B( u1_L12_27 ) , .Z( u1_N442 ) , .A( u1_out13_27 ) );
  XOR2_X1 u1_U101 (.B( u1_L12_26 ) , .Z( u1_N441 ) , .A( u1_out13_26 ) );
  XOR2_X1 u1_U102 (.B( u1_L12_25 ) , .Z( u1_N440 ) , .A( u1_out13_25 ) );
  XOR2_X1 u1_U103 (.B( u1_L0_13 ) , .Z( u1_N44 ) , .A( u1_out1_13 ) );
  XOR2_X1 u1_U104 (.B( u1_L12_24 ) , .Z( u1_N439 ) , .A( u1_out13_24 ) );
  XOR2_X1 u1_U105 (.B( u1_L12_23 ) , .Z( u1_N438 ) , .A( u1_out13_23 ) );
  XOR2_X1 u1_U106 (.B( u1_L12_22 ) , .Z( u1_N437 ) , .A( u1_out13_22 ) );
  XOR2_X1 u1_U107 (.B( u1_L12_21 ) , .Z( u1_N436 ) , .A( u1_out13_21 ) );
  XOR2_X1 u1_U108 (.B( u1_L12_20 ) , .Z( u1_N435 ) , .A( u1_out13_20 ) );
  XOR2_X1 u1_U109 (.B( u1_L12_19 ) , .Z( u1_N434 ) , .A( u1_out13_19 ) );
  XOR2_X1 u1_U11 (.B( u1_L1_28 ) , .Z( u1_N91 ) , .A( u1_out2_28 ) );
  XOR2_X1 u1_U110 (.B( u1_L12_18 ) , .Z( u1_N433 ) , .A( u1_out13_18 ) );
  XOR2_X1 u1_U111 (.B( u1_L12_17 ) , .Z( u1_N432 ) , .A( u1_out13_17 ) );
  XOR2_X1 u1_U112 (.B( u1_L12_16 ) , .Z( u1_N431 ) , .A( u1_out13_16 ) );
  XOR2_X1 u1_U113 (.B( u1_L12_15 ) , .Z( u1_N430 ) , .A( u1_out13_15 ) );
  XOR2_X1 u1_U114 (.B( u1_L0_12 ) , .Z( u1_N43 ) , .A( u1_out1_12 ) );
  XOR2_X1 u1_U115 (.B( u1_L12_14 ) , .Z( u1_N429 ) , .A( u1_out13_14 ) );
  XOR2_X1 u1_U116 (.B( u1_L12_13 ) , .Z( u1_N428 ) , .A( u1_out13_13 ) );
  XOR2_X1 u1_U117 (.B( u1_L12_12 ) , .Z( u1_N427 ) , .A( u1_out13_12 ) );
  XOR2_X1 u1_U118 (.B( u1_L12_11 ) , .Z( u1_N426 ) , .A( u1_out13_11 ) );
  XOR2_X1 u1_U119 (.B( u1_L12_10 ) , .Z( u1_N425 ) , .A( u1_out13_10 ) );
  XOR2_X1 u1_U12 (.B( u1_L1_27 ) , .Z( u1_N90 ) , .A( u1_out2_27 ) );
  XOR2_X1 u1_U120 (.B( u1_L12_9 ) , .Z( u1_N424 ) , .A( u1_out13_9 ) );
  XOR2_X1 u1_U121 (.B( u1_L12_8 ) , .Z( u1_N423 ) , .A( u1_out13_8 ) );
  XOR2_X1 u1_U122 (.B( u1_L12_7 ) , .Z( u1_N422 ) , .A( u1_out13_7 ) );
  XOR2_X1 u1_U123 (.B( u1_L12_6 ) , .Z( u1_N421 ) , .A( u1_out13_6 ) );
  XOR2_X1 u1_U124 (.B( u1_L12_5 ) , .Z( u1_N420 ) , .A( u1_out13_5 ) );
  XOR2_X1 u1_U125 (.B( u1_L0_11 ) , .Z( u1_N42 ) , .A( u1_out1_11 ) );
  XOR2_X1 u1_U126 (.B( u1_L12_4 ) , .Z( u1_N419 ) , .A( u1_out13_4 ) );
  XOR2_X1 u1_U127 (.B( u1_L12_3 ) , .Z( u1_N418 ) , .A( u1_out13_3 ) );
  XOR2_X1 u1_U128 (.B( u1_L12_2 ) , .Z( u1_N417 ) , .A( u1_out13_2 ) );
  XOR2_X1 u1_U129 (.B( u1_L12_1 ) , .Z( u1_N416 ) , .A( u1_out13_1 ) );
  XOR2_X1 u1_U13 (.Z( u1_N9 ) , .B( u1_desIn_r_12 ) , .A( u1_out0_10 ) );
  XOR2_X1 u1_U130 (.B( u1_L11_32 ) , .Z( u1_N415 ) , .A( u1_out12_32 ) );
  XOR2_X1 u1_U131 (.B( u1_L11_31 ) , .Z( u1_N414 ) , .A( u1_out12_31 ) );
  XOR2_X1 u1_U132 (.B( u1_L11_30 ) , .Z( u1_N413 ) , .A( u1_out12_30 ) );
  XOR2_X1 u1_U133 (.B( u1_L11_29 ) , .Z( u1_N412 ) , .A( u1_out12_29 ) );
  XOR2_X1 u1_U134 (.B( u1_L11_28 ) , .Z( u1_N411 ) , .A( u1_out12_28 ) );
  XOR2_X1 u1_U135 (.B( u1_L11_27 ) , .Z( u1_N410 ) , .A( u1_out12_27 ) );
  XOR2_X1 u1_U136 (.B( u1_L0_10 ) , .Z( u1_N41 ) , .A( u1_out1_10 ) );
  XOR2_X1 u1_U137 (.B( u1_L11_26 ) , .Z( u1_N409 ) , .A( u1_out12_26 ) );
  XOR2_X1 u1_U138 (.B( u1_L11_25 ) , .Z( u1_N408 ) , .A( u1_out12_25 ) );
  XOR2_X1 u1_U139 (.B( u1_L11_24 ) , .Z( u1_N407 ) , .A( u1_out12_24 ) );
  XOR2_X1 u1_U14 (.B( u1_L1_26 ) , .Z( u1_N89 ) , .A( u1_out2_26 ) );
  XOR2_X1 u1_U140 (.B( u1_L11_23 ) , .Z( u1_N406 ) , .A( u1_out12_23 ) );
  XOR2_X1 u1_U141 (.B( u1_L11_22 ) , .Z( u1_N405 ) , .A( u1_out12_22 ) );
  XOR2_X1 u1_U142 (.B( u1_L11_21 ) , .Z( u1_N404 ) , .A( u1_out12_21 ) );
  XOR2_X1 u1_U143 (.B( u1_L11_20 ) , .Z( u1_N403 ) , .A( u1_out12_20 ) );
  XOR2_X1 u1_U144 (.B( u1_L11_19 ) , .Z( u1_N402 ) , .A( u1_out12_19 ) );
  XOR2_X1 u1_U145 (.B( u1_L11_18 ) , .Z( u1_N401 ) , .A( u1_out12_18 ) );
  XOR2_X1 u1_U146 (.B( u1_L11_17 ) , .Z( u1_N400 ) , .A( u1_out12_17 ) );
  XOR2_X1 u1_U147 (.B( u1_L0_9 ) , .Z( u1_N40 ) , .A( u1_out1_9 ) );
  XOR2_X1 u1_U148 (.Z( u1_N4 ) , .B( u1_desIn_r_38 ) , .A( u1_out0_5 ) );
  XOR2_X1 u1_U149 (.B( u1_L11_16 ) , .Z( u1_N399 ) , .A( u1_out12_16 ) );
  XOR2_X1 u1_U15 (.B( u1_L1_25 ) , .Z( u1_N88 ) , .A( u1_out2_25 ) );
  XOR2_X1 u1_U150 (.B( u1_L11_15 ) , .Z( u1_N398 ) , .A( u1_out12_15 ) );
  XOR2_X1 u1_U151 (.B( u1_L11_14 ) , .Z( u1_N397 ) , .A( u1_out12_14 ) );
  XOR2_X1 u1_U152 (.B( u1_L11_13 ) , .Z( u1_N396 ) , .A( u1_out12_13 ) );
  XOR2_X1 u1_U153 (.B( u1_L11_12 ) , .Z( u1_N395 ) , .A( u1_out12_12 ) );
  XOR2_X1 u1_U154 (.B( u1_L11_11 ) , .Z( u1_N394 ) , .A( u1_out12_11 ) );
  XOR2_X1 u1_U155 (.B( u1_L11_10 ) , .Z( u1_N393 ) , .A( u1_out12_10 ) );
  XOR2_X1 u1_U156 (.B( u1_L11_9 ) , .Z( u1_N392 ) , .A( u1_out12_9 ) );
  XOR2_X1 u1_U157 (.B( u1_L11_8 ) , .Z( u1_N391 ) , .A( u1_out12_8 ) );
  XOR2_X1 u1_U158 (.B( u1_L11_7 ) , .Z( u1_N390 ) , .A( u1_out12_7 ) );
  XOR2_X1 u1_U159 (.B( u1_L0_8 ) , .Z( u1_N39 ) , .A( u1_out1_8 ) );
  XOR2_X1 u1_U16 (.B( u1_L1_24 ) , .Z( u1_N87 ) , .A( u1_out2_24 ) );
  XOR2_X1 u1_U160 (.B( u1_L11_6 ) , .Z( u1_N389 ) , .A( u1_out12_6 ) );
  XOR2_X1 u1_U161 (.B( u1_L11_5 ) , .Z( u1_N388 ) , .A( u1_out12_5 ) );
  XOR2_X1 u1_U162 (.B( u1_L11_4 ) , .Z( u1_N387 ) , .A( u1_out12_4 ) );
  XOR2_X1 u1_U163 (.B( u1_L11_3 ) , .Z( u1_N386 ) , .A( u1_out12_3 ) );
  XOR2_X1 u1_U164 (.B( u1_L11_2 ) , .Z( u1_N385 ) , .A( u1_out12_2 ) );
  XOR2_X1 u1_U165 (.B( u1_L11_1 ) , .Z( u1_N384 ) , .A( u1_out12_1 ) );
  XOR2_X1 u1_U166 (.B( u1_L10_32 ) , .Z( u1_N383 ) , .A( u1_out11_32 ) );
  XOR2_X1 u1_U167 (.B( u1_L10_31 ) , .Z( u1_N382 ) , .A( u1_out11_31 ) );
  XOR2_X1 u1_U168 (.B( u1_L10_30 ) , .Z( u1_N381 ) , .A( u1_out11_30 ) );
  XOR2_X1 u1_U169 (.B( u1_L10_29 ) , .Z( u1_N380 ) , .A( u1_out11_29 ) );
  XOR2_X1 u1_U17 (.B( u1_L1_23 ) , .Z( u1_N86 ) , .A( u1_out2_23 ) );
  XOR2_X1 u1_U170 (.B( u1_L0_7 ) , .Z( u1_N38 ) , .A( u1_out1_7 ) );
  XOR2_X1 u1_U171 (.B( u1_L10_28 ) , .Z( u1_N379 ) , .A( u1_out11_28 ) );
  XOR2_X1 u1_U172 (.B( u1_L10_27 ) , .Z( u1_N378 ) , .A( u1_out11_27 ) );
  XOR2_X1 u1_U173 (.B( u1_L10_26 ) , .Z( u1_N377 ) , .A( u1_out11_26 ) );
  XOR2_X1 u1_U174 (.B( u1_L10_25 ) , .Z( u1_N376 ) , .A( u1_out11_25 ) );
  XOR2_X1 u1_U175 (.B( u1_L10_24 ) , .Z( u1_N375 ) , .A( u1_out11_24 ) );
  XOR2_X1 u1_U176 (.B( u1_L10_23 ) , .Z( u1_N374 ) , .A( u1_out11_23 ) );
  XOR2_X1 u1_U177 (.B( u1_L10_22 ) , .Z( u1_N373 ) , .A( u1_out11_22 ) );
  XOR2_X1 u1_U178 (.B( u1_L10_21 ) , .Z( u1_N372 ) , .A( u1_out11_21 ) );
  XOR2_X1 u1_U179 (.B( u1_L10_20 ) , .Z( u1_N371 ) , .A( u1_out11_20 ) );
  XOR2_X1 u1_U18 (.B( u1_L1_22 ) , .Z( u1_N85 ) , .A( u1_out2_22 ) );
  XOR2_X1 u1_U180 (.B( u1_L10_19 ) , .Z( u1_N370 ) , .A( u1_out11_19 ) );
  XOR2_X1 u1_U181 (.B( u1_L0_6 ) , .Z( u1_N37 ) , .A( u1_out1_6 ) );
  XOR2_X1 u1_U182 (.B( u1_L10_18 ) , .Z( u1_N369 ) , .A( u1_out11_18 ) );
  XOR2_X1 u1_U183 (.B( u1_L10_17 ) , .Z( u1_N368 ) , .A( u1_out11_17 ) );
  XOR2_X1 u1_U184 (.B( u1_L10_16 ) , .Z( u1_N367 ) , .A( u1_out11_16 ) );
  XOR2_X1 u1_U185 (.B( u1_L10_15 ) , .Z( u1_N366 ) , .A( u1_out11_15 ) );
  XOR2_X1 u1_U186 (.B( u1_L10_14 ) , .Z( u1_N365 ) , .A( u1_out11_14 ) );
  XOR2_X1 u1_U187 (.B( u1_L10_13 ) , .Z( u1_N364 ) , .A( u1_out11_13 ) );
  XOR2_X1 u1_U188 (.B( u1_L10_12 ) , .Z( u1_N363 ) , .A( u1_out11_12 ) );
  XOR2_X1 u1_U189 (.B( u1_L10_11 ) , .Z( u1_N362 ) , .A( u1_out11_11 ) );
  XOR2_X1 u1_U19 (.B( u1_L1_21 ) , .Z( u1_N84 ) , .A( u1_out2_21 ) );
  XOR2_X1 u1_U190 (.B( u1_L10_10 ) , .Z( u1_N361 ) , .A( u1_out11_10 ) );
  XOR2_X1 u1_U191 (.B( u1_L10_9 ) , .Z( u1_N360 ) , .A( u1_out11_9 ) );
  XOR2_X1 u1_U192 (.B( u1_L0_5 ) , .Z( u1_N36 ) , .A( u1_out1_5 ) );
  XOR2_X1 u1_U193 (.B( u1_L10_8 ) , .Z( u1_N359 ) , .A( u1_out11_8 ) );
  XOR2_X1 u1_U194 (.B( u1_L10_7 ) , .Z( u1_N358 ) , .A( u1_out11_7 ) );
  XOR2_X1 u1_U195 (.B( u1_L10_6 ) , .Z( u1_N357 ) , .A( u1_out11_6 ) );
  XOR2_X1 u1_U196 (.B( u1_L10_5 ) , .Z( u1_N356 ) , .A( u1_out11_5 ) );
  XOR2_X1 u1_U197 (.B( u1_L10_4 ) , .Z( u1_N355 ) , .A( u1_out11_4 ) );
  XOR2_X1 u1_U198 (.B( u1_L10_3 ) , .Z( u1_N354 ) , .A( u1_out11_3 ) );
  XOR2_X1 u1_U199 (.B( u1_L10_2 ) , .Z( u1_N353 ) , .A( u1_out11_2 ) );
  XOR2_X1 u1_U20 (.B( u1_L1_20 ) , .Z( u1_N83 ) , .A( u1_out2_20 ) );
  XOR2_X1 u1_U200 (.B( u1_L10_1 ) , .Z( u1_N352 ) , .A( u1_out11_1 ) );
  XOR2_X1 u1_U201 (.B( u1_L9_32 ) , .Z( u1_N351 ) , .A( u1_out10_32 ) );
  XOR2_X1 u1_U202 (.B( u1_L9_31 ) , .Z( u1_N350 ) , .A( u1_out10_31 ) );
  XOR2_X1 u1_U203 (.B( u1_L0_4 ) , .Z( u1_N35 ) , .A( u1_out1_4 ) );
  XOR2_X1 u1_U204 (.B( u1_L9_30 ) , .Z( u1_N349 ) , .A( u1_out10_30 ) );
  XOR2_X1 u1_U205 (.B( u1_L9_29 ) , .Z( u1_N348 ) , .A( u1_out10_29 ) );
  XOR2_X1 u1_U206 (.B( u1_L9_28 ) , .Z( u1_N347 ) , .A( u1_out10_28 ) );
  XOR2_X1 u1_U207 (.B( u1_L9_27 ) , .Z( u1_N346 ) , .A( u1_out10_27 ) );
  XOR2_X1 u1_U208 (.B( u1_L9_26 ) , .Z( u1_N345 ) , .A( u1_out10_26 ) );
  XOR2_X1 u1_U209 (.B( u1_L9_25 ) , .Z( u1_N344 ) , .A( u1_out10_25 ) );
  XOR2_X1 u1_U21 (.B( u1_L1_19 ) , .Z( u1_N82 ) , .A( u1_out2_19 ) );
  XOR2_X1 u1_U210 (.B( u1_L9_24 ) , .Z( u1_N343 ) , .A( u1_out10_24 ) );
  XOR2_X1 u1_U211 (.B( u1_L9_23 ) , .Z( u1_N342 ) , .A( u1_out10_23 ) );
  XOR2_X1 u1_U212 (.B( u1_L9_22 ) , .Z( u1_N341 ) , .A( u1_out10_22 ) );
  XOR2_X1 u1_U213 (.B( u1_L9_21 ) , .Z( u1_N340 ) , .A( u1_out10_21 ) );
  XOR2_X1 u1_U214 (.B( u1_L0_3 ) , .Z( u1_N34 ) , .A( u1_out1_3 ) );
  XOR2_X1 u1_U215 (.B( u1_L9_20 ) , .Z( u1_N339 ) , .A( u1_out10_20 ) );
  XOR2_X1 u1_U216 (.B( u1_L9_19 ) , .Z( u1_N338 ) , .A( u1_out10_19 ) );
  XOR2_X1 u1_U217 (.B( u1_L9_18 ) , .Z( u1_N337 ) , .A( u1_out10_18 ) );
  XOR2_X1 u1_U218 (.B( u1_L9_17 ) , .Z( u1_N336 ) , .A( u1_out10_17 ) );
  XOR2_X1 u1_U219 (.B( u1_L9_16 ) , .Z( u1_N335 ) , .A( u1_out10_16 ) );
  XOR2_X1 u1_U22 (.B( u1_L1_18 ) , .Z( u1_N81 ) , .A( u1_out2_18 ) );
  XOR2_X1 u1_U220 (.B( u1_L9_15 ) , .Z( u1_N334 ) , .A( u1_out10_15 ) );
  XOR2_X1 u1_U221 (.B( u1_L9_14 ) , .Z( u1_N333 ) , .A( u1_out10_14 ) );
  XOR2_X1 u1_U222 (.B( u1_L9_13 ) , .Z( u1_N332 ) , .A( u1_out10_13 ) );
  XOR2_X1 u1_U223 (.B( u1_L9_12 ) , .Z( u1_N331 ) , .A( u1_out10_12 ) );
  XOR2_X1 u1_U224 (.B( u1_L9_11 ) , .Z( u1_N330 ) , .A( u1_out10_11 ) );
  XOR2_X1 u1_U225 (.B( u1_L0_2 ) , .Z( u1_N33 ) , .A( u1_out1_2 ) );
  XOR2_X1 u1_U226 (.B( u1_L9_10 ) , .Z( u1_N329 ) , .A( u1_out10_10 ) );
  XOR2_X1 u1_U227 (.B( u1_L9_9 ) , .Z( u1_N328 ) , .A( u1_out10_9 ) );
  XOR2_X1 u1_U228 (.B( u1_L9_8 ) , .Z( u1_N327 ) , .A( u1_out10_8 ) );
  XOR2_X1 u1_U229 (.B( u1_L9_7 ) , .Z( u1_N326 ) , .A( u1_out10_7 ) );
  XOR2_X1 u1_U23 (.B( u1_L1_17 ) , .Z( u1_N80 ) , .A( u1_out2_17 ) );
  XOR2_X1 u1_U230 (.B( u1_L9_6 ) , .Z( u1_N325 ) , .A( u1_out10_6 ) );
  XOR2_X1 u1_U231 (.B( u1_L9_5 ) , .Z( u1_N324 ) , .A( u1_out10_5 ) );
  XOR2_X1 u1_U232 (.B( u1_L9_4 ) , .Z( u1_N323 ) , .A( u1_out10_4 ) );
  XOR2_X1 u1_U233 (.B( u1_L9_3 ) , .Z( u1_N322 ) , .A( u1_out10_3 ) );
  XOR2_X1 u1_U234 (.B( u1_L9_2 ) , .Z( u1_N321 ) , .A( u1_out10_2 ) );
  XOR2_X1 u1_U235 (.B( u1_L9_1 ) , .Z( u1_N320 ) , .A( u1_out10_1 ) );
  XOR2_X1 u1_U236 (.B( u1_L0_1 ) , .Z( u1_N32 ) , .A( u1_out1_1 ) );
  XOR2_X1 u1_U237 (.B( u1_L8_32 ) , .Z( u1_N319 ) , .A( u1_out9_32 ) );
  XOR2_X1 u1_U238 (.B( u1_L8_31 ) , .Z( u1_N318 ) , .A( u1_out9_31 ) );
  XOR2_X1 u1_U239 (.B( u1_L8_30 ) , .Z( u1_N317 ) , .A( u1_out9_30 ) );
  XOR2_X1 u1_U24 (.Z( u1_N8 ) , .B( u1_desIn_r_4 ) , .A( u1_out0_9 ) );
  XOR2_X1 u1_U240 (.B( u1_L8_29 ) , .Z( u1_N316 ) , .A( u1_out9_29 ) );
  XOR2_X1 u1_U241 (.B( u1_L8_28 ) , .Z( u1_N315 ) , .A( u1_out9_28 ) );
  XOR2_X1 u1_U242 (.B( u1_L8_27 ) , .Z( u1_N314 ) , .A( u1_out9_27 ) );
  XOR2_X1 u1_U243 (.B( u1_L8_26 ) , .Z( u1_N313 ) , .A( u1_out9_26 ) );
  XOR2_X1 u1_U244 (.B( u1_L8_25 ) , .Z( u1_N312 ) , .A( u1_out9_25 ) );
  XOR2_X1 u1_U245 (.B( u1_L8_24 ) , .Z( u1_N311 ) , .A( u1_out9_24 ) );
  XOR2_X1 u1_U246 (.B( u1_L8_23 ) , .Z( u1_N310 ) , .A( u1_out9_23 ) );
  XOR2_X1 u1_U247 (.Z( u1_N31 ) , .B( u1_desIn_r_56 ) , .A( u1_out0_32 ) );
  XOR2_X1 u1_U248 (.B( u1_L8_22 ) , .Z( u1_N309 ) , .A( u1_out9_22 ) );
  XOR2_X1 u1_U249 (.B( u1_L8_21 ) , .Z( u1_N308 ) , .A( u1_out9_21 ) );
  XOR2_X1 u1_U25 (.B( u1_L1_16 ) , .Z( u1_N79 ) , .A( u1_out2_16 ) );
  XOR2_X1 u1_U250 (.B( u1_L8_20 ) , .Z( u1_N307 ) , .A( u1_out9_20 ) );
  XOR2_X1 u1_U251 (.B( u1_L8_19 ) , .Z( u1_N306 ) , .A( u1_out9_19 ) );
  XOR2_X1 u1_U252 (.B( u1_L8_18 ) , .Z( u1_N305 ) , .A( u1_out9_18 ) );
  XOR2_X1 u1_U253 (.B( u1_L8_17 ) , .Z( u1_N304 ) , .A( u1_out9_17 ) );
  XOR2_X1 u1_U254 (.B( u1_L8_16 ) , .Z( u1_N303 ) , .A( u1_out9_16 ) );
  XOR2_X1 u1_U255 (.B( u1_L8_15 ) , .Z( u1_N302 ) , .A( u1_out9_15 ) );
  XOR2_X1 u1_U256 (.B( u1_L8_14 ) , .Z( u1_N301 ) , .A( u1_out9_14 ) );
  XOR2_X1 u1_U257 (.B( u1_L8_13 ) , .Z( u1_N300 ) , .A( u1_out9_13 ) );
  XOR2_X1 u1_U258 (.Z( u1_N30 ) , .B( u1_desIn_r_48 ) , .A( u1_out0_31 ) );
  XOR2_X1 u1_U259 (.Z( u1_N3 ) , .B( u1_desIn_r_30 ) , .A( u1_out0_4 ) );
  XOR2_X1 u1_U26 (.B( u1_L1_15 ) , .Z( u1_N78 ) , .A( u1_out2_15 ) );
  XOR2_X1 u1_U260 (.B( u1_L8_12 ) , .Z( u1_N299 ) , .A( u1_out9_12 ) );
  XOR2_X1 u1_U261 (.B( u1_L8_11 ) , .Z( u1_N298 ) , .A( u1_out9_11 ) );
  XOR2_X1 u1_U262 (.B( u1_L8_10 ) , .Z( u1_N297 ) , .A( u1_out9_10 ) );
  XOR2_X1 u1_U263 (.B( u1_L8_9 ) , .Z( u1_N296 ) , .A( u1_out9_9 ) );
  XOR2_X1 u1_U264 (.B( u1_L8_8 ) , .Z( u1_N295 ) , .A( u1_out9_8 ) );
  XOR2_X1 u1_U265 (.B( u1_L8_7 ) , .Z( u1_N294 ) , .A( u1_out9_7 ) );
  XOR2_X1 u1_U266 (.B( u1_L8_6 ) , .Z( u1_N293 ) , .A( u1_out9_6 ) );
  XOR2_X1 u1_U267 (.B( u1_L8_5 ) , .Z( u1_N292 ) , .A( u1_out9_5 ) );
  XOR2_X1 u1_U268 (.B( u1_L8_4 ) , .Z( u1_N291 ) , .A( u1_out9_4 ) );
  XOR2_X1 u1_U269 (.B( u1_L8_3 ) , .Z( u1_N290 ) , .A( u1_out9_3 ) );
  XOR2_X1 u1_U27 (.B( u1_L1_14 ) , .Z( u1_N77 ) , .A( u1_out2_14 ) );
  XOR2_X1 u1_U270 (.Z( u1_N29 ) , .B( u1_desIn_r_40 ) , .A( u1_out0_30 ) );
  XOR2_X1 u1_U271 (.B( u1_L8_2 ) , .Z( u1_N289 ) , .A( u1_out9_2 ) );
  XOR2_X1 u1_U272 (.B( u1_L8_1 ) , .Z( u1_N288 ) , .A( u1_out9_1 ) );
  XOR2_X1 u1_U273 (.B( u1_L7_32 ) , .Z( u1_N287 ) , .A( u1_out8_32 ) );
  XOR2_X1 u1_U274 (.B( u1_L7_31 ) , .Z( u1_N286 ) , .A( u1_out8_31 ) );
  XOR2_X1 u1_U275 (.B( u1_L7_30 ) , .Z( u1_N285 ) , .A( u1_out8_30 ) );
  XOR2_X1 u1_U276 (.B( u1_L7_29 ) , .Z( u1_N284 ) , .A( u1_out8_29 ) );
  XOR2_X1 u1_U277 (.B( u1_L7_28 ) , .Z( u1_N283 ) , .A( u1_out8_28 ) );
  XOR2_X1 u1_U278 (.B( u1_L7_27 ) , .Z( u1_N282 ) , .A( u1_out8_27 ) );
  XOR2_X1 u1_U279 (.B( u1_L7_26 ) , .Z( u1_N281 ) , .A( u1_out8_26 ) );
  XOR2_X1 u1_U28 (.B( u1_L1_13 ) , .Z( u1_N76 ) , .A( u1_out2_13 ) );
  XOR2_X1 u1_U280 (.B( u1_L7_25 ) , .Z( u1_N280 ) , .A( u1_out8_25 ) );
  XOR2_X1 u1_U281 (.Z( u1_N28 ) , .B( u1_desIn_r_32 ) , .A( u1_out0_29 ) );
  XOR2_X1 u1_U282 (.B( u1_L7_24 ) , .Z( u1_N279 ) , .A( u1_out8_24 ) );
  XOR2_X1 u1_U283 (.B( u1_L7_23 ) , .Z( u1_N278 ) , .A( u1_out8_23 ) );
  XOR2_X1 u1_U284 (.B( u1_L7_22 ) , .Z( u1_N277 ) , .A( u1_out8_22 ) );
  XOR2_X1 u1_U285 (.B( u1_L7_21 ) , .Z( u1_N276 ) , .A( u1_out8_21 ) );
  XOR2_X1 u1_U286 (.B( u1_L7_20 ) , .Z( u1_N275 ) , .A( u1_out8_20 ) );
  XOR2_X1 u1_U287 (.B( u1_L7_19 ) , .Z( u1_N274 ) , .A( u1_out8_19 ) );
  XOR2_X1 u1_U288 (.B( u1_L7_18 ) , .Z( u1_N273 ) , .A( u1_out8_18 ) );
  XOR2_X1 u1_U289 (.B( u1_L7_17 ) , .Z( u1_N272 ) , .A( u1_out8_17 ) );
  XOR2_X1 u1_U29 (.B( u1_L1_12 ) , .Z( u1_N75 ) , .A( u1_out2_12 ) );
  XOR2_X1 u1_U290 (.B( u1_L7_16 ) , .Z( u1_N271 ) , .A( u1_out8_16 ) );
  XOR2_X1 u1_U291 (.B( u1_L7_15 ) , .Z( u1_N270 ) , .A( u1_out8_15 ) );
  XOR2_X1 u1_U292 (.Z( u1_N27 ) , .B( u1_desIn_r_24 ) , .A( u1_out0_28 ) );
  XOR2_X1 u1_U293 (.B( u1_L7_14 ) , .Z( u1_N269 ) , .A( u1_out8_14 ) );
  XOR2_X1 u1_U294 (.B( u1_L7_13 ) , .Z( u1_N268 ) , .A( u1_out8_13 ) );
  XOR2_X1 u1_U295 (.B( u1_L7_12 ) , .Z( u1_N267 ) , .A( u1_out8_12 ) );
  XOR2_X1 u1_U296 (.B( u1_L7_11 ) , .Z( u1_N266 ) , .A( u1_out8_11 ) );
  XOR2_X1 u1_U297 (.B( u1_L7_10 ) , .Z( u1_N265 ) , .A( u1_out8_10 ) );
  XOR2_X1 u1_U298 (.B( u1_L7_9 ) , .Z( u1_N264 ) , .A( u1_out8_9 ) );
  XOR2_X1 u1_U299 (.B( u1_L7_8 ) , .Z( u1_N263 ) , .A( u1_out8_8 ) );
  XOR2_X1 u1_U3 (.B( u1_L2_4 ) , .Z( u1_N99 ) , .A( u1_out3_4 ) );
  XOR2_X1 u1_U30 (.B( u1_L1_11 ) , .Z( u1_N74 ) , .A( u1_out2_11 ) );
  XOR2_X1 u1_U300 (.B( u1_L7_7 ) , .Z( u1_N262 ) , .A( u1_out8_7 ) );
  XOR2_X1 u1_U301 (.B( u1_L7_6 ) , .Z( u1_N261 ) , .A( u1_out8_6 ) );
  XOR2_X1 u1_U302 (.B( u1_L7_5 ) , .Z( u1_N260 ) , .A( u1_out8_5 ) );
  XOR2_X1 u1_U303 (.Z( u1_N26 ) , .B( u1_desIn_r_16 ) , .A( u1_out0_27 ) );
  XOR2_X1 u1_U304 (.B( u1_L7_4 ) , .Z( u1_N259 ) , .A( u1_out8_4 ) );
  XOR2_X1 u1_U305 (.B( u1_L7_3 ) , .Z( u1_N258 ) , .A( u1_out8_3 ) );
  XOR2_X1 u1_U306 (.B( u1_L7_2 ) , .Z( u1_N257 ) , .A( u1_out8_2 ) );
  XOR2_X1 u1_U307 (.B( u1_L7_1 ) , .Z( u1_N256 ) , .A( u1_out8_1 ) );
  XOR2_X1 u1_U308 (.B( u1_L6_32 ) , .Z( u1_N255 ) , .A( u1_out7_32 ) );
  XOR2_X1 u1_U309 (.B( u1_L6_31 ) , .Z( u1_N254 ) , .A( u1_out7_31 ) );
  XOR2_X1 u1_U31 (.B( u1_L1_10 ) , .Z( u1_N73 ) , .A( u1_out2_10 ) );
  XOR2_X1 u1_U310 (.B( u1_L6_30 ) , .Z( u1_N253 ) , .A( u1_out7_30 ) );
  XOR2_X1 u1_U311 (.B( u1_L6_29 ) , .Z( u1_N252 ) , .A( u1_out7_29 ) );
  XOR2_X1 u1_U312 (.B( u1_L6_28 ) , .Z( u1_N251 ) , .A( u1_out7_28 ) );
  XOR2_X1 u1_U313 (.B( u1_L6_27 ) , .Z( u1_N250 ) , .A( u1_out7_27 ) );
  XOR2_X1 u1_U314 (.Z( u1_N25 ) , .B( u1_desIn_r_8 ) , .A( u1_out0_26 ) );
  XOR2_X1 u1_U315 (.B( u1_L6_26 ) , .Z( u1_N249 ) , .A( u1_out7_26 ) );
  XOR2_X1 u1_U316 (.B( u1_L6_25 ) , .Z( u1_N248 ) , .A( u1_out7_25 ) );
  XOR2_X1 u1_U317 (.B( u1_L6_24 ) , .Z( u1_N247 ) , .A( u1_out7_24 ) );
  XOR2_X1 u1_U318 (.B( u1_L6_23 ) , .Z( u1_N246 ) , .A( u1_out7_23 ) );
  XOR2_X1 u1_U319 (.B( u1_L6_22 ) , .Z( u1_N245 ) , .A( u1_out7_22 ) );
  XOR2_X1 u1_U32 (.B( u1_L1_9 ) , .Z( u1_N72 ) , .A( u1_out2_9 ) );
  XOR2_X1 u1_U320 (.B( u1_L6_21 ) , .Z( u1_N244 ) , .A( u1_out7_21 ) );
  XOR2_X1 u1_U321 (.B( u1_L6_20 ) , .Z( u1_N243 ) , .A( u1_out7_20 ) );
  XOR2_X1 u1_U322 (.B( u1_L6_19 ) , .Z( u1_N242 ) , .A( u1_out7_19 ) );
  XOR2_X1 u1_U323 (.B( u1_L6_18 ) , .Z( u1_N241 ) , .A( u1_out7_18 ) );
  XOR2_X1 u1_U324 (.B( u1_L6_17 ) , .Z( u1_N240 ) , .A( u1_out7_17 ) );
  XOR2_X1 u1_U325 (.Z( u1_N24 ) , .B( u1_desIn_r_0 ) , .A( u1_out0_25 ) );
  XOR2_X1 u1_U326 (.B( u1_L6_16 ) , .Z( u1_N239 ) , .A( u1_out7_16 ) );
  XOR2_X1 u1_U327 (.B( u1_L6_15 ) , .Z( u1_N238 ) , .A( u1_out7_15 ) );
  XOR2_X1 u1_U328 (.B( u1_L6_14 ) , .Z( u1_N237 ) , .A( u1_out7_14 ) );
  XOR2_X1 u1_U329 (.B( u1_L6_13 ) , .Z( u1_N236 ) , .A( u1_out7_13 ) );
  XOR2_X1 u1_U33 (.B( u1_L1_8 ) , .Z( u1_N71 ) , .A( u1_out2_8 ) );
  XOR2_X1 u1_U330 (.B( u1_L6_12 ) , .Z( u1_N235 ) , .A( u1_out7_12 ) );
  XOR2_X1 u1_U331 (.B( u1_L6_11 ) , .Z( u1_N234 ) , .A( u1_out7_11 ) );
  XOR2_X1 u1_U332 (.B( u1_L6_10 ) , .Z( u1_N233 ) , .A( u1_out7_10 ) );
  XOR2_X1 u1_U333 (.B( u1_L6_9 ) , .Z( u1_N232 ) , .A( u1_out7_9 ) );
  XOR2_X1 u1_U334 (.B( u1_L6_8 ) , .Z( u1_N231 ) , .A( u1_out7_8 ) );
  XOR2_X1 u1_U335 (.B( u1_L6_7 ) , .Z( u1_N230 ) , .A( u1_out7_7 ) );
  XOR2_X1 u1_U336 (.Z( u1_N23 ) , .B( u1_desIn_r_58 ) , .A( u1_out0_24 ) );
  XOR2_X1 u1_U337 (.B( u1_L6_6 ) , .Z( u1_N229 ) , .A( u1_out7_6 ) );
  XOR2_X1 u1_U338 (.B( u1_L6_5 ) , .Z( u1_N228 ) , .A( u1_out7_5 ) );
  XOR2_X1 u1_U339 (.B( u1_L6_4 ) , .Z( u1_N227 ) , .A( u1_out7_4 ) );
  XOR2_X1 u1_U34 (.B( u1_L1_7 ) , .Z( u1_N70 ) , .A( u1_out2_7 ) );
  XOR2_X1 u1_U340 (.B( u1_L6_3 ) , .Z( u1_N226 ) , .A( u1_out7_3 ) );
  XOR2_X1 u1_U341 (.B( u1_L6_2 ) , .Z( u1_N225 ) , .A( u1_out7_2 ) );
  XOR2_X1 u1_U342 (.B( u1_L6_1 ) , .Z( u1_N224 ) , .A( u1_out7_1 ) );
  XOR2_X1 u1_U343 (.B( u1_L5_32 ) , .Z( u1_N223 ) , .A( u1_out6_32 ) );
  XOR2_X1 u1_U344 (.B( u1_L5_31 ) , .Z( u1_N222 ) , .A( u1_out6_31 ) );
  XOR2_X1 u1_U345 (.B( u1_L5_30 ) , .Z( u1_N221 ) , .A( u1_out6_30 ) );
  XOR2_X1 u1_U346 (.B( u1_L5_29 ) , .Z( u1_N220 ) , .A( u1_out6_29 ) );
  XOR2_X1 u1_U347 (.Z( u1_N22 ) , .B( u1_desIn_r_50 ) , .A( u1_out0_23 ) );
  XOR2_X1 u1_U348 (.B( u1_L5_28 ) , .Z( u1_N219 ) , .A( u1_out6_28 ) );
  XOR2_X1 u1_U349 (.B( u1_L5_27 ) , .Z( u1_N218 ) , .A( u1_out6_27 ) );
  XOR2_X1 u1_U35 (.Z( u1_N7 ) , .B( u1_desIn_r_62 ) , .A( u1_out0_8 ) );
  XOR2_X1 u1_U350 (.B( u1_L5_26 ) , .Z( u1_N217 ) , .A( u1_out6_26 ) );
  XOR2_X1 u1_U351 (.B( u1_L5_25 ) , .Z( u1_N216 ) , .A( u1_out6_25 ) );
  XOR2_X1 u1_U352 (.B( u1_L5_24 ) , .Z( u1_N215 ) , .A( u1_out6_24 ) );
  XOR2_X1 u1_U353 (.B( u1_L5_23 ) , .Z( u1_N214 ) , .A( u1_out6_23 ) );
  XOR2_X1 u1_U354 (.B( u1_L5_22 ) , .Z( u1_N213 ) , .A( u1_out6_22 ) );
  XOR2_X1 u1_U355 (.B( u1_L5_21 ) , .Z( u1_N212 ) , .A( u1_out6_21 ) );
  XOR2_X1 u1_U356 (.B( u1_L5_20 ) , .Z( u1_N211 ) , .A( u1_out6_20 ) );
  XOR2_X1 u1_U357 (.B( u1_L5_19 ) , .Z( u1_N210 ) , .A( u1_out6_19 ) );
  XOR2_X1 u1_U358 (.Z( u1_N21 ) , .B( u1_desIn_r_42 ) , .A( u1_out0_22 ) );
  XOR2_X1 u1_U359 (.B( u1_L5_18 ) , .Z( u1_N209 ) , .A( u1_out6_18 ) );
  XOR2_X1 u1_U36 (.B( u1_L1_6 ) , .Z( u1_N69 ) , .A( u1_out2_6 ) );
  XOR2_X1 u1_U360 (.B( u1_L5_17 ) , .Z( u1_N208 ) , .A( u1_out6_17 ) );
  XOR2_X1 u1_U361 (.B( u1_L5_16 ) , .Z( u1_N207 ) , .A( u1_out6_16 ) );
  XOR2_X1 u1_U362 (.B( u1_L5_15 ) , .Z( u1_N206 ) , .A( u1_out6_15 ) );
  XOR2_X1 u1_U363 (.B( u1_L5_14 ) , .Z( u1_N205 ) , .A( u1_out6_14 ) );
  XOR2_X1 u1_U364 (.B( u1_L5_13 ) , .Z( u1_N204 ) , .A( u1_out6_13 ) );
  XOR2_X1 u1_U365 (.B( u1_L5_12 ) , .Z( u1_N203 ) , .A( u1_out6_12 ) );
  XOR2_X1 u1_U366 (.B( u1_L5_11 ) , .Z( u1_N202 ) , .A( u1_out6_11 ) );
  XOR2_X1 u1_U367 (.B( u1_L5_10 ) , .Z( u1_N201 ) , .A( u1_out6_10 ) );
  XOR2_X1 u1_U368 (.B( u1_L5_9 ) , .Z( u1_N200 ) , .A( u1_out6_9 ) );
  XOR2_X1 u1_U369 (.Z( u1_N20 ) , .B( u1_desIn_r_34 ) , .A( u1_out0_21 ) );
  XOR2_X1 u1_U37 (.B( u1_L1_5 ) , .Z( u1_N68 ) , .A( u1_out2_5 ) );
  XOR2_X1 u1_U370 (.Z( u1_N2 ) , .B( u1_desIn_r_22 ) , .A( u1_out0_3 ) );
  XOR2_X1 u1_U371 (.B( u1_L5_8 ) , .Z( u1_N199 ) , .A( u1_out6_8 ) );
  XOR2_X1 u1_U372 (.B( u1_L5_7 ) , .Z( u1_N198 ) , .A( u1_out6_7 ) );
  XOR2_X1 u1_U373 (.B( u1_L5_6 ) , .Z( u1_N197 ) , .A( u1_out6_6 ) );
  XOR2_X1 u1_U374 (.B( u1_L5_5 ) , .Z( u1_N196 ) , .A( u1_out6_5 ) );
  XOR2_X1 u1_U375 (.B( u1_L5_4 ) , .Z( u1_N195 ) , .A( u1_out6_4 ) );
  XOR2_X1 u1_U376 (.B( u1_L5_3 ) , .Z( u1_N194 ) , .A( u1_out6_3 ) );
  XOR2_X1 u1_U377 (.B( u1_L5_2 ) , .Z( u1_N193 ) , .A( u1_out6_2 ) );
  XOR2_X1 u1_U378 (.B( u1_L5_1 ) , .Z( u1_N192 ) , .A( u1_out6_1 ) );
  XOR2_X1 u1_U379 (.B( u1_L4_32 ) , .Z( u1_N191 ) , .A( u1_out5_32 ) );
  XOR2_X1 u1_U38 (.B( u1_L1_4 ) , .Z( u1_N67 ) , .A( u1_out2_4 ) );
  XOR2_X1 u1_U380 (.B( u1_L4_31 ) , .Z( u1_N190 ) , .A( u1_out5_31 ) );
  XOR2_X1 u1_U381 (.Z( u1_N19 ) , .B( u1_desIn_r_26 ) , .A( u1_out0_20 ) );
  XOR2_X1 u1_U382 (.B( u1_L4_30 ) , .Z( u1_N189 ) , .A( u1_out5_30 ) );
  XOR2_X1 u1_U383 (.B( u1_L4_29 ) , .Z( u1_N188 ) , .A( u1_out5_29 ) );
  XOR2_X1 u1_U384 (.B( u1_L4_28 ) , .Z( u1_N187 ) , .A( u1_out5_28 ) );
  XOR2_X1 u1_U385 (.B( u1_L4_27 ) , .Z( u1_N186 ) , .A( u1_out5_27 ) );
  XOR2_X1 u1_U386 (.B( u1_L4_26 ) , .Z( u1_N185 ) , .A( u1_out5_26 ) );
  XOR2_X1 u1_U387 (.B( u1_L4_25 ) , .Z( u1_N184 ) , .A( u1_out5_25 ) );
  XOR2_X1 u1_U388 (.B( u1_L4_24 ) , .Z( u1_N183 ) , .A( u1_out5_24 ) );
  XOR2_X1 u1_U389 (.B( u1_L4_23 ) , .Z( u1_N182 ) , .A( u1_out5_23 ) );
  XOR2_X1 u1_U39 (.B( u1_L1_3 ) , .Z( u1_N66 ) , .A( u1_out2_3 ) );
  XOR2_X1 u1_U390 (.B( u1_L4_22 ) , .Z( u1_N181 ) , .A( u1_out5_22 ) );
  XOR2_X1 u1_U391 (.B( u1_L4_21 ) , .Z( u1_N180 ) , .A( u1_out5_21 ) );
  XOR2_X1 u1_U392 (.Z( u1_N18 ) , .B( u1_desIn_r_18 ) , .A( u1_out0_19 ) );
  XOR2_X1 u1_U393 (.B( u1_L4_20 ) , .Z( u1_N179 ) , .A( u1_out5_20 ) );
  XOR2_X1 u1_U394 (.B( u1_L4_19 ) , .Z( u1_N178 ) , .A( u1_out5_19 ) );
  XOR2_X1 u1_U395 (.B( u1_L4_18 ) , .Z( u1_N177 ) , .A( u1_out5_18 ) );
  XOR2_X1 u1_U396 (.B( u1_L4_17 ) , .Z( u1_N176 ) , .A( u1_out5_17 ) );
  XOR2_X1 u1_U397 (.B( u1_L4_16 ) , .Z( u1_N175 ) , .A( u1_out5_16 ) );
  XOR2_X1 u1_U398 (.B( u1_L4_15 ) , .Z( u1_N174 ) , .A( u1_out5_15 ) );
  XOR2_X1 u1_U399 (.B( u1_L4_14 ) , .Z( u1_N173 ) , .A( u1_out5_14 ) );
  XOR2_X1 u1_U4 (.B( u1_L2_3 ) , .Z( u1_N98 ) , .A( u1_out3_3 ) );
  XOR2_X1 u1_U40 (.B( u1_L1_2 ) , .Z( u1_N65 ) , .A( u1_out2_2 ) );
  XOR2_X1 u1_U400 (.B( u1_L4_13 ) , .Z( u1_N172 ) , .A( u1_out5_13 ) );
  XOR2_X1 u1_U401 (.B( u1_L4_12 ) , .Z( u1_N171 ) , .A( u1_out5_12 ) );
  XOR2_X1 u1_U402 (.B( u1_L4_11 ) , .Z( u1_N170 ) , .A( u1_out5_11 ) );
  XOR2_X1 u1_U403 (.Z( u1_N17 ) , .B( u1_desIn_r_10 ) , .A( u1_out0_18 ) );
  XOR2_X1 u1_U404 (.B( u1_L4_10 ) , .Z( u1_N169 ) , .A( u1_out5_10 ) );
  XOR2_X1 u1_U405 (.B( u1_L4_9 ) , .Z( u1_N168 ) , .A( u1_out5_9 ) );
  XOR2_X1 u1_U406 (.B( u1_L4_8 ) , .Z( u1_N167 ) , .A( u1_out5_8 ) );
  XOR2_X1 u1_U407 (.B( u1_L4_7 ) , .Z( u1_N166 ) , .A( u1_out5_7 ) );
  XOR2_X1 u1_U408 (.B( u1_L4_6 ) , .Z( u1_N165 ) , .A( u1_out5_6 ) );
  XOR2_X1 u1_U409 (.B( u1_L4_5 ) , .Z( u1_N164 ) , .A( u1_out5_5 ) );
  XOR2_X1 u1_U41 (.B( u1_L1_1 ) , .Z( u1_N64 ) , .A( u1_out2_1 ) );
  XOR2_X1 u1_U410 (.B( u1_L4_4 ) , .Z( u1_N163 ) , .A( u1_out5_4 ) );
  XOR2_X1 u1_U411 (.B( u1_L4_3 ) , .Z( u1_N162 ) , .A( u1_out5_3 ) );
  XOR2_X1 u1_U412 (.B( u1_L4_2 ) , .Z( u1_N161 ) , .A( u1_out5_2 ) );
  XOR2_X1 u1_U413 (.B( u1_L4_1 ) , .Z( u1_N160 ) , .A( u1_out5_1 ) );
  XOR2_X1 u1_U414 (.Z( u1_N16 ) , .B( u1_desIn_r_2 ) , .A( u1_out0_17 ) );
  XOR2_X1 u1_U415 (.B( u1_L3_32 ) , .Z( u1_N159 ) , .A( u1_out4_32 ) );
  XOR2_X1 u1_U416 (.B( u1_L3_31 ) , .Z( u1_N158 ) , .A( u1_out4_31 ) );
  XOR2_X1 u1_U417 (.B( u1_L3_30 ) , .Z( u1_N157 ) , .A( u1_out4_30 ) );
  XOR2_X1 u1_U418 (.B( u1_L3_29 ) , .Z( u1_N156 ) , .A( u1_out4_29 ) );
  XOR2_X1 u1_U419 (.B( u1_L3_28 ) , .Z( u1_N155 ) , .A( u1_out4_28 ) );
  XOR2_X1 u1_U42 (.B( u1_L0_32 ) , .Z( u1_N63 ) , .A( u1_out1_32 ) );
  XOR2_X1 u1_U420 (.B( u1_L3_27 ) , .Z( u1_N154 ) , .A( u1_out4_27 ) );
  XOR2_X1 u1_U421 (.B( u1_L3_26 ) , .Z( u1_N153 ) , .A( u1_out4_26 ) );
  XOR2_X1 u1_U422 (.B( u1_L3_25 ) , .Z( u1_N152 ) , .A( u1_out4_25 ) );
  XOR2_X1 u1_U423 (.B( u1_L3_24 ) , .Z( u1_N151 ) , .A( u1_out4_24 ) );
  XOR2_X1 u1_U424 (.B( u1_L3_23 ) , .Z( u1_N150 ) , .A( u1_out4_23 ) );
  XOR2_X1 u1_U425 (.Z( u1_N15 ) , .B( u1_desIn_r_60 ) , .A( u1_out0_16 ) );
  XOR2_X1 u1_U426 (.B( u1_L3_22 ) , .Z( u1_N149 ) , .A( u1_out4_22 ) );
  XOR2_X1 u1_U427 (.B( u1_L3_21 ) , .Z( u1_N148 ) , .A( u1_out4_21 ) );
  XOR2_X1 u1_U428 (.B( u1_L3_20 ) , .Z( u1_N147 ) , .A( u1_out4_20 ) );
  XOR2_X1 u1_U429 (.B( u1_L3_19 ) , .Z( u1_N146 ) , .A( u1_out4_19 ) );
  XOR2_X1 u1_U43 (.B( u1_L0_31 ) , .Z( u1_N62 ) , .A( u1_out1_31 ) );
  XOR2_X1 u1_U430 (.B( u1_L3_18 ) , .Z( u1_N145 ) , .A( u1_out4_18 ) );
  XOR2_X1 u1_U431 (.B( u1_L3_17 ) , .Z( u1_N144 ) , .A( u1_out4_17 ) );
  XOR2_X1 u1_U432 (.B( u1_L3_16 ) , .Z( u1_N143 ) , .A( u1_out4_16 ) );
  XOR2_X1 u1_U433 (.B( u1_L3_15 ) , .Z( u1_N142 ) , .A( u1_out4_15 ) );
  XOR2_X1 u1_U434 (.B( u1_L3_14 ) , .Z( u1_N141 ) , .A( u1_out4_14 ) );
  XOR2_X1 u1_U435 (.B( u1_L3_13 ) , .Z( u1_N140 ) , .A( u1_out4_13 ) );
  XOR2_X1 u1_U436 (.Z( u1_N14 ) , .B( u1_desIn_r_52 ) , .A( u1_out0_15 ) );
  XOR2_X1 u1_U437 (.B( u1_L3_12 ) , .Z( u1_N139 ) , .A( u1_out4_12 ) );
  XOR2_X1 u1_U438 (.B( u1_L3_11 ) , .Z( u1_N138 ) , .A( u1_out4_11 ) );
  XOR2_X1 u1_U439 (.B( u1_L3_10 ) , .Z( u1_N137 ) , .A( u1_out4_10 ) );
  XOR2_X1 u1_U44 (.B( u1_L0_30 ) , .Z( u1_N61 ) , .A( u1_out1_30 ) );
  XOR2_X1 u1_U440 (.B( u1_L3_9 ) , .Z( u1_N136 ) , .A( u1_out4_9 ) );
  XOR2_X1 u1_U441 (.B( u1_L3_8 ) , .Z( u1_N135 ) , .A( u1_out4_8 ) );
  XOR2_X1 u1_U442 (.B( u1_L3_7 ) , .Z( u1_N134 ) , .A( u1_out4_7 ) );
  XOR2_X1 u1_U443 (.B( u1_L3_6 ) , .Z( u1_N133 ) , .A( u1_out4_6 ) );
  XOR2_X1 u1_U444 (.B( u1_L3_5 ) , .Z( u1_N132 ) , .A( u1_out4_5 ) );
  XOR2_X1 u1_U445 (.B( u1_L3_4 ) , .Z( u1_N131 ) , .A( u1_out4_4 ) );
  XOR2_X1 u1_U446 (.B( u1_L3_3 ) , .Z( u1_N130 ) , .A( u1_out4_3 ) );
  XOR2_X1 u1_U447 (.Z( u1_N13 ) , .B( u1_desIn_r_44 ) , .A( u1_out0_14 ) );
  XOR2_X1 u1_U448 (.B( u1_L3_2 ) , .Z( u1_N129 ) , .A( u1_out4_2 ) );
  XOR2_X1 u1_U449 (.B( u1_L3_1 ) , .Z( u1_N128 ) , .A( u1_out4_1 ) );
  XOR2_X1 u1_U45 (.B( u1_L0_29 ) , .Z( u1_N60 ) , .A( u1_out1_29 ) );
  XOR2_X1 u1_U450 (.B( u1_L2_32 ) , .Z( u1_N127 ) , .A( u1_out3_32 ) );
  XOR2_X1 u1_U451 (.B( u1_L2_31 ) , .Z( u1_N126 ) , .A( u1_out3_31 ) );
  XOR2_X1 u1_U452 (.B( u1_L2_30 ) , .Z( u1_N125 ) , .A( u1_out3_30 ) );
  XOR2_X1 u1_U453 (.B( u1_L2_29 ) , .Z( u1_N124 ) , .A( u1_out3_29 ) );
  XOR2_X1 u1_U454 (.B( u1_L2_28 ) , .Z( u1_N123 ) , .A( u1_out3_28 ) );
  XOR2_X1 u1_U455 (.B( u1_L2_27 ) , .Z( u1_N122 ) , .A( u1_out3_27 ) );
  XOR2_X1 u1_U456 (.B( u1_L2_26 ) , .Z( u1_N121 ) , .A( u1_out3_26 ) );
  XOR2_X1 u1_U457 (.B( u1_L2_25 ) , .Z( u1_N120 ) , .A( u1_out3_25 ) );
  XOR2_X1 u1_U458 (.Z( u1_N12 ) , .B( u1_desIn_r_36 ) , .A( u1_out0_13 ) );
  XOR2_X1 u1_U459 (.B( u1_L2_24 ) , .Z( u1_N119 ) , .A( u1_out3_24 ) );
  XOR2_X1 u1_U46 (.Z( u1_N6 ) , .B( u1_desIn_r_54 ) , .A( u1_out0_7 ) );
  XOR2_X1 u1_U460 (.B( u1_L2_23 ) , .Z( u1_N118 ) , .A( u1_out3_23 ) );
  XOR2_X1 u1_U461 (.B( u1_L2_22 ) , .Z( u1_N117 ) , .A( u1_out3_22 ) );
  XOR2_X1 u1_U462 (.B( u1_L2_21 ) , .Z( u1_N116 ) , .A( u1_out3_21 ) );
  XOR2_X1 u1_U463 (.B( u1_L2_20 ) , .Z( u1_N115 ) , .A( u1_out3_20 ) );
  XOR2_X1 u1_U464 (.B( u1_L2_19 ) , .Z( u1_N114 ) , .A( u1_out3_19 ) );
  XOR2_X1 u1_U465 (.B( u1_L2_18 ) , .Z( u1_N113 ) , .A( u1_out3_18 ) );
  XOR2_X1 u1_U466 (.B( u1_L2_17 ) , .Z( u1_N112 ) , .A( u1_out3_17 ) );
  XOR2_X1 u1_U467 (.B( u1_L2_16 ) , .Z( u1_N111 ) , .A( u1_out3_16 ) );
  XOR2_X1 u1_U468 (.B( u1_L2_15 ) , .Z( u1_N110 ) , .A( u1_out3_15 ) );
  XOR2_X1 u1_U469 (.Z( u1_N11 ) , .B( u1_desIn_r_28 ) , .A( u1_out0_12 ) );
  XOR2_X1 u1_U47 (.B( u1_L0_28 ) , .Z( u1_N59 ) , .A( u1_out1_28 ) );
  XOR2_X1 u1_U470 (.B( u1_L2_14 ) , .Z( u1_N109 ) , .A( u1_out3_14 ) );
  XOR2_X1 u1_U471 (.B( u1_L2_13 ) , .Z( u1_N108 ) , .A( u1_out3_13 ) );
  XOR2_X1 u1_U472 (.B( u1_L2_12 ) , .Z( u1_N107 ) , .A( u1_out3_12 ) );
  XOR2_X1 u1_U473 (.B( u1_L2_11 ) , .Z( u1_N106 ) , .A( u1_out3_11 ) );
  XOR2_X1 u1_U474 (.B( u1_L2_10 ) , .Z( u1_N105 ) , .A( u1_out3_10 ) );
  XOR2_X1 u1_U475 (.B( u1_L2_9 ) , .Z( u1_N104 ) , .A( u1_out3_9 ) );
  XOR2_X1 u1_U476 (.B( u1_L2_8 ) , .Z( u1_N103 ) , .A( u1_out3_8 ) );
  XOR2_X1 u1_U477 (.B( u1_L2_7 ) , .Z( u1_N102 ) , .A( u1_out3_7 ) );
  XOR2_X1 u1_U478 (.B( u1_L2_6 ) , .Z( u1_N101 ) , .A( u1_out3_6 ) );
  XOR2_X1 u1_U479 (.B( u1_L2_5 ) , .Z( u1_N100 ) , .A( u1_out3_5 ) );
  XOR2_X1 u1_U48 (.B( u1_L0_27 ) , .Z( u1_N58 ) , .A( u1_out1_27 ) );
  XOR2_X1 u1_U480 (.Z( u1_N10 ) , .B( u1_desIn_r_20 ) , .A( u1_out0_11 ) );
  XOR2_X1 u1_U481 (.Z( u1_N1 ) , .B( u1_desIn_r_14 ) , .A( u1_out0_2 ) );
  XOR2_X1 u1_U482 (.Z( u1_N0 ) , .B( u1_desIn_r_6 ) , .A( u1_out0_1 ) );
  XOR2_X1 u1_U483 (.Z( u1_FP_9 ) , .B( u1_L14_9 ) , .A( u1_out15_9 ) );
  XOR2_X1 u1_U484 (.Z( u1_FP_8 ) , .B( u1_L14_8 ) , .A( u1_out15_8 ) );
  XOR2_X1 u1_U485 (.Z( u1_FP_7 ) , .B( u1_L14_7 ) , .A( u1_out15_7 ) );
  XOR2_X1 u1_U486 (.Z( u1_FP_6 ) , .B( u1_L14_6 ) , .A( u1_out15_6 ) );
  XOR2_X1 u1_U487 (.Z( u1_FP_5 ) , .B( u1_L14_5 ) , .A( u1_out15_5 ) );
  XOR2_X1 u1_U488 (.Z( u1_FP_4 ) , .B( u1_L14_4 ) , .A( u1_out15_4 ) );
  XOR2_X1 u1_U489 (.Z( u1_FP_3 ) , .B( u1_L14_3 ) , .A( u1_out15_3 ) );
  XOR2_X1 u1_U49 (.B( u1_L0_26 ) , .Z( u1_N57 ) , .A( u1_out1_26 ) );
  XOR2_X1 u1_U490 (.Z( u1_FP_32 ) , .B( u1_L14_32 ) , .A( u1_out15_32 ) );
  XOR2_X1 u1_U491 (.Z( u1_FP_31 ) , .B( u1_L14_31 ) , .A( u1_out15_31 ) );
  XOR2_X1 u1_U492 (.Z( u1_FP_30 ) , .B( u1_L14_30 ) , .A( u1_out15_30 ) );
  XOR2_X1 u1_U493 (.Z( u1_FP_2 ) , .B( u1_L14_2 ) , .A( u1_out15_2 ) );
  XOR2_X1 u1_U494 (.Z( u1_FP_29 ) , .B( u1_L14_29 ) , .A( u1_out15_29 ) );
  XOR2_X1 u1_U495 (.Z( u1_FP_28 ) , .B( u1_L14_28 ) , .A( u1_out15_28 ) );
  XOR2_X1 u1_U496 (.Z( u1_FP_27 ) , .B( u1_L14_27 ) , .A( u1_out15_27 ) );
  XOR2_X1 u1_U497 (.Z( u1_FP_26 ) , .B( u1_L14_26 ) , .A( u1_out15_26 ) );
  XOR2_X1 u1_U498 (.Z( u1_FP_25 ) , .B( u1_L14_25 ) , .A( u1_out15_25 ) );
  XOR2_X1 u1_U499 (.Z( u1_FP_24 ) , .B( u1_L14_24 ) , .A( u1_out15_24 ) );
  XOR2_X1 u1_U5 (.B( u1_L2_2 ) , .Z( u1_N97 ) , .A( u1_out3_2 ) );
  XOR2_X1 u1_U50 (.B( u1_L0_25 ) , .Z( u1_N56 ) , .A( u1_out1_25 ) );
  XOR2_X1 u1_U500 (.Z( u1_FP_23 ) , .B( u1_L14_23 ) , .A( u1_out15_23 ) );
  XOR2_X1 u1_U501 (.Z( u1_FP_22 ) , .B( u1_L14_22 ) , .A( u1_out15_22 ) );
  XOR2_X1 u1_U502 (.Z( u1_FP_21 ) , .B( u1_L14_21 ) , .A( u1_out15_21 ) );
  XOR2_X1 u1_U503 (.Z( u1_FP_20 ) , .B( u1_L14_20 ) , .A( u1_out15_20 ) );
  XOR2_X1 u1_U504 (.Z( u1_FP_1 ) , .B( u1_L14_1 ) , .A( u1_out15_1 ) );
  XOR2_X1 u1_U505 (.Z( u1_FP_19 ) , .B( u1_L14_19 ) , .A( u1_out15_19 ) );
  XOR2_X1 u1_U506 (.Z( u1_FP_18 ) , .B( u1_L14_18 ) , .A( u1_out15_18 ) );
  XOR2_X1 u1_U507 (.Z( u1_FP_17 ) , .B( u1_L14_17 ) , .A( u1_out15_17 ) );
  XOR2_X1 u1_U508 (.Z( u1_FP_16 ) , .B( u1_L14_16 ) , .A( u1_out15_16 ) );
  XOR2_X1 u1_U509 (.Z( u1_FP_15 ) , .B( u1_L14_15 ) , .A( u1_out15_15 ) );
  XOR2_X1 u1_U51 (.B( u1_L0_24 ) , .Z( u1_N55 ) , .A( u1_out1_24 ) );
  XOR2_X1 u1_U510 (.Z( u1_FP_14 ) , .B( u1_L14_14 ) , .A( u1_out15_14 ) );
  XOR2_X1 u1_U511 (.Z( u1_FP_13 ) , .B( u1_L14_13 ) , .A( u1_out15_13 ) );
  XOR2_X1 u1_U512 (.Z( u1_FP_12 ) , .B( u1_L14_12 ) , .A( u1_out15_12 ) );
  XOR2_X1 u1_U513 (.Z( u1_FP_11 ) , .B( u1_L14_11 ) , .A( u1_out15_11 ) );
  XOR2_X1 u1_U514 (.Z( u1_FP_10 ) , .B( u1_L14_10 ) , .A( u1_out15_10 ) );
  XOR2_X1 u1_U52 (.B( u1_L0_23 ) , .Z( u1_N54 ) , .A( u1_out1_23 ) );
  XOR2_X1 u1_U53 (.B( u1_L0_22 ) , .Z( u1_N53 ) , .A( u1_out1_22 ) );
  XOR2_X1 u1_U54 (.B( u1_L0_21 ) , .Z( u1_N52 ) , .A( u1_out1_21 ) );
  XOR2_X1 u1_U55 (.B( u1_L0_20 ) , .Z( u1_N51 ) , .A( u1_out1_20 ) );
  XOR2_X1 u1_U56 (.B( u1_L0_19 ) , .Z( u1_N50 ) , .A( u1_out1_19 ) );
  XOR2_X1 u1_U57 (.Z( u1_N5 ) , .B( u1_desIn_r_46 ) , .A( u1_out0_6 ) );
  XOR2_X1 u1_U58 (.B( u1_L0_18 ) , .Z( u1_N49 ) , .A( u1_out1_18 ) );
  XOR2_X1 u1_U59 (.B( u1_L0_17 ) , .Z( u1_N48 ) , .A( u1_out1_17 ) );
  XOR2_X1 u1_U6 (.B( u1_L2_1 ) , .Z( u1_N96 ) , .A( u1_out3_1 ) );
  XOR2_X1 u1_U60 (.B( u1_L13_32 ) , .Z( u1_N479 ) , .A( u1_out14_32 ) );
  XOR2_X1 u1_U61 (.B( u1_L13_31 ) , .Z( u1_N478 ) , .A( u1_out14_31 ) );
  XOR2_X1 u1_U62 (.B( u1_L13_30 ) , .Z( u1_N477 ) , .A( u1_out14_30 ) );
  XOR2_X1 u1_U63 (.B( u1_L13_29 ) , .Z( u1_N476 ) , .A( u1_out14_29 ) );
  XOR2_X1 u1_U64 (.B( u1_L13_28 ) , .Z( u1_N475 ) , .A( u1_out14_28 ) );
  XOR2_X1 u1_U65 (.B( u1_L13_27 ) , .Z( u1_N474 ) , .A( u1_out14_27 ) );
  XOR2_X1 u1_U66 (.B( u1_L13_26 ) , .Z( u1_N473 ) , .A( u1_out14_26 ) );
  XOR2_X1 u1_U67 (.B( u1_L13_25 ) , .Z( u1_N472 ) , .A( u1_out14_25 ) );
  XOR2_X1 u1_U68 (.B( u1_L13_24 ) , .Z( u1_N471 ) , .A( u1_out14_24 ) );
  XOR2_X1 u1_U69 (.B( u1_L13_23 ) , .Z( u1_N470 ) , .A( u1_out14_23 ) );
  XOR2_X1 u1_U7 (.B( u1_L1_32 ) , .Z( u1_N95 ) , .A( u1_out2_32 ) );
  XOR2_X1 u1_U70 (.B( u1_L0_16 ) , .Z( u1_N47 ) , .A( u1_out1_16 ) );
  XOR2_X1 u1_U71 (.B( u1_L13_22 ) , .Z( u1_N469 ) , .A( u1_out14_22 ) );
  XOR2_X1 u1_U72 (.B( u1_L13_21 ) , .Z( u1_N468 ) , .A( u1_out14_21 ) );
  XOR2_X1 u1_U73 (.B( u1_L13_20 ) , .Z( u1_N467 ) , .A( u1_out14_20 ) );
  XOR2_X1 u1_U74 (.B( u1_L13_19 ) , .Z( u1_N466 ) , .A( u1_out14_19 ) );
  XOR2_X1 u1_U75 (.B( u1_L13_18 ) , .Z( u1_N465 ) , .A( u1_out14_18 ) );
  XOR2_X1 u1_U76 (.B( u1_L13_17 ) , .Z( u1_N464 ) , .A( u1_out14_17 ) );
  XOR2_X1 u1_U77 (.B( u1_L13_16 ) , .Z( u1_N463 ) , .A( u1_out14_16 ) );
  XOR2_X1 u1_U78 (.B( u1_L13_15 ) , .Z( u1_N462 ) , .A( u1_out14_15 ) );
  XOR2_X1 u1_U79 (.B( u1_L13_14 ) , .Z( u1_N461 ) , .A( u1_out14_14 ) );
  XOR2_X1 u1_U8 (.B( u1_L1_31 ) , .Z( u1_N94 ) , .A( u1_out2_31 ) );
  XOR2_X1 u1_U80 (.B( u1_L13_13 ) , .Z( u1_N460 ) , .A( u1_out14_13 ) );
  XOR2_X1 u1_U81 (.B( u1_L0_15 ) , .Z( u1_N46 ) , .A( u1_out1_15 ) );
  XOR2_X1 u1_U82 (.B( u1_L13_12 ) , .Z( u1_N459 ) , .A( u1_out14_12 ) );
  XOR2_X1 u1_U83 (.B( u1_L13_11 ) , .Z( u1_N458 ) , .A( u1_out14_11 ) );
  XOR2_X1 u1_U84 (.B( u1_L13_10 ) , .Z( u1_N457 ) , .A( u1_out14_10 ) );
  XOR2_X1 u1_U85 (.B( u1_L13_9 ) , .Z( u1_N456 ) , .A( u1_out14_9 ) );
  XOR2_X1 u1_U86 (.B( u1_L13_8 ) , .Z( u1_N455 ) , .A( u1_out14_8 ) );
  XOR2_X1 u1_U87 (.B( u1_L13_7 ) , .Z( u1_N454 ) , .A( u1_out14_7 ) );
  XOR2_X1 u1_U88 (.B( u1_L13_6 ) , .Z( u1_N453 ) , .A( u1_out14_6 ) );
  XOR2_X1 u1_U89 (.B( u1_L13_5 ) , .Z( u1_N452 ) , .A( u1_out14_5 ) );
  XOR2_X1 u1_U9 (.B( u1_L1_30 ) , .Z( u1_N93 ) , .A( u1_out2_30 ) );
  XOR2_X1 u1_U90 (.B( u1_L13_4 ) , .Z( u1_N451 ) , .A( u1_out14_4 ) );
  XOR2_X1 u1_U91 (.B( u1_L13_3 ) , .Z( u1_N450 ) , .A( u1_out14_3 ) );
  XOR2_X1 u1_U92 (.B( u1_L0_14 ) , .Z( u1_N45 ) , .A( u1_out1_14 ) );
  XOR2_X1 u1_U93 (.B( u1_L13_2 ) , .Z( u1_N449 ) , .A( u1_out14_2 ) );
  XOR2_X1 u1_U94 (.B( u1_L13_1 ) , .Z( u1_N448 ) , .A( u1_out14_1 ) );
  XOR2_X1 u1_U95 (.B( u1_L12_32 ) , .Z( u1_N447 ) , .A( u1_out13_32 ) );
  XOR2_X1 u1_U96 (.B( u1_L12_31 ) , .Z( u1_N446 ) , .A( u1_out13_31 ) );
  XOR2_X1 u1_U97 (.B( u1_L12_30 ) , .Z( u1_N445 ) , .A( u1_out13_30 ) );
  XOR2_X1 u1_U98 (.B( u1_L12_29 ) , .Z( u1_N444 ) , .A( u1_out13_29 ) );
  XOR2_X1 u1_U99 (.B( u1_L12_28 ) , .Z( u1_N443 ) , .A( u1_out13_28 ) );
  DFF_X1 u1_desIn_r_reg_0 (.CK( clk ) , .D( stage1_out_0 ) , .Q( u1_desIn_r_0 ) );
  DFF_X1 u1_desIn_r_reg_1 (.CK( clk ) , .D( stage1_out_1 ) , .Q( u1_desIn_r_1 ) );
  DFF_X1 u1_desIn_r_reg_10 (.CK( clk ) , .D( stage1_out_10 ) , .Q( u1_desIn_r_10 ) );
  DFF_X1 u1_desIn_r_reg_11 (.CK( clk ) , .D( stage1_out_11 ) , .Q( u1_desIn_r_11 ) );
  DFF_X1 u1_desIn_r_reg_12 (.CK( clk ) , .D( stage1_out_12 ) , .Q( u1_desIn_r_12 ) );
  DFF_X1 u1_desIn_r_reg_13 (.CK( clk ) , .D( stage1_out_13 ) , .Q( u1_desIn_r_13 ) );
  DFF_X1 u1_desIn_r_reg_14 (.CK( clk ) , .D( stage1_out_14 ) , .Q( u1_desIn_r_14 ) );
  DFF_X1 u1_desIn_r_reg_15 (.CK( clk ) , .D( stage1_out_15 ) , .Q( u1_desIn_r_15 ) );
  DFF_X1 u1_desIn_r_reg_16 (.CK( clk ) , .D( stage1_out_16 ) , .Q( u1_desIn_r_16 ) );
  DFF_X1 u1_desIn_r_reg_17 (.CK( clk ) , .D( stage1_out_17 ) , .Q( u1_desIn_r_17 ) );
  DFF_X1 u1_desIn_r_reg_18 (.CK( clk ) , .D( stage1_out_18 ) , .Q( u1_desIn_r_18 ) );
  DFF_X1 u1_desIn_r_reg_19 (.CK( clk ) , .D( stage1_out_19 ) , .Q( u1_desIn_r_19 ) );
  DFF_X1 u1_desIn_r_reg_2 (.CK( clk ) , .D( stage1_out_2 ) , .Q( u1_desIn_r_2 ) );
  DFF_X1 u1_desIn_r_reg_20 (.CK( clk ) , .D( stage1_out_20 ) , .Q( u1_desIn_r_20 ) );
  DFF_X1 u1_desIn_r_reg_21 (.CK( clk ) , .D( stage1_out_21 ) , .Q( u1_desIn_r_21 ) );
  DFF_X1 u1_desIn_r_reg_22 (.CK( clk ) , .D( stage1_out_22 ) , .Q( u1_desIn_r_22 ) );
  DFF_X1 u1_desIn_r_reg_23 (.CK( clk ) , .D( stage1_out_23 ) , .Q( u1_desIn_r_23 ) );
  DFF_X1 u1_desIn_r_reg_24 (.CK( clk ) , .D( stage1_out_24 ) , .Q( u1_desIn_r_24 ) );
  DFF_X1 u1_desIn_r_reg_25 (.CK( clk ) , .D( stage1_out_25 ) , .Q( u1_desIn_r_25 ) );
  DFF_X1 u1_desIn_r_reg_26 (.CK( clk ) , .D( stage1_out_26 ) , .Q( u1_desIn_r_26 ) );
  DFF_X1 u1_desIn_r_reg_27 (.CK( clk ) , .D( stage1_out_27 ) , .Q( u1_desIn_r_27 ) );
  DFF_X1 u1_desIn_r_reg_28 (.CK( clk ) , .D( stage1_out_28 ) , .Q( u1_desIn_r_28 ) );
  DFF_X1 u1_desIn_r_reg_29 (.CK( clk ) , .D( stage1_out_29 ) , .Q( u1_desIn_r_29 ) );
  DFF_X1 u1_desIn_r_reg_3 (.CK( clk ) , .D( stage1_out_3 ) , .Q( u1_desIn_r_3 ) );
  DFF_X1 u1_desIn_r_reg_30 (.CK( clk ) , .D( stage1_out_30 ) , .Q( u1_desIn_r_30 ) );
  DFF_X1 u1_desIn_r_reg_31 (.CK( clk ) , .D( stage1_out_31 ) , .Q( u1_desIn_r_31 ) );
  DFF_X1 u1_desIn_r_reg_32 (.CK( clk ) , .D( stage1_out_32 ) , .Q( u1_desIn_r_32 ) );
  DFF_X1 u1_desIn_r_reg_33 (.CK( clk ) , .D( stage1_out_33 ) , .Q( u1_desIn_r_33 ) );
  DFF_X1 u1_desIn_r_reg_34 (.CK( clk ) , .D( stage1_out_34 ) , .Q( u1_desIn_r_34 ) );
  DFF_X1 u1_desIn_r_reg_35 (.CK( clk ) , .D( stage1_out_35 ) , .Q( u1_desIn_r_35 ) );
  DFF_X1 u1_desIn_r_reg_36 (.CK( clk ) , .D( stage1_out_36 ) , .Q( u1_desIn_r_36 ) );
  DFF_X1 u1_desIn_r_reg_37 (.CK( clk ) , .D( stage1_out_37 ) , .Q( u1_desIn_r_37 ) );
  DFF_X1 u1_desIn_r_reg_38 (.CK( clk ) , .D( stage1_out_38 ) , .Q( u1_desIn_r_38 ) );
  DFF_X1 u1_desIn_r_reg_39 (.CK( clk ) , .D( stage1_out_39 ) , .Q( u1_desIn_r_39 ) );
  DFF_X1 u1_desIn_r_reg_4 (.CK( clk ) , .D( stage1_out_4 ) , .Q( u1_desIn_r_4 ) );
  DFF_X1 u1_desIn_r_reg_40 (.CK( clk ) , .D( stage1_out_40 ) , .Q( u1_desIn_r_40 ) );
  DFF_X1 u1_desIn_r_reg_41 (.CK( clk ) , .D( stage1_out_41 ) , .Q( u1_desIn_r_41 ) );
  DFF_X1 u1_desIn_r_reg_42 (.CK( clk ) , .D( stage1_out_42 ) , .Q( u1_desIn_r_42 ) );
  DFF_X1 u1_desIn_r_reg_43 (.CK( clk ) , .D( stage1_out_43 ) , .Q( u1_desIn_r_43 ) );
  DFF_X1 u1_desIn_r_reg_44 (.CK( clk ) , .D( stage1_out_44 ) , .Q( u1_desIn_r_44 ) );
  DFF_X1 u1_desIn_r_reg_45 (.CK( clk ) , .D( stage1_out_45 ) , .Q( u1_desIn_r_45 ) );
  DFF_X1 u1_desIn_r_reg_46 (.CK( clk ) , .D( stage1_out_46 ) , .Q( u1_desIn_r_46 ) );
  DFF_X1 u1_desIn_r_reg_47 (.CK( clk ) , .D( stage1_out_47 ) , .Q( u1_desIn_r_47 ) );
  DFF_X1 u1_desIn_r_reg_48 (.CK( clk ) , .D( stage1_out_48 ) , .Q( u1_desIn_r_48 ) );
  DFF_X1 u1_desIn_r_reg_49 (.CK( clk ) , .D( stage1_out_49 ) , .Q( u1_desIn_r_49 ) );
  DFF_X1 u1_desIn_r_reg_5 (.CK( clk ) , .D( stage1_out_5 ) , .Q( u1_desIn_r_5 ) );
  DFF_X1 u1_desIn_r_reg_50 (.CK( clk ) , .D( stage1_out_50 ) , .Q( u1_desIn_r_50 ) );
  DFF_X1 u1_desIn_r_reg_51 (.CK( clk ) , .D( stage1_out_51 ) , .Q( u1_desIn_r_51 ) );
  DFF_X1 u1_desIn_r_reg_52 (.CK( clk ) , .D( stage1_out_52 ) , .Q( u1_desIn_r_52 ) );
  DFF_X1 u1_desIn_r_reg_53 (.CK( clk ) , .D( stage1_out_53 ) , .Q( u1_desIn_r_53 ) );
  DFF_X1 u1_desIn_r_reg_54 (.CK( clk ) , .D( stage1_out_54 ) , .Q( u1_desIn_r_54 ) );
  DFF_X1 u1_desIn_r_reg_55 (.CK( clk ) , .D( stage1_out_55 ) , .Q( u1_desIn_r_55 ) );
  DFF_X1 u1_desIn_r_reg_56 (.CK( clk ) , .D( stage1_out_56 ) , .Q( u1_desIn_r_56 ) );
  DFF_X1 u1_desIn_r_reg_57 (.CK( clk ) , .D( stage1_out_57 ) , .Q( u1_desIn_r_57 ) );
  DFF_X1 u1_desIn_r_reg_58 (.CK( clk ) , .D( stage1_out_58 ) , .Q( u1_desIn_r_58 ) );
  DFF_X1 u1_desIn_r_reg_59 (.CK( clk ) , .D( stage1_out_59 ) , .Q( u1_desIn_r_59 ) );
  DFF_X1 u1_desIn_r_reg_6 (.CK( clk ) , .D( stage1_out_6 ) , .Q( u1_desIn_r_6 ) );
  DFF_X1 u1_desIn_r_reg_60 (.CK( clk ) , .D( stage1_out_60 ) , .Q( u1_desIn_r_60 ) );
  DFF_X1 u1_desIn_r_reg_61 (.CK( clk ) , .D( stage1_out_61 ) , .Q( u1_desIn_r_61 ) );
  DFF_X1 u1_desIn_r_reg_62 (.CK( clk ) , .D( stage1_out_62 ) , .Q( u1_desIn_r_62 ) );
  DFF_X1 u1_desIn_r_reg_63 (.CK( clk ) , .D( stage1_out_63 ) , .Q( u1_desIn_r_63 ) );
  DFF_X1 u1_desIn_r_reg_7 (.CK( clk ) , .D( stage1_out_7 ) , .Q( u1_desIn_r_7 ) );
  DFF_X1 u1_desIn_r_reg_8 (.CK( clk ) , .D( stage1_out_8 ) , .Q( u1_desIn_r_8 ) );
  DFF_X1 u1_desIn_r_reg_9 (.CK( clk ) , .D( stage1_out_9 ) , .Q( u1_desIn_r_9 ) );
  DFF_X1 u1_desOut_reg_0 (.CK( clk ) , .Q( stage2_out_0 ) , .D( u1_FP_25 ) );
  DFF_X1 u1_desOut_reg_1 (.CK( clk ) , .Q( stage2_out_1 ) , .D( u1_FP_57 ) );
  DFF_X1 u1_desOut_reg_10 (.CK( clk ) , .Q( stage2_out_10 ) , .D( u1_FP_18 ) );
  DFF_X1 u1_desOut_reg_11 (.CK( clk ) , .Q( stage2_out_11 ) , .D( u1_FP_50 ) );
  DFF_X1 u1_desOut_reg_12 (.CK( clk ) , .Q( stage2_out_12 ) , .D( u1_FP_10 ) );
  DFF_X1 u1_desOut_reg_13 (.CK( clk ) , .Q( stage2_out_13 ) , .D( u1_FP_42 ) );
  DFF_X1 u1_desOut_reg_14 (.CK( clk ) , .Q( stage2_out_14 ) , .D( u1_FP_2 ) );
  DFF_X1 u1_desOut_reg_15 (.CK( clk ) , .Q( stage2_out_15 ) , .D( u1_FP_34 ) );
  DFF_X1 u1_desOut_reg_16 (.CK( clk ) , .Q( stage2_out_16 ) , .D( u1_FP_27 ) );
  DFF_X1 u1_desOut_reg_17 (.CK( clk ) , .Q( stage2_out_17 ) , .D( u1_FP_59 ) );
  DFF_X1 u1_desOut_reg_18 (.CK( clk ) , .Q( stage2_out_18 ) , .D( u1_FP_19 ) );
  DFF_X1 u1_desOut_reg_19 (.CK( clk ) , .Q( stage2_out_19 ) , .D( u1_FP_51 ) );
  DFF_X1 u1_desOut_reg_2 (.CK( clk ) , .Q( stage2_out_2 ) , .D( u1_FP_17 ) );
  DFF_X1 u1_desOut_reg_20 (.CK( clk ) , .Q( stage2_out_20 ) , .D( u1_FP_11 ) );
  DFF_X1 u1_desOut_reg_21 (.CK( clk ) , .Q( stage2_out_21 ) , .D( u1_FP_43 ) );
  DFF_X1 u1_desOut_reg_22 (.CK( clk ) , .Q( stage2_out_22 ) , .D( u1_FP_3 ) );
  DFF_X1 u1_desOut_reg_23 (.CK( clk ) , .Q( stage2_out_23 ) , .D( u1_FP_35 ) );
  DFF_X1 u1_desOut_reg_24 (.CK( clk ) , .Q( stage2_out_24 ) , .D( u1_FP_28 ) );
  DFF_X1 u1_desOut_reg_25 (.CK( clk ) , .Q( stage2_out_25 ) , .D( u1_FP_60 ) );
  DFF_X1 u1_desOut_reg_26 (.CK( clk ) , .Q( stage2_out_26 ) , .D( u1_FP_20 ) );
  DFF_X1 u1_desOut_reg_27 (.CK( clk ) , .Q( stage2_out_27 ) , .D( u1_FP_52 ) );
  DFF_X1 u1_desOut_reg_28 (.CK( clk ) , .Q( stage2_out_28 ) , .D( u1_FP_12 ) );
  DFF_X1 u1_desOut_reg_29 (.CK( clk ) , .Q( stage2_out_29 ) , .D( u1_FP_44 ) );
  DFF_X1 u1_desOut_reg_3 (.CK( clk ) , .Q( stage2_out_3 ) , .D( u1_FP_49 ) );
  DFF_X1 u1_desOut_reg_30 (.CK( clk ) , .Q( stage2_out_30 ) , .D( u1_FP_4 ) );
  DFF_X1 u1_desOut_reg_31 (.CK( clk ) , .Q( stage2_out_31 ) , .D( u1_FP_36 ) );
  DFF_X1 u1_desOut_reg_32 (.CK( clk ) , .Q( stage2_out_32 ) , .D( u1_FP_29 ) );
  DFF_X1 u1_desOut_reg_33 (.CK( clk ) , .Q( stage2_out_33 ) , .D( u1_FP_61 ) );
  DFF_X1 u1_desOut_reg_34 (.CK( clk ) , .Q( stage2_out_34 ) , .D( u1_FP_21 ) );
  DFF_X1 u1_desOut_reg_35 (.CK( clk ) , .Q( stage2_out_35 ) , .D( u1_FP_53 ) );
  DFF_X1 u1_desOut_reg_36 (.CK( clk ) , .Q( stage2_out_36 ) , .D( u1_FP_13 ) );
  DFF_X1 u1_desOut_reg_37 (.CK( clk ) , .Q( stage2_out_37 ) , .D( u1_FP_45 ) );
  DFF_X1 u1_desOut_reg_38 (.CK( clk ) , .Q( stage2_out_38 ) , .D( u1_FP_5 ) );
  DFF_X1 u1_desOut_reg_39 (.CK( clk ) , .Q( stage2_out_39 ) , .D( u1_FP_37 ) );
  DFF_X1 u1_desOut_reg_4 (.CK( clk ) , .Q( stage2_out_4 ) , .D( u1_FP_9 ) );
  DFF_X1 u1_desOut_reg_40 (.CK( clk ) , .Q( stage2_out_40 ) , .D( u1_FP_30 ) );
  DFF_X1 u1_desOut_reg_41 (.CK( clk ) , .Q( stage2_out_41 ) , .D( u1_FP_62 ) );
  DFF_X1 u1_desOut_reg_42 (.CK( clk ) , .Q( stage2_out_42 ) , .D( u1_FP_22 ) );
  DFF_X1 u1_desOut_reg_43 (.CK( clk ) , .Q( stage2_out_43 ) , .D( u1_FP_54 ) );
  DFF_X1 u1_desOut_reg_44 (.CK( clk ) , .Q( stage2_out_44 ) , .D( u1_FP_14 ) );
  DFF_X1 u1_desOut_reg_45 (.CK( clk ) , .Q( stage2_out_45 ) , .D( u1_FP_46 ) );
  DFF_X1 u1_desOut_reg_46 (.CK( clk ) , .Q( stage2_out_46 ) , .D( u1_FP_6 ) );
  DFF_X1 u1_desOut_reg_47 (.CK( clk ) , .Q( stage2_out_47 ) , .D( u1_FP_38 ) );
  DFF_X1 u1_desOut_reg_48 (.CK( clk ) , .Q( stage2_out_48 ) , .D( u1_FP_31 ) );
  DFF_X1 u1_desOut_reg_49 (.CK( clk ) , .Q( stage2_out_49 ) , .D( u1_FP_63 ) );
  DFF_X1 u1_desOut_reg_5 (.CK( clk ) , .Q( stage2_out_5 ) , .D( u1_FP_41 ) );
  DFF_X1 u1_desOut_reg_50 (.CK( clk ) , .Q( stage2_out_50 ) , .D( u1_FP_23 ) );
  DFF_X1 u1_desOut_reg_51 (.CK( clk ) , .Q( stage2_out_51 ) , .D( u1_FP_55 ) );
  DFF_X1 u1_desOut_reg_52 (.CK( clk ) , .Q( stage2_out_52 ) , .D( u1_FP_15 ) );
  DFF_X1 u1_desOut_reg_53 (.CK( clk ) , .Q( stage2_out_53 ) , .D( u1_FP_47 ) );
  DFF_X1 u1_desOut_reg_54 (.CK( clk ) , .Q( stage2_out_54 ) , .D( u1_FP_7 ) );
  DFF_X1 u1_desOut_reg_55 (.CK( clk ) , .Q( stage2_out_55 ) , .D( u1_FP_39 ) );
  DFF_X1 u1_desOut_reg_56 (.CK( clk ) , .Q( stage2_out_56 ) , .D( u1_FP_32 ) );
  DFF_X1 u1_desOut_reg_57 (.CK( clk ) , .Q( stage2_out_57 ) , .D( u1_FP_64 ) );
  DFF_X1 u1_desOut_reg_58 (.CK( clk ) , .Q( stage2_out_58 ) , .D( u1_FP_24 ) );
  DFF_X1 u1_desOut_reg_59 (.CK( clk ) , .Q( stage2_out_59 ) , .D( u1_FP_56 ) );
  DFF_X1 u1_desOut_reg_6 (.CK( clk ) , .Q( stage2_out_6 ) , .D( u1_FP_1 ) );
  DFF_X1 u1_desOut_reg_60 (.CK( clk ) , .Q( stage2_out_60 ) , .D( u1_FP_16 ) );
  DFF_X1 u1_desOut_reg_61 (.CK( clk ) , .Q( stage2_out_61 ) , .D( u1_FP_48 ) );
  DFF_X1 u1_desOut_reg_62 (.CK( clk ) , .Q( stage2_out_62 ) , .D( u1_FP_8 ) );
  DFF_X1 u1_desOut_reg_63 (.CK( clk ) , .Q( stage2_out_63 ) , .D( u1_FP_40 ) );
  DFF_X1 u1_desOut_reg_7 (.CK( clk ) , .Q( stage2_out_7 ) , .D( u1_FP_33 ) );
  DFF_X1 u1_desOut_reg_8 (.CK( clk ) , .Q( stage2_out_8 ) , .D( u1_FP_26 ) );
  DFF_X1 u1_desOut_reg_9 (.CK( clk ) , .Q( stage2_out_9 ) , .D( u1_FP_58 ) );
  DFF_X1 u1_key_r_reg_0 (.CK( clk ) , .D( key_b_r_16_0 ) , .Q( u1_key_r_0 ) );
  DFF_X1 u1_key_r_reg_1 (.CK( clk ) , .D( key_b_r_16_1 ) , .Q( u1_key_r_1 ) );
  DFF_X1 u1_key_r_reg_10 (.CK( clk ) , .D( key_b_r_16_10 ) , .Q( u1_key_r_10 ) );
  DFF_X1 u1_key_r_reg_11 (.CK( clk ) , .D( key_b_r_16_11 ) , .Q( u1_key_r_11 ) );
  DFF_X1 u1_key_r_reg_12 (.CK( clk ) , .D( key_b_r_16_12 ) , .Q( u1_key_r_12 ) );
  DFF_X1 u1_key_r_reg_13 (.CK( clk ) , .D( key_b_r_16_13 ) , .Q( u1_key_r_13 ) );
  DFF_X1 u1_key_r_reg_14 (.CK( clk ) , .D( key_b_r_16_14 ) , .Q( u1_key_r_14 ) );
  DFF_X1 u1_key_r_reg_15 (.CK( clk ) , .D( key_b_r_16_15 ) , .Q( u1_key_r_15 ) );
  DFF_X1 u1_key_r_reg_16 (.CK( clk ) , .D( key_b_r_16_16 ) , .Q( u1_key_r_16 ) );
  DFF_X1 u1_key_r_reg_17 (.CK( clk ) , .D( key_b_r_16_17 ) , .Q( u1_key_r_17 ) );
  DFF_X1 u1_key_r_reg_18 (.CK( clk ) , .D( key_b_r_16_18 ) , .Q( u1_key_r_18 ) );
  DFF_X1 u1_key_r_reg_19 (.CK( clk ) , .D( key_b_r_16_19 ) , .Q( u1_key_r_19 ) );
  DFF_X1 u1_key_r_reg_2 (.CK( clk ) , .D( key_b_r_16_2 ) , .Q( u1_key_r_2 ) );
  DFF_X1 u1_key_r_reg_20 (.CK( clk ) , .D( key_b_r_16_20 ) , .Q( u1_key_r_20 ) );
  DFF_X1 u1_key_r_reg_21 (.CK( clk ) , .D( key_b_r_16_21 ) , .Q( u1_key_r_21 ) );
  DFF_X1 u1_key_r_reg_22 (.CK( clk ) , .D( key_b_r_16_22 ) , .Q( u1_key_r_22 ) );
  DFF_X1 u1_key_r_reg_23 (.CK( clk ) , .D( key_b_r_16_23 ) , .Q( u1_key_r_23 ) );
  DFF_X1 u1_key_r_reg_24 (.CK( clk ) , .D( key_b_r_16_24 ) , .Q( u1_key_r_24 ) );
  DFF_X1 u1_key_r_reg_25 (.CK( clk ) , .D( key_b_r_16_25 ) , .Q( u1_key_r_25 ) );
  DFF_X1 u1_key_r_reg_26 (.CK( clk ) , .D( key_b_r_16_26 ) , .Q( u1_key_r_26 ) );
  DFF_X1 u1_key_r_reg_27 (.CK( clk ) , .D( key_b_r_16_27 ) , .Q( u1_key_r_27 ) );
  DFF_X1 u1_key_r_reg_28 (.CK( clk ) , .D( key_b_r_16_28 ) , .Q( u1_key_r_28 ) );
  DFF_X1 u1_key_r_reg_29 (.CK( clk ) , .D( key_b_r_16_29 ) , .Q( u1_key_r_29 ) );
  DFF_X1 u1_key_r_reg_3 (.CK( clk ) , .D( key_b_r_16_3 ) , .Q( u1_key_r_3 ) );
  DFF_X1 u1_key_r_reg_30 (.CK( clk ) , .D( key_b_r_16_30 ) , .Q( u1_key_r_30 ) );
  DFF_X1 u1_key_r_reg_31 (.CK( clk ) , .D( key_b_r_16_31 ) , .Q( u1_key_r_31 ) );
  DFF_X1 u1_key_r_reg_32 (.CK( clk ) , .D( key_b_r_16_32 ) , .Q( u1_key_r_32 ) );
  DFF_X1 u1_key_r_reg_33 (.CK( clk ) , .D( key_b_r_16_33 ) , .Q( u1_key_r_33 ) );
  DFF_X1 u1_key_r_reg_34 (.CK( clk ) , .D( key_b_r_16_34 ) , .Q( u1_key_r_34 ) );
  DFF_X1 u1_key_r_reg_35 (.CK( clk ) , .D( key_b_r_16_35 ) , .Q( u1_key_r_35 ) );
  DFF_X1 u1_key_r_reg_36 (.CK( clk ) , .D( key_b_r_16_36 ) , .Q( u1_key_r_36 ) );
  DFF_X1 u1_key_r_reg_37 (.CK( clk ) , .D( key_b_r_16_37 ) , .Q( u1_key_r_37 ) );
  DFF_X1 u1_key_r_reg_38 (.CK( clk ) , .D( key_b_r_16_38 ) , .Q( u1_key_r_38 ) );
  DFF_X1 u1_key_r_reg_39 (.CK( clk ) , .D( key_b_r_16_39 ) , .Q( u1_key_r_39 ) );
  DFF_X1 u1_key_r_reg_4 (.CK( clk ) , .D( key_b_r_16_4 ) , .Q( u1_key_r_4 ) );
  DFF_X1 u1_key_r_reg_40 (.CK( clk ) , .D( key_b_r_16_40 ) , .Q( u1_key_r_40 ) );
  DFF_X1 u1_key_r_reg_41 (.CK( clk ) , .D( key_b_r_16_41 ) , .Q( u1_key_r_41 ) );
  DFF_X1 u1_key_r_reg_42 (.CK( clk ) , .D( key_b_r_16_42 ) , .Q( u1_key_r_42 ) );
  DFF_X1 u1_key_r_reg_43 (.CK( clk ) , .D( key_b_r_16_43 ) , .Q( u1_key_r_43 ) );
  DFF_X1 u1_key_r_reg_44 (.CK( clk ) , .D( key_b_r_16_44 ) , .Q( u1_key_r_44 ) );
  DFF_X1 u1_key_r_reg_45 (.CK( clk ) , .D( key_b_r_16_45 ) , .Q( u1_key_r_45 ) );
  DFF_X1 u1_key_r_reg_46 (.CK( clk ) , .D( key_b_r_16_46 ) , .Q( u1_key_r_46 ) );
  DFF_X1 u1_key_r_reg_47 (.CK( clk ) , .D( key_b_r_16_47 ) , .Q( u1_key_r_47 ) );
  DFF_X1 u1_key_r_reg_48 (.CK( clk ) , .D( key_b_r_16_48 ) , .Q( u1_key_r_48 ) );
  DFF_X1 u1_key_r_reg_49 (.CK( clk ) , .D( key_b_r_16_49 ) , .Q( u1_key_r_49 ) );
  DFF_X1 u1_key_r_reg_5 (.CK( clk ) , .D( key_b_r_16_5 ) , .Q( u1_key_r_5 ) );
  DFF_X1 u1_key_r_reg_50 (.CK( clk ) , .D( key_b_r_16_50 ) , .Q( u1_key_r_50 ) );
  DFF_X1 u1_key_r_reg_51 (.CK( clk ) , .D( key_b_r_16_51 ) , .Q( u1_key_r_51 ) );
  DFF_X1 u1_key_r_reg_52 (.CK( clk ) , .D( key_b_r_16_52 ) , .Q( u1_key_r_52 ) );
  DFF_X1 u1_key_r_reg_53 (.CK( clk ) , .D( key_b_r_16_53 ) , .Q( u1_key_r_53 ) );
  DFF_X1 u1_key_r_reg_54 (.CK( clk ) , .D( key_b_r_16_54 ) , .Q( u1_key_r_54 ) );
  DFF_X1 u1_key_r_reg_55 (.CK( clk ) , .D( key_b_r_16_55 ) , .Q( u1_key_r_55 ) );
  DFF_X1 u1_key_r_reg_6 (.CK( clk ) , .D( key_b_r_16_6 ) , .Q( u1_key_r_6 ) );
  DFF_X1 u1_key_r_reg_7 (.CK( clk ) , .D( key_b_r_16_7 ) , .Q( u1_key_r_7 ) );
  DFF_X1 u1_key_r_reg_8 (.CK( clk ) , .D( key_b_r_16_8 ) , .Q( u1_key_r_8 ) );
  DFF_X1 u1_key_r_reg_9 (.CK( clk ) , .D( key_b_r_16_9 ) , .Q( u1_key_r_9 ) );
  XOR2_X1 u1_u0_U1 (.B( u1_K1_9 ) , .A( u1_desIn_r_47 ) , .Z( u1_u0_X_9 ) );
  XOR2_X1 u1_u0_U10 (.B( u1_K1_45 ) , .A( u1_desIn_r_41 ) , .Z( u1_u0_X_45 ) );
  XOR2_X1 u1_u0_U11 (.B( u1_K1_44 ) , .A( u1_desIn_r_33 ) , .Z( u1_u0_X_44 ) );
  XOR2_X1 u1_u0_U13 (.B( u1_K1_42 ) , .A( u1_desIn_r_33 ) , .Z( u1_u0_X_42 ) );
  XOR2_X1 u1_u0_U15 (.B( u1_K1_40 ) , .A( u1_desIn_r_17 ) , .Z( u1_u0_X_40 ) );
  XOR2_X1 u1_u0_U16 (.B( u1_K1_3 ) , .A( u1_desIn_r_15 ) , .Z( u1_u0_X_3 ) );
  XOR2_X1 u1_u0_U17 (.B( u1_K1_39 ) , .A( u1_desIn_r_9 ) , .Z( u1_u0_X_39 ) );
  XOR2_X1 u1_u0_U18 (.B( u1_K1_38 ) , .A( u1_desIn_r_1 ) , .Z( u1_u0_X_38 ) );
  XOR2_X1 u1_u0_U19 (.B( u1_K1_37 ) , .A( u1_desIn_r_59 ) , .Z( u1_u0_X_37 ) );
  XOR2_X1 u1_u0_U20 (.B( u1_K1_36 ) , .A( u1_desIn_r_1 ) , .Z( u1_u0_X_36 ) );
  XOR2_X1 u1_u0_U21 (.B( u1_K1_35 ) , .A( u1_desIn_r_59 ) , .Z( u1_u0_X_35 ) );
  XOR2_X1 u1_u0_U22 (.B( u1_K1_34 ) , .A( u1_desIn_r_51 ) , .Z( u1_u0_X_34 ) );
  XOR2_X1 u1_u0_U23 (.B( u1_K1_33 ) , .A( u1_desIn_r_43 ) , .Z( u1_u0_X_33 ) );
  XOR2_X1 u1_u0_U24 (.B( u1_K1_32 ) , .A( u1_desIn_r_35 ) , .Z( u1_u0_X_32 ) );
  XOR2_X1 u1_u0_U25 (.B( u1_K1_31 ) , .A( u1_desIn_r_27 ) , .Z( u1_u0_X_31 ) );
  XOR2_X1 u1_u0_U26 (.B( u1_K1_30 ) , .A( u1_desIn_r_35 ) , .Z( u1_u0_X_30 ) );
  XOR2_X1 u1_u0_U27 (.B( u1_K1_2 ) , .A( u1_desIn_r_7 ) , .Z( u1_u0_X_2 ) );
  XOR2_X1 u1_u0_U28 (.B( u1_K1_29 ) , .A( u1_desIn_r_27 ) , .Z( u1_u0_X_29 ) );
  XOR2_X1 u1_u0_U29 (.B( u1_K1_28 ) , .A( u1_desIn_r_19 ) , .Z( u1_u0_X_28 ) );
  XOR2_X1 u1_u0_U3 (.B( u1_K1_7 ) , .A( u1_desIn_r_31 ) , .Z( u1_u0_X_7 ) );
  XOR2_X1 u1_u0_U30 (.B( u1_K1_27 ) , .A( u1_desIn_r_11 ) , .Z( u1_u0_X_27 ) );
  XOR2_X1 u1_u0_U31 (.B( u1_K1_26 ) , .A( u1_desIn_r_3 ) , .Z( u1_u0_X_26 ) );
  XOR2_X1 u1_u0_U32 (.B( u1_K1_25 ) , .A( u1_desIn_r_61 ) , .Z( u1_u0_X_25 ) );
  XOR2_X1 u1_u0_U33 (.B( u1_K1_24 ) , .A( u1_desIn_r_3 ) , .Z( u1_u0_X_24 ) );
  XOR2_X1 u1_u0_U34 (.B( u1_K1_23 ) , .A( u1_desIn_r_61 ) , .Z( u1_u0_X_23 ) );
  XOR2_X1 u1_u0_U35 (.B( u1_K1_22 ) , .A( u1_desIn_r_53 ) , .Z( u1_u0_X_22 ) );
  XOR2_X1 u1_u0_U36 (.B( u1_K1_21 ) , .A( u1_desIn_r_45 ) , .Z( u1_u0_X_21 ) );
  XOR2_X1 u1_u0_U42 (.B( u1_K1_16 ) , .A( u1_desIn_r_21 ) , .Z( u1_u0_X_16 ) );
  XOR2_X1 u1_u0_U43 (.B( u1_K1_15 ) , .A( u1_desIn_r_13 ) , .Z( u1_u0_X_15 ) );
  XOR2_X1 u1_u0_U44 (.B( u1_K1_14 ) , .A( u1_desIn_r_5 ) , .Z( u1_u0_X_14 ) );
  XOR2_X1 u1_u0_U45 (.B( u1_K1_13 ) , .A( u1_desIn_r_63 ) , .Z( u1_u0_X_13 ) );
  XOR2_X1 u1_u0_U46 (.B( u1_K1_12 ) , .A( u1_desIn_r_5 ) , .Z( u1_u0_X_12 ) );
  XOR2_X1 u1_u0_U47 (.B( u1_K1_11 ) , .A( u1_desIn_r_63 ) , .Z( u1_u0_X_11 ) );
  XOR2_X1 u1_u0_U48 (.B( u1_K1_10 ) , .A( u1_desIn_r_55 ) , .Z( u1_u0_X_10 ) );
  XOR2_X1 u1_u0_U5 (.B( u1_K1_5 ) , .A( u1_desIn_r_31 ) , .Z( u1_u0_X_5 ) );
  XOR2_X1 u1_u0_U6 (.B( u1_K1_4 ) , .A( u1_desIn_r_23 ) , .Z( u1_u0_X_4 ) );
  XOR2_X1 u1_u0_U7 (.B( u1_K1_48 ) , .A( u1_desIn_r_7 ) , .Z( u1_u0_X_48 ) );
  XOR2_X1 u1_u0_U9 (.B( u1_K1_46 ) , .A( u1_desIn_r_49 ) , .Z( u1_u0_X_46 ) );
  XOR2_X1 u1_u10_U1 (.B( u1_K11_9 ) , .A( u1_R9_6 ) , .Z( u1_u10_X_9 ) );
  XOR2_X1 u1_u10_U10 (.B( u1_K11_45 ) , .A( u1_R9_30 ) , .Z( u1_u10_X_45 ) );
  XOR2_X1 u1_u10_U11 (.B( u1_K11_44 ) , .A( u1_R9_29 ) , .Z( u1_u10_X_44 ) );
  XOR2_X1 u1_u10_U12 (.B( u1_K11_43 ) , .A( u1_R9_28 ) , .Z( u1_u10_X_43 ) );
  XOR2_X1 u1_u10_U13 (.B( u1_K11_42 ) , .A( u1_R9_29 ) , .Z( u1_u10_X_42 ) );
  XOR2_X1 u1_u10_U14 (.B( u1_K11_41 ) , .A( u1_R9_28 ) , .Z( u1_u10_X_41 ) );
  XOR2_X1 u1_u10_U15 (.B( u1_K11_40 ) , .A( u1_R9_27 ) , .Z( u1_u10_X_40 ) );
  XOR2_X1 u1_u10_U16 (.B( u1_K11_3 ) , .A( u1_R9_2 ) , .Z( u1_u10_X_3 ) );
  XOR2_X1 u1_u10_U17 (.B( u1_K11_39 ) , .A( u1_R9_26 ) , .Z( u1_u10_X_39 ) );
  XOR2_X1 u1_u10_U2 (.B( u1_K11_8 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_8 ) );
  XOR2_X1 u1_u10_U23 (.B( u1_K11_33 ) , .A( u1_R9_22 ) , .Z( u1_u10_X_33 ) );
  XOR2_X1 u1_u10_U29 (.B( u1_K11_28 ) , .A( u1_R9_19 ) , .Z( u1_u10_X_28 ) );
  XOR2_X1 u1_u10_U30 (.B( u1_K11_27 ) , .A( u1_R9_18 ) , .Z( u1_u10_X_27 ) );
  XOR2_X1 u1_u10_U31 (.B( u1_K11_26 ) , .A( u1_R9_17 ) , .Z( u1_u10_X_26 ) );
  XOR2_X1 u1_u10_U33 (.B( u1_K11_24 ) , .A( u1_R9_17 ) , .Z( u1_u10_X_24 ) );
  XOR2_X1 u1_u10_U36 (.B( u1_K11_21 ) , .A( u1_R9_14 ) , .Z( u1_u10_X_21 ) );
  XOR2_X1 u1_u10_U37 (.B( u1_K11_20 ) , .A( u1_R9_13 ) , .Z( u1_u10_X_20 ) );
  XOR2_X1 u1_u10_U38 (.B( u1_K11_1 ) , .A( u1_R9_32 ) , .Z( u1_u10_X_1 ) );
  XOR2_X1 u1_u10_U4 (.B( u1_K11_6 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_6 ) );
  XOR2_X1 u1_u10_U40 (.B( u1_K11_18 ) , .A( u1_R9_13 ) , .Z( u1_u10_X_18 ) );
  XOR2_X1 u1_u10_U42 (.B( u1_K11_16 ) , .A( u1_R9_11 ) , .Z( u1_u10_X_16 ) );
  XOR2_X1 u1_u10_U43 (.B( u1_K11_15 ) , .A( u1_R9_10 ) , .Z( u1_u10_X_15 ) );
  XOR2_X1 u1_u10_U48 (.B( u1_K11_10 ) , .A( u1_R9_7 ) , .Z( u1_u10_X_10 ) );
  XOR2_X1 u1_u10_U6 (.B( u1_K11_4 ) , .A( u1_R9_3 ) , .Z( u1_u10_X_4 ) );
  XOR2_X1 u1_u10_U8 (.B( u1_K11_47 ) , .A( u1_R9_32 ) , .Z( u1_u10_X_47 ) );
  XOR2_X1 u1_u10_U9 (.B( u1_K11_46 ) , .A( u1_R9_31 ) , .Z( u1_u10_X_46 ) );
  XOR2_X1 u1_u11_U1 (.B( u1_K12_9 ) , .A( u1_R10_6 ) , .Z( u1_u11_X_9 ) );
  XOR2_X1 u1_u11_U10 (.B( u1_K12_45 ) , .A( u1_R10_30 ) , .Z( u1_u11_X_45 ) );
  XOR2_X1 u1_u11_U15 (.B( u1_K12_40 ) , .A( u1_R10_27 ) , .Z( u1_u11_X_40 ) );
  XOR2_X1 u1_u11_U16 (.B( u1_K12_3 ) , .A( u1_R10_2 ) , .Z( u1_u11_X_3 ) );
  XOR2_X1 u1_u11_U17 (.B( u1_K12_39 ) , .A( u1_R10_26 ) , .Z( u1_u11_X_39 ) );
  XOR2_X1 u1_u11_U22 (.B( u1_K12_34 ) , .A( u1_R10_23 ) , .Z( u1_u11_X_34 ) );
  XOR2_X1 u1_u11_U23 (.B( u1_K12_33 ) , .A( u1_R10_22 ) , .Z( u1_u11_X_33 ) );
  XOR2_X1 u1_u11_U24 (.B( u1_K12_32 ) , .A( u1_R10_21 ) , .Z( u1_u11_X_32 ) );
  XOR2_X1 u1_u11_U25 (.B( u1_K12_31 ) , .A( u1_R10_20 ) , .Z( u1_u11_X_31 ) );
  XOR2_X1 u1_u11_U26 (.B( u1_K12_30 ) , .A( u1_R10_21 ) , .Z( u1_u11_X_30 ) );
  XOR2_X1 u1_u11_U28 (.B( u1_K12_29 ) , .A( u1_R10_20 ) , .Z( u1_u11_X_29 ) );
  XOR2_X1 u1_u11_U29 (.B( u1_K12_28 ) , .A( u1_R10_19 ) , .Z( u1_u11_X_28 ) );
  XOR2_X1 u1_u11_U3 (.B( u1_K12_7 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_7 ) );
  XOR2_X1 u1_u11_U30 (.B( u1_K12_27 ) , .A( u1_R10_18 ) , .Z( u1_u11_X_27 ) );
  XOR2_X1 u1_u11_U35 (.B( u1_K12_22 ) , .A( u1_R10_15 ) , .Z( u1_u11_X_22 ) );
  XOR2_X1 u1_u11_U42 (.B( u1_K12_16 ) , .A( u1_R10_11 ) , .Z( u1_u11_X_16 ) );
  XOR2_X1 u1_u11_U44 (.B( u1_K12_14 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_14 ) );
  XOR2_X1 u1_u11_U45 (.B( u1_K12_13 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_13 ) );
  XOR2_X1 u1_u11_U46 (.B( u1_K12_12 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_12 ) );
  XOR2_X1 u1_u11_U47 (.B( u1_K12_11 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_11 ) );
  XOR2_X1 u1_u11_U48 (.B( u1_K12_10 ) , .A( u1_R10_7 ) , .Z( u1_u11_X_10 ) );
  XOR2_X1 u1_u11_U5 (.B( u1_K12_5 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_5 ) );
  XOR2_X1 u1_u11_U6 (.B( u1_K12_4 ) , .A( u1_R10_3 ) , .Z( u1_u11_X_4 ) );
  XOR2_X1 u1_u11_U9 (.B( u1_K12_46 ) , .A( u1_R10_31 ) , .Z( u1_u11_X_46 ) );
  XOR2_X1 u1_u12_U1 (.B( u1_K13_9 ) , .A( u1_R11_6 ) , .Z( u1_u12_X_9 ) );
  XOR2_X1 u1_u12_U10 (.B( u1_K13_45 ) , .A( u1_R11_30 ) , .Z( u1_u12_X_45 ) );
  XOR2_X1 u1_u12_U11 (.B( u1_K13_44 ) , .A( u1_R11_29 ) , .Z( u1_u12_X_44 ) );
  XOR2_X1 u1_u12_U12 (.B( u1_K13_43 ) , .A( u1_R11_28 ) , .Z( u1_u12_X_43 ) );
  XOR2_X1 u1_u12_U13 (.B( u1_K13_42 ) , .A( u1_R11_29 ) , .Z( u1_u12_X_42 ) );
  XOR2_X1 u1_u12_U14 (.B( u1_K13_41 ) , .A( u1_R11_28 ) , .Z( u1_u12_X_41 ) );
  XOR2_X1 u1_u12_U15 (.B( u1_K13_40 ) , .A( u1_R11_27 ) , .Z( u1_u12_X_40 ) );
  XOR2_X1 u1_u12_U16 (.B( u1_K13_3 ) , .A( u1_R11_2 ) , .Z( u1_u12_X_3 ) );
  XOR2_X1 u1_u12_U17 (.B( u1_K13_39 ) , .A( u1_R11_26 ) , .Z( u1_u12_X_39 ) );
  XOR2_X1 u1_u12_U18 (.B( u1_K13_38 ) , .A( u1_R11_25 ) , .Z( u1_u12_X_38 ) );
  XOR2_X1 u1_u12_U20 (.B( u1_K13_36 ) , .A( u1_R11_25 ) , .Z( u1_u12_X_36 ) );
  XOR2_X1 u1_u12_U22 (.B( u1_K13_34 ) , .A( u1_R11_23 ) , .Z( u1_u12_X_34 ) );
  XOR2_X1 u1_u12_U23 (.B( u1_K13_33 ) , .A( u1_R11_22 ) , .Z( u1_u12_X_33 ) );
  XOR2_X1 u1_u12_U29 (.B( u1_K13_28 ) , .A( u1_R11_19 ) , .Z( u1_u12_X_28 ) );
  XOR2_X1 u1_u12_U30 (.B( u1_K13_27 ) , .A( u1_R11_18 ) , .Z( u1_u12_X_27 ) );
  XOR2_X1 u1_u12_U31 (.B( u1_K13_26 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_26 ) );
  XOR2_X1 u1_u12_U32 (.B( u1_K13_25 ) , .A( u1_R11_16 ) , .Z( u1_u12_X_25 ) );
  XOR2_X1 u1_u12_U33 (.B( u1_K13_24 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_24 ) );
  XOR2_X1 u1_u12_U34 (.B( u1_K13_23 ) , .A( u1_R11_16 ) , .Z( u1_u12_X_23 ) );
  XOR2_X1 u1_u12_U35 (.B( u1_K13_22 ) , .A( u1_R11_15 ) , .Z( u1_u12_X_22 ) );
  XOR2_X1 u1_u12_U36 (.B( u1_K13_21 ) , .A( u1_R11_14 ) , .Z( u1_u12_X_21 ) );
  XOR2_X1 u1_u12_U38 (.B( u1_K13_1 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_1 ) );
  XOR2_X1 u1_u12_U42 (.B( u1_K13_16 ) , .A( u1_R11_11 ) , .Z( u1_u12_X_16 ) );
  XOR2_X1 u1_u12_U48 (.B( u1_K13_10 ) , .A( u1_R11_7 ) , .Z( u1_u12_X_10 ) );
  XOR2_X1 u1_u12_U6 (.B( u1_K13_4 ) , .A( u1_R11_3 ) , .Z( u1_u12_X_4 ) );
  XOR2_X1 u1_u12_U8 (.B( u1_K13_47 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_47 ) );
  XOR2_X1 u1_u12_U9 (.B( u1_K13_46 ) , .A( u1_R11_31 ) , .Z( u1_u12_X_46 ) );
  XOR2_X1 u1_u13_U1 (.B( u1_K14_9 ) , .A( u1_R12_6 ) , .Z( u1_u13_X_9 ) );
  XOR2_X1 u1_u13_U10 (.B( u1_K14_45 ) , .A( u1_R12_30 ) , .Z( u1_u13_X_45 ) );
  XOR2_X1 u1_u13_U12 (.B( u1_K14_43 ) , .A( u1_R12_28 ) , .Z( u1_u13_X_43 ) );
  XOR2_X1 u1_u13_U14 (.B( u1_K14_41 ) , .A( u1_R12_28 ) , .Z( u1_u13_X_41 ) );
  XOR2_X1 u1_u13_U15 (.B( u1_K14_40 ) , .A( u1_R12_27 ) , .Z( u1_u13_X_40 ) );
  XOR2_X1 u1_u13_U16 (.B( u1_K14_3 ) , .A( u1_R12_2 ) , .Z( u1_u13_X_3 ) );
  XOR2_X1 u1_u13_U17 (.B( u1_K14_39 ) , .A( u1_R12_26 ) , .Z( u1_u13_X_39 ) );
  XOR2_X1 u1_u13_U18 (.B( u1_K14_38 ) , .A( u1_R12_25 ) , .Z( u1_u13_X_38 ) );
  XOR2_X1 u1_u13_U19 (.B( u1_K14_37 ) , .A( u1_R12_24 ) , .Z( u1_u13_X_37 ) );
  XOR2_X1 u1_u13_U2 (.B( u1_K14_8 ) , .A( u1_R12_5 ) , .Z( u1_u13_X_8 ) );
  XOR2_X1 u1_u13_U20 (.B( u1_K14_36 ) , .A( u1_R12_25 ) , .Z( u1_u13_X_36 ) );
  XOR2_X1 u1_u13_U21 (.B( u1_K14_35 ) , .A( u1_R12_24 ) , .Z( u1_u13_X_35 ) );
  XOR2_X1 u1_u13_U23 (.B( u1_K14_33 ) , .A( u1_R12_22 ) , .Z( u1_u13_X_33 ) );
  XOR2_X1 u1_u13_U29 (.B( u1_K14_28 ) , .A( u1_R12_19 ) , .Z( u1_u13_X_28 ) );
  XOR2_X1 u1_u13_U3 (.B( u1_K14_7 ) , .A( u1_R12_4 ) , .Z( u1_u13_X_7 ) );
  XOR2_X1 u1_u13_U30 (.B( u1_K14_27 ) , .A( u1_R12_18 ) , .Z( u1_u13_X_27 ) );
  XOR2_X1 u1_u13_U31 (.B( u1_K14_26 ) , .A( u1_R12_17 ) , .Z( u1_u13_X_26 ) );
  XOR2_X1 u1_u13_U32 (.B( u1_K14_25 ) , .A( u1_R12_16 ) , .Z( u1_u13_X_25 ) );
  XOR2_X1 u1_u13_U33 (.B( u1_K14_24 ) , .A( u1_R12_17 ) , .Z( u1_u13_X_24 ) );
  XOR2_X1 u1_u13_U34 (.B( u1_K14_23 ) , .A( u1_R12_16 ) , .Z( u1_u13_X_23 ) );
  XOR2_X1 u1_u13_U35 (.B( u1_K14_22 ) , .A( u1_R12_15 ) , .Z( u1_u13_X_22 ) );
  XOR2_X1 u1_u13_U36 (.B( u1_K14_21 ) , .A( u1_R12_14 ) , .Z( u1_u13_X_21 ) );
  XOR2_X1 u1_u13_U37 (.B( u1_K14_20 ) , .A( u1_R12_13 ) , .Z( u1_u13_X_20 ) );
  XOR2_X1 u1_u13_U39 (.B( u1_K14_19 ) , .A( u1_R12_12 ) , .Z( u1_u13_X_19 ) );
  XOR2_X1 u1_u13_U4 (.B( u1_K14_6 ) , .A( u1_R12_5 ) , .Z( u1_u13_X_6 ) );
  XOR2_X1 u1_u13_U40 (.B( u1_K14_18 ) , .A( u1_R12_13 ) , .Z( u1_u13_X_18 ) );
  XOR2_X1 u1_u13_U41 (.B( u1_K14_17 ) , .A( u1_R12_12 ) , .Z( u1_u13_X_17 ) );
  XOR2_X1 u1_u13_U42 (.B( u1_K14_16 ) , .A( u1_R12_11 ) , .Z( u1_u13_X_16 ) );
  XOR2_X1 u1_u13_U43 (.B( u1_K14_15 ) , .A( u1_R12_10 ) , .Z( u1_u13_X_15 ) );
  XOR2_X1 u1_u13_U44 (.B( u1_K14_14 ) , .A( u1_R12_9 ) , .Z( u1_u13_X_14 ) );
  XOR2_X1 u1_u13_U45 (.B( u1_K14_13 ) , .A( u1_R12_8 ) , .Z( u1_u13_X_13 ) );
  XOR2_X1 u1_u13_U46 (.B( u1_K14_12 ) , .A( u1_R12_9 ) , .Z( u1_u13_X_12 ) );
  XOR2_X1 u1_u13_U47 (.B( u1_K14_11 ) , .A( u1_R12_8 ) , .Z( u1_u13_X_11 ) );
  XOR2_X1 u1_u13_U48 (.B( u1_K14_10 ) , .A( u1_R12_7 ) , .Z( u1_u13_X_10 ) );
  XOR2_X1 u1_u13_U5 (.B( u1_K14_5 ) , .A( u1_R12_4 ) , .Z( u1_u13_X_5 ) );
  XOR2_X1 u1_u13_U6 (.B( u1_K14_4 ) , .A( u1_R12_3 ) , .Z( u1_u13_X_4 ) );
  XOR2_X1 u1_u13_U9 (.B( u1_K14_46 ) , .A( u1_R12_31 ) , .Z( u1_u13_X_46 ) );
  XOR2_X1 u1_u14_U1 (.B( u1_K15_9 ) , .A( u1_R13_6 ) , .Z( u1_u14_X_9 ) );
  XOR2_X1 u1_u14_U10 (.B( u1_K15_45 ) , .A( u1_R13_30 ) , .Z( u1_u14_X_45 ) );
  XOR2_X1 u1_u14_U15 (.B( u1_K15_40 ) , .A( u1_R13_27 ) , .Z( u1_u14_X_40 ) );
  XOR2_X1 u1_u14_U16 (.B( u1_K15_3 ) , .A( u1_R13_2 ) , .Z( u1_u14_X_3 ) );
  XOR2_X1 u1_u14_U17 (.B( u1_K15_39 ) , .A( u1_R13_26 ) , .Z( u1_u14_X_39 ) );
  XOR2_X1 u1_u14_U22 (.B( u1_K15_34 ) , .A( u1_R13_23 ) , .Z( u1_u14_X_34 ) );
  XOR2_X1 u1_u14_U23 (.B( u1_K15_33 ) , .A( u1_R13_22 ) , .Z( u1_u14_X_33 ) );
  XOR2_X1 u1_u14_U29 (.B( u1_K15_28 ) , .A( u1_R13_19 ) , .Z( u1_u14_X_28 ) );
  XOR2_X1 u1_u14_U30 (.B( u1_K15_27 ) , .A( u1_R13_18 ) , .Z( u1_u14_X_27 ) );
  XOR2_X1 u1_u14_U35 (.B( u1_K15_22 ) , .A( u1_R13_15 ) , .Z( u1_u14_X_22 ) );
  XOR2_X1 u1_u14_U36 (.B( u1_K15_21 ) , .A( u1_R13_14 ) , .Z( u1_u14_X_21 ) );
  XOR2_X1 u1_u14_U38 (.B( u1_K15_1 ) , .A( u1_R13_32 ) , .Z( u1_u14_X_1 ) );
  XOR2_X1 u1_u14_U39 (.B( u1_K15_19 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_19 ) );
  XOR2_X1 u1_u14_U41 (.B( u1_K15_17 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_17 ) );
  XOR2_X1 u1_u14_U42 (.B( u1_K15_16 ) , .A( u1_R13_11 ) , .Z( u1_u14_X_16 ) );
  XOR2_X1 u1_u14_U43 (.B( u1_K15_15 ) , .A( u1_R13_10 ) , .Z( u1_u14_X_15 ) );
  XOR2_X1 u1_u14_U48 (.B( u1_K15_10 ) , .A( u1_R13_7 ) , .Z( u1_u14_X_10 ) );
  XOR2_X1 u1_u14_U6 (.B( u1_K15_4 ) , .A( u1_R13_3 ) , .Z( u1_u14_X_4 ) );
  XOR2_X1 u1_u14_U8 (.B( u1_K15_47 ) , .A( u1_R13_32 ) , .Z( u1_u14_X_47 ) );
  XOR2_X1 u1_u14_U9 (.B( u1_K15_46 ) , .A( u1_R13_31 ) , .Z( u1_u14_X_46 ) );
  XOR2_X1 u1_u15_U1 (.A( u1_FP_38 ) , .B( u1_K16_9 ) , .Z( u1_u15_X_9 ) );
  XOR2_X1 u1_u15_U10 (.A( u1_FP_62 ) , .B( u1_K16_45 ) , .Z( u1_u15_X_45 ) );
  XOR2_X1 u1_u15_U15 (.A( u1_FP_59 ) , .B( u1_K16_40 ) , .Z( u1_u15_X_40 ) );
  XOR2_X1 u1_u15_U16 (.A( u1_FP_34 ) , .B( u1_K16_3 ) , .Z( u1_u15_X_3 ) );
  XOR2_X1 u1_u15_U17 (.A( u1_FP_58 ) , .B( u1_K16_39 ) , .Z( u1_u15_X_39 ) );
  XOR2_X1 u1_u15_U18 (.A( u1_FP_57 ) , .B( u1_K16_38 ) , .Z( u1_u15_X_38 ) );
  XOR2_X1 u1_u15_U20 (.A( u1_FP_57 ) , .B( u1_K16_36 ) , .Z( u1_u15_X_36 ) );
  XOR2_X1 u1_u15_U23 (.A( u1_FP_54 ) , .B( u1_K16_33 ) , .Z( u1_u15_X_33 ) );
  XOR2_X1 u1_u15_U29 (.A( u1_FP_51 ) , .B( u1_K16_28 ) , .Z( u1_u15_X_28 ) );
  XOR2_X1 u1_u15_U3 (.A( u1_FP_36 ) , .B( u1_K16_7 ) , .Z( u1_u15_X_7 ) );
  XOR2_X1 u1_u15_U30 (.A( u1_FP_50 ) , .B( u1_K16_27 ) , .Z( u1_u15_X_27 ) );
  XOR2_X1 u1_u15_U31 (.A( u1_FP_49 ) , .B( u1_K16_26 ) , .Z( u1_u15_X_26 ) );
  XOR2_X1 u1_u15_U32 (.A( u1_FP_48 ) , .B( u1_K16_25 ) , .Z( u1_u15_X_25 ) );
  XOR2_X1 u1_u15_U33 (.A( u1_FP_49 ) , .B( u1_K16_24 ) , .Z( u1_u15_X_24 ) );
  XOR2_X1 u1_u15_U34 (.A( u1_FP_48 ) , .B( u1_K16_23 ) , .Z( u1_u15_X_23 ) );
  XOR2_X1 u1_u15_U35 (.A( u1_FP_47 ) , .B( u1_K16_22 ) , .Z( u1_u15_X_22 ) );
  XOR2_X1 u1_u15_U36 (.A( u1_FP_46 ) , .B( u1_K16_21 ) , .Z( u1_u15_X_21 ) );
  XOR2_X1 u1_u15_U38 (.A( u1_FP_64 ) , .B( u1_K16_1 ) , .Z( u1_u15_X_1 ) );
  XOR2_X1 u1_u15_U42 (.A( u1_FP_43 ) , .B( u1_K16_16 ) , .Z( u1_u15_X_16 ) );
  XOR2_X1 u1_u15_U43 (.A( u1_FP_42 ) , .B( u1_K16_15 ) , .Z( u1_u15_X_15 ) );
  XOR2_X1 u1_u15_U48 (.A( u1_FP_39 ) , .B( u1_K16_10 ) , .Z( u1_u15_X_10 ) );
  XOR2_X1 u1_u15_U5 (.A( u1_FP_36 ) , .B( u1_K16_5 ) , .Z( u1_u15_X_5 ) );
  XOR2_X1 u1_u15_U6 (.A( u1_FP_35 ) , .B( u1_K16_4 ) , .Z( u1_u15_X_4 ) );
  XOR2_X1 u1_u15_U8 (.A( u1_FP_64 ) , .B( u1_K16_47 ) , .Z( u1_u15_X_47 ) );
  XOR2_X1 u1_u15_U9 (.A( u1_FP_63 ) , .B( u1_K16_46 ) , .Z( u1_u15_X_46 ) );
  XOR2_X1 u1_u1_U1 (.B( u1_K2_9 ) , .A( u1_R0_6 ) , .Z( u1_u1_X_9 ) );
  XOR2_X1 u1_u1_U10 (.B( u1_K2_45 ) , .A( u1_R0_30 ) , .Z( u1_u1_X_45 ) );
  XOR2_X1 u1_u1_U15 (.B( u1_K2_40 ) , .A( u1_R0_27 ) , .Z( u1_u1_X_40 ) );
  XOR2_X1 u1_u1_U16 (.B( u1_K2_3 ) , .A( u1_R0_2 ) , .Z( u1_u1_X_3 ) );
  XOR2_X1 u1_u1_U17 (.B( u1_K2_39 ) , .A( u1_R0_26 ) , .Z( u1_u1_X_39 ) );
  XOR2_X1 u1_u1_U18 (.B( u1_K2_38 ) , .A( u1_R0_25 ) , .Z( u1_u1_X_38 ) );
  XOR2_X1 u1_u1_U19 (.B( u1_K2_37 ) , .A( u1_R0_24 ) , .Z( u1_u1_X_37 ) );
  XOR2_X1 u1_u1_U20 (.B( u1_K2_36 ) , .A( u1_R0_25 ) , .Z( u1_u1_X_36 ) );
  XOR2_X1 u1_u1_U21 (.B( u1_K2_35 ) , .A( u1_R0_24 ) , .Z( u1_u1_X_35 ) );
  XOR2_X1 u1_u1_U22 (.B( u1_K2_34 ) , .A( u1_R0_23 ) , .Z( u1_u1_X_34 ) );
  XOR2_X1 u1_u1_U23 (.B( u1_K2_33 ) , .A( u1_R0_22 ) , .Z( u1_u1_X_33 ) );
  XOR2_X1 u1_u1_U29 (.B( u1_K2_28 ) , .A( u1_R0_19 ) , .Z( u1_u1_X_28 ) );
  XOR2_X1 u1_u1_U30 (.B( u1_K2_27 ) , .A( u1_R0_18 ) , .Z( u1_u1_X_27 ) );
  XOR2_X1 u1_u1_U35 (.B( u1_K2_22 ) , .A( u1_R0_15 ) , .Z( u1_u1_X_22 ) );
  XOR2_X1 u1_u1_U36 (.B( u1_K2_21 ) , .A( u1_R0_14 ) , .Z( u1_u1_X_21 ) );
  XOR2_X1 u1_u1_U42 (.B( u1_K2_16 ) , .A( u1_R0_11 ) , .Z( u1_u1_X_16 ) );
  XOR2_X1 u1_u1_U43 (.B( u1_K2_15 ) , .A( u1_R0_10 ) , .Z( u1_u1_X_15 ) );
  XOR2_X1 u1_u1_U6 (.B( u1_K2_4 ) , .A( u1_R0_3 ) , .Z( u1_u1_X_4 ) );
  XOR2_X1 u1_u1_U9 (.B( u1_K2_46 ) , .A( u1_R0_31 ) , .Z( u1_u1_X_46 ) );
  XOR2_X1 u1_u2_U1 (.B( u1_K3_9 ) , .A( u1_R1_6 ) , .Z( u1_u2_X_9 ) );
  XOR2_X1 u1_u2_U10 (.B( u1_K3_45 ) , .A( u1_R1_30 ) , .Z( u1_u2_X_45 ) );
  XOR2_X1 u1_u2_U15 (.B( u1_K3_40 ) , .A( u1_R1_27 ) , .Z( u1_u2_X_40 ) );
  XOR2_X1 u1_u2_U16 (.B( u1_K3_3 ) , .A( u1_R1_2 ) , .Z( u1_u2_X_3 ) );
  XOR2_X1 u1_u2_U17 (.B( u1_K3_39 ) , .A( u1_R1_26 ) , .Z( u1_u2_X_39 ) );
  XOR2_X1 u1_u2_U22 (.B( u1_K3_34 ) , .A( u1_R1_23 ) , .Z( u1_u2_X_34 ) );
  XOR2_X1 u1_u2_U23 (.B( u1_K3_33 ) , .A( u1_R1_22 ) , .Z( u1_u2_X_33 ) );
  XOR2_X1 u1_u2_U24 (.B( u1_K3_32 ) , .A( u1_R1_21 ) , .Z( u1_u2_X_32 ) );
  XOR2_X1 u1_u2_U26 (.B( u1_K3_30 ) , .A( u1_R1_21 ) , .Z( u1_u2_X_30 ) );
  XOR2_X1 u1_u2_U29 (.B( u1_K3_28 ) , .A( u1_R1_19 ) , .Z( u1_u2_X_28 ) );
  XOR2_X1 u1_u2_U30 (.B( u1_K3_27 ) , .A( u1_R1_18 ) , .Z( u1_u2_X_27 ) );
  XOR2_X1 u1_u2_U35 (.B( u1_K3_22 ) , .A( u1_R1_15 ) , .Z( u1_u2_X_22 ) );
  XOR2_X1 u1_u2_U36 (.B( u1_K3_21 ) , .A( u1_R1_14 ) , .Z( u1_u2_X_21 ) );
  XOR2_X1 u1_u2_U42 (.B( u1_K3_16 ) , .A( u1_R1_11 ) , .Z( u1_u2_X_16 ) );
  XOR2_X1 u1_u2_U43 (.B( u1_K3_15 ) , .A( u1_R1_10 ) , .Z( u1_u2_X_15 ) );
  XOR2_X1 u1_u2_U45 (.B( u1_K3_13 ) , .A( u1_R1_8 ) , .Z( u1_u2_X_13 ) );
  XOR2_X1 u1_u2_U47 (.B( u1_K3_11 ) , .A( u1_R1_8 ) , .Z( u1_u2_X_11 ) );
  XOR2_X1 u1_u2_U48 (.B( u1_K3_10 ) , .A( u1_R1_7 ) , .Z( u1_u2_X_10 ) );
  XOR2_X1 u1_u2_U6 (.B( u1_K3_4 ) , .A( u1_R1_3 ) , .Z( u1_u2_X_4 ) );
  XOR2_X1 u1_u2_U9 (.B( u1_K3_46 ) , .A( u1_R1_31 ) , .Z( u1_u2_X_46 ) );
  XOR2_X1 u1_u3_U1 (.B( u1_K4_9 ) , .A( u1_R2_6 ) , .Z( u1_u3_X_9 ) );
  XOR2_X1 u1_u3_U10 (.B( u1_K4_45 ) , .A( u1_R2_30 ) , .Z( u1_u3_X_45 ) );
  XOR2_X1 u1_u3_U15 (.B( u1_K4_40 ) , .A( u1_R2_27 ) , .Z( u1_u3_X_40 ) );
  XOR2_X1 u1_u3_U17 (.B( u1_K4_39 ) , .A( u1_R2_26 ) , .Z( u1_u3_X_39 ) );
  XOR2_X1 u1_u3_U22 (.B( u1_K4_34 ) , .A( u1_R2_23 ) , .Z( u1_u3_X_34 ) );
  XOR2_X1 u1_u3_U23 (.B( u1_K4_33 ) , .A( u1_R2_22 ) , .Z( u1_u3_X_33 ) );
  XOR2_X1 u1_u3_U29 (.B( u1_K4_28 ) , .A( u1_R2_19 ) , .Z( u1_u3_X_28 ) );
  XOR2_X1 u1_u3_U3 (.B( u1_K4_7 ) , .A( u1_R2_4 ) , .Z( u1_u3_X_7 ) );
  XOR2_X1 u1_u3_U30 (.B( u1_K4_27 ) , .A( u1_R2_18 ) , .Z( u1_u3_X_27 ) );
  XOR2_X1 u1_u3_U35 (.B( u1_K4_22 ) , .A( u1_R2_15 ) , .Z( u1_u3_X_22 ) );
  XOR2_X1 u1_u3_U36 (.B( u1_K4_21 ) , .A( u1_R2_14 ) , .Z( u1_u3_X_21 ) );
  XOR2_X1 u1_u3_U42 (.B( u1_K4_16 ) , .A( u1_R2_11 ) , .Z( u1_u3_X_16 ) );
  XOR2_X1 u1_u3_U43 (.B( u1_K4_15 ) , .A( u1_R2_10 ) , .Z( u1_u3_X_15 ) );
  XOR2_X1 u1_u3_U5 (.B( u1_K4_5 ) , .A( u1_R2_4 ) , .Z( u1_u3_X_5 ) );
  XOR2_X1 u1_u3_U6 (.B( u1_K4_4 ) , .A( u1_R2_3 ) , .Z( u1_u3_X_4 ) );
  XOR2_X1 u1_u3_U9 (.B( u1_K4_46 ) , .A( u1_R2_31 ) , .Z( u1_u3_X_46 ) );
  XOR2_X1 u1_u4_U1 (.B( u1_K5_9 ) , .A( u1_R3_6 ) , .Z( u1_u4_X_9 ) );
  XOR2_X1 u1_u4_U10 (.B( u1_K5_45 ) , .A( u1_R3_30 ) , .Z( u1_u4_X_45 ) );
  XOR2_X1 u1_u4_U15 (.B( u1_K5_40 ) , .A( u1_R3_27 ) , .Z( u1_u4_X_40 ) );
  XOR2_X1 u1_u4_U16 (.B( u1_K5_3 ) , .A( u1_R3_2 ) , .Z( u1_u4_X_3 ) );
  XOR2_X1 u1_u4_U17 (.B( u1_K5_39 ) , .A( u1_R3_26 ) , .Z( u1_u4_X_39 ) );
  XOR2_X1 u1_u4_U22 (.B( u1_K5_34 ) , .A( u1_R3_23 ) , .Z( u1_u4_X_34 ) );
  XOR2_X1 u1_u4_U23 (.B( u1_K5_33 ) , .A( u1_R3_22 ) , .Z( u1_u4_X_33 ) );
  XOR2_X1 u1_u4_U29 (.B( u1_K5_28 ) , .A( u1_R3_19 ) , .Z( u1_u4_X_28 ) );
  XOR2_X1 u1_u4_U36 (.B( u1_K5_21 ) , .A( u1_R3_14 ) , .Z( u1_u4_X_21 ) );
  XOR2_X1 u1_u4_U42 (.B( u1_K5_16 ) , .A( u1_R3_11 ) , .Z( u1_u4_X_16 ) );
  XOR2_X1 u1_u4_U43 (.B( u1_K5_15 ) , .A( u1_R3_10 ) , .Z( u1_u4_X_15 ) );
  XOR2_X1 u1_u4_U48 (.B( u1_K5_10 ) , .A( u1_R3_7 ) , .Z( u1_u4_X_10 ) );
  XOR2_X1 u1_u4_U6 (.B( u1_K5_4 ) , .A( u1_R3_3 ) , .Z( u1_u4_X_4 ) );
  XOR2_X1 u1_u4_U9 (.B( u1_K5_46 ) , .A( u1_R3_31 ) , .Z( u1_u4_X_46 ) );
  XOR2_X1 u1_u5_U10 (.B( u1_K6_45 ) , .A( u1_R4_30 ) , .Z( u1_u5_X_45 ) );
  XOR2_X1 u1_u5_U15 (.B( u1_K6_40 ) , .A( u1_R4_27 ) , .Z( u1_u5_X_40 ) );
  XOR2_X1 u1_u5_U16 (.B( u1_K6_3 ) , .A( u1_R4_2 ) , .Z( u1_u5_X_3 ) );
  XOR2_X1 u1_u5_U17 (.B( u1_K6_39 ) , .A( u1_R4_26 ) , .Z( u1_u5_X_39 ) );
  XOR2_X1 u1_u5_U22 (.B( u1_K6_34 ) , .A( u1_R4_23 ) , .Z( u1_u5_X_34 ) );
  XOR2_X1 u1_u5_U23 (.B( u1_K6_33 ) , .A( u1_R4_22 ) , .Z( u1_u5_X_33 ) );
  XOR2_X1 u1_u5_U29 (.B( u1_K6_28 ) , .A( u1_R4_19 ) , .Z( u1_u5_X_28 ) );
  XOR2_X1 u1_u5_U30 (.B( u1_K6_27 ) , .A( u1_R4_18 ) , .Z( u1_u5_X_27 ) );
  XOR2_X1 u1_u5_U35 (.B( u1_K6_22 ) , .A( u1_R4_15 ) , .Z( u1_u5_X_22 ) );
  XOR2_X1 u1_u5_U39 (.B( u1_K6_19 ) , .A( u1_R4_12 ) , .Z( u1_u5_X_19 ) );
  XOR2_X1 u1_u5_U41 (.B( u1_K6_17 ) , .A( u1_R4_12 ) , .Z( u1_u5_X_17 ) );
  XOR2_X1 u1_u5_U42 (.B( u1_K6_16 ) , .A( u1_R4_11 ) , .Z( u1_u5_X_16 ) );
  XOR2_X1 u1_u5_U43 (.B( u1_K6_15 ) , .A( u1_R4_10 ) , .Z( u1_u5_X_15 ) );
  XOR2_X1 u1_u5_U9 (.B( u1_K6_46 ) , .A( u1_R4_31 ) , .Z( u1_u5_X_46 ) );
  XOR2_X1 u1_u6_U1 (.B( u1_K7_9 ) , .A( u1_R5_6 ) , .Z( u1_u6_X_9 ) );
  XOR2_X1 u1_u6_U10 (.B( u1_K7_45 ) , .A( u1_R5_30 ) , .Z( u1_u6_X_45 ) );
  XOR2_X1 u1_u6_U15 (.B( u1_K7_40 ) , .A( u1_R5_27 ) , .Z( u1_u6_X_40 ) );
  XOR2_X1 u1_u6_U16 (.B( u1_K7_3 ) , .A( u1_R5_2 ) , .Z( u1_u6_X_3 ) );
  XOR2_X1 u1_u6_U17 (.B( u1_K7_39 ) , .A( u1_R5_26 ) , .Z( u1_u6_X_39 ) );
  XOR2_X1 u1_u6_U23 (.B( u1_K7_33 ) , .A( u1_R5_22 ) , .Z( u1_u6_X_33 ) );
  XOR2_X1 u1_u6_U29 (.B( u1_K7_28 ) , .A( u1_R5_19 ) , .Z( u1_u6_X_28 ) );
  XOR2_X1 u1_u6_U35 (.B( u1_K7_22 ) , .A( u1_R5_15 ) , .Z( u1_u6_X_22 ) );
  XOR2_X1 u1_u6_U36 (.B( u1_K7_21 ) , .A( u1_R5_14 ) , .Z( u1_u6_X_21 ) );
  XOR2_X1 u1_u6_U42 (.B( u1_K7_16 ) , .A( u1_R5_11 ) , .Z( u1_u6_X_16 ) );
  XOR2_X1 u1_u6_U43 (.B( u1_K7_15 ) , .A( u1_R5_10 ) , .Z( u1_u6_X_15 ) );
  XOR2_X1 u1_u6_U48 (.B( u1_K7_10 ) , .A( u1_R5_7 ) , .Z( u1_u6_X_10 ) );
  XOR2_X1 u1_u6_U6 (.B( u1_K7_4 ) , .A( u1_R5_3 ) , .Z( u1_u6_X_4 ) );
  XOR2_X1 u1_u7_U1 (.B( u1_K8_9 ) , .A( u1_R6_6 ) , .Z( u1_u7_X_9 ) );
  XOR2_X1 u1_u7_U10 (.B( u1_K8_45 ) , .A( u1_R6_30 ) , .Z( u1_u7_X_45 ) );
  XOR2_X1 u1_u7_U15 (.B( u1_K8_40 ) , .A( u1_R6_27 ) , .Z( u1_u7_X_40 ) );
  XOR2_X1 u1_u7_U17 (.B( u1_K8_39 ) , .A( u1_R6_26 ) , .Z( u1_u7_X_39 ) );
  XOR2_X1 u1_u7_U2 (.B( u1_K8_8 ) , .A( u1_R6_5 ) , .Z( u1_u7_X_8 ) );
  XOR2_X1 u1_u7_U22 (.B( u1_K8_34 ) , .A( u1_R6_23 ) , .Z( u1_u7_X_34 ) );
  XOR2_X1 u1_u7_U23 (.B( u1_K8_33 ) , .A( u1_R6_22 ) , .Z( u1_u7_X_33 ) );
  XOR2_X1 u1_u7_U29 (.B( u1_K8_28 ) , .A( u1_R6_19 ) , .Z( u1_u7_X_28 ) );
  XOR2_X1 u1_u7_U30 (.B( u1_K8_27 ) , .A( u1_R6_18 ) , .Z( u1_u7_X_27 ) );
  XOR2_X1 u1_u7_U35 (.B( u1_K8_22 ) , .A( u1_R6_15 ) , .Z( u1_u7_X_22 ) );
  XOR2_X1 u1_u7_U36 (.B( u1_K8_21 ) , .A( u1_R6_14 ) , .Z( u1_u7_X_21 ) );
  XOR2_X1 u1_u7_U39 (.B( u1_K8_19 ) , .A( u1_R6_12 ) , .Z( u1_u7_X_19 ) );
  XOR2_X1 u1_u7_U4 (.B( u1_K8_6 ) , .A( u1_R6_5 ) , .Z( u1_u7_X_6 ) );
  XOR2_X1 u1_u7_U41 (.B( u1_K8_17 ) , .A( u1_R6_12 ) , .Z( u1_u7_X_17 ) );
  XOR2_X1 u1_u7_U42 (.B( u1_K8_16 ) , .A( u1_R6_11 ) , .Z( u1_u7_X_16 ) );
  XOR2_X1 u1_u7_U48 (.B( u1_K8_10 ) , .A( u1_R6_7 ) , .Z( u1_u7_X_10 ) );
  XOR2_X1 u1_u7_U6 (.B( u1_K8_4 ) , .A( u1_R6_3 ) , .Z( u1_u7_X_4 ) );
  XOR2_X1 u1_u7_U9 (.B( u1_K8_46 ) , .A( u1_R6_31 ) , .Z( u1_u7_X_46 ) );
  XOR2_X1 u1_u8_U10 (.B( u1_K9_45 ) , .A( u1_R7_30 ) , .Z( u1_u8_X_45 ) );
  XOR2_X1 u1_u8_U15 (.B( u1_K9_40 ) , .A( u1_R7_27 ) , .Z( u1_u8_X_40 ) );
  XOR2_X1 u1_u8_U16 (.B( u1_K9_3 ) , .A( u1_R7_2 ) , .Z( u1_u8_X_3 ) );
  XOR2_X1 u1_u8_U17 (.B( u1_K9_39 ) , .A( u1_R7_26 ) , .Z( u1_u8_X_39 ) );
  XOR2_X1 u1_u8_U22 (.B( u1_K9_34 ) , .A( u1_R7_23 ) , .Z( u1_u8_X_34 ) );
  XOR2_X1 u1_u8_U23 (.B( u1_K9_33 ) , .A( u1_R7_22 ) , .Z( u1_u8_X_33 ) );
  XOR2_X1 u1_u8_U24 (.B( u1_K9_32 ) , .A( u1_R7_21 ) , .Z( u1_u8_X_32 ) );
  XOR2_X1 u1_u8_U26 (.B( u1_K9_30 ) , .A( u1_R7_21 ) , .Z( u1_u8_X_30 ) );
  XOR2_X1 u1_u8_U29 (.B( u1_K9_28 ) , .A( u1_R7_19 ) , .Z( u1_u8_X_28 ) );
  XOR2_X1 u1_u8_U36 (.B( u1_K9_21 ) , .A( u1_R7_14 ) , .Z( u1_u8_X_21 ) );
  XOR2_X1 u1_u8_U42 (.B( u1_K9_16 ) , .A( u1_R7_11 ) , .Z( u1_u8_X_16 ) );
  XOR2_X1 u1_u8_U43 (.B( u1_K9_15 ) , .A( u1_R7_10 ) , .Z( u1_u8_X_15 ) );
  XOR2_X1 u1_u8_U6 (.B( u1_K9_4 ) , .A( u1_R7_3 ) , .Z( u1_u8_X_4 ) );
  XOR2_X1 u1_u8_U9 (.B( u1_K9_46 ) , .A( u1_R7_31 ) , .Z( u1_u8_X_46 ) );
  XOR2_X1 u1_u9_U10 (.B( u1_K10_45 ) , .A( u1_R8_30 ) , .Z( u1_u9_X_45 ) );
  XOR2_X1 u1_u9_U15 (.B( u1_K10_40 ) , .A( u1_R8_27 ) , .Z( u1_u9_X_40 ) );
  XOR2_X1 u1_u9_U16 (.B( u1_K10_3 ) , .A( u1_R8_2 ) , .Z( u1_u9_X_3 ) );
  XOR2_X1 u1_u9_U17 (.B( u1_K10_39 ) , .A( u1_R8_26 ) , .Z( u1_u9_X_39 ) );
  XOR2_X1 u1_u9_U22 (.B( u1_K10_34 ) , .A( u1_R8_23 ) , .Z( u1_u9_X_34 ) );
  XOR2_X1 u1_u9_U29 (.B( u1_K10_28 ) , .A( u1_R8_19 ) , .Z( u1_u9_X_28 ) );
  XOR2_X1 u1_u9_U30 (.B( u1_K10_27 ) , .A( u1_R8_18 ) , .Z( u1_u9_X_27 ) );
  XOR2_X1 u1_u9_U36 (.B( u1_K10_21 ) , .A( u1_R8_14 ) , .Z( u1_u9_X_21 ) );
  XOR2_X1 u1_u9_U39 (.B( u1_K10_19 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_19 ) );
  XOR2_X1 u1_u9_U41 (.B( u1_K10_17 ) , .A( u1_R8_12 ) , .Z( u1_u9_X_17 ) );
  XOR2_X1 u1_u9_U42 (.B( u1_K10_16 ) , .A( u1_R8_11 ) , .Z( u1_u9_X_16 ) );
  XOR2_X1 u1_u9_U43 (.B( u1_K10_15 ) , .A( u1_R8_10 ) , .Z( u1_u9_X_15 ) );
  XOR2_X1 u1_u9_U48 (.B( u1_K10_10 ) , .A( u1_R8_7 ) , .Z( u1_u9_X_10 ) );
  XOR2_X1 u1_u9_U6 (.B( u1_K10_4 ) , .A( u1_R8_3 ) , .Z( u1_u9_X_4 ) );
  XOR2_X1 u1_u9_U9 (.B( u1_K10_46 ) , .A( u1_R8_31 ) , .Z( u1_u9_X_46 ) );
  DFF_X1 u1_uk_K_r0_reg_0 (.CK( clk ) , .D( u1_key_r_0 ) , .Q( u1_uk_K_r0_0 ) , .QN( u1_uk_n1260 ) );
  DFF_X1 u1_uk_K_r0_reg_1 (.CK( clk ) , .D( u1_key_r_1 ) , .Q( u1_uk_K_r0_1 ) );
  DFF_X1 u1_uk_K_r0_reg_10 (.CK( clk ) , .D( u1_key_r_10 ) , .Q( u1_uk_K_r0_10 ) , .QN( u1_uk_n1268 ) );
  DFF_X1 u1_uk_K_r0_reg_11 (.CK( clk ) , .D( u1_key_r_11 ) , .Q( u1_uk_K_r0_11 ) );
  DFF_X1 u1_uk_K_r0_reg_12 (.CK( clk ) , .D( u1_key_r_12 ) , .Q( u1_uk_K_r0_12 ) , .QN( u1_uk_n1269 ) );
  DFF_X1 u1_uk_K_r0_reg_13 (.CK( clk ) , .D( u1_key_r_13 ) , .Q( u1_uk_K_r0_13 ) , .QN( u1_uk_n1270 ) );
  DFF_X1 u1_uk_K_r0_reg_14 (.CK( clk ) , .D( u1_key_r_14 ) , .Q( u1_uk_K_r0_14 ) , .QN( u1_uk_n1271 ) );
  DFF_X1 u1_uk_K_r0_reg_15 (.CK( clk ) , .D( u1_key_r_15 ) , .Q( u1_uk_K_r0_15 ) );
  DFF_X1 u1_uk_K_r0_reg_16 (.CK( clk ) , .D( u1_key_r_16 ) , .Q( u1_uk_K_r0_16 ) , .QN( u1_uk_n1272 ) );
  DFF_X1 u1_uk_K_r0_reg_17 (.CK( clk ) , .D( u1_key_r_17 ) , .Q( u1_uk_K_r0_17 ) );
  DFF_X1 u1_uk_K_r0_reg_18 (.CK( clk ) , .D( u1_key_r_18 ) , .Q( u1_uk_K_r0_18 ) , .QN( u1_uk_n1273 ) );
  DFF_X1 u1_uk_K_r0_reg_19 (.CK( clk ) , .D( u1_key_r_19 ) , .Q( u1_uk_K_r0_19 ) );
  DFF_X1 u1_uk_K_r0_reg_2 (.CK( clk ) , .D( u1_key_r_2 ) , .Q( u1_uk_K_r0_2 ) );
  DFF_X1 u1_uk_K_r0_reg_20 (.CK( clk ) , .D( u1_key_r_20 ) , .Q( u1_uk_K_r0_20 ) , .QN( u1_uk_n1274 ) );
  DFF_X1 u1_uk_K_r0_reg_21 (.CK( clk ) , .D( u1_key_r_21 ) , .Q( u1_uk_K_r0_21 ) , .QN( u1_uk_n1275 ) );
  DFF_X1 u1_uk_K_r0_reg_22 (.CK( clk ) , .D( u1_key_r_22 ) , .Q( u1_uk_K_r0_22 ) );
  DFF_X1 u1_uk_K_r0_reg_23 (.CK( clk ) , .D( u1_key_r_23 ) , .Q( u1_uk_K_r0_23 ) , .QN( u1_uk_n1276 ) );
  DFF_X1 u1_uk_K_r0_reg_24 (.CK( clk ) , .D( u1_key_r_24 ) , .Q( u1_uk_K_r0_24 ) , .QN( u1_uk_n1277 ) );
  DFF_X1 u1_uk_K_r0_reg_25 (.CK( clk ) , .D( u1_key_r_25 ) , .Q( u1_uk_K_r0_25 ) );
  DFF_X1 u1_uk_K_r0_reg_26 (.CK( clk ) , .D( u1_key_r_26 ) , .Q( u1_uk_K_r0_26 ) , .QN( u1_uk_n1278 ) );
  DFF_X1 u1_uk_K_r0_reg_27 (.CK( clk ) , .D( u1_key_r_27 ) , .Q( u1_uk_K_r0_27 ) , .QN( u1_uk_n1279 ) );
  DFF_X1 u1_uk_K_r0_reg_28 (.CK( clk ) , .D( u1_key_r_28 ) , .Q( u1_uk_K_r0_28 ) );
  DFF_X1 u1_uk_K_r0_reg_29 (.CK( clk ) , .D( u1_key_r_29 ) , .Q( u1_uk_K_r0_29 ) , .QN( u1_uk_n1281 ) );
  DFF_X1 u1_uk_K_r0_reg_3 (.CK( clk ) , .D( u1_key_r_3 ) , .Q( u1_uk_K_r0_3 ) , .QN( u1_uk_n1261 ) );
  DFF_X1 u1_uk_K_r0_reg_30 (.CK( clk ) , .D( u1_key_r_30 ) , .Q( u1_uk_K_r0_30 ) , .QN( u1_uk_n1282 ) );
  DFF_X1 u1_uk_K_r0_reg_31 (.CK( clk ) , .D( u1_key_r_31 ) , .Q( u1_uk_K_r0_31 ) );
  DFF_X1 u1_uk_K_r0_reg_32 (.CK( clk ) , .D( u1_key_r_32 ) , .Q( u1_uk_K_r0_32 ) );
  DFF_X1 u1_uk_K_r0_reg_33 (.CK( clk ) , .D( u1_key_r_33 ) , .Q( u1_uk_K_r0_33 ) , .QN( u1_uk_n1284 ) );
  DFF_X1 u1_uk_K_r0_reg_34 (.CK( clk ) , .D( u1_key_r_34 ) , .Q( u1_uk_K_r0_34 ) );
  DFF_X1 u1_uk_K_r0_reg_35 (.CK( clk ) , .D( u1_key_r_35 ) , .Q( u1_uk_K_r0_35 ) , .QN( u1_uk_n1286 ) );
  DFF_X1 u1_uk_K_r0_reg_36 (.CK( clk ) , .D( u1_key_r_36 ) , .Q( u1_uk_K_r0_36 ) );
  DFF_X1 u1_uk_K_r0_reg_37 (.CK( clk ) , .D( u1_key_r_37 ) , .Q( u1_uk_K_r0_37 ) , .QN( u1_uk_n1288 ) );
  DFF_X1 u1_uk_K_r0_reg_38 (.CK( clk ) , .D( u1_key_r_38 ) , .Q( u1_uk_K_r0_38 ) , .QN( u1_uk_n1289 ) );
  DFF_X1 u1_uk_K_r0_reg_39 (.CK( clk ) , .D( u1_key_r_39 ) , .Q( u1_uk_K_r0_39 ) , .QN( u1_uk_n1290 ) );
  DFF_X1 u1_uk_K_r0_reg_4 (.CK( clk ) , .D( u1_key_r_4 ) , .Q( u1_uk_K_r0_4 ) , .QN( u1_uk_n1262 ) );
  DFF_X1 u1_uk_K_r0_reg_40 (.CK( clk ) , .D( u1_key_r_40 ) , .Q( u1_uk_K_r0_40 ) , .QN( u1_uk_n1291 ) );
  DFF_X1 u1_uk_K_r0_reg_41 (.CK( clk ) , .D( u1_key_r_41 ) , .Q( u1_uk_K_r0_41 ) , .QN( u1_uk_n1292 ) );
  DFF_X1 u1_uk_K_r0_reg_42 (.CK( clk ) , .D( u1_key_r_42 ) , .Q( u1_uk_K_r0_42 ) , .QN( u1_uk_n1293 ) );
  DFF_X1 u1_uk_K_r0_reg_43 (.CK( clk ) , .D( u1_key_r_43 ) , .Q( u1_uk_K_r0_43 ) , .QN( u1_uk_n1294 ) );
  DFF_X1 u1_uk_K_r0_reg_44 (.CK( clk ) , .D( u1_key_r_44 ) , .Q( u1_uk_K_r0_44 ) , .QN( u1_uk_n1295 ) );
  DFF_X1 u1_uk_K_r0_reg_45 (.CK( clk ) , .D( u1_key_r_45 ) , .Q( u1_uk_K_r0_45 ) , .QN( u1_uk_n1296 ) );
  DFF_X1 u1_uk_K_r0_reg_46 (.CK( clk ) , .D( u1_key_r_46 ) , .Q( u1_uk_K_r0_46 ) , .QN( u1_uk_n1297 ) );
  DFF_X1 u1_uk_K_r0_reg_47 (.CK( clk ) , .D( u1_key_r_47 ) , .Q( u1_uk_K_r0_47 ) , .QN( u1_uk_n1299 ) );
  DFF_X1 u1_uk_K_r0_reg_48 (.CK( clk ) , .D( u1_key_r_48 ) , .Q( u1_uk_K_r0_48 ) , .QN( u1_uk_n1300 ) );
  DFF_X1 u1_uk_K_r0_reg_49 (.CK( clk ) , .D( u1_key_r_49 ) , .Q( u1_uk_K_r0_49 ) );
  DFF_X1 u1_uk_K_r0_reg_5 (.CK( clk ) , .D( u1_key_r_5 ) , .Q( u1_uk_K_r0_5 ) , .QN( u1_uk_n1263 ) );
  DFF_X1 u1_uk_K_r0_reg_50 (.CK( clk ) , .D( u1_key_r_50 ) , .Q( u1_uk_K_r0_50 ) , .QN( u1_uk_n1303 ) );
  DFF_X1 u1_uk_K_r0_reg_51 (.CK( clk ) , .D( u1_key_r_51 ) , .Q( u1_uk_K_r0_51 ) , .QN( u1_uk_n1304 ) );
  DFF_X1 u1_uk_K_r0_reg_52 (.CK( clk ) , .D( u1_key_r_52 ) , .Q( u1_uk_K_r0_52 ) );
  DFF_X1 u1_uk_K_r0_reg_53 (.CK( clk ) , .D( u1_key_r_53 ) , .Q( u1_uk_K_r0_53 ) );
  DFF_X1 u1_uk_K_r0_reg_54 (.CK( clk ) , .D( u1_key_r_54 ) , .Q( u1_uk_K_r0_54 ) , .QN( u1_uk_n1305 ) );
  DFF_X1 u1_uk_K_r0_reg_55 (.CK( clk ) , .D( u1_key_r_55 ) , .Q( u1_uk_K_r0_55 ) );
  DFF_X1 u1_uk_K_r0_reg_6 (.CK( clk ) , .D( u1_key_r_6 ) , .Q( u1_uk_K_r0_6 ) , .QN( u1_uk_n1264 ) );
  DFF_X1 u1_uk_K_r0_reg_7 (.CK( clk ) , .D( u1_key_r_7 ) , .Q( u1_uk_K_r0_7 ) , .QN( u1_uk_n1265 ) );
  DFF_X1 u1_uk_K_r0_reg_8 (.CK( clk ) , .D( u1_key_r_8 ) , .Q( u1_uk_K_r0_8 ) , .QN( u1_uk_n1266 ) );
  DFF_X1 u1_uk_K_r0_reg_9 (.CK( clk ) , .D( u1_key_r_9 ) , .Q( u1_uk_K_r0_9 ) , .QN( u1_uk_n1267 ) );
  DFF_X1 u1_uk_K_r10_reg_0 (.CK( clk ) , .Q( u1_uk_K_r10_0 ) , .D( u1_uk_K_r9_0 ) , .QN( u1_uk_n1708 ) );
  DFF_X1 u1_uk_K_r10_reg_1 (.CK( clk ) , .Q( u1_uk_K_r10_1 ) , .D( u1_uk_K_r9_1 ) , .QN( u1_uk_n1709 ) );
  DFF_X1 u1_uk_K_r10_reg_10 (.CK( clk ) , .Q( u1_uk_K_r10_10 ) , .D( u1_uk_K_r9_10 ) );
  DFF_X1 u1_uk_K_r10_reg_11 (.CK( clk ) , .Q( u1_uk_K_r10_11 ) , .D( u1_uk_K_r9_11 ) );
  DFF_X1 u1_uk_K_r10_reg_12 (.CK( clk ) , .Q( u1_uk_K_r10_12 ) , .D( u1_uk_K_r9_12 ) , .QN( u1_uk_n1716 ) );
  DFF_X1 u1_uk_K_r10_reg_13 (.CK( clk ) , .Q( u1_uk_K_r10_13 ) , .D( u1_uk_K_r9_13 ) );
  DFF_X1 u1_uk_K_r10_reg_14 (.CK( clk ) , .Q( u1_uk_K_r10_14 ) , .D( u1_uk_K_r9_14 ) );
  DFF_X1 u1_uk_K_r10_reg_15 (.CK( clk ) , .Q( u1_uk_K_r10_15 ) , .D( u1_uk_K_r9_15 ) , .QN( u1_uk_n1717 ) );
  DFF_X1 u1_uk_K_r10_reg_16 (.CK( clk ) , .Q( u1_uk_K_r10_16 ) , .D( u1_uk_K_r9_16 ) );
  DFF_X1 u1_uk_K_r10_reg_17 (.CK( clk ) , .Q( u1_uk_K_r10_17 ) , .D( u1_uk_K_r9_17 ) , .QN( u1_uk_n1718 ) );
  DFF_X1 u1_uk_K_r10_reg_18 (.CK( clk ) , .Q( u1_uk_K_r10_18 ) , .D( u1_uk_K_r9_18 ) );
  DFF_X1 u1_uk_K_r10_reg_19 (.CK( clk ) , .Q( u1_uk_K_r10_19 ) , .D( u1_uk_K_r9_19 ) );
  DFF_X1 u1_uk_K_r10_reg_2 (.CK( clk ) , .Q( u1_uk_K_r10_2 ) , .D( u1_uk_K_r9_2 ) , .QN( u1_uk_n1710 ) );
  DFF_X1 u1_uk_K_r10_reg_20 (.CK( clk ) , .Q( u1_uk_K_r10_20 ) , .D( u1_uk_K_r9_20 ) , .QN( u1_uk_n1719 ) );
  DFF_X1 u1_uk_K_r10_reg_21 (.CK( clk ) , .Q( u1_uk_K_r10_21 ) , .D( u1_uk_K_r9_21 ) , .QN( u1_uk_n1720 ) );
  DFF_X1 u1_uk_K_r10_reg_22 (.CK( clk ) , .Q( u1_uk_K_r10_22 ) , .D( u1_uk_K_r9_22 ) , .QN( u1_uk_n1721 ) );
  DFF_X1 u1_uk_K_r10_reg_23 (.CK( clk ) , .Q( u1_uk_K_r10_23 ) , .D( u1_uk_K_r9_23 ) );
  DFF_X1 u1_uk_K_r10_reg_24 (.CK( clk ) , .Q( u1_uk_K_r10_24 ) , .D( u1_uk_K_r9_24 ) , .QN( u1_uk_n1722 ) );
  DFF_X1 u1_uk_K_r10_reg_25 (.CK( clk ) , .Q( u1_uk_K_r10_25 ) , .D( u1_uk_K_r9_25 ) );
  DFF_X1 u1_uk_K_r10_reg_26 (.CK( clk ) , .Q( u1_uk_K_r10_26 ) , .D( u1_uk_K_r9_26 ) , .QN( u1_uk_n1723 ) );
  DFF_X1 u1_uk_K_r10_reg_27 (.CK( clk ) , .Q( u1_uk_K_r10_27 ) , .D( u1_uk_K_r9_27 ) );
  DFF_X1 u1_uk_K_r10_reg_28 (.CK( clk ) , .Q( u1_uk_K_r10_28 ) , .D( u1_uk_K_r9_28 ) );
  DFF_X1 u1_uk_K_r10_reg_29 (.CK( clk ) , .Q( u1_uk_K_r10_29 ) , .D( u1_uk_K_r9_29 ) , .QN( u1_uk_n1728 ) );
  DFF_X1 u1_uk_K_r10_reg_3 (.CK( clk ) , .Q( u1_uk_K_r10_3 ) , .D( u1_uk_K_r9_3 ) , .QN( u1_uk_n1711 ) );
  DFF_X1 u1_uk_K_r10_reg_30 (.CK( clk ) , .Q( u1_uk_K_r10_30 ) , .D( u1_uk_K_r9_30 ) , .QN( u1_uk_n1729 ) );
  DFF_X1 u1_uk_K_r10_reg_31 (.CK( clk ) , .Q( u1_uk_K_r10_31 ) , .D( u1_uk_K_r9_31 ) , .QN( u1_uk_n1730 ) );
  DFF_X1 u1_uk_K_r10_reg_32 (.CK( clk ) , .Q( u1_uk_K_r10_32 ) , .D( u1_uk_K_r9_32 ) , .QN( u1_uk_n1731 ) );
  DFF_X1 u1_uk_K_r10_reg_33 (.CK( clk ) , .Q( u1_uk_K_r10_33 ) , .D( u1_uk_K_r9_33 ) , .QN( u1_uk_n1732 ) );
  DFF_X1 u1_uk_K_r10_reg_34 (.CK( clk ) , .Q( u1_uk_K_r10_34 ) , .D( u1_uk_K_r9_34 ) );
  DFF_X1 u1_uk_K_r10_reg_35 (.CK( clk ) , .Q( u1_uk_K_r10_35 ) , .D( u1_uk_K_r9_35 ) , .QN( u1_uk_n1734 ) );
  DFF_X1 u1_uk_K_r10_reg_36 (.CK( clk ) , .Q( u1_uk_K_r10_36 ) , .D( u1_uk_K_r9_36 ) , .QN( u1_uk_n1735 ) );
  DFF_X1 u1_uk_K_r10_reg_37 (.CK( clk ) , .Q( u1_uk_K_r10_37 ) , .D( u1_uk_K_r9_37 ) , .QN( u1_uk_n1736 ) );
  DFF_X1 u1_uk_K_r10_reg_38 (.CK( clk ) , .Q( u1_uk_K_r10_38 ) , .D( u1_uk_K_r9_38 ) , .QN( u1_uk_n1737 ) );
  DFF_X1 u1_uk_K_r10_reg_39 (.CK( clk ) , .Q( u1_uk_K_r10_39 ) , .D( u1_uk_K_r9_39 ) , .QN( u1_uk_n1738 ) );
  DFF_X1 u1_uk_K_r10_reg_4 (.CK( clk ) , .Q( u1_uk_K_r10_4 ) , .D( u1_uk_K_r9_4 ) );
  DFF_X1 u1_uk_K_r10_reg_40 (.CK( clk ) , .Q( u1_uk_K_r10_40 ) , .D( u1_uk_K_r9_40 ) , .QN( u1_uk_n1739 ) );
  DFF_X1 u1_uk_K_r10_reg_41 (.CK( clk ) , .Q( u1_uk_K_r10_41 ) , .D( u1_uk_K_r9_41 ) );
  DFF_X1 u1_uk_K_r10_reg_42 (.CK( clk ) , .Q( u1_uk_K_r10_42 ) , .D( u1_uk_K_r9_42 ) );
  DFF_X1 u1_uk_K_r10_reg_43 (.CK( clk ) , .Q( u1_uk_K_r10_43 ) , .D( u1_uk_K_r9_43 ) );
  DFF_X1 u1_uk_K_r10_reg_44 (.CK( clk ) , .Q( u1_uk_K_r10_44 ) , .D( u1_uk_K_r9_44 ) );
  DFF_X1 u1_uk_K_r10_reg_45 (.CK( clk ) , .Q( u1_uk_K_r10_45 ) , .D( u1_uk_K_r9_45 ) , .QN( u1_uk_n1744 ) );
  DFF_X1 u1_uk_K_r10_reg_46 (.CK( clk ) , .Q( u1_uk_K_r10_46 ) , .D( u1_uk_K_r9_46 ) , .QN( u1_uk_n1745 ) );
  DFF_X1 u1_uk_K_r10_reg_47 (.CK( clk ) , .Q( u1_uk_K_r10_47 ) , .D( u1_uk_K_r9_47 ) );
  DFF_X1 u1_uk_K_r10_reg_48 (.CK( clk ) , .Q( u1_uk_K_r10_48 ) , .D( u1_uk_K_r9_48 ) );
  DFF_X1 u1_uk_K_r10_reg_49 (.CK( clk ) , .Q( u1_uk_K_r10_49 ) , .D( u1_uk_K_r9_49 ) );
  DFF_X1 u1_uk_K_r10_reg_5 (.CK( clk ) , .Q( u1_uk_K_r10_5 ) , .D( u1_uk_K_r9_5 ) , .QN( u1_uk_n1712 ) );
  DFF_X1 u1_uk_K_r10_reg_50 (.CK( clk ) , .Q( u1_uk_K_r10_50 ) , .D( u1_uk_K_r9_50 ) , .QN( u1_uk_n1748 ) );
  DFF_X1 u1_uk_K_r10_reg_51 (.CK( clk ) , .Q( u1_uk_K_r10_51 ) , .D( u1_uk_K_r9_51 ) , .QN( u1_uk_n1749 ) );
  DFF_X1 u1_uk_K_r10_reg_52 (.CK( clk ) , .Q( u1_uk_K_r10_52 ) , .D( u1_uk_K_r9_52 ) );
  DFF_X1 u1_uk_K_r10_reg_53 (.CK( clk ) , .Q( u1_uk_K_r10_53 ) , .D( u1_uk_K_r9_53 ) , .QN( u1_uk_n1750 ) );
  DFF_X1 u1_uk_K_r10_reg_54 (.CK( clk ) , .Q( u1_uk_K_r10_54 ) , .D( u1_uk_K_r9_54 ) , .QN( u1_uk_n1751 ) );
  DFF_X1 u1_uk_K_r10_reg_55 (.CK( clk ) , .Q( u1_uk_K_r10_55 ) , .D( u1_uk_K_r9_55 ) , .QN( u1_uk_n1752 ) );
  DFF_X1 u1_uk_K_r10_reg_6 (.CK( clk ) , .Q( u1_uk_K_r10_6 ) , .D( u1_uk_K_r9_6 ) , .QN( u1_uk_n1713 ) );
  DFF_X1 u1_uk_K_r10_reg_7 (.CK( clk ) , .Q( u1_uk_K_r10_7 ) , .D( u1_uk_K_r9_7 ) , .QN( u1_uk_n1714 ) );
  DFF_X1 u1_uk_K_r10_reg_8 (.CK( clk ) , .Q( u1_uk_K_r10_8 ) , .D( u1_uk_K_r9_8 ) , .QN( u1_uk_n1715 ) );
  DFF_X1 u1_uk_K_r10_reg_9 (.CK( clk ) , .Q( u1_uk_K_r10_9 ) , .D( u1_uk_K_r9_9 ) );
  DFF_X1 u1_uk_K_r11_reg_0 (.CK( clk ) , .D( u1_uk_K_r10_0 ) , .Q( u1_uk_K_r11_0 ) , .QN( u1_uk_n1753 ) );
  DFF_X1 u1_uk_K_r11_reg_1 (.CK( clk ) , .D( u1_uk_K_r10_1 ) , .Q( u1_uk_K_r11_1 ) , .QN( u1_uk_n1754 ) );
  DFF_X1 u1_uk_K_r11_reg_10 (.CK( clk ) , .D( u1_uk_K_r10_10 ) , .Q( u1_uk_K_r11_10 ) );
  DFF_X1 u1_uk_K_r11_reg_11 (.CK( clk ) , .D( u1_uk_K_r10_11 ) , .Q( u1_uk_K_r11_11 ) );
  DFF_X1 u1_uk_K_r11_reg_12 (.CK( clk ) , .D( u1_uk_K_r10_12 ) , .Q( u1_uk_K_r11_12 ) , .QN( u1_uk_n1761 ) );
  DFF_X1 u1_uk_K_r11_reg_13 (.CK( clk ) , .D( u1_uk_K_r10_13 ) , .Q( u1_uk_K_r11_13 ) , .QN( u1_uk_n1762 ) );
  DFF_X1 u1_uk_K_r11_reg_14 (.CK( clk ) , .D( u1_uk_K_r10_14 ) , .Q( u1_uk_K_r11_14 ) , .QN( u1_uk_n1763 ) );
  DFF_X1 u1_uk_K_r11_reg_15 (.CK( clk ) , .D( u1_uk_K_r10_15 ) , .Q( u1_uk_K_r11_15 ) , .QN( u1_uk_n1764 ) );
  DFF_X1 u1_uk_K_r11_reg_16 (.CK( clk ) , .D( u1_uk_K_r10_16 ) , .Q( u1_uk_K_r11_16 ) , .QN( u1_uk_n1765 ) );
  DFF_X1 u1_uk_K_r11_reg_17 (.CK( clk ) , .D( u1_uk_K_r10_17 ) , .Q( u1_uk_K_r11_17 ) , .QN( u1_uk_n1766 ) );
  DFF_X1 u1_uk_K_r11_reg_18 (.CK( clk ) , .D( u1_uk_K_r10_18 ) , .Q( u1_uk_K_r11_18 ) , .QN( u1_uk_n1767 ) );
  DFF_X1 u1_uk_K_r11_reg_19 (.CK( clk ) , .D( u1_uk_K_r10_19 ) , .Q( u1_uk_K_r11_19 ) );
  DFF_X1 u1_uk_K_r11_reg_2 (.CK( clk ) , .D( u1_uk_K_r10_2 ) , .Q( u1_uk_K_r11_2 ) , .QN( u1_uk_n1755 ) );
  DFF_X1 u1_uk_K_r11_reg_20 (.CK( clk ) , .D( u1_uk_K_r10_20 ) , .Q( u1_uk_K_r11_20 ) );
  DFF_X1 u1_uk_K_r11_reg_21 (.CK( clk ) , .D( u1_uk_K_r10_21 ) , .Q( u1_uk_K_r11_21 ) );
  DFF_X1 u1_uk_K_r11_reg_22 (.CK( clk ) , .D( u1_uk_K_r10_22 ) , .Q( u1_uk_K_r11_22 ) , .QN( u1_uk_n1768 ) );
  DFF_X1 u1_uk_K_r11_reg_23 (.CK( clk ) , .D( u1_uk_K_r10_23 ) , .Q( u1_uk_K_r11_23 ) , .QN( u1_uk_n1769 ) );
  DFF_X1 u1_uk_K_r11_reg_24 (.CK( clk ) , .D( u1_uk_K_r10_24 ) , .Q( u1_uk_K_r11_24 ) );
  DFF_X1 u1_uk_K_r11_reg_25 (.CK( clk ) , .D( u1_uk_K_r10_25 ) , .Q( u1_uk_K_r11_25 ) );
  DFF_X1 u1_uk_K_r11_reg_26 (.CK( clk ) , .D( u1_uk_K_r10_26 ) , .Q( u1_uk_K_r11_26 ) );
  DFF_X1 u1_uk_K_r11_reg_27 (.CK( clk ) , .D( u1_uk_K_r10_27 ) , .Q( u1_uk_K_r11_27 ) );
  DFF_X1 u1_uk_K_r11_reg_28 (.CK( clk ) , .D( u1_uk_K_r10_28 ) , .Q( u1_uk_K_r11_28 ) );
  DFF_X1 u1_uk_K_r11_reg_29 (.CK( clk ) , .D( u1_uk_K_r10_29 ) , .Q( u1_uk_K_r11_29 ) );
  DFF_X1 u1_uk_K_r11_reg_3 (.CK( clk ) , .D( u1_uk_K_r10_3 ) , .Q( u1_uk_K_r11_3 ) , .QN( u1_uk_n1756 ) );
  DFF_X1 u1_uk_K_r11_reg_30 (.CK( clk ) , .D( u1_uk_K_r10_30 ) , .Q( u1_uk_K_r11_30 ) );
  DFF_X1 u1_uk_K_r11_reg_31 (.CK( clk ) , .D( u1_uk_K_r10_31 ) , .Q( u1_uk_K_r11_31 ) , .QN( u1_uk_n1772 ) );
  DFF_X1 u1_uk_K_r11_reg_32 (.CK( clk ) , .D( u1_uk_K_r10_32 ) , .Q( u1_uk_K_r11_32 ) , .QN( u1_uk_n1773 ) );
  DFF_X1 u1_uk_K_r11_reg_33 (.CK( clk ) , .D( u1_uk_K_r10_33 ) , .Q( u1_uk_K_r11_33 ) );
  DFF_X1 u1_uk_K_r11_reg_34 (.CK( clk ) , .D( u1_uk_K_r10_34 ) , .Q( u1_uk_K_r11_34 ) );
  DFF_X1 u1_uk_K_r11_reg_35 (.CK( clk ) , .D( u1_uk_K_r10_35 ) , .Q( u1_uk_K_r11_35 ) , .QN( u1_uk_n1774 ) );
  DFF_X1 u1_uk_K_r11_reg_36 (.CK( clk ) , .D( u1_uk_K_r10_36 ) , .Q( u1_uk_K_r11_36 ) , .QN( u1_uk_n1775 ) );
  DFF_X1 u1_uk_K_r11_reg_37 (.CK( clk ) , .D( u1_uk_K_r10_37 ) , .Q( u1_uk_K_r11_37 ) , .QN( u1_uk_n1776 ) );
  DFF_X1 u1_uk_K_r11_reg_38 (.CK( clk ) , .D( u1_uk_K_r10_38 ) , .Q( u1_uk_K_r11_38 ) , .QN( u1_uk_n1777 ) );
  DFF_X1 u1_uk_K_r11_reg_39 (.CK( clk ) , .D( u1_uk_K_r10_39 ) , .Q( u1_uk_K_r11_39 ) );
  DFF_X1 u1_uk_K_r11_reg_4 (.CK( clk ) , .D( u1_uk_K_r10_4 ) , .Q( u1_uk_K_r11_4 ) );
  DFF_X1 u1_uk_K_r11_reg_40 (.CK( clk ) , .D( u1_uk_K_r10_40 ) , .Q( u1_uk_K_r11_40 ) , .QN( u1_uk_n1780 ) );
  DFF_X1 u1_uk_K_r11_reg_41 (.CK( clk ) , .D( u1_uk_K_r10_41 ) , .Q( u1_uk_K_r11_41 ) , .QN( u1_uk_n1781 ) );
  DFF_X1 u1_uk_K_r11_reg_42 (.CK( clk ) , .D( u1_uk_K_r10_42 ) , .Q( u1_uk_K_r11_42 ) , .QN( u1_uk_n1782 ) );
  DFF_X1 u1_uk_K_r11_reg_43 (.CK( clk ) , .D( u1_uk_K_r10_43 ) , .Q( u1_uk_K_r11_43 ) , .QN( u1_uk_n1783 ) );
  DFF_X1 u1_uk_K_r11_reg_44 (.CK( clk ) , .D( u1_uk_K_r10_44 ) , .Q( u1_uk_K_r11_44 ) , .QN( u1_uk_n1784 ) );
  DFF_X1 u1_uk_K_r11_reg_45 (.CK( clk ) , .D( u1_uk_K_r10_45 ) , .Q( u1_uk_K_r11_45 ) , .QN( u1_uk_n1785 ) );
  DFF_X1 u1_uk_K_r11_reg_46 (.CK( clk ) , .D( u1_uk_K_r10_46 ) , .Q( u1_uk_K_r11_46 ) , .QN( u1_uk_n1787 ) );
  DFF_X1 u1_uk_K_r11_reg_47 (.CK( clk ) , .D( u1_uk_K_r10_47 ) , .Q( u1_uk_K_r11_47 ) );
  DFF_X1 u1_uk_K_r11_reg_48 (.CK( clk ) , .D( u1_uk_K_r10_48 ) , .Q( u1_uk_K_r11_48 ) );
  DFF_X1 u1_uk_K_r11_reg_49 (.CK( clk ) , .D( u1_uk_K_r10_49 ) , .Q( u1_uk_K_r11_49 ) , .QN( u1_uk_n1790 ) );
  DFF_X1 u1_uk_K_r11_reg_5 (.CK( clk ) , .D( u1_uk_K_r10_5 ) , .Q( u1_uk_K_r11_5 ) , .QN( u1_uk_n1757 ) );
  DFF_X1 u1_uk_K_r11_reg_50 (.CK( clk ) , .D( u1_uk_K_r10_50 ) , .Q( u1_uk_K_r11_50 ) , .QN( u1_uk_n1791 ) );
  DFF_X1 u1_uk_K_r11_reg_51 (.CK( clk ) , .D( u1_uk_K_r10_51 ) , .Q( u1_uk_K_r11_51 ) , .QN( u1_uk_n1792 ) );
  DFF_X1 u1_uk_K_r11_reg_52 (.CK( clk ) , .D( u1_uk_K_r10_52 ) , .Q( u1_uk_K_r11_52 ) , .QN( u1_uk_n1793 ) );
  DFF_X1 u1_uk_K_r11_reg_53 (.CK( clk ) , .D( u1_uk_K_r10_53 ) , .Q( u1_uk_K_r11_53 ) );
  DFF_X1 u1_uk_K_r11_reg_54 (.CK( clk ) , .D( u1_uk_K_r10_54 ) , .Q( u1_uk_K_r11_54 ) );
  DFF_X1 u1_uk_K_r11_reg_55 (.CK( clk ) , .D( u1_uk_K_r10_55 ) , .Q( u1_uk_K_r11_55 ) , .QN( u1_uk_n1797 ) );
  DFF_X1 u1_uk_K_r11_reg_6 (.CK( clk ) , .D( u1_uk_K_r10_6 ) , .Q( u1_uk_K_r11_6 ) );
  DFF_X1 u1_uk_K_r11_reg_7 (.CK( clk ) , .D( u1_uk_K_r10_7 ) , .Q( u1_uk_K_r11_7 ) );
  DFF_X1 u1_uk_K_r11_reg_8 (.CK( clk ) , .D( u1_uk_K_r10_8 ) , .Q( u1_uk_K_r11_8 ) );
  DFF_X1 u1_uk_K_r11_reg_9 (.CK( clk ) , .D( u1_uk_K_r10_9 ) , .Q( u1_uk_K_r11_9 ) , .QN( u1_uk_n1758 ) );
  DFF_X1 u1_uk_K_r12_reg_0 (.CK( clk ) , .D( u1_uk_K_r11_0 ) , .Q( u1_uk_K_r12_0 ) , .QN( u1_uk_n1798 ) );
  DFF_X1 u1_uk_K_r12_reg_1 (.CK( clk ) , .D( u1_uk_K_r11_1 ) , .Q( u1_uk_K_r12_1 ) , .QN( u1_uk_n1799 ) );
  DFF_X1 u1_uk_K_r12_reg_10 (.CK( clk ) , .D( u1_uk_K_r11_10 ) , .Q( u1_uk_K_r12_10 ) );
  DFF_X1 u1_uk_K_r12_reg_11 (.CK( clk ) , .D( u1_uk_K_r11_11 ) , .Q( u1_uk_K_r12_11 ) , .QN( u1_uk_n1808 ) );
  DFF_X1 u1_uk_K_r12_reg_12 (.CK( clk ) , .D( u1_uk_K_r11_12 ) , .Q( u1_uk_K_r12_12 ) , .QN( u1_uk_n1809 ) );
  DFF_X1 u1_uk_K_r12_reg_13 (.CK( clk ) , .D( u1_uk_K_r11_13 ) , .Q( u1_uk_K_r12_13 ) , .QN( u1_uk_n1810 ) );
  DFF_X1 u1_uk_K_r12_reg_14 (.CK( clk ) , .D( u1_uk_K_r11_14 ) , .Q( u1_uk_K_r12_14 ) , .QN( u1_uk_n1811 ) );
  DFF_X1 u1_uk_K_r12_reg_15 (.CK( clk ) , .D( u1_uk_K_r11_15 ) , .Q( u1_uk_K_r12_15 ) );
  DFF_X1 u1_uk_K_r12_reg_16 (.CK( clk ) , .D( u1_uk_K_r11_16 ) , .Q( u1_uk_K_r12_16 ) );
  DFF_X1 u1_uk_K_r12_reg_17 (.CK( clk ) , .D( u1_uk_K_r11_17 ) , .Q( u1_uk_K_r12_17 ) , .QN( u1_uk_n1812 ) );
  DFF_X1 u1_uk_K_r12_reg_18 (.CK( clk ) , .D( u1_uk_K_r11_18 ) , .Q( u1_uk_K_r12_18 ) );
  DFF_X1 u1_uk_K_r12_reg_19 (.CK( clk ) , .D( u1_uk_K_r11_19 ) , .Q( u1_uk_K_r12_19 ) , .QN( u1_uk_n1813 ) );
  DFF_X1 u1_uk_K_r12_reg_2 (.CK( clk ) , .D( u1_uk_K_r11_2 ) , .Q( u1_uk_K_r12_2 ) , .QN( u1_uk_n1800 ) );
  DFF_X1 u1_uk_K_r12_reg_20 (.CK( clk ) , .D( u1_uk_K_r11_20 ) , .Q( u1_uk_K_r12_20 ) , .QN( u1_uk_n1814 ) );
  DFF_X1 u1_uk_K_r12_reg_21 (.CK( clk ) , .D( u1_uk_K_r11_21 ) , .Q( u1_uk_K_r12_21 ) );
  DFF_X1 u1_uk_K_r12_reg_22 (.CK( clk ) , .D( u1_uk_K_r11_22 ) , .Q( u1_uk_K_r12_22 ) );
  DFF_X1 u1_uk_K_r12_reg_23 (.CK( clk ) , .D( u1_uk_K_r11_23 ) , .Q( u1_uk_K_r12_23 ) , .QN( u1_uk_n1815 ) );
  DFF_X1 u1_uk_K_r12_reg_24 (.CK( clk ) , .D( u1_uk_K_r11_24 ) , .Q( u1_uk_K_r12_24 ) , .QN( u1_uk_n1816 ) );
  DFF_X1 u1_uk_K_r12_reg_25 (.CK( clk ) , .D( u1_uk_K_r11_25 ) , .Q( u1_uk_K_r12_25 ) , .QN( u1_uk_n1817 ) );
  DFF_X1 u1_uk_K_r12_reg_26 (.CK( clk ) , .D( u1_uk_K_r11_26 ) , .Q( u1_uk_K_r12_26 ) , .QN( u1_uk_n1818 ) );
  DFF_X1 u1_uk_K_r12_reg_27 (.CK( clk ) , .D( u1_uk_K_r11_27 ) , .Q( u1_uk_K_r12_27 ) , .QN( u1_uk_n1819 ) );
  DFF_X1 u1_uk_K_r12_reg_28 (.CK( clk ) , .D( u1_uk_K_r11_28 ) , .Q( u1_uk_K_r12_28 ) , .QN( u1_uk_n1820 ) );
  DFF_X1 u1_uk_K_r12_reg_29 (.CK( clk ) , .D( u1_uk_K_r11_29 ) , .Q( u1_uk_K_r12_29 ) , .QN( u1_uk_n1821 ) );
  DFF_X1 u1_uk_K_r12_reg_3 (.CK( clk ) , .D( u1_uk_K_r11_3 ) , .Q( u1_uk_K_r12_3 ) , .QN( u1_uk_n1801 ) );
  DFF_X1 u1_uk_K_r12_reg_30 (.CK( clk ) , .D( u1_uk_K_r11_30 ) , .Q( u1_uk_K_r12_30 ) , .QN( u1_uk_n1822 ) );
  DFF_X1 u1_uk_K_r12_reg_31 (.CK( clk ) , .D( u1_uk_K_r11_31 ) , .Q( u1_uk_K_r12_31 ) , .QN( u1_uk_n1823 ) );
  DFF_X1 u1_uk_K_r12_reg_32 (.CK( clk ) , .D( u1_uk_K_r11_32 ) , .Q( u1_uk_K_r12_32 ) , .QN( u1_uk_n1824 ) );
  DFF_X1 u1_uk_K_r12_reg_33 (.CK( clk ) , .D( u1_uk_K_r11_33 ) , .Q( u1_uk_K_r12_33 ) );
  DFF_X1 u1_uk_K_r12_reg_34 (.CK( clk ) , .D( u1_uk_K_r11_34 ) , .Q( u1_uk_K_r12_34 ) , .QN( u1_uk_n1826 ) );
  DFF_X1 u1_uk_K_r12_reg_35 (.CK( clk ) , .D( u1_uk_K_r11_35 ) , .Q( u1_uk_K_r12_35 ) , .QN( u1_uk_n1827 ) );
  DFF_X1 u1_uk_K_r12_reg_36 (.CK( clk ) , .D( u1_uk_K_r11_36 ) , .Q( u1_uk_K_r12_36 ) );
  DFF_X1 u1_uk_K_r12_reg_37 (.CK( clk ) , .D( u1_uk_K_r11_37 ) , .Q( u1_uk_K_r12_37 ) , .QN( u1_uk_n1829 ) );
  DFF_X1 u1_uk_K_r12_reg_38 (.CK( clk ) , .D( u1_uk_K_r11_38 ) , .Q( u1_uk_K_r12_38 ) , .QN( u1_uk_n1830 ) );
  DFF_X1 u1_uk_K_r12_reg_39 (.CK( clk ) , .D( u1_uk_K_r11_39 ) , .Q( u1_uk_K_r12_39 ) );
  DFF_X1 u1_uk_K_r12_reg_4 (.CK( clk ) , .D( u1_uk_K_r11_4 ) , .Q( u1_uk_K_r12_4 ) , .QN( u1_uk_n1802 ) );
  DFF_X1 u1_uk_K_r12_reg_40 (.CK( clk ) , .D( u1_uk_K_r11_40 ) , .Q( u1_uk_K_r12_40 ) , .QN( u1_uk_n1831 ) );
  DFF_X1 u1_uk_K_r12_reg_41 (.CK( clk ) , .D( u1_uk_K_r11_41 ) , .Q( u1_uk_K_r12_41 ) );
  DFF_X1 u1_uk_K_r12_reg_42 (.CK( clk ) , .D( u1_uk_K_r11_42 ) , .Q( u1_uk_K_r12_42 ) );
  DFF_X1 u1_uk_K_r12_reg_43 (.CK( clk ) , .D( u1_uk_K_r11_43 ) , .Q( u1_uk_K_r12_43 ) , .QN( u1_uk_n1832 ) );
  DFF_X1 u1_uk_K_r12_reg_44 (.CK( clk ) , .D( u1_uk_K_r11_44 ) , .Q( u1_uk_K_r12_44 ) );
  DFF_X1 u1_uk_K_r12_reg_45 (.CK( clk ) , .D( u1_uk_K_r11_45 ) , .Q( u1_uk_K_r12_45 ) , .QN( u1_uk_n1833 ) );
  DFF_X1 u1_uk_K_r12_reg_46 (.CK( clk ) , .D( u1_uk_K_r11_46 ) , .Q( u1_uk_K_r12_46 ) , .QN( u1_uk_n1834 ) );
  DFF_X1 u1_uk_K_r12_reg_47 (.CK( clk ) , .D( u1_uk_K_r11_47 ) , .Q( u1_uk_K_r12_47 ) );
  DFF_X1 u1_uk_K_r12_reg_48 (.CK( clk ) , .D( u1_uk_K_r11_48 ) , .Q( u1_uk_K_r12_48 ) , .QN( u1_uk_n1835 ) );
  DFF_X1 u1_uk_K_r12_reg_49 (.CK( clk ) , .D( u1_uk_K_r11_49 ) , .Q( u1_uk_K_r12_49 ) , .QN( u1_uk_n1836 ) );
  DFF_X1 u1_uk_K_r12_reg_5 (.CK( clk ) , .D( u1_uk_K_r11_5 ) , .Q( u1_uk_K_r12_5 ) , .QN( u1_uk_n1803 ) );
  DFF_X1 u1_uk_K_r12_reg_50 (.CK( clk ) , .D( u1_uk_K_r11_50 ) , .Q( u1_uk_K_r12_50 ) , .QN( u1_uk_n1837 ) );
  DFF_X1 u1_uk_K_r12_reg_51 (.CK( clk ) , .D( u1_uk_K_r11_51 ) , .Q( u1_uk_K_r12_51 ) , .QN( u1_uk_n1838 ) );
  DFF_X1 u1_uk_K_r12_reg_52 (.CK( clk ) , .D( u1_uk_K_r11_52 ) , .Q( u1_uk_K_r12_52 ) , .QN( u1_uk_n1839 ) );
  DFF_X1 u1_uk_K_r12_reg_53 (.CK( clk ) , .D( u1_uk_K_r11_53 ) , .Q( u1_uk_K_r12_53 ) , .QN( u1_uk_n1840 ) );
  DFF_X1 u1_uk_K_r12_reg_54 (.CK( clk ) , .D( u1_uk_K_r11_54 ) , .Q( u1_uk_K_r12_54 ) , .QN( u1_uk_n1841 ) );
  DFF_X1 u1_uk_K_r12_reg_55 (.CK( clk ) , .D( u1_uk_K_r11_55 ) , .Q( u1_uk_K_r12_55 ) , .QN( u1_uk_n1842 ) );
  DFF_X1 u1_uk_K_r12_reg_6 (.CK( clk ) , .D( u1_uk_K_r11_6 ) , .Q( u1_uk_K_r12_6 ) , .QN( u1_uk_n1804 ) );
  DFF_X1 u1_uk_K_r12_reg_7 (.CK( clk ) , .D( u1_uk_K_r11_7 ) , .Q( u1_uk_K_r12_7 ) );
  DFF_X1 u1_uk_K_r12_reg_8 (.CK( clk ) , .D( u1_uk_K_r11_8 ) , .Q( u1_uk_K_r12_8 ) , .QN( u1_uk_n1806 ) );
  DFF_X1 u1_uk_K_r12_reg_9 (.CK( clk ) , .D( u1_uk_K_r11_9 ) , .Q( u1_uk_K_r12_9 ) , .QN( u1_uk_n1807 ) );
  DFF_X1 u1_uk_K_r13_reg_0 (.CK( clk ) , .D( u1_uk_K_r12_0 ) , .Q( u1_uk_K_r13_0 ) , .QN( u1_uk_n1843 ) );
  DFF_X1 u1_uk_K_r13_reg_1 (.CK( clk ) , .D( u1_uk_K_r12_1 ) , .Q( u1_uk_K_r13_1 ) );
  DFF_X1 u1_uk_K_r13_reg_10 (.CK( clk ) , .D( u1_uk_K_r12_10 ) , .Q( u1_uk_K_r13_10 ) , .QN( u1_uk_n1850 ) );
  DFF_X1 u1_uk_K_r13_reg_11 (.CK( clk ) , .D( u1_uk_K_r12_11 ) , .Q( u1_uk_K_r13_11 ) , .QN( u1_uk_n1851 ) );
  DFF_X1 u1_uk_K_r13_reg_12 (.CK( clk ) , .D( u1_uk_K_r12_12 ) , .Q( u1_uk_K_r13_12 ) , .QN( u1_uk_n1852 ) );
  DFF_X1 u1_uk_K_r13_reg_13 (.CK( clk ) , .D( u1_uk_K_r12_13 ) , .Q( u1_uk_K_r13_13 ) , .QN( u1_uk_n1853 ) );
  DFF_X1 u1_uk_K_r13_reg_14 (.CK( clk ) , .D( u1_uk_K_r12_14 ) , .Q( u1_uk_K_r13_14 ) , .QN( u1_uk_n1854 ) );
  DFF_X1 u1_uk_K_r13_reg_15 (.CK( clk ) , .D( u1_uk_K_r12_15 ) , .Q( u1_uk_K_r13_15 ) , .QN( u1_uk_n1855 ) );
  DFF_X1 u1_uk_K_r13_reg_16 (.CK( clk ) , .D( u1_uk_K_r12_16 ) , .Q( u1_uk_K_r13_16 ) , .QN( u1_uk_n1856 ) );
  DFF_X1 u1_uk_K_r13_reg_17 (.CK( clk ) , .D( u1_uk_K_r12_17 ) , .Q( u1_uk_K_r13_17 ) );
  DFF_X1 u1_uk_K_r13_reg_18 (.CK( clk ) , .D( u1_uk_K_r12_18 ) , .Q( u1_uk_K_r13_18 ) , .QN( u1_uk_n1858 ) );
  DFF_X1 u1_uk_K_r13_reg_19 (.CK( clk ) , .D( u1_uk_K_r12_19 ) , .Q( u1_uk_K_r13_19 ) );
  DFF_X1 u1_uk_K_r13_reg_2 (.CK( clk ) , .D( u1_uk_K_r12_2 ) , .Q( u1_uk_K_r13_2 ) );
  DFF_X1 u1_uk_K_r13_reg_20 (.CK( clk ) , .D( u1_uk_K_r12_20 ) , .Q( u1_uk_K_r13_20 ) , .QN( u1_uk_n1859 ) );
  DFF_X1 u1_uk_K_r13_reg_21 (.CK( clk ) , .D( u1_uk_K_r12_21 ) , .Q( u1_uk_K_r13_21 ) , .QN( u1_uk_n1860 ) );
  DFF_X1 u1_uk_K_r13_reg_22 (.CK( clk ) , .D( u1_uk_K_r12_22 ) , .Q( u1_uk_K_r13_22 ) );
  DFF_X1 u1_uk_K_r13_reg_23 (.CK( clk ) , .D( u1_uk_K_r12_23 ) , .Q( u1_uk_K_r13_23 ) );
  DFF_X1 u1_uk_K_r13_reg_24 (.CK( clk ) , .D( u1_uk_K_r12_24 ) , .Q( u1_uk_K_r13_24 ) , .QN( u1_uk_n1862 ) );
  DFF_X1 u1_uk_K_r13_reg_25 (.CK( clk ) , .D( u1_uk_K_r12_25 ) , .Q( u1_uk_K_r13_25 ) );
  DFF_X1 u1_uk_K_r13_reg_26 (.CK( clk ) , .D( u1_uk_K_r12_26 ) , .Q( u1_uk_K_r13_26 ) , .QN( u1_uk_n1863 ) );
  DFF_X1 u1_uk_K_r13_reg_27 (.CK( clk ) , .D( u1_uk_K_r12_27 ) , .Q( u1_uk_K_r13_27 ) , .QN( u1_uk_n1864 ) );
  DFF_X1 u1_uk_K_r13_reg_28 (.CK( clk ) , .D( u1_uk_K_r12_28 ) , .Q( u1_uk_K_r13_28 ) , .QN( u1_uk_n1865 ) );
  DFF_X1 u1_uk_K_r13_reg_29 (.CK( clk ) , .D( u1_uk_K_r12_29 ) , .Q( u1_uk_K_r13_29 ) , .QN( u1_uk_n1866 ) );
  DFF_X1 u1_uk_K_r13_reg_3 (.CK( clk ) , .D( u1_uk_K_r12_3 ) , .Q( u1_uk_K_r13_3 ) , .QN( u1_uk_n1844 ) );
  DFF_X1 u1_uk_K_r13_reg_30 (.CK( clk ) , .D( u1_uk_K_r12_30 ) , .Q( u1_uk_K_r13_30 ) , .QN( u1_uk_n1867 ) );
  DFF_X1 u1_uk_K_r13_reg_31 (.CK( clk ) , .D( u1_uk_K_r12_31 ) , .Q( u1_uk_K_r13_31 ) );
  DFF_X1 u1_uk_K_r13_reg_32 (.CK( clk ) , .D( u1_uk_K_r12_32 ) , .Q( u1_uk_K_r13_32 ) );
  DFF_X1 u1_uk_K_r13_reg_33 (.CK( clk ) , .D( u1_uk_K_r12_33 ) , .Q( u1_uk_K_r13_33 ) , .QN( u1_uk_n1868 ) );
  DFF_X1 u1_uk_K_r13_reg_34 (.CK( clk ) , .D( u1_uk_K_r12_34 ) , .Q( u1_uk_K_r13_34 ) , .QN( u1_uk_n1869 ) );
  DFF_X1 u1_uk_K_r13_reg_35 (.CK( clk ) , .D( u1_uk_K_r12_35 ) , .Q( u1_uk_K_r13_35 ) );
  DFF_X1 u1_uk_K_r13_reg_36 (.CK( clk ) , .D( u1_uk_K_r12_36 ) , .Q( u1_uk_K_r13_36 ) );
  DFF_X1 u1_uk_K_r13_reg_37 (.CK( clk ) , .D( u1_uk_K_r12_37 ) , .Q( u1_uk_K_r13_37 ) , .QN( u1_uk_n1870 ) );
  DFF_X1 u1_uk_K_r13_reg_38 (.CK( clk ) , .D( u1_uk_K_r12_38 ) , .Q( u1_uk_K_r13_38 ) );
  DFF_X1 u1_uk_K_r13_reg_39 (.CK( clk ) , .D( u1_uk_K_r12_39 ) , .Q( u1_uk_K_r13_39 ) , .QN( u1_uk_n1872 ) );
  DFF_X1 u1_uk_K_r13_reg_4 (.CK( clk ) , .D( u1_uk_K_r12_4 ) , .Q( u1_uk_K_r13_4 ) );
  DFF_X1 u1_uk_K_r13_reg_40 (.CK( clk ) , .D( u1_uk_K_r12_40 ) , .Q( u1_uk_K_r13_40 ) , .QN( u1_uk_n1873 ) );
  DFF_X1 u1_uk_K_r13_reg_41 (.CK( clk ) , .D( u1_uk_K_r12_41 ) , .Q( u1_uk_K_r13_41 ) , .QN( u1_uk_n1874 ) );
  DFF_X1 u1_uk_K_r13_reg_42 (.CK( clk ) , .D( u1_uk_K_r12_42 ) , .Q( u1_uk_K_r13_42 ) , .QN( u1_uk_n1875 ) );
  DFF_X1 u1_uk_K_r13_reg_43 (.CK( clk ) , .D( u1_uk_K_r12_43 ) , .Q( u1_uk_K_r13_43 ) , .QN( u1_uk_n1876 ) );
  DFF_X1 u1_uk_K_r13_reg_44 (.CK( clk ) , .D( u1_uk_K_r12_44 ) , .Q( u1_uk_K_r13_44 ) );
  DFF_X1 u1_uk_K_r13_reg_45 (.CK( clk ) , .D( u1_uk_K_r12_45 ) , .Q( u1_uk_K_r13_45 ) , .QN( u1_uk_n1879 ) );
  DFF_X1 u1_uk_K_r13_reg_46 (.CK( clk ) , .D( u1_uk_K_r12_46 ) , .Q( u1_uk_K_r13_46 ) , .QN( u1_uk_n1880 ) );
  DFF_X1 u1_uk_K_r13_reg_47 (.CK( clk ) , .D( u1_uk_K_r12_47 ) , .Q( u1_uk_K_r13_47 ) , .QN( u1_uk_n1881 ) );
  DFF_X1 u1_uk_K_r13_reg_48 (.CK( clk ) , .D( u1_uk_K_r12_48 ) , .Q( u1_uk_K_r13_48 ) , .QN( u1_uk_n1882 ) );
  DFF_X1 u1_uk_K_r13_reg_49 (.CK( clk ) , .D( u1_uk_K_r12_49 ) , .Q( u1_uk_K_r13_49 ) , .QN( u1_uk_n1883 ) );
  DFF_X1 u1_uk_K_r13_reg_5 (.CK( clk ) , .D( u1_uk_K_r12_5 ) , .Q( u1_uk_K_r13_5 ) , .QN( u1_uk_n1845 ) );
  DFF_X1 u1_uk_K_r13_reg_50 (.CK( clk ) , .D( u1_uk_K_r12_50 ) , .Q( u1_uk_K_r13_50 ) , .QN( u1_uk_n1884 ) );
  DFF_X1 u1_uk_K_r13_reg_51 (.CK( clk ) , .D( u1_uk_K_r12_51 ) , .Q( u1_uk_K_r13_51 ) , .QN( u1_uk_n1885 ) );
  DFF_X1 u1_uk_K_r13_reg_52 (.CK( clk ) , .D( u1_uk_K_r12_52 ) , .Q( u1_uk_K_r13_52 ) , .QN( u1_uk_n1886 ) );
  DFF_X1 u1_uk_K_r13_reg_53 (.CK( clk ) , .D( u1_uk_K_r12_53 ) , .Q( u1_uk_K_r13_53 ) );
  DFF_X1 u1_uk_K_r13_reg_54 (.CK( clk ) , .D( u1_uk_K_r12_54 ) , .Q( u1_uk_K_r13_54 ) , .QN( u1_uk_n1887 ) );
  DFF_X1 u1_uk_K_r13_reg_55 (.CK( clk ) , .D( u1_uk_K_r12_55 ) , .Q( u1_uk_K_r13_55 ) );
  DFF_X1 u1_uk_K_r13_reg_6 (.CK( clk ) , .D( u1_uk_K_r12_6 ) , .Q( u1_uk_K_r13_6 ) , .QN( u1_uk_n1846 ) );
  DFF_X1 u1_uk_K_r13_reg_7 (.CK( clk ) , .D( u1_uk_K_r12_7 ) , .Q( u1_uk_K_r13_7 ) , .QN( u1_uk_n1847 ) );
  DFF_X1 u1_uk_K_r13_reg_8 (.CK( clk ) , .D( u1_uk_K_r12_8 ) , .Q( u1_uk_K_r13_8 ) , .QN( u1_uk_n1848 ) );
  DFF_X1 u1_uk_K_r13_reg_9 (.CK( clk ) , .D( u1_uk_K_r12_9 ) , .Q( u1_uk_K_r13_9 ) , .QN( u1_uk_n1849 ) );
  DFF_X1 u1_uk_K_r14_reg_0 (.CK( clk ) , .D( u1_uk_K_r13_0 ) , .QN( u1_uk_n1218 ) );
  DFF_X1 u1_uk_K_r14_reg_1 (.CK( clk ) , .D( u1_uk_K_r13_1 ) , .QN( u1_uk_n1219 ) );
  DFF_X1 u1_uk_K_r14_reg_10 (.CK( clk ) , .D( u1_uk_K_r13_10 ) , .Q( u1_uk_K_r14_10 ) );
  DFF_X1 u1_uk_K_r14_reg_11 (.CK( clk ) , .D( u1_uk_K_r13_11 ) , .Q( u1_uk_K_r14_11 ) );
  DFF_X1 u1_uk_K_r14_reg_12 (.CK( clk ) , .D( u1_uk_K_r13_12 ) , .Q( u1_uk_K_r14_12 ) );
  DFF_X1 u1_uk_K_r14_reg_13 (.CK( clk ) , .D( u1_uk_K_r13_13 ) , .QN( u1_uk_n1224 ) );
  DFF_X1 u1_uk_K_r14_reg_14 (.CK( clk ) , .D( u1_uk_K_r13_14 ) , .QN( u1_uk_n1225 ) );
  DFF_X1 u1_uk_K_r14_reg_15 (.CK( clk ) , .D( u1_uk_K_r13_15 ) , .Q( u1_uk_K_r14_15 ) );
  DFF_X1 u1_uk_K_r14_reg_16 (.CK( clk ) , .D( u1_uk_K_r13_16 ) , .Q( u1_uk_K_r14_16 ) );
  DFF_X1 u1_uk_K_r14_reg_17 (.CK( clk ) , .D( u1_uk_K_r13_17 ) , .QN( u1_uk_n1227 ) );
  DFF_X1 u1_uk_K_r14_reg_18 (.CK( clk ) , .D( u1_uk_K_r13_18 ) , .Q( u1_uk_K_r14_18 ) );
  DFF_X1 u1_uk_K_r14_reg_19 (.CK( clk ) , .D( u1_uk_K_r13_19 ) , .QN( u1_uk_n1228 ) );
  DFF_X1 u1_uk_K_r14_reg_2 (.CK( clk ) , .D( u1_uk_K_r13_2 ) , .Q( u1_uk_K_r14_2 ) );
  DFF_X1 u1_uk_K_r14_reg_20 (.CK( clk ) , .D( u1_uk_K_r13_20 ) , .QN( u1_uk_n1229 ) );
  DFF_X1 u1_uk_K_r14_reg_21 (.CK( clk ) , .D( u1_uk_K_r13_21 ) , .QN( u1_uk_n1230 ) );
  DFF_X1 u1_uk_K_r14_reg_22 (.CK( clk ) , .D( u1_uk_K_r13_22 ) , .QN( u1_uk_n1231 ) );
  DFF_X1 u1_uk_K_r14_reg_23 (.CK( clk ) , .D( u1_uk_K_r13_23 ) , .Q( u1_uk_K_r14_23 ) , .QN( u1_uk_n1233 ) );
  DFF_X1 u1_uk_K_r14_reg_24 (.CK( clk ) , .D( u1_uk_K_r13_24 ) , .QN( u1_uk_n1234 ) );
  DFF_X1 u1_uk_K_r14_reg_25 (.CK( clk ) , .D( u1_uk_K_r13_25 ) , .QN( u1_uk_n1235 ) );
  DFF_X1 u1_uk_K_r14_reg_26 (.CK( clk ) , .D( u1_uk_K_r13_26 ) , .QN( u1_uk_n1236 ) );
  DFF_X1 u1_uk_K_r14_reg_27 (.CK( clk ) , .D( u1_uk_K_r13_27 ) , .QN( u1_uk_n1237 ) );
  DFF_X1 u1_uk_K_r14_reg_28 (.CK( clk ) , .D( u1_uk_K_r13_28 ) , .QN( u1_uk_n1238 ) );
  DFF_X1 u1_uk_K_r14_reg_29 (.CK( clk ) , .D( u1_uk_K_r13_29 ) , .QN( u1_uk_n1239 ) );
  DFF_X1 u1_uk_K_r14_reg_3 (.CK( clk ) , .D( u1_uk_K_r13_3 ) , .Q( u1_uk_K_r14_3 ) );
  DFF_X1 u1_uk_K_r14_reg_30 (.CK( clk ) , .D( u1_uk_K_r13_30 ) , .QN( u1_uk_n1240 ) );
  DFF_X1 u1_uk_K_r14_reg_31 (.CK( clk ) , .D( u1_uk_K_r13_31 ) , .QN( u1_uk_n1241 ) );
  DFF_X1 u1_uk_K_r14_reg_32 (.CK( clk ) , .D( u1_uk_K_r13_32 ) , .QN( u1_uk_n1242 ) );
  DFF_X1 u1_uk_K_r14_reg_33 (.CK( clk ) , .D( u1_uk_K_r13_33 ) , .QN( u1_uk_n1243 ) );
  DFF_X1 u1_uk_K_r14_reg_34 (.CK( clk ) , .D( u1_uk_K_r13_34 ) , .QN( u1_uk_n1244 ) );
  DFF_X1 u1_uk_K_r14_reg_35 (.CK( clk ) , .D( u1_uk_K_r13_35 ) , .QN( u1_uk_n1245 ) );
  DFF_X1 u1_uk_K_r14_reg_36 (.CK( clk ) , .D( u1_uk_K_r13_36 ) , .QN( u1_uk_n1246 ) );
  DFF_X1 u1_uk_K_r14_reg_37 (.CK( clk ) , .D( u1_uk_K_r13_37 ) , .QN( u1_uk_n1247 ) );
  DFF_X1 u1_uk_K_r14_reg_38 (.CK( clk ) , .D( u1_uk_K_r13_38 ) , .Q( u1_uk_K_r14_38 ) );
  DFF_X1 u1_uk_K_r14_reg_39 (.CK( clk ) , .D( u1_uk_K_r13_39 ) , .Q( u1_uk_K_r14_39 ) );
  DFF_X1 u1_uk_K_r14_reg_4 (.CK( clk ) , .D( u1_uk_K_r13_4 ) , .QN( u1_uk_n1220 ) );
  DFF_X1 u1_uk_K_r14_reg_40 (.CK( clk ) , .D( u1_uk_K_r13_40 ) , .QN( u1_uk_n1248 ) );
  DFF_X1 u1_uk_K_r14_reg_41 (.CK( clk ) , .D( u1_uk_K_r13_41 ) , .QN( u1_uk_n1249 ) );
  DFF_X1 u1_uk_K_r14_reg_42 (.CK( clk ) , .D( u1_uk_K_r13_42 ) , .Q( u1_uk_K_r14_42 ) );
  DFF_X1 u1_uk_K_r14_reg_43 (.CK( clk ) , .D( u1_uk_K_r13_43 ) , .Q( u1_uk_K_r14_43 ) );
  DFF_X1 u1_uk_K_r14_reg_44 (.CK( clk ) , .D( u1_uk_K_r13_44 ) , .QN( u1_uk_n1250 ) );
  DFF_X1 u1_uk_K_r14_reg_45 (.CK( clk ) , .D( u1_uk_K_r13_45 ) , .Q( u1_uk_K_r14_45 ) );
  DFF_X1 u1_uk_K_r14_reg_46 (.CK( clk ) , .D( u1_uk_K_r13_46 ) , .Q( u1_uk_K_r14_46 ) );
  DFF_X1 u1_uk_K_r14_reg_47 (.CK( clk ) , .D( u1_uk_K_r13_47 ) , .QN( u1_uk_n1251 ) );
  DFF_X1 u1_uk_K_r14_reg_48 (.CK( clk ) , .D( u1_uk_K_r13_48 ) , .QN( u1_uk_n1252 ) );
  DFF_X1 u1_uk_K_r14_reg_49 (.CK( clk ) , .D( u1_uk_K_r13_49 ) , .QN( u1_uk_n1253 ) );
  DFF_X1 u1_uk_K_r14_reg_5 (.CK( clk ) , .D( u1_uk_K_r13_5 ) , .Q( u1_uk_K_r14_5 ) );
  DFF_X1 u1_uk_K_r14_reg_50 (.CK( clk ) , .D( u1_uk_K_r13_50 ) , .Q( u1_uk_K_r14_50 ) );
  DFF_X1 u1_uk_K_r14_reg_51 (.CK( clk ) , .D( u1_uk_K_r13_51 ) , .QN( u1_uk_n1255 ) );
  DFF_X1 u1_uk_K_r14_reg_52 (.CK( clk ) , .D( u1_uk_K_r13_52 ) , .QN( u1_uk_n1256 ) );
  DFF_X1 u1_uk_K_r14_reg_53 (.CK( clk ) , .D( u1_uk_K_r13_53 ) , .QN( u1_uk_n1257 ) );
  DFF_X1 u1_uk_K_r14_reg_54 (.CK( clk ) , .D( u1_uk_K_r13_54 ) , .QN( u1_uk_n1258 ) );
  DFF_X1 u1_uk_K_r14_reg_55 (.CK( clk ) , .D( u1_uk_K_r13_55 ) , .QN( u1_uk_n1259 ) );
  DFF_X1 u1_uk_K_r14_reg_6 (.CK( clk ) , .D( u1_uk_K_r13_6 ) , .QN( u1_uk_n1221 ) );
  DFF_X1 u1_uk_K_r14_reg_7 (.CK( clk ) , .D( u1_uk_K_r13_7 ) , .QN( u1_uk_n1222 ) );
  DFF_X1 u1_uk_K_r14_reg_8 (.CK( clk ) , .D( u1_uk_K_r13_8 ) , .Q( u1_uk_K_r14_8 ) );
  DFF_X1 u1_uk_K_r14_reg_9 (.CK( clk ) , .D( u1_uk_K_r13_9 ) , .Q( u1_uk_K_r14_9 ) );
  DFF_X1 u1_uk_K_r1_reg_0 (.CK( clk ) , .D( u1_uk_K_r0_0 ) , .Q( u1_uk_K_r1_0 ) , .QN( u1_uk_n1307 ) );
  DFF_X1 u1_uk_K_r1_reg_1 (.CK( clk ) , .D( u1_uk_K_r0_1 ) , .Q( u1_uk_K_r1_1 ) , .QN( u1_uk_n1308 ) );
  DFF_X1 u1_uk_K_r1_reg_10 (.CK( clk ) , .D( u1_uk_K_r0_10 ) , .Q( u1_uk_K_r1_10 ) );
  DFF_X1 u1_uk_K_r1_reg_11 (.CK( clk ) , .D( u1_uk_K_r0_11 ) , .Q( u1_uk_K_r1_11 ) , .QN( u1_uk_n1315 ) );
  DFF_X1 u1_uk_K_r1_reg_12 (.CK( clk ) , .D( u1_uk_K_r0_12 ) , .Q( u1_uk_K_r1_12 ) , .QN( u1_uk_n1316 ) );
  DFF_X1 u1_uk_K_r1_reg_13 (.CK( clk ) , .D( u1_uk_K_r0_13 ) , .Q( u1_uk_K_r1_13 ) , .QN( u1_uk_n1317 ) );
  DFF_X1 u1_uk_K_r1_reg_14 (.CK( clk ) , .D( u1_uk_K_r0_14 ) , .Q( u1_uk_K_r1_14 ) , .QN( u1_uk_n1318 ) );
  DFF_X1 u1_uk_K_r1_reg_15 (.CK( clk ) , .D( u1_uk_K_r0_15 ) , .Q( u1_uk_K_r1_15 ) );
  DFF_X1 u1_uk_K_r1_reg_16 (.CK( clk ) , .D( u1_uk_K_r0_16 ) , .Q( u1_uk_K_r1_16 ) );
  DFF_X1 u1_uk_K_r1_reg_17 (.CK( clk ) , .D( u1_uk_K_r0_17 ) , .Q( u1_uk_K_r1_17 ) , .QN( u1_uk_n1319 ) );
  DFF_X1 u1_uk_K_r1_reg_18 (.CK( clk ) , .D( u1_uk_K_r0_18 ) , .Q( u1_uk_K_r1_18 ) );
  DFF_X1 u1_uk_K_r1_reg_19 (.CK( clk ) , .D( u1_uk_K_r0_19 ) , .Q( u1_uk_K_r1_19 ) , .QN( u1_uk_n1320 ) );
  DFF_X1 u1_uk_K_r1_reg_2 (.CK( clk ) , .D( u1_uk_K_r0_2 ) , .Q( u1_uk_K_r1_2 ) , .QN( u1_uk_n1309 ) );
  DFF_X1 u1_uk_K_r1_reg_20 (.CK( clk ) , .D( u1_uk_K_r0_20 ) , .Q( u1_uk_K_r1_20 ) , .QN( u1_uk_n1321 ) );
  DFF_X1 u1_uk_K_r1_reg_21 (.CK( clk ) , .D( u1_uk_K_r0_21 ) , .Q( u1_uk_K_r1_21 ) );
  DFF_X1 u1_uk_K_r1_reg_22 (.CK( clk ) , .D( u1_uk_K_r0_22 ) , .Q( u1_uk_K_r1_22 ) );
  DFF_X1 u1_uk_K_r1_reg_23 (.CK( clk ) , .D( u1_uk_K_r0_23 ) , .Q( u1_uk_K_r1_23 ) , .QN( u1_uk_n1322 ) );
  DFF_X1 u1_uk_K_r1_reg_24 (.CK( clk ) , .D( u1_uk_K_r0_24 ) , .Q( u1_uk_K_r1_24 ) , .QN( u1_uk_n1323 ) );
  DFF_X1 u1_uk_K_r1_reg_25 (.CK( clk ) , .D( u1_uk_K_r0_25 ) , .Q( u1_uk_K_r1_25 ) , .QN( u1_uk_n1324 ) );
  DFF_X1 u1_uk_K_r1_reg_26 (.CK( clk ) , .D( u1_uk_K_r0_26 ) , .Q( u1_uk_K_r1_26 ) , .QN( u1_uk_n1325 ) );
  DFF_X1 u1_uk_K_r1_reg_27 (.CK( clk ) , .D( u1_uk_K_r0_27 ) , .Q( u1_uk_K_r1_27 ) , .QN( u1_uk_n1326 ) );
  DFF_X1 u1_uk_K_r1_reg_28 (.CK( clk ) , .D( u1_uk_K_r0_28 ) , .Q( u1_uk_K_r1_28 ) , .QN( u1_uk_n1327 ) );
  DFF_X1 u1_uk_K_r1_reg_29 (.CK( clk ) , .D( u1_uk_K_r0_29 ) , .Q( u1_uk_K_r1_29 ) , .QN( u1_uk_n1328 ) );
  DFF_X1 u1_uk_K_r1_reg_3 (.CK( clk ) , .D( u1_uk_K_r0_3 ) , .Q( u1_uk_K_r1_3 ) , .QN( u1_uk_n1310 ) );
  DFF_X1 u1_uk_K_r1_reg_30 (.CK( clk ) , .D( u1_uk_K_r0_30 ) , .Q( u1_uk_K_r1_30 ) , .QN( u1_uk_n1329 ) );
  DFF_X1 u1_uk_K_r1_reg_31 (.CK( clk ) , .D( u1_uk_K_r0_31 ) , .Q( u1_uk_K_r1_31 ) , .QN( u1_uk_n1330 ) );
  DFF_X1 u1_uk_K_r1_reg_32 (.CK( clk ) , .D( u1_uk_K_r0_32 ) , .Q( u1_uk_K_r1_32 ) , .QN( u1_uk_n1331 ) );
  DFF_X1 u1_uk_K_r1_reg_33 (.CK( clk ) , .D( u1_uk_K_r0_33 ) , .Q( u1_uk_K_r1_33 ) );
  DFF_X1 u1_uk_K_r1_reg_34 (.CK( clk ) , .D( u1_uk_K_r0_34 ) , .Q( u1_uk_K_r1_34 ) , .QN( u1_uk_n1332 ) );
  DFF_X1 u1_uk_K_r1_reg_35 (.CK( clk ) , .D( u1_uk_K_r0_35 ) , .Q( u1_uk_K_r1_35 ) , .QN( u1_uk_n1333 ) );
  DFF_X1 u1_uk_K_r1_reg_36 (.CK( clk ) , .D( u1_uk_K_r0_36 ) , .Q( u1_uk_K_r1_36 ) );
  DFF_X1 u1_uk_K_r1_reg_37 (.CK( clk ) , .D( u1_uk_K_r0_37 ) , .Q( u1_uk_K_r1_37 ) , .QN( u1_uk_n1334 ) );
  DFF_X1 u1_uk_K_r1_reg_38 (.CK( clk ) , .D( u1_uk_K_r0_38 ) , .Q( u1_uk_K_r1_38 ) , .QN( u1_uk_n1335 ) );
  DFF_X1 u1_uk_K_r1_reg_39 (.CK( clk ) , .D( u1_uk_K_r0_39 ) , .Q( u1_uk_K_r1_39 ) );
  DFF_X1 u1_uk_K_r1_reg_4 (.CK( clk ) , .D( u1_uk_K_r0_4 ) , .Q( u1_uk_K_r1_4 ) , .QN( u1_uk_n1311 ) );
  DFF_X1 u1_uk_K_r1_reg_40 (.CK( clk ) , .D( u1_uk_K_r0_40 ) , .Q( u1_uk_K_r1_40 ) , .QN( u1_uk_n1336 ) );
  DFF_X1 u1_uk_K_r1_reg_41 (.CK( clk ) , .D( u1_uk_K_r0_41 ) , .Q( u1_uk_K_r1_41 ) );
  DFF_X1 u1_uk_K_r1_reg_42 (.CK( clk ) , .D( u1_uk_K_r0_42 ) , .Q( u1_uk_K_r1_42 ) );
  DFF_X1 u1_uk_K_r1_reg_43 (.CK( clk ) , .D( u1_uk_K_r0_43 ) , .Q( u1_uk_K_r1_43 ) , .QN( u1_uk_n1338 ) );
  DFF_X1 u1_uk_K_r1_reg_44 (.CK( clk ) , .D( u1_uk_K_r0_44 ) , .Q( u1_uk_K_r1_44 ) );
  DFF_X1 u1_uk_K_r1_reg_45 (.CK( clk ) , .D( u1_uk_K_r0_45 ) , .Q( u1_uk_K_r1_45 ) , .QN( u1_uk_n1339 ) );
  DFF_X1 u1_uk_K_r1_reg_46 (.CK( clk ) , .D( u1_uk_K_r0_46 ) , .Q( u1_uk_K_r1_46 ) , .QN( u1_uk_n1340 ) );
  DFF_X1 u1_uk_K_r1_reg_47 (.CK( clk ) , .D( u1_uk_K_r0_47 ) , .Q( u1_uk_K_r1_47 ) );
  DFF_X1 u1_uk_K_r1_reg_48 (.CK( clk ) , .D( u1_uk_K_r0_48 ) , .Q( u1_uk_K_r1_48 ) , .QN( u1_uk_n1341 ) );
  DFF_X1 u1_uk_K_r1_reg_49 (.CK( clk ) , .D( u1_uk_K_r0_49 ) , .Q( u1_uk_K_r1_49 ) , .QN( u1_uk_n1342 ) );
  DFF_X1 u1_uk_K_r1_reg_5 (.CK( clk ) , .D( u1_uk_K_r0_5 ) , .Q( u1_uk_K_r1_5 ) , .QN( u1_uk_n1312 ) );
  DFF_X1 u1_uk_K_r1_reg_50 (.CK( clk ) , .D( u1_uk_K_r0_50 ) , .Q( u1_uk_K_r1_50 ) , .QN( u1_uk_n1343 ) );
  DFF_X1 u1_uk_K_r1_reg_51 (.CK( clk ) , .D( u1_uk_K_r0_51 ) , .Q( u1_uk_K_r1_51 ) , .QN( u1_uk_n1344 ) );
  DFF_X1 u1_uk_K_r1_reg_52 (.CK( clk ) , .D( u1_uk_K_r0_52 ) , .Q( u1_uk_K_r1_52 ) , .QN( u1_uk_n1345 ) );
  DFF_X1 u1_uk_K_r1_reg_53 (.CK( clk ) , .D( u1_uk_K_r0_53 ) , .Q( u1_uk_K_r1_53 ) , .QN( u1_uk_n1346 ) );
  DFF_X1 u1_uk_K_r1_reg_54 (.CK( clk ) , .D( u1_uk_K_r0_54 ) , .Q( u1_uk_K_r1_54 ) , .QN( u1_uk_n1347 ) );
  DFF_X1 u1_uk_K_r1_reg_55 (.CK( clk ) , .D( u1_uk_K_r0_55 ) , .Q( u1_uk_K_r1_55 ) , .QN( u1_uk_n1348 ) );
  DFF_X1 u1_uk_K_r1_reg_6 (.CK( clk ) , .D( u1_uk_K_r0_6 ) , .Q( u1_uk_K_r1_6 ) );
  DFF_X1 u1_uk_K_r1_reg_7 (.CK( clk ) , .D( u1_uk_K_r0_7 ) , .Q( u1_uk_K_r1_7 ) );
  DFF_X1 u1_uk_K_r1_reg_8 (.CK( clk ) , .D( u1_uk_K_r0_8 ) , .Q( u1_uk_K_r1_8 ) , .QN( u1_uk_n1313 ) );
  DFF_X1 u1_uk_K_r1_reg_9 (.CK( clk ) , .D( u1_uk_K_r0_9 ) , .Q( u1_uk_K_r1_9 ) , .QN( u1_uk_n1314 ) );
  DFF_X1 u1_uk_K_r2_reg_0 (.CK( clk ) , .D( u1_uk_K_r1_0 ) , .Q( u1_uk_K_r2_0 ) , .QN( u1_uk_n1349 ) );
  DFF_X1 u1_uk_K_r2_reg_1 (.CK( clk ) , .D( u1_uk_K_r1_1 ) , .Q( u1_uk_K_r2_1 ) , .QN( u1_uk_n1350 ) );
  DFF_X1 u1_uk_K_r2_reg_10 (.CK( clk ) , .D( u1_uk_K_r1_10 ) , .Q( u1_uk_K_r2_10 ) , .QN( u1_uk_n1357 ) );
  DFF_X1 u1_uk_K_r2_reg_11 (.CK( clk ) , .D( u1_uk_K_r1_11 ) , .Q( u1_uk_K_r2_11 ) , .QN( u1_uk_n1358 ) );
  DFF_X1 u1_uk_K_r2_reg_12 (.CK( clk ) , .D( u1_uk_K_r1_12 ) , .Q( u1_uk_K_r2_12 ) , .QN( u1_uk_n1359 ) );
  DFF_X1 u1_uk_K_r2_reg_13 (.CK( clk ) , .D( u1_uk_K_r1_13 ) , .Q( u1_uk_K_r2_13 ) );
  DFF_X1 u1_uk_K_r2_reg_14 (.CK( clk ) , .D( u1_uk_K_r1_14 ) , .Q( u1_uk_K_r2_14 ) , .QN( u1_uk_n1360 ) );
  DFF_X1 u1_uk_K_r2_reg_15 (.CK( clk ) , .D( u1_uk_K_r1_15 ) , .Q( u1_uk_K_r2_15 ) , .QN( u1_uk_n1361 ) );
  DFF_X1 u1_uk_K_r2_reg_16 (.CK( clk ) , .D( u1_uk_K_r1_16 ) , .Q( u1_uk_K_r2_16 ) );
  DFF_X1 u1_uk_K_r2_reg_17 (.CK( clk ) , .D( u1_uk_K_r1_17 ) , .Q( u1_uk_K_r2_17 ) , .QN( u1_uk_n1363 ) );
  DFF_X1 u1_uk_K_r2_reg_18 (.CK( clk ) , .D( u1_uk_K_r1_18 ) , .Q( u1_uk_K_r2_18 ) );
  DFF_X1 u1_uk_K_r2_reg_19 (.CK( clk ) , .D( u1_uk_K_r1_19 ) , .Q( u1_uk_K_r2_19 ) , .QN( u1_uk_n1365 ) );
  DFF_X1 u1_uk_K_r2_reg_2 (.CK( clk ) , .D( u1_uk_K_r1_2 ) , .Q( u1_uk_K_r2_2 ) , .QN( u1_uk_n1351 ) );
  DFF_X1 u1_uk_K_r2_reg_20 (.CK( clk ) , .D( u1_uk_K_r1_20 ) , .Q( u1_uk_K_r2_20 ) );
  DFF_X1 u1_uk_K_r2_reg_21 (.CK( clk ) , .D( u1_uk_K_r1_21 ) , .Q( u1_uk_K_r2_21 ) );
  DFF_X1 u1_uk_K_r2_reg_22 (.CK( clk ) , .D( u1_uk_K_r1_22 ) , .Q( u1_uk_K_r2_22 ) , .QN( u1_uk_n1366 ) );
  DFF_X1 u1_uk_K_r2_reg_23 (.CK( clk ) , .D( u1_uk_K_r1_23 ) , .Q( u1_uk_K_r2_23 ) , .QN( u1_uk_n1367 ) );
  DFF_X1 u1_uk_K_r2_reg_24 (.CK( clk ) , .D( u1_uk_K_r1_24 ) , .Q( u1_uk_K_r2_24 ) );
  DFF_X1 u1_uk_K_r2_reg_25 (.CK( clk ) , .D( u1_uk_K_r1_25 ) , .Q( u1_uk_K_r2_25 ) );
  DFF_X1 u1_uk_K_r2_reg_26 (.CK( clk ) , .D( u1_uk_K_r1_26 ) , .Q( u1_uk_K_r2_26 ) );
  DFF_X1 u1_uk_K_r2_reg_27 (.CK( clk ) , .D( u1_uk_K_r1_27 ) , .Q( u1_uk_K_r2_27 ) );
  DFF_X1 u1_uk_K_r2_reg_28 (.CK( clk ) , .D( u1_uk_K_r1_28 ) , .Q( u1_uk_K_r2_28 ) );
  DFF_X1 u1_uk_K_r2_reg_29 (.CK( clk ) , .D( u1_uk_K_r1_29 ) , .Q( u1_uk_K_r2_29 ) );
  DFF_X1 u1_uk_K_r2_reg_3 (.CK( clk ) , .D( u1_uk_K_r1_3 ) , .Q( u1_uk_K_r2_3 ) , .QN( u1_uk_n1352 ) );
  DFF_X1 u1_uk_K_r2_reg_30 (.CK( clk ) , .D( u1_uk_K_r1_30 ) , .Q( u1_uk_K_r2_30 ) );
  DFF_X1 u1_uk_K_r2_reg_31 (.CK( clk ) , .D( u1_uk_K_r1_31 ) , .Q( u1_uk_K_r2_31 ) );
  DFF_X1 u1_uk_K_r2_reg_32 (.CK( clk ) , .D( u1_uk_K_r1_32 ) , .Q( u1_uk_K_r2_32 ) , .QN( u1_uk_n1369 ) );
  DFF_X1 u1_uk_K_r2_reg_33 (.CK( clk ) , .D( u1_uk_K_r1_33 ) , .Q( u1_uk_K_r2_33 ) );
  DFF_X1 u1_uk_K_r2_reg_34 (.CK( clk ) , .D( u1_uk_K_r1_34 ) , .Q( u1_uk_K_r2_34 ) , .QN( u1_uk_n1371 ) );
  DFF_X1 u1_uk_K_r2_reg_35 (.CK( clk ) , .D( u1_uk_K_r1_35 ) , .Q( u1_uk_K_r2_35 ) , .QN( u1_uk_n1372 ) );
  DFF_X1 u1_uk_K_r2_reg_36 (.CK( clk ) , .D( u1_uk_K_r1_36 ) , .Q( u1_uk_K_r2_36 ) , .QN( u1_uk_n1374 ) );
  DFF_X1 u1_uk_K_r2_reg_37 (.CK( clk ) , .D( u1_uk_K_r1_37 ) , .Q( u1_uk_K_r2_37 ) , .QN( u1_uk_n1375 ) );
  DFF_X1 u1_uk_K_r2_reg_38 (.CK( clk ) , .D( u1_uk_K_r1_38 ) , .Q( u1_uk_K_r2_38 ) , .QN( u1_uk_n1376 ) );
  DFF_X1 u1_uk_K_r2_reg_39 (.CK( clk ) , .D( u1_uk_K_r1_39 ) , .Q( u1_uk_K_r2_39 ) , .QN( u1_uk_n1377 ) );
  DFF_X1 u1_uk_K_r2_reg_4 (.CK( clk ) , .D( u1_uk_K_r1_4 ) , .Q( u1_uk_K_r2_4 ) );
  DFF_X1 u1_uk_K_r2_reg_40 (.CK( clk ) , .D( u1_uk_K_r1_40 ) , .Q( u1_uk_K_r2_40 ) , .QN( u1_uk_n1378 ) );
  DFF_X1 u1_uk_K_r2_reg_41 (.CK( clk ) , .D( u1_uk_K_r1_41 ) , .Q( u1_uk_K_r2_41 ) );
  DFF_X1 u1_uk_K_r2_reg_42 (.CK( clk ) , .D( u1_uk_K_r1_42 ) , .Q( u1_uk_K_r2_42 ) , .QN( u1_uk_n1380 ) );
  DFF_X1 u1_uk_K_r2_reg_43 (.CK( clk ) , .D( u1_uk_K_r1_43 ) , .Q( u1_uk_K_r2_43 ) , .QN( u1_uk_n1381 ) );
  DFF_X1 u1_uk_K_r2_reg_44 (.CK( clk ) , .D( u1_uk_K_r1_44 ) , .Q( u1_uk_K_r2_44 ) , .QN( u1_uk_n1382 ) );
  DFF_X1 u1_uk_K_r2_reg_45 (.CK( clk ) , .D( u1_uk_K_r1_45 ) , .Q( u1_uk_K_r2_45 ) , .QN( u1_uk_n1383 ) );
  DFF_X1 u1_uk_K_r2_reg_46 (.CK( clk ) , .D( u1_uk_K_r1_46 ) , .Q( u1_uk_K_r2_46 ) );
  DFF_X1 u1_uk_K_r2_reg_47 (.CK( clk ) , .D( u1_uk_K_r1_47 ) , .Q( u1_uk_K_r2_47 ) );
  DFF_X1 u1_uk_K_r2_reg_48 (.CK( clk ) , .D( u1_uk_K_r1_48 ) , .Q( u1_uk_K_r2_48 ) , .QN( u1_uk_n1386 ) );
  DFF_X1 u1_uk_K_r2_reg_49 (.CK( clk ) , .D( u1_uk_K_r1_49 ) , .Q( u1_uk_K_r2_49 ) );
  DFF_X1 u1_uk_K_r2_reg_5 (.CK( clk ) , .D( u1_uk_K_r1_5 ) , .Q( u1_uk_K_r2_5 ) , .QN( u1_uk_n1353 ) );
  DFF_X1 u1_uk_K_r2_reg_50 (.CK( clk ) , .D( u1_uk_K_r1_50 ) , .Q( u1_uk_K_r2_50 ) );
  DFF_X1 u1_uk_K_r2_reg_51 (.CK( clk ) , .D( u1_uk_K_r1_51 ) , .Q( u1_uk_K_r2_51 ) , .QN( u1_uk_n1389 ) );
  DFF_X1 u1_uk_K_r2_reg_52 (.CK( clk ) , .D( u1_uk_K_r1_52 ) , .Q( u1_uk_K_r2_52 ) , .QN( u1_uk_n1390 ) );
  DFF_X1 u1_uk_K_r2_reg_53 (.CK( clk ) , .D( u1_uk_K_r1_53 ) , .Q( u1_uk_K_r2_53 ) );
  DFF_X1 u1_uk_K_r2_reg_54 (.CK( clk ) , .D( u1_uk_K_r1_54 ) , .Q( u1_uk_K_r2_54 ) , .QN( u1_uk_n1391 ) );
  DFF_X1 u1_uk_K_r2_reg_55 (.CK( clk ) , .D( u1_uk_K_r1_55 ) , .Q( u1_uk_K_r2_55 ) , .QN( u1_uk_n1393 ) );
  DFF_X1 u1_uk_K_r2_reg_6 (.CK( clk ) , .D( u1_uk_K_r1_6 ) , .Q( u1_uk_K_r2_6 ) , .QN( u1_uk_n1354 ) );
  DFF_X1 u1_uk_K_r2_reg_7 (.CK( clk ) , .D( u1_uk_K_r1_7 ) , .Q( u1_uk_K_r2_7 ) );
  DFF_X1 u1_uk_K_r2_reg_8 (.CK( clk ) , .D( u1_uk_K_r1_8 ) , .Q( u1_uk_K_r2_8 ) , .QN( u1_uk_n1355 ) );
  DFF_X1 u1_uk_K_r2_reg_9 (.CK( clk ) , .D( u1_uk_K_r1_9 ) , .Q( u1_uk_K_r2_9 ) , .QN( u1_uk_n1356 ) );
  DFF_X1 u1_uk_K_r3_reg_0 (.CK( clk ) , .D( u1_uk_K_r2_0 ) , .Q( u1_uk_K_r3_0 ) , .QN( u1_uk_n1394 ) );
  DFF_X1 u1_uk_K_r3_reg_1 (.CK( clk ) , .D( u1_uk_K_r2_1 ) , .Q( u1_uk_K_r3_1 ) , .QN( u1_uk_n1395 ) );
  DFF_X1 u1_uk_K_r3_reg_10 (.CK( clk ) , .D( u1_uk_K_r2_10 ) , .Q( u1_uk_K_r3_10 ) );
  DFF_X1 u1_uk_K_r3_reg_11 (.CK( clk ) , .D( u1_uk_K_r2_11 ) , .Q( u1_uk_K_r3_11 ) );
  DFF_X1 u1_uk_K_r3_reg_12 (.CK( clk ) , .D( u1_uk_K_r2_12 ) , .Q( u1_uk_K_r3_12 ) , .QN( u1_uk_n1402 ) );
  DFF_X1 u1_uk_K_r3_reg_13 (.CK( clk ) , .D( u1_uk_K_r2_13 ) , .Q( u1_uk_K_r3_13 ) );
  DFF_X1 u1_uk_K_r3_reg_14 (.CK( clk ) , .D( u1_uk_K_r2_14 ) , .Q( u1_uk_K_r3_14 ) );
  DFF_X1 u1_uk_K_r3_reg_15 (.CK( clk ) , .D( u1_uk_K_r2_15 ) , .Q( u1_uk_K_r3_15 ) );
  DFF_X1 u1_uk_K_r3_reg_16 (.CK( clk ) , .D( u1_uk_K_r2_16 ) , .Q( u1_uk_K_r3_16 ) );
  DFF_X1 u1_uk_K_r3_reg_17 (.CK( clk ) , .D( u1_uk_K_r2_17 ) , .Q( u1_uk_K_r3_17 ) , .QN( u1_uk_n1403 ) );
  DFF_X1 u1_uk_K_r3_reg_18 (.CK( clk ) , .D( u1_uk_K_r2_18 ) , .Q( u1_uk_K_r3_18 ) , .QN( u1_uk_n1404 ) );
  DFF_X1 u1_uk_K_r3_reg_19 (.CK( clk ) , .D( u1_uk_K_r2_19 ) , .Q( u1_uk_K_r3_19 ) );
  DFF_X1 u1_uk_K_r3_reg_2 (.CK( clk ) , .D( u1_uk_K_r2_2 ) , .Q( u1_uk_K_r3_2 ) , .QN( u1_uk_n1396 ) );
  DFF_X1 u1_uk_K_r3_reg_20 (.CK( clk ) , .D( u1_uk_K_r2_20 ) , .Q( u1_uk_K_r3_20 ) , .QN( u1_uk_n1405 ) );
  DFF_X1 u1_uk_K_r3_reg_21 (.CK( clk ) , .D( u1_uk_K_r2_21 ) , .Q( u1_uk_K_r3_21 ) , .QN( u1_uk_n1406 ) );
  DFF_X1 u1_uk_K_r3_reg_22 (.CK( clk ) , .D( u1_uk_K_r2_22 ) , .Q( u1_uk_K_r3_22 ) , .QN( u1_uk_n1407 ) );
  DFF_X1 u1_uk_K_r3_reg_23 (.CK( clk ) , .D( u1_uk_K_r2_23 ) , .Q( u1_uk_K_r3_23 ) , .QN( u1_uk_n1408 ) );
  DFF_X1 u1_uk_K_r3_reg_24 (.CK( clk ) , .D( u1_uk_K_r2_24 ) , .Q( u1_uk_K_r3_24 ) );
  DFF_X1 u1_uk_K_r3_reg_25 (.CK( clk ) , .D( u1_uk_K_r2_25 ) , .Q( u1_uk_K_r3_25 ) , .QN( u1_uk_n1409 ) );
  DFF_X1 u1_uk_K_r3_reg_26 (.CK( clk ) , .D( u1_uk_K_r2_26 ) , .Q( u1_uk_K_r3_26 ) , .QN( u1_uk_n1410 ) );
  DFF_X1 u1_uk_K_r3_reg_27 (.CK( clk ) , .D( u1_uk_K_r2_27 ) , .Q( u1_uk_K_r3_27 ) , .QN( u1_uk_n1411 ) );
  DFF_X1 u1_uk_K_r3_reg_28 (.CK( clk ) , .D( u1_uk_K_r2_28 ) , .Q( u1_uk_K_r3_28 ) , .QN( u1_uk_n1412 ) );
  DFF_X1 u1_uk_K_r3_reg_29 (.CK( clk ) , .D( u1_uk_K_r2_29 ) , .Q( u1_uk_K_r3_29 ) );
  DFF_X1 u1_uk_K_r3_reg_3 (.CK( clk ) , .D( u1_uk_K_r2_3 ) , .Q( u1_uk_K_r3_3 ) , .QN( u1_uk_n1397 ) );
  DFF_X1 u1_uk_K_r3_reg_30 (.CK( clk ) , .D( u1_uk_K_r2_30 ) , .Q( u1_uk_K_r3_30 ) , .QN( u1_uk_n1413 ) );
  DFF_X1 u1_uk_K_r3_reg_31 (.CK( clk ) , .D( u1_uk_K_r2_31 ) , .Q( u1_uk_K_r3_31 ) , .QN( u1_uk_n1414 ) );
  DFF_X1 u1_uk_K_r3_reg_32 (.CK( clk ) , .D( u1_uk_K_r2_32 ) , .Q( u1_uk_K_r3_32 ) , .QN( u1_uk_n1415 ) );
  DFF_X1 u1_uk_K_r3_reg_33 (.CK( clk ) , .D( u1_uk_K_r2_33 ) , .Q( u1_uk_K_r3_33 ) , .QN( u1_uk_n1417 ) );
  DFF_X1 u1_uk_K_r3_reg_34 (.CK( clk ) , .D( u1_uk_K_r2_34 ) , .Q( u1_uk_K_r3_34 ) );
  DFF_X1 u1_uk_K_r3_reg_35 (.CK( clk ) , .D( u1_uk_K_r2_35 ) , .Q( u1_uk_K_r3_35 ) );
  DFF_X1 u1_uk_K_r3_reg_36 (.CK( clk ) , .D( u1_uk_K_r2_36 ) , .Q( u1_uk_K_r3_36 ) , .QN( u1_uk_n1418 ) );
  DFF_X1 u1_uk_K_r3_reg_37 (.CK( clk ) , .D( u1_uk_K_r2_37 ) , .Q( u1_uk_K_r3_37 ) , .QN( u1_uk_n1419 ) );
  DFF_X1 u1_uk_K_r3_reg_38 (.CK( clk ) , .D( u1_uk_K_r2_38 ) , .Q( u1_uk_K_r3_38 ) );
  DFF_X1 u1_uk_K_r3_reg_39 (.CK( clk ) , .D( u1_uk_K_r2_39 ) , .Q( u1_uk_K_r3_39 ) , .QN( u1_uk_n1422 ) );
  DFF_X1 u1_uk_K_r3_reg_4 (.CK( clk ) , .D( u1_uk_K_r2_4 ) , .Q( u1_uk_K_r3_4 ) );
  DFF_X1 u1_uk_K_r3_reg_40 (.CK( clk ) , .D( u1_uk_K_r2_40 ) , .Q( u1_uk_K_r3_40 ) , .QN( u1_uk_n1423 ) );
  DFF_X1 u1_uk_K_r3_reg_41 (.CK( clk ) , .D( u1_uk_K_r2_41 ) , .Q( u1_uk_K_r3_41 ) , .QN( u1_uk_n1424 ) );
  DFF_X1 u1_uk_K_r3_reg_42 (.CK( clk ) , .D( u1_uk_K_r2_42 ) , .Q( u1_uk_K_r3_42 ) , .QN( u1_uk_n1425 ) );
  DFF_X1 u1_uk_K_r3_reg_43 (.CK( clk ) , .D( u1_uk_K_r2_43 ) , .Q( u1_uk_K_r3_43 ) );
  DFF_X1 u1_uk_K_r3_reg_44 (.CK( clk ) , .D( u1_uk_K_r2_44 ) , .Q( u1_uk_K_r3_44 ) );
  DFF_X1 u1_uk_K_r3_reg_45 (.CK( clk ) , .D( u1_uk_K_r2_45 ) , .Q( u1_uk_K_r3_45 ) , .QN( u1_uk_n1426 ) );
  DFF_X1 u1_uk_K_r3_reg_46 (.CK( clk ) , .D( u1_uk_K_r2_46 ) , .Q( u1_uk_K_r3_46 ) , .QN( u1_uk_n1427 ) );
  DFF_X1 u1_uk_K_r3_reg_47 (.CK( clk ) , .D( u1_uk_K_r2_47 ) , .Q( u1_uk_K_r3_47 ) );
  DFF_X1 u1_uk_K_r3_reg_48 (.CK( clk ) , .D( u1_uk_K_r2_48 ) , .Q( u1_uk_K_r3_48 ) , .QN( u1_uk_n1429 ) );
  DFF_X1 u1_uk_K_r3_reg_49 (.CK( clk ) , .D( u1_uk_K_r2_49 ) , .Q( u1_uk_K_r3_49 ) , .QN( u1_uk_n1430 ) );
  DFF_X1 u1_uk_K_r3_reg_5 (.CK( clk ) , .D( u1_uk_K_r2_5 ) , .Q( u1_uk_K_r3_5 ) , .QN( u1_uk_n1398 ) );
  DFF_X1 u1_uk_K_r3_reg_50 (.CK( clk ) , .D( u1_uk_K_r2_50 ) , .Q( u1_uk_K_r3_50 ) , .QN( u1_uk_n1431 ) );
  DFF_X1 u1_uk_K_r3_reg_51 (.CK( clk ) , .D( u1_uk_K_r2_51 ) , .Q( u1_uk_K_r3_51 ) , .QN( u1_uk_n1433 ) );
  DFF_X1 u1_uk_K_r3_reg_52 (.CK( clk ) , .D( u1_uk_K_r2_52 ) , .Q( u1_uk_K_r3_52 ) );
  DFF_X1 u1_uk_K_r3_reg_53 (.CK( clk ) , .D( u1_uk_K_r2_53 ) , .Q( u1_uk_K_r3_53 ) , .QN( u1_uk_n1435 ) );
  DFF_X1 u1_uk_K_r3_reg_54 (.CK( clk ) , .D( u1_uk_K_r2_54 ) , .Q( u1_uk_K_r3_54 ) , .QN( u1_uk_n1436 ) );
  DFF_X1 u1_uk_K_r3_reg_55 (.CK( clk ) , .D( u1_uk_K_r2_55 ) , .Q( u1_uk_K_r3_55 ) , .QN( u1_uk_n1437 ) );
  DFF_X1 u1_uk_K_r3_reg_6 (.CK( clk ) , .D( u1_uk_K_r2_6 ) , .Q( u1_uk_K_r3_6 ) , .QN( u1_uk_n1399 ) );
  DFF_X1 u1_uk_K_r3_reg_7 (.CK( clk ) , .D( u1_uk_K_r2_7 ) , .Q( u1_uk_K_r3_7 ) , .QN( u1_uk_n1400 ) );
  DFF_X1 u1_uk_K_r3_reg_8 (.CK( clk ) , .D( u1_uk_K_r2_8 ) , .Q( u1_uk_K_r3_8 ) , .QN( u1_uk_n1401 ) );
  DFF_X1 u1_uk_K_r3_reg_9 (.CK( clk ) , .D( u1_uk_K_r2_9 ) , .Q( u1_uk_K_r3_9 ) );
  DFF_X1 u1_uk_K_r4_reg_0 (.CK( clk ) , .D( u1_uk_K_r3_0 ) , .Q( u1_uk_K_r4_0 ) );
  DFF_X1 u1_uk_K_r4_reg_1 (.CK( clk ) , .D( u1_uk_K_r3_1 ) , .Q( u1_uk_K_r4_1 ) , .QN( u1_uk_n1438 ) );
  DFF_X1 u1_uk_K_r4_reg_10 (.CK( clk ) , .D( u1_uk_K_r3_10 ) , .Q( u1_uk_K_r4_10 ) , .QN( u1_uk_n1444 ) );
  DFF_X1 u1_uk_K_r4_reg_11 (.CK( clk ) , .D( u1_uk_K_r3_11 ) , .Q( u1_uk_K_r4_11 ) );
  DFF_X1 u1_uk_K_r4_reg_12 (.CK( clk ) , .D( u1_uk_K_r3_12 ) , .Q( u1_uk_K_r4_12 ) , .QN( u1_uk_n1446 ) );
  DFF_X1 u1_uk_K_r4_reg_13 (.CK( clk ) , .D( u1_uk_K_r3_13 ) , .Q( u1_uk_K_r4_13 ) , .QN( u1_uk_n1447 ) );
  DFF_X1 u1_uk_K_r4_reg_14 (.CK( clk ) , .D( u1_uk_K_r3_14 ) , .Q( u1_uk_K_r4_14 ) , .QN( u1_uk_n1448 ) );
  DFF_X1 u1_uk_K_r4_reg_15 (.CK( clk ) , .D( u1_uk_K_r3_15 ) , .Q( u1_uk_K_r4_15 ) , .QN( u1_uk_n1449 ) );
  DFF_X1 u1_uk_K_r4_reg_16 (.CK( clk ) , .D( u1_uk_K_r3_16 ) , .Q( u1_uk_K_r4_16 ) , .QN( u1_uk_n1450 ) );
  DFF_X1 u1_uk_K_r4_reg_17 (.CK( clk ) , .D( u1_uk_K_r3_17 ) , .Q( u1_uk_K_r4_17 ) );
  DFF_X1 u1_uk_K_r4_reg_18 (.CK( clk ) , .D( u1_uk_K_r3_18 ) , .Q( u1_uk_K_r4_18 ) );
  DFF_X1 u1_uk_K_r4_reg_19 (.CK( clk ) , .D( u1_uk_K_r3_19 ) , .Q( u1_uk_K_r4_19 ) , .QN( u1_uk_n1452 ) );
  DFF_X1 u1_uk_K_r4_reg_2 (.CK( clk ) , .D( u1_uk_K_r3_2 ) , .Q( u1_uk_K_r4_2 ) );
  DFF_X1 u1_uk_K_r4_reg_20 (.CK( clk ) , .D( u1_uk_K_r3_20 ) , .Q( u1_uk_K_r4_20 ) , .QN( u1_uk_n1453 ) );
  DFF_X1 u1_uk_K_r4_reg_21 (.CK( clk ) , .D( u1_uk_K_r3_21 ) , .Q( u1_uk_K_r4_21 ) , .QN( u1_uk_n1454 ) );
  DFF_X1 u1_uk_K_r4_reg_22 (.CK( clk ) , .D( u1_uk_K_r3_22 ) , .Q( u1_uk_K_r4_22 ) , .QN( u1_uk_n1455 ) );
  DFF_X1 u1_uk_K_r4_reg_23 (.CK( clk ) , .D( u1_uk_K_r3_23 ) , .Q( u1_uk_K_r4_23 ) );
  DFF_X1 u1_uk_K_r4_reg_24 (.CK( clk ) , .D( u1_uk_K_r3_24 ) , .Q( u1_uk_K_r4_24 ) );
  DFF_X1 u1_uk_K_r4_reg_25 (.CK( clk ) , .D( u1_uk_K_r3_25 ) , .Q( u1_uk_K_r4_25 ) , .QN( u1_uk_n1456 ) );
  DFF_X1 u1_uk_K_r4_reg_26 (.CK( clk ) , .D( u1_uk_K_r3_26 ) , .Q( u1_uk_K_r4_26 ) , .QN( u1_uk_n1457 ) );
  DFF_X1 u1_uk_K_r4_reg_27 (.CK( clk ) , .D( u1_uk_K_r3_27 ) , .Q( u1_uk_K_r4_27 ) );
  DFF_X1 u1_uk_K_r4_reg_28 (.CK( clk ) , .D( u1_uk_K_r3_28 ) , .Q( u1_uk_K_r4_28 ) , .QN( u1_uk_n1458 ) );
  DFF_X1 u1_uk_K_r4_reg_29 (.CK( clk ) , .D( u1_uk_K_r3_29 ) , .Q( u1_uk_K_r4_29 ) , .QN( u1_uk_n1459 ) );
  DFF_X1 u1_uk_K_r4_reg_3 (.CK( clk ) , .D( u1_uk_K_r3_3 ) , .Q( u1_uk_K_r4_3 ) );
  DFF_X1 u1_uk_K_r4_reg_30 (.CK( clk ) , .D( u1_uk_K_r3_30 ) , .Q( u1_uk_K_r4_30 ) , .QN( u1_uk_n1460 ) );
  DFF_X1 u1_uk_K_r4_reg_31 (.CK( clk ) , .D( u1_uk_K_r3_31 ) , .Q( u1_uk_K_r4_31 ) );
  DFF_X1 u1_uk_K_r4_reg_32 (.CK( clk ) , .D( u1_uk_K_r3_32 ) , .Q( u1_uk_K_r4_32 ) , .QN( u1_uk_n1461 ) );
  DFF_X1 u1_uk_K_r4_reg_33 (.CK( clk ) , .D( u1_uk_K_r3_33 ) , .Q( u1_uk_K_r4_33 ) );
  DFF_X1 u1_uk_K_r4_reg_34 (.CK( clk ) , .D( u1_uk_K_r3_34 ) , .Q( u1_uk_K_r4_34 ) , .QN( u1_uk_n1462 ) );
  DFF_X1 u1_uk_K_r4_reg_35 (.CK( clk ) , .D( u1_uk_K_r3_35 ) , .Q( u1_uk_K_r4_35 ) );
  DFF_X1 u1_uk_K_r4_reg_36 (.CK( clk ) , .D( u1_uk_K_r3_36 ) , .Q( u1_uk_K_r4_36 ) , .QN( u1_uk_n1463 ) );
  DFF_X1 u1_uk_K_r4_reg_37 (.CK( clk ) , .D( u1_uk_K_r3_37 ) , .Q( u1_uk_K_r4_37 ) , .QN( u1_uk_n1464 ) );
  DFF_X1 u1_uk_K_r4_reg_38 (.CK( clk ) , .D( u1_uk_K_r3_38 ) , .Q( u1_uk_K_r4_38 ) );
  DFF_X1 u1_uk_K_r4_reg_39 (.CK( clk ) , .D( u1_uk_K_r3_39 ) , .Q( u1_uk_K_r4_39 ) , .QN( u1_uk_n1465 ) );
  DFF_X1 u1_uk_K_r4_reg_4 (.CK( clk ) , .D( u1_uk_K_r3_4 ) , .Q( u1_uk_K_r4_4 ) , .QN( u1_uk_n1439 ) );
  DFF_X1 u1_uk_K_r4_reg_40 (.CK( clk ) , .D( u1_uk_K_r3_40 ) , .Q( u1_uk_K_r4_40 ) , .QN( u1_uk_n1466 ) );
  DFF_X1 u1_uk_K_r4_reg_41 (.CK( clk ) , .D( u1_uk_K_r3_41 ) , .Q( u1_uk_K_r4_41 ) );
  DFF_X1 u1_uk_K_r4_reg_42 (.CK( clk ) , .D( u1_uk_K_r3_42 ) , .Q( u1_uk_K_r4_42 ) , .QN( u1_uk_n1468 ) );
  DFF_X1 u1_uk_K_r4_reg_43 (.CK( clk ) , .D( u1_uk_K_r3_43 ) , .Q( u1_uk_K_r4_43 ) , .QN( u1_uk_n1469 ) );
  DFF_X1 u1_uk_K_r4_reg_44 (.CK( clk ) , .D( u1_uk_K_r3_44 ) , .Q( u1_uk_K_r4_44 ) , .QN( u1_uk_n1470 ) );
  DFF_X1 u1_uk_K_r4_reg_45 (.CK( clk ) , .D( u1_uk_K_r3_45 ) , .Q( u1_uk_K_r4_45 ) , .QN( u1_uk_n1471 ) );
  DFF_X1 u1_uk_K_r4_reg_46 (.CK( clk ) , .D( u1_uk_K_r3_46 ) , .Q( u1_uk_K_r4_46 ) , .QN( u1_uk_n1472 ) );
  DFF_X1 u1_uk_K_r4_reg_47 (.CK( clk ) , .D( u1_uk_K_r3_47 ) , .Q( u1_uk_K_r4_47 ) , .QN( u1_uk_n1474 ) );
  DFF_X1 u1_uk_K_r4_reg_48 (.CK( clk ) , .D( u1_uk_K_r3_48 ) , .Q( u1_uk_K_r4_48 ) );
  DFF_X1 u1_uk_K_r4_reg_49 (.CK( clk ) , .D( u1_uk_K_r3_49 ) , .Q( u1_uk_K_r4_49 ) );
  DFF_X1 u1_uk_K_r4_reg_5 (.CK( clk ) , .D( u1_uk_K_r3_5 ) , .Q( u1_uk_K_r4_5 ) );
  DFF_X1 u1_uk_K_r4_reg_50 (.CK( clk ) , .D( u1_uk_K_r3_50 ) , .Q( u1_uk_K_r4_50 ) , .QN( u1_uk_n1475 ) );
  DFF_X1 u1_uk_K_r4_reg_51 (.CK( clk ) , .D( u1_uk_K_r3_51 ) , .Q( u1_uk_K_r4_51 ) , .QN( u1_uk_n1476 ) );
  DFF_X1 u1_uk_K_r4_reg_52 (.CK( clk ) , .D( u1_uk_K_r3_52 ) , .Q( u1_uk_K_r4_52 ) , .QN( u1_uk_n1477 ) );
  DFF_X1 u1_uk_K_r4_reg_53 (.CK( clk ) , .D( u1_uk_K_r3_53 ) , .Q( u1_uk_K_r4_53 ) , .QN( u1_uk_n1478 ) );
  DFF_X1 u1_uk_K_r4_reg_54 (.CK( clk ) , .D( u1_uk_K_r3_54 ) , .Q( u1_uk_K_r4_54 ) );
  DFF_X1 u1_uk_K_r4_reg_55 (.CK( clk ) , .D( u1_uk_K_r3_55 ) , .Q( u1_uk_K_r4_55 ) );
  DFF_X1 u1_uk_K_r4_reg_6 (.CK( clk ) , .D( u1_uk_K_r3_6 ) , .Q( u1_uk_K_r4_6 ) , .QN( u1_uk_n1440 ) );
  DFF_X1 u1_uk_K_r4_reg_7 (.CK( clk ) , .D( u1_uk_K_r3_7 ) , .Q( u1_uk_K_r4_7 ) , .QN( u1_uk_n1441 ) );
  DFF_X1 u1_uk_K_r4_reg_8 (.CK( clk ) , .D( u1_uk_K_r3_8 ) , .Q( u1_uk_K_r4_8 ) , .QN( u1_uk_n1442 ) );
  DFF_X1 u1_uk_K_r4_reg_9 (.CK( clk ) , .D( u1_uk_K_r3_9 ) , .Q( u1_uk_K_r4_9 ) , .QN( u1_uk_n1443 ) );
  DFF_X1 u1_uk_K_r5_reg_0 (.CK( clk ) , .D( u1_uk_K_r4_0 ) , .Q( u1_uk_K_r5_0 ) );
  DFF_X1 u1_uk_K_r5_reg_1 (.CK( clk ) , .D( u1_uk_K_r4_1 ) , .Q( u1_uk_K_r5_1 ) );
  DFF_X1 u1_uk_K_r5_reg_10 (.CK( clk ) , .D( u1_uk_K_r4_10 ) , .Q( u1_uk_K_r5_10 ) );
  DFF_X1 u1_uk_K_r5_reg_11 (.CK( clk ) , .D( u1_uk_K_r4_11 ) , .Q( u1_uk_K_r5_11 ) , .QN( u1_uk_n1487 ) );
  DFF_X1 u1_uk_K_r5_reg_12 (.CK( clk ) , .D( u1_uk_K_r4_12 ) , .Q( u1_uk_K_r5_12 ) , .QN( u1_uk_n1488 ) );
  DFF_X1 u1_uk_K_r5_reg_13 (.CK( clk ) , .D( u1_uk_K_r4_13 ) , .Q( u1_uk_K_r5_13 ) );
  DFF_X1 u1_uk_K_r5_reg_14 (.CK( clk ) , .D( u1_uk_K_r4_14 ) , .Q( u1_uk_K_r5_14 ) , .QN( u1_uk_n1489 ) );
  DFF_X1 u1_uk_K_r5_reg_15 (.CK( clk ) , .D( u1_uk_K_r4_15 ) , .Q( u1_uk_K_r5_15 ) , .QN( u1_uk_n1490 ) );
  DFF_X1 u1_uk_K_r5_reg_16 (.CK( clk ) , .D( u1_uk_K_r4_16 ) , .Q( u1_uk_K_r5_16 ) );
  DFF_X1 u1_uk_K_r5_reg_17 (.CK( clk ) , .D( u1_uk_K_r4_17 ) , .Q( u1_uk_K_r5_17 ) , .QN( u1_uk_n1491 ) );
  DFF_X1 u1_uk_K_r5_reg_18 (.CK( clk ) , .D( u1_uk_K_r4_18 ) , .Q( u1_uk_K_r5_18 ) );
  DFF_X1 u1_uk_K_r5_reg_19 (.CK( clk ) , .D( u1_uk_K_r4_19 ) , .Q( u1_uk_K_r5_19 ) );
  DFF_X1 u1_uk_K_r5_reg_2 (.CK( clk ) , .D( u1_uk_K_r4_2 ) , .Q( u1_uk_K_r5_2 ) , .QN( u1_uk_n1482 ) );
  DFF_X1 u1_uk_K_r5_reg_20 (.CK( clk ) , .D( u1_uk_K_r4_20 ) , .Q( u1_uk_K_r5_20 ) , .QN( u1_uk_n1492 ) );
  DFF_X1 u1_uk_K_r5_reg_21 (.CK( clk ) , .D( u1_uk_K_r4_21 ) , .Q( u1_uk_K_r5_21 ) );
  DFF_X1 u1_uk_K_r5_reg_22 (.CK( clk ) , .D( u1_uk_K_r4_22 ) , .Q( u1_uk_K_r5_22 ) , .QN( u1_uk_n1494 ) );
  DFF_X1 u1_uk_K_r5_reg_23 (.CK( clk ) , .D( u1_uk_K_r4_23 ) , .Q( u1_uk_K_r5_23 ) );
  DFF_X1 u1_uk_K_r5_reg_24 (.CK( clk ) , .D( u1_uk_K_r4_24 ) , .Q( u1_uk_K_r5_24 ) , .QN( u1_uk_n1495 ) );
  DFF_X1 u1_uk_K_r5_reg_25 (.CK( clk ) , .D( u1_uk_K_r4_25 ) , .Q( u1_uk_K_r5_25 ) , .QN( u1_uk_n1496 ) );
  DFF_X1 u1_uk_K_r5_reg_26 (.CK( clk ) , .D( u1_uk_K_r4_26 ) , .Q( u1_uk_K_r5_26 ) );
  DFF_X1 u1_uk_K_r5_reg_27 (.CK( clk ) , .D( u1_uk_K_r4_27 ) , .Q( u1_uk_K_r5_27 ) , .QN( u1_uk_n1498 ) );
  DFF_X1 u1_uk_K_r5_reg_28 (.CK( clk ) , .D( u1_uk_K_r4_28 ) , .Q( u1_uk_K_r5_28 ) , .QN( u1_uk_n1499 ) );
  DFF_X1 u1_uk_K_r5_reg_29 (.CK( clk ) , .D( u1_uk_K_r4_29 ) , .Q( u1_uk_K_r5_29 ) , .QN( u1_uk_n1500 ) );
  DFF_X1 u1_uk_K_r5_reg_3 (.CK( clk ) , .D( u1_uk_K_r4_3 ) , .Q( u1_uk_K_r5_3 ) , .QN( u1_uk_n1483 ) );
  DFF_X1 u1_uk_K_r5_reg_30 (.CK( clk ) , .D( u1_uk_K_r4_30 ) , .Q( u1_uk_K_r5_30 ) , .QN( u1_uk_n1501 ) );
  DFF_X1 u1_uk_K_r5_reg_31 (.CK( clk ) , .D( u1_uk_K_r4_31 ) , .Q( u1_uk_K_r5_31 ) );
  DFF_X1 u1_uk_K_r5_reg_32 (.CK( clk ) , .D( u1_uk_K_r4_32 ) , .Q( u1_uk_K_r5_32 ) );
  DFF_X1 u1_uk_K_r5_reg_33 (.CK( clk ) , .D( u1_uk_K_r4_33 ) , .Q( u1_uk_K_r5_33 ) , .QN( u1_uk_n1504 ) );
  DFF_X1 u1_uk_K_r5_reg_34 (.CK( clk ) , .D( u1_uk_K_r4_34 ) , .Q( u1_uk_K_r5_34 ) , .QN( u1_uk_n1505 ) );
  DFF_X1 u1_uk_K_r5_reg_35 (.CK( clk ) , .D( u1_uk_K_r4_35 ) , .Q( u1_uk_K_r5_35 ) , .QN( u1_uk_n1507 ) );
  DFF_X1 u1_uk_K_r5_reg_36 (.CK( clk ) , .D( u1_uk_K_r4_36 ) , .Q( u1_uk_K_r5_36 ) , .QN( u1_uk_n1508 ) );
  DFF_X1 u1_uk_K_r5_reg_37 (.CK( clk ) , .D( u1_uk_K_r4_37 ) , .Q( u1_uk_K_r5_37 ) );
  DFF_X1 u1_uk_K_r5_reg_38 (.CK( clk ) , .D( u1_uk_K_r4_38 ) , .Q( u1_uk_K_r5_38 ) , .QN( u1_uk_n1510 ) );
  DFF_X1 u1_uk_K_r5_reg_39 (.CK( clk ) , .D( u1_uk_K_r4_39 ) , .Q( u1_uk_K_r5_39 ) );
  DFF_X1 u1_uk_K_r5_reg_4 (.CK( clk ) , .D( u1_uk_K_r4_4 ) , .Q( u1_uk_K_r5_4 ) );
  DFF_X1 u1_uk_K_r5_reg_40 (.CK( clk ) , .D( u1_uk_K_r4_40 ) , .Q( u1_uk_K_r5_40 ) );
  DFF_X1 u1_uk_K_r5_reg_41 (.CK( clk ) , .D( u1_uk_K_r4_41 ) , .Q( u1_uk_K_r5_41 ) );
  DFF_X1 u1_uk_K_r5_reg_42 (.CK( clk ) , .D( u1_uk_K_r4_42 ) , .Q( u1_uk_K_r5_42 ) , .QN( u1_uk_n1514 ) );
  DFF_X1 u1_uk_K_r5_reg_43 (.CK( clk ) , .D( u1_uk_K_r4_43 ) , .Q( u1_uk_K_r5_43 ) );
  DFF_X1 u1_uk_K_r5_reg_44 (.CK( clk ) , .D( u1_uk_K_r4_44 ) , .Q( u1_uk_K_r5_44 ) , .QN( u1_uk_n1516 ) );
  DFF_X1 u1_uk_K_r5_reg_45 (.CK( clk ) , .D( u1_uk_K_r4_45 ) , .Q( u1_uk_K_r5_45 ) );
  DFF_X1 u1_uk_K_r5_reg_46 (.CK( clk ) , .D( u1_uk_K_r4_46 ) , .Q( u1_uk_K_r5_46 ) , .QN( u1_uk_n1517 ) );
  DFF_X1 u1_uk_K_r5_reg_47 (.CK( clk ) , .D( u1_uk_K_r4_47 ) , .Q( u1_uk_K_r5_47 ) , .QN( u1_uk_n1518 ) );
  DFF_X1 u1_uk_K_r5_reg_48 (.CK( clk ) , .D( u1_uk_K_r4_48 ) , .Q( u1_uk_K_r5_48 ) );
  DFF_X1 u1_uk_K_r5_reg_49 (.CK( clk ) , .D( u1_uk_K_r4_49 ) , .Q( u1_uk_K_r5_49 ) , .QN( u1_uk_n1520 ) );
  DFF_X1 u1_uk_K_r5_reg_5 (.CK( clk ) , .D( u1_uk_K_r4_5 ) , .Q( u1_uk_K_r5_5 ) );
  DFF_X1 u1_uk_K_r5_reg_50 (.CK( clk ) , .D( u1_uk_K_r4_50 ) , .Q( u1_uk_K_r5_50 ) , .QN( u1_uk_n1521 ) );
  DFF_X1 u1_uk_K_r5_reg_51 (.CK( clk ) , .D( u1_uk_K_r4_51 ) , .Q( u1_uk_K_r5_51 ) );
  DFF_X1 u1_uk_K_r5_reg_52 (.CK( clk ) , .D( u1_uk_K_r4_52 ) , .Q( u1_uk_K_r5_52 ) , .QN( u1_uk_n1523 ) );
  DFF_X1 u1_uk_K_r5_reg_53 (.CK( clk ) , .D( u1_uk_K_r4_53 ) , .Q( u1_uk_K_r5_53 ) , .QN( u1_uk_n1524 ) );
  DFF_X1 u1_uk_K_r5_reg_54 (.CK( clk ) , .D( u1_uk_K_r4_54 ) , .Q( u1_uk_K_r5_54 ) , .QN( u1_uk_n1526 ) );
  DFF_X1 u1_uk_K_r5_reg_55 (.CK( clk ) , .D( u1_uk_K_r4_55 ) , .Q( u1_uk_K_r5_55 ) , .QN( u1_uk_n1527 ) );
  DFF_X1 u1_uk_K_r5_reg_6 (.CK( clk ) , .D( u1_uk_K_r4_6 ) , .Q( u1_uk_K_r5_6 ) , .QN( u1_uk_n1484 ) );
  DFF_X1 u1_uk_K_r5_reg_7 (.CK( clk ) , .D( u1_uk_K_r4_7 ) , .Q( u1_uk_K_r5_7 ) , .QN( u1_uk_n1485 ) );
  DFF_X1 u1_uk_K_r5_reg_8 (.CK( clk ) , .D( u1_uk_K_r4_8 ) , .Q( u1_uk_K_r5_8 ) );
  DFF_X1 u1_uk_K_r5_reg_9 (.CK( clk ) , .D( u1_uk_K_r4_9 ) , .Q( u1_uk_K_r5_9 ) , .QN( u1_uk_n1486 ) );
  DFF_X1 u1_uk_K_r6_reg_0 (.CK( clk ) , .D( u1_uk_K_r5_0 ) , .Q( u1_uk_K_r6_0 ) );
  DFF_X1 u1_uk_K_r6_reg_1 (.CK( clk ) , .D( u1_uk_K_r5_1 ) , .Q( u1_uk_K_r6_1 ) , .QN( u1_uk_n1528 ) );
  DFF_X1 u1_uk_K_r6_reg_10 (.CK( clk ) , .D( u1_uk_K_r5_10 ) , .Q( u1_uk_K_r6_10 ) );
  DFF_X1 u1_uk_K_r6_reg_11 (.CK( clk ) , .D( u1_uk_K_r5_11 ) , .Q( u1_uk_K_r6_11 ) , .QN( u1_uk_n1536 ) );
  DFF_X1 u1_uk_K_r6_reg_12 (.CK( clk ) , .D( u1_uk_K_r5_12 ) , .Q( u1_uk_K_r6_12 ) , .QN( u1_uk_n1537 ) );
  DFF_X1 u1_uk_K_r6_reg_13 (.CK( clk ) , .D( u1_uk_K_r5_13 ) , .Q( u1_uk_K_r6_13 ) , .QN( u1_uk_n1538 ) );
  DFF_X1 u1_uk_K_r6_reg_14 (.CK( clk ) , .D( u1_uk_K_r5_14 ) , .Q( u1_uk_K_r6_14 ) );
  DFF_X1 u1_uk_K_r6_reg_15 (.CK( clk ) , .D( u1_uk_K_r5_15 ) , .Q( u1_uk_K_r6_15 ) , .QN( u1_uk_n1540 ) );
  DFF_X1 u1_uk_K_r6_reg_16 (.CK( clk ) , .D( u1_uk_K_r5_16 ) , .Q( u1_uk_K_r6_16 ) , .QN( u1_uk_n1541 ) );
  DFF_X1 u1_uk_K_r6_reg_17 (.CK( clk ) , .D( u1_uk_K_r5_17 ) , .Q( u1_uk_K_r6_17 ) , .QN( u1_uk_n1543 ) );
  DFF_X1 u1_uk_K_r6_reg_18 (.CK( clk ) , .D( u1_uk_K_r5_18 ) , .Q( u1_uk_K_r6_18 ) , .QN( u1_uk_n1544 ) );
  DFF_X1 u1_uk_K_r6_reg_19 (.CK( clk ) , .D( u1_uk_K_r5_19 ) , .Q( u1_uk_K_r6_19 ) );
  DFF_X1 u1_uk_K_r6_reg_2 (.CK( clk ) , .D( u1_uk_K_r5_2 ) , .Q( u1_uk_K_r6_2 ) , .QN( u1_uk_n1529 ) );
  DFF_X1 u1_uk_K_r6_reg_20 (.CK( clk ) , .D( u1_uk_K_r5_20 ) , .Q( u1_uk_K_r6_20 ) , .QN( u1_uk_n1545 ) );
  DFF_X1 u1_uk_K_r6_reg_21 (.CK( clk ) , .D( u1_uk_K_r5_21 ) , .Q( u1_uk_K_r6_21 ) );
  DFF_X1 u1_uk_K_r6_reg_22 (.CK( clk ) , .D( u1_uk_K_r5_22 ) , .Q( u1_uk_K_r6_22 ) );
  DFF_X1 u1_uk_K_r6_reg_23 (.CK( clk ) , .D( u1_uk_K_r5_23 ) , .Q( u1_uk_K_r6_23 ) , .QN( u1_uk_n1547 ) );
  DFF_X1 u1_uk_K_r6_reg_24 (.CK( clk ) , .D( u1_uk_K_r5_24 ) , .Q( u1_uk_K_r6_24 ) , .QN( u1_uk_n1548 ) );
  DFF_X1 u1_uk_K_r6_reg_25 (.CK( clk ) , .D( u1_uk_K_r5_25 ) , .Q( u1_uk_K_r6_25 ) , .QN( u1_uk_n1549 ) );
  DFF_X1 u1_uk_K_r6_reg_26 (.CK( clk ) , .D( u1_uk_K_r5_26 ) , .Q( u1_uk_K_r6_26 ) );
  DFF_X1 u1_uk_K_r6_reg_27 (.CK( clk ) , .D( u1_uk_K_r5_27 ) , .Q( u1_uk_K_r6_27 ) );
  DFF_X1 u1_uk_K_r6_reg_28 (.CK( clk ) , .D( u1_uk_K_r5_28 ) , .Q( u1_uk_K_r6_28 ) );
  DFF_X1 u1_uk_K_r6_reg_29 (.CK( clk ) , .D( u1_uk_K_r5_29 ) , .Q( u1_uk_K_r6_29 ) );
  DFF_X1 u1_uk_K_r6_reg_3 (.CK( clk ) , .D( u1_uk_K_r5_3 ) , .Q( u1_uk_K_r6_3 ) );
  DFF_X1 u1_uk_K_r6_reg_30 (.CK( clk ) , .D( u1_uk_K_r5_30 ) , .Q( u1_uk_K_r6_30 ) );
  DFF_X1 u1_uk_K_r6_reg_31 (.CK( clk ) , .D( u1_uk_K_r5_31 ) , .Q( u1_uk_K_r6_31 ) );
  DFF_X1 u1_uk_K_r6_reg_32 (.CK( clk ) , .D( u1_uk_K_r5_32 ) , .Q( u1_uk_K_r6_32 ) , .QN( u1_uk_n1551 ) );
  DFF_X1 u1_uk_K_r6_reg_33 (.CK( clk ) , .D( u1_uk_K_r5_33 ) , .Q( u1_uk_K_r6_33 ) , .QN( u1_uk_n1552 ) );
  DFF_X1 u1_uk_K_r6_reg_34 (.CK( clk ) , .D( u1_uk_K_r5_34 ) , .Q( u1_uk_K_r6_34 ) );
  DFF_X1 u1_uk_K_r6_reg_35 (.CK( clk ) , .D( u1_uk_K_r5_35 ) , .Q( u1_uk_K_r6_35 ) , .QN( u1_uk_n1554 ) );
  DFF_X1 u1_uk_K_r6_reg_36 (.CK( clk ) , .D( u1_uk_K_r5_36 ) , .Q( u1_uk_K_r6_36 ) , .QN( u1_uk_n1555 ) );
  DFF_X1 u1_uk_K_r6_reg_37 (.CK( clk ) , .D( u1_uk_K_r5_37 ) , .Q( u1_uk_K_r6_37 ) );
  DFF_X1 u1_uk_K_r6_reg_38 (.CK( clk ) , .D( u1_uk_K_r5_38 ) , .Q( u1_uk_K_r6_38 ) , .QN( u1_uk_n1556 ) );
  DFF_X1 u1_uk_K_r6_reg_39 (.CK( clk ) , .D( u1_uk_K_r5_39 ) , .Q( u1_uk_K_r6_39 ) , .QN( u1_uk_n1557 ) );
  DFF_X1 u1_uk_K_r6_reg_4 (.CK( clk ) , .D( u1_uk_K_r5_4 ) , .Q( u1_uk_K_r6_4 ) , .QN( u1_uk_n1530 ) );
  DFF_X1 u1_uk_K_r6_reg_40 (.CK( clk ) , .D( u1_uk_K_r5_40 ) , .Q( u1_uk_K_r6_40 ) , .QN( u1_uk_n1558 ) );
  DFF_X1 u1_uk_K_r6_reg_41 (.CK( clk ) , .D( u1_uk_K_r5_41 ) , .Q( u1_uk_K_r6_41 ) , .QN( u1_uk_n1559 ) );
  DFF_X1 u1_uk_K_r6_reg_42 (.CK( clk ) , .D( u1_uk_K_r5_42 ) , .Q( u1_uk_K_r6_42 ) , .QN( u1_uk_n1560 ) );
  DFF_X1 u1_uk_K_r6_reg_43 (.CK( clk ) , .D( u1_uk_K_r5_43 ) , .Q( u1_uk_K_r6_43 ) , .QN( u1_uk_n1561 ) );
  DFF_X1 u1_uk_K_r6_reg_44 (.CK( clk ) , .D( u1_uk_K_r5_44 ) , .Q( u1_uk_K_r6_44 ) , .QN( u1_uk_n1562 ) );
  DFF_X1 u1_uk_K_r6_reg_45 (.CK( clk ) , .D( u1_uk_K_r5_45 ) , .Q( u1_uk_K_r6_45 ) , .QN( u1_uk_n1563 ) );
  DFF_X1 u1_uk_K_r6_reg_46 (.CK( clk ) , .D( u1_uk_K_r5_46 ) , .Q( u1_uk_K_r6_46 ) );
  DFF_X1 u1_uk_K_r6_reg_47 (.CK( clk ) , .D( u1_uk_K_r5_47 ) , .Q( u1_uk_K_r6_47 ) , .QN( u1_uk_n1564 ) );
  DFF_X1 u1_uk_K_r6_reg_48 (.CK( clk ) , .D( u1_uk_K_r5_48 ) , .Q( u1_uk_K_r6_48 ) , .QN( u1_uk_n1565 ) );
  DFF_X1 u1_uk_K_r6_reg_49 (.CK( clk ) , .D( u1_uk_K_r5_49 ) , .Q( u1_uk_K_r6_49 ) , .QN( u1_uk_n1566 ) );
  DFF_X1 u1_uk_K_r6_reg_5 (.CK( clk ) , .D( u1_uk_K_r5_5 ) , .Q( u1_uk_K_r6_5 ) , .QN( u1_uk_n1531 ) );
  DFF_X1 u1_uk_K_r6_reg_50 (.CK( clk ) , .D( u1_uk_K_r5_50 ) , .Q( u1_uk_K_r6_50 ) , .QN( u1_uk_n1567 ) );
  DFF_X1 u1_uk_K_r6_reg_51 (.CK( clk ) , .D( u1_uk_K_r5_51 ) , .Q( u1_uk_K_r6_51 ) );
  DFF_X1 u1_uk_K_r6_reg_52 (.CK( clk ) , .D( u1_uk_K_r5_52 ) , .Q( u1_uk_K_r6_52 ) , .QN( u1_uk_n1568 ) );
  DFF_X1 u1_uk_K_r6_reg_53 (.CK( clk ) , .D( u1_uk_K_r5_53 ) , .Q( u1_uk_K_r6_53 ) );
  DFF_X1 u1_uk_K_r6_reg_54 (.CK( clk ) , .D( u1_uk_K_r5_54 ) , .Q( u1_uk_K_r6_54 ) , .QN( u1_uk_n1570 ) );
  DFF_X1 u1_uk_K_r6_reg_55 (.CK( clk ) , .D( u1_uk_K_r5_55 ) , .Q( u1_uk_K_r6_55 ) );
  DFF_X1 u1_uk_K_r6_reg_6 (.CK( clk ) , .D( u1_uk_K_r5_6 ) , .Q( u1_uk_K_r6_6 ) , .QN( u1_uk_n1532 ) );
  DFF_X1 u1_uk_K_r6_reg_7 (.CK( clk ) , .D( u1_uk_K_r5_7 ) , .Q( u1_uk_K_r6_7 ) );
  DFF_X1 u1_uk_K_r6_reg_8 (.CK( clk ) , .D( u1_uk_K_r5_8 ) , .Q( u1_uk_K_r6_8 ) , .QN( u1_uk_n1533 ) );
  DFF_X1 u1_uk_K_r6_reg_9 (.CK( clk ) , .D( u1_uk_K_r5_9 ) , .Q( u1_uk_K_r6_9 ) , .QN( u1_uk_n1534 ) );
  DFF_X1 u1_uk_K_r7_reg_0 (.CK( clk ) , .D( u1_uk_K_r6_0 ) , .Q( u1_uk_K_r7_0 ) );
  DFF_X1 u1_uk_K_r7_reg_1 (.CK( clk ) , .D( u1_uk_K_r6_1 ) , .Q( u1_uk_K_r7_1 ) , .QN( u1_uk_n1571 ) );
  DFF_X1 u1_uk_K_r7_reg_10 (.CK( clk ) , .D( u1_uk_K_r6_10 ) , .Q( u1_uk_K_r7_10 ) , .QN( u1_uk_n1577 ) );
  DFF_X1 u1_uk_K_r7_reg_11 (.CK( clk ) , .D( u1_uk_K_r6_11 ) , .Q( u1_uk_K_r7_11 ) , .QN( u1_uk_n1578 ) );
  DFF_X1 u1_uk_K_r7_reg_12 (.CK( clk ) , .D( u1_uk_K_r6_12 ) , .Q( u1_uk_K_r7_12 ) , .QN( u1_uk_n1579 ) );
  DFF_X1 u1_uk_K_r7_reg_13 (.CK( clk ) , .D( u1_uk_K_r6_13 ) , .Q( u1_uk_K_r7_13 ) );
  DFF_X1 u1_uk_K_r7_reg_14 (.CK( clk ) , .D( u1_uk_K_r6_14 ) , .Q( u1_uk_K_r7_14 ) , .QN( u1_uk_n1581 ) );
  DFF_X1 u1_uk_K_r7_reg_15 (.CK( clk ) , .D( u1_uk_K_r6_15 ) , .Q( u1_uk_K_r7_15 ) );
  DFF_X1 u1_uk_K_r7_reg_16 (.CK( clk ) , .D( u1_uk_K_r6_16 ) , .Q( u1_uk_K_r7_16 ) );
  DFF_X1 u1_uk_K_r7_reg_17 (.CK( clk ) , .D( u1_uk_K_r6_17 ) , .Q( u1_uk_K_r7_17 ) , .QN( u1_uk_n1584 ) );
  DFF_X1 u1_uk_K_r7_reg_18 (.CK( clk ) , .D( u1_uk_K_r6_18 ) , .Q( u1_uk_K_r7_18 ) , .QN( u1_uk_n1585 ) );
  DFF_X1 u1_uk_K_r7_reg_19 (.CK( clk ) , .D( u1_uk_K_r6_19 ) , .Q( u1_uk_K_r7_19 ) , .QN( u1_uk_n1586 ) );
  DFF_X1 u1_uk_K_r7_reg_2 (.CK( clk ) , .D( u1_uk_K_r6_2 ) , .Q( u1_uk_K_r7_2 ) , .QN( u1_uk_n1572 ) );
  DFF_X1 u1_uk_K_r7_reg_20 (.CK( clk ) , .D( u1_uk_K_r6_20 ) , .Q( u1_uk_K_r7_20 ) );
  DFF_X1 u1_uk_K_r7_reg_21 (.CK( clk ) , .D( u1_uk_K_r6_21 ) , .Q( u1_uk_K_r7_21 ) , .QN( u1_uk_n1588 ) );
  DFF_X1 u1_uk_K_r7_reg_22 (.CK( clk ) , .D( u1_uk_K_r6_22 ) , .Q( u1_uk_K_r7_22 ) );
  DFF_X1 u1_uk_K_r7_reg_23 (.CK( clk ) , .D( u1_uk_K_r6_23 ) , .Q( u1_uk_K_r7_23 ) );
  DFF_X1 u1_uk_K_r7_reg_24 (.CK( clk ) , .D( u1_uk_K_r6_24 ) , .Q( u1_uk_K_r7_24 ) , .QN( u1_uk_n1592 ) );
  DFF_X1 u1_uk_K_r7_reg_25 (.CK( clk ) , .D( u1_uk_K_r6_25 ) , .Q( u1_uk_K_r7_25 ) , .QN( u1_uk_n1593 ) );
  DFF_X1 u1_uk_K_r7_reg_26 (.CK( clk ) , .D( u1_uk_K_r6_26 ) , .Q( u1_uk_K_r7_26 ) );
  DFF_X1 u1_uk_K_r7_reg_27 (.CK( clk ) , .D( u1_uk_K_r6_27 ) , .Q( u1_uk_K_r7_27 ) );
  DFF_X1 u1_uk_K_r7_reg_28 (.CK( clk ) , .D( u1_uk_K_r6_28 ) , .Q( u1_uk_K_r7_28 ) , .QN( u1_uk_n1595 ) );
  DFF_X1 u1_uk_K_r7_reg_29 (.CK( clk ) , .D( u1_uk_K_r6_29 ) , .Q( u1_uk_K_r7_29 ) );
  DFF_X1 u1_uk_K_r7_reg_3 (.CK( clk ) , .D( u1_uk_K_r6_3 ) , .Q( u1_uk_K_r7_3 ) , .QN( u1_uk_n1573 ) );
  DFF_X1 u1_uk_K_r7_reg_30 (.CK( clk ) , .D( u1_uk_K_r6_30 ) , .Q( u1_uk_K_r7_30 ) );
  DFF_X1 u1_uk_K_r7_reg_31 (.CK( clk ) , .D( u1_uk_K_r6_31 ) , .Q( u1_uk_K_r7_31 ) );
  DFF_X1 u1_uk_K_r7_reg_32 (.CK( clk ) , .D( u1_uk_K_r6_32 ) , .Q( u1_uk_K_r7_32 ) );
  DFF_X1 u1_uk_K_r7_reg_33 (.CK( clk ) , .D( u1_uk_K_r6_33 ) , .Q( u1_uk_K_r7_33 ) , .QN( u1_uk_n1598 ) );
  DFF_X1 u1_uk_K_r7_reg_34 (.CK( clk ) , .D( u1_uk_K_r6_34 ) , .Q( u1_uk_K_r7_34 ) );
  DFF_X1 u1_uk_K_r7_reg_35 (.CK( clk ) , .D( u1_uk_K_r6_35 ) , .Q( u1_uk_K_r7_35 ) , .QN( u1_uk_n1599 ) );
  DFF_X1 u1_uk_K_r7_reg_36 (.CK( clk ) , .D( u1_uk_K_r6_36 ) , .Q( u1_uk_K_r7_36 ) , .QN( u1_uk_n1600 ) );
  DFF_X1 u1_uk_K_r7_reg_37 (.CK( clk ) , .D( u1_uk_K_r6_37 ) , .Q( u1_uk_K_r7_37 ) );
  DFF_X1 u1_uk_K_r7_reg_38 (.CK( clk ) , .D( u1_uk_K_r6_38 ) , .Q( u1_uk_K_r7_38 ) , .QN( u1_uk_n1601 ) );
  DFF_X1 u1_uk_K_r7_reg_39 (.CK( clk ) , .D( u1_uk_K_r6_39 ) , .Q( u1_uk_K_r7_39 ) );
  DFF_X1 u1_uk_K_r7_reg_4 (.CK( clk ) , .D( u1_uk_K_r6_4 ) , .Q( u1_uk_K_r7_4 ) , .QN( u1_uk_n1574 ) );
  DFF_X1 u1_uk_K_r7_reg_40 (.CK( clk ) , .D( u1_uk_K_r6_40 ) , .Q( u1_uk_K_r7_40 ) , .QN( u1_uk_n1603 ) );
  DFF_X1 u1_uk_K_r7_reg_41 (.CK( clk ) , .D( u1_uk_K_r6_41 ) , .Q( u1_uk_K_r7_41 ) , .QN( u1_uk_n1604 ) );
  DFF_X1 u1_uk_K_r7_reg_42 (.CK( clk ) , .D( u1_uk_K_r6_42 ) , .Q( u1_uk_K_r7_42 ) , .QN( u1_uk_n1605 ) );
  DFF_X1 u1_uk_K_r7_reg_43 (.CK( clk ) , .D( u1_uk_K_r6_43 ) , .Q( u1_uk_K_r7_43 ) , .QN( u1_uk_n1606 ) );
  DFF_X1 u1_uk_K_r7_reg_44 (.CK( clk ) , .D( u1_uk_K_r6_44 ) , .Q( u1_uk_K_r7_44 ) , .QN( u1_uk_n1607 ) );
  DFF_X1 u1_uk_K_r7_reg_45 (.CK( clk ) , .D( u1_uk_K_r6_45 ) , .Q( u1_uk_K_r7_45 ) , .QN( u1_uk_n1608 ) );
  DFF_X1 u1_uk_K_r7_reg_46 (.CK( clk ) , .D( u1_uk_K_r6_46 ) , .Q( u1_uk_K_r7_46 ) );
  DFF_X1 u1_uk_K_r7_reg_47 (.CK( clk ) , .D( u1_uk_K_r6_47 ) , .Q( u1_uk_K_r7_47 ) , .QN( u1_uk_n1610 ) );
  DFF_X1 u1_uk_K_r7_reg_48 (.CK( clk ) , .D( u1_uk_K_r6_48 ) , .Q( u1_uk_K_r7_48 ) );
  DFF_X1 u1_uk_K_r7_reg_49 (.CK( clk ) , .D( u1_uk_K_r6_49 ) , .Q( u1_uk_K_r7_49 ) , .QN( u1_uk_n1612 ) );
  DFF_X1 u1_uk_K_r7_reg_5 (.CK( clk ) , .D( u1_uk_K_r6_5 ) , .Q( u1_uk_K_r7_5 ) );
  DFF_X1 u1_uk_K_r7_reg_50 (.CK( clk ) , .D( u1_uk_K_r6_50 ) , .Q( u1_uk_K_r7_50 ) , .QN( u1_uk_n1613 ) );
  DFF_X1 u1_uk_K_r7_reg_51 (.CK( clk ) , .D( u1_uk_K_r6_51 ) , .Q( u1_uk_K_r7_51 ) , .QN( u1_uk_n1614 ) );
  DFF_X1 u1_uk_K_r7_reg_52 (.CK( clk ) , .D( u1_uk_K_r6_52 ) , .Q( u1_uk_K_r7_52 ) , .QN( u1_uk_n1615 ) );
  DFF_X1 u1_uk_K_r7_reg_53 (.CK( clk ) , .D( u1_uk_K_r6_53 ) , .Q( u1_uk_K_r7_53 ) );
  DFF_X1 u1_uk_K_r7_reg_54 (.CK( clk ) , .D( u1_uk_K_r6_54 ) , .Q( u1_uk_K_r7_54 ) , .QN( u1_uk_n1616 ) );
  DFF_X1 u1_uk_K_r7_reg_55 (.CK( clk ) , .D( u1_uk_K_r6_55 ) , .Q( u1_uk_K_r7_55 ) );
  DFF_X1 u1_uk_K_r7_reg_6 (.CK( clk ) , .D( u1_uk_K_r6_6 ) , .Q( u1_uk_K_r7_6 ) );
  DFF_X1 u1_uk_K_r7_reg_7 (.CK( clk ) , .D( u1_uk_K_r6_7 ) , .Q( u1_uk_K_r7_7 ) );
  DFF_X1 u1_uk_K_r7_reg_8 (.CK( clk ) , .D( u1_uk_K_r6_8 ) , .Q( u1_uk_K_r7_8 ) );
  DFF_X1 u1_uk_K_r7_reg_9 (.CK( clk ) , .D( u1_uk_K_r6_9 ) , .Q( u1_uk_K_r7_9 ) );
  DFF_X1 u1_uk_K_r8_reg_0 (.CK( clk ) , .D( u1_uk_K_r7_0 ) , .Q( u1_uk_K_r8_0 ) , .QN( u1_uk_n1618 ) );
  DFF_X1 u1_uk_K_r8_reg_1 (.CK( clk ) , .D( u1_uk_K_r7_1 ) , .Q( u1_uk_K_r8_1 ) , .QN( u1_uk_n1619 ) );
  DFF_X1 u1_uk_K_r8_reg_10 (.CK( clk ) , .D( u1_uk_K_r7_10 ) , .Q( u1_uk_K_r8_10 ) );
  DFF_X1 u1_uk_K_r8_reg_11 (.CK( clk ) , .D( u1_uk_K_r7_11 ) , .Q( u1_uk_K_r8_11 ) , .QN( u1_uk_n1625 ) );
  DFF_X1 u1_uk_K_r8_reg_12 (.CK( clk ) , .D( u1_uk_K_r7_12 ) , .Q( u1_uk_K_r8_12 ) , .QN( u1_uk_n1626 ) );
  DFF_X1 u1_uk_K_r8_reg_13 (.CK( clk ) , .D( u1_uk_K_r7_13 ) , .Q( u1_uk_K_r8_13 ) );
  DFF_X1 u1_uk_K_r8_reg_14 (.CK( clk ) , .D( u1_uk_K_r7_14 ) , .Q( u1_uk_K_r8_14 ) , .QN( u1_uk_n1627 ) );
  DFF_X1 u1_uk_K_r8_reg_15 (.CK( clk ) , .D( u1_uk_K_r7_15 ) , .Q( u1_uk_K_r8_15 ) , .QN( u1_uk_n1628 ) );
  DFF_X1 u1_uk_K_r8_reg_16 (.CK( clk ) , .D( u1_uk_K_r7_16 ) , .Q( u1_uk_K_r8_16 ) );
  DFF_X1 u1_uk_K_r8_reg_17 (.CK( clk ) , .D( u1_uk_K_r7_17 ) , .Q( u1_uk_K_r8_17 ) );
  DFF_X1 u1_uk_K_r8_reg_18 (.CK( clk ) , .D( u1_uk_K_r7_18 ) , .Q( u1_uk_K_r8_18 ) , .QN( u1_uk_n1629 ) );
  DFF_X1 u1_uk_K_r8_reg_19 (.CK( clk ) , .D( u1_uk_K_r7_19 ) , .Q( u1_uk_K_r8_19 ) );
  DFF_X1 u1_uk_K_r8_reg_2 (.CK( clk ) , .D( u1_uk_K_r7_2 ) , .Q( u1_uk_K_r8_2 ) );
  DFF_X1 u1_uk_K_r8_reg_20 (.CK( clk ) , .D( u1_uk_K_r7_20 ) , .Q( u1_uk_K_r8_20 ) , .QN( u1_uk_n1630 ) );
  DFF_X1 u1_uk_K_r8_reg_21 (.CK( clk ) , .D( u1_uk_K_r7_21 ) , .Q( u1_uk_K_r8_21 ) );
  DFF_X1 u1_uk_K_r8_reg_22 (.CK( clk ) , .D( u1_uk_K_r7_22 ) , .Q( u1_uk_K_r8_22 ) );
  DFF_X1 u1_uk_K_r8_reg_23 (.CK( clk ) , .D( u1_uk_K_r7_23 ) , .Q( u1_uk_K_r8_23 ) , .QN( u1_uk_n1632 ) );
  DFF_X1 u1_uk_K_r8_reg_24 (.CK( clk ) , .D( u1_uk_K_r7_24 ) , .Q( u1_uk_K_r8_24 ) , .QN( u1_uk_n1633 ) );
  DFF_X1 u1_uk_K_r8_reg_25 (.CK( clk ) , .D( u1_uk_K_r7_25 ) , .Q( u1_uk_K_r8_25 ) , .QN( u1_uk_n1634 ) );
  DFF_X1 u1_uk_K_r8_reg_26 (.CK( clk ) , .D( u1_uk_K_r7_26 ) , .Q( u1_uk_K_r8_26 ) , .QN( u1_uk_n1635 ) );
  DFF_X1 u1_uk_K_r8_reg_27 (.CK( clk ) , .D( u1_uk_K_r7_27 ) , .Q( u1_uk_K_r8_27 ) );
  DFF_X1 u1_uk_K_r8_reg_28 (.CK( clk ) , .D( u1_uk_K_r7_28 ) , .Q( u1_uk_K_r8_28 ) );
  DFF_X1 u1_uk_K_r8_reg_29 (.CK( clk ) , .D( u1_uk_K_r7_29 ) , .Q( u1_uk_K_r8_29 ) , .QN( u1_uk_n1639 ) );
  DFF_X1 u1_uk_K_r8_reg_3 (.CK( clk ) , .D( u1_uk_K_r7_3 ) , .Q( u1_uk_K_r8_3 ) , .QN( u1_uk_n1620 ) );
  DFF_X1 u1_uk_K_r8_reg_30 (.CK( clk ) , .D( u1_uk_K_r7_30 ) , .Q( u1_uk_K_r8_30 ) , .QN( u1_uk_n1640 ) );
  DFF_X1 u1_uk_K_r8_reg_31 (.CK( clk ) , .D( u1_uk_K_r7_31 ) , .Q( u1_uk_K_r8_31 ) , .QN( u1_uk_n1641 ) );
  DFF_X1 u1_uk_K_r8_reg_32 (.CK( clk ) , .D( u1_uk_K_r7_32 ) , .Q( u1_uk_K_r8_32 ) );
  DFF_X1 u1_uk_K_r8_reg_33 (.CK( clk ) , .D( u1_uk_K_r7_33 ) , .Q( u1_uk_K_r8_33 ) , .QN( u1_uk_n1642 ) );
  DFF_X1 u1_uk_K_r8_reg_34 (.CK( clk ) , .D( u1_uk_K_r7_34 ) , .Q( u1_uk_K_r8_34 ) , .QN( u1_uk_n1643 ) );
  DFF_X1 u1_uk_K_r8_reg_35 (.CK( clk ) , .D( u1_uk_K_r7_35 ) , .Q( u1_uk_K_r8_35 ) , .QN( u1_uk_n1644 ) );
  DFF_X1 u1_uk_K_r8_reg_36 (.CK( clk ) , .D( u1_uk_K_r7_36 ) , .Q( u1_uk_K_r8_36 ) , .QN( u1_uk_n1645 ) );
  DFF_X1 u1_uk_K_r8_reg_37 (.CK( clk ) , .D( u1_uk_K_r7_37 ) , .Q( u1_uk_K_r8_37 ) );
  DFF_X1 u1_uk_K_r8_reg_38 (.CK( clk ) , .D( u1_uk_K_r7_38 ) , .Q( u1_uk_K_r8_38 ) , .QN( u1_uk_n1647 ) );
  DFF_X1 u1_uk_K_r8_reg_39 (.CK( clk ) , .D( u1_uk_K_r7_39 ) , .Q( u1_uk_K_r8_39 ) , .QN( u1_uk_n1649 ) );
  DFF_X1 u1_uk_K_r8_reg_4 (.CK( clk ) , .D( u1_uk_K_r7_4 ) , .Q( u1_uk_K_r8_4 ) , .QN( u1_uk_n1621 ) );
  DFF_X1 u1_uk_K_r8_reg_40 (.CK( clk ) , .D( u1_uk_K_r7_40 ) , .Q( u1_uk_K_r8_40 ) );
  DFF_X1 u1_uk_K_r8_reg_41 (.CK( clk ) , .D( u1_uk_K_r7_41 ) , .Q( u1_uk_K_r8_41 ) );
  DFF_X1 u1_uk_K_r8_reg_42 (.CK( clk ) , .D( u1_uk_K_r7_42 ) , .Q( u1_uk_K_r8_42 ) , .QN( u1_uk_n1651 ) );
  DFF_X1 u1_uk_K_r8_reg_43 (.CK( clk ) , .D( u1_uk_K_r7_43 ) , .Q( u1_uk_K_r8_43 ) );
  DFF_X1 u1_uk_K_r8_reg_44 (.CK( clk ) , .D( u1_uk_K_r7_44 ) , .Q( u1_uk_K_r8_44 ) , .QN( u1_uk_n1652 ) );
  DFF_X1 u1_uk_K_r8_reg_45 (.CK( clk ) , .D( u1_uk_K_r7_45 ) , .Q( u1_uk_K_r8_45 ) );
  DFF_X1 u1_uk_K_r8_reg_46 (.CK( clk ) , .D( u1_uk_K_r7_46 ) , .Q( u1_uk_K_r8_46 ) , .QN( u1_uk_n1653 ) );
  DFF_X1 u1_uk_K_r8_reg_47 (.CK( clk ) , .D( u1_uk_K_r7_47 ) , .Q( u1_uk_K_r8_47 ) , .QN( u1_uk_n1654 ) );
  DFF_X1 u1_uk_K_r8_reg_48 (.CK( clk ) , .D( u1_uk_K_r7_48 ) , .Q( u1_uk_K_r8_48 ) );
  DFF_X1 u1_uk_K_r8_reg_49 (.CK( clk ) , .D( u1_uk_K_r7_49 ) , .Q( u1_uk_K_r8_49 ) , .QN( u1_uk_n1655 ) );
  DFF_X1 u1_uk_K_r8_reg_5 (.CK( clk ) , .D( u1_uk_K_r7_5 ) , .Q( u1_uk_K_r8_5 ) );
  DFF_X1 u1_uk_K_r8_reg_50 (.CK( clk ) , .D( u1_uk_K_r7_50 ) , .Q( u1_uk_K_r8_50 ) , .QN( u1_uk_n1656 ) );
  DFF_X1 u1_uk_K_r8_reg_51 (.CK( clk ) , .D( u1_uk_K_r7_51 ) , .Q( u1_uk_K_r8_51 ) );
  DFF_X1 u1_uk_K_r8_reg_52 (.CK( clk ) , .D( u1_uk_K_r7_52 ) , .Q( u1_uk_K_r8_52 ) );
  DFF_X1 u1_uk_K_r8_reg_53 (.CK( clk ) , .D( u1_uk_K_r7_53 ) , .Q( u1_uk_K_r8_53 ) , .QN( u1_uk_n1659 ) );
  DFF_X1 u1_uk_K_r8_reg_54 (.CK( clk ) , .D( u1_uk_K_r7_54 ) , .Q( u1_uk_K_r8_54 ) , .QN( u1_uk_n1660 ) );
  DFF_X1 u1_uk_K_r8_reg_55 (.CK( clk ) , .D( u1_uk_K_r7_55 ) , .Q( u1_uk_K_r8_55 ) , .QN( u1_uk_n1661 ) );
  DFF_X1 u1_uk_K_r8_reg_6 (.CK( clk ) , .D( u1_uk_K_r7_6 ) , .Q( u1_uk_K_r8_6 ) , .QN( u1_uk_n1622 ) );
  DFF_X1 u1_uk_K_r8_reg_7 (.CK( clk ) , .D( u1_uk_K_r7_7 ) , .Q( u1_uk_K_r8_7 ) , .QN( u1_uk_n1623 ) );
  DFF_X1 u1_uk_K_r8_reg_8 (.CK( clk ) , .D( u1_uk_K_r7_8 ) , .Q( u1_uk_K_r8_8 ) );
  DFF_X1 u1_uk_K_r8_reg_9 (.CK( clk ) , .D( u1_uk_K_r7_9 ) , .Q( u1_uk_K_r8_9 ) , .QN( u1_uk_n1624 ) );
  DFF_X1 u1_uk_K_r9_reg_0 (.CK( clk ) , .D( u1_uk_K_r8_0 ) , .Q( u1_uk_K_r9_0 ) );
  DFF_X1 u1_uk_K_r9_reg_1 (.CK( clk ) , .D( u1_uk_K_r8_1 ) , .Q( u1_uk_K_r9_1 ) , .QN( u1_uk_n1662 ) );
  DFF_X1 u1_uk_K_r9_reg_10 (.CK( clk ) , .D( u1_uk_K_r8_10 ) , .Q( u1_uk_K_r9_10 ) );
  DFF_X1 u1_uk_K_r9_reg_11 (.CK( clk ) , .D( u1_uk_K_r8_11 ) , .Q( u1_uk_K_r9_11 ) , .QN( u1_uk_n1667 ) );
  DFF_X1 u1_uk_K_r9_reg_12 (.CK( clk ) , .D( u1_uk_K_r8_12 ) , .Q( u1_uk_K_r9_12 ) );
  DFF_X1 u1_uk_K_r9_reg_13 (.CK( clk ) , .D( u1_uk_K_r8_13 ) , .Q( u1_uk_K_r9_13 ) , .QN( u1_uk_n1669 ) );
  DFF_X1 u1_uk_K_r9_reg_14 (.CK( clk ) , .D( u1_uk_K_r8_14 ) , .Q( u1_uk_K_r9_14 ) , .QN( u1_uk_n1670 ) );
  DFF_X1 u1_uk_K_r9_reg_15 (.CK( clk ) , .D( u1_uk_K_r8_15 ) , .Q( u1_uk_K_r9_15 ) );
  DFF_X1 u1_uk_K_r9_reg_16 (.CK( clk ) , .D( u1_uk_K_r8_16 ) , .Q( u1_uk_K_r9_16 ) , .QN( u1_uk_n1672 ) );
  DFF_X1 u1_uk_K_r9_reg_17 (.CK( clk ) , .D( u1_uk_K_r8_17 ) , .Q( u1_uk_K_r9_17 ) , .QN( u1_uk_n1673 ) );
  DFF_X1 u1_uk_K_r9_reg_18 (.CK( clk ) , .D( u1_uk_K_r8_18 ) , .Q( u1_uk_K_r9_18 ) );
  DFF_X1 u1_uk_K_r9_reg_19 (.CK( clk ) , .D( u1_uk_K_r8_19 ) , .Q( u1_uk_K_r9_19 ) );
  DFF_X1 u1_uk_K_r9_reg_2 (.CK( clk ) , .D( u1_uk_K_r8_2 ) , .Q( u1_uk_K_r9_2 ) );
  DFF_X1 u1_uk_K_r9_reg_20 (.CK( clk ) , .D( u1_uk_K_r8_20 ) , .Q( u1_uk_K_r9_20 ) , .QN( u1_uk_n1676 ) );
  DFF_X1 u1_uk_K_r9_reg_21 (.CK( clk ) , .D( u1_uk_K_r8_21 ) , .Q( u1_uk_K_r9_21 ) , .QN( u1_uk_n1677 ) );
  DFF_X1 u1_uk_K_r9_reg_22 (.CK( clk ) , .D( u1_uk_K_r8_22 ) , .Q( u1_uk_K_r9_22 ) , .QN( u1_uk_n1678 ) );
  DFF_X1 u1_uk_K_r9_reg_23 (.CK( clk ) , .D( u1_uk_K_r8_23 ) , .Q( u1_uk_K_r9_23 ) );
  DFF_X1 u1_uk_K_r9_reg_24 (.CK( clk ) , .D( u1_uk_K_r8_24 ) , .Q( u1_uk_K_r9_24 ) );
  DFF_X1 u1_uk_K_r9_reg_25 (.CK( clk ) , .D( u1_uk_K_r8_25 ) , .Q( u1_uk_K_r9_25 ) );
  DFF_X1 u1_uk_K_r9_reg_26 (.CK( clk ) , .D( u1_uk_K_r8_26 ) , .Q( u1_uk_K_r9_26 ) , .QN( u1_uk_n1682 ) );
  DFF_X1 u1_uk_K_r9_reg_27 (.CK( clk ) , .D( u1_uk_K_r8_27 ) , .Q( u1_uk_K_r9_27 ) );
  DFF_X1 u1_uk_K_r9_reg_28 (.CK( clk ) , .D( u1_uk_K_r8_28 ) , .Q( u1_uk_K_r9_28 ) , .QN( u1_uk_n1683 ) );
  DFF_X1 u1_uk_K_r9_reg_29 (.CK( clk ) , .D( u1_uk_K_r8_29 ) , .Q( u1_uk_K_r9_29 ) , .QN( u1_uk_n1684 ) );
  DFF_X1 u1_uk_K_r9_reg_3 (.CK( clk ) , .D( u1_uk_K_r8_3 ) , .Q( u1_uk_K_r9_3 ) , .QN( u1_uk_n1663 ) );
  DFF_X1 u1_uk_K_r9_reg_30 (.CK( clk ) , .D( u1_uk_K_r8_30 ) , .Q( u1_uk_K_r9_30 ) );
  DFF_X1 u1_uk_K_r9_reg_31 (.CK( clk ) , .D( u1_uk_K_r8_31 ) , .Q( u1_uk_K_r9_31 ) );
  DFF_X1 u1_uk_K_r9_reg_32 (.CK( clk ) , .D( u1_uk_K_r8_32 ) , .Q( u1_uk_K_r9_32 ) , .QN( u1_uk_n1687 ) );
  DFF_X1 u1_uk_K_r9_reg_33 (.CK( clk ) , .D( u1_uk_K_r8_33 ) , .Q( u1_uk_K_r9_33 ) );
  DFF_X1 u1_uk_K_r9_reg_34 (.CK( clk ) , .D( u1_uk_K_r8_34 ) , .Q( u1_uk_K_r9_34 ) , .QN( u1_uk_n1688 ) );
  DFF_X1 u1_uk_K_r9_reg_35 (.CK( clk ) , .D( u1_uk_K_r8_35 ) , .Q( u1_uk_K_r9_35 ) );
  DFF_X1 u1_uk_K_r9_reg_36 (.CK( clk ) , .D( u1_uk_K_r8_36 ) , .Q( u1_uk_K_r9_36 ) , .QN( u1_uk_n1689 ) );
  DFF_X1 u1_uk_K_r9_reg_37 (.CK( clk ) , .D( u1_uk_K_r8_37 ) , .Q( u1_uk_K_r9_37 ) , .QN( u1_uk_n1690 ) );
  DFF_X1 u1_uk_K_r9_reg_38 (.CK( clk ) , .D( u1_uk_K_r8_38 ) , .Q( u1_uk_K_r9_38 ) );
  DFF_X1 u1_uk_K_r9_reg_39 (.CK( clk ) , .D( u1_uk_K_r8_39 ) , .Q( u1_uk_K_r9_39 ) , .QN( u1_uk_n1691 ) );
  DFF_X1 u1_uk_K_r9_reg_4 (.CK( clk ) , .D( u1_uk_K_r8_4 ) , .Q( u1_uk_K_r9_4 ) );
  DFF_X1 u1_uk_K_r9_reg_40 (.CK( clk ) , .D( u1_uk_K_r8_40 ) , .Q( u1_uk_K_r9_40 ) , .QN( u1_uk_n1692 ) );
  DFF_X1 u1_uk_K_r9_reg_41 (.CK( clk ) , .D( u1_uk_K_r8_41 ) , .Q( u1_uk_K_r9_41 ) , .QN( u1_uk_n1693 ) );
  DFF_X1 u1_uk_K_r9_reg_42 (.CK( clk ) , .D( u1_uk_K_r8_42 ) , .Q( u1_uk_K_r9_42 ) , .QN( u1_uk_n1694 ) );
  DFF_X1 u1_uk_K_r9_reg_43 (.CK( clk ) , .D( u1_uk_K_r8_43 ) , .Q( u1_uk_K_r9_43 ) , .QN( u1_uk_n1695 ) );
  DFF_X1 u1_uk_K_r9_reg_44 (.CK( clk ) , .D( u1_uk_K_r8_44 ) , .Q( u1_uk_K_r9_44 ) , .QN( u1_uk_n1696 ) );
  DFF_X1 u1_uk_K_r9_reg_45 (.CK( clk ) , .D( u1_uk_K_r8_45 ) , .Q( u1_uk_K_r9_45 ) );
  DFF_X1 u1_uk_K_r9_reg_46 (.CK( clk ) , .D( u1_uk_K_r8_46 ) , .Q( u1_uk_K_r9_46 ) , .QN( u1_uk_n1698 ) );
  DFF_X1 u1_uk_K_r9_reg_47 (.CK( clk ) , .D( u1_uk_K_r8_47 ) , .Q( u1_uk_K_r9_47 ) , .QN( u1_uk_n1699 ) );
  DFF_X1 u1_uk_K_r9_reg_48 (.CK( clk ) , .D( u1_uk_K_r8_48 ) , .Q( u1_uk_K_r9_48 ) );
  DFF_X1 u1_uk_K_r9_reg_49 (.CK( clk ) , .D( u1_uk_K_r8_49 ) , .Q( u1_uk_K_r9_49 ) );
  DFF_X1 u1_uk_K_r9_reg_5 (.CK( clk ) , .D( u1_uk_K_r8_5 ) , .Q( u1_uk_K_r9_5 ) );
  DFF_X1 u1_uk_K_r9_reg_50 (.CK( clk ) , .D( u1_uk_K_r8_50 ) , .Q( u1_uk_K_r9_50 ) , .QN( u1_uk_n1702 ) );
  DFF_X1 u1_uk_K_r9_reg_51 (.CK( clk ) , .D( u1_uk_K_r8_51 ) , .Q( u1_uk_K_r9_51 ) , .QN( u1_uk_n1703 ) );
  DFF_X1 u1_uk_K_r9_reg_52 (.CK( clk ) , .D( u1_uk_K_r8_52 ) , .Q( u1_uk_K_r9_52 ) , .QN( u1_uk_n1704 ) );
  DFF_X1 u1_uk_K_r9_reg_53 (.CK( clk ) , .D( u1_uk_K_r8_53 ) , .Q( u1_uk_K_r9_53 ) , .QN( u1_uk_n1705 ) );
  DFF_X1 u1_uk_K_r9_reg_54 (.CK( clk ) , .D( u1_uk_K_r8_54 ) , .Q( u1_uk_K_r9_54 ) );
  DFF_X1 u1_uk_K_r9_reg_55 (.CK( clk ) , .D( u1_uk_K_r8_55 ) , .Q( u1_uk_K_r9_55 ) , .QN( u1_uk_n1707 ) );
  DFF_X1 u1_uk_K_r9_reg_6 (.CK( clk ) , .D( u1_uk_K_r8_6 ) , .Q( u1_uk_K_r9_6 ) );
  DFF_X1 u1_uk_K_r9_reg_7 (.CK( clk ) , .D( u1_uk_K_r8_7 ) , .Q( u1_uk_K_r9_7 ) );
  DFF_X1 u1_uk_K_r9_reg_8 (.CK( clk ) , .D( u1_uk_K_r8_8 ) , .Q( u1_uk_K_r9_8 ) , .QN( u1_uk_n1664 ) );
  DFF_X1 u1_uk_K_r9_reg_9 (.CK( clk ) , .D( u1_uk_K_r8_9 ) , .Q( u1_uk_K_r9_9 ) );
  INV_X1 u1_uk_U10 (.A( u1_uk_n209 ) , .ZN( u1_uk_n83 ) );
  AOI22_X1 u1_uk_U100 (.B2( u1_uk_K_r0_28 ) , .A2( u1_uk_K_r0_49 ) , .ZN( u1_uk_n1031 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1000 (.ZN( u1_K6_23 ) , .A( u1_uk_n1093 ) , .B2( u1_uk_n1472 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1001 (.A1( u1_uk_K_r4_27 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1093 ) );
  OAI21_X1 u1_uk_U1002 (.ZN( u1_K3_35 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1042 ) , .B2( u1_uk_n1308 ) );
  NAND2_X1 u1_uk_U1003 (.A1( u1_uk_K_r1_7 ) , .ZN( u1_uk_n1042 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U1004 (.ZN( u1_K14_46 ) , .B2( u1_uk_n1820 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n961 ) );
  NAND2_X1 u1_uk_U1005 (.A1( u1_uk_K_r12_22 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n961 ) );
  OAI21_X1 u1_uk_U1006 (.ZN( u1_K16_4 ) , .B2( u1_uk_n1257 ) , .B1( u1_uk_n99 ) , .A( u1_uk_n995 ) );
  NAND2_X1 u1_uk_U1007 (.A1( u1_uk_K_r14_3 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n995 ) );
  OAI21_X1 u1_uk_U1008 (.ZN( u1_K8_4 ) , .A( u1_uk_n1146 ) , .B2( u1_uk_n1537 ) , .B1( u1_uk_n17 ) );
  NAND2_X1 u1_uk_U1009 (.A1( u1_uk_K_r6_19 ) , .ZN( u1_uk_n1146 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U101 (.ZN( u1_K15_41 ) , .B2( u1_uk_n1865 ) , .A2( u1_uk_n1883 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1010 (.ZN( u1_K5_4 ) , .A( u1_uk_n1085 ) , .B2( u1_uk_n1411 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1011 (.A1( u1_uk_K_r3_4 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1085 ) );
  OAI21_X1 u1_uk_U1012 (.ZN( u1_K4_5 ) , .A( u1_uk_n1068 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1386 ) );
  NAND2_X1 u1_uk_U1013 (.A1( u1_uk_K_r2_53 ) , .ZN( u1_uk_n1068 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1014 (.ZN( u1_K3_5 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1048 ) , .B2( u1_uk_n1332 ) );
  NAND2_X1 u1_uk_U1015 (.A1( u1_uk_K_r1_10 ) , .ZN( u1_uk_n1048 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1016 (.ZN( u1_K5_45 ) , .A( u1_uk_n1084 ) , .B2( u1_uk_n1400 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1017 (.A1( u1_uk_K_r3_43 ) , .ZN( u1_uk_n1084 ) , .A2( u1_uk_n11 ) );
  OAI21_X1 u1_uk_U1018 (.ZN( u1_K3_45 ) , .A( u1_uk_n1046 ) , .B2( u1_uk_n1335 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U1019 (.A1( u1_uk_K_r1_16 ) , .ZN( u1_uk_n1046 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U102 (.ZN( u1_K13_41 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1753 ) , .A2( u1_uk_n1768 ) , .A1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U1020 (.ZN( u1_K1_13 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1214 ) , .A( u1_uk_n999 ) );
  NAND2_X1 u1_uk_U1021 (.A1( u1_key_r_46 ) , .A2( u1_uk_n146 ) , .ZN( u1_uk_n999 ) );
  OAI21_X1 u1_uk_U1022 (.ZN( u1_K1_17 ) , .A( u1_uk_n1001 ) , .B2( u1_uk_n1183 ) , .B1( u1_uk_n129 ) );
  NAND2_X1 u1_uk_U1023 (.A1( u1_key_r_10 ) , .ZN( u1_uk_n1001 ) , .A2( u1_uk_n187 ) );
  OAI21_X1 u1_uk_U1024 (.ZN( u1_K10_21 ) , .B2( u1_uk_n1660 ) , .A( u1_uk_n308 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1025 (.A1( u1_uk_K_r8_19 ) , .ZN( u1_uk_n308 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1026 (.ZN( u1_K1_37 ) , .A( u1_uk_n1013 ) , .B2( u1_uk_n1174 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U1027 (.A1( u1_key_r_50 ) , .ZN( u1_uk_n1013 ) , .A2( u1_uk_n162 ) );
  OAI21_X1 u1_uk_U1028 (.ZN( u1_K9_39 ) , .A( u1_uk_n1165 ) , .B2( u1_uk_n1601 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1029 (.A1( u1_uk_K_r7_31 ) , .ZN( u1_uk_n1165 ) , .A2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U103 (.ZN( u1_K7_41 ) , .A2( u1_uk_n1486 ) , .B2( u1_uk_n1516 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U1030 (.ZN( u1_K14_44 ) , .B2( u1_uk_n1807 ) , .B1( u1_uk_n251 ) , .A( u1_uk_n959 ) );
  NAND2_X1 u1_uk_U1031 (.A1( u1_uk_K_r12_15 ) , .A2( u1_uk_n279 ) , .ZN( u1_uk_n959 ) );
  OAI21_X1 u1_uk_U1032 (.ZN( u1_K9_44 ) , .A( u1_uk_n1168 ) , .B2( u1_uk_n1615 ) , .B1( u1_uk_n223 ) );
  NAND2_X1 u1_uk_U1033 (.A1( u1_uk_K_r7_0 ) , .ZN( u1_uk_n1168 ) , .A2( u1_uk_n207 ) );
  OAI21_X1 u1_uk_U1034 (.ZN( u1_K12_6 ) , .B2( u1_uk_n1732 ) , .B1( u1_uk_n230 ) , .A( u1_uk_n662 ) );
  NAND2_X1 u1_uk_U1035 (.A1( u1_uk_K_r10_10 ) , .A2( u1_uk_n251 ) , .ZN( u1_uk_n662 ) );
  OAI21_X1 u1_uk_U1036 (.ZN( u1_K8_46 ) , .A( u1_uk_n1145 ) , .B2( u1_uk_n1562 ) , .B1( u1_uk_n188 ) );
  NAND2_X1 u1_uk_U1037 (.A1( u1_uk_K_r6_37 ) , .ZN( u1_uk_n1145 ) , .A2( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U1038 (.ZN( u1_K10_13 ) , .B2( u1_uk_n1635 ) , .A( u1_uk_n301 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1039 (.A1( u1_uk_K_r8_48 ) , .ZN( u1_uk_n301 ) , .A2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U104 (.ZN( u1_K4_41 ) , .B2( u1_uk_n1349 ) , .A2( u1_uk_n1366 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U1040 (.ZN( u1_K12_36 ) , .B2( u1_uk_n1728 ) , .A( u1_uk_n587 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1041 (.A1( u1_uk_K_r10_52 ) , .A2( u1_uk_n110 ) , .ZN( u1_uk_n587 ) );
  OAI21_X1 u1_uk_U1042 (.ZN( u1_K16_41 ) , .B2( u1_uk_n1245 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n991 ) );
  NAND2_X1 u1_uk_U1043 (.A1( u1_uk_K_r14_42 ) , .A2( u1_uk_n141 ) , .ZN( u1_uk_n991 ) );
  OAI21_X1 u1_uk_U1044 (.ZN( u1_K8_41 ) , .A( u1_uk_n1141 ) , .B2( u1_uk_n1547 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U1045 (.A1( u1_uk_K_r6_30 ) , .ZN( u1_uk_n1141 ) , .A2( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U1046 (.ZN( u1_K6_41 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1099 ) , .B2( u1_uk_n1475 ) );
  NAND2_X1 u1_uk_U1047 (.A1( u1_uk_K_r4_31 ) , .ZN( u1_uk_n1099 ) , .A2( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1048 (.ZN( u1_K16_28 ) , .B2( u1_uk_n1219 ) , .A( u1_uk_n984 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1049 (.A1( u1_uk_K_r14_8 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n984 ) );
  OAI21_X1 u1_uk_U1050 (.ZN( u1_K8_28 ) , .A( u1_uk_n1133 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1562 ) );
  NAND2_X1 u1_uk_U1051 (.A1( u1_uk_K_r6_51 ) , .ZN( u1_uk_n1133 ) , .A2( u1_uk_n145 ) );
  OAI21_X1 u1_uk_U1052 (.ZN( u1_K4_28 ) , .A( u1_uk_n1059 ) , .B2( u1_uk_n1381 ) , .B1( u1_uk_n148 ) );
  NAND2_X1 u1_uk_U1053 (.A1( u1_uk_K_r2_21 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1059 ) );
  OAI21_X1 u1_uk_U1054 (.ZN( u1_K9_14 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1151 ) , .B2( u1_uk_n1604 ) );
  NAND2_X1 u1_uk_U1055 (.A1( u1_uk_K_r7_34 ) , .A2( u1_uk_n100 ) , .ZN( u1_uk_n1151 ) );
  OAI21_X1 u1_uk_U1056 (.ZN( u1_K7_31 ) , .A( u1_uk_n1117 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1508 ) );
  NAND2_X1 u1_uk_U1057 (.A1( u1_uk_K_r5_16 ) , .ZN( u1_uk_n1117 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1058 (.ZN( u1_K14_40 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1823 ) , .A( u1_uk_n958 ) );
  NAND2_X1 u1_uk_U1059 (.A1( u1_uk_K_r12_21 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n958 ) );
  AOI22_X1 u1_uk_U106 (.B2( u1_uk_K_r9_19 ) , .A2( u1_uk_K_r9_25 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n250 ) , .ZN( u1_uk_n496 ) );
  OAI21_X1 u1_uk_U1060 (.ZN( u1_K12_40 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1729 ) , .A( u1_uk_n603 ) );
  NAND2_X1 u1_uk_U1061 (.A1( u1_uk_K_r10_49 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n603 ) );
  OAI21_X1 u1_uk_U1062 (.ZN( u1_K15_14 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1851 ) , .A( u1_uk_n966 ) );
  NAND2_X1 u1_uk_U1063 (.A1( u1_uk_K_r13_32 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n966 ) );
  OAI21_X1 u1_uk_U1064 (.ZN( u1_K10_32 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1618 ) , .A( u1_uk_n346 ) );
  NAND2_X1 u1_uk_U1065 (.A1( u1_uk_K_r8_51 ) , .A2( u1_uk_n142 ) , .ZN( u1_uk_n346 ) );
  OAI21_X1 u1_uk_U1066 (.ZN( u1_K15_32 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1855 ) , .A( u1_uk_n971 ) );
  NAND2_X1 u1_uk_U1067 (.A1( u1_uk_K_r13_36 ) , .A2( u1_uk_n147 ) , .ZN( u1_uk_n971 ) );
  OAI21_X1 u1_uk_U1068 (.ZN( u1_K16_42 ) , .B2( u1_uk_n1241 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n992 ) );
  NAND2_X1 u1_uk_U1069 (.A1( u1_uk_K_r14_38 ) , .A2( u1_uk_n31 ) , .ZN( u1_uk_n992 ) );
  OAI22_X1 u1_uk_U107 (.ZN( u1_K1_5 ) , .A2( u1_uk_n1176 ) , .B2( u1_uk_n1180 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U1070 (.ZN( u1_K8_42 ) , .A( u1_uk_n1142 ) , .B2( u1_uk_n1540 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U1071 (.A1( u1_uk_K_r6_22 ) , .ZN( u1_uk_n1142 ) , .A2( u1_uk_n117 ) );
  OAI21_X1 u1_uk_U1072 (.ZN( u1_K7_38 ) , .A( u1_uk_n1122 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1499 ) );
  NAND2_X1 u1_uk_U1073 (.A1( u1_uk_K_r5_8 ) , .ZN( u1_uk_n1122 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1074 (.ZN( u1_K5_42 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1082 ) , .B2( u1_uk_n1412 ) );
  NAND2_X1 u1_uk_U1075 (.A1( u1_uk_K_r3_9 ) , .ZN( u1_uk_n1082 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1076 (.ZN( u1_K4_38 ) , .A( u1_uk_n1064 ) , .B2( u1_uk_n1383 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U1077 (.A1( u1_uk_K_r2_50 ) , .ZN( u1_uk_n1064 ) , .A2( u1_uk_n155 ) );
  INV_X1 u1_uk_U1078 (.A( u1_key_r_9 ) , .ZN( u1_uk_n1179 ) );
  INV_X1 u1_uk_U1079 (.A( u1_key_r_7 ) , .ZN( u1_uk_n1177 ) );
  OAI22_X1 u1_uk_U108 (.ZN( u1_K16_5 ) , .A2( u1_uk_n1221 ) , .B2( u1_uk_n1224 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n294 ) );
  INV_X1 u1_uk_U1080 (.A( u1_key_r_6 ) , .ZN( u1_uk_n1176 ) );
  INV_X1 u1_uk_U1081 (.A( u1_key_r_54 ) , .ZN( u1_uk_n1215 ) );
  INV_X1 u1_uk_U1082 (.A( u1_key_r_33 ) , .ZN( u1_uk_n1197 ) );
  INV_X1 u1_uk_U1083 (.A( u1_key_r_23 ) , .ZN( u1_uk_n1188 ) );
  INV_X1 u1_uk_U1084 (.A( u1_key_r_26 ) , .ZN( u1_uk_n1191 ) );
  INV_X1 u1_uk_U1085 (.A( u1_key_r_40 ) , .ZN( u1_uk_n1204 ) );
  INV_X1 u1_uk_U1086 (.A( u1_key_r_30 ) , .ZN( u1_uk_n1195 ) );
  INV_X1 u1_uk_U1087 (.A( u1_key_r_47 ) , .ZN( u1_uk_n1209 ) );
  INV_X1 u1_uk_U1088 (.A( u1_key_r_34 ) , .ZN( u1_uk_n1198 ) );
  INV_X1 u1_uk_U1089 (.A( u1_key_r_27 ) , .ZN( u1_uk_n1192 ) );
  OAI22_X1 u1_uk_U109 (.ZN( u1_K15_5 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1859 ) , .A2( u1_uk_n1862 ) , .B1( u1_uk_n217 ) );
  INV_X1 u1_uk_U1090 (.A( u1_key_r_24 ) , .ZN( u1_uk_n1189 ) );
  INV_X1 u1_uk_U1091 (.A( u1_key_r_20 ) , .ZN( u1_uk_n1185 ) );
  INV_X1 u1_uk_U1092 (.A( u1_key_r_37 ) , .ZN( u1_uk_n1201 ) );
  INV_X1 u1_uk_U1093 (.A( u1_key_r_52 ) , .ZN( u1_uk_n1213 ) );
  INV_X1 u1_uk_U1094 (.A( u1_key_r_0 ) , .ZN( u1_uk_n1172 ) );
  INV_X1 u1_uk_U1095 (.A( u1_key_r_16 ) , .ZN( u1_uk_n1182 ) );
  INV_X1 u1_uk_U1096 (.A( u1_key_r_13 ) , .ZN( u1_uk_n1180 ) );
  INV_X1 u1_uk_U1097 (.A( u1_key_r_1 ) , .ZN( u1_uk_n1173 ) );
  INV_X1 u1_uk_U1098 (.A( u1_key_r_2 ) , .ZN( u1_uk_n1174 ) );
  INV_X1 u1_uk_U1099 (.A( u1_key_r_19 ) , .ZN( u1_uk_n1184 ) );
  INV_X1 u1_uk_U11 (.A( u1_uk_n298 ) , .ZN( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U110 (.ZN( u1_K14_5 ) , .B2( u1_uk_n1826 ) , .B1( u1_uk_n250 ) , .A( u1_uk_n962 ) );
  INV_X1 u1_uk_U1100 (.A( u1_key_r_4 ) , .ZN( u1_uk_n1175 ) );
  INV_X1 u1_uk_U1101 (.A( u1_key_r_17 ) , .ZN( u1_uk_n1183 ) );
  INV_X1 u1_uk_U1102 (.A( u1_key_r_53 ) , .ZN( u1_uk_n1214 ) );
  OAI21_X1 u1_uk_U1103 (.ZN( u1_K13_28 ) , .B2( u1_uk_n1783 ) , .B1( u1_uk_n230 ) , .A( u1_uk_n695 ) );
  NAND2_X1 u1_uk_U1104 (.A1( u1_uk_K_r11_21 ) , .A2( u1_uk_n277 ) , .ZN( u1_uk_n695 ) );
  OAI21_X1 u1_uk_U1105 (.ZN( u1_K8_14 ) , .A( u1_uk_n1129 ) , .B2( u1_uk_n1559 ) , .B1( u1_uk_n203 ) );
  NAND2_X1 u1_uk_U1106 (.A1( u1_uk_K_r6_34 ) , .ZN( u1_uk_n1129 ) , .A2( u1_uk_n291 ) );
  OAI21_X1 u1_uk_U1107 (.ZN( u1_K16_14 ) , .B2( u1_uk_n1235 ) , .B1( u1_uk_n252 ) , .A( u1_uk_n981 ) );
  NAND2_X1 u1_uk_U1108 (.A1( u1_uk_K_r14_18 ) , .A2( u1_uk_n291 ) , .ZN( u1_uk_n981 ) );
  OAI21_X1 u1_uk_U1109 (.ZN( u1_K3_40 ) , .A( u1_uk_n1044 ) , .B2( u1_uk_n1330 ) , .B1( u1_uk_n209 ) );
  NAND2_X1 u1_uk_U111 (.A1( u1_uk_K_r12_10 ) , .A2( u1_uk_n298 ) , .ZN( u1_uk_n962 ) );
  NAND2_X1 u1_uk_U1110 (.A1( u1_uk_K_r1_21 ) , .ZN( u1_uk_n1044 ) , .A2( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U1111 (.ZN( u1_K16_39 ) , .B2( u1_uk_n1231 ) , .B1( u1_uk_n291 ) , .A( u1_uk_n990 ) );
  NAND2_X1 u1_uk_U1112 (.A1( u1_uk_K_r14_15 ) , .A2( u1_uk_n214 ) , .ZN( u1_uk_n990 ) );
  OAI21_X1 u1_uk_U1113 (.ZN( u1_K8_39 ) , .A( u1_uk_n1139 ) , .B2( u1_uk_n1556 ) , .B1( u1_uk_n203 ) );
  NAND2_X1 u1_uk_U1114 (.A1( u1_uk_K_r6_31 ) , .ZN( u1_uk_n1139 ) , .A2( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U1115 (.ZN( u1_K5_39 ) , .A( u1_uk_n1081 ) , .B2( u1_uk_n1406 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U1116 (.A1( u1_uk_K_r3_16 ) , .ZN( u1_uk_n1081 ) , .A2( u1_uk_n242 ) );
  INV_X1 u1_uk_U1117 (.ZN( u1_K13_10 ) , .A( u1_uk_n671 ) );
  AOI22_X1 u1_uk_U1118 (.B2( u1_uk_K_r11_26 ) , .A2( u1_uk_K_r11_6 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n203 ) , .ZN( u1_uk_n671 ) );
  AOI22_X1 u1_uk_U1120 (.B2( u1_uk_K_r7_48 ) , .A2( u1_uk_K_r7_55 ) , .B1( u1_uk_n109 ) , .ZN( u1_uk_n1148 ) , .A1( u1_uk_n220 ) );
  AOI22_X1 u1_uk_U1122 (.B2( u1_uk_K_r0_34 ) , .A2( u1_uk_K_r0_55 ) , .ZN( u1_uk_n1021 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) );
  INV_X1 u1_uk_U1123 (.ZN( u1_K1_11 ) , .A( u1_uk_n997 ) );
  AOI22_X1 u1_uk_U1124 (.B2( u1_key_r_32 ) , .A2( u1_key_r_39 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n277 ) , .ZN( u1_uk_n997 ) );
  AOI22_X1 u1_uk_U1126 (.A2( u1_key_r_5 ) , .B2( u1_key_r_55 ) , .ZN( u1_uk_n1002 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n294 ) );
  AOI22_X1 u1_uk_U1128 (.B2( u1_key_r_35 ) , .A2( u1_key_r_42 ) , .ZN( u1_uk_n1015 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n298 ) );
  INV_X1 u1_uk_U1129 (.ZN( u1_K11_8 ) , .A( u1_uk_n501 ) );
  AOI22_X1 u1_uk_U113 (.B2( u1_uk_K_r11_48 ) , .A2( u1_uk_K_r11_53 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n223 ) , .ZN( u1_uk_n948 ) );
  AOI22_X1 u1_uk_U1130 (.B2( u1_uk_K_r9_12 ) , .A2( u1_uk_K_r9_18 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n501 ) );
  AOI22_X1 u1_uk_U1132 (.B2( u1_uk_K_r9_25 ) , .A2( u1_uk_K_r9_6 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n291 ) , .ZN( u1_uk_n379 ) );
  AOI22_X1 u1_uk_U1134 (.B2( u1_uk_K_r6_3 ) , .A2( u1_uk_K_r6_53 ) , .ZN( u1_uk_n1128 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) );
  AOI22_X1 u1_uk_U1136 (.B2( u1_uk_K_r0_13 ) , .A2( u1_uk_K_r0_34 ) , .ZN( u1_uk_n1034 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n27 ) );
  AOI22_X1 u1_uk_U1138 (.B2( u1_key_r_48 ) , .A2( u1_key_r_55 ) , .ZN( u1_uk_n1003 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U114 (.ZN( u1_K12_5 ) , .A2( u1_uk_n1712 ) , .B2( u1_uk_n1738 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n99 ) );
  AOI22_X1 u1_uk_U1140 (.B2( u1_uk_K_r9_1 ) , .A2( u1_uk_K_r9_9 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n421 ) );
  INV_X1 u1_uk_U1141 (.ZN( u1_K12_32 ) , .A( u1_uk_n582 ) );
  AOI22_X1 u1_uk_U1142 (.B2( u1_uk_K_r10_23 ) , .A2( u1_uk_K_r10_28 ) , .B1( u1_uk_n10 ) , .A1( u1_uk_n294 ) , .ZN( u1_uk_n582 ) );
  AOI22_X1 u1_uk_U1144 (.B2( u1_uk_K_r0_15 ) , .A2( u1_uk_K_r0_36 ) , .ZN( u1_uk_n1029 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n271 ) );
  AOI22_X1 u1_uk_U1146 (.B2( u1_uk_K_r7_32 ) , .A2( u1_uk_K_r7_39 ) , .B1( u1_uk_n11 ) , .ZN( u1_uk_n1156 ) , .A1( u1_uk_n294 ) );
  AOI22_X1 u1_uk_U1148 (.B2( u1_uk_K_r2_13 ) , .A2( u1_uk_K_r2_33 ) , .ZN( u1_uk_n1054 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U115 (.ZN( u1_K9_5 ) , .B2( u1_uk_n1610 ) , .A2( u1_uk_n1616 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n188 ) );
  AOI22_X1 u1_uk_U1150 (.B2( u1_uk_K_r5_26 ) , .A2( u1_uk_K_r5_48 ) , .ZN( u1_uk_n1106 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n217 ) );
  INV_X1 u1_uk_U1151 (.ZN( u1_K1_32 ) , .A( u1_uk_n1010 ) );
  AOI22_X1 u1_uk_U1152 (.B2( u1_key_r_22 ) , .A2( u1_key_r_29 ) , .ZN( u1_uk_n1010 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) );
  AOI22_X1 u1_uk_U1154 (.B2( u1_uk_K_r5_0 ) , .A2( u1_uk_K_r5_51 ) , .ZN( u1_uk_n1118 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n222 ) );
  AOI22_X1 u1_uk_U1156 (.B2( u1_uk_K_r4_17 ) , .A2( u1_uk_K_r4_55 ) , .ZN( u1_uk_n1096 ) , .B1( u1_uk_n257 ) , .A1( u1_uk_n27 ) );
  AOI22_X1 u1_uk_U1158 (.B2( u1_uk_K_r8_17 ) , .A2( u1_uk_K_r8_39 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n297 ) , .ZN( u1_uk_n299 ) );
  OAI22_X1 u1_uk_U116 (.ZN( u1_K7_5 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1487 ) , .A2( u1_uk_n1504 ) , .B1( u1_uk_n242 ) );
  AOI22_X1 u1_uk_U1160 (.B2( u1_uk_K_r6_10 ) , .A2( u1_uk_K_r6_17 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1130 ) , .B1( u1_uk_n207 ) );
  AOI22_X1 u1_uk_U1162 (.B2( u1_uk_K_r5_31 ) , .A2( u1_uk_K_r5_7 ) , .A1( u1_uk_n10 ) , .ZN( u1_uk_n1114 ) , .B1( u1_uk_n208 ) );
  AOI22_X1 u1_uk_U1164 (.B2( u1_uk_K_r11_34 ) , .A2( u1_uk_K_r11_54 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n252 ) , .ZN( u1_uk_n676 ) );
  AOI22_X1 u1_uk_U1165 (.B1( n116 ) , .A2( u1_uk_K_r13_2 ) , .B2( u1_uk_K_r13_23 ) , .A1( u1_uk_n286 ) , .ZN( u1_uk_n974 ) );
  AOI22_X1 u1_uk_U1167 (.B2( u1_uk_K_r11_26 ) , .A2( u1_uk_K_r11_46 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n27 ) , .ZN( u1_uk_n702 ) );
  OAI22_X1 u1_uk_U117 (.ZN( u1_K5_5 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1398 ) , .B2( u1_uk_n1422 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U118 (.ZN( u1_K2_5 ) , .B2( u1_uk_n1274 ) , .A2( u1_uk_n1277 ) , .A1( u1_uk_n291 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U119 (.ZN( u1_K10_41 ) , .A2( u1_uk_n1624 ) , .B2( u1_uk_n1652 ) , .A1( u1_uk_n223 ) , .B1( u1_uk_n31 ) );
  INV_X1 u1_uk_U12 (.A( u1_uk_n208 ) , .ZN( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U120 (.ZN( u1_K14_41 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1806 ) , .B2( u1_uk_n1811 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U121 (.ZN( u1_K12_41 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1735 ) , .A2( u1_uk_n1744 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U122 (.ZN( u1_K3_41 ) , .A2( u1_uk_n1313 ) , .B2( u1_uk_n1318 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U123 (.ZN( u1_K16_47 ) , .B2( u1_uk_n1218 ) , .A2( u1_uk_n1222 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U124 (.ZN( u1_K13_47 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1782 ) , .A2( u1_uk_n1792 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U125 (.ZN( u1_K12_47 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1709 ) , .A2( u1_uk_n1736 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U126 (.ZN( u1_K11_47 ) , .A( u1_uk_n472 ) );
  AOI22_X1 u1_uk_U127 (.B2( u1_uk_K_r9_15 ) , .A2( u1_uk_K_r9_23 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n223 ) , .ZN( u1_uk_n472 ) );
  OAI22_X1 u1_uk_U128 (.ZN( u1_K10_47 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1624 ) , .B2( u1_uk_n1639 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U129 (.ZN( u1_K8_47 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1561 ) , .A2( u1_uk_n1567 ) , .A1( u1_uk_n294 ) );
  INV_X1 u1_uk_U13 (.A( u1_uk_n222 ) , .ZN( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U130 (.ZN( u1_K7_47 ) , .A2( u1_uk_n1486 ) , .B2( u1_uk_n1500 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U131 (.ZN( u1_K6_47 ) , .A( u1_uk_n1100 ) , .B1( u1_uk_n142 ) , .B2( u1_uk_n1449 ) );
  NAND2_X1 u1_uk_U132 (.A1( u1_uk_K_r4_23 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1100 ) );
  OAI22_X1 u1_uk_U133 (.ZN( u1_K5_47 ) , .B2( u1_uk_n1395 ) , .A2( u1_uk_n1419 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U134 (.ZN( u1_K4_47 ) , .B2( u1_uk_n1380 ) , .A2( u1_uk_n1389 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U135 (.ZN( u1_K2_47 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1033 ) , .B2( u1_uk_n1271 ) );
  NAND2_X1 u1_uk_U136 (.A1( u1_uk_K_r0_52 ) , .ZN( u1_uk_n1033 ) , .A2( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U137 (.ZN( u1_K1_15 ) , .B2( u1_uk_n1191 ) , .A2( u1_uk_n1197 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U138 (.ZN( u1_K4_15 ) , .B2( u1_uk_n1358 ) , .A2( u1_uk_n1386 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U139 (.ZN( u1_K5_15 ) , .A( u1_uk_n1072 ) , .B2( u1_uk_n1409 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U14 (.ZN( u1_uk_n100 ) , .A( u1_uk_n213 ) );
  NAND2_X1 u1_uk_U140 (.A1( u1_uk_K_r3_34 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1072 ) );
  AOI22_X1 u1_uk_U142 (.B2( u1_uk_K_r11_11 ) , .A2( u1_uk_K_r11_48 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n678 ) );
  OAI22_X1 u1_uk_U143 (.ZN( u1_K7_15 ) , .A2( u1_uk_n1484 ) , .B2( u1_uk_n1524 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n92 ) );
  AOI22_X1 u1_uk_U145 (.B2( u1_uk_K_r10_25 ) , .A2( u1_uk_K_r10_34 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n252 ) , .ZN( u1_uk_n504 ) );
  OAI22_X1 u1_uk_U146 (.ZN( u1_K3_15 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1312 ) , .B2( u1_uk_n1347 ) , .A1( u1_uk_n286 ) );
  AOI22_X1 u1_uk_U148 (.B2( u1_uk_K_r11_19 ) , .A2( u1_uk_K_r11_39 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n252 ) , .ZN( u1_uk_n685 ) );
  OAI22_X1 u1_uk_U149 (.ZN( u1_K11_15 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1676 ) , .A2( u1_uk_n1691 ) , .A1( u1_uk_n297 ) );
  INV_X1 u1_uk_U15 (.A( u1_uk_n188 ) , .ZN( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U150 (.ZN( u1_K6_19 ) , .A( u1_uk_n1091 ) , .B2( u1_uk_n1444 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U151 (.A1( u1_uk_K_r4_48 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1091 ) );
  OAI21_X1 u1_uk_U152 (.ZN( u1_K2_15 ) , .A( u1_uk_n1024 ) , .B2( u1_uk_n1291 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U153 (.A1( u1_uk_K_r0_19 ) , .ZN( u1_uk_n1024 ) , .A2( u1_uk_n118 ) );
  OAI22_X1 u1_uk_U154 (.ZN( u1_K1_19 ) , .B2( u1_uk_n1175 ) , .A2( u1_uk_n1215 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U155 (.ZN( u1_K16_15 ) , .B2( u1_uk_n1236 ) , .A2( u1_uk_n1243 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U156 (.ZN( u1_K10_15 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1622 ) , .B2( u1_uk_n1659 ) , .B1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U157 (.ZN( u1_K15_15 ) , .B2( u1_uk_n1873 ) , .B1( u1_uk_n222 ) , .A( u1_uk_n967 ) );
  NAND2_X1 u1_uk_U158 (.A1( u1_uk_K_r13_19 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n967 ) );
  INV_X1 u1_uk_U159 (.ZN( u1_K14_19 ) , .A( u1_uk_n951 ) );
  INV_X1 u1_uk_U16 (.ZN( u1_uk_n109 ) , .A( u1_uk_n231 ) );
  AOI22_X1 u1_uk_U160 (.B2( u1_uk_K_r12_25 ) , .A2( u1_uk_K_r12_33 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n951 ) );
  AOI22_X1 u1_uk_U162 (.B2( u1_uk_K_r9_10 ) , .A2( u1_uk_K_r9_48 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n222 ) , .ZN( u1_uk_n386 ) );
  AOI22_X1 u1_uk_U164 (.B1( u1_uk_K_r7_13 ) , .A2( u1_uk_K_r7_20 ) , .ZN( u1_uk_n1154 ) , .A1( u1_uk_n291 ) , .B2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U165 (.ZN( u1_K7_19 ) , .B2( u1_uk_n1495 ) , .A2( u1_uk_n1505 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U166 (.ZN( u1_K4_19 ) , .B2( u1_uk_n1365 ) , .A2( u1_uk_n1377 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U167 (.ZN( u1_K3_19 ) , .A( u1_uk_n1037 ) , .B2( u1_uk_n1324 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U168 (.A1( u1_uk_K_r1_33 ) , .ZN( u1_uk_n1037 ) , .A2( u1_uk_n63 ) );
  INV_X1 u1_uk_U17 (.ZN( u1_uk_n110 ) , .A( u1_uk_n209 ) );
  AOI22_X1 u1_uk_U170 (.B2( u1_uk_K_r0_11 ) , .A2( u1_uk_K_r0_47 ) , .ZN( u1_uk_n1025 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U171 (.ZN( u1_K14_15 ) , .A1( u1_uk_n146 ) , .A2( u1_uk_n1803 ) , .B2( u1_uk_n1841 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U172 (.ZN( u1_K8_19 ) , .B2( u1_uk_n1538 ) , .A2( u1_uk_n1545 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U173 (.ZN( u1_K10_19 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1633 ) , .A2( u1_uk_n1643 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U174 (.ZN( u1_K5_30 ) , .B2( u1_uk_n1408 ) , .A2( u1_uk_n1425 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U175 (.ZN( u1_K2_30 ) , .B2( u1_uk_n1260 ) , .A2( u1_uk_n1289 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U176 (.ZN( u1_K14_30 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1811 ) , .A2( u1_uk_n1838 ) , .B1( u1_uk_n223 ) );
  INV_X1 u1_uk_U177 (.ZN( u1_K12_30 ) , .A( u1_uk_n526 ) );
  AOI22_X1 u1_uk_U178 (.B2( u1_uk_K_r10_23 ) , .A2( u1_uk_K_r10_42 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n271 ) , .ZN( u1_uk_n526 ) );
  OAI22_X1 u1_uk_U179 (.ZN( u1_K10_30 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1628 ) , .A2( u1_uk_n1656 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U18 (.ZN( u1_uk_n118 ) , .A( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U180 (.ZN( u1_K12_24 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1716 ) , .A2( u1_uk_n1745 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U181 (.ZN( u1_K1_14 ) , .A( u1_uk_n1000 ) , .B2( u1_uk_n1190 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U182 (.A1( u1_key_r_18 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1000 ) );
  INV_X1 u1_uk_U183 (.A( u1_key_r_25 ) , .ZN( u1_uk_n1190 ) );
  OAI21_X1 u1_uk_U184 (.ZN( u1_K8_30 ) , .A( u1_uk_n1136 ) , .B2( u1_uk_n1555 ) , .B1( u1_uk_n207 ) );
  NAND2_X1 u1_uk_U185 (.A1( u1_uk_K_r6_29 ) , .ZN( u1_uk_n1136 ) , .A2( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U186 (.ZN( u1_K16_30 ) , .B2( u1_uk_n1256 ) , .B1( u1_uk_n222 ) , .A( u1_uk_n987 ) );
  NAND2_X1 u1_uk_U187 (.A1( u1_uk_K_r14_45 ) , .A2( u1_uk_n279 ) , .ZN( u1_uk_n987 ) );
  OAI22_X1 u1_uk_U188 (.ZN( u1_K13_14 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1756 ) , .A2( u1_uk_n1780 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U189 (.ZN( u1_K12_14 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1718 ) , .A2( u1_uk_n1723 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U19 (.ZN( u1_uk_n141 ) , .A( u1_uk_n238 ) );
  AOI22_X1 u1_uk_U191 (.B2( u1_uk_K_r9_12 ) , .A2( u1_uk_K_r9_6 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n207 ) , .ZN( u1_uk_n382 ) );
  OAI21_X1 u1_uk_U192 (.ZN( u1_K10_24 ) , .B2( u1_uk_n1629 ) , .B1( u1_uk_n17 ) , .A( u1_uk_n319 ) );
  NAND2_X1 u1_uk_U193 (.A1( u1_uk_K_r8_40 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n319 ) );
  OAI22_X1 u1_uk_U194 (.ZN( u1_K6_14 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1440 ) , .B2( u1_uk_n1446 ) , .B1( u1_uk_n257 ) );
  AOI22_X1 u1_uk_U196 (.B2( u1_uk_K_r0_11 ) , .A2( u1_uk_K_r0_32 ) , .ZN( u1_uk_n1023 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U197 (.ZN( u1_K1_24 ) , .B2( u1_uk_n1180 ) , .A2( u1_uk_n1185 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U198 (.ZN( u1_K10_14 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1630 ) , .A2( u1_uk_n1661 ) , .B1( u1_uk_n213 ) );
  OAI21_X1 u1_uk_U199 (.ZN( u1_K13_30 ) , .B2( u1_uk_n1776 ) , .A( u1_uk_n717 ) , .B1( u1_uk_n83 ) );
  INV_X1 u1_uk_U20 (.ZN( u1_uk_n142 ) , .A( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U200 (.A1( u1_uk_K_r11_28 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n717 ) );
  OAI21_X1 u1_uk_U201 (.ZN( u1_K14_24 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1812 ) , .A( u1_uk_n952 ) );
  NAND2_X1 u1_uk_U202 (.A1( u1_uk_K_r12_41 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n952 ) );
  AOI22_X1 u1_uk_U204 (.B2( u1_uk_K_r5_18 ) , .A2( u1_uk_K_r5_40 ) , .ZN( u1_uk_n1113 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U205 (.ZN( u1_K4_24 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1352 ) , .A2( u1_uk_n1393 ) , .B1( u1_uk_n213 ) );
  AOI22_X1 u1_uk_U207 (.B2( u1_uk_K_r1_17 ) , .A2( u1_uk_K_r1_41 ) , .ZN( u1_uk_n1038 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U208 (.ZN( u1_K15_24 ) , .A1( u1_uk_n146 ) , .A2( u1_uk_n1846 ) , .B2( u1_uk_n1864 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U209 (.ZN( u1_K1_30 ) , .A( u1_uk_n1009 ) , .B2( u1_uk_n1213 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U21 (.ZN( u1_uk_n128 ) , .A( u1_uk_n297 ) );
  NAND2_X1 u1_uk_U210 (.A1( u1_key_r_45 ) , .ZN( u1_uk_n1009 ) , .A2( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U211 (.ZN( u1_K9_30 ) , .A( u1_uk_n1161 ) , .B2( u1_uk_n1600 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U212 (.A1( u1_uk_K_r7_29 ) , .ZN( u1_uk_n1161 ) , .A2( u1_uk_n187 ) );
  OAI21_X1 u1_uk_U213 (.ZN( u1_K4_30 ) , .A( u1_uk_n1062 ) , .B2( u1_uk_n1375 ) , .B1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U214 (.A1( u1_uk_K_r2_28 ) , .ZN( u1_uk_n1062 ) , .A2( u1_uk_n230 ) );
  AOI22_X1 u1_uk_U216 (.B2( u1_uk_K_r13_0 ) , .A2( u1_uk_K_r13_38 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n970 ) );
  OAI22_X1 u1_uk_U217 (.ZN( u1_K3_14 ) , .B2( u1_uk_n1340 ) , .A2( u1_uk_n1347 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n31 ) );
  AOI22_X1 u1_uk_U219 (.B2( u1_uk_K_r2_31 ) , .A2( u1_uk_K_r2_49 ) , .ZN( u1_uk_n1063 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U22 (.ZN( u1_uk_n147 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U220 (.ZN( u1_K1_31 ) , .A2( u1_uk_n1177 ) , .B2( u1_uk_n1181 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U221 (.A( u1_key_r_14 ) , .ZN( u1_uk_n1181 ) );
  OAI22_X1 u1_uk_U222 (.ZN( u1_K16_31 ) , .A2( u1_uk_n1222 ) , .B2( u1_uk_n1225 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U223 (.ZN( u1_K8_31 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1529 ) , .A2( u1_uk_n1567 ) , .B1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U224 (.ZN( u1_K12_31 ) , .B2( u1_uk_n1715 ) , .B1( u1_uk_n207 ) , .A( u1_uk_n551 ) );
  NAND2_X1 u1_uk_U225 (.A1( u1_uk_K_r10_44 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n551 ) );
  AOI22_X1 u1_uk_U227 (.B2( u1_uk_K_r9_22 ) , .A2( u1_uk_K_r9_30 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n251 ) , .ZN( u1_uk_n437 ) );
  OAI22_X1 u1_uk_U228 (.ZN( u1_K2_31 ) , .B2( u1_uk_n1260 ) , .A2( u1_uk_n1275 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n220 ) );
  INV_X1 u1_uk_U229 (.ZN( u1_K11_39 ) , .A( u1_uk_n460 ) );
  INV_X1 u1_uk_U23 (.ZN( u1_uk_n117 ) , .A( u1_uk_n277 ) );
  AOI22_X1 u1_uk_U230 (.B2( u1_uk_K_r9_30 ) , .A2( u1_uk_K_r9_7 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n292 ) , .ZN( u1_uk_n460 ) );
  INV_X1 u1_uk_U231 (.ZN( u1_K10_39 ) , .A( u1_uk_n373 ) );
  AOI22_X1 u1_uk_U232 (.B2( u1_uk_K_r8_44 ) , .A2( u1_uk_K_r8_52 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n209 ) , .ZN( u1_uk_n373 ) );
  OAI22_X1 u1_uk_U233 (.ZN( u1_K13_31 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1772 ) , .A2( u1_uk_n1790 ) , .A1( u1_uk_n207 ) );
  OAI21_X1 u1_uk_U234 (.ZN( u1_K10_31 ) , .B2( u1_uk_n1645 ) , .B1( u1_uk_n298 ) , .A( u1_uk_n342 ) );
  NAND2_X1 u1_uk_U235 (.A1( u1_uk_K_r8_16 ) , .A2( u1_uk_n277 ) , .ZN( u1_uk_n342 ) );
  OAI22_X1 u1_uk_U236 (.ZN( u1_K6_31 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1455 ) , .A2( u1_uk_n1460 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U237 (.ZN( u1_K3_31 ) , .B2( u1_uk_n1333 ) , .A2( u1_uk_n1339 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U238 (.ZN( u1_K5_31 ) , .B1( u1_uk_n100 ) , .A( u1_uk_n1077 ) , .B2( u1_uk_n1401 ) );
  NAND2_X1 u1_uk_U239 (.A1( u1_uk_K_r3_44 ) , .ZN( u1_uk_n1077 ) , .A2( u1_uk_n27 ) );
  INV_X1 u1_uk_U24 (.ZN( u1_uk_n129 ) , .A( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U240 (.ZN( u1_K15_31 ) , .B2( u1_uk_n1843 ) , .A2( u1_uk_n1860 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U241 (.ZN( u1_K1_39 ) , .A( u1_uk_n1014 ) , .B2( u1_uk_n1187 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U242 (.A1( u1_key_r_15 ) , .ZN( u1_uk_n1014 ) , .A2( u1_uk_n155 ) );
  INV_X1 u1_uk_U243 (.A( u1_key_r_22 ) , .ZN( u1_uk_n1187 ) );
  OAI22_X1 u1_uk_U244 (.ZN( u1_K14_31 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1827 ) , .A2( u1_uk_n1833 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U245 (.ZN( u1_K9_31 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1572 ) , .A2( u1_uk_n1613 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U246 (.ZN( u1_K15_39 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1848 ) , .B2( u1_uk_n1866 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U247 (.ZN( u1_K14_39 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1832 ) , .A2( u1_uk_n1836 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U248 (.ZN( u1_K13_39 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1755 ) , .A2( u1_uk_n1774 ) , .B1( u1_uk_n240 ) );
  OAI21_X1 u1_uk_U249 (.ZN( u1_K12_39 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1720 ) , .A( u1_uk_n590 ) );
  INV_X1 u1_uk_U25 (.ZN( u1_uk_n146 ) , .A( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U250 (.A1( u1_uk_K_r10_16 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n590 ) );
  OAI22_X1 u1_uk_U251 (.ZN( u1_K16_48 ) , .B2( u1_uk_n1230 ) , .A2( u1_uk_n1238 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U252 (.ZN( u1_K16_44 ) , .B2( u1_uk_n1246 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n994 ) );
  NAND2_X1 u1_uk_U253 (.A1( u1_uk_K_r14_43 ) , .A2( u1_uk_n94 ) , .ZN( u1_uk_n994 ) );
  OAI21_X1 u1_uk_U254 (.ZN( u1_K8_44 ) , .A( u1_uk_n1144 ) , .B1( u1_uk_n141 ) , .B2( u1_uk_n1568 ) );
  NAND2_X1 u1_uk_U255 (.A1( u1_uk_K_r6_0 ) , .ZN( u1_uk_n1144 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U256 (.ZN( u1_K8_48 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1534 ) , .B2( u1_uk_n1541 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U257 (.ZN( u1_K5_44 ) , .B2( u1_uk_n1419 ) , .A2( u1_uk_n1425 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U258 (.ZN( u1_K5_48 ) , .B2( u1_uk_n1407 ) , .A2( u1_uk_n1414 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U259 (.ZN( u1_K1_48 ) , .A( u1_uk_n1019 ) );
  INV_X1 u1_uk_U26 (.ZN( u1_uk_n145 ) , .A( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U260 (.B2( u1_key_r_21 ) , .A2( u1_key_r_28 ) , .ZN( u1_uk_n1019 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n291 ) );
  INV_X1 u1_uk_U261 (.ZN( u1_K1_44 ) , .A( u1_uk_n1017 ) );
  AOI22_X1 u1_uk_U262 (.B2( u1_key_r_36 ) , .A2( u1_key_r_43 ) , .ZN( u1_uk_n1017 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U263 (.ZN( u1_K15_44 ) , .B2( u1_uk_n1866 ) , .A2( u1_uk_n1884 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U264 (.ZN( u1_K15_48 ) , .B1( u1_uk_n10 ) , .B2( u1_uk_n1854 ) , .A( u1_uk_n975 ) );
  NAND2_X1 u1_uk_U265 (.A1( u1_uk_K_r13_35 ) , .A2( u1_uk_n148 ) , .ZN( u1_uk_n975 ) );
  OAI22_X1 u1_uk_U266 (.ZN( u1_K14_48 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1798 ) , .A2( u1_uk_n1836 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U267 (.ZN( u1_K13_44 ) , .B2( u1_uk_n1754 ) , .A2( u1_uk_n1769 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U268 (.ZN( u1_K13_48 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1785 ) , .A( u1_uk_n947 ) );
  NAND2_X1 u1_uk_U269 (.A1( u1_uk_K_r11_8 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n947 ) );
  INV_X1 u1_uk_U27 (.ZN( u1_uk_n148 ) , .A( u1_uk_n214 ) );
  AOI22_X1 u1_uk_U271 (.B2( u1_uk_K_r10_37 ) , .A2( u1_uk_K_r10_42 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n271 ) , .ZN( u1_uk_n608 ) );
  OAI22_X1 u1_uk_U272 (.ZN( u1_K12_48 ) , .B2( u1_uk_n1721 ) , .A2( u1_uk_n1730 ) , .B1( u1_uk_n207 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U273 (.ZN( u1_K11_44 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1683 ) , .A2( u1_uk_n1703 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U274 (.ZN( u1_K10_44 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1627 ) , .A2( u1_uk_n1647 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U275 (.ZN( u1_K10_48 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1640 ) , .A2( u1_uk_n1656 ) , .A1( u1_uk_n240 ) );
  AOI22_X1 u1_uk_U277 (.B2( u1_uk_K_r7_16 ) , .A2( u1_uk_K_r7_9 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1170 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U278 (.ZN( u1_K7_44 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1489 ) , .A2( u1_uk_n1510 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U279 (.ZN( u1_K7_48 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1501 ) , .A2( u1_uk_n1521 ) , .B1( u1_uk_n291 ) );
  INV_X1 u1_uk_U28 (.A( u1_uk_n202 ) , .ZN( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U280 (.ZN( u1_K6_44 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1458 ) , .A2( u1_uk_n1476 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U281 (.ZN( u1_K6_48 ) , .B2( u1_uk_n1463 ) , .A2( u1_uk_n1470 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U282 (.ZN( u1_K4_44 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1350 ) , .A2( u1_uk_n1367 ) , .B1( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U283 (.ZN( u1_K3_44 ) , .A( u1_uk_n1045 ) , .B2( u1_uk_n1314 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U284 (.A1( u1_uk_K_r1_15 ) , .ZN( u1_uk_n1045 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U285 (.ZN( u1_K3_48 ) , .B2( u1_uk_n1307 ) , .A2( u1_uk_n1342 ) , .A1( u1_uk_n148 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U286 (.ZN( u1_K2_44 ) , .B2( u1_uk_n1281 ) , .A2( u1_uk_n1303 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U287 (.ZN( u1_K16_6 ) , .B2( u1_uk_n1244 ) , .A2( u1_uk_n1249 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U288 (.ZN( u1_K10_6 ) , .B1( u1_uk_n129 ) , .A2( u1_uk_n1621 ) , .B2( u1_uk_n1649 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U289 (.ZN( u1_K8_6 ) , .B2( u1_uk_n1544 ) , .A2( u1_uk_n1549 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n92 ) );
  INV_X1 u1_uk_U29 (.ZN( u1_uk_n10 ) , .A( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U290 (.ZN( u1_K6_6 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1474 ) , .A2( u1_uk_n1478 ) , .A1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U291 (.ZN( u1_K6_8 ) , .A( u1_uk_n1103 ) , .B2( u1_uk_n1446 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U292 (.A1( u1_uk_K_r4_18 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1103 ) );
  OAI21_X1 u1_uk_U293 (.ZN( u1_K5_6 ) , .A( u1_uk_n1086 ) , .B2( u1_uk_n1417 ) , .B1( u1_uk_n93 ) );
  NAND2_X1 u1_uk_U294 (.A1( u1_uk_K_r3_10 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1086 ) );
  OAI21_X1 u1_uk_U295 (.ZN( u1_K4_6 ) , .A( u1_uk_n1069 ) , .B2( u1_uk_n1365 ) , .B1( u1_uk_n83 ) );
  NAND2_X1 u1_uk_U296 (.A1( u1_uk_K_r2_24 ) , .ZN( u1_uk_n1069 ) , .A2( u1_uk_n145 ) );
  OAI22_X1 u1_uk_U297 (.ZN( u1_K2_6 ) , .B2( u1_uk_n1279 ) , .A2( u1_uk_n1300 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U298 (.ZN( u1_K1_8 ) , .A1( u1_uk_n100 ) , .A2( u1_uk_n1176 ) , .B2( u1_uk_n1189 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U3 (.A( u1_uk_n191 ) , .ZN( u1_uk_n31 ) );
  INV_X1 u1_uk_U30 (.ZN( u1_uk_n17 ) , .A( u1_uk_n214 ) );
  AOI22_X1 u1_uk_U300 (.B2( u1_uk_K_r13_13 ) , .A2( u1_uk_K_r13_17 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n976 ) );
  OAI22_X1 u1_uk_U301 (.ZN( u1_K12_8 ) , .B2( u1_uk_n1731 ) , .A2( u1_uk_n1752 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U302 (.ZN( u1_K8_8 ) , .B2( u1_uk_n1558 ) , .A2( u1_uk_n1564 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n94 ) );
  AOI22_X1 u1_uk_U304 (.B2( u1_uk_K_r5_26 ) , .A2( u1_uk_K_r5_4 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1126 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U305 (.ZN( u1_K5_8 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1415 ) , .A2( u1_uk_n1437 ) , .B1( u1_uk_n277 ) );
  AOI22_X1 u1_uk_U307 (.B2( u1_uk_K_r2_41 ) , .A2( u1_uk_K_r2_46 ) , .ZN( u1_uk_n1070 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U308 (.ZN( u1_K3_8 ) , .A2( u1_uk_n1310 ) , .B2( u1_uk_n1326 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U309 (.ZN( u1_K2_8 ) , .A( u1_uk_n1035 ) , .B2( u1_uk_n1270 ) , .B1( u1_uk_n148 ) );
  INV_X1 u1_uk_U31 (.ZN( u1_uk_n11 ) , .A( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U310 (.A1( u1_uk_K_r0_17 ) , .ZN( u1_uk_n1035 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U311 (.ZN( u1_K7_26 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1500 ) , .A2( u1_uk_n1520 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U312 (.ZN( u1_K1_26 ) , .A( u1_uk_n1006 ) );
  AOI22_X1 u1_uk_U313 (.B2( u1_key_r_31 ) , .A2( u1_key_r_51 ) , .ZN( u1_uk_n1006 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U314 (.ZN( u1_K16_8 ) , .A2( u1_uk_n1221 ) , .B2( u1_uk_n1234 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n60 ) );
  AOI22_X1 u1_uk_U316 (.B2( u1_uk_K_r7_15 ) , .A2( u1_uk_K_r7_8 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1158 ) , .B1( u1_uk_n208 ) );
  AOI22_X1 u1_uk_U318 (.B2( u1_uk_K_r2_16 ) , .A2( u1_uk_K_r2_7 ) , .ZN( u1_uk_n1058 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n207 ) );
  INV_X1 u1_uk_U32 (.ZN( u1_uk_n155 ) , .A( u1_uk_n271 ) );
  AOI22_X1 u1_uk_U320 (.B2( u1_uk_K_r13_38 ) , .A2( u1_uk_K_r13_44 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n291 ) , .ZN( u1_uk_n969 ) );
  OAI21_X1 u1_uk_U321 (.ZN( u1_K6_26 ) , .A( u1_uk_n1094 ) , .B2( u1_uk_n1469 ) , .B1( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U322 (.A1( u1_uk_K_r4_35 ) , .ZN( u1_uk_n1094 ) , .A2( u1_uk_n297 ) );
  OAI21_X1 u1_uk_U323 (.ZN( u1_K11_26 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1695 ) , .A( u1_uk_n409 ) );
  NAND2_X1 u1_uk_U324 (.A1( u1_uk_K_r9_35 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n409 ) );
  OAI21_X1 u1_uk_U325 (.ZN( u1_K13_26 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1765 ) , .A( u1_uk_n694 ) );
  NAND2_X1 u1_uk_U326 (.A1( u1_uk_K_r11_7 ) , .A2( u1_uk_n31 ) , .ZN( u1_uk_n694 ) );
  OAI22_X1 u1_uk_U327 (.ZN( u1_K5_26 ) , .A2( u1_uk_n1396 ) , .B2( u1_uk_n1406 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U328 (.ZN( u1_K2_26 ) , .B2( u1_uk_n1289 ) , .A2( u1_uk_n1295 ) , .A1( u1_uk_n214 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U329 (.ZN( u1_K16_26 ) , .B2( u1_uk_n1241 ) , .A2( u1_uk_n1255 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n279 ) );
  INV_X1 u1_uk_U33 (.ZN( u1_uk_n161 ) , .A( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U330 (.ZN( u1_K14_26 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1822 ) , .A2( u1_uk_n1839 ) , .A1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U331 (.ZN( u1_K12_26 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1710 ) , .B2( u1_uk_n1720 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U332 (.ZN( u1_K10_26 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1639 ) , .A2( u1_uk_n1655 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U333 (.ZN( u1_K8_26 ) , .A1( u1_uk_n10 ) , .A2( u1_uk_n1533 ) , .B2( u1_uk_n1540 ) , .B1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U334 (.ZN( u1_K3_26 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1329 ) , .A2( u1_uk_n1345 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U335 (.ZN( u1_K5_46 ) , .B2( u1_uk_n1394 ) , .A1( u1_uk_n141 ) , .A2( u1_uk_n1431 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U336 (.ZN( u1_K15_46 ) , .A2( u1_uk_n1848 ) , .B2( u1_uk_n1875 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U337 (.ZN( u1_K13_46 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1763 ) , .A2( u1_uk_n1775 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U338 (.ZN( u1_K12_46 ) , .B2( u1_uk_n1708 ) , .A2( u1_uk_n1748 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U339 (.ZN( u1_K4_46 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1360 ) , .A2( u1_uk_n1374 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U34 (.ZN( u1_uk_n162 ) , .A( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U340 (.ZN( u1_K3_46 ) , .A( u1_uk_n1047 ) , .B2( u1_uk_n1327 ) , .B1( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U341 (.A1( u1_uk_K_r1_22 ) , .ZN( u1_uk_n1047 ) , .A2( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U342 (.ZN( u1_K2_46 ) , .A2( u1_uk_n1266 ) , .B2( u1_uk_n1293 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U343 (.ZN( u1_K1_46 ) , .A( u1_uk_n1018 ) , .B2( u1_uk_n1173 ) , .B1( u1_uk_n17 ) );
  NAND2_X1 u1_uk_U344 (.A1( u1_key_r_49 ) , .ZN( u1_uk_n1018 ) , .A2( u1_uk_n142 ) );
  OAI22_X1 u1_uk_U345 (.ZN( u1_K11_4 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1693 ) , .A2( u1_uk_n1699 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U346 (.ZN( u1_K15_4 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1850 ) , .A2( u1_uk_n1880 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U347 (.ZN( u1_K14_4 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1816 ) , .A2( u1_uk_n1824 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U348 (.ZN( u1_K7_4 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1504 ) , .A2( u1_uk_n1527 ) , .B1( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U349 (.ZN( u1_K1_4 ) , .A( u1_uk_n1020 ) , .B2( u1_uk_n1214 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U35 (.ZN( u1_uk_n187 ) , .A( u1_uk_n213 ) );
  NAND2_X1 u1_uk_U350 (.A1( u1_key_r_3 ) , .ZN( u1_uk_n1020 ) , .A2( u1_uk_n223 ) );
  AOI22_X1 u1_uk_U352 (.B2( u1_uk_K_r4_41 ) , .A2( u1_uk_K_r4_47 ) , .ZN( u1_uk_n1101 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n297 ) );
  INV_X1 u1_uk_U353 (.ZN( u1_K4_4 ) , .A( u1_uk_n1067 ) );
  AOI22_X1 u1_uk_U354 (.B2( u1_uk_K_r2_13 ) , .A2( u1_uk_K_r2_18 ) , .ZN( u1_uk_n1067 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U355 (.ZN( u1_K3_4 ) , .B2( u1_uk_n1323 ) , .A2( u1_uk_n1331 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U356 (.ZN( u1_K2_4 ) , .B2( u1_uk_n1268 ) , .A2( u1_uk_n1297 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U357 (.ZN( u1_K1_40 ) , .B2( u1_uk_n1172 ) , .A2( u1_uk_n1213 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U358 (.ZN( u1_K16_40 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1218 ) , .A2( u1_uk_n1256 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U359 (.ZN( u1_K12_4 ) , .A( u1_uk_n656 ) );
  BUF_X1 u1_uk_U36 (.Z( u1_uk_n230 ) , .A( u1_uk_n277 ) );
  AOI22_X1 u1_uk_U360 (.B2( u1_uk_K_r10_27 ) , .A2( u1_uk_K_r10_4 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n31 ) , .ZN( u1_uk_n656 ) );
  OAI22_X1 u1_uk_U361 (.ZN( u1_K10_4 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1642 ) , .A2( u1_uk_n1661 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U362 (.ZN( u1_K15_40 ) , .A2( u1_uk_n1847 ) , .B2( u1_uk_n1879 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U363 (.ZN( u1_K13_40 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1774 ) , .A2( u1_uk_n1784 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U364 (.ZN( u1_K6_40 ) , .A2( u1_uk_n1442 ) , .B2( u1_uk_n1450 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n240 ) );
  INV_X1 u1_uk_U365 (.ZN( u1_K11_46 ) , .A( u1_uk_n468 ) );
  AOI22_X1 u1_uk_U366 (.B2( u1_uk_K_r9_45 ) , .A2( u1_uk_K_r9_9 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n292 ) , .ZN( u1_uk_n468 ) );
  OAI21_X1 u1_uk_U367 (.ZN( u1_K9_46 ) , .B1( u1_uk_n11 ) , .A( u1_uk_n1169 ) , .B2( u1_uk_n1607 ) );
  NAND2_X1 u1_uk_U368 (.A1( u1_uk_K_r7_37 ) , .ZN( u1_uk_n1169 ) , .A2( u1_uk_n31 ) );
  BUF_X1 u1_uk_U37 (.Z( u1_uk_n213 ) , .A( u1_uk_n286 ) );
  AOI22_X1 u1_uk_U370 (.B2( u1_uk_K_r5_23 ) , .A2( u1_uk_K_r5_31 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1124 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U371 (.ZN( u1_K10_40 ) , .A( u1_uk_n375 ) );
  AOI22_X1 u1_uk_U372 (.A2( u1_uk_K_r8_2 ) , .B2( u1_uk_K_r8_22 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n250 ) , .ZN( u1_uk_n375 ) );
  OAI22_X1 u1_uk_U373 (.ZN( u1_K11_40 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1664 ) , .B2( u1_uk_n1672 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U374 (.ZN( u1_K8_40 ) , .B2( u1_uk_n1555 ) , .A2( u1_uk_n1561 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U375 (.ZN( u1_K7_40 ) , .A2( u1_uk_n1482 ) , .B2( u1_uk_n1494 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U376 (.ZN( u1_K4_40 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1372 ) , .A2( u1_uk_n1382 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U377 (.ZN( u1_K2_40 ) , .A2( u1_uk_n1265 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1296 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U378 (.ZN( u1_K15_33 ) , .B2( u1_uk_n1870 ) , .B1( u1_uk_n83 ) , .A( u1_uk_n972 ) );
  NAND2_X1 u1_uk_U379 (.A1( u1_uk_K_r13_31 ) , .A2( u1_uk_n60 ) , .ZN( u1_uk_n972 ) );
  BUF_X1 u1_uk_U38 (.Z( u1_uk_n208 ) , .A( u1_uk_n291 ) );
  OAI21_X1 u1_uk_U380 (.ZN( u1_K2_33 ) , .A( u1_uk_n1030 ) , .B2( u1_uk_n1288 ) , .B1( u1_uk_n223 ) );
  NAND2_X1 u1_uk_U381 (.A1( u1_uk_K_r0_31 ) , .ZN( u1_uk_n1030 ) , .A2( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U382 (.ZN( u1_K1_28 ) , .B2( u1_uk_n1173 ) , .A2( u1_uk_n1178 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U383 (.A( u1_key_r_8 ) , .ZN( u1_uk_n1178 ) );
  OAI22_X1 u1_uk_U384 (.ZN( u1_K14_28 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1821 ) , .A2( u1_uk_n1827 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U385 (.ZN( u1_K11_28 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1672 ) , .A2( u1_uk_n1704 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U386 (.ZN( u1_K6_28 ) , .B2( u1_uk_n1450 ) , .A2( u1_uk_n1477 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U387 (.ZN( u1_K3_28 ) , .B2( u1_uk_n1328 ) , .A2( u1_uk_n1333 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U388 (.ZN( u1_K5_33 ) , .A( u1_uk_n1078 ) , .B2( u1_uk_n1431 ) , .B1( u1_uk_n214 ) );
  NAND2_X1 u1_uk_U389 (.A1( u1_uk_K_r3_14 ) , .ZN( u1_uk_n1078 ) , .A2( u1_uk_n252 ) );
  BUF_X1 u1_uk_U39 (.Z( u1_uk_n202 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U390 (.ZN( u1_K15_28 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1855 ) , .A2( u1_uk_n1883 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U391 (.ZN( u1_K12_28 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1710 ) , .A2( u1_uk_n1714 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U392 (.ZN( u1_K10_28 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1640 ) , .A2( u1_uk_n1647 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U393 (.ZN( u1_K9_28 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1607 ) , .A2( u1_uk_n1614 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U394 (.ZN( u1_K7_28 ) , .B2( u1_uk_n1501 ) , .A2( u1_uk_n1510 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U395 (.ZN( u1_K5_28 ) , .B2( u1_uk_n1396 ) , .A2( u1_uk_n1400 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U396 (.ZN( u1_K14_1 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1808 ) , .A2( u1_uk_n1813 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U397 (.ZN( u1_K11_1 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1688 ) , .A2( u1_uk_n1705 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U398 (.ZN( u1_K3_1 ) , .B2( u1_uk_n1315 ) , .A2( u1_uk_n1320 ) , .A1( u1_uk_n279 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U399 (.ZN( u1_K2_1 ) , .B2( u1_uk_n1284 ) , .A2( u1_uk_n1305 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U4 (.ZN( u1_uk_n164 ) , .A( u1_uk_n203 ) );
  BUF_X1 u1_uk_U40 (.Z( u1_uk_n209 ) , .A( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U400 (.ZN( u1_K7_1 ) , .A( u1_uk_n1108 ) , .B2( u1_uk_n1492 ) , .B1( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U401 (.A1( u1_uk_K_r5_10 ) , .ZN( u1_uk_n1108 ) , .A2( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U402 (.ZN( u1_K5_1 ) , .B2( u1_uk_n1422 ) , .A2( u1_uk_n1429 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U403 (.ZN( u1_K1_9 ) , .B2( u1_uk_n1209 ) , .A2( u1_uk_n1215 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U404 (.ZN( u1_K13_16 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1761 ) , .A2( u1_uk_n1766 ) , .B1( u1_uk_n202 ) );
  OAI21_X1 u1_uk_U405 (.ZN( u1_K10_16 ) , .B2( u1_uk_n1660 ) , .B1( u1_uk_n286 ) , .A( u1_uk_n305 ) );
  NAND2_X1 u1_uk_U406 (.A1( u1_uk_K_r8_32 ) , .A2( u1_uk_n203 ) , .ZN( u1_uk_n305 ) );
  OAI22_X1 u1_uk_U407 (.ZN( u1_K9_16 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1578 ) , .A2( u1_uk_n1585 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U408 (.ZN( u1_K8_16 ) , .B2( u1_uk_n1536 ) , .A2( u1_uk_n1544 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U409 (.ZN( u1_K7_16 ) , .A( u1_uk_n1107 ) , .B2( u1_uk_n1526 ) , .B1( u1_uk_n161 ) );
  BUF_X1 u1_uk_U41 (.Z( u1_uk_n203 ) , .A( u1_uk_n291 ) );
  NAND2_X1 u1_uk_U410 (.A1( u1_uk_K_r5_32 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1107 ) );
  OAI22_X1 u1_uk_U411 (.ZN( u1_K6_16 ) , .B2( u1_uk_n1466 ) , .A2( u1_uk_n1472 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U412 (.ZN( u1_K4_16 ) , .B2( u1_uk_n1359 ) , .A2( u1_uk_n1363 ) , .B1( u1_uk_n145 ) , .A1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U413 (.ZN( u1_K3_16 ) , .A( u1_uk_n1036 ) , .B2( u1_uk_n1348 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U414 (.A1( u1_uk_K_r1_6 ) , .ZN( u1_uk_n1036 ) , .A2( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U415 (.ZN( u1_K1_16 ) , .B2( u1_uk_n1192 ) , .A2( u1_uk_n1198 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U416 (.ZN( u1_K15_9 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1873 ) , .A( u1_uk_n977 ) );
  NAND2_X1 u1_uk_U417 (.A1( u1_uk_K_r13_4 ) , .A2( u1_uk_n63 ) , .ZN( u1_uk_n977 ) );
  OAI21_X1 u1_uk_U418 (.ZN( u1_K14_9 ) , .B2( u1_uk_n1818 ) , .B1( u1_uk_n83 ) , .A( u1_uk_n963 ) );
  NAND2_X1 u1_uk_U419 (.A1( u1_uk_K_r12_18 ) , .ZN( u1_uk_n963 ) , .A2( u1_uk_n99 ) );
  BUF_X1 u1_uk_U42 (.Z( u1_uk_n242 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U420 (.ZN( u1_K13_9 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1761 ) , .A2( u1_uk_n1773 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U421 (.ZN( u1_K12_9 ) , .A1( u1_uk_n10 ) , .B2( u1_uk_n1745 ) , .A2( u1_uk_n1752 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U422 (.ZN( u1_K11_9 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1663 ) , .A2( u1_uk_n1693 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U423 (.ZN( u1_K8_9 ) , .A1( u1_uk_n109 ) , .A2( u1_uk_n1532 ) , .B2( u1_uk_n1538 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U424 (.ZN( u1_K5_9 ) , .B2( u1_uk_n1427 ) , .A2( u1_uk_n1437 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U425 (.ZN( u1_K4_9 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1359 ) , .A2( u1_uk_n1369 ) , .B1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U426 (.ZN( u1_K3_9 ) , .A( u1_uk_n1049 ) , .B2( u1_uk_n1325 ) , .B1( u1_uk_n277 ) );
  NAND2_X1 u1_uk_U427 (.A1( u1_uk_K_r1_18 ) , .ZN( u1_uk_n1049 ) , .A2( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U428 (.ZN( u1_K2_9 ) , .A2( u1_uk_n1262 ) , .B2( u1_uk_n1291 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U429 (.ZN( u1_K16_9 ) , .B2( u1_uk_n1251 ) , .A2( u1_uk_n1258 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n60 ) );
  BUF_X1 u1_uk_U43 (.Z( u1_uk_n220 ) , .A( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U430 (.ZN( u1_K12_33 ) , .B2( u1_uk_n1748 ) , .A( u1_uk_n586 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U431 (.A1( u1_uk_K_r10_14 ) , .A2( u1_uk_n117 ) , .ZN( u1_uk_n586 ) );
  OAI22_X1 u1_uk_U432 (.ZN( u1_K16_16 ) , .B2( u1_uk_n1237 ) , .A2( u1_uk_n1244 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U433 (.ZN( u1_K15_16 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1859 ) , .A2( u1_uk_n1874 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U434 (.ZN( u1_K5_16 ) , .B1( u1_uk_n129 ) , .A2( u1_uk_n1397 ) , .B2( u1_uk_n1410 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U435 (.ZN( u1_K2_16 ) , .B2( u1_uk_n1274 ) , .A2( u1_uk_n1292 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U436 (.ZN( u1_K2_28 ) , .A( u1_uk_n1028 ) );
  AOI22_X1 u1_uk_U437 (.B2( u1_uk_K_r0_15 ) , .A2( u1_uk_K_r0_49 ) , .ZN( u1_uk_n1028 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U438 (.ZN( u1_K14_37 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1815 ) , .A2( u1_uk_n1821 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U439 (.ZN( u1_K5_37 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1395 ) , .A2( u1_uk_n1433 ) , .B1( u1_uk_n257 ) );
  BUF_X1 u1_uk_U44 (.Z( u1_uk_n214 ) , .A( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U440 (.ZN( u1_K4_37 ) , .B2( u1_uk_n1361 ) , .A2( u1_uk_n1375 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n209 ) );
  AOI22_X1 u1_uk_U442 (.B2( u1_uk_K_r8_28 ) , .A2( u1_uk_K_r8_52 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n208 ) , .ZN( u1_uk_n366 ) );
  AOI22_X1 u1_uk_U444 (.B2( u1_uk_K_r6_14 ) , .A2( u1_uk_K_r6_7 ) , .ZN( u1_uk_n1138 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n203 ) );
  AOI22_X1 u1_uk_U446 (.B2( u1_uk_K_r8_17 ) , .A2( u1_uk_K_r8_27 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n297 ) , .ZN( u1_uk_n376 ) );
  AOI22_X1 u1_uk_U448 (.B2( u1_uk_K_r7_13 ) , .A1( u1_uk_K_r7_6 ) , .ZN( u1_uk_n1171 ) , .A2( u1_uk_n148 ) , .B1( u1_uk_n207 ) );
  BUF_X1 u1_uk_U45 (.Z( u1_uk_n240 ) , .A( u1_uk_n271 ) );
  AOI22_X1 u1_uk_U450 (.B2( u1_uk_K_r4_3 ) , .A2( u1_uk_K_r4_41 ) , .ZN( u1_uk_n1104 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U451 (.ZN( u1_K7_9 ) , .B2( u1_uk_n1491 ) , .A2( u1_uk_n1498 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U452 (.ZN( u1_K15_1 ) , .B2( u1_uk_n1868 ) , .A2( u1_uk_n1887 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n99 ) );
  AOI22_X1 u1_uk_U454 (.B2( u1_uk_K_r14_2 ) , .A2( u1_uk_K_r14_50 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n989 ) );
  OAI22_X1 u1_uk_U455 (.ZN( u1_K16_33 ) , .B2( u1_uk_n1250 ) , .A2( u1_uk_n1255 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U456 (.ZN( u1_K14_33 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1815 ) , .A2( u1_uk_n1833 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U457 (.ZN( u1_K13_33 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1753 ) , .A2( u1_uk_n1758 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U458 (.ZN( u1_K11_33 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1683 ) , .A2( u1_uk_n1689 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U459 (.ZN( u1_K7_33 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1494 ) , .A2( u1_uk_n1514 ) , .B1( u1_uk_n279 ) );
  BUF_X1 u1_uk_U46 (.Z( u1_uk_n238 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U460 (.ZN( u1_K3_33 ) , .B2( u1_uk_n1322 ) , .A2( u1_uk_n1339 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n203 ) );
  INV_X1 u1_uk_U461 (.ZN( u1_K9_33 ) , .A( u1_uk_n1162 ) );
  AOI22_X1 u1_uk_U462 (.B2( u1_uk_K_r7_1 ) , .A2( u1_uk_K_r7_8 ) , .ZN( u1_uk_n1162 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n286 ) );
  AOI22_X1 u1_uk_U464 (.B2( u1_uk_K_r8_22 ) , .A2( u1_uk_K_r8_42 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n297 ) , .ZN( u1_uk_n349 ) );
  INV_X1 u1_uk_U465 (.ZN( u1_K1_33 ) , .A( u1_uk_n1011 ) );
  AOI22_X1 u1_uk_U466 (.B2( u1_key_r_44 ) , .A2( u1_key_r_51 ) , .ZN( u1_uk_n1011 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U467 (.ZN( u1_K8_33 ) , .B2( u1_uk_n1528 ) , .A2( u1_uk_n1533 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U468 (.ZN( u1_K6_33 ) , .B2( u1_uk_n1458 ) , .A2( u1_uk_n1463 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U469 (.ZN( u1_K4_33 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1349 ) , .A2( u1_uk_n1356 ) , .A1( u1_uk_n250 ) );
  BUF_X1 u1_uk_U47 (.Z( u1_uk_n217 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U470 (.ZN( u1_K15_37 ) , .A2( u1_uk_n1849 ) , .B2( u1_uk_n1876 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U471 (.ZN( u1_K13_37 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1764 ) , .A2( u1_uk_n1776 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U472 (.ZN( u1_K12_37 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1709 ) , .A2( u1_uk_n1749 ) , .A1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U473 (.ZN( u1_K11_37 ) , .B2( u1_uk_n1694 ) , .A( u1_uk_n456 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U474 (.A1( u1_uk_K_r9_38 ) , .ZN( u1_uk_n456 ) , .A2( u1_uk_n63 ) );
  OAI21_X1 u1_uk_U475 (.ZN( u1_K9_37 ) , .A( u1_uk_n1164 ) , .B2( u1_uk_n1581 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U476 (.A1( u1_uk_K_r7_7 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n1164 ) );
  OAI21_X1 u1_uk_U477 (.ZN( u1_K6_37 ) , .A( u1_uk_n1098 ) , .B2( u1_uk_n1468 ) , .B1( u1_uk_n271 ) );
  NAND2_X1 u1_uk_U478 (.A1( u1_uk_K_r4_38 ) , .ZN( u1_uk_n1098 ) , .A2( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U479 (.ZN( u1_K3_37 ) , .B2( u1_uk_n1322 ) , .A2( u1_uk_n1328 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n94 ) );
  BUF_X1 u1_uk_U48 (.Z( u1_uk_n223 ) , .A( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U480 (.ZN( u1_K1_29 ) , .B2( u1_uk_n1182 ) , .A2( u1_uk_n1188 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U481 (.ZN( u1_K10_36 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1619 ) , .A( u1_uk_n363 ) );
  NAND2_X1 u1_uk_U482 (.A1( u1_uk_K_r8_21 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n363 ) );
  OAI21_X1 u1_uk_U483 (.ZN( u1_K14_29 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1837 ) , .A( u1_uk_n954 ) );
  NAND2_X1 u1_uk_U484 (.A1( u1_uk_K_r12_44 ) , .A2( u1_uk_n164 ) , .ZN( u1_uk_n954 ) );
  OAI22_X1 u1_uk_U485 (.ZN( u1_K13_29 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1772 ) , .A2( u1_uk_n1775 ) , .B1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U486 (.ZN( u1_K11_29 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1664 ) , .A( u1_uk_n415 ) );
  NAND2_X1 u1_uk_U487 (.A1( u1_uk_K_r9_0 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n415 ) );
  OAI21_X1 u1_uk_U488 (.ZN( u1_K3_29 ) , .A( u1_uk_n1040 ) , .B2( u1_uk_n1343 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U489 (.A1( u1_uk_K_r1_44 ) , .ZN( u1_uk_n1040 ) , .A2( u1_uk_n294 ) );
  BUF_X1 u1_uk_U49 (.Z( u1_uk_n231 ) , .A( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U490 (.ZN( u1_K2_29 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1267 ) , .B2( u1_uk_n1282 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U491 (.ZN( u1_K15_29 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1849 ) , .B2( u1_uk_n1867 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U492 (.ZN( u1_K10_29 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1627 ) , .A2( u1_uk_n1655 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U493 (.ZN( u1_K9_29 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1595 ) , .A2( u1_uk_n1599 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U494 (.ZN( u1_K5_29 ) , .B2( u1_uk_n1407 ) , .A1( u1_uk_n142 ) , .A2( u1_uk_n1426 ) , .B1( u1_uk_n277 ) );
  AOI22_X1 u1_uk_U496 (.B2( u1_uk_K_r14_16 ) , .A2( u1_uk_K_r14_23 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n277 ) , .ZN( u1_uk_n985 ) );
  AOI22_X1 u1_uk_U498 (.B2( u1_uk_K_r6_28 ) , .A2( u1_uk_K_r6_35 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1134 ) , .B1( u1_uk_n230 ) );
  OAI21_X1 u1_uk_U499 (.ZN( u1_K6_29 ) , .A( u1_uk_n1095 ) , .B2( u1_uk_n1442 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U5 (.ZN( u1_uk_n163 ) , .A( u1_uk_n202 ) );
  BUF_X1 u1_uk_U50 (.Z( u1_uk_n191 ) , .A( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U500 (.A1( u1_uk_K_r4_0 ) , .ZN( u1_uk_n1095 ) , .A2( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U502 (.B2( u1_uk_K_r2_31 ) , .A2( u1_uk_K_r2_36 ) , .ZN( u1_uk_n1060 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U503 (.ZN( u1_K12_29 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1721 ) , .A2( u1_uk_n1744 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U504 (.ZN( u1_K7_29 ) , .B2( u1_uk_n1489 ) , .A2( u1_uk_n1520 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U505 (.ZN( u1_K14_2 ) , .A1( u1_uk_n182 ) , .B2( u1_uk_n1824 ) , .A2( u1_uk_n1831 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U506 (.ZN( u1_K11_2 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1673 ) , .A2( u1_uk_n1707 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U507 (.ZN( u1_K3_2 ) , .B2( u1_uk_n1331 ) , .A2( u1_uk_n1336 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U508 (.ZN( u1_K2_2 ) , .B2( u1_uk_n1273 ) , .A2( u1_uk_n1305 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U509 (.ZN( u1_K8_2 ) , .A( u1_uk_n1135 ) , .B2( u1_uk_n1545 ) , .B1( u1_uk_n155 ) );
  BUF_X1 u1_uk_U51 (.Z( u1_uk_n207 ) , .A( u1_uk_n291 ) );
  NAND2_X1 u1_uk_U510 (.A1( u1_uk_K_r6_27 ) , .ZN( u1_uk_n1135 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U511 (.ZN( u1_K7_2 ) , .A( u1_uk_n1116 ) , .B2( u1_uk_n1484 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U512 (.A1( u1_uk_K_r5_41 ) , .ZN( u1_uk_n1116 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U513 (.ZN( u1_K5_2 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1397 ) , .B2( u1_uk_n1402 ) , .B1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U514 (.ZN( u1_K9_12 ) , .A( u1_uk_n1149 ) , .B2( u1_uk_n1573 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U515 (.A1( u1_uk_K_r7_53 ) , .ZN( u1_uk_n1149 ) , .A2( u1_uk_n142 ) );
  OAI21_X1 u1_uk_U516 (.ZN( u1_K1_12 ) , .B2( u1_uk_n1184 ) , .B1( u1_uk_n148 ) , .A( u1_uk_n998 ) );
  NAND2_X1 u1_uk_U517 (.A1( u1_key_r_12 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n998 ) );
  OAI21_X1 u1_uk_U518 (.ZN( u1_K13_17 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1773 ) , .A( u1_uk_n681 ) );
  NAND2_X1 u1_uk_U519 (.A1( u1_uk_K_r11_27 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n681 ) );
  BUF_X1 u1_uk_U52 (.Z( u1_uk_n222 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U520 (.ZN( u1_K10_17 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1626 ) , .A2( u1_uk_n1654 ) , .B1( u1_uk_n251 ) );
  OAI21_X1 u1_uk_U521 (.ZN( u1_K9_17 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1152 ) , .B2( u1_uk_n1598 ) );
  NAND2_X1 u1_uk_U522 (.A1( u1_uk_K_r7_26 ) , .ZN( u1_uk_n1152 ) , .A2( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U523 (.ZN( u1_K8_17 ) , .A( u1_uk_n1131 ) , .B2( u1_uk_n1552 ) , .B1( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U524 (.A1( u1_uk_K_r6_26 ) , .ZN( u1_uk_n1131 ) , .A2( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U525 (.ZN( u1_K7_17 ) , .B2( u1_uk_n1488 ) , .A2( u1_uk_n1518 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U526 (.ZN( u1_K4_17 ) , .A( u1_uk_n1051 ) , .B2( u1_uk_n1369 ) , .B1( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U527 (.A1( u1_uk_K_r2_27 ) , .ZN( u1_uk_n1051 ) , .A2( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U528 (.ZN( u1_K3_17 ) , .B2( u1_uk_n1317 ) , .A2( u1_uk_n1340 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U529 (.ZN( u1_K15_12 ) , .A1( u1_uk_n147 ) , .A2( u1_uk_n1845 ) , .B2( u1_uk_n1863 ) , .B1( u1_uk_n240 ) );
  BUF_X1 u1_uk_U53 (.Z( u1_uk_n188 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U530 (.ZN( u1_K14_12 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1831 ) , .A2( u1_uk_n1835 ) , .B1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U531 (.ZN( u1_K12_12 ) , .B2( u1_uk_n1719 ) , .A( u1_uk_n503 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U532 (.A1( u1_uk_K_r10_11 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n503 ) );
  OAI22_X1 u1_uk_U533 (.ZN( u1_K15_2 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1858 ) , .A2( u1_uk_n1887 ) , .B1( u1_uk_n213 ) );
  AOI22_X1 u1_uk_U535 (.B2( u1_uk_K_r10_18 ) , .A2( u1_uk_K_r10_41 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n257 ) , .ZN( u1_uk_n509 ) );
  AOI22_X1 u1_uk_U537 (.B2( u1_uk_K_r9_4 ) , .A2( u1_uk_K_r9_55 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n188 ) , .ZN( u1_uk_n385 ) );
  AOI22_X1 u1_uk_U539 (.B2( u1_uk_K_r5_17 ) , .A2( u1_uk_K_r5_39 ) , .ZN( u1_uk_n1105 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n242 ) );
  BUF_X1 u1_uk_U54 (.Z( u1_uk_n250 ) , .A( u1_uk_n257 ) );
  OAI21_X1 u1_uk_U540 (.ZN( u1_K5_12 ) , .A( u1_uk_n1071 ) , .B2( u1_uk_n1405 ) , .B1( u1_uk_n230 ) );
  NAND2_X1 u1_uk_U541 (.A1( u1_uk_K_r3_11 ) , .ZN( u1_uk_n1071 ) , .A2( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U542 (.ZN( u1_K4_12 ) , .B2( u1_uk_n1371 ) , .A2( u1_uk_n1391 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U543 (.ZN( u1_K3_12 ) , .B2( u1_uk_n1336 ) , .A2( u1_uk_n1341 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U544 (.ZN( u1_K2_12 ) , .A2( u1_uk_n1263 ) , .B2( u1_uk_n1278 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U545 (.ZN( u1_K1_36 ) , .B2( u1_uk_n1188 ) , .A2( u1_uk_n1195 ) , .A1( u1_uk_n148 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U546 (.ZN( u1_K16_12 ) , .B2( u1_uk_n1228 ) , .B1( u1_uk_n223 ) , .A( u1_uk_n979 ) );
  NAND2_X1 u1_uk_U547 (.A1( u1_uk_K_r14_12 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n979 ) );
  OAI21_X1 u1_uk_U548 (.ZN( u1_K16_17 ) , .B2( u1_uk_n1227 ) , .B1( u1_uk_n202 ) , .A( u1_uk_n982 ) );
  NAND2_X1 u1_uk_U549 (.A1( u1_uk_K_r14_10 ) , .A2( u1_uk_n257 ) , .ZN( u1_uk_n982 ) );
  BUF_X1 u1_uk_U55 (.Z( u1_uk_n251 ) , .A( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U550 (.ZN( u1_K9_36 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1599 ) , .A2( u1_uk_n1605 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U551 (.ZN( u1_K15_17 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1844 ) , .B2( u1_uk_n1862 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U552 (.ZN( u1_K14_17 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1810 ) , .A2( u1_uk_n1834 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U553 (.ZN( u1_K5_17 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1404 ) , .A2( u1_uk_n1424 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U554 (.ZN( u1_K6_17 ) , .A( u1_uk_n1089 ) );
  AOI22_X1 u1_uk_U555 (.B2( u1_uk_K_r4_4 ) , .A2( u1_uk_K_r4_55 ) , .ZN( u1_uk_n1089 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U556 (.ZN( u1_K15_36 ) , .B2( u1_uk_n1856 ) , .A2( u1_uk_n1870 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U557 (.ZN( u1_K14_36 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1800 ) , .A2( u1_uk_n1838 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U558 (.ZN( u1_K13_36 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1777 ) , .A2( u1_uk_n1783 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U559 (.ZN( u1_K3_36 ) , .B2( u1_uk_n1309 ) , .A2( u1_uk_n1344 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n203 ) );
  BUF_X1 u1_uk_U56 (.A( u1_uk_n251 ) , .Z( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U560 (.ZN( u1_K2_36 ) , .B2( u1_uk_n1272 ) , .A2( u1_uk_n1288 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U561 (.ZN( u1_K1_38 ) , .B2( u1_uk_n1195 ) , .A2( u1_uk_n1201 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U562 (.ZN( u1_K16_36 ) , .B2( u1_uk_n1233 ) , .A2( u1_uk_n1240 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U563 (.ZN( u1_K12_38 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1708 ) , .A2( u1_uk_n1735 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U564 (.ZN( u1_K11_38 ) , .B2( u1_uk_n1670 ) , .A2( u1_uk_n1678 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U565 (.ZN( u1_K9_38 ) , .B2( u1_uk_n1605 ) , .A2( u1_uk_n1612 ) , .B1( u1_uk_n214 ) , .A1( u1_uk_n92 ) );
  AOI22_X1 u1_uk_U567 (.B2( u1_uk_K_r5_1 ) , .A2( u1_uk_K_r5_21 ) , .ZN( u1_uk_n1121 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n220 ) );
  AOI22_X1 u1_uk_U569 (.B2( u1_uk_K_r9_15 ) , .A2( u1_uk_K_r9_7 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n202 ) , .ZN( u1_uk_n454 ) );
  BUF_X1 u1_uk_U57 (.Z( u1_uk_n286 ) , .A( u1_uk_n294 ) );
  AOI22_X1 u1_uk_U571 (.B2( u1_uk_K_r3_29 ) , .A2( u1_uk_K_r3_52 ) , .ZN( u1_uk_n1080 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n257 ) );
  AOI22_X1 u1_uk_U573 (.B2( u1_uk_K_r13_23 ) , .A2( u1_uk_K_r13_44 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n220 ) , .ZN( u1_uk_n973 ) );
  AOI22_X1 u1_uk_U575 (.B2( u1_uk_K_r8_28 ) , .A2( u1_uk_K_r8_8 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n369 ) );
  OAI22_X1 u1_uk_U576 (.ZN( u1_K8_36 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1554 ) , .A2( u1_uk_n1560 ) , .A1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U577 (.ZN( u1_K6_38 ) , .B2( u1_uk_n1448 ) , .B1( u1_uk_n145 ) , .A2( u1_uk_n1455 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U578 (.ZN( u1_K5_38 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1394 ) , .A2( u1_uk_n1418 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U579 (.ZN( u1_K16_10 ) , .B2( u1_uk_n1249 ) , .A2( u1_uk_n1252 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n83 ) );
  BUF_X1 u1_uk_U58 (.Z( u1_uk_n291 ) , .A( u1_uk_n294 ) );
  OAI21_X1 u1_uk_U580 (.ZN( u1_K15_10 ) , .B2( u1_uk_n1869 ) , .B1( u1_uk_n94 ) , .A( u1_uk_n964 ) );
  NAND2_X1 u1_uk_U581 (.A1( u1_uk_K_r13_55 ) , .A2( u1_uk_n92 ) , .ZN( u1_uk_n964 ) );
  OAI22_X1 u1_uk_U582 (.ZN( u1_K14_10 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1809 ) , .A2( u1_uk_n1814 ) , .B1( u1_uk_n213 ) );
  OAI21_X1 u1_uk_U583 (.ZN( u1_K11_10 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1663 ) , .A( u1_uk_n377 ) );
  NAND2_X1 u1_uk_U584 (.A1( u1_uk_K_r9_54 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n377 ) );
  OAI22_X1 u1_uk_U585 (.ZN( u1_K10_10 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1625 ) , .A2( u1_uk_n1653 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U586 (.ZN( u1_K5_10 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1403 ) , .A2( u1_uk_n1423 ) , .B1( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U588 (.B1( n116 ) , .B2( u1_uk_K_r7_25 ) , .A2( u1_uk_K_r7_32 ) , .ZN( u1_uk_n1147 ) , .A1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U589 (.ZN( u1_K8_10 ) , .B2( u1_uk_n1549 ) , .A2( u1_uk_n1551 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n92 ) );
  BUF_X1 u1_uk_U59 (.Z( u1_uk_n279 ) , .A( u1_uk_n297 ) );
  AOI22_X1 u1_uk_U591 (.B2( u1_uk_K_r4_3 ) , .A2( u1_uk_K_r4_54 ) , .ZN( u1_uk_n1088 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n208 ) );
  AOI22_X1 u1_uk_U593 (.B2( u1_uk_K_r2_26 ) , .A2( u1_uk_K_r2_6 ) , .ZN( u1_uk_n1050 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U594 (.ZN( u1_K1_10 ) , .A( u1_uk_n996 ) );
  AOI22_X1 u1_uk_U595 (.B2( u1_key_r_41 ) , .A2( u1_key_r_48 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n298 ) , .ZN( u1_uk_n996 ) );
  OAI22_X1 u1_uk_U596 (.ZN( u1_K16_22 ) , .B2( u1_uk_n1235 ) , .A2( u1_uk_n1242 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U597 (.ZN( u1_K12_22 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1722 ) , .A2( u1_uk_n1732 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U598 (.ZN( u1_K3_22 ) , .B2( u1_uk_n1311 ) , .A2( u1_uk_n1346 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U599 (.ZN( u1_K13_22 ) , .A( u1_uk_n692 ) );
  INV_X1 u1_uk_U6 (.ZN( u1_uk_n182 ) , .A( u1_uk_n223 ) );
  BUF_X1 u1_uk_U60 (.Z( u1_uk_n271 ) , .A( u1_uk_n297 ) );
  AOI22_X1 u1_uk_U600 (.B2( u1_uk_K_r11_10 ) , .A2( u1_uk_K_r11_47 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n238 ) , .ZN( u1_uk_n692 ) );
  AOI22_X1 u1_uk_U602 (.B2( u1_uk_K_r9_13 ) , .A2( u1_uk_K_r9_19 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n230 ) , .ZN( u1_uk_n407 ) );
  AOI22_X1 u1_uk_U604 (.B2( u1_uk_K_r8_27 ) , .A2( u1_uk_K_r8_5 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n279 ) , .ZN( u1_uk_n312 ) );
  AOI22_X1 u1_uk_U606 (.B2( u1_uk_K_r7_41 ) , .A2( u1_uk_K_r7_48 ) , .ZN( u1_uk_n1157 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U607 (.ZN( u1_K8_22 ) , .B2( u1_uk_n1559 ) , .A2( u1_uk_n1565 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n60 ) );
  AOI22_X1 u1_uk_U609 (.B2( u1_uk_K_r3_24 ) , .A2( u1_uk_K_r3_33 ) , .ZN( u1_uk_n1074 ) , .B1( u1_uk_n222 ) , .A1( u1_uk_n31 ) );
  BUF_X1 u1_uk_U61 (.Z( u1_uk_n277 ) , .A( u1_uk_n297 ) );
  INV_X1 u1_uk_U610 (.ZN( u1_K1_22 ) , .A( u1_uk_n1004 ) );
  AOI22_X1 u1_uk_U611 (.B2( u1_key_r_25 ) , .A2( u1_key_r_32 ) , .ZN( u1_uk_n1004 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U612 (.ZN( u1_K16_35 ) , .B2( u1_uk_n1238 ) , .A2( u1_uk_n1245 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U613 (.ZN( u1_K11_35 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1695 ) , .A2( u1_uk_n1703 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U614 (.ZN( u1_K8_35 ) , .B2( u1_uk_n1541 ) , .A2( u1_uk_n1547 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U615 (.ZN( u1_K7_35 ) , .A( u1_uk_n1120 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1482 ) );
  NAND2_X1 u1_uk_U616 (.A1( u1_uk_K_r5_37 ) , .ZN( u1_uk_n1120 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U617 (.ZN( u1_K15_35 ) , .B2( u1_uk_n1860 ) , .A2( u1_uk_n1875 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U618 (.ZN( u1_K13_35 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1764 ) , .A2( u1_uk_n1793 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U619 (.ZN( u1_K12_35 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1728 ) , .A2( u1_uk_n1737 ) , .B1( u1_uk_n213 ) );
  BUF_X1 u1_uk_U62 (.Z( u1_uk_n292 ) , .A( u1_uk_n294 ) );
  INV_X1 u1_uk_U620 (.ZN( u1_K14_35 ) , .A( u1_uk_n956 ) );
  AOI22_X1 u1_uk_U621 (.B2( u1_uk_K_r12_1 ) , .A2( u1_uk_K_r12_7 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n242 ) , .ZN( u1_uk_n956 ) );
  AOI22_X1 u1_uk_U623 (.B2( u1_uk_K_r8_2 ) , .A2( u1_uk_K_r8_37 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n252 ) , .ZN( u1_uk_n353 ) );
  AOI22_X1 u1_uk_U625 (.B2( u1_uk_K_r7_16 ) , .A2( u1_uk_K_r7_23 ) , .ZN( u1_uk_n1163 ) , .B1( u1_uk_n129 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U626 (.ZN( u1_K6_35 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1469 ) , .A2( u1_uk_n1476 ) , .A1( u1_uk_n203 ) );
  AOI22_X1 u1_uk_U628 (.B2( u1_uk_K_r3_29 ) , .A2( u1_uk_K_r3_38 ) , .ZN( u1_uk_n1079 ) , .B1( u1_uk_n251 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U629 (.ZN( u1_K4_35 ) , .B2( u1_uk_n1361 ) , .A2( u1_uk_n1390 ) , .B1( u1_uk_n142 ) , .A1( u1_uk_n271 ) );
  BUF_X1 u1_uk_U63 (.Z( u1_uk_n257 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U630 (.ZN( u1_K2_35 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1275 ) , .A2( u1_uk_n1293 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U631 (.ZN( u1_K1_35 ) , .A( u1_uk_n1012 ) );
  AOI22_X1 u1_uk_U632 (.B2( u1_key_r_28 ) , .A2( u1_key_r_35 ) , .ZN( u1_uk_n1012 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U633 (.ZN( u1_K16_11 ) , .B2( u1_uk_n1242 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n978 ) );
  NAND2_X1 u1_uk_U634 (.A1( u1_uk_K_r14_39 ) , .A2( u1_uk_n94 ) , .ZN( u1_uk_n978 ) );
  OAI21_X1 u1_uk_U635 (.ZN( u1_K15_11 ) , .B2( u1_uk_n1880 ) , .B1( u1_uk_n250 ) , .A( u1_uk_n965 ) );
  NAND2_X1 u1_uk_U636 (.A1( u1_uk_K_r13_25 ) , .A2( u1_uk_n230 ) , .ZN( u1_uk_n965 ) );
  OAI22_X1 u1_uk_U637 (.ZN( u1_K14_11 ) , .A2( u1_uk_n1801 ) , .B2( u1_uk_n1808 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U638 (.ZN( u1_K11_11 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1676 ) , .A2( u1_uk_n1682 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U639 (.ZN( u1_K3_11 ) , .A2( u1_uk_n1310 ) , .B2( u1_uk_n1315 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n191 ) );
  BUF_X1 u1_uk_U64 (.Z( u1_uk_n294 ) , .A( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U640 (.ZN( u1_K2_11 ) , .A( u1_uk_n1022 ) , .B2( u1_uk_n1297 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U641 (.A1( u1_uk_K_r0_25 ) , .ZN( u1_uk_n1022 ) , .A2( u1_uk_n141 ) );
  AOI22_X1 u1_uk_U643 (.B2( u1_uk_K_r11_17 ) , .A2( u1_uk_K_r11_54 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n191 ) , .ZN( u1_uk_n672 ) );
  OAI22_X1 u1_uk_U644 (.ZN( u1_K10_11 ) , .B2( u1_uk_n1626 ) , .A2( u1_uk_n1643 ) , .A1( u1_uk_n214 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U645 (.ZN( u1_K8_11 ) , .A( u1_uk_n1127 ) , .B2( u1_uk_n1565 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U646 (.A1( u1_uk_K_r6_55 ) , .ZN( u1_uk_n1127 ) , .A2( u1_uk_n147 ) );
  OAI22_X1 u1_uk_U647 (.ZN( u1_K7_11 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1488 ) , .A2( u1_uk_n1505 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U648 (.ZN( u1_K6_11 ) , .B2( u1_uk_n1453 ) , .A2( u1_uk_n1457 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U649 (.ZN( u1_K5_11 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1399 ) , .B2( u1_uk_n1423 ) , .B1( u1_uk_n220 ) );
  BUF_X1 u1_uk_U65 (.Z( u1_uk_n297 ) , .A( u1_uk_n298 ) );
  AOI22_X1 u1_uk_U651 (.B2( u1_uk_K_r2_18 ) , .A2( u1_uk_K_r2_55 ) , .ZN( u1_uk_n1056 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U652 (.ZN( u1_K16_45 ) , .B2( u1_uk_n1247 ) , .A2( u1_uk_n1250 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U653 (.ZN( u1_K1_45 ) , .B2( u1_uk_n1201 ) , .A2( u1_uk_n1208 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n242 ) );
  INV_X1 u1_uk_U654 (.A( u1_key_r_44 ) , .ZN( u1_uk_n1208 ) );
  OAI22_X1 u1_uk_U655 (.ZN( u1_K14_43 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1829 ) , .A2( u1_uk_n1832 ) , .B1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U656 (.ZN( u1_K4_43 ) , .A( u1_uk_n1066 ) , .B2( u1_uk_n1389 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U657 (.A1( u1_uk_K_r2_29 ) , .ZN( u1_uk_n1066 ) , .A2( u1_uk_n128 ) );
  OAI22_X1 u1_uk_U658 (.ZN( u1_K3_43 ) , .B2( u1_uk_n1334 ) , .A2( u1_uk_n1338 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U659 (.ZN( u1_K2_43 ) , .A( u1_uk_n1032 ) , .B2( u1_uk_n1276 ) , .B1( u1_uk_n162 ) );
  INV_X1 u1_uk_U66 (.A( n116 ) , .ZN( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U660 (.A1( u1_uk_K_r0_2 ) , .ZN( u1_uk_n1032 ) , .A2( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U661 (.ZN( u1_K11_3 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1669 ) , .A2( u1_uk_n1687 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U662 (.ZN( u1_K1_7 ) , .B2( u1_uk_n1185 ) , .A2( u1_uk_n1192 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U663 (.ZN( u1_K4_7 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1353 ) , .B2( u1_uk_n1357 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U664 (.ZN( u1_K9_25 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1608 ) , .A2( u1_uk_n1615 ) , .B1( u1_uk_n292 ) );
  AOI22_X1 u1_uk_U666 (.B2( u1_uk_K_r14_16 ) , .A2( u1_uk_K_r14_9 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) , .ZN( u1_uk_n993 ) );
  AOI22_X1 u1_uk_U668 (.B2( u1_uk_K_r3_15 ) , .A2( u1_uk_K_r3_38 ) , .ZN( u1_uk_n1083 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U669 (.ZN( u1_K14_45 ) , .B2( u1_uk_n1830 ) , .B1( u1_uk_n251 ) , .A( u1_uk_n960 ) );
  NAND2_X1 u1_uk_U670 (.A1( u1_uk_K_r12_16 ) , .A2( u1_uk_n292 ) , .ZN( u1_uk_n960 ) );
  OAI21_X1 u1_uk_U671 (.ZN( u1_K13_43 ) , .B2( u1_uk_n1792 ) , .B1( u1_uk_n191 ) , .A( u1_uk_n946 ) );
  NAND2_X1 u1_uk_U672 (.A1( u1_uk_K_r11_29 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n946 ) );
  OAI21_X1 u1_uk_U673 (.ZN( u1_K12_45 ) , .B2( u1_uk_n1714 ) , .B1( u1_uk_n191 ) , .A( u1_uk_n634 ) );
  NAND2_X1 u1_uk_U674 (.A1( u1_uk_K_r10_43 ) , .A2( u1_uk_n214 ) , .ZN( u1_uk_n634 ) );
  OAI22_X1 u1_uk_U675 (.ZN( u1_K11_43 ) , .B1( u1_uk_n146 ) , .B2( u1_uk_n1662 ) , .A2( u1_uk_n1704 ) , .A1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U676 (.ZN( u1_K10_43 ) , .A2( u1_uk_n1623 ) , .B2( u1_uk_n1651 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U677 (.ZN( u1_K10_45 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1628 ) , .A2( u1_uk_n1644 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U678 (.ZN( u1_K9_43 ) , .A1( u1_uk_n11 ) , .B2( u1_uk_n1588 ) , .A2( u1_uk_n1595 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U679 (.ZN( u1_K9_45 ) , .B2( u1_uk_n1571 ) , .A2( u1_uk_n1612 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U68 (.A1( n116 ) , .B2( u1_uk_K_r14_2 ) , .A2( u1_uk_K_r14_9 ) , .B1( u1_uk_n213 ) , .ZN( u1_uk_n988 ) );
  OAI22_X1 u1_uk_U680 (.ZN( u1_K7_43 ) , .A1( u1_uk_n141 ) , .A2( u1_uk_n1485 ) , .B2( u1_uk_n1514 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U681 (.ZN( u1_K10_7 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1634 ) , .A2( u1_uk_n1654 ) , .A1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U682 (.ZN( u1_K6_7 ) , .A( u1_uk_n1102 ) , .B2( u1_uk_n1465 ) , .B1( u1_uk_n222 ) );
  NAND2_X1 u1_uk_U683 (.A1( u1_uk_K_r4_33 ) , .ZN( u1_uk_n1102 ) , .A2( u1_uk_n208 ) );
  OAI21_X1 u1_uk_U684 (.ZN( u1_K12_7 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1750 ) , .A( u1_uk_n665 ) );
  NAND2_X1 u1_uk_U685 (.A1( u1_uk_K_r10_19 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n665 ) );
  OAI21_X1 u1_uk_U686 (.ZN( u1_K11_7 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1691 ) , .A( u1_uk_n500 ) );
  NAND2_X1 u1_uk_U687 (.A1( u1_uk_K_r9_33 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n500 ) );
  OAI21_X1 u1_uk_U688 (.ZN( u1_K15_25 ) , .B2( u1_uk_n1876 ) , .B1( u1_uk_n223 ) , .A( u1_uk_n968 ) );
  NAND2_X1 u1_uk_U689 (.A1( u1_uk_K_r13_22 ) , .A2( u1_uk_n213 ) , .ZN( u1_uk_n968 ) );
  OAI22_X1 u1_uk_U690 (.ZN( u1_K11_25 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1677 ) , .A2( u1_uk_n1696 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U691 (.ZN( u1_K13_25 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1765 ) , .A2( u1_uk_n1790 ) , .B1( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U692 (.ZN( u1_K2_25 ) , .A( u1_uk_n1026 ) , .B2( u1_uk_n1294 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U693 (.A1( u1_uk_K_r0_22 ) , .ZN( u1_uk_n1026 ) , .A2( u1_uk_n109 ) );
  OAI22_X1 u1_uk_U694 (.ZN( u1_K16_25 ) , .B2( u1_uk_n1239 ) , .A2( u1_uk_n1246 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U695 (.ZN( u1_K12_25 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1729 ) , .A2( u1_uk_n1734 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U696 (.ZN( u1_K10_25 ) , .A1( u1_uk_n109 ) , .A2( u1_uk_n1623 ) , .B2( u1_uk_n1641 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U697 (.ZN( u1_K8_25 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1563 ) , .A2( u1_uk_n1568 ) , .A1( u1_uk_n214 ) );
  AOI22_X1 u1_uk_U699 (.B2( u1_uk_K_r6_21 ) , .A2( u1_uk_K_r6_28 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1143 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U7 (.ZN( u1_uk_n102 ) , .A( u1_uk_n230 ) );
  AOI22_X1 u1_uk_U70 (.B2( u1_uk_K_r9_45 ) , .A2( u1_uk_K_r9_49 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n443 ) );
  OAI22_X1 u1_uk_U700 (.ZN( u1_K16_3 ) , .B2( u1_uk_n1228 ) , .A2( u1_uk_n1236 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U701 (.ZN( u1_K15_7 ) , .B2( u1_uk_n1853 ) , .A2( u1_uk_n1869 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U702 (.ZN( u1_K16_7 ) , .B2( u1_uk_n1229 ) , .A2( u1_uk_n1237 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U703 (.ZN( u1_K12_3 ) , .A( u1_uk_n601 ) );
  AOI22_X1 u1_uk_U704 (.B2( u1_uk_K_r10_18 ) , .A2( u1_uk_K_r10_27 ) , .B1( u1_uk_n129 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n601 ) );
  AOI22_X1 u1_uk_U706 (.B2( u1_uk_K_r6_10 ) , .A2( u1_uk_K_r6_3 ) , .ZN( u1_uk_n1140 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n294 ) );
  AOI22_X1 u1_uk_U708 (.A2( u1_uk_K_r2_4 ) , .B2( u1_uk_K_r2_41 ) , .ZN( u1_uk_n1065 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n188 ) );
  INV_X1 u1_uk_U71 (.ZN( u1_K8_34 ) , .A( u1_uk_n1137 ) );
  AOI22_X1 u1_uk_U710 (.B2( u1_uk_K_r11_10 ) , .A2( u1_uk_K_r11_5 ) , .B1( u1_uk_n207 ) , .A1( u1_uk_n93 ) , .ZN( u1_uk_n950 ) );
  OAI21_X1 u1_uk_U711 (.ZN( u1_K5_7 ) , .A( u1_uk_n1087 ) , .B2( u1_uk_n1435 ) , .B1( u1_uk_n250 ) );
  NAND2_X1 u1_uk_U712 (.A1( u1_uk_K_r3_19 ) , .ZN( u1_uk_n1087 ) , .A2( u1_uk_n188 ) );
  INV_X1 u1_uk_U713 (.ZN( u1_K1_25 ) , .A( u1_uk_n1005 ) );
  AOI22_X1 u1_uk_U714 (.B2( u1_key_r_29 ) , .A2( u1_key_r_36 ) , .ZN( u1_uk_n1005 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n250 ) );
  AOI22_X1 u1_uk_U716 (.B2( u1_uk_K_r2_16 ) , .A2( u1_uk_K_r2_49 ) , .ZN( u1_uk_n1057 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U717 (.ZN( u1_K12_2 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1711 ) , .B2( u1_uk_n1716 ) , .A1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U718 (.ZN( u1_K10_2 ) , .B2( u1_uk_n1622 ) , .B1( u1_uk_n257 ) , .A( u1_uk_n338 ) );
  NAND2_X1 u1_uk_U719 (.A1( u1_uk_K_r8_41 ) , .A2( u1_uk_n188 ) , .ZN( u1_uk_n338 ) );
  AOI22_X1 u1_uk_U72 (.B2( u1_uk_K_r6_14 ) , .A2( u1_uk_K_r6_21 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1137 ) , .B1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U720 (.ZN( u1_K1_2 ) , .A( u1_uk_n1008 ) , .B2( u1_uk_n1175 ) , .B1( u1_uk_n242 ) );
  NAND2_X1 u1_uk_U721 (.A1( u1_key_r_11 ) , .ZN( u1_uk_n1008 ) , .A2( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U722 (.ZN( u1_K4_32 ) , .A1( u1_uk_n110 ) , .A2( u1_uk_n1356 ) , .B2( u1_uk_n1380 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U723 (.ZN( u1_K16_32 ) , .B2( u1_uk_n1231 ) , .A2( u1_uk_n1239 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U724 (.ZN( u1_K8_32 ) , .B2( u1_uk_n1556 ) , .A2( u1_uk_n1563 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U725 (.ZN( u1_K11_32 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1670 ) , .A2( u1_uk_n1690 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U726 (.ZN( u1_K13_32 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1758 ) , .B2( u1_uk_n1782 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U727 (.ZN( u1_K6_32 ) , .B2( u1_uk_n1448 ) , .A2( u1_uk_n1464 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U728 (.ZN( u1_K3_32 ) , .B2( u1_uk_n1308 ) , .A2( u1_uk_n1343 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U729 (.ZN( u1_K5_32 ) , .B2( u1_uk_n1408 ) , .A2( u1_uk_n1412 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U730 (.ZN( u1_K14_32 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1799 ) , .A2( u1_uk_n1837 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U731 (.ZN( u1_K9_32 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1601 ) , .A2( u1_uk_n1608 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U732 (.ZN( u1_K15_42 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1879 ) , .A2( u1_uk_n1885 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U733 (.ZN( u1_K14_42 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1798 ) , .A2( u1_uk_n1829 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U734 (.ZN( u1_K13_42 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1763 ) , .A2( u1_uk_n1769 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U735 (.ZN( u1_K11_42 ) , .A1( u1_uk_n164 ) , .B2( u1_uk_n1694 ) , .A2( u1_uk_n1702 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U736 (.ZN( u1_K10_42 ) , .B2( u1_uk_n1619 ) , .A1( u1_uk_n162 ) , .A2( u1_uk_n1645 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U737 (.ZN( u1_K4_42 ) , .B2( u1_uk_n1360 ) , .A2( u1_uk_n1367 ) , .B1( u1_uk_n141 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U738 (.ZN( u1_K3_42 ) , .B2( u1_uk_n1307 ) , .A2( u1_uk_n1334 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U739 (.ZN( u1_K2_42 ) , .B2( u1_uk_n1296 ) , .A2( u1_uk_n1304 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U74 (.B2( u1_uk_K_r5_0 ) , .A2( u1_uk_K_r5_35 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1119 ) , .B1( u1_uk_n209 ) );
  AOI22_X1 u1_uk_U741 (.B2( u1_uk_K_r10_28 ) , .A2( u1_uk_K_r10_9 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n294 ) , .ZN( u1_uk_n605 ) );
  AOI22_X1 u1_uk_U743 (.B2( u1_uk_K_r7_15 ) , .A2( u1_uk_K_r7_22 ) , .ZN( u1_uk_n1167 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n291 ) );
  AOI22_X1 u1_uk_U745 (.B2( u1_uk_K_r5_1 ) , .A2( u1_uk_K_r5_36 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1123 ) , .B1( u1_uk_n297 ) );
  INV_X1 u1_uk_U746 (.ZN( u1_K1_42 ) , .A( u1_uk_n1016 ) );
  AOI22_X1 u1_uk_U747 (.B2( u1_key_r_31 ) , .A2( u1_key_r_38 ) , .ZN( u1_uk_n1016 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U748 (.ZN( u1_K14_27 ) , .B2( u1_uk_n1839 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n953 ) );
  NAND2_X1 u1_uk_U749 (.A1( u1_uk_K_r12_42 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n953 ) );
  OAI22_X1 u1_uk_U75 (.ZN( u1_K15_34 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1856 ) , .A2( u1_uk_n1884 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U750 (.ZN( u1_K12_27 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1717 ) , .A2( u1_uk_n1749 ) , .B1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U751 (.ZN( u1_K10_27 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1632 ) , .A( u1_uk_n335 ) );
  NAND2_X1 u1_uk_U752 (.A1( u1_uk_K_r8_43 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n335 ) );
  OAI22_X1 u1_uk_U753 (.ZN( u1_K8_27 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1529 ) , .A2( u1_uk_n1534 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U754 (.ZN( u1_K16_27 ) , .B2( u1_uk_n1225 ) , .A2( u1_uk_n1230 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U755 (.ZN( u1_K12_13 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1719 ) , .A2( u1_uk_n1751 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U756 (.ZN( u1_K11_13 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1688 ) , .A2( u1_uk_n1692 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U757 (.ZN( u1_K8_13 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1531 ) , .B2( u1_uk_n1537 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U758 (.ZN( u1_K6_13 ) , .B2( u1_uk_n1462 ) , .A2( u1_uk_n1466 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U759 (.ZN( u1_K2_13 ) , .A2( u1_uk_n1261 ) , .B2( u1_uk_n1290 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U760 (.ZN( u1_K1_21 ) , .B2( u1_uk_n1183 ) , .A2( u1_uk_n1189 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U761 (.ZN( u1_K9_13 ) , .A( u1_uk_n1150 ) , .B2( u1_uk_n1579 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U762 (.A1( u1_uk_K_r7_5 ) , .ZN( u1_uk_n1150 ) , .A2( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U763 (.ZN( u1_K11_27 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1684 ) , .A2( u1_uk_n1690 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U764 (.ZN( u1_K13_27 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1754 ) , .A2( u1_uk_n1777 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U765 (.ZN( u1_K14_21 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1814 ) , .A2( u1_uk_n1840 ) , .B1( u1_uk_n220 ) );
  OAI21_X1 u1_uk_U766 (.ZN( u1_K11_21 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1667 ) , .A( u1_uk_n395 ) );
  NAND2_X1 u1_uk_U767 (.A1( u1_uk_K_r9_5 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n395 ) );
  OAI22_X1 u1_uk_U768 (.ZN( u1_K9_21 ) , .B2( u1_uk_n1598 ) , .A2( u1_uk_n1603 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U769 (.ZN( u1_K5_21 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1409 ) , .A2( u1_uk_n1429 ) , .B1( u1_uk_n202 ) );
  AOI22_X1 u1_uk_U77 (.B2( u1_uk_K_r12_30 ) , .A2( u1_uk_K_r12_36 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n279 ) , .ZN( u1_uk_n955 ) );
  OAI22_X1 u1_uk_U770 (.ZN( u1_K2_21 ) , .A2( u1_uk_n1264 ) , .B2( u1_uk_n1268 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U771 (.ZN( u1_K7_21 ) , .A( u1_uk_n1110 ) , .B2( u1_uk_n1526 ) , .B1( u1_uk_n271 ) );
  NAND2_X1 u1_uk_U772 (.A1( u1_uk_K_r5_19 ) , .ZN( u1_uk_n1110 ) , .A2( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U773 (.ZN( u1_K4_21 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1371 ) , .A2( u1_uk_n1377 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U774 (.ZN( u1_K15_21 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1846 ) , .B2( u1_uk_n1850 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U775 (.ZN( u1_K14_13 ) , .B2( u1_uk_n1812 ) , .A2( u1_uk_n1817 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U776 (.ZN( u1_K4_27 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1350 ) , .A2( u1_uk_n1376 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U777 (.ZN( u1_K15_27 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1847 ) , .B2( u1_uk_n1865 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U778 (.ZN( u1_K4_13 ) , .A2( u1_uk_n1354 ) , .B2( u1_uk_n1358 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U78 (.ZN( u1_K12_34 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1715 ) , .B2( u1_uk_n1730 ) , .B1( u1_uk_n213 ) );
  AOI22_X1 u1_uk_U780 (.B2( u1_uk_K_r10_25 ) , .A2( u1_uk_K_r10_48 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n250 ) , .ZN( u1_uk_n520 ) );
  AOI22_X1 u1_uk_U782 (.B2( u1_uk_K_r11_11 ) , .A2( u1_uk_K_r11_6 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n240 ) , .ZN( u1_uk_n677 ) );
  INV_X1 u1_uk_U783 (.ZN( u1_K13_21 ) , .A( u1_uk_n689 ) );
  AOI22_X1 u1_uk_U784 (.B2( u1_uk_K_r11_34 ) , .A2( u1_uk_K_r11_39 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n230 ) , .ZN( u1_uk_n689 ) );
  AOI22_X1 u1_uk_U786 (.B2( u1_uk_K_r4_11 ) , .A2( u1_uk_K_r4_5 ) , .ZN( u1_uk_n1092 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U787 (.ZN( u1_K16_13 ) , .B2( u1_uk_n1257 ) , .B1( u1_uk_n297 ) , .A( u1_uk_n980 ) );
  NAND2_X1 u1_uk_U788 (.A1( u1_uk_K_r14_46 ) , .A2( u1_uk_n242 ) , .ZN( u1_uk_n980 ) );
  OAI22_X1 u1_uk_U789 (.ZN( u1_K6_27 ) , .B2( u1_uk_n1459 ) , .A2( u1_uk_n1464 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U79 (.ZN( u1_K6_34 ) , .A( u1_uk_n1097 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1471 ) );
  AOI22_X1 u1_uk_U791 (.B2( u1_uk_K_r3_15 ) , .A2( u1_uk_K_r3_51 ) , .ZN( u1_uk_n1076 ) , .B1( u1_uk_n240 ) , .A1( u1_uk_n83 ) );
  INV_X1 u1_uk_U792 (.ZN( u1_K2_27 ) , .A( u1_uk_n1027 ) );
  AOI22_X1 u1_uk_U793 (.B2( u1_uk_K_r0_28 ) , .A2( u1_uk_K_r0_7 ) , .ZN( u1_uk_n1027 ) , .A1( u1_uk_n129 ) , .B1( u1_uk_n252 ) );
  OAI21_X1 u1_uk_U794 (.ZN( u1_K3_27 ) , .A( u1_uk_n1039 ) , .B2( u1_uk_n1345 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U795 (.A1( u1_uk_K_r1_42 ) , .ZN( u1_uk_n1039 ) , .A2( u1_uk_n298 ) );
  AOI22_X1 u1_uk_U797 (.B2( u1_uk_K_r5_23 ) , .A2( u1_uk_K_r5_43 ) , .ZN( u1_uk_n1115 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n203 ) );
  INV_X1 u1_uk_U798 (.ZN( u1_K1_27 ) , .A( u1_uk_n1007 ) );
  AOI22_X1 u1_uk_U799 (.B2( u1_key_r_14 ) , .A2( u1_key_r_21 ) , .ZN( u1_uk_n1007 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U8 (.A( u1_uk_n203 ) , .ZN( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U80 (.A1( u1_uk_K_r4_49 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1097 ) );
  AOI22_X1 u1_uk_U801 (.B2( u1_uk_K_r7_2 ) , .A2( u1_uk_K_r7_9 ) , .B1( u1_uk_n100 ) , .ZN( u1_uk_n1159 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U802 (.ZN( u1_K16_1 ) , .B2( u1_uk_n1248 ) , .A2( u1_uk_n1251 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U803 (.ZN( u1_K13_1 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1757 ) , .A( u1_uk_n686 ) );
  NAND2_X1 u1_uk_U804 (.A1( u1_uk_K_r11_25 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n686 ) );
  OAI22_X1 u1_uk_U805 (.ZN( u1_K6_1 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1462 ) , .A2( u1_uk_n1478 ) , .B1( u1_uk_n188 ) );
  AOI22_X1 u1_uk_U807 (.B2( u1_uk_K_r7_24 ) , .A2( u1_uk_K_r7_6 ) , .ZN( u1_uk_n1155 ) , .B1( u1_uk_n155 ) , .A1( u1_uk_n250 ) );
  OAI21_X1 u1_uk_U808 (.ZN( u1_K4_1 ) , .A( u1_uk_n1053 ) , .B2( u1_uk_n1353 ) , .B1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U809 (.A1( u1_uk_K_r2_25 ) , .ZN( u1_uk_n1053 ) , .A2( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U81 (.ZN( u1_K4_34 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1366 ) , .A2( u1_uk_n1382 ) , .B1( u1_uk_n202 ) );
  OAI21_X1 u1_uk_U810 (.ZN( u1_K4_18 ) , .A( u1_uk_n1052 ) , .B2( u1_uk_n1378 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U811 (.A1( u1_uk_K_r2_20 ) , .ZN( u1_uk_n1052 ) , .A2( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U812 (.ZN( u1_K5_18 ) , .A2( u1_uk_n1399 ) , .B2( u1_uk_n1436 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U813 (.ZN( u1_K13_20 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1762 ) , .A( u1_uk_n688 ) );
  NAND2_X1 u1_uk_U814 (.A1( u1_uk_K_r11_33 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n688 ) );
  OAI21_X1 u1_uk_U815 (.ZN( u1_K13_18 ) , .B2( u1_uk_n1780 ) , .B1( u1_uk_n231 ) , .A( u1_uk_n682 ) );
  NAND2_X1 u1_uk_U816 (.A1( u1_uk_K_r11_20 ) , .A2( u1_uk_n291 ) , .ZN( u1_uk_n682 ) );
  OAI22_X1 u1_uk_U817 (.ZN( u1_K7_18 ) , .A2( u1_uk_n1483 ) , .B2( u1_uk_n1496 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U818 (.ZN( u1_K8_18 ) , .A( u1_uk_n1132 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1557 ) );
  NAND2_X1 u1_uk_U819 (.A1( u1_uk_K_r6_46 ) , .ZN( u1_uk_n1132 ) , .A2( u1_uk_n146 ) );
  OAI21_X1 u1_uk_U82 (.ZN( u1_K3_34 ) , .B1( u1_uk_n100 ) , .A( u1_uk_n1041 ) , .B2( u1_uk_n1329 ) );
  OAI22_X1 u1_uk_U820 (.ZN( u1_K2_18 ) , .B2( u1_uk_n1269 ) , .A2( u1_uk_n1300 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U821 (.ZN( u1_K16_18 ) , .B2( u1_uk_n1259 ) , .B1( u1_uk_n94 ) , .A( u1_uk_n983 ) );
  NAND2_X1 u1_uk_U822 (.A1( u1_uk_K_r14_5 ) , .A2( u1_uk_n118 ) , .ZN( u1_uk_n983 ) );
  OAI22_X1 u1_uk_U823 (.ZN( u1_K10_18 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1620 ) , .B2( u1_uk_n1634 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U824 (.ZN( u1_K15_18 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1852 ) , .A2( u1_uk_n1882 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U825 (.ZN( u1_K3_20 ) , .B2( u1_uk_n1320 ) , .A2( u1_uk_n1326 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U826 (.ZN( u1_K12_20 ) , .B1( u1_uk_n162 ) , .B2( u1_uk_n1722 ) , .A( u1_uk_n518 ) );
  NAND2_X1 u1_uk_U827 (.A1( u1_uk_K_r10_47 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n518 ) );
  OAI22_X1 u1_uk_U828 (.ZN( u1_K16_20 ) , .B2( u1_uk_n1252 ) , .A2( u1_uk_n1259 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U829 (.ZN( u1_K15_20 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1845 ) , .B2( u1_uk_n1874 ) , .A1( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U83 (.A1( u1_uk_K_r1_36 ) , .ZN( u1_uk_n1041 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U830 (.ZN( u1_K8_20 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1551 ) , .A2( u1_uk_n1557 ) , .A1( u1_uk_n222 ) );
  AOI22_X1 u1_uk_U832 (.B2( u1_uk_K_r7_39 ) , .A2( u1_uk_K_r7_46 ) , .ZN( u1_uk_n1153 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n230 ) );
  AOI22_X1 u1_uk_U834 (.B2( u1_uk_K_r4_11 ) , .A2( u1_uk_K_r4_17 ) , .ZN( u1_uk_n1090 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n252 ) );
  INV_X1 u1_uk_U835 (.ZN( u1_K11_20 ) , .A( u1_uk_n391 ) );
  AOI22_X1 u1_uk_U836 (.B2( u1_uk_K_r9_10 ) , .A2( u1_uk_K_r9_4 ) , .A1( u1_uk_n100 ) , .B1( u1_uk_n292 ) , .ZN( u1_uk_n391 ) );
  AOI22_X1 u1_uk_U838 (.B2( u1_uk_K_r5_18 ) , .A2( u1_uk_K_r5_53 ) , .A1( u1_uk_n11 ) , .ZN( u1_uk_n1109 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U84 (.ZN( u1_K2_34 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1272 ) , .A2( u1_uk_n1303 ) , .A1( u1_uk_n217 ) );
  AOI22_X1 u1_uk_U840 (.B2( u1_uk_K_r3_24 ) , .A2( u1_uk_K_r3_47 ) , .ZN( u1_uk_n1073 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U841 (.ZN( u1_K4_22 ) , .A( u1_uk_n1055 ) , .B2( u1_uk_n1357 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U842 (.A1( u1_uk_K_r2_47 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n1055 ) );
  OAI22_X1 u1_uk_U843 (.ZN( u1_K1_6 ) , .B2( u1_uk_n1198 ) , .A2( u1_uk_n1205 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n240 ) );
  INV_X1 u1_uk_U844 (.A( u1_key_r_41 ) , .ZN( u1_uk_n1205 ) );
  OAI22_X1 u1_uk_U845 (.ZN( u1_K15_6 ) , .B2( u1_uk_n1864 ) , .A2( u1_uk_n1882 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U846 (.ZN( u1_K1_43 ) , .A2( u1_uk_n1179 ) , .B2( u1_uk_n1182 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U847 (.ZN( u1_K13_3 ) , .B2( u1_uk_n1781 ) , .B1( u1_uk_n27 ) , .A( u1_uk_n945 ) );
  NAND2_X1 u1_uk_U848 (.A1( u1_uk_K_r11_4 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n945 ) );
  OAI22_X1 u1_uk_U849 (.ZN( u1_K7_3 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1495 ) , .A2( u1_uk_n1517 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U85 (.ZN( u1_K16_23 ) , .B2( u1_uk_n1243 ) , .A2( u1_uk_n1248 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U850 (.ZN( u1_K15_3 ) , .B2( u1_uk_n1852 ) , .A2( u1_uk_n1868 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n83 ) );
  AOI22_X1 u1_uk_U852 (.B2( u1_uk_K_r5_39 ) , .A2( u1_uk_K_r5_4 ) , .ZN( u1_uk_n1125 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U853 (.ZN( u1_K14_3 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1842 ) , .A( u1_uk_n957 ) );
  NAND2_X1 u1_uk_U854 (.A1( u1_uk_K_r12_47 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n957 ) );
  OAI21_X1 u1_uk_U855 (.ZN( u1_K3_3 ) , .A( u1_uk_n1043 ) , .B2( u1_uk_n1348 ) , .B1( u1_uk_n242 ) );
  NAND2_X1 u1_uk_U856 (.A1( u1_uk_K_r1_47 ) , .ZN( u1_uk_n1043 ) , .A2( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U857 (.ZN( u1_K16_2 ) , .B2( u1_uk_n1220 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n986 ) );
  NAND2_X1 u1_uk_U858 (.A1( u1_uk_K_r14_11 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n986 ) );
  AOI22_X1 u1_uk_U859 (.B2( u1_uk_K_r7_20 ) , .A2( u1_uk_K_r7_27 ) , .ZN( u1_uk_n1160 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n286 ) );
  AOI22_X1 u1_uk_U860 (.B2( u1_uk_K_r2_26 ) , .A2( u1_uk_K_r2_46 ) , .ZN( u1_uk_n1061 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U861 (.ZN( u1_K10_1 ) , .B2( u1_uk_n1630 ) , .A( u1_uk_n306 ) , .B1( u1_uk_n31 ) );
  NAND2_X1 u1_uk_U862 (.A1( u1_uk_K_r8_10 ) , .A2( u1_uk_n118 ) , .ZN( u1_uk_n306 ) );
  OAI22_X1 u1_uk_U863 (.ZN( u1_K1_1 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1204 ) , .A2( u1_uk_n1209 ) , .B1( u1_uk_n240 ) );
  AOI22_X1 u1_uk_U864 (.B2( u1_uk_K_r10_39 ) , .A2( u1_uk_K_r10_48 ) , .B1( u1_uk_n155 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n515 ) );
  AOI22_X1 u1_uk_U865 (.B2( u1_uk_K_r11_19 ) , .A2( u1_uk_K_r11_24 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) , .ZN( u1_uk_n949 ) );
  OAI22_X1 u1_uk_U866 (.ZN( u1_K3_18 ) , .B2( u1_uk_n1325 ) , .A2( u1_uk_n1332 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U867 (.ZN( u1_K14_22 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1802 ) , .A2( u1_uk_n1840 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U868 (.ZN( u1_K10_5 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1625 ) , .A2( u1_uk_n1642 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U869 (.ZN( u1_K5_41 ) , .B2( u1_uk_n1418 ) , .A2( u1_uk_n1426 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U87 (.B2( u1_uk_K_r10_32 ) , .A2( u1_uk_K_r10_41 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n238 ) , .ZN( u1_uk_n524 ) );
  OAI22_X1 u1_uk_U870 (.ZN( u1_K15_22 ) , .B2( u1_uk_n1858 ) , .A2( u1_uk_n1872 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U871 (.ZN( u1_K6_22 ) , .B2( u1_uk_n1447 ) , .A2( u1_uk_n1452 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U872 (.ZN( u1_K15_23 ) , .B2( u1_uk_n1863 ) , .A2( u1_uk_n1881 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U873 (.ZN( u1_K14_23 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1802 ) , .B2( u1_uk_n1809 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U874 (.ZN( u1_K5_23 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1415 ) , .A2( u1_uk_n1424 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U875 (.ZN( u1_K13_34 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1768 ) , .A2( u1_uk_n1784 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U876 (.ZN( u1_K5_34 ) , .B1( u1_uk_n118 ) , .A2( u1_uk_n1401 ) , .B2( u1_uk_n1414 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U877 (.ZN( u1_K3_47 ) , .B2( u1_uk_n1327 ) , .A2( u1_uk_n1335 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U878 (.ZN( u1_K8_5 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1564 ) , .A2( u1_uk_n1570 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U879 (.ZN( u1_K6_5 ) , .B2( u1_uk_n1452 ) , .A2( u1_uk_n1456 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U88 (.ZN( u1_K11_23 ) , .B2( u1_uk_n1698 ) , .B1( u1_uk_n292 ) , .A( u1_uk_n408 ) );
  OAI22_X1 u1_uk_U880 (.ZN( u1_K12_10 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1718 ) , .A2( u1_uk_n1739 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U881 (.ZN( u1_K12_11 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1713 ) , .B2( u1_uk_n1739 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U882 (.ZN( u1_K7_10 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1487 ) , .A2( u1_uk_n1517 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U883 (.B1( n116 ) , .ZN( u1_K4_11 ) , .B2( u1_uk_n1363 ) , .A2( u1_uk_n1391 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U884 (.ZN( u1_K3_10 ) , .B2( u1_uk_n1316 ) , .A2( u1_uk_n1321 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U885 (.ZN( u1_K15_45 ) , .B2( u1_uk_n1867 ) , .A2( u1_uk_n1885 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U886 (.ZN( u1_K13_45 ) , .B1( u1_uk_n162 ) , .B2( u1_uk_n1755 ) , .A2( u1_uk_n1793 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U887 (.ZN( u1_K12_43 ) , .B2( u1_uk_n1717 ) , .A2( u1_uk_n1737 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U888 (.ZN( u1_K6_45 ) , .B2( u1_uk_n1454 ) , .A2( u1_uk_n1459 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U889 (.ZN( u1_K3_30 ) , .B2( u1_uk_n1318 ) , .A2( u1_uk_n1344 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U89 (.A1( u1_uk_K_r9_27 ) , .A2( u1_uk_n298 ) , .ZN( u1_uk_n408 ) );
  OAI22_X1 u1_uk_U890 (.ZN( u1_K8_1 ) , .B1( u1_uk_n146 ) , .A2( u1_uk_n1532 ) , .B2( u1_uk_n1548 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U891 (.ZN( u1_K14_6 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1803 ) , .B2( u1_uk_n1810 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U892 (.ZN( u1_K10_3 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1633 ) , .A2( u1_uk_n1653 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U893 (.ZN( u1_K9_3 ) , .B1( u1_uk_n147 ) , .A2( u1_uk_n1573 ) , .B2( u1_uk_n1577 ) , .A1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U894 (.ZN( u1_K9_7 ) , .B1( u1_uk_n146 ) , .A2( u1_uk_n1574 ) , .B2( u1_uk_n1578 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U895 (.ZN( u1_K6_12 ) , .A2( u1_uk_n1440 ) , .B2( u1_uk_n1456 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U896 (.ZN( u1_K5_3 ) , .B2( u1_uk_n1404 ) , .A2( u1_uk_n1411 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U897 (.ZN( u1_K7_14 ) , .B2( u1_uk_n1492 ) , .A2( u1_uk_n1527 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U898 (.ZN( u1_K14_7 ) , .B2( u1_uk_n1816 ) , .A2( u1_uk_n1835 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U899 (.ZN( u1_K13_24 ) , .B2( u1_uk_n1756 ) , .A2( u1_uk_n1797 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n99 ) );
  INV_X1 u1_uk_U9 (.A( u1_uk_n209 ) , .ZN( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U90 (.ZN( u1_K10_23 ) , .B2( u1_uk_n1620 ) , .B1( u1_uk_n294 ) , .A( u1_uk_n313 ) );
  OAI22_X1 u1_uk_U900 (.ZN( u1_K6_24 ) , .B2( u1_uk_n1457 ) , .A2( u1_uk_n1461 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U901 (.ZN( u1_K15_13 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1844 ) , .B2( u1_uk_n1872 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U902 (.ZN( u1_K3_21 ) , .B2( u1_uk_n1321 ) , .A2( u1_uk_n1346 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U903 (.ZN( u1_K9_24 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1574 ) , .A2( u1_uk_n1616 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U904 (.ZN( u1_K5_19 ) , .A2( u1_uk_n1398 ) , .B2( u1_uk_n1435 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U905 (.ZN( u1_K5_24 ) , .B2( u1_uk_n1402 ) , .A2( u1_uk_n1427 ) , .B1( u1_uk_n145 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U906 (.ZN( u1_K2_24 ) , .A2( u1_uk_n1264 ) , .B2( u1_uk_n1279 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U907 (.ZN( u1_K16_21 ) , .B2( u1_uk_n1227 ) , .A2( u1_uk_n1234 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U908 (.ZN( u1_K8_21 ) , .B2( u1_uk_n1552 ) , .A2( u1_uk_n1558 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U909 (.ZN( u1_K16_24 ) , .B2( u1_uk_n1224 ) , .A2( u1_uk_n1229 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U91 (.A1( u1_uk_K_r8_13 ) , .A2( u1_uk_n271 ) , .ZN( u1_uk_n313 ) );
  OAI22_X1 u1_uk_U910 (.ZN( u1_K7_30 ) , .B2( u1_uk_n1490 ) , .A2( u1_uk_n1521 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U911 (.ZN( u1_K5_13 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1405 ) , .A2( u1_uk_n1436 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U912 (.ZN( u1_K5_14 ) , .B2( u1_uk_n1403 ) , .B1( u1_uk_n141 ) , .A2( u1_uk_n1410 ) , .A1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U913 (.ZN( u1_K4_14 ) , .B1( u1_uk_n110 ) , .B2( u1_uk_n1352 ) , .A2( u1_uk_n1378 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U914 (.ZN( u1_K3_13 ) , .B2( u1_uk_n1319 ) , .A2( u1_uk_n1324 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U915 (.ZN( u1_K4_36 ) , .B2( u1_uk_n1376 ) , .A2( u1_uk_n1381 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U916 (.ZN( u1_K2_17 ) , .A2( u1_uk_n1261 ) , .B2( u1_uk_n1277 ) , .A1( u1_uk_n291 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U917 (.ZN( u1_K6_30 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1438 ) , .A2( u1_uk_n1443 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U918 (.ZN( u1_K3_25 ) , .B2( u1_uk_n1309 ) , .A2( u1_uk_n1313 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U919 (.ZN( u1_K16_38 ) , .B2( u1_uk_n1240 ) , .A2( u1_uk_n1247 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U92 (.ZN( u1_K8_23 ) , .B2( u1_uk_n1543 ) , .A2( u1_uk_n1548 ) , .A1( u1_uk_n279 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U920 (.ZN( u1_K8_38 ) , .B1( u1_uk_n145 ) , .B2( u1_uk_n1560 ) , .A2( u1_uk_n1566 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U921 (.ZN( u1_K7_39 ) , .B2( u1_uk_n1516 ) , .A2( u1_uk_n1523 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U922 (.ZN( u1_K6_42 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1468 ) , .A2( u1_uk_n1475 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U923 (.ZN( u1_K6_39 ) , .A2( u1_uk_n1441 ) , .B2( u1_uk_n1460 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U924 (.ZN( u1_K4_39 ) , .B2( u1_uk_n1351 ) , .A2( u1_uk_n1372 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U925 (.ZN( u1_K3_38 ) , .A2( u1_uk_n1314 ) , .B2( u1_uk_n1330 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U926 (.ZN( u1_K3_39 ) , .B2( u1_uk_n1338 ) , .A2( u1_uk_n1342 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U927 (.ZN( u1_K2_39 ) , .A2( u1_uk_n1266 ) , .B2( u1_uk_n1281 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U928 (.ZN( u1_K13_23 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1767 ) , .A2( u1_uk_n1797 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U929 (.ZN( u1_K9_23 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1584 ) , .A2( u1_uk_n1592 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U93 (.ZN( u1_K3_23 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1311 ) , .B2( u1_uk_n1316 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U930 (.ZN( u1_K9_47 ) , .B2( u1_uk_n1606 ) , .A2( u1_uk_n1613 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U931 (.ZN( u1_K12_16 ) , .A2( u1_uk_n1711 ) , .B2( u1_uk_n1723 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U932 (.ZN( u1_K11_16 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1692 ) , .A2( u1_uk_n1698 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U933 (.ZN( u1_K11_48 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1689 ) , .A2( u1_uk_n1696 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U934 (.ZN( u1_K11_6 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1699 ) , .A2( u1_uk_n1705 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U935 (.ZN( u1_K9_6 ) , .B2( u1_uk_n1585 ) , .A2( u1_uk_n1593 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U936 (.ZN( u1_K9_8 ) , .B2( u1_uk_n1603 ) , .A2( u1_uk_n1610 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U937 (.ZN( u1_K14_8 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1801 ) , .B2( u1_uk_n1819 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U938 (.ZN( u1_K12_18 ) , .A1( u1_uk_n164 ) , .A2( u1_uk_n1713 ) , .B2( u1_uk_n1751 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U939 (.ZN( u1_K14_20 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1813 ) , .A2( u1_uk_n1819 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U94 (.ZN( u1_K2_23 ) , .B2( u1_uk_n1278 ) , .A2( u1_uk_n1299 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U940 (.ZN( u1_K2_20 ) , .A2( u1_uk_n1263 ) , .B2( u1_uk_n1292 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U941 (.ZN( u1_K11_24 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1682 ) , .A2( u1_uk_n1687 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U942 (.ZN( u1_K14_14 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1834 ) , .A2( u1_uk_n1841 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U943 (.ZN( u1_K8_24 ) , .B2( u1_uk_n1530 ) , .A1( u1_uk_n155 ) , .A2( u1_uk_n1570 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U944 (.ZN( u1_K16_46 ) , .B2( u1_uk_n1219 ) , .A2( u1_uk_n1253 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U945 (.ZN( u1_K15_47 ) , .B2( u1_uk_n1854 ) , .A2( u1_uk_n1886 ) , .B1( u1_uk_n208 ) , .A1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U946 (.ZN( u1_K14_47 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1820 ) , .A2( u1_uk_n1830 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U947 (.ZN( u1_K10_46 ) , .B2( u1_uk_n1632 ) , .A2( u1_uk_n1641 ) , .B1( u1_uk_n279 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U948 (.ZN( u1_K10_34 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1618 ) , .A2( u1_uk_n1644 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U949 (.ZN( u1_K9_34 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1581 ) , .A2( u1_uk_n1588 ) , .B1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U95 (.ZN( u1_K11_41 ) , .B2( u1_uk_n1702 ) , .B1( u1_uk_n217 ) , .A( u1_uk_n467 ) );
  OAI22_X1 u1_uk_U950 (.ZN( u1_K6_46 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1443 ) , .B2( u1_uk_n1471 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U951 (.ZN( u1_K13_4 ) , .A1( u1_uk_n155 ) , .B2( u1_uk_n1762 ) , .A2( u1_uk_n1767 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U952 (.ZN( u1_K9_4 ) , .A1( u1_uk_n10 ) , .B2( u1_uk_n1579 ) , .A2( u1_uk_n1586 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U953 (.ZN( u1_K4_48 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1355 ) , .B2( u1_uk_n1383 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U954 (.ZN( u1_K2_48 ) , .B2( u1_uk_n1271 ) , .A2( u1_uk_n1286 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U955 (.ZN( u1_K10_8 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1621 ) , .B2( u1_uk_n1635 ) , .B1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U956 (.ZN( u1_K13_8 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1781 ) , .A2( u1_uk_n1787 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U957 (.ZN( u1_K6_20 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1439 ) , .B2( u1_uk_n1444 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U958 (.ZN( u1_K11_18 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1667 ) , .A2( u1_uk_n1673 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U959 (.ZN( u1_K14_18 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1818 ) , .A2( u1_uk_n1826 ) , .B1( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U96 (.A1( u1_uk_K_r9_31 ) , .A2( u1_uk_n203 ) , .ZN( u1_uk_n467 ) );
  OAI22_X1 u1_uk_U960 (.ZN( u1_K12_19 ) , .A1( u1_uk_n110 ) , .A2( u1_uk_n1712 ) , .B2( u1_uk_n1750 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U961 (.ZN( u1_K16_19 ) , .B2( u1_uk_n1220 ) , .A2( u1_uk_n1258 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U962 (.ZN( u1_K15_19 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1851 ) , .A2( u1_uk_n1881 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U963 (.ZN( u1_K10_20 ) , .B2( u1_uk_n1629 ) , .A1( u1_uk_n163 ) , .A2( u1_uk_n1659 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U964 (.ZN( u1_K14_16 ) , .A1( u1_uk_n142 ) , .A2( u1_uk_n1804 ) , .B2( u1_uk_n1842 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U965 (.ZN( u1_K6_36 ) , .A1( u1_uk_n11 ) , .A2( u1_uk_n1441 ) , .B2( u1_uk_n1449 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U966 (.ZN( u1_K14_38 ) , .A2( u1_uk_n1807 ) , .B2( u1_uk_n1823 ) , .B1( u1_uk_n230 ) , .A1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U967 (.ZN( u1_K13_38 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1785 ) , .A2( u1_uk_n1791 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U968 (.ZN( u1_K2_38 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1276 ) , .A2( u1_uk_n1295 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U969 (.ZN( u1_K7_37 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1499 ) , .A2( u1_uk_n1523 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U970 (.ZN( u1_K2_37 ) , .A2( u1_uk_n1267 ) , .B2( u1_uk_n1294 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U971 (.ZN( u1_K9_40 ) , .B2( u1_uk_n1600 ) , .A2( u1_uk_n1606 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U972 (.ZN( u1_K5_40 ) , .B2( u1_uk_n1413 ) , .A2( u1_uk_n1430 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U973 (.ZN( u1_K2_22 ) , .B2( u1_uk_n1273 ) , .A2( u1_uk_n1290 ) , .B1( u1_uk_n222 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U974 (.ZN( u1_K8_45 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1528 ) , .A2( u1_uk_n1566 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U975 (.ZN( u1_K11_45 ) , .A1( u1_uk_n161 ) , .B2( u1_uk_n1677 ) , .A2( u1_uk_n1684 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U976 (.ZN( u1_K7_45 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1490 ) , .A2( u1_uk_n1507 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U977 (.ZN( u1_K6_43 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1438 ) , .A2( u1_uk_n1477 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U978 (.ZN( u1_K4_45 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1351 ) , .A2( u1_uk_n1390 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U979 (.ZN( u1_K2_45 ) , .B2( u1_uk_n1282 ) , .A2( u1_uk_n1304 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U98 (.B2( u1_uk_K_r7_23 ) , .A2( u1_uk_K_r7_30 ) , .ZN( u1_uk_n1166 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U980 (.ZN( u1_K2_3 ) , .B2( u1_uk_n1269 ) , .A2( u1_uk_n1284 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U981 (.ZN( u1_K6_3 ) , .B2( u1_uk_n1447 ) , .A2( u1_uk_n1461 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U982 (.ZN( u1_K3_6 ) , .A2( u1_uk_n1312 ) , .B2( u1_uk_n1317 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U983 (.ZN( u1_K8_7 ) , .A2( u1_uk_n1530 ) , .B2( u1_uk_n1536 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U984 (.ZN( u1_K7_7 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1496 ) , .A2( u1_uk_n1518 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U985 (.ZN( u1_K3_7 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1323 ) , .A2( u1_uk_n1341 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U986 (.ZN( u1_K9_15 ) , .B2( u1_uk_n1577 ) , .A2( u1_uk_n1584 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U987 (.ZN( u1_K6_15 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1453 ) , .A2( u1_uk_n1465 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U988 (.ZN( u1_K6_25 ) , .B2( u1_uk_n1454 ) , .A2( u1_uk_n1470 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U989 (.ZN( u1_K14_25 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1800 ) , .A2( u1_uk_n1806 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U990 (.ZN( u1_K1_23 ) , .B2( u1_uk_n1197 ) , .A2( u1_uk_n1204 ) , .A1( u1_uk_n128 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U991 (.ZN( u1_K1_34 ) , .B2( u1_uk_n1174 ) , .A2( u1_uk_n1179 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U992 (.ZN( u1_K1_47 ) , .B2( u1_uk_n1172 ) , .A2( u1_uk_n1177 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U993 (.ZN( u1_K1_3 ) , .B2( u1_uk_n1184 ) , .A2( u1_uk_n1191 ) , .A1( u1_uk_n128 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U994 (.ZN( u1_K5_25 ) , .A( u1_uk_n1075 ) , .B2( u1_uk_n1413 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U995 (.A1( u1_uk_K_r3_35 ) , .ZN( u1_uk_n1075 ) , .A2( u1_uk_n63 ) );
  OAI21_X1 u1_uk_U996 (.ZN( u1_K7_22 ) , .A( u1_uk_n1111 ) , .B2( u1_uk_n1498 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U997 (.A1( u1_uk_K_r5_5 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1111 ) );
  OAI21_X1 u1_uk_U998 (.ZN( u1_K7_23 ) , .A( u1_uk_n1112 ) , .B2( u1_uk_n1483 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U999 (.A1( u1_uk_K_r5_13 ) , .ZN( u1_uk_n1112 ) , .A2( u1_uk_n17 ) );
  DFF_X1 u2_L0_reg_1 (.CK( clk ) , .Q( u2_L0_1 ) , .D( u2_desIn_r_7 ) );
  DFF_X1 u2_L0_reg_10 (.CK( clk ) , .Q( u2_L0_10 ) , .D( u2_desIn_r_13 ) );
  DFF_X1 u2_L0_reg_11 (.CK( clk ) , .Q( u2_L0_11 ) , .D( u2_desIn_r_21 ) );
  DFF_X1 u2_L0_reg_12 (.CK( clk ) , .Q( u2_L0_12 ) , .D( u2_desIn_r_29 ) );
  DFF_X1 u2_L0_reg_13 (.CK( clk ) , .Q( u2_L0_13 ) , .D( u2_desIn_r_37 ) );
  DFF_X1 u2_L0_reg_14 (.CK( clk ) , .Q( u2_L0_14 ) , .D( u2_desIn_r_45 ) );
  DFF_X1 u2_L0_reg_15 (.CK( clk ) , .Q( u2_L0_15 ) , .D( u2_desIn_r_53 ) );
  DFF_X1 u2_L0_reg_16 (.CK( clk ) , .Q( u2_L0_16 ) , .D( u2_desIn_r_61 ) );
  DFF_X1 u2_L0_reg_17 (.CK( clk ) , .Q( u2_L0_17 ) , .D( u2_desIn_r_3 ) );
  DFF_X1 u2_L0_reg_18 (.CK( clk ) , .Q( u2_L0_18 ) , .D( u2_desIn_r_11 ) );
  DFF_X1 u2_L0_reg_19 (.CK( clk ) , .Q( u2_L0_19 ) , .D( u2_desIn_r_19 ) );
  DFF_X1 u2_L0_reg_2 (.CK( clk ) , .Q( u2_L0_2 ) , .D( u2_desIn_r_15 ) );
  DFF_X1 u2_L0_reg_20 (.CK( clk ) , .Q( u2_L0_20 ) , .D( u2_desIn_r_27 ) );
  DFF_X1 u2_L0_reg_21 (.CK( clk ) , .Q( u2_L0_21 ) , .D( u2_desIn_r_35 ) );
  DFF_X1 u2_L0_reg_22 (.CK( clk ) , .Q( u2_L0_22 ) , .D( u2_desIn_r_43 ) );
  DFF_X1 u2_L0_reg_23 (.CK( clk ) , .Q( u2_L0_23 ) , .D( u2_desIn_r_51 ) );
  DFF_X1 u2_L0_reg_24 (.CK( clk ) , .Q( u2_L0_24 ) , .D( u2_desIn_r_59 ) );
  DFF_X1 u2_L0_reg_25 (.CK( clk ) , .Q( u2_L0_25 ) , .D( u2_desIn_r_1 ) );
  DFF_X1 u2_L0_reg_26 (.CK( clk ) , .Q( u2_L0_26 ) , .D( u2_desIn_r_9 ) );
  DFF_X1 u2_L0_reg_27 (.CK( clk ) , .Q( u2_L0_27 ) , .D( u2_desIn_r_17 ) );
  DFF_X1 u2_L0_reg_28 (.CK( clk ) , .Q( u2_L0_28 ) , .D( u2_desIn_r_25 ) );
  DFF_X1 u2_L0_reg_29 (.CK( clk ) , .Q( u2_L0_29 ) , .D( u2_desIn_r_33 ) );
  DFF_X1 u2_L0_reg_3 (.CK( clk ) , .Q( u2_L0_3 ) , .D( u2_desIn_r_23 ) );
  DFF_X1 u2_L0_reg_30 (.CK( clk ) , .Q( u2_L0_30 ) , .D( u2_desIn_r_41 ) );
  DFF_X1 u2_L0_reg_31 (.CK( clk ) , .Q( u2_L0_31 ) , .D( u2_desIn_r_49 ) );
  DFF_X1 u2_L0_reg_32 (.CK( clk ) , .Q( u2_L0_32 ) , .D( u2_desIn_r_57 ) );
  DFF_X1 u2_L0_reg_4 (.CK( clk ) , .Q( u2_L0_4 ) , .D( u2_desIn_r_31 ) );
  DFF_X1 u2_L0_reg_5 (.CK( clk ) , .Q( u2_L0_5 ) , .D( u2_desIn_r_39 ) );
  DFF_X1 u2_L0_reg_6 (.CK( clk ) , .Q( u2_L0_6 ) , .D( u2_desIn_r_47 ) );
  DFF_X1 u2_L0_reg_7 (.CK( clk ) , .Q( u2_L0_7 ) , .D( u2_desIn_r_55 ) );
  DFF_X1 u2_L0_reg_8 (.CK( clk ) , .Q( u2_L0_8 ) , .D( u2_desIn_r_63 ) );
  DFF_X1 u2_L0_reg_9 (.CK( clk ) , .Q( u2_L0_9 ) , .D( u2_desIn_r_5 ) );
  DFF_X1 u2_L10_reg_1 (.CK( clk ) , .Q( u2_L10_1 ) , .D( u2_R9_1 ) );
  DFF_X1 u2_L10_reg_10 (.CK( clk ) , .Q( u2_L10_10 ) , .D( u2_R9_10 ) );
  DFF_X1 u2_L10_reg_11 (.CK( clk ) , .Q( u2_L10_11 ) , .D( u2_R9_11 ) );
  DFF_X1 u2_L10_reg_12 (.CK( clk ) , .Q( u2_L10_12 ) , .D( u2_R9_12 ) );
  DFF_X1 u2_L10_reg_13 (.CK( clk ) , .Q( u2_L10_13 ) , .D( u2_R9_13 ) );
  DFF_X1 u2_L10_reg_14 (.CK( clk ) , .Q( u2_L10_14 ) , .D( u2_R9_14 ) );
  DFF_X1 u2_L10_reg_15 (.CK( clk ) , .Q( u2_L10_15 ) , .D( u2_R9_15 ) );
  DFF_X1 u2_L10_reg_16 (.CK( clk ) , .Q( u2_L10_16 ) , .D( u2_R9_16 ) );
  DFF_X1 u2_L10_reg_17 (.CK( clk ) , .Q( u2_L10_17 ) , .D( u2_R9_17 ) );
  DFF_X1 u2_L10_reg_18 (.CK( clk ) , .Q( u2_L10_18 ) , .D( u2_R9_18 ) );
  DFF_X1 u2_L10_reg_19 (.CK( clk ) , .Q( u2_L10_19 ) , .D( u2_R9_19 ) );
  DFF_X1 u2_L10_reg_2 (.CK( clk ) , .Q( u2_L10_2 ) , .D( u2_R9_2 ) );
  DFF_X1 u2_L10_reg_20 (.CK( clk ) , .Q( u2_L10_20 ) , .D( u2_R9_20 ) );
  DFF_X1 u2_L10_reg_21 (.CK( clk ) , .Q( u2_L10_21 ) , .D( u2_R9_21 ) );
  DFF_X1 u2_L10_reg_22 (.CK( clk ) , .Q( u2_L10_22 ) , .D( u2_R9_22 ) );
  DFF_X1 u2_L10_reg_23 (.CK( clk ) , .Q( u2_L10_23 ) , .D( u2_R9_23 ) );
  DFF_X1 u2_L10_reg_24 (.CK( clk ) , .Q( u2_L10_24 ) , .D( u2_R9_24 ) );
  DFF_X1 u2_L10_reg_25 (.CK( clk ) , .Q( u2_L10_25 ) , .D( u2_R9_25 ) );
  DFF_X1 u2_L10_reg_26 (.CK( clk ) , .Q( u2_L10_26 ) , .D( u2_R9_26 ) );
  DFF_X1 u2_L10_reg_27 (.CK( clk ) , .Q( u2_L10_27 ) , .D( u2_R9_27 ) );
  DFF_X1 u2_L10_reg_28 (.CK( clk ) , .Q( u2_L10_28 ) , .D( u2_R9_28 ) );
  DFF_X1 u2_L10_reg_29 (.CK( clk ) , .Q( u2_L10_29 ) , .D( u2_R9_29 ) );
  DFF_X1 u2_L10_reg_3 (.CK( clk ) , .Q( u2_L10_3 ) , .D( u2_R9_3 ) );
  DFF_X1 u2_L10_reg_30 (.CK( clk ) , .Q( u2_L10_30 ) , .D( u2_R9_30 ) );
  DFF_X1 u2_L10_reg_31 (.CK( clk ) , .Q( u2_L10_31 ) , .D( u2_R9_31 ) );
  DFF_X1 u2_L10_reg_32 (.CK( clk ) , .Q( u2_L10_32 ) , .D( u2_R9_32 ) );
  DFF_X1 u2_L10_reg_4 (.CK( clk ) , .Q( u2_L10_4 ) , .D( u2_R9_4 ) );
  DFF_X1 u2_L10_reg_5 (.CK( clk ) , .Q( u2_L10_5 ) , .D( u2_R9_5 ) );
  DFF_X1 u2_L10_reg_6 (.CK( clk ) , .Q( u2_L10_6 ) , .D( u2_R9_6 ) );
  DFF_X1 u2_L10_reg_7 (.CK( clk ) , .Q( u2_L10_7 ) , .D( u2_R9_7 ) );
  DFF_X1 u2_L10_reg_8 (.CK( clk ) , .Q( u2_L10_8 ) , .D( u2_R9_8 ) );
  DFF_X1 u2_L10_reg_9 (.CK( clk ) , .Q( u2_L10_9 ) , .D( u2_R9_9 ) );
  DFF_X1 u2_L11_reg_1 (.CK( clk ) , .Q( u2_L11_1 ) , .D( u2_R10_1 ) );
  DFF_X1 u2_L11_reg_10 (.CK( clk ) , .Q( u2_L11_10 ) , .D( u2_R10_10 ) );
  DFF_X1 u2_L11_reg_11 (.CK( clk ) , .Q( u2_L11_11 ) , .D( u2_R10_11 ) );
  DFF_X1 u2_L11_reg_12 (.CK( clk ) , .Q( u2_L11_12 ) , .D( u2_R10_12 ) );
  DFF_X1 u2_L11_reg_13 (.CK( clk ) , .Q( u2_L11_13 ) , .D( u2_R10_13 ) );
  DFF_X1 u2_L11_reg_14 (.CK( clk ) , .Q( u2_L11_14 ) , .D( u2_R10_14 ) );
  DFF_X1 u2_L11_reg_15 (.CK( clk ) , .Q( u2_L11_15 ) , .D( u2_R10_15 ) );
  DFF_X1 u2_L11_reg_16 (.CK( clk ) , .Q( u2_L11_16 ) , .D( u2_R10_16 ) );
  DFF_X1 u2_L11_reg_17 (.CK( clk ) , .Q( u2_L11_17 ) , .D( u2_R10_17 ) );
  DFF_X1 u2_L11_reg_18 (.CK( clk ) , .Q( u2_L11_18 ) , .D( u2_R10_18 ) );
  DFF_X1 u2_L11_reg_19 (.CK( clk ) , .Q( u2_L11_19 ) , .D( u2_R10_19 ) );
  DFF_X1 u2_L11_reg_2 (.CK( clk ) , .Q( u2_L11_2 ) , .D( u2_R10_2 ) );
  DFF_X1 u2_L11_reg_20 (.CK( clk ) , .Q( u2_L11_20 ) , .D( u2_R10_20 ) );
  DFF_X1 u2_L11_reg_21 (.CK( clk ) , .Q( u2_L11_21 ) , .D( u2_R10_21 ) );
  DFF_X1 u2_L11_reg_22 (.CK( clk ) , .Q( u2_L11_22 ) , .D( u2_R10_22 ) );
  DFF_X1 u2_L11_reg_23 (.CK( clk ) , .Q( u2_L11_23 ) , .D( u2_R10_23 ) );
  DFF_X1 u2_L11_reg_24 (.CK( clk ) , .Q( u2_L11_24 ) , .D( u2_R10_24 ) );
  DFF_X1 u2_L11_reg_25 (.CK( clk ) , .Q( u2_L11_25 ) , .D( u2_R10_25 ) );
  DFF_X1 u2_L11_reg_26 (.CK( clk ) , .Q( u2_L11_26 ) , .D( u2_R10_26 ) );
  DFF_X1 u2_L11_reg_27 (.CK( clk ) , .Q( u2_L11_27 ) , .D( u2_R10_27 ) );
  DFF_X1 u2_L11_reg_28 (.CK( clk ) , .Q( u2_L11_28 ) , .D( u2_R10_28 ) );
  DFF_X1 u2_L11_reg_29 (.CK( clk ) , .Q( u2_L11_29 ) , .D( u2_R10_29 ) );
  DFF_X1 u2_L11_reg_3 (.CK( clk ) , .Q( u2_L11_3 ) , .D( u2_R10_3 ) );
  DFF_X1 u2_L11_reg_30 (.CK( clk ) , .Q( u2_L11_30 ) , .D( u2_R10_30 ) );
  DFF_X1 u2_L11_reg_31 (.CK( clk ) , .Q( u2_L11_31 ) , .D( u2_R10_31 ) );
  DFF_X1 u2_L11_reg_32 (.CK( clk ) , .Q( u2_L11_32 ) , .D( u2_R10_32 ) );
  DFF_X1 u2_L11_reg_4 (.CK( clk ) , .Q( u2_L11_4 ) , .D( u2_R10_4 ) );
  DFF_X1 u2_L11_reg_5 (.CK( clk ) , .Q( u2_L11_5 ) , .D( u2_R10_5 ) );
  DFF_X1 u2_L11_reg_6 (.CK( clk ) , .Q( u2_L11_6 ) , .D( u2_R10_6 ) );
  DFF_X1 u2_L11_reg_7 (.CK( clk ) , .Q( u2_L11_7 ) , .D( u2_R10_7 ) );
  DFF_X1 u2_L11_reg_8 (.CK( clk ) , .Q( u2_L11_8 ) , .D( u2_R10_8 ) );
  DFF_X1 u2_L11_reg_9 (.CK( clk ) , .Q( u2_L11_9 ) , .D( u2_R10_9 ) );
  DFF_X1 u2_L12_reg_1 (.CK( clk ) , .Q( u2_L12_1 ) , .D( u2_R11_1 ) );
  DFF_X1 u2_L12_reg_10 (.CK( clk ) , .Q( u2_L12_10 ) , .D( u2_R11_10 ) );
  DFF_X1 u2_L12_reg_11 (.CK( clk ) , .Q( u2_L12_11 ) , .D( u2_R11_11 ) );
  DFF_X1 u2_L12_reg_12 (.CK( clk ) , .Q( u2_L12_12 ) , .D( u2_R11_12 ) );
  DFF_X1 u2_L12_reg_13 (.CK( clk ) , .Q( u2_L12_13 ) , .D( u2_R11_13 ) );
  DFF_X1 u2_L12_reg_14 (.CK( clk ) , .Q( u2_L12_14 ) , .D( u2_R11_14 ) );
  DFF_X1 u2_L12_reg_15 (.CK( clk ) , .Q( u2_L12_15 ) , .D( u2_R11_15 ) );
  DFF_X1 u2_L12_reg_16 (.CK( clk ) , .Q( u2_L12_16 ) , .D( u2_R11_16 ) );
  DFF_X1 u2_L12_reg_17 (.CK( clk ) , .Q( u2_L12_17 ) , .D( u2_R11_17 ) );
  DFF_X1 u2_L12_reg_18 (.CK( clk ) , .Q( u2_L12_18 ) , .D( u2_R11_18 ) );
  DFF_X1 u2_L12_reg_19 (.CK( clk ) , .Q( u2_L12_19 ) , .D( u2_R11_19 ) );
  DFF_X1 u2_L12_reg_2 (.CK( clk ) , .Q( u2_L12_2 ) , .D( u2_R11_2 ) );
  DFF_X1 u2_L12_reg_20 (.CK( clk ) , .Q( u2_L12_20 ) , .D( u2_R11_20 ) );
  DFF_X1 u2_L12_reg_21 (.CK( clk ) , .Q( u2_L12_21 ) , .D( u2_R11_21 ) );
  DFF_X1 u2_L12_reg_22 (.CK( clk ) , .Q( u2_L12_22 ) , .D( u2_R11_22 ) );
  DFF_X1 u2_L12_reg_23 (.CK( clk ) , .Q( u2_L12_23 ) , .D( u2_R11_23 ) );
  DFF_X1 u2_L12_reg_24 (.CK( clk ) , .Q( u2_L12_24 ) , .D( u2_R11_24 ) );
  DFF_X1 u2_L12_reg_25 (.CK( clk ) , .Q( u2_L12_25 ) , .D( u2_R11_25 ) );
  DFF_X1 u2_L12_reg_26 (.CK( clk ) , .Q( u2_L12_26 ) , .D( u2_R11_26 ) );
  DFF_X1 u2_L12_reg_27 (.CK( clk ) , .Q( u2_L12_27 ) , .D( u2_R11_27 ) );
  DFF_X1 u2_L12_reg_28 (.CK( clk ) , .Q( u2_L12_28 ) , .D( u2_R11_28 ) );
  DFF_X1 u2_L12_reg_29 (.CK( clk ) , .Q( u2_L12_29 ) , .D( u2_R11_29 ) );
  DFF_X1 u2_L12_reg_3 (.CK( clk ) , .Q( u2_L12_3 ) , .D( u2_R11_3 ) );
  DFF_X1 u2_L12_reg_30 (.CK( clk ) , .Q( u2_L12_30 ) , .D( u2_R11_30 ) );
  DFF_X1 u2_L12_reg_31 (.CK( clk ) , .Q( u2_L12_31 ) , .D( u2_R11_31 ) );
  DFF_X1 u2_L12_reg_32 (.CK( clk ) , .Q( u2_L12_32 ) , .D( u2_R11_32 ) );
  DFF_X1 u2_L12_reg_4 (.CK( clk ) , .Q( u2_L12_4 ) , .D( u2_R11_4 ) );
  DFF_X1 u2_L12_reg_5 (.CK( clk ) , .Q( u2_L12_5 ) , .D( u2_R11_5 ) );
  DFF_X1 u2_L12_reg_6 (.CK( clk ) , .Q( u2_L12_6 ) , .D( u2_R11_6 ) );
  DFF_X1 u2_L12_reg_7 (.CK( clk ) , .Q( u2_L12_7 ) , .D( u2_R11_7 ) );
  DFF_X1 u2_L12_reg_8 (.CK( clk ) , .Q( u2_L12_8 ) , .D( u2_R11_8 ) );
  DFF_X1 u2_L12_reg_9 (.CK( clk ) , .Q( u2_L12_9 ) , .D( u2_R11_9 ) );
  DFF_X1 u2_L13_reg_1 (.CK( clk ) , .Q( u2_L13_1 ) , .D( u2_R12_1 ) );
  DFF_X1 u2_L13_reg_10 (.CK( clk ) , .Q( u2_L13_10 ) , .D( u2_R12_10 ) );
  DFF_X1 u2_L13_reg_11 (.CK( clk ) , .Q( u2_L13_11 ) , .D( u2_R12_11 ) );
  DFF_X1 u2_L13_reg_12 (.CK( clk ) , .Q( u2_L13_12 ) , .D( u2_R12_12 ) );
  DFF_X1 u2_L13_reg_13 (.CK( clk ) , .Q( u2_L13_13 ) , .D( u2_R12_13 ) );
  DFF_X1 u2_L13_reg_14 (.CK( clk ) , .Q( u2_L13_14 ) , .D( u2_R12_14 ) );
  DFF_X1 u2_L13_reg_15 (.CK( clk ) , .Q( u2_L13_15 ) , .D( u2_R12_15 ) );
  DFF_X1 u2_L13_reg_16 (.CK( clk ) , .Q( u2_L13_16 ) , .D( u2_R12_16 ) );
  DFF_X1 u2_L13_reg_17 (.CK( clk ) , .Q( u2_L13_17 ) , .D( u2_R12_17 ) );
  DFF_X1 u2_L13_reg_18 (.CK( clk ) , .Q( u2_L13_18 ) , .D( u2_R12_18 ) );
  DFF_X1 u2_L13_reg_19 (.CK( clk ) , .Q( u2_L13_19 ) , .D( u2_R12_19 ) );
  DFF_X1 u2_L13_reg_2 (.CK( clk ) , .Q( u2_L13_2 ) , .D( u2_R12_2 ) );
  DFF_X1 u2_L13_reg_20 (.CK( clk ) , .Q( u2_L13_20 ) , .D( u2_R12_20 ) );
  DFF_X1 u2_L13_reg_21 (.CK( clk ) , .Q( u2_L13_21 ) , .D( u2_R12_21 ) );
  DFF_X1 u2_L13_reg_22 (.CK( clk ) , .Q( u2_L13_22 ) , .D( u2_R12_22 ) );
  DFF_X1 u2_L13_reg_23 (.CK( clk ) , .Q( u2_L13_23 ) , .D( u2_R12_23 ) );
  DFF_X1 u2_L13_reg_24 (.CK( clk ) , .Q( u2_L13_24 ) , .D( u2_R12_24 ) );
  DFF_X1 u2_L13_reg_25 (.CK( clk ) , .Q( u2_L13_25 ) , .D( u2_R12_25 ) );
  DFF_X1 u2_L13_reg_26 (.CK( clk ) , .Q( u2_L13_26 ) , .D( u2_R12_26 ) );
  DFF_X1 u2_L13_reg_27 (.CK( clk ) , .Q( u2_L13_27 ) , .D( u2_R12_27 ) );
  DFF_X1 u2_L13_reg_28 (.CK( clk ) , .Q( u2_L13_28 ) , .D( u2_R12_28 ) );
  DFF_X1 u2_L13_reg_29 (.CK( clk ) , .Q( u2_L13_29 ) , .D( u2_R12_29 ) );
  DFF_X1 u2_L13_reg_3 (.CK( clk ) , .Q( u2_L13_3 ) , .D( u2_R12_3 ) );
  DFF_X1 u2_L13_reg_30 (.CK( clk ) , .Q( u2_L13_30 ) , .D( u2_R12_30 ) );
  DFF_X1 u2_L13_reg_31 (.CK( clk ) , .Q( u2_L13_31 ) , .D( u2_R12_31 ) );
  DFF_X1 u2_L13_reg_32 (.CK( clk ) , .Q( u2_L13_32 ) , .D( u2_R12_32 ) );
  DFF_X1 u2_L13_reg_4 (.CK( clk ) , .Q( u2_L13_4 ) , .D( u2_R12_4 ) );
  DFF_X1 u2_L13_reg_5 (.CK( clk ) , .Q( u2_L13_5 ) , .D( u2_R12_5 ) );
  DFF_X1 u2_L13_reg_6 (.CK( clk ) , .Q( u2_L13_6 ) , .D( u2_R12_6 ) );
  DFF_X1 u2_L13_reg_7 (.CK( clk ) , .Q( u2_L13_7 ) , .D( u2_R12_7 ) );
  DFF_X1 u2_L13_reg_8 (.CK( clk ) , .Q( u2_L13_8 ) , .D( u2_R12_8 ) );
  DFF_X1 u2_L13_reg_9 (.CK( clk ) , .Q( u2_L13_9 ) , .D( u2_R12_9 ) );
  DFF_X1 u2_L14_reg_1 (.CK( clk ) , .Q( u2_L14_1 ) , .D( u2_R13_1 ) );
  DFF_X1 u2_L14_reg_10 (.CK( clk ) , .Q( u2_L14_10 ) , .D( u2_R13_10 ) );
  DFF_X1 u2_L14_reg_11 (.CK( clk ) , .Q( u2_L14_11 ) , .D( u2_R13_11 ) );
  DFF_X1 u2_L14_reg_12 (.CK( clk ) , .Q( u2_L14_12 ) , .D( u2_R13_12 ) );
  DFF_X1 u2_L14_reg_13 (.CK( clk ) , .Q( u2_L14_13 ) , .D( u2_R13_13 ) );
  DFF_X1 u2_L14_reg_14 (.CK( clk ) , .Q( u2_L14_14 ) , .D( u2_R13_14 ) );
  DFF_X1 u2_L14_reg_15 (.CK( clk ) , .Q( u2_L14_15 ) , .D( u2_R13_15 ) );
  DFF_X1 u2_L14_reg_16 (.CK( clk ) , .Q( u2_L14_16 ) , .D( u2_R13_16 ) );
  DFF_X1 u2_L14_reg_17 (.CK( clk ) , .Q( u2_L14_17 ) , .D( u2_R13_17 ) );
  DFF_X1 u2_L14_reg_18 (.CK( clk ) , .Q( u2_L14_18 ) , .D( u2_R13_18 ) );
  DFF_X1 u2_L14_reg_19 (.CK( clk ) , .Q( u2_L14_19 ) , .D( u2_R13_19 ) );
  DFF_X1 u2_L14_reg_2 (.CK( clk ) , .Q( u2_L14_2 ) , .D( u2_R13_2 ) );
  DFF_X1 u2_L14_reg_20 (.CK( clk ) , .Q( u2_L14_20 ) , .D( u2_R13_20 ) );
  DFF_X1 u2_L14_reg_21 (.CK( clk ) , .Q( u2_L14_21 ) , .D( u2_R13_21 ) );
  DFF_X1 u2_L14_reg_22 (.CK( clk ) , .Q( u2_L14_22 ) , .D( u2_R13_22 ) );
  DFF_X1 u2_L14_reg_23 (.CK( clk ) , .Q( u2_L14_23 ) , .D( u2_R13_23 ) );
  DFF_X1 u2_L14_reg_24 (.CK( clk ) , .Q( u2_L14_24 ) , .D( u2_R13_24 ) );
  DFF_X1 u2_L14_reg_25 (.CK( clk ) , .Q( u2_L14_25 ) , .D( u2_R13_25 ) );
  DFF_X1 u2_L14_reg_26 (.CK( clk ) , .Q( u2_L14_26 ) , .D( u2_R13_26 ) );
  DFF_X1 u2_L14_reg_27 (.CK( clk ) , .Q( u2_L14_27 ) , .D( u2_R13_27 ) );
  DFF_X1 u2_L14_reg_28 (.CK( clk ) , .Q( u2_L14_28 ) , .D( u2_R13_28 ) );
  DFF_X1 u2_L14_reg_29 (.CK( clk ) , .Q( u2_L14_29 ) , .D( u2_R13_29 ) );
  DFF_X1 u2_L14_reg_3 (.CK( clk ) , .Q( u2_L14_3 ) , .D( u2_R13_3 ) );
  DFF_X1 u2_L14_reg_30 (.CK( clk ) , .Q( u2_L14_30 ) , .D( u2_R13_30 ) );
  DFF_X1 u2_L14_reg_31 (.CK( clk ) , .Q( u2_L14_31 ) , .D( u2_R13_31 ) );
  DFF_X1 u2_L14_reg_32 (.CK( clk ) , .Q( u2_L14_32 ) , .D( u2_R13_32 ) );
  DFF_X1 u2_L14_reg_4 (.CK( clk ) , .Q( u2_L14_4 ) , .D( u2_R13_4 ) );
  DFF_X1 u2_L14_reg_5 (.CK( clk ) , .Q( u2_L14_5 ) , .D( u2_R13_5 ) );
  DFF_X1 u2_L14_reg_6 (.CK( clk ) , .Q( u2_L14_6 ) , .D( u2_R13_6 ) );
  DFF_X1 u2_L14_reg_7 (.CK( clk ) , .Q( u2_L14_7 ) , .D( u2_R13_7 ) );
  DFF_X1 u2_L14_reg_8 (.CK( clk ) , .Q( u2_L14_8 ) , .D( u2_R13_8 ) );
  DFF_X1 u2_L14_reg_9 (.CK( clk ) , .Q( u2_L14_9 ) , .D( u2_R13_9 ) );
  DFF_X1 u2_L1_reg_1 (.CK( clk ) , .Q( u2_L1_1 ) , .D( u2_R0_1 ) );
  DFF_X1 u2_L1_reg_10 (.CK( clk ) , .Q( u2_L1_10 ) , .D( u2_R0_10 ) );
  DFF_X1 u2_L1_reg_11 (.CK( clk ) , .Q( u2_L1_11 ) , .D( u2_R0_11 ) );
  DFF_X1 u2_L1_reg_12 (.CK( clk ) , .Q( u2_L1_12 ) , .D( u2_R0_12 ) );
  DFF_X1 u2_L1_reg_13 (.CK( clk ) , .Q( u2_L1_13 ) , .D( u2_R0_13 ) );
  DFF_X1 u2_L1_reg_14 (.CK( clk ) , .Q( u2_L1_14 ) , .D( u2_R0_14 ) );
  DFF_X1 u2_L1_reg_15 (.CK( clk ) , .Q( u2_L1_15 ) , .D( u2_R0_15 ) );
  DFF_X1 u2_L1_reg_16 (.CK( clk ) , .Q( u2_L1_16 ) , .D( u2_R0_16 ) );
  DFF_X1 u2_L1_reg_17 (.CK( clk ) , .Q( u2_L1_17 ) , .D( u2_R0_17 ) );
  DFF_X1 u2_L1_reg_18 (.CK( clk ) , .Q( u2_L1_18 ) , .D( u2_R0_18 ) );
  DFF_X1 u2_L1_reg_19 (.CK( clk ) , .Q( u2_L1_19 ) , .D( u2_R0_19 ) );
  DFF_X1 u2_L1_reg_2 (.CK( clk ) , .Q( u2_L1_2 ) , .D( u2_R0_2 ) );
  DFF_X1 u2_L1_reg_20 (.CK( clk ) , .Q( u2_L1_20 ) , .D( u2_R0_20 ) );
  DFF_X1 u2_L1_reg_21 (.CK( clk ) , .Q( u2_L1_21 ) , .D( u2_R0_21 ) );
  DFF_X1 u2_L1_reg_22 (.CK( clk ) , .Q( u2_L1_22 ) , .D( u2_R0_22 ) );
  DFF_X1 u2_L1_reg_23 (.CK( clk ) , .Q( u2_L1_23 ) , .D( u2_R0_23 ) );
  DFF_X1 u2_L1_reg_24 (.CK( clk ) , .Q( u2_L1_24 ) , .D( u2_R0_24 ) );
  DFF_X1 u2_L1_reg_25 (.CK( clk ) , .Q( u2_L1_25 ) , .D( u2_R0_25 ) );
  DFF_X1 u2_L1_reg_26 (.CK( clk ) , .Q( u2_L1_26 ) , .D( u2_R0_26 ) );
  DFF_X1 u2_L1_reg_27 (.CK( clk ) , .Q( u2_L1_27 ) , .D( u2_R0_27 ) );
  DFF_X1 u2_L1_reg_28 (.CK( clk ) , .Q( u2_L1_28 ) , .D( u2_R0_28 ) );
  DFF_X1 u2_L1_reg_29 (.CK( clk ) , .Q( u2_L1_29 ) , .D( u2_R0_29 ) );
  DFF_X1 u2_L1_reg_3 (.CK( clk ) , .Q( u2_L1_3 ) , .D( u2_R0_3 ) );
  DFF_X1 u2_L1_reg_30 (.CK( clk ) , .Q( u2_L1_30 ) , .D( u2_R0_30 ) );
  DFF_X1 u2_L1_reg_31 (.CK( clk ) , .Q( u2_L1_31 ) , .D( u2_R0_31 ) );
  DFF_X1 u2_L1_reg_32 (.CK( clk ) , .Q( u2_L1_32 ) , .D( u2_R0_32 ) );
  DFF_X1 u2_L1_reg_4 (.CK( clk ) , .Q( u2_L1_4 ) , .D( u2_R0_4 ) );
  DFF_X1 u2_L1_reg_5 (.CK( clk ) , .Q( u2_L1_5 ) , .D( u2_R0_5 ) );
  DFF_X1 u2_L1_reg_6 (.CK( clk ) , .Q( u2_L1_6 ) , .D( u2_R0_6 ) );
  DFF_X1 u2_L1_reg_7 (.CK( clk ) , .Q( u2_L1_7 ) , .D( u2_R0_7 ) );
  DFF_X1 u2_L1_reg_8 (.CK( clk ) , .Q( u2_L1_8 ) , .D( u2_R0_8 ) );
  DFF_X1 u2_L1_reg_9 (.CK( clk ) , .Q( u2_L1_9 ) , .D( u2_R0_9 ) );
  DFF_X1 u2_L2_reg_1 (.CK( clk ) , .Q( u2_L2_1 ) , .D( u2_R1_1 ) );
  DFF_X1 u2_L2_reg_10 (.CK( clk ) , .Q( u2_L2_10 ) , .D( u2_R1_10 ) );
  DFF_X1 u2_L2_reg_11 (.CK( clk ) , .Q( u2_L2_11 ) , .D( u2_R1_11 ) );
  DFF_X1 u2_L2_reg_12 (.CK( clk ) , .Q( u2_L2_12 ) , .D( u2_R1_12 ) );
  DFF_X1 u2_L2_reg_13 (.CK( clk ) , .Q( u2_L2_13 ) , .D( u2_R1_13 ) );
  DFF_X1 u2_L2_reg_14 (.CK( clk ) , .Q( u2_L2_14 ) , .D( u2_R1_14 ) );
  DFF_X1 u2_L2_reg_15 (.CK( clk ) , .Q( u2_L2_15 ) , .D( u2_R1_15 ) );
  DFF_X1 u2_L2_reg_16 (.CK( clk ) , .Q( u2_L2_16 ) , .D( u2_R1_16 ) );
  DFF_X1 u2_L2_reg_17 (.CK( clk ) , .Q( u2_L2_17 ) , .D( u2_R1_17 ) );
  DFF_X1 u2_L2_reg_18 (.CK( clk ) , .Q( u2_L2_18 ) , .D( u2_R1_18 ) );
  DFF_X1 u2_L2_reg_19 (.CK( clk ) , .Q( u2_L2_19 ) , .D( u2_R1_19 ) );
  DFF_X1 u2_L2_reg_2 (.CK( clk ) , .Q( u2_L2_2 ) , .D( u2_R1_2 ) );
  DFF_X1 u2_L2_reg_20 (.CK( clk ) , .Q( u2_L2_20 ) , .D( u2_R1_20 ) );
  DFF_X1 u2_L2_reg_21 (.CK( clk ) , .Q( u2_L2_21 ) , .D( u2_R1_21 ) );
  DFF_X1 u2_L2_reg_22 (.CK( clk ) , .Q( u2_L2_22 ) , .D( u2_R1_22 ) );
  DFF_X1 u2_L2_reg_23 (.CK( clk ) , .Q( u2_L2_23 ) , .D( u2_R1_23 ) );
  DFF_X1 u2_L2_reg_24 (.CK( clk ) , .Q( u2_L2_24 ) , .D( u2_R1_24 ) );
  DFF_X1 u2_L2_reg_25 (.CK( clk ) , .Q( u2_L2_25 ) , .D( u2_R1_25 ) );
  DFF_X1 u2_L2_reg_26 (.CK( clk ) , .Q( u2_L2_26 ) , .D( u2_R1_26 ) );
  DFF_X1 u2_L2_reg_27 (.CK( clk ) , .Q( u2_L2_27 ) , .D( u2_R1_27 ) );
  DFF_X1 u2_L2_reg_28 (.CK( clk ) , .Q( u2_L2_28 ) , .D( u2_R1_28 ) );
  DFF_X1 u2_L2_reg_29 (.CK( clk ) , .Q( u2_L2_29 ) , .D( u2_R1_29 ) );
  DFF_X1 u2_L2_reg_3 (.CK( clk ) , .Q( u2_L2_3 ) , .D( u2_R1_3 ) );
  DFF_X1 u2_L2_reg_30 (.CK( clk ) , .Q( u2_L2_30 ) , .D( u2_R1_30 ) );
  DFF_X1 u2_L2_reg_31 (.CK( clk ) , .Q( u2_L2_31 ) , .D( u2_R1_31 ) );
  DFF_X1 u2_L2_reg_32 (.CK( clk ) , .Q( u2_L2_32 ) , .D( u2_R1_32 ) );
  DFF_X1 u2_L2_reg_4 (.CK( clk ) , .Q( u2_L2_4 ) , .D( u2_R1_4 ) );
  DFF_X1 u2_L2_reg_5 (.CK( clk ) , .Q( u2_L2_5 ) , .D( u2_R1_5 ) );
  DFF_X1 u2_L2_reg_6 (.CK( clk ) , .Q( u2_L2_6 ) , .D( u2_R1_6 ) );
  DFF_X1 u2_L2_reg_7 (.CK( clk ) , .Q( u2_L2_7 ) , .D( u2_R1_7 ) );
  DFF_X1 u2_L2_reg_8 (.CK( clk ) , .Q( u2_L2_8 ) , .D( u2_R1_8 ) );
  DFF_X1 u2_L2_reg_9 (.CK( clk ) , .Q( u2_L2_9 ) , .D( u2_R1_9 ) );
  DFF_X1 u2_L3_reg_1 (.CK( clk ) , .Q( u2_L3_1 ) , .D( u2_R2_1 ) );
  DFF_X1 u2_L3_reg_10 (.CK( clk ) , .Q( u2_L3_10 ) , .D( u2_R2_10 ) );
  DFF_X1 u2_L3_reg_11 (.CK( clk ) , .Q( u2_L3_11 ) , .D( u2_R2_11 ) );
  DFF_X1 u2_L3_reg_12 (.CK( clk ) , .Q( u2_L3_12 ) , .D( u2_R2_12 ) );
  DFF_X1 u2_L3_reg_13 (.CK( clk ) , .Q( u2_L3_13 ) , .D( u2_R2_13 ) );
  DFF_X1 u2_L3_reg_14 (.CK( clk ) , .Q( u2_L3_14 ) , .D( u2_R2_14 ) );
  DFF_X1 u2_L3_reg_15 (.CK( clk ) , .Q( u2_L3_15 ) , .D( u2_R2_15 ) );
  DFF_X1 u2_L3_reg_16 (.CK( clk ) , .Q( u2_L3_16 ) , .D( u2_R2_16 ) );
  DFF_X1 u2_L3_reg_17 (.CK( clk ) , .Q( u2_L3_17 ) , .D( u2_R2_17 ) );
  DFF_X1 u2_L3_reg_18 (.CK( clk ) , .Q( u2_L3_18 ) , .D( u2_R2_18 ) );
  DFF_X1 u2_L3_reg_19 (.CK( clk ) , .Q( u2_L3_19 ) , .D( u2_R2_19 ) );
  DFF_X1 u2_L3_reg_2 (.CK( clk ) , .Q( u2_L3_2 ) , .D( u2_R2_2 ) );
  DFF_X1 u2_L3_reg_20 (.CK( clk ) , .Q( u2_L3_20 ) , .D( u2_R2_20 ) );
  DFF_X1 u2_L3_reg_21 (.CK( clk ) , .Q( u2_L3_21 ) , .D( u2_R2_21 ) );
  DFF_X1 u2_L3_reg_22 (.CK( clk ) , .Q( u2_L3_22 ) , .D( u2_R2_22 ) );
  DFF_X1 u2_L3_reg_23 (.CK( clk ) , .Q( u2_L3_23 ) , .D( u2_R2_23 ) );
  DFF_X1 u2_L3_reg_24 (.CK( clk ) , .Q( u2_L3_24 ) , .D( u2_R2_24 ) );
  DFF_X1 u2_L3_reg_25 (.CK( clk ) , .Q( u2_L3_25 ) , .D( u2_R2_25 ) );
  DFF_X1 u2_L3_reg_26 (.CK( clk ) , .Q( u2_L3_26 ) , .D( u2_R2_26 ) );
  DFF_X1 u2_L3_reg_27 (.CK( clk ) , .Q( u2_L3_27 ) , .D( u2_R2_27 ) );
  DFF_X1 u2_L3_reg_28 (.CK( clk ) , .Q( u2_L3_28 ) , .D( u2_R2_28 ) );
  DFF_X1 u2_L3_reg_29 (.CK( clk ) , .Q( u2_L3_29 ) , .D( u2_R2_29 ) );
  DFF_X1 u2_L3_reg_3 (.CK( clk ) , .Q( u2_L3_3 ) , .D( u2_R2_3 ) );
  DFF_X1 u2_L3_reg_30 (.CK( clk ) , .Q( u2_L3_30 ) , .D( u2_R2_30 ) );
  DFF_X1 u2_L3_reg_31 (.CK( clk ) , .Q( u2_L3_31 ) , .D( u2_R2_31 ) );
  DFF_X1 u2_L3_reg_32 (.CK( clk ) , .Q( u2_L3_32 ) , .D( u2_R2_32 ) );
  DFF_X1 u2_L3_reg_4 (.CK( clk ) , .Q( u2_L3_4 ) , .D( u2_R2_4 ) );
  DFF_X1 u2_L3_reg_5 (.CK( clk ) , .Q( u2_L3_5 ) , .D( u2_R2_5 ) );
  DFF_X1 u2_L3_reg_6 (.CK( clk ) , .Q( u2_L3_6 ) , .D( u2_R2_6 ) );
  DFF_X1 u2_L3_reg_7 (.CK( clk ) , .Q( u2_L3_7 ) , .D( u2_R2_7 ) );
  DFF_X1 u2_L3_reg_8 (.CK( clk ) , .Q( u2_L3_8 ) , .D( u2_R2_8 ) );
  DFF_X1 u2_L3_reg_9 (.CK( clk ) , .Q( u2_L3_9 ) , .D( u2_R2_9 ) );
  DFF_X1 u2_L4_reg_1 (.CK( clk ) , .Q( u2_L4_1 ) , .D( u2_R3_1 ) );
  DFF_X1 u2_L4_reg_10 (.CK( clk ) , .Q( u2_L4_10 ) , .D( u2_R3_10 ) );
  DFF_X1 u2_L4_reg_11 (.CK( clk ) , .Q( u2_L4_11 ) , .D( u2_R3_11 ) );
  DFF_X1 u2_L4_reg_12 (.CK( clk ) , .Q( u2_L4_12 ) , .D( u2_R3_12 ) );
  DFF_X1 u2_L4_reg_13 (.CK( clk ) , .Q( u2_L4_13 ) , .D( u2_R3_13 ) );
  DFF_X1 u2_L4_reg_14 (.CK( clk ) , .Q( u2_L4_14 ) , .D( u2_R3_14 ) );
  DFF_X1 u2_L4_reg_15 (.CK( clk ) , .Q( u2_L4_15 ) , .D( u2_R3_15 ) );
  DFF_X1 u2_L4_reg_16 (.CK( clk ) , .Q( u2_L4_16 ) , .D( u2_R3_16 ) );
  DFF_X1 u2_L4_reg_17 (.CK( clk ) , .Q( u2_L4_17 ) , .D( u2_R3_17 ) );
  DFF_X1 u2_L4_reg_18 (.CK( clk ) , .Q( u2_L4_18 ) , .D( u2_R3_18 ) );
  DFF_X1 u2_L4_reg_19 (.CK( clk ) , .Q( u2_L4_19 ) , .D( u2_R3_19 ) );
  DFF_X1 u2_L4_reg_2 (.CK( clk ) , .Q( u2_L4_2 ) , .D( u2_R3_2 ) );
  DFF_X1 u2_L4_reg_20 (.CK( clk ) , .Q( u2_L4_20 ) , .D( u2_R3_20 ) );
  DFF_X1 u2_L4_reg_21 (.CK( clk ) , .Q( u2_L4_21 ) , .D( u2_R3_21 ) );
  DFF_X1 u2_L4_reg_22 (.CK( clk ) , .Q( u2_L4_22 ) , .D( u2_R3_22 ) );
  DFF_X1 u2_L4_reg_23 (.CK( clk ) , .Q( u2_L4_23 ) , .D( u2_R3_23 ) );
  DFF_X1 u2_L4_reg_24 (.CK( clk ) , .Q( u2_L4_24 ) , .D( u2_R3_24 ) );
  DFF_X1 u2_L4_reg_25 (.CK( clk ) , .Q( u2_L4_25 ) , .D( u2_R3_25 ) );
  DFF_X1 u2_L4_reg_26 (.CK( clk ) , .Q( u2_L4_26 ) , .D( u2_R3_26 ) );
  DFF_X1 u2_L4_reg_27 (.CK( clk ) , .Q( u2_L4_27 ) , .D( u2_R3_27 ) );
  DFF_X1 u2_L4_reg_28 (.CK( clk ) , .Q( u2_L4_28 ) , .D( u2_R3_28 ) );
  DFF_X1 u2_L4_reg_29 (.CK( clk ) , .Q( u2_L4_29 ) , .D( u2_R3_29 ) );
  DFF_X1 u2_L4_reg_3 (.CK( clk ) , .Q( u2_L4_3 ) , .D( u2_R3_3 ) );
  DFF_X1 u2_L4_reg_30 (.CK( clk ) , .Q( u2_L4_30 ) , .D( u2_R3_30 ) );
  DFF_X1 u2_L4_reg_31 (.CK( clk ) , .Q( u2_L4_31 ) , .D( u2_R3_31 ) );
  DFF_X1 u2_L4_reg_32 (.CK( clk ) , .Q( u2_L4_32 ) , .D( u2_R3_32 ) );
  DFF_X1 u2_L4_reg_4 (.CK( clk ) , .Q( u2_L4_4 ) , .D( u2_R3_4 ) );
  DFF_X1 u2_L4_reg_5 (.CK( clk ) , .Q( u2_L4_5 ) , .D( u2_R3_5 ) );
  DFF_X1 u2_L4_reg_6 (.CK( clk ) , .Q( u2_L4_6 ) , .D( u2_R3_6 ) );
  DFF_X1 u2_L4_reg_7 (.CK( clk ) , .Q( u2_L4_7 ) , .D( u2_R3_7 ) );
  DFF_X1 u2_L4_reg_8 (.CK( clk ) , .Q( u2_L4_8 ) , .D( u2_R3_8 ) );
  DFF_X1 u2_L4_reg_9 (.CK( clk ) , .Q( u2_L4_9 ) , .D( u2_R3_9 ) );
  DFF_X1 u2_L5_reg_1 (.CK( clk ) , .Q( u2_L5_1 ) , .D( u2_R4_1 ) );
  DFF_X1 u2_L5_reg_10 (.CK( clk ) , .Q( u2_L5_10 ) , .D( u2_R4_10 ) );
  DFF_X1 u2_L5_reg_11 (.CK( clk ) , .Q( u2_L5_11 ) , .D( u2_R4_11 ) );
  DFF_X1 u2_L5_reg_12 (.CK( clk ) , .Q( u2_L5_12 ) , .D( u2_R4_12 ) );
  DFF_X1 u2_L5_reg_13 (.CK( clk ) , .Q( u2_L5_13 ) , .D( u2_R4_13 ) );
  DFF_X1 u2_L5_reg_14 (.CK( clk ) , .Q( u2_L5_14 ) , .D( u2_R4_14 ) );
  DFF_X1 u2_L5_reg_15 (.CK( clk ) , .Q( u2_L5_15 ) , .D( u2_R4_15 ) );
  DFF_X1 u2_L5_reg_16 (.CK( clk ) , .Q( u2_L5_16 ) , .D( u2_R4_16 ) );
  DFF_X1 u2_L5_reg_17 (.CK( clk ) , .Q( u2_L5_17 ) , .D( u2_R4_17 ) );
  DFF_X1 u2_L5_reg_18 (.CK( clk ) , .Q( u2_L5_18 ) , .D( u2_R4_18 ) );
  DFF_X1 u2_L5_reg_19 (.CK( clk ) , .Q( u2_L5_19 ) , .D( u2_R4_19 ) );
  DFF_X1 u2_L5_reg_2 (.CK( clk ) , .Q( u2_L5_2 ) , .D( u2_R4_2 ) );
  DFF_X1 u2_L5_reg_20 (.CK( clk ) , .Q( u2_L5_20 ) , .D( u2_R4_20 ) );
  DFF_X1 u2_L5_reg_21 (.CK( clk ) , .Q( u2_L5_21 ) , .D( u2_R4_21 ) );
  DFF_X1 u2_L5_reg_22 (.CK( clk ) , .Q( u2_L5_22 ) , .D( u2_R4_22 ) );
  DFF_X1 u2_L5_reg_23 (.CK( clk ) , .Q( u2_L5_23 ) , .D( u2_R4_23 ) );
  DFF_X1 u2_L5_reg_24 (.CK( clk ) , .Q( u2_L5_24 ) , .D( u2_R4_24 ) );
  DFF_X1 u2_L5_reg_25 (.CK( clk ) , .Q( u2_L5_25 ) , .D( u2_R4_25 ) );
  DFF_X1 u2_L5_reg_26 (.CK( clk ) , .Q( u2_L5_26 ) , .D( u2_R4_26 ) );
  DFF_X1 u2_L5_reg_27 (.CK( clk ) , .Q( u2_L5_27 ) , .D( u2_R4_27 ) );
  DFF_X1 u2_L5_reg_28 (.CK( clk ) , .Q( u2_L5_28 ) , .D( u2_R4_28 ) );
  DFF_X1 u2_L5_reg_29 (.CK( clk ) , .Q( u2_L5_29 ) , .D( u2_R4_29 ) );
  DFF_X1 u2_L5_reg_3 (.CK( clk ) , .Q( u2_L5_3 ) , .D( u2_R4_3 ) );
  DFF_X1 u2_L5_reg_30 (.CK( clk ) , .Q( u2_L5_30 ) , .D( u2_R4_30 ) );
  DFF_X1 u2_L5_reg_31 (.CK( clk ) , .Q( u2_L5_31 ) , .D( u2_R4_31 ) );
  DFF_X1 u2_L5_reg_32 (.CK( clk ) , .Q( u2_L5_32 ) , .D( u2_R4_32 ) );
  DFF_X1 u2_L5_reg_4 (.CK( clk ) , .Q( u2_L5_4 ) , .D( u2_R4_4 ) );
  DFF_X1 u2_L5_reg_5 (.CK( clk ) , .Q( u2_L5_5 ) , .D( u2_R4_5 ) );
  DFF_X1 u2_L5_reg_6 (.CK( clk ) , .Q( u2_L5_6 ) , .D( u2_R4_6 ) );
  DFF_X1 u2_L5_reg_7 (.CK( clk ) , .Q( u2_L5_7 ) , .D( u2_R4_7 ) );
  DFF_X1 u2_L5_reg_8 (.CK( clk ) , .Q( u2_L5_8 ) , .D( u2_R4_8 ) );
  DFF_X1 u2_L5_reg_9 (.CK( clk ) , .Q( u2_L5_9 ) , .D( u2_R4_9 ) );
  DFF_X1 u2_L6_reg_1 (.CK( clk ) , .Q( u2_L6_1 ) , .D( u2_R5_1 ) );
  DFF_X1 u2_L6_reg_10 (.CK( clk ) , .Q( u2_L6_10 ) , .D( u2_R5_10 ) );
  DFF_X1 u2_L6_reg_11 (.CK( clk ) , .Q( u2_L6_11 ) , .D( u2_R5_11 ) );
  DFF_X1 u2_L6_reg_12 (.CK( clk ) , .Q( u2_L6_12 ) , .D( u2_R5_12 ) );
  DFF_X1 u2_L6_reg_13 (.CK( clk ) , .Q( u2_L6_13 ) , .D( u2_R5_13 ) );
  DFF_X1 u2_L6_reg_14 (.CK( clk ) , .Q( u2_L6_14 ) , .D( u2_R5_14 ) );
  DFF_X1 u2_L6_reg_15 (.CK( clk ) , .Q( u2_L6_15 ) , .D( u2_R5_15 ) );
  DFF_X1 u2_L6_reg_16 (.CK( clk ) , .Q( u2_L6_16 ) , .D( u2_R5_16 ) );
  DFF_X1 u2_L6_reg_17 (.CK( clk ) , .Q( u2_L6_17 ) , .D( u2_R5_17 ) );
  DFF_X1 u2_L6_reg_18 (.CK( clk ) , .Q( u2_L6_18 ) , .D( u2_R5_18 ) );
  DFF_X1 u2_L6_reg_19 (.CK( clk ) , .Q( u2_L6_19 ) , .D( u2_R5_19 ) );
  DFF_X1 u2_L6_reg_2 (.CK( clk ) , .Q( u2_L6_2 ) , .D( u2_R5_2 ) );
  DFF_X1 u2_L6_reg_20 (.CK( clk ) , .Q( u2_L6_20 ) , .D( u2_R5_20 ) );
  DFF_X1 u2_L6_reg_21 (.CK( clk ) , .Q( u2_L6_21 ) , .D( u2_R5_21 ) );
  DFF_X1 u2_L6_reg_22 (.CK( clk ) , .Q( u2_L6_22 ) , .D( u2_R5_22 ) );
  DFF_X1 u2_L6_reg_23 (.CK( clk ) , .Q( u2_L6_23 ) , .D( u2_R5_23 ) );
  DFF_X1 u2_L6_reg_24 (.CK( clk ) , .Q( u2_L6_24 ) , .D( u2_R5_24 ) );
  DFF_X1 u2_L6_reg_25 (.CK( clk ) , .Q( u2_L6_25 ) , .D( u2_R5_25 ) );
  DFF_X1 u2_L6_reg_26 (.CK( clk ) , .Q( u2_L6_26 ) , .D( u2_R5_26 ) );
  DFF_X1 u2_L6_reg_27 (.CK( clk ) , .Q( u2_L6_27 ) , .D( u2_R5_27 ) );
  DFF_X1 u2_L6_reg_28 (.CK( clk ) , .Q( u2_L6_28 ) , .D( u2_R5_28 ) );
  DFF_X1 u2_L6_reg_29 (.CK( clk ) , .Q( u2_L6_29 ) , .D( u2_R5_29 ) );
  DFF_X1 u2_L6_reg_3 (.CK( clk ) , .Q( u2_L6_3 ) , .D( u2_R5_3 ) );
  DFF_X1 u2_L6_reg_30 (.CK( clk ) , .Q( u2_L6_30 ) , .D( u2_R5_30 ) );
  DFF_X1 u2_L6_reg_31 (.CK( clk ) , .Q( u2_L6_31 ) , .D( u2_R5_31 ) );
  DFF_X1 u2_L6_reg_32 (.CK( clk ) , .Q( u2_L6_32 ) , .D( u2_R5_32 ) );
  DFF_X1 u2_L6_reg_4 (.CK( clk ) , .Q( u2_L6_4 ) , .D( u2_R5_4 ) );
  DFF_X1 u2_L6_reg_5 (.CK( clk ) , .Q( u2_L6_5 ) , .D( u2_R5_5 ) );
  DFF_X1 u2_L6_reg_6 (.CK( clk ) , .Q( u2_L6_6 ) , .D( u2_R5_6 ) );
  DFF_X1 u2_L6_reg_7 (.CK( clk ) , .Q( u2_L6_7 ) , .D( u2_R5_7 ) );
  DFF_X1 u2_L6_reg_8 (.CK( clk ) , .Q( u2_L6_8 ) , .D( u2_R5_8 ) );
  DFF_X1 u2_L6_reg_9 (.CK( clk ) , .Q( u2_L6_9 ) , .D( u2_R5_9 ) );
  DFF_X1 u2_L7_reg_1 (.CK( clk ) , .Q( u2_L7_1 ) , .D( u2_R6_1 ) );
  DFF_X1 u2_L7_reg_10 (.CK( clk ) , .Q( u2_L7_10 ) , .D( u2_R6_10 ) );
  DFF_X1 u2_L7_reg_11 (.CK( clk ) , .Q( u2_L7_11 ) , .D( u2_R6_11 ) );
  DFF_X1 u2_L7_reg_12 (.CK( clk ) , .Q( u2_L7_12 ) , .D( u2_R6_12 ) );
  DFF_X1 u2_L7_reg_13 (.CK( clk ) , .Q( u2_L7_13 ) , .D( u2_R6_13 ) );
  DFF_X1 u2_L7_reg_14 (.CK( clk ) , .Q( u2_L7_14 ) , .D( u2_R6_14 ) );
  DFF_X1 u2_L7_reg_15 (.CK( clk ) , .Q( u2_L7_15 ) , .D( u2_R6_15 ) );
  DFF_X1 u2_L7_reg_16 (.CK( clk ) , .Q( u2_L7_16 ) , .D( u2_R6_16 ) );
  DFF_X1 u2_L7_reg_17 (.CK( clk ) , .Q( u2_L7_17 ) , .D( u2_R6_17 ) );
  DFF_X1 u2_L7_reg_18 (.CK( clk ) , .Q( u2_L7_18 ) , .D( u2_R6_18 ) );
  DFF_X1 u2_L7_reg_19 (.CK( clk ) , .Q( u2_L7_19 ) , .D( u2_R6_19 ) );
  DFF_X1 u2_L7_reg_2 (.CK( clk ) , .Q( u2_L7_2 ) , .D( u2_R6_2 ) );
  DFF_X1 u2_L7_reg_20 (.CK( clk ) , .Q( u2_L7_20 ) , .D( u2_R6_20 ) );
  DFF_X1 u2_L7_reg_21 (.CK( clk ) , .Q( u2_L7_21 ) , .D( u2_R6_21 ) );
  DFF_X1 u2_L7_reg_22 (.CK( clk ) , .Q( u2_L7_22 ) , .D( u2_R6_22 ) );
  DFF_X1 u2_L7_reg_23 (.CK( clk ) , .Q( u2_L7_23 ) , .D( u2_R6_23 ) );
  DFF_X1 u2_L7_reg_24 (.CK( clk ) , .Q( u2_L7_24 ) , .D( u2_R6_24 ) );
  DFF_X1 u2_L7_reg_25 (.CK( clk ) , .Q( u2_L7_25 ) , .D( u2_R6_25 ) );
  DFF_X1 u2_L7_reg_26 (.CK( clk ) , .Q( u2_L7_26 ) , .D( u2_R6_26 ) );
  DFF_X1 u2_L7_reg_27 (.CK( clk ) , .Q( u2_L7_27 ) , .D( u2_R6_27 ) );
  DFF_X1 u2_L7_reg_28 (.CK( clk ) , .Q( u2_L7_28 ) , .D( u2_R6_28 ) );
  DFF_X1 u2_L7_reg_29 (.CK( clk ) , .Q( u2_L7_29 ) , .D( u2_R6_29 ) );
  DFF_X1 u2_L7_reg_3 (.CK( clk ) , .Q( u2_L7_3 ) , .D( u2_R6_3 ) );
  DFF_X1 u2_L7_reg_30 (.CK( clk ) , .Q( u2_L7_30 ) , .D( u2_R6_30 ) );
  DFF_X1 u2_L7_reg_31 (.CK( clk ) , .Q( u2_L7_31 ) , .D( u2_R6_31 ) );
  DFF_X1 u2_L7_reg_32 (.CK( clk ) , .Q( u2_L7_32 ) , .D( u2_R6_32 ) );
  DFF_X1 u2_L7_reg_4 (.CK( clk ) , .Q( u2_L7_4 ) , .D( u2_R6_4 ) );
  DFF_X1 u2_L7_reg_5 (.CK( clk ) , .Q( u2_L7_5 ) , .D( u2_R6_5 ) );
  DFF_X1 u2_L7_reg_6 (.CK( clk ) , .Q( u2_L7_6 ) , .D( u2_R6_6 ) );
  DFF_X1 u2_L7_reg_7 (.CK( clk ) , .Q( u2_L7_7 ) , .D( u2_R6_7 ) );
  DFF_X1 u2_L7_reg_8 (.CK( clk ) , .Q( u2_L7_8 ) , .D( u2_R6_8 ) );
  DFF_X1 u2_L7_reg_9 (.CK( clk ) , .Q( u2_L7_9 ) , .D( u2_R6_9 ) );
  DFF_X1 u2_L8_reg_1 (.CK( clk ) , .Q( u2_L8_1 ) , .D( u2_R7_1 ) );
  DFF_X1 u2_L8_reg_10 (.CK( clk ) , .Q( u2_L8_10 ) , .D( u2_R7_10 ) );
  DFF_X1 u2_L8_reg_11 (.CK( clk ) , .Q( u2_L8_11 ) , .D( u2_R7_11 ) );
  DFF_X1 u2_L8_reg_12 (.CK( clk ) , .Q( u2_L8_12 ) , .D( u2_R7_12 ) );
  DFF_X1 u2_L8_reg_13 (.CK( clk ) , .Q( u2_L8_13 ) , .D( u2_R7_13 ) );
  DFF_X1 u2_L8_reg_14 (.CK( clk ) , .Q( u2_L8_14 ) , .D( u2_R7_14 ) );
  DFF_X1 u2_L8_reg_15 (.CK( clk ) , .Q( u2_L8_15 ) , .D( u2_R7_15 ) );
  DFF_X1 u2_L8_reg_16 (.CK( clk ) , .Q( u2_L8_16 ) , .D( u2_R7_16 ) );
  DFF_X1 u2_L8_reg_17 (.CK( clk ) , .Q( u2_L8_17 ) , .D( u2_R7_17 ) );
  DFF_X1 u2_L8_reg_18 (.CK( clk ) , .Q( u2_L8_18 ) , .D( u2_R7_18 ) );
  DFF_X1 u2_L8_reg_19 (.CK( clk ) , .Q( u2_L8_19 ) , .D( u2_R7_19 ) );
  DFF_X1 u2_L8_reg_2 (.CK( clk ) , .Q( u2_L8_2 ) , .D( u2_R7_2 ) );
  DFF_X1 u2_L8_reg_20 (.CK( clk ) , .Q( u2_L8_20 ) , .D( u2_R7_20 ) );
  DFF_X1 u2_L8_reg_21 (.CK( clk ) , .Q( u2_L8_21 ) , .D( u2_R7_21 ) );
  DFF_X1 u2_L8_reg_22 (.CK( clk ) , .Q( u2_L8_22 ) , .D( u2_R7_22 ) );
  DFF_X1 u2_L8_reg_23 (.CK( clk ) , .Q( u2_L8_23 ) , .D( u2_R7_23 ) );
  DFF_X1 u2_L8_reg_24 (.CK( clk ) , .Q( u2_L8_24 ) , .D( u2_R7_24 ) );
  DFF_X1 u2_L8_reg_25 (.CK( clk ) , .Q( u2_L8_25 ) , .D( u2_R7_25 ) );
  DFF_X1 u2_L8_reg_26 (.CK( clk ) , .Q( u2_L8_26 ) , .D( u2_R7_26 ) );
  DFF_X1 u2_L8_reg_27 (.CK( clk ) , .Q( u2_L8_27 ) , .D( u2_R7_27 ) );
  DFF_X1 u2_L8_reg_28 (.CK( clk ) , .Q( u2_L8_28 ) , .D( u2_R7_28 ) );
  DFF_X1 u2_L8_reg_29 (.CK( clk ) , .Q( u2_L8_29 ) , .D( u2_R7_29 ) );
  DFF_X1 u2_L8_reg_3 (.CK( clk ) , .Q( u2_L8_3 ) , .D( u2_R7_3 ) );
  DFF_X1 u2_L8_reg_30 (.CK( clk ) , .Q( u2_L8_30 ) , .D( u2_R7_30 ) );
  DFF_X1 u2_L8_reg_31 (.CK( clk ) , .Q( u2_L8_31 ) , .D( u2_R7_31 ) );
  DFF_X1 u2_L8_reg_32 (.CK( clk ) , .Q( u2_L8_32 ) , .D( u2_R7_32 ) );
  DFF_X1 u2_L8_reg_4 (.CK( clk ) , .Q( u2_L8_4 ) , .D( u2_R7_4 ) );
  DFF_X1 u2_L8_reg_5 (.CK( clk ) , .Q( u2_L8_5 ) , .D( u2_R7_5 ) );
  DFF_X1 u2_L8_reg_6 (.CK( clk ) , .Q( u2_L8_6 ) , .D( u2_R7_6 ) );
  DFF_X1 u2_L8_reg_7 (.CK( clk ) , .Q( u2_L8_7 ) , .D( u2_R7_7 ) );
  DFF_X1 u2_L8_reg_8 (.CK( clk ) , .Q( u2_L8_8 ) , .D( u2_R7_8 ) );
  DFF_X1 u2_L8_reg_9 (.CK( clk ) , .Q( u2_L8_9 ) , .D( u2_R7_9 ) );
  DFF_X1 u2_L9_reg_1 (.CK( clk ) , .Q( u2_L9_1 ) , .D( u2_R8_1 ) );
  DFF_X1 u2_L9_reg_10 (.CK( clk ) , .Q( u2_L9_10 ) , .D( u2_R8_10 ) );
  DFF_X1 u2_L9_reg_11 (.CK( clk ) , .Q( u2_L9_11 ) , .D( u2_R8_11 ) );
  DFF_X1 u2_L9_reg_12 (.CK( clk ) , .Q( u2_L9_12 ) , .D( u2_R8_12 ) );
  DFF_X1 u2_L9_reg_13 (.CK( clk ) , .Q( u2_L9_13 ) , .D( u2_R8_13 ) );
  DFF_X1 u2_L9_reg_14 (.CK( clk ) , .Q( u2_L9_14 ) , .D( u2_R8_14 ) );
  DFF_X1 u2_L9_reg_15 (.CK( clk ) , .Q( u2_L9_15 ) , .D( u2_R8_15 ) );
  DFF_X1 u2_L9_reg_16 (.CK( clk ) , .Q( u2_L9_16 ) , .D( u2_R8_16 ) );
  DFF_X1 u2_L9_reg_17 (.CK( clk ) , .Q( u2_L9_17 ) , .D( u2_R8_17 ) );
  DFF_X1 u2_L9_reg_18 (.CK( clk ) , .Q( u2_L9_18 ) , .D( u2_R8_18 ) );
  DFF_X1 u2_L9_reg_19 (.CK( clk ) , .Q( u2_L9_19 ) , .D( u2_R8_19 ) );
  DFF_X1 u2_L9_reg_2 (.CK( clk ) , .Q( u2_L9_2 ) , .D( u2_R8_2 ) );
  DFF_X1 u2_L9_reg_20 (.CK( clk ) , .Q( u2_L9_20 ) , .D( u2_R8_20 ) );
  DFF_X1 u2_L9_reg_21 (.CK( clk ) , .Q( u2_L9_21 ) , .D( u2_R8_21 ) );
  DFF_X1 u2_L9_reg_22 (.CK( clk ) , .Q( u2_L9_22 ) , .D( u2_R8_22 ) );
  DFF_X1 u2_L9_reg_23 (.CK( clk ) , .Q( u2_L9_23 ) , .D( u2_R8_23 ) );
  DFF_X1 u2_L9_reg_24 (.CK( clk ) , .Q( u2_L9_24 ) , .D( u2_R8_24 ) );
  DFF_X1 u2_L9_reg_25 (.CK( clk ) , .Q( u2_L9_25 ) , .D( u2_R8_25 ) );
  DFF_X1 u2_L9_reg_26 (.CK( clk ) , .Q( u2_L9_26 ) , .D( u2_R8_26 ) );
  DFF_X1 u2_L9_reg_27 (.CK( clk ) , .Q( u2_L9_27 ) , .D( u2_R8_27 ) );
  DFF_X1 u2_L9_reg_28 (.CK( clk ) , .Q( u2_L9_28 ) , .D( u2_R8_28 ) );
  DFF_X1 u2_L9_reg_29 (.CK( clk ) , .Q( u2_L9_29 ) , .D( u2_R8_29 ) );
  DFF_X1 u2_L9_reg_3 (.CK( clk ) , .Q( u2_L9_3 ) , .D( u2_R8_3 ) );
  DFF_X1 u2_L9_reg_30 (.CK( clk ) , .Q( u2_L9_30 ) , .D( u2_R8_30 ) );
  DFF_X1 u2_L9_reg_31 (.CK( clk ) , .Q( u2_L9_31 ) , .D( u2_R8_31 ) );
  DFF_X1 u2_L9_reg_32 (.CK( clk ) , .Q( u2_L9_32 ) , .D( u2_R8_32 ) );
  DFF_X1 u2_L9_reg_4 (.CK( clk ) , .Q( u2_L9_4 ) , .D( u2_R8_4 ) );
  DFF_X1 u2_L9_reg_5 (.CK( clk ) , .Q( u2_L9_5 ) , .D( u2_R8_5 ) );
  DFF_X1 u2_L9_reg_6 (.CK( clk ) , .Q( u2_L9_6 ) , .D( u2_R8_6 ) );
  DFF_X1 u2_L9_reg_7 (.CK( clk ) , .Q( u2_L9_7 ) , .D( u2_R8_7 ) );
  DFF_X1 u2_L9_reg_8 (.CK( clk ) , .Q( u2_L9_8 ) , .D( u2_R8_8 ) );
  DFF_X1 u2_L9_reg_9 (.CK( clk ) , .Q( u2_L9_9 ) , .D( u2_R8_9 ) );
  DFF_X1 u2_R0_reg_1 (.CK( clk ) , .D( u2_N0 ) , .Q( u2_R0_1 ) );
  DFF_X1 u2_R0_reg_10 (.CK( clk ) , .D( u2_N9 ) , .Q( u2_R0_10 ) );
  DFF_X1 u2_R0_reg_11 (.CK( clk ) , .D( u2_N10 ) , .Q( u2_R0_11 ) );
  DFF_X1 u2_R0_reg_12 (.CK( clk ) , .D( u2_N11 ) , .Q( u2_R0_12 ) );
  DFF_X1 u2_R0_reg_13 (.CK( clk ) , .D( u2_N12 ) , .Q( u2_R0_13 ) );
  DFF_X1 u2_R0_reg_14 (.CK( clk ) , .D( u2_N13 ) , .Q( u2_R0_14 ) );
  DFF_X1 u2_R0_reg_15 (.CK( clk ) , .D( u2_N14 ) , .Q( u2_R0_15 ) );
  DFF_X1 u2_R0_reg_16 (.CK( clk ) , .D( u2_N15 ) , .Q( u2_R0_16 ) );
  DFF_X1 u2_R0_reg_17 (.CK( clk ) , .D( u2_N16 ) , .Q( u2_R0_17 ) );
  DFF_X1 u2_R0_reg_18 (.CK( clk ) , .D( u2_N17 ) , .Q( u2_R0_18 ) );
  DFF_X1 u2_R0_reg_19 (.CK( clk ) , .D( u2_N18 ) , .Q( u2_R0_19 ) );
  DFF_X1 u2_R0_reg_2 (.CK( clk ) , .D( u2_N1 ) , .Q( u2_R0_2 ) );
  DFF_X1 u2_R0_reg_20 (.CK( clk ) , .D( u2_N19 ) , .Q( u2_R0_20 ) );
  DFF_X1 u2_R0_reg_21 (.CK( clk ) , .D( u2_N20 ) , .Q( u2_R0_21 ) );
  DFF_X1 u2_R0_reg_22 (.CK( clk ) , .D( u2_N21 ) , .Q( u2_R0_22 ) );
  DFF_X1 u2_R0_reg_23 (.CK( clk ) , .D( u2_N22 ) , .Q( u2_R0_23 ) );
  DFF_X1 u2_R0_reg_24 (.CK( clk ) , .D( u2_N23 ) , .Q( u2_R0_24 ) );
  DFF_X1 u2_R0_reg_25 (.CK( clk ) , .D( u2_N24 ) , .Q( u2_R0_25 ) );
  DFF_X1 u2_R0_reg_26 (.CK( clk ) , .D( u2_N25 ) , .Q( u2_R0_26 ) );
  DFF_X1 u2_R0_reg_27 (.CK( clk ) , .D( u2_N26 ) , .Q( u2_R0_27 ) );
  DFF_X1 u2_R0_reg_28 (.CK( clk ) , .D( u2_N27 ) , .Q( u2_R0_28 ) );
  DFF_X1 u2_R0_reg_29 (.CK( clk ) , .D( u2_N28 ) , .Q( u2_R0_29 ) );
  DFF_X1 u2_R0_reg_3 (.CK( clk ) , .D( u2_N2 ) , .Q( u2_R0_3 ) );
  DFF_X1 u2_R0_reg_30 (.CK( clk ) , .D( u2_N29 ) , .Q( u2_R0_30 ) );
  DFF_X1 u2_R0_reg_31 (.CK( clk ) , .D( u2_N30 ) , .Q( u2_R0_31 ) );
  DFF_X1 u2_R0_reg_32 (.CK( clk ) , .D( u2_N31 ) , .Q( u2_R0_32 ) );
  DFF_X1 u2_R0_reg_4 (.CK( clk ) , .D( u2_N3 ) , .Q( u2_R0_4 ) );
  DFF_X1 u2_R0_reg_5 (.CK( clk ) , .D( u2_N4 ) , .Q( u2_R0_5 ) );
  DFF_X1 u2_R0_reg_6 (.CK( clk ) , .D( u2_N5 ) , .Q( u2_R0_6 ) );
  DFF_X1 u2_R0_reg_7 (.CK( clk ) , .D( u2_N6 ) , .Q( u2_R0_7 ) );
  DFF_X1 u2_R0_reg_8 (.CK( clk ) , .D( u2_N7 ) , .Q( u2_R0_8 ) );
  DFF_X1 u2_R0_reg_9 (.CK( clk ) , .D( u2_N8 ) , .Q( u2_R0_9 ) );
  DFF_X1 u2_R10_reg_1 (.CK( clk ) , .D( u2_N320 ) , .Q( u2_R10_1 ) );
  DFF_X1 u2_R10_reg_10 (.CK( clk ) , .D( u2_N329 ) , .Q( u2_R10_10 ) );
  DFF_X1 u2_R10_reg_11 (.CK( clk ) , .D( u2_N330 ) , .Q( u2_R10_11 ) );
  DFF_X1 u2_R10_reg_12 (.CK( clk ) , .D( u2_N331 ) , .Q( u2_R10_12 ) );
  DFF_X1 u2_R10_reg_13 (.CK( clk ) , .D( u2_N332 ) , .Q( u2_R10_13 ) );
  DFF_X1 u2_R10_reg_14 (.CK( clk ) , .D( u2_N333 ) , .Q( u2_R10_14 ) );
  DFF_X1 u2_R10_reg_15 (.CK( clk ) , .D( u2_N334 ) , .Q( u2_R10_15 ) );
  DFF_X1 u2_R10_reg_16 (.CK( clk ) , .D( u2_N335 ) , .Q( u2_R10_16 ) );
  DFF_X1 u2_R10_reg_17 (.CK( clk ) , .D( u2_N336 ) , .Q( u2_R10_17 ) );
  DFF_X1 u2_R10_reg_18 (.CK( clk ) , .D( u2_N337 ) , .Q( u2_R10_18 ) );
  DFF_X1 u2_R10_reg_19 (.CK( clk ) , .D( u2_N338 ) , .Q( u2_R10_19 ) );
  DFF_X1 u2_R10_reg_2 (.CK( clk ) , .D( u2_N321 ) , .Q( u2_R10_2 ) );
  DFF_X1 u2_R10_reg_20 (.CK( clk ) , .D( u2_N339 ) , .Q( u2_R10_20 ) );
  DFF_X1 u2_R10_reg_21 (.CK( clk ) , .D( u2_N340 ) , .Q( u2_R10_21 ) );
  DFF_X1 u2_R10_reg_22 (.CK( clk ) , .D( u2_N341 ) , .Q( u2_R10_22 ) );
  DFF_X1 u2_R10_reg_23 (.CK( clk ) , .D( u2_N342 ) , .Q( u2_R10_23 ) );
  DFF_X1 u2_R10_reg_24 (.CK( clk ) , .D( u2_N343 ) , .Q( u2_R10_24 ) );
  DFF_X1 u2_R10_reg_25 (.CK( clk ) , .D( u2_N344 ) , .Q( u2_R10_25 ) );
  DFF_X1 u2_R10_reg_26 (.CK( clk ) , .D( u2_N345 ) , .Q( u2_R10_26 ) );
  DFF_X1 u2_R10_reg_27 (.CK( clk ) , .D( u2_N346 ) , .Q( u2_R10_27 ) );
  DFF_X1 u2_R10_reg_28 (.CK( clk ) , .D( u2_N347 ) , .Q( u2_R10_28 ) );
  DFF_X1 u2_R10_reg_29 (.CK( clk ) , .D( u2_N348 ) , .Q( u2_R10_29 ) );
  DFF_X1 u2_R10_reg_3 (.CK( clk ) , .D( u2_N322 ) , .Q( u2_R10_3 ) );
  DFF_X1 u2_R10_reg_30 (.CK( clk ) , .D( u2_N349 ) , .Q( u2_R10_30 ) );
  DFF_X1 u2_R10_reg_31 (.CK( clk ) , .D( u2_N350 ) , .Q( u2_R10_31 ) );
  DFF_X1 u2_R10_reg_32 (.CK( clk ) , .D( u2_N351 ) , .Q( u2_R10_32 ) );
  DFF_X1 u2_R10_reg_4 (.CK( clk ) , .D( u2_N323 ) , .Q( u2_R10_4 ) );
  DFF_X1 u2_R10_reg_5 (.CK( clk ) , .D( u2_N324 ) , .Q( u2_R10_5 ) );
  DFF_X1 u2_R10_reg_6 (.CK( clk ) , .D( u2_N325 ) , .Q( u2_R10_6 ) );
  DFF_X1 u2_R10_reg_7 (.CK( clk ) , .D( u2_N326 ) , .Q( u2_R10_7 ) );
  DFF_X1 u2_R10_reg_8 (.CK( clk ) , .D( u2_N327 ) , .Q( u2_R10_8 ) );
  DFF_X1 u2_R10_reg_9 (.CK( clk ) , .D( u2_N328 ) , .Q( u2_R10_9 ) );
  DFF_X1 u2_R11_reg_1 (.CK( clk ) , .D( u2_N352 ) , .Q( u2_R11_1 ) );
  DFF_X1 u2_R11_reg_10 (.CK( clk ) , .D( u2_N361 ) , .Q( u2_R11_10 ) );
  DFF_X1 u2_R11_reg_11 (.CK( clk ) , .D( u2_N362 ) , .Q( u2_R11_11 ) );
  DFF_X1 u2_R11_reg_12 (.CK( clk ) , .D( u2_N363 ) , .Q( u2_R11_12 ) );
  DFF_X1 u2_R11_reg_13 (.CK( clk ) , .D( u2_N364 ) , .Q( u2_R11_13 ) );
  DFF_X1 u2_R11_reg_14 (.CK( clk ) , .D( u2_N365 ) , .Q( u2_R11_14 ) );
  DFF_X1 u2_R11_reg_15 (.CK( clk ) , .D( u2_N366 ) , .Q( u2_R11_15 ) );
  DFF_X1 u2_R11_reg_16 (.CK( clk ) , .D( u2_N367 ) , .Q( u2_R11_16 ) );
  DFF_X1 u2_R11_reg_17 (.CK( clk ) , .D( u2_N368 ) , .Q( u2_R11_17 ) );
  DFF_X1 u2_R11_reg_18 (.CK( clk ) , .D( u2_N369 ) , .Q( u2_R11_18 ) );
  DFF_X1 u2_R11_reg_19 (.CK( clk ) , .D( u2_N370 ) , .Q( u2_R11_19 ) );
  DFF_X1 u2_R11_reg_2 (.CK( clk ) , .D( u2_N353 ) , .Q( u2_R11_2 ) );
  DFF_X1 u2_R11_reg_20 (.CK( clk ) , .D( u2_N371 ) , .Q( u2_R11_20 ) );
  DFF_X1 u2_R11_reg_21 (.CK( clk ) , .D( u2_N372 ) , .Q( u2_R11_21 ) );
  DFF_X1 u2_R11_reg_22 (.CK( clk ) , .D( u2_N373 ) , .Q( u2_R11_22 ) );
  DFF_X1 u2_R11_reg_23 (.CK( clk ) , .D( u2_N374 ) , .Q( u2_R11_23 ) );
  DFF_X1 u2_R11_reg_24 (.CK( clk ) , .D( u2_N375 ) , .Q( u2_R11_24 ) );
  DFF_X1 u2_R11_reg_25 (.CK( clk ) , .D( u2_N376 ) , .Q( u2_R11_25 ) );
  DFF_X1 u2_R11_reg_26 (.CK( clk ) , .D( u2_N377 ) , .Q( u2_R11_26 ) );
  DFF_X1 u2_R11_reg_27 (.CK( clk ) , .D( u2_N378 ) , .Q( u2_R11_27 ) );
  DFF_X1 u2_R11_reg_28 (.CK( clk ) , .D( u2_N379 ) , .Q( u2_R11_28 ) );
  DFF_X1 u2_R11_reg_29 (.CK( clk ) , .D( u2_N380 ) , .Q( u2_R11_29 ) );
  DFF_X1 u2_R11_reg_3 (.CK( clk ) , .D( u2_N354 ) , .Q( u2_R11_3 ) );
  DFF_X1 u2_R11_reg_30 (.CK( clk ) , .D( u2_N381 ) , .Q( u2_R11_30 ) );
  DFF_X1 u2_R11_reg_31 (.CK( clk ) , .D( u2_N382 ) , .Q( u2_R11_31 ) );
  DFF_X1 u2_R11_reg_32 (.CK( clk ) , .D( u2_N383 ) , .Q( u2_R11_32 ) );
  DFF_X1 u2_R11_reg_4 (.CK( clk ) , .D( u2_N355 ) , .Q( u2_R11_4 ) );
  DFF_X1 u2_R11_reg_5 (.CK( clk ) , .D( u2_N356 ) , .Q( u2_R11_5 ) );
  DFF_X1 u2_R11_reg_6 (.CK( clk ) , .D( u2_N357 ) , .Q( u2_R11_6 ) );
  DFF_X1 u2_R11_reg_7 (.CK( clk ) , .D( u2_N358 ) , .Q( u2_R11_7 ) );
  DFF_X1 u2_R11_reg_8 (.CK( clk ) , .D( u2_N359 ) , .Q( u2_R11_8 ) );
  DFF_X1 u2_R11_reg_9 (.CK( clk ) , .D( u2_N360 ) , .Q( u2_R11_9 ) );
  DFF_X1 u2_R12_reg_1 (.CK( clk ) , .D( u2_N384 ) , .Q( u2_R12_1 ) );
  DFF_X1 u2_R12_reg_10 (.CK( clk ) , .D( u2_N393 ) , .Q( u2_R12_10 ) );
  DFF_X1 u2_R12_reg_11 (.CK( clk ) , .D( u2_N394 ) , .Q( u2_R12_11 ) );
  DFF_X1 u2_R12_reg_12 (.CK( clk ) , .D( u2_N395 ) , .Q( u2_R12_12 ) );
  DFF_X1 u2_R12_reg_13 (.CK( clk ) , .D( u2_N396 ) , .Q( u2_R12_13 ) );
  DFF_X1 u2_R12_reg_14 (.CK( clk ) , .D( u2_N397 ) , .Q( u2_R12_14 ) );
  DFF_X1 u2_R12_reg_15 (.CK( clk ) , .D( u2_N398 ) , .Q( u2_R12_15 ) );
  DFF_X1 u2_R12_reg_16 (.CK( clk ) , .D( u2_N399 ) , .Q( u2_R12_16 ) );
  DFF_X1 u2_R12_reg_17 (.CK( clk ) , .D( u2_N400 ) , .Q( u2_R12_17 ) );
  DFF_X1 u2_R12_reg_18 (.CK( clk ) , .D( u2_N401 ) , .Q( u2_R12_18 ) );
  DFF_X1 u2_R12_reg_19 (.CK( clk ) , .D( u2_N402 ) , .Q( u2_R12_19 ) );
  DFF_X1 u2_R12_reg_2 (.CK( clk ) , .D( u2_N385 ) , .Q( u2_R12_2 ) );
  DFF_X1 u2_R12_reg_20 (.CK( clk ) , .D( u2_N403 ) , .Q( u2_R12_20 ) );
  DFF_X1 u2_R12_reg_21 (.CK( clk ) , .D( u2_N404 ) , .Q( u2_R12_21 ) );
  DFF_X1 u2_R12_reg_22 (.CK( clk ) , .D( u2_N405 ) , .Q( u2_R12_22 ) );
  DFF_X1 u2_R12_reg_23 (.CK( clk ) , .D( u2_N406 ) , .Q( u2_R12_23 ) );
  DFF_X1 u2_R12_reg_24 (.CK( clk ) , .D( u2_N407 ) , .Q( u2_R12_24 ) );
  DFF_X1 u2_R12_reg_25 (.CK( clk ) , .D( u2_N408 ) , .Q( u2_R12_25 ) );
  DFF_X1 u2_R12_reg_26 (.CK( clk ) , .D( u2_N409 ) , .Q( u2_R12_26 ) );
  DFF_X1 u2_R12_reg_27 (.CK( clk ) , .D( u2_N410 ) , .Q( u2_R12_27 ) );
  DFF_X1 u2_R12_reg_28 (.CK( clk ) , .D( u2_N411 ) , .Q( u2_R12_28 ) );
  DFF_X1 u2_R12_reg_29 (.CK( clk ) , .D( u2_N412 ) , .Q( u2_R12_29 ) );
  DFF_X1 u2_R12_reg_3 (.CK( clk ) , .D( u2_N386 ) , .Q( u2_R12_3 ) );
  DFF_X1 u2_R12_reg_30 (.CK( clk ) , .D( u2_N413 ) , .Q( u2_R12_30 ) );
  DFF_X1 u2_R12_reg_31 (.CK( clk ) , .D( u2_N414 ) , .Q( u2_R12_31 ) );
  DFF_X1 u2_R12_reg_32 (.CK( clk ) , .D( u2_N415 ) , .Q( u2_R12_32 ) );
  DFF_X1 u2_R12_reg_4 (.CK( clk ) , .D( u2_N387 ) , .Q( u2_R12_4 ) );
  DFF_X1 u2_R12_reg_5 (.CK( clk ) , .D( u2_N388 ) , .Q( u2_R12_5 ) );
  DFF_X1 u2_R12_reg_6 (.CK( clk ) , .D( u2_N389 ) , .Q( u2_R12_6 ) );
  DFF_X1 u2_R12_reg_7 (.CK( clk ) , .D( u2_N390 ) , .Q( u2_R12_7 ) );
  DFF_X1 u2_R12_reg_8 (.CK( clk ) , .D( u2_N391 ) , .Q( u2_R12_8 ) );
  DFF_X1 u2_R12_reg_9 (.CK( clk ) , .D( u2_N392 ) , .Q( u2_R12_9 ) );
  DFF_X1 u2_R13_reg_1 (.CK( clk ) , .D( u2_N416 ) , .Q( u2_R13_1 ) );
  DFF_X1 u2_R13_reg_10 (.CK( clk ) , .D( u2_N425 ) , .Q( u2_R13_10 ) );
  DFF_X1 u2_R13_reg_11 (.CK( clk ) , .D( u2_N426 ) , .Q( u2_R13_11 ) );
  DFF_X1 u2_R13_reg_12 (.CK( clk ) , .D( u2_N427 ) , .Q( u2_R13_12 ) );
  DFF_X1 u2_R13_reg_13 (.CK( clk ) , .D( u2_N428 ) , .Q( u2_R13_13 ) );
  DFF_X1 u2_R13_reg_14 (.CK( clk ) , .D( u2_N429 ) , .Q( u2_R13_14 ) );
  DFF_X1 u2_R13_reg_15 (.CK( clk ) , .D( u2_N430 ) , .Q( u2_R13_15 ) );
  DFF_X1 u2_R13_reg_16 (.CK( clk ) , .D( u2_N431 ) , .Q( u2_R13_16 ) );
  DFF_X1 u2_R13_reg_17 (.CK( clk ) , .D( u2_N432 ) , .Q( u2_R13_17 ) );
  DFF_X1 u2_R13_reg_18 (.CK( clk ) , .D( u2_N433 ) , .Q( u2_R13_18 ) );
  DFF_X1 u2_R13_reg_19 (.CK( clk ) , .D( u2_N434 ) , .Q( u2_R13_19 ) );
  DFF_X1 u2_R13_reg_2 (.CK( clk ) , .D( u2_N417 ) , .Q( u2_R13_2 ) );
  DFF_X1 u2_R13_reg_20 (.CK( clk ) , .D( u2_N435 ) , .Q( u2_R13_20 ) );
  DFF_X1 u2_R13_reg_21 (.CK( clk ) , .D( u2_N436 ) , .Q( u2_R13_21 ) );
  DFF_X1 u2_R13_reg_22 (.CK( clk ) , .D( u2_N437 ) , .Q( u2_R13_22 ) );
  DFF_X1 u2_R13_reg_23 (.CK( clk ) , .D( u2_N438 ) , .Q( u2_R13_23 ) );
  DFF_X1 u2_R13_reg_24 (.CK( clk ) , .D( u2_N439 ) , .Q( u2_R13_24 ) );
  DFF_X1 u2_R13_reg_25 (.CK( clk ) , .D( u2_N440 ) , .Q( u2_R13_25 ) );
  DFF_X1 u2_R13_reg_26 (.CK( clk ) , .D( u2_N441 ) , .Q( u2_R13_26 ) );
  DFF_X1 u2_R13_reg_27 (.CK( clk ) , .D( u2_N442 ) , .Q( u2_R13_27 ) );
  DFF_X1 u2_R13_reg_28 (.CK( clk ) , .D( u2_N443 ) , .Q( u2_R13_28 ) );
  DFF_X1 u2_R13_reg_29 (.CK( clk ) , .D( u2_N444 ) , .Q( u2_R13_29 ) );
  DFF_X1 u2_R13_reg_3 (.CK( clk ) , .D( u2_N418 ) , .Q( u2_R13_3 ) );
  DFF_X1 u2_R13_reg_30 (.CK( clk ) , .D( u2_N445 ) , .Q( u2_R13_30 ) );
  DFF_X1 u2_R13_reg_31 (.CK( clk ) , .D( u2_N446 ) , .Q( u2_R13_31 ) );
  DFF_X1 u2_R13_reg_32 (.CK( clk ) , .D( u2_N447 ) , .Q( u2_R13_32 ) );
  DFF_X1 u2_R13_reg_4 (.CK( clk ) , .D( u2_N419 ) , .Q( u2_R13_4 ) );
  DFF_X1 u2_R13_reg_5 (.CK( clk ) , .D( u2_N420 ) , .Q( u2_R13_5 ) );
  DFF_X1 u2_R13_reg_6 (.CK( clk ) , .D( u2_N421 ) , .Q( u2_R13_6 ) );
  DFF_X1 u2_R13_reg_7 (.CK( clk ) , .D( u2_N422 ) , .Q( u2_R13_7 ) );
  DFF_X1 u2_R13_reg_8 (.CK( clk ) , .D( u2_N423 ) , .Q( u2_R13_8 ) );
  DFF_X1 u2_R13_reg_9 (.CK( clk ) , .D( u2_N424 ) , .Q( u2_R13_9 ) );
  DFF_X1 u2_R14_reg_1 (.CK( clk ) , .Q( u2_FP_33 ) , .D( u2_N448 ) );
  DFF_X1 u2_R14_reg_10 (.CK( clk ) , .Q( u2_FP_42 ) , .D( u2_N457 ) );
  DFF_X1 u2_R14_reg_11 (.CK( clk ) , .Q( u2_FP_43 ) , .D( u2_N458 ) );
  DFF_X1 u2_R14_reg_12 (.CK( clk ) , .Q( u2_FP_44 ) , .D( u2_N459 ) );
  DFF_X1 u2_R14_reg_13 (.CK( clk ) , .Q( u2_FP_45 ) , .D( u2_N460 ) );
  DFF_X1 u2_R14_reg_14 (.CK( clk ) , .Q( u2_FP_46 ) , .D( u2_N461 ) );
  DFF_X1 u2_R14_reg_15 (.CK( clk ) , .Q( u2_FP_47 ) , .D( u2_N462 ) );
  DFF_X1 u2_R14_reg_16 (.CK( clk ) , .Q( u2_FP_48 ) , .D( u2_N463 ) );
  DFF_X1 u2_R14_reg_17 (.CK( clk ) , .Q( u2_FP_49 ) , .D( u2_N464 ) );
  DFF_X1 u2_R14_reg_18 (.CK( clk ) , .Q( u2_FP_50 ) , .D( u2_N465 ) );
  DFF_X1 u2_R14_reg_19 (.CK( clk ) , .Q( u2_FP_51 ) , .D( u2_N466 ) );
  DFF_X1 u2_R14_reg_2 (.CK( clk ) , .Q( u2_FP_34 ) , .D( u2_N449 ) );
  DFF_X1 u2_R14_reg_20 (.CK( clk ) , .Q( u2_FP_52 ) , .D( u2_N467 ) );
  DFF_X1 u2_R14_reg_21 (.CK( clk ) , .Q( u2_FP_53 ) , .D( u2_N468 ) );
  DFF_X1 u2_R14_reg_22 (.CK( clk ) , .Q( u2_FP_54 ) , .D( u2_N469 ) );
  DFF_X1 u2_R14_reg_23 (.CK( clk ) , .Q( u2_FP_55 ) , .D( u2_N470 ) );
  DFF_X1 u2_R14_reg_24 (.CK( clk ) , .Q( u2_FP_56 ) , .D( u2_N471 ) );
  DFF_X1 u2_R14_reg_25 (.CK( clk ) , .Q( u2_FP_57 ) , .D( u2_N472 ) );
  DFF_X1 u2_R14_reg_26 (.CK( clk ) , .Q( u2_FP_58 ) , .D( u2_N473 ) );
  DFF_X1 u2_R14_reg_27 (.CK( clk ) , .Q( u2_FP_59 ) , .D( u2_N474 ) );
  DFF_X1 u2_R14_reg_28 (.CK( clk ) , .Q( u2_FP_60 ) , .D( u2_N475 ) );
  DFF_X1 u2_R14_reg_29 (.CK( clk ) , .Q( u2_FP_61 ) , .D( u2_N476 ) );
  DFF_X1 u2_R14_reg_3 (.CK( clk ) , .Q( u2_FP_35 ) , .D( u2_N450 ) );
  DFF_X1 u2_R14_reg_30 (.CK( clk ) , .Q( u2_FP_62 ) , .D( u2_N477 ) );
  DFF_X1 u2_R14_reg_31 (.CK( clk ) , .Q( u2_FP_63 ) , .D( u2_N478 ) );
  DFF_X1 u2_R14_reg_32 (.CK( clk ) , .Q( u2_FP_64 ) , .D( u2_N479 ) );
  DFF_X1 u2_R14_reg_4 (.CK( clk ) , .Q( u2_FP_36 ) , .D( u2_N451 ) );
  DFF_X1 u2_R14_reg_5 (.CK( clk ) , .Q( u2_FP_37 ) , .D( u2_N452 ) );
  DFF_X1 u2_R14_reg_6 (.CK( clk ) , .Q( u2_FP_38 ) , .D( u2_N453 ) );
  DFF_X1 u2_R14_reg_7 (.CK( clk ) , .Q( u2_FP_39 ) , .D( u2_N454 ) );
  DFF_X1 u2_R14_reg_8 (.CK( clk ) , .Q( u2_FP_40 ) , .D( u2_N455 ) );
  DFF_X1 u2_R14_reg_9 (.CK( clk ) , .Q( u2_FP_41 ) , .D( u2_N456 ) );
  DFF_X1 u2_R1_reg_1 (.CK( clk ) , .D( u2_N32 ) , .Q( u2_R1_1 ) );
  DFF_X1 u2_R1_reg_10 (.CK( clk ) , .D( u2_N41 ) , .Q( u2_R1_10 ) );
  DFF_X1 u2_R1_reg_11 (.CK( clk ) , .D( u2_N42 ) , .Q( u2_R1_11 ) );
  DFF_X1 u2_R1_reg_12 (.CK( clk ) , .D( u2_N43 ) , .Q( u2_R1_12 ) );
  DFF_X1 u2_R1_reg_13 (.CK( clk ) , .D( u2_N44 ) , .Q( u2_R1_13 ) );
  DFF_X1 u2_R1_reg_14 (.CK( clk ) , .D( u2_N45 ) , .Q( u2_R1_14 ) );
  DFF_X1 u2_R1_reg_15 (.CK( clk ) , .D( u2_N46 ) , .Q( u2_R1_15 ) );
  DFF_X1 u2_R1_reg_16 (.CK( clk ) , .D( u2_N47 ) , .Q( u2_R1_16 ) );
  DFF_X1 u2_R1_reg_17 (.CK( clk ) , .D( u2_N48 ) , .Q( u2_R1_17 ) );
  DFF_X1 u2_R1_reg_18 (.CK( clk ) , .D( u2_N49 ) , .Q( u2_R1_18 ) );
  DFF_X1 u2_R1_reg_19 (.CK( clk ) , .D( u2_N50 ) , .Q( u2_R1_19 ) );
  DFF_X1 u2_R1_reg_2 (.CK( clk ) , .D( u2_N33 ) , .Q( u2_R1_2 ) );
  DFF_X1 u2_R1_reg_20 (.CK( clk ) , .D( u2_N51 ) , .Q( u2_R1_20 ) );
  DFF_X1 u2_R1_reg_21 (.CK( clk ) , .D( u2_N52 ) , .Q( u2_R1_21 ) );
  DFF_X1 u2_R1_reg_22 (.CK( clk ) , .D( u2_N53 ) , .Q( u2_R1_22 ) );
  DFF_X1 u2_R1_reg_23 (.CK( clk ) , .D( u2_N54 ) , .Q( u2_R1_23 ) );
  DFF_X1 u2_R1_reg_24 (.CK( clk ) , .D( u2_N55 ) , .Q( u2_R1_24 ) );
  DFF_X1 u2_R1_reg_25 (.CK( clk ) , .D( u2_N56 ) , .Q( u2_R1_25 ) );
  DFF_X1 u2_R1_reg_26 (.CK( clk ) , .D( u2_N57 ) , .Q( u2_R1_26 ) );
  DFF_X1 u2_R1_reg_27 (.CK( clk ) , .D( u2_N58 ) , .Q( u2_R1_27 ) );
  DFF_X1 u2_R1_reg_28 (.CK( clk ) , .D( u2_N59 ) , .Q( u2_R1_28 ) );
  DFF_X1 u2_R1_reg_29 (.CK( clk ) , .D( u2_N60 ) , .Q( u2_R1_29 ) );
  DFF_X1 u2_R1_reg_3 (.CK( clk ) , .D( u2_N34 ) , .Q( u2_R1_3 ) );
  DFF_X1 u2_R1_reg_30 (.CK( clk ) , .D( u2_N61 ) , .Q( u2_R1_30 ) );
  DFF_X1 u2_R1_reg_31 (.CK( clk ) , .D( u2_N62 ) , .Q( u2_R1_31 ) );
  DFF_X1 u2_R1_reg_32 (.CK( clk ) , .D( u2_N63 ) , .Q( u2_R1_32 ) );
  DFF_X1 u2_R1_reg_4 (.CK( clk ) , .D( u2_N35 ) , .Q( u2_R1_4 ) );
  DFF_X1 u2_R1_reg_5 (.CK( clk ) , .D( u2_N36 ) , .Q( u2_R1_5 ) );
  DFF_X1 u2_R1_reg_6 (.CK( clk ) , .D( u2_N37 ) , .Q( u2_R1_6 ) );
  DFF_X1 u2_R1_reg_7 (.CK( clk ) , .D( u2_N38 ) , .Q( u2_R1_7 ) );
  DFF_X1 u2_R1_reg_8 (.CK( clk ) , .D( u2_N39 ) , .Q( u2_R1_8 ) );
  DFF_X1 u2_R1_reg_9 (.CK( clk ) , .D( u2_N40 ) , .Q( u2_R1_9 ) );
  DFF_X1 u2_R2_reg_1 (.CK( clk ) , .D( u2_N64 ) , .Q( u2_R2_1 ) );
  DFF_X1 u2_R2_reg_10 (.CK( clk ) , .D( u2_N73 ) , .Q( u2_R2_10 ) );
  DFF_X1 u2_R2_reg_11 (.CK( clk ) , .D( u2_N74 ) , .Q( u2_R2_11 ) );
  DFF_X1 u2_R2_reg_12 (.CK( clk ) , .D( u2_N75 ) , .Q( u2_R2_12 ) );
  DFF_X1 u2_R2_reg_13 (.CK( clk ) , .D( u2_N76 ) , .Q( u2_R2_13 ) );
  DFF_X1 u2_R2_reg_14 (.CK( clk ) , .D( u2_N77 ) , .Q( u2_R2_14 ) );
  DFF_X1 u2_R2_reg_15 (.CK( clk ) , .D( u2_N78 ) , .Q( u2_R2_15 ) );
  DFF_X1 u2_R2_reg_16 (.CK( clk ) , .D( u2_N79 ) , .Q( u2_R2_16 ) );
  DFF_X1 u2_R2_reg_17 (.CK( clk ) , .D( u2_N80 ) , .Q( u2_R2_17 ) );
  DFF_X1 u2_R2_reg_18 (.CK( clk ) , .D( u2_N81 ) , .Q( u2_R2_18 ) );
  DFF_X1 u2_R2_reg_19 (.CK( clk ) , .D( u2_N82 ) , .Q( u2_R2_19 ) );
  DFF_X1 u2_R2_reg_2 (.CK( clk ) , .D( u2_N65 ) , .Q( u2_R2_2 ) );
  DFF_X1 u2_R2_reg_20 (.CK( clk ) , .D( u2_N83 ) , .Q( u2_R2_20 ) );
  DFF_X1 u2_R2_reg_21 (.CK( clk ) , .D( u2_N84 ) , .Q( u2_R2_21 ) );
  DFF_X1 u2_R2_reg_22 (.CK( clk ) , .D( u2_N85 ) , .Q( u2_R2_22 ) );
  DFF_X1 u2_R2_reg_23 (.CK( clk ) , .D( u2_N86 ) , .Q( u2_R2_23 ) );
  DFF_X1 u2_R2_reg_24 (.CK( clk ) , .D( u2_N87 ) , .Q( u2_R2_24 ) );
  DFF_X1 u2_R2_reg_25 (.CK( clk ) , .D( u2_N88 ) , .Q( u2_R2_25 ) );
  DFF_X1 u2_R2_reg_26 (.CK( clk ) , .D( u2_N89 ) , .Q( u2_R2_26 ) );
  DFF_X1 u2_R2_reg_27 (.CK( clk ) , .D( u2_N90 ) , .Q( u2_R2_27 ) );
  DFF_X1 u2_R2_reg_28 (.CK( clk ) , .D( u2_N91 ) , .Q( u2_R2_28 ) );
  DFF_X1 u2_R2_reg_29 (.CK( clk ) , .D( u2_N92 ) , .Q( u2_R2_29 ) );
  DFF_X1 u2_R2_reg_3 (.CK( clk ) , .D( u2_N66 ) , .Q( u2_R2_3 ) );
  DFF_X1 u2_R2_reg_30 (.CK( clk ) , .D( u2_N93 ) , .Q( u2_R2_30 ) );
  DFF_X1 u2_R2_reg_31 (.CK( clk ) , .D( u2_N94 ) , .Q( u2_R2_31 ) );
  DFF_X1 u2_R2_reg_32 (.CK( clk ) , .D( u2_N95 ) , .Q( u2_R2_32 ) );
  DFF_X1 u2_R2_reg_4 (.CK( clk ) , .D( u2_N67 ) , .Q( u2_R2_4 ) );
  DFF_X1 u2_R2_reg_5 (.CK( clk ) , .D( u2_N68 ) , .Q( u2_R2_5 ) );
  DFF_X1 u2_R2_reg_6 (.CK( clk ) , .D( u2_N69 ) , .Q( u2_R2_6 ) );
  DFF_X1 u2_R2_reg_7 (.CK( clk ) , .D( u2_N70 ) , .Q( u2_R2_7 ) );
  DFF_X1 u2_R2_reg_8 (.CK( clk ) , .D( u2_N71 ) , .Q( u2_R2_8 ) );
  DFF_X1 u2_R2_reg_9 (.CK( clk ) , .D( u2_N72 ) , .Q( u2_R2_9 ) );
  DFF_X1 u2_R3_reg_1 (.CK( clk ) , .D( u2_N96 ) , .Q( u2_R3_1 ) );
  DFF_X1 u2_R3_reg_10 (.CK( clk ) , .D( u2_N105 ) , .Q( u2_R3_10 ) );
  DFF_X1 u2_R3_reg_11 (.CK( clk ) , .D( u2_N106 ) , .Q( u2_R3_11 ) );
  DFF_X1 u2_R3_reg_12 (.CK( clk ) , .D( u2_N107 ) , .Q( u2_R3_12 ) );
  DFF_X1 u2_R3_reg_13 (.CK( clk ) , .D( u2_N108 ) , .Q( u2_R3_13 ) );
  DFF_X1 u2_R3_reg_14 (.CK( clk ) , .D( u2_N109 ) , .Q( u2_R3_14 ) );
  DFF_X1 u2_R3_reg_15 (.CK( clk ) , .D( u2_N110 ) , .Q( u2_R3_15 ) );
  DFF_X1 u2_R3_reg_16 (.CK( clk ) , .D( u2_N111 ) , .Q( u2_R3_16 ) );
  DFF_X1 u2_R3_reg_17 (.CK( clk ) , .D( u2_N112 ) , .Q( u2_R3_17 ) );
  DFF_X1 u2_R3_reg_18 (.CK( clk ) , .D( u2_N113 ) , .Q( u2_R3_18 ) );
  DFF_X1 u2_R3_reg_19 (.CK( clk ) , .D( u2_N114 ) , .Q( u2_R3_19 ) );
  DFF_X1 u2_R3_reg_2 (.CK( clk ) , .D( u2_N97 ) , .Q( u2_R3_2 ) );
  DFF_X1 u2_R3_reg_20 (.CK( clk ) , .D( u2_N115 ) , .Q( u2_R3_20 ) );
  DFF_X1 u2_R3_reg_21 (.CK( clk ) , .D( u2_N116 ) , .Q( u2_R3_21 ) );
  DFF_X1 u2_R3_reg_22 (.CK( clk ) , .D( u2_N117 ) , .Q( u2_R3_22 ) );
  DFF_X1 u2_R3_reg_23 (.CK( clk ) , .D( u2_N118 ) , .Q( u2_R3_23 ) );
  DFF_X1 u2_R3_reg_24 (.CK( clk ) , .D( u2_N119 ) , .Q( u2_R3_24 ) );
  DFF_X1 u2_R3_reg_25 (.CK( clk ) , .D( u2_N120 ) , .Q( u2_R3_25 ) );
  DFF_X1 u2_R3_reg_26 (.CK( clk ) , .D( u2_N121 ) , .Q( u2_R3_26 ) );
  DFF_X1 u2_R3_reg_27 (.CK( clk ) , .D( u2_N122 ) , .Q( u2_R3_27 ) );
  DFF_X1 u2_R3_reg_28 (.CK( clk ) , .D( u2_N123 ) , .Q( u2_R3_28 ) );
  DFF_X1 u2_R3_reg_29 (.CK( clk ) , .D( u2_N124 ) , .Q( u2_R3_29 ) );
  DFF_X1 u2_R3_reg_3 (.CK( clk ) , .D( u2_N98 ) , .Q( u2_R3_3 ) );
  DFF_X1 u2_R3_reg_30 (.CK( clk ) , .D( u2_N125 ) , .Q( u2_R3_30 ) );
  DFF_X1 u2_R3_reg_31 (.CK( clk ) , .D( u2_N126 ) , .Q( u2_R3_31 ) );
  DFF_X1 u2_R3_reg_32 (.CK( clk ) , .D( u2_N127 ) , .Q( u2_R3_32 ) );
  DFF_X1 u2_R3_reg_4 (.CK( clk ) , .D( u2_N99 ) , .Q( u2_R3_4 ) );
  DFF_X1 u2_R3_reg_5 (.CK( clk ) , .D( u2_N100 ) , .Q( u2_R3_5 ) );
  DFF_X1 u2_R3_reg_6 (.CK( clk ) , .D( u2_N101 ) , .Q( u2_R3_6 ) );
  DFF_X1 u2_R3_reg_7 (.CK( clk ) , .D( u2_N102 ) , .Q( u2_R3_7 ) );
  DFF_X1 u2_R3_reg_8 (.CK( clk ) , .D( u2_N103 ) , .Q( u2_R3_8 ) );
  DFF_X1 u2_R3_reg_9 (.CK( clk ) , .D( u2_N104 ) , .Q( u2_R3_9 ) );
  DFF_X1 u2_R4_reg_1 (.CK( clk ) , .D( u2_N128 ) , .Q( u2_R4_1 ) );
  DFF_X1 u2_R4_reg_10 (.CK( clk ) , .D( u2_N137 ) , .Q( u2_R4_10 ) );
  DFF_X1 u2_R4_reg_11 (.CK( clk ) , .D( u2_N138 ) , .Q( u2_R4_11 ) );
  DFF_X1 u2_R4_reg_12 (.CK( clk ) , .D( u2_N139 ) , .Q( u2_R4_12 ) );
  DFF_X1 u2_R4_reg_13 (.CK( clk ) , .D( u2_N140 ) , .Q( u2_R4_13 ) );
  DFF_X1 u2_R4_reg_14 (.CK( clk ) , .D( u2_N141 ) , .Q( u2_R4_14 ) );
  DFF_X1 u2_R4_reg_15 (.CK( clk ) , .D( u2_N142 ) , .Q( u2_R4_15 ) );
  DFF_X1 u2_R4_reg_16 (.CK( clk ) , .D( u2_N143 ) , .Q( u2_R4_16 ) );
  DFF_X1 u2_R4_reg_17 (.CK( clk ) , .D( u2_N144 ) , .Q( u2_R4_17 ) );
  DFF_X1 u2_R4_reg_18 (.CK( clk ) , .D( u2_N145 ) , .Q( u2_R4_18 ) );
  DFF_X1 u2_R4_reg_19 (.CK( clk ) , .D( u2_N146 ) , .Q( u2_R4_19 ) );
  DFF_X1 u2_R4_reg_2 (.CK( clk ) , .D( u2_N129 ) , .Q( u2_R4_2 ) );
  DFF_X1 u2_R4_reg_20 (.CK( clk ) , .D( u2_N147 ) , .Q( u2_R4_20 ) );
  DFF_X1 u2_R4_reg_21 (.CK( clk ) , .D( u2_N148 ) , .Q( u2_R4_21 ) );
  DFF_X1 u2_R4_reg_22 (.CK( clk ) , .D( u2_N149 ) , .Q( u2_R4_22 ) );
  DFF_X1 u2_R4_reg_23 (.CK( clk ) , .D( u2_N150 ) , .Q( u2_R4_23 ) );
  DFF_X1 u2_R4_reg_24 (.CK( clk ) , .D( u2_N151 ) , .Q( u2_R4_24 ) );
  DFF_X1 u2_R4_reg_25 (.CK( clk ) , .D( u2_N152 ) , .Q( u2_R4_25 ) );
  DFF_X1 u2_R4_reg_26 (.CK( clk ) , .D( u2_N153 ) , .Q( u2_R4_26 ) );
  DFF_X1 u2_R4_reg_27 (.CK( clk ) , .D( u2_N154 ) , .Q( u2_R4_27 ) );
  DFF_X1 u2_R4_reg_28 (.CK( clk ) , .D( u2_N155 ) , .Q( u2_R4_28 ) );
  DFF_X1 u2_R4_reg_29 (.CK( clk ) , .D( u2_N156 ) , .Q( u2_R4_29 ) );
  DFF_X1 u2_R4_reg_3 (.CK( clk ) , .D( u2_N130 ) , .Q( u2_R4_3 ) );
  DFF_X1 u2_R4_reg_30 (.CK( clk ) , .D( u2_N157 ) , .Q( u2_R4_30 ) );
  DFF_X1 u2_R4_reg_31 (.CK( clk ) , .D( u2_N158 ) , .Q( u2_R4_31 ) );
  DFF_X1 u2_R4_reg_32 (.CK( clk ) , .D( u2_N159 ) , .Q( u2_R4_32 ) );
  DFF_X1 u2_R4_reg_4 (.CK( clk ) , .D( u2_N131 ) , .Q( u2_R4_4 ) );
  DFF_X1 u2_R4_reg_5 (.CK( clk ) , .D( u2_N132 ) , .Q( u2_R4_5 ) );
  DFF_X1 u2_R4_reg_6 (.CK( clk ) , .D( u2_N133 ) , .Q( u2_R4_6 ) );
  DFF_X1 u2_R4_reg_7 (.CK( clk ) , .D( u2_N134 ) , .Q( u2_R4_7 ) );
  DFF_X1 u2_R4_reg_8 (.CK( clk ) , .D( u2_N135 ) , .Q( u2_R4_8 ) );
  DFF_X1 u2_R4_reg_9 (.CK( clk ) , .D( u2_N136 ) , .Q( u2_R4_9 ) );
  DFF_X1 u2_R5_reg_1 (.CK( clk ) , .D( u2_N160 ) , .Q( u2_R5_1 ) );
  DFF_X1 u2_R5_reg_10 (.CK( clk ) , .D( u2_N169 ) , .Q( u2_R5_10 ) );
  DFF_X1 u2_R5_reg_11 (.CK( clk ) , .D( u2_N170 ) , .Q( u2_R5_11 ) );
  DFF_X1 u2_R5_reg_12 (.CK( clk ) , .D( u2_N171 ) , .Q( u2_R5_12 ) );
  DFF_X1 u2_R5_reg_13 (.CK( clk ) , .D( u2_N172 ) , .Q( u2_R5_13 ) );
  DFF_X1 u2_R5_reg_14 (.CK( clk ) , .D( u2_N173 ) , .Q( u2_R5_14 ) );
  DFF_X1 u2_R5_reg_15 (.CK( clk ) , .D( u2_N174 ) , .Q( u2_R5_15 ) );
  DFF_X1 u2_R5_reg_16 (.CK( clk ) , .D( u2_N175 ) , .Q( u2_R5_16 ) );
  DFF_X1 u2_R5_reg_17 (.CK( clk ) , .D( u2_N176 ) , .Q( u2_R5_17 ) );
  DFF_X1 u2_R5_reg_18 (.CK( clk ) , .D( u2_N177 ) , .Q( u2_R5_18 ) );
  DFF_X1 u2_R5_reg_19 (.CK( clk ) , .D( u2_N178 ) , .Q( u2_R5_19 ) );
  DFF_X1 u2_R5_reg_2 (.CK( clk ) , .D( u2_N161 ) , .Q( u2_R5_2 ) );
  DFF_X1 u2_R5_reg_20 (.CK( clk ) , .D( u2_N179 ) , .Q( u2_R5_20 ) );
  DFF_X1 u2_R5_reg_21 (.CK( clk ) , .D( u2_N180 ) , .Q( u2_R5_21 ) );
  DFF_X1 u2_R5_reg_22 (.CK( clk ) , .D( u2_N181 ) , .Q( u2_R5_22 ) );
  DFF_X1 u2_R5_reg_23 (.CK( clk ) , .D( u2_N182 ) , .Q( u2_R5_23 ) );
  DFF_X1 u2_R5_reg_24 (.CK( clk ) , .D( u2_N183 ) , .Q( u2_R5_24 ) );
  DFF_X1 u2_R5_reg_25 (.CK( clk ) , .D( u2_N184 ) , .Q( u2_R5_25 ) );
  DFF_X1 u2_R5_reg_26 (.CK( clk ) , .D( u2_N185 ) , .Q( u2_R5_26 ) );
  DFF_X1 u2_R5_reg_27 (.CK( clk ) , .D( u2_N186 ) , .Q( u2_R5_27 ) );
  DFF_X1 u2_R5_reg_28 (.CK( clk ) , .D( u2_N187 ) , .Q( u2_R5_28 ) );
  DFF_X1 u2_R5_reg_29 (.CK( clk ) , .D( u2_N188 ) , .Q( u2_R5_29 ) );
  DFF_X1 u2_R5_reg_3 (.CK( clk ) , .D( u2_N162 ) , .Q( u2_R5_3 ) );
  DFF_X1 u2_R5_reg_30 (.CK( clk ) , .D( u2_N189 ) , .Q( u2_R5_30 ) );
  DFF_X1 u2_R5_reg_31 (.CK( clk ) , .D( u2_N190 ) , .Q( u2_R5_31 ) );
  DFF_X1 u2_R5_reg_32 (.CK( clk ) , .D( u2_N191 ) , .Q( u2_R5_32 ) );
  DFF_X1 u2_R5_reg_4 (.CK( clk ) , .D( u2_N163 ) , .Q( u2_R5_4 ) );
  DFF_X1 u2_R5_reg_5 (.CK( clk ) , .D( u2_N164 ) , .Q( u2_R5_5 ) );
  DFF_X1 u2_R5_reg_6 (.CK( clk ) , .D( u2_N165 ) , .Q( u2_R5_6 ) );
  DFF_X1 u2_R5_reg_7 (.CK( clk ) , .D( u2_N166 ) , .Q( u2_R5_7 ) );
  DFF_X1 u2_R5_reg_8 (.CK( clk ) , .D( u2_N167 ) , .Q( u2_R5_8 ) );
  DFF_X1 u2_R5_reg_9 (.CK( clk ) , .D( u2_N168 ) , .Q( u2_R5_9 ) );
  DFF_X1 u2_R6_reg_1 (.CK( clk ) , .D( u2_N192 ) , .Q( u2_R6_1 ) );
  DFF_X1 u2_R6_reg_10 (.CK( clk ) , .D( u2_N201 ) , .Q( u2_R6_10 ) );
  DFF_X1 u2_R6_reg_11 (.CK( clk ) , .D( u2_N202 ) , .Q( u2_R6_11 ) );
  DFF_X1 u2_R6_reg_12 (.CK( clk ) , .D( u2_N203 ) , .Q( u2_R6_12 ) );
  DFF_X1 u2_R6_reg_13 (.CK( clk ) , .D( u2_N204 ) , .Q( u2_R6_13 ) );
  DFF_X1 u2_R6_reg_14 (.CK( clk ) , .D( u2_N205 ) , .Q( u2_R6_14 ) );
  DFF_X1 u2_R6_reg_15 (.CK( clk ) , .D( u2_N206 ) , .Q( u2_R6_15 ) );
  DFF_X1 u2_R6_reg_16 (.CK( clk ) , .D( u2_N207 ) , .Q( u2_R6_16 ) );
  DFF_X1 u2_R6_reg_17 (.CK( clk ) , .D( u2_N208 ) , .Q( u2_R6_17 ) );
  DFF_X1 u2_R6_reg_18 (.CK( clk ) , .D( u2_N209 ) , .Q( u2_R6_18 ) );
  DFF_X1 u2_R6_reg_19 (.CK( clk ) , .D( u2_N210 ) , .Q( u2_R6_19 ) );
  DFF_X1 u2_R6_reg_2 (.CK( clk ) , .D( u2_N193 ) , .Q( u2_R6_2 ) );
  DFF_X1 u2_R6_reg_20 (.CK( clk ) , .D( u2_N211 ) , .Q( u2_R6_20 ) );
  DFF_X1 u2_R6_reg_21 (.CK( clk ) , .D( u2_N212 ) , .Q( u2_R6_21 ) );
  DFF_X1 u2_R6_reg_22 (.CK( clk ) , .D( u2_N213 ) , .Q( u2_R6_22 ) );
  DFF_X1 u2_R6_reg_23 (.CK( clk ) , .D( u2_N214 ) , .Q( u2_R6_23 ) );
  DFF_X1 u2_R6_reg_24 (.CK( clk ) , .D( u2_N215 ) , .Q( u2_R6_24 ) );
  DFF_X1 u2_R6_reg_25 (.CK( clk ) , .D( u2_N216 ) , .Q( u2_R6_25 ) );
  DFF_X1 u2_R6_reg_26 (.CK( clk ) , .D( u2_N217 ) , .Q( u2_R6_26 ) );
  DFF_X1 u2_R6_reg_27 (.CK( clk ) , .D( u2_N218 ) , .Q( u2_R6_27 ) );
  DFF_X1 u2_R6_reg_28 (.CK( clk ) , .D( u2_N219 ) , .Q( u2_R6_28 ) );
  DFF_X1 u2_R6_reg_29 (.CK( clk ) , .D( u2_N220 ) , .Q( u2_R6_29 ) );
  DFF_X1 u2_R6_reg_3 (.CK( clk ) , .D( u2_N194 ) , .Q( u2_R6_3 ) );
  DFF_X1 u2_R6_reg_30 (.CK( clk ) , .D( u2_N221 ) , .Q( u2_R6_30 ) );
  DFF_X1 u2_R6_reg_31 (.CK( clk ) , .D( u2_N222 ) , .Q( u2_R6_31 ) );
  DFF_X1 u2_R6_reg_32 (.CK( clk ) , .D( u2_N223 ) , .Q( u2_R6_32 ) );
  DFF_X1 u2_R6_reg_4 (.CK( clk ) , .D( u2_N195 ) , .Q( u2_R6_4 ) );
  DFF_X1 u2_R6_reg_5 (.CK( clk ) , .D( u2_N196 ) , .Q( u2_R6_5 ) );
  DFF_X1 u2_R6_reg_6 (.CK( clk ) , .D( u2_N197 ) , .Q( u2_R6_6 ) );
  DFF_X1 u2_R6_reg_7 (.CK( clk ) , .D( u2_N198 ) , .Q( u2_R6_7 ) );
  DFF_X1 u2_R6_reg_8 (.CK( clk ) , .D( u2_N199 ) , .Q( u2_R6_8 ) );
  DFF_X1 u2_R6_reg_9 (.CK( clk ) , .D( u2_N200 ) , .Q( u2_R6_9 ) );
  DFF_X1 u2_R7_reg_1 (.CK( clk ) , .D( u2_N224 ) , .Q( u2_R7_1 ) );
  DFF_X1 u2_R7_reg_10 (.CK( clk ) , .D( u2_N233 ) , .Q( u2_R7_10 ) );
  DFF_X1 u2_R7_reg_11 (.CK( clk ) , .D( u2_N234 ) , .Q( u2_R7_11 ) );
  DFF_X1 u2_R7_reg_12 (.CK( clk ) , .D( u2_N235 ) , .Q( u2_R7_12 ) );
  DFF_X1 u2_R7_reg_13 (.CK( clk ) , .D( u2_N236 ) , .Q( u2_R7_13 ) );
  DFF_X1 u2_R7_reg_14 (.CK( clk ) , .D( u2_N237 ) , .Q( u2_R7_14 ) );
  DFF_X1 u2_R7_reg_15 (.CK( clk ) , .D( u2_N238 ) , .Q( u2_R7_15 ) );
  DFF_X1 u2_R7_reg_16 (.CK( clk ) , .D( u2_N239 ) , .Q( u2_R7_16 ) );
  DFF_X1 u2_R7_reg_17 (.CK( clk ) , .D( u2_N240 ) , .Q( u2_R7_17 ) );
  DFF_X1 u2_R7_reg_18 (.CK( clk ) , .D( u2_N241 ) , .Q( u2_R7_18 ) );
  DFF_X1 u2_R7_reg_19 (.CK( clk ) , .D( u2_N242 ) , .Q( u2_R7_19 ) );
  DFF_X1 u2_R7_reg_2 (.CK( clk ) , .D( u2_N225 ) , .Q( u2_R7_2 ) );
  DFF_X1 u2_R7_reg_20 (.CK( clk ) , .D( u2_N243 ) , .Q( u2_R7_20 ) );
  DFF_X1 u2_R7_reg_21 (.CK( clk ) , .D( u2_N244 ) , .Q( u2_R7_21 ) );
  DFF_X1 u2_R7_reg_22 (.CK( clk ) , .D( u2_N245 ) , .Q( u2_R7_22 ) );
  DFF_X1 u2_R7_reg_23 (.CK( clk ) , .D( u2_N246 ) , .Q( u2_R7_23 ) );
  DFF_X1 u2_R7_reg_24 (.CK( clk ) , .D( u2_N247 ) , .Q( u2_R7_24 ) );
  DFF_X1 u2_R7_reg_25 (.CK( clk ) , .D( u2_N248 ) , .Q( u2_R7_25 ) );
  DFF_X1 u2_R7_reg_26 (.CK( clk ) , .D( u2_N249 ) , .Q( u2_R7_26 ) );
  DFF_X1 u2_R7_reg_27 (.CK( clk ) , .D( u2_N250 ) , .Q( u2_R7_27 ) );
  DFF_X1 u2_R7_reg_28 (.CK( clk ) , .D( u2_N251 ) , .Q( u2_R7_28 ) );
  DFF_X1 u2_R7_reg_29 (.CK( clk ) , .D( u2_N252 ) , .Q( u2_R7_29 ) );
  DFF_X1 u2_R7_reg_3 (.CK( clk ) , .D( u2_N226 ) , .Q( u2_R7_3 ) );
  DFF_X1 u2_R7_reg_30 (.CK( clk ) , .D( u2_N253 ) , .Q( u2_R7_30 ) );
  DFF_X1 u2_R7_reg_31 (.CK( clk ) , .D( u2_N254 ) , .Q( u2_R7_31 ) );
  DFF_X1 u2_R7_reg_32 (.CK( clk ) , .D( u2_N255 ) , .Q( u2_R7_32 ) );
  DFF_X1 u2_R7_reg_4 (.CK( clk ) , .D( u2_N227 ) , .Q( u2_R7_4 ) );
  DFF_X1 u2_R7_reg_5 (.CK( clk ) , .D( u2_N228 ) , .Q( u2_R7_5 ) );
  DFF_X1 u2_R7_reg_6 (.CK( clk ) , .D( u2_N229 ) , .Q( u2_R7_6 ) );
  DFF_X1 u2_R7_reg_7 (.CK( clk ) , .D( u2_N230 ) , .Q( u2_R7_7 ) );
  DFF_X1 u2_R7_reg_8 (.CK( clk ) , .D( u2_N231 ) , .Q( u2_R7_8 ) );
  DFF_X1 u2_R7_reg_9 (.CK( clk ) , .D( u2_N232 ) , .Q( u2_R7_9 ) );
  DFF_X1 u2_R8_reg_1 (.CK( clk ) , .D( u2_N256 ) , .Q( u2_R8_1 ) );
  DFF_X1 u2_R8_reg_10 (.CK( clk ) , .D( u2_N265 ) , .Q( u2_R8_10 ) );
  DFF_X1 u2_R8_reg_11 (.CK( clk ) , .D( u2_N266 ) , .Q( u2_R8_11 ) );
  DFF_X1 u2_R8_reg_12 (.CK( clk ) , .D( u2_N267 ) , .Q( u2_R8_12 ) );
  DFF_X1 u2_R8_reg_13 (.CK( clk ) , .D( u2_N268 ) , .Q( u2_R8_13 ) );
  DFF_X1 u2_R8_reg_14 (.CK( clk ) , .D( u2_N269 ) , .Q( u2_R8_14 ) );
  DFF_X1 u2_R8_reg_15 (.CK( clk ) , .D( u2_N270 ) , .Q( u2_R8_15 ) );
  DFF_X1 u2_R8_reg_16 (.CK( clk ) , .D( u2_N271 ) , .Q( u2_R8_16 ) );
  DFF_X1 u2_R8_reg_17 (.CK( clk ) , .D( u2_N272 ) , .Q( u2_R8_17 ) );
  DFF_X1 u2_R8_reg_18 (.CK( clk ) , .D( u2_N273 ) , .Q( u2_R8_18 ) );
  DFF_X1 u2_R8_reg_19 (.CK( clk ) , .D( u2_N274 ) , .Q( u2_R8_19 ) );
  DFF_X1 u2_R8_reg_2 (.CK( clk ) , .D( u2_N257 ) , .Q( u2_R8_2 ) );
  DFF_X1 u2_R8_reg_20 (.CK( clk ) , .D( u2_N275 ) , .Q( u2_R8_20 ) );
  DFF_X1 u2_R8_reg_21 (.CK( clk ) , .D( u2_N276 ) , .Q( u2_R8_21 ) );
  DFF_X1 u2_R8_reg_22 (.CK( clk ) , .D( u2_N277 ) , .Q( u2_R8_22 ) );
  DFF_X1 u2_R8_reg_23 (.CK( clk ) , .D( u2_N278 ) , .Q( u2_R8_23 ) );
  DFF_X1 u2_R8_reg_24 (.CK( clk ) , .D( u2_N279 ) , .Q( u2_R8_24 ) );
  DFF_X1 u2_R8_reg_25 (.CK( clk ) , .D( u2_N280 ) , .Q( u2_R8_25 ) );
  DFF_X1 u2_R8_reg_26 (.CK( clk ) , .D( u2_N281 ) , .Q( u2_R8_26 ) );
  DFF_X1 u2_R8_reg_27 (.CK( clk ) , .D( u2_N282 ) , .Q( u2_R8_27 ) );
  DFF_X1 u2_R8_reg_28 (.CK( clk ) , .D( u2_N283 ) , .Q( u2_R8_28 ) );
  DFF_X1 u2_R8_reg_29 (.CK( clk ) , .D( u2_N284 ) , .Q( u2_R8_29 ) );
  DFF_X1 u2_R8_reg_3 (.CK( clk ) , .D( u2_N258 ) , .Q( u2_R8_3 ) );
  DFF_X1 u2_R8_reg_30 (.CK( clk ) , .D( u2_N285 ) , .Q( u2_R8_30 ) );
  DFF_X1 u2_R8_reg_31 (.CK( clk ) , .D( u2_N286 ) , .Q( u2_R8_31 ) );
  DFF_X1 u2_R8_reg_32 (.CK( clk ) , .D( u2_N287 ) , .Q( u2_R8_32 ) );
  DFF_X1 u2_R8_reg_4 (.CK( clk ) , .D( u2_N259 ) , .Q( u2_R8_4 ) );
  DFF_X1 u2_R8_reg_5 (.CK( clk ) , .D( u2_N260 ) , .Q( u2_R8_5 ) );
  DFF_X1 u2_R8_reg_6 (.CK( clk ) , .D( u2_N261 ) , .Q( u2_R8_6 ) );
  DFF_X1 u2_R8_reg_7 (.CK( clk ) , .D( u2_N262 ) , .Q( u2_R8_7 ) );
  DFF_X1 u2_R8_reg_8 (.CK( clk ) , .D( u2_N263 ) , .Q( u2_R8_8 ) );
  DFF_X1 u2_R8_reg_9 (.CK( clk ) , .D( u2_N264 ) , .Q( u2_R8_9 ) );
  DFF_X1 u2_R9_reg_1 (.CK( clk ) , .D( u2_N288 ) , .Q( u2_R9_1 ) );
  DFF_X1 u2_R9_reg_10 (.CK( clk ) , .D( u2_N297 ) , .Q( u2_R9_10 ) );
  DFF_X1 u2_R9_reg_11 (.CK( clk ) , .D( u2_N298 ) , .Q( u2_R9_11 ) );
  DFF_X1 u2_R9_reg_12 (.CK( clk ) , .D( u2_N299 ) , .Q( u2_R9_12 ) );
  DFF_X1 u2_R9_reg_13 (.CK( clk ) , .D( u2_N300 ) , .Q( u2_R9_13 ) );
  DFF_X1 u2_R9_reg_14 (.CK( clk ) , .D( u2_N301 ) , .Q( u2_R9_14 ) );
  DFF_X1 u2_R9_reg_15 (.CK( clk ) , .D( u2_N302 ) , .Q( u2_R9_15 ) );
  DFF_X1 u2_R9_reg_16 (.CK( clk ) , .D( u2_N303 ) , .Q( u2_R9_16 ) );
  DFF_X1 u2_R9_reg_17 (.CK( clk ) , .D( u2_N304 ) , .Q( u2_R9_17 ) );
  DFF_X1 u2_R9_reg_18 (.CK( clk ) , .D( u2_N305 ) , .Q( u2_R9_18 ) );
  DFF_X1 u2_R9_reg_19 (.CK( clk ) , .D( u2_N306 ) , .Q( u2_R9_19 ) );
  DFF_X1 u2_R9_reg_2 (.CK( clk ) , .D( u2_N289 ) , .Q( u2_R9_2 ) );
  DFF_X1 u2_R9_reg_20 (.CK( clk ) , .D( u2_N307 ) , .Q( u2_R9_20 ) );
  DFF_X1 u2_R9_reg_21 (.CK( clk ) , .D( u2_N308 ) , .Q( u2_R9_21 ) );
  DFF_X1 u2_R9_reg_22 (.CK( clk ) , .D( u2_N309 ) , .Q( u2_R9_22 ) );
  DFF_X1 u2_R9_reg_23 (.CK( clk ) , .D( u2_N310 ) , .Q( u2_R9_23 ) );
  DFF_X1 u2_R9_reg_24 (.CK( clk ) , .D( u2_N311 ) , .Q( u2_R9_24 ) );
  DFF_X1 u2_R9_reg_25 (.CK( clk ) , .D( u2_N312 ) , .Q( u2_R9_25 ) );
  DFF_X1 u2_R9_reg_26 (.CK( clk ) , .D( u2_N313 ) , .Q( u2_R9_26 ) );
  DFF_X1 u2_R9_reg_27 (.CK( clk ) , .D( u2_N314 ) , .Q( u2_R9_27 ) );
  DFF_X1 u2_R9_reg_28 (.CK( clk ) , .D( u2_N315 ) , .Q( u2_R9_28 ) );
  DFF_X1 u2_R9_reg_29 (.CK( clk ) , .D( u2_N316 ) , .Q( u2_R9_29 ) );
  DFF_X1 u2_R9_reg_3 (.CK( clk ) , .D( u2_N290 ) , .Q( u2_R9_3 ) );
  DFF_X1 u2_R9_reg_30 (.CK( clk ) , .D( u2_N317 ) , .Q( u2_R9_30 ) );
  DFF_X1 u2_R9_reg_31 (.CK( clk ) , .D( u2_N318 ) , .Q( u2_R9_31 ) );
  DFF_X1 u2_R9_reg_32 (.CK( clk ) , .D( u2_N319 ) , .Q( u2_R9_32 ) );
  DFF_X1 u2_R9_reg_4 (.CK( clk ) , .D( u2_N291 ) , .Q( u2_R9_4 ) );
  DFF_X1 u2_R9_reg_5 (.CK( clk ) , .D( u2_N292 ) , .Q( u2_R9_5 ) );
  DFF_X1 u2_R9_reg_6 (.CK( clk ) , .D( u2_N293 ) , .Q( u2_R9_6 ) );
  DFF_X1 u2_R9_reg_7 (.CK( clk ) , .D( u2_N294 ) , .Q( u2_R9_7 ) );
  DFF_X1 u2_R9_reg_8 (.CK( clk ) , .D( u2_N295 ) , .Q( u2_R9_8 ) );
  DFF_X1 u2_R9_reg_9 (.CK( clk ) , .D( u2_N296 ) , .Q( u2_R9_9 ) );
  XOR2_X1 u2_U10 (.B( u2_L1_29 ) , .Z( u2_N92 ) , .A( u2_out2_29 ) );
  XOR2_X1 u2_U100 (.B( u2_L12_27 ) , .Z( u2_N442 ) , .A( u2_out13_27 ) );
  XOR2_X1 u2_U101 (.B( u2_L12_26 ) , .Z( u2_N441 ) , .A( u2_out13_26 ) );
  XOR2_X1 u2_U102 (.B( u2_L12_25 ) , .Z( u2_N440 ) , .A( u2_out13_25 ) );
  XOR2_X1 u2_U103 (.B( u2_L0_13 ) , .Z( u2_N44 ) , .A( u2_out1_13 ) );
  XOR2_X1 u2_U104 (.B( u2_L12_24 ) , .Z( u2_N439 ) , .A( u2_out13_24 ) );
  XOR2_X1 u2_U105 (.B( u2_L12_23 ) , .Z( u2_N438 ) , .A( u2_out13_23 ) );
  XOR2_X1 u2_U106 (.B( u2_L12_22 ) , .Z( u2_N437 ) , .A( u2_out13_22 ) );
  XOR2_X1 u2_U107 (.B( u2_L12_21 ) , .Z( u2_N436 ) , .A( u2_out13_21 ) );
  XOR2_X1 u2_U108 (.B( u2_L12_20 ) , .Z( u2_N435 ) , .A( u2_out13_20 ) );
  XOR2_X1 u2_U109 (.B( u2_L12_19 ) , .Z( u2_N434 ) , .A( u2_out13_19 ) );
  XOR2_X1 u2_U11 (.B( u2_L1_28 ) , .Z( u2_N91 ) , .A( u2_out2_28 ) );
  XOR2_X1 u2_U110 (.B( u2_L12_18 ) , .Z( u2_N433 ) , .A( u2_out13_18 ) );
  XOR2_X1 u2_U111 (.B( u2_L12_17 ) , .Z( u2_N432 ) , .A( u2_out13_17 ) );
  XOR2_X1 u2_U112 (.B( u2_L12_16 ) , .Z( u2_N431 ) , .A( u2_out13_16 ) );
  XOR2_X1 u2_U113 (.B( u2_L12_15 ) , .Z( u2_N430 ) , .A( u2_out13_15 ) );
  XOR2_X1 u2_U114 (.B( u2_L0_12 ) , .Z( u2_N43 ) , .A( u2_out1_12 ) );
  XOR2_X1 u2_U115 (.B( u2_L12_14 ) , .Z( u2_N429 ) , .A( u2_out13_14 ) );
  XOR2_X1 u2_U116 (.B( u2_L12_13 ) , .Z( u2_N428 ) , .A( u2_out13_13 ) );
  XOR2_X1 u2_U117 (.B( u2_L12_12 ) , .Z( u2_N427 ) , .A( u2_out13_12 ) );
  XOR2_X1 u2_U118 (.B( u2_L12_11 ) , .Z( u2_N426 ) , .A( u2_out13_11 ) );
  XOR2_X1 u2_U119 (.B( u2_L12_10 ) , .Z( u2_N425 ) , .A( u2_out13_10 ) );
  XOR2_X1 u2_U12 (.B( u2_L1_27 ) , .Z( u2_N90 ) , .A( u2_out2_27 ) );
  XOR2_X1 u2_U120 (.B( u2_L12_9 ) , .Z( u2_N424 ) , .A( u2_out13_9 ) );
  XOR2_X1 u2_U121 (.B( u2_L12_8 ) , .Z( u2_N423 ) , .A( u2_out13_8 ) );
  XOR2_X1 u2_U122 (.B( u2_L12_7 ) , .Z( u2_N422 ) , .A( u2_out13_7 ) );
  XOR2_X1 u2_U123 (.B( u2_L12_6 ) , .Z( u2_N421 ) , .A( u2_out13_6 ) );
  XOR2_X1 u2_U124 (.B( u2_L12_5 ) , .Z( u2_N420 ) , .A( u2_out13_5 ) );
  XOR2_X1 u2_U125 (.B( u2_L0_11 ) , .Z( u2_N42 ) , .A( u2_out1_11 ) );
  XOR2_X1 u2_U126 (.B( u2_L12_4 ) , .Z( u2_N419 ) , .A( u2_out13_4 ) );
  XOR2_X1 u2_U127 (.B( u2_L12_3 ) , .Z( u2_N418 ) , .A( u2_out13_3 ) );
  XOR2_X1 u2_U128 (.B( u2_L12_2 ) , .Z( u2_N417 ) , .A( u2_out13_2 ) );
  XOR2_X1 u2_U129 (.B( u2_L12_1 ) , .Z( u2_N416 ) , .A( u2_out13_1 ) );
  XOR2_X1 u2_U13 (.Z( u2_N9 ) , .B( u2_desIn_r_12 ) , .A( u2_out0_10 ) );
  XOR2_X1 u2_U130 (.B( u2_L11_32 ) , .Z( u2_N415 ) , .A( u2_out12_32 ) );
  XOR2_X1 u2_U131 (.B( u2_L11_31 ) , .Z( u2_N414 ) , .A( u2_out12_31 ) );
  XOR2_X1 u2_U132 (.B( u2_L11_30 ) , .Z( u2_N413 ) , .A( u2_out12_30 ) );
  XOR2_X1 u2_U133 (.B( u2_L11_29 ) , .Z( u2_N412 ) , .A( u2_out12_29 ) );
  XOR2_X1 u2_U134 (.B( u2_L11_28 ) , .Z( u2_N411 ) , .A( u2_out12_28 ) );
  XOR2_X1 u2_U135 (.B( u2_L11_27 ) , .Z( u2_N410 ) , .A( u2_out12_27 ) );
  XOR2_X1 u2_U136 (.B( u2_L0_10 ) , .Z( u2_N41 ) , .A( u2_out1_10 ) );
  XOR2_X1 u2_U137 (.B( u2_L11_26 ) , .Z( u2_N409 ) , .A( u2_out12_26 ) );
  XOR2_X1 u2_U138 (.B( u2_L11_25 ) , .Z( u2_N408 ) , .A( u2_out12_25 ) );
  XOR2_X1 u2_U139 (.B( u2_L11_24 ) , .Z( u2_N407 ) , .A( u2_out12_24 ) );
  XOR2_X1 u2_U14 (.B( u2_L1_26 ) , .Z( u2_N89 ) , .A( u2_out2_26 ) );
  XOR2_X1 u2_U140 (.B( u2_L11_23 ) , .Z( u2_N406 ) , .A( u2_out12_23 ) );
  XOR2_X1 u2_U141 (.B( u2_L11_22 ) , .Z( u2_N405 ) , .A( u2_out12_22 ) );
  XOR2_X1 u2_U142 (.B( u2_L11_21 ) , .Z( u2_N404 ) , .A( u2_out12_21 ) );
  XOR2_X1 u2_U143 (.B( u2_L11_20 ) , .Z( u2_N403 ) , .A( u2_out12_20 ) );
  XOR2_X1 u2_U144 (.B( u2_L11_19 ) , .Z( u2_N402 ) , .A( u2_out12_19 ) );
  XOR2_X1 u2_U145 (.B( u2_L11_18 ) , .Z( u2_N401 ) , .A( u2_out12_18 ) );
  XOR2_X1 u2_U146 (.B( u2_L11_17 ) , .Z( u2_N400 ) , .A( u2_out12_17 ) );
  XOR2_X1 u2_U147 (.B( u2_L0_9 ) , .Z( u2_N40 ) , .A( u2_out1_9 ) );
  XOR2_X1 u2_U148 (.Z( u2_N4 ) , .B( u2_desIn_r_38 ) , .A( u2_out0_5 ) );
  XOR2_X1 u2_U149 (.B( u2_L11_16 ) , .Z( u2_N399 ) , .A( u2_out12_16 ) );
  XOR2_X1 u2_U15 (.B( u2_L1_25 ) , .Z( u2_N88 ) , .A( u2_out2_25 ) );
  XOR2_X1 u2_U150 (.B( u2_L11_15 ) , .Z( u2_N398 ) , .A( u2_out12_15 ) );
  XOR2_X1 u2_U151 (.B( u2_L11_14 ) , .Z( u2_N397 ) , .A( u2_out12_14 ) );
  XOR2_X1 u2_U152 (.B( u2_L11_13 ) , .Z( u2_N396 ) , .A( u2_out12_13 ) );
  XOR2_X1 u2_U153 (.B( u2_L11_12 ) , .Z( u2_N395 ) , .A( u2_out12_12 ) );
  XOR2_X1 u2_U154 (.B( u2_L11_11 ) , .Z( u2_N394 ) , .A( u2_out12_11 ) );
  XOR2_X1 u2_U155 (.B( u2_L11_10 ) , .Z( u2_N393 ) , .A( u2_out12_10 ) );
  XOR2_X1 u2_U156 (.B( u2_L11_9 ) , .Z( u2_N392 ) , .A( u2_out12_9 ) );
  XOR2_X1 u2_U157 (.B( u2_L11_8 ) , .Z( u2_N391 ) , .A( u2_out12_8 ) );
  XOR2_X1 u2_U158 (.B( u2_L11_7 ) , .Z( u2_N390 ) , .A( u2_out12_7 ) );
  XOR2_X1 u2_U159 (.B( u2_L0_8 ) , .Z( u2_N39 ) , .A( u2_out1_8 ) );
  XOR2_X1 u2_U16 (.B( u2_L1_24 ) , .Z( u2_N87 ) , .A( u2_out2_24 ) );
  XOR2_X1 u2_U160 (.B( u2_L11_6 ) , .Z( u2_N389 ) , .A( u2_out12_6 ) );
  XOR2_X1 u2_U161 (.B( u2_L11_5 ) , .Z( u2_N388 ) , .A( u2_out12_5 ) );
  XOR2_X1 u2_U162 (.B( u2_L11_4 ) , .Z( u2_N387 ) , .A( u2_out12_4 ) );
  XOR2_X1 u2_U163 (.B( u2_L11_3 ) , .Z( u2_N386 ) , .A( u2_out12_3 ) );
  XOR2_X1 u2_U164 (.B( u2_L11_2 ) , .Z( u2_N385 ) , .A( u2_out12_2 ) );
  XOR2_X1 u2_U165 (.B( u2_L11_1 ) , .Z( u2_N384 ) , .A( u2_out12_1 ) );
  XOR2_X1 u2_U166 (.B( u2_L10_32 ) , .Z( u2_N383 ) , .A( u2_out11_32 ) );
  XOR2_X1 u2_U167 (.B( u2_L10_31 ) , .Z( u2_N382 ) , .A( u2_out11_31 ) );
  XOR2_X1 u2_U168 (.B( u2_L10_30 ) , .Z( u2_N381 ) , .A( u2_out11_30 ) );
  XOR2_X1 u2_U169 (.B( u2_L10_29 ) , .Z( u2_N380 ) , .A( u2_out11_29 ) );
  XOR2_X1 u2_U17 (.B( u2_L1_23 ) , .Z( u2_N86 ) , .A( u2_out2_23 ) );
  XOR2_X1 u2_U170 (.B( u2_L0_7 ) , .Z( u2_N38 ) , .A( u2_out1_7 ) );
  XOR2_X1 u2_U171 (.B( u2_L10_28 ) , .Z( u2_N379 ) , .A( u2_out11_28 ) );
  XOR2_X1 u2_U172 (.B( u2_L10_27 ) , .Z( u2_N378 ) , .A( u2_out11_27 ) );
  XOR2_X1 u2_U173 (.B( u2_L10_26 ) , .Z( u2_N377 ) , .A( u2_out11_26 ) );
  XOR2_X1 u2_U174 (.B( u2_L10_25 ) , .Z( u2_N376 ) , .A( u2_out11_25 ) );
  XOR2_X1 u2_U175 (.B( u2_L10_24 ) , .Z( u2_N375 ) , .A( u2_out11_24 ) );
  XOR2_X1 u2_U176 (.B( u2_L10_23 ) , .Z( u2_N374 ) , .A( u2_out11_23 ) );
  XOR2_X1 u2_U177 (.B( u2_L10_22 ) , .Z( u2_N373 ) , .A( u2_out11_22 ) );
  XOR2_X1 u2_U178 (.B( u2_L10_21 ) , .Z( u2_N372 ) , .A( u2_out11_21 ) );
  XOR2_X1 u2_U179 (.B( u2_L10_20 ) , .Z( u2_N371 ) , .A( u2_out11_20 ) );
  XOR2_X1 u2_U18 (.B( u2_L1_22 ) , .Z( u2_N85 ) , .A( u2_out2_22 ) );
  XOR2_X1 u2_U180 (.B( u2_L10_19 ) , .Z( u2_N370 ) , .A( u2_out11_19 ) );
  XOR2_X1 u2_U181 (.B( u2_L0_6 ) , .Z( u2_N37 ) , .A( u2_out1_6 ) );
  XOR2_X1 u2_U182 (.B( u2_L10_18 ) , .Z( u2_N369 ) , .A( u2_out11_18 ) );
  XOR2_X1 u2_U183 (.B( u2_L10_17 ) , .Z( u2_N368 ) , .A( u2_out11_17 ) );
  XOR2_X1 u2_U184 (.B( u2_L10_16 ) , .Z( u2_N367 ) , .A( u2_out11_16 ) );
  XOR2_X1 u2_U185 (.B( u2_L10_15 ) , .Z( u2_N366 ) , .A( u2_out11_15 ) );
  XOR2_X1 u2_U186 (.B( u2_L10_14 ) , .Z( u2_N365 ) , .A( u2_out11_14 ) );
  XOR2_X1 u2_U187 (.B( u2_L10_13 ) , .Z( u2_N364 ) , .A( u2_out11_13 ) );
  XOR2_X1 u2_U188 (.B( u2_L10_12 ) , .Z( u2_N363 ) , .A( u2_out11_12 ) );
  XOR2_X1 u2_U189 (.B( u2_L10_11 ) , .Z( u2_N362 ) , .A( u2_out11_11 ) );
  XOR2_X1 u2_U19 (.B( u2_L1_21 ) , .Z( u2_N84 ) , .A( u2_out2_21 ) );
  XOR2_X1 u2_U190 (.B( u2_L10_10 ) , .Z( u2_N361 ) , .A( u2_out11_10 ) );
  XOR2_X1 u2_U191 (.B( u2_L10_9 ) , .Z( u2_N360 ) , .A( u2_out11_9 ) );
  XOR2_X1 u2_U192 (.B( u2_L0_5 ) , .Z( u2_N36 ) , .A( u2_out1_5 ) );
  XOR2_X1 u2_U193 (.B( u2_L10_8 ) , .Z( u2_N359 ) , .A( u2_out11_8 ) );
  XOR2_X1 u2_U194 (.B( u2_L10_7 ) , .Z( u2_N358 ) , .A( u2_out11_7 ) );
  XOR2_X1 u2_U195 (.B( u2_L10_6 ) , .Z( u2_N357 ) , .A( u2_out11_6 ) );
  XOR2_X1 u2_U196 (.B( u2_L10_5 ) , .Z( u2_N356 ) , .A( u2_out11_5 ) );
  XOR2_X1 u2_U197 (.B( u2_L10_4 ) , .Z( u2_N355 ) , .A( u2_out11_4 ) );
  XOR2_X1 u2_U198 (.B( u2_L10_3 ) , .Z( u2_N354 ) , .A( u2_out11_3 ) );
  XOR2_X1 u2_U199 (.B( u2_L10_2 ) , .Z( u2_N353 ) , .A( u2_out11_2 ) );
  XOR2_X1 u2_U20 (.B( u2_L1_20 ) , .Z( u2_N83 ) , .A( u2_out2_20 ) );
  XOR2_X1 u2_U200 (.B( u2_L10_1 ) , .Z( u2_N352 ) , .A( u2_out11_1 ) );
  XOR2_X1 u2_U201 (.B( u2_L9_32 ) , .Z( u2_N351 ) , .A( u2_out10_32 ) );
  XOR2_X1 u2_U202 (.B( u2_L9_31 ) , .Z( u2_N350 ) , .A( u2_out10_31 ) );
  XOR2_X1 u2_U203 (.B( u2_L0_4 ) , .Z( u2_N35 ) , .A( u2_out1_4 ) );
  XOR2_X1 u2_U204 (.B( u2_L9_30 ) , .Z( u2_N349 ) , .A( u2_out10_30 ) );
  XOR2_X1 u2_U205 (.B( u2_L9_29 ) , .Z( u2_N348 ) , .A( u2_out10_29 ) );
  XOR2_X1 u2_U206 (.B( u2_L9_28 ) , .Z( u2_N347 ) , .A( u2_out10_28 ) );
  XOR2_X1 u2_U207 (.B( u2_L9_27 ) , .Z( u2_N346 ) , .A( u2_out10_27 ) );
  XOR2_X1 u2_U208 (.B( u2_L9_26 ) , .Z( u2_N345 ) , .A( u2_out10_26 ) );
  XOR2_X1 u2_U209 (.B( u2_L9_25 ) , .Z( u2_N344 ) , .A( u2_out10_25 ) );
  XOR2_X1 u2_U21 (.B( u2_L1_19 ) , .Z( u2_N82 ) , .A( u2_out2_19 ) );
  XOR2_X1 u2_U210 (.B( u2_L9_24 ) , .Z( u2_N343 ) , .A( u2_out10_24 ) );
  XOR2_X1 u2_U211 (.B( u2_L9_23 ) , .Z( u2_N342 ) , .A( u2_out10_23 ) );
  XOR2_X1 u2_U212 (.B( u2_L9_22 ) , .Z( u2_N341 ) , .A( u2_out10_22 ) );
  XOR2_X1 u2_U213 (.B( u2_L9_21 ) , .Z( u2_N340 ) , .A( u2_out10_21 ) );
  XOR2_X1 u2_U214 (.B( u2_L0_3 ) , .Z( u2_N34 ) , .A( u2_out1_3 ) );
  XOR2_X1 u2_U215 (.B( u2_L9_20 ) , .Z( u2_N339 ) , .A( u2_out10_20 ) );
  XOR2_X1 u2_U216 (.B( u2_L9_19 ) , .Z( u2_N338 ) , .A( u2_out10_19 ) );
  XOR2_X1 u2_U217 (.B( u2_L9_18 ) , .Z( u2_N337 ) , .A( u2_out10_18 ) );
  XOR2_X1 u2_U218 (.B( u2_L9_17 ) , .Z( u2_N336 ) , .A( u2_out10_17 ) );
  XOR2_X1 u2_U219 (.B( u2_L9_16 ) , .Z( u2_N335 ) , .A( u2_out10_16 ) );
  XOR2_X1 u2_U22 (.B( u2_L1_18 ) , .Z( u2_N81 ) , .A( u2_out2_18 ) );
  XOR2_X1 u2_U220 (.B( u2_L9_15 ) , .Z( u2_N334 ) , .A( u2_out10_15 ) );
  XOR2_X1 u2_U221 (.B( u2_L9_14 ) , .Z( u2_N333 ) , .A( u2_out10_14 ) );
  XOR2_X1 u2_U222 (.B( u2_L9_13 ) , .Z( u2_N332 ) , .A( u2_out10_13 ) );
  XOR2_X1 u2_U223 (.B( u2_L9_12 ) , .Z( u2_N331 ) , .A( u2_out10_12 ) );
  XOR2_X1 u2_U224 (.B( u2_L9_11 ) , .Z( u2_N330 ) , .A( u2_out10_11 ) );
  XOR2_X1 u2_U225 (.B( u2_L0_2 ) , .Z( u2_N33 ) , .A( u2_out1_2 ) );
  XOR2_X1 u2_U226 (.B( u2_L9_10 ) , .Z( u2_N329 ) , .A( u2_out10_10 ) );
  XOR2_X1 u2_U227 (.B( u2_L9_9 ) , .Z( u2_N328 ) , .A( u2_out10_9 ) );
  XOR2_X1 u2_U228 (.B( u2_L9_8 ) , .Z( u2_N327 ) , .A( u2_out10_8 ) );
  XOR2_X1 u2_U229 (.B( u2_L9_7 ) , .Z( u2_N326 ) , .A( u2_out10_7 ) );
  XOR2_X1 u2_U23 (.B( u2_L1_17 ) , .Z( u2_N80 ) , .A( u2_out2_17 ) );
  XOR2_X1 u2_U230 (.B( u2_L9_6 ) , .Z( u2_N325 ) , .A( u2_out10_6 ) );
  XOR2_X1 u2_U231 (.B( u2_L9_5 ) , .Z( u2_N324 ) , .A( u2_out10_5 ) );
  XOR2_X1 u2_U232 (.B( u2_L9_4 ) , .Z( u2_N323 ) , .A( u2_out10_4 ) );
  XOR2_X1 u2_U233 (.B( u2_L9_3 ) , .Z( u2_N322 ) , .A( u2_out10_3 ) );
  XOR2_X1 u2_U234 (.B( u2_L9_2 ) , .Z( u2_N321 ) , .A( u2_out10_2 ) );
  XOR2_X1 u2_U235 (.B( u2_L9_1 ) , .Z( u2_N320 ) , .A( u2_out10_1 ) );
  XOR2_X1 u2_U236 (.B( u2_L0_1 ) , .Z( u2_N32 ) , .A( u2_out1_1 ) );
  XOR2_X1 u2_U237 (.B( u2_L8_32 ) , .Z( u2_N319 ) , .A( u2_out9_32 ) );
  XOR2_X1 u2_U238 (.B( u2_L8_31 ) , .Z( u2_N318 ) , .A( u2_out9_31 ) );
  XOR2_X1 u2_U239 (.B( u2_L8_30 ) , .Z( u2_N317 ) , .A( u2_out9_30 ) );
  XOR2_X1 u2_U24 (.Z( u2_N8 ) , .B( u2_desIn_r_4 ) , .A( u2_out0_9 ) );
  XOR2_X1 u2_U240 (.B( u2_L8_29 ) , .Z( u2_N316 ) , .A( u2_out9_29 ) );
  XOR2_X1 u2_U241 (.B( u2_L8_28 ) , .Z( u2_N315 ) , .A( u2_out9_28 ) );
  XOR2_X1 u2_U242 (.B( u2_L8_27 ) , .Z( u2_N314 ) , .A( u2_out9_27 ) );
  XOR2_X1 u2_U243 (.B( u2_L8_26 ) , .Z( u2_N313 ) , .A( u2_out9_26 ) );
  XOR2_X1 u2_U244 (.B( u2_L8_25 ) , .Z( u2_N312 ) , .A( u2_out9_25 ) );
  XOR2_X1 u2_U245 (.B( u2_L8_24 ) , .Z( u2_N311 ) , .A( u2_out9_24 ) );
  XOR2_X1 u2_U246 (.B( u2_L8_23 ) , .Z( u2_N310 ) , .A( u2_out9_23 ) );
  XOR2_X1 u2_U247 (.Z( u2_N31 ) , .B( u2_desIn_r_56 ) , .A( u2_out0_32 ) );
  XOR2_X1 u2_U248 (.B( u2_L8_22 ) , .Z( u2_N309 ) , .A( u2_out9_22 ) );
  XOR2_X1 u2_U249 (.B( u2_L8_21 ) , .Z( u2_N308 ) , .A( u2_out9_21 ) );
  XOR2_X1 u2_U25 (.B( u2_L1_16 ) , .Z( u2_N79 ) , .A( u2_out2_16 ) );
  XOR2_X1 u2_U250 (.B( u2_L8_20 ) , .Z( u2_N307 ) , .A( u2_out9_20 ) );
  XOR2_X1 u2_U251 (.B( u2_L8_19 ) , .Z( u2_N306 ) , .A( u2_out9_19 ) );
  XOR2_X1 u2_U252 (.B( u2_L8_18 ) , .Z( u2_N305 ) , .A( u2_out9_18 ) );
  XOR2_X1 u2_U253 (.B( u2_L8_17 ) , .Z( u2_N304 ) , .A( u2_out9_17 ) );
  XOR2_X1 u2_U254 (.B( u2_L8_16 ) , .Z( u2_N303 ) , .A( u2_out9_16 ) );
  XOR2_X1 u2_U255 (.B( u2_L8_15 ) , .Z( u2_N302 ) , .A( u2_out9_15 ) );
  XOR2_X1 u2_U256 (.B( u2_L8_14 ) , .Z( u2_N301 ) , .A( u2_out9_14 ) );
  XOR2_X1 u2_U257 (.B( u2_L8_13 ) , .Z( u2_N300 ) , .A( u2_out9_13 ) );
  XOR2_X1 u2_U258 (.Z( u2_N30 ) , .B( u2_desIn_r_48 ) , .A( u2_out0_31 ) );
  XOR2_X1 u2_U259 (.Z( u2_N3 ) , .B( u2_desIn_r_30 ) , .A( u2_out0_4 ) );
  XOR2_X1 u2_U26 (.B( u2_L1_15 ) , .Z( u2_N78 ) , .A( u2_out2_15 ) );
  XOR2_X1 u2_U260 (.B( u2_L8_12 ) , .Z( u2_N299 ) , .A( u2_out9_12 ) );
  XOR2_X1 u2_U261 (.B( u2_L8_11 ) , .Z( u2_N298 ) , .A( u2_out9_11 ) );
  XOR2_X1 u2_U262 (.B( u2_L8_10 ) , .Z( u2_N297 ) , .A( u2_out9_10 ) );
  XOR2_X1 u2_U263 (.B( u2_L8_9 ) , .Z( u2_N296 ) , .A( u2_out9_9 ) );
  XOR2_X1 u2_U264 (.B( u2_L8_8 ) , .Z( u2_N295 ) , .A( u2_out9_8 ) );
  XOR2_X1 u2_U265 (.B( u2_L8_7 ) , .Z( u2_N294 ) , .A( u2_out9_7 ) );
  XOR2_X1 u2_U266 (.B( u2_L8_6 ) , .Z( u2_N293 ) , .A( u2_out9_6 ) );
  XOR2_X1 u2_U267 (.B( u2_L8_5 ) , .Z( u2_N292 ) , .A( u2_out9_5 ) );
  XOR2_X1 u2_U268 (.B( u2_L8_4 ) , .Z( u2_N291 ) , .A( u2_out9_4 ) );
  XOR2_X1 u2_U269 (.B( u2_L8_3 ) , .Z( u2_N290 ) , .A( u2_out9_3 ) );
  XOR2_X1 u2_U27 (.B( u2_L1_14 ) , .Z( u2_N77 ) , .A( u2_out2_14 ) );
  XOR2_X1 u2_U270 (.Z( u2_N29 ) , .B( u2_desIn_r_40 ) , .A( u2_out0_30 ) );
  XOR2_X1 u2_U271 (.B( u2_L8_2 ) , .Z( u2_N289 ) , .A( u2_out9_2 ) );
  XOR2_X1 u2_U272 (.B( u2_L8_1 ) , .Z( u2_N288 ) , .A( u2_out9_1 ) );
  XOR2_X1 u2_U273 (.B( u2_L7_32 ) , .Z( u2_N287 ) , .A( u2_out8_32 ) );
  XOR2_X1 u2_U274 (.B( u2_L7_31 ) , .Z( u2_N286 ) , .A( u2_out8_31 ) );
  XOR2_X1 u2_U275 (.B( u2_L7_30 ) , .Z( u2_N285 ) , .A( u2_out8_30 ) );
  XOR2_X1 u2_U276 (.B( u2_L7_29 ) , .Z( u2_N284 ) , .A( u2_out8_29 ) );
  XOR2_X1 u2_U277 (.B( u2_L7_28 ) , .Z( u2_N283 ) , .A( u2_out8_28 ) );
  XOR2_X1 u2_U278 (.B( u2_L7_27 ) , .Z( u2_N282 ) , .A( u2_out8_27 ) );
  XOR2_X1 u2_U279 (.B( u2_L7_26 ) , .Z( u2_N281 ) , .A( u2_out8_26 ) );
  XOR2_X1 u2_U28 (.B( u2_L1_13 ) , .Z( u2_N76 ) , .A( u2_out2_13 ) );
  XOR2_X1 u2_U280 (.B( u2_L7_25 ) , .Z( u2_N280 ) , .A( u2_out8_25 ) );
  XOR2_X1 u2_U281 (.Z( u2_N28 ) , .B( u2_desIn_r_32 ) , .A( u2_out0_29 ) );
  XOR2_X1 u2_U282 (.B( u2_L7_24 ) , .Z( u2_N279 ) , .A( u2_out8_24 ) );
  XOR2_X1 u2_U283 (.B( u2_L7_23 ) , .Z( u2_N278 ) , .A( u2_out8_23 ) );
  XOR2_X1 u2_U284 (.B( u2_L7_22 ) , .Z( u2_N277 ) , .A( u2_out8_22 ) );
  XOR2_X1 u2_U285 (.B( u2_L7_21 ) , .Z( u2_N276 ) , .A( u2_out8_21 ) );
  XOR2_X1 u2_U286 (.B( u2_L7_20 ) , .Z( u2_N275 ) , .A( u2_out8_20 ) );
  XOR2_X1 u2_U287 (.B( u2_L7_19 ) , .Z( u2_N274 ) , .A( u2_out8_19 ) );
  XOR2_X1 u2_U288 (.B( u2_L7_18 ) , .Z( u2_N273 ) , .A( u2_out8_18 ) );
  XOR2_X1 u2_U289 (.B( u2_L7_17 ) , .Z( u2_N272 ) , .A( u2_out8_17 ) );
  XOR2_X1 u2_U29 (.B( u2_L1_12 ) , .Z( u2_N75 ) , .A( u2_out2_12 ) );
  XOR2_X1 u2_U290 (.B( u2_L7_16 ) , .Z( u2_N271 ) , .A( u2_out8_16 ) );
  XOR2_X1 u2_U291 (.B( u2_L7_15 ) , .Z( u2_N270 ) , .A( u2_out8_15 ) );
  XOR2_X1 u2_U292 (.Z( u2_N27 ) , .B( u2_desIn_r_24 ) , .A( u2_out0_28 ) );
  XOR2_X1 u2_U293 (.B( u2_L7_14 ) , .Z( u2_N269 ) , .A( u2_out8_14 ) );
  XOR2_X1 u2_U294 (.B( u2_L7_13 ) , .Z( u2_N268 ) , .A( u2_out8_13 ) );
  XOR2_X1 u2_U295 (.B( u2_L7_12 ) , .Z( u2_N267 ) , .A( u2_out8_12 ) );
  XOR2_X1 u2_U296 (.B( u2_L7_11 ) , .Z( u2_N266 ) , .A( u2_out8_11 ) );
  XOR2_X1 u2_U297 (.B( u2_L7_10 ) , .Z( u2_N265 ) , .A( u2_out8_10 ) );
  XOR2_X1 u2_U298 (.B( u2_L7_9 ) , .Z( u2_N264 ) , .A( u2_out8_9 ) );
  XOR2_X1 u2_U299 (.B( u2_L7_8 ) , .Z( u2_N263 ) , .A( u2_out8_8 ) );
  XOR2_X1 u2_U3 (.B( u2_L2_4 ) , .Z( u2_N99 ) , .A( u2_out3_4 ) );
  XOR2_X1 u2_U30 (.B( u2_L1_11 ) , .Z( u2_N74 ) , .A( u2_out2_11 ) );
  XOR2_X1 u2_U300 (.B( u2_L7_7 ) , .Z( u2_N262 ) , .A( u2_out8_7 ) );
  XOR2_X1 u2_U301 (.B( u2_L7_6 ) , .Z( u2_N261 ) , .A( u2_out8_6 ) );
  XOR2_X1 u2_U302 (.B( u2_L7_5 ) , .Z( u2_N260 ) , .A( u2_out8_5 ) );
  XOR2_X1 u2_U303 (.Z( u2_N26 ) , .B( u2_desIn_r_16 ) , .A( u2_out0_27 ) );
  XOR2_X1 u2_U304 (.B( u2_L7_4 ) , .Z( u2_N259 ) , .A( u2_out8_4 ) );
  XOR2_X1 u2_U305 (.B( u2_L7_3 ) , .Z( u2_N258 ) , .A( u2_out8_3 ) );
  XOR2_X1 u2_U306 (.B( u2_L7_2 ) , .Z( u2_N257 ) , .A( u2_out8_2 ) );
  XOR2_X1 u2_U307 (.B( u2_L7_1 ) , .Z( u2_N256 ) , .A( u2_out8_1 ) );
  XOR2_X1 u2_U308 (.B( u2_L6_32 ) , .Z( u2_N255 ) , .A( u2_out7_32 ) );
  XOR2_X1 u2_U309 (.B( u2_L6_31 ) , .Z( u2_N254 ) , .A( u2_out7_31 ) );
  XOR2_X1 u2_U31 (.B( u2_L1_10 ) , .Z( u2_N73 ) , .A( u2_out2_10 ) );
  XOR2_X1 u2_U310 (.B( u2_L6_30 ) , .Z( u2_N253 ) , .A( u2_out7_30 ) );
  XOR2_X1 u2_U311 (.B( u2_L6_29 ) , .Z( u2_N252 ) , .A( u2_out7_29 ) );
  XOR2_X1 u2_U312 (.B( u2_L6_28 ) , .Z( u2_N251 ) , .A( u2_out7_28 ) );
  XOR2_X1 u2_U313 (.B( u2_L6_27 ) , .Z( u2_N250 ) , .A( u2_out7_27 ) );
  XOR2_X1 u2_U314 (.Z( u2_N25 ) , .B( u2_desIn_r_8 ) , .A( u2_out0_26 ) );
  XOR2_X1 u2_U315 (.B( u2_L6_26 ) , .Z( u2_N249 ) , .A( u2_out7_26 ) );
  XOR2_X1 u2_U316 (.B( u2_L6_25 ) , .Z( u2_N248 ) , .A( u2_out7_25 ) );
  XOR2_X1 u2_U317 (.B( u2_L6_24 ) , .Z( u2_N247 ) , .A( u2_out7_24 ) );
  XOR2_X1 u2_U318 (.B( u2_L6_23 ) , .Z( u2_N246 ) , .A( u2_out7_23 ) );
  XOR2_X1 u2_U319 (.B( u2_L6_22 ) , .Z( u2_N245 ) , .A( u2_out7_22 ) );
  XOR2_X1 u2_U32 (.B( u2_L1_9 ) , .Z( u2_N72 ) , .A( u2_out2_9 ) );
  XOR2_X1 u2_U320 (.B( u2_L6_21 ) , .Z( u2_N244 ) , .A( u2_out7_21 ) );
  XOR2_X1 u2_U321 (.B( u2_L6_20 ) , .Z( u2_N243 ) , .A( u2_out7_20 ) );
  XOR2_X1 u2_U322 (.B( u2_L6_19 ) , .Z( u2_N242 ) , .A( u2_out7_19 ) );
  XOR2_X1 u2_U323 (.B( u2_L6_18 ) , .Z( u2_N241 ) , .A( u2_out7_18 ) );
  XOR2_X1 u2_U324 (.B( u2_L6_17 ) , .Z( u2_N240 ) , .A( u2_out7_17 ) );
  XOR2_X1 u2_U325 (.Z( u2_N24 ) , .B( u2_desIn_r_0 ) , .A( u2_out0_25 ) );
  XOR2_X1 u2_U326 (.B( u2_L6_16 ) , .Z( u2_N239 ) , .A( u2_out7_16 ) );
  XOR2_X1 u2_U327 (.B( u2_L6_15 ) , .Z( u2_N238 ) , .A( u2_out7_15 ) );
  XOR2_X1 u2_U328 (.B( u2_L6_14 ) , .Z( u2_N237 ) , .A( u2_out7_14 ) );
  XOR2_X1 u2_U329 (.B( u2_L6_13 ) , .Z( u2_N236 ) , .A( u2_out7_13 ) );
  XOR2_X1 u2_U33 (.B( u2_L1_8 ) , .Z( u2_N71 ) , .A( u2_out2_8 ) );
  XOR2_X1 u2_U330 (.B( u2_L6_12 ) , .Z( u2_N235 ) , .A( u2_out7_12 ) );
  XOR2_X1 u2_U331 (.B( u2_L6_11 ) , .Z( u2_N234 ) , .A( u2_out7_11 ) );
  XOR2_X1 u2_U332 (.B( u2_L6_10 ) , .Z( u2_N233 ) , .A( u2_out7_10 ) );
  XOR2_X1 u2_U333 (.B( u2_L6_9 ) , .Z( u2_N232 ) , .A( u2_out7_9 ) );
  XOR2_X1 u2_U334 (.B( u2_L6_8 ) , .Z( u2_N231 ) , .A( u2_out7_8 ) );
  XOR2_X1 u2_U335 (.B( u2_L6_7 ) , .Z( u2_N230 ) , .A( u2_out7_7 ) );
  XOR2_X1 u2_U336 (.Z( u2_N23 ) , .B( u2_desIn_r_58 ) , .A( u2_out0_24 ) );
  XOR2_X1 u2_U337 (.B( u2_L6_6 ) , .Z( u2_N229 ) , .A( u2_out7_6 ) );
  XOR2_X1 u2_U338 (.B( u2_L6_5 ) , .Z( u2_N228 ) , .A( u2_out7_5 ) );
  XOR2_X1 u2_U339 (.B( u2_L6_4 ) , .Z( u2_N227 ) , .A( u2_out7_4 ) );
  XOR2_X1 u2_U34 (.B( u2_L1_7 ) , .Z( u2_N70 ) , .A( u2_out2_7 ) );
  XOR2_X1 u2_U340 (.B( u2_L6_3 ) , .Z( u2_N226 ) , .A( u2_out7_3 ) );
  XOR2_X1 u2_U341 (.B( u2_L6_2 ) , .Z( u2_N225 ) , .A( u2_out7_2 ) );
  XOR2_X1 u2_U342 (.B( u2_L6_1 ) , .Z( u2_N224 ) , .A( u2_out7_1 ) );
  XOR2_X1 u2_U343 (.B( u2_L5_32 ) , .Z( u2_N223 ) , .A( u2_out6_32 ) );
  XOR2_X1 u2_U344 (.B( u2_L5_31 ) , .Z( u2_N222 ) , .A( u2_out6_31 ) );
  XOR2_X1 u2_U345 (.B( u2_L5_30 ) , .Z( u2_N221 ) , .A( u2_out6_30 ) );
  XOR2_X1 u2_U346 (.B( u2_L5_29 ) , .Z( u2_N220 ) , .A( u2_out6_29 ) );
  XOR2_X1 u2_U347 (.Z( u2_N22 ) , .B( u2_desIn_r_50 ) , .A( u2_out0_23 ) );
  XOR2_X1 u2_U348 (.B( u2_L5_28 ) , .Z( u2_N219 ) , .A( u2_out6_28 ) );
  XOR2_X1 u2_U349 (.B( u2_L5_27 ) , .Z( u2_N218 ) , .A( u2_out6_27 ) );
  XOR2_X1 u2_U35 (.Z( u2_N7 ) , .B( u2_desIn_r_62 ) , .A( u2_out0_8 ) );
  XOR2_X1 u2_U350 (.B( u2_L5_26 ) , .Z( u2_N217 ) , .A( u2_out6_26 ) );
  XOR2_X1 u2_U351 (.B( u2_L5_25 ) , .Z( u2_N216 ) , .A( u2_out6_25 ) );
  XOR2_X1 u2_U352 (.B( u2_L5_24 ) , .Z( u2_N215 ) , .A( u2_out6_24 ) );
  XOR2_X1 u2_U353 (.B( u2_L5_23 ) , .Z( u2_N214 ) , .A( u2_out6_23 ) );
  XOR2_X1 u2_U354 (.B( u2_L5_22 ) , .Z( u2_N213 ) , .A( u2_out6_22 ) );
  XOR2_X1 u2_U355 (.B( u2_L5_21 ) , .Z( u2_N212 ) , .A( u2_out6_21 ) );
  XOR2_X1 u2_U356 (.B( u2_L5_20 ) , .Z( u2_N211 ) , .A( u2_out6_20 ) );
  XOR2_X1 u2_U357 (.B( u2_L5_19 ) , .Z( u2_N210 ) , .A( u2_out6_19 ) );
  XOR2_X1 u2_U358 (.Z( u2_N21 ) , .B( u2_desIn_r_42 ) , .A( u2_out0_22 ) );
  XOR2_X1 u2_U359 (.B( u2_L5_18 ) , .Z( u2_N209 ) , .A( u2_out6_18 ) );
  XOR2_X1 u2_U36 (.B( u2_L1_6 ) , .Z( u2_N69 ) , .A( u2_out2_6 ) );
  XOR2_X1 u2_U360 (.B( u2_L5_17 ) , .Z( u2_N208 ) , .A( u2_out6_17 ) );
  XOR2_X1 u2_U361 (.B( u2_L5_16 ) , .Z( u2_N207 ) , .A( u2_out6_16 ) );
  XOR2_X1 u2_U362 (.B( u2_L5_15 ) , .Z( u2_N206 ) , .A( u2_out6_15 ) );
  XOR2_X1 u2_U363 (.B( u2_L5_14 ) , .Z( u2_N205 ) , .A( u2_out6_14 ) );
  XOR2_X1 u2_U364 (.B( u2_L5_13 ) , .Z( u2_N204 ) , .A( u2_out6_13 ) );
  XOR2_X1 u2_U365 (.B( u2_L5_12 ) , .Z( u2_N203 ) , .A( u2_out6_12 ) );
  XOR2_X1 u2_U366 (.B( u2_L5_11 ) , .Z( u2_N202 ) , .A( u2_out6_11 ) );
  XOR2_X1 u2_U367 (.B( u2_L5_10 ) , .Z( u2_N201 ) , .A( u2_out6_10 ) );
  XOR2_X1 u2_U368 (.B( u2_L5_9 ) , .Z( u2_N200 ) , .A( u2_out6_9 ) );
  XOR2_X1 u2_U369 (.Z( u2_N20 ) , .B( u2_desIn_r_34 ) , .A( u2_out0_21 ) );
  XOR2_X1 u2_U37 (.B( u2_L1_5 ) , .Z( u2_N68 ) , .A( u2_out2_5 ) );
  XOR2_X1 u2_U370 (.Z( u2_N2 ) , .B( u2_desIn_r_22 ) , .A( u2_out0_3 ) );
  XOR2_X1 u2_U371 (.B( u2_L5_8 ) , .Z( u2_N199 ) , .A( u2_out6_8 ) );
  XOR2_X1 u2_U372 (.B( u2_L5_7 ) , .Z( u2_N198 ) , .A( u2_out6_7 ) );
  XOR2_X1 u2_U373 (.B( u2_L5_6 ) , .Z( u2_N197 ) , .A( u2_out6_6 ) );
  XOR2_X1 u2_U374 (.B( u2_L5_5 ) , .Z( u2_N196 ) , .A( u2_out6_5 ) );
  XOR2_X1 u2_U375 (.B( u2_L5_4 ) , .Z( u2_N195 ) , .A( u2_out6_4 ) );
  XOR2_X1 u2_U376 (.B( u2_L5_3 ) , .Z( u2_N194 ) , .A( u2_out6_3 ) );
  XOR2_X1 u2_U377 (.B( u2_L5_2 ) , .Z( u2_N193 ) , .A( u2_out6_2 ) );
  XOR2_X1 u2_U378 (.B( u2_L5_1 ) , .Z( u2_N192 ) , .A( u2_out6_1 ) );
  XOR2_X1 u2_U379 (.B( u2_L4_32 ) , .Z( u2_N191 ) , .A( u2_out5_32 ) );
  XOR2_X1 u2_U38 (.B( u2_L1_4 ) , .Z( u2_N67 ) , .A( u2_out2_4 ) );
  XOR2_X1 u2_U380 (.B( u2_L4_31 ) , .Z( u2_N190 ) , .A( u2_out5_31 ) );
  XOR2_X1 u2_U381 (.Z( u2_N19 ) , .B( u2_desIn_r_26 ) , .A( u2_out0_20 ) );
  XOR2_X1 u2_U382 (.B( u2_L4_30 ) , .Z( u2_N189 ) , .A( u2_out5_30 ) );
  XOR2_X1 u2_U383 (.B( u2_L4_29 ) , .Z( u2_N188 ) , .A( u2_out5_29 ) );
  XOR2_X1 u2_U384 (.B( u2_L4_28 ) , .Z( u2_N187 ) , .A( u2_out5_28 ) );
  XOR2_X1 u2_U385 (.B( u2_L4_27 ) , .Z( u2_N186 ) , .A( u2_out5_27 ) );
  XOR2_X1 u2_U386 (.B( u2_L4_26 ) , .Z( u2_N185 ) , .A( u2_out5_26 ) );
  XOR2_X1 u2_U387 (.B( u2_L4_25 ) , .Z( u2_N184 ) , .A( u2_out5_25 ) );
  XOR2_X1 u2_U388 (.B( u2_L4_24 ) , .Z( u2_N183 ) , .A( u2_out5_24 ) );
  XOR2_X1 u2_U389 (.B( u2_L4_23 ) , .Z( u2_N182 ) , .A( u2_out5_23 ) );
  XOR2_X1 u2_U39 (.B( u2_L1_3 ) , .Z( u2_N66 ) , .A( u2_out2_3 ) );
  XOR2_X1 u2_U390 (.B( u2_L4_22 ) , .Z( u2_N181 ) , .A( u2_out5_22 ) );
  XOR2_X1 u2_U391 (.B( u2_L4_21 ) , .Z( u2_N180 ) , .A( u2_out5_21 ) );
  XOR2_X1 u2_U392 (.Z( u2_N18 ) , .B( u2_desIn_r_18 ) , .A( u2_out0_19 ) );
  XOR2_X1 u2_U393 (.B( u2_L4_20 ) , .Z( u2_N179 ) , .A( u2_out5_20 ) );
  XOR2_X1 u2_U394 (.B( u2_L4_19 ) , .Z( u2_N178 ) , .A( u2_out5_19 ) );
  XOR2_X1 u2_U395 (.B( u2_L4_18 ) , .Z( u2_N177 ) , .A( u2_out5_18 ) );
  XOR2_X1 u2_U396 (.B( u2_L4_17 ) , .Z( u2_N176 ) , .A( u2_out5_17 ) );
  XOR2_X1 u2_U397 (.B( u2_L4_16 ) , .Z( u2_N175 ) , .A( u2_out5_16 ) );
  XOR2_X1 u2_U398 (.B( u2_L4_15 ) , .Z( u2_N174 ) , .A( u2_out5_15 ) );
  XOR2_X1 u2_U399 (.B( u2_L4_14 ) , .Z( u2_N173 ) , .A( u2_out5_14 ) );
  XOR2_X1 u2_U4 (.B( u2_L2_3 ) , .Z( u2_N98 ) , .A( u2_out3_3 ) );
  XOR2_X1 u2_U40 (.B( u2_L1_2 ) , .Z( u2_N65 ) , .A( u2_out2_2 ) );
  XOR2_X1 u2_U400 (.B( u2_L4_13 ) , .Z( u2_N172 ) , .A( u2_out5_13 ) );
  XOR2_X1 u2_U401 (.B( u2_L4_12 ) , .Z( u2_N171 ) , .A( u2_out5_12 ) );
  XOR2_X1 u2_U402 (.B( u2_L4_11 ) , .Z( u2_N170 ) , .A( u2_out5_11 ) );
  XOR2_X1 u2_U403 (.Z( u2_N17 ) , .B( u2_desIn_r_10 ) , .A( u2_out0_18 ) );
  XOR2_X1 u2_U404 (.B( u2_L4_10 ) , .Z( u2_N169 ) , .A( u2_out5_10 ) );
  XOR2_X1 u2_U405 (.B( u2_L4_9 ) , .Z( u2_N168 ) , .A( u2_out5_9 ) );
  XOR2_X1 u2_U406 (.B( u2_L4_8 ) , .Z( u2_N167 ) , .A( u2_out5_8 ) );
  XOR2_X1 u2_U407 (.B( u2_L4_7 ) , .Z( u2_N166 ) , .A( u2_out5_7 ) );
  XOR2_X1 u2_U408 (.B( u2_L4_6 ) , .Z( u2_N165 ) , .A( u2_out5_6 ) );
  XOR2_X1 u2_U409 (.B( u2_L4_5 ) , .Z( u2_N164 ) , .A( u2_out5_5 ) );
  XOR2_X1 u2_U41 (.B( u2_L1_1 ) , .Z( u2_N64 ) , .A( u2_out2_1 ) );
  XOR2_X1 u2_U410 (.B( u2_L4_4 ) , .Z( u2_N163 ) , .A( u2_out5_4 ) );
  XOR2_X1 u2_U411 (.B( u2_L4_3 ) , .Z( u2_N162 ) , .A( u2_out5_3 ) );
  XOR2_X1 u2_U412 (.B( u2_L4_2 ) , .Z( u2_N161 ) , .A( u2_out5_2 ) );
  XOR2_X1 u2_U413 (.B( u2_L4_1 ) , .Z( u2_N160 ) , .A( u2_out5_1 ) );
  XOR2_X1 u2_U414 (.Z( u2_N16 ) , .B( u2_desIn_r_2 ) , .A( u2_out0_17 ) );
  XOR2_X1 u2_U415 (.B( u2_L3_32 ) , .Z( u2_N159 ) , .A( u2_out4_32 ) );
  XOR2_X1 u2_U416 (.B( u2_L3_31 ) , .Z( u2_N158 ) , .A( u2_out4_31 ) );
  XOR2_X1 u2_U417 (.B( u2_L3_30 ) , .Z( u2_N157 ) , .A( u2_out4_30 ) );
  XOR2_X1 u2_U418 (.B( u2_L3_29 ) , .Z( u2_N156 ) , .A( u2_out4_29 ) );
  XOR2_X1 u2_U419 (.B( u2_L3_28 ) , .Z( u2_N155 ) , .A( u2_out4_28 ) );
  XOR2_X1 u2_U42 (.B( u2_L0_32 ) , .Z( u2_N63 ) , .A( u2_out1_32 ) );
  XOR2_X1 u2_U420 (.B( u2_L3_27 ) , .Z( u2_N154 ) , .A( u2_out4_27 ) );
  XOR2_X1 u2_U421 (.B( u2_L3_26 ) , .Z( u2_N153 ) , .A( u2_out4_26 ) );
  XOR2_X1 u2_U422 (.B( u2_L3_25 ) , .Z( u2_N152 ) , .A( u2_out4_25 ) );
  XOR2_X1 u2_U423 (.B( u2_L3_24 ) , .Z( u2_N151 ) , .A( u2_out4_24 ) );
  XOR2_X1 u2_U424 (.B( u2_L3_23 ) , .Z( u2_N150 ) , .A( u2_out4_23 ) );
  XOR2_X1 u2_U425 (.Z( u2_N15 ) , .B( u2_desIn_r_60 ) , .A( u2_out0_16 ) );
  XOR2_X1 u2_U426 (.B( u2_L3_22 ) , .Z( u2_N149 ) , .A( u2_out4_22 ) );
  XOR2_X1 u2_U427 (.B( u2_L3_21 ) , .Z( u2_N148 ) , .A( u2_out4_21 ) );
  XOR2_X1 u2_U428 (.B( u2_L3_20 ) , .Z( u2_N147 ) , .A( u2_out4_20 ) );
  XOR2_X1 u2_U429 (.B( u2_L3_19 ) , .Z( u2_N146 ) , .A( u2_out4_19 ) );
  XOR2_X1 u2_U43 (.B( u2_L0_31 ) , .Z( u2_N62 ) , .A( u2_out1_31 ) );
  XOR2_X1 u2_U430 (.B( u2_L3_18 ) , .Z( u2_N145 ) , .A( u2_out4_18 ) );
  XOR2_X1 u2_U431 (.B( u2_L3_17 ) , .Z( u2_N144 ) , .A( u2_out4_17 ) );
  XOR2_X1 u2_U432 (.B( u2_L3_16 ) , .Z( u2_N143 ) , .A( u2_out4_16 ) );
  XOR2_X1 u2_U433 (.B( u2_L3_15 ) , .Z( u2_N142 ) , .A( u2_out4_15 ) );
  XOR2_X1 u2_U434 (.B( u2_L3_14 ) , .Z( u2_N141 ) , .A( u2_out4_14 ) );
  XOR2_X1 u2_U435 (.B( u2_L3_13 ) , .Z( u2_N140 ) , .A( u2_out4_13 ) );
  XOR2_X1 u2_U436 (.Z( u2_N14 ) , .B( u2_desIn_r_52 ) , .A( u2_out0_15 ) );
  XOR2_X1 u2_U437 (.B( u2_L3_12 ) , .Z( u2_N139 ) , .A( u2_out4_12 ) );
  XOR2_X1 u2_U438 (.B( u2_L3_11 ) , .Z( u2_N138 ) , .A( u2_out4_11 ) );
  XOR2_X1 u2_U439 (.B( u2_L3_10 ) , .Z( u2_N137 ) , .A( u2_out4_10 ) );
  XOR2_X1 u2_U44 (.B( u2_L0_30 ) , .Z( u2_N61 ) , .A( u2_out1_30 ) );
  XOR2_X1 u2_U440 (.B( u2_L3_9 ) , .Z( u2_N136 ) , .A( u2_out4_9 ) );
  XOR2_X1 u2_U441 (.B( u2_L3_8 ) , .Z( u2_N135 ) , .A( u2_out4_8 ) );
  XOR2_X1 u2_U442 (.B( u2_L3_7 ) , .Z( u2_N134 ) , .A( u2_out4_7 ) );
  XOR2_X1 u2_U443 (.B( u2_L3_6 ) , .Z( u2_N133 ) , .A( u2_out4_6 ) );
  XOR2_X1 u2_U444 (.B( u2_L3_5 ) , .Z( u2_N132 ) , .A( u2_out4_5 ) );
  XOR2_X1 u2_U445 (.B( u2_L3_4 ) , .Z( u2_N131 ) , .A( u2_out4_4 ) );
  XOR2_X1 u2_U446 (.B( u2_L3_3 ) , .Z( u2_N130 ) , .A( u2_out4_3 ) );
  XOR2_X1 u2_U447 (.Z( u2_N13 ) , .B( u2_desIn_r_44 ) , .A( u2_out0_14 ) );
  XOR2_X1 u2_U448 (.B( u2_L3_2 ) , .Z( u2_N129 ) , .A( u2_out4_2 ) );
  XOR2_X1 u2_U449 (.B( u2_L3_1 ) , .Z( u2_N128 ) , .A( u2_out4_1 ) );
  XOR2_X1 u2_U45 (.B( u2_L0_29 ) , .Z( u2_N60 ) , .A( u2_out1_29 ) );
  XOR2_X1 u2_U450 (.B( u2_L2_32 ) , .Z( u2_N127 ) , .A( u2_out3_32 ) );
  XOR2_X1 u2_U451 (.B( u2_L2_31 ) , .Z( u2_N126 ) , .A( u2_out3_31 ) );
  XOR2_X1 u2_U452 (.B( u2_L2_30 ) , .Z( u2_N125 ) , .A( u2_out3_30 ) );
  XOR2_X1 u2_U453 (.B( u2_L2_29 ) , .Z( u2_N124 ) , .A( u2_out3_29 ) );
  XOR2_X1 u2_U454 (.B( u2_L2_28 ) , .Z( u2_N123 ) , .A( u2_out3_28 ) );
  XOR2_X1 u2_U455 (.B( u2_L2_27 ) , .Z( u2_N122 ) , .A( u2_out3_27 ) );
  XOR2_X1 u2_U456 (.B( u2_L2_26 ) , .Z( u2_N121 ) , .A( u2_out3_26 ) );
  XOR2_X1 u2_U457 (.B( u2_L2_25 ) , .Z( u2_N120 ) , .A( u2_out3_25 ) );
  XOR2_X1 u2_U458 (.Z( u2_N12 ) , .B( u2_desIn_r_36 ) , .A( u2_out0_13 ) );
  XOR2_X1 u2_U459 (.B( u2_L2_24 ) , .Z( u2_N119 ) , .A( u2_out3_24 ) );
  XOR2_X1 u2_U46 (.Z( u2_N6 ) , .B( u2_desIn_r_54 ) , .A( u2_out0_7 ) );
  XOR2_X1 u2_U460 (.B( u2_L2_23 ) , .Z( u2_N118 ) , .A( u2_out3_23 ) );
  XOR2_X1 u2_U461 (.B( u2_L2_22 ) , .Z( u2_N117 ) , .A( u2_out3_22 ) );
  XOR2_X1 u2_U462 (.B( u2_L2_21 ) , .Z( u2_N116 ) , .A( u2_out3_21 ) );
  XOR2_X1 u2_U463 (.B( u2_L2_20 ) , .Z( u2_N115 ) , .A( u2_out3_20 ) );
  XOR2_X1 u2_U464 (.B( u2_L2_19 ) , .Z( u2_N114 ) , .A( u2_out3_19 ) );
  XOR2_X1 u2_U465 (.B( u2_L2_18 ) , .Z( u2_N113 ) , .A( u2_out3_18 ) );
  XOR2_X1 u2_U466 (.B( u2_L2_17 ) , .Z( u2_N112 ) , .A( u2_out3_17 ) );
  XOR2_X1 u2_U467 (.B( u2_L2_16 ) , .Z( u2_N111 ) , .A( u2_out3_16 ) );
  XOR2_X1 u2_U468 (.B( u2_L2_15 ) , .Z( u2_N110 ) , .A( u2_out3_15 ) );
  XOR2_X1 u2_U469 (.Z( u2_N11 ) , .B( u2_desIn_r_28 ) , .A( u2_out0_12 ) );
  XOR2_X1 u2_U47 (.B( u2_L0_28 ) , .Z( u2_N59 ) , .A( u2_out1_28 ) );
  XOR2_X1 u2_U470 (.B( u2_L2_14 ) , .Z( u2_N109 ) , .A( u2_out3_14 ) );
  XOR2_X1 u2_U471 (.B( u2_L2_13 ) , .Z( u2_N108 ) , .A( u2_out3_13 ) );
  XOR2_X1 u2_U472 (.B( u2_L2_12 ) , .Z( u2_N107 ) , .A( u2_out3_12 ) );
  XOR2_X1 u2_U473 (.B( u2_L2_11 ) , .Z( u2_N106 ) , .A( u2_out3_11 ) );
  XOR2_X1 u2_U474 (.B( u2_L2_10 ) , .Z( u2_N105 ) , .A( u2_out3_10 ) );
  XOR2_X1 u2_U475 (.B( u2_L2_9 ) , .Z( u2_N104 ) , .A( u2_out3_9 ) );
  XOR2_X1 u2_U476 (.B( u2_L2_8 ) , .Z( u2_N103 ) , .A( u2_out3_8 ) );
  XOR2_X1 u2_U477 (.B( u2_L2_7 ) , .Z( u2_N102 ) , .A( u2_out3_7 ) );
  XOR2_X1 u2_U478 (.B( u2_L2_6 ) , .Z( u2_N101 ) , .A( u2_out3_6 ) );
  XOR2_X1 u2_U479 (.B( u2_L2_5 ) , .Z( u2_N100 ) , .A( u2_out3_5 ) );
  XOR2_X1 u2_U48 (.B( u2_L0_27 ) , .Z( u2_N58 ) , .A( u2_out1_27 ) );
  XOR2_X1 u2_U480 (.Z( u2_N10 ) , .B( u2_desIn_r_20 ) , .A( u2_out0_11 ) );
  XOR2_X1 u2_U481 (.Z( u2_N1 ) , .B( u2_desIn_r_14 ) , .A( u2_out0_2 ) );
  XOR2_X1 u2_U482 (.Z( u2_N0 ) , .B( u2_desIn_r_6 ) , .A( u2_out0_1 ) );
  XOR2_X1 u2_U483 (.Z( u2_FP_9 ) , .B( u2_L14_9 ) , .A( u2_out15_9 ) );
  XOR2_X1 u2_U484 (.Z( u2_FP_8 ) , .B( u2_L14_8 ) , .A( u2_out15_8 ) );
  XOR2_X1 u2_U485 (.Z( u2_FP_7 ) , .B( u2_L14_7 ) , .A( u2_out15_7 ) );
  XOR2_X1 u2_U486 (.Z( u2_FP_6 ) , .B( u2_L14_6 ) , .A( u2_out15_6 ) );
  XOR2_X1 u2_U487 (.Z( u2_FP_5 ) , .B( u2_L14_5 ) , .A( u2_out15_5 ) );
  XOR2_X1 u2_U488 (.Z( u2_FP_4 ) , .B( u2_L14_4 ) , .A( u2_out15_4 ) );
  XOR2_X1 u2_U489 (.Z( u2_FP_3 ) , .B( u2_L14_3 ) , .A( u2_out15_3 ) );
  XOR2_X1 u2_U49 (.B( u2_L0_26 ) , .Z( u2_N57 ) , .A( u2_out1_26 ) );
  XOR2_X1 u2_U490 (.Z( u2_FP_32 ) , .B( u2_L14_32 ) , .A( u2_out15_32 ) );
  XOR2_X1 u2_U491 (.Z( u2_FP_31 ) , .B( u2_L14_31 ) , .A( u2_out15_31 ) );
  XOR2_X1 u2_U492 (.Z( u2_FP_30 ) , .B( u2_L14_30 ) , .A( u2_out15_30 ) );
  XOR2_X1 u2_U493 (.Z( u2_FP_2 ) , .B( u2_L14_2 ) , .A( u2_out15_2 ) );
  XOR2_X1 u2_U494 (.Z( u2_FP_29 ) , .B( u2_L14_29 ) , .A( u2_out15_29 ) );
  XOR2_X1 u2_U495 (.Z( u2_FP_28 ) , .B( u2_L14_28 ) , .A( u2_out15_28 ) );
  XOR2_X1 u2_U496 (.Z( u2_FP_27 ) , .B( u2_L14_27 ) , .A( u2_out15_27 ) );
  XOR2_X1 u2_U497 (.Z( u2_FP_26 ) , .B( u2_L14_26 ) , .A( u2_out15_26 ) );
  XOR2_X1 u2_U498 (.Z( u2_FP_25 ) , .B( u2_L14_25 ) , .A( u2_out15_25 ) );
  XOR2_X1 u2_U499 (.Z( u2_FP_24 ) , .B( u2_L14_24 ) , .A( u2_out15_24 ) );
  XOR2_X1 u2_U5 (.B( u2_L2_2 ) , .Z( u2_N97 ) , .A( u2_out3_2 ) );
  XOR2_X1 u2_U50 (.B( u2_L0_25 ) , .Z( u2_N56 ) , .A( u2_out1_25 ) );
  XOR2_X1 u2_U500 (.Z( u2_FP_23 ) , .B( u2_L14_23 ) , .A( u2_out15_23 ) );
  XOR2_X1 u2_U501 (.Z( u2_FP_22 ) , .B( u2_L14_22 ) , .A( u2_out15_22 ) );
  XOR2_X1 u2_U502 (.Z( u2_FP_21 ) , .B( u2_L14_21 ) , .A( u2_out15_21 ) );
  XOR2_X1 u2_U503 (.Z( u2_FP_20 ) , .B( u2_L14_20 ) , .A( u2_out15_20 ) );
  XOR2_X1 u2_U504 (.Z( u2_FP_1 ) , .B( u2_L14_1 ) , .A( u2_out15_1 ) );
  XOR2_X1 u2_U505 (.Z( u2_FP_19 ) , .B( u2_L14_19 ) , .A( u2_out15_19 ) );
  XOR2_X1 u2_U506 (.Z( u2_FP_18 ) , .B( u2_L14_18 ) , .A( u2_out15_18 ) );
  XOR2_X1 u2_U507 (.Z( u2_FP_17 ) , .B( u2_L14_17 ) , .A( u2_out15_17 ) );
  XOR2_X1 u2_U508 (.Z( u2_FP_16 ) , .B( u2_L14_16 ) , .A( u2_out15_16 ) );
  XOR2_X1 u2_U509 (.Z( u2_FP_15 ) , .B( u2_L14_15 ) , .A( u2_out15_15 ) );
  XOR2_X1 u2_U51 (.B( u2_L0_24 ) , .Z( u2_N55 ) , .A( u2_out1_24 ) );
  XOR2_X1 u2_U510 (.Z( u2_FP_14 ) , .B( u2_L14_14 ) , .A( u2_out15_14 ) );
  XOR2_X1 u2_U511 (.Z( u2_FP_13 ) , .B( u2_L14_13 ) , .A( u2_out15_13 ) );
  XOR2_X1 u2_U512 (.Z( u2_FP_12 ) , .B( u2_L14_12 ) , .A( u2_out15_12 ) );
  XOR2_X1 u2_U513 (.Z( u2_FP_11 ) , .B( u2_L14_11 ) , .A( u2_out15_11 ) );
  XOR2_X1 u2_U514 (.Z( u2_FP_10 ) , .B( u2_L14_10 ) , .A( u2_out15_10 ) );
  XOR2_X1 u2_U52 (.B( u2_L0_23 ) , .Z( u2_N54 ) , .A( u2_out1_23 ) );
  XOR2_X1 u2_U53 (.B( u2_L0_22 ) , .Z( u2_N53 ) , .A( u2_out1_22 ) );
  XOR2_X1 u2_U54 (.B( u2_L0_21 ) , .Z( u2_N52 ) , .A( u2_out1_21 ) );
  XOR2_X1 u2_U55 (.B( u2_L0_20 ) , .Z( u2_N51 ) , .A( u2_out1_20 ) );
  XOR2_X1 u2_U56 (.B( u2_L0_19 ) , .Z( u2_N50 ) , .A( u2_out1_19 ) );
  XOR2_X1 u2_U57 (.Z( u2_N5 ) , .B( u2_desIn_r_46 ) , .A( u2_out0_6 ) );
  XOR2_X1 u2_U58 (.B( u2_L0_18 ) , .Z( u2_N49 ) , .A( u2_out1_18 ) );
  XOR2_X1 u2_U59 (.B( u2_L0_17 ) , .Z( u2_N48 ) , .A( u2_out1_17 ) );
  XOR2_X1 u2_U6 (.B( u2_L2_1 ) , .Z( u2_N96 ) , .A( u2_out3_1 ) );
  XOR2_X1 u2_U60 (.B( u2_L13_32 ) , .Z( u2_N479 ) , .A( u2_out14_32 ) );
  XOR2_X1 u2_U61 (.B( u2_L13_31 ) , .Z( u2_N478 ) , .A( u2_out14_31 ) );
  XOR2_X1 u2_U62 (.B( u2_L13_30 ) , .Z( u2_N477 ) , .A( u2_out14_30 ) );
  XOR2_X1 u2_U63 (.B( u2_L13_29 ) , .Z( u2_N476 ) , .A( u2_out14_29 ) );
  XOR2_X1 u2_U64 (.B( u2_L13_28 ) , .Z( u2_N475 ) , .A( u2_out14_28 ) );
  XOR2_X1 u2_U65 (.B( u2_L13_27 ) , .Z( u2_N474 ) , .A( u2_out14_27 ) );
  XOR2_X1 u2_U66 (.B( u2_L13_26 ) , .Z( u2_N473 ) , .A( u2_out14_26 ) );
  XOR2_X1 u2_U67 (.B( u2_L13_25 ) , .Z( u2_N472 ) , .A( u2_out14_25 ) );
  XOR2_X1 u2_U68 (.B( u2_L13_24 ) , .Z( u2_N471 ) , .A( u2_out14_24 ) );
  XOR2_X1 u2_U69 (.B( u2_L13_23 ) , .Z( u2_N470 ) , .A( u2_out14_23 ) );
  XOR2_X1 u2_U7 (.B( u2_L1_32 ) , .Z( u2_N95 ) , .A( u2_out2_32 ) );
  XOR2_X1 u2_U70 (.B( u2_L0_16 ) , .Z( u2_N47 ) , .A( u2_out1_16 ) );
  XOR2_X1 u2_U71 (.B( u2_L13_22 ) , .Z( u2_N469 ) , .A( u2_out14_22 ) );
  XOR2_X1 u2_U72 (.B( u2_L13_21 ) , .Z( u2_N468 ) , .A( u2_out14_21 ) );
  XOR2_X1 u2_U73 (.B( u2_L13_20 ) , .Z( u2_N467 ) , .A( u2_out14_20 ) );
  XOR2_X1 u2_U74 (.B( u2_L13_19 ) , .Z( u2_N466 ) , .A( u2_out14_19 ) );
  XOR2_X1 u2_U75 (.B( u2_L13_18 ) , .Z( u2_N465 ) , .A( u2_out14_18 ) );
  XOR2_X1 u2_U76 (.B( u2_L13_17 ) , .Z( u2_N464 ) , .A( u2_out14_17 ) );
  XOR2_X1 u2_U77 (.B( u2_L13_16 ) , .Z( u2_N463 ) , .A( u2_out14_16 ) );
  XOR2_X1 u2_U78 (.B( u2_L13_15 ) , .Z( u2_N462 ) , .A( u2_out14_15 ) );
  XOR2_X1 u2_U79 (.B( u2_L13_14 ) , .Z( u2_N461 ) , .A( u2_out14_14 ) );
  XOR2_X1 u2_U8 (.B( u2_L1_31 ) , .Z( u2_N94 ) , .A( u2_out2_31 ) );
  XOR2_X1 u2_U80 (.B( u2_L13_13 ) , .Z( u2_N460 ) , .A( u2_out14_13 ) );
  XOR2_X1 u2_U81 (.B( u2_L0_15 ) , .Z( u2_N46 ) , .A( u2_out1_15 ) );
  XOR2_X1 u2_U82 (.B( u2_L13_12 ) , .Z( u2_N459 ) , .A( u2_out14_12 ) );
  XOR2_X1 u2_U83 (.B( u2_L13_11 ) , .Z( u2_N458 ) , .A( u2_out14_11 ) );
  XOR2_X1 u2_U84 (.B( u2_L13_10 ) , .Z( u2_N457 ) , .A( u2_out14_10 ) );
  XOR2_X1 u2_U85 (.B( u2_L13_9 ) , .Z( u2_N456 ) , .A( u2_out14_9 ) );
  XOR2_X1 u2_U86 (.B( u2_L13_8 ) , .Z( u2_N455 ) , .A( u2_out14_8 ) );
  XOR2_X1 u2_U87 (.B( u2_L13_7 ) , .Z( u2_N454 ) , .A( u2_out14_7 ) );
  XOR2_X1 u2_U88 (.B( u2_L13_6 ) , .Z( u2_N453 ) , .A( u2_out14_6 ) );
  XOR2_X1 u2_U89 (.B( u2_L13_5 ) , .Z( u2_N452 ) , .A( u2_out14_5 ) );
  XOR2_X1 u2_U9 (.B( u2_L1_30 ) , .Z( u2_N93 ) , .A( u2_out2_30 ) );
  XOR2_X1 u2_U90 (.B( u2_L13_4 ) , .Z( u2_N451 ) , .A( u2_out14_4 ) );
  XOR2_X1 u2_U91 (.B( u2_L13_3 ) , .Z( u2_N450 ) , .A( u2_out14_3 ) );
  XOR2_X1 u2_U92 (.B( u2_L0_14 ) , .Z( u2_N45 ) , .A( u2_out1_14 ) );
  XOR2_X1 u2_U93 (.B( u2_L13_2 ) , .Z( u2_N449 ) , .A( u2_out14_2 ) );
  XOR2_X1 u2_U94 (.B( u2_L13_1 ) , .Z( u2_N448 ) , .A( u2_out14_1 ) );
  XOR2_X1 u2_U95 (.B( u2_L12_32 ) , .Z( u2_N447 ) , .A( u2_out13_32 ) );
  XOR2_X1 u2_U96 (.B( u2_L12_31 ) , .Z( u2_N446 ) , .A( u2_out13_31 ) );
  XOR2_X1 u2_U97 (.B( u2_L12_30 ) , .Z( u2_N445 ) , .A( u2_out13_30 ) );
  XOR2_X1 u2_U98 (.B( u2_L12_29 ) , .Z( u2_N444 ) , .A( u2_out13_29 ) );
  XOR2_X1 u2_U99 (.B( u2_L12_28 ) , .Z( u2_N443 ) , .A( u2_out13_28 ) );
  DFF_X1 u2_desIn_r_reg_0 (.CK( clk ) , .D( stage2_out_0 ) , .Q( u2_desIn_r_0 ) );
  DFF_X1 u2_desIn_r_reg_1 (.CK( clk ) , .D( stage2_out_1 ) , .Q( u2_desIn_r_1 ) );
  DFF_X1 u2_desIn_r_reg_10 (.CK( clk ) , .D( stage2_out_10 ) , .Q( u2_desIn_r_10 ) );
  DFF_X1 u2_desIn_r_reg_11 (.CK( clk ) , .D( stage2_out_11 ) , .Q( u2_desIn_r_11 ) );
  DFF_X1 u2_desIn_r_reg_12 (.CK( clk ) , .D( stage2_out_12 ) , .Q( u2_desIn_r_12 ) );
  DFF_X1 u2_desIn_r_reg_13 (.CK( clk ) , .D( stage2_out_13 ) , .Q( u2_desIn_r_13 ) );
  DFF_X1 u2_desIn_r_reg_14 (.CK( clk ) , .D( stage2_out_14 ) , .Q( u2_desIn_r_14 ) );
  DFF_X1 u2_desIn_r_reg_15 (.CK( clk ) , .D( stage2_out_15 ) , .Q( u2_desIn_r_15 ) );
  DFF_X1 u2_desIn_r_reg_16 (.CK( clk ) , .D( stage2_out_16 ) , .Q( u2_desIn_r_16 ) );
  DFF_X1 u2_desIn_r_reg_17 (.CK( clk ) , .D( stage2_out_17 ) , .Q( u2_desIn_r_17 ) );
  DFF_X1 u2_desIn_r_reg_18 (.CK( clk ) , .D( stage2_out_18 ) , .Q( u2_desIn_r_18 ) );
  DFF_X1 u2_desIn_r_reg_19 (.CK( clk ) , .D( stage2_out_19 ) , .Q( u2_desIn_r_19 ) );
  DFF_X1 u2_desIn_r_reg_2 (.CK( clk ) , .D( stage2_out_2 ) , .Q( u2_desIn_r_2 ) );
  DFF_X1 u2_desIn_r_reg_20 (.CK( clk ) , .D( stage2_out_20 ) , .Q( u2_desIn_r_20 ) );
  DFF_X1 u2_desIn_r_reg_21 (.CK( clk ) , .D( stage2_out_21 ) , .Q( u2_desIn_r_21 ) );
  DFF_X1 u2_desIn_r_reg_22 (.CK( clk ) , .D( stage2_out_22 ) , .Q( u2_desIn_r_22 ) );
  DFF_X1 u2_desIn_r_reg_23 (.CK( clk ) , .D( stage2_out_23 ) , .Q( u2_desIn_r_23 ) );
  DFF_X1 u2_desIn_r_reg_24 (.CK( clk ) , .D( stage2_out_24 ) , .Q( u2_desIn_r_24 ) );
  DFF_X1 u2_desIn_r_reg_25 (.CK( clk ) , .D( stage2_out_25 ) , .Q( u2_desIn_r_25 ) );
  DFF_X1 u2_desIn_r_reg_26 (.CK( clk ) , .D( stage2_out_26 ) , .Q( u2_desIn_r_26 ) );
  DFF_X1 u2_desIn_r_reg_27 (.CK( clk ) , .D( stage2_out_27 ) , .Q( u2_desIn_r_27 ) );
  DFF_X1 u2_desIn_r_reg_28 (.CK( clk ) , .D( stage2_out_28 ) , .Q( u2_desIn_r_28 ) );
  DFF_X1 u2_desIn_r_reg_29 (.CK( clk ) , .D( stage2_out_29 ) , .Q( u2_desIn_r_29 ) );
  DFF_X1 u2_desIn_r_reg_3 (.CK( clk ) , .D( stage2_out_3 ) , .Q( u2_desIn_r_3 ) );
  DFF_X1 u2_desIn_r_reg_30 (.CK( clk ) , .D( stage2_out_30 ) , .Q( u2_desIn_r_30 ) );
  DFF_X1 u2_desIn_r_reg_31 (.CK( clk ) , .D( stage2_out_31 ) , .Q( u2_desIn_r_31 ) );
  DFF_X1 u2_desIn_r_reg_32 (.CK( clk ) , .D( stage2_out_32 ) , .Q( u2_desIn_r_32 ) );
  DFF_X1 u2_desIn_r_reg_33 (.CK( clk ) , .D( stage2_out_33 ) , .Q( u2_desIn_r_33 ) );
  DFF_X1 u2_desIn_r_reg_34 (.CK( clk ) , .D( stage2_out_34 ) , .Q( u2_desIn_r_34 ) );
  DFF_X1 u2_desIn_r_reg_35 (.CK( clk ) , .D( stage2_out_35 ) , .Q( u2_desIn_r_35 ) );
  DFF_X1 u2_desIn_r_reg_36 (.CK( clk ) , .D( stage2_out_36 ) , .Q( u2_desIn_r_36 ) );
  DFF_X1 u2_desIn_r_reg_37 (.CK( clk ) , .D( stage2_out_37 ) , .Q( u2_desIn_r_37 ) );
  DFF_X1 u2_desIn_r_reg_38 (.CK( clk ) , .D( stage2_out_38 ) , .Q( u2_desIn_r_38 ) );
  DFF_X1 u2_desIn_r_reg_39 (.CK( clk ) , .D( stage2_out_39 ) , .Q( u2_desIn_r_39 ) );
  DFF_X1 u2_desIn_r_reg_4 (.CK( clk ) , .D( stage2_out_4 ) , .Q( u2_desIn_r_4 ) );
  DFF_X1 u2_desIn_r_reg_40 (.CK( clk ) , .D( stage2_out_40 ) , .Q( u2_desIn_r_40 ) );
  DFF_X1 u2_desIn_r_reg_41 (.CK( clk ) , .D( stage2_out_41 ) , .Q( u2_desIn_r_41 ) );
  DFF_X1 u2_desIn_r_reg_42 (.CK( clk ) , .D( stage2_out_42 ) , .Q( u2_desIn_r_42 ) );
  DFF_X1 u2_desIn_r_reg_43 (.CK( clk ) , .D( stage2_out_43 ) , .Q( u2_desIn_r_43 ) );
  DFF_X1 u2_desIn_r_reg_44 (.CK( clk ) , .D( stage2_out_44 ) , .Q( u2_desIn_r_44 ) );
  DFF_X1 u2_desIn_r_reg_45 (.CK( clk ) , .D( stage2_out_45 ) , .Q( u2_desIn_r_45 ) );
  DFF_X1 u2_desIn_r_reg_46 (.CK( clk ) , .D( stage2_out_46 ) , .Q( u2_desIn_r_46 ) );
  DFF_X1 u2_desIn_r_reg_47 (.CK( clk ) , .D( stage2_out_47 ) , .Q( u2_desIn_r_47 ) );
  DFF_X1 u2_desIn_r_reg_48 (.CK( clk ) , .D( stage2_out_48 ) , .Q( u2_desIn_r_48 ) );
  DFF_X1 u2_desIn_r_reg_49 (.CK( clk ) , .D( stage2_out_49 ) , .Q( u2_desIn_r_49 ) );
  DFF_X1 u2_desIn_r_reg_5 (.CK( clk ) , .D( stage2_out_5 ) , .Q( u2_desIn_r_5 ) );
  DFF_X1 u2_desIn_r_reg_50 (.CK( clk ) , .D( stage2_out_50 ) , .Q( u2_desIn_r_50 ) );
  DFF_X1 u2_desIn_r_reg_51 (.CK( clk ) , .D( stage2_out_51 ) , .Q( u2_desIn_r_51 ) );
  DFF_X1 u2_desIn_r_reg_52 (.CK( clk ) , .D( stage2_out_52 ) , .Q( u2_desIn_r_52 ) );
  DFF_X1 u2_desIn_r_reg_53 (.CK( clk ) , .D( stage2_out_53 ) , .Q( u2_desIn_r_53 ) );
  DFF_X1 u2_desIn_r_reg_54 (.CK( clk ) , .D( stage2_out_54 ) , .Q( u2_desIn_r_54 ) );
  DFF_X1 u2_desIn_r_reg_55 (.CK( clk ) , .D( stage2_out_55 ) , .Q( u2_desIn_r_55 ) );
  DFF_X1 u2_desIn_r_reg_56 (.CK( clk ) , .D( stage2_out_56 ) , .Q( u2_desIn_r_56 ) );
  DFF_X1 u2_desIn_r_reg_57 (.CK( clk ) , .D( stage2_out_57 ) , .Q( u2_desIn_r_57 ) );
  DFF_X1 u2_desIn_r_reg_58 (.CK( clk ) , .D( stage2_out_58 ) , .Q( u2_desIn_r_58 ) );
  DFF_X1 u2_desIn_r_reg_59 (.CK( clk ) , .D( stage2_out_59 ) , .Q( u2_desIn_r_59 ) );
  DFF_X1 u2_desIn_r_reg_6 (.CK( clk ) , .D( stage2_out_6 ) , .Q( u2_desIn_r_6 ) );
  DFF_X1 u2_desIn_r_reg_60 (.CK( clk ) , .D( stage2_out_60 ) , .Q( u2_desIn_r_60 ) );
  DFF_X1 u2_desIn_r_reg_61 (.CK( clk ) , .D( stage2_out_61 ) , .Q( u2_desIn_r_61 ) );
  DFF_X1 u2_desIn_r_reg_62 (.CK( clk ) , .D( stage2_out_62 ) , .Q( u2_desIn_r_62 ) );
  DFF_X1 u2_desIn_r_reg_63 (.CK( clk ) , .D( stage2_out_63 ) , .Q( u2_desIn_r_63 ) );
  DFF_X1 u2_desIn_r_reg_7 (.CK( clk ) , .D( stage2_out_7 ) , .Q( u2_desIn_r_7 ) );
  DFF_X1 u2_desIn_r_reg_8 (.CK( clk ) , .D( stage2_out_8 ) , .Q( u2_desIn_r_8 ) );
  DFF_X1 u2_desIn_r_reg_9 (.CK( clk ) , .D( stage2_out_9 ) , .Q( u2_desIn_r_9 ) );
  DFF_X1 u2_desOut_reg_0 (.CK( clk ) , .Q( desOut[0] ) , .D( u2_FP_25 ) );
  DFF_X1 u2_desOut_reg_1 (.CK( clk ) , .Q( desOut[1] ) , .D( u2_FP_57 ) );
  DFF_X1 u2_desOut_reg_10 (.CK( clk ) , .Q( desOut[10] ) , .D( u2_FP_18 ) );
  DFF_X1 u2_desOut_reg_11 (.CK( clk ) , .Q( desOut[11] ) , .D( u2_FP_50 ) );
  DFF_X1 u2_desOut_reg_12 (.CK( clk ) , .Q( desOut[12] ) , .D( u2_FP_10 ) );
  DFF_X1 u2_desOut_reg_13 (.CK( clk ) , .Q( desOut[13] ) , .D( u2_FP_42 ) );
  DFF_X1 u2_desOut_reg_14 (.CK( clk ) , .Q( desOut[14] ) , .D( u2_FP_2 ) );
  DFF_X1 u2_desOut_reg_15 (.CK( clk ) , .Q( desOut[15] ) , .D( u2_FP_34 ) );
  DFF_X1 u2_desOut_reg_16 (.CK( clk ) , .Q( desOut[16] ) , .D( u2_FP_27 ) );
  DFF_X1 u2_desOut_reg_17 (.CK( clk ) , .Q( desOut[17] ) , .D( u2_FP_59 ) );
  DFF_X1 u2_desOut_reg_18 (.CK( clk ) , .Q( desOut[18] ) , .D( u2_FP_19 ) );
  DFF_X1 u2_desOut_reg_19 (.CK( clk ) , .Q( desOut[19] ) , .D( u2_FP_51 ) );
  DFF_X1 u2_desOut_reg_2 (.CK( clk ) , .Q( desOut[2] ) , .D( u2_FP_17 ) );
  DFF_X1 u2_desOut_reg_20 (.CK( clk ) , .Q( desOut[20] ) , .D( u2_FP_11 ) );
  DFF_X1 u2_desOut_reg_21 (.CK( clk ) , .Q( desOut[21] ) , .D( u2_FP_43 ) );
  DFF_X1 u2_desOut_reg_22 (.CK( clk ) , .Q( desOut[22] ) , .D( u2_FP_3 ) );
  DFF_X1 u2_desOut_reg_23 (.CK( clk ) , .Q( desOut[23] ) , .D( u2_FP_35 ) );
  DFF_X1 u2_desOut_reg_24 (.CK( clk ) , .Q( desOut[24] ) , .D( u2_FP_28 ) );
  DFF_X1 u2_desOut_reg_25 (.CK( clk ) , .Q( desOut[25] ) , .D( u2_FP_60 ) );
  DFF_X1 u2_desOut_reg_26 (.CK( clk ) , .Q( desOut[26] ) , .D( u2_FP_20 ) );
  DFF_X1 u2_desOut_reg_27 (.CK( clk ) , .Q( desOut[27] ) , .D( u2_FP_52 ) );
  DFF_X1 u2_desOut_reg_28 (.CK( clk ) , .Q( desOut[28] ) , .D( u2_FP_12 ) );
  DFF_X1 u2_desOut_reg_29 (.CK( clk ) , .Q( desOut[29] ) , .D( u2_FP_44 ) );
  DFF_X1 u2_desOut_reg_3 (.CK( clk ) , .Q( desOut[3] ) , .D( u2_FP_49 ) );
  DFF_X1 u2_desOut_reg_30 (.CK( clk ) , .Q( desOut[30] ) , .D( u2_FP_4 ) );
  DFF_X1 u2_desOut_reg_31 (.CK( clk ) , .Q( desOut[31] ) , .D( u2_FP_36 ) );
  DFF_X1 u2_desOut_reg_32 (.CK( clk ) , .Q( desOut[32] ) , .D( u2_FP_29 ) );
  DFF_X1 u2_desOut_reg_33 (.CK( clk ) , .Q( desOut[33] ) , .D( u2_FP_61 ) );
  DFF_X1 u2_desOut_reg_34 (.CK( clk ) , .Q( desOut[34] ) , .D( u2_FP_21 ) );
  DFF_X1 u2_desOut_reg_35 (.CK( clk ) , .Q( desOut[35] ) , .D( u2_FP_53 ) );
  DFF_X1 u2_desOut_reg_36 (.CK( clk ) , .Q( desOut[36] ) , .D( u2_FP_13 ) );
  DFF_X1 u2_desOut_reg_37 (.CK( clk ) , .Q( desOut[37] ) , .D( u2_FP_45 ) );
  DFF_X1 u2_desOut_reg_38 (.CK( clk ) , .Q( desOut[38] ) , .D( u2_FP_5 ) );
  DFF_X1 u2_desOut_reg_39 (.CK( clk ) , .Q( desOut[39] ) , .D( u2_FP_37 ) );
  DFF_X1 u2_desOut_reg_4 (.CK( clk ) , .Q( desOut[4] ) , .D( u2_FP_9 ) );
  DFF_X1 u2_desOut_reg_40 (.CK( clk ) , .Q( desOut[40] ) , .D( u2_FP_30 ) );
  DFF_X1 u2_desOut_reg_41 (.CK( clk ) , .Q( desOut[41] ) , .D( u2_FP_62 ) );
  DFF_X1 u2_desOut_reg_42 (.CK( clk ) , .Q( desOut[42] ) , .D( u2_FP_22 ) );
  DFF_X1 u2_desOut_reg_43 (.CK( clk ) , .Q( desOut[43] ) , .D( u2_FP_54 ) );
  DFF_X1 u2_desOut_reg_44 (.CK( clk ) , .Q( desOut[44] ) , .D( u2_FP_14 ) );
  DFF_X1 u2_desOut_reg_45 (.CK( clk ) , .Q( desOut[45] ) , .D( u2_FP_46 ) );
  DFF_X1 u2_desOut_reg_46 (.CK( clk ) , .Q( desOut[46] ) , .D( u2_FP_6 ) );
  DFF_X1 u2_desOut_reg_47 (.CK( clk ) , .Q( desOut[47] ) , .D( u2_FP_38 ) );
  DFF_X1 u2_desOut_reg_48 (.CK( clk ) , .Q( desOut[48] ) , .D( u2_FP_31 ) );
  DFF_X1 u2_desOut_reg_49 (.CK( clk ) , .Q( desOut[49] ) , .D( u2_FP_63 ) );
  DFF_X1 u2_desOut_reg_5 (.CK( clk ) , .Q( desOut[5] ) , .D( u2_FP_41 ) );
  DFF_X1 u2_desOut_reg_50 (.CK( clk ) , .Q( desOut[50] ) , .D( u2_FP_23 ) );
  DFF_X1 u2_desOut_reg_51 (.CK( clk ) , .Q( desOut[51] ) , .D( u2_FP_55 ) );
  DFF_X1 u2_desOut_reg_52 (.CK( clk ) , .Q( desOut[52] ) , .D( u2_FP_15 ) );
  DFF_X1 u2_desOut_reg_53 (.CK( clk ) , .Q( desOut[53] ) , .D( u2_FP_47 ) );
  DFF_X1 u2_desOut_reg_54 (.CK( clk ) , .Q( desOut[54] ) , .D( u2_FP_7 ) );
  DFF_X1 u2_desOut_reg_55 (.CK( clk ) , .Q( desOut[55] ) , .D( u2_FP_39 ) );
  DFF_X1 u2_desOut_reg_56 (.CK( clk ) , .Q( desOut[56] ) , .D( u2_FP_32 ) );
  DFF_X1 u2_desOut_reg_57 (.CK( clk ) , .Q( desOut[57] ) , .D( u2_FP_64 ) );
  DFF_X1 u2_desOut_reg_58 (.CK( clk ) , .Q( desOut[58] ) , .D( u2_FP_24 ) );
  DFF_X1 u2_desOut_reg_59 (.CK( clk ) , .Q( desOut[59] ) , .D( u2_FP_56 ) );
  DFF_X1 u2_desOut_reg_6 (.CK( clk ) , .Q( desOut[6] ) , .D( u2_FP_1 ) );
  DFF_X1 u2_desOut_reg_60 (.CK( clk ) , .Q( desOut[60] ) , .D( u2_FP_16 ) );
  DFF_X1 u2_desOut_reg_61 (.CK( clk ) , .Q( desOut[61] ) , .D( u2_FP_48 ) );
  DFF_X1 u2_desOut_reg_62 (.CK( clk ) , .Q( desOut[62] ) , .D( u2_FP_8 ) );
  DFF_X1 u2_desOut_reg_63 (.CK( clk ) , .Q( desOut[63] ) , .D( u2_FP_40 ) );
  DFF_X1 u2_desOut_reg_7 (.CK( clk ) , .Q( desOut[7] ) , .D( u2_FP_33 ) );
  DFF_X1 u2_desOut_reg_8 (.CK( clk ) , .Q( desOut[8] ) , .D( u2_FP_26 ) );
  DFF_X1 u2_desOut_reg_9 (.CK( clk ) , .Q( desOut[9] ) , .D( u2_FP_58 ) );
  DFF_X1 u2_key_r_reg_0 (.CK( clk ) , .D( key_c_r_33_0 ) , .Q( u2_key_r_0 ) );
  DFF_X1 u2_key_r_reg_1 (.CK( clk ) , .D( key_c_r_33_1 ) , .Q( u2_key_r_1 ) );
  DFF_X1 u2_key_r_reg_10 (.CK( clk ) , .D( key_c_r_33_10 ) , .Q( u2_key_r_10 ) );
  DFF_X1 u2_key_r_reg_11 (.CK( clk ) , .D( key_c_r_33_11 ) , .Q( u2_key_r_11 ) );
  DFF_X1 u2_key_r_reg_12 (.CK( clk ) , .D( key_c_r_33_12 ) , .Q( u2_key_r_12 ) );
  DFF_X1 u2_key_r_reg_13 (.CK( clk ) , .D( key_c_r_33_13 ) , .Q( u2_key_r_13 ) );
  DFF_X1 u2_key_r_reg_14 (.CK( clk ) , .D( key_c_r_33_14 ) , .Q( u2_key_r_14 ) );
  DFF_X1 u2_key_r_reg_15 (.CK( clk ) , .D( key_c_r_33_15 ) , .Q( u2_key_r_15 ) );
  DFF_X1 u2_key_r_reg_16 (.CK( clk ) , .D( key_c_r_33_16 ) , .Q( u2_key_r_16 ) );
  DFF_X1 u2_key_r_reg_17 (.CK( clk ) , .D( key_c_r_33_17 ) , .Q( u2_key_r_17 ) );
  DFF_X1 u2_key_r_reg_18 (.CK( clk ) , .D( key_c_r_33_18 ) , .Q( u2_key_r_18 ) );
  DFF_X1 u2_key_r_reg_19 (.CK( clk ) , .D( key_c_r_33_19 ) , .Q( u2_key_r_19 ) );
  DFF_X1 u2_key_r_reg_2 (.CK( clk ) , .D( key_c_r_33_2 ) , .Q( u2_key_r_2 ) );
  DFF_X1 u2_key_r_reg_20 (.CK( clk ) , .D( key_c_r_33_20 ) , .Q( u2_key_r_20 ) );
  DFF_X1 u2_key_r_reg_21 (.CK( clk ) , .D( key_c_r_33_21 ) , .Q( u2_key_r_21 ) );
  DFF_X1 u2_key_r_reg_22 (.CK( clk ) , .D( key_c_r_33_22 ) , .Q( u2_key_r_22 ) );
  DFF_X1 u2_key_r_reg_23 (.CK( clk ) , .D( key_c_r_33_23 ) , .Q( u2_key_r_23 ) );
  DFF_X1 u2_key_r_reg_24 (.CK( clk ) , .D( key_c_r_33_24 ) , .Q( u2_key_r_24 ) );
  DFF_X1 u2_key_r_reg_25 (.CK( clk ) , .D( key_c_r_33_25 ) , .Q( u2_key_r_25 ) );
  DFF_X1 u2_key_r_reg_26 (.CK( clk ) , .D( key_c_r_33_26 ) , .Q( u2_key_r_26 ) );
  DFF_X1 u2_key_r_reg_27 (.CK( clk ) , .D( key_c_r_33_27 ) , .Q( u2_key_r_27 ) );
  DFF_X1 u2_key_r_reg_28 (.CK( clk ) , .D( key_c_r_33_28 ) , .Q( u2_key_r_28 ) );
  DFF_X1 u2_key_r_reg_29 (.CK( clk ) , .D( key_c_r_33_29 ) , .Q( u2_key_r_29 ) );
  DFF_X1 u2_key_r_reg_3 (.CK( clk ) , .D( key_c_r_33_3 ) , .Q( u2_key_r_3 ) );
  DFF_X1 u2_key_r_reg_30 (.CK( clk ) , .D( key_c_r_33_30 ) , .Q( u2_key_r_30 ) );
  DFF_X1 u2_key_r_reg_31 (.CK( clk ) , .D( key_c_r_33_31 ) , .Q( u2_key_r_31 ) );
  DFF_X1 u2_key_r_reg_32 (.CK( clk ) , .D( key_c_r_33_32 ) , .Q( u2_key_r_32 ) );
  DFF_X1 u2_key_r_reg_33 (.CK( clk ) , .D( key_c_r_33_33 ) , .Q( u2_key_r_33 ) );
  DFF_X1 u2_key_r_reg_34 (.CK( clk ) , .D( key_c_r_33_34 ) , .Q( u2_key_r_34 ) );
  DFF_X1 u2_key_r_reg_35 (.CK( clk ) , .D( key_c_r_33_35 ) , .Q( u2_key_r_35 ) );
  DFF_X1 u2_key_r_reg_36 (.CK( clk ) , .D( key_c_r_33_36 ) , .Q( u2_key_r_36 ) );
  DFF_X1 u2_key_r_reg_37 (.CK( clk ) , .D( key_c_r_33_37 ) , .Q( u2_key_r_37 ) );
  DFF_X1 u2_key_r_reg_38 (.CK( clk ) , .D( key_c_r_33_38 ) , .Q( u2_key_r_38 ) );
  DFF_X1 u2_key_r_reg_39 (.CK( clk ) , .D( key_c_r_33_39 ) , .Q( u2_key_r_39 ) );
  DFF_X1 u2_key_r_reg_4 (.CK( clk ) , .D( key_c_r_33_4 ) , .Q( u2_key_r_4 ) );
  DFF_X1 u2_key_r_reg_40 (.CK( clk ) , .D( key_c_r_33_40 ) , .Q( u2_key_r_40 ) );
  DFF_X1 u2_key_r_reg_41 (.CK( clk ) , .D( key_c_r_33_41 ) , .Q( u2_key_r_41 ) );
  DFF_X1 u2_key_r_reg_42 (.CK( clk ) , .D( key_c_r_33_42 ) , .Q( u2_key_r_42 ) );
  DFF_X1 u2_key_r_reg_43 (.CK( clk ) , .D( key_c_r_33_43 ) , .Q( u2_key_r_43 ) );
  DFF_X1 u2_key_r_reg_44 (.CK( clk ) , .D( key_c_r_33_44 ) , .Q( u2_key_r_44 ) );
  DFF_X1 u2_key_r_reg_45 (.CK( clk ) , .D( key_c_r_33_45 ) , .Q( u2_key_r_45 ) );
  DFF_X1 u2_key_r_reg_46 (.CK( clk ) , .D( key_c_r_33_46 ) , .Q( u2_key_r_46 ) );
  DFF_X1 u2_key_r_reg_47 (.CK( clk ) , .D( key_c_r_33_47 ) , .Q( u2_key_r_47 ) );
  DFF_X1 u2_key_r_reg_48 (.CK( clk ) , .D( key_c_r_33_48 ) , .Q( u2_key_r_48 ) );
  DFF_X1 u2_key_r_reg_49 (.CK( clk ) , .D( key_c_r_33_49 ) , .Q( u2_key_r_49 ) );
  DFF_X1 u2_key_r_reg_5 (.CK( clk ) , .D( key_c_r_33_5 ) , .Q( u2_key_r_5 ) );
  DFF_X1 u2_key_r_reg_50 (.CK( clk ) , .D( key_c_r_33_50 ) , .Q( u2_key_r_50 ) );
  DFF_X1 u2_key_r_reg_51 (.CK( clk ) , .D( key_c_r_33_51 ) , .Q( u2_key_r_51 ) );
  DFF_X1 u2_key_r_reg_52 (.CK( clk ) , .D( key_c_r_33_52 ) , .Q( u2_key_r_52 ) );
  DFF_X1 u2_key_r_reg_53 (.CK( clk ) , .D( key_c_r_33_53 ) , .Q( u2_key_r_53 ) );
  DFF_X1 u2_key_r_reg_54 (.CK( clk ) , .D( key_c_r_33_54 ) , .Q( u2_key_r_54 ) );
  DFF_X1 u2_key_r_reg_55 (.CK( clk ) , .D( key_c_r_33_55 ) , .Q( u2_key_r_55 ) );
  DFF_X1 u2_key_r_reg_6 (.CK( clk ) , .D( key_c_r_33_6 ) , .Q( u2_key_r_6 ) );
  DFF_X1 u2_key_r_reg_7 (.CK( clk ) , .D( key_c_r_33_7 ) , .Q( u2_key_r_7 ) );
  DFF_X1 u2_key_r_reg_8 (.CK( clk ) , .D( key_c_r_33_8 ) , .Q( u2_key_r_8 ) );
  DFF_X1 u2_key_r_reg_9 (.CK( clk ) , .D( key_c_r_33_9 ) , .Q( u2_key_r_9 ) );
  XOR2_X1 u2_u0_U1 (.B( u2_K1_9 ) , .A( u2_desIn_r_47 ) , .Z( u2_u0_X_9 ) );
  XOR2_X1 u2_u0_U10 (.B( u2_K1_45 ) , .A( u2_desIn_r_41 ) , .Z( u2_u0_X_45 ) );
  XOR2_X1 u2_u0_U15 (.B( u2_K1_40 ) , .A( u2_desIn_r_17 ) , .Z( u2_u0_X_40 ) );
  XOR2_X1 u2_u0_U16 (.B( u2_K1_3 ) , .A( u2_desIn_r_15 ) , .Z( u2_u0_X_3 ) );
  XOR2_X1 u2_u0_U17 (.B( u2_K1_39 ) , .A( u2_desIn_r_9 ) , .Z( u2_u0_X_39 ) );
  XOR2_X1 u2_u0_U19 (.B( u2_K1_37 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_37 ) );
  XOR2_X1 u2_u0_U2 (.B( u2_K1_8 ) , .A( u2_desIn_r_39 ) , .Z( u2_u0_X_8 ) );
  XOR2_X1 u2_u0_U21 (.B( u2_K1_35 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_35 ) );
  XOR2_X1 u2_u0_U22 (.B( u2_K1_34 ) , .A( u2_desIn_r_51 ) , .Z( u2_u0_X_34 ) );
  XOR2_X1 u2_u0_U23 (.B( u2_K1_33 ) , .A( u2_desIn_r_43 ) , .Z( u2_u0_X_33 ) );
  XOR2_X1 u2_u0_U24 (.B( u2_K1_32 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_32 ) );
  XOR2_X1 u2_u0_U26 (.B( u2_K1_30 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_30 ) );
  XOR2_X1 u2_u0_U27 (.B( u2_K1_2 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_2 ) );
  XOR2_X1 u2_u0_U29 (.B( u2_K1_28 ) , .A( u2_desIn_r_19 ) , .Z( u2_u0_X_28 ) );
  XOR2_X1 u2_u0_U3 (.B( u2_K1_7 ) , .A( u2_desIn_r_31 ) , .Z( u2_u0_X_7 ) );
  XOR2_X1 u2_u0_U30 (.B( u2_K1_27 ) , .A( u2_desIn_r_11 ) , .Z( u2_u0_X_27 ) );
  XOR2_X1 u2_u0_U31 (.B( u2_K1_26 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_26 ) );
  XOR2_X1 u2_u0_U32 (.B( u2_K1_25 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_25 ) );
  XOR2_X1 u2_u0_U33 (.B( u2_K1_24 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_24 ) );
  XOR2_X1 u2_u0_U34 (.B( u2_K1_23 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_23 ) );
  XOR2_X1 u2_u0_U35 (.B( u2_K1_22 ) , .A( u2_desIn_r_53 ) , .Z( u2_u0_X_22 ) );
  XOR2_X1 u2_u0_U36 (.B( u2_K1_21 ) , .A( u2_desIn_r_45 ) , .Z( u2_u0_X_21 ) );
  XOR2_X1 u2_u0_U37 (.B( u2_K1_20 ) , .A( u2_desIn_r_37 ) , .Z( u2_u0_X_20 ) );
  XOR2_X1 u2_u0_U38 (.B( u2_K1_1 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_1 ) );
  XOR2_X1 u2_u0_U39 (.B( u2_K1_19 ) , .A( u2_desIn_r_29 ) , .Z( u2_u0_X_19 ) );
  XOR2_X1 u2_u0_U4 (.B( u2_K1_6 ) , .A( u2_desIn_r_39 ) , .Z( u2_u0_X_6 ) );
  XOR2_X1 u2_u0_U40 (.B( u2_K1_18 ) , .A( u2_desIn_r_37 ) , .Z( u2_u0_X_18 ) );
  XOR2_X1 u2_u0_U41 (.B( u2_K1_17 ) , .A( u2_desIn_r_29 ) , .Z( u2_u0_X_17 ) );
  XOR2_X1 u2_u0_U42 (.B( u2_K1_16 ) , .A( u2_desIn_r_21 ) , .Z( u2_u0_X_16 ) );
  XOR2_X1 u2_u0_U43 (.B( u2_K1_15 ) , .A( u2_desIn_r_13 ) , .Z( u2_u0_X_15 ) );
  XOR2_X1 u2_u0_U44 (.B( u2_K1_14 ) , .A( u2_desIn_r_5 ) , .Z( u2_u0_X_14 ) );
  XOR2_X1 u2_u0_U45 (.B( u2_K1_13 ) , .A( u2_desIn_r_63 ) , .Z( u2_u0_X_13 ) );
  XOR2_X1 u2_u0_U46 (.B( u2_K1_12 ) , .A( u2_desIn_r_5 ) , .Z( u2_u0_X_12 ) );
  XOR2_X1 u2_u0_U47 (.B( u2_K1_11 ) , .A( u2_desIn_r_63 ) , .Z( u2_u0_X_11 ) );
  XOR2_X1 u2_u0_U48 (.B( u2_K1_10 ) , .A( u2_desIn_r_55 ) , .Z( u2_u0_X_10 ) );
  XOR2_X1 u2_u0_U5 (.B( u2_K1_5 ) , .A( u2_desIn_r_31 ) , .Z( u2_u0_X_5 ) );
  XOR2_X1 u2_u0_U6 (.B( u2_K1_4 ) , .A( u2_desIn_r_23 ) , .Z( u2_u0_X_4 ) );
  XOR2_X1 u2_u0_U7 (.B( u2_K1_48 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_48 ) );
  XOR2_X1 u2_u0_U9 (.B( u2_K1_46 ) , .A( u2_desIn_r_49 ) , .Z( u2_u0_X_46 ) );
  AND3_X1 u2_u0_u0_U10 (.A2( u2_u0_u0_n112 ) , .ZN( u2_u0_u0_n127 ) , .A3( u2_u0_u0_n130 ) , .A1( u2_u0_u0_n148 ) );
  NAND2_X1 u2_u0_u0_U11 (.ZN( u2_u0_u0_n113 ) , .A1( u2_u0_u0_n139 ) , .A2( u2_u0_u0_n149 ) );
  AND2_X1 u2_u0_u0_U12 (.ZN( u2_u0_u0_n107 ) , .A1( u2_u0_u0_n130 ) , .A2( u2_u0_u0_n140 ) );
  AND2_X1 u2_u0_u0_U13 (.A2( u2_u0_u0_n129 ) , .A1( u2_u0_u0_n130 ) , .ZN( u2_u0_u0_n151 ) );
  AND2_X1 u2_u0_u0_U14 (.A1( u2_u0_u0_n108 ) , .A2( u2_u0_u0_n125 ) , .ZN( u2_u0_u0_n145 ) );
  INV_X1 u2_u0_u0_U15 (.A( u2_u0_u0_n143 ) , .ZN( u2_u0_u0_n173 ) );
  NOR2_X1 u2_u0_u0_U16 (.A2( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n147 ) , .A1( u2_u0_u0_n160 ) );
  OAI22_X1 u2_u0_u0_U17 (.B1( u2_u0_u0_n125 ) , .ZN( u2_u0_u0_n126 ) , .A1( u2_u0_u0_n138 ) , .A2( u2_u0_u0_n146 ) , .B2( u2_u0_u0_n147 ) );
  OAI22_X1 u2_u0_u0_U18 (.B1( u2_u0_u0_n131 ) , .A1( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n147 ) , .A2( u2_u0_u0_n90 ) , .ZN( u2_u0_u0_n91 ) );
  AND3_X1 u2_u0_u0_U19 (.A3( u2_u0_u0_n121 ) , .A2( u2_u0_u0_n125 ) , .A1( u2_u0_u0_n148 ) , .ZN( u2_u0_u0_n90 ) );
  NOR2_X1 u2_u0_u0_U20 (.A1( u2_u0_u0_n163 ) , .A2( u2_u0_u0_n164 ) , .ZN( u2_u0_u0_n95 ) );
  AOI22_X1 u2_u0_u0_U21 (.B2( u2_u0_u0_n109 ) , .A2( u2_u0_u0_n110 ) , .ZN( u2_u0_u0_n111 ) , .B1( u2_u0_u0_n118 ) , .A1( u2_u0_u0_n160 ) );
  NAND2_X1 u2_u0_u0_U22 (.A1( u2_u0_u0_n100 ) , .A2( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n125 ) );
  NAND2_X1 u2_u0_u0_U23 (.A1( u2_u0_u0_n101 ) , .A2( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n150 ) );
  INV_X1 u2_u0_u0_U24 (.A( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n161 ) );
  INV_X1 u2_u0_u0_U25 (.A( u2_u0_u0_n118 ) , .ZN( u2_u0_u0_n158 ) );
  AOI21_X1 u2_u0_u0_U26 (.B1( u2_u0_u0_n127 ) , .B2( u2_u0_u0_n129 ) , .A( u2_u0_u0_n138 ) , .ZN( u2_u0_u0_n96 ) );
  AOI21_X1 u2_u0_u0_U27 (.ZN( u2_u0_u0_n104 ) , .B1( u2_u0_u0_n107 ) , .B2( u2_u0_u0_n141 ) , .A( u2_u0_u0_n144 ) );
  NAND2_X1 u2_u0_u0_U28 (.A2( u2_u0_u0_n100 ) , .A1( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n139 ) );
  NAND2_X1 u2_u0_u0_U29 (.A2( u2_u0_u0_n100 ) , .ZN( u2_u0_u0_n131 ) , .A1( u2_u0_u0_n92 ) );
  INV_X1 u2_u0_u0_U3 (.A( u2_u0_u0_n113 ) , .ZN( u2_u0_u0_n166 ) );
  NAND2_X1 u2_u0_u0_U30 (.A2( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n114 ) , .A1( u2_u0_u0_n92 ) );
  NOR2_X1 u2_u0_u0_U31 (.A1( u2_u0_u0_n120 ) , .ZN( u2_u0_u0_n143 ) , .A2( u2_u0_u0_n167 ) );
  OAI221_X1 u2_u0_u0_U32 (.C1( u2_u0_u0_n112 ) , .ZN( u2_u0_u0_n120 ) , .B1( u2_u0_u0_n138 ) , .B2( u2_u0_u0_n141 ) , .C2( u2_u0_u0_n147 ) , .A( u2_u0_u0_n172 ) );
  AOI211_X1 u2_u0_u0_U33 (.B( u2_u0_u0_n115 ) , .A( u2_u0_u0_n116 ) , .C2( u2_u0_u0_n117 ) , .C1( u2_u0_u0_n118 ) , .ZN( u2_u0_u0_n119 ) );
  INV_X1 u2_u0_u0_U34 (.A( u2_u0_u0_n138 ) , .ZN( u2_u0_u0_n160 ) );
  NAND2_X1 u2_u0_u0_U35 (.A2( u2_u0_u0_n102 ) , .A1( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n149 ) );
  NAND2_X1 u2_u0_u0_U36 (.A2( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n121 ) , .A1( u2_u0_u0_n93 ) );
  NAND2_X1 u2_u0_u0_U37 (.ZN( u2_u0_u0_n112 ) , .A2( u2_u0_u0_n92 ) , .A1( u2_u0_u0_n93 ) );
  INV_X1 u2_u0_u0_U38 (.ZN( u2_u0_u0_n172 ) , .A( u2_u0_u0_n88 ) );
  OAI222_X1 u2_u0_u0_U39 (.C1( u2_u0_u0_n108 ) , .A1( u2_u0_u0_n125 ) , .B2( u2_u0_u0_n128 ) , .B1( u2_u0_u0_n144 ) , .A2( u2_u0_u0_n158 ) , .C2( u2_u0_u0_n161 ) , .ZN( u2_u0_u0_n88 ) );
  AOI21_X1 u2_u0_u0_U4 (.B1( u2_u0_u0_n114 ) , .ZN( u2_u0_u0_n115 ) , .B2( u2_u0_u0_n129 ) , .A( u2_u0_u0_n161 ) );
  AOI21_X1 u2_u0_u0_U40 (.B1( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n132 ) , .A( u2_u0_u0_n165 ) , .B2( u2_u0_u0_n93 ) );
  OR3_X1 u2_u0_u0_U41 (.A3( u2_u0_u0_n152 ) , .A2( u2_u0_u0_n153 ) , .A1( u2_u0_u0_n154 ) , .ZN( u2_u0_u0_n155 ) );
  AOI21_X1 u2_u0_u0_U42 (.B2( u2_u0_u0_n150 ) , .B1( u2_u0_u0_n151 ) , .ZN( u2_u0_u0_n152 ) , .A( u2_u0_u0_n158 ) );
  AOI21_X1 u2_u0_u0_U43 (.A( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n145 ) , .B1( u2_u0_u0_n146 ) , .ZN( u2_u0_u0_n154 ) );
  AOI21_X1 u2_u0_u0_U44 (.A( u2_u0_u0_n147 ) , .B2( u2_u0_u0_n148 ) , .B1( u2_u0_u0_n149 ) , .ZN( u2_u0_u0_n153 ) );
  INV_X1 u2_u0_u0_U45 (.ZN( u2_u0_u0_n171 ) , .A( u2_u0_u0_n99 ) );
  OAI211_X1 u2_u0_u0_U46 (.C2( u2_u0_u0_n140 ) , .C1( u2_u0_u0_n161 ) , .A( u2_u0_u0_n169 ) , .B( u2_u0_u0_n98 ) , .ZN( u2_u0_u0_n99 ) );
  INV_X1 u2_u0_u0_U47 (.ZN( u2_u0_u0_n169 ) , .A( u2_u0_u0_n91 ) );
  AOI211_X1 u2_u0_u0_U48 (.C1( u2_u0_u0_n118 ) , .A( u2_u0_u0_n123 ) , .B( u2_u0_u0_n96 ) , .C2( u2_u0_u0_n97 ) , .ZN( u2_u0_u0_n98 ) );
  NOR2_X1 u2_u0_u0_U49 (.A2( u2_u0_X_4 ) , .A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n118 ) );
  NOR2_X1 u2_u0_u0_U5 (.A1( u2_u0_u0_n108 ) , .ZN( u2_u0_u0_n123 ) , .A2( u2_u0_u0_n158 ) );
  NOR2_X1 u2_u0_u0_U50 (.A2( u2_u0_X_2 ) , .ZN( u2_u0_u0_n103 ) , .A1( u2_u0_u0_n164 ) );
  NAND2_X1 u2_u0_u0_U51 (.A2( u2_u0_X_4 ) , .A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n144 ) );
  NOR2_X1 u2_u0_u0_U52 (.A2( u2_u0_X_5 ) , .ZN( u2_u0_u0_n136 ) , .A1( u2_u0_u0_n159 ) );
  NAND2_X1 u2_u0_u0_U53 (.A1( u2_u0_X_5 ) , .ZN( u2_u0_u0_n138 ) , .A2( u2_u0_u0_n159 ) );
  AND2_X1 u2_u0_u0_U54 (.A2( u2_u0_X_3 ) , .A1( u2_u0_X_6 ) , .ZN( u2_u0_u0_n102 ) );
  INV_X1 u2_u0_u0_U55 (.A( u2_u0_X_4 ) , .ZN( u2_u0_u0_n159 ) );
  INV_X1 u2_u0_u0_U56 (.A( u2_u0_X_2 ) , .ZN( u2_u0_u0_n163 ) );
  INV_X1 u2_u0_u0_U57 (.A( u2_u0_X_3 ) , .ZN( u2_u0_u0_n162 ) );
  INV_X1 u2_u0_u0_U58 (.A( u2_u0_u0_n126 ) , .ZN( u2_u0_u0_n168 ) );
  AOI211_X1 u2_u0_u0_U59 (.B( u2_u0_u0_n133 ) , .A( u2_u0_u0_n134 ) , .C2( u2_u0_u0_n135 ) , .C1( u2_u0_u0_n136 ) , .ZN( u2_u0_u0_n137 ) );
  AOI21_X1 u2_u0_u0_U6 (.B2( u2_u0_u0_n131 ) , .ZN( u2_u0_u0_n134 ) , .B1( u2_u0_u0_n151 ) , .A( u2_u0_u0_n158 ) );
  OR4_X1 u2_u0_u0_U60 (.ZN( u2_out0_17 ) , .A4( u2_u0_u0_n122 ) , .A2( u2_u0_u0_n123 ) , .A1( u2_u0_u0_n124 ) , .A3( u2_u0_u0_n170 ) );
  AOI21_X1 u2_u0_u0_U61 (.B2( u2_u0_u0_n107 ) , .ZN( u2_u0_u0_n124 ) , .B1( u2_u0_u0_n128 ) , .A( u2_u0_u0_n161 ) );
  INV_X1 u2_u0_u0_U62 (.A( u2_u0_u0_n111 ) , .ZN( u2_u0_u0_n170 ) );
  OR4_X1 u2_u0_u0_U63 (.ZN( u2_out0_31 ) , .A4( u2_u0_u0_n155 ) , .A2( u2_u0_u0_n156 ) , .A1( u2_u0_u0_n157 ) , .A3( u2_u0_u0_n173 ) );
  AOI21_X1 u2_u0_u0_U64 (.A( u2_u0_u0_n138 ) , .B2( u2_u0_u0_n139 ) , .B1( u2_u0_u0_n140 ) , .ZN( u2_u0_u0_n157 ) );
  INV_X1 u2_u0_u0_U65 (.ZN( u2_u0_u0_n174 ) , .A( u2_u0_u0_n89 ) );
  AOI211_X1 u2_u0_u0_U66 (.B( u2_u0_u0_n104 ) , .A( u2_u0_u0_n105 ) , .ZN( u2_u0_u0_n106 ) , .C2( u2_u0_u0_n113 ) , .C1( u2_u0_u0_n160 ) );
  AOI21_X1 u2_u0_u0_U67 (.B2( u2_u0_u0_n141 ) , .B1( u2_u0_u0_n142 ) , .ZN( u2_u0_u0_n156 ) , .A( u2_u0_u0_n161 ) );
  AOI21_X1 u2_u0_u0_U68 (.ZN( u2_u0_u0_n116 ) , .B2( u2_u0_u0_n142 ) , .A( u2_u0_u0_n144 ) , .B1( u2_u0_u0_n166 ) );
  NAND2_X1 u2_u0_u0_U69 (.ZN( u2_u0_u0_n148 ) , .A1( u2_u0_u0_n93 ) , .A2( u2_u0_u0_n95 ) );
  OAI21_X1 u2_u0_u0_U7 (.B1( u2_u0_u0_n150 ) , .B2( u2_u0_u0_n158 ) , .A( u2_u0_u0_n172 ) , .ZN( u2_u0_u0_n89 ) );
  NAND2_X1 u2_u0_u0_U70 (.A1( u2_u0_u0_n100 ) , .ZN( u2_u0_u0_n129 ) , .A2( u2_u0_u0_n95 ) );
  NAND2_X1 u2_u0_u0_U71 (.A1( u2_u0_u0_n102 ) , .ZN( u2_u0_u0_n128 ) , .A2( u2_u0_u0_n95 ) );
  INV_X1 u2_u0_u0_U72 (.A( u2_u0_u0_n142 ) , .ZN( u2_u0_u0_n165 ) );
  NOR2_X1 u2_u0_u0_U73 (.A2( u2_u0_X_1 ) , .A1( u2_u0_X_2 ) , .ZN( u2_u0_u0_n92 ) );
  NOR2_X1 u2_u0_u0_U74 (.A2( u2_u0_X_1 ) , .ZN( u2_u0_u0_n101 ) , .A1( u2_u0_u0_n163 ) );
  INV_X1 u2_u0_u0_U75 (.A( u2_u0_X_1 ) , .ZN( u2_u0_u0_n164 ) );
  AND2_X1 u2_u0_u0_U76 (.A1( u2_u0_X_6 ) , .A2( u2_u0_u0_n162 ) , .ZN( u2_u0_u0_n93 ) );
  NOR2_X1 u2_u0_u0_U77 (.A2( u2_u0_X_3 ) , .A1( u2_u0_X_6 ) , .ZN( u2_u0_u0_n94 ) );
  NOR2_X1 u2_u0_u0_U78 (.A2( u2_u0_X_6 ) , .ZN( u2_u0_u0_n100 ) , .A1( u2_u0_u0_n162 ) );
  OAI221_X1 u2_u0_u0_U79 (.C1( u2_u0_u0_n121 ) , .ZN( u2_u0_u0_n122 ) , .B2( u2_u0_u0_n127 ) , .A( u2_u0_u0_n143 ) , .B1( u2_u0_u0_n144 ) , .C2( u2_u0_u0_n147 ) );
  AND2_X1 u2_u0_u0_U8 (.A1( u2_u0_u0_n114 ) , .A2( u2_u0_u0_n121 ) , .ZN( u2_u0_u0_n146 ) );
  AOI21_X1 u2_u0_u0_U80 (.B1( u2_u0_u0_n132 ) , .ZN( u2_u0_u0_n133 ) , .A( u2_u0_u0_n144 ) , .B2( u2_u0_u0_n166 ) );
  OAI22_X1 u2_u0_u0_U81 (.ZN( u2_u0_u0_n105 ) , .A2( u2_u0_u0_n132 ) , .B1( u2_u0_u0_n146 ) , .A1( u2_u0_u0_n147 ) , .B2( u2_u0_u0_n161 ) );
  NAND2_X1 u2_u0_u0_U82 (.ZN( u2_u0_u0_n110 ) , .A2( u2_u0_u0_n132 ) , .A1( u2_u0_u0_n145 ) );
  INV_X1 u2_u0_u0_U83 (.A( u2_u0_u0_n119 ) , .ZN( u2_u0_u0_n167 ) );
  NAND2_X1 u2_u0_u0_U84 (.A2( u2_u0_u0_n103 ) , .ZN( u2_u0_u0_n140 ) , .A1( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U85 (.A1( u2_u0_u0_n101 ) , .ZN( u2_u0_u0_n130 ) , .A2( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U86 (.ZN( u2_u0_u0_n108 ) , .A1( u2_u0_u0_n92 ) , .A2( u2_u0_u0_n94 ) );
  NAND2_X1 u2_u0_u0_U87 (.ZN( u2_u0_u0_n142 ) , .A1( u2_u0_u0_n94 ) , .A2( u2_u0_u0_n95 ) );
  NAND3_X1 u2_u0_u0_U88 (.ZN( u2_out0_23 ) , .A3( u2_u0_u0_n137 ) , .A1( u2_u0_u0_n168 ) , .A2( u2_u0_u0_n171 ) );
  NAND3_X1 u2_u0_u0_U89 (.A3( u2_u0_u0_n127 ) , .A2( u2_u0_u0_n128 ) , .ZN( u2_u0_u0_n135 ) , .A1( u2_u0_u0_n150 ) );
  AND2_X1 u2_u0_u0_U9 (.A1( u2_u0_u0_n131 ) , .ZN( u2_u0_u0_n141 ) , .A2( u2_u0_u0_n150 ) );
  NAND3_X1 u2_u0_u0_U90 (.ZN( u2_u0_u0_n117 ) , .A3( u2_u0_u0_n132 ) , .A2( u2_u0_u0_n139 ) , .A1( u2_u0_u0_n148 ) );
  NAND3_X1 u2_u0_u0_U91 (.ZN( u2_u0_u0_n109 ) , .A2( u2_u0_u0_n114 ) , .A3( u2_u0_u0_n140 ) , .A1( u2_u0_u0_n149 ) );
  NAND3_X1 u2_u0_u0_U92 (.ZN( u2_out0_9 ) , .A3( u2_u0_u0_n106 ) , .A2( u2_u0_u0_n171 ) , .A1( u2_u0_u0_n174 ) );
  NAND3_X1 u2_u0_u0_U93 (.A2( u2_u0_u0_n128 ) , .A1( u2_u0_u0_n132 ) , .A3( u2_u0_u0_n146 ) , .ZN( u2_u0_u0_n97 ) );
  OAI22_X1 u2_u0_u2_U10 (.B1( u2_u0_u2_n151 ) , .A2( u2_u0_u2_n152 ) , .A1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n160 ) , .B2( u2_u0_u2_n168 ) );
  NAND3_X1 u2_u0_u2_U100 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n98 ) );
  NOR3_X1 u2_u0_u2_U11 (.A1( u2_u0_u2_n150 ) , .ZN( u2_u0_u2_n151 ) , .A3( u2_u0_u2_n175 ) , .A2( u2_u0_u2_n188 ) );
  AOI21_X1 u2_u0_u2_U12 (.B2( u2_u0_u2_n123 ) , .ZN( u2_u0_u2_n125 ) , .A( u2_u0_u2_n171 ) , .B1( u2_u0_u2_n184 ) );
  INV_X1 u2_u0_u2_U13 (.A( u2_u0_u2_n150 ) , .ZN( u2_u0_u2_n184 ) );
  AOI21_X1 u2_u0_u2_U14 (.ZN( u2_u0_u2_n144 ) , .B2( u2_u0_u2_n155 ) , .A( u2_u0_u2_n172 ) , .B1( u2_u0_u2_n185 ) );
  AOI21_X1 u2_u0_u2_U15 (.B2( u2_u0_u2_n143 ) , .ZN( u2_u0_u2_n145 ) , .B1( u2_u0_u2_n152 ) , .A( u2_u0_u2_n171 ) );
  INV_X1 u2_u0_u2_U16 (.A( u2_u0_u2_n156 ) , .ZN( u2_u0_u2_n171 ) );
  INV_X1 u2_u0_u2_U17 (.A( u2_u0_u2_n120 ) , .ZN( u2_u0_u2_n188 ) );
  NAND2_X1 u2_u0_u2_U18 (.A2( u2_u0_u2_n122 ) , .ZN( u2_u0_u2_n150 ) , .A1( u2_u0_u2_n152 ) );
  INV_X1 u2_u0_u2_U19 (.A( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n170 ) );
  INV_X1 u2_u0_u2_U20 (.A( u2_u0_u2_n137 ) , .ZN( u2_u0_u2_n173 ) );
  NAND2_X1 u2_u0_u2_U21 (.A1( u2_u0_u2_n132 ) , .A2( u2_u0_u2_n139 ) , .ZN( u2_u0_u2_n157 ) );
  INV_X1 u2_u0_u2_U22 (.A( u2_u0_u2_n113 ) , .ZN( u2_u0_u2_n178 ) );
  INV_X1 u2_u0_u2_U23 (.A( u2_u0_u2_n139 ) , .ZN( u2_u0_u2_n175 ) );
  INV_X1 u2_u0_u2_U24 (.A( u2_u0_u2_n155 ) , .ZN( u2_u0_u2_n181 ) );
  INV_X1 u2_u0_u2_U25 (.A( u2_u0_u2_n119 ) , .ZN( u2_u0_u2_n177 ) );
  INV_X1 u2_u0_u2_U26 (.A( u2_u0_u2_n116 ) , .ZN( u2_u0_u2_n180 ) );
  INV_X1 u2_u0_u2_U27 (.A( u2_u0_u2_n131 ) , .ZN( u2_u0_u2_n179 ) );
  INV_X1 u2_u0_u2_U28 (.A( u2_u0_u2_n154 ) , .ZN( u2_u0_u2_n176 ) );
  NAND2_X1 u2_u0_u2_U29 (.A2( u2_u0_u2_n116 ) , .A1( u2_u0_u2_n117 ) , .ZN( u2_u0_u2_n118 ) );
  NOR2_X1 u2_u0_u2_U3 (.ZN( u2_u0_u2_n121 ) , .A2( u2_u0_u2_n177 ) , .A1( u2_u0_u2_n180 ) );
  INV_X1 u2_u0_u2_U30 (.A( u2_u0_u2_n132 ) , .ZN( u2_u0_u2_n182 ) );
  INV_X1 u2_u0_u2_U31 (.A( u2_u0_u2_n158 ) , .ZN( u2_u0_u2_n183 ) );
  OAI21_X1 u2_u0_u2_U32 (.A( u2_u0_u2_n156 ) , .B1( u2_u0_u2_n157 ) , .ZN( u2_u0_u2_n158 ) , .B2( u2_u0_u2_n179 ) );
  NOR2_X1 u2_u0_u2_U33 (.ZN( u2_u0_u2_n156 ) , .A1( u2_u0_u2_n166 ) , .A2( u2_u0_u2_n169 ) );
  NOR2_X1 u2_u0_u2_U34 (.A2( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n137 ) , .A1( u2_u0_u2_n140 ) );
  NOR2_X1 u2_u0_u2_U35 (.A2( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n153 ) , .A1( u2_u0_u2_n156 ) );
  AOI211_X1 u2_u0_u2_U36 (.ZN( u2_u0_u2_n130 ) , .C1( u2_u0_u2_n138 ) , .C2( u2_u0_u2_n179 ) , .B( u2_u0_u2_n96 ) , .A( u2_u0_u2_n97 ) );
  OAI22_X1 u2_u0_u2_U37 (.B1( u2_u0_u2_n133 ) , .A2( u2_u0_u2_n137 ) , .A1( u2_u0_u2_n152 ) , .B2( u2_u0_u2_n168 ) , .ZN( u2_u0_u2_n97 ) );
  OAI221_X1 u2_u0_u2_U38 (.B1( u2_u0_u2_n113 ) , .C1( u2_u0_u2_n132 ) , .A( u2_u0_u2_n149 ) , .B2( u2_u0_u2_n171 ) , .C2( u2_u0_u2_n172 ) , .ZN( u2_u0_u2_n96 ) );
  OAI221_X1 u2_u0_u2_U39 (.A( u2_u0_u2_n115 ) , .C2( u2_u0_u2_n123 ) , .B2( u2_u0_u2_n143 ) , .B1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n163 ) , .C1( u2_u0_u2_n168 ) );
  INV_X1 u2_u0_u2_U4 (.A( u2_u0_u2_n134 ) , .ZN( u2_u0_u2_n185 ) );
  OAI21_X1 u2_u0_u2_U40 (.A( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n115 ) , .B1( u2_u0_u2_n176 ) , .B2( u2_u0_u2_n178 ) );
  OAI221_X1 u2_u0_u2_U41 (.A( u2_u0_u2_n135 ) , .B2( u2_u0_u2_n136 ) , .B1( u2_u0_u2_n137 ) , .ZN( u2_u0_u2_n162 ) , .C2( u2_u0_u2_n167 ) , .C1( u2_u0_u2_n185 ) );
  AND3_X1 u2_u0_u2_U42 (.A3( u2_u0_u2_n131 ) , .A2( u2_u0_u2_n132 ) , .A1( u2_u0_u2_n133 ) , .ZN( u2_u0_u2_n136 ) );
  AOI22_X1 u2_u0_u2_U43 (.ZN( u2_u0_u2_n135 ) , .B1( u2_u0_u2_n140 ) , .A1( u2_u0_u2_n156 ) , .B2( u2_u0_u2_n180 ) , .A2( u2_u0_u2_n188 ) );
  AOI21_X1 u2_u0_u2_U44 (.ZN( u2_u0_u2_n149 ) , .B1( u2_u0_u2_n173 ) , .B2( u2_u0_u2_n188 ) , .A( u2_u0_u2_n95 ) );
  AND3_X1 u2_u0_u2_U45 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n156 ) , .ZN( u2_u0_u2_n95 ) );
  OAI21_X1 u2_u0_u2_U46 (.A( u2_u0_u2_n141 ) , .B2( u2_u0_u2_n142 ) , .ZN( u2_u0_u2_n146 ) , .B1( u2_u0_u2_n153 ) );
  OAI21_X1 u2_u0_u2_U47 (.A( u2_u0_u2_n140 ) , .ZN( u2_u0_u2_n141 ) , .B1( u2_u0_u2_n176 ) , .B2( u2_u0_u2_n177 ) );
  NOR3_X1 u2_u0_u2_U48 (.ZN( u2_u0_u2_n142 ) , .A3( u2_u0_u2_n175 ) , .A2( u2_u0_u2_n178 ) , .A1( u2_u0_u2_n181 ) );
  OAI21_X1 u2_u0_u2_U49 (.A( u2_u0_u2_n101 ) , .B2( u2_u0_u2_n121 ) , .B1( u2_u0_u2_n153 ) , .ZN( u2_u0_u2_n164 ) );
  NOR4_X1 u2_u0_u2_U5 (.A4( u2_u0_u2_n124 ) , .A3( u2_u0_u2_n125 ) , .A2( u2_u0_u2_n126 ) , .A1( u2_u0_u2_n127 ) , .ZN( u2_u0_u2_n128 ) );
  NAND2_X1 u2_u0_u2_U50 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n155 ) );
  NAND2_X1 u2_u0_u2_U51 (.A2( u2_u0_u2_n105 ) , .A1( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n143 ) );
  NAND2_X1 u2_u0_u2_U52 (.A1( u2_u0_u2_n104 ) , .A2( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n152 ) );
  NAND2_X1 u2_u0_u2_U53 (.A1( u2_u0_u2_n100 ) , .A2( u2_u0_u2_n105 ) , .ZN( u2_u0_u2_n132 ) );
  INV_X1 u2_u0_u2_U54 (.A( u2_u0_u2_n140 ) , .ZN( u2_u0_u2_n168 ) );
  INV_X1 u2_u0_u2_U55 (.A( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n167 ) );
  NAND2_X1 u2_u0_u2_U56 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n113 ) );
  NAND2_X1 u2_u0_u2_U57 (.A1( u2_u0_u2_n106 ) , .A2( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n131 ) );
  NAND2_X1 u2_u0_u2_U58 (.A1( u2_u0_u2_n103 ) , .A2( u2_u0_u2_n107 ) , .ZN( u2_u0_u2_n139 ) );
  NAND2_X1 u2_u0_u2_U59 (.A1( u2_u0_u2_n103 ) , .A2( u2_u0_u2_n105 ) , .ZN( u2_u0_u2_n133 ) );
  AOI21_X1 u2_u0_u2_U6 (.B2( u2_u0_u2_n119 ) , .ZN( u2_u0_u2_n127 ) , .A( u2_u0_u2_n137 ) , .B1( u2_u0_u2_n155 ) );
  NAND2_X1 u2_u0_u2_U60 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n103 ) , .ZN( u2_u0_u2_n154 ) );
  NAND2_X1 u2_u0_u2_U61 (.A2( u2_u0_u2_n103 ) , .A1( u2_u0_u2_n104 ) , .ZN( u2_u0_u2_n119 ) );
  NAND2_X1 u2_u0_u2_U62 (.A2( u2_u0_u2_n107 ) , .A1( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n123 ) );
  NAND2_X1 u2_u0_u2_U63 (.A1( u2_u0_u2_n104 ) , .A2( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n122 ) );
  INV_X1 u2_u0_u2_U64 (.A( u2_u0_u2_n114 ) , .ZN( u2_u0_u2_n172 ) );
  NAND2_X1 u2_u0_u2_U65 (.A2( u2_u0_u2_n100 ) , .A1( u2_u0_u2_n102 ) , .ZN( u2_u0_u2_n116 ) );
  NAND2_X1 u2_u0_u2_U66 (.A1( u2_u0_u2_n102 ) , .A2( u2_u0_u2_n108 ) , .ZN( u2_u0_u2_n120 ) );
  NAND2_X1 u2_u0_u2_U67 (.A2( u2_u0_u2_n105 ) , .A1( u2_u0_u2_n106 ) , .ZN( u2_u0_u2_n117 ) );
  INV_X1 u2_u0_u2_U68 (.ZN( u2_u0_u2_n187 ) , .A( u2_u0_u2_n99 ) );
  OAI21_X1 u2_u0_u2_U69 (.B1( u2_u0_u2_n137 ) , .B2( u2_u0_u2_n143 ) , .A( u2_u0_u2_n98 ) , .ZN( u2_u0_u2_n99 ) );
  AOI21_X1 u2_u0_u2_U7 (.ZN( u2_u0_u2_n124 ) , .B1( u2_u0_u2_n131 ) , .B2( u2_u0_u2_n143 ) , .A( u2_u0_u2_n172 ) );
  NOR2_X1 u2_u0_u2_U70 (.A2( u2_u0_X_16 ) , .ZN( u2_u0_u2_n140 ) , .A1( u2_u0_u2_n166 ) );
  NOR2_X1 u2_u0_u2_U71 (.A2( u2_u0_X_13 ) , .A1( u2_u0_X_14 ) , .ZN( u2_u0_u2_n100 ) );
  NOR2_X1 u2_u0_u2_U72 (.A2( u2_u0_X_16 ) , .A1( u2_u0_X_17 ) , .ZN( u2_u0_u2_n138 ) );
  NOR2_X1 u2_u0_u2_U73 (.A2( u2_u0_X_15 ) , .A1( u2_u0_X_18 ) , .ZN( u2_u0_u2_n104 ) );
  NOR2_X1 u2_u0_u2_U74 (.A2( u2_u0_X_14 ) , .ZN( u2_u0_u2_n103 ) , .A1( u2_u0_u2_n174 ) );
  NOR2_X1 u2_u0_u2_U75 (.A2( u2_u0_X_15 ) , .ZN( u2_u0_u2_n102 ) , .A1( u2_u0_u2_n165 ) );
  NOR2_X1 u2_u0_u2_U76 (.A2( u2_u0_X_17 ) , .ZN( u2_u0_u2_n114 ) , .A1( u2_u0_u2_n169 ) );
  AND2_X1 u2_u0_u2_U77 (.A1( u2_u0_X_15 ) , .ZN( u2_u0_u2_n105 ) , .A2( u2_u0_u2_n165 ) );
  AND2_X1 u2_u0_u2_U78 (.A2( u2_u0_X_15 ) , .A1( u2_u0_X_18 ) , .ZN( u2_u0_u2_n107 ) );
  AND2_X1 u2_u0_u2_U79 (.A1( u2_u0_X_14 ) , .ZN( u2_u0_u2_n106 ) , .A2( u2_u0_u2_n174 ) );
  AOI21_X1 u2_u0_u2_U8 (.B2( u2_u0_u2_n120 ) , .B1( u2_u0_u2_n121 ) , .ZN( u2_u0_u2_n126 ) , .A( u2_u0_u2_n167 ) );
  AND2_X1 u2_u0_u2_U80 (.A1( u2_u0_X_13 ) , .A2( u2_u0_X_14 ) , .ZN( u2_u0_u2_n108 ) );
  INV_X1 u2_u0_u2_U81 (.A( u2_u0_X_16 ) , .ZN( u2_u0_u2_n169 ) );
  INV_X1 u2_u0_u2_U82 (.A( u2_u0_X_17 ) , .ZN( u2_u0_u2_n166 ) );
  INV_X1 u2_u0_u2_U83 (.A( u2_u0_X_13 ) , .ZN( u2_u0_u2_n174 ) );
  INV_X1 u2_u0_u2_U84 (.A( u2_u0_X_18 ) , .ZN( u2_u0_u2_n165 ) );
  NAND4_X1 u2_u0_u2_U85 (.ZN( u2_out0_30 ) , .A4( u2_u0_u2_n147 ) , .A3( u2_u0_u2_n148 ) , .A2( u2_u0_u2_n149 ) , .A1( u2_u0_u2_n187 ) );
  NOR3_X1 u2_u0_u2_U86 (.A3( u2_u0_u2_n144 ) , .A2( u2_u0_u2_n145 ) , .A1( u2_u0_u2_n146 ) , .ZN( u2_u0_u2_n147 ) );
  AOI21_X1 u2_u0_u2_U87 (.B2( u2_u0_u2_n138 ) , .ZN( u2_u0_u2_n148 ) , .A( u2_u0_u2_n162 ) , .B1( u2_u0_u2_n182 ) );
  NAND4_X1 u2_u0_u2_U88 (.ZN( u2_out0_24 ) , .A4( u2_u0_u2_n111 ) , .A3( u2_u0_u2_n112 ) , .A1( u2_u0_u2_n130 ) , .A2( u2_u0_u2_n187 ) );
  AOI221_X1 u2_u0_u2_U89 (.A( u2_u0_u2_n109 ) , .B1( u2_u0_u2_n110 ) , .ZN( u2_u0_u2_n111 ) , .C1( u2_u0_u2_n134 ) , .C2( u2_u0_u2_n170 ) , .B2( u2_u0_u2_n173 ) );
  OAI22_X1 u2_u0_u2_U9 (.ZN( u2_u0_u2_n109 ) , .A2( u2_u0_u2_n113 ) , .B2( u2_u0_u2_n133 ) , .B1( u2_u0_u2_n167 ) , .A1( u2_u0_u2_n168 ) );
  AOI21_X1 u2_u0_u2_U90 (.ZN( u2_u0_u2_n112 ) , .B2( u2_u0_u2_n156 ) , .A( u2_u0_u2_n164 ) , .B1( u2_u0_u2_n181 ) );
  NAND4_X1 u2_u0_u2_U91 (.ZN( u2_out0_16 ) , .A4( u2_u0_u2_n128 ) , .A3( u2_u0_u2_n129 ) , .A1( u2_u0_u2_n130 ) , .A2( u2_u0_u2_n186 ) );
  AOI22_X1 u2_u0_u2_U92 (.A2( u2_u0_u2_n118 ) , .ZN( u2_u0_u2_n129 ) , .A1( u2_u0_u2_n140 ) , .B1( u2_u0_u2_n157 ) , .B2( u2_u0_u2_n170 ) );
  INV_X1 u2_u0_u2_U93 (.A( u2_u0_u2_n163 ) , .ZN( u2_u0_u2_n186 ) );
  OR4_X1 u2_u0_u2_U94 (.ZN( u2_out0_6 ) , .A4( u2_u0_u2_n161 ) , .A3( u2_u0_u2_n162 ) , .A2( u2_u0_u2_n163 ) , .A1( u2_u0_u2_n164 ) );
  OR3_X1 u2_u0_u2_U95 (.A2( u2_u0_u2_n159 ) , .A1( u2_u0_u2_n160 ) , .ZN( u2_u0_u2_n161 ) , .A3( u2_u0_u2_n183 ) );
  AOI21_X1 u2_u0_u2_U96 (.B2( u2_u0_u2_n154 ) , .B1( u2_u0_u2_n155 ) , .ZN( u2_u0_u2_n159 ) , .A( u2_u0_u2_n167 ) );
  NAND3_X1 u2_u0_u2_U97 (.A2( u2_u0_u2_n117 ) , .A1( u2_u0_u2_n122 ) , .A3( u2_u0_u2_n123 ) , .ZN( u2_u0_u2_n134 ) );
  NAND3_X1 u2_u0_u2_U98 (.ZN( u2_u0_u2_n110 ) , .A2( u2_u0_u2_n131 ) , .A3( u2_u0_u2_n139 ) , .A1( u2_u0_u2_n154 ) );
  NAND3_X1 u2_u0_u2_U99 (.A2( u2_u0_u2_n100 ) , .ZN( u2_u0_u2_n101 ) , .A1( u2_u0_u2_n104 ) , .A3( u2_u0_u2_n114 ) );
  OAI211_X1 u2_u0_u3_U10 (.B( u2_u0_u3_n106 ) , .ZN( u2_u0_u3_n119 ) , .C2( u2_u0_u3_n128 ) , .C1( u2_u0_u3_n167 ) , .A( u2_u0_u3_n181 ) );
  AOI221_X1 u2_u0_u3_U11 (.C1( u2_u0_u3_n105 ) , .ZN( u2_u0_u3_n106 ) , .A( u2_u0_u3_n131 ) , .B2( u2_u0_u3_n132 ) , .C2( u2_u0_u3_n133 ) , .B1( u2_u0_u3_n169 ) );
  INV_X1 u2_u0_u3_U12 (.ZN( u2_u0_u3_n181 ) , .A( u2_u0_u3_n98 ) );
  NAND2_X1 u2_u0_u3_U13 (.ZN( u2_u0_u3_n105 ) , .A2( u2_u0_u3_n130 ) , .A1( u2_u0_u3_n155 ) );
  AOI22_X1 u2_u0_u3_U14 (.B1( u2_u0_u3_n115 ) , .A2( u2_u0_u3_n116 ) , .ZN( u2_u0_u3_n123 ) , .B2( u2_u0_u3_n133 ) , .A1( u2_u0_u3_n169 ) );
  NAND2_X1 u2_u0_u3_U15 (.ZN( u2_u0_u3_n116 ) , .A2( u2_u0_u3_n151 ) , .A1( u2_u0_u3_n182 ) );
  NOR2_X1 u2_u0_u3_U16 (.ZN( u2_u0_u3_n126 ) , .A2( u2_u0_u3_n150 ) , .A1( u2_u0_u3_n164 ) );
  AOI21_X1 u2_u0_u3_U17 (.ZN( u2_u0_u3_n112 ) , .B2( u2_u0_u3_n146 ) , .B1( u2_u0_u3_n155 ) , .A( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U18 (.A1( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n142 ) , .A2( u2_u0_u3_n164 ) );
  NAND2_X1 u2_u0_u3_U19 (.ZN( u2_u0_u3_n132 ) , .A2( u2_u0_u3_n152 ) , .A1( u2_u0_u3_n156 ) );
  INV_X1 u2_u0_u3_U20 (.A( u2_u0_u3_n133 ) , .ZN( u2_u0_u3_n165 ) );
  AND2_X1 u2_u0_u3_U21 (.A2( u2_u0_u3_n113 ) , .A1( u2_u0_u3_n114 ) , .ZN( u2_u0_u3_n151 ) );
  INV_X1 u2_u0_u3_U22 (.A( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n170 ) );
  NAND2_X1 u2_u0_u3_U23 (.A1( u2_u0_u3_n107 ) , .A2( u2_u0_u3_n108 ) , .ZN( u2_u0_u3_n140 ) );
  NAND2_X1 u2_u0_u3_U24 (.ZN( u2_u0_u3_n117 ) , .A1( u2_u0_u3_n124 ) , .A2( u2_u0_u3_n148 ) );
  INV_X1 u2_u0_u3_U25 (.A( u2_u0_u3_n128 ) , .ZN( u2_u0_u3_n176 ) );
  INV_X1 u2_u0_u3_U26 (.A( u2_u0_u3_n155 ) , .ZN( u2_u0_u3_n174 ) );
  INV_X1 u2_u0_u3_U27 (.A( u2_u0_u3_n130 ) , .ZN( u2_u0_u3_n177 ) );
  INV_X1 u2_u0_u3_U28 (.A( u2_u0_u3_n139 ) , .ZN( u2_u0_u3_n185 ) );
  NOR2_X1 u2_u0_u3_U29 (.ZN( u2_u0_u3_n135 ) , .A2( u2_u0_u3_n141 ) , .A1( u2_u0_u3_n169 ) );
  INV_X1 u2_u0_u3_U3 (.A( u2_u0_u3_n140 ) , .ZN( u2_u0_u3_n182 ) );
  OAI222_X1 u2_u0_u3_U30 (.C2( u2_u0_u3_n107 ) , .A2( u2_u0_u3_n108 ) , .B1( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n138 ) , .B2( u2_u0_u3_n146 ) , .C1( u2_u0_u3_n154 ) , .A1( u2_u0_u3_n164 ) );
  NOR4_X1 u2_u0_u3_U31 (.A4( u2_u0_u3_n157 ) , .A3( u2_u0_u3_n158 ) , .A2( u2_u0_u3_n159 ) , .A1( u2_u0_u3_n160 ) , .ZN( u2_u0_u3_n161 ) );
  AOI21_X1 u2_u0_u3_U32 (.B2( u2_u0_u3_n152 ) , .B1( u2_u0_u3_n153 ) , .ZN( u2_u0_u3_n158 ) , .A( u2_u0_u3_n164 ) );
  AOI21_X1 u2_u0_u3_U33 (.A( u2_u0_u3_n154 ) , .B2( u2_u0_u3_n155 ) , .B1( u2_u0_u3_n156 ) , .ZN( u2_u0_u3_n157 ) );
  AOI21_X1 u2_u0_u3_U34 (.A( u2_u0_u3_n149 ) , .B2( u2_u0_u3_n150 ) , .B1( u2_u0_u3_n151 ) , .ZN( u2_u0_u3_n159 ) );
  AOI211_X1 u2_u0_u3_U35 (.ZN( u2_u0_u3_n109 ) , .A( u2_u0_u3_n119 ) , .C2( u2_u0_u3_n129 ) , .B( u2_u0_u3_n138 ) , .C1( u2_u0_u3_n141 ) );
  AOI211_X1 u2_u0_u3_U36 (.B( u2_u0_u3_n119 ) , .A( u2_u0_u3_n120 ) , .C2( u2_u0_u3_n121 ) , .ZN( u2_u0_u3_n122 ) , .C1( u2_u0_u3_n179 ) );
  INV_X1 u2_u0_u3_U37 (.A( u2_u0_u3_n156 ) , .ZN( u2_u0_u3_n179 ) );
  OAI22_X1 u2_u0_u3_U38 (.B1( u2_u0_u3_n118 ) , .ZN( u2_u0_u3_n120 ) , .A1( u2_u0_u3_n135 ) , .B2( u2_u0_u3_n154 ) , .A2( u2_u0_u3_n178 ) );
  AND3_X1 u2_u0_u3_U39 (.ZN( u2_u0_u3_n118 ) , .A2( u2_u0_u3_n124 ) , .A1( u2_u0_u3_n144 ) , .A3( u2_u0_u3_n152 ) );
  INV_X1 u2_u0_u3_U4 (.A( u2_u0_u3_n129 ) , .ZN( u2_u0_u3_n183 ) );
  INV_X1 u2_u0_u3_U40 (.A( u2_u0_u3_n121 ) , .ZN( u2_u0_u3_n164 ) );
  OAI211_X1 u2_u0_u3_U41 (.B( u2_u0_u3_n127 ) , .ZN( u2_u0_u3_n139 ) , .C1( u2_u0_u3_n150 ) , .C2( u2_u0_u3_n154 ) , .A( u2_u0_u3_n184 ) );
  INV_X1 u2_u0_u3_U42 (.A( u2_u0_u3_n125 ) , .ZN( u2_u0_u3_n184 ) );
  AOI221_X1 u2_u0_u3_U43 (.A( u2_u0_u3_n126 ) , .ZN( u2_u0_u3_n127 ) , .C2( u2_u0_u3_n132 ) , .C1( u2_u0_u3_n169 ) , .B2( u2_u0_u3_n170 ) , .B1( u2_u0_u3_n174 ) );
  OAI22_X1 u2_u0_u3_U44 (.A1( u2_u0_u3_n124 ) , .ZN( u2_u0_u3_n125 ) , .B2( u2_u0_u3_n145 ) , .A2( u2_u0_u3_n165 ) , .B1( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U45 (.A1( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n150 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U46 (.A2( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n155 ) , .A1( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U47 (.ZN( u2_u0_u3_n133 ) , .A1( u2_u0_u3_n154 ) , .A2( u2_u0_u3_n164 ) );
  NOR2_X1 u2_u0_u3_U48 (.A1( u2_u0_u3_n113 ) , .ZN( u2_u0_u3_n131 ) , .A2( u2_u0_u3_n154 ) );
  AOI21_X1 u2_u0_u3_U49 (.B2( u2_u0_u3_n114 ) , .B1( u2_u0_u3_n146 ) , .A( u2_u0_u3_n154 ) , .ZN( u2_u0_u3_n94 ) );
  INV_X1 u2_u0_u3_U5 (.A( u2_u0_u3_n117 ) , .ZN( u2_u0_u3_n178 ) );
  AOI21_X1 u2_u0_u3_U50 (.ZN( u2_u0_u3_n110 ) , .B2( u2_u0_u3_n142 ) , .B1( u2_u0_u3_n186 ) , .A( u2_u0_u3_n95 ) );
  INV_X1 u2_u0_u3_U51 (.A( u2_u0_u3_n145 ) , .ZN( u2_u0_u3_n186 ) );
  AOI21_X1 u2_u0_u3_U52 (.B1( u2_u0_u3_n124 ) , .A( u2_u0_u3_n149 ) , .B2( u2_u0_u3_n155 ) , .ZN( u2_u0_u3_n95 ) );
  INV_X1 u2_u0_u3_U53 (.A( u2_u0_u3_n141 ) , .ZN( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U54 (.ZN( u2_u0_u3_n124 ) , .A1( u2_u0_u3_n96 ) , .A2( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U55 (.A2( u2_u0_u3_n100 ) , .ZN( u2_u0_u3_n146 ) , .A1( u2_u0_u3_n96 ) );
  INV_X1 u2_u0_u3_U56 (.A( u2_u0_u3_n149 ) , .ZN( u2_u0_u3_n169 ) );
  NAND2_X1 u2_u0_u3_U57 (.A1( u2_u0_u3_n101 ) , .ZN( u2_u0_u3_n145 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U58 (.A1( u2_u0_u3_n100 ) , .ZN( u2_u0_u3_n156 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U59 (.A2( u2_u0_u3_n101 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n148 ) );
  OAI22_X1 u2_u0_u3_U6 (.B2( u2_u0_u3_n147 ) , .A2( u2_u0_u3_n148 ) , .ZN( u2_u0_u3_n160 ) , .B1( u2_u0_u3_n165 ) , .A1( u2_u0_u3_n168 ) );
  NAND2_X1 u2_u0_u3_U60 (.A1( u2_u0_u3_n100 ) , .A2( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n128 ) );
  NAND2_X1 u2_u0_u3_U61 (.A2( u2_u0_u3_n101 ) , .A1( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n152 ) );
  NAND2_X1 u2_u0_u3_U62 (.A2( u2_u0_u3_n101 ) , .ZN( u2_u0_u3_n114 ) , .A1( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U63 (.ZN( u2_u0_u3_n107 ) , .A1( u2_u0_u3_n97 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U64 (.A2( u2_u0_u3_n100 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n113 ) );
  NAND2_X1 u2_u0_u3_U65 (.A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n153 ) , .A2( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U66 (.A2( u2_u0_u3_n103 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n130 ) );
  NAND2_X1 u2_u0_u3_U67 (.A2( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n144 ) , .A1( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U68 (.A1( u2_u0_u3_n102 ) , .A2( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n108 ) );
  NOR2_X1 u2_u0_u3_U69 (.A2( u2_u0_X_19 ) , .A1( u2_u0_X_20 ) , .ZN( u2_u0_u3_n99 ) );
  AND3_X1 u2_u0_u3_U7 (.A3( u2_u0_u3_n144 ) , .A2( u2_u0_u3_n145 ) , .A1( u2_u0_u3_n146 ) , .ZN( u2_u0_u3_n147 ) );
  NOR2_X1 u2_u0_u3_U70 (.A2( u2_u0_X_21 ) , .A1( u2_u0_X_24 ) , .ZN( u2_u0_u3_n103 ) );
  NOR2_X1 u2_u0_u3_U71 (.A2( u2_u0_X_24 ) , .A1( u2_u0_u3_n171 ) , .ZN( u2_u0_u3_n97 ) );
  NOR2_X1 u2_u0_u3_U72 (.A2( u2_u0_X_23 ) , .ZN( u2_u0_u3_n141 ) , .A1( u2_u0_u3_n166 ) );
  NOR2_X1 u2_u0_u3_U73 (.A2( u2_u0_X_19 ) , .A1( u2_u0_u3_n172 ) , .ZN( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U74 (.A1( u2_u0_X_22 ) , .A2( u2_u0_X_23 ) , .ZN( u2_u0_u3_n154 ) );
  NOR2_X1 u2_u0_u3_U75 (.A2( u2_u0_X_22 ) , .A1( u2_u0_X_23 ) , .ZN( u2_u0_u3_n121 ) );
  AND2_X1 u2_u0_u3_U76 (.A1( u2_u0_X_24 ) , .ZN( u2_u0_u3_n101 ) , .A2( u2_u0_u3_n171 ) );
  NAND2_X1 u2_u0_u3_U77 (.A1( u2_u0_X_23 ) , .ZN( u2_u0_u3_n149 ) , .A2( u2_u0_u3_n166 ) );
  AND2_X1 u2_u0_u3_U78 (.A1( u2_u0_X_19 ) , .ZN( u2_u0_u3_n102 ) , .A2( u2_u0_u3_n172 ) );
  AND2_X1 u2_u0_u3_U79 (.A1( u2_u0_X_21 ) , .A2( u2_u0_X_24 ) , .ZN( u2_u0_u3_n100 ) );
  INV_X1 u2_u0_u3_U8 (.A( u2_u0_u3_n143 ) , .ZN( u2_u0_u3_n168 ) );
  AND2_X1 u2_u0_u3_U80 (.A2( u2_u0_X_19 ) , .A1( u2_u0_X_20 ) , .ZN( u2_u0_u3_n104 ) );
  INV_X1 u2_u0_u3_U81 (.A( u2_u0_X_22 ) , .ZN( u2_u0_u3_n166 ) );
  INV_X1 u2_u0_u3_U82 (.A( u2_u0_X_21 ) , .ZN( u2_u0_u3_n171 ) );
  INV_X1 u2_u0_u3_U83 (.A( u2_u0_X_20 ) , .ZN( u2_u0_u3_n172 ) );
  NAND4_X1 u2_u0_u3_U84 (.ZN( u2_out0_26 ) , .A4( u2_u0_u3_n109 ) , .A3( u2_u0_u3_n110 ) , .A2( u2_u0_u3_n111 ) , .A1( u2_u0_u3_n173 ) );
  INV_X1 u2_u0_u3_U85 (.ZN( u2_u0_u3_n173 ) , .A( u2_u0_u3_n94 ) );
  OAI21_X1 u2_u0_u3_U86 (.ZN( u2_u0_u3_n111 ) , .B2( u2_u0_u3_n117 ) , .A( u2_u0_u3_n133 ) , .B1( u2_u0_u3_n176 ) );
  NAND4_X1 u2_u0_u3_U87 (.ZN( u2_out0_20 ) , .A4( u2_u0_u3_n122 ) , .A3( u2_u0_u3_n123 ) , .A1( u2_u0_u3_n175 ) , .A2( u2_u0_u3_n180 ) );
  INV_X1 u2_u0_u3_U88 (.A( u2_u0_u3_n126 ) , .ZN( u2_u0_u3_n180 ) );
  INV_X1 u2_u0_u3_U89 (.A( u2_u0_u3_n112 ) , .ZN( u2_u0_u3_n175 ) );
  OAI22_X1 u2_u0_u3_U9 (.B1( u2_u0_u3_n113 ) , .A2( u2_u0_u3_n135 ) , .A1( u2_u0_u3_n150 ) , .B2( u2_u0_u3_n164 ) , .ZN( u2_u0_u3_n98 ) );
  NAND4_X1 u2_u0_u3_U90 (.ZN( u2_out0_1 ) , .A4( u2_u0_u3_n161 ) , .A3( u2_u0_u3_n162 ) , .A2( u2_u0_u3_n163 ) , .A1( u2_u0_u3_n185 ) );
  NAND2_X1 u2_u0_u3_U91 (.ZN( u2_u0_u3_n163 ) , .A2( u2_u0_u3_n170 ) , .A1( u2_u0_u3_n176 ) );
  AOI22_X1 u2_u0_u3_U92 (.B2( u2_u0_u3_n140 ) , .B1( u2_u0_u3_n141 ) , .A2( u2_u0_u3_n142 ) , .ZN( u2_u0_u3_n162 ) , .A1( u2_u0_u3_n177 ) );
  OR4_X1 u2_u0_u3_U93 (.ZN( u2_out0_10 ) , .A4( u2_u0_u3_n136 ) , .A3( u2_u0_u3_n137 ) , .A1( u2_u0_u3_n138 ) , .A2( u2_u0_u3_n139 ) );
  OAI222_X1 u2_u0_u3_U94 (.C1( u2_u0_u3_n128 ) , .ZN( u2_u0_u3_n137 ) , .B1( u2_u0_u3_n148 ) , .A2( u2_u0_u3_n150 ) , .B2( u2_u0_u3_n154 ) , .C2( u2_u0_u3_n164 ) , .A1( u2_u0_u3_n167 ) );
  OAI221_X1 u2_u0_u3_U95 (.A( u2_u0_u3_n134 ) , .B2( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n136 ) , .C1( u2_u0_u3_n149 ) , .B1( u2_u0_u3_n151 ) , .C2( u2_u0_u3_n183 ) );
  AOI221_X1 u2_u0_u3_U96 (.A( u2_u0_u3_n131 ) , .C2( u2_u0_u3_n132 ) , .C1( u2_u0_u3_n133 ) , .ZN( u2_u0_u3_n134 ) , .B1( u2_u0_u3_n143 ) , .B2( u2_u0_u3_n177 ) );
  NAND2_X1 u2_u0_u3_U97 (.ZN( u2_u0_u3_n143 ) , .A1( u2_u0_u3_n165 ) , .A2( u2_u0_u3_n167 ) );
  NAND3_X1 u2_u0_u3_U98 (.A1( u2_u0_u3_n114 ) , .ZN( u2_u0_u3_n115 ) , .A2( u2_u0_u3_n145 ) , .A3( u2_u0_u3_n153 ) );
  NAND3_X1 u2_u0_u3_U99 (.ZN( u2_u0_u3_n129 ) , .A2( u2_u0_u3_n144 ) , .A1( u2_u0_u3_n153 ) , .A3( u2_u0_u3_n182 ) );
  XOR2_X1 u2_u10_U1 (.B( u2_K11_9 ) , .A( u2_R9_6 ) , .Z( u2_u10_X_9 ) );
  XOR2_X1 u2_u10_U10 (.B( u2_K11_45 ) , .A( u2_R9_30 ) , .Z( u2_u10_X_45 ) );
  XOR2_X1 u2_u10_U11 (.B( u2_K11_44 ) , .A( u2_R9_29 ) , .Z( u2_u10_X_44 ) );
  XOR2_X1 u2_u10_U12 (.B( u2_K11_43 ) , .A( u2_R9_28 ) , .Z( u2_u10_X_43 ) );
  XOR2_X1 u2_u10_U13 (.B( u2_K11_42 ) , .A( u2_R9_29 ) , .Z( u2_u10_X_42 ) );
  XOR2_X1 u2_u10_U14 (.B( u2_K11_41 ) , .A( u2_R9_28 ) , .Z( u2_u10_X_41 ) );
  XOR2_X1 u2_u10_U15 (.B( u2_K11_40 ) , .A( u2_R9_27 ) , .Z( u2_u10_X_40 ) );
  XOR2_X1 u2_u10_U16 (.B( u2_K11_3 ) , .A( u2_R9_2 ) , .Z( u2_u10_X_3 ) );
  XOR2_X1 u2_u10_U17 (.B( u2_K11_39 ) , .A( u2_R9_26 ) , .Z( u2_u10_X_39 ) );
  XOR2_X1 u2_u10_U18 (.B( u2_K11_38 ) , .A( u2_R9_25 ) , .Z( u2_u10_X_38 ) );
  XOR2_X1 u2_u10_U19 (.B( u2_K11_37 ) , .A( u2_R9_24 ) , .Z( u2_u10_X_37 ) );
  XOR2_X1 u2_u10_U2 (.B( u2_K11_8 ) , .A( u2_R9_5 ) , .Z( u2_u10_X_8 ) );
  XOR2_X1 u2_u10_U20 (.B( u2_K11_36 ) , .A( u2_R9_25 ) , .Z( u2_u10_X_36 ) );
  XOR2_X1 u2_u10_U21 (.B( u2_K11_35 ) , .A( u2_R9_24 ) , .Z( u2_u10_X_35 ) );
  XOR2_X1 u2_u10_U22 (.B( u2_K11_34 ) , .A( u2_R9_23 ) , .Z( u2_u10_X_34 ) );
  XOR2_X1 u2_u10_U23 (.B( u2_K11_33 ) , .A( u2_R9_22 ) , .Z( u2_u10_X_33 ) );
  XOR2_X1 u2_u10_U24 (.B( u2_K11_32 ) , .A( u2_R9_21 ) , .Z( u2_u10_X_32 ) );
  XOR2_X1 u2_u10_U26 (.B( u2_K11_30 ) , .A( u2_R9_21 ) , .Z( u2_u10_X_30 ) );
  XOR2_X1 u2_u10_U27 (.B( u2_K11_2 ) , .A( u2_R9_1 ) , .Z( u2_u10_X_2 ) );
  XOR2_X1 u2_u10_U29 (.B( u2_K11_28 ) , .A( u2_R9_19 ) , .Z( u2_u10_X_28 ) );
  XOR2_X1 u2_u10_U3 (.B( u2_K11_7 ) , .A( u2_R9_4 ) , .Z( u2_u10_X_7 ) );
  XOR2_X1 u2_u10_U30 (.B( u2_K11_27 ) , .A( u2_R9_18 ) , .Z( u2_u10_X_27 ) );
  XOR2_X1 u2_u10_U32 (.B( u2_K11_25 ) , .A( u2_R9_16 ) , .Z( u2_u10_X_25 ) );
  XOR2_X1 u2_u10_U34 (.B( u2_K11_23 ) , .A( u2_R9_16 ) , .Z( u2_u10_X_23 ) );
  XOR2_X1 u2_u10_U35 (.B( u2_K11_22 ) , .A( u2_R9_15 ) , .Z( u2_u10_X_22 ) );
  XOR2_X1 u2_u10_U36 (.B( u2_K11_21 ) , .A( u2_R9_14 ) , .Z( u2_u10_X_21 ) );
  XOR2_X1 u2_u10_U38 (.B( u2_K11_1 ) , .A( u2_R9_32 ) , .Z( u2_u10_X_1 ) );
  XOR2_X1 u2_u10_U4 (.B( u2_K11_6 ) , .A( u2_R9_5 ) , .Z( u2_u10_X_6 ) );
  XOR2_X1 u2_u10_U40 (.B( u2_K11_18 ) , .A( u2_R9_13 ) , .Z( u2_u10_X_18 ) );
  XOR2_X1 u2_u10_U42 (.B( u2_K11_16 ) , .A( u2_R9_11 ) , .Z( u2_u10_X_16 ) );
  XOR2_X1 u2_u10_U43 (.B( u2_K11_15 ) , .A( u2_R9_10 ) , .Z( u2_u10_X_15 ) );
  XOR2_X1 u2_u10_U48 (.B( u2_K11_10 ) , .A( u2_R9_7 ) , .Z( u2_u10_X_10 ) );
  XOR2_X1 u2_u10_U5 (.B( u2_K11_5 ) , .A( u2_R9_4 ) , .Z( u2_u10_X_5 ) );
  XOR2_X1 u2_u10_U6 (.B( u2_K11_4 ) , .A( u2_R9_3 ) , .Z( u2_u10_X_4 ) );
  XOR2_X1 u2_u10_U7 (.B( u2_K11_48 ) , .A( u2_R9_1 ) , .Z( u2_u10_X_48 ) );
  XOR2_X1 u2_u10_U9 (.B( u2_K11_46 ) , .A( u2_R9_31 ) , .Z( u2_u10_X_46 ) );
  AND3_X1 u2_u10_u0_U10 (.A2( u2_u10_u0_n112 ) , .ZN( u2_u10_u0_n127 ) , .A3( u2_u10_u0_n130 ) , .A1( u2_u10_u0_n148 ) );
  NAND2_X1 u2_u10_u0_U11 (.ZN( u2_u10_u0_n113 ) , .A1( u2_u10_u0_n139 ) , .A2( u2_u10_u0_n149 ) );
  AND2_X1 u2_u10_u0_U12 (.ZN( u2_u10_u0_n107 ) , .A1( u2_u10_u0_n130 ) , .A2( u2_u10_u0_n140 ) );
  AND2_X1 u2_u10_u0_U13 (.A2( u2_u10_u0_n129 ) , .A1( u2_u10_u0_n130 ) , .ZN( u2_u10_u0_n151 ) );
  AND2_X1 u2_u10_u0_U14 (.A1( u2_u10_u0_n108 ) , .A2( u2_u10_u0_n125 ) , .ZN( u2_u10_u0_n145 ) );
  INV_X1 u2_u10_u0_U15 (.A( u2_u10_u0_n143 ) , .ZN( u2_u10_u0_n173 ) );
  NOR2_X1 u2_u10_u0_U16 (.A2( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n147 ) , .A1( u2_u10_u0_n160 ) );
  NOR2_X1 u2_u10_u0_U17 (.A1( u2_u10_u0_n163 ) , .A2( u2_u10_u0_n164 ) , .ZN( u2_u10_u0_n95 ) );
  AOI21_X1 u2_u10_u0_U18 (.B1( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n132 ) , .A( u2_u10_u0_n165 ) , .B2( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U19 (.A( u2_u10_u0_n142 ) , .ZN( u2_u10_u0_n165 ) );
  OAI221_X1 u2_u10_u0_U20 (.C1( u2_u10_u0_n121 ) , .ZN( u2_u10_u0_n122 ) , .B2( u2_u10_u0_n127 ) , .A( u2_u10_u0_n143 ) , .B1( u2_u10_u0_n144 ) , .C2( u2_u10_u0_n147 ) );
  OAI22_X1 u2_u10_u0_U21 (.B1( u2_u10_u0_n125 ) , .ZN( u2_u10_u0_n126 ) , .A1( u2_u10_u0_n138 ) , .A2( u2_u10_u0_n146 ) , .B2( u2_u10_u0_n147 ) );
  OAI22_X1 u2_u10_u0_U22 (.B1( u2_u10_u0_n131 ) , .A1( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n147 ) , .A2( u2_u10_u0_n90 ) , .ZN( u2_u10_u0_n91 ) );
  AND3_X1 u2_u10_u0_U23 (.A3( u2_u10_u0_n121 ) , .A2( u2_u10_u0_n125 ) , .A1( u2_u10_u0_n148 ) , .ZN( u2_u10_u0_n90 ) );
  NAND2_X1 u2_u10_u0_U24 (.A1( u2_u10_u0_n100 ) , .A2( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n125 ) );
  INV_X1 u2_u10_u0_U25 (.A( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n161 ) );
  NOR2_X1 u2_u10_u0_U26 (.A1( u2_u10_u0_n120 ) , .ZN( u2_u10_u0_n143 ) , .A2( u2_u10_u0_n167 ) );
  OAI221_X1 u2_u10_u0_U27 (.C1( u2_u10_u0_n112 ) , .ZN( u2_u10_u0_n120 ) , .B1( u2_u10_u0_n138 ) , .B2( u2_u10_u0_n141 ) , .C2( u2_u10_u0_n147 ) , .A( u2_u10_u0_n172 ) );
  AOI211_X1 u2_u10_u0_U28 (.B( u2_u10_u0_n115 ) , .A( u2_u10_u0_n116 ) , .C2( u2_u10_u0_n117 ) , .C1( u2_u10_u0_n118 ) , .ZN( u2_u10_u0_n119 ) );
  AOI22_X1 u2_u10_u0_U29 (.B2( u2_u10_u0_n109 ) , .A2( u2_u10_u0_n110 ) , .ZN( u2_u10_u0_n111 ) , .B1( u2_u10_u0_n118 ) , .A1( u2_u10_u0_n160 ) );
  INV_X1 u2_u10_u0_U3 (.A( u2_u10_u0_n113 ) , .ZN( u2_u10_u0_n166 ) );
  NAND2_X1 u2_u10_u0_U30 (.A1( u2_u10_u0_n100 ) , .ZN( u2_u10_u0_n129 ) , .A2( u2_u10_u0_n95 ) );
  INV_X1 u2_u10_u0_U31 (.A( u2_u10_u0_n118 ) , .ZN( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U32 (.ZN( u2_u10_u0_n104 ) , .B1( u2_u10_u0_n107 ) , .B2( u2_u10_u0_n141 ) , .A( u2_u10_u0_n144 ) );
  AOI21_X1 u2_u10_u0_U33 (.B1( u2_u10_u0_n127 ) , .B2( u2_u10_u0_n129 ) , .A( u2_u10_u0_n138 ) , .ZN( u2_u10_u0_n96 ) );
  AOI21_X1 u2_u10_u0_U34 (.ZN( u2_u10_u0_n116 ) , .B2( u2_u10_u0_n142 ) , .A( u2_u10_u0_n144 ) , .B1( u2_u10_u0_n166 ) );
  NAND2_X1 u2_u10_u0_U35 (.A2( u2_u10_u0_n100 ) , .A1( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n139 ) );
  NAND2_X1 u2_u10_u0_U36 (.A2( u2_u10_u0_n100 ) , .ZN( u2_u10_u0_n131 ) , .A1( u2_u10_u0_n92 ) );
  NAND2_X1 u2_u10_u0_U37 (.A1( u2_u10_u0_n101 ) , .A2( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n150 ) );
  INV_X1 u2_u10_u0_U38 (.A( u2_u10_u0_n138 ) , .ZN( u2_u10_u0_n160 ) );
  NAND2_X1 u2_u10_u0_U39 (.A1( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n128 ) , .A2( u2_u10_u0_n95 ) );
  AOI21_X1 u2_u10_u0_U4 (.B1( u2_u10_u0_n114 ) , .ZN( u2_u10_u0_n115 ) , .B2( u2_u10_u0_n129 ) , .A( u2_u10_u0_n161 ) );
  NAND2_X1 u2_u10_u0_U40 (.ZN( u2_u10_u0_n148 ) , .A1( u2_u10_u0_n93 ) , .A2( u2_u10_u0_n95 ) );
  NAND2_X1 u2_u10_u0_U41 (.A2( u2_u10_u0_n102 ) , .A1( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n149 ) );
  NAND2_X1 u2_u10_u0_U42 (.A2( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n114 ) , .A1( u2_u10_u0_n92 ) );
  NAND2_X1 u2_u10_u0_U43 (.A2( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n121 ) , .A1( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U44 (.ZN( u2_u10_u0_n172 ) , .A( u2_u10_u0_n88 ) );
  OAI222_X1 u2_u10_u0_U45 (.C1( u2_u10_u0_n108 ) , .A1( u2_u10_u0_n125 ) , .B2( u2_u10_u0_n128 ) , .B1( u2_u10_u0_n144 ) , .A2( u2_u10_u0_n158 ) , .C2( u2_u10_u0_n161 ) , .ZN( u2_u10_u0_n88 ) );
  NAND2_X1 u2_u10_u0_U46 (.ZN( u2_u10_u0_n112 ) , .A2( u2_u10_u0_n92 ) , .A1( u2_u10_u0_n93 ) );
  OR3_X1 u2_u10_u0_U47 (.A3( u2_u10_u0_n152 ) , .A2( u2_u10_u0_n153 ) , .A1( u2_u10_u0_n154 ) , .ZN( u2_u10_u0_n155 ) );
  AOI21_X1 u2_u10_u0_U48 (.A( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n145 ) , .B1( u2_u10_u0_n146 ) , .ZN( u2_u10_u0_n154 ) );
  AOI21_X1 u2_u10_u0_U49 (.B2( u2_u10_u0_n150 ) , .B1( u2_u10_u0_n151 ) , .ZN( u2_u10_u0_n152 ) , .A( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U5 (.B2( u2_u10_u0_n131 ) , .ZN( u2_u10_u0_n134 ) , .B1( u2_u10_u0_n151 ) , .A( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U50 (.A( u2_u10_u0_n147 ) , .B2( u2_u10_u0_n148 ) , .B1( u2_u10_u0_n149 ) , .ZN( u2_u10_u0_n153 ) );
  INV_X1 u2_u10_u0_U51 (.ZN( u2_u10_u0_n171 ) , .A( u2_u10_u0_n99 ) );
  OAI211_X1 u2_u10_u0_U52 (.C2( u2_u10_u0_n140 ) , .C1( u2_u10_u0_n161 ) , .A( u2_u10_u0_n169 ) , .B( u2_u10_u0_n98 ) , .ZN( u2_u10_u0_n99 ) );
  AOI211_X1 u2_u10_u0_U53 (.C1( u2_u10_u0_n118 ) , .A( u2_u10_u0_n123 ) , .B( u2_u10_u0_n96 ) , .C2( u2_u10_u0_n97 ) , .ZN( u2_u10_u0_n98 ) );
  INV_X1 u2_u10_u0_U54 (.ZN( u2_u10_u0_n169 ) , .A( u2_u10_u0_n91 ) );
  NOR2_X1 u2_u10_u0_U55 (.A2( u2_u10_X_4 ) , .A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n118 ) );
  NOR2_X1 u2_u10_u0_U56 (.A2( u2_u10_X_2 ) , .ZN( u2_u10_u0_n103 ) , .A1( u2_u10_u0_n164 ) );
  NOR2_X1 u2_u10_u0_U57 (.A2( u2_u10_X_1 ) , .A1( u2_u10_X_2 ) , .ZN( u2_u10_u0_n92 ) );
  NOR2_X1 u2_u10_u0_U58 (.A2( u2_u10_X_1 ) , .ZN( u2_u10_u0_n101 ) , .A1( u2_u10_u0_n163 ) );
  NAND2_X1 u2_u10_u0_U59 (.A2( u2_u10_X_4 ) , .A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n144 ) );
  NOR2_X1 u2_u10_u0_U6 (.A1( u2_u10_u0_n108 ) , .ZN( u2_u10_u0_n123 ) , .A2( u2_u10_u0_n158 ) );
  NOR2_X1 u2_u10_u0_U60 (.A2( u2_u10_X_5 ) , .ZN( u2_u10_u0_n136 ) , .A1( u2_u10_u0_n159 ) );
  NAND2_X1 u2_u10_u0_U61 (.A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n138 ) , .A2( u2_u10_u0_n159 ) );
  AND2_X1 u2_u10_u0_U62 (.A2( u2_u10_X_3 ) , .A1( u2_u10_X_6 ) , .ZN( u2_u10_u0_n102 ) );
  AND2_X1 u2_u10_u0_U63 (.A1( u2_u10_X_6 ) , .A2( u2_u10_u0_n162 ) , .ZN( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U64 (.A( u2_u10_X_4 ) , .ZN( u2_u10_u0_n159 ) );
  INV_X1 u2_u10_u0_U65 (.A( u2_u10_X_1 ) , .ZN( u2_u10_u0_n164 ) );
  INV_X1 u2_u10_u0_U66 (.A( u2_u10_X_2 ) , .ZN( u2_u10_u0_n163 ) );
  INV_X1 u2_u10_u0_U67 (.A( u2_u10_X_3 ) , .ZN( u2_u10_u0_n162 ) );
  INV_X1 u2_u10_u0_U68 (.A( u2_u10_u0_n126 ) , .ZN( u2_u10_u0_n168 ) );
  AOI211_X1 u2_u10_u0_U69 (.B( u2_u10_u0_n133 ) , .A( u2_u10_u0_n134 ) , .C2( u2_u10_u0_n135 ) , .C1( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n137 ) );
  OAI21_X1 u2_u10_u0_U7 (.B1( u2_u10_u0_n150 ) , .B2( u2_u10_u0_n158 ) , .A( u2_u10_u0_n172 ) , .ZN( u2_u10_u0_n89 ) );
  INV_X1 u2_u10_u0_U70 (.ZN( u2_u10_u0_n174 ) , .A( u2_u10_u0_n89 ) );
  AOI211_X1 u2_u10_u0_U71 (.B( u2_u10_u0_n104 ) , .A( u2_u10_u0_n105 ) , .ZN( u2_u10_u0_n106 ) , .C2( u2_u10_u0_n113 ) , .C1( u2_u10_u0_n160 ) );
  OR4_X1 u2_u10_u0_U72 (.ZN( u2_out10_17 ) , .A4( u2_u10_u0_n122 ) , .A2( u2_u10_u0_n123 ) , .A1( u2_u10_u0_n124 ) , .A3( u2_u10_u0_n170 ) );
  AOI21_X1 u2_u10_u0_U73 (.B2( u2_u10_u0_n107 ) , .ZN( u2_u10_u0_n124 ) , .B1( u2_u10_u0_n128 ) , .A( u2_u10_u0_n161 ) );
  INV_X1 u2_u10_u0_U74 (.A( u2_u10_u0_n111 ) , .ZN( u2_u10_u0_n170 ) );
  OR4_X1 u2_u10_u0_U75 (.ZN( u2_out10_31 ) , .A4( u2_u10_u0_n155 ) , .A2( u2_u10_u0_n156 ) , .A1( u2_u10_u0_n157 ) , .A3( u2_u10_u0_n173 ) );
  AOI21_X1 u2_u10_u0_U76 (.A( u2_u10_u0_n138 ) , .B2( u2_u10_u0_n139 ) , .B1( u2_u10_u0_n140 ) , .ZN( u2_u10_u0_n157 ) );
  AOI21_X1 u2_u10_u0_U77 (.B2( u2_u10_u0_n141 ) , .B1( u2_u10_u0_n142 ) , .ZN( u2_u10_u0_n156 ) , .A( u2_u10_u0_n161 ) );
  AOI21_X1 u2_u10_u0_U78 (.B1( u2_u10_u0_n132 ) , .ZN( u2_u10_u0_n133 ) , .A( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n166 ) );
  OAI22_X1 u2_u10_u0_U79 (.ZN( u2_u10_u0_n105 ) , .A2( u2_u10_u0_n132 ) , .B1( u2_u10_u0_n146 ) , .A1( u2_u10_u0_n147 ) , .B2( u2_u10_u0_n161 ) );
  AND2_X1 u2_u10_u0_U8 (.A1( u2_u10_u0_n114 ) , .A2( u2_u10_u0_n121 ) , .ZN( u2_u10_u0_n146 ) );
  NAND2_X1 u2_u10_u0_U80 (.ZN( u2_u10_u0_n110 ) , .A2( u2_u10_u0_n132 ) , .A1( u2_u10_u0_n145 ) );
  INV_X1 u2_u10_u0_U81 (.A( u2_u10_u0_n119 ) , .ZN( u2_u10_u0_n167 ) );
  NAND2_X1 u2_u10_u0_U82 (.A2( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n140 ) , .A1( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U83 (.A1( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n130 ) , .A2( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U84 (.ZN( u2_u10_u0_n108 ) , .A1( u2_u10_u0_n92 ) , .A2( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U85 (.ZN( u2_u10_u0_n142 ) , .A1( u2_u10_u0_n94 ) , .A2( u2_u10_u0_n95 ) );
  NOR2_X1 u2_u10_u0_U86 (.A2( u2_u10_X_6 ) , .ZN( u2_u10_u0_n100 ) , .A1( u2_u10_u0_n162 ) );
  NOR2_X1 u2_u10_u0_U87 (.A2( u2_u10_X_3 ) , .A1( u2_u10_X_6 ) , .ZN( u2_u10_u0_n94 ) );
  NAND3_X1 u2_u10_u0_U88 (.ZN( u2_out10_23 ) , .A3( u2_u10_u0_n137 ) , .A1( u2_u10_u0_n168 ) , .A2( u2_u10_u0_n171 ) );
  NAND3_X1 u2_u10_u0_U89 (.A3( u2_u10_u0_n127 ) , .A2( u2_u10_u0_n128 ) , .ZN( u2_u10_u0_n135 ) , .A1( u2_u10_u0_n150 ) );
  AND2_X1 u2_u10_u0_U9 (.A1( u2_u10_u0_n131 ) , .ZN( u2_u10_u0_n141 ) , .A2( u2_u10_u0_n150 ) );
  NAND3_X1 u2_u10_u0_U90 (.ZN( u2_u10_u0_n117 ) , .A3( u2_u10_u0_n132 ) , .A2( u2_u10_u0_n139 ) , .A1( u2_u10_u0_n148 ) );
  NAND3_X1 u2_u10_u0_U91 (.ZN( u2_u10_u0_n109 ) , .A2( u2_u10_u0_n114 ) , .A3( u2_u10_u0_n140 ) , .A1( u2_u10_u0_n149 ) );
  NAND3_X1 u2_u10_u0_U92 (.ZN( u2_out10_9 ) , .A3( u2_u10_u0_n106 ) , .A2( u2_u10_u0_n171 ) , .A1( u2_u10_u0_n174 ) );
  NAND3_X1 u2_u10_u0_U93 (.A2( u2_u10_u0_n128 ) , .A1( u2_u10_u0_n132 ) , .A3( u2_u10_u0_n146 ) , .ZN( u2_u10_u0_n97 ) );
  XOR2_X1 u2_u11_U1 (.B( u2_K12_9 ) , .A( u2_R10_6 ) , .Z( u2_u11_X_9 ) );
  XOR2_X1 u2_u11_U10 (.B( u2_K12_45 ) , .A( u2_R10_30 ) , .Z( u2_u11_X_45 ) );
  XOR2_X1 u2_u11_U12 (.B( u2_K12_43 ) , .A( u2_R10_28 ) , .Z( u2_u11_X_43 ) );
  XOR2_X1 u2_u11_U14 (.B( u2_K12_41 ) , .A( u2_R10_28 ) , .Z( u2_u11_X_41 ) );
  XOR2_X1 u2_u11_U15 (.B( u2_K12_40 ) , .A( u2_R10_27 ) , .Z( u2_u11_X_40 ) );
  XOR2_X1 u2_u11_U16 (.B( u2_K12_3 ) , .A( u2_R10_2 ) , .Z( u2_u11_X_3 ) );
  XOR2_X1 u2_u11_U17 (.B( u2_K12_39 ) , .A( u2_R10_26 ) , .Z( u2_u11_X_39 ) );
  XOR2_X1 u2_u11_U19 (.B( u2_K12_37 ) , .A( u2_R10_24 ) , .Z( u2_u11_X_37 ) );
  XOR2_X1 u2_u11_U2 (.B( u2_K12_8 ) , .A( u2_R10_5 ) , .Z( u2_u11_X_8 ) );
  XOR2_X1 u2_u11_U21 (.B( u2_K12_35 ) , .A( u2_R10_24 ) , .Z( u2_u11_X_35 ) );
  XOR2_X1 u2_u11_U22 (.B( u2_K12_34 ) , .A( u2_R10_23 ) , .Z( u2_u11_X_34 ) );
  XOR2_X1 u2_u11_U23 (.B( u2_K12_33 ) , .A( u2_R10_22 ) , .Z( u2_u11_X_33 ) );
  XOR2_X1 u2_u11_U25 (.B( u2_K12_31 ) , .A( u2_R10_20 ) , .Z( u2_u11_X_31 ) );
  XOR2_X1 u2_u11_U28 (.B( u2_K12_29 ) , .A( u2_R10_20 ) , .Z( u2_u11_X_29 ) );
  XOR2_X1 u2_u11_U29 (.B( u2_K12_28 ) , .A( u2_R10_19 ) , .Z( u2_u11_X_28 ) );
  XOR2_X1 u2_u11_U30 (.B( u2_K12_27 ) , .A( u2_R10_18 ) , .Z( u2_u11_X_27 ) );
  XOR2_X1 u2_u11_U31 (.B( u2_K12_26 ) , .A( u2_R10_17 ) , .Z( u2_u11_X_26 ) );
  XOR2_X1 u2_u11_U33 (.B( u2_K12_24 ) , .A( u2_R10_17 ) , .Z( u2_u11_X_24 ) );
  XOR2_X1 u2_u11_U35 (.B( u2_K12_22 ) , .A( u2_R10_15 ) , .Z( u2_u11_X_22 ) );
  XOR2_X1 u2_u11_U36 (.B( u2_K12_21 ) , .A( u2_R10_14 ) , .Z( u2_u11_X_21 ) );
  XOR2_X1 u2_u11_U4 (.B( u2_K12_6 ) , .A( u2_R10_5 ) , .Z( u2_u11_X_6 ) );
  XOR2_X1 u2_u11_U42 (.B( u2_K12_16 ) , .A( u2_R10_11 ) , .Z( u2_u11_X_16 ) );
  XOR2_X1 u2_u11_U43 (.B( u2_K12_15 ) , .A( u2_R10_10 ) , .Z( u2_u11_X_15 ) );
  XOR2_X1 u2_u11_U9 (.B( u2_K12_46 ) , .A( u2_R10_31 ) , .Z( u2_u11_X_46 ) );
  XOR2_X1 u2_u12_U1 (.B( u2_K13_9 ) , .A( u2_R11_6 ) , .Z( u2_u12_X_9 ) );
  XOR2_X1 u2_u12_U10 (.B( u2_K13_45 ) , .A( u2_R11_30 ) , .Z( u2_u12_X_45 ) );
  XOR2_X1 u2_u12_U11 (.B( u2_K13_44 ) , .A( u2_R11_29 ) , .Z( u2_u12_X_44 ) );
  XOR2_X1 u2_u12_U12 (.B( u2_K13_43 ) , .A( u2_R11_28 ) , .Z( u2_u12_X_43 ) );
  XOR2_X1 u2_u12_U13 (.B( u2_K13_42 ) , .A( u2_R11_29 ) , .Z( u2_u12_X_42 ) );
  XOR2_X1 u2_u12_U14 (.B( u2_K13_41 ) , .A( u2_R11_28 ) , .Z( u2_u12_X_41 ) );
  XOR2_X1 u2_u12_U15 (.B( u2_K13_40 ) , .A( u2_R11_27 ) , .Z( u2_u12_X_40 ) );
  XOR2_X1 u2_u12_U16 (.B( u2_K13_3 ) , .A( u2_R11_2 ) , .Z( u2_u12_X_3 ) );
  XOR2_X1 u2_u12_U17 (.B( u2_K13_39 ) , .A( u2_R11_26 ) , .Z( u2_u12_X_39 ) );
  XOR2_X1 u2_u12_U18 (.B( u2_K13_38 ) , .A( u2_R11_25 ) , .Z( u2_u12_X_38 ) );
  XOR2_X1 u2_u12_U2 (.B( u2_K13_8 ) , .A( u2_R11_5 ) , .Z( u2_u12_X_8 ) );
  XOR2_X1 u2_u12_U20 (.B( u2_K13_36 ) , .A( u2_R11_25 ) , .Z( u2_u12_X_36 ) );
  XOR2_X1 u2_u12_U22 (.B( u2_K13_34 ) , .A( u2_R11_23 ) , .Z( u2_u12_X_34 ) );
  XOR2_X1 u2_u12_U23 (.B( u2_K13_33 ) , .A( u2_R11_22 ) , .Z( u2_u12_X_33 ) );
  XOR2_X1 u2_u12_U25 (.B( u2_K13_31 ) , .A( u2_R11_20 ) , .Z( u2_u12_X_31 ) );
  XOR2_X1 u2_u12_U28 (.B( u2_K13_29 ) , .A( u2_R11_20 ) , .Z( u2_u12_X_29 ) );
  XOR2_X1 u2_u12_U29 (.B( u2_K13_28 ) , .A( u2_R11_19 ) , .Z( u2_u12_X_28 ) );
  XOR2_X1 u2_u12_U30 (.B( u2_K13_27 ) , .A( u2_R11_18 ) , .Z( u2_u12_X_27 ) );
  XOR2_X1 u2_u12_U31 (.B( u2_K13_26 ) , .A( u2_R11_17 ) , .Z( u2_u12_X_26 ) );
  XOR2_X1 u2_u12_U32 (.B( u2_K13_25 ) , .A( u2_R11_16 ) , .Z( u2_u12_X_25 ) );
  XOR2_X1 u2_u12_U33 (.B( u2_K13_24 ) , .A( u2_R11_17 ) , .Z( u2_u12_X_24 ) );
  XOR2_X1 u2_u12_U34 (.B( u2_K13_23 ) , .A( u2_R11_16 ) , .Z( u2_u12_X_23 ) );
  XOR2_X1 u2_u12_U35 (.B( u2_K13_22 ) , .A( u2_R11_15 ) , .Z( u2_u12_X_22 ) );
  XOR2_X1 u2_u12_U36 (.B( u2_K13_21 ) , .A( u2_R11_14 ) , .Z( u2_u12_X_21 ) );
  XOR2_X1 u2_u12_U37 (.B( u2_K13_20 ) , .A( u2_R11_13 ) , .Z( u2_u12_X_20 ) );
  XOR2_X1 u2_u12_U38 (.B( u2_K13_1 ) , .A( u2_R11_32 ) , .Z( u2_u12_X_1 ) );
  XOR2_X1 u2_u12_U39 (.B( u2_K13_19 ) , .A( u2_R11_12 ) , .Z( u2_u12_X_19 ) );
  XOR2_X1 u2_u12_U4 (.B( u2_K13_6 ) , .A( u2_R11_5 ) , .Z( u2_u12_X_6 ) );
  XOR2_X1 u2_u12_U40 (.B( u2_K13_18 ) , .A( u2_R11_13 ) , .Z( u2_u12_X_18 ) );
  XOR2_X1 u2_u12_U41 (.B( u2_K13_17 ) , .A( u2_R11_12 ) , .Z( u2_u12_X_17 ) );
  XOR2_X1 u2_u12_U42 (.B( u2_K13_16 ) , .A( u2_R11_11 ) , .Z( u2_u12_X_16 ) );
  XOR2_X1 u2_u12_U43 (.B( u2_K13_15 ) , .A( u2_R11_10 ) , .Z( u2_u12_X_15 ) );
  XOR2_X1 u2_u12_U44 (.B( u2_K13_14 ) , .A( u2_R11_9 ) , .Z( u2_u12_X_14 ) );
  XOR2_X1 u2_u12_U45 (.B( u2_K13_13 ) , .A( u2_R11_8 ) , .Z( u2_u12_X_13 ) );
  XOR2_X1 u2_u12_U46 (.B( u2_K13_12 ) , .A( u2_R11_9 ) , .Z( u2_u12_X_12 ) );
  XOR2_X1 u2_u12_U47 (.B( u2_K13_11 ) , .A( u2_R11_8 ) , .Z( u2_u12_X_11 ) );
  XOR2_X1 u2_u12_U48 (.B( u2_K13_10 ) , .A( u2_R11_7 ) , .Z( u2_u12_X_10 ) );
  XOR2_X1 u2_u12_U6 (.B( u2_K13_4 ) , .A( u2_R11_3 ) , .Z( u2_u12_X_4 ) );
  XOR2_X1 u2_u12_U8 (.B( u2_K13_47 ) , .A( u2_R11_32 ) , .Z( u2_u12_X_47 ) );
  XOR2_X1 u2_u12_U9 (.B( u2_K13_46 ) , .A( u2_R11_31 ) , .Z( u2_u12_X_46 ) );
  OAI22_X1 u2_u12_u2_U10 (.B1( u2_u12_u2_n151 ) , .A2( u2_u12_u2_n152 ) , .A1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n160 ) , .B2( u2_u12_u2_n168 ) );
  NAND3_X1 u2_u12_u2_U100 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n98 ) );
  NOR3_X1 u2_u12_u2_U11 (.A1( u2_u12_u2_n150 ) , .ZN( u2_u12_u2_n151 ) , .A3( u2_u12_u2_n175 ) , .A2( u2_u12_u2_n188 ) );
  AOI21_X1 u2_u12_u2_U12 (.B2( u2_u12_u2_n123 ) , .ZN( u2_u12_u2_n125 ) , .A( u2_u12_u2_n171 ) , .B1( u2_u12_u2_n184 ) );
  INV_X1 u2_u12_u2_U13 (.A( u2_u12_u2_n150 ) , .ZN( u2_u12_u2_n184 ) );
  AOI21_X1 u2_u12_u2_U14 (.ZN( u2_u12_u2_n144 ) , .B2( u2_u12_u2_n155 ) , .A( u2_u12_u2_n172 ) , .B1( u2_u12_u2_n185 ) );
  AOI21_X1 u2_u12_u2_U15 (.B2( u2_u12_u2_n143 ) , .ZN( u2_u12_u2_n145 ) , .B1( u2_u12_u2_n152 ) , .A( u2_u12_u2_n171 ) );
  INV_X1 u2_u12_u2_U16 (.A( u2_u12_u2_n156 ) , .ZN( u2_u12_u2_n171 ) );
  INV_X1 u2_u12_u2_U17 (.A( u2_u12_u2_n120 ) , .ZN( u2_u12_u2_n188 ) );
  NAND2_X1 u2_u12_u2_U18 (.A2( u2_u12_u2_n122 ) , .ZN( u2_u12_u2_n150 ) , .A1( u2_u12_u2_n152 ) );
  INV_X1 u2_u12_u2_U19 (.A( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n170 ) );
  INV_X1 u2_u12_u2_U20 (.A( u2_u12_u2_n137 ) , .ZN( u2_u12_u2_n173 ) );
  NAND2_X1 u2_u12_u2_U21 (.A1( u2_u12_u2_n132 ) , .A2( u2_u12_u2_n139 ) , .ZN( u2_u12_u2_n157 ) );
  INV_X1 u2_u12_u2_U22 (.A( u2_u12_u2_n113 ) , .ZN( u2_u12_u2_n178 ) );
  INV_X1 u2_u12_u2_U23 (.A( u2_u12_u2_n139 ) , .ZN( u2_u12_u2_n175 ) );
  INV_X1 u2_u12_u2_U24 (.A( u2_u12_u2_n155 ) , .ZN( u2_u12_u2_n181 ) );
  INV_X1 u2_u12_u2_U25 (.A( u2_u12_u2_n119 ) , .ZN( u2_u12_u2_n177 ) );
  INV_X1 u2_u12_u2_U26 (.A( u2_u12_u2_n116 ) , .ZN( u2_u12_u2_n180 ) );
  INV_X1 u2_u12_u2_U27 (.A( u2_u12_u2_n131 ) , .ZN( u2_u12_u2_n179 ) );
  INV_X1 u2_u12_u2_U28 (.A( u2_u12_u2_n154 ) , .ZN( u2_u12_u2_n176 ) );
  NAND2_X1 u2_u12_u2_U29 (.A2( u2_u12_u2_n116 ) , .A1( u2_u12_u2_n117 ) , .ZN( u2_u12_u2_n118 ) );
  NOR2_X1 u2_u12_u2_U3 (.ZN( u2_u12_u2_n121 ) , .A2( u2_u12_u2_n177 ) , .A1( u2_u12_u2_n180 ) );
  INV_X1 u2_u12_u2_U30 (.A( u2_u12_u2_n132 ) , .ZN( u2_u12_u2_n182 ) );
  INV_X1 u2_u12_u2_U31 (.A( u2_u12_u2_n158 ) , .ZN( u2_u12_u2_n183 ) );
  OAI21_X1 u2_u12_u2_U32 (.A( u2_u12_u2_n156 ) , .B1( u2_u12_u2_n157 ) , .ZN( u2_u12_u2_n158 ) , .B2( u2_u12_u2_n179 ) );
  NOR2_X1 u2_u12_u2_U33 (.ZN( u2_u12_u2_n156 ) , .A1( u2_u12_u2_n166 ) , .A2( u2_u12_u2_n169 ) );
  NOR2_X1 u2_u12_u2_U34 (.A2( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n137 ) , .A1( u2_u12_u2_n140 ) );
  NOR2_X1 u2_u12_u2_U35 (.A2( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n153 ) , .A1( u2_u12_u2_n156 ) );
  AOI211_X1 u2_u12_u2_U36 (.ZN( u2_u12_u2_n130 ) , .C1( u2_u12_u2_n138 ) , .C2( u2_u12_u2_n179 ) , .B( u2_u12_u2_n96 ) , .A( u2_u12_u2_n97 ) );
  OAI22_X1 u2_u12_u2_U37 (.B1( u2_u12_u2_n133 ) , .A2( u2_u12_u2_n137 ) , .A1( u2_u12_u2_n152 ) , .B2( u2_u12_u2_n168 ) , .ZN( u2_u12_u2_n97 ) );
  OAI221_X1 u2_u12_u2_U38 (.B1( u2_u12_u2_n113 ) , .C1( u2_u12_u2_n132 ) , .A( u2_u12_u2_n149 ) , .B2( u2_u12_u2_n171 ) , .C2( u2_u12_u2_n172 ) , .ZN( u2_u12_u2_n96 ) );
  OAI221_X1 u2_u12_u2_U39 (.A( u2_u12_u2_n115 ) , .C2( u2_u12_u2_n123 ) , .B2( u2_u12_u2_n143 ) , .B1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n163 ) , .C1( u2_u12_u2_n168 ) );
  INV_X1 u2_u12_u2_U4 (.A( u2_u12_u2_n134 ) , .ZN( u2_u12_u2_n185 ) );
  OAI21_X1 u2_u12_u2_U40 (.A( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n115 ) , .B1( u2_u12_u2_n176 ) , .B2( u2_u12_u2_n178 ) );
  OAI221_X1 u2_u12_u2_U41 (.A( u2_u12_u2_n135 ) , .B2( u2_u12_u2_n136 ) , .B1( u2_u12_u2_n137 ) , .ZN( u2_u12_u2_n162 ) , .C2( u2_u12_u2_n167 ) , .C1( u2_u12_u2_n185 ) );
  AND3_X1 u2_u12_u2_U42 (.A3( u2_u12_u2_n131 ) , .A2( u2_u12_u2_n132 ) , .A1( u2_u12_u2_n133 ) , .ZN( u2_u12_u2_n136 ) );
  AOI22_X1 u2_u12_u2_U43 (.ZN( u2_u12_u2_n135 ) , .B1( u2_u12_u2_n140 ) , .A1( u2_u12_u2_n156 ) , .B2( u2_u12_u2_n180 ) , .A2( u2_u12_u2_n188 ) );
  AOI21_X1 u2_u12_u2_U44 (.ZN( u2_u12_u2_n149 ) , .B1( u2_u12_u2_n173 ) , .B2( u2_u12_u2_n188 ) , .A( u2_u12_u2_n95 ) );
  AND3_X1 u2_u12_u2_U45 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n156 ) , .ZN( u2_u12_u2_n95 ) );
  OAI21_X1 u2_u12_u2_U46 (.A( u2_u12_u2_n101 ) , .B2( u2_u12_u2_n121 ) , .B1( u2_u12_u2_n153 ) , .ZN( u2_u12_u2_n164 ) );
  NAND2_X1 u2_u12_u2_U47 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n155 ) );
  NAND2_X1 u2_u12_u2_U48 (.A2( u2_u12_u2_n105 ) , .A1( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n143 ) );
  NAND2_X1 u2_u12_u2_U49 (.A1( u2_u12_u2_n104 ) , .A2( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n152 ) );
  NOR4_X1 u2_u12_u2_U5 (.A4( u2_u12_u2_n124 ) , .A3( u2_u12_u2_n125 ) , .A2( u2_u12_u2_n126 ) , .A1( u2_u12_u2_n127 ) , .ZN( u2_u12_u2_n128 ) );
  NAND2_X1 u2_u12_u2_U50 (.A1( u2_u12_u2_n100 ) , .A2( u2_u12_u2_n105 ) , .ZN( u2_u12_u2_n132 ) );
  INV_X1 u2_u12_u2_U51 (.A( u2_u12_u2_n140 ) , .ZN( u2_u12_u2_n168 ) );
  INV_X1 u2_u12_u2_U52 (.A( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n167 ) );
  OAI21_X1 u2_u12_u2_U53 (.A( u2_u12_u2_n141 ) , .B2( u2_u12_u2_n142 ) , .ZN( u2_u12_u2_n146 ) , .B1( u2_u12_u2_n153 ) );
  OAI21_X1 u2_u12_u2_U54 (.A( u2_u12_u2_n140 ) , .ZN( u2_u12_u2_n141 ) , .B1( u2_u12_u2_n176 ) , .B2( u2_u12_u2_n177 ) );
  NOR3_X1 u2_u12_u2_U55 (.ZN( u2_u12_u2_n142 ) , .A3( u2_u12_u2_n175 ) , .A2( u2_u12_u2_n178 ) , .A1( u2_u12_u2_n181 ) );
  NAND2_X1 u2_u12_u2_U56 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n113 ) );
  NAND2_X1 u2_u12_u2_U57 (.A1( u2_u12_u2_n106 ) , .A2( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n131 ) );
  NAND2_X1 u2_u12_u2_U58 (.A1( u2_u12_u2_n103 ) , .A2( u2_u12_u2_n107 ) , .ZN( u2_u12_u2_n139 ) );
  NAND2_X1 u2_u12_u2_U59 (.A1( u2_u12_u2_n103 ) , .A2( u2_u12_u2_n105 ) , .ZN( u2_u12_u2_n133 ) );
  AOI21_X1 u2_u12_u2_U6 (.B2( u2_u12_u2_n119 ) , .ZN( u2_u12_u2_n127 ) , .A( u2_u12_u2_n137 ) , .B1( u2_u12_u2_n155 ) );
  NAND2_X1 u2_u12_u2_U60 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n103 ) , .ZN( u2_u12_u2_n154 ) );
  NAND2_X1 u2_u12_u2_U61 (.A2( u2_u12_u2_n103 ) , .A1( u2_u12_u2_n104 ) , .ZN( u2_u12_u2_n119 ) );
  NAND2_X1 u2_u12_u2_U62 (.A2( u2_u12_u2_n107 ) , .A1( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n123 ) );
  NAND2_X1 u2_u12_u2_U63 (.A1( u2_u12_u2_n104 ) , .A2( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n122 ) );
  INV_X1 u2_u12_u2_U64 (.A( u2_u12_u2_n114 ) , .ZN( u2_u12_u2_n172 ) );
  NAND2_X1 u2_u12_u2_U65 (.A2( u2_u12_u2_n100 ) , .A1( u2_u12_u2_n102 ) , .ZN( u2_u12_u2_n116 ) );
  NAND2_X1 u2_u12_u2_U66 (.A1( u2_u12_u2_n102 ) , .A2( u2_u12_u2_n108 ) , .ZN( u2_u12_u2_n120 ) );
  NAND2_X1 u2_u12_u2_U67 (.A2( u2_u12_u2_n105 ) , .A1( u2_u12_u2_n106 ) , .ZN( u2_u12_u2_n117 ) );
  INV_X1 u2_u12_u2_U68 (.ZN( u2_u12_u2_n187 ) , .A( u2_u12_u2_n99 ) );
  OAI21_X1 u2_u12_u2_U69 (.B1( u2_u12_u2_n137 ) , .B2( u2_u12_u2_n143 ) , .A( u2_u12_u2_n98 ) , .ZN( u2_u12_u2_n99 ) );
  AOI21_X1 u2_u12_u2_U7 (.ZN( u2_u12_u2_n124 ) , .B1( u2_u12_u2_n131 ) , .B2( u2_u12_u2_n143 ) , .A( u2_u12_u2_n172 ) );
  NOR2_X1 u2_u12_u2_U70 (.A2( u2_u12_X_16 ) , .ZN( u2_u12_u2_n140 ) , .A1( u2_u12_u2_n166 ) );
  NOR2_X1 u2_u12_u2_U71 (.A2( u2_u12_X_13 ) , .A1( u2_u12_X_14 ) , .ZN( u2_u12_u2_n100 ) );
  NOR2_X1 u2_u12_u2_U72 (.A2( u2_u12_X_16 ) , .A1( u2_u12_X_17 ) , .ZN( u2_u12_u2_n138 ) );
  NOR2_X1 u2_u12_u2_U73 (.A2( u2_u12_X_15 ) , .A1( u2_u12_X_18 ) , .ZN( u2_u12_u2_n104 ) );
  NOR2_X1 u2_u12_u2_U74 (.A2( u2_u12_X_14 ) , .ZN( u2_u12_u2_n103 ) , .A1( u2_u12_u2_n174 ) );
  NOR2_X1 u2_u12_u2_U75 (.A2( u2_u12_X_15 ) , .ZN( u2_u12_u2_n102 ) , .A1( u2_u12_u2_n165 ) );
  NOR2_X1 u2_u12_u2_U76 (.A2( u2_u12_X_17 ) , .ZN( u2_u12_u2_n114 ) , .A1( u2_u12_u2_n169 ) );
  AND2_X1 u2_u12_u2_U77 (.A1( u2_u12_X_15 ) , .ZN( u2_u12_u2_n105 ) , .A2( u2_u12_u2_n165 ) );
  AND2_X1 u2_u12_u2_U78 (.A2( u2_u12_X_15 ) , .A1( u2_u12_X_18 ) , .ZN( u2_u12_u2_n107 ) );
  AND2_X1 u2_u12_u2_U79 (.A1( u2_u12_X_14 ) , .ZN( u2_u12_u2_n106 ) , .A2( u2_u12_u2_n174 ) );
  AOI21_X1 u2_u12_u2_U8 (.B2( u2_u12_u2_n120 ) , .B1( u2_u12_u2_n121 ) , .ZN( u2_u12_u2_n126 ) , .A( u2_u12_u2_n167 ) );
  AND2_X1 u2_u12_u2_U80 (.A1( u2_u12_X_13 ) , .A2( u2_u12_X_14 ) , .ZN( u2_u12_u2_n108 ) );
  INV_X1 u2_u12_u2_U81 (.A( u2_u12_X_16 ) , .ZN( u2_u12_u2_n169 ) );
  INV_X1 u2_u12_u2_U82 (.A( u2_u12_X_17 ) , .ZN( u2_u12_u2_n166 ) );
  INV_X1 u2_u12_u2_U83 (.A( u2_u12_X_13 ) , .ZN( u2_u12_u2_n174 ) );
  INV_X1 u2_u12_u2_U84 (.A( u2_u12_X_18 ) , .ZN( u2_u12_u2_n165 ) );
  NAND4_X1 u2_u12_u2_U85 (.ZN( u2_out12_30 ) , .A4( u2_u12_u2_n147 ) , .A3( u2_u12_u2_n148 ) , .A2( u2_u12_u2_n149 ) , .A1( u2_u12_u2_n187 ) );
  AOI21_X1 u2_u12_u2_U86 (.B2( u2_u12_u2_n138 ) , .ZN( u2_u12_u2_n148 ) , .A( u2_u12_u2_n162 ) , .B1( u2_u12_u2_n182 ) );
  NOR3_X1 u2_u12_u2_U87 (.A3( u2_u12_u2_n144 ) , .A2( u2_u12_u2_n145 ) , .A1( u2_u12_u2_n146 ) , .ZN( u2_u12_u2_n147 ) );
  NAND4_X1 u2_u12_u2_U88 (.ZN( u2_out12_24 ) , .A4( u2_u12_u2_n111 ) , .A3( u2_u12_u2_n112 ) , .A1( u2_u12_u2_n130 ) , .A2( u2_u12_u2_n187 ) );
  AOI221_X1 u2_u12_u2_U89 (.A( u2_u12_u2_n109 ) , .B1( u2_u12_u2_n110 ) , .ZN( u2_u12_u2_n111 ) , .C1( u2_u12_u2_n134 ) , .C2( u2_u12_u2_n170 ) , .B2( u2_u12_u2_n173 ) );
  OAI22_X1 u2_u12_u2_U9 (.ZN( u2_u12_u2_n109 ) , .A2( u2_u12_u2_n113 ) , .B2( u2_u12_u2_n133 ) , .B1( u2_u12_u2_n167 ) , .A1( u2_u12_u2_n168 ) );
  AOI21_X1 u2_u12_u2_U90 (.ZN( u2_u12_u2_n112 ) , .B2( u2_u12_u2_n156 ) , .A( u2_u12_u2_n164 ) , .B1( u2_u12_u2_n181 ) );
  NAND4_X1 u2_u12_u2_U91 (.ZN( u2_out12_16 ) , .A4( u2_u12_u2_n128 ) , .A3( u2_u12_u2_n129 ) , .A1( u2_u12_u2_n130 ) , .A2( u2_u12_u2_n186 ) );
  AOI22_X1 u2_u12_u2_U92 (.A2( u2_u12_u2_n118 ) , .ZN( u2_u12_u2_n129 ) , .A1( u2_u12_u2_n140 ) , .B1( u2_u12_u2_n157 ) , .B2( u2_u12_u2_n170 ) );
  INV_X1 u2_u12_u2_U93 (.A( u2_u12_u2_n163 ) , .ZN( u2_u12_u2_n186 ) );
  OR4_X1 u2_u12_u2_U94 (.ZN( u2_out12_6 ) , .A4( u2_u12_u2_n161 ) , .A3( u2_u12_u2_n162 ) , .A2( u2_u12_u2_n163 ) , .A1( u2_u12_u2_n164 ) );
  OR3_X1 u2_u12_u2_U95 (.A2( u2_u12_u2_n159 ) , .A1( u2_u12_u2_n160 ) , .ZN( u2_u12_u2_n161 ) , .A3( u2_u12_u2_n183 ) );
  AOI21_X1 u2_u12_u2_U96 (.B2( u2_u12_u2_n154 ) , .B1( u2_u12_u2_n155 ) , .ZN( u2_u12_u2_n159 ) , .A( u2_u12_u2_n167 ) );
  NAND3_X1 u2_u12_u2_U97 (.A2( u2_u12_u2_n117 ) , .A1( u2_u12_u2_n122 ) , .A3( u2_u12_u2_n123 ) , .ZN( u2_u12_u2_n134 ) );
  NAND3_X1 u2_u12_u2_U98 (.ZN( u2_u12_u2_n110 ) , .A2( u2_u12_u2_n131 ) , .A3( u2_u12_u2_n139 ) , .A1( u2_u12_u2_n154 ) );
  NAND3_X1 u2_u12_u2_U99 (.A2( u2_u12_u2_n100 ) , .ZN( u2_u12_u2_n101 ) , .A1( u2_u12_u2_n104 ) , .A3( u2_u12_u2_n114 ) );
  OAI22_X1 u2_u12_u3_U10 (.B1( u2_u12_u3_n113 ) , .A2( u2_u12_u3_n135 ) , .A1( u2_u12_u3_n150 ) , .B2( u2_u12_u3_n164 ) , .ZN( u2_u12_u3_n98 ) );
  OAI211_X1 u2_u12_u3_U11 (.B( u2_u12_u3_n106 ) , .ZN( u2_u12_u3_n119 ) , .C2( u2_u12_u3_n128 ) , .C1( u2_u12_u3_n167 ) , .A( u2_u12_u3_n181 ) );
  AOI221_X1 u2_u12_u3_U12 (.C1( u2_u12_u3_n105 ) , .ZN( u2_u12_u3_n106 ) , .A( u2_u12_u3_n131 ) , .B2( u2_u12_u3_n132 ) , .C2( u2_u12_u3_n133 ) , .B1( u2_u12_u3_n169 ) );
  INV_X1 u2_u12_u3_U13 (.ZN( u2_u12_u3_n181 ) , .A( u2_u12_u3_n98 ) );
  NAND2_X1 u2_u12_u3_U14 (.ZN( u2_u12_u3_n105 ) , .A2( u2_u12_u3_n130 ) , .A1( u2_u12_u3_n155 ) );
  AOI22_X1 u2_u12_u3_U15 (.B1( u2_u12_u3_n115 ) , .A2( u2_u12_u3_n116 ) , .ZN( u2_u12_u3_n123 ) , .B2( u2_u12_u3_n133 ) , .A1( u2_u12_u3_n169 ) );
  NAND2_X1 u2_u12_u3_U16 (.ZN( u2_u12_u3_n116 ) , .A2( u2_u12_u3_n151 ) , .A1( u2_u12_u3_n182 ) );
  NOR2_X1 u2_u12_u3_U17 (.ZN( u2_u12_u3_n126 ) , .A2( u2_u12_u3_n150 ) , .A1( u2_u12_u3_n164 ) );
  AOI21_X1 u2_u12_u3_U18 (.ZN( u2_u12_u3_n112 ) , .B2( u2_u12_u3_n146 ) , .B1( u2_u12_u3_n155 ) , .A( u2_u12_u3_n167 ) );
  NAND2_X1 u2_u12_u3_U19 (.A1( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n142 ) , .A2( u2_u12_u3_n164 ) );
  NAND2_X1 u2_u12_u3_U20 (.ZN( u2_u12_u3_n132 ) , .A2( u2_u12_u3_n152 ) , .A1( u2_u12_u3_n156 ) );
  AND2_X1 u2_u12_u3_U21 (.A2( u2_u12_u3_n113 ) , .A1( u2_u12_u3_n114 ) , .ZN( u2_u12_u3_n151 ) );
  INV_X1 u2_u12_u3_U22 (.A( u2_u12_u3_n133 ) , .ZN( u2_u12_u3_n165 ) );
  INV_X1 u2_u12_u3_U23 (.A( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n170 ) );
  NAND2_X1 u2_u12_u3_U24 (.A1( u2_u12_u3_n107 ) , .A2( u2_u12_u3_n108 ) , .ZN( u2_u12_u3_n140 ) );
  NAND2_X1 u2_u12_u3_U25 (.ZN( u2_u12_u3_n117 ) , .A1( u2_u12_u3_n124 ) , .A2( u2_u12_u3_n148 ) );
  NAND2_X1 u2_u12_u3_U26 (.ZN( u2_u12_u3_n143 ) , .A1( u2_u12_u3_n165 ) , .A2( u2_u12_u3_n167 ) );
  INV_X1 u2_u12_u3_U27 (.A( u2_u12_u3_n130 ) , .ZN( u2_u12_u3_n177 ) );
  INV_X1 u2_u12_u3_U28 (.A( u2_u12_u3_n128 ) , .ZN( u2_u12_u3_n176 ) );
  INV_X1 u2_u12_u3_U29 (.A( u2_u12_u3_n155 ) , .ZN( u2_u12_u3_n174 ) );
  INV_X1 u2_u12_u3_U3 (.A( u2_u12_u3_n129 ) , .ZN( u2_u12_u3_n183 ) );
  INV_X1 u2_u12_u3_U30 (.A( u2_u12_u3_n139 ) , .ZN( u2_u12_u3_n185 ) );
  NOR2_X1 u2_u12_u3_U31 (.ZN( u2_u12_u3_n135 ) , .A2( u2_u12_u3_n141 ) , .A1( u2_u12_u3_n169 ) );
  OAI222_X1 u2_u12_u3_U32 (.C2( u2_u12_u3_n107 ) , .A2( u2_u12_u3_n108 ) , .B1( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n138 ) , .B2( u2_u12_u3_n146 ) , .C1( u2_u12_u3_n154 ) , .A1( u2_u12_u3_n164 ) );
  NOR4_X1 u2_u12_u3_U33 (.A4( u2_u12_u3_n157 ) , .A3( u2_u12_u3_n158 ) , .A2( u2_u12_u3_n159 ) , .A1( u2_u12_u3_n160 ) , .ZN( u2_u12_u3_n161 ) );
  AOI21_X1 u2_u12_u3_U34 (.B2( u2_u12_u3_n152 ) , .B1( u2_u12_u3_n153 ) , .ZN( u2_u12_u3_n158 ) , .A( u2_u12_u3_n164 ) );
  AOI21_X1 u2_u12_u3_U35 (.A( u2_u12_u3_n154 ) , .B2( u2_u12_u3_n155 ) , .B1( u2_u12_u3_n156 ) , .ZN( u2_u12_u3_n157 ) );
  AOI21_X1 u2_u12_u3_U36 (.A( u2_u12_u3_n149 ) , .B2( u2_u12_u3_n150 ) , .B1( u2_u12_u3_n151 ) , .ZN( u2_u12_u3_n159 ) );
  AOI211_X1 u2_u12_u3_U37 (.ZN( u2_u12_u3_n109 ) , .A( u2_u12_u3_n119 ) , .C2( u2_u12_u3_n129 ) , .B( u2_u12_u3_n138 ) , .C1( u2_u12_u3_n141 ) );
  AOI211_X1 u2_u12_u3_U38 (.B( u2_u12_u3_n119 ) , .A( u2_u12_u3_n120 ) , .C2( u2_u12_u3_n121 ) , .ZN( u2_u12_u3_n122 ) , .C1( u2_u12_u3_n179 ) );
  INV_X1 u2_u12_u3_U39 (.A( u2_u12_u3_n156 ) , .ZN( u2_u12_u3_n179 ) );
  INV_X1 u2_u12_u3_U4 (.A( u2_u12_u3_n140 ) , .ZN( u2_u12_u3_n182 ) );
  OAI22_X1 u2_u12_u3_U40 (.B1( u2_u12_u3_n118 ) , .ZN( u2_u12_u3_n120 ) , .A1( u2_u12_u3_n135 ) , .B2( u2_u12_u3_n154 ) , .A2( u2_u12_u3_n178 ) );
  AND3_X1 u2_u12_u3_U41 (.ZN( u2_u12_u3_n118 ) , .A2( u2_u12_u3_n124 ) , .A1( u2_u12_u3_n144 ) , .A3( u2_u12_u3_n152 ) );
  INV_X1 u2_u12_u3_U42 (.A( u2_u12_u3_n121 ) , .ZN( u2_u12_u3_n164 ) );
  NAND2_X1 u2_u12_u3_U43 (.ZN( u2_u12_u3_n133 ) , .A1( u2_u12_u3_n154 ) , .A2( u2_u12_u3_n164 ) );
  OAI211_X1 u2_u12_u3_U44 (.B( u2_u12_u3_n127 ) , .ZN( u2_u12_u3_n139 ) , .C1( u2_u12_u3_n150 ) , .C2( u2_u12_u3_n154 ) , .A( u2_u12_u3_n184 ) );
  INV_X1 u2_u12_u3_U45 (.A( u2_u12_u3_n125 ) , .ZN( u2_u12_u3_n184 ) );
  AOI221_X1 u2_u12_u3_U46 (.A( u2_u12_u3_n126 ) , .ZN( u2_u12_u3_n127 ) , .C2( u2_u12_u3_n132 ) , .C1( u2_u12_u3_n169 ) , .B2( u2_u12_u3_n170 ) , .B1( u2_u12_u3_n174 ) );
  OAI22_X1 u2_u12_u3_U47 (.A1( u2_u12_u3_n124 ) , .ZN( u2_u12_u3_n125 ) , .B2( u2_u12_u3_n145 ) , .A2( u2_u12_u3_n165 ) , .B1( u2_u12_u3_n167 ) );
  NOR2_X1 u2_u12_u3_U48 (.A1( u2_u12_u3_n113 ) , .ZN( u2_u12_u3_n131 ) , .A2( u2_u12_u3_n154 ) );
  NAND2_X1 u2_u12_u3_U49 (.A1( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n150 ) , .A2( u2_u12_u3_n99 ) );
  INV_X1 u2_u12_u3_U5 (.A( u2_u12_u3_n117 ) , .ZN( u2_u12_u3_n178 ) );
  NAND2_X1 u2_u12_u3_U50 (.A2( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n155 ) , .A1( u2_u12_u3_n97 ) );
  INV_X1 u2_u12_u3_U51 (.A( u2_u12_u3_n141 ) , .ZN( u2_u12_u3_n167 ) );
  AOI21_X1 u2_u12_u3_U52 (.B2( u2_u12_u3_n114 ) , .B1( u2_u12_u3_n146 ) , .A( u2_u12_u3_n154 ) , .ZN( u2_u12_u3_n94 ) );
  AOI21_X1 u2_u12_u3_U53 (.ZN( u2_u12_u3_n110 ) , .B2( u2_u12_u3_n142 ) , .B1( u2_u12_u3_n186 ) , .A( u2_u12_u3_n95 ) );
  INV_X1 u2_u12_u3_U54 (.A( u2_u12_u3_n145 ) , .ZN( u2_u12_u3_n186 ) );
  AOI21_X1 u2_u12_u3_U55 (.B1( u2_u12_u3_n124 ) , .A( u2_u12_u3_n149 ) , .B2( u2_u12_u3_n155 ) , .ZN( u2_u12_u3_n95 ) );
  INV_X1 u2_u12_u3_U56 (.A( u2_u12_u3_n149 ) , .ZN( u2_u12_u3_n169 ) );
  NAND2_X1 u2_u12_u3_U57 (.ZN( u2_u12_u3_n124 ) , .A1( u2_u12_u3_n96 ) , .A2( u2_u12_u3_n97 ) );
  NAND2_X1 u2_u12_u3_U58 (.A2( u2_u12_u3_n100 ) , .ZN( u2_u12_u3_n146 ) , .A1( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U59 (.A1( u2_u12_u3_n101 ) , .ZN( u2_u12_u3_n145 ) , .A2( u2_u12_u3_n99 ) );
  AOI221_X1 u2_u12_u3_U6 (.A( u2_u12_u3_n131 ) , .C2( u2_u12_u3_n132 ) , .C1( u2_u12_u3_n133 ) , .ZN( u2_u12_u3_n134 ) , .B1( u2_u12_u3_n143 ) , .B2( u2_u12_u3_n177 ) );
  NAND2_X1 u2_u12_u3_U60 (.A1( u2_u12_u3_n100 ) , .ZN( u2_u12_u3_n156 ) , .A2( u2_u12_u3_n99 ) );
  NAND2_X1 u2_u12_u3_U61 (.A2( u2_u12_u3_n101 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n148 ) );
  NAND2_X1 u2_u12_u3_U62 (.A1( u2_u12_u3_n100 ) , .A2( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n128 ) );
  NAND2_X1 u2_u12_u3_U63 (.A2( u2_u12_u3_n101 ) , .A1( u2_u12_u3_n102 ) , .ZN( u2_u12_u3_n152 ) );
  NAND2_X1 u2_u12_u3_U64 (.A2( u2_u12_u3_n101 ) , .ZN( u2_u12_u3_n114 ) , .A1( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U65 (.ZN( u2_u12_u3_n107 ) , .A1( u2_u12_u3_n97 ) , .A2( u2_u12_u3_n99 ) );
  NAND2_X1 u2_u12_u3_U66 (.A2( u2_u12_u3_n100 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n113 ) );
  NAND2_X1 u2_u12_u3_U67 (.A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n153 ) , .A2( u2_u12_u3_n97 ) );
  NAND2_X1 u2_u12_u3_U68 (.A2( u2_u12_u3_n103 ) , .A1( u2_u12_u3_n104 ) , .ZN( u2_u12_u3_n130 ) );
  NAND2_X1 u2_u12_u3_U69 (.A2( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n144 ) , .A1( u2_u12_u3_n96 ) );
  OAI22_X1 u2_u12_u3_U7 (.B2( u2_u12_u3_n147 ) , .A2( u2_u12_u3_n148 ) , .ZN( u2_u12_u3_n160 ) , .B1( u2_u12_u3_n165 ) , .A1( u2_u12_u3_n168 ) );
  NAND2_X1 u2_u12_u3_U70 (.A1( u2_u12_u3_n102 ) , .A2( u2_u12_u3_n103 ) , .ZN( u2_u12_u3_n108 ) );
  NOR2_X1 u2_u12_u3_U71 (.A2( u2_u12_X_19 ) , .A1( u2_u12_X_20 ) , .ZN( u2_u12_u3_n99 ) );
  NOR2_X1 u2_u12_u3_U72 (.A2( u2_u12_X_21 ) , .A1( u2_u12_X_24 ) , .ZN( u2_u12_u3_n103 ) );
  NOR2_X1 u2_u12_u3_U73 (.A2( u2_u12_X_24 ) , .A1( u2_u12_u3_n171 ) , .ZN( u2_u12_u3_n97 ) );
  NOR2_X1 u2_u12_u3_U74 (.A2( u2_u12_X_23 ) , .ZN( u2_u12_u3_n141 ) , .A1( u2_u12_u3_n166 ) );
  NOR2_X1 u2_u12_u3_U75 (.A2( u2_u12_X_19 ) , .A1( u2_u12_u3_n172 ) , .ZN( u2_u12_u3_n96 ) );
  NAND2_X1 u2_u12_u3_U76 (.A1( u2_u12_X_22 ) , .A2( u2_u12_X_23 ) , .ZN( u2_u12_u3_n154 ) );
  NAND2_X1 u2_u12_u3_U77 (.A1( u2_u12_X_23 ) , .ZN( u2_u12_u3_n149 ) , .A2( u2_u12_u3_n166 ) );
  NOR2_X1 u2_u12_u3_U78 (.A2( u2_u12_X_22 ) , .A1( u2_u12_X_23 ) , .ZN( u2_u12_u3_n121 ) );
  AND2_X1 u2_u12_u3_U79 (.A1( u2_u12_X_24 ) , .ZN( u2_u12_u3_n101 ) , .A2( u2_u12_u3_n171 ) );
  AND3_X1 u2_u12_u3_U8 (.A3( u2_u12_u3_n144 ) , .A2( u2_u12_u3_n145 ) , .A1( u2_u12_u3_n146 ) , .ZN( u2_u12_u3_n147 ) );
  AND2_X1 u2_u12_u3_U80 (.A1( u2_u12_X_19 ) , .ZN( u2_u12_u3_n102 ) , .A2( u2_u12_u3_n172 ) );
  AND2_X1 u2_u12_u3_U81 (.A1( u2_u12_X_21 ) , .A2( u2_u12_X_24 ) , .ZN( u2_u12_u3_n100 ) );
  AND2_X1 u2_u12_u3_U82 (.A2( u2_u12_X_19 ) , .A1( u2_u12_X_20 ) , .ZN( u2_u12_u3_n104 ) );
  INV_X1 u2_u12_u3_U83 (.A( u2_u12_X_22 ) , .ZN( u2_u12_u3_n166 ) );
  INV_X1 u2_u12_u3_U84 (.A( u2_u12_X_21 ) , .ZN( u2_u12_u3_n171 ) );
  INV_X1 u2_u12_u3_U85 (.A( u2_u12_X_20 ) , .ZN( u2_u12_u3_n172 ) );
  OR4_X1 u2_u12_u3_U86 (.ZN( u2_out12_10 ) , .A4( u2_u12_u3_n136 ) , .A3( u2_u12_u3_n137 ) , .A1( u2_u12_u3_n138 ) , .A2( u2_u12_u3_n139 ) );
  OAI222_X1 u2_u12_u3_U87 (.C1( u2_u12_u3_n128 ) , .ZN( u2_u12_u3_n137 ) , .B1( u2_u12_u3_n148 ) , .A2( u2_u12_u3_n150 ) , .B2( u2_u12_u3_n154 ) , .C2( u2_u12_u3_n164 ) , .A1( u2_u12_u3_n167 ) );
  OAI221_X1 u2_u12_u3_U88 (.A( u2_u12_u3_n134 ) , .B2( u2_u12_u3_n135 ) , .ZN( u2_u12_u3_n136 ) , .C1( u2_u12_u3_n149 ) , .B1( u2_u12_u3_n151 ) , .C2( u2_u12_u3_n183 ) );
  NAND4_X1 u2_u12_u3_U89 (.ZN( u2_out12_26 ) , .A4( u2_u12_u3_n109 ) , .A3( u2_u12_u3_n110 ) , .A2( u2_u12_u3_n111 ) , .A1( u2_u12_u3_n173 ) );
  INV_X1 u2_u12_u3_U9 (.A( u2_u12_u3_n143 ) , .ZN( u2_u12_u3_n168 ) );
  INV_X1 u2_u12_u3_U90 (.ZN( u2_u12_u3_n173 ) , .A( u2_u12_u3_n94 ) );
  OAI21_X1 u2_u12_u3_U91 (.ZN( u2_u12_u3_n111 ) , .B2( u2_u12_u3_n117 ) , .A( u2_u12_u3_n133 ) , .B1( u2_u12_u3_n176 ) );
  NAND4_X1 u2_u12_u3_U92 (.ZN( u2_out12_20 ) , .A4( u2_u12_u3_n122 ) , .A3( u2_u12_u3_n123 ) , .A1( u2_u12_u3_n175 ) , .A2( u2_u12_u3_n180 ) );
  INV_X1 u2_u12_u3_U93 (.A( u2_u12_u3_n126 ) , .ZN( u2_u12_u3_n180 ) );
  INV_X1 u2_u12_u3_U94 (.A( u2_u12_u3_n112 ) , .ZN( u2_u12_u3_n175 ) );
  NAND4_X1 u2_u12_u3_U95 (.ZN( u2_out12_1 ) , .A4( u2_u12_u3_n161 ) , .A3( u2_u12_u3_n162 ) , .A2( u2_u12_u3_n163 ) , .A1( u2_u12_u3_n185 ) );
  NAND2_X1 u2_u12_u3_U96 (.ZN( u2_u12_u3_n163 ) , .A2( u2_u12_u3_n170 ) , .A1( u2_u12_u3_n176 ) );
  AOI22_X1 u2_u12_u3_U97 (.B2( u2_u12_u3_n140 ) , .B1( u2_u12_u3_n141 ) , .A2( u2_u12_u3_n142 ) , .ZN( u2_u12_u3_n162 ) , .A1( u2_u12_u3_n177 ) );
  NAND3_X1 u2_u12_u3_U98 (.A1( u2_u12_u3_n114 ) , .ZN( u2_u12_u3_n115 ) , .A2( u2_u12_u3_n145 ) , .A3( u2_u12_u3_n153 ) );
  NAND3_X1 u2_u12_u3_U99 (.ZN( u2_u12_u3_n129 ) , .A2( u2_u12_u3_n144 ) , .A1( u2_u12_u3_n153 ) , .A3( u2_u12_u3_n182 ) );
  XOR2_X1 u2_u13_U1 (.B( u2_K14_9 ) , .A( u2_R12_6 ) , .Z( u2_u13_X_9 ) );
  XOR2_X1 u2_u13_U10 (.B( u2_K14_45 ) , .A( u2_R12_30 ) , .Z( u2_u13_X_45 ) );
  XOR2_X1 u2_u13_U11 (.B( u2_K14_44 ) , .A( u2_R12_29 ) , .Z( u2_u13_X_44 ) );
  XOR2_X1 u2_u13_U12 (.B( u2_K14_43 ) , .A( u2_R12_28 ) , .Z( u2_u13_X_43 ) );
  XOR2_X1 u2_u13_U13 (.B( u2_K14_42 ) , .A( u2_R12_29 ) , .Z( u2_u13_X_42 ) );
  XOR2_X1 u2_u13_U14 (.B( u2_K14_41 ) , .A( u2_R12_28 ) , .Z( u2_u13_X_41 ) );
  XOR2_X1 u2_u13_U15 (.B( u2_K14_40 ) , .A( u2_R12_27 ) , .Z( u2_u13_X_40 ) );
  XOR2_X1 u2_u13_U16 (.B( u2_K14_3 ) , .A( u2_R12_2 ) , .Z( u2_u13_X_3 ) );
  XOR2_X1 u2_u13_U17 (.B( u2_K14_39 ) , .A( u2_R12_26 ) , .Z( u2_u13_X_39 ) );
  XOR2_X1 u2_u13_U19 (.B( u2_K14_37 ) , .A( u2_R12_24 ) , .Z( u2_u13_X_37 ) );
  XOR2_X1 u2_u13_U2 (.B( u2_K14_8 ) , .A( u2_R12_5 ) , .Z( u2_u13_X_8 ) );
  XOR2_X1 u2_u13_U21 (.B( u2_K14_35 ) , .A( u2_R12_24 ) , .Z( u2_u13_X_35 ) );
  XOR2_X1 u2_u13_U22 (.B( u2_K14_34 ) , .A( u2_R12_23 ) , .Z( u2_u13_X_34 ) );
  XOR2_X1 u2_u13_U27 (.B( u2_K14_2 ) , .A( u2_R12_1 ) , .Z( u2_u13_X_2 ) );
  XOR2_X1 u2_u13_U29 (.B( u2_K14_28 ) , .A( u2_R12_19 ) , .Z( u2_u13_X_28 ) );
  XOR2_X1 u2_u13_U3 (.B( u2_K14_7 ) , .A( u2_R12_4 ) , .Z( u2_u13_X_7 ) );
  XOR2_X1 u2_u13_U30 (.B( u2_K14_27 ) , .A( u2_R12_18 ) , .Z( u2_u13_X_27 ) );
  XOR2_X1 u2_u13_U31 (.B( u2_K14_26 ) , .A( u2_R12_17 ) , .Z( u2_u13_X_26 ) );
  XOR2_X1 u2_u13_U32 (.B( u2_K14_25 ) , .A( u2_R12_16 ) , .Z( u2_u13_X_25 ) );
  XOR2_X1 u2_u13_U33 (.B( u2_K14_24 ) , .A( u2_R12_17 ) , .Z( u2_u13_X_24 ) );
  XOR2_X1 u2_u13_U34 (.B( u2_K14_23 ) , .A( u2_R12_16 ) , .Z( u2_u13_X_23 ) );
  XOR2_X1 u2_u13_U35 (.B( u2_K14_22 ) , .A( u2_R12_15 ) , .Z( u2_u13_X_22 ) );
  XOR2_X1 u2_u13_U36 (.B( u2_K14_21 ) , .A( u2_R12_14 ) , .Z( u2_u13_X_21 ) );
  XOR2_X1 u2_u13_U37 (.B( u2_K14_20 ) , .A( u2_R12_13 ) , .Z( u2_u13_X_20 ) );
  XOR2_X1 u2_u13_U38 (.B( u2_K14_1 ) , .A( u2_R12_32 ) , .Z( u2_u13_X_1 ) );
  XOR2_X1 u2_u13_U39 (.B( u2_K14_19 ) , .A( u2_R12_12 ) , .Z( u2_u13_X_19 ) );
  XOR2_X1 u2_u13_U4 (.B( u2_K14_6 ) , .A( u2_R12_5 ) , .Z( u2_u13_X_6 ) );
  XOR2_X1 u2_u13_U40 (.B( u2_K14_18 ) , .A( u2_R12_13 ) , .Z( u2_u13_X_18 ) );
  XOR2_X1 u2_u13_U41 (.B( u2_K14_17 ) , .A( u2_R12_12 ) , .Z( u2_u13_X_17 ) );
  XOR2_X1 u2_u13_U42 (.B( u2_K14_16 ) , .A( u2_R12_11 ) , .Z( u2_u13_X_16 ) );
  XOR2_X1 u2_u13_U43 (.B( u2_K14_15 ) , .A( u2_R12_10 ) , .Z( u2_u13_X_15 ) );
  XOR2_X1 u2_u13_U44 (.B( u2_K14_14 ) , .A( u2_R12_9 ) , .Z( u2_u13_X_14 ) );
  XOR2_X1 u2_u13_U45 (.B( u2_K14_13 ) , .A( u2_R12_8 ) , .Z( u2_u13_X_13 ) );
  XOR2_X1 u2_u13_U46 (.B( u2_K14_12 ) , .A( u2_R12_9 ) , .Z( u2_u13_X_12 ) );
  XOR2_X1 u2_u13_U47 (.B( u2_K14_11 ) , .A( u2_R12_8 ) , .Z( u2_u13_X_11 ) );
  XOR2_X1 u2_u13_U48 (.B( u2_K14_10 ) , .A( u2_R12_7 ) , .Z( u2_u13_X_10 ) );
  XOR2_X1 u2_u13_U5 (.B( u2_K14_5 ) , .A( u2_R12_4 ) , .Z( u2_u13_X_5 ) );
  XOR2_X1 u2_u13_U6 (.B( u2_K14_4 ) , .A( u2_R12_3 ) , .Z( u2_u13_X_4 ) );
  XOR2_X1 u2_u13_U7 (.B( u2_K14_48 ) , .A( u2_R12_1 ) , .Z( u2_u13_X_48 ) );
  XOR2_X1 u2_u13_U8 (.B( u2_K14_47 ) , .A( u2_R12_32 ) , .Z( u2_u13_X_47 ) );
  XOR2_X1 u2_u13_U9 (.B( u2_K14_46 ) , .A( u2_R12_31 ) , .Z( u2_u13_X_46 ) );
  AND3_X1 u2_u13_u0_U10 (.A2( u2_u13_u0_n112 ) , .ZN( u2_u13_u0_n127 ) , .A3( u2_u13_u0_n130 ) , .A1( u2_u13_u0_n148 ) );
  NAND2_X1 u2_u13_u0_U11 (.ZN( u2_u13_u0_n113 ) , .A1( u2_u13_u0_n139 ) , .A2( u2_u13_u0_n149 ) );
  AND2_X1 u2_u13_u0_U12 (.ZN( u2_u13_u0_n107 ) , .A1( u2_u13_u0_n130 ) , .A2( u2_u13_u0_n140 ) );
  AND2_X1 u2_u13_u0_U13 (.A2( u2_u13_u0_n129 ) , .A1( u2_u13_u0_n130 ) , .ZN( u2_u13_u0_n151 ) );
  AND2_X1 u2_u13_u0_U14 (.A1( u2_u13_u0_n108 ) , .A2( u2_u13_u0_n125 ) , .ZN( u2_u13_u0_n145 ) );
  INV_X1 u2_u13_u0_U15 (.A( u2_u13_u0_n143 ) , .ZN( u2_u13_u0_n173 ) );
  NOR2_X1 u2_u13_u0_U16 (.A2( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n147 ) , .A1( u2_u13_u0_n160 ) );
  INV_X1 u2_u13_u0_U17 (.ZN( u2_u13_u0_n172 ) , .A( u2_u13_u0_n88 ) );
  OAI222_X1 u2_u13_u0_U18 (.C1( u2_u13_u0_n108 ) , .A1( u2_u13_u0_n125 ) , .B2( u2_u13_u0_n128 ) , .B1( u2_u13_u0_n144 ) , .A2( u2_u13_u0_n158 ) , .C2( u2_u13_u0_n161 ) , .ZN( u2_u13_u0_n88 ) );
  NOR2_X1 u2_u13_u0_U19 (.A1( u2_u13_u0_n163 ) , .A2( u2_u13_u0_n164 ) , .ZN( u2_u13_u0_n95 ) );
  AOI21_X1 u2_u13_u0_U20 (.B1( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n132 ) , .A( u2_u13_u0_n165 ) , .B2( u2_u13_u0_n93 ) );
  INV_X1 u2_u13_u0_U21 (.A( u2_u13_u0_n142 ) , .ZN( u2_u13_u0_n165 ) );
  OAI221_X1 u2_u13_u0_U22 (.C1( u2_u13_u0_n121 ) , .ZN( u2_u13_u0_n122 ) , .B2( u2_u13_u0_n127 ) , .A( u2_u13_u0_n143 ) , .B1( u2_u13_u0_n144 ) , .C2( u2_u13_u0_n147 ) );
  OAI22_X1 u2_u13_u0_U23 (.B1( u2_u13_u0_n125 ) , .ZN( u2_u13_u0_n126 ) , .A1( u2_u13_u0_n138 ) , .A2( u2_u13_u0_n146 ) , .B2( u2_u13_u0_n147 ) );
  OAI22_X1 u2_u13_u0_U24 (.B1( u2_u13_u0_n131 ) , .A1( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n147 ) , .A2( u2_u13_u0_n90 ) , .ZN( u2_u13_u0_n91 ) );
  AND3_X1 u2_u13_u0_U25 (.A3( u2_u13_u0_n121 ) , .A2( u2_u13_u0_n125 ) , .A1( u2_u13_u0_n148 ) , .ZN( u2_u13_u0_n90 ) );
  INV_X1 u2_u13_u0_U26 (.A( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n161 ) );
  NOR2_X1 u2_u13_u0_U27 (.A1( u2_u13_u0_n120 ) , .ZN( u2_u13_u0_n143 ) , .A2( u2_u13_u0_n167 ) );
  OAI221_X1 u2_u13_u0_U28 (.C1( u2_u13_u0_n112 ) , .ZN( u2_u13_u0_n120 ) , .B1( u2_u13_u0_n138 ) , .B2( u2_u13_u0_n141 ) , .C2( u2_u13_u0_n147 ) , .A( u2_u13_u0_n172 ) );
  AOI211_X1 u2_u13_u0_U29 (.B( u2_u13_u0_n115 ) , .A( u2_u13_u0_n116 ) , .C2( u2_u13_u0_n117 ) , .C1( u2_u13_u0_n118 ) , .ZN( u2_u13_u0_n119 ) );
  INV_X1 u2_u13_u0_U3 (.A( u2_u13_u0_n113 ) , .ZN( u2_u13_u0_n166 ) );
  AOI22_X1 u2_u13_u0_U30 (.B2( u2_u13_u0_n109 ) , .A2( u2_u13_u0_n110 ) , .ZN( u2_u13_u0_n111 ) , .B1( u2_u13_u0_n118 ) , .A1( u2_u13_u0_n160 ) );
  INV_X1 u2_u13_u0_U31 (.A( u2_u13_u0_n118 ) , .ZN( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U32 (.ZN( u2_u13_u0_n104 ) , .B1( u2_u13_u0_n107 ) , .B2( u2_u13_u0_n141 ) , .A( u2_u13_u0_n144 ) );
  AOI21_X1 u2_u13_u0_U33 (.B1( u2_u13_u0_n127 ) , .B2( u2_u13_u0_n129 ) , .A( u2_u13_u0_n138 ) , .ZN( u2_u13_u0_n96 ) );
  AOI21_X1 u2_u13_u0_U34 (.ZN( u2_u13_u0_n116 ) , .B2( u2_u13_u0_n142 ) , .A( u2_u13_u0_n144 ) , .B1( u2_u13_u0_n166 ) );
  NAND2_X1 u2_u13_u0_U35 (.A1( u2_u13_u0_n100 ) , .A2( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n125 ) );
  NAND2_X1 u2_u13_u0_U36 (.A1( u2_u13_u0_n101 ) , .A2( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n150 ) );
  INV_X1 u2_u13_u0_U37 (.A( u2_u13_u0_n138 ) , .ZN( u2_u13_u0_n160 ) );
  NAND2_X1 u2_u13_u0_U38 (.A1( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n128 ) , .A2( u2_u13_u0_n95 ) );
  NAND2_X1 u2_u13_u0_U39 (.A1( u2_u13_u0_n100 ) , .ZN( u2_u13_u0_n129 ) , .A2( u2_u13_u0_n95 ) );
  AOI21_X1 u2_u13_u0_U4 (.B1( u2_u13_u0_n114 ) , .ZN( u2_u13_u0_n115 ) , .B2( u2_u13_u0_n129 ) , .A( u2_u13_u0_n161 ) );
  NAND2_X1 u2_u13_u0_U40 (.A2( u2_u13_u0_n100 ) , .ZN( u2_u13_u0_n131 ) , .A1( u2_u13_u0_n92 ) );
  NAND2_X1 u2_u13_u0_U41 (.A2( u2_u13_u0_n100 ) , .A1( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n139 ) );
  NAND2_X1 u2_u13_u0_U42 (.ZN( u2_u13_u0_n148 ) , .A1( u2_u13_u0_n93 ) , .A2( u2_u13_u0_n95 ) );
  NAND2_X1 u2_u13_u0_U43 (.A2( u2_u13_u0_n102 ) , .A1( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n149 ) );
  NAND2_X1 u2_u13_u0_U44 (.A2( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n114 ) , .A1( u2_u13_u0_n92 ) );
  NAND2_X1 u2_u13_u0_U45 (.A2( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n121 ) , .A1( u2_u13_u0_n93 ) );
  NAND2_X1 u2_u13_u0_U46 (.ZN( u2_u13_u0_n112 ) , .A2( u2_u13_u0_n92 ) , .A1( u2_u13_u0_n93 ) );
  OR3_X1 u2_u13_u0_U47 (.A3( u2_u13_u0_n152 ) , .A2( u2_u13_u0_n153 ) , .A1( u2_u13_u0_n154 ) , .ZN( u2_u13_u0_n155 ) );
  AOI21_X1 u2_u13_u0_U48 (.B2( u2_u13_u0_n150 ) , .B1( u2_u13_u0_n151 ) , .ZN( u2_u13_u0_n152 ) , .A( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U49 (.A( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n145 ) , .B1( u2_u13_u0_n146 ) , .ZN( u2_u13_u0_n154 ) );
  AOI21_X1 u2_u13_u0_U5 (.B2( u2_u13_u0_n131 ) , .ZN( u2_u13_u0_n134 ) , .B1( u2_u13_u0_n151 ) , .A( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U50 (.A( u2_u13_u0_n147 ) , .B2( u2_u13_u0_n148 ) , .B1( u2_u13_u0_n149 ) , .ZN( u2_u13_u0_n153 ) );
  INV_X1 u2_u13_u0_U51 (.ZN( u2_u13_u0_n171 ) , .A( u2_u13_u0_n99 ) );
  OAI211_X1 u2_u13_u0_U52 (.C2( u2_u13_u0_n140 ) , .C1( u2_u13_u0_n161 ) , .A( u2_u13_u0_n169 ) , .B( u2_u13_u0_n98 ) , .ZN( u2_u13_u0_n99 ) );
  INV_X1 u2_u13_u0_U53 (.ZN( u2_u13_u0_n169 ) , .A( u2_u13_u0_n91 ) );
  AOI211_X1 u2_u13_u0_U54 (.C1( u2_u13_u0_n118 ) , .A( u2_u13_u0_n123 ) , .B( u2_u13_u0_n96 ) , .C2( u2_u13_u0_n97 ) , .ZN( u2_u13_u0_n98 ) );
  NOR2_X1 u2_u13_u0_U55 (.A2( u2_u13_X_6 ) , .ZN( u2_u13_u0_n100 ) , .A1( u2_u13_u0_n162 ) );
  NOR2_X1 u2_u13_u0_U56 (.A2( u2_u13_X_4 ) , .A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n118 ) );
  NOR2_X1 u2_u13_u0_U57 (.A2( u2_u13_X_2 ) , .ZN( u2_u13_u0_n103 ) , .A1( u2_u13_u0_n164 ) );
  NOR2_X1 u2_u13_u0_U58 (.A2( u2_u13_X_1 ) , .A1( u2_u13_X_2 ) , .ZN( u2_u13_u0_n92 ) );
  NOR2_X1 u2_u13_u0_U59 (.A2( u2_u13_X_1 ) , .ZN( u2_u13_u0_n101 ) , .A1( u2_u13_u0_n163 ) );
  NOR2_X1 u2_u13_u0_U6 (.A1( u2_u13_u0_n108 ) , .ZN( u2_u13_u0_n123 ) , .A2( u2_u13_u0_n158 ) );
  NAND2_X1 u2_u13_u0_U60 (.A2( u2_u13_X_4 ) , .A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n144 ) );
  NOR2_X1 u2_u13_u0_U61 (.A2( u2_u13_X_5 ) , .ZN( u2_u13_u0_n136 ) , .A1( u2_u13_u0_n159 ) );
  NAND2_X1 u2_u13_u0_U62 (.A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n138 ) , .A2( u2_u13_u0_n159 ) );
  NOR2_X1 u2_u13_u0_U63 (.A2( u2_u13_X_3 ) , .A1( u2_u13_X_6 ) , .ZN( u2_u13_u0_n94 ) );
  AND2_X1 u2_u13_u0_U64 (.A2( u2_u13_X_3 ) , .A1( u2_u13_X_6 ) , .ZN( u2_u13_u0_n102 ) );
  AND2_X1 u2_u13_u0_U65 (.A1( u2_u13_X_6 ) , .A2( u2_u13_u0_n162 ) , .ZN( u2_u13_u0_n93 ) );
  INV_X1 u2_u13_u0_U66 (.A( u2_u13_X_4 ) , .ZN( u2_u13_u0_n159 ) );
  INV_X1 u2_u13_u0_U67 (.A( u2_u13_X_1 ) , .ZN( u2_u13_u0_n164 ) );
  INV_X1 u2_u13_u0_U68 (.A( u2_u13_X_2 ) , .ZN( u2_u13_u0_n163 ) );
  INV_X1 u2_u13_u0_U69 (.A( u2_u13_X_3 ) , .ZN( u2_u13_u0_n162 ) );
  OAI21_X1 u2_u13_u0_U7 (.B1( u2_u13_u0_n150 ) , .B2( u2_u13_u0_n158 ) , .A( u2_u13_u0_n172 ) , .ZN( u2_u13_u0_n89 ) );
  INV_X1 u2_u13_u0_U70 (.A( u2_u13_u0_n126 ) , .ZN( u2_u13_u0_n168 ) );
  AOI211_X1 u2_u13_u0_U71 (.B( u2_u13_u0_n133 ) , .A( u2_u13_u0_n134 ) , .C2( u2_u13_u0_n135 ) , .C1( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n137 ) );
  INV_X1 u2_u13_u0_U72 (.ZN( u2_u13_u0_n174 ) , .A( u2_u13_u0_n89 ) );
  AOI211_X1 u2_u13_u0_U73 (.B( u2_u13_u0_n104 ) , .A( u2_u13_u0_n105 ) , .ZN( u2_u13_u0_n106 ) , .C2( u2_u13_u0_n113 ) , .C1( u2_u13_u0_n160 ) );
  OR4_X1 u2_u13_u0_U74 (.ZN( u2_out13_17 ) , .A4( u2_u13_u0_n122 ) , .A2( u2_u13_u0_n123 ) , .A1( u2_u13_u0_n124 ) , .A3( u2_u13_u0_n170 ) );
  AOI21_X1 u2_u13_u0_U75 (.B2( u2_u13_u0_n107 ) , .ZN( u2_u13_u0_n124 ) , .B1( u2_u13_u0_n128 ) , .A( u2_u13_u0_n161 ) );
  INV_X1 u2_u13_u0_U76 (.A( u2_u13_u0_n111 ) , .ZN( u2_u13_u0_n170 ) );
  OR4_X1 u2_u13_u0_U77 (.ZN( u2_out13_31 ) , .A4( u2_u13_u0_n155 ) , .A2( u2_u13_u0_n156 ) , .A1( u2_u13_u0_n157 ) , .A3( u2_u13_u0_n173 ) );
  AOI21_X1 u2_u13_u0_U78 (.A( u2_u13_u0_n138 ) , .B2( u2_u13_u0_n139 ) , .B1( u2_u13_u0_n140 ) , .ZN( u2_u13_u0_n157 ) );
  AOI21_X1 u2_u13_u0_U79 (.B2( u2_u13_u0_n141 ) , .B1( u2_u13_u0_n142 ) , .ZN( u2_u13_u0_n156 ) , .A( u2_u13_u0_n161 ) );
  AND2_X1 u2_u13_u0_U8 (.A1( u2_u13_u0_n114 ) , .A2( u2_u13_u0_n121 ) , .ZN( u2_u13_u0_n146 ) );
  AOI21_X1 u2_u13_u0_U80 (.B1( u2_u13_u0_n132 ) , .ZN( u2_u13_u0_n133 ) , .A( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n166 ) );
  OAI22_X1 u2_u13_u0_U81 (.ZN( u2_u13_u0_n105 ) , .A2( u2_u13_u0_n132 ) , .B1( u2_u13_u0_n146 ) , .A1( u2_u13_u0_n147 ) , .B2( u2_u13_u0_n161 ) );
  NAND2_X1 u2_u13_u0_U82 (.ZN( u2_u13_u0_n110 ) , .A2( u2_u13_u0_n132 ) , .A1( u2_u13_u0_n145 ) );
  INV_X1 u2_u13_u0_U83 (.A( u2_u13_u0_n119 ) , .ZN( u2_u13_u0_n167 ) );
  NAND2_X1 u2_u13_u0_U84 (.A2( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n140 ) , .A1( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U85 (.A1( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n130 ) , .A2( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U86 (.ZN( u2_u13_u0_n108 ) , .A1( u2_u13_u0_n92 ) , .A2( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U87 (.ZN( u2_u13_u0_n142 ) , .A1( u2_u13_u0_n94 ) , .A2( u2_u13_u0_n95 ) );
  NAND3_X1 u2_u13_u0_U88 (.ZN( u2_out13_23 ) , .A3( u2_u13_u0_n137 ) , .A1( u2_u13_u0_n168 ) , .A2( u2_u13_u0_n171 ) );
  NAND3_X1 u2_u13_u0_U89 (.A3( u2_u13_u0_n127 ) , .A2( u2_u13_u0_n128 ) , .ZN( u2_u13_u0_n135 ) , .A1( u2_u13_u0_n150 ) );
  AND2_X1 u2_u13_u0_U9 (.A1( u2_u13_u0_n131 ) , .ZN( u2_u13_u0_n141 ) , .A2( u2_u13_u0_n150 ) );
  NAND3_X1 u2_u13_u0_U90 (.ZN( u2_u13_u0_n117 ) , .A3( u2_u13_u0_n132 ) , .A2( u2_u13_u0_n139 ) , .A1( u2_u13_u0_n148 ) );
  NAND3_X1 u2_u13_u0_U91 (.ZN( u2_u13_u0_n109 ) , .A2( u2_u13_u0_n114 ) , .A3( u2_u13_u0_n140 ) , .A1( u2_u13_u0_n149 ) );
  NAND3_X1 u2_u13_u0_U92 (.ZN( u2_out13_9 ) , .A3( u2_u13_u0_n106 ) , .A2( u2_u13_u0_n171 ) , .A1( u2_u13_u0_n174 ) );
  NAND3_X1 u2_u13_u0_U93 (.A2( u2_u13_u0_n128 ) , .A1( u2_u13_u0_n132 ) , .A3( u2_u13_u0_n146 ) , .ZN( u2_u13_u0_n97 ) );
  AOI21_X1 u2_u13_u1_U10 (.B2( u2_u13_u1_n155 ) , .B1( u2_u13_u1_n156 ) , .ZN( u2_u13_u1_n157 ) , .A( u2_u13_u1_n174 ) );
  NAND3_X1 u2_u13_u1_U100 (.ZN( u2_u13_u1_n113 ) , .A1( u2_u13_u1_n120 ) , .A3( u2_u13_u1_n133 ) , .A2( u2_u13_u1_n155 ) );
  NAND2_X1 u2_u13_u1_U11 (.ZN( u2_u13_u1_n140 ) , .A2( u2_u13_u1_n150 ) , .A1( u2_u13_u1_n155 ) );
  NAND2_X1 u2_u13_u1_U12 (.A1( u2_u13_u1_n131 ) , .ZN( u2_u13_u1_n147 ) , .A2( u2_u13_u1_n153 ) );
  INV_X1 u2_u13_u1_U13 (.A( u2_u13_u1_n139 ) , .ZN( u2_u13_u1_n174 ) );
  OR4_X1 u2_u13_u1_U14 (.A4( u2_u13_u1_n106 ) , .A3( u2_u13_u1_n107 ) , .ZN( u2_u13_u1_n108 ) , .A1( u2_u13_u1_n117 ) , .A2( u2_u13_u1_n184 ) );
  AOI21_X1 u2_u13_u1_U15 (.ZN( u2_u13_u1_n106 ) , .A( u2_u13_u1_n112 ) , .B1( u2_u13_u1_n154 ) , .B2( u2_u13_u1_n156 ) );
  AOI21_X1 u2_u13_u1_U16 (.ZN( u2_u13_u1_n107 ) , .B1( u2_u13_u1_n134 ) , .B2( u2_u13_u1_n149 ) , .A( u2_u13_u1_n174 ) );
  INV_X1 u2_u13_u1_U17 (.A( u2_u13_u1_n101 ) , .ZN( u2_u13_u1_n184 ) );
  INV_X1 u2_u13_u1_U18 (.A( u2_u13_u1_n112 ) , .ZN( u2_u13_u1_n171 ) );
  NAND2_X1 u2_u13_u1_U19 (.ZN( u2_u13_u1_n141 ) , .A1( u2_u13_u1_n153 ) , .A2( u2_u13_u1_n156 ) );
  AND2_X1 u2_u13_u1_U20 (.A1( u2_u13_u1_n123 ) , .ZN( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n161 ) );
  NAND2_X1 u2_u13_u1_U21 (.A2( u2_u13_u1_n115 ) , .A1( u2_u13_u1_n116 ) , .ZN( u2_u13_u1_n148 ) );
  NAND2_X1 u2_u13_u1_U22 (.A2( u2_u13_u1_n133 ) , .A1( u2_u13_u1_n135 ) , .ZN( u2_u13_u1_n159 ) );
  NAND2_X1 u2_u13_u1_U23 (.A2( u2_u13_u1_n115 ) , .A1( u2_u13_u1_n120 ) , .ZN( u2_u13_u1_n132 ) );
  INV_X1 u2_u13_u1_U24 (.A( u2_u13_u1_n154 ) , .ZN( u2_u13_u1_n178 ) );
  AOI22_X1 u2_u13_u1_U25 (.B2( u2_u13_u1_n113 ) , .A2( u2_u13_u1_n114 ) , .ZN( u2_u13_u1_n125 ) , .A1( u2_u13_u1_n171 ) , .B1( u2_u13_u1_n173 ) );
  NAND2_X1 u2_u13_u1_U26 (.ZN( u2_u13_u1_n114 ) , .A1( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n156 ) );
  INV_X1 u2_u13_u1_U27 (.A( u2_u13_u1_n151 ) , .ZN( u2_u13_u1_n183 ) );
  AND2_X1 u2_u13_u1_U28 (.A1( u2_u13_u1_n129 ) , .A2( u2_u13_u1_n133 ) , .ZN( u2_u13_u1_n149 ) );
  INV_X1 u2_u13_u1_U29 (.A( u2_u13_u1_n131 ) , .ZN( u2_u13_u1_n180 ) );
  INV_X1 u2_u13_u1_U3 (.A( u2_u13_u1_n159 ) , .ZN( u2_u13_u1_n182 ) );
  OAI221_X1 u2_u13_u1_U30 (.A( u2_u13_u1_n119 ) , .C2( u2_u13_u1_n129 ) , .ZN( u2_u13_u1_n138 ) , .B2( u2_u13_u1_n152 ) , .C1( u2_u13_u1_n174 ) , .B1( u2_u13_u1_n187 ) );
  INV_X1 u2_u13_u1_U31 (.A( u2_u13_u1_n148 ) , .ZN( u2_u13_u1_n187 ) );
  AOI211_X1 u2_u13_u1_U32 (.B( u2_u13_u1_n117 ) , .A( u2_u13_u1_n118 ) , .ZN( u2_u13_u1_n119 ) , .C2( u2_u13_u1_n146 ) , .C1( u2_u13_u1_n159 ) );
  NOR2_X1 u2_u13_u1_U33 (.A1( u2_u13_u1_n168 ) , .A2( u2_u13_u1_n176 ) , .ZN( u2_u13_u1_n98 ) );
  AOI211_X1 u2_u13_u1_U34 (.B( u2_u13_u1_n162 ) , .A( u2_u13_u1_n163 ) , .C2( u2_u13_u1_n164 ) , .ZN( u2_u13_u1_n165 ) , .C1( u2_u13_u1_n171 ) );
  AOI21_X1 u2_u13_u1_U35 (.A( u2_u13_u1_n160 ) , .B2( u2_u13_u1_n161 ) , .ZN( u2_u13_u1_n162 ) , .B1( u2_u13_u1_n182 ) );
  OR2_X1 u2_u13_u1_U36 (.A2( u2_u13_u1_n157 ) , .A1( u2_u13_u1_n158 ) , .ZN( u2_u13_u1_n163 ) );
  OAI21_X1 u2_u13_u1_U37 (.B2( u2_u13_u1_n123 ) , .ZN( u2_u13_u1_n145 ) , .B1( u2_u13_u1_n160 ) , .A( u2_u13_u1_n185 ) );
  INV_X1 u2_u13_u1_U38 (.A( u2_u13_u1_n122 ) , .ZN( u2_u13_u1_n185 ) );
  AOI21_X1 u2_u13_u1_U39 (.B2( u2_u13_u1_n120 ) , .B1( u2_u13_u1_n121 ) , .ZN( u2_u13_u1_n122 ) , .A( u2_u13_u1_n128 ) );
  AOI221_X1 u2_u13_u1_U4 (.A( u2_u13_u1_n138 ) , .C2( u2_u13_u1_n139 ) , .C1( u2_u13_u1_n140 ) , .B2( u2_u13_u1_n141 ) , .ZN( u2_u13_u1_n142 ) , .B1( u2_u13_u1_n175 ) );
  NAND2_X1 u2_u13_u1_U40 (.A1( u2_u13_u1_n128 ) , .ZN( u2_u13_u1_n146 ) , .A2( u2_u13_u1_n160 ) );
  NAND2_X1 u2_u13_u1_U41 (.A2( u2_u13_u1_n112 ) , .ZN( u2_u13_u1_n139 ) , .A1( u2_u13_u1_n152 ) );
  NAND2_X1 u2_u13_u1_U42 (.A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n156 ) , .A2( u2_u13_u1_n99 ) );
  AOI221_X1 u2_u13_u1_U43 (.B1( u2_u13_u1_n140 ) , .ZN( u2_u13_u1_n167 ) , .B2( u2_u13_u1_n172 ) , .C2( u2_u13_u1_n175 ) , .C1( u2_u13_u1_n178 ) , .A( u2_u13_u1_n188 ) );
  INV_X1 u2_u13_u1_U44 (.ZN( u2_u13_u1_n188 ) , .A( u2_u13_u1_n97 ) );
  AOI211_X1 u2_u13_u1_U45 (.A( u2_u13_u1_n118 ) , .C1( u2_u13_u1_n132 ) , .C2( u2_u13_u1_n139 ) , .B( u2_u13_u1_n96 ) , .ZN( u2_u13_u1_n97 ) );
  AOI21_X1 u2_u13_u1_U46 (.B2( u2_u13_u1_n121 ) , .B1( u2_u13_u1_n135 ) , .A( u2_u13_u1_n152 ) , .ZN( u2_u13_u1_n96 ) );
  NOR2_X1 u2_u13_u1_U47 (.ZN( u2_u13_u1_n117 ) , .A1( u2_u13_u1_n121 ) , .A2( u2_u13_u1_n160 ) );
  AOI21_X1 u2_u13_u1_U48 (.A( u2_u13_u1_n128 ) , .B2( u2_u13_u1_n129 ) , .ZN( u2_u13_u1_n130 ) , .B1( u2_u13_u1_n150 ) );
  NAND2_X1 u2_u13_u1_U49 (.ZN( u2_u13_u1_n112 ) , .A1( u2_u13_u1_n169 ) , .A2( u2_u13_u1_n170 ) );
  AOI211_X1 u2_u13_u1_U5 (.ZN( u2_u13_u1_n124 ) , .A( u2_u13_u1_n138 ) , .C2( u2_u13_u1_n139 ) , .B( u2_u13_u1_n145 ) , .C1( u2_u13_u1_n147 ) );
  NAND2_X1 u2_u13_u1_U50 (.ZN( u2_u13_u1_n129 ) , .A2( u2_u13_u1_n95 ) , .A1( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U51 (.A1( u2_u13_u1_n102 ) , .ZN( u2_u13_u1_n154 ) , .A2( u2_u13_u1_n99 ) );
  NAND2_X1 u2_u13_u1_U52 (.A2( u2_u13_u1_n100 ) , .ZN( u2_u13_u1_n135 ) , .A1( u2_u13_u1_n99 ) );
  AOI21_X1 u2_u13_u1_U53 (.A( u2_u13_u1_n152 ) , .B2( u2_u13_u1_n153 ) , .B1( u2_u13_u1_n154 ) , .ZN( u2_u13_u1_n158 ) );
  INV_X1 u2_u13_u1_U54 (.A( u2_u13_u1_n160 ) , .ZN( u2_u13_u1_n175 ) );
  NAND2_X1 u2_u13_u1_U55 (.A1( u2_u13_u1_n100 ) , .ZN( u2_u13_u1_n116 ) , .A2( u2_u13_u1_n95 ) );
  NAND2_X1 u2_u13_u1_U56 (.A1( u2_u13_u1_n102 ) , .ZN( u2_u13_u1_n131 ) , .A2( u2_u13_u1_n95 ) );
  NAND2_X1 u2_u13_u1_U57 (.A2( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n121 ) , .A1( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U58 (.A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n153 ) , .A2( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U59 (.A2( u2_u13_u1_n104 ) , .A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n133 ) );
  AOI22_X1 u2_u13_u1_U6 (.B2( u2_u13_u1_n136 ) , .A2( u2_u13_u1_n137 ) , .ZN( u2_u13_u1_n143 ) , .A1( u2_u13_u1_n171 ) , .B1( u2_u13_u1_n173 ) );
  NAND2_X1 u2_u13_u1_U60 (.ZN( u2_u13_u1_n150 ) , .A2( u2_u13_u1_n98 ) , .A1( u2_u13_u1_n99 ) );
  NAND2_X1 u2_u13_u1_U61 (.A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n155 ) , .A2( u2_u13_u1_n95 ) );
  OAI21_X1 u2_u13_u1_U62 (.ZN( u2_u13_u1_n109 ) , .B1( u2_u13_u1_n129 ) , .B2( u2_u13_u1_n160 ) , .A( u2_u13_u1_n167 ) );
  NAND2_X1 u2_u13_u1_U63 (.A2( u2_u13_u1_n100 ) , .A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n120 ) );
  NAND2_X1 u2_u13_u1_U64 (.A1( u2_u13_u1_n102 ) , .A2( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n115 ) );
  NAND2_X1 u2_u13_u1_U65 (.A2( u2_u13_u1_n100 ) , .A1( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n151 ) );
  NAND2_X1 u2_u13_u1_U66 (.A2( u2_u13_u1_n103 ) , .A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n161 ) );
  INV_X1 u2_u13_u1_U67 (.A( u2_u13_u1_n152 ) , .ZN( u2_u13_u1_n173 ) );
  INV_X1 u2_u13_u1_U68 (.A( u2_u13_u1_n128 ) , .ZN( u2_u13_u1_n172 ) );
  NAND2_X1 u2_u13_u1_U69 (.A2( u2_u13_u1_n102 ) , .A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n123 ) );
  INV_X1 u2_u13_u1_U7 (.A( u2_u13_u1_n147 ) , .ZN( u2_u13_u1_n181 ) );
  NOR2_X1 u2_u13_u1_U70 (.A2( u2_u13_X_7 ) , .A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n95 ) );
  NOR2_X1 u2_u13_u1_U71 (.A1( u2_u13_X_12 ) , .A2( u2_u13_X_9 ) , .ZN( u2_u13_u1_n100 ) );
  NOR2_X1 u2_u13_u1_U72 (.A2( u2_u13_X_8 ) , .A1( u2_u13_u1_n177 ) , .ZN( u2_u13_u1_n99 ) );
  NOR2_X1 u2_u13_u1_U73 (.A2( u2_u13_X_12 ) , .ZN( u2_u13_u1_n102 ) , .A1( u2_u13_u1_n176 ) );
  NOR2_X1 u2_u13_u1_U74 (.A2( u2_u13_X_9 ) , .ZN( u2_u13_u1_n105 ) , .A1( u2_u13_u1_n168 ) );
  NAND2_X1 u2_u13_u1_U75 (.A1( u2_u13_X_10 ) , .ZN( u2_u13_u1_n160 ) , .A2( u2_u13_u1_n169 ) );
  NAND2_X1 u2_u13_u1_U76 (.A2( u2_u13_X_10 ) , .A1( u2_u13_X_11 ) , .ZN( u2_u13_u1_n152 ) );
  NAND2_X1 u2_u13_u1_U77 (.A1( u2_u13_X_11 ) , .ZN( u2_u13_u1_n128 ) , .A2( u2_u13_u1_n170 ) );
  AND2_X1 u2_u13_u1_U78 (.A2( u2_u13_X_7 ) , .A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n104 ) );
  AND2_X1 u2_u13_u1_U79 (.A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n103 ) , .A2( u2_u13_u1_n177 ) );
  NOR2_X1 u2_u13_u1_U8 (.A1( u2_u13_u1_n112 ) , .A2( u2_u13_u1_n116 ) , .ZN( u2_u13_u1_n118 ) );
  INV_X1 u2_u13_u1_U80 (.A( u2_u13_X_10 ) , .ZN( u2_u13_u1_n170 ) );
  INV_X1 u2_u13_u1_U81 (.A( u2_u13_X_9 ) , .ZN( u2_u13_u1_n176 ) );
  INV_X1 u2_u13_u1_U82 (.A( u2_u13_X_11 ) , .ZN( u2_u13_u1_n169 ) );
  INV_X1 u2_u13_u1_U83 (.A( u2_u13_X_12 ) , .ZN( u2_u13_u1_n168 ) );
  INV_X1 u2_u13_u1_U84 (.A( u2_u13_X_7 ) , .ZN( u2_u13_u1_n177 ) );
  NAND4_X1 u2_u13_u1_U85 (.ZN( u2_out13_28 ) , .A4( u2_u13_u1_n124 ) , .A3( u2_u13_u1_n125 ) , .A2( u2_u13_u1_n126 ) , .A1( u2_u13_u1_n127 ) );
  OAI21_X1 u2_u13_u1_U86 (.ZN( u2_u13_u1_n127 ) , .B2( u2_u13_u1_n139 ) , .B1( u2_u13_u1_n175 ) , .A( u2_u13_u1_n183 ) );
  OAI21_X1 u2_u13_u1_U87 (.ZN( u2_u13_u1_n126 ) , .B2( u2_u13_u1_n140 ) , .A( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n178 ) );
  NAND4_X1 u2_u13_u1_U88 (.ZN( u2_out13_18 ) , .A4( u2_u13_u1_n165 ) , .A3( u2_u13_u1_n166 ) , .A1( u2_u13_u1_n167 ) , .A2( u2_u13_u1_n186 ) );
  AOI22_X1 u2_u13_u1_U89 (.B2( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n147 ) , .A2( u2_u13_u1_n148 ) , .ZN( u2_u13_u1_n166 ) , .A1( u2_u13_u1_n172 ) );
  OAI21_X1 u2_u13_u1_U9 (.ZN( u2_u13_u1_n101 ) , .B1( u2_u13_u1_n141 ) , .A( u2_u13_u1_n146 ) , .B2( u2_u13_u1_n183 ) );
  INV_X1 u2_u13_u1_U90 (.A( u2_u13_u1_n145 ) , .ZN( u2_u13_u1_n186 ) );
  NAND4_X1 u2_u13_u1_U91 (.ZN( u2_out13_2 ) , .A4( u2_u13_u1_n142 ) , .A3( u2_u13_u1_n143 ) , .A2( u2_u13_u1_n144 ) , .A1( u2_u13_u1_n179 ) );
  OAI21_X1 u2_u13_u1_U92 (.B2( u2_u13_u1_n132 ) , .ZN( u2_u13_u1_n144 ) , .A( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n180 ) );
  INV_X1 u2_u13_u1_U93 (.A( u2_u13_u1_n130 ) , .ZN( u2_u13_u1_n179 ) );
  OR4_X1 u2_u13_u1_U94 (.ZN( u2_out13_13 ) , .A4( u2_u13_u1_n108 ) , .A3( u2_u13_u1_n109 ) , .A2( u2_u13_u1_n110 ) , .A1( u2_u13_u1_n111 ) );
  AOI21_X1 u2_u13_u1_U95 (.ZN( u2_u13_u1_n111 ) , .A( u2_u13_u1_n128 ) , .B2( u2_u13_u1_n131 ) , .B1( u2_u13_u1_n135 ) );
  AOI21_X1 u2_u13_u1_U96 (.ZN( u2_u13_u1_n110 ) , .A( u2_u13_u1_n116 ) , .B1( u2_u13_u1_n152 ) , .B2( u2_u13_u1_n160 ) );
  NAND3_X1 u2_u13_u1_U97 (.A3( u2_u13_u1_n149 ) , .A2( u2_u13_u1_n150 ) , .A1( u2_u13_u1_n151 ) , .ZN( u2_u13_u1_n164 ) );
  NAND3_X1 u2_u13_u1_U98 (.A3( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n135 ) , .ZN( u2_u13_u1_n136 ) , .A1( u2_u13_u1_n151 ) );
  NAND3_X1 u2_u13_u1_U99 (.A1( u2_u13_u1_n133 ) , .ZN( u2_u13_u1_n137 ) , .A2( u2_u13_u1_n154 ) , .A3( u2_u13_u1_n181 ) );
  OAI22_X1 u2_u13_u2_U10 (.B1( u2_u13_u2_n151 ) , .A2( u2_u13_u2_n152 ) , .A1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n160 ) , .B2( u2_u13_u2_n168 ) );
  NAND3_X1 u2_u13_u2_U100 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n98 ) );
  NOR3_X1 u2_u13_u2_U11 (.A1( u2_u13_u2_n150 ) , .ZN( u2_u13_u2_n151 ) , .A3( u2_u13_u2_n175 ) , .A2( u2_u13_u2_n188 ) );
  AOI21_X1 u2_u13_u2_U12 (.B2( u2_u13_u2_n123 ) , .ZN( u2_u13_u2_n125 ) , .A( u2_u13_u2_n171 ) , .B1( u2_u13_u2_n184 ) );
  INV_X1 u2_u13_u2_U13 (.A( u2_u13_u2_n150 ) , .ZN( u2_u13_u2_n184 ) );
  AOI21_X1 u2_u13_u2_U14 (.ZN( u2_u13_u2_n144 ) , .B2( u2_u13_u2_n155 ) , .A( u2_u13_u2_n172 ) , .B1( u2_u13_u2_n185 ) );
  AOI21_X1 u2_u13_u2_U15 (.B2( u2_u13_u2_n143 ) , .ZN( u2_u13_u2_n145 ) , .B1( u2_u13_u2_n152 ) , .A( u2_u13_u2_n171 ) );
  INV_X1 u2_u13_u2_U16 (.A( u2_u13_u2_n156 ) , .ZN( u2_u13_u2_n171 ) );
  INV_X1 u2_u13_u2_U17 (.A( u2_u13_u2_n120 ) , .ZN( u2_u13_u2_n188 ) );
  NAND2_X1 u2_u13_u2_U18 (.A2( u2_u13_u2_n122 ) , .ZN( u2_u13_u2_n150 ) , .A1( u2_u13_u2_n152 ) );
  INV_X1 u2_u13_u2_U19 (.A( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n170 ) );
  INV_X1 u2_u13_u2_U20 (.A( u2_u13_u2_n137 ) , .ZN( u2_u13_u2_n173 ) );
  NAND2_X1 u2_u13_u2_U21 (.A1( u2_u13_u2_n132 ) , .A2( u2_u13_u2_n139 ) , .ZN( u2_u13_u2_n157 ) );
  INV_X1 u2_u13_u2_U22 (.A( u2_u13_u2_n113 ) , .ZN( u2_u13_u2_n178 ) );
  INV_X1 u2_u13_u2_U23 (.A( u2_u13_u2_n139 ) , .ZN( u2_u13_u2_n175 ) );
  INV_X1 u2_u13_u2_U24 (.A( u2_u13_u2_n155 ) , .ZN( u2_u13_u2_n181 ) );
  INV_X1 u2_u13_u2_U25 (.A( u2_u13_u2_n119 ) , .ZN( u2_u13_u2_n177 ) );
  INV_X1 u2_u13_u2_U26 (.A( u2_u13_u2_n116 ) , .ZN( u2_u13_u2_n180 ) );
  INV_X1 u2_u13_u2_U27 (.A( u2_u13_u2_n131 ) , .ZN( u2_u13_u2_n179 ) );
  INV_X1 u2_u13_u2_U28 (.A( u2_u13_u2_n154 ) , .ZN( u2_u13_u2_n176 ) );
  NAND2_X1 u2_u13_u2_U29 (.A2( u2_u13_u2_n116 ) , .A1( u2_u13_u2_n117 ) , .ZN( u2_u13_u2_n118 ) );
  NOR2_X1 u2_u13_u2_U3 (.ZN( u2_u13_u2_n121 ) , .A2( u2_u13_u2_n177 ) , .A1( u2_u13_u2_n180 ) );
  INV_X1 u2_u13_u2_U30 (.A( u2_u13_u2_n132 ) , .ZN( u2_u13_u2_n182 ) );
  INV_X1 u2_u13_u2_U31 (.A( u2_u13_u2_n158 ) , .ZN( u2_u13_u2_n183 ) );
  OAI21_X1 u2_u13_u2_U32 (.A( u2_u13_u2_n156 ) , .B1( u2_u13_u2_n157 ) , .ZN( u2_u13_u2_n158 ) , .B2( u2_u13_u2_n179 ) );
  NOR2_X1 u2_u13_u2_U33 (.ZN( u2_u13_u2_n156 ) , .A1( u2_u13_u2_n166 ) , .A2( u2_u13_u2_n169 ) );
  NOR2_X1 u2_u13_u2_U34 (.A2( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n137 ) , .A1( u2_u13_u2_n140 ) );
  NOR2_X1 u2_u13_u2_U35 (.A2( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n153 ) , .A1( u2_u13_u2_n156 ) );
  AOI211_X1 u2_u13_u2_U36 (.ZN( u2_u13_u2_n130 ) , .C1( u2_u13_u2_n138 ) , .C2( u2_u13_u2_n179 ) , .B( u2_u13_u2_n96 ) , .A( u2_u13_u2_n97 ) );
  OAI22_X1 u2_u13_u2_U37 (.B1( u2_u13_u2_n133 ) , .A2( u2_u13_u2_n137 ) , .A1( u2_u13_u2_n152 ) , .B2( u2_u13_u2_n168 ) , .ZN( u2_u13_u2_n97 ) );
  OAI221_X1 u2_u13_u2_U38 (.B1( u2_u13_u2_n113 ) , .C1( u2_u13_u2_n132 ) , .A( u2_u13_u2_n149 ) , .B2( u2_u13_u2_n171 ) , .C2( u2_u13_u2_n172 ) , .ZN( u2_u13_u2_n96 ) );
  OAI221_X1 u2_u13_u2_U39 (.A( u2_u13_u2_n115 ) , .C2( u2_u13_u2_n123 ) , .B2( u2_u13_u2_n143 ) , .B1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n163 ) , .C1( u2_u13_u2_n168 ) );
  INV_X1 u2_u13_u2_U4 (.A( u2_u13_u2_n134 ) , .ZN( u2_u13_u2_n185 ) );
  OAI21_X1 u2_u13_u2_U40 (.A( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n115 ) , .B1( u2_u13_u2_n176 ) , .B2( u2_u13_u2_n178 ) );
  OAI221_X1 u2_u13_u2_U41 (.A( u2_u13_u2_n135 ) , .B2( u2_u13_u2_n136 ) , .B1( u2_u13_u2_n137 ) , .ZN( u2_u13_u2_n162 ) , .C2( u2_u13_u2_n167 ) , .C1( u2_u13_u2_n185 ) );
  AND3_X1 u2_u13_u2_U42 (.A3( u2_u13_u2_n131 ) , .A2( u2_u13_u2_n132 ) , .A1( u2_u13_u2_n133 ) , .ZN( u2_u13_u2_n136 ) );
  AOI22_X1 u2_u13_u2_U43 (.ZN( u2_u13_u2_n135 ) , .B1( u2_u13_u2_n140 ) , .A1( u2_u13_u2_n156 ) , .B2( u2_u13_u2_n180 ) , .A2( u2_u13_u2_n188 ) );
  AOI21_X1 u2_u13_u2_U44 (.ZN( u2_u13_u2_n149 ) , .B1( u2_u13_u2_n173 ) , .B2( u2_u13_u2_n188 ) , .A( u2_u13_u2_n95 ) );
  AND3_X1 u2_u13_u2_U45 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n156 ) , .ZN( u2_u13_u2_n95 ) );
  OAI21_X1 u2_u13_u2_U46 (.A( u2_u13_u2_n141 ) , .B2( u2_u13_u2_n142 ) , .ZN( u2_u13_u2_n146 ) , .B1( u2_u13_u2_n153 ) );
  OAI21_X1 u2_u13_u2_U47 (.A( u2_u13_u2_n140 ) , .ZN( u2_u13_u2_n141 ) , .B1( u2_u13_u2_n176 ) , .B2( u2_u13_u2_n177 ) );
  NOR3_X1 u2_u13_u2_U48 (.ZN( u2_u13_u2_n142 ) , .A3( u2_u13_u2_n175 ) , .A2( u2_u13_u2_n178 ) , .A1( u2_u13_u2_n181 ) );
  OAI21_X1 u2_u13_u2_U49 (.A( u2_u13_u2_n101 ) , .B2( u2_u13_u2_n121 ) , .B1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n164 ) );
  NOR4_X1 u2_u13_u2_U5 (.A4( u2_u13_u2_n124 ) , .A3( u2_u13_u2_n125 ) , .A2( u2_u13_u2_n126 ) , .A1( u2_u13_u2_n127 ) , .ZN( u2_u13_u2_n128 ) );
  NAND2_X1 u2_u13_u2_U50 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n155 ) );
  NAND2_X1 u2_u13_u2_U51 (.A2( u2_u13_u2_n105 ) , .A1( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n143 ) );
  NAND2_X1 u2_u13_u2_U52 (.A1( u2_u13_u2_n104 ) , .A2( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n152 ) );
  NAND2_X1 u2_u13_u2_U53 (.A1( u2_u13_u2_n100 ) , .A2( u2_u13_u2_n105 ) , .ZN( u2_u13_u2_n132 ) );
  INV_X1 u2_u13_u2_U54 (.A( u2_u13_u2_n140 ) , .ZN( u2_u13_u2_n168 ) );
  INV_X1 u2_u13_u2_U55 (.A( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n167 ) );
  NAND2_X1 u2_u13_u2_U56 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n113 ) );
  NAND2_X1 u2_u13_u2_U57 (.A1( u2_u13_u2_n106 ) , .A2( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n131 ) );
  NAND2_X1 u2_u13_u2_U58 (.A1( u2_u13_u2_n103 ) , .A2( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n139 ) );
  NAND2_X1 u2_u13_u2_U59 (.A1( u2_u13_u2_n103 ) , .A2( u2_u13_u2_n105 ) , .ZN( u2_u13_u2_n133 ) );
  AOI21_X1 u2_u13_u2_U6 (.B2( u2_u13_u2_n119 ) , .ZN( u2_u13_u2_n127 ) , .A( u2_u13_u2_n137 ) , .B1( u2_u13_u2_n155 ) );
  NAND2_X1 u2_u13_u2_U60 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n103 ) , .ZN( u2_u13_u2_n154 ) );
  NAND2_X1 u2_u13_u2_U61 (.A2( u2_u13_u2_n103 ) , .A1( u2_u13_u2_n104 ) , .ZN( u2_u13_u2_n119 ) );
  NAND2_X1 u2_u13_u2_U62 (.A2( u2_u13_u2_n107 ) , .A1( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n123 ) );
  NAND2_X1 u2_u13_u2_U63 (.A1( u2_u13_u2_n104 ) , .A2( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n122 ) );
  INV_X1 u2_u13_u2_U64 (.A( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n172 ) );
  NAND2_X1 u2_u13_u2_U65 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n102 ) , .ZN( u2_u13_u2_n116 ) );
  NAND2_X1 u2_u13_u2_U66 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n120 ) );
  NAND2_X1 u2_u13_u2_U67 (.A2( u2_u13_u2_n105 ) , .A1( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n117 ) );
  INV_X1 u2_u13_u2_U68 (.ZN( u2_u13_u2_n187 ) , .A( u2_u13_u2_n99 ) );
  OAI21_X1 u2_u13_u2_U69 (.B1( u2_u13_u2_n137 ) , .B2( u2_u13_u2_n143 ) , .A( u2_u13_u2_n98 ) , .ZN( u2_u13_u2_n99 ) );
  AOI21_X1 u2_u13_u2_U7 (.ZN( u2_u13_u2_n124 ) , .B1( u2_u13_u2_n131 ) , .B2( u2_u13_u2_n143 ) , .A( u2_u13_u2_n172 ) );
  NOR2_X1 u2_u13_u2_U70 (.A2( u2_u13_X_16 ) , .ZN( u2_u13_u2_n140 ) , .A1( u2_u13_u2_n166 ) );
  NOR2_X1 u2_u13_u2_U71 (.A2( u2_u13_X_13 ) , .A1( u2_u13_X_14 ) , .ZN( u2_u13_u2_n100 ) );
  NOR2_X1 u2_u13_u2_U72 (.A2( u2_u13_X_16 ) , .A1( u2_u13_X_17 ) , .ZN( u2_u13_u2_n138 ) );
  NOR2_X1 u2_u13_u2_U73 (.A2( u2_u13_X_15 ) , .A1( u2_u13_X_18 ) , .ZN( u2_u13_u2_n104 ) );
  NOR2_X1 u2_u13_u2_U74 (.A2( u2_u13_X_14 ) , .ZN( u2_u13_u2_n103 ) , .A1( u2_u13_u2_n174 ) );
  NOR2_X1 u2_u13_u2_U75 (.A2( u2_u13_X_15 ) , .ZN( u2_u13_u2_n102 ) , .A1( u2_u13_u2_n165 ) );
  NOR2_X1 u2_u13_u2_U76 (.A2( u2_u13_X_17 ) , .ZN( u2_u13_u2_n114 ) , .A1( u2_u13_u2_n169 ) );
  AND2_X1 u2_u13_u2_U77 (.A1( u2_u13_X_15 ) , .ZN( u2_u13_u2_n105 ) , .A2( u2_u13_u2_n165 ) );
  AND2_X1 u2_u13_u2_U78 (.A2( u2_u13_X_15 ) , .A1( u2_u13_X_18 ) , .ZN( u2_u13_u2_n107 ) );
  AND2_X1 u2_u13_u2_U79 (.A1( u2_u13_X_14 ) , .ZN( u2_u13_u2_n106 ) , .A2( u2_u13_u2_n174 ) );
  AOI21_X1 u2_u13_u2_U8 (.B2( u2_u13_u2_n120 ) , .B1( u2_u13_u2_n121 ) , .ZN( u2_u13_u2_n126 ) , .A( u2_u13_u2_n167 ) );
  AND2_X1 u2_u13_u2_U80 (.A1( u2_u13_X_13 ) , .A2( u2_u13_X_14 ) , .ZN( u2_u13_u2_n108 ) );
  INV_X1 u2_u13_u2_U81 (.A( u2_u13_X_16 ) , .ZN( u2_u13_u2_n169 ) );
  INV_X1 u2_u13_u2_U82 (.A( u2_u13_X_17 ) , .ZN( u2_u13_u2_n166 ) );
  INV_X1 u2_u13_u2_U83 (.A( u2_u13_X_13 ) , .ZN( u2_u13_u2_n174 ) );
  INV_X1 u2_u13_u2_U84 (.A( u2_u13_X_18 ) , .ZN( u2_u13_u2_n165 ) );
  NAND4_X1 u2_u13_u2_U85 (.ZN( u2_out13_30 ) , .A4( u2_u13_u2_n147 ) , .A3( u2_u13_u2_n148 ) , .A2( u2_u13_u2_n149 ) , .A1( u2_u13_u2_n187 ) );
  AOI21_X1 u2_u13_u2_U86 (.B2( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n148 ) , .A( u2_u13_u2_n162 ) , .B1( u2_u13_u2_n182 ) );
  NOR3_X1 u2_u13_u2_U87 (.A3( u2_u13_u2_n144 ) , .A2( u2_u13_u2_n145 ) , .A1( u2_u13_u2_n146 ) , .ZN( u2_u13_u2_n147 ) );
  NAND4_X1 u2_u13_u2_U88 (.ZN( u2_out13_24 ) , .A4( u2_u13_u2_n111 ) , .A3( u2_u13_u2_n112 ) , .A1( u2_u13_u2_n130 ) , .A2( u2_u13_u2_n187 ) );
  AOI221_X1 u2_u13_u2_U89 (.A( u2_u13_u2_n109 ) , .B1( u2_u13_u2_n110 ) , .ZN( u2_u13_u2_n111 ) , .C1( u2_u13_u2_n134 ) , .C2( u2_u13_u2_n170 ) , .B2( u2_u13_u2_n173 ) );
  OAI22_X1 u2_u13_u2_U9 (.ZN( u2_u13_u2_n109 ) , .A2( u2_u13_u2_n113 ) , .B2( u2_u13_u2_n133 ) , .B1( u2_u13_u2_n167 ) , .A1( u2_u13_u2_n168 ) );
  AOI21_X1 u2_u13_u2_U90 (.ZN( u2_u13_u2_n112 ) , .B2( u2_u13_u2_n156 ) , .A( u2_u13_u2_n164 ) , .B1( u2_u13_u2_n181 ) );
  NAND4_X1 u2_u13_u2_U91 (.ZN( u2_out13_16 ) , .A4( u2_u13_u2_n128 ) , .A3( u2_u13_u2_n129 ) , .A1( u2_u13_u2_n130 ) , .A2( u2_u13_u2_n186 ) );
  AOI22_X1 u2_u13_u2_U92 (.A2( u2_u13_u2_n118 ) , .ZN( u2_u13_u2_n129 ) , .A1( u2_u13_u2_n140 ) , .B1( u2_u13_u2_n157 ) , .B2( u2_u13_u2_n170 ) );
  INV_X1 u2_u13_u2_U93 (.A( u2_u13_u2_n163 ) , .ZN( u2_u13_u2_n186 ) );
  OR4_X1 u2_u13_u2_U94 (.ZN( u2_out13_6 ) , .A4( u2_u13_u2_n161 ) , .A3( u2_u13_u2_n162 ) , .A2( u2_u13_u2_n163 ) , .A1( u2_u13_u2_n164 ) );
  OR3_X1 u2_u13_u2_U95 (.A2( u2_u13_u2_n159 ) , .A1( u2_u13_u2_n160 ) , .ZN( u2_u13_u2_n161 ) , .A3( u2_u13_u2_n183 ) );
  AOI21_X1 u2_u13_u2_U96 (.B2( u2_u13_u2_n154 ) , .B1( u2_u13_u2_n155 ) , .ZN( u2_u13_u2_n159 ) , .A( u2_u13_u2_n167 ) );
  NAND3_X1 u2_u13_u2_U97 (.A2( u2_u13_u2_n117 ) , .A1( u2_u13_u2_n122 ) , .A3( u2_u13_u2_n123 ) , .ZN( u2_u13_u2_n134 ) );
  NAND3_X1 u2_u13_u2_U98 (.ZN( u2_u13_u2_n110 ) , .A2( u2_u13_u2_n131 ) , .A3( u2_u13_u2_n139 ) , .A1( u2_u13_u2_n154 ) );
  NAND3_X1 u2_u13_u2_U99 (.A2( u2_u13_u2_n100 ) , .ZN( u2_u13_u2_n101 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n114 ) );
  OAI22_X1 u2_u13_u3_U10 (.B1( u2_u13_u3_n113 ) , .A2( u2_u13_u3_n135 ) , .A1( u2_u13_u3_n150 ) , .B2( u2_u13_u3_n164 ) , .ZN( u2_u13_u3_n98 ) );
  OAI211_X1 u2_u13_u3_U11 (.B( u2_u13_u3_n106 ) , .ZN( u2_u13_u3_n119 ) , .C2( u2_u13_u3_n128 ) , .C1( u2_u13_u3_n167 ) , .A( u2_u13_u3_n181 ) );
  AOI221_X1 u2_u13_u3_U12 (.C1( u2_u13_u3_n105 ) , .ZN( u2_u13_u3_n106 ) , .A( u2_u13_u3_n131 ) , .B2( u2_u13_u3_n132 ) , .C2( u2_u13_u3_n133 ) , .B1( u2_u13_u3_n169 ) );
  INV_X1 u2_u13_u3_U13 (.ZN( u2_u13_u3_n181 ) , .A( u2_u13_u3_n98 ) );
  NAND2_X1 u2_u13_u3_U14 (.ZN( u2_u13_u3_n105 ) , .A2( u2_u13_u3_n130 ) , .A1( u2_u13_u3_n155 ) );
  AOI22_X1 u2_u13_u3_U15 (.B1( u2_u13_u3_n115 ) , .A2( u2_u13_u3_n116 ) , .ZN( u2_u13_u3_n123 ) , .B2( u2_u13_u3_n133 ) , .A1( u2_u13_u3_n169 ) );
  NAND2_X1 u2_u13_u3_U16 (.ZN( u2_u13_u3_n116 ) , .A2( u2_u13_u3_n151 ) , .A1( u2_u13_u3_n182 ) );
  NOR2_X1 u2_u13_u3_U17 (.ZN( u2_u13_u3_n126 ) , .A2( u2_u13_u3_n150 ) , .A1( u2_u13_u3_n164 ) );
  AOI21_X1 u2_u13_u3_U18 (.ZN( u2_u13_u3_n112 ) , .B2( u2_u13_u3_n146 ) , .B1( u2_u13_u3_n155 ) , .A( u2_u13_u3_n167 ) );
  NAND2_X1 u2_u13_u3_U19 (.A1( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n142 ) , .A2( u2_u13_u3_n164 ) );
  NAND2_X1 u2_u13_u3_U20 (.ZN( u2_u13_u3_n132 ) , .A2( u2_u13_u3_n152 ) , .A1( u2_u13_u3_n156 ) );
  AND2_X1 u2_u13_u3_U21 (.A2( u2_u13_u3_n113 ) , .A1( u2_u13_u3_n114 ) , .ZN( u2_u13_u3_n151 ) );
  INV_X1 u2_u13_u3_U22 (.A( u2_u13_u3_n133 ) , .ZN( u2_u13_u3_n165 ) );
  INV_X1 u2_u13_u3_U23 (.A( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n170 ) );
  NAND2_X1 u2_u13_u3_U24 (.A1( u2_u13_u3_n107 ) , .A2( u2_u13_u3_n108 ) , .ZN( u2_u13_u3_n140 ) );
  NAND2_X1 u2_u13_u3_U25 (.ZN( u2_u13_u3_n117 ) , .A1( u2_u13_u3_n124 ) , .A2( u2_u13_u3_n148 ) );
  NAND2_X1 u2_u13_u3_U26 (.ZN( u2_u13_u3_n143 ) , .A1( u2_u13_u3_n165 ) , .A2( u2_u13_u3_n167 ) );
  INV_X1 u2_u13_u3_U27 (.A( u2_u13_u3_n130 ) , .ZN( u2_u13_u3_n177 ) );
  INV_X1 u2_u13_u3_U28 (.A( u2_u13_u3_n128 ) , .ZN( u2_u13_u3_n176 ) );
  INV_X1 u2_u13_u3_U29 (.A( u2_u13_u3_n155 ) , .ZN( u2_u13_u3_n174 ) );
  INV_X1 u2_u13_u3_U3 (.A( u2_u13_u3_n129 ) , .ZN( u2_u13_u3_n183 ) );
  INV_X1 u2_u13_u3_U30 (.A( u2_u13_u3_n139 ) , .ZN( u2_u13_u3_n185 ) );
  NOR2_X1 u2_u13_u3_U31 (.ZN( u2_u13_u3_n135 ) , .A2( u2_u13_u3_n141 ) , .A1( u2_u13_u3_n169 ) );
  OAI222_X1 u2_u13_u3_U32 (.C2( u2_u13_u3_n107 ) , .A2( u2_u13_u3_n108 ) , .B1( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n138 ) , .B2( u2_u13_u3_n146 ) , .C1( u2_u13_u3_n154 ) , .A1( u2_u13_u3_n164 ) );
  NOR4_X1 u2_u13_u3_U33 (.A4( u2_u13_u3_n157 ) , .A3( u2_u13_u3_n158 ) , .A2( u2_u13_u3_n159 ) , .A1( u2_u13_u3_n160 ) , .ZN( u2_u13_u3_n161 ) );
  AOI21_X1 u2_u13_u3_U34 (.B2( u2_u13_u3_n152 ) , .B1( u2_u13_u3_n153 ) , .ZN( u2_u13_u3_n158 ) , .A( u2_u13_u3_n164 ) );
  AOI21_X1 u2_u13_u3_U35 (.A( u2_u13_u3_n154 ) , .B2( u2_u13_u3_n155 ) , .B1( u2_u13_u3_n156 ) , .ZN( u2_u13_u3_n157 ) );
  AOI21_X1 u2_u13_u3_U36 (.A( u2_u13_u3_n149 ) , .B2( u2_u13_u3_n150 ) , .B1( u2_u13_u3_n151 ) , .ZN( u2_u13_u3_n159 ) );
  AOI211_X1 u2_u13_u3_U37 (.ZN( u2_u13_u3_n109 ) , .A( u2_u13_u3_n119 ) , .C2( u2_u13_u3_n129 ) , .B( u2_u13_u3_n138 ) , .C1( u2_u13_u3_n141 ) );
  AOI211_X1 u2_u13_u3_U38 (.B( u2_u13_u3_n119 ) , .A( u2_u13_u3_n120 ) , .C2( u2_u13_u3_n121 ) , .ZN( u2_u13_u3_n122 ) , .C1( u2_u13_u3_n179 ) );
  INV_X1 u2_u13_u3_U39 (.A( u2_u13_u3_n156 ) , .ZN( u2_u13_u3_n179 ) );
  INV_X1 u2_u13_u3_U4 (.A( u2_u13_u3_n140 ) , .ZN( u2_u13_u3_n182 ) );
  OAI22_X1 u2_u13_u3_U40 (.B1( u2_u13_u3_n118 ) , .ZN( u2_u13_u3_n120 ) , .A1( u2_u13_u3_n135 ) , .B2( u2_u13_u3_n154 ) , .A2( u2_u13_u3_n178 ) );
  AND3_X1 u2_u13_u3_U41 (.ZN( u2_u13_u3_n118 ) , .A2( u2_u13_u3_n124 ) , .A1( u2_u13_u3_n144 ) , .A3( u2_u13_u3_n152 ) );
  INV_X1 u2_u13_u3_U42 (.A( u2_u13_u3_n121 ) , .ZN( u2_u13_u3_n164 ) );
  NAND2_X1 u2_u13_u3_U43 (.ZN( u2_u13_u3_n133 ) , .A1( u2_u13_u3_n154 ) , .A2( u2_u13_u3_n164 ) );
  OAI211_X1 u2_u13_u3_U44 (.B( u2_u13_u3_n127 ) , .ZN( u2_u13_u3_n139 ) , .C1( u2_u13_u3_n150 ) , .C2( u2_u13_u3_n154 ) , .A( u2_u13_u3_n184 ) );
  INV_X1 u2_u13_u3_U45 (.A( u2_u13_u3_n125 ) , .ZN( u2_u13_u3_n184 ) );
  AOI221_X1 u2_u13_u3_U46 (.A( u2_u13_u3_n126 ) , .ZN( u2_u13_u3_n127 ) , .C2( u2_u13_u3_n132 ) , .C1( u2_u13_u3_n169 ) , .B2( u2_u13_u3_n170 ) , .B1( u2_u13_u3_n174 ) );
  OAI22_X1 u2_u13_u3_U47 (.A1( u2_u13_u3_n124 ) , .ZN( u2_u13_u3_n125 ) , .B2( u2_u13_u3_n145 ) , .A2( u2_u13_u3_n165 ) , .B1( u2_u13_u3_n167 ) );
  NOR2_X1 u2_u13_u3_U48 (.A1( u2_u13_u3_n113 ) , .ZN( u2_u13_u3_n131 ) , .A2( u2_u13_u3_n154 ) );
  NAND2_X1 u2_u13_u3_U49 (.A1( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n150 ) , .A2( u2_u13_u3_n99 ) );
  INV_X1 u2_u13_u3_U5 (.A( u2_u13_u3_n117 ) , .ZN( u2_u13_u3_n178 ) );
  NAND2_X1 u2_u13_u3_U50 (.A2( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n155 ) , .A1( u2_u13_u3_n97 ) );
  INV_X1 u2_u13_u3_U51 (.A( u2_u13_u3_n141 ) , .ZN( u2_u13_u3_n167 ) );
  AOI21_X1 u2_u13_u3_U52 (.B2( u2_u13_u3_n114 ) , .B1( u2_u13_u3_n146 ) , .A( u2_u13_u3_n154 ) , .ZN( u2_u13_u3_n94 ) );
  AOI21_X1 u2_u13_u3_U53 (.ZN( u2_u13_u3_n110 ) , .B2( u2_u13_u3_n142 ) , .B1( u2_u13_u3_n186 ) , .A( u2_u13_u3_n95 ) );
  INV_X1 u2_u13_u3_U54 (.A( u2_u13_u3_n145 ) , .ZN( u2_u13_u3_n186 ) );
  AOI21_X1 u2_u13_u3_U55 (.B1( u2_u13_u3_n124 ) , .A( u2_u13_u3_n149 ) , .B2( u2_u13_u3_n155 ) , .ZN( u2_u13_u3_n95 ) );
  INV_X1 u2_u13_u3_U56 (.A( u2_u13_u3_n149 ) , .ZN( u2_u13_u3_n169 ) );
  NAND2_X1 u2_u13_u3_U57 (.ZN( u2_u13_u3_n124 ) , .A1( u2_u13_u3_n96 ) , .A2( u2_u13_u3_n97 ) );
  NAND2_X1 u2_u13_u3_U58 (.A2( u2_u13_u3_n100 ) , .ZN( u2_u13_u3_n146 ) , .A1( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U59 (.A1( u2_u13_u3_n101 ) , .ZN( u2_u13_u3_n145 ) , .A2( u2_u13_u3_n99 ) );
  AOI221_X1 u2_u13_u3_U6 (.A( u2_u13_u3_n131 ) , .C2( u2_u13_u3_n132 ) , .C1( u2_u13_u3_n133 ) , .ZN( u2_u13_u3_n134 ) , .B1( u2_u13_u3_n143 ) , .B2( u2_u13_u3_n177 ) );
  NAND2_X1 u2_u13_u3_U60 (.A1( u2_u13_u3_n100 ) , .ZN( u2_u13_u3_n156 ) , .A2( u2_u13_u3_n99 ) );
  NAND2_X1 u2_u13_u3_U61 (.A2( u2_u13_u3_n101 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n148 ) );
  NAND2_X1 u2_u13_u3_U62 (.A1( u2_u13_u3_n100 ) , .A2( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n128 ) );
  NAND2_X1 u2_u13_u3_U63 (.A2( u2_u13_u3_n101 ) , .A1( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n152 ) );
  NAND2_X1 u2_u13_u3_U64 (.A2( u2_u13_u3_n101 ) , .ZN( u2_u13_u3_n114 ) , .A1( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U65 (.ZN( u2_u13_u3_n107 ) , .A1( u2_u13_u3_n97 ) , .A2( u2_u13_u3_n99 ) );
  NAND2_X1 u2_u13_u3_U66 (.A2( u2_u13_u3_n100 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n113 ) );
  NAND2_X1 u2_u13_u3_U67 (.A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n153 ) , .A2( u2_u13_u3_n97 ) );
  NAND2_X1 u2_u13_u3_U68 (.A2( u2_u13_u3_n103 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n130 ) );
  NAND2_X1 u2_u13_u3_U69 (.A2( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n144 ) , .A1( u2_u13_u3_n96 ) );
  OAI22_X1 u2_u13_u3_U7 (.B2( u2_u13_u3_n147 ) , .A2( u2_u13_u3_n148 ) , .ZN( u2_u13_u3_n160 ) , .B1( u2_u13_u3_n165 ) , .A1( u2_u13_u3_n168 ) );
  NAND2_X1 u2_u13_u3_U70 (.A1( u2_u13_u3_n102 ) , .A2( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n108 ) );
  NOR2_X1 u2_u13_u3_U71 (.A2( u2_u13_X_19 ) , .A1( u2_u13_X_20 ) , .ZN( u2_u13_u3_n99 ) );
  NOR2_X1 u2_u13_u3_U72 (.A2( u2_u13_X_21 ) , .A1( u2_u13_X_24 ) , .ZN( u2_u13_u3_n103 ) );
  NOR2_X1 u2_u13_u3_U73 (.A2( u2_u13_X_24 ) , .A1( u2_u13_u3_n171 ) , .ZN( u2_u13_u3_n97 ) );
  NOR2_X1 u2_u13_u3_U74 (.A2( u2_u13_X_23 ) , .ZN( u2_u13_u3_n141 ) , .A1( u2_u13_u3_n166 ) );
  NOR2_X1 u2_u13_u3_U75 (.A2( u2_u13_X_19 ) , .A1( u2_u13_u3_n172 ) , .ZN( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U76 (.A1( u2_u13_X_22 ) , .A2( u2_u13_X_23 ) , .ZN( u2_u13_u3_n154 ) );
  NAND2_X1 u2_u13_u3_U77 (.A1( u2_u13_X_23 ) , .ZN( u2_u13_u3_n149 ) , .A2( u2_u13_u3_n166 ) );
  NOR2_X1 u2_u13_u3_U78 (.A2( u2_u13_X_22 ) , .A1( u2_u13_X_23 ) , .ZN( u2_u13_u3_n121 ) );
  AND2_X1 u2_u13_u3_U79 (.A1( u2_u13_X_24 ) , .ZN( u2_u13_u3_n101 ) , .A2( u2_u13_u3_n171 ) );
  AND3_X1 u2_u13_u3_U8 (.A3( u2_u13_u3_n144 ) , .A2( u2_u13_u3_n145 ) , .A1( u2_u13_u3_n146 ) , .ZN( u2_u13_u3_n147 ) );
  AND2_X1 u2_u13_u3_U80 (.A1( u2_u13_X_19 ) , .ZN( u2_u13_u3_n102 ) , .A2( u2_u13_u3_n172 ) );
  AND2_X1 u2_u13_u3_U81 (.A1( u2_u13_X_21 ) , .A2( u2_u13_X_24 ) , .ZN( u2_u13_u3_n100 ) );
  AND2_X1 u2_u13_u3_U82 (.A2( u2_u13_X_19 ) , .A1( u2_u13_X_20 ) , .ZN( u2_u13_u3_n104 ) );
  INV_X1 u2_u13_u3_U83 (.A( u2_u13_X_22 ) , .ZN( u2_u13_u3_n166 ) );
  INV_X1 u2_u13_u3_U84 (.A( u2_u13_X_21 ) , .ZN( u2_u13_u3_n171 ) );
  INV_X1 u2_u13_u3_U85 (.A( u2_u13_X_20 ) , .ZN( u2_u13_u3_n172 ) );
  NAND4_X1 u2_u13_u3_U86 (.ZN( u2_out13_26 ) , .A4( u2_u13_u3_n109 ) , .A3( u2_u13_u3_n110 ) , .A2( u2_u13_u3_n111 ) , .A1( u2_u13_u3_n173 ) );
  INV_X1 u2_u13_u3_U87 (.ZN( u2_u13_u3_n173 ) , .A( u2_u13_u3_n94 ) );
  OAI21_X1 u2_u13_u3_U88 (.ZN( u2_u13_u3_n111 ) , .B2( u2_u13_u3_n117 ) , .A( u2_u13_u3_n133 ) , .B1( u2_u13_u3_n176 ) );
  NAND4_X1 u2_u13_u3_U89 (.ZN( u2_out13_20 ) , .A4( u2_u13_u3_n122 ) , .A3( u2_u13_u3_n123 ) , .A1( u2_u13_u3_n175 ) , .A2( u2_u13_u3_n180 ) );
  INV_X1 u2_u13_u3_U9 (.A( u2_u13_u3_n143 ) , .ZN( u2_u13_u3_n168 ) );
  INV_X1 u2_u13_u3_U90 (.A( u2_u13_u3_n112 ) , .ZN( u2_u13_u3_n175 ) );
  INV_X1 u2_u13_u3_U91 (.A( u2_u13_u3_n126 ) , .ZN( u2_u13_u3_n180 ) );
  NAND4_X1 u2_u13_u3_U92 (.ZN( u2_out13_1 ) , .A4( u2_u13_u3_n161 ) , .A3( u2_u13_u3_n162 ) , .A2( u2_u13_u3_n163 ) , .A1( u2_u13_u3_n185 ) );
  NAND2_X1 u2_u13_u3_U93 (.ZN( u2_u13_u3_n163 ) , .A2( u2_u13_u3_n170 ) , .A1( u2_u13_u3_n176 ) );
  AOI22_X1 u2_u13_u3_U94 (.B2( u2_u13_u3_n140 ) , .B1( u2_u13_u3_n141 ) , .A2( u2_u13_u3_n142 ) , .ZN( u2_u13_u3_n162 ) , .A1( u2_u13_u3_n177 ) );
  OR4_X1 u2_u13_u3_U95 (.ZN( u2_out13_10 ) , .A4( u2_u13_u3_n136 ) , .A3( u2_u13_u3_n137 ) , .A1( u2_u13_u3_n138 ) , .A2( u2_u13_u3_n139 ) );
  OAI222_X1 u2_u13_u3_U96 (.C1( u2_u13_u3_n128 ) , .ZN( u2_u13_u3_n137 ) , .B1( u2_u13_u3_n148 ) , .A2( u2_u13_u3_n150 ) , .B2( u2_u13_u3_n154 ) , .C2( u2_u13_u3_n164 ) , .A1( u2_u13_u3_n167 ) );
  OAI221_X1 u2_u13_u3_U97 (.A( u2_u13_u3_n134 ) , .B2( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n136 ) , .C1( u2_u13_u3_n149 ) , .B1( u2_u13_u3_n151 ) , .C2( u2_u13_u3_n183 ) );
  NAND3_X1 u2_u13_u3_U98 (.A1( u2_u13_u3_n114 ) , .ZN( u2_u13_u3_n115 ) , .A2( u2_u13_u3_n145 ) , .A3( u2_u13_u3_n153 ) );
  NAND3_X1 u2_u13_u3_U99 (.ZN( u2_u13_u3_n129 ) , .A2( u2_u13_u3_n144 ) , .A1( u2_u13_u3_n153 ) , .A3( u2_u13_u3_n182 ) );
  XOR2_X1 u2_u14_U1 (.B( u2_K15_9 ) , .A( u2_R13_6 ) , .Z( u2_u14_X_9 ) );
  XOR2_X1 u2_u14_U10 (.B( u2_K15_45 ) , .A( u2_R13_30 ) , .Z( u2_u14_X_45 ) );
  XOR2_X1 u2_u14_U12 (.B( u2_K15_43 ) , .A( u2_R13_28 ) , .Z( u2_u14_X_43 ) );
  XOR2_X1 u2_u14_U14 (.B( u2_K15_41 ) , .A( u2_R13_28 ) , .Z( u2_u14_X_41 ) );
  XOR2_X1 u2_u14_U16 (.B( u2_K15_3 ) , .A( u2_R13_2 ) , .Z( u2_u14_X_3 ) );
  XOR2_X1 u2_u14_U17 (.B( u2_K15_39 ) , .A( u2_R13_26 ) , .Z( u2_u14_X_39 ) );
  XOR2_X1 u2_u14_U22 (.B( u2_K15_34 ) , .A( u2_R13_23 ) , .Z( u2_u14_X_34 ) );
  XOR2_X1 u2_u14_U24 (.B( u2_K15_32 ) , .A( u2_R13_21 ) , .Z( u2_u14_X_32 ) );
  XOR2_X1 u2_u14_U26 (.B( u2_K15_30 ) , .A( u2_R13_21 ) , .Z( u2_u14_X_30 ) );
  XOR2_X1 u2_u14_U29 (.B( u2_K15_28 ) , .A( u2_R13_19 ) , .Z( u2_u14_X_28 ) );
  XOR2_X1 u2_u14_U3 (.B( u2_K15_7 ) , .A( u2_R13_4 ) , .Z( u2_u14_X_7 ) );
  XOR2_X1 u2_u14_U30 (.B( u2_K15_27 ) , .A( u2_R13_18 ) , .Z( u2_u14_X_27 ) );
  XOR2_X1 u2_u14_U35 (.B( u2_K15_22 ) , .A( u2_R13_15 ) , .Z( u2_u14_X_22 ) );
  XOR2_X1 u2_u14_U36 (.B( u2_K15_21 ) , .A( u2_R13_14 ) , .Z( u2_u14_X_21 ) );
  XOR2_X1 u2_u14_U37 (.B( u2_K15_20 ) , .A( u2_R13_13 ) , .Z( u2_u14_X_20 ) );
  XOR2_X1 u2_u14_U40 (.B( u2_K15_18 ) , .A( u2_R13_13 ) , .Z( u2_u14_X_18 ) );
  XOR2_X1 u2_u14_U42 (.B( u2_K15_16 ) , .A( u2_R13_11 ) , .Z( u2_u14_X_16 ) );
  XOR2_X1 u2_u14_U43 (.B( u2_K15_15 ) , .A( u2_R13_10 ) , .Z( u2_u14_X_15 ) );
  XOR2_X1 u2_u14_U45 (.B( u2_K15_13 ) , .A( u2_R13_8 ) , .Z( u2_u14_X_13 ) );
  XOR2_X1 u2_u14_U47 (.B( u2_K15_11 ) , .A( u2_R13_8 ) , .Z( u2_u14_X_11 ) );
  XOR2_X1 u2_u14_U48 (.B( u2_K15_10 ) , .A( u2_R13_7 ) , .Z( u2_u14_X_10 ) );
  XOR2_X1 u2_u14_U5 (.B( u2_K15_5 ) , .A( u2_R13_4 ) , .Z( u2_u14_X_5 ) );
  XOR2_X1 u2_u14_U6 (.B( u2_K15_4 ) , .A( u2_R13_3 ) , .Z( u2_u14_X_4 ) );
  XOR2_X1 u2_u14_U9 (.B( u2_K15_46 ) , .A( u2_R13_31 ) , .Z( u2_u14_X_46 ) );
  XOR2_X1 u2_u15_U1 (.A( u2_FP_38 ) , .B( u2_K16_9 ) , .Z( u2_u15_X_9 ) );
  XOR2_X1 u2_u15_U10 (.A( u2_FP_62 ) , .B( u2_K16_45 ) , .Z( u2_u15_X_45 ) );
  XOR2_X1 u2_u15_U15 (.A( u2_FP_59 ) , .B( u2_K16_40 ) , .Z( u2_u15_X_40 ) );
  XOR2_X1 u2_u15_U16 (.A( u2_FP_34 ) , .B( u2_K16_3 ) , .Z( u2_u15_X_3 ) );
  XOR2_X1 u2_u15_U17 (.A( u2_FP_58 ) , .B( u2_K16_39 ) , .Z( u2_u15_X_39 ) );
  XOR2_X1 u2_u15_U23 (.A( u2_FP_54 ) , .B( u2_K16_33 ) , .Z( u2_u15_X_33 ) );
  XOR2_X1 u2_u15_U29 (.A( u2_FP_51 ) , .B( u2_K16_28 ) , .Z( u2_u15_X_28 ) );
  XOR2_X1 u2_u15_U30 (.A( u2_FP_50 ) , .B( u2_K16_27 ) , .Z( u2_u15_X_27 ) );
  XOR2_X1 u2_u15_U35 (.A( u2_FP_47 ) , .B( u2_K16_22 ) , .Z( u2_u15_X_22 ) );
  XOR2_X1 u2_u15_U36 (.A( u2_FP_46 ) , .B( u2_K16_21 ) , .Z( u2_u15_X_21 ) );
  XOR2_X1 u2_u15_U42 (.A( u2_FP_43 ) , .B( u2_K16_16 ) , .Z( u2_u15_X_16 ) );
  XOR2_X1 u2_u15_U43 (.A( u2_FP_42 ) , .B( u2_K16_15 ) , .Z( u2_u15_X_15 ) );
  XOR2_X1 u2_u15_U48 (.A( u2_FP_39 ) , .B( u2_K16_10 ) , .Z( u2_u15_X_10 ) );
  XOR2_X1 u2_u15_U6 (.A( u2_FP_35 ) , .B( u2_K16_4 ) , .Z( u2_u15_X_4 ) );
  XOR2_X1 u2_u15_U9 (.A( u2_FP_63 ) , .B( u2_K16_46 ) , .Z( u2_u15_X_46 ) );
  XOR2_X1 u2_u1_U1 (.B( u2_K2_9 ) , .A( u2_R0_6 ) , .Z( u2_u1_X_9 ) );
  XOR2_X1 u2_u1_U10 (.B( u2_K2_45 ) , .A( u2_R0_30 ) , .Z( u2_u1_X_45 ) );
  XOR2_X1 u2_u1_U12 (.B( u2_K2_43 ) , .A( u2_R0_28 ) , .Z( u2_u1_X_43 ) );
  XOR2_X1 u2_u1_U14 (.B( u2_K2_41 ) , .A( u2_R0_28 ) , .Z( u2_u1_X_41 ) );
  XOR2_X1 u2_u1_U15 (.B( u2_K2_40 ) , .A( u2_R0_27 ) , .Z( u2_u1_X_40 ) );
  XOR2_X1 u2_u1_U16 (.B( u2_K2_3 ) , .A( u2_R0_2 ) , .Z( u2_u1_X_3 ) );
  XOR2_X1 u2_u1_U17 (.B( u2_K2_39 ) , .A( u2_R0_26 ) , .Z( u2_u1_X_39 ) );
  XOR2_X1 u2_u1_U22 (.B( u2_K2_34 ) , .A( u2_R0_23 ) , .Z( u2_u1_X_34 ) );
  XOR2_X1 u2_u1_U23 (.B( u2_K2_33 ) , .A( u2_R0_22 ) , .Z( u2_u1_X_33 ) );
  XOR2_X1 u2_u1_U30 (.B( u2_K2_27 ) , .A( u2_R0_18 ) , .Z( u2_u1_X_27 ) );
  XOR2_X1 u2_u1_U35 (.B( u2_K2_22 ) , .A( u2_R0_15 ) , .Z( u2_u1_X_22 ) );
  XOR2_X1 u2_u1_U36 (.B( u2_K2_21 ) , .A( u2_R0_14 ) , .Z( u2_u1_X_21 ) );
  XOR2_X1 u2_u1_U42 (.B( u2_K2_16 ) , .A( u2_R0_11 ) , .Z( u2_u1_X_16 ) );
  XOR2_X1 u2_u1_U43 (.B( u2_K2_15 ) , .A( u2_R0_10 ) , .Z( u2_u1_X_15 ) );
  XOR2_X1 u2_u1_U6 (.B( u2_K2_4 ) , .A( u2_R0_3 ) , .Z( u2_u1_X_4 ) );
  XOR2_X1 u2_u1_U9 (.B( u2_K2_46 ) , .A( u2_R0_31 ) , .Z( u2_u1_X_46 ) );
  XOR2_X1 u2_u2_U17 (.B( u2_K3_39 ) , .A( u2_R1_26 ) , .Z( u2_u2_X_39 ) );
  XOR2_X1 u2_u2_U19 (.B( u2_K3_37 ) , .A( u2_R1_24 ) , .Z( u2_u2_X_37 ) );
  XOR2_X1 u2_u2_U21 (.B( u2_K3_35 ) , .A( u2_R1_24 ) , .Z( u2_u2_X_35 ) );
  XOR2_X1 u2_u2_U22 (.B( u2_K3_34 ) , .A( u2_R1_23 ) , .Z( u2_u2_X_34 ) );
  XOR2_X1 u2_u2_U23 (.B( u2_K3_33 ) , .A( u2_R1_22 ) , .Z( u2_u2_X_33 ) );
  XOR2_X1 u2_u2_U24 (.B( u2_K3_32 ) , .A( u2_R1_21 ) , .Z( u2_u2_X_32 ) );
  XOR2_X1 u2_u2_U25 (.B( u2_K3_31 ) , .A( u2_R1_20 ) , .Z( u2_u2_X_31 ) );
  XOR2_X1 u2_u2_U26 (.B( u2_K3_30 ) , .A( u2_R1_21 ) , .Z( u2_u2_X_30 ) );
  XOR2_X1 u2_u2_U28 (.B( u2_K3_29 ) , .A( u2_R1_20 ) , .Z( u2_u2_X_29 ) );
  XOR2_X1 u2_u2_U29 (.B( u2_K3_28 ) , .A( u2_R1_19 ) , .Z( u2_u2_X_28 ) );
  XOR2_X1 u2_u2_U3 (.B( u2_K3_7 ) , .A( u2_R1_4 ) , .Z( u2_u2_X_7 ) );
  XOR2_X1 u2_u2_U30 (.B( u2_K3_27 ) , .A( u2_R1_18 ) , .Z( u2_u2_X_27 ) );
  XOR2_X1 u2_u2_U42 (.B( u2_K3_16 ) , .A( u2_R1_11 ) , .Z( u2_u2_X_16 ) );
  XOR2_X1 u2_u2_U43 (.B( u2_K3_15 ) , .A( u2_R1_10 ) , .Z( u2_u2_X_15 ) );
  XOR2_X1 u2_u2_U5 (.B( u2_K3_5 ) , .A( u2_R1_4 ) , .Z( u2_u2_X_5 ) );
  XOR2_X1 u2_u3_U10 (.B( u2_K4_45 ) , .A( u2_R2_30 ) , .Z( u2_u3_X_45 ) );
  XOR2_X1 u2_u3_U11 (.B( u2_K4_44 ) , .A( u2_R2_29 ) , .Z( u2_u3_X_44 ) );
  XOR2_X1 u2_u3_U12 (.B( u2_K4_43 ) , .A( u2_R2_28 ) , .Z( u2_u3_X_43 ) );
  XOR2_X1 u2_u3_U13 (.B( u2_K4_42 ) , .A( u2_R2_29 ) , .Z( u2_u3_X_42 ) );
  XOR2_X1 u2_u3_U14 (.B( u2_K4_41 ) , .A( u2_R2_28 ) , .Z( u2_u3_X_41 ) );
  XOR2_X1 u2_u3_U15 (.B( u2_K4_40 ) , .A( u2_R2_27 ) , .Z( u2_u3_X_40 ) );
  XOR2_X1 u2_u3_U17 (.B( u2_K4_39 ) , .A( u2_R2_26 ) , .Z( u2_u3_X_39 ) );
  XOR2_X1 u2_u3_U18 (.B( u2_K4_38 ) , .A( u2_R2_25 ) , .Z( u2_u3_X_38 ) );
  XOR2_X1 u2_u3_U19 (.B( u2_K4_37 ) , .A( u2_R2_24 ) , .Z( u2_u3_X_37 ) );
  XOR2_X1 u2_u3_U21 (.B( u2_K4_35 ) , .A( u2_R2_24 ) , .Z( u2_u3_X_35 ) );
  XOR2_X1 u2_u3_U22 (.B( u2_K4_34 ) , .A( u2_R2_23 ) , .Z( u2_u3_X_34 ) );
  XOR2_X1 u2_u3_U23 (.B( u2_K4_33 ) , .A( u2_R2_22 ) , .Z( u2_u3_X_33 ) );
  XOR2_X1 u2_u3_U30 (.B( u2_K4_27 ) , .A( u2_R2_18 ) , .Z( u2_u3_X_27 ) );
  XOR2_X1 u2_u3_U35 (.B( u2_K4_22 ) , .A( u2_R2_15 ) , .Z( u2_u3_X_22 ) );
  XOR2_X1 u2_u3_U36 (.B( u2_K4_21 ) , .A( u2_R2_14 ) , .Z( u2_u3_X_21 ) );
  XOR2_X1 u2_u3_U9 (.B( u2_K4_46 ) , .A( u2_R2_31 ) , .Z( u2_u3_X_46 ) );
  INV_X1 u2_u3_u6_U10 (.ZN( u2_u3_u6_n172 ) , .A( u2_u3_u6_n88 ) );
  OAI21_X1 u2_u3_u6_U11 (.A( u2_u3_u6_n159 ) , .B1( u2_u3_u6_n169 ) , .B2( u2_u3_u6_n173 ) , .ZN( u2_u3_u6_n90 ) );
  AOI22_X1 u2_u3_u6_U12 (.A2( u2_u3_u6_n151 ) , .B2( u2_u3_u6_n161 ) , .A1( u2_u3_u6_n167 ) , .B1( u2_u3_u6_n170 ) , .ZN( u2_u3_u6_n89 ) );
  AOI21_X1 u2_u3_u6_U13 (.ZN( u2_u3_u6_n106 ) , .A( u2_u3_u6_n142 ) , .B2( u2_u3_u6_n159 ) , .B1( u2_u3_u6_n164 ) );
  INV_X1 u2_u3_u6_U14 (.A( u2_u3_u6_n155 ) , .ZN( u2_u3_u6_n161 ) );
  INV_X1 u2_u3_u6_U15 (.A( u2_u3_u6_n128 ) , .ZN( u2_u3_u6_n164 ) );
  NAND2_X1 u2_u3_u6_U16 (.ZN( u2_u3_u6_n110 ) , .A1( u2_u3_u6_n122 ) , .A2( u2_u3_u6_n129 ) );
  NAND2_X1 u2_u3_u6_U17 (.ZN( u2_u3_u6_n124 ) , .A2( u2_u3_u6_n146 ) , .A1( u2_u3_u6_n148 ) );
  INV_X1 u2_u3_u6_U18 (.A( u2_u3_u6_n132 ) , .ZN( u2_u3_u6_n171 ) );
  AND2_X1 u2_u3_u6_U19 (.A1( u2_u3_u6_n100 ) , .ZN( u2_u3_u6_n130 ) , .A2( u2_u3_u6_n147 ) );
  INV_X1 u2_u3_u6_U20 (.A( u2_u3_u6_n127 ) , .ZN( u2_u3_u6_n173 ) );
  INV_X1 u2_u3_u6_U21 (.A( u2_u3_u6_n121 ) , .ZN( u2_u3_u6_n167 ) );
  INV_X1 u2_u3_u6_U22 (.A( u2_u3_u6_n100 ) , .ZN( u2_u3_u6_n169 ) );
  INV_X1 u2_u3_u6_U23 (.A( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n170 ) );
  INV_X1 u2_u3_u6_U24 (.A( u2_u3_u6_n113 ) , .ZN( u2_u3_u6_n168 ) );
  AND2_X1 u2_u3_u6_U25 (.A1( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n119 ) , .ZN( u2_u3_u6_n133 ) );
  AND2_X1 u2_u3_u6_U26 (.A2( u2_u3_u6_n121 ) , .A1( u2_u3_u6_n122 ) , .ZN( u2_u3_u6_n131 ) );
  AND3_X1 u2_u3_u6_U27 (.ZN( u2_u3_u6_n120 ) , .A2( u2_u3_u6_n127 ) , .A1( u2_u3_u6_n132 ) , .A3( u2_u3_u6_n145 ) );
  INV_X1 u2_u3_u6_U28 (.A( u2_u3_u6_n146 ) , .ZN( u2_u3_u6_n163 ) );
  AOI222_X1 u2_u3_u6_U29 (.ZN( u2_u3_u6_n114 ) , .A1( u2_u3_u6_n118 ) , .A2( u2_u3_u6_n126 ) , .B2( u2_u3_u6_n151 ) , .C2( u2_u3_u6_n159 ) , .C1( u2_u3_u6_n168 ) , .B1( u2_u3_u6_n169 ) );
  INV_X1 u2_u3_u6_U3 (.A( u2_u3_u6_n110 ) , .ZN( u2_u3_u6_n166 ) );
  NOR2_X1 u2_u3_u6_U30 (.A1( u2_u3_u6_n162 ) , .A2( u2_u3_u6_n165 ) , .ZN( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U31 (.A1( u2_u3_u6_n144 ) , .ZN( u2_u3_u6_n151 ) , .A2( u2_u3_u6_n158 ) );
  NAND2_X1 u2_u3_u6_U32 (.ZN( u2_u3_u6_n132 ) , .A1( u2_u3_u6_n91 ) , .A2( u2_u3_u6_n97 ) );
  AOI22_X1 u2_u3_u6_U33 (.B2( u2_u3_u6_n110 ) , .B1( u2_u3_u6_n111 ) , .A1( u2_u3_u6_n112 ) , .ZN( u2_u3_u6_n115 ) , .A2( u2_u3_u6_n161 ) );
  NAND4_X1 u2_u3_u6_U34 (.A3( u2_u3_u6_n109 ) , .ZN( u2_u3_u6_n112 ) , .A4( u2_u3_u6_n132 ) , .A2( u2_u3_u6_n147 ) , .A1( u2_u3_u6_n166 ) );
  NOR2_X1 u2_u3_u6_U35 (.ZN( u2_u3_u6_n109 ) , .A1( u2_u3_u6_n170 ) , .A2( u2_u3_u6_n173 ) );
  NOR2_X1 u2_u3_u6_U36 (.A2( u2_u3_u6_n126 ) , .ZN( u2_u3_u6_n155 ) , .A1( u2_u3_u6_n160 ) );
  NAND2_X1 u2_u3_u6_U37 (.ZN( u2_u3_u6_n146 ) , .A2( u2_u3_u6_n94 ) , .A1( u2_u3_u6_n99 ) );
  AOI21_X1 u2_u3_u6_U38 (.A( u2_u3_u6_n144 ) , .B2( u2_u3_u6_n145 ) , .B1( u2_u3_u6_n146 ) , .ZN( u2_u3_u6_n150 ) );
  AOI211_X1 u2_u3_u6_U39 (.B( u2_u3_u6_n134 ) , .A( u2_u3_u6_n135 ) , .C1( u2_u3_u6_n136 ) , .ZN( u2_u3_u6_n137 ) , .C2( u2_u3_u6_n151 ) );
  INV_X1 u2_u3_u6_U4 (.A( u2_u3_u6_n142 ) , .ZN( u2_u3_u6_n174 ) );
  AOI21_X1 u2_u3_u6_U40 (.B2( u2_u3_u6_n132 ) , .B1( u2_u3_u6_n133 ) , .ZN( u2_u3_u6_n134 ) , .A( u2_u3_u6_n158 ) );
  NAND4_X1 u2_u3_u6_U41 (.A4( u2_u3_u6_n127 ) , .A3( u2_u3_u6_n128 ) , .A2( u2_u3_u6_n129 ) , .A1( u2_u3_u6_n130 ) , .ZN( u2_u3_u6_n136 ) );
  AOI21_X1 u2_u3_u6_U42 (.B1( u2_u3_u6_n131 ) , .ZN( u2_u3_u6_n135 ) , .A( u2_u3_u6_n144 ) , .B2( u2_u3_u6_n146 ) );
  INV_X1 u2_u3_u6_U43 (.A( u2_u3_u6_n111 ) , .ZN( u2_u3_u6_n158 ) );
  NAND2_X1 u2_u3_u6_U44 (.ZN( u2_u3_u6_n127 ) , .A1( u2_u3_u6_n91 ) , .A2( u2_u3_u6_n92 ) );
  NAND2_X1 u2_u3_u6_U45 (.ZN( u2_u3_u6_n129 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n96 ) );
  INV_X1 u2_u3_u6_U46 (.A( u2_u3_u6_n144 ) , .ZN( u2_u3_u6_n159 ) );
  NAND2_X1 u2_u3_u6_U47 (.ZN( u2_u3_u6_n145 ) , .A2( u2_u3_u6_n97 ) , .A1( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U48 (.ZN( u2_u3_u6_n148 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n94 ) );
  NAND2_X1 u2_u3_u6_U49 (.ZN( u2_u3_u6_n108 ) , .A2( u2_u3_u6_n139 ) , .A1( u2_u3_u6_n144 ) );
  NAND2_X1 u2_u3_u6_U5 (.A2( u2_u3_u6_n143 ) , .ZN( u2_u3_u6_n152 ) , .A1( u2_u3_u6_n166 ) );
  NAND2_X1 u2_u3_u6_U50 (.ZN( u2_u3_u6_n121 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n97 ) );
  NAND2_X1 u2_u3_u6_U51 (.ZN( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n95 ) );
  AND2_X1 u2_u3_u6_U52 (.ZN( u2_u3_u6_n118 ) , .A2( u2_u3_u6_n91 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U53 (.ZN( u2_u3_u6_n147 ) , .A2( u2_u3_u6_n98 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U54 (.ZN( u2_u3_u6_n128 ) , .A1( u2_u3_u6_n94 ) , .A2( u2_u3_u6_n96 ) );
  NAND2_X1 u2_u3_u6_U55 (.ZN( u2_u3_u6_n119 ) , .A2( u2_u3_u6_n95 ) , .A1( u2_u3_u6_n99 ) );
  NAND2_X1 u2_u3_u6_U56 (.ZN( u2_u3_u6_n123 ) , .A2( u2_u3_u6_n91 ) , .A1( u2_u3_u6_n96 ) );
  NAND2_X1 u2_u3_u6_U57 (.ZN( u2_u3_u6_n100 ) , .A2( u2_u3_u6_n92 ) , .A1( u2_u3_u6_n98 ) );
  NAND2_X1 u2_u3_u6_U58 (.ZN( u2_u3_u6_n122 ) , .A1( u2_u3_u6_n94 ) , .A2( u2_u3_u6_n97 ) );
  INV_X1 u2_u3_u6_U59 (.A( u2_u3_u6_n139 ) , .ZN( u2_u3_u6_n160 ) );
  AOI22_X1 u2_u3_u6_U6 (.B2( u2_u3_u6_n101 ) , .A1( u2_u3_u6_n102 ) , .ZN( u2_u3_u6_n103 ) , .B1( u2_u3_u6_n160 ) , .A2( u2_u3_u6_n161 ) );
  NAND2_X1 u2_u3_u6_U60 (.ZN( u2_u3_u6_n113 ) , .A1( u2_u3_u6_n96 ) , .A2( u2_u3_u6_n98 ) );
  NOR2_X1 u2_u3_u6_U61 (.A2( u2_u3_X_40 ) , .A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n126 ) );
  NOR2_X1 u2_u3_u6_U62 (.A2( u2_u3_X_39 ) , .A1( u2_u3_X_42 ) , .ZN( u2_u3_u6_n92 ) );
  NOR2_X1 u2_u3_u6_U63 (.A2( u2_u3_X_39 ) , .A1( u2_u3_u6_n156 ) , .ZN( u2_u3_u6_n97 ) );
  NOR2_X1 u2_u3_u6_U64 (.A2( u2_u3_X_38 ) , .A1( u2_u3_u6_n165 ) , .ZN( u2_u3_u6_n95 ) );
  NOR2_X1 u2_u3_u6_U65 (.A2( u2_u3_X_41 ) , .ZN( u2_u3_u6_n111 ) , .A1( u2_u3_u6_n157 ) );
  NOR2_X1 u2_u3_u6_U66 (.A2( u2_u3_X_37 ) , .A1( u2_u3_u6_n162 ) , .ZN( u2_u3_u6_n94 ) );
  NOR2_X1 u2_u3_u6_U67 (.A2( u2_u3_X_37 ) , .A1( u2_u3_X_38 ) , .ZN( u2_u3_u6_n91 ) );
  NAND2_X1 u2_u3_u6_U68 (.A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n144 ) , .A2( u2_u3_u6_n157 ) );
  NAND2_X1 u2_u3_u6_U69 (.A2( u2_u3_X_40 ) , .A1( u2_u3_X_41 ) , .ZN( u2_u3_u6_n139 ) );
  NOR2_X1 u2_u3_u6_U7 (.A1( u2_u3_u6_n118 ) , .ZN( u2_u3_u6_n143 ) , .A2( u2_u3_u6_n168 ) );
  AND2_X1 u2_u3_u6_U70 (.A1( u2_u3_X_39 ) , .A2( u2_u3_u6_n156 ) , .ZN( u2_u3_u6_n96 ) );
  AND2_X1 u2_u3_u6_U71 (.A1( u2_u3_X_39 ) , .A2( u2_u3_X_42 ) , .ZN( u2_u3_u6_n99 ) );
  INV_X1 u2_u3_u6_U72 (.A( u2_u3_X_40 ) , .ZN( u2_u3_u6_n157 ) );
  INV_X1 u2_u3_u6_U73 (.A( u2_u3_X_37 ) , .ZN( u2_u3_u6_n165 ) );
  INV_X1 u2_u3_u6_U74 (.A( u2_u3_X_38 ) , .ZN( u2_u3_u6_n162 ) );
  INV_X1 u2_u3_u6_U75 (.A( u2_u3_X_42 ) , .ZN( u2_u3_u6_n156 ) );
  NAND4_X1 u2_u3_u6_U76 (.ZN( u2_out3_32 ) , .A4( u2_u3_u6_n103 ) , .A3( u2_u3_u6_n104 ) , .A2( u2_u3_u6_n105 ) , .A1( u2_u3_u6_n106 ) );
  AOI22_X1 u2_u3_u6_U77 (.ZN( u2_u3_u6_n105 ) , .A2( u2_u3_u6_n108 ) , .A1( u2_u3_u6_n118 ) , .B2( u2_u3_u6_n126 ) , .B1( u2_u3_u6_n171 ) );
  AOI22_X1 u2_u3_u6_U78 (.ZN( u2_u3_u6_n104 ) , .A1( u2_u3_u6_n111 ) , .B1( u2_u3_u6_n124 ) , .B2( u2_u3_u6_n151 ) , .A2( u2_u3_u6_n93 ) );
  NAND4_X1 u2_u3_u6_U79 (.ZN( u2_out3_12 ) , .A4( u2_u3_u6_n114 ) , .A3( u2_u3_u6_n115 ) , .A2( u2_u3_u6_n116 ) , .A1( u2_u3_u6_n117 ) );
  AOI21_X1 u2_u3_u6_U8 (.B1( u2_u3_u6_n107 ) , .B2( u2_u3_u6_n132 ) , .A( u2_u3_u6_n158 ) , .ZN( u2_u3_u6_n88 ) );
  OAI22_X1 u2_u3_u6_U80 (.B2( u2_u3_u6_n111 ) , .ZN( u2_u3_u6_n116 ) , .B1( u2_u3_u6_n126 ) , .A2( u2_u3_u6_n164 ) , .A1( u2_u3_u6_n167 ) );
  OAI21_X1 u2_u3_u6_U81 (.A( u2_u3_u6_n108 ) , .ZN( u2_u3_u6_n117 ) , .B2( u2_u3_u6_n141 ) , .B1( u2_u3_u6_n163 ) );
  OAI211_X1 u2_u3_u6_U82 (.ZN( u2_out3_22 ) , .B( u2_u3_u6_n137 ) , .A( u2_u3_u6_n138 ) , .C2( u2_u3_u6_n139 ) , .C1( u2_u3_u6_n140 ) );
  AOI22_X1 u2_u3_u6_U83 (.B1( u2_u3_u6_n124 ) , .A2( u2_u3_u6_n125 ) , .A1( u2_u3_u6_n126 ) , .ZN( u2_u3_u6_n138 ) , .B2( u2_u3_u6_n161 ) );
  AND4_X1 u2_u3_u6_U84 (.A3( u2_u3_u6_n119 ) , .A1( u2_u3_u6_n120 ) , .A4( u2_u3_u6_n129 ) , .ZN( u2_u3_u6_n140 ) , .A2( u2_u3_u6_n143 ) );
  OAI211_X1 u2_u3_u6_U85 (.ZN( u2_out3_7 ) , .B( u2_u3_u6_n153 ) , .C2( u2_u3_u6_n154 ) , .C1( u2_u3_u6_n155 ) , .A( u2_u3_u6_n174 ) );
  NOR3_X1 u2_u3_u6_U86 (.A1( u2_u3_u6_n141 ) , .ZN( u2_u3_u6_n154 ) , .A3( u2_u3_u6_n164 ) , .A2( u2_u3_u6_n171 ) );
  AOI211_X1 u2_u3_u6_U87 (.B( u2_u3_u6_n149 ) , .A( u2_u3_u6_n150 ) , .C2( u2_u3_u6_n151 ) , .C1( u2_u3_u6_n152 ) , .ZN( u2_u3_u6_n153 ) );
  NAND3_X1 u2_u3_u6_U88 (.A2( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n125 ) , .A1( u2_u3_u6_n130 ) , .A3( u2_u3_u6_n131 ) );
  NAND3_X1 u2_u3_u6_U89 (.A3( u2_u3_u6_n133 ) , .ZN( u2_u3_u6_n141 ) , .A1( u2_u3_u6_n145 ) , .A2( u2_u3_u6_n148 ) );
  AOI21_X1 u2_u3_u6_U9 (.B2( u2_u3_u6_n147 ) , .B1( u2_u3_u6_n148 ) , .ZN( u2_u3_u6_n149 ) , .A( u2_u3_u6_n158 ) );
  NAND3_X1 u2_u3_u6_U90 (.ZN( u2_u3_u6_n101 ) , .A3( u2_u3_u6_n107 ) , .A2( u2_u3_u6_n121 ) , .A1( u2_u3_u6_n127 ) );
  NAND3_X1 u2_u3_u6_U91 (.ZN( u2_u3_u6_n102 ) , .A3( u2_u3_u6_n130 ) , .A2( u2_u3_u6_n145 ) , .A1( u2_u3_u6_n166 ) );
  NAND3_X1 u2_u3_u6_U92 (.A3( u2_u3_u6_n113 ) , .A1( u2_u3_u6_n119 ) , .A2( u2_u3_u6_n123 ) , .ZN( u2_u3_u6_n93 ) );
  NAND3_X1 u2_u3_u6_U93 (.ZN( u2_u3_u6_n142 ) , .A2( u2_u3_u6_n172 ) , .A3( u2_u3_u6_n89 ) , .A1( u2_u3_u6_n90 ) );
  XOR2_X1 u2_u4_U1 (.B( u2_K5_9 ) , .A( u2_R3_6 ) , .Z( u2_u4_X_9 ) );
  XOR2_X1 u2_u4_U15 (.B( u2_K5_40 ) , .A( u2_R3_27 ) , .Z( u2_u4_X_40 ) );
  XOR2_X1 u2_u4_U16 (.B( u2_K5_3 ) , .A( u2_R3_2 ) , .Z( u2_u4_X_3 ) );
  XOR2_X1 u2_u4_U17 (.B( u2_K5_39 ) , .A( u2_R3_26 ) , .Z( u2_u4_X_39 ) );
  XOR2_X1 u2_u4_U22 (.B( u2_K5_34 ) , .A( u2_R3_23 ) , .Z( u2_u4_X_34 ) );
  XOR2_X1 u2_u4_U29 (.B( u2_K5_28 ) , .A( u2_R3_19 ) , .Z( u2_u4_X_28 ) );
  XOR2_X1 u2_u4_U35 (.B( u2_K5_22 ) , .A( u2_R3_15 ) , .Z( u2_u4_X_22 ) );
  XOR2_X1 u2_u4_U36 (.B( u2_K5_21 ) , .A( u2_R3_14 ) , .Z( u2_u4_X_21 ) );
  XOR2_X1 u2_u4_U38 (.B( u2_K5_1 ) , .A( u2_R3_32 ) , .Z( u2_u4_X_1 ) );
  XOR2_X1 u2_u4_U42 (.B( u2_K5_16 ) , .A( u2_R3_11 ) , .Z( u2_u4_X_16 ) );
  XOR2_X1 u2_u4_U43 (.B( u2_K5_15 ) , .A( u2_R3_10 ) , .Z( u2_u4_X_15 ) );
  XOR2_X1 u2_u4_U48 (.B( u2_K5_10 ) , .A( u2_R3_7 ) , .Z( u2_u4_X_10 ) );
  XOR2_X1 u2_u4_U6 (.B( u2_K5_4 ) , .A( u2_R3_3 ) , .Z( u2_u4_X_4 ) );
  XOR2_X1 u2_u4_U8 (.B( u2_K5_47 ) , .A( u2_R3_32 ) , .Z( u2_u4_X_47 ) );
  XOR2_X1 u2_u4_U9 (.B( u2_K5_46 ) , .A( u2_R3_31 ) , .Z( u2_u4_X_46 ) );
  XOR2_X1 u2_u5_U10 (.B( u2_K6_45 ) , .A( u2_R4_30 ) , .Z( u2_u5_X_45 ) );
  XOR2_X1 u2_u5_U15 (.B( u2_K6_40 ) , .A( u2_R4_27 ) , .Z( u2_u5_X_40 ) );
  XOR2_X1 u2_u5_U16 (.B( u2_K6_3 ) , .A( u2_R4_2 ) , .Z( u2_u5_X_3 ) );
  XOR2_X1 u2_u5_U17 (.B( u2_K6_39 ) , .A( u2_R4_26 ) , .Z( u2_u5_X_39 ) );
  XOR2_X1 u2_u5_U18 (.B( u2_K6_38 ) , .A( u2_R4_25 ) , .Z( u2_u5_X_38 ) );
  XOR2_X1 u2_u5_U20 (.B( u2_K6_36 ) , .A( u2_R4_25 ) , .Z( u2_u5_X_36 ) );
  XOR2_X1 u2_u5_U22 (.B( u2_K6_34 ) , .A( u2_R4_23 ) , .Z( u2_u5_X_34 ) );
  XOR2_X1 u2_u5_U25 (.B( u2_K6_31 ) , .A( u2_R4_20 ) , .Z( u2_u5_X_31 ) );
  XOR2_X1 u2_u5_U28 (.B( u2_K6_29 ) , .A( u2_R4_20 ) , .Z( u2_u5_X_29 ) );
  XOR2_X1 u2_u5_U29 (.B( u2_K6_28 ) , .A( u2_R4_19 ) , .Z( u2_u5_X_28 ) );
  XOR2_X1 u2_u5_U30 (.B( u2_K6_27 ) , .A( u2_R4_18 ) , .Z( u2_u5_X_27 ) );
  XOR2_X1 u2_u5_U32 (.B( u2_K6_25 ) , .A( u2_R4_16 ) , .Z( u2_u5_X_25 ) );
  XOR2_X1 u2_u5_U34 (.B( u2_K6_23 ) , .A( u2_R4_16 ) , .Z( u2_u5_X_23 ) );
  XOR2_X1 u2_u5_U35 (.B( u2_K6_22 ) , .A( u2_R4_15 ) , .Z( u2_u5_X_22 ) );
  XOR2_X1 u2_u5_U42 (.B( u2_K6_16 ) , .A( u2_R4_11 ) , .Z( u2_u5_X_16 ) );
  XOR2_X1 u2_u5_U43 (.B( u2_K6_15 ) , .A( u2_R4_10 ) , .Z( u2_u5_X_15 ) );
  XOR2_X1 u2_u5_U48 (.B( u2_K6_10 ) , .A( u2_R4_7 ) , .Z( u2_u5_X_10 ) );
  XOR2_X1 u2_u5_U6 (.B( u2_K6_4 ) , .A( u2_R4_3 ) , .Z( u2_u5_X_4 ) );
  XOR2_X1 u2_u6_U1 (.B( u2_K7_9 ) , .A( u2_R5_6 ) , .Z( u2_u6_X_9 ) );
  XOR2_X1 u2_u6_U10 (.B( u2_K7_45 ) , .A( u2_R5_30 ) , .Z( u2_u6_X_45 ) );
  XOR2_X1 u2_u6_U15 (.B( u2_K7_40 ) , .A( u2_R5_27 ) , .Z( u2_u6_X_40 ) );
  XOR2_X1 u2_u6_U16 (.B( u2_K7_3 ) , .A( u2_R5_2 ) , .Z( u2_u6_X_3 ) );
  XOR2_X1 u2_u6_U23 (.B( u2_K7_33 ) , .A( u2_R5_22 ) , .Z( u2_u6_X_33 ) );
  XOR2_X1 u2_u6_U29 (.B( u2_K7_28 ) , .A( u2_R5_19 ) , .Z( u2_u6_X_28 ) );
  XOR2_X1 u2_u6_U30 (.B( u2_K7_27 ) , .A( u2_R5_18 ) , .Z( u2_u6_X_27 ) );
  XOR2_X1 u2_u6_U35 (.B( u2_K7_22 ) , .A( u2_R5_15 ) , .Z( u2_u6_X_22 ) );
  XOR2_X1 u2_u6_U48 (.B( u2_K7_10 ) , .A( u2_R5_7 ) , .Z( u2_u6_X_10 ) );
  XOR2_X1 u2_u6_U6 (.B( u2_K7_4 ) , .A( u2_R5_3 ) , .Z( u2_u6_X_4 ) );
  XOR2_X1 u2_u6_U9 (.B( u2_K7_46 ) , .A( u2_R5_31 ) , .Z( u2_u6_X_46 ) );
  XOR2_X1 u2_u7_U1 (.B( u2_K8_9 ) , .A( u2_R6_6 ) , .Z( u2_u7_X_9 ) );
  XOR2_X1 u2_u7_U10 (.B( u2_K8_45 ) , .A( u2_R6_30 ) , .Z( u2_u7_X_45 ) );
  XOR2_X1 u2_u7_U11 (.B( u2_K8_44 ) , .A( u2_R6_29 ) , .Z( u2_u7_X_44 ) );
  XOR2_X1 u2_u7_U13 (.B( u2_K8_42 ) , .A( u2_R6_29 ) , .Z( u2_u7_X_42 ) );
  XOR2_X1 u2_u7_U14 (.B( u2_K8_41 ) , .A( u2_R6_28 ) , .Z( u2_u7_X_41 ) );
  XOR2_X1 u2_u7_U15 (.B( u2_K8_40 ) , .A( u2_R6_27 ) , .Z( u2_u7_X_40 ) );
  XOR2_X1 u2_u7_U17 (.B( u2_K8_39 ) , .A( u2_R6_26 ) , .Z( u2_u7_X_39 ) );
  XOR2_X1 u2_u7_U18 (.B( u2_K8_38 ) , .A( u2_R6_25 ) , .Z( u2_u7_X_38 ) );
  XOR2_X1 u2_u7_U19 (.B( u2_K8_37 ) , .A( u2_R6_24 ) , .Z( u2_u7_X_37 ) );
  XOR2_X1 u2_u7_U20 (.B( u2_K8_36 ) , .A( u2_R6_25 ) , .Z( u2_u7_X_36 ) );
  XOR2_X1 u2_u7_U21 (.B( u2_K8_35 ) , .A( u2_R6_24 ) , .Z( u2_u7_X_35 ) );
  XOR2_X1 u2_u7_U22 (.B( u2_K8_34 ) , .A( u2_R6_23 ) , .Z( u2_u7_X_34 ) );
  XOR2_X1 u2_u7_U23 (.B( u2_K8_33 ) , .A( u2_R6_22 ) , .Z( u2_u7_X_33 ) );
  XOR2_X1 u2_u7_U24 (.B( u2_K8_32 ) , .A( u2_R6_21 ) , .Z( u2_u7_X_32 ) );
  XOR2_X1 u2_u7_U25 (.B( u2_K8_31 ) , .A( u2_R6_20 ) , .Z( u2_u7_X_31 ) );
  XOR2_X1 u2_u7_U26 (.B( u2_K8_30 ) , .A( u2_R6_21 ) , .Z( u2_u7_X_30 ) );
  XOR2_X1 u2_u7_U28 (.B( u2_K8_29 ) , .A( u2_R6_20 ) , .Z( u2_u7_X_29 ) );
  XOR2_X1 u2_u7_U29 (.B( u2_K8_28 ) , .A( u2_R6_19 ) , .Z( u2_u7_X_28 ) );
  XOR2_X1 u2_u7_U30 (.B( u2_K8_27 ) , .A( u2_R6_18 ) , .Z( u2_u7_X_27 ) );
  XOR2_X1 u2_u7_U31 (.B( u2_K8_26 ) , .A( u2_R6_17 ) , .Z( u2_u7_X_26 ) );
  XOR2_X1 u2_u7_U32 (.B( u2_K8_25 ) , .A( u2_R6_16 ) , .Z( u2_u7_X_25 ) );
  XOR2_X1 u2_u7_U33 (.B( u2_K8_24 ) , .A( u2_R6_17 ) , .Z( u2_u7_X_24 ) );
  XOR2_X1 u2_u7_U34 (.B( u2_K8_23 ) , .A( u2_R6_16 ) , .Z( u2_u7_X_23 ) );
  XOR2_X1 u2_u7_U35 (.B( u2_K8_22 ) , .A( u2_R6_15 ) , .Z( u2_u7_X_22 ) );
  XOR2_X1 u2_u7_U36 (.B( u2_K8_21 ) , .A( u2_R6_14 ) , .Z( u2_u7_X_21 ) );
  XOR2_X1 u2_u7_U42 (.B( u2_K8_16 ) , .A( u2_R6_11 ) , .Z( u2_u7_X_16 ) );
  XOR2_X1 u2_u7_U43 (.B( u2_K8_15 ) , .A( u2_R6_10 ) , .Z( u2_u7_X_15 ) );
  XOR2_X1 u2_u7_U48 (.B( u2_K8_10 ) , .A( u2_R6_7 ) , .Z( u2_u7_X_10 ) );
  XOR2_X1 u2_u7_U6 (.B( u2_K8_4 ) , .A( u2_R6_3 ) , .Z( u2_u7_X_4 ) );
  XOR2_X1 u2_u7_U9 (.B( u2_K8_46 ) , .A( u2_R6_31 ) , .Z( u2_u7_X_46 ) );
  OAI22_X1 u2_u7_u4_U10 (.B2( u2_u7_u4_n135 ) , .ZN( u2_u7_u4_n137 ) , .B1( u2_u7_u4_n153 ) , .A1( u2_u7_u4_n155 ) , .A2( u2_u7_u4_n171 ) );
  AND3_X1 u2_u7_u4_U11 (.A2( u2_u7_u4_n134 ) , .ZN( u2_u7_u4_n135 ) , .A3( u2_u7_u4_n145 ) , .A1( u2_u7_u4_n157 ) );
  OR3_X1 u2_u7_u4_U12 (.A3( u2_u7_u4_n114 ) , .A2( u2_u7_u4_n115 ) , .A1( u2_u7_u4_n116 ) , .ZN( u2_u7_u4_n136 ) );
  AOI21_X1 u2_u7_u4_U13 (.A( u2_u7_u4_n113 ) , .ZN( u2_u7_u4_n116 ) , .B2( u2_u7_u4_n173 ) , .B1( u2_u7_u4_n174 ) );
  AOI21_X1 u2_u7_u4_U14 (.ZN( u2_u7_u4_n115 ) , .B2( u2_u7_u4_n145 ) , .B1( u2_u7_u4_n146 ) , .A( u2_u7_u4_n156 ) );
  OAI22_X1 u2_u7_u4_U15 (.ZN( u2_u7_u4_n114 ) , .A2( u2_u7_u4_n121 ) , .B1( u2_u7_u4_n160 ) , .B2( u2_u7_u4_n170 ) , .A1( u2_u7_u4_n171 ) );
  NAND2_X1 u2_u7_u4_U16 (.ZN( u2_u7_u4_n132 ) , .A2( u2_u7_u4_n170 ) , .A1( u2_u7_u4_n173 ) );
  AOI21_X1 u2_u7_u4_U17 (.B2( u2_u7_u4_n160 ) , .B1( u2_u7_u4_n161 ) , .ZN( u2_u7_u4_n162 ) , .A( u2_u7_u4_n170 ) );
  AOI21_X1 u2_u7_u4_U18 (.ZN( u2_u7_u4_n107 ) , .B2( u2_u7_u4_n143 ) , .A( u2_u7_u4_n174 ) , .B1( u2_u7_u4_n184 ) );
  AOI21_X1 u2_u7_u4_U19 (.B2( u2_u7_u4_n158 ) , .B1( u2_u7_u4_n159 ) , .ZN( u2_u7_u4_n163 ) , .A( u2_u7_u4_n174 ) );
  AOI21_X1 u2_u7_u4_U20 (.A( u2_u7_u4_n153 ) , .B2( u2_u7_u4_n154 ) , .B1( u2_u7_u4_n155 ) , .ZN( u2_u7_u4_n165 ) );
  AOI21_X1 u2_u7_u4_U21 (.A( u2_u7_u4_n156 ) , .B2( u2_u7_u4_n157 ) , .ZN( u2_u7_u4_n164 ) , .B1( u2_u7_u4_n184 ) );
  INV_X1 u2_u7_u4_U22 (.A( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n170 ) );
  AND2_X1 u2_u7_u4_U23 (.A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n155 ) , .A1( u2_u7_u4_n160 ) );
  INV_X1 u2_u7_u4_U24 (.A( u2_u7_u4_n156 ) , .ZN( u2_u7_u4_n175 ) );
  NAND2_X1 u2_u7_u4_U25 (.A2( u2_u7_u4_n118 ) , .ZN( u2_u7_u4_n131 ) , .A1( u2_u7_u4_n147 ) );
  NAND2_X1 u2_u7_u4_U26 (.A1( u2_u7_u4_n119 ) , .A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n130 ) );
  NAND2_X1 u2_u7_u4_U27 (.ZN( u2_u7_u4_n117 ) , .A2( u2_u7_u4_n118 ) , .A1( u2_u7_u4_n148 ) );
  NAND2_X1 u2_u7_u4_U28 (.ZN( u2_u7_u4_n129 ) , .A1( u2_u7_u4_n134 ) , .A2( u2_u7_u4_n148 ) );
  AND3_X1 u2_u7_u4_U29 (.A1( u2_u7_u4_n119 ) , .A2( u2_u7_u4_n143 ) , .A3( u2_u7_u4_n154 ) , .ZN( u2_u7_u4_n161 ) );
  NOR2_X1 u2_u7_u4_U3 (.ZN( u2_u7_u4_n121 ) , .A1( u2_u7_u4_n181 ) , .A2( u2_u7_u4_n182 ) );
  AND2_X1 u2_u7_u4_U30 (.A1( u2_u7_u4_n145 ) , .A2( u2_u7_u4_n147 ) , .ZN( u2_u7_u4_n159 ) );
  INV_X1 u2_u7_u4_U31 (.A( u2_u7_u4_n158 ) , .ZN( u2_u7_u4_n182 ) );
  INV_X1 u2_u7_u4_U32 (.ZN( u2_u7_u4_n181 ) , .A( u2_u7_u4_n96 ) );
  INV_X1 u2_u7_u4_U33 (.A( u2_u7_u4_n144 ) , .ZN( u2_u7_u4_n179 ) );
  INV_X1 u2_u7_u4_U34 (.A( u2_u7_u4_n157 ) , .ZN( u2_u7_u4_n178 ) );
  NAND2_X1 u2_u7_u4_U35 (.A2( u2_u7_u4_n154 ) , .A1( u2_u7_u4_n96 ) , .ZN( u2_u7_u4_n97 ) );
  INV_X1 u2_u7_u4_U36 (.ZN( u2_u7_u4_n186 ) , .A( u2_u7_u4_n95 ) );
  OAI221_X1 u2_u7_u4_U37 (.C1( u2_u7_u4_n134 ) , .B1( u2_u7_u4_n158 ) , .B2( u2_u7_u4_n171 ) , .C2( u2_u7_u4_n173 ) , .A( u2_u7_u4_n94 ) , .ZN( u2_u7_u4_n95 ) );
  AOI222_X1 u2_u7_u4_U38 (.B2( u2_u7_u4_n132 ) , .A1( u2_u7_u4_n138 ) , .C2( u2_u7_u4_n175 ) , .A2( u2_u7_u4_n179 ) , .C1( u2_u7_u4_n181 ) , .B1( u2_u7_u4_n185 ) , .ZN( u2_u7_u4_n94 ) );
  INV_X1 u2_u7_u4_U39 (.A( u2_u7_u4_n113 ) , .ZN( u2_u7_u4_n185 ) );
  INV_X1 u2_u7_u4_U4 (.A( u2_u7_u4_n117 ) , .ZN( u2_u7_u4_n184 ) );
  INV_X1 u2_u7_u4_U40 (.A( u2_u7_u4_n143 ) , .ZN( u2_u7_u4_n183 ) );
  NOR2_X1 u2_u7_u4_U41 (.ZN( u2_u7_u4_n138 ) , .A1( u2_u7_u4_n168 ) , .A2( u2_u7_u4_n169 ) );
  NOR2_X1 u2_u7_u4_U42 (.A1( u2_u7_u4_n150 ) , .A2( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n153 ) );
  NOR2_X1 u2_u7_u4_U43 (.A2( u2_u7_u4_n128 ) , .A1( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n156 ) );
  AOI22_X1 u2_u7_u4_U44 (.B2( u2_u7_u4_n122 ) , .A1( u2_u7_u4_n123 ) , .ZN( u2_u7_u4_n124 ) , .B1( u2_u7_u4_n128 ) , .A2( u2_u7_u4_n172 ) );
  NAND2_X1 u2_u7_u4_U45 (.A2( u2_u7_u4_n120 ) , .ZN( u2_u7_u4_n123 ) , .A1( u2_u7_u4_n161 ) );
  INV_X1 u2_u7_u4_U46 (.A( u2_u7_u4_n153 ) , .ZN( u2_u7_u4_n172 ) );
  AOI22_X1 u2_u7_u4_U47 (.B2( u2_u7_u4_n132 ) , .A2( u2_u7_u4_n133 ) , .ZN( u2_u7_u4_n140 ) , .A1( u2_u7_u4_n150 ) , .B1( u2_u7_u4_n179 ) );
  NAND2_X1 u2_u7_u4_U48 (.ZN( u2_u7_u4_n133 ) , .A2( u2_u7_u4_n146 ) , .A1( u2_u7_u4_n154 ) );
  NAND2_X1 u2_u7_u4_U49 (.A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n154 ) , .A2( u2_u7_u4_n98 ) );
  NOR4_X1 u2_u7_u4_U5 (.A4( u2_u7_u4_n106 ) , .A3( u2_u7_u4_n107 ) , .A2( u2_u7_u4_n108 ) , .A1( u2_u7_u4_n109 ) , .ZN( u2_u7_u4_n110 ) );
  NAND2_X1 u2_u7_u4_U50 (.A1( u2_u7_u4_n101 ) , .ZN( u2_u7_u4_n158 ) , .A2( u2_u7_u4_n99 ) );
  AOI21_X1 u2_u7_u4_U51 (.ZN( u2_u7_u4_n127 ) , .A( u2_u7_u4_n136 ) , .B2( u2_u7_u4_n150 ) , .B1( u2_u7_u4_n180 ) );
  INV_X1 u2_u7_u4_U52 (.A( u2_u7_u4_n160 ) , .ZN( u2_u7_u4_n180 ) );
  NAND2_X1 u2_u7_u4_U53 (.A2( u2_u7_u4_n104 ) , .A1( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n146 ) );
  NAND2_X1 u2_u7_u4_U54 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n160 ) );
  NAND2_X1 u2_u7_u4_U55 (.ZN( u2_u7_u4_n134 ) , .A1( u2_u7_u4_n98 ) , .A2( u2_u7_u4_n99 ) );
  NAND2_X1 u2_u7_u4_U56 (.A1( u2_u7_u4_n103 ) , .A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n143 ) );
  NAND2_X1 u2_u7_u4_U57 (.A2( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n145 ) , .A1( u2_u7_u4_n98 ) );
  NAND2_X1 u2_u7_u4_U58 (.A1( u2_u7_u4_n100 ) , .A2( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n120 ) );
  NAND2_X1 u2_u7_u4_U59 (.A1( u2_u7_u4_n102 ) , .A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n148 ) );
  AOI21_X1 u2_u7_u4_U6 (.ZN( u2_u7_u4_n106 ) , .B2( u2_u7_u4_n146 ) , .B1( u2_u7_u4_n158 ) , .A( u2_u7_u4_n170 ) );
  NAND2_X1 u2_u7_u4_U60 (.A2( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n157 ) );
  INV_X1 u2_u7_u4_U61 (.A( u2_u7_u4_n150 ) , .ZN( u2_u7_u4_n173 ) );
  INV_X1 u2_u7_u4_U62 (.A( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n171 ) );
  NAND2_X1 u2_u7_u4_U63 (.A1( u2_u7_u4_n100 ) , .ZN( u2_u7_u4_n118 ) , .A2( u2_u7_u4_n99 ) );
  NAND2_X1 u2_u7_u4_U64 (.A2( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n144 ) );
  NAND2_X1 u2_u7_u4_U65 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n105 ) , .ZN( u2_u7_u4_n96 ) );
  INV_X1 u2_u7_u4_U66 (.A( u2_u7_u4_n128 ) , .ZN( u2_u7_u4_n174 ) );
  NAND2_X1 u2_u7_u4_U67 (.A2( u2_u7_u4_n102 ) , .ZN( u2_u7_u4_n119 ) , .A1( u2_u7_u4_n98 ) );
  NAND2_X1 u2_u7_u4_U68 (.A2( u2_u7_u4_n101 ) , .A1( u2_u7_u4_n103 ) , .ZN( u2_u7_u4_n147 ) );
  NAND2_X1 u2_u7_u4_U69 (.A2( u2_u7_u4_n104 ) , .ZN( u2_u7_u4_n113 ) , .A1( u2_u7_u4_n99 ) );
  AOI21_X1 u2_u7_u4_U7 (.ZN( u2_u7_u4_n108 ) , .B2( u2_u7_u4_n134 ) , .B1( u2_u7_u4_n155 ) , .A( u2_u7_u4_n156 ) );
  NOR2_X1 u2_u7_u4_U70 (.A2( u2_u7_X_28 ) , .ZN( u2_u7_u4_n150 ) , .A1( u2_u7_u4_n168 ) );
  NOR2_X1 u2_u7_u4_U71 (.A2( u2_u7_X_29 ) , .ZN( u2_u7_u4_n152 ) , .A1( u2_u7_u4_n169 ) );
  NOR2_X1 u2_u7_u4_U72 (.A2( u2_u7_X_26 ) , .ZN( u2_u7_u4_n100 ) , .A1( u2_u7_u4_n177 ) );
  NOR2_X1 u2_u7_u4_U73 (.A2( u2_u7_X_30 ) , .ZN( u2_u7_u4_n105 ) , .A1( u2_u7_u4_n176 ) );
  NOR2_X1 u2_u7_u4_U74 (.A2( u2_u7_X_28 ) , .A1( u2_u7_X_29 ) , .ZN( u2_u7_u4_n128 ) );
  NOR2_X1 u2_u7_u4_U75 (.A2( u2_u7_X_25 ) , .A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n98 ) );
  NOR2_X1 u2_u7_u4_U76 (.A2( u2_u7_X_27 ) , .A1( u2_u7_X_30 ) , .ZN( u2_u7_u4_n102 ) );
  AND2_X1 u2_u7_u4_U77 (.A2( u2_u7_X_25 ) , .A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n104 ) );
  AND2_X1 u2_u7_u4_U78 (.A1( u2_u7_X_30 ) , .A2( u2_u7_u4_n176 ) , .ZN( u2_u7_u4_n99 ) );
  AND2_X1 u2_u7_u4_U79 (.A1( u2_u7_X_26 ) , .ZN( u2_u7_u4_n101 ) , .A2( u2_u7_u4_n177 ) );
  AOI21_X1 u2_u7_u4_U8 (.ZN( u2_u7_u4_n109 ) , .A( u2_u7_u4_n153 ) , .B1( u2_u7_u4_n159 ) , .B2( u2_u7_u4_n184 ) );
  AND2_X1 u2_u7_u4_U80 (.A1( u2_u7_X_27 ) , .A2( u2_u7_X_30 ) , .ZN( u2_u7_u4_n103 ) );
  INV_X1 u2_u7_u4_U81 (.A( u2_u7_X_28 ) , .ZN( u2_u7_u4_n169 ) );
  INV_X1 u2_u7_u4_U82 (.A( u2_u7_X_29 ) , .ZN( u2_u7_u4_n168 ) );
  INV_X1 u2_u7_u4_U83 (.A( u2_u7_X_25 ) , .ZN( u2_u7_u4_n177 ) );
  INV_X1 u2_u7_u4_U84 (.A( u2_u7_X_27 ) , .ZN( u2_u7_u4_n176 ) );
  NAND4_X1 u2_u7_u4_U85 (.ZN( u2_out7_25 ) , .A4( u2_u7_u4_n139 ) , .A3( u2_u7_u4_n140 ) , .A2( u2_u7_u4_n141 ) , .A1( u2_u7_u4_n142 ) );
  OAI21_X1 u2_u7_u4_U86 (.A( u2_u7_u4_n128 ) , .B2( u2_u7_u4_n129 ) , .B1( u2_u7_u4_n130 ) , .ZN( u2_u7_u4_n142 ) );
  OAI21_X1 u2_u7_u4_U87 (.B2( u2_u7_u4_n131 ) , .ZN( u2_u7_u4_n141 ) , .A( u2_u7_u4_n175 ) , .B1( u2_u7_u4_n183 ) );
  NAND4_X1 u2_u7_u4_U88 (.ZN( u2_out7_14 ) , .A4( u2_u7_u4_n124 ) , .A3( u2_u7_u4_n125 ) , .A2( u2_u7_u4_n126 ) , .A1( u2_u7_u4_n127 ) );
  AOI22_X1 u2_u7_u4_U89 (.B2( u2_u7_u4_n117 ) , .ZN( u2_u7_u4_n126 ) , .A1( u2_u7_u4_n129 ) , .B1( u2_u7_u4_n152 ) , .A2( u2_u7_u4_n175 ) );
  AOI211_X1 u2_u7_u4_U9 (.B( u2_u7_u4_n136 ) , .A( u2_u7_u4_n137 ) , .C2( u2_u7_u4_n138 ) , .ZN( u2_u7_u4_n139 ) , .C1( u2_u7_u4_n182 ) );
  AOI22_X1 u2_u7_u4_U90 (.ZN( u2_u7_u4_n125 ) , .B2( u2_u7_u4_n131 ) , .A2( u2_u7_u4_n132 ) , .B1( u2_u7_u4_n138 ) , .A1( u2_u7_u4_n178 ) );
  NAND4_X1 u2_u7_u4_U91 (.ZN( u2_out7_8 ) , .A4( u2_u7_u4_n110 ) , .A3( u2_u7_u4_n111 ) , .A2( u2_u7_u4_n112 ) , .A1( u2_u7_u4_n186 ) );
  NAND2_X1 u2_u7_u4_U92 (.ZN( u2_u7_u4_n112 ) , .A2( u2_u7_u4_n130 ) , .A1( u2_u7_u4_n150 ) );
  AOI22_X1 u2_u7_u4_U93 (.ZN( u2_u7_u4_n111 ) , .B2( u2_u7_u4_n132 ) , .A1( u2_u7_u4_n152 ) , .B1( u2_u7_u4_n178 ) , .A2( u2_u7_u4_n97 ) );
  AOI22_X1 u2_u7_u4_U94 (.B2( u2_u7_u4_n149 ) , .B1( u2_u7_u4_n150 ) , .A2( u2_u7_u4_n151 ) , .A1( u2_u7_u4_n152 ) , .ZN( u2_u7_u4_n167 ) );
  NOR4_X1 u2_u7_u4_U95 (.A4( u2_u7_u4_n162 ) , .A3( u2_u7_u4_n163 ) , .A2( u2_u7_u4_n164 ) , .A1( u2_u7_u4_n165 ) , .ZN( u2_u7_u4_n166 ) );
  NAND3_X1 u2_u7_u4_U96 (.ZN( u2_out7_3 ) , .A3( u2_u7_u4_n166 ) , .A1( u2_u7_u4_n167 ) , .A2( u2_u7_u4_n186 ) );
  NAND3_X1 u2_u7_u4_U97 (.A3( u2_u7_u4_n146 ) , .A2( u2_u7_u4_n147 ) , .A1( u2_u7_u4_n148 ) , .ZN( u2_u7_u4_n149 ) );
  NAND3_X1 u2_u7_u4_U98 (.A3( u2_u7_u4_n143 ) , .A2( u2_u7_u4_n144 ) , .A1( u2_u7_u4_n145 ) , .ZN( u2_u7_u4_n151 ) );
  NAND3_X1 u2_u7_u4_U99 (.A3( u2_u7_u4_n121 ) , .ZN( u2_u7_u4_n122 ) , .A2( u2_u7_u4_n144 ) , .A1( u2_u7_u4_n154 ) );
  INV_X1 u2_u7_u5_U10 (.A( u2_u7_u5_n121 ) , .ZN( u2_u7_u5_n177 ) );
  NOR3_X1 u2_u7_u5_U100 (.A3( u2_u7_u5_n141 ) , .A1( u2_u7_u5_n142 ) , .ZN( u2_u7_u5_n143 ) , .A2( u2_u7_u5_n191 ) );
  NAND4_X1 u2_u7_u5_U101 (.ZN( u2_out7_4 ) , .A4( u2_u7_u5_n112 ) , .A2( u2_u7_u5_n113 ) , .A1( u2_u7_u5_n114 ) , .A3( u2_u7_u5_n195 ) );
  AOI211_X1 u2_u7_u5_U102 (.A( u2_u7_u5_n110 ) , .C1( u2_u7_u5_n111 ) , .ZN( u2_u7_u5_n112 ) , .B( u2_u7_u5_n118 ) , .C2( u2_u7_u5_n177 ) );
  AOI222_X1 u2_u7_u5_U103 (.ZN( u2_u7_u5_n113 ) , .A1( u2_u7_u5_n131 ) , .C1( u2_u7_u5_n148 ) , .B2( u2_u7_u5_n174 ) , .C2( u2_u7_u5_n178 ) , .A2( u2_u7_u5_n179 ) , .B1( u2_u7_u5_n99 ) );
  NAND3_X1 u2_u7_u5_U104 (.A2( u2_u7_u5_n154 ) , .A3( u2_u7_u5_n158 ) , .A1( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n99 ) );
  NOR2_X1 u2_u7_u5_U11 (.ZN( u2_u7_u5_n160 ) , .A2( u2_u7_u5_n173 ) , .A1( u2_u7_u5_n177 ) );
  INV_X1 u2_u7_u5_U12 (.A( u2_u7_u5_n150 ) , .ZN( u2_u7_u5_n174 ) );
  AOI21_X1 u2_u7_u5_U13 (.A( u2_u7_u5_n160 ) , .B2( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n162 ) , .B1( u2_u7_u5_n192 ) );
  INV_X1 u2_u7_u5_U14 (.A( u2_u7_u5_n159 ) , .ZN( u2_u7_u5_n192 ) );
  AOI21_X1 u2_u7_u5_U15 (.A( u2_u7_u5_n156 ) , .B2( u2_u7_u5_n157 ) , .B1( u2_u7_u5_n158 ) , .ZN( u2_u7_u5_n163 ) );
  AOI21_X1 u2_u7_u5_U16 (.B2( u2_u7_u5_n139 ) , .B1( u2_u7_u5_n140 ) , .ZN( u2_u7_u5_n141 ) , .A( u2_u7_u5_n150 ) );
  OAI21_X1 u2_u7_u5_U17 (.A( u2_u7_u5_n133 ) , .B2( u2_u7_u5_n134 ) , .B1( u2_u7_u5_n135 ) , .ZN( u2_u7_u5_n142 ) );
  OAI21_X1 u2_u7_u5_U18 (.ZN( u2_u7_u5_n133 ) , .B2( u2_u7_u5_n147 ) , .A( u2_u7_u5_n173 ) , .B1( u2_u7_u5_n188 ) );
  NAND2_X1 u2_u7_u5_U19 (.A2( u2_u7_u5_n119 ) , .A1( u2_u7_u5_n123 ) , .ZN( u2_u7_u5_n137 ) );
  INV_X1 u2_u7_u5_U20 (.A( u2_u7_u5_n155 ) , .ZN( u2_u7_u5_n194 ) );
  NAND2_X1 u2_u7_u5_U21 (.A1( u2_u7_u5_n121 ) , .ZN( u2_u7_u5_n132 ) , .A2( u2_u7_u5_n172 ) );
  NAND2_X1 u2_u7_u5_U22 (.A2( u2_u7_u5_n122 ) , .ZN( u2_u7_u5_n136 ) , .A1( u2_u7_u5_n154 ) );
  NAND2_X1 u2_u7_u5_U23 (.A2( u2_u7_u5_n119 ) , .A1( u2_u7_u5_n120 ) , .ZN( u2_u7_u5_n159 ) );
  INV_X1 u2_u7_u5_U24 (.A( u2_u7_u5_n156 ) , .ZN( u2_u7_u5_n175 ) );
  INV_X1 u2_u7_u5_U25 (.A( u2_u7_u5_n158 ) , .ZN( u2_u7_u5_n188 ) );
  INV_X1 u2_u7_u5_U26 (.A( u2_u7_u5_n152 ) , .ZN( u2_u7_u5_n179 ) );
  INV_X1 u2_u7_u5_U27 (.A( u2_u7_u5_n140 ) , .ZN( u2_u7_u5_n182 ) );
  INV_X1 u2_u7_u5_U28 (.A( u2_u7_u5_n151 ) , .ZN( u2_u7_u5_n183 ) );
  INV_X1 u2_u7_u5_U29 (.A( u2_u7_u5_n123 ) , .ZN( u2_u7_u5_n185 ) );
  NOR2_X1 u2_u7_u5_U3 (.ZN( u2_u7_u5_n134 ) , .A1( u2_u7_u5_n183 ) , .A2( u2_u7_u5_n190 ) );
  INV_X1 u2_u7_u5_U30 (.A( u2_u7_u5_n161 ) , .ZN( u2_u7_u5_n184 ) );
  INV_X1 u2_u7_u5_U31 (.A( u2_u7_u5_n139 ) , .ZN( u2_u7_u5_n189 ) );
  INV_X1 u2_u7_u5_U32 (.A( u2_u7_u5_n157 ) , .ZN( u2_u7_u5_n190 ) );
  INV_X1 u2_u7_u5_U33 (.A( u2_u7_u5_n120 ) , .ZN( u2_u7_u5_n193 ) );
  NAND2_X1 u2_u7_u5_U34 (.ZN( u2_u7_u5_n111 ) , .A1( u2_u7_u5_n140 ) , .A2( u2_u7_u5_n155 ) );
  NOR2_X1 u2_u7_u5_U35 (.ZN( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n170 ) , .A2( u2_u7_u5_n180 ) );
  INV_X1 u2_u7_u5_U36 (.A( u2_u7_u5_n117 ) , .ZN( u2_u7_u5_n196 ) );
  OAI221_X1 u2_u7_u5_U37 (.A( u2_u7_u5_n116 ) , .ZN( u2_u7_u5_n117 ) , .B2( u2_u7_u5_n119 ) , .C1( u2_u7_u5_n153 ) , .C2( u2_u7_u5_n158 ) , .B1( u2_u7_u5_n172 ) );
  AOI222_X1 u2_u7_u5_U38 (.ZN( u2_u7_u5_n116 ) , .B2( u2_u7_u5_n145 ) , .C1( u2_u7_u5_n148 ) , .A2( u2_u7_u5_n174 ) , .C2( u2_u7_u5_n177 ) , .B1( u2_u7_u5_n187 ) , .A1( u2_u7_u5_n193 ) );
  INV_X1 u2_u7_u5_U39 (.A( u2_u7_u5_n115 ) , .ZN( u2_u7_u5_n187 ) );
  INV_X1 u2_u7_u5_U4 (.A( u2_u7_u5_n138 ) , .ZN( u2_u7_u5_n191 ) );
  AOI22_X1 u2_u7_u5_U40 (.B2( u2_u7_u5_n131 ) , .A2( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n169 ) , .B1( u2_u7_u5_n174 ) , .A1( u2_u7_u5_n185 ) );
  NOR2_X1 u2_u7_u5_U41 (.A1( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n150 ) , .A2( u2_u7_u5_n173 ) );
  AOI21_X1 u2_u7_u5_U42 (.A( u2_u7_u5_n118 ) , .B2( u2_u7_u5_n145 ) , .ZN( u2_u7_u5_n168 ) , .B1( u2_u7_u5_n186 ) );
  INV_X1 u2_u7_u5_U43 (.A( u2_u7_u5_n122 ) , .ZN( u2_u7_u5_n186 ) );
  NOR2_X1 u2_u7_u5_U44 (.A1( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n152 ) , .A2( u2_u7_u5_n176 ) );
  NOR2_X1 u2_u7_u5_U45 (.A1( u2_u7_u5_n115 ) , .ZN( u2_u7_u5_n118 ) , .A2( u2_u7_u5_n153 ) );
  NOR2_X1 u2_u7_u5_U46 (.A2( u2_u7_u5_n145 ) , .ZN( u2_u7_u5_n156 ) , .A1( u2_u7_u5_n174 ) );
  NOR2_X1 u2_u7_u5_U47 (.ZN( u2_u7_u5_n121 ) , .A2( u2_u7_u5_n145 ) , .A1( u2_u7_u5_n176 ) );
  AOI22_X1 u2_u7_u5_U48 (.ZN( u2_u7_u5_n114 ) , .A2( u2_u7_u5_n137 ) , .A1( u2_u7_u5_n145 ) , .B2( u2_u7_u5_n175 ) , .B1( u2_u7_u5_n193 ) );
  OAI211_X1 u2_u7_u5_U49 (.B( u2_u7_u5_n124 ) , .A( u2_u7_u5_n125 ) , .C2( u2_u7_u5_n126 ) , .C1( u2_u7_u5_n127 ) , .ZN( u2_u7_u5_n128 ) );
  OAI21_X1 u2_u7_u5_U5 (.B2( u2_u7_u5_n136 ) , .B1( u2_u7_u5_n137 ) , .ZN( u2_u7_u5_n138 ) , .A( u2_u7_u5_n177 ) );
  NOR3_X1 u2_u7_u5_U50 (.ZN( u2_u7_u5_n127 ) , .A1( u2_u7_u5_n136 ) , .A3( u2_u7_u5_n148 ) , .A2( u2_u7_u5_n182 ) );
  OAI21_X1 u2_u7_u5_U51 (.ZN( u2_u7_u5_n124 ) , .A( u2_u7_u5_n177 ) , .B2( u2_u7_u5_n183 ) , .B1( u2_u7_u5_n189 ) );
  OAI21_X1 u2_u7_u5_U52 (.ZN( u2_u7_u5_n125 ) , .A( u2_u7_u5_n174 ) , .B2( u2_u7_u5_n185 ) , .B1( u2_u7_u5_n190 ) );
  AOI21_X1 u2_u7_u5_U53 (.A( u2_u7_u5_n153 ) , .B2( u2_u7_u5_n154 ) , .B1( u2_u7_u5_n155 ) , .ZN( u2_u7_u5_n164 ) );
  AOI21_X1 u2_u7_u5_U54 (.ZN( u2_u7_u5_n110 ) , .B1( u2_u7_u5_n122 ) , .B2( u2_u7_u5_n139 ) , .A( u2_u7_u5_n153 ) );
  INV_X1 u2_u7_u5_U55 (.A( u2_u7_u5_n153 ) , .ZN( u2_u7_u5_n176 ) );
  INV_X1 u2_u7_u5_U56 (.A( u2_u7_u5_n126 ) , .ZN( u2_u7_u5_n173 ) );
  AND2_X1 u2_u7_u5_U57 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n147 ) );
  AND2_X1 u2_u7_u5_U58 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n148 ) );
  NAND2_X1 u2_u7_u5_U59 (.A1( u2_u7_u5_n105 ) , .A2( u2_u7_u5_n106 ) , .ZN( u2_u7_u5_n158 ) );
  INV_X1 u2_u7_u5_U6 (.A( u2_u7_u5_n135 ) , .ZN( u2_u7_u5_n178 ) );
  NAND2_X1 u2_u7_u5_U60 (.A2( u2_u7_u5_n108 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n139 ) );
  NAND2_X1 u2_u7_u5_U61 (.A1( u2_u7_u5_n106 ) , .A2( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n119 ) );
  NAND2_X1 u2_u7_u5_U62 (.A2( u2_u7_u5_n103 ) , .A1( u2_u7_u5_n105 ) , .ZN( u2_u7_u5_n140 ) );
  NAND2_X1 u2_u7_u5_U63 (.A2( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n105 ) , .ZN( u2_u7_u5_n155 ) );
  NAND2_X1 u2_u7_u5_U64 (.A2( u2_u7_u5_n106 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n122 ) );
  NAND2_X1 u2_u7_u5_U65 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n106 ) , .ZN( u2_u7_u5_n115 ) );
  NAND2_X1 u2_u7_u5_U66 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n103 ) , .ZN( u2_u7_u5_n161 ) );
  NAND2_X1 u2_u7_u5_U67 (.A1( u2_u7_u5_n105 ) , .A2( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n154 ) );
  INV_X1 u2_u7_u5_U68 (.A( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n172 ) );
  NAND2_X1 u2_u7_u5_U69 (.A1( u2_u7_u5_n103 ) , .A2( u2_u7_u5_n108 ) , .ZN( u2_u7_u5_n123 ) );
  OAI22_X1 u2_u7_u5_U7 (.B2( u2_u7_u5_n149 ) , .B1( u2_u7_u5_n150 ) , .A2( u2_u7_u5_n151 ) , .A1( u2_u7_u5_n152 ) , .ZN( u2_u7_u5_n165 ) );
  NAND2_X1 u2_u7_u5_U70 (.A2( u2_u7_u5_n103 ) , .A1( u2_u7_u5_n107 ) , .ZN( u2_u7_u5_n151 ) );
  NAND2_X1 u2_u7_u5_U71 (.A2( u2_u7_u5_n107 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n120 ) );
  NAND2_X1 u2_u7_u5_U72 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n109 ) , .ZN( u2_u7_u5_n157 ) );
  AND2_X1 u2_u7_u5_U73 (.A2( u2_u7_u5_n100 ) , .A1( u2_u7_u5_n104 ) , .ZN( u2_u7_u5_n131 ) );
  INV_X1 u2_u7_u5_U74 (.A( u2_u7_u5_n102 ) , .ZN( u2_u7_u5_n195 ) );
  OAI221_X1 u2_u7_u5_U75 (.A( u2_u7_u5_n101 ) , .ZN( u2_u7_u5_n102 ) , .C2( u2_u7_u5_n115 ) , .C1( u2_u7_u5_n126 ) , .B1( u2_u7_u5_n134 ) , .B2( u2_u7_u5_n160 ) );
  OAI21_X1 u2_u7_u5_U76 (.ZN( u2_u7_u5_n101 ) , .B1( u2_u7_u5_n137 ) , .A( u2_u7_u5_n146 ) , .B2( u2_u7_u5_n147 ) );
  NOR2_X1 u2_u7_u5_U77 (.A2( u2_u7_X_34 ) , .A1( u2_u7_X_35 ) , .ZN( u2_u7_u5_n145 ) );
  NOR2_X1 u2_u7_u5_U78 (.A2( u2_u7_X_34 ) , .ZN( u2_u7_u5_n146 ) , .A1( u2_u7_u5_n171 ) );
  NOR2_X1 u2_u7_u5_U79 (.A2( u2_u7_X_31 ) , .A1( u2_u7_X_32 ) , .ZN( u2_u7_u5_n103 ) );
  NOR3_X1 u2_u7_u5_U8 (.A2( u2_u7_u5_n147 ) , .A1( u2_u7_u5_n148 ) , .ZN( u2_u7_u5_n149 ) , .A3( u2_u7_u5_n194 ) );
  NOR2_X1 u2_u7_u5_U80 (.A2( u2_u7_X_36 ) , .ZN( u2_u7_u5_n105 ) , .A1( u2_u7_u5_n180 ) );
  NOR2_X1 u2_u7_u5_U81 (.A2( u2_u7_X_33 ) , .ZN( u2_u7_u5_n108 ) , .A1( u2_u7_u5_n170 ) );
  NOR2_X1 u2_u7_u5_U82 (.A2( u2_u7_X_33 ) , .A1( u2_u7_X_36 ) , .ZN( u2_u7_u5_n107 ) );
  NOR2_X1 u2_u7_u5_U83 (.A2( u2_u7_X_31 ) , .ZN( u2_u7_u5_n104 ) , .A1( u2_u7_u5_n181 ) );
  NAND2_X1 u2_u7_u5_U84 (.A2( u2_u7_X_34 ) , .A1( u2_u7_X_35 ) , .ZN( u2_u7_u5_n153 ) );
  NAND2_X1 u2_u7_u5_U85 (.A1( u2_u7_X_34 ) , .ZN( u2_u7_u5_n126 ) , .A2( u2_u7_u5_n171 ) );
  AND2_X1 u2_u7_u5_U86 (.A1( u2_u7_X_31 ) , .A2( u2_u7_X_32 ) , .ZN( u2_u7_u5_n106 ) );
  AND2_X1 u2_u7_u5_U87 (.A1( u2_u7_X_31 ) , .ZN( u2_u7_u5_n109 ) , .A2( u2_u7_u5_n181 ) );
  INV_X1 u2_u7_u5_U88 (.A( u2_u7_X_33 ) , .ZN( u2_u7_u5_n180 ) );
  INV_X1 u2_u7_u5_U89 (.A( u2_u7_X_35 ) , .ZN( u2_u7_u5_n171 ) );
  NOR2_X1 u2_u7_u5_U9 (.ZN( u2_u7_u5_n135 ) , .A1( u2_u7_u5_n173 ) , .A2( u2_u7_u5_n176 ) );
  INV_X1 u2_u7_u5_U90 (.A( u2_u7_X_36 ) , .ZN( u2_u7_u5_n170 ) );
  INV_X1 u2_u7_u5_U91 (.A( u2_u7_X_32 ) , .ZN( u2_u7_u5_n181 ) );
  NAND4_X1 u2_u7_u5_U92 (.ZN( u2_out7_29 ) , .A4( u2_u7_u5_n129 ) , .A3( u2_u7_u5_n130 ) , .A2( u2_u7_u5_n168 ) , .A1( u2_u7_u5_n196 ) );
  AOI221_X1 u2_u7_u5_U93 (.A( u2_u7_u5_n128 ) , .ZN( u2_u7_u5_n129 ) , .C2( u2_u7_u5_n132 ) , .B2( u2_u7_u5_n159 ) , .B1( u2_u7_u5_n176 ) , .C1( u2_u7_u5_n184 ) );
  AOI222_X1 u2_u7_u5_U94 (.ZN( u2_u7_u5_n130 ) , .A2( u2_u7_u5_n146 ) , .B1( u2_u7_u5_n147 ) , .C2( u2_u7_u5_n175 ) , .B2( u2_u7_u5_n179 ) , .A1( u2_u7_u5_n188 ) , .C1( u2_u7_u5_n194 ) );
  NAND4_X1 u2_u7_u5_U95 (.ZN( u2_out7_19 ) , .A4( u2_u7_u5_n166 ) , .A3( u2_u7_u5_n167 ) , .A2( u2_u7_u5_n168 ) , .A1( u2_u7_u5_n169 ) );
  AOI22_X1 u2_u7_u5_U96 (.B2( u2_u7_u5_n145 ) , .A2( u2_u7_u5_n146 ) , .ZN( u2_u7_u5_n167 ) , .B1( u2_u7_u5_n182 ) , .A1( u2_u7_u5_n189 ) );
  NOR4_X1 u2_u7_u5_U97 (.A4( u2_u7_u5_n162 ) , .A3( u2_u7_u5_n163 ) , .A2( u2_u7_u5_n164 ) , .A1( u2_u7_u5_n165 ) , .ZN( u2_u7_u5_n166 ) );
  NAND4_X1 u2_u7_u5_U98 (.ZN( u2_out7_11 ) , .A4( u2_u7_u5_n143 ) , .A3( u2_u7_u5_n144 ) , .A2( u2_u7_u5_n169 ) , .A1( u2_u7_u5_n196 ) );
  AOI22_X1 u2_u7_u5_U99 (.A2( u2_u7_u5_n132 ) , .ZN( u2_u7_u5_n144 ) , .B2( u2_u7_u5_n145 ) , .B1( u2_u7_u5_n184 ) , .A1( u2_u7_u5_n194 ) );
  INV_X1 u2_u7_u6_U10 (.ZN( u2_u7_u6_n172 ) , .A( u2_u7_u6_n88 ) );
  OAI21_X1 u2_u7_u6_U11 (.A( u2_u7_u6_n159 ) , .B1( u2_u7_u6_n169 ) , .B2( u2_u7_u6_n173 ) , .ZN( u2_u7_u6_n90 ) );
  AOI22_X1 u2_u7_u6_U12 (.A2( u2_u7_u6_n151 ) , .B2( u2_u7_u6_n161 ) , .A1( u2_u7_u6_n167 ) , .B1( u2_u7_u6_n170 ) , .ZN( u2_u7_u6_n89 ) );
  AOI21_X1 u2_u7_u6_U13 (.ZN( u2_u7_u6_n106 ) , .A( u2_u7_u6_n142 ) , .B2( u2_u7_u6_n159 ) , .B1( u2_u7_u6_n164 ) );
  INV_X1 u2_u7_u6_U14 (.A( u2_u7_u6_n155 ) , .ZN( u2_u7_u6_n161 ) );
  INV_X1 u2_u7_u6_U15 (.A( u2_u7_u6_n128 ) , .ZN( u2_u7_u6_n164 ) );
  NAND2_X1 u2_u7_u6_U16 (.ZN( u2_u7_u6_n110 ) , .A1( u2_u7_u6_n122 ) , .A2( u2_u7_u6_n129 ) );
  NAND2_X1 u2_u7_u6_U17 (.ZN( u2_u7_u6_n124 ) , .A2( u2_u7_u6_n146 ) , .A1( u2_u7_u6_n148 ) );
  INV_X1 u2_u7_u6_U18 (.A( u2_u7_u6_n132 ) , .ZN( u2_u7_u6_n171 ) );
  AND2_X1 u2_u7_u6_U19 (.A1( u2_u7_u6_n100 ) , .ZN( u2_u7_u6_n130 ) , .A2( u2_u7_u6_n147 ) );
  INV_X1 u2_u7_u6_U20 (.A( u2_u7_u6_n127 ) , .ZN( u2_u7_u6_n173 ) );
  INV_X1 u2_u7_u6_U21 (.A( u2_u7_u6_n121 ) , .ZN( u2_u7_u6_n167 ) );
  INV_X1 u2_u7_u6_U22 (.A( u2_u7_u6_n100 ) , .ZN( u2_u7_u6_n169 ) );
  INV_X1 u2_u7_u6_U23 (.A( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n170 ) );
  INV_X1 u2_u7_u6_U24 (.A( u2_u7_u6_n113 ) , .ZN( u2_u7_u6_n168 ) );
  AND2_X1 u2_u7_u6_U25 (.A1( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n119 ) , .ZN( u2_u7_u6_n133 ) );
  AND2_X1 u2_u7_u6_U26 (.A2( u2_u7_u6_n121 ) , .A1( u2_u7_u6_n122 ) , .ZN( u2_u7_u6_n131 ) );
  AND3_X1 u2_u7_u6_U27 (.ZN( u2_u7_u6_n120 ) , .A2( u2_u7_u6_n127 ) , .A1( u2_u7_u6_n132 ) , .A3( u2_u7_u6_n145 ) );
  INV_X1 u2_u7_u6_U28 (.A( u2_u7_u6_n146 ) , .ZN( u2_u7_u6_n163 ) );
  AOI222_X1 u2_u7_u6_U29 (.ZN( u2_u7_u6_n114 ) , .A1( u2_u7_u6_n118 ) , .A2( u2_u7_u6_n126 ) , .B2( u2_u7_u6_n151 ) , .C2( u2_u7_u6_n159 ) , .C1( u2_u7_u6_n168 ) , .B1( u2_u7_u6_n169 ) );
  INV_X1 u2_u7_u6_U3 (.A( u2_u7_u6_n110 ) , .ZN( u2_u7_u6_n166 ) );
  NOR2_X1 u2_u7_u6_U30 (.A1( u2_u7_u6_n162 ) , .A2( u2_u7_u6_n165 ) , .ZN( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U31 (.A1( u2_u7_u6_n144 ) , .ZN( u2_u7_u6_n151 ) , .A2( u2_u7_u6_n158 ) );
  NAND2_X1 u2_u7_u6_U32 (.ZN( u2_u7_u6_n132 ) , .A1( u2_u7_u6_n91 ) , .A2( u2_u7_u6_n97 ) );
  AOI22_X1 u2_u7_u6_U33 (.B2( u2_u7_u6_n110 ) , .B1( u2_u7_u6_n111 ) , .A1( u2_u7_u6_n112 ) , .ZN( u2_u7_u6_n115 ) , .A2( u2_u7_u6_n161 ) );
  NAND4_X1 u2_u7_u6_U34 (.A3( u2_u7_u6_n109 ) , .ZN( u2_u7_u6_n112 ) , .A4( u2_u7_u6_n132 ) , .A2( u2_u7_u6_n147 ) , .A1( u2_u7_u6_n166 ) );
  NOR2_X1 u2_u7_u6_U35 (.ZN( u2_u7_u6_n109 ) , .A1( u2_u7_u6_n170 ) , .A2( u2_u7_u6_n173 ) );
  NOR2_X1 u2_u7_u6_U36 (.A2( u2_u7_u6_n126 ) , .ZN( u2_u7_u6_n155 ) , .A1( u2_u7_u6_n160 ) );
  NAND2_X1 u2_u7_u6_U37 (.ZN( u2_u7_u6_n146 ) , .A2( u2_u7_u6_n94 ) , .A1( u2_u7_u6_n99 ) );
  AOI21_X1 u2_u7_u6_U38 (.A( u2_u7_u6_n144 ) , .B2( u2_u7_u6_n145 ) , .B1( u2_u7_u6_n146 ) , .ZN( u2_u7_u6_n150 ) );
  AOI211_X1 u2_u7_u6_U39 (.B( u2_u7_u6_n134 ) , .A( u2_u7_u6_n135 ) , .C1( u2_u7_u6_n136 ) , .ZN( u2_u7_u6_n137 ) , .C2( u2_u7_u6_n151 ) );
  INV_X1 u2_u7_u6_U4 (.A( u2_u7_u6_n142 ) , .ZN( u2_u7_u6_n174 ) );
  NAND4_X1 u2_u7_u6_U40 (.A4( u2_u7_u6_n127 ) , .A3( u2_u7_u6_n128 ) , .A2( u2_u7_u6_n129 ) , .A1( u2_u7_u6_n130 ) , .ZN( u2_u7_u6_n136 ) );
  AOI21_X1 u2_u7_u6_U41 (.B2( u2_u7_u6_n132 ) , .B1( u2_u7_u6_n133 ) , .ZN( u2_u7_u6_n134 ) , .A( u2_u7_u6_n158 ) );
  AOI21_X1 u2_u7_u6_U42 (.B1( u2_u7_u6_n131 ) , .ZN( u2_u7_u6_n135 ) , .A( u2_u7_u6_n144 ) , .B2( u2_u7_u6_n146 ) );
  INV_X1 u2_u7_u6_U43 (.A( u2_u7_u6_n111 ) , .ZN( u2_u7_u6_n158 ) );
  NAND2_X1 u2_u7_u6_U44 (.ZN( u2_u7_u6_n127 ) , .A1( u2_u7_u6_n91 ) , .A2( u2_u7_u6_n92 ) );
  NAND2_X1 u2_u7_u6_U45 (.ZN( u2_u7_u6_n129 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n96 ) );
  INV_X1 u2_u7_u6_U46 (.A( u2_u7_u6_n144 ) , .ZN( u2_u7_u6_n159 ) );
  NAND2_X1 u2_u7_u6_U47 (.ZN( u2_u7_u6_n145 ) , .A2( u2_u7_u6_n97 ) , .A1( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U48 (.ZN( u2_u7_u6_n148 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n94 ) );
  NAND2_X1 u2_u7_u6_U49 (.ZN( u2_u7_u6_n108 ) , .A2( u2_u7_u6_n139 ) , .A1( u2_u7_u6_n144 ) );
  NAND2_X1 u2_u7_u6_U5 (.A2( u2_u7_u6_n143 ) , .ZN( u2_u7_u6_n152 ) , .A1( u2_u7_u6_n166 ) );
  NAND2_X1 u2_u7_u6_U50 (.ZN( u2_u7_u6_n121 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n97 ) );
  NAND2_X1 u2_u7_u6_U51 (.ZN( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n95 ) );
  AND2_X1 u2_u7_u6_U52 (.ZN( u2_u7_u6_n118 ) , .A2( u2_u7_u6_n91 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U53 (.ZN( u2_u7_u6_n147 ) , .A2( u2_u7_u6_n98 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U54 (.ZN( u2_u7_u6_n128 ) , .A1( u2_u7_u6_n94 ) , .A2( u2_u7_u6_n96 ) );
  NAND2_X1 u2_u7_u6_U55 (.ZN( u2_u7_u6_n119 ) , .A2( u2_u7_u6_n95 ) , .A1( u2_u7_u6_n99 ) );
  NAND2_X1 u2_u7_u6_U56 (.ZN( u2_u7_u6_n123 ) , .A2( u2_u7_u6_n91 ) , .A1( u2_u7_u6_n96 ) );
  NAND2_X1 u2_u7_u6_U57 (.ZN( u2_u7_u6_n100 ) , .A2( u2_u7_u6_n92 ) , .A1( u2_u7_u6_n98 ) );
  NAND2_X1 u2_u7_u6_U58 (.ZN( u2_u7_u6_n122 ) , .A1( u2_u7_u6_n94 ) , .A2( u2_u7_u6_n97 ) );
  INV_X1 u2_u7_u6_U59 (.A( u2_u7_u6_n139 ) , .ZN( u2_u7_u6_n160 ) );
  AOI22_X1 u2_u7_u6_U6 (.B2( u2_u7_u6_n101 ) , .A1( u2_u7_u6_n102 ) , .ZN( u2_u7_u6_n103 ) , .B1( u2_u7_u6_n160 ) , .A2( u2_u7_u6_n161 ) );
  NAND2_X1 u2_u7_u6_U60 (.ZN( u2_u7_u6_n113 ) , .A1( u2_u7_u6_n96 ) , .A2( u2_u7_u6_n98 ) );
  NOR2_X1 u2_u7_u6_U61 (.A2( u2_u7_X_40 ) , .A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n126 ) );
  NOR2_X1 u2_u7_u6_U62 (.A2( u2_u7_X_39 ) , .A1( u2_u7_X_42 ) , .ZN( u2_u7_u6_n92 ) );
  NOR2_X1 u2_u7_u6_U63 (.A2( u2_u7_X_39 ) , .A1( u2_u7_u6_n156 ) , .ZN( u2_u7_u6_n97 ) );
  NOR2_X1 u2_u7_u6_U64 (.A2( u2_u7_X_38 ) , .A1( u2_u7_u6_n165 ) , .ZN( u2_u7_u6_n95 ) );
  NOR2_X1 u2_u7_u6_U65 (.A2( u2_u7_X_41 ) , .ZN( u2_u7_u6_n111 ) , .A1( u2_u7_u6_n157 ) );
  NOR2_X1 u2_u7_u6_U66 (.A2( u2_u7_X_37 ) , .A1( u2_u7_u6_n162 ) , .ZN( u2_u7_u6_n94 ) );
  NOR2_X1 u2_u7_u6_U67 (.A2( u2_u7_X_37 ) , .A1( u2_u7_X_38 ) , .ZN( u2_u7_u6_n91 ) );
  NAND2_X1 u2_u7_u6_U68 (.A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n144 ) , .A2( u2_u7_u6_n157 ) );
  NAND2_X1 u2_u7_u6_U69 (.A2( u2_u7_X_40 ) , .A1( u2_u7_X_41 ) , .ZN( u2_u7_u6_n139 ) );
  NOR2_X1 u2_u7_u6_U7 (.A1( u2_u7_u6_n118 ) , .ZN( u2_u7_u6_n143 ) , .A2( u2_u7_u6_n168 ) );
  AND2_X1 u2_u7_u6_U70 (.A1( u2_u7_X_39 ) , .A2( u2_u7_u6_n156 ) , .ZN( u2_u7_u6_n96 ) );
  AND2_X1 u2_u7_u6_U71 (.A1( u2_u7_X_39 ) , .A2( u2_u7_X_42 ) , .ZN( u2_u7_u6_n99 ) );
  INV_X1 u2_u7_u6_U72 (.A( u2_u7_X_40 ) , .ZN( u2_u7_u6_n157 ) );
  INV_X1 u2_u7_u6_U73 (.A( u2_u7_X_37 ) , .ZN( u2_u7_u6_n165 ) );
  INV_X1 u2_u7_u6_U74 (.A( u2_u7_X_38 ) , .ZN( u2_u7_u6_n162 ) );
  INV_X1 u2_u7_u6_U75 (.A( u2_u7_X_42 ) , .ZN( u2_u7_u6_n156 ) );
  NAND4_X1 u2_u7_u6_U76 (.ZN( u2_out7_12 ) , .A4( u2_u7_u6_n114 ) , .A3( u2_u7_u6_n115 ) , .A2( u2_u7_u6_n116 ) , .A1( u2_u7_u6_n117 ) );
  OAI22_X1 u2_u7_u6_U77 (.B2( u2_u7_u6_n111 ) , .ZN( u2_u7_u6_n116 ) , .B1( u2_u7_u6_n126 ) , .A2( u2_u7_u6_n164 ) , .A1( u2_u7_u6_n167 ) );
  OAI21_X1 u2_u7_u6_U78 (.A( u2_u7_u6_n108 ) , .ZN( u2_u7_u6_n117 ) , .B2( u2_u7_u6_n141 ) , .B1( u2_u7_u6_n163 ) );
  NAND4_X1 u2_u7_u6_U79 (.ZN( u2_out7_32 ) , .A4( u2_u7_u6_n103 ) , .A3( u2_u7_u6_n104 ) , .A2( u2_u7_u6_n105 ) , .A1( u2_u7_u6_n106 ) );
  AOI21_X1 u2_u7_u6_U8 (.B1( u2_u7_u6_n107 ) , .B2( u2_u7_u6_n132 ) , .A( u2_u7_u6_n158 ) , .ZN( u2_u7_u6_n88 ) );
  AOI22_X1 u2_u7_u6_U80 (.ZN( u2_u7_u6_n105 ) , .A2( u2_u7_u6_n108 ) , .A1( u2_u7_u6_n118 ) , .B2( u2_u7_u6_n126 ) , .B1( u2_u7_u6_n171 ) );
  AOI22_X1 u2_u7_u6_U81 (.ZN( u2_u7_u6_n104 ) , .A1( u2_u7_u6_n111 ) , .B1( u2_u7_u6_n124 ) , .B2( u2_u7_u6_n151 ) , .A2( u2_u7_u6_n93 ) );
  OAI211_X1 u2_u7_u6_U82 (.ZN( u2_out7_22 ) , .B( u2_u7_u6_n137 ) , .A( u2_u7_u6_n138 ) , .C2( u2_u7_u6_n139 ) , .C1( u2_u7_u6_n140 ) );
  AOI22_X1 u2_u7_u6_U83 (.B1( u2_u7_u6_n124 ) , .A2( u2_u7_u6_n125 ) , .A1( u2_u7_u6_n126 ) , .ZN( u2_u7_u6_n138 ) , .B2( u2_u7_u6_n161 ) );
  AND4_X1 u2_u7_u6_U84 (.A3( u2_u7_u6_n119 ) , .A1( u2_u7_u6_n120 ) , .A4( u2_u7_u6_n129 ) , .ZN( u2_u7_u6_n140 ) , .A2( u2_u7_u6_n143 ) );
  OAI211_X1 u2_u7_u6_U85 (.ZN( u2_out7_7 ) , .B( u2_u7_u6_n153 ) , .C2( u2_u7_u6_n154 ) , .C1( u2_u7_u6_n155 ) , .A( u2_u7_u6_n174 ) );
  NOR3_X1 u2_u7_u6_U86 (.A1( u2_u7_u6_n141 ) , .ZN( u2_u7_u6_n154 ) , .A3( u2_u7_u6_n164 ) , .A2( u2_u7_u6_n171 ) );
  AOI211_X1 u2_u7_u6_U87 (.B( u2_u7_u6_n149 ) , .A( u2_u7_u6_n150 ) , .C2( u2_u7_u6_n151 ) , .C1( u2_u7_u6_n152 ) , .ZN( u2_u7_u6_n153 ) );
  NAND3_X1 u2_u7_u6_U88 (.A2( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n125 ) , .A1( u2_u7_u6_n130 ) , .A3( u2_u7_u6_n131 ) );
  NAND3_X1 u2_u7_u6_U89 (.A3( u2_u7_u6_n133 ) , .ZN( u2_u7_u6_n141 ) , .A1( u2_u7_u6_n145 ) , .A2( u2_u7_u6_n148 ) );
  AOI21_X1 u2_u7_u6_U9 (.B2( u2_u7_u6_n147 ) , .B1( u2_u7_u6_n148 ) , .ZN( u2_u7_u6_n149 ) , .A( u2_u7_u6_n158 ) );
  NAND3_X1 u2_u7_u6_U90 (.ZN( u2_u7_u6_n101 ) , .A3( u2_u7_u6_n107 ) , .A2( u2_u7_u6_n121 ) , .A1( u2_u7_u6_n127 ) );
  NAND3_X1 u2_u7_u6_U91 (.ZN( u2_u7_u6_n102 ) , .A3( u2_u7_u6_n130 ) , .A2( u2_u7_u6_n145 ) , .A1( u2_u7_u6_n166 ) );
  NAND3_X1 u2_u7_u6_U92 (.A3( u2_u7_u6_n113 ) , .A1( u2_u7_u6_n119 ) , .A2( u2_u7_u6_n123 ) , .ZN( u2_u7_u6_n93 ) );
  NAND3_X1 u2_u7_u6_U93 (.ZN( u2_u7_u6_n142 ) , .A2( u2_u7_u6_n172 ) , .A3( u2_u7_u6_n89 ) , .A1( u2_u7_u6_n90 ) );
  XOR2_X1 u2_u8_U10 (.B( u2_K9_45 ) , .A( u2_R7_30 ) , .Z( u2_u8_X_45 ) );
  XOR2_X1 u2_u8_U15 (.B( u2_K9_40 ) , .A( u2_R7_27 ) , .Z( u2_u8_X_40 ) );
  XOR2_X1 u2_u8_U16 (.B( u2_K9_3 ) , .A( u2_R7_2 ) , .Z( u2_u8_X_3 ) );
  XOR2_X1 u2_u8_U17 (.B( u2_K9_39 ) , .A( u2_R7_26 ) , .Z( u2_u8_X_39 ) );
  XOR2_X1 u2_u8_U22 (.B( u2_K9_34 ) , .A( u2_R7_23 ) , .Z( u2_u8_X_34 ) );
  XOR2_X1 u2_u8_U24 (.B( u2_K9_32 ) , .A( u2_R7_21 ) , .Z( u2_u8_X_32 ) );
  XOR2_X1 u2_u8_U25 (.B( u2_K9_31 ) , .A( u2_R7_20 ) , .Z( u2_u8_X_31 ) );
  XOR2_X1 u2_u8_U26 (.B( u2_K9_30 ) , .A( u2_R7_21 ) , .Z( u2_u8_X_30 ) );
  XOR2_X1 u2_u8_U28 (.B( u2_K9_29 ) , .A( u2_R7_20 ) , .Z( u2_u8_X_29 ) );
  XOR2_X1 u2_u8_U29 (.B( u2_K9_28 ) , .A( u2_R7_19 ) , .Z( u2_u8_X_28 ) );
  XOR2_X1 u2_u8_U30 (.B( u2_K9_27 ) , .A( u2_R7_18 ) , .Z( u2_u8_X_27 ) );
  XOR2_X1 u2_u8_U38 (.B( u2_K9_1 ) , .A( u2_R7_32 ) , .Z( u2_u8_X_1 ) );
  XOR2_X1 u2_u8_U43 (.B( u2_K9_15 ) , .A( u2_R7_10 ) , .Z( u2_u8_X_15 ) );
  XOR2_X1 u2_u8_U8 (.B( u2_K9_47 ) , .A( u2_R7_32 ) , .Z( u2_u8_X_47 ) );
  XOR2_X1 u2_u8_U9 (.B( u2_K9_46 ) , .A( u2_R7_31 ) , .Z( u2_u8_X_46 ) );
  XOR2_X1 u2_u9_U10 (.B( u2_K10_45 ) , .A( u2_R8_30 ) , .Z( u2_u9_X_45 ) );
  XOR2_X1 u2_u9_U16 (.B( u2_K10_3 ) , .A( u2_R8_2 ) , .Z( u2_u9_X_3 ) );
  XOR2_X1 u2_u9_U22 (.B( u2_K10_34 ) , .A( u2_R8_23 ) , .Z( u2_u9_X_34 ) );
  XOR2_X1 u2_u9_U24 (.B( u2_K10_32 ) , .A( u2_R8_21 ) , .Z( u2_u9_X_32 ) );
  XOR2_X1 u2_u9_U26 (.B( u2_K10_30 ) , .A( u2_R8_21 ) , .Z( u2_u9_X_30 ) );
  XOR2_X1 u2_u9_U28 (.B( u2_K10_29 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_29 ) );
  XOR2_X1 u2_u9_U29 (.B( u2_K10_28 ) , .A( u2_R8_19 ) , .Z( u2_u9_X_28 ) );
  XOR2_X1 u2_u9_U30 (.B( u2_K10_27 ) , .A( u2_R8_18 ) , .Z( u2_u9_X_27 ) );
  XOR2_X1 u2_u9_U36 (.B( u2_K10_21 ) , .A( u2_R8_14 ) , .Z( u2_u9_X_21 ) );
  XOR2_X1 u2_u9_U4 (.B( u2_K10_6 ) , .A( u2_R8_5 ) , .Z( u2_u9_X_6 ) );
  XOR2_X1 u2_u9_U42 (.B( u2_K10_16 ) , .A( u2_R8_11 ) , .Z( u2_u9_X_16 ) );
  XOR2_X1 u2_u9_U43 (.B( u2_K10_15 ) , .A( u2_R8_10 ) , .Z( u2_u9_X_15 ) );
  XOR2_X1 u2_u9_U48 (.B( u2_K10_10 ) , .A( u2_R8_7 ) , .Z( u2_u9_X_10 ) );
  XOR2_X1 u2_u9_U6 (.B( u2_K10_4 ) , .A( u2_R8_3 ) , .Z( u2_u9_X_4 ) );
  XOR2_X1 u2_u9_U9 (.B( u2_K10_46 ) , .A( u2_R8_31 ) , .Z( u2_u9_X_46 ) );
  DFF_X1 u2_uk_K_r0_reg_0 (.CK( clk ) , .D( u2_key_r_0 ) , .Q( u2_uk_K_r0_0 ) , .QN( u2_uk_n1230 ) );
  DFF_X1 u2_uk_K_r0_reg_1 (.CK( clk ) , .D( u2_key_r_1 ) , .Q( u2_uk_K_r0_1 ) );
  DFF_X1 u2_uk_K_r0_reg_10 (.CK( clk ) , .D( u2_key_r_10 ) , .Q( u2_uk_K_r0_10 ) , .QN( u2_uk_n1238 ) );
  DFF_X1 u2_uk_K_r0_reg_11 (.CK( clk ) , .D( u2_key_r_11 ) , .Q( u2_uk_K_r0_11 ) );
  DFF_X1 u2_uk_K_r0_reg_12 (.CK( clk ) , .D( u2_key_r_12 ) , .Q( u2_uk_K_r0_12 ) , .QN( u2_uk_n1239 ) );
  DFF_X1 u2_uk_K_r0_reg_13 (.CK( clk ) , .D( u2_key_r_13 ) , .Q( u2_uk_K_r0_13 ) , .QN( u2_uk_n1240 ) );
  DFF_X1 u2_uk_K_r0_reg_14 (.CK( clk ) , .D( u2_key_r_14 ) , .Q( u2_uk_K_r0_14 ) , .QN( u2_uk_n1241 ) );
  DFF_X1 u2_uk_K_r0_reg_15 (.CK( clk ) , .D( u2_key_r_15 ) , .Q( u2_uk_K_r0_15 ) );
  DFF_X1 u2_uk_K_r0_reg_16 (.CK( clk ) , .D( u2_key_r_16 ) , .Q( u2_uk_K_r0_16 ) , .QN( u2_uk_n1242 ) );
  DFF_X1 u2_uk_K_r0_reg_17 (.CK( clk ) , .D( u2_key_r_17 ) , .Q( u2_uk_K_r0_17 ) );
  DFF_X1 u2_uk_K_r0_reg_18 (.CK( clk ) , .D( u2_key_r_18 ) , .Q( u2_uk_K_r0_18 ) , .QN( u2_uk_n1243 ) );
  DFF_X1 u2_uk_K_r0_reg_19 (.CK( clk ) , .D( u2_key_r_19 ) , .Q( u2_uk_K_r0_19 ) );
  DFF_X1 u2_uk_K_r0_reg_2 (.CK( clk ) , .D( u2_key_r_2 ) , .Q( u2_uk_K_r0_2 ) );
  DFF_X1 u2_uk_K_r0_reg_20 (.CK( clk ) , .D( u2_key_r_20 ) , .Q( u2_uk_K_r0_20 ) , .QN( u2_uk_n1244 ) );
  DFF_X1 u2_uk_K_r0_reg_21 (.CK( clk ) , .D( u2_key_r_21 ) , .Q( u2_uk_K_r0_21 ) , .QN( u2_uk_n1245 ) );
  DFF_X1 u2_uk_K_r0_reg_22 (.CK( clk ) , .D( u2_key_r_22 ) , .Q( u2_uk_K_r0_22 ) );
  DFF_X1 u2_uk_K_r0_reg_23 (.CK( clk ) , .D( u2_key_r_23 ) , .Q( u2_uk_K_r0_23 ) , .QN( u2_uk_n1246 ) );
  DFF_X1 u2_uk_K_r0_reg_24 (.CK( clk ) , .D( u2_key_r_24 ) , .Q( u2_uk_K_r0_24 ) , .QN( u2_uk_n1247 ) );
  DFF_X1 u2_uk_K_r0_reg_25 (.CK( clk ) , .D( u2_key_r_25 ) , .Q( u2_uk_K_r0_25 ) );
  DFF_X1 u2_uk_K_r0_reg_26 (.CK( clk ) , .D( u2_key_r_26 ) , .Q( u2_uk_K_r0_26 ) , .QN( u2_uk_n1248 ) );
  DFF_X1 u2_uk_K_r0_reg_27 (.CK( clk ) , .D( u2_key_r_27 ) , .Q( u2_uk_K_r0_27 ) , .QN( u2_uk_n1249 ) );
  DFF_X1 u2_uk_K_r0_reg_28 (.CK( clk ) , .D( u2_key_r_28 ) , .Q( u2_uk_K_r0_28 ) );
  DFF_X1 u2_uk_K_r0_reg_29 (.CK( clk ) , .D( u2_key_r_29 ) , .Q( u2_uk_K_r0_29 ) , .QN( u2_uk_n1251 ) );
  DFF_X1 u2_uk_K_r0_reg_3 (.CK( clk ) , .D( u2_key_r_3 ) , .Q( u2_uk_K_r0_3 ) , .QN( u2_uk_n1231 ) );
  DFF_X1 u2_uk_K_r0_reg_30 (.CK( clk ) , .D( u2_key_r_30 ) , .Q( u2_uk_K_r0_30 ) , .QN( u2_uk_n1252 ) );
  DFF_X1 u2_uk_K_r0_reg_31 (.CK( clk ) , .D( u2_key_r_31 ) , .Q( u2_uk_K_r0_31 ) );
  DFF_X1 u2_uk_K_r0_reg_32 (.CK( clk ) , .D( u2_key_r_32 ) , .Q( u2_uk_K_r0_32 ) );
  DFF_X1 u2_uk_K_r0_reg_33 (.CK( clk ) , .D( u2_key_r_33 ) , .Q( u2_uk_K_r0_33 ) , .QN( u2_uk_n1254 ) );
  DFF_X1 u2_uk_K_r0_reg_34 (.CK( clk ) , .D( u2_key_r_34 ) , .Q( u2_uk_K_r0_34 ) );
  DFF_X1 u2_uk_K_r0_reg_35 (.CK( clk ) , .D( u2_key_r_35 ) , .Q( u2_uk_K_r0_35 ) , .QN( u2_uk_n1256 ) );
  DFF_X1 u2_uk_K_r0_reg_36 (.CK( clk ) , .D( u2_key_r_36 ) , .Q( u2_uk_K_r0_36 ) );
  DFF_X1 u2_uk_K_r0_reg_37 (.CK( clk ) , .D( u2_key_r_37 ) , .Q( u2_uk_K_r0_37 ) , .QN( u2_uk_n1258 ) );
  DFF_X1 u2_uk_K_r0_reg_38 (.CK( clk ) , .D( u2_key_r_38 ) , .Q( u2_uk_K_r0_38 ) , .QN( u2_uk_n1259 ) );
  DFF_X1 u2_uk_K_r0_reg_39 (.CK( clk ) , .D( u2_key_r_39 ) , .Q( u2_uk_K_r0_39 ) , .QN( u2_uk_n1260 ) );
  DFF_X1 u2_uk_K_r0_reg_4 (.CK( clk ) , .D( u2_key_r_4 ) , .Q( u2_uk_K_r0_4 ) , .QN( u2_uk_n1232 ) );
  DFF_X1 u2_uk_K_r0_reg_40 (.CK( clk ) , .D( u2_key_r_40 ) , .Q( u2_uk_K_r0_40 ) , .QN( u2_uk_n1261 ) );
  DFF_X1 u2_uk_K_r0_reg_41 (.CK( clk ) , .D( u2_key_r_41 ) , .Q( u2_uk_K_r0_41 ) , .QN( u2_uk_n1262 ) );
  DFF_X1 u2_uk_K_r0_reg_42 (.CK( clk ) , .D( u2_key_r_42 ) , .Q( u2_uk_K_r0_42 ) , .QN( u2_uk_n1263 ) );
  DFF_X1 u2_uk_K_r0_reg_43 (.CK( clk ) , .D( u2_key_r_43 ) , .Q( u2_uk_K_r0_43 ) , .QN( u2_uk_n1264 ) );
  DFF_X1 u2_uk_K_r0_reg_44 (.CK( clk ) , .D( u2_key_r_44 ) , .Q( u2_uk_K_r0_44 ) , .QN( u2_uk_n1265 ) );
  DFF_X1 u2_uk_K_r0_reg_45 (.CK( clk ) , .D( u2_key_r_45 ) , .Q( u2_uk_K_r0_45 ) , .QN( u2_uk_n1266 ) );
  DFF_X1 u2_uk_K_r0_reg_46 (.CK( clk ) , .D( u2_key_r_46 ) , .Q( u2_uk_K_r0_46 ) , .QN( u2_uk_n1267 ) );
  DFF_X1 u2_uk_K_r0_reg_47 (.CK( clk ) , .D( u2_key_r_47 ) , .Q( u2_uk_K_r0_47 ) , .QN( u2_uk_n1269 ) );
  DFF_X1 u2_uk_K_r0_reg_48 (.CK( clk ) , .D( u2_key_r_48 ) , .Q( u2_uk_K_r0_48 ) , .QN( u2_uk_n1270 ) );
  DFF_X1 u2_uk_K_r0_reg_49 (.CK( clk ) , .D( u2_key_r_49 ) , .Q( u2_uk_K_r0_49 ) );
  DFF_X1 u2_uk_K_r0_reg_5 (.CK( clk ) , .D( u2_key_r_5 ) , .Q( u2_uk_K_r0_5 ) , .QN( u2_uk_n1233 ) );
  DFF_X1 u2_uk_K_r0_reg_50 (.CK( clk ) , .D( u2_key_r_50 ) , .Q( u2_uk_K_r0_50 ) , .QN( u2_uk_n1273 ) );
  DFF_X1 u2_uk_K_r0_reg_51 (.CK( clk ) , .D( u2_key_r_51 ) , .Q( u2_uk_K_r0_51 ) , .QN( u2_uk_n1274 ) );
  DFF_X1 u2_uk_K_r0_reg_52 (.CK( clk ) , .D( u2_key_r_52 ) , .Q( u2_uk_K_r0_52 ) );
  DFF_X1 u2_uk_K_r0_reg_53 (.CK( clk ) , .D( u2_key_r_53 ) , .Q( u2_uk_K_r0_53 ) );
  DFF_X1 u2_uk_K_r0_reg_54 (.CK( clk ) , .D( u2_key_r_54 ) , .Q( u2_uk_K_r0_54 ) , .QN( u2_uk_n1275 ) );
  DFF_X1 u2_uk_K_r0_reg_55 (.CK( clk ) , .D( u2_key_r_55 ) , .Q( u2_uk_K_r0_55 ) );
  DFF_X1 u2_uk_K_r0_reg_6 (.CK( clk ) , .D( u2_key_r_6 ) , .Q( u2_uk_K_r0_6 ) , .QN( u2_uk_n1234 ) );
  DFF_X1 u2_uk_K_r0_reg_7 (.CK( clk ) , .D( u2_key_r_7 ) , .Q( u2_uk_K_r0_7 ) , .QN( u2_uk_n1235 ) );
  DFF_X1 u2_uk_K_r0_reg_8 (.CK( clk ) , .D( u2_key_r_8 ) , .Q( u2_uk_K_r0_8 ) , .QN( u2_uk_n1236 ) );
  DFF_X1 u2_uk_K_r0_reg_9 (.CK( clk ) , .D( u2_key_r_9 ) , .Q( u2_uk_K_r0_9 ) , .QN( u2_uk_n1237 ) );
  DFF_X1 u2_uk_K_r10_reg_0 (.CK( clk ) , .Q( u2_uk_K_r10_0 ) , .D( u2_uk_K_r9_0 ) , .QN( u2_uk_n1678 ) );
  DFF_X1 u2_uk_K_r10_reg_1 (.CK( clk ) , .Q( u2_uk_K_r10_1 ) , .D( u2_uk_K_r9_1 ) , .QN( u2_uk_n1679 ) );
  DFF_X1 u2_uk_K_r10_reg_10 (.CK( clk ) , .Q( u2_uk_K_r10_10 ) , .D( u2_uk_K_r9_10 ) );
  DFF_X1 u2_uk_K_r10_reg_11 (.CK( clk ) , .Q( u2_uk_K_r10_11 ) , .D( u2_uk_K_r9_11 ) );
  DFF_X1 u2_uk_K_r10_reg_12 (.CK( clk ) , .Q( u2_uk_K_r10_12 ) , .D( u2_uk_K_r9_12 ) , .QN( u2_uk_n1686 ) );
  DFF_X1 u2_uk_K_r10_reg_13 (.CK( clk ) , .Q( u2_uk_K_r10_13 ) , .D( u2_uk_K_r9_13 ) );
  DFF_X1 u2_uk_K_r10_reg_14 (.CK( clk ) , .Q( u2_uk_K_r10_14 ) , .D( u2_uk_K_r9_14 ) );
  DFF_X1 u2_uk_K_r10_reg_15 (.CK( clk ) , .Q( u2_uk_K_r10_15 ) , .D( u2_uk_K_r9_15 ) , .QN( u2_uk_n1687 ) );
  DFF_X1 u2_uk_K_r10_reg_16 (.CK( clk ) , .Q( u2_uk_K_r10_16 ) , .D( u2_uk_K_r9_16 ) );
  DFF_X1 u2_uk_K_r10_reg_17 (.CK( clk ) , .Q( u2_uk_K_r10_17 ) , .D( u2_uk_K_r9_17 ) , .QN( u2_uk_n1688 ) );
  DFF_X1 u2_uk_K_r10_reg_18 (.CK( clk ) , .Q( u2_uk_K_r10_18 ) , .D( u2_uk_K_r9_18 ) );
  DFF_X1 u2_uk_K_r10_reg_19 (.CK( clk ) , .Q( u2_uk_K_r10_19 ) , .D( u2_uk_K_r9_19 ) );
  DFF_X1 u2_uk_K_r10_reg_2 (.CK( clk ) , .Q( u2_uk_K_r10_2 ) , .D( u2_uk_K_r9_2 ) , .QN( u2_uk_n1680 ) );
  DFF_X1 u2_uk_K_r10_reg_20 (.CK( clk ) , .Q( u2_uk_K_r10_20 ) , .D( u2_uk_K_r9_20 ) , .QN( u2_uk_n1689 ) );
  DFF_X1 u2_uk_K_r10_reg_21 (.CK( clk ) , .Q( u2_uk_K_r10_21 ) , .D( u2_uk_K_r9_21 ) , .QN( u2_uk_n1690 ) );
  DFF_X1 u2_uk_K_r10_reg_22 (.CK( clk ) , .Q( u2_uk_K_r10_22 ) , .D( u2_uk_K_r9_22 ) , .QN( u2_uk_n1691 ) );
  DFF_X1 u2_uk_K_r10_reg_23 (.CK( clk ) , .Q( u2_uk_K_r10_23 ) , .D( u2_uk_K_r9_23 ) );
  DFF_X1 u2_uk_K_r10_reg_24 (.CK( clk ) , .Q( u2_uk_K_r10_24 ) , .D( u2_uk_K_r9_24 ) , .QN( u2_uk_n1692 ) );
  DFF_X1 u2_uk_K_r10_reg_25 (.CK( clk ) , .Q( u2_uk_K_r10_25 ) , .D( u2_uk_K_r9_25 ) );
  DFF_X1 u2_uk_K_r10_reg_26 (.CK( clk ) , .Q( u2_uk_K_r10_26 ) , .D( u2_uk_K_r9_26 ) , .QN( u2_uk_n1693 ) );
  DFF_X1 u2_uk_K_r10_reg_27 (.CK( clk ) , .Q( u2_uk_K_r10_27 ) , .D( u2_uk_K_r9_27 ) );
  DFF_X1 u2_uk_K_r10_reg_28 (.CK( clk ) , .Q( u2_uk_K_r10_28 ) , .D( u2_uk_K_r9_28 ) );
  DFF_X1 u2_uk_K_r10_reg_29 (.CK( clk ) , .Q( u2_uk_K_r10_29 ) , .D( u2_uk_K_r9_29 ) , .QN( u2_uk_n1698 ) );
  DFF_X1 u2_uk_K_r10_reg_3 (.CK( clk ) , .Q( u2_uk_K_r10_3 ) , .D( u2_uk_K_r9_3 ) , .QN( u2_uk_n1681 ) );
  DFF_X1 u2_uk_K_r10_reg_30 (.CK( clk ) , .Q( u2_uk_K_r10_30 ) , .D( u2_uk_K_r9_30 ) , .QN( u2_uk_n1699 ) );
  DFF_X1 u2_uk_K_r10_reg_31 (.CK( clk ) , .Q( u2_uk_K_r10_31 ) , .D( u2_uk_K_r9_31 ) , .QN( u2_uk_n1700 ) );
  DFF_X1 u2_uk_K_r10_reg_32 (.CK( clk ) , .Q( u2_uk_K_r10_32 ) , .D( u2_uk_K_r9_32 ) , .QN( u2_uk_n1701 ) );
  DFF_X1 u2_uk_K_r10_reg_33 (.CK( clk ) , .Q( u2_uk_K_r10_33 ) , .D( u2_uk_K_r9_33 ) , .QN( u2_uk_n1702 ) );
  DFF_X1 u2_uk_K_r10_reg_34 (.CK( clk ) , .Q( u2_uk_K_r10_34 ) , .D( u2_uk_K_r9_34 ) );
  DFF_X1 u2_uk_K_r10_reg_35 (.CK( clk ) , .Q( u2_uk_K_r10_35 ) , .D( u2_uk_K_r9_35 ) , .QN( u2_uk_n1704 ) );
  DFF_X1 u2_uk_K_r10_reg_36 (.CK( clk ) , .Q( u2_uk_K_r10_36 ) , .D( u2_uk_K_r9_36 ) , .QN( u2_uk_n1705 ) );
  DFF_X1 u2_uk_K_r10_reg_37 (.CK( clk ) , .Q( u2_uk_K_r10_37 ) , .D( u2_uk_K_r9_37 ) , .QN( u2_uk_n1706 ) );
  DFF_X1 u2_uk_K_r10_reg_38 (.CK( clk ) , .Q( u2_uk_K_r10_38 ) , .D( u2_uk_K_r9_38 ) , .QN( u2_uk_n1707 ) );
  DFF_X1 u2_uk_K_r10_reg_39 (.CK( clk ) , .Q( u2_uk_K_r10_39 ) , .D( u2_uk_K_r9_39 ) , .QN( u2_uk_n1708 ) );
  DFF_X1 u2_uk_K_r10_reg_4 (.CK( clk ) , .Q( u2_uk_K_r10_4 ) , .D( u2_uk_K_r9_4 ) );
  DFF_X1 u2_uk_K_r10_reg_40 (.CK( clk ) , .Q( u2_uk_K_r10_40 ) , .D( u2_uk_K_r9_40 ) , .QN( u2_uk_n1709 ) );
  DFF_X1 u2_uk_K_r10_reg_41 (.CK( clk ) , .Q( u2_uk_K_r10_41 ) , .D( u2_uk_K_r9_41 ) );
  DFF_X1 u2_uk_K_r10_reg_42 (.CK( clk ) , .Q( u2_uk_K_r10_42 ) , .D( u2_uk_K_r9_42 ) );
  DFF_X1 u2_uk_K_r10_reg_43 (.CK( clk ) , .Q( u2_uk_K_r10_43 ) , .D( u2_uk_K_r9_43 ) );
  DFF_X1 u2_uk_K_r10_reg_44 (.CK( clk ) , .Q( u2_uk_K_r10_44 ) , .D( u2_uk_K_r9_44 ) );
  DFF_X1 u2_uk_K_r10_reg_45 (.CK( clk ) , .Q( u2_uk_K_r10_45 ) , .D( u2_uk_K_r9_45 ) , .QN( u2_uk_n1714 ) );
  DFF_X1 u2_uk_K_r10_reg_46 (.CK( clk ) , .Q( u2_uk_K_r10_46 ) , .D( u2_uk_K_r9_46 ) , .QN( u2_uk_n1715 ) );
  DFF_X1 u2_uk_K_r10_reg_47 (.CK( clk ) , .Q( u2_uk_K_r10_47 ) , .D( u2_uk_K_r9_47 ) );
  DFF_X1 u2_uk_K_r10_reg_48 (.CK( clk ) , .Q( u2_uk_K_r10_48 ) , .D( u2_uk_K_r9_48 ) );
  DFF_X1 u2_uk_K_r10_reg_49 (.CK( clk ) , .Q( u2_uk_K_r10_49 ) , .D( u2_uk_K_r9_49 ) );
  DFF_X1 u2_uk_K_r10_reg_5 (.CK( clk ) , .Q( u2_uk_K_r10_5 ) , .D( u2_uk_K_r9_5 ) , .QN( u2_uk_n1682 ) );
  DFF_X1 u2_uk_K_r10_reg_50 (.CK( clk ) , .Q( u2_uk_K_r10_50 ) , .D( u2_uk_K_r9_50 ) , .QN( u2_uk_n1718 ) );
  DFF_X1 u2_uk_K_r10_reg_51 (.CK( clk ) , .Q( u2_uk_K_r10_51 ) , .D( u2_uk_K_r9_51 ) , .QN( u2_uk_n1719 ) );
  DFF_X1 u2_uk_K_r10_reg_52 (.CK( clk ) , .Q( u2_uk_K_r10_52 ) , .D( u2_uk_K_r9_52 ) );
  DFF_X1 u2_uk_K_r10_reg_53 (.CK( clk ) , .Q( u2_uk_K_r10_53 ) , .D( u2_uk_K_r9_53 ) , .QN( u2_uk_n1720 ) );
  DFF_X1 u2_uk_K_r10_reg_54 (.CK( clk ) , .Q( u2_uk_K_r10_54 ) , .D( u2_uk_K_r9_54 ) , .QN( u2_uk_n1721 ) );
  DFF_X1 u2_uk_K_r10_reg_55 (.CK( clk ) , .Q( u2_uk_K_r10_55 ) , .D( u2_uk_K_r9_55 ) , .QN( u2_uk_n1722 ) );
  DFF_X1 u2_uk_K_r10_reg_6 (.CK( clk ) , .Q( u2_uk_K_r10_6 ) , .D( u2_uk_K_r9_6 ) , .QN( u2_uk_n1683 ) );
  DFF_X1 u2_uk_K_r10_reg_7 (.CK( clk ) , .Q( u2_uk_K_r10_7 ) , .D( u2_uk_K_r9_7 ) , .QN( u2_uk_n1684 ) );
  DFF_X1 u2_uk_K_r10_reg_8 (.CK( clk ) , .Q( u2_uk_K_r10_8 ) , .D( u2_uk_K_r9_8 ) , .QN( u2_uk_n1685 ) );
  DFF_X1 u2_uk_K_r10_reg_9 (.CK( clk ) , .Q( u2_uk_K_r10_9 ) , .D( u2_uk_K_r9_9 ) );
  DFF_X1 u2_uk_K_r11_reg_0 (.CK( clk ) , .D( u2_uk_K_r10_0 ) , .Q( u2_uk_K_r11_0 ) , .QN( u2_uk_n1723 ) );
  DFF_X1 u2_uk_K_r11_reg_1 (.CK( clk ) , .D( u2_uk_K_r10_1 ) , .Q( u2_uk_K_r11_1 ) , .QN( u2_uk_n1724 ) );
  DFF_X1 u2_uk_K_r11_reg_10 (.CK( clk ) , .D( u2_uk_K_r10_10 ) , .Q( u2_uk_K_r11_10 ) );
  DFF_X1 u2_uk_K_r11_reg_11 (.CK( clk ) , .D( u2_uk_K_r10_11 ) , .Q( u2_uk_K_r11_11 ) );
  DFF_X1 u2_uk_K_r11_reg_12 (.CK( clk ) , .D( u2_uk_K_r10_12 ) , .Q( u2_uk_K_r11_12 ) , .QN( u2_uk_n1731 ) );
  DFF_X1 u2_uk_K_r11_reg_13 (.CK( clk ) , .D( u2_uk_K_r10_13 ) , .Q( u2_uk_K_r11_13 ) , .QN( u2_uk_n1732 ) );
  DFF_X1 u2_uk_K_r11_reg_14 (.CK( clk ) , .D( u2_uk_K_r10_14 ) , .Q( u2_uk_K_r11_14 ) , .QN( u2_uk_n1733 ) );
  DFF_X1 u2_uk_K_r11_reg_15 (.CK( clk ) , .D( u2_uk_K_r10_15 ) , .Q( u2_uk_K_r11_15 ) , .QN( u2_uk_n1734 ) );
  DFF_X1 u2_uk_K_r11_reg_16 (.CK( clk ) , .D( u2_uk_K_r10_16 ) , .Q( u2_uk_K_r11_16 ) , .QN( u2_uk_n1735 ) );
  DFF_X1 u2_uk_K_r11_reg_17 (.CK( clk ) , .D( u2_uk_K_r10_17 ) , .Q( u2_uk_K_r11_17 ) , .QN( u2_uk_n1736 ) );
  DFF_X1 u2_uk_K_r11_reg_18 (.CK( clk ) , .D( u2_uk_K_r10_18 ) , .Q( u2_uk_K_r11_18 ) , .QN( u2_uk_n1737 ) );
  DFF_X1 u2_uk_K_r11_reg_19 (.CK( clk ) , .D( u2_uk_K_r10_19 ) , .Q( u2_uk_K_r11_19 ) );
  DFF_X1 u2_uk_K_r11_reg_2 (.CK( clk ) , .D( u2_uk_K_r10_2 ) , .Q( u2_uk_K_r11_2 ) , .QN( u2_uk_n1725 ) );
  DFF_X1 u2_uk_K_r11_reg_20 (.CK( clk ) , .D( u2_uk_K_r10_20 ) , .Q( u2_uk_K_r11_20 ) );
  DFF_X1 u2_uk_K_r11_reg_21 (.CK( clk ) , .D( u2_uk_K_r10_21 ) , .Q( u2_uk_K_r11_21 ) );
  DFF_X1 u2_uk_K_r11_reg_22 (.CK( clk ) , .D( u2_uk_K_r10_22 ) , .Q( u2_uk_K_r11_22 ) , .QN( u2_uk_n1738 ) );
  DFF_X1 u2_uk_K_r11_reg_23 (.CK( clk ) , .D( u2_uk_K_r10_23 ) , .Q( u2_uk_K_r11_23 ) , .QN( u2_uk_n1739 ) );
  DFF_X1 u2_uk_K_r11_reg_24 (.CK( clk ) , .D( u2_uk_K_r10_24 ) , .Q( u2_uk_K_r11_24 ) );
  DFF_X1 u2_uk_K_r11_reg_25 (.CK( clk ) , .D( u2_uk_K_r10_25 ) , .Q( u2_uk_K_r11_25 ) );
  DFF_X1 u2_uk_K_r11_reg_26 (.CK( clk ) , .D( u2_uk_K_r10_26 ) , .Q( u2_uk_K_r11_26 ) );
  DFF_X1 u2_uk_K_r11_reg_27 (.CK( clk ) , .D( u2_uk_K_r10_27 ) , .Q( u2_uk_K_r11_27 ) );
  DFF_X1 u2_uk_K_r11_reg_28 (.CK( clk ) , .D( u2_uk_K_r10_28 ) , .Q( u2_uk_K_r11_28 ) );
  DFF_X1 u2_uk_K_r11_reg_29 (.CK( clk ) , .D( u2_uk_K_r10_29 ) , .Q( u2_uk_K_r11_29 ) );
  DFF_X1 u2_uk_K_r11_reg_3 (.CK( clk ) , .D( u2_uk_K_r10_3 ) , .Q( u2_uk_K_r11_3 ) , .QN( u2_uk_n1726 ) );
  DFF_X1 u2_uk_K_r11_reg_30 (.CK( clk ) , .D( u2_uk_K_r10_30 ) , .Q( u2_uk_K_r11_30 ) );
  DFF_X1 u2_uk_K_r11_reg_31 (.CK( clk ) , .D( u2_uk_K_r10_31 ) , .Q( u2_uk_K_r11_31 ) , .QN( u2_uk_n1742 ) );
  DFF_X1 u2_uk_K_r11_reg_32 (.CK( clk ) , .D( u2_uk_K_r10_32 ) , .Q( u2_uk_K_r11_32 ) , .QN( u2_uk_n1743 ) );
  DFF_X1 u2_uk_K_r11_reg_33 (.CK( clk ) , .D( u2_uk_K_r10_33 ) , .Q( u2_uk_K_r11_33 ) );
  DFF_X1 u2_uk_K_r11_reg_34 (.CK( clk ) , .D( u2_uk_K_r10_34 ) , .Q( u2_uk_K_r11_34 ) );
  DFF_X1 u2_uk_K_r11_reg_35 (.CK( clk ) , .D( u2_uk_K_r10_35 ) , .Q( u2_uk_K_r11_35 ) , .QN( u2_uk_n1744 ) );
  DFF_X1 u2_uk_K_r11_reg_36 (.CK( clk ) , .D( u2_uk_K_r10_36 ) , .Q( u2_uk_K_r11_36 ) , .QN( u2_uk_n1745 ) );
  DFF_X1 u2_uk_K_r11_reg_37 (.CK( clk ) , .D( u2_uk_K_r10_37 ) , .Q( u2_uk_K_r11_37 ) , .QN( u2_uk_n1746 ) );
  DFF_X1 u2_uk_K_r11_reg_38 (.CK( clk ) , .D( u2_uk_K_r10_38 ) , .Q( u2_uk_K_r11_38 ) , .QN( u2_uk_n1747 ) );
  DFF_X1 u2_uk_K_r11_reg_39 (.CK( clk ) , .D( u2_uk_K_r10_39 ) , .Q( u2_uk_K_r11_39 ) );
  DFF_X1 u2_uk_K_r11_reg_4 (.CK( clk ) , .D( u2_uk_K_r10_4 ) , .Q( u2_uk_K_r11_4 ) );
  DFF_X1 u2_uk_K_r11_reg_40 (.CK( clk ) , .D( u2_uk_K_r10_40 ) , .Q( u2_uk_K_r11_40 ) , .QN( u2_uk_n1750 ) );
  DFF_X1 u2_uk_K_r11_reg_41 (.CK( clk ) , .D( u2_uk_K_r10_41 ) , .Q( u2_uk_K_r11_41 ) , .QN( u2_uk_n1751 ) );
  DFF_X1 u2_uk_K_r11_reg_42 (.CK( clk ) , .D( u2_uk_K_r10_42 ) , .Q( u2_uk_K_r11_42 ) , .QN( u2_uk_n1752 ) );
  DFF_X1 u2_uk_K_r11_reg_43 (.CK( clk ) , .D( u2_uk_K_r10_43 ) , .Q( u2_uk_K_r11_43 ) , .QN( u2_uk_n1753 ) );
  DFF_X1 u2_uk_K_r11_reg_44 (.CK( clk ) , .D( u2_uk_K_r10_44 ) , .Q( u2_uk_K_r11_44 ) , .QN( u2_uk_n1754 ) );
  DFF_X1 u2_uk_K_r11_reg_45 (.CK( clk ) , .D( u2_uk_K_r10_45 ) , .Q( u2_uk_K_r11_45 ) , .QN( u2_uk_n1755 ) );
  DFF_X1 u2_uk_K_r11_reg_46 (.CK( clk ) , .D( u2_uk_K_r10_46 ) , .Q( u2_uk_K_r11_46 ) , .QN( u2_uk_n1757 ) );
  DFF_X1 u2_uk_K_r11_reg_47 (.CK( clk ) , .D( u2_uk_K_r10_47 ) , .Q( u2_uk_K_r11_47 ) );
  DFF_X1 u2_uk_K_r11_reg_48 (.CK( clk ) , .D( u2_uk_K_r10_48 ) , .Q( u2_uk_K_r11_48 ) );
  DFF_X1 u2_uk_K_r11_reg_49 (.CK( clk ) , .D( u2_uk_K_r10_49 ) , .Q( u2_uk_K_r11_49 ) , .QN( u2_uk_n1760 ) );
  DFF_X1 u2_uk_K_r11_reg_5 (.CK( clk ) , .D( u2_uk_K_r10_5 ) , .Q( u2_uk_K_r11_5 ) , .QN( u2_uk_n1727 ) );
  DFF_X1 u2_uk_K_r11_reg_50 (.CK( clk ) , .D( u2_uk_K_r10_50 ) , .Q( u2_uk_K_r11_50 ) , .QN( u2_uk_n1761 ) );
  DFF_X1 u2_uk_K_r11_reg_51 (.CK( clk ) , .D( u2_uk_K_r10_51 ) , .Q( u2_uk_K_r11_51 ) , .QN( u2_uk_n1762 ) );
  DFF_X1 u2_uk_K_r11_reg_52 (.CK( clk ) , .D( u2_uk_K_r10_52 ) , .Q( u2_uk_K_r11_52 ) , .QN( u2_uk_n1763 ) );
  DFF_X1 u2_uk_K_r11_reg_53 (.CK( clk ) , .D( u2_uk_K_r10_53 ) , .Q( u2_uk_K_r11_53 ) );
  DFF_X1 u2_uk_K_r11_reg_54 (.CK( clk ) , .D( u2_uk_K_r10_54 ) , .Q( u2_uk_K_r11_54 ) );
  DFF_X1 u2_uk_K_r11_reg_55 (.CK( clk ) , .D( u2_uk_K_r10_55 ) , .Q( u2_uk_K_r11_55 ) , .QN( u2_uk_n1767 ) );
  DFF_X1 u2_uk_K_r11_reg_6 (.CK( clk ) , .D( u2_uk_K_r10_6 ) , .Q( u2_uk_K_r11_6 ) );
  DFF_X1 u2_uk_K_r11_reg_7 (.CK( clk ) , .D( u2_uk_K_r10_7 ) , .Q( u2_uk_K_r11_7 ) );
  DFF_X1 u2_uk_K_r11_reg_8 (.CK( clk ) , .D( u2_uk_K_r10_8 ) , .Q( u2_uk_K_r11_8 ) );
  DFF_X1 u2_uk_K_r11_reg_9 (.CK( clk ) , .D( u2_uk_K_r10_9 ) , .Q( u2_uk_K_r11_9 ) , .QN( u2_uk_n1728 ) );
  DFF_X1 u2_uk_K_r12_reg_0 (.CK( clk ) , .D( u2_uk_K_r11_0 ) , .Q( u2_uk_K_r12_0 ) , .QN( u2_uk_n1768 ) );
  DFF_X1 u2_uk_K_r12_reg_1 (.CK( clk ) , .D( u2_uk_K_r11_1 ) , .Q( u2_uk_K_r12_1 ) , .QN( u2_uk_n1769 ) );
  DFF_X1 u2_uk_K_r12_reg_10 (.CK( clk ) , .D( u2_uk_K_r11_10 ) , .Q( u2_uk_K_r12_10 ) );
  DFF_X1 u2_uk_K_r12_reg_11 (.CK( clk ) , .D( u2_uk_K_r11_11 ) , .Q( u2_uk_K_r12_11 ) , .QN( u2_uk_n1778 ) );
  DFF_X1 u2_uk_K_r12_reg_12 (.CK( clk ) , .D( u2_uk_K_r11_12 ) , .Q( u2_uk_K_r12_12 ) , .QN( u2_uk_n1779 ) );
  DFF_X1 u2_uk_K_r12_reg_13 (.CK( clk ) , .D( u2_uk_K_r11_13 ) , .Q( u2_uk_K_r12_13 ) , .QN( u2_uk_n1780 ) );
  DFF_X1 u2_uk_K_r12_reg_14 (.CK( clk ) , .D( u2_uk_K_r11_14 ) , .Q( u2_uk_K_r12_14 ) , .QN( u2_uk_n1781 ) );
  DFF_X1 u2_uk_K_r12_reg_15 (.CK( clk ) , .D( u2_uk_K_r11_15 ) , .Q( u2_uk_K_r12_15 ) );
  DFF_X1 u2_uk_K_r12_reg_16 (.CK( clk ) , .D( u2_uk_K_r11_16 ) , .Q( u2_uk_K_r12_16 ) );
  DFF_X1 u2_uk_K_r12_reg_17 (.CK( clk ) , .D( u2_uk_K_r11_17 ) , .Q( u2_uk_K_r12_17 ) , .QN( u2_uk_n1782 ) );
  DFF_X1 u2_uk_K_r12_reg_18 (.CK( clk ) , .D( u2_uk_K_r11_18 ) , .Q( u2_uk_K_r12_18 ) );
  DFF_X1 u2_uk_K_r12_reg_19 (.CK( clk ) , .D( u2_uk_K_r11_19 ) , .Q( u2_uk_K_r12_19 ) , .QN( u2_uk_n1783 ) );
  DFF_X1 u2_uk_K_r12_reg_2 (.CK( clk ) , .D( u2_uk_K_r11_2 ) , .Q( u2_uk_K_r12_2 ) , .QN( u2_uk_n1770 ) );
  DFF_X1 u2_uk_K_r12_reg_20 (.CK( clk ) , .D( u2_uk_K_r11_20 ) , .Q( u2_uk_K_r12_20 ) , .QN( u2_uk_n1784 ) );
  DFF_X1 u2_uk_K_r12_reg_21 (.CK( clk ) , .D( u2_uk_K_r11_21 ) , .Q( u2_uk_K_r12_21 ) );
  DFF_X1 u2_uk_K_r12_reg_22 (.CK( clk ) , .D( u2_uk_K_r11_22 ) , .Q( u2_uk_K_r12_22 ) );
  DFF_X1 u2_uk_K_r12_reg_23 (.CK( clk ) , .D( u2_uk_K_r11_23 ) , .Q( u2_uk_K_r12_23 ) , .QN( u2_uk_n1785 ) );
  DFF_X1 u2_uk_K_r12_reg_24 (.CK( clk ) , .D( u2_uk_K_r11_24 ) , .Q( u2_uk_K_r12_24 ) , .QN( u2_uk_n1786 ) );
  DFF_X1 u2_uk_K_r12_reg_25 (.CK( clk ) , .D( u2_uk_K_r11_25 ) , .Q( u2_uk_K_r12_25 ) , .QN( u2_uk_n1787 ) );
  DFF_X1 u2_uk_K_r12_reg_26 (.CK( clk ) , .D( u2_uk_K_r11_26 ) , .Q( u2_uk_K_r12_26 ) , .QN( u2_uk_n1788 ) );
  DFF_X1 u2_uk_K_r12_reg_27 (.CK( clk ) , .D( u2_uk_K_r11_27 ) , .Q( u2_uk_K_r12_27 ) , .QN( u2_uk_n1789 ) );
  DFF_X1 u2_uk_K_r12_reg_28 (.CK( clk ) , .D( u2_uk_K_r11_28 ) , .Q( u2_uk_K_r12_28 ) , .QN( u2_uk_n1790 ) );
  DFF_X1 u2_uk_K_r12_reg_29 (.CK( clk ) , .D( u2_uk_K_r11_29 ) , .Q( u2_uk_K_r12_29 ) , .QN( u2_uk_n1791 ) );
  DFF_X1 u2_uk_K_r12_reg_3 (.CK( clk ) , .D( u2_uk_K_r11_3 ) , .Q( u2_uk_K_r12_3 ) , .QN( u2_uk_n1771 ) );
  DFF_X1 u2_uk_K_r12_reg_30 (.CK( clk ) , .D( u2_uk_K_r11_30 ) , .Q( u2_uk_K_r12_30 ) , .QN( u2_uk_n1792 ) );
  DFF_X1 u2_uk_K_r12_reg_31 (.CK( clk ) , .D( u2_uk_K_r11_31 ) , .Q( u2_uk_K_r12_31 ) , .QN( u2_uk_n1793 ) );
  DFF_X1 u2_uk_K_r12_reg_32 (.CK( clk ) , .D( u2_uk_K_r11_32 ) , .Q( u2_uk_K_r12_32 ) , .QN( u2_uk_n1794 ) );
  DFF_X1 u2_uk_K_r12_reg_33 (.CK( clk ) , .D( u2_uk_K_r11_33 ) , .Q( u2_uk_K_r12_33 ) );
  DFF_X1 u2_uk_K_r12_reg_34 (.CK( clk ) , .D( u2_uk_K_r11_34 ) , .Q( u2_uk_K_r12_34 ) , .QN( u2_uk_n1796 ) );
  DFF_X1 u2_uk_K_r12_reg_35 (.CK( clk ) , .D( u2_uk_K_r11_35 ) , .Q( u2_uk_K_r12_35 ) , .QN( u2_uk_n1797 ) );
  DFF_X1 u2_uk_K_r12_reg_36 (.CK( clk ) , .D( u2_uk_K_r11_36 ) , .Q( u2_uk_K_r12_36 ) );
  DFF_X1 u2_uk_K_r12_reg_37 (.CK( clk ) , .D( u2_uk_K_r11_37 ) , .Q( u2_uk_K_r12_37 ) , .QN( u2_uk_n1799 ) );
  DFF_X1 u2_uk_K_r12_reg_38 (.CK( clk ) , .D( u2_uk_K_r11_38 ) , .Q( u2_uk_K_r12_38 ) , .QN( u2_uk_n1800 ) );
  DFF_X1 u2_uk_K_r12_reg_39 (.CK( clk ) , .D( u2_uk_K_r11_39 ) , .Q( u2_uk_K_r12_39 ) );
  DFF_X1 u2_uk_K_r12_reg_4 (.CK( clk ) , .D( u2_uk_K_r11_4 ) , .Q( u2_uk_K_r12_4 ) , .QN( u2_uk_n1772 ) );
  DFF_X1 u2_uk_K_r12_reg_40 (.CK( clk ) , .D( u2_uk_K_r11_40 ) , .Q( u2_uk_K_r12_40 ) , .QN( u2_uk_n1801 ) );
  DFF_X1 u2_uk_K_r12_reg_41 (.CK( clk ) , .D( u2_uk_K_r11_41 ) , .Q( u2_uk_K_r12_41 ) );
  DFF_X1 u2_uk_K_r12_reg_42 (.CK( clk ) , .D( u2_uk_K_r11_42 ) , .Q( u2_uk_K_r12_42 ) );
  DFF_X1 u2_uk_K_r12_reg_43 (.CK( clk ) , .D( u2_uk_K_r11_43 ) , .Q( u2_uk_K_r12_43 ) , .QN( u2_uk_n1802 ) );
  DFF_X1 u2_uk_K_r12_reg_44 (.CK( clk ) , .D( u2_uk_K_r11_44 ) , .Q( u2_uk_K_r12_44 ) );
  DFF_X1 u2_uk_K_r12_reg_45 (.CK( clk ) , .D( u2_uk_K_r11_45 ) , .Q( u2_uk_K_r12_45 ) , .QN( u2_uk_n1803 ) );
  DFF_X1 u2_uk_K_r12_reg_46 (.CK( clk ) , .D( u2_uk_K_r11_46 ) , .Q( u2_uk_K_r12_46 ) , .QN( u2_uk_n1804 ) );
  DFF_X1 u2_uk_K_r12_reg_47 (.CK( clk ) , .D( u2_uk_K_r11_47 ) , .Q( u2_uk_K_r12_47 ) );
  DFF_X1 u2_uk_K_r12_reg_48 (.CK( clk ) , .D( u2_uk_K_r11_48 ) , .Q( u2_uk_K_r12_48 ) , .QN( u2_uk_n1805 ) );
  DFF_X1 u2_uk_K_r12_reg_49 (.CK( clk ) , .D( u2_uk_K_r11_49 ) , .Q( u2_uk_K_r12_49 ) , .QN( u2_uk_n1806 ) );
  DFF_X1 u2_uk_K_r12_reg_5 (.CK( clk ) , .D( u2_uk_K_r11_5 ) , .Q( u2_uk_K_r12_5 ) , .QN( u2_uk_n1773 ) );
  DFF_X1 u2_uk_K_r12_reg_50 (.CK( clk ) , .D( u2_uk_K_r11_50 ) , .Q( u2_uk_K_r12_50 ) , .QN( u2_uk_n1807 ) );
  DFF_X1 u2_uk_K_r12_reg_51 (.CK( clk ) , .D( u2_uk_K_r11_51 ) , .Q( u2_uk_K_r12_51 ) , .QN( u2_uk_n1808 ) );
  DFF_X1 u2_uk_K_r12_reg_52 (.CK( clk ) , .D( u2_uk_K_r11_52 ) , .Q( u2_uk_K_r12_52 ) , .QN( u2_uk_n1809 ) );
  DFF_X1 u2_uk_K_r12_reg_53 (.CK( clk ) , .D( u2_uk_K_r11_53 ) , .Q( u2_uk_K_r12_53 ) , .QN( u2_uk_n1810 ) );
  DFF_X1 u2_uk_K_r12_reg_54 (.CK( clk ) , .D( u2_uk_K_r11_54 ) , .Q( u2_uk_K_r12_54 ) , .QN( u2_uk_n1811 ) );
  DFF_X1 u2_uk_K_r12_reg_55 (.CK( clk ) , .D( u2_uk_K_r11_55 ) , .Q( u2_uk_K_r12_55 ) , .QN( u2_uk_n1812 ) );
  DFF_X1 u2_uk_K_r12_reg_6 (.CK( clk ) , .D( u2_uk_K_r11_6 ) , .Q( u2_uk_K_r12_6 ) , .QN( u2_uk_n1774 ) );
  DFF_X1 u2_uk_K_r12_reg_7 (.CK( clk ) , .D( u2_uk_K_r11_7 ) , .Q( u2_uk_K_r12_7 ) );
  DFF_X1 u2_uk_K_r12_reg_8 (.CK( clk ) , .D( u2_uk_K_r11_8 ) , .Q( u2_uk_K_r12_8 ) , .QN( u2_uk_n1776 ) );
  DFF_X1 u2_uk_K_r12_reg_9 (.CK( clk ) , .D( u2_uk_K_r11_9 ) , .Q( u2_uk_K_r12_9 ) , .QN( u2_uk_n1777 ) );
  DFF_X1 u2_uk_K_r13_reg_0 (.CK( clk ) , .D( u2_uk_K_r12_0 ) , .Q( u2_uk_K_r13_0 ) , .QN( u2_uk_n1813 ) );
  DFF_X1 u2_uk_K_r13_reg_1 (.CK( clk ) , .D( u2_uk_K_r12_1 ) , .Q( u2_uk_K_r13_1 ) );
  DFF_X1 u2_uk_K_r13_reg_10 (.CK( clk ) , .D( u2_uk_K_r12_10 ) , .Q( u2_uk_K_r13_10 ) , .QN( u2_uk_n1820 ) );
  DFF_X1 u2_uk_K_r13_reg_11 (.CK( clk ) , .D( u2_uk_K_r12_11 ) , .Q( u2_uk_K_r13_11 ) , .QN( u2_uk_n1821 ) );
  DFF_X1 u2_uk_K_r13_reg_12 (.CK( clk ) , .D( u2_uk_K_r12_12 ) , .Q( u2_uk_K_r13_12 ) , .QN( u2_uk_n1822 ) );
  DFF_X1 u2_uk_K_r13_reg_13 (.CK( clk ) , .D( u2_uk_K_r12_13 ) , .Q( u2_uk_K_r13_13 ) , .QN( u2_uk_n1823 ) );
  DFF_X1 u2_uk_K_r13_reg_14 (.CK( clk ) , .D( u2_uk_K_r12_14 ) , .Q( u2_uk_K_r13_14 ) , .QN( u2_uk_n1824 ) );
  DFF_X1 u2_uk_K_r13_reg_15 (.CK( clk ) , .D( u2_uk_K_r12_15 ) , .Q( u2_uk_K_r13_15 ) , .QN( u2_uk_n1825 ) );
  DFF_X1 u2_uk_K_r13_reg_16 (.CK( clk ) , .D( u2_uk_K_r12_16 ) , .Q( u2_uk_K_r13_16 ) , .QN( u2_uk_n1826 ) );
  DFF_X1 u2_uk_K_r13_reg_17 (.CK( clk ) , .D( u2_uk_K_r12_17 ) , .Q( u2_uk_K_r13_17 ) );
  DFF_X1 u2_uk_K_r13_reg_18 (.CK( clk ) , .D( u2_uk_K_r12_18 ) , .Q( u2_uk_K_r13_18 ) , .QN( u2_uk_n1828 ) );
  DFF_X1 u2_uk_K_r13_reg_19 (.CK( clk ) , .D( u2_uk_K_r12_19 ) , .Q( u2_uk_K_r13_19 ) );
  DFF_X1 u2_uk_K_r13_reg_2 (.CK( clk ) , .D( u2_uk_K_r12_2 ) , .Q( u2_uk_K_r13_2 ) );
  DFF_X1 u2_uk_K_r13_reg_20 (.CK( clk ) , .D( u2_uk_K_r12_20 ) , .Q( u2_uk_K_r13_20 ) , .QN( u2_uk_n1829 ) );
  DFF_X1 u2_uk_K_r13_reg_21 (.CK( clk ) , .D( u2_uk_K_r12_21 ) , .Q( u2_uk_K_r13_21 ) , .QN( u2_uk_n1830 ) );
  DFF_X1 u2_uk_K_r13_reg_22 (.CK( clk ) , .D( u2_uk_K_r12_22 ) , .Q( u2_uk_K_r13_22 ) );
  DFF_X1 u2_uk_K_r13_reg_23 (.CK( clk ) , .D( u2_uk_K_r12_23 ) , .Q( u2_uk_K_r13_23 ) );
  DFF_X1 u2_uk_K_r13_reg_24 (.CK( clk ) , .D( u2_uk_K_r12_24 ) , .Q( u2_uk_K_r13_24 ) , .QN( u2_uk_n1832 ) );
  DFF_X1 u2_uk_K_r13_reg_25 (.CK( clk ) , .D( u2_uk_K_r12_25 ) , .Q( u2_uk_K_r13_25 ) );
  DFF_X1 u2_uk_K_r13_reg_26 (.CK( clk ) , .D( u2_uk_K_r12_26 ) , .Q( u2_uk_K_r13_26 ) , .QN( u2_uk_n1833 ) );
  DFF_X1 u2_uk_K_r13_reg_27 (.CK( clk ) , .D( u2_uk_K_r12_27 ) , .Q( u2_uk_K_r13_27 ) , .QN( u2_uk_n1834 ) );
  DFF_X1 u2_uk_K_r13_reg_28 (.CK( clk ) , .D( u2_uk_K_r12_28 ) , .Q( u2_uk_K_r13_28 ) , .QN( u2_uk_n1835 ) );
  DFF_X1 u2_uk_K_r13_reg_29 (.CK( clk ) , .D( u2_uk_K_r12_29 ) , .Q( u2_uk_K_r13_29 ) , .QN( u2_uk_n1836 ) );
  DFF_X1 u2_uk_K_r13_reg_3 (.CK( clk ) , .D( u2_uk_K_r12_3 ) , .Q( u2_uk_K_r13_3 ) , .QN( u2_uk_n1814 ) );
  DFF_X1 u2_uk_K_r13_reg_30 (.CK( clk ) , .D( u2_uk_K_r12_30 ) , .Q( u2_uk_K_r13_30 ) , .QN( u2_uk_n1837 ) );
  DFF_X1 u2_uk_K_r13_reg_31 (.CK( clk ) , .D( u2_uk_K_r12_31 ) , .Q( u2_uk_K_r13_31 ) );
  DFF_X1 u2_uk_K_r13_reg_32 (.CK( clk ) , .D( u2_uk_K_r12_32 ) , .Q( u2_uk_K_r13_32 ) );
  DFF_X1 u2_uk_K_r13_reg_33 (.CK( clk ) , .D( u2_uk_K_r12_33 ) , .Q( u2_uk_K_r13_33 ) , .QN( u2_uk_n1838 ) );
  DFF_X1 u2_uk_K_r13_reg_34 (.CK( clk ) , .D( u2_uk_K_r12_34 ) , .Q( u2_uk_K_r13_34 ) , .QN( u2_uk_n1839 ) );
  DFF_X1 u2_uk_K_r13_reg_35 (.CK( clk ) , .D( u2_uk_K_r12_35 ) , .Q( u2_uk_K_r13_35 ) );
  DFF_X1 u2_uk_K_r13_reg_36 (.CK( clk ) , .D( u2_uk_K_r12_36 ) , .Q( u2_uk_K_r13_36 ) );
  DFF_X1 u2_uk_K_r13_reg_37 (.CK( clk ) , .D( u2_uk_K_r12_37 ) , .Q( u2_uk_K_r13_37 ) , .QN( u2_uk_n1840 ) );
  DFF_X1 u2_uk_K_r13_reg_38 (.CK( clk ) , .D( u2_uk_K_r12_38 ) , .Q( u2_uk_K_r13_38 ) );
  DFF_X1 u2_uk_K_r13_reg_39 (.CK( clk ) , .D( u2_uk_K_r12_39 ) , .Q( u2_uk_K_r13_39 ) , .QN( u2_uk_n1842 ) );
  DFF_X1 u2_uk_K_r13_reg_4 (.CK( clk ) , .D( u2_uk_K_r12_4 ) , .Q( u2_uk_K_r13_4 ) );
  DFF_X1 u2_uk_K_r13_reg_40 (.CK( clk ) , .D( u2_uk_K_r12_40 ) , .Q( u2_uk_K_r13_40 ) , .QN( u2_uk_n1843 ) );
  DFF_X1 u2_uk_K_r13_reg_41 (.CK( clk ) , .D( u2_uk_K_r12_41 ) , .Q( u2_uk_K_r13_41 ) , .QN( u2_uk_n1844 ) );
  DFF_X1 u2_uk_K_r13_reg_42 (.CK( clk ) , .D( u2_uk_K_r12_42 ) , .Q( u2_uk_K_r13_42 ) , .QN( u2_uk_n1845 ) );
  DFF_X1 u2_uk_K_r13_reg_43 (.CK( clk ) , .D( u2_uk_K_r12_43 ) , .Q( u2_uk_K_r13_43 ) , .QN( u2_uk_n1846 ) );
  DFF_X1 u2_uk_K_r13_reg_44 (.CK( clk ) , .D( u2_uk_K_r12_44 ) , .Q( u2_uk_K_r13_44 ) );
  DFF_X1 u2_uk_K_r13_reg_45 (.CK( clk ) , .D( u2_uk_K_r12_45 ) , .Q( u2_uk_K_r13_45 ) , .QN( u2_uk_n1849 ) );
  DFF_X1 u2_uk_K_r13_reg_46 (.CK( clk ) , .D( u2_uk_K_r12_46 ) , .Q( u2_uk_K_r13_46 ) , .QN( u2_uk_n1850 ) );
  DFF_X1 u2_uk_K_r13_reg_47 (.CK( clk ) , .D( u2_uk_K_r12_47 ) , .Q( u2_uk_K_r13_47 ) , .QN( u2_uk_n1851 ) );
  DFF_X1 u2_uk_K_r13_reg_48 (.CK( clk ) , .D( u2_uk_K_r12_48 ) , .Q( u2_uk_K_r13_48 ) , .QN( u2_uk_n1852 ) );
  DFF_X1 u2_uk_K_r13_reg_49 (.CK( clk ) , .D( u2_uk_K_r12_49 ) , .Q( u2_uk_K_r13_49 ) , .QN( u2_uk_n1853 ) );
  DFF_X1 u2_uk_K_r13_reg_5 (.CK( clk ) , .D( u2_uk_K_r12_5 ) , .Q( u2_uk_K_r13_5 ) , .QN( u2_uk_n1815 ) );
  DFF_X1 u2_uk_K_r13_reg_50 (.CK( clk ) , .D( u2_uk_K_r12_50 ) , .Q( u2_uk_K_r13_50 ) , .QN( u2_uk_n1854 ) );
  DFF_X1 u2_uk_K_r13_reg_51 (.CK( clk ) , .D( u2_uk_K_r12_51 ) , .Q( u2_uk_K_r13_51 ) , .QN( u2_uk_n1855 ) );
  DFF_X1 u2_uk_K_r13_reg_52 (.CK( clk ) , .D( u2_uk_K_r12_52 ) , .Q( u2_uk_K_r13_52 ) , .QN( u2_uk_n1856 ) );
  DFF_X1 u2_uk_K_r13_reg_53 (.CK( clk ) , .D( u2_uk_K_r12_53 ) , .Q( u2_uk_K_r13_53 ) );
  DFF_X1 u2_uk_K_r13_reg_54 (.CK( clk ) , .D( u2_uk_K_r12_54 ) , .Q( u2_uk_K_r13_54 ) , .QN( u2_uk_n1857 ) );
  DFF_X1 u2_uk_K_r13_reg_55 (.CK( clk ) , .D( u2_uk_K_r12_55 ) , .Q( u2_uk_K_r13_55 ) );
  DFF_X1 u2_uk_K_r13_reg_6 (.CK( clk ) , .D( u2_uk_K_r12_6 ) , .Q( u2_uk_K_r13_6 ) , .QN( u2_uk_n1816 ) );
  DFF_X1 u2_uk_K_r13_reg_7 (.CK( clk ) , .D( u2_uk_K_r12_7 ) , .Q( u2_uk_K_r13_7 ) , .QN( u2_uk_n1817 ) );
  DFF_X1 u2_uk_K_r13_reg_8 (.CK( clk ) , .D( u2_uk_K_r12_8 ) , .Q( u2_uk_K_r13_8 ) , .QN( u2_uk_n1818 ) );
  DFF_X1 u2_uk_K_r13_reg_9 (.CK( clk ) , .D( u2_uk_K_r12_9 ) , .Q( u2_uk_K_r13_9 ) , .QN( u2_uk_n1819 ) );
  DFF_X1 u2_uk_K_r14_reg_0 (.CK( clk ) , .D( u2_uk_K_r13_0 ) , .QN( u2_uk_n1188 ) );
  DFF_X1 u2_uk_K_r14_reg_1 (.CK( clk ) , .D( u2_uk_K_r13_1 ) , .QN( u2_uk_n1189 ) );
  DFF_X1 u2_uk_K_r14_reg_10 (.CK( clk ) , .D( u2_uk_K_r13_10 ) , .Q( u2_uk_K_r14_10 ) );
  DFF_X1 u2_uk_K_r14_reg_11 (.CK( clk ) , .D( u2_uk_K_r13_11 ) , .Q( u2_uk_K_r14_11 ) );
  DFF_X1 u2_uk_K_r14_reg_12 (.CK( clk ) , .D( u2_uk_K_r13_12 ) , .Q( u2_uk_K_r14_12 ) );
  DFF_X1 u2_uk_K_r14_reg_13 (.CK( clk ) , .D( u2_uk_K_r13_13 ) , .QN( u2_uk_n1194 ) );
  DFF_X1 u2_uk_K_r14_reg_14 (.CK( clk ) , .D( u2_uk_K_r13_14 ) , .QN( u2_uk_n1195 ) );
  DFF_X1 u2_uk_K_r14_reg_15 (.CK( clk ) , .D( u2_uk_K_r13_15 ) , .Q( u2_uk_K_r14_15 ) );
  DFF_X1 u2_uk_K_r14_reg_16 (.CK( clk ) , .D( u2_uk_K_r13_16 ) , .Q( u2_uk_K_r14_16 ) );
  DFF_X1 u2_uk_K_r14_reg_17 (.CK( clk ) , .D( u2_uk_K_r13_17 ) , .QN( u2_uk_n1197 ) );
  DFF_X1 u2_uk_K_r14_reg_18 (.CK( clk ) , .D( u2_uk_K_r13_18 ) , .Q( u2_uk_K_r14_18 ) );
  DFF_X1 u2_uk_K_r14_reg_19 (.CK( clk ) , .D( u2_uk_K_r13_19 ) , .QN( u2_uk_n1198 ) );
  DFF_X1 u2_uk_K_r14_reg_2 (.CK( clk ) , .D( u2_uk_K_r13_2 ) , .Q( u2_uk_K_r14_2 ) );
  DFF_X1 u2_uk_K_r14_reg_20 (.CK( clk ) , .D( u2_uk_K_r13_20 ) , .QN( u2_uk_n1199 ) );
  DFF_X1 u2_uk_K_r14_reg_21 (.CK( clk ) , .D( u2_uk_K_r13_21 ) , .QN( u2_uk_n1200 ) );
  DFF_X1 u2_uk_K_r14_reg_22 (.CK( clk ) , .D( u2_uk_K_r13_22 ) , .QN( u2_uk_n1201 ) );
  DFF_X1 u2_uk_K_r14_reg_23 (.CK( clk ) , .D( u2_uk_K_r13_23 ) , .Q( u2_uk_K_r14_23 ) , .QN( u2_uk_n1203 ) );
  DFF_X1 u2_uk_K_r14_reg_24 (.CK( clk ) , .D( u2_uk_K_r13_24 ) , .QN( u2_uk_n1204 ) );
  DFF_X1 u2_uk_K_r14_reg_25 (.CK( clk ) , .D( u2_uk_K_r13_25 ) , .QN( u2_uk_n1205 ) );
  DFF_X1 u2_uk_K_r14_reg_26 (.CK( clk ) , .D( u2_uk_K_r13_26 ) , .QN( u2_uk_n1206 ) );
  DFF_X1 u2_uk_K_r14_reg_27 (.CK( clk ) , .D( u2_uk_K_r13_27 ) , .QN( u2_uk_n1207 ) );
  DFF_X1 u2_uk_K_r14_reg_28 (.CK( clk ) , .D( u2_uk_K_r13_28 ) , .QN( u2_uk_n1208 ) );
  DFF_X1 u2_uk_K_r14_reg_29 (.CK( clk ) , .D( u2_uk_K_r13_29 ) , .QN( u2_uk_n1209 ) );
  DFF_X1 u2_uk_K_r14_reg_3 (.CK( clk ) , .D( u2_uk_K_r13_3 ) , .Q( u2_uk_K_r14_3 ) );
  DFF_X1 u2_uk_K_r14_reg_30 (.CK( clk ) , .D( u2_uk_K_r13_30 ) , .QN( u2_uk_n1210 ) );
  DFF_X1 u2_uk_K_r14_reg_31 (.CK( clk ) , .D( u2_uk_K_r13_31 ) , .QN( u2_uk_n1211 ) );
  DFF_X1 u2_uk_K_r14_reg_32 (.CK( clk ) , .D( u2_uk_K_r13_32 ) , .QN( u2_uk_n1212 ) );
  DFF_X1 u2_uk_K_r14_reg_33 (.CK( clk ) , .D( u2_uk_K_r13_33 ) , .QN( u2_uk_n1213 ) );
  DFF_X1 u2_uk_K_r14_reg_34 (.CK( clk ) , .D( u2_uk_K_r13_34 ) , .QN( u2_uk_n1214 ) );
  DFF_X1 u2_uk_K_r14_reg_35 (.CK( clk ) , .D( u2_uk_K_r13_35 ) , .QN( u2_uk_n1215 ) );
  DFF_X1 u2_uk_K_r14_reg_36 (.CK( clk ) , .D( u2_uk_K_r13_36 ) , .QN( u2_uk_n1216 ) );
  DFF_X1 u2_uk_K_r14_reg_37 (.CK( clk ) , .D( u2_uk_K_r13_37 ) , .QN( u2_uk_n1217 ) );
  DFF_X1 u2_uk_K_r14_reg_38 (.CK( clk ) , .D( u2_uk_K_r13_38 ) , .Q( u2_uk_K_r14_38 ) );
  DFF_X1 u2_uk_K_r14_reg_39 (.CK( clk ) , .D( u2_uk_K_r13_39 ) , .Q( u2_uk_K_r14_39 ) );
  DFF_X1 u2_uk_K_r14_reg_4 (.CK( clk ) , .D( u2_uk_K_r13_4 ) , .QN( u2_uk_n1190 ) );
  DFF_X1 u2_uk_K_r14_reg_40 (.CK( clk ) , .D( u2_uk_K_r13_40 ) , .QN( u2_uk_n1218 ) );
  DFF_X1 u2_uk_K_r14_reg_41 (.CK( clk ) , .D( u2_uk_K_r13_41 ) , .QN( u2_uk_n1219 ) );
  DFF_X1 u2_uk_K_r14_reg_42 (.CK( clk ) , .D( u2_uk_K_r13_42 ) , .Q( u2_uk_K_r14_42 ) );
  DFF_X1 u2_uk_K_r14_reg_43 (.CK( clk ) , .D( u2_uk_K_r13_43 ) , .Q( u2_uk_K_r14_43 ) );
  DFF_X1 u2_uk_K_r14_reg_44 (.CK( clk ) , .D( u2_uk_K_r13_44 ) , .QN( u2_uk_n1220 ) );
  DFF_X1 u2_uk_K_r14_reg_45 (.CK( clk ) , .D( u2_uk_K_r13_45 ) , .Q( u2_uk_K_r14_45 ) );
  DFF_X1 u2_uk_K_r14_reg_46 (.CK( clk ) , .D( u2_uk_K_r13_46 ) , .Q( u2_uk_K_r14_46 ) );
  DFF_X1 u2_uk_K_r14_reg_47 (.CK( clk ) , .D( u2_uk_K_r13_47 ) , .QN( u2_uk_n1221 ) );
  DFF_X1 u2_uk_K_r14_reg_48 (.CK( clk ) , .D( u2_uk_K_r13_48 ) , .QN( u2_uk_n1222 ) );
  DFF_X1 u2_uk_K_r14_reg_49 (.CK( clk ) , .D( u2_uk_K_r13_49 ) , .QN( u2_uk_n1223 ) );
  DFF_X1 u2_uk_K_r14_reg_5 (.CK( clk ) , .D( u2_uk_K_r13_5 ) , .Q( u2_uk_K_r14_5 ) );
  DFF_X1 u2_uk_K_r14_reg_50 (.CK( clk ) , .D( u2_uk_K_r13_50 ) , .Q( u2_uk_K_r14_50 ) );
  DFF_X1 u2_uk_K_r14_reg_51 (.CK( clk ) , .D( u2_uk_K_r13_51 ) , .QN( u2_uk_n1225 ) );
  DFF_X1 u2_uk_K_r14_reg_52 (.CK( clk ) , .D( u2_uk_K_r13_52 ) , .QN( u2_uk_n1226 ) );
  DFF_X1 u2_uk_K_r14_reg_53 (.CK( clk ) , .D( u2_uk_K_r13_53 ) , .QN( u2_uk_n1227 ) );
  DFF_X1 u2_uk_K_r14_reg_54 (.CK( clk ) , .D( u2_uk_K_r13_54 ) , .QN( u2_uk_n1228 ) );
  DFF_X1 u2_uk_K_r14_reg_55 (.CK( clk ) , .D( u2_uk_K_r13_55 ) , .QN( u2_uk_n1229 ) );
  DFF_X1 u2_uk_K_r14_reg_6 (.CK( clk ) , .D( u2_uk_K_r13_6 ) , .QN( u2_uk_n1191 ) );
  DFF_X1 u2_uk_K_r14_reg_7 (.CK( clk ) , .D( u2_uk_K_r13_7 ) , .QN( u2_uk_n1192 ) );
  DFF_X1 u2_uk_K_r14_reg_8 (.CK( clk ) , .D( u2_uk_K_r13_8 ) , .Q( u2_uk_K_r14_8 ) );
  DFF_X1 u2_uk_K_r14_reg_9 (.CK( clk ) , .D( u2_uk_K_r13_9 ) , .Q( u2_uk_K_r14_9 ) );
  DFF_X1 u2_uk_K_r1_reg_0 (.CK( clk ) , .D( u2_uk_K_r0_0 ) , .Q( u2_uk_K_r1_0 ) , .QN( u2_uk_n1277 ) );
  DFF_X1 u2_uk_K_r1_reg_1 (.CK( clk ) , .D( u2_uk_K_r0_1 ) , .Q( u2_uk_K_r1_1 ) , .QN( u2_uk_n1278 ) );
  DFF_X1 u2_uk_K_r1_reg_10 (.CK( clk ) , .D( u2_uk_K_r0_10 ) , .Q( u2_uk_K_r1_10 ) );
  DFF_X1 u2_uk_K_r1_reg_11 (.CK( clk ) , .D( u2_uk_K_r0_11 ) , .Q( u2_uk_K_r1_11 ) , .QN( u2_uk_n1285 ) );
  DFF_X1 u2_uk_K_r1_reg_12 (.CK( clk ) , .D( u2_uk_K_r0_12 ) , .Q( u2_uk_K_r1_12 ) , .QN( u2_uk_n1286 ) );
  DFF_X1 u2_uk_K_r1_reg_13 (.CK( clk ) , .D( u2_uk_K_r0_13 ) , .Q( u2_uk_K_r1_13 ) , .QN( u2_uk_n1287 ) );
  DFF_X1 u2_uk_K_r1_reg_14 (.CK( clk ) , .D( u2_uk_K_r0_14 ) , .Q( u2_uk_K_r1_14 ) , .QN( u2_uk_n1288 ) );
  DFF_X1 u2_uk_K_r1_reg_15 (.CK( clk ) , .D( u2_uk_K_r0_15 ) , .Q( u2_uk_K_r1_15 ) );
  DFF_X1 u2_uk_K_r1_reg_16 (.CK( clk ) , .D( u2_uk_K_r0_16 ) , .Q( u2_uk_K_r1_16 ) );
  DFF_X1 u2_uk_K_r1_reg_17 (.CK( clk ) , .D( u2_uk_K_r0_17 ) , .Q( u2_uk_K_r1_17 ) , .QN( u2_uk_n1289 ) );
  DFF_X1 u2_uk_K_r1_reg_18 (.CK( clk ) , .D( u2_uk_K_r0_18 ) , .Q( u2_uk_K_r1_18 ) );
  DFF_X1 u2_uk_K_r1_reg_19 (.CK( clk ) , .D( u2_uk_K_r0_19 ) , .Q( u2_uk_K_r1_19 ) , .QN( u2_uk_n1290 ) );
  DFF_X1 u2_uk_K_r1_reg_2 (.CK( clk ) , .D( u2_uk_K_r0_2 ) , .Q( u2_uk_K_r1_2 ) , .QN( u2_uk_n1279 ) );
  DFF_X1 u2_uk_K_r1_reg_20 (.CK( clk ) , .D( u2_uk_K_r0_20 ) , .Q( u2_uk_K_r1_20 ) , .QN( u2_uk_n1291 ) );
  DFF_X1 u2_uk_K_r1_reg_21 (.CK( clk ) , .D( u2_uk_K_r0_21 ) , .Q( u2_uk_K_r1_21 ) );
  DFF_X1 u2_uk_K_r1_reg_22 (.CK( clk ) , .D( u2_uk_K_r0_22 ) , .Q( u2_uk_K_r1_22 ) );
  DFF_X1 u2_uk_K_r1_reg_23 (.CK( clk ) , .D( u2_uk_K_r0_23 ) , .Q( u2_uk_K_r1_23 ) , .QN( u2_uk_n1292 ) );
  DFF_X1 u2_uk_K_r1_reg_24 (.CK( clk ) , .D( u2_uk_K_r0_24 ) , .Q( u2_uk_K_r1_24 ) , .QN( u2_uk_n1293 ) );
  DFF_X1 u2_uk_K_r1_reg_25 (.CK( clk ) , .D( u2_uk_K_r0_25 ) , .Q( u2_uk_K_r1_25 ) , .QN( u2_uk_n1294 ) );
  DFF_X1 u2_uk_K_r1_reg_26 (.CK( clk ) , .D( u2_uk_K_r0_26 ) , .Q( u2_uk_K_r1_26 ) , .QN( u2_uk_n1295 ) );
  DFF_X1 u2_uk_K_r1_reg_27 (.CK( clk ) , .D( u2_uk_K_r0_27 ) , .Q( u2_uk_K_r1_27 ) , .QN( u2_uk_n1296 ) );
  DFF_X1 u2_uk_K_r1_reg_28 (.CK( clk ) , .D( u2_uk_K_r0_28 ) , .Q( u2_uk_K_r1_28 ) , .QN( u2_uk_n1297 ) );
  DFF_X1 u2_uk_K_r1_reg_29 (.CK( clk ) , .D( u2_uk_K_r0_29 ) , .Q( u2_uk_K_r1_29 ) , .QN( u2_uk_n1298 ) );
  DFF_X1 u2_uk_K_r1_reg_3 (.CK( clk ) , .D( u2_uk_K_r0_3 ) , .Q( u2_uk_K_r1_3 ) , .QN( u2_uk_n1280 ) );
  DFF_X1 u2_uk_K_r1_reg_30 (.CK( clk ) , .D( u2_uk_K_r0_30 ) , .Q( u2_uk_K_r1_30 ) , .QN( u2_uk_n1299 ) );
  DFF_X1 u2_uk_K_r1_reg_31 (.CK( clk ) , .D( u2_uk_K_r0_31 ) , .Q( u2_uk_K_r1_31 ) , .QN( u2_uk_n1300 ) );
  DFF_X1 u2_uk_K_r1_reg_32 (.CK( clk ) , .D( u2_uk_K_r0_32 ) , .Q( u2_uk_K_r1_32 ) , .QN( u2_uk_n1301 ) );
  DFF_X1 u2_uk_K_r1_reg_33 (.CK( clk ) , .D( u2_uk_K_r0_33 ) , .Q( u2_uk_K_r1_33 ) );
  DFF_X1 u2_uk_K_r1_reg_34 (.CK( clk ) , .D( u2_uk_K_r0_34 ) , .Q( u2_uk_K_r1_34 ) , .QN( u2_uk_n1302 ) );
  DFF_X1 u2_uk_K_r1_reg_35 (.CK( clk ) , .D( u2_uk_K_r0_35 ) , .Q( u2_uk_K_r1_35 ) , .QN( u2_uk_n1303 ) );
  DFF_X1 u2_uk_K_r1_reg_36 (.CK( clk ) , .D( u2_uk_K_r0_36 ) , .Q( u2_uk_K_r1_36 ) );
  DFF_X1 u2_uk_K_r1_reg_37 (.CK( clk ) , .D( u2_uk_K_r0_37 ) , .Q( u2_uk_K_r1_37 ) , .QN( u2_uk_n1304 ) );
  DFF_X1 u2_uk_K_r1_reg_38 (.CK( clk ) , .D( u2_uk_K_r0_38 ) , .Q( u2_uk_K_r1_38 ) , .QN( u2_uk_n1305 ) );
  DFF_X1 u2_uk_K_r1_reg_39 (.CK( clk ) , .D( u2_uk_K_r0_39 ) , .Q( u2_uk_K_r1_39 ) );
  DFF_X1 u2_uk_K_r1_reg_4 (.CK( clk ) , .D( u2_uk_K_r0_4 ) , .Q( u2_uk_K_r1_4 ) , .QN( u2_uk_n1281 ) );
  DFF_X1 u2_uk_K_r1_reg_40 (.CK( clk ) , .D( u2_uk_K_r0_40 ) , .Q( u2_uk_K_r1_40 ) , .QN( u2_uk_n1306 ) );
  DFF_X1 u2_uk_K_r1_reg_41 (.CK( clk ) , .D( u2_uk_K_r0_41 ) , .Q( u2_uk_K_r1_41 ) );
  DFF_X1 u2_uk_K_r1_reg_42 (.CK( clk ) , .D( u2_uk_K_r0_42 ) , .Q( u2_uk_K_r1_42 ) );
  DFF_X1 u2_uk_K_r1_reg_43 (.CK( clk ) , .D( u2_uk_K_r0_43 ) , .Q( u2_uk_K_r1_43 ) , .QN( u2_uk_n1308 ) );
  DFF_X1 u2_uk_K_r1_reg_44 (.CK( clk ) , .D( u2_uk_K_r0_44 ) , .Q( u2_uk_K_r1_44 ) );
  DFF_X1 u2_uk_K_r1_reg_45 (.CK( clk ) , .D( u2_uk_K_r0_45 ) , .Q( u2_uk_K_r1_45 ) , .QN( u2_uk_n1309 ) );
  DFF_X1 u2_uk_K_r1_reg_46 (.CK( clk ) , .D( u2_uk_K_r0_46 ) , .Q( u2_uk_K_r1_46 ) , .QN( u2_uk_n1310 ) );
  DFF_X1 u2_uk_K_r1_reg_47 (.CK( clk ) , .D( u2_uk_K_r0_47 ) , .Q( u2_uk_K_r1_47 ) );
  DFF_X1 u2_uk_K_r1_reg_48 (.CK( clk ) , .D( u2_uk_K_r0_48 ) , .Q( u2_uk_K_r1_48 ) , .QN( u2_uk_n1311 ) );
  DFF_X1 u2_uk_K_r1_reg_49 (.CK( clk ) , .D( u2_uk_K_r0_49 ) , .Q( u2_uk_K_r1_49 ) , .QN( u2_uk_n1312 ) );
  DFF_X1 u2_uk_K_r1_reg_5 (.CK( clk ) , .D( u2_uk_K_r0_5 ) , .Q( u2_uk_K_r1_5 ) , .QN( u2_uk_n1282 ) );
  DFF_X1 u2_uk_K_r1_reg_50 (.CK( clk ) , .D( u2_uk_K_r0_50 ) , .Q( u2_uk_K_r1_50 ) , .QN( u2_uk_n1313 ) );
  DFF_X1 u2_uk_K_r1_reg_51 (.CK( clk ) , .D( u2_uk_K_r0_51 ) , .Q( u2_uk_K_r1_51 ) , .QN( u2_uk_n1314 ) );
  DFF_X1 u2_uk_K_r1_reg_52 (.CK( clk ) , .D( u2_uk_K_r0_52 ) , .Q( u2_uk_K_r1_52 ) , .QN( u2_uk_n1315 ) );
  DFF_X1 u2_uk_K_r1_reg_53 (.CK( clk ) , .D( u2_uk_K_r0_53 ) , .Q( u2_uk_K_r1_53 ) , .QN( u2_uk_n1316 ) );
  DFF_X1 u2_uk_K_r1_reg_54 (.CK( clk ) , .D( u2_uk_K_r0_54 ) , .Q( u2_uk_K_r1_54 ) , .QN( u2_uk_n1317 ) );
  DFF_X1 u2_uk_K_r1_reg_55 (.CK( clk ) , .D( u2_uk_K_r0_55 ) , .Q( u2_uk_K_r1_55 ) , .QN( u2_uk_n1318 ) );
  DFF_X1 u2_uk_K_r1_reg_6 (.CK( clk ) , .D( u2_uk_K_r0_6 ) , .Q( u2_uk_K_r1_6 ) );
  DFF_X1 u2_uk_K_r1_reg_7 (.CK( clk ) , .D( u2_uk_K_r0_7 ) , .Q( u2_uk_K_r1_7 ) );
  DFF_X1 u2_uk_K_r1_reg_8 (.CK( clk ) , .D( u2_uk_K_r0_8 ) , .Q( u2_uk_K_r1_8 ) , .QN( u2_uk_n1283 ) );
  DFF_X1 u2_uk_K_r1_reg_9 (.CK( clk ) , .D( u2_uk_K_r0_9 ) , .Q( u2_uk_K_r1_9 ) , .QN( u2_uk_n1284 ) );
  DFF_X1 u2_uk_K_r2_reg_0 (.CK( clk ) , .D( u2_uk_K_r1_0 ) , .Q( u2_uk_K_r2_0 ) , .QN( u2_uk_n1319 ) );
  DFF_X1 u2_uk_K_r2_reg_1 (.CK( clk ) , .D( u2_uk_K_r1_1 ) , .Q( u2_uk_K_r2_1 ) , .QN( u2_uk_n1320 ) );
  DFF_X1 u2_uk_K_r2_reg_10 (.CK( clk ) , .D( u2_uk_K_r1_10 ) , .Q( u2_uk_K_r2_10 ) , .QN( u2_uk_n1327 ) );
  DFF_X1 u2_uk_K_r2_reg_11 (.CK( clk ) , .D( u2_uk_K_r1_11 ) , .Q( u2_uk_K_r2_11 ) , .QN( u2_uk_n1328 ) );
  DFF_X1 u2_uk_K_r2_reg_12 (.CK( clk ) , .D( u2_uk_K_r1_12 ) , .Q( u2_uk_K_r2_12 ) , .QN( u2_uk_n1329 ) );
  DFF_X1 u2_uk_K_r2_reg_13 (.CK( clk ) , .D( u2_uk_K_r1_13 ) , .Q( u2_uk_K_r2_13 ) );
  DFF_X1 u2_uk_K_r2_reg_14 (.CK( clk ) , .D( u2_uk_K_r1_14 ) , .Q( u2_uk_K_r2_14 ) , .QN( u2_uk_n1330 ) );
  DFF_X1 u2_uk_K_r2_reg_15 (.CK( clk ) , .D( u2_uk_K_r1_15 ) , .Q( u2_uk_K_r2_15 ) , .QN( u2_uk_n1331 ) );
  DFF_X1 u2_uk_K_r2_reg_16 (.CK( clk ) , .D( u2_uk_K_r1_16 ) , .Q( u2_uk_K_r2_16 ) );
  DFF_X1 u2_uk_K_r2_reg_17 (.CK( clk ) , .D( u2_uk_K_r1_17 ) , .Q( u2_uk_K_r2_17 ) , .QN( u2_uk_n1333 ) );
  DFF_X1 u2_uk_K_r2_reg_18 (.CK( clk ) , .D( u2_uk_K_r1_18 ) , .Q( u2_uk_K_r2_18 ) );
  DFF_X1 u2_uk_K_r2_reg_19 (.CK( clk ) , .D( u2_uk_K_r1_19 ) , .Q( u2_uk_K_r2_19 ) , .QN( u2_uk_n1335 ) );
  DFF_X1 u2_uk_K_r2_reg_2 (.CK( clk ) , .D( u2_uk_K_r1_2 ) , .Q( u2_uk_K_r2_2 ) , .QN( u2_uk_n1321 ) );
  DFF_X1 u2_uk_K_r2_reg_20 (.CK( clk ) , .D( u2_uk_K_r1_20 ) , .Q( u2_uk_K_r2_20 ) );
  DFF_X1 u2_uk_K_r2_reg_21 (.CK( clk ) , .D( u2_uk_K_r1_21 ) , .Q( u2_uk_K_r2_21 ) );
  DFF_X1 u2_uk_K_r2_reg_22 (.CK( clk ) , .D( u2_uk_K_r1_22 ) , .Q( u2_uk_K_r2_22 ) , .QN( u2_uk_n1336 ) );
  DFF_X1 u2_uk_K_r2_reg_23 (.CK( clk ) , .D( u2_uk_K_r1_23 ) , .Q( u2_uk_K_r2_23 ) , .QN( u2_uk_n1337 ) );
  DFF_X1 u2_uk_K_r2_reg_24 (.CK( clk ) , .D( u2_uk_K_r1_24 ) , .Q( u2_uk_K_r2_24 ) );
  DFF_X1 u2_uk_K_r2_reg_25 (.CK( clk ) , .D( u2_uk_K_r1_25 ) , .Q( u2_uk_K_r2_25 ) );
  DFF_X1 u2_uk_K_r2_reg_26 (.CK( clk ) , .D( u2_uk_K_r1_26 ) , .Q( u2_uk_K_r2_26 ) );
  DFF_X1 u2_uk_K_r2_reg_27 (.CK( clk ) , .D( u2_uk_K_r1_27 ) , .Q( u2_uk_K_r2_27 ) );
  DFF_X1 u2_uk_K_r2_reg_28 (.CK( clk ) , .D( u2_uk_K_r1_28 ) , .Q( u2_uk_K_r2_28 ) );
  DFF_X1 u2_uk_K_r2_reg_29 (.CK( clk ) , .D( u2_uk_K_r1_29 ) , .Q( u2_uk_K_r2_29 ) );
  DFF_X1 u2_uk_K_r2_reg_3 (.CK( clk ) , .D( u2_uk_K_r1_3 ) , .Q( u2_uk_K_r2_3 ) , .QN( u2_uk_n1322 ) );
  DFF_X1 u2_uk_K_r2_reg_30 (.CK( clk ) , .D( u2_uk_K_r1_30 ) , .Q( u2_uk_K_r2_30 ) );
  DFF_X1 u2_uk_K_r2_reg_31 (.CK( clk ) , .D( u2_uk_K_r1_31 ) , .Q( u2_uk_K_r2_31 ) );
  DFF_X1 u2_uk_K_r2_reg_32 (.CK( clk ) , .D( u2_uk_K_r1_32 ) , .Q( u2_uk_K_r2_32 ) , .QN( u2_uk_n1339 ) );
  DFF_X1 u2_uk_K_r2_reg_33 (.CK( clk ) , .D( u2_uk_K_r1_33 ) , .Q( u2_uk_K_r2_33 ) );
  DFF_X1 u2_uk_K_r2_reg_34 (.CK( clk ) , .D( u2_uk_K_r1_34 ) , .Q( u2_uk_K_r2_34 ) , .QN( u2_uk_n1341 ) );
  DFF_X1 u2_uk_K_r2_reg_35 (.CK( clk ) , .D( u2_uk_K_r1_35 ) , .Q( u2_uk_K_r2_35 ) , .QN( u2_uk_n1342 ) );
  DFF_X1 u2_uk_K_r2_reg_36 (.CK( clk ) , .D( u2_uk_K_r1_36 ) , .Q( u2_uk_K_r2_36 ) , .QN( u2_uk_n1344 ) );
  DFF_X1 u2_uk_K_r2_reg_37 (.CK( clk ) , .D( u2_uk_K_r1_37 ) , .Q( u2_uk_K_r2_37 ) , .QN( u2_uk_n1345 ) );
  DFF_X1 u2_uk_K_r2_reg_38 (.CK( clk ) , .D( u2_uk_K_r1_38 ) , .Q( u2_uk_K_r2_38 ) , .QN( u2_uk_n1346 ) );
  DFF_X1 u2_uk_K_r2_reg_39 (.CK( clk ) , .D( u2_uk_K_r1_39 ) , .Q( u2_uk_K_r2_39 ) , .QN( u2_uk_n1347 ) );
  DFF_X1 u2_uk_K_r2_reg_4 (.CK( clk ) , .D( u2_uk_K_r1_4 ) , .Q( u2_uk_K_r2_4 ) );
  DFF_X1 u2_uk_K_r2_reg_40 (.CK( clk ) , .D( u2_uk_K_r1_40 ) , .Q( u2_uk_K_r2_40 ) , .QN( u2_uk_n1348 ) );
  DFF_X1 u2_uk_K_r2_reg_41 (.CK( clk ) , .D( u2_uk_K_r1_41 ) , .Q( u2_uk_K_r2_41 ) );
  DFF_X1 u2_uk_K_r2_reg_42 (.CK( clk ) , .D( u2_uk_K_r1_42 ) , .Q( u2_uk_K_r2_42 ) , .QN( u2_uk_n1350 ) );
  DFF_X1 u2_uk_K_r2_reg_43 (.CK( clk ) , .D( u2_uk_K_r1_43 ) , .Q( u2_uk_K_r2_43 ) , .QN( u2_uk_n1351 ) );
  DFF_X1 u2_uk_K_r2_reg_44 (.CK( clk ) , .D( u2_uk_K_r1_44 ) , .Q( u2_uk_K_r2_44 ) , .QN( u2_uk_n1352 ) );
  DFF_X1 u2_uk_K_r2_reg_45 (.CK( clk ) , .D( u2_uk_K_r1_45 ) , .Q( u2_uk_K_r2_45 ) , .QN( u2_uk_n1353 ) );
  DFF_X1 u2_uk_K_r2_reg_46 (.CK( clk ) , .D( u2_uk_K_r1_46 ) , .Q( u2_uk_K_r2_46 ) );
  DFF_X1 u2_uk_K_r2_reg_47 (.CK( clk ) , .D( u2_uk_K_r1_47 ) , .Q( u2_uk_K_r2_47 ) );
  DFF_X1 u2_uk_K_r2_reg_48 (.CK( clk ) , .D( u2_uk_K_r1_48 ) , .Q( u2_uk_K_r2_48 ) , .QN( u2_uk_n1356 ) );
  DFF_X1 u2_uk_K_r2_reg_49 (.CK( clk ) , .D( u2_uk_K_r1_49 ) , .Q( u2_uk_K_r2_49 ) );
  DFF_X1 u2_uk_K_r2_reg_5 (.CK( clk ) , .D( u2_uk_K_r1_5 ) , .Q( u2_uk_K_r2_5 ) , .QN( u2_uk_n1323 ) );
  DFF_X1 u2_uk_K_r2_reg_50 (.CK( clk ) , .D( u2_uk_K_r1_50 ) , .Q( u2_uk_K_r2_50 ) );
  DFF_X1 u2_uk_K_r2_reg_51 (.CK( clk ) , .D( u2_uk_K_r1_51 ) , .Q( u2_uk_K_r2_51 ) , .QN( u2_uk_n1359 ) );
  DFF_X1 u2_uk_K_r2_reg_52 (.CK( clk ) , .D( u2_uk_K_r1_52 ) , .Q( u2_uk_K_r2_52 ) , .QN( u2_uk_n1360 ) );
  DFF_X1 u2_uk_K_r2_reg_53 (.CK( clk ) , .D( u2_uk_K_r1_53 ) , .Q( u2_uk_K_r2_53 ) );
  DFF_X1 u2_uk_K_r2_reg_54 (.CK( clk ) , .D( u2_uk_K_r1_54 ) , .Q( u2_uk_K_r2_54 ) , .QN( u2_uk_n1361 ) );
  DFF_X1 u2_uk_K_r2_reg_55 (.CK( clk ) , .D( u2_uk_K_r1_55 ) , .Q( u2_uk_K_r2_55 ) , .QN( u2_uk_n1363 ) );
  DFF_X1 u2_uk_K_r2_reg_6 (.CK( clk ) , .D( u2_uk_K_r1_6 ) , .Q( u2_uk_K_r2_6 ) , .QN( u2_uk_n1324 ) );
  DFF_X1 u2_uk_K_r2_reg_7 (.CK( clk ) , .D( u2_uk_K_r1_7 ) , .Q( u2_uk_K_r2_7 ) );
  DFF_X1 u2_uk_K_r2_reg_8 (.CK( clk ) , .D( u2_uk_K_r1_8 ) , .Q( u2_uk_K_r2_8 ) , .QN( u2_uk_n1325 ) );
  DFF_X1 u2_uk_K_r2_reg_9 (.CK( clk ) , .D( u2_uk_K_r1_9 ) , .Q( u2_uk_K_r2_9 ) , .QN( u2_uk_n1326 ) );
  DFF_X1 u2_uk_K_r3_reg_0 (.CK( clk ) , .D( u2_uk_K_r2_0 ) , .Q( u2_uk_K_r3_0 ) , .QN( u2_uk_n1364 ) );
  DFF_X1 u2_uk_K_r3_reg_1 (.CK( clk ) , .D( u2_uk_K_r2_1 ) , .Q( u2_uk_K_r3_1 ) , .QN( u2_uk_n1365 ) );
  DFF_X1 u2_uk_K_r3_reg_10 (.CK( clk ) , .D( u2_uk_K_r2_10 ) , .Q( u2_uk_K_r3_10 ) );
  DFF_X1 u2_uk_K_r3_reg_11 (.CK( clk ) , .D( u2_uk_K_r2_11 ) , .Q( u2_uk_K_r3_11 ) );
  DFF_X1 u2_uk_K_r3_reg_12 (.CK( clk ) , .D( u2_uk_K_r2_12 ) , .Q( u2_uk_K_r3_12 ) , .QN( u2_uk_n1372 ) );
  DFF_X1 u2_uk_K_r3_reg_13 (.CK( clk ) , .D( u2_uk_K_r2_13 ) , .Q( u2_uk_K_r3_13 ) );
  DFF_X1 u2_uk_K_r3_reg_14 (.CK( clk ) , .D( u2_uk_K_r2_14 ) , .Q( u2_uk_K_r3_14 ) );
  DFF_X1 u2_uk_K_r3_reg_15 (.CK( clk ) , .D( u2_uk_K_r2_15 ) , .Q( u2_uk_K_r3_15 ) );
  DFF_X1 u2_uk_K_r3_reg_16 (.CK( clk ) , .D( u2_uk_K_r2_16 ) , .Q( u2_uk_K_r3_16 ) );
  DFF_X1 u2_uk_K_r3_reg_17 (.CK( clk ) , .D( u2_uk_K_r2_17 ) , .Q( u2_uk_K_r3_17 ) , .QN( u2_uk_n1373 ) );
  DFF_X1 u2_uk_K_r3_reg_18 (.CK( clk ) , .D( u2_uk_K_r2_18 ) , .Q( u2_uk_K_r3_18 ) , .QN( u2_uk_n1374 ) );
  DFF_X1 u2_uk_K_r3_reg_19 (.CK( clk ) , .D( u2_uk_K_r2_19 ) , .Q( u2_uk_K_r3_19 ) );
  DFF_X1 u2_uk_K_r3_reg_2 (.CK( clk ) , .D( u2_uk_K_r2_2 ) , .Q( u2_uk_K_r3_2 ) , .QN( u2_uk_n1366 ) );
  DFF_X1 u2_uk_K_r3_reg_20 (.CK( clk ) , .D( u2_uk_K_r2_20 ) , .Q( u2_uk_K_r3_20 ) , .QN( u2_uk_n1375 ) );
  DFF_X1 u2_uk_K_r3_reg_21 (.CK( clk ) , .D( u2_uk_K_r2_21 ) , .Q( u2_uk_K_r3_21 ) , .QN( u2_uk_n1376 ) );
  DFF_X1 u2_uk_K_r3_reg_22 (.CK( clk ) , .D( u2_uk_K_r2_22 ) , .Q( u2_uk_K_r3_22 ) , .QN( u2_uk_n1377 ) );
  DFF_X1 u2_uk_K_r3_reg_23 (.CK( clk ) , .D( u2_uk_K_r2_23 ) , .Q( u2_uk_K_r3_23 ) , .QN( u2_uk_n1378 ) );
  DFF_X1 u2_uk_K_r3_reg_24 (.CK( clk ) , .D( u2_uk_K_r2_24 ) , .Q( u2_uk_K_r3_24 ) );
  DFF_X1 u2_uk_K_r3_reg_25 (.CK( clk ) , .D( u2_uk_K_r2_25 ) , .Q( u2_uk_K_r3_25 ) , .QN( u2_uk_n1379 ) );
  DFF_X1 u2_uk_K_r3_reg_26 (.CK( clk ) , .D( u2_uk_K_r2_26 ) , .Q( u2_uk_K_r3_26 ) , .QN( u2_uk_n1380 ) );
  DFF_X1 u2_uk_K_r3_reg_27 (.CK( clk ) , .D( u2_uk_K_r2_27 ) , .Q( u2_uk_K_r3_27 ) , .QN( u2_uk_n1381 ) );
  DFF_X1 u2_uk_K_r3_reg_28 (.CK( clk ) , .D( u2_uk_K_r2_28 ) , .Q( u2_uk_K_r3_28 ) , .QN( u2_uk_n1382 ) );
  DFF_X1 u2_uk_K_r3_reg_29 (.CK( clk ) , .D( u2_uk_K_r2_29 ) , .Q( u2_uk_K_r3_29 ) );
  DFF_X1 u2_uk_K_r3_reg_3 (.CK( clk ) , .D( u2_uk_K_r2_3 ) , .Q( u2_uk_K_r3_3 ) , .QN( u2_uk_n1367 ) );
  DFF_X1 u2_uk_K_r3_reg_30 (.CK( clk ) , .D( u2_uk_K_r2_30 ) , .Q( u2_uk_K_r3_30 ) , .QN( u2_uk_n1383 ) );
  DFF_X1 u2_uk_K_r3_reg_31 (.CK( clk ) , .D( u2_uk_K_r2_31 ) , .Q( u2_uk_K_r3_31 ) , .QN( u2_uk_n1384 ) );
  DFF_X1 u2_uk_K_r3_reg_32 (.CK( clk ) , .D( u2_uk_K_r2_32 ) , .Q( u2_uk_K_r3_32 ) , .QN( u2_uk_n1385 ) );
  DFF_X1 u2_uk_K_r3_reg_33 (.CK( clk ) , .D( u2_uk_K_r2_33 ) , .Q( u2_uk_K_r3_33 ) , .QN( u2_uk_n1387 ) );
  DFF_X1 u2_uk_K_r3_reg_34 (.CK( clk ) , .D( u2_uk_K_r2_34 ) , .Q( u2_uk_K_r3_34 ) );
  DFF_X1 u2_uk_K_r3_reg_35 (.CK( clk ) , .D( u2_uk_K_r2_35 ) , .Q( u2_uk_K_r3_35 ) );
  DFF_X1 u2_uk_K_r3_reg_36 (.CK( clk ) , .D( u2_uk_K_r2_36 ) , .Q( u2_uk_K_r3_36 ) , .QN( u2_uk_n1388 ) );
  DFF_X1 u2_uk_K_r3_reg_37 (.CK( clk ) , .D( u2_uk_K_r2_37 ) , .Q( u2_uk_K_r3_37 ) , .QN( u2_uk_n1389 ) );
  DFF_X1 u2_uk_K_r3_reg_38 (.CK( clk ) , .D( u2_uk_K_r2_38 ) , .Q( u2_uk_K_r3_38 ) );
  DFF_X1 u2_uk_K_r3_reg_39 (.CK( clk ) , .D( u2_uk_K_r2_39 ) , .Q( u2_uk_K_r3_39 ) , .QN( u2_uk_n1392 ) );
  DFF_X1 u2_uk_K_r3_reg_4 (.CK( clk ) , .D( u2_uk_K_r2_4 ) , .Q( u2_uk_K_r3_4 ) );
  DFF_X1 u2_uk_K_r3_reg_40 (.CK( clk ) , .D( u2_uk_K_r2_40 ) , .Q( u2_uk_K_r3_40 ) , .QN( u2_uk_n1393 ) );
  DFF_X1 u2_uk_K_r3_reg_41 (.CK( clk ) , .D( u2_uk_K_r2_41 ) , .Q( u2_uk_K_r3_41 ) , .QN( u2_uk_n1394 ) );
  DFF_X1 u2_uk_K_r3_reg_42 (.CK( clk ) , .D( u2_uk_K_r2_42 ) , .Q( u2_uk_K_r3_42 ) , .QN( u2_uk_n1395 ) );
  DFF_X1 u2_uk_K_r3_reg_43 (.CK( clk ) , .D( u2_uk_K_r2_43 ) , .Q( u2_uk_K_r3_43 ) );
  DFF_X1 u2_uk_K_r3_reg_44 (.CK( clk ) , .D( u2_uk_K_r2_44 ) , .Q( u2_uk_K_r3_44 ) );
  DFF_X1 u2_uk_K_r3_reg_45 (.CK( clk ) , .D( u2_uk_K_r2_45 ) , .Q( u2_uk_K_r3_45 ) , .QN( u2_uk_n1396 ) );
  DFF_X1 u2_uk_K_r3_reg_46 (.CK( clk ) , .D( u2_uk_K_r2_46 ) , .Q( u2_uk_K_r3_46 ) , .QN( u2_uk_n1397 ) );
  DFF_X1 u2_uk_K_r3_reg_47 (.CK( clk ) , .D( u2_uk_K_r2_47 ) , .Q( u2_uk_K_r3_47 ) );
  DFF_X1 u2_uk_K_r3_reg_48 (.CK( clk ) , .D( u2_uk_K_r2_48 ) , .Q( u2_uk_K_r3_48 ) , .QN( u2_uk_n1399 ) );
  DFF_X1 u2_uk_K_r3_reg_49 (.CK( clk ) , .D( u2_uk_K_r2_49 ) , .Q( u2_uk_K_r3_49 ) , .QN( u2_uk_n1400 ) );
  DFF_X1 u2_uk_K_r3_reg_5 (.CK( clk ) , .D( u2_uk_K_r2_5 ) , .Q( u2_uk_K_r3_5 ) , .QN( u2_uk_n1368 ) );
  DFF_X1 u2_uk_K_r3_reg_50 (.CK( clk ) , .D( u2_uk_K_r2_50 ) , .Q( u2_uk_K_r3_50 ) , .QN( u2_uk_n1401 ) );
  DFF_X1 u2_uk_K_r3_reg_51 (.CK( clk ) , .D( u2_uk_K_r2_51 ) , .Q( u2_uk_K_r3_51 ) , .QN( u2_uk_n1403 ) );
  DFF_X1 u2_uk_K_r3_reg_52 (.CK( clk ) , .D( u2_uk_K_r2_52 ) , .Q( u2_uk_K_r3_52 ) );
  DFF_X1 u2_uk_K_r3_reg_53 (.CK( clk ) , .D( u2_uk_K_r2_53 ) , .Q( u2_uk_K_r3_53 ) , .QN( u2_uk_n1405 ) );
  DFF_X1 u2_uk_K_r3_reg_54 (.CK( clk ) , .D( u2_uk_K_r2_54 ) , .Q( u2_uk_K_r3_54 ) , .QN( u2_uk_n1406 ) );
  DFF_X1 u2_uk_K_r3_reg_55 (.CK( clk ) , .D( u2_uk_K_r2_55 ) , .Q( u2_uk_K_r3_55 ) , .QN( u2_uk_n1407 ) );
  DFF_X1 u2_uk_K_r3_reg_6 (.CK( clk ) , .D( u2_uk_K_r2_6 ) , .Q( u2_uk_K_r3_6 ) , .QN( u2_uk_n1369 ) );
  DFF_X1 u2_uk_K_r3_reg_7 (.CK( clk ) , .D( u2_uk_K_r2_7 ) , .Q( u2_uk_K_r3_7 ) , .QN( u2_uk_n1370 ) );
  DFF_X1 u2_uk_K_r3_reg_8 (.CK( clk ) , .D( u2_uk_K_r2_8 ) , .Q( u2_uk_K_r3_8 ) , .QN( u2_uk_n1371 ) );
  DFF_X1 u2_uk_K_r3_reg_9 (.CK( clk ) , .D( u2_uk_K_r2_9 ) , .Q( u2_uk_K_r3_9 ) );
  DFF_X1 u2_uk_K_r4_reg_0 (.CK( clk ) , .D( u2_uk_K_r3_0 ) , .Q( u2_uk_K_r4_0 ) );
  DFF_X1 u2_uk_K_r4_reg_1 (.CK( clk ) , .D( u2_uk_K_r3_1 ) , .Q( u2_uk_K_r4_1 ) , .QN( u2_uk_n1408 ) );
  DFF_X1 u2_uk_K_r4_reg_10 (.CK( clk ) , .D( u2_uk_K_r3_10 ) , .Q( u2_uk_K_r4_10 ) , .QN( u2_uk_n1414 ) );
  DFF_X1 u2_uk_K_r4_reg_11 (.CK( clk ) , .D( u2_uk_K_r3_11 ) , .Q( u2_uk_K_r4_11 ) );
  DFF_X1 u2_uk_K_r4_reg_12 (.CK( clk ) , .D( u2_uk_K_r3_12 ) , .Q( u2_uk_K_r4_12 ) , .QN( u2_uk_n1416 ) );
  DFF_X1 u2_uk_K_r4_reg_13 (.CK( clk ) , .D( u2_uk_K_r3_13 ) , .Q( u2_uk_K_r4_13 ) , .QN( u2_uk_n1417 ) );
  DFF_X1 u2_uk_K_r4_reg_14 (.CK( clk ) , .D( u2_uk_K_r3_14 ) , .Q( u2_uk_K_r4_14 ) , .QN( u2_uk_n1418 ) );
  DFF_X1 u2_uk_K_r4_reg_15 (.CK( clk ) , .D( u2_uk_K_r3_15 ) , .Q( u2_uk_K_r4_15 ) , .QN( u2_uk_n1419 ) );
  DFF_X1 u2_uk_K_r4_reg_16 (.CK( clk ) , .D( u2_uk_K_r3_16 ) , .Q( u2_uk_K_r4_16 ) , .QN( u2_uk_n1420 ) );
  DFF_X1 u2_uk_K_r4_reg_17 (.CK( clk ) , .D( u2_uk_K_r3_17 ) , .Q( u2_uk_K_r4_17 ) );
  DFF_X1 u2_uk_K_r4_reg_18 (.CK( clk ) , .D( u2_uk_K_r3_18 ) , .Q( u2_uk_K_r4_18 ) );
  DFF_X1 u2_uk_K_r4_reg_19 (.CK( clk ) , .D( u2_uk_K_r3_19 ) , .Q( u2_uk_K_r4_19 ) , .QN( u2_uk_n1422 ) );
  DFF_X1 u2_uk_K_r4_reg_2 (.CK( clk ) , .D( u2_uk_K_r3_2 ) , .Q( u2_uk_K_r4_2 ) );
  DFF_X1 u2_uk_K_r4_reg_20 (.CK( clk ) , .D( u2_uk_K_r3_20 ) , .Q( u2_uk_K_r4_20 ) , .QN( u2_uk_n1423 ) );
  DFF_X1 u2_uk_K_r4_reg_21 (.CK( clk ) , .D( u2_uk_K_r3_21 ) , .Q( u2_uk_K_r4_21 ) , .QN( u2_uk_n1424 ) );
  DFF_X1 u2_uk_K_r4_reg_22 (.CK( clk ) , .D( u2_uk_K_r3_22 ) , .Q( u2_uk_K_r4_22 ) , .QN( u2_uk_n1425 ) );
  DFF_X1 u2_uk_K_r4_reg_23 (.CK( clk ) , .D( u2_uk_K_r3_23 ) , .Q( u2_uk_K_r4_23 ) );
  DFF_X1 u2_uk_K_r4_reg_24 (.CK( clk ) , .D( u2_uk_K_r3_24 ) , .Q( u2_uk_K_r4_24 ) );
  DFF_X1 u2_uk_K_r4_reg_25 (.CK( clk ) , .D( u2_uk_K_r3_25 ) , .Q( u2_uk_K_r4_25 ) , .QN( u2_uk_n1426 ) );
  DFF_X1 u2_uk_K_r4_reg_26 (.CK( clk ) , .D( u2_uk_K_r3_26 ) , .Q( u2_uk_K_r4_26 ) , .QN( u2_uk_n1427 ) );
  DFF_X1 u2_uk_K_r4_reg_27 (.CK( clk ) , .D( u2_uk_K_r3_27 ) , .Q( u2_uk_K_r4_27 ) );
  DFF_X1 u2_uk_K_r4_reg_28 (.CK( clk ) , .D( u2_uk_K_r3_28 ) , .Q( u2_uk_K_r4_28 ) , .QN( u2_uk_n1428 ) );
  DFF_X1 u2_uk_K_r4_reg_29 (.CK( clk ) , .D( u2_uk_K_r3_29 ) , .Q( u2_uk_K_r4_29 ) , .QN( u2_uk_n1429 ) );
  DFF_X1 u2_uk_K_r4_reg_3 (.CK( clk ) , .D( u2_uk_K_r3_3 ) , .Q( u2_uk_K_r4_3 ) );
  DFF_X1 u2_uk_K_r4_reg_30 (.CK( clk ) , .D( u2_uk_K_r3_30 ) , .Q( u2_uk_K_r4_30 ) , .QN( u2_uk_n1430 ) );
  DFF_X1 u2_uk_K_r4_reg_31 (.CK( clk ) , .D( u2_uk_K_r3_31 ) , .Q( u2_uk_K_r4_31 ) );
  DFF_X1 u2_uk_K_r4_reg_32 (.CK( clk ) , .D( u2_uk_K_r3_32 ) , .Q( u2_uk_K_r4_32 ) , .QN( u2_uk_n1431 ) );
  DFF_X1 u2_uk_K_r4_reg_33 (.CK( clk ) , .D( u2_uk_K_r3_33 ) , .Q( u2_uk_K_r4_33 ) );
  DFF_X1 u2_uk_K_r4_reg_34 (.CK( clk ) , .D( u2_uk_K_r3_34 ) , .Q( u2_uk_K_r4_34 ) , .QN( u2_uk_n1432 ) );
  DFF_X1 u2_uk_K_r4_reg_35 (.CK( clk ) , .D( u2_uk_K_r3_35 ) , .Q( u2_uk_K_r4_35 ) );
  DFF_X1 u2_uk_K_r4_reg_36 (.CK( clk ) , .D( u2_uk_K_r3_36 ) , .Q( u2_uk_K_r4_36 ) , .QN( u2_uk_n1433 ) );
  DFF_X1 u2_uk_K_r4_reg_37 (.CK( clk ) , .D( u2_uk_K_r3_37 ) , .Q( u2_uk_K_r4_37 ) , .QN( u2_uk_n1434 ) );
  DFF_X1 u2_uk_K_r4_reg_38 (.CK( clk ) , .D( u2_uk_K_r3_38 ) , .Q( u2_uk_K_r4_38 ) );
  DFF_X1 u2_uk_K_r4_reg_39 (.CK( clk ) , .D( u2_uk_K_r3_39 ) , .Q( u2_uk_K_r4_39 ) , .QN( u2_uk_n1435 ) );
  DFF_X1 u2_uk_K_r4_reg_4 (.CK( clk ) , .D( u2_uk_K_r3_4 ) , .Q( u2_uk_K_r4_4 ) , .QN( u2_uk_n1409 ) );
  DFF_X1 u2_uk_K_r4_reg_40 (.CK( clk ) , .D( u2_uk_K_r3_40 ) , .Q( u2_uk_K_r4_40 ) , .QN( u2_uk_n1436 ) );
  DFF_X1 u2_uk_K_r4_reg_41 (.CK( clk ) , .D( u2_uk_K_r3_41 ) , .Q( u2_uk_K_r4_41 ) );
  DFF_X1 u2_uk_K_r4_reg_42 (.CK( clk ) , .D( u2_uk_K_r3_42 ) , .Q( u2_uk_K_r4_42 ) , .QN( u2_uk_n1438 ) );
  DFF_X1 u2_uk_K_r4_reg_43 (.CK( clk ) , .D( u2_uk_K_r3_43 ) , .Q( u2_uk_K_r4_43 ) , .QN( u2_uk_n1439 ) );
  DFF_X1 u2_uk_K_r4_reg_44 (.CK( clk ) , .D( u2_uk_K_r3_44 ) , .Q( u2_uk_K_r4_44 ) , .QN( u2_uk_n1440 ) );
  DFF_X1 u2_uk_K_r4_reg_45 (.CK( clk ) , .D( u2_uk_K_r3_45 ) , .Q( u2_uk_K_r4_45 ) , .QN( u2_uk_n1441 ) );
  DFF_X1 u2_uk_K_r4_reg_46 (.CK( clk ) , .D( u2_uk_K_r3_46 ) , .Q( u2_uk_K_r4_46 ) , .QN( u2_uk_n1442 ) );
  DFF_X1 u2_uk_K_r4_reg_47 (.CK( clk ) , .D( u2_uk_K_r3_47 ) , .Q( u2_uk_K_r4_47 ) , .QN( u2_uk_n1444 ) );
  DFF_X1 u2_uk_K_r4_reg_48 (.CK( clk ) , .D( u2_uk_K_r3_48 ) , .Q( u2_uk_K_r4_48 ) );
  DFF_X1 u2_uk_K_r4_reg_49 (.CK( clk ) , .D( u2_uk_K_r3_49 ) , .Q( u2_uk_K_r4_49 ) );
  DFF_X1 u2_uk_K_r4_reg_5 (.CK( clk ) , .D( u2_uk_K_r3_5 ) , .Q( u2_uk_K_r4_5 ) );
  DFF_X1 u2_uk_K_r4_reg_50 (.CK( clk ) , .D( u2_uk_K_r3_50 ) , .Q( u2_uk_K_r4_50 ) , .QN( u2_uk_n1445 ) );
  DFF_X1 u2_uk_K_r4_reg_51 (.CK( clk ) , .D( u2_uk_K_r3_51 ) , .Q( u2_uk_K_r4_51 ) , .QN( u2_uk_n1446 ) );
  DFF_X1 u2_uk_K_r4_reg_52 (.CK( clk ) , .D( u2_uk_K_r3_52 ) , .Q( u2_uk_K_r4_52 ) , .QN( u2_uk_n1447 ) );
  DFF_X1 u2_uk_K_r4_reg_53 (.CK( clk ) , .D( u2_uk_K_r3_53 ) , .Q( u2_uk_K_r4_53 ) , .QN( u2_uk_n1448 ) );
  DFF_X1 u2_uk_K_r4_reg_54 (.CK( clk ) , .D( u2_uk_K_r3_54 ) , .Q( u2_uk_K_r4_54 ) );
  DFF_X1 u2_uk_K_r4_reg_55 (.CK( clk ) , .D( u2_uk_K_r3_55 ) , .Q( u2_uk_K_r4_55 ) );
  DFF_X1 u2_uk_K_r4_reg_6 (.CK( clk ) , .D( u2_uk_K_r3_6 ) , .Q( u2_uk_K_r4_6 ) , .QN( u2_uk_n1410 ) );
  DFF_X1 u2_uk_K_r4_reg_7 (.CK( clk ) , .D( u2_uk_K_r3_7 ) , .Q( u2_uk_K_r4_7 ) , .QN( u2_uk_n1411 ) );
  DFF_X1 u2_uk_K_r4_reg_8 (.CK( clk ) , .D( u2_uk_K_r3_8 ) , .Q( u2_uk_K_r4_8 ) , .QN( u2_uk_n1412 ) );
  DFF_X1 u2_uk_K_r4_reg_9 (.CK( clk ) , .D( u2_uk_K_r3_9 ) , .Q( u2_uk_K_r4_9 ) , .QN( u2_uk_n1413 ) );
  DFF_X1 u2_uk_K_r5_reg_0 (.CK( clk ) , .D( u2_uk_K_r4_0 ) , .Q( u2_uk_K_r5_0 ) );
  DFF_X1 u2_uk_K_r5_reg_1 (.CK( clk ) , .D( u2_uk_K_r4_1 ) , .Q( u2_uk_K_r5_1 ) );
  DFF_X1 u2_uk_K_r5_reg_10 (.CK( clk ) , .D( u2_uk_K_r4_10 ) , .Q( u2_uk_K_r5_10 ) );
  DFF_X1 u2_uk_K_r5_reg_11 (.CK( clk ) , .D( u2_uk_K_r4_11 ) , .Q( u2_uk_K_r5_11 ) , .QN( u2_uk_n1457 ) );
  DFF_X1 u2_uk_K_r5_reg_12 (.CK( clk ) , .D( u2_uk_K_r4_12 ) , .Q( u2_uk_K_r5_12 ) , .QN( u2_uk_n1458 ) );
  DFF_X1 u2_uk_K_r5_reg_13 (.CK( clk ) , .D( u2_uk_K_r4_13 ) , .Q( u2_uk_K_r5_13 ) );
  DFF_X1 u2_uk_K_r5_reg_14 (.CK( clk ) , .D( u2_uk_K_r4_14 ) , .Q( u2_uk_K_r5_14 ) , .QN( u2_uk_n1459 ) );
  DFF_X1 u2_uk_K_r5_reg_15 (.CK( clk ) , .D( u2_uk_K_r4_15 ) , .Q( u2_uk_K_r5_15 ) , .QN( u2_uk_n1460 ) );
  DFF_X1 u2_uk_K_r5_reg_16 (.CK( clk ) , .D( u2_uk_K_r4_16 ) , .Q( u2_uk_K_r5_16 ) );
  DFF_X1 u2_uk_K_r5_reg_17 (.CK( clk ) , .D( u2_uk_K_r4_17 ) , .Q( u2_uk_K_r5_17 ) , .QN( u2_uk_n1461 ) );
  DFF_X1 u2_uk_K_r5_reg_18 (.CK( clk ) , .D( u2_uk_K_r4_18 ) , .Q( u2_uk_K_r5_18 ) );
  DFF_X1 u2_uk_K_r5_reg_19 (.CK( clk ) , .D( u2_uk_K_r4_19 ) , .Q( u2_uk_K_r5_19 ) );
  DFF_X1 u2_uk_K_r5_reg_2 (.CK( clk ) , .D( u2_uk_K_r4_2 ) , .Q( u2_uk_K_r5_2 ) , .QN( u2_uk_n1452 ) );
  DFF_X1 u2_uk_K_r5_reg_20 (.CK( clk ) , .D( u2_uk_K_r4_20 ) , .Q( u2_uk_K_r5_20 ) , .QN( u2_uk_n1462 ) );
  DFF_X1 u2_uk_K_r5_reg_21 (.CK( clk ) , .D( u2_uk_K_r4_21 ) , .Q( u2_uk_K_r5_21 ) );
  DFF_X1 u2_uk_K_r5_reg_22 (.CK( clk ) , .D( u2_uk_K_r4_22 ) , .Q( u2_uk_K_r5_22 ) , .QN( u2_uk_n1464 ) );
  DFF_X1 u2_uk_K_r5_reg_23 (.CK( clk ) , .D( u2_uk_K_r4_23 ) , .Q( u2_uk_K_r5_23 ) );
  DFF_X1 u2_uk_K_r5_reg_24 (.CK( clk ) , .D( u2_uk_K_r4_24 ) , .Q( u2_uk_K_r5_24 ) , .QN( u2_uk_n1465 ) );
  DFF_X1 u2_uk_K_r5_reg_25 (.CK( clk ) , .D( u2_uk_K_r4_25 ) , .Q( u2_uk_K_r5_25 ) , .QN( u2_uk_n1466 ) );
  DFF_X1 u2_uk_K_r5_reg_26 (.CK( clk ) , .D( u2_uk_K_r4_26 ) , .Q( u2_uk_K_r5_26 ) );
  DFF_X1 u2_uk_K_r5_reg_27 (.CK( clk ) , .D( u2_uk_K_r4_27 ) , .Q( u2_uk_K_r5_27 ) , .QN( u2_uk_n1468 ) );
  DFF_X1 u2_uk_K_r5_reg_28 (.CK( clk ) , .D( u2_uk_K_r4_28 ) , .Q( u2_uk_K_r5_28 ) , .QN( u2_uk_n1469 ) );
  DFF_X1 u2_uk_K_r5_reg_29 (.CK( clk ) , .D( u2_uk_K_r4_29 ) , .Q( u2_uk_K_r5_29 ) , .QN( u2_uk_n1470 ) );
  DFF_X1 u2_uk_K_r5_reg_3 (.CK( clk ) , .D( u2_uk_K_r4_3 ) , .Q( u2_uk_K_r5_3 ) , .QN( u2_uk_n1453 ) );
  DFF_X1 u2_uk_K_r5_reg_30 (.CK( clk ) , .D( u2_uk_K_r4_30 ) , .Q( u2_uk_K_r5_30 ) , .QN( u2_uk_n1471 ) );
  DFF_X1 u2_uk_K_r5_reg_31 (.CK( clk ) , .D( u2_uk_K_r4_31 ) , .Q( u2_uk_K_r5_31 ) );
  DFF_X1 u2_uk_K_r5_reg_32 (.CK( clk ) , .D( u2_uk_K_r4_32 ) , .Q( u2_uk_K_r5_32 ) );
  DFF_X1 u2_uk_K_r5_reg_33 (.CK( clk ) , .D( u2_uk_K_r4_33 ) , .Q( u2_uk_K_r5_33 ) , .QN( u2_uk_n1474 ) );
  DFF_X1 u2_uk_K_r5_reg_34 (.CK( clk ) , .D( u2_uk_K_r4_34 ) , .Q( u2_uk_K_r5_34 ) , .QN( u2_uk_n1475 ) );
  DFF_X1 u2_uk_K_r5_reg_35 (.CK( clk ) , .D( u2_uk_K_r4_35 ) , .Q( u2_uk_K_r5_35 ) , .QN( u2_uk_n1477 ) );
  DFF_X1 u2_uk_K_r5_reg_36 (.CK( clk ) , .D( u2_uk_K_r4_36 ) , .Q( u2_uk_K_r5_36 ) , .QN( u2_uk_n1478 ) );
  DFF_X1 u2_uk_K_r5_reg_37 (.CK( clk ) , .D( u2_uk_K_r4_37 ) , .Q( u2_uk_K_r5_37 ) );
  DFF_X1 u2_uk_K_r5_reg_38 (.CK( clk ) , .D( u2_uk_K_r4_38 ) , .Q( u2_uk_K_r5_38 ) , .QN( u2_uk_n1480 ) );
  DFF_X1 u2_uk_K_r5_reg_39 (.CK( clk ) , .D( u2_uk_K_r4_39 ) , .Q( u2_uk_K_r5_39 ) );
  DFF_X1 u2_uk_K_r5_reg_4 (.CK( clk ) , .D( u2_uk_K_r4_4 ) , .Q( u2_uk_K_r5_4 ) );
  DFF_X1 u2_uk_K_r5_reg_40 (.CK( clk ) , .D( u2_uk_K_r4_40 ) , .Q( u2_uk_K_r5_40 ) );
  DFF_X1 u2_uk_K_r5_reg_41 (.CK( clk ) , .D( u2_uk_K_r4_41 ) , .Q( u2_uk_K_r5_41 ) );
  DFF_X1 u2_uk_K_r5_reg_42 (.CK( clk ) , .D( u2_uk_K_r4_42 ) , .Q( u2_uk_K_r5_42 ) , .QN( u2_uk_n1484 ) );
  DFF_X1 u2_uk_K_r5_reg_43 (.CK( clk ) , .D( u2_uk_K_r4_43 ) , .Q( u2_uk_K_r5_43 ) );
  DFF_X1 u2_uk_K_r5_reg_44 (.CK( clk ) , .D( u2_uk_K_r4_44 ) , .Q( u2_uk_K_r5_44 ) , .QN( u2_uk_n1486 ) );
  DFF_X1 u2_uk_K_r5_reg_45 (.CK( clk ) , .D( u2_uk_K_r4_45 ) , .Q( u2_uk_K_r5_45 ) );
  DFF_X1 u2_uk_K_r5_reg_46 (.CK( clk ) , .D( u2_uk_K_r4_46 ) , .Q( u2_uk_K_r5_46 ) , .QN( u2_uk_n1487 ) );
  DFF_X1 u2_uk_K_r5_reg_47 (.CK( clk ) , .D( u2_uk_K_r4_47 ) , .Q( u2_uk_K_r5_47 ) , .QN( u2_uk_n1488 ) );
  DFF_X1 u2_uk_K_r5_reg_48 (.CK( clk ) , .D( u2_uk_K_r4_48 ) , .Q( u2_uk_K_r5_48 ) );
  DFF_X1 u2_uk_K_r5_reg_49 (.CK( clk ) , .D( u2_uk_K_r4_49 ) , .Q( u2_uk_K_r5_49 ) , .QN( u2_uk_n1490 ) );
  DFF_X1 u2_uk_K_r5_reg_5 (.CK( clk ) , .D( u2_uk_K_r4_5 ) , .Q( u2_uk_K_r5_5 ) );
  DFF_X1 u2_uk_K_r5_reg_50 (.CK( clk ) , .D( u2_uk_K_r4_50 ) , .Q( u2_uk_K_r5_50 ) , .QN( u2_uk_n1491 ) );
  DFF_X1 u2_uk_K_r5_reg_51 (.CK( clk ) , .D( u2_uk_K_r4_51 ) , .Q( u2_uk_K_r5_51 ) );
  DFF_X1 u2_uk_K_r5_reg_52 (.CK( clk ) , .D( u2_uk_K_r4_52 ) , .Q( u2_uk_K_r5_52 ) , .QN( u2_uk_n1493 ) );
  DFF_X1 u2_uk_K_r5_reg_53 (.CK( clk ) , .D( u2_uk_K_r4_53 ) , .Q( u2_uk_K_r5_53 ) , .QN( u2_uk_n1494 ) );
  DFF_X1 u2_uk_K_r5_reg_54 (.CK( clk ) , .D( u2_uk_K_r4_54 ) , .Q( u2_uk_K_r5_54 ) , .QN( u2_uk_n1496 ) );
  DFF_X1 u2_uk_K_r5_reg_55 (.CK( clk ) , .D( u2_uk_K_r4_55 ) , .Q( u2_uk_K_r5_55 ) , .QN( u2_uk_n1497 ) );
  DFF_X1 u2_uk_K_r5_reg_6 (.CK( clk ) , .D( u2_uk_K_r4_6 ) , .Q( u2_uk_K_r5_6 ) , .QN( u2_uk_n1454 ) );
  DFF_X1 u2_uk_K_r5_reg_7 (.CK( clk ) , .D( u2_uk_K_r4_7 ) , .Q( u2_uk_K_r5_7 ) , .QN( u2_uk_n1455 ) );
  DFF_X1 u2_uk_K_r5_reg_8 (.CK( clk ) , .D( u2_uk_K_r4_8 ) , .Q( u2_uk_K_r5_8 ) );
  DFF_X1 u2_uk_K_r5_reg_9 (.CK( clk ) , .D( u2_uk_K_r4_9 ) , .Q( u2_uk_K_r5_9 ) , .QN( u2_uk_n1456 ) );
  DFF_X1 u2_uk_K_r6_reg_0 (.CK( clk ) , .D( u2_uk_K_r5_0 ) , .Q( u2_uk_K_r6_0 ) );
  DFF_X1 u2_uk_K_r6_reg_1 (.CK( clk ) , .D( u2_uk_K_r5_1 ) , .Q( u2_uk_K_r6_1 ) , .QN( u2_uk_n1498 ) );
  DFF_X1 u2_uk_K_r6_reg_10 (.CK( clk ) , .D( u2_uk_K_r5_10 ) , .Q( u2_uk_K_r6_10 ) );
  DFF_X1 u2_uk_K_r6_reg_11 (.CK( clk ) , .D( u2_uk_K_r5_11 ) , .Q( u2_uk_K_r6_11 ) , .QN( u2_uk_n1506 ) );
  DFF_X1 u2_uk_K_r6_reg_12 (.CK( clk ) , .D( u2_uk_K_r5_12 ) , .Q( u2_uk_K_r6_12 ) , .QN( u2_uk_n1507 ) );
  DFF_X1 u2_uk_K_r6_reg_13 (.CK( clk ) , .D( u2_uk_K_r5_13 ) , .Q( u2_uk_K_r6_13 ) , .QN( u2_uk_n1508 ) );
  DFF_X1 u2_uk_K_r6_reg_14 (.CK( clk ) , .D( u2_uk_K_r5_14 ) , .Q( u2_uk_K_r6_14 ) );
  DFF_X1 u2_uk_K_r6_reg_15 (.CK( clk ) , .D( u2_uk_K_r5_15 ) , .Q( u2_uk_K_r6_15 ) , .QN( u2_uk_n1510 ) );
  DFF_X1 u2_uk_K_r6_reg_16 (.CK( clk ) , .D( u2_uk_K_r5_16 ) , .Q( u2_uk_K_r6_16 ) , .QN( u2_uk_n1511 ) );
  DFF_X1 u2_uk_K_r6_reg_17 (.CK( clk ) , .D( u2_uk_K_r5_17 ) , .Q( u2_uk_K_r6_17 ) , .QN( u2_uk_n1513 ) );
  DFF_X1 u2_uk_K_r6_reg_18 (.CK( clk ) , .D( u2_uk_K_r5_18 ) , .Q( u2_uk_K_r6_18 ) , .QN( u2_uk_n1514 ) );
  DFF_X1 u2_uk_K_r6_reg_19 (.CK( clk ) , .D( u2_uk_K_r5_19 ) , .Q( u2_uk_K_r6_19 ) );
  DFF_X1 u2_uk_K_r6_reg_2 (.CK( clk ) , .D( u2_uk_K_r5_2 ) , .Q( u2_uk_K_r6_2 ) , .QN( u2_uk_n1499 ) );
  DFF_X1 u2_uk_K_r6_reg_20 (.CK( clk ) , .D( u2_uk_K_r5_20 ) , .Q( u2_uk_K_r6_20 ) , .QN( u2_uk_n1515 ) );
  DFF_X1 u2_uk_K_r6_reg_21 (.CK( clk ) , .D( u2_uk_K_r5_21 ) , .Q( u2_uk_K_r6_21 ) );
  DFF_X1 u2_uk_K_r6_reg_22 (.CK( clk ) , .D( u2_uk_K_r5_22 ) , .Q( u2_uk_K_r6_22 ) );
  DFF_X1 u2_uk_K_r6_reg_23 (.CK( clk ) , .D( u2_uk_K_r5_23 ) , .Q( u2_uk_K_r6_23 ) , .QN( u2_uk_n1517 ) );
  DFF_X1 u2_uk_K_r6_reg_24 (.CK( clk ) , .D( u2_uk_K_r5_24 ) , .Q( u2_uk_K_r6_24 ) , .QN( u2_uk_n1518 ) );
  DFF_X1 u2_uk_K_r6_reg_25 (.CK( clk ) , .D( u2_uk_K_r5_25 ) , .Q( u2_uk_K_r6_25 ) , .QN( u2_uk_n1519 ) );
  DFF_X1 u2_uk_K_r6_reg_26 (.CK( clk ) , .D( u2_uk_K_r5_26 ) , .Q( u2_uk_K_r6_26 ) );
  DFF_X1 u2_uk_K_r6_reg_27 (.CK( clk ) , .D( u2_uk_K_r5_27 ) , .Q( u2_uk_K_r6_27 ) );
  DFF_X1 u2_uk_K_r6_reg_28 (.CK( clk ) , .D( u2_uk_K_r5_28 ) , .Q( u2_uk_K_r6_28 ) );
  DFF_X1 u2_uk_K_r6_reg_29 (.CK( clk ) , .D( u2_uk_K_r5_29 ) , .Q( u2_uk_K_r6_29 ) );
  DFF_X1 u2_uk_K_r6_reg_3 (.CK( clk ) , .D( u2_uk_K_r5_3 ) , .Q( u2_uk_K_r6_3 ) );
  DFF_X1 u2_uk_K_r6_reg_30 (.CK( clk ) , .D( u2_uk_K_r5_30 ) , .Q( u2_uk_K_r6_30 ) );
  DFF_X1 u2_uk_K_r6_reg_31 (.CK( clk ) , .D( u2_uk_K_r5_31 ) , .Q( u2_uk_K_r6_31 ) );
  DFF_X1 u2_uk_K_r6_reg_32 (.CK( clk ) , .D( u2_uk_K_r5_32 ) , .Q( u2_uk_K_r6_32 ) , .QN( u2_uk_n1521 ) );
  DFF_X1 u2_uk_K_r6_reg_33 (.CK( clk ) , .D( u2_uk_K_r5_33 ) , .Q( u2_uk_K_r6_33 ) , .QN( u2_uk_n1522 ) );
  DFF_X1 u2_uk_K_r6_reg_34 (.CK( clk ) , .D( u2_uk_K_r5_34 ) , .Q( u2_uk_K_r6_34 ) );
  DFF_X1 u2_uk_K_r6_reg_35 (.CK( clk ) , .D( u2_uk_K_r5_35 ) , .Q( u2_uk_K_r6_35 ) , .QN( u2_uk_n1524 ) );
  DFF_X1 u2_uk_K_r6_reg_36 (.CK( clk ) , .D( u2_uk_K_r5_36 ) , .Q( u2_uk_K_r6_36 ) , .QN( u2_uk_n1525 ) );
  DFF_X1 u2_uk_K_r6_reg_37 (.CK( clk ) , .D( u2_uk_K_r5_37 ) , .Q( u2_uk_K_r6_37 ) );
  DFF_X1 u2_uk_K_r6_reg_38 (.CK( clk ) , .D( u2_uk_K_r5_38 ) , .Q( u2_uk_K_r6_38 ) , .QN( u2_uk_n1526 ) );
  DFF_X1 u2_uk_K_r6_reg_39 (.CK( clk ) , .D( u2_uk_K_r5_39 ) , .Q( u2_uk_K_r6_39 ) , .QN( u2_uk_n1527 ) );
  DFF_X1 u2_uk_K_r6_reg_4 (.CK( clk ) , .D( u2_uk_K_r5_4 ) , .Q( u2_uk_K_r6_4 ) , .QN( u2_uk_n1500 ) );
  DFF_X1 u2_uk_K_r6_reg_40 (.CK( clk ) , .D( u2_uk_K_r5_40 ) , .Q( u2_uk_K_r6_40 ) , .QN( u2_uk_n1528 ) );
  DFF_X1 u2_uk_K_r6_reg_41 (.CK( clk ) , .D( u2_uk_K_r5_41 ) , .Q( u2_uk_K_r6_41 ) , .QN( u2_uk_n1529 ) );
  DFF_X1 u2_uk_K_r6_reg_42 (.CK( clk ) , .D( u2_uk_K_r5_42 ) , .Q( u2_uk_K_r6_42 ) , .QN( u2_uk_n1530 ) );
  DFF_X1 u2_uk_K_r6_reg_43 (.CK( clk ) , .D( u2_uk_K_r5_43 ) , .Q( u2_uk_K_r6_43 ) , .QN( u2_uk_n1531 ) );
  DFF_X1 u2_uk_K_r6_reg_44 (.CK( clk ) , .D( u2_uk_K_r5_44 ) , .Q( u2_uk_K_r6_44 ) , .QN( u2_uk_n1532 ) );
  DFF_X1 u2_uk_K_r6_reg_45 (.CK( clk ) , .D( u2_uk_K_r5_45 ) , .Q( u2_uk_K_r6_45 ) , .QN( u2_uk_n1533 ) );
  DFF_X1 u2_uk_K_r6_reg_46 (.CK( clk ) , .D( u2_uk_K_r5_46 ) , .Q( u2_uk_K_r6_46 ) );
  DFF_X1 u2_uk_K_r6_reg_47 (.CK( clk ) , .D( u2_uk_K_r5_47 ) , .Q( u2_uk_K_r6_47 ) , .QN( u2_uk_n1534 ) );
  DFF_X1 u2_uk_K_r6_reg_48 (.CK( clk ) , .D( u2_uk_K_r5_48 ) , .Q( u2_uk_K_r6_48 ) , .QN( u2_uk_n1535 ) );
  DFF_X1 u2_uk_K_r6_reg_49 (.CK( clk ) , .D( u2_uk_K_r5_49 ) , .Q( u2_uk_K_r6_49 ) , .QN( u2_uk_n1536 ) );
  DFF_X1 u2_uk_K_r6_reg_5 (.CK( clk ) , .D( u2_uk_K_r5_5 ) , .Q( u2_uk_K_r6_5 ) , .QN( u2_uk_n1501 ) );
  DFF_X1 u2_uk_K_r6_reg_50 (.CK( clk ) , .D( u2_uk_K_r5_50 ) , .Q( u2_uk_K_r6_50 ) , .QN( u2_uk_n1537 ) );
  DFF_X1 u2_uk_K_r6_reg_51 (.CK( clk ) , .D( u2_uk_K_r5_51 ) , .Q( u2_uk_K_r6_51 ) );
  DFF_X1 u2_uk_K_r6_reg_52 (.CK( clk ) , .D( u2_uk_K_r5_52 ) , .Q( u2_uk_K_r6_52 ) , .QN( u2_uk_n1538 ) );
  DFF_X1 u2_uk_K_r6_reg_53 (.CK( clk ) , .D( u2_uk_K_r5_53 ) , .Q( u2_uk_K_r6_53 ) );
  DFF_X1 u2_uk_K_r6_reg_54 (.CK( clk ) , .D( u2_uk_K_r5_54 ) , .Q( u2_uk_K_r6_54 ) , .QN( u2_uk_n1540 ) );
  DFF_X1 u2_uk_K_r6_reg_55 (.CK( clk ) , .D( u2_uk_K_r5_55 ) , .Q( u2_uk_K_r6_55 ) );
  DFF_X1 u2_uk_K_r6_reg_6 (.CK( clk ) , .D( u2_uk_K_r5_6 ) , .Q( u2_uk_K_r6_6 ) , .QN( u2_uk_n1502 ) );
  DFF_X1 u2_uk_K_r6_reg_7 (.CK( clk ) , .D( u2_uk_K_r5_7 ) , .Q( u2_uk_K_r6_7 ) );
  DFF_X1 u2_uk_K_r6_reg_8 (.CK( clk ) , .D( u2_uk_K_r5_8 ) , .Q( u2_uk_K_r6_8 ) , .QN( u2_uk_n1503 ) );
  DFF_X1 u2_uk_K_r6_reg_9 (.CK( clk ) , .D( u2_uk_K_r5_9 ) , .Q( u2_uk_K_r6_9 ) , .QN( u2_uk_n1504 ) );
  DFF_X1 u2_uk_K_r7_reg_0 (.CK( clk ) , .D( u2_uk_K_r6_0 ) , .Q( u2_uk_K_r7_0 ) );
  DFF_X1 u2_uk_K_r7_reg_1 (.CK( clk ) , .D( u2_uk_K_r6_1 ) , .Q( u2_uk_K_r7_1 ) , .QN( u2_uk_n1541 ) );
  DFF_X1 u2_uk_K_r7_reg_10 (.CK( clk ) , .D( u2_uk_K_r6_10 ) , .Q( u2_uk_K_r7_10 ) , .QN( u2_uk_n1547 ) );
  DFF_X1 u2_uk_K_r7_reg_11 (.CK( clk ) , .D( u2_uk_K_r6_11 ) , .Q( u2_uk_K_r7_11 ) , .QN( u2_uk_n1548 ) );
  DFF_X1 u2_uk_K_r7_reg_12 (.CK( clk ) , .D( u2_uk_K_r6_12 ) , .Q( u2_uk_K_r7_12 ) , .QN( u2_uk_n1549 ) );
  DFF_X1 u2_uk_K_r7_reg_13 (.CK( clk ) , .D( u2_uk_K_r6_13 ) , .Q( u2_uk_K_r7_13 ) );
  DFF_X1 u2_uk_K_r7_reg_14 (.CK( clk ) , .D( u2_uk_K_r6_14 ) , .Q( u2_uk_K_r7_14 ) , .QN( u2_uk_n1551 ) );
  DFF_X1 u2_uk_K_r7_reg_15 (.CK( clk ) , .D( u2_uk_K_r6_15 ) , .Q( u2_uk_K_r7_15 ) );
  DFF_X1 u2_uk_K_r7_reg_16 (.CK( clk ) , .D( u2_uk_K_r6_16 ) , .Q( u2_uk_K_r7_16 ) );
  DFF_X1 u2_uk_K_r7_reg_17 (.CK( clk ) , .D( u2_uk_K_r6_17 ) , .Q( u2_uk_K_r7_17 ) , .QN( u2_uk_n1554 ) );
  DFF_X1 u2_uk_K_r7_reg_18 (.CK( clk ) , .D( u2_uk_K_r6_18 ) , .Q( u2_uk_K_r7_18 ) , .QN( u2_uk_n1555 ) );
  DFF_X1 u2_uk_K_r7_reg_19 (.CK( clk ) , .D( u2_uk_K_r6_19 ) , .Q( u2_uk_K_r7_19 ) , .QN( u2_uk_n1556 ) );
  DFF_X1 u2_uk_K_r7_reg_2 (.CK( clk ) , .D( u2_uk_K_r6_2 ) , .Q( u2_uk_K_r7_2 ) , .QN( u2_uk_n1542 ) );
  DFF_X1 u2_uk_K_r7_reg_20 (.CK( clk ) , .D( u2_uk_K_r6_20 ) , .Q( u2_uk_K_r7_20 ) );
  DFF_X1 u2_uk_K_r7_reg_21 (.CK( clk ) , .D( u2_uk_K_r6_21 ) , .Q( u2_uk_K_r7_21 ) , .QN( u2_uk_n1558 ) );
  DFF_X1 u2_uk_K_r7_reg_22 (.CK( clk ) , .D( u2_uk_K_r6_22 ) , .Q( u2_uk_K_r7_22 ) );
  DFF_X1 u2_uk_K_r7_reg_23 (.CK( clk ) , .D( u2_uk_K_r6_23 ) , .Q( u2_uk_K_r7_23 ) );
  DFF_X1 u2_uk_K_r7_reg_24 (.CK( clk ) , .D( u2_uk_K_r6_24 ) , .Q( u2_uk_K_r7_24 ) , .QN( u2_uk_n1562 ) );
  DFF_X1 u2_uk_K_r7_reg_25 (.CK( clk ) , .D( u2_uk_K_r6_25 ) , .Q( u2_uk_K_r7_25 ) , .QN( u2_uk_n1563 ) );
  DFF_X1 u2_uk_K_r7_reg_26 (.CK( clk ) , .D( u2_uk_K_r6_26 ) , .Q( u2_uk_K_r7_26 ) );
  DFF_X1 u2_uk_K_r7_reg_27 (.CK( clk ) , .D( u2_uk_K_r6_27 ) , .Q( u2_uk_K_r7_27 ) );
  DFF_X1 u2_uk_K_r7_reg_28 (.CK( clk ) , .D( u2_uk_K_r6_28 ) , .Q( u2_uk_K_r7_28 ) , .QN( u2_uk_n1565 ) );
  DFF_X1 u2_uk_K_r7_reg_29 (.CK( clk ) , .D( u2_uk_K_r6_29 ) , .Q( u2_uk_K_r7_29 ) );
  DFF_X1 u2_uk_K_r7_reg_3 (.CK( clk ) , .D( u2_uk_K_r6_3 ) , .Q( u2_uk_K_r7_3 ) , .QN( u2_uk_n1543 ) );
  DFF_X1 u2_uk_K_r7_reg_30 (.CK( clk ) , .D( u2_uk_K_r6_30 ) , .Q( u2_uk_K_r7_30 ) );
  DFF_X1 u2_uk_K_r7_reg_31 (.CK( clk ) , .D( u2_uk_K_r6_31 ) , .Q( u2_uk_K_r7_31 ) );
  DFF_X1 u2_uk_K_r7_reg_32 (.CK( clk ) , .D( u2_uk_K_r6_32 ) , .Q( u2_uk_K_r7_32 ) );
  DFF_X1 u2_uk_K_r7_reg_33 (.CK( clk ) , .D( u2_uk_K_r6_33 ) , .Q( u2_uk_K_r7_33 ) , .QN( u2_uk_n1568 ) );
  DFF_X1 u2_uk_K_r7_reg_34 (.CK( clk ) , .D( u2_uk_K_r6_34 ) , .Q( u2_uk_K_r7_34 ) );
  DFF_X1 u2_uk_K_r7_reg_35 (.CK( clk ) , .D( u2_uk_K_r6_35 ) , .Q( u2_uk_K_r7_35 ) , .QN( u2_uk_n1569 ) );
  DFF_X1 u2_uk_K_r7_reg_36 (.CK( clk ) , .D( u2_uk_K_r6_36 ) , .Q( u2_uk_K_r7_36 ) , .QN( u2_uk_n1570 ) );
  DFF_X1 u2_uk_K_r7_reg_37 (.CK( clk ) , .D( u2_uk_K_r6_37 ) , .Q( u2_uk_K_r7_37 ) );
  DFF_X1 u2_uk_K_r7_reg_38 (.CK( clk ) , .D( u2_uk_K_r6_38 ) , .Q( u2_uk_K_r7_38 ) , .QN( u2_uk_n1571 ) );
  DFF_X1 u2_uk_K_r7_reg_39 (.CK( clk ) , .D( u2_uk_K_r6_39 ) , .Q( u2_uk_K_r7_39 ) );
  DFF_X1 u2_uk_K_r7_reg_4 (.CK( clk ) , .D( u2_uk_K_r6_4 ) , .Q( u2_uk_K_r7_4 ) , .QN( u2_uk_n1544 ) );
  DFF_X1 u2_uk_K_r7_reg_40 (.CK( clk ) , .D( u2_uk_K_r6_40 ) , .Q( u2_uk_K_r7_40 ) , .QN( u2_uk_n1573 ) );
  DFF_X1 u2_uk_K_r7_reg_41 (.CK( clk ) , .D( u2_uk_K_r6_41 ) , .Q( u2_uk_K_r7_41 ) , .QN( u2_uk_n1574 ) );
  DFF_X1 u2_uk_K_r7_reg_42 (.CK( clk ) , .D( u2_uk_K_r6_42 ) , .Q( u2_uk_K_r7_42 ) , .QN( u2_uk_n1575 ) );
  DFF_X1 u2_uk_K_r7_reg_43 (.CK( clk ) , .D( u2_uk_K_r6_43 ) , .Q( u2_uk_K_r7_43 ) , .QN( u2_uk_n1576 ) );
  DFF_X1 u2_uk_K_r7_reg_44 (.CK( clk ) , .D( u2_uk_K_r6_44 ) , .Q( u2_uk_K_r7_44 ) , .QN( u2_uk_n1577 ) );
  DFF_X1 u2_uk_K_r7_reg_45 (.CK( clk ) , .D( u2_uk_K_r6_45 ) , .Q( u2_uk_K_r7_45 ) , .QN( u2_uk_n1578 ) );
  DFF_X1 u2_uk_K_r7_reg_46 (.CK( clk ) , .D( u2_uk_K_r6_46 ) , .Q( u2_uk_K_r7_46 ) );
  DFF_X1 u2_uk_K_r7_reg_47 (.CK( clk ) , .D( u2_uk_K_r6_47 ) , .Q( u2_uk_K_r7_47 ) , .QN( u2_uk_n1580 ) );
  DFF_X1 u2_uk_K_r7_reg_48 (.CK( clk ) , .D( u2_uk_K_r6_48 ) , .Q( u2_uk_K_r7_48 ) );
  DFF_X1 u2_uk_K_r7_reg_49 (.CK( clk ) , .D( u2_uk_K_r6_49 ) , .Q( u2_uk_K_r7_49 ) , .QN( u2_uk_n1582 ) );
  DFF_X1 u2_uk_K_r7_reg_5 (.CK( clk ) , .D( u2_uk_K_r6_5 ) , .Q( u2_uk_K_r7_5 ) );
  DFF_X1 u2_uk_K_r7_reg_50 (.CK( clk ) , .D( u2_uk_K_r6_50 ) , .Q( u2_uk_K_r7_50 ) , .QN( u2_uk_n1583 ) );
  DFF_X1 u2_uk_K_r7_reg_51 (.CK( clk ) , .D( u2_uk_K_r6_51 ) , .Q( u2_uk_K_r7_51 ) , .QN( u2_uk_n1584 ) );
  DFF_X1 u2_uk_K_r7_reg_52 (.CK( clk ) , .D( u2_uk_K_r6_52 ) , .Q( u2_uk_K_r7_52 ) , .QN( u2_uk_n1585 ) );
  DFF_X1 u2_uk_K_r7_reg_53 (.CK( clk ) , .D( u2_uk_K_r6_53 ) , .Q( u2_uk_K_r7_53 ) );
  DFF_X1 u2_uk_K_r7_reg_54 (.CK( clk ) , .D( u2_uk_K_r6_54 ) , .Q( u2_uk_K_r7_54 ) , .QN( u2_uk_n1586 ) );
  DFF_X1 u2_uk_K_r7_reg_55 (.CK( clk ) , .D( u2_uk_K_r6_55 ) , .Q( u2_uk_K_r7_55 ) );
  DFF_X1 u2_uk_K_r7_reg_6 (.CK( clk ) , .D( u2_uk_K_r6_6 ) , .Q( u2_uk_K_r7_6 ) );
  DFF_X1 u2_uk_K_r7_reg_7 (.CK( clk ) , .D( u2_uk_K_r6_7 ) , .Q( u2_uk_K_r7_7 ) );
  DFF_X1 u2_uk_K_r7_reg_8 (.CK( clk ) , .D( u2_uk_K_r6_8 ) , .Q( u2_uk_K_r7_8 ) );
  DFF_X1 u2_uk_K_r7_reg_9 (.CK( clk ) , .D( u2_uk_K_r6_9 ) , .Q( u2_uk_K_r7_9 ) );
  DFF_X1 u2_uk_K_r8_reg_0 (.CK( clk ) , .D( u2_uk_K_r7_0 ) , .Q( u2_uk_K_r8_0 ) , .QN( u2_uk_n1588 ) );
  DFF_X1 u2_uk_K_r8_reg_1 (.CK( clk ) , .D( u2_uk_K_r7_1 ) , .Q( u2_uk_K_r8_1 ) , .QN( u2_uk_n1589 ) );
  DFF_X1 u2_uk_K_r8_reg_10 (.CK( clk ) , .D( u2_uk_K_r7_10 ) , .Q( u2_uk_K_r8_10 ) );
  DFF_X1 u2_uk_K_r8_reg_11 (.CK( clk ) , .D( u2_uk_K_r7_11 ) , .Q( u2_uk_K_r8_11 ) , .QN( u2_uk_n1595 ) );
  DFF_X1 u2_uk_K_r8_reg_12 (.CK( clk ) , .D( u2_uk_K_r7_12 ) , .Q( u2_uk_K_r8_12 ) , .QN( u2_uk_n1596 ) );
  DFF_X1 u2_uk_K_r8_reg_13 (.CK( clk ) , .D( u2_uk_K_r7_13 ) , .Q( u2_uk_K_r8_13 ) );
  DFF_X1 u2_uk_K_r8_reg_14 (.CK( clk ) , .D( u2_uk_K_r7_14 ) , .Q( u2_uk_K_r8_14 ) , .QN( u2_uk_n1597 ) );
  DFF_X1 u2_uk_K_r8_reg_15 (.CK( clk ) , .D( u2_uk_K_r7_15 ) , .Q( u2_uk_K_r8_15 ) , .QN( u2_uk_n1598 ) );
  DFF_X1 u2_uk_K_r8_reg_16 (.CK( clk ) , .D( u2_uk_K_r7_16 ) , .Q( u2_uk_K_r8_16 ) );
  DFF_X1 u2_uk_K_r8_reg_17 (.CK( clk ) , .D( u2_uk_K_r7_17 ) , .Q( u2_uk_K_r8_17 ) );
  DFF_X1 u2_uk_K_r8_reg_18 (.CK( clk ) , .D( u2_uk_K_r7_18 ) , .Q( u2_uk_K_r8_18 ) , .QN( u2_uk_n1599 ) );
  DFF_X1 u2_uk_K_r8_reg_19 (.CK( clk ) , .D( u2_uk_K_r7_19 ) , .Q( u2_uk_K_r8_19 ) );
  DFF_X1 u2_uk_K_r8_reg_2 (.CK( clk ) , .D( u2_uk_K_r7_2 ) , .Q( u2_uk_K_r8_2 ) );
  DFF_X1 u2_uk_K_r8_reg_20 (.CK( clk ) , .D( u2_uk_K_r7_20 ) , .Q( u2_uk_K_r8_20 ) , .QN( u2_uk_n1600 ) );
  DFF_X1 u2_uk_K_r8_reg_21 (.CK( clk ) , .D( u2_uk_K_r7_21 ) , .Q( u2_uk_K_r8_21 ) );
  DFF_X1 u2_uk_K_r8_reg_22 (.CK( clk ) , .D( u2_uk_K_r7_22 ) , .Q( u2_uk_K_r8_22 ) );
  DFF_X1 u2_uk_K_r8_reg_23 (.CK( clk ) , .D( u2_uk_K_r7_23 ) , .Q( u2_uk_K_r8_23 ) , .QN( u2_uk_n1602 ) );
  DFF_X1 u2_uk_K_r8_reg_24 (.CK( clk ) , .D( u2_uk_K_r7_24 ) , .Q( u2_uk_K_r8_24 ) , .QN( u2_uk_n1603 ) );
  DFF_X1 u2_uk_K_r8_reg_25 (.CK( clk ) , .D( u2_uk_K_r7_25 ) , .Q( u2_uk_K_r8_25 ) , .QN( u2_uk_n1604 ) );
  DFF_X1 u2_uk_K_r8_reg_26 (.CK( clk ) , .D( u2_uk_K_r7_26 ) , .Q( u2_uk_K_r8_26 ) , .QN( u2_uk_n1605 ) );
  DFF_X1 u2_uk_K_r8_reg_27 (.CK( clk ) , .D( u2_uk_K_r7_27 ) , .Q( u2_uk_K_r8_27 ) );
  DFF_X1 u2_uk_K_r8_reg_28 (.CK( clk ) , .D( u2_uk_K_r7_28 ) , .Q( u2_uk_K_r8_28 ) );
  DFF_X1 u2_uk_K_r8_reg_29 (.CK( clk ) , .D( u2_uk_K_r7_29 ) , .Q( u2_uk_K_r8_29 ) , .QN( u2_uk_n1609 ) );
  DFF_X1 u2_uk_K_r8_reg_3 (.CK( clk ) , .D( u2_uk_K_r7_3 ) , .Q( u2_uk_K_r8_3 ) , .QN( u2_uk_n1590 ) );
  DFF_X1 u2_uk_K_r8_reg_30 (.CK( clk ) , .D( u2_uk_K_r7_30 ) , .Q( u2_uk_K_r8_30 ) , .QN( u2_uk_n1610 ) );
  DFF_X1 u2_uk_K_r8_reg_31 (.CK( clk ) , .D( u2_uk_K_r7_31 ) , .Q( u2_uk_K_r8_31 ) , .QN( u2_uk_n1611 ) );
  DFF_X1 u2_uk_K_r8_reg_32 (.CK( clk ) , .D( u2_uk_K_r7_32 ) , .Q( u2_uk_K_r8_32 ) );
  DFF_X1 u2_uk_K_r8_reg_33 (.CK( clk ) , .D( u2_uk_K_r7_33 ) , .Q( u2_uk_K_r8_33 ) , .QN( u2_uk_n1612 ) );
  DFF_X1 u2_uk_K_r8_reg_34 (.CK( clk ) , .D( u2_uk_K_r7_34 ) , .Q( u2_uk_K_r8_34 ) , .QN( u2_uk_n1613 ) );
  DFF_X1 u2_uk_K_r8_reg_35 (.CK( clk ) , .D( u2_uk_K_r7_35 ) , .Q( u2_uk_K_r8_35 ) , .QN( u2_uk_n1614 ) );
  DFF_X1 u2_uk_K_r8_reg_36 (.CK( clk ) , .D( u2_uk_K_r7_36 ) , .Q( u2_uk_K_r8_36 ) , .QN( u2_uk_n1615 ) );
  DFF_X1 u2_uk_K_r8_reg_37 (.CK( clk ) , .D( u2_uk_K_r7_37 ) , .Q( u2_uk_K_r8_37 ) );
  DFF_X1 u2_uk_K_r8_reg_38 (.CK( clk ) , .D( u2_uk_K_r7_38 ) , .Q( u2_uk_K_r8_38 ) , .QN( u2_uk_n1617 ) );
  DFF_X1 u2_uk_K_r8_reg_39 (.CK( clk ) , .D( u2_uk_K_r7_39 ) , .Q( u2_uk_K_r8_39 ) , .QN( u2_uk_n1619 ) );
  DFF_X1 u2_uk_K_r8_reg_4 (.CK( clk ) , .D( u2_uk_K_r7_4 ) , .Q( u2_uk_K_r8_4 ) , .QN( u2_uk_n1591 ) );
  DFF_X1 u2_uk_K_r8_reg_40 (.CK( clk ) , .D( u2_uk_K_r7_40 ) , .Q( u2_uk_K_r8_40 ) );
  DFF_X1 u2_uk_K_r8_reg_41 (.CK( clk ) , .D( u2_uk_K_r7_41 ) , .Q( u2_uk_K_r8_41 ) );
  DFF_X1 u2_uk_K_r8_reg_42 (.CK( clk ) , .D( u2_uk_K_r7_42 ) , .Q( u2_uk_K_r8_42 ) , .QN( u2_uk_n1621 ) );
  DFF_X1 u2_uk_K_r8_reg_43 (.CK( clk ) , .D( u2_uk_K_r7_43 ) , .Q( u2_uk_K_r8_43 ) );
  DFF_X1 u2_uk_K_r8_reg_44 (.CK( clk ) , .D( u2_uk_K_r7_44 ) , .Q( u2_uk_K_r8_44 ) , .QN( u2_uk_n1622 ) );
  DFF_X1 u2_uk_K_r8_reg_45 (.CK( clk ) , .D( u2_uk_K_r7_45 ) , .Q( u2_uk_K_r8_45 ) );
  DFF_X1 u2_uk_K_r8_reg_46 (.CK( clk ) , .D( u2_uk_K_r7_46 ) , .Q( u2_uk_K_r8_46 ) , .QN( u2_uk_n1623 ) );
  DFF_X1 u2_uk_K_r8_reg_47 (.CK( clk ) , .D( u2_uk_K_r7_47 ) , .Q( u2_uk_K_r8_47 ) , .QN( u2_uk_n1624 ) );
  DFF_X1 u2_uk_K_r8_reg_48 (.CK( clk ) , .D( u2_uk_K_r7_48 ) , .Q( u2_uk_K_r8_48 ) );
  DFF_X1 u2_uk_K_r8_reg_49 (.CK( clk ) , .D( u2_uk_K_r7_49 ) , .Q( u2_uk_K_r8_49 ) , .QN( u2_uk_n1625 ) );
  DFF_X1 u2_uk_K_r8_reg_5 (.CK( clk ) , .D( u2_uk_K_r7_5 ) , .Q( u2_uk_K_r8_5 ) );
  DFF_X1 u2_uk_K_r8_reg_50 (.CK( clk ) , .D( u2_uk_K_r7_50 ) , .Q( u2_uk_K_r8_50 ) , .QN( u2_uk_n1626 ) );
  DFF_X1 u2_uk_K_r8_reg_51 (.CK( clk ) , .D( u2_uk_K_r7_51 ) , .Q( u2_uk_K_r8_51 ) );
  DFF_X1 u2_uk_K_r8_reg_52 (.CK( clk ) , .D( u2_uk_K_r7_52 ) , .Q( u2_uk_K_r8_52 ) );
  DFF_X1 u2_uk_K_r8_reg_53 (.CK( clk ) , .D( u2_uk_K_r7_53 ) , .Q( u2_uk_K_r8_53 ) , .QN( u2_uk_n1629 ) );
  DFF_X1 u2_uk_K_r8_reg_54 (.CK( clk ) , .D( u2_uk_K_r7_54 ) , .Q( u2_uk_K_r8_54 ) , .QN( u2_uk_n1630 ) );
  DFF_X1 u2_uk_K_r8_reg_55 (.CK( clk ) , .D( u2_uk_K_r7_55 ) , .Q( u2_uk_K_r8_55 ) , .QN( u2_uk_n1631 ) );
  DFF_X1 u2_uk_K_r8_reg_6 (.CK( clk ) , .D( u2_uk_K_r7_6 ) , .Q( u2_uk_K_r8_6 ) , .QN( u2_uk_n1592 ) );
  DFF_X1 u2_uk_K_r8_reg_7 (.CK( clk ) , .D( u2_uk_K_r7_7 ) , .Q( u2_uk_K_r8_7 ) , .QN( u2_uk_n1593 ) );
  DFF_X1 u2_uk_K_r8_reg_8 (.CK( clk ) , .D( u2_uk_K_r7_8 ) , .Q( u2_uk_K_r8_8 ) );
  DFF_X1 u2_uk_K_r8_reg_9 (.CK( clk ) , .D( u2_uk_K_r7_9 ) , .Q( u2_uk_K_r8_9 ) , .QN( u2_uk_n1594 ) );
  DFF_X1 u2_uk_K_r9_reg_0 (.CK( clk ) , .D( u2_uk_K_r8_0 ) , .Q( u2_uk_K_r9_0 ) );
  DFF_X1 u2_uk_K_r9_reg_1 (.CK( clk ) , .D( u2_uk_K_r8_1 ) , .Q( u2_uk_K_r9_1 ) , .QN( u2_uk_n1632 ) );
  DFF_X1 u2_uk_K_r9_reg_10 (.CK( clk ) , .D( u2_uk_K_r8_10 ) , .Q( u2_uk_K_r9_10 ) );
  DFF_X1 u2_uk_K_r9_reg_11 (.CK( clk ) , .D( u2_uk_K_r8_11 ) , .Q( u2_uk_K_r9_11 ) , .QN( u2_uk_n1637 ) );
  DFF_X1 u2_uk_K_r9_reg_12 (.CK( clk ) , .D( u2_uk_K_r8_12 ) , .Q( u2_uk_K_r9_12 ) );
  DFF_X1 u2_uk_K_r9_reg_13 (.CK( clk ) , .D( u2_uk_K_r8_13 ) , .Q( u2_uk_K_r9_13 ) , .QN( u2_uk_n1639 ) );
  DFF_X1 u2_uk_K_r9_reg_14 (.CK( clk ) , .D( u2_uk_K_r8_14 ) , .Q( u2_uk_K_r9_14 ) , .QN( u2_uk_n1640 ) );
  DFF_X1 u2_uk_K_r9_reg_15 (.CK( clk ) , .D( u2_uk_K_r8_15 ) , .Q( u2_uk_K_r9_15 ) );
  DFF_X1 u2_uk_K_r9_reg_16 (.CK( clk ) , .D( u2_uk_K_r8_16 ) , .Q( u2_uk_K_r9_16 ) , .QN( u2_uk_n1642 ) );
  DFF_X1 u2_uk_K_r9_reg_17 (.CK( clk ) , .D( u2_uk_K_r8_17 ) , .Q( u2_uk_K_r9_17 ) , .QN( u2_uk_n1643 ) );
  DFF_X1 u2_uk_K_r9_reg_18 (.CK( clk ) , .D( u2_uk_K_r8_18 ) , .Q( u2_uk_K_r9_18 ) );
  DFF_X1 u2_uk_K_r9_reg_19 (.CK( clk ) , .D( u2_uk_K_r8_19 ) , .Q( u2_uk_K_r9_19 ) );
  DFF_X1 u2_uk_K_r9_reg_2 (.CK( clk ) , .D( u2_uk_K_r8_2 ) , .Q( u2_uk_K_r9_2 ) );
  DFF_X1 u2_uk_K_r9_reg_20 (.CK( clk ) , .D( u2_uk_K_r8_20 ) , .Q( u2_uk_K_r9_20 ) , .QN( u2_uk_n1646 ) );
  DFF_X1 u2_uk_K_r9_reg_21 (.CK( clk ) , .D( u2_uk_K_r8_21 ) , .Q( u2_uk_K_r9_21 ) , .QN( u2_uk_n1647 ) );
  DFF_X1 u2_uk_K_r9_reg_22 (.CK( clk ) , .D( u2_uk_K_r8_22 ) , .Q( u2_uk_K_r9_22 ) , .QN( u2_uk_n1648 ) );
  DFF_X1 u2_uk_K_r9_reg_23 (.CK( clk ) , .D( u2_uk_K_r8_23 ) , .Q( u2_uk_K_r9_23 ) );
  DFF_X1 u2_uk_K_r9_reg_24 (.CK( clk ) , .D( u2_uk_K_r8_24 ) , .Q( u2_uk_K_r9_24 ) );
  DFF_X1 u2_uk_K_r9_reg_25 (.CK( clk ) , .D( u2_uk_K_r8_25 ) , .Q( u2_uk_K_r9_25 ) );
  DFF_X1 u2_uk_K_r9_reg_26 (.CK( clk ) , .D( u2_uk_K_r8_26 ) , .Q( u2_uk_K_r9_26 ) , .QN( u2_uk_n1652 ) );
  DFF_X1 u2_uk_K_r9_reg_27 (.CK( clk ) , .D( u2_uk_K_r8_27 ) , .Q( u2_uk_K_r9_27 ) );
  DFF_X1 u2_uk_K_r9_reg_28 (.CK( clk ) , .D( u2_uk_K_r8_28 ) , .Q( u2_uk_K_r9_28 ) , .QN( u2_uk_n1653 ) );
  DFF_X1 u2_uk_K_r9_reg_29 (.CK( clk ) , .D( u2_uk_K_r8_29 ) , .Q( u2_uk_K_r9_29 ) , .QN( u2_uk_n1654 ) );
  DFF_X1 u2_uk_K_r9_reg_3 (.CK( clk ) , .D( u2_uk_K_r8_3 ) , .Q( u2_uk_K_r9_3 ) , .QN( u2_uk_n1633 ) );
  DFF_X1 u2_uk_K_r9_reg_30 (.CK( clk ) , .D( u2_uk_K_r8_30 ) , .Q( u2_uk_K_r9_30 ) );
  DFF_X1 u2_uk_K_r9_reg_31 (.CK( clk ) , .D( u2_uk_K_r8_31 ) , .Q( u2_uk_K_r9_31 ) );
  DFF_X1 u2_uk_K_r9_reg_32 (.CK( clk ) , .D( u2_uk_K_r8_32 ) , .Q( u2_uk_K_r9_32 ) , .QN( u2_uk_n1657 ) );
  DFF_X1 u2_uk_K_r9_reg_33 (.CK( clk ) , .D( u2_uk_K_r8_33 ) , .Q( u2_uk_K_r9_33 ) );
  DFF_X1 u2_uk_K_r9_reg_34 (.CK( clk ) , .D( u2_uk_K_r8_34 ) , .Q( u2_uk_K_r9_34 ) , .QN( u2_uk_n1658 ) );
  DFF_X1 u2_uk_K_r9_reg_35 (.CK( clk ) , .D( u2_uk_K_r8_35 ) , .Q( u2_uk_K_r9_35 ) );
  DFF_X1 u2_uk_K_r9_reg_36 (.CK( clk ) , .D( u2_uk_K_r8_36 ) , .Q( u2_uk_K_r9_36 ) , .QN( u2_uk_n1659 ) );
  DFF_X1 u2_uk_K_r9_reg_37 (.CK( clk ) , .D( u2_uk_K_r8_37 ) , .Q( u2_uk_K_r9_37 ) , .QN( u2_uk_n1660 ) );
  DFF_X1 u2_uk_K_r9_reg_38 (.CK( clk ) , .D( u2_uk_K_r8_38 ) , .Q( u2_uk_K_r9_38 ) );
  DFF_X1 u2_uk_K_r9_reg_39 (.CK( clk ) , .D( u2_uk_K_r8_39 ) , .Q( u2_uk_K_r9_39 ) , .QN( u2_uk_n1661 ) );
  DFF_X1 u2_uk_K_r9_reg_4 (.CK( clk ) , .D( u2_uk_K_r8_4 ) , .Q( u2_uk_K_r9_4 ) );
  DFF_X1 u2_uk_K_r9_reg_40 (.CK( clk ) , .D( u2_uk_K_r8_40 ) , .Q( u2_uk_K_r9_40 ) , .QN( u2_uk_n1662 ) );
  DFF_X1 u2_uk_K_r9_reg_41 (.CK( clk ) , .D( u2_uk_K_r8_41 ) , .Q( u2_uk_K_r9_41 ) , .QN( u2_uk_n1663 ) );
  DFF_X1 u2_uk_K_r9_reg_42 (.CK( clk ) , .D( u2_uk_K_r8_42 ) , .Q( u2_uk_K_r9_42 ) , .QN( u2_uk_n1664 ) );
  DFF_X1 u2_uk_K_r9_reg_43 (.CK( clk ) , .D( u2_uk_K_r8_43 ) , .Q( u2_uk_K_r9_43 ) , .QN( u2_uk_n1665 ) );
  DFF_X1 u2_uk_K_r9_reg_44 (.CK( clk ) , .D( u2_uk_K_r8_44 ) , .Q( u2_uk_K_r9_44 ) , .QN( u2_uk_n1666 ) );
  DFF_X1 u2_uk_K_r9_reg_45 (.CK( clk ) , .D( u2_uk_K_r8_45 ) , .Q( u2_uk_K_r9_45 ) );
  DFF_X1 u2_uk_K_r9_reg_46 (.CK( clk ) , .D( u2_uk_K_r8_46 ) , .Q( u2_uk_K_r9_46 ) , .QN( u2_uk_n1668 ) );
  DFF_X1 u2_uk_K_r9_reg_47 (.CK( clk ) , .D( u2_uk_K_r8_47 ) , .Q( u2_uk_K_r9_47 ) , .QN( u2_uk_n1669 ) );
  DFF_X1 u2_uk_K_r9_reg_48 (.CK( clk ) , .D( u2_uk_K_r8_48 ) , .Q( u2_uk_K_r9_48 ) );
  DFF_X1 u2_uk_K_r9_reg_49 (.CK( clk ) , .D( u2_uk_K_r8_49 ) , .Q( u2_uk_K_r9_49 ) );
  DFF_X1 u2_uk_K_r9_reg_5 (.CK( clk ) , .D( u2_uk_K_r8_5 ) , .Q( u2_uk_K_r9_5 ) );
  DFF_X1 u2_uk_K_r9_reg_50 (.CK( clk ) , .D( u2_uk_K_r8_50 ) , .Q( u2_uk_K_r9_50 ) , .QN( u2_uk_n1672 ) );
  DFF_X1 u2_uk_K_r9_reg_51 (.CK( clk ) , .D( u2_uk_K_r8_51 ) , .Q( u2_uk_K_r9_51 ) , .QN( u2_uk_n1673 ) );
  DFF_X1 u2_uk_K_r9_reg_52 (.CK( clk ) , .D( u2_uk_K_r8_52 ) , .Q( u2_uk_K_r9_52 ) , .QN( u2_uk_n1674 ) );
  DFF_X1 u2_uk_K_r9_reg_53 (.CK( clk ) , .D( u2_uk_K_r8_53 ) , .Q( u2_uk_K_r9_53 ) , .QN( u2_uk_n1675 ) );
  DFF_X1 u2_uk_K_r9_reg_54 (.CK( clk ) , .D( u2_uk_K_r8_54 ) , .Q( u2_uk_K_r9_54 ) );
  DFF_X1 u2_uk_K_r9_reg_55 (.CK( clk ) , .D( u2_uk_K_r8_55 ) , .Q( u2_uk_K_r9_55 ) , .QN( u2_uk_n1677 ) );
  DFF_X1 u2_uk_K_r9_reg_6 (.CK( clk ) , .D( u2_uk_K_r8_6 ) , .Q( u2_uk_K_r9_6 ) );
  DFF_X1 u2_uk_K_r9_reg_7 (.CK( clk ) , .D( u2_uk_K_r8_7 ) , .Q( u2_uk_K_r9_7 ) );
  DFF_X1 u2_uk_K_r9_reg_8 (.CK( clk ) , .D( u2_uk_K_r8_8 ) , .Q( u2_uk_K_r9_8 ) , .QN( u2_uk_n1634 ) );
  DFF_X1 u2_uk_K_r9_reg_9 (.CK( clk ) , .D( u2_uk_K_r8_9 ) , .Q( u2_uk_K_r9_9 ) );
  AOI22_X1 u2_uk_U100 (.B2( u2_uk_K_r9_19 ) , .A2( u2_uk_K_r9_25 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n391 ) );
  NAND2_X1 u2_uk_U1000 (.A1( u2_key_r_46 ) , .A2( u2_uk_n100 ) , .ZN( u2_uk_n969 ) );
  OAI21_X1 u2_uk_U1001 (.ZN( u2_K1_17 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1153 ) , .A( u2_uk_n971 ) );
  NAND2_X1 u2_uk_U1002 (.A1( u2_key_r_10 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n971 ) );
  NAND2_X1 u2_uk_U1004 (.A2( decrypt ) , .A1( u2_uk_K_r10_19 ) , .ZN( u2_uk_n520 ) );
  OAI21_X1 u2_uk_U1005 (.ZN( u2_K10_21 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1630 ) , .A( u2_uk_n252 ) );
  NAND2_X1 u2_uk_U1006 (.A1( u2_uk_K_r8_19 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n252 ) );
  OAI21_X1 u2_uk_U1007 (.B1( decrypt ) , .ZN( u2_K1_37 ) , .B2( u2_uk_n1144 ) , .A( u2_uk_n983 ) );
  NAND2_X1 u2_uk_U1008 (.A1( u2_key_r_50 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n983 ) );
  OAI21_X1 u2_uk_U1009 (.ZN( u2_K9_39 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1135 ) , .B2( u2_uk_n1571 ) );
  OAI22_X1 u2_uk_U101 (.A1( decrypt ) , .ZN( u2_K9_5 ) , .B2( u2_uk_n1580 ) , .A2( u2_uk_n1586 ) , .B1( u2_uk_n191 ) );
  NAND2_X1 u2_uk_U1010 (.A1( u2_uk_K_r7_31 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n1135 ) );
  OAI21_X1 u2_uk_U1011 (.ZN( u2_K14_44 ) , .B2( u2_uk_n1777 ) , .B1( u2_uk_n238 ) , .A( u2_uk_n717 ) );
  NAND2_X1 u2_uk_U1012 (.A1( u2_uk_K_r12_15 ) , .A2( u2_uk_n214 ) , .ZN( u2_uk_n717 ) );
  OAI21_X1 u2_uk_U1015 (.ZN( u2_K8_46 ) , .A( u2_uk_n1115 ) , .B2( u2_uk_n1532 ) , .B1( u2_uk_n182 ) );
  NAND2_X1 u2_uk_U1016 (.A1( u2_uk_K_r6_37 ) , .ZN( u2_uk_n1115 ) , .A2( u2_uk_n155 ) );
  OAI21_X1 u2_uk_U1017 (.ZN( u2_K10_13 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1605 ) , .A( u2_uk_n242 ) );
  NAND2_X1 u2_uk_U1018 (.A1( u2_uk_K_r8_48 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n242 ) );
  OAI21_X1 u2_uk_U1019 (.ZN( u2_K12_36 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1698 ) , .A( u2_uk_n472 ) );
  OAI22_X1 u2_uk_U102 (.A1( decrypt ) , .ZN( u2_K7_5 ) , .B2( u2_uk_n1457 ) , .A2( u2_uk_n1474 ) , .B1( u2_uk_n155 ) );
  NAND2_X1 u2_uk_U1020 (.A2( decrypt ) , .A1( u2_uk_K_r10_52 ) , .ZN( u2_uk_n472 ) );
  NAND2_X1 u2_uk_U1022 (.A2( decrypt ) , .A1( u2_uk_K_r4_31 ) , .ZN( u2_uk_n1069 ) );
  OAI21_X1 u2_uk_U1023 (.ZN( u2_K8_28 ) , .A( u2_uk_n1103 ) , .B2( u2_uk_n1532 ) , .B1( u2_uk_n27 ) );
  NAND2_X1 u2_uk_U1024 (.A1( u2_uk_K_r6_51 ) , .ZN( u2_uk_n1103 ) , .A2( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U1027 (.B1( decrypt ) , .ZN( u2_K7_31 ) , .A( u2_uk_n1087 ) , .B2( u2_uk_n1478 ) );
  NAND2_X1 u2_uk_U1028 (.A1( u2_uk_K_r5_16 ) , .ZN( u2_uk_n1087 ) , .A2( u2_uk_n17 ) );
  OAI21_X1 u2_uk_U1029 (.ZN( u2_K12_40 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1699 ) , .A( u2_uk_n501 ) );
  OAI22_X1 u2_uk_U103 (.A1( decrypt ) , .ZN( u2_K5_5 ) , .A2( u2_uk_n1368 ) , .B2( u2_uk_n1392 ) , .B1( u2_uk_n146 ) );
  NAND2_X1 u2_uk_U1030 (.A1( u2_uk_K_r10_49 ) , .A2( u2_uk_n102 ) , .ZN( u2_uk_n501 ) );
  OAI21_X1 u2_uk_U1033 (.ZN( u2_K15_32 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1825 ) , .A( u2_uk_n941 ) );
  NAND2_X1 u2_uk_U1034 (.A2( decrypt ) , .A1( u2_uk_K_r13_36 ) , .ZN( u2_uk_n941 ) );
  OAI21_X1 u2_uk_U1035 (.B1( decrypt ) , .ZN( u2_K7_38 ) , .A( u2_uk_n1092 ) , .B2( u2_uk_n1469 ) );
  NAND2_X1 u2_uk_U1036 (.A2( decrypt ) , .A1( u2_uk_K_r5_8 ) , .ZN( u2_uk_n1092 ) );
  OAI21_X1 u2_uk_U1039 (.B1( decrypt ) , .ZN( u2_K4_38 ) , .A( u2_uk_n1034 ) , .B2( u2_uk_n1353 ) );
  OAI22_X1 u2_uk_U104 (.ZN( u2_K2_5 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1244 ) , .A2( u2_uk_n1247 ) , .A1( u2_uk_n220 ) );
  NAND2_X1 u2_uk_U1040 (.A1( u2_uk_K_r2_50 ) , .A2( u2_uk_n102 ) , .ZN( u2_uk_n1034 ) );
  OAI21_X1 u2_uk_U1041 (.B1( decrypt ) , .ZN( u2_K11_29 ) , .B2( u2_uk_n1634 ) , .A( u2_uk_n366 ) );
  NAND2_X1 u2_uk_U1042 (.A1( u2_uk_K_r9_0 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n366 ) );
  INV_X1 u2_uk_U1043 (.A( u2_key_r_9 ) , .ZN( u2_uk_n1149 ) );
  INV_X1 u2_uk_U1045 (.A( u2_key_r_6 ) , .ZN( u2_uk_n1146 ) );
  INV_X1 u2_uk_U1046 (.A( u2_key_r_54 ) , .ZN( u2_uk_n1185 ) );
  INV_X1 u2_uk_U1048 (.A( u2_key_r_26 ) , .ZN( u2_uk_n1161 ) );
  OAI22_X1 u2_uk_U105 (.B1( decrypt ) , .ZN( u2_K1_5 ) , .A2( u2_uk_n1146 ) , .B2( u2_uk_n1150 ) , .A1( u2_uk_n147 ) );
  INV_X1 u2_uk_U1050 (.A( u2_key_r_47 ) , .ZN( u2_uk_n1179 ) );
  INV_X1 u2_uk_U1051 (.A( u2_key_r_34 ) , .ZN( u2_uk_n1168 ) );
  INV_X1 u2_uk_U1052 (.A( u2_key_r_27 ) , .ZN( u2_uk_n1162 ) );
  INV_X1 u2_uk_U1053 (.A( u2_key_r_24 ) , .ZN( u2_uk_n1159 ) );
  INV_X1 u2_uk_U1054 (.A( u2_key_r_20 ) , .ZN( u2_uk_n1155 ) );
  INV_X1 u2_uk_U1055 (.A( u2_key_r_37 ) , .ZN( u2_uk_n1171 ) );
  INV_X1 u2_uk_U1056 (.A( u2_key_r_52 ) , .ZN( u2_uk_n1183 ) );
  INV_X1 u2_uk_U1057 (.A( u2_key_r_0 ) , .ZN( u2_uk_n1142 ) );
  INV_X1 u2_uk_U1058 (.A( u2_key_r_16 ) , .ZN( u2_uk_n1152 ) );
  INV_X1 u2_uk_U1059 (.A( u2_key_r_13 ) , .ZN( u2_uk_n1150 ) );
  INV_X1 u2_uk_U1060 (.A( u2_key_r_1 ) , .ZN( u2_uk_n1143 ) );
  INV_X1 u2_uk_U1061 (.A( u2_key_r_2 ) , .ZN( u2_uk_n1144 ) );
  INV_X1 u2_uk_U1062 (.A( u2_key_r_19 ) , .ZN( u2_uk_n1154 ) );
  INV_X1 u2_uk_U1063 (.A( u2_key_r_4 ) , .ZN( u2_uk_n1145 ) );
  INV_X1 u2_uk_U1064 (.A( u2_key_r_17 ) , .ZN( u2_uk_n1153 ) );
  INV_X1 u2_uk_U1065 (.A( u2_key_r_53 ) , .ZN( u2_uk_n1184 ) );
  OAI21_X1 u2_uk_U1066 (.ZN( u2_K13_28 ) , .B2( u2_uk_n1753 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n662 ) );
  NAND2_X1 u2_uk_U1067 (.A1( u2_uk_K_r11_21 ) , .A2( u2_uk_n238 ) , .ZN( u2_uk_n662 ) );
  OAI21_X1 u2_uk_U1068 (.ZN( u2_K8_14 ) , .A( u2_uk_n1099 ) , .B2( u2_uk_n1529 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U1069 (.A1( u2_uk_K_r6_34 ) , .ZN( u2_uk_n1099 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U107 (.ZN( u2_K14_41 ) , .A1( u2_uk_n147 ) , .A2( u2_uk_n1776 ) , .B2( u2_uk_n1781 ) , .B1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U1070 (.ZN( u2_K16_14 ) , .B2( u2_uk_n1205 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n951 ) );
  NAND2_X1 u2_uk_U1071 (.A1( u2_uk_K_r14_18 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n951 ) );
  OAI21_X1 u2_uk_U1074 (.ZN( u2_K16_39 ) , .B2( u2_uk_n1201 ) , .B1( u2_uk_n202 ) , .A( u2_uk_n960 ) );
  NAND2_X1 u2_uk_U1075 (.A1( u2_uk_K_r14_15 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n960 ) );
  OAI21_X1 u2_uk_U1076 (.ZN( u2_K8_39 ) , .A( u2_uk_n1109 ) , .B2( u2_uk_n1526 ) , .B1( u2_uk_n202 ) );
  NAND2_X1 u2_uk_U1077 (.A1( u2_uk_K_r6_31 ) , .ZN( u2_uk_n1109 ) , .A2( u2_uk_n155 ) );
  OAI21_X1 u2_uk_U1078 (.ZN( u2_K5_39 ) , .A( u2_uk_n1051 ) , .B2( u2_uk_n1376 ) , .B1( u2_uk_n162 ) );
  NAND2_X1 u2_uk_U1079 (.A1( u2_uk_K_r3_16 ) , .ZN( u2_uk_n1051 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U108 (.A1( decrypt ) , .ZN( u2_K12_41 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1705 ) , .A2( u2_uk_n1714 ) );
  INV_X1 u2_uk_U1080 (.A( u2_key_r_40 ) , .ZN( u2_uk_n1174 ) );
  INV_X1 u2_uk_U1081 (.ZN( u2_K13_10 ) , .A( u2_uk_n524 ) );
  AOI22_X1 u2_uk_U1083 (.B2( u2_uk_K_r0_34 ) , .A2( u2_uk_K_r0_55 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n147 ) , .ZN( u2_uk_n991 ) );
  INV_X1 u2_uk_U1084 (.ZN( u2_K1_11 ) , .A( u2_uk_n967 ) );
  AOI22_X1 u2_uk_U1085 (.B1( decrypt ) , .B2( u2_key_r_32 ) , .A2( u2_key_r_39 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n967 ) );
  INV_X1 u2_uk_U1086 (.ZN( u2_K1_18 ) , .A( u2_uk_n972 ) );
  AOI22_X1 u2_uk_U1087 (.B1( decrypt ) , .A2( u2_key_r_5 ) , .B2( u2_key_r_55 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n972 ) );
  AOI22_X1 u2_uk_U1089 (.B2( u2_uk_K_r6_10 ) , .A2( u2_uk_K_r6_3 ) , .ZN( u2_uk_n1110 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n162 ) );
  AOI22_X1 u2_uk_U1093 (.B2( u2_key_r_35 ) , .A2( u2_key_r_42 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) , .ZN( u2_uk_n985 ) );
  INV_X1 u2_uk_U1094 (.ZN( u2_K11_8 ) , .A( u2_uk_n407 ) );
  AOI22_X1 u2_uk_U1095 (.B2( u2_uk_K_r9_12 ) , .A2( u2_uk_K_r9_18 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n230 ) , .ZN( u2_uk_n407 ) );
  AOI22_X1 u2_uk_U1097 (.B1( decrypt ) , .B2( u2_uk_K_r9_25 ) , .A2( u2_uk_K_r9_6 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n313 ) );
  AOI22_X1 u2_uk_U1099 (.B2( u2_uk_K_r6_3 ) , .A2( u2_uk_K_r6_53 ) , .ZN( u2_uk_n1098 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U110 (.B1( decrypt ) , .ZN( u2_K16_47 ) , .B2( u2_uk_n1188 ) , .A2( u2_uk_n1192 ) , .A1( u2_uk_n207 ) );
  INV_X1 u2_uk_U1100 (.ZN( u2_K1_20 ) , .A( u2_uk_n973 ) );
  AOI22_X1 u2_uk_U1101 (.B2( u2_key_r_48 ) , .A2( u2_key_r_55 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n63 ) , .ZN( u2_uk_n973 ) );
  AOI22_X1 u2_uk_U1103 (.B2( u2_uk_K_r0_15 ) , .A2( u2_uk_K_r0_36 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n155 ) , .ZN( u2_uk_n999 ) );
  AOI22_X1 u2_uk_U1105 (.B1( decrypt ) , .A2( u2_uk_K_r2_4 ) , .B2( u2_uk_K_r2_41 ) , .ZN( u2_uk_n1035 ) , .A1( u2_uk_n230 ) );
  AOI22_X1 u2_uk_U1107 (.B2( u2_uk_K_r10_32 ) , .A2( u2_uk_K_r10_41 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n454 ) );
  AOI22_X1 u2_uk_U1109 (.B2( u2_uk_K_r0_13 ) , .A2( u2_uk_K_r0_34 ) , .ZN( u2_uk_n1004 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U111 (.A1( decrypt ) , .ZN( u2_K13_47 ) , .B2( u2_uk_n1752 ) , .A2( u2_uk_n1762 ) , .B1( u2_uk_n202 ) );
  AOI22_X1 u2_uk_U1111 (.B1( decrypt ) , .B2( u2_uk_K_r10_23 ) , .A2( u2_uk_K_r10_28 ) , .A1( u2_uk_n220 ) , .ZN( u2_uk_n467 ) );
  AOI22_X1 u2_uk_U1115 (.B1( decrypt ) , .B2( u2_uk_K_r3_24 ) , .A2( u2_uk_K_r3_47 ) , .ZN( u2_uk_n1043 ) , .A1( u2_uk_n155 ) );
  AOI22_X1 u2_uk_U1117 (.B2( u2_uk_K_r5_26 ) , .A2( u2_uk_K_r5_48 ) , .ZN( u2_uk_n1076 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n145 ) );
  INV_X1 u2_uk_U1118 (.ZN( u2_K1_32 ) , .A( u2_uk_n980 ) );
  AOI22_X1 u2_uk_U1119 (.B2( u2_key_r_22 ) , .A2( u2_key_r_29 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n980 ) );
  OAI22_X1 u2_uk_U112 (.A1( decrypt ) , .ZN( u2_K12_47 ) , .B2( u2_uk_n1679 ) , .A2( u2_uk_n1706 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U1121 (.B2( u2_uk_K_r5_0 ) , .A2( u2_uk_K_r5_51 ) , .ZN( u2_uk_n1088 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n231 ) );
  AOI22_X1 u2_uk_U1123 (.B1( decrypt ) , .B2( u2_uk_K_r2_13 ) , .A2( u2_uk_K_r2_33 ) , .ZN( u2_uk_n1024 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U1127 (.A1( decrypt ) , .B2( u2_uk_K_r3_29 ) , .A2( u2_uk_K_r3_38 ) , .ZN( u2_uk_n1049 ) , .B1( u2_uk_n163 ) );
  INV_X1 u2_uk_U1128 (.ZN( u2_K6_4 ) , .A( u2_uk_n1071 ) );
  AOI22_X1 u2_uk_U1129 (.B2( u2_uk_K_r4_41 ) , .A2( u2_uk_K_r4_47 ) , .ZN( u2_uk_n1071 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n60 ) );
  AOI22_X1 u2_uk_U1131 (.B2( u2_uk_K_r2_26 ) , .A2( u2_uk_K_r2_6 ) , .ZN( u2_uk_n1020 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n60 ) );
  AOI22_X1 u2_uk_U1133 (.A1( decrypt ) , .B2( u2_uk_K_r8_17 ) , .A2( u2_uk_K_r8_39 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n240 ) );
  INV_X1 u2_uk_U1134 (.ZN( u2_K13_12 ) , .A( u2_uk_n551 ) );
  AOI22_X1 u2_uk_U1135 (.A1( decrypt ) , .B2( u2_uk_K_r11_34 ) , .A2( u2_uk_K_r11_54 ) , .B1( u2_uk_n238 ) , .ZN( u2_uk_n551 ) );
  INV_X1 u2_uk_U1136 (.ZN( u2_K8_15 ) , .A( u2_uk_n1100 ) );
  AOI22_X1 u2_uk_U1137 (.A1( decrypt ) , .B2( u2_uk_K_r6_10 ) , .A2( u2_uk_K_r6_17 ) , .ZN( u2_uk_n1100 ) , .B1( u2_uk_n188 ) );
  AOI22_X1 u2_uk_U1138 (.A1( decrypt ) , .B2( u2_uk_K_r6_21 ) , .A2( u2_uk_K_r6_28 ) , .ZN( u2_uk_n1113 ) , .B1( u2_uk_n238 ) );
  AOI22_X1 u2_uk_U114 (.B2( u2_uk_K_r9_15 ) , .A2( u2_uk_K_r9_23 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n223 ) , .ZN( u2_uk_n386 ) );
  OAI21_X1 u2_uk_U1140 (.ZN( u2_K16_2 ) , .B2( u2_uk_n1190 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n956 ) );
  NAND2_X1 u2_uk_U1141 (.A2( decrypt ) , .A1( u2_uk_K_r14_11 ) , .ZN( u2_uk_n956 ) );
  AOI22_X1 u2_uk_U1142 (.B1( decrypt ) , .A2( u2_uk_K_r13_2 ) , .B2( u2_uk_K_r13_23 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n944 ) );
  INV_X1 u2_uk_U1143 (.ZN( u2_K15_43 ) , .A( u2_uk_n944 ) );
  AOI22_X1 u2_uk_U1144 (.B1( decrypt ) , .B2( u2_uk_K_r10_39 ) , .A2( u2_uk_K_r10_48 ) , .A1( u2_uk_n209 ) , .ZN( u2_uk_n421 ) );
  AOI22_X1 u2_uk_U1147 (.B2( u2_uk_K_r11_26 ) , .A2( u2_uk_K_r11_6 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n524 ) );
  AOI22_X1 u2_uk_U1148 (.A1( decrypt ) , .B2( u2_uk_K_r11_26 ) , .A2( u2_uk_K_r11_46 ) , .B1( u2_uk_n209 ) , .ZN( u2_uk_n665 ) );
  INV_X1 u2_uk_U1149 (.ZN( u2_K13_6 ) , .A( u2_uk_n681 ) );
  OAI22_X1 u2_uk_U1150 (.ZN( u2_K1_23 ) , .B2( u2_uk_n1167 ) , .A2( u2_uk_n1174 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U1151 (.A( u2_key_r_33 ) , .ZN( u2_uk_n1167 ) );
  AOI22_X1 u2_uk_U1152 (.B1( decrypt ) , .B2( u2_uk_K_r7_20 ) , .A2( u2_uk_K_r7_27 ) , .ZN( u2_uk_n1130 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U1156 (.B1( decrypt ) , .B2( u2_uk_K_r2_26 ) , .A2( u2_uk_K_r2_46 ) , .ZN( u2_uk_n1031 ) , .A1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U116 (.ZN( u2_K8_47 ) , .B2( u2_uk_n1531 ) , .A2( u2_uk_n1537 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n223 ) );
  OAI21_X1 u2_uk_U118 (.ZN( u2_K6_47 ) , .A( u2_uk_n1070 ) , .B2( u2_uk_n1419 ) , .B1( u2_uk_n60 ) );
  NAND2_X1 u2_uk_U119 (.A2( decrypt ) , .A1( u2_uk_K_r4_23 ) , .ZN( u2_uk_n1070 ) );
  OAI22_X1 u2_uk_U120 (.B1( decrypt ) , .ZN( u2_K5_47 ) , .B2( u2_uk_n1365 ) , .A2( u2_uk_n1389 ) , .A1( u2_uk_n213 ) );
  OAI21_X1 u2_uk_U122 (.B1( decrypt ) , .ZN( u2_K2_47 ) , .A( u2_uk_n1003 ) , .B2( u2_uk_n1241 ) );
  NAND2_X1 u2_uk_U123 (.A2( decrypt ) , .A1( u2_uk_K_r0_52 ) , .ZN( u2_uk_n1003 ) );
  OAI22_X1 u2_uk_U124 (.A1( decrypt ) , .ZN( u2_K1_15 ) , .B2( u2_uk_n1161 ) , .A2( u2_uk_n1167 ) , .B1( u2_uk_n209 ) );
  OAI21_X1 u2_uk_U126 (.ZN( u2_K5_15 ) , .A( u2_uk_n1042 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1379 ) );
  NAND2_X1 u2_uk_U127 (.A2( decrypt ) , .A1( u2_uk_K_r3_34 ) , .ZN( u2_uk_n1042 ) );
  INV_X1 u2_uk_U128 (.ZN( u2_K13_15 ) , .A( u2_uk_n586 ) );
  AOI22_X1 u2_uk_U129 (.B1( decrypt ) , .B2( u2_uk_K_r11_11 ) , .A2( u2_uk_K_r11_48 ) , .A1( u2_uk_n141 ) , .ZN( u2_uk_n586 ) );
  INV_X1 u2_uk_U131 (.ZN( u2_K12_15 ) , .A( u2_uk_n409 ) );
  AOI22_X1 u2_uk_U132 (.B2( u2_uk_K_r10_25 ) , .A2( u2_uk_K_r10_34 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n222 ) , .ZN( u2_uk_n409 ) );
  OAI22_X1 u2_uk_U133 (.B1( decrypt ) , .ZN( u2_K3_15 ) , .A2( u2_uk_n1282 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1317 ) );
  INV_X1 u2_uk_U134 (.ZN( u2_K13_19 ) , .A( u2_uk_n601 ) );
  AOI22_X1 u2_uk_U135 (.B2( u2_uk_K_r11_19 ) , .A2( u2_uk_K_r11_39 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n601 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U136 (.ZN( u2_K11_15 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1646 ) , .A2( u2_uk_n1661 ) , .B1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U137 (.ZN( u2_K6_19 ) , .A( u2_uk_n1061 ) , .B2( u2_uk_n1414 ) , .B1( u2_uk_n63 ) );
  NAND2_X1 u2_uk_U138 (.A2( decrypt ) , .A1( u2_uk_K_r4_48 ) , .ZN( u2_uk_n1061 ) );
  OAI21_X1 u2_uk_U139 (.ZN( u2_K2_15 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1261 ) , .A( u2_uk_n994 ) );
  NAND2_X1 u2_uk_U140 (.A2( decrypt ) , .A1( u2_uk_K_r0_19 ) , .ZN( u2_uk_n994 ) );
  OAI22_X1 u2_uk_U141 (.B1( decrypt ) , .ZN( u2_K1_19 ) , .B2( u2_uk_n1145 ) , .A2( u2_uk_n1185 ) , .A1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U142 (.ZN( u2_K16_15 ) , .B2( u2_uk_n1206 ) , .A2( u2_uk_n1213 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U143 (.A1( decrypt ) , .ZN( u2_K10_15 ) , .A2( u2_uk_n1592 ) , .B2( u2_uk_n1629 ) , .B1( u2_uk_n182 ) );
  OAI21_X1 u2_uk_U144 (.ZN( u2_K15_15 ) , .B2( u2_uk_n1843 ) , .B1( u2_uk_n188 ) , .A( u2_uk_n937 ) );
  NAND2_X1 u2_uk_U145 (.A1( u2_uk_K_r13_19 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n937 ) );
  OAI22_X1 u2_uk_U146 (.ZN( u2_K14_15 ) , .A2( u2_uk_n1773 ) , .B2( u2_uk_n1811 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U147 (.ZN( u2_K14_19 ) , .A( u2_uk_n685 ) );
  AOI22_X1 u2_uk_U148 (.B2( u2_uk_K_r12_25 ) , .A2( u2_uk_K_r12_33 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n685 ) );
  AOI22_X1 u2_uk_U152 (.B1( u2_uk_K_r7_13 ) , .A2( u2_uk_K_r7_20 ) , .B2( u2_uk_n10 ) , .ZN( u2_uk_n1124 ) , .A1( u2_uk_n162 ) );
  OAI21_X1 u2_uk_U154 (.ZN( u2_K3_19 ) , .A( u2_uk_n1007 ) , .B2( u2_uk_n1294 ) , .B1( u2_uk_n83 ) );
  NAND2_X1 u2_uk_U155 (.A2( decrypt ) , .A1( u2_uk_K_r1_33 ) , .ZN( u2_uk_n1007 ) );
  AOI22_X1 u2_uk_U157 (.B2( u2_uk_K_r0_11 ) , .A2( u2_uk_K_r0_47 ) , .A1( u2_uk_n128 ) , .B1( u2_uk_n231 ) , .ZN( u2_uk_n995 ) );
  OAI22_X1 u2_uk_U158 (.ZN( u2_K16_19 ) , .B2( u2_uk_n1190 ) , .A2( u2_uk_n1228 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U159 (.ZN( u2_K8_19 ) , .B2( u2_uk_n1508 ) , .A2( u2_uk_n1515 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U160 (.ZN( u2_K10_19 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1603 ) , .A2( u2_uk_n1613 ) , .B1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U161 (.ZN( u2_K5_30 ) , .B2( u2_uk_n1378 ) , .A2( u2_uk_n1395 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U162 (.ZN( u2_K2_30 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1230 ) , .A2( u2_uk_n1259 ) , .A1( u2_uk_n162 ) );
  AOI22_X1 u2_uk_U165 (.A1( decrypt ) , .B2( u2_uk_K_r10_23 ) , .A2( u2_uk_K_r10_42 ) , .B1( u2_uk_n191 ) , .ZN( u2_uk_n456 ) );
  OAI22_X1 u2_uk_U166 (.A1( decrypt ) , .ZN( u2_K10_30 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1598 ) , .A2( u2_uk_n1626 ) );
  OAI22_X1 u2_uk_U167 (.A1( decrypt ) , .ZN( u2_K12_24 ) , .B1( u2_uk_n155 ) , .B2( u2_uk_n1686 ) , .A2( u2_uk_n1715 ) );
  OAI21_X1 u2_uk_U168 (.ZN( u2_K1_14 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1160 ) , .A( u2_uk_n970 ) );
  NAND2_X1 u2_uk_U169 (.A2( decrypt ) , .A1( u2_key_r_18 ) , .ZN( u2_uk_n970 ) );
  INV_X1 u2_uk_U170 (.A( u2_key_r_25 ) , .ZN( u2_uk_n1160 ) );
  OAI21_X1 u2_uk_U171 (.ZN( u2_K8_30 ) , .A( u2_uk_n1106 ) , .B2( u2_uk_n1525 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U172 (.A1( u2_uk_K_r6_29 ) , .ZN( u2_uk_n1106 ) , .A2( u2_uk_n191 ) );
  OAI21_X1 u2_uk_U173 (.ZN( u2_K16_30 ) , .B2( u2_uk_n1226 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n957 ) );
  NAND2_X1 u2_uk_U174 (.A1( u2_uk_K_r14_45 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n957 ) );
  OAI22_X1 u2_uk_U175 (.A1( decrypt ) , .ZN( u2_K13_14 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1726 ) , .A2( u2_uk_n1750 ) );
  AOI22_X1 u2_uk_U178 (.A1( decrypt ) , .B2( u2_uk_K_r9_12 ) , .A2( u2_uk_K_r9_6 ) , .B1( u2_uk_n188 ) , .ZN( u2_uk_n319 ) );
  OAI21_X1 u2_uk_U179 (.ZN( u2_K10_24 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1599 ) , .A( u2_uk_n277 ) );
  NAND2_X1 u2_uk_U180 (.A1( u2_uk_K_r8_40 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n277 ) );
  OAI21_X1 u2_uk_U181 (.ZN( u2_K9_14 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1121 ) , .B2( u2_uk_n1574 ) );
  NAND2_X1 u2_uk_U182 (.A2( decrypt ) , .A1( u2_uk_K_r7_34 ) , .ZN( u2_uk_n1121 ) );
  OAI22_X1 u2_uk_U183 (.A1( decrypt ) , .ZN( u2_K6_14 ) , .A2( u2_uk_n1410 ) , .B2( u2_uk_n1416 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U185 (.B2( u2_uk_K_r0_11 ) , .A2( u2_uk_K_r0_32 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n993 ) );
  OAI22_X1 u2_uk_U186 (.A1( decrypt ) , .ZN( u2_K1_24 ) , .B2( u2_uk_n1150 ) , .A2( u2_uk_n1155 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U187 (.ZN( u2_K11_30 ) , .A( u2_uk_n369 ) );
  AOI22_X1 u2_uk_U188 (.B2( u2_uk_K_r9_1 ) , .A2( u2_uk_K_r9_9 ) , .B1( u2_uk_n110 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n369 ) );
  OAI22_X1 u2_uk_U189 (.ZN( u2_K10_14 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1600 ) , .A2( u2_uk_n1631 ) , .B1( u2_uk_n238 ) );
  OAI21_X1 u2_uk_U192 (.ZN( u2_K14_24 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1782 ) , .A( u2_uk_n686 ) );
  NAND2_X1 u2_uk_U193 (.A1( u2_uk_K_r12_41 ) , .A2( u2_uk_n17 ) , .ZN( u2_uk_n686 ) );
  AOI22_X1 u2_uk_U195 (.B2( u2_uk_K_r5_18 ) , .A2( u2_uk_K_r5_40 ) , .ZN( u2_uk_n1083 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U196 (.ZN( u2_K4_24 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1322 ) , .A2( u2_uk_n1363 ) , .B1( u2_uk_n142 ) );
  AOI22_X1 u2_uk_U198 (.B2( u2_uk_K_r1_17 ) , .A2( u2_uk_K_r1_41 ) , .ZN( u2_uk_n1008 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U200 (.ZN( u2_K1_30 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1183 ) , .A( u2_uk_n979 ) );
  NAND2_X1 u2_uk_U201 (.A2( decrypt ) , .A1( u2_key_r_45 ) , .ZN( u2_uk_n979 ) );
  OAI21_X1 u2_uk_U202 (.ZN( u2_K9_30 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1131 ) , .B2( u2_uk_n1570 ) );
  NAND2_X1 u2_uk_U203 (.A2( decrypt ) , .A1( u2_uk_K_r7_29 ) , .ZN( u2_uk_n1131 ) );
  INV_X1 u2_uk_U206 (.ZN( u2_K15_30 ) , .A( u2_uk_n940 ) );
  AOI22_X1 u2_uk_U207 (.B2( u2_uk_K_r13_0 ) , .A2( u2_uk_K_r13_38 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n940 ) );
  OAI22_X1 u2_uk_U213 (.A1( decrypt ) , .ZN( u2_K16_31 ) , .A2( u2_uk_n1192 ) , .B2( u2_uk_n1195 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U214 (.A1( decrypt ) , .ZN( u2_K8_31 ) , .B2( u2_uk_n1499 ) , .A2( u2_uk_n1537 ) , .B1( u2_uk_n208 ) );
  OAI21_X1 u2_uk_U215 (.ZN( u2_K12_31 ) , .B2( u2_uk_n1685 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n460 ) );
  NAND2_X1 u2_uk_U216 (.A1( u2_uk_K_r10_44 ) , .A2( u2_uk_n217 ) , .ZN( u2_uk_n460 ) );
  AOI22_X1 u2_uk_U218 (.B1( decrypt ) , .B2( u2_uk_K_r9_22 ) , .A2( u2_uk_K_r9_30 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n373 ) );
  OAI22_X1 u2_uk_U219 (.ZN( u2_K2_31 ) , .B2( u2_uk_n1230 ) , .A2( u2_uk_n1245 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U220 (.ZN( u2_K11_39 ) , .A( u2_uk_n379 ) );
  AOI22_X1 u2_uk_U221 (.B1( decrypt ) , .B2( u2_uk_K_r9_30 ) , .A2( u2_uk_K_r9_7 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n379 ) );
  AOI22_X1 u2_uk_U223 (.B2( u2_uk_K_r8_44 ) , .A2( u2_uk_K_r8_52 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n305 ) );
  OAI22_X1 u2_uk_U224 (.B1( decrypt ) , .ZN( u2_K13_31 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1742 ) , .A2( u2_uk_n1760 ) );
  OAI22_X1 u2_uk_U227 (.ZN( u2_K6_31 ) , .B2( u2_uk_n1425 ) , .A2( u2_uk_n1430 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U228 (.ZN( u2_K3_31 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1303 ) , .A2( u2_uk_n1309 ) , .A1( u2_uk_n213 ) );
  OAI21_X1 u2_uk_U229 (.B1( decrypt ) , .ZN( u2_K5_31 ) , .A( u2_uk_n1047 ) , .B2( u2_uk_n1371 ) );
  NAND2_X1 u2_uk_U230 (.A2( decrypt ) , .A1( u2_uk_K_r3_44 ) , .ZN( u2_uk_n1047 ) );
  OAI22_X1 u2_uk_U231 (.B1( decrypt ) , .ZN( u2_K15_31 ) , .B2( u2_uk_n1813 ) , .A2( u2_uk_n1830 ) , .A1( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U232 (.ZN( u2_K1_39 ) , .B2( u2_uk_n1157 ) , .B1( u2_uk_n63 ) , .A( u2_uk_n984 ) );
  NAND2_X1 u2_uk_U233 (.A2( decrypt ) , .A1( u2_key_r_15 ) , .ZN( u2_uk_n984 ) );
  INV_X1 u2_uk_U234 (.A( u2_key_r_22 ) , .ZN( u2_uk_n1157 ) );
  OAI22_X1 u2_uk_U236 (.ZN( u2_K9_31 ) , .B2( u2_uk_n1542 ) , .A2( u2_uk_n1583 ) , .A1( u2_uk_n230 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U237 (.A1( decrypt ) , .ZN( u2_K15_39 ) , .A2( u2_uk_n1818 ) , .B2( u2_uk_n1836 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U238 (.A1( decrypt ) , .ZN( u2_K14_39 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1802 ) , .A2( u2_uk_n1806 ) );
  OAI22_X1 u2_uk_U239 (.ZN( u2_K13_39 ) , .B1( u2_uk_n161 ) , .B2( u2_uk_n1725 ) , .A2( u2_uk_n1744 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U240 (.ZN( u2_K12_39 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1690 ) , .A( u2_uk_n496 ) );
  NAND2_X1 u2_uk_U241 (.A1( u2_uk_K_r10_16 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n496 ) );
  OAI22_X1 u2_uk_U242 (.ZN( u2_K16_48 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1200 ) , .A2( u2_uk_n1208 ) , .A1( u2_uk_n213 ) );
  OAI21_X1 u2_uk_U243 (.B1( decrypt ) , .ZN( u2_K16_44 ) , .B2( u2_uk_n1216 ) , .A( u2_uk_n964 ) );
  NAND2_X1 u2_uk_U244 (.A2( decrypt ) , .A1( u2_uk_K_r14_43 ) , .ZN( u2_uk_n964 ) );
  OAI22_X1 u2_uk_U245 (.B1( decrypt ) , .ZN( u2_K5_44 ) , .B2( u2_uk_n1389 ) , .A2( u2_uk_n1395 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U246 (.B1( decrypt ) , .ZN( u2_K5_48 ) , .B2( u2_uk_n1377 ) , .A2( u2_uk_n1384 ) , .A1( u2_uk_n213 ) );
  INV_X1 u2_uk_U247 (.ZN( u2_K1_48 ) , .A( u2_uk_n989 ) );
  AOI22_X1 u2_uk_U248 (.B2( u2_key_r_21 ) , .A2( u2_key_r_28 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n217 ) , .ZN( u2_uk_n989 ) );
  OAI22_X1 u2_uk_U249 (.ZN( u2_K15_44 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1836 ) , .A2( u2_uk_n1854 ) , .A1( u2_uk_n230 ) );
  NAND2_X1 u2_uk_U251 (.A2( decrypt ) , .A1( u2_uk_K_r13_35 ) , .ZN( u2_uk_n945 ) );
  OAI22_X1 u2_uk_U252 (.ZN( u2_K14_48 ) , .B2( u2_uk_n1768 ) , .A2( u2_uk_n1806 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U253 (.B1( decrypt ) , .ZN( u2_K13_44 ) , .B2( u2_uk_n1724 ) , .A2( u2_uk_n1739 ) , .A1( u2_uk_n220 ) );
  OAI21_X1 u2_uk_U254 (.ZN( u2_K13_48 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1755 ) , .A( u2_uk_n677 ) );
  NAND2_X1 u2_uk_U255 (.A2( decrypt ) , .A1( u2_uk_K_r11_8 ) , .ZN( u2_uk_n677 ) );
  AOI22_X1 u2_uk_U257 (.B1( decrypt ) , .B2( u2_uk_K_r10_37 ) , .A2( u2_uk_K_r10_42 ) , .A1( u2_uk_n230 ) , .ZN( u2_uk_n504 ) );
  OAI22_X1 u2_uk_U258 (.ZN( u2_K12_48 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1691 ) , .A2( u2_uk_n1700 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U259 (.ZN( u2_K11_44 ) , .A1( u2_uk_n142 ) , .B2( u2_uk_n1653 ) , .A2( u2_uk_n1673 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U260 (.B1( decrypt ) , .ZN( u2_K10_44 ) , .B2( u2_uk_n1597 ) , .A2( u2_uk_n1617 ) , .A1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U261 (.ZN( u2_K10_48 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1610 ) , .A2( u2_uk_n1626 ) , .B1( u2_uk_n83 ) );
  AOI22_X1 u2_uk_U263 (.A1( decrypt ) , .B2( u2_uk_K_r7_16 ) , .A2( u2_uk_K_r7_9 ) , .ZN( u2_uk_n1140 ) , .B1( u2_uk_n231 ) );
  OAI21_X1 u2_uk_U264 (.ZN( u2_K8_44 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1114 ) , .B2( u2_uk_n1538 ) );
  NAND2_X1 u2_uk_U265 (.A1( u2_uk_K_r6_0 ) , .ZN( u2_uk_n1114 ) , .A2( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U266 (.ZN( u2_K8_48 ) , .A2( u2_uk_n1504 ) , .B2( u2_uk_n1511 ) , .B1( u2_uk_n217 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U268 (.A1( decrypt ) , .ZN( u2_K7_48 ) , .B2( u2_uk_n1471 ) , .A2( u2_uk_n1491 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U271 (.ZN( u2_K4_44 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1320 ) , .A2( u2_uk_n1337 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U274 (.A1( decrypt ) , .ZN( u2_K3_48 ) , .B2( u2_uk_n1277 ) , .A2( u2_uk_n1312 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U275 (.A1( decrypt ) , .ZN( u2_K2_44 ) , .B2( u2_uk_n1251 ) , .A2( u2_uk_n1273 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U276 (.B1( decrypt ) , .ZN( u2_K16_6 ) , .B2( u2_uk_n1214 ) , .A2( u2_uk_n1219 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U278 (.B1( decrypt ) , .ZN( u2_K14_6 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1773 ) , .B2( u2_uk_n1780 ) );
  OAI22_X1 u2_uk_U279 (.B1( decrypt ) , .ZN( u2_K10_6 ) , .A1( u2_uk_n147 ) , .A2( u2_uk_n1591 ) , .B2( u2_uk_n1619 ) );
  OAI22_X1 u2_uk_U280 (.ZN( u2_K6_6 ) , .B2( u2_uk_n1444 ) , .A2( u2_uk_n1448 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) );
  OAI21_X1 u2_uk_U281 (.ZN( u2_K6_8 ) , .A( u2_uk_n1073 ) , .B2( u2_uk_n1416 ) , .B1( u2_uk_n31 ) );
  NAND2_X1 u2_uk_U282 (.A2( decrypt ) , .A1( u2_uk_K_r4_18 ) , .ZN( u2_uk_n1073 ) );
  OAI22_X1 u2_uk_U284 (.ZN( u2_K1_8 ) , .A2( u2_uk_n1146 ) , .B2( u2_uk_n1159 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  AOI22_X1 u2_uk_U286 (.B2( u2_uk_K_r13_13 ) , .A2( u2_uk_K_r13_17 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n141 ) , .ZN( u2_uk_n946 ) );
  OAI22_X1 u2_uk_U287 (.B1( decrypt ) , .ZN( u2_K12_8 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1701 ) , .A2( u2_uk_n1722 ) );
  OAI22_X1 u2_uk_U288 (.B1( decrypt ) , .ZN( u2_K8_8 ) , .B2( u2_uk_n1528 ) , .A2( u2_uk_n1534 ) , .A1( u2_uk_n203 ) );
  AOI22_X1 u2_uk_U290 (.A1( decrypt ) , .B2( u2_uk_K_r5_26 ) , .A2( u2_uk_K_r5_4 ) , .ZN( u2_uk_n1096 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U291 (.A1( decrypt ) , .ZN( u2_K5_8 ) , .B2( u2_uk_n1385 ) , .A2( u2_uk_n1407 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U293 (.A1( decrypt ) , .B2( u2_uk_K_r2_41 ) , .A2( u2_uk_K_r2_46 ) , .ZN( u2_uk_n1040 ) , .B1( u2_uk_n188 ) );
  OAI21_X1 u2_uk_U295 (.ZN( u2_K2_8 ) , .A( u2_uk_n1005 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1240 ) );
  NAND2_X1 u2_uk_U296 (.A1( u2_uk_K_r0_17 ) , .ZN( u2_uk_n1005 ) , .A2( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U297 (.A1( decrypt ) , .ZN( u2_K7_26 ) , .B2( u2_uk_n1470 ) , .A2( u2_uk_n1490 ) , .B1( u2_uk_n209 ) );
  INV_X1 u2_uk_U298 (.ZN( u2_K1_26 ) , .A( u2_uk_n976 ) );
  AOI22_X1 u2_uk_U299 (.B2( u2_key_r_31 ) , .A2( u2_key_r_51 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n976 ) );
  OAI22_X1 u2_uk_U300 (.B1( decrypt ) , .ZN( u2_K16_8 ) , .A2( u2_uk_n1191 ) , .B2( u2_uk_n1204 ) , .A1( u2_uk_n230 ) );
  AOI22_X1 u2_uk_U302 (.A1( decrypt ) , .B2( u2_uk_K_r7_15 ) , .A2( u2_uk_K_r7_8 ) , .ZN( u2_uk_n1128 ) , .B1( u2_uk_n238 ) );
  AOI22_X1 u2_uk_U304 (.B1( decrypt ) , .B2( u2_uk_K_r2_16 ) , .A2( u2_uk_K_r2_7 ) , .ZN( u2_uk_n1028 ) , .A1( u2_uk_n163 ) );
  AOI22_X1 u2_uk_U306 (.B1( decrypt ) , .B2( u2_uk_K_r13_38 ) , .A2( u2_uk_K_r13_44 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n939 ) );
  OAI21_X1 u2_uk_U309 (.ZN( u2_K11_26 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1665 ) , .A( u2_uk_n363 ) );
  NAND2_X1 u2_uk_U310 (.A2( decrypt ) , .A1( u2_uk_K_r9_35 ) , .ZN( u2_uk_n363 ) );
  OAI21_X1 u2_uk_U311 (.B1( decrypt ) , .ZN( u2_K13_26 ) , .B2( u2_uk_n1735 ) , .A( u2_uk_n656 ) );
  NAND2_X1 u2_uk_U312 (.A1( u2_uk_K_r11_7 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n656 ) );
  OAI22_X1 u2_uk_U313 (.B1( decrypt ) , .ZN( u2_K5_26 ) , .A2( u2_uk_n1366 ) , .B2( u2_uk_n1376 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U314 (.ZN( u2_K2_26 ) , .B2( u2_uk_n1259 ) , .A2( u2_uk_n1265 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U315 (.A1( decrypt ) , .ZN( u2_K16_26 ) , .B2( u2_uk_n1211 ) , .A2( u2_uk_n1225 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U316 (.ZN( u2_K14_26 ) , .B2( u2_uk_n1792 ) , .A2( u2_uk_n1809 ) , .A1( u2_uk_n191 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U317 (.A1( decrypt ) , .ZN( u2_K12_26 ) , .B1( u2_uk_n146 ) , .A2( u2_uk_n1680 ) , .B2( u2_uk_n1690 ) );
  OAI22_X1 u2_uk_U318 (.B1( decrypt ) , .ZN( u2_K10_26 ) , .B2( u2_uk_n1609 ) , .A2( u2_uk_n1625 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U319 (.A1( decrypt ) , .ZN( u2_K8_26 ) , .A2( u2_uk_n1503 ) , .B2( u2_uk_n1510 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U320 (.ZN( u2_K3_26 ) , .B2( u2_uk_n1299 ) , .A2( u2_uk_n1315 ) , .B1( u2_uk_n141 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U321 (.ZN( u2_K5_46 ) , .B2( u2_uk_n1364 ) , .A2( u2_uk_n1401 ) , .B1( u2_uk_n146 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U322 (.ZN( u2_K15_46 ) , .B1( u2_uk_n17 ) , .A2( u2_uk_n1818 ) , .B2( u2_uk_n1845 ) , .A1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U323 (.B1( decrypt ) , .ZN( u2_K13_46 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1733 ) , .A2( u2_uk_n1745 ) );
  OAI22_X1 u2_uk_U324 (.B1( decrypt ) , .ZN( u2_K12_46 ) , .B2( u2_uk_n1678 ) , .A2( u2_uk_n1718 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U325 (.ZN( u2_K4_46 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1330 ) , .A2( u2_uk_n1344 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U328 (.A1( decrypt ) , .ZN( u2_K2_46 ) , .A2( u2_uk_n1236 ) , .B2( u2_uk_n1263 ) , .B1( u2_uk_n163 ) );
  OAI21_X1 u2_uk_U329 (.B1( decrypt ) , .ZN( u2_K1_46 ) , .B2( u2_uk_n1143 ) , .A( u2_uk_n988 ) );
  NAND2_X1 u2_uk_U330 (.A1( u2_key_r_49 ) , .A2( u2_uk_n94 ) , .ZN( u2_uk_n988 ) );
  OAI22_X1 u2_uk_U331 (.ZN( u2_K15_4 ) , .B2( u2_uk_n1820 ) , .A2( u2_uk_n1850 ) , .B1( u2_uk_n208 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U332 (.ZN( u2_K14_4 ) , .B2( u2_uk_n1786 ) , .A2( u2_uk_n1794 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U333 (.A1( decrypt ) , .ZN( u2_K11_4 ) , .B2( u2_uk_n1663 ) , .A2( u2_uk_n1669 ) , .B1( u2_uk_n214 ) );
  INV_X1 u2_uk_U334 (.ZN( u2_K11_46 ) , .A( u2_uk_n385 ) );
  AOI22_X1 u2_uk_U335 (.A1( decrypt ) , .B2( u2_uk_K_r9_45 ) , .A2( u2_uk_K_r9_9 ) , .B1( u2_uk_n188 ) , .ZN( u2_uk_n385 ) );
  OAI21_X1 u2_uk_U336 (.ZN( u2_K9_46 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1139 ) , .B2( u2_uk_n1577 ) );
  NAND2_X1 u2_uk_U337 (.A1( u2_uk_K_r7_37 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n1139 ) );
  AOI22_X1 u2_uk_U339 (.B2( u2_uk_K_r10_27 ) , .A2( u2_uk_K_r10_4 ) , .B1( u2_uk_n10 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n515 ) );
  OAI22_X1 u2_uk_U340 (.B1( decrypt ) , .ZN( u2_K10_4 ) , .B2( u2_uk_n1612 ) , .A2( u2_uk_n1631 ) , .A1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U341 (.A1( decrypt ) , .ZN( u2_K7_4 ) , .B2( u2_uk_n1474 ) , .A2( u2_uk_n1497 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U343 (.ZN( u2_K2_4 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1238 ) , .A2( u2_uk_n1267 ) , .A1( u2_uk_n129 ) );
  OAI21_X1 u2_uk_U344 (.ZN( u2_K1_4 ) , .B2( u2_uk_n1184 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n990 ) );
  NAND2_X1 u2_uk_U345 (.A1( u2_key_r_3 ) , .A2( u2_uk_n207 ) , .ZN( u2_uk_n990 ) );
  OAI22_X1 u2_uk_U346 (.B1( decrypt ) , .ZN( u2_K1_40 ) , .B2( u2_uk_n1142 ) , .A2( u2_uk_n1183 ) , .A1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U347 (.A1( decrypt ) , .ZN( u2_K6_40 ) , .A2( u2_uk_n1412 ) , .B2( u2_uk_n1420 ) , .B1( u2_uk_n146 ) );
  INV_X1 u2_uk_U348 (.ZN( u2_K7_46 ) , .A( u2_uk_n1094 ) );
  AOI22_X1 u2_uk_U349 (.A1( decrypt ) , .B2( u2_uk_K_r5_23 ) , .A2( u2_uk_K_r5_31 ) , .ZN( u2_uk_n1094 ) , .B1( u2_uk_n148 ) );
  OAI21_X1 u2_uk_U352 (.ZN( u2_K14_40 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1793 ) , .A( u2_uk_n702 ) );
  NAND2_X1 u2_uk_U353 (.A2( decrypt ) , .A1( u2_uk_K_r12_21 ) , .ZN( u2_uk_n702 ) );
  OAI22_X1 u2_uk_U354 (.ZN( u2_K16_40 ) , .B2( u2_uk_n1188 ) , .A2( u2_uk_n1226 ) , .B1( u2_uk_n238 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U356 (.A1( decrypt ) , .ZN( u2_K13_40 ) , .B2( u2_uk_n1744 ) , .A2( u2_uk_n1754 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U357 (.ZN( u2_K11_40 ) , .A1( u2_uk_n161 ) , .A2( u2_uk_n1634 ) , .B2( u2_uk_n1642 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U358 (.ZN( u2_K8_40 ) , .B2( u2_uk_n1525 ) , .A2( u2_uk_n1531 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U359 (.ZN( u2_K7_40 ) , .A2( u2_uk_n1452 ) , .B2( u2_uk_n1464 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U360 (.ZN( u2_K4_40 ) , .B2( u2_uk_n1342 ) , .A2( u2_uk_n1352 ) , .A1( u2_uk_n146 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U361 (.A1( decrypt ) , .ZN( u2_K2_40 ) , .A2( u2_uk_n1235 ) , .B2( u2_uk_n1266 ) , .B1( u2_uk_n163 ) );
  NAND2_X1 u2_uk_U363 (.A2( decrypt ) , .A1( u2_uk_K_r13_31 ) , .ZN( u2_uk_n942 ) );
  OAI21_X1 u2_uk_U364 (.ZN( u2_K2_33 ) , .A( u2_uk_n1000 ) , .B2( u2_uk_n1258 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U365 (.A1( u2_uk_K_r0_31 ) , .ZN( u2_uk_n1000 ) , .A2( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U366 (.A1( decrypt ) , .ZN( u2_K1_28 ) , .B2( u2_uk_n1143 ) , .A2( u2_uk_n1148 ) , .B1( u2_uk_n214 ) );
  INV_X1 u2_uk_U367 (.A( u2_key_r_8 ) , .ZN( u2_uk_n1148 ) );
  OAI21_X1 u2_uk_U368 (.ZN( u2_K16_28 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1189 ) , .A( u2_uk_n954 ) );
  NAND2_X1 u2_uk_U369 (.A2( decrypt ) , .A1( u2_uk_K_r14_8 ) , .ZN( u2_uk_n954 ) );
  OAI22_X1 u2_uk_U370 (.A1( decrypt ) , .ZN( u2_K14_28 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1791 ) , .A2( u2_uk_n1797 ) );
  OAI22_X1 u2_uk_U371 (.ZN( u2_K11_28 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1642 ) , .A2( u2_uk_n1674 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U372 (.ZN( u2_K6_28 ) , .B2( u2_uk_n1420 ) , .A2( u2_uk_n1447 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U373 (.ZN( u2_K3_28 ) , .B2( u2_uk_n1298 ) , .A2( u2_uk_n1303 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U376 (.A1( decrypt ) , .ZN( u2_K15_28 ) , .B2( u2_uk_n1825 ) , .A2( u2_uk_n1853 ) , .B1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U377 (.ZN( u2_K12_28 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1680 ) , .A2( u2_uk_n1684 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U378 (.ZN( u2_K10_28 ) , .B2( u2_uk_n1610 ) , .A2( u2_uk_n1617 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U379 (.A1( decrypt ) , .ZN( u2_K9_28 ) , .B2( u2_uk_n1577 ) , .A2( u2_uk_n1584 ) , .B1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U380 (.ZN( u2_K7_28 ) , .B2( u2_uk_n1471 ) , .A2( u2_uk_n1480 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U381 (.B1( decrypt ) , .ZN( u2_K5_28 ) , .B2( u2_uk_n1366 ) , .A2( u2_uk_n1370 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U382 (.B1( decrypt ) , .ZN( u2_K15_1 ) , .B2( u2_uk_n1838 ) , .A2( u2_uk_n1857 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U383 (.ZN( u2_K14_1 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1778 ) , .A2( u2_uk_n1783 ) );
  OAI21_X1 u2_uk_U384 (.ZN( u2_K10_1 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1600 ) , .A( u2_uk_n251 ) );
  NAND2_X1 u2_uk_U385 (.A2( decrypt ) , .A1( u2_uk_K_r8_10 ) , .ZN( u2_uk_n251 ) );
  OAI22_X1 u2_uk_U386 (.A1( decrypt ) , .ZN( u2_K6_1 ) , .B2( u2_uk_n1432 ) , .A2( u2_uk_n1448 ) , .B1( u2_uk_n146 ) );
  OAI22_X1 u2_uk_U387 (.B1( decrypt ) , .ZN( u2_K5_1 ) , .B2( u2_uk_n1392 ) , .A2( u2_uk_n1399 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U391 (.ZN( u2_K16_1 ) , .B2( u2_uk_n1218 ) , .A2( u2_uk_n1221 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U394 (.A1( decrypt ) , .ZN( u2_K1_9 ) , .B2( u2_uk_n1179 ) , .A2( u2_uk_n1185 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U395 (.ZN( u2_K13_16 ) , .B2( u2_uk_n1731 ) , .A2( u2_uk_n1736 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U396 (.ZN( u2_K10_16 ) , .B2( u2_uk_n1630 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n250 ) );
  NAND2_X1 u2_uk_U397 (.A1( u2_uk_K_r8_32 ) , .A2( u2_uk_n230 ) , .ZN( u2_uk_n250 ) );
  OAI22_X1 u2_uk_U399 (.ZN( u2_K8_16 ) , .B2( u2_uk_n1506 ) , .A2( u2_uk_n1514 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  NAND2_X1 u2_uk_U401 (.A2( decrypt ) , .A1( u2_uk_K_r5_32 ) , .ZN( u2_uk_n1077 ) );
  OAI22_X1 u2_uk_U402 (.B1( decrypt ) , .ZN( u2_K6_16 ) , .B2( u2_uk_n1436 ) , .A2( u2_uk_n1442 ) , .A1( u2_uk_n148 ) );
  OAI21_X1 u2_uk_U404 (.B1( decrypt ) , .ZN( u2_K3_16 ) , .A( u2_uk_n1006 ) , .B2( u2_uk_n1318 ) );
  NAND2_X1 u2_uk_U405 (.A2( decrypt ) , .A1( u2_uk_K_r1_6 ) , .ZN( u2_uk_n1006 ) );
  OAI22_X1 u2_uk_U406 (.A1( decrypt ) , .ZN( u2_K1_16 ) , .B2( u2_uk_n1162 ) , .A2( u2_uk_n1168 ) , .B1( u2_uk_n214 ) );
  OAI21_X1 u2_uk_U407 (.ZN( u2_K15_9 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1843 ) , .A( u2_uk_n947 ) );
  NAND2_X1 u2_uk_U408 (.A2( decrypt ) , .A1( u2_uk_K_r13_4 ) , .ZN( u2_uk_n947 ) );
  OAI21_X1 u2_uk_U409 (.ZN( u2_K14_9 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1788 ) , .A( u2_uk_n933 ) );
  NAND2_X1 u2_uk_U410 (.A2( decrypt ) , .A1( u2_uk_K_r12_18 ) , .ZN( u2_uk_n933 ) );
  OAI22_X1 u2_uk_U411 (.ZN( u2_K13_9 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1731 ) , .A2( u2_uk_n1743 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U412 (.ZN( u2_K12_9 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1715 ) , .A2( u2_uk_n1722 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U413 (.A1( decrypt ) , .ZN( u2_K11_9 ) , .B2( u2_uk_n1633 ) , .A2( u2_uk_n1663 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U414 (.ZN( u2_K8_9 ) , .A2( u2_uk_n1502 ) , .B2( u2_uk_n1508 ) , .B1( u2_uk_n161 ) , .A1( u2_uk_n92 ) );
  AOI22_X1 u2_uk_U417 (.A1( decrypt ) , .B2( u2_uk_K_r8_28 ) , .A2( u2_uk_K_r8_52 ) , .B1( u2_uk_n147 ) , .ZN( u2_uk_n299 ) );
  INV_X1 u2_uk_U418 (.ZN( u2_K8_37 ) , .A( u2_uk_n1108 ) );
  AOI22_X1 u2_uk_U419 (.B2( u2_uk_K_r6_14 ) , .A2( u2_uk_K_r6_7 ) , .ZN( u2_uk_n1108 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n162 ) );
  AOI22_X1 u2_uk_U421 (.B2( u2_uk_K_r8_17 ) , .A2( u2_uk_K_r8_27 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n308 ) );
  AOI22_X1 u2_uk_U423 (.A2( decrypt ) , .B2( u2_uk_K_r7_13 ) , .A1( u2_uk_K_r7_6 ) , .ZN( u2_uk_n1141 ) , .B1( u2_uk_n217 ) );
  AOI22_X1 u2_uk_U425 (.A1( decrypt ) , .B2( u2_uk_K_r4_3 ) , .A2( u2_uk_K_r4_41 ) , .ZN( u2_uk_n1074 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U426 (.ZN( u2_K7_9 ) , .B2( u2_uk_n1461 ) , .A2( u2_uk_n1468 ) , .A1( u2_uk_n231 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U427 (.B1( decrypt ) , .ZN( u2_K5_9 ) , .B2( u2_uk_n1397 ) , .A2( u2_uk_n1407 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U430 (.ZN( u2_K2_9 ) , .A2( u2_uk_n1232 ) , .B2( u2_uk_n1261 ) , .B1( u2_uk_n145 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U431 (.ZN( u2_K11_1 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1658 ) , .A2( u2_uk_n1675 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U432 (.A1( decrypt ) , .ZN( u2_K2_1 ) , .B2( u2_uk_n1254 ) , .A2( u2_uk_n1275 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U433 (.B1( decrypt ) , .ZN( u2_K16_9 ) , .B2( u2_uk_n1221 ) , .A2( u2_uk_n1228 ) , .A1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U434 (.ZN( u2_K16_16 ) , .B2( u2_uk_n1207 ) , .A2( u2_uk_n1214 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U435 (.B1( decrypt ) , .ZN( u2_K15_16 ) , .A1( u2_uk_n145 ) , .B2( u2_uk_n1829 ) , .A2( u2_uk_n1844 ) );
  OAI22_X1 u2_uk_U436 (.B1( decrypt ) , .ZN( u2_K5_16 ) , .A2( u2_uk_n1367 ) , .B2( u2_uk_n1380 ) , .A1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U437 (.A1( decrypt ) , .ZN( u2_K2_16 ) , .B2( u2_uk_n1244 ) , .A2( u2_uk_n1262 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U438 (.ZN( u2_K4_37 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1331 ) , .A2( u2_uk_n1345 ) , .B1( u2_uk_n238 ) );
  AOI22_X1 u2_uk_U440 (.B2( u2_uk_K_r0_15 ) , .A2( u2_uk_K_r0_49 ) , .A1( u2_uk_n102 ) , .B1( u2_uk_n208 ) , .ZN( u2_uk_n998 ) );
  AOI22_X1 u2_uk_U442 (.B2( u2_uk_K_r14_2 ) , .A2( u2_uk_K_r14_50 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n959 ) );
  OAI22_X1 u2_uk_U443 (.A1( decrypt ) , .ZN( u2_K7_33 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1464 ) , .A2( u2_uk_n1484 ) );
  AOI22_X1 u2_uk_U445 (.B1( decrypt ) , .B2( u2_uk_K_r7_1 ) , .A2( u2_uk_K_r7_8 ) , .ZN( u2_uk_n1132 ) , .A1( u2_uk_n207 ) );
  INV_X1 u2_uk_U448 (.ZN( u2_K1_33 ) , .A( u2_uk_n981 ) );
  AOI22_X1 u2_uk_U449 (.B2( u2_key_r_44 ) , .A2( u2_key_r_51 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n981 ) );
  OAI21_X1 u2_uk_U450 (.ZN( u2_K12_33 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1718 ) , .A( u2_uk_n468 ) );
  NAND2_X1 u2_uk_U451 (.A2( decrypt ) , .A1( u2_uk_K_r10_14 ) , .ZN( u2_uk_n468 ) );
  OAI22_X1 u2_uk_U452 (.ZN( u2_K16_33 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1220 ) , .A2( u2_uk_n1225 ) , .A1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U454 (.ZN( u2_K13_33 ) , .B2( u2_uk_n1723 ) , .A2( u2_uk_n1728 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U455 (.ZN( u2_K11_33 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1653 ) , .A2( u2_uk_n1659 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U456 (.ZN( u2_K8_33 ) , .B2( u2_uk_n1498 ) , .A2( u2_uk_n1503 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U458 (.B1( decrypt ) , .ZN( u2_K4_33 ) , .B2( u2_uk_n1319 ) , .A2( u2_uk_n1326 ) , .A1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U459 (.ZN( u2_K3_33 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1292 ) , .A2( u2_uk_n1309 ) , .B1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U461 (.ZN( u2_K14_37 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1785 ) , .A2( u2_uk_n1791 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U462 (.B1( decrypt ) , .ZN( u2_K13_37 ) , .B2( u2_uk_n1734 ) , .A2( u2_uk_n1746 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U463 (.B1( decrypt ) , .ZN( u2_K12_37 ) , .B2( u2_uk_n1679 ) , .A2( u2_uk_n1719 ) , .A1( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U464 (.ZN( u2_K11_37 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1664 ) , .A( u2_uk_n377 ) );
  NAND2_X1 u2_uk_U465 (.A2( decrypt ) , .A1( u2_uk_K_r9_38 ) , .ZN( u2_uk_n377 ) );
  OAI21_X1 u2_uk_U466 (.ZN( u2_K9_37 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1134 ) , .B2( u2_uk_n1551 ) );
  NAND2_X1 u2_uk_U467 (.A2( decrypt ) , .A1( u2_uk_K_r7_7 ) , .ZN( u2_uk_n1134 ) );
  OAI22_X1 u2_uk_U470 (.ZN( u2_K5_37 ) , .B2( u2_uk_n1365 ) , .A2( u2_uk_n1403 ) , .B1( u2_uk_n147 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U471 (.ZN( u2_K3_37 ) , .B2( u2_uk_n1292 ) , .A2( u2_uk_n1298 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U473 (.B1( decrypt ) , .ZN( u2_K10_36 ) , .B2( u2_uk_n1589 ) , .A( u2_uk_n298 ) );
  NAND2_X1 u2_uk_U474 (.A1( u2_uk_K_r8_21 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n298 ) );
  NAND2_X1 u2_uk_U476 (.A2( decrypt ) , .A1( u2_uk_K_r12_44 ) , .ZN( u2_uk_n689 ) );
  OAI22_X1 u2_uk_U477 (.ZN( u2_K13_29 ) , .B2( u2_uk_n1742 ) , .A2( u2_uk_n1745 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U478 (.ZN( u2_K6_29 ) , .A( u2_uk_n1065 ) , .B2( u2_uk_n1412 ) , .B1( u2_uk_n161 ) );
  NAND2_X1 u2_uk_U479 (.A1( u2_uk_K_r4_0 ) , .ZN( u2_uk_n1065 ) , .A2( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U480 (.A1( decrypt ) , .ZN( u2_K15_29 ) , .A2( u2_uk_n1819 ) , .B2( u2_uk_n1837 ) , .B1( u2_uk_n222 ) );
  AOI22_X1 u2_uk_U482 (.A1( decrypt ) , .B2( u2_uk_K_r14_16 ) , .A2( u2_uk_K_r14_23 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n955 ) );
  OAI21_X1 u2_uk_U485 (.ZN( u2_K3_29 ) , .A( u2_uk_n1010 ) , .B2( u2_uk_n1313 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U486 (.A1( u2_uk_K_r1_44 ) , .ZN( u2_uk_n1010 ) , .A2( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U487 (.ZN( u2_K2_29 ) , .A2( u2_uk_n1237 ) , .B2( u2_uk_n1252 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U488 (.B1( decrypt ) , .ZN( u2_K12_29 ) , .B2( u2_uk_n1691 ) , .A2( u2_uk_n1714 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U489 (.ZN( u2_K10_29 ) , .B2( u2_uk_n1597 ) , .A2( u2_uk_n1625 ) , .B1( u2_uk_n202 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U490 (.A1( decrypt ) , .ZN( u2_K9_29 ) , .B2( u2_uk_n1565 ) , .A2( u2_uk_n1569 ) , .B1( u2_uk_n163 ) );
  INV_X1 u2_uk_U491 (.ZN( u2_K8_29 ) , .A( u2_uk_n1104 ) );
  AOI22_X1 u2_uk_U492 (.A1( decrypt ) , .B2( u2_uk_K_r6_28 ) , .A2( u2_uk_K_r6_35 ) , .ZN( u2_uk_n1104 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U494 (.ZN( u2_K5_29 ) , .B2( u2_uk_n1377 ) , .A2( u2_uk_n1396 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U495 (.A1( decrypt ) , .ZN( u2_K15_2 ) , .B2( u2_uk_n1828 ) , .A2( u2_uk_n1857 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U496 (.ZN( u2_K14_2 ) , .B2( u2_uk_n1794 ) , .A2( u2_uk_n1801 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U499 (.ZN( u2_K8_2 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1105 ) , .B2( u2_uk_n1515 ) );
  NAND2_X1 u2_uk_U500 (.A2( decrypt ) , .A1( u2_uk_K_r6_27 ) , .ZN( u2_uk_n1105 ) );
  OAI22_X1 u2_uk_U501 (.ZN( u2_K5_2 ) , .A2( u2_uk_n1367 ) , .B2( u2_uk_n1372 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U505 (.ZN( u2_K9_12 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1119 ) , .B2( u2_uk_n1543 ) );
  NAND2_X1 u2_uk_U506 (.A2( decrypt ) , .A1( u2_uk_K_r7_53 ) , .ZN( u2_uk_n1119 ) );
  OAI21_X1 u2_uk_U507 (.ZN( u2_K1_12 ) , .B2( u2_uk_n1154 ) , .B1( u2_uk_n93 ) , .A( u2_uk_n968 ) );
  NAND2_X1 u2_uk_U508 (.A1( u2_key_r_12 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n968 ) );
  OAI21_X1 u2_uk_U509 (.ZN( u2_K13_17 ) , .B2( u2_uk_n1743 ) , .A( u2_uk_n587 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U51 (.A( decrypt ) , .ZN( u2_uk_n238 ) );
  NAND2_X1 u2_uk_U510 (.A1( u2_uk_K_r11_27 ) , .ZN( u2_uk_n587 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U511 (.A1( decrypt ) , .ZN( u2_K10_17 ) , .B2( u2_uk_n1596 ) , .A2( u2_uk_n1624 ) , .B1( u2_uk_n187 ) );
  OAI21_X1 u2_uk_U514 (.ZN( u2_K8_17 ) , .A( u2_uk_n1101 ) , .B2( u2_uk_n1522 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U515 (.A1( u2_uk_K_r6_26 ) , .ZN( u2_uk_n1101 ) , .A2( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U520 (.ZN( u2_K11_2 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1643 ) , .A2( u2_uk_n1677 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U521 (.ZN( u2_K15_12 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1815 ) , .B2( u2_uk_n1833 ) );
  OAI22_X1 u2_uk_U522 (.A1( decrypt ) , .ZN( u2_K14_12 ) , .B2( u2_uk_n1801 ) , .A2( u2_uk_n1805 ) , .B1( u2_uk_n223 ) );
  NAND2_X1 u2_uk_U524 (.A2( decrypt ) , .A1( u2_uk_K_r10_11 ) , .ZN( u2_uk_n408 ) );
  AOI22_X1 u2_uk_U53 (.B2( u2_uk_K_r14_2 ) , .A2( u2_uk_K_r14_9 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n238 ) , .ZN( u2_uk_n958 ) );
  OAI22_X1 u2_uk_U531 (.ZN( u2_K2_12 ) , .A2( u2_uk_n1233 ) , .B2( u2_uk_n1248 ) , .A1( u2_uk_n141 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U532 (.ZN( u2_K2_2 ) , .B2( u2_uk_n1243 ) , .A2( u2_uk_n1275 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n31 ) );
  OAI21_X1 u2_uk_U534 (.ZN( u2_K16_12 ) , .B2( u2_uk_n1198 ) , .B1( u2_uk_n208 ) , .A( u2_uk_n949 ) );
  NAND2_X1 u2_uk_U535 (.A1( u2_uk_K_r14_12 ) , .A2( u2_uk_n145 ) , .ZN( u2_uk_n949 ) );
  OAI21_X1 u2_uk_U536 (.ZN( u2_K16_17 ) , .B2( u2_uk_n1197 ) , .B1( u2_uk_n188 ) , .A( u2_uk_n952 ) );
  NAND2_X1 u2_uk_U537 (.A1( u2_uk_K_r14_10 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n952 ) );
  OAI22_X1 u2_uk_U538 (.A1( decrypt ) , .ZN( u2_K9_36 ) , .B2( u2_uk_n1569 ) , .A2( u2_uk_n1575 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U539 (.ZN( u2_K15_17 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1814 ) , .B2( u2_uk_n1832 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U54 (.ZN( u2_K11_34 ) , .A( u2_uk_n375 ) );
  OAI22_X1 u2_uk_U540 (.A1( decrypt ) , .ZN( u2_K14_17 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1780 ) , .A2( u2_uk_n1804 ) );
  OAI22_X1 u2_uk_U541 (.A1( decrypt ) , .ZN( u2_K5_17 ) , .B2( u2_uk_n1374 ) , .A2( u2_uk_n1394 ) , .B1( u2_uk_n148 ) );
  AOI22_X1 u2_uk_U543 (.A1( decrypt ) , .B2( u2_uk_K_r10_18 ) , .A2( u2_uk_K_r10_41 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n415 ) );
  AOI22_X1 u2_uk_U545 (.B2( u2_uk_K_r9_4 ) , .A2( u2_uk_K_r9_55 ) , .A1( u2_uk_n109 ) , .B1( u2_uk_n231 ) , .ZN( u2_uk_n335 ) );
  AOI22_X1 u2_uk_U55 (.B2( u2_uk_K_r9_45 ) , .A2( u2_uk_K_r9_49 ) , .B1( u2_uk_n10 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n375 ) );
  OAI22_X1 u2_uk_U550 (.ZN( u2_K13_36 ) , .B2( u2_uk_n1747 ) , .A2( u2_uk_n1753 ) , .B1( u2_uk_n202 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U552 (.A1( decrypt ) , .ZN( u2_K2_36 ) , .B2( u2_uk_n1242 ) , .A2( u2_uk_n1258 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U554 (.ZN( u2_K12_38 ) , .A1( u2_uk_n10 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1678 ) , .A2( u2_uk_n1705 ) );
  OAI22_X1 u2_uk_U555 (.A1( decrypt ) , .ZN( u2_K11_38 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1640 ) , .A2( u2_uk_n1648 ) );
  OAI22_X1 u2_uk_U556 (.A1( decrypt ) , .ZN( u2_K9_38 ) , .B2( u2_uk_n1575 ) , .A2( u2_uk_n1582 ) , .B1( u2_uk_n188 ) );
  AOI22_X1 u2_uk_U558 (.B2( u2_uk_K_r5_1 ) , .A2( u2_uk_K_r5_21 ) , .ZN( u2_uk_n1091 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n202 ) );
  INV_X1 u2_uk_U559 (.ZN( u2_K11_36 ) , .A( u2_uk_n376 ) );
  INV_X1 u2_uk_U56 (.ZN( u2_K8_34 ) , .A( u2_uk_n1107 ) );
  AOI22_X1 u2_uk_U560 (.A1( decrypt ) , .B2( u2_uk_K_r9_15 ) , .A2( u2_uk_K_r9_7 ) , .B1( u2_uk_n162 ) , .ZN( u2_uk_n376 ) );
  AOI22_X1 u2_uk_U562 (.B2( u2_uk_K_r3_29 ) , .A2( u2_uk_K_r3_52 ) , .ZN( u2_uk_n1050 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U563 (.ZN( u2_K16_36 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1203 ) , .A2( u2_uk_n1210 ) , .A1( u2_uk_n129 ) );
  AOI22_X1 u2_uk_U565 (.A1( decrypt ) , .B2( u2_uk_K_r13_23 ) , .A2( u2_uk_K_r13_44 ) , .B1( u2_uk_n163 ) , .ZN( u2_uk_n943 ) );
  AOI22_X1 u2_uk_U567 (.B2( u2_uk_K_r8_28 ) , .A2( u2_uk_K_r8_8 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n301 ) );
  OAI22_X1 u2_uk_U568 (.ZN( u2_K8_36 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1524 ) , .A2( u2_uk_n1530 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U569 (.ZN( u2_K6_38 ) , .B2( u2_uk_n1418 ) , .A2( u2_uk_n1425 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  AOI22_X1 u2_uk_U57 (.A1( decrypt ) , .B2( u2_uk_K_r6_14 ) , .A2( u2_uk_K_r6_21 ) , .ZN( u2_uk_n1107 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U570 (.B1( decrypt ) , .ZN( u2_K5_38 ) , .B2( u2_uk_n1364 ) , .A2( u2_uk_n1388 ) , .A1( u2_uk_n213 ) );
  OAI21_X1 u2_uk_U571 (.ZN( u2_K15_10 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1839 ) , .A( u2_uk_n934 ) );
  NAND2_X1 u2_uk_U572 (.A1( u2_uk_K_r13_55 ) , .A2( u2_uk_n11 ) , .ZN( u2_uk_n934 ) );
  OAI22_X1 u2_uk_U573 (.A1( decrypt ) , .ZN( u2_K14_10 ) , .B2( u2_uk_n1779 ) , .A2( u2_uk_n1784 ) , .B1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U574 (.ZN( u2_K11_10 ) , .B2( u2_uk_n1633 ) , .A( u2_uk_n312 ) , .B1( u2_uk_n83 ) );
  NAND2_X1 u2_uk_U575 (.A1( u2_uk_K_r9_54 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n312 ) );
  OAI22_X1 u2_uk_U576 (.A1( decrypt ) , .ZN( u2_K10_10 ) , .B1( u2_uk_n155 ) , .B2( u2_uk_n1595 ) , .A2( u2_uk_n1623 ) );
  OAI22_X1 u2_uk_U577 (.A1( decrypt ) , .ZN( u2_K5_10 ) , .B2( u2_uk_n1373 ) , .A2( u2_uk_n1393 ) , .B1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U578 (.ZN( u2_K16_10 ) , .B2( u2_uk_n1219 ) , .A2( u2_uk_n1222 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U581 (.ZN( u2_K8_10 ) , .B2( u2_uk_n1519 ) , .A2( u2_uk_n1521 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U582 (.ZN( u2_K6_10 ) , .A( u2_uk_n1058 ) );
  AOI22_X1 u2_uk_U583 (.B2( u2_uk_K_r4_3 ) , .A2( u2_uk_K_r4_54 ) , .ZN( u2_uk_n1058 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n148 ) );
  INV_X1 u2_uk_U584 (.ZN( u2_K1_10 ) , .A( u2_uk_n966 ) );
  AOI22_X1 u2_uk_U585 (.B2( u2_key_r_41 ) , .A2( u2_key_r_48 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n161 ) , .ZN( u2_uk_n966 ) );
  OAI22_X1 u2_uk_U586 (.A1( decrypt ) , .ZN( u2_K12_22 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1692 ) , .A2( u2_uk_n1702 ) );
  OAI22_X1 u2_uk_U588 (.ZN( u2_K16_22 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1205 ) , .A2( u2_uk_n1212 ) , .A1( u2_uk_n213 ) );
  INV_X1 u2_uk_U589 (.ZN( u2_K13_22 ) , .A( u2_uk_n634 ) );
  AOI22_X1 u2_uk_U59 (.A1( decrypt ) , .B2( u2_uk_K_r5_0 ) , .A2( u2_uk_K_r5_35 ) , .ZN( u2_uk_n1089 ) , .B1( u2_uk_n217 ) );
  AOI22_X1 u2_uk_U590 (.B2( u2_uk_K_r11_10 ) , .A2( u2_uk_K_r11_47 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n634 ) , .B1( u2_uk_n94 ) );
  INV_X1 u2_uk_U591 (.ZN( u2_K11_22 ) , .A( u2_uk_n349 ) );
  AOI22_X1 u2_uk_U592 (.B2( u2_uk_K_r9_13 ) , .A2( u2_uk_K_r9_19 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n349 ) );
  AOI22_X1 u2_uk_U594 (.B1( decrypt ) , .B2( u2_uk_K_r8_27 ) , .A2( u2_uk_K_r8_5 ) , .A1( u2_uk_n220 ) , .ZN( u2_uk_n257 ) );
  OAI22_X1 u2_uk_U597 (.ZN( u2_K8_22 ) , .B2( u2_uk_n1529 ) , .A2( u2_uk_n1535 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U598 (.ZN( u2_K7_22 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1081 ) , .B2( u2_uk_n1468 ) );
  NAND2_X1 u2_uk_U599 (.A2( decrypt ) , .A1( u2_uk_K_r5_5 ) , .ZN( u2_uk_n1081 ) );
  OAI22_X1 u2_uk_U60 (.A1( decrypt ) , .ZN( u2_K15_34 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1826 ) , .A2( u2_uk_n1854 ) );
  INV_X1 u2_uk_U600 (.ZN( u2_K5_22 ) , .A( u2_uk_n1044 ) );
  AOI22_X1 u2_uk_U601 (.A1( decrypt ) , .B2( u2_uk_K_r3_24 ) , .A2( u2_uk_K_r3_33 ) , .ZN( u2_uk_n1044 ) , .B1( u2_uk_n214 ) );
  INV_X1 u2_uk_U602 (.ZN( u2_K1_22 ) , .A( u2_uk_n974 ) );
  AOI22_X1 u2_uk_U603 (.B2( u2_key_r_25 ) , .A2( u2_key_r_32 ) , .B1( u2_uk_n109 ) , .A1( u2_uk_n191 ) , .ZN( u2_uk_n974 ) );
  OAI22_X1 u2_uk_U604 (.ZN( u2_K16_35 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1208 ) , .A2( u2_uk_n1215 ) , .A1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U605 (.ZN( u2_K11_35 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1665 ) , .A2( u2_uk_n1673 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U606 (.ZN( u2_K8_35 ) , .B2( u2_uk_n1511 ) , .A2( u2_uk_n1517 ) , .A1( u2_uk_n203 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U607 (.B1( decrypt ) , .ZN( u2_K7_35 ) , .A( u2_uk_n1090 ) , .B2( u2_uk_n1452 ) );
  NAND2_X1 u2_uk_U608 (.A1( u2_uk_K_r5_37 ) , .ZN( u2_uk_n1090 ) , .A2( u2_uk_n11 ) );
  OAI22_X1 u2_uk_U609 (.B1( decrypt ) , .ZN( u2_K15_35 ) , .B2( u2_uk_n1830 ) , .A2( u2_uk_n1845 ) , .A1( u2_uk_n188 ) );
  INV_X1 u2_uk_U61 (.ZN( u2_K14_34 ) , .A( u2_uk_n692 ) );
  OAI22_X1 u2_uk_U610 (.ZN( u2_K13_35 ) , .B2( u2_uk_n1734 ) , .A2( u2_uk_n1763 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U611 (.ZN( u2_K12_35 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1698 ) , .A2( u2_uk_n1707 ) , .B1( u2_uk_n230 ) );
  INV_X1 u2_uk_U612 (.ZN( u2_K14_35 ) , .A( u2_uk_n694 ) );
  AOI22_X1 u2_uk_U613 (.B2( u2_uk_K_r12_1 ) , .A2( u2_uk_K_r12_7 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n694 ) );
  AOI22_X1 u2_uk_U617 (.B2( u2_uk_K_r7_16 ) , .A2( u2_uk_K_r7_23 ) , .B1( u2_uk_n102 ) , .ZN( u2_uk_n1133 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U619 (.B1( decrypt ) , .ZN( u2_K4_35 ) , .B2( u2_uk_n1331 ) , .A2( u2_uk_n1360 ) , .A1( u2_uk_n164 ) );
  AOI22_X1 u2_uk_U62 (.B2( u2_uk_K_r12_30 ) , .A2( u2_uk_K_r12_36 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n692 ) );
  OAI22_X1 u2_uk_U620 (.A1( decrypt ) , .ZN( u2_K2_35 ) , .B2( u2_uk_n1245 ) , .A2( u2_uk_n1263 ) , .B1( u2_uk_n164 ) );
  INV_X1 u2_uk_U621 (.ZN( u2_K1_35 ) , .A( u2_uk_n982 ) );
  AOI22_X1 u2_uk_U622 (.B2( u2_key_r_28 ) , .A2( u2_key_r_35 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n982 ) );
  OAI21_X1 u2_uk_U623 (.ZN( u2_K16_11 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1212 ) , .A( u2_uk_n948 ) );
  NAND2_X1 u2_uk_U624 (.A2( decrypt ) , .A1( u2_uk_K_r14_39 ) , .ZN( u2_uk_n948 ) );
  OAI21_X1 u2_uk_U626 (.ZN( u2_K15_11 ) , .B2( u2_uk_n1850 ) , .B1( u2_uk_n231 ) , .A( u2_uk_n935 ) );
  NAND2_X1 u2_uk_U627 (.A1( u2_uk_K_r13_25 ) , .A2( u2_uk_n207 ) , .ZN( u2_uk_n935 ) );
  OAI22_X1 u2_uk_U628 (.B1( decrypt ) , .ZN( u2_K14_11 ) , .A1( u2_uk_n142 ) , .A2( u2_uk_n1771 ) , .B2( u2_uk_n1778 ) );
  OAI22_X1 u2_uk_U629 (.A1( decrypt ) , .ZN( u2_K11_11 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1646 ) , .A2( u2_uk_n1652 ) );
  OAI22_X1 u2_uk_U63 (.A1( decrypt ) , .ZN( u2_K12_34 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1685 ) , .B2( u2_uk_n1700 ) );
  INV_X1 u2_uk_U630 (.ZN( u2_K13_11 ) , .A( u2_uk_n526 ) );
  AOI22_X1 u2_uk_U631 (.B1( decrypt ) , .B2( u2_uk_K_r11_17 ) , .A2( u2_uk_K_r11_54 ) , .A1( u2_uk_n231 ) , .ZN( u2_uk_n526 ) );
  OAI22_X1 u2_uk_U632 (.B1( decrypt ) , .ZN( u2_K10_11 ) , .B2( u2_uk_n1596 ) , .A2( u2_uk_n1613 ) , .A1( u2_uk_n187 ) );
  OAI21_X1 u2_uk_U633 (.ZN( u2_K8_11 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1097 ) , .B2( u2_uk_n1535 ) );
  NAND2_X1 u2_uk_U634 (.A2( decrypt ) , .A1( u2_uk_K_r6_55 ) , .ZN( u2_uk_n1097 ) );
  OAI22_X1 u2_uk_U637 (.B1( decrypt ) , .ZN( u2_K6_11 ) , .B2( u2_uk_n1423 ) , .A2( u2_uk_n1427 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U638 (.A1( decrypt ) , .ZN( u2_K5_11 ) , .A2( u2_uk_n1369 ) , .B2( u2_uk_n1393 ) , .B1( u2_uk_n147 ) );
  OAI21_X1 u2_uk_U64 (.B1( decrypt ) , .ZN( u2_K6_34 ) , .A( u2_uk_n1067 ) , .B2( u2_uk_n1441 ) );
  OAI21_X1 u2_uk_U640 (.ZN( u2_K2_11 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1267 ) , .A( u2_uk_n992 ) );
  NAND2_X1 u2_uk_U641 (.A1( u2_uk_K_r0_25 ) , .A2( u2_uk_n100 ) , .ZN( u2_uk_n992 ) );
  OAI21_X1 u2_uk_U642 (.B1( decrypt ) , .ZN( u2_K4_6 ) , .A( u2_uk_n1039 ) , .B2( u2_uk_n1335 ) );
  NAND2_X1 u2_uk_U643 (.A1( u2_uk_K_r2_24 ) , .ZN( u2_uk_n1039 ) , .A2( u2_uk_n60 ) );
  AOI22_X1 u2_uk_U645 (.B2( u2_key_r_36 ) , .A2( u2_key_r_43 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n182 ) , .ZN( u2_uk_n987 ) );
  OAI21_X1 u2_uk_U646 (.ZN( u2_K12_6 ) , .B1( u2_uk_n162 ) , .B2( u2_uk_n1702 ) , .A( u2_uk_n518 ) );
  NAND2_X1 u2_uk_U647 (.A1( u2_uk_K_r10_10 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n518 ) );
  OAI22_X1 u2_uk_U648 (.ZN( u2_K16_45 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1217 ) , .A2( u2_uk_n1220 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U649 (.A1( decrypt ) , .ZN( u2_K1_45 ) , .B2( u2_uk_n1171 ) , .A2( u2_uk_n1178 ) , .B1( u2_uk_n230 ) );
  NAND2_X1 u2_uk_U65 (.A2( decrypt ) , .A1( u2_uk_K_r4_49 ) , .ZN( u2_uk_n1067 ) );
  INV_X1 u2_uk_U650 (.A( u2_key_r_44 ) , .ZN( u2_uk_n1178 ) );
  OAI22_X1 u2_uk_U651 (.ZN( u2_K14_43 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1799 ) , .A2( u2_uk_n1802 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U652 (.ZN( u2_K9_43 ) , .A1( u2_uk_n102 ) , .B2( u2_uk_n1558 ) , .A2( u2_uk_n1565 ) , .B1( u2_uk_n214 ) );
  OAI21_X1 u2_uk_U653 (.ZN( u2_K4_43 ) , .A( u2_uk_n1036 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1359 ) );
  NAND2_X1 u2_uk_U654 (.A2( decrypt ) , .A1( u2_uk_K_r2_29 ) , .ZN( u2_uk_n1036 ) );
  OAI22_X1 u2_uk_U655 (.B1( decrypt ) , .ZN( u2_K3_43 ) , .B2( u2_uk_n1304 ) , .A2( u2_uk_n1308 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U656 (.B1( decrypt ) , .ZN( u2_K2_43 ) , .A( u2_uk_n1002 ) , .B2( u2_uk_n1246 ) );
  NAND2_X1 u2_uk_U657 (.A2( decrypt ) , .A1( u2_uk_K_r0_2 ) , .ZN( u2_uk_n1002 ) );
  OAI22_X1 u2_uk_U658 (.ZN( u2_K1_7 ) , .B2( u2_uk_n1155 ) , .A2( u2_uk_n1162 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U659 (.A1( decrypt ) , .ZN( u2_K4_7 ) , .A2( u2_uk_n1323 ) , .B2( u2_uk_n1327 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U66 (.A1( decrypt ) , .ZN( u2_K4_34 ) , .B2( u2_uk_n1336 ) , .A2( u2_uk_n1352 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U660 (.A1( decrypt ) , .ZN( u2_K9_25 ) , .B2( u2_uk_n1578 ) , .A2( u2_uk_n1585 ) , .B1( u2_uk_n238 ) );
  AOI22_X1 u2_uk_U662 (.B2( u2_uk_K_r14_16 ) , .A2( u2_uk_K_r14_9 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n161 ) , .ZN( u2_uk_n963 ) );
  AOI22_X1 u2_uk_U664 (.B2( u2_uk_K_r3_15 ) , .A2( u2_uk_K_r3_38 ) , .ZN( u2_uk_n1053 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n155 ) );
  OAI21_X1 u2_uk_U665 (.ZN( u2_K14_45 ) , .B2( u2_uk_n1800 ) , .B1( u2_uk_n238 ) , .A( u2_uk_n930 ) );
  NAND2_X1 u2_uk_U666 (.A1( u2_uk_K_r12_16 ) , .A2( u2_uk_n220 ) , .ZN( u2_uk_n930 ) );
  OAI21_X1 u2_uk_U667 (.ZN( u2_K13_43 ) , .B2( u2_uk_n1762 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n676 ) );
  NAND2_X1 u2_uk_U668 (.A1( u2_uk_K_r11_29 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n676 ) );
  OAI21_X1 u2_uk_U669 (.ZN( u2_K12_45 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1684 ) , .A( u2_uk_n509 ) );
  OAI21_X1 u2_uk_U67 (.ZN( u2_K3_34 ) , .A( u2_uk_n1011 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1299 ) );
  NAND2_X1 u2_uk_U670 (.A1( u2_uk_K_r10_43 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n509 ) );
  OAI22_X1 u2_uk_U671 (.ZN( u2_K11_43 ) , .A1( u2_uk_n161 ) , .B2( u2_uk_n1632 ) , .A2( u2_uk_n1674 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U672 (.B1( decrypt ) , .ZN( u2_K10_43 ) , .A2( u2_uk_n1593 ) , .B2( u2_uk_n1621 ) , .A1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U673 (.ZN( u2_K10_45 ) , .B2( u2_uk_n1598 ) , .A2( u2_uk_n1614 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U674 (.B1( decrypt ) , .ZN( u2_K9_45 ) , .B2( u2_uk_n1541 ) , .A2( u2_uk_n1582 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U675 (.A1( decrypt ) , .ZN( u2_K7_43 ) , .A2( u2_uk_n1455 ) , .B2( u2_uk_n1484 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U676 (.ZN( u2_K16_3 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1198 ) , .A2( u2_uk_n1206 ) , .A1( u2_uk_n191 ) );
  OAI21_X1 u2_uk_U677 (.B1( decrypt ) , .ZN( u2_K14_3 ) , .B2( u2_uk_n1812 ) , .A( u2_uk_n695 ) );
  NAND2_X1 u2_uk_U678 (.A2( decrypt ) , .A1( u2_uk_K_r12_47 ) , .ZN( u2_uk_n695 ) );
  OAI22_X1 u2_uk_U679 (.ZN( u2_K10_7 ) , .B2( u2_uk_n1604 ) , .A2( u2_uk_n1624 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n83 ) );
  NAND2_X1 u2_uk_U68 (.A2( decrypt ) , .A1( u2_uk_K_r1_36 ) , .ZN( u2_uk_n1011 ) );
  OAI22_X1 u2_uk_U684 (.ZN( u2_K15_7 ) , .A1( u2_uk_n163 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1823 ) , .A2( u2_uk_n1839 ) );
  OAI21_X1 u2_uk_U685 (.B1( decrypt ) , .ZN( u2_K11_7 ) , .B2( u2_uk_n1661 ) , .A( u2_uk_n395 ) );
  NAND2_X1 u2_uk_U686 (.A1( u2_uk_K_r9_33 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n395 ) );
  OAI22_X1 u2_uk_U687 (.ZN( u2_K16_7 ) , .B2( u2_uk_n1199 ) , .A2( u2_uk_n1207 ) , .A1( u2_uk_n141 ) , .B1( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U688 (.ZN( u2_K11_25 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1647 ) , .A2( u2_uk_n1666 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U689 (.ZN( u2_K13_25 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1735 ) , .A2( u2_uk_n1760 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U69 (.B1( decrypt ) , .ZN( u2_K2_34 ) , .B2( u2_uk_n1242 ) , .A2( u2_uk_n1273 ) , .A1( u2_uk_n161 ) );
  OAI21_X1 u2_uk_U690 (.B1( decrypt ) , .ZN( u2_K5_25 ) , .A( u2_uk_n1045 ) , .B2( u2_uk_n1383 ) );
  NAND2_X1 u2_uk_U691 (.A2( decrypt ) , .A1( u2_uk_K_r3_35 ) , .ZN( u2_uk_n1045 ) );
  OAI21_X1 u2_uk_U692 (.ZN( u2_K2_25 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1264 ) , .A( u2_uk_n996 ) );
  NAND2_X1 u2_uk_U693 (.A2( decrypt ) , .A1( u2_uk_K_r0_22 ) , .ZN( u2_uk_n996 ) );
  OAI22_X1 u2_uk_U694 (.A1( decrypt ) , .ZN( u2_K12_25 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1699 ) , .A2( u2_uk_n1704 ) );
  OAI22_X1 u2_uk_U695 (.A1( decrypt ) , .ZN( u2_K10_25 ) , .B1( u2_uk_n146 ) , .A2( u2_uk_n1593 ) , .B2( u2_uk_n1611 ) );
  OAI22_X1 u2_uk_U696 (.ZN( u2_K8_25 ) , .B2( u2_uk_n1533 ) , .A2( u2_uk_n1538 ) , .A1( u2_uk_n222 ) , .B1( u2_uk_n27 ) );
  AOI22_X1 u2_uk_U698 (.A1( decrypt ) , .B2( u2_uk_K_r11_10 ) , .A2( u2_uk_K_r11_5 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n682 ) );
  OAI22_X1 u2_uk_U70 (.ZN( u2_K16_23 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1213 ) , .A2( u2_uk_n1218 ) , .A1( u2_uk_n164 ) );
  AOI22_X1 u2_uk_U702 (.B2( u2_uk_K_r5_31 ) , .A2( u2_uk_K_r5_7 ) , .A1( u2_uk_n10 ) , .ZN( u2_uk_n1084 ) , .B1( u2_uk_n217 ) );
  INV_X1 u2_uk_U703 (.ZN( u2_K1_25 ) , .A( u2_uk_n975 ) );
  AOI22_X1 u2_uk_U704 (.B2( u2_key_r_29 ) , .A2( u2_key_r_36 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n975 ) );
  AOI22_X1 u2_uk_U706 (.A1( decrypt ) , .B2( u2_uk_K_r2_16 ) , .A2( u2_uk_K_r2_49 ) , .ZN( u2_uk_n1027 ) , .B1( u2_uk_n148 ) );
  OAI22_X1 u2_uk_U709 (.ZN( u2_K16_25 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1209 ) , .A2( u2_uk_n1216 ) , .A1( u2_uk_n208 ) );
  OAI21_X1 u2_uk_U71 (.ZN( u2_K11_23 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1668 ) , .A( u2_uk_n353 ) );
  OAI22_X1 u2_uk_U710 (.B1( decrypt ) , .ZN( u2_K12_2 ) , .A2( u2_uk_n1681 ) , .B2( u2_uk_n1686 ) , .A1( u2_uk_n182 ) );
  OAI21_X1 u2_uk_U711 (.ZN( u2_K1_2 ) , .B2( u2_uk_n1145 ) , .B1( u2_uk_n220 ) , .A( u2_uk_n978 ) );
  NAND2_X1 u2_uk_U712 (.A1( u2_key_r_11 ) , .A2( u2_uk_n191 ) , .ZN( u2_uk_n978 ) );
  OAI22_X1 u2_uk_U714 (.ZN( u2_K16_32 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1201 ) , .A2( u2_uk_n1209 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U715 (.ZN( u2_K8_32 ) , .B2( u2_uk_n1526 ) , .A2( u2_uk_n1533 ) , .A1( u2_uk_n238 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U716 (.ZN( u2_K11_32 ) , .B2( u2_uk_n1640 ) , .A2( u2_uk_n1660 ) , .A1( u2_uk_n203 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U717 (.B1( decrypt ) , .ZN( u2_K13_32 ) , .A2( u2_uk_n1728 ) , .B2( u2_uk_n1752 ) , .A1( u2_uk_n220 ) );
  OAI21_X1 u2_uk_U718 (.B1( decrypt ) , .ZN( u2_K10_32 ) , .B2( u2_uk_n1588 ) , .A( u2_uk_n292 ) );
  NAND2_X1 u2_uk_U719 (.A2( decrypt ) , .A1( u2_uk_K_r8_51 ) , .ZN( u2_uk_n292 ) );
  NAND2_X1 u2_uk_U72 (.A1( u2_uk_K_r9_27 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n353 ) );
  OAI22_X1 u2_uk_U720 (.A1( decrypt ) , .ZN( u2_K6_32 ) , .B2( u2_uk_n1418 ) , .A2( u2_uk_n1434 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U721 (.A1( decrypt ) , .ZN( u2_K3_32 ) , .B2( u2_uk_n1278 ) , .A2( u2_uk_n1313 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U722 (.B1( decrypt ) , .ZN( u2_K5_32 ) , .B2( u2_uk_n1378 ) , .A2( u2_uk_n1382 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U724 (.A1( decrypt ) , .ZN( u2_K9_32 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1571 ) , .A2( u2_uk_n1578 ) );
  OAI21_X1 u2_uk_U725 (.B1( decrypt ) , .ZN( u2_K16_42 ) , .B2( u2_uk_n1211 ) , .A( u2_uk_n962 ) );
  NAND2_X1 u2_uk_U726 (.A2( decrypt ) , .A1( u2_uk_K_r14_38 ) , .ZN( u2_uk_n962 ) );
  OAI22_X1 u2_uk_U728 (.A1( decrypt ) , .ZN( u2_K14_42 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1768 ) , .A2( u2_uk_n1799 ) );
  OAI22_X1 u2_uk_U729 (.A1( decrypt ) , .ZN( u2_K13_42 ) , .B2( u2_uk_n1733 ) , .A2( u2_uk_n1739 ) , .B1( u2_uk_n203 ) );
  OAI21_X1 u2_uk_U73 (.ZN( u2_K10_23 ) , .B2( u2_uk_n1590 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n271 ) );
  OAI22_X1 u2_uk_U730 (.A1( decrypt ) , .ZN( u2_K11_42 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1664 ) , .A2( u2_uk_n1672 ) );
  OAI22_X1 u2_uk_U731 (.A1( decrypt ) , .ZN( u2_K10_42 ) , .B2( u2_uk_n1589 ) , .A2( u2_uk_n1615 ) , .B1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U732 (.ZN( u2_K8_42 ) , .A( u2_uk_n1112 ) , .B2( u2_uk_n1510 ) , .B1( u2_uk_n17 ) );
  NAND2_X1 u2_uk_U733 (.A2( decrypt ) , .A1( u2_uk_K_r6_22 ) , .ZN( u2_uk_n1112 ) );
  OAI22_X1 u2_uk_U734 (.B1( decrypt ) , .ZN( u2_K4_42 ) , .B2( u2_uk_n1330 ) , .A2( u2_uk_n1337 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U735 (.B1( decrypt ) , .ZN( u2_K3_42 ) , .B2( u2_uk_n1277 ) , .A2( u2_uk_n1304 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U736 (.ZN( u2_K2_42 ) , .B2( u2_uk_n1266 ) , .A2( u2_uk_n1274 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  AOI22_X1 u2_uk_U738 (.A1( decrypt ) , .B2( u2_uk_K_r5_1 ) , .A2( u2_uk_K_r5_36 ) , .ZN( u2_uk_n1093 ) , .B1( u2_uk_n147 ) );
  NAND2_X1 u2_uk_U74 (.A1( u2_uk_K_r8_13 ) , .A2( u2_uk_n129 ) , .ZN( u2_uk_n271 ) );
  AOI22_X1 u2_uk_U740 (.B1( decrypt ) , .B2( u2_key_r_31 ) , .A2( u2_key_r_38 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n986 ) );
  OAI21_X1 u2_uk_U741 (.ZN( u2_K14_27 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1809 ) , .A( u2_uk_n688 ) );
  NAND2_X1 u2_uk_U742 (.A1( u2_uk_K_r12_42 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n688 ) );
  OAI22_X1 u2_uk_U743 (.A1( decrypt ) , .ZN( u2_K12_27 ) , .B1( u2_uk_n129 ) , .B2( u2_uk_n1687 ) , .A2( u2_uk_n1719 ) );
  OAI21_X1 u2_uk_U744 (.ZN( u2_K10_27 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1602 ) , .A( u2_uk_n279 ) );
  NAND2_X1 u2_uk_U745 (.A1( u2_uk_K_r8_43 ) , .ZN( u2_uk_n279 ) , .A2( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U746 (.ZN( u2_K8_27 ) , .B2( u2_uk_n1499 ) , .A2( u2_uk_n1504 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U747 (.ZN( u2_K16_27 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1195 ) , .A2( u2_uk_n1200 ) , .A1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U749 (.A1( decrypt ) , .ZN( u2_K11_13 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1658 ) , .A2( u2_uk_n1662 ) );
  OAI22_X1 u2_uk_U75 (.ZN( u2_K8_23 ) , .B2( u2_uk_n1513 ) , .A2( u2_uk_n1518 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U750 (.ZN( u2_K8_13 ) , .A2( u2_uk_n1501 ) , .B2( u2_uk_n1507 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U751 (.B1( decrypt ) , .ZN( u2_K6_13 ) , .B2( u2_uk_n1432 ) , .A2( u2_uk_n1436 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U752 (.ZN( u2_K2_13 ) , .A2( u2_uk_n1231 ) , .B2( u2_uk_n1260 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U753 (.ZN( u2_K1_21 ) , .B2( u2_uk_n1153 ) , .A2( u2_uk_n1159 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n83 ) );
  NAND2_X1 u2_uk_U755 (.A2( decrypt ) , .A1( u2_uk_K_r7_5 ) , .ZN( u2_uk_n1120 ) );
  OAI22_X1 u2_uk_U756 (.ZN( u2_K11_27 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1654 ) , .A2( u2_uk_n1660 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U757 (.ZN( u2_K13_27 ) , .A1( u2_uk_n128 ) , .B2( u2_uk_n1724 ) , .A2( u2_uk_n1747 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U758 (.A1( decrypt ) , .ZN( u2_K14_21 ) , .B2( u2_uk_n1784 ) , .A2( u2_uk_n1810 ) , .B1( u2_uk_n230 ) );
  OAI21_X1 u2_uk_U759 (.B1( decrypt ) , .ZN( u2_K11_21 ) , .B2( u2_uk_n1637 ) , .A( u2_uk_n346 ) );
  NAND2_X1 u2_uk_U760 (.A1( u2_uk_K_r9_5 ) , .A2( u2_uk_n27 ) , .ZN( u2_uk_n346 ) );
  OAI22_X1 u2_uk_U762 (.A1( decrypt ) , .ZN( u2_K5_21 ) , .B2( u2_uk_n1379 ) , .A2( u2_uk_n1399 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U763 (.B1( decrypt ) , .ZN( u2_K4_21 ) , .B2( u2_uk_n1341 ) , .A2( u2_uk_n1347 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U764 (.ZN( u2_K2_21 ) , .A2( u2_uk_n1234 ) , .B2( u2_uk_n1238 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U765 (.A1( decrypt ) , .ZN( u2_K14_13 ) , .B2( u2_uk_n1782 ) , .A2( u2_uk_n1787 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U766 (.B1( decrypt ) , .ZN( u2_K15_21 ) , .A1( u2_uk_n148 ) , .A2( u2_uk_n1816 ) , .B2( u2_uk_n1820 ) );
  OAI22_X1 u2_uk_U767 (.ZN( u2_K15_27 ) , .A2( u2_uk_n1817 ) , .B2( u2_uk_n1835 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U768 (.ZN( u2_K2_27 ) , .A( u2_uk_n997 ) );
  AOI22_X1 u2_uk_U769 (.A1( decrypt ) , .B2( u2_uk_K_r0_28 ) , .A2( u2_uk_K_r0_7 ) , .B1( u2_uk_n188 ) , .ZN( u2_uk_n997 ) );
  INV_X1 u2_uk_U770 (.ZN( u2_K12_21 ) , .A( u2_uk_n443 ) );
  AOI22_X1 u2_uk_U771 (.A1( decrypt ) , .B2( u2_uk_K_r10_25 ) , .A2( u2_uk_K_r10_48 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n443 ) );
  OAI21_X1 u2_uk_U772 (.ZN( u2_K3_27 ) , .A( u2_uk_n1009 ) , .B2( u2_uk_n1315 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U773 (.A1( u2_uk_K_r1_42 ) , .ZN( u2_uk_n1009 ) , .A2( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U774 (.B1( decrypt ) , .ZN( u2_K4_27 ) , .B2( u2_uk_n1320 ) , .A2( u2_uk_n1346 ) , .A1( u2_uk_n182 ) );
  INV_X1 u2_uk_U776 (.ZN( u2_K13_21 ) , .A( u2_uk_n608 ) );
  AOI22_X1 u2_uk_U777 (.B1( decrypt ) , .B2( u2_uk_K_r11_34 ) , .A2( u2_uk_K_r11_39 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n608 ) );
  OAI22_X1 u2_uk_U78 (.A1( decrypt ) , .ZN( u2_K3_23 ) , .A2( u2_uk_n1281 ) , .B2( u2_uk_n1286 ) , .B1( u2_uk_n141 ) );
  OAI21_X1 u2_uk_U780 (.ZN( u2_K16_13 ) , .B2( u2_uk_n1227 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n950 ) );
  NAND2_X1 u2_uk_U781 (.A1( u2_uk_K_r14_46 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n950 ) );
  OAI22_X1 u2_uk_U784 (.B1( decrypt ) , .ZN( u2_K6_27 ) , .B2( u2_uk_n1429 ) , .A2( u2_uk_n1434 ) , .A1( u2_uk_n231 ) );
  AOI22_X1 u2_uk_U786 (.A1( decrypt ) , .B2( u2_uk_K_r3_15 ) , .A2( u2_uk_K_r3_51 ) , .ZN( u2_uk_n1046 ) , .B1( u2_uk_n209 ) );
  INV_X1 u2_uk_U787 (.ZN( u2_K13_13 ) , .A( u2_uk_n582 ) );
  AOI22_X1 u2_uk_U788 (.B2( u2_uk_K_r11_11 ) , .A2( u2_uk_K_r11_6 ) , .B1( u2_uk_n214 ) , .ZN( u2_uk_n582 ) , .A1( u2_uk_n83 ) );
  INV_X1 u2_uk_U789 (.ZN( u2_K7_27 ) , .A( u2_uk_n1085 ) );
  OAI22_X1 u2_uk_U79 (.ZN( u2_K2_23 ) , .B2( u2_uk_n1248 ) , .A2( u2_uk_n1269 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  AOI22_X1 u2_uk_U790 (.B2( u2_uk_K_r5_23 ) , .A2( u2_uk_K_r5_43 ) , .ZN( u2_uk_n1085 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n141 ) );
  INV_X1 u2_uk_U791 (.ZN( u2_K1_27 ) , .A( u2_uk_n977 ) );
  AOI22_X1 u2_uk_U792 (.B2( u2_key_r_14 ) , .A2( u2_key_r_21 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n977 ) );
  INV_X1 u2_uk_U793 (.ZN( u2_K9_27 ) , .A( u2_uk_n1129 ) );
  AOI22_X1 u2_uk_U794 (.B2( u2_uk_K_r7_2 ) , .A2( u2_uk_K_r7_9 ) , .B1( u2_uk_n109 ) , .ZN( u2_uk_n1129 ) , .A1( u2_uk_n163 ) );
  OAI21_X1 u2_uk_U795 (.ZN( u2_K13_1 ) , .B1( u2_uk_n109 ) , .B2( u2_uk_n1727 ) , .A( u2_uk_n603 ) );
  NAND2_X1 u2_uk_U796 (.A1( u2_uk_K_r11_25 ) , .ZN( u2_uk_n603 ) , .A2( u2_uk_n93 ) );
  INV_X1 u2_uk_U797 (.ZN( u2_K9_1 ) , .A( u2_uk_n1125 ) );
  AOI22_X1 u2_uk_U798 (.B1( decrypt ) , .B2( u2_uk_K_r7_24 ) , .A2( u2_uk_K_r7_6 ) , .ZN( u2_uk_n1125 ) , .A1( u2_uk_n162 ) );
  OAI21_X1 u2_uk_U799 (.ZN( u2_K4_18 ) , .B1( u2_uk_n10 ) , .A( u2_uk_n1022 ) , .B2( u2_uk_n1348 ) );
  OAI21_X1 u2_uk_U80 (.ZN( u2_K16_41 ) , .B2( u2_uk_n1215 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n961 ) );
  NAND2_X1 u2_uk_U800 (.A2( decrypt ) , .A1( u2_uk_K_r2_20 ) , .ZN( u2_uk_n1022 ) );
  OAI22_X1 u2_uk_U801 (.B1( decrypt ) , .ZN( u2_K5_18 ) , .A2( u2_uk_n1369 ) , .B2( u2_uk_n1406 ) , .A1( u2_uk_n207 ) );
  OAI21_X1 u2_uk_U803 (.B1( decrypt ) , .ZN( u2_K13_20 ) , .B2( u2_uk_n1732 ) , .A( u2_uk_n605 ) );
  NAND2_X1 u2_uk_U804 (.A1( u2_uk_K_r11_33 ) , .ZN( u2_uk_n605 ) , .A2( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U805 (.B1( decrypt ) , .ZN( u2_K8_18 ) , .A( u2_uk_n1102 ) , .B2( u2_uk_n1527 ) );
  NAND2_X1 u2_uk_U806 (.A1( u2_uk_K_r6_46 ) , .ZN( u2_uk_n1102 ) , .A2( u2_uk_n17 ) );
  OAI22_X1 u2_uk_U807 (.B1( decrypt ) , .ZN( u2_K2_18 ) , .B2( u2_uk_n1239 ) , .A2( u2_uk_n1270 ) , .A1( u2_uk_n223 ) );
  OAI21_X1 u2_uk_U808 (.ZN( u2_K16_18 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1229 ) , .A( u2_uk_n953 ) );
  NAND2_X1 u2_uk_U809 (.A1( u2_uk_K_r14_5 ) , .A2( u2_uk_n109 ) , .ZN( u2_uk_n953 ) );
  NAND2_X1 u2_uk_U81 (.A2( decrypt ) , .A1( u2_uk_K_r14_42 ) , .ZN( u2_uk_n961 ) );
  OAI22_X1 u2_uk_U810 (.ZN( u2_K10_18 ) , .A1( u2_uk_n110 ) , .A2( u2_uk_n1590 ) , .B2( u2_uk_n1604 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U811 (.A1( decrypt ) , .ZN( u2_K15_18 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1822 ) , .A2( u2_uk_n1852 ) );
  OAI21_X1 u2_uk_U812 (.ZN( u2_K13_18 ) , .B2( u2_uk_n1750 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n590 ) );
  NAND2_X1 u2_uk_U813 (.A1( u2_uk_K_r11_20 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n590 ) );
  OAI22_X1 u2_uk_U814 (.B1( decrypt ) , .ZN( u2_K3_20 ) , .B2( u2_uk_n1290 ) , .A2( u2_uk_n1296 ) , .A1( u2_uk_n202 ) );
  OAI21_X1 u2_uk_U815 (.B1( decrypt ) , .ZN( u2_K12_20 ) , .B2( u2_uk_n1692 ) , .A( u2_uk_n437 ) );
  NAND2_X1 u2_uk_U816 (.A2( decrypt ) , .A1( u2_uk_K_r10_47 ) , .ZN( u2_uk_n437 ) );
  OAI22_X1 u2_uk_U817 (.ZN( u2_K16_20 ) , .B2( u2_uk_n1222 ) , .A2( u2_uk_n1229 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U818 (.B1( decrypt ) , .ZN( u2_K15_20 ) , .A2( u2_uk_n1815 ) , .B2( u2_uk_n1844 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U819 (.ZN( u2_K8_20 ) , .B2( u2_uk_n1521 ) , .A2( u2_uk_n1527 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U82 (.ZN( u2_K11_41 ) , .B2( u2_uk_n1672 ) , .B1( u2_uk_n214 ) , .A( u2_uk_n382 ) );
  AOI22_X1 u2_uk_U821 (.B2( u2_uk_K_r7_39 ) , .A2( u2_uk_K_r7_46 ) , .B1( u2_uk_n110 ) , .ZN( u2_uk_n1123 ) , .A1( u2_uk_n163 ) );
  AOI22_X1 u2_uk_U827 (.A1( decrypt ) , .B2( u2_uk_K_r5_18 ) , .A2( u2_uk_K_r5_53 ) , .ZN( u2_uk_n1079 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U828 (.ZN( u2_K8_6 ) , .B2( u2_uk_n1514 ) , .A2( u2_uk_n1519 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U829 (.A1( decrypt ) , .ZN( u2_K11_6 ) , .B2( u2_uk_n1669 ) , .A2( u2_uk_n1675 ) , .B1( u2_uk_n209 ) );
  NAND2_X1 u2_uk_U83 (.A1( u2_uk_K_r9_31 ) , .A2( u2_uk_n203 ) , .ZN( u2_uk_n382 ) );
  OAI22_X1 u2_uk_U830 (.ZN( u2_K2_6 ) , .B2( u2_uk_n1249 ) , .A2( u2_uk_n1270 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U831 (.ZN( u2_K12_3 ) , .A( u2_uk_n500 ) );
  AOI22_X1 u2_uk_U832 (.B1( decrypt ) , .B2( u2_uk_K_r10_18 ) , .A2( u2_uk_K_r10_27 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n500 ) );
  OAI21_X1 u2_uk_U833 (.B1( decrypt ) , .ZN( u2_K13_3 ) , .B2( u2_uk_n1751 ) , .A( u2_uk_n672 ) );
  NAND2_X1 u2_uk_U834 (.A1( u2_uk_K_r11_4 ) , .A2( u2_uk_n128 ) , .ZN( u2_uk_n672 ) );
  OAI22_X1 u2_uk_U835 (.B1( decrypt ) , .ZN( u2_K5_3 ) , .B2( u2_uk_n1374 ) , .A2( u2_uk_n1381 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U836 (.ZN( u2_K2_3 ) , .B2( u2_uk_n1239 ) , .A2( u2_uk_n1254 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U837 (.ZN( u2_K11_3 ) , .B2( u2_uk_n1639 ) , .A2( u2_uk_n1657 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U838 (.ZN( u2_K1_6 ) , .B2( u2_uk_n1168 ) , .A2( u2_uk_n1175 ) , .B1( u2_uk_n145 ) , .A1( u2_uk_n94 ) );
  INV_X1 u2_uk_U839 (.A( u2_key_r_41 ) , .ZN( u2_uk_n1175 ) );
  OAI21_X1 u2_uk_U84 (.B1( decrypt ) , .ZN( u2_K8_41 ) , .A( u2_uk_n1111 ) , .B2( u2_uk_n1517 ) );
  OAI21_X1 u2_uk_U840 (.B1( decrypt ) , .ZN( u2_K5_6 ) , .A( u2_uk_n1056 ) , .B2( u2_uk_n1387 ) );
  NAND2_X1 u2_uk_U841 (.A1( u2_uk_K_r3_10 ) , .ZN( u2_uk_n1056 ) , .A2( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U842 (.A1( decrypt ) , .ZN( u2_K7_3 ) , .B2( u2_uk_n1465 ) , .A2( u2_uk_n1487 ) , .B1( u2_uk_n187 ) );
  OAI22_X1 u2_uk_U843 (.B1( decrypt ) , .ZN( u2_K1_43 ) , .A2( u2_uk_n1149 ) , .B2( u2_uk_n1152 ) , .A1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U844 (.ZN( u2_K1_1 ) , .A1( u2_uk_n11 ) , .B2( u2_uk_n1174 ) , .A2( u2_uk_n1179 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U846 (.ZN( u2_K14_22 ) , .A1( u2_uk_n162 ) , .B2( u2_uk_n1772 ) , .A2( u2_uk_n1810 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U847 (.ZN( u2_K10_5 ) , .B2( u2_uk_n1595 ) , .A2( u2_uk_n1612 ) , .A1( u2_uk_n231 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U848 (.B1( decrypt ) , .ZN( u2_K5_41 ) , .B2( u2_uk_n1388 ) , .A2( u2_uk_n1396 ) , .A1( u2_uk_n145 ) );
  OAI22_X1 u2_uk_U849 (.ZN( u2_K15_22 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1828 ) , .A2( u2_uk_n1842 ) );
  NAND2_X1 u2_uk_U85 (.A2( decrypt ) , .A1( u2_uk_K_r6_30 ) , .ZN( u2_uk_n1111 ) );
  OAI22_X1 u2_uk_U850 (.B1( decrypt ) , .ZN( u2_K6_22 ) , .B2( u2_uk_n1417 ) , .A2( u2_uk_n1422 ) , .A1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U851 (.B1( decrypt ) , .ZN( u2_K15_23 ) , .B2( u2_uk_n1833 ) , .A2( u2_uk_n1851 ) , .A1( u2_uk_n207 ) );
  OAI22_X1 u2_uk_U852 (.ZN( u2_K14_23 ) , .A1( u2_uk_n163 ) , .A2( u2_uk_n1772 ) , .B2( u2_uk_n1779 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U853 (.B1( decrypt ) , .ZN( u2_K5_23 ) , .B2( u2_uk_n1385 ) , .A2( u2_uk_n1394 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U854 (.B1( decrypt ) , .ZN( u2_K13_34 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1738 ) , .A2( u2_uk_n1754 ) );
  OAI22_X1 u2_uk_U855 (.B1( decrypt ) , .ZN( u2_K5_34 ) , .A2( u2_uk_n1371 ) , .B2( u2_uk_n1384 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U856 (.B1( decrypt ) , .ZN( u2_K3_47 ) , .B2( u2_uk_n1297 ) , .A2( u2_uk_n1305 ) , .A1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U857 (.B1( decrypt ) , .ZN( u2_K8_5 ) , .B2( u2_uk_n1534 ) , .A2( u2_uk_n1540 ) , .A1( u2_uk_n231 ) );
  INV_X1 u2_uk_U86 (.ZN( u2_K2_41 ) , .A( u2_uk_n1001 ) );
  OAI22_X1 u2_uk_U861 (.ZN( u2_K7_10 ) , .B2( u2_uk_n1457 ) , .A2( u2_uk_n1487 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U864 (.ZN( u2_K15_45 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1837 ) , .A2( u2_uk_n1855 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U865 (.B1( decrypt ) , .ZN( u2_K13_45 ) , .B2( u2_uk_n1725 ) , .A2( u2_uk_n1763 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U866 (.ZN( u2_K12_43 ) , .B2( u2_uk_n1687 ) , .A2( u2_uk_n1707 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U867 (.ZN( u2_K6_45 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1424 ) , .A2( u2_uk_n1429 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U868 (.B1( decrypt ) , .ZN( u2_K3_30 ) , .B2( u2_uk_n1288 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1314 ) );
  OAI22_X1 u2_uk_U869 (.ZN( u2_K15_3 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1822 ) , .A2( u2_uk_n1838 ) , .A1( u2_uk_n231 ) );
  AOI22_X1 u2_uk_U87 (.B1( decrypt ) , .B2( u2_uk_K_r0_28 ) , .A2( u2_uk_K_r0_49 ) , .ZN( u2_uk_n1001 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U870 (.ZN( u2_K8_1 ) , .A2( u2_uk_n1502 ) , .B2( u2_uk_n1518 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U871 (.ZN( u2_K10_3 ) , .A1( u2_uk_n148 ) , .B2( u2_uk_n1603 ) , .A2( u2_uk_n1623 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U872 (.B1( decrypt ) , .ZN( u2_K9_3 ) , .A2( u2_uk_n1543 ) , .B2( u2_uk_n1547 ) , .A1( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U876 (.ZN( u2_K14_7 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1786 ) , .A2( u2_uk_n1805 ) );
  OAI22_X1 u2_uk_U877 (.ZN( u2_K13_24 ) , .B2( u2_uk_n1726 ) , .A2( u2_uk_n1767 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U878 (.B1( decrypt ) , .ZN( u2_K6_24 ) , .B2( u2_uk_n1427 ) , .A2( u2_uk_n1431 ) , .A1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U879 (.B1( decrypt ) , .ZN( u2_K15_13 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1814 ) , .B2( u2_uk_n1842 ) );
  OAI22_X1 u2_uk_U88 (.ZN( u2_K15_41 ) , .B1( u2_uk_n17 ) , .B2( u2_uk_n1835 ) , .A2( u2_uk_n1853 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U882 (.B1( decrypt ) , .ZN( u2_K5_19 ) , .A2( u2_uk_n1368 ) , .B2( u2_uk_n1405 ) , .A1( u2_uk_n203 ) );
  OAI22_X1 u2_uk_U883 (.B1( decrypt ) , .ZN( u2_K5_24 ) , .B2( u2_uk_n1372 ) , .A2( u2_uk_n1397 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U884 (.ZN( u2_K2_24 ) , .A2( u2_uk_n1234 ) , .B2( u2_uk_n1249 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U885 (.ZN( u2_K16_21 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1197 ) , .A2( u2_uk_n1204 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U886 (.ZN( u2_K8_21 ) , .B2( u2_uk_n1522 ) , .A2( u2_uk_n1528 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U887 (.ZN( u2_K16_24 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1194 ) , .A2( u2_uk_n1199 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U888 (.ZN( u2_K7_30 ) , .B2( u2_uk_n1460 ) , .A2( u2_uk_n1491 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U889 (.B1( decrypt ) , .ZN( u2_K5_13 ) , .B2( u2_uk_n1375 ) , .A2( u2_uk_n1406 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U89 (.ZN( u2_K13_41 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1723 ) , .A2( u2_uk_n1738 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U890 (.B1( decrypt ) , .ZN( u2_K5_14 ) , .B2( u2_uk_n1373 ) , .A2( u2_uk_n1380 ) , .A1( u2_uk_n213 ) );
  OAI22_X1 u2_uk_U891 (.B1( decrypt ) , .ZN( u2_K4_14 ) , .B2( u2_uk_n1322 ) , .A2( u2_uk_n1348 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U892 (.B1( decrypt ) , .ZN( u2_K3_13 ) , .B2( u2_uk_n1289 ) , .A2( u2_uk_n1294 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U894 (.ZN( u2_K2_17 ) , .A2( u2_uk_n1231 ) , .B2( u2_uk_n1247 ) , .A1( u2_uk_n145 ) , .B1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U897 (.ZN( u2_K16_38 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1210 ) , .A2( u2_uk_n1217 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U898 (.ZN( u2_K8_38 ) , .B1( u2_uk_n118 ) , .B2( u2_uk_n1530 ) , .A2( u2_uk_n1536 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U901 (.ZN( u2_K6_39 ) , .A1( u2_uk_n129 ) , .A2( u2_uk_n1411 ) , .B2( u2_uk_n1430 ) , .B1( u2_uk_n60 ) );
  OAI22_X1 u2_uk_U902 (.B1( decrypt ) , .ZN( u2_K4_39 ) , .B2( u2_uk_n1321 ) , .A2( u2_uk_n1342 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U904 (.ZN( u2_K3_39 ) , .B1( u2_uk_n118 ) , .B2( u2_uk_n1308 ) , .A2( u2_uk_n1312 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U905 (.ZN( u2_K2_39 ) , .B1( u2_uk_n11 ) , .A2( u2_uk_n1236 ) , .B2( u2_uk_n1251 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U906 (.A1( decrypt ) , .ZN( u2_K14_18 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1788 ) , .A2( u2_uk_n1796 ) );
  OAI22_X1 u2_uk_U907 (.ZN( u2_K13_23 ) , .A1( u2_uk_n110 ) , .B2( u2_uk_n1737 ) , .A2( u2_uk_n1767 ) , .B1( u2_uk_n223 ) );
  OAI22_X1 u2_uk_U908 (.A1( decrypt ) , .ZN( u2_K9_23 ) , .B2( u2_uk_n1554 ) , .A2( u2_uk_n1562 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U909 (.ZN( u2_K9_47 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1576 ) , .A2( u2_uk_n1583 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U91 (.ZN( u2_K4_41 ) , .B2( u2_uk_n1319 ) , .A2( u2_uk_n1336 ) , .B1( u2_uk_n162 ) , .A1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U910 (.ZN( u2_K12_16 ) , .A2( u2_uk_n1681 ) , .B2( u2_uk_n1693 ) , .B1( u2_uk_n209 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U911 (.A1( decrypt ) , .ZN( u2_K11_16 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1662 ) , .A2( u2_uk_n1668 ) );
  OAI22_X1 u2_uk_U912 (.A1( decrypt ) , .ZN( u2_K11_48 ) , .B2( u2_uk_n1659 ) , .A2( u2_uk_n1666 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U915 (.A1( decrypt ) , .ZN( u2_K14_8 ) , .B1( u2_uk_n142 ) , .A2( u2_uk_n1771 ) , .B2( u2_uk_n1789 ) );
  OAI22_X1 u2_uk_U917 (.ZN( u2_K14_20 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1783 ) , .A2( u2_uk_n1789 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U918 (.A1( decrypt ) , .ZN( u2_K2_20 ) , .A2( u2_uk_n1233 ) , .B2( u2_uk_n1262 ) , .B1( u2_uk_n142 ) );
  OAI22_X1 u2_uk_U919 (.A1( decrypt ) , .ZN( u2_K14_14 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1804 ) , .A2( u2_uk_n1811 ) );
  OAI22_X1 u2_uk_U92 (.A1( decrypt ) , .ZN( u2_K16_5 ) , .A2( u2_uk_n1191 ) , .B2( u2_uk_n1194 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U920 (.ZN( u2_K11_24 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1652 ) , .A2( u2_uk_n1657 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U921 (.A1( decrypt ) , .ZN( u2_K8_24 ) , .B2( u2_uk_n1500 ) , .A2( u2_uk_n1540 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U922 (.ZN( u2_K16_46 ) , .B2( u2_uk_n1189 ) , .A2( u2_uk_n1223 ) , .B1( u2_uk_n217 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U924 (.ZN( u2_K14_47 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1790 ) , .A2( u2_uk_n1800 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U925 (.A1( decrypt ) , .ZN( u2_K10_46 ) , .B2( u2_uk_n1602 ) , .A2( u2_uk_n1611 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U926 (.A1( decrypt ) , .ZN( u2_K10_34 ) , .B2( u2_uk_n1588 ) , .A2( u2_uk_n1614 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U927 (.ZN( u2_K9_34 ) , .A1( u2_uk_n100 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1551 ) , .A2( u2_uk_n1558 ) );
  OAI22_X1 u2_uk_U929 (.ZN( u2_K13_4 ) , .B2( u2_uk_n1732 ) , .A2( u2_uk_n1737 ) , .B1( u2_uk_n187 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U93 (.A1( decrypt ) , .ZN( u2_K15_5 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1829 ) , .A2( u2_uk_n1832 ) );
  OAI22_X1 u2_uk_U931 (.ZN( u2_K4_48 ) , .A1( u2_uk_n109 ) , .A2( u2_uk_n1325 ) , .B2( u2_uk_n1353 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U932 (.A1( decrypt ) , .ZN( u2_K2_48 ) , .B2( u2_uk_n1241 ) , .A2( u2_uk_n1256 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U933 (.ZN( u2_K10_8 ) , .A2( u2_uk_n1591 ) , .B2( u2_uk_n1605 ) , .B1( u2_uk_n161 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U934 (.A1( decrypt ) , .ZN( u2_K13_8 ) , .B2( u2_uk_n1751 ) , .A2( u2_uk_n1757 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U935 (.A1( decrypt ) , .ZN( u2_K6_20 ) , .A2( u2_uk_n1409 ) , .B2( u2_uk_n1414 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U936 (.A1( decrypt ) , .ZN( u2_K11_18 ) , .B2( u2_uk_n1637 ) , .A2( u2_uk_n1643 ) , .B1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U937 (.ZN( u2_K4_19 ) , .B2( u2_uk_n1335 ) , .A2( u2_uk_n1347 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U94 (.ZN( u2_K14_5 ) , .B2( u2_uk_n1796 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n932 ) );
  OAI22_X1 u2_uk_U940 (.ZN( u2_K10_20 ) , .A1( u2_uk_n118 ) , .B2( u2_uk_n1599 ) , .A2( u2_uk_n1629 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U941 (.A1( decrypt ) , .ZN( u2_K14_16 ) , .B1( u2_uk_n141 ) , .A2( u2_uk_n1774 ) , .B2( u2_uk_n1812 ) );
  OAI22_X1 u2_uk_U942 (.A1( decrypt ) , .ZN( u2_K6_36 ) , .A2( u2_uk_n1411 ) , .B2( u2_uk_n1419 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U943 (.ZN( u2_K14_38 ) , .B1( u2_uk_n145 ) , .A2( u2_uk_n1777 ) , .B2( u2_uk_n1793 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U944 (.ZN( u2_K13_38 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1755 ) , .A2( u2_uk_n1761 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U945 (.ZN( u2_K2_38 ) , .B2( u2_uk_n1246 ) , .A2( u2_uk_n1265 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U946 (.A1( decrypt ) , .ZN( u2_K7_37 ) , .B2( u2_uk_n1469 ) , .A2( u2_uk_n1493 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U947 (.ZN( u2_K2_37 ) , .A2( u2_uk_n1237 ) , .B2( u2_uk_n1264 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U948 (.A1( decrypt ) , .ZN( u2_K9_40 ) , .B2( u2_uk_n1570 ) , .A2( u2_uk_n1576 ) , .B1( u2_uk_n188 ) );
  OAI22_X1 u2_uk_U949 (.ZN( u2_K5_40 ) , .B2( u2_uk_n1383 ) , .A2( u2_uk_n1400 ) , .B1( u2_uk_n146 ) , .A1( u2_uk_n92 ) );
  NAND2_X1 u2_uk_U95 (.A1( u2_uk_K_r12_10 ) , .A2( u2_uk_n223 ) , .ZN( u2_uk_n932 ) );
  OAI22_X1 u2_uk_U950 (.ZN( u2_K2_22 ) , .B2( u2_uk_n1243 ) , .A2( u2_uk_n1260 ) , .B1( u2_uk_n230 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U951 (.A1( decrypt ) , .ZN( u2_K11_45 ) , .B2( u2_uk_n1647 ) , .A2( u2_uk_n1654 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U952 (.A1( decrypt ) , .ZN( u2_K8_45 ) , .B2( u2_uk_n1498 ) , .A2( u2_uk_n1536 ) , .B1( u2_uk_n191 ) );
  OAI22_X1 u2_uk_U953 (.A1( decrypt ) , .ZN( u2_K7_45 ) , .B2( u2_uk_n1460 ) , .A2( u2_uk_n1477 ) , .B1( u2_uk_n222 ) );
  OAI22_X1 u2_uk_U955 (.ZN( u2_K4_45 ) , .A1( u2_uk_n102 ) , .B2( u2_uk_n1321 ) , .A2( u2_uk_n1360 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U956 (.A1( decrypt ) , .ZN( u2_K2_45 ) , .B2( u2_uk_n1252 ) , .A2( u2_uk_n1274 ) , .B1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U957 (.A1( decrypt ) , .ZN( u2_K6_3 ) , .B2( u2_uk_n1417 ) , .A2( u2_uk_n1431 ) , .B1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U958 (.ZN( u2_K8_7 ) , .A2( u2_uk_n1500 ) , .B2( u2_uk_n1506 ) , .B1( u2_uk_n164 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U959 (.A1( decrypt ) , .ZN( u2_K7_7 ) , .B2( u2_uk_n1466 ) , .B1( u2_uk_n148 ) , .A2( u2_uk_n1488 ) );
  OAI22_X1 u2_uk_U960 (.A1( decrypt ) , .ZN( u2_K3_7 ) , .B2( u2_uk_n1293 ) , .A2( u2_uk_n1311 ) , .B1( u2_uk_n230 ) );
  OAI22_X1 u2_uk_U961 (.A1( decrypt ) , .ZN( u2_K9_15 ) , .B2( u2_uk_n1547 ) , .A2( u2_uk_n1554 ) , .B1( u2_uk_n209 ) );
  OAI22_X1 u2_uk_U962 (.A1( decrypt ) , .ZN( u2_K6_15 ) , .B2( u2_uk_n1423 ) , .A2( u2_uk_n1435 ) , .B1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U963 (.A1( decrypt ) , .ZN( u2_K6_25 ) , .B2( u2_uk_n1424 ) , .A2( u2_uk_n1440 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U964 (.A1( decrypt ) , .ZN( u2_K14_25 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1770 ) , .A2( u2_uk_n1776 ) );
  OAI22_X1 u2_uk_U965 (.ZN( u2_K1_34 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1144 ) , .A2( u2_uk_n1149 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U967 (.ZN( u2_K1_3 ) , .B2( u2_uk_n1154 ) , .A2( u2_uk_n1161 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n207 ) );
  AOI22_X1 u2_uk_U969 (.B1( decrypt ) , .B2( u2_uk_K_r7_23 ) , .A2( u2_uk_K_r7_30 ) , .ZN( u2_uk_n1136 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U971 (.B1( decrypt ) , .B2( u2_uk_K_r10_28 ) , .A2( u2_uk_K_r10_9 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n503 ) );
  AOI22_X1 u2_uk_U973 (.B1( decrypt ) , .B2( u2_uk_K_r7_15 ) , .A2( u2_uk_K_r7_22 ) , .ZN( u2_uk_n1137 ) , .A1( u2_uk_n161 ) );
  AOI22_X1 u2_uk_U974 (.B2( u2_uk_K_r11_19 ) , .A2( u2_uk_K_r11_24 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n681 ) );
  OAI21_X1 u2_uk_U975 (.B1( decrypt ) , .ZN( u2_K4_22 ) , .A( u2_uk_n1025 ) , .B2( u2_uk_n1327 ) );
  NAND2_X1 u2_uk_U976 (.A2( decrypt ) , .A1( u2_uk_K_r2_47 ) , .ZN( u2_uk_n1025 ) );
  NAND2_X1 u2_uk_U978 (.A2( decrypt ) , .A1( u2_uk_K_r5_13 ) , .ZN( u2_uk_n1082 ) );
  OAI21_X1 u2_uk_U979 (.ZN( u2_K6_23 ) , .A( u2_uk_n1063 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1442 ) );
  NAND2_X1 u2_uk_U980 (.A2( decrypt ) , .A1( u2_uk_K_r4_27 ) , .ZN( u2_uk_n1063 ) );
  OAI21_X1 u2_uk_U981 (.B1( decrypt ) , .ZN( u2_K3_35 ) , .A( u2_uk_n1012 ) , .B2( u2_uk_n1278 ) );
  NAND2_X1 u2_uk_U982 (.A1( u2_uk_K_r1_7 ) , .ZN( u2_uk_n1012 ) , .A2( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U983 (.ZN( u2_K14_46 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1790 ) , .A( u2_uk_n931 ) );
  NAND2_X1 u2_uk_U984 (.A2( decrypt ) , .A1( u2_uk_K_r12_22 ) , .ZN( u2_uk_n931 ) );
  NAND2_X1 u2_uk_U986 (.A2( decrypt ) , .A1( u2_uk_K_r2_53 ) , .ZN( u2_uk_n1038 ) );
  OAI21_X1 u2_uk_U987 (.ZN( u2_K16_4 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1227 ) , .A( u2_uk_n965 ) );
  NAND2_X1 u2_uk_U988 (.A1( u2_uk_K_r14_3 ) , .A2( u2_uk_n92 ) , .ZN( u2_uk_n965 ) );
  OAI21_X1 u2_uk_U989 (.ZN( u2_K8_4 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1116 ) , .B2( u2_uk_n1507 ) );
  INV_X1 u2_uk_U99 (.ZN( u2_K11_5 ) , .A( u2_uk_n391 ) );
  NAND2_X1 u2_uk_U990 (.A2( decrypt ) , .A1( u2_uk_K_r6_19 ) , .ZN( u2_uk_n1116 ) );
  OAI21_X1 u2_uk_U991 (.ZN( u2_K5_4 ) , .A( u2_uk_n1055 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1381 ) );
  NAND2_X1 u2_uk_U992 (.A1( u2_uk_K_r3_4 ) , .ZN( u2_uk_n1055 ) , .A2( u2_uk_n63 ) );
  OAI21_X1 u2_uk_U993 (.ZN( u2_K3_5 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1018 ) , .B2( u2_uk_n1302 ) );
  NAND2_X1 u2_uk_U994 (.A2( decrypt ) , .A1( u2_uk_K_r1_10 ) , .ZN( u2_uk_n1018 ) );
  OAI21_X1 u2_uk_U999 (.ZN( u2_K1_13 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1184 ) , .A( u2_uk_n969 ) );
endmodule
