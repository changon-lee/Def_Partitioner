module aes_aes_die_6 ( sa03_0, sa03_1, sa03_2, sa03_3, sa03_6, sa03_7, sa33_0, sa33_1, sa33_2, 
       sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, us03_n446, us03_n447, us03_n667, us03_n697, 
       us03_n706, us03_n747, us03_n778, us03_n782, us03_n784, us03_n789, us03_n810, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa30_sr_0, 
        sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, us03_n445, us03_n450, 
        us03_n458, us03_n462 );
  input sa03_0, sa03_1, sa03_2, sa03_3, sa03_6, sa03_7, sa33_0, sa33_1, sa33_2, 
        sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, us03_n446, us03_n447, us03_n667, us03_n697, 
        us03_n706, us03_n747, us03_n778, us03_n782, us03_n784, us03_n789, us03_n810;
  output sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa30_sr_0, 
        sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, us03_n445, us03_n450, 
        us03_n458, us03_n462;
  wire us03_n438, us03_n440, us03_n441, us03_n442, us03_n443, us03_n444, us03_n448, us03_n449, us03_n451, 
       us03_n452, us03_n453, us03_n454, us03_n455, us03_n456, us03_n457, us03_n459, us03_n460, us03_n461, 
       us03_n464, us03_n465, us03_n466, us03_n467, us03_n468, us03_n469, us03_n470, us03_n471, us03_n472, 
       us03_n473, us03_n474, us03_n475, us03_n476, us03_n477, us03_n478, us03_n479, us03_n480, us03_n481, 
       us03_n482, us03_n483, us03_n484, us03_n485, us03_n486, us03_n487, us03_n488, us03_n489, us03_n490, 
       us03_n491, us03_n492, us03_n493, us03_n494, us03_n495, us03_n496, us03_n497, us03_n498, us03_n499, 
       us03_n500, us03_n501, us03_n502, us03_n503, us03_n504, us03_n505, us03_n506, us03_n507, us03_n508, 
       us03_n509, us03_n510, us03_n511, us03_n512, us03_n513, us03_n514, us03_n515, us03_n516, us03_n517, 
       us03_n518, us03_n519, us03_n520, us03_n521, us03_n522, us03_n523, us03_n524, us03_n525, us03_n526, 
       us03_n527, us03_n528, us03_n529, us03_n530, us03_n531, us03_n532, us03_n533, us03_n534, us03_n535, 
       us03_n536, us03_n537, us03_n538, us03_n539, us03_n540, us03_n541, us03_n542, us03_n543, us03_n544, 
       us03_n545, us03_n546, us03_n547, us03_n548, us03_n549, us03_n550, us03_n551, us03_n552, us03_n553, 
       us03_n554, us03_n555, us03_n556, us03_n557, us03_n558, us03_n559, us03_n560, us03_n561, us03_n562, 
       us03_n563, us03_n564, us03_n565, us03_n566, us03_n567, us03_n568, us03_n569, us03_n570, us03_n571, 
       us03_n572, us03_n573, us03_n574, us03_n575, us03_n576, us03_n577, us03_n578, us03_n579, us03_n580, 
       us03_n581, us03_n582, us03_n583, us03_n584, us03_n585, us03_n586, us03_n587, us03_n588, us03_n589, 
       us03_n590, us03_n591, us03_n592, us03_n593, us03_n594, us03_n595, us03_n596, us03_n597, us03_n598, 
       us03_n599, us03_n600, us03_n601, us03_n602, us03_n603, us03_n604, us03_n605, us03_n606, us03_n607, 
       us03_n608, us03_n609, us03_n610, us03_n611, us03_n612, us03_n613, us03_n614, us03_n615, us03_n616, 
       us03_n617, us03_n618, us03_n619, us03_n620, us03_n621, us03_n622, us03_n623, us03_n624, us03_n625, 
       us03_n626, us03_n627, us03_n628, us03_n629, us03_n630, us03_n631, us03_n632, us03_n633, us03_n634, 
       us03_n635, us03_n636, us03_n637, us03_n638, us03_n639, us03_n640, us03_n641, us03_n642, us03_n643, 
       us03_n644, us03_n645, us03_n646, us03_n647, us03_n648, us03_n649, us03_n650, us03_n651, us03_n652, 
       us03_n653, us03_n654, us03_n655, us03_n656, us03_n657, us03_n658, us03_n659, us03_n660, us03_n661, 
       us03_n662, us03_n663, us03_n664, us03_n665, us03_n666, us03_n668, us03_n669, us03_n670, us03_n671, 
       us03_n672, us03_n673, us03_n674, us03_n675, us03_n676, us03_n677, us03_n678, us03_n679, us03_n680, 
       us03_n681, us03_n682, us03_n683, us03_n684, us03_n685, us03_n686, us03_n687, us03_n688, us03_n689, 
       us03_n690, us03_n691, us03_n692, us03_n693, us03_n694, us03_n695, us03_n696, us03_n698, us03_n699, 
       us03_n700, us03_n701, us03_n702, us03_n703, us03_n704, us03_n705, us03_n707, us03_n708, us03_n709, 
       us03_n710, us03_n711, us03_n712, us03_n713, us03_n714, us03_n715, us03_n716, us03_n717, us03_n718, 
       us03_n719, us03_n720, us03_n721, us03_n722, us03_n723, us03_n724, us03_n725, us03_n726, us03_n727, 
       us03_n728, us03_n729, us03_n730, us03_n731, us03_n732, us03_n733, us03_n734, us03_n735, us03_n736, 
       us03_n737, us03_n738, us03_n739, us03_n740, us03_n741, us03_n742, us03_n743, us03_n744, us03_n745, 
       us03_n746, us03_n748, us03_n749, us03_n750, us03_n751, us03_n752, us03_n753, us03_n754, us03_n755, 
       us03_n756, us03_n757, us03_n758, us03_n759, us03_n760, us03_n761, us03_n762, us03_n763, us03_n764, 
       us03_n765, us03_n766, us03_n767, us03_n768, us03_n769, us03_n770, us03_n771, us03_n772, us03_n773, 
       us03_n774, us03_n775, us03_n776, us03_n777, us03_n779, us03_n780, us03_n781, us03_n783, us03_n785, 
       us03_n786, us03_n787, us03_n788, us03_n790, us03_n791, us03_n792, us03_n793, us03_n794, us03_n795, 
       us03_n796, us03_n797, us03_n798, us03_n799, us03_n800, us03_n801, us03_n802, us03_n803, us03_n804, 
       us03_n805, us03_n806, us03_n807, us03_n808, us03_n809, us03_n811, us03_n812, us03_n813, us03_n814, 
       us03_n815, us03_n816, us03_n817, us03_n818, us03_n819, us03_n820, us03_n821, us03_n822, us03_n823, 
       us03_n824, us03_n825, us03_n826, us03_n827, us03_n828, us03_n829, us03_n830, us03_n831, us03_n832, 
       us03_n833, us03_n834, us03_n835, us03_n836, us03_n837, us03_n838, us03_n839, us03_n840, us03_n841, 
       us03_n842, us03_n843, us03_n844, us03_n847, us03_n848, us03_n849, us03_n850, us03_n851, us03_n852, 
       us03_n853, us03_n854, us03_n855, us03_n856, us03_n857, us03_n858, us03_n859, us03_n860, us03_n861, 
       us03_n862, us03_n863, us03_n864, us03_n865, us03_n866, us03_n867, us03_n868, us03_n869, us03_n870, 
       us03_n871, us03_n872, us03_n873, us03_n874, us33_n438, us33_n439, us33_n440, us33_n441, us33_n442, 
       us33_n443, us33_n444, us33_n445, us33_n446, us33_n447, us33_n448, us33_n449, us33_n450, us33_n451, 
       us33_n452, us33_n453, us33_n454, us33_n455, us33_n456, us33_n457, us33_n458, us33_n459, us33_n460, 
       us33_n461, us33_n462, us33_n463, us33_n464, us33_n465, us33_n466, us33_n467, us33_n468, us33_n469, 
       us33_n470, us33_n471, us33_n472, us33_n473, us33_n474, us33_n475, us33_n476, us33_n477, us33_n478, 
       us33_n479, us33_n480, us33_n481, us33_n482, us33_n483, us33_n484, us33_n485, us33_n486, us33_n487, 
       us33_n488, us33_n489, us33_n490, us33_n491, us33_n492, us33_n493, us33_n494, us33_n495, us33_n496, 
       us33_n497, us33_n498, us33_n499, us33_n500, us33_n501, us33_n502, us33_n503, us33_n504, us33_n505, 
       us33_n506, us33_n507, us33_n508, us33_n509, us33_n510, us33_n511, us33_n512, us33_n513, us33_n514, 
       us33_n515, us33_n516, us33_n517, us33_n518, us33_n519, us33_n520, us33_n521, us33_n522, us33_n523, 
       us33_n524, us33_n525, us33_n526, us33_n527, us33_n528, us33_n529, us33_n530, us33_n531, us33_n532, 
       us33_n533, us33_n534, us33_n535, us33_n536, us33_n537, us33_n538, us33_n539, us33_n540, us33_n541, 
       us33_n542, us33_n543, us33_n544, us33_n545, us33_n546, us33_n547, us33_n548, us33_n549, us33_n550, 
       us33_n551, us33_n552, us33_n553, us33_n554, us33_n555, us33_n556, us33_n557, us33_n558, us33_n559, 
       us33_n560, us33_n561, us33_n562, us33_n563, us33_n564, us33_n565, us33_n566, us33_n567, us33_n568, 
       us33_n569, us33_n570, us33_n571, us33_n572, us33_n573, us33_n574, us33_n575, us33_n576, us33_n577, 
       us33_n578, us33_n579, us33_n580, us33_n581, us33_n582, us33_n583, us33_n584, us33_n585, us33_n586, 
       us33_n587, us33_n588, us33_n589, us33_n590, us33_n591, us33_n592, us33_n593, us33_n594, us33_n595, 
       us33_n596, us33_n597, us33_n598, us33_n599, us33_n600, us33_n601, us33_n602, us33_n603, us33_n604, 
       us33_n605, us33_n606, us33_n607, us33_n608, us33_n609, us33_n610, us33_n611, us33_n612, us33_n613, 
       us33_n614, us33_n615, us33_n616, us33_n617, us33_n618, us33_n619, us33_n620, us33_n621, us33_n622, 
       us33_n623, us33_n624, us33_n625, us33_n626, us33_n627, us33_n628, us33_n629, us33_n630, us33_n631, 
       us33_n632, us33_n633, us33_n634, us33_n635, us33_n636, us33_n637, us33_n638, us33_n639, us33_n640, 
       us33_n641, us33_n642, us33_n643, us33_n644, us33_n645, us33_n646, us33_n647, us33_n648, us33_n649, 
       us33_n650, us33_n651, us33_n652, us33_n653, us33_n654, us33_n655, us33_n656, us33_n657, us33_n658, 
       us33_n659, us33_n660, us33_n661, us33_n662, us33_n663, us33_n664, us33_n665, us33_n666, us33_n667, 
       us33_n668, us33_n669, us33_n670, us33_n671, us33_n672, us33_n673, us33_n674, us33_n675, us33_n676, 
       us33_n677, us33_n678, us33_n679, us33_n680, us33_n681, us33_n682, us33_n683, us33_n684, us33_n685, 
       us33_n686, us33_n687, us33_n688, us33_n689, us33_n690, us33_n691, us33_n692, us33_n693, us33_n694, 
       us33_n695, us33_n696, us33_n697, us33_n698, us33_n699, us33_n700, us33_n701, us33_n702, us33_n703, 
       us33_n704, us33_n705, us33_n706, us33_n707, us33_n708, us33_n709, us33_n710, us33_n711, us33_n712, 
       us33_n713, us33_n714, us33_n715, us33_n716, us33_n717, us33_n718, us33_n719, us33_n720, us33_n721, 
       us33_n722, us33_n723, us33_n724, us33_n725, us33_n726, us33_n727, us33_n728, us33_n729, us33_n730, 
       us33_n731, us33_n732, us33_n733, us33_n734, us33_n735, us33_n736, us33_n737, us33_n738, us33_n739, 
       us33_n740, us33_n741, us33_n742, us33_n743, us33_n744, us33_n745, us33_n746, us33_n747, us33_n748, 
       us33_n749, us33_n750, us33_n751, us33_n752, us33_n753, us33_n754, us33_n755, us33_n756, us33_n757, 
       us33_n758, us33_n759, us33_n760, us33_n761, us33_n762, us33_n763, us33_n764, us33_n765, us33_n766, 
       us33_n767, us33_n768, us33_n769, us33_n770, us33_n771, us33_n772, us33_n773, us33_n774, us33_n775, 
       us33_n776, us33_n777, us33_n778, us33_n779, us33_n780, us33_n781, us33_n782, us33_n783, us33_n784, 
       us33_n785, us33_n786, us33_n787, us33_n788, us33_n789, us33_n790, us33_n791, us33_n792, us33_n793, 
       us33_n794, us33_n795, us33_n796, us33_n797, us33_n798, us33_n799, us33_n800, us33_n801, us33_n802, 
       us33_n803, us33_n804, us33_n805, us33_n806, us33_n807, us33_n808, us33_n809, us33_n810, us33_n811, 
       us33_n812, us33_n813, us33_n814, us33_n815, us33_n816, us33_n817, us33_n818, us33_n819, us33_n820, 
       us33_n821, us33_n822, us33_n823, us33_n824, us33_n825, us33_n826, us33_n827, us33_n828, us33_n829, 
       us33_n830, us33_n831, us33_n832, us33_n833, us33_n834, us33_n835, us33_n836, us33_n837, us33_n838, 
       us33_n839, us33_n840, us33_n841, us33_n842, us33_n843, us33_n844, us33_n845, us33_n846, us33_n847, 
       us33_n848, us33_n849, us33_n850, us33_n851, us33_n852, us33_n853, us33_n854, us33_n855, us33_n856, 
       us33_n857, us33_n858, us33_n859, us33_n860, us33_n861, us33_n862, us33_n863, us33_n864, us33_n865, 
       us33_n866, us33_n867, us33_n868, us33_n869, us33_n870, us33_n871, us33_n872, us33_n873, us33_n874, 
       us33_n875,  us33_n876;
  INV_X1 us03_U10 (.A( us03_n678 ) , .ZN( us03_n838 ) );
  NOR4_X1 us03_U100 (.A4( us03_n607 ) , .A3( us03_n608 ) , .A2( us03_n609 ) , .A1( us03_n610 ) , .ZN( us03_n617 ) );
  NOR4_X1 us03_U101 (.A4( us03_n612 ) , .A3( us03_n613 ) , .A2( us03_n614 ) , .A1( us03_n615 ) , .ZN( us03_n616 ) );
  NOR2_X1 us03_U102 (.ZN( us03_n684 ) , .A1( us03_n829 ) , .A2( us03_n830 ) );
  NAND4_X1 us03_U103 (.A4( us03_n471 ) , .A3( us03_n472 ) , .A2( us03_n473 ) , .A1( us03_n474 ) , .ZN( us03_n676 ) );
  NOR4_X1 us03_U104 (.A4( us03_n468 ) , .ZN( us03_n474 ) , .A3( us03_n554 ) , .A1( us03_n733 ) , .A2( us03_n753 ) );
  NOR4_X1 us03_U105 (.ZN( us03_n473 ) , .A1( us03_n529 ) , .A3( us03_n566 ) , .A4( us03_n598 ) , .A2( us03_n640 ) );
  NOR4_X1 us03_U106 (.ZN( us03_n472 ) , .A1( us03_n504 ) , .A3( us03_n542 ) , .A2( us03_n581 ) , .A4( us03_n714 ) );
  NAND4_X1 us03_U107 (.ZN( sa03_sr_1 ) , .A4( us03_n593 ) , .A3( us03_n594 ) , .A2( us03_n595 ) , .A1( us03_n596 ) );
  AOI211_X1 us03_U108 (.B( us03_n587 ) , .A( us03_n588 ) , .ZN( us03_n594 ) , .C2( us03_n809 ) , .C1( us03_n831 ) );
  NOR4_X1 us03_U109 (.A4( us03_n589 ) , .A3( us03_n590 ) , .A2( us03_n591 ) , .A1( us03_n592 ) , .ZN( us03_n593 ) );
  NOR4_X1 us03_U11 (.A4( us03_n443 ) , .A3( us03_n444 ) , .A2( us03_n514 ) , .A1( us03_n539 ) , .ZN( us03_n704 ) );
  AOI211_X1 us03_U110 (.A( us03_n586 ) , .ZN( us03_n595 ) , .B( us03_n619 ) , .C1( us03_n843 ) , .C2( us03_n853 ) );
  NAND4_X1 us03_U111 (.ZN( sa03_sr_0 ) , .A4( us03_n499 ) , .A3( us03_n500 ) , .A2( us03_n501 ) , .A1( us03_n502 ) );
  NOR4_X1 us03_U112 (.A4( us03_n496 ) , .A3( us03_n497 ) , .A2( us03_n498 ) , .ZN( us03_n499 ) , .A1( us03_n525 ) );
  AOI221_X1 us03_U113 (.A( us03_n495 ) , .ZN( us03_n500 ) , .B2( us03_n841 ) , .C1( us03_n844 ) , .C2( us03_n858 ) , .B1( us03_n860 ) );
  AOI211_X1 us03_U114 (.A( us03_n494 ) , .ZN( us03_n501 ) , .B( us03_n800 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NAND4_X1 us03_U115 (.A4( us03_n689 ) , .A3( us03_n690 ) , .A1( us03_n691 ) , .ZN( us03_n774 ) , .A2( us03_n870 ) );
  INV_X1 us03_U116 (.A( us03_n677 ) , .ZN( us03_n870 ) );
  AOI221_X1 us03_U117 (.A( us03_n679 ) , .ZN( us03_n690 ) , .B2( us03_n838 ) , .C1( us03_n840 ) , .C2( us03_n860 ) , .B1( us03_n863 ) );
  NOR4_X1 us03_U118 (.A4( us03_n685 ) , .A3( us03_n686 ) , .A2( us03_n687 ) , .A1( us03_n688 ) , .ZN( us03_n689 ) );
  NOR2_X1 us03_U119 (.ZN( us03_n731 ) , .A2( us03_n830 ) , .A1( us03_n843 ) );
  OR3_X1 us03_U12 (.ZN( us03_n444 ) , .A1( us03_n526 ) , .A3( us03_n575 ) , .A2( us03_n873 ) );
  NAND4_X1 us03_U120 (.A4( us03_n717 ) , .A3( us03_n718 ) , .A2( us03_n719 ) , .ZN( us03_n739 ) , .A1( us03_n855 ) );
  INV_X1 us03_U121 (.A( us03_n707 ) , .ZN( us03_n855 ) );
  NOR4_X1 us03_U122 (.A4( us03_n713 ) , .A3( us03_n714 ) , .A2( us03_n715 ) , .A1( us03_n716 ) , .ZN( us03_n717 ) );
  AOI221_X1 us03_U123 (.A( us03_n708 ) , .ZN( us03_n719 ) , .C2( us03_n842 ) , .B2( us03_n843 ) , .C1( us03_n859 ) , .B1( us03_n860 ) );
  NOR2_X1 us03_U124 (.ZN( us03_n645 ) , .A1( us03_n852 ) , .A2( us03_n866 ) );
  NAND4_X1 us03_U125 (.A4( us03_n571 ) , .A3( us03_n572 ) , .A1( us03_n573 ) , .ZN( us03_n721 ) , .A2( us03_n872 ) );
  NOR4_X1 us03_U126 (.A4( us03_n567 ) , .A3( us03_n568 ) , .A2( us03_n569 ) , .A1( us03_n570 ) , .ZN( us03_n571 ) );
  AOI221_X1 us03_U127 (.A( us03_n562 ) , .C2( us03_n563 ) , .ZN( us03_n572 ) , .B2( us03_n843 ) , .B1( us03_n850 ) , .C1( us03_n851 ) );
  INV_X1 us03_U128 (.A( us03_n605 ) , .ZN( us03_n872 ) );
  NAND4_X1 us03_U129 (.A4( us03_n491 ) , .A3( us03_n492 ) , .A1( us03_n493 ) , .ZN( us03_n800 ) , .A2( us03_n865 ) );
  OR4_X1 us03_U13 (.A4( us03_n440 ) , .A2( us03_n441 ) , .A1( us03_n442 ) , .ZN( us03_n443 ) , .A3( us03_n551 ) );
  AOI221_X1 us03_U130 (.A( us03_n487 ) , .ZN( us03_n492 ) , .B2( us03_n834 ) , .C2( us03_n839 ) , .C1( us03_n849 ) , .B1( us03_n858 ) );
  INV_X1 us03_U131 (.A( us03_n776 ) , .ZN( us03_n865 ) );
  NOR2_X1 us03_U132 (.ZN( us03_n493 ) , .A1( us03_n676 ) , .A2( us03_n692 ) );
  INV_X1 us03_U133 (.A( us03_n760 ) , .ZN( us03_n828 ) );
  INV_X1 us03_U134 (.A( us03_n461 ) , .ZN( us03_n862 ) );
  OAI21_X1 us03_U135 (.ZN( us03_n461 ) , .B1( us03_n807 ) , .A( us03_n832 ) , .B2( us03_n849 ) );
  OR4_X1 us03_U136 (.A4( us03_n578 ) , .A3( us03_n579 ) , .A2( us03_n580 ) , .A1( us03_n581 ) , .ZN( us03_n582 ) );
  OR4_X1 us03_U137 (.A4( us03_n564 ) , .A3( us03_n565 ) , .A2( us03_n566 ) , .ZN( us03_n570 ) , .A1( us03_n663 ) );
  OR4_X1 us03_U138 (.A4( us03_n516 ) , .A2( us03_n517 ) , .A1( us03_n518 ) , .ZN( us03_n520 ) , .A3( us03_n819 ) );
  OR4_X1 us03_U139 (.A4( us03_n680 ) , .A3( us03_n681 ) , .A2( us03_n682 ) , .A1( us03_n683 ) , .ZN( us03_n688 ) );
  INV_X1 us03_U14 (.A( us03_n611 ) , .ZN( us03_n873 ) );
  OR4_X1 us03_U140 (.ZN( us03_n464 ) , .A4( us03_n516 ) , .A3( us03_n527 ) , .A2( us03_n576 ) , .A1( us03_n710 ) );
  NAND2_X1 us03_U141 (.ZN( us03_n611 ) , .A2( us03_n835 ) , .A1( us03_n871 ) );
  OR3_X1 us03_U142 (.A3( us03_n504 ) , .A2( us03_n505 ) , .A1( us03_n506 ) , .ZN( us03_n509 ) );
  AOI221_X1 us03_U143 (.A( us03_n711 ) , .B2( us03_n712 ) , .ZN( us03_n718 ) , .C1( us03_n830 ) , .B1( us03_n837 ) , .C2( us03_n861 ) );
  OR2_X1 us03_U144 (.A2( us03_n709 ) , .A1( us03_n710 ) , .ZN( us03_n711 ) );
  INV_X1 us03_U145 (.A( us03_n752 ) , .ZN( us03_n867 ) );
  OAI21_X1 us03_U146 (.B1( us03_n751 ) , .ZN( us03_n752 ) , .A( us03_n843 ) , .B2( us03_n866 ) );
  INV_X1 us03_U147 (.A( us03_n670 ) , .ZN( us03_n857 ) );
  AOI21_X1 us03_U148 (.A( us03_n668 ) , .B1( us03_n669 ) , .ZN( us03_n670 ) , .B2( us03_n854 ) );
  AOI222_X1 us03_U149 (.ZN( us03_n658 ) , .A2( us03_n837 ) , .B1( us03_n839 ) , .C2( us03_n843 ) , .A1( us03_n858 ) , .C1( us03_n861 ) , .B2( us03_n868 ) );
  INV_X1 us03_U15 (.A( us03_n747 ) , .ZN( us03_n861 ) );
  INV_X1 us03_U150 (.A( us03_n645 ) , .ZN( us03_n868 ) );
  OAI22_X1 us03_U151 (.ZN( us03_n481 ) , .A1( us03_n706 ) , .B2( us03_n783 ) , .A2( us03_n804 ) , .B1( us03_n810 ) );
  OAI222_X1 us03_U153 (.B2( us03_n745 ) , .B1( us03_n746 ) , .A2( us03_n747 ) , .ZN( us03_n755 ) , .C2( us03_n803 ) , .C1( us03_n812 ) , .A1( us03_n815 ) );
  OAI222_X1 us03_U154 (.B2( us03_n706 ) , .ZN( us03_n707 ) , .C2( us03_n722 ) , .B1( us03_n745 ) , .A1( us03_n804 ) , .C1( us03_n812 ) , .A2( us03_n813 ) );
  OAI222_X1 us03_U155 (.ZN( us03_n615 ) , .B1( us03_n695 ) , .C1( us03_n722 ) , .C2( us03_n745 ) , .B2( us03_n784 ) , .A2( us03_n790 ) , .A1( us03_n814 ) );
  OAI222_X1 us03_U156 (.ZN( us03_n503 ) , .C2( us03_n623 ) , .B2( us03_n645 ) , .B1( us03_n745 ) , .A2( us03_n746 ) , .C1( us03_n803 ) , .A1( us03_n804 ) );
  AOI22_X1 us03_U157 (.ZN( us03_n694 ) , .A1( us03_n828 ) , .B2( us03_n841 ) , .A2( us03_n863 ) , .B1( us03_n866 ) );
  INV_X1 us03_U158 (.A( us03_n728 ) , .ZN( us03_n837 ) );
  AOI221_X1 us03_U159 (.A( us03_n762 ) , .ZN( us03_n772 ) , .C2( us03_n808 ) , .B2( us03_n833 ) , .C1( us03_n853 ) , .B1( us03_n864 ) );
  AOI222_X1 us03_U16 (.ZN( us03_n561 ) , .B1( us03_n828 ) , .C1( us03_n839 ) , .A2( us03_n841 ) , .A1( us03_n852 ) , .B2( us03_n861 ) , .C2( us03_n871 ) );
  AOI21_X1 us03_U160 (.B2( us03_n761 ) , .ZN( us03_n762 ) , .A( us03_n786 ) , .B1( us03_n790 ) );
  INV_X1 us03_U161 (.A( us03_n759 ) , .ZN( us03_n833 ) );
  NAND2_X1 us03_U162 (.A1( us03_n449 ) , .A2( us03_n451 ) , .ZN( us03_n760 ) );
  INV_X1 us03_U163 (.A( us03_n788 ) , .ZN( us03_n830 ) );
  OAI22_X1 us03_U164 (.ZN( us03_n635 ) , .A1( us03_n697 ) , .B2( us03_n726 ) , .A2( us03_n760 ) , .B1( us03_n814 ) );
  OAI221_X1 us03_U165 (.A( us03_n725 ) , .C2( us03_n726 ) , .B2( us03_n727 ) , .B1( us03_n728 ) , .ZN( us03_n735 ) , .C1( us03_n815 ) );
  AOI22_X1 us03_U166 (.ZN( us03_n725 ) , .B1( us03_n830 ) , .A2( us03_n836 ) , .A1( us03_n861 ) , .B2( us03_n864 ) );
  OAI22_X1 us03_U167 (.ZN( us03_n487 ) , .A1( us03_n722 ) , .B2( us03_n726 ) , .B1( us03_n728 ) , .A2( us03_n777 ) );
  OAI22_X1 us03_U168 (.ZN( us03_n622 ) , .B1( us03_n667 ) , .B2( us03_n745 ) , .A1( us03_n813 ) , .A2( us03_n814 ) );
  OAI22_X1 us03_U169 (.A1( us03_n722 ) , .ZN( us03_n724 ) , .B2( us03_n748 ) , .B1( us03_n810 ) , .A2( us03_n814 ) );
  NOR4_X1 us03_U17 (.ZN( us03_n471 ) , .A2( us03_n519 ) , .A4( us03_n592 ) , .A1( us03_n607 ) , .A3( us03_n627 ) );
  OAI22_X1 us03_U170 (.B2( us03_n777 ) , .B1( us03_n778 ) , .ZN( us03_n779 ) , .A2( us03_n812 ) , .A1( us03_n813 ) );
  OAI22_X1 us03_U171 (.B2( us03_n742 ) , .ZN( us03_n744 ) , .A2( us03_n760 ) , .B1( us03_n778 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U172 (.B2( us03_n801 ) , .B1( us03_n802 ) , .A2( us03_n803 ) , .A1( us03_n804 ) , .ZN( us03_n806 ) );
  OAI22_X1 us03_U173 (.ZN( us03_n494 ) , .A2( us03_n742 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n804 ) );
  INV_X1 us03_U174 (.A( us03_n742 ) , .ZN( us03_n835 ) );
  INV_X1 us03_U175 (.A( us03_n814 ) , .ZN( us03_n829 ) );
  INV_X1 us03_U176 (.A( us03_n786 ) , .ZN( us03_n843 ) );
  INV_X1 us03_U177 (.A( us03_n812 ) , .ZN( us03_n831 ) );
  OAI22_X1 us03_U178 (.ZN( us03_n588 ) , .B1( us03_n728 ) , .B2( us03_n747 ) , .A2( us03_n784 ) , .A1( us03_n801 ) );
  OAI22_X1 us03_U179 (.ZN( us03_n693 ) , .A2( us03_n728 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n815 ) );
  NOR4_X1 us03_U18 (.ZN( us03_n477 ) , .A1( us03_n518 ) , .A4( us03_n555 ) , .A3( us03_n580 ) , .A2( us03_n628 ) );
  OAI22_X1 us03_U180 (.ZN( us03_n708 ) , .A2( us03_n726 ) , .B2( us03_n727 ) , .A1( us03_n742 ) , .B1( us03_n811 ) );
  INV_X1 us03_U181 (.A( us03_n667 ) , .ZN( us03_n863 ) );
  NOR2_X1 us03_U182 (.A1( us03_n695 ) , .ZN( us03_n768 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U183 (.ZN( us03_n664 ) , .A1( us03_n726 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U184 (.ZN( us03_n592 ) , .A2( us03_n695 ) , .A1( us03_n726 ) );
  NOR2_X1 us03_U185 (.ZN( us03_n568 ) , .A1( us03_n726 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U186 (.ZN( us03_n716 ) , .A2( us03_n722 ) , .A1( us03_n742 ) );
  NOR2_X1 us03_U187 (.ZN( us03_n544 ) , .A2( us03_n778 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U188 (.ZN( us03_n575 ) , .A2( us03_n697 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U189 (.ZN( us03_n652 ) , .A1( us03_n726 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U19 (.A4( us03_n530 ) , .A3( us03_n531 ) , .A2( us03_n532 ) , .ZN( us03_n533 ) , .A1( us03_n818 ) );
  NOR2_X1 us03_U190 (.ZN( us03_n610 ) , .A1( us03_n777 ) , .A2( us03_n784 ) );
  INV_X1 us03_U191 (.A( us03_n748 ) , .ZN( us03_n840 ) );
  NOR2_X1 us03_U192 (.ZN( us03_n530 ) , .A2( us03_n747 ) , .A1( us03_n748 ) );
  NOR2_X1 us03_U193 (.ZN( us03_n627 ) , .A2( us03_n726 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U194 (.ZN( us03_n613 ) , .A1( us03_n783 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U195 (.ZN( us03_n599 ) , .A2( us03_n778 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U196 (.ZN( us03_n609 ) , .A2( us03_n778 ) , .A1( us03_n804 ) );
  INV_X1 us03_U197 (.A( us03_n745 ) , .ZN( us03_n832 ) );
  NOR2_X1 us03_U198 (.A2( us03_n742 ) , .ZN( us03_n767 ) , .A1( us03_n810 ) );
  NOR2_X1 us03_U199 (.ZN( us03_n526 ) , .A2( us03_n722 ) , .A1( us03_n801 ) );
  NOR4_X1 us03_U20 (.ZN( us03_n454 ) , .A2( us03_n515 ) , .A1( us03_n541 ) , .A3( us03_n577 ) , .A4( us03_n613 ) );
  NOR2_X1 us03_U200 (.ZN( us03_n529 ) , .A2( us03_n778 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U201 (.ZN( us03_n626 ) , .A2( us03_n667 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U202 (.ZN( us03_n597 ) , .A2( us03_n789 ) , .A1( us03_n814 ) );
  INV_X1 us03_U203 (.A( us03_n790 ) , .ZN( us03_n849 ) );
  NOR2_X1 us03_U204 (.ZN( us03_n650 ) , .A1( us03_n667 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U205 (.A1( us03_n667 ) , .ZN( us03_n671 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U206 (.ZN( us03_n600 ) , .A1( us03_n667 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U207 (.A1( us03_n667 ) , .ZN( us03_n686 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U208 (.A2( us03_n706 ) , .A1( us03_n748 ) , .ZN( us03_n769 ) );
  NOR2_X1 us03_U209 (.A1( us03_n667 ) , .ZN( us03_n764 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U21 (.A4( us03_n539 ) , .A3( us03_n540 ) , .A2( us03_n541 ) , .ZN( us03_n548 ) , .A1( us03_n686 ) );
  NOR2_X1 us03_U210 (.A1( us03_n697 ) , .ZN( us03_n766 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U211 (.ZN( us03_n539 ) , .A2( us03_n695 ) , .A1( us03_n697 ) );
  NOR2_X1 us03_U212 (.ZN( us03_n525 ) , .A1( us03_n667 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U213 (.ZN( us03_n665 ) , .A1( us03_n748 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U214 (.ZN( us03_n553 ) , .A1( us03_n748 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U215 (.ZN( us03_n506 ) , .A2( us03_n778 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U216 (.ZN( us03_n541 ) , .A2( us03_n706 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U217 (.ZN( us03_n662 ) , .A1( us03_n783 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U218 (.A2( us03_n695 ) , .ZN( us03_n714 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U219 (.B1( us03_n438 ) , .ZN( us03_n442 ) , .A2( us03_n726 ) , .A1( us03_n742 ) , .B2( us03_n747 ) );
  NOR2_X1 us03_U22 (.ZN( us03_n678 ) , .A2( us03_n832 ) , .A1( us03_n837 ) );
  NOR3_X1 us03_U220 (.ZN( us03_n438 ) , .A2( us03_n834 ) , .A3( us03_n835 ) , .A1( us03_n844 ) );
  NOR2_X1 us03_U221 (.ZN( us03_n505 ) , .A1( us03_n810 ) , .A2( us03_n815 ) );
  INV_X1 us03_U222 (.A( us03_n804 ) , .ZN( us03_n839 ) );
  NOR2_X1 us03_U223 (.ZN( us03_n659 ) , .A1( us03_n727 ) , .A2( us03_n788 ) );
  NOR2_X1 us03_U224 (.ZN( us03_n660 ) , .A2( us03_n695 ) , .A1( us03_n727 ) );
  NOR2_X1 us03_U225 (.ZN( us03_n555 ) , .A1( us03_n790 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U226 (.ZN( us03_n543 ) , .A1( us03_n747 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U227 (.ZN( us03_n507 ) , .A1( us03_n727 ) , .A2( us03_n777 ) );
  INV_X1 us03_U228 (.A( us03_n801 ) , .ZN( us03_n841 ) );
  NOR2_X1 us03_U229 (.A2( us03_n695 ) , .A1( us03_n778 ) , .ZN( us03_n818 ) );
  NOR4_X1 us03_U23 (.A4( us03_n512 ) , .A3( us03_n513 ) , .A2( us03_n514 ) , .A1( us03_n515 ) , .ZN( us03_n522 ) );
  NOR2_X1 us03_U230 (.ZN( us03_n528 ) , .A2( us03_n742 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U231 (.B2( us03_n748 ) , .B1( us03_n749 ) , .A1( us03_n750 ) , .ZN( us03_n754 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U232 (.ZN( us03_n749 ) , .A2( us03_n850 ) , .A1( us03_n858 ) );
  NOR3_X1 us03_U233 (.ZN( us03_n750 ) , .A2( us03_n851 ) , .A1( us03_n861 ) , .A3( us03_n863 ) );
  NOR2_X1 us03_U234 (.A1( us03_n747 ) , .ZN( us03_n765 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U235 (.A2( us03_n742 ) , .ZN( us03_n753 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U236 (.ZN( us03_n542 ) , .A2( us03_n783 ) , .A1( us03_n790 ) );
  NOR2_X1 us03_U237 (.ZN( us03_n661 ) , .A1( us03_n727 ) , .A2( us03_n783 ) );
  INV_X1 us03_U238 (.A( us03_n726 ) , .ZN( us03_n850 ) );
  NOR2_X1 us03_U239 (.ZN( us03_n629 ) , .A1( us03_n722 ) , .A2( us03_n811 ) );
  AOI222_X1 us03_U24 (.ZN( us03_n523 ) , .A1( us03_n832 ) , .B2( us03_n835 ) , .C1( us03_n842 ) , .C2( us03_n848 ) , .A2( us03_n850 ) , .B1( us03_n864 ) );
  NOR2_X1 us03_U240 (.ZN( us03_n733 ) , .A2( us03_n801 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U241 (.ZN( us03_n612 ) , .A1( us03_n760 ) , .A2( us03_n810 ) );
  NOR4_X1 us03_U242 (.A2( us03_n489 ) , .A1( us03_n490 ) , .ZN( us03_n491 ) , .A3( us03_n578 ) , .A4( us03_n610 ) );
  OR4_X1 us03_U243 (.ZN( us03_n490 ) , .A4( us03_n532 ) , .A2( us03_n545 ) , .A1( us03_n557 ) , .A3( us03_n630 ) );
  OAI22_X1 us03_U244 (.B1( us03_n488 ) , .ZN( us03_n489 ) , .A1( us03_n684 ) , .A2( us03_n761 ) , .B2( us03_n815 ) );
  NOR3_X1 us03_U245 (.ZN( us03_n488 ) , .A1( us03_n780 ) , .A2( us03_n848 ) , .A3( us03_n861 ) );
  NOR2_X1 us03_U246 (.ZN( us03_n504 ) , .A2( us03_n726 ) , .A1( us03_n760 ) );
  NOR2_X1 us03_U247 (.ZN( us03_n514 ) , .A1( us03_n706 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U248 (.ZN( us03_n715 ) , .A2( us03_n742 ) , .A1( us03_n784 ) );
  NOR2_X1 us03_U249 (.ZN( us03_n552 ) , .A1( us03_n784 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U25 (.A3( us03_n519 ) , .A1( us03_n520 ) , .ZN( us03_n521 ) , .A2( us03_n671 ) , .A4( us03_n767 ) );
  NOR2_X1 us03_U250 (.ZN( us03_n515 ) , .A1( us03_n706 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U251 (.ZN( us03_n556 ) , .A1( us03_n706 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U252 (.ZN( us03_n519 ) , .A1( us03_n788 ) , .A2( us03_n810 ) );
  INV_X1 us03_U253 (.A( us03_n803 ) , .ZN( us03_n858 ) );
  NOR2_X1 us03_U254 (.ZN( us03_n628 ) , .A1( us03_n745 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U255 (.ZN( us03_n713 ) , .A1( us03_n803 ) , .A2( us03_n815 ) );
  AOI21_X1 us03_U256 (.ZN( us03_n569 ) , .B2( us03_n695 ) , .B1( us03_n804 ) , .A( us03_n810 ) );
  NOR2_X1 us03_U257 (.ZN( us03_n653 ) , .A1( us03_n788 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U258 (.ZN( us03_n666 ) , .A2( us03_n706 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U259 (.ZN( us03_n654 ) , .A1( us03_n745 ) , .A2( us03_n778 ) );
  AOI222_X1 us03_U26 (.B2( us03_n636 ) , .ZN( us03_n642 ) , .B1( us03_n839 ) , .A1( us03_n840 ) , .C2( us03_n844 ) , .C1( us03_n861 ) , .A2( us03_n863 ) );
  NOR2_X1 us03_U260 (.ZN( us03_n554 ) , .A1( us03_n760 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U261 (.ZN( us03_n540 ) , .A1( us03_n760 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U262 (.ZN( us03_n699 ) , .A2( us03_n784 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U263 (.ZN( us03_n607 ) , .A2( us03_n722 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U264 (.A1( us03_n728 ) , .ZN( us03_n763 ) , .A2( us03_n784 ) );
  AOI21_X1 us03_U265 (.A( us03_n813 ) , .B2( us03_n814 ) , .B1( us03_n815 ) , .ZN( us03_n816 ) );
  NOR2_X1 us03_U266 (.ZN( us03_n577 ) , .A2( us03_n706 ) , .A1( us03_n728 ) );
  NOR2_X1 us03_U267 (.ZN( us03_n531 ) , .A2( us03_n722 ) , .A1( us03_n728 ) );
  AOI21_X1 us03_U268 (.B1( us03_n623 ) , .ZN( us03_n625 ) , .A( us03_n761 ) , .B2( us03_n812 ) );
  AOI21_X1 us03_U269 (.A( us03_n810 ) , .B2( us03_n811 ) , .B1( us03_n812 ) , .ZN( us03_n817 ) );
  NOR4_X1 us03_U27 (.A4( us03_n637 ) , .A3( us03_n638 ) , .A2( us03_n639 ) , .A1( us03_n640 ) , .ZN( us03_n641 ) );
  AOI21_X1 us03_U270 (.ZN( us03_n513 ) , .A( us03_n727 ) , .B1( us03_n748 ) , .B2( us03_n801 ) );
  AOI21_X1 us03_U271 (.ZN( us03_n497 ) , .B1( us03_n678 ) , .A( us03_n810 ) , .B2( us03_n814 ) );
  AOI21_X1 us03_U272 (.ZN( us03_n476 ) , .B2( us03_n695 ) , .A( us03_n747 ) , .B1( us03_n777 ) );
  NOR2_X1 us03_U273 (.ZN( us03_n580 ) , .A1( us03_n742 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U274 (.ZN( us03_n640 ) , .A2( us03_n786 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U275 (.ZN( us03_n591 ) , .B1( us03_n748 ) , .A( us03_n790 ) , .B2( us03_n811 ) );
  NOR2_X1 us03_U276 (.A2( us03_n706 ) , .A1( us03_n760 ) , .ZN( us03_n792 ) );
  AOI21_X1 us03_U277 (.ZN( us03_n624 ) , .B2( us03_n667 ) , .A( us03_n788 ) , .B1( us03_n789 ) );
  NOR2_X1 us03_U278 (.ZN( us03_n668 ) , .A1( us03_n788 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U279 (.ZN( us03_n518 ) , .A2( us03_n706 ) , .A1( us03_n812 ) );
  NOR3_X1 us03_U28 (.A2( us03_n605 ) , .A1( us03_n606 ) , .ZN( us03_n644 ) , .A3( us03_n720 ) );
  AOI21_X1 us03_U280 (.ZN( us03_n475 ) , .A( us03_n667 ) , .B1( us03_n748 ) , .B2( us03_n804 ) );
  NOR2_X1 us03_U281 (.ZN( us03_n557 ) , .A2( us03_n789 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U282 (.ZN( us03_n517 ) , .A2( us03_n697 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U283 (.ZN( us03_n681 ) , .A2( us03_n697 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U284 (.ZN( us03_n651 ) , .A1( us03_n760 ) , .A2( us03_n784 ) );
  INV_X1 us03_U285 (.A( us03_n811 ) , .ZN( us03_n834 ) );
  AOI21_X1 us03_U286 (.ZN( us03_n508 ) , .B2( us03_n667 ) , .A( us03_n728 ) , .B1( us03_n813 ) );
  AOI21_X1 us03_U287 (.ZN( us03_n537 ) , .B2( us03_n810 ) , .A( us03_n812 ) , .B1( us03_n813 ) );
  INV_X1 us03_U288 (.A( us03_n761 ) , .ZN( us03_n864 ) );
  AOI21_X1 us03_U289 (.ZN( us03_n538 ) , .A( us03_n761 ) , .B2( us03_n777 ) , .B1( us03_n815 ) );
  AOI221_X1 us03_U29 (.A( us03_n779 ) , .ZN( us03_n796 ) , .C2( us03_n835 ) , .B2( us03_n836 ) , .B1( us03_n863 ) , .C1( us03_n864 ) );
  NOR2_X1 us03_U290 (.ZN( us03_n579 ) , .A1( us03_n667 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U291 (.ZN( us03_n587 ) , .B2( us03_n697 ) , .B1( us03_n813 ) , .A( us03_n815 ) );
  AOI21_X1 us03_U292 (.B1( us03_n697 ) , .ZN( us03_n698 ) , .A( us03_n730 ) , .B2( us03_n761 ) );
  AOI21_X1 us03_U293 (.ZN( us03_n589 ) , .B2( us03_n761 ) , .A( us03_n783 ) , .B1( us03_n810 ) );
  AOI21_X1 us03_U294 (.ZN( us03_n496 ) , .A( us03_n722 ) , .B2( us03_n760 ) , .B1( us03_n812 ) );
  AOI21_X1 us03_U295 (.ZN( us03_n550 ) , .B1( us03_n667 ) , .A( us03_n695 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U296 (.ZN( us03_n545 ) , .A1( us03_n697 ) , .A2( us03_n742 ) );
  INV_X1 us03_U297 (.A( us03_n727 ) , .ZN( us03_n866 ) );
  INV_X1 us03_U298 (.A( us03_n789 ) , .ZN( us03_n871 ) );
  INV_X1 us03_U299 (.A( us03_n810 ) , .ZN( us03_n852 ) );
  NOR3_X1 us03_U3 (.ZN( us03_n596 ) , .A1( us03_n606 ) , .A3( us03_n721 ) , .A2( us03_n740 ) );
  NOR4_X1 us03_U30 (.A4( us03_n791 ) , .A3( us03_n792 ) , .A2( us03_n793 ) , .A1( us03_n794 ) , .ZN( us03_n795 ) );
  AOI21_X1 us03_U300 (.ZN( us03_n638 ) , .B2( us03_n745 ) , .A( us03_n790 ) , .B1( us03_n801 ) );
  AOI21_X1 us03_U301 (.ZN( us03_n647 ) , .B1( us03_n727 ) , .B2( us03_n761 ) , .A( us03_n811 ) );
  INV_X1 us03_U302 (.A( us03_n784 ) , .ZN( us03_n860 ) );
  NOR2_X1 us03_U303 (.ZN( us03_n683 ) , .A1( us03_n727 ) , .A2( us03_n814 ) );
  AOI21_X1 us03_U304 (.B1( us03_n684 ) , .ZN( us03_n685 ) , .A( us03_n726 ) , .B2( us03_n759 ) );
  AOI21_X1 us03_U305 (.ZN( us03_n567 ) , .B1( us03_n748 ) , .B2( us03_n760 ) , .A( us03_n778 ) );
  AOI21_X1 us03_U306 (.ZN( us03_n498 ) , .A( us03_n695 ) , .B1( us03_n706 ) , .B2( us03_n784 ) );
  NOR2_X1 us03_U307 (.ZN( us03_n566 ) , .A1( us03_n727 ) , .A2( us03_n760 ) );
  AOI21_X1 us03_U308 (.ZN( us03_n637 ) , .B2( us03_n747 ) , .A( us03_n786 ) , .B1( us03_n810 ) );
  NOR2_X1 us03_U309 (.ZN( us03_n564 ) , .A2( us03_n695 ) , .A1( us03_n761 ) );
  NOR4_X1 us03_U31 (.A4( us03_n774 ) , .A3( us03_n775 ) , .A1( us03_n776 ) , .ZN( us03_n797 ) , .A2( us03_n799 ) );
  NOR2_X1 us03_U310 (.ZN( us03_n578 ) , .A2( us03_n695 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U311 (.ZN( us03_n512 ) , .A( us03_n777 ) , .B2( us03_n790 ) , .B1( us03_n810 ) );
  INV_X1 us03_U312 (.A( us03_n697 ) , .ZN( us03_n851 ) );
  NOR2_X1 us03_U313 (.ZN( us03_n663 ) , .A1( us03_n778 ) , .A2( us03_n811 ) );
  AOI21_X1 us03_U314 (.ZN( us03_n448 ) , .B2( us03_n790 ) , .A( us03_n801 ) , .B1( us03_n813 ) );
  NOR2_X1 us03_U315 (.ZN( us03_n630 ) , .A2( us03_n695 ) , .A1( us03_n722 ) );
  AOI21_X1 us03_U316 (.ZN( us03_n562 ) , .B1( us03_n722 ) , .A( us03_n777 ) , .B2( us03_n789 ) );
  AOI21_X1 us03_U317 (.ZN( us03_n687 ) , .B2( us03_n747 ) , .B1( us03_n761 ) , .A( us03_n804 ) );
  NOR2_X1 us03_U318 (.ZN( us03_n527 ) , .A1( us03_n706 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U319 (.ZN( us03_n576 ) , .A1( us03_n706 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U32 (.ZN( us03_n802 ) , .A1( us03_n852 ) , .A2( us03_n859 ) );
  AOI21_X1 us03_U320 (.ZN( us03_n648 ) , .A( us03_n777 ) , .B1( us03_n790 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U321 (.ZN( us03_n682 ) , .A1( us03_n789 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U322 (.A2( us03_n811 ) , .A1( us03_n813 ) , .ZN( us03_n819 ) );
  AOI21_X1 us03_U323 (.A( us03_n788 ) , .B2( us03_n789 ) , .B1( us03_n790 ) , .ZN( us03_n791 ) );
  AOI21_X1 us03_U324 (.A( us03_n731 ) , .ZN( us03_n732 ) , .B2( us03_n778 ) , .B1( us03_n790 ) );
  NOR2_X1 us03_U325 (.ZN( us03_n565 ) , .A1( us03_n745 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U326 (.ZN( us03_n581 ) , .A1( us03_n790 ) , .A2( us03_n815 ) );
  NOR2_X1 us03_U327 (.ZN( us03_n532 ) , .A1( us03_n722 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U328 (.ZN( us03_n639 ) , .B1( us03_n678 ) , .A( us03_n789 ) , .B2( us03_n815 ) );
  NOR2_X1 us03_U329 (.ZN( us03_n709 ) , .A1( us03_n760 ) , .A2( us03_n761 ) );
  NAND4_X1 us03_U33 (.ZN( sa03_sr_7 ) , .A4( us03_n820 ) , .A3( us03_n821 ) , .A2( us03_n822 ) , .A1( us03_n823 ) );
  NOR2_X1 us03_U330 (.ZN( us03_n680 ) , .A2( us03_n706 ) , .A1( us03_n815 ) );
  INV_X1 us03_U331 (.A( us03_n695 ) , .ZN( us03_n836 ) );
  INV_X1 us03_U332 (.A( us03_n813 ) , .ZN( us03_n853 ) );
  AOI21_X1 us03_U333 (.ZN( us03_n440 ) , .A( us03_n697 ) , .B1( us03_n731 ) , .B2( us03_n748 ) );
  OAI21_X1 us03_U334 (.A( us03_n696 ) , .ZN( us03_n700 ) , .B2( us03_n748 ) , .B1( us03_n802 ) );
  OAI21_X1 us03_U335 (.ZN( us03_n696 ) , .B2( us03_n831 ) , .B1( us03_n836 ) , .A( us03_n858 ) );
  INV_X1 us03_U336 (.A( us03_n778 ) , .ZN( us03_n848 ) );
  AOI22_X1 us03_U337 (.A2( us03_n780 ) , .ZN( us03_n781 ) , .B2( us03_n829 ) , .A1( us03_n832 ) , .B1( us03_n861 ) );
  NAND2_X1 us03_U338 (.ZN( us03_n712 ) , .A1( us03_n726 ) , .A2( us03_n778 ) );
  NAND2_X1 us03_U339 (.ZN( us03_n751 ) , .A1( us03_n761 ) , .A2( us03_n803 ) );
  NOR4_X1 us03_U34 (.A4( us03_n816 ) , .A3( us03_n817 ) , .A2( us03_n818 ) , .A1( us03_n819 ) , .ZN( us03_n820 ) );
  NAND2_X1 us03_U340 (.A2( us03_n760 ) , .A1( us03_n804 ) , .ZN( us03_n808 ) );
  AOI21_X1 us03_U341 (.ZN( us03_n441 ) , .B1( us03_n787 ) , .B2( us03_n789 ) , .A( us03_n812 ) );
  NAND2_X2 us03_U342 (.A1( us03_n449 ) , .A2( us03_n460 ) , .ZN( us03_n788 ) );
  OAI21_X1 us03_U343 (.A( us03_n785 ) , .B2( us03_n786 ) , .B1( us03_n787 ) , .ZN( us03_n793 ) );
  OAI21_X1 us03_U344 (.ZN( us03_n785 ) , .A( us03_n837 ) , .B1( us03_n861 ) , .B2( us03_n871 ) );
  AOI21_X1 us03_U345 (.ZN( us03_n495 ) , .A( us03_n777 ) , .B2( us03_n789 ) , .B1( us03_n802 ) );
  INV_X1 us03_U347 (.A( us03_n783 ) , .ZN( us03_n844 ) );
  NOR2_X1 us03_U348 (.ZN( us03_n468 ) , .A2( us03_n777 ) , .A1( us03_n813 ) );
  OAI21_X1 us03_U349 (.A( us03_n729 ) , .B1( us03_n730 ) , .ZN( us03_n734 ) , .B2( us03_n803 ) );
  AOI222_X1 us03_U35 (.C2( us03_n807 ) , .B2( us03_n808 ) , .A2( us03_n809 ) , .ZN( us03_n821 ) , .C1( us03_n830 ) , .A1( us03_n837 ) , .B1( us03_n851 ) );
  OAI21_X1 us03_U350 (.ZN( us03_n729 ) , .A( us03_n831 ) , .B2( us03_n850 ) , .B1( us03_n871 ) );
  NOR2_X1 us03_U351 (.ZN( us03_n524 ) , .A1( us03_n722 ) , .A2( us03_n748 ) );
  NOR2_X1 us03_U352 (.ZN( us03_n710 ) , .A2( us03_n722 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U353 (.ZN( us03_n482 ) , .A1( us03_n786 ) , .A2( us03_n803 ) );
  NAND2_X1 us03_U354 (.A1( us03_n697 ) , .A2( us03_n727 ) , .ZN( us03_n780 ) );
  NOR2_X1 us03_U355 (.ZN( us03_n516 ) , .A1( us03_n706 ) , .A2( us03_n786 ) );
  NAND2_X1 us03_U356 (.ZN( us03_n669 ) , .A1( us03_n804 ) , .A2( us03_n814 ) );
  NAND2_X1 us03_U357 (.A2( us03_n747 ) , .A1( us03_n784 ) , .ZN( us03_n807 ) );
  INV_X1 us03_U358 (.A( us03_n722 ) , .ZN( us03_n854 ) );
  INV_X1 us03_U359 (.A( us03_n815 ) , .ZN( us03_n842 ) );
  AOI211_X1 us03_U36 (.B( us03_n805 ) , .A( us03_n806 ) , .ZN( us03_n822 ) , .C1( us03_n840 ) , .C2( us03_n848 ) );
  AND2_X1 us03_U360 (.ZN( us03_n730 ) , .A1( us03_n777 ) , .A2( us03_n783 ) );
  NAND2_X1 us03_U361 (.A1( us03_n453 ) , .A2( us03_n469 ) , .ZN( us03_n801 ) );
  NAND2_X1 us03_U362 (.A1( us03_n449 ) , .A2( us03_n452 ) , .ZN( us03_n812 ) );
  NAND2_X1 us03_U363 (.A1( us03_n449 ) , .A2( us03_n469 ) , .ZN( us03_n814 ) );
  NAND2_X1 us03_U364 (.A1( us03_n452 ) , .A2( us03_n459 ) , .ZN( us03_n811 ) );
  NAND2_X1 us03_U365 (.A1( us03_n451 ) , .A2( us03_n459 ) , .ZN( us03_n742 ) );
  NAND2_X1 us03_U367 (.A2( us03_n446 ) , .A1( us03_n458 ) , .ZN( us03_n726 ) );
  NAND2_X1 us03_U368 (.A1( us03_n453 ) , .A2( us03_n460 ) , .ZN( us03_n748 ) );
  NAND2_X1 us03_U369 (.A2( us03_n451 ) , .A1( us03_n453 ) , .ZN( us03_n804 ) );
  NOR2_X1 us03_U37 (.ZN( us03_n746 ) , .A1( us03_n859 ) , .A2( us03_n860 ) );
  NAND2_X1 us03_U370 (.A2( us03_n452 ) , .A1( us03_n470 ) , .ZN( us03_n777 ) );
  NAND2_X1 us03_U371 (.A1( us03_n451 ) , .A2( us03_n470 ) , .ZN( us03_n783 ) );
  NAND2_X1 us03_U374 (.A2( us03_n447 ) , .A1( us03_n450 ) , .ZN( us03_n761 ) );
  NAND2_X1 us03_U375 (.A2( us03_n446 ) , .A1( us03_n450 ) , .ZN( us03_n727 ) );
  NOR2_X1 us03_U376 (.ZN( us03_n445 ) , .A2( us03_n847 ) , .A1( us03_n856 ) );
  NAND2_X1 us03_U377 (.A2( us03_n459 ) , .A1( us03_n460 ) , .ZN( us03_n745 ) );
  NAND2_X1 us03_U378 (.A1( us03_n460 ) , .A2( us03_n470 ) , .ZN( us03_n786 ) );
  NOR2_X1 us03_U38 (.ZN( us03_n623 ) , .A2( us03_n834 ) , .A1( us03_n837 ) );
  NAND2_X2 us03_U380 (.A2( us03_n459 ) , .A1( us03_n469 ) , .ZN( us03_n695 ) );
  NOR2_X1 us03_U381 (.ZN( us03_n451 ) , .A1( us03_n824 ) , .A2( us03_n825 ) );
  NOR2_X1 us03_U382 (.ZN( us03_n449 ) , .A1( us03_n826 ) , .A2( us03_n827 ) );
  NAND2_X1 us03_U383 (.A2( us03_n452 ) , .A1( us03_n453 ) , .ZN( us03_n728 ) );
  NAND2_X2 us03_U384 (.A2( us03_n446 ) , .A1( us03_n462 ) , .ZN( us03_n813 ) );
  NAND2_X2 us03_U386 (.A1( us03_n447 ) , .A2( us03_n462 ) , .ZN( us03_n722 ) );
  NAND2_X2 us03_U387 (.A1( us03_n447 ) , .A2( us03_n458 ) , .ZN( us03_n790 ) );
  NAND2_X2 us03_U389 (.A2( us03_n469 ) , .A1( us03_n470 ) , .ZN( us03_n815 ) );
  NAND4_X1 us03_U39 (.A4( us03_n601 ) , .A3( us03_n602 ) , .A2( us03_n603 ) , .A1( us03_n604 ) , .ZN( us03_n720 ) );
  NAND2_X1 us03_U391 (.A1( us03_n445 ) , .A2( us03_n447 ) , .ZN( us03_n803 ) );
  NOR2_X1 us03_U393 (.A2( sa03_6 ) , .A1( sa03_7 ) , .ZN( us03_n462 ) );
  NOR2_X1 us03_U396 (.A2( sa03_7 ) , .ZN( us03_n458 ) , .A1( us03_n847 ) );
  NOR2_X1 us03_U398 (.A2( sa03_1 ) , .ZN( us03_n469 ) , .A1( us03_n824 ) );
  NOR2_X1 us03_U399 (.A2( sa03_2 ) , .A1( sa03_3 ) , .ZN( us03_n470 ) );
  NOR3_X1 us03_U4 (.A3( us03_n798 ) , .A2( us03_n799 ) , .A1( us03_n800 ) , .ZN( us03_n823 ) );
  NOR3_X1 us03_U40 (.A1( us03_n597 ) , .ZN( us03_n602 ) , .A3( us03_n661 ) , .A2( us03_n768 ) );
  NOR2_X1 us03_U400 (.A2( sa03_6 ) , .ZN( us03_n450 ) , .A1( us03_n856 ) );
  NOR2_X1 us03_U401 (.A2( sa03_2 ) , .ZN( us03_n459 ) , .A1( us03_n827 ) );
  NOR2_X1 us03_U402 (.A2( sa03_0 ) , .ZN( us03_n452 ) , .A1( us03_n825 ) );
  NOR2_X1 us03_U403 (.A2( sa03_0 ) , .A1( sa03_1 ) , .ZN( us03_n460 ) );
  NOR2_X1 us03_U404 (.A2( sa03_3 ) , .ZN( us03_n453 ) , .A1( us03_n826 ) );
  INV_X1 us03_U405 (.A( sa03_6 ) , .ZN( us03_n847 ) );
  INV_X1 us03_U406 (.A( sa03_3 ) , .ZN( us03_n827 ) );
  INV_X1 us03_U407 (.A( sa03_1 ) , .ZN( us03_n825 ) );
  INV_X1 us03_U408 (.A( sa03_0 ) , .ZN( us03_n824 ) );
  INV_X1 us03_U409 (.A( sa03_2 ) , .ZN( us03_n826 ) );
  NOR4_X1 us03_U41 (.A3( us03_n598 ) , .A2( us03_n599 ) , .A1( us03_n600 ) , .ZN( us03_n601 ) , .A4( us03_n653 ) );
  INV_X1 us03_U410 (.A( sa03_7 ) , .ZN( us03_n856 ) );
  AOI222_X1 us03_U412 (.ZN( us03_n603 ) , .B2( us03_n669 ) , .B1( us03_n751 ) , .C2( us03_n829 ) , .A1( us03_n831 ) , .A2( us03_n860 ) , .C1( us03_n861 ) );
  AOI222_X1 us03_U413 (.ZN( us03_n511 ) , .C1( us03_n830 ) , .B2( us03_n835 ) , .A2( us03_n841 ) , .C2( us03_n860 ) , .B1( us03_n861 ) , .A1( us03_n864 ) );
  AOI221_X1 us03_U414 (.A( us03_n481 ) , .ZN( us03_n486 ) , .B1( us03_n829 ) , .C2( us03_n842 ) , .C1( us03_n850 ) , .B2( us03_n860 ) );
  NOR2_X1 us03_U415 (.ZN( us03_n787 ) , .A2( us03_n860 ) , .A1( us03_n866 ) );
  NAND4_X1 us03_U416 (.ZN( sa03_sr_2 ) , .A4( us03_n641 ) , .A3( us03_n642 ) , .A2( us03_n643 ) , .A1( us03_n644 ) );
  OAI221_X1 us03_U417 (.A( us03_n781 ) , .C2( us03_n782 ) , .B2( us03_n783 ) , .B1( us03_n784 ) , .ZN( us03_n794 ) , .C1( us03_n811 ) );
  NAND2_X1 us03_U418 (.A1( us03_n727 ) , .A2( us03_n782 ) , .ZN( us03_n809 ) );
  OAI22_X1 us03_U419 (.ZN( us03_n586 ) , .A2( us03_n745 ) , .B2( us03_n760 ) , .A1( us03_n761 ) , .B1( us03_n782 ) );
  AOI222_X1 us03_U42 (.ZN( us03_n604 ) , .A1( us03_n828 ) , .C2( us03_n835 ) , .B1( us03_n840 ) , .A2( us03_n854 ) , .B2( us03_n859 ) , .C1( us03_n866 ) );
  OAI221_X1 us03_U420 (.A( us03_n694 ) , .ZN( us03_n701 ) , .C2( us03_n782 ) , .C1( us03_n783 ) , .B1( us03_n784 ) , .B2( us03_n804 ) );
  AOI21_X1 us03_U421 (.ZN( us03_n590 ) , .B1( us03_n726 ) , .B2( us03_n782 ) , .A( us03_n788 ) );
  AOI21_X1 us03_U422 (.ZN( us03_n621 ) , .B1( us03_n697 ) , .A( us03_n777 ) , .B2( us03_n782 ) );
  AOI21_X1 us03_U423 (.ZN( us03_n646 ) , .A( us03_n760 ) , .B2( us03_n782 ) , .B1( us03_n790 ) );
  OAI22_X1 us03_U424 (.ZN( us03_n679 ) , .A1( us03_n697 ) , .A2( us03_n728 ) , .B2( us03_n782 ) , .B1( us03_n815 ) );
  OAI21_X1 us03_U425 (.A( us03_n611 ) , .ZN( us03_n614 ) , .B1( us03_n623 ) , .B2( us03_n782 ) );
  NOR2_X1 us03_U426 (.ZN( us03_n608 ) , .A1( us03_n782 ) , .A2( us03_n814 ) );
  OAI222_X1 us03_U427 (.A2( us03_n667 ) , .ZN( us03_n672 ) , .B1( us03_n745 ) , .B2( us03_n782 ) , .C2( us03_n786 ) , .C1( us03_n813 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U428 (.ZN( us03_n649 ) , .A1( us03_n782 ) , .A2( us03_n786 ) );
  NOR2_X1 us03_U429 (.ZN( us03_n598 ) , .A2( us03_n695 ) , .A1( us03_n782 ) );
  NAND4_X1 us03_U43 (.ZN( sa03_sr_3 ) , .A4( us03_n702 ) , .A3( us03_n703 ) , .A2( us03_n704 ) , .A1( us03_n705 ) );
  NOR2_X1 us03_U430 (.ZN( us03_n551 ) , .A2( us03_n742 ) , .A1( us03_n782 ) );
  INV_X1 us03_U431 (.A( us03_n782 ) , .ZN( us03_n859 ) );
  AOI221_X1 us03_U432 (.A( us03_n574 ) , .ZN( us03_n585 ) , .B2( us03_n829 ) , .C2( us03_n841 ) , .B1( us03_n852 ) , .C1( us03_n859 ) );
  AOI21_X1 us03_U433 (.ZN( us03_n574 ) , .B2( us03_n722 ) , .B1( us03_n746 ) , .A( us03_n783 ) );
  AOI211_X1 us03_U434 (.A( us03_n635 ) , .ZN( us03_n643 ) , .B( us03_n741 ) , .C2( us03_n837 ) , .C1( us03_n852 ) );
  NAND4_X1 us03_U435 (.A4( us03_n631 ) , .A3( us03_n632 ) , .A2( us03_n633 ) , .A1( us03_n634 ) , .ZN( us03_n741 ) );
  NAND3_X1 us03_U437 (.ZN( sa03_sr_6 ) , .A3( us03_n795 ) , .A2( us03_n796 ) , .A1( us03_n797 ) );
  NAND3_X1 us03_U438 (.ZN( sa03_sr_5 ) , .A3( us03_n756 ) , .A2( us03_n757 ) , .A1( us03_n758 ) );
  NAND3_X1 us03_U439 (.ZN( sa03_sr_4 ) , .A3( us03_n736 ) , .A2( us03_n737 ) , .A1( us03_n738 ) );
  NOR4_X1 us03_U44 (.A4( us03_n698 ) , .A3( us03_n699 ) , .A2( us03_n700 ) , .A1( us03_n701 ) , .ZN( us03_n702 ) );
  NAND3_X1 us03_U440 (.A3( us03_n673 ) , .A2( us03_n674 ) , .A1( us03_n675 ) , .ZN( us03_n805 ) );
  NAND3_X1 us03_U441 (.ZN( us03_n636 ) , .A3( us03_n706 ) , .A2( us03_n722 ) , .A1( us03_n790 ) );
  NAND3_X1 us03_U442 (.A3( us03_n616 ) , .A2( us03_n617 ) , .A1( us03_n618 ) , .ZN( us03_n723 ) );
  NAND3_X1 us03_U443 (.A3( us03_n583 ) , .A2( us03_n584 ) , .A1( us03_n585 ) , .ZN( us03_n619 ) );
  NAND3_X1 us03_U444 (.ZN( us03_n563 ) , .A3( us03_n678 ) , .A2( us03_n748 ) , .A1( us03_n783 ) );
  NAND3_X1 us03_U445 (.A3( us03_n521 ) , .A2( us03_n522 ) , .A1( us03_n523 ) , .ZN( us03_n740 ) );
  NAND3_X1 us03_U446 (.A3( us03_n510 ) , .A1( us03_n511 ) , .ZN( us03_n606 ) , .A2( us03_n869 ) );
  NAND3_X1 us03_U447 (.A3( us03_n465 ) , .A2( us03_n466 ) , .A1( us03_n467 ) , .ZN( us03_n775 ) );
  AOI211_X1 us03_U45 (.B( us03_n692 ) , .A( us03_n693 ) , .ZN( us03_n703 ) , .C2( us03_n829 ) , .C1( us03_n849 ) );
  NOR2_X1 us03_U46 (.ZN( us03_n705 ) , .A2( us03_n774 ) , .A1( us03_n798 ) );
  AOI222_X1 us03_U47 (.ZN( us03_n467 ) , .B1( us03_n830 ) , .A1( us03_n837 ) , .C1( us03_n840 ) , .C2( us03_n849 ) , .A2( us03_n853 ) , .B2( us03_n863 ) );
  NOR4_X1 us03_U48 (.A1( us03_n464 ) , .ZN( us03_n465 ) , .A4( us03_n540 ) , .A2( us03_n552 ) , .A3( us03_n612 ) );
  AOI221_X1 us03_U49 (.ZN( us03_n466 ) , .C2( us03_n712 ) , .B2( us03_n829 ) , .C1( us03_n843 ) , .B1( us03_n858 ) , .A( us03_n862 ) );
  NOR3_X1 us03_U5 (.ZN( us03_n502 ) , .A2( us03_n677 ) , .A3( us03_n775 ) , .A1( us03_n874 ) );
  NOR4_X1 us03_U50 (.A4( us03_n575 ) , .A3( us03_n576 ) , .A2( us03_n577 ) , .ZN( us03_n584 ) , .A1( us03_n681 ) );
  NOR4_X1 us03_U51 (.A1( us03_n582 ) , .ZN( us03_n583 ) , .A3( us03_n650 ) , .A2( us03_n660 ) , .A4( us03_n765 ) );
  NAND4_X1 us03_U52 (.A4( us03_n483 ) , .A3( us03_n484 ) , .A2( us03_n485 ) , .A1( us03_n486 ) , .ZN( us03_n776 ) );
  NOR4_X1 us03_U53 (.A4( us03_n482 ) , .ZN( us03_n485 ) , .A1( us03_n564 ) , .A2( us03_n579 ) , .A3( us03_n600 ) );
  NOR4_X1 us03_U54 (.ZN( us03_n484 ) , .A1( us03_n505 ) , .A2( us03_n517 ) , .A4( us03_n544 ) , .A3( us03_n609 ) );
  NOR4_X1 us03_U55 (.ZN( us03_n483 ) , .A2( us03_n531 ) , .A1( us03_n556 ) , .A3( us03_n629 ) , .A4( us03_n716 ) );
  AOI211_X1 us03_U56 (.B( us03_n621 ) , .A( us03_n622 ) , .ZN( us03_n633 ) , .C2( us03_n834 ) , .C1( us03_n861 ) );
  NOR4_X1 us03_U57 (.A4( us03_n627 ) , .A3( us03_n628 ) , .A2( us03_n629 ) , .A1( us03_n630 ) , .ZN( us03_n631 ) );
  NOR4_X1 us03_U58 (.A4( us03_n624 ) , .A3( us03_n625 ) , .A2( us03_n626 ) , .ZN( us03_n632 ) , .A1( us03_n662 ) );
  NAND4_X1 us03_U59 (.A4( us03_n655 ) , .A3( us03_n656 ) , .A2( us03_n657 ) , .A1( us03_n658 ) , .ZN( us03_n798 ) );
  INV_X1 us03_U6 (.A( us03_n704 ) , .ZN( us03_n874 ) );
  NOR3_X1 us03_U60 (.A3( us03_n646 ) , .A2( us03_n647 ) , .A1( us03_n648 ) , .ZN( us03_n657 ) );
  NOR3_X1 us03_U61 (.A3( us03_n649 ) , .A2( us03_n650 ) , .A1( us03_n651 ) , .ZN( us03_n656 ) );
  NOR3_X1 us03_U62 (.A3( us03_n652 ) , .A2( us03_n653 ) , .A1( us03_n654 ) , .ZN( us03_n655 ) );
  NAND4_X1 us03_U63 (.A4( us03_n558 ) , .A3( us03_n559 ) , .A2( us03_n560 ) , .A1( us03_n561 ) , .ZN( us03_n605 ) );
  NOR4_X1 us03_U64 (.A4( us03_n554 ) , .A3( us03_n555 ) , .A2( us03_n556 ) , .A1( us03_n557 ) , .ZN( us03_n558 ) );
  NOR4_X1 us03_U65 (.ZN( us03_n559 ) , .A1( us03_n651 ) , .A3( us03_n659 ) , .A4( us03_n683 ) , .A2( us03_n766 ) );
  NOR4_X1 us03_U66 (.A4( us03_n550 ) , .A3( us03_n551 ) , .A2( us03_n552 ) , .A1( us03_n553 ) , .ZN( us03_n560 ) );
  NAND4_X1 us03_U67 (.A4( us03_n770 ) , .A3( us03_n771 ) , .A2( us03_n772 ) , .A1( us03_n773 ) , .ZN( us03_n799 ) );
  NOR3_X1 us03_U68 (.A3( us03_n763 ) , .A2( us03_n764 ) , .A1( us03_n765 ) , .ZN( us03_n771 ) );
  NOR4_X1 us03_U69 (.A4( us03_n766 ) , .A3( us03_n767 ) , .A2( us03_n768 ) , .A1( us03_n769 ) , .ZN( us03_n770 ) );
  NOR3_X1 us03_U7 (.A3( us03_n619 ) , .A2( us03_n620 ) , .ZN( us03_n634 ) , .A1( us03_n723 ) );
  AOI222_X1 us03_U70 (.ZN( us03_n773 ) , .A1( us03_n828 ) , .C1( us03_n832 ) , .B2( us03_n839 ) , .A2( us03_n848 ) , .B1( us03_n859 ) , .C2( us03_n871 ) );
  NOR4_X1 us03_U71 (.A4( us03_n507 ) , .A2( us03_n508 ) , .A1( us03_n509 ) , .ZN( us03_n510 ) , .A3( us03_n668 ) );
  INV_X1 us03_U72 (.A( us03_n503 ) , .ZN( us03_n869 ) );
  NOR4_X1 us03_U73 (.A4( us03_n663 ) , .A3( us03_n664 ) , .A2( us03_n665 ) , .A1( us03_n666 ) , .ZN( us03_n674 ) );
  NOR4_X1 us03_U74 (.A4( us03_n659 ) , .A3( us03_n660 ) , .A2( us03_n661 ) , .A1( us03_n662 ) , .ZN( us03_n675 ) );
  NOR4_X1 us03_U75 (.A3( us03_n671 ) , .A1( us03_n672 ) , .ZN( us03_n673 ) , .A4( us03_n713 ) , .A2( us03_n857 ) );
  NOR2_X1 us03_U76 (.ZN( us03_n759 ) , .A1( us03_n831 ) , .A2( us03_n832 ) );
  NOR4_X1 us03_U77 (.A4( us03_n732 ) , .A3( us03_n733 ) , .A2( us03_n734 ) , .A1( us03_n735 ) , .ZN( us03_n736 ) );
  AOI211_X1 us03_U78 (.B( us03_n723 ) , .A( us03_n724 ) , .ZN( us03_n737 ) , .C1( us03_n841 ) , .C2( us03_n853 ) );
  NOR3_X1 us03_U79 (.A3( us03_n720 ) , .A1( us03_n721 ) , .ZN( us03_n738 ) , .A2( us03_n739 ) );
  NOR2_X1 us03_U8 (.ZN( us03_n573 ) , .A1( us03_n620 ) , .A2( us03_n743 ) );
  NOR4_X1 us03_U80 (.A3( us03_n753 ) , .A2( us03_n754 ) , .A1( us03_n755 ) , .ZN( us03_n756 ) , .A4( us03_n867 ) );
  AOI211_X1 us03_U81 (.B( us03_n743 ) , .A( us03_n744 ) , .ZN( us03_n757 ) , .C1( us03_n830 ) , .C2( us03_n851 ) );
  NOR3_X1 us03_U82 (.A3( us03_n739 ) , .A2( us03_n740 ) , .A1( us03_n741 ) , .ZN( us03_n758 ) );
  NAND4_X1 us03_U83 (.A4( us03_n454 ) , .A3( us03_n455 ) , .A2( us03_n456 ) , .A1( us03_n457 ) , .ZN( us03_n677 ) );
  NOR3_X1 us03_U84 (.ZN( us03_n455 ) , .A3( us03_n528 ) , .A1( us03_n553 ) , .A2( us03_n568 ) );
  AOI221_X1 us03_U85 (.A( us03_n448 ) , .ZN( us03_n457 ) , .C2( us03_n751 ) , .B1( us03_n830 ) , .C1( us03_n840 ) , .B2( us03_n859 ) );
  NOR4_X1 us03_U86 (.ZN( us03_n456 ) , .A2( us03_n507 ) , .A1( us03_n597 ) , .A4( us03_n626 ) , .A3( us03_n709 ) );
  NAND4_X1 us03_U87 (.A4( us03_n533 ) , .A3( us03_n534 ) , .A2( us03_n535 ) , .A1( us03_n536 ) , .ZN( us03_n620 ) );
  NOR4_X1 us03_U88 (.A4( us03_n524 ) , .A2( us03_n525 ) , .A1( us03_n526 ) , .ZN( us03_n536 ) , .A3( us03_n699 ) );
  NOR4_X1 us03_U89 (.A1( us03_n529 ) , .ZN( us03_n534 ) , .A2( us03_n652 ) , .A4( us03_n666 ) , .A3( us03_n763 ) );
  NOR2_X1 us03_U9 (.A1( us03_n676 ) , .ZN( us03_n691 ) , .A2( us03_n805 ) );
  NOR4_X1 us03_U90 (.A4( us03_n527 ) , .A3( us03_n528 ) , .ZN( us03_n535 ) , .A2( us03_n682 ) , .A1( us03_n792 ) );
  NAND4_X1 us03_U91 (.A4( us03_n477 ) , .A3( us03_n478 ) , .A2( us03_n479 ) , .A1( us03_n480 ) , .ZN( us03_n692 ) );
  NOR3_X1 us03_U92 (.ZN( us03_n478 ) , .A2( us03_n506 ) , .A3( us03_n599 ) , .A1( us03_n608 ) );
  AOI211_X1 us03_U93 (.B( us03_n475 ) , .A( us03_n476 ) , .ZN( us03_n480 ) , .C2( us03_n831 ) , .C1( us03_n859 ) );
  NOR4_X1 us03_U94 (.ZN( us03_n479 ) , .A3( us03_n530 ) , .A4( us03_n543 ) , .A2( us03_n565 ) , .A1( us03_n715 ) );
  NAND4_X1 us03_U95 (.A4( us03_n546 ) , .A3( us03_n547 ) , .A2( us03_n548 ) , .A1( us03_n549 ) , .ZN( us03_n743 ) );
  NOR3_X1 us03_U96 (.ZN( us03_n547 ) , .A2( us03_n649 ) , .A1( us03_n665 ) , .A3( us03_n769 ) );
  AOI211_X1 us03_U97 (.B( us03_n537 ) , .A( us03_n538 ) , .ZN( us03_n549 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NOR4_X1 us03_U98 (.A4( us03_n542 ) , .A3( us03_n543 ) , .A2( us03_n544 ) , .A1( us03_n545 ) , .ZN( us03_n546 ) );
  NOR4_X1 us03_U99 (.ZN( us03_n618 ) , .A1( us03_n654 ) , .A3( us03_n664 ) , .A4( us03_n680 ) , .A2( us03_n764 ) );
  NOR2_X1 us33_U10 (.ZN( us33_n495 ) , .A1( us33_n678 ) , .A2( us33_n694 ) );
  NAND4_X1 us33_U100 (.A4( us33_n479 ) , .A3( us33_n480 ) , .A2( us33_n481 ) , .A1( us33_n482 ) , .ZN( us33_n694 ) );
  NOR3_X1 us33_U101 (.ZN( us33_n480 ) , .A2( us33_n508 ) , .A3( us33_n601 ) , .A1( us33_n610 ) );
  AOI211_X1 us33_U102 (.B( us33_n477 ) , .A( us33_n478 ) , .ZN( us33_n482 ) , .C2( us33_n833 ) , .C1( us33_n861 ) );
  NOR4_X1 us33_U103 (.ZN( us33_n481 ) , .A3( us33_n532 ) , .A4( us33_n545 ) , .A2( us33_n567 ) , .A1( us33_n717 ) );
  NAND4_X1 us33_U104 (.A4( us33_n548 ) , .A3( us33_n549 ) , .A2( us33_n550 ) , .A1( us33_n551 ) , .ZN( us33_n745 ) );
  NOR3_X1 us33_U105 (.ZN( us33_n549 ) , .A2( us33_n651 ) , .A1( us33_n667 ) , .A3( us33_n771 ) );
  AOI211_X1 us33_U106 (.B( us33_n539 ) , .A( us33_n540 ) , .ZN( us33_n551 ) , .C2( us33_n839 ) , .C1( us33_n851 ) );
  NOR4_X1 us33_U107 (.A4( us33_n544 ) , .A3( us33_n545 ) , .A2( us33_n546 ) , .A1( us33_n547 ) , .ZN( us33_n548 ) );
  NOR4_X1 us33_U108 (.ZN( us33_n620 ) , .A1( us33_n656 ) , .A3( us33_n666 ) , .A4( us33_n682 ) , .A2( us33_n766 ) );
  NOR4_X1 us33_U109 (.A4( us33_n609 ) , .A3( us33_n610 ) , .A2( us33_n611 ) , .A1( us33_n612 ) , .ZN( us33_n619 ) );
  NOR2_X1 us33_U11 (.A1( us33_n678 ) , .ZN( us33_n693 ) , .A2( us33_n807 ) );
  NOR4_X1 us33_U110 (.A4( us33_n614 ) , .A3( us33_n615 ) , .A2( us33_n616 ) , .A1( us33_n617 ) , .ZN( us33_n618 ) );
  NOR2_X1 us33_U111 (.ZN( us33_n686 ) , .A1( us33_n831 ) , .A2( us33_n832 ) );
  NAND4_X1 us33_U112 (.A4( us33_n485 ) , .A3( us33_n486 ) , .A2( us33_n487 ) , .A1( us33_n488 ) , .ZN( us33_n778 ) );
  NOR4_X1 us33_U113 (.A4( us33_n484 ) , .ZN( us33_n487 ) , .A1( us33_n566 ) , .A2( us33_n581 ) , .A3( us33_n602 ) );
  NOR4_X1 us33_U114 (.ZN( us33_n486 ) , .A1( us33_n507 ) , .A2( us33_n519 ) , .A4( us33_n546 ) , .A3( us33_n611 ) );
  NOR4_X1 us33_U115 (.ZN( us33_n485 ) , .A2( us33_n533 ) , .A1( us33_n558 ) , .A3( us33_n631 ) , .A4( us33_n718 ) );
  NAND4_X1 us33_U116 (.A4( us33_n691 ) , .A3( us33_n692 ) , .A1( us33_n693 ) , .ZN( us33_n776 ) , .A2( us33_n872 ) );
  AOI221_X1 us33_U117 (.A( us33_n681 ) , .ZN( us33_n692 ) , .B2( us33_n840 ) , .C1( us33_n842 ) , .C2( us33_n862 ) , .B1( us33_n865 ) );
  INV_X1 us33_U118 (.A( us33_n679 ) , .ZN( us33_n872 ) );
  NOR4_X1 us33_U119 (.A4( us33_n687 ) , .A3( us33_n688 ) , .A2( us33_n689 ) , .A1( us33_n690 ) , .ZN( us33_n691 ) );
  NOR3_X1 us33_U12 (.ZN( us33_n504 ) , .A2( us33_n679 ) , .A3( us33_n777 ) , .A1( us33_n876 ) );
  NAND4_X1 us33_U120 (.A4( us33_n719 ) , .A3( us33_n720 ) , .A2( us33_n721 ) , .ZN( us33_n741 ) , .A1( us33_n857 ) );
  INV_X1 us33_U121 (.A( us33_n709 ) , .ZN( us33_n857 ) );
  AOI221_X1 us33_U122 (.A( us33_n710 ) , .ZN( us33_n721 ) , .C2( us33_n844 ) , .B2( us33_n845 ) , .C1( us33_n861 ) , .B1( us33_n862 ) );
  NOR4_X1 us33_U123 (.A4( us33_n715 ) , .A3( us33_n716 ) , .A2( us33_n717 ) , .A1( us33_n718 ) , .ZN( us33_n719 ) );
  NAND4_X1 us33_U124 (.A4( us33_n473 ) , .A3( us33_n474 ) , .A2( us33_n475 ) , .A1( us33_n476 ) , .ZN( us33_n678 ) );
  NOR4_X1 us33_U125 (.ZN( us33_n475 ) , .A1( us33_n531 ) , .A3( us33_n568 ) , .A4( us33_n600 ) , .A2( us33_n642 ) );
  NOR4_X1 us33_U126 (.A4( us33_n470 ) , .ZN( us33_n476 ) , .A3( us33_n556 ) , .A1( us33_n735 ) , .A2( us33_n755 ) );
  NOR4_X1 us33_U127 (.ZN( us33_n474 ) , .A1( us33_n506 ) , .A3( us33_n544 ) , .A2( us33_n583 ) , .A4( us33_n716 ) );
  NOR2_X1 us33_U128 (.ZN( us33_n733 ) , .A2( us33_n832 ) , .A1( us33_n845 ) );
  NOR2_X1 us33_U129 (.ZN( us33_n789 ) , .A2( us33_n862 ) , .A1( us33_n868 ) );
  INV_X1 us33_U13 (.A( us33_n706 ) , .ZN( us33_n876 ) );
  NAND4_X1 us33_U130 (.A4( us33_n573 ) , .A3( us33_n574 ) , .A1( us33_n575 ) , .ZN( us33_n723 ) , .A2( us33_n874 ) );
  AOI221_X1 us33_U131 (.A( us33_n564 ) , .C2( us33_n565 ) , .ZN( us33_n574 ) , .B2( us33_n845 ) , .B1( us33_n852 ) , .C1( us33_n853 ) );
  NOR4_X1 us33_U132 (.A4( us33_n569 ) , .A3( us33_n570 ) , .A2( us33_n571 ) , .A1( us33_n572 ) , .ZN( us33_n573 ) );
  INV_X1 us33_U133 (.A( us33_n607 ) , .ZN( us33_n874 ) );
  NAND4_X1 us33_U134 (.A4( us33_n633 ) , .A3( us33_n634 ) , .A2( us33_n635 ) , .A1( us33_n636 ) , .ZN( us33_n743 ) );
  AOI211_X1 us33_U135 (.B( us33_n623 ) , .A( us33_n624 ) , .ZN( us33_n635 ) , .C2( us33_n836 ) , .C1( us33_n863 ) );
  NOR4_X1 us33_U136 (.A4( us33_n629 ) , .A3( us33_n630 ) , .A2( us33_n631 ) , .A1( us33_n632 ) , .ZN( us33_n633 ) );
  NOR4_X1 us33_U137 (.A4( us33_n626 ) , .A3( us33_n627 ) , .A2( us33_n628 ) , .ZN( us33_n634 ) , .A1( us33_n664 ) );
  NAND4_X1 us33_U138 (.A4( us33_n493 ) , .A3( us33_n494 ) , .A1( us33_n495 ) , .ZN( us33_n802 ) , .A2( us33_n867 ) );
  AOI221_X1 us33_U139 (.A( us33_n489 ) , .ZN( us33_n494 ) , .B2( us33_n836 ) , .C2( us33_n841 ) , .C1( us33_n851 ) , .B1( us33_n860 ) );
  INV_X1 us33_U14 (.A( us33_n680 ) , .ZN( us33_n840 ) );
  INV_X1 us33_U140 (.A( us33_n778 ) , .ZN( us33_n867 ) );
  NOR4_X1 us33_U141 (.A2( us33_n491 ) , .A1( us33_n492 ) , .ZN( us33_n493 ) , .A3( us33_n580 ) , .A4( us33_n612 ) );
  NOR4_X1 us33_U142 (.A4( us33_n734 ) , .A3( us33_n735 ) , .A2( us33_n736 ) , .A1( us33_n737 ) , .ZN( us33_n738 ) );
  AOI211_X1 us33_U143 (.B( us33_n725 ) , .A( us33_n726 ) , .ZN( us33_n739 ) , .C1( us33_n843 ) , .C2( us33_n855 ) );
  NOR3_X1 us33_U144 (.A3( us33_n722 ) , .A1( us33_n723 ) , .ZN( us33_n740 ) , .A2( us33_n741 ) );
  INV_X1 us33_U145 (.A( us33_n762 ) , .ZN( us33_n830 ) );
  OR4_X1 us33_U146 (.A4( us33_n566 ) , .A3( us33_n567 ) , .A2( us33_n568 ) , .ZN( us33_n572 ) , .A1( us33_n665 ) );
  OR4_X1 us33_U147 (.A4( us33_n682 ) , .A3( us33_n683 ) , .A2( us33_n684 ) , .A1( us33_n685 ) , .ZN( us33_n690 ) );
  OR4_X1 us33_U148 (.ZN( us33_n466 ) , .A4( us33_n518 ) , .A3( us33_n529 ) , .A2( us33_n578 ) , .A1( us33_n712 ) );
  OR4_X1 us33_U149 (.A4( us33_n518 ) , .A2( us33_n519 ) , .A1( us33_n520 ) , .ZN( us33_n522 ) , .A3( us33_n821 ) );
  NOR4_X1 us33_U15 (.A4( us33_n445 ) , .A3( us33_n446 ) , .A2( us33_n516 ) , .A1( us33_n541 ) , .ZN( us33_n706 ) );
  OR4_X1 us33_U150 (.ZN( us33_n492 ) , .A4( us33_n534 ) , .A2( us33_n547 ) , .A1( us33_n559 ) , .A3( us33_n632 ) );
  OR4_X1 us33_U151 (.A4( us33_n580 ) , .A3( us33_n581 ) , .A2( us33_n582 ) , .A1( us33_n583 ) , .ZN( us33_n584 ) );
  INV_X1 us33_U152 (.A( us33_n697 ) , .ZN( us33_n838 ) );
  NAND2_X1 us33_U153 (.ZN( us33_n613 ) , .A2( us33_n837 ) , .A1( us33_n873 ) );
  OR3_X1 us33_U154 (.A3( us33_n506 ) , .A2( us33_n507 ) , .A1( us33_n508 ) , .ZN( us33_n511 ) );
  INV_X1 us33_U155 (.A( us33_n754 ) , .ZN( us33_n869 ) );
  OAI21_X1 us33_U156 (.B1( us33_n753 ) , .ZN( us33_n754 ) , .A( us33_n845 ) , .B2( us33_n868 ) );
  INV_X1 us33_U157 (.A( us33_n463 ) , .ZN( us33_n864 ) );
  OAI21_X1 us33_U158 (.ZN( us33_n463 ) , .B1( us33_n809 ) , .A( us33_n834 ) , .B2( us33_n851 ) );
  INV_X1 us33_U159 (.A( us33_n672 ) , .ZN( us33_n859 ) );
  OR3_X1 us33_U16 (.ZN( us33_n446 ) , .A1( us33_n528 ) , .A3( us33_n577 ) , .A2( us33_n875 ) );
  AOI21_X1 us33_U160 (.A( us33_n670 ) , .B1( us33_n671 ) , .ZN( us33_n672 ) , .B2( us33_n856 ) );
  OAI222_X1 us33_U161 (.B2( us33_n747 ) , .B1( us33_n748 ) , .A2( us33_n749 ) , .ZN( us33_n757 ) , .C2( us33_n805 ) , .C1( us33_n814 ) , .A1( us33_n817 ) );
  OAI222_X1 us33_U162 (.ZN( us33_n505 ) , .C2( us33_n625 ) , .B2( us33_n647 ) , .B1( us33_n747 ) , .A2( us33_n748 ) , .C1( us33_n805 ) , .A1( us33_n806 ) );
  OAI222_X1 us33_U163 (.B2( us33_n708 ) , .ZN( us33_n709 ) , .C2( us33_n724 ) , .B1( us33_n747 ) , .A1( us33_n806 ) , .C1( us33_n814 ) , .A2( us33_n815 ) );
  NAND2_X1 us33_U164 (.A1( us33_n447 ) , .A2( us33_n465 ) , .ZN( us33_n749 ) );
  AOI22_X1 us33_U165 (.ZN( us33_n696 ) , .A1( us33_n830 ) , .B2( us33_n843 ) , .A2( us33_n865 ) , .B1( us33_n868 ) );
  AOI22_X1 us33_U166 (.A2( us33_n782 ) , .ZN( us33_n783 ) , .B2( us33_n831 ) , .A1( us33_n834 ) , .B1( us33_n863 ) );
  INV_X1 us33_U167 (.A( us33_n730 ) , .ZN( us33_n839 ) );
  AOI221_X1 us33_U168 (.A( us33_n764 ) , .ZN( us33_n774 ) , .C2( us33_n810 ) , .B2( us33_n835 ) , .C1( us33_n855 ) , .B1( us33_n866 ) );
  AOI21_X1 us33_U169 (.B2( us33_n763 ) , .ZN( us33_n764 ) , .A( us33_n788 ) , .B1( us33_n792 ) );
  OR4_X1 us33_U17 (.A4( us33_n442 ) , .A2( us33_n443 ) , .A1( us33_n444 ) , .ZN( us33_n445 ) , .A3( us33_n553 ) );
  INV_X1 us33_U170 (.A( us33_n761 ) , .ZN( us33_n835 ) );
  AOI221_X1 us33_U171 (.A( us33_n483 ) , .ZN( us33_n488 ) , .B1( us33_n831 ) , .C2( us33_n844 ) , .C1( us33_n852 ) , .B2( us33_n862 ) );
  OAI22_X1 us33_U172 (.ZN( us33_n483 ) , .A1( us33_n708 ) , .B2( us33_n785 ) , .A2( us33_n806 ) , .B1( us33_n812 ) );
  INV_X1 us33_U173 (.A( us33_n790 ) , .ZN( us33_n832 ) );
  NAND2_X1 us33_U174 (.A1( us33_n451 ) , .A2( us33_n453 ) , .ZN( us33_n762 ) );
  OAI221_X1 us33_U175 (.A( us33_n727 ) , .C2( us33_n728 ) , .B2( us33_n729 ) , .B1( us33_n730 ) , .ZN( us33_n737 ) , .C1( us33_n817 ) );
  AOI22_X1 us33_U176 (.ZN( us33_n727 ) , .B1( us33_n832 ) , .A2( us33_n838 ) , .A1( us33_n863 ) , .B2( us33_n866 ) );
  INV_X1 us33_U177 (.A( us33_n786 ) , .ZN( us33_n862 ) );
  OAI22_X1 us33_U178 (.ZN( us33_n710 ) , .A2( us33_n728 ) , .B2( us33_n729 ) , .A1( us33_n744 ) , .B1( us33_n813 ) );
  INV_X1 us33_U179 (.A( us33_n816 ) , .ZN( us33_n831 ) );
  INV_X1 us33_U18 (.A( us33_n613 ) , .ZN( us33_n875 ) );
  OAI22_X1 us33_U180 (.ZN( us33_n489 ) , .A1( us33_n724 ) , .B2( us33_n728 ) , .B1( us33_n730 ) , .A2( us33_n779 ) );
  OAI22_X1 us33_U181 (.ZN( us33_n624 ) , .B1( us33_n669 ) , .B2( us33_n747 ) , .A1( us33_n815 ) , .A2( us33_n816 ) );
  INV_X1 us33_U182 (.A( us33_n744 ) , .ZN( us33_n837 ) );
  INV_X1 us33_U183 (.A( us33_n788 ) , .ZN( us33_n845 ) );
  OAI22_X1 us33_U184 (.B2( us33_n779 ) , .B1( us33_n780 ) , .ZN( us33_n781 ) , .A2( us33_n814 ) , .A1( us33_n815 ) );
  OAI22_X1 us33_U185 (.A1( us33_n724 ) , .ZN( us33_n726 ) , .B2( us33_n750 ) , .B1( us33_n812 ) , .A2( us33_n816 ) );
  INV_X1 us33_U186 (.A( us33_n805 ) , .ZN( us33_n860 ) );
  INV_X1 us33_U187 (.A( us33_n814 ) , .ZN( us33_n833 ) );
  INV_X1 us33_U188 (.A( us33_n669 ) , .ZN( us33_n865 ) );
  OAI22_X1 us33_U189 (.B2( us33_n744 ) , .ZN( us33_n746 ) , .A2( us33_n762 ) , .B1( us33_n780 ) , .A1( us33_n792 ) );
  INV_X1 us33_U19 (.A( us33_n749 ) , .ZN( us33_n863 ) );
  OAI22_X1 us33_U190 (.ZN( us33_n496 ) , .A2( us33_n744 ) , .A1( us33_n780 ) , .B1( us33_n791 ) , .B2( us33_n806 ) );
  OAI22_X1 us33_U191 (.B2( us33_n803 ) , .B1( us33_n804 ) , .A2( us33_n805 ) , .A1( us33_n806 ) , .ZN( us33_n808 ) );
  AOI211_X1 us33_U192 (.A( us33_n637 ) , .ZN( us33_n645 ) , .B( us33_n743 ) , .C2( us33_n839 ) , .C1( us33_n854 ) );
  OAI22_X1 us33_U193 (.ZN( us33_n637 ) , .A1( us33_n699 ) , .B2( us33_n728 ) , .A2( us33_n762 ) , .B1( us33_n816 ) );
  OAI22_X1 us33_U194 (.B1( us33_n490 ) , .ZN( us33_n491 ) , .A1( us33_n686 ) , .A2( us33_n763 ) , .B2( us33_n817 ) );
  NOR3_X1 us33_U195 (.ZN( us33_n490 ) , .A1( us33_n782 ) , .A2( us33_n850 ) , .A3( us33_n863 ) );
  INV_X1 us33_U196 (.A( us33_n750 ) , .ZN( us33_n842 ) );
  OAI22_X1 us33_U197 (.ZN( us33_n695 ) , .A2( us33_n730 ) , .A1( us33_n780 ) , .B1( us33_n791 ) , .B2( us33_n817 ) );
  NOR2_X1 us33_U198 (.ZN( us33_n715 ) , .A1( us33_n805 ) , .A2( us33_n817 ) );
  NOR2_X1 us33_U199 (.ZN( us33_n666 ) , .A1( us33_n728 ) , .A2( us33_n803 ) );
  AOI222_X1 us33_U20 (.ZN( us33_n605 ) , .B2( us33_n671 ) , .B1( us33_n753 ) , .C2( us33_n831 ) , .A1( us33_n833 ) , .A2( us33_n862 ) , .C1( us33_n863 ) );
  NOR2_X1 us33_U200 (.ZN( us33_n594 ) , .A2( us33_n697 ) , .A1( us33_n728 ) );
  NOR2_X1 us33_U201 (.ZN( us33_n570 ) , .A1( us33_n728 ) , .A2( us33_n806 ) );
  NOR2_X1 us33_U202 (.A2( us33_n744 ) , .ZN( us33_n755 ) , .A1( us33_n805 ) );
  NOR2_X1 us33_U203 (.ZN( us33_n735 ) , .A2( us33_n803 ) , .A1( us33_n805 ) );
  NOR2_X1 us33_U204 (.ZN( us33_n546 ) , .A2( us33_n780 ) , .A1( us33_n814 ) );
  NOR2_X1 us33_U205 (.ZN( us33_n577 ) , .A2( us33_n699 ) , .A1( us33_n814 ) );
  NOR2_X1 us33_U206 (.ZN( us33_n654 ) , .A1( us33_n728 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U207 (.ZN( us33_n718 ) , .A2( us33_n724 ) , .A1( us33_n744 ) );
  NOR2_X1 us33_U208 (.ZN( us33_n532 ) , .A2( us33_n749 ) , .A1( us33_n750 ) );
  NOR2_X1 us33_U209 (.ZN( us33_n615 ) , .A1( us33_n785 ) , .A2( us33_n815 ) );
  AOI222_X1 us33_U21 (.ZN( us33_n563 ) , .B1( us33_n830 ) , .C1( us33_n841 ) , .A2( us33_n843 ) , .A1( us33_n854 ) , .B2( us33_n863 ) , .C2( us33_n873 ) );
  NOR2_X1 us33_U210 (.ZN( us33_n629 ) , .A2( us33_n728 ) , .A1( us33_n785 ) );
  NOR2_X1 us33_U211 (.ZN( us33_n611 ) , .A2( us33_n780 ) , .A1( us33_n806 ) );
  NOR2_X1 us33_U212 (.ZN( us33_n628 ) , .A2( us33_n669 ) , .A1( us33_n785 ) );
  INV_X1 us33_U213 (.A( us33_n747 ) , .ZN( us33_n834 ) );
  INV_X1 us33_U214 (.A( us33_n728 ) , .ZN( us33_n852 ) );
  NOR2_X1 us33_U215 (.ZN( us33_n652 ) , .A1( us33_n669 ) , .A2( us33_n814 ) );
  NOR2_X1 us33_U216 (.A1( us33_n669 ) , .ZN( us33_n673 ) , .A2( us33_n744 ) );
  NOR2_X1 us33_U217 (.ZN( us33_n602 ) , .A1( us33_n669 ) , .A2( us33_n803 ) );
  NOR2_X1 us33_U218 (.A1( us33_n669 ) , .ZN( us33_n688 ) , .A2( us33_n816 ) );
  NOR2_X1 us33_U219 (.A2( us33_n744 ) , .ZN( us33_n769 ) , .A1( us33_n812 ) );
  AOI222_X1 us33_U22 (.ZN( us33_n660 ) , .A2( us33_n839 ) , .B1( us33_n841 ) , .C2( us33_n845 ) , .A1( us33_n860 ) , .C1( us33_n863 ) , .B2( us33_n870 ) );
  NOR2_X1 us33_U220 (.ZN( us33_n531 ) , .A2( us33_n780 ) , .A1( us33_n816 ) );
  INV_X1 us33_U221 (.A( us33_n792 ) , .ZN( us33_n851 ) );
  NOR2_X1 us33_U222 (.A2( us33_n708 ) , .A1( us33_n750 ) , .ZN( us33_n771 ) );
  NOR2_X1 us33_U223 (.ZN( us33_n599 ) , .A2( us33_n791 ) , .A1( us33_n816 ) );
  NOR2_X1 us33_U224 (.A1( us33_n669 ) , .ZN( us33_n766 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U225 (.ZN( us33_n601 ) , .A2( us33_n780 ) , .A1( us33_n803 ) );
  NOR2_X1 us33_U226 (.A1( us33_n699 ) , .ZN( us33_n768 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U227 (.ZN( us33_n541 ) , .A2( us33_n697 ) , .A1( us33_n699 ) );
  NOR2_X1 us33_U228 (.ZN( us33_n527 ) , .A1( us33_n669 ) , .A2( us33_n779 ) );
  NOR2_X1 us33_U229 (.ZN( us33_n667 ) , .A1( us33_n750 ) , .A2( us33_n815 ) );
  INV_X1 us33_U23 (.A( us33_n647 ) , .ZN( us33_n870 ) );
  NOR2_X1 us33_U230 (.ZN( us33_n555 ) , .A1( us33_n750 ) , .A2( us33_n791 ) );
  NOR2_X1 us33_U231 (.ZN( us33_n508 ) , .A2( us33_n780 ) , .A1( us33_n785 ) );
  NOR2_X1 us33_U232 (.ZN( us33_n543 ) , .A2( us33_n708 ) , .A1( us33_n785 ) );
  NOR2_X1 us33_U233 (.ZN( us33_n528 ) , .A2( us33_n724 ) , .A1( us33_n803 ) );
  NOR2_X1 us33_U234 (.ZN( us33_n664 ) , .A1( us33_n785 ) , .A2( us33_n791 ) );
  NOR2_X1 us33_U235 (.ZN( us33_n556 ) , .A1( us33_n762 ) , .A2( us33_n805 ) );
  INV_X1 us33_U236 (.A( us33_n806 ) , .ZN( us33_n841 ) );
  NOR2_X1 us33_U237 (.ZN( us33_n661 ) , .A1( us33_n729 ) , .A2( us33_n790 ) );
  OAI22_X1 us33_U238 (.B1( us33_n440 ) , .ZN( us33_n444 ) , .A2( us33_n728 ) , .A1( us33_n744 ) , .B2( us33_n749 ) );
  NOR3_X1 us33_U239 (.ZN( us33_n440 ) , .A2( us33_n836 ) , .A3( us33_n837 ) , .A1( us33_n846 ) );
  NOR4_X1 us33_U24 (.ZN( us33_n473 ) , .A2( us33_n521 ) , .A4( us33_n594 ) , .A1( us33_n609 ) , .A3( us33_n629 ) );
  NOR2_X1 us33_U240 (.ZN( us33_n507 ) , .A1( us33_n812 ) , .A2( us33_n817 ) );
  NOR2_X1 us33_U241 (.ZN( us33_n557 ) , .A1( us33_n792 ) , .A2( us33_n814 ) );
  NOR2_X1 us33_U242 (.ZN( us33_n545 ) , .A1( us33_n749 ) , .A2( us33_n814 ) );
  NOR2_X1 us33_U243 (.ZN( us33_n509 ) , .A1( us33_n729 ) , .A2( us33_n779 ) );
  NOR2_X1 us33_U244 (.ZN( us33_n662 ) , .A2( us33_n697 ) , .A1( us33_n729 ) );
  OAI22_X1 us33_U245 (.B2( us33_n750 ) , .B1( us33_n751 ) , .A1( us33_n752 ) , .ZN( us33_n756 ) , .A2( us33_n806 ) );
  NOR2_X1 us33_U246 (.ZN( us33_n751 ) , .A2( us33_n852 ) , .A1( us33_n860 ) );
  NOR3_X1 us33_U247 (.ZN( us33_n752 ) , .A2( us33_n853 ) , .A1( us33_n863 ) , .A3( us33_n865 ) );
  NOR2_X1 us33_U248 (.ZN( us33_n544 ) , .A2( us33_n785 ) , .A1( us33_n792 ) );
  NOR2_X1 us33_U249 (.ZN( us33_n663 ) , .A1( us33_n729 ) , .A2( us33_n785 ) );
  NOR4_X1 us33_U25 (.ZN( us33_n479 ) , .A1( us33_n520 ) , .A4( us33_n557 ) , .A3( us33_n582 ) , .A2( us33_n630 ) );
  NOR2_X1 us33_U250 (.ZN( us33_n530 ) , .A2( us33_n744 ) , .A1( us33_n792 ) );
  NOR2_X1 us33_U251 (.ZN( us33_n506 ) , .A2( us33_n728 ) , .A1( us33_n762 ) );
  NOR2_X1 us33_U252 (.ZN( us33_n631 ) , .A1( us33_n724 ) , .A2( us33_n813 ) );
  NOR2_X1 us33_U253 (.ZN( us33_n614 ) , .A1( us33_n762 ) , .A2( us33_n812 ) );
  NOR2_X1 us33_U254 (.A1( us33_n749 ) , .ZN( us33_n767 ) , .A2( us33_n803 ) );
  NOR2_X1 us33_U255 (.ZN( us33_n516 ) , .A1( us33_n708 ) , .A2( us33_n744 ) );
  NOR2_X1 us33_U256 (.ZN( us33_n670 ) , .A1( us33_n790 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U257 (.ZN( us33_n558 ) , .A1( us33_n708 ) , .A2( us33_n816 ) );
  NOR2_X1 us33_U258 (.A2( us33_n697 ) , .ZN( us33_n716 ) , .A1( us33_n792 ) );
  NOR2_X1 us33_U259 (.ZN( us33_n517 ) , .A1( us33_n708 ) , .A2( us33_n803 ) );
  NOR4_X1 us33_U26 (.A4( us33_n532 ) , .A3( us33_n533 ) , .A2( us33_n534 ) , .ZN( us33_n535 ) , .A1( us33_n820 ) );
  NOR2_X1 us33_U260 (.ZN( us33_n521 ) , .A1( us33_n790 ) , .A2( us33_n812 ) );
  NOR2_X1 us33_U261 (.ZN( us33_n630 ) , .A1( us33_n747 ) , .A2( us33_n815 ) );
  NOR2_X1 us33_U262 (.ZN( us33_n655 ) , .A1( us33_n790 ) , .A2( us33_n815 ) );
  INV_X1 us33_U263 (.A( us33_n763 ) , .ZN( us33_n866 ) );
  AOI21_X1 us33_U264 (.ZN( us33_n552 ) , .B1( us33_n669 ) , .A( us33_n697 ) , .B2( us33_n805 ) );
  NOR2_X1 us33_U265 (.ZN( us33_n668 ) , .A2( us33_n708 ) , .A1( us33_n790 ) );
  NOR2_X1 us33_U266 (.ZN( us33_n542 ) , .A1( us33_n762 ) , .A2( us33_n791 ) );
  NOR2_X1 us33_U267 (.ZN( us33_n656 ) , .A1( us33_n747 ) , .A2( us33_n780 ) );
  NOR2_X1 us33_U268 (.ZN( us33_n609 ) , .A2( us33_n724 ) , .A1( us33_n817 ) );
  INV_X1 us33_U269 (.A( us33_n729 ) , .ZN( us33_n868 ) );
  NOR4_X1 us33_U27 (.ZN( us33_n456 ) , .A2( us33_n517 ) , .A1( us33_n543 ) , .A3( us33_n579 ) , .A4( us33_n615 ) );
  AOI21_X1 us33_U270 (.B1( us33_n625 ) , .ZN( us33_n627 ) , .A( us33_n763 ) , .B2( us33_n814 ) );
  AOI21_X1 us33_U271 (.ZN( us33_n650 ) , .A( us33_n779 ) , .B1( us33_n792 ) , .B2( us33_n805 ) );
  AOI21_X1 us33_U272 (.A( us33_n815 ) , .B2( us33_n816 ) , .B1( us33_n817 ) , .ZN( us33_n818 ) );
  NOR2_X1 us33_U273 (.ZN( us33_n579 ) , .A2( us33_n708 ) , .A1( us33_n730 ) );
  NOR2_X1 us33_U274 (.ZN( us33_n533 ) , .A2( us33_n724 ) , .A1( us33_n730 ) );
  NOR2_X1 us33_U275 (.ZN( us33_n642 ) , .A2( us33_n788 ) , .A1( us33_n791 ) );
  AOI21_X1 us33_U276 (.A( us33_n812 ) , .B2( us33_n813 ) , .B1( us33_n814 ) , .ZN( us33_n819 ) );
  NOR2_X1 us33_U277 (.A2( us33_n708 ) , .A1( us33_n762 ) , .ZN( us33_n794 ) );
  NOR2_X1 us33_U278 (.A2( us33_n697 ) , .A1( us33_n780 ) , .ZN( us33_n820 ) );
  AOI21_X1 us33_U279 (.ZN( us33_n626 ) , .B2( us33_n669 ) , .A( us33_n790 ) , .B1( us33_n791 ) );
  NOR4_X1 us33_U28 (.A4( us33_n541 ) , .A3( us33_n542 ) , .A2( us33_n543 ) , .ZN( us33_n550 ) , .A1( us33_n688 ) );
  AOI21_X1 us33_U280 (.ZN( us33_n499 ) , .B1( us33_n680 ) , .A( us33_n812 ) , .B2( us33_n816 ) );
  NOR2_X1 us33_U281 (.ZN( us33_n520 ) , .A2( us33_n708 ) , .A1( us33_n814 ) );
  AOI21_X1 us33_U282 (.ZN( us33_n477 ) , .A( us33_n669 ) , .B1( us33_n750 ) , .B2( us33_n806 ) );
  NOR2_X1 us33_U283 (.ZN( us33_n582 ) , .A1( us33_n744 ) , .A2( us33_n815 ) );
  AOI21_X1 us33_U284 (.ZN( us33_n593 ) , .B1( us33_n750 ) , .A( us33_n792 ) , .B2( us33_n813 ) );
  AOI21_X1 us33_U285 (.ZN( us33_n515 ) , .A( us33_n729 ) , .B1( us33_n750 ) , .B2( us33_n803 ) );
  NOR2_X1 us33_U286 (.A1( us33_n697 ) , .ZN( us33_n770 ) , .A2( us33_n815 ) );
  AOI21_X1 us33_U287 (.ZN( us33_n510 ) , .B2( us33_n669 ) , .A( us33_n730 ) , .B1( us33_n815 ) );
  NOR2_X1 us33_U288 (.ZN( us33_n519 ) , .A2( us33_n699 ) , .A1( us33_n816 ) );
  NOR2_X1 us33_U289 (.ZN( us33_n559 ) , .A2( us33_n791 ) , .A1( us33_n803 ) );
  AOI221_X1 us33_U29 (.A( us33_n713 ) , .B2( us33_n714 ) , .ZN( us33_n720 ) , .C1( us33_n832 ) , .B1( us33_n839 ) , .C2( us33_n863 ) );
  NOR2_X1 us33_U290 (.ZN( us33_n581 ) , .A1( us33_n669 ) , .A2( us33_n788 ) );
  INV_X1 us33_U291 (.A( us33_n813 ) , .ZN( us33_n836 ) );
  NOR2_X1 us33_U292 (.ZN( us33_n683 ) , .A2( us33_n699 ) , .A1( us33_n803 ) );
  AOI21_X1 us33_U293 (.ZN( us33_n589 ) , .B2( us33_n699 ) , .B1( us33_n815 ) , .A( us33_n817 ) );
  AOI21_X1 us33_U294 (.ZN( us33_n539 ) , .B2( us33_n812 ) , .A( us33_n814 ) , .B1( us33_n815 ) );
  AOI21_X1 us33_U295 (.ZN( us33_n540 ) , .A( us33_n763 ) , .B2( us33_n779 ) , .B1( us33_n817 ) );
  AOI21_X1 us33_U296 (.B1( us33_n699 ) , .ZN( us33_n700 ) , .A( us33_n732 ) , .B2( us33_n763 ) );
  AOI21_X1 us33_U297 (.ZN( us33_n591 ) , .B2( us33_n763 ) , .A( us33_n785 ) , .B1( us33_n812 ) );
  AOI21_X1 us33_U298 (.ZN( us33_n498 ) , .A( us33_n724 ) , .B2( us33_n762 ) , .B1( us33_n814 ) );
  NOR2_X1 us33_U299 (.ZN( us33_n547 ) , .A1( us33_n699 ) , .A2( us33_n744 ) );
  NAND2_X1 us33_U3 (.A1( us33_n441 ) , .A2( us33_n464 ) , .ZN( us33_n708 ) );
  OR2_X1 us33_U30 (.A2( us33_n711 ) , .A1( us33_n712 ) , .ZN( us33_n713 ) );
  INV_X1 us33_U300 (.A( us33_n791 ) , .ZN( us33_n873 ) );
  AOI21_X1 us33_U301 (.ZN( us33_n649 ) , .B1( us33_n729 ) , .B2( us33_n763 ) , .A( us33_n813 ) );
  NOR2_X1 us33_U302 (.ZN( us33_n685 ) , .A1( us33_n729 ) , .A2( us33_n816 ) );
  AOI21_X1 us33_U303 (.B1( us33_n686 ) , .ZN( us33_n687 ) , .A( us33_n728 ) , .B2( us33_n761 ) );
  AOI21_X1 us33_U304 (.ZN( us33_n569 ) , .B1( us33_n750 ) , .B2( us33_n762 ) , .A( us33_n780 ) );
  AOI21_X1 us33_U305 (.ZN( us33_n571 ) , .B2( us33_n697 ) , .B1( us33_n806 ) , .A( us33_n812 ) );
  NOR2_X1 us33_U306 (.ZN( us33_n568 ) , .A1( us33_n729 ) , .A2( us33_n762 ) );
  NOR2_X1 us33_U307 (.ZN( us33_n566 ) , .A2( us33_n697 ) , .A1( us33_n763 ) );
  AOI21_X1 us33_U308 (.ZN( us33_n640 ) , .B2( us33_n747 ) , .A( us33_n792 ) , .B1( us33_n803 ) );
  INV_X1 us33_U309 (.A( us33_n699 ) , .ZN( us33_n853 ) );
  NOR2_X1 us33_U31 (.ZN( us33_n680 ) , .A2( us33_n834 ) , .A1( us33_n839 ) );
  AOI21_X1 us33_U310 (.ZN( us33_n514 ) , .A( us33_n779 ) , .B2( us33_n792 ) , .B1( us33_n812 ) );
  AOI21_X1 us33_U311 (.ZN( us33_n639 ) , .B2( us33_n749 ) , .A( us33_n788 ) , .B1( us33_n812 ) );
  NAND2_X1 us33_U312 (.ZN( us33_n753 ) , .A1( us33_n763 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U313 (.ZN( us33_n665 ) , .A1( us33_n780 ) , .A2( us33_n813 ) );
  AOI21_X1 us33_U314 (.ZN( us33_n564 ) , .B1( us33_n724 ) , .A( us33_n779 ) , .B2( us33_n791 ) );
  AOI21_X1 us33_U315 (.ZN( us33_n497 ) , .A( us33_n779 ) , .B2( us33_n791 ) , .B1( us33_n804 ) );
  AOI21_X1 us33_U316 (.ZN( us33_n689 ) , .B2( us33_n749 ) , .B1( us33_n763 ) , .A( us33_n806 ) );
  AOI21_X1 us33_U317 (.ZN( us33_n450 ) , .B2( us33_n792 ) , .A( us33_n803 ) , .B1( us33_n815 ) );
  NOR2_X1 us33_U318 (.ZN( us33_n567 ) , .A1( us33_n747 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U319 (.ZN( us33_n529 ) , .A1( us33_n708 ) , .A2( us33_n779 ) );
  AOI222_X1 us33_U32 (.ZN( us33_n469 ) , .B1( us33_n832 ) , .A1( us33_n839 ) , .C1( us33_n842 ) , .C2( us33_n851 ) , .A2( us33_n855 ) , .B2( us33_n865 ) );
  NOR2_X1 us33_U320 (.ZN( us33_n578 ) , .A1( us33_n708 ) , .A2( us33_n813 ) );
  AOI21_X1 us33_U321 (.ZN( us33_n478 ) , .B2( us33_n697 ) , .A( us33_n749 ) , .B1( us33_n779 ) );
  AOI21_X1 us33_U322 (.A( us33_n790 ) , .B2( us33_n791 ) , .B1( us33_n792 ) , .ZN( us33_n793 ) );
  NOR2_X1 us33_U323 (.ZN( us33_n684 ) , .A1( us33_n791 ) , .A2( us33_n813 ) );
  AOI21_X1 us33_U324 (.A( us33_n733 ) , .ZN( us33_n734 ) , .B2( us33_n780 ) , .B1( us33_n792 ) );
  NOR2_X1 us33_U325 (.A2( us33_n813 ) , .A1( us33_n815 ) , .ZN( us33_n821 ) );
  AOI21_X1 us33_U326 (.ZN( us33_n641 ) , .B1( us33_n680 ) , .A( us33_n791 ) , .B2( us33_n817 ) );
  NOR2_X1 us33_U327 (.ZN( us33_n711 ) , .A1( us33_n762 ) , .A2( us33_n763 ) );
  NOR2_X1 us33_U328 (.ZN( us33_n583 ) , .A1( us33_n792 ) , .A2( us33_n817 ) );
  NOR2_X1 us33_U329 (.ZN( us33_n534 ) , .A1( us33_n724 ) , .A2( us33_n788 ) );
  NOR4_X1 us33_U33 (.A1( us33_n466 ) , .ZN( us33_n467 ) , .A4( us33_n542 ) , .A2( us33_n554 ) , .A3( us33_n614 ) );
  NOR2_X1 us33_U330 (.ZN( us33_n632 ) , .A2( us33_n697 ) , .A1( us33_n724 ) );
  NOR2_X1 us33_U331 (.ZN( us33_n682 ) , .A2( us33_n708 ) , .A1( us33_n817 ) );
  NOR2_X1 us33_U332 (.ZN( us33_n580 ) , .A2( us33_n697 ) , .A1( us33_n791 ) );
  INV_X1 us33_U333 (.A( us33_n815 ) , .ZN( us33_n855 ) );
  AOI21_X1 us33_U334 (.ZN( us33_n442 ) , .A( us33_n699 ) , .B1( us33_n733 ) , .B2( us33_n750 ) );
  INV_X1 us33_U335 (.A( us33_n780 ) , .ZN( us33_n850 ) );
  INV_X1 us33_U336 (.A( us33_n785 ) , .ZN( us33_n846 ) );
  NAND2_X1 us33_U337 (.ZN( us33_n714 ) , .A1( us33_n728 ) , .A2( us33_n780 ) );
  NAND2_X1 us33_U338 (.A2( us33_n762 ) , .A1( us33_n806 ) , .ZN( us33_n810 ) );
  AOI21_X1 us33_U339 (.ZN( us33_n443 ) , .B1( us33_n789 ) , .B2( us33_n791 ) , .A( us33_n814 ) );
  AOI221_X1 us33_U34 (.ZN( us33_n468 ) , .C2( us33_n714 ) , .B2( us33_n831 ) , .C1( us33_n845 ) , .B1( us33_n860 ) , .A( us33_n864 ) );
  NAND2_X1 us33_U340 (.ZN( us33_n671 ) , .A1( us33_n806 ) , .A2( us33_n816 ) );
  NOR2_X1 us33_U341 (.ZN( us33_n484 ) , .A1( us33_n788 ) , .A2( us33_n805 ) );
  NOR2_X1 us33_U342 (.ZN( us33_n470 ) , .A2( us33_n779 ) , .A1( us33_n815 ) );
  NOR2_X1 us33_U343 (.ZN( us33_n712 ) , .A2( us33_n724 ) , .A1( us33_n790 ) );
  OAI21_X1 us33_U344 (.A( us33_n787 ) , .B2( us33_n788 ) , .B1( us33_n789 ) , .ZN( us33_n795 ) );
  OAI21_X1 us33_U345 (.ZN( us33_n787 ) , .A( us33_n839 ) , .B1( us33_n863 ) , .B2( us33_n873 ) );
  NOR2_X1 us33_U346 (.ZN( us33_n526 ) , .A1( us33_n724 ) , .A2( us33_n750 ) );
  NAND2_X1 us33_U347 (.A1( us33_n699 ) , .A2( us33_n729 ) , .ZN( us33_n782 ) );
  NOR2_X1 us33_U348 (.ZN( us33_n518 ) , .A1( us33_n708 ) , .A2( us33_n788 ) );
  OAI21_X1 us33_U349 (.A( us33_n698 ) , .ZN( us33_n702 ) , .B2( us33_n750 ) , .B1( us33_n804 ) );
  NOR4_X1 us33_U35 (.A4( us33_n514 ) , .A3( us33_n515 ) , .A2( us33_n516 ) , .A1( us33_n517 ) , .ZN( us33_n524 ) );
  OAI21_X1 us33_U350 (.ZN( us33_n698 ) , .B2( us33_n833 ) , .B1( us33_n838 ) , .A( us33_n860 ) );
  OAI21_X1 us33_U351 (.A( us33_n731 ) , .B1( us33_n732 ) , .ZN( us33_n736 ) , .B2( us33_n805 ) );
  OAI21_X1 us33_U352 (.ZN( us33_n731 ) , .A( us33_n833 ) , .B2( us33_n852 ) , .B1( us33_n873 ) );
  INV_X1 us33_U353 (.A( us33_n817 ) , .ZN( us33_n844 ) );
  INV_X1 us33_U354 (.A( us33_n724 ) , .ZN( us33_n856 ) );
  AND2_X1 us33_U355 (.ZN( us33_n732 ) , .A1( us33_n779 ) , .A2( us33_n785 ) );
  NAND2_X1 us33_U356 (.A1( us33_n447 ) , .A2( us33_n449 ) , .ZN( us33_n805 ) );
  NAND2_X1 us33_U357 (.A1( us33_n451 ) , .A2( us33_n454 ) , .ZN( us33_n814 ) );
  NAND2_X1 us33_U358 (.A1( us33_n452 ) , .A2( us33_n465 ) , .ZN( us33_n669 ) );
  NAND2_X1 us33_U359 (.A2( us33_n448 ) , .A1( us33_n460 ) , .ZN( us33_n728 ) );
  AOI222_X1 us33_U36 (.ZN( us33_n525 ) , .A1( us33_n834 ) , .B2( us33_n837 ) , .C1( us33_n844 ) , .C2( us33_n850 ) , .A2( us33_n852 ) , .B1( us33_n866 ) );
  NAND2_X1 us33_U360 (.A1( us33_n455 ) , .A2( us33_n462 ) , .ZN( us33_n750 ) );
  NAND2_X1 us33_U361 (.A2( us33_n453 ) , .A1( us33_n455 ) , .ZN( us33_n806 ) );
  NAND2_X1 us33_U362 (.A1( us33_n451 ) , .A2( us33_n471 ) , .ZN( us33_n816 ) );
  NAND2_X1 us33_U363 (.A1( us33_n454 ) , .A2( us33_n461 ) , .ZN( us33_n813 ) );
  NAND2_X1 us33_U364 (.A1( us33_n455 ) , .A2( us33_n471 ) , .ZN( us33_n803 ) );
  NAND2_X1 us33_U365 (.A1( us33_n453 ) , .A2( us33_n461 ) , .ZN( us33_n744 ) );
  NAND2_X1 us33_U366 (.A1( us33_n453 ) , .A2( us33_n472 ) , .ZN( us33_n785 ) );
  NAND2_X1 us33_U367 (.A2( us33_n454 ) , .A1( us33_n472 ) , .ZN( us33_n779 ) );
  NAND2_X1 us33_U368 (.A2( us33_n464 ) , .A1( us33_n465 ) , .ZN( us33_n812 ) );
  NAND2_X1 us33_U369 (.A1( us33_n441 ) , .A2( us33_n460 ) , .ZN( us33_n699 ) );
  NOR4_X1 us33_U37 (.A3( us33_n521 ) , .A1( us33_n522 ) , .ZN( us33_n523 ) , .A2( us33_n673 ) , .A4( us33_n769 ) );
  NAND2_X1 us33_U370 (.A2( us33_n449 ) , .A1( us33_n452 ) , .ZN( us33_n763 ) );
  NAND2_X1 us33_U371 (.A2( us33_n448 ) , .A1( us33_n452 ) , .ZN( us33_n729 ) );
  NAND2_X1 us33_U372 (.A2( us33_n461 ) , .A1( us33_n462 ) , .ZN( us33_n747 ) );
  NAND2_X1 us33_U373 (.A1( us33_n462 ) , .A2( us33_n472 ) , .ZN( us33_n788 ) );
  NOR2_X1 us33_U374 (.ZN( us33_n465 ) , .A2( us33_n847 ) , .A1( us33_n848 ) );
  NOR2_X1 us33_U375 (.ZN( us33_n453 ) , .A1( us33_n826 ) , .A2( us33_n827 ) );
  NOR2_X1 us33_U376 (.ZN( us33_n451 ) , .A1( us33_n828 ) , .A2( us33_n829 ) );
  NAND2_X1 us33_U377 (.A1( us33_n451 ) , .A2( us33_n462 ) , .ZN( us33_n790 ) );
  NAND2_X2 us33_U378 (.A2( us33_n448 ) , .A1( us33_n464 ) , .ZN( us33_n815 ) );
  NAND2_X1 us33_U379 (.A2( us33_n441 ) , .A1( us33_n447 ) , .ZN( us33_n784 ) );
  AOI221_X1 us33_U38 (.A( us33_n781 ) , .ZN( us33_n798 ) , .C2( us33_n837 ) , .B2( us33_n838 ) , .B1( us33_n865 ) , .C1( us33_n866 ) );
  NAND2_X1 us33_U380 (.A2( us33_n454 ) , .A1( us33_n455 ) , .ZN( us33_n730 ) );
  NAND2_X2 us33_U381 (.A1( us33_n449 ) , .A2( us33_n464 ) , .ZN( us33_n724 ) );
  NAND2_X2 us33_U382 (.A1( us33_n449 ) , .A2( us33_n460 ) , .ZN( us33_n792 ) );
  NAND2_X2 us33_U383 (.A2( us33_n460 ) , .A1( us33_n465 ) , .ZN( us33_n780 ) );
  NOR2_X1 us33_U384 (.ZN( us33_n447 ) , .A2( us33_n849 ) , .A1( us33_n858 ) );
  NAND2_X1 us33_U385 (.A1( us33_n447 ) , .A2( us33_n448 ) , .ZN( us33_n786 ) );
  NOR2_X1 us33_U386 (.A2( sa33_6 ) , .A1( sa33_7 ) , .ZN( us33_n464 ) );
  NOR2_X1 us33_U387 (.A2( sa33_7 ) , .ZN( us33_n460 ) , .A1( us33_n849 ) );
  NOR2_X1 us33_U388 (.A2( sa33_4 ) , .ZN( us33_n449 ) , .A1( us33_n848 ) );
  NOR2_X1 us33_U389 (.A2( sa33_4 ) , .A1( sa33_5 ) , .ZN( us33_n441 ) );
  NOR4_X1 us33_U39 (.A4( us33_n793 ) , .A3( us33_n794 ) , .A2( us33_n795 ) , .A1( us33_n796 ) , .ZN( us33_n797 ) );
  NOR2_X1 us33_U390 (.A2( sa33_5 ) , .ZN( us33_n448 ) , .A1( us33_n847 ) );
  NOR2_X1 us33_U391 (.A2( sa33_2 ) , .A1( sa33_3 ) , .ZN( us33_n472 ) );
  NOR2_X1 us33_U392 (.A2( sa33_6 ) , .ZN( us33_n452 ) , .A1( us33_n858 ) );
  NOR2_X1 us33_U393 (.A2( sa33_1 ) , .ZN( us33_n471 ) , .A1( us33_n826 ) );
  NOR2_X1 us33_U394 (.A2( sa33_0 ) , .ZN( us33_n454 ) , .A1( us33_n827 ) );
  NOR2_X1 us33_U395 (.A2( sa33_0 ) , .A1( sa33_1 ) , .ZN( us33_n462 ) );
  NOR2_X1 us33_U396 (.A2( sa33_3 ) , .ZN( us33_n455 ) , .A1( us33_n828 ) );
  NOR2_X1 us33_U397 (.A2( sa33_2 ) , .ZN( us33_n461 ) , .A1( us33_n829 ) );
  INV_X1 us33_U398 (.A( sa33_6 ) , .ZN( us33_n849 ) );
  INV_X1 us33_U399 (.A( sa33_4 ) , .ZN( us33_n847 ) );
  NAND2_X1 us33_U4 (.A2( us33_n441 ) , .A1( us33_n452 ) , .ZN( us33_n791 ) );
  NOR4_X1 us33_U40 (.A4( us33_n776 ) , .A3( us33_n777 ) , .A1( us33_n778 ) , .ZN( us33_n799 ) , .A2( us33_n801 ) );
  INV_X1 us33_U400 (.A( sa33_3 ) , .ZN( us33_n829 ) );
  INV_X1 us33_U401 (.A( sa33_1 ) , .ZN( us33_n827 ) );
  INV_X1 us33_U402 (.A( sa33_0 ) , .ZN( us33_n826 ) );
  INV_X1 us33_U403 (.A( sa33_2 ) , .ZN( us33_n828 ) );
  INV_X1 us33_U404 (.A( sa33_7 ) , .ZN( us33_n858 ) );
  INV_X1 us33_U405 (.A( sa33_5 ) , .ZN( us33_n848 ) );
  NAND2_X1 us33_U406 (.A2( us33_n461 ) , .A1( us33_n471 ) , .ZN( us33_n697 ) );
  OAI221_X1 us33_U407 (.A( us33_n783 ) , .C2( us33_n784 ) , .B2( us33_n785 ) , .B1( us33_n786 ) , .ZN( us33_n796 ) , .C1( us33_n813 ) );
  NAND2_X1 us33_U408 (.A1( us33_n729 ) , .A2( us33_n784 ) , .ZN( us33_n811 ) );
  OAI22_X1 us33_U409 (.ZN( us33_n588 ) , .A2( us33_n747 ) , .B2( us33_n762 ) , .A1( us33_n763 ) , .B1( us33_n784 ) );
  NOR4_X1 us33_U41 (.A3( us33_n755 ) , .A2( us33_n756 ) , .A1( us33_n757 ) , .ZN( us33_n758 ) , .A4( us33_n869 ) );
  AOI21_X1 us33_U410 (.ZN( us33_n592 ) , .B1( us33_n728 ) , .B2( us33_n784 ) , .A( us33_n790 ) );
  AOI21_X1 us33_U411 (.ZN( us33_n623 ) , .B1( us33_n699 ) , .A( us33_n779 ) , .B2( us33_n784 ) );
  AOI21_X1 us33_U412 (.ZN( us33_n648 ) , .A( us33_n762 ) , .B2( us33_n784 ) , .B1( us33_n792 ) );
  OAI22_X1 us33_U413 (.ZN( us33_n681 ) , .A1( us33_n699 ) , .A2( us33_n730 ) , .B2( us33_n784 ) , .B1( us33_n817 ) );
  OAI21_X1 us33_U414 (.A( us33_n613 ) , .ZN( us33_n616 ) , .B1( us33_n625 ) , .B2( us33_n784 ) );
  NOR2_X1 us33_U415 (.ZN( us33_n610 ) , .A1( us33_n784 ) , .A2( us33_n816 ) );
  OAI222_X1 us33_U416 (.A2( us33_n669 ) , .ZN( us33_n674 ) , .B1( us33_n747 ) , .B2( us33_n784 ) , .C2( us33_n788 ) , .C1( us33_n815 ) , .A1( us33_n817 ) );
  NOR2_X1 us33_U417 (.ZN( us33_n651 ) , .A1( us33_n784 ) , .A2( us33_n788 ) );
  NOR2_X1 us33_U418 (.ZN( us33_n600 ) , .A2( us33_n697 ) , .A1( us33_n784 ) );
  NOR2_X1 us33_U419 (.ZN( us33_n553 ) , .A2( us33_n744 ) , .A1( us33_n784 ) );
  AOI211_X1 us33_U42 (.B( us33_n745 ) , .A( us33_n746 ) , .ZN( us33_n759 ) , .C1( us33_n832 ) , .C2( us33_n853 ) );
  INV_X1 us33_U420 (.A( us33_n784 ) , .ZN( us33_n861 ) );
  AOI21_X1 us33_U421 (.ZN( us33_n500 ) , .A( us33_n697 ) , .B1( us33_n708 ) , .B2( us33_n786 ) );
  OAI221_X1 us33_U422 (.A( us33_n696 ) , .ZN( us33_n703 ) , .C2( us33_n784 ) , .C1( us33_n785 ) , .B1( us33_n786 ) , .B2( us33_n806 ) );
  OAI22_X1 us33_U423 (.ZN( us33_n590 ) , .B1( us33_n730 ) , .B2( us33_n749 ) , .A2( us33_n786 ) , .A1( us33_n803 ) );
  NOR2_X1 us33_U424 (.ZN( us33_n612 ) , .A1( us33_n779 ) , .A2( us33_n786 ) );
  NAND2_X1 us33_U425 (.A2( us33_n749 ) , .A1( us33_n786 ) , .ZN( us33_n809 ) );
  OAI222_X1 us33_U426 (.ZN( us33_n617 ) , .B1( us33_n697 ) , .C1( us33_n724 ) , .C2( us33_n747 ) , .B2( us33_n786 ) , .A2( us33_n792 ) , .A1( us33_n816 ) );
  NOR2_X1 us33_U427 (.ZN( us33_n717 ) , .A2( us33_n744 ) , .A1( us33_n786 ) );
  NOR2_X1 us33_U428 (.ZN( us33_n653 ) , .A1( us33_n762 ) , .A2( us33_n786 ) );
  NOR2_X1 us33_U429 (.ZN( us33_n554 ) , .A1( us33_n786 ) , .A2( us33_n813 ) );
  NOR3_X1 us33_U43 (.A3( us33_n741 ) , .A2( us33_n742 ) , .A1( us33_n743 ) , .ZN( us33_n760 ) );
  NOR2_X1 us33_U430 (.ZN( us33_n701 ) , .A2( us33_n786 ) , .A1( us33_n817 ) );
  NOR2_X1 us33_U431 (.A1( us33_n730 ) , .ZN( us33_n765 ) , .A2( us33_n786 ) );
  AND2_X1 us33_U432 (.ZN( us33_n438 ) , .A2( us33_n831 ) , .A1( us33_n854 ) );
  AND2_X1 us33_U433 (.ZN( us33_n439 ) , .A2( us33_n843 ) , .A1( us33_n861 ) );
  NOR3_X1 us33_U434 (.A1( us33_n438 ) , .A2( us33_n439 ) , .A3( us33_n576 ) , .ZN( us33_n587 ) );
  NAND4_X1 us33_U435 (.ZN( sa30_sr_2 ) , .A4( us33_n643 ) , .A3( us33_n644 ) , .A2( us33_n645 ) , .A1( us33_n646 ) );
  INV_X1 us33_U436 (.A( us33_n812 ) , .ZN( us33_n854 ) );
  NAND3_X1 us33_U437 (.ZN( sa30_sr_6 ) , .A3( us33_n797 ) , .A2( us33_n798 ) , .A1( us33_n799 ) );
  NAND3_X1 us33_U438 (.ZN( sa30_sr_5 ) , .A3( us33_n758 ) , .A2( us33_n759 ) , .A1( us33_n760 ) );
  NAND3_X1 us33_U439 (.ZN( sa30_sr_4 ) , .A3( us33_n738 ) , .A2( us33_n739 ) , .A1( us33_n740 ) );
  NAND4_X1 us33_U44 (.ZN( sa30_sr_3 ) , .A4( us33_n704 ) , .A3( us33_n705 ) , .A2( us33_n706 ) , .A1( us33_n707 ) );
  NAND3_X1 us33_U440 (.A3( us33_n675 ) , .A2( us33_n676 ) , .A1( us33_n677 ) , .ZN( us33_n807 ) );
  NAND3_X1 us33_U441 (.ZN( us33_n638 ) , .A3( us33_n708 ) , .A2( us33_n724 ) , .A1( us33_n792 ) );
  NAND3_X1 us33_U442 (.A3( us33_n618 ) , .A2( us33_n619 ) , .A1( us33_n620 ) , .ZN( us33_n725 ) );
  NAND3_X1 us33_U443 (.A3( us33_n585 ) , .A2( us33_n586 ) , .A1( us33_n587 ) , .ZN( us33_n621 ) );
  NAND3_X1 us33_U444 (.ZN( us33_n565 ) , .A3( us33_n680 ) , .A2( us33_n750 ) , .A1( us33_n785 ) );
  NAND3_X1 us33_U445 (.A3( us33_n523 ) , .A2( us33_n524 ) , .A1( us33_n525 ) , .ZN( us33_n742 ) );
  NAND3_X1 us33_U446 (.A3( us33_n512 ) , .A1( us33_n513 ) , .ZN( us33_n608 ) , .A2( us33_n871 ) );
  NAND3_X1 us33_U447 (.A3( us33_n467 ) , .A2( us33_n468 ) , .A1( us33_n469 ) , .ZN( us33_n777 ) );
  INV_X1 us33_U448 (.A( us33_n803 ) , .ZN( us33_n843 ) );
  AOI21_X1 us33_U449 (.ZN( us33_n576 ) , .B2( us33_n724 ) , .B1( us33_n748 ) , .A( us33_n785 ) );
  NOR4_X1 us33_U45 (.A4( us33_n700 ) , .A3( us33_n701 ) , .A2( us33_n702 ) , .A1( us33_n703 ) , .ZN( us33_n704 ) );
  AOI211_X1 us33_U46 (.B( us33_n694 ) , .A( us33_n695 ) , .ZN( us33_n705 ) , .C2( us33_n831 ) , .C1( us33_n851 ) );
  NOR2_X1 us33_U47 (.ZN( us33_n707 ) , .A2( us33_n776 ) , .A1( us33_n800 ) );
  AOI222_X1 us33_U48 (.B2( us33_n638 ) , .ZN( us33_n644 ) , .B1( us33_n841 ) , .A1( us33_n842 ) , .C2( us33_n846 ) , .C1( us33_n863 ) , .A2( us33_n865 ) );
  NOR4_X1 us33_U49 (.A4( us33_n639 ) , .A3( us33_n640 ) , .A2( us33_n641 ) , .A1( us33_n642 ) , .ZN( us33_n643 ) );
  NAND2_X1 us33_U5 (.A2( us33_n471 ) , .A1( us33_n472 ) , .ZN( us33_n817 ) );
  NOR3_X1 us33_U50 (.A2( us33_n607 ) , .A1( us33_n608 ) , .ZN( us33_n646 ) , .A3( us33_n722 ) );
  NOR2_X1 us33_U51 (.ZN( us33_n804 ) , .A1( us33_n854 ) , .A2( us33_n861 ) );
  NAND4_X1 us33_U52 (.ZN( sa30_sr_7 ) , .A4( us33_n822 ) , .A3( us33_n823 ) , .A2( us33_n824 ) , .A1( us33_n825 ) );
  NOR4_X1 us33_U53 (.A4( us33_n818 ) , .A3( us33_n819 ) , .A2( us33_n820 ) , .A1( us33_n821 ) , .ZN( us33_n822 ) );
  AOI222_X1 us33_U54 (.C2( us33_n809 ) , .B2( us33_n810 ) , .A2( us33_n811 ) , .ZN( us33_n823 ) , .C1( us33_n832 ) , .A1( us33_n839 ) , .B1( us33_n853 ) );
  AOI211_X1 us33_U55 (.B( us33_n807 ) , .A( us33_n808 ) , .ZN( us33_n824 ) , .C1( us33_n842 ) , .C2( us33_n850 ) );
  NAND4_X1 us33_U56 (.ZN( sa30_sr_0 ) , .A4( us33_n501 ) , .A3( us33_n502 ) , .A2( us33_n503 ) , .A1( us33_n504 ) );
  AOI221_X1 us33_U57 (.A( us33_n497 ) , .ZN( us33_n502 ) , .B2( us33_n843 ) , .C1( us33_n846 ) , .C2( us33_n860 ) , .B1( us33_n862 ) );
  NOR4_X1 us33_U58 (.A4( us33_n498 ) , .A3( us33_n499 ) , .A2( us33_n500 ) , .ZN( us33_n501 ) , .A1( us33_n527 ) );
  AOI211_X1 us33_U59 (.A( us33_n496 ) , .ZN( us33_n503 ) , .B( us33_n802 ) , .C2( us33_n839 ) , .C1( us33_n851 ) );
  NOR3_X1 us33_U6 (.ZN( us33_n598 ) , .A1( us33_n608 ) , .A3( us33_n723 ) , .A2( us33_n742 ) );
  NAND4_X1 us33_U60 (.ZN( sa30_sr_1 ) , .A4( us33_n595 ) , .A3( us33_n596 ) , .A2( us33_n597 ) , .A1( us33_n598 ) );
  NOR4_X1 us33_U61 (.A4( us33_n591 ) , .A3( us33_n592 ) , .A2( us33_n593 ) , .A1( us33_n594 ) , .ZN( us33_n595 ) );
  AOI211_X1 us33_U62 (.B( us33_n589 ) , .A( us33_n590 ) , .ZN( us33_n596 ) , .C2( us33_n811 ) , .C1( us33_n833 ) );
  AOI211_X1 us33_U63 (.A( us33_n588 ) , .ZN( us33_n597 ) , .B( us33_n621 ) , .C1( us33_n845 ) , .C2( us33_n855 ) );
  NOR2_X1 us33_U64 (.ZN( us33_n748 ) , .A1( us33_n861 ) , .A2( us33_n862 ) );
  NOR2_X1 us33_U65 (.ZN( us33_n625 ) , .A2( us33_n836 ) , .A1( us33_n839 ) );
  NAND4_X1 us33_U66 (.A4( us33_n603 ) , .A3( us33_n604 ) , .A2( us33_n605 ) , .A1( us33_n606 ) , .ZN( us33_n722 ) );
  NOR3_X1 us33_U67 (.A1( us33_n599 ) , .ZN( us33_n604 ) , .A3( us33_n663 ) , .A2( us33_n770 ) );
  NOR4_X1 us33_U68 (.A3( us33_n600 ) , .A2( us33_n601 ) , .A1( us33_n602 ) , .ZN( us33_n603 ) , .A4( us33_n655 ) );
  AOI222_X1 us33_U69 (.ZN( us33_n606 ) , .A1( us33_n830 ) , .C2( us33_n837 ) , .B1( us33_n842 ) , .A2( us33_n856 ) , .B2( us33_n861 ) , .C1( us33_n868 ) );
  NOR3_X1 us33_U7 (.A3( us33_n800 ) , .A2( us33_n801 ) , .A1( us33_n802 ) , .ZN( us33_n825 ) );
  NAND4_X1 us33_U70 (.A4( us33_n657 ) , .A3( us33_n658 ) , .A2( us33_n659 ) , .A1( us33_n660 ) , .ZN( us33_n800 ) );
  NOR3_X1 us33_U71 (.A3( us33_n648 ) , .A2( us33_n649 ) , .A1( us33_n650 ) , .ZN( us33_n659 ) );
  NOR3_X1 us33_U72 (.A3( us33_n651 ) , .A2( us33_n652 ) , .A1( us33_n653 ) , .ZN( us33_n658 ) );
  NOR3_X1 us33_U73 (.A3( us33_n654 ) , .A2( us33_n655 ) , .A1( us33_n656 ) , .ZN( us33_n657 ) );
  NAND4_X1 us33_U74 (.A4( us33_n560 ) , .A3( us33_n561 ) , .A2( us33_n562 ) , .A1( us33_n563 ) , .ZN( us33_n607 ) );
  NOR4_X1 us33_U75 (.ZN( us33_n561 ) , .A1( us33_n653 ) , .A3( us33_n661 ) , .A4( us33_n685 ) , .A2( us33_n768 ) );
  NOR4_X1 us33_U76 (.A4( us33_n552 ) , .A3( us33_n553 ) , .A2( us33_n554 ) , .A1( us33_n555 ) , .ZN( us33_n562 ) );
  NOR4_X1 us33_U77 (.A4( us33_n556 ) , .A3( us33_n557 ) , .A2( us33_n558 ) , .A1( us33_n559 ) , .ZN( us33_n560 ) );
  NAND4_X1 us33_U78 (.A4( us33_n772 ) , .A3( us33_n773 ) , .A2( us33_n774 ) , .A1( us33_n775 ) , .ZN( us33_n801 ) );
  NOR3_X1 us33_U79 (.A3( us33_n765 ) , .A2( us33_n766 ) , .A1( us33_n767 ) , .ZN( us33_n773 ) );
  NOR3_X1 us33_U8 (.A3( us33_n621 ) , .A2( us33_n622 ) , .ZN( us33_n636 ) , .A1( us33_n725 ) );
  NOR4_X1 us33_U80 (.A4( us33_n768 ) , .A3( us33_n769 ) , .A2( us33_n770 ) , .A1( us33_n771 ) , .ZN( us33_n772 ) );
  AOI222_X1 us33_U81 (.ZN( us33_n775 ) , .A1( us33_n830 ) , .C1( us33_n834 ) , .B2( us33_n841 ) , .A2( us33_n850 ) , .B1( us33_n861 ) , .C2( us33_n873 ) );
  NOR4_X1 us33_U82 (.A4( us33_n665 ) , .A3( us33_n666 ) , .A2( us33_n667 ) , .A1( us33_n668 ) , .ZN( us33_n676 ) );
  NOR4_X1 us33_U83 (.A4( us33_n661 ) , .A3( us33_n662 ) , .A2( us33_n663 ) , .A1( us33_n664 ) , .ZN( us33_n677 ) );
  NOR4_X1 us33_U84 (.A3( us33_n673 ) , .A1( us33_n674 ) , .ZN( us33_n675 ) , .A4( us33_n715 ) , .A2( us33_n859 ) );
  NOR2_X1 us33_U85 (.ZN( us33_n761 ) , .A1( us33_n833 ) , .A2( us33_n834 ) );
  NOR4_X1 us33_U86 (.A4( us33_n577 ) , .A3( us33_n578 ) , .A2( us33_n579 ) , .ZN( us33_n586 ) , .A1( us33_n683 ) );
  NOR4_X1 us33_U87 (.A1( us33_n584 ) , .ZN( us33_n585 ) , .A3( us33_n652 ) , .A2( us33_n662 ) , .A4( us33_n767 ) );
  AOI222_X1 us33_U88 (.ZN( us33_n513 ) , .C1( us33_n832 ) , .B2( us33_n837 ) , .A2( us33_n843 ) , .C2( us33_n862 ) , .B1( us33_n863 ) , .A1( us33_n866 ) );
  NOR4_X1 us33_U89 (.A4( us33_n509 ) , .A2( us33_n510 ) , .A1( us33_n511 ) , .ZN( us33_n512 ) , .A3( us33_n670 ) );
  NOR2_X1 us33_U9 (.ZN( us33_n575 ) , .A1( us33_n622 ) , .A2( us33_n745 ) );
  INV_X1 us33_U90 (.A( us33_n505 ) , .ZN( us33_n871 ) );
  NAND4_X1 us33_U91 (.A4( us33_n456 ) , .A3( us33_n457 ) , .A2( us33_n458 ) , .A1( us33_n459 ) , .ZN( us33_n679 ) );
  NOR3_X1 us33_U92 (.ZN( us33_n457 ) , .A3( us33_n530 ) , .A1( us33_n555 ) , .A2( us33_n570 ) );
  AOI221_X1 us33_U93 (.A( us33_n450 ) , .ZN( us33_n459 ) , .C2( us33_n753 ) , .B1( us33_n832 ) , .C1( us33_n842 ) , .B2( us33_n861 ) );
  NOR4_X1 us33_U94 (.ZN( us33_n458 ) , .A2( us33_n509 ) , .A1( us33_n599 ) , .A4( us33_n628 ) , .A3( us33_n711 ) );
  NAND4_X1 us33_U95 (.A4( us33_n535 ) , .A3( us33_n536 ) , .A2( us33_n537 ) , .A1( us33_n538 ) , .ZN( us33_n622 ) );
  NOR4_X1 us33_U96 (.A4( us33_n526 ) , .A2( us33_n527 ) , .A1( us33_n528 ) , .ZN( us33_n538 ) , .A3( us33_n701 ) );
  NOR4_X1 us33_U97 (.A1( us33_n531 ) , .ZN( us33_n536 ) , .A2( us33_n654 ) , .A4( us33_n668 ) , .A3( us33_n765 ) );
  NOR4_X1 us33_U98 (.A4( us33_n529 ) , .A3( us33_n530 ) , .ZN( us33_n537 ) , .A2( us33_n684 ) , .A1( us33_n794 ) );
  NOR2_X1 us33_U99 (.ZN( us33_n647 ) , .A1( us33_n854 ) , .A2( us33_n868 ) );
endmodule

