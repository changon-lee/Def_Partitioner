module aes_aes_die_1 ( sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa13_0, 
       sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa21_0, sa21_1, 
       sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa22_0, sa22_1, sa22_2, 
       sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa32_0, sa32_1, sa32_2, sa32_3, 
       sa32_4, sa32_5, sa32_6, sa32_7, us00_n417, us00_n425, us00_n430, us13_n447, us13_n448, 
       us13_n449, us13_n452, us13_n460, us13_n465, us13_n669, us13_n728, us13_n852, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa12_sr_0, 
        sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, sa20_sr_1, 
        sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, 
        sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
        sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7 );
  input sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa13_0, 
        sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa21_0, sa21_1, 
        sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa22_0, sa22_1, sa22_2, 
        sa22_3, sa22_4, sa22_5, sa22_6, sa22_7, sa32_0, sa32_1, sa32_2, sa32_3, 
        sa32_4, sa32_5, sa32_6, sa32_7, us00_n417, us00_n425, us00_n430, us13_n447, us13_n448, 
        us13_n449, us13_n452, us13_n460, us13_n465, us13_n669, us13_n728, us13_n852;
  output sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa12_sr_0, 
        sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa20_sr_0, sa20_sr_1, 
        sa20_sr_2, sa20_sr_3, sa20_sr_4, sa20_sr_5, sa20_sr_6, sa20_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, 
        sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
        sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7;
  wire us00_n1, us00_n10, us00_n100, us00_n101, us00_n102, us00_n103, us00_n104, us00_n105, us00_n106, 
       us00_n107, us00_n108, us00_n109, us00_n11, us00_n110, us00_n111, us00_n112, us00_n113, us00_n114, 
       us00_n115, us00_n116, us00_n117, us00_n118, us00_n119, us00_n12, us00_n120, us00_n121, us00_n122, 
       us00_n123, us00_n124, us00_n125, us00_n126, us00_n127, us00_n128, us00_n129, us00_n13, us00_n130, 
       us00_n131, us00_n132, us00_n133, us00_n134, us00_n135, us00_n136, us00_n137, us00_n138, us00_n139, 
       us00_n14, us00_n140, us00_n141, us00_n142, us00_n143, us00_n144, us00_n145, us00_n146, us00_n147, 
       us00_n148, us00_n149, us00_n15, us00_n150, us00_n151, us00_n152, us00_n153, us00_n154, us00_n155, 
       us00_n156, us00_n157, us00_n158, us00_n159, us00_n16, us00_n160, us00_n161, us00_n162, us00_n163, 
       us00_n164, us00_n165, us00_n166, us00_n167, us00_n168, us00_n169, us00_n17, us00_n170, us00_n171, 
       us00_n172, us00_n173, us00_n174, us00_n175, us00_n176, us00_n177, us00_n178, us00_n179, us00_n18, 
       us00_n180, us00_n181, us00_n182, us00_n183, us00_n184, us00_n185, us00_n186, us00_n187, us00_n188, 
       us00_n189, us00_n190, us00_n191, us00_n192, us00_n193, us00_n194, us00_n195, us00_n196, us00_n197, 
       us00_n198, us00_n199, us00_n2, us00_n20, us00_n200, us00_n201, us00_n202, us00_n203, us00_n204, 
       us00_n205, us00_n206, us00_n207, us00_n208, us00_n209, us00_n21, us00_n210, us00_n211, us00_n212, 
       us00_n213, us00_n214, us00_n215, us00_n216, us00_n217, us00_n218, us00_n219, us00_n22, us00_n220, 
       us00_n221, us00_n222, us00_n223, us00_n224, us00_n225, us00_n226, us00_n227, us00_n228, us00_n229, 
       us00_n23, us00_n230, us00_n231, us00_n232, us00_n233, us00_n234, us00_n235, us00_n236, us00_n237, 
       us00_n238, us00_n239, us00_n24, us00_n240, us00_n241, us00_n242, us00_n243, us00_n244, us00_n245, 
       us00_n246, us00_n247, us00_n248, us00_n249, us00_n25, us00_n250, us00_n251, us00_n252, us00_n253, 
       us00_n254, us00_n255, us00_n256, us00_n257, us00_n258, us00_n259, us00_n26, us00_n260, us00_n261, 
       us00_n262, us00_n263, us00_n264, us00_n265, us00_n266, us00_n267, us00_n268, us00_n269, us00_n27, 
       us00_n270, us00_n271, us00_n272, us00_n273, us00_n274, us00_n275, us00_n276, us00_n277, us00_n278, 
       us00_n279, us00_n280, us00_n281, us00_n282, us00_n283, us00_n284, us00_n285, us00_n286, us00_n287, 
       us00_n288, us00_n289, us00_n29, us00_n290, us00_n291, us00_n292, us00_n293, us00_n294, us00_n295, 
       us00_n296, us00_n297, us00_n298, us00_n299, us00_n3, us00_n30, us00_n300, us00_n301, us00_n302, 
       us00_n303, us00_n304, us00_n305, us00_n306, us00_n307, us00_n308, us00_n309, us00_n31, us00_n310, 
       us00_n311, us00_n312, us00_n313, us00_n314, us00_n315, us00_n316, us00_n317, us00_n318, us00_n319, 
       us00_n32, us00_n320, us00_n321, us00_n322, us00_n323, us00_n324, us00_n325, us00_n326, us00_n327, 
       us00_n328, us00_n329, us00_n33, us00_n330, us00_n331, us00_n332, us00_n333, us00_n334, us00_n335, 
       us00_n336, us00_n337, us00_n338, us00_n339, us00_n34, us00_n340, us00_n341, us00_n342, us00_n343, 
       us00_n344, us00_n345, us00_n346, us00_n347, us00_n348, us00_n349, us00_n35, us00_n350, us00_n351, 
       us00_n352, us00_n353, us00_n354, us00_n355, us00_n356, us00_n357, us00_n358, us00_n359, us00_n36, 
       us00_n360, us00_n361, us00_n362, us00_n363, us00_n364, us00_n365, us00_n366, us00_n367, us00_n368, 
       us00_n369, us00_n37, us00_n370, us00_n371, us00_n372, us00_n373, us00_n374, us00_n375, us00_n376, 
       us00_n377, us00_n378, us00_n379, us00_n38, us00_n380, us00_n381, us00_n382, us00_n383, us00_n384, 
       us00_n385, us00_n386, us00_n387, us00_n388, us00_n389, us00_n39, us00_n390, us00_n391, us00_n392, 
       us00_n393, us00_n394, us00_n395, us00_n396, us00_n397, us00_n398, us00_n399, us00_n4, us00_n40, 
       us00_n400, us00_n401, us00_n402, us00_n403, us00_n404, us00_n405, us00_n406, us00_n407, us00_n408, 
       us00_n409, us00_n41, us00_n410, us00_n411, us00_n412, us00_n413, us00_n414, us00_n415, us00_n416, 
       us00_n418, us00_n419, us00_n42, us00_n420, us00_n421, us00_n422, us00_n423, us00_n424, us00_n426, 
       us00_n427, us00_n428, us00_n429, us00_n43, us00_n431, us00_n432, us00_n433, us00_n434, us00_n435, 
       us00_n436, us00_n437, us00_n44, us00_n45, us00_n46, us00_n47, us00_n48, us00_n49, us00_n5, 
       us00_n50, us00_n51, us00_n52, us00_n53, us00_n54, us00_n55, us00_n56, us00_n57, us00_n58, 
       us00_n59, us00_n6, us00_n60, us00_n61, us00_n62, us00_n63, us00_n64, us00_n65, us00_n66, 
       us00_n67, us00_n68, us00_n69, us00_n7, us00_n70, us00_n71, us00_n72, us00_n73, us00_n74, 
       us00_n75, us00_n76, us00_n77, us00_n78, us00_n79, us00_n8, us00_n80, us00_n81, us00_n82, 
       us00_n83, us00_n84, us00_n85, us00_n86, us00_n87, us00_n88, us00_n89, us00_n9, us00_n90, 
       us00_n91, us00_n92, us00_n93, us00_n94, us00_n95, us00_n96, us00_n97, us00_n98, us00_n99, 
       us13_n438, us13_n439, us13_n440, us13_n441, us13_n442, us13_n443, us13_n444, us13_n445, us13_n446, 
       us13_n450, us13_n451, us13_n453, us13_n454, us13_n455, us13_n456, us13_n457, us13_n458, us13_n459, 
       us13_n461, us13_n462, us13_n463, us13_n464, us13_n466, us13_n467, us13_n468, us13_n469, us13_n470, 
       us13_n471, us13_n472, us13_n473, us13_n474, us13_n475, us13_n476, us13_n477, us13_n478, us13_n479, 
       us13_n480, us13_n481, us13_n482, us13_n483, us13_n484, us13_n485, us13_n486, us13_n487, us13_n488, 
       us13_n489, us13_n490, us13_n491, us13_n492, us13_n493, us13_n494, us13_n495, us13_n496, us13_n497, 
       us13_n498, us13_n499, us13_n500, us13_n501, us13_n502, us13_n503, us13_n504, us13_n505, us13_n506, 
       us13_n507, us13_n508, us13_n509, us13_n510, us13_n511, us13_n512, us13_n513, us13_n514, us13_n515, 
       us13_n516, us13_n517, us13_n518, us13_n519, us13_n520, us13_n521, us13_n522, us13_n523, us13_n524, 
       us13_n525, us13_n526, us13_n527, us13_n528, us13_n529, us13_n530, us13_n531, us13_n532, us13_n533, 
       us13_n534, us13_n535, us13_n536, us13_n537, us13_n538, us13_n539, us13_n540, us13_n541, us13_n542, 
       us13_n543, us13_n544, us13_n545, us13_n546, us13_n547, us13_n548, us13_n549, us13_n550, us13_n551, 
       us13_n552, us13_n553, us13_n554, us13_n555, us13_n556, us13_n557, us13_n558, us13_n559, us13_n560, 
       us13_n561, us13_n562, us13_n563, us13_n564, us13_n565, us13_n566, us13_n567, us13_n568, us13_n569, 
       us13_n570, us13_n571, us13_n572, us13_n573, us13_n574, us13_n575, us13_n576, us13_n577, us13_n578, 
       us13_n579, us13_n580, us13_n581, us13_n582, us13_n583, us13_n584, us13_n585, us13_n586, us13_n587, 
       us13_n588, us13_n589, us13_n590, us13_n591, us13_n592, us13_n593, us13_n594, us13_n595, us13_n596, 
       us13_n597, us13_n598, us13_n599, us13_n600, us13_n601, us13_n602, us13_n603, us13_n604, us13_n605, 
       us13_n606, us13_n607, us13_n608, us13_n609, us13_n610, us13_n611, us13_n612, us13_n613, us13_n614, 
       us13_n615, us13_n616, us13_n617, us13_n618, us13_n619, us13_n620, us13_n621, us13_n622, us13_n623, 
       us13_n624, us13_n625, us13_n626, us13_n627, us13_n628, us13_n629, us13_n630, us13_n631, us13_n632, 
       us13_n633, us13_n634, us13_n635, us13_n636, us13_n637, us13_n638, us13_n639, us13_n640, us13_n641, 
       us13_n642, us13_n643, us13_n644, us13_n645, us13_n646, us13_n647, us13_n648, us13_n649, us13_n650, 
       us13_n651, us13_n652, us13_n653, us13_n654, us13_n655, us13_n656, us13_n657, us13_n658, us13_n659, 
       us13_n660, us13_n661, us13_n662, us13_n663, us13_n664, us13_n665, us13_n666, us13_n667, us13_n668, 
       us13_n670, us13_n671, us13_n672, us13_n673, us13_n674, us13_n675, us13_n676, us13_n677, us13_n678, 
       us13_n679, us13_n680, us13_n681, us13_n682, us13_n683, us13_n684, us13_n685, us13_n686, us13_n687, 
       us13_n688, us13_n689, us13_n690, us13_n691, us13_n692, us13_n693, us13_n694, us13_n695, us13_n696, 
       us13_n697, us13_n698, us13_n699, us13_n700, us13_n701, us13_n702, us13_n703, us13_n704, us13_n705, 
       us13_n706, us13_n707, us13_n708, us13_n709, us13_n710, us13_n711, us13_n712, us13_n713, us13_n714, 
       us13_n715, us13_n716, us13_n717, us13_n718, us13_n719, us13_n720, us13_n721, us13_n722, us13_n723, 
       us13_n724, us13_n725, us13_n726, us13_n727, us13_n729, us13_n730, us13_n731, us13_n732, us13_n733, 
       us13_n734, us13_n735, us13_n736, us13_n737, us13_n738, us13_n739, us13_n740, us13_n741, us13_n742, 
       us13_n743, us13_n744, us13_n745, us13_n746, us13_n747, us13_n748, us13_n749, us13_n750, us13_n751, 
       us13_n752, us13_n753, us13_n754, us13_n755, us13_n756, us13_n757, us13_n758, us13_n759, us13_n760, 
       us13_n761, us13_n762, us13_n763, us13_n764, us13_n765, us13_n766, us13_n767, us13_n768, us13_n769, 
       us13_n770, us13_n771, us13_n772, us13_n773, us13_n774, us13_n775, us13_n776, us13_n777, us13_n778, 
       us13_n779, us13_n780, us13_n781, us13_n782, us13_n783, us13_n784, us13_n785, us13_n786, us13_n787, 
       us13_n788, us13_n789, us13_n790, us13_n791, us13_n792, us13_n793, us13_n794, us13_n795, us13_n796, 
       us13_n797, us13_n798, us13_n799, us13_n800, us13_n801, us13_n802, us13_n803, us13_n804, us13_n805, 
       us13_n806, us13_n807, us13_n808, us13_n809, us13_n810, us13_n811, us13_n812, us13_n813, us13_n814, 
       us13_n815, us13_n816, us13_n817, us13_n818, us13_n819, us13_n820, us13_n821, us13_n822, us13_n823, 
       us13_n824, us13_n825, us13_n826, us13_n827, us13_n828, us13_n829, us13_n830, us13_n831, us13_n832, 
       us13_n833, us13_n834, us13_n835, us13_n836, us13_n837, us13_n838, us13_n839, us13_n840, us13_n841, 
       us13_n842, us13_n843, us13_n844, us13_n845, us13_n846, us13_n850, us13_n851, us13_n853, us13_n854, 
       us13_n855, us13_n856, us13_n857, us13_n859, us13_n860, us13_n861, us13_n862, us13_n863, us13_n864, 
       us13_n865, us13_n866, us13_n867, us13_n868, us13_n869, us13_n870, us13_n871, us13_n872, us13_n873, 
       us13_n874, us13_n875, us13_n876, us21_n438, us21_n439, us21_n440, us21_n441, us21_n442, us21_n443, 
       us21_n444, us21_n445, us21_n446, us21_n447, us21_n448, us21_n449, us21_n450, us21_n451, us21_n452, 
       us21_n453, us21_n454, us21_n455, us21_n456, us21_n457, us21_n458, us21_n459, us21_n460, us21_n461, 
       us21_n462, us21_n463, us21_n464, us21_n465, us21_n466, us21_n467, us21_n468, us21_n469, us21_n470, 
       us21_n471, us21_n472, us21_n473, us21_n474, us21_n475, us21_n476, us21_n477, us21_n478, us21_n479, 
       us21_n480, us21_n481, us21_n482, us21_n483, us21_n484, us21_n485, us21_n486, us21_n487, us21_n488, 
       us21_n489, us21_n490, us21_n491, us21_n492, us21_n493, us21_n494, us21_n495, us21_n496, us21_n497, 
       us21_n498, us21_n499, us21_n500, us21_n501, us21_n502, us21_n503, us21_n504, us21_n505, us21_n506, 
       us21_n507, us21_n508, us21_n509, us21_n510, us21_n511, us21_n512, us21_n513, us21_n514, us21_n515, 
       us21_n516, us21_n517, us21_n518, us21_n519, us21_n520, us21_n521, us21_n522, us21_n523, us21_n524, 
       us21_n525, us21_n526, us21_n527, us21_n528, us21_n529, us21_n530, us21_n531, us21_n532, us21_n533, 
       us21_n534, us21_n535, us21_n536, us21_n537, us21_n538, us21_n539, us21_n540, us21_n541, us21_n542, 
       us21_n543, us21_n544, us21_n545, us21_n546, us21_n547, us21_n548, us21_n549, us21_n550, us21_n551, 
       us21_n552, us21_n553, us21_n554, us21_n555, us21_n556, us21_n557, us21_n558, us21_n559, us21_n560, 
       us21_n561, us21_n562, us21_n563, us21_n564, us21_n565, us21_n566, us21_n567, us21_n568, us21_n569, 
       us21_n570, us21_n571, us21_n572, us21_n573, us21_n574, us21_n575, us21_n576, us21_n577, us21_n578, 
       us21_n579, us21_n580, us21_n581, us21_n582, us21_n583, us21_n584, us21_n585, us21_n586, us21_n587, 
       us21_n588, us21_n589, us21_n590, us21_n591, us21_n592, us21_n593, us21_n594, us21_n595, us21_n596, 
       us21_n597, us21_n598, us21_n599, us21_n600, us21_n601, us21_n602, us21_n603, us21_n604, us21_n605, 
       us21_n606, us21_n607, us21_n608, us21_n609, us21_n610, us21_n611, us21_n612, us21_n613, us21_n614, 
       us21_n615, us21_n616, us21_n617, us21_n618, us21_n619, us21_n620, us21_n621, us21_n622, us21_n623, 
       us21_n624, us21_n625, us21_n626, us21_n627, us21_n628, us21_n629, us21_n630, us21_n631, us21_n632, 
       us21_n633, us21_n634, us21_n635, us21_n636, us21_n637, us21_n638, us21_n639, us21_n640, us21_n641, 
       us21_n642, us21_n643, us21_n644, us21_n645, us21_n646, us21_n647, us21_n648, us21_n649, us21_n650, 
       us21_n651, us21_n652, us21_n653, us21_n654, us21_n655, us21_n656, us21_n657, us21_n658, us21_n659, 
       us21_n660, us21_n661, us21_n662, us21_n663, us21_n664, us21_n665, us21_n666, us21_n667, us21_n668, 
       us21_n669, us21_n670, us21_n671, us21_n672, us21_n673, us21_n674, us21_n675, us21_n676, us21_n677, 
       us21_n678, us21_n679, us21_n680, us21_n681, us21_n682, us21_n683, us21_n684, us21_n685, us21_n686, 
       us21_n687, us21_n688, us21_n689, us21_n690, us21_n691, us21_n692, us21_n693, us21_n694, us21_n695, 
       us21_n696, us21_n697, us21_n698, us21_n699, us21_n700, us21_n701, us21_n702, us21_n703, us21_n704, 
       us21_n705, us21_n706, us21_n707, us21_n708, us21_n709, us21_n710, us21_n711, us21_n712, us21_n713, 
       us21_n714, us21_n715, us21_n716, us21_n717, us21_n718, us21_n719, us21_n720, us21_n721, us21_n722, 
       us21_n723, us21_n724, us21_n725, us21_n726, us21_n727, us21_n728, us21_n729, us21_n730, us21_n731, 
       us21_n732, us21_n733, us21_n734, us21_n735, us21_n736, us21_n737, us21_n738, us21_n739, us21_n740, 
       us21_n741, us21_n742, us21_n743, us21_n744, us21_n745, us21_n746, us21_n747, us21_n748, us21_n749, 
       us21_n750, us21_n751, us21_n752, us21_n753, us21_n754, us21_n755, us21_n756, us21_n757, us21_n758, 
       us21_n759, us21_n760, us21_n761, us21_n762, us21_n763, us21_n764, us21_n765, us21_n766, us21_n767, 
       us21_n768, us21_n769, us21_n770, us21_n771, us21_n772, us21_n773, us21_n774, us21_n775, us21_n776, 
       us21_n777, us21_n778, us21_n779, us21_n780, us21_n781, us21_n782, us21_n783, us21_n784, us21_n785, 
       us21_n786, us21_n787, us21_n788, us21_n789, us21_n790, us21_n791, us21_n792, us21_n793, us21_n794, 
       us21_n795, us21_n796, us21_n797, us21_n798, us21_n799, us21_n800, us21_n801, us21_n802, us21_n803, 
       us21_n804, us21_n805, us21_n806, us21_n807, us21_n808, us21_n809, us21_n810, us21_n811, us21_n812, 
       us21_n813, us21_n814, us21_n815, us21_n816, us21_n817, us21_n818, us21_n819, us21_n820, us21_n821, 
       us21_n822, us21_n823, us21_n824, us21_n825, us21_n826, us21_n827, us21_n828, us21_n829, us21_n830, 
       us21_n831, us21_n832, us21_n833, us21_n834, us21_n835, us21_n836, us21_n837, us21_n838, us21_n839, 
       us21_n840, us21_n841, us21_n842, us21_n843, us21_n844, us21_n845, us21_n846, us21_n847, us21_n848, 
       us21_n849, us21_n850, us21_n851, us21_n852, us21_n853, us21_n854, us21_n855, us21_n856, us21_n857, 
       us21_n858, us21_n859, us21_n860, us21_n861, us21_n862, us21_n863, us21_n864, us21_n865, us21_n866, 
       us21_n867, us21_n868, us21_n869, us21_n870, us21_n871, us21_n872, us21_n873, us21_n874, us22_n438, 
       us22_n439, us22_n440, us22_n441, us22_n442, us22_n443, us22_n444, us22_n445, us22_n446, us22_n447, 
       us22_n448, us22_n449, us22_n450, us22_n451, us22_n452, us22_n453, us22_n454, us22_n455, us22_n456, 
       us22_n457, us22_n458, us22_n459, us22_n460, us22_n461, us22_n462, us22_n463, us22_n464, us22_n465, 
       us22_n466, us22_n467, us22_n468, us22_n469, us22_n470, us22_n471, us22_n472, us22_n473, us22_n474, 
       us22_n475, us22_n476, us22_n477, us22_n478, us22_n479, us22_n480, us22_n481, us22_n482, us22_n483, 
       us22_n484, us22_n485, us22_n486, us22_n487, us22_n488, us22_n489, us22_n490, us22_n491, us22_n492, 
       us22_n493, us22_n494, us22_n495, us22_n496, us22_n497, us22_n498, us22_n499, us22_n500, us22_n501, 
       us22_n502, us22_n503, us22_n504, us22_n505, us22_n506, us22_n507, us22_n508, us22_n509, us22_n510, 
       us22_n511, us22_n512, us22_n513, us22_n514, us22_n515, us22_n516, us22_n517, us22_n518, us22_n519, 
       us22_n520, us22_n521, us22_n522, us22_n523, us22_n524, us22_n525, us22_n526, us22_n527, us22_n528, 
       us22_n529, us22_n530, us22_n531, us22_n532, us22_n533, us22_n534, us22_n535, us22_n536, us22_n537, 
       us22_n538, us22_n539, us22_n540, us22_n541, us22_n542, us22_n543, us22_n544, us22_n545, us22_n546, 
       us22_n547, us22_n548, us22_n549, us22_n550, us22_n551, us22_n552, us22_n553, us22_n554, us22_n555, 
       us22_n556, us22_n557, us22_n558, us22_n559, us22_n560, us22_n561, us22_n562, us22_n563, us22_n564, 
       us22_n565, us22_n566, us22_n567, us22_n568, us22_n569, us22_n570, us22_n571, us22_n572, us22_n573, 
       us22_n574, us22_n575, us22_n576, us22_n577, us22_n578, us22_n579, us22_n580, us22_n581, us22_n582, 
       us22_n583, us22_n584, us22_n585, us22_n586, us22_n587, us22_n588, us22_n589, us22_n590, us22_n591, 
       us22_n592, us22_n593, us22_n594, us22_n595, us22_n596, us22_n597, us22_n598, us22_n599, us22_n600, 
       us22_n601, us22_n602, us22_n603, us22_n604, us22_n605, us22_n606, us22_n607, us22_n608, us22_n609, 
       us22_n610, us22_n611, us22_n612, us22_n613, us22_n614, us22_n615, us22_n616, us22_n617, us22_n618, 
       us22_n619, us22_n620, us22_n621, us22_n622, us22_n623, us22_n624, us22_n625, us22_n626, us22_n627, 
       us22_n628, us22_n629, us22_n630, us22_n631, us22_n632, us22_n633, us22_n634, us22_n635, us22_n636, 
       us22_n637, us22_n638, us22_n639, us22_n640, us22_n641, us22_n642, us22_n643, us22_n644, us22_n645, 
       us22_n646, us22_n647, us22_n648, us22_n649, us22_n650, us22_n651, us22_n652, us22_n653, us22_n654, 
       us22_n655, us22_n656, us22_n657, us22_n658, us22_n659, us22_n660, us22_n661, us22_n662, us22_n663, 
       us22_n664, us22_n665, us22_n666, us22_n667, us22_n668, us22_n669, us22_n670, us22_n671, us22_n672, 
       us22_n673, us22_n674, us22_n675, us22_n676, us22_n677, us22_n678, us22_n679, us22_n680, us22_n681, 
       us22_n682, us22_n683, us22_n684, us22_n685, us22_n686, us22_n687, us22_n688, us22_n689, us22_n690, 
       us22_n691, us22_n692, us22_n693, us22_n694, us22_n695, us22_n696, us22_n697, us22_n698, us22_n699, 
       us22_n700, us22_n701, us22_n702, us22_n703, us22_n704, us22_n705, us22_n706, us22_n707, us22_n708, 
       us22_n709, us22_n710, us22_n711, us22_n712, us22_n713, us22_n714, us22_n715, us22_n716, us22_n717, 
       us22_n718, us22_n719, us22_n720, us22_n721, us22_n722, us22_n723, us22_n724, us22_n725, us22_n726, 
       us22_n727, us22_n728, us22_n729, us22_n730, us22_n731, us22_n732, us22_n733, us22_n734, us22_n735, 
       us22_n736, us22_n737, us22_n738, us22_n739, us22_n740, us22_n741, us22_n742, us22_n743, us22_n744, 
       us22_n745, us22_n746, us22_n747, us22_n748, us22_n749, us22_n750, us22_n751, us22_n752, us22_n753, 
       us22_n754, us22_n755, us22_n756, us22_n757, us22_n758, us22_n759, us22_n760, us22_n761, us22_n762, 
       us22_n763, us22_n764, us22_n765, us22_n766, us22_n767, us22_n768, us22_n769, us22_n770, us22_n771, 
       us22_n772, us22_n773, us22_n774, us22_n775, us22_n776, us22_n777, us22_n778, us22_n779, us22_n780, 
       us22_n781, us22_n782, us22_n783, us22_n784, us22_n785, us22_n786, us22_n787, us22_n788, us22_n789, 
       us22_n790, us22_n791, us22_n792, us22_n793, us22_n794, us22_n795, us22_n796, us22_n797, us22_n798, 
       us22_n799, us22_n800, us22_n801, us22_n802, us22_n803, us22_n804, us22_n805, us22_n806, us22_n807, 
       us22_n808, us22_n809, us22_n810, us22_n811, us22_n812, us22_n813, us22_n814, us22_n815, us22_n816, 
       us22_n817, us22_n818, us22_n819, us22_n820, us22_n821, us22_n822, us22_n823, us22_n824, us22_n825, 
       us22_n826, us22_n827, us22_n828, us22_n829, us22_n830, us22_n831, us22_n832, us22_n833, us22_n834, 
       us22_n835, us22_n836, us22_n837, us22_n838, us22_n839, us22_n840, us22_n841, us22_n842, us22_n843, 
       us22_n844, us22_n845, us22_n846, us22_n847, us22_n848, us22_n849, us22_n850, us22_n851, us22_n852, 
       us22_n853, us22_n854, us22_n855, us22_n856, us22_n857, us22_n858, us22_n859, us22_n860, us22_n861, 
       us22_n862, us22_n863, us22_n864, us22_n865, us22_n866, us22_n867, us22_n868, us22_n869, us22_n870, 
       us22_n871, us22_n872, us22_n873, us22_n874, us32_n438, us32_n439, us32_n440, us32_n441, us32_n442, 
       us32_n443, us32_n444, us32_n445, us32_n446, us32_n447, us32_n448, us32_n449, us32_n450, us32_n451, 
       us32_n452, us32_n453, us32_n454, us32_n455, us32_n456, us32_n457, us32_n458, us32_n459, us32_n460, 
       us32_n461, us32_n462, us32_n463, us32_n464, us32_n465, us32_n466, us32_n467, us32_n468, us32_n469, 
       us32_n470, us32_n471, us32_n472, us32_n473, us32_n474, us32_n475, us32_n476, us32_n477, us32_n478, 
       us32_n479, us32_n480, us32_n481, us32_n482, us32_n483, us32_n484, us32_n485, us32_n486, us32_n487, 
       us32_n488, us32_n489, us32_n490, us32_n491, us32_n492, us32_n493, us32_n494, us32_n495, us32_n496, 
       us32_n497, us32_n498, us32_n499, us32_n500, us32_n501, us32_n502, us32_n503, us32_n504, us32_n505, 
       us32_n506, us32_n507, us32_n508, us32_n509, us32_n510, us32_n511, us32_n512, us32_n513, us32_n514, 
       us32_n515, us32_n516, us32_n517, us32_n518, us32_n519, us32_n520, us32_n521, us32_n522, us32_n523, 
       us32_n524, us32_n525, us32_n526, us32_n527, us32_n528, us32_n529, us32_n530, us32_n531, us32_n532, 
       us32_n533, us32_n534, us32_n535, us32_n536, us32_n537, us32_n538, us32_n539, us32_n540, us32_n541, 
       us32_n542, us32_n543, us32_n544, us32_n545, us32_n546, us32_n547, us32_n548, us32_n549, us32_n550, 
       us32_n551, us32_n552, us32_n553, us32_n554, us32_n555, us32_n556, us32_n557, us32_n558, us32_n559, 
       us32_n560, us32_n561, us32_n562, us32_n563, us32_n564, us32_n565, us32_n566, us32_n567, us32_n568, 
       us32_n569, us32_n570, us32_n571, us32_n572, us32_n573, us32_n574, us32_n575, us32_n576, us32_n577, 
       us32_n578, us32_n579, us32_n580, us32_n581, us32_n582, us32_n583, us32_n584, us32_n585, us32_n586, 
       us32_n587, us32_n588, us32_n589, us32_n590, us32_n591, us32_n592, us32_n593, us32_n594, us32_n595, 
       us32_n596, us32_n597, us32_n598, us32_n599, us32_n600, us32_n601, us32_n602, us32_n603, us32_n604, 
       us32_n605, us32_n606, us32_n607, us32_n608, us32_n609, us32_n610, us32_n611, us32_n612, us32_n613, 
       us32_n614, us32_n615, us32_n616, us32_n617, us32_n618, us32_n619, us32_n620, us32_n621, us32_n622, 
       us32_n623, us32_n624, us32_n625, us32_n626, us32_n627, us32_n628, us32_n629, us32_n630, us32_n631, 
       us32_n632, us32_n633, us32_n634, us32_n635, us32_n636, us32_n637, us32_n638, us32_n639, us32_n640, 
       us32_n641, us32_n642, us32_n643, us32_n644, us32_n645, us32_n646, us32_n647, us32_n648, us32_n649, 
       us32_n650, us32_n651, us32_n652, us32_n653, us32_n654, us32_n655, us32_n656, us32_n657, us32_n658, 
       us32_n659, us32_n660, us32_n661, us32_n662, us32_n663, us32_n664, us32_n665, us32_n666, us32_n667, 
       us32_n668, us32_n669, us32_n670, us32_n671, us32_n672, us32_n673, us32_n674, us32_n675, us32_n676, 
       us32_n677, us32_n678, us32_n679, us32_n680, us32_n681, us32_n682, us32_n683, us32_n684, us32_n685, 
       us32_n686, us32_n687, us32_n688, us32_n689, us32_n690, us32_n691, us32_n692, us32_n693, us32_n694, 
       us32_n695, us32_n696, us32_n697, us32_n698, us32_n699, us32_n700, us32_n701, us32_n702, us32_n703, 
       us32_n704, us32_n705, us32_n706, us32_n707, us32_n708, us32_n709, us32_n710, us32_n711, us32_n712, 
       us32_n713, us32_n714, us32_n715, us32_n716, us32_n717, us32_n718, us32_n719, us32_n720, us32_n721, 
       us32_n722, us32_n723, us32_n724, us32_n725, us32_n726, us32_n727, us32_n728, us32_n729, us32_n730, 
       us32_n731, us32_n732, us32_n733, us32_n734, us32_n735, us32_n736, us32_n737, us32_n738, us32_n739, 
       us32_n740, us32_n741, us32_n742, us32_n743, us32_n744, us32_n745, us32_n746, us32_n747, us32_n748, 
       us32_n749, us32_n750, us32_n751, us32_n752, us32_n753, us32_n754, us32_n755, us32_n756, us32_n757, 
       us32_n758, us32_n759, us32_n760, us32_n761, us32_n762, us32_n763, us32_n764, us32_n765, us32_n766, 
       us32_n767, us32_n768, us32_n769, us32_n770, us32_n771, us32_n772, us32_n773, us32_n774, us32_n775, 
       us32_n776, us32_n777, us32_n778, us32_n779, us32_n780, us32_n781, us32_n782, us32_n783, us32_n784, 
       us32_n785, us32_n786, us32_n787, us32_n788, us32_n789, us32_n790, us32_n791, us32_n792, us32_n793, 
       us32_n794, us32_n795, us32_n796, us32_n797, us32_n798, us32_n799, us32_n800, us32_n801, us32_n802, 
       us32_n803, us32_n804, us32_n805, us32_n806, us32_n807, us32_n808, us32_n809, us32_n810, us32_n811, 
       us32_n812, us32_n813, us32_n814, us32_n815, us32_n816, us32_n817, us32_n818, us32_n819, us32_n820, 
       us32_n821, us32_n822, us32_n823, us32_n824, us32_n825, us32_n826, us32_n827, us32_n828, us32_n829, 
       us32_n830, us32_n831, us32_n832, us32_n833, us32_n834, us32_n835, us32_n836, us32_n837, us32_n838, 
       us32_n839, us32_n840, us32_n841, us32_n842, us32_n843, us32_n844, us32_n845, us32_n846, us32_n847, 
       us32_n848, us32_n849, us32_n850, us32_n851, us32_n852, us32_n853, us32_n854, us32_n855, us32_n856, 
       us32_n857, us32_n858, us32_n859, us32_n860, us32_n861, us32_n862, us32_n863, us32_n864, us32_n865, 
       us32_n866, us32_n867, us32_n868, us32_n869, us32_n870, us32_n871, us32_n872, us32_n873, us32_n874, 
       us32_n875,  us32_n876;
  NOR2_X1 us00_U10 (.A2( us00_n132 ) , .A1( us00_n255 ) , .ZN( us00_n302 ) );
  NOR4_X1 us00_U100 (.A2( us00_n193 ) , .ZN( us00_n340 ) , .A3( us00_n347 ) , .A4( us00_n348 ) , .A1( us00_n83 ) );
  NAND4_X1 us00_U101 (.ZN( us00_n183 ) , .A1( us00_n395 ) , .A2( us00_n396 ) , .A3( us00_n397 ) , .A4( us00_n398 ) );
  NOR3_X1 us00_U102 (.A1( us00_n267 ) , .A3( us00_n276 ) , .A2( us00_n369 ) , .ZN( us00_n397 ) );
  AOI211_X1 us00_U103 (.C1( us00_n16 ) , .ZN( us00_n395 ) , .A( us00_n399 ) , .B( us00_n400 ) , .C2( us00_n44 ) );
  NOR4_X1 us00_U104 (.A1( us00_n160 ) , .A2( us00_n310 ) , .A4( us00_n332 ) , .A3( us00_n345 ) , .ZN( us00_n396 ) );
  NAND4_X1 us00_U105 (.ZN( us00_n132 ) , .A1( us00_n326 ) , .A2( us00_n327 ) , .A3( us00_n328 ) , .A4( us00_n329 ) );
  NOR3_X1 us00_U106 (.A3( us00_n106 ) , .A1( us00_n210 ) , .A2( us00_n226 ) , .ZN( us00_n328 ) );
  AOI211_X1 us00_U107 (.C1( us00_n26 ) , .ZN( us00_n326 ) , .A( us00_n337 ) , .B( us00_n338 ) , .C2( us00_n38 ) );
  NOR4_X1 us00_U108 (.ZN( us00_n329 ) , .A1( us00_n330 ) , .A2( us00_n331 ) , .A3( us00_n332 ) , .A4( us00_n333 ) );
  NOR2_X1 us00_U109 (.ZN( us00_n191 ) , .A2( us00_n45 ) , .A1( us00_n46 ) );
  NOR2_X1 us00_U11 (.ZN( us00_n184 ) , .A1( us00_n199 ) , .A2( us00_n70 ) );
  NOR4_X1 us00_U110 (.A2( us00_n111 ) , .A4( us00_n195 ) , .A3( us00_n211 ) , .A1( us00_n221 ) , .ZN( us00_n257 ) );
  NOR4_X1 us00_U111 (.ZN( us00_n258 ) , .A1( us00_n265 ) , .A2( us00_n266 ) , .A3( us00_n267 ) , .A4( us00_n268 ) );
  NOR4_X1 us00_U112 (.ZN( us00_n259 ) , .A1( us00_n260 ) , .A2( us00_n261 ) , .A3( us00_n262 ) , .A4( us00_n263 ) );
  NAND4_X1 us00_U113 (.A1( us00_n389 ) , .A2( us00_n390 ) , .A3( us00_n391 ) , .A4( us00_n392 ) , .ZN( us00_n99 ) );
  NOR4_X1 us00_U114 (.A3( us00_n275 ) , .A2( us00_n296 ) , .A1( us00_n311 ) , .ZN( us00_n390 ) , .A4( us00_n393 ) );
  NOR4_X1 us00_U115 (.A3( us00_n266 ) , .A4( us00_n331 ) , .A2( us00_n358 ) , .A1( us00_n370 ) , .ZN( us00_n391 ) );
  NOR4_X1 us00_U116 (.A4( us00_n159 ) , .A3( us00_n246 ) , .A1( us00_n319 ) , .A2( us00_n344 ) , .ZN( us00_n392 ) );
  NAND4_X1 us00_U117 (.ZN( us00_n101 ) , .A1( us00_n184 ) , .A3( us00_n185 ) , .A4( us00_n186 ) , .A2( us00_n5 ) );
  AOI221_X1 us00_U118 (.B1( us00_n12 ) , .C2( us00_n15 ) , .ZN( us00_n185 ) , .A( us00_n196 ) , .C1( us00_n35 ) , .B2( us00_n37 ) );
  INV_X1 us00_U119 (.A( us00_n198 ) , .ZN( us00_n5 ) );
  INV_X1 us00_U12 (.A( us00_n197 ) , .ZN( us00_n37 ) );
  NOR4_X1 us00_U120 (.ZN( us00_n186 ) , .A1( us00_n187 ) , .A2( us00_n188 ) , .A3( us00_n189 ) , .A4( us00_n190 ) );
  NAND4_X1 us00_U121 (.ZN( us00_n136 ) , .A2( us00_n156 ) , .A3( us00_n157 ) , .A4( us00_n158 ) , .A1( us00_n20 ) );
  INV_X1 us00_U122 (.A( us00_n168 ) , .ZN( us00_n20 ) );
  AOI221_X1 us00_U123 (.B1( us00_n15 ) , .ZN( us00_n156 ) , .C1( us00_n16 ) , .A( us00_n167 ) , .B2( us00_n32 ) , .C2( us00_n33 ) );
  NOR4_X1 us00_U124 (.ZN( us00_n158 ) , .A1( us00_n159 ) , .A2( us00_n160 ) , .A3( us00_n161 ) , .A4( us00_n162 ) );
  NAND4_X1 us00_U125 (.ZN( us00_n199 ) , .A1( us00_n401 ) , .A2( us00_n402 ) , .A3( us00_n403 ) , .A4( us00_n404 ) );
  NOR4_X1 us00_U126 (.A2( us00_n122 ) , .A1( us00_n142 ) , .A3( us00_n321 ) , .ZN( us00_n401 ) , .A4( us00_n407 ) );
  NOR4_X1 us00_U127 (.A2( us00_n235 ) , .A4( us00_n277 ) , .A3( us00_n309 ) , .A1( us00_n346 ) , .ZN( us00_n402 ) );
  NOR4_X1 us00_U128 (.A4( us00_n161 ) , .A2( us00_n294 ) , .A3( us00_n333 ) , .A1( us00_n371 ) , .ZN( us00_n403 ) );
  NOR2_X1 us00_U129 (.ZN( us00_n144 ) , .A1( us00_n32 ) , .A2( us00_n45 ) );
  NOR4_X1 us00_U13 (.ZN( us00_n171 ) , .A1( us00_n336 ) , .A2( us00_n361 ) , .A3( us00_n431 ) , .A4( us00_n432 ) );
  NOR2_X1 us00_U130 (.A2( us00_n15 ) , .ZN( us00_n88 ) , .A1( us00_n9 ) );
  NOR2_X1 us00_U131 (.A1( us00_n23 ) , .ZN( us00_n230 ) , .A2( us00_n9 ) );
  NAND4_X1 us00_U132 (.ZN( us00_n154 ) , .A2( us00_n3 ) , .A1( us00_n302 ) , .A3( us00_n303 ) , .A4( us00_n304 ) );
  NOR4_X1 us00_U133 (.ZN( us00_n304 ) , .A1( us00_n305 ) , .A2( us00_n306 ) , .A3( us00_n307 ) , .A4( us00_n308 ) );
  AOI221_X1 us00_U134 (.C1( us00_n24 ) , .B1( us00_n25 ) , .ZN( us00_n303 ) , .C2( us00_n312 ) , .A( us00_n313 ) , .B2( us00_n32 ) );
  INV_X1 us00_U135 (.A( us00_n270 ) , .ZN( us00_n3 ) );
  NAND4_X1 us00_U136 (.A2( us00_n10 ) , .A1( us00_n382 ) , .A3( us00_n383 ) , .A4( us00_n384 ) , .ZN( us00_n75 ) );
  AOI221_X1 us00_U137 (.B1( us00_n17 ) , .C1( us00_n26 ) , .C2( us00_n36 ) , .ZN( us00_n383 ) , .A( us00_n388 ) , .B2( us00_n41 ) );
  INV_X1 us00_U138 (.ZN( us00_n10 ) , .A( us00_n99 ) );
  NOR2_X1 us00_U139 (.A2( us00_n183 ) , .A1( us00_n199 ) , .ZN( us00_n382 ) );
  OR3_X1 us00_U14 (.A2( us00_n2 ) , .A3( us00_n300 ) , .A1( us00_n349 ) , .ZN( us00_n431 ) );
  INV_X1 us00_U140 (.A( us00_n115 ) , .ZN( us00_n47 ) );
  INV_X1 us00_U141 (.ZN( us00_n13 ) , .A( us00_n414 ) );
  OAI21_X1 us00_U142 (.B2( us00_n26 ) , .ZN( us00_n414 ) , .A( us00_n43 ) , .B1( us00_n68 ) );
  OR4_X1 us00_U143 (.A1( us00_n212 ) , .ZN( us00_n305 ) , .A2( us00_n309 ) , .A3( us00_n310 ) , .A4( us00_n311 ) );
  OR4_X1 us00_U144 (.ZN( us00_n355 ) , .A1( us00_n357 ) , .A2( us00_n358 ) , .A4( us00_n359 ) , .A3( us00_n56 ) );
  OR4_X1 us00_U145 (.A1( us00_n165 ) , .A2( us00_n299 ) , .A3( us00_n348 ) , .A4( us00_n359 ) , .ZN( us00_n411 ) );
  OR4_X1 us00_U146 (.ZN( us00_n187 ) , .A1( us00_n192 ) , .A2( us00_n193 ) , .A3( us00_n194 ) , .A4( us00_n195 ) );
  OR4_X1 us00_U147 (.ZN( us00_n293 ) , .A1( us00_n294 ) , .A2( us00_n295 ) , .A3( us00_n296 ) , .A4( us00_n297 ) );
  NAND2_X1 us00_U148 (.ZN( us00_n264 ) , .A1( us00_n4 ) , .A2( us00_n40 ) );
  OR3_X1 us00_U149 (.ZN( us00_n366 ) , .A1( us00_n369 ) , .A2( us00_n370 ) , .A3( us00_n371 ) );
  OR4_X1 us00_U15 (.A3( us00_n324 ) , .ZN( us00_n432 ) , .A1( us00_n433 ) , .A2( us00_n434 ) , .A4( us00_n435 ) );
  AOI221_X1 us00_U150 (.C2( us00_n14 ) , .ZN( us00_n157 ) , .B2( us00_n163 ) , .A( us00_n164 ) , .B1( us00_n38 ) , .C1( us00_n45 ) );
  OR2_X1 us00_U151 (.ZN( us00_n164 ) , .A1( us00_n165 ) , .A2( us00_n166 ) );
  INV_X1 us00_U152 (.A( us00_n123 ) , .ZN( us00_n8 ) );
  OAI21_X1 us00_U153 (.ZN( us00_n123 ) , .B1( us00_n124 ) , .A( us00_n32 ) , .B2( us00_n9 ) );
  INV_X1 us00_U154 (.ZN( us00_n18 ) , .A( us00_n205 ) );
  AOI21_X1 us00_U155 (.ZN( us00_n205 ) , .B1( us00_n206 ) , .A( us00_n207 ) , .B2( us00_n21 ) );
  NAND2_X1 us00_U156 (.ZN( us00_n128 ) , .A2( us00_n412 ) , .A1( us00_n430 ) );
  OAI222_X1 us00_U157 (.ZN( us00_n120 ) , .A2( us00_n128 ) , .B1( us00_n129 ) , .B2( us00_n130 ) , .A1( us00_n60 ) , .C1( us00_n63 ) , .C2( us00_n72 ) );
  OAI222_X1 us00_U158 (.A2( us00_n129 ) , .B1( us00_n130 ) , .B2( us00_n230 ) , .C2( us00_n252 ) , .ZN( us00_n372 ) , .A1( us00_n71 ) , .C1( us00_n72 ) );
  OAI222_X1 us00_U159 (.B1( us00_n130 ) , .C2( us00_n153 ) , .ZN( us00_n168 ) , .B2( us00_n169 ) , .A2( us00_n62 ) , .C1( us00_n63 ) , .A1( us00_n71 ) );
  INV_X1 us00_U16 (.ZN( us00_n2 ) , .A( us00_n264 ) );
  OAI222_X1 us00_U160 (.C2( us00_n130 ) , .C1( us00_n153 ) , .B1( us00_n180 ) , .ZN( us00_n260 ) , .A1( us00_n61 ) , .A2( us00_n85 ) , .B2( us00_n91 ) );
  NOR4_X1 us00_U161 (.A4( us00_n265 ) , .A3( us00_n297 ) , .ZN( us00_n384 ) , .A1( us00_n385 ) , .A2( us00_n386 ) );
  OR4_X1 us00_U162 (.A3( us00_n245 ) , .A1( us00_n318 ) , .A2( us00_n330 ) , .A4( us00_n343 ) , .ZN( us00_n385 ) );
  OAI22_X1 us00_U163 (.A2( us00_n114 ) , .A1( us00_n191 ) , .ZN( us00_n386 ) , .B1( us00_n387 ) , .B2( us00_n60 ) );
  NOR3_X1 us00_U164 (.A3( us00_n14 ) , .A2( us00_n27 ) , .ZN( us00_n387 ) , .A1( us00_n95 ) );
  AOI22_X1 us00_U165 (.A2( us00_n12 ) , .ZN( us00_n181 ) , .B2( us00_n34 ) , .A1( us00_n47 ) , .B1( us00_n9 ) );
  INV_X1 us00_U166 (.A( us00_n147 ) , .ZN( us00_n38 ) );
  AOI221_X1 us00_U167 (.B2( us00_n15 ) , .C1( us00_n25 ) , .C2( us00_n33 ) , .ZN( us00_n389 ) , .A( us00_n394 ) , .B1( us00_n46 ) );
  OAI22_X1 us00_U168 (.A1( us00_n169 ) , .ZN( us00_n394 ) , .B1( us00_n65 ) , .A2( us00_n71 ) , .B2( us00_n92 ) );
  INV_X1 us00_U169 (.ZN( us00_n45 ) , .A( us00_n87 ) );
  INV_X1 us00_U17 (.A( us00_n128 ) , .ZN( us00_n14 ) );
  NAND2_X1 us00_U170 (.ZN( us00_n115 ) , .A2( us00_n424 ) , .A1( us00_n426 ) );
  OAI22_X1 us00_U171 (.A2( us00_n115 ) , .B2( us00_n149 ) , .A1( us00_n178 ) , .ZN( us00_n240 ) , .B1( us00_n61 ) );
  OAI221_X1 us00_U172 (.ZN( us00_n140 ) , .B1( us00_n147 ) , .B2( us00_n148 ) , .C2( us00_n149 ) , .A( us00_n150 ) , .C1( us00_n60 ) );
  AOI22_X1 us00_U173 (.B2( us00_n11 ) , .A1( us00_n14 ) , .ZN( us00_n150 ) , .A2( us00_n39 ) , .B1( us00_n45 ) );
  INV_X1 us00_U174 (.ZN( us00_n15 ) , .A( us00_n91 ) );
  OAI22_X1 us00_U175 (.A1( us00_n133 ) , .B2( us00_n148 ) , .A2( us00_n149 ) , .ZN( us00_n167 ) , .B1( us00_n64 ) );
  INV_X1 us00_U176 (.ZN( us00_n46 ) , .A( us00_n61 ) );
  OAI22_X1 us00_U177 (.B1( us00_n147 ) , .B2( us00_n149 ) , .A1( us00_n153 ) , .ZN( us00_n388 ) , .A2( us00_n98 ) );
  OAI22_X1 us00_U178 (.B2( us00_n130 ) , .B1( us00_n208 ) , .ZN( us00_n253 ) , .A2( us00_n61 ) , .A1( us00_n62 ) );
  INV_X1 us00_U179 (.A( us00_n133 ) , .ZN( us00_n40 ) );
  AOI222_X1 us00_U18 (.B1( us00_n124 ) , .C1( us00_n14 ) , .A2( us00_n15 ) , .B2( us00_n206 ) , .ZN( us00_n272 ) , .A1( us00_n44 ) , .C2( us00_n46 ) );
  OAI22_X1 us00_U180 (.B2( us00_n127 ) , .ZN( us00_n151 ) , .A1( us00_n153 ) , .A2( us00_n61 ) , .B1( us00_n65 ) );
  OAI22_X1 us00_U181 (.A1( us00_n62 ) , .A2( us00_n63 ) , .ZN( us00_n96 ) , .B1( us00_n97 ) , .B2( us00_n98 ) );
  INV_X1 us00_U182 (.ZN( us00_n32 ) , .A( us00_n89 ) );
  INV_X1 us00_U183 (.ZN( us00_n17 ) , .A( us00_n72 ) );
  INV_X1 us00_U184 (.ZN( us00_n44 ) , .A( us00_n63 ) );
  OAI22_X1 us00_U185 (.A2( us00_n115 ) , .ZN( us00_n131 ) , .B2( us00_n133 ) , .A1( us00_n85 ) , .B1( us00_n97 ) );
  OAI22_X1 us00_U186 (.ZN( us00_n69 ) , .A1( us00_n71 ) , .A2( us00_n72 ) , .B1( us00_n73 ) , .B2( us00_n74 ) );
  INV_X1 us00_U187 (.ZN( us00_n12 ) , .A( us00_n208 ) );
  OAI22_X1 us00_U188 (.A2( us00_n133 ) , .ZN( us00_n381 ) , .B2( us00_n71 ) , .B1( us00_n86 ) , .A1( us00_n97 ) );
  INV_X1 us00_U189 (.A( us00_n127 ) , .ZN( us00_n35 ) );
  AOI222_X1 us00_U19 (.B2( us00_n14 ) , .A1( us00_n23 ) , .ZN( us00_n314 ) , .A2( us00_n34 ) , .C1( us00_n36 ) , .C2( us00_n4 ) , .B1( us00_n47 ) );
  OAI22_X1 us00_U190 (.B2( us00_n128 ) , .B1( us00_n147 ) , .ZN( us00_n287 ) , .A1( us00_n74 ) , .A2( us00_n91 ) );
  OAI22_X1 us00_U191 (.A2( us00_n147 ) , .ZN( us00_n182 ) , .B2( us00_n60 ) , .B1( us00_n86 ) , .A1( us00_n97 ) );
  INV_X1 us00_U192 (.ZN( us00_n34 ) , .A( us00_n74 ) );
  NOR2_X1 us00_U193 (.ZN( us00_n162 ) , .A2( us00_n60 ) , .A1( us00_n72 ) );
  NOR2_X1 us00_U194 (.ZN( us00_n107 ) , .A1( us00_n180 ) , .A2( us00_n62 ) );
  NOR2_X1 us00_U195 (.A1( us00_n149 ) , .ZN( us00_n211 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U196 (.A1( us00_n149 ) , .A2( us00_n180 ) , .ZN( us00_n283 ) );
  NOR2_X1 us00_U197 (.A1( us00_n149 ) , .ZN( us00_n307 ) , .A2( us00_n71 ) );
  NOR2_X1 us00_U198 (.ZN( us00_n122 ) , .A2( us00_n133 ) , .A1( us00_n72 ) );
  NOR2_X1 us00_U199 (.A1( us00_n133 ) , .A2( us00_n153 ) , .ZN( us00_n159 ) );
  AOI222_X1 us00_U20 (.C1( us00_n14 ) , .A1( us00_n17 ) , .ZN( us00_n217 ) , .C2( us00_n32 ) , .B1( us00_n36 ) , .A2( us00_n38 ) , .B2( us00_n7 ) );
  NOR2_X1 us00_U200 (.ZN( us00_n142 ) , .A1( us00_n72 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U201 (.ZN( us00_n331 ) , .A1( us00_n63 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U202 (.A2( us00_n178 ) , .ZN( us00_n300 ) , .A1( us00_n63 ) );
  NOR2_X1 us00_U203 (.A1( us00_n149 ) , .ZN( us00_n223 ) , .A2( us00_n64 ) );
  NOR2_X1 us00_U204 (.ZN( us00_n265 ) , .A2( us00_n91 ) , .A1( us00_n98 ) );
  NOR2_X1 us00_U205 (.A1( us00_n127 ) , .A2( us00_n128 ) , .ZN( us00_n345 ) );
  NOR2_X1 us00_U206 (.ZN( us00_n262 ) , .A2( us00_n62 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U207 (.A2( us00_n149 ) , .ZN( us00_n248 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U208 (.ZN( us00_n276 ) , .A1( us00_n74 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U209 (.ZN( us00_n266 ) , .A1( us00_n71 ) , .A2( us00_n97 ) );
  INV_X1 us00_U21 (.A( us00_n230 ) , .ZN( us00_n7 ) );
  INV_X1 us00_U210 (.A( us00_n130 ) , .ZN( us00_n43 ) );
  NOR2_X1 us00_U211 (.ZN( us00_n108 ) , .A2( us00_n133 ) , .A1( us00_n65 ) );
  NOR2_X1 us00_U212 (.A2( us00_n153 ) , .ZN( us00_n349 ) , .A1( us00_n74 ) );
  NOR2_X1 us00_U213 (.ZN( us00_n346 ) , .A1( us00_n61 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U214 (.A2( us00_n208 ) , .ZN( us00_n249 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U215 (.ZN( us00_n278 ) , .A1( us00_n61 ) , .A2( us00_n86 ) );
  INV_X1 us00_U216 (.A( us00_n149 ) , .ZN( us00_n25 ) );
  NOR2_X1 us00_U217 (.A1( us00_n208 ) , .ZN( us00_n225 ) , .A2( us00_n63 ) );
  NOR2_X1 us00_U218 (.A2( us00_n133 ) , .ZN( us00_n204 ) , .A1( us00_n208 ) );
  NOR2_X1 us00_U219 (.A1( us00_n208 ) , .ZN( us00_n275 ) , .A2( us00_n74 ) );
  NOR4_X1 us00_U22 (.A3( us00_n248 ) , .A1( us00_n268 ) , .A4( us00_n283 ) , .A2( us00_n356 ) , .ZN( us00_n404 ) );
  NOR2_X1 us00_U220 (.ZN( us00_n189 ) , .A1( us00_n208 ) , .A2( us00_n61 ) );
  INV_X1 us00_U221 (.ZN( us00_n26 ) , .A( us00_n85 ) );
  NOR2_X1 us00_U222 (.ZN( us00_n106 ) , .A1( us00_n127 ) , .A2( us00_n169 ) );
  NOR2_X1 us00_U223 (.ZN( us00_n111 ) , .A1( us00_n208 ) , .A2( us00_n64 ) );
  NOR2_X1 us00_U224 (.ZN( us00_n109 ) , .A1( us00_n178 ) , .A2( us00_n64 ) );
  NOR2_X1 us00_U225 (.A1( us00_n178 ) , .A2( us00_n180 ) , .ZN( us00_n336 ) );
  NOR2_X1 us00_U226 (.A1( us00_n208 ) , .ZN( us00_n350 ) , .A2( us00_n98 ) );
  NOR2_X1 us00_U227 (.A1( us00_n127 ) , .ZN( us00_n210 ) , .A2( us00_n62 ) );
  NOR2_X1 us00_U228 (.A1( us00_n127 ) , .ZN( us00_n322 ) , .A2( us00_n86 ) );
  NOR2_X1 us00_U229 (.ZN( us00_n369 ) , .A1( us00_n92 ) , .A2( us00_n97 ) );
  NOR4_X1 us00_U23 (.A2( us00_n247 ) , .A3( us00_n295 ) , .A4( us00_n320 ) , .A1( us00_n357 ) , .ZN( us00_n398 ) );
  NOR2_X1 us00_U230 (.A2( us00_n169 ) , .ZN( us00_n334 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U231 (.ZN( us00_n213 ) , .A2( us00_n86 ) , .A1( us00_n92 ) );
  NOR2_X1 us00_U232 (.ZN( us00_n161 ) , .A2( us00_n180 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U233 (.ZN( us00_n370 ) , .A2( us00_n60 ) , .A1( us00_n65 ) );
  NOR2_X1 us00_U234 (.A1( us00_n115 ) , .ZN( us00_n321 ) , .A2( us00_n72 ) );
  INV_X1 us00_U235 (.ZN( us00_n36 ) , .A( us00_n71 ) );
  NOR2_X1 us00_U236 (.A1( us00_n148 ) , .ZN( us00_n216 ) , .A2( us00_n87 ) );
  NOR2_X1 us00_U237 (.A1( us00_n148 ) , .A2( us00_n180 ) , .ZN( us00_n215 ) );
  NOR2_X1 us00_U238 (.ZN( us00_n320 ) , .A2( us00_n63 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U239 (.A1( us00_n128 ) , .ZN( us00_n332 ) , .A2( us00_n63 ) );
  NOR4_X1 us00_U24 (.ZN( us00_n342 ) , .A2( us00_n343 ) , .A3( us00_n344 ) , .A4( us00_n345 ) , .A1( us00_n57 ) );
  NOR2_X1 us00_U240 (.A1( us00_n148 ) , .ZN( us00_n368 ) , .A2( us00_n98 ) );
  NOR2_X1 us00_U241 (.A2( us00_n180 ) , .ZN( us00_n57 ) , .A1( us00_n97 ) );
  OAI22_X1 us00_U242 (.ZN( us00_n121 ) , .A1( us00_n125 ) , .B1( us00_n126 ) , .B2( us00_n127 ) , .A2( us00_n71 ) );
  NOR2_X1 us00_U243 (.ZN( us00_n126 ) , .A1( us00_n17 ) , .A2( us00_n25 ) );
  NOR3_X1 us00_U244 (.A3( us00_n12 ) , .ZN( us00_n125 ) , .A1( us00_n14 ) , .A2( us00_n24 ) );
  NOR2_X1 us00_U245 (.A2( us00_n133 ) , .ZN( us00_n347 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U246 (.ZN( us00_n110 ) , .A1( us00_n128 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U247 (.ZN( us00_n333 ) , .A1( us00_n85 ) , .A2( us00_n92 ) );
  NOR2_X1 us00_U248 (.A1( us00_n148 ) , .ZN( us00_n214 ) , .A2( us00_n92 ) );
  NOR2_X1 us00_U249 (.A1( us00_n153 ) , .ZN( us00_n246 ) , .A2( us00_n64 ) );
  NOR4_X1 us00_U25 (.A4( us00_n262 ) , .A3( us00_n298 ) , .A1( us00_n334 ) , .A2( us00_n360 ) , .ZN( us00_n421 ) );
  NOR2_X1 us00_U250 (.A1( us00_n115 ) , .ZN( us00_n263 ) , .A2( us00_n65 ) );
  OAI22_X1 us00_U251 (.B2( us00_n128 ) , .A1( us00_n133 ) , .A2( us00_n149 ) , .ZN( us00_n433 ) , .B1( us00_n437 ) );
  NOR3_X1 us00_U252 (.A1( us00_n31 ) , .A3( us00_n40 ) , .A2( us00_n41 ) , .ZN( us00_n437 ) );
  NOR2_X1 us00_U253 (.A1( us00_n115 ) , .A2( us00_n149 ) , .ZN( us00_n371 ) );
  NOR2_X1 us00_U254 (.A2( us00_n133 ) , .A1( us00_n169 ) , .ZN( us00_n361 ) );
  NOR2_X1 us00_U255 (.A2( us00_n133 ) , .ZN( us00_n160 ) , .A1( us00_n91 ) );
  NOR2_X1 us00_U256 (.ZN( us00_n323 ) , .A2( us00_n64 ) , .A1( us00_n91 ) );
  NOR2_X1 us00_U257 (.A1( us00_n169 ) , .ZN( us00_n360 ) , .A2( us00_n74 ) );
  NOR2_X1 us00_U258 (.A1( us00_n169 ) , .ZN( us00_n319 ) , .A2( us00_n61 ) );
  NOR2_X1 us00_U259 (.ZN( us00_n207 ) , .A2( us00_n72 ) , .A1( us00_n87 ) );
  NOR4_X1 us00_U26 (.A1( us00_n189 ) , .ZN( us00_n327 ) , .A2( us00_n334 ) , .A3( us00_n335 ) , .A4( us00_n336 ) );
  NOR2_X1 us00_U260 (.ZN( us00_n356 ) , .A2( us00_n65 ) , .A1( us00_n87 ) );
  NOR2_X1 us00_U261 (.A1( us00_n130 ) , .ZN( us00_n247 ) , .A2( us00_n62 ) );
  AOI21_X1 us00_U262 (.B2( us00_n180 ) , .ZN( us00_n306 ) , .A( us00_n65 ) , .B1( us00_n71 ) );
  NOR2_X1 us00_U263 (.ZN( us00_n222 ) , .A2( us00_n62 ) , .A1( us00_n87 ) );
  INV_X1 us00_U264 (.ZN( us00_n11 ) , .A( us00_n114 ) );
  AOI21_X1 us00_U265 (.A( us00_n180 ) , .B1( us00_n208 ) , .ZN( us00_n325 ) , .B2( us00_n72 ) );
  NOR2_X1 us00_U266 (.A2( us00_n169 ) , .ZN( us00_n209 ) , .A1( us00_n87 ) );
  NOR2_X1 us00_U267 (.A1( us00_n130 ) , .ZN( us00_n221 ) , .A2( us00_n97 ) );
  NOR2_X1 us00_U268 (.A1( us00_n115 ) , .ZN( us00_n335 ) , .A2( us00_n86 ) );
  NOR2_X1 us00_U269 (.ZN( us00_n176 ) , .A1( us00_n60 ) , .A2( us00_n91 ) );
  NOR2_X1 us00_U27 (.ZN( us00_n197 ) , .A1( us00_n38 ) , .A2( us00_n43 ) );
  NOR2_X1 us00_U270 (.A2( us00_n153 ) , .ZN( us00_n268 ) , .A1( us00_n60 ) );
  NOR2_X1 us00_U271 (.ZN( us00_n112 ) , .A1( us00_n147 ) , .A2( us00_n91 ) );
  AOI21_X1 us00_U272 (.ZN( us00_n59 ) , .B1( us00_n60 ) , .B2( us00_n61 ) , .A( us00_n62 ) );
  INV_X1 us00_U273 (.A( us00_n148 ) , .ZN( us00_n9 ) );
  NOR2_X1 us00_U274 (.A1( us00_n147 ) , .A2( us00_n169 ) , .ZN( us00_n298 ) );
  NOR2_X1 us00_U275 (.A1( us00_n147 ) , .A2( us00_n153 ) , .ZN( us00_n344 ) );
  AOI21_X1 us00_U276 (.A( us00_n114 ) , .ZN( us00_n250 ) , .B1( us00_n252 ) , .B2( us00_n63 ) );
  AOI21_X1 us00_U277 (.ZN( us00_n58 ) , .B1( us00_n63 ) , .B2( us00_n64 ) , .A( us00_n65 ) );
  AOI21_X1 us00_U278 (.B1( us00_n127 ) , .A( us00_n148 ) , .ZN( us00_n362 ) , .B2( us00_n74 ) );
  AOI21_X1 us00_U279 (.B1( us00_n197 ) , .ZN( us00_n378 ) , .B2( us00_n61 ) , .A( us00_n65 ) );
  AOI222_X1 us00_U28 (.B2( us00_n12 ) , .A2( us00_n22 ) , .C2( us00_n26 ) , .C1( us00_n35 ) , .A1( us00_n38 ) , .ZN( us00_n408 ) , .B1( us00_n45 ) );
  AOI21_X1 us00_U280 (.ZN( us00_n227 ) , .B2( us00_n72 ) , .B1( us00_n85 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U281 (.A( us00_n128 ) , .B2( us00_n180 ) , .ZN( us00_n399 ) , .B1( us00_n98 ) );
  NOR2_X1 us00_U282 (.A1( us00_n133 ) , .ZN( us00_n295 ) , .A2( us00_n62 ) );
  NOR2_X1 us00_U283 (.ZN( us00_n235 ) , .A1( us00_n86 ) , .A2( us00_n89 ) );
  AOI21_X1 us00_U284 (.B1( us00_n127 ) , .ZN( us00_n284 ) , .B2( us00_n64 ) , .A( us00_n85 ) );
  NOR2_X1 us00_U285 (.A1( us00_n115 ) , .A2( us00_n169 ) , .ZN( us00_n83 ) );
  AOI21_X1 us00_U286 (.B2( us00_n208 ) , .ZN( us00_n251 ) , .B1( us00_n86 ) , .A( us00_n87 ) );
  NOR2_X1 us00_U287 (.A2( us00_n169 ) , .ZN( us00_n357 ) , .A1( us00_n63 ) );
  AOI21_X1 us00_U288 (.B1( us00_n127 ) , .A( us00_n208 ) , .ZN( us00_n400 ) , .B2( us00_n71 ) );
  NOR2_X1 us00_U289 (.ZN( us00_n318 ) , .A1( us00_n74 ) , .A2( us00_n86 ) );
  NOR4_X1 us00_U29 (.A3( us00_n263 ) , .A2( us00_n323 ) , .A4( us00_n335 ) , .ZN( us00_n410 ) , .A1( us00_n411 ) );
  NOR2_X1 us00_U290 (.A2( us00_n178 ) , .ZN( us00_n358 ) , .A1( us00_n61 ) );
  NOR2_X1 us00_U291 (.A2( us00_n178 ) , .ZN( us00_n194 ) , .A1( us00_n74 ) );
  NOR2_X1 us00_U292 (.A1( us00_n115 ) , .ZN( us00_n224 ) , .A2( us00_n91 ) );
  INV_X1 us00_U293 (.ZN( us00_n41 ) , .A( us00_n64 ) );
  AOI21_X1 us00_U294 (.A( us00_n147 ) , .B2( us00_n208 ) , .ZN( us00_n367 ) , .B1( us00_n62 ) );
  AOI21_X1 us00_U295 (.ZN( us00_n338 ) , .B1( us00_n62 ) , .A( us00_n63 ) , .B2( us00_n65 ) );
  AOI21_X1 us00_U296 (.A( us00_n114 ) , .ZN( us00_n337 ) , .B1( us00_n60 ) , .B2( us00_n98 ) );
  NOR2_X1 us00_U297 (.A1( us00_n208 ) , .ZN( us00_n296 ) , .A2( us00_n89 ) );
  AOI21_X1 us00_U298 (.B2( us00_n178 ) , .ZN( us00_n288 ) , .A( us00_n60 ) , .B1( us00_n62 ) );
  AOI21_X1 us00_U299 (.B2( us00_n114 ) , .A( us00_n145 ) , .ZN( us00_n177 ) , .B1( us00_n178 ) );
  NAND2_X1 us00_U3 (.ZN( us00_n169 ) , .A2( us00_n413 ) , .A1( us00_n436 ) );
  AOI221_X1 us00_U30 (.A( us00_n13 ) , .C2( us00_n163 ) , .B1( us00_n17 ) , .C1( us00_n32 ) , .ZN( us00_n409 ) , .B2( us00_n46 ) );
  AOI21_X1 us00_U300 (.B2( us00_n114 ) , .ZN( us00_n286 ) , .B1( us00_n65 ) , .A( us00_n92 ) );
  AOI21_X1 us00_U301 (.B2( us00_n115 ) , .A( us00_n153 ) , .ZN( us00_n379 ) , .B1( us00_n63 ) );
  NOR2_X1 us00_U302 (.A2( us00_n133 ) , .A1( us00_n178 ) , .ZN( us00_n330 ) );
  INV_X1 us00_U303 (.ZN( us00_n4 ) , .A( us00_n86 ) );
  INV_X1 us00_U304 (.ZN( us00_n23 ) , .A( us00_n65 ) );
  AOI21_X1 us00_U305 (.B2( us00_n130 ) , .ZN( us00_n237 ) , .B1( us00_n74 ) , .A( us00_n85 ) );
  AOI21_X1 us00_U306 (.B2( us00_n114 ) , .B1( us00_n148 ) , .ZN( us00_n228 ) , .A( us00_n64 ) );
  NOR2_X1 us00_U307 (.A1( us00_n148 ) , .ZN( us00_n192 ) , .A2( us00_n61 ) );
  AOI21_X1 us00_U308 (.B2( us00_n116 ) , .A( us00_n149 ) , .ZN( us00_n190 ) , .B1( us00_n191 ) );
  AOI21_X1 us00_U309 (.B2( us00_n115 ) , .B1( us00_n127 ) , .ZN( us00_n308 ) , .A( us00_n97 ) );
  NOR4_X1 us00_U31 (.ZN( us00_n353 ) , .A1( us00_n360 ) , .A2( us00_n361 ) , .A3( us00_n362 ) , .A4( us00_n363 ) );
  AOI21_X1 us00_U310 (.B1( us00_n169 ) , .A( us00_n180 ) , .ZN( us00_n377 ) , .B2( us00_n91 ) );
  NOR2_X1 us00_U311 (.A2( us00_n115 ) , .A1( us00_n148 ) , .ZN( us00_n309 ) );
  NOR2_X1 us00_U312 (.A2( us00_n180 ) , .ZN( us00_n297 ) , .A1( us00_n86 ) );
  NOR2_X1 us00_U313 (.A1( us00_n114 ) , .A2( us00_n180 ) , .ZN( us00_n311 ) );
  AOI21_X1 us00_U314 (.ZN( us00_n363 ) , .B1( us00_n65 ) , .B2( us00_n85 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U315 (.B2( us00_n128 ) , .ZN( us00_n238 ) , .B1( us00_n65 ) , .A( us00_n89 ) );
  INV_X1 us00_U316 (.A( us00_n178 ) , .ZN( us00_n24 ) );
  NOR2_X1 us00_U317 (.ZN( us00_n212 ) , .A2( us00_n64 ) , .A1( us00_n97 ) );
  AOI21_X1 us00_U318 (.ZN( us00_n427 ) , .B1( us00_n62 ) , .A( us00_n74 ) , .B2( us00_n85 ) );
  NOR2_X1 us00_U319 (.A1( us00_n153 ) , .A2( us00_n180 ) , .ZN( us00_n245 ) );
  AOI222_X1 us00_U32 (.B1( us00_n11 ) , .A2( us00_n25 ) , .C2( us00_n27 ) , .C1( us00_n33 ) , .ZN( us00_n352 ) , .B2( us00_n40 ) , .A1( us00_n43 ) );
  AOI21_X1 us00_U320 (.B1( us00_n153 ) , .ZN( us00_n313 ) , .B2( us00_n86 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U321 (.ZN( us00_n380 ) , .B1( us00_n73 ) , .B2( us00_n86 ) , .A( us00_n98 ) );
  NAND2_X1 us00_U322 (.A1( us00_n114 ) , .ZN( us00_n124 ) , .A2( us00_n72 ) );
  NOR2_X1 us00_U323 (.A1( us00_n169 ) , .ZN( us00_n348 ) , .A2( us00_n98 ) );
  NOR2_X1 us00_U324 (.A1( us00_n169 ) , .ZN( us00_n299 ) , .A2( us00_n64 ) );
  AOI21_X1 us00_U325 (.B1( us00_n114 ) , .B2( us00_n128 ) , .ZN( us00_n188 ) , .A( us00_n71 ) );
  NOR2_X1 us00_U326 (.A1( us00_n130 ) , .ZN( us00_n310 ) , .A2( us00_n72 ) );
  NOR2_X1 us00_U327 (.ZN( us00_n193 ) , .A2( us00_n64 ) , .A1( us00_n86 ) );
  NOR2_X1 us00_U328 (.ZN( us00_n56 ) , .A1( us00_n62 ) , .A2( us00_n64 ) );
  AOI21_X1 us00_U329 (.ZN( us00_n84 ) , .B1( us00_n85 ) , .B2( us00_n86 ) , .A( us00_n87 ) );
  NOR4_X1 us00_U33 (.A4( us00_n108 ) , .A2( us00_n204 ) , .ZN( us00_n354 ) , .A1( us00_n355 ) , .A3( us00_n356 ) );
  AOI21_X1 us00_U330 (.ZN( us00_n143 ) , .A( us00_n144 ) , .B1( us00_n85 ) , .B2( us00_n97 ) );
  AOI21_X1 us00_U331 (.B1( us00_n197 ) , .ZN( us00_n236 ) , .B2( us00_n60 ) , .A( us00_n86 ) );
  NOR2_X1 us00_U332 (.A2( us00_n114 ) , .A1( us00_n115 ) , .ZN( us00_n166 ) );
  NOR2_X1 us00_U333 (.ZN( us00_n294 ) , .A2( us00_n60 ) , .A1( us00_n85 ) );
  NOR2_X1 us00_U334 (.A1( us00_n153 ) , .ZN( us00_n343 ) , .A2( us00_n89 ) );
  NOR2_X1 us00_U335 (.A2( us00_n169 ) , .ZN( us00_n195 ) , .A1( us00_n60 ) );
  INV_X1 us00_U336 (.A( us00_n180 ) , .ZN( us00_n39 ) );
  INV_X1 us00_U337 (.ZN( us00_n22 ) , .A( us00_n62 ) );
  AOI21_X1 us00_U338 (.B2( us00_n127 ) , .B1( us00_n144 ) , .A( us00_n178 ) , .ZN( us00_n435 ) );
  OAI21_X1 us00_U339 (.B2( us00_n127 ) , .ZN( us00_n175 ) , .A( us00_n179 ) , .B1( us00_n73 ) );
  NOR4_X1 us00_U34 (.ZN( us00_n139 ) , .A1( us00_n140 ) , .A2( us00_n141 ) , .A3( us00_n142 ) , .A4( us00_n143 ) );
  OAI21_X1 us00_U340 (.A( us00_n17 ) , .ZN( us00_n179 ) , .B1( us00_n39 ) , .B2( us00_n44 ) );
  INV_X1 us00_U341 (.ZN( us00_n27 ) , .A( us00_n97 ) );
  INV_X1 us00_U342 (.ZN( us00_n31 ) , .A( us00_n92 ) );
  AOI22_X1 us00_U343 (.B1( us00_n14 ) , .A1( us00_n43 ) , .B2( us00_n46 ) , .ZN( us00_n94 ) , .A2( us00_n95 ) );
  NAND2_X1 us00_U344 (.ZN( us00_n206 ) , .A2( us00_n61 ) , .A1( us00_n71 ) );
  NAND2_X1 us00_U345 (.A1( us00_n149 ) , .ZN( us00_n163 ) , .A2( us00_n97 ) );
  NAND2_X1 us00_U346 (.A2( us00_n115 ) , .ZN( us00_n67 ) , .A1( us00_n71 ) );
  AOI21_X1 us00_U347 (.ZN( us00_n434 ) , .A( us00_n63 ) , .B2( us00_n86 ) , .B1( us00_n88 ) );
  NOR2_X1 us00_U348 (.ZN( us00_n393 ) , .A2( us00_n72 ) , .A1( us00_n89 ) );
  NOR2_X1 us00_U349 (.ZN( us00_n407 ) , .A1( us00_n62 ) , .A2( us00_n98 ) );
  AOI211_X1 us00_U35 (.ZN( us00_n138 ) , .A( us00_n151 ) , .B( us00_n152 ) , .C2( us00_n22 ) , .C1( us00_n34 ) );
  OAI21_X1 us00_U350 (.ZN( us00_n82 ) , .B1( us00_n88 ) , .B2( us00_n89 ) , .A( us00_n90 ) );
  OAI21_X1 us00_U351 (.B1( us00_n14 ) , .A( us00_n38 ) , .B2( us00_n4 ) , .ZN( us00_n90 ) );
  NOR2_X1 us00_U352 (.A2( us00_n153 ) , .ZN( us00_n165 ) , .A1( us00_n87 ) );
  NOR2_X1 us00_U353 (.A2( us00_n127 ) , .A1( us00_n153 ) , .ZN( us00_n351 ) );
  NAND2_X1 us00_U354 (.A2( us00_n148 ) , .A1( us00_n178 ) , .ZN( us00_n95 ) );
  NOR2_X1 us00_U355 (.A1( us00_n169 ) , .ZN( us00_n359 ) , .A2( us00_n89 ) );
  OAI21_X1 us00_U356 (.ZN( us00_n141 ) , .B1( us00_n145 ) , .A( us00_n146 ) , .B2( us00_n72 ) );
  OAI21_X1 us00_U357 (.ZN( us00_n146 ) , .B2( us00_n25 ) , .B1( us00_n4 ) , .A( us00_n44 ) );
  NAND2_X1 us00_U358 (.A2( us00_n128 ) , .ZN( us00_n68 ) , .A1( us00_n91 ) );
  INV_X1 us00_U359 (.ZN( us00_n33 ) , .A( us00_n60 ) );
  NOR3_X1 us00_U36 (.A2( us00_n136 ) , .ZN( us00_n137 ) , .A1( us00_n154 ) , .A3( us00_n155 ) );
  INV_X1 us00_U360 (.A( us00_n153 ) , .ZN( us00_n21 ) );
  AND2_X1 us00_U361 (.ZN( us00_n145 ) , .A2( us00_n92 ) , .A1( us00_n98 ) );
  AOI221_X1 us00_U362 (.ZN( us00_n103 ) , .B1( us00_n11 ) , .A( us00_n113 ) , .C1( us00_n22 ) , .B2( us00_n42 ) , .C2( us00_n67 ) );
  AOI21_X1 us00_U363 (.ZN( us00_n113 ) , .B2( us00_n114 ) , .B1( us00_n85 ) , .A( us00_n89 ) );
  INV_X1 us00_U364 (.A( us00_n116 ) , .ZN( us00_n42 ) );
  NAND2_X1 us00_U365 (.A2( us00_n428 ) , .A1( us00_n430 ) , .ZN( us00_n72 ) );
  NAND2_X1 us00_U366 (.A2( us00_n406 ) , .A1( us00_n422 ) , .ZN( us00_n74 ) );
  NAND2_X1 us00_U367 (.A2( us00_n423 ) , .A1( us00_n426 ) , .ZN( us00_n63 ) );
  NAND2_X1 us00_U368 (.A2( us00_n406 ) , .A1( us00_n426 ) , .ZN( us00_n61 ) );
  NAND2_X1 us00_U369 (.A2( us00_n416 ) , .A1( us00_n423 ) , .ZN( us00_n64 ) );
  NOR4_X1 us00_U37 (.ZN( us00_n119 ) , .A1( us00_n120 ) , .A2( us00_n121 ) , .A3( us00_n122 ) , .A4( us00_n8 ) );
  NAND2_X1 us00_U370 (.ZN( us00_n133 ) , .A2( us00_n416 ) , .A1( us00_n424 ) );
  NAND2_X1 us00_U371 (.ZN( us00_n208 ) , .A2( us00_n412 ) , .A1( us00_n425 ) );
  NAND2_X1 us00_U372 (.ZN( us00_n149 ) , .A1( us00_n417 ) , .A2( us00_n429 ) );
  NAND2_X1 us00_U373 (.ZN( us00_n127 ) , .A2( us00_n415 ) , .A1( us00_n422 ) );
  NAND2_X1 us00_U374 (.A1( us00_n422 ) , .A2( us00_n424 ) , .ZN( us00_n71 ) );
  NAND2_X1 us00_U375 (.A1( us00_n405 ) , .A2( us00_n423 ) , .ZN( us00_n98 ) );
  NAND2_X1 us00_U376 (.A2( us00_n405 ) , .A1( us00_n424 ) , .ZN( us00_n92 ) );
  NAND2_X1 us00_U377 (.A1( us00_n412 ) , .A2( us00_n413 ) , .ZN( us00_n65 ) );
  NAND2_X1 us00_U378 (.ZN( us00_n178 ) , .A2( us00_n417 ) , .A1( us00_n436 ) );
  NAND2_X1 us00_U379 (.ZN( us00_n114 ) , .A1( us00_n425 ) , .A2( us00_n428 ) );
  AOI211_X1 us00_U38 (.ZN( us00_n118 ) , .A( us00_n131 ) , .B( us00_n132 ) , .C2( us00_n24 ) , .C1( us00_n45 ) );
  NAND2_X2 us00_U380 (.ZN( us00_n180 ) , .A1( us00_n406 ) , .A2( us00_n416 ) );
  NAND2_X1 us00_U381 (.ZN( us00_n148 ) , .A1( us00_n425 ) , .A2( us00_n429 ) );
  NAND2_X1 us00_U382 (.ZN( us00_n130 ) , .A1( us00_n415 ) , .A2( us00_n416 ) );
  NAND2_X1 us00_U383 (.A2( us00_n405 ) , .A1( us00_n415 ) , .ZN( us00_n89 ) );
  NOR2_X1 us00_U384 (.A1( us00_n29 ) , .A2( us00_n30 ) , .ZN( us00_n412 ) );
  NOR2_X1 us00_U385 (.ZN( us00_n424 ) , .A2( us00_n50 ) , .A1( us00_n51 ) );
  NOR2_X1 us00_U386 (.ZN( us00_n426 ) , .A2( us00_n48 ) , .A1( us00_n49 ) );
  NAND2_X1 us00_U388 (.ZN( us00_n147 ) , .A1( us00_n422 ) , .A2( us00_n423 ) );
  NAND2_X1 us00_U389 (.A2( us00_n415 ) , .A1( us00_n426 ) , .ZN( us00_n87 ) );
  NOR3_X1 us00_U39 (.ZN( us00_n117 ) , .A1( us00_n134 ) , .A2( us00_n135 ) , .A3( us00_n136 ) );
  NAND2_X2 us00_U390 (.A1( us00_n413 ) , .A2( us00_n429 ) , .ZN( us00_n62 ) );
  NAND2_X2 us00_U391 (.A1( us00_n425 ) , .A2( us00_n436 ) , .ZN( us00_n86 ) );
  NAND2_X2 us00_U392 (.ZN( us00_n153 ) , .A2( us00_n413 ) , .A1( us00_n428 ) );
  NAND2_X1 us00_U393 (.A1( us00_n430 ) , .A2( us00_n436 ) , .ZN( us00_n93 ) );
  NAND2_X2 us00_U394 (.A2( us00_n417 ) , .A1( us00_n428 ) , .ZN( us00_n85 ) );
  NAND2_X2 us00_U395 (.A1( us00_n412 ) , .A2( us00_n417 ) , .ZN( us00_n97 ) );
  NAND2_X1 us00_U396 (.A2( us00_n429 ) , .A1( us00_n430 ) , .ZN( us00_n91 ) );
  NOR2_X1 us00_U397 (.A2( sa00_6 ) , .A1( sa00_7 ) , .ZN( us00_n413 ) );
  NOR2_X1 us00_U398 (.A2( sa00_5 ) , .A1( us00_n30 ) , .ZN( us00_n429 ) );
  NAND2_X1 us00_U4 (.A1( us00_n405 ) , .A2( us00_n406 ) , .ZN( us00_n60 ) );
  AOI221_X1 us00_U40 (.C1( us00_n11 ) , .B1( us00_n12 ) , .B2( us00_n39 ) , .C2( us00_n40 ) , .ZN( us00_n79 ) , .A( us00_n96 ) );
  NOR2_X1 us00_U400 (.A2( sa00_4 ) , .A1( us00_n29 ) , .ZN( us00_n428 ) );
  NOR2_X1 us00_U401 (.A2( sa00_4 ) , .A1( sa00_5 ) , .ZN( us00_n436 ) );
  NOR2_X1 us00_U402 (.A2( sa00_1 ) , .ZN( us00_n406 ) , .A1( us00_n51 ) );
  NOR2_X1 us00_U403 (.A2( sa00_2 ) , .A1( sa00_3 ) , .ZN( us00_n405 ) );
  NOR2_X1 us00_U405 (.A2( sa00_2 ) , .ZN( us00_n416 ) , .A1( us00_n48 ) );
  NOR2_X1 us00_U406 (.A2( sa00_0 ) , .ZN( us00_n423 ) , .A1( us00_n50 ) );
  NOR2_X1 us00_U407 (.A2( sa00_0 ) , .A1( sa00_1 ) , .ZN( us00_n415 ) );
  NOR2_X1 us00_U408 (.A2( sa00_3 ) , .ZN( us00_n422 ) , .A1( us00_n49 ) );
  NOR4_X1 us00_U41 (.ZN( us00_n80 ) , .A1( us00_n81 ) , .A2( us00_n82 ) , .A3( us00_n83 ) , .A4( us00_n84 ) );
  INV_X1 us00_U410 (.A( sa00_1 ) , .ZN( us00_n50 ) );
  INV_X1 us00_U411 (.A( sa00_3 ) , .ZN( us00_n48 ) );
  INV_X1 us00_U412 (.A( sa00_2 ) , .ZN( us00_n49 ) );
  INV_X1 us00_U413 (.A( sa00_0 ) , .ZN( us00_n51 ) );
  INV_X1 us00_U414 (.A( sa00_5 ) , .ZN( us00_n29 ) );
  OAI221_X1 us00_U416 (.C1( us00_n64 ) , .ZN( us00_n81 ) , .B1( us00_n91 ) , .B2( us00_n92 ) , .C2( us00_n93 ) , .A( us00_n94 ) );
  NAND2_X1 us00_U417 (.A1( us00_n148 ) , .ZN( us00_n66 ) , .A2( us00_n93 ) );
  OAI22_X1 us00_U418 (.A1( us00_n114 ) , .B2( us00_n115 ) , .A2( us00_n130 ) , .ZN( us00_n289 ) , .B1( us00_n93 ) );
  OAI221_X1 us00_U419 (.ZN( us00_n174 ) , .A( us00_n181 ) , .B2( us00_n71 ) , .B1( us00_n91 ) , .C1( us00_n92 ) , .C2( us00_n93 ) );
  NOR4_X1 us00_U42 (.A3( us00_n100 ) , .A4( us00_n101 ) , .A2( us00_n76 ) , .ZN( us00_n78 ) , .A1( us00_n99 ) );
  AOI21_X1 us00_U420 (.B1( us00_n149 ) , .ZN( us00_n285 ) , .A( us00_n87 ) , .B2( us00_n93 ) );
  AOI21_X1 us00_U421 (.B1( us00_n178 ) , .ZN( us00_n254 ) , .B2( us00_n93 ) , .A( us00_n98 ) );
  AOI21_X1 us00_U422 (.A( us00_n115 ) , .ZN( us00_n229 ) , .B1( us00_n85 ) , .B2( us00_n93 ) );
  OAI22_X1 us00_U423 (.A2( us00_n147 ) , .A1( us00_n178 ) , .ZN( us00_n196 ) , .B1( us00_n60 ) , .B2( us00_n93 ) );
  OAI21_X1 us00_U424 (.B1( us00_n252 ) , .ZN( us00_n261 ) , .A( us00_n264 ) , .B2( us00_n93 ) );
  NOR2_X1 us00_U425 (.ZN( us00_n267 ) , .A2( us00_n61 ) , .A1( us00_n93 ) );
  OAI222_X1 us00_U426 (.B1( us00_n130 ) , .ZN( us00_n203 ) , .A2( us00_n208 ) , .A1( us00_n60 ) , .C1( us00_n62 ) , .C2( us00_n89 ) , .B2( us00_n93 ) );
  NOR2_X1 us00_U427 (.ZN( us00_n226 ) , .A2( us00_n89 ) , .A1( us00_n93 ) );
  NOR2_X1 us00_U428 (.A2( us00_n180 ) , .ZN( us00_n277 ) , .A1( us00_n93 ) );
  NOR2_X1 us00_U429 (.A2( us00_n133 ) , .ZN( us00_n324 ) , .A1( us00_n93 ) );
  NOR2_X1 us00_U43 (.A2( us00_n16 ) , .A1( us00_n23 ) , .ZN( us00_n73 ) );
  INV_X1 us00_U430 (.ZN( us00_n16 ) , .A( us00_n93 ) );
  NAND4_X1 us00_U431 (.ZN( sa00_sr_2 ) , .A2( us00_n231 ) , .A1( us00_n232 ) , .A3( us00_n233 ) , .A4( us00_n234 ) );
  AOI221_X1 us00_U432 (.C1( us00_n16 ) , .B1( us00_n23 ) , .ZN( us00_n290 ) , .A( us00_n301 ) , .C2( us00_n34 ) , .B2( us00_n46 ) );
  AOI21_X1 us00_U433 (.B1( us00_n129 ) , .B2( us00_n153 ) , .ZN( us00_n301 ) , .A( us00_n92 ) );
  AOI211_X1 us00_U434 (.B( us00_n134 ) , .C1( us00_n23 ) , .ZN( us00_n232 ) , .A( us00_n240 ) , .C2( us00_n38 ) );
  NAND4_X1 us00_U435 (.ZN( us00_n134 ) , .A1( us00_n241 ) , .A2( us00_n242 ) , .A3( us00_n243 ) , .A4( us00_n244 ) );
  INV_X1 us00_U436 (.A( sa00_4 ) , .ZN( us00_n30 ) );
  NAND3_X1 us00_U437 (.ZN( sa00_sr_6 ) , .A1( us00_n78 ) , .A2( us00_n79 ) , .A3( us00_n80 ) );
  NAND3_X1 us00_U438 (.ZN( sa00_sr_5 ) , .A1( us00_n117 ) , .A2( us00_n118 ) , .A3( us00_n119 ) );
  NAND3_X1 us00_U439 (.ZN( sa00_sr_4 ) , .A1( us00_n137 ) , .A2( us00_n138 ) , .A3( us00_n139 ) );
  NAND4_X1 us00_U44 (.ZN( sa00_sr_3 ) , .A1( us00_n170 ) , .A2( us00_n171 ) , .A3( us00_n172 ) , .A4( us00_n173 ) );
  NAND3_X1 us00_U440 (.A1( us00_n200 ) , .A2( us00_n201 ) , .A3( us00_n202 ) , .ZN( us00_n70 ) );
  NAND3_X1 us00_U441 (.A2( us00_n153 ) , .A3( us00_n169 ) , .ZN( us00_n239 ) , .A1( us00_n85 ) );
  NAND3_X1 us00_U442 (.ZN( us00_n152 ) , .A1( us00_n257 ) , .A2( us00_n258 ) , .A3( us00_n259 ) );
  NAND3_X1 us00_U443 (.ZN( us00_n256 ) , .A1( us00_n290 ) , .A2( us00_n291 ) , .A3( us00_n292 ) );
  NAND3_X1 us00_U444 (.A2( us00_n127 ) , .A3( us00_n197 ) , .ZN( us00_n312 ) , .A1( us00_n92 ) );
  NAND3_X1 us00_U445 (.ZN( us00_n135 ) , .A1( us00_n352 ) , .A2( us00_n353 ) , .A3( us00_n354 ) );
  NAND3_X1 us00_U446 (.ZN( us00_n269 ) , .A1( us00_n364 ) , .A3( us00_n365 ) , .A2( us00_n6 ) );
  NAND3_X1 us00_U447 (.ZN( us00_n100 ) , .A1( us00_n408 ) , .A2( us00_n409 ) , .A3( us00_n410 ) );
  NOR4_X1 us00_U45 (.ZN( us00_n173 ) , .A1( us00_n174 ) , .A2( us00_n175 ) , .A3( us00_n176 ) , .A4( us00_n177 ) );
  AOI211_X1 us00_U46 (.ZN( us00_n172 ) , .A( us00_n182 ) , .B( us00_n183 ) , .C1( us00_n26 ) , .C2( us00_n46 ) );
  NOR2_X1 us00_U47 (.A2( us00_n101 ) , .ZN( us00_n170 ) , .A1( us00_n77 ) );
  NAND4_X1 us00_U48 (.ZN( sa00_sr_7 ) , .A1( us00_n52 ) , .A2( us00_n53 ) , .A3( us00_n54 ) , .A4( us00_n55 ) );
  NOR4_X1 us00_U49 (.ZN( us00_n55 ) , .A1( us00_n56 ) , .A2( us00_n57 ) , .A3( us00_n58 ) , .A4( us00_n59 ) );
  NOR3_X1 us00_U5 (.A2( us00_n135 ) , .A3( us00_n154 ) , .A1( us00_n269 ) , .ZN( us00_n279 ) );
  AOI222_X1 us00_U50 (.B1( us00_n24 ) , .A1( us00_n38 ) , .C1( us00_n45 ) , .ZN( us00_n54 ) , .A2( us00_n66 ) , .B2( us00_n67 ) , .C2( us00_n68 ) );
  AOI211_X1 us00_U51 (.C2( us00_n27 ) , .C1( us00_n35 ) , .ZN( us00_n53 ) , .A( us00_n69 ) , .B( us00_n70 ) );
  NOR2_X1 us00_U52 (.ZN( us00_n129 ) , .A2( us00_n15 ) , .A1( us00_n16 ) );
  NAND4_X1 us00_U53 (.ZN( sa00_sr_0 ) , .A1( us00_n373 ) , .A2( us00_n374 ) , .A3( us00_n375 ) , .A4( us00_n376 ) );
  AOI221_X1 us00_U54 (.B1( us00_n15 ) , .C2( us00_n17 ) , .C1( us00_n31 ) , .B2( us00_n34 ) , .ZN( us00_n375 ) , .A( us00_n380 ) );
  NOR4_X1 us00_U55 (.A1( us00_n350 ) , .ZN( us00_n376 ) , .A2( us00_n377 ) , .A3( us00_n378 ) , .A4( us00_n379 ) );
  AOI211_X1 us00_U56 (.C1( us00_n26 ) , .ZN( us00_n374 ) , .C2( us00_n38 ) , .A( us00_n381 ) , .B( us00_n75 ) );
  NAND4_X1 us00_U57 (.ZN( sa00_sr_1 ) , .A1( us00_n279 ) , .A2( us00_n280 ) , .A3( us00_n281 ) , .A4( us00_n282 ) );
  NOR4_X1 us00_U58 (.ZN( us00_n282 ) , .A1( us00_n283 ) , .A2( us00_n284 ) , .A3( us00_n285 ) , .A4( us00_n286 ) );
  AOI211_X1 us00_U59 (.ZN( us00_n281 ) , .A( us00_n287 ) , .B( us00_n288 ) , .C1( us00_n44 ) , .C2( us00_n66 ) );
  NOR3_X1 us00_U6 (.ZN( us00_n52 ) , .A1( us00_n75 ) , .A2( us00_n76 ) , .A3( us00_n77 ) );
  AOI211_X1 us00_U60 (.C2( us00_n22 ) , .B( us00_n256 ) , .ZN( us00_n280 ) , .A( us00_n289 ) , .C1( us00_n32 ) );
  NOR2_X1 us00_U61 (.ZN( us00_n252 ) , .A1( us00_n38 ) , .A2( us00_n41 ) );
  NAND4_X1 us00_U62 (.ZN( us00_n155 ) , .A1( us00_n271 ) , .A2( us00_n272 ) , .A3( us00_n273 ) , .A4( us00_n274 ) );
  NOR3_X1 us00_U63 (.A2( us00_n107 ) , .A3( us00_n214 ) , .ZN( us00_n273 ) , .A1( us00_n278 ) );
  NOR4_X1 us00_U64 (.A4( us00_n222 ) , .ZN( us00_n274 ) , .A1( us00_n275 ) , .A2( us00_n276 ) , .A3( us00_n277 ) );
  AOI222_X1 us00_U65 (.B2( us00_n16 ) , .A2( us00_n21 ) , .ZN( us00_n271 ) , .B1( us00_n35 ) , .C2( us00_n40 ) , .A1( us00_n47 ) , .C1( us00_n9 ) );
  NOR4_X1 us00_U66 (.A1( us00_n194 ) , .ZN( us00_n291 ) , .A2( us00_n298 ) , .A3( us00_n299 ) , .A4( us00_n300 ) );
  NOR4_X1 us00_U67 (.A4( us00_n110 ) , .A2( us00_n215 ) , .A3( us00_n225 ) , .ZN( us00_n292 ) , .A1( us00_n293 ) );
  AOI211_X1 us00_U68 (.C1( us00_n14 ) , .ZN( us00_n242 ) , .A( us00_n253 ) , .B( us00_n254 ) , .C2( us00_n41 ) );
  NOR4_X1 us00_U69 (.ZN( us00_n244 ) , .A1( us00_n245 ) , .A2( us00_n246 ) , .A3( us00_n247 ) , .A4( us00_n248 ) );
  NOR3_X1 us00_U7 (.A1( us00_n1 ) , .A3( us00_n100 ) , .A2( us00_n198 ) , .ZN( us00_n373 ) );
  NOR4_X1 us00_U70 (.A1( us00_n213 ) , .ZN( us00_n243 ) , .A2( us00_n249 ) , .A3( us00_n250 ) , .A4( us00_n251 ) );
  NAND4_X1 us00_U71 (.A1( us00_n217 ) , .A2( us00_n218 ) , .A3( us00_n219 ) , .A4( us00_n220 ) , .ZN( us00_n77 ) );
  NOR3_X1 us00_U72 (.ZN( us00_n218 ) , .A1( us00_n227 ) , .A2( us00_n228 ) , .A3( us00_n229 ) );
  NOR3_X1 us00_U73 (.ZN( us00_n219 ) , .A1( us00_n224 ) , .A2( us00_n225 ) , .A3( us00_n226 ) );
  NOR3_X1 us00_U74 (.ZN( us00_n220 ) , .A1( us00_n221 ) , .A2( us00_n222 ) , .A3( us00_n223 ) );
  NAND4_X1 us00_U75 (.ZN( us00_n270 ) , .A1( us00_n314 ) , .A2( us00_n315 ) , .A3( us00_n316 ) , .A4( us00_n317 ) );
  NOR4_X1 us00_U76 (.A2( us00_n109 ) , .A4( us00_n192 ) , .A3( us00_n216 ) , .A1( us00_n224 ) , .ZN( us00_n316 ) );
  NOR4_X1 us00_U77 (.ZN( us00_n315 ) , .A1( us00_n322 ) , .A2( us00_n323 ) , .A3( us00_n324 ) , .A4( us00_n325 ) );
  NOR4_X1 us00_U78 (.ZN( us00_n317 ) , .A1( us00_n318 ) , .A2( us00_n319 ) , .A3( us00_n320 ) , .A4( us00_n321 ) );
  NAND4_X1 us00_U79 (.A1( us00_n102 ) , .A2( us00_n103 ) , .A3( us00_n104 ) , .A4( us00_n105 ) , .ZN( us00_n76 ) );
  INV_X1 us00_U8 (.ZN( us00_n1 ) , .A( us00_n171 ) );
  NOR3_X1 us00_U80 (.ZN( us00_n104 ) , .A1( us00_n110 ) , .A2( us00_n111 ) , .A3( us00_n112 ) );
  NOR4_X1 us00_U81 (.ZN( us00_n105 ) , .A1( us00_n106 ) , .A2( us00_n107 ) , .A3( us00_n108 ) , .A4( us00_n109 ) );
  AOI222_X1 us00_U82 (.ZN( us00_n102 ) , .B1( us00_n16 ) , .A2( us00_n27 ) , .B2( us00_n36 ) , .C2( us00_n4 ) , .C1( us00_n43 ) , .A1( us00_n47 ) );
  NOR4_X1 us00_U83 (.ZN( us00_n201 ) , .A1( us00_n209 ) , .A2( us00_n210 ) , .A3( us00_n211 ) , .A4( us00_n212 ) );
  NOR4_X1 us00_U84 (.ZN( us00_n200 ) , .A1( us00_n213 ) , .A2( us00_n214 ) , .A3( us00_n215 ) , .A4( us00_n216 ) );
  NOR4_X1 us00_U85 (.A4( us00_n162 ) , .A2( us00_n18 ) , .ZN( us00_n202 ) , .A1( us00_n203 ) , .A3( us00_n204 ) );
  NOR2_X1 us00_U86 (.ZN( us00_n116 ) , .A2( us00_n43 ) , .A1( us00_n44 ) );
  AOI222_X1 us00_U87 (.A2( us00_n12 ) , .C1( us00_n14 ) , .ZN( us00_n233 ) , .B2( us00_n239 ) , .C2( us00_n31 ) , .A1( us00_n35 ) , .B1( us00_n36 ) );
  NOR4_X1 us00_U88 (.ZN( us00_n234 ) , .A1( us00_n235 ) , .A2( us00_n236 ) , .A3( us00_n237 ) , .A4( us00_n238 ) );
  NOR3_X1 us00_U89 (.A3( us00_n155 ) , .ZN( us00_n231 ) , .A1( us00_n269 ) , .A2( us00_n270 ) );
  NOR3_X1 us00_U9 (.A1( us00_n152 ) , .ZN( us00_n241 ) , .A2( us00_n255 ) , .A3( us00_n256 ) );
  AOI222_X1 us00_U90 (.A1( us00_n11 ) , .B1( us00_n14 ) , .C2( us00_n15 ) , .A2( us00_n34 ) , .ZN( us00_n364 ) , .B2( us00_n40 ) , .C1( us00_n45 ) );
  NOR4_X1 us00_U91 (.A3( us00_n207 ) , .ZN( us00_n365 ) , .A1( us00_n366 ) , .A2( us00_n367 ) , .A4( us00_n368 ) );
  INV_X1 us00_U92 (.A( us00_n372 ) , .ZN( us00_n6 ) );
  NAND4_X1 us00_U93 (.ZN( us00_n198 ) , .A1( us00_n418 ) , .A2( us00_n419 ) , .A3( us00_n420 ) , .A4( us00_n421 ) );
  NOR3_X1 us00_U94 (.A2( us00_n307 ) , .A1( us00_n322 ) , .A3( us00_n347 ) , .ZN( us00_n420 ) );
  AOI221_X1 us00_U95 (.C2( us00_n124 ) , .B2( us00_n16 ) , .C1( us00_n35 ) , .ZN( us00_n418 ) , .A( us00_n427 ) , .B1( us00_n45 ) );
  NOR4_X1 us00_U96 (.A3( us00_n166 ) , .A4( us00_n249 ) , .A1( us00_n278 ) , .A2( us00_n368 ) , .ZN( us00_n419 ) );
  NAND4_X1 us00_U97 (.ZN( us00_n255 ) , .A1( us00_n339 ) , .A2( us00_n340 ) , .A3( us00_n341 ) , .A4( us00_n342 ) );
  NOR4_X1 us00_U98 (.A3( us00_n176 ) , .ZN( us00_n339 ) , .A1( us00_n349 ) , .A2( us00_n350 ) , .A4( us00_n351 ) );
  NOR4_X1 us00_U99 (.A3( us00_n112 ) , .A4( us00_n209 ) , .A2( us00_n223 ) , .ZN( us00_n341 ) , .A1( us00_n346 ) );
  NOR3_X1 us13_U10 (.A3( us13_n621 ) , .A2( us13_n622 ) , .ZN( us13_n636 ) , .A1( us13_n725 ) );
  NOR4_X1 us13_U100 (.ZN( us13_n458 ) , .A2( us13_n509 ) , .A1( us13_n599 ) , .A4( us13_n628 ) , .A3( us13_n711 ) );
  NAND4_X1 us13_U101 (.A4( us13_n535 ) , .A3( us13_n536 ) , .A2( us13_n537 ) , .A1( us13_n538 ) , .ZN( us13_n622 ) );
  NOR4_X1 us13_U102 (.A4( us13_n526 ) , .A2( us13_n527 ) , .A1( us13_n528 ) , .ZN( us13_n538 ) , .A3( us13_n701 ) );
  NOR4_X1 us13_U103 (.A4( us13_n529 ) , .A3( us13_n530 ) , .ZN( us13_n537 ) , .A2( us13_n684 ) , .A1( us13_n794 ) );
  NOR4_X1 us13_U104 (.A4( us13_n532 ) , .A3( us13_n533 ) , .A2( us13_n534 ) , .ZN( us13_n535 ) , .A1( us13_n820 ) );
  NAND4_X1 us13_U105 (.A4( us13_n548 ) , .A3( us13_n549 ) , .A2( us13_n550 ) , .A1( us13_n551 ) , .ZN( us13_n745 ) );
  NOR3_X1 us13_U106 (.ZN( us13_n549 ) , .A2( us13_n651 ) , .A1( us13_n667 ) , .A3( us13_n771 ) );
  AOI211_X1 us13_U107 (.B( us13_n539 ) , .A( us13_n540 ) , .ZN( us13_n551 ) , .C2( us13_n839 ) , .C1( us13_n851 ) );
  NOR4_X1 us13_U108 (.A4( us13_n541 ) , .A3( us13_n542 ) , .A2( us13_n543 ) , .ZN( us13_n550 ) , .A1( us13_n688 ) );
  NAND4_X1 us13_U109 (.A4( us13_n479 ) , .A3( us13_n480 ) , .A2( us13_n481 ) , .A1( us13_n482 ) , .ZN( us13_n694 ) );
  NOR2_X1 us13_U11 (.A1( us13_n678 ) , .ZN( us13_n693 ) , .A2( us13_n807 ) );
  NOR3_X1 us13_U110 (.ZN( us13_n480 ) , .A2( us13_n508 ) , .A3( us13_n601 ) , .A1( us13_n610 ) );
  AOI211_X1 us13_U111 (.B( us13_n477 ) , .A( us13_n478 ) , .ZN( us13_n482 ) , .C2( us13_n833 ) , .C1( us13_n861 ) );
  NOR4_X1 us13_U112 (.ZN( us13_n481 ) , .A3( us13_n532 ) , .A4( us13_n545 ) , .A2( us13_n567 ) , .A1( us13_n717 ) );
  NOR2_X1 us13_U113 (.ZN( us13_n647 ) , .A1( us13_n854 ) , .A2( us13_n868 ) );
  NOR4_X1 us13_U114 (.ZN( us13_n620 ) , .A1( us13_n656 ) , .A3( us13_n666 ) , .A4( us13_n682 ) , .A2( us13_n766 ) );
  NOR4_X1 us13_U115 (.A4( us13_n609 ) , .A3( us13_n610 ) , .A2( us13_n611 ) , .A1( us13_n612 ) , .ZN( us13_n619 ) );
  NOR4_X1 us13_U116 (.A4( us13_n614 ) , .A3( us13_n615 ) , .A2( us13_n616 ) , .A1( us13_n617 ) , .ZN( us13_n618 ) );
  NOR2_X1 us13_U117 (.ZN( us13_n686 ) , .A1( us13_n831 ) , .A2( us13_n832 ) );
  NAND4_X1 us13_U118 (.A4( us13_n473 ) , .A3( us13_n474 ) , .A2( us13_n475 ) , .A1( us13_n476 ) , .ZN( us13_n678 ) );
  NOR4_X1 us13_U119 (.ZN( us13_n475 ) , .A1( us13_n531 ) , .A3( us13_n568 ) , .A4( us13_n600 ) , .A2( us13_n642 ) );
  INV_X1 us13_U12 (.A( us13_n607 ) , .ZN( us13_n874 ) );
  NOR4_X1 us13_U120 (.A4( us13_n470 ) , .ZN( us13_n476 ) , .A3( us13_n556 ) , .A1( us13_n735 ) , .A2( us13_n755 ) );
  NOR4_X1 us13_U121 (.ZN( us13_n474 ) , .A1( us13_n506 ) , .A3( us13_n544 ) , .A2( us13_n583 ) , .A4( us13_n716 ) );
  NOR2_X1 us13_U122 (.ZN( us13_n733 ) , .A2( us13_n832 ) , .A1( us13_n845 ) );
  NAND4_X1 us13_U123 (.A4( us13_n719 ) , .A3( us13_n720 ) , .A2( us13_n721 ) , .ZN( us13_n741 ) , .A1( us13_n857 ) );
  INV_X1 us13_U124 (.A( us13_n709 ) , .ZN( us13_n857 ) );
  NOR4_X1 us13_U125 (.A4( us13_n715 ) , .A3( us13_n716 ) , .A2( us13_n717 ) , .A1( us13_n718 ) , .ZN( us13_n719 ) );
  AOI221_X1 us13_U126 (.A( us13_n710 ) , .ZN( us13_n721 ) , .C2( us13_n844 ) , .B2( us13_n845 ) , .C1( us13_n861 ) , .B1( us13_n862 ) );
  NAND4_X1 us13_U127 (.A4( us13_n573 ) , .A3( us13_n574 ) , .A1( us13_n575 ) , .ZN( us13_n723 ) , .A2( us13_n874 ) );
  NOR4_X1 us13_U128 (.A4( us13_n569 ) , .A3( us13_n570 ) , .A2( us13_n571 ) , .A1( us13_n572 ) , .ZN( us13_n573 ) );
  AOI221_X1 us13_U129 (.A( us13_n564 ) , .C2( us13_n565 ) , .ZN( us13_n574 ) , .B2( us13_n845 ) , .B1( us13_n852 ) , .C1( us13_n853 ) );
  INV_X1 us13_U13 (.A( us13_n680 ) , .ZN( us13_n840 ) );
  NOR2_X1 us13_U130 (.ZN( us13_n575 ) , .A1( us13_n622 ) , .A2( us13_n745 ) );
  NAND4_X1 us13_U131 (.A4( us13_n633 ) , .A3( us13_n634 ) , .A2( us13_n635 ) , .A1( us13_n636 ) , .ZN( us13_n743 ) );
  AOI211_X1 us13_U132 (.B( us13_n623 ) , .A( us13_n624 ) , .ZN( us13_n635 ) , .C2( us13_n836 ) , .C1( us13_n863 ) );
  NOR4_X1 us13_U133 (.A4( us13_n629 ) , .A3( us13_n630 ) , .A2( us13_n631 ) , .A1( us13_n632 ) , .ZN( us13_n633 ) );
  NOR4_X1 us13_U134 (.A4( us13_n626 ) , .A3( us13_n627 ) , .A2( us13_n628 ) , .ZN( us13_n634 ) , .A1( us13_n664 ) );
  NAND4_X1 us13_U135 (.A4( us13_n493 ) , .A3( us13_n494 ) , .A1( us13_n495 ) , .ZN( us13_n802 ) , .A2( us13_n867 ) );
  AOI221_X1 us13_U136 (.A( us13_n489 ) , .ZN( us13_n494 ) , .B2( us13_n836 ) , .C2( us13_n841 ) , .C1( us13_n851 ) , .B1( us13_n860 ) );
  INV_X1 us13_U137 (.A( us13_n778 ) , .ZN( us13_n867 ) );
  NOR2_X1 us13_U138 (.ZN( us13_n495 ) , .A1( us13_n678 ) , .A2( us13_n694 ) );
  INV_X1 us13_U139 (.A( us13_n762 ) , .ZN( us13_n830 ) );
  NOR4_X1 us13_U14 (.A4( us13_n445 ) , .A3( us13_n446 ) , .A2( us13_n516 ) , .A1( us13_n541 ) , .ZN( us13_n706 ) );
  OR4_X1 us13_U140 (.A4( us13_n566 ) , .A3( us13_n567 ) , .A2( us13_n568 ) , .ZN( us13_n572 ) , .A1( us13_n665 ) );
  OR4_X1 us13_U141 (.A4( us13_n518 ) , .A2( us13_n519 ) , .A1( us13_n520 ) , .ZN( us13_n522 ) , .A3( us13_n821 ) );
  OR4_X1 us13_U142 (.ZN( us13_n466 ) , .A4( us13_n518 ) , .A3( us13_n529 ) , .A2( us13_n578 ) , .A1( us13_n712 ) );
  OR4_X1 us13_U143 (.A4( us13_n682 ) , .A3( us13_n683 ) , .A2( us13_n684 ) , .A1( us13_n685 ) , .ZN( us13_n690 ) );
  OR4_X1 us13_U144 (.A4( us13_n580 ) , .A3( us13_n581 ) , .A2( us13_n582 ) , .A1( us13_n583 ) , .ZN( us13_n584 ) );
  NAND2_X1 us13_U145 (.ZN( us13_n613 ) , .A2( us13_n837 ) , .A1( us13_n873 ) );
  OR3_X1 us13_U146 (.A3( us13_n506 ) , .A2( us13_n507 ) , .A1( us13_n508 ) , .ZN( us13_n511 ) );
  AOI221_X1 us13_U147 (.A( us13_n713 ) , .B2( us13_n714 ) , .ZN( us13_n720 ) , .C1( us13_n832 ) , .B1( us13_n839 ) , .C2( us13_n863 ) );
  OR2_X1 us13_U148 (.A2( us13_n711 ) , .A1( us13_n712 ) , .ZN( us13_n713 ) );
  INV_X1 us13_U149 (.A( us13_n463 ) , .ZN( us13_n864 ) );
  OR3_X1 us13_U15 (.ZN( us13_n446 ) , .A1( us13_n528 ) , .A3( us13_n577 ) , .A2( us13_n875 ) );
  OAI21_X1 us13_U150 (.ZN( us13_n463 ) , .B1( us13_n809 ) , .A( us13_n834 ) , .B2( us13_n851 ) );
  INV_X1 us13_U151 (.A( us13_n754 ) , .ZN( us13_n869 ) );
  OAI21_X1 us13_U152 (.B1( us13_n753 ) , .ZN( us13_n754 ) , .A( us13_n845 ) , .B2( us13_n868 ) );
  INV_X1 us13_U153 (.A( us13_n672 ) , .ZN( us13_n859 ) );
  AOI21_X1 us13_U154 (.A( us13_n670 ) , .B1( us13_n671 ) , .ZN( us13_n672 ) , .B2( us13_n856 ) );
  NAND2_X1 us13_U155 (.A1( us13_n447 ) , .A2( us13_n465 ) , .ZN( us13_n749 ) );
  OAI222_X1 us13_U156 (.B2( us13_n747 ) , .B1( us13_n748 ) , .A2( us13_n749 ) , .ZN( us13_n757 ) , .C2( us13_n805 ) , .C1( us13_n814 ) , .A1( us13_n817 ) );
  OAI222_X1 us13_U157 (.B2( us13_n708 ) , .ZN( us13_n709 ) , .C2( us13_n724 ) , .B1( us13_n747 ) , .A1( us13_n806 ) , .C1( us13_n814 ) , .A2( us13_n815 ) );
  OAI222_X1 us13_U158 (.ZN( us13_n505 ) , .C2( us13_n625 ) , .B2( us13_n647 ) , .B1( us13_n747 ) , .A2( us13_n748 ) , .C1( us13_n805 ) , .A1( us13_n806 ) );
  NOR4_X1 us13_U159 (.A2( us13_n491 ) , .A1( us13_n492 ) , .ZN( us13_n493 ) , .A3( us13_n580 ) , .A4( us13_n612 ) );
  OR4_X1 us13_U16 (.A4( us13_n442 ) , .A2( us13_n443 ) , .A1( us13_n444 ) , .ZN( us13_n445 ) , .A3( us13_n553 ) );
  OR4_X1 us13_U160 (.ZN( us13_n492 ) , .A4( us13_n534 ) , .A2( us13_n547 ) , .A1( us13_n559 ) , .A3( us13_n632 ) );
  OAI22_X1 us13_U161 (.B1( us13_n490 ) , .ZN( us13_n491 ) , .A1( us13_n686 ) , .A2( us13_n763 ) , .B2( us13_n817 ) );
  NOR3_X1 us13_U162 (.ZN( us13_n490 ) , .A1( us13_n782 ) , .A2( us13_n850 ) , .A3( us13_n863 ) );
  INV_X1 us13_U163 (.A( us13_n730 ) , .ZN( us13_n839 ) );
  INV_X1 us13_U164 (.A( us13_n790 ) , .ZN( us13_n832 ) );
  NAND2_X1 us13_U165 (.A1( us13_n451 ) , .A2( us13_n453 ) , .ZN( us13_n762 ) );
  AOI211_X1 us13_U166 (.A( us13_n637 ) , .ZN( us13_n645 ) , .B( us13_n743 ) , .C2( us13_n839 ) , .C1( us13_n854 ) );
  OAI22_X1 us13_U167 (.ZN( us13_n637 ) , .A1( us13_n699 ) , .B2( us13_n728 ) , .A2( us13_n762 ) , .B1( us13_n816 ) );
  OAI221_X1 us13_U168 (.A( us13_n727 ) , .C2( us13_n728 ) , .B2( us13_n729 ) , .B1( us13_n730 ) , .ZN( us13_n737 ) , .C1( us13_n817 ) );
  AOI22_X1 us13_U169 (.ZN( us13_n727 ) , .B1( us13_n832 ) , .A2( us13_n838 ) , .A1( us13_n863 ) , .B2( us13_n866 ) );
  INV_X1 us13_U17 (.A( us13_n613 ) , .ZN( us13_n875 ) );
  INV_X1 us13_U170 (.A( us13_n744 ) , .ZN( us13_n837 ) );
  OAI22_X1 us13_U171 (.ZN( us13_n489 ) , .A1( us13_n724 ) , .B2( us13_n728 ) , .B1( us13_n730 ) , .A2( us13_n779 ) );
  OAI22_X1 us13_U172 (.ZN( us13_n624 ) , .B1( us13_n669 ) , .B2( us13_n747 ) , .A1( us13_n815 ) , .A2( us13_n816 ) );
  OAI22_X1 us13_U173 (.B2( us13_n779 ) , .B1( us13_n780 ) , .ZN( us13_n781 ) , .A2( us13_n814 ) , .A1( us13_n815 ) );
  OAI22_X1 us13_U174 (.A1( us13_n724 ) , .ZN( us13_n726 ) , .B2( us13_n750 ) , .B1( us13_n812 ) , .A2( us13_n816 ) );
  INV_X1 us13_U175 (.A( us13_n805 ) , .ZN( us13_n860 ) );
  OAI22_X1 us13_U176 (.B2( us13_n744 ) , .ZN( us13_n746 ) , .A2( us13_n762 ) , .B1( us13_n780 ) , .A1( us13_n792 ) );
  OAI22_X1 us13_U177 (.B2( us13_n803 ) , .B1( us13_n804 ) , .A2( us13_n805 ) , .A1( us13_n806 ) , .ZN( us13_n808 ) );
  OAI22_X1 us13_U178 (.ZN( us13_n496 ) , .A2( us13_n744 ) , .A1( us13_n780 ) , .B1( us13_n791 ) , .B2( us13_n806 ) );
  OAI22_X1 us13_U179 (.ZN( us13_n710 ) , .A2( us13_n728 ) , .B2( us13_n729 ) , .A1( us13_n744 ) , .B1( us13_n813 ) );
  INV_X1 us13_U18 (.A( us13_n749 ) , .ZN( us13_n863 ) );
  INV_X1 us13_U180 (.A( us13_n788 ) , .ZN( us13_n845 ) );
  INV_X1 us13_U181 (.A( us13_n814 ) , .ZN( us13_n833 ) );
  OAI22_X1 us13_U182 (.ZN( us13_n590 ) , .B1( us13_n730 ) , .B2( us13_n749 ) , .A2( us13_n786 ) , .A1( us13_n803 ) );
  OAI22_X1 us13_U183 (.ZN( us13_n695 ) , .A2( us13_n730 ) , .A1( us13_n780 ) , .B1( us13_n791 ) , .B2( us13_n817 ) );
  INV_X1 us13_U184 (.A( us13_n816 ) , .ZN( us13_n831 ) );
  INV_X1 us13_U185 (.A( us13_n669 ) , .ZN( us13_n865 ) );
  NOR2_X1 us13_U186 (.ZN( us13_n715 ) , .A1( us13_n805 ) , .A2( us13_n817 ) );
  NOR2_X1 us13_U187 (.ZN( us13_n718 ) , .A2( us13_n724 ) , .A1( us13_n744 ) );
  NOR2_X1 us13_U188 (.ZN( us13_n666 ) , .A1( us13_n728 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U189 (.ZN( us13_n546 ) , .A2( us13_n780 ) , .A1( us13_n814 ) );
  AOI222_X1 us13_U19 (.ZN( us13_n563 ) , .B1( us13_n830 ) , .C1( us13_n841 ) , .A2( us13_n843 ) , .A1( us13_n854 ) , .B2( us13_n863 ) , .C2( us13_n873 ) );
  NOR2_X1 us13_U190 (.ZN( us13_n577 ) , .A2( us13_n699 ) , .A1( us13_n814 ) );
  NOR2_X1 us13_U191 (.ZN( us13_n570 ) , .A1( us13_n728 ) , .A2( us13_n806 ) );
  NOR2_X1 us13_U192 (.A2( us13_n744 ) , .ZN( us13_n755 ) , .A1( us13_n805 ) );
  INV_X1 us13_U193 (.A( us13_n750 ) , .ZN( us13_n842 ) );
  NOR2_X1 us13_U194 (.ZN( us13_n735 ) , .A2( us13_n803 ) , .A1( us13_n805 ) );
  NOR2_X1 us13_U195 (.ZN( us13_n532 ) , .A2( us13_n749 ) , .A1( us13_n750 ) );
  NOR2_X1 us13_U196 (.ZN( us13_n654 ) , .A1( us13_n728 ) , .A2( us13_n813 ) );
  OAI22_X1 us13_U197 (.ZN( us13_n483 ) , .A1( us13_n708 ) , .B2( us13_n785 ) , .A2( us13_n806 ) , .B1( us13_n812 ) );
  NOR2_X1 us13_U198 (.ZN( us13_n629 ) , .A2( us13_n728 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U199 (.ZN( us13_n615 ) , .A1( us13_n785 ) , .A2( us13_n815 ) );
  AOI222_X1 us13_U20 (.ZN( us13_n660 ) , .A2( us13_n839 ) , .B1( us13_n841 ) , .C2( us13_n845 ) , .A1( us13_n860 ) , .C1( us13_n863 ) , .B2( us13_n870 ) );
  NOR2_X1 us13_U200 (.ZN( us13_n612 ) , .A1( us13_n779 ) , .A2( us13_n786 ) );
  NOR2_X1 us13_U201 (.ZN( us13_n628 ) , .A2( us13_n669 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U202 (.ZN( us13_n611 ) , .A2( us13_n780 ) , .A1( us13_n806 ) );
  NOR2_X1 us13_U203 (.ZN( us13_n601 ) , .A2( us13_n780 ) , .A1( us13_n803 ) );
  INV_X1 us13_U204 (.A( us13_n747 ) , .ZN( us13_n834 ) );
  NOR2_X1 us13_U205 (.ZN( us13_n528 ) , .A2( us13_n724 ) , .A1( us13_n803 ) );
  NOR2_X1 us13_U206 (.ZN( us13_n531 ) , .A2( us13_n780 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U207 (.A2( us13_n708 ) , .A1( us13_n750 ) , .ZN( us13_n771 ) );
  NOR2_X1 us13_U208 (.ZN( us13_n599 ) , .A2( us13_n791 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U209 (.ZN( us13_n652 ) , .A1( us13_n669 ) , .A2( us13_n814 ) );
  INV_X1 us13_U21 (.A( us13_n647 ) , .ZN( us13_n870 ) );
  INV_X1 us13_U210 (.A( us13_n792 ) , .ZN( us13_n851 ) );
  NOR2_X1 us13_U211 (.A1( us13_n669 ) , .ZN( us13_n673 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U212 (.ZN( us13_n602 ) , .A1( us13_n669 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U213 (.A1( us13_n669 ) , .ZN( us13_n688 ) , .A2( us13_n816 ) );
  NOR2_X1 us13_U214 (.ZN( us13_n667 ) , .A1( us13_n750 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U215 (.A2( us13_n744 ) , .ZN( us13_n769 ) , .A1( us13_n812 ) );
  NOR2_X1 us13_U216 (.ZN( us13_n555 ) , .A1( us13_n750 ) , .A2( us13_n791 ) );
  NOR2_X1 us13_U217 (.ZN( us13_n508 ) , .A2( us13_n780 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U218 (.ZN( us13_n543 ) , .A2( us13_n708 ) , .A1( us13_n785 ) );
  NOR2_X1 us13_U219 (.ZN( us13_n664 ) , .A1( us13_n785 ) , .A2( us13_n791 ) );
  NOR4_X1 us13_U22 (.ZN( us13_n473 ) , .A2( us13_n521 ) , .A4( us13_n594 ) , .A1( us13_n609 ) , .A3( us13_n629 ) );
  NOR2_X1 us13_U220 (.A1( us13_n669 ) , .ZN( us13_n766 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U221 (.A1( us13_n699 ) , .ZN( us13_n768 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U222 (.ZN( us13_n527 ) , .A1( us13_n669 ) , .A2( us13_n779 ) );
  NOR2_X1 us13_U223 (.ZN( us13_n557 ) , .A1( us13_n792 ) , .A2( us13_n814 ) );
  NOR2_X1 us13_U224 (.ZN( us13_n545 ) , .A1( us13_n749 ) , .A2( us13_n814 ) );
  NOR2_X1 us13_U225 (.ZN( us13_n556 ) , .A1( us13_n762 ) , .A2( us13_n805 ) );
  NOR2_X1 us13_U226 (.ZN( us13_n661 ) , .A1( us13_n729 ) , .A2( us13_n790 ) );
  NOR2_X1 us13_U227 (.ZN( us13_n507 ) , .A1( us13_n812 ) , .A2( us13_n817 ) );
  INV_X1 us13_U228 (.A( us13_n806 ) , .ZN( us13_n841 ) );
  NOR2_X1 us13_U229 (.ZN( us13_n554 ) , .A1( us13_n786 ) , .A2( us13_n813 ) );
  NOR4_X1 us13_U23 (.A4( us13_n544 ) , .A3( us13_n545 ) , .A2( us13_n546 ) , .A1( us13_n547 ) , .ZN( us13_n548 ) );
  NOR2_X1 us13_U230 (.ZN( us13_n509 ) , .A1( us13_n729 ) , .A2( us13_n779 ) );
  NOR2_X1 us13_U231 (.ZN( us13_n530 ) , .A2( us13_n744 ) , .A1( us13_n792 ) );
  OAI22_X1 us13_U232 (.B2( us13_n750 ) , .B1( us13_n751 ) , .A1( us13_n752 ) , .ZN( us13_n756 ) , .A2( us13_n806 ) );
  NOR2_X1 us13_U233 (.ZN( us13_n751 ) , .A2( us13_n852 ) , .A1( us13_n860 ) );
  NOR3_X1 us13_U234 (.ZN( us13_n752 ) , .A2( us13_n853 ) , .A1( us13_n863 ) , .A3( us13_n865 ) );
  NOR2_X1 us13_U235 (.ZN( us13_n544 ) , .A2( us13_n785 ) , .A1( us13_n792 ) );
  NOR2_X1 us13_U236 (.A1( us13_n749 ) , .ZN( us13_n767 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U237 (.ZN( us13_n516 ) , .A1( us13_n708 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U238 (.ZN( us13_n663 ) , .A1( us13_n729 ) , .A2( us13_n785 ) );
  OAI22_X1 us13_U239 (.B1( us13_n440 ) , .ZN( us13_n444 ) , .A2( us13_n728 ) , .A1( us13_n744 ) , .B2( us13_n749 ) );
  NOR4_X1 us13_U24 (.ZN( us13_n479 ) , .A1( us13_n520 ) , .A4( us13_n557 ) , .A3( us13_n582 ) , .A2( us13_n630 ) );
  NOR3_X1 us13_U240 (.ZN( us13_n440 ) , .A2( us13_n836 ) , .A3( us13_n837 ) , .A1( us13_n846 ) );
  NOR2_X1 us13_U241 (.ZN( us13_n717 ) , .A2( us13_n744 ) , .A1( us13_n786 ) );
  NOR2_X1 us13_U243 (.ZN( us13_n506 ) , .A2( us13_n728 ) , .A1( us13_n762 ) );
  NOR2_X1 us13_U244 (.ZN( us13_n614 ) , .A1( us13_n762 ) , .A2( us13_n812 ) );
  NOR2_X1 us13_U245 (.ZN( us13_n517 ) , .A1( us13_n708 ) , .A2( us13_n803 ) );
  NOR2_X1 us13_U246 (.ZN( us13_n558 ) , .A1( us13_n708 ) , .A2( us13_n816 ) );
  AOI21_X1 us13_U247 (.A( us13_n812 ) , .B2( us13_n813 ) , .B1( us13_n814 ) , .ZN( us13_n819 ) );
  NOR2_X1 us13_U248 (.ZN( us13_n670 ) , .A1( us13_n790 ) , .A2( us13_n805 ) );
  NOR2_X1 us13_U249 (.ZN( us13_n630 ) , .A1( us13_n747 ) , .A2( us13_n815 ) );
  NOR4_X1 us13_U25 (.ZN( us13_n456 ) , .A2( us13_n517 ) , .A1( us13_n543 ) , .A3( us13_n579 ) , .A4( us13_n615 ) );
  NOR2_X1 us13_U250 (.ZN( us13_n655 ) , .A1( us13_n790 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U251 (.ZN( us13_n521 ) , .A1( us13_n790 ) , .A2( us13_n812 ) );
  NOR2_X1 us13_U252 (.ZN( us13_n668 ) , .A2( us13_n708 ) , .A1( us13_n790 ) );
  NOR2_X1 us13_U253 (.ZN( us13_n542 ) , .A1( us13_n762 ) , .A2( us13_n791 ) );
  NOR2_X1 us13_U254 (.ZN( us13_n701 ) , .A2( us13_n786 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U255 (.ZN( us13_n631 ) , .A1( us13_n724 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U256 (.ZN( us13_n656 ) , .A1( us13_n747 ) , .A2( us13_n780 ) );
  INV_X1 us13_U257 (.A( us13_n763 ) , .ZN( us13_n866 ) );
  NOR2_X1 us13_U258 (.ZN( us13_n609 ) , .A2( us13_n724 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U259 (.A1( us13_n730 ) , .ZN( us13_n765 ) , .A2( us13_n786 ) );
  NOR4_X1 us13_U26 (.ZN( us13_n485 ) , .A2( us13_n533 ) , .A1( us13_n558 ) , .A3( us13_n631 ) , .A4( us13_n718 ) );
  NOR2_X1 us13_U260 (.ZN( us13_n533 ) , .A2( us13_n724 ) , .A1( us13_n730 ) );
  NOR2_X1 us13_U261 (.ZN( us13_n579 ) , .A2( us13_n708 ) , .A1( us13_n730 ) );
  AOI21_X1 us13_U262 (.B1( us13_n625 ) , .ZN( us13_n627 ) , .A( us13_n763 ) , .B2( us13_n814 ) );
  AOI21_X1 us13_U263 (.A( us13_n815 ) , .B2( us13_n816 ) , .B1( us13_n817 ) , .ZN( us13_n818 ) );
  NOR2_X1 us13_U264 (.ZN( us13_n582 ) , .A1( us13_n744 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U265 (.A2( us13_n708 ) , .A1( us13_n762 ) , .ZN( us13_n794 ) );
  AOI21_X1 us13_U266 (.ZN( us13_n515 ) , .A( us13_n729 ) , .B1( us13_n750 ) , .B2( us13_n803 ) );
  NOR2_X1 us13_U267 (.ZN( us13_n642 ) , .A2( us13_n788 ) , .A1( us13_n791 ) );
  AOI21_X1 us13_U268 (.ZN( us13_n499 ) , .B1( us13_n680 ) , .A( us13_n812 ) , .B2( us13_n816 ) );
  AOI21_X1 us13_U269 (.ZN( us13_n650 ) , .A( us13_n779 ) , .B1( us13_n792 ) , .B2( us13_n805 ) );
  NOR4_X1 us13_U27 (.A1( us13_n531 ) , .ZN( us13_n536 ) , .A2( us13_n654 ) , .A4( us13_n668 ) , .A3( us13_n765 ) );
  NOR2_X1 us13_U270 (.ZN( us13_n520 ) , .A2( us13_n708 ) , .A1( us13_n814 ) );
  AOI21_X1 us13_U271 (.ZN( us13_n626 ) , .B2( us13_n669 ) , .A( us13_n790 ) , .B1( us13_n791 ) );
  NOR2_X1 us13_U272 (.ZN( us13_n653 ) , .A1( us13_n762 ) , .A2( us13_n786 ) );
  AOI21_X1 us13_U273 (.ZN( us13_n477 ) , .A( us13_n669 ) , .B1( us13_n750 ) , .B2( us13_n806 ) );
  NOR2_X1 us13_U274 (.ZN( us13_n559 ) , .A2( us13_n791 ) , .A1( us13_n803 ) );
  NOR2_X1 us13_U275 (.ZN( us13_n519 ) , .A2( us13_n699 ) , .A1( us13_n816 ) );
  NOR2_X1 us13_U276 (.ZN( us13_n683 ) , .A2( us13_n699 ) , .A1( us13_n803 ) );
  AOI21_X1 us13_U277 (.ZN( us13_n510 ) , .B2( us13_n669 ) , .A( us13_n730 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U278 (.ZN( us13_n540 ) , .A( us13_n763 ) , .B2( us13_n779 ) , .B1( us13_n817 ) );
  NOR2_X1 us13_U279 (.ZN( us13_n581 ) , .A1( us13_n669 ) , .A2( us13_n788 ) );
  NOR2_X1 us13_U28 (.ZN( us13_n680 ) , .A2( us13_n834 ) , .A1( us13_n839 ) );
  AOI21_X1 us13_U280 (.ZN( us13_n589 ) , .B2( us13_n699 ) , .B1( us13_n815 ) , .A( us13_n817 ) );
  AOI21_X1 us13_U281 (.ZN( us13_n498 ) , .A( us13_n724 ) , .B2( us13_n762 ) , .B1( us13_n814 ) );
  AOI21_X1 us13_U282 (.ZN( us13_n539 ) , .B2( us13_n812 ) , .A( us13_n814 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U283 (.B1( us13_n699 ) , .ZN( us13_n700 ) , .A( us13_n732 ) , .B2( us13_n763 ) );
  AOI21_X1 us13_U284 (.ZN( us13_n591 ) , .B2( us13_n763 ) , .A( us13_n785 ) , .B1( us13_n812 ) );
  INV_X1 us13_U285 (.A( us13_n791 ) , .ZN( us13_n873 ) );
  NOR2_X1 us13_U286 (.ZN( us13_n547 ) , .A1( us13_n699 ) , .A2( us13_n744 ) );
  NOR2_X1 us13_U287 (.ZN( us13_n665 ) , .A1( us13_n780 ) , .A2( us13_n813 ) );
  INV_X1 us13_U288 (.A( us13_n729 ) , .ZN( us13_n868 ) );
  AOI21_X1 us13_U289 (.ZN( us13_n640 ) , .B2( us13_n747 ) , .A( us13_n792 ) , .B1( us13_n803 ) );
  AOI221_X1 us13_U29 (.A( us13_n781 ) , .ZN( us13_n798 ) , .C2( us13_n837 ) , .B2( us13_n838 ) , .B1( us13_n865 ) , .C1( us13_n866 ) );
  AOI21_X1 us13_U290 (.ZN( us13_n569 ) , .B1( us13_n750 ) , .B2( us13_n762 ) , .A( us13_n780 ) );
  AOI21_X1 us13_U291 (.ZN( us13_n649 ) , .B1( us13_n729 ) , .B2( us13_n763 ) , .A( us13_n813 ) );
  NOR2_X1 us13_U292 (.ZN( us13_n685 ) , .A1( us13_n729 ) , .A2( us13_n816 ) );
  AOI21_X1 us13_U293 (.B1( us13_n686 ) , .ZN( us13_n687 ) , .A( us13_n728 ) , .B2( us13_n761 ) );
  NOR2_X1 us13_U294 (.ZN( us13_n568 ) , .A1( us13_n729 ) , .A2( us13_n762 ) );
  NOR2_X1 us13_U295 (.ZN( us13_n684 ) , .A1( us13_n791 ) , .A2( us13_n813 ) );
  AOI21_X1 us13_U296 (.ZN( us13_n514 ) , .A( us13_n779 ) , .B2( us13_n792 ) , .B1( us13_n812 ) );
  AOI21_X1 us13_U297 (.ZN( us13_n593 ) , .B1( us13_n750 ) , .A( us13_n792 ) , .B2( us13_n813 ) );
  AOI21_X1 us13_U298 (.ZN( us13_n450 ) , .B2( us13_n792 ) , .A( us13_n803 ) , .B1( us13_n815 ) );
  AOI21_X1 us13_U299 (.ZN( us13_n639 ) , .B2( us13_n749 ) , .A( us13_n788 ) , .B1( us13_n812 ) );
  NAND4_X1 us13_U3 (.ZN( sa12_sr_2 ) , .A4( us13_n643 ) , .A3( us13_n644 ) , .A2( us13_n645 ) , .A1( us13_n646 ) );
  NOR4_X1 us13_U30 (.A4( us13_n793 ) , .A3( us13_n794 ) , .A2( us13_n795 ) , .A1( us13_n796 ) , .ZN( us13_n797 ) );
  INV_X1 us13_U300 (.A( us13_n699 ) , .ZN( us13_n853 ) );
  AOI21_X1 us13_U301 (.ZN( us13_n564 ) , .B1( us13_n724 ) , .A( us13_n779 ) , .B2( us13_n791 ) );
  AOI21_X1 us13_U302 (.ZN( us13_n497 ) , .A( us13_n779 ) , .B2( us13_n791 ) , .B1( us13_n804 ) );
  NOR2_X1 us13_U303 (.ZN( us13_n529 ) , .A1( us13_n708 ) , .A2( us13_n779 ) );
  AOI21_X1 us13_U304 (.ZN( us13_n689 ) , .B2( us13_n749 ) , .B1( us13_n763 ) , .A( us13_n806 ) );
  NOR2_X1 us13_U305 (.ZN( us13_n567 ) , .A1( us13_n747 ) , .A2( us13_n805 ) );
  AOI21_X1 us13_U306 (.A( us13_n790 ) , .B2( us13_n791 ) , .B1( us13_n792 ) , .ZN( us13_n793 ) );
  AOI21_X1 us13_U307 (.A( us13_n733 ) , .ZN( us13_n734 ) , .B2( us13_n780 ) , .B1( us13_n792 ) );
  NOR2_X1 us13_U308 (.A2( us13_n813 ) , .A1( us13_n815 ) , .ZN( us13_n821 ) );
  AOI21_X1 us13_U309 (.ZN( us13_n641 ) , .B1( us13_n680 ) , .A( us13_n791 ) , .B2( us13_n817 ) );
  NOR4_X1 us13_U31 (.A4( us13_n776 ) , .A3( us13_n777 ) , .A1( us13_n778 ) , .ZN( us13_n799 ) , .A2( us13_n801 ) );
  NOR2_X1 us13_U310 (.ZN( us13_n578 ) , .A1( us13_n708 ) , .A2( us13_n813 ) );
  NOR2_X1 us13_U311 (.ZN( us13_n682 ) , .A2( us13_n708 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U312 (.ZN( us13_n711 ) , .A1( us13_n762 ) , .A2( us13_n763 ) );
  NOR2_X1 us13_U313 (.ZN( us13_n583 ) , .A1( us13_n792 ) , .A2( us13_n817 ) );
  NOR2_X1 us13_U314 (.ZN( us13_n534 ) , .A1( us13_n724 ) , .A2( us13_n788 ) );
  NAND2_X1 us13_U315 (.ZN( us13_n753 ) , .A1( us13_n763 ) , .A2( us13_n805 ) );
  INV_X1 us13_U316 (.A( us13_n815 ) , .ZN( us13_n855 ) );
  AOI21_X1 us13_U317 (.ZN( us13_n442 ) , .A( us13_n699 ) , .B1( us13_n733 ) , .B2( us13_n750 ) );
  OAI21_X1 us13_U318 (.A( us13_n731 ) , .B1( us13_n732 ) , .ZN( us13_n736 ) , .B2( us13_n805 ) );
  OAI21_X1 us13_U319 (.ZN( us13_n731 ) , .A( us13_n833 ) , .B2( us13_n852 ) , .B1( us13_n873 ) );
  NOR4_X1 us13_U32 (.A3( us13_n755 ) , .A2( us13_n756 ) , .A1( us13_n757 ) , .ZN( us13_n758 ) , .A4( us13_n869 ) );
  INV_X1 us13_U320 (.A( us13_n780 ) , .ZN( us13_n850 ) );
  INV_X1 us13_U321 (.A( us13_n785 ) , .ZN( us13_n846 ) );
  AOI22_X1 us13_U322 (.ZN( us13_n696 ) , .A1( us13_n830 ) , .B2( us13_n843 ) , .A2( us13_n865 ) , .B1( us13_n868 ) );
  AOI22_X1 us13_U323 (.A2( us13_n782 ) , .ZN( us13_n783 ) , .B2( us13_n831 ) , .A1( us13_n834 ) , .B1( us13_n863 ) );
  AOI21_X1 us13_U324 (.ZN( us13_n443 ) , .B1( us13_n789 ) , .B2( us13_n791 ) , .A( us13_n814 ) );
  NAND2_X1 us13_U325 (.ZN( us13_n714 ) , .A1( us13_n728 ) , .A2( us13_n780 ) );
  OAI21_X1 us13_U326 (.A( us13_n787 ) , .B2( us13_n788 ) , .B1( us13_n789 ) , .ZN( us13_n795 ) );
  OAI21_X1 us13_U327 (.ZN( us13_n787 ) , .A( us13_n839 ) , .B1( us13_n863 ) , .B2( us13_n873 ) );
  NAND2_X1 us13_U328 (.A2( us13_n762 ) , .A1( us13_n806 ) , .ZN( us13_n810 ) );
  NOR2_X1 us13_U329 (.ZN( us13_n484 ) , .A1( us13_n788 ) , .A2( us13_n805 ) );
  AOI211_X1 us13_U33 (.B( us13_n745 ) , .A( us13_n746 ) , .ZN( us13_n759 ) , .C1( us13_n832 ) , .C2( us13_n853 ) );
  NOR2_X1 us13_U330 (.ZN( us13_n470 ) , .A2( us13_n779 ) , .A1( us13_n815 ) );
  NOR2_X1 us13_U331 (.ZN( us13_n712 ) , .A2( us13_n724 ) , .A1( us13_n790 ) );
  NOR2_X1 us13_U332 (.ZN( us13_n526 ) , .A1( us13_n724 ) , .A2( us13_n750 ) );
  NAND2_X1 us13_U333 (.A1( us13_n699 ) , .A2( us13_n729 ) , .ZN( us13_n782 ) );
  NOR2_X1 us13_U334 (.ZN( us13_n518 ) , .A1( us13_n708 ) , .A2( us13_n788 ) );
  INV_X1 us13_U335 (.A( us13_n813 ) , .ZN( us13_n836 ) );
  NAND2_X1 us13_U336 (.ZN( us13_n671 ) , .A1( us13_n806 ) , .A2( us13_n816 ) );
  OAI21_X1 us13_U337 (.A( us13_n698 ) , .ZN( us13_n702 ) , .B2( us13_n750 ) , .B1( us13_n804 ) );
  OAI21_X1 us13_U338 (.ZN( us13_n698 ) , .B2( us13_n833 ) , .B1( us13_n838 ) , .A( us13_n860 ) );
  NAND2_X1 us13_U339 (.A2( us13_n749 ) , .A1( us13_n786 ) , .ZN( us13_n809 ) );
  NOR3_X1 us13_U34 (.A3( us13_n741 ) , .A2( us13_n742 ) , .A1( us13_n743 ) , .ZN( us13_n760 ) );
  INV_X1 us13_U340 (.A( us13_n724 ) , .ZN( us13_n856 ) );
  INV_X1 us13_U341 (.A( us13_n817 ) , .ZN( us13_n844 ) );
  NAND2_X2 us13_U342 (.A1( us13_n451 ) , .A2( us13_n462 ) , .ZN( us13_n790 ) );
  AND2_X1 us13_U343 (.ZN( us13_n732 ) , .A1( us13_n779 ) , .A2( us13_n785 ) );
  OAI222_X1 us13_U344 (.ZN( us13_n617 ) , .B1( us13_n697 ) , .C1( us13_n724 ) , .C2( us13_n747 ) , .B2( us13_n786 ) , .A2( us13_n792 ) , .A1( us13_n816 ) );
  AOI221_X1 us13_U345 (.A( us13_n764 ) , .ZN( us13_n774 ) , .C2( us13_n810 ) , .B2( us13_n835 ) , .C1( us13_n855 ) , .B1( us13_n866 ) );
  AOI21_X1 us13_U346 (.B2( us13_n763 ) , .ZN( us13_n764 ) , .A( us13_n788 ) , .B1( us13_n792 ) );
  INV_X1 us13_U347 (.A( us13_n761 ) , .ZN( us13_n835 ) );
  NAND2_X1 us13_U348 (.A1( us13_n451 ) , .A2( us13_n454 ) , .ZN( us13_n814 ) );
  NAND2_X1 us13_U349 (.A1( us13_n447 ) , .A2( us13_n449 ) , .ZN( us13_n805 ) );
  NOR4_X1 us13_U35 (.A4( us13_n734 ) , .A3( us13_n735 ) , .A2( us13_n736 ) , .A1( us13_n737 ) , .ZN( us13_n738 ) );
  NAND2_X1 us13_U350 (.A1( us13_n453 ) , .A2( us13_n461 ) , .ZN( us13_n744 ) );
  NAND2_X1 us13_U351 (.A1( us13_n455 ) , .A2( us13_n471 ) , .ZN( us13_n803 ) );
  NAND2_X1 us13_U352 (.A1( us13_n455 ) , .A2( us13_n462 ) , .ZN( us13_n750 ) );
  NAND2_X1 us13_U353 (.A1( us13_n451 ) , .A2( us13_n471 ) , .ZN( us13_n816 ) );
  NAND2_X1 us13_U356 (.A2( us13_n453 ) , .A1( us13_n455 ) , .ZN( us13_n806 ) );
  NAND2_X1 us13_U357 (.A1( us13_n453 ) , .A2( us13_n472 ) , .ZN( us13_n785 ) );
  NAND2_X1 us13_U358 (.A2( us13_n454 ) , .A1( us13_n472 ) , .ZN( us13_n779 ) );
  NAND2_X1 us13_U359 (.A2( us13_n464 ) , .A1( us13_n465 ) , .ZN( us13_n812 ) );
  AOI211_X1 us13_U36 (.B( us13_n725 ) , .A( us13_n726 ) , .ZN( us13_n739 ) , .C1( us13_n843 ) , .C2( us13_n855 ) );
  NAND2_X1 us13_U360 (.A1( us13_n441 ) , .A2( us13_n460 ) , .ZN( us13_n699 ) );
  NAND2_X1 us13_U361 (.A2( us13_n449 ) , .A1( us13_n452 ) , .ZN( us13_n763 ) );
  NAND2_X1 us13_U362 (.A2( us13_n448 ) , .A1( us13_n452 ) , .ZN( us13_n729 ) );
  NAND2_X1 us13_U363 (.A1( us13_n447 ) , .A2( us13_n448 ) , .ZN( us13_n786 ) );
  NAND2_X1 us13_U364 (.A2( us13_n461 ) , .A1( us13_n462 ) , .ZN( us13_n747 ) );
  NAND2_X1 us13_U365 (.A1( us13_n462 ) , .A2( us13_n472 ) , .ZN( us13_n788 ) );
  NOR2_X1 us13_U367 (.ZN( us13_n453 ) , .A1( us13_n826 ) , .A2( us13_n827 ) );
  NOR2_X1 us13_U368 (.ZN( us13_n451 ) , .A1( us13_n828 ) , .A2( us13_n829 ) );
  NAND2_X1 us13_U369 (.A2( us13_n461 ) , .A1( us13_n471 ) , .ZN( us13_n697 ) );
  NOR3_X1 us13_U37 (.A3( us13_n722 ) , .A1( us13_n723 ) , .ZN( us13_n740 ) , .A2( us13_n741 ) );
  NAND2_X1 us13_U370 (.A2( us13_n454 ) , .A1( us13_n455 ) , .ZN( us13_n730 ) );
  NAND2_X1 us13_U371 (.A2( us13_n441 ) , .A1( us13_n447 ) , .ZN( us13_n784 ) );
  NAND2_X2 us13_U372 (.A2( us13_n448 ) , .A1( us13_n464 ) , .ZN( us13_n815 ) );
  NAND2_X2 us13_U373 (.A2( us13_n441 ) , .A1( us13_n452 ) , .ZN( us13_n791 ) );
  NAND2_X2 us13_U374 (.A1( us13_n449 ) , .A2( us13_n460 ) , .ZN( us13_n792 ) );
  NAND2_X2 us13_U375 (.A1( us13_n441 ) , .A2( us13_n464 ) , .ZN( us13_n708 ) );
  NAND2_X2 us13_U376 (.A2( us13_n460 ) , .A1( us13_n465 ) , .ZN( us13_n780 ) );
  NOR2_X1 us13_U378 (.A2( sa13_6 ) , .A1( sa13_7 ) , .ZN( us13_n464 ) );
  NAND4_X1 us13_U38 (.ZN( sa12_sr_3 ) , .A4( us13_n704 ) , .A3( us13_n705 ) , .A2( us13_n706 ) , .A1( us13_n707 ) );
  NOR2_X1 us13_U381 (.A2( sa13_4 ) , .A1( sa13_5 ) , .ZN( us13_n441 ) );
  NOR2_X1 us13_U383 (.A2( sa13_1 ) , .ZN( us13_n471 ) , .A1( us13_n826 ) );
  NOR2_X1 us13_U384 (.A2( sa13_2 ) , .A1( sa13_3 ) , .ZN( us13_n472 ) );
  NOR2_X1 us13_U386 (.A2( sa13_0 ) , .A1( sa13_1 ) , .ZN( us13_n462 ) );
  NOR2_X1 us13_U387 (.A2( sa13_3 ) , .ZN( us13_n455 ) , .A1( us13_n828 ) );
  NOR2_X1 us13_U388 (.A2( sa13_2 ) , .ZN( us13_n461 ) , .A1( us13_n829 ) );
  NOR2_X1 us13_U389 (.A2( sa13_0 ) , .ZN( us13_n454 ) , .A1( us13_n827 ) );
  NOR4_X1 us13_U39 (.A4( us13_n700 ) , .A3( us13_n701 ) , .A2( us13_n702 ) , .A1( us13_n703 ) , .ZN( us13_n704 ) );
  INV_X1 us13_U392 (.A( sa13_1 ) , .ZN( us13_n827 ) );
  INV_X1 us13_U393 (.A( sa13_3 ) , .ZN( us13_n829 ) );
  INV_X1 us13_U394 (.A( sa13_0 ) , .ZN( us13_n826 ) );
  INV_X1 us13_U395 (.A( sa13_2 ) , .ZN( us13_n828 ) );
  AOI21_X1 us13_U398 (.ZN( us13_n500 ) , .A( us13_n697 ) , .B1( us13_n708 ) , .B2( us13_n786 ) );
  INV_X1 us13_U399 (.A( us13_n697 ) , .ZN( us13_n838 ) );
  NAND2_X1 us13_U4 (.A1( us13_n449 ) , .A2( us13_n464 ) , .ZN( us13_n724 ) );
  AOI211_X1 us13_U40 (.B( us13_n694 ) , .A( us13_n695 ) , .ZN( us13_n705 ) , .C2( us13_n831 ) , .C1( us13_n851 ) );
  AOI21_X1 us13_U400 (.ZN( us13_n571 ) , .B2( us13_n697 ) , .B1( us13_n806 ) , .A( us13_n812 ) );
  NOR2_X1 us13_U401 (.A1( us13_n697 ) , .ZN( us13_n770 ) , .A2( us13_n815 ) );
  NOR2_X1 us13_U402 (.ZN( us13_n566 ) , .A2( us13_n697 ) , .A1( us13_n763 ) );
  AOI21_X1 us13_U403 (.ZN( us13_n552 ) , .B1( us13_n669 ) , .A( us13_n697 ) , .B2( us13_n805 ) );
  NOR2_X1 us13_U404 (.ZN( us13_n632 ) , .A2( us13_n697 ) , .A1( us13_n724 ) );
  NOR2_X1 us13_U405 (.ZN( us13_n541 ) , .A2( us13_n697 ) , .A1( us13_n699 ) );
  AOI21_X1 us13_U406 (.ZN( us13_n478 ) , .B2( us13_n697 ) , .A( us13_n749 ) , .B1( us13_n779 ) );
  NOR2_X1 us13_U407 (.A2( us13_n697 ) , .A1( us13_n780 ) , .ZN( us13_n820 ) );
  NOR2_X1 us13_U408 (.ZN( us13_n662 ) , .A2( us13_n697 ) , .A1( us13_n729 ) );
  NOR2_X1 us13_U409 (.A2( us13_n697 ) , .ZN( us13_n716 ) , .A1( us13_n792 ) );
  NOR2_X1 us13_U41 (.ZN( us13_n707 ) , .A2( us13_n776 ) , .A1( us13_n800 ) );
  NOR2_X1 us13_U410 (.ZN( us13_n594 ) , .A2( us13_n697 ) , .A1( us13_n728 ) );
  NOR2_X1 us13_U411 (.ZN( us13_n580 ) , .A2( us13_n697 ) , .A1( us13_n791 ) );
  OAI221_X1 us13_U412 (.A( us13_n783 ) , .C2( us13_n784 ) , .B2( us13_n785 ) , .B1( us13_n786 ) , .ZN( us13_n796 ) , .C1( us13_n813 ) );
  OAI22_X1 us13_U413 (.ZN( us13_n588 ) , .A2( us13_n747 ) , .B2( us13_n762 ) , .A1( us13_n763 ) , .B1( us13_n784 ) );
  AOI21_X1 us13_U414 (.ZN( us13_n592 ) , .B1( us13_n728 ) , .B2( us13_n784 ) , .A( us13_n790 ) );
  OAI221_X1 us13_U415 (.A( us13_n696 ) , .ZN( us13_n703 ) , .C2( us13_n784 ) , .C1( us13_n785 ) , .B1( us13_n786 ) , .B2( us13_n806 ) );
  NAND2_X1 us13_U416 (.A1( us13_n729 ) , .A2( us13_n784 ) , .ZN( us13_n811 ) );
  AOI21_X1 us13_U417 (.ZN( us13_n623 ) , .B1( us13_n699 ) , .A( us13_n779 ) , .B2( us13_n784 ) );
  AOI21_X1 us13_U418 (.ZN( us13_n648 ) , .A( us13_n762 ) , .B2( us13_n784 ) , .B1( us13_n792 ) );
  OAI22_X1 us13_U419 (.ZN( us13_n681 ) , .A1( us13_n699 ) , .A2( us13_n730 ) , .B2( us13_n784 ) , .B1( us13_n817 ) );
  NOR2_X1 us13_U42 (.ZN( us13_n804 ) , .A1( us13_n854 ) , .A2( us13_n861 ) );
  NOR2_X1 us13_U420 (.ZN( us13_n651 ) , .A1( us13_n784 ) , .A2( us13_n788 ) );
  NOR2_X1 us13_U421 (.ZN( us13_n553 ) , .A2( us13_n744 ) , .A1( us13_n784 ) );
  OAI21_X1 us13_U422 (.A( us13_n613 ) , .ZN( us13_n616 ) , .B1( us13_n625 ) , .B2( us13_n784 ) );
  NOR2_X1 us13_U423 (.ZN( us13_n610 ) , .A1( us13_n784 ) , .A2( us13_n816 ) );
  OAI222_X1 us13_U424 (.A2( us13_n669 ) , .ZN( us13_n674 ) , .B1( us13_n747 ) , .B2( us13_n784 ) , .C2( us13_n788 ) , .C1( us13_n815 ) , .A1( us13_n817 ) );
  NOR2_X1 us13_U425 (.ZN( us13_n600 ) , .A2( us13_n697 ) , .A1( us13_n784 ) );
  INV_X1 us13_U426 (.A( us13_n784 ) , .ZN( us13_n861 ) );
  NAND2_X1 us13_U427 (.A1( us13_n454 ) , .A2( us13_n461 ) , .ZN( us13_n813 ) );
  NOR2_X1 us13_U428 (.ZN( us13_n789 ) , .A2( us13_n862 ) , .A1( us13_n868 ) );
  AOI221_X1 us13_U429 (.A( us13_n483 ) , .ZN( us13_n488 ) , .B1( us13_n831 ) , .C2( us13_n844 ) , .C1( us13_n852 ) , .B2( us13_n862 ) );
  AOI222_X1 us13_U43 (.B2( us13_n638 ) , .ZN( us13_n644 ) , .B1( us13_n841 ) , .A1( us13_n842 ) , .C2( us13_n846 ) , .C1( us13_n863 ) , .A2( us13_n865 ) );
  AOI221_X1 us13_U430 (.A( us13_n681 ) , .ZN( us13_n692 ) , .B2( us13_n840 ) , .C1( us13_n842 ) , .C2( us13_n862 ) , .B1( us13_n865 ) );
  AOI222_X1 us13_U431 (.ZN( us13_n605 ) , .B2( us13_n671 ) , .B1( us13_n753 ) , .C2( us13_n831 ) , .A1( us13_n833 ) , .A2( us13_n862 ) , .C1( us13_n863 ) );
  INV_X1 us13_U432 (.A( us13_n786 ) , .ZN( us13_n862 ) );
  AND2_X1 us13_U433 (.ZN( us13_n438 ) , .A2( us13_n831 ) , .A1( us13_n854 ) );
  AND2_X1 us13_U434 (.ZN( us13_n439 ) , .A2( us13_n843 ) , .A1( us13_n861 ) );
  NOR3_X1 us13_U435 (.A1( us13_n438 ) , .A2( us13_n439 ) , .A3( us13_n576 ) , .ZN( us13_n587 ) );
  INV_X1 us13_U436 (.A( us13_n812 ) , .ZN( us13_n854 ) );
  NAND3_X1 us13_U437 (.ZN( sa12_sr_6 ) , .A3( us13_n797 ) , .A2( us13_n798 ) , .A1( us13_n799 ) );
  NAND3_X1 us13_U438 (.ZN( sa12_sr_5 ) , .A3( us13_n758 ) , .A2( us13_n759 ) , .A1( us13_n760 ) );
  NAND3_X1 us13_U439 (.ZN( sa12_sr_4 ) , .A3( us13_n738 ) , .A2( us13_n739 ) , .A1( us13_n740 ) );
  NOR4_X1 us13_U44 (.A4( us13_n639 ) , .A3( us13_n640 ) , .A2( us13_n641 ) , .A1( us13_n642 ) , .ZN( us13_n643 ) );
  NAND3_X1 us13_U440 (.A3( us13_n675 ) , .A2( us13_n676 ) , .A1( us13_n677 ) , .ZN( us13_n807 ) );
  NAND3_X1 us13_U441 (.ZN( us13_n638 ) , .A3( us13_n708 ) , .A2( us13_n724 ) , .A1( us13_n792 ) );
  NAND3_X1 us13_U442 (.A3( us13_n618 ) , .A2( us13_n619 ) , .A1( us13_n620 ) , .ZN( us13_n725 ) );
  NAND3_X1 us13_U443 (.A3( us13_n585 ) , .A2( us13_n586 ) , .A1( us13_n587 ) , .ZN( us13_n621 ) );
  NAND3_X1 us13_U444 (.ZN( us13_n565 ) , .A3( us13_n680 ) , .A2( us13_n750 ) , .A1( us13_n785 ) );
  NAND3_X1 us13_U445 (.A3( us13_n523 ) , .A2( us13_n524 ) , .A1( us13_n525 ) , .ZN( us13_n742 ) );
  NAND3_X1 us13_U446 (.A3( us13_n512 ) , .A1( us13_n513 ) , .ZN( us13_n608 ) , .A2( us13_n871 ) );
  NAND3_X1 us13_U447 (.A3( us13_n467 ) , .A2( us13_n468 ) , .A1( us13_n469 ) , .ZN( us13_n777 ) );
  INV_X1 us13_U448 (.A( us13_n803 ) , .ZN( us13_n843 ) );
  AOI21_X1 us13_U449 (.ZN( us13_n576 ) , .B2( us13_n724 ) , .B1( us13_n748 ) , .A( us13_n785 ) );
  NOR3_X1 us13_U45 (.A2( us13_n607 ) , .A1( us13_n608 ) , .ZN( us13_n646 ) , .A3( us13_n722 ) );
  NAND4_X1 us13_U46 (.ZN( sa12_sr_0 ) , .A4( us13_n501 ) , .A3( us13_n502 ) , .A2( us13_n503 ) , .A1( us13_n504 ) );
  AOI221_X1 us13_U47 (.A( us13_n497 ) , .ZN( us13_n502 ) , .B2( us13_n843 ) , .C1( us13_n846 ) , .C2( us13_n860 ) , .B1( us13_n862 ) );
  NOR4_X1 us13_U48 (.A4( us13_n498 ) , .A3( us13_n499 ) , .A2( us13_n500 ) , .ZN( us13_n501 ) , .A1( us13_n527 ) );
  AOI211_X1 us13_U49 (.A( us13_n496 ) , .ZN( us13_n503 ) , .B( us13_n802 ) , .C2( us13_n839 ) , .C1( us13_n851 ) );
  NAND2_X1 us13_U5 (.A2( us13_n471 ) , .A1( us13_n472 ) , .ZN( us13_n817 ) );
  NAND4_X1 us13_U50 (.ZN( sa12_sr_1 ) , .A4( us13_n595 ) , .A3( us13_n596 ) , .A2( us13_n597 ) , .A1( us13_n598 ) );
  AOI211_X1 us13_U51 (.B( us13_n589 ) , .A( us13_n590 ) , .ZN( us13_n596 ) , .C2( us13_n811 ) , .C1( us13_n833 ) );
  NOR4_X1 us13_U52 (.A4( us13_n591 ) , .A3( us13_n592 ) , .A2( us13_n593 ) , .A1( us13_n594 ) , .ZN( us13_n595 ) );
  AOI211_X1 us13_U53 (.A( us13_n588 ) , .ZN( us13_n597 ) , .B( us13_n621 ) , .C1( us13_n845 ) , .C2( us13_n855 ) );
  NOR2_X1 us13_U54 (.ZN( us13_n748 ) , .A1( us13_n861 ) , .A2( us13_n862 ) );
  NAND4_X1 us13_U55 (.ZN( sa12_sr_7 ) , .A4( us13_n822 ) , .A3( us13_n823 ) , .A2( us13_n824 ) , .A1( us13_n825 ) );
  AOI222_X1 us13_U56 (.C2( us13_n809 ) , .B2( us13_n810 ) , .A2( us13_n811 ) , .ZN( us13_n823 ) , .C1( us13_n832 ) , .A1( us13_n839 ) , .B1( us13_n853 ) );
  NOR4_X1 us13_U57 (.A4( us13_n818 ) , .A3( us13_n819 ) , .A2( us13_n820 ) , .A1( us13_n821 ) , .ZN( us13_n822 ) );
  AOI211_X1 us13_U58 (.B( us13_n807 ) , .A( us13_n808 ) , .ZN( us13_n824 ) , .C1( us13_n842 ) , .C2( us13_n850 ) );
  NOR2_X1 us13_U59 (.ZN( us13_n625 ) , .A2( us13_n836 ) , .A1( us13_n839 ) );
  NOR3_X1 us13_U6 (.ZN( us13_n598 ) , .A1( us13_n608 ) , .A3( us13_n723 ) , .A2( us13_n742 ) );
  NAND4_X1 us13_U60 (.A4( us13_n603 ) , .A3( us13_n604 ) , .A2( us13_n605 ) , .A1( us13_n606 ) , .ZN( us13_n722 ) );
  NOR3_X1 us13_U61 (.A1( us13_n599 ) , .ZN( us13_n604 ) , .A3( us13_n663 ) , .A2( us13_n770 ) );
  NOR4_X1 us13_U62 (.A3( us13_n600 ) , .A2( us13_n601 ) , .A1( us13_n602 ) , .ZN( us13_n603 ) , .A4( us13_n655 ) );
  AOI222_X1 us13_U63 (.ZN( us13_n606 ) , .A1( us13_n830 ) , .C2( us13_n837 ) , .B1( us13_n842 ) , .A2( us13_n856 ) , .B2( us13_n861 ) , .C1( us13_n868 ) );
  AOI222_X1 us13_U64 (.ZN( us13_n469 ) , .B1( us13_n832 ) , .A1( us13_n839 ) , .C1( us13_n842 ) , .C2( us13_n851 ) , .A2( us13_n855 ) , .B2( us13_n865 ) );
  NOR4_X1 us13_U65 (.A1( us13_n466 ) , .ZN( us13_n467 ) , .A4( us13_n542 ) , .A2( us13_n554 ) , .A3( us13_n614 ) );
  AOI221_X1 us13_U66 (.ZN( us13_n468 ) , .C2( us13_n714 ) , .B2( us13_n831 ) , .C1( us13_n845 ) , .B1( us13_n860 ) , .A( us13_n864 ) );
  NAND4_X1 us13_U67 (.A4( us13_n485 ) , .A3( us13_n486 ) , .A2( us13_n487 ) , .A1( us13_n488 ) , .ZN( us13_n778 ) );
  NOR4_X1 us13_U68 (.A4( us13_n484 ) , .ZN( us13_n487 ) , .A1( us13_n566 ) , .A2( us13_n581 ) , .A3( us13_n602 ) );
  NOR4_X1 us13_U69 (.ZN( us13_n486 ) , .A1( us13_n507 ) , .A2( us13_n519 ) , .A4( us13_n546 ) , .A3( us13_n611 ) );
  NOR3_X1 us13_U7 (.A3( us13_n800 ) , .A2( us13_n801 ) , .A1( us13_n802 ) , .ZN( us13_n825 ) );
  NOR4_X1 us13_U70 (.A4( us13_n514 ) , .A3( us13_n515 ) , .A2( us13_n516 ) , .A1( us13_n517 ) , .ZN( us13_n524 ) );
  AOI222_X1 us13_U71 (.ZN( us13_n525 ) , .A1( us13_n834 ) , .B2( us13_n837 ) , .C1( us13_n844 ) , .C2( us13_n850 ) , .A2( us13_n852 ) , .B1( us13_n866 ) );
  NOR4_X1 us13_U72 (.A3( us13_n521 ) , .A1( us13_n522 ) , .ZN( us13_n523 ) , .A2( us13_n673 ) , .A4( us13_n769 ) );
  NAND4_X1 us13_U73 (.A4( us13_n657 ) , .A3( us13_n658 ) , .A2( us13_n659 ) , .A1( us13_n660 ) , .ZN( us13_n800 ) );
  NOR3_X1 us13_U74 (.A3( us13_n651 ) , .A2( us13_n652 ) , .A1( us13_n653 ) , .ZN( us13_n658 ) );
  NOR3_X1 us13_U75 (.A3( us13_n648 ) , .A2( us13_n649 ) , .A1( us13_n650 ) , .ZN( us13_n659 ) );
  NOR3_X1 us13_U76 (.A3( us13_n654 ) , .A2( us13_n655 ) , .A1( us13_n656 ) , .ZN( us13_n657 ) );
  NAND4_X1 us13_U77 (.A4( us13_n560 ) , .A3( us13_n561 ) , .A2( us13_n562 ) , .A1( us13_n563 ) , .ZN( us13_n607 ) );
  NOR4_X1 us13_U78 (.A4( us13_n552 ) , .A3( us13_n553 ) , .A2( us13_n554 ) , .A1( us13_n555 ) , .ZN( us13_n562 ) );
  NOR4_X1 us13_U79 (.ZN( us13_n561 ) , .A1( us13_n653 ) , .A3( us13_n661 ) , .A4( us13_n685 ) , .A2( us13_n768 ) );
  NOR3_X1 us13_U8 (.ZN( us13_n504 ) , .A2( us13_n679 ) , .A3( us13_n777 ) , .A1( us13_n876 ) );
  NOR4_X1 us13_U80 (.A4( us13_n556 ) , .A3( us13_n557 ) , .A2( us13_n558 ) , .A1( us13_n559 ) , .ZN( us13_n560 ) );
  NAND4_X1 us13_U81 (.A4( us13_n772 ) , .A3( us13_n773 ) , .A2( us13_n774 ) , .A1( us13_n775 ) , .ZN( us13_n801 ) );
  NOR3_X1 us13_U82 (.A3( us13_n765 ) , .A2( us13_n766 ) , .A1( us13_n767 ) , .ZN( us13_n773 ) );
  AOI222_X1 us13_U83 (.ZN( us13_n775 ) , .A1( us13_n830 ) , .C1( us13_n834 ) , .B2( us13_n841 ) , .A2( us13_n850 ) , .B1( us13_n861 ) , .C2( us13_n873 ) );
  NOR4_X1 us13_U84 (.A4( us13_n768 ) , .A3( us13_n769 ) , .A2( us13_n770 ) , .A1( us13_n771 ) , .ZN( us13_n772 ) );
  NAND4_X1 us13_U85 (.A4( us13_n691 ) , .A3( us13_n692 ) , .A1( us13_n693 ) , .ZN( us13_n776 ) , .A2( us13_n872 ) );
  INV_X1 us13_U86 (.A( us13_n679 ) , .ZN( us13_n872 ) );
  NOR4_X1 us13_U87 (.A4( us13_n687 ) , .A3( us13_n688 ) , .A2( us13_n689 ) , .A1( us13_n690 ) , .ZN( us13_n691 ) );
  NOR4_X1 us13_U88 (.A4( us13_n661 ) , .A3( us13_n662 ) , .A2( us13_n663 ) , .A1( us13_n664 ) , .ZN( us13_n677 ) );
  NOR4_X1 us13_U89 (.A4( us13_n665 ) , .A3( us13_n666 ) , .A2( us13_n667 ) , .A1( us13_n668 ) , .ZN( us13_n676 ) );
  INV_X1 us13_U9 (.A( us13_n706 ) , .ZN( us13_n876 ) );
  NOR4_X1 us13_U90 (.A3( us13_n673 ) , .A1( us13_n674 ) , .ZN( us13_n675 ) , .A4( us13_n715 ) , .A2( us13_n859 ) );
  NOR2_X1 us13_U91 (.ZN( us13_n761 ) , .A1( us13_n833 ) , .A2( us13_n834 ) );
  NOR4_X1 us13_U92 (.A4( us13_n577 ) , .A3( us13_n578 ) , .A2( us13_n579 ) , .ZN( us13_n586 ) , .A1( us13_n683 ) );
  NOR4_X1 us13_U93 (.A1( us13_n584 ) , .ZN( us13_n585 ) , .A3( us13_n652 ) , .A2( us13_n662 ) , .A4( us13_n767 ) );
  AOI222_X1 us13_U94 (.ZN( us13_n513 ) , .C1( us13_n832 ) , .B2( us13_n837 ) , .A2( us13_n843 ) , .C2( us13_n862 ) , .B1( us13_n863 ) , .A1( us13_n866 ) );
  NOR4_X1 us13_U95 (.A4( us13_n509 ) , .A2( us13_n510 ) , .A1( us13_n511 ) , .ZN( us13_n512 ) , .A3( us13_n670 ) );
  INV_X1 us13_U96 (.A( us13_n505 ) , .ZN( us13_n871 ) );
  NAND4_X1 us13_U97 (.A4( us13_n456 ) , .A3( us13_n457 ) , .A2( us13_n458 ) , .A1( us13_n459 ) , .ZN( us13_n679 ) );
  NOR3_X1 us13_U98 (.ZN( us13_n457 ) , .A3( us13_n530 ) , .A1( us13_n555 ) , .A2( us13_n570 ) );
  AOI221_X1 us13_U99 (.A( us13_n450 ) , .ZN( us13_n459 ) , .C2( us13_n753 ) , .B1( us13_n832 ) , .C1( us13_n842 ) , .B2( us13_n861 ) );
  NOR3_X1 us21_U10 (.A3( us21_n619 ) , .A2( us21_n620 ) , .ZN( us21_n634 ) , .A1( us21_n723 ) );
  NOR4_X1 us21_U100 (.A4( us21_n524 ) , .A2( us21_n525 ) , .A1( us21_n526 ) , .ZN( us21_n536 ) , .A3( us21_n699 ) );
  NOR4_X1 us21_U101 (.A1( us21_n529 ) , .ZN( us21_n534 ) , .A2( us21_n652 ) , .A4( us21_n666 ) , .A3( us21_n763 ) );
  NOR4_X1 us21_U102 (.A4( us21_n527 ) , .A3( us21_n528 ) , .ZN( us21_n535 ) , .A2( us21_n682 ) , .A1( us21_n792 ) );
  NAND4_X1 us21_U103 (.A4( us21_n546 ) , .A3( us21_n547 ) , .A2( us21_n548 ) , .A1( us21_n549 ) , .ZN( us21_n743 ) );
  NOR3_X1 us21_U104 (.ZN( us21_n547 ) , .A2( us21_n649 ) , .A1( us21_n665 ) , .A3( us21_n769 ) );
  AOI211_X1 us21_U105 (.B( us21_n537 ) , .A( us21_n538 ) , .ZN( us21_n549 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NOR4_X1 us21_U106 (.A4( us21_n539 ) , .A3( us21_n540 ) , .A2( us21_n541 ) , .ZN( us21_n548 ) , .A1( us21_n686 ) );
  NAND4_X1 us21_U107 (.A4( us21_n477 ) , .A3( us21_n478 ) , .A2( us21_n479 ) , .A1( us21_n480 ) , .ZN( us21_n692 ) );
  NOR3_X1 us21_U108 (.ZN( us21_n478 ) , .A2( us21_n506 ) , .A3( us21_n599 ) , .A1( us21_n608 ) );
  AOI211_X1 us21_U109 (.B( us21_n475 ) , .A( us21_n476 ) , .ZN( us21_n480 ) , .C2( us21_n831 ) , .C1( us21_n859 ) );
  NOR2_X1 us21_U11 (.ZN( us21_n493 ) , .A1( us21_n676 ) , .A2( us21_n692 ) );
  NOR4_X1 us21_U110 (.ZN( us21_n479 ) , .A3( us21_n530 ) , .A4( us21_n543 ) , .A2( us21_n565 ) , .A1( us21_n715 ) );
  NOR4_X1 us21_U111 (.A4( us21_n607 ) , .A3( us21_n608 ) , .A2( us21_n609 ) , .A1( us21_n610 ) , .ZN( us21_n617 ) );
  NOR4_X1 us21_U112 (.ZN( us21_n618 ) , .A1( us21_n654 ) , .A3( us21_n664 ) , .A4( us21_n680 ) , .A2( us21_n764 ) );
  NOR4_X1 us21_U113 (.A4( us21_n612 ) , .A3( us21_n613 ) , .A2( us21_n614 ) , .A1( us21_n615 ) , .ZN( us21_n616 ) );
  NOR2_X1 us21_U114 (.ZN( us21_n684 ) , .A1( us21_n829 ) , .A2( us21_n830 ) );
  NAND4_X1 us21_U115 (.A4( us21_n471 ) , .A3( us21_n472 ) , .A2( us21_n473 ) , .A1( us21_n474 ) , .ZN( us21_n676 ) );
  NOR4_X1 us21_U116 (.A4( us21_n468 ) , .ZN( us21_n474 ) , .A3( us21_n554 ) , .A1( us21_n733 ) , .A2( us21_n753 ) );
  NOR4_X1 us21_U117 (.ZN( us21_n473 ) , .A1( us21_n529 ) , .A3( us21_n566 ) , .A4( us21_n598 ) , .A2( us21_n640 ) );
  NOR4_X1 us21_U118 (.ZN( us21_n472 ) , .A1( us21_n504 ) , .A3( us21_n542 ) , .A2( us21_n581 ) , .A4( us21_n714 ) );
  NAND4_X1 us21_U119 (.A4( us21_n689 ) , .A3( us21_n690 ) , .A1( us21_n691 ) , .ZN( us21_n774 ) , .A2( us21_n870 ) );
  NOR2_X1 us21_U12 (.A1( us21_n676 ) , .ZN( us21_n691 ) , .A2( us21_n805 ) );
  INV_X1 us21_U120 (.A( us21_n677 ) , .ZN( us21_n870 ) );
  AOI221_X1 us21_U121 (.A( us21_n679 ) , .ZN( us21_n690 ) , .B2( us21_n838 ) , .C1( us21_n840 ) , .C2( us21_n860 ) , .B1( us21_n863 ) );
  NOR4_X1 us21_U122 (.A4( us21_n685 ) , .A3( us21_n686 ) , .A2( us21_n687 ) , .A1( us21_n688 ) , .ZN( us21_n689 ) );
  NOR2_X1 us21_U123 (.ZN( us21_n731 ) , .A2( us21_n830 ) , .A1( us21_n843 ) );
  NAND4_X1 us21_U124 (.A4( us21_n717 ) , .A3( us21_n718 ) , .A2( us21_n719 ) , .ZN( us21_n739 ) , .A1( us21_n855 ) );
  INV_X1 us21_U125 (.A( us21_n707 ) , .ZN( us21_n855 ) );
  NOR4_X1 us21_U126 (.A4( us21_n713 ) , .A3( us21_n714 ) , .A2( us21_n715 ) , .A1( us21_n716 ) , .ZN( us21_n717 ) );
  AOI221_X1 us21_U127 (.A( us21_n708 ) , .ZN( us21_n719 ) , .C2( us21_n842 ) , .B2( us21_n843 ) , .C1( us21_n859 ) , .B1( us21_n860 ) );
  NAND4_X1 us21_U128 (.A4( us21_n571 ) , .A3( us21_n572 ) , .A1( us21_n573 ) , .ZN( us21_n721 ) , .A2( us21_n872 ) );
  NOR4_X1 us21_U129 (.A4( us21_n567 ) , .A3( us21_n568 ) , .A2( us21_n569 ) , .A1( us21_n570 ) , .ZN( us21_n571 ) );
  INV_X1 us21_U13 (.A( us21_n605 ) , .ZN( us21_n872 ) );
  AOI221_X1 us21_U130 (.A( us21_n562 ) , .C2( us21_n563 ) , .ZN( us21_n572 ) , .B2( us21_n843 ) , .B1( us21_n850 ) , .C1( us21_n851 ) );
  NOR2_X1 us21_U131 (.ZN( us21_n573 ) , .A1( us21_n620 ) , .A2( us21_n743 ) );
  NAND4_X1 us21_U132 (.A4( us21_n491 ) , .A3( us21_n492 ) , .A1( us21_n493 ) , .ZN( us21_n800 ) , .A2( us21_n865 ) );
  AOI221_X1 us21_U133 (.A( us21_n487 ) , .ZN( us21_n492 ) , .B2( us21_n834 ) , .C2( us21_n839 ) , .C1( us21_n849 ) , .B1( us21_n858 ) );
  INV_X1 us21_U134 (.A( us21_n776 ) , .ZN( us21_n865 ) );
  NOR4_X1 us21_U135 (.A2( us21_n489 ) , .A1( us21_n490 ) , .ZN( us21_n491 ) , .A3( us21_n578 ) , .A4( us21_n610 ) );
  INV_X1 us21_U136 (.A( us21_n760 ) , .ZN( us21_n828 ) );
  NOR2_X1 us21_U137 (.ZN( us21_n645 ) , .A1( us21_n852 ) , .A2( us21_n866 ) );
  INV_X1 us21_U138 (.A( us21_n461 ) , .ZN( us21_n862 ) );
  OAI21_X1 us21_U139 (.ZN( us21_n461 ) , .B1( us21_n807 ) , .A( us21_n832 ) , .B2( us21_n849 ) );
  INV_X1 us21_U14 (.A( us21_n678 ) , .ZN( us21_n838 ) );
  OR4_X1 us21_U140 (.ZN( us21_n490 ) , .A4( us21_n532 ) , .A2( us21_n545 ) , .A1( us21_n557 ) , .A3( us21_n630 ) );
  OR4_X1 us21_U141 (.A4( us21_n564 ) , .A3( us21_n565 ) , .A2( us21_n566 ) , .ZN( us21_n570 ) , .A1( us21_n663 ) );
  OR4_X1 us21_U142 (.A4( us21_n680 ) , .A3( us21_n681 ) , .A2( us21_n682 ) , .A1( us21_n683 ) , .ZN( us21_n688 ) );
  OR4_X1 us21_U143 (.ZN( us21_n464 ) , .A4( us21_n516 ) , .A3( us21_n527 ) , .A2( us21_n576 ) , .A1( us21_n710 ) );
  OR4_X1 us21_U144 (.A4( us21_n516 ) , .A2( us21_n517 ) , .A1( us21_n518 ) , .ZN( us21_n520 ) , .A3( us21_n819 ) );
  OR4_X1 us21_U145 (.A4( us21_n578 ) , .A3( us21_n579 ) , .A2( us21_n580 ) , .A1( us21_n581 ) , .ZN( us21_n582 ) );
  NAND2_X1 us21_U146 (.ZN( us21_n611 ) , .A2( us21_n835 ) , .A1( us21_n871 ) );
  OR3_X1 us21_U147 (.A3( us21_n504 ) , .A2( us21_n505 ) , .A1( us21_n506 ) , .ZN( us21_n509 ) );
  AOI221_X1 us21_U148 (.A( us21_n711 ) , .B2( us21_n712 ) , .ZN( us21_n718 ) , .C1( us21_n830 ) , .B1( us21_n837 ) , .C2( us21_n861 ) );
  OR2_X1 us21_U149 (.A2( us21_n709 ) , .A1( us21_n710 ) , .ZN( us21_n711 ) );
  NOR4_X1 us21_U15 (.A4( us21_n443 ) , .A3( us21_n444 ) , .A2( us21_n514 ) , .A1( us21_n539 ) , .ZN( us21_n704 ) );
  INV_X1 us21_U150 (.A( us21_n752 ) , .ZN( us21_n867 ) );
  OAI21_X1 us21_U151 (.B1( us21_n751 ) , .ZN( us21_n752 ) , .A( us21_n843 ) , .B2( us21_n866 ) );
  INV_X1 us21_U152 (.A( us21_n670 ) , .ZN( us21_n857 ) );
  AOI21_X1 us21_U153 (.A( us21_n668 ) , .B1( us21_n669 ) , .ZN( us21_n670 ) , .B2( us21_n854 ) );
  AOI222_X1 us21_U154 (.ZN( us21_n658 ) , .A2( us21_n837 ) , .B1( us21_n839 ) , .C2( us21_n843 ) , .A1( us21_n858 ) , .C1( us21_n861 ) , .B2( us21_n868 ) );
  INV_X1 us21_U155 (.A( us21_n645 ) , .ZN( us21_n868 ) );
  OAI22_X1 us21_U156 (.ZN( us21_n481 ) , .A1( us21_n706 ) , .B2( us21_n783 ) , .A2( us21_n804 ) , .B1( us21_n810 ) );
  OAI22_X1 us21_U157 (.ZN( us21_n635 ) , .A1( us21_n697 ) , .B2( us21_n726 ) , .A2( us21_n760 ) , .B1( us21_n814 ) );
  OAI222_X1 us21_U158 (.B2( us21_n706 ) , .ZN( us21_n707 ) , .C2( us21_n722 ) , .B1( us21_n745 ) , .A1( us21_n804 ) , .C1( us21_n812 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U159 (.A1( us21_n445 ) , .A2( us21_n463 ) , .ZN( us21_n747 ) );
  OR3_X1 us21_U16 (.ZN( us21_n444 ) , .A1( us21_n526 ) , .A3( us21_n575 ) , .A2( us21_n873 ) );
  AOI22_X1 us21_U160 (.ZN( us21_n694 ) , .A1( us21_n828 ) , .B2( us21_n841 ) , .A2( us21_n863 ) , .B1( us21_n866 ) );
  INV_X1 us21_U161 (.A( us21_n728 ) , .ZN( us21_n837 ) );
  NAND2_X1 us21_U162 (.A1( us21_n449 ) , .A2( us21_n451 ) , .ZN( us21_n760 ) );
  INV_X1 us21_U163 (.A( us21_n788 ) , .ZN( us21_n830 ) );
  OAI221_X1 us21_U164 (.A( us21_n725 ) , .C2( us21_n726 ) , .B2( us21_n727 ) , .B1( us21_n728 ) , .ZN( us21_n735 ) , .C1( us21_n815 ) );
  AOI22_X1 us21_U165 (.ZN( us21_n725 ) , .B1( us21_n830 ) , .A2( us21_n836 ) , .A1( us21_n861 ) , .B2( us21_n864 ) );
  AND2_X1 us21_U166 (.ZN( us21_n746 ) , .A1( us21_n782 ) , .A2( us21_n784 ) );
  OAI22_X1 us21_U167 (.ZN( us21_n487 ) , .A1( us21_n722 ) , .B2( us21_n726 ) , .B1( us21_n728 ) , .A2( us21_n777 ) );
  OAI22_X1 us21_U168 (.ZN( us21_n622 ) , .B1( us21_n667 ) , .B2( us21_n745 ) , .A1( us21_n813 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U169 (.B2( us21_n777 ) , .B1( us21_n778 ) , .ZN( us21_n779 ) , .A2( us21_n812 ) , .A1( us21_n813 ) );
  OR4_X1 us21_U17 (.A4( us21_n440 ) , .A2( us21_n441 ) , .A1( us21_n442 ) , .ZN( us21_n443 ) , .A3( us21_n551 ) );
  OAI22_X1 us21_U170 (.A1( us21_n722 ) , .ZN( us21_n724 ) , .B2( us21_n748 ) , .B1( us21_n810 ) , .A2( us21_n814 ) );
  OAI22_X1 us21_U171 (.B2( us21_n742 ) , .ZN( us21_n744 ) , .A2( us21_n760 ) , .B1( us21_n778 ) , .A1( us21_n790 ) );
  OAI22_X1 us21_U172 (.B2( us21_n801 ) , .B1( us21_n802 ) , .A2( us21_n803 ) , .A1( us21_n804 ) , .ZN( us21_n806 ) );
  OAI22_X1 us21_U173 (.ZN( us21_n494 ) , .A2( us21_n742 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n804 ) );
  INV_X1 us21_U174 (.A( us21_n742 ) , .ZN( us21_n835 ) );
  INV_X1 us21_U175 (.A( us21_n786 ) , .ZN( us21_n843 ) );
  INV_X1 us21_U176 (.A( us21_n814 ) , .ZN( us21_n829 ) );
  OAI22_X1 us21_U177 (.B1( us21_n488 ) , .ZN( us21_n489 ) , .A1( us21_n684 ) , .A2( us21_n761 ) , .B2( us21_n815 ) );
  NOR3_X1 us21_U178 (.ZN( us21_n488 ) , .A1( us21_n780 ) , .A2( us21_n848 ) , .A3( us21_n861 ) );
  OAI22_X1 us21_U179 (.ZN( us21_n588 ) , .B1( us21_n728 ) , .B2( us21_n747 ) , .A2( us21_n784 ) , .A1( us21_n801 ) );
  INV_X1 us21_U18 (.A( us21_n611 ) , .ZN( us21_n873 ) );
  OAI22_X1 us21_U180 (.ZN( us21_n693 ) , .A2( us21_n728 ) , .A1( us21_n778 ) , .B1( us21_n789 ) , .B2( us21_n815 ) );
  OAI22_X1 us21_U181 (.ZN( us21_n708 ) , .A2( us21_n726 ) , .B2( us21_n727 ) , .A1( us21_n742 ) , .B1( us21_n811 ) );
  INV_X1 us21_U182 (.A( us21_n812 ) , .ZN( us21_n831 ) );
  INV_X1 us21_U183 (.A( us21_n667 ) , .ZN( us21_n863 ) );
  NOR2_X1 us21_U184 (.ZN( us21_n716 ) , .A2( us21_n722 ) , .A1( us21_n742 ) );
  NOR2_X1 us21_U185 (.ZN( us21_n664 ) , .A1( us21_n726 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U186 (.ZN( us21_n568 ) , .A1( us21_n726 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U187 (.ZN( us21_n544 ) , .A2( us21_n778 ) , .A1( us21_n812 ) );
  INV_X1 us21_U188 (.A( us21_n748 ) , .ZN( us21_n840 ) );
  NOR2_X1 us21_U189 (.ZN( us21_n530 ) , .A2( us21_n747 ) , .A1( us21_n748 ) );
  INV_X1 us21_U19 (.A( us21_n747 ) , .ZN( us21_n861 ) );
  NOR2_X1 us21_U190 (.ZN( us21_n575 ) , .A2( us21_n697 ) , .A1( us21_n812 ) );
  NOR2_X1 us21_U191 (.ZN( us21_n652 ) , .A1( us21_n726 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U192 (.ZN( us21_n613 ) , .A1( us21_n783 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U193 (.ZN( us21_n627 ) , .A2( us21_n726 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U194 (.ZN( us21_n599 ) , .A2( us21_n778 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U195 (.ZN( us21_n610 ) , .A1( us21_n777 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U196 (.ZN( us21_n526 ) , .A2( us21_n722 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U197 (.ZN( us21_n626 ) , .A2( us21_n667 ) , .A1( us21_n783 ) );
  INV_X1 us21_U198 (.A( us21_n790 ) , .ZN( us21_n849 ) );
  NOR2_X1 us21_U199 (.A2( us21_n742 ) , .ZN( us21_n767 ) , .A1( us21_n810 ) );
  AOI222_X1 us21_U20 (.ZN( us21_n561 ) , .B1( us21_n828 ) , .C1( us21_n839 ) , .A2( us21_n841 ) , .A1( us21_n852 ) , .B2( us21_n861 ) , .C2( us21_n871 ) );
  NOR2_X1 us21_U200 (.ZN( us21_n529 ) , .A2( us21_n778 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U201 (.A2( us21_n706 ) , .A1( us21_n748 ) , .ZN( us21_n769 ) );
  NOR2_X1 us21_U202 (.ZN( us21_n597 ) , .A2( us21_n789 ) , .A1( us21_n814 ) );
  NOR2_X1 us21_U203 (.ZN( us21_n609 ) , .A2( us21_n778 ) , .A1( us21_n804 ) );
  NOR2_X1 us21_U204 (.ZN( us21_n650 ) , .A1( us21_n667 ) , .A2( us21_n812 ) );
  INV_X1 us21_U205 (.A( us21_n745 ) , .ZN( us21_n832 ) );
  NOR2_X1 us21_U206 (.A1( us21_n667 ) , .ZN( us21_n671 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U207 (.ZN( us21_n600 ) , .A1( us21_n667 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U208 (.A1( us21_n667 ) , .ZN( us21_n686 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U209 (.ZN( us21_n665 ) , .A1( us21_n748 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U21 (.ZN( us21_n471 ) , .A2( us21_n519 ) , .A4( us21_n592 ) , .A1( us21_n607 ) , .A3( us21_n627 ) );
  NOR2_X1 us21_U210 (.ZN( us21_n553 ) , .A1( us21_n748 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U211 (.ZN( us21_n506 ) , .A2( us21_n778 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U212 (.ZN( us21_n541 ) , .A2( us21_n706 ) , .A1( us21_n783 ) );
  NOR2_X1 us21_U213 (.ZN( us21_n662 ) , .A1( us21_n783 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U214 (.A1( us21_n667 ) , .ZN( us21_n764 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U215 (.A1( us21_n697 ) , .ZN( us21_n766 ) , .A2( us21_n811 ) );
  OAI22_X1 us21_U216 (.B1( us21_n438 ) , .ZN( us21_n442 ) , .A2( us21_n726 ) , .A1( us21_n742 ) , .B2( us21_n747 ) );
  NOR3_X1 us21_U217 (.ZN( us21_n438 ) , .A2( us21_n834 ) , .A3( us21_n835 ) , .A1( us21_n844 ) );
  NOR2_X1 us21_U218 (.ZN( us21_n525 ) , .A1( us21_n667 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U219 (.ZN( us21_n505 ) , .A1( us21_n810 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U22 (.A4( us21_n542 ) , .A3( us21_n543 ) , .A2( us21_n544 ) , .A1( us21_n545 ) , .ZN( us21_n546 ) );
  NOR2_X1 us21_U220 (.ZN( us21_n659 ) , .A1( us21_n727 ) , .A2( us21_n788 ) );
  INV_X1 us21_U221 (.A( us21_n801 ) , .ZN( us21_n841 ) );
  NOR2_X1 us21_U222 (.ZN( us21_n555 ) , .A1( us21_n790 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U223 (.ZN( us21_n543 ) , .A1( us21_n747 ) , .A2( us21_n812 ) );
  NOR2_X1 us21_U224 (.ZN( us21_n507 ) , .A1( us21_n727 ) , .A2( us21_n777 ) );
  NOR2_X1 us21_U225 (.ZN( us21_n528 ) , .A2( us21_n742 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U226 (.A1( us21_n747 ) , .ZN( us21_n765 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U227 (.A2( us21_n742 ) , .ZN( us21_n753 ) , .A1( us21_n803 ) );
  OAI22_X1 us21_U228 (.B2( us21_n748 ) , .B1( us21_n749 ) , .A1( us21_n750 ) , .ZN( us21_n754 ) , .A2( us21_n804 ) );
  NOR2_X1 us21_U229 (.ZN( us21_n749 ) , .A2( us21_n850 ) , .A1( us21_n858 ) );
  NOR4_X1 us21_U23 (.ZN( us21_n477 ) , .A1( us21_n518 ) , .A4( us21_n555 ) , .A3( us21_n580 ) , .A2( us21_n628 ) );
  NOR3_X1 us21_U230 (.ZN( us21_n750 ) , .A2( us21_n851 ) , .A1( us21_n861 ) , .A3( us21_n863 ) );
  NOR2_X1 us21_U231 (.ZN( us21_n542 ) , .A2( us21_n783 ) , .A1( us21_n790 ) );
  INV_X1 us21_U232 (.A( us21_n804 ) , .ZN( us21_n839 ) );
  NOR2_X1 us21_U233 (.ZN( us21_n629 ) , .A1( us21_n722 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U234 (.ZN( us21_n733 ) , .A2( us21_n801 ) , .A1( us21_n803 ) );
  NOR2_X1 us21_U235 (.ZN( us21_n514 ) , .A1( us21_n706 ) , .A2( us21_n742 ) );
  NOR2_X1 us21_U236 (.ZN( us21_n661 ) , .A1( us21_n727 ) , .A2( us21_n783 ) );
  NOR2_X1 us21_U237 (.ZN( us21_n715 ) , .A2( us21_n742 ) , .A1( us21_n784 ) );
  NOR2_X1 us21_U238 (.ZN( us21_n612 ) , .A1( us21_n760 ) , .A2( us21_n810 ) );
  INV_X1 us21_U239 (.A( us21_n726 ) , .ZN( us21_n850 ) );
  NOR4_X1 us21_U24 (.ZN( us21_n454 ) , .A2( us21_n515 ) , .A1( us21_n541 ) , .A3( us21_n577 ) , .A4( us21_n613 ) );
  NOR2_X1 us21_U240 (.ZN( us21_n552 ) , .A1( us21_n784 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U241 (.ZN( us21_n515 ) , .A1( us21_n706 ) , .A2( us21_n801 ) );
  NOR2_X1 us21_U242 (.ZN( us21_n504 ) , .A2( us21_n726 ) , .A1( us21_n760 ) );
  NOR2_X1 us21_U243 (.ZN( us21_n556 ) , .A1( us21_n706 ) , .A2( us21_n814 ) );
  NOR2_X1 us21_U244 (.ZN( us21_n519 ) , .A1( us21_n788 ) , .A2( us21_n810 ) );
  INV_X1 us21_U245 (.A( us21_n803 ) , .ZN( us21_n858 ) );
  NOR2_X1 us21_U246 (.ZN( us21_n713 ) , .A1( us21_n803 ) , .A2( us21_n815 ) );
  NOR2_X1 us21_U247 (.ZN( us21_n653 ) , .A1( us21_n788 ) , .A2( us21_n813 ) );
  NOR2_X1 us21_U248 (.ZN( us21_n666 ) , .A2( us21_n706 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U249 (.ZN( us21_n628 ) , .A1( us21_n745 ) , .A2( us21_n813 ) );
  NOR4_X1 us21_U25 (.A4( us21_n530 ) , .A3( us21_n531 ) , .A2( us21_n532 ) , .ZN( us21_n533 ) , .A1( us21_n818 ) );
  NOR2_X1 us21_U250 (.ZN( us21_n554 ) , .A1( us21_n760 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U251 (.ZN( us21_n540 ) , .A1( us21_n760 ) , .A2( us21_n789 ) );
  NOR2_X1 us21_U252 (.ZN( us21_n699 ) , .A2( us21_n784 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U253 (.A1( us21_n728 ) , .ZN( us21_n763 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U254 (.ZN( us21_n607 ) , .A2( us21_n722 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U255 (.ZN( us21_n577 ) , .A2( us21_n706 ) , .A1( us21_n728 ) );
  NOR2_X1 us21_U256 (.ZN( us21_n531 ) , .A2( us21_n722 ) , .A1( us21_n728 ) );
  AOI21_X1 us21_U257 (.A( us21_n810 ) , .B2( us21_n811 ) , .B1( us21_n812 ) , .ZN( us21_n817 ) );
  AOI21_X1 us21_U258 (.ZN( us21_n513 ) , .A( us21_n727 ) , .B1( us21_n748 ) , .B2( us21_n801 ) );
  NOR2_X1 us21_U259 (.ZN( us21_n654 ) , .A1( us21_n745 ) , .A2( us21_n778 ) );
  NOR2_X1 us21_U26 (.ZN( us21_n678 ) , .A2( us21_n832 ) , .A1( us21_n837 ) );
  AOI21_X1 us21_U260 (.A( us21_n813 ) , .B2( us21_n814 ) , .B1( us21_n815 ) , .ZN( us21_n816 ) );
  NOR2_X1 us21_U261 (.ZN( us21_n580 ) , .A1( us21_n742 ) , .A2( us21_n813 ) );
  AOI21_X1 us21_U262 (.ZN( us21_n591 ) , .B1( us21_n748 ) , .A( us21_n790 ) , .B2( us21_n811 ) );
  AOI21_X1 us21_U263 (.B1( us21_n623 ) , .ZN( us21_n625 ) , .A( us21_n761 ) , .B2( us21_n812 ) );
  NOR2_X1 us21_U264 (.A2( us21_n706 ) , .A1( us21_n760 ) , .ZN( us21_n792 ) );
  NOR2_X1 us21_U265 (.ZN( us21_n640 ) , .A2( us21_n786 ) , .A1( us21_n789 ) );
  AOI21_X1 us21_U266 (.ZN( us21_n497 ) , .B1( us21_n678 ) , .A( us21_n810 ) , .B2( us21_n814 ) );
  NOR2_X1 us21_U267 (.ZN( us21_n668 ) , .A1( us21_n788 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U268 (.ZN( us21_n557 ) , .A2( us21_n789 ) , .A1( us21_n801 ) );
  AOI21_X1 us21_U269 (.ZN( us21_n624 ) , .B2( us21_n667 ) , .A( us21_n788 ) , .B1( us21_n789 ) );
  NOR4_X1 us21_U27 (.A4( us21_n575 ) , .A3( us21_n576 ) , .A2( us21_n577 ) , .ZN( us21_n584 ) , .A1( us21_n681 ) );
  NOR2_X1 us21_U270 (.ZN( us21_n681 ) , .A2( us21_n697 ) , .A1( us21_n801 ) );
  NOR2_X1 us21_U271 (.ZN( us21_n651 ) , .A1( us21_n760 ) , .A2( us21_n784 ) );
  NOR2_X1 us21_U272 (.ZN( us21_n518 ) , .A2( us21_n706 ) , .A1( us21_n812 ) );
  INV_X1 us21_U273 (.A( us21_n811 ) , .ZN( us21_n834 ) );
  NOR2_X1 us21_U274 (.ZN( us21_n517 ) , .A2( us21_n697 ) , .A1( us21_n814 ) );
  AOI21_X1 us21_U275 (.ZN( us21_n475 ) , .A( us21_n667 ) , .B1( us21_n748 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U276 (.ZN( us21_n508 ) , .B2( us21_n667 ) , .A( us21_n728 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U277 (.ZN( us21_n537 ) , .B2( us21_n810 ) , .A( us21_n812 ) , .B1( us21_n813 ) );
  INV_X1 us21_U278 (.A( us21_n761 ) , .ZN( us21_n864 ) );
  AOI21_X1 us21_U279 (.ZN( us21_n538 ) , .A( us21_n761 ) , .B2( us21_n777 ) , .B1( us21_n815 ) );
  NOR4_X1 us21_U28 (.A1( us21_n582 ) , .ZN( us21_n583 ) , .A3( us21_n650 ) , .A2( us21_n660 ) , .A4( us21_n765 ) );
  NOR2_X1 us21_U280 (.ZN( us21_n579 ) , .A1( us21_n667 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U281 (.ZN( us21_n587 ) , .B2( us21_n697 ) , .B1( us21_n813 ) , .A( us21_n815 ) );
  AOI21_X1 us21_U282 (.ZN( us21_n589 ) , .B2( us21_n761 ) , .A( us21_n783 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U283 (.B1( us21_n697 ) , .ZN( us21_n698 ) , .A( us21_n730 ) , .B2( us21_n761 ) );
  AOI21_X1 us21_U284 (.ZN( us21_n638 ) , .B2( us21_n745 ) , .A( us21_n790 ) , .B1( us21_n801 ) );
  AOI21_X1 us21_U285 (.ZN( us21_n496 ) , .A( us21_n722 ) , .B2( us21_n760 ) , .B1( us21_n812 ) );
  INV_X1 us21_U286 (.A( us21_n789 ) , .ZN( us21_n871 ) );
  NOR2_X1 us21_U287 (.ZN( us21_n545 ) , .A1( us21_n697 ) , .A2( us21_n742 ) );
  INV_X1 us21_U288 (.A( us21_n727 ) , .ZN( us21_n866 ) );
  AOI21_X1 us21_U289 (.ZN( us21_n647 ) , .B1( us21_n727 ) , .B2( us21_n761 ) , .A( us21_n811 ) );
  AOI221_X1 us21_U29 (.A( us21_n779 ) , .ZN( us21_n796 ) , .C2( us21_n835 ) , .B2( us21_n836 ) , .B1( us21_n863 ) , .C1( us21_n864 ) );
  AOI21_X1 us21_U290 (.ZN( us21_n567 ) , .B1( us21_n748 ) , .B2( us21_n760 ) , .A( us21_n778 ) );
  INV_X1 us21_U291 (.A( us21_n810 ) , .ZN( us21_n852 ) );
  NOR2_X1 us21_U292 (.ZN( us21_n683 ) , .A1( us21_n727 ) , .A2( us21_n814 ) );
  AOI21_X1 us21_U293 (.B1( us21_n684 ) , .ZN( us21_n685 ) , .A( us21_n726 ) , .B2( us21_n759 ) );
  NOR2_X1 us21_U294 (.ZN( us21_n566 ) , .A1( us21_n727 ) , .A2( us21_n760 ) );
  NOR2_X1 us21_U295 (.ZN( us21_n663 ) , .A1( us21_n778 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U296 (.ZN( us21_n448 ) , .B2( us21_n790 ) , .A( us21_n801 ) , .B1( us21_n813 ) );
  AOI21_X1 us21_U297 (.ZN( us21_n512 ) , .A( us21_n777 ) , .B2( us21_n790 ) , .B1( us21_n810 ) );
  AOI21_X1 us21_U298 (.ZN( us21_n637 ) , .B2( us21_n747 ) , .A( us21_n786 ) , .B1( us21_n810 ) );
  INV_X1 us21_U299 (.A( us21_n697 ) , .ZN( us21_n851 ) );
  NAND2_X2 us21_U3 (.A2( us21_n458 ) , .A1( us21_n463 ) , .ZN( us21_n778 ) );
  NOR4_X1 us21_U30 (.A4( us21_n791 ) , .A3( us21_n792 ) , .A2( us21_n793 ) , .A1( us21_n794 ) , .ZN( us21_n795 ) );
  AOI21_X1 us21_U300 (.ZN( us21_n562 ) , .B1( us21_n722 ) , .A( us21_n777 ) , .B2( us21_n789 ) );
  NOR2_X1 us21_U301 (.ZN( us21_n576 ) , .A1( us21_n706 ) , .A2( us21_n811 ) );
  NOR2_X1 us21_U302 (.ZN( us21_n527 ) , .A1( us21_n706 ) , .A2( us21_n777 ) );
  AOI21_X1 us21_U303 (.ZN( us21_n687 ) , .B2( us21_n747 ) , .B1( us21_n761 ) , .A( us21_n804 ) );
  NOR2_X1 us21_U304 (.ZN( us21_n682 ) , .A1( us21_n789 ) , .A2( us21_n811 ) );
  AOI21_X1 us21_U305 (.ZN( us21_n648 ) , .A( us21_n777 ) , .B1( us21_n790 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U306 (.A2( us21_n811 ) , .A1( us21_n813 ) , .ZN( us21_n819 ) );
  AOI21_X1 us21_U307 (.A( us21_n788 ) , .B2( us21_n789 ) , .B1( us21_n790 ) , .ZN( us21_n791 ) );
  AOI21_X1 us21_U308 (.A( us21_n731 ) , .ZN( us21_n732 ) , .B2( us21_n778 ) , .B1( us21_n790 ) );
  NOR2_X1 us21_U309 (.ZN( us21_n581 ) , .A1( us21_n790 ) , .A2( us21_n815 ) );
  NOR4_X1 us21_U31 (.A4( us21_n774 ) , .A3( us21_n775 ) , .A1( us21_n776 ) , .ZN( us21_n797 ) , .A2( us21_n799 ) );
  NOR2_X1 us21_U310 (.ZN( us21_n532 ) , .A1( us21_n722 ) , .A2( us21_n786 ) );
  AOI21_X1 us21_U311 (.ZN( us21_n639 ) , .B1( us21_n678 ) , .A( us21_n789 ) , .B2( us21_n815 ) );
  NOR2_X1 us21_U312 (.ZN( us21_n709 ) , .A1( us21_n760 ) , .A2( us21_n761 ) );
  NOR2_X1 us21_U313 (.ZN( us21_n565 ) , .A1( us21_n745 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U314 (.ZN( us21_n680 ) , .A2( us21_n706 ) , .A1( us21_n815 ) );
  INV_X1 us21_U315 (.A( us21_n813 ) , .ZN( us21_n853 ) );
  AOI21_X1 us21_U316 (.ZN( us21_n440 ) , .A( us21_n697 ) , .B1( us21_n731 ) , .B2( us21_n748 ) );
  INV_X1 us21_U317 (.A( us21_n778 ) , .ZN( us21_n848 ) );
  AOI22_X1 us21_U318 (.A2( us21_n780 ) , .ZN( us21_n781 ) , .B2( us21_n829 ) , .A1( us21_n832 ) , .B1( us21_n861 ) );
  NAND2_X1 us21_U319 (.ZN( us21_n712 ) , .A1( us21_n726 ) , .A2( us21_n778 ) );
  NOR4_X1 us21_U32 (.A3( us21_n753 ) , .A2( us21_n754 ) , .A1( us21_n755 ) , .ZN( us21_n756 ) , .A4( us21_n867 ) );
  NAND2_X1 us21_U320 (.ZN( us21_n751 ) , .A1( us21_n761 ) , .A2( us21_n803 ) );
  AOI21_X1 us21_U321 (.ZN( us21_n441 ) , .B1( us21_n787 ) , .B2( us21_n789 ) , .A( us21_n812 ) );
  INV_X1 us21_U322 (.A( us21_n783 ) , .ZN( us21_n844 ) );
  AOI21_X1 us21_U323 (.ZN( us21_n495 ) , .A( us21_n777 ) , .B2( us21_n789 ) , .B1( us21_n802 ) );
  NAND2_X1 us21_U324 (.A2( us21_n760 ) , .A1( us21_n804 ) , .ZN( us21_n808 ) );
  NOR2_X1 us21_U325 (.ZN( us21_n468 ) , .A2( us21_n777 ) , .A1( us21_n813 ) );
  NOR2_X1 us21_U326 (.ZN( us21_n710 ) , .A2( us21_n722 ) , .A1( us21_n788 ) );
  NOR2_X1 us21_U327 (.ZN( us21_n482 ) , .A1( us21_n786 ) , .A2( us21_n803 ) );
  NOR2_X1 us21_U328 (.ZN( us21_n524 ) , .A1( us21_n722 ) , .A2( us21_n748 ) );
  OAI21_X1 us21_U329 (.A( us21_n729 ) , .B1( us21_n730 ) , .ZN( us21_n734 ) , .B2( us21_n803 ) );
  AOI211_X1 us21_U33 (.B( us21_n743 ) , .A( us21_n744 ) , .ZN( us21_n757 ) , .C1( us21_n830 ) , .C2( us21_n851 ) );
  OAI21_X1 us21_U330 (.ZN( us21_n729 ) , .A( us21_n831 ) , .B2( us21_n850 ) , .B1( us21_n871 ) );
  OAI21_X1 us21_U331 (.A( us21_n785 ) , .B2( us21_n786 ) , .B1( us21_n787 ) , .ZN( us21_n793 ) );
  OAI21_X1 us21_U332 (.ZN( us21_n785 ) , .A( us21_n837 ) , .B1( us21_n861 ) , .B2( us21_n871 ) );
  NAND2_X1 us21_U333 (.A1( us21_n697 ) , .A2( us21_n727 ) , .ZN( us21_n780 ) );
  NOR2_X1 us21_U334 (.ZN( us21_n516 ) , .A1( us21_n706 ) , .A2( us21_n786 ) );
  NAND2_X1 us21_U335 (.ZN( us21_n669 ) , .A1( us21_n804 ) , .A2( us21_n814 ) );
  OAI21_X1 us21_U336 (.A( us21_n696 ) , .ZN( us21_n700 ) , .B2( us21_n748 ) , .B1( us21_n802 ) );
  OAI21_X1 us21_U337 (.ZN( us21_n696 ) , .B2( us21_n831 ) , .B1( us21_n836 ) , .A( us21_n858 ) );
  NAND2_X1 us21_U338 (.A2( us21_n747 ) , .A1( us21_n784 ) , .ZN( us21_n807 ) );
  INV_X1 us21_U339 (.A( us21_n722 ) , .ZN( us21_n854 ) );
  NOR3_X1 us21_U34 (.A3( us21_n739 ) , .A2( us21_n740 ) , .A1( us21_n741 ) , .ZN( us21_n758 ) );
  INV_X1 us21_U340 (.A( us21_n815 ) , .ZN( us21_n842 ) );
  AND2_X1 us21_U341 (.ZN( us21_n730 ) , .A1( us21_n777 ) , .A2( us21_n783 ) );
  OAI222_X1 us21_U342 (.ZN( us21_n615 ) , .B1( us21_n695 ) , .C1( us21_n722 ) , .C2( us21_n745 ) , .B2( us21_n784 ) , .A2( us21_n790 ) , .A1( us21_n814 ) );
  AOI221_X1 us21_U343 (.A( us21_n762 ) , .ZN( us21_n772 ) , .C2( us21_n808 ) , .B2( us21_n833 ) , .C1( us21_n853 ) , .B1( us21_n864 ) );
  AOI21_X1 us21_U344 (.B2( us21_n761 ) , .ZN( us21_n762 ) , .A( us21_n786 ) , .B1( us21_n790 ) );
  INV_X1 us21_U345 (.A( us21_n759 ) , .ZN( us21_n833 ) );
  NAND2_X2 us21_U346 (.A2( us21_n439 ) , .A1( us21_n445 ) , .ZN( us21_n782 ) );
  NAND2_X1 us21_U347 (.A1( us21_n453 ) , .A2( us21_n469 ) , .ZN( us21_n801 ) );
  NAND2_X1 us21_U348 (.A1( us21_n452 ) , .A2( us21_n459 ) , .ZN( us21_n811 ) );
  NAND2_X1 us21_U349 (.A1( us21_n451 ) , .A2( us21_n459 ) , .ZN( us21_n742 ) );
  NOR4_X1 us21_U35 (.A4( us21_n732 ) , .A3( us21_n733 ) , .A2( us21_n734 ) , .A1( us21_n735 ) , .ZN( us21_n736 ) );
  NAND2_X1 us21_U350 (.A1( us21_n449 ) , .A2( us21_n452 ) , .ZN( us21_n812 ) );
  NAND2_X1 us21_U351 (.A1( us21_n453 ) , .A2( us21_n460 ) , .ZN( us21_n748 ) );
  NAND2_X1 us21_U352 (.A1( us21_n449 ) , .A2( us21_n469 ) , .ZN( us21_n814 ) );
  NAND2_X1 us21_U353 (.A1( us21_n450 ) , .A2( us21_n463 ) , .ZN( us21_n667 ) );
  NAND2_X1 us21_U354 (.A2( us21_n446 ) , .A1( us21_n458 ) , .ZN( us21_n726 ) );
  NAND2_X1 us21_U355 (.A1( us21_n451 ) , .A2( us21_n470 ) , .ZN( us21_n783 ) );
  NAND2_X1 us21_U356 (.A2( us21_n452 ) , .A1( us21_n470 ) , .ZN( us21_n777 ) );
  NAND2_X1 us21_U357 (.A2( us21_n451 ) , .A1( us21_n453 ) , .ZN( us21_n804 ) );
  NAND2_X1 us21_U358 (.A2( us21_n462 ) , .A1( us21_n463 ) , .ZN( us21_n810 ) );
  NAND2_X1 us21_U359 (.A1( us21_n439 ) , .A2( us21_n458 ) , .ZN( us21_n697 ) );
  AOI211_X1 us21_U36 (.B( us21_n723 ) , .A( us21_n724 ) , .ZN( us21_n737 ) , .C1( us21_n841 ) , .C2( us21_n853 ) );
  NAND2_X1 us21_U360 (.A2( us21_n447 ) , .A1( us21_n450 ) , .ZN( us21_n761 ) );
  NAND2_X1 us21_U361 (.A2( us21_n446 ) , .A1( us21_n450 ) , .ZN( us21_n727 ) );
  NOR2_X1 us21_U362 (.ZN( us21_n445 ) , .A2( us21_n847 ) , .A1( us21_n856 ) );
  NAND2_X1 us21_U363 (.A1( us21_n460 ) , .A2( us21_n470 ) , .ZN( us21_n786 ) );
  NOR2_X1 us21_U364 (.ZN( us21_n463 ) , .A2( us21_n845 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U365 (.ZN( us21_n451 ) , .A1( us21_n824 ) , .A2( us21_n825 ) );
  NAND2_X1 us21_U366 (.A2( us21_n459 ) , .A1( us21_n460 ) , .ZN( us21_n745 ) );
  NOR2_X1 us21_U367 (.ZN( us21_n449 ) , .A1( us21_n826 ) , .A2( us21_n827 ) );
  NAND2_X1 us21_U368 (.A2( us21_n459 ) , .A1( us21_n469 ) , .ZN( us21_n695 ) );
  NAND2_X1 us21_U369 (.A2( us21_n452 ) , .A1( us21_n453 ) , .ZN( us21_n728 ) );
  NOR3_X1 us21_U37 (.A3( us21_n720 ) , .A1( us21_n721 ) , .ZN( us21_n738 ) , .A2( us21_n739 ) );
  NAND2_X1 us21_U370 (.A1( us21_n449 ) , .A2( us21_n460 ) , .ZN( us21_n788 ) );
  NAND2_X2 us21_U371 (.A2( us21_n446 ) , .A1( us21_n462 ) , .ZN( us21_n813 ) );
  NAND2_X2 us21_U372 (.A2( us21_n439 ) , .A1( us21_n450 ) , .ZN( us21_n789 ) );
  NAND2_X2 us21_U373 (.A1( us21_n447 ) , .A2( us21_n458 ) , .ZN( us21_n790 ) );
  NAND2_X2 us21_U374 (.A1( us21_n439 ) , .A2( us21_n462 ) , .ZN( us21_n706 ) );
  NAND2_X2 us21_U375 (.A2( us21_n469 ) , .A1( us21_n470 ) , .ZN( us21_n815 ) );
  NAND2_X2 us21_U376 (.A1( us21_n445 ) , .A2( us21_n446 ) , .ZN( us21_n784 ) );
  NOR2_X1 us21_U377 (.A2( sa21_6 ) , .A1( sa21_7 ) , .ZN( us21_n462 ) );
  NOR2_X1 us21_U378 (.A2( sa21_4 ) , .ZN( us21_n447 ) , .A1( us21_n846 ) );
  NOR2_X1 us21_U379 (.A2( sa21_5 ) , .ZN( us21_n446 ) , .A1( us21_n845 ) );
  NAND4_X1 us21_U38 (.ZN( sa23_sr_3 ) , .A4( us21_n702 ) , .A3( us21_n703 ) , .A2( us21_n704 ) , .A1( us21_n705 ) );
  NOR2_X1 us21_U380 (.A2( sa21_7 ) , .ZN( us21_n458 ) , .A1( us21_n847 ) );
  NOR2_X1 us21_U381 (.A2( sa21_4 ) , .A1( sa21_5 ) , .ZN( us21_n439 ) );
  NOR2_X1 us21_U382 (.A2( sa21_1 ) , .ZN( us21_n469 ) , .A1( us21_n824 ) );
  NOR2_X1 us21_U383 (.A2( sa21_2 ) , .A1( sa21_3 ) , .ZN( us21_n470 ) );
  NOR2_X1 us21_U384 (.A2( sa21_6 ) , .ZN( us21_n450 ) , .A1( us21_n856 ) );
  NOR2_X1 us21_U385 (.A2( sa21_2 ) , .ZN( us21_n459 ) , .A1( us21_n827 ) );
  NOR2_X1 us21_U386 (.A2( sa21_0 ) , .ZN( us21_n452 ) , .A1( us21_n825 ) );
  NOR2_X1 us21_U387 (.A2( sa21_0 ) , .A1( sa21_1 ) , .ZN( us21_n460 ) );
  NOR2_X1 us21_U388 (.A2( sa21_3 ) , .ZN( us21_n453 ) , .A1( us21_n826 ) );
  INV_X1 us21_U389 (.A( sa21_6 ) , .ZN( us21_n847 ) );
  NOR4_X1 us21_U39 (.A4( us21_n698 ) , .A3( us21_n699 ) , .A2( us21_n700 ) , .A1( us21_n701 ) , .ZN( us21_n702 ) );
  INV_X1 us21_U390 (.A( sa21_3 ) , .ZN( us21_n827 ) );
  INV_X1 us21_U391 (.A( sa21_1 ) , .ZN( us21_n825 ) );
  INV_X1 us21_U392 (.A( sa21_0 ) , .ZN( us21_n824 ) );
  INV_X1 us21_U393 (.A( sa21_2 ) , .ZN( us21_n826 ) );
  INV_X1 us21_U394 (.A( sa21_5 ) , .ZN( us21_n846 ) );
  INV_X1 us21_U395 (.A( sa21_7 ) , .ZN( us21_n856 ) );
  INV_X1 us21_U396 (.A( us21_n784 ) , .ZN( us21_n860 ) );
  AOI21_X1 us21_U397 (.ZN( us21_n498 ) , .A( us21_n695 ) , .B1( us21_n706 ) , .B2( us21_n784 ) );
  INV_X1 us21_U398 (.A( us21_n695 ) , .ZN( us21_n836 ) );
  NOR2_X1 us21_U399 (.A1( us21_n695 ) , .ZN( us21_n768 ) , .A2( us21_n813 ) );
  NAND2_X1 us21_U4 (.A1( us21_n447 ) , .A2( us21_n462 ) , .ZN( us21_n722 ) );
  AOI211_X1 us21_U40 (.B( us21_n692 ) , .A( us21_n693 ) , .ZN( us21_n703 ) , .C2( us21_n829 ) , .C1( us21_n849 ) );
  AOI21_X1 us21_U400 (.ZN( us21_n569 ) , .B2( us21_n695 ) , .B1( us21_n804 ) , .A( us21_n810 ) );
  NOR2_X1 us21_U401 (.ZN( us21_n630 ) , .A2( us21_n695 ) , .A1( us21_n722 ) );
  AOI21_X1 us21_U402 (.ZN( us21_n476 ) , .B2( us21_n695 ) , .A( us21_n747 ) , .B1( us21_n777 ) );
  NOR2_X1 us21_U403 (.ZN( us21_n660 ) , .A2( us21_n695 ) , .A1( us21_n727 ) );
  NOR2_X1 us21_U404 (.A2( us21_n695 ) , .A1( us21_n778 ) , .ZN( us21_n818 ) );
  NOR2_X1 us21_U405 (.A2( us21_n695 ) , .ZN( us21_n714 ) , .A1( us21_n790 ) );
  NOR2_X1 us21_U406 (.ZN( us21_n564 ) , .A2( us21_n695 ) , .A1( us21_n761 ) );
  NOR2_X1 us21_U407 (.ZN( us21_n592 ) , .A2( us21_n695 ) , .A1( us21_n726 ) );
  AOI21_X1 us21_U408 (.ZN( us21_n550 ) , .B1( us21_n667 ) , .A( us21_n695 ) , .B2( us21_n803 ) );
  NOR2_X1 us21_U409 (.ZN( us21_n539 ) , .A2( us21_n695 ) , .A1( us21_n697 ) );
  NOR2_X1 us21_U41 (.ZN( us21_n705 ) , .A2( us21_n774 ) , .A1( us21_n798 ) );
  NOR2_X1 us21_U410 (.ZN( us21_n578 ) , .A2( us21_n695 ) , .A1( us21_n789 ) );
  OAI222_X1 us21_U411 (.B2( us21_n745 ) , .B1( us21_n746 ) , .A2( us21_n747 ) , .ZN( us21_n755 ) , .C2( us21_n803 ) , .C1( us21_n812 ) , .A1( us21_n815 ) );
  OAI222_X1 us21_U412 (.ZN( us21_n503 ) , .C2( us21_n623 ) , .B2( us21_n645 ) , .B1( us21_n745 ) , .A2( us21_n746 ) , .C1( us21_n803 ) , .A1( us21_n804 ) );
  AOI222_X1 us21_U413 (.ZN( us21_n511 ) , .C1( us21_n830 ) , .B2( us21_n835 ) , .A2( us21_n841 ) , .C2( us21_n860 ) , .B1( us21_n861 ) , .A1( us21_n864 ) );
  AOI222_X1 us21_U414 (.ZN( us21_n603 ) , .B2( us21_n669 ) , .B1( us21_n751 ) , .C2( us21_n829 ) , .A1( us21_n831 ) , .A2( us21_n860 ) , .C1( us21_n861 ) );
  AOI221_X1 us21_U415 (.A( us21_n481 ) , .ZN( us21_n486 ) , .B1( us21_n829 ) , .C2( us21_n842 ) , .C1( us21_n850 ) , .B2( us21_n860 ) );
  NOR2_X1 us21_U416 (.ZN( us21_n787 ) , .A2( us21_n860 ) , .A1( us21_n866 ) );
  OAI221_X1 us21_U417 (.A( us21_n781 ) , .C2( us21_n782 ) , .B2( us21_n783 ) , .B1( us21_n784 ) , .ZN( us21_n794 ) , .C1( us21_n811 ) );
  NAND2_X1 us21_U418 (.A1( us21_n727 ) , .A2( us21_n782 ) , .ZN( us21_n809 ) );
  OAI22_X1 us21_U419 (.ZN( us21_n586 ) , .A2( us21_n745 ) , .B2( us21_n760 ) , .A1( us21_n761 ) , .B1( us21_n782 ) );
  NOR2_X1 us21_U42 (.ZN( us21_n802 ) , .A1( us21_n852 ) , .A2( us21_n859 ) );
  OAI221_X1 us21_U420 (.A( us21_n694 ) , .ZN( us21_n701 ) , .C2( us21_n782 ) , .C1( us21_n783 ) , .B1( us21_n784 ) , .B2( us21_n804 ) );
  AOI21_X1 us21_U421 (.ZN( us21_n590 ) , .B1( us21_n726 ) , .B2( us21_n782 ) , .A( us21_n788 ) );
  AOI21_X1 us21_U422 (.ZN( us21_n646 ) , .A( us21_n760 ) , .B2( us21_n782 ) , .B1( us21_n790 ) );
  AOI21_X1 us21_U423 (.ZN( us21_n621 ) , .B1( us21_n697 ) , .A( us21_n777 ) , .B2( us21_n782 ) );
  OAI22_X1 us21_U424 (.ZN( us21_n679 ) , .A1( us21_n697 ) , .A2( us21_n728 ) , .B2( us21_n782 ) , .B1( us21_n815 ) );
  OAI21_X1 us21_U425 (.A( us21_n611 ) , .ZN( us21_n614 ) , .B1( us21_n623 ) , .B2( us21_n782 ) );
  NOR2_X1 us21_U426 (.ZN( us21_n608 ) , .A1( us21_n782 ) , .A2( us21_n814 ) );
  OAI222_X1 us21_U427 (.A2( us21_n667 ) , .ZN( us21_n672 ) , .B1( us21_n745 ) , .B2( us21_n782 ) , .C2( us21_n786 ) , .C1( us21_n813 ) , .A1( us21_n815 ) );
  NOR2_X1 us21_U428 (.ZN( us21_n649 ) , .A1( us21_n782 ) , .A2( us21_n786 ) );
  NOR2_X1 us21_U429 (.ZN( us21_n598 ) , .A2( us21_n695 ) , .A1( us21_n782 ) );
  NAND4_X1 us21_U43 (.ZN( sa23_sr_2 ) , .A4( us21_n641 ) , .A3( us21_n642 ) , .A2( us21_n643 ) , .A1( us21_n644 ) );
  NOR2_X1 us21_U430 (.ZN( us21_n551 ) , .A2( us21_n742 ) , .A1( us21_n782 ) );
  INV_X1 us21_U431 (.A( us21_n782 ) , .ZN( us21_n859 ) );
  AOI221_X1 us21_U432 (.A( us21_n574 ) , .ZN( us21_n585 ) , .B2( us21_n829 ) , .C2( us21_n841 ) , .B1( us21_n852 ) , .C1( us21_n859 ) );
  AOI21_X1 us21_U433 (.ZN( us21_n574 ) , .B2( us21_n722 ) , .B1( us21_n746 ) , .A( us21_n783 ) );
  INV_X1 us21_U434 (.A( sa21_4 ) , .ZN( us21_n845 ) );
  AOI211_X1 us21_U435 (.A( us21_n635 ) , .ZN( us21_n643 ) , .B( us21_n741 ) , .C2( us21_n837 ) , .C1( us21_n852 ) );
  NAND4_X1 us21_U436 (.A4( us21_n631 ) , .A3( us21_n632 ) , .A2( us21_n633 ) , .A1( us21_n634 ) , .ZN( us21_n741 ) );
  NAND3_X1 us21_U437 (.ZN( sa23_sr_6 ) , .A3( us21_n795 ) , .A2( us21_n796 ) , .A1( us21_n797 ) );
  NAND3_X1 us21_U438 (.ZN( sa23_sr_5 ) , .A3( us21_n756 ) , .A2( us21_n757 ) , .A1( us21_n758 ) );
  NAND3_X1 us21_U439 (.ZN( sa23_sr_4 ) , .A3( us21_n736 ) , .A2( us21_n737 ) , .A1( us21_n738 ) );
  AOI222_X1 us21_U44 (.B2( us21_n636 ) , .ZN( us21_n642 ) , .B1( us21_n839 ) , .A1( us21_n840 ) , .C2( us21_n844 ) , .C1( us21_n861 ) , .A2( us21_n863 ) );
  NAND3_X1 us21_U440 (.A3( us21_n673 ) , .A2( us21_n674 ) , .A1( us21_n675 ) , .ZN( us21_n805 ) );
  NAND3_X1 us21_U441 (.ZN( us21_n636 ) , .A3( us21_n706 ) , .A2( us21_n722 ) , .A1( us21_n790 ) );
  NAND3_X1 us21_U442 (.A3( us21_n616 ) , .A2( us21_n617 ) , .A1( us21_n618 ) , .ZN( us21_n723 ) );
  NAND3_X1 us21_U443 (.A3( us21_n583 ) , .A2( us21_n584 ) , .A1( us21_n585 ) , .ZN( us21_n619 ) );
  NAND3_X1 us21_U444 (.ZN( us21_n563 ) , .A3( us21_n678 ) , .A2( us21_n748 ) , .A1( us21_n783 ) );
  NAND3_X1 us21_U445 (.A3( us21_n521 ) , .A2( us21_n522 ) , .A1( us21_n523 ) , .ZN( us21_n740 ) );
  NAND3_X1 us21_U446 (.A3( us21_n510 ) , .A1( us21_n511 ) , .ZN( us21_n606 ) , .A2( us21_n869 ) );
  NAND3_X1 us21_U447 (.A3( us21_n465 ) , .A2( us21_n466 ) , .A1( us21_n467 ) , .ZN( us21_n775 ) );
  NOR4_X1 us21_U45 (.A4( us21_n637 ) , .A3( us21_n638 ) , .A2( us21_n639 ) , .A1( us21_n640 ) , .ZN( us21_n641 ) );
  NOR3_X1 us21_U46 (.A2( us21_n605 ) , .A1( us21_n606 ) , .ZN( us21_n644 ) , .A3( us21_n720 ) );
  NAND4_X1 us21_U47 (.ZN( sa23_sr_0 ) , .A4( us21_n499 ) , .A3( us21_n500 ) , .A2( us21_n501 ) , .A1( us21_n502 ) );
  NOR4_X1 us21_U48 (.A4( us21_n496 ) , .A3( us21_n497 ) , .A2( us21_n498 ) , .ZN( us21_n499 ) , .A1( us21_n525 ) );
  AOI221_X1 us21_U49 (.A( us21_n495 ) , .ZN( us21_n500 ) , .B2( us21_n841 ) , .C1( us21_n844 ) , .C2( us21_n858 ) , .B1( us21_n860 ) );
  NAND2_X1 us21_U5 (.A1( us21_n445 ) , .A2( us21_n447 ) , .ZN( us21_n803 ) );
  AOI211_X1 us21_U50 (.A( us21_n494 ) , .ZN( us21_n501 ) , .B( us21_n800 ) , .C2( us21_n837 ) , .C1( us21_n849 ) );
  NAND4_X1 us21_U51 (.ZN( sa23_sr_1 ) , .A4( us21_n593 ) , .A3( us21_n594 ) , .A2( us21_n595 ) , .A1( us21_n596 ) );
  AOI211_X1 us21_U52 (.B( us21_n587 ) , .A( us21_n588 ) , .ZN( us21_n594 ) , .C2( us21_n809 ) , .C1( us21_n831 ) );
  NOR4_X1 us21_U53 (.A4( us21_n589 ) , .A3( us21_n590 ) , .A2( us21_n591 ) , .A1( us21_n592 ) , .ZN( us21_n593 ) );
  AOI211_X1 us21_U54 (.A( us21_n586 ) , .ZN( us21_n595 ) , .B( us21_n619 ) , .C1( us21_n843 ) , .C2( us21_n853 ) );
  NAND4_X1 us21_U55 (.A4( us21_n601 ) , .A3( us21_n602 ) , .A2( us21_n603 ) , .A1( us21_n604 ) , .ZN( us21_n720 ) );
  NOR3_X1 us21_U56 (.A1( us21_n597 ) , .ZN( us21_n602 ) , .A3( us21_n661 ) , .A2( us21_n768 ) );
  NOR4_X1 us21_U57 (.A3( us21_n598 ) , .A2( us21_n599 ) , .A1( us21_n600 ) , .ZN( us21_n601 ) , .A4( us21_n653 ) );
  AOI222_X1 us21_U58 (.ZN( us21_n604 ) , .A1( us21_n828 ) , .C2( us21_n835 ) , .B1( us21_n840 ) , .A2( us21_n854 ) , .B2( us21_n859 ) , .C1( us21_n866 ) );
  AOI222_X1 us21_U59 (.ZN( us21_n467 ) , .B1( us21_n830 ) , .A1( us21_n837 ) , .C1( us21_n840 ) , .C2( us21_n849 ) , .A2( us21_n853 ) , .B2( us21_n863 ) );
  NOR3_X1 us21_U6 (.ZN( us21_n596 ) , .A1( us21_n606 ) , .A3( us21_n721 ) , .A2( us21_n740 ) );
  NOR4_X1 us21_U60 (.A1( us21_n464 ) , .ZN( us21_n465 ) , .A4( us21_n540 ) , .A2( us21_n552 ) , .A3( us21_n612 ) );
  AOI221_X1 us21_U61 (.ZN( us21_n466 ) , .C2( us21_n712 ) , .B2( us21_n829 ) , .C1( us21_n843 ) , .B1( us21_n858 ) , .A( us21_n862 ) );
  NAND4_X1 us21_U62 (.A4( us21_n483 ) , .A3( us21_n484 ) , .A2( us21_n485 ) , .A1( us21_n486 ) , .ZN( us21_n776 ) );
  NOR4_X1 us21_U63 (.ZN( us21_n484 ) , .A1( us21_n505 ) , .A2( us21_n517 ) , .A4( us21_n544 ) , .A3( us21_n609 ) );
  NOR4_X1 us21_U64 (.A4( us21_n482 ) , .ZN( us21_n485 ) , .A1( us21_n564 ) , .A2( us21_n579 ) , .A3( us21_n600 ) );
  NOR4_X1 us21_U65 (.ZN( us21_n483 ) , .A2( us21_n531 ) , .A1( us21_n556 ) , .A3( us21_n629 ) , .A4( us21_n716 ) );
  AOI211_X1 us21_U66 (.B( us21_n621 ) , .A( us21_n622 ) , .ZN( us21_n633 ) , .C2( us21_n834 ) , .C1( us21_n861 ) );
  NOR4_X1 us21_U67 (.A4( us21_n627 ) , .A3( us21_n628 ) , .A2( us21_n629 ) , .A1( us21_n630 ) , .ZN( us21_n631 ) );
  NOR4_X1 us21_U68 (.A4( us21_n624 ) , .A3( us21_n625 ) , .A2( us21_n626 ) , .ZN( us21_n632 ) , .A1( us21_n662 ) );
  NOR4_X1 us21_U69 (.A4( us21_n512 ) , .A3( us21_n513 ) , .A2( us21_n514 ) , .A1( us21_n515 ) , .ZN( us21_n522 ) );
  NOR3_X1 us21_U7 (.A3( us21_n798 ) , .A2( us21_n799 ) , .A1( us21_n800 ) , .ZN( us21_n823 ) );
  AOI222_X1 us21_U70 (.ZN( us21_n523 ) , .A1( us21_n832 ) , .B2( us21_n835 ) , .C1( us21_n842 ) , .C2( us21_n848 ) , .A2( us21_n850 ) , .B1( us21_n864 ) );
  NOR4_X1 us21_U71 (.A3( us21_n519 ) , .A1( us21_n520 ) , .ZN( us21_n521 ) , .A2( us21_n671 ) , .A4( us21_n767 ) );
  NAND4_X1 us21_U72 (.A4( us21_n655 ) , .A3( us21_n656 ) , .A2( us21_n657 ) , .A1( us21_n658 ) , .ZN( us21_n798 ) );
  NOR3_X1 us21_U73 (.A3( us21_n646 ) , .A2( us21_n647 ) , .A1( us21_n648 ) , .ZN( us21_n657 ) );
  NOR3_X1 us21_U74 (.A3( us21_n649 ) , .A2( us21_n650 ) , .A1( us21_n651 ) , .ZN( us21_n656 ) );
  NOR3_X1 us21_U75 (.A3( us21_n652 ) , .A2( us21_n653 ) , .A1( us21_n654 ) , .ZN( us21_n655 ) );
  NAND4_X1 us21_U76 (.A4( us21_n558 ) , .A3( us21_n559 ) , .A2( us21_n560 ) , .A1( us21_n561 ) , .ZN( us21_n605 ) );
  NOR4_X1 us21_U77 (.A4( us21_n550 ) , .A3( us21_n551 ) , .A2( us21_n552 ) , .A1( us21_n553 ) , .ZN( us21_n560 ) );
  NOR4_X1 us21_U78 (.A4( us21_n554 ) , .A3( us21_n555 ) , .A2( us21_n556 ) , .A1( us21_n557 ) , .ZN( us21_n558 ) );
  NOR4_X1 us21_U79 (.ZN( us21_n559 ) , .A1( us21_n651 ) , .A3( us21_n659 ) , .A4( us21_n683 ) , .A2( us21_n766 ) );
  NOR3_X1 us21_U8 (.ZN( us21_n502 ) , .A2( us21_n677 ) , .A3( us21_n775 ) , .A1( us21_n874 ) );
  NAND4_X1 us21_U80 (.A4( us21_n770 ) , .A3( us21_n771 ) , .A2( us21_n772 ) , .A1( us21_n773 ) , .ZN( us21_n799 ) );
  NOR3_X1 us21_U81 (.A3( us21_n763 ) , .A2( us21_n764 ) , .A1( us21_n765 ) , .ZN( us21_n771 ) );
  NOR4_X1 us21_U82 (.A4( us21_n766 ) , .A3( us21_n767 ) , .A2( us21_n768 ) , .A1( us21_n769 ) , .ZN( us21_n770 ) );
  AOI222_X1 us21_U83 (.ZN( us21_n773 ) , .A1( us21_n828 ) , .C1( us21_n832 ) , .B2( us21_n839 ) , .A2( us21_n848 ) , .B1( us21_n859 ) , .C2( us21_n871 ) );
  NOR4_X1 us21_U84 (.A4( us21_n507 ) , .A2( us21_n508 ) , .A1( us21_n509 ) , .ZN( us21_n510 ) , .A3( us21_n668 ) );
  INV_X1 us21_U85 (.A( us21_n503 ) , .ZN( us21_n869 ) );
  NOR4_X1 us21_U86 (.A4( us21_n659 ) , .A3( us21_n660 ) , .A2( us21_n661 ) , .A1( us21_n662 ) , .ZN( us21_n675 ) );
  NOR4_X1 us21_U87 (.A4( us21_n663 ) , .A3( us21_n664 ) , .A2( us21_n665 ) , .A1( us21_n666 ) , .ZN( us21_n674 ) );
  NOR4_X1 us21_U88 (.A3( us21_n671 ) , .A1( us21_n672 ) , .ZN( us21_n673 ) , .A4( us21_n713 ) , .A2( us21_n857 ) );
  NOR2_X1 us21_U89 (.ZN( us21_n623 ) , .A2( us21_n834 ) , .A1( us21_n837 ) );
  INV_X1 us21_U9 (.A( us21_n704 ) , .ZN( us21_n874 ) );
  NOR2_X1 us21_U90 (.ZN( us21_n759 ) , .A1( us21_n831 ) , .A2( us21_n832 ) );
  NAND4_X1 us21_U91 (.A4( us21_n454 ) , .A3( us21_n455 ) , .A2( us21_n456 ) , .A1( us21_n457 ) , .ZN( us21_n677 ) );
  NOR3_X1 us21_U92 (.ZN( us21_n455 ) , .A3( us21_n528 ) , .A1( us21_n553 ) , .A2( us21_n568 ) );
  AOI221_X1 us21_U93 (.A( us21_n448 ) , .ZN( us21_n457 ) , .C2( us21_n751 ) , .B1( us21_n830 ) , .C1( us21_n840 ) , .B2( us21_n859 ) );
  NOR4_X1 us21_U94 (.ZN( us21_n456 ) , .A2( us21_n507 ) , .A1( us21_n597 ) , .A4( us21_n626 ) , .A3( us21_n709 ) );
  NAND4_X1 us21_U95 (.ZN( sa23_sr_7 ) , .A4( us21_n820 ) , .A3( us21_n821 ) , .A2( us21_n822 ) , .A1( us21_n823 ) );
  NOR4_X1 us21_U96 (.A4( us21_n816 ) , .A3( us21_n817 ) , .A2( us21_n818 ) , .A1( us21_n819 ) , .ZN( us21_n820 ) );
  AOI222_X1 us21_U97 (.C2( us21_n807 ) , .B2( us21_n808 ) , .A2( us21_n809 ) , .ZN( us21_n821 ) , .C1( us21_n830 ) , .A1( us21_n837 ) , .B1( us21_n851 ) );
  AOI211_X1 us21_U98 (.B( us21_n805 ) , .A( us21_n806 ) , .ZN( us21_n822 ) , .C1( us21_n840 ) , .C2( us21_n848 ) );
  NAND4_X1 us21_U99 (.A4( us21_n533 ) , .A3( us21_n534 ) , .A2( us21_n535 ) , .A1( us21_n536 ) , .ZN( us21_n620 ) );
  NOR2_X1 us22_U10 (.ZN( us22_n573 ) , .A1( us22_n620 ) , .A2( us22_n743 ) );
  NOR4_X1 us22_U100 (.A4( us22_n527 ) , .A3( us22_n528 ) , .ZN( us22_n535 ) , .A2( us22_n682 ) , .A1( us22_n792 ) );
  NAND4_X1 us22_U101 (.A4( us22_n477 ) , .A3( us22_n478 ) , .A2( us22_n479 ) , .A1( us22_n480 ) , .ZN( us22_n692 ) );
  NOR3_X1 us22_U102 (.ZN( us22_n478 ) , .A2( us22_n506 ) , .A3( us22_n599 ) , .A1( us22_n608 ) );
  AOI211_X1 us22_U103 (.B( us22_n475 ) , .A( us22_n476 ) , .ZN( us22_n480 ) , .C2( us22_n831 ) , .C1( us22_n859 ) );
  NOR4_X1 us22_U104 (.ZN( us22_n479 ) , .A3( us22_n530 ) , .A4( us22_n543 ) , .A2( us22_n565 ) , .A1( us22_n715 ) );
  NAND4_X1 us22_U105 (.A4( us22_n546 ) , .A3( us22_n547 ) , .A2( us22_n548 ) , .A1( us22_n549 ) , .ZN( us22_n743 ) );
  NOR3_X1 us22_U106 (.ZN( us22_n547 ) , .A2( us22_n649 ) , .A1( us22_n665 ) , .A3( us22_n769 ) );
  AOI211_X1 us22_U107 (.B( us22_n537 ) , .A( us22_n538 ) , .ZN( us22_n549 ) , .C2( us22_n837 ) , .C1( us22_n849 ) );
  NOR4_X1 us22_U108 (.A4( us22_n542 ) , .A3( us22_n543 ) , .A2( us22_n544 ) , .A1( us22_n545 ) , .ZN( us22_n546 ) );
  NOR2_X1 us22_U109 (.ZN( us22_n684 ) , .A1( us22_n829 ) , .A2( us22_n830 ) );
  NOR2_X1 us22_U11 (.A1( us22_n676 ) , .ZN( us22_n691 ) , .A2( us22_n805 ) );
  NOR4_X1 us22_U110 (.ZN( us22_n618 ) , .A1( us22_n654 ) , .A3( us22_n664 ) , .A4( us22_n680 ) , .A2( us22_n764 ) );
  NOR4_X1 us22_U111 (.A4( us22_n607 ) , .A3( us22_n608 ) , .A2( us22_n609 ) , .A1( us22_n610 ) , .ZN( us22_n617 ) );
  NOR4_X1 us22_U112 (.A4( us22_n612 ) , .A3( us22_n613 ) , .A2( us22_n614 ) , .A1( us22_n615 ) , .ZN( us22_n616 ) );
  NAND4_X1 us22_U113 (.A4( us22_n483 ) , .A3( us22_n484 ) , .A2( us22_n485 ) , .A1( us22_n486 ) , .ZN( us22_n776 ) );
  NOR4_X1 us22_U114 (.A4( us22_n482 ) , .ZN( us22_n485 ) , .A1( us22_n564 ) , .A2( us22_n579 ) , .A3( us22_n600 ) );
  NOR4_X1 us22_U115 (.ZN( us22_n484 ) , .A1( us22_n505 ) , .A2( us22_n517 ) , .A4( us22_n544 ) , .A3( us22_n609 ) );
  NOR4_X1 us22_U116 (.ZN( us22_n483 ) , .A2( us22_n531 ) , .A1( us22_n556 ) , .A3( us22_n629 ) , .A4( us22_n716 ) );
  NAND4_X1 us22_U117 (.A4( us22_n689 ) , .A3( us22_n690 ) , .A1( us22_n691 ) , .ZN( us22_n774 ) , .A2( us22_n870 ) );
  AOI221_X1 us22_U118 (.A( us22_n679 ) , .ZN( us22_n690 ) , .B2( us22_n838 ) , .C1( us22_n840 ) , .C2( us22_n860 ) , .B1( us22_n863 ) );
  INV_X1 us22_U119 (.A( us22_n677 ) , .ZN( us22_n870 ) );
  INV_X1 us22_U12 (.A( us22_n678 ) , .ZN( us22_n838 ) );
  NOR4_X1 us22_U120 (.A4( us22_n685 ) , .A3( us22_n686 ) , .A2( us22_n687 ) , .A1( us22_n688 ) , .ZN( us22_n689 ) );
  NAND4_X1 us22_U121 (.A4( us22_n717 ) , .A3( us22_n718 ) , .A2( us22_n719 ) , .ZN( us22_n739 ) , .A1( us22_n855 ) );
  INV_X1 us22_U122 (.A( us22_n707 ) , .ZN( us22_n855 ) );
  AOI221_X1 us22_U123 (.A( us22_n708 ) , .ZN( us22_n719 ) , .C2( us22_n842 ) , .B2( us22_n843 ) , .C1( us22_n859 ) , .B1( us22_n860 ) );
  NOR4_X1 us22_U124 (.A4( us22_n713 ) , .A3( us22_n714 ) , .A2( us22_n715 ) , .A1( us22_n716 ) , .ZN( us22_n717 ) );
  NAND4_X1 us22_U125 (.A4( us22_n471 ) , .A3( us22_n472 ) , .A2( us22_n473 ) , .A1( us22_n474 ) , .ZN( us22_n676 ) );
  NOR4_X1 us22_U126 (.A4( us22_n468 ) , .ZN( us22_n474 ) , .A3( us22_n554 ) , .A1( us22_n733 ) , .A2( us22_n753 ) );
  NOR4_X1 us22_U127 (.ZN( us22_n473 ) , .A1( us22_n529 ) , .A3( us22_n566 ) , .A4( us22_n598 ) , .A2( us22_n640 ) );
  NOR4_X1 us22_U128 (.ZN( us22_n472 ) , .A1( us22_n504 ) , .A3( us22_n542 ) , .A2( us22_n581 ) , .A4( us22_n714 ) );
  NOR2_X1 us22_U129 (.ZN( us22_n731 ) , .A2( us22_n830 ) , .A1( us22_n843 ) );
  NOR4_X1 us22_U13 (.A4( us22_n443 ) , .A3( us22_n444 ) , .A2( us22_n514 ) , .A1( us22_n539 ) , .ZN( us22_n704 ) );
  NOR2_X1 us22_U130 (.ZN( us22_n787 ) , .A2( us22_n860 ) , .A1( us22_n866 ) );
  NOR2_X1 us22_U131 (.ZN( us22_n645 ) , .A1( us22_n852 ) , .A2( us22_n866 ) );
  NAND4_X1 us22_U132 (.A4( us22_n571 ) , .A3( us22_n572 ) , .A1( us22_n573 ) , .ZN( us22_n721 ) , .A2( us22_n872 ) );
  NOR4_X1 us22_U133 (.A4( us22_n567 ) , .A3( us22_n568 ) , .A2( us22_n569 ) , .A1( us22_n570 ) , .ZN( us22_n571 ) );
  AOI221_X1 us22_U134 (.A( us22_n562 ) , .C2( us22_n563 ) , .ZN( us22_n572 ) , .B2( us22_n843 ) , .B1( us22_n850 ) , .C1( us22_n851 ) );
  INV_X1 us22_U135 (.A( us22_n605 ) , .ZN( us22_n872 ) );
  NAND4_X1 us22_U136 (.A4( us22_n491 ) , .A3( us22_n492 ) , .A1( us22_n493 ) , .ZN( us22_n800 ) , .A2( us22_n865 ) );
  AOI221_X1 us22_U137 (.A( us22_n487 ) , .ZN( us22_n492 ) , .B2( us22_n834 ) , .C2( us22_n839 ) , .C1( us22_n849 ) , .B1( us22_n858 ) );
  INV_X1 us22_U138 (.A( us22_n776 ) , .ZN( us22_n865 ) );
  NOR2_X1 us22_U139 (.ZN( us22_n493 ) , .A1( us22_n676 ) , .A2( us22_n692 ) );
  OR3_X1 us22_U14 (.ZN( us22_n444 ) , .A1( us22_n526 ) , .A3( us22_n575 ) , .A2( us22_n873 ) );
  INV_X1 us22_U140 (.A( us22_n760 ) , .ZN( us22_n828 ) );
  INV_X1 us22_U141 (.A( us22_n461 ) , .ZN( us22_n862 ) );
  OAI21_X1 us22_U142 (.ZN( us22_n461 ) , .B1( us22_n807 ) , .A( us22_n832 ) , .B2( us22_n849 ) );
  OR4_X1 us22_U143 (.A4( us22_n578 ) , .A3( us22_n579 ) , .A2( us22_n580 ) , .A1( us22_n581 ) , .ZN( us22_n582 ) );
  OR4_X1 us22_U144 (.A4( us22_n680 ) , .A3( us22_n681 ) , .A2( us22_n682 ) , .A1( us22_n683 ) , .ZN( us22_n688 ) );
  OR4_X1 us22_U145 (.A4( us22_n564 ) , .A3( us22_n565 ) , .A2( us22_n566 ) , .ZN( us22_n570 ) , .A1( us22_n663 ) );
  OR4_X1 us22_U146 (.A4( us22_n516 ) , .A2( us22_n517 ) , .A1( us22_n518 ) , .ZN( us22_n520 ) , .A3( us22_n819 ) );
  OR4_X1 us22_U147 (.ZN( us22_n464 ) , .A4( us22_n516 ) , .A3( us22_n527 ) , .A2( us22_n576 ) , .A1( us22_n710 ) );
  NAND2_X1 us22_U148 (.ZN( us22_n611 ) , .A2( us22_n835 ) , .A1( us22_n871 ) );
  OR3_X1 us22_U149 (.A3( us22_n504 ) , .A2( us22_n505 ) , .A1( us22_n506 ) , .ZN( us22_n509 ) );
  OR4_X1 us22_U15 (.A4( us22_n440 ) , .A2( us22_n441 ) , .A1( us22_n442 ) , .ZN( us22_n443 ) , .A3( us22_n551 ) );
  AOI221_X1 us22_U150 (.A( us22_n711 ) , .B2( us22_n712 ) , .ZN( us22_n718 ) , .C1( us22_n830 ) , .B1( us22_n837 ) , .C2( us22_n861 ) );
  OR2_X1 us22_U151 (.A2( us22_n709 ) , .A1( us22_n710 ) , .ZN( us22_n711 ) );
  INV_X1 us22_U152 (.A( us22_n752 ) , .ZN( us22_n867 ) );
  OAI21_X1 us22_U153 (.B1( us22_n751 ) , .ZN( us22_n752 ) , .A( us22_n843 ) , .B2( us22_n866 ) );
  INV_X1 us22_U154 (.A( us22_n670 ) , .ZN( us22_n857 ) );
  AOI21_X1 us22_U155 (.A( us22_n668 ) , .B1( us22_n669 ) , .ZN( us22_n670 ) , .B2( us22_n854 ) );
  NAND2_X1 us22_U156 (.A1( us22_n445 ) , .A2( us22_n463 ) , .ZN( us22_n747 ) );
  OAI222_X1 us22_U157 (.B2( us22_n745 ) , .B1( us22_n746 ) , .A2( us22_n747 ) , .ZN( us22_n755 ) , .C2( us22_n803 ) , .C1( us22_n812 ) , .A1( us22_n815 ) );
  OAI222_X1 us22_U158 (.B2( us22_n706 ) , .ZN( us22_n707 ) , .C2( us22_n722 ) , .B1( us22_n745 ) , .A1( us22_n804 ) , .C1( us22_n812 ) , .A2( us22_n813 ) );
  OAI222_X1 us22_U159 (.ZN( us22_n615 ) , .B1( us22_n695 ) , .C1( us22_n722 ) , .C2( us22_n745 ) , .B2( us22_n784 ) , .A2( us22_n790 ) , .A1( us22_n814 ) );
  INV_X1 us22_U16 (.A( us22_n611 ) , .ZN( us22_n873 ) );
  OAI222_X1 us22_U160 (.ZN( us22_n503 ) , .C2( us22_n623 ) , .B2( us22_n645 ) , .B1( us22_n745 ) , .A2( us22_n746 ) , .C1( us22_n803 ) , .A1( us22_n804 ) );
  NOR4_X1 us22_U161 (.A2( us22_n489 ) , .A1( us22_n490 ) , .ZN( us22_n491 ) , .A3( us22_n578 ) , .A4( us22_n610 ) );
  OR4_X1 us22_U162 (.ZN( us22_n490 ) , .A4( us22_n532 ) , .A2( us22_n545 ) , .A1( us22_n557 ) , .A3( us22_n630 ) );
  OAI22_X1 us22_U163 (.B1( us22_n488 ) , .ZN( us22_n489 ) , .A1( us22_n684 ) , .A2( us22_n761 ) , .B2( us22_n815 ) );
  NOR3_X1 us22_U164 (.ZN( us22_n488 ) , .A1( us22_n780 ) , .A2( us22_n848 ) , .A3( us22_n861 ) );
  AOI22_X1 us22_U165 (.ZN( us22_n694 ) , .A1( us22_n828 ) , .B2( us22_n841 ) , .A2( us22_n863 ) , .B1( us22_n866 ) );
  AOI22_X1 us22_U166 (.A2( us22_n780 ) , .ZN( us22_n781 ) , .B2( us22_n829 ) , .A1( us22_n832 ) , .B1( us22_n861 ) );
  INV_X1 us22_U167 (.A( us22_n728 ) , .ZN( us22_n837 ) );
  AOI221_X1 us22_U168 (.A( us22_n481 ) , .ZN( us22_n486 ) , .B1( us22_n829 ) , .C2( us22_n842 ) , .C1( us22_n850 ) , .B2( us22_n860 ) );
  OAI22_X1 us22_U169 (.ZN( us22_n481 ) , .A1( us22_n706 ) , .B2( us22_n783 ) , .A2( us22_n804 ) , .B1( us22_n810 ) );
  INV_X1 us22_U17 (.A( us22_n747 ) , .ZN( us22_n861 ) );
  INV_X1 us22_U170 (.A( us22_n788 ) , .ZN( us22_n830 ) );
  NAND2_X1 us22_U171 (.A1( us22_n449 ) , .A2( us22_n451 ) , .ZN( us22_n760 ) );
  OAI22_X1 us22_U172 (.ZN( us22_n635 ) , .A1( us22_n697 ) , .B2( us22_n726 ) , .A2( us22_n760 ) , .B1( us22_n814 ) );
  OAI221_X1 us22_U173 (.A( us22_n725 ) , .C2( us22_n726 ) , .B2( us22_n727 ) , .B1( us22_n728 ) , .ZN( us22_n735 ) , .C1( us22_n815 ) );
  AOI22_X1 us22_U174 (.ZN( us22_n725 ) , .B1( us22_n830 ) , .A2( us22_n836 ) , .A1( us22_n861 ) , .B2( us22_n864 ) );
  OAI22_X1 us22_U175 (.ZN( us22_n708 ) , .A2( us22_n726 ) , .B2( us22_n727 ) , .A1( us22_n742 ) , .B1( us22_n811 ) );
  INV_X1 us22_U176 (.A( us22_n814 ) , .ZN( us22_n829 ) );
  OAI22_X1 us22_U177 (.ZN( us22_n487 ) , .A1( us22_n722 ) , .B2( us22_n726 ) , .B1( us22_n728 ) , .A2( us22_n777 ) );
  OAI22_X1 us22_U178 (.ZN( us22_n622 ) , .B1( us22_n667 ) , .B2( us22_n745 ) , .A1( us22_n813 ) , .A2( us22_n814 ) );
  INV_X1 us22_U179 (.A( us22_n742 ) , .ZN( us22_n835 ) );
  AOI222_X1 us22_U18 (.ZN( us22_n603 ) , .B2( us22_n669 ) , .B1( us22_n751 ) , .C2( us22_n829 ) , .A1( us22_n831 ) , .A2( us22_n860 ) , .C1( us22_n861 ) );
  OAI22_X1 us22_U180 (.A1( us22_n722 ) , .ZN( us22_n724 ) , .B2( us22_n748 ) , .B1( us22_n810 ) , .A2( us22_n814 ) );
  OAI22_X1 us22_U181 (.B2( us22_n777 ) , .B1( us22_n778 ) , .ZN( us22_n779 ) , .A2( us22_n812 ) , .A1( us22_n813 ) );
  INV_X1 us22_U182 (.A( us22_n786 ) , .ZN( us22_n843 ) );
  INV_X1 us22_U183 (.A( us22_n812 ) , .ZN( us22_n831 ) );
  OAI22_X1 us22_U184 (.B2( us22_n742 ) , .ZN( us22_n744 ) , .A2( us22_n760 ) , .B1( us22_n778 ) , .A1( us22_n790 ) );
  OAI22_X1 us22_U185 (.B2( us22_n801 ) , .B1( us22_n802 ) , .A2( us22_n803 ) , .A1( us22_n804 ) , .ZN( us22_n806 ) );
  INV_X1 us22_U186 (.A( us22_n667 ) , .ZN( us22_n863 ) );
  OAI22_X1 us22_U187 (.ZN( us22_n494 ) , .A2( us22_n742 ) , .A1( us22_n778 ) , .B1( us22_n789 ) , .B2( us22_n804 ) );
  INV_X1 us22_U188 (.A( us22_n748 ) , .ZN( us22_n840 ) );
  OAI22_X1 us22_U189 (.ZN( us22_n588 ) , .B1( us22_n728 ) , .B2( us22_n747 ) , .A2( us22_n784 ) , .A1( us22_n801 ) );
  AOI222_X1 us22_U19 (.ZN( us22_n561 ) , .B1( us22_n828 ) , .C1( us22_n839 ) , .A2( us22_n841 ) , .A1( us22_n852 ) , .B2( us22_n861 ) , .C2( us22_n871 ) );
  OAI22_X1 us22_U190 (.ZN( us22_n693 ) , .A2( us22_n728 ) , .A1( us22_n778 ) , .B1( us22_n789 ) , .B2( us22_n815 ) );
  INV_X1 us22_U191 (.A( us22_n801 ) , .ZN( us22_n841 ) );
  NOR2_X1 us22_U192 (.A1( us22_n695 ) , .ZN( us22_n768 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U193 (.ZN( us22_n664 ) , .A1( us22_n726 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U194 (.ZN( us22_n592 ) , .A2( us22_n695 ) , .A1( us22_n726 ) );
  NOR2_X1 us22_U195 (.ZN( us22_n568 ) , .A1( us22_n726 ) , .A2( us22_n804 ) );
  NOR2_X1 us22_U196 (.ZN( us22_n716 ) , .A2( us22_n722 ) , .A1( us22_n742 ) );
  NOR2_X1 us22_U197 (.ZN( us22_n544 ) , .A2( us22_n778 ) , .A1( us22_n812 ) );
  NOR2_X1 us22_U198 (.ZN( us22_n575 ) , .A2( us22_n697 ) , .A1( us22_n812 ) );
  NOR2_X1 us22_U199 (.ZN( us22_n652 ) , .A1( us22_n726 ) , .A2( us22_n811 ) );
  AOI222_X1 us22_U20 (.ZN( us22_n658 ) , .A2( us22_n837 ) , .B1( us22_n839 ) , .C2( us22_n843 ) , .A1( us22_n858 ) , .C1( us22_n861 ) , .B2( us22_n868 ) );
  NOR2_X1 us22_U200 (.ZN( us22_n610 ) , .A1( us22_n777 ) , .A2( us22_n784 ) );
  NOR2_X1 us22_U201 (.ZN( us22_n530 ) , .A2( us22_n747 ) , .A1( us22_n748 ) );
  NOR2_X1 us22_U202 (.ZN( us22_n627 ) , .A2( us22_n726 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U203 (.ZN( us22_n613 ) , .A1( us22_n783 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U204 (.ZN( us22_n599 ) , .A2( us22_n778 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U205 (.ZN( us22_n609 ) , .A2( us22_n778 ) , .A1( us22_n804 ) );
  INV_X1 us22_U206 (.A( us22_n745 ) , .ZN( us22_n832 ) );
  NOR2_X1 us22_U207 (.A2( us22_n742 ) , .ZN( us22_n767 ) , .A1( us22_n810 ) );
  NOR2_X1 us22_U208 (.ZN( us22_n526 ) , .A2( us22_n722 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U209 (.ZN( us22_n529 ) , .A2( us22_n778 ) , .A1( us22_n814 ) );
  INV_X1 us22_U21 (.A( us22_n645 ) , .ZN( us22_n868 ) );
  NOR2_X1 us22_U210 (.ZN( us22_n626 ) , .A2( us22_n667 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U211 (.ZN( us22_n597 ) , .A2( us22_n789 ) , .A1( us22_n814 ) );
  INV_X1 us22_U212 (.A( us22_n790 ) , .ZN( us22_n849 ) );
  INV_X1 us22_U213 (.A( us22_n726 ) , .ZN( us22_n850 ) );
  NOR2_X1 us22_U214 (.ZN( us22_n650 ) , .A1( us22_n667 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U215 (.A1( us22_n667 ) , .ZN( us22_n671 ) , .A2( us22_n742 ) );
  INV_X1 us22_U216 (.A( us22_n803 ) , .ZN( us22_n858 ) );
  NOR2_X1 us22_U217 (.ZN( us22_n600 ) , .A1( us22_n667 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U218 (.A1( us22_n667 ) , .ZN( us22_n686 ) , .A2( us22_n814 ) );
  NOR2_X1 us22_U219 (.A2( us22_n706 ) , .A1( us22_n748 ) , .ZN( us22_n769 ) );
  NOR4_X1 us22_U22 (.ZN( us22_n471 ) , .A2( us22_n519 ) , .A4( us22_n592 ) , .A1( us22_n607 ) , .A3( us22_n627 ) );
  NOR2_X1 us22_U220 (.A1( us22_n667 ) , .ZN( us22_n764 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U221 (.A1( us22_n697 ) , .ZN( us22_n766 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U222 (.ZN( us22_n539 ) , .A2( us22_n695 ) , .A1( us22_n697 ) );
  NOR2_X1 us22_U223 (.ZN( us22_n525 ) , .A1( us22_n667 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U224 (.ZN( us22_n665 ) , .A1( us22_n748 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U225 (.ZN( us22_n553 ) , .A1( us22_n748 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U226 (.ZN( us22_n506 ) , .A2( us22_n778 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U227 (.ZN( us22_n541 ) , .A2( us22_n706 ) , .A1( us22_n783 ) );
  NOR2_X1 us22_U228 (.ZN( us22_n662 ) , .A1( us22_n783 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U229 (.A2( us22_n695 ) , .ZN( us22_n714 ) , .A1( us22_n790 ) );
  NOR4_X1 us22_U23 (.ZN( us22_n477 ) , .A1( us22_n518 ) , .A4( us22_n555 ) , .A3( us22_n580 ) , .A2( us22_n628 ) );
  NOR2_X1 us22_U230 (.ZN( us22_n505 ) , .A1( us22_n810 ) , .A2( us22_n815 ) );
  INV_X1 us22_U231 (.A( us22_n804 ) , .ZN( us22_n839 ) );
  NOR2_X1 us22_U232 (.ZN( us22_n659 ) , .A1( us22_n727 ) , .A2( us22_n788 ) );
  NOR2_X1 us22_U233 (.ZN( us22_n660 ) , .A2( us22_n695 ) , .A1( us22_n727 ) );
  NOR2_X1 us22_U234 (.ZN( us22_n555 ) , .A1( us22_n790 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U235 (.ZN( us22_n543 ) , .A1( us22_n747 ) , .A2( us22_n812 ) );
  NOR2_X1 us22_U236 (.ZN( us22_n507 ) , .A1( us22_n727 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U237 (.A2( us22_n695 ) , .A1( us22_n778 ) , .ZN( us22_n818 ) );
  OAI22_X1 us22_U238 (.B2( us22_n748 ) , .B1( us22_n749 ) , .A1( us22_n750 ) , .ZN( us22_n754 ) , .A2( us22_n804 ) );
  NOR2_X1 us22_U239 (.ZN( us22_n749 ) , .A2( us22_n850 ) , .A1( us22_n858 ) );
  NOR4_X1 us22_U24 (.ZN( us22_n454 ) , .A2( us22_n515 ) , .A1( us22_n541 ) , .A3( us22_n577 ) , .A4( us22_n613 ) );
  NOR3_X1 us22_U240 (.ZN( us22_n750 ) , .A2( us22_n851 ) , .A1( us22_n861 ) , .A3( us22_n863 ) );
  NOR2_X1 us22_U241 (.ZN( us22_n528 ) , .A2( us22_n742 ) , .A1( us22_n790 ) );
  NOR2_X1 us22_U242 (.A1( us22_n747 ) , .ZN( us22_n765 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U243 (.A2( us22_n742 ) , .ZN( us22_n753 ) , .A1( us22_n803 ) );
  NOR2_X1 us22_U244 (.ZN( us22_n542 ) , .A2( us22_n783 ) , .A1( us22_n790 ) );
  NOR2_X1 us22_U245 (.ZN( us22_n661 ) , .A1( us22_n727 ) , .A2( us22_n783 ) );
  NOR2_X1 us22_U246 (.ZN( us22_n629 ) , .A1( us22_n722 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U247 (.ZN( us22_n733 ) , .A2( us22_n801 ) , .A1( us22_n803 ) );
  NOR2_X1 us22_U248 (.ZN( us22_n612 ) , .A1( us22_n760 ) , .A2( us22_n810 ) );
  OAI22_X1 us22_U249 (.B1( us22_n438 ) , .ZN( us22_n442 ) , .A2( us22_n726 ) , .A1( us22_n742 ) , .B2( us22_n747 ) );
  NOR4_X1 us22_U25 (.A4( us22_n530 ) , .A3( us22_n531 ) , .A2( us22_n532 ) , .ZN( us22_n533 ) , .A1( us22_n818 ) );
  NOR3_X1 us22_U250 (.ZN( us22_n438 ) , .A2( us22_n834 ) , .A3( us22_n835 ) , .A1( us22_n844 ) );
  NOR2_X1 us22_U251 (.ZN( us22_n504 ) , .A2( us22_n726 ) , .A1( us22_n760 ) );
  NOR2_X1 us22_U252 (.ZN( us22_n514 ) , .A1( us22_n706 ) , .A2( us22_n742 ) );
  NOR2_X1 us22_U253 (.ZN( us22_n715 ) , .A2( us22_n742 ) , .A1( us22_n784 ) );
  NOR2_X1 us22_U254 (.ZN( us22_n552 ) , .A1( us22_n784 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U255 (.ZN( us22_n515 ) , .A1( us22_n706 ) , .A2( us22_n801 ) );
  NOR2_X1 us22_U256 (.ZN( us22_n556 ) , .A1( us22_n706 ) , .A2( us22_n814 ) );
  NOR2_X1 us22_U257 (.ZN( us22_n519 ) , .A1( us22_n788 ) , .A2( us22_n810 ) );
  NOR2_X1 us22_U258 (.ZN( us22_n628 ) , .A1( us22_n745 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U259 (.ZN( us22_n713 ) , .A1( us22_n803 ) , .A2( us22_n815 ) );
  NOR4_X1 us22_U26 (.A4( us22_n539 ) , .A3( us22_n540 ) , .A2( us22_n541 ) , .ZN( us22_n548 ) , .A1( us22_n686 ) );
  AOI21_X1 us22_U260 (.ZN( us22_n569 ) , .B2( us22_n695 ) , .B1( us22_n804 ) , .A( us22_n810 ) );
  INV_X1 us22_U261 (.A( us22_n761 ) , .ZN( us22_n864 ) );
  NOR2_X1 us22_U262 (.ZN( us22_n653 ) , .A1( us22_n788 ) , .A2( us22_n813 ) );
  NOR2_X1 us22_U263 (.ZN( us22_n666 ) , .A2( us22_n706 ) , .A1( us22_n788 ) );
  NOR2_X1 us22_U264 (.ZN( us22_n654 ) , .A1( us22_n745 ) , .A2( us22_n778 ) );
  NOR2_X1 us22_U265 (.ZN( us22_n554 ) , .A1( us22_n760 ) , .A2( us22_n803 ) );
  NOR2_X1 us22_U266 (.ZN( us22_n540 ) , .A1( us22_n760 ) , .A2( us22_n789 ) );
  NOR2_X1 us22_U267 (.ZN( us22_n699 ) , .A2( us22_n784 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U268 (.ZN( us22_n607 ) , .A2( us22_n722 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U269 (.A1( us22_n728 ) , .ZN( us22_n763 ) , .A2( us22_n784 ) );
  NOR2_X1 us22_U27 (.ZN( us22_n678 ) , .A2( us22_n832 ) , .A1( us22_n837 ) );
  AOI21_X1 us22_U270 (.A( us22_n813 ) , .B2( us22_n814 ) , .B1( us22_n815 ) , .ZN( us22_n816 ) );
  INV_X1 us22_U271 (.A( us22_n727 ) , .ZN( us22_n866 ) );
  NOR2_X1 us22_U272 (.ZN( us22_n577 ) , .A2( us22_n706 ) , .A1( us22_n728 ) );
  NOR2_X1 us22_U273 (.ZN( us22_n531 ) , .A2( us22_n722 ) , .A1( us22_n728 ) );
  AOI21_X1 us22_U274 (.B1( us22_n623 ) , .ZN( us22_n625 ) , .A( us22_n761 ) , .B2( us22_n812 ) );
  AOI21_X1 us22_U275 (.A( us22_n810 ) , .B2( us22_n811 ) , .B1( us22_n812 ) , .ZN( us22_n817 ) );
  AOI21_X1 us22_U276 (.ZN( us22_n513 ) , .A( us22_n727 ) , .B1( us22_n748 ) , .B2( us22_n801 ) );
  AOI21_X1 us22_U277 (.ZN( us22_n497 ) , .B1( us22_n678 ) , .A( us22_n810 ) , .B2( us22_n814 ) );
  AOI21_X1 us22_U278 (.ZN( us22_n476 ) , .B2( us22_n695 ) , .A( us22_n747 ) , .B1( us22_n777 ) );
  NOR2_X1 us22_U279 (.ZN( us22_n580 ) , .A1( us22_n742 ) , .A2( us22_n813 ) );
  NOR4_X1 us22_U28 (.A4( us22_n512 ) , .A3( us22_n513 ) , .A2( us22_n514 ) , .A1( us22_n515 ) , .ZN( us22_n522 ) );
  NOR2_X1 us22_U280 (.ZN( us22_n640 ) , .A2( us22_n786 ) , .A1( us22_n789 ) );
  AOI21_X1 us22_U281 (.ZN( us22_n591 ) , .B1( us22_n748 ) , .A( us22_n790 ) , .B2( us22_n811 ) );
  NOR2_X1 us22_U282 (.A2( us22_n706 ) , .A1( us22_n760 ) , .ZN( us22_n792 ) );
  AOI21_X1 us22_U283 (.ZN( us22_n624 ) , .B2( us22_n667 ) , .A( us22_n788 ) , .B1( us22_n789 ) );
  NOR2_X1 us22_U284 (.ZN( us22_n668 ) , .A1( us22_n788 ) , .A2( us22_n803 ) );
  NOR2_X1 us22_U285 (.ZN( us22_n518 ) , .A2( us22_n706 ) , .A1( us22_n812 ) );
  AOI21_X1 us22_U286 (.ZN( us22_n475 ) , .A( us22_n667 ) , .B1( us22_n748 ) , .B2( us22_n804 ) );
  NOR2_X1 us22_U287 (.ZN( us22_n557 ) , .A2( us22_n789 ) , .A1( us22_n801 ) );
  NOR2_X1 us22_U288 (.ZN( us22_n517 ) , .A2( us22_n697 ) , .A1( us22_n814 ) );
  NOR2_X1 us22_U289 (.ZN( us22_n681 ) , .A2( us22_n697 ) , .A1( us22_n801 ) );
  AOI222_X1 us22_U29 (.ZN( us22_n523 ) , .A1( us22_n832 ) , .B2( us22_n835 ) , .C1( us22_n842 ) , .C2( us22_n848 ) , .A2( us22_n850 ) , .B1( us22_n864 ) );
  NOR2_X1 us22_U290 (.ZN( us22_n651 ) , .A1( us22_n760 ) , .A2( us22_n784 ) );
  INV_X1 us22_U291 (.A( us22_n811 ) , .ZN( us22_n834 ) );
  AOI21_X1 us22_U292 (.ZN( us22_n508 ) , .B2( us22_n667 ) , .A( us22_n728 ) , .B1( us22_n813 ) );
  AOI21_X1 us22_U293 (.ZN( us22_n537 ) , .B2( us22_n810 ) , .A( us22_n812 ) , .B1( us22_n813 ) );
  AOI21_X1 us22_U294 (.ZN( us22_n538 ) , .A( us22_n761 ) , .B2( us22_n777 ) , .B1( us22_n815 ) );
  NOR2_X1 us22_U295 (.ZN( us22_n579 ) , .A1( us22_n667 ) , .A2( us22_n786 ) );
  AOI21_X1 us22_U296 (.ZN( us22_n587 ) , .B2( us22_n697 ) , .B1( us22_n813 ) , .A( us22_n815 ) );
  AOI21_X1 us22_U297 (.B1( us22_n697 ) , .ZN( us22_n698 ) , .A( us22_n730 ) , .B2( us22_n761 ) );
  AOI21_X1 us22_U298 (.ZN( us22_n589 ) , .B2( us22_n761 ) , .A( us22_n783 ) , .B1( us22_n810 ) );
  AOI21_X1 us22_U299 (.ZN( us22_n496 ) , .A( us22_n722 ) , .B2( us22_n760 ) , .B1( us22_n812 ) );
  NAND2_X2 us22_U3 (.A1( us22_n445 ) , .A2( us22_n446 ) , .ZN( us22_n784 ) );
  NOR4_X1 us22_U30 (.A3( us22_n519 ) , .A1( us22_n520 ) , .ZN( us22_n521 ) , .A2( us22_n671 ) , .A4( us22_n767 ) );
  AOI21_X1 us22_U300 (.ZN( us22_n550 ) , .B1( us22_n667 ) , .A( us22_n695 ) , .B2( us22_n803 ) );
  NOR2_X1 us22_U301 (.ZN( us22_n545 ) , .A1( us22_n697 ) , .A2( us22_n742 ) );
  INV_X1 us22_U302 (.A( us22_n789 ) , .ZN( us22_n871 ) );
  INV_X1 us22_U303 (.A( us22_n810 ) , .ZN( us22_n852 ) );
  AOI21_X1 us22_U304 (.ZN( us22_n638 ) , .B2( us22_n745 ) , .A( us22_n790 ) , .B1( us22_n801 ) );
  AOI21_X1 us22_U305 (.ZN( us22_n647 ) , .B1( us22_n727 ) , .B2( us22_n761 ) , .A( us22_n811 ) );
  NOR2_X1 us22_U306 (.ZN( us22_n683 ) , .A1( us22_n727 ) , .A2( us22_n814 ) );
  AOI21_X1 us22_U307 (.B1( us22_n684 ) , .ZN( us22_n685 ) , .A( us22_n726 ) , .B2( us22_n759 ) );
  AOI21_X1 us22_U308 (.ZN( us22_n567 ) , .B1( us22_n748 ) , .B2( us22_n760 ) , .A( us22_n778 ) );
  AOI21_X1 us22_U309 (.ZN( us22_n498 ) , .A( us22_n695 ) , .B1( us22_n706 ) , .B2( us22_n784 ) );
  AOI221_X1 us22_U31 (.A( us22_n779 ) , .ZN( us22_n796 ) , .C2( us22_n835 ) , .B2( us22_n836 ) , .B1( us22_n863 ) , .C1( us22_n864 ) );
  NOR2_X1 us22_U310 (.ZN( us22_n566 ) , .A1( us22_n727 ) , .A2( us22_n760 ) );
  AOI21_X1 us22_U311 (.ZN( us22_n637 ) , .B2( us22_n747 ) , .A( us22_n786 ) , .B1( us22_n810 ) );
  NOR2_X1 us22_U312 (.ZN( us22_n564 ) , .A2( us22_n695 ) , .A1( us22_n761 ) );
  NOR2_X1 us22_U313 (.ZN( us22_n578 ) , .A2( us22_n695 ) , .A1( us22_n789 ) );
  AOI21_X1 us22_U314 (.ZN( us22_n512 ) , .A( us22_n777 ) , .B2( us22_n790 ) , .B1( us22_n810 ) );
  INV_X1 us22_U315 (.A( us22_n697 ) , .ZN( us22_n851 ) );
  NOR2_X1 us22_U316 (.ZN( us22_n663 ) , .A1( us22_n778 ) , .A2( us22_n811 ) );
  AOI21_X1 us22_U317 (.ZN( us22_n448 ) , .B2( us22_n790 ) , .A( us22_n801 ) , .B1( us22_n813 ) );
  NOR2_X1 us22_U318 (.ZN( us22_n630 ) , .A2( us22_n695 ) , .A1( us22_n722 ) );
  AOI21_X1 us22_U319 (.ZN( us22_n562 ) , .B1( us22_n722 ) , .A( us22_n777 ) , .B2( us22_n789 ) );
  NOR4_X1 us22_U32 (.A4( us22_n791 ) , .A3( us22_n792 ) , .A2( us22_n793 ) , .A1( us22_n794 ) , .ZN( us22_n795 ) );
  AOI21_X1 us22_U320 (.ZN( us22_n495 ) , .A( us22_n777 ) , .B2( us22_n789 ) , .B1( us22_n802 ) );
  AOI21_X1 us22_U321 (.ZN( us22_n687 ) , .B2( us22_n747 ) , .B1( us22_n761 ) , .A( us22_n804 ) );
  NOR2_X1 us22_U322 (.ZN( us22_n527 ) , .A1( us22_n706 ) , .A2( us22_n777 ) );
  NOR2_X1 us22_U323 (.ZN( us22_n576 ) , .A1( us22_n706 ) , .A2( us22_n811 ) );
  AOI21_X1 us22_U324 (.ZN( us22_n648 ) , .A( us22_n777 ) , .B1( us22_n790 ) , .B2( us22_n803 ) );
  NOR2_X1 us22_U325 (.ZN( us22_n682 ) , .A1( us22_n789 ) , .A2( us22_n811 ) );
  NOR2_X1 us22_U326 (.A2( us22_n811 ) , .A1( us22_n813 ) , .ZN( us22_n819 ) );
  AOI21_X1 us22_U327 (.A( us22_n788 ) , .B2( us22_n789 ) , .B1( us22_n790 ) , .ZN( us22_n791 ) );
  AOI21_X1 us22_U328 (.A( us22_n731 ) , .ZN( us22_n732 ) , .B2( us22_n778 ) , .B1( us22_n790 ) );
  NOR2_X1 us22_U329 (.ZN( us22_n565 ) , .A1( us22_n745 ) , .A2( us22_n803 ) );
  NOR4_X1 us22_U33 (.A4( us22_n774 ) , .A3( us22_n775 ) , .A1( us22_n776 ) , .ZN( us22_n797 ) , .A2( us22_n799 ) );
  NOR2_X1 us22_U330 (.ZN( us22_n581 ) , .A1( us22_n790 ) , .A2( us22_n815 ) );
  NOR2_X1 us22_U331 (.ZN( us22_n532 ) , .A1( us22_n722 ) , .A2( us22_n786 ) );
  AOI21_X1 us22_U332 (.ZN( us22_n639 ) , .B1( us22_n678 ) , .A( us22_n789 ) , .B2( us22_n815 ) );
  NOR2_X1 us22_U333 (.ZN( us22_n709 ) , .A1( us22_n760 ) , .A2( us22_n761 ) );
  NOR2_X1 us22_U334 (.ZN( us22_n680 ) , .A2( us22_n706 ) , .A1( us22_n815 ) );
  INV_X1 us22_U335 (.A( us22_n695 ) , .ZN( us22_n836 ) );
  INV_X1 us22_U336 (.A( us22_n813 ) , .ZN( us22_n853 ) );
  AOI21_X1 us22_U337 (.ZN( us22_n440 ) , .A( us22_n697 ) , .B1( us22_n731 ) , .B2( us22_n748 ) );
  OAI21_X1 us22_U338 (.A( us22_n696 ) , .ZN( us22_n700 ) , .B2( us22_n748 ) , .B1( us22_n802 ) );
  OAI21_X1 us22_U339 (.ZN( us22_n696 ) , .B2( us22_n831 ) , .B1( us22_n836 ) , .A( us22_n858 ) );
  NOR4_X1 us22_U34 (.A3( us22_n753 ) , .A2( us22_n754 ) , .A1( us22_n755 ) , .ZN( us22_n756 ) , .A4( us22_n867 ) );
  NAND2_X1 us22_U340 (.ZN( us22_n751 ) , .A1( us22_n761 ) , .A2( us22_n803 ) );
  INV_X1 us22_U341 (.A( us22_n778 ) , .ZN( us22_n848 ) );
  INV_X1 us22_U342 (.A( us22_n783 ) , .ZN( us22_n844 ) );
  NAND2_X1 us22_U343 (.ZN( us22_n669 ) , .A1( us22_n804 ) , .A2( us22_n814 ) );
  NAND2_X1 us22_U344 (.ZN( us22_n712 ) , .A1( us22_n726 ) , .A2( us22_n778 ) );
  NAND2_X1 us22_U345 (.A2( us22_n760 ) , .A1( us22_n804 ) , .ZN( us22_n808 ) );
  NAND2_X2 us22_U346 (.A2( us22_n439 ) , .A1( us22_n445 ) , .ZN( us22_n782 ) );
  AOI21_X1 us22_U347 (.ZN( us22_n441 ) , .B1( us22_n787 ) , .B2( us22_n789 ) , .A( us22_n812 ) );
  NOR2_X1 us22_U348 (.ZN( us22_n468 ) , .A2( us22_n777 ) , .A1( us22_n813 ) );
  OAI21_X1 us22_U349 (.A( us22_n785 ) , .B2( us22_n786 ) , .B1( us22_n787 ) , .ZN( us22_n793 ) );
  AOI211_X1 us22_U35 (.B( us22_n743 ) , .A( us22_n744 ) , .ZN( us22_n757 ) , .C1( us22_n830 ) , .C2( us22_n851 ) );
  OAI21_X1 us22_U350 (.ZN( us22_n785 ) , .A( us22_n837 ) , .B1( us22_n861 ) , .B2( us22_n871 ) );
  NOR2_X1 us22_U351 (.ZN( us22_n524 ) , .A1( us22_n722 ) , .A2( us22_n748 ) );
  NOR2_X1 us22_U352 (.ZN( us22_n710 ) , .A2( us22_n722 ) , .A1( us22_n788 ) );
  NOR2_X1 us22_U353 (.ZN( us22_n482 ) , .A1( us22_n786 ) , .A2( us22_n803 ) );
  NAND2_X1 us22_U354 (.A1( us22_n697 ) , .A2( us22_n727 ) , .ZN( us22_n780 ) );
  NOR2_X1 us22_U355 (.ZN( us22_n516 ) , .A1( us22_n706 ) , .A2( us22_n786 ) );
  NAND2_X1 us22_U356 (.A2( us22_n747 ) , .A1( us22_n784 ) , .ZN( us22_n807 ) );
  OAI21_X1 us22_U357 (.A( us22_n729 ) , .B1( us22_n730 ) , .ZN( us22_n734 ) , .B2( us22_n803 ) );
  OAI21_X1 us22_U358 (.ZN( us22_n729 ) , .A( us22_n831 ) , .B2( us22_n850 ) , .B1( us22_n871 ) );
  INV_X1 us22_U359 (.A( us22_n815 ) , .ZN( us22_n842 ) );
  NOR3_X1 us22_U36 (.A3( us22_n739 ) , .A2( us22_n740 ) , .A1( us22_n741 ) , .ZN( us22_n758 ) );
  INV_X1 us22_U360 (.A( us22_n722 ) , .ZN( us22_n854 ) );
  AND2_X1 us22_U361 (.ZN( us22_n730 ) , .A1( us22_n777 ) , .A2( us22_n783 ) );
  AOI221_X1 us22_U362 (.A( us22_n762 ) , .ZN( us22_n772 ) , .C2( us22_n808 ) , .B2( us22_n833 ) , .C1( us22_n853 ) , .B1( us22_n864 ) );
  AOI21_X1 us22_U363 (.B2( us22_n761 ) , .ZN( us22_n762 ) , .A( us22_n786 ) , .B1( us22_n790 ) );
  INV_X1 us22_U364 (.A( us22_n759 ) , .ZN( us22_n833 ) );
  NAND2_X1 us22_U365 (.A1( us22_n453 ) , .A2( us22_n469 ) , .ZN( us22_n801 ) );
  NAND2_X1 us22_U366 (.A1( us22_n449 ) , .A2( us22_n452 ) , .ZN( us22_n812 ) );
  NAND2_X1 us22_U367 (.A1( us22_n449 ) , .A2( us22_n469 ) , .ZN( us22_n814 ) );
  NAND2_X1 us22_U368 (.A1( us22_n452 ) , .A2( us22_n459 ) , .ZN( us22_n811 ) );
  NAND2_X1 us22_U369 (.A1( us22_n451 ) , .A2( us22_n459 ) , .ZN( us22_n742 ) );
  NOR4_X1 us22_U37 (.A4( us22_n732 ) , .A3( us22_n733 ) , .A2( us22_n734 ) , .A1( us22_n735 ) , .ZN( us22_n736 ) );
  NAND2_X1 us22_U370 (.A1( us22_n450 ) , .A2( us22_n463 ) , .ZN( us22_n667 ) );
  NAND2_X1 us22_U371 (.A2( us22_n446 ) , .A1( us22_n458 ) , .ZN( us22_n726 ) );
  NAND2_X1 us22_U372 (.A1( us22_n453 ) , .A2( us22_n460 ) , .ZN( us22_n748 ) );
  NAND2_X1 us22_U373 (.A2( us22_n451 ) , .A1( us22_n453 ) , .ZN( us22_n804 ) );
  NAND2_X1 us22_U374 (.A2( us22_n452 ) , .A1( us22_n470 ) , .ZN( us22_n777 ) );
  NAND2_X1 us22_U375 (.A1( us22_n451 ) , .A2( us22_n470 ) , .ZN( us22_n783 ) );
  NAND2_X1 us22_U376 (.A2( us22_n462 ) , .A1( us22_n463 ) , .ZN( us22_n810 ) );
  NAND2_X1 us22_U377 (.A1( us22_n439 ) , .A2( us22_n458 ) , .ZN( us22_n697 ) );
  NAND2_X1 us22_U378 (.A2( us22_n447 ) , .A1( us22_n450 ) , .ZN( us22_n761 ) );
  NAND2_X1 us22_U379 (.A2( us22_n446 ) , .A1( us22_n450 ) , .ZN( us22_n727 ) );
  AOI211_X1 us22_U38 (.B( us22_n723 ) , .A( us22_n724 ) , .ZN( us22_n737 ) , .C1( us22_n841 ) , .C2( us22_n853 ) );
  NAND2_X2 us22_U380 (.A2( us22_n459 ) , .A1( us22_n469 ) , .ZN( us22_n695 ) );
  NOR2_X1 us22_U381 (.ZN( us22_n445 ) , .A2( us22_n847 ) , .A1( us22_n856 ) );
  NAND2_X1 us22_U382 (.A2( us22_n459 ) , .A1( us22_n460 ) , .ZN( us22_n745 ) );
  NAND2_X1 us22_U383 (.A1( us22_n460 ) , .A2( us22_n470 ) , .ZN( us22_n786 ) );
  NOR2_X1 us22_U384 (.ZN( us22_n463 ) , .A2( us22_n845 ) , .A1( us22_n846 ) );
  NOR2_X1 us22_U385 (.ZN( us22_n451 ) , .A1( us22_n824 ) , .A2( us22_n825 ) );
  NOR2_X1 us22_U386 (.ZN( us22_n449 ) , .A1( us22_n826 ) , .A2( us22_n827 ) );
  NAND2_X1 us22_U387 (.A2( us22_n452 ) , .A1( us22_n453 ) , .ZN( us22_n728 ) );
  NAND2_X1 us22_U388 (.A1( us22_n449 ) , .A2( us22_n460 ) , .ZN( us22_n788 ) );
  NAND2_X2 us22_U389 (.A2( us22_n446 ) , .A1( us22_n462 ) , .ZN( us22_n813 ) );
  NOR3_X1 us22_U39 (.A3( us22_n720 ) , .A1( us22_n721 ) , .ZN( us22_n738 ) , .A2( us22_n739 ) );
  NAND2_X2 us22_U390 (.A2( us22_n439 ) , .A1( us22_n450 ) , .ZN( us22_n789 ) );
  NAND2_X2 us22_U391 (.A1( us22_n447 ) , .A2( us22_n462 ) , .ZN( us22_n722 ) );
  NAND2_X2 us22_U392 (.A1( us22_n447 ) , .A2( us22_n458 ) , .ZN( us22_n790 ) );
  NAND2_X2 us22_U393 (.A1( us22_n439 ) , .A2( us22_n462 ) , .ZN( us22_n706 ) );
  NAND2_X2 us22_U394 (.A2( us22_n469 ) , .A1( us22_n470 ) , .ZN( us22_n815 ) );
  NAND2_X2 us22_U395 (.A2( us22_n458 ) , .A1( us22_n463 ) , .ZN( us22_n778 ) );
  NAND2_X1 us22_U396 (.A1( us22_n445 ) , .A2( us22_n447 ) , .ZN( us22_n803 ) );
  NOR2_X1 us22_U397 (.A2( sa22_6 ) , .A1( sa22_7 ) , .ZN( us22_n462 ) );
  NOR2_X1 us22_U398 (.A2( sa22_4 ) , .ZN( us22_n447 ) , .A1( us22_n846 ) );
  NOR2_X1 us22_U399 (.A2( sa22_5 ) , .ZN( us22_n446 ) , .A1( us22_n845 ) );
  INV_X1 us22_U4 (.A( us22_n784 ) , .ZN( us22_n860 ) );
  NAND4_X1 us22_U40 (.ZN( sa20_sr_3 ) , .A4( us22_n702 ) , .A3( us22_n703 ) , .A2( us22_n704 ) , .A1( us22_n705 ) );
  NOR2_X1 us22_U400 (.A2( sa22_7 ) , .ZN( us22_n458 ) , .A1( us22_n847 ) );
  NOR2_X1 us22_U401 (.A2( sa22_4 ) , .A1( sa22_5 ) , .ZN( us22_n439 ) );
  NOR2_X1 us22_U402 (.A2( sa22_1 ) , .ZN( us22_n469 ) , .A1( us22_n824 ) );
  NOR2_X1 us22_U403 (.A2( sa22_2 ) , .A1( sa22_3 ) , .ZN( us22_n470 ) );
  NOR2_X1 us22_U404 (.A2( sa22_6 ) , .ZN( us22_n450 ) , .A1( us22_n856 ) );
  NOR2_X1 us22_U405 (.A2( sa22_2 ) , .ZN( us22_n459 ) , .A1( us22_n827 ) );
  NOR2_X1 us22_U406 (.A2( sa22_0 ) , .ZN( us22_n452 ) , .A1( us22_n825 ) );
  NOR2_X1 us22_U407 (.A2( sa22_0 ) , .A1( sa22_1 ) , .ZN( us22_n460 ) );
  NOR2_X1 us22_U408 (.A2( sa22_3 ) , .ZN( us22_n453 ) , .A1( us22_n826 ) );
  INV_X1 us22_U409 (.A( sa22_6 ) , .ZN( us22_n847 ) );
  NOR4_X1 us22_U41 (.A4( us22_n698 ) , .A3( us22_n699 ) , .A2( us22_n700 ) , .A1( us22_n701 ) , .ZN( us22_n702 ) );
  INV_X1 us22_U410 (.A( sa22_3 ) , .ZN( us22_n827 ) );
  INV_X1 us22_U411 (.A( sa22_1 ) , .ZN( us22_n825 ) );
  INV_X1 us22_U412 (.A( sa22_2 ) , .ZN( us22_n826 ) );
  INV_X1 us22_U413 (.A( sa22_0 ) , .ZN( us22_n824 ) );
  INV_X1 us22_U414 (.A( sa22_7 ) , .ZN( us22_n856 ) );
  INV_X1 us22_U415 (.A( sa22_5 ) , .ZN( us22_n846 ) );
  OAI221_X1 us22_U416 (.A( us22_n781 ) , .C2( us22_n782 ) , .B2( us22_n783 ) , .B1( us22_n784 ) , .ZN( us22_n794 ) , .C1( us22_n811 ) );
  NAND2_X1 us22_U417 (.A1( us22_n727 ) , .A2( us22_n782 ) , .ZN( us22_n809 ) );
  OAI22_X1 us22_U418 (.ZN( us22_n586 ) , .A2( us22_n745 ) , .B2( us22_n760 ) , .A1( us22_n761 ) , .B1( us22_n782 ) );
  OAI221_X1 us22_U419 (.A( us22_n694 ) , .ZN( us22_n701 ) , .C2( us22_n782 ) , .C1( us22_n783 ) , .B1( us22_n784 ) , .B2( us22_n804 ) );
  AOI211_X1 us22_U42 (.B( us22_n692 ) , .A( us22_n693 ) , .ZN( us22_n703 ) , .C2( us22_n829 ) , .C1( us22_n849 ) );
  AOI21_X1 us22_U420 (.ZN( us22_n590 ) , .B1( us22_n726 ) , .B2( us22_n782 ) , .A( us22_n788 ) );
  AOI21_X1 us22_U421 (.ZN( us22_n621 ) , .B1( us22_n697 ) , .A( us22_n777 ) , .B2( us22_n782 ) );
  AOI21_X1 us22_U422 (.ZN( us22_n646 ) , .A( us22_n760 ) , .B2( us22_n782 ) , .B1( us22_n790 ) );
  OAI22_X1 us22_U423 (.ZN( us22_n679 ) , .A1( us22_n697 ) , .A2( us22_n728 ) , .B2( us22_n782 ) , .B1( us22_n815 ) );
  OAI21_X1 us22_U424 (.A( us22_n611 ) , .ZN( us22_n614 ) , .B1( us22_n623 ) , .B2( us22_n782 ) );
  NOR2_X1 us22_U425 (.ZN( us22_n608 ) , .A1( us22_n782 ) , .A2( us22_n814 ) );
  OAI222_X1 us22_U426 (.A2( us22_n667 ) , .ZN( us22_n672 ) , .B1( us22_n745 ) , .B2( us22_n782 ) , .C2( us22_n786 ) , .C1( us22_n813 ) , .A1( us22_n815 ) );
  NOR2_X1 us22_U427 (.ZN( us22_n649 ) , .A1( us22_n782 ) , .A2( us22_n786 ) );
  NOR2_X1 us22_U428 (.ZN( us22_n598 ) , .A2( us22_n695 ) , .A1( us22_n782 ) );
  NOR2_X1 us22_U429 (.ZN( us22_n551 ) , .A2( us22_n742 ) , .A1( us22_n782 ) );
  NOR2_X1 us22_U43 (.ZN( us22_n705 ) , .A2( us22_n774 ) , .A1( us22_n798 ) );
  INV_X1 us22_U430 (.A( us22_n782 ) , .ZN( us22_n859 ) );
  NAND4_X1 us22_U431 (.ZN( sa20_sr_2 ) , .A4( us22_n641 ) , .A3( us22_n642 ) , .A1( us22_n643 ) , .A2( us22_n644 ) );
  AOI221_X1 us22_U432 (.A( us22_n574 ) , .ZN( us22_n585 ) , .B2( us22_n829 ) , .C2( us22_n841 ) , .B1( us22_n852 ) , .C1( us22_n859 ) );
  AOI21_X1 us22_U433 (.ZN( us22_n574 ) , .B2( us22_n722 ) , .B1( us22_n746 ) , .A( us22_n783 ) );
  AOI211_X1 us22_U434 (.A( us22_n635 ) , .ZN( us22_n643 ) , .B( us22_n741 ) , .C2( us22_n837 ) , .C1( us22_n852 ) );
  NAND4_X1 us22_U435 (.A4( us22_n631 ) , .A3( us22_n632 ) , .A2( us22_n633 ) , .A1( us22_n634 ) , .ZN( us22_n741 ) );
  INV_X1 us22_U436 (.A( sa22_4 ) , .ZN( us22_n845 ) );
  NAND3_X1 us22_U437 (.ZN( sa20_sr_6 ) , .A3( us22_n795 ) , .A2( us22_n796 ) , .A1( us22_n797 ) );
  NAND3_X1 us22_U438 (.ZN( sa20_sr_5 ) , .A3( us22_n756 ) , .A2( us22_n757 ) , .A1( us22_n758 ) );
  NAND3_X1 us22_U439 (.ZN( sa20_sr_4 ) , .A3( us22_n736 ) , .A2( us22_n737 ) , .A1( us22_n738 ) );
  AOI222_X1 us22_U44 (.B2( us22_n636 ) , .ZN( us22_n642 ) , .B1( us22_n839 ) , .A1( us22_n840 ) , .C2( us22_n844 ) , .C1( us22_n861 ) , .A2( us22_n863 ) );
  NAND3_X1 us22_U440 (.A3( us22_n673 ) , .A2( us22_n674 ) , .A1( us22_n675 ) , .ZN( us22_n805 ) );
  NAND3_X1 us22_U441 (.ZN( us22_n636 ) , .A3( us22_n706 ) , .A2( us22_n722 ) , .A1( us22_n790 ) );
  NAND3_X1 us22_U442 (.A3( us22_n616 ) , .A2( us22_n617 ) , .A1( us22_n618 ) , .ZN( us22_n723 ) );
  NAND3_X1 us22_U443 (.A3( us22_n583 ) , .A2( us22_n584 ) , .A1( us22_n585 ) , .ZN( us22_n619 ) );
  NAND3_X1 us22_U444 (.ZN( us22_n563 ) , .A3( us22_n678 ) , .A2( us22_n748 ) , .A1( us22_n783 ) );
  NAND3_X1 us22_U445 (.A3( us22_n521 ) , .A2( us22_n522 ) , .A1( us22_n523 ) , .ZN( us22_n740 ) );
  NAND3_X1 us22_U446 (.A3( us22_n510 ) , .A1( us22_n511 ) , .ZN( us22_n606 ) , .A2( us22_n869 ) );
  NAND3_X1 us22_U447 (.A3( us22_n465 ) , .A2( us22_n466 ) , .A1( us22_n467 ) , .ZN( us22_n775 ) );
  NOR4_X1 us22_U45 (.A4( us22_n637 ) , .A3( us22_n638 ) , .A2( us22_n639 ) , .A1( us22_n640 ) , .ZN( us22_n641 ) );
  NOR3_X1 us22_U46 (.A2( us22_n605 ) , .A1( us22_n606 ) , .ZN( us22_n644 ) , .A3( us22_n720 ) );
  NOR2_X1 us22_U47 (.ZN( us22_n802 ) , .A1( us22_n852 ) , .A2( us22_n859 ) );
  NAND4_X1 us22_U48 (.ZN( sa20_sr_7 ) , .A4( us22_n820 ) , .A3( us22_n821 ) , .A2( us22_n822 ) , .A1( us22_n823 ) );
  NOR4_X1 us22_U49 (.A4( us22_n816 ) , .A3( us22_n817 ) , .A2( us22_n818 ) , .A1( us22_n819 ) , .ZN( us22_n820 ) );
  NOR3_X1 us22_U5 (.ZN( us22_n596 ) , .A1( us22_n606 ) , .A3( us22_n721 ) , .A2( us22_n740 ) );
  AOI222_X1 us22_U50 (.C2( us22_n807 ) , .B2( us22_n808 ) , .A2( us22_n809 ) , .ZN( us22_n821 ) , .C1( us22_n830 ) , .A1( us22_n837 ) , .B1( us22_n851 ) );
  AOI211_X1 us22_U51 (.B( us22_n805 ) , .A( us22_n806 ) , .ZN( us22_n822 ) , .C1( us22_n840 ) , .C2( us22_n848 ) );
  NAND4_X1 us22_U52 (.ZN( sa20_sr_0 ) , .A4( us22_n499 ) , .A3( us22_n500 ) , .A2( us22_n501 ) , .A1( us22_n502 ) );
  AOI221_X1 us22_U53 (.A( us22_n495 ) , .ZN( us22_n500 ) , .B2( us22_n841 ) , .C1( us22_n844 ) , .C2( us22_n858 ) , .B1( us22_n860 ) );
  NOR4_X1 us22_U54 (.A4( us22_n496 ) , .A3( us22_n497 ) , .A2( us22_n498 ) , .ZN( us22_n499 ) , .A1( us22_n525 ) );
  AOI211_X1 us22_U55 (.A( us22_n494 ) , .ZN( us22_n501 ) , .B( us22_n800 ) , .C2( us22_n837 ) , .C1( us22_n849 ) );
  NOR2_X1 us22_U56 (.ZN( us22_n746 ) , .A1( us22_n859 ) , .A2( us22_n860 ) );
  NAND4_X1 us22_U57 (.ZN( sa20_sr_1 ) , .A4( us22_n593 ) , .A3( us22_n594 ) , .A2( us22_n595 ) , .A1( us22_n596 ) );
  NOR4_X1 us22_U58 (.A4( us22_n589 ) , .A3( us22_n590 ) , .A2( us22_n591 ) , .A1( us22_n592 ) , .ZN( us22_n593 ) );
  AOI211_X1 us22_U59 (.B( us22_n587 ) , .A( us22_n588 ) , .ZN( us22_n594 ) , .C2( us22_n809 ) , .C1( us22_n831 ) );
  NOR3_X1 us22_U6 (.A3( us22_n798 ) , .A2( us22_n799 ) , .A1( us22_n800 ) , .ZN( us22_n823 ) );
  AOI211_X1 us22_U60 (.A( us22_n586 ) , .ZN( us22_n595 ) , .B( us22_n619 ) , .C1( us22_n843 ) , .C2( us22_n853 ) );
  NOR2_X1 us22_U61 (.ZN( us22_n623 ) , .A2( us22_n834 ) , .A1( us22_n837 ) );
  AOI222_X1 us22_U62 (.ZN( us22_n467 ) , .B1( us22_n830 ) , .A1( us22_n837 ) , .C1( us22_n840 ) , .C2( us22_n849 ) , .A2( us22_n853 ) , .B2( us22_n863 ) );
  NOR4_X1 us22_U63 (.A1( us22_n464 ) , .ZN( us22_n465 ) , .A4( us22_n540 ) , .A2( us22_n552 ) , .A3( us22_n612 ) );
  AOI221_X1 us22_U64 (.ZN( us22_n466 ) , .C2( us22_n712 ) , .B2( us22_n829 ) , .C1( us22_n843 ) , .B1( us22_n858 ) , .A( us22_n862 ) );
  NAND4_X1 us22_U65 (.A4( us22_n601 ) , .A3( us22_n602 ) , .A2( us22_n603 ) , .A1( us22_n604 ) , .ZN( us22_n720 ) );
  NOR3_X1 us22_U66 (.A1( us22_n597 ) , .ZN( us22_n602 ) , .A3( us22_n661 ) , .A2( us22_n768 ) );
  NOR4_X1 us22_U67 (.A3( us22_n598 ) , .A2( us22_n599 ) , .A1( us22_n600 ) , .ZN( us22_n601 ) , .A4( us22_n653 ) );
  AOI222_X1 us22_U68 (.ZN( us22_n604 ) , .A1( us22_n828 ) , .C2( us22_n835 ) , .B1( us22_n840 ) , .A2( us22_n854 ) , .B2( us22_n859 ) , .C1( us22_n866 ) );
  NOR4_X1 us22_U69 (.A4( us22_n575 ) , .A3( us22_n576 ) , .A2( us22_n577 ) , .ZN( us22_n584 ) , .A1( us22_n681 ) );
  NOR3_X1 us22_U7 (.ZN( us22_n502 ) , .A2( us22_n677 ) , .A3( us22_n775 ) , .A1( us22_n874 ) );
  NOR4_X1 us22_U70 (.A1( us22_n582 ) , .ZN( us22_n583 ) , .A3( us22_n650 ) , .A2( us22_n660 ) , .A4( us22_n765 ) );
  AOI211_X1 us22_U71 (.B( us22_n621 ) , .A( us22_n622 ) , .ZN( us22_n633 ) , .C2( us22_n834 ) , .C1( us22_n861 ) );
  NOR4_X1 us22_U72 (.A4( us22_n627 ) , .A3( us22_n628 ) , .A2( us22_n629 ) , .A1( us22_n630 ) , .ZN( us22_n631 ) );
  NOR4_X1 us22_U73 (.A4( us22_n624 ) , .A3( us22_n625 ) , .A2( us22_n626 ) , .ZN( us22_n632 ) , .A1( us22_n662 ) );
  NAND4_X1 us22_U74 (.A4( us22_n655 ) , .A3( us22_n656 ) , .A2( us22_n657 ) , .A1( us22_n658 ) , .ZN( us22_n798 ) );
  NOR3_X1 us22_U75 (.A3( us22_n646 ) , .A2( us22_n647 ) , .A1( us22_n648 ) , .ZN( us22_n657 ) );
  NOR3_X1 us22_U76 (.A3( us22_n649 ) , .A2( us22_n650 ) , .A1( us22_n651 ) , .ZN( us22_n656 ) );
  NOR3_X1 us22_U77 (.A3( us22_n652 ) , .A2( us22_n653 ) , .A1( us22_n654 ) , .ZN( us22_n655 ) );
  NAND4_X1 us22_U78 (.A4( us22_n558 ) , .A3( us22_n559 ) , .A2( us22_n560 ) , .A1( us22_n561 ) , .ZN( us22_n605 ) );
  NOR4_X1 us22_U79 (.A4( us22_n554 ) , .A3( us22_n555 ) , .A2( us22_n556 ) , .A1( us22_n557 ) , .ZN( us22_n558 ) );
  INV_X1 us22_U8 (.A( us22_n704 ) , .ZN( us22_n874 ) );
  NOR4_X1 us22_U80 (.ZN( us22_n559 ) , .A1( us22_n651 ) , .A3( us22_n659 ) , .A4( us22_n683 ) , .A2( us22_n766 ) );
  NOR4_X1 us22_U81 (.A4( us22_n550 ) , .A3( us22_n551 ) , .A2( us22_n552 ) , .A1( us22_n553 ) , .ZN( us22_n560 ) );
  NAND4_X1 us22_U82 (.A4( us22_n770 ) , .A3( us22_n771 ) , .A2( us22_n772 ) , .A1( us22_n773 ) , .ZN( us22_n799 ) );
  NOR3_X1 us22_U83 (.A3( us22_n763 ) , .A2( us22_n764 ) , .A1( us22_n765 ) , .ZN( us22_n771 ) );
  NOR4_X1 us22_U84 (.A4( us22_n766 ) , .A3( us22_n767 ) , .A2( us22_n768 ) , .A1( us22_n769 ) , .ZN( us22_n770 ) );
  AOI222_X1 us22_U85 (.ZN( us22_n773 ) , .A1( us22_n828 ) , .C1( us22_n832 ) , .B2( us22_n839 ) , .A2( us22_n848 ) , .B1( us22_n859 ) , .C2( us22_n871 ) );
  NOR4_X1 us22_U86 (.A4( us22_n663 ) , .A3( us22_n664 ) , .A2( us22_n665 ) , .A1( us22_n666 ) , .ZN( us22_n674 ) );
  NOR4_X1 us22_U87 (.A4( us22_n659 ) , .A3( us22_n660 ) , .A2( us22_n661 ) , .A1( us22_n662 ) , .ZN( us22_n675 ) );
  NOR4_X1 us22_U88 (.A3( us22_n671 ) , .A1( us22_n672 ) , .ZN( us22_n673 ) , .A4( us22_n713 ) , .A2( us22_n857 ) );
  NOR2_X1 us22_U89 (.ZN( us22_n759 ) , .A1( us22_n831 ) , .A2( us22_n832 ) );
  NOR3_X1 us22_U9 (.A3( us22_n619 ) , .A2( us22_n620 ) , .ZN( us22_n634 ) , .A1( us22_n723 ) );
  AOI222_X1 us22_U90 (.ZN( us22_n511 ) , .C1( us22_n830 ) , .B2( us22_n835 ) , .A2( us22_n841 ) , .C2( us22_n860 ) , .B1( us22_n861 ) , .A1( us22_n864 ) );
  NOR4_X1 us22_U91 (.A4( us22_n507 ) , .A2( us22_n508 ) , .A1( us22_n509 ) , .ZN( us22_n510 ) , .A3( us22_n668 ) );
  INV_X1 us22_U92 (.A( us22_n503 ) , .ZN( us22_n869 ) );
  NAND4_X1 us22_U93 (.A4( us22_n454 ) , .A3( us22_n455 ) , .A2( us22_n456 ) , .A1( us22_n457 ) , .ZN( us22_n677 ) );
  NOR3_X1 us22_U94 (.ZN( us22_n455 ) , .A3( us22_n528 ) , .A1( us22_n553 ) , .A2( us22_n568 ) );
  AOI221_X1 us22_U95 (.A( us22_n448 ) , .ZN( us22_n457 ) , .C2( us22_n751 ) , .B1( us22_n830 ) , .C1( us22_n840 ) , .B2( us22_n859 ) );
  NOR4_X1 us22_U96 (.ZN( us22_n456 ) , .A2( us22_n507 ) , .A1( us22_n597 ) , .A4( us22_n626 ) , .A3( us22_n709 ) );
  NAND4_X1 us22_U97 (.A4( us22_n533 ) , .A3( us22_n534 ) , .A2( us22_n535 ) , .A1( us22_n536 ) , .ZN( us22_n620 ) );
  NOR4_X1 us22_U98 (.A4( us22_n524 ) , .A2( us22_n525 ) , .A1( us22_n526 ) , .ZN( us22_n536 ) , .A3( us22_n699 ) );
  NOR4_X1 us22_U99 (.A1( us22_n529 ) , .ZN( us22_n534 ) , .A2( us22_n652 ) , .A4( us22_n666 ) , .A3( us22_n763 ) );
  NOR2_X1 us32_U10 (.A1( us32_n678 ) , .ZN( us32_n693 ) , .A2( us32_n807 ) );
  AOI211_X1 us32_U100 (.B( us32_n477 ) , .A( us32_n478 ) , .ZN( us32_n482 ) , .C2( us32_n833 ) , .C1( us32_n861 ) );
  NOR4_X1 us32_U101 (.ZN( us32_n481 ) , .A3( us32_n532 ) , .A4( us32_n545 ) , .A2( us32_n567 ) , .A1( us32_n717 ) );
  NAND4_X1 us32_U102 (.A4( us32_n548 ) , .A3( us32_n549 ) , .A2( us32_n550 ) , .A1( us32_n551 ) , .ZN( us32_n745 ) );
  NOR3_X1 us32_U103 (.ZN( us32_n549 ) , .A2( us32_n651 ) , .A1( us32_n667 ) , .A3( us32_n771 ) );
  AOI211_X1 us32_U104 (.B( us32_n539 ) , .A( us32_n540 ) , .ZN( us32_n551 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NOR4_X1 us32_U105 (.A4( us32_n541 ) , .A3( us32_n542 ) , .A2( us32_n543 ) , .ZN( us32_n550 ) , .A1( us32_n688 ) );
  NOR4_X1 us32_U106 (.ZN( us32_n620 ) , .A1( us32_n656 ) , .A3( us32_n666 ) , .A4( us32_n682 ) , .A2( us32_n766 ) );
  NOR4_X1 us32_U107 (.A4( us32_n609 ) , .A3( us32_n610 ) , .A2( us32_n611 ) , .A1( us32_n612 ) , .ZN( us32_n619 ) );
  NOR4_X1 us32_U108 (.A4( us32_n614 ) , .A3( us32_n615 ) , .A2( us32_n616 ) , .A1( us32_n617 ) , .ZN( us32_n618 ) );
  NOR2_X1 us32_U109 (.ZN( us32_n686 ) , .A1( us32_n831 ) , .A2( us32_n832 ) );
  NOR3_X1 us32_U11 (.ZN( us32_n504 ) , .A2( us32_n679 ) , .A3( us32_n777 ) , .A1( us32_n876 ) );
  NAND4_X1 us32_U110 (.A4( us32_n485 ) , .A3( us32_n486 ) , .A2( us32_n487 ) , .A1( us32_n488 ) , .ZN( us32_n778 ) );
  NOR4_X1 us32_U111 (.A4( us32_n484 ) , .ZN( us32_n487 ) , .A1( us32_n566 ) , .A2( us32_n581 ) , .A3( us32_n602 ) );
  NOR4_X1 us32_U112 (.ZN( us32_n486 ) , .A1( us32_n507 ) , .A2( us32_n519 ) , .A4( us32_n546 ) , .A3( us32_n611 ) );
  NOR4_X1 us32_U113 (.ZN( us32_n485 ) , .A2( us32_n533 ) , .A1( us32_n558 ) , .A3( us32_n631 ) , .A4( us32_n718 ) );
  NAND4_X1 us32_U114 (.A4( us32_n691 ) , .A3( us32_n692 ) , .A1( us32_n693 ) , .ZN( us32_n776 ) , .A2( us32_n872 ) );
  AOI221_X1 us32_U115 (.A( us32_n681 ) , .ZN( us32_n692 ) , .B2( us32_n840 ) , .C1( us32_n842 ) , .C2( us32_n862 ) , .B1( us32_n865 ) );
  INV_X1 us32_U116 (.A( us32_n679 ) , .ZN( us32_n872 ) );
  NOR4_X1 us32_U117 (.A4( us32_n687 ) , .A3( us32_n688 ) , .A2( us32_n689 ) , .A1( us32_n690 ) , .ZN( us32_n691 ) );
  NAND4_X1 us32_U118 (.A4( us32_n473 ) , .A3( us32_n474 ) , .A2( us32_n475 ) , .A1( us32_n476 ) , .ZN( us32_n678 ) );
  NOR4_X1 us32_U119 (.ZN( us32_n475 ) , .A1( us32_n531 ) , .A3( us32_n568 ) , .A4( us32_n600 ) , .A2( us32_n642 ) );
  INV_X1 us32_U12 (.A( us32_n706 ) , .ZN( us32_n876 ) );
  NOR4_X1 us32_U120 (.A4( us32_n470 ) , .ZN( us32_n476 ) , .A3( us32_n556 ) , .A1( us32_n735 ) , .A2( us32_n755 ) );
  NOR4_X1 us32_U121 (.ZN( us32_n473 ) , .A2( us32_n521 ) , .A4( us32_n594 ) , .A1( us32_n609 ) , .A3( us32_n629 ) );
  NAND4_X1 us32_U122 (.A4( us32_n719 ) , .A3( us32_n720 ) , .A2( us32_n721 ) , .ZN( us32_n741 ) , .A1( us32_n857 ) );
  INV_X1 us32_U123 (.A( us32_n709 ) , .ZN( us32_n857 ) );
  AOI221_X1 us32_U124 (.A( us32_n710 ) , .ZN( us32_n721 ) , .C2( us32_n844 ) , .B2( us32_n845 ) , .C1( us32_n861 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U125 (.A4( us32_n715 ) , .A3( us32_n716 ) , .A2( us32_n717 ) , .A1( us32_n718 ) , .ZN( us32_n719 ) );
  NOR2_X1 us32_U126 (.ZN( us32_n733 ) , .A2( us32_n832 ) , .A1( us32_n845 ) );
  NOR2_X1 us32_U127 (.ZN( us32_n789 ) , .A2( us32_n862 ) , .A1( us32_n868 ) );
  NAND4_X1 us32_U128 (.A4( us32_n573 ) , .A3( us32_n574 ) , .A1( us32_n575 ) , .ZN( us32_n723 ) , .A2( us32_n874 ) );
  AOI221_X1 us32_U129 (.A( us32_n564 ) , .C2( us32_n565 ) , .ZN( us32_n574 ) , .B2( us32_n845 ) , .B1( us32_n852 ) , .C1( us32_n853 ) );
  INV_X1 us32_U13 (.A( us32_n607 ) , .ZN( us32_n874 ) );
  NOR4_X1 us32_U130 (.A4( us32_n569 ) , .A3( us32_n570 ) , .A2( us32_n571 ) , .A1( us32_n572 ) , .ZN( us32_n573 ) );
  NOR2_X1 us32_U131 (.ZN( us32_n575 ) , .A1( us32_n622 ) , .A2( us32_n745 ) );
  NOR2_X1 us32_U132 (.ZN( us32_n748 ) , .A1( us32_n861 ) , .A2( us32_n862 ) );
  NAND4_X1 us32_U133 (.A4( us32_n633 ) , .A3( us32_n634 ) , .A2( us32_n635 ) , .A1( us32_n636 ) , .ZN( us32_n743 ) );
  AOI211_X1 us32_U134 (.B( us32_n623 ) , .A( us32_n624 ) , .ZN( us32_n635 ) , .C2( us32_n836 ) , .C1( us32_n863 ) );
  NOR4_X1 us32_U135 (.A4( us32_n629 ) , .A3( us32_n630 ) , .A2( us32_n631 ) , .A1( us32_n632 ) , .ZN( us32_n633 ) );
  NOR4_X1 us32_U136 (.A4( us32_n626 ) , .A3( us32_n627 ) , .A2( us32_n628 ) , .ZN( us32_n634 ) , .A1( us32_n664 ) );
  NAND4_X1 us32_U137 (.A4( us32_n493 ) , .A3( us32_n494 ) , .A1( us32_n495 ) , .ZN( us32_n802 ) , .A2( us32_n867 ) );
  AOI221_X1 us32_U138 (.A( us32_n489 ) , .ZN( us32_n494 ) , .B2( us32_n836 ) , .C2( us32_n841 ) , .C1( us32_n851 ) , .B1( us32_n860 ) );
  INV_X1 us32_U139 (.A( us32_n778 ) , .ZN( us32_n867 ) );
  INV_X1 us32_U14 (.A( us32_n680 ) , .ZN( us32_n840 ) );
  NOR4_X1 us32_U140 (.A2( us32_n491 ) , .A1( us32_n492 ) , .ZN( us32_n493 ) , .A3( us32_n580 ) , .A4( us32_n612 ) );
  NOR4_X1 us32_U141 (.A4( us32_n734 ) , .A3( us32_n735 ) , .A2( us32_n736 ) , .A1( us32_n737 ) , .ZN( us32_n738 ) );
  AOI211_X1 us32_U142 (.B( us32_n725 ) , .A( us32_n726 ) , .ZN( us32_n739 ) , .C1( us32_n843 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U143 (.A3( us32_n722 ) , .A1( us32_n723 ) , .ZN( us32_n740 ) , .A2( us32_n741 ) );
  NOR2_X1 us32_U144 (.ZN( us32_n647 ) , .A1( us32_n854 ) , .A2( us32_n868 ) );
  INV_X1 us32_U145 (.A( us32_n762 ) , .ZN( us32_n830 ) );
  INV_X1 us32_U146 (.A( us32_n754 ) , .ZN( us32_n869 ) );
  OAI21_X1 us32_U147 (.B1( us32_n753 ) , .ZN( us32_n754 ) , .A( us32_n845 ) , .B2( us32_n868 ) );
  INV_X1 us32_U148 (.A( us32_n697 ) , .ZN( us32_n838 ) );
  OR4_X1 us32_U149 (.ZN( us32_n492 ) , .A4( us32_n534 ) , .A2( us32_n547 ) , .A1( us32_n559 ) , .A3( us32_n632 ) );
  NOR4_X1 us32_U15 (.A4( us32_n445 ) , .A3( us32_n446 ) , .A2( us32_n516 ) , .A1( us32_n541 ) , .ZN( us32_n706 ) );
  OR4_X1 us32_U150 (.A4( us32_n566 ) , .A3( us32_n567 ) , .A2( us32_n568 ) , .ZN( us32_n572 ) , .A1( us32_n665 ) );
  OR4_X1 us32_U151 (.A4( us32_n682 ) , .A3( us32_n683 ) , .A2( us32_n684 ) , .A1( us32_n685 ) , .ZN( us32_n690 ) );
  OR4_X1 us32_U152 (.ZN( us32_n466 ) , .A4( us32_n518 ) , .A3( us32_n529 ) , .A2( us32_n578 ) , .A1( us32_n712 ) );
  OR4_X1 us32_U153 (.A4( us32_n518 ) , .A2( us32_n519 ) , .A1( us32_n520 ) , .ZN( us32_n522 ) , .A3( us32_n821 ) );
  OR4_X1 us32_U154 (.A4( us32_n580 ) , .A3( us32_n581 ) , .A2( us32_n582 ) , .A1( us32_n583 ) , .ZN( us32_n584 ) );
  NAND2_X1 us32_U155 (.ZN( us32_n613 ) , .A2( us32_n837 ) , .A1( us32_n873 ) );
  OR3_X1 us32_U156 (.A3( us32_n506 ) , .A2( us32_n507 ) , .A1( us32_n508 ) , .ZN( us32_n511 ) );
  INV_X1 us32_U157 (.A( us32_n672 ) , .ZN( us32_n859 ) );
  AOI21_X1 us32_U158 (.A( us32_n670 ) , .B1( us32_n671 ) , .ZN( us32_n672 ) , .B2( us32_n856 ) );
  INV_X1 us32_U159 (.A( us32_n463 ) , .ZN( us32_n864 ) );
  OR3_X1 us32_U16 (.ZN( us32_n446 ) , .A1( us32_n528 ) , .A3( us32_n577 ) , .A2( us32_n875 ) );
  OAI21_X1 us32_U160 (.ZN( us32_n463 ) , .B1( us32_n809 ) , .A( us32_n834 ) , .B2( us32_n851 ) );
  OAI222_X1 us32_U161 (.B2( us32_n708 ) , .ZN( us32_n709 ) , .C2( us32_n724 ) , .B1( us32_n747 ) , .A1( us32_n806 ) , .C1( us32_n814 ) , .A2( us32_n815 ) );
  NAND2_X1 us32_U162 (.A1( us32_n447 ) , .A2( us32_n465 ) , .ZN( us32_n749 ) );
  AOI22_X1 us32_U163 (.A2( us32_n782 ) , .ZN( us32_n783 ) , .B2( us32_n831 ) , .A1( us32_n834 ) , .B1( us32_n863 ) );
  AOI22_X1 us32_U164 (.ZN( us32_n696 ) , .A1( us32_n830 ) , .B2( us32_n843 ) , .A2( us32_n865 ) , .B1( us32_n868 ) );
  INV_X1 us32_U165 (.A( us32_n730 ) , .ZN( us32_n839 ) );
  AOI221_X1 us32_U166 (.A( us32_n483 ) , .ZN( us32_n488 ) , .B1( us32_n831 ) , .C2( us32_n844 ) , .C1( us32_n852 ) , .B2( us32_n862 ) );
  OAI22_X1 us32_U167 (.ZN( us32_n483 ) , .A1( us32_n708 ) , .B2( us32_n785 ) , .A2( us32_n806 ) , .B1( us32_n812 ) );
  INV_X1 us32_U168 (.A( us32_n790 ) , .ZN( us32_n832 ) );
  OAI221_X1 us32_U169 (.A( us32_n727 ) , .C2( us32_n728 ) , .B2( us32_n729 ) , .B1( us32_n730 ) , .ZN( us32_n737 ) , .C1( us32_n817 ) );
  OR4_X1 us32_U17 (.A4( us32_n442 ) , .A2( us32_n443 ) , .A1( us32_n444 ) , .ZN( us32_n445 ) , .A3( us32_n553 ) );
  AOI22_X1 us32_U170 (.ZN( us32_n727 ) , .B1( us32_n832 ) , .A2( us32_n838 ) , .A1( us32_n863 ) , .B2( us32_n866 ) );
  NAND2_X1 us32_U171 (.A1( us32_n451 ) , .A2( us32_n453 ) , .ZN( us32_n762 ) );
  INV_X1 us32_U172 (.A( us32_n786 ) , .ZN( us32_n862 ) );
  OAI22_X1 us32_U173 (.ZN( us32_n710 ) , .A2( us32_n728 ) , .B2( us32_n729 ) , .A1( us32_n744 ) , .B1( us32_n813 ) );
  INV_X1 us32_U174 (.A( us32_n816 ) , .ZN( us32_n831 ) );
  OAI22_X1 us32_U175 (.ZN( us32_n489 ) , .A1( us32_n724 ) , .B2( us32_n728 ) , .B1( us32_n730 ) , .A2( us32_n779 ) );
  OAI22_X1 us32_U176 (.ZN( us32_n624 ) , .B1( us32_n669 ) , .B2( us32_n747 ) , .A1( us32_n815 ) , .A2( us32_n816 ) );
  INV_X1 us32_U177 (.A( us32_n788 ) , .ZN( us32_n845 ) );
  OAI22_X1 us32_U178 (.A1( us32_n724 ) , .ZN( us32_n726 ) , .B2( us32_n750 ) , .B1( us32_n812 ) , .A2( us32_n816 ) );
  INV_X1 us32_U179 (.A( us32_n744 ) , .ZN( us32_n837 ) );
  INV_X1 us32_U18 (.A( us32_n613 ) , .ZN( us32_n875 ) );
  OAI22_X1 us32_U180 (.B2( us32_n779 ) , .B1( us32_n780 ) , .ZN( us32_n781 ) , .A2( us32_n814 ) , .A1( us32_n815 ) );
  INV_X1 us32_U181 (.A( us32_n814 ) , .ZN( us32_n833 ) );
  INV_X1 us32_U182 (.A( us32_n669 ) , .ZN( us32_n865 ) );
  OAI22_X1 us32_U183 (.B2( us32_n744 ) , .ZN( us32_n746 ) , .A2( us32_n762 ) , .B1( us32_n780 ) , .A1( us32_n792 ) );
  OAI22_X1 us32_U184 (.ZN( us32_n496 ) , .A2( us32_n744 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n806 ) );
  AOI211_X1 us32_U185 (.A( us32_n637 ) , .ZN( us32_n645 ) , .B( us32_n743 ) , .C2( us32_n839 ) , .C1( us32_n854 ) );
  OAI22_X1 us32_U186 (.ZN( us32_n637 ) , .A1( us32_n699 ) , .B2( us32_n728 ) , .A2( us32_n762 ) , .B1( us32_n816 ) );
  INV_X1 us32_U187 (.A( us32_n750 ) , .ZN( us32_n842 ) );
  OAI22_X1 us32_U188 (.B1( us32_n490 ) , .ZN( us32_n491 ) , .A1( us32_n686 ) , .A2( us32_n763 ) , .B2( us32_n817 ) );
  NOR3_X1 us32_U189 (.ZN( us32_n490 ) , .A1( us32_n782 ) , .A2( us32_n850 ) , .A3( us32_n863 ) );
  INV_X1 us32_U19 (.A( us32_n749 ) , .ZN( us32_n863 ) );
  OAI22_X1 us32_U190 (.ZN( us32_n695 ) , .A2( us32_n730 ) , .A1( us32_n780 ) , .B1( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U191 (.ZN( us32_n666 ) , .A1( us32_n728 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U192 (.ZN( us32_n594 ) , .A2( us32_n697 ) , .A1( us32_n728 ) );
  NOR2_X1 us32_U193 (.ZN( us32_n570 ) , .A1( us32_n728 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U194 (.ZN( us32_n654 ) , .A1( us32_n728 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U195 (.ZN( us32_n546 ) , .A2( us32_n780 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U196 (.ZN( us32_n532 ) , .A2( us32_n749 ) , .A1( us32_n750 ) );
  NOR2_X1 us32_U197 (.ZN( us32_n577 ) , .A2( us32_n699 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U198 (.ZN( us32_n615 ) , .A1( us32_n785 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U199 (.ZN( us32_n629 ) , .A2( us32_n728 ) , .A1( us32_n785 ) );
  AOI222_X1 us32_U20 (.ZN( us32_n605 ) , .B2( us32_n671 ) , .B1( us32_n753 ) , .C2( us32_n831 ) , .A1( us32_n833 ) , .A2( us32_n862 ) , .C1( us32_n863 ) );
  NOR2_X1 us32_U200 (.ZN( us32_n718 ) , .A2( us32_n724 ) , .A1( us32_n744 ) );
  NOR2_X1 us32_U201 (.ZN( us32_n628 ) , .A2( us32_n669 ) , .A1( us32_n785 ) );
  INV_X1 us32_U202 (.A( us32_n728 ) , .ZN( us32_n852 ) );
  NOR2_X1 us32_U203 (.A2( us32_n744 ) , .ZN( us32_n769 ) , .A1( us32_n812 ) );
  NOR2_X1 us32_U204 (.ZN( us32_n531 ) , .A2( us32_n780 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U205 (.A2( us32_n708 ) , .A1( us32_n750 ) , .ZN( us32_n771 ) );
  NOR2_X1 us32_U206 (.ZN( us32_n599 ) , .A2( us32_n791 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U207 (.ZN( us32_n611 ) , .A2( us32_n780 ) , .A1( us32_n806 ) );
  NOR2_X1 us32_U208 (.ZN( us32_n652 ) , .A1( us32_n669 ) , .A2( us32_n814 ) );
  INV_X1 us32_U209 (.A( us32_n792 ) , .ZN( us32_n851 ) );
  AOI222_X1 us32_U21 (.ZN( us32_n563 ) , .B1( us32_n830 ) , .C1( us32_n841 ) , .A2( us32_n843 ) , .A1( us32_n854 ) , .B2( us32_n863 ) , .C2( us32_n873 ) );
  NOR2_X1 us32_U210 (.A1( us32_n699 ) , .ZN( us32_n768 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U211 (.A1( us32_n669 ) , .ZN( us32_n673 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U212 (.ZN( us32_n541 ) , .A2( us32_n697 ) , .A1( us32_n699 ) );
  NOR2_X1 us32_U213 (.ZN( us32_n602 ) , .A1( us32_n669 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U214 (.A1( us32_n669 ) , .ZN( us32_n688 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U215 (.ZN( us32_n667 ) , .A1( us32_n750 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U216 (.ZN( us32_n555 ) , .A1( us32_n750 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U217 (.ZN( us32_n508 ) , .A2( us32_n780 ) , .A1( us32_n785 ) );
  NOR2_X1 us32_U218 (.ZN( us32_n543 ) , .A2( us32_n708 ) , .A1( us32_n785 ) );
  INV_X1 us32_U219 (.A( us32_n747 ) , .ZN( us32_n834 ) );
  AOI222_X1 us32_U22 (.ZN( us32_n660 ) , .A2( us32_n839 ) , .B1( us32_n841 ) , .C2( us32_n845 ) , .A1( us32_n860 ) , .C1( us32_n863 ) , .B2( us32_n870 ) );
  NOR2_X1 us32_U220 (.ZN( us32_n664 ) , .A1( us32_n785 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U221 (.A1( us32_n669 ) , .ZN( us32_n766 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U222 (.ZN( us32_n527 ) , .A1( us32_n669 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U223 (.ZN( us32_n661 ) , .A1( us32_n729 ) , .A2( us32_n790 ) );
  NOR2_X1 us32_U224 (.ZN( us32_n601 ) , .A2( us32_n780 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U225 (.ZN( us32_n507 ) , .A1( us32_n812 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U226 (.ZN( us32_n528 ) , .A2( us32_n724 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U227 (.ZN( us32_n509 ) , .A1( us32_n729 ) , .A2( us32_n779 ) );
  NOR2_X1 us32_U228 (.ZN( us32_n557 ) , .A1( us32_n792 ) , .A2( us32_n814 ) );
  NOR2_X1 us32_U229 (.ZN( us32_n545 ) , .A1( us32_n749 ) , .A2( us32_n814 ) );
  INV_X1 us32_U23 (.A( us32_n647 ) , .ZN( us32_n870 ) );
  OAI22_X1 us32_U230 (.B1( us32_n440 ) , .ZN( us32_n444 ) , .A2( us32_n728 ) , .A1( us32_n744 ) , .B2( us32_n749 ) );
  NOR3_X1 us32_U231 (.ZN( us32_n440 ) , .A2( us32_n836 ) , .A3( us32_n837 ) , .A1( us32_n846 ) );
  NOR2_X1 us32_U232 (.ZN( us32_n662 ) , .A2( us32_n697 ) , .A1( us32_n729 ) );
  OAI22_X1 us32_U233 (.B2( us32_n750 ) , .B1( us32_n751 ) , .A1( us32_n752 ) , .ZN( us32_n756 ) , .A2( us32_n806 ) );
  NOR2_X1 us32_U234 (.ZN( us32_n751 ) , .A2( us32_n852 ) , .A1( us32_n860 ) );
  NOR3_X1 us32_U235 (.ZN( us32_n752 ) , .A2( us32_n853 ) , .A1( us32_n863 ) , .A3( us32_n865 ) );
  NOR2_X1 us32_U236 (.ZN( us32_n544 ) , .A2( us32_n785 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U237 (.ZN( us32_n663 ) , .A1( us32_n729 ) , .A2( us32_n785 ) );
  INV_X1 us32_U238 (.A( us32_n806 ) , .ZN( us32_n841 ) );
  NOR2_X1 us32_U239 (.ZN( us32_n506 ) , .A2( us32_n728 ) , .A1( us32_n762 ) );
  NOR4_X1 us32_U24 (.A4( us32_n544 ) , .A3( us32_n545 ) , .A2( us32_n546 ) , .A1( us32_n547 ) , .ZN( us32_n548 ) );
  NOR2_X1 us32_U240 (.ZN( us32_n631 ) , .A1( us32_n724 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U241 (.ZN( us32_n614 ) , .A1( us32_n762 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U242 (.ZN( us32_n530 ) , .A2( us32_n744 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U243 (.ZN( us32_n558 ) , .A1( us32_n708 ) , .A2( us32_n816 ) );
  NOR2_X1 us32_U244 (.ZN( us32_n516 ) , .A1( us32_n708 ) , .A2( us32_n744 ) );
  NOR2_X1 us32_U245 (.A2( us32_n697 ) , .ZN( us32_n716 ) , .A1( us32_n792 ) );
  NOR2_X1 us32_U246 (.A1( us32_n749 ) , .ZN( us32_n767 ) , .A2( us32_n803 ) );
  NOR2_X1 us32_U247 (.ZN( us32_n521 ) , .A1( us32_n790 ) , .A2( us32_n812 ) );
  NOR2_X1 us32_U248 (.ZN( us32_n655 ) , .A1( us32_n790 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U249 (.ZN( us32_n668 ) , .A2( us32_n708 ) , .A1( us32_n790 ) );
  NOR4_X1 us32_U25 (.ZN( us32_n479 ) , .A1( us32_n520 ) , .A4( us32_n557 ) , .A3( us32_n582 ) , .A2( us32_n630 ) );
  NOR2_X1 us32_U250 (.ZN( us32_n517 ) , .A1( us32_n708 ) , .A2( us32_n803 ) );
  INV_X1 us32_U251 (.A( us32_n763 ) , .ZN( us32_n866 ) );
  NOR2_X1 us32_U252 (.ZN( us32_n542 ) , .A1( us32_n762 ) , .A2( us32_n791 ) );
  NOR2_X1 us32_U253 (.ZN( us32_n630 ) , .A1( us32_n747 ) , .A2( us32_n815 ) );
  INV_X1 us32_U254 (.A( us32_n729 ) , .ZN( us32_n868 ) );
  NOR2_X1 us32_U255 (.ZN( us32_n609 ) , .A2( us32_n724 ) , .A1( us32_n817 ) );
  AOI21_X1 us32_U256 (.A( us32_n815 ) , .B2( us32_n816 ) , .B1( us32_n817 ) , .ZN( us32_n818 ) );
  NOR2_X1 us32_U257 (.ZN( us32_n579 ) , .A2( us32_n708 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U258 (.ZN( us32_n533 ) , .A2( us32_n724 ) , .A1( us32_n730 ) );
  NOR2_X1 us32_U259 (.ZN( us32_n642 ) , .A2( us32_n788 ) , .A1( us32_n791 ) );
  NOR4_X1 us32_U26 (.ZN( us32_n456 ) , .A2( us32_n517 ) , .A1( us32_n543 ) , .A3( us32_n579 ) , .A4( us32_n615 ) );
  AOI21_X1 us32_U260 (.B1( us32_n625 ) , .ZN( us32_n627 ) , .A( us32_n763 ) , .B2( us32_n814 ) );
  NOR2_X1 us32_U261 (.ZN( us32_n656 ) , .A1( us32_n747 ) , .A2( us32_n780 ) );
  AOI21_X1 us32_U262 (.A( us32_n812 ) , .B2( us32_n813 ) , .B1( us32_n814 ) , .ZN( us32_n819 ) );
  NOR2_X1 us32_U263 (.A2( us32_n697 ) , .A1( us32_n780 ) , .ZN( us32_n820 ) );
  AOI21_X1 us32_U264 (.ZN( us32_n499 ) , .B1( us32_n680 ) , .A( us32_n812 ) , .B2( us32_n816 ) );
  NOR2_X1 us32_U265 (.A2( us32_n708 ) , .A1( us32_n762 ) , .ZN( us32_n794 ) );
  AOI21_X1 us32_U266 (.ZN( us32_n593 ) , .B1( us32_n750 ) , .A( us32_n792 ) , .B2( us32_n813 ) );
  AOI21_X1 us32_U267 (.ZN( us32_n626 ) , .B2( us32_n669 ) , .A( us32_n790 ) , .B1( us32_n791 ) );
  NOR2_X1 us32_U268 (.ZN( us32_n520 ) , .A2( us32_n708 ) , .A1( us32_n814 ) );
  NOR2_X1 us32_U269 (.A1( us32_n697 ) , .ZN( us32_n770 ) , .A2( us32_n815 ) );
  NOR4_X1 us32_U27 (.A4( us32_n532 ) , .A3( us32_n533 ) , .A2( us32_n534 ) , .ZN( us32_n535 ) , .A1( us32_n820 ) );
  NOR2_X1 us32_U270 (.ZN( us32_n582 ) , .A1( us32_n744 ) , .A2( us32_n815 ) );
  NOR2_X1 us32_U271 (.ZN( us32_n519 ) , .A2( us32_n699 ) , .A1( us32_n816 ) );
  AOI21_X1 us32_U272 (.ZN( us32_n477 ) , .A( us32_n669 ) , .B1( us32_n750 ) , .B2( us32_n806 ) );
  AOI21_X1 us32_U273 (.ZN( us32_n510 ) , .B2( us32_n669 ) , .A( us32_n730 ) , .B1( us32_n815 ) );
  INV_X1 us32_U274 (.A( us32_n813 ) , .ZN( us32_n836 ) );
  AOI21_X1 us32_U275 (.ZN( us32_n589 ) , .B2( us32_n699 ) , .B1( us32_n815 ) , .A( us32_n817 ) );
  AOI21_X1 us32_U276 (.ZN( us32_n515 ) , .A( us32_n729 ) , .B1( us32_n750 ) , .B2( us32_n803 ) );
  AOI21_X1 us32_U277 (.ZN( us32_n539 ) , .B2( us32_n812 ) , .A( us32_n814 ) , .B1( us32_n815 ) );
  NOR2_X1 us32_U278 (.ZN( us32_n581 ) , .A1( us32_n669 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U279 (.ZN( us32_n547 ) , .A1( us32_n699 ) , .A2( us32_n744 ) );
  NOR4_X1 us32_U28 (.ZN( us32_n474 ) , .A1( us32_n506 ) , .A3( us32_n544 ) , .A2( us32_n583 ) , .A4( us32_n716 ) );
  AOI21_X1 us32_U280 (.ZN( us32_n540 ) , .A( us32_n763 ) , .B2( us32_n779 ) , .B1( us32_n817 ) );
  AOI21_X1 us32_U281 (.B1( us32_n699 ) , .ZN( us32_n700 ) , .A( us32_n732 ) , .B2( us32_n763 ) );
  AOI21_X1 us32_U282 (.ZN( us32_n591 ) , .B2( us32_n763 ) , .A( us32_n785 ) , .B1( us32_n812 ) );
  INV_X1 us32_U283 (.A( us32_n791 ) , .ZN( us32_n873 ) );
  NOR2_X1 us32_U284 (.ZN( us32_n559 ) , .A2( us32_n791 ) , .A1( us32_n803 ) );
  AOI21_X1 us32_U285 (.ZN( us32_n498 ) , .A( us32_n724 ) , .B2( us32_n762 ) , .B1( us32_n814 ) );
  NOR2_X1 us32_U286 (.ZN( us32_n683 ) , .A2( us32_n699 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U287 (.ZN( us32_n685 ) , .A1( us32_n729 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U288 (.B1( us32_n686 ) , .ZN( us32_n687 ) , .A( us32_n728 ) , .B2( us32_n761 ) );
  AOI21_X1 us32_U289 (.ZN( us32_n569 ) , .B1( us32_n750 ) , .B2( us32_n762 ) , .A( us32_n780 ) );
  AOI221_X1 us32_U29 (.A( us32_n713 ) , .B2( us32_n714 ) , .ZN( us32_n720 ) , .C1( us32_n832 ) , .B1( us32_n839 ) , .C2( us32_n863 ) );
  AOI21_X1 us32_U290 (.ZN( us32_n649 ) , .B1( us32_n729 ) , .B2( us32_n763 ) , .A( us32_n813 ) );
  NOR2_X1 us32_U291 (.ZN( us32_n568 ) , .A1( us32_n729 ) , .A2( us32_n762 ) );
  INV_X1 us32_U292 (.A( us32_n699 ) , .ZN( us32_n853 ) );
  NOR2_X1 us32_U293 (.ZN( us32_n566 ) , .A2( us32_n697 ) , .A1( us32_n763 ) );
  AOI21_X1 us32_U294 (.ZN( us32_n514 ) , .A( us32_n779 ) , .B2( us32_n792 ) , .B1( us32_n812 ) );
  AOI21_X1 us32_U295 (.ZN( us32_n639 ) , .B2( us32_n749 ) , .A( us32_n788 ) , .B1( us32_n812 ) );
  NOR2_X1 us32_U296 (.ZN( us32_n665 ) , .A1( us32_n780 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U297 (.ZN( us32_n571 ) , .B2( us32_n697 ) , .B1( us32_n806 ) , .A( us32_n812 ) );
  AOI21_X1 us32_U298 (.ZN( us32_n564 ) , .B1( us32_n724 ) , .A( us32_n779 ) , .B2( us32_n791 ) );
  AOI21_X1 us32_U299 (.ZN( us32_n497 ) , .A( us32_n779 ) , .B2( us32_n791 ) , .B1( us32_n804 ) );
  NAND2_X1 us32_U3 (.A1( us32_n449 ) , .A2( us32_n464 ) , .ZN( us32_n724 ) );
  OR2_X1 us32_U30 (.A2( us32_n711 ) , .A1( us32_n712 ) , .ZN( us32_n713 ) );
  AOI21_X1 us32_U300 (.ZN( us32_n640 ) , .B2( us32_n747 ) , .A( us32_n792 ) , .B1( us32_n803 ) );
  NOR2_X1 us32_U301 (.ZN( us32_n578 ) , .A1( us32_n708 ) , .A2( us32_n813 ) );
  NOR2_X1 us32_U302 (.ZN( us32_n529 ) , .A1( us32_n708 ) , .A2( us32_n779 ) );
  AOI21_X1 us32_U303 (.ZN( us32_n689 ) , .B2( us32_n749 ) , .B1( us32_n763 ) , .A( us32_n806 ) );
  AOI21_X1 us32_U304 (.A( us32_n790 ) , .B2( us32_n791 ) , .B1( us32_n792 ) , .ZN( us32_n793 ) );
  AOI21_X1 us32_U305 (.ZN( us32_n478 ) , .B2( us32_n697 ) , .A( us32_n749 ) , .B1( us32_n779 ) );
  NOR2_X1 us32_U306 (.ZN( us32_n684 ) , .A1( us32_n791 ) , .A2( us32_n813 ) );
  AOI21_X1 us32_U307 (.ZN( us32_n450 ) , .B2( us32_n792 ) , .A( us32_n803 ) , .B1( us32_n815 ) );
  AOI21_X1 us32_U308 (.A( us32_n733 ) , .ZN( us32_n734 ) , .B2( us32_n780 ) , .B1( us32_n792 ) );
  NOR2_X1 us32_U309 (.A2( us32_n813 ) , .A1( us32_n815 ) , .ZN( us32_n821 ) );
  NOR2_X1 us32_U31 (.ZN( us32_n680 ) , .A2( us32_n834 ) , .A1( us32_n839 ) );
  AOI21_X1 us32_U310 (.ZN( us32_n641 ) , .B1( us32_n680 ) , .A( us32_n791 ) , .B2( us32_n817 ) );
  NOR2_X1 us32_U311 (.ZN( us32_n583 ) , .A1( us32_n792 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U312 (.ZN( us32_n711 ) , .A1( us32_n762 ) , .A2( us32_n763 ) );
  NOR2_X1 us32_U313 (.ZN( us32_n534 ) , .A1( us32_n724 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U314 (.ZN( us32_n632 ) , .A2( us32_n697 ) , .A1( us32_n724 ) );
  NOR2_X1 us32_U315 (.ZN( us32_n580 ) , .A2( us32_n697 ) , .A1( us32_n791 ) );
  NOR2_X1 us32_U316 (.ZN( us32_n682 ) , .A2( us32_n708 ) , .A1( us32_n817 ) );
  INV_X1 us32_U317 (.A( us32_n815 ) , .ZN( us32_n855 ) );
  AOI21_X1 us32_U318 (.ZN( us32_n442 ) , .A( us32_n699 ) , .B1( us32_n733 ) , .B2( us32_n750 ) );
  INV_X1 us32_U319 (.A( us32_n780 ) , .ZN( us32_n850 ) );
  NOR4_X1 us32_U32 (.A4( us32_n514 ) , .A3( us32_n515 ) , .A2( us32_n516 ) , .A1( us32_n517 ) , .ZN( us32_n524 ) );
  INV_X1 us32_U320 (.A( us32_n785 ) , .ZN( us32_n846 ) );
  NAND2_X1 us32_U321 (.ZN( us32_n714 ) , .A1( us32_n728 ) , .A2( us32_n780 ) );
  NAND2_X1 us32_U322 (.ZN( us32_n671 ) , .A1( us32_n806 ) , .A2( us32_n816 ) );
  AOI21_X1 us32_U323 (.ZN( us32_n443 ) , .B1( us32_n789 ) , .B2( us32_n791 ) , .A( us32_n814 ) );
  NOR2_X1 us32_U324 (.ZN( us32_n470 ) , .A2( us32_n779 ) , .A1( us32_n815 ) );
  NAND2_X1 us32_U325 (.A2( us32_n762 ) , .A1( us32_n806 ) , .ZN( us32_n810 ) );
  NOR2_X1 us32_U326 (.ZN( us32_n526 ) , .A1( us32_n724 ) , .A2( us32_n750 ) );
  OAI21_X1 us32_U327 (.A( us32_n787 ) , .B2( us32_n788 ) , .B1( us32_n789 ) , .ZN( us32_n795 ) );
  OAI21_X1 us32_U328 (.ZN( us32_n787 ) , .A( us32_n839 ) , .B1( us32_n863 ) , .B2( us32_n873 ) );
  NAND2_X1 us32_U329 (.A1( us32_n699 ) , .A2( us32_n729 ) , .ZN( us32_n782 ) );
  AOI222_X1 us32_U33 (.ZN( us32_n525 ) , .A1( us32_n834 ) , .B2( us32_n837 ) , .C1( us32_n844 ) , .C2( us32_n850 ) , .A2( us32_n852 ) , .B1( us32_n866 ) );
  NOR2_X1 us32_U330 (.ZN( us32_n712 ) , .A2( us32_n724 ) , .A1( us32_n790 ) );
  NOR2_X1 us32_U331 (.ZN( us32_n518 ) , .A1( us32_n708 ) , .A2( us32_n788 ) );
  OAI21_X1 us32_U332 (.A( us32_n698 ) , .ZN( us32_n702 ) , .B2( us32_n750 ) , .B1( us32_n804 ) );
  OAI21_X1 us32_U333 (.ZN( us32_n698 ) , .B2( us32_n833 ) , .B1( us32_n838 ) , .A( us32_n860 ) );
  INV_X1 us32_U334 (.A( us32_n817 ) , .ZN( us32_n844 ) );
  INV_X1 us32_U335 (.A( us32_n724 ) , .ZN( us32_n856 ) );
  OAI21_X1 us32_U336 (.ZN( us32_n731 ) , .A( us32_n833 ) , .B2( us32_n852 ) , .B1( us32_n873 ) );
  AND2_X1 us32_U337 (.ZN( us32_n732 ) , .A1( us32_n779 ) , .A2( us32_n785 ) );
  AOI221_X1 us32_U338 (.A( us32_n764 ) , .ZN( us32_n774 ) , .C2( us32_n810 ) , .B2( us32_n835 ) , .C1( us32_n855 ) , .B1( us32_n866 ) );
  AOI21_X1 us32_U339 (.B2( us32_n763 ) , .ZN( us32_n764 ) , .A( us32_n788 ) , .B1( us32_n792 ) );
  NOR4_X1 us32_U34 (.A3( us32_n521 ) , .A1( us32_n522 ) , .ZN( us32_n523 ) , .A2( us32_n673 ) , .A4( us32_n769 ) );
  INV_X1 us32_U340 (.A( us32_n761 ) , .ZN( us32_n835 ) );
  NAND2_X1 us32_U341 (.A2( us32_n448 ) , .A1( us32_n460 ) , .ZN( us32_n728 ) );
  NAND2_X1 us32_U342 (.A1( us32_n451 ) , .A2( us32_n454 ) , .ZN( us32_n814 ) );
  NAND2_X1 us32_U343 (.A1( us32_n455 ) , .A2( us32_n462 ) , .ZN( us32_n750 ) );
  NAND2_X1 us32_U344 (.A1( us32_n451 ) , .A2( us32_n471 ) , .ZN( us32_n816 ) );
  NAND2_X1 us32_U345 (.A1( us32_n454 ) , .A2( us32_n461 ) , .ZN( us32_n813 ) );
  NAND2_X1 us32_U346 (.A1( us32_n452 ) , .A2( us32_n465 ) , .ZN( us32_n669 ) );
  NAND2_X1 us32_U347 (.A1( us32_n453 ) , .A2( us32_n472 ) , .ZN( us32_n785 ) );
  NAND2_X1 us32_U348 (.A1( us32_n453 ) , .A2( us32_n461 ) , .ZN( us32_n744 ) );
  NAND2_X1 us32_U349 (.A2( us32_n453 ) , .A1( us32_n455 ) , .ZN( us32_n806 ) );
  AOI221_X1 us32_U35 (.A( us32_n781 ) , .ZN( us32_n798 ) , .C2( us32_n837 ) , .B2( us32_n838 ) , .B1( us32_n865 ) , .C1( us32_n866 ) );
  NAND2_X1 us32_U350 (.A1( us32_n455 ) , .A2( us32_n471 ) , .ZN( us32_n803 ) );
  NAND2_X1 us32_U351 (.A2( us32_n454 ) , .A1( us32_n472 ) , .ZN( us32_n779 ) );
  NAND2_X1 us32_U352 (.A2( us32_n464 ) , .A1( us32_n465 ) , .ZN( us32_n812 ) );
  NAND2_X1 us32_U353 (.A1( us32_n441 ) , .A2( us32_n460 ) , .ZN( us32_n699 ) );
  NAND2_X1 us32_U354 (.A2( us32_n448 ) , .A1( us32_n452 ) , .ZN( us32_n729 ) );
  NAND2_X1 us32_U355 (.A2( us32_n449 ) , .A1( us32_n452 ) , .ZN( us32_n763 ) );
  NOR2_X1 us32_U356 (.ZN( us32_n465 ) , .A2( us32_n847 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U357 (.ZN( us32_n453 ) , .A1( us32_n826 ) , .A2( us32_n827 ) );
  NAND2_X1 us32_U358 (.A1( us32_n462 ) , .A2( us32_n472 ) , .ZN( us32_n788 ) );
  NOR2_X1 us32_U359 (.ZN( us32_n451 ) , .A1( us32_n828 ) , .A2( us32_n829 ) );
  NOR4_X1 us32_U36 (.A4( us32_n793 ) , .A3( us32_n794 ) , .A2( us32_n795 ) , .A1( us32_n796 ) , .ZN( us32_n797 ) );
  NAND2_X1 us32_U360 (.A2( us32_n461 ) , .A1( us32_n462 ) , .ZN( us32_n747 ) );
  NAND2_X1 us32_U361 (.A1( us32_n451 ) , .A2( us32_n462 ) , .ZN( us32_n790 ) );
  NAND2_X2 us32_U362 (.A2( us32_n448 ) , .A1( us32_n464 ) , .ZN( us32_n815 ) );
  NAND2_X1 us32_U363 (.A2( us32_n441 ) , .A1( us32_n447 ) , .ZN( us32_n784 ) );
  NAND2_X1 us32_U364 (.A1( us32_n447 ) , .A2( us32_n449 ) , .ZN( us32_n805 ) );
  NAND2_X1 us32_U365 (.A2( us32_n454 ) , .A1( us32_n455 ) , .ZN( us32_n730 ) );
  NAND2_X2 us32_U366 (.A1( us32_n449 ) , .A2( us32_n460 ) , .ZN( us32_n792 ) );
  NAND2_X2 us32_U367 (.A2( us32_n460 ) , .A1( us32_n465 ) , .ZN( us32_n780 ) );
  NOR2_X1 us32_U368 (.ZN( us32_n447 ) , .A2( us32_n849 ) , .A1( us32_n858 ) );
  NAND2_X1 us32_U369 (.A1( us32_n447 ) , .A2( us32_n448 ) , .ZN( us32_n786 ) );
  NOR4_X1 us32_U37 (.A4( us32_n776 ) , .A3( us32_n777 ) , .A1( us32_n778 ) , .ZN( us32_n799 ) , .A2( us32_n801 ) );
  NAND2_X1 us32_U370 (.A2( us32_n471 ) , .A1( us32_n472 ) , .ZN( us32_n817 ) );
  NOR2_X1 us32_U371 (.A2( sa32_6 ) , .A1( sa32_7 ) , .ZN( us32_n464 ) );
  NOR2_X1 us32_U372 (.A2( sa32_7 ) , .ZN( us32_n460 ) , .A1( us32_n849 ) );
  NOR2_X1 us32_U373 (.A2( sa32_4 ) , .ZN( us32_n449 ) , .A1( us32_n848 ) );
  NOR2_X1 us32_U374 (.A2( sa32_4 ) , .A1( sa32_5 ) , .ZN( us32_n441 ) );
  NOR2_X1 us32_U375 (.A2( sa32_5 ) , .ZN( us32_n448 ) , .A1( us32_n847 ) );
  NOR2_X1 us32_U376 (.A2( sa32_2 ) , .A1( sa32_3 ) , .ZN( us32_n472 ) );
  NOR2_X1 us32_U377 (.A2( sa32_6 ) , .ZN( us32_n452 ) , .A1( us32_n858 ) );
  NOR2_X1 us32_U378 (.A2( sa32_1 ) , .ZN( us32_n471 ) , .A1( us32_n826 ) );
  NOR2_X1 us32_U379 (.A2( sa32_0 ) , .ZN( us32_n454 ) , .A1( us32_n827 ) );
  NOR4_X1 us32_U38 (.A3( us32_n755 ) , .A2( us32_n756 ) , .A1( us32_n757 ) , .ZN( us32_n758 ) , .A4( us32_n869 ) );
  NOR2_X1 us32_U380 (.A2( sa32_0 ) , .A1( sa32_1 ) , .ZN( us32_n462 ) );
  NOR2_X1 us32_U381 (.A2( sa32_3 ) , .ZN( us32_n455 ) , .A1( us32_n828 ) );
  NOR2_X1 us32_U382 (.A2( sa32_2 ) , .ZN( us32_n461 ) , .A1( us32_n829 ) );
  INV_X1 us32_U383 (.A( sa32_4 ) , .ZN( us32_n847 ) );
  INV_X1 us32_U384 (.A( sa32_6 ) , .ZN( us32_n849 ) );
  INV_X1 us32_U385 (.A( sa32_3 ) , .ZN( us32_n829 ) );
  INV_X1 us32_U386 (.A( sa32_1 ) , .ZN( us32_n827 ) );
  INV_X1 us32_U387 (.A( sa32_0 ) , .ZN( us32_n826 ) );
  INV_X1 us32_U388 (.A( sa32_2 ) , .ZN( us32_n828 ) );
  INV_X1 us32_U389 (.A( sa32_5 ) , .ZN( us32_n848 ) );
  AOI211_X1 us32_U39 (.B( us32_n745 ) , .A( us32_n746 ) , .ZN( us32_n759 ) , .C1( us32_n832 ) , .C2( us32_n853 ) );
  INV_X1 us32_U390 (.A( sa32_7 ) , .ZN( us32_n858 ) );
  NAND2_X1 us32_U391 (.A2( us32_n461 ) , .A1( us32_n471 ) , .ZN( us32_n697 ) );
  OAI222_X1 us32_U392 (.B2( us32_n747 ) , .B1( us32_n748 ) , .A2( us32_n749 ) , .ZN( us32_n757 ) , .C2( us32_n805 ) , .C1( us32_n814 ) , .A1( us32_n817 ) );
  OAI22_X1 us32_U393 (.B2( us32_n803 ) , .B1( us32_n804 ) , .A2( us32_n805 ) , .A1( us32_n806 ) , .ZN( us32_n808 ) );
  OAI21_X1 us32_U394 (.A( us32_n731 ) , .B1( us32_n732 ) , .ZN( us32_n736 ) , .B2( us32_n805 ) );
  OAI222_X1 us32_U395 (.ZN( us32_n505 ) , .C2( us32_n625 ) , .B2( us32_n647 ) , .B1( us32_n747 ) , .A2( us32_n748 ) , .C1( us32_n805 ) , .A1( us32_n806 ) );
  AOI21_X1 us32_U396 (.ZN( us32_n650 ) , .A( us32_n779 ) , .B1( us32_n792 ) , .B2( us32_n805 ) );
  INV_X1 us32_U397 (.A( us32_n805 ) , .ZN( us32_n860 ) );
  NOR2_X1 us32_U398 (.ZN( us32_n735 ) , .A2( us32_n803 ) , .A1( us32_n805 ) );
  NOR2_X1 us32_U399 (.ZN( us32_n484 ) , .A1( us32_n788 ) , .A2( us32_n805 ) );
  NAND2_X1 us32_U4 (.A1( us32_n441 ) , .A2( us32_n464 ) , .ZN( us32_n708 ) );
  NOR3_X1 us32_U40 (.A3( us32_n741 ) , .A2( us32_n742 ) , .A1( us32_n743 ) , .ZN( us32_n760 ) );
  NOR2_X1 us32_U400 (.A2( us32_n744 ) , .ZN( us32_n755 ) , .A1( us32_n805 ) );
  NAND2_X1 us32_U401 (.ZN( us32_n753 ) , .A1( us32_n763 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U402 (.ZN( us32_n715 ) , .A1( us32_n805 ) , .A2( us32_n817 ) );
  NOR2_X1 us32_U403 (.ZN( us32_n567 ) , .A1( us32_n747 ) , .A2( us32_n805 ) );
  AOI21_X1 us32_U404 (.ZN( us32_n552 ) , .B1( us32_n669 ) , .A( us32_n697 ) , .B2( us32_n805 ) );
  NOR2_X1 us32_U405 (.ZN( us32_n556 ) , .A1( us32_n762 ) , .A2( us32_n805 ) );
  NOR2_X1 us32_U406 (.ZN( us32_n670 ) , .A1( us32_n790 ) , .A2( us32_n805 ) );
  OAI221_X1 us32_U407 (.A( us32_n783 ) , .C2( us32_n784 ) , .B2( us32_n785 ) , .B1( us32_n786 ) , .ZN( us32_n796 ) , .C1( us32_n813 ) );
  NAND2_X1 us32_U408 (.A1( us32_n729 ) , .A2( us32_n784 ) , .ZN( us32_n811 ) );
  OAI22_X1 us32_U409 (.ZN( us32_n588 ) , .A2( us32_n747 ) , .B2( us32_n762 ) , .A1( us32_n763 ) , .B1( us32_n784 ) );
  NAND4_X1 us32_U41 (.ZN( sa33_sr_3 ) , .A4( us32_n704 ) , .A3( us32_n705 ) , .A2( us32_n706 ) , .A1( us32_n707 ) );
  AOI21_X1 us32_U410 (.ZN( us32_n592 ) , .B1( us32_n728 ) , .B2( us32_n784 ) , .A( us32_n790 ) );
  AOI21_X1 us32_U411 (.ZN( us32_n623 ) , .B1( us32_n699 ) , .A( us32_n779 ) , .B2( us32_n784 ) );
  AOI21_X1 us32_U412 (.ZN( us32_n648 ) , .A( us32_n762 ) , .B2( us32_n784 ) , .B1( us32_n792 ) );
  OAI22_X1 us32_U413 (.ZN( us32_n681 ) , .A1( us32_n699 ) , .A2( us32_n730 ) , .B2( us32_n784 ) , .B1( us32_n817 ) );
  OAI21_X1 us32_U414 (.A( us32_n613 ) , .ZN( us32_n616 ) , .B1( us32_n625 ) , .B2( us32_n784 ) );
  NOR2_X1 us32_U415 (.ZN( us32_n610 ) , .A1( us32_n784 ) , .A2( us32_n816 ) );
  OAI222_X1 us32_U416 (.A2( us32_n669 ) , .ZN( us32_n674 ) , .B1( us32_n747 ) , .B2( us32_n784 ) , .C2( us32_n788 ) , .C1( us32_n815 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U417 (.ZN( us32_n651 ) , .A1( us32_n784 ) , .A2( us32_n788 ) );
  NOR2_X1 us32_U418 (.ZN( us32_n600 ) , .A2( us32_n697 ) , .A1( us32_n784 ) );
  NOR2_X1 us32_U419 (.ZN( us32_n553 ) , .A2( us32_n744 ) , .A1( us32_n784 ) );
  NOR4_X1 us32_U42 (.A4( us32_n700 ) , .A3( us32_n701 ) , .A2( us32_n702 ) , .A1( us32_n703 ) , .ZN( us32_n704 ) );
  INV_X1 us32_U420 (.A( us32_n784 ) , .ZN( us32_n861 ) );
  AOI21_X1 us32_U421 (.ZN( us32_n500 ) , .A( us32_n697 ) , .B1( us32_n708 ) , .B2( us32_n786 ) );
  OAI221_X1 us32_U422 (.A( us32_n696 ) , .ZN( us32_n703 ) , .C2( us32_n784 ) , .C1( us32_n785 ) , .B1( us32_n786 ) , .B2( us32_n806 ) );
  OAI22_X1 us32_U423 (.ZN( us32_n590 ) , .B1( us32_n730 ) , .B2( us32_n749 ) , .A2( us32_n786 ) , .A1( us32_n803 ) );
  NOR2_X1 us32_U424 (.ZN( us32_n612 ) , .A1( us32_n779 ) , .A2( us32_n786 ) );
  NAND2_X1 us32_U425 (.A2( us32_n749 ) , .A1( us32_n786 ) , .ZN( us32_n809 ) );
  OAI222_X1 us32_U426 (.ZN( us32_n617 ) , .B1( us32_n697 ) , .C1( us32_n724 ) , .C2( us32_n747 ) , .B2( us32_n786 ) , .A2( us32_n792 ) , .A1( us32_n816 ) );
  NOR2_X1 us32_U427 (.ZN( us32_n717 ) , .A2( us32_n744 ) , .A1( us32_n786 ) );
  NOR2_X1 us32_U428 (.ZN( us32_n653 ) , .A1( us32_n762 ) , .A2( us32_n786 ) );
  NOR2_X1 us32_U429 (.ZN( us32_n554 ) , .A1( us32_n786 ) , .A2( us32_n813 ) );
  AOI211_X1 us32_U43 (.B( us32_n694 ) , .A( us32_n695 ) , .ZN( us32_n705 ) , .C2( us32_n831 ) , .C1( us32_n851 ) );
  NOR2_X1 us32_U430 (.ZN( us32_n701 ) , .A2( us32_n786 ) , .A1( us32_n817 ) );
  NOR2_X1 us32_U431 (.A1( us32_n730 ) , .ZN( us32_n765 ) , .A2( us32_n786 ) );
  AND2_X1 us32_U432 (.ZN( us32_n438 ) , .A2( us32_n831 ) , .A1( us32_n854 ) );
  AND2_X1 us32_U433 (.ZN( us32_n439 ) , .A2( us32_n843 ) , .A1( us32_n861 ) );
  NOR3_X1 us32_U434 (.A1( us32_n438 ) , .A2( us32_n439 ) , .A3( us32_n576 ) , .ZN( us32_n587 ) );
  NAND4_X1 us32_U435 (.ZN( sa33_sr_2 ) , .A4( us32_n643 ) , .A3( us32_n644 ) , .A2( us32_n645 ) , .A1( us32_n646 ) );
  INV_X1 us32_U436 (.A( us32_n812 ) , .ZN( us32_n854 ) );
  NAND3_X1 us32_U437 (.ZN( sa33_sr_6 ) , .A3( us32_n797 ) , .A2( us32_n798 ) , .A1( us32_n799 ) );
  NAND3_X1 us32_U438 (.ZN( sa33_sr_5 ) , .A3( us32_n758 ) , .A2( us32_n759 ) , .A1( us32_n760 ) );
  NAND3_X1 us32_U439 (.ZN( sa33_sr_4 ) , .A3( us32_n738 ) , .A2( us32_n739 ) , .A1( us32_n740 ) );
  NOR2_X1 us32_U44 (.ZN( us32_n707 ) , .A2( us32_n776 ) , .A1( us32_n800 ) );
  NAND3_X1 us32_U440 (.A3( us32_n675 ) , .A2( us32_n676 ) , .A1( us32_n677 ) , .ZN( us32_n807 ) );
  NAND3_X1 us32_U441 (.ZN( us32_n638 ) , .A3( us32_n708 ) , .A2( us32_n724 ) , .A1( us32_n792 ) );
  NAND3_X1 us32_U442 (.A3( us32_n618 ) , .A2( us32_n619 ) , .A1( us32_n620 ) , .ZN( us32_n725 ) );
  NAND3_X1 us32_U443 (.A3( us32_n585 ) , .A2( us32_n586 ) , .A1( us32_n587 ) , .ZN( us32_n621 ) );
  NAND3_X1 us32_U444 (.ZN( us32_n565 ) , .A3( us32_n680 ) , .A2( us32_n750 ) , .A1( us32_n785 ) );
  NAND3_X1 us32_U445 (.A3( us32_n523 ) , .A2( us32_n524 ) , .A1( us32_n525 ) , .ZN( us32_n742 ) );
  NAND3_X1 us32_U446 (.A3( us32_n512 ) , .A1( us32_n513 ) , .ZN( us32_n608 ) , .A2( us32_n871 ) );
  NAND3_X1 us32_U447 (.A3( us32_n467 ) , .A2( us32_n468 ) , .A1( us32_n469 ) , .ZN( us32_n777 ) );
  INV_X1 us32_U448 (.A( us32_n803 ) , .ZN( us32_n843 ) );
  AOI21_X1 us32_U449 (.ZN( us32_n576 ) , .B2( us32_n724 ) , .B1( us32_n748 ) , .A( us32_n785 ) );
  AOI222_X1 us32_U45 (.B2( us32_n638 ) , .ZN( us32_n644 ) , .B1( us32_n841 ) , .A1( us32_n842 ) , .C2( us32_n846 ) , .C1( us32_n863 ) , .A2( us32_n865 ) );
  NOR4_X1 us32_U46 (.A4( us32_n639 ) , .A3( us32_n640 ) , .A2( us32_n641 ) , .A1( us32_n642 ) , .ZN( us32_n643 ) );
  NOR3_X1 us32_U47 (.A2( us32_n607 ) , .A1( us32_n608 ) , .ZN( us32_n646 ) , .A3( us32_n722 ) );
  NAND4_X1 us32_U48 (.ZN( sa33_sr_7 ) , .A4( us32_n822 ) , .A3( us32_n823 ) , .A2( us32_n824 ) , .A1( us32_n825 ) );
  NOR4_X1 us32_U49 (.A4( us32_n818 ) , .A3( us32_n819 ) , .A2( us32_n820 ) , .A1( us32_n821 ) , .ZN( us32_n822 ) );
  NAND2_X1 us32_U5 (.A2( us32_n441 ) , .A1( us32_n452 ) , .ZN( us32_n791 ) );
  AOI222_X1 us32_U50 (.C2( us32_n809 ) , .B2( us32_n810 ) , .A2( us32_n811 ) , .ZN( us32_n823 ) , .C1( us32_n832 ) , .A1( us32_n839 ) , .B1( us32_n853 ) );
  AOI211_X1 us32_U51 (.B( us32_n807 ) , .A( us32_n808 ) , .ZN( us32_n824 ) , .C1( us32_n842 ) , .C2( us32_n850 ) );
  NAND4_X1 us32_U52 (.ZN( sa33_sr_0 ) , .A4( us32_n501 ) , .A3( us32_n502 ) , .A2( us32_n503 ) , .A1( us32_n504 ) );
  AOI221_X1 us32_U53 (.A( us32_n497 ) , .ZN( us32_n502 ) , .B2( us32_n843 ) , .C1( us32_n846 ) , .C2( us32_n860 ) , .B1( us32_n862 ) );
  NOR4_X1 us32_U54 (.A4( us32_n498 ) , .A3( us32_n499 ) , .A2( us32_n500 ) , .ZN( us32_n501 ) , .A1( us32_n527 ) );
  AOI211_X1 us32_U55 (.A( us32_n496 ) , .ZN( us32_n503 ) , .B( us32_n802 ) , .C2( us32_n839 ) , .C1( us32_n851 ) );
  NAND4_X1 us32_U56 (.ZN( sa33_sr_1 ) , .A4( us32_n595 ) , .A3( us32_n596 ) , .A2( us32_n597 ) , .A1( us32_n598 ) );
  NOR4_X1 us32_U57 (.A4( us32_n591 ) , .A3( us32_n592 ) , .A2( us32_n593 ) , .A1( us32_n594 ) , .ZN( us32_n595 ) );
  AOI211_X1 us32_U58 (.B( us32_n589 ) , .A( us32_n590 ) , .ZN( us32_n596 ) , .C2( us32_n811 ) , .C1( us32_n833 ) );
  AOI211_X1 us32_U59 (.A( us32_n588 ) , .ZN( us32_n597 ) , .B( us32_n621 ) , .C1( us32_n845 ) , .C2( us32_n855 ) );
  NOR3_X1 us32_U6 (.ZN( us32_n598 ) , .A1( us32_n608 ) , .A3( us32_n723 ) , .A2( us32_n742 ) );
  NOR2_X1 us32_U60 (.ZN( us32_n804 ) , .A1( us32_n854 ) , .A2( us32_n861 ) );
  AOI222_X1 us32_U61 (.ZN( us32_n469 ) , .B1( us32_n832 ) , .A1( us32_n839 ) , .C1( us32_n842 ) , .C2( us32_n851 ) , .A2( us32_n855 ) , .B2( us32_n865 ) );
  NOR4_X1 us32_U62 (.A1( us32_n466 ) , .ZN( us32_n467 ) , .A4( us32_n542 ) , .A2( us32_n554 ) , .A3( us32_n614 ) );
  AOI221_X1 us32_U63 (.ZN( us32_n468 ) , .C2( us32_n714 ) , .B2( us32_n831 ) , .C1( us32_n845 ) , .B1( us32_n860 ) , .A( us32_n864 ) );
  NAND4_X1 us32_U64 (.A4( us32_n603 ) , .A3( us32_n604 ) , .A2( us32_n605 ) , .A1( us32_n606 ) , .ZN( us32_n722 ) );
  NOR3_X1 us32_U65 (.A1( us32_n599 ) , .ZN( us32_n604 ) , .A3( us32_n663 ) , .A2( us32_n770 ) );
  NOR4_X1 us32_U66 (.A3( us32_n600 ) , .A2( us32_n601 ) , .A1( us32_n602 ) , .ZN( us32_n603 ) , .A4( us32_n655 ) );
  AOI222_X1 us32_U67 (.ZN( us32_n606 ) , .A1( us32_n830 ) , .C2( us32_n837 ) , .B1( us32_n842 ) , .A2( us32_n856 ) , .B2( us32_n861 ) , .C1( us32_n868 ) );
  NAND4_X1 us32_U68 (.A4( us32_n657 ) , .A3( us32_n658 ) , .A2( us32_n659 ) , .A1( us32_n660 ) , .ZN( us32_n800 ) );
  NOR3_X1 us32_U69 (.A3( us32_n648 ) , .A2( us32_n649 ) , .A1( us32_n650 ) , .ZN( us32_n659 ) );
  NOR3_X1 us32_U7 (.A3( us32_n800 ) , .A2( us32_n801 ) , .A1( us32_n802 ) , .ZN( us32_n825 ) );
  NOR3_X1 us32_U70 (.A3( us32_n651 ) , .A2( us32_n652 ) , .A1( us32_n653 ) , .ZN( us32_n658 ) );
  NOR3_X1 us32_U71 (.A3( us32_n654 ) , .A2( us32_n655 ) , .A1( us32_n656 ) , .ZN( us32_n657 ) );
  NAND4_X1 us32_U72 (.A4( us32_n560 ) , .A3( us32_n561 ) , .A2( us32_n562 ) , .A1( us32_n563 ) , .ZN( us32_n607 ) );
  NOR4_X1 us32_U73 (.A4( us32_n556 ) , .A3( us32_n557 ) , .A2( us32_n558 ) , .A1( us32_n559 ) , .ZN( us32_n560 ) );
  NOR4_X1 us32_U74 (.ZN( us32_n561 ) , .A1( us32_n653 ) , .A3( us32_n661 ) , .A4( us32_n685 ) , .A2( us32_n768 ) );
  NOR4_X1 us32_U75 (.A4( us32_n552 ) , .A3( us32_n553 ) , .A2( us32_n554 ) , .A1( us32_n555 ) , .ZN( us32_n562 ) );
  NAND4_X1 us32_U76 (.A4( us32_n772 ) , .A3( us32_n773 ) , .A2( us32_n774 ) , .A1( us32_n775 ) , .ZN( us32_n801 ) );
  NOR3_X1 us32_U77 (.A3( us32_n765 ) , .A2( us32_n766 ) , .A1( us32_n767 ) , .ZN( us32_n773 ) );
  NOR4_X1 us32_U78 (.A4( us32_n768 ) , .A3( us32_n769 ) , .A2( us32_n770 ) , .A1( us32_n771 ) , .ZN( us32_n772 ) );
  AOI222_X1 us32_U79 (.ZN( us32_n775 ) , .A1( us32_n830 ) , .C1( us32_n834 ) , .B2( us32_n841 ) , .A2( us32_n850 ) , .B1( us32_n861 ) , .C2( us32_n873 ) );
  NOR3_X1 us32_U8 (.A3( us32_n621 ) , .A2( us32_n622 ) , .ZN( us32_n636 ) , .A1( us32_n725 ) );
  NOR4_X1 us32_U80 (.A4( us32_n665 ) , .A3( us32_n666 ) , .A2( us32_n667 ) , .A1( us32_n668 ) , .ZN( us32_n676 ) );
  NOR4_X1 us32_U81 (.A4( us32_n661 ) , .A3( us32_n662 ) , .A2( us32_n663 ) , .A1( us32_n664 ) , .ZN( us32_n677 ) );
  NOR4_X1 us32_U82 (.A3( us32_n673 ) , .A1( us32_n674 ) , .ZN( us32_n675 ) , .A4( us32_n715 ) , .A2( us32_n859 ) );
  NOR2_X1 us32_U83 (.ZN( us32_n625 ) , .A2( us32_n836 ) , .A1( us32_n839 ) );
  NOR2_X1 us32_U84 (.ZN( us32_n761 ) , .A1( us32_n833 ) , .A2( us32_n834 ) );
  NOR4_X1 us32_U85 (.A4( us32_n577 ) , .A3( us32_n578 ) , .A2( us32_n579 ) , .ZN( us32_n586 ) , .A1( us32_n683 ) );
  NOR4_X1 us32_U86 (.A1( us32_n584 ) , .ZN( us32_n585 ) , .A3( us32_n652 ) , .A2( us32_n662 ) , .A4( us32_n767 ) );
  AOI222_X1 us32_U87 (.ZN( us32_n513 ) , .C1( us32_n832 ) , .B2( us32_n837 ) , .A2( us32_n843 ) , .C2( us32_n862 ) , .B1( us32_n863 ) , .A1( us32_n866 ) );
  NOR4_X1 us32_U88 (.A4( us32_n509 ) , .A2( us32_n510 ) , .A1( us32_n511 ) , .ZN( us32_n512 ) , .A3( us32_n670 ) );
  INV_X1 us32_U89 (.A( us32_n505 ) , .ZN( us32_n871 ) );
  NOR2_X1 us32_U9 (.ZN( us32_n495 ) , .A1( us32_n678 ) , .A2( us32_n694 ) );
  NAND4_X1 us32_U90 (.A4( us32_n456 ) , .A3( us32_n457 ) , .A2( us32_n458 ) , .A1( us32_n459 ) , .ZN( us32_n679 ) );
  NOR3_X1 us32_U91 (.ZN( us32_n457 ) , .A3( us32_n530 ) , .A1( us32_n555 ) , .A2( us32_n570 ) );
  AOI221_X1 us32_U92 (.A( us32_n450 ) , .ZN( us32_n459 ) , .C2( us32_n753 ) , .B1( us32_n832 ) , .C1( us32_n842 ) , .B2( us32_n861 ) );
  NOR4_X1 us32_U93 (.ZN( us32_n458 ) , .A2( us32_n509 ) , .A1( us32_n599 ) , .A4( us32_n628 ) , .A3( us32_n711 ) );
  NAND4_X1 us32_U94 (.A4( us32_n535 ) , .A3( us32_n536 ) , .A2( us32_n537 ) , .A1( us32_n538 ) , .ZN( us32_n622 ) );
  NOR4_X1 us32_U95 (.A4( us32_n526 ) , .A2( us32_n527 ) , .A1( us32_n528 ) , .ZN( us32_n538 ) , .A3( us32_n701 ) );
  NOR4_X1 us32_U96 (.A1( us32_n531 ) , .ZN( us32_n536 ) , .A2( us32_n654 ) , .A4( us32_n668 ) , .A3( us32_n765 ) );
  NOR4_X1 us32_U97 (.A4( us32_n529 ) , .A3( us32_n530 ) , .ZN( us32_n537 ) , .A2( us32_n684 ) , .A1( us32_n794 ) );
  NAND4_X1 us32_U98 (.A4( us32_n479 ) , .A3( us32_n480 ) , .A2( us32_n481 ) , .A1( us32_n482 ) , .ZN( us32_n694 ) );
  NOR3_X1 us32_U99 (.ZN( us32_n480 ) , .A2( us32_n508 ) , .A3( us32_n601 ) , .A1( us32_n610 ) );
endmodule

