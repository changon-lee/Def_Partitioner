module des_des_die_5 ( u0_FP_40, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_47, u0_FP_48, 
       u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_K11_37, u0_K12_39, u0_K12_40, u0_K12_7, 
       u0_K12_9, u0_K16_18, u0_K16_19, u0_K16_22, u0_K16_24, u0_K16_26, u0_K2_11, u0_K2_12, u0_K2_4, 
       u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_10, u0_K3_12, u0_K3_14, u0_K3_15, u0_K3_17, u0_K3_18, 
       u0_K3_19, u0_K3_23, u0_K3_34, u0_K3_5, u0_K4_35, u0_K7_2, u0_L0_12, u0_L0_13, u0_L0_16, 
       u0_L0_17, u0_L0_18, u0_L0_2, u0_L0_22, u0_L0_23, u0_L0_24, u0_L0_28, u0_L0_30, u0_L0_31, 
       u0_L0_32, u0_L0_6, u0_L0_7, u0_L0_9, u0_L10_12, u0_L10_13, u0_L10_16, u0_L10_18, u0_L10_2, 
       u0_L10_22, u0_L10_24, u0_L10_28, u0_L10_30, u0_L10_32, u0_L10_6, u0_L10_7, u0_L14_1, u0_L14_10, 
       u0_L14_14, u0_L14_16, u0_L14_20, u0_L14_24, u0_L14_25, u0_L14_26, u0_L14_3, u0_L14_30, u0_L14_6, 
       u0_L14_8, u0_L1_1, u0_L1_10, u0_L1_11, u0_L1_13, u0_L1_16, u0_L1_17, u0_L1_18, u0_L1_19, 
       u0_L1_2, u0_L1_20, u0_L1_23, u0_L1_24, u0_L1_26, u0_L1_28, u0_L1_29, u0_L1_30, u0_L1_31, 
       u0_L1_4, u0_L1_6, u0_L1_9, u0_L2_11, u0_L2_19, u0_L2_29, u0_L2_4, u0_L5_11, u0_L5_12, 
       u0_L5_15, u0_L5_17, u0_L5_19, u0_L5_21, u0_L5_22, u0_L5_23, u0_L5_27, u0_L5_29, u0_L5_31, 
       u0_L5_32, u0_L5_4, u0_L5_5, u0_L5_7, u0_L5_9, u0_L8_17, u0_L8_23, u0_L8_31, u0_L8_9, 
       u0_L9_11, u0_L9_12, u0_L9_13, u0_L9_17, u0_L9_18, u0_L9_19, u0_L9_2, u0_L9_22, u0_L9_23, 
       u0_L9_28, u0_L9_29, u0_L9_31, u0_L9_32, u0_L9_4, u0_L9_7, u0_L9_9, u0_R0_1, u0_R0_10, 
       u0_R0_11, u0_R0_12, u0_R0_13, u0_R0_2, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, u0_R0_28, 
       u0_R0_29, u0_R0_3, u0_R0_32, u0_R0_4, u0_R0_5, u0_R0_6, u0_R0_7, u0_R0_8, u0_R0_9, 
       u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_24, u0_R10_25, u0_R10_26, u0_R10_27, u0_R10_28, 
       u0_R10_29, u0_R10_4, u0_R10_5, u0_R10_6, u0_R10_7, u0_R10_8, u0_R10_9, u0_R1_1, u0_R1_10, 
       u0_R1_11, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, u0_R1_17, u0_R1_2, u0_R1_20, 
       u0_R1_21, u0_R1_22, u0_R1_23, u0_R1_24, u0_R1_25, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, 
       u0_R1_6, u0_R1_7, u0_R1_8, u0_R1_9, u0_R2_20, u0_R2_21, u0_R2_22, u0_R2_23, u0_R2_24, 
       u0_R2_25, u0_R5_1, u0_R5_2, u0_R5_20, u0_R5_21, u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, 
       u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, 
       u0_R8_1, u0_R8_2, u0_R8_3, u0_R8_32, u0_R8_4, u0_R8_5, u0_R9_1, u0_R9_2, u0_R9_20, 
       u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_28, u0_R9_29, 
       u0_R9_3, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_u6_X_6, 
       u0_uk_K_r0_11, u0_uk_K_r0_19, u0_uk_K_r0_22, u0_uk_K_r0_25, u0_uk_K_r0_28, u0_uk_K_r0_32, u0_uk_K_r0_34, u0_uk_K_r0_49, u0_uk_K_r0_55, 
       u0_uk_K_r10_18, u0_uk_K_r10_25, u0_uk_K_r10_28, u0_uk_K_r10_34, u0_uk_K_r10_41, u0_uk_K_r10_9, u0_uk_K_r14_10, u0_uk_K_r14_18, u0_uk_K_r14_45, 
       u0_uk_K_r14_46, u0_uk_K_r14_8, u0_uk_K_r1_10, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_41, u0_uk_K_r1_47, u0_uk_K_r1_7, u0_uk_K_r2_29, 
       u0_uk_K_r5_0, u0_uk_K_r5_1, u0_uk_K_r5_10, u0_uk_K_r5_16, u0_uk_K_r5_21, u0_uk_K_r5_37, u0_uk_K_r5_5, u0_uk_K_r5_51, u0_uk_K_r5_8, 
       u0_uk_K_r8_41, u0_uk_K_r9_12, u0_uk_K_r9_18, u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_25, u0_uk_K_r9_30, u0_uk_K_r9_31, u0_uk_K_r9_33, 
       u0_uk_K_r9_45, u0_uk_K_r9_49, u0_uk_K_r9_6, u0_uk_K_r9_7, u0_uk_n10, u0_uk_n1004, u0_uk_n102, u0_uk_n1021, u0_uk_n11, 
       u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n141, u0_uk_n144, u0_uk_n145, 
       u0_uk_n149, u0_uk_n153, u0_uk_n157, u0_uk_n161, u0_uk_n162, u0_uk_n165, u0_uk_n169, u0_uk_n170, u0_uk_n175, 
       u0_uk_n177, u0_uk_n179, u0_uk_n180, u0_uk_n181, u0_uk_n182, u0_uk_n183, u0_uk_n185, u0_uk_n186, u0_uk_n187, 
       u0_uk_n188, u0_uk_n189, u0_uk_n193, u0_uk_n194, u0_uk_n195, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n200, 
       u0_uk_n201, u0_uk_n202, u0_uk_n205, u0_uk_n206, u0_uk_n207, u0_uk_n209, u0_uk_n210, u0_uk_n212, u0_uk_n213, 
       u0_uk_n215, u0_uk_n216, u0_uk_n218, u0_uk_n219, u0_uk_n223, u0_uk_n224, u0_uk_n225, u0_uk_n227, u0_uk_n235, 
       u0_uk_n238, u0_uk_n239, u0_uk_n242, u0_uk_n246, u0_uk_n255, u0_uk_n257, u0_uk_n258, u0_uk_n263, u0_uk_n266, 
       u0_uk_n267, u0_uk_n31, u0_uk_n361, u0_uk_n365, u0_uk_n367, u0_uk_n371, u0_uk_n372, u0_uk_n374, u0_uk_n378, 
       u0_uk_n380, u0_uk_n381, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n393, u0_uk_n394, u0_uk_n396, 
       u0_uk_n398, u0_uk_n399, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n406, u0_uk_n506, u0_uk_n507, u0_uk_n508, 
       u0_uk_n512, u0_uk_n522, u0_uk_n532, u0_uk_n539, u0_uk_n540, u0_uk_n542, u0_uk_n544, u0_uk_n545, u0_uk_n547, 
       u0_uk_n549, u0_uk_n552, u0_uk_n555, u0_uk_n557, u0_uk_n562, u0_uk_n563, u0_uk_n564, u0_uk_n565, u0_uk_n566, 
       u0_uk_n567, u0_uk_n568, u0_uk_n569, u0_uk_n571, u0_uk_n573, u0_uk_n576, u0_uk_n577, u0_uk_n578, u0_uk_n579, 
       u0_uk_n580, u0_uk_n583, u0_uk_n584, u0_uk_n588, u0_uk_n592, u0_uk_n593, u0_uk_n594, u0_uk_n596, u0_uk_n597, 
       u0_uk_n598, u0_uk_n60, u0_uk_n604, u0_uk_n607, u0_uk_n611, u0_uk_n612, u0_uk_n614, u0_uk_n615, u0_uk_n619, 
       u0_uk_n621, u0_uk_n622, u0_uk_n623, u0_uk_n626, u0_uk_n627, u0_uk_n629, u0_uk_n63, u0_uk_n631, u0_uk_n632, 
       u0_uk_n636, u0_uk_n640, u0_uk_n642, u0_uk_n644, u0_uk_n645, u0_uk_n649, u0_uk_n651, u0_uk_n652, u0_uk_n653, 
       u0_uk_n654, u0_uk_n658, u0_uk_n661, u0_uk_n663, u0_uk_n669, u0_uk_n765, u0_uk_n766, u0_uk_n770, u0_uk_n826, 
       u0_uk_n853, u0_uk_n855, u0_uk_n904, u0_uk_n92, u0_uk_n981, u0_uk_n99, u0_uk_n990, u1_FP_62, u1_FP_63, 
       u1_K13_16, u1_K13_33, u1_K13_34, u1_K13_9, u1_K14_15, u1_K14_16, u1_K14_3, u1_K14_4, u1_K15_10, 
       u1_K15_9, u1_K16_45, u1_K16_46, u1_K2_33, u1_K2_34, u1_K3_27, u1_K3_28, u1_K3_3, u1_K3_4, 
       u1_K4_15, u1_K4_16, u1_K4_27, u1_K4_28, u1_K4_30, u1_K4_32, u1_K4_33, u1_K4_34, u1_K4_45, 
       u1_K4_46, u1_K8_33, u1_L0_11, u1_L0_19, u1_L0_29, u1_L0_4, u1_L11_11, u1_L11_13, u1_L11_16, 
       u1_L11_18, u1_L11_19, u1_L11_2, u1_L11_24, u1_L11_28, u1_L11_29, u1_L11_30, u1_L11_4, u1_L11_6, 
       u1_L12_16, u1_L12_17, u1_L12_23, u1_L12_24, u1_L12_30, u1_L12_31, u1_L12_6, u1_L12_9, u1_L13_13, 
       u1_L13_18, u1_L13_2, u1_L13_28, u1_L14_15, u1_L14_21, u1_L14_27, u1_L14_5, u1_L1_14, u1_L1_17, 
       u1_L1_23, u1_L1_25, u1_L1_3, u1_L1_31, u1_L1_8, u1_L1_9, u1_L2_11, u1_L2_14, u1_L2_15, 
       u1_L2_16, u1_L2_19, u1_L2_21, u1_L2_24, u1_L2_25, u1_L2_27, u1_L2_29, u1_L2_3, u1_L2_30, 
       u1_L2_4, u1_L2_5, u1_L2_6, u1_L2_8, u1_L4_13, u1_L4_18, u1_L4_2, u1_L4_28, u1_L6_11, 
       u1_L6_19, u1_L6_29, u1_L6_4, u1_R0_22, u1_R0_23, u1_R11_10, u1_R11_11, u1_R11_22, u1_R11_23, 
       u1_R11_6, u1_R11_7, u1_R11_8, u1_R12_10, u1_R12_11, u1_R12_2, u1_R12_3, u1_R13_6, u1_R13_7, 
       u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_3, u1_R2_10, u1_R2_11, u1_R2_18, u1_R2_19, u1_R2_20, 
       u1_R2_21, u1_R2_22, u1_R2_23, u1_R2_30, u1_R2_31, u1_R4_6, u1_R4_7, u1_R6_22, u1_R6_23, 
       u1_u12_X_12, u1_u12_X_14, u1_u12_X_17, u1_u12_X_18, u1_u12_X_31, u1_u12_X_32, u1_u12_X_35, u1_u12_X_36, u1_u12_X_7, 
       u1_u12_X_8, u1_u13_X_1, u1_u13_X_13, u1_u13_X_14, u1_u13_X_17, u1_u13_X_18, u1_u13_X_2, u1_u13_X_5, u1_u13_X_6, 
       u1_u14_X_11, u1_u14_X_12, u1_u14_X_7, u1_u14_X_8, u1_u15_X_43, u1_u15_X_44, u1_u15_X_47, u1_u15_X_48, u1_u1_X_31, 
       u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u2_X_1, u1_u2_X_2, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, 
       u1_u2_X_5, u1_u2_X_6, u1_u3_X_13, u1_u3_X_14, u1_u3_X_17, u1_u3_X_18, u1_u3_X_25, u1_u3_X_26, u1_u3_X_35, 
       u1_u3_X_36, u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, u1_u3_X_48, u1_u5_X_11, u1_u5_X_12, u1_u5_X_7, u1_u5_X_8, 
       u1_u7_X_31, u1_u7_X_32, u1_u7_X_35, u1_u7_X_36, u1_uk_n1060, u1_uk_n1063, u1_uk_n1088, u1_uk_n1104, u1_uk_n1137, 
       u1_uk_n671, u1_uk_n672, u1_uk_n677, u1_uk_n678, u2_K6_13, u2_K6_14, u2_K6_15, u2_K6_16, u2_K8_5, 
       u2_L4_16, u2_L4_24, u2_L4_30, u2_L4_6, u2_L6_17, u2_L6_23, u2_L6_31, u2_L6_9, u2_R4_10, 
       u2_R4_11, u2_R4_12, u2_R4_13, u2_R4_8, u2_R4_9, u2_R6_1, u2_R6_2, u2_R6_3, u2_R6_32, 
       u2_R6_4, u2_R6_5, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_4, u2_uk_K_r4_55, u2_uk_K_r6_10, u2_uk_K_r6_3, u2_uk_n100, 
       u2_uk_n102, u2_uk_n1105, u2_uk_n1116, u2_uk_n117, u2_uk_n118, u2_uk_n147, u2_uk_n1502, u2_uk_n1507, u2_uk_n1514, 
       u2_uk_n1515, u2_uk_n1518, u2_uk_n1519, u2_uk_n155, u2_uk_n162, u2_uk_n182, u2_uk_n188, u2_uk_n27, u2_uk_n83, u0_FP_1, u0_FP_10, u0_FP_14, u0_FP_16, u0_FP_20, u0_FP_24, u0_FP_25, u0_FP_26, u0_FP_3, 
        u0_FP_30, u0_FP_6, u0_FP_8, u0_N106, u0_N114, u0_N124, u0_N195, u0_N196, u0_N198, 
        u0_N200, u0_N202, u0_N203, u0_N206, u0_N208, u0_N210, u0_N212, u0_N213, u0_N214, 
        u0_N218, u0_N220, u0_N222, u0_N223, u0_N296, u0_N304, u0_N310, u0_N318, u0_N321, 
        u0_N323, u0_N326, u0_N328, u0_N33, u0_N330, u0_N331, u0_N332, u0_N336, u0_N337, 
        u0_N338, u0_N341, u0_N342, u0_N347, u0_N348, u0_N350, u0_N351, u0_N353, u0_N357, 
        u0_N358, u0_N363, u0_N364, u0_N367, u0_N369, u0_N37, u0_N373, u0_N375, u0_N379, 
        u0_N38, u0_N381, u0_N383, u0_N40, u0_N43, u0_N44, u0_N47, u0_N48, u0_N49, 
        u0_N53, u0_N54, u0_N55, u0_N59, u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, 
        u0_N67, u0_N69, u0_N72, u0_N73, u0_N74, u0_N76, u0_N79, u0_N80, u0_N81, 
        u0_N82, u0_N83, u0_N86, u0_N87, u0_N89, u0_N91, u0_N92, u0_N93, u0_N94, 
        u0_N99, u0_uk_n100, u0_uk_n109, u0_uk_n110, u0_uk_n129, u0_uk_n142, u0_uk_n146, u0_uk_n147, u0_uk_n148, 
        u0_uk_n155, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n191, u0_uk_n203, u0_uk_n208, u0_uk_n214, u0_uk_n217, 
        u0_uk_n220, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n240, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n778, 
        u0_uk_n823, u0_uk_n83, u0_uk_n841, u0_uk_n863, u0_uk_n867, u0_uk_n93, u0_uk_n94, u1_FP_15, u1_FP_21, 
        u1_FP_27, u1_FP_5, u1_N100, u1_N101, u1_N103, u1_N106, u1_N109, u1_N110, u1_N111, 
        u1_N114, u1_N116, u1_N119, u1_N120, u1_N122, u1_N124, u1_N125, u1_N161, u1_N172, 
        u1_N177, u1_N187, u1_N227, u1_N234, u1_N242, u1_N252, u1_N35, u1_N385, u1_N387, 
        u1_N389, u1_N394, u1_N396, u1_N399, u1_N401, u1_N402, u1_N407, u1_N411, u1_N412, 
        u1_N413, u1_N42, u1_N421, u1_N424, u1_N431, u1_N432, u1_N438, u1_N439, u1_N445, 
        u1_N446, u1_N449, u1_N460, u1_N465, u1_N475, u1_N50, u1_N60, u1_N66, u1_N71, 
        u1_N72, u1_N77, u1_N80, u1_N86, u1_N88, u1_N94, u1_N98, u1_N99, u2_N165, 
        u2_N175, u2_N183, u2_N189, u2_N232, u2_N240, u2_N246, u2_N254 );
  input u0_FP_40, u0_FP_41, u0_FP_42, u0_FP_43, u0_FP_44, u0_FP_45, u0_FP_46, u0_FP_47, u0_FP_48, 
        u0_FP_49, u0_FP_50, u0_FP_51, u0_FP_52, u0_FP_53, u0_K11_37, u0_K12_39, u0_K12_40, u0_K12_7, 
        u0_K12_9, u0_K16_18, u0_K16_19, u0_K16_22, u0_K16_24, u0_K16_26, u0_K2_11, u0_K2_12, u0_K2_4, 
        u0_K2_5, u0_K2_6, u0_K2_8, u0_K3_10, u0_K3_12, u0_K3_14, u0_K3_15, u0_K3_17, u0_K3_18, 
        u0_K3_19, u0_K3_23, u0_K3_34, u0_K3_5, u0_K4_35, u0_K7_2, u0_L0_12, u0_L0_13, u0_L0_16, 
        u0_L0_17, u0_L0_18, u0_L0_2, u0_L0_22, u0_L0_23, u0_L0_24, u0_L0_28, u0_L0_30, u0_L0_31, 
        u0_L0_32, u0_L0_6, u0_L0_7, u0_L0_9, u0_L10_12, u0_L10_13, u0_L10_16, u0_L10_18, u0_L10_2, 
        u0_L10_22, u0_L10_24, u0_L10_28, u0_L10_30, u0_L10_32, u0_L10_6, u0_L10_7, u0_L14_1, u0_L14_10, 
        u0_L14_14, u0_L14_16, u0_L14_20, u0_L14_24, u0_L14_25, u0_L14_26, u0_L14_3, u0_L14_30, u0_L14_6, 
        u0_L14_8, u0_L1_1, u0_L1_10, u0_L1_11, u0_L1_13, u0_L1_16, u0_L1_17, u0_L1_18, u0_L1_19, 
        u0_L1_2, u0_L1_20, u0_L1_23, u0_L1_24, u0_L1_26, u0_L1_28, u0_L1_29, u0_L1_30, u0_L1_31, 
        u0_L1_4, u0_L1_6, u0_L1_9, u0_L2_11, u0_L2_19, u0_L2_29, u0_L2_4, u0_L5_11, u0_L5_12, 
        u0_L5_15, u0_L5_17, u0_L5_19, u0_L5_21, u0_L5_22, u0_L5_23, u0_L5_27, u0_L5_29, u0_L5_31, 
        u0_L5_32, u0_L5_4, u0_L5_5, u0_L5_7, u0_L5_9, u0_L8_17, u0_L8_23, u0_L8_31, u0_L8_9, 
        u0_L9_11, u0_L9_12, u0_L9_13, u0_L9_17, u0_L9_18, u0_L9_19, u0_L9_2, u0_L9_22, u0_L9_23, 
        u0_L9_28, u0_L9_29, u0_L9_31, u0_L9_32, u0_L9_4, u0_L9_7, u0_L9_9, u0_R0_1, u0_R0_10, 
        u0_R0_11, u0_R0_12, u0_R0_13, u0_R0_2, u0_R0_24, u0_R0_25, u0_R0_26, u0_R0_27, u0_R0_28, 
        u0_R0_29, u0_R0_3, u0_R0_32, u0_R0_4, u0_R0_5, u0_R0_6, u0_R0_7, u0_R0_8, u0_R0_9, 
        u0_R10_10, u0_R10_11, u0_R10_12, u0_R10_13, u0_R10_24, u0_R10_25, u0_R10_26, u0_R10_27, u0_R10_28, 
        u0_R10_29, u0_R10_4, u0_R10_5, u0_R10_6, u0_R10_7, u0_R10_8, u0_R10_9, u0_R1_1, u0_R1_10, 
        u0_R1_11, u0_R1_12, u0_R1_13, u0_R1_14, u0_R1_15, u0_R1_16, u0_R1_17, u0_R1_2, u0_R1_20, 
        u0_R1_21, u0_R1_22, u0_R1_23, u0_R1_24, u0_R1_25, u0_R1_3, u0_R1_32, u0_R1_4, u0_R1_5, 
        u0_R1_6, u0_R1_7, u0_R1_8, u0_R1_9, u0_R2_20, u0_R2_21, u0_R2_22, u0_R2_23, u0_R2_24, 
        u0_R2_25, u0_R5_1, u0_R5_2, u0_R5_20, u0_R5_21, u0_R5_22, u0_R5_23, u0_R5_24, u0_R5_25, 
        u0_R5_26, u0_R5_27, u0_R5_28, u0_R5_29, u0_R5_3, u0_R5_30, u0_R5_31, u0_R5_32, u0_R5_4, 
        u0_R8_1, u0_R8_2, u0_R8_3, u0_R8_32, u0_R8_4, u0_R8_5, u0_R9_1, u0_R9_2, u0_R9_20, 
        u0_R9_21, u0_R9_22, u0_R9_23, u0_R9_24, u0_R9_25, u0_R9_26, u0_R9_27, u0_R9_28, u0_R9_29, 
        u0_R9_3, u0_R9_32, u0_R9_4, u0_R9_5, u0_R9_6, u0_R9_7, u0_R9_8, u0_R9_9, u0_u6_X_6, 
        u0_uk_K_r0_11, u0_uk_K_r0_19, u0_uk_K_r0_22, u0_uk_K_r0_25, u0_uk_K_r0_28, u0_uk_K_r0_32, u0_uk_K_r0_34, u0_uk_K_r0_49, u0_uk_K_r0_55, 
        u0_uk_K_r10_18, u0_uk_K_r10_25, u0_uk_K_r10_28, u0_uk_K_r10_34, u0_uk_K_r10_41, u0_uk_K_r10_9, u0_uk_K_r14_10, u0_uk_K_r14_18, u0_uk_K_r14_45, 
        u0_uk_K_r14_46, u0_uk_K_r14_8, u0_uk_K_r1_10, u0_uk_K_r1_17, u0_uk_K_r1_18, u0_uk_K_r1_41, u0_uk_K_r1_47, u0_uk_K_r1_7, u0_uk_K_r2_29, 
        u0_uk_K_r5_0, u0_uk_K_r5_1, u0_uk_K_r5_10, u0_uk_K_r5_16, u0_uk_K_r5_21, u0_uk_K_r5_37, u0_uk_K_r5_5, u0_uk_K_r5_51, u0_uk_K_r5_8, 
        u0_uk_K_r8_41, u0_uk_K_r9_12, u0_uk_K_r9_18, u0_uk_K_r9_19, u0_uk_K_r9_22, u0_uk_K_r9_25, u0_uk_K_r9_30, u0_uk_K_r9_31, u0_uk_K_r9_33, 
        u0_uk_K_r9_45, u0_uk_K_r9_49, u0_uk_K_r9_6, u0_uk_K_r9_7, u0_uk_n10, u0_uk_n1004, u0_uk_n102, u0_uk_n1021, u0_uk_n11, 
        u0_uk_n117, u0_uk_n118, u0_uk_n128, u0_uk_n136, u0_uk_n137, u0_uk_n139, u0_uk_n141, u0_uk_n144, u0_uk_n145, 
        u0_uk_n149, u0_uk_n153, u0_uk_n157, u0_uk_n161, u0_uk_n162, u0_uk_n165, u0_uk_n169, u0_uk_n170, u0_uk_n175, 
        u0_uk_n177, u0_uk_n179, u0_uk_n180, u0_uk_n181, u0_uk_n182, u0_uk_n183, u0_uk_n185, u0_uk_n186, u0_uk_n187, 
        u0_uk_n188, u0_uk_n189, u0_uk_n193, u0_uk_n194, u0_uk_n195, u0_uk_n197, u0_uk_n198, u0_uk_n199, u0_uk_n200, 
        u0_uk_n201, u0_uk_n202, u0_uk_n205, u0_uk_n206, u0_uk_n207, u0_uk_n209, u0_uk_n210, u0_uk_n212, u0_uk_n213, 
        u0_uk_n215, u0_uk_n216, u0_uk_n218, u0_uk_n219, u0_uk_n223, u0_uk_n224, u0_uk_n225, u0_uk_n227, u0_uk_n235, 
        u0_uk_n238, u0_uk_n239, u0_uk_n242, u0_uk_n246, u0_uk_n255, u0_uk_n257, u0_uk_n258, u0_uk_n263, u0_uk_n266, 
        u0_uk_n267, u0_uk_n31, u0_uk_n361, u0_uk_n365, u0_uk_n367, u0_uk_n371, u0_uk_n372, u0_uk_n374, u0_uk_n378, 
        u0_uk_n380, u0_uk_n381, u0_uk_n384, u0_uk_n387, u0_uk_n388, u0_uk_n389, u0_uk_n393, u0_uk_n394, u0_uk_n396, 
        u0_uk_n398, u0_uk_n399, u0_uk_n401, u0_uk_n402, u0_uk_n403, u0_uk_n406, u0_uk_n506, u0_uk_n507, u0_uk_n508, 
        u0_uk_n512, u0_uk_n522, u0_uk_n532, u0_uk_n539, u0_uk_n540, u0_uk_n542, u0_uk_n544, u0_uk_n545, u0_uk_n547, 
        u0_uk_n549, u0_uk_n552, u0_uk_n555, u0_uk_n557, u0_uk_n562, u0_uk_n563, u0_uk_n564, u0_uk_n565, u0_uk_n566, 
        u0_uk_n567, u0_uk_n568, u0_uk_n569, u0_uk_n571, u0_uk_n573, u0_uk_n576, u0_uk_n577, u0_uk_n578, u0_uk_n579, 
        u0_uk_n580, u0_uk_n583, u0_uk_n584, u0_uk_n588, u0_uk_n592, u0_uk_n593, u0_uk_n594, u0_uk_n596, u0_uk_n597, 
        u0_uk_n598, u0_uk_n60, u0_uk_n604, u0_uk_n607, u0_uk_n611, u0_uk_n612, u0_uk_n614, u0_uk_n615, u0_uk_n619, 
        u0_uk_n621, u0_uk_n622, u0_uk_n623, u0_uk_n626, u0_uk_n627, u0_uk_n629, u0_uk_n63, u0_uk_n631, u0_uk_n632, 
        u0_uk_n636, u0_uk_n640, u0_uk_n642, u0_uk_n644, u0_uk_n645, u0_uk_n649, u0_uk_n651, u0_uk_n652, u0_uk_n653, 
        u0_uk_n654, u0_uk_n658, u0_uk_n661, u0_uk_n663, u0_uk_n669, u0_uk_n765, u0_uk_n766, u0_uk_n770, u0_uk_n826, 
        u0_uk_n853, u0_uk_n855, u0_uk_n904, u0_uk_n92, u0_uk_n981, u0_uk_n99, u0_uk_n990, u1_FP_62, u1_FP_63, 
        u1_K13_16, u1_K13_33, u1_K13_34, u1_K13_9, u1_K14_15, u1_K14_16, u1_K14_3, u1_K14_4, u1_K15_10, 
        u1_K15_9, u1_K16_45, u1_K16_46, u1_K2_33, u1_K2_34, u1_K3_27, u1_K3_28, u1_K3_3, u1_K3_4, 
        u1_K4_15, u1_K4_16, u1_K4_27, u1_K4_28, u1_K4_30, u1_K4_32, u1_K4_33, u1_K4_34, u1_K4_45, 
        u1_K4_46, u1_K8_33, u1_L0_11, u1_L0_19, u1_L0_29, u1_L0_4, u1_L11_11, u1_L11_13, u1_L11_16, 
        u1_L11_18, u1_L11_19, u1_L11_2, u1_L11_24, u1_L11_28, u1_L11_29, u1_L11_30, u1_L11_4, u1_L11_6, 
        u1_L12_16, u1_L12_17, u1_L12_23, u1_L12_24, u1_L12_30, u1_L12_31, u1_L12_6, u1_L12_9, u1_L13_13, 
        u1_L13_18, u1_L13_2, u1_L13_28, u1_L14_15, u1_L14_21, u1_L14_27, u1_L14_5, u1_L1_14, u1_L1_17, 
        u1_L1_23, u1_L1_25, u1_L1_3, u1_L1_31, u1_L1_8, u1_L1_9, u1_L2_11, u1_L2_14, u1_L2_15, 
        u1_L2_16, u1_L2_19, u1_L2_21, u1_L2_24, u1_L2_25, u1_L2_27, u1_L2_29, u1_L2_3, u1_L2_30, 
        u1_L2_4, u1_L2_5, u1_L2_6, u1_L2_8, u1_L4_13, u1_L4_18, u1_L4_2, u1_L4_28, u1_L6_11, 
        u1_L6_19, u1_L6_29, u1_L6_4, u1_R0_22, u1_R0_23, u1_R11_10, u1_R11_11, u1_R11_22, u1_R11_23, 
        u1_R11_6, u1_R11_7, u1_R11_8, u1_R12_10, u1_R12_11, u1_R12_2, u1_R12_3, u1_R13_6, u1_R13_7, 
        u1_R1_18, u1_R1_19, u1_R1_2, u1_R1_3, u1_R2_10, u1_R2_11, u1_R2_18, u1_R2_19, u1_R2_20, 
        u1_R2_21, u1_R2_22, u1_R2_23, u1_R2_30, u1_R2_31, u1_R4_6, u1_R4_7, u1_R6_22, u1_R6_23, 
        u1_u12_X_12, u1_u12_X_14, u1_u12_X_17, u1_u12_X_18, u1_u12_X_31, u1_u12_X_32, u1_u12_X_35, u1_u12_X_36, u1_u12_X_7, 
        u1_u12_X_8, u1_u13_X_1, u1_u13_X_13, u1_u13_X_14, u1_u13_X_17, u1_u13_X_18, u1_u13_X_2, u1_u13_X_5, u1_u13_X_6, 
        u1_u14_X_11, u1_u14_X_12, u1_u14_X_7, u1_u14_X_8, u1_u15_X_43, u1_u15_X_44, u1_u15_X_47, u1_u15_X_48, u1_u1_X_31, 
        u1_u1_X_32, u1_u1_X_35, u1_u1_X_36, u1_u2_X_1, u1_u2_X_2, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, 
        u1_u2_X_5, u1_u2_X_6, u1_u3_X_13, u1_u3_X_14, u1_u3_X_17, u1_u3_X_18, u1_u3_X_25, u1_u3_X_26, u1_u3_X_35, 
        u1_u3_X_36, u1_u3_X_43, u1_u3_X_44, u1_u3_X_47, u1_u3_X_48, u1_u5_X_11, u1_u5_X_12, u1_u5_X_7, u1_u5_X_8, 
        u1_u7_X_31, u1_u7_X_32, u1_u7_X_35, u1_u7_X_36, u1_uk_n1060, u1_uk_n1063, u1_uk_n1088, u1_uk_n1104, u1_uk_n1137, 
        u1_uk_n671, u1_uk_n672, u1_uk_n677, u1_uk_n678, u2_K6_13, u2_K6_14, u2_K6_15, u2_K6_16, u2_K8_5, 
        u2_L4_16, u2_L4_24, u2_L4_30, u2_L4_6, u2_L6_17, u2_L6_23, u2_L6_31, u2_L6_9, u2_R4_10, 
        u2_R4_11, u2_R4_12, u2_R4_13, u2_R4_8, u2_R4_9, u2_R6_1, u2_R6_2, u2_R6_3, u2_R6_32, 
        u2_R6_4, u2_R6_5, u2_uk_K_r4_11, u2_uk_K_r4_17, u2_uk_K_r4_4, u2_uk_K_r4_55, u2_uk_K_r6_10, u2_uk_K_r6_3, u2_uk_n100, 
        u2_uk_n102, u2_uk_n1105, u2_uk_n1116, u2_uk_n117, u2_uk_n118, u2_uk_n147, u2_uk_n1502, u2_uk_n1507, u2_uk_n1514, 
        u2_uk_n1515, u2_uk_n1518, u2_uk_n1519, u2_uk_n155, u2_uk_n162, u2_uk_n182, u2_uk_n188, u2_uk_n27, u2_uk_n83;
  output u0_FP_1, u0_FP_10, u0_FP_14, u0_FP_16, u0_FP_20, u0_FP_24, u0_FP_25, u0_FP_26, u0_FP_3, 
        u0_FP_30, u0_FP_6, u0_FP_8, u0_N106, u0_N114, u0_N124, u0_N195, u0_N196, u0_N198, 
        u0_N200, u0_N202, u0_N203, u0_N206, u0_N208, u0_N210, u0_N212, u0_N213, u0_N214, 
        u0_N218, u0_N220, u0_N222, u0_N223, u0_N296, u0_N304, u0_N310, u0_N318, u0_N321, 
        u0_N323, u0_N326, u0_N328, u0_N33, u0_N330, u0_N331, u0_N332, u0_N336, u0_N337, 
        u0_N338, u0_N341, u0_N342, u0_N347, u0_N348, u0_N350, u0_N351, u0_N353, u0_N357, 
        u0_N358, u0_N363, u0_N364, u0_N367, u0_N369, u0_N37, u0_N373, u0_N375, u0_N379, 
        u0_N38, u0_N381, u0_N383, u0_N40, u0_N43, u0_N44, u0_N47, u0_N48, u0_N49, 
        u0_N53, u0_N54, u0_N55, u0_N59, u0_N61, u0_N62, u0_N63, u0_N64, u0_N65, 
        u0_N67, u0_N69, u0_N72, u0_N73, u0_N74, u0_N76, u0_N79, u0_N80, u0_N81, 
        u0_N82, u0_N83, u0_N86, u0_N87, u0_N89, u0_N91, u0_N92, u0_N93, u0_N94, 
        u0_N99, u0_uk_n100, u0_uk_n109, u0_uk_n110, u0_uk_n129, u0_uk_n142, u0_uk_n146, u0_uk_n147, u0_uk_n148, 
        u0_uk_n155, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n191, u0_uk_n203, u0_uk_n208, u0_uk_n214, u0_uk_n217, 
        u0_uk_n220, u0_uk_n222, u0_uk_n230, u0_uk_n231, u0_uk_n240, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n778, 
        u0_uk_n823, u0_uk_n83, u0_uk_n841, u0_uk_n863, u0_uk_n867, u0_uk_n93, u0_uk_n94, u1_FP_15, u1_FP_21, 
        u1_FP_27, u1_FP_5, u1_N100, u1_N101, u1_N103, u1_N106, u1_N109, u1_N110, u1_N111, 
        u1_N114, u1_N116, u1_N119, u1_N120, u1_N122, u1_N124, u1_N125, u1_N161, u1_N172, 
        u1_N177, u1_N187, u1_N227, u1_N234, u1_N242, u1_N252, u1_N35, u1_N385, u1_N387, 
        u1_N389, u1_N394, u1_N396, u1_N399, u1_N401, u1_N402, u1_N407, u1_N411, u1_N412, 
        u1_N413, u1_N42, u1_N421, u1_N424, u1_N431, u1_N432, u1_N438, u1_N439, u1_N445, 
        u1_N446, u1_N449, u1_N460, u1_N465, u1_N475, u1_N50, u1_N60, u1_N66, u1_N71, 
        u1_N72, u1_N77, u1_N80, u1_N86, u1_N88, u1_N94, u1_N98, u1_N99, u2_N165, 
        u2_N175, u2_N183, u2_N189, u2_N232, u2_N240, u2_N246, u2_N254;
  wire u0_K10_1, u0_K10_2, u0_K10_3, u0_K10_4, u0_K10_5, u0_K10_6, u0_K11_1, u0_K11_10, u0_K11_11, 
       u0_K11_12, u0_K11_2, u0_K11_3, u0_K11_31, u0_K11_32, u0_K11_33, u0_K11_34, u0_K11_35, u0_K11_36, 
       u0_K11_38, u0_K11_39, u0_K11_4, u0_K11_40, u0_K11_41, u0_K11_42, u0_K11_5, u0_K11_6, u0_K11_7, 
       u0_K11_8, u0_K11_9, u0_K12_10, u0_K12_11, u0_K12_12, u0_K12_13, u0_K12_14, u0_K12_15, u0_K12_16, 
       u0_K12_17, u0_K12_18, u0_K12_37, u0_K12_38, u0_K12_41, u0_K12_42, u0_K12_8, u0_K16_13, u0_K16_14, 
       u0_K16_15, u0_K16_16, u0_K16_17, u0_K16_20, u0_K16_21, u0_K16_23, u0_K16_25, u0_K16_27, u0_K16_28, 
       u0_K16_29, u0_K16_30, u0_K2_1, u0_K2_10, u0_K2_13, u0_K2_14, u0_K2_15, u0_K2_16, u0_K2_17, 
       u0_K2_18, u0_K2_2, u0_K2_3, u0_K2_37, u0_K2_38, u0_K2_39, u0_K2_40, u0_K2_41, u0_K2_42, 
       u0_K2_7, u0_K2_9, u0_K3_1, u0_K3_11, u0_K3_13, u0_K3_16, u0_K3_2, u0_K3_20, u0_K3_21, 
       u0_K3_22, u0_K3_24, u0_K3_3, u0_K3_31, u0_K3_32, u0_K3_33, u0_K3_35, u0_K3_36, u0_K3_4, 
       u0_K3_6, u0_K3_7, u0_K3_8, u0_K3_9, u0_K4_31, u0_K4_32, u0_K4_33, u0_K4_34, u0_K4_36, 
       u0_K7_1, u0_K7_3, u0_K7_31, u0_K7_32, u0_K7_33, u0_K7_34, u0_K7_35, u0_K7_36, u0_K7_37, 
       u0_K7_38, u0_K7_39, u0_K7_4, u0_K7_40, u0_K7_41, u0_K7_42, u0_K7_43, u0_K7_44, u0_K7_45, 
       u0_K7_46, u0_K7_47, u0_K7_48, u0_K7_5, u0_out10_11, u0_out10_12, u0_out10_13, u0_out10_17, u0_out10_18, 
       u0_out10_19, u0_out10_2, u0_out10_22, u0_out10_23, u0_out10_28, u0_out10_29, u0_out10_31, u0_out10_32, u0_out10_4, 
       u0_out10_7, u0_out10_9, u0_out11_12, u0_out11_13, u0_out11_16, u0_out11_18, u0_out11_2, u0_out11_22, u0_out11_24, 
       u0_out11_28, u0_out11_30, u0_out11_32, u0_out11_6, u0_out11_7, u0_out15_1, u0_out15_10, u0_out15_14, u0_out15_16, 
       u0_out15_20, u0_out15_24, u0_out15_25, u0_out15_26, u0_out15_3, u0_out15_30, u0_out15_6, u0_out15_8, u0_out1_12, 
       u0_out1_13, u0_out1_16, u0_out1_17, u0_out1_18, u0_out1_2, u0_out1_22, u0_out1_23, u0_out1_24, u0_out1_28, 
       u0_out1_30, u0_out1_31, u0_out1_32, u0_out1_6, u0_out1_7, u0_out1_9, u0_out2_1, u0_out2_10, u0_out2_11, 
       u0_out2_13, u0_out2_16, u0_out2_17, u0_out2_18, u0_out2_19, u0_out2_2, u0_out2_20, u0_out2_23, u0_out2_24, 
       u0_out2_26, u0_out2_28, u0_out2_29, u0_out2_30, u0_out2_31, u0_out2_4, u0_out2_6, u0_out2_9, u0_out3_11, 
       u0_out3_19, u0_out3_29, u0_out3_4, u0_out6_11, u0_out6_12, u0_out6_15, u0_out6_17, u0_out6_19, u0_out6_21, 
       u0_out6_22, u0_out6_23, u0_out6_27, u0_out6_29, u0_out6_31, u0_out6_32, u0_out6_4, u0_out6_5, u0_out6_7, 
       u0_out6_9, u0_out9_17, u0_out9_23, u0_out9_31, u0_out9_9, u0_u10_X_1, u0_u10_X_10, u0_u10_X_11, u0_u10_X_12, 
       u0_u10_X_2, u0_u10_X_3, u0_u10_X_31, u0_u10_X_32, u0_u10_X_33, u0_u10_X_34, u0_u10_X_35, u0_u10_X_36, u0_u10_X_37, 
       u0_u10_X_38, u0_u10_X_39, u0_u10_X_4, u0_u10_X_40, u0_u10_X_41, u0_u10_X_42, u0_u10_X_5, u0_u10_X_6, u0_u10_X_7, 
       u0_u10_X_8, u0_u10_X_9, u0_u10_u0_n100, u0_u10_u0_n101, u0_u10_u0_n102, u0_u10_u0_n103, u0_u10_u0_n104, u0_u10_u0_n105, u0_u10_u0_n106, 
       u0_u10_u0_n107, u0_u10_u0_n108, u0_u10_u0_n109, u0_u10_u0_n110, u0_u10_u0_n111, u0_u10_u0_n112, u0_u10_u0_n113, u0_u10_u0_n114, u0_u10_u0_n115, 
       u0_u10_u0_n116, u0_u10_u0_n117, u0_u10_u0_n118, u0_u10_u0_n119, u0_u10_u0_n120, u0_u10_u0_n121, u0_u10_u0_n122, u0_u10_u0_n123, u0_u10_u0_n124, 
       u0_u10_u0_n125, u0_u10_u0_n126, u0_u10_u0_n127, u0_u10_u0_n128, u0_u10_u0_n129, u0_u10_u0_n130, u0_u10_u0_n131, u0_u10_u0_n132, u0_u10_u0_n133, 
       u0_u10_u0_n134, u0_u10_u0_n135, u0_u10_u0_n136, u0_u10_u0_n137, u0_u10_u0_n138, u0_u10_u0_n139, u0_u10_u0_n140, u0_u10_u0_n141, u0_u10_u0_n142, 
       u0_u10_u0_n143, u0_u10_u0_n144, u0_u10_u0_n145, u0_u10_u0_n146, u0_u10_u0_n147, u0_u10_u0_n148, u0_u10_u0_n149, u0_u10_u0_n150, u0_u10_u0_n151, 
       u0_u10_u0_n152, u0_u10_u0_n153, u0_u10_u0_n154, u0_u10_u0_n155, u0_u10_u0_n156, u0_u10_u0_n157, u0_u10_u0_n158, u0_u10_u0_n159, u0_u10_u0_n160, 
       u0_u10_u0_n161, u0_u10_u0_n162, u0_u10_u0_n163, u0_u10_u0_n164, u0_u10_u0_n165, u0_u10_u0_n166, u0_u10_u0_n167, u0_u10_u0_n168, u0_u10_u0_n169, 
       u0_u10_u0_n170, u0_u10_u0_n171, u0_u10_u0_n172, u0_u10_u0_n173, u0_u10_u0_n174, u0_u10_u0_n88, u0_u10_u0_n89, u0_u10_u0_n90, u0_u10_u0_n91, 
       u0_u10_u0_n92, u0_u10_u0_n93, u0_u10_u0_n94, u0_u10_u0_n95, u0_u10_u0_n96, u0_u10_u0_n97, u0_u10_u0_n98, u0_u10_u0_n99, u0_u10_u1_n100, 
       u0_u10_u1_n101, u0_u10_u1_n102, u0_u10_u1_n103, u0_u10_u1_n104, u0_u10_u1_n105, u0_u10_u1_n106, u0_u10_u1_n107, u0_u10_u1_n108, u0_u10_u1_n109, 
       u0_u10_u1_n110, u0_u10_u1_n111, u0_u10_u1_n112, u0_u10_u1_n113, u0_u10_u1_n114, u0_u10_u1_n115, u0_u10_u1_n116, u0_u10_u1_n117, u0_u10_u1_n118, 
       u0_u10_u1_n119, u0_u10_u1_n120, u0_u10_u1_n121, u0_u10_u1_n122, u0_u10_u1_n123, u0_u10_u1_n124, u0_u10_u1_n125, u0_u10_u1_n126, u0_u10_u1_n127, 
       u0_u10_u1_n128, u0_u10_u1_n129, u0_u10_u1_n130, u0_u10_u1_n131, u0_u10_u1_n132, u0_u10_u1_n133, u0_u10_u1_n134, u0_u10_u1_n135, u0_u10_u1_n136, 
       u0_u10_u1_n137, u0_u10_u1_n138, u0_u10_u1_n139, u0_u10_u1_n140, u0_u10_u1_n141, u0_u10_u1_n142, u0_u10_u1_n143, u0_u10_u1_n144, u0_u10_u1_n145, 
       u0_u10_u1_n146, u0_u10_u1_n147, u0_u10_u1_n148, u0_u10_u1_n149, u0_u10_u1_n150, u0_u10_u1_n151, u0_u10_u1_n152, u0_u10_u1_n153, u0_u10_u1_n154, 
       u0_u10_u1_n155, u0_u10_u1_n156, u0_u10_u1_n157, u0_u10_u1_n158, u0_u10_u1_n159, u0_u10_u1_n160, u0_u10_u1_n161, u0_u10_u1_n162, u0_u10_u1_n163, 
       u0_u10_u1_n164, u0_u10_u1_n165, u0_u10_u1_n166, u0_u10_u1_n167, u0_u10_u1_n168, u0_u10_u1_n169, u0_u10_u1_n170, u0_u10_u1_n171, u0_u10_u1_n172, 
       u0_u10_u1_n173, u0_u10_u1_n174, u0_u10_u1_n175, u0_u10_u1_n176, u0_u10_u1_n177, u0_u10_u1_n178, u0_u10_u1_n179, u0_u10_u1_n180, u0_u10_u1_n181, 
       u0_u10_u1_n182, u0_u10_u1_n183, u0_u10_u1_n184, u0_u10_u1_n185, u0_u10_u1_n186, u0_u10_u1_n187, u0_u10_u1_n188, u0_u10_u1_n95, u0_u10_u1_n96, 
       u0_u10_u1_n97, u0_u10_u1_n98, u0_u10_u1_n99, u0_u10_u5_n100, u0_u10_u5_n101, u0_u10_u5_n102, u0_u10_u5_n103, u0_u10_u5_n104, u0_u10_u5_n105, 
       u0_u10_u5_n106, u0_u10_u5_n107, u0_u10_u5_n108, u0_u10_u5_n109, u0_u10_u5_n110, u0_u10_u5_n111, u0_u10_u5_n112, u0_u10_u5_n113, u0_u10_u5_n114, 
       u0_u10_u5_n115, u0_u10_u5_n116, u0_u10_u5_n117, u0_u10_u5_n118, u0_u10_u5_n119, u0_u10_u5_n120, u0_u10_u5_n121, u0_u10_u5_n122, u0_u10_u5_n123, 
       u0_u10_u5_n124, u0_u10_u5_n125, u0_u10_u5_n126, u0_u10_u5_n127, u0_u10_u5_n128, u0_u10_u5_n129, u0_u10_u5_n130, u0_u10_u5_n131, u0_u10_u5_n132, 
       u0_u10_u5_n133, u0_u10_u5_n134, u0_u10_u5_n135, u0_u10_u5_n136, u0_u10_u5_n137, u0_u10_u5_n138, u0_u10_u5_n139, u0_u10_u5_n140, u0_u10_u5_n141, 
       u0_u10_u5_n142, u0_u10_u5_n143, u0_u10_u5_n144, u0_u10_u5_n145, u0_u10_u5_n146, u0_u10_u5_n147, u0_u10_u5_n148, u0_u10_u5_n149, u0_u10_u5_n150, 
       u0_u10_u5_n151, u0_u10_u5_n152, u0_u10_u5_n153, u0_u10_u5_n154, u0_u10_u5_n155, u0_u10_u5_n156, u0_u10_u5_n157, u0_u10_u5_n158, u0_u10_u5_n159, 
       u0_u10_u5_n160, u0_u10_u5_n161, u0_u10_u5_n162, u0_u10_u5_n163, u0_u10_u5_n164, u0_u10_u5_n165, u0_u10_u5_n166, u0_u10_u5_n167, u0_u10_u5_n168, 
       u0_u10_u5_n169, u0_u10_u5_n170, u0_u10_u5_n171, u0_u10_u5_n172, u0_u10_u5_n173, u0_u10_u5_n174, u0_u10_u5_n175, u0_u10_u5_n176, u0_u10_u5_n177, 
       u0_u10_u5_n178, u0_u10_u5_n179, u0_u10_u5_n180, u0_u10_u5_n181, u0_u10_u5_n182, u0_u10_u5_n183, u0_u10_u5_n184, u0_u10_u5_n185, u0_u10_u5_n186, 
       u0_u10_u5_n187, u0_u10_u5_n188, u0_u10_u5_n189, u0_u10_u5_n190, u0_u10_u5_n191, u0_u10_u5_n192, u0_u10_u5_n193, u0_u10_u5_n194, u0_u10_u5_n195, 
       u0_u10_u5_n196, u0_u10_u5_n99, u0_u10_u6_n100, u0_u10_u6_n101, u0_u10_u6_n102, u0_u10_u6_n103, u0_u10_u6_n104, u0_u10_u6_n105, u0_u10_u6_n106, 
       u0_u10_u6_n107, u0_u10_u6_n108, u0_u10_u6_n109, u0_u10_u6_n110, u0_u10_u6_n111, u0_u10_u6_n112, u0_u10_u6_n113, u0_u10_u6_n114, u0_u10_u6_n115, 
       u0_u10_u6_n116, u0_u10_u6_n117, u0_u10_u6_n118, u0_u10_u6_n119, u0_u10_u6_n120, u0_u10_u6_n121, u0_u10_u6_n122, u0_u10_u6_n123, u0_u10_u6_n124, 
       u0_u10_u6_n125, u0_u10_u6_n126, u0_u10_u6_n127, u0_u10_u6_n128, u0_u10_u6_n129, u0_u10_u6_n130, u0_u10_u6_n131, u0_u10_u6_n132, u0_u10_u6_n133, 
       u0_u10_u6_n134, u0_u10_u6_n135, u0_u10_u6_n136, u0_u10_u6_n137, u0_u10_u6_n138, u0_u10_u6_n139, u0_u10_u6_n140, u0_u10_u6_n141, u0_u10_u6_n142, 
       u0_u10_u6_n143, u0_u10_u6_n144, u0_u10_u6_n145, u0_u10_u6_n146, u0_u10_u6_n147, u0_u10_u6_n148, u0_u10_u6_n149, u0_u10_u6_n150, u0_u10_u6_n151, 
       u0_u10_u6_n152, u0_u10_u6_n153, u0_u10_u6_n154, u0_u10_u6_n155, u0_u10_u6_n156, u0_u10_u6_n157, u0_u10_u6_n158, u0_u10_u6_n159, u0_u10_u6_n160, 
       u0_u10_u6_n161, u0_u10_u6_n162, u0_u10_u6_n163, u0_u10_u6_n164, u0_u10_u6_n165, u0_u10_u6_n166, u0_u10_u6_n167, u0_u10_u6_n168, u0_u10_u6_n169, 
       u0_u10_u6_n170, u0_u10_u6_n171, u0_u10_u6_n172, u0_u10_u6_n173, u0_u10_u6_n174, u0_u10_u6_n88, u0_u10_u6_n89, u0_u10_u6_n90, u0_u10_u6_n91, 
       u0_u10_u6_n92, u0_u10_u6_n93, u0_u10_u6_n94, u0_u10_u6_n95, u0_u10_u6_n96, u0_u10_u6_n97, u0_u10_u6_n98, u0_u10_u6_n99, u0_u11_X_10, 
       u0_u11_X_11, u0_u11_X_12, u0_u11_X_13, u0_u11_X_14, u0_u11_X_15, u0_u11_X_16, u0_u11_X_17, u0_u11_X_18, u0_u11_X_37, 
       u0_u11_X_38, u0_u11_X_39, u0_u11_X_40, u0_u11_X_41, u0_u11_X_42, u0_u11_X_7, u0_u11_X_8, u0_u11_X_9, u0_u11_u1_n100, 
       u0_u11_u1_n101, u0_u11_u1_n102, u0_u11_u1_n103, u0_u11_u1_n104, u0_u11_u1_n105, u0_u11_u1_n106, u0_u11_u1_n107, u0_u11_u1_n108, u0_u11_u1_n109, 
       u0_u11_u1_n110, u0_u11_u1_n111, u0_u11_u1_n112, u0_u11_u1_n113, u0_u11_u1_n114, u0_u11_u1_n115, u0_u11_u1_n116, u0_u11_u1_n117, u0_u11_u1_n118, 
       u0_u11_u1_n119, u0_u11_u1_n120, u0_u11_u1_n121, u0_u11_u1_n122, u0_u11_u1_n123, u0_u11_u1_n124, u0_u11_u1_n125, u0_u11_u1_n126, u0_u11_u1_n127, 
       u0_u11_u1_n128, u0_u11_u1_n129, u0_u11_u1_n130, u0_u11_u1_n131, u0_u11_u1_n132, u0_u11_u1_n133, u0_u11_u1_n134, u0_u11_u1_n135, u0_u11_u1_n136, 
       u0_u11_u1_n137, u0_u11_u1_n138, u0_u11_u1_n139, u0_u11_u1_n140, u0_u11_u1_n141, u0_u11_u1_n142, u0_u11_u1_n143, u0_u11_u1_n144, u0_u11_u1_n145, 
       u0_u11_u1_n146, u0_u11_u1_n147, u0_u11_u1_n148, u0_u11_u1_n149, u0_u11_u1_n150, u0_u11_u1_n151, u0_u11_u1_n152, u0_u11_u1_n153, u0_u11_u1_n154, 
       u0_u11_u1_n155, u0_u11_u1_n156, u0_u11_u1_n157, u0_u11_u1_n158, u0_u11_u1_n159, u0_u11_u1_n160, u0_u11_u1_n161, u0_u11_u1_n162, u0_u11_u1_n163, 
       u0_u11_u1_n164, u0_u11_u1_n165, u0_u11_u1_n166, u0_u11_u1_n167, u0_u11_u1_n168, u0_u11_u1_n169, u0_u11_u1_n170, u0_u11_u1_n171, u0_u11_u1_n172, 
       u0_u11_u1_n173, u0_u11_u1_n174, u0_u11_u1_n175, u0_u11_u1_n176, u0_u11_u1_n177, u0_u11_u1_n178, u0_u11_u1_n179, u0_u11_u1_n180, u0_u11_u1_n181, 
       u0_u11_u1_n182, u0_u11_u1_n183, u0_u11_u1_n184, u0_u11_u1_n185, u0_u11_u1_n186, u0_u11_u1_n187, u0_u11_u1_n188, u0_u11_u1_n95, u0_u11_u1_n96, 
       u0_u11_u1_n97, u0_u11_u1_n98, u0_u11_u1_n99, u0_u11_u2_n100, u0_u11_u2_n101, u0_u11_u2_n102, u0_u11_u2_n103, u0_u11_u2_n104, u0_u11_u2_n105, 
       u0_u11_u2_n106, u0_u11_u2_n107, u0_u11_u2_n108, u0_u11_u2_n109, u0_u11_u2_n110, u0_u11_u2_n111, u0_u11_u2_n112, u0_u11_u2_n113, u0_u11_u2_n114, 
       u0_u11_u2_n115, u0_u11_u2_n116, u0_u11_u2_n117, u0_u11_u2_n118, u0_u11_u2_n119, u0_u11_u2_n120, u0_u11_u2_n121, u0_u11_u2_n122, u0_u11_u2_n123, 
       u0_u11_u2_n124, u0_u11_u2_n125, u0_u11_u2_n126, u0_u11_u2_n127, u0_u11_u2_n128, u0_u11_u2_n129, u0_u11_u2_n130, u0_u11_u2_n131, u0_u11_u2_n132, 
       u0_u11_u2_n133, u0_u11_u2_n134, u0_u11_u2_n135, u0_u11_u2_n136, u0_u11_u2_n137, u0_u11_u2_n138, u0_u11_u2_n139, u0_u11_u2_n140, u0_u11_u2_n141, 
       u0_u11_u2_n142, u0_u11_u2_n143, u0_u11_u2_n144, u0_u11_u2_n145, u0_u11_u2_n146, u0_u11_u2_n147, u0_u11_u2_n148, u0_u11_u2_n149, u0_u11_u2_n150, 
       u0_u11_u2_n151, u0_u11_u2_n152, u0_u11_u2_n153, u0_u11_u2_n154, u0_u11_u2_n155, u0_u11_u2_n156, u0_u11_u2_n157, u0_u11_u2_n158, u0_u11_u2_n159, 
       u0_u11_u2_n160, u0_u11_u2_n161, u0_u11_u2_n162, u0_u11_u2_n163, u0_u11_u2_n164, u0_u11_u2_n165, u0_u11_u2_n166, u0_u11_u2_n167, u0_u11_u2_n168, 
       u0_u11_u2_n169, u0_u11_u2_n170, u0_u11_u2_n171, u0_u11_u2_n172, u0_u11_u2_n173, u0_u11_u2_n174, u0_u11_u2_n175, u0_u11_u2_n176, u0_u11_u2_n177, 
       u0_u11_u2_n178, u0_u11_u2_n179, u0_u11_u2_n180, u0_u11_u2_n181, u0_u11_u2_n182, u0_u11_u2_n183, u0_u11_u2_n184, u0_u11_u2_n185, u0_u11_u2_n186, 
       u0_u11_u2_n187, u0_u11_u2_n188, u0_u11_u2_n95, u0_u11_u2_n96, u0_u11_u2_n97, u0_u11_u2_n98, u0_u11_u2_n99, u0_u11_u6_n100, u0_u11_u6_n101, 
       u0_u11_u6_n102, u0_u11_u6_n103, u0_u11_u6_n104, u0_u11_u6_n105, u0_u11_u6_n106, u0_u11_u6_n107, u0_u11_u6_n108, u0_u11_u6_n109, u0_u11_u6_n110, 
       u0_u11_u6_n111, u0_u11_u6_n112, u0_u11_u6_n113, u0_u11_u6_n114, u0_u11_u6_n115, u0_u11_u6_n116, u0_u11_u6_n117, u0_u11_u6_n118, u0_u11_u6_n119, 
       u0_u11_u6_n120, u0_u11_u6_n121, u0_u11_u6_n122, u0_u11_u6_n123, u0_u11_u6_n124, u0_u11_u6_n125, u0_u11_u6_n126, u0_u11_u6_n127, u0_u11_u6_n128, 
       u0_u11_u6_n129, u0_u11_u6_n130, u0_u11_u6_n131, u0_u11_u6_n132, u0_u11_u6_n133, u0_u11_u6_n134, u0_u11_u6_n135, u0_u11_u6_n136, u0_u11_u6_n137, 
       u0_u11_u6_n138, u0_u11_u6_n139, u0_u11_u6_n140, u0_u11_u6_n141, u0_u11_u6_n142, u0_u11_u6_n143, u0_u11_u6_n144, u0_u11_u6_n145, u0_u11_u6_n146, 
       u0_u11_u6_n147, u0_u11_u6_n148, u0_u11_u6_n149, u0_u11_u6_n150, u0_u11_u6_n151, u0_u11_u6_n152, u0_u11_u6_n153, u0_u11_u6_n154, u0_u11_u6_n155, 
       u0_u11_u6_n156, u0_u11_u6_n157, u0_u11_u6_n158, u0_u11_u6_n159, u0_u11_u6_n160, u0_u11_u6_n161, u0_u11_u6_n162, u0_u11_u6_n163, u0_u11_u6_n164, 
       u0_u11_u6_n165, u0_u11_u6_n166, u0_u11_u6_n167, u0_u11_u6_n168, u0_u11_u6_n169, u0_u11_u6_n170, u0_u11_u6_n171, u0_u11_u6_n172, u0_u11_u6_n173, 
       u0_u11_u6_n174, u0_u11_u6_n88, u0_u11_u6_n89, u0_u11_u6_n90, u0_u11_u6_n91, u0_u11_u6_n92, u0_u11_u6_n93, u0_u11_u6_n94, u0_u11_u6_n95, 
       u0_u11_u6_n96, u0_u11_u6_n97, u0_u11_u6_n98, u0_u11_u6_n99, u0_u15_X_13, u0_u15_X_14, u0_u15_X_15, u0_u15_X_16, u0_u15_X_17, 
       u0_u15_X_18, u0_u15_X_19, u0_u15_X_20, u0_u15_X_21, u0_u15_X_22, u0_u15_X_23, u0_u15_X_24, u0_u15_X_25, u0_u15_X_26, 
       u0_u15_X_27, u0_u15_X_28, u0_u15_X_29, u0_u15_X_30, u0_u15_u2_n100, u0_u15_u2_n101, u0_u15_u2_n102, u0_u15_u2_n103, u0_u15_u2_n104, 
       u0_u15_u2_n105, u0_u15_u2_n106, u0_u15_u2_n107, u0_u15_u2_n108, u0_u15_u2_n109, u0_u15_u2_n110, u0_u15_u2_n111, u0_u15_u2_n112, u0_u15_u2_n113, 
       u0_u15_u2_n114, u0_u15_u2_n115, u0_u15_u2_n116, u0_u15_u2_n117, u0_u15_u2_n118, u0_u15_u2_n119, u0_u15_u2_n120, u0_u15_u2_n121, u0_u15_u2_n122, 
       u0_u15_u2_n123, u0_u15_u2_n124, u0_u15_u2_n125, u0_u15_u2_n126, u0_u15_u2_n127, u0_u15_u2_n128, u0_u15_u2_n129, u0_u15_u2_n130, u0_u15_u2_n131, 
       u0_u15_u2_n132, u0_u15_u2_n133, u0_u15_u2_n134, u0_u15_u2_n135, u0_u15_u2_n136, u0_u15_u2_n137, u0_u15_u2_n138, u0_u15_u2_n139, u0_u15_u2_n140, 
       u0_u15_u2_n141, u0_u15_u2_n142, u0_u15_u2_n143, u0_u15_u2_n144, u0_u15_u2_n145, u0_u15_u2_n146, u0_u15_u2_n147, u0_u15_u2_n148, u0_u15_u2_n149, 
       u0_u15_u2_n150, u0_u15_u2_n151, u0_u15_u2_n152, u0_u15_u2_n153, u0_u15_u2_n154, u0_u15_u2_n155, u0_u15_u2_n156, u0_u15_u2_n157, u0_u15_u2_n158, 
       u0_u15_u2_n159, u0_u15_u2_n160, u0_u15_u2_n161, u0_u15_u2_n162, u0_u15_u2_n163, u0_u15_u2_n164, u0_u15_u2_n165, u0_u15_u2_n166, u0_u15_u2_n167, 
       u0_u15_u2_n168, u0_u15_u2_n169, u0_u15_u2_n170, u0_u15_u2_n171, u0_u15_u2_n172, u0_u15_u2_n173, u0_u15_u2_n174, u0_u15_u2_n175, u0_u15_u2_n176, 
       u0_u15_u2_n177, u0_u15_u2_n178, u0_u15_u2_n179, u0_u15_u2_n180, u0_u15_u2_n181, u0_u15_u2_n182, u0_u15_u2_n183, u0_u15_u2_n184, u0_u15_u2_n185, 
       u0_u15_u2_n186, u0_u15_u2_n187, u0_u15_u2_n188, u0_u15_u2_n95, u0_u15_u2_n96, u0_u15_u2_n97, u0_u15_u2_n98, u0_u15_u2_n99, u0_u15_u3_n100, 
       u0_u15_u3_n101, u0_u15_u3_n102, u0_u15_u3_n103, u0_u15_u3_n104, u0_u15_u3_n105, u0_u15_u3_n106, u0_u15_u3_n107, u0_u15_u3_n108, u0_u15_u3_n109, 
       u0_u15_u3_n110, u0_u15_u3_n111, u0_u15_u3_n112, u0_u15_u3_n113, u0_u15_u3_n114, u0_u15_u3_n115, u0_u15_u3_n116, u0_u15_u3_n117, u0_u15_u3_n118, 
       u0_u15_u3_n119, u0_u15_u3_n120, u0_u15_u3_n121, u0_u15_u3_n122, u0_u15_u3_n123, u0_u15_u3_n124, u0_u15_u3_n125, u0_u15_u3_n126, u0_u15_u3_n127, 
       u0_u15_u3_n128, u0_u15_u3_n129, u0_u15_u3_n130, u0_u15_u3_n131, u0_u15_u3_n132, u0_u15_u3_n133, u0_u15_u3_n134, u0_u15_u3_n135, u0_u15_u3_n136, 
       u0_u15_u3_n137, u0_u15_u3_n138, u0_u15_u3_n139, u0_u15_u3_n140, u0_u15_u3_n141, u0_u15_u3_n142, u0_u15_u3_n143, u0_u15_u3_n144, u0_u15_u3_n145, 
       u0_u15_u3_n146, u0_u15_u3_n147, u0_u15_u3_n148, u0_u15_u3_n149, u0_u15_u3_n150, u0_u15_u3_n151, u0_u15_u3_n152, u0_u15_u3_n153, u0_u15_u3_n154, 
       u0_u15_u3_n155, u0_u15_u3_n156, u0_u15_u3_n157, u0_u15_u3_n158, u0_u15_u3_n159, u0_u15_u3_n160, u0_u15_u3_n161, u0_u15_u3_n162, u0_u15_u3_n163, 
       u0_u15_u3_n164, u0_u15_u3_n165, u0_u15_u3_n166, u0_u15_u3_n167, u0_u15_u3_n168, u0_u15_u3_n169, u0_u15_u3_n170, u0_u15_u3_n171, u0_u15_u3_n172, 
       u0_u15_u3_n173, u0_u15_u3_n174, u0_u15_u3_n175, u0_u15_u3_n176, u0_u15_u3_n177, u0_u15_u3_n178, u0_u15_u3_n179, u0_u15_u3_n180, u0_u15_u3_n181, 
       u0_u15_u3_n182, u0_u15_u3_n183, u0_u15_u3_n184, u0_u15_u3_n185, u0_u15_u3_n186, u0_u15_u3_n94, u0_u15_u3_n95, u0_u15_u3_n96, u0_u15_u3_n97, 
       u0_u15_u3_n98, u0_u15_u3_n99, u0_u15_u4_n100, u0_u15_u4_n101, u0_u15_u4_n102, u0_u15_u4_n103, u0_u15_u4_n104, u0_u15_u4_n105, u0_u15_u4_n106, 
       u0_u15_u4_n107, u0_u15_u4_n108, u0_u15_u4_n109, u0_u15_u4_n110, u0_u15_u4_n111, u0_u15_u4_n112, u0_u15_u4_n113, u0_u15_u4_n114, u0_u15_u4_n115, 
       u0_u15_u4_n116, u0_u15_u4_n117, u0_u15_u4_n118, u0_u15_u4_n119, u0_u15_u4_n120, u0_u15_u4_n121, u0_u15_u4_n122, u0_u15_u4_n123, u0_u15_u4_n124, 
       u0_u15_u4_n125, u0_u15_u4_n126, u0_u15_u4_n127, u0_u15_u4_n128, u0_u15_u4_n129, u0_u15_u4_n130, u0_u15_u4_n131, u0_u15_u4_n132, u0_u15_u4_n133, 
       u0_u15_u4_n134, u0_u15_u4_n135, u0_u15_u4_n136, u0_u15_u4_n137, u0_u15_u4_n138, u0_u15_u4_n139, u0_u15_u4_n140, u0_u15_u4_n141, u0_u15_u4_n142, 
       u0_u15_u4_n143, u0_u15_u4_n144, u0_u15_u4_n145, u0_u15_u4_n146, u0_u15_u4_n147, u0_u15_u4_n148, u0_u15_u4_n149, u0_u15_u4_n150, u0_u15_u4_n151, 
       u0_u15_u4_n152, u0_u15_u4_n153, u0_u15_u4_n154, u0_u15_u4_n155, u0_u15_u4_n156, u0_u15_u4_n157, u0_u15_u4_n158, u0_u15_u4_n159, u0_u15_u4_n160, 
       u0_u15_u4_n161, u0_u15_u4_n162, u0_u15_u4_n163, u0_u15_u4_n164, u0_u15_u4_n165, u0_u15_u4_n166, u0_u15_u4_n167, u0_u15_u4_n168, u0_u15_u4_n169, 
       u0_u15_u4_n170, u0_u15_u4_n171, u0_u15_u4_n172, u0_u15_u4_n173, u0_u15_u4_n174, u0_u15_u4_n175, u0_u15_u4_n176, u0_u15_u4_n177, u0_u15_u4_n178, 
       u0_u15_u4_n179, u0_u15_u4_n180, u0_u15_u4_n181, u0_u15_u4_n182, u0_u15_u4_n183, u0_u15_u4_n184, u0_u15_u4_n185, u0_u15_u4_n186, u0_u15_u4_n94, 
       u0_u15_u4_n95, u0_u15_u4_n96, u0_u15_u4_n97, u0_u15_u4_n98, u0_u15_u4_n99, u0_u1_X_1, u0_u1_X_10, u0_u1_X_11, u0_u1_X_12, 
       u0_u1_X_13, u0_u1_X_14, u0_u1_X_15, u0_u1_X_16, u0_u1_X_17, u0_u1_X_18, u0_u1_X_2, u0_u1_X_3, u0_u1_X_37, 
       u0_u1_X_38, u0_u1_X_39, u0_u1_X_4, u0_u1_X_40, u0_u1_X_41, u0_u1_X_42, u0_u1_X_5, u0_u1_X_6, u0_u1_X_7, 
       u0_u1_X_8, u0_u1_X_9, u0_u1_u0_n100, u0_u1_u0_n101, u0_u1_u0_n102, u0_u1_u0_n103, u0_u1_u0_n104, u0_u1_u0_n105, u0_u1_u0_n106, 
       u0_u1_u0_n107, u0_u1_u0_n108, u0_u1_u0_n109, u0_u1_u0_n110, u0_u1_u0_n111, u0_u1_u0_n112, u0_u1_u0_n113, u0_u1_u0_n114, u0_u1_u0_n115, 
       u0_u1_u0_n116, u0_u1_u0_n117, u0_u1_u0_n118, u0_u1_u0_n119, u0_u1_u0_n120, u0_u1_u0_n121, u0_u1_u0_n122, u0_u1_u0_n123, u0_u1_u0_n124, 
       u0_u1_u0_n125, u0_u1_u0_n126, u0_u1_u0_n127, u0_u1_u0_n128, u0_u1_u0_n129, u0_u1_u0_n130, u0_u1_u0_n131, u0_u1_u0_n132, u0_u1_u0_n133, 
       u0_u1_u0_n134, u0_u1_u0_n135, u0_u1_u0_n136, u0_u1_u0_n137, u0_u1_u0_n138, u0_u1_u0_n139, u0_u1_u0_n140, u0_u1_u0_n141, u0_u1_u0_n142, 
       u0_u1_u0_n143, u0_u1_u0_n144, u0_u1_u0_n145, u0_u1_u0_n146, u0_u1_u0_n147, u0_u1_u0_n148, u0_u1_u0_n149, u0_u1_u0_n150, u0_u1_u0_n151, 
       u0_u1_u0_n152, u0_u1_u0_n153, u0_u1_u0_n154, u0_u1_u0_n155, u0_u1_u0_n156, u0_u1_u0_n157, u0_u1_u0_n158, u0_u1_u0_n159, u0_u1_u0_n160, 
       u0_u1_u0_n161, u0_u1_u0_n162, u0_u1_u0_n163, u0_u1_u0_n164, u0_u1_u0_n165, u0_u1_u0_n166, u0_u1_u0_n167, u0_u1_u0_n168, u0_u1_u0_n169, 
       u0_u1_u0_n170, u0_u1_u0_n171, u0_u1_u0_n172, u0_u1_u0_n173, u0_u1_u0_n174, u0_u1_u0_n88, u0_u1_u0_n89, u0_u1_u0_n90, u0_u1_u0_n91, 
       u0_u1_u0_n92, u0_u1_u0_n93, u0_u1_u0_n94, u0_u1_u0_n95, u0_u1_u0_n96, u0_u1_u0_n97, u0_u1_u0_n98, u0_u1_u0_n99, u0_u1_u1_n100, 
       u0_u1_u1_n101, u0_u1_u1_n102, u0_u1_u1_n103, u0_u1_u1_n104, u0_u1_u1_n105, u0_u1_u1_n106, u0_u1_u1_n107, u0_u1_u1_n108, u0_u1_u1_n109, 
       u0_u1_u1_n110, u0_u1_u1_n111, u0_u1_u1_n112, u0_u1_u1_n113, u0_u1_u1_n114, u0_u1_u1_n115, u0_u1_u1_n116, u0_u1_u1_n117, u0_u1_u1_n118, 
       u0_u1_u1_n119, u0_u1_u1_n120, u0_u1_u1_n121, u0_u1_u1_n122, u0_u1_u1_n123, u0_u1_u1_n124, u0_u1_u1_n125, u0_u1_u1_n126, u0_u1_u1_n127, 
       u0_u1_u1_n128, u0_u1_u1_n129, u0_u1_u1_n130, u0_u1_u1_n131, u0_u1_u1_n132, u0_u1_u1_n133, u0_u1_u1_n134, u0_u1_u1_n135, u0_u1_u1_n136, 
       u0_u1_u1_n137, u0_u1_u1_n138, u0_u1_u1_n139, u0_u1_u1_n140, u0_u1_u1_n141, u0_u1_u1_n142, u0_u1_u1_n143, u0_u1_u1_n144, u0_u1_u1_n145, 
       u0_u1_u1_n146, u0_u1_u1_n147, u0_u1_u1_n148, u0_u1_u1_n149, u0_u1_u1_n150, u0_u1_u1_n151, u0_u1_u1_n152, u0_u1_u1_n153, u0_u1_u1_n154, 
       u0_u1_u1_n155, u0_u1_u1_n156, u0_u1_u1_n157, u0_u1_u1_n158, u0_u1_u1_n159, u0_u1_u1_n160, u0_u1_u1_n161, u0_u1_u1_n162, u0_u1_u1_n163, 
       u0_u1_u1_n164, u0_u1_u1_n165, u0_u1_u1_n166, u0_u1_u1_n167, u0_u1_u1_n168, u0_u1_u1_n169, u0_u1_u1_n170, u0_u1_u1_n171, u0_u1_u1_n172, 
       u0_u1_u1_n173, u0_u1_u1_n174, u0_u1_u1_n175, u0_u1_u1_n176, u0_u1_u1_n177, u0_u1_u1_n178, u0_u1_u1_n179, u0_u1_u1_n180, u0_u1_u1_n181, 
       u0_u1_u1_n182, u0_u1_u1_n183, u0_u1_u1_n184, u0_u1_u1_n185, u0_u1_u1_n186, u0_u1_u1_n187, u0_u1_u1_n188, u0_u1_u1_n95, u0_u1_u1_n96, 
       u0_u1_u1_n97, u0_u1_u1_n98, u0_u1_u1_n99, u0_u1_u2_n100, u0_u1_u2_n101, u0_u1_u2_n102, u0_u1_u2_n103, u0_u1_u2_n104, u0_u1_u2_n105, 
       u0_u1_u2_n106, u0_u1_u2_n107, u0_u1_u2_n108, u0_u1_u2_n109, u0_u1_u2_n110, u0_u1_u2_n111, u0_u1_u2_n112, u0_u1_u2_n113, u0_u1_u2_n114, 
       u0_u1_u2_n115, u0_u1_u2_n116, u0_u1_u2_n117, u0_u1_u2_n118, u0_u1_u2_n119, u0_u1_u2_n120, u0_u1_u2_n121, u0_u1_u2_n122, u0_u1_u2_n123, 
       u0_u1_u2_n124, u0_u1_u2_n125, u0_u1_u2_n126, u0_u1_u2_n127, u0_u1_u2_n128, u0_u1_u2_n129, u0_u1_u2_n130, u0_u1_u2_n131, u0_u1_u2_n132, 
       u0_u1_u2_n133, u0_u1_u2_n134, u0_u1_u2_n135, u0_u1_u2_n136, u0_u1_u2_n137, u0_u1_u2_n138, u0_u1_u2_n139, u0_u1_u2_n140, u0_u1_u2_n141, 
       u0_u1_u2_n142, u0_u1_u2_n143, u0_u1_u2_n144, u0_u1_u2_n145, u0_u1_u2_n146, u0_u1_u2_n147, u0_u1_u2_n148, u0_u1_u2_n149, u0_u1_u2_n150, 
       u0_u1_u2_n151, u0_u1_u2_n152, u0_u1_u2_n153, u0_u1_u2_n154, u0_u1_u2_n155, u0_u1_u2_n156, u0_u1_u2_n157, u0_u1_u2_n158, u0_u1_u2_n159, 
       u0_u1_u2_n160, u0_u1_u2_n161, u0_u1_u2_n162, u0_u1_u2_n163, u0_u1_u2_n164, u0_u1_u2_n165, u0_u1_u2_n166, u0_u1_u2_n167, u0_u1_u2_n168, 
       u0_u1_u2_n169, u0_u1_u2_n170, u0_u1_u2_n171, u0_u1_u2_n172, u0_u1_u2_n173, u0_u1_u2_n174, u0_u1_u2_n175, u0_u1_u2_n176, u0_u1_u2_n177, 
       u0_u1_u2_n178, u0_u1_u2_n179, u0_u1_u2_n180, u0_u1_u2_n181, u0_u1_u2_n182, u0_u1_u2_n183, u0_u1_u2_n184, u0_u1_u2_n185, u0_u1_u2_n186, 
       u0_u1_u2_n187, u0_u1_u2_n188, u0_u1_u2_n95, u0_u1_u2_n96, u0_u1_u2_n97, u0_u1_u2_n98, u0_u1_u2_n99, u0_u1_u6_n100, u0_u1_u6_n101, 
       u0_u1_u6_n102, u0_u1_u6_n103, u0_u1_u6_n104, u0_u1_u6_n105, u0_u1_u6_n106, u0_u1_u6_n107, u0_u1_u6_n108, u0_u1_u6_n109, u0_u1_u6_n110, 
       u0_u1_u6_n111, u0_u1_u6_n112, u0_u1_u6_n113, u0_u1_u6_n114, u0_u1_u6_n115, u0_u1_u6_n116, u0_u1_u6_n117, u0_u1_u6_n118, u0_u1_u6_n119, 
       u0_u1_u6_n120, u0_u1_u6_n121, u0_u1_u6_n122, u0_u1_u6_n123, u0_u1_u6_n124, u0_u1_u6_n125, u0_u1_u6_n126, u0_u1_u6_n127, u0_u1_u6_n128, 
       u0_u1_u6_n129, u0_u1_u6_n130, u0_u1_u6_n131, u0_u1_u6_n132, u0_u1_u6_n133, u0_u1_u6_n134, u0_u1_u6_n135, u0_u1_u6_n136, u0_u1_u6_n137, 
       u0_u1_u6_n138, u0_u1_u6_n139, u0_u1_u6_n140, u0_u1_u6_n141, u0_u1_u6_n142, u0_u1_u6_n143, u0_u1_u6_n144, u0_u1_u6_n145, u0_u1_u6_n146, 
       u0_u1_u6_n147, u0_u1_u6_n148, u0_u1_u6_n149, u0_u1_u6_n150, u0_u1_u6_n151, u0_u1_u6_n152, u0_u1_u6_n153, u0_u1_u6_n154, u0_u1_u6_n155, 
       u0_u1_u6_n156, u0_u1_u6_n157, u0_u1_u6_n158, u0_u1_u6_n159, u0_u1_u6_n160, u0_u1_u6_n161, u0_u1_u6_n162, u0_u1_u6_n163, u0_u1_u6_n164, 
       u0_u1_u6_n165, u0_u1_u6_n166, u0_u1_u6_n167, u0_u1_u6_n168, u0_u1_u6_n169, u0_u1_u6_n170, u0_u1_u6_n171, u0_u1_u6_n172, u0_u1_u6_n173, 
       u0_u1_u6_n174, u0_u1_u6_n88, u0_u1_u6_n89, u0_u1_u6_n90, u0_u1_u6_n91, u0_u1_u6_n92, u0_u1_u6_n93, u0_u1_u6_n94, u0_u1_u6_n95, 
       u0_u1_u6_n96, u0_u1_u6_n97, u0_u1_u6_n98, u0_u1_u6_n99, u0_u2_X_1, u0_u2_X_10, u0_u2_X_11, u0_u2_X_12, u0_u2_X_13, 
       u0_u2_X_14, u0_u2_X_15, u0_u2_X_16, u0_u2_X_17, u0_u2_X_18, u0_u2_X_19, u0_u2_X_2, u0_u2_X_20, u0_u2_X_21, 
       u0_u2_X_22, u0_u2_X_23, u0_u2_X_24, u0_u2_X_3, u0_u2_X_31, u0_u2_X_32, u0_u2_X_33, u0_u2_X_34, u0_u2_X_35, 
       u0_u2_X_36, u0_u2_X_4, u0_u2_X_5, u0_u2_X_6, u0_u2_X_7, u0_u2_X_8, u0_u2_X_9, u0_u2_u0_n100, u0_u2_u0_n101, 
       u0_u2_u0_n102, u0_u2_u0_n103, u0_u2_u0_n104, u0_u2_u0_n105, u0_u2_u0_n106, u0_u2_u0_n107, u0_u2_u0_n108, u0_u2_u0_n109, u0_u2_u0_n110, 
       u0_u2_u0_n111, u0_u2_u0_n112, u0_u2_u0_n113, u0_u2_u0_n114, u0_u2_u0_n115, u0_u2_u0_n116, u0_u2_u0_n117, u0_u2_u0_n118, u0_u2_u0_n119, 
       u0_u2_u0_n120, u0_u2_u0_n121, u0_u2_u0_n122, u0_u2_u0_n123, u0_u2_u0_n124, u0_u2_u0_n125, u0_u2_u0_n126, u0_u2_u0_n127, u0_u2_u0_n128, 
       u0_u2_u0_n129, u0_u2_u0_n130, u0_u2_u0_n131, u0_u2_u0_n132, u0_u2_u0_n133, u0_u2_u0_n134, u0_u2_u0_n135, u0_u2_u0_n136, u0_u2_u0_n137, 
       u0_u2_u0_n138, u0_u2_u0_n139, u0_u2_u0_n140, u0_u2_u0_n141, u0_u2_u0_n142, u0_u2_u0_n143, u0_u2_u0_n144, u0_u2_u0_n145, u0_u2_u0_n146, 
       u0_u2_u0_n147, u0_u2_u0_n148, u0_u2_u0_n149, u0_u2_u0_n150, u0_u2_u0_n151, u0_u2_u0_n152, u0_u2_u0_n153, u0_u2_u0_n154, u0_u2_u0_n155, 
       u0_u2_u0_n156, u0_u2_u0_n157, u0_u2_u0_n158, u0_u2_u0_n159, u0_u2_u0_n160, u0_u2_u0_n161, u0_u2_u0_n162, u0_u2_u0_n163, u0_u2_u0_n164, 
       u0_u2_u0_n165, u0_u2_u0_n166, u0_u2_u0_n167, u0_u2_u0_n168, u0_u2_u0_n169, u0_u2_u0_n170, u0_u2_u0_n171, u0_u2_u0_n172, u0_u2_u0_n173, 
       u0_u2_u0_n174, u0_u2_u0_n88, u0_u2_u0_n89, u0_u2_u0_n90, u0_u2_u0_n91, u0_u2_u0_n92, u0_u2_u0_n93, u0_u2_u0_n94, u0_u2_u0_n95, 
       u0_u2_u0_n96, u0_u2_u0_n97, u0_u2_u0_n98, u0_u2_u0_n99, u0_u2_u1_n100, u0_u2_u1_n101, u0_u2_u1_n102, u0_u2_u1_n103, u0_u2_u1_n104, 
       u0_u2_u1_n105, u0_u2_u1_n106, u0_u2_u1_n107, u0_u2_u1_n108, u0_u2_u1_n109, u0_u2_u1_n110, u0_u2_u1_n111, u0_u2_u1_n112, u0_u2_u1_n113, 
       u0_u2_u1_n114, u0_u2_u1_n115, u0_u2_u1_n116, u0_u2_u1_n117, u0_u2_u1_n118, u0_u2_u1_n119, u0_u2_u1_n120, u0_u2_u1_n121, u0_u2_u1_n122, 
       u0_u2_u1_n123, u0_u2_u1_n124, u0_u2_u1_n125, u0_u2_u1_n126, u0_u2_u1_n127, u0_u2_u1_n128, u0_u2_u1_n129, u0_u2_u1_n130, u0_u2_u1_n131, 
       u0_u2_u1_n132, u0_u2_u1_n133, u0_u2_u1_n134, u0_u2_u1_n135, u0_u2_u1_n136, u0_u2_u1_n137, u0_u2_u1_n138, u0_u2_u1_n139, u0_u2_u1_n140, 
       u0_u2_u1_n141, u0_u2_u1_n142, u0_u2_u1_n143, u0_u2_u1_n144, u0_u2_u1_n145, u0_u2_u1_n146, u0_u2_u1_n147, u0_u2_u1_n148, u0_u2_u1_n149, 
       u0_u2_u1_n150, u0_u2_u1_n151, u0_u2_u1_n152, u0_u2_u1_n153, u0_u2_u1_n154, u0_u2_u1_n155, u0_u2_u1_n156, u0_u2_u1_n157, u0_u2_u1_n158, 
       u0_u2_u1_n159, u0_u2_u1_n160, u0_u2_u1_n161, u0_u2_u1_n162, u0_u2_u1_n163, u0_u2_u1_n164, u0_u2_u1_n165, u0_u2_u1_n166, u0_u2_u1_n167, 
       u0_u2_u1_n168, u0_u2_u1_n169, u0_u2_u1_n170, u0_u2_u1_n171, u0_u2_u1_n172, u0_u2_u1_n173, u0_u2_u1_n174, u0_u2_u1_n175, u0_u2_u1_n176, 
       u0_u2_u1_n177, u0_u2_u1_n178, u0_u2_u1_n179, u0_u2_u1_n180, u0_u2_u1_n181, u0_u2_u1_n182, u0_u2_u1_n183, u0_u2_u1_n184, u0_u2_u1_n185, 
       u0_u2_u1_n186, u0_u2_u1_n187, u0_u2_u1_n188, u0_u2_u1_n95, u0_u2_u1_n96, u0_u2_u1_n97, u0_u2_u1_n98, u0_u2_u1_n99, u0_u2_u2_n100, 
       u0_u2_u2_n101, u0_u2_u2_n102, u0_u2_u2_n103, u0_u2_u2_n104, u0_u2_u2_n105, u0_u2_u2_n106, u0_u2_u2_n107, u0_u2_u2_n108, u0_u2_u2_n109, 
       u0_u2_u2_n110, u0_u2_u2_n111, u0_u2_u2_n112, u0_u2_u2_n113, u0_u2_u2_n114, u0_u2_u2_n115, u0_u2_u2_n116, u0_u2_u2_n117, u0_u2_u2_n118, 
       u0_u2_u2_n119, u0_u2_u2_n120, u0_u2_u2_n121, u0_u2_u2_n122, u0_u2_u2_n123, u0_u2_u2_n124, u0_u2_u2_n125, u0_u2_u2_n126, u0_u2_u2_n127, 
       u0_u2_u2_n128, u0_u2_u2_n129, u0_u2_u2_n130, u0_u2_u2_n131, u0_u2_u2_n132, u0_u2_u2_n133, u0_u2_u2_n134, u0_u2_u2_n135, u0_u2_u2_n136, 
       u0_u2_u2_n137, u0_u2_u2_n138, u0_u2_u2_n139, u0_u2_u2_n140, u0_u2_u2_n141, u0_u2_u2_n142, u0_u2_u2_n143, u0_u2_u2_n144, u0_u2_u2_n145, 
       u0_u2_u2_n146, u0_u2_u2_n147, u0_u2_u2_n148, u0_u2_u2_n149, u0_u2_u2_n150, u0_u2_u2_n151, u0_u2_u2_n152, u0_u2_u2_n153, u0_u2_u2_n154, 
       u0_u2_u2_n155, u0_u2_u2_n156, u0_u2_u2_n157, u0_u2_u2_n158, u0_u2_u2_n159, u0_u2_u2_n160, u0_u2_u2_n161, u0_u2_u2_n162, u0_u2_u2_n163, 
       u0_u2_u2_n164, u0_u2_u2_n165, u0_u2_u2_n166, u0_u2_u2_n167, u0_u2_u2_n168, u0_u2_u2_n169, u0_u2_u2_n170, u0_u2_u2_n171, u0_u2_u2_n172, 
       u0_u2_u2_n173, u0_u2_u2_n174, u0_u2_u2_n175, u0_u2_u2_n176, u0_u2_u2_n177, u0_u2_u2_n178, u0_u2_u2_n179, u0_u2_u2_n180, u0_u2_u2_n181, 
       u0_u2_u2_n182, u0_u2_u2_n183, u0_u2_u2_n184, u0_u2_u2_n185, u0_u2_u2_n186, u0_u2_u2_n187, u0_u2_u2_n188, u0_u2_u2_n95, u0_u2_u2_n96, 
       u0_u2_u2_n97, u0_u2_u2_n98, u0_u2_u2_n99, u0_u2_u3_n100, u0_u2_u3_n101, u0_u2_u3_n102, u0_u2_u3_n103, u0_u2_u3_n104, u0_u2_u3_n105, 
       u0_u2_u3_n106, u0_u2_u3_n107, u0_u2_u3_n108, u0_u2_u3_n109, u0_u2_u3_n110, u0_u2_u3_n111, u0_u2_u3_n112, u0_u2_u3_n113, u0_u2_u3_n114, 
       u0_u2_u3_n115, u0_u2_u3_n116, u0_u2_u3_n117, u0_u2_u3_n118, u0_u2_u3_n119, u0_u2_u3_n120, u0_u2_u3_n121, u0_u2_u3_n122, u0_u2_u3_n123, 
       u0_u2_u3_n124, u0_u2_u3_n125, u0_u2_u3_n126, u0_u2_u3_n127, u0_u2_u3_n128, u0_u2_u3_n129, u0_u2_u3_n130, u0_u2_u3_n131, u0_u2_u3_n132, 
       u0_u2_u3_n133, u0_u2_u3_n134, u0_u2_u3_n135, u0_u2_u3_n136, u0_u2_u3_n137, u0_u2_u3_n138, u0_u2_u3_n139, u0_u2_u3_n140, u0_u2_u3_n141, 
       u0_u2_u3_n142, u0_u2_u3_n143, u0_u2_u3_n144, u0_u2_u3_n145, u0_u2_u3_n146, u0_u2_u3_n147, u0_u2_u3_n148, u0_u2_u3_n149, u0_u2_u3_n150, 
       u0_u2_u3_n151, u0_u2_u3_n152, u0_u2_u3_n153, u0_u2_u3_n154, u0_u2_u3_n155, u0_u2_u3_n156, u0_u2_u3_n157, u0_u2_u3_n158, u0_u2_u3_n159, 
       u0_u2_u3_n160, u0_u2_u3_n161, u0_u2_u3_n162, u0_u2_u3_n163, u0_u2_u3_n164, u0_u2_u3_n165, u0_u2_u3_n166, u0_u2_u3_n167, u0_u2_u3_n168, 
       u0_u2_u3_n169, u0_u2_u3_n170, u0_u2_u3_n171, u0_u2_u3_n172, u0_u2_u3_n173, u0_u2_u3_n174, u0_u2_u3_n175, u0_u2_u3_n176, u0_u2_u3_n177, 
       u0_u2_u3_n178, u0_u2_u3_n179, u0_u2_u3_n180, u0_u2_u3_n181, u0_u2_u3_n182, u0_u2_u3_n183, u0_u2_u3_n184, u0_u2_u3_n185, u0_u2_u3_n186, 
       u0_u2_u3_n94, u0_u2_u3_n95, u0_u2_u3_n96, u0_u2_u3_n97, u0_u2_u3_n98, u0_u2_u3_n99, u0_u2_u5_n100, u0_u2_u5_n101, u0_u2_u5_n102, 
       u0_u2_u5_n103, u0_u2_u5_n104, u0_u2_u5_n105, u0_u2_u5_n106, u0_u2_u5_n107, u0_u2_u5_n108, u0_u2_u5_n109, u0_u2_u5_n110, u0_u2_u5_n111, 
       u0_u2_u5_n112, u0_u2_u5_n113, u0_u2_u5_n114, u0_u2_u5_n115, u0_u2_u5_n116, u0_u2_u5_n117, u0_u2_u5_n118, u0_u2_u5_n119, u0_u2_u5_n120, 
       u0_u2_u5_n121, u0_u2_u5_n122, u0_u2_u5_n123, u0_u2_u5_n124, u0_u2_u5_n125, u0_u2_u5_n126, u0_u2_u5_n127, u0_u2_u5_n128, u0_u2_u5_n129, 
       u0_u2_u5_n130, u0_u2_u5_n131, u0_u2_u5_n132, u0_u2_u5_n133, u0_u2_u5_n134, u0_u2_u5_n135, u0_u2_u5_n136, u0_u2_u5_n137, u0_u2_u5_n138, 
       u0_u2_u5_n139, u0_u2_u5_n140, u0_u2_u5_n141, u0_u2_u5_n142, u0_u2_u5_n143, u0_u2_u5_n144, u0_u2_u5_n145, u0_u2_u5_n146, u0_u2_u5_n147, 
       u0_u2_u5_n148, u0_u2_u5_n149, u0_u2_u5_n150, u0_u2_u5_n151, u0_u2_u5_n152, u0_u2_u5_n153, u0_u2_u5_n154, u0_u2_u5_n155, u0_u2_u5_n156, 
       u0_u2_u5_n157, u0_u2_u5_n158, u0_u2_u5_n159, u0_u2_u5_n160, u0_u2_u5_n161, u0_u2_u5_n162, u0_u2_u5_n163, u0_u2_u5_n164, u0_u2_u5_n165, 
       u0_u2_u5_n166, u0_u2_u5_n167, u0_u2_u5_n168, u0_u2_u5_n169, u0_u2_u5_n170, u0_u2_u5_n171, u0_u2_u5_n172, u0_u2_u5_n173, u0_u2_u5_n174, 
       u0_u2_u5_n175, u0_u2_u5_n176, u0_u2_u5_n177, u0_u2_u5_n178, u0_u2_u5_n179, u0_u2_u5_n180, u0_u2_u5_n181, u0_u2_u5_n182, u0_u2_u5_n183, 
       u0_u2_u5_n184, u0_u2_u5_n185, u0_u2_u5_n186, u0_u2_u5_n187, u0_u2_u5_n188, u0_u2_u5_n189, u0_u2_u5_n190, u0_u2_u5_n191, u0_u2_u5_n192, 
       u0_u2_u5_n193, u0_u2_u5_n194, u0_u2_u5_n195, u0_u2_u5_n196, u0_u2_u5_n99, u0_u3_X_31, u0_u3_X_32, u0_u3_X_33, u0_u3_X_34, 
       u0_u3_X_35, u0_u3_X_36, u0_u3_u5_n100, u0_u3_u5_n101, u0_u3_u5_n102, u0_u3_u5_n103, u0_u3_u5_n104, u0_u3_u5_n105, u0_u3_u5_n106, 
       u0_u3_u5_n107, u0_u3_u5_n108, u0_u3_u5_n109, u0_u3_u5_n110, u0_u3_u5_n111, u0_u3_u5_n112, u0_u3_u5_n113, u0_u3_u5_n114, u0_u3_u5_n115, 
       u0_u3_u5_n116, u0_u3_u5_n117, u0_u3_u5_n118, u0_u3_u5_n119, u0_u3_u5_n120, u0_u3_u5_n121, u0_u3_u5_n122, u0_u3_u5_n123, u0_u3_u5_n124, 
       u0_u3_u5_n125, u0_u3_u5_n126, u0_u3_u5_n127, u0_u3_u5_n128, u0_u3_u5_n129, u0_u3_u5_n130, u0_u3_u5_n131, u0_u3_u5_n132, u0_u3_u5_n133, 
       u0_u3_u5_n134, u0_u3_u5_n135, u0_u3_u5_n136, u0_u3_u5_n137, u0_u3_u5_n138, u0_u3_u5_n139, u0_u3_u5_n140, u0_u3_u5_n141, u0_u3_u5_n142, 
       u0_u3_u5_n143, u0_u3_u5_n144, u0_u3_u5_n145, u0_u3_u5_n146, u0_u3_u5_n147, u0_u3_u5_n148, u0_u3_u5_n149, u0_u3_u5_n150, u0_u3_u5_n151, 
       u0_u3_u5_n152, u0_u3_u5_n153, u0_u3_u5_n154, u0_u3_u5_n155, u0_u3_u5_n156, u0_u3_u5_n157, u0_u3_u5_n158, u0_u3_u5_n159, u0_u3_u5_n160, 
       u0_u3_u5_n161, u0_u3_u5_n162, u0_u3_u5_n163, u0_u3_u5_n164, u0_u3_u5_n165, u0_u3_u5_n166, u0_u3_u5_n167, u0_u3_u5_n168, u0_u3_u5_n169, 
       u0_u3_u5_n170, u0_u3_u5_n171, u0_u3_u5_n172, u0_u3_u5_n173, u0_u3_u5_n174, u0_u3_u5_n175, u0_u3_u5_n176, u0_u3_u5_n177, u0_u3_u5_n178, 
       u0_u3_u5_n179, u0_u3_u5_n180, u0_u3_u5_n181, u0_u3_u5_n182, u0_u3_u5_n183, u0_u3_u5_n184, u0_u3_u5_n185, u0_u3_u5_n186, u0_u3_u5_n187, 
       u0_u3_u5_n188, u0_u3_u5_n189, u0_u3_u5_n190, u0_u3_u5_n191, u0_u3_u5_n192, u0_u3_u5_n193, u0_u3_u5_n194, u0_u3_u5_n195, u0_u3_u5_n196, 
       u0_u3_u5_n99, u0_u6_X_1, u0_u6_X_2, u0_u6_X_3, u0_u6_X_31, u0_u6_X_32, u0_u6_X_33, u0_u6_X_34, u0_u6_X_35, 
       u0_u6_X_36, u0_u6_X_37, u0_u6_X_38, u0_u6_X_39, u0_u6_X_4, u0_u6_X_40, u0_u6_X_41, u0_u6_X_42, u0_u6_X_43, 
       u0_u6_X_44, u0_u6_X_45, u0_u6_X_46, u0_u6_X_47, u0_u6_X_48, u0_u6_X_5, u0_u6_u0_n100, u0_u6_u0_n101, u0_u6_u0_n102, 
       u0_u6_u0_n103, u0_u6_u0_n104, u0_u6_u0_n105, u0_u6_u0_n106, u0_u6_u0_n107, u0_u6_u0_n108, u0_u6_u0_n109, u0_u6_u0_n110, u0_u6_u0_n111, 
       u0_u6_u0_n112, u0_u6_u0_n113, u0_u6_u0_n114, u0_u6_u0_n115, u0_u6_u0_n116, u0_u6_u0_n117, u0_u6_u0_n118, u0_u6_u0_n119, u0_u6_u0_n120, 
       u0_u6_u0_n121, u0_u6_u0_n122, u0_u6_u0_n123, u0_u6_u0_n124, u0_u6_u0_n125, u0_u6_u0_n126, u0_u6_u0_n127, u0_u6_u0_n128, u0_u6_u0_n129, 
       u0_u6_u0_n130, u0_u6_u0_n131, u0_u6_u0_n132, u0_u6_u0_n133, u0_u6_u0_n134, u0_u6_u0_n135, u0_u6_u0_n136, u0_u6_u0_n137, u0_u6_u0_n138, 
       u0_u6_u0_n139, u0_u6_u0_n140, u0_u6_u0_n141, u0_u6_u0_n142, u0_u6_u0_n143, u0_u6_u0_n144, u0_u6_u0_n145, u0_u6_u0_n146, u0_u6_u0_n147, 
       u0_u6_u0_n148, u0_u6_u0_n149, u0_u6_u0_n150, u0_u6_u0_n151, u0_u6_u0_n152, u0_u6_u0_n153, u0_u6_u0_n154, u0_u6_u0_n155, u0_u6_u0_n156, 
       u0_u6_u0_n157, u0_u6_u0_n158, u0_u6_u0_n159, u0_u6_u0_n160, u0_u6_u0_n161, u0_u6_u0_n162, u0_u6_u0_n163, u0_u6_u0_n164, u0_u6_u0_n165, 
       u0_u6_u0_n166, u0_u6_u0_n167, u0_u6_u0_n168, u0_u6_u0_n169, u0_u6_u0_n170, u0_u6_u0_n171, u0_u6_u0_n172, u0_u6_u0_n173, u0_u6_u0_n174, 
       u0_u6_u0_n88, u0_u6_u0_n89, u0_u6_u0_n90, u0_u6_u0_n91, u0_u6_u0_n92, u0_u6_u0_n93, u0_u6_u0_n94, u0_u6_u0_n95, u0_u6_u0_n96, 
       u0_u6_u0_n97, u0_u6_u0_n98, u0_u6_u0_n99, u0_u6_u5_n100, u0_u6_u5_n101, u0_u6_u5_n102, u0_u6_u5_n103, u0_u6_u5_n104, u0_u6_u5_n105, 
       u0_u6_u5_n106, u0_u6_u5_n107, u0_u6_u5_n108, u0_u6_u5_n109, u0_u6_u5_n110, u0_u6_u5_n111, u0_u6_u5_n112, u0_u6_u5_n113, u0_u6_u5_n114, 
       u0_u6_u5_n115, u0_u6_u5_n116, u0_u6_u5_n117, u0_u6_u5_n118, u0_u6_u5_n119, u0_u6_u5_n120, u0_u6_u5_n121, u0_u6_u5_n122, u0_u6_u5_n123, 
       u0_u6_u5_n124, u0_u6_u5_n125, u0_u6_u5_n126, u0_u6_u5_n127, u0_u6_u5_n128, u0_u6_u5_n129, u0_u6_u5_n130, u0_u6_u5_n131, u0_u6_u5_n132, 
       u0_u6_u5_n133, u0_u6_u5_n134, u0_u6_u5_n135, u0_u6_u5_n136, u0_u6_u5_n137, u0_u6_u5_n138, u0_u6_u5_n139, u0_u6_u5_n140, u0_u6_u5_n141, 
       u0_u6_u5_n142, u0_u6_u5_n143, u0_u6_u5_n144, u0_u6_u5_n145, u0_u6_u5_n146, u0_u6_u5_n147, u0_u6_u5_n148, u0_u6_u5_n149, u0_u6_u5_n150, 
       u0_u6_u5_n151, u0_u6_u5_n152, u0_u6_u5_n153, u0_u6_u5_n154, u0_u6_u5_n155, u0_u6_u5_n156, u0_u6_u5_n157, u0_u6_u5_n158, u0_u6_u5_n159, 
       u0_u6_u5_n160, u0_u6_u5_n161, u0_u6_u5_n162, u0_u6_u5_n163, u0_u6_u5_n164, u0_u6_u5_n165, u0_u6_u5_n166, u0_u6_u5_n167, u0_u6_u5_n168, 
       u0_u6_u5_n169, u0_u6_u5_n170, u0_u6_u5_n171, u0_u6_u5_n172, u0_u6_u5_n173, u0_u6_u5_n174, u0_u6_u5_n175, u0_u6_u5_n176, u0_u6_u5_n177, 
       u0_u6_u5_n178, u0_u6_u5_n179, u0_u6_u5_n180, u0_u6_u5_n181, u0_u6_u5_n182, u0_u6_u5_n183, u0_u6_u5_n184, u0_u6_u5_n185, u0_u6_u5_n186, 
       u0_u6_u5_n187, u0_u6_u5_n188, u0_u6_u5_n189, u0_u6_u5_n190, u0_u6_u5_n191, u0_u6_u5_n192, u0_u6_u5_n193, u0_u6_u5_n194, u0_u6_u5_n195, 
       u0_u6_u5_n196, u0_u6_u5_n99, u0_u6_u6_n100, u0_u6_u6_n101, u0_u6_u6_n102, u0_u6_u6_n103, u0_u6_u6_n104, u0_u6_u6_n105, u0_u6_u6_n106, 
       u0_u6_u6_n107, u0_u6_u6_n108, u0_u6_u6_n109, u0_u6_u6_n110, u0_u6_u6_n111, u0_u6_u6_n112, u0_u6_u6_n113, u0_u6_u6_n114, u0_u6_u6_n115, 
       u0_u6_u6_n116, u0_u6_u6_n117, u0_u6_u6_n118, u0_u6_u6_n119, u0_u6_u6_n120, u0_u6_u6_n121, u0_u6_u6_n122, u0_u6_u6_n123, u0_u6_u6_n124, 
       u0_u6_u6_n125, u0_u6_u6_n126, u0_u6_u6_n127, u0_u6_u6_n128, u0_u6_u6_n129, u0_u6_u6_n130, u0_u6_u6_n131, u0_u6_u6_n132, u0_u6_u6_n133, 
       u0_u6_u6_n134, u0_u6_u6_n135, u0_u6_u6_n136, u0_u6_u6_n137, u0_u6_u6_n138, u0_u6_u6_n139, u0_u6_u6_n140, u0_u6_u6_n141, u0_u6_u6_n142, 
       u0_u6_u6_n143, u0_u6_u6_n144, u0_u6_u6_n145, u0_u6_u6_n146, u0_u6_u6_n147, u0_u6_u6_n148, u0_u6_u6_n149, u0_u6_u6_n150, u0_u6_u6_n151, 
       u0_u6_u6_n152, u0_u6_u6_n153, u0_u6_u6_n154, u0_u6_u6_n155, u0_u6_u6_n156, u0_u6_u6_n157, u0_u6_u6_n158, u0_u6_u6_n159, u0_u6_u6_n160, 
       u0_u6_u6_n161, u0_u6_u6_n162, u0_u6_u6_n163, u0_u6_u6_n164, u0_u6_u6_n165, u0_u6_u6_n166, u0_u6_u6_n167, u0_u6_u6_n168, u0_u6_u6_n169, 
       u0_u6_u6_n170, u0_u6_u6_n171, u0_u6_u6_n172, u0_u6_u6_n173, u0_u6_u6_n174, u0_u6_u6_n88, u0_u6_u6_n89, u0_u6_u6_n90, u0_u6_u6_n91, 
       u0_u6_u6_n92, u0_u6_u6_n93, u0_u6_u6_n94, u0_u6_u6_n95, u0_u6_u6_n96, u0_u6_u6_n97, u0_u6_u6_n98, u0_u6_u6_n99, u0_u6_u7_n100, 
       u0_u6_u7_n101, u0_u6_u7_n102, u0_u6_u7_n103, u0_u6_u7_n104, u0_u6_u7_n105, u0_u6_u7_n106, u0_u6_u7_n107, u0_u6_u7_n108, u0_u6_u7_n109, 
       u0_u6_u7_n110, u0_u6_u7_n111, u0_u6_u7_n112, u0_u6_u7_n113, u0_u6_u7_n114, u0_u6_u7_n115, u0_u6_u7_n116, u0_u6_u7_n117, u0_u6_u7_n118, 
       u0_u6_u7_n119, u0_u6_u7_n120, u0_u6_u7_n121, u0_u6_u7_n122, u0_u6_u7_n123, u0_u6_u7_n124, u0_u6_u7_n125, u0_u6_u7_n126, u0_u6_u7_n127, 
       u0_u6_u7_n128, u0_u6_u7_n129, u0_u6_u7_n130, u0_u6_u7_n131, u0_u6_u7_n132, u0_u6_u7_n133, u0_u6_u7_n134, u0_u6_u7_n135, u0_u6_u7_n136, 
       u0_u6_u7_n137, u0_u6_u7_n138, u0_u6_u7_n139, u0_u6_u7_n140, u0_u6_u7_n141, u0_u6_u7_n142, u0_u6_u7_n143, u0_u6_u7_n144, u0_u6_u7_n145, 
       u0_u6_u7_n146, u0_u6_u7_n147, u0_u6_u7_n148, u0_u6_u7_n149, u0_u6_u7_n150, u0_u6_u7_n151, u0_u6_u7_n152, u0_u6_u7_n153, u0_u6_u7_n154, 
       u0_u6_u7_n155, u0_u6_u7_n156, u0_u6_u7_n157, u0_u6_u7_n158, u0_u6_u7_n159, u0_u6_u7_n160, u0_u6_u7_n161, u0_u6_u7_n162, u0_u6_u7_n163, 
       u0_u6_u7_n164, u0_u6_u7_n165, u0_u6_u7_n166, u0_u6_u7_n167, u0_u6_u7_n168, u0_u6_u7_n169, u0_u6_u7_n170, u0_u6_u7_n171, u0_u6_u7_n172, 
       u0_u6_u7_n173, u0_u6_u7_n174, u0_u6_u7_n175, u0_u6_u7_n176, u0_u6_u7_n177, u0_u6_u7_n178, u0_u6_u7_n179, u0_u6_u7_n180, u0_u6_u7_n91, 
       u0_u6_u7_n92, u0_u6_u7_n93, u0_u6_u7_n94, u0_u6_u7_n95, u0_u6_u7_n96, u0_u6_u7_n97, u0_u6_u7_n98, u0_u6_u7_n99, u0_u9_X_1, 
       u0_u9_X_2, u0_u9_X_3, u0_u9_X_4, u0_u9_X_5, u0_u9_X_6, u0_u9_u0_n100, u0_u9_u0_n101, u0_u9_u0_n102, u0_u9_u0_n103, 
       u0_u9_u0_n104, u0_u9_u0_n105, u0_u9_u0_n106, u0_u9_u0_n107, u0_u9_u0_n108, u0_u9_u0_n109, u0_u9_u0_n110, u0_u9_u0_n111, u0_u9_u0_n112, 
       u0_u9_u0_n113, u0_u9_u0_n114, u0_u9_u0_n115, u0_u9_u0_n116, u0_u9_u0_n117, u0_u9_u0_n118, u0_u9_u0_n119, u0_u9_u0_n120, u0_u9_u0_n121, 
       u0_u9_u0_n122, u0_u9_u0_n123, u0_u9_u0_n124, u0_u9_u0_n125, u0_u9_u0_n126, u0_u9_u0_n127, u0_u9_u0_n128, u0_u9_u0_n129, u0_u9_u0_n130, 
       u0_u9_u0_n131, u0_u9_u0_n132, u0_u9_u0_n133, u0_u9_u0_n134, u0_u9_u0_n135, u0_u9_u0_n136, u0_u9_u0_n137, u0_u9_u0_n138, u0_u9_u0_n139, 
       u0_u9_u0_n140, u0_u9_u0_n141, u0_u9_u0_n142, u0_u9_u0_n143, u0_u9_u0_n144, u0_u9_u0_n145, u0_u9_u0_n146, u0_u9_u0_n147, u0_u9_u0_n148, 
       u0_u9_u0_n149, u0_u9_u0_n150, u0_u9_u0_n151, u0_u9_u0_n152, u0_u9_u0_n153, u0_u9_u0_n154, u0_u9_u0_n155, u0_u9_u0_n156, u0_u9_u0_n157, 
       u0_u9_u0_n158, u0_u9_u0_n159, u0_u9_u0_n160, u0_u9_u0_n161, u0_u9_u0_n162, u0_u9_u0_n163, u0_u9_u0_n164, u0_u9_u0_n165, u0_u9_u0_n166, 
       u0_u9_u0_n167, u0_u9_u0_n168, u0_u9_u0_n169, u0_u9_u0_n170, u0_u9_u0_n171, u0_u9_u0_n172, u0_u9_u0_n173, u0_u9_u0_n174, u0_u9_u0_n88, 
       u0_u9_u0_n89, u0_u9_u0_n90, u0_u9_u0_n91, u0_u9_u0_n92, u0_u9_u0_n93, u0_u9_u0_n94, u0_u9_u0_n95, u0_u9_u0_n96, u0_u9_u0_n97, 
       u0_u9_u0_n98, u0_u9_u0_n99, u0_uk_n1003, u0_uk_n1015, u0_uk_n767, u0_uk_n768, u0_uk_n769, u0_uk_n771, u0_uk_n772, 
       u0_uk_n781, u0_uk_n840, u0_uk_n846, u0_uk_n847, u0_uk_n851, u0_uk_n858, u0_uk_n865, u0_uk_n866, u0_uk_n868, 
       u0_uk_n902, u0_uk_n905, u0_uk_n907, u0_uk_n908, u0_uk_n909, u0_uk_n966, u0_uk_n979, u0_uk_n980, u0_uk_n982, 
       u0_uk_n983, u0_uk_n984, u0_uk_n987, u0_uk_n988, u0_uk_n991, u0_uk_n992, u1_K13_10, u1_K13_11, u1_K13_13, 
       u1_K13_15, u1_K4_29, u1_K4_31, u1_K6_10, u1_K6_9, u1_K8_34, u1_out12_11, u1_out12_13, u1_out12_16, 
       u1_out12_18, u1_out12_19, u1_out12_2, u1_out12_24, u1_out12_28, u1_out12_29, u1_out12_30, u1_out12_4, u1_out12_6, 
       u1_out13_16, u1_out13_17, u1_out13_23, u1_out13_24, u1_out13_30, u1_out13_31, u1_out13_6, u1_out13_9, u1_out14_13, 
       u1_out14_18, u1_out14_2, u1_out14_28, u1_out15_15, u1_out15_21, u1_out15_27, u1_out15_5, u1_out1_11, u1_out1_19, 
       u1_out1_29, u1_out1_4, u1_out2_14, u1_out2_17, u1_out2_23, u1_out2_25, u1_out2_3, u1_out2_31, u1_out2_8, 
       u1_out2_9, u1_out3_11, u1_out3_14, u1_out3_15, u1_out3_16, u1_out3_19, u1_out3_21, u1_out3_24, u1_out3_25, 
       u1_out3_27, u1_out3_29, u1_out3_3, u1_out3_30, u1_out3_4, u1_out3_5, u1_out3_6, u1_out3_8, u1_out5_13, 
       u1_out5_18, u1_out5_2, u1_out5_28, u1_out7_11, u1_out7_19, u1_out7_29, u1_out7_4, u1_u12_X_10, u1_u12_X_11, 
       u1_u12_X_13, u1_u12_X_15, u1_u12_X_16, u1_u12_X_33, u1_u12_X_34, u1_u12_X_9, u1_u12_u1_n100, u1_u12_u1_n101, u1_u12_u1_n102, 
       u1_u12_u1_n103, u1_u12_u1_n104, u1_u12_u1_n105, u1_u12_u1_n106, u1_u12_u1_n107, u1_u12_u1_n108, u1_u12_u1_n109, u1_u12_u1_n110, u1_u12_u1_n111, 
       u1_u12_u1_n112, u1_u12_u1_n113, u1_u12_u1_n114, u1_u12_u1_n115, u1_u12_u1_n116, u1_u12_u1_n117, u1_u12_u1_n118, u1_u12_u1_n119, u1_u12_u1_n120, 
       u1_u12_u1_n121, u1_u12_u1_n122, u1_u12_u1_n123, u1_u12_u1_n124, u1_u12_u1_n125, u1_u12_u1_n126, u1_u12_u1_n127, u1_u12_u1_n128, u1_u12_u1_n129, 
       u1_u12_u1_n130, u1_u12_u1_n131, u1_u12_u1_n132, u1_u12_u1_n133, u1_u12_u1_n134, u1_u12_u1_n135, u1_u12_u1_n136, u1_u12_u1_n137, u1_u12_u1_n138, 
       u1_u12_u1_n139, u1_u12_u1_n140, u1_u12_u1_n141, u1_u12_u1_n142, u1_u12_u1_n143, u1_u12_u1_n144, u1_u12_u1_n145, u1_u12_u1_n146, u1_u12_u1_n147, 
       u1_u12_u1_n148, u1_u12_u1_n149, u1_u12_u1_n150, u1_u12_u1_n151, u1_u12_u1_n152, u1_u12_u1_n153, u1_u12_u1_n154, u1_u12_u1_n155, u1_u12_u1_n156, 
       u1_u12_u1_n157, u1_u12_u1_n158, u1_u12_u1_n159, u1_u12_u1_n160, u1_u12_u1_n161, u1_u12_u1_n162, u1_u12_u1_n163, u1_u12_u1_n164, u1_u12_u1_n165, 
       u1_u12_u1_n166, u1_u12_u1_n167, u1_u12_u1_n168, u1_u12_u1_n169, u1_u12_u1_n170, u1_u12_u1_n171, u1_u12_u1_n172, u1_u12_u1_n173, u1_u12_u1_n174, 
       u1_u12_u1_n175, u1_u12_u1_n176, u1_u12_u1_n177, u1_u12_u1_n178, u1_u12_u1_n179, u1_u12_u1_n180, u1_u12_u1_n181, u1_u12_u1_n182, u1_u12_u1_n183, 
       u1_u12_u1_n184, u1_u12_u1_n185, u1_u12_u1_n186, u1_u12_u1_n187, u1_u12_u1_n188, u1_u12_u1_n95, u1_u12_u1_n96, u1_u12_u1_n97, u1_u12_u1_n98, 
       u1_u12_u1_n99, u1_u12_u2_n100, u1_u12_u2_n101, u1_u12_u2_n102, u1_u12_u2_n103, u1_u12_u2_n104, u1_u12_u2_n105, u1_u12_u2_n106, u1_u12_u2_n107, 
       u1_u12_u2_n108, u1_u12_u2_n109, u1_u12_u2_n110, u1_u12_u2_n111, u1_u12_u2_n112, u1_u12_u2_n113, u1_u12_u2_n114, u1_u12_u2_n115, u1_u12_u2_n116, 
       u1_u12_u2_n117, u1_u12_u2_n118, u1_u12_u2_n119, u1_u12_u2_n120, u1_u12_u2_n121, u1_u12_u2_n122, u1_u12_u2_n123, u1_u12_u2_n124, u1_u12_u2_n125, 
       u1_u12_u2_n126, u1_u12_u2_n127, u1_u12_u2_n128, u1_u12_u2_n129, u1_u12_u2_n130, u1_u12_u2_n131, u1_u12_u2_n132, u1_u12_u2_n133, u1_u12_u2_n134, 
       u1_u12_u2_n135, u1_u12_u2_n136, u1_u12_u2_n137, u1_u12_u2_n138, u1_u12_u2_n139, u1_u12_u2_n140, u1_u12_u2_n141, u1_u12_u2_n142, u1_u12_u2_n143, 
       u1_u12_u2_n144, u1_u12_u2_n145, u1_u12_u2_n146, u1_u12_u2_n147, u1_u12_u2_n148, u1_u12_u2_n149, u1_u12_u2_n150, u1_u12_u2_n151, u1_u12_u2_n152, 
       u1_u12_u2_n153, u1_u12_u2_n154, u1_u12_u2_n155, u1_u12_u2_n156, u1_u12_u2_n157, u1_u12_u2_n158, u1_u12_u2_n159, u1_u12_u2_n160, u1_u12_u2_n161, 
       u1_u12_u2_n162, u1_u12_u2_n163, u1_u12_u2_n164, u1_u12_u2_n165, u1_u12_u2_n166, u1_u12_u2_n167, u1_u12_u2_n168, u1_u12_u2_n169, u1_u12_u2_n170, 
       u1_u12_u2_n171, u1_u12_u2_n172, u1_u12_u2_n173, u1_u12_u2_n174, u1_u12_u2_n175, u1_u12_u2_n176, u1_u12_u2_n177, u1_u12_u2_n178, u1_u12_u2_n179, 
       u1_u12_u2_n180, u1_u12_u2_n181, u1_u12_u2_n182, u1_u12_u2_n183, u1_u12_u2_n184, u1_u12_u2_n185, u1_u12_u2_n186, u1_u12_u2_n187, u1_u12_u2_n188, 
       u1_u12_u2_n95, u1_u12_u2_n96, u1_u12_u2_n97, u1_u12_u2_n98, u1_u12_u2_n99, u1_u12_u5_n100, u1_u12_u5_n101, u1_u12_u5_n102, u1_u12_u5_n103, 
       u1_u12_u5_n104, u1_u12_u5_n105, u1_u12_u5_n106, u1_u12_u5_n107, u1_u12_u5_n108, u1_u12_u5_n109, u1_u12_u5_n110, u1_u12_u5_n111, u1_u12_u5_n112, 
       u1_u12_u5_n113, u1_u12_u5_n114, u1_u12_u5_n115, u1_u12_u5_n116, u1_u12_u5_n117, u1_u12_u5_n118, u1_u12_u5_n119, u1_u12_u5_n120, u1_u12_u5_n121, 
       u1_u12_u5_n122, u1_u12_u5_n123, u1_u12_u5_n124, u1_u12_u5_n125, u1_u12_u5_n126, u1_u12_u5_n127, u1_u12_u5_n128, u1_u12_u5_n129, u1_u12_u5_n130, 
       u1_u12_u5_n131, u1_u12_u5_n132, u1_u12_u5_n133, u1_u12_u5_n134, u1_u12_u5_n135, u1_u12_u5_n136, u1_u12_u5_n137, u1_u12_u5_n138, u1_u12_u5_n139, 
       u1_u12_u5_n140, u1_u12_u5_n141, u1_u12_u5_n142, u1_u12_u5_n143, u1_u12_u5_n144, u1_u12_u5_n145, u1_u12_u5_n146, u1_u12_u5_n147, u1_u12_u5_n148, 
       u1_u12_u5_n149, u1_u12_u5_n150, u1_u12_u5_n151, u1_u12_u5_n152, u1_u12_u5_n153, u1_u12_u5_n154, u1_u12_u5_n155, u1_u12_u5_n156, u1_u12_u5_n157, 
       u1_u12_u5_n158, u1_u12_u5_n159, u1_u12_u5_n160, u1_u12_u5_n161, u1_u12_u5_n162, u1_u12_u5_n163, u1_u12_u5_n164, u1_u12_u5_n165, u1_u12_u5_n166, 
       u1_u12_u5_n167, u1_u12_u5_n168, u1_u12_u5_n169, u1_u12_u5_n170, u1_u12_u5_n171, u1_u12_u5_n172, u1_u12_u5_n173, u1_u12_u5_n174, u1_u12_u5_n175, 
       u1_u12_u5_n176, u1_u12_u5_n177, u1_u12_u5_n178, u1_u12_u5_n179, u1_u12_u5_n180, u1_u12_u5_n181, u1_u12_u5_n182, u1_u12_u5_n183, u1_u12_u5_n184, 
       u1_u12_u5_n185, u1_u12_u5_n186, u1_u12_u5_n187, u1_u12_u5_n188, u1_u12_u5_n189, u1_u12_u5_n190, u1_u12_u5_n191, u1_u12_u5_n192, u1_u12_u5_n193, 
       u1_u12_u5_n194, u1_u12_u5_n195, u1_u12_u5_n196, u1_u12_u5_n99, u1_u13_X_15, u1_u13_X_16, u1_u13_X_3, u1_u13_X_4, u1_u13_u0_n100, 
       u1_u13_u0_n101, u1_u13_u0_n102, u1_u13_u0_n103, u1_u13_u0_n104, u1_u13_u0_n105, u1_u13_u0_n106, u1_u13_u0_n107, u1_u13_u0_n108, u1_u13_u0_n109, 
       u1_u13_u0_n110, u1_u13_u0_n111, u1_u13_u0_n112, u1_u13_u0_n113, u1_u13_u0_n114, u1_u13_u0_n115, u1_u13_u0_n116, u1_u13_u0_n117, u1_u13_u0_n118, 
       u1_u13_u0_n119, u1_u13_u0_n120, u1_u13_u0_n121, u1_u13_u0_n122, u1_u13_u0_n123, u1_u13_u0_n124, u1_u13_u0_n125, u1_u13_u0_n126, u1_u13_u0_n127, 
       u1_u13_u0_n128, u1_u13_u0_n129, u1_u13_u0_n130, u1_u13_u0_n131, u1_u13_u0_n132, u1_u13_u0_n133, u1_u13_u0_n134, u1_u13_u0_n135, u1_u13_u0_n136, 
       u1_u13_u0_n137, u1_u13_u0_n138, u1_u13_u0_n139, u1_u13_u0_n140, u1_u13_u0_n141, u1_u13_u0_n142, u1_u13_u0_n143, u1_u13_u0_n144, u1_u13_u0_n145, 
       u1_u13_u0_n146, u1_u13_u0_n147, u1_u13_u0_n148, u1_u13_u0_n149, u1_u13_u0_n150, u1_u13_u0_n151, u1_u13_u0_n152, u1_u13_u0_n153, u1_u13_u0_n154, 
       u1_u13_u0_n155, u1_u13_u0_n156, u1_u13_u0_n157, u1_u13_u0_n158, u1_u13_u0_n159, u1_u13_u0_n160, u1_u13_u0_n161, u1_u13_u0_n162, u1_u13_u0_n163, 
       u1_u13_u0_n164, u1_u13_u0_n165, u1_u13_u0_n166, u1_u13_u0_n167, u1_u13_u0_n168, u1_u13_u0_n169, u1_u13_u0_n170, u1_u13_u0_n171, u1_u13_u0_n172, 
       u1_u13_u0_n173, u1_u13_u0_n174, u1_u13_u0_n88, u1_u13_u0_n89, u1_u13_u0_n90, u1_u13_u0_n91, u1_u13_u0_n92, u1_u13_u0_n93, u1_u13_u0_n94, 
       u1_u13_u0_n95, u1_u13_u0_n96, u1_u13_u0_n97, u1_u13_u0_n98, u1_u13_u0_n99, u1_u13_u2_n100, u1_u13_u2_n101, u1_u13_u2_n102, u1_u13_u2_n103, 
       u1_u13_u2_n104, u1_u13_u2_n105, u1_u13_u2_n106, u1_u13_u2_n107, u1_u13_u2_n108, u1_u13_u2_n109, u1_u13_u2_n110, u1_u13_u2_n111, u1_u13_u2_n112, 
       u1_u13_u2_n113, u1_u13_u2_n114, u1_u13_u2_n115, u1_u13_u2_n116, u1_u13_u2_n117, u1_u13_u2_n118, u1_u13_u2_n119, u1_u13_u2_n120, u1_u13_u2_n121, 
       u1_u13_u2_n122, u1_u13_u2_n123, u1_u13_u2_n124, u1_u13_u2_n125, u1_u13_u2_n126, u1_u13_u2_n127, u1_u13_u2_n128, u1_u13_u2_n129, u1_u13_u2_n130, 
       u1_u13_u2_n131, u1_u13_u2_n132, u1_u13_u2_n133, u1_u13_u2_n134, u1_u13_u2_n135, u1_u13_u2_n136, u1_u13_u2_n137, u1_u13_u2_n138, u1_u13_u2_n139, 
       u1_u13_u2_n140, u1_u13_u2_n141, u1_u13_u2_n142, u1_u13_u2_n143, u1_u13_u2_n144, u1_u13_u2_n145, u1_u13_u2_n146, u1_u13_u2_n147, u1_u13_u2_n148, 
       u1_u13_u2_n149, u1_u13_u2_n150, u1_u13_u2_n151, u1_u13_u2_n152, u1_u13_u2_n153, u1_u13_u2_n154, u1_u13_u2_n155, u1_u13_u2_n156, u1_u13_u2_n157, 
       u1_u13_u2_n158, u1_u13_u2_n159, u1_u13_u2_n160, u1_u13_u2_n161, u1_u13_u2_n162, u1_u13_u2_n163, u1_u13_u2_n164, u1_u13_u2_n165, u1_u13_u2_n166, 
       u1_u13_u2_n167, u1_u13_u2_n168, u1_u13_u2_n169, u1_u13_u2_n170, u1_u13_u2_n171, u1_u13_u2_n172, u1_u13_u2_n173, u1_u13_u2_n174, u1_u13_u2_n175, 
       u1_u13_u2_n176, u1_u13_u2_n177, u1_u13_u2_n178, u1_u13_u2_n179, u1_u13_u2_n180, u1_u13_u2_n181, u1_u13_u2_n182, u1_u13_u2_n183, u1_u13_u2_n184, 
       u1_u13_u2_n185, u1_u13_u2_n186, u1_u13_u2_n187, u1_u13_u2_n188, u1_u13_u2_n95, u1_u13_u2_n96, u1_u13_u2_n97, u1_u13_u2_n98, u1_u13_u2_n99, 
       u1_u14_X_10, u1_u14_X_9, u1_u14_u1_n100, u1_u14_u1_n101, u1_u14_u1_n102, u1_u14_u1_n103, u1_u14_u1_n104, u1_u14_u1_n105, u1_u14_u1_n106, 
       u1_u14_u1_n107, u1_u14_u1_n108, u1_u14_u1_n109, u1_u14_u1_n110, u1_u14_u1_n111, u1_u14_u1_n112, u1_u14_u1_n113, u1_u14_u1_n114, u1_u14_u1_n115, 
       u1_u14_u1_n116, u1_u14_u1_n117, u1_u14_u1_n118, u1_u14_u1_n119, u1_u14_u1_n120, u1_u14_u1_n121, u1_u14_u1_n122, u1_u14_u1_n123, u1_u14_u1_n124, 
       u1_u14_u1_n125, u1_u14_u1_n126, u1_u14_u1_n127, u1_u14_u1_n128, u1_u14_u1_n129, u1_u14_u1_n130, u1_u14_u1_n131, u1_u14_u1_n132, u1_u14_u1_n133, 
       u1_u14_u1_n134, u1_u14_u1_n135, u1_u14_u1_n136, u1_u14_u1_n137, u1_u14_u1_n138, u1_u14_u1_n139, u1_u14_u1_n140, u1_u14_u1_n141, u1_u14_u1_n142, 
       u1_u14_u1_n143, u1_u14_u1_n144, u1_u14_u1_n145, u1_u14_u1_n146, u1_u14_u1_n147, u1_u14_u1_n148, u1_u14_u1_n149, u1_u14_u1_n150, u1_u14_u1_n151, 
       u1_u14_u1_n152, u1_u14_u1_n153, u1_u14_u1_n154, u1_u14_u1_n155, u1_u14_u1_n156, u1_u14_u1_n157, u1_u14_u1_n158, u1_u14_u1_n159, u1_u14_u1_n160, 
       u1_u14_u1_n161, u1_u14_u1_n162, u1_u14_u1_n163, u1_u14_u1_n164, u1_u14_u1_n165, u1_u14_u1_n166, u1_u14_u1_n167, u1_u14_u1_n168, u1_u14_u1_n169, 
       u1_u14_u1_n170, u1_u14_u1_n171, u1_u14_u1_n172, u1_u14_u1_n173, u1_u14_u1_n174, u1_u14_u1_n175, u1_u14_u1_n176, u1_u14_u1_n177, u1_u14_u1_n178, 
       u1_u14_u1_n179, u1_u14_u1_n180, u1_u14_u1_n181, u1_u14_u1_n182, u1_u14_u1_n183, u1_u14_u1_n184, u1_u14_u1_n185, u1_u14_u1_n186, u1_u14_u1_n187, 
       u1_u14_u1_n188, u1_u14_u1_n95, u1_u14_u1_n96, u1_u14_u1_n97, u1_u14_u1_n98, u1_u14_u1_n99, u1_u15_X_45, u1_u15_X_46, u1_u15_u7_n100, 
       u1_u15_u7_n101, u1_u15_u7_n102, u1_u15_u7_n103, u1_u15_u7_n104, u1_u15_u7_n105, u1_u15_u7_n106, u1_u15_u7_n107, u1_u15_u7_n108, u1_u15_u7_n109, 
       u1_u15_u7_n110, u1_u15_u7_n111, u1_u15_u7_n112, u1_u15_u7_n113, u1_u15_u7_n114, u1_u15_u7_n115, u1_u15_u7_n116, u1_u15_u7_n117, u1_u15_u7_n118, 
       u1_u15_u7_n119, u1_u15_u7_n120, u1_u15_u7_n121, u1_u15_u7_n122, u1_u15_u7_n123, u1_u15_u7_n124, u1_u15_u7_n125, u1_u15_u7_n126, u1_u15_u7_n127, 
       u1_u15_u7_n128, u1_u15_u7_n129, u1_u15_u7_n130, u1_u15_u7_n131, u1_u15_u7_n132, u1_u15_u7_n133, u1_u15_u7_n134, u1_u15_u7_n135, u1_u15_u7_n136, 
       u1_u15_u7_n137, u1_u15_u7_n138, u1_u15_u7_n139, u1_u15_u7_n140, u1_u15_u7_n141, u1_u15_u7_n142, u1_u15_u7_n143, u1_u15_u7_n144, u1_u15_u7_n145, 
       u1_u15_u7_n146, u1_u15_u7_n147, u1_u15_u7_n148, u1_u15_u7_n149, u1_u15_u7_n150, u1_u15_u7_n151, u1_u15_u7_n152, u1_u15_u7_n153, u1_u15_u7_n154, 
       u1_u15_u7_n155, u1_u15_u7_n156, u1_u15_u7_n157, u1_u15_u7_n158, u1_u15_u7_n159, u1_u15_u7_n160, u1_u15_u7_n161, u1_u15_u7_n162, u1_u15_u7_n163, 
       u1_u15_u7_n164, u1_u15_u7_n165, u1_u15_u7_n166, u1_u15_u7_n167, u1_u15_u7_n168, u1_u15_u7_n169, u1_u15_u7_n170, u1_u15_u7_n171, u1_u15_u7_n172, 
       u1_u15_u7_n173, u1_u15_u7_n174, u1_u15_u7_n175, u1_u15_u7_n176, u1_u15_u7_n177, u1_u15_u7_n178, u1_u15_u7_n179, u1_u15_u7_n180, u1_u15_u7_n91, 
       u1_u15_u7_n92, u1_u15_u7_n93, u1_u15_u7_n94, u1_u15_u7_n95, u1_u15_u7_n96, u1_u15_u7_n97, u1_u15_u7_n98, u1_u15_u7_n99, u1_u1_X_33, 
       u1_u1_X_34, u1_u1_u5_n100, u1_u1_u5_n101, u1_u1_u5_n102, u1_u1_u5_n103, u1_u1_u5_n104, u1_u1_u5_n105, u1_u1_u5_n106, u1_u1_u5_n107, 
       u1_u1_u5_n108, u1_u1_u5_n109, u1_u1_u5_n110, u1_u1_u5_n111, u1_u1_u5_n112, u1_u1_u5_n113, u1_u1_u5_n114, u1_u1_u5_n115, u1_u1_u5_n116, 
       u1_u1_u5_n117, u1_u1_u5_n118, u1_u1_u5_n119, u1_u1_u5_n120, u1_u1_u5_n121, u1_u1_u5_n122, u1_u1_u5_n123, u1_u1_u5_n124, u1_u1_u5_n125, 
       u1_u1_u5_n126, u1_u1_u5_n127, u1_u1_u5_n128, u1_u1_u5_n129, u1_u1_u5_n130, u1_u1_u5_n131, u1_u1_u5_n132, u1_u1_u5_n133, u1_u1_u5_n134, 
       u1_u1_u5_n135, u1_u1_u5_n136, u1_u1_u5_n137, u1_u1_u5_n138, u1_u1_u5_n139, u1_u1_u5_n140, u1_u1_u5_n141, u1_u1_u5_n142, u1_u1_u5_n143, 
       u1_u1_u5_n144, u1_u1_u5_n145, u1_u1_u5_n146, u1_u1_u5_n147, u1_u1_u5_n148, u1_u1_u5_n149, u1_u1_u5_n150, u1_u1_u5_n151, u1_u1_u5_n152, 
       u1_u1_u5_n153, u1_u1_u5_n154, u1_u1_u5_n155, u1_u1_u5_n156, u1_u1_u5_n157, u1_u1_u5_n158, u1_u1_u5_n159, u1_u1_u5_n160, u1_u1_u5_n161, 
       u1_u1_u5_n162, u1_u1_u5_n163, u1_u1_u5_n164, u1_u1_u5_n165, u1_u1_u5_n166, u1_u1_u5_n167, u1_u1_u5_n168, u1_u1_u5_n169, u1_u1_u5_n170, 
       u1_u1_u5_n171, u1_u1_u5_n172, u1_u1_u5_n173, u1_u1_u5_n174, u1_u1_u5_n175, u1_u1_u5_n176, u1_u1_u5_n177, u1_u1_u5_n178, u1_u1_u5_n179, 
       u1_u1_u5_n180, u1_u1_u5_n181, u1_u1_u5_n182, u1_u1_u5_n183, u1_u1_u5_n184, u1_u1_u5_n185, u1_u1_u5_n186, u1_u1_u5_n187, u1_u1_u5_n188, 
       u1_u1_u5_n189, u1_u1_u5_n190, u1_u1_u5_n191, u1_u1_u5_n192, u1_u1_u5_n193, u1_u1_u5_n194, u1_u1_u5_n195, u1_u1_u5_n196, u1_u1_u5_n99, 
       u1_u2_X_27, u1_u2_X_28, u1_u2_X_3, u1_u2_X_4, u1_u2_u0_n100, u1_u2_u0_n101, u1_u2_u0_n102, u1_u2_u0_n103, u1_u2_u0_n104, 
       u1_u2_u0_n105, u1_u2_u0_n106, u1_u2_u0_n107, u1_u2_u0_n108, u1_u2_u0_n109, u1_u2_u0_n110, u1_u2_u0_n111, u1_u2_u0_n112, u1_u2_u0_n113, 
       u1_u2_u0_n114, u1_u2_u0_n115, u1_u2_u0_n116, u1_u2_u0_n117, u1_u2_u0_n118, u1_u2_u0_n119, u1_u2_u0_n120, u1_u2_u0_n121, u1_u2_u0_n122, 
       u1_u2_u0_n123, u1_u2_u0_n124, u1_u2_u0_n125, u1_u2_u0_n126, u1_u2_u0_n127, u1_u2_u0_n128, u1_u2_u0_n129, u1_u2_u0_n130, u1_u2_u0_n131, 
       u1_u2_u0_n132, u1_u2_u0_n133, u1_u2_u0_n134, u1_u2_u0_n135, u1_u2_u0_n136, u1_u2_u0_n137, u1_u2_u0_n138, u1_u2_u0_n139, u1_u2_u0_n140, 
       u1_u2_u0_n141, u1_u2_u0_n142, u1_u2_u0_n143, u1_u2_u0_n144, u1_u2_u0_n145, u1_u2_u0_n146, u1_u2_u0_n147, u1_u2_u0_n148, u1_u2_u0_n149, 
       u1_u2_u0_n150, u1_u2_u0_n151, u1_u2_u0_n152, u1_u2_u0_n153, u1_u2_u0_n154, u1_u2_u0_n155, u1_u2_u0_n156, u1_u2_u0_n157, u1_u2_u0_n158, 
       u1_u2_u0_n159, u1_u2_u0_n160, u1_u2_u0_n161, u1_u2_u0_n162, u1_u2_u0_n163, u1_u2_u0_n164, u1_u2_u0_n165, u1_u2_u0_n166, u1_u2_u0_n167, 
       u1_u2_u0_n168, u1_u2_u0_n169, u1_u2_u0_n170, u1_u2_u0_n171, u1_u2_u0_n172, u1_u2_u0_n173, u1_u2_u0_n174, u1_u2_u0_n88, u1_u2_u0_n89, 
       u1_u2_u0_n90, u1_u2_u0_n91, u1_u2_u0_n92, u1_u2_u0_n93, u1_u2_u0_n94, u1_u2_u0_n95, u1_u2_u0_n96, u1_u2_u0_n97, u1_u2_u0_n98, 
       u1_u2_u0_n99, u1_u2_u4_n100, u1_u2_u4_n101, u1_u2_u4_n102, u1_u2_u4_n103, u1_u2_u4_n104, u1_u2_u4_n105, u1_u2_u4_n106, u1_u2_u4_n107, 
       u1_u2_u4_n108, u1_u2_u4_n109, u1_u2_u4_n110, u1_u2_u4_n111, u1_u2_u4_n112, u1_u2_u4_n113, u1_u2_u4_n114, u1_u2_u4_n115, u1_u2_u4_n116, 
       u1_u2_u4_n117, u1_u2_u4_n118, u1_u2_u4_n119, u1_u2_u4_n120, u1_u2_u4_n121, u1_u2_u4_n122, u1_u2_u4_n123, u1_u2_u4_n124, u1_u2_u4_n125, 
       u1_u2_u4_n126, u1_u2_u4_n127, u1_u2_u4_n128, u1_u2_u4_n129, u1_u2_u4_n130, u1_u2_u4_n131, u1_u2_u4_n132, u1_u2_u4_n133, u1_u2_u4_n134, 
       u1_u2_u4_n135, u1_u2_u4_n136, u1_u2_u4_n137, u1_u2_u4_n138, u1_u2_u4_n139, u1_u2_u4_n140, u1_u2_u4_n141, u1_u2_u4_n142, u1_u2_u4_n143, 
       u1_u2_u4_n144, u1_u2_u4_n145, u1_u2_u4_n146, u1_u2_u4_n147, u1_u2_u4_n148, u1_u2_u4_n149, u1_u2_u4_n150, u1_u2_u4_n151, u1_u2_u4_n152, 
       u1_u2_u4_n153, u1_u2_u4_n154, u1_u2_u4_n155, u1_u2_u4_n156, u1_u2_u4_n157, u1_u2_u4_n158, u1_u2_u4_n159, u1_u2_u4_n160, u1_u2_u4_n161, 
       u1_u2_u4_n162, u1_u2_u4_n163, u1_u2_u4_n164, u1_u2_u4_n165, u1_u2_u4_n166, u1_u2_u4_n167, u1_u2_u4_n168, u1_u2_u4_n169, u1_u2_u4_n170, 
       u1_u2_u4_n171, u1_u2_u4_n172, u1_u2_u4_n173, u1_u2_u4_n174, u1_u2_u4_n175, u1_u2_u4_n176, u1_u2_u4_n177, u1_u2_u4_n178, u1_u2_u4_n179, 
       u1_u2_u4_n180, u1_u2_u4_n181, u1_u2_u4_n182, u1_u2_u4_n183, u1_u2_u4_n184, u1_u2_u4_n185, u1_u2_u4_n186, u1_u2_u4_n94, u1_u2_u4_n95, 
       u1_u2_u4_n96, u1_u2_u4_n97, u1_u2_u4_n98, u1_u2_u4_n99, u1_u3_X_15, u1_u3_X_16, u1_u3_X_27, u1_u3_X_28, u1_u3_X_29, 
       u1_u3_X_30, u1_u3_X_31, u1_u3_X_32, u1_u3_X_33, u1_u3_X_34, u1_u3_X_45, u1_u3_X_46, u1_u3_u2_n100, u1_u3_u2_n101, 
       u1_u3_u2_n102, u1_u3_u2_n103, u1_u3_u2_n104, u1_u3_u2_n105, u1_u3_u2_n106, u1_u3_u2_n107, u1_u3_u2_n108, u1_u3_u2_n109, u1_u3_u2_n110, 
       u1_u3_u2_n111, u1_u3_u2_n112, u1_u3_u2_n113, u1_u3_u2_n114, u1_u3_u2_n115, u1_u3_u2_n116, u1_u3_u2_n117, u1_u3_u2_n118, u1_u3_u2_n119, 
       u1_u3_u2_n120, u1_u3_u2_n121, u1_u3_u2_n122, u1_u3_u2_n123, u1_u3_u2_n124, u1_u3_u2_n125, u1_u3_u2_n126, u1_u3_u2_n127, u1_u3_u2_n128, 
       u1_u3_u2_n129, u1_u3_u2_n130, u1_u3_u2_n131, u1_u3_u2_n132, u1_u3_u2_n133, u1_u3_u2_n134, u1_u3_u2_n135, u1_u3_u2_n136, u1_u3_u2_n137, 
       u1_u3_u2_n138, u1_u3_u2_n139, u1_u3_u2_n140, u1_u3_u2_n141, u1_u3_u2_n142, u1_u3_u2_n143, u1_u3_u2_n144, u1_u3_u2_n145, u1_u3_u2_n146, 
       u1_u3_u2_n147, u1_u3_u2_n148, u1_u3_u2_n149, u1_u3_u2_n150, u1_u3_u2_n151, u1_u3_u2_n152, u1_u3_u2_n153, u1_u3_u2_n154, u1_u3_u2_n155, 
       u1_u3_u2_n156, u1_u3_u2_n157, u1_u3_u2_n158, u1_u3_u2_n159, u1_u3_u2_n160, u1_u3_u2_n161, u1_u3_u2_n162, u1_u3_u2_n163, u1_u3_u2_n164, 
       u1_u3_u2_n165, u1_u3_u2_n166, u1_u3_u2_n167, u1_u3_u2_n168, u1_u3_u2_n169, u1_u3_u2_n170, u1_u3_u2_n171, u1_u3_u2_n172, u1_u3_u2_n173, 
       u1_u3_u2_n174, u1_u3_u2_n175, u1_u3_u2_n176, u1_u3_u2_n177, u1_u3_u2_n178, u1_u3_u2_n179, u1_u3_u2_n180, u1_u3_u2_n181, u1_u3_u2_n182, 
       u1_u3_u2_n183, u1_u3_u2_n184, u1_u3_u2_n185, u1_u3_u2_n186, u1_u3_u2_n187, u1_u3_u2_n188, u1_u3_u2_n95, u1_u3_u2_n96, u1_u3_u2_n97, 
       u1_u3_u2_n98, u1_u3_u2_n99, u1_u3_u4_n100, u1_u3_u4_n101, u1_u3_u4_n102, u1_u3_u4_n103, u1_u3_u4_n104, u1_u3_u4_n105, u1_u3_u4_n106, 
       u1_u3_u4_n107, u1_u3_u4_n108, u1_u3_u4_n109, u1_u3_u4_n110, u1_u3_u4_n111, u1_u3_u4_n112, u1_u3_u4_n113, u1_u3_u4_n114, u1_u3_u4_n115, 
       u1_u3_u4_n116, u1_u3_u4_n117, u1_u3_u4_n118, u1_u3_u4_n119, u1_u3_u4_n120, u1_u3_u4_n121, u1_u3_u4_n122, u1_u3_u4_n123, u1_u3_u4_n124, 
       u1_u3_u4_n125, u1_u3_u4_n126, u1_u3_u4_n127, u1_u3_u4_n128, u1_u3_u4_n129, u1_u3_u4_n130, u1_u3_u4_n131, u1_u3_u4_n132, u1_u3_u4_n133, 
       u1_u3_u4_n134, u1_u3_u4_n135, u1_u3_u4_n136, u1_u3_u4_n137, u1_u3_u4_n138, u1_u3_u4_n139, u1_u3_u4_n140, u1_u3_u4_n141, u1_u3_u4_n142, 
       u1_u3_u4_n143, u1_u3_u4_n144, u1_u3_u4_n145, u1_u3_u4_n146, u1_u3_u4_n147, u1_u3_u4_n148, u1_u3_u4_n149, u1_u3_u4_n150, u1_u3_u4_n151, 
       u1_u3_u4_n152, u1_u3_u4_n153, u1_u3_u4_n154, u1_u3_u4_n155, u1_u3_u4_n156, u1_u3_u4_n157, u1_u3_u4_n158, u1_u3_u4_n159, u1_u3_u4_n160, 
       u1_u3_u4_n161, u1_u3_u4_n162, u1_u3_u4_n163, u1_u3_u4_n164, u1_u3_u4_n165, u1_u3_u4_n166, u1_u3_u4_n167, u1_u3_u4_n168, u1_u3_u4_n169, 
       u1_u3_u4_n170, u1_u3_u4_n171, u1_u3_u4_n172, u1_u3_u4_n173, u1_u3_u4_n174, u1_u3_u4_n175, u1_u3_u4_n176, u1_u3_u4_n177, u1_u3_u4_n178, 
       u1_u3_u4_n179, u1_u3_u4_n180, u1_u3_u4_n181, u1_u3_u4_n182, u1_u3_u4_n183, u1_u3_u4_n184, u1_u3_u4_n185, u1_u3_u4_n186, u1_u3_u4_n94, 
       u1_u3_u4_n95, u1_u3_u4_n96, u1_u3_u4_n97, u1_u3_u4_n98, u1_u3_u4_n99, u1_u3_u5_n100, u1_u3_u5_n101, u1_u3_u5_n102, u1_u3_u5_n103, 
       u1_u3_u5_n104, u1_u3_u5_n105, u1_u3_u5_n106, u1_u3_u5_n107, u1_u3_u5_n108, u1_u3_u5_n109, u1_u3_u5_n110, u1_u3_u5_n111, u1_u3_u5_n112, 
       u1_u3_u5_n113, u1_u3_u5_n114, u1_u3_u5_n115, u1_u3_u5_n116, u1_u3_u5_n117, u1_u3_u5_n118, u1_u3_u5_n119, u1_u3_u5_n120, u1_u3_u5_n121, 
       u1_u3_u5_n122, u1_u3_u5_n123, u1_u3_u5_n124, u1_u3_u5_n125, u1_u3_u5_n126, u1_u3_u5_n127, u1_u3_u5_n128, u1_u3_u5_n129, u1_u3_u5_n130, 
       u1_u3_u5_n131, u1_u3_u5_n132, u1_u3_u5_n133, u1_u3_u5_n134, u1_u3_u5_n135, u1_u3_u5_n136, u1_u3_u5_n137, u1_u3_u5_n138, u1_u3_u5_n139, 
       u1_u3_u5_n140, u1_u3_u5_n141, u1_u3_u5_n142, u1_u3_u5_n143, u1_u3_u5_n144, u1_u3_u5_n145, u1_u3_u5_n146, u1_u3_u5_n147, u1_u3_u5_n148, 
       u1_u3_u5_n149, u1_u3_u5_n150, u1_u3_u5_n151, u1_u3_u5_n152, u1_u3_u5_n153, u1_u3_u5_n154, u1_u3_u5_n155, u1_u3_u5_n156, u1_u3_u5_n157, 
       u1_u3_u5_n158, u1_u3_u5_n159, u1_u3_u5_n160, u1_u3_u5_n161, u1_u3_u5_n162, u1_u3_u5_n163, u1_u3_u5_n164, u1_u3_u5_n165, u1_u3_u5_n166, 
       u1_u3_u5_n167, u1_u3_u5_n168, u1_u3_u5_n169, u1_u3_u5_n170, u1_u3_u5_n171, u1_u3_u5_n172, u1_u3_u5_n173, u1_u3_u5_n174, u1_u3_u5_n175, 
       u1_u3_u5_n176, u1_u3_u5_n177, u1_u3_u5_n178, u1_u3_u5_n179, u1_u3_u5_n180, u1_u3_u5_n181, u1_u3_u5_n182, u1_u3_u5_n183, u1_u3_u5_n184, 
       u1_u3_u5_n185, u1_u3_u5_n186, u1_u3_u5_n187, u1_u3_u5_n188, u1_u3_u5_n189, u1_u3_u5_n190, u1_u3_u5_n191, u1_u3_u5_n192, u1_u3_u5_n193, 
       u1_u3_u5_n194, u1_u3_u5_n195, u1_u3_u5_n196, u1_u3_u5_n99, u1_u3_u7_n100, u1_u3_u7_n101, u1_u3_u7_n102, u1_u3_u7_n103, u1_u3_u7_n104, 
       u1_u3_u7_n105, u1_u3_u7_n106, u1_u3_u7_n107, u1_u3_u7_n108, u1_u3_u7_n109, u1_u3_u7_n110, u1_u3_u7_n111, u1_u3_u7_n112, u1_u3_u7_n113, 
       u1_u3_u7_n114, u1_u3_u7_n115, u1_u3_u7_n116, u1_u3_u7_n117, u1_u3_u7_n118, u1_u3_u7_n119, u1_u3_u7_n120, u1_u3_u7_n121, u1_u3_u7_n122, 
       u1_u3_u7_n123, u1_u3_u7_n124, u1_u3_u7_n125, u1_u3_u7_n126, u1_u3_u7_n127, u1_u3_u7_n128, u1_u3_u7_n129, u1_u3_u7_n130, u1_u3_u7_n131, 
       u1_u3_u7_n132, u1_u3_u7_n133, u1_u3_u7_n134, u1_u3_u7_n135, u1_u3_u7_n136, u1_u3_u7_n137, u1_u3_u7_n138, u1_u3_u7_n139, u1_u3_u7_n140, 
       u1_u3_u7_n141, u1_u3_u7_n142, u1_u3_u7_n143, u1_u3_u7_n144, u1_u3_u7_n145, u1_u3_u7_n146, u1_u3_u7_n147, u1_u3_u7_n148, u1_u3_u7_n149, 
       u1_u3_u7_n150, u1_u3_u7_n151, u1_u3_u7_n152, u1_u3_u7_n153, u1_u3_u7_n154, u1_u3_u7_n155, u1_u3_u7_n156, u1_u3_u7_n157, u1_u3_u7_n158, 
       u1_u3_u7_n159, u1_u3_u7_n160, u1_u3_u7_n161, u1_u3_u7_n162, u1_u3_u7_n163, u1_u3_u7_n164, u1_u3_u7_n165, u1_u3_u7_n166, u1_u3_u7_n167, 
       u1_u3_u7_n168, u1_u3_u7_n169, u1_u3_u7_n170, u1_u3_u7_n171, u1_u3_u7_n172, u1_u3_u7_n173, u1_u3_u7_n174, u1_u3_u7_n175, u1_u3_u7_n176, 
       u1_u3_u7_n177, u1_u3_u7_n178, u1_u3_u7_n179, u1_u3_u7_n180, u1_u3_u7_n91, u1_u3_u7_n92, u1_u3_u7_n93, u1_u3_u7_n94, u1_u3_u7_n95, 
       u1_u3_u7_n96, u1_u3_u7_n97, u1_u3_u7_n98, u1_u3_u7_n99, u1_u5_X_10, u1_u5_X_9, u1_u5_u1_n100, u1_u5_u1_n101, u1_u5_u1_n102, 
       u1_u5_u1_n103, u1_u5_u1_n104, u1_u5_u1_n105, u1_u5_u1_n106, u1_u5_u1_n107, u1_u5_u1_n108, u1_u5_u1_n109, u1_u5_u1_n110, u1_u5_u1_n111, 
       u1_u5_u1_n112, u1_u5_u1_n113, u1_u5_u1_n114, u1_u5_u1_n115, u1_u5_u1_n116, u1_u5_u1_n117, u1_u5_u1_n118, u1_u5_u1_n119, u1_u5_u1_n120, 
       u1_u5_u1_n121, u1_u5_u1_n122, u1_u5_u1_n123, u1_u5_u1_n124, u1_u5_u1_n125, u1_u5_u1_n126, u1_u5_u1_n127, u1_u5_u1_n128, u1_u5_u1_n129, 
       u1_u5_u1_n130, u1_u5_u1_n131, u1_u5_u1_n132, u1_u5_u1_n133, u1_u5_u1_n134, u1_u5_u1_n135, u1_u5_u1_n136, u1_u5_u1_n137, u1_u5_u1_n138, 
       u1_u5_u1_n139, u1_u5_u1_n140, u1_u5_u1_n141, u1_u5_u1_n142, u1_u5_u1_n143, u1_u5_u1_n144, u1_u5_u1_n145, u1_u5_u1_n146, u1_u5_u1_n147, 
       u1_u5_u1_n148, u1_u5_u1_n149, u1_u5_u1_n150, u1_u5_u1_n151, u1_u5_u1_n152, u1_u5_u1_n153, u1_u5_u1_n154, u1_u5_u1_n155, u1_u5_u1_n156, 
       u1_u5_u1_n157, u1_u5_u1_n158, u1_u5_u1_n159, u1_u5_u1_n160, u1_u5_u1_n161, u1_u5_u1_n162, u1_u5_u1_n163, u1_u5_u1_n164, u1_u5_u1_n165, 
       u1_u5_u1_n166, u1_u5_u1_n167, u1_u5_u1_n168, u1_u5_u1_n169, u1_u5_u1_n170, u1_u5_u1_n171, u1_u5_u1_n172, u1_u5_u1_n173, u1_u5_u1_n174, 
       u1_u5_u1_n175, u1_u5_u1_n176, u1_u5_u1_n177, u1_u5_u1_n178, u1_u5_u1_n179, u1_u5_u1_n180, u1_u5_u1_n181, u1_u5_u1_n182, u1_u5_u1_n183, 
       u1_u5_u1_n184, u1_u5_u1_n185, u1_u5_u1_n186, u1_u5_u1_n187, u1_u5_u1_n188, u1_u5_u1_n95, u1_u5_u1_n96, u1_u5_u1_n97, u1_u5_u1_n98, 
       u1_u5_u1_n99, u1_u7_X_33, u1_u7_X_34, u1_u7_u5_n100, u1_u7_u5_n101, u1_u7_u5_n102, u1_u7_u5_n103, u1_u7_u5_n104, u1_u7_u5_n105, 
       u1_u7_u5_n106, u1_u7_u5_n107, u1_u7_u5_n108, u1_u7_u5_n109, u1_u7_u5_n110, u1_u7_u5_n111, u1_u7_u5_n112, u1_u7_u5_n113, u1_u7_u5_n114, 
       u1_u7_u5_n115, u1_u7_u5_n116, u1_u7_u5_n117, u1_u7_u5_n118, u1_u7_u5_n119, u1_u7_u5_n120, u1_u7_u5_n121, u1_u7_u5_n122, u1_u7_u5_n123, 
       u1_u7_u5_n124, u1_u7_u5_n125, u1_u7_u5_n126, u1_u7_u5_n127, u1_u7_u5_n128, u1_u7_u5_n129, u1_u7_u5_n130, u1_u7_u5_n131, u1_u7_u5_n132, 
       u1_u7_u5_n133, u1_u7_u5_n134, u1_u7_u5_n135, u1_u7_u5_n136, u1_u7_u5_n137, u1_u7_u5_n138, u1_u7_u5_n139, u1_u7_u5_n140, u1_u7_u5_n141, 
       u1_u7_u5_n142, u1_u7_u5_n143, u1_u7_u5_n144, u1_u7_u5_n145, u1_u7_u5_n146, u1_u7_u5_n147, u1_u7_u5_n148, u1_u7_u5_n149, u1_u7_u5_n150, 
       u1_u7_u5_n151, u1_u7_u5_n152, u1_u7_u5_n153, u1_u7_u5_n154, u1_u7_u5_n155, u1_u7_u5_n156, u1_u7_u5_n157, u1_u7_u5_n158, u1_u7_u5_n159, 
       u1_u7_u5_n160, u1_u7_u5_n161, u1_u7_u5_n162, u1_u7_u5_n163, u1_u7_u5_n164, u1_u7_u5_n165, u1_u7_u5_n166, u1_u7_u5_n167, u1_u7_u5_n168, 
       u1_u7_u5_n169, u1_u7_u5_n170, u1_u7_u5_n171, u1_u7_u5_n172, u1_u7_u5_n173, u1_u7_u5_n174, u1_u7_u5_n175, u1_u7_u5_n176, u1_u7_u5_n177, 
       u1_u7_u5_n178, u1_u7_u5_n179, u1_u7_u5_n180, u1_u7_u5_n181, u1_u7_u5_n182, u1_u7_u5_n183, u1_u7_u5_n184, u1_u7_u5_n185, u1_u7_u5_n186, 
       u1_u7_u5_n187, u1_u7_u5_n188, u1_u7_u5_n189, u1_u7_u5_n190, u1_u7_u5_n191, u1_u7_u5_n192, u1_u7_u5_n193, u1_u7_u5_n194, u1_u7_u5_n195, 
       u1_u7_u5_n196, u1_u7_u5_n99, u2_K6_17, u2_K6_18, u2_K8_1, u2_K8_2, u2_K8_3, u2_K8_4, u2_K8_6, 
       u2_out5_16, u2_out5_24, u2_out5_30, u2_out5_6, u2_out7_17, u2_out7_23, u2_out7_31, u2_out7_9, u2_u5_X_13, 
       u2_u5_X_14, u2_u5_X_15, u2_u5_X_16, u2_u5_X_17, u2_u5_X_18, u2_u5_u2_n100, u2_u5_u2_n101, u2_u5_u2_n102, u2_u5_u2_n103, 
       u2_u5_u2_n104, u2_u5_u2_n105, u2_u5_u2_n106, u2_u5_u2_n107, u2_u5_u2_n108, u2_u5_u2_n109, u2_u5_u2_n110, u2_u5_u2_n111, u2_u5_u2_n112, 
       u2_u5_u2_n113, u2_u5_u2_n114, u2_u5_u2_n115, u2_u5_u2_n116, u2_u5_u2_n117, u2_u5_u2_n118, u2_u5_u2_n119, u2_u5_u2_n120, u2_u5_u2_n121, 
       u2_u5_u2_n122, u2_u5_u2_n123, u2_u5_u2_n124, u2_u5_u2_n125, u2_u5_u2_n126, u2_u5_u2_n127, u2_u5_u2_n128, u2_u5_u2_n129, u2_u5_u2_n130, 
       u2_u5_u2_n131, u2_u5_u2_n132, u2_u5_u2_n133, u2_u5_u2_n134, u2_u5_u2_n135, u2_u5_u2_n136, u2_u5_u2_n137, u2_u5_u2_n138, u2_u5_u2_n139, 
       u2_u5_u2_n140, u2_u5_u2_n141, u2_u5_u2_n142, u2_u5_u2_n143, u2_u5_u2_n144, u2_u5_u2_n145, u2_u5_u2_n146, u2_u5_u2_n147, u2_u5_u2_n148, 
       u2_u5_u2_n149, u2_u5_u2_n150, u2_u5_u2_n151, u2_u5_u2_n152, u2_u5_u2_n153, u2_u5_u2_n154, u2_u5_u2_n155, u2_u5_u2_n156, u2_u5_u2_n157, 
       u2_u5_u2_n158, u2_u5_u2_n159, u2_u5_u2_n160, u2_u5_u2_n161, u2_u5_u2_n162, u2_u5_u2_n163, u2_u5_u2_n164, u2_u5_u2_n165, u2_u5_u2_n166, 
       u2_u5_u2_n167, u2_u5_u2_n168, u2_u5_u2_n169, u2_u5_u2_n170, u2_u5_u2_n171, u2_u5_u2_n172, u2_u5_u2_n173, u2_u5_u2_n174, u2_u5_u2_n175, 
       u2_u5_u2_n176, u2_u5_u2_n177, u2_u5_u2_n178, u2_u5_u2_n179, u2_u5_u2_n180, u2_u5_u2_n181, u2_u5_u2_n182, u2_u5_u2_n183, u2_u5_u2_n184, 
       u2_u5_u2_n185, u2_u5_u2_n186, u2_u5_u2_n187, u2_u5_u2_n188, u2_u5_u2_n95, u2_u5_u2_n96, u2_u5_u2_n97, u2_u5_u2_n98, u2_u5_u2_n99, 
       u2_u7_X_1, u2_u7_X_2, u2_u7_X_3, u2_u7_X_4, u2_u7_X_5, u2_u7_X_6, u2_u7_u0_n100, u2_u7_u0_n101, u2_u7_u0_n102, 
       u2_u7_u0_n103, u2_u7_u0_n104, u2_u7_u0_n105, u2_u7_u0_n106, u2_u7_u0_n107, u2_u7_u0_n108, u2_u7_u0_n109, u2_u7_u0_n110, u2_u7_u0_n111, 
       u2_u7_u0_n112, u2_u7_u0_n113, u2_u7_u0_n114, u2_u7_u0_n115, u2_u7_u0_n116, u2_u7_u0_n117, u2_u7_u0_n118, u2_u7_u0_n119, u2_u7_u0_n120, 
       u2_u7_u0_n121, u2_u7_u0_n122, u2_u7_u0_n123, u2_u7_u0_n124, u2_u7_u0_n125, u2_u7_u0_n126, u2_u7_u0_n127, u2_u7_u0_n128, u2_u7_u0_n129, 
       u2_u7_u0_n130, u2_u7_u0_n131, u2_u7_u0_n132, u2_u7_u0_n133, u2_u7_u0_n134, u2_u7_u0_n135, u2_u7_u0_n136, u2_u7_u0_n137, u2_u7_u0_n138, 
       u2_u7_u0_n139, u2_u7_u0_n140, u2_u7_u0_n141, u2_u7_u0_n142, u2_u7_u0_n143, u2_u7_u0_n144, u2_u7_u0_n145, u2_u7_u0_n146, u2_u7_u0_n147, 
       u2_u7_u0_n148, u2_u7_u0_n149, u2_u7_u0_n150, u2_u7_u0_n151, u2_u7_u0_n152, u2_u7_u0_n153, u2_u7_u0_n154, u2_u7_u0_n155, u2_u7_u0_n156, 
       u2_u7_u0_n157, u2_u7_u0_n158, u2_u7_u0_n159, u2_u7_u0_n160, u2_u7_u0_n161, u2_u7_u0_n162, u2_u7_u0_n163, u2_u7_u0_n164, u2_u7_u0_n165, 
       u2_u7_u0_n166, u2_u7_u0_n167, u2_u7_u0_n168, u2_u7_u0_n169, u2_u7_u0_n170, u2_u7_u0_n171, u2_u7_u0_n172, u2_u7_u0_n173, u2_u7_u0_n174, 
       u2_u7_u0_n88, u2_u7_u0_n89, u2_u7_u0_n90, u2_u7_u0_n91, u2_u7_u0_n92, u2_u7_u0_n93, u2_u7_u0_n94, u2_u7_u0_n95, u2_u7_u0_n96, 
       u2_u7_u0_n97, u2_u7_u0_n98, u2_u7_u0_n99, u2_uk_n1059, u2_uk_n1060,  u2_uk_n1110;
  XOR2_X1 u0_U10 (.B( u0_L1_29 ) , .Z( u0_N92 ) , .A( u0_out2_29 ) );
  XOR2_X1 u0_U103 (.B( u0_L0_13 ) , .Z( u0_N44 ) , .A( u0_out1_13 ) );
  XOR2_X1 u0_U11 (.B( u0_L1_28 ) , .Z( u0_N91 ) , .A( u0_out2_28 ) );
  XOR2_X1 u0_U114 (.B( u0_L0_12 ) , .Z( u0_N43 ) , .A( u0_out1_12 ) );
  XOR2_X1 u0_U14 (.B( u0_L1_26 ) , .Z( u0_N89 ) , .A( u0_out2_26 ) );
  XOR2_X1 u0_U147 (.B( u0_L0_9 ) , .Z( u0_N40 ) , .A( u0_out1_9 ) );
  XOR2_X1 u0_U16 (.B( u0_L1_24 ) , .Z( u0_N87 ) , .A( u0_out2_24 ) );
  XOR2_X1 u0_U166 (.B( u0_L10_32 ) , .Z( u0_N383 ) , .A( u0_out11_32 ) );
  XOR2_X1 u0_U168 (.B( u0_L10_30 ) , .Z( u0_N381 ) , .A( u0_out11_30 ) );
  XOR2_X1 u0_U17 (.B( u0_L1_23 ) , .Z( u0_N86 ) , .A( u0_out2_23 ) );
  XOR2_X1 u0_U170 (.B( u0_L0_7 ) , .Z( u0_N38 ) , .A( u0_out1_7 ) );
  XOR2_X1 u0_U171 (.B( u0_L10_28 ) , .Z( u0_N379 ) , .A( u0_out11_28 ) );
  XOR2_X1 u0_U175 (.B( u0_L10_24 ) , .Z( u0_N375 ) , .A( u0_out11_24 ) );
  XOR2_X1 u0_U177 (.B( u0_L10_22 ) , .Z( u0_N373 ) , .A( u0_out11_22 ) );
  XOR2_X1 u0_U181 (.B( u0_L0_6 ) , .Z( u0_N37 ) , .A( u0_out1_6 ) );
  XOR2_X1 u0_U182 (.B( u0_L10_18 ) , .Z( u0_N369 ) , .A( u0_out11_18 ) );
  XOR2_X1 u0_U184 (.B( u0_L10_16 ) , .Z( u0_N367 ) , .A( u0_out11_16 ) );
  XOR2_X1 u0_U187 (.B( u0_L10_13 ) , .Z( u0_N364 ) , .A( u0_out11_13 ) );
  XOR2_X1 u0_U188 (.B( u0_L10_12 ) , .Z( u0_N363 ) , .A( u0_out11_12 ) );
  XOR2_X1 u0_U194 (.B( u0_L10_7 ) , .Z( u0_N358 ) , .A( u0_out11_7 ) );
  XOR2_X1 u0_U195 (.B( u0_L10_6 ) , .Z( u0_N357 ) , .A( u0_out11_6 ) );
  XOR2_X1 u0_U199 (.B( u0_L10_2 ) , .Z( u0_N353 ) , .A( u0_out11_2 ) );
  XOR2_X1 u0_U20 (.B( u0_L1_20 ) , .Z( u0_N83 ) , .A( u0_out2_20 ) );
  XOR2_X1 u0_U201 (.B( u0_L9_32 ) , .Z( u0_N351 ) , .A( u0_out10_32 ) );
  XOR2_X1 u0_U202 (.B( u0_L9_31 ) , .Z( u0_N350 ) , .A( u0_out10_31 ) );
  XOR2_X1 u0_U205 (.B( u0_L9_29 ) , .Z( u0_N348 ) , .A( u0_out10_29 ) );
  XOR2_X1 u0_U206 (.B( u0_L9_28 ) , .Z( u0_N347 ) , .A( u0_out10_28 ) );
  XOR2_X1 u0_U21 (.B( u0_L1_19 ) , .Z( u0_N82 ) , .A( u0_out2_19 ) );
  XOR2_X1 u0_U211 (.B( u0_L9_23 ) , .Z( u0_N342 ) , .A( u0_out10_23 ) );
  XOR2_X1 u0_U212 (.B( u0_L9_22 ) , .Z( u0_N341 ) , .A( u0_out10_22 ) );
  XOR2_X1 u0_U216 (.B( u0_L9_19 ) , .Z( u0_N338 ) , .A( u0_out10_19 ) );
  XOR2_X1 u0_U217 (.B( u0_L9_18 ) , .Z( u0_N337 ) , .A( u0_out10_18 ) );
  XOR2_X1 u0_U218 (.B( u0_L9_17 ) , .Z( u0_N336 ) , .A( u0_out10_17 ) );
  XOR2_X1 u0_U22 (.B( u0_L1_18 ) , .Z( u0_N81 ) , .A( u0_out2_18 ) );
  XOR2_X1 u0_U222 (.B( u0_L9_13 ) , .Z( u0_N332 ) , .A( u0_out10_13 ) );
  XOR2_X1 u0_U223 (.B( u0_L9_12 ) , .Z( u0_N331 ) , .A( u0_out10_12 ) );
  XOR2_X1 u0_U224 (.B( u0_L9_11 ) , .Z( u0_N330 ) , .A( u0_out10_11 ) );
  XOR2_X1 u0_U225 (.B( u0_L0_2 ) , .Z( u0_N33 ) , .A( u0_out1_2 ) );
  XOR2_X1 u0_U227 (.B( u0_L9_9 ) , .Z( u0_N328 ) , .A( u0_out10_9 ) );
  XOR2_X1 u0_U229 (.B( u0_L9_7 ) , .Z( u0_N326 ) , .A( u0_out10_7 ) );
  XOR2_X1 u0_U23 (.B( u0_L1_17 ) , .Z( u0_N80 ) , .A( u0_out2_17 ) );
  XOR2_X1 u0_U232 (.B( u0_L9_4 ) , .Z( u0_N323 ) , .A( u0_out10_4 ) );
  XOR2_X1 u0_U234 (.B( u0_L9_2 ) , .Z( u0_N321 ) , .A( u0_out10_2 ) );
  XOR2_X1 u0_U238 (.B( u0_L8_31 ) , .Z( u0_N318 ) , .A( u0_out9_31 ) );
  XOR2_X1 u0_U246 (.B( u0_L8_23 ) , .Z( u0_N310 ) , .A( u0_out9_23 ) );
  XOR2_X1 u0_U25 (.B( u0_L1_16 ) , .Z( u0_N79 ) , .A( u0_out2_16 ) );
  XOR2_X1 u0_U253 (.B( u0_L8_17 ) , .Z( u0_N304 ) , .A( u0_out9_17 ) );
  XOR2_X1 u0_U263 (.B( u0_L8_9 ) , .Z( u0_N296 ) , .A( u0_out9_9 ) );
  XOR2_X1 u0_U28 (.B( u0_L1_13 ) , .Z( u0_N76 ) , .A( u0_out2_13 ) );
  XOR2_X1 u0_U3 (.B( u0_L2_4 ) , .Z( u0_N99 ) , .A( u0_out3_4 ) );
  XOR2_X1 u0_U30 (.B( u0_L1_11 ) , .Z( u0_N74 ) , .A( u0_out2_11 ) );
  XOR2_X1 u0_U31 (.B( u0_L1_10 ) , .Z( u0_N73 ) , .A( u0_out2_10 ) );
  XOR2_X1 u0_U32 (.B( u0_L1_9 ) , .Z( u0_N72 ) , .A( u0_out2_9 ) );
  XOR2_X1 u0_U343 (.B( u0_L5_32 ) , .Z( u0_N223 ) , .A( u0_out6_32 ) );
  XOR2_X1 u0_U344 (.B( u0_L5_31 ) , .Z( u0_N222 ) , .A( u0_out6_31 ) );
  XOR2_X1 u0_U346 (.B( u0_L5_29 ) , .Z( u0_N220 ) , .A( u0_out6_29 ) );
  XOR2_X1 u0_U349 (.B( u0_L5_27 ) , .Z( u0_N218 ) , .A( u0_out6_27 ) );
  XOR2_X1 u0_U353 (.B( u0_L5_23 ) , .Z( u0_N214 ) , .A( u0_out6_23 ) );
  XOR2_X1 u0_U354 (.B( u0_L5_22 ) , .Z( u0_N213 ) , .A( u0_out6_22 ) );
  XOR2_X1 u0_U355 (.B( u0_L5_21 ) , .Z( u0_N212 ) , .A( u0_out6_21 ) );
  XOR2_X1 u0_U357 (.B( u0_L5_19 ) , .Z( u0_N210 ) , .A( u0_out6_19 ) );
  XOR2_X1 u0_U36 (.B( u0_L1_6 ) , .Z( u0_N69 ) , .A( u0_out2_6 ) );
  XOR2_X1 u0_U360 (.B( u0_L5_17 ) , .Z( u0_N208 ) , .A( u0_out6_17 ) );
  XOR2_X1 u0_U362 (.B( u0_L5_15 ) , .Z( u0_N206 ) , .A( u0_out6_15 ) );
  XOR2_X1 u0_U365 (.B( u0_L5_12 ) , .Z( u0_N203 ) , .A( u0_out6_12 ) );
  XOR2_X1 u0_U366 (.B( u0_L5_11 ) , .Z( u0_N202 ) , .A( u0_out6_11 ) );
  XOR2_X1 u0_U368 (.B( u0_L5_9 ) , .Z( u0_N200 ) , .A( u0_out6_9 ) );
  XOR2_X1 u0_U372 (.B( u0_L5_7 ) , .Z( u0_N198 ) , .A( u0_out6_7 ) );
  XOR2_X1 u0_U374 (.B( u0_L5_5 ) , .Z( u0_N196 ) , .A( u0_out6_5 ) );
  XOR2_X1 u0_U375 (.B( u0_L5_4 ) , .Z( u0_N195 ) , .A( u0_out6_4 ) );
  XOR2_X1 u0_U38 (.B( u0_L1_4 ) , .Z( u0_N67 ) , .A( u0_out2_4 ) );
  XOR2_X1 u0_U40 (.B( u0_L1_2 ) , .Z( u0_N65 ) , .A( u0_out2_2 ) );
  XOR2_X1 u0_U41 (.B( u0_L1_1 ) , .Z( u0_N64 ) , .A( u0_out2_1 ) );
  XOR2_X1 u0_U42 (.B( u0_L0_32 ) , .Z( u0_N63 ) , .A( u0_out1_32 ) );
  XOR2_X1 u0_U43 (.B( u0_L0_31 ) , .Z( u0_N62 ) , .A( u0_out1_31 ) );
  XOR2_X1 u0_U44 (.B( u0_L0_30 ) , .Z( u0_N61 ) , .A( u0_out1_30 ) );
  XOR2_X1 u0_U453 (.B( u0_L2_29 ) , .Z( u0_N124 ) , .A( u0_out3_29 ) );
  XOR2_X1 u0_U464 (.B( u0_L2_19 ) , .Z( u0_N114 ) , .A( u0_out3_19 ) );
  XOR2_X1 u0_U47 (.B( u0_L0_28 ) , .Z( u0_N59 ) , .A( u0_out1_28 ) );
  XOR2_X1 u0_U473 (.B( u0_L2_11 ) , .Z( u0_N106 ) , .A( u0_out3_11 ) );
  XOR2_X1 u0_U484 (.Z( u0_FP_8 ) , .B( u0_L14_8 ) , .A( u0_out15_8 ) );
  XOR2_X1 u0_U486 (.Z( u0_FP_6 ) , .B( u0_L14_6 ) , .A( u0_out15_6 ) );
  XOR2_X1 u0_U489 (.Z( u0_FP_3 ) , .B( u0_L14_3 ) , .A( u0_out15_3 ) );
  XOR2_X1 u0_U492 (.Z( u0_FP_30 ) , .B( u0_L14_30 ) , .A( u0_out15_30 ) );
  XOR2_X1 u0_U497 (.Z( u0_FP_26 ) , .B( u0_L14_26 ) , .A( u0_out15_26 ) );
  XOR2_X1 u0_U498 (.Z( u0_FP_25 ) , .B( u0_L14_25 ) , .A( u0_out15_25 ) );
  XOR2_X1 u0_U499 (.Z( u0_FP_24 ) , .B( u0_L14_24 ) , .A( u0_out15_24 ) );
  XOR2_X1 u0_U503 (.Z( u0_FP_20 ) , .B( u0_L14_20 ) , .A( u0_out15_20 ) );
  XOR2_X1 u0_U504 (.Z( u0_FP_1 ) , .B( u0_L14_1 ) , .A( u0_out15_1 ) );
  XOR2_X1 u0_U508 (.Z( u0_FP_16 ) , .B( u0_L14_16 ) , .A( u0_out15_16 ) );
  XOR2_X1 u0_U51 (.B( u0_L0_24 ) , .Z( u0_N55 ) , .A( u0_out1_24 ) );
  XOR2_X1 u0_U510 (.Z( u0_FP_14 ) , .B( u0_L14_14 ) , .A( u0_out15_14 ) );
  XOR2_X1 u0_U514 (.Z( u0_FP_10 ) , .B( u0_L14_10 ) , .A( u0_out15_10 ) );
  XOR2_X1 u0_U52 (.B( u0_L0_23 ) , .Z( u0_N54 ) , .A( u0_out1_23 ) );
  XOR2_X1 u0_U53 (.B( u0_L0_22 ) , .Z( u0_N53 ) , .A( u0_out1_22 ) );
  XOR2_X1 u0_U58 (.B( u0_L0_18 ) , .Z( u0_N49 ) , .A( u0_out1_18 ) );
  XOR2_X1 u0_U59 (.B( u0_L0_17 ) , .Z( u0_N48 ) , .A( u0_out1_17 ) );
  XOR2_X1 u0_U70 (.B( u0_L0_16 ) , .Z( u0_N47 ) , .A( u0_out1_16 ) );
  XOR2_X1 u0_U8 (.B( u0_L1_31 ) , .Z( u0_N94 ) , .A( u0_out2_31 ) );
  XOR2_X1 u0_U9 (.B( u0_L1_30 ) , .Z( u0_N93 ) , .A( u0_out2_30 ) );
  XOR2_X1 u0_u10_U1 (.B( u0_K11_9 ) , .A( u0_R9_6 ) , .Z( u0_u10_X_9 ) );
  XOR2_X1 u0_u10_U13 (.B( u0_K11_42 ) , .A( u0_R9_29 ) , .Z( u0_u10_X_42 ) );
  XOR2_X1 u0_u10_U14 (.B( u0_K11_41 ) , .A( u0_R9_28 ) , .Z( u0_u10_X_41 ) );
  XOR2_X1 u0_u10_U15 (.B( u0_K11_40 ) , .A( u0_R9_27 ) , .Z( u0_u10_X_40 ) );
  XOR2_X1 u0_u10_U16 (.B( u0_K11_3 ) , .A( u0_R9_2 ) , .Z( u0_u10_X_3 ) );
  XOR2_X1 u0_u10_U17 (.B( u0_K11_39 ) , .A( u0_R9_26 ) , .Z( u0_u10_X_39 ) );
  XOR2_X1 u0_u10_U18 (.B( u0_K11_38 ) , .A( u0_R9_25 ) , .Z( u0_u10_X_38 ) );
  XOR2_X1 u0_u10_U19 (.B( u0_K11_37 ) , .A( u0_R9_24 ) , .Z( u0_u10_X_37 ) );
  XOR2_X1 u0_u10_U2 (.B( u0_K11_8 ) , .A( u0_R9_5 ) , .Z( u0_u10_X_8 ) );
  XOR2_X1 u0_u10_U20 (.B( u0_K11_36 ) , .A( u0_R9_25 ) , .Z( u0_u10_X_36 ) );
  XOR2_X1 u0_u10_U21 (.B( u0_K11_35 ) , .A( u0_R9_24 ) , .Z( u0_u10_X_35 ) );
  XOR2_X1 u0_u10_U22 (.B( u0_K11_34 ) , .A( u0_R9_23 ) , .Z( u0_u10_X_34 ) );
  XOR2_X1 u0_u10_U23 (.B( u0_K11_33 ) , .A( u0_R9_22 ) , .Z( u0_u10_X_33 ) );
  XOR2_X1 u0_u10_U24 (.B( u0_K11_32 ) , .A( u0_R9_21 ) , .Z( u0_u10_X_32 ) );
  XOR2_X1 u0_u10_U25 (.B( u0_K11_31 ) , .A( u0_R9_20 ) , .Z( u0_u10_X_31 ) );
  XOR2_X1 u0_u10_U27 (.B( u0_K11_2 ) , .A( u0_R9_1 ) , .Z( u0_u10_X_2 ) );
  XOR2_X1 u0_u10_U3 (.B( u0_K11_7 ) , .A( u0_R9_4 ) , .Z( u0_u10_X_7 ) );
  XOR2_X1 u0_u10_U38 (.B( u0_K11_1 ) , .A( u0_R9_32 ) , .Z( u0_u10_X_1 ) );
  XOR2_X1 u0_u10_U4 (.B( u0_K11_6 ) , .A( u0_R9_5 ) , .Z( u0_u10_X_6 ) );
  XOR2_X1 u0_u10_U46 (.B( u0_K11_12 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_12 ) );
  XOR2_X1 u0_u10_U47 (.B( u0_K11_11 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_11 ) );
  XOR2_X1 u0_u10_U48 (.B( u0_K11_10 ) , .A( u0_R9_7 ) , .Z( u0_u10_X_10 ) );
  XOR2_X1 u0_u10_U5 (.B( u0_K11_5 ) , .A( u0_R9_4 ) , .Z( u0_u10_X_5 ) );
  XOR2_X1 u0_u10_U6 (.B( u0_K11_4 ) , .A( u0_R9_3 ) , .Z( u0_u10_X_4 ) );
  AND3_X1 u0_u10_u0_U10 (.A2( u0_u10_u0_n112 ) , .ZN( u0_u10_u0_n127 ) , .A3( u0_u10_u0_n130 ) , .A1( u0_u10_u0_n148 ) );
  NAND2_X1 u0_u10_u0_U11 (.ZN( u0_u10_u0_n113 ) , .A1( u0_u10_u0_n139 ) , .A2( u0_u10_u0_n149 ) );
  AND2_X1 u0_u10_u0_U12 (.ZN( u0_u10_u0_n107 ) , .A1( u0_u10_u0_n130 ) , .A2( u0_u10_u0_n140 ) );
  AND2_X1 u0_u10_u0_U13 (.A2( u0_u10_u0_n129 ) , .A1( u0_u10_u0_n130 ) , .ZN( u0_u10_u0_n151 ) );
  AND2_X1 u0_u10_u0_U14 (.A1( u0_u10_u0_n108 ) , .A2( u0_u10_u0_n125 ) , .ZN( u0_u10_u0_n145 ) );
  INV_X1 u0_u10_u0_U15 (.A( u0_u10_u0_n143 ) , .ZN( u0_u10_u0_n173 ) );
  NOR2_X1 u0_u10_u0_U16 (.A2( u0_u10_u0_n136 ) , .ZN( u0_u10_u0_n147 ) , .A1( u0_u10_u0_n160 ) );
  NOR2_X1 u0_u10_u0_U17 (.A1( u0_u10_u0_n163 ) , .A2( u0_u10_u0_n164 ) , .ZN( u0_u10_u0_n95 ) );
  AOI21_X1 u0_u10_u0_U18 (.B1( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n132 ) , .A( u0_u10_u0_n165 ) , .B2( u0_u10_u0_n93 ) );
  INV_X1 u0_u10_u0_U19 (.A( u0_u10_u0_n142 ) , .ZN( u0_u10_u0_n165 ) );
  OAI221_X1 u0_u10_u0_U20 (.C1( u0_u10_u0_n121 ) , .ZN( u0_u10_u0_n122 ) , .B2( u0_u10_u0_n127 ) , .A( u0_u10_u0_n143 ) , .B1( u0_u10_u0_n144 ) , .C2( u0_u10_u0_n147 ) );
  OAI22_X1 u0_u10_u0_U21 (.B1( u0_u10_u0_n125 ) , .ZN( u0_u10_u0_n126 ) , .A1( u0_u10_u0_n138 ) , .A2( u0_u10_u0_n146 ) , .B2( u0_u10_u0_n147 ) );
  OAI22_X1 u0_u10_u0_U22 (.B1( u0_u10_u0_n131 ) , .A1( u0_u10_u0_n144 ) , .B2( u0_u10_u0_n147 ) , .A2( u0_u10_u0_n90 ) , .ZN( u0_u10_u0_n91 ) );
  AND3_X1 u0_u10_u0_U23 (.A3( u0_u10_u0_n121 ) , .A2( u0_u10_u0_n125 ) , .A1( u0_u10_u0_n148 ) , .ZN( u0_u10_u0_n90 ) );
  INV_X1 u0_u10_u0_U24 (.A( u0_u10_u0_n136 ) , .ZN( u0_u10_u0_n161 ) );
  NOR2_X1 u0_u10_u0_U25 (.A1( u0_u10_u0_n120 ) , .ZN( u0_u10_u0_n143 ) , .A2( u0_u10_u0_n167 ) );
  OAI221_X1 u0_u10_u0_U26 (.C1( u0_u10_u0_n112 ) , .ZN( u0_u10_u0_n120 ) , .B1( u0_u10_u0_n138 ) , .B2( u0_u10_u0_n141 ) , .C2( u0_u10_u0_n147 ) , .A( u0_u10_u0_n172 ) );
  AOI22_X1 u0_u10_u0_U27 (.B2( u0_u10_u0_n109 ) , .A2( u0_u10_u0_n110 ) , .ZN( u0_u10_u0_n111 ) , .B1( u0_u10_u0_n118 ) , .A1( u0_u10_u0_n160 ) );
  INV_X1 u0_u10_u0_U28 (.A( u0_u10_u0_n118 ) , .ZN( u0_u10_u0_n158 ) );
  AOI21_X1 u0_u10_u0_U29 (.B1( u0_u10_u0_n132 ) , .ZN( u0_u10_u0_n133 ) , .A( u0_u10_u0_n144 ) , .B2( u0_u10_u0_n166 ) );
  INV_X1 u0_u10_u0_U3 (.A( u0_u10_u0_n113 ) , .ZN( u0_u10_u0_n166 ) );
  AOI21_X1 u0_u10_u0_U30 (.ZN( u0_u10_u0_n104 ) , .B1( u0_u10_u0_n107 ) , .B2( u0_u10_u0_n141 ) , .A( u0_u10_u0_n144 ) );
  AOI21_X1 u0_u10_u0_U31 (.B1( u0_u10_u0_n127 ) , .B2( u0_u10_u0_n129 ) , .A( u0_u10_u0_n138 ) , .ZN( u0_u10_u0_n96 ) );
  AOI21_X1 u0_u10_u0_U32 (.ZN( u0_u10_u0_n116 ) , .B2( u0_u10_u0_n142 ) , .A( u0_u10_u0_n144 ) , .B1( u0_u10_u0_n166 ) );
  NAND2_X1 u0_u10_u0_U33 (.A1( u0_u10_u0_n100 ) , .A2( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n125 ) );
  NAND2_X1 u0_u10_u0_U34 (.A2( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n140 ) , .A1( u0_u10_u0_n94 ) );
  NAND2_X1 u0_u10_u0_U35 (.A1( u0_u10_u0_n101 ) , .A2( u0_u10_u0_n102 ) , .ZN( u0_u10_u0_n150 ) );
  INV_X1 u0_u10_u0_U36 (.A( u0_u10_u0_n138 ) , .ZN( u0_u10_u0_n160 ) );
  NAND2_X1 u0_u10_u0_U37 (.ZN( u0_u10_u0_n142 ) , .A1( u0_u10_u0_n94 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U38 (.A1( u0_u10_u0_n102 ) , .ZN( u0_u10_u0_n128 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U39 (.A2( u0_u10_u0_n102 ) , .A1( u0_u10_u0_n103 ) , .ZN( u0_u10_u0_n149 ) );
  AOI21_X1 u0_u10_u0_U4 (.B2( u0_u10_u0_n131 ) , .ZN( u0_u10_u0_n134 ) , .B1( u0_u10_u0_n151 ) , .A( u0_u10_u0_n158 ) );
  NAND2_X1 u0_u10_u0_U40 (.A1( u0_u10_u0_n100 ) , .ZN( u0_u10_u0_n129 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U41 (.A2( u0_u10_u0_n100 ) , .A1( u0_u10_u0_n101 ) , .ZN( u0_u10_u0_n139 ) );
  NAND2_X1 u0_u10_u0_U42 (.A2( u0_u10_u0_n100 ) , .ZN( u0_u10_u0_n131 ) , .A1( u0_u10_u0_n92 ) );
  NAND2_X1 u0_u10_u0_U43 (.ZN( u0_u10_u0_n108 ) , .A1( u0_u10_u0_n92 ) , .A2( u0_u10_u0_n94 ) );
  NAND2_X1 u0_u10_u0_U44 (.ZN( u0_u10_u0_n148 ) , .A1( u0_u10_u0_n93 ) , .A2( u0_u10_u0_n95 ) );
  NAND2_X1 u0_u10_u0_U45 (.A2( u0_u10_u0_n102 ) , .ZN( u0_u10_u0_n114 ) , .A1( u0_u10_u0_n92 ) );
  NAND2_X1 u0_u10_u0_U46 (.A1( u0_u10_u0_n101 ) , .ZN( u0_u10_u0_n130 ) , .A2( u0_u10_u0_n94 ) );
  NAND2_X1 u0_u10_u0_U47 (.A2( u0_u10_u0_n101 ) , .ZN( u0_u10_u0_n121 ) , .A1( u0_u10_u0_n93 ) );
  INV_X1 u0_u10_u0_U48 (.ZN( u0_u10_u0_n172 ) , .A( u0_u10_u0_n88 ) );
  OAI222_X1 u0_u10_u0_U49 (.C1( u0_u10_u0_n108 ) , .A1( u0_u10_u0_n125 ) , .B2( u0_u10_u0_n128 ) , .B1( u0_u10_u0_n144 ) , .A2( u0_u10_u0_n158 ) , .C2( u0_u10_u0_n161 ) , .ZN( u0_u10_u0_n88 ) );
  NOR2_X1 u0_u10_u0_U5 (.A1( u0_u10_u0_n108 ) , .ZN( u0_u10_u0_n123 ) , .A2( u0_u10_u0_n158 ) );
  NAND2_X1 u0_u10_u0_U50 (.ZN( u0_u10_u0_n112 ) , .A2( u0_u10_u0_n92 ) , .A1( u0_u10_u0_n93 ) );
  OR3_X1 u0_u10_u0_U51 (.A3( u0_u10_u0_n152 ) , .A2( u0_u10_u0_n153 ) , .A1( u0_u10_u0_n154 ) , .ZN( u0_u10_u0_n155 ) );
  AOI21_X1 u0_u10_u0_U52 (.A( u0_u10_u0_n144 ) , .B2( u0_u10_u0_n145 ) , .B1( u0_u10_u0_n146 ) , .ZN( u0_u10_u0_n154 ) );
  AOI21_X1 u0_u10_u0_U53 (.B2( u0_u10_u0_n150 ) , .B1( u0_u10_u0_n151 ) , .ZN( u0_u10_u0_n152 ) , .A( u0_u10_u0_n158 ) );
  AOI21_X1 u0_u10_u0_U54 (.A( u0_u10_u0_n147 ) , .B2( u0_u10_u0_n148 ) , .B1( u0_u10_u0_n149 ) , .ZN( u0_u10_u0_n153 ) );
  INV_X1 u0_u10_u0_U55 (.ZN( u0_u10_u0_n171 ) , .A( u0_u10_u0_n99 ) );
  OAI211_X1 u0_u10_u0_U56 (.C2( u0_u10_u0_n140 ) , .C1( u0_u10_u0_n161 ) , .A( u0_u10_u0_n169 ) , .B( u0_u10_u0_n98 ) , .ZN( u0_u10_u0_n99 ) );
  INV_X1 u0_u10_u0_U57 (.ZN( u0_u10_u0_n169 ) , .A( u0_u10_u0_n91 ) );
  AOI211_X1 u0_u10_u0_U58 (.C1( u0_u10_u0_n118 ) , .A( u0_u10_u0_n123 ) , .B( u0_u10_u0_n96 ) , .C2( u0_u10_u0_n97 ) , .ZN( u0_u10_u0_n98 ) );
  NOR2_X1 u0_u10_u0_U59 (.A2( u0_u10_X_2 ) , .ZN( u0_u10_u0_n103 ) , .A1( u0_u10_u0_n164 ) );
  OAI21_X1 u0_u10_u0_U6 (.B1( u0_u10_u0_n150 ) , .B2( u0_u10_u0_n158 ) , .A( u0_u10_u0_n172 ) , .ZN( u0_u10_u0_n89 ) );
  NOR2_X1 u0_u10_u0_U60 (.A2( u0_u10_X_3 ) , .A1( u0_u10_X_6 ) , .ZN( u0_u10_u0_n94 ) );
  NOR2_X1 u0_u10_u0_U61 (.A2( u0_u10_X_6 ) , .ZN( u0_u10_u0_n100 ) , .A1( u0_u10_u0_n162 ) );
  NOR2_X1 u0_u10_u0_U62 (.A2( u0_u10_X_1 ) , .A1( u0_u10_X_2 ) , .ZN( u0_u10_u0_n92 ) );
  NOR2_X1 u0_u10_u0_U63 (.A2( u0_u10_X_1 ) , .ZN( u0_u10_u0_n101 ) , .A1( u0_u10_u0_n163 ) );
  NOR2_X1 u0_u10_u0_U64 (.A2( u0_u10_X_4 ) , .A1( u0_u10_X_5 ) , .ZN( u0_u10_u0_n118 ) );
  NAND2_X1 u0_u10_u0_U65 (.A2( u0_u10_X_4 ) , .A1( u0_u10_X_5 ) , .ZN( u0_u10_u0_n144 ) );
  NOR2_X1 u0_u10_u0_U66 (.A2( u0_u10_X_5 ) , .ZN( u0_u10_u0_n136 ) , .A1( u0_u10_u0_n159 ) );
  NAND2_X1 u0_u10_u0_U67 (.A1( u0_u10_X_5 ) , .ZN( u0_u10_u0_n138 ) , .A2( u0_u10_u0_n159 ) );
  AND2_X1 u0_u10_u0_U68 (.A2( u0_u10_X_3 ) , .A1( u0_u10_X_6 ) , .ZN( u0_u10_u0_n102 ) );
  AND2_X1 u0_u10_u0_U69 (.A1( u0_u10_X_6 ) , .A2( u0_u10_u0_n162 ) , .ZN( u0_u10_u0_n93 ) );
  AOI21_X1 u0_u10_u0_U7 (.B1( u0_u10_u0_n114 ) , .ZN( u0_u10_u0_n115 ) , .B2( u0_u10_u0_n129 ) , .A( u0_u10_u0_n161 ) );
  INV_X1 u0_u10_u0_U70 (.A( u0_u10_X_4 ) , .ZN( u0_u10_u0_n159 ) );
  INV_X1 u0_u10_u0_U71 (.A( u0_u10_X_1 ) , .ZN( u0_u10_u0_n164 ) );
  INV_X1 u0_u10_u0_U72 (.A( u0_u10_X_2 ) , .ZN( u0_u10_u0_n163 ) );
  INV_X1 u0_u10_u0_U73 (.A( u0_u10_X_3 ) , .ZN( u0_u10_u0_n162 ) );
  INV_X1 u0_u10_u0_U74 (.A( u0_u10_u0_n126 ) , .ZN( u0_u10_u0_n168 ) );
  AOI211_X1 u0_u10_u0_U75 (.B( u0_u10_u0_n133 ) , .A( u0_u10_u0_n134 ) , .C2( u0_u10_u0_n135 ) , .C1( u0_u10_u0_n136 ) , .ZN( u0_u10_u0_n137 ) );
  INV_X1 u0_u10_u0_U76 (.ZN( u0_u10_u0_n174 ) , .A( u0_u10_u0_n89 ) );
  AOI211_X1 u0_u10_u0_U77 (.B( u0_u10_u0_n104 ) , .A( u0_u10_u0_n105 ) , .ZN( u0_u10_u0_n106 ) , .C2( u0_u10_u0_n113 ) , .C1( u0_u10_u0_n160 ) );
  OR4_X1 u0_u10_u0_U78 (.ZN( u0_out10_31 ) , .A4( u0_u10_u0_n155 ) , .A2( u0_u10_u0_n156 ) , .A1( u0_u10_u0_n157 ) , .A3( u0_u10_u0_n173 ) );
  AOI21_X1 u0_u10_u0_U79 (.A( u0_u10_u0_n138 ) , .B2( u0_u10_u0_n139 ) , .B1( u0_u10_u0_n140 ) , .ZN( u0_u10_u0_n157 ) );
  AND2_X1 u0_u10_u0_U8 (.A1( u0_u10_u0_n114 ) , .A2( u0_u10_u0_n121 ) , .ZN( u0_u10_u0_n146 ) );
  AOI21_X1 u0_u10_u0_U80 (.B2( u0_u10_u0_n141 ) , .B1( u0_u10_u0_n142 ) , .ZN( u0_u10_u0_n156 ) , .A( u0_u10_u0_n161 ) );
  OR4_X1 u0_u10_u0_U81 (.ZN( u0_out10_17 ) , .A4( u0_u10_u0_n122 ) , .A2( u0_u10_u0_n123 ) , .A1( u0_u10_u0_n124 ) , .A3( u0_u10_u0_n170 ) );
  AOI21_X1 u0_u10_u0_U82 (.B2( u0_u10_u0_n107 ) , .ZN( u0_u10_u0_n124 ) , .B1( u0_u10_u0_n128 ) , .A( u0_u10_u0_n161 ) );
  INV_X1 u0_u10_u0_U83 (.A( u0_u10_u0_n111 ) , .ZN( u0_u10_u0_n170 ) );
  AOI211_X1 u0_u10_u0_U84 (.B( u0_u10_u0_n115 ) , .A( u0_u10_u0_n116 ) , .C2( u0_u10_u0_n117 ) , .C1( u0_u10_u0_n118 ) , .ZN( u0_u10_u0_n119 ) );
  INV_X1 u0_u10_u0_U85 (.A( u0_u10_u0_n119 ) , .ZN( u0_u10_u0_n167 ) );
  NAND2_X1 u0_u10_u0_U86 (.ZN( u0_u10_u0_n110 ) , .A2( u0_u10_u0_n132 ) , .A1( u0_u10_u0_n145 ) );
  OAI22_X1 u0_u10_u0_U87 (.ZN( u0_u10_u0_n105 ) , .A2( u0_u10_u0_n132 ) , .B1( u0_u10_u0_n146 ) , .A1( u0_u10_u0_n147 ) , .B2( u0_u10_u0_n161 ) );
  NAND3_X1 u0_u10_u0_U88 (.ZN( u0_out10_23 ) , .A3( u0_u10_u0_n137 ) , .A1( u0_u10_u0_n168 ) , .A2( u0_u10_u0_n171 ) );
  NAND3_X1 u0_u10_u0_U89 (.A3( u0_u10_u0_n127 ) , .A2( u0_u10_u0_n128 ) , .ZN( u0_u10_u0_n135 ) , .A1( u0_u10_u0_n150 ) );
  AND2_X1 u0_u10_u0_U9 (.A1( u0_u10_u0_n131 ) , .ZN( u0_u10_u0_n141 ) , .A2( u0_u10_u0_n150 ) );
  NAND3_X1 u0_u10_u0_U90 (.ZN( u0_u10_u0_n117 ) , .A3( u0_u10_u0_n132 ) , .A2( u0_u10_u0_n139 ) , .A1( u0_u10_u0_n148 ) );
  NAND3_X1 u0_u10_u0_U91 (.ZN( u0_u10_u0_n109 ) , .A2( u0_u10_u0_n114 ) , .A3( u0_u10_u0_n140 ) , .A1( u0_u10_u0_n149 ) );
  NAND3_X1 u0_u10_u0_U92 (.ZN( u0_out10_9 ) , .A3( u0_u10_u0_n106 ) , .A2( u0_u10_u0_n171 ) , .A1( u0_u10_u0_n174 ) );
  NAND3_X1 u0_u10_u0_U93 (.A2( u0_u10_u0_n128 ) , .A1( u0_u10_u0_n132 ) , .A3( u0_u10_u0_n146 ) , .ZN( u0_u10_u0_n97 ) );
  AOI21_X1 u0_u10_u1_U10 (.B2( u0_u10_u1_n155 ) , .B1( u0_u10_u1_n156 ) , .ZN( u0_u10_u1_n157 ) , .A( u0_u10_u1_n174 ) );
  NAND3_X1 u0_u10_u1_U100 (.ZN( u0_u10_u1_n113 ) , .A1( u0_u10_u1_n120 ) , .A3( u0_u10_u1_n133 ) , .A2( u0_u10_u1_n155 ) );
  NAND2_X1 u0_u10_u1_U11 (.ZN( u0_u10_u1_n140 ) , .A2( u0_u10_u1_n150 ) , .A1( u0_u10_u1_n155 ) );
  NAND2_X1 u0_u10_u1_U12 (.A1( u0_u10_u1_n131 ) , .ZN( u0_u10_u1_n147 ) , .A2( u0_u10_u1_n153 ) );
  AOI22_X1 u0_u10_u1_U13 (.B2( u0_u10_u1_n136 ) , .A2( u0_u10_u1_n137 ) , .ZN( u0_u10_u1_n143 ) , .A1( u0_u10_u1_n171 ) , .B1( u0_u10_u1_n173 ) );
  INV_X1 u0_u10_u1_U14 (.A( u0_u10_u1_n147 ) , .ZN( u0_u10_u1_n181 ) );
  INV_X1 u0_u10_u1_U15 (.A( u0_u10_u1_n139 ) , .ZN( u0_u10_u1_n174 ) );
  OR4_X1 u0_u10_u1_U16 (.A4( u0_u10_u1_n106 ) , .A3( u0_u10_u1_n107 ) , .ZN( u0_u10_u1_n108 ) , .A1( u0_u10_u1_n117 ) , .A2( u0_u10_u1_n184 ) );
  AOI21_X1 u0_u10_u1_U17 (.ZN( u0_u10_u1_n106 ) , .A( u0_u10_u1_n112 ) , .B1( u0_u10_u1_n154 ) , .B2( u0_u10_u1_n156 ) );
  AOI21_X1 u0_u10_u1_U18 (.ZN( u0_u10_u1_n107 ) , .B1( u0_u10_u1_n134 ) , .B2( u0_u10_u1_n149 ) , .A( u0_u10_u1_n174 ) );
  INV_X1 u0_u10_u1_U19 (.A( u0_u10_u1_n101 ) , .ZN( u0_u10_u1_n184 ) );
  INV_X1 u0_u10_u1_U20 (.A( u0_u10_u1_n112 ) , .ZN( u0_u10_u1_n171 ) );
  NAND2_X1 u0_u10_u1_U21 (.ZN( u0_u10_u1_n141 ) , .A1( u0_u10_u1_n153 ) , .A2( u0_u10_u1_n156 ) );
  AND2_X1 u0_u10_u1_U22 (.A1( u0_u10_u1_n123 ) , .ZN( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n161 ) );
  NAND2_X1 u0_u10_u1_U23 (.A2( u0_u10_u1_n115 ) , .A1( u0_u10_u1_n116 ) , .ZN( u0_u10_u1_n148 ) );
  NAND2_X1 u0_u10_u1_U24 (.A2( u0_u10_u1_n133 ) , .A1( u0_u10_u1_n135 ) , .ZN( u0_u10_u1_n159 ) );
  NAND2_X1 u0_u10_u1_U25 (.A2( u0_u10_u1_n115 ) , .A1( u0_u10_u1_n120 ) , .ZN( u0_u10_u1_n132 ) );
  INV_X1 u0_u10_u1_U26 (.A( u0_u10_u1_n154 ) , .ZN( u0_u10_u1_n178 ) );
  INV_X1 u0_u10_u1_U27 (.A( u0_u10_u1_n151 ) , .ZN( u0_u10_u1_n183 ) );
  AND2_X1 u0_u10_u1_U28 (.A1( u0_u10_u1_n129 ) , .A2( u0_u10_u1_n133 ) , .ZN( u0_u10_u1_n149 ) );
  INV_X1 u0_u10_u1_U29 (.A( u0_u10_u1_n131 ) , .ZN( u0_u10_u1_n180 ) );
  INV_X1 u0_u10_u1_U3 (.A( u0_u10_u1_n159 ) , .ZN( u0_u10_u1_n182 ) );
  OAI221_X1 u0_u10_u1_U30 (.A( u0_u10_u1_n119 ) , .C2( u0_u10_u1_n129 ) , .ZN( u0_u10_u1_n138 ) , .B2( u0_u10_u1_n152 ) , .C1( u0_u10_u1_n174 ) , .B1( u0_u10_u1_n187 ) );
  INV_X1 u0_u10_u1_U31 (.A( u0_u10_u1_n148 ) , .ZN( u0_u10_u1_n187 ) );
  AOI211_X1 u0_u10_u1_U32 (.B( u0_u10_u1_n117 ) , .A( u0_u10_u1_n118 ) , .ZN( u0_u10_u1_n119 ) , .C2( u0_u10_u1_n146 ) , .C1( u0_u10_u1_n159 ) );
  NOR2_X1 u0_u10_u1_U33 (.A1( u0_u10_u1_n168 ) , .A2( u0_u10_u1_n176 ) , .ZN( u0_u10_u1_n98 ) );
  OAI21_X1 u0_u10_u1_U34 (.B2( u0_u10_u1_n123 ) , .ZN( u0_u10_u1_n145 ) , .B1( u0_u10_u1_n160 ) , .A( u0_u10_u1_n185 ) );
  INV_X1 u0_u10_u1_U35 (.A( u0_u10_u1_n122 ) , .ZN( u0_u10_u1_n185 ) );
  AOI21_X1 u0_u10_u1_U36 (.B2( u0_u10_u1_n120 ) , .B1( u0_u10_u1_n121 ) , .ZN( u0_u10_u1_n122 ) , .A( u0_u10_u1_n128 ) );
  NAND2_X1 u0_u10_u1_U37 (.A1( u0_u10_u1_n128 ) , .ZN( u0_u10_u1_n146 ) , .A2( u0_u10_u1_n160 ) );
  NAND2_X1 u0_u10_u1_U38 (.A2( u0_u10_u1_n112 ) , .ZN( u0_u10_u1_n139 ) , .A1( u0_u10_u1_n152 ) );
  NAND2_X1 u0_u10_u1_U39 (.A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n156 ) , .A2( u0_u10_u1_n99 ) );
  AOI221_X1 u0_u10_u1_U4 (.A( u0_u10_u1_n138 ) , .C2( u0_u10_u1_n139 ) , .C1( u0_u10_u1_n140 ) , .B2( u0_u10_u1_n141 ) , .ZN( u0_u10_u1_n142 ) , .B1( u0_u10_u1_n175 ) );
  AOI221_X1 u0_u10_u1_U40 (.B1( u0_u10_u1_n140 ) , .ZN( u0_u10_u1_n167 ) , .B2( u0_u10_u1_n172 ) , .C2( u0_u10_u1_n175 ) , .C1( u0_u10_u1_n178 ) , .A( u0_u10_u1_n188 ) );
  INV_X1 u0_u10_u1_U41 (.ZN( u0_u10_u1_n188 ) , .A( u0_u10_u1_n97 ) );
  AOI211_X1 u0_u10_u1_U42 (.A( u0_u10_u1_n118 ) , .C1( u0_u10_u1_n132 ) , .C2( u0_u10_u1_n139 ) , .B( u0_u10_u1_n96 ) , .ZN( u0_u10_u1_n97 ) );
  AOI21_X1 u0_u10_u1_U43 (.B2( u0_u10_u1_n121 ) , .B1( u0_u10_u1_n135 ) , .A( u0_u10_u1_n152 ) , .ZN( u0_u10_u1_n96 ) );
  NOR2_X1 u0_u10_u1_U44 (.ZN( u0_u10_u1_n117 ) , .A1( u0_u10_u1_n121 ) , .A2( u0_u10_u1_n160 ) );
  AOI21_X1 u0_u10_u1_U45 (.A( u0_u10_u1_n128 ) , .B2( u0_u10_u1_n129 ) , .ZN( u0_u10_u1_n130 ) , .B1( u0_u10_u1_n150 ) );
  NAND2_X1 u0_u10_u1_U46 (.ZN( u0_u10_u1_n112 ) , .A1( u0_u10_u1_n169 ) , .A2( u0_u10_u1_n170 ) );
  NAND2_X1 u0_u10_u1_U47 (.ZN( u0_u10_u1_n129 ) , .A2( u0_u10_u1_n95 ) , .A1( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U48 (.A1( u0_u10_u1_n102 ) , .ZN( u0_u10_u1_n154 ) , .A2( u0_u10_u1_n99 ) );
  NAND2_X1 u0_u10_u1_U49 (.A2( u0_u10_u1_n100 ) , .ZN( u0_u10_u1_n135 ) , .A1( u0_u10_u1_n99 ) );
  AOI211_X1 u0_u10_u1_U5 (.ZN( u0_u10_u1_n124 ) , .A( u0_u10_u1_n138 ) , .C2( u0_u10_u1_n139 ) , .B( u0_u10_u1_n145 ) , .C1( u0_u10_u1_n147 ) );
  AOI21_X1 u0_u10_u1_U50 (.A( u0_u10_u1_n152 ) , .B2( u0_u10_u1_n153 ) , .B1( u0_u10_u1_n154 ) , .ZN( u0_u10_u1_n158 ) );
  INV_X1 u0_u10_u1_U51 (.A( u0_u10_u1_n160 ) , .ZN( u0_u10_u1_n175 ) );
  NAND2_X1 u0_u10_u1_U52 (.A1( u0_u10_u1_n100 ) , .ZN( u0_u10_u1_n116 ) , .A2( u0_u10_u1_n95 ) );
  NAND2_X1 u0_u10_u1_U53 (.A1( u0_u10_u1_n102 ) , .ZN( u0_u10_u1_n131 ) , .A2( u0_u10_u1_n95 ) );
  NAND2_X1 u0_u10_u1_U54 (.A2( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n121 ) , .A1( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U55 (.A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n153 ) , .A2( u0_u10_u1_n98 ) );
  NAND2_X1 u0_u10_u1_U56 (.A2( u0_u10_u1_n104 ) , .A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n133 ) );
  NAND2_X1 u0_u10_u1_U57 (.ZN( u0_u10_u1_n150 ) , .A2( u0_u10_u1_n98 ) , .A1( u0_u10_u1_n99 ) );
  NAND2_X1 u0_u10_u1_U58 (.A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n155 ) , .A2( u0_u10_u1_n95 ) );
  OAI21_X1 u0_u10_u1_U59 (.ZN( u0_u10_u1_n109 ) , .B1( u0_u10_u1_n129 ) , .B2( u0_u10_u1_n160 ) , .A( u0_u10_u1_n167 ) );
  AOI22_X1 u0_u10_u1_U6 (.B2( u0_u10_u1_n113 ) , .A2( u0_u10_u1_n114 ) , .ZN( u0_u10_u1_n125 ) , .A1( u0_u10_u1_n171 ) , .B1( u0_u10_u1_n173 ) );
  NAND2_X1 u0_u10_u1_U60 (.A2( u0_u10_u1_n100 ) , .A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n120 ) );
  NAND2_X1 u0_u10_u1_U61 (.A1( u0_u10_u1_n102 ) , .A2( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n115 ) );
  NAND2_X1 u0_u10_u1_U62 (.A2( u0_u10_u1_n100 ) , .A1( u0_u10_u1_n104 ) , .ZN( u0_u10_u1_n151 ) );
  NAND2_X1 u0_u10_u1_U63 (.A2( u0_u10_u1_n103 ) , .A1( u0_u10_u1_n105 ) , .ZN( u0_u10_u1_n161 ) );
  INV_X1 u0_u10_u1_U64 (.A( u0_u10_u1_n152 ) , .ZN( u0_u10_u1_n173 ) );
  INV_X1 u0_u10_u1_U65 (.A( u0_u10_u1_n128 ) , .ZN( u0_u10_u1_n172 ) );
  NAND2_X1 u0_u10_u1_U66 (.A2( u0_u10_u1_n102 ) , .A1( u0_u10_u1_n103 ) , .ZN( u0_u10_u1_n123 ) );
  AOI211_X1 u0_u10_u1_U67 (.B( u0_u10_u1_n162 ) , .A( u0_u10_u1_n163 ) , .C2( u0_u10_u1_n164 ) , .ZN( u0_u10_u1_n165 ) , .C1( u0_u10_u1_n171 ) );
  AOI21_X1 u0_u10_u1_U68 (.A( u0_u10_u1_n160 ) , .B2( u0_u10_u1_n161 ) , .ZN( u0_u10_u1_n162 ) , .B1( u0_u10_u1_n182 ) );
  OR2_X1 u0_u10_u1_U69 (.A2( u0_u10_u1_n157 ) , .A1( u0_u10_u1_n158 ) , .ZN( u0_u10_u1_n163 ) );
  NAND2_X1 u0_u10_u1_U7 (.ZN( u0_u10_u1_n114 ) , .A1( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n156 ) );
  NOR2_X1 u0_u10_u1_U70 (.A2( u0_u10_X_7 ) , .A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n95 ) );
  NOR2_X1 u0_u10_u1_U71 (.A1( u0_u10_X_12 ) , .A2( u0_u10_X_9 ) , .ZN( u0_u10_u1_n100 ) );
  NOR2_X1 u0_u10_u1_U72 (.A2( u0_u10_X_8 ) , .A1( u0_u10_u1_n177 ) , .ZN( u0_u10_u1_n99 ) );
  NOR2_X1 u0_u10_u1_U73 (.A2( u0_u10_X_12 ) , .ZN( u0_u10_u1_n102 ) , .A1( u0_u10_u1_n176 ) );
  NOR2_X1 u0_u10_u1_U74 (.A2( u0_u10_X_9 ) , .ZN( u0_u10_u1_n105 ) , .A1( u0_u10_u1_n168 ) );
  NAND2_X1 u0_u10_u1_U75 (.A1( u0_u10_X_10 ) , .ZN( u0_u10_u1_n160 ) , .A2( u0_u10_u1_n169 ) );
  NAND2_X1 u0_u10_u1_U76 (.A2( u0_u10_X_10 ) , .A1( u0_u10_X_11 ) , .ZN( u0_u10_u1_n152 ) );
  NAND2_X1 u0_u10_u1_U77 (.A1( u0_u10_X_11 ) , .ZN( u0_u10_u1_n128 ) , .A2( u0_u10_u1_n170 ) );
  AND2_X1 u0_u10_u1_U78 (.A2( u0_u10_X_7 ) , .A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n104 ) );
  AND2_X1 u0_u10_u1_U79 (.A1( u0_u10_X_8 ) , .ZN( u0_u10_u1_n103 ) , .A2( u0_u10_u1_n177 ) );
  NOR2_X1 u0_u10_u1_U8 (.A1( u0_u10_u1_n112 ) , .A2( u0_u10_u1_n116 ) , .ZN( u0_u10_u1_n118 ) );
  INV_X1 u0_u10_u1_U80 (.A( u0_u10_X_10 ) , .ZN( u0_u10_u1_n170 ) );
  INV_X1 u0_u10_u1_U81 (.A( u0_u10_X_9 ) , .ZN( u0_u10_u1_n176 ) );
  INV_X1 u0_u10_u1_U82 (.A( u0_u10_X_11 ) , .ZN( u0_u10_u1_n169 ) );
  INV_X1 u0_u10_u1_U83 (.A( u0_u10_X_12 ) , .ZN( u0_u10_u1_n168 ) );
  INV_X1 u0_u10_u1_U84 (.A( u0_u10_X_7 ) , .ZN( u0_u10_u1_n177 ) );
  NAND4_X1 u0_u10_u1_U85 (.ZN( u0_out10_28 ) , .A4( u0_u10_u1_n124 ) , .A3( u0_u10_u1_n125 ) , .A2( u0_u10_u1_n126 ) , .A1( u0_u10_u1_n127 ) );
  OAI21_X1 u0_u10_u1_U86 (.ZN( u0_u10_u1_n127 ) , .B2( u0_u10_u1_n139 ) , .B1( u0_u10_u1_n175 ) , .A( u0_u10_u1_n183 ) );
  OAI21_X1 u0_u10_u1_U87 (.ZN( u0_u10_u1_n126 ) , .B2( u0_u10_u1_n140 ) , .A( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n178 ) );
  NAND4_X1 u0_u10_u1_U88 (.ZN( u0_out10_18 ) , .A4( u0_u10_u1_n165 ) , .A3( u0_u10_u1_n166 ) , .A1( u0_u10_u1_n167 ) , .A2( u0_u10_u1_n186 ) );
  AOI22_X1 u0_u10_u1_U89 (.B2( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n147 ) , .A2( u0_u10_u1_n148 ) , .ZN( u0_u10_u1_n166 ) , .A1( u0_u10_u1_n172 ) );
  OAI21_X1 u0_u10_u1_U9 (.ZN( u0_u10_u1_n101 ) , .B1( u0_u10_u1_n141 ) , .A( u0_u10_u1_n146 ) , .B2( u0_u10_u1_n183 ) );
  INV_X1 u0_u10_u1_U90 (.A( u0_u10_u1_n145 ) , .ZN( u0_u10_u1_n186 ) );
  NAND4_X1 u0_u10_u1_U91 (.ZN( u0_out10_2 ) , .A4( u0_u10_u1_n142 ) , .A3( u0_u10_u1_n143 ) , .A2( u0_u10_u1_n144 ) , .A1( u0_u10_u1_n179 ) );
  OAI21_X1 u0_u10_u1_U92 (.B2( u0_u10_u1_n132 ) , .ZN( u0_u10_u1_n144 ) , .A( u0_u10_u1_n146 ) , .B1( u0_u10_u1_n180 ) );
  INV_X1 u0_u10_u1_U93 (.A( u0_u10_u1_n130 ) , .ZN( u0_u10_u1_n179 ) );
  OR4_X1 u0_u10_u1_U94 (.ZN( u0_out10_13 ) , .A4( u0_u10_u1_n108 ) , .A3( u0_u10_u1_n109 ) , .A2( u0_u10_u1_n110 ) , .A1( u0_u10_u1_n111 ) );
  AOI21_X1 u0_u10_u1_U95 (.ZN( u0_u10_u1_n111 ) , .A( u0_u10_u1_n128 ) , .B2( u0_u10_u1_n131 ) , .B1( u0_u10_u1_n135 ) );
  AOI21_X1 u0_u10_u1_U96 (.ZN( u0_u10_u1_n110 ) , .A( u0_u10_u1_n116 ) , .B1( u0_u10_u1_n152 ) , .B2( u0_u10_u1_n160 ) );
  NAND3_X1 u0_u10_u1_U97 (.A3( u0_u10_u1_n149 ) , .A2( u0_u10_u1_n150 ) , .A1( u0_u10_u1_n151 ) , .ZN( u0_u10_u1_n164 ) );
  NAND3_X1 u0_u10_u1_U98 (.A3( u0_u10_u1_n134 ) , .A2( u0_u10_u1_n135 ) , .ZN( u0_u10_u1_n136 ) , .A1( u0_u10_u1_n151 ) );
  NAND3_X1 u0_u10_u1_U99 (.A1( u0_u10_u1_n133 ) , .ZN( u0_u10_u1_n137 ) , .A2( u0_u10_u1_n154 ) , .A3( u0_u10_u1_n181 ) );
  INV_X1 u0_u10_u5_U10 (.A( u0_u10_u5_n121 ) , .ZN( u0_u10_u5_n177 ) );
  NOR3_X1 u0_u10_u5_U100 (.A3( u0_u10_u5_n141 ) , .A1( u0_u10_u5_n142 ) , .ZN( u0_u10_u5_n143 ) , .A2( u0_u10_u5_n191 ) );
  NAND4_X1 u0_u10_u5_U101 (.ZN( u0_out10_4 ) , .A4( u0_u10_u5_n112 ) , .A2( u0_u10_u5_n113 ) , .A1( u0_u10_u5_n114 ) , .A3( u0_u10_u5_n195 ) );
  AOI211_X1 u0_u10_u5_U102 (.A( u0_u10_u5_n110 ) , .C1( u0_u10_u5_n111 ) , .ZN( u0_u10_u5_n112 ) , .B( u0_u10_u5_n118 ) , .C2( u0_u10_u5_n177 ) );
  AOI222_X1 u0_u10_u5_U103 (.ZN( u0_u10_u5_n113 ) , .A1( u0_u10_u5_n131 ) , .C1( u0_u10_u5_n148 ) , .B2( u0_u10_u5_n174 ) , .C2( u0_u10_u5_n178 ) , .A2( u0_u10_u5_n179 ) , .B1( u0_u10_u5_n99 ) );
  NAND3_X1 u0_u10_u5_U104 (.A2( u0_u10_u5_n154 ) , .A3( u0_u10_u5_n158 ) , .A1( u0_u10_u5_n161 ) , .ZN( u0_u10_u5_n99 ) );
  NOR2_X1 u0_u10_u5_U11 (.ZN( u0_u10_u5_n160 ) , .A2( u0_u10_u5_n173 ) , .A1( u0_u10_u5_n177 ) );
  INV_X1 u0_u10_u5_U12 (.A( u0_u10_u5_n150 ) , .ZN( u0_u10_u5_n174 ) );
  AOI21_X1 u0_u10_u5_U13 (.A( u0_u10_u5_n160 ) , .B2( u0_u10_u5_n161 ) , .ZN( u0_u10_u5_n162 ) , .B1( u0_u10_u5_n192 ) );
  INV_X1 u0_u10_u5_U14 (.A( u0_u10_u5_n159 ) , .ZN( u0_u10_u5_n192 ) );
  AOI21_X1 u0_u10_u5_U15 (.A( u0_u10_u5_n156 ) , .B2( u0_u10_u5_n157 ) , .B1( u0_u10_u5_n158 ) , .ZN( u0_u10_u5_n163 ) );
  AOI21_X1 u0_u10_u5_U16 (.B2( u0_u10_u5_n139 ) , .B1( u0_u10_u5_n140 ) , .ZN( u0_u10_u5_n141 ) , .A( u0_u10_u5_n150 ) );
  OAI21_X1 u0_u10_u5_U17 (.A( u0_u10_u5_n133 ) , .B2( u0_u10_u5_n134 ) , .B1( u0_u10_u5_n135 ) , .ZN( u0_u10_u5_n142 ) );
  OAI21_X1 u0_u10_u5_U18 (.ZN( u0_u10_u5_n133 ) , .B2( u0_u10_u5_n147 ) , .A( u0_u10_u5_n173 ) , .B1( u0_u10_u5_n188 ) );
  NAND2_X1 u0_u10_u5_U19 (.A2( u0_u10_u5_n119 ) , .A1( u0_u10_u5_n123 ) , .ZN( u0_u10_u5_n137 ) );
  INV_X1 u0_u10_u5_U20 (.A( u0_u10_u5_n155 ) , .ZN( u0_u10_u5_n194 ) );
  NAND2_X1 u0_u10_u5_U21 (.A1( u0_u10_u5_n121 ) , .ZN( u0_u10_u5_n132 ) , .A2( u0_u10_u5_n172 ) );
  NAND2_X1 u0_u10_u5_U22 (.A2( u0_u10_u5_n122 ) , .ZN( u0_u10_u5_n136 ) , .A1( u0_u10_u5_n154 ) );
  NAND2_X1 u0_u10_u5_U23 (.A2( u0_u10_u5_n119 ) , .A1( u0_u10_u5_n120 ) , .ZN( u0_u10_u5_n159 ) );
  INV_X1 u0_u10_u5_U24 (.A( u0_u10_u5_n156 ) , .ZN( u0_u10_u5_n175 ) );
  INV_X1 u0_u10_u5_U25 (.A( u0_u10_u5_n158 ) , .ZN( u0_u10_u5_n188 ) );
  INV_X1 u0_u10_u5_U26 (.A( u0_u10_u5_n152 ) , .ZN( u0_u10_u5_n179 ) );
  INV_X1 u0_u10_u5_U27 (.A( u0_u10_u5_n140 ) , .ZN( u0_u10_u5_n182 ) );
  INV_X1 u0_u10_u5_U28 (.A( u0_u10_u5_n151 ) , .ZN( u0_u10_u5_n183 ) );
  INV_X1 u0_u10_u5_U29 (.A( u0_u10_u5_n123 ) , .ZN( u0_u10_u5_n185 ) );
  NOR2_X1 u0_u10_u5_U3 (.ZN( u0_u10_u5_n134 ) , .A1( u0_u10_u5_n183 ) , .A2( u0_u10_u5_n190 ) );
  INV_X1 u0_u10_u5_U30 (.A( u0_u10_u5_n161 ) , .ZN( u0_u10_u5_n184 ) );
  INV_X1 u0_u10_u5_U31 (.A( u0_u10_u5_n139 ) , .ZN( u0_u10_u5_n189 ) );
  INV_X1 u0_u10_u5_U32 (.A( u0_u10_u5_n157 ) , .ZN( u0_u10_u5_n190 ) );
  INV_X1 u0_u10_u5_U33 (.A( u0_u10_u5_n120 ) , .ZN( u0_u10_u5_n193 ) );
  NAND2_X1 u0_u10_u5_U34 (.ZN( u0_u10_u5_n111 ) , .A1( u0_u10_u5_n140 ) , .A2( u0_u10_u5_n155 ) );
  NOR2_X1 u0_u10_u5_U35 (.ZN( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n170 ) , .A2( u0_u10_u5_n180 ) );
  INV_X1 u0_u10_u5_U36 (.A( u0_u10_u5_n117 ) , .ZN( u0_u10_u5_n196 ) );
  OAI221_X1 u0_u10_u5_U37 (.A( u0_u10_u5_n116 ) , .ZN( u0_u10_u5_n117 ) , .B2( u0_u10_u5_n119 ) , .C1( u0_u10_u5_n153 ) , .C2( u0_u10_u5_n158 ) , .B1( u0_u10_u5_n172 ) );
  AOI222_X1 u0_u10_u5_U38 (.ZN( u0_u10_u5_n116 ) , .B2( u0_u10_u5_n145 ) , .C1( u0_u10_u5_n148 ) , .A2( u0_u10_u5_n174 ) , .C2( u0_u10_u5_n177 ) , .B1( u0_u10_u5_n187 ) , .A1( u0_u10_u5_n193 ) );
  INV_X1 u0_u10_u5_U39 (.A( u0_u10_u5_n115 ) , .ZN( u0_u10_u5_n187 ) );
  INV_X1 u0_u10_u5_U4 (.A( u0_u10_u5_n138 ) , .ZN( u0_u10_u5_n191 ) );
  AOI22_X1 u0_u10_u5_U40 (.B2( u0_u10_u5_n131 ) , .A2( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n169 ) , .B1( u0_u10_u5_n174 ) , .A1( u0_u10_u5_n185 ) );
  NOR2_X1 u0_u10_u5_U41 (.A1( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n150 ) , .A2( u0_u10_u5_n173 ) );
  AOI21_X1 u0_u10_u5_U42 (.A( u0_u10_u5_n118 ) , .B2( u0_u10_u5_n145 ) , .ZN( u0_u10_u5_n168 ) , .B1( u0_u10_u5_n186 ) );
  INV_X1 u0_u10_u5_U43 (.A( u0_u10_u5_n122 ) , .ZN( u0_u10_u5_n186 ) );
  NOR2_X1 u0_u10_u5_U44 (.A1( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n152 ) , .A2( u0_u10_u5_n176 ) );
  NOR2_X1 u0_u10_u5_U45 (.A1( u0_u10_u5_n115 ) , .ZN( u0_u10_u5_n118 ) , .A2( u0_u10_u5_n153 ) );
  NOR2_X1 u0_u10_u5_U46 (.A2( u0_u10_u5_n145 ) , .ZN( u0_u10_u5_n156 ) , .A1( u0_u10_u5_n174 ) );
  NOR2_X1 u0_u10_u5_U47 (.ZN( u0_u10_u5_n121 ) , .A2( u0_u10_u5_n145 ) , .A1( u0_u10_u5_n176 ) );
  AOI22_X1 u0_u10_u5_U48 (.ZN( u0_u10_u5_n114 ) , .A2( u0_u10_u5_n137 ) , .A1( u0_u10_u5_n145 ) , .B2( u0_u10_u5_n175 ) , .B1( u0_u10_u5_n193 ) );
  OAI211_X1 u0_u10_u5_U49 (.B( u0_u10_u5_n124 ) , .A( u0_u10_u5_n125 ) , .C2( u0_u10_u5_n126 ) , .C1( u0_u10_u5_n127 ) , .ZN( u0_u10_u5_n128 ) );
  OAI21_X1 u0_u10_u5_U5 (.B2( u0_u10_u5_n136 ) , .B1( u0_u10_u5_n137 ) , .ZN( u0_u10_u5_n138 ) , .A( u0_u10_u5_n177 ) );
  NOR3_X1 u0_u10_u5_U50 (.ZN( u0_u10_u5_n127 ) , .A1( u0_u10_u5_n136 ) , .A3( u0_u10_u5_n148 ) , .A2( u0_u10_u5_n182 ) );
  OAI21_X1 u0_u10_u5_U51 (.ZN( u0_u10_u5_n124 ) , .A( u0_u10_u5_n177 ) , .B2( u0_u10_u5_n183 ) , .B1( u0_u10_u5_n189 ) );
  OAI21_X1 u0_u10_u5_U52 (.ZN( u0_u10_u5_n125 ) , .A( u0_u10_u5_n174 ) , .B2( u0_u10_u5_n185 ) , .B1( u0_u10_u5_n190 ) );
  AOI21_X1 u0_u10_u5_U53 (.A( u0_u10_u5_n153 ) , .B2( u0_u10_u5_n154 ) , .B1( u0_u10_u5_n155 ) , .ZN( u0_u10_u5_n164 ) );
  AOI21_X1 u0_u10_u5_U54 (.ZN( u0_u10_u5_n110 ) , .B1( u0_u10_u5_n122 ) , .B2( u0_u10_u5_n139 ) , .A( u0_u10_u5_n153 ) );
  INV_X1 u0_u10_u5_U55 (.A( u0_u10_u5_n153 ) , .ZN( u0_u10_u5_n176 ) );
  INV_X1 u0_u10_u5_U56 (.A( u0_u10_u5_n126 ) , .ZN( u0_u10_u5_n173 ) );
  AND2_X1 u0_u10_u5_U57 (.A2( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n107 ) , .ZN( u0_u10_u5_n147 ) );
  AND2_X1 u0_u10_u5_U58 (.A2( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n108 ) , .ZN( u0_u10_u5_n148 ) );
  NAND2_X1 u0_u10_u5_U59 (.A1( u0_u10_u5_n105 ) , .A2( u0_u10_u5_n106 ) , .ZN( u0_u10_u5_n158 ) );
  INV_X1 u0_u10_u5_U6 (.A( u0_u10_u5_n135 ) , .ZN( u0_u10_u5_n178 ) );
  NAND2_X1 u0_u10_u5_U60 (.A2( u0_u10_u5_n108 ) , .A1( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n139 ) );
  NAND2_X1 u0_u10_u5_U61 (.A1( u0_u10_u5_n106 ) , .A2( u0_u10_u5_n108 ) , .ZN( u0_u10_u5_n119 ) );
  NAND2_X1 u0_u10_u5_U62 (.A2( u0_u10_u5_n103 ) , .A1( u0_u10_u5_n105 ) , .ZN( u0_u10_u5_n140 ) );
  NAND2_X1 u0_u10_u5_U63 (.A2( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n105 ) , .ZN( u0_u10_u5_n155 ) );
  NAND2_X1 u0_u10_u5_U64 (.A2( u0_u10_u5_n106 ) , .A1( u0_u10_u5_n107 ) , .ZN( u0_u10_u5_n122 ) );
  NAND2_X1 u0_u10_u5_U65 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n106 ) , .ZN( u0_u10_u5_n115 ) );
  NAND2_X1 u0_u10_u5_U66 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n103 ) , .ZN( u0_u10_u5_n161 ) );
  NAND2_X1 u0_u10_u5_U67 (.A1( u0_u10_u5_n105 ) , .A2( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n154 ) );
  INV_X1 u0_u10_u5_U68 (.A( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n172 ) );
  NAND2_X1 u0_u10_u5_U69 (.A1( u0_u10_u5_n103 ) , .A2( u0_u10_u5_n108 ) , .ZN( u0_u10_u5_n123 ) );
  OAI22_X1 u0_u10_u5_U7 (.B2( u0_u10_u5_n149 ) , .B1( u0_u10_u5_n150 ) , .A2( u0_u10_u5_n151 ) , .A1( u0_u10_u5_n152 ) , .ZN( u0_u10_u5_n165 ) );
  NAND2_X1 u0_u10_u5_U70 (.A2( u0_u10_u5_n103 ) , .A1( u0_u10_u5_n107 ) , .ZN( u0_u10_u5_n151 ) );
  NAND2_X1 u0_u10_u5_U71 (.A2( u0_u10_u5_n107 ) , .A1( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n120 ) );
  NAND2_X1 u0_u10_u5_U72 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n109 ) , .ZN( u0_u10_u5_n157 ) );
  AND2_X1 u0_u10_u5_U73 (.A2( u0_u10_u5_n100 ) , .A1( u0_u10_u5_n104 ) , .ZN( u0_u10_u5_n131 ) );
  INV_X1 u0_u10_u5_U74 (.A( u0_u10_u5_n102 ) , .ZN( u0_u10_u5_n195 ) );
  OAI221_X1 u0_u10_u5_U75 (.A( u0_u10_u5_n101 ) , .ZN( u0_u10_u5_n102 ) , .C2( u0_u10_u5_n115 ) , .C1( u0_u10_u5_n126 ) , .B1( u0_u10_u5_n134 ) , .B2( u0_u10_u5_n160 ) );
  OAI21_X1 u0_u10_u5_U76 (.ZN( u0_u10_u5_n101 ) , .B1( u0_u10_u5_n137 ) , .A( u0_u10_u5_n146 ) , .B2( u0_u10_u5_n147 ) );
  NOR2_X1 u0_u10_u5_U77 (.A2( u0_u10_X_34 ) , .A1( u0_u10_X_35 ) , .ZN( u0_u10_u5_n145 ) );
  NOR2_X1 u0_u10_u5_U78 (.A2( u0_u10_X_34 ) , .ZN( u0_u10_u5_n146 ) , .A1( u0_u10_u5_n171 ) );
  NOR2_X1 u0_u10_u5_U79 (.A2( u0_u10_X_31 ) , .A1( u0_u10_X_32 ) , .ZN( u0_u10_u5_n103 ) );
  NOR3_X1 u0_u10_u5_U8 (.A2( u0_u10_u5_n147 ) , .A1( u0_u10_u5_n148 ) , .ZN( u0_u10_u5_n149 ) , .A3( u0_u10_u5_n194 ) );
  NOR2_X1 u0_u10_u5_U80 (.A2( u0_u10_X_36 ) , .ZN( u0_u10_u5_n105 ) , .A1( u0_u10_u5_n180 ) );
  NOR2_X1 u0_u10_u5_U81 (.A2( u0_u10_X_33 ) , .ZN( u0_u10_u5_n108 ) , .A1( u0_u10_u5_n170 ) );
  NOR2_X1 u0_u10_u5_U82 (.A2( u0_u10_X_33 ) , .A1( u0_u10_X_36 ) , .ZN( u0_u10_u5_n107 ) );
  NOR2_X1 u0_u10_u5_U83 (.A2( u0_u10_X_31 ) , .ZN( u0_u10_u5_n104 ) , .A1( u0_u10_u5_n181 ) );
  NAND2_X1 u0_u10_u5_U84 (.A2( u0_u10_X_34 ) , .A1( u0_u10_X_35 ) , .ZN( u0_u10_u5_n153 ) );
  NAND2_X1 u0_u10_u5_U85 (.A1( u0_u10_X_34 ) , .ZN( u0_u10_u5_n126 ) , .A2( u0_u10_u5_n171 ) );
  AND2_X1 u0_u10_u5_U86 (.A1( u0_u10_X_31 ) , .A2( u0_u10_X_32 ) , .ZN( u0_u10_u5_n106 ) );
  AND2_X1 u0_u10_u5_U87 (.A1( u0_u10_X_31 ) , .ZN( u0_u10_u5_n109 ) , .A2( u0_u10_u5_n181 ) );
  INV_X1 u0_u10_u5_U88 (.A( u0_u10_X_33 ) , .ZN( u0_u10_u5_n180 ) );
  INV_X1 u0_u10_u5_U89 (.A( u0_u10_X_35 ) , .ZN( u0_u10_u5_n171 ) );
  NOR2_X1 u0_u10_u5_U9 (.ZN( u0_u10_u5_n135 ) , .A1( u0_u10_u5_n173 ) , .A2( u0_u10_u5_n176 ) );
  INV_X1 u0_u10_u5_U90 (.A( u0_u10_X_36 ) , .ZN( u0_u10_u5_n170 ) );
  INV_X1 u0_u10_u5_U91 (.A( u0_u10_X_32 ) , .ZN( u0_u10_u5_n181 ) );
  NAND4_X1 u0_u10_u5_U92 (.ZN( u0_out10_29 ) , .A4( u0_u10_u5_n129 ) , .A3( u0_u10_u5_n130 ) , .A2( u0_u10_u5_n168 ) , .A1( u0_u10_u5_n196 ) );
  AOI221_X1 u0_u10_u5_U93 (.A( u0_u10_u5_n128 ) , .ZN( u0_u10_u5_n129 ) , .C2( u0_u10_u5_n132 ) , .B2( u0_u10_u5_n159 ) , .B1( u0_u10_u5_n176 ) , .C1( u0_u10_u5_n184 ) );
  AOI222_X1 u0_u10_u5_U94 (.ZN( u0_u10_u5_n130 ) , .A2( u0_u10_u5_n146 ) , .B1( u0_u10_u5_n147 ) , .C2( u0_u10_u5_n175 ) , .B2( u0_u10_u5_n179 ) , .A1( u0_u10_u5_n188 ) , .C1( u0_u10_u5_n194 ) );
  NAND4_X1 u0_u10_u5_U95 (.ZN( u0_out10_19 ) , .A4( u0_u10_u5_n166 ) , .A3( u0_u10_u5_n167 ) , .A2( u0_u10_u5_n168 ) , .A1( u0_u10_u5_n169 ) );
  AOI22_X1 u0_u10_u5_U96 (.B2( u0_u10_u5_n145 ) , .A2( u0_u10_u5_n146 ) , .ZN( u0_u10_u5_n167 ) , .B1( u0_u10_u5_n182 ) , .A1( u0_u10_u5_n189 ) );
  NOR4_X1 u0_u10_u5_U97 (.A4( u0_u10_u5_n162 ) , .A3( u0_u10_u5_n163 ) , .A2( u0_u10_u5_n164 ) , .A1( u0_u10_u5_n165 ) , .ZN( u0_u10_u5_n166 ) );
  NAND4_X1 u0_u10_u5_U98 (.ZN( u0_out10_11 ) , .A4( u0_u10_u5_n143 ) , .A3( u0_u10_u5_n144 ) , .A2( u0_u10_u5_n169 ) , .A1( u0_u10_u5_n196 ) );
  AOI22_X1 u0_u10_u5_U99 (.A2( u0_u10_u5_n132 ) , .ZN( u0_u10_u5_n144 ) , .B2( u0_u10_u5_n145 ) , .B1( u0_u10_u5_n184 ) , .A1( u0_u10_u5_n194 ) );
  AOI22_X1 u0_u10_u6_U10 (.A2( u0_u10_u6_n151 ) , .B2( u0_u10_u6_n161 ) , .A1( u0_u10_u6_n167 ) , .B1( u0_u10_u6_n170 ) , .ZN( u0_u10_u6_n89 ) );
  AOI21_X1 u0_u10_u6_U11 (.B1( u0_u10_u6_n107 ) , .B2( u0_u10_u6_n132 ) , .A( u0_u10_u6_n158 ) , .ZN( u0_u10_u6_n88 ) );
  AOI21_X1 u0_u10_u6_U12 (.B2( u0_u10_u6_n147 ) , .B1( u0_u10_u6_n148 ) , .ZN( u0_u10_u6_n149 ) , .A( u0_u10_u6_n158 ) );
  AOI21_X1 u0_u10_u6_U13 (.ZN( u0_u10_u6_n106 ) , .A( u0_u10_u6_n142 ) , .B2( u0_u10_u6_n159 ) , .B1( u0_u10_u6_n164 ) );
  INV_X1 u0_u10_u6_U14 (.A( u0_u10_u6_n155 ) , .ZN( u0_u10_u6_n161 ) );
  INV_X1 u0_u10_u6_U15 (.A( u0_u10_u6_n128 ) , .ZN( u0_u10_u6_n164 ) );
  NAND2_X1 u0_u10_u6_U16 (.ZN( u0_u10_u6_n110 ) , .A1( u0_u10_u6_n122 ) , .A2( u0_u10_u6_n129 ) );
  NAND2_X1 u0_u10_u6_U17 (.ZN( u0_u10_u6_n124 ) , .A2( u0_u10_u6_n146 ) , .A1( u0_u10_u6_n148 ) );
  INV_X1 u0_u10_u6_U18 (.A( u0_u10_u6_n132 ) , .ZN( u0_u10_u6_n171 ) );
  AND2_X1 u0_u10_u6_U19 (.A1( u0_u10_u6_n100 ) , .ZN( u0_u10_u6_n130 ) , .A2( u0_u10_u6_n147 ) );
  INV_X1 u0_u10_u6_U20 (.A( u0_u10_u6_n127 ) , .ZN( u0_u10_u6_n173 ) );
  INV_X1 u0_u10_u6_U21 (.A( u0_u10_u6_n121 ) , .ZN( u0_u10_u6_n167 ) );
  INV_X1 u0_u10_u6_U22 (.A( u0_u10_u6_n100 ) , .ZN( u0_u10_u6_n169 ) );
  INV_X1 u0_u10_u6_U23 (.A( u0_u10_u6_n123 ) , .ZN( u0_u10_u6_n170 ) );
  INV_X1 u0_u10_u6_U24 (.A( u0_u10_u6_n113 ) , .ZN( u0_u10_u6_n168 ) );
  AND2_X1 u0_u10_u6_U25 (.A1( u0_u10_u6_n107 ) , .A2( u0_u10_u6_n119 ) , .ZN( u0_u10_u6_n133 ) );
  AND2_X1 u0_u10_u6_U26 (.A2( u0_u10_u6_n121 ) , .A1( u0_u10_u6_n122 ) , .ZN( u0_u10_u6_n131 ) );
  AND3_X1 u0_u10_u6_U27 (.ZN( u0_u10_u6_n120 ) , .A2( u0_u10_u6_n127 ) , .A1( u0_u10_u6_n132 ) , .A3( u0_u10_u6_n145 ) );
  INV_X1 u0_u10_u6_U28 (.A( u0_u10_u6_n146 ) , .ZN( u0_u10_u6_n163 ) );
  AOI222_X1 u0_u10_u6_U29 (.ZN( u0_u10_u6_n114 ) , .A1( u0_u10_u6_n118 ) , .A2( u0_u10_u6_n126 ) , .B2( u0_u10_u6_n151 ) , .C2( u0_u10_u6_n159 ) , .C1( u0_u10_u6_n168 ) , .B1( u0_u10_u6_n169 ) );
  INV_X1 u0_u10_u6_U3 (.A( u0_u10_u6_n110 ) , .ZN( u0_u10_u6_n166 ) );
  NOR2_X1 u0_u10_u6_U30 (.A1( u0_u10_u6_n162 ) , .A2( u0_u10_u6_n165 ) , .ZN( u0_u10_u6_n98 ) );
  AOI211_X1 u0_u10_u6_U31 (.B( u0_u10_u6_n134 ) , .A( u0_u10_u6_n135 ) , .C1( u0_u10_u6_n136 ) , .ZN( u0_u10_u6_n137 ) , .C2( u0_u10_u6_n151 ) );
  NAND4_X1 u0_u10_u6_U32 (.A4( u0_u10_u6_n127 ) , .A3( u0_u10_u6_n128 ) , .A2( u0_u10_u6_n129 ) , .A1( u0_u10_u6_n130 ) , .ZN( u0_u10_u6_n136 ) );
  AOI21_X1 u0_u10_u6_U33 (.B2( u0_u10_u6_n132 ) , .B1( u0_u10_u6_n133 ) , .ZN( u0_u10_u6_n134 ) , .A( u0_u10_u6_n158 ) );
  AOI21_X1 u0_u10_u6_U34 (.B1( u0_u10_u6_n131 ) , .ZN( u0_u10_u6_n135 ) , .A( u0_u10_u6_n144 ) , .B2( u0_u10_u6_n146 ) );
  NAND2_X1 u0_u10_u6_U35 (.A1( u0_u10_u6_n144 ) , .ZN( u0_u10_u6_n151 ) , .A2( u0_u10_u6_n158 ) );
  NAND2_X1 u0_u10_u6_U36 (.ZN( u0_u10_u6_n132 ) , .A1( u0_u10_u6_n91 ) , .A2( u0_u10_u6_n97 ) );
  AOI22_X1 u0_u10_u6_U37 (.B2( u0_u10_u6_n110 ) , .B1( u0_u10_u6_n111 ) , .A1( u0_u10_u6_n112 ) , .ZN( u0_u10_u6_n115 ) , .A2( u0_u10_u6_n161 ) );
  NAND4_X1 u0_u10_u6_U38 (.A3( u0_u10_u6_n109 ) , .ZN( u0_u10_u6_n112 ) , .A4( u0_u10_u6_n132 ) , .A2( u0_u10_u6_n147 ) , .A1( u0_u10_u6_n166 ) );
  NOR2_X1 u0_u10_u6_U39 (.ZN( u0_u10_u6_n109 ) , .A1( u0_u10_u6_n170 ) , .A2( u0_u10_u6_n173 ) );
  INV_X1 u0_u10_u6_U4 (.A( u0_u10_u6_n142 ) , .ZN( u0_u10_u6_n174 ) );
  NOR2_X1 u0_u10_u6_U40 (.A2( u0_u10_u6_n126 ) , .ZN( u0_u10_u6_n155 ) , .A1( u0_u10_u6_n160 ) );
  NAND2_X1 u0_u10_u6_U41 (.ZN( u0_u10_u6_n146 ) , .A2( u0_u10_u6_n94 ) , .A1( u0_u10_u6_n99 ) );
  AOI21_X1 u0_u10_u6_U42 (.A( u0_u10_u6_n144 ) , .B2( u0_u10_u6_n145 ) , .B1( u0_u10_u6_n146 ) , .ZN( u0_u10_u6_n150 ) );
  INV_X1 u0_u10_u6_U43 (.A( u0_u10_u6_n111 ) , .ZN( u0_u10_u6_n158 ) );
  NAND2_X1 u0_u10_u6_U44 (.ZN( u0_u10_u6_n127 ) , .A1( u0_u10_u6_n91 ) , .A2( u0_u10_u6_n92 ) );
  NAND2_X1 u0_u10_u6_U45 (.ZN( u0_u10_u6_n129 ) , .A2( u0_u10_u6_n95 ) , .A1( u0_u10_u6_n96 ) );
  INV_X1 u0_u10_u6_U46 (.A( u0_u10_u6_n144 ) , .ZN( u0_u10_u6_n159 ) );
  NAND2_X1 u0_u10_u6_U47 (.ZN( u0_u10_u6_n145 ) , .A2( u0_u10_u6_n97 ) , .A1( u0_u10_u6_n98 ) );
  NAND2_X1 u0_u10_u6_U48 (.ZN( u0_u10_u6_n148 ) , .A2( u0_u10_u6_n92 ) , .A1( u0_u10_u6_n94 ) );
  NAND2_X1 u0_u10_u6_U49 (.ZN( u0_u10_u6_n108 ) , .A2( u0_u10_u6_n139 ) , .A1( u0_u10_u6_n144 ) );
  NAND2_X1 u0_u10_u6_U5 (.A2( u0_u10_u6_n143 ) , .ZN( u0_u10_u6_n152 ) , .A1( u0_u10_u6_n166 ) );
  NAND2_X1 u0_u10_u6_U50 (.ZN( u0_u10_u6_n121 ) , .A2( u0_u10_u6_n95 ) , .A1( u0_u10_u6_n97 ) );
  NAND2_X1 u0_u10_u6_U51 (.ZN( u0_u10_u6_n107 ) , .A2( u0_u10_u6_n92 ) , .A1( u0_u10_u6_n95 ) );
  AND2_X1 u0_u10_u6_U52 (.ZN( u0_u10_u6_n118 ) , .A2( u0_u10_u6_n91 ) , .A1( u0_u10_u6_n99 ) );
  NAND2_X1 u0_u10_u6_U53 (.ZN( u0_u10_u6_n147 ) , .A2( u0_u10_u6_n98 ) , .A1( u0_u10_u6_n99 ) );
  NAND2_X1 u0_u10_u6_U54 (.ZN( u0_u10_u6_n128 ) , .A1( u0_u10_u6_n94 ) , .A2( u0_u10_u6_n96 ) );
  NAND2_X1 u0_u10_u6_U55 (.ZN( u0_u10_u6_n119 ) , .A2( u0_u10_u6_n95 ) , .A1( u0_u10_u6_n99 ) );
  NAND2_X1 u0_u10_u6_U56 (.ZN( u0_u10_u6_n123 ) , .A2( u0_u10_u6_n91 ) , .A1( u0_u10_u6_n96 ) );
  NAND2_X1 u0_u10_u6_U57 (.ZN( u0_u10_u6_n100 ) , .A2( u0_u10_u6_n92 ) , .A1( u0_u10_u6_n98 ) );
  NAND2_X1 u0_u10_u6_U58 (.ZN( u0_u10_u6_n122 ) , .A1( u0_u10_u6_n94 ) , .A2( u0_u10_u6_n97 ) );
  INV_X1 u0_u10_u6_U59 (.A( u0_u10_u6_n139 ) , .ZN( u0_u10_u6_n160 ) );
  AOI22_X1 u0_u10_u6_U6 (.B2( u0_u10_u6_n101 ) , .A1( u0_u10_u6_n102 ) , .ZN( u0_u10_u6_n103 ) , .B1( u0_u10_u6_n160 ) , .A2( u0_u10_u6_n161 ) );
  NAND2_X1 u0_u10_u6_U60 (.ZN( u0_u10_u6_n113 ) , .A1( u0_u10_u6_n96 ) , .A2( u0_u10_u6_n98 ) );
  NOR2_X1 u0_u10_u6_U61 (.A2( u0_u10_X_40 ) , .A1( u0_u10_X_41 ) , .ZN( u0_u10_u6_n126 ) );
  NOR2_X1 u0_u10_u6_U62 (.A2( u0_u10_X_39 ) , .A1( u0_u10_X_42 ) , .ZN( u0_u10_u6_n92 ) );
  NOR2_X1 u0_u10_u6_U63 (.A2( u0_u10_X_39 ) , .A1( u0_u10_u6_n156 ) , .ZN( u0_u10_u6_n97 ) );
  NOR2_X1 u0_u10_u6_U64 (.A2( u0_u10_X_38 ) , .A1( u0_u10_u6_n165 ) , .ZN( u0_u10_u6_n95 ) );
  NOR2_X1 u0_u10_u6_U65 (.A2( u0_u10_X_41 ) , .ZN( u0_u10_u6_n111 ) , .A1( u0_u10_u6_n157 ) );
  NOR2_X1 u0_u10_u6_U66 (.A2( u0_u10_X_37 ) , .A1( u0_u10_u6_n162 ) , .ZN( u0_u10_u6_n94 ) );
  NOR2_X1 u0_u10_u6_U67 (.A2( u0_u10_X_37 ) , .A1( u0_u10_X_38 ) , .ZN( u0_u10_u6_n91 ) );
  NAND2_X1 u0_u10_u6_U68 (.A1( u0_u10_X_41 ) , .ZN( u0_u10_u6_n144 ) , .A2( u0_u10_u6_n157 ) );
  NAND2_X1 u0_u10_u6_U69 (.A2( u0_u10_X_40 ) , .A1( u0_u10_X_41 ) , .ZN( u0_u10_u6_n139 ) );
  NOR2_X1 u0_u10_u6_U7 (.A1( u0_u10_u6_n118 ) , .ZN( u0_u10_u6_n143 ) , .A2( u0_u10_u6_n168 ) );
  AND2_X1 u0_u10_u6_U70 (.A1( u0_u10_X_39 ) , .A2( u0_u10_u6_n156 ) , .ZN( u0_u10_u6_n96 ) );
  AND2_X1 u0_u10_u6_U71 (.A1( u0_u10_X_39 ) , .A2( u0_u10_X_42 ) , .ZN( u0_u10_u6_n99 ) );
  INV_X1 u0_u10_u6_U72 (.A( u0_u10_X_40 ) , .ZN( u0_u10_u6_n157 ) );
  INV_X1 u0_u10_u6_U73 (.A( u0_u10_X_37 ) , .ZN( u0_u10_u6_n165 ) );
  INV_X1 u0_u10_u6_U74 (.A( u0_u10_X_38 ) , .ZN( u0_u10_u6_n162 ) );
  INV_X1 u0_u10_u6_U75 (.A( u0_u10_X_42 ) , .ZN( u0_u10_u6_n156 ) );
  NAND4_X1 u0_u10_u6_U76 (.ZN( u0_out10_32 ) , .A4( u0_u10_u6_n103 ) , .A3( u0_u10_u6_n104 ) , .A2( u0_u10_u6_n105 ) , .A1( u0_u10_u6_n106 ) );
  AOI22_X1 u0_u10_u6_U77 (.ZN( u0_u10_u6_n105 ) , .A2( u0_u10_u6_n108 ) , .A1( u0_u10_u6_n118 ) , .B2( u0_u10_u6_n126 ) , .B1( u0_u10_u6_n171 ) );
  AOI22_X1 u0_u10_u6_U78 (.ZN( u0_u10_u6_n104 ) , .A1( u0_u10_u6_n111 ) , .B1( u0_u10_u6_n124 ) , .B2( u0_u10_u6_n151 ) , .A2( u0_u10_u6_n93 ) );
  NAND4_X1 u0_u10_u6_U79 (.ZN( u0_out10_12 ) , .A4( u0_u10_u6_n114 ) , .A3( u0_u10_u6_n115 ) , .A2( u0_u10_u6_n116 ) , .A1( u0_u10_u6_n117 ) );
  INV_X1 u0_u10_u6_U8 (.ZN( u0_u10_u6_n172 ) , .A( u0_u10_u6_n88 ) );
  OAI22_X1 u0_u10_u6_U80 (.B2( u0_u10_u6_n111 ) , .ZN( u0_u10_u6_n116 ) , .B1( u0_u10_u6_n126 ) , .A2( u0_u10_u6_n164 ) , .A1( u0_u10_u6_n167 ) );
  OAI21_X1 u0_u10_u6_U81 (.A( u0_u10_u6_n108 ) , .ZN( u0_u10_u6_n117 ) , .B2( u0_u10_u6_n141 ) , .B1( u0_u10_u6_n163 ) );
  OAI211_X1 u0_u10_u6_U82 (.ZN( u0_out10_7 ) , .B( u0_u10_u6_n153 ) , .C2( u0_u10_u6_n154 ) , .C1( u0_u10_u6_n155 ) , .A( u0_u10_u6_n174 ) );
  NOR3_X1 u0_u10_u6_U83 (.A1( u0_u10_u6_n141 ) , .ZN( u0_u10_u6_n154 ) , .A3( u0_u10_u6_n164 ) , .A2( u0_u10_u6_n171 ) );
  AOI211_X1 u0_u10_u6_U84 (.B( u0_u10_u6_n149 ) , .A( u0_u10_u6_n150 ) , .C2( u0_u10_u6_n151 ) , .C1( u0_u10_u6_n152 ) , .ZN( u0_u10_u6_n153 ) );
  OAI211_X1 u0_u10_u6_U85 (.ZN( u0_out10_22 ) , .B( u0_u10_u6_n137 ) , .A( u0_u10_u6_n138 ) , .C2( u0_u10_u6_n139 ) , .C1( u0_u10_u6_n140 ) );
  AOI22_X1 u0_u10_u6_U86 (.B1( u0_u10_u6_n124 ) , .A2( u0_u10_u6_n125 ) , .A1( u0_u10_u6_n126 ) , .ZN( u0_u10_u6_n138 ) , .B2( u0_u10_u6_n161 ) );
  AND4_X1 u0_u10_u6_U87 (.A3( u0_u10_u6_n119 ) , .A1( u0_u10_u6_n120 ) , .A4( u0_u10_u6_n129 ) , .ZN( u0_u10_u6_n140 ) , .A2( u0_u10_u6_n143 ) );
  NAND3_X1 u0_u10_u6_U88 (.A2( u0_u10_u6_n123 ) , .ZN( u0_u10_u6_n125 ) , .A1( u0_u10_u6_n130 ) , .A3( u0_u10_u6_n131 ) );
  NAND3_X1 u0_u10_u6_U89 (.A3( u0_u10_u6_n133 ) , .ZN( u0_u10_u6_n141 ) , .A1( u0_u10_u6_n145 ) , .A2( u0_u10_u6_n148 ) );
  OAI21_X1 u0_u10_u6_U9 (.A( u0_u10_u6_n159 ) , .B1( u0_u10_u6_n169 ) , .B2( u0_u10_u6_n173 ) , .ZN( u0_u10_u6_n90 ) );
  NAND3_X1 u0_u10_u6_U90 (.ZN( u0_u10_u6_n101 ) , .A3( u0_u10_u6_n107 ) , .A2( u0_u10_u6_n121 ) , .A1( u0_u10_u6_n127 ) );
  NAND3_X1 u0_u10_u6_U91 (.ZN( u0_u10_u6_n102 ) , .A3( u0_u10_u6_n130 ) , .A2( u0_u10_u6_n145 ) , .A1( u0_u10_u6_n166 ) );
  NAND3_X1 u0_u10_u6_U92 (.A3( u0_u10_u6_n113 ) , .A1( u0_u10_u6_n119 ) , .A2( u0_u10_u6_n123 ) , .ZN( u0_u10_u6_n93 ) );
  NAND3_X1 u0_u10_u6_U93 (.ZN( u0_u10_u6_n142 ) , .A2( u0_u10_u6_n172 ) , .A3( u0_u10_u6_n89 ) , .A1( u0_u10_u6_n90 ) );
  XOR2_X1 u0_u11_U1 (.B( u0_K12_9 ) , .A( u0_R10_6 ) , .Z( u0_u11_X_9 ) );
  XOR2_X1 u0_u11_U13 (.B( u0_K12_42 ) , .A( u0_R10_29 ) , .Z( u0_u11_X_42 ) );
  XOR2_X1 u0_u11_U14 (.B( u0_K12_41 ) , .A( u0_R10_28 ) , .Z( u0_u11_X_41 ) );
  XOR2_X1 u0_u11_U15 (.B( u0_K12_40 ) , .A( u0_R10_27 ) , .Z( u0_u11_X_40 ) );
  XOR2_X1 u0_u11_U17 (.B( u0_K12_39 ) , .A( u0_R10_26 ) , .Z( u0_u11_X_39 ) );
  XOR2_X1 u0_u11_U18 (.B( u0_K12_38 ) , .A( u0_R10_25 ) , .Z( u0_u11_X_38 ) );
  XOR2_X1 u0_u11_U19 (.B( u0_K12_37 ) , .A( u0_R10_24 ) , .Z( u0_u11_X_37 ) );
  XOR2_X1 u0_u11_U2 (.B( u0_K12_8 ) , .A( u0_R10_5 ) , .Z( u0_u11_X_8 ) );
  XOR2_X1 u0_u11_U3 (.B( u0_K12_7 ) , .A( u0_R10_4 ) , .Z( u0_u11_X_7 ) );
  XOR2_X1 u0_u11_U40 (.B( u0_K12_18 ) , .A( u0_R10_13 ) , .Z( u0_u11_X_18 ) );
  XOR2_X1 u0_u11_U41 (.B( u0_K12_17 ) , .A( u0_R10_12 ) , .Z( u0_u11_X_17 ) );
  XOR2_X1 u0_u11_U42 (.B( u0_K12_16 ) , .A( u0_R10_11 ) , .Z( u0_u11_X_16 ) );
  XOR2_X1 u0_u11_U43 (.B( u0_K12_15 ) , .A( u0_R10_10 ) , .Z( u0_u11_X_15 ) );
  XOR2_X1 u0_u11_U44 (.B( u0_K12_14 ) , .A( u0_R10_9 ) , .Z( u0_u11_X_14 ) );
  XOR2_X1 u0_u11_U45 (.B( u0_K12_13 ) , .A( u0_R10_8 ) , .Z( u0_u11_X_13 ) );
  XOR2_X1 u0_u11_U46 (.B( u0_K12_12 ) , .A( u0_R10_9 ) , .Z( u0_u11_X_12 ) );
  XOR2_X1 u0_u11_U47 (.B( u0_K12_11 ) , .A( u0_R10_8 ) , .Z( u0_u11_X_11 ) );
  XOR2_X1 u0_u11_U48 (.B( u0_K12_10 ) , .A( u0_R10_7 ) , .Z( u0_u11_X_10 ) );
  NOR2_X1 u0_u11_u1_U10 (.A1( u0_u11_u1_n112 ) , .A2( u0_u11_u1_n116 ) , .ZN( u0_u11_u1_n118 ) );
  NAND3_X1 u0_u11_u1_U100 (.ZN( u0_u11_u1_n113 ) , .A1( u0_u11_u1_n120 ) , .A3( u0_u11_u1_n133 ) , .A2( u0_u11_u1_n155 ) );
  OAI21_X1 u0_u11_u1_U11 (.ZN( u0_u11_u1_n101 ) , .B1( u0_u11_u1_n141 ) , .A( u0_u11_u1_n146 ) , .B2( u0_u11_u1_n183 ) );
  AOI21_X1 u0_u11_u1_U12 (.B2( u0_u11_u1_n155 ) , .B1( u0_u11_u1_n156 ) , .ZN( u0_u11_u1_n157 ) , .A( u0_u11_u1_n174 ) );
  NAND2_X1 u0_u11_u1_U13 (.ZN( u0_u11_u1_n140 ) , .A2( u0_u11_u1_n150 ) , .A1( u0_u11_u1_n155 ) );
  NAND2_X1 u0_u11_u1_U14 (.A1( u0_u11_u1_n131 ) , .ZN( u0_u11_u1_n147 ) , .A2( u0_u11_u1_n153 ) );
  INV_X1 u0_u11_u1_U15 (.A( u0_u11_u1_n139 ) , .ZN( u0_u11_u1_n174 ) );
  OR4_X1 u0_u11_u1_U16 (.A4( u0_u11_u1_n106 ) , .A3( u0_u11_u1_n107 ) , .ZN( u0_u11_u1_n108 ) , .A1( u0_u11_u1_n117 ) , .A2( u0_u11_u1_n184 ) );
  AOI21_X1 u0_u11_u1_U17 (.ZN( u0_u11_u1_n106 ) , .A( u0_u11_u1_n112 ) , .B1( u0_u11_u1_n154 ) , .B2( u0_u11_u1_n156 ) );
  AOI21_X1 u0_u11_u1_U18 (.ZN( u0_u11_u1_n107 ) , .B1( u0_u11_u1_n134 ) , .B2( u0_u11_u1_n149 ) , .A( u0_u11_u1_n174 ) );
  INV_X1 u0_u11_u1_U19 (.A( u0_u11_u1_n101 ) , .ZN( u0_u11_u1_n184 ) );
  INV_X1 u0_u11_u1_U20 (.A( u0_u11_u1_n112 ) , .ZN( u0_u11_u1_n171 ) );
  NAND2_X1 u0_u11_u1_U21 (.ZN( u0_u11_u1_n141 ) , .A1( u0_u11_u1_n153 ) , .A2( u0_u11_u1_n156 ) );
  AND2_X1 u0_u11_u1_U22 (.A1( u0_u11_u1_n123 ) , .ZN( u0_u11_u1_n134 ) , .A2( u0_u11_u1_n161 ) );
  NAND2_X1 u0_u11_u1_U23 (.A2( u0_u11_u1_n115 ) , .A1( u0_u11_u1_n116 ) , .ZN( u0_u11_u1_n148 ) );
  NAND2_X1 u0_u11_u1_U24 (.A2( u0_u11_u1_n133 ) , .A1( u0_u11_u1_n135 ) , .ZN( u0_u11_u1_n159 ) );
  NAND2_X1 u0_u11_u1_U25 (.A2( u0_u11_u1_n115 ) , .A1( u0_u11_u1_n120 ) , .ZN( u0_u11_u1_n132 ) );
  INV_X1 u0_u11_u1_U26 (.A( u0_u11_u1_n154 ) , .ZN( u0_u11_u1_n178 ) );
  INV_X1 u0_u11_u1_U27 (.A( u0_u11_u1_n151 ) , .ZN( u0_u11_u1_n183 ) );
  AND2_X1 u0_u11_u1_U28 (.A1( u0_u11_u1_n129 ) , .A2( u0_u11_u1_n133 ) , .ZN( u0_u11_u1_n149 ) );
  INV_X1 u0_u11_u1_U29 (.A( u0_u11_u1_n131 ) , .ZN( u0_u11_u1_n180 ) );
  INV_X1 u0_u11_u1_U3 (.A( u0_u11_u1_n159 ) , .ZN( u0_u11_u1_n182 ) );
  OAI221_X1 u0_u11_u1_U30 (.A( u0_u11_u1_n119 ) , .C2( u0_u11_u1_n129 ) , .ZN( u0_u11_u1_n138 ) , .B2( u0_u11_u1_n152 ) , .C1( u0_u11_u1_n174 ) , .B1( u0_u11_u1_n187 ) );
  INV_X1 u0_u11_u1_U31 (.A( u0_u11_u1_n148 ) , .ZN( u0_u11_u1_n187 ) );
  AOI211_X1 u0_u11_u1_U32 (.B( u0_u11_u1_n117 ) , .A( u0_u11_u1_n118 ) , .ZN( u0_u11_u1_n119 ) , .C2( u0_u11_u1_n146 ) , .C1( u0_u11_u1_n159 ) );
  NOR2_X1 u0_u11_u1_U33 (.A1( u0_u11_u1_n168 ) , .A2( u0_u11_u1_n176 ) , .ZN( u0_u11_u1_n98 ) );
  AOI211_X1 u0_u11_u1_U34 (.B( u0_u11_u1_n162 ) , .A( u0_u11_u1_n163 ) , .C2( u0_u11_u1_n164 ) , .ZN( u0_u11_u1_n165 ) , .C1( u0_u11_u1_n171 ) );
  AOI21_X1 u0_u11_u1_U35 (.A( u0_u11_u1_n160 ) , .B2( u0_u11_u1_n161 ) , .ZN( u0_u11_u1_n162 ) , .B1( u0_u11_u1_n182 ) );
  OR2_X1 u0_u11_u1_U36 (.A2( u0_u11_u1_n157 ) , .A1( u0_u11_u1_n158 ) , .ZN( u0_u11_u1_n163 ) );
  NAND2_X1 u0_u11_u1_U37 (.A1( u0_u11_u1_n128 ) , .ZN( u0_u11_u1_n146 ) , .A2( u0_u11_u1_n160 ) );
  NAND2_X1 u0_u11_u1_U38 (.A2( u0_u11_u1_n112 ) , .ZN( u0_u11_u1_n139 ) , .A1( u0_u11_u1_n152 ) );
  NAND2_X1 u0_u11_u1_U39 (.A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n156 ) , .A2( u0_u11_u1_n99 ) );
  AOI221_X1 u0_u11_u1_U4 (.A( u0_u11_u1_n138 ) , .C2( u0_u11_u1_n139 ) , .C1( u0_u11_u1_n140 ) , .B2( u0_u11_u1_n141 ) , .ZN( u0_u11_u1_n142 ) , .B1( u0_u11_u1_n175 ) );
  AOI221_X1 u0_u11_u1_U40 (.B1( u0_u11_u1_n140 ) , .ZN( u0_u11_u1_n167 ) , .B2( u0_u11_u1_n172 ) , .C2( u0_u11_u1_n175 ) , .C1( u0_u11_u1_n178 ) , .A( u0_u11_u1_n188 ) );
  INV_X1 u0_u11_u1_U41 (.ZN( u0_u11_u1_n188 ) , .A( u0_u11_u1_n97 ) );
  AOI211_X1 u0_u11_u1_U42 (.A( u0_u11_u1_n118 ) , .C1( u0_u11_u1_n132 ) , .C2( u0_u11_u1_n139 ) , .B( u0_u11_u1_n96 ) , .ZN( u0_u11_u1_n97 ) );
  AOI21_X1 u0_u11_u1_U43 (.B2( u0_u11_u1_n121 ) , .B1( u0_u11_u1_n135 ) , .A( u0_u11_u1_n152 ) , .ZN( u0_u11_u1_n96 ) );
  NOR2_X1 u0_u11_u1_U44 (.ZN( u0_u11_u1_n117 ) , .A1( u0_u11_u1_n121 ) , .A2( u0_u11_u1_n160 ) );
  OAI21_X1 u0_u11_u1_U45 (.B2( u0_u11_u1_n123 ) , .ZN( u0_u11_u1_n145 ) , .B1( u0_u11_u1_n160 ) , .A( u0_u11_u1_n185 ) );
  INV_X1 u0_u11_u1_U46 (.A( u0_u11_u1_n122 ) , .ZN( u0_u11_u1_n185 ) );
  AOI21_X1 u0_u11_u1_U47 (.B2( u0_u11_u1_n120 ) , .B1( u0_u11_u1_n121 ) , .ZN( u0_u11_u1_n122 ) , .A( u0_u11_u1_n128 ) );
  AOI21_X1 u0_u11_u1_U48 (.A( u0_u11_u1_n128 ) , .B2( u0_u11_u1_n129 ) , .ZN( u0_u11_u1_n130 ) , .B1( u0_u11_u1_n150 ) );
  NAND2_X1 u0_u11_u1_U49 (.ZN( u0_u11_u1_n112 ) , .A1( u0_u11_u1_n169 ) , .A2( u0_u11_u1_n170 ) );
  AOI211_X1 u0_u11_u1_U5 (.ZN( u0_u11_u1_n124 ) , .A( u0_u11_u1_n138 ) , .C2( u0_u11_u1_n139 ) , .B( u0_u11_u1_n145 ) , .C1( u0_u11_u1_n147 ) );
  NAND2_X1 u0_u11_u1_U50 (.ZN( u0_u11_u1_n129 ) , .A2( u0_u11_u1_n95 ) , .A1( u0_u11_u1_n98 ) );
  NAND2_X1 u0_u11_u1_U51 (.A1( u0_u11_u1_n102 ) , .ZN( u0_u11_u1_n154 ) , .A2( u0_u11_u1_n99 ) );
  NAND2_X1 u0_u11_u1_U52 (.A2( u0_u11_u1_n100 ) , .ZN( u0_u11_u1_n135 ) , .A1( u0_u11_u1_n99 ) );
  AOI21_X1 u0_u11_u1_U53 (.A( u0_u11_u1_n152 ) , .B2( u0_u11_u1_n153 ) , .B1( u0_u11_u1_n154 ) , .ZN( u0_u11_u1_n158 ) );
  INV_X1 u0_u11_u1_U54 (.A( u0_u11_u1_n160 ) , .ZN( u0_u11_u1_n175 ) );
  NAND2_X1 u0_u11_u1_U55 (.A1( u0_u11_u1_n100 ) , .ZN( u0_u11_u1_n116 ) , .A2( u0_u11_u1_n95 ) );
  NAND2_X1 u0_u11_u1_U56 (.A1( u0_u11_u1_n102 ) , .ZN( u0_u11_u1_n131 ) , .A2( u0_u11_u1_n95 ) );
  NAND2_X1 u0_u11_u1_U57 (.A2( u0_u11_u1_n104 ) , .ZN( u0_u11_u1_n121 ) , .A1( u0_u11_u1_n98 ) );
  NAND2_X1 u0_u11_u1_U58 (.A1( u0_u11_u1_n103 ) , .ZN( u0_u11_u1_n153 ) , .A2( u0_u11_u1_n98 ) );
  NAND2_X1 u0_u11_u1_U59 (.A2( u0_u11_u1_n104 ) , .A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n133 ) );
  AOI22_X1 u0_u11_u1_U6 (.B2( u0_u11_u1_n113 ) , .A2( u0_u11_u1_n114 ) , .ZN( u0_u11_u1_n125 ) , .A1( u0_u11_u1_n171 ) , .B1( u0_u11_u1_n173 ) );
  NAND2_X1 u0_u11_u1_U60 (.ZN( u0_u11_u1_n150 ) , .A2( u0_u11_u1_n98 ) , .A1( u0_u11_u1_n99 ) );
  NAND2_X1 u0_u11_u1_U61 (.A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n155 ) , .A2( u0_u11_u1_n95 ) );
  OAI21_X1 u0_u11_u1_U62 (.ZN( u0_u11_u1_n109 ) , .B1( u0_u11_u1_n129 ) , .B2( u0_u11_u1_n160 ) , .A( u0_u11_u1_n167 ) );
  NAND2_X1 u0_u11_u1_U63 (.A2( u0_u11_u1_n100 ) , .A1( u0_u11_u1_n103 ) , .ZN( u0_u11_u1_n120 ) );
  NAND2_X1 u0_u11_u1_U64 (.A1( u0_u11_u1_n102 ) , .A2( u0_u11_u1_n104 ) , .ZN( u0_u11_u1_n115 ) );
  NAND2_X1 u0_u11_u1_U65 (.A2( u0_u11_u1_n100 ) , .A1( u0_u11_u1_n104 ) , .ZN( u0_u11_u1_n151 ) );
  NAND2_X1 u0_u11_u1_U66 (.A2( u0_u11_u1_n103 ) , .A1( u0_u11_u1_n105 ) , .ZN( u0_u11_u1_n161 ) );
  INV_X1 u0_u11_u1_U67 (.A( u0_u11_u1_n152 ) , .ZN( u0_u11_u1_n173 ) );
  INV_X1 u0_u11_u1_U68 (.A( u0_u11_u1_n128 ) , .ZN( u0_u11_u1_n172 ) );
  NAND2_X1 u0_u11_u1_U69 (.A2( u0_u11_u1_n102 ) , .A1( u0_u11_u1_n103 ) , .ZN( u0_u11_u1_n123 ) );
  NAND2_X1 u0_u11_u1_U7 (.ZN( u0_u11_u1_n114 ) , .A1( u0_u11_u1_n134 ) , .A2( u0_u11_u1_n156 ) );
  NOR2_X1 u0_u11_u1_U70 (.A2( u0_u11_X_7 ) , .A1( u0_u11_X_8 ) , .ZN( u0_u11_u1_n95 ) );
  NOR2_X1 u0_u11_u1_U71 (.A1( u0_u11_X_12 ) , .A2( u0_u11_X_9 ) , .ZN( u0_u11_u1_n100 ) );
  NOR2_X1 u0_u11_u1_U72 (.A2( u0_u11_X_8 ) , .A1( u0_u11_u1_n177 ) , .ZN( u0_u11_u1_n99 ) );
  NOR2_X1 u0_u11_u1_U73 (.A2( u0_u11_X_12 ) , .ZN( u0_u11_u1_n102 ) , .A1( u0_u11_u1_n176 ) );
  NOR2_X1 u0_u11_u1_U74 (.A2( u0_u11_X_9 ) , .ZN( u0_u11_u1_n105 ) , .A1( u0_u11_u1_n168 ) );
  NAND2_X1 u0_u11_u1_U75 (.A1( u0_u11_X_10 ) , .ZN( u0_u11_u1_n160 ) , .A2( u0_u11_u1_n169 ) );
  NAND2_X1 u0_u11_u1_U76 (.A2( u0_u11_X_10 ) , .A1( u0_u11_X_11 ) , .ZN( u0_u11_u1_n152 ) );
  NAND2_X1 u0_u11_u1_U77 (.A1( u0_u11_X_11 ) , .ZN( u0_u11_u1_n128 ) , .A2( u0_u11_u1_n170 ) );
  AND2_X1 u0_u11_u1_U78 (.A2( u0_u11_X_7 ) , .A1( u0_u11_X_8 ) , .ZN( u0_u11_u1_n104 ) );
  AND2_X1 u0_u11_u1_U79 (.A1( u0_u11_X_8 ) , .ZN( u0_u11_u1_n103 ) , .A2( u0_u11_u1_n177 ) );
  AOI22_X1 u0_u11_u1_U8 (.B2( u0_u11_u1_n136 ) , .A2( u0_u11_u1_n137 ) , .ZN( u0_u11_u1_n143 ) , .A1( u0_u11_u1_n171 ) , .B1( u0_u11_u1_n173 ) );
  INV_X1 u0_u11_u1_U80 (.A( u0_u11_X_10 ) , .ZN( u0_u11_u1_n170 ) );
  INV_X1 u0_u11_u1_U81 (.A( u0_u11_X_9 ) , .ZN( u0_u11_u1_n176 ) );
  INV_X1 u0_u11_u1_U82 (.A( u0_u11_X_11 ) , .ZN( u0_u11_u1_n169 ) );
  INV_X1 u0_u11_u1_U83 (.A( u0_u11_X_12 ) , .ZN( u0_u11_u1_n168 ) );
  INV_X1 u0_u11_u1_U84 (.A( u0_u11_X_7 ) , .ZN( u0_u11_u1_n177 ) );
  NAND4_X1 u0_u11_u1_U85 (.ZN( u0_out11_28 ) , .A4( u0_u11_u1_n124 ) , .A3( u0_u11_u1_n125 ) , .A2( u0_u11_u1_n126 ) , .A1( u0_u11_u1_n127 ) );
  OAI21_X1 u0_u11_u1_U86 (.ZN( u0_u11_u1_n127 ) , .B2( u0_u11_u1_n139 ) , .B1( u0_u11_u1_n175 ) , .A( u0_u11_u1_n183 ) );
  OAI21_X1 u0_u11_u1_U87 (.ZN( u0_u11_u1_n126 ) , .B2( u0_u11_u1_n140 ) , .A( u0_u11_u1_n146 ) , .B1( u0_u11_u1_n178 ) );
  NAND4_X1 u0_u11_u1_U88 (.ZN( u0_out11_18 ) , .A4( u0_u11_u1_n165 ) , .A3( u0_u11_u1_n166 ) , .A1( u0_u11_u1_n167 ) , .A2( u0_u11_u1_n186 ) );
  AOI22_X1 u0_u11_u1_U89 (.B2( u0_u11_u1_n146 ) , .B1( u0_u11_u1_n147 ) , .A2( u0_u11_u1_n148 ) , .ZN( u0_u11_u1_n166 ) , .A1( u0_u11_u1_n172 ) );
  INV_X1 u0_u11_u1_U9 (.A( u0_u11_u1_n147 ) , .ZN( u0_u11_u1_n181 ) );
  INV_X1 u0_u11_u1_U90 (.A( u0_u11_u1_n145 ) , .ZN( u0_u11_u1_n186 ) );
  NAND4_X1 u0_u11_u1_U91 (.ZN( u0_out11_2 ) , .A4( u0_u11_u1_n142 ) , .A3( u0_u11_u1_n143 ) , .A2( u0_u11_u1_n144 ) , .A1( u0_u11_u1_n179 ) );
  OAI21_X1 u0_u11_u1_U92 (.B2( u0_u11_u1_n132 ) , .ZN( u0_u11_u1_n144 ) , .A( u0_u11_u1_n146 ) , .B1( u0_u11_u1_n180 ) );
  INV_X1 u0_u11_u1_U93 (.A( u0_u11_u1_n130 ) , .ZN( u0_u11_u1_n179 ) );
  OR4_X1 u0_u11_u1_U94 (.ZN( u0_out11_13 ) , .A4( u0_u11_u1_n108 ) , .A3( u0_u11_u1_n109 ) , .A2( u0_u11_u1_n110 ) , .A1( u0_u11_u1_n111 ) );
  AOI21_X1 u0_u11_u1_U95 (.ZN( u0_u11_u1_n111 ) , .A( u0_u11_u1_n128 ) , .B2( u0_u11_u1_n131 ) , .B1( u0_u11_u1_n135 ) );
  AOI21_X1 u0_u11_u1_U96 (.ZN( u0_u11_u1_n110 ) , .A( u0_u11_u1_n116 ) , .B1( u0_u11_u1_n152 ) , .B2( u0_u11_u1_n160 ) );
  NAND3_X1 u0_u11_u1_U97 (.A3( u0_u11_u1_n149 ) , .A2( u0_u11_u1_n150 ) , .A1( u0_u11_u1_n151 ) , .ZN( u0_u11_u1_n164 ) );
  NAND3_X1 u0_u11_u1_U98 (.A3( u0_u11_u1_n134 ) , .A2( u0_u11_u1_n135 ) , .ZN( u0_u11_u1_n136 ) , .A1( u0_u11_u1_n151 ) );
  NAND3_X1 u0_u11_u1_U99 (.A1( u0_u11_u1_n133 ) , .ZN( u0_u11_u1_n137 ) , .A2( u0_u11_u1_n154 ) , .A3( u0_u11_u1_n181 ) );
  OAI22_X1 u0_u11_u2_U10 (.ZN( u0_u11_u2_n109 ) , .A2( u0_u11_u2_n113 ) , .B2( u0_u11_u2_n133 ) , .B1( u0_u11_u2_n167 ) , .A1( u0_u11_u2_n168 ) );
  NAND3_X1 u0_u11_u2_U100 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n98 ) );
  OAI22_X1 u0_u11_u2_U11 (.B1( u0_u11_u2_n151 ) , .A2( u0_u11_u2_n152 ) , .A1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n160 ) , .B2( u0_u11_u2_n168 ) );
  NOR3_X1 u0_u11_u2_U12 (.A1( u0_u11_u2_n150 ) , .ZN( u0_u11_u2_n151 ) , .A3( u0_u11_u2_n175 ) , .A2( u0_u11_u2_n188 ) );
  AOI21_X1 u0_u11_u2_U13 (.ZN( u0_u11_u2_n144 ) , .B2( u0_u11_u2_n155 ) , .A( u0_u11_u2_n172 ) , .B1( u0_u11_u2_n185 ) );
  AOI21_X1 u0_u11_u2_U14 (.B2( u0_u11_u2_n143 ) , .ZN( u0_u11_u2_n145 ) , .B1( u0_u11_u2_n152 ) , .A( u0_u11_u2_n171 ) );
  AOI21_X1 u0_u11_u2_U15 (.B2( u0_u11_u2_n120 ) , .B1( u0_u11_u2_n121 ) , .ZN( u0_u11_u2_n126 ) , .A( u0_u11_u2_n167 ) );
  INV_X1 u0_u11_u2_U16 (.A( u0_u11_u2_n156 ) , .ZN( u0_u11_u2_n171 ) );
  INV_X1 u0_u11_u2_U17 (.A( u0_u11_u2_n120 ) , .ZN( u0_u11_u2_n188 ) );
  NAND2_X1 u0_u11_u2_U18 (.A2( u0_u11_u2_n122 ) , .ZN( u0_u11_u2_n150 ) , .A1( u0_u11_u2_n152 ) );
  INV_X1 u0_u11_u2_U19 (.A( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n170 ) );
  INV_X1 u0_u11_u2_U20 (.A( u0_u11_u2_n137 ) , .ZN( u0_u11_u2_n173 ) );
  NAND2_X1 u0_u11_u2_U21 (.A1( u0_u11_u2_n132 ) , .A2( u0_u11_u2_n139 ) , .ZN( u0_u11_u2_n157 ) );
  INV_X1 u0_u11_u2_U22 (.A( u0_u11_u2_n113 ) , .ZN( u0_u11_u2_n178 ) );
  INV_X1 u0_u11_u2_U23 (.A( u0_u11_u2_n139 ) , .ZN( u0_u11_u2_n175 ) );
  INV_X1 u0_u11_u2_U24 (.A( u0_u11_u2_n155 ) , .ZN( u0_u11_u2_n181 ) );
  INV_X1 u0_u11_u2_U25 (.A( u0_u11_u2_n119 ) , .ZN( u0_u11_u2_n177 ) );
  INV_X1 u0_u11_u2_U26 (.A( u0_u11_u2_n116 ) , .ZN( u0_u11_u2_n180 ) );
  INV_X1 u0_u11_u2_U27 (.A( u0_u11_u2_n131 ) , .ZN( u0_u11_u2_n179 ) );
  INV_X1 u0_u11_u2_U28 (.A( u0_u11_u2_n154 ) , .ZN( u0_u11_u2_n176 ) );
  NAND2_X1 u0_u11_u2_U29 (.A2( u0_u11_u2_n116 ) , .A1( u0_u11_u2_n117 ) , .ZN( u0_u11_u2_n118 ) );
  NOR2_X1 u0_u11_u2_U3 (.ZN( u0_u11_u2_n121 ) , .A2( u0_u11_u2_n177 ) , .A1( u0_u11_u2_n180 ) );
  INV_X1 u0_u11_u2_U30 (.A( u0_u11_u2_n132 ) , .ZN( u0_u11_u2_n182 ) );
  INV_X1 u0_u11_u2_U31 (.A( u0_u11_u2_n158 ) , .ZN( u0_u11_u2_n183 ) );
  OAI21_X1 u0_u11_u2_U32 (.A( u0_u11_u2_n156 ) , .B1( u0_u11_u2_n157 ) , .ZN( u0_u11_u2_n158 ) , .B2( u0_u11_u2_n179 ) );
  NOR2_X1 u0_u11_u2_U33 (.ZN( u0_u11_u2_n156 ) , .A1( u0_u11_u2_n166 ) , .A2( u0_u11_u2_n169 ) );
  NOR2_X1 u0_u11_u2_U34 (.A2( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n137 ) , .A1( u0_u11_u2_n140 ) );
  NOR2_X1 u0_u11_u2_U35 (.A2( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n153 ) , .A1( u0_u11_u2_n156 ) );
  AOI211_X1 u0_u11_u2_U36 (.ZN( u0_u11_u2_n130 ) , .C1( u0_u11_u2_n138 ) , .C2( u0_u11_u2_n179 ) , .B( u0_u11_u2_n96 ) , .A( u0_u11_u2_n97 ) );
  OAI22_X1 u0_u11_u2_U37 (.B1( u0_u11_u2_n133 ) , .A2( u0_u11_u2_n137 ) , .A1( u0_u11_u2_n152 ) , .B2( u0_u11_u2_n168 ) , .ZN( u0_u11_u2_n97 ) );
  OAI221_X1 u0_u11_u2_U38 (.B1( u0_u11_u2_n113 ) , .C1( u0_u11_u2_n132 ) , .A( u0_u11_u2_n149 ) , .B2( u0_u11_u2_n171 ) , .C2( u0_u11_u2_n172 ) , .ZN( u0_u11_u2_n96 ) );
  OAI221_X1 u0_u11_u2_U39 (.A( u0_u11_u2_n115 ) , .C2( u0_u11_u2_n123 ) , .B2( u0_u11_u2_n143 ) , .B1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n163 ) , .C1( u0_u11_u2_n168 ) );
  INV_X1 u0_u11_u2_U4 (.A( u0_u11_u2_n134 ) , .ZN( u0_u11_u2_n185 ) );
  OAI21_X1 u0_u11_u2_U40 (.A( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n115 ) , .B1( u0_u11_u2_n176 ) , .B2( u0_u11_u2_n178 ) );
  OAI221_X1 u0_u11_u2_U41 (.A( u0_u11_u2_n135 ) , .B2( u0_u11_u2_n136 ) , .B1( u0_u11_u2_n137 ) , .ZN( u0_u11_u2_n162 ) , .C2( u0_u11_u2_n167 ) , .C1( u0_u11_u2_n185 ) );
  AND3_X1 u0_u11_u2_U42 (.A3( u0_u11_u2_n131 ) , .A2( u0_u11_u2_n132 ) , .A1( u0_u11_u2_n133 ) , .ZN( u0_u11_u2_n136 ) );
  AOI22_X1 u0_u11_u2_U43 (.ZN( u0_u11_u2_n135 ) , .B1( u0_u11_u2_n140 ) , .A1( u0_u11_u2_n156 ) , .B2( u0_u11_u2_n180 ) , .A2( u0_u11_u2_n188 ) );
  AOI21_X1 u0_u11_u2_U44 (.ZN( u0_u11_u2_n149 ) , .B1( u0_u11_u2_n173 ) , .B2( u0_u11_u2_n188 ) , .A( u0_u11_u2_n95 ) );
  AND3_X1 u0_u11_u2_U45 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n156 ) , .ZN( u0_u11_u2_n95 ) );
  OAI21_X1 u0_u11_u2_U46 (.A( u0_u11_u2_n101 ) , .B2( u0_u11_u2_n121 ) , .B1( u0_u11_u2_n153 ) , .ZN( u0_u11_u2_n164 ) );
  NAND2_X1 u0_u11_u2_U47 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n155 ) );
  NAND2_X1 u0_u11_u2_U48 (.A2( u0_u11_u2_n105 ) , .A1( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n143 ) );
  NAND2_X1 u0_u11_u2_U49 (.A1( u0_u11_u2_n104 ) , .A2( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n152 ) );
  INV_X1 u0_u11_u2_U5 (.A( u0_u11_u2_n150 ) , .ZN( u0_u11_u2_n184 ) );
  NAND2_X1 u0_u11_u2_U50 (.A1( u0_u11_u2_n100 ) , .A2( u0_u11_u2_n105 ) , .ZN( u0_u11_u2_n132 ) );
  INV_X1 u0_u11_u2_U51 (.A( u0_u11_u2_n140 ) , .ZN( u0_u11_u2_n168 ) );
  INV_X1 u0_u11_u2_U52 (.A( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n167 ) );
  OAI21_X1 u0_u11_u2_U53 (.A( u0_u11_u2_n141 ) , .B2( u0_u11_u2_n142 ) , .ZN( u0_u11_u2_n146 ) , .B1( u0_u11_u2_n153 ) );
  OAI21_X1 u0_u11_u2_U54 (.A( u0_u11_u2_n140 ) , .ZN( u0_u11_u2_n141 ) , .B1( u0_u11_u2_n176 ) , .B2( u0_u11_u2_n177 ) );
  NOR3_X1 u0_u11_u2_U55 (.ZN( u0_u11_u2_n142 ) , .A3( u0_u11_u2_n175 ) , .A2( u0_u11_u2_n178 ) , .A1( u0_u11_u2_n181 ) );
  NAND2_X1 u0_u11_u2_U56 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n113 ) );
  NAND2_X1 u0_u11_u2_U57 (.A1( u0_u11_u2_n106 ) , .A2( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n131 ) );
  NAND2_X1 u0_u11_u2_U58 (.A1( u0_u11_u2_n103 ) , .A2( u0_u11_u2_n107 ) , .ZN( u0_u11_u2_n139 ) );
  NAND2_X1 u0_u11_u2_U59 (.A1( u0_u11_u2_n103 ) , .A2( u0_u11_u2_n105 ) , .ZN( u0_u11_u2_n133 ) );
  NOR4_X1 u0_u11_u2_U6 (.A4( u0_u11_u2_n124 ) , .A3( u0_u11_u2_n125 ) , .A2( u0_u11_u2_n126 ) , .A1( u0_u11_u2_n127 ) , .ZN( u0_u11_u2_n128 ) );
  NAND2_X1 u0_u11_u2_U60 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n103 ) , .ZN( u0_u11_u2_n154 ) );
  NAND2_X1 u0_u11_u2_U61 (.A2( u0_u11_u2_n103 ) , .A1( u0_u11_u2_n104 ) , .ZN( u0_u11_u2_n119 ) );
  NAND2_X1 u0_u11_u2_U62 (.A2( u0_u11_u2_n107 ) , .A1( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n123 ) );
  NAND2_X1 u0_u11_u2_U63 (.A1( u0_u11_u2_n104 ) , .A2( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n122 ) );
  INV_X1 u0_u11_u2_U64 (.A( u0_u11_u2_n114 ) , .ZN( u0_u11_u2_n172 ) );
  NAND2_X1 u0_u11_u2_U65 (.A2( u0_u11_u2_n100 ) , .A1( u0_u11_u2_n102 ) , .ZN( u0_u11_u2_n116 ) );
  NAND2_X1 u0_u11_u2_U66 (.A1( u0_u11_u2_n102 ) , .A2( u0_u11_u2_n108 ) , .ZN( u0_u11_u2_n120 ) );
  NAND2_X1 u0_u11_u2_U67 (.A2( u0_u11_u2_n105 ) , .A1( u0_u11_u2_n106 ) , .ZN( u0_u11_u2_n117 ) );
  INV_X1 u0_u11_u2_U68 (.ZN( u0_u11_u2_n187 ) , .A( u0_u11_u2_n99 ) );
  OAI21_X1 u0_u11_u2_U69 (.B1( u0_u11_u2_n137 ) , .B2( u0_u11_u2_n143 ) , .A( u0_u11_u2_n98 ) , .ZN( u0_u11_u2_n99 ) );
  AOI21_X1 u0_u11_u2_U7 (.ZN( u0_u11_u2_n124 ) , .B1( u0_u11_u2_n131 ) , .B2( u0_u11_u2_n143 ) , .A( u0_u11_u2_n172 ) );
  NOR2_X1 u0_u11_u2_U70 (.A2( u0_u11_X_16 ) , .ZN( u0_u11_u2_n140 ) , .A1( u0_u11_u2_n166 ) );
  NOR2_X1 u0_u11_u2_U71 (.A2( u0_u11_X_13 ) , .A1( u0_u11_X_14 ) , .ZN( u0_u11_u2_n100 ) );
  NOR2_X1 u0_u11_u2_U72 (.A2( u0_u11_X_16 ) , .A1( u0_u11_X_17 ) , .ZN( u0_u11_u2_n138 ) );
  NOR2_X1 u0_u11_u2_U73 (.A2( u0_u11_X_15 ) , .A1( u0_u11_X_18 ) , .ZN( u0_u11_u2_n104 ) );
  NOR2_X1 u0_u11_u2_U74 (.A2( u0_u11_X_14 ) , .ZN( u0_u11_u2_n103 ) , .A1( u0_u11_u2_n174 ) );
  NOR2_X1 u0_u11_u2_U75 (.A2( u0_u11_X_15 ) , .ZN( u0_u11_u2_n102 ) , .A1( u0_u11_u2_n165 ) );
  NOR2_X1 u0_u11_u2_U76 (.A2( u0_u11_X_17 ) , .ZN( u0_u11_u2_n114 ) , .A1( u0_u11_u2_n169 ) );
  AND2_X1 u0_u11_u2_U77 (.A1( u0_u11_X_15 ) , .ZN( u0_u11_u2_n105 ) , .A2( u0_u11_u2_n165 ) );
  AND2_X1 u0_u11_u2_U78 (.A2( u0_u11_X_15 ) , .A1( u0_u11_X_18 ) , .ZN( u0_u11_u2_n107 ) );
  AND2_X1 u0_u11_u2_U79 (.A1( u0_u11_X_14 ) , .ZN( u0_u11_u2_n106 ) , .A2( u0_u11_u2_n174 ) );
  AOI21_X1 u0_u11_u2_U8 (.B2( u0_u11_u2_n119 ) , .ZN( u0_u11_u2_n127 ) , .A( u0_u11_u2_n137 ) , .B1( u0_u11_u2_n155 ) );
  AND2_X1 u0_u11_u2_U80 (.A1( u0_u11_X_13 ) , .A2( u0_u11_X_14 ) , .ZN( u0_u11_u2_n108 ) );
  INV_X1 u0_u11_u2_U81 (.A( u0_u11_X_16 ) , .ZN( u0_u11_u2_n169 ) );
  INV_X1 u0_u11_u2_U82 (.A( u0_u11_X_17 ) , .ZN( u0_u11_u2_n166 ) );
  INV_X1 u0_u11_u2_U83 (.A( u0_u11_X_13 ) , .ZN( u0_u11_u2_n174 ) );
  INV_X1 u0_u11_u2_U84 (.A( u0_u11_X_18 ) , .ZN( u0_u11_u2_n165 ) );
  NAND4_X1 u0_u11_u2_U85 (.ZN( u0_out11_30 ) , .A4( u0_u11_u2_n147 ) , .A3( u0_u11_u2_n148 ) , .A2( u0_u11_u2_n149 ) , .A1( u0_u11_u2_n187 ) );
  NOR3_X1 u0_u11_u2_U86 (.A3( u0_u11_u2_n144 ) , .A2( u0_u11_u2_n145 ) , .A1( u0_u11_u2_n146 ) , .ZN( u0_u11_u2_n147 ) );
  AOI21_X1 u0_u11_u2_U87 (.B2( u0_u11_u2_n138 ) , .ZN( u0_u11_u2_n148 ) , .A( u0_u11_u2_n162 ) , .B1( u0_u11_u2_n182 ) );
  NAND4_X1 u0_u11_u2_U88 (.ZN( u0_out11_24 ) , .A4( u0_u11_u2_n111 ) , .A3( u0_u11_u2_n112 ) , .A1( u0_u11_u2_n130 ) , .A2( u0_u11_u2_n187 ) );
  AOI221_X1 u0_u11_u2_U89 (.A( u0_u11_u2_n109 ) , .B1( u0_u11_u2_n110 ) , .ZN( u0_u11_u2_n111 ) , .C1( u0_u11_u2_n134 ) , .C2( u0_u11_u2_n170 ) , .B2( u0_u11_u2_n173 ) );
  AOI21_X1 u0_u11_u2_U9 (.B2( u0_u11_u2_n123 ) , .ZN( u0_u11_u2_n125 ) , .A( u0_u11_u2_n171 ) , .B1( u0_u11_u2_n184 ) );
  AOI21_X1 u0_u11_u2_U90 (.ZN( u0_u11_u2_n112 ) , .B2( u0_u11_u2_n156 ) , .A( u0_u11_u2_n164 ) , .B1( u0_u11_u2_n181 ) );
  NAND4_X1 u0_u11_u2_U91 (.ZN( u0_out11_16 ) , .A4( u0_u11_u2_n128 ) , .A3( u0_u11_u2_n129 ) , .A1( u0_u11_u2_n130 ) , .A2( u0_u11_u2_n186 ) );
  AOI22_X1 u0_u11_u2_U92 (.A2( u0_u11_u2_n118 ) , .ZN( u0_u11_u2_n129 ) , .A1( u0_u11_u2_n140 ) , .B1( u0_u11_u2_n157 ) , .B2( u0_u11_u2_n170 ) );
  INV_X1 u0_u11_u2_U93 (.A( u0_u11_u2_n163 ) , .ZN( u0_u11_u2_n186 ) );
  OR4_X1 u0_u11_u2_U94 (.ZN( u0_out11_6 ) , .A4( u0_u11_u2_n161 ) , .A3( u0_u11_u2_n162 ) , .A2( u0_u11_u2_n163 ) , .A1( u0_u11_u2_n164 ) );
  OR3_X1 u0_u11_u2_U95 (.A2( u0_u11_u2_n159 ) , .A1( u0_u11_u2_n160 ) , .ZN( u0_u11_u2_n161 ) , .A3( u0_u11_u2_n183 ) );
  AOI21_X1 u0_u11_u2_U96 (.B2( u0_u11_u2_n154 ) , .B1( u0_u11_u2_n155 ) , .ZN( u0_u11_u2_n159 ) , .A( u0_u11_u2_n167 ) );
  NAND3_X1 u0_u11_u2_U97 (.A2( u0_u11_u2_n117 ) , .A1( u0_u11_u2_n122 ) , .A3( u0_u11_u2_n123 ) , .ZN( u0_u11_u2_n134 ) );
  NAND3_X1 u0_u11_u2_U98 (.ZN( u0_u11_u2_n110 ) , .A2( u0_u11_u2_n131 ) , .A3( u0_u11_u2_n139 ) , .A1( u0_u11_u2_n154 ) );
  NAND3_X1 u0_u11_u2_U99 (.A2( u0_u11_u2_n100 ) , .ZN( u0_u11_u2_n101 ) , .A1( u0_u11_u2_n104 ) , .A3( u0_u11_u2_n114 ) );
  OAI21_X1 u0_u11_u6_U10 (.A( u0_u11_u6_n159 ) , .B1( u0_u11_u6_n169 ) , .B2( u0_u11_u6_n173 ) , .ZN( u0_u11_u6_n90 ) );
  INV_X1 u0_u11_u6_U11 (.ZN( u0_u11_u6_n172 ) , .A( u0_u11_u6_n88 ) );
  AOI22_X1 u0_u11_u6_U12 (.A2( u0_u11_u6_n151 ) , .B2( u0_u11_u6_n161 ) , .A1( u0_u11_u6_n167 ) , .B1( u0_u11_u6_n170 ) , .ZN( u0_u11_u6_n89 ) );
  AOI21_X1 u0_u11_u6_U13 (.ZN( u0_u11_u6_n106 ) , .A( u0_u11_u6_n142 ) , .B2( u0_u11_u6_n159 ) , .B1( u0_u11_u6_n164 ) );
  INV_X1 u0_u11_u6_U14 (.A( u0_u11_u6_n155 ) , .ZN( u0_u11_u6_n161 ) );
  INV_X1 u0_u11_u6_U15 (.A( u0_u11_u6_n128 ) , .ZN( u0_u11_u6_n164 ) );
  NAND2_X1 u0_u11_u6_U16 (.ZN( u0_u11_u6_n110 ) , .A1( u0_u11_u6_n122 ) , .A2( u0_u11_u6_n129 ) );
  NAND2_X1 u0_u11_u6_U17 (.ZN( u0_u11_u6_n124 ) , .A2( u0_u11_u6_n146 ) , .A1( u0_u11_u6_n148 ) );
  INV_X1 u0_u11_u6_U18 (.A( u0_u11_u6_n132 ) , .ZN( u0_u11_u6_n171 ) );
  AND2_X1 u0_u11_u6_U19 (.A1( u0_u11_u6_n100 ) , .ZN( u0_u11_u6_n130 ) , .A2( u0_u11_u6_n147 ) );
  INV_X1 u0_u11_u6_U20 (.A( u0_u11_u6_n127 ) , .ZN( u0_u11_u6_n173 ) );
  INV_X1 u0_u11_u6_U21 (.A( u0_u11_u6_n121 ) , .ZN( u0_u11_u6_n167 ) );
  INV_X1 u0_u11_u6_U22 (.A( u0_u11_u6_n100 ) , .ZN( u0_u11_u6_n169 ) );
  INV_X1 u0_u11_u6_U23 (.A( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n170 ) );
  INV_X1 u0_u11_u6_U24 (.A( u0_u11_u6_n113 ) , .ZN( u0_u11_u6_n168 ) );
  AND2_X1 u0_u11_u6_U25 (.A1( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n119 ) , .ZN( u0_u11_u6_n133 ) );
  AND2_X1 u0_u11_u6_U26 (.A2( u0_u11_u6_n121 ) , .A1( u0_u11_u6_n122 ) , .ZN( u0_u11_u6_n131 ) );
  AND3_X1 u0_u11_u6_U27 (.ZN( u0_u11_u6_n120 ) , .A2( u0_u11_u6_n127 ) , .A1( u0_u11_u6_n132 ) , .A3( u0_u11_u6_n145 ) );
  INV_X1 u0_u11_u6_U28 (.A( u0_u11_u6_n146 ) , .ZN( u0_u11_u6_n163 ) );
  AOI222_X1 u0_u11_u6_U29 (.ZN( u0_u11_u6_n114 ) , .A1( u0_u11_u6_n118 ) , .A2( u0_u11_u6_n126 ) , .B2( u0_u11_u6_n151 ) , .C2( u0_u11_u6_n159 ) , .C1( u0_u11_u6_n168 ) , .B1( u0_u11_u6_n169 ) );
  INV_X1 u0_u11_u6_U3 (.A( u0_u11_u6_n110 ) , .ZN( u0_u11_u6_n166 ) );
  NOR2_X1 u0_u11_u6_U30 (.A1( u0_u11_u6_n162 ) , .A2( u0_u11_u6_n165 ) , .ZN( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U31 (.A1( u0_u11_u6_n144 ) , .ZN( u0_u11_u6_n151 ) , .A2( u0_u11_u6_n158 ) );
  NAND2_X1 u0_u11_u6_U32 (.ZN( u0_u11_u6_n132 ) , .A1( u0_u11_u6_n91 ) , .A2( u0_u11_u6_n97 ) );
  AOI22_X1 u0_u11_u6_U33 (.B2( u0_u11_u6_n110 ) , .B1( u0_u11_u6_n111 ) , .A1( u0_u11_u6_n112 ) , .ZN( u0_u11_u6_n115 ) , .A2( u0_u11_u6_n161 ) );
  NAND4_X1 u0_u11_u6_U34 (.A3( u0_u11_u6_n109 ) , .ZN( u0_u11_u6_n112 ) , .A4( u0_u11_u6_n132 ) , .A2( u0_u11_u6_n147 ) , .A1( u0_u11_u6_n166 ) );
  NOR2_X1 u0_u11_u6_U35 (.ZN( u0_u11_u6_n109 ) , .A1( u0_u11_u6_n170 ) , .A2( u0_u11_u6_n173 ) );
  NOR2_X1 u0_u11_u6_U36 (.A2( u0_u11_u6_n126 ) , .ZN( u0_u11_u6_n155 ) , .A1( u0_u11_u6_n160 ) );
  NAND2_X1 u0_u11_u6_U37 (.ZN( u0_u11_u6_n146 ) , .A2( u0_u11_u6_n94 ) , .A1( u0_u11_u6_n99 ) );
  AOI21_X1 u0_u11_u6_U38 (.A( u0_u11_u6_n144 ) , .B2( u0_u11_u6_n145 ) , .B1( u0_u11_u6_n146 ) , .ZN( u0_u11_u6_n150 ) );
  AOI211_X1 u0_u11_u6_U39 (.B( u0_u11_u6_n134 ) , .A( u0_u11_u6_n135 ) , .C1( u0_u11_u6_n136 ) , .ZN( u0_u11_u6_n137 ) , .C2( u0_u11_u6_n151 ) );
  INV_X1 u0_u11_u6_U4 (.A( u0_u11_u6_n142 ) , .ZN( u0_u11_u6_n174 ) );
  NAND4_X1 u0_u11_u6_U40 (.A4( u0_u11_u6_n127 ) , .A3( u0_u11_u6_n128 ) , .A2( u0_u11_u6_n129 ) , .A1( u0_u11_u6_n130 ) , .ZN( u0_u11_u6_n136 ) );
  AOI21_X1 u0_u11_u6_U41 (.B2( u0_u11_u6_n132 ) , .B1( u0_u11_u6_n133 ) , .ZN( u0_u11_u6_n134 ) , .A( u0_u11_u6_n158 ) );
  AOI21_X1 u0_u11_u6_U42 (.B1( u0_u11_u6_n131 ) , .ZN( u0_u11_u6_n135 ) , .A( u0_u11_u6_n144 ) , .B2( u0_u11_u6_n146 ) );
  INV_X1 u0_u11_u6_U43 (.A( u0_u11_u6_n111 ) , .ZN( u0_u11_u6_n158 ) );
  NAND2_X1 u0_u11_u6_U44 (.ZN( u0_u11_u6_n127 ) , .A1( u0_u11_u6_n91 ) , .A2( u0_u11_u6_n92 ) );
  NAND2_X1 u0_u11_u6_U45 (.ZN( u0_u11_u6_n129 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n96 ) );
  INV_X1 u0_u11_u6_U46 (.A( u0_u11_u6_n144 ) , .ZN( u0_u11_u6_n159 ) );
  NAND2_X1 u0_u11_u6_U47 (.ZN( u0_u11_u6_n145 ) , .A2( u0_u11_u6_n97 ) , .A1( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U48 (.ZN( u0_u11_u6_n148 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n94 ) );
  NAND2_X1 u0_u11_u6_U49 (.ZN( u0_u11_u6_n108 ) , .A2( u0_u11_u6_n139 ) , .A1( u0_u11_u6_n144 ) );
  NAND2_X1 u0_u11_u6_U5 (.A2( u0_u11_u6_n143 ) , .ZN( u0_u11_u6_n152 ) , .A1( u0_u11_u6_n166 ) );
  NAND2_X1 u0_u11_u6_U50 (.ZN( u0_u11_u6_n121 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n97 ) );
  NAND2_X1 u0_u11_u6_U51 (.ZN( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n95 ) );
  AND2_X1 u0_u11_u6_U52 (.ZN( u0_u11_u6_n118 ) , .A2( u0_u11_u6_n91 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U53 (.ZN( u0_u11_u6_n147 ) , .A2( u0_u11_u6_n98 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U54 (.ZN( u0_u11_u6_n128 ) , .A1( u0_u11_u6_n94 ) , .A2( u0_u11_u6_n96 ) );
  NAND2_X1 u0_u11_u6_U55 (.ZN( u0_u11_u6_n119 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U56 (.ZN( u0_u11_u6_n123 ) , .A2( u0_u11_u6_n91 ) , .A1( u0_u11_u6_n96 ) );
  NAND2_X1 u0_u11_u6_U57 (.ZN( u0_u11_u6_n100 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U58 (.ZN( u0_u11_u6_n122 ) , .A1( u0_u11_u6_n94 ) , .A2( u0_u11_u6_n97 ) );
  INV_X1 u0_u11_u6_U59 (.A( u0_u11_u6_n139 ) , .ZN( u0_u11_u6_n160 ) );
  AOI22_X1 u0_u11_u6_U6 (.B2( u0_u11_u6_n101 ) , .A1( u0_u11_u6_n102 ) , .ZN( u0_u11_u6_n103 ) , .B1( u0_u11_u6_n160 ) , .A2( u0_u11_u6_n161 ) );
  NAND2_X1 u0_u11_u6_U60 (.ZN( u0_u11_u6_n113 ) , .A1( u0_u11_u6_n96 ) , .A2( u0_u11_u6_n98 ) );
  NOR2_X1 u0_u11_u6_U61 (.A2( u0_u11_X_40 ) , .A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n126 ) );
  NOR2_X1 u0_u11_u6_U62 (.A2( u0_u11_X_39 ) , .A1( u0_u11_X_42 ) , .ZN( u0_u11_u6_n92 ) );
  NOR2_X1 u0_u11_u6_U63 (.A2( u0_u11_X_39 ) , .A1( u0_u11_u6_n156 ) , .ZN( u0_u11_u6_n97 ) );
  NOR2_X1 u0_u11_u6_U64 (.A2( u0_u11_X_38 ) , .A1( u0_u11_u6_n165 ) , .ZN( u0_u11_u6_n95 ) );
  NOR2_X1 u0_u11_u6_U65 (.A2( u0_u11_X_41 ) , .ZN( u0_u11_u6_n111 ) , .A1( u0_u11_u6_n157 ) );
  NOR2_X1 u0_u11_u6_U66 (.A2( u0_u11_X_37 ) , .A1( u0_u11_u6_n162 ) , .ZN( u0_u11_u6_n94 ) );
  NOR2_X1 u0_u11_u6_U67 (.A2( u0_u11_X_37 ) , .A1( u0_u11_X_38 ) , .ZN( u0_u11_u6_n91 ) );
  NAND2_X1 u0_u11_u6_U68 (.A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n144 ) , .A2( u0_u11_u6_n157 ) );
  NAND2_X1 u0_u11_u6_U69 (.A2( u0_u11_X_40 ) , .A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n139 ) );
  NOR2_X1 u0_u11_u6_U7 (.A1( u0_u11_u6_n118 ) , .ZN( u0_u11_u6_n143 ) , .A2( u0_u11_u6_n168 ) );
  AND2_X1 u0_u11_u6_U70 (.A1( u0_u11_X_39 ) , .A2( u0_u11_u6_n156 ) , .ZN( u0_u11_u6_n96 ) );
  AND2_X1 u0_u11_u6_U71 (.A1( u0_u11_X_39 ) , .A2( u0_u11_X_42 ) , .ZN( u0_u11_u6_n99 ) );
  INV_X1 u0_u11_u6_U72 (.A( u0_u11_X_40 ) , .ZN( u0_u11_u6_n157 ) );
  INV_X1 u0_u11_u6_U73 (.A( u0_u11_X_37 ) , .ZN( u0_u11_u6_n165 ) );
  INV_X1 u0_u11_u6_U74 (.A( u0_u11_X_38 ) , .ZN( u0_u11_u6_n162 ) );
  INV_X1 u0_u11_u6_U75 (.A( u0_u11_X_42 ) , .ZN( u0_u11_u6_n156 ) );
  NAND4_X1 u0_u11_u6_U76 (.ZN( u0_out11_32 ) , .A4( u0_u11_u6_n103 ) , .A3( u0_u11_u6_n104 ) , .A2( u0_u11_u6_n105 ) , .A1( u0_u11_u6_n106 ) );
  AOI22_X1 u0_u11_u6_U77 (.ZN( u0_u11_u6_n105 ) , .A2( u0_u11_u6_n108 ) , .A1( u0_u11_u6_n118 ) , .B2( u0_u11_u6_n126 ) , .B1( u0_u11_u6_n171 ) );
  AOI22_X1 u0_u11_u6_U78 (.ZN( u0_u11_u6_n104 ) , .A1( u0_u11_u6_n111 ) , .B1( u0_u11_u6_n124 ) , .B2( u0_u11_u6_n151 ) , .A2( u0_u11_u6_n93 ) );
  NAND4_X1 u0_u11_u6_U79 (.ZN( u0_out11_12 ) , .A4( u0_u11_u6_n114 ) , .A3( u0_u11_u6_n115 ) , .A2( u0_u11_u6_n116 ) , .A1( u0_u11_u6_n117 ) );
  AOI21_X1 u0_u11_u6_U8 (.B1( u0_u11_u6_n107 ) , .B2( u0_u11_u6_n132 ) , .A( u0_u11_u6_n158 ) , .ZN( u0_u11_u6_n88 ) );
  OAI22_X1 u0_u11_u6_U80 (.B2( u0_u11_u6_n111 ) , .ZN( u0_u11_u6_n116 ) , .B1( u0_u11_u6_n126 ) , .A2( u0_u11_u6_n164 ) , .A1( u0_u11_u6_n167 ) );
  OAI21_X1 u0_u11_u6_U81 (.A( u0_u11_u6_n108 ) , .ZN( u0_u11_u6_n117 ) , .B2( u0_u11_u6_n141 ) , .B1( u0_u11_u6_n163 ) );
  OAI211_X1 u0_u11_u6_U82 (.ZN( u0_out11_7 ) , .B( u0_u11_u6_n153 ) , .C2( u0_u11_u6_n154 ) , .C1( u0_u11_u6_n155 ) , .A( u0_u11_u6_n174 ) );
  NOR3_X1 u0_u11_u6_U83 (.A1( u0_u11_u6_n141 ) , .ZN( u0_u11_u6_n154 ) , .A3( u0_u11_u6_n164 ) , .A2( u0_u11_u6_n171 ) );
  AOI211_X1 u0_u11_u6_U84 (.B( u0_u11_u6_n149 ) , .A( u0_u11_u6_n150 ) , .C2( u0_u11_u6_n151 ) , .C1( u0_u11_u6_n152 ) , .ZN( u0_u11_u6_n153 ) );
  OAI211_X1 u0_u11_u6_U85 (.ZN( u0_out11_22 ) , .B( u0_u11_u6_n137 ) , .A( u0_u11_u6_n138 ) , .C2( u0_u11_u6_n139 ) , .C1( u0_u11_u6_n140 ) );
  AOI22_X1 u0_u11_u6_U86 (.B1( u0_u11_u6_n124 ) , .A2( u0_u11_u6_n125 ) , .A1( u0_u11_u6_n126 ) , .ZN( u0_u11_u6_n138 ) , .B2( u0_u11_u6_n161 ) );
  AND4_X1 u0_u11_u6_U87 (.A3( u0_u11_u6_n119 ) , .A1( u0_u11_u6_n120 ) , .A4( u0_u11_u6_n129 ) , .ZN( u0_u11_u6_n140 ) , .A2( u0_u11_u6_n143 ) );
  NAND3_X1 u0_u11_u6_U88 (.A2( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n125 ) , .A1( u0_u11_u6_n130 ) , .A3( u0_u11_u6_n131 ) );
  NAND3_X1 u0_u11_u6_U89 (.A3( u0_u11_u6_n133 ) , .ZN( u0_u11_u6_n141 ) , .A1( u0_u11_u6_n145 ) , .A2( u0_u11_u6_n148 ) );
  AOI21_X1 u0_u11_u6_U9 (.B2( u0_u11_u6_n147 ) , .B1( u0_u11_u6_n148 ) , .ZN( u0_u11_u6_n149 ) , .A( u0_u11_u6_n158 ) );
  NAND3_X1 u0_u11_u6_U90 (.ZN( u0_u11_u6_n101 ) , .A3( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n121 ) , .A1( u0_u11_u6_n127 ) );
  NAND3_X1 u0_u11_u6_U91 (.ZN( u0_u11_u6_n102 ) , .A3( u0_u11_u6_n130 ) , .A2( u0_u11_u6_n145 ) , .A1( u0_u11_u6_n166 ) );
  NAND3_X1 u0_u11_u6_U92 (.A3( u0_u11_u6_n113 ) , .A1( u0_u11_u6_n119 ) , .A2( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n93 ) );
  NAND3_X1 u0_u11_u6_U93 (.ZN( u0_u11_u6_n142 ) , .A2( u0_u11_u6_n172 ) , .A3( u0_u11_u6_n89 ) , .A1( u0_u11_u6_n90 ) );
  XOR2_X1 u0_u15_U26 (.A( u0_FP_53 ) , .B( u0_K16_30 ) , .Z( u0_u15_X_30 ) );
  XOR2_X1 u0_u15_U28 (.A( u0_FP_52 ) , .B( u0_K16_29 ) , .Z( u0_u15_X_29 ) );
  XOR2_X1 u0_u15_U29 (.A( u0_FP_51 ) , .B( u0_K16_28 ) , .Z( u0_u15_X_28 ) );
  XOR2_X1 u0_u15_U30 (.A( u0_FP_50 ) , .B( u0_K16_27 ) , .Z( u0_u15_X_27 ) );
  XOR2_X1 u0_u15_U31 (.A( u0_FP_49 ) , .B( u0_K16_26 ) , .Z( u0_u15_X_26 ) );
  XOR2_X1 u0_u15_U32 (.A( u0_FP_48 ) , .B( u0_K16_25 ) , .Z( u0_u15_X_25 ) );
  XOR2_X1 u0_u15_U33 (.A( u0_FP_49 ) , .B( u0_K16_24 ) , .Z( u0_u15_X_24 ) );
  XOR2_X1 u0_u15_U34 (.A( u0_FP_48 ) , .B( u0_K16_23 ) , .Z( u0_u15_X_23 ) );
  XOR2_X1 u0_u15_U35 (.A( u0_FP_47 ) , .B( u0_K16_22 ) , .Z( u0_u15_X_22 ) );
  XOR2_X1 u0_u15_U36 (.A( u0_FP_46 ) , .B( u0_K16_21 ) , .Z( u0_u15_X_21 ) );
  XOR2_X1 u0_u15_U37 (.A( u0_FP_45 ) , .B( u0_K16_20 ) , .Z( u0_u15_X_20 ) );
  XOR2_X1 u0_u15_U39 (.A( u0_FP_44 ) , .B( u0_K16_19 ) , .Z( u0_u15_X_19 ) );
  XOR2_X1 u0_u15_U40 (.A( u0_FP_45 ) , .B( u0_K16_18 ) , .Z( u0_u15_X_18 ) );
  XOR2_X1 u0_u15_U41 (.A( u0_FP_44 ) , .B( u0_K16_17 ) , .Z( u0_u15_X_17 ) );
  XOR2_X1 u0_u15_U42 (.A( u0_FP_43 ) , .B( u0_K16_16 ) , .Z( u0_u15_X_16 ) );
  XOR2_X1 u0_u15_U43 (.A( u0_FP_42 ) , .B( u0_K16_15 ) , .Z( u0_u15_X_15 ) );
  XOR2_X1 u0_u15_U44 (.A( u0_FP_41 ) , .B( u0_K16_14 ) , .Z( u0_u15_X_14 ) );
  XOR2_X1 u0_u15_U45 (.A( u0_FP_40 ) , .B( u0_K16_13 ) , .Z( u0_u15_X_13 ) );
  OAI22_X1 u0_u15_u2_U10 (.B1( u0_u15_u2_n151 ) , .A2( u0_u15_u2_n152 ) , .A1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n160 ) , .B2( u0_u15_u2_n168 ) );
  NAND3_X1 u0_u15_u2_U100 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n98 ) );
  NOR3_X1 u0_u15_u2_U11 (.A1( u0_u15_u2_n150 ) , .ZN( u0_u15_u2_n151 ) , .A3( u0_u15_u2_n175 ) , .A2( u0_u15_u2_n188 ) );
  AOI21_X1 u0_u15_u2_U12 (.B2( u0_u15_u2_n123 ) , .ZN( u0_u15_u2_n125 ) , .A( u0_u15_u2_n171 ) , .B1( u0_u15_u2_n184 ) );
  INV_X1 u0_u15_u2_U13 (.A( u0_u15_u2_n150 ) , .ZN( u0_u15_u2_n184 ) );
  AOI21_X1 u0_u15_u2_U14 (.ZN( u0_u15_u2_n144 ) , .B2( u0_u15_u2_n155 ) , .A( u0_u15_u2_n172 ) , .B1( u0_u15_u2_n185 ) );
  AOI21_X1 u0_u15_u2_U15 (.B2( u0_u15_u2_n143 ) , .ZN( u0_u15_u2_n145 ) , .B1( u0_u15_u2_n152 ) , .A( u0_u15_u2_n171 ) );
  INV_X1 u0_u15_u2_U16 (.A( u0_u15_u2_n156 ) , .ZN( u0_u15_u2_n171 ) );
  INV_X1 u0_u15_u2_U17 (.A( u0_u15_u2_n120 ) , .ZN( u0_u15_u2_n188 ) );
  NAND2_X1 u0_u15_u2_U18 (.A2( u0_u15_u2_n122 ) , .ZN( u0_u15_u2_n150 ) , .A1( u0_u15_u2_n152 ) );
  INV_X1 u0_u15_u2_U19 (.A( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n170 ) );
  INV_X1 u0_u15_u2_U20 (.A( u0_u15_u2_n137 ) , .ZN( u0_u15_u2_n173 ) );
  NAND2_X1 u0_u15_u2_U21 (.A1( u0_u15_u2_n132 ) , .A2( u0_u15_u2_n139 ) , .ZN( u0_u15_u2_n157 ) );
  INV_X1 u0_u15_u2_U22 (.A( u0_u15_u2_n113 ) , .ZN( u0_u15_u2_n178 ) );
  INV_X1 u0_u15_u2_U23 (.A( u0_u15_u2_n139 ) , .ZN( u0_u15_u2_n175 ) );
  INV_X1 u0_u15_u2_U24 (.A( u0_u15_u2_n155 ) , .ZN( u0_u15_u2_n181 ) );
  INV_X1 u0_u15_u2_U25 (.A( u0_u15_u2_n119 ) , .ZN( u0_u15_u2_n177 ) );
  INV_X1 u0_u15_u2_U26 (.A( u0_u15_u2_n116 ) , .ZN( u0_u15_u2_n180 ) );
  INV_X1 u0_u15_u2_U27 (.A( u0_u15_u2_n131 ) , .ZN( u0_u15_u2_n179 ) );
  INV_X1 u0_u15_u2_U28 (.A( u0_u15_u2_n154 ) , .ZN( u0_u15_u2_n176 ) );
  NAND2_X1 u0_u15_u2_U29 (.A2( u0_u15_u2_n116 ) , .A1( u0_u15_u2_n117 ) , .ZN( u0_u15_u2_n118 ) );
  NOR2_X1 u0_u15_u2_U3 (.ZN( u0_u15_u2_n121 ) , .A2( u0_u15_u2_n177 ) , .A1( u0_u15_u2_n180 ) );
  INV_X1 u0_u15_u2_U30 (.A( u0_u15_u2_n132 ) , .ZN( u0_u15_u2_n182 ) );
  INV_X1 u0_u15_u2_U31 (.A( u0_u15_u2_n158 ) , .ZN( u0_u15_u2_n183 ) );
  OAI21_X1 u0_u15_u2_U32 (.A( u0_u15_u2_n156 ) , .B1( u0_u15_u2_n157 ) , .ZN( u0_u15_u2_n158 ) , .B2( u0_u15_u2_n179 ) );
  NOR2_X1 u0_u15_u2_U33 (.ZN( u0_u15_u2_n156 ) , .A1( u0_u15_u2_n166 ) , .A2( u0_u15_u2_n169 ) );
  NOR2_X1 u0_u15_u2_U34 (.A2( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n137 ) , .A1( u0_u15_u2_n140 ) );
  NOR2_X1 u0_u15_u2_U35 (.A2( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n153 ) , .A1( u0_u15_u2_n156 ) );
  AOI211_X1 u0_u15_u2_U36 (.ZN( u0_u15_u2_n130 ) , .C1( u0_u15_u2_n138 ) , .C2( u0_u15_u2_n179 ) , .B( u0_u15_u2_n96 ) , .A( u0_u15_u2_n97 ) );
  OAI22_X1 u0_u15_u2_U37 (.B1( u0_u15_u2_n133 ) , .A2( u0_u15_u2_n137 ) , .A1( u0_u15_u2_n152 ) , .B2( u0_u15_u2_n168 ) , .ZN( u0_u15_u2_n97 ) );
  OAI221_X1 u0_u15_u2_U38 (.B1( u0_u15_u2_n113 ) , .C1( u0_u15_u2_n132 ) , .A( u0_u15_u2_n149 ) , .B2( u0_u15_u2_n171 ) , .C2( u0_u15_u2_n172 ) , .ZN( u0_u15_u2_n96 ) );
  OAI221_X1 u0_u15_u2_U39 (.A( u0_u15_u2_n115 ) , .C2( u0_u15_u2_n123 ) , .B2( u0_u15_u2_n143 ) , .B1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n163 ) , .C1( u0_u15_u2_n168 ) );
  INV_X1 u0_u15_u2_U4 (.A( u0_u15_u2_n134 ) , .ZN( u0_u15_u2_n185 ) );
  OAI21_X1 u0_u15_u2_U40 (.A( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n115 ) , .B1( u0_u15_u2_n176 ) , .B2( u0_u15_u2_n178 ) );
  OAI221_X1 u0_u15_u2_U41 (.A( u0_u15_u2_n135 ) , .B2( u0_u15_u2_n136 ) , .B1( u0_u15_u2_n137 ) , .ZN( u0_u15_u2_n162 ) , .C2( u0_u15_u2_n167 ) , .C1( u0_u15_u2_n185 ) );
  AND3_X1 u0_u15_u2_U42 (.A3( u0_u15_u2_n131 ) , .A2( u0_u15_u2_n132 ) , .A1( u0_u15_u2_n133 ) , .ZN( u0_u15_u2_n136 ) );
  AOI22_X1 u0_u15_u2_U43 (.ZN( u0_u15_u2_n135 ) , .B1( u0_u15_u2_n140 ) , .A1( u0_u15_u2_n156 ) , .B2( u0_u15_u2_n180 ) , .A2( u0_u15_u2_n188 ) );
  AOI21_X1 u0_u15_u2_U44 (.ZN( u0_u15_u2_n149 ) , .B1( u0_u15_u2_n173 ) , .B2( u0_u15_u2_n188 ) , .A( u0_u15_u2_n95 ) );
  AND3_X1 u0_u15_u2_U45 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n156 ) , .ZN( u0_u15_u2_n95 ) );
  OAI21_X1 u0_u15_u2_U46 (.A( u0_u15_u2_n141 ) , .B2( u0_u15_u2_n142 ) , .ZN( u0_u15_u2_n146 ) , .B1( u0_u15_u2_n153 ) );
  OAI21_X1 u0_u15_u2_U47 (.A( u0_u15_u2_n140 ) , .ZN( u0_u15_u2_n141 ) , .B1( u0_u15_u2_n176 ) , .B2( u0_u15_u2_n177 ) );
  NOR3_X1 u0_u15_u2_U48 (.ZN( u0_u15_u2_n142 ) , .A3( u0_u15_u2_n175 ) , .A2( u0_u15_u2_n178 ) , .A1( u0_u15_u2_n181 ) );
  OAI21_X1 u0_u15_u2_U49 (.A( u0_u15_u2_n101 ) , .B2( u0_u15_u2_n121 ) , .B1( u0_u15_u2_n153 ) , .ZN( u0_u15_u2_n164 ) );
  NOR4_X1 u0_u15_u2_U5 (.A4( u0_u15_u2_n124 ) , .A3( u0_u15_u2_n125 ) , .A2( u0_u15_u2_n126 ) , .A1( u0_u15_u2_n127 ) , .ZN( u0_u15_u2_n128 ) );
  NAND2_X1 u0_u15_u2_U50 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n155 ) );
  NAND2_X1 u0_u15_u2_U51 (.A2( u0_u15_u2_n105 ) , .A1( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n143 ) );
  NAND2_X1 u0_u15_u2_U52 (.A1( u0_u15_u2_n104 ) , .A2( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n152 ) );
  NAND2_X1 u0_u15_u2_U53 (.A1( u0_u15_u2_n100 ) , .A2( u0_u15_u2_n105 ) , .ZN( u0_u15_u2_n132 ) );
  INV_X1 u0_u15_u2_U54 (.A( u0_u15_u2_n140 ) , .ZN( u0_u15_u2_n168 ) );
  INV_X1 u0_u15_u2_U55 (.A( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n167 ) );
  INV_X1 u0_u15_u2_U56 (.ZN( u0_u15_u2_n187 ) , .A( u0_u15_u2_n99 ) );
  OAI21_X1 u0_u15_u2_U57 (.B1( u0_u15_u2_n137 ) , .B2( u0_u15_u2_n143 ) , .A( u0_u15_u2_n98 ) , .ZN( u0_u15_u2_n99 ) );
  NAND2_X1 u0_u15_u2_U58 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n113 ) );
  NAND2_X1 u0_u15_u2_U59 (.A1( u0_u15_u2_n106 ) , .A2( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n131 ) );
  AOI21_X1 u0_u15_u2_U6 (.B2( u0_u15_u2_n119 ) , .ZN( u0_u15_u2_n127 ) , .A( u0_u15_u2_n137 ) , .B1( u0_u15_u2_n155 ) );
  NAND2_X1 u0_u15_u2_U60 (.A1( u0_u15_u2_n103 ) , .A2( u0_u15_u2_n107 ) , .ZN( u0_u15_u2_n139 ) );
  NAND2_X1 u0_u15_u2_U61 (.A1( u0_u15_u2_n103 ) , .A2( u0_u15_u2_n105 ) , .ZN( u0_u15_u2_n133 ) );
  NAND2_X1 u0_u15_u2_U62 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n103 ) , .ZN( u0_u15_u2_n154 ) );
  NAND2_X1 u0_u15_u2_U63 (.A2( u0_u15_u2_n103 ) , .A1( u0_u15_u2_n104 ) , .ZN( u0_u15_u2_n119 ) );
  NAND2_X1 u0_u15_u2_U64 (.A2( u0_u15_u2_n107 ) , .A1( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n123 ) );
  NAND2_X1 u0_u15_u2_U65 (.A1( u0_u15_u2_n104 ) , .A2( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n122 ) );
  INV_X1 u0_u15_u2_U66 (.A( u0_u15_u2_n114 ) , .ZN( u0_u15_u2_n172 ) );
  NAND2_X1 u0_u15_u2_U67 (.A2( u0_u15_u2_n100 ) , .A1( u0_u15_u2_n102 ) , .ZN( u0_u15_u2_n116 ) );
  NAND2_X1 u0_u15_u2_U68 (.A1( u0_u15_u2_n102 ) , .A2( u0_u15_u2_n108 ) , .ZN( u0_u15_u2_n120 ) );
  NAND2_X1 u0_u15_u2_U69 (.A2( u0_u15_u2_n105 ) , .A1( u0_u15_u2_n106 ) , .ZN( u0_u15_u2_n117 ) );
  AOI21_X1 u0_u15_u2_U7 (.ZN( u0_u15_u2_n124 ) , .B1( u0_u15_u2_n131 ) , .B2( u0_u15_u2_n143 ) , .A( u0_u15_u2_n172 ) );
  NOR2_X1 u0_u15_u2_U70 (.A2( u0_u15_X_16 ) , .ZN( u0_u15_u2_n140 ) , .A1( u0_u15_u2_n166 ) );
  NOR2_X1 u0_u15_u2_U71 (.A2( u0_u15_X_13 ) , .A1( u0_u15_X_14 ) , .ZN( u0_u15_u2_n100 ) );
  NOR2_X1 u0_u15_u2_U72 (.A2( u0_u15_X_16 ) , .A1( u0_u15_X_17 ) , .ZN( u0_u15_u2_n138 ) );
  NOR2_X1 u0_u15_u2_U73 (.A2( u0_u15_X_15 ) , .A1( u0_u15_X_18 ) , .ZN( u0_u15_u2_n104 ) );
  NOR2_X1 u0_u15_u2_U74 (.A2( u0_u15_X_14 ) , .ZN( u0_u15_u2_n103 ) , .A1( u0_u15_u2_n174 ) );
  NOR2_X1 u0_u15_u2_U75 (.A2( u0_u15_X_15 ) , .ZN( u0_u15_u2_n102 ) , .A1( u0_u15_u2_n165 ) );
  NOR2_X1 u0_u15_u2_U76 (.A2( u0_u15_X_17 ) , .ZN( u0_u15_u2_n114 ) , .A1( u0_u15_u2_n169 ) );
  AND2_X1 u0_u15_u2_U77 (.A1( u0_u15_X_15 ) , .ZN( u0_u15_u2_n105 ) , .A2( u0_u15_u2_n165 ) );
  AND2_X1 u0_u15_u2_U78 (.A2( u0_u15_X_15 ) , .A1( u0_u15_X_18 ) , .ZN( u0_u15_u2_n107 ) );
  AND2_X1 u0_u15_u2_U79 (.A1( u0_u15_X_14 ) , .ZN( u0_u15_u2_n106 ) , .A2( u0_u15_u2_n174 ) );
  AOI21_X1 u0_u15_u2_U8 (.B2( u0_u15_u2_n120 ) , .B1( u0_u15_u2_n121 ) , .ZN( u0_u15_u2_n126 ) , .A( u0_u15_u2_n167 ) );
  AND2_X1 u0_u15_u2_U80 (.A1( u0_u15_X_13 ) , .A2( u0_u15_X_14 ) , .ZN( u0_u15_u2_n108 ) );
  INV_X1 u0_u15_u2_U81 (.A( u0_u15_X_16 ) , .ZN( u0_u15_u2_n169 ) );
  INV_X1 u0_u15_u2_U82 (.A( u0_u15_X_17 ) , .ZN( u0_u15_u2_n166 ) );
  INV_X1 u0_u15_u2_U83 (.A( u0_u15_X_13 ) , .ZN( u0_u15_u2_n174 ) );
  INV_X1 u0_u15_u2_U84 (.A( u0_u15_X_18 ) , .ZN( u0_u15_u2_n165 ) );
  NAND4_X1 u0_u15_u2_U85 (.ZN( u0_out15_30 ) , .A4( u0_u15_u2_n147 ) , .A3( u0_u15_u2_n148 ) , .A2( u0_u15_u2_n149 ) , .A1( u0_u15_u2_n187 ) );
  NOR3_X1 u0_u15_u2_U86 (.A3( u0_u15_u2_n144 ) , .A2( u0_u15_u2_n145 ) , .A1( u0_u15_u2_n146 ) , .ZN( u0_u15_u2_n147 ) );
  AOI21_X1 u0_u15_u2_U87 (.B2( u0_u15_u2_n138 ) , .ZN( u0_u15_u2_n148 ) , .A( u0_u15_u2_n162 ) , .B1( u0_u15_u2_n182 ) );
  NAND4_X1 u0_u15_u2_U88 (.ZN( u0_out15_24 ) , .A4( u0_u15_u2_n111 ) , .A3( u0_u15_u2_n112 ) , .A1( u0_u15_u2_n130 ) , .A2( u0_u15_u2_n187 ) );
  AOI221_X1 u0_u15_u2_U89 (.A( u0_u15_u2_n109 ) , .B1( u0_u15_u2_n110 ) , .ZN( u0_u15_u2_n111 ) , .C1( u0_u15_u2_n134 ) , .C2( u0_u15_u2_n170 ) , .B2( u0_u15_u2_n173 ) );
  OAI22_X1 u0_u15_u2_U9 (.ZN( u0_u15_u2_n109 ) , .A2( u0_u15_u2_n113 ) , .B2( u0_u15_u2_n133 ) , .B1( u0_u15_u2_n167 ) , .A1( u0_u15_u2_n168 ) );
  AOI21_X1 u0_u15_u2_U90 (.ZN( u0_u15_u2_n112 ) , .B2( u0_u15_u2_n156 ) , .A( u0_u15_u2_n164 ) , .B1( u0_u15_u2_n181 ) );
  NAND4_X1 u0_u15_u2_U91 (.ZN( u0_out15_16 ) , .A4( u0_u15_u2_n128 ) , .A3( u0_u15_u2_n129 ) , .A1( u0_u15_u2_n130 ) , .A2( u0_u15_u2_n186 ) );
  AOI22_X1 u0_u15_u2_U92 (.A2( u0_u15_u2_n118 ) , .ZN( u0_u15_u2_n129 ) , .A1( u0_u15_u2_n140 ) , .B1( u0_u15_u2_n157 ) , .B2( u0_u15_u2_n170 ) );
  INV_X1 u0_u15_u2_U93 (.A( u0_u15_u2_n163 ) , .ZN( u0_u15_u2_n186 ) );
  OR4_X1 u0_u15_u2_U94 (.ZN( u0_out15_6 ) , .A4( u0_u15_u2_n161 ) , .A3( u0_u15_u2_n162 ) , .A2( u0_u15_u2_n163 ) , .A1( u0_u15_u2_n164 ) );
  OR3_X1 u0_u15_u2_U95 (.A2( u0_u15_u2_n159 ) , .A1( u0_u15_u2_n160 ) , .ZN( u0_u15_u2_n161 ) , .A3( u0_u15_u2_n183 ) );
  AOI21_X1 u0_u15_u2_U96 (.B2( u0_u15_u2_n154 ) , .B1( u0_u15_u2_n155 ) , .ZN( u0_u15_u2_n159 ) , .A( u0_u15_u2_n167 ) );
  NAND3_X1 u0_u15_u2_U97 (.A2( u0_u15_u2_n117 ) , .A1( u0_u15_u2_n122 ) , .A3( u0_u15_u2_n123 ) , .ZN( u0_u15_u2_n134 ) );
  NAND3_X1 u0_u15_u2_U98 (.ZN( u0_u15_u2_n110 ) , .A2( u0_u15_u2_n131 ) , .A3( u0_u15_u2_n139 ) , .A1( u0_u15_u2_n154 ) );
  NAND3_X1 u0_u15_u2_U99 (.A2( u0_u15_u2_n100 ) , .ZN( u0_u15_u2_n101 ) , .A1( u0_u15_u2_n104 ) , .A3( u0_u15_u2_n114 ) );
  OAI22_X1 u0_u15_u3_U10 (.B1( u0_u15_u3_n113 ) , .A2( u0_u15_u3_n135 ) , .A1( u0_u15_u3_n150 ) , .B2( u0_u15_u3_n164 ) , .ZN( u0_u15_u3_n98 ) );
  OAI211_X1 u0_u15_u3_U11 (.B( u0_u15_u3_n106 ) , .ZN( u0_u15_u3_n119 ) , .C2( u0_u15_u3_n128 ) , .C1( u0_u15_u3_n167 ) , .A( u0_u15_u3_n181 ) );
  AOI221_X1 u0_u15_u3_U12 (.C1( u0_u15_u3_n105 ) , .ZN( u0_u15_u3_n106 ) , .A( u0_u15_u3_n131 ) , .B2( u0_u15_u3_n132 ) , .C2( u0_u15_u3_n133 ) , .B1( u0_u15_u3_n169 ) );
  INV_X1 u0_u15_u3_U13 (.ZN( u0_u15_u3_n181 ) , .A( u0_u15_u3_n98 ) );
  NAND2_X1 u0_u15_u3_U14 (.ZN( u0_u15_u3_n105 ) , .A2( u0_u15_u3_n130 ) , .A1( u0_u15_u3_n155 ) );
  AOI22_X1 u0_u15_u3_U15 (.B1( u0_u15_u3_n115 ) , .A2( u0_u15_u3_n116 ) , .ZN( u0_u15_u3_n123 ) , .B2( u0_u15_u3_n133 ) , .A1( u0_u15_u3_n169 ) );
  NAND2_X1 u0_u15_u3_U16 (.ZN( u0_u15_u3_n116 ) , .A2( u0_u15_u3_n151 ) , .A1( u0_u15_u3_n182 ) );
  NOR2_X1 u0_u15_u3_U17 (.ZN( u0_u15_u3_n126 ) , .A2( u0_u15_u3_n150 ) , .A1( u0_u15_u3_n164 ) );
  AOI21_X1 u0_u15_u3_U18 (.ZN( u0_u15_u3_n112 ) , .B2( u0_u15_u3_n146 ) , .B1( u0_u15_u3_n155 ) , .A( u0_u15_u3_n167 ) );
  NAND2_X1 u0_u15_u3_U19 (.A1( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n142 ) , .A2( u0_u15_u3_n164 ) );
  NAND2_X1 u0_u15_u3_U20 (.ZN( u0_u15_u3_n132 ) , .A2( u0_u15_u3_n152 ) , .A1( u0_u15_u3_n156 ) );
  AND2_X1 u0_u15_u3_U21 (.A2( u0_u15_u3_n113 ) , .A1( u0_u15_u3_n114 ) , .ZN( u0_u15_u3_n151 ) );
  INV_X1 u0_u15_u3_U22 (.A( u0_u15_u3_n133 ) , .ZN( u0_u15_u3_n165 ) );
  INV_X1 u0_u15_u3_U23 (.A( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n170 ) );
  NAND2_X1 u0_u15_u3_U24 (.A1( u0_u15_u3_n107 ) , .A2( u0_u15_u3_n108 ) , .ZN( u0_u15_u3_n140 ) );
  NAND2_X1 u0_u15_u3_U25 (.ZN( u0_u15_u3_n117 ) , .A1( u0_u15_u3_n124 ) , .A2( u0_u15_u3_n148 ) );
  NAND2_X1 u0_u15_u3_U26 (.ZN( u0_u15_u3_n143 ) , .A1( u0_u15_u3_n165 ) , .A2( u0_u15_u3_n167 ) );
  INV_X1 u0_u15_u3_U27 (.A( u0_u15_u3_n130 ) , .ZN( u0_u15_u3_n177 ) );
  INV_X1 u0_u15_u3_U28 (.A( u0_u15_u3_n128 ) , .ZN( u0_u15_u3_n176 ) );
  INV_X1 u0_u15_u3_U29 (.A( u0_u15_u3_n155 ) , .ZN( u0_u15_u3_n174 ) );
  INV_X1 u0_u15_u3_U3 (.A( u0_u15_u3_n129 ) , .ZN( u0_u15_u3_n183 ) );
  INV_X1 u0_u15_u3_U30 (.A( u0_u15_u3_n139 ) , .ZN( u0_u15_u3_n185 ) );
  NOR2_X1 u0_u15_u3_U31 (.ZN( u0_u15_u3_n135 ) , .A2( u0_u15_u3_n141 ) , .A1( u0_u15_u3_n169 ) );
  OAI222_X1 u0_u15_u3_U32 (.C2( u0_u15_u3_n107 ) , .A2( u0_u15_u3_n108 ) , .B1( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n138 ) , .B2( u0_u15_u3_n146 ) , .C1( u0_u15_u3_n154 ) , .A1( u0_u15_u3_n164 ) );
  NOR4_X1 u0_u15_u3_U33 (.A4( u0_u15_u3_n157 ) , .A3( u0_u15_u3_n158 ) , .A2( u0_u15_u3_n159 ) , .A1( u0_u15_u3_n160 ) , .ZN( u0_u15_u3_n161 ) );
  AOI21_X1 u0_u15_u3_U34 (.B2( u0_u15_u3_n152 ) , .B1( u0_u15_u3_n153 ) , .ZN( u0_u15_u3_n158 ) , .A( u0_u15_u3_n164 ) );
  AOI21_X1 u0_u15_u3_U35 (.A( u0_u15_u3_n154 ) , .B2( u0_u15_u3_n155 ) , .B1( u0_u15_u3_n156 ) , .ZN( u0_u15_u3_n157 ) );
  AOI21_X1 u0_u15_u3_U36 (.A( u0_u15_u3_n149 ) , .B2( u0_u15_u3_n150 ) , .B1( u0_u15_u3_n151 ) , .ZN( u0_u15_u3_n159 ) );
  AOI211_X1 u0_u15_u3_U37 (.ZN( u0_u15_u3_n109 ) , .A( u0_u15_u3_n119 ) , .C2( u0_u15_u3_n129 ) , .B( u0_u15_u3_n138 ) , .C1( u0_u15_u3_n141 ) );
  AOI211_X1 u0_u15_u3_U38 (.B( u0_u15_u3_n119 ) , .A( u0_u15_u3_n120 ) , .C2( u0_u15_u3_n121 ) , .ZN( u0_u15_u3_n122 ) , .C1( u0_u15_u3_n179 ) );
  INV_X1 u0_u15_u3_U39 (.A( u0_u15_u3_n156 ) , .ZN( u0_u15_u3_n179 ) );
  INV_X1 u0_u15_u3_U4 (.A( u0_u15_u3_n140 ) , .ZN( u0_u15_u3_n182 ) );
  OAI22_X1 u0_u15_u3_U40 (.B1( u0_u15_u3_n118 ) , .ZN( u0_u15_u3_n120 ) , .A1( u0_u15_u3_n135 ) , .B2( u0_u15_u3_n154 ) , .A2( u0_u15_u3_n178 ) );
  AND3_X1 u0_u15_u3_U41 (.ZN( u0_u15_u3_n118 ) , .A2( u0_u15_u3_n124 ) , .A1( u0_u15_u3_n144 ) , .A3( u0_u15_u3_n152 ) );
  INV_X1 u0_u15_u3_U42 (.A( u0_u15_u3_n121 ) , .ZN( u0_u15_u3_n164 ) );
  NAND2_X1 u0_u15_u3_U43 (.ZN( u0_u15_u3_n133 ) , .A1( u0_u15_u3_n154 ) , .A2( u0_u15_u3_n164 ) );
  OAI211_X1 u0_u15_u3_U44 (.B( u0_u15_u3_n127 ) , .ZN( u0_u15_u3_n139 ) , .C1( u0_u15_u3_n150 ) , .C2( u0_u15_u3_n154 ) , .A( u0_u15_u3_n184 ) );
  INV_X1 u0_u15_u3_U45 (.A( u0_u15_u3_n125 ) , .ZN( u0_u15_u3_n184 ) );
  AOI221_X1 u0_u15_u3_U46 (.A( u0_u15_u3_n126 ) , .ZN( u0_u15_u3_n127 ) , .C2( u0_u15_u3_n132 ) , .C1( u0_u15_u3_n169 ) , .B2( u0_u15_u3_n170 ) , .B1( u0_u15_u3_n174 ) );
  OAI22_X1 u0_u15_u3_U47 (.A1( u0_u15_u3_n124 ) , .ZN( u0_u15_u3_n125 ) , .B2( u0_u15_u3_n145 ) , .A2( u0_u15_u3_n165 ) , .B1( u0_u15_u3_n167 ) );
  NOR2_X1 u0_u15_u3_U48 (.A1( u0_u15_u3_n113 ) , .ZN( u0_u15_u3_n131 ) , .A2( u0_u15_u3_n154 ) );
  NAND2_X1 u0_u15_u3_U49 (.A1( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n150 ) , .A2( u0_u15_u3_n99 ) );
  INV_X1 u0_u15_u3_U5 (.A( u0_u15_u3_n117 ) , .ZN( u0_u15_u3_n178 ) );
  NAND2_X1 u0_u15_u3_U50 (.A2( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n155 ) , .A1( u0_u15_u3_n97 ) );
  INV_X1 u0_u15_u3_U51 (.A( u0_u15_u3_n141 ) , .ZN( u0_u15_u3_n167 ) );
  AOI21_X1 u0_u15_u3_U52 (.B2( u0_u15_u3_n114 ) , .B1( u0_u15_u3_n146 ) , .A( u0_u15_u3_n154 ) , .ZN( u0_u15_u3_n94 ) );
  AOI21_X1 u0_u15_u3_U53 (.ZN( u0_u15_u3_n110 ) , .B2( u0_u15_u3_n142 ) , .B1( u0_u15_u3_n186 ) , .A( u0_u15_u3_n95 ) );
  INV_X1 u0_u15_u3_U54 (.A( u0_u15_u3_n145 ) , .ZN( u0_u15_u3_n186 ) );
  AOI21_X1 u0_u15_u3_U55 (.B1( u0_u15_u3_n124 ) , .A( u0_u15_u3_n149 ) , .B2( u0_u15_u3_n155 ) , .ZN( u0_u15_u3_n95 ) );
  INV_X1 u0_u15_u3_U56 (.A( u0_u15_u3_n149 ) , .ZN( u0_u15_u3_n169 ) );
  NAND2_X1 u0_u15_u3_U57 (.ZN( u0_u15_u3_n124 ) , .A1( u0_u15_u3_n96 ) , .A2( u0_u15_u3_n97 ) );
  NAND2_X1 u0_u15_u3_U58 (.A2( u0_u15_u3_n100 ) , .ZN( u0_u15_u3_n146 ) , .A1( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U59 (.A1( u0_u15_u3_n101 ) , .ZN( u0_u15_u3_n145 ) , .A2( u0_u15_u3_n99 ) );
  AOI221_X1 u0_u15_u3_U6 (.A( u0_u15_u3_n131 ) , .C2( u0_u15_u3_n132 ) , .C1( u0_u15_u3_n133 ) , .ZN( u0_u15_u3_n134 ) , .B1( u0_u15_u3_n143 ) , .B2( u0_u15_u3_n177 ) );
  NAND2_X1 u0_u15_u3_U60 (.A1( u0_u15_u3_n100 ) , .ZN( u0_u15_u3_n156 ) , .A2( u0_u15_u3_n99 ) );
  NAND2_X1 u0_u15_u3_U61 (.A2( u0_u15_u3_n101 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n148 ) );
  NAND2_X1 u0_u15_u3_U62 (.A1( u0_u15_u3_n100 ) , .A2( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n128 ) );
  NAND2_X1 u0_u15_u3_U63 (.A2( u0_u15_u3_n101 ) , .A1( u0_u15_u3_n102 ) , .ZN( u0_u15_u3_n152 ) );
  NAND2_X1 u0_u15_u3_U64 (.A2( u0_u15_u3_n101 ) , .ZN( u0_u15_u3_n114 ) , .A1( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U65 (.ZN( u0_u15_u3_n107 ) , .A1( u0_u15_u3_n97 ) , .A2( u0_u15_u3_n99 ) );
  NAND2_X1 u0_u15_u3_U66 (.A2( u0_u15_u3_n100 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n113 ) );
  NAND2_X1 u0_u15_u3_U67 (.A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n153 ) , .A2( u0_u15_u3_n97 ) );
  NAND2_X1 u0_u15_u3_U68 (.A2( u0_u15_u3_n103 ) , .A1( u0_u15_u3_n104 ) , .ZN( u0_u15_u3_n130 ) );
  NAND2_X1 u0_u15_u3_U69 (.A2( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n144 ) , .A1( u0_u15_u3_n96 ) );
  OAI22_X1 u0_u15_u3_U7 (.B2( u0_u15_u3_n147 ) , .A2( u0_u15_u3_n148 ) , .ZN( u0_u15_u3_n160 ) , .B1( u0_u15_u3_n165 ) , .A1( u0_u15_u3_n168 ) );
  NAND2_X1 u0_u15_u3_U70 (.A1( u0_u15_u3_n102 ) , .A2( u0_u15_u3_n103 ) , .ZN( u0_u15_u3_n108 ) );
  NOR2_X1 u0_u15_u3_U71 (.A2( u0_u15_X_19 ) , .A1( u0_u15_X_20 ) , .ZN( u0_u15_u3_n99 ) );
  NOR2_X1 u0_u15_u3_U72 (.A2( u0_u15_X_21 ) , .A1( u0_u15_X_24 ) , .ZN( u0_u15_u3_n103 ) );
  NOR2_X1 u0_u15_u3_U73 (.A2( u0_u15_X_24 ) , .A1( u0_u15_u3_n171 ) , .ZN( u0_u15_u3_n97 ) );
  NOR2_X1 u0_u15_u3_U74 (.A2( u0_u15_X_23 ) , .ZN( u0_u15_u3_n141 ) , .A1( u0_u15_u3_n166 ) );
  NOR2_X1 u0_u15_u3_U75 (.A2( u0_u15_X_19 ) , .A1( u0_u15_u3_n172 ) , .ZN( u0_u15_u3_n96 ) );
  NAND2_X1 u0_u15_u3_U76 (.A1( u0_u15_X_22 ) , .A2( u0_u15_X_23 ) , .ZN( u0_u15_u3_n154 ) );
  NAND2_X1 u0_u15_u3_U77 (.A1( u0_u15_X_23 ) , .ZN( u0_u15_u3_n149 ) , .A2( u0_u15_u3_n166 ) );
  NOR2_X1 u0_u15_u3_U78 (.A2( u0_u15_X_22 ) , .A1( u0_u15_X_23 ) , .ZN( u0_u15_u3_n121 ) );
  AND2_X1 u0_u15_u3_U79 (.A1( u0_u15_X_24 ) , .ZN( u0_u15_u3_n101 ) , .A2( u0_u15_u3_n171 ) );
  AND3_X1 u0_u15_u3_U8 (.A3( u0_u15_u3_n144 ) , .A2( u0_u15_u3_n145 ) , .A1( u0_u15_u3_n146 ) , .ZN( u0_u15_u3_n147 ) );
  AND2_X1 u0_u15_u3_U80 (.A1( u0_u15_X_19 ) , .ZN( u0_u15_u3_n102 ) , .A2( u0_u15_u3_n172 ) );
  AND2_X1 u0_u15_u3_U81 (.A1( u0_u15_X_21 ) , .A2( u0_u15_X_24 ) , .ZN( u0_u15_u3_n100 ) );
  AND2_X1 u0_u15_u3_U82 (.A2( u0_u15_X_19 ) , .A1( u0_u15_X_20 ) , .ZN( u0_u15_u3_n104 ) );
  INV_X1 u0_u15_u3_U83 (.A( u0_u15_X_22 ) , .ZN( u0_u15_u3_n166 ) );
  INV_X1 u0_u15_u3_U84 (.A( u0_u15_X_21 ) , .ZN( u0_u15_u3_n171 ) );
  INV_X1 u0_u15_u3_U85 (.A( u0_u15_X_20 ) , .ZN( u0_u15_u3_n172 ) );
  OR4_X1 u0_u15_u3_U86 (.ZN( u0_out15_10 ) , .A4( u0_u15_u3_n136 ) , .A3( u0_u15_u3_n137 ) , .A1( u0_u15_u3_n138 ) , .A2( u0_u15_u3_n139 ) );
  OAI222_X1 u0_u15_u3_U87 (.C1( u0_u15_u3_n128 ) , .ZN( u0_u15_u3_n137 ) , .B1( u0_u15_u3_n148 ) , .A2( u0_u15_u3_n150 ) , .B2( u0_u15_u3_n154 ) , .C2( u0_u15_u3_n164 ) , .A1( u0_u15_u3_n167 ) );
  OAI221_X1 u0_u15_u3_U88 (.A( u0_u15_u3_n134 ) , .B2( u0_u15_u3_n135 ) , .ZN( u0_u15_u3_n136 ) , .C1( u0_u15_u3_n149 ) , .B1( u0_u15_u3_n151 ) , .C2( u0_u15_u3_n183 ) );
  NAND4_X1 u0_u15_u3_U89 (.ZN( u0_out15_26 ) , .A4( u0_u15_u3_n109 ) , .A3( u0_u15_u3_n110 ) , .A2( u0_u15_u3_n111 ) , .A1( u0_u15_u3_n173 ) );
  INV_X1 u0_u15_u3_U9 (.A( u0_u15_u3_n143 ) , .ZN( u0_u15_u3_n168 ) );
  INV_X1 u0_u15_u3_U90 (.ZN( u0_u15_u3_n173 ) , .A( u0_u15_u3_n94 ) );
  OAI21_X1 u0_u15_u3_U91 (.ZN( u0_u15_u3_n111 ) , .B2( u0_u15_u3_n117 ) , .A( u0_u15_u3_n133 ) , .B1( u0_u15_u3_n176 ) );
  NAND4_X1 u0_u15_u3_U92 (.ZN( u0_out15_20 ) , .A4( u0_u15_u3_n122 ) , .A3( u0_u15_u3_n123 ) , .A1( u0_u15_u3_n175 ) , .A2( u0_u15_u3_n180 ) );
  INV_X1 u0_u15_u3_U93 (.A( u0_u15_u3_n126 ) , .ZN( u0_u15_u3_n180 ) );
  INV_X1 u0_u15_u3_U94 (.A( u0_u15_u3_n112 ) , .ZN( u0_u15_u3_n175 ) );
  NAND4_X1 u0_u15_u3_U95 (.ZN( u0_out15_1 ) , .A4( u0_u15_u3_n161 ) , .A3( u0_u15_u3_n162 ) , .A2( u0_u15_u3_n163 ) , .A1( u0_u15_u3_n185 ) );
  NAND2_X1 u0_u15_u3_U96 (.ZN( u0_u15_u3_n163 ) , .A2( u0_u15_u3_n170 ) , .A1( u0_u15_u3_n176 ) );
  AOI22_X1 u0_u15_u3_U97 (.B2( u0_u15_u3_n140 ) , .B1( u0_u15_u3_n141 ) , .A2( u0_u15_u3_n142 ) , .ZN( u0_u15_u3_n162 ) , .A1( u0_u15_u3_n177 ) );
  NAND3_X1 u0_u15_u3_U98 (.A1( u0_u15_u3_n114 ) , .ZN( u0_u15_u3_n115 ) , .A2( u0_u15_u3_n145 ) , .A3( u0_u15_u3_n153 ) );
  NAND3_X1 u0_u15_u3_U99 (.ZN( u0_u15_u3_n129 ) , .A2( u0_u15_u3_n144 ) , .A1( u0_u15_u3_n153 ) , .A3( u0_u15_u3_n182 ) );
  OAI22_X1 u0_u15_u4_U10 (.B2( u0_u15_u4_n135 ) , .ZN( u0_u15_u4_n137 ) , .B1( u0_u15_u4_n153 ) , .A1( u0_u15_u4_n155 ) , .A2( u0_u15_u4_n171 ) );
  AND3_X1 u0_u15_u4_U11 (.A2( u0_u15_u4_n134 ) , .ZN( u0_u15_u4_n135 ) , .A3( u0_u15_u4_n145 ) , .A1( u0_u15_u4_n157 ) );
  OR3_X1 u0_u15_u4_U12 (.A3( u0_u15_u4_n114 ) , .A2( u0_u15_u4_n115 ) , .A1( u0_u15_u4_n116 ) , .ZN( u0_u15_u4_n136 ) );
  AOI21_X1 u0_u15_u4_U13 (.A( u0_u15_u4_n113 ) , .ZN( u0_u15_u4_n116 ) , .B2( u0_u15_u4_n173 ) , .B1( u0_u15_u4_n174 ) );
  AOI21_X1 u0_u15_u4_U14 (.ZN( u0_u15_u4_n115 ) , .B2( u0_u15_u4_n145 ) , .B1( u0_u15_u4_n146 ) , .A( u0_u15_u4_n156 ) );
  OAI22_X1 u0_u15_u4_U15 (.ZN( u0_u15_u4_n114 ) , .A2( u0_u15_u4_n121 ) , .B1( u0_u15_u4_n160 ) , .B2( u0_u15_u4_n170 ) , .A1( u0_u15_u4_n171 ) );
  NAND2_X1 u0_u15_u4_U16 (.ZN( u0_u15_u4_n132 ) , .A2( u0_u15_u4_n170 ) , .A1( u0_u15_u4_n173 ) );
  AOI21_X1 u0_u15_u4_U17 (.B2( u0_u15_u4_n160 ) , .B1( u0_u15_u4_n161 ) , .ZN( u0_u15_u4_n162 ) , .A( u0_u15_u4_n170 ) );
  AOI21_X1 u0_u15_u4_U18 (.ZN( u0_u15_u4_n107 ) , .B2( u0_u15_u4_n143 ) , .A( u0_u15_u4_n174 ) , .B1( u0_u15_u4_n184 ) );
  AOI21_X1 u0_u15_u4_U19 (.B2( u0_u15_u4_n158 ) , .B1( u0_u15_u4_n159 ) , .ZN( u0_u15_u4_n163 ) , .A( u0_u15_u4_n174 ) );
  AOI21_X1 u0_u15_u4_U20 (.A( u0_u15_u4_n153 ) , .B2( u0_u15_u4_n154 ) , .B1( u0_u15_u4_n155 ) , .ZN( u0_u15_u4_n165 ) );
  AOI21_X1 u0_u15_u4_U21 (.A( u0_u15_u4_n156 ) , .B2( u0_u15_u4_n157 ) , .ZN( u0_u15_u4_n164 ) , .B1( u0_u15_u4_n184 ) );
  INV_X1 u0_u15_u4_U22 (.A( u0_u15_u4_n138 ) , .ZN( u0_u15_u4_n170 ) );
  AND2_X1 u0_u15_u4_U23 (.A2( u0_u15_u4_n120 ) , .ZN( u0_u15_u4_n155 ) , .A1( u0_u15_u4_n160 ) );
  INV_X1 u0_u15_u4_U24 (.A( u0_u15_u4_n156 ) , .ZN( u0_u15_u4_n175 ) );
  NAND2_X1 u0_u15_u4_U25 (.A2( u0_u15_u4_n118 ) , .ZN( u0_u15_u4_n131 ) , .A1( u0_u15_u4_n147 ) );
  NAND2_X1 u0_u15_u4_U26 (.A1( u0_u15_u4_n119 ) , .A2( u0_u15_u4_n120 ) , .ZN( u0_u15_u4_n130 ) );
  NAND2_X1 u0_u15_u4_U27 (.ZN( u0_u15_u4_n117 ) , .A2( u0_u15_u4_n118 ) , .A1( u0_u15_u4_n148 ) );
  NAND2_X1 u0_u15_u4_U28 (.ZN( u0_u15_u4_n129 ) , .A1( u0_u15_u4_n134 ) , .A2( u0_u15_u4_n148 ) );
  AND3_X1 u0_u15_u4_U29 (.A1( u0_u15_u4_n119 ) , .A2( u0_u15_u4_n143 ) , .A3( u0_u15_u4_n154 ) , .ZN( u0_u15_u4_n161 ) );
  NOR2_X1 u0_u15_u4_U3 (.ZN( u0_u15_u4_n121 ) , .A1( u0_u15_u4_n181 ) , .A2( u0_u15_u4_n182 ) );
  AND2_X1 u0_u15_u4_U30 (.A1( u0_u15_u4_n145 ) , .A2( u0_u15_u4_n147 ) , .ZN( u0_u15_u4_n159 ) );
  INV_X1 u0_u15_u4_U31 (.A( u0_u15_u4_n158 ) , .ZN( u0_u15_u4_n182 ) );
  INV_X1 u0_u15_u4_U32 (.ZN( u0_u15_u4_n181 ) , .A( u0_u15_u4_n96 ) );
  INV_X1 u0_u15_u4_U33 (.A( u0_u15_u4_n144 ) , .ZN( u0_u15_u4_n179 ) );
  INV_X1 u0_u15_u4_U34 (.A( u0_u15_u4_n157 ) , .ZN( u0_u15_u4_n178 ) );
  NAND2_X1 u0_u15_u4_U35 (.A2( u0_u15_u4_n154 ) , .A1( u0_u15_u4_n96 ) , .ZN( u0_u15_u4_n97 ) );
  INV_X1 u0_u15_u4_U36 (.ZN( u0_u15_u4_n186 ) , .A( u0_u15_u4_n95 ) );
  OAI221_X1 u0_u15_u4_U37 (.C1( u0_u15_u4_n134 ) , .B1( u0_u15_u4_n158 ) , .B2( u0_u15_u4_n171 ) , .C2( u0_u15_u4_n173 ) , .A( u0_u15_u4_n94 ) , .ZN( u0_u15_u4_n95 ) );
  AOI222_X1 u0_u15_u4_U38 (.B2( u0_u15_u4_n132 ) , .A1( u0_u15_u4_n138 ) , .C2( u0_u15_u4_n175 ) , .A2( u0_u15_u4_n179 ) , .C1( u0_u15_u4_n181 ) , .B1( u0_u15_u4_n185 ) , .ZN( u0_u15_u4_n94 ) );
  INV_X1 u0_u15_u4_U39 (.A( u0_u15_u4_n113 ) , .ZN( u0_u15_u4_n185 ) );
  INV_X1 u0_u15_u4_U4 (.A( u0_u15_u4_n117 ) , .ZN( u0_u15_u4_n184 ) );
  INV_X1 u0_u15_u4_U40 (.A( u0_u15_u4_n143 ) , .ZN( u0_u15_u4_n183 ) );
  NOR2_X1 u0_u15_u4_U41 (.ZN( u0_u15_u4_n138 ) , .A1( u0_u15_u4_n168 ) , .A2( u0_u15_u4_n169 ) );
  NOR2_X1 u0_u15_u4_U42 (.A1( u0_u15_u4_n150 ) , .A2( u0_u15_u4_n152 ) , .ZN( u0_u15_u4_n153 ) );
  NOR2_X1 u0_u15_u4_U43 (.A2( u0_u15_u4_n128 ) , .A1( u0_u15_u4_n138 ) , .ZN( u0_u15_u4_n156 ) );
  AOI22_X1 u0_u15_u4_U44 (.B2( u0_u15_u4_n122 ) , .A1( u0_u15_u4_n123 ) , .ZN( u0_u15_u4_n124 ) , .B1( u0_u15_u4_n128 ) , .A2( u0_u15_u4_n172 ) );
  NAND2_X1 u0_u15_u4_U45 (.A2( u0_u15_u4_n120 ) , .ZN( u0_u15_u4_n123 ) , .A1( u0_u15_u4_n161 ) );
  INV_X1 u0_u15_u4_U46 (.A( u0_u15_u4_n153 ) , .ZN( u0_u15_u4_n172 ) );
  AOI22_X1 u0_u15_u4_U47 (.B2( u0_u15_u4_n132 ) , .A2( u0_u15_u4_n133 ) , .ZN( u0_u15_u4_n140 ) , .A1( u0_u15_u4_n150 ) , .B1( u0_u15_u4_n179 ) );
  NAND2_X1 u0_u15_u4_U48 (.ZN( u0_u15_u4_n133 ) , .A2( u0_u15_u4_n146 ) , .A1( u0_u15_u4_n154 ) );
  NAND2_X1 u0_u15_u4_U49 (.A1( u0_u15_u4_n103 ) , .ZN( u0_u15_u4_n154 ) , .A2( u0_u15_u4_n98 ) );
  NOR4_X1 u0_u15_u4_U5 (.A4( u0_u15_u4_n106 ) , .A3( u0_u15_u4_n107 ) , .A2( u0_u15_u4_n108 ) , .A1( u0_u15_u4_n109 ) , .ZN( u0_u15_u4_n110 ) );
  NAND2_X1 u0_u15_u4_U50 (.A1( u0_u15_u4_n101 ) , .ZN( u0_u15_u4_n158 ) , .A2( u0_u15_u4_n99 ) );
  AOI21_X1 u0_u15_u4_U51 (.ZN( u0_u15_u4_n127 ) , .A( u0_u15_u4_n136 ) , .B2( u0_u15_u4_n150 ) , .B1( u0_u15_u4_n180 ) );
  INV_X1 u0_u15_u4_U52 (.A( u0_u15_u4_n160 ) , .ZN( u0_u15_u4_n180 ) );
  NAND2_X1 u0_u15_u4_U53 (.A2( u0_u15_u4_n104 ) , .A1( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n146 ) );
  NAND2_X1 u0_u15_u4_U54 (.A2( u0_u15_u4_n101 ) , .A1( u0_u15_u4_n102 ) , .ZN( u0_u15_u4_n160 ) );
  NAND2_X1 u0_u15_u4_U55 (.ZN( u0_u15_u4_n134 ) , .A1( u0_u15_u4_n98 ) , .A2( u0_u15_u4_n99 ) );
  NAND2_X1 u0_u15_u4_U56 (.A1( u0_u15_u4_n103 ) , .A2( u0_u15_u4_n104 ) , .ZN( u0_u15_u4_n143 ) );
  NAND2_X1 u0_u15_u4_U57 (.A2( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n145 ) , .A1( u0_u15_u4_n98 ) );
  NAND2_X1 u0_u15_u4_U58 (.A1( u0_u15_u4_n100 ) , .A2( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n120 ) );
  NAND2_X1 u0_u15_u4_U59 (.A1( u0_u15_u4_n102 ) , .A2( u0_u15_u4_n104 ) , .ZN( u0_u15_u4_n148 ) );
  AOI21_X1 u0_u15_u4_U6 (.ZN( u0_u15_u4_n106 ) , .B2( u0_u15_u4_n146 ) , .B1( u0_u15_u4_n158 ) , .A( u0_u15_u4_n170 ) );
  NAND2_X1 u0_u15_u4_U60 (.A2( u0_u15_u4_n100 ) , .A1( u0_u15_u4_n103 ) , .ZN( u0_u15_u4_n157 ) );
  INV_X1 u0_u15_u4_U61 (.A( u0_u15_u4_n150 ) , .ZN( u0_u15_u4_n173 ) );
  INV_X1 u0_u15_u4_U62 (.A( u0_u15_u4_n152 ) , .ZN( u0_u15_u4_n171 ) );
  NAND2_X1 u0_u15_u4_U63 (.A1( u0_u15_u4_n100 ) , .ZN( u0_u15_u4_n118 ) , .A2( u0_u15_u4_n99 ) );
  NAND2_X1 u0_u15_u4_U64 (.A2( u0_u15_u4_n100 ) , .A1( u0_u15_u4_n102 ) , .ZN( u0_u15_u4_n144 ) );
  NAND2_X1 u0_u15_u4_U65 (.A2( u0_u15_u4_n101 ) , .A1( u0_u15_u4_n105 ) , .ZN( u0_u15_u4_n96 ) );
  INV_X1 u0_u15_u4_U66 (.A( u0_u15_u4_n128 ) , .ZN( u0_u15_u4_n174 ) );
  NAND2_X1 u0_u15_u4_U67 (.A2( u0_u15_u4_n102 ) , .ZN( u0_u15_u4_n119 ) , .A1( u0_u15_u4_n98 ) );
  NAND2_X1 u0_u15_u4_U68 (.A2( u0_u15_u4_n101 ) , .A1( u0_u15_u4_n103 ) , .ZN( u0_u15_u4_n147 ) );
  NAND2_X1 u0_u15_u4_U69 (.A2( u0_u15_u4_n104 ) , .ZN( u0_u15_u4_n113 ) , .A1( u0_u15_u4_n99 ) );
  AOI21_X1 u0_u15_u4_U7 (.ZN( u0_u15_u4_n108 ) , .B2( u0_u15_u4_n134 ) , .B1( u0_u15_u4_n155 ) , .A( u0_u15_u4_n156 ) );
  NOR2_X1 u0_u15_u4_U70 (.A2( u0_u15_X_28 ) , .ZN( u0_u15_u4_n150 ) , .A1( u0_u15_u4_n168 ) );
  NOR2_X1 u0_u15_u4_U71 (.A2( u0_u15_X_29 ) , .ZN( u0_u15_u4_n152 ) , .A1( u0_u15_u4_n169 ) );
  NOR2_X1 u0_u15_u4_U72 (.A2( u0_u15_X_26 ) , .ZN( u0_u15_u4_n100 ) , .A1( u0_u15_u4_n177 ) );
  NOR2_X1 u0_u15_u4_U73 (.A2( u0_u15_X_30 ) , .ZN( u0_u15_u4_n105 ) , .A1( u0_u15_u4_n176 ) );
  NOR2_X1 u0_u15_u4_U74 (.A2( u0_u15_X_28 ) , .A1( u0_u15_X_29 ) , .ZN( u0_u15_u4_n128 ) );
  NOR2_X1 u0_u15_u4_U75 (.A2( u0_u15_X_25 ) , .A1( u0_u15_X_26 ) , .ZN( u0_u15_u4_n98 ) );
  NOR2_X1 u0_u15_u4_U76 (.A2( u0_u15_X_27 ) , .A1( u0_u15_X_30 ) , .ZN( u0_u15_u4_n102 ) );
  AND2_X1 u0_u15_u4_U77 (.A2( u0_u15_X_25 ) , .A1( u0_u15_X_26 ) , .ZN( u0_u15_u4_n104 ) );
  AND2_X1 u0_u15_u4_U78 (.A1( u0_u15_X_30 ) , .A2( u0_u15_u4_n176 ) , .ZN( u0_u15_u4_n99 ) );
  AND2_X1 u0_u15_u4_U79 (.A1( u0_u15_X_26 ) , .ZN( u0_u15_u4_n101 ) , .A2( u0_u15_u4_n177 ) );
  AOI21_X1 u0_u15_u4_U8 (.ZN( u0_u15_u4_n109 ) , .A( u0_u15_u4_n153 ) , .B1( u0_u15_u4_n159 ) , .B2( u0_u15_u4_n184 ) );
  AND2_X1 u0_u15_u4_U80 (.A1( u0_u15_X_27 ) , .A2( u0_u15_X_30 ) , .ZN( u0_u15_u4_n103 ) );
  INV_X1 u0_u15_u4_U81 (.A( u0_u15_X_28 ) , .ZN( u0_u15_u4_n169 ) );
  INV_X1 u0_u15_u4_U82 (.A( u0_u15_X_29 ) , .ZN( u0_u15_u4_n168 ) );
  INV_X1 u0_u15_u4_U83 (.A( u0_u15_X_25 ) , .ZN( u0_u15_u4_n177 ) );
  INV_X1 u0_u15_u4_U84 (.A( u0_u15_X_27 ) , .ZN( u0_u15_u4_n176 ) );
  NAND4_X1 u0_u15_u4_U85 (.ZN( u0_out15_25 ) , .A4( u0_u15_u4_n139 ) , .A3( u0_u15_u4_n140 ) , .A2( u0_u15_u4_n141 ) , .A1( u0_u15_u4_n142 ) );
  OAI21_X1 u0_u15_u4_U86 (.A( u0_u15_u4_n128 ) , .B2( u0_u15_u4_n129 ) , .B1( u0_u15_u4_n130 ) , .ZN( u0_u15_u4_n142 ) );
  OAI21_X1 u0_u15_u4_U87 (.B2( u0_u15_u4_n131 ) , .ZN( u0_u15_u4_n141 ) , .A( u0_u15_u4_n175 ) , .B1( u0_u15_u4_n183 ) );
  NAND4_X1 u0_u15_u4_U88 (.ZN( u0_out15_14 ) , .A4( u0_u15_u4_n124 ) , .A3( u0_u15_u4_n125 ) , .A2( u0_u15_u4_n126 ) , .A1( u0_u15_u4_n127 ) );
  AOI22_X1 u0_u15_u4_U89 (.B2( u0_u15_u4_n117 ) , .ZN( u0_u15_u4_n126 ) , .A1( u0_u15_u4_n129 ) , .B1( u0_u15_u4_n152 ) , .A2( u0_u15_u4_n175 ) );
  AOI211_X1 u0_u15_u4_U9 (.B( u0_u15_u4_n136 ) , .A( u0_u15_u4_n137 ) , .C2( u0_u15_u4_n138 ) , .ZN( u0_u15_u4_n139 ) , .C1( u0_u15_u4_n182 ) );
  AOI22_X1 u0_u15_u4_U90 (.ZN( u0_u15_u4_n125 ) , .B2( u0_u15_u4_n131 ) , .A2( u0_u15_u4_n132 ) , .B1( u0_u15_u4_n138 ) , .A1( u0_u15_u4_n178 ) );
  AOI22_X1 u0_u15_u4_U91 (.B2( u0_u15_u4_n149 ) , .B1( u0_u15_u4_n150 ) , .A2( u0_u15_u4_n151 ) , .A1( u0_u15_u4_n152 ) , .ZN( u0_u15_u4_n167 ) );
  NOR4_X1 u0_u15_u4_U92 (.A4( u0_u15_u4_n162 ) , .A3( u0_u15_u4_n163 ) , .A2( u0_u15_u4_n164 ) , .A1( u0_u15_u4_n165 ) , .ZN( u0_u15_u4_n166 ) );
  NAND4_X1 u0_u15_u4_U93 (.ZN( u0_out15_8 ) , .A4( u0_u15_u4_n110 ) , .A3( u0_u15_u4_n111 ) , .A2( u0_u15_u4_n112 ) , .A1( u0_u15_u4_n186 ) );
  NAND2_X1 u0_u15_u4_U94 (.ZN( u0_u15_u4_n112 ) , .A2( u0_u15_u4_n130 ) , .A1( u0_u15_u4_n150 ) );
  AOI22_X1 u0_u15_u4_U95 (.ZN( u0_u15_u4_n111 ) , .B2( u0_u15_u4_n132 ) , .A1( u0_u15_u4_n152 ) , .B1( u0_u15_u4_n178 ) , .A2( u0_u15_u4_n97 ) );
  NAND3_X1 u0_u15_u4_U96 (.ZN( u0_out15_3 ) , .A3( u0_u15_u4_n166 ) , .A1( u0_u15_u4_n167 ) , .A2( u0_u15_u4_n186 ) );
  NAND3_X1 u0_u15_u4_U97 (.A3( u0_u15_u4_n146 ) , .A2( u0_u15_u4_n147 ) , .A1( u0_u15_u4_n148 ) , .ZN( u0_u15_u4_n149 ) );
  NAND3_X1 u0_u15_u4_U98 (.A3( u0_u15_u4_n143 ) , .A2( u0_u15_u4_n144 ) , .A1( u0_u15_u4_n145 ) , .ZN( u0_u15_u4_n151 ) );
  NAND3_X1 u0_u15_u4_U99 (.A3( u0_u15_u4_n121 ) , .ZN( u0_u15_u4_n122 ) , .A2( u0_u15_u4_n144 ) , .A1( u0_u15_u4_n154 ) );
  XOR2_X1 u0_u1_U1 (.B( u0_K2_9 ) , .A( u0_R0_6 ) , .Z( u0_u1_X_9 ) );
  XOR2_X1 u0_u1_U13 (.B( u0_K2_42 ) , .A( u0_R0_29 ) , .Z( u0_u1_X_42 ) );
  XOR2_X1 u0_u1_U14 (.B( u0_K2_41 ) , .A( u0_R0_28 ) , .Z( u0_u1_X_41 ) );
  XOR2_X1 u0_u1_U15 (.B( u0_K2_40 ) , .A( u0_R0_27 ) , .Z( u0_u1_X_40 ) );
  XOR2_X1 u0_u1_U16 (.B( u0_K2_3 ) , .A( u0_R0_2 ) , .Z( u0_u1_X_3 ) );
  XOR2_X1 u0_u1_U17 (.B( u0_K2_39 ) , .A( u0_R0_26 ) , .Z( u0_u1_X_39 ) );
  XOR2_X1 u0_u1_U18 (.B( u0_K2_38 ) , .A( u0_R0_25 ) , .Z( u0_u1_X_38 ) );
  XOR2_X1 u0_u1_U19 (.B( u0_K2_37 ) , .A( u0_R0_24 ) , .Z( u0_u1_X_37 ) );
  XOR2_X1 u0_u1_U2 (.B( u0_K2_8 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_8 ) );
  XOR2_X1 u0_u1_U27 (.B( u0_K2_2 ) , .A( u0_R0_1 ) , .Z( u0_u1_X_2 ) );
  XOR2_X1 u0_u1_U3 (.B( u0_K2_7 ) , .A( u0_R0_4 ) , .Z( u0_u1_X_7 ) );
  XOR2_X1 u0_u1_U38 (.B( u0_K2_1 ) , .A( u0_R0_32 ) , .Z( u0_u1_X_1 ) );
  XOR2_X1 u0_u1_U4 (.B( u0_K2_6 ) , .A( u0_R0_5 ) , .Z( u0_u1_X_6 ) );
  XOR2_X1 u0_u1_U40 (.B( u0_K2_18 ) , .A( u0_R0_13 ) , .Z( u0_u1_X_18 ) );
  XOR2_X1 u0_u1_U41 (.B( u0_K2_17 ) , .A( u0_R0_12 ) , .Z( u0_u1_X_17 ) );
  XOR2_X1 u0_u1_U42 (.B( u0_K2_16 ) , .A( u0_R0_11 ) , .Z( u0_u1_X_16 ) );
  XOR2_X1 u0_u1_U43 (.B( u0_K2_15 ) , .A( u0_R0_10 ) , .Z( u0_u1_X_15 ) );
  XOR2_X1 u0_u1_U44 (.B( u0_K2_14 ) , .A( u0_R0_9 ) , .Z( u0_u1_X_14 ) );
  XOR2_X1 u0_u1_U45 (.B( u0_K2_13 ) , .A( u0_R0_8 ) , .Z( u0_u1_X_13 ) );
  XOR2_X1 u0_u1_U46 (.B( u0_K2_12 ) , .A( u0_R0_9 ) , .Z( u0_u1_X_12 ) );
  XOR2_X1 u0_u1_U47 (.B( u0_K2_11 ) , .A( u0_R0_8 ) , .Z( u0_u1_X_11 ) );
  XOR2_X1 u0_u1_U48 (.B( u0_K2_10 ) , .A( u0_R0_7 ) , .Z( u0_u1_X_10 ) );
  XOR2_X1 u0_u1_U5 (.B( u0_K2_5 ) , .A( u0_R0_4 ) , .Z( u0_u1_X_5 ) );
  XOR2_X1 u0_u1_U6 (.B( u0_K2_4 ) , .A( u0_R0_3 ) , .Z( u0_u1_X_4 ) );
  AND3_X1 u0_u1_u0_U10 (.A2( u0_u1_u0_n112 ) , .ZN( u0_u1_u0_n127 ) , .A3( u0_u1_u0_n130 ) , .A1( u0_u1_u0_n148 ) );
  NAND2_X1 u0_u1_u0_U11 (.ZN( u0_u1_u0_n113 ) , .A1( u0_u1_u0_n139 ) , .A2( u0_u1_u0_n149 ) );
  AND2_X1 u0_u1_u0_U12 (.ZN( u0_u1_u0_n107 ) , .A1( u0_u1_u0_n130 ) , .A2( u0_u1_u0_n140 ) );
  AND2_X1 u0_u1_u0_U13 (.A2( u0_u1_u0_n129 ) , .A1( u0_u1_u0_n130 ) , .ZN( u0_u1_u0_n151 ) );
  AND2_X1 u0_u1_u0_U14 (.A1( u0_u1_u0_n108 ) , .A2( u0_u1_u0_n125 ) , .ZN( u0_u1_u0_n145 ) );
  INV_X1 u0_u1_u0_U15 (.A( u0_u1_u0_n143 ) , .ZN( u0_u1_u0_n173 ) );
  NOR2_X1 u0_u1_u0_U16 (.A2( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n147 ) , .A1( u0_u1_u0_n160 ) );
  NOR2_X1 u0_u1_u0_U17 (.A1( u0_u1_u0_n163 ) , .A2( u0_u1_u0_n164 ) , .ZN( u0_u1_u0_n95 ) );
  AOI21_X1 u0_u1_u0_U18 (.B1( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n132 ) , .A( u0_u1_u0_n165 ) , .B2( u0_u1_u0_n93 ) );
  INV_X1 u0_u1_u0_U19 (.A( u0_u1_u0_n142 ) , .ZN( u0_u1_u0_n165 ) );
  OAI221_X1 u0_u1_u0_U20 (.C1( u0_u1_u0_n121 ) , .ZN( u0_u1_u0_n122 ) , .B2( u0_u1_u0_n127 ) , .A( u0_u1_u0_n143 ) , .B1( u0_u1_u0_n144 ) , .C2( u0_u1_u0_n147 ) );
  OAI22_X1 u0_u1_u0_U21 (.B1( u0_u1_u0_n125 ) , .ZN( u0_u1_u0_n126 ) , .A1( u0_u1_u0_n138 ) , .A2( u0_u1_u0_n146 ) , .B2( u0_u1_u0_n147 ) );
  OAI22_X1 u0_u1_u0_U22 (.B1( u0_u1_u0_n131 ) , .A1( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n147 ) , .A2( u0_u1_u0_n90 ) , .ZN( u0_u1_u0_n91 ) );
  AND3_X1 u0_u1_u0_U23 (.A3( u0_u1_u0_n121 ) , .A2( u0_u1_u0_n125 ) , .A1( u0_u1_u0_n148 ) , .ZN( u0_u1_u0_n90 ) );
  INV_X1 u0_u1_u0_U24 (.A( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n161 ) );
  NOR2_X1 u0_u1_u0_U25 (.A1( u0_u1_u0_n120 ) , .ZN( u0_u1_u0_n143 ) , .A2( u0_u1_u0_n167 ) );
  OAI221_X1 u0_u1_u0_U26 (.C1( u0_u1_u0_n112 ) , .ZN( u0_u1_u0_n120 ) , .B1( u0_u1_u0_n138 ) , .B2( u0_u1_u0_n141 ) , .C2( u0_u1_u0_n147 ) , .A( u0_u1_u0_n172 ) );
  AOI211_X1 u0_u1_u0_U27 (.B( u0_u1_u0_n115 ) , .A( u0_u1_u0_n116 ) , .C2( u0_u1_u0_n117 ) , .C1( u0_u1_u0_n118 ) , .ZN( u0_u1_u0_n119 ) );
  AOI22_X1 u0_u1_u0_U28 (.B2( u0_u1_u0_n109 ) , .A2( u0_u1_u0_n110 ) , .ZN( u0_u1_u0_n111 ) , .B1( u0_u1_u0_n118 ) , .A1( u0_u1_u0_n160 ) );
  INV_X1 u0_u1_u0_U29 (.A( u0_u1_u0_n118 ) , .ZN( u0_u1_u0_n158 ) );
  INV_X1 u0_u1_u0_U3 (.A( u0_u1_u0_n113 ) , .ZN( u0_u1_u0_n166 ) );
  AOI21_X1 u0_u1_u0_U30 (.ZN( u0_u1_u0_n104 ) , .B1( u0_u1_u0_n107 ) , .B2( u0_u1_u0_n141 ) , .A( u0_u1_u0_n144 ) );
  AOI21_X1 u0_u1_u0_U31 (.B1( u0_u1_u0_n127 ) , .B2( u0_u1_u0_n129 ) , .A( u0_u1_u0_n138 ) , .ZN( u0_u1_u0_n96 ) );
  AOI21_X1 u0_u1_u0_U32 (.ZN( u0_u1_u0_n116 ) , .B2( u0_u1_u0_n142 ) , .A( u0_u1_u0_n144 ) , .B1( u0_u1_u0_n166 ) );
  NAND2_X1 u0_u1_u0_U33 (.A1( u0_u1_u0_n100 ) , .A2( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n125 ) );
  NAND2_X1 u0_u1_u0_U34 (.A2( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n140 ) , .A1( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U35 (.A1( u0_u1_u0_n101 ) , .A2( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n150 ) );
  INV_X1 u0_u1_u0_U36 (.A( u0_u1_u0_n138 ) , .ZN( u0_u1_u0_n160 ) );
  NAND2_X1 u0_u1_u0_U37 (.ZN( u0_u1_u0_n142 ) , .A1( u0_u1_u0_n94 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U38 (.A1( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n128 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U39 (.A2( u0_u1_u0_n102 ) , .A1( u0_u1_u0_n103 ) , .ZN( u0_u1_u0_n149 ) );
  AOI21_X1 u0_u1_u0_U4 (.B1( u0_u1_u0_n114 ) , .ZN( u0_u1_u0_n115 ) , .B2( u0_u1_u0_n129 ) , .A( u0_u1_u0_n161 ) );
  NAND2_X1 u0_u1_u0_U40 (.A1( u0_u1_u0_n100 ) , .ZN( u0_u1_u0_n129 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U41 (.A2( u0_u1_u0_n100 ) , .A1( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n139 ) );
  NAND2_X1 u0_u1_u0_U42 (.A2( u0_u1_u0_n100 ) , .ZN( u0_u1_u0_n131 ) , .A1( u0_u1_u0_n92 ) );
  NAND2_X1 u0_u1_u0_U43 (.ZN( u0_u1_u0_n108 ) , .A1( u0_u1_u0_n92 ) , .A2( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U44 (.ZN( u0_u1_u0_n148 ) , .A1( u0_u1_u0_n93 ) , .A2( u0_u1_u0_n95 ) );
  NAND2_X1 u0_u1_u0_U45 (.A2( u0_u1_u0_n102 ) , .ZN( u0_u1_u0_n114 ) , .A1( u0_u1_u0_n92 ) );
  NAND2_X1 u0_u1_u0_U46 (.A1( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n130 ) , .A2( u0_u1_u0_n94 ) );
  NAND2_X1 u0_u1_u0_U47 (.A2( u0_u1_u0_n101 ) , .ZN( u0_u1_u0_n121 ) , .A1( u0_u1_u0_n93 ) );
  INV_X1 u0_u1_u0_U48 (.ZN( u0_u1_u0_n172 ) , .A( u0_u1_u0_n88 ) );
  OAI222_X1 u0_u1_u0_U49 (.C1( u0_u1_u0_n108 ) , .A1( u0_u1_u0_n125 ) , .B2( u0_u1_u0_n128 ) , .B1( u0_u1_u0_n144 ) , .A2( u0_u1_u0_n158 ) , .C2( u0_u1_u0_n161 ) , .ZN( u0_u1_u0_n88 ) );
  AOI21_X1 u0_u1_u0_U5 (.B2( u0_u1_u0_n131 ) , .ZN( u0_u1_u0_n134 ) , .B1( u0_u1_u0_n151 ) , .A( u0_u1_u0_n158 ) );
  NAND2_X1 u0_u1_u0_U50 (.ZN( u0_u1_u0_n112 ) , .A2( u0_u1_u0_n92 ) , .A1( u0_u1_u0_n93 ) );
  OR3_X1 u0_u1_u0_U51 (.A3( u0_u1_u0_n152 ) , .A2( u0_u1_u0_n153 ) , .A1( u0_u1_u0_n154 ) , .ZN( u0_u1_u0_n155 ) );
  AOI21_X1 u0_u1_u0_U52 (.B2( u0_u1_u0_n150 ) , .B1( u0_u1_u0_n151 ) , .ZN( u0_u1_u0_n152 ) , .A( u0_u1_u0_n158 ) );
  AOI21_X1 u0_u1_u0_U53 (.A( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n145 ) , .B1( u0_u1_u0_n146 ) , .ZN( u0_u1_u0_n154 ) );
  AOI21_X1 u0_u1_u0_U54 (.A( u0_u1_u0_n147 ) , .B2( u0_u1_u0_n148 ) , .B1( u0_u1_u0_n149 ) , .ZN( u0_u1_u0_n153 ) );
  INV_X1 u0_u1_u0_U55 (.ZN( u0_u1_u0_n171 ) , .A( u0_u1_u0_n99 ) );
  OAI211_X1 u0_u1_u0_U56 (.C2( u0_u1_u0_n140 ) , .C1( u0_u1_u0_n161 ) , .A( u0_u1_u0_n169 ) , .B( u0_u1_u0_n98 ) , .ZN( u0_u1_u0_n99 ) );
  INV_X1 u0_u1_u0_U57 (.ZN( u0_u1_u0_n169 ) , .A( u0_u1_u0_n91 ) );
  AOI211_X1 u0_u1_u0_U58 (.C1( u0_u1_u0_n118 ) , .A( u0_u1_u0_n123 ) , .B( u0_u1_u0_n96 ) , .C2( u0_u1_u0_n97 ) , .ZN( u0_u1_u0_n98 ) );
  NOR2_X1 u0_u1_u0_U59 (.A2( u0_u1_X_2 ) , .ZN( u0_u1_u0_n103 ) , .A1( u0_u1_u0_n164 ) );
  NOR2_X1 u0_u1_u0_U6 (.A1( u0_u1_u0_n108 ) , .ZN( u0_u1_u0_n123 ) , .A2( u0_u1_u0_n158 ) );
  NOR2_X1 u0_u1_u0_U60 (.A2( u0_u1_X_3 ) , .A1( u0_u1_X_6 ) , .ZN( u0_u1_u0_n94 ) );
  NOR2_X1 u0_u1_u0_U61 (.A2( u0_u1_X_6 ) , .ZN( u0_u1_u0_n100 ) , .A1( u0_u1_u0_n162 ) );
  NOR2_X1 u0_u1_u0_U62 (.A2( u0_u1_X_4 ) , .A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n118 ) );
  NOR2_X1 u0_u1_u0_U63 (.A2( u0_u1_X_1 ) , .A1( u0_u1_X_2 ) , .ZN( u0_u1_u0_n92 ) );
  NOR2_X1 u0_u1_u0_U64 (.A2( u0_u1_X_1 ) , .ZN( u0_u1_u0_n101 ) , .A1( u0_u1_u0_n163 ) );
  NAND2_X1 u0_u1_u0_U65 (.A2( u0_u1_X_4 ) , .A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n144 ) );
  NOR2_X1 u0_u1_u0_U66 (.A2( u0_u1_X_5 ) , .ZN( u0_u1_u0_n136 ) , .A1( u0_u1_u0_n159 ) );
  NAND2_X1 u0_u1_u0_U67 (.A1( u0_u1_X_5 ) , .ZN( u0_u1_u0_n138 ) , .A2( u0_u1_u0_n159 ) );
  AND2_X1 u0_u1_u0_U68 (.A2( u0_u1_X_3 ) , .A1( u0_u1_X_6 ) , .ZN( u0_u1_u0_n102 ) );
  AND2_X1 u0_u1_u0_U69 (.A1( u0_u1_X_6 ) , .A2( u0_u1_u0_n162 ) , .ZN( u0_u1_u0_n93 ) );
  OAI21_X1 u0_u1_u0_U7 (.B1( u0_u1_u0_n150 ) , .B2( u0_u1_u0_n158 ) , .A( u0_u1_u0_n172 ) , .ZN( u0_u1_u0_n89 ) );
  INV_X1 u0_u1_u0_U70 (.A( u0_u1_X_4 ) , .ZN( u0_u1_u0_n159 ) );
  INV_X1 u0_u1_u0_U71 (.A( u0_u1_X_1 ) , .ZN( u0_u1_u0_n164 ) );
  INV_X1 u0_u1_u0_U72 (.A( u0_u1_X_2 ) , .ZN( u0_u1_u0_n163 ) );
  INV_X1 u0_u1_u0_U73 (.A( u0_u1_X_3 ) , .ZN( u0_u1_u0_n162 ) );
  INV_X1 u0_u1_u0_U74 (.ZN( u0_u1_u0_n174 ) , .A( u0_u1_u0_n89 ) );
  AOI211_X1 u0_u1_u0_U75 (.B( u0_u1_u0_n104 ) , .A( u0_u1_u0_n105 ) , .ZN( u0_u1_u0_n106 ) , .C2( u0_u1_u0_n113 ) , .C1( u0_u1_u0_n160 ) );
  INV_X1 u0_u1_u0_U76 (.A( u0_u1_u0_n126 ) , .ZN( u0_u1_u0_n168 ) );
  AOI211_X1 u0_u1_u0_U77 (.B( u0_u1_u0_n133 ) , .A( u0_u1_u0_n134 ) , .C2( u0_u1_u0_n135 ) , .C1( u0_u1_u0_n136 ) , .ZN( u0_u1_u0_n137 ) );
  OR4_X1 u0_u1_u0_U78 (.ZN( u0_out1_31 ) , .A4( u0_u1_u0_n155 ) , .A2( u0_u1_u0_n156 ) , .A1( u0_u1_u0_n157 ) , .A3( u0_u1_u0_n173 ) );
  AOI21_X1 u0_u1_u0_U79 (.A( u0_u1_u0_n138 ) , .B2( u0_u1_u0_n139 ) , .B1( u0_u1_u0_n140 ) , .ZN( u0_u1_u0_n157 ) );
  AND2_X1 u0_u1_u0_U8 (.A1( u0_u1_u0_n114 ) , .A2( u0_u1_u0_n121 ) , .ZN( u0_u1_u0_n146 ) );
  AOI21_X1 u0_u1_u0_U80 (.B2( u0_u1_u0_n141 ) , .B1( u0_u1_u0_n142 ) , .ZN( u0_u1_u0_n156 ) , .A( u0_u1_u0_n161 ) );
  OR4_X1 u0_u1_u0_U81 (.ZN( u0_out1_17 ) , .A4( u0_u1_u0_n122 ) , .A2( u0_u1_u0_n123 ) , .A1( u0_u1_u0_n124 ) , .A3( u0_u1_u0_n170 ) );
  AOI21_X1 u0_u1_u0_U82 (.B2( u0_u1_u0_n107 ) , .ZN( u0_u1_u0_n124 ) , .B1( u0_u1_u0_n128 ) , .A( u0_u1_u0_n161 ) );
  INV_X1 u0_u1_u0_U83 (.A( u0_u1_u0_n111 ) , .ZN( u0_u1_u0_n170 ) );
  AOI21_X1 u0_u1_u0_U84 (.B1( u0_u1_u0_n132 ) , .ZN( u0_u1_u0_n133 ) , .A( u0_u1_u0_n144 ) , .B2( u0_u1_u0_n166 ) );
  OAI22_X1 u0_u1_u0_U85 (.ZN( u0_u1_u0_n105 ) , .A2( u0_u1_u0_n132 ) , .B1( u0_u1_u0_n146 ) , .A1( u0_u1_u0_n147 ) , .B2( u0_u1_u0_n161 ) );
  NAND2_X1 u0_u1_u0_U86 (.ZN( u0_u1_u0_n110 ) , .A2( u0_u1_u0_n132 ) , .A1( u0_u1_u0_n145 ) );
  INV_X1 u0_u1_u0_U87 (.A( u0_u1_u0_n119 ) , .ZN( u0_u1_u0_n167 ) );
  NAND3_X1 u0_u1_u0_U88 (.ZN( u0_out1_23 ) , .A3( u0_u1_u0_n137 ) , .A1( u0_u1_u0_n168 ) , .A2( u0_u1_u0_n171 ) );
  NAND3_X1 u0_u1_u0_U89 (.A3( u0_u1_u0_n127 ) , .A2( u0_u1_u0_n128 ) , .ZN( u0_u1_u0_n135 ) , .A1( u0_u1_u0_n150 ) );
  AND2_X1 u0_u1_u0_U9 (.A1( u0_u1_u0_n131 ) , .ZN( u0_u1_u0_n141 ) , .A2( u0_u1_u0_n150 ) );
  NAND3_X1 u0_u1_u0_U90 (.ZN( u0_u1_u0_n117 ) , .A3( u0_u1_u0_n132 ) , .A2( u0_u1_u0_n139 ) , .A1( u0_u1_u0_n148 ) );
  NAND3_X1 u0_u1_u0_U91 (.ZN( u0_u1_u0_n109 ) , .A2( u0_u1_u0_n114 ) , .A3( u0_u1_u0_n140 ) , .A1( u0_u1_u0_n149 ) );
  NAND3_X1 u0_u1_u0_U92 (.ZN( u0_out1_9 ) , .A3( u0_u1_u0_n106 ) , .A2( u0_u1_u0_n171 ) , .A1( u0_u1_u0_n174 ) );
  NAND3_X1 u0_u1_u0_U93 (.A2( u0_u1_u0_n128 ) , .A1( u0_u1_u0_n132 ) , .A3( u0_u1_u0_n146 ) , .ZN( u0_u1_u0_n97 ) );
  NOR2_X1 u0_u1_u1_U10 (.A1( u0_u1_u1_n112 ) , .A2( u0_u1_u1_n116 ) , .ZN( u0_u1_u1_n118 ) );
  NAND3_X1 u0_u1_u1_U100 (.ZN( u0_u1_u1_n113 ) , .A1( u0_u1_u1_n120 ) , .A3( u0_u1_u1_n133 ) , .A2( u0_u1_u1_n155 ) );
  OAI21_X1 u0_u1_u1_U11 (.ZN( u0_u1_u1_n101 ) , .B1( u0_u1_u1_n141 ) , .A( u0_u1_u1_n146 ) , .B2( u0_u1_u1_n183 ) );
  AOI21_X1 u0_u1_u1_U12 (.B2( u0_u1_u1_n155 ) , .B1( u0_u1_u1_n156 ) , .ZN( u0_u1_u1_n157 ) , .A( u0_u1_u1_n174 ) );
  OR4_X1 u0_u1_u1_U13 (.A4( u0_u1_u1_n106 ) , .A3( u0_u1_u1_n107 ) , .ZN( u0_u1_u1_n108 ) , .A1( u0_u1_u1_n117 ) , .A2( u0_u1_u1_n184 ) );
  AOI21_X1 u0_u1_u1_U14 (.ZN( u0_u1_u1_n106 ) , .A( u0_u1_u1_n112 ) , .B1( u0_u1_u1_n154 ) , .B2( u0_u1_u1_n156 ) );
  INV_X1 u0_u1_u1_U15 (.A( u0_u1_u1_n101 ) , .ZN( u0_u1_u1_n184 ) );
  AOI21_X1 u0_u1_u1_U16 (.ZN( u0_u1_u1_n107 ) , .B1( u0_u1_u1_n134 ) , .B2( u0_u1_u1_n149 ) , .A( u0_u1_u1_n174 ) );
  NAND2_X1 u0_u1_u1_U17 (.ZN( u0_u1_u1_n140 ) , .A2( u0_u1_u1_n150 ) , .A1( u0_u1_u1_n155 ) );
  NAND2_X1 u0_u1_u1_U18 (.A1( u0_u1_u1_n131 ) , .ZN( u0_u1_u1_n147 ) , .A2( u0_u1_u1_n153 ) );
  INV_X1 u0_u1_u1_U19 (.A( u0_u1_u1_n139 ) , .ZN( u0_u1_u1_n174 ) );
  INV_X1 u0_u1_u1_U20 (.A( u0_u1_u1_n112 ) , .ZN( u0_u1_u1_n171 ) );
  NAND2_X1 u0_u1_u1_U21 (.ZN( u0_u1_u1_n141 ) , .A1( u0_u1_u1_n153 ) , .A2( u0_u1_u1_n156 ) );
  AND2_X1 u0_u1_u1_U22 (.A1( u0_u1_u1_n123 ) , .ZN( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n161 ) );
  NAND2_X1 u0_u1_u1_U23 (.A2( u0_u1_u1_n115 ) , .A1( u0_u1_u1_n116 ) , .ZN( u0_u1_u1_n148 ) );
  NAND2_X1 u0_u1_u1_U24 (.A2( u0_u1_u1_n133 ) , .A1( u0_u1_u1_n135 ) , .ZN( u0_u1_u1_n159 ) );
  NAND2_X1 u0_u1_u1_U25 (.A2( u0_u1_u1_n115 ) , .A1( u0_u1_u1_n120 ) , .ZN( u0_u1_u1_n132 ) );
  INV_X1 u0_u1_u1_U26 (.A( u0_u1_u1_n154 ) , .ZN( u0_u1_u1_n178 ) );
  INV_X1 u0_u1_u1_U27 (.A( u0_u1_u1_n151 ) , .ZN( u0_u1_u1_n183 ) );
  AND2_X1 u0_u1_u1_U28 (.A1( u0_u1_u1_n129 ) , .A2( u0_u1_u1_n133 ) , .ZN( u0_u1_u1_n149 ) );
  INV_X1 u0_u1_u1_U29 (.A( u0_u1_u1_n131 ) , .ZN( u0_u1_u1_n180 ) );
  INV_X1 u0_u1_u1_U3 (.A( u0_u1_u1_n159 ) , .ZN( u0_u1_u1_n182 ) );
  AOI221_X1 u0_u1_u1_U30 (.B1( u0_u1_u1_n140 ) , .ZN( u0_u1_u1_n167 ) , .B2( u0_u1_u1_n172 ) , .C2( u0_u1_u1_n175 ) , .C1( u0_u1_u1_n178 ) , .A( u0_u1_u1_n188 ) );
  INV_X1 u0_u1_u1_U31 (.ZN( u0_u1_u1_n188 ) , .A( u0_u1_u1_n97 ) );
  AOI211_X1 u0_u1_u1_U32 (.A( u0_u1_u1_n118 ) , .C1( u0_u1_u1_n132 ) , .C2( u0_u1_u1_n139 ) , .B( u0_u1_u1_n96 ) , .ZN( u0_u1_u1_n97 ) );
  AOI21_X1 u0_u1_u1_U33 (.B2( u0_u1_u1_n121 ) , .B1( u0_u1_u1_n135 ) , .A( u0_u1_u1_n152 ) , .ZN( u0_u1_u1_n96 ) );
  OAI221_X1 u0_u1_u1_U34 (.A( u0_u1_u1_n119 ) , .C2( u0_u1_u1_n129 ) , .ZN( u0_u1_u1_n138 ) , .B2( u0_u1_u1_n152 ) , .C1( u0_u1_u1_n174 ) , .B1( u0_u1_u1_n187 ) );
  INV_X1 u0_u1_u1_U35 (.A( u0_u1_u1_n148 ) , .ZN( u0_u1_u1_n187 ) );
  AOI211_X1 u0_u1_u1_U36 (.B( u0_u1_u1_n117 ) , .A( u0_u1_u1_n118 ) , .ZN( u0_u1_u1_n119 ) , .C2( u0_u1_u1_n146 ) , .C1( u0_u1_u1_n159 ) );
  NOR2_X1 u0_u1_u1_U37 (.A1( u0_u1_u1_n168 ) , .A2( u0_u1_u1_n176 ) , .ZN( u0_u1_u1_n98 ) );
  AOI211_X1 u0_u1_u1_U38 (.B( u0_u1_u1_n162 ) , .A( u0_u1_u1_n163 ) , .C2( u0_u1_u1_n164 ) , .ZN( u0_u1_u1_n165 ) , .C1( u0_u1_u1_n171 ) );
  AOI21_X1 u0_u1_u1_U39 (.A( u0_u1_u1_n160 ) , .B2( u0_u1_u1_n161 ) , .ZN( u0_u1_u1_n162 ) , .B1( u0_u1_u1_n182 ) );
  AOI221_X1 u0_u1_u1_U4 (.A( u0_u1_u1_n138 ) , .C2( u0_u1_u1_n139 ) , .C1( u0_u1_u1_n140 ) , .B2( u0_u1_u1_n141 ) , .ZN( u0_u1_u1_n142 ) , .B1( u0_u1_u1_n175 ) );
  OR2_X1 u0_u1_u1_U40 (.A2( u0_u1_u1_n157 ) , .A1( u0_u1_u1_n158 ) , .ZN( u0_u1_u1_n163 ) );
  OAI21_X1 u0_u1_u1_U41 (.B2( u0_u1_u1_n123 ) , .ZN( u0_u1_u1_n145 ) , .B1( u0_u1_u1_n160 ) , .A( u0_u1_u1_n185 ) );
  INV_X1 u0_u1_u1_U42 (.A( u0_u1_u1_n122 ) , .ZN( u0_u1_u1_n185 ) );
  AOI21_X1 u0_u1_u1_U43 (.B2( u0_u1_u1_n120 ) , .B1( u0_u1_u1_n121 ) , .ZN( u0_u1_u1_n122 ) , .A( u0_u1_u1_n128 ) );
  NAND2_X1 u0_u1_u1_U44 (.A1( u0_u1_u1_n128 ) , .ZN( u0_u1_u1_n146 ) , .A2( u0_u1_u1_n160 ) );
  NAND2_X1 u0_u1_u1_U45 (.A2( u0_u1_u1_n112 ) , .ZN( u0_u1_u1_n139 ) , .A1( u0_u1_u1_n152 ) );
  NAND2_X1 u0_u1_u1_U46 (.A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n156 ) , .A2( u0_u1_u1_n99 ) );
  NOR2_X1 u0_u1_u1_U47 (.ZN( u0_u1_u1_n117 ) , .A1( u0_u1_u1_n121 ) , .A2( u0_u1_u1_n160 ) );
  AOI21_X1 u0_u1_u1_U48 (.A( u0_u1_u1_n128 ) , .B2( u0_u1_u1_n129 ) , .ZN( u0_u1_u1_n130 ) , .B1( u0_u1_u1_n150 ) );
  NAND2_X1 u0_u1_u1_U49 (.ZN( u0_u1_u1_n112 ) , .A1( u0_u1_u1_n169 ) , .A2( u0_u1_u1_n170 ) );
  AOI211_X1 u0_u1_u1_U5 (.ZN( u0_u1_u1_n124 ) , .A( u0_u1_u1_n138 ) , .C2( u0_u1_u1_n139 ) , .B( u0_u1_u1_n145 ) , .C1( u0_u1_u1_n147 ) );
  NAND2_X1 u0_u1_u1_U50 (.ZN( u0_u1_u1_n129 ) , .A2( u0_u1_u1_n95 ) , .A1( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U51 (.A1( u0_u1_u1_n102 ) , .ZN( u0_u1_u1_n154 ) , .A2( u0_u1_u1_n99 ) );
  NAND2_X1 u0_u1_u1_U52 (.A2( u0_u1_u1_n100 ) , .ZN( u0_u1_u1_n135 ) , .A1( u0_u1_u1_n99 ) );
  AOI21_X1 u0_u1_u1_U53 (.A( u0_u1_u1_n152 ) , .B2( u0_u1_u1_n153 ) , .B1( u0_u1_u1_n154 ) , .ZN( u0_u1_u1_n158 ) );
  INV_X1 u0_u1_u1_U54 (.A( u0_u1_u1_n160 ) , .ZN( u0_u1_u1_n175 ) );
  NAND2_X1 u0_u1_u1_U55 (.A1( u0_u1_u1_n100 ) , .ZN( u0_u1_u1_n116 ) , .A2( u0_u1_u1_n95 ) );
  NAND2_X1 u0_u1_u1_U56 (.A1( u0_u1_u1_n102 ) , .ZN( u0_u1_u1_n131 ) , .A2( u0_u1_u1_n95 ) );
  NAND2_X1 u0_u1_u1_U57 (.A2( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n121 ) , .A1( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U58 (.A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n153 ) , .A2( u0_u1_u1_n98 ) );
  NAND2_X1 u0_u1_u1_U59 (.A2( u0_u1_u1_n104 ) , .A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n133 ) );
  AOI22_X1 u0_u1_u1_U6 (.B2( u0_u1_u1_n113 ) , .A2( u0_u1_u1_n114 ) , .ZN( u0_u1_u1_n125 ) , .A1( u0_u1_u1_n171 ) , .B1( u0_u1_u1_n173 ) );
  NAND2_X1 u0_u1_u1_U60 (.ZN( u0_u1_u1_n150 ) , .A2( u0_u1_u1_n98 ) , .A1( u0_u1_u1_n99 ) );
  NAND2_X1 u0_u1_u1_U61 (.A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n155 ) , .A2( u0_u1_u1_n95 ) );
  OAI21_X1 u0_u1_u1_U62 (.ZN( u0_u1_u1_n109 ) , .B1( u0_u1_u1_n129 ) , .B2( u0_u1_u1_n160 ) , .A( u0_u1_u1_n167 ) );
  NAND2_X1 u0_u1_u1_U63 (.A2( u0_u1_u1_n100 ) , .A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n120 ) );
  NAND2_X1 u0_u1_u1_U64 (.A1( u0_u1_u1_n102 ) , .A2( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n115 ) );
  NAND2_X1 u0_u1_u1_U65 (.A2( u0_u1_u1_n100 ) , .A1( u0_u1_u1_n104 ) , .ZN( u0_u1_u1_n151 ) );
  NAND2_X1 u0_u1_u1_U66 (.A2( u0_u1_u1_n103 ) , .A1( u0_u1_u1_n105 ) , .ZN( u0_u1_u1_n161 ) );
  INV_X1 u0_u1_u1_U67 (.A( u0_u1_u1_n152 ) , .ZN( u0_u1_u1_n173 ) );
  INV_X1 u0_u1_u1_U68 (.A( u0_u1_u1_n128 ) , .ZN( u0_u1_u1_n172 ) );
  NAND2_X1 u0_u1_u1_U69 (.A2( u0_u1_u1_n102 ) , .A1( u0_u1_u1_n103 ) , .ZN( u0_u1_u1_n123 ) );
  NAND2_X1 u0_u1_u1_U7 (.ZN( u0_u1_u1_n114 ) , .A1( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n156 ) );
  NOR2_X1 u0_u1_u1_U70 (.A2( u0_u1_X_7 ) , .A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n95 ) );
  NOR2_X1 u0_u1_u1_U71 (.A1( u0_u1_X_12 ) , .A2( u0_u1_X_9 ) , .ZN( u0_u1_u1_n100 ) );
  NOR2_X1 u0_u1_u1_U72 (.A2( u0_u1_X_8 ) , .A1( u0_u1_u1_n177 ) , .ZN( u0_u1_u1_n99 ) );
  NOR2_X1 u0_u1_u1_U73 (.A2( u0_u1_X_12 ) , .ZN( u0_u1_u1_n102 ) , .A1( u0_u1_u1_n176 ) );
  NOR2_X1 u0_u1_u1_U74 (.A2( u0_u1_X_9 ) , .ZN( u0_u1_u1_n105 ) , .A1( u0_u1_u1_n168 ) );
  NAND2_X1 u0_u1_u1_U75 (.A1( u0_u1_X_10 ) , .ZN( u0_u1_u1_n160 ) , .A2( u0_u1_u1_n169 ) );
  NAND2_X1 u0_u1_u1_U76 (.A2( u0_u1_X_10 ) , .A1( u0_u1_X_11 ) , .ZN( u0_u1_u1_n152 ) );
  NAND2_X1 u0_u1_u1_U77 (.A1( u0_u1_X_11 ) , .ZN( u0_u1_u1_n128 ) , .A2( u0_u1_u1_n170 ) );
  AND2_X1 u0_u1_u1_U78 (.A2( u0_u1_X_7 ) , .A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n104 ) );
  AND2_X1 u0_u1_u1_U79 (.A1( u0_u1_X_8 ) , .ZN( u0_u1_u1_n103 ) , .A2( u0_u1_u1_n177 ) );
  AOI22_X1 u0_u1_u1_U8 (.B2( u0_u1_u1_n136 ) , .A2( u0_u1_u1_n137 ) , .ZN( u0_u1_u1_n143 ) , .A1( u0_u1_u1_n171 ) , .B1( u0_u1_u1_n173 ) );
  INV_X1 u0_u1_u1_U80 (.A( u0_u1_X_10 ) , .ZN( u0_u1_u1_n170 ) );
  INV_X1 u0_u1_u1_U81 (.A( u0_u1_X_9 ) , .ZN( u0_u1_u1_n176 ) );
  INV_X1 u0_u1_u1_U82 (.A( u0_u1_X_11 ) , .ZN( u0_u1_u1_n169 ) );
  INV_X1 u0_u1_u1_U83 (.A( u0_u1_X_12 ) , .ZN( u0_u1_u1_n168 ) );
  INV_X1 u0_u1_u1_U84 (.A( u0_u1_X_7 ) , .ZN( u0_u1_u1_n177 ) );
  NAND4_X1 u0_u1_u1_U85 (.ZN( u0_out1_28 ) , .A4( u0_u1_u1_n124 ) , .A3( u0_u1_u1_n125 ) , .A2( u0_u1_u1_n126 ) , .A1( u0_u1_u1_n127 ) );
  OAI21_X1 u0_u1_u1_U86 (.ZN( u0_u1_u1_n127 ) , .B2( u0_u1_u1_n139 ) , .B1( u0_u1_u1_n175 ) , .A( u0_u1_u1_n183 ) );
  OAI21_X1 u0_u1_u1_U87 (.ZN( u0_u1_u1_n126 ) , .B2( u0_u1_u1_n140 ) , .A( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n178 ) );
  NAND4_X1 u0_u1_u1_U88 (.ZN( u0_out1_18 ) , .A4( u0_u1_u1_n165 ) , .A3( u0_u1_u1_n166 ) , .A1( u0_u1_u1_n167 ) , .A2( u0_u1_u1_n186 ) );
  AOI22_X1 u0_u1_u1_U89 (.B2( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n147 ) , .A2( u0_u1_u1_n148 ) , .ZN( u0_u1_u1_n166 ) , .A1( u0_u1_u1_n172 ) );
  INV_X1 u0_u1_u1_U9 (.A( u0_u1_u1_n147 ) , .ZN( u0_u1_u1_n181 ) );
  INV_X1 u0_u1_u1_U90 (.A( u0_u1_u1_n145 ) , .ZN( u0_u1_u1_n186 ) );
  NAND4_X1 u0_u1_u1_U91 (.ZN( u0_out1_2 ) , .A4( u0_u1_u1_n142 ) , .A3( u0_u1_u1_n143 ) , .A2( u0_u1_u1_n144 ) , .A1( u0_u1_u1_n179 ) );
  INV_X1 u0_u1_u1_U92 (.A( u0_u1_u1_n130 ) , .ZN( u0_u1_u1_n179 ) );
  OAI21_X1 u0_u1_u1_U93 (.B2( u0_u1_u1_n132 ) , .ZN( u0_u1_u1_n144 ) , .A( u0_u1_u1_n146 ) , .B1( u0_u1_u1_n180 ) );
  OR4_X1 u0_u1_u1_U94 (.ZN( u0_out1_13 ) , .A4( u0_u1_u1_n108 ) , .A3( u0_u1_u1_n109 ) , .A2( u0_u1_u1_n110 ) , .A1( u0_u1_u1_n111 ) );
  AOI21_X1 u0_u1_u1_U95 (.ZN( u0_u1_u1_n111 ) , .A( u0_u1_u1_n128 ) , .B2( u0_u1_u1_n131 ) , .B1( u0_u1_u1_n135 ) );
  AOI21_X1 u0_u1_u1_U96 (.ZN( u0_u1_u1_n110 ) , .A( u0_u1_u1_n116 ) , .B1( u0_u1_u1_n152 ) , .B2( u0_u1_u1_n160 ) );
  NAND3_X1 u0_u1_u1_U97 (.A3( u0_u1_u1_n149 ) , .A2( u0_u1_u1_n150 ) , .A1( u0_u1_u1_n151 ) , .ZN( u0_u1_u1_n164 ) );
  NAND3_X1 u0_u1_u1_U98 (.A3( u0_u1_u1_n134 ) , .A2( u0_u1_u1_n135 ) , .ZN( u0_u1_u1_n136 ) , .A1( u0_u1_u1_n151 ) );
  NAND3_X1 u0_u1_u1_U99 (.A1( u0_u1_u1_n133 ) , .ZN( u0_u1_u1_n137 ) , .A2( u0_u1_u1_n154 ) , .A3( u0_u1_u1_n181 ) );
  OAI22_X1 u0_u1_u2_U10 (.ZN( u0_u1_u2_n109 ) , .A2( u0_u1_u2_n113 ) , .B2( u0_u1_u2_n133 ) , .B1( u0_u1_u2_n167 ) , .A1( u0_u1_u2_n168 ) );
  NAND3_X1 u0_u1_u2_U100 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n104 ) , .A3( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n98 ) );
  OAI22_X1 u0_u1_u2_U11 (.B1( u0_u1_u2_n151 ) , .A2( u0_u1_u2_n152 ) , .A1( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n160 ) , .B2( u0_u1_u2_n168 ) );
  NOR3_X1 u0_u1_u2_U12 (.A1( u0_u1_u2_n150 ) , .ZN( u0_u1_u2_n151 ) , .A3( u0_u1_u2_n175 ) , .A2( u0_u1_u2_n188 ) );
  AOI21_X1 u0_u1_u2_U13 (.ZN( u0_u1_u2_n144 ) , .B2( u0_u1_u2_n155 ) , .A( u0_u1_u2_n172 ) , .B1( u0_u1_u2_n185 ) );
  AOI21_X1 u0_u1_u2_U14 (.B2( u0_u1_u2_n143 ) , .ZN( u0_u1_u2_n145 ) , .B1( u0_u1_u2_n152 ) , .A( u0_u1_u2_n171 ) );
  AOI21_X1 u0_u1_u2_U15 (.B2( u0_u1_u2_n120 ) , .B1( u0_u1_u2_n121 ) , .ZN( u0_u1_u2_n126 ) , .A( u0_u1_u2_n167 ) );
  INV_X1 u0_u1_u2_U16 (.A( u0_u1_u2_n156 ) , .ZN( u0_u1_u2_n171 ) );
  INV_X1 u0_u1_u2_U17 (.A( u0_u1_u2_n120 ) , .ZN( u0_u1_u2_n188 ) );
  NAND2_X1 u0_u1_u2_U18 (.A2( u0_u1_u2_n122 ) , .ZN( u0_u1_u2_n150 ) , .A1( u0_u1_u2_n152 ) );
  INV_X1 u0_u1_u2_U19 (.A( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n170 ) );
  INV_X1 u0_u1_u2_U20 (.A( u0_u1_u2_n137 ) , .ZN( u0_u1_u2_n173 ) );
  NAND2_X1 u0_u1_u2_U21 (.A1( u0_u1_u2_n132 ) , .A2( u0_u1_u2_n139 ) , .ZN( u0_u1_u2_n157 ) );
  INV_X1 u0_u1_u2_U22 (.A( u0_u1_u2_n113 ) , .ZN( u0_u1_u2_n178 ) );
  INV_X1 u0_u1_u2_U23 (.A( u0_u1_u2_n139 ) , .ZN( u0_u1_u2_n175 ) );
  INV_X1 u0_u1_u2_U24 (.A( u0_u1_u2_n155 ) , .ZN( u0_u1_u2_n181 ) );
  INV_X1 u0_u1_u2_U25 (.A( u0_u1_u2_n119 ) , .ZN( u0_u1_u2_n177 ) );
  INV_X1 u0_u1_u2_U26 (.A( u0_u1_u2_n116 ) , .ZN( u0_u1_u2_n180 ) );
  INV_X1 u0_u1_u2_U27 (.A( u0_u1_u2_n131 ) , .ZN( u0_u1_u2_n179 ) );
  INV_X1 u0_u1_u2_U28 (.A( u0_u1_u2_n154 ) , .ZN( u0_u1_u2_n176 ) );
  NAND2_X1 u0_u1_u2_U29 (.A2( u0_u1_u2_n116 ) , .A1( u0_u1_u2_n117 ) , .ZN( u0_u1_u2_n118 ) );
  NOR2_X1 u0_u1_u2_U3 (.ZN( u0_u1_u2_n121 ) , .A2( u0_u1_u2_n177 ) , .A1( u0_u1_u2_n180 ) );
  INV_X1 u0_u1_u2_U30 (.A( u0_u1_u2_n132 ) , .ZN( u0_u1_u2_n182 ) );
  INV_X1 u0_u1_u2_U31 (.A( u0_u1_u2_n158 ) , .ZN( u0_u1_u2_n183 ) );
  OAI21_X1 u0_u1_u2_U32 (.A( u0_u1_u2_n156 ) , .B1( u0_u1_u2_n157 ) , .ZN( u0_u1_u2_n158 ) , .B2( u0_u1_u2_n179 ) );
  NOR2_X1 u0_u1_u2_U33 (.ZN( u0_u1_u2_n156 ) , .A1( u0_u1_u2_n166 ) , .A2( u0_u1_u2_n169 ) );
  NOR2_X1 u0_u1_u2_U34 (.A2( u0_u1_u2_n114 ) , .ZN( u0_u1_u2_n137 ) , .A1( u0_u1_u2_n140 ) );
  NOR2_X1 u0_u1_u2_U35 (.A2( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n153 ) , .A1( u0_u1_u2_n156 ) );
  AOI211_X1 u0_u1_u2_U36 (.ZN( u0_u1_u2_n130 ) , .C1( u0_u1_u2_n138 ) , .C2( u0_u1_u2_n179 ) , .B( u0_u1_u2_n96 ) , .A( u0_u1_u2_n97 ) );
  OAI22_X1 u0_u1_u2_U37 (.B1( u0_u1_u2_n133 ) , .A2( u0_u1_u2_n137 ) , .A1( u0_u1_u2_n152 ) , .B2( u0_u1_u2_n168 ) , .ZN( u0_u1_u2_n97 ) );
  OAI221_X1 u0_u1_u2_U38 (.B1( u0_u1_u2_n113 ) , .C1( u0_u1_u2_n132 ) , .A( u0_u1_u2_n149 ) , .B2( u0_u1_u2_n171 ) , .C2( u0_u1_u2_n172 ) , .ZN( u0_u1_u2_n96 ) );
  OAI221_X1 u0_u1_u2_U39 (.A( u0_u1_u2_n115 ) , .C2( u0_u1_u2_n123 ) , .B2( u0_u1_u2_n143 ) , .B1( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n163 ) , .C1( u0_u1_u2_n168 ) );
  INV_X1 u0_u1_u2_U4 (.A( u0_u1_u2_n134 ) , .ZN( u0_u1_u2_n185 ) );
  OAI21_X1 u0_u1_u2_U40 (.A( u0_u1_u2_n114 ) , .ZN( u0_u1_u2_n115 ) , .B1( u0_u1_u2_n176 ) , .B2( u0_u1_u2_n178 ) );
  OAI221_X1 u0_u1_u2_U41 (.A( u0_u1_u2_n135 ) , .B2( u0_u1_u2_n136 ) , .B1( u0_u1_u2_n137 ) , .ZN( u0_u1_u2_n162 ) , .C2( u0_u1_u2_n167 ) , .C1( u0_u1_u2_n185 ) );
  AND3_X1 u0_u1_u2_U42 (.A3( u0_u1_u2_n131 ) , .A2( u0_u1_u2_n132 ) , .A1( u0_u1_u2_n133 ) , .ZN( u0_u1_u2_n136 ) );
  AOI22_X1 u0_u1_u2_U43 (.ZN( u0_u1_u2_n135 ) , .B1( u0_u1_u2_n140 ) , .A1( u0_u1_u2_n156 ) , .B2( u0_u1_u2_n180 ) , .A2( u0_u1_u2_n188 ) );
  AOI21_X1 u0_u1_u2_U44 (.ZN( u0_u1_u2_n149 ) , .B1( u0_u1_u2_n173 ) , .B2( u0_u1_u2_n188 ) , .A( u0_u1_u2_n95 ) );
  AND3_X1 u0_u1_u2_U45 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n104 ) , .A3( u0_u1_u2_n156 ) , .ZN( u0_u1_u2_n95 ) );
  OAI21_X1 u0_u1_u2_U46 (.A( u0_u1_u2_n101 ) , .B2( u0_u1_u2_n121 ) , .B1( u0_u1_u2_n153 ) , .ZN( u0_u1_u2_n164 ) );
  NAND2_X1 u0_u1_u2_U47 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n107 ) , .ZN( u0_u1_u2_n155 ) );
  NAND2_X1 u0_u1_u2_U48 (.A2( u0_u1_u2_n105 ) , .A1( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n143 ) );
  NAND2_X1 u0_u1_u2_U49 (.A1( u0_u1_u2_n104 ) , .A2( u0_u1_u2_n106 ) , .ZN( u0_u1_u2_n152 ) );
  INV_X1 u0_u1_u2_U5 (.A( u0_u1_u2_n150 ) , .ZN( u0_u1_u2_n184 ) );
  NAND2_X1 u0_u1_u2_U50 (.A1( u0_u1_u2_n100 ) , .A2( u0_u1_u2_n105 ) , .ZN( u0_u1_u2_n132 ) );
  INV_X1 u0_u1_u2_U51 (.A( u0_u1_u2_n140 ) , .ZN( u0_u1_u2_n168 ) );
  INV_X1 u0_u1_u2_U52 (.A( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n167 ) );
  OAI21_X1 u0_u1_u2_U53 (.A( u0_u1_u2_n141 ) , .B2( u0_u1_u2_n142 ) , .ZN( u0_u1_u2_n146 ) , .B1( u0_u1_u2_n153 ) );
  OAI21_X1 u0_u1_u2_U54 (.A( u0_u1_u2_n140 ) , .ZN( u0_u1_u2_n141 ) , .B1( u0_u1_u2_n176 ) , .B2( u0_u1_u2_n177 ) );
  NOR3_X1 u0_u1_u2_U55 (.ZN( u0_u1_u2_n142 ) , .A3( u0_u1_u2_n175 ) , .A2( u0_u1_u2_n178 ) , .A1( u0_u1_u2_n181 ) );
  NAND2_X1 u0_u1_u2_U56 (.A1( u0_u1_u2_n102 ) , .A2( u0_u1_u2_n106 ) , .ZN( u0_u1_u2_n113 ) );
  NAND2_X1 u0_u1_u2_U57 (.A1( u0_u1_u2_n106 ) , .A2( u0_u1_u2_n107 ) , .ZN( u0_u1_u2_n131 ) );
  NAND2_X1 u0_u1_u2_U58 (.A1( u0_u1_u2_n103 ) , .A2( u0_u1_u2_n107 ) , .ZN( u0_u1_u2_n139 ) );
  NAND2_X1 u0_u1_u2_U59 (.A1( u0_u1_u2_n103 ) , .A2( u0_u1_u2_n105 ) , .ZN( u0_u1_u2_n133 ) );
  NOR4_X1 u0_u1_u2_U6 (.A4( u0_u1_u2_n124 ) , .A3( u0_u1_u2_n125 ) , .A2( u0_u1_u2_n126 ) , .A1( u0_u1_u2_n127 ) , .ZN( u0_u1_u2_n128 ) );
  NAND2_X1 u0_u1_u2_U60 (.A1( u0_u1_u2_n102 ) , .A2( u0_u1_u2_n103 ) , .ZN( u0_u1_u2_n154 ) );
  NAND2_X1 u0_u1_u2_U61 (.A2( u0_u1_u2_n103 ) , .A1( u0_u1_u2_n104 ) , .ZN( u0_u1_u2_n119 ) );
  NAND2_X1 u0_u1_u2_U62 (.A2( u0_u1_u2_n107 ) , .A1( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n123 ) );
  NAND2_X1 u0_u1_u2_U63 (.A1( u0_u1_u2_n104 ) , .A2( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n122 ) );
  INV_X1 u0_u1_u2_U64 (.A( u0_u1_u2_n114 ) , .ZN( u0_u1_u2_n172 ) );
  NAND2_X1 u0_u1_u2_U65 (.A2( u0_u1_u2_n100 ) , .A1( u0_u1_u2_n102 ) , .ZN( u0_u1_u2_n116 ) );
  NAND2_X1 u0_u1_u2_U66 (.A1( u0_u1_u2_n102 ) , .A2( u0_u1_u2_n108 ) , .ZN( u0_u1_u2_n120 ) );
  NAND2_X1 u0_u1_u2_U67 (.A2( u0_u1_u2_n105 ) , .A1( u0_u1_u2_n106 ) , .ZN( u0_u1_u2_n117 ) );
  INV_X1 u0_u1_u2_U68 (.ZN( u0_u1_u2_n187 ) , .A( u0_u1_u2_n99 ) );
  OAI21_X1 u0_u1_u2_U69 (.B1( u0_u1_u2_n137 ) , .B2( u0_u1_u2_n143 ) , .A( u0_u1_u2_n98 ) , .ZN( u0_u1_u2_n99 ) );
  AOI21_X1 u0_u1_u2_U7 (.B2( u0_u1_u2_n119 ) , .ZN( u0_u1_u2_n127 ) , .A( u0_u1_u2_n137 ) , .B1( u0_u1_u2_n155 ) );
  NOR2_X1 u0_u1_u2_U70 (.A2( u0_u1_X_16 ) , .ZN( u0_u1_u2_n140 ) , .A1( u0_u1_u2_n166 ) );
  NOR2_X1 u0_u1_u2_U71 (.A2( u0_u1_X_13 ) , .A1( u0_u1_X_14 ) , .ZN( u0_u1_u2_n100 ) );
  NOR2_X1 u0_u1_u2_U72 (.A2( u0_u1_X_16 ) , .A1( u0_u1_X_17 ) , .ZN( u0_u1_u2_n138 ) );
  NOR2_X1 u0_u1_u2_U73 (.A2( u0_u1_X_15 ) , .A1( u0_u1_X_18 ) , .ZN( u0_u1_u2_n104 ) );
  NOR2_X1 u0_u1_u2_U74 (.A2( u0_u1_X_14 ) , .ZN( u0_u1_u2_n103 ) , .A1( u0_u1_u2_n174 ) );
  NOR2_X1 u0_u1_u2_U75 (.A2( u0_u1_X_15 ) , .ZN( u0_u1_u2_n102 ) , .A1( u0_u1_u2_n165 ) );
  NOR2_X1 u0_u1_u2_U76 (.A2( u0_u1_X_17 ) , .ZN( u0_u1_u2_n114 ) , .A1( u0_u1_u2_n169 ) );
  AND2_X1 u0_u1_u2_U77 (.A1( u0_u1_X_15 ) , .ZN( u0_u1_u2_n105 ) , .A2( u0_u1_u2_n165 ) );
  AND2_X1 u0_u1_u2_U78 (.A2( u0_u1_X_15 ) , .A1( u0_u1_X_18 ) , .ZN( u0_u1_u2_n107 ) );
  AND2_X1 u0_u1_u2_U79 (.A1( u0_u1_X_14 ) , .ZN( u0_u1_u2_n106 ) , .A2( u0_u1_u2_n174 ) );
  AOI21_X1 u0_u1_u2_U8 (.ZN( u0_u1_u2_n124 ) , .B1( u0_u1_u2_n131 ) , .B2( u0_u1_u2_n143 ) , .A( u0_u1_u2_n172 ) );
  AND2_X1 u0_u1_u2_U80 (.A1( u0_u1_X_13 ) , .A2( u0_u1_X_14 ) , .ZN( u0_u1_u2_n108 ) );
  INV_X1 u0_u1_u2_U81 (.A( u0_u1_X_16 ) , .ZN( u0_u1_u2_n169 ) );
  INV_X1 u0_u1_u2_U82 (.A( u0_u1_X_17 ) , .ZN( u0_u1_u2_n166 ) );
  INV_X1 u0_u1_u2_U83 (.A( u0_u1_X_13 ) , .ZN( u0_u1_u2_n174 ) );
  INV_X1 u0_u1_u2_U84 (.A( u0_u1_X_18 ) , .ZN( u0_u1_u2_n165 ) );
  NAND4_X1 u0_u1_u2_U85 (.ZN( u0_out1_30 ) , .A4( u0_u1_u2_n147 ) , .A3( u0_u1_u2_n148 ) , .A2( u0_u1_u2_n149 ) , .A1( u0_u1_u2_n187 ) );
  NOR3_X1 u0_u1_u2_U86 (.A3( u0_u1_u2_n144 ) , .A2( u0_u1_u2_n145 ) , .A1( u0_u1_u2_n146 ) , .ZN( u0_u1_u2_n147 ) );
  AOI21_X1 u0_u1_u2_U87 (.B2( u0_u1_u2_n138 ) , .ZN( u0_u1_u2_n148 ) , .A( u0_u1_u2_n162 ) , .B1( u0_u1_u2_n182 ) );
  NAND4_X1 u0_u1_u2_U88 (.ZN( u0_out1_24 ) , .A4( u0_u1_u2_n111 ) , .A3( u0_u1_u2_n112 ) , .A1( u0_u1_u2_n130 ) , .A2( u0_u1_u2_n187 ) );
  AOI221_X1 u0_u1_u2_U89 (.A( u0_u1_u2_n109 ) , .B1( u0_u1_u2_n110 ) , .ZN( u0_u1_u2_n111 ) , .C1( u0_u1_u2_n134 ) , .C2( u0_u1_u2_n170 ) , .B2( u0_u1_u2_n173 ) );
  AOI21_X1 u0_u1_u2_U9 (.B2( u0_u1_u2_n123 ) , .ZN( u0_u1_u2_n125 ) , .A( u0_u1_u2_n171 ) , .B1( u0_u1_u2_n184 ) );
  AOI21_X1 u0_u1_u2_U90 (.ZN( u0_u1_u2_n112 ) , .B2( u0_u1_u2_n156 ) , .A( u0_u1_u2_n164 ) , .B1( u0_u1_u2_n181 ) );
  NAND4_X1 u0_u1_u2_U91 (.ZN( u0_out1_16 ) , .A4( u0_u1_u2_n128 ) , .A3( u0_u1_u2_n129 ) , .A1( u0_u1_u2_n130 ) , .A2( u0_u1_u2_n186 ) );
  AOI22_X1 u0_u1_u2_U92 (.A2( u0_u1_u2_n118 ) , .ZN( u0_u1_u2_n129 ) , .A1( u0_u1_u2_n140 ) , .B1( u0_u1_u2_n157 ) , .B2( u0_u1_u2_n170 ) );
  INV_X1 u0_u1_u2_U93 (.A( u0_u1_u2_n163 ) , .ZN( u0_u1_u2_n186 ) );
  OR4_X1 u0_u1_u2_U94 (.ZN( u0_out1_6 ) , .A4( u0_u1_u2_n161 ) , .A3( u0_u1_u2_n162 ) , .A2( u0_u1_u2_n163 ) , .A1( u0_u1_u2_n164 ) );
  OR3_X1 u0_u1_u2_U95 (.A2( u0_u1_u2_n159 ) , .A1( u0_u1_u2_n160 ) , .ZN( u0_u1_u2_n161 ) , .A3( u0_u1_u2_n183 ) );
  AOI21_X1 u0_u1_u2_U96 (.B2( u0_u1_u2_n154 ) , .B1( u0_u1_u2_n155 ) , .ZN( u0_u1_u2_n159 ) , .A( u0_u1_u2_n167 ) );
  NAND3_X1 u0_u1_u2_U97 (.A2( u0_u1_u2_n117 ) , .A1( u0_u1_u2_n122 ) , .A3( u0_u1_u2_n123 ) , .ZN( u0_u1_u2_n134 ) );
  NAND3_X1 u0_u1_u2_U98 (.ZN( u0_u1_u2_n110 ) , .A2( u0_u1_u2_n131 ) , .A3( u0_u1_u2_n139 ) , .A1( u0_u1_u2_n154 ) );
  NAND3_X1 u0_u1_u2_U99 (.A2( u0_u1_u2_n100 ) , .ZN( u0_u1_u2_n101 ) , .A1( u0_u1_u2_n104 ) , .A3( u0_u1_u2_n114 ) );
  AOI22_X1 u0_u1_u6_U10 (.A2( u0_u1_u6_n151 ) , .B2( u0_u1_u6_n161 ) , .A1( u0_u1_u6_n167 ) , .B1( u0_u1_u6_n170 ) , .ZN( u0_u1_u6_n89 ) );
  AOI21_X1 u0_u1_u6_U11 (.B1( u0_u1_u6_n107 ) , .B2( u0_u1_u6_n132 ) , .A( u0_u1_u6_n158 ) , .ZN( u0_u1_u6_n88 ) );
  AOI21_X1 u0_u1_u6_U12 (.B2( u0_u1_u6_n147 ) , .B1( u0_u1_u6_n148 ) , .ZN( u0_u1_u6_n149 ) , .A( u0_u1_u6_n158 ) );
  AOI21_X1 u0_u1_u6_U13 (.ZN( u0_u1_u6_n106 ) , .A( u0_u1_u6_n142 ) , .B2( u0_u1_u6_n159 ) , .B1( u0_u1_u6_n164 ) );
  INV_X1 u0_u1_u6_U14 (.A( u0_u1_u6_n155 ) , .ZN( u0_u1_u6_n161 ) );
  INV_X1 u0_u1_u6_U15 (.A( u0_u1_u6_n128 ) , .ZN( u0_u1_u6_n164 ) );
  NAND2_X1 u0_u1_u6_U16 (.ZN( u0_u1_u6_n110 ) , .A1( u0_u1_u6_n122 ) , .A2( u0_u1_u6_n129 ) );
  NAND2_X1 u0_u1_u6_U17 (.ZN( u0_u1_u6_n124 ) , .A2( u0_u1_u6_n146 ) , .A1( u0_u1_u6_n148 ) );
  INV_X1 u0_u1_u6_U18 (.A( u0_u1_u6_n132 ) , .ZN( u0_u1_u6_n171 ) );
  AND2_X1 u0_u1_u6_U19 (.A1( u0_u1_u6_n100 ) , .ZN( u0_u1_u6_n130 ) , .A2( u0_u1_u6_n147 ) );
  INV_X1 u0_u1_u6_U20 (.A( u0_u1_u6_n127 ) , .ZN( u0_u1_u6_n173 ) );
  INV_X1 u0_u1_u6_U21 (.A( u0_u1_u6_n121 ) , .ZN( u0_u1_u6_n167 ) );
  INV_X1 u0_u1_u6_U22 (.A( u0_u1_u6_n100 ) , .ZN( u0_u1_u6_n169 ) );
  INV_X1 u0_u1_u6_U23 (.A( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n170 ) );
  INV_X1 u0_u1_u6_U24 (.A( u0_u1_u6_n113 ) , .ZN( u0_u1_u6_n168 ) );
  AND2_X1 u0_u1_u6_U25 (.A1( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n119 ) , .ZN( u0_u1_u6_n133 ) );
  AND2_X1 u0_u1_u6_U26 (.A2( u0_u1_u6_n121 ) , .A1( u0_u1_u6_n122 ) , .ZN( u0_u1_u6_n131 ) );
  AND3_X1 u0_u1_u6_U27 (.ZN( u0_u1_u6_n120 ) , .A2( u0_u1_u6_n127 ) , .A1( u0_u1_u6_n132 ) , .A3( u0_u1_u6_n145 ) );
  INV_X1 u0_u1_u6_U28 (.A( u0_u1_u6_n146 ) , .ZN( u0_u1_u6_n163 ) );
  AOI222_X1 u0_u1_u6_U29 (.ZN( u0_u1_u6_n114 ) , .A1( u0_u1_u6_n118 ) , .A2( u0_u1_u6_n126 ) , .B2( u0_u1_u6_n151 ) , .C2( u0_u1_u6_n159 ) , .C1( u0_u1_u6_n168 ) , .B1( u0_u1_u6_n169 ) );
  INV_X1 u0_u1_u6_U3 (.A( u0_u1_u6_n110 ) , .ZN( u0_u1_u6_n166 ) );
  NOR2_X1 u0_u1_u6_U30 (.A1( u0_u1_u6_n162 ) , .A2( u0_u1_u6_n165 ) , .ZN( u0_u1_u6_n98 ) );
  AOI211_X1 u0_u1_u6_U31 (.B( u0_u1_u6_n134 ) , .A( u0_u1_u6_n135 ) , .C1( u0_u1_u6_n136 ) , .ZN( u0_u1_u6_n137 ) , .C2( u0_u1_u6_n151 ) );
  AOI21_X1 u0_u1_u6_U32 (.B1( u0_u1_u6_n131 ) , .ZN( u0_u1_u6_n135 ) , .A( u0_u1_u6_n144 ) , .B2( u0_u1_u6_n146 ) );
  NAND4_X1 u0_u1_u6_U33 (.A4( u0_u1_u6_n127 ) , .A3( u0_u1_u6_n128 ) , .A2( u0_u1_u6_n129 ) , .A1( u0_u1_u6_n130 ) , .ZN( u0_u1_u6_n136 ) );
  AOI21_X1 u0_u1_u6_U34 (.B2( u0_u1_u6_n132 ) , .B1( u0_u1_u6_n133 ) , .ZN( u0_u1_u6_n134 ) , .A( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U35 (.A1( u0_u1_u6_n144 ) , .ZN( u0_u1_u6_n151 ) , .A2( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U36 (.ZN( u0_u1_u6_n132 ) , .A1( u0_u1_u6_n91 ) , .A2( u0_u1_u6_n97 ) );
  AOI22_X1 u0_u1_u6_U37 (.B2( u0_u1_u6_n110 ) , .B1( u0_u1_u6_n111 ) , .A1( u0_u1_u6_n112 ) , .ZN( u0_u1_u6_n115 ) , .A2( u0_u1_u6_n161 ) );
  NAND4_X1 u0_u1_u6_U38 (.A3( u0_u1_u6_n109 ) , .ZN( u0_u1_u6_n112 ) , .A4( u0_u1_u6_n132 ) , .A2( u0_u1_u6_n147 ) , .A1( u0_u1_u6_n166 ) );
  NOR2_X1 u0_u1_u6_U39 (.ZN( u0_u1_u6_n109 ) , .A1( u0_u1_u6_n170 ) , .A2( u0_u1_u6_n173 ) );
  INV_X1 u0_u1_u6_U4 (.A( u0_u1_u6_n142 ) , .ZN( u0_u1_u6_n174 ) );
  NOR2_X1 u0_u1_u6_U40 (.A2( u0_u1_u6_n126 ) , .ZN( u0_u1_u6_n155 ) , .A1( u0_u1_u6_n160 ) );
  NAND2_X1 u0_u1_u6_U41 (.ZN( u0_u1_u6_n146 ) , .A2( u0_u1_u6_n94 ) , .A1( u0_u1_u6_n99 ) );
  AOI21_X1 u0_u1_u6_U42 (.A( u0_u1_u6_n144 ) , .B2( u0_u1_u6_n145 ) , .B1( u0_u1_u6_n146 ) , .ZN( u0_u1_u6_n150 ) );
  INV_X1 u0_u1_u6_U43 (.A( u0_u1_u6_n111 ) , .ZN( u0_u1_u6_n158 ) );
  NAND2_X1 u0_u1_u6_U44 (.ZN( u0_u1_u6_n127 ) , .A1( u0_u1_u6_n91 ) , .A2( u0_u1_u6_n92 ) );
  NAND2_X1 u0_u1_u6_U45 (.ZN( u0_u1_u6_n129 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n96 ) );
  INV_X1 u0_u1_u6_U46 (.A( u0_u1_u6_n144 ) , .ZN( u0_u1_u6_n159 ) );
  NAND2_X1 u0_u1_u6_U47 (.ZN( u0_u1_u6_n145 ) , .A2( u0_u1_u6_n97 ) , .A1( u0_u1_u6_n98 ) );
  NAND2_X1 u0_u1_u6_U48 (.ZN( u0_u1_u6_n148 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n94 ) );
  NAND2_X1 u0_u1_u6_U49 (.ZN( u0_u1_u6_n108 ) , .A2( u0_u1_u6_n139 ) , .A1( u0_u1_u6_n144 ) );
  NAND2_X1 u0_u1_u6_U5 (.A2( u0_u1_u6_n143 ) , .ZN( u0_u1_u6_n152 ) , .A1( u0_u1_u6_n166 ) );
  NAND2_X1 u0_u1_u6_U50 (.ZN( u0_u1_u6_n121 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n97 ) );
  NAND2_X1 u0_u1_u6_U51 (.ZN( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n95 ) );
  AND2_X1 u0_u1_u6_U52 (.ZN( u0_u1_u6_n118 ) , .A2( u0_u1_u6_n91 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U53 (.ZN( u0_u1_u6_n147 ) , .A2( u0_u1_u6_n98 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U54 (.ZN( u0_u1_u6_n128 ) , .A1( u0_u1_u6_n94 ) , .A2( u0_u1_u6_n96 ) );
  NAND2_X1 u0_u1_u6_U55 (.ZN( u0_u1_u6_n119 ) , .A2( u0_u1_u6_n95 ) , .A1( u0_u1_u6_n99 ) );
  NAND2_X1 u0_u1_u6_U56 (.ZN( u0_u1_u6_n123 ) , .A2( u0_u1_u6_n91 ) , .A1( u0_u1_u6_n96 ) );
  NAND2_X1 u0_u1_u6_U57 (.ZN( u0_u1_u6_n100 ) , .A2( u0_u1_u6_n92 ) , .A1( u0_u1_u6_n98 ) );
  NAND2_X1 u0_u1_u6_U58 (.ZN( u0_u1_u6_n122 ) , .A1( u0_u1_u6_n94 ) , .A2( u0_u1_u6_n97 ) );
  INV_X1 u0_u1_u6_U59 (.A( u0_u1_u6_n139 ) , .ZN( u0_u1_u6_n160 ) );
  AOI22_X1 u0_u1_u6_U6 (.B2( u0_u1_u6_n101 ) , .A1( u0_u1_u6_n102 ) , .ZN( u0_u1_u6_n103 ) , .B1( u0_u1_u6_n160 ) , .A2( u0_u1_u6_n161 ) );
  NAND2_X1 u0_u1_u6_U60 (.ZN( u0_u1_u6_n113 ) , .A1( u0_u1_u6_n96 ) , .A2( u0_u1_u6_n98 ) );
  NOR2_X1 u0_u1_u6_U61 (.A2( u0_u1_X_40 ) , .A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n126 ) );
  NOR2_X1 u0_u1_u6_U62 (.A2( u0_u1_X_39 ) , .A1( u0_u1_X_42 ) , .ZN( u0_u1_u6_n92 ) );
  NOR2_X1 u0_u1_u6_U63 (.A2( u0_u1_X_39 ) , .A1( u0_u1_u6_n156 ) , .ZN( u0_u1_u6_n97 ) );
  NOR2_X1 u0_u1_u6_U64 (.A2( u0_u1_X_38 ) , .A1( u0_u1_u6_n165 ) , .ZN( u0_u1_u6_n95 ) );
  NOR2_X1 u0_u1_u6_U65 (.A2( u0_u1_X_41 ) , .ZN( u0_u1_u6_n111 ) , .A1( u0_u1_u6_n157 ) );
  NOR2_X1 u0_u1_u6_U66 (.A2( u0_u1_X_37 ) , .A1( u0_u1_u6_n162 ) , .ZN( u0_u1_u6_n94 ) );
  NOR2_X1 u0_u1_u6_U67 (.A2( u0_u1_X_37 ) , .A1( u0_u1_X_38 ) , .ZN( u0_u1_u6_n91 ) );
  NAND2_X1 u0_u1_u6_U68 (.A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n144 ) , .A2( u0_u1_u6_n157 ) );
  NAND2_X1 u0_u1_u6_U69 (.A2( u0_u1_X_40 ) , .A1( u0_u1_X_41 ) , .ZN( u0_u1_u6_n139 ) );
  NOR2_X1 u0_u1_u6_U7 (.A1( u0_u1_u6_n118 ) , .ZN( u0_u1_u6_n143 ) , .A2( u0_u1_u6_n168 ) );
  AND2_X1 u0_u1_u6_U70 (.A1( u0_u1_X_39 ) , .A2( u0_u1_u6_n156 ) , .ZN( u0_u1_u6_n96 ) );
  AND2_X1 u0_u1_u6_U71 (.A1( u0_u1_X_39 ) , .A2( u0_u1_X_42 ) , .ZN( u0_u1_u6_n99 ) );
  INV_X1 u0_u1_u6_U72 (.A( u0_u1_X_40 ) , .ZN( u0_u1_u6_n157 ) );
  INV_X1 u0_u1_u6_U73 (.A( u0_u1_X_37 ) , .ZN( u0_u1_u6_n165 ) );
  INV_X1 u0_u1_u6_U74 (.A( u0_u1_X_38 ) , .ZN( u0_u1_u6_n162 ) );
  INV_X1 u0_u1_u6_U75 (.A( u0_u1_X_42 ) , .ZN( u0_u1_u6_n156 ) );
  NAND4_X1 u0_u1_u6_U76 (.ZN( u0_out1_12 ) , .A4( u0_u1_u6_n114 ) , .A3( u0_u1_u6_n115 ) , .A2( u0_u1_u6_n116 ) , .A1( u0_u1_u6_n117 ) );
  OAI22_X1 u0_u1_u6_U77 (.B2( u0_u1_u6_n111 ) , .ZN( u0_u1_u6_n116 ) , .B1( u0_u1_u6_n126 ) , .A2( u0_u1_u6_n164 ) , .A1( u0_u1_u6_n167 ) );
  OAI21_X1 u0_u1_u6_U78 (.A( u0_u1_u6_n108 ) , .ZN( u0_u1_u6_n117 ) , .B2( u0_u1_u6_n141 ) , .B1( u0_u1_u6_n163 ) );
  NAND4_X1 u0_u1_u6_U79 (.ZN( u0_out1_32 ) , .A4( u0_u1_u6_n103 ) , .A3( u0_u1_u6_n104 ) , .A2( u0_u1_u6_n105 ) , .A1( u0_u1_u6_n106 ) );
  OAI21_X1 u0_u1_u6_U8 (.A( u0_u1_u6_n159 ) , .B1( u0_u1_u6_n169 ) , .B2( u0_u1_u6_n173 ) , .ZN( u0_u1_u6_n90 ) );
  AOI22_X1 u0_u1_u6_U80 (.ZN( u0_u1_u6_n105 ) , .A2( u0_u1_u6_n108 ) , .A1( u0_u1_u6_n118 ) , .B2( u0_u1_u6_n126 ) , .B1( u0_u1_u6_n171 ) );
  AOI22_X1 u0_u1_u6_U81 (.ZN( u0_u1_u6_n104 ) , .A1( u0_u1_u6_n111 ) , .B1( u0_u1_u6_n124 ) , .B2( u0_u1_u6_n151 ) , .A2( u0_u1_u6_n93 ) );
  OAI211_X1 u0_u1_u6_U82 (.ZN( u0_out1_22 ) , .B( u0_u1_u6_n137 ) , .A( u0_u1_u6_n138 ) , .C2( u0_u1_u6_n139 ) , .C1( u0_u1_u6_n140 ) );
  AND4_X1 u0_u1_u6_U83 (.A3( u0_u1_u6_n119 ) , .A1( u0_u1_u6_n120 ) , .A4( u0_u1_u6_n129 ) , .ZN( u0_u1_u6_n140 ) , .A2( u0_u1_u6_n143 ) );
  AOI22_X1 u0_u1_u6_U84 (.B1( u0_u1_u6_n124 ) , .A2( u0_u1_u6_n125 ) , .A1( u0_u1_u6_n126 ) , .ZN( u0_u1_u6_n138 ) , .B2( u0_u1_u6_n161 ) );
  OAI211_X1 u0_u1_u6_U85 (.ZN( u0_out1_7 ) , .B( u0_u1_u6_n153 ) , .C2( u0_u1_u6_n154 ) , .C1( u0_u1_u6_n155 ) , .A( u0_u1_u6_n174 ) );
  NOR3_X1 u0_u1_u6_U86 (.A1( u0_u1_u6_n141 ) , .ZN( u0_u1_u6_n154 ) , .A3( u0_u1_u6_n164 ) , .A2( u0_u1_u6_n171 ) );
  AOI211_X1 u0_u1_u6_U87 (.B( u0_u1_u6_n149 ) , .A( u0_u1_u6_n150 ) , .C2( u0_u1_u6_n151 ) , .C1( u0_u1_u6_n152 ) , .ZN( u0_u1_u6_n153 ) );
  NAND3_X1 u0_u1_u6_U88 (.A2( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n125 ) , .A1( u0_u1_u6_n130 ) , .A3( u0_u1_u6_n131 ) );
  NAND3_X1 u0_u1_u6_U89 (.A3( u0_u1_u6_n133 ) , .ZN( u0_u1_u6_n141 ) , .A1( u0_u1_u6_n145 ) , .A2( u0_u1_u6_n148 ) );
  INV_X1 u0_u1_u6_U9 (.ZN( u0_u1_u6_n172 ) , .A( u0_u1_u6_n88 ) );
  NAND3_X1 u0_u1_u6_U90 (.ZN( u0_u1_u6_n101 ) , .A3( u0_u1_u6_n107 ) , .A2( u0_u1_u6_n121 ) , .A1( u0_u1_u6_n127 ) );
  NAND3_X1 u0_u1_u6_U91 (.ZN( u0_u1_u6_n102 ) , .A3( u0_u1_u6_n130 ) , .A2( u0_u1_u6_n145 ) , .A1( u0_u1_u6_n166 ) );
  NAND3_X1 u0_u1_u6_U92 (.A3( u0_u1_u6_n113 ) , .A1( u0_u1_u6_n119 ) , .A2( u0_u1_u6_n123 ) , .ZN( u0_u1_u6_n93 ) );
  NAND3_X1 u0_u1_u6_U93 (.ZN( u0_u1_u6_n142 ) , .A2( u0_u1_u6_n172 ) , .A3( u0_u1_u6_n89 ) , .A1( u0_u1_u6_n90 ) );
  XOR2_X1 u0_u2_U1 (.B( u0_K3_9 ) , .A( u0_R1_6 ) , .Z( u0_u2_X_9 ) );
  XOR2_X1 u0_u2_U16 (.B( u0_K3_3 ) , .A( u0_R1_2 ) , .Z( u0_u2_X_3 ) );
  XOR2_X1 u0_u2_U2 (.B( u0_K3_8 ) , .A( u0_R1_5 ) , .Z( u0_u2_X_8 ) );
  XOR2_X1 u0_u2_U20 (.B( u0_K3_36 ) , .A( u0_R1_25 ) , .Z( u0_u2_X_36 ) );
  XOR2_X1 u0_u2_U21 (.B( u0_K3_35 ) , .A( u0_R1_24 ) , .Z( u0_u2_X_35 ) );
  XOR2_X1 u0_u2_U22 (.B( u0_K3_34 ) , .A( u0_R1_23 ) , .Z( u0_u2_X_34 ) );
  XOR2_X1 u0_u2_U23 (.B( u0_K3_33 ) , .A( u0_R1_22 ) , .Z( u0_u2_X_33 ) );
  XOR2_X1 u0_u2_U24 (.B( u0_K3_32 ) , .A( u0_R1_21 ) , .Z( u0_u2_X_32 ) );
  XOR2_X1 u0_u2_U25 (.B( u0_K3_31 ) , .A( u0_R1_20 ) , .Z( u0_u2_X_31 ) );
  XOR2_X1 u0_u2_U27 (.B( u0_K3_2 ) , .A( u0_R1_1 ) , .Z( u0_u2_X_2 ) );
  XOR2_X1 u0_u2_U3 (.B( u0_K3_7 ) , .A( u0_R1_4 ) , .Z( u0_u2_X_7 ) );
  XOR2_X1 u0_u2_U33 (.B( u0_K3_24 ) , .A( u0_R1_17 ) , .Z( u0_u2_X_24 ) );
  XOR2_X1 u0_u2_U34 (.B( u0_K3_23 ) , .A( u0_R1_16 ) , .Z( u0_u2_X_23 ) );
  XOR2_X1 u0_u2_U35 (.B( u0_K3_22 ) , .A( u0_R1_15 ) , .Z( u0_u2_X_22 ) );
  XOR2_X1 u0_u2_U36 (.B( u0_K3_21 ) , .A( u0_R1_14 ) , .Z( u0_u2_X_21 ) );
  XOR2_X1 u0_u2_U37 (.B( u0_K3_20 ) , .A( u0_R1_13 ) , .Z( u0_u2_X_20 ) );
  XOR2_X1 u0_u2_U38 (.B( u0_K3_1 ) , .A( u0_R1_32 ) , .Z( u0_u2_X_1 ) );
  XOR2_X1 u0_u2_U39 (.B( u0_K3_19 ) , .A( u0_R1_12 ) , .Z( u0_u2_X_19 ) );
  XOR2_X1 u0_u2_U4 (.B( u0_K3_6 ) , .A( u0_R1_5 ) , .Z( u0_u2_X_6 ) );
  XOR2_X1 u0_u2_U40 (.B( u0_K3_18 ) , .A( u0_R1_13 ) , .Z( u0_u2_X_18 ) );
  XOR2_X1 u0_u2_U41 (.B( u0_K3_17 ) , .A( u0_R1_12 ) , .Z( u0_u2_X_17 ) );
  XOR2_X1 u0_u2_U42 (.B( u0_K3_16 ) , .A( u0_R1_11 ) , .Z( u0_u2_X_16 ) );
  XOR2_X1 u0_u2_U43 (.B( u0_K3_15 ) , .A( u0_R1_10 ) , .Z( u0_u2_X_15 ) );
  XOR2_X1 u0_u2_U44 (.B( u0_K3_14 ) , .A( u0_R1_9 ) , .Z( u0_u2_X_14 ) );
  XOR2_X1 u0_u2_U45 (.B( u0_K3_13 ) , .A( u0_R1_8 ) , .Z( u0_u2_X_13 ) );
  XOR2_X1 u0_u2_U46 (.B( u0_K3_12 ) , .A( u0_R1_9 ) , .Z( u0_u2_X_12 ) );
  XOR2_X1 u0_u2_U47 (.B( u0_K3_11 ) , .A( u0_R1_8 ) , .Z( u0_u2_X_11 ) );
  XOR2_X1 u0_u2_U48 (.B( u0_K3_10 ) , .A( u0_R1_7 ) , .Z( u0_u2_X_10 ) );
  XOR2_X1 u0_u2_U5 (.B( u0_K3_5 ) , .A( u0_R1_4 ) , .Z( u0_u2_X_5 ) );
  XOR2_X1 u0_u2_U6 (.B( u0_K3_4 ) , .A( u0_R1_3 ) , .Z( u0_u2_X_4 ) );
  AND3_X1 u0_u2_u0_U10 (.A2( u0_u2_u0_n112 ) , .ZN( u0_u2_u0_n127 ) , .A3( u0_u2_u0_n130 ) , .A1( u0_u2_u0_n148 ) );
  NAND2_X1 u0_u2_u0_U11 (.ZN( u0_u2_u0_n113 ) , .A1( u0_u2_u0_n139 ) , .A2( u0_u2_u0_n149 ) );
  AND2_X1 u0_u2_u0_U12 (.ZN( u0_u2_u0_n107 ) , .A1( u0_u2_u0_n130 ) , .A2( u0_u2_u0_n140 ) );
  AND2_X1 u0_u2_u0_U13 (.A2( u0_u2_u0_n129 ) , .A1( u0_u2_u0_n130 ) , .ZN( u0_u2_u0_n151 ) );
  AND2_X1 u0_u2_u0_U14 (.A1( u0_u2_u0_n108 ) , .A2( u0_u2_u0_n125 ) , .ZN( u0_u2_u0_n145 ) );
  INV_X1 u0_u2_u0_U15 (.A( u0_u2_u0_n143 ) , .ZN( u0_u2_u0_n173 ) );
  NOR2_X1 u0_u2_u0_U16 (.A2( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n147 ) , .A1( u0_u2_u0_n160 ) );
  INV_X1 u0_u2_u0_U17 (.ZN( u0_u2_u0_n172 ) , .A( u0_u2_u0_n88 ) );
  OAI222_X1 u0_u2_u0_U18 (.C1( u0_u2_u0_n108 ) , .A1( u0_u2_u0_n125 ) , .B2( u0_u2_u0_n128 ) , .B1( u0_u2_u0_n144 ) , .A2( u0_u2_u0_n158 ) , .C2( u0_u2_u0_n161 ) , .ZN( u0_u2_u0_n88 ) );
  NOR2_X1 u0_u2_u0_U19 (.A1( u0_u2_u0_n163 ) , .A2( u0_u2_u0_n164 ) , .ZN( u0_u2_u0_n95 ) );
  AOI21_X1 u0_u2_u0_U20 (.B1( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n132 ) , .A( u0_u2_u0_n165 ) , .B2( u0_u2_u0_n93 ) );
  INV_X1 u0_u2_u0_U21 (.A( u0_u2_u0_n142 ) , .ZN( u0_u2_u0_n165 ) );
  OAI221_X1 u0_u2_u0_U22 (.C1( u0_u2_u0_n121 ) , .ZN( u0_u2_u0_n122 ) , .B2( u0_u2_u0_n127 ) , .A( u0_u2_u0_n143 ) , .B1( u0_u2_u0_n144 ) , .C2( u0_u2_u0_n147 ) );
  OAI22_X1 u0_u2_u0_U23 (.B1( u0_u2_u0_n125 ) , .ZN( u0_u2_u0_n126 ) , .A1( u0_u2_u0_n138 ) , .A2( u0_u2_u0_n146 ) , .B2( u0_u2_u0_n147 ) );
  OAI22_X1 u0_u2_u0_U24 (.B1( u0_u2_u0_n131 ) , .A1( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n147 ) , .A2( u0_u2_u0_n90 ) , .ZN( u0_u2_u0_n91 ) );
  AND3_X1 u0_u2_u0_U25 (.A3( u0_u2_u0_n121 ) , .A2( u0_u2_u0_n125 ) , .A1( u0_u2_u0_n148 ) , .ZN( u0_u2_u0_n90 ) );
  INV_X1 u0_u2_u0_U26 (.A( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n161 ) );
  NOR2_X1 u0_u2_u0_U27 (.A1( u0_u2_u0_n120 ) , .ZN( u0_u2_u0_n143 ) , .A2( u0_u2_u0_n167 ) );
  OAI221_X1 u0_u2_u0_U28 (.C1( u0_u2_u0_n112 ) , .ZN( u0_u2_u0_n120 ) , .B1( u0_u2_u0_n138 ) , .B2( u0_u2_u0_n141 ) , .C2( u0_u2_u0_n147 ) , .A( u0_u2_u0_n172 ) );
  AOI211_X1 u0_u2_u0_U29 (.B( u0_u2_u0_n115 ) , .A( u0_u2_u0_n116 ) , .C2( u0_u2_u0_n117 ) , .C1( u0_u2_u0_n118 ) , .ZN( u0_u2_u0_n119 ) );
  INV_X1 u0_u2_u0_U3 (.A( u0_u2_u0_n113 ) , .ZN( u0_u2_u0_n166 ) );
  AOI22_X1 u0_u2_u0_U30 (.B2( u0_u2_u0_n109 ) , .A2( u0_u2_u0_n110 ) , .ZN( u0_u2_u0_n111 ) , .B1( u0_u2_u0_n118 ) , .A1( u0_u2_u0_n160 ) );
  INV_X1 u0_u2_u0_U31 (.A( u0_u2_u0_n118 ) , .ZN( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U32 (.ZN( u0_u2_u0_n104 ) , .B1( u0_u2_u0_n107 ) , .B2( u0_u2_u0_n141 ) , .A( u0_u2_u0_n144 ) );
  AOI21_X1 u0_u2_u0_U33 (.B1( u0_u2_u0_n127 ) , .B2( u0_u2_u0_n129 ) , .A( u0_u2_u0_n138 ) , .ZN( u0_u2_u0_n96 ) );
  AOI21_X1 u0_u2_u0_U34 (.ZN( u0_u2_u0_n116 ) , .B2( u0_u2_u0_n142 ) , .A( u0_u2_u0_n144 ) , .B1( u0_u2_u0_n166 ) );
  NAND2_X1 u0_u2_u0_U35 (.A1( u0_u2_u0_n100 ) , .A2( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n125 ) );
  NAND2_X1 u0_u2_u0_U36 (.A1( u0_u2_u0_n101 ) , .A2( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n150 ) );
  INV_X1 u0_u2_u0_U37 (.A( u0_u2_u0_n138 ) , .ZN( u0_u2_u0_n160 ) );
  NAND2_X1 u0_u2_u0_U38 (.A1( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n128 ) , .A2( u0_u2_u0_n95 ) );
  NAND2_X1 u0_u2_u0_U39 (.A1( u0_u2_u0_n100 ) , .ZN( u0_u2_u0_n129 ) , .A2( u0_u2_u0_n95 ) );
  AOI21_X1 u0_u2_u0_U4 (.B1( u0_u2_u0_n114 ) , .ZN( u0_u2_u0_n115 ) , .B2( u0_u2_u0_n129 ) , .A( u0_u2_u0_n161 ) );
  NAND2_X1 u0_u2_u0_U40 (.A2( u0_u2_u0_n100 ) , .ZN( u0_u2_u0_n131 ) , .A1( u0_u2_u0_n92 ) );
  NAND2_X1 u0_u2_u0_U41 (.A2( u0_u2_u0_n100 ) , .A1( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n139 ) );
  NAND2_X1 u0_u2_u0_U42 (.ZN( u0_u2_u0_n148 ) , .A1( u0_u2_u0_n93 ) , .A2( u0_u2_u0_n95 ) );
  NAND2_X1 u0_u2_u0_U43 (.A2( u0_u2_u0_n102 ) , .A1( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n149 ) );
  NAND2_X1 u0_u2_u0_U44 (.A2( u0_u2_u0_n102 ) , .ZN( u0_u2_u0_n114 ) , .A1( u0_u2_u0_n92 ) );
  NAND2_X1 u0_u2_u0_U45 (.A2( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n121 ) , .A1( u0_u2_u0_n93 ) );
  NAND2_X1 u0_u2_u0_U46 (.ZN( u0_u2_u0_n112 ) , .A2( u0_u2_u0_n92 ) , .A1( u0_u2_u0_n93 ) );
  OR3_X1 u0_u2_u0_U47 (.A3( u0_u2_u0_n152 ) , .A2( u0_u2_u0_n153 ) , .A1( u0_u2_u0_n154 ) , .ZN( u0_u2_u0_n155 ) );
  AOI21_X1 u0_u2_u0_U48 (.B2( u0_u2_u0_n150 ) , .B1( u0_u2_u0_n151 ) , .ZN( u0_u2_u0_n152 ) , .A( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U49 (.A( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n145 ) , .B1( u0_u2_u0_n146 ) , .ZN( u0_u2_u0_n154 ) );
  AOI21_X1 u0_u2_u0_U5 (.B2( u0_u2_u0_n131 ) , .ZN( u0_u2_u0_n134 ) , .B1( u0_u2_u0_n151 ) , .A( u0_u2_u0_n158 ) );
  AOI21_X1 u0_u2_u0_U50 (.A( u0_u2_u0_n147 ) , .B2( u0_u2_u0_n148 ) , .B1( u0_u2_u0_n149 ) , .ZN( u0_u2_u0_n153 ) );
  INV_X1 u0_u2_u0_U51 (.ZN( u0_u2_u0_n171 ) , .A( u0_u2_u0_n99 ) );
  OAI211_X1 u0_u2_u0_U52 (.C2( u0_u2_u0_n140 ) , .C1( u0_u2_u0_n161 ) , .A( u0_u2_u0_n169 ) , .B( u0_u2_u0_n98 ) , .ZN( u0_u2_u0_n99 ) );
  AOI211_X1 u0_u2_u0_U53 (.C1( u0_u2_u0_n118 ) , .A( u0_u2_u0_n123 ) , .B( u0_u2_u0_n96 ) , .C2( u0_u2_u0_n97 ) , .ZN( u0_u2_u0_n98 ) );
  INV_X1 u0_u2_u0_U54 (.ZN( u0_u2_u0_n169 ) , .A( u0_u2_u0_n91 ) );
  NOR2_X1 u0_u2_u0_U55 (.A2( u0_u2_X_6 ) , .ZN( u0_u2_u0_n100 ) , .A1( u0_u2_u0_n162 ) );
  NOR2_X1 u0_u2_u0_U56 (.A2( u0_u2_X_4 ) , .A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n118 ) );
  NOR2_X1 u0_u2_u0_U57 (.A2( u0_u2_X_2 ) , .ZN( u0_u2_u0_n103 ) , .A1( u0_u2_u0_n164 ) );
  NOR2_X1 u0_u2_u0_U58 (.A2( u0_u2_X_1 ) , .A1( u0_u2_X_2 ) , .ZN( u0_u2_u0_n92 ) );
  NOR2_X1 u0_u2_u0_U59 (.A2( u0_u2_X_1 ) , .ZN( u0_u2_u0_n101 ) , .A1( u0_u2_u0_n163 ) );
  NOR2_X1 u0_u2_u0_U6 (.A1( u0_u2_u0_n108 ) , .ZN( u0_u2_u0_n123 ) , .A2( u0_u2_u0_n158 ) );
  NAND2_X1 u0_u2_u0_U60 (.A2( u0_u2_X_4 ) , .A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n144 ) );
  NOR2_X1 u0_u2_u0_U61 (.A2( u0_u2_X_5 ) , .ZN( u0_u2_u0_n136 ) , .A1( u0_u2_u0_n159 ) );
  NAND2_X1 u0_u2_u0_U62 (.A1( u0_u2_X_5 ) , .ZN( u0_u2_u0_n138 ) , .A2( u0_u2_u0_n159 ) );
  AND2_X1 u0_u2_u0_U63 (.A2( u0_u2_X_3 ) , .A1( u0_u2_X_6 ) , .ZN( u0_u2_u0_n102 ) );
  AND2_X1 u0_u2_u0_U64 (.A1( u0_u2_X_6 ) , .A2( u0_u2_u0_n162 ) , .ZN( u0_u2_u0_n93 ) );
  INV_X1 u0_u2_u0_U65 (.A( u0_u2_X_4 ) , .ZN( u0_u2_u0_n159 ) );
  INV_X1 u0_u2_u0_U66 (.A( u0_u2_X_1 ) , .ZN( u0_u2_u0_n164 ) );
  INV_X1 u0_u2_u0_U67 (.A( u0_u2_X_2 ) , .ZN( u0_u2_u0_n163 ) );
  INV_X1 u0_u2_u0_U68 (.ZN( u0_u2_u0_n174 ) , .A( u0_u2_u0_n89 ) );
  AOI211_X1 u0_u2_u0_U69 (.B( u0_u2_u0_n104 ) , .A( u0_u2_u0_n105 ) , .ZN( u0_u2_u0_n106 ) , .C2( u0_u2_u0_n113 ) , .C1( u0_u2_u0_n160 ) );
  OAI21_X1 u0_u2_u0_U7 (.B1( u0_u2_u0_n150 ) , .B2( u0_u2_u0_n158 ) , .A( u0_u2_u0_n172 ) , .ZN( u0_u2_u0_n89 ) );
  INV_X1 u0_u2_u0_U70 (.A( u0_u2_u0_n126 ) , .ZN( u0_u2_u0_n168 ) );
  AOI211_X1 u0_u2_u0_U71 (.B( u0_u2_u0_n133 ) , .A( u0_u2_u0_n134 ) , .C2( u0_u2_u0_n135 ) , .C1( u0_u2_u0_n136 ) , .ZN( u0_u2_u0_n137 ) );
  OR4_X1 u0_u2_u0_U72 (.ZN( u0_out2_31 ) , .A4( u0_u2_u0_n155 ) , .A2( u0_u2_u0_n156 ) , .A1( u0_u2_u0_n157 ) , .A3( u0_u2_u0_n173 ) );
  AOI21_X1 u0_u2_u0_U73 (.A( u0_u2_u0_n138 ) , .B2( u0_u2_u0_n139 ) , .B1( u0_u2_u0_n140 ) , .ZN( u0_u2_u0_n157 ) );
  AOI21_X1 u0_u2_u0_U74 (.B2( u0_u2_u0_n141 ) , .B1( u0_u2_u0_n142 ) , .ZN( u0_u2_u0_n156 ) , .A( u0_u2_u0_n161 ) );
  OR4_X1 u0_u2_u0_U75 (.ZN( u0_out2_17 ) , .A4( u0_u2_u0_n122 ) , .A2( u0_u2_u0_n123 ) , .A1( u0_u2_u0_n124 ) , .A3( u0_u2_u0_n170 ) );
  AOI21_X1 u0_u2_u0_U76 (.B2( u0_u2_u0_n107 ) , .ZN( u0_u2_u0_n124 ) , .B1( u0_u2_u0_n128 ) , .A( u0_u2_u0_n161 ) );
  INV_X1 u0_u2_u0_U77 (.A( u0_u2_u0_n111 ) , .ZN( u0_u2_u0_n170 ) );
  AOI21_X1 u0_u2_u0_U78 (.B1( u0_u2_u0_n132 ) , .ZN( u0_u2_u0_n133 ) , .A( u0_u2_u0_n144 ) , .B2( u0_u2_u0_n166 ) );
  OAI22_X1 u0_u2_u0_U79 (.ZN( u0_u2_u0_n105 ) , .A2( u0_u2_u0_n132 ) , .B1( u0_u2_u0_n146 ) , .A1( u0_u2_u0_n147 ) , .B2( u0_u2_u0_n161 ) );
  AND2_X1 u0_u2_u0_U8 (.A1( u0_u2_u0_n114 ) , .A2( u0_u2_u0_n121 ) , .ZN( u0_u2_u0_n146 ) );
  NAND2_X1 u0_u2_u0_U80 (.ZN( u0_u2_u0_n110 ) , .A2( u0_u2_u0_n132 ) , .A1( u0_u2_u0_n145 ) );
  INV_X1 u0_u2_u0_U81 (.A( u0_u2_u0_n119 ) , .ZN( u0_u2_u0_n167 ) );
  NAND2_X1 u0_u2_u0_U82 (.A2( u0_u2_u0_n103 ) , .ZN( u0_u2_u0_n140 ) , .A1( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U83 (.A1( u0_u2_u0_n101 ) , .ZN( u0_u2_u0_n130 ) , .A2( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U84 (.ZN( u0_u2_u0_n108 ) , .A1( u0_u2_u0_n92 ) , .A2( u0_u2_u0_n94 ) );
  NAND2_X1 u0_u2_u0_U85 (.ZN( u0_u2_u0_n142 ) , .A1( u0_u2_u0_n94 ) , .A2( u0_u2_u0_n95 ) );
  INV_X1 u0_u2_u0_U86 (.A( u0_u2_X_3 ) , .ZN( u0_u2_u0_n162 ) );
  NOR2_X1 u0_u2_u0_U87 (.A2( u0_u2_X_3 ) , .A1( u0_u2_X_6 ) , .ZN( u0_u2_u0_n94 ) );
  NAND3_X1 u0_u2_u0_U88 (.ZN( u0_out2_23 ) , .A3( u0_u2_u0_n137 ) , .A1( u0_u2_u0_n168 ) , .A2( u0_u2_u0_n171 ) );
  NAND3_X1 u0_u2_u0_U89 (.A3( u0_u2_u0_n127 ) , .A2( u0_u2_u0_n128 ) , .ZN( u0_u2_u0_n135 ) , .A1( u0_u2_u0_n150 ) );
  AND2_X1 u0_u2_u0_U9 (.A1( u0_u2_u0_n131 ) , .ZN( u0_u2_u0_n141 ) , .A2( u0_u2_u0_n150 ) );
  NAND3_X1 u0_u2_u0_U90 (.ZN( u0_u2_u0_n117 ) , .A3( u0_u2_u0_n132 ) , .A2( u0_u2_u0_n139 ) , .A1( u0_u2_u0_n148 ) );
  NAND3_X1 u0_u2_u0_U91 (.ZN( u0_u2_u0_n109 ) , .A2( u0_u2_u0_n114 ) , .A3( u0_u2_u0_n140 ) , .A1( u0_u2_u0_n149 ) );
  NAND3_X1 u0_u2_u0_U92 (.ZN( u0_out2_9 ) , .A3( u0_u2_u0_n106 ) , .A2( u0_u2_u0_n171 ) , .A1( u0_u2_u0_n174 ) );
  NAND3_X1 u0_u2_u0_U93 (.A2( u0_u2_u0_n128 ) , .A1( u0_u2_u0_n132 ) , .A3( u0_u2_u0_n146 ) , .ZN( u0_u2_u0_n97 ) );
  NOR2_X1 u0_u2_u1_U10 (.A1( u0_u2_u1_n112 ) , .A2( u0_u2_u1_n116 ) , .ZN( u0_u2_u1_n118 ) );
  NAND3_X1 u0_u2_u1_U100 (.ZN( u0_u2_u1_n113 ) , .A1( u0_u2_u1_n120 ) , .A3( u0_u2_u1_n133 ) , .A2( u0_u2_u1_n155 ) );
  OAI21_X1 u0_u2_u1_U11 (.ZN( u0_u2_u1_n101 ) , .B1( u0_u2_u1_n141 ) , .A( u0_u2_u1_n146 ) , .B2( u0_u2_u1_n183 ) );
  AOI21_X1 u0_u2_u1_U12 (.B2( u0_u2_u1_n155 ) , .B1( u0_u2_u1_n156 ) , .ZN( u0_u2_u1_n157 ) , .A( u0_u2_u1_n174 ) );
  OR4_X1 u0_u2_u1_U13 (.A4( u0_u2_u1_n106 ) , .A3( u0_u2_u1_n107 ) , .ZN( u0_u2_u1_n108 ) , .A1( u0_u2_u1_n117 ) , .A2( u0_u2_u1_n184 ) );
  AOI21_X1 u0_u2_u1_U14 (.ZN( u0_u2_u1_n106 ) , .A( u0_u2_u1_n112 ) , .B1( u0_u2_u1_n154 ) , .B2( u0_u2_u1_n156 ) );
  INV_X1 u0_u2_u1_U15 (.A( u0_u2_u1_n101 ) , .ZN( u0_u2_u1_n184 ) );
  AOI21_X1 u0_u2_u1_U16 (.ZN( u0_u2_u1_n107 ) , .B1( u0_u2_u1_n134 ) , .B2( u0_u2_u1_n149 ) , .A( u0_u2_u1_n174 ) );
  NAND2_X1 u0_u2_u1_U17 (.ZN( u0_u2_u1_n140 ) , .A2( u0_u2_u1_n150 ) , .A1( u0_u2_u1_n155 ) );
  NAND2_X1 u0_u2_u1_U18 (.A1( u0_u2_u1_n131 ) , .ZN( u0_u2_u1_n147 ) , .A2( u0_u2_u1_n153 ) );
  INV_X1 u0_u2_u1_U19 (.A( u0_u2_u1_n139 ) , .ZN( u0_u2_u1_n174 ) );
  INV_X1 u0_u2_u1_U20 (.A( u0_u2_u1_n112 ) , .ZN( u0_u2_u1_n171 ) );
  NAND2_X1 u0_u2_u1_U21 (.ZN( u0_u2_u1_n141 ) , .A1( u0_u2_u1_n153 ) , .A2( u0_u2_u1_n156 ) );
  AND2_X1 u0_u2_u1_U22 (.A1( u0_u2_u1_n123 ) , .ZN( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n161 ) );
  NAND2_X1 u0_u2_u1_U23 (.A2( u0_u2_u1_n115 ) , .A1( u0_u2_u1_n116 ) , .ZN( u0_u2_u1_n148 ) );
  NAND2_X1 u0_u2_u1_U24 (.A2( u0_u2_u1_n133 ) , .A1( u0_u2_u1_n135 ) , .ZN( u0_u2_u1_n159 ) );
  NAND2_X1 u0_u2_u1_U25 (.A2( u0_u2_u1_n115 ) , .A1( u0_u2_u1_n120 ) , .ZN( u0_u2_u1_n132 ) );
  INV_X1 u0_u2_u1_U26 (.A( u0_u2_u1_n154 ) , .ZN( u0_u2_u1_n178 ) );
  INV_X1 u0_u2_u1_U27 (.A( u0_u2_u1_n151 ) , .ZN( u0_u2_u1_n183 ) );
  AND2_X1 u0_u2_u1_U28 (.A1( u0_u2_u1_n129 ) , .A2( u0_u2_u1_n133 ) , .ZN( u0_u2_u1_n149 ) );
  INV_X1 u0_u2_u1_U29 (.A( u0_u2_u1_n131 ) , .ZN( u0_u2_u1_n180 ) );
  INV_X1 u0_u2_u1_U3 (.A( u0_u2_u1_n159 ) , .ZN( u0_u2_u1_n182 ) );
  OAI221_X1 u0_u2_u1_U30 (.A( u0_u2_u1_n119 ) , .C2( u0_u2_u1_n129 ) , .ZN( u0_u2_u1_n138 ) , .B2( u0_u2_u1_n152 ) , .C1( u0_u2_u1_n174 ) , .B1( u0_u2_u1_n187 ) );
  INV_X1 u0_u2_u1_U31 (.A( u0_u2_u1_n148 ) , .ZN( u0_u2_u1_n187 ) );
  AOI211_X1 u0_u2_u1_U32 (.B( u0_u2_u1_n117 ) , .A( u0_u2_u1_n118 ) , .ZN( u0_u2_u1_n119 ) , .C2( u0_u2_u1_n146 ) , .C1( u0_u2_u1_n159 ) );
  NOR2_X1 u0_u2_u1_U33 (.A1( u0_u2_u1_n168 ) , .A2( u0_u2_u1_n176 ) , .ZN( u0_u2_u1_n98 ) );
  AOI211_X1 u0_u2_u1_U34 (.B( u0_u2_u1_n162 ) , .A( u0_u2_u1_n163 ) , .C2( u0_u2_u1_n164 ) , .ZN( u0_u2_u1_n165 ) , .C1( u0_u2_u1_n171 ) );
  AOI21_X1 u0_u2_u1_U35 (.A( u0_u2_u1_n160 ) , .B2( u0_u2_u1_n161 ) , .ZN( u0_u2_u1_n162 ) , .B1( u0_u2_u1_n182 ) );
  OR2_X1 u0_u2_u1_U36 (.A2( u0_u2_u1_n157 ) , .A1( u0_u2_u1_n158 ) , .ZN( u0_u2_u1_n163 ) );
  OAI21_X1 u0_u2_u1_U37 (.B2( u0_u2_u1_n123 ) , .ZN( u0_u2_u1_n145 ) , .B1( u0_u2_u1_n160 ) , .A( u0_u2_u1_n185 ) );
  INV_X1 u0_u2_u1_U38 (.A( u0_u2_u1_n122 ) , .ZN( u0_u2_u1_n185 ) );
  AOI21_X1 u0_u2_u1_U39 (.B2( u0_u2_u1_n120 ) , .B1( u0_u2_u1_n121 ) , .ZN( u0_u2_u1_n122 ) , .A( u0_u2_u1_n128 ) );
  AOI221_X1 u0_u2_u1_U4 (.A( u0_u2_u1_n138 ) , .C2( u0_u2_u1_n139 ) , .C1( u0_u2_u1_n140 ) , .B2( u0_u2_u1_n141 ) , .ZN( u0_u2_u1_n142 ) , .B1( u0_u2_u1_n175 ) );
  NAND2_X1 u0_u2_u1_U40 (.A1( u0_u2_u1_n128 ) , .ZN( u0_u2_u1_n146 ) , .A2( u0_u2_u1_n160 ) );
  NAND2_X1 u0_u2_u1_U41 (.A2( u0_u2_u1_n112 ) , .ZN( u0_u2_u1_n139 ) , .A1( u0_u2_u1_n152 ) );
  NAND2_X1 u0_u2_u1_U42 (.A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n156 ) , .A2( u0_u2_u1_n99 ) );
  AOI221_X1 u0_u2_u1_U43 (.B1( u0_u2_u1_n140 ) , .ZN( u0_u2_u1_n167 ) , .B2( u0_u2_u1_n172 ) , .C2( u0_u2_u1_n175 ) , .C1( u0_u2_u1_n178 ) , .A( u0_u2_u1_n188 ) );
  INV_X1 u0_u2_u1_U44 (.ZN( u0_u2_u1_n188 ) , .A( u0_u2_u1_n97 ) );
  AOI211_X1 u0_u2_u1_U45 (.A( u0_u2_u1_n118 ) , .C1( u0_u2_u1_n132 ) , .C2( u0_u2_u1_n139 ) , .B( u0_u2_u1_n96 ) , .ZN( u0_u2_u1_n97 ) );
  AOI21_X1 u0_u2_u1_U46 (.B2( u0_u2_u1_n121 ) , .B1( u0_u2_u1_n135 ) , .A( u0_u2_u1_n152 ) , .ZN( u0_u2_u1_n96 ) );
  NOR2_X1 u0_u2_u1_U47 (.ZN( u0_u2_u1_n117 ) , .A1( u0_u2_u1_n121 ) , .A2( u0_u2_u1_n160 ) );
  AOI21_X1 u0_u2_u1_U48 (.A( u0_u2_u1_n128 ) , .B2( u0_u2_u1_n129 ) , .ZN( u0_u2_u1_n130 ) , .B1( u0_u2_u1_n150 ) );
  NAND2_X1 u0_u2_u1_U49 (.ZN( u0_u2_u1_n112 ) , .A1( u0_u2_u1_n169 ) , .A2( u0_u2_u1_n170 ) );
  AOI211_X1 u0_u2_u1_U5 (.ZN( u0_u2_u1_n124 ) , .A( u0_u2_u1_n138 ) , .C2( u0_u2_u1_n139 ) , .B( u0_u2_u1_n145 ) , .C1( u0_u2_u1_n147 ) );
  NAND2_X1 u0_u2_u1_U50 (.ZN( u0_u2_u1_n129 ) , .A2( u0_u2_u1_n95 ) , .A1( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U51 (.A1( u0_u2_u1_n102 ) , .ZN( u0_u2_u1_n154 ) , .A2( u0_u2_u1_n99 ) );
  NAND2_X1 u0_u2_u1_U52 (.A2( u0_u2_u1_n100 ) , .ZN( u0_u2_u1_n135 ) , .A1( u0_u2_u1_n99 ) );
  AOI21_X1 u0_u2_u1_U53 (.A( u0_u2_u1_n152 ) , .B2( u0_u2_u1_n153 ) , .B1( u0_u2_u1_n154 ) , .ZN( u0_u2_u1_n158 ) );
  INV_X1 u0_u2_u1_U54 (.A( u0_u2_u1_n160 ) , .ZN( u0_u2_u1_n175 ) );
  NAND2_X1 u0_u2_u1_U55 (.A1( u0_u2_u1_n100 ) , .ZN( u0_u2_u1_n116 ) , .A2( u0_u2_u1_n95 ) );
  NAND2_X1 u0_u2_u1_U56 (.A1( u0_u2_u1_n102 ) , .ZN( u0_u2_u1_n131 ) , .A2( u0_u2_u1_n95 ) );
  NAND2_X1 u0_u2_u1_U57 (.A2( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n121 ) , .A1( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U58 (.A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n153 ) , .A2( u0_u2_u1_n98 ) );
  NAND2_X1 u0_u2_u1_U59 (.A2( u0_u2_u1_n104 ) , .A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n133 ) );
  AOI22_X1 u0_u2_u1_U6 (.B2( u0_u2_u1_n113 ) , .A2( u0_u2_u1_n114 ) , .ZN( u0_u2_u1_n125 ) , .A1( u0_u2_u1_n171 ) , .B1( u0_u2_u1_n173 ) );
  NAND2_X1 u0_u2_u1_U60 (.ZN( u0_u2_u1_n150 ) , .A2( u0_u2_u1_n98 ) , .A1( u0_u2_u1_n99 ) );
  NAND2_X1 u0_u2_u1_U61 (.A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n155 ) , .A2( u0_u2_u1_n95 ) );
  OAI21_X1 u0_u2_u1_U62 (.ZN( u0_u2_u1_n109 ) , .B1( u0_u2_u1_n129 ) , .B2( u0_u2_u1_n160 ) , .A( u0_u2_u1_n167 ) );
  NAND2_X1 u0_u2_u1_U63 (.A2( u0_u2_u1_n100 ) , .A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n120 ) );
  NAND2_X1 u0_u2_u1_U64 (.A1( u0_u2_u1_n102 ) , .A2( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n115 ) );
  NAND2_X1 u0_u2_u1_U65 (.A2( u0_u2_u1_n100 ) , .A1( u0_u2_u1_n104 ) , .ZN( u0_u2_u1_n151 ) );
  NAND2_X1 u0_u2_u1_U66 (.A2( u0_u2_u1_n103 ) , .A1( u0_u2_u1_n105 ) , .ZN( u0_u2_u1_n161 ) );
  INV_X1 u0_u2_u1_U67 (.A( u0_u2_u1_n152 ) , .ZN( u0_u2_u1_n173 ) );
  INV_X1 u0_u2_u1_U68 (.A( u0_u2_u1_n128 ) , .ZN( u0_u2_u1_n172 ) );
  NAND2_X1 u0_u2_u1_U69 (.A2( u0_u2_u1_n102 ) , .A1( u0_u2_u1_n103 ) , .ZN( u0_u2_u1_n123 ) );
  NAND2_X1 u0_u2_u1_U7 (.ZN( u0_u2_u1_n114 ) , .A1( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n156 ) );
  NOR2_X1 u0_u2_u1_U70 (.A2( u0_u2_X_7 ) , .A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n95 ) );
  NOR2_X1 u0_u2_u1_U71 (.A1( u0_u2_X_12 ) , .A2( u0_u2_X_9 ) , .ZN( u0_u2_u1_n100 ) );
  NOR2_X1 u0_u2_u1_U72 (.A2( u0_u2_X_8 ) , .A1( u0_u2_u1_n177 ) , .ZN( u0_u2_u1_n99 ) );
  NOR2_X1 u0_u2_u1_U73 (.A2( u0_u2_X_12 ) , .ZN( u0_u2_u1_n102 ) , .A1( u0_u2_u1_n176 ) );
  NOR2_X1 u0_u2_u1_U74 (.A2( u0_u2_X_9 ) , .ZN( u0_u2_u1_n105 ) , .A1( u0_u2_u1_n168 ) );
  NAND2_X1 u0_u2_u1_U75 (.A1( u0_u2_X_10 ) , .ZN( u0_u2_u1_n160 ) , .A2( u0_u2_u1_n169 ) );
  NAND2_X1 u0_u2_u1_U76 (.A2( u0_u2_X_10 ) , .A1( u0_u2_X_11 ) , .ZN( u0_u2_u1_n152 ) );
  NAND2_X1 u0_u2_u1_U77 (.A1( u0_u2_X_11 ) , .ZN( u0_u2_u1_n128 ) , .A2( u0_u2_u1_n170 ) );
  AND2_X1 u0_u2_u1_U78 (.A2( u0_u2_X_7 ) , .A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n104 ) );
  AND2_X1 u0_u2_u1_U79 (.A1( u0_u2_X_8 ) , .ZN( u0_u2_u1_n103 ) , .A2( u0_u2_u1_n177 ) );
  AOI22_X1 u0_u2_u1_U8 (.B2( u0_u2_u1_n136 ) , .A2( u0_u2_u1_n137 ) , .ZN( u0_u2_u1_n143 ) , .A1( u0_u2_u1_n171 ) , .B1( u0_u2_u1_n173 ) );
  INV_X1 u0_u2_u1_U80 (.A( u0_u2_X_10 ) , .ZN( u0_u2_u1_n170 ) );
  INV_X1 u0_u2_u1_U81 (.A( u0_u2_X_9 ) , .ZN( u0_u2_u1_n176 ) );
  INV_X1 u0_u2_u1_U82 (.A( u0_u2_X_11 ) , .ZN( u0_u2_u1_n169 ) );
  INV_X1 u0_u2_u1_U83 (.A( u0_u2_X_12 ) , .ZN( u0_u2_u1_n168 ) );
  INV_X1 u0_u2_u1_U84 (.A( u0_u2_X_7 ) , .ZN( u0_u2_u1_n177 ) );
  NAND4_X1 u0_u2_u1_U85 (.ZN( u0_out2_28 ) , .A4( u0_u2_u1_n124 ) , .A3( u0_u2_u1_n125 ) , .A2( u0_u2_u1_n126 ) , .A1( u0_u2_u1_n127 ) );
  OAI21_X1 u0_u2_u1_U86 (.ZN( u0_u2_u1_n127 ) , .B2( u0_u2_u1_n139 ) , .B1( u0_u2_u1_n175 ) , .A( u0_u2_u1_n183 ) );
  OAI21_X1 u0_u2_u1_U87 (.ZN( u0_u2_u1_n126 ) , .B2( u0_u2_u1_n140 ) , .A( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n178 ) );
  NAND4_X1 u0_u2_u1_U88 (.ZN( u0_out2_18 ) , .A4( u0_u2_u1_n165 ) , .A3( u0_u2_u1_n166 ) , .A1( u0_u2_u1_n167 ) , .A2( u0_u2_u1_n186 ) );
  AOI22_X1 u0_u2_u1_U89 (.B2( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n147 ) , .A2( u0_u2_u1_n148 ) , .ZN( u0_u2_u1_n166 ) , .A1( u0_u2_u1_n172 ) );
  INV_X1 u0_u2_u1_U9 (.A( u0_u2_u1_n147 ) , .ZN( u0_u2_u1_n181 ) );
  INV_X1 u0_u2_u1_U90 (.A( u0_u2_u1_n145 ) , .ZN( u0_u2_u1_n186 ) );
  NAND4_X1 u0_u2_u1_U91 (.ZN( u0_out2_2 ) , .A4( u0_u2_u1_n142 ) , .A3( u0_u2_u1_n143 ) , .A2( u0_u2_u1_n144 ) , .A1( u0_u2_u1_n179 ) );
  OAI21_X1 u0_u2_u1_U92 (.B2( u0_u2_u1_n132 ) , .ZN( u0_u2_u1_n144 ) , .A( u0_u2_u1_n146 ) , .B1( u0_u2_u1_n180 ) );
  INV_X1 u0_u2_u1_U93 (.A( u0_u2_u1_n130 ) , .ZN( u0_u2_u1_n179 ) );
  OR4_X1 u0_u2_u1_U94 (.ZN( u0_out2_13 ) , .A4( u0_u2_u1_n108 ) , .A3( u0_u2_u1_n109 ) , .A2( u0_u2_u1_n110 ) , .A1( u0_u2_u1_n111 ) );
  AOI21_X1 u0_u2_u1_U95 (.ZN( u0_u2_u1_n111 ) , .A( u0_u2_u1_n128 ) , .B2( u0_u2_u1_n131 ) , .B1( u0_u2_u1_n135 ) );
  AOI21_X1 u0_u2_u1_U96 (.ZN( u0_u2_u1_n110 ) , .A( u0_u2_u1_n116 ) , .B1( u0_u2_u1_n152 ) , .B2( u0_u2_u1_n160 ) );
  NAND3_X1 u0_u2_u1_U97 (.A3( u0_u2_u1_n149 ) , .A2( u0_u2_u1_n150 ) , .A1( u0_u2_u1_n151 ) , .ZN( u0_u2_u1_n164 ) );
  NAND3_X1 u0_u2_u1_U98 (.A3( u0_u2_u1_n134 ) , .A2( u0_u2_u1_n135 ) , .ZN( u0_u2_u1_n136 ) , .A1( u0_u2_u1_n151 ) );
  NAND3_X1 u0_u2_u1_U99 (.A1( u0_u2_u1_n133 ) , .ZN( u0_u2_u1_n137 ) , .A2( u0_u2_u1_n154 ) , .A3( u0_u2_u1_n181 ) );
  OAI22_X1 u0_u2_u2_U10 (.B1( u0_u2_u2_n151 ) , .A2( u0_u2_u2_n152 ) , .A1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n160 ) , .B2( u0_u2_u2_n168 ) );
  NAND3_X1 u0_u2_u2_U100 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n98 ) );
  NOR3_X1 u0_u2_u2_U11 (.A1( u0_u2_u2_n150 ) , .ZN( u0_u2_u2_n151 ) , .A3( u0_u2_u2_n175 ) , .A2( u0_u2_u2_n188 ) );
  AOI21_X1 u0_u2_u2_U12 (.B2( u0_u2_u2_n123 ) , .ZN( u0_u2_u2_n125 ) , .A( u0_u2_u2_n171 ) , .B1( u0_u2_u2_n184 ) );
  INV_X1 u0_u2_u2_U13 (.A( u0_u2_u2_n150 ) , .ZN( u0_u2_u2_n184 ) );
  AOI21_X1 u0_u2_u2_U14 (.ZN( u0_u2_u2_n144 ) , .B2( u0_u2_u2_n155 ) , .A( u0_u2_u2_n172 ) , .B1( u0_u2_u2_n185 ) );
  AOI21_X1 u0_u2_u2_U15 (.B2( u0_u2_u2_n143 ) , .ZN( u0_u2_u2_n145 ) , .B1( u0_u2_u2_n152 ) , .A( u0_u2_u2_n171 ) );
  INV_X1 u0_u2_u2_U16 (.A( u0_u2_u2_n156 ) , .ZN( u0_u2_u2_n171 ) );
  INV_X1 u0_u2_u2_U17 (.A( u0_u2_u2_n120 ) , .ZN( u0_u2_u2_n188 ) );
  NAND2_X1 u0_u2_u2_U18 (.A2( u0_u2_u2_n122 ) , .ZN( u0_u2_u2_n150 ) , .A1( u0_u2_u2_n152 ) );
  INV_X1 u0_u2_u2_U19 (.A( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n170 ) );
  INV_X1 u0_u2_u2_U20 (.A( u0_u2_u2_n137 ) , .ZN( u0_u2_u2_n173 ) );
  NAND2_X1 u0_u2_u2_U21 (.A1( u0_u2_u2_n132 ) , .A2( u0_u2_u2_n139 ) , .ZN( u0_u2_u2_n157 ) );
  INV_X1 u0_u2_u2_U22 (.A( u0_u2_u2_n113 ) , .ZN( u0_u2_u2_n178 ) );
  INV_X1 u0_u2_u2_U23 (.A( u0_u2_u2_n139 ) , .ZN( u0_u2_u2_n175 ) );
  INV_X1 u0_u2_u2_U24 (.A( u0_u2_u2_n155 ) , .ZN( u0_u2_u2_n181 ) );
  INV_X1 u0_u2_u2_U25 (.A( u0_u2_u2_n119 ) , .ZN( u0_u2_u2_n177 ) );
  INV_X1 u0_u2_u2_U26 (.A( u0_u2_u2_n116 ) , .ZN( u0_u2_u2_n180 ) );
  INV_X1 u0_u2_u2_U27 (.A( u0_u2_u2_n131 ) , .ZN( u0_u2_u2_n179 ) );
  INV_X1 u0_u2_u2_U28 (.A( u0_u2_u2_n154 ) , .ZN( u0_u2_u2_n176 ) );
  NAND2_X1 u0_u2_u2_U29 (.A2( u0_u2_u2_n116 ) , .A1( u0_u2_u2_n117 ) , .ZN( u0_u2_u2_n118 ) );
  NOR2_X1 u0_u2_u2_U3 (.ZN( u0_u2_u2_n121 ) , .A2( u0_u2_u2_n177 ) , .A1( u0_u2_u2_n180 ) );
  INV_X1 u0_u2_u2_U30 (.A( u0_u2_u2_n132 ) , .ZN( u0_u2_u2_n182 ) );
  INV_X1 u0_u2_u2_U31 (.A( u0_u2_u2_n158 ) , .ZN( u0_u2_u2_n183 ) );
  OAI21_X1 u0_u2_u2_U32 (.A( u0_u2_u2_n156 ) , .B1( u0_u2_u2_n157 ) , .ZN( u0_u2_u2_n158 ) , .B2( u0_u2_u2_n179 ) );
  NOR2_X1 u0_u2_u2_U33 (.ZN( u0_u2_u2_n156 ) , .A1( u0_u2_u2_n166 ) , .A2( u0_u2_u2_n169 ) );
  NOR2_X1 u0_u2_u2_U34 (.A2( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n137 ) , .A1( u0_u2_u2_n140 ) );
  NOR2_X1 u0_u2_u2_U35 (.A2( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n153 ) , .A1( u0_u2_u2_n156 ) );
  AOI211_X1 u0_u2_u2_U36 (.ZN( u0_u2_u2_n130 ) , .C1( u0_u2_u2_n138 ) , .C2( u0_u2_u2_n179 ) , .B( u0_u2_u2_n96 ) , .A( u0_u2_u2_n97 ) );
  OAI22_X1 u0_u2_u2_U37 (.B1( u0_u2_u2_n133 ) , .A2( u0_u2_u2_n137 ) , .A1( u0_u2_u2_n152 ) , .B2( u0_u2_u2_n168 ) , .ZN( u0_u2_u2_n97 ) );
  OAI221_X1 u0_u2_u2_U38 (.B1( u0_u2_u2_n113 ) , .C1( u0_u2_u2_n132 ) , .A( u0_u2_u2_n149 ) , .B2( u0_u2_u2_n171 ) , .C2( u0_u2_u2_n172 ) , .ZN( u0_u2_u2_n96 ) );
  OAI221_X1 u0_u2_u2_U39 (.A( u0_u2_u2_n115 ) , .C2( u0_u2_u2_n123 ) , .B2( u0_u2_u2_n143 ) , .B1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n163 ) , .C1( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U4 (.A( u0_u2_u2_n134 ) , .ZN( u0_u2_u2_n185 ) );
  OAI21_X1 u0_u2_u2_U40 (.A( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n115 ) , .B1( u0_u2_u2_n176 ) , .B2( u0_u2_u2_n178 ) );
  OAI221_X1 u0_u2_u2_U41 (.A( u0_u2_u2_n135 ) , .B2( u0_u2_u2_n136 ) , .B1( u0_u2_u2_n137 ) , .ZN( u0_u2_u2_n162 ) , .C2( u0_u2_u2_n167 ) , .C1( u0_u2_u2_n185 ) );
  AND3_X1 u0_u2_u2_U42 (.A3( u0_u2_u2_n131 ) , .A2( u0_u2_u2_n132 ) , .A1( u0_u2_u2_n133 ) , .ZN( u0_u2_u2_n136 ) );
  AOI22_X1 u0_u2_u2_U43 (.ZN( u0_u2_u2_n135 ) , .B1( u0_u2_u2_n140 ) , .A1( u0_u2_u2_n156 ) , .B2( u0_u2_u2_n180 ) , .A2( u0_u2_u2_n188 ) );
  AOI21_X1 u0_u2_u2_U44 (.ZN( u0_u2_u2_n149 ) , .B1( u0_u2_u2_n173 ) , .B2( u0_u2_u2_n188 ) , .A( u0_u2_u2_n95 ) );
  AND3_X1 u0_u2_u2_U45 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n156 ) , .ZN( u0_u2_u2_n95 ) );
  OAI21_X1 u0_u2_u2_U46 (.A( u0_u2_u2_n141 ) , .B2( u0_u2_u2_n142 ) , .ZN( u0_u2_u2_n146 ) , .B1( u0_u2_u2_n153 ) );
  OAI21_X1 u0_u2_u2_U47 (.A( u0_u2_u2_n140 ) , .ZN( u0_u2_u2_n141 ) , .B1( u0_u2_u2_n176 ) , .B2( u0_u2_u2_n177 ) );
  NOR3_X1 u0_u2_u2_U48 (.ZN( u0_u2_u2_n142 ) , .A3( u0_u2_u2_n175 ) , .A2( u0_u2_u2_n178 ) , .A1( u0_u2_u2_n181 ) );
  OAI21_X1 u0_u2_u2_U49 (.A( u0_u2_u2_n101 ) , .B2( u0_u2_u2_n121 ) , .B1( u0_u2_u2_n153 ) , .ZN( u0_u2_u2_n164 ) );
  NOR4_X1 u0_u2_u2_U5 (.A4( u0_u2_u2_n124 ) , .A3( u0_u2_u2_n125 ) , .A2( u0_u2_u2_n126 ) , .A1( u0_u2_u2_n127 ) , .ZN( u0_u2_u2_n128 ) );
  NAND2_X1 u0_u2_u2_U50 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n155 ) );
  NAND2_X1 u0_u2_u2_U51 (.A2( u0_u2_u2_n105 ) , .A1( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n143 ) );
  NAND2_X1 u0_u2_u2_U52 (.A1( u0_u2_u2_n104 ) , .A2( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n152 ) );
  NAND2_X1 u0_u2_u2_U53 (.A1( u0_u2_u2_n100 ) , .A2( u0_u2_u2_n105 ) , .ZN( u0_u2_u2_n132 ) );
  INV_X1 u0_u2_u2_U54 (.A( u0_u2_u2_n140 ) , .ZN( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U55 (.A( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n167 ) );
  INV_X1 u0_u2_u2_U56 (.ZN( u0_u2_u2_n187 ) , .A( u0_u2_u2_n99 ) );
  OAI21_X1 u0_u2_u2_U57 (.B1( u0_u2_u2_n137 ) , .B2( u0_u2_u2_n143 ) , .A( u0_u2_u2_n98 ) , .ZN( u0_u2_u2_n99 ) );
  NAND2_X1 u0_u2_u2_U58 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n113 ) );
  NAND2_X1 u0_u2_u2_U59 (.A1( u0_u2_u2_n106 ) , .A2( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n131 ) );
  AOI21_X1 u0_u2_u2_U6 (.B2( u0_u2_u2_n119 ) , .ZN( u0_u2_u2_n127 ) , .A( u0_u2_u2_n137 ) , .B1( u0_u2_u2_n155 ) );
  NAND2_X1 u0_u2_u2_U60 (.A1( u0_u2_u2_n103 ) , .A2( u0_u2_u2_n107 ) , .ZN( u0_u2_u2_n139 ) );
  NAND2_X1 u0_u2_u2_U61 (.A1( u0_u2_u2_n103 ) , .A2( u0_u2_u2_n105 ) , .ZN( u0_u2_u2_n133 ) );
  NAND2_X1 u0_u2_u2_U62 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n103 ) , .ZN( u0_u2_u2_n154 ) );
  NAND2_X1 u0_u2_u2_U63 (.A2( u0_u2_u2_n103 ) , .A1( u0_u2_u2_n104 ) , .ZN( u0_u2_u2_n119 ) );
  NAND2_X1 u0_u2_u2_U64 (.A2( u0_u2_u2_n107 ) , .A1( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n123 ) );
  NAND2_X1 u0_u2_u2_U65 (.A1( u0_u2_u2_n104 ) , .A2( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n122 ) );
  INV_X1 u0_u2_u2_U66 (.A( u0_u2_u2_n114 ) , .ZN( u0_u2_u2_n172 ) );
  NAND2_X1 u0_u2_u2_U67 (.A2( u0_u2_u2_n100 ) , .A1( u0_u2_u2_n102 ) , .ZN( u0_u2_u2_n116 ) );
  NAND2_X1 u0_u2_u2_U68 (.A1( u0_u2_u2_n102 ) , .A2( u0_u2_u2_n108 ) , .ZN( u0_u2_u2_n120 ) );
  NAND2_X1 u0_u2_u2_U69 (.A2( u0_u2_u2_n105 ) , .A1( u0_u2_u2_n106 ) , .ZN( u0_u2_u2_n117 ) );
  AOI21_X1 u0_u2_u2_U7 (.ZN( u0_u2_u2_n124 ) , .B1( u0_u2_u2_n131 ) , .B2( u0_u2_u2_n143 ) , .A( u0_u2_u2_n172 ) );
  NOR2_X1 u0_u2_u2_U70 (.A2( u0_u2_X_16 ) , .ZN( u0_u2_u2_n140 ) , .A1( u0_u2_u2_n166 ) );
  NOR2_X1 u0_u2_u2_U71 (.A2( u0_u2_X_13 ) , .A1( u0_u2_X_14 ) , .ZN( u0_u2_u2_n100 ) );
  NOR2_X1 u0_u2_u2_U72 (.A2( u0_u2_X_16 ) , .A1( u0_u2_X_17 ) , .ZN( u0_u2_u2_n138 ) );
  NOR2_X1 u0_u2_u2_U73 (.A2( u0_u2_X_15 ) , .A1( u0_u2_X_18 ) , .ZN( u0_u2_u2_n104 ) );
  NOR2_X1 u0_u2_u2_U74 (.A2( u0_u2_X_14 ) , .ZN( u0_u2_u2_n103 ) , .A1( u0_u2_u2_n174 ) );
  NOR2_X1 u0_u2_u2_U75 (.A2( u0_u2_X_15 ) , .ZN( u0_u2_u2_n102 ) , .A1( u0_u2_u2_n165 ) );
  NOR2_X1 u0_u2_u2_U76 (.A2( u0_u2_X_17 ) , .ZN( u0_u2_u2_n114 ) , .A1( u0_u2_u2_n169 ) );
  AND2_X1 u0_u2_u2_U77 (.A1( u0_u2_X_15 ) , .ZN( u0_u2_u2_n105 ) , .A2( u0_u2_u2_n165 ) );
  AND2_X1 u0_u2_u2_U78 (.A2( u0_u2_X_15 ) , .A1( u0_u2_X_18 ) , .ZN( u0_u2_u2_n107 ) );
  AND2_X1 u0_u2_u2_U79 (.A1( u0_u2_X_14 ) , .ZN( u0_u2_u2_n106 ) , .A2( u0_u2_u2_n174 ) );
  AOI21_X1 u0_u2_u2_U8 (.B2( u0_u2_u2_n120 ) , .B1( u0_u2_u2_n121 ) , .ZN( u0_u2_u2_n126 ) , .A( u0_u2_u2_n167 ) );
  AND2_X1 u0_u2_u2_U80 (.A1( u0_u2_X_13 ) , .A2( u0_u2_X_14 ) , .ZN( u0_u2_u2_n108 ) );
  INV_X1 u0_u2_u2_U81 (.A( u0_u2_X_16 ) , .ZN( u0_u2_u2_n169 ) );
  INV_X1 u0_u2_u2_U82 (.A( u0_u2_X_17 ) , .ZN( u0_u2_u2_n166 ) );
  INV_X1 u0_u2_u2_U83 (.A( u0_u2_X_13 ) , .ZN( u0_u2_u2_n174 ) );
  INV_X1 u0_u2_u2_U84 (.A( u0_u2_X_18 ) , .ZN( u0_u2_u2_n165 ) );
  NAND4_X1 u0_u2_u2_U85 (.ZN( u0_out2_24 ) , .A4( u0_u2_u2_n111 ) , .A3( u0_u2_u2_n112 ) , .A1( u0_u2_u2_n130 ) , .A2( u0_u2_u2_n187 ) );
  AOI21_X1 u0_u2_u2_U86 (.ZN( u0_u2_u2_n112 ) , .B2( u0_u2_u2_n156 ) , .A( u0_u2_u2_n164 ) , .B1( u0_u2_u2_n181 ) );
  AOI221_X1 u0_u2_u2_U87 (.A( u0_u2_u2_n109 ) , .B1( u0_u2_u2_n110 ) , .ZN( u0_u2_u2_n111 ) , .C1( u0_u2_u2_n134 ) , .C2( u0_u2_u2_n170 ) , .B2( u0_u2_u2_n173 ) );
  NAND4_X1 u0_u2_u2_U88 (.ZN( u0_out2_16 ) , .A4( u0_u2_u2_n128 ) , .A3( u0_u2_u2_n129 ) , .A1( u0_u2_u2_n130 ) , .A2( u0_u2_u2_n186 ) );
  AOI22_X1 u0_u2_u2_U89 (.A2( u0_u2_u2_n118 ) , .ZN( u0_u2_u2_n129 ) , .A1( u0_u2_u2_n140 ) , .B1( u0_u2_u2_n157 ) , .B2( u0_u2_u2_n170 ) );
  OAI22_X1 u0_u2_u2_U9 (.ZN( u0_u2_u2_n109 ) , .A2( u0_u2_u2_n113 ) , .B2( u0_u2_u2_n133 ) , .B1( u0_u2_u2_n167 ) , .A1( u0_u2_u2_n168 ) );
  INV_X1 u0_u2_u2_U90 (.A( u0_u2_u2_n163 ) , .ZN( u0_u2_u2_n186 ) );
  NAND4_X1 u0_u2_u2_U91 (.ZN( u0_out2_30 ) , .A4( u0_u2_u2_n147 ) , .A3( u0_u2_u2_n148 ) , .A2( u0_u2_u2_n149 ) , .A1( u0_u2_u2_n187 ) );
  NOR3_X1 u0_u2_u2_U92 (.A3( u0_u2_u2_n144 ) , .A2( u0_u2_u2_n145 ) , .A1( u0_u2_u2_n146 ) , .ZN( u0_u2_u2_n147 ) );
  AOI21_X1 u0_u2_u2_U93 (.B2( u0_u2_u2_n138 ) , .ZN( u0_u2_u2_n148 ) , .A( u0_u2_u2_n162 ) , .B1( u0_u2_u2_n182 ) );
  OR4_X1 u0_u2_u2_U94 (.ZN( u0_out2_6 ) , .A4( u0_u2_u2_n161 ) , .A3( u0_u2_u2_n162 ) , .A2( u0_u2_u2_n163 ) , .A1( u0_u2_u2_n164 ) );
  OR3_X1 u0_u2_u2_U95 (.A2( u0_u2_u2_n159 ) , .A1( u0_u2_u2_n160 ) , .ZN( u0_u2_u2_n161 ) , .A3( u0_u2_u2_n183 ) );
  AOI21_X1 u0_u2_u2_U96 (.B2( u0_u2_u2_n154 ) , .B1( u0_u2_u2_n155 ) , .ZN( u0_u2_u2_n159 ) , .A( u0_u2_u2_n167 ) );
  NAND3_X1 u0_u2_u2_U97 (.A2( u0_u2_u2_n117 ) , .A1( u0_u2_u2_n122 ) , .A3( u0_u2_u2_n123 ) , .ZN( u0_u2_u2_n134 ) );
  NAND3_X1 u0_u2_u2_U98 (.ZN( u0_u2_u2_n110 ) , .A2( u0_u2_u2_n131 ) , .A3( u0_u2_u2_n139 ) , .A1( u0_u2_u2_n154 ) );
  NAND3_X1 u0_u2_u2_U99 (.A2( u0_u2_u2_n100 ) , .ZN( u0_u2_u2_n101 ) , .A1( u0_u2_u2_n104 ) , .A3( u0_u2_u2_n114 ) );
  OAI22_X1 u0_u2_u3_U10 (.B1( u0_u2_u3_n113 ) , .A2( u0_u2_u3_n135 ) , .A1( u0_u2_u3_n150 ) , .B2( u0_u2_u3_n164 ) , .ZN( u0_u2_u3_n98 ) );
  OAI211_X1 u0_u2_u3_U11 (.B( u0_u2_u3_n106 ) , .ZN( u0_u2_u3_n119 ) , .C2( u0_u2_u3_n128 ) , .C1( u0_u2_u3_n167 ) , .A( u0_u2_u3_n181 ) );
  AOI221_X1 u0_u2_u3_U12 (.C1( u0_u2_u3_n105 ) , .ZN( u0_u2_u3_n106 ) , .A( u0_u2_u3_n131 ) , .B2( u0_u2_u3_n132 ) , .C2( u0_u2_u3_n133 ) , .B1( u0_u2_u3_n169 ) );
  INV_X1 u0_u2_u3_U13 (.ZN( u0_u2_u3_n181 ) , .A( u0_u2_u3_n98 ) );
  NAND2_X1 u0_u2_u3_U14 (.ZN( u0_u2_u3_n105 ) , .A2( u0_u2_u3_n130 ) , .A1( u0_u2_u3_n155 ) );
  AOI22_X1 u0_u2_u3_U15 (.B1( u0_u2_u3_n115 ) , .A2( u0_u2_u3_n116 ) , .ZN( u0_u2_u3_n123 ) , .B2( u0_u2_u3_n133 ) , .A1( u0_u2_u3_n169 ) );
  NAND2_X1 u0_u2_u3_U16 (.ZN( u0_u2_u3_n116 ) , .A2( u0_u2_u3_n151 ) , .A1( u0_u2_u3_n182 ) );
  NOR2_X1 u0_u2_u3_U17 (.ZN( u0_u2_u3_n126 ) , .A2( u0_u2_u3_n150 ) , .A1( u0_u2_u3_n164 ) );
  AOI21_X1 u0_u2_u3_U18 (.ZN( u0_u2_u3_n112 ) , .B2( u0_u2_u3_n146 ) , .B1( u0_u2_u3_n155 ) , .A( u0_u2_u3_n167 ) );
  NAND2_X1 u0_u2_u3_U19 (.A1( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n142 ) , .A2( u0_u2_u3_n164 ) );
  NAND2_X1 u0_u2_u3_U20 (.ZN( u0_u2_u3_n132 ) , .A2( u0_u2_u3_n152 ) , .A1( u0_u2_u3_n156 ) );
  AND2_X1 u0_u2_u3_U21 (.A2( u0_u2_u3_n113 ) , .A1( u0_u2_u3_n114 ) , .ZN( u0_u2_u3_n151 ) );
  INV_X1 u0_u2_u3_U22 (.A( u0_u2_u3_n133 ) , .ZN( u0_u2_u3_n165 ) );
  INV_X1 u0_u2_u3_U23 (.A( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n170 ) );
  NAND2_X1 u0_u2_u3_U24 (.A1( u0_u2_u3_n107 ) , .A2( u0_u2_u3_n108 ) , .ZN( u0_u2_u3_n140 ) );
  NAND2_X1 u0_u2_u3_U25 (.ZN( u0_u2_u3_n117 ) , .A1( u0_u2_u3_n124 ) , .A2( u0_u2_u3_n148 ) );
  NAND2_X1 u0_u2_u3_U26 (.ZN( u0_u2_u3_n143 ) , .A1( u0_u2_u3_n165 ) , .A2( u0_u2_u3_n167 ) );
  INV_X1 u0_u2_u3_U27 (.A( u0_u2_u3_n130 ) , .ZN( u0_u2_u3_n177 ) );
  INV_X1 u0_u2_u3_U28 (.A( u0_u2_u3_n128 ) , .ZN( u0_u2_u3_n176 ) );
  INV_X1 u0_u2_u3_U29 (.A( u0_u2_u3_n155 ) , .ZN( u0_u2_u3_n174 ) );
  INV_X1 u0_u2_u3_U3 (.A( u0_u2_u3_n129 ) , .ZN( u0_u2_u3_n183 ) );
  INV_X1 u0_u2_u3_U30 (.A( u0_u2_u3_n139 ) , .ZN( u0_u2_u3_n185 ) );
  NOR2_X1 u0_u2_u3_U31 (.ZN( u0_u2_u3_n135 ) , .A2( u0_u2_u3_n141 ) , .A1( u0_u2_u3_n169 ) );
  OAI222_X1 u0_u2_u3_U32 (.C2( u0_u2_u3_n107 ) , .A2( u0_u2_u3_n108 ) , .B1( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n138 ) , .B2( u0_u2_u3_n146 ) , .C1( u0_u2_u3_n154 ) , .A1( u0_u2_u3_n164 ) );
  NOR4_X1 u0_u2_u3_U33 (.A4( u0_u2_u3_n157 ) , .A3( u0_u2_u3_n158 ) , .A2( u0_u2_u3_n159 ) , .A1( u0_u2_u3_n160 ) , .ZN( u0_u2_u3_n161 ) );
  AOI21_X1 u0_u2_u3_U34 (.B2( u0_u2_u3_n152 ) , .B1( u0_u2_u3_n153 ) , .ZN( u0_u2_u3_n158 ) , .A( u0_u2_u3_n164 ) );
  AOI21_X1 u0_u2_u3_U35 (.A( u0_u2_u3_n154 ) , .B2( u0_u2_u3_n155 ) , .B1( u0_u2_u3_n156 ) , .ZN( u0_u2_u3_n157 ) );
  AOI21_X1 u0_u2_u3_U36 (.A( u0_u2_u3_n149 ) , .B2( u0_u2_u3_n150 ) , .B1( u0_u2_u3_n151 ) , .ZN( u0_u2_u3_n159 ) );
  AOI211_X1 u0_u2_u3_U37 (.ZN( u0_u2_u3_n109 ) , .A( u0_u2_u3_n119 ) , .C2( u0_u2_u3_n129 ) , .B( u0_u2_u3_n138 ) , .C1( u0_u2_u3_n141 ) );
  AOI211_X1 u0_u2_u3_U38 (.B( u0_u2_u3_n119 ) , .A( u0_u2_u3_n120 ) , .C2( u0_u2_u3_n121 ) , .ZN( u0_u2_u3_n122 ) , .C1( u0_u2_u3_n179 ) );
  INV_X1 u0_u2_u3_U39 (.A( u0_u2_u3_n156 ) , .ZN( u0_u2_u3_n179 ) );
  INV_X1 u0_u2_u3_U4 (.A( u0_u2_u3_n140 ) , .ZN( u0_u2_u3_n182 ) );
  OAI22_X1 u0_u2_u3_U40 (.B1( u0_u2_u3_n118 ) , .ZN( u0_u2_u3_n120 ) , .A1( u0_u2_u3_n135 ) , .B2( u0_u2_u3_n154 ) , .A2( u0_u2_u3_n178 ) );
  AND3_X1 u0_u2_u3_U41 (.ZN( u0_u2_u3_n118 ) , .A2( u0_u2_u3_n124 ) , .A1( u0_u2_u3_n144 ) , .A3( u0_u2_u3_n152 ) );
  INV_X1 u0_u2_u3_U42 (.A( u0_u2_u3_n121 ) , .ZN( u0_u2_u3_n164 ) );
  NAND2_X1 u0_u2_u3_U43 (.ZN( u0_u2_u3_n133 ) , .A1( u0_u2_u3_n154 ) , .A2( u0_u2_u3_n164 ) );
  OAI211_X1 u0_u2_u3_U44 (.B( u0_u2_u3_n127 ) , .ZN( u0_u2_u3_n139 ) , .C1( u0_u2_u3_n150 ) , .C2( u0_u2_u3_n154 ) , .A( u0_u2_u3_n184 ) );
  INV_X1 u0_u2_u3_U45 (.A( u0_u2_u3_n125 ) , .ZN( u0_u2_u3_n184 ) );
  AOI221_X1 u0_u2_u3_U46 (.A( u0_u2_u3_n126 ) , .ZN( u0_u2_u3_n127 ) , .C2( u0_u2_u3_n132 ) , .C1( u0_u2_u3_n169 ) , .B2( u0_u2_u3_n170 ) , .B1( u0_u2_u3_n174 ) );
  OAI22_X1 u0_u2_u3_U47 (.A1( u0_u2_u3_n124 ) , .ZN( u0_u2_u3_n125 ) , .B2( u0_u2_u3_n145 ) , .A2( u0_u2_u3_n165 ) , .B1( u0_u2_u3_n167 ) );
  NOR2_X1 u0_u2_u3_U48 (.A1( u0_u2_u3_n113 ) , .ZN( u0_u2_u3_n131 ) , .A2( u0_u2_u3_n154 ) );
  NAND2_X1 u0_u2_u3_U49 (.A1( u0_u2_u3_n103 ) , .ZN( u0_u2_u3_n150 ) , .A2( u0_u2_u3_n99 ) );
  INV_X1 u0_u2_u3_U5 (.A( u0_u2_u3_n117 ) , .ZN( u0_u2_u3_n178 ) );
  NAND2_X1 u0_u2_u3_U50 (.A2( u0_u2_u3_n102 ) , .ZN( u0_u2_u3_n155 ) , .A1( u0_u2_u3_n97 ) );
  INV_X1 u0_u2_u3_U51 (.A( u0_u2_u3_n141 ) , .ZN( u0_u2_u3_n167 ) );
  AOI21_X1 u0_u2_u3_U52 (.B2( u0_u2_u3_n114 ) , .B1( u0_u2_u3_n146 ) , .A( u0_u2_u3_n154 ) , .ZN( u0_u2_u3_n94 ) );
  AOI21_X1 u0_u2_u3_U53 (.ZN( u0_u2_u3_n110 ) , .B2( u0_u2_u3_n142 ) , .B1( u0_u2_u3_n186 ) , .A( u0_u2_u3_n95 ) );
  INV_X1 u0_u2_u3_U54 (.A( u0_u2_u3_n145 ) , .ZN( u0_u2_u3_n186 ) );
  AOI21_X1 u0_u2_u3_U55 (.B1( u0_u2_u3_n124 ) , .A( u0_u2_u3_n149 ) , .B2( u0_u2_u3_n155 ) , .ZN( u0_u2_u3_n95 ) );
  INV_X1 u0_u2_u3_U56 (.A( u0_u2_u3_n149 ) , .ZN( u0_u2_u3_n169 ) );
  NAND2_X1 u0_u2_u3_U57 (.ZN( u0_u2_u3_n124 ) , .A1( u0_u2_u3_n96 ) , .A2( u0_u2_u3_n97 ) );
  NAND2_X1 u0_u2_u3_U58 (.A2( u0_u2_u3_n100 ) , .ZN( u0_u2_u3_n146 ) , .A1( u0_u2_u3_n96 ) );
  NAND2_X1 u0_u2_u3_U59 (.A1( u0_u2_u3_n101 ) , .ZN( u0_u2_u3_n145 ) , .A2( u0_u2_u3_n99 ) );
  AOI221_X1 u0_u2_u3_U6 (.A( u0_u2_u3_n131 ) , .C2( u0_u2_u3_n132 ) , .C1( u0_u2_u3_n133 ) , .ZN( u0_u2_u3_n134 ) , .B1( u0_u2_u3_n143 ) , .B2( u0_u2_u3_n177 ) );
  NAND2_X1 u0_u2_u3_U60 (.A1( u0_u2_u3_n100 ) , .ZN( u0_u2_u3_n156 ) , .A2( u0_u2_u3_n99 ) );
  NAND2_X1 u0_u2_u3_U61 (.A2( u0_u2_u3_n101 ) , .A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n148 ) );
  NAND2_X1 u0_u2_u3_U62 (.A1( u0_u2_u3_n100 ) , .A2( u0_u2_u3_n102 ) , .ZN( u0_u2_u3_n128 ) );
  NAND2_X1 u0_u2_u3_U63 (.A2( u0_u2_u3_n101 ) , .A1( u0_u2_u3_n102 ) , .ZN( u0_u2_u3_n152 ) );
  NAND2_X1 u0_u2_u3_U64 (.A2( u0_u2_u3_n101 ) , .ZN( u0_u2_u3_n114 ) , .A1( u0_u2_u3_n96 ) );
  NAND2_X1 u0_u2_u3_U65 (.ZN( u0_u2_u3_n107 ) , .A1( u0_u2_u3_n97 ) , .A2( u0_u2_u3_n99 ) );
  NAND2_X1 u0_u2_u3_U66 (.A2( u0_u2_u3_n100 ) , .A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n113 ) );
  NAND2_X1 u0_u2_u3_U67 (.A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n153 ) , .A2( u0_u2_u3_n97 ) );
  NAND2_X1 u0_u2_u3_U68 (.A2( u0_u2_u3_n103 ) , .A1( u0_u2_u3_n104 ) , .ZN( u0_u2_u3_n130 ) );
  NAND2_X1 u0_u2_u3_U69 (.A2( u0_u2_u3_n103 ) , .ZN( u0_u2_u3_n144 ) , .A1( u0_u2_u3_n96 ) );
  OAI22_X1 u0_u2_u3_U7 (.B2( u0_u2_u3_n147 ) , .A2( u0_u2_u3_n148 ) , .ZN( u0_u2_u3_n160 ) , .B1( u0_u2_u3_n165 ) , .A1( u0_u2_u3_n168 ) );
  NAND2_X1 u0_u2_u3_U70 (.A1( u0_u2_u3_n102 ) , .A2( u0_u2_u3_n103 ) , .ZN( u0_u2_u3_n108 ) );
  NOR2_X1 u0_u2_u3_U71 (.A2( u0_u2_X_19 ) , .A1( u0_u2_X_20 ) , .ZN( u0_u2_u3_n99 ) );
  NOR2_X1 u0_u2_u3_U72 (.A2( u0_u2_X_21 ) , .A1( u0_u2_X_24 ) , .ZN( u0_u2_u3_n103 ) );
  NOR2_X1 u0_u2_u3_U73 (.A2( u0_u2_X_24 ) , .A1( u0_u2_u3_n171 ) , .ZN( u0_u2_u3_n97 ) );
  NOR2_X1 u0_u2_u3_U74 (.A2( u0_u2_X_23 ) , .ZN( u0_u2_u3_n141 ) , .A1( u0_u2_u3_n166 ) );
  NOR2_X1 u0_u2_u3_U75 (.A2( u0_u2_X_19 ) , .A1( u0_u2_u3_n172 ) , .ZN( u0_u2_u3_n96 ) );
  NAND2_X1 u0_u2_u3_U76 (.A1( u0_u2_X_22 ) , .A2( u0_u2_X_23 ) , .ZN( u0_u2_u3_n154 ) );
  NAND2_X1 u0_u2_u3_U77 (.A1( u0_u2_X_23 ) , .ZN( u0_u2_u3_n149 ) , .A2( u0_u2_u3_n166 ) );
  NOR2_X1 u0_u2_u3_U78 (.A2( u0_u2_X_22 ) , .A1( u0_u2_X_23 ) , .ZN( u0_u2_u3_n121 ) );
  AND2_X1 u0_u2_u3_U79 (.A1( u0_u2_X_24 ) , .ZN( u0_u2_u3_n101 ) , .A2( u0_u2_u3_n171 ) );
  AND3_X1 u0_u2_u3_U8 (.A3( u0_u2_u3_n144 ) , .A2( u0_u2_u3_n145 ) , .A1( u0_u2_u3_n146 ) , .ZN( u0_u2_u3_n147 ) );
  AND2_X1 u0_u2_u3_U80 (.A1( u0_u2_X_19 ) , .ZN( u0_u2_u3_n102 ) , .A2( u0_u2_u3_n172 ) );
  AND2_X1 u0_u2_u3_U81 (.A1( u0_u2_X_21 ) , .A2( u0_u2_X_24 ) , .ZN( u0_u2_u3_n100 ) );
  AND2_X1 u0_u2_u3_U82 (.A2( u0_u2_X_19 ) , .A1( u0_u2_X_20 ) , .ZN( u0_u2_u3_n104 ) );
  INV_X1 u0_u2_u3_U83 (.A( u0_u2_X_22 ) , .ZN( u0_u2_u3_n166 ) );
  INV_X1 u0_u2_u3_U84 (.A( u0_u2_X_21 ) , .ZN( u0_u2_u3_n171 ) );
  INV_X1 u0_u2_u3_U85 (.A( u0_u2_X_20 ) , .ZN( u0_u2_u3_n172 ) );
  OR4_X1 u0_u2_u3_U86 (.ZN( u0_out2_10 ) , .A4( u0_u2_u3_n136 ) , .A3( u0_u2_u3_n137 ) , .A1( u0_u2_u3_n138 ) , .A2( u0_u2_u3_n139 ) );
  OAI222_X1 u0_u2_u3_U87 (.C1( u0_u2_u3_n128 ) , .ZN( u0_u2_u3_n137 ) , .B1( u0_u2_u3_n148 ) , .A2( u0_u2_u3_n150 ) , .B2( u0_u2_u3_n154 ) , .C2( u0_u2_u3_n164 ) , .A1( u0_u2_u3_n167 ) );
  OAI221_X1 u0_u2_u3_U88 (.A( u0_u2_u3_n134 ) , .B2( u0_u2_u3_n135 ) , .ZN( u0_u2_u3_n136 ) , .C1( u0_u2_u3_n149 ) , .B1( u0_u2_u3_n151 ) , .C2( u0_u2_u3_n183 ) );
  NAND4_X1 u0_u2_u3_U89 (.ZN( u0_out2_26 ) , .A4( u0_u2_u3_n109 ) , .A3( u0_u2_u3_n110 ) , .A2( u0_u2_u3_n111 ) , .A1( u0_u2_u3_n173 ) );
  INV_X1 u0_u2_u3_U9 (.A( u0_u2_u3_n143 ) , .ZN( u0_u2_u3_n168 ) );
  INV_X1 u0_u2_u3_U90 (.ZN( u0_u2_u3_n173 ) , .A( u0_u2_u3_n94 ) );
  OAI21_X1 u0_u2_u3_U91 (.ZN( u0_u2_u3_n111 ) , .B2( u0_u2_u3_n117 ) , .A( u0_u2_u3_n133 ) , .B1( u0_u2_u3_n176 ) );
  NAND4_X1 u0_u2_u3_U92 (.ZN( u0_out2_20 ) , .A4( u0_u2_u3_n122 ) , .A3( u0_u2_u3_n123 ) , .A1( u0_u2_u3_n175 ) , .A2( u0_u2_u3_n180 ) );
  INV_X1 u0_u2_u3_U93 (.A( u0_u2_u3_n112 ) , .ZN( u0_u2_u3_n175 ) );
  INV_X1 u0_u2_u3_U94 (.A( u0_u2_u3_n126 ) , .ZN( u0_u2_u3_n180 ) );
  NAND4_X1 u0_u2_u3_U95 (.ZN( u0_out2_1 ) , .A4( u0_u2_u3_n161 ) , .A3( u0_u2_u3_n162 ) , .A2( u0_u2_u3_n163 ) , .A1( u0_u2_u3_n185 ) );
  NAND2_X1 u0_u2_u3_U96 (.ZN( u0_u2_u3_n163 ) , .A2( u0_u2_u3_n170 ) , .A1( u0_u2_u3_n176 ) );
  AOI22_X1 u0_u2_u3_U97 (.B2( u0_u2_u3_n140 ) , .B1( u0_u2_u3_n141 ) , .A2( u0_u2_u3_n142 ) , .ZN( u0_u2_u3_n162 ) , .A1( u0_u2_u3_n177 ) );
  NAND3_X1 u0_u2_u3_U98 (.A1( u0_u2_u3_n114 ) , .ZN( u0_u2_u3_n115 ) , .A2( u0_u2_u3_n145 ) , .A3( u0_u2_u3_n153 ) );
  NAND3_X1 u0_u2_u3_U99 (.ZN( u0_u2_u3_n129 ) , .A2( u0_u2_u3_n144 ) , .A1( u0_u2_u3_n153 ) , .A3( u0_u2_u3_n182 ) );
  INV_X1 u0_u2_u5_U10 (.A( u0_u2_u5_n121 ) , .ZN( u0_u2_u5_n177 ) );
  AOI222_X1 u0_u2_u5_U100 (.ZN( u0_u2_u5_n113 ) , .A1( u0_u2_u5_n131 ) , .C1( u0_u2_u5_n148 ) , .B2( u0_u2_u5_n174 ) , .C2( u0_u2_u5_n178 ) , .A2( u0_u2_u5_n179 ) , .B1( u0_u2_u5_n99 ) );
  NAND4_X1 u0_u2_u5_U101 (.ZN( u0_out2_29 ) , .A4( u0_u2_u5_n129 ) , .A3( u0_u2_u5_n130 ) , .A2( u0_u2_u5_n168 ) , .A1( u0_u2_u5_n196 ) );
  AOI221_X1 u0_u2_u5_U102 (.A( u0_u2_u5_n128 ) , .ZN( u0_u2_u5_n129 ) , .C2( u0_u2_u5_n132 ) , .B2( u0_u2_u5_n159 ) , .B1( u0_u2_u5_n176 ) , .C1( u0_u2_u5_n184 ) );
  AOI222_X1 u0_u2_u5_U103 (.ZN( u0_u2_u5_n130 ) , .A2( u0_u2_u5_n146 ) , .B1( u0_u2_u5_n147 ) , .C2( u0_u2_u5_n175 ) , .B2( u0_u2_u5_n179 ) , .A1( u0_u2_u5_n188 ) , .C1( u0_u2_u5_n194 ) );
  NAND3_X1 u0_u2_u5_U104 (.A2( u0_u2_u5_n154 ) , .A3( u0_u2_u5_n158 ) , .A1( u0_u2_u5_n161 ) , .ZN( u0_u2_u5_n99 ) );
  NOR2_X1 u0_u2_u5_U11 (.ZN( u0_u2_u5_n160 ) , .A2( u0_u2_u5_n173 ) , .A1( u0_u2_u5_n177 ) );
  INV_X1 u0_u2_u5_U12 (.A( u0_u2_u5_n150 ) , .ZN( u0_u2_u5_n174 ) );
  AOI21_X1 u0_u2_u5_U13 (.A( u0_u2_u5_n160 ) , .B2( u0_u2_u5_n161 ) , .ZN( u0_u2_u5_n162 ) , .B1( u0_u2_u5_n192 ) );
  INV_X1 u0_u2_u5_U14 (.A( u0_u2_u5_n159 ) , .ZN( u0_u2_u5_n192 ) );
  AOI21_X1 u0_u2_u5_U15 (.A( u0_u2_u5_n156 ) , .B2( u0_u2_u5_n157 ) , .B1( u0_u2_u5_n158 ) , .ZN( u0_u2_u5_n163 ) );
  AOI21_X1 u0_u2_u5_U16 (.B2( u0_u2_u5_n139 ) , .B1( u0_u2_u5_n140 ) , .ZN( u0_u2_u5_n141 ) , .A( u0_u2_u5_n150 ) );
  OAI21_X1 u0_u2_u5_U17 (.A( u0_u2_u5_n133 ) , .B2( u0_u2_u5_n134 ) , .B1( u0_u2_u5_n135 ) , .ZN( u0_u2_u5_n142 ) );
  OAI21_X1 u0_u2_u5_U18 (.ZN( u0_u2_u5_n133 ) , .B2( u0_u2_u5_n147 ) , .A( u0_u2_u5_n173 ) , .B1( u0_u2_u5_n188 ) );
  NAND2_X1 u0_u2_u5_U19 (.A2( u0_u2_u5_n119 ) , .A1( u0_u2_u5_n123 ) , .ZN( u0_u2_u5_n137 ) );
  INV_X1 u0_u2_u5_U20 (.A( u0_u2_u5_n155 ) , .ZN( u0_u2_u5_n194 ) );
  NAND2_X1 u0_u2_u5_U21 (.A1( u0_u2_u5_n121 ) , .ZN( u0_u2_u5_n132 ) , .A2( u0_u2_u5_n172 ) );
  NAND2_X1 u0_u2_u5_U22 (.A2( u0_u2_u5_n122 ) , .ZN( u0_u2_u5_n136 ) , .A1( u0_u2_u5_n154 ) );
  NAND2_X1 u0_u2_u5_U23 (.A2( u0_u2_u5_n119 ) , .A1( u0_u2_u5_n120 ) , .ZN( u0_u2_u5_n159 ) );
  INV_X1 u0_u2_u5_U24 (.A( u0_u2_u5_n156 ) , .ZN( u0_u2_u5_n175 ) );
  INV_X1 u0_u2_u5_U25 (.A( u0_u2_u5_n158 ) , .ZN( u0_u2_u5_n188 ) );
  INV_X1 u0_u2_u5_U26 (.A( u0_u2_u5_n152 ) , .ZN( u0_u2_u5_n179 ) );
  INV_X1 u0_u2_u5_U27 (.A( u0_u2_u5_n140 ) , .ZN( u0_u2_u5_n182 ) );
  INV_X1 u0_u2_u5_U28 (.A( u0_u2_u5_n151 ) , .ZN( u0_u2_u5_n183 ) );
  INV_X1 u0_u2_u5_U29 (.A( u0_u2_u5_n123 ) , .ZN( u0_u2_u5_n185 ) );
  NOR2_X1 u0_u2_u5_U3 (.ZN( u0_u2_u5_n134 ) , .A1( u0_u2_u5_n183 ) , .A2( u0_u2_u5_n190 ) );
  INV_X1 u0_u2_u5_U30 (.A( u0_u2_u5_n161 ) , .ZN( u0_u2_u5_n184 ) );
  INV_X1 u0_u2_u5_U31 (.A( u0_u2_u5_n139 ) , .ZN( u0_u2_u5_n189 ) );
  INV_X1 u0_u2_u5_U32 (.A( u0_u2_u5_n157 ) , .ZN( u0_u2_u5_n190 ) );
  INV_X1 u0_u2_u5_U33 (.A( u0_u2_u5_n120 ) , .ZN( u0_u2_u5_n193 ) );
  NAND2_X1 u0_u2_u5_U34 (.ZN( u0_u2_u5_n111 ) , .A1( u0_u2_u5_n140 ) , .A2( u0_u2_u5_n155 ) );
  INV_X1 u0_u2_u5_U35 (.A( u0_u2_u5_n117 ) , .ZN( u0_u2_u5_n196 ) );
  OAI221_X1 u0_u2_u5_U36 (.A( u0_u2_u5_n116 ) , .ZN( u0_u2_u5_n117 ) , .B2( u0_u2_u5_n119 ) , .C1( u0_u2_u5_n153 ) , .C2( u0_u2_u5_n158 ) , .B1( u0_u2_u5_n172 ) );
  AOI222_X1 u0_u2_u5_U37 (.ZN( u0_u2_u5_n116 ) , .B2( u0_u2_u5_n145 ) , .C1( u0_u2_u5_n148 ) , .A2( u0_u2_u5_n174 ) , .C2( u0_u2_u5_n177 ) , .B1( u0_u2_u5_n187 ) , .A1( u0_u2_u5_n193 ) );
  INV_X1 u0_u2_u5_U38 (.A( u0_u2_u5_n115 ) , .ZN( u0_u2_u5_n187 ) );
  NOR2_X1 u0_u2_u5_U39 (.ZN( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n170 ) , .A2( u0_u2_u5_n180 ) );
  INV_X1 u0_u2_u5_U4 (.A( u0_u2_u5_n138 ) , .ZN( u0_u2_u5_n191 ) );
  AOI22_X1 u0_u2_u5_U40 (.B2( u0_u2_u5_n131 ) , .A2( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n169 ) , .B1( u0_u2_u5_n174 ) , .A1( u0_u2_u5_n185 ) );
  NOR2_X1 u0_u2_u5_U41 (.A1( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n150 ) , .A2( u0_u2_u5_n173 ) );
  AOI21_X1 u0_u2_u5_U42 (.A( u0_u2_u5_n118 ) , .B2( u0_u2_u5_n145 ) , .ZN( u0_u2_u5_n168 ) , .B1( u0_u2_u5_n186 ) );
  INV_X1 u0_u2_u5_U43 (.A( u0_u2_u5_n122 ) , .ZN( u0_u2_u5_n186 ) );
  NOR2_X1 u0_u2_u5_U44 (.A1( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n152 ) , .A2( u0_u2_u5_n176 ) );
  NOR2_X1 u0_u2_u5_U45 (.A1( u0_u2_u5_n115 ) , .ZN( u0_u2_u5_n118 ) , .A2( u0_u2_u5_n153 ) );
  NOR2_X1 u0_u2_u5_U46 (.A2( u0_u2_u5_n145 ) , .ZN( u0_u2_u5_n156 ) , .A1( u0_u2_u5_n174 ) );
  NOR2_X1 u0_u2_u5_U47 (.ZN( u0_u2_u5_n121 ) , .A2( u0_u2_u5_n145 ) , .A1( u0_u2_u5_n176 ) );
  AOI22_X1 u0_u2_u5_U48 (.ZN( u0_u2_u5_n114 ) , .A2( u0_u2_u5_n137 ) , .A1( u0_u2_u5_n145 ) , .B2( u0_u2_u5_n175 ) , .B1( u0_u2_u5_n193 ) );
  AOI21_X1 u0_u2_u5_U49 (.A( u0_u2_u5_n153 ) , .B2( u0_u2_u5_n154 ) , .B1( u0_u2_u5_n155 ) , .ZN( u0_u2_u5_n164 ) );
  OAI21_X1 u0_u2_u5_U5 (.B2( u0_u2_u5_n136 ) , .B1( u0_u2_u5_n137 ) , .ZN( u0_u2_u5_n138 ) , .A( u0_u2_u5_n177 ) );
  AOI21_X1 u0_u2_u5_U50 (.ZN( u0_u2_u5_n110 ) , .B1( u0_u2_u5_n122 ) , .B2( u0_u2_u5_n139 ) , .A( u0_u2_u5_n153 ) );
  INV_X1 u0_u2_u5_U51 (.A( u0_u2_u5_n153 ) , .ZN( u0_u2_u5_n176 ) );
  INV_X1 u0_u2_u5_U52 (.A( u0_u2_u5_n126 ) , .ZN( u0_u2_u5_n173 ) );
  AND2_X1 u0_u2_u5_U53 (.A2( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n107 ) , .ZN( u0_u2_u5_n147 ) );
  AND2_X1 u0_u2_u5_U54 (.A2( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n108 ) , .ZN( u0_u2_u5_n148 ) );
  NAND2_X1 u0_u2_u5_U55 (.A1( u0_u2_u5_n105 ) , .A2( u0_u2_u5_n106 ) , .ZN( u0_u2_u5_n158 ) );
  NAND2_X1 u0_u2_u5_U56 (.A2( u0_u2_u5_n108 ) , .A1( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n139 ) );
  NAND2_X1 u0_u2_u5_U57 (.A1( u0_u2_u5_n106 ) , .A2( u0_u2_u5_n108 ) , .ZN( u0_u2_u5_n119 ) );
  OAI211_X1 u0_u2_u5_U58 (.B( u0_u2_u5_n124 ) , .A( u0_u2_u5_n125 ) , .C2( u0_u2_u5_n126 ) , .C1( u0_u2_u5_n127 ) , .ZN( u0_u2_u5_n128 ) );
  NOR3_X1 u0_u2_u5_U59 (.ZN( u0_u2_u5_n127 ) , .A1( u0_u2_u5_n136 ) , .A3( u0_u2_u5_n148 ) , .A2( u0_u2_u5_n182 ) );
  INV_X1 u0_u2_u5_U6 (.A( u0_u2_u5_n135 ) , .ZN( u0_u2_u5_n178 ) );
  OAI21_X1 u0_u2_u5_U60 (.ZN( u0_u2_u5_n124 ) , .A( u0_u2_u5_n177 ) , .B2( u0_u2_u5_n183 ) , .B1( u0_u2_u5_n189 ) );
  OAI21_X1 u0_u2_u5_U61 (.ZN( u0_u2_u5_n125 ) , .A( u0_u2_u5_n174 ) , .B2( u0_u2_u5_n185 ) , .B1( u0_u2_u5_n190 ) );
  NAND2_X1 u0_u2_u5_U62 (.A2( u0_u2_u5_n103 ) , .A1( u0_u2_u5_n105 ) , .ZN( u0_u2_u5_n140 ) );
  NAND2_X1 u0_u2_u5_U63 (.A2( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n105 ) , .ZN( u0_u2_u5_n155 ) );
  NAND2_X1 u0_u2_u5_U64 (.A2( u0_u2_u5_n106 ) , .A1( u0_u2_u5_n107 ) , .ZN( u0_u2_u5_n122 ) );
  NAND2_X1 u0_u2_u5_U65 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n106 ) , .ZN( u0_u2_u5_n115 ) );
  NAND2_X1 u0_u2_u5_U66 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n103 ) , .ZN( u0_u2_u5_n161 ) );
  NAND2_X1 u0_u2_u5_U67 (.A1( u0_u2_u5_n105 ) , .A2( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n154 ) );
  INV_X1 u0_u2_u5_U68 (.A( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n172 ) );
  NAND2_X1 u0_u2_u5_U69 (.A1( u0_u2_u5_n103 ) , .A2( u0_u2_u5_n108 ) , .ZN( u0_u2_u5_n123 ) );
  OAI22_X1 u0_u2_u5_U7 (.B2( u0_u2_u5_n149 ) , .B1( u0_u2_u5_n150 ) , .A2( u0_u2_u5_n151 ) , .A1( u0_u2_u5_n152 ) , .ZN( u0_u2_u5_n165 ) );
  NAND2_X1 u0_u2_u5_U70 (.A2( u0_u2_u5_n103 ) , .A1( u0_u2_u5_n107 ) , .ZN( u0_u2_u5_n151 ) );
  NAND2_X1 u0_u2_u5_U71 (.A2( u0_u2_u5_n107 ) , .A1( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n120 ) );
  NAND2_X1 u0_u2_u5_U72 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n109 ) , .ZN( u0_u2_u5_n157 ) );
  AND2_X1 u0_u2_u5_U73 (.A2( u0_u2_u5_n100 ) , .A1( u0_u2_u5_n104 ) , .ZN( u0_u2_u5_n131 ) );
  INV_X1 u0_u2_u5_U74 (.A( u0_u2_u5_n102 ) , .ZN( u0_u2_u5_n195 ) );
  OAI221_X1 u0_u2_u5_U75 (.A( u0_u2_u5_n101 ) , .ZN( u0_u2_u5_n102 ) , .C2( u0_u2_u5_n115 ) , .C1( u0_u2_u5_n126 ) , .B1( u0_u2_u5_n134 ) , .B2( u0_u2_u5_n160 ) );
  OAI21_X1 u0_u2_u5_U76 (.ZN( u0_u2_u5_n101 ) , .B1( u0_u2_u5_n137 ) , .A( u0_u2_u5_n146 ) , .B2( u0_u2_u5_n147 ) );
  NOR2_X1 u0_u2_u5_U77 (.A2( u0_u2_X_34 ) , .A1( u0_u2_X_35 ) , .ZN( u0_u2_u5_n145 ) );
  NOR2_X1 u0_u2_u5_U78 (.A2( u0_u2_X_34 ) , .ZN( u0_u2_u5_n146 ) , .A1( u0_u2_u5_n171 ) );
  NOR2_X1 u0_u2_u5_U79 (.A2( u0_u2_X_31 ) , .A1( u0_u2_X_32 ) , .ZN( u0_u2_u5_n103 ) );
  NOR3_X1 u0_u2_u5_U8 (.A2( u0_u2_u5_n147 ) , .A1( u0_u2_u5_n148 ) , .ZN( u0_u2_u5_n149 ) , .A3( u0_u2_u5_n194 ) );
  NOR2_X1 u0_u2_u5_U80 (.A2( u0_u2_X_36 ) , .ZN( u0_u2_u5_n105 ) , .A1( u0_u2_u5_n180 ) );
  NOR2_X1 u0_u2_u5_U81 (.A2( u0_u2_X_33 ) , .ZN( u0_u2_u5_n108 ) , .A1( u0_u2_u5_n170 ) );
  NOR2_X1 u0_u2_u5_U82 (.A2( u0_u2_X_33 ) , .A1( u0_u2_X_36 ) , .ZN( u0_u2_u5_n107 ) );
  NOR2_X1 u0_u2_u5_U83 (.A2( u0_u2_X_31 ) , .ZN( u0_u2_u5_n104 ) , .A1( u0_u2_u5_n181 ) );
  NAND2_X1 u0_u2_u5_U84 (.A2( u0_u2_X_34 ) , .A1( u0_u2_X_35 ) , .ZN( u0_u2_u5_n153 ) );
  NAND2_X1 u0_u2_u5_U85 (.A1( u0_u2_X_34 ) , .ZN( u0_u2_u5_n126 ) , .A2( u0_u2_u5_n171 ) );
  AND2_X1 u0_u2_u5_U86 (.A1( u0_u2_X_31 ) , .A2( u0_u2_X_32 ) , .ZN( u0_u2_u5_n106 ) );
  AND2_X1 u0_u2_u5_U87 (.A1( u0_u2_X_31 ) , .ZN( u0_u2_u5_n109 ) , .A2( u0_u2_u5_n181 ) );
  INV_X1 u0_u2_u5_U88 (.A( u0_u2_X_33 ) , .ZN( u0_u2_u5_n180 ) );
  INV_X1 u0_u2_u5_U89 (.A( u0_u2_X_35 ) , .ZN( u0_u2_u5_n171 ) );
  NOR2_X1 u0_u2_u5_U9 (.ZN( u0_u2_u5_n135 ) , .A1( u0_u2_u5_n173 ) , .A2( u0_u2_u5_n176 ) );
  INV_X1 u0_u2_u5_U90 (.A( u0_u2_X_36 ) , .ZN( u0_u2_u5_n170 ) );
  INV_X1 u0_u2_u5_U91 (.A( u0_u2_X_32 ) , .ZN( u0_u2_u5_n181 ) );
  NAND4_X1 u0_u2_u5_U92 (.ZN( u0_out2_19 ) , .A4( u0_u2_u5_n166 ) , .A3( u0_u2_u5_n167 ) , .A2( u0_u2_u5_n168 ) , .A1( u0_u2_u5_n169 ) );
  AOI22_X1 u0_u2_u5_U93 (.B2( u0_u2_u5_n145 ) , .A2( u0_u2_u5_n146 ) , .ZN( u0_u2_u5_n167 ) , .B1( u0_u2_u5_n182 ) , .A1( u0_u2_u5_n189 ) );
  NOR4_X1 u0_u2_u5_U94 (.A4( u0_u2_u5_n162 ) , .A3( u0_u2_u5_n163 ) , .A2( u0_u2_u5_n164 ) , .A1( u0_u2_u5_n165 ) , .ZN( u0_u2_u5_n166 ) );
  NAND4_X1 u0_u2_u5_U95 (.ZN( u0_out2_11 ) , .A4( u0_u2_u5_n143 ) , .A3( u0_u2_u5_n144 ) , .A2( u0_u2_u5_n169 ) , .A1( u0_u2_u5_n196 ) );
  AOI22_X1 u0_u2_u5_U96 (.A2( u0_u2_u5_n132 ) , .ZN( u0_u2_u5_n144 ) , .B2( u0_u2_u5_n145 ) , .B1( u0_u2_u5_n184 ) , .A1( u0_u2_u5_n194 ) );
  NOR3_X1 u0_u2_u5_U97 (.A3( u0_u2_u5_n141 ) , .A1( u0_u2_u5_n142 ) , .ZN( u0_u2_u5_n143 ) , .A2( u0_u2_u5_n191 ) );
  NAND4_X1 u0_u2_u5_U98 (.ZN( u0_out2_4 ) , .A4( u0_u2_u5_n112 ) , .A2( u0_u2_u5_n113 ) , .A1( u0_u2_u5_n114 ) , .A3( u0_u2_u5_n195 ) );
  AOI211_X1 u0_u2_u5_U99 (.A( u0_u2_u5_n110 ) , .C1( u0_u2_u5_n111 ) , .ZN( u0_u2_u5_n112 ) , .B( u0_u2_u5_n118 ) , .C2( u0_u2_u5_n177 ) );
  XOR2_X1 u0_u3_U20 (.B( u0_K4_36 ) , .A( u0_R2_25 ) , .Z( u0_u3_X_36 ) );
  XOR2_X1 u0_u3_U21 (.B( u0_K4_35 ) , .A( u0_R2_24 ) , .Z( u0_u3_X_35 ) );
  XOR2_X1 u0_u3_U22 (.B( u0_K4_34 ) , .A( u0_R2_23 ) , .Z( u0_u3_X_34 ) );
  XOR2_X1 u0_u3_U23 (.B( u0_K4_33 ) , .A( u0_R2_22 ) , .Z( u0_u3_X_33 ) );
  XOR2_X1 u0_u3_U24 (.B( u0_K4_32 ) , .A( u0_R2_21 ) , .Z( u0_u3_X_32 ) );
  XOR2_X1 u0_u3_U25 (.B( u0_K4_31 ) , .A( u0_R2_20 ) , .Z( u0_u3_X_31 ) );
  INV_X1 u0_u3_u5_U10 (.A( u0_u3_u5_n121 ) , .ZN( u0_u3_u5_n177 ) );
  NOR3_X1 u0_u3_u5_U100 (.A3( u0_u3_u5_n141 ) , .A1( u0_u3_u5_n142 ) , .ZN( u0_u3_u5_n143 ) , .A2( u0_u3_u5_n191 ) );
  NAND4_X1 u0_u3_u5_U101 (.ZN( u0_out3_4 ) , .A4( u0_u3_u5_n112 ) , .A2( u0_u3_u5_n113 ) , .A1( u0_u3_u5_n114 ) , .A3( u0_u3_u5_n195 ) );
  AOI211_X1 u0_u3_u5_U102 (.A( u0_u3_u5_n110 ) , .C1( u0_u3_u5_n111 ) , .ZN( u0_u3_u5_n112 ) , .B( u0_u3_u5_n118 ) , .C2( u0_u3_u5_n177 ) );
  AOI222_X1 u0_u3_u5_U103 (.ZN( u0_u3_u5_n113 ) , .A1( u0_u3_u5_n131 ) , .C1( u0_u3_u5_n148 ) , .B2( u0_u3_u5_n174 ) , .C2( u0_u3_u5_n178 ) , .A2( u0_u3_u5_n179 ) , .B1( u0_u3_u5_n99 ) );
  NAND3_X1 u0_u3_u5_U104 (.A2( u0_u3_u5_n154 ) , .A3( u0_u3_u5_n158 ) , .A1( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n99 ) );
  NOR2_X1 u0_u3_u5_U11 (.ZN( u0_u3_u5_n160 ) , .A2( u0_u3_u5_n173 ) , .A1( u0_u3_u5_n177 ) );
  INV_X1 u0_u3_u5_U12 (.A( u0_u3_u5_n150 ) , .ZN( u0_u3_u5_n174 ) );
  AOI21_X1 u0_u3_u5_U13 (.A( u0_u3_u5_n160 ) , .B2( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n162 ) , .B1( u0_u3_u5_n192 ) );
  INV_X1 u0_u3_u5_U14 (.A( u0_u3_u5_n159 ) , .ZN( u0_u3_u5_n192 ) );
  AOI21_X1 u0_u3_u5_U15 (.A( u0_u3_u5_n156 ) , .B2( u0_u3_u5_n157 ) , .B1( u0_u3_u5_n158 ) , .ZN( u0_u3_u5_n163 ) );
  AOI21_X1 u0_u3_u5_U16 (.B2( u0_u3_u5_n139 ) , .B1( u0_u3_u5_n140 ) , .ZN( u0_u3_u5_n141 ) , .A( u0_u3_u5_n150 ) );
  OAI21_X1 u0_u3_u5_U17 (.A( u0_u3_u5_n133 ) , .B2( u0_u3_u5_n134 ) , .B1( u0_u3_u5_n135 ) , .ZN( u0_u3_u5_n142 ) );
  OAI21_X1 u0_u3_u5_U18 (.ZN( u0_u3_u5_n133 ) , .B2( u0_u3_u5_n147 ) , .A( u0_u3_u5_n173 ) , .B1( u0_u3_u5_n188 ) );
  NAND2_X1 u0_u3_u5_U19 (.A2( u0_u3_u5_n119 ) , .A1( u0_u3_u5_n123 ) , .ZN( u0_u3_u5_n137 ) );
  INV_X1 u0_u3_u5_U20 (.A( u0_u3_u5_n155 ) , .ZN( u0_u3_u5_n194 ) );
  NAND2_X1 u0_u3_u5_U21 (.A1( u0_u3_u5_n121 ) , .ZN( u0_u3_u5_n132 ) , .A2( u0_u3_u5_n172 ) );
  NAND2_X1 u0_u3_u5_U22 (.A2( u0_u3_u5_n122 ) , .ZN( u0_u3_u5_n136 ) , .A1( u0_u3_u5_n154 ) );
  NAND2_X1 u0_u3_u5_U23 (.A2( u0_u3_u5_n119 ) , .A1( u0_u3_u5_n120 ) , .ZN( u0_u3_u5_n159 ) );
  INV_X1 u0_u3_u5_U24 (.A( u0_u3_u5_n156 ) , .ZN( u0_u3_u5_n175 ) );
  INV_X1 u0_u3_u5_U25 (.A( u0_u3_u5_n158 ) , .ZN( u0_u3_u5_n188 ) );
  INV_X1 u0_u3_u5_U26 (.A( u0_u3_u5_n152 ) , .ZN( u0_u3_u5_n179 ) );
  INV_X1 u0_u3_u5_U27 (.A( u0_u3_u5_n140 ) , .ZN( u0_u3_u5_n182 ) );
  INV_X1 u0_u3_u5_U28 (.A( u0_u3_u5_n151 ) , .ZN( u0_u3_u5_n183 ) );
  INV_X1 u0_u3_u5_U29 (.A( u0_u3_u5_n123 ) , .ZN( u0_u3_u5_n185 ) );
  NOR2_X1 u0_u3_u5_U3 (.ZN( u0_u3_u5_n134 ) , .A1( u0_u3_u5_n183 ) , .A2( u0_u3_u5_n190 ) );
  INV_X1 u0_u3_u5_U30 (.A( u0_u3_u5_n161 ) , .ZN( u0_u3_u5_n184 ) );
  INV_X1 u0_u3_u5_U31 (.A( u0_u3_u5_n139 ) , .ZN( u0_u3_u5_n189 ) );
  INV_X1 u0_u3_u5_U32 (.A( u0_u3_u5_n157 ) , .ZN( u0_u3_u5_n190 ) );
  INV_X1 u0_u3_u5_U33 (.A( u0_u3_u5_n120 ) , .ZN( u0_u3_u5_n193 ) );
  NAND2_X1 u0_u3_u5_U34 (.ZN( u0_u3_u5_n111 ) , .A1( u0_u3_u5_n140 ) , .A2( u0_u3_u5_n155 ) );
  INV_X1 u0_u3_u5_U35 (.A( u0_u3_u5_n117 ) , .ZN( u0_u3_u5_n196 ) );
  OAI221_X1 u0_u3_u5_U36 (.A( u0_u3_u5_n116 ) , .ZN( u0_u3_u5_n117 ) , .B2( u0_u3_u5_n119 ) , .C1( u0_u3_u5_n153 ) , .C2( u0_u3_u5_n158 ) , .B1( u0_u3_u5_n172 ) );
  AOI222_X1 u0_u3_u5_U37 (.ZN( u0_u3_u5_n116 ) , .B2( u0_u3_u5_n145 ) , .C1( u0_u3_u5_n148 ) , .A2( u0_u3_u5_n174 ) , .C2( u0_u3_u5_n177 ) , .B1( u0_u3_u5_n187 ) , .A1( u0_u3_u5_n193 ) );
  INV_X1 u0_u3_u5_U38 (.A( u0_u3_u5_n115 ) , .ZN( u0_u3_u5_n187 ) );
  NOR2_X1 u0_u3_u5_U39 (.ZN( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n170 ) , .A2( u0_u3_u5_n180 ) );
  INV_X1 u0_u3_u5_U4 (.A( u0_u3_u5_n138 ) , .ZN( u0_u3_u5_n191 ) );
  AOI22_X1 u0_u3_u5_U40 (.B2( u0_u3_u5_n131 ) , .A2( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n169 ) , .B1( u0_u3_u5_n174 ) , .A1( u0_u3_u5_n185 ) );
  NOR2_X1 u0_u3_u5_U41 (.A1( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n150 ) , .A2( u0_u3_u5_n173 ) );
  AOI21_X1 u0_u3_u5_U42 (.A( u0_u3_u5_n118 ) , .B2( u0_u3_u5_n145 ) , .ZN( u0_u3_u5_n168 ) , .B1( u0_u3_u5_n186 ) );
  INV_X1 u0_u3_u5_U43 (.A( u0_u3_u5_n122 ) , .ZN( u0_u3_u5_n186 ) );
  NOR2_X1 u0_u3_u5_U44 (.A1( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n152 ) , .A2( u0_u3_u5_n176 ) );
  NOR2_X1 u0_u3_u5_U45 (.A1( u0_u3_u5_n115 ) , .ZN( u0_u3_u5_n118 ) , .A2( u0_u3_u5_n153 ) );
  NOR2_X1 u0_u3_u5_U46 (.A2( u0_u3_u5_n145 ) , .ZN( u0_u3_u5_n156 ) , .A1( u0_u3_u5_n174 ) );
  NOR2_X1 u0_u3_u5_U47 (.ZN( u0_u3_u5_n121 ) , .A2( u0_u3_u5_n145 ) , .A1( u0_u3_u5_n176 ) );
  AOI22_X1 u0_u3_u5_U48 (.ZN( u0_u3_u5_n114 ) , .A2( u0_u3_u5_n137 ) , .A1( u0_u3_u5_n145 ) , .B2( u0_u3_u5_n175 ) , .B1( u0_u3_u5_n193 ) );
  OAI211_X1 u0_u3_u5_U49 (.B( u0_u3_u5_n124 ) , .A( u0_u3_u5_n125 ) , .C2( u0_u3_u5_n126 ) , .C1( u0_u3_u5_n127 ) , .ZN( u0_u3_u5_n128 ) );
  OAI21_X1 u0_u3_u5_U5 (.B2( u0_u3_u5_n136 ) , .B1( u0_u3_u5_n137 ) , .ZN( u0_u3_u5_n138 ) , .A( u0_u3_u5_n177 ) );
  NOR3_X1 u0_u3_u5_U50 (.ZN( u0_u3_u5_n127 ) , .A1( u0_u3_u5_n136 ) , .A3( u0_u3_u5_n148 ) , .A2( u0_u3_u5_n182 ) );
  OAI21_X1 u0_u3_u5_U51 (.ZN( u0_u3_u5_n124 ) , .A( u0_u3_u5_n177 ) , .B2( u0_u3_u5_n183 ) , .B1( u0_u3_u5_n189 ) );
  OAI21_X1 u0_u3_u5_U52 (.ZN( u0_u3_u5_n125 ) , .A( u0_u3_u5_n174 ) , .B2( u0_u3_u5_n185 ) , .B1( u0_u3_u5_n190 ) );
  AOI21_X1 u0_u3_u5_U53 (.A( u0_u3_u5_n153 ) , .B2( u0_u3_u5_n154 ) , .B1( u0_u3_u5_n155 ) , .ZN( u0_u3_u5_n164 ) );
  AOI21_X1 u0_u3_u5_U54 (.ZN( u0_u3_u5_n110 ) , .B1( u0_u3_u5_n122 ) , .B2( u0_u3_u5_n139 ) , .A( u0_u3_u5_n153 ) );
  INV_X1 u0_u3_u5_U55 (.A( u0_u3_u5_n153 ) , .ZN( u0_u3_u5_n176 ) );
  INV_X1 u0_u3_u5_U56 (.A( u0_u3_u5_n126 ) , .ZN( u0_u3_u5_n173 ) );
  AND2_X1 u0_u3_u5_U57 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n147 ) );
  AND2_X1 u0_u3_u5_U58 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n148 ) );
  NAND2_X1 u0_u3_u5_U59 (.A1( u0_u3_u5_n105 ) , .A2( u0_u3_u5_n106 ) , .ZN( u0_u3_u5_n158 ) );
  INV_X1 u0_u3_u5_U6 (.A( u0_u3_u5_n135 ) , .ZN( u0_u3_u5_n178 ) );
  NAND2_X1 u0_u3_u5_U60 (.A2( u0_u3_u5_n108 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n139 ) );
  NAND2_X1 u0_u3_u5_U61 (.A1( u0_u3_u5_n106 ) , .A2( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n119 ) );
  NAND2_X1 u0_u3_u5_U62 (.A2( u0_u3_u5_n103 ) , .A1( u0_u3_u5_n105 ) , .ZN( u0_u3_u5_n140 ) );
  NAND2_X1 u0_u3_u5_U63 (.A2( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n105 ) , .ZN( u0_u3_u5_n155 ) );
  NAND2_X1 u0_u3_u5_U64 (.A2( u0_u3_u5_n106 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n122 ) );
  NAND2_X1 u0_u3_u5_U65 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n106 ) , .ZN( u0_u3_u5_n115 ) );
  NAND2_X1 u0_u3_u5_U66 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n103 ) , .ZN( u0_u3_u5_n161 ) );
  NAND2_X1 u0_u3_u5_U67 (.A1( u0_u3_u5_n105 ) , .A2( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n154 ) );
  INV_X1 u0_u3_u5_U68 (.A( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n172 ) );
  NAND2_X1 u0_u3_u5_U69 (.A1( u0_u3_u5_n103 ) , .A2( u0_u3_u5_n108 ) , .ZN( u0_u3_u5_n123 ) );
  OAI22_X1 u0_u3_u5_U7 (.B2( u0_u3_u5_n149 ) , .B1( u0_u3_u5_n150 ) , .A2( u0_u3_u5_n151 ) , .A1( u0_u3_u5_n152 ) , .ZN( u0_u3_u5_n165 ) );
  NAND2_X1 u0_u3_u5_U70 (.A2( u0_u3_u5_n103 ) , .A1( u0_u3_u5_n107 ) , .ZN( u0_u3_u5_n151 ) );
  NAND2_X1 u0_u3_u5_U71 (.A2( u0_u3_u5_n107 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n120 ) );
  NAND2_X1 u0_u3_u5_U72 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n109 ) , .ZN( u0_u3_u5_n157 ) );
  AND2_X1 u0_u3_u5_U73 (.A2( u0_u3_u5_n100 ) , .A1( u0_u3_u5_n104 ) , .ZN( u0_u3_u5_n131 ) );
  INV_X1 u0_u3_u5_U74 (.A( u0_u3_u5_n102 ) , .ZN( u0_u3_u5_n195 ) );
  OAI221_X1 u0_u3_u5_U75 (.A( u0_u3_u5_n101 ) , .ZN( u0_u3_u5_n102 ) , .C2( u0_u3_u5_n115 ) , .C1( u0_u3_u5_n126 ) , .B1( u0_u3_u5_n134 ) , .B2( u0_u3_u5_n160 ) );
  OAI21_X1 u0_u3_u5_U76 (.ZN( u0_u3_u5_n101 ) , .B1( u0_u3_u5_n137 ) , .A( u0_u3_u5_n146 ) , .B2( u0_u3_u5_n147 ) );
  NOR2_X1 u0_u3_u5_U77 (.A2( u0_u3_X_34 ) , .A1( u0_u3_X_35 ) , .ZN( u0_u3_u5_n145 ) );
  NOR2_X1 u0_u3_u5_U78 (.A2( u0_u3_X_34 ) , .ZN( u0_u3_u5_n146 ) , .A1( u0_u3_u5_n171 ) );
  NOR2_X1 u0_u3_u5_U79 (.A2( u0_u3_X_31 ) , .A1( u0_u3_X_32 ) , .ZN( u0_u3_u5_n103 ) );
  NOR3_X1 u0_u3_u5_U8 (.A2( u0_u3_u5_n147 ) , .A1( u0_u3_u5_n148 ) , .ZN( u0_u3_u5_n149 ) , .A3( u0_u3_u5_n194 ) );
  NOR2_X1 u0_u3_u5_U80 (.A2( u0_u3_X_36 ) , .ZN( u0_u3_u5_n105 ) , .A1( u0_u3_u5_n180 ) );
  NOR2_X1 u0_u3_u5_U81 (.A2( u0_u3_X_33 ) , .ZN( u0_u3_u5_n108 ) , .A1( u0_u3_u5_n170 ) );
  NOR2_X1 u0_u3_u5_U82 (.A2( u0_u3_X_33 ) , .A1( u0_u3_X_36 ) , .ZN( u0_u3_u5_n107 ) );
  NOR2_X1 u0_u3_u5_U83 (.A2( u0_u3_X_31 ) , .ZN( u0_u3_u5_n104 ) , .A1( u0_u3_u5_n181 ) );
  NAND2_X1 u0_u3_u5_U84 (.A2( u0_u3_X_34 ) , .A1( u0_u3_X_35 ) , .ZN( u0_u3_u5_n153 ) );
  NAND2_X1 u0_u3_u5_U85 (.A1( u0_u3_X_34 ) , .ZN( u0_u3_u5_n126 ) , .A2( u0_u3_u5_n171 ) );
  AND2_X1 u0_u3_u5_U86 (.A1( u0_u3_X_31 ) , .A2( u0_u3_X_32 ) , .ZN( u0_u3_u5_n106 ) );
  AND2_X1 u0_u3_u5_U87 (.A1( u0_u3_X_31 ) , .ZN( u0_u3_u5_n109 ) , .A2( u0_u3_u5_n181 ) );
  INV_X1 u0_u3_u5_U88 (.A( u0_u3_X_33 ) , .ZN( u0_u3_u5_n180 ) );
  INV_X1 u0_u3_u5_U89 (.A( u0_u3_X_35 ) , .ZN( u0_u3_u5_n171 ) );
  NOR2_X1 u0_u3_u5_U9 (.ZN( u0_u3_u5_n135 ) , .A1( u0_u3_u5_n173 ) , .A2( u0_u3_u5_n176 ) );
  INV_X1 u0_u3_u5_U90 (.A( u0_u3_X_36 ) , .ZN( u0_u3_u5_n170 ) );
  INV_X1 u0_u3_u5_U91 (.A( u0_u3_X_32 ) , .ZN( u0_u3_u5_n181 ) );
  NAND4_X1 u0_u3_u5_U92 (.ZN( u0_out3_29 ) , .A4( u0_u3_u5_n129 ) , .A3( u0_u3_u5_n130 ) , .A2( u0_u3_u5_n168 ) , .A1( u0_u3_u5_n196 ) );
  AOI221_X1 u0_u3_u5_U93 (.A( u0_u3_u5_n128 ) , .ZN( u0_u3_u5_n129 ) , .C2( u0_u3_u5_n132 ) , .B2( u0_u3_u5_n159 ) , .B1( u0_u3_u5_n176 ) , .C1( u0_u3_u5_n184 ) );
  AOI222_X1 u0_u3_u5_U94 (.ZN( u0_u3_u5_n130 ) , .A2( u0_u3_u5_n146 ) , .B1( u0_u3_u5_n147 ) , .C2( u0_u3_u5_n175 ) , .B2( u0_u3_u5_n179 ) , .A1( u0_u3_u5_n188 ) , .C1( u0_u3_u5_n194 ) );
  NAND4_X1 u0_u3_u5_U95 (.ZN( u0_out3_19 ) , .A4( u0_u3_u5_n166 ) , .A3( u0_u3_u5_n167 ) , .A2( u0_u3_u5_n168 ) , .A1( u0_u3_u5_n169 ) );
  AOI22_X1 u0_u3_u5_U96 (.B2( u0_u3_u5_n145 ) , .A2( u0_u3_u5_n146 ) , .ZN( u0_u3_u5_n167 ) , .B1( u0_u3_u5_n182 ) , .A1( u0_u3_u5_n189 ) );
  NOR4_X1 u0_u3_u5_U97 (.A4( u0_u3_u5_n162 ) , .A3( u0_u3_u5_n163 ) , .A2( u0_u3_u5_n164 ) , .A1( u0_u3_u5_n165 ) , .ZN( u0_u3_u5_n166 ) );
  NAND4_X1 u0_u3_u5_U98 (.ZN( u0_out3_11 ) , .A4( u0_u3_u5_n143 ) , .A3( u0_u3_u5_n144 ) , .A2( u0_u3_u5_n169 ) , .A1( u0_u3_u5_n196 ) );
  AOI22_X1 u0_u3_u5_U99 (.A2( u0_u3_u5_n132 ) , .ZN( u0_u3_u5_n144 ) , .B2( u0_u3_u5_n145 ) , .B1( u0_u3_u5_n184 ) , .A1( u0_u3_u5_n194 ) );
  XOR2_X1 u0_u6_U10 (.B( u0_K7_45 ) , .A( u0_R5_30 ) , .Z( u0_u6_X_45 ) );
  XOR2_X1 u0_u6_U11 (.B( u0_K7_44 ) , .A( u0_R5_29 ) , .Z( u0_u6_X_44 ) );
  XOR2_X1 u0_u6_U12 (.B( u0_K7_43 ) , .A( u0_R5_28 ) , .Z( u0_u6_X_43 ) );
  XOR2_X1 u0_u6_U13 (.B( u0_K7_42 ) , .A( u0_R5_29 ) , .Z( u0_u6_X_42 ) );
  XOR2_X1 u0_u6_U14 (.B( u0_K7_41 ) , .A( u0_R5_28 ) , .Z( u0_u6_X_41 ) );
  XOR2_X1 u0_u6_U15 (.B( u0_K7_40 ) , .A( u0_R5_27 ) , .Z( u0_u6_X_40 ) );
  XOR2_X1 u0_u6_U16 (.B( u0_K7_3 ) , .A( u0_R5_2 ) , .Z( u0_u6_X_3 ) );
  XOR2_X1 u0_u6_U17 (.B( u0_K7_39 ) , .A( u0_R5_26 ) , .Z( u0_u6_X_39 ) );
  XOR2_X1 u0_u6_U18 (.B( u0_K7_38 ) , .A( u0_R5_25 ) , .Z( u0_u6_X_38 ) );
  XOR2_X1 u0_u6_U19 (.B( u0_K7_37 ) , .A( u0_R5_24 ) , .Z( u0_u6_X_37 ) );
  XOR2_X1 u0_u6_U20 (.B( u0_K7_36 ) , .A( u0_R5_25 ) , .Z( u0_u6_X_36 ) );
  XOR2_X1 u0_u6_U21 (.B( u0_K7_35 ) , .A( u0_R5_24 ) , .Z( u0_u6_X_35 ) );
  XOR2_X1 u0_u6_U22 (.B( u0_K7_34 ) , .A( u0_R5_23 ) , .Z( u0_u6_X_34 ) );
  XOR2_X1 u0_u6_U23 (.B( u0_K7_33 ) , .A( u0_R5_22 ) , .Z( u0_u6_X_33 ) );
  XOR2_X1 u0_u6_U24 (.B( u0_K7_32 ) , .A( u0_R5_21 ) , .Z( u0_u6_X_32 ) );
  XOR2_X1 u0_u6_U25 (.B( u0_K7_31 ) , .A( u0_R5_20 ) , .Z( u0_u6_X_31 ) );
  XOR2_X1 u0_u6_U27 (.B( u0_K7_2 ) , .A( u0_R5_1 ) , .Z( u0_u6_X_2 ) );
  XOR2_X1 u0_u6_U38 (.B( u0_K7_1 ) , .A( u0_R5_32 ) , .Z( u0_u6_X_1 ) );
  XOR2_X1 u0_u6_U5 (.B( u0_K7_5 ) , .A( u0_R5_4 ) , .Z( u0_u6_X_5 ) );
  XOR2_X1 u0_u6_U6 (.B( u0_K7_4 ) , .A( u0_R5_3 ) , .Z( u0_u6_X_4 ) );
  XOR2_X1 u0_u6_U7 (.B( u0_K7_48 ) , .A( u0_R5_1 ) , .Z( u0_u6_X_48 ) );
  XOR2_X1 u0_u6_U8 (.B( u0_K7_47 ) , .A( u0_R5_32 ) , .Z( u0_u6_X_47 ) );
  XOR2_X1 u0_u6_U9 (.B( u0_K7_46 ) , .A( u0_R5_31 ) , .Z( u0_u6_X_46 ) );
  NAND2_X1 u0_u6_u0_U10 (.ZN( u0_u6_u0_n113 ) , .A1( u0_u6_u0_n139 ) , .A2( u0_u6_u0_n149 ) );
  AND2_X1 u0_u6_u0_U11 (.A1( u0_u6_u0_n131 ) , .ZN( u0_u6_u0_n141 ) , .A2( u0_u6_u0_n150 ) );
  AND2_X1 u0_u6_u0_U12 (.ZN( u0_u6_u0_n107 ) , .A1( u0_u6_u0_n130 ) , .A2( u0_u6_u0_n140 ) );
  AND2_X1 u0_u6_u0_U13 (.A2( u0_u6_u0_n129 ) , .A1( u0_u6_u0_n130 ) , .ZN( u0_u6_u0_n151 ) );
  AND2_X1 u0_u6_u0_U14 (.A1( u0_u6_u0_n108 ) , .A2( u0_u6_u0_n125 ) , .ZN( u0_u6_u0_n145 ) );
  INV_X1 u0_u6_u0_U15 (.A( u0_u6_u0_n143 ) , .ZN( u0_u6_u0_n173 ) );
  NOR2_X1 u0_u6_u0_U16 (.A2( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n147 ) , .A1( u0_u6_u0_n160 ) );
  AOI21_X1 u0_u6_u0_U17 (.B1( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n132 ) , .A( u0_u6_u0_n165 ) , .B2( u0_u6_u0_n93 ) );
  OAI221_X1 u0_u6_u0_U18 (.C1( u0_u6_u0_n121 ) , .ZN( u0_u6_u0_n122 ) , .B2( u0_u6_u0_n127 ) , .A( u0_u6_u0_n143 ) , .B1( u0_u6_u0_n144 ) , .C2( u0_u6_u0_n147 ) );
  OAI22_X1 u0_u6_u0_U19 (.B1( u0_u6_u0_n125 ) , .ZN( u0_u6_u0_n126 ) , .A1( u0_u6_u0_n138 ) , .A2( u0_u6_u0_n146 ) , .B2( u0_u6_u0_n147 ) );
  OAI22_X1 u0_u6_u0_U20 (.B1( u0_u6_u0_n131 ) , .A1( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n147 ) , .A2( u0_u6_u0_n90 ) , .ZN( u0_u6_u0_n91 ) );
  AND3_X1 u0_u6_u0_U21 (.A3( u0_u6_u0_n121 ) , .A2( u0_u6_u0_n125 ) , .A1( u0_u6_u0_n148 ) , .ZN( u0_u6_u0_n90 ) );
  NOR2_X1 u0_u6_u0_U22 (.A1( u0_u6_u0_n163 ) , .A2( u0_u6_u0_n164 ) , .ZN( u0_u6_u0_n95 ) );
  NOR2_X1 u0_u6_u0_U23 (.A1( u0_u6_u0_n120 ) , .ZN( u0_u6_u0_n143 ) , .A2( u0_u6_u0_n167 ) );
  OAI221_X1 u0_u6_u0_U24 (.C1( u0_u6_u0_n112 ) , .ZN( u0_u6_u0_n120 ) , .B1( u0_u6_u0_n138 ) , .B2( u0_u6_u0_n141 ) , .C2( u0_u6_u0_n147 ) , .A( u0_u6_u0_n172 ) );
  AOI211_X1 u0_u6_u0_U25 (.B( u0_u6_u0_n115 ) , .A( u0_u6_u0_n116 ) , .C2( u0_u6_u0_n117 ) , .C1( u0_u6_u0_n118 ) , .ZN( u0_u6_u0_n119 ) );
  AOI22_X1 u0_u6_u0_U26 (.B2( u0_u6_u0_n109 ) , .A2( u0_u6_u0_n110 ) , .ZN( u0_u6_u0_n111 ) , .B1( u0_u6_u0_n118 ) , .A1( u0_u6_u0_n160 ) );
  NAND2_X1 u0_u6_u0_U27 (.A1( u0_u6_u0_n100 ) , .A2( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n125 ) );
  INV_X1 u0_u6_u0_U28 (.A( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U29 (.A( u0_u6_u0_n118 ) , .ZN( u0_u6_u0_n158 ) );
  INV_X1 u0_u6_u0_U3 (.A( u0_u6_u0_n113 ) , .ZN( u0_u6_u0_n166 ) );
  AOI21_X1 u0_u6_u0_U30 (.B1( u0_u6_u0_n127 ) , .B2( u0_u6_u0_n129 ) , .A( u0_u6_u0_n138 ) , .ZN( u0_u6_u0_n96 ) );
  AOI21_X1 u0_u6_u0_U31 (.ZN( u0_u6_u0_n104 ) , .B1( u0_u6_u0_n107 ) , .B2( u0_u6_u0_n141 ) , .A( u0_u6_u0_n144 ) );
  NAND2_X1 u0_u6_u0_U32 (.A2( u0_u6_u0_n102 ) , .A1( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n149 ) );
  NAND2_X1 u0_u6_u0_U33 (.A2( u0_u6_u0_n100 ) , .ZN( u0_u6_u0_n131 ) , .A1( u0_u6_u0_n92 ) );
  NAND2_X1 u0_u6_u0_U34 (.A2( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n114 ) , .A1( u0_u6_u0_n92 ) );
  NAND2_X1 u0_u6_u0_U35 (.A1( u0_u6_u0_n101 ) , .A2( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n150 ) );
  INV_X1 u0_u6_u0_U36 (.A( u0_u6_u0_n138 ) , .ZN( u0_u6_u0_n160 ) );
  NAND2_X1 u0_u6_u0_U37 (.A2( u0_u6_u0_n100 ) , .A1( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n139 ) );
  NAND2_X1 u0_u6_u0_U38 (.ZN( u0_u6_u0_n112 ) , .A2( u0_u6_u0_n92 ) , .A1( u0_u6_u0_n93 ) );
  NAND2_X1 u0_u6_u0_U39 (.A2( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n121 ) , .A1( u0_u6_u0_n93 ) );
  AOI21_X1 u0_u6_u0_U4 (.B1( u0_u6_u0_n114 ) , .ZN( u0_u6_u0_n115 ) , .B2( u0_u6_u0_n129 ) , .A( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U40 (.ZN( u0_u6_u0_n172 ) , .A( u0_u6_u0_n88 ) );
  OAI222_X1 u0_u6_u0_U41 (.C1( u0_u6_u0_n108 ) , .A1( u0_u6_u0_n125 ) , .B2( u0_u6_u0_n128 ) , .B1( u0_u6_u0_n144 ) , .A2( u0_u6_u0_n158 ) , .C2( u0_u6_u0_n161 ) , .ZN( u0_u6_u0_n88 ) );
  OR3_X1 u0_u6_u0_U42 (.A3( u0_u6_u0_n152 ) , .A2( u0_u6_u0_n153 ) , .A1( u0_u6_u0_n154 ) , .ZN( u0_u6_u0_n155 ) );
  AOI21_X1 u0_u6_u0_U43 (.A( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n145 ) , .B1( u0_u6_u0_n146 ) , .ZN( u0_u6_u0_n154 ) );
  AOI21_X1 u0_u6_u0_U44 (.B2( u0_u6_u0_n150 ) , .B1( u0_u6_u0_n151 ) , .ZN( u0_u6_u0_n152 ) , .A( u0_u6_u0_n158 ) );
  AOI21_X1 u0_u6_u0_U45 (.A( u0_u6_u0_n147 ) , .B2( u0_u6_u0_n148 ) , .B1( u0_u6_u0_n149 ) , .ZN( u0_u6_u0_n153 ) );
  INV_X1 u0_u6_u0_U46 (.ZN( u0_u6_u0_n171 ) , .A( u0_u6_u0_n99 ) );
  OAI211_X1 u0_u6_u0_U47 (.C2( u0_u6_u0_n140 ) , .C1( u0_u6_u0_n161 ) , .A( u0_u6_u0_n169 ) , .B( u0_u6_u0_n98 ) , .ZN( u0_u6_u0_n99 ) );
  AOI211_X1 u0_u6_u0_U48 (.C1( u0_u6_u0_n118 ) , .A( u0_u6_u0_n123 ) , .B( u0_u6_u0_n96 ) , .C2( u0_u6_u0_n97 ) , .ZN( u0_u6_u0_n98 ) );
  INV_X1 u0_u6_u0_U49 (.ZN( u0_u6_u0_n169 ) , .A( u0_u6_u0_n91 ) );
  NOR2_X1 u0_u6_u0_U5 (.A1( u0_u6_u0_n108 ) , .ZN( u0_u6_u0_n123 ) , .A2( u0_u6_u0_n158 ) );
  NOR2_X1 u0_u6_u0_U50 (.A2( u0_u6_X_4 ) , .A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n118 ) );
  NOR2_X1 u0_u6_u0_U51 (.A2( u0_u6_X_1 ) , .ZN( u0_u6_u0_n101 ) , .A1( u0_u6_u0_n163 ) );
  NAND2_X1 u0_u6_u0_U52 (.A2( u0_u6_X_4 ) , .A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n144 ) );
  NOR2_X1 u0_u6_u0_U53 (.A2( u0_u6_X_5 ) , .ZN( u0_u6_u0_n136 ) , .A1( u0_u6_u0_n159 ) );
  NAND2_X1 u0_u6_u0_U54 (.A1( u0_u6_X_5 ) , .ZN( u0_u6_u0_n138 ) , .A2( u0_u6_u0_n159 ) );
  AND2_X1 u0_u6_u0_U55 (.A2( u0_u6_X_3 ) , .A1( u0_u6_X_6 ) , .ZN( u0_u6_u0_n102 ) );
  INV_X1 u0_u6_u0_U56 (.A( u0_u6_X_4 ) , .ZN( u0_u6_u0_n159 ) );
  INV_X1 u0_u6_u0_U57 (.A( u0_u6_X_1 ) , .ZN( u0_u6_u0_n164 ) );
  INV_X1 u0_u6_u0_U58 (.A( u0_u6_X_3 ) , .ZN( u0_u6_u0_n162 ) );
  INV_X1 u0_u6_u0_U59 (.A( u0_u6_u0_n126 ) , .ZN( u0_u6_u0_n168 ) );
  AOI21_X1 u0_u6_u0_U6 (.B2( u0_u6_u0_n131 ) , .ZN( u0_u6_u0_n134 ) , .B1( u0_u6_u0_n151 ) , .A( u0_u6_u0_n158 ) );
  AOI211_X1 u0_u6_u0_U60 (.B( u0_u6_u0_n133 ) , .A( u0_u6_u0_n134 ) , .C2( u0_u6_u0_n135 ) , .C1( u0_u6_u0_n136 ) , .ZN( u0_u6_u0_n137 ) );
  INV_X1 u0_u6_u0_U61 (.ZN( u0_u6_u0_n174 ) , .A( u0_u6_u0_n89 ) );
  AOI211_X1 u0_u6_u0_U62 (.B( u0_u6_u0_n104 ) , .A( u0_u6_u0_n105 ) , .ZN( u0_u6_u0_n106 ) , .C2( u0_u6_u0_n113 ) , .C1( u0_u6_u0_n160 ) );
  OR4_X1 u0_u6_u0_U63 (.ZN( u0_out6_31 ) , .A4( u0_u6_u0_n155 ) , .A2( u0_u6_u0_n156 ) , .A1( u0_u6_u0_n157 ) , .A3( u0_u6_u0_n173 ) );
  AOI21_X1 u0_u6_u0_U64 (.A( u0_u6_u0_n138 ) , .B2( u0_u6_u0_n139 ) , .B1( u0_u6_u0_n140 ) , .ZN( u0_u6_u0_n157 ) );
  OR4_X1 u0_u6_u0_U65 (.ZN( u0_out6_17 ) , .A4( u0_u6_u0_n122 ) , .A2( u0_u6_u0_n123 ) , .A1( u0_u6_u0_n124 ) , .A3( u0_u6_u0_n170 ) );
  AOI21_X1 u0_u6_u0_U66 (.B2( u0_u6_u0_n107 ) , .ZN( u0_u6_u0_n124 ) , .B1( u0_u6_u0_n128 ) , .A( u0_u6_u0_n161 ) );
  INV_X1 u0_u6_u0_U67 (.A( u0_u6_u0_n111 ) , .ZN( u0_u6_u0_n170 ) );
  AOI21_X1 u0_u6_u0_U68 (.B2( u0_u6_u0_n141 ) , .B1( u0_u6_u0_n142 ) , .ZN( u0_u6_u0_n156 ) , .A( u0_u6_u0_n161 ) );
  AOI21_X1 u0_u6_u0_U69 (.ZN( u0_u6_u0_n116 ) , .B2( u0_u6_u0_n142 ) , .A( u0_u6_u0_n144 ) , .B1( u0_u6_u0_n166 ) );
  OAI21_X1 u0_u6_u0_U7 (.B1( u0_u6_u0_n150 ) , .B2( u0_u6_u0_n158 ) , .A( u0_u6_u0_n172 ) , .ZN( u0_u6_u0_n89 ) );
  NAND2_X1 u0_u6_u0_U70 (.ZN( u0_u6_u0_n148 ) , .A1( u0_u6_u0_n93 ) , .A2( u0_u6_u0_n95 ) );
  NAND2_X1 u0_u6_u0_U71 (.A1( u0_u6_u0_n100 ) , .ZN( u0_u6_u0_n129 ) , .A2( u0_u6_u0_n95 ) );
  NAND2_X1 u0_u6_u0_U72 (.A1( u0_u6_u0_n102 ) , .ZN( u0_u6_u0_n128 ) , .A2( u0_u6_u0_n95 ) );
  INV_X1 u0_u6_u0_U73 (.A( u0_u6_u0_n142 ) , .ZN( u0_u6_u0_n165 ) );
  NOR2_X1 u0_u6_u0_U74 (.A2( u0_u6_X_1 ) , .A1( u0_u6_X_2 ) , .ZN( u0_u6_u0_n92 ) );
  NOR2_X1 u0_u6_u0_U75 (.A2( u0_u6_X_2 ) , .ZN( u0_u6_u0_n103 ) , .A1( u0_u6_u0_n164 ) );
  INV_X1 u0_u6_u0_U76 (.A( u0_u6_X_2 ) , .ZN( u0_u6_u0_n163 ) );
  AOI21_X1 u0_u6_u0_U77 (.B1( u0_u6_u0_n132 ) , .ZN( u0_u6_u0_n133 ) , .A( u0_u6_u0_n144 ) , .B2( u0_u6_u0_n166 ) );
  OAI22_X1 u0_u6_u0_U78 (.ZN( u0_u6_u0_n105 ) , .A2( u0_u6_u0_n132 ) , .B1( u0_u6_u0_n146 ) , .A1( u0_u6_u0_n147 ) , .B2( u0_u6_u0_n161 ) );
  NAND2_X1 u0_u6_u0_U79 (.ZN( u0_u6_u0_n110 ) , .A2( u0_u6_u0_n132 ) , .A1( u0_u6_u0_n145 ) );
  AND2_X1 u0_u6_u0_U8 (.A1( u0_u6_u0_n114 ) , .A2( u0_u6_u0_n121 ) , .ZN( u0_u6_u0_n146 ) );
  INV_X1 u0_u6_u0_U80 (.A( u0_u6_u0_n119 ) , .ZN( u0_u6_u0_n167 ) );
  NAND2_X1 u0_u6_u0_U81 (.A2( u0_u6_u0_n103 ) , .ZN( u0_u6_u0_n140 ) , .A1( u0_u6_u0_n94 ) );
  NAND2_X1 u0_u6_u0_U82 (.A1( u0_u6_u0_n101 ) , .ZN( u0_u6_u0_n130 ) , .A2( u0_u6_u0_n94 ) );
  NAND2_X1 u0_u6_u0_U83 (.ZN( u0_u6_u0_n108 ) , .A1( u0_u6_u0_n92 ) , .A2( u0_u6_u0_n94 ) );
  AND2_X1 u0_u6_u0_U84 (.A1( u0_u6_X_6 ) , .A2( u0_u6_u0_n162 ) , .ZN( u0_u6_u0_n93 ) );
  NAND2_X1 u0_u6_u0_U85 (.ZN( u0_u6_u0_n142 ) , .A1( u0_u6_u0_n94 ) , .A2( u0_u6_u0_n95 ) );
  NOR2_X1 u0_u6_u0_U86 (.A2( u0_u6_X_6 ) , .ZN( u0_u6_u0_n100 ) , .A1( u0_u6_u0_n162 ) );
  NOR2_X1 u0_u6_u0_U87 (.A2( u0_u6_X_3 ) , .A1( u0_u6_X_6 ) , .ZN( u0_u6_u0_n94 ) );
  NAND3_X1 u0_u6_u0_U88 (.ZN( u0_out6_23 ) , .A3( u0_u6_u0_n137 ) , .A1( u0_u6_u0_n168 ) , .A2( u0_u6_u0_n171 ) );
  NAND3_X1 u0_u6_u0_U89 (.A3( u0_u6_u0_n127 ) , .A2( u0_u6_u0_n128 ) , .ZN( u0_u6_u0_n135 ) , .A1( u0_u6_u0_n150 ) );
  AND3_X1 u0_u6_u0_U9 (.A2( u0_u6_u0_n112 ) , .ZN( u0_u6_u0_n127 ) , .A3( u0_u6_u0_n130 ) , .A1( u0_u6_u0_n148 ) );
  NAND3_X1 u0_u6_u0_U90 (.ZN( u0_u6_u0_n117 ) , .A3( u0_u6_u0_n132 ) , .A2( u0_u6_u0_n139 ) , .A1( u0_u6_u0_n148 ) );
  NAND3_X1 u0_u6_u0_U91 (.ZN( u0_u6_u0_n109 ) , .A2( u0_u6_u0_n114 ) , .A3( u0_u6_u0_n140 ) , .A1( u0_u6_u0_n149 ) );
  NAND3_X1 u0_u6_u0_U92 (.ZN( u0_out6_9 ) , .A3( u0_u6_u0_n106 ) , .A2( u0_u6_u0_n171 ) , .A1( u0_u6_u0_n174 ) );
  NAND3_X1 u0_u6_u0_U93 (.A2( u0_u6_u0_n128 ) , .A1( u0_u6_u0_n132 ) , .A3( u0_u6_u0_n146 ) , .ZN( u0_u6_u0_n97 ) );
  INV_X1 u0_u6_u5_U10 (.A( u0_u6_u5_n121 ) , .ZN( u0_u6_u5_n177 ) );
  NOR3_X1 u0_u6_u5_U100 (.A3( u0_u6_u5_n141 ) , .A1( u0_u6_u5_n142 ) , .ZN( u0_u6_u5_n143 ) , .A2( u0_u6_u5_n191 ) );
  NAND4_X1 u0_u6_u5_U101 (.ZN( u0_out6_4 ) , .A4( u0_u6_u5_n112 ) , .A2( u0_u6_u5_n113 ) , .A1( u0_u6_u5_n114 ) , .A3( u0_u6_u5_n195 ) );
  AOI211_X1 u0_u6_u5_U102 (.A( u0_u6_u5_n110 ) , .C1( u0_u6_u5_n111 ) , .ZN( u0_u6_u5_n112 ) , .B( u0_u6_u5_n118 ) , .C2( u0_u6_u5_n177 ) );
  AOI222_X1 u0_u6_u5_U103 (.ZN( u0_u6_u5_n113 ) , .A1( u0_u6_u5_n131 ) , .C1( u0_u6_u5_n148 ) , .B2( u0_u6_u5_n174 ) , .C2( u0_u6_u5_n178 ) , .A2( u0_u6_u5_n179 ) , .B1( u0_u6_u5_n99 ) );
  NAND3_X1 u0_u6_u5_U104 (.A2( u0_u6_u5_n154 ) , .A3( u0_u6_u5_n158 ) , .A1( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n99 ) );
  NOR2_X1 u0_u6_u5_U11 (.ZN( u0_u6_u5_n160 ) , .A2( u0_u6_u5_n173 ) , .A1( u0_u6_u5_n177 ) );
  INV_X1 u0_u6_u5_U12 (.A( u0_u6_u5_n150 ) , .ZN( u0_u6_u5_n174 ) );
  AOI21_X1 u0_u6_u5_U13 (.A( u0_u6_u5_n160 ) , .B2( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n162 ) , .B1( u0_u6_u5_n192 ) );
  INV_X1 u0_u6_u5_U14 (.A( u0_u6_u5_n159 ) , .ZN( u0_u6_u5_n192 ) );
  AOI21_X1 u0_u6_u5_U15 (.A( u0_u6_u5_n156 ) , .B2( u0_u6_u5_n157 ) , .B1( u0_u6_u5_n158 ) , .ZN( u0_u6_u5_n163 ) );
  AOI21_X1 u0_u6_u5_U16 (.B2( u0_u6_u5_n139 ) , .B1( u0_u6_u5_n140 ) , .ZN( u0_u6_u5_n141 ) , .A( u0_u6_u5_n150 ) );
  OAI21_X1 u0_u6_u5_U17 (.A( u0_u6_u5_n133 ) , .B2( u0_u6_u5_n134 ) , .B1( u0_u6_u5_n135 ) , .ZN( u0_u6_u5_n142 ) );
  OAI21_X1 u0_u6_u5_U18 (.ZN( u0_u6_u5_n133 ) , .B2( u0_u6_u5_n147 ) , .A( u0_u6_u5_n173 ) , .B1( u0_u6_u5_n188 ) );
  NAND2_X1 u0_u6_u5_U19 (.A2( u0_u6_u5_n119 ) , .A1( u0_u6_u5_n123 ) , .ZN( u0_u6_u5_n137 ) );
  INV_X1 u0_u6_u5_U20 (.A( u0_u6_u5_n155 ) , .ZN( u0_u6_u5_n194 ) );
  NAND2_X1 u0_u6_u5_U21 (.A1( u0_u6_u5_n121 ) , .ZN( u0_u6_u5_n132 ) , .A2( u0_u6_u5_n172 ) );
  NAND2_X1 u0_u6_u5_U22 (.A2( u0_u6_u5_n122 ) , .ZN( u0_u6_u5_n136 ) , .A1( u0_u6_u5_n154 ) );
  NAND2_X1 u0_u6_u5_U23 (.A2( u0_u6_u5_n119 ) , .A1( u0_u6_u5_n120 ) , .ZN( u0_u6_u5_n159 ) );
  INV_X1 u0_u6_u5_U24 (.A( u0_u6_u5_n156 ) , .ZN( u0_u6_u5_n175 ) );
  INV_X1 u0_u6_u5_U25 (.A( u0_u6_u5_n158 ) , .ZN( u0_u6_u5_n188 ) );
  INV_X1 u0_u6_u5_U26 (.A( u0_u6_u5_n152 ) , .ZN( u0_u6_u5_n179 ) );
  INV_X1 u0_u6_u5_U27 (.A( u0_u6_u5_n140 ) , .ZN( u0_u6_u5_n182 ) );
  INV_X1 u0_u6_u5_U28 (.A( u0_u6_u5_n151 ) , .ZN( u0_u6_u5_n183 ) );
  INV_X1 u0_u6_u5_U29 (.A( u0_u6_u5_n123 ) , .ZN( u0_u6_u5_n185 ) );
  NOR2_X1 u0_u6_u5_U3 (.ZN( u0_u6_u5_n134 ) , .A1( u0_u6_u5_n183 ) , .A2( u0_u6_u5_n190 ) );
  INV_X1 u0_u6_u5_U30 (.A( u0_u6_u5_n161 ) , .ZN( u0_u6_u5_n184 ) );
  INV_X1 u0_u6_u5_U31 (.A( u0_u6_u5_n139 ) , .ZN( u0_u6_u5_n189 ) );
  INV_X1 u0_u6_u5_U32 (.A( u0_u6_u5_n157 ) , .ZN( u0_u6_u5_n190 ) );
  INV_X1 u0_u6_u5_U33 (.A( u0_u6_u5_n120 ) , .ZN( u0_u6_u5_n193 ) );
  NAND2_X1 u0_u6_u5_U34 (.ZN( u0_u6_u5_n111 ) , .A1( u0_u6_u5_n140 ) , .A2( u0_u6_u5_n155 ) );
  INV_X1 u0_u6_u5_U35 (.A( u0_u6_u5_n117 ) , .ZN( u0_u6_u5_n196 ) );
  OAI221_X1 u0_u6_u5_U36 (.A( u0_u6_u5_n116 ) , .ZN( u0_u6_u5_n117 ) , .B2( u0_u6_u5_n119 ) , .C1( u0_u6_u5_n153 ) , .C2( u0_u6_u5_n158 ) , .B1( u0_u6_u5_n172 ) );
  AOI222_X1 u0_u6_u5_U37 (.ZN( u0_u6_u5_n116 ) , .B2( u0_u6_u5_n145 ) , .C1( u0_u6_u5_n148 ) , .A2( u0_u6_u5_n174 ) , .C2( u0_u6_u5_n177 ) , .B1( u0_u6_u5_n187 ) , .A1( u0_u6_u5_n193 ) );
  INV_X1 u0_u6_u5_U38 (.A( u0_u6_u5_n115 ) , .ZN( u0_u6_u5_n187 ) );
  NOR2_X1 u0_u6_u5_U39 (.ZN( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n170 ) , .A2( u0_u6_u5_n180 ) );
  INV_X1 u0_u6_u5_U4 (.A( u0_u6_u5_n138 ) , .ZN( u0_u6_u5_n191 ) );
  AOI22_X1 u0_u6_u5_U40 (.B2( u0_u6_u5_n131 ) , .A2( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n169 ) , .B1( u0_u6_u5_n174 ) , .A1( u0_u6_u5_n185 ) );
  NOR2_X1 u0_u6_u5_U41 (.A1( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n150 ) , .A2( u0_u6_u5_n173 ) );
  AOI21_X1 u0_u6_u5_U42 (.A( u0_u6_u5_n118 ) , .B2( u0_u6_u5_n145 ) , .ZN( u0_u6_u5_n168 ) , .B1( u0_u6_u5_n186 ) );
  INV_X1 u0_u6_u5_U43 (.A( u0_u6_u5_n122 ) , .ZN( u0_u6_u5_n186 ) );
  NOR2_X1 u0_u6_u5_U44 (.A1( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n152 ) , .A2( u0_u6_u5_n176 ) );
  NOR2_X1 u0_u6_u5_U45 (.A1( u0_u6_u5_n115 ) , .ZN( u0_u6_u5_n118 ) , .A2( u0_u6_u5_n153 ) );
  NOR2_X1 u0_u6_u5_U46 (.A2( u0_u6_u5_n145 ) , .ZN( u0_u6_u5_n156 ) , .A1( u0_u6_u5_n174 ) );
  NOR2_X1 u0_u6_u5_U47 (.ZN( u0_u6_u5_n121 ) , .A2( u0_u6_u5_n145 ) , .A1( u0_u6_u5_n176 ) );
  AOI22_X1 u0_u6_u5_U48 (.ZN( u0_u6_u5_n114 ) , .A2( u0_u6_u5_n137 ) , .A1( u0_u6_u5_n145 ) , .B2( u0_u6_u5_n175 ) , .B1( u0_u6_u5_n193 ) );
  OAI211_X1 u0_u6_u5_U49 (.B( u0_u6_u5_n124 ) , .A( u0_u6_u5_n125 ) , .C2( u0_u6_u5_n126 ) , .C1( u0_u6_u5_n127 ) , .ZN( u0_u6_u5_n128 ) );
  OAI21_X1 u0_u6_u5_U5 (.B2( u0_u6_u5_n136 ) , .B1( u0_u6_u5_n137 ) , .ZN( u0_u6_u5_n138 ) , .A( u0_u6_u5_n177 ) );
  NOR3_X1 u0_u6_u5_U50 (.ZN( u0_u6_u5_n127 ) , .A1( u0_u6_u5_n136 ) , .A3( u0_u6_u5_n148 ) , .A2( u0_u6_u5_n182 ) );
  OAI21_X1 u0_u6_u5_U51 (.ZN( u0_u6_u5_n124 ) , .A( u0_u6_u5_n177 ) , .B2( u0_u6_u5_n183 ) , .B1( u0_u6_u5_n189 ) );
  OAI21_X1 u0_u6_u5_U52 (.ZN( u0_u6_u5_n125 ) , .A( u0_u6_u5_n174 ) , .B2( u0_u6_u5_n185 ) , .B1( u0_u6_u5_n190 ) );
  AOI21_X1 u0_u6_u5_U53 (.A( u0_u6_u5_n153 ) , .B2( u0_u6_u5_n154 ) , .B1( u0_u6_u5_n155 ) , .ZN( u0_u6_u5_n164 ) );
  AOI21_X1 u0_u6_u5_U54 (.ZN( u0_u6_u5_n110 ) , .B1( u0_u6_u5_n122 ) , .B2( u0_u6_u5_n139 ) , .A( u0_u6_u5_n153 ) );
  INV_X1 u0_u6_u5_U55 (.A( u0_u6_u5_n153 ) , .ZN( u0_u6_u5_n176 ) );
  INV_X1 u0_u6_u5_U56 (.A( u0_u6_u5_n126 ) , .ZN( u0_u6_u5_n173 ) );
  AND2_X1 u0_u6_u5_U57 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n147 ) );
  AND2_X1 u0_u6_u5_U58 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n148 ) );
  NAND2_X1 u0_u6_u5_U59 (.A1( u0_u6_u5_n105 ) , .A2( u0_u6_u5_n106 ) , .ZN( u0_u6_u5_n158 ) );
  INV_X1 u0_u6_u5_U6 (.A( u0_u6_u5_n135 ) , .ZN( u0_u6_u5_n178 ) );
  NAND2_X1 u0_u6_u5_U60 (.A2( u0_u6_u5_n108 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n139 ) );
  NAND2_X1 u0_u6_u5_U61 (.A1( u0_u6_u5_n106 ) , .A2( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n119 ) );
  NAND2_X1 u0_u6_u5_U62 (.A2( u0_u6_u5_n103 ) , .A1( u0_u6_u5_n105 ) , .ZN( u0_u6_u5_n140 ) );
  NAND2_X1 u0_u6_u5_U63 (.A2( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n105 ) , .ZN( u0_u6_u5_n155 ) );
  NAND2_X1 u0_u6_u5_U64 (.A2( u0_u6_u5_n106 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n122 ) );
  NAND2_X1 u0_u6_u5_U65 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n106 ) , .ZN( u0_u6_u5_n115 ) );
  NAND2_X1 u0_u6_u5_U66 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n103 ) , .ZN( u0_u6_u5_n161 ) );
  NAND2_X1 u0_u6_u5_U67 (.A1( u0_u6_u5_n105 ) , .A2( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n154 ) );
  INV_X1 u0_u6_u5_U68 (.A( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n172 ) );
  NAND2_X1 u0_u6_u5_U69 (.A1( u0_u6_u5_n103 ) , .A2( u0_u6_u5_n108 ) , .ZN( u0_u6_u5_n123 ) );
  OAI22_X1 u0_u6_u5_U7 (.B2( u0_u6_u5_n149 ) , .B1( u0_u6_u5_n150 ) , .A2( u0_u6_u5_n151 ) , .A1( u0_u6_u5_n152 ) , .ZN( u0_u6_u5_n165 ) );
  NAND2_X1 u0_u6_u5_U70 (.A2( u0_u6_u5_n103 ) , .A1( u0_u6_u5_n107 ) , .ZN( u0_u6_u5_n151 ) );
  NAND2_X1 u0_u6_u5_U71 (.A2( u0_u6_u5_n107 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n120 ) );
  NAND2_X1 u0_u6_u5_U72 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n109 ) , .ZN( u0_u6_u5_n157 ) );
  AND2_X1 u0_u6_u5_U73 (.A2( u0_u6_u5_n100 ) , .A1( u0_u6_u5_n104 ) , .ZN( u0_u6_u5_n131 ) );
  INV_X1 u0_u6_u5_U74 (.A( u0_u6_u5_n102 ) , .ZN( u0_u6_u5_n195 ) );
  OAI221_X1 u0_u6_u5_U75 (.A( u0_u6_u5_n101 ) , .ZN( u0_u6_u5_n102 ) , .C2( u0_u6_u5_n115 ) , .C1( u0_u6_u5_n126 ) , .B1( u0_u6_u5_n134 ) , .B2( u0_u6_u5_n160 ) );
  OAI21_X1 u0_u6_u5_U76 (.ZN( u0_u6_u5_n101 ) , .B1( u0_u6_u5_n137 ) , .A( u0_u6_u5_n146 ) , .B2( u0_u6_u5_n147 ) );
  NOR2_X1 u0_u6_u5_U77 (.A2( u0_u6_X_34 ) , .A1( u0_u6_X_35 ) , .ZN( u0_u6_u5_n145 ) );
  NOR2_X1 u0_u6_u5_U78 (.A2( u0_u6_X_34 ) , .ZN( u0_u6_u5_n146 ) , .A1( u0_u6_u5_n171 ) );
  NOR2_X1 u0_u6_u5_U79 (.A2( u0_u6_X_31 ) , .A1( u0_u6_X_32 ) , .ZN( u0_u6_u5_n103 ) );
  NOR3_X1 u0_u6_u5_U8 (.A2( u0_u6_u5_n147 ) , .A1( u0_u6_u5_n148 ) , .ZN( u0_u6_u5_n149 ) , .A3( u0_u6_u5_n194 ) );
  NOR2_X1 u0_u6_u5_U80 (.A2( u0_u6_X_36 ) , .ZN( u0_u6_u5_n105 ) , .A1( u0_u6_u5_n180 ) );
  NOR2_X1 u0_u6_u5_U81 (.A2( u0_u6_X_33 ) , .ZN( u0_u6_u5_n108 ) , .A1( u0_u6_u5_n170 ) );
  NOR2_X1 u0_u6_u5_U82 (.A2( u0_u6_X_33 ) , .A1( u0_u6_X_36 ) , .ZN( u0_u6_u5_n107 ) );
  NOR2_X1 u0_u6_u5_U83 (.A2( u0_u6_X_31 ) , .ZN( u0_u6_u5_n104 ) , .A1( u0_u6_u5_n181 ) );
  NAND2_X1 u0_u6_u5_U84 (.A2( u0_u6_X_34 ) , .A1( u0_u6_X_35 ) , .ZN( u0_u6_u5_n153 ) );
  NAND2_X1 u0_u6_u5_U85 (.A1( u0_u6_X_34 ) , .ZN( u0_u6_u5_n126 ) , .A2( u0_u6_u5_n171 ) );
  AND2_X1 u0_u6_u5_U86 (.A1( u0_u6_X_31 ) , .A2( u0_u6_X_32 ) , .ZN( u0_u6_u5_n106 ) );
  AND2_X1 u0_u6_u5_U87 (.A1( u0_u6_X_31 ) , .ZN( u0_u6_u5_n109 ) , .A2( u0_u6_u5_n181 ) );
  INV_X1 u0_u6_u5_U88 (.A( u0_u6_X_33 ) , .ZN( u0_u6_u5_n180 ) );
  INV_X1 u0_u6_u5_U89 (.A( u0_u6_X_35 ) , .ZN( u0_u6_u5_n171 ) );
  NOR2_X1 u0_u6_u5_U9 (.ZN( u0_u6_u5_n135 ) , .A1( u0_u6_u5_n173 ) , .A2( u0_u6_u5_n176 ) );
  INV_X1 u0_u6_u5_U90 (.A( u0_u6_X_36 ) , .ZN( u0_u6_u5_n170 ) );
  INV_X1 u0_u6_u5_U91 (.A( u0_u6_X_32 ) , .ZN( u0_u6_u5_n181 ) );
  NAND4_X1 u0_u6_u5_U92 (.ZN( u0_out6_29 ) , .A4( u0_u6_u5_n129 ) , .A3( u0_u6_u5_n130 ) , .A2( u0_u6_u5_n168 ) , .A1( u0_u6_u5_n196 ) );
  AOI221_X1 u0_u6_u5_U93 (.A( u0_u6_u5_n128 ) , .ZN( u0_u6_u5_n129 ) , .C2( u0_u6_u5_n132 ) , .B2( u0_u6_u5_n159 ) , .B1( u0_u6_u5_n176 ) , .C1( u0_u6_u5_n184 ) );
  AOI222_X1 u0_u6_u5_U94 (.ZN( u0_u6_u5_n130 ) , .A2( u0_u6_u5_n146 ) , .B1( u0_u6_u5_n147 ) , .C2( u0_u6_u5_n175 ) , .B2( u0_u6_u5_n179 ) , .A1( u0_u6_u5_n188 ) , .C1( u0_u6_u5_n194 ) );
  NAND4_X1 u0_u6_u5_U95 (.ZN( u0_out6_19 ) , .A4( u0_u6_u5_n166 ) , .A3( u0_u6_u5_n167 ) , .A2( u0_u6_u5_n168 ) , .A1( u0_u6_u5_n169 ) );
  AOI22_X1 u0_u6_u5_U96 (.B2( u0_u6_u5_n145 ) , .A2( u0_u6_u5_n146 ) , .ZN( u0_u6_u5_n167 ) , .B1( u0_u6_u5_n182 ) , .A1( u0_u6_u5_n189 ) );
  NOR4_X1 u0_u6_u5_U97 (.A4( u0_u6_u5_n162 ) , .A3( u0_u6_u5_n163 ) , .A2( u0_u6_u5_n164 ) , .A1( u0_u6_u5_n165 ) , .ZN( u0_u6_u5_n166 ) );
  NAND4_X1 u0_u6_u5_U98 (.ZN( u0_out6_11 ) , .A4( u0_u6_u5_n143 ) , .A3( u0_u6_u5_n144 ) , .A2( u0_u6_u5_n169 ) , .A1( u0_u6_u5_n196 ) );
  AOI22_X1 u0_u6_u5_U99 (.A2( u0_u6_u5_n132 ) , .ZN( u0_u6_u5_n144 ) , .B2( u0_u6_u5_n145 ) , .B1( u0_u6_u5_n184 ) , .A1( u0_u6_u5_n194 ) );
  AOI21_X1 u0_u6_u6_U10 (.ZN( u0_u6_u6_n106 ) , .A( u0_u6_u6_n142 ) , .B2( u0_u6_u6_n159 ) , .B1( u0_u6_u6_n164 ) );
  INV_X1 u0_u6_u6_U11 (.A( u0_u6_u6_n155 ) , .ZN( u0_u6_u6_n161 ) );
  INV_X1 u0_u6_u6_U12 (.A( u0_u6_u6_n128 ) , .ZN( u0_u6_u6_n164 ) );
  NAND2_X1 u0_u6_u6_U13 (.ZN( u0_u6_u6_n110 ) , .A1( u0_u6_u6_n122 ) , .A2( u0_u6_u6_n129 ) );
  NAND2_X1 u0_u6_u6_U14 (.ZN( u0_u6_u6_n124 ) , .A2( u0_u6_u6_n146 ) , .A1( u0_u6_u6_n148 ) );
  INV_X1 u0_u6_u6_U15 (.A( u0_u6_u6_n132 ) , .ZN( u0_u6_u6_n171 ) );
  AND2_X1 u0_u6_u6_U16 (.A1( u0_u6_u6_n100 ) , .ZN( u0_u6_u6_n130 ) , .A2( u0_u6_u6_n147 ) );
  INV_X1 u0_u6_u6_U17 (.A( u0_u6_u6_n127 ) , .ZN( u0_u6_u6_n173 ) );
  INV_X1 u0_u6_u6_U18 (.A( u0_u6_u6_n121 ) , .ZN( u0_u6_u6_n167 ) );
  INV_X1 u0_u6_u6_U19 (.A( u0_u6_u6_n100 ) , .ZN( u0_u6_u6_n169 ) );
  INV_X1 u0_u6_u6_U20 (.A( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n170 ) );
  INV_X1 u0_u6_u6_U21 (.A( u0_u6_u6_n113 ) , .ZN( u0_u6_u6_n168 ) );
  AND2_X1 u0_u6_u6_U22 (.A1( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n119 ) , .ZN( u0_u6_u6_n133 ) );
  AND2_X1 u0_u6_u6_U23 (.A2( u0_u6_u6_n121 ) , .A1( u0_u6_u6_n122 ) , .ZN( u0_u6_u6_n131 ) );
  AND3_X1 u0_u6_u6_U24 (.ZN( u0_u6_u6_n120 ) , .A2( u0_u6_u6_n127 ) , .A1( u0_u6_u6_n132 ) , .A3( u0_u6_u6_n145 ) );
  INV_X1 u0_u6_u6_U25 (.A( u0_u6_u6_n146 ) , .ZN( u0_u6_u6_n163 ) );
  AOI222_X1 u0_u6_u6_U26 (.ZN( u0_u6_u6_n114 ) , .A1( u0_u6_u6_n118 ) , .A2( u0_u6_u6_n126 ) , .B2( u0_u6_u6_n151 ) , .C2( u0_u6_u6_n159 ) , .C1( u0_u6_u6_n168 ) , .B1( u0_u6_u6_n169 ) );
  NOR2_X1 u0_u6_u6_U27 (.A1( u0_u6_u6_n162 ) , .A2( u0_u6_u6_n165 ) , .ZN( u0_u6_u6_n98 ) );
  AOI211_X1 u0_u6_u6_U28 (.B( u0_u6_u6_n149 ) , .A( u0_u6_u6_n150 ) , .C2( u0_u6_u6_n151 ) , .C1( u0_u6_u6_n152 ) , .ZN( u0_u6_u6_n153 ) );
  AOI21_X1 u0_u6_u6_U29 (.B2( u0_u6_u6_n147 ) , .B1( u0_u6_u6_n148 ) , .ZN( u0_u6_u6_n149 ) , .A( u0_u6_u6_n158 ) );
  INV_X1 u0_u6_u6_U3 (.A( u0_u6_u6_n110 ) , .ZN( u0_u6_u6_n166 ) );
  AOI21_X1 u0_u6_u6_U30 (.A( u0_u6_u6_n144 ) , .B2( u0_u6_u6_n145 ) , .B1( u0_u6_u6_n146 ) , .ZN( u0_u6_u6_n150 ) );
  NAND2_X1 u0_u6_u6_U31 (.A2( u0_u6_u6_n143 ) , .ZN( u0_u6_u6_n152 ) , .A1( u0_u6_u6_n166 ) );
  NAND2_X1 u0_u6_u6_U32 (.A1( u0_u6_u6_n144 ) , .ZN( u0_u6_u6_n151 ) , .A2( u0_u6_u6_n158 ) );
  NAND2_X1 u0_u6_u6_U33 (.ZN( u0_u6_u6_n132 ) , .A1( u0_u6_u6_n91 ) , .A2( u0_u6_u6_n97 ) );
  AOI22_X1 u0_u6_u6_U34 (.B2( u0_u6_u6_n110 ) , .B1( u0_u6_u6_n111 ) , .A1( u0_u6_u6_n112 ) , .ZN( u0_u6_u6_n115 ) , .A2( u0_u6_u6_n161 ) );
  NAND4_X1 u0_u6_u6_U35 (.A3( u0_u6_u6_n109 ) , .ZN( u0_u6_u6_n112 ) , .A4( u0_u6_u6_n132 ) , .A2( u0_u6_u6_n147 ) , .A1( u0_u6_u6_n166 ) );
  NOR2_X1 u0_u6_u6_U36 (.ZN( u0_u6_u6_n109 ) , .A1( u0_u6_u6_n170 ) , .A2( u0_u6_u6_n173 ) );
  NOR2_X1 u0_u6_u6_U37 (.A2( u0_u6_u6_n126 ) , .ZN( u0_u6_u6_n155 ) , .A1( u0_u6_u6_n160 ) );
  NAND2_X1 u0_u6_u6_U38 (.ZN( u0_u6_u6_n146 ) , .A2( u0_u6_u6_n94 ) , .A1( u0_u6_u6_n99 ) );
  AOI211_X1 u0_u6_u6_U39 (.B( u0_u6_u6_n134 ) , .A( u0_u6_u6_n135 ) , .C1( u0_u6_u6_n136 ) , .ZN( u0_u6_u6_n137 ) , .C2( u0_u6_u6_n151 ) );
  AOI22_X1 u0_u6_u6_U4 (.B2( u0_u6_u6_n101 ) , .A1( u0_u6_u6_n102 ) , .ZN( u0_u6_u6_n103 ) , .B1( u0_u6_u6_n160 ) , .A2( u0_u6_u6_n161 ) );
  NAND4_X1 u0_u6_u6_U40 (.A4( u0_u6_u6_n127 ) , .A3( u0_u6_u6_n128 ) , .A2( u0_u6_u6_n129 ) , .A1( u0_u6_u6_n130 ) , .ZN( u0_u6_u6_n136 ) );
  AOI21_X1 u0_u6_u6_U41 (.B2( u0_u6_u6_n132 ) , .B1( u0_u6_u6_n133 ) , .ZN( u0_u6_u6_n134 ) , .A( u0_u6_u6_n158 ) );
  AOI21_X1 u0_u6_u6_U42 (.B1( u0_u6_u6_n131 ) , .ZN( u0_u6_u6_n135 ) , .A( u0_u6_u6_n144 ) , .B2( u0_u6_u6_n146 ) );
  INV_X1 u0_u6_u6_U43 (.A( u0_u6_u6_n111 ) , .ZN( u0_u6_u6_n158 ) );
  NAND2_X1 u0_u6_u6_U44 (.ZN( u0_u6_u6_n127 ) , .A1( u0_u6_u6_n91 ) , .A2( u0_u6_u6_n92 ) );
  NAND2_X1 u0_u6_u6_U45 (.ZN( u0_u6_u6_n129 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n96 ) );
  INV_X1 u0_u6_u6_U46 (.A( u0_u6_u6_n144 ) , .ZN( u0_u6_u6_n159 ) );
  NAND2_X1 u0_u6_u6_U47 (.ZN( u0_u6_u6_n145 ) , .A2( u0_u6_u6_n97 ) , .A1( u0_u6_u6_n98 ) );
  NAND2_X1 u0_u6_u6_U48 (.ZN( u0_u6_u6_n148 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n94 ) );
  NAND2_X1 u0_u6_u6_U49 (.ZN( u0_u6_u6_n108 ) , .A2( u0_u6_u6_n139 ) , .A1( u0_u6_u6_n144 ) );
  NOR2_X1 u0_u6_u6_U5 (.A1( u0_u6_u6_n118 ) , .ZN( u0_u6_u6_n143 ) , .A2( u0_u6_u6_n168 ) );
  NAND2_X1 u0_u6_u6_U50 (.ZN( u0_u6_u6_n121 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n97 ) );
  NAND2_X1 u0_u6_u6_U51 (.ZN( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n95 ) );
  AND2_X1 u0_u6_u6_U52 (.ZN( u0_u6_u6_n118 ) , .A2( u0_u6_u6_n91 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U53 (.ZN( u0_u6_u6_n147 ) , .A2( u0_u6_u6_n98 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U54 (.ZN( u0_u6_u6_n128 ) , .A1( u0_u6_u6_n94 ) , .A2( u0_u6_u6_n96 ) );
  NAND2_X1 u0_u6_u6_U55 (.ZN( u0_u6_u6_n119 ) , .A2( u0_u6_u6_n95 ) , .A1( u0_u6_u6_n99 ) );
  NAND2_X1 u0_u6_u6_U56 (.ZN( u0_u6_u6_n123 ) , .A2( u0_u6_u6_n91 ) , .A1( u0_u6_u6_n96 ) );
  NAND2_X1 u0_u6_u6_U57 (.ZN( u0_u6_u6_n100 ) , .A2( u0_u6_u6_n92 ) , .A1( u0_u6_u6_n98 ) );
  NAND2_X1 u0_u6_u6_U58 (.ZN( u0_u6_u6_n122 ) , .A1( u0_u6_u6_n94 ) , .A2( u0_u6_u6_n97 ) );
  INV_X1 u0_u6_u6_U59 (.A( u0_u6_u6_n139 ) , .ZN( u0_u6_u6_n160 ) );
  AOI21_X1 u0_u6_u6_U6 (.B1( u0_u6_u6_n107 ) , .B2( u0_u6_u6_n132 ) , .A( u0_u6_u6_n158 ) , .ZN( u0_u6_u6_n88 ) );
  NAND2_X1 u0_u6_u6_U60 (.ZN( u0_u6_u6_n113 ) , .A1( u0_u6_u6_n96 ) , .A2( u0_u6_u6_n98 ) );
  NOR2_X1 u0_u6_u6_U61 (.A2( u0_u6_X_40 ) , .A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n126 ) );
  NOR2_X1 u0_u6_u6_U62 (.A2( u0_u6_X_39 ) , .A1( u0_u6_X_42 ) , .ZN( u0_u6_u6_n92 ) );
  NOR2_X1 u0_u6_u6_U63 (.A2( u0_u6_X_39 ) , .A1( u0_u6_u6_n156 ) , .ZN( u0_u6_u6_n97 ) );
  NOR2_X1 u0_u6_u6_U64 (.A2( u0_u6_X_38 ) , .A1( u0_u6_u6_n165 ) , .ZN( u0_u6_u6_n95 ) );
  NOR2_X1 u0_u6_u6_U65 (.A2( u0_u6_X_41 ) , .ZN( u0_u6_u6_n111 ) , .A1( u0_u6_u6_n157 ) );
  NOR2_X1 u0_u6_u6_U66 (.A2( u0_u6_X_37 ) , .A1( u0_u6_u6_n162 ) , .ZN( u0_u6_u6_n94 ) );
  NOR2_X1 u0_u6_u6_U67 (.A2( u0_u6_X_37 ) , .A1( u0_u6_X_38 ) , .ZN( u0_u6_u6_n91 ) );
  NAND2_X1 u0_u6_u6_U68 (.A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n144 ) , .A2( u0_u6_u6_n157 ) );
  NAND2_X1 u0_u6_u6_U69 (.A2( u0_u6_X_40 ) , .A1( u0_u6_X_41 ) , .ZN( u0_u6_u6_n139 ) );
  OAI21_X1 u0_u6_u6_U7 (.A( u0_u6_u6_n159 ) , .B1( u0_u6_u6_n169 ) , .B2( u0_u6_u6_n173 ) , .ZN( u0_u6_u6_n90 ) );
  AND2_X1 u0_u6_u6_U70 (.A1( u0_u6_X_39 ) , .A2( u0_u6_u6_n156 ) , .ZN( u0_u6_u6_n96 ) );
  AND2_X1 u0_u6_u6_U71 (.A1( u0_u6_X_39 ) , .A2( u0_u6_X_42 ) , .ZN( u0_u6_u6_n99 ) );
  INV_X1 u0_u6_u6_U72 (.A( u0_u6_X_40 ) , .ZN( u0_u6_u6_n157 ) );
  INV_X1 u0_u6_u6_U73 (.A( u0_u6_X_37 ) , .ZN( u0_u6_u6_n165 ) );
  INV_X1 u0_u6_u6_U74 (.A( u0_u6_X_38 ) , .ZN( u0_u6_u6_n162 ) );
  INV_X1 u0_u6_u6_U75 (.A( u0_u6_X_42 ) , .ZN( u0_u6_u6_n156 ) );
  NAND4_X1 u0_u6_u6_U76 (.ZN( u0_out6_32 ) , .A4( u0_u6_u6_n103 ) , .A3( u0_u6_u6_n104 ) , .A2( u0_u6_u6_n105 ) , .A1( u0_u6_u6_n106 ) );
  AOI22_X1 u0_u6_u6_U77 (.ZN( u0_u6_u6_n104 ) , .A1( u0_u6_u6_n111 ) , .B1( u0_u6_u6_n124 ) , .B2( u0_u6_u6_n151 ) , .A2( u0_u6_u6_n93 ) );
  AOI22_X1 u0_u6_u6_U78 (.ZN( u0_u6_u6_n105 ) , .A2( u0_u6_u6_n108 ) , .A1( u0_u6_u6_n118 ) , .B2( u0_u6_u6_n126 ) , .B1( u0_u6_u6_n171 ) );
  NAND4_X1 u0_u6_u6_U79 (.ZN( u0_out6_12 ) , .A4( u0_u6_u6_n114 ) , .A3( u0_u6_u6_n115 ) , .A2( u0_u6_u6_n116 ) , .A1( u0_u6_u6_n117 ) );
  INV_X1 u0_u6_u6_U8 (.ZN( u0_u6_u6_n172 ) , .A( u0_u6_u6_n88 ) );
  OAI22_X1 u0_u6_u6_U80 (.B2( u0_u6_u6_n111 ) , .ZN( u0_u6_u6_n116 ) , .B1( u0_u6_u6_n126 ) , .A2( u0_u6_u6_n164 ) , .A1( u0_u6_u6_n167 ) );
  OAI21_X1 u0_u6_u6_U81 (.A( u0_u6_u6_n108 ) , .ZN( u0_u6_u6_n117 ) , .B2( u0_u6_u6_n141 ) , .B1( u0_u6_u6_n163 ) );
  OAI211_X1 u0_u6_u6_U82 (.ZN( u0_out6_22 ) , .B( u0_u6_u6_n137 ) , .A( u0_u6_u6_n138 ) , .C2( u0_u6_u6_n139 ) , .C1( u0_u6_u6_n140 ) );
  AOI22_X1 u0_u6_u6_U83 (.B1( u0_u6_u6_n124 ) , .A2( u0_u6_u6_n125 ) , .A1( u0_u6_u6_n126 ) , .ZN( u0_u6_u6_n138 ) , .B2( u0_u6_u6_n161 ) );
  AND4_X1 u0_u6_u6_U84 (.A3( u0_u6_u6_n119 ) , .A1( u0_u6_u6_n120 ) , .A4( u0_u6_u6_n129 ) , .ZN( u0_u6_u6_n140 ) , .A2( u0_u6_u6_n143 ) );
  OAI211_X1 u0_u6_u6_U85 (.ZN( u0_out6_7 ) , .B( u0_u6_u6_n153 ) , .C2( u0_u6_u6_n154 ) , .C1( u0_u6_u6_n155 ) , .A( u0_u6_u6_n174 ) );
  NOR3_X1 u0_u6_u6_U86 (.A1( u0_u6_u6_n141 ) , .ZN( u0_u6_u6_n154 ) , .A3( u0_u6_u6_n164 ) , .A2( u0_u6_u6_n171 ) );
  INV_X1 u0_u6_u6_U87 (.A( u0_u6_u6_n142 ) , .ZN( u0_u6_u6_n174 ) );
  NAND3_X1 u0_u6_u6_U88 (.A2( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n125 ) , .A1( u0_u6_u6_n130 ) , .A3( u0_u6_u6_n131 ) );
  NAND3_X1 u0_u6_u6_U89 (.A3( u0_u6_u6_n133 ) , .ZN( u0_u6_u6_n141 ) , .A1( u0_u6_u6_n145 ) , .A2( u0_u6_u6_n148 ) );
  AOI22_X1 u0_u6_u6_U9 (.A2( u0_u6_u6_n151 ) , .B2( u0_u6_u6_n161 ) , .A1( u0_u6_u6_n167 ) , .B1( u0_u6_u6_n170 ) , .ZN( u0_u6_u6_n89 ) );
  NAND3_X1 u0_u6_u6_U90 (.ZN( u0_u6_u6_n101 ) , .A3( u0_u6_u6_n107 ) , .A2( u0_u6_u6_n121 ) , .A1( u0_u6_u6_n127 ) );
  NAND3_X1 u0_u6_u6_U91 (.ZN( u0_u6_u6_n102 ) , .A3( u0_u6_u6_n130 ) , .A2( u0_u6_u6_n145 ) , .A1( u0_u6_u6_n166 ) );
  NAND3_X1 u0_u6_u6_U92 (.A3( u0_u6_u6_n113 ) , .A1( u0_u6_u6_n119 ) , .A2( u0_u6_u6_n123 ) , .ZN( u0_u6_u6_n93 ) );
  NAND3_X1 u0_u6_u6_U93 (.ZN( u0_u6_u6_n142 ) , .A2( u0_u6_u6_n172 ) , .A3( u0_u6_u6_n89 ) , .A1( u0_u6_u6_n90 ) );
  AND3_X1 u0_u6_u7_U10 (.A3( u0_u6_u7_n110 ) , .A2( u0_u6_u7_n127 ) , .A1( u0_u6_u7_n132 ) , .ZN( u0_u6_u7_n92 ) );
  OAI21_X1 u0_u6_u7_U11 (.A( u0_u6_u7_n161 ) , .B1( u0_u6_u7_n168 ) , .B2( u0_u6_u7_n173 ) , .ZN( u0_u6_u7_n91 ) );
  AOI211_X1 u0_u6_u7_U12 (.A( u0_u6_u7_n117 ) , .ZN( u0_u6_u7_n118 ) , .C2( u0_u6_u7_n126 ) , .C1( u0_u6_u7_n177 ) , .B( u0_u6_u7_n180 ) );
  OAI22_X1 u0_u6_u7_U13 (.B1( u0_u6_u7_n115 ) , .ZN( u0_u6_u7_n117 ) , .A2( u0_u6_u7_n133 ) , .A1( u0_u6_u7_n137 ) , .B2( u0_u6_u7_n162 ) );
  INV_X1 u0_u6_u7_U14 (.A( u0_u6_u7_n116 ) , .ZN( u0_u6_u7_n180 ) );
  NOR3_X1 u0_u6_u7_U15 (.ZN( u0_u6_u7_n115 ) , .A3( u0_u6_u7_n145 ) , .A2( u0_u6_u7_n168 ) , .A1( u0_u6_u7_n169 ) );
  OAI211_X1 u0_u6_u7_U16 (.B( u0_u6_u7_n122 ) , .A( u0_u6_u7_n123 ) , .C2( u0_u6_u7_n124 ) , .ZN( u0_u6_u7_n154 ) , .C1( u0_u6_u7_n162 ) );
  AOI222_X1 u0_u6_u7_U17 (.ZN( u0_u6_u7_n122 ) , .C2( u0_u6_u7_n126 ) , .C1( u0_u6_u7_n145 ) , .B1( u0_u6_u7_n161 ) , .A2( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n170 ) , .A1( u0_u6_u7_n176 ) );
  INV_X1 u0_u6_u7_U18 (.A( u0_u6_u7_n133 ) , .ZN( u0_u6_u7_n176 ) );
  NOR3_X1 u0_u6_u7_U19 (.A2( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n135 ) , .ZN( u0_u6_u7_n136 ) , .A3( u0_u6_u7_n171 ) );
  NOR2_X1 u0_u6_u7_U20 (.A1( u0_u6_u7_n130 ) , .A2( u0_u6_u7_n134 ) , .ZN( u0_u6_u7_n153 ) );
  INV_X1 u0_u6_u7_U21 (.A( u0_u6_u7_n101 ) , .ZN( u0_u6_u7_n165 ) );
  NOR2_X1 u0_u6_u7_U22 (.ZN( u0_u6_u7_n111 ) , .A2( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n169 ) );
  AOI21_X1 u0_u6_u7_U23 (.ZN( u0_u6_u7_n104 ) , .B2( u0_u6_u7_n112 ) , .B1( u0_u6_u7_n127 ) , .A( u0_u6_u7_n164 ) );
  AOI21_X1 u0_u6_u7_U24 (.ZN( u0_u6_u7_n106 ) , .B1( u0_u6_u7_n133 ) , .B2( u0_u6_u7_n146 ) , .A( u0_u6_u7_n162 ) );
  AOI21_X1 u0_u6_u7_U25 (.A( u0_u6_u7_n101 ) , .ZN( u0_u6_u7_n107 ) , .B2( u0_u6_u7_n128 ) , .B1( u0_u6_u7_n175 ) );
  INV_X1 u0_u6_u7_U26 (.A( u0_u6_u7_n138 ) , .ZN( u0_u6_u7_n171 ) );
  INV_X1 u0_u6_u7_U27 (.A( u0_u6_u7_n131 ) , .ZN( u0_u6_u7_n177 ) );
  INV_X1 u0_u6_u7_U28 (.A( u0_u6_u7_n110 ) , .ZN( u0_u6_u7_n174 ) );
  NAND2_X1 u0_u6_u7_U29 (.A1( u0_u6_u7_n129 ) , .A2( u0_u6_u7_n132 ) , .ZN( u0_u6_u7_n149 ) );
  OAI21_X1 u0_u6_u7_U3 (.ZN( u0_u6_u7_n159 ) , .A( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n171 ) , .B1( u0_u6_u7_n174 ) );
  NAND2_X1 u0_u6_u7_U30 (.A1( u0_u6_u7_n113 ) , .A2( u0_u6_u7_n124 ) , .ZN( u0_u6_u7_n130 ) );
  INV_X1 u0_u6_u7_U31 (.A( u0_u6_u7_n112 ) , .ZN( u0_u6_u7_n173 ) );
  INV_X1 u0_u6_u7_U32 (.A( u0_u6_u7_n128 ) , .ZN( u0_u6_u7_n168 ) );
  INV_X1 u0_u6_u7_U33 (.A( u0_u6_u7_n148 ) , .ZN( u0_u6_u7_n169 ) );
  INV_X1 u0_u6_u7_U34 (.A( u0_u6_u7_n127 ) , .ZN( u0_u6_u7_n179 ) );
  NOR2_X1 u0_u6_u7_U35 (.ZN( u0_u6_u7_n101 ) , .A2( u0_u6_u7_n150 ) , .A1( u0_u6_u7_n156 ) );
  AOI211_X1 u0_u6_u7_U36 (.B( u0_u6_u7_n154 ) , .A( u0_u6_u7_n155 ) , .C1( u0_u6_u7_n156 ) , .ZN( u0_u6_u7_n157 ) , .C2( u0_u6_u7_n172 ) );
  INV_X1 u0_u6_u7_U37 (.A( u0_u6_u7_n153 ) , .ZN( u0_u6_u7_n172 ) );
  AOI211_X1 u0_u6_u7_U38 (.B( u0_u6_u7_n139 ) , .A( u0_u6_u7_n140 ) , .C2( u0_u6_u7_n141 ) , .ZN( u0_u6_u7_n142 ) , .C1( u0_u6_u7_n156 ) );
  NAND4_X1 u0_u6_u7_U39 (.A3( u0_u6_u7_n127 ) , .A2( u0_u6_u7_n128 ) , .A1( u0_u6_u7_n129 ) , .ZN( u0_u6_u7_n141 ) , .A4( u0_u6_u7_n147 ) );
  INV_X1 u0_u6_u7_U4 (.A( u0_u6_u7_n111 ) , .ZN( u0_u6_u7_n170 ) );
  AOI21_X1 u0_u6_u7_U40 (.A( u0_u6_u7_n137 ) , .B1( u0_u6_u7_n138 ) , .ZN( u0_u6_u7_n139 ) , .B2( u0_u6_u7_n146 ) );
  OAI22_X1 u0_u6_u7_U41 (.B1( u0_u6_u7_n136 ) , .ZN( u0_u6_u7_n140 ) , .A1( u0_u6_u7_n153 ) , .B2( u0_u6_u7_n162 ) , .A2( u0_u6_u7_n164 ) );
  AOI21_X1 u0_u6_u7_U42 (.ZN( u0_u6_u7_n123 ) , .B1( u0_u6_u7_n165 ) , .B2( u0_u6_u7_n177 ) , .A( u0_u6_u7_n97 ) );
  AOI21_X1 u0_u6_u7_U43 (.B2( u0_u6_u7_n113 ) , .B1( u0_u6_u7_n124 ) , .A( u0_u6_u7_n125 ) , .ZN( u0_u6_u7_n97 ) );
  INV_X1 u0_u6_u7_U44 (.A( u0_u6_u7_n125 ) , .ZN( u0_u6_u7_n161 ) );
  INV_X1 u0_u6_u7_U45 (.A( u0_u6_u7_n152 ) , .ZN( u0_u6_u7_n162 ) );
  AOI22_X1 u0_u6_u7_U46 (.A2( u0_u6_u7_n114 ) , .ZN( u0_u6_u7_n119 ) , .B1( u0_u6_u7_n130 ) , .A1( u0_u6_u7_n156 ) , .B2( u0_u6_u7_n165 ) );
  NAND2_X1 u0_u6_u7_U47 (.A2( u0_u6_u7_n112 ) , .ZN( u0_u6_u7_n114 ) , .A1( u0_u6_u7_n175 ) );
  AND2_X1 u0_u6_u7_U48 (.ZN( u0_u6_u7_n145 ) , .A2( u0_u6_u7_n98 ) , .A1( u0_u6_u7_n99 ) );
  NOR2_X1 u0_u6_u7_U49 (.ZN( u0_u6_u7_n137 ) , .A1( u0_u6_u7_n150 ) , .A2( u0_u6_u7_n161 ) );
  INV_X1 u0_u6_u7_U5 (.A( u0_u6_u7_n149 ) , .ZN( u0_u6_u7_n175 ) );
  AOI21_X1 u0_u6_u7_U50 (.ZN( u0_u6_u7_n105 ) , .B2( u0_u6_u7_n110 ) , .A( u0_u6_u7_n125 ) , .B1( u0_u6_u7_n147 ) );
  NAND2_X1 u0_u6_u7_U51 (.ZN( u0_u6_u7_n146 ) , .A1( u0_u6_u7_n95 ) , .A2( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U52 (.A2( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n147 ) , .A1( u0_u6_u7_n93 ) );
  NAND2_X1 u0_u6_u7_U53 (.A1( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n127 ) , .A2( u0_u6_u7_n99 ) );
  OR2_X1 u0_u6_u7_U54 (.ZN( u0_u6_u7_n126 ) , .A2( u0_u6_u7_n152 ) , .A1( u0_u6_u7_n156 ) );
  NAND2_X1 u0_u6_u7_U55 (.A2( u0_u6_u7_n102 ) , .A1( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n133 ) );
  NAND2_X1 u0_u6_u7_U56 (.ZN( u0_u6_u7_n112 ) , .A2( u0_u6_u7_n96 ) , .A1( u0_u6_u7_n99 ) );
  NAND2_X1 u0_u6_u7_U57 (.A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n128 ) , .A1( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U58 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n113 ) , .A2( u0_u6_u7_n93 ) );
  NAND2_X1 u0_u6_u7_U59 (.A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n124 ) , .A1( u0_u6_u7_n96 ) );
  INV_X1 u0_u6_u7_U6 (.A( u0_u6_u7_n154 ) , .ZN( u0_u6_u7_n178 ) );
  NAND2_X1 u0_u6_u7_U60 (.ZN( u0_u6_u7_n110 ) , .A1( u0_u6_u7_n95 ) , .A2( u0_u6_u7_n96 ) );
  INV_X1 u0_u6_u7_U61 (.A( u0_u6_u7_n150 ) , .ZN( u0_u6_u7_n164 ) );
  AND2_X1 u0_u6_u7_U62 (.ZN( u0_u6_u7_n134 ) , .A1( u0_u6_u7_n93 ) , .A2( u0_u6_u7_n98 ) );
  NAND2_X1 u0_u6_u7_U63 (.A1( u0_u6_u7_n100 ) , .A2( u0_u6_u7_n102 ) , .ZN( u0_u6_u7_n129 ) );
  NAND2_X1 u0_u6_u7_U64 (.A2( u0_u6_u7_n103 ) , .ZN( u0_u6_u7_n131 ) , .A1( u0_u6_u7_n95 ) );
  NAND2_X1 u0_u6_u7_U65 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n138 ) , .A2( u0_u6_u7_n99 ) );
  NAND2_X1 u0_u6_u7_U66 (.ZN( u0_u6_u7_n132 ) , .A1( u0_u6_u7_n93 ) , .A2( u0_u6_u7_n96 ) );
  NAND2_X1 u0_u6_u7_U67 (.A1( u0_u6_u7_n100 ) , .ZN( u0_u6_u7_n148 ) , .A2( u0_u6_u7_n95 ) );
  NOR2_X1 u0_u6_u7_U68 (.A2( u0_u6_X_47 ) , .ZN( u0_u6_u7_n150 ) , .A1( u0_u6_u7_n163 ) );
  NOR2_X1 u0_u6_u7_U69 (.A2( u0_u6_X_43 ) , .A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n103 ) );
  AOI211_X1 u0_u6_u7_U7 (.ZN( u0_u6_u7_n116 ) , .A( u0_u6_u7_n155 ) , .C1( u0_u6_u7_n161 ) , .C2( u0_u6_u7_n171 ) , .B( u0_u6_u7_n94 ) );
  NOR2_X1 u0_u6_u7_U70 (.A2( u0_u6_X_48 ) , .A1( u0_u6_u7_n166 ) , .ZN( u0_u6_u7_n95 ) );
  NOR2_X1 u0_u6_u7_U71 (.A2( u0_u6_X_45 ) , .A1( u0_u6_X_48 ) , .ZN( u0_u6_u7_n99 ) );
  NOR2_X1 u0_u6_u7_U72 (.A2( u0_u6_X_44 ) , .A1( u0_u6_u7_n167 ) , .ZN( u0_u6_u7_n98 ) );
  NOR2_X1 u0_u6_u7_U73 (.A2( u0_u6_X_46 ) , .A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n152 ) );
  AND2_X1 u0_u6_u7_U74 (.A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n156 ) , .A2( u0_u6_u7_n163 ) );
  NAND2_X1 u0_u6_u7_U75 (.A2( u0_u6_X_46 ) , .A1( u0_u6_X_47 ) , .ZN( u0_u6_u7_n125 ) );
  AND2_X1 u0_u6_u7_U76 (.A2( u0_u6_X_45 ) , .A1( u0_u6_X_48 ) , .ZN( u0_u6_u7_n102 ) );
  AND2_X1 u0_u6_u7_U77 (.A2( u0_u6_X_43 ) , .A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n96 ) );
  AND2_X1 u0_u6_u7_U78 (.A1( u0_u6_X_44 ) , .ZN( u0_u6_u7_n100 ) , .A2( u0_u6_u7_n167 ) );
  AND2_X1 u0_u6_u7_U79 (.A1( u0_u6_X_48 ) , .A2( u0_u6_u7_n166 ) , .ZN( u0_u6_u7_n93 ) );
  OAI222_X1 u0_u6_u7_U8 (.C2( u0_u6_u7_n101 ) , .B2( u0_u6_u7_n111 ) , .A1( u0_u6_u7_n113 ) , .C1( u0_u6_u7_n146 ) , .A2( u0_u6_u7_n162 ) , .B1( u0_u6_u7_n164 ) , .ZN( u0_u6_u7_n94 ) );
  INV_X1 u0_u6_u7_U80 (.A( u0_u6_X_46 ) , .ZN( u0_u6_u7_n163 ) );
  INV_X1 u0_u6_u7_U81 (.A( u0_u6_X_43 ) , .ZN( u0_u6_u7_n167 ) );
  INV_X1 u0_u6_u7_U82 (.A( u0_u6_X_45 ) , .ZN( u0_u6_u7_n166 ) );
  NAND4_X1 u0_u6_u7_U83 (.ZN( u0_out6_5 ) , .A4( u0_u6_u7_n108 ) , .A3( u0_u6_u7_n109 ) , .A1( u0_u6_u7_n116 ) , .A2( u0_u6_u7_n123 ) );
  AOI22_X1 u0_u6_u7_U84 (.ZN( u0_u6_u7_n109 ) , .A2( u0_u6_u7_n126 ) , .B2( u0_u6_u7_n145 ) , .B1( u0_u6_u7_n156 ) , .A1( u0_u6_u7_n171 ) );
  NOR4_X1 u0_u6_u7_U85 (.A4( u0_u6_u7_n104 ) , .A3( u0_u6_u7_n105 ) , .A2( u0_u6_u7_n106 ) , .A1( u0_u6_u7_n107 ) , .ZN( u0_u6_u7_n108 ) );
  NAND4_X1 u0_u6_u7_U86 (.ZN( u0_out6_27 ) , .A4( u0_u6_u7_n118 ) , .A3( u0_u6_u7_n119 ) , .A2( u0_u6_u7_n120 ) , .A1( u0_u6_u7_n121 ) );
  OAI21_X1 u0_u6_u7_U87 (.ZN( u0_u6_u7_n121 ) , .B2( u0_u6_u7_n145 ) , .A( u0_u6_u7_n150 ) , .B1( u0_u6_u7_n174 ) );
  OAI21_X1 u0_u6_u7_U88 (.ZN( u0_u6_u7_n120 ) , .A( u0_u6_u7_n161 ) , .B2( u0_u6_u7_n170 ) , .B1( u0_u6_u7_n179 ) );
  NAND4_X1 u0_u6_u7_U89 (.ZN( u0_out6_21 ) , .A4( u0_u6_u7_n157 ) , .A3( u0_u6_u7_n158 ) , .A2( u0_u6_u7_n159 ) , .A1( u0_u6_u7_n160 ) );
  OAI221_X1 u0_u6_u7_U9 (.C1( u0_u6_u7_n101 ) , .C2( u0_u6_u7_n147 ) , .ZN( u0_u6_u7_n155 ) , .B2( u0_u6_u7_n162 ) , .A( u0_u6_u7_n91 ) , .B1( u0_u6_u7_n92 ) );
  OAI21_X1 u0_u6_u7_U90 (.B1( u0_u6_u7_n145 ) , .ZN( u0_u6_u7_n160 ) , .A( u0_u6_u7_n161 ) , .B2( u0_u6_u7_n177 ) );
  AOI22_X1 u0_u6_u7_U91 (.B2( u0_u6_u7_n149 ) , .B1( u0_u6_u7_n150 ) , .A2( u0_u6_u7_n151 ) , .A1( u0_u6_u7_n152 ) , .ZN( u0_u6_u7_n158 ) );
  NAND4_X1 u0_u6_u7_U92 (.ZN( u0_out6_15 ) , .A4( u0_u6_u7_n142 ) , .A3( u0_u6_u7_n143 ) , .A2( u0_u6_u7_n144 ) , .A1( u0_u6_u7_n178 ) );
  OR2_X1 u0_u6_u7_U93 (.A2( u0_u6_u7_n125 ) , .A1( u0_u6_u7_n129 ) , .ZN( u0_u6_u7_n144 ) );
  AOI22_X1 u0_u6_u7_U94 (.A2( u0_u6_u7_n126 ) , .ZN( u0_u6_u7_n143 ) , .B2( u0_u6_u7_n165 ) , .B1( u0_u6_u7_n173 ) , .A1( u0_u6_u7_n174 ) );
  NAND3_X1 u0_u6_u7_U95 (.A3( u0_u6_u7_n146 ) , .A2( u0_u6_u7_n147 ) , .A1( u0_u6_u7_n148 ) , .ZN( u0_u6_u7_n151 ) );
  NAND3_X1 u0_u6_u7_U96 (.A3( u0_u6_u7_n131 ) , .A2( u0_u6_u7_n132 ) , .A1( u0_u6_u7_n133 ) , .ZN( u0_u6_u7_n135 ) );
  XOR2_X1 u0_u9_U16 (.B( u0_K10_3 ) , .A( u0_R8_2 ) , .Z( u0_u9_X_3 ) );
  XOR2_X1 u0_u9_U27 (.B( u0_K10_2 ) , .A( u0_R8_1 ) , .Z( u0_u9_X_2 ) );
  XOR2_X1 u0_u9_U38 (.B( u0_K10_1 ) , .A( u0_R8_32 ) , .Z( u0_u9_X_1 ) );
  XOR2_X1 u0_u9_U4 (.B( u0_K10_6 ) , .A( u0_R8_5 ) , .Z( u0_u9_X_6 ) );
  XOR2_X1 u0_u9_U5 (.B( u0_K10_5 ) , .A( u0_R8_4 ) , .Z( u0_u9_X_5 ) );
  XOR2_X1 u0_u9_U6 (.B( u0_K10_4 ) , .A( u0_R8_3 ) , .Z( u0_u9_X_4 ) );
  AND3_X1 u0_u9_u0_U10 (.A2( u0_u9_u0_n112 ) , .ZN( u0_u9_u0_n127 ) , .A3( u0_u9_u0_n130 ) , .A1( u0_u9_u0_n148 ) );
  NAND2_X1 u0_u9_u0_U11 (.ZN( u0_u9_u0_n113 ) , .A1( u0_u9_u0_n139 ) , .A2( u0_u9_u0_n149 ) );
  AND2_X1 u0_u9_u0_U12 (.ZN( u0_u9_u0_n107 ) , .A1( u0_u9_u0_n130 ) , .A2( u0_u9_u0_n140 ) );
  AND2_X1 u0_u9_u0_U13 (.A2( u0_u9_u0_n129 ) , .A1( u0_u9_u0_n130 ) , .ZN( u0_u9_u0_n151 ) );
  AND2_X1 u0_u9_u0_U14 (.A1( u0_u9_u0_n108 ) , .A2( u0_u9_u0_n125 ) , .ZN( u0_u9_u0_n145 ) );
  INV_X1 u0_u9_u0_U15 (.A( u0_u9_u0_n143 ) , .ZN( u0_u9_u0_n173 ) );
  NOR2_X1 u0_u9_u0_U16 (.A2( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n147 ) , .A1( u0_u9_u0_n160 ) );
  AOI21_X1 u0_u9_u0_U17 (.B1( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n132 ) , .A( u0_u9_u0_n165 ) , .B2( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U18 (.A( u0_u9_u0_n142 ) , .ZN( u0_u9_u0_n165 ) );
  OAI221_X1 u0_u9_u0_U19 (.C1( u0_u9_u0_n121 ) , .ZN( u0_u9_u0_n122 ) , .B2( u0_u9_u0_n127 ) , .A( u0_u9_u0_n143 ) , .B1( u0_u9_u0_n144 ) , .C2( u0_u9_u0_n147 ) );
  OAI22_X1 u0_u9_u0_U20 (.B1( u0_u9_u0_n131 ) , .A1( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n147 ) , .A2( u0_u9_u0_n90 ) , .ZN( u0_u9_u0_n91 ) );
  AND3_X1 u0_u9_u0_U21 (.A3( u0_u9_u0_n121 ) , .A2( u0_u9_u0_n125 ) , .A1( u0_u9_u0_n148 ) , .ZN( u0_u9_u0_n90 ) );
  OAI22_X1 u0_u9_u0_U22 (.B1( u0_u9_u0_n125 ) , .ZN( u0_u9_u0_n126 ) , .A1( u0_u9_u0_n138 ) , .A2( u0_u9_u0_n146 ) , .B2( u0_u9_u0_n147 ) );
  NOR2_X1 u0_u9_u0_U23 (.A1( u0_u9_u0_n163 ) , .A2( u0_u9_u0_n164 ) , .ZN( u0_u9_u0_n95 ) );
  INV_X1 u0_u9_u0_U24 (.A( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n161 ) );
  NOR2_X1 u0_u9_u0_U25 (.A1( u0_u9_u0_n120 ) , .ZN( u0_u9_u0_n143 ) , .A2( u0_u9_u0_n167 ) );
  OAI221_X1 u0_u9_u0_U26 (.C1( u0_u9_u0_n112 ) , .ZN( u0_u9_u0_n120 ) , .B1( u0_u9_u0_n138 ) , .B2( u0_u9_u0_n141 ) , .C2( u0_u9_u0_n147 ) , .A( u0_u9_u0_n172 ) );
  AOI211_X1 u0_u9_u0_U27 (.B( u0_u9_u0_n115 ) , .A( u0_u9_u0_n116 ) , .C2( u0_u9_u0_n117 ) , .C1( u0_u9_u0_n118 ) , .ZN( u0_u9_u0_n119 ) );
  NAND2_X1 u0_u9_u0_U28 (.A1( u0_u9_u0_n101 ) , .A2( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n150 ) );
  AOI22_X1 u0_u9_u0_U29 (.B2( u0_u9_u0_n109 ) , .A2( u0_u9_u0_n110 ) , .ZN( u0_u9_u0_n111 ) , .B1( u0_u9_u0_n118 ) , .A1( u0_u9_u0_n160 ) );
  INV_X1 u0_u9_u0_U3 (.A( u0_u9_u0_n113 ) , .ZN( u0_u9_u0_n166 ) );
  INV_X1 u0_u9_u0_U30 (.A( u0_u9_u0_n118 ) , .ZN( u0_u9_u0_n158 ) );
  NAND2_X1 u0_u9_u0_U31 (.A2( u0_u9_u0_n100 ) , .A1( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n139 ) );
  NAND2_X1 u0_u9_u0_U32 (.A2( u0_u9_u0_n100 ) , .ZN( u0_u9_u0_n131 ) , .A1( u0_u9_u0_n92 ) );
  NAND2_X1 u0_u9_u0_U33 (.ZN( u0_u9_u0_n108 ) , .A1( u0_u9_u0_n92 ) , .A2( u0_u9_u0_n94 ) );
  AOI21_X1 u0_u9_u0_U34 (.ZN( u0_u9_u0_n104 ) , .B1( u0_u9_u0_n107 ) , .B2( u0_u9_u0_n141 ) , .A( u0_u9_u0_n144 ) );
  AOI21_X1 u0_u9_u0_U35 (.B1( u0_u9_u0_n127 ) , .B2( u0_u9_u0_n129 ) , .A( u0_u9_u0_n138 ) , .ZN( u0_u9_u0_n96 ) );
  NAND2_X1 u0_u9_u0_U36 (.A2( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n114 ) , .A1( u0_u9_u0_n92 ) );
  AOI21_X1 u0_u9_u0_U37 (.ZN( u0_u9_u0_n116 ) , .B2( u0_u9_u0_n142 ) , .A( u0_u9_u0_n144 ) , .B1( u0_u9_u0_n166 ) );
  NAND2_X1 u0_u9_u0_U38 (.A1( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n130 ) , .A2( u0_u9_u0_n94 ) );
  NAND2_X1 u0_u9_u0_U39 (.A1( u0_u9_u0_n100 ) , .A2( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n125 ) );
  AOI21_X1 u0_u9_u0_U4 (.B1( u0_u9_u0_n114 ) , .ZN( u0_u9_u0_n115 ) , .B2( u0_u9_u0_n129 ) , .A( u0_u9_u0_n161 ) );
  NAND2_X1 u0_u9_u0_U40 (.A2( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n140 ) , .A1( u0_u9_u0_n94 ) );
  INV_X1 u0_u9_u0_U41 (.A( u0_u9_u0_n138 ) , .ZN( u0_u9_u0_n160 ) );
  NAND2_X1 u0_u9_u0_U42 (.A2( u0_u9_u0_n102 ) , .A1( u0_u9_u0_n103 ) , .ZN( u0_u9_u0_n149 ) );
  NAND2_X1 u0_u9_u0_U43 (.A2( u0_u9_u0_n101 ) , .ZN( u0_u9_u0_n121 ) , .A1( u0_u9_u0_n93 ) );
  NAND2_X1 u0_u9_u0_U44 (.ZN( u0_u9_u0_n112 ) , .A2( u0_u9_u0_n92 ) , .A1( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U45 (.ZN( u0_u9_u0_n172 ) , .A( u0_u9_u0_n88 ) );
  OAI222_X1 u0_u9_u0_U46 (.C1( u0_u9_u0_n108 ) , .A1( u0_u9_u0_n125 ) , .B2( u0_u9_u0_n128 ) , .B1( u0_u9_u0_n144 ) , .A2( u0_u9_u0_n158 ) , .C2( u0_u9_u0_n161 ) , .ZN( u0_u9_u0_n88 ) );
  OR3_X1 u0_u9_u0_U47 (.A3( u0_u9_u0_n152 ) , .A2( u0_u9_u0_n153 ) , .A1( u0_u9_u0_n154 ) , .ZN( u0_u9_u0_n155 ) );
  AOI21_X1 u0_u9_u0_U48 (.A( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n145 ) , .B1( u0_u9_u0_n146 ) , .ZN( u0_u9_u0_n154 ) );
  AOI21_X1 u0_u9_u0_U49 (.B2( u0_u9_u0_n150 ) , .B1( u0_u9_u0_n151 ) , .ZN( u0_u9_u0_n152 ) , .A( u0_u9_u0_n158 ) );
  AOI21_X1 u0_u9_u0_U5 (.B2( u0_u9_u0_n131 ) , .ZN( u0_u9_u0_n134 ) , .B1( u0_u9_u0_n151 ) , .A( u0_u9_u0_n158 ) );
  AOI21_X1 u0_u9_u0_U50 (.A( u0_u9_u0_n147 ) , .B2( u0_u9_u0_n148 ) , .B1( u0_u9_u0_n149 ) , .ZN( u0_u9_u0_n153 ) );
  INV_X1 u0_u9_u0_U51 (.ZN( u0_u9_u0_n171 ) , .A( u0_u9_u0_n99 ) );
  OAI211_X1 u0_u9_u0_U52 (.C2( u0_u9_u0_n140 ) , .C1( u0_u9_u0_n161 ) , .A( u0_u9_u0_n169 ) , .B( u0_u9_u0_n98 ) , .ZN( u0_u9_u0_n99 ) );
  INV_X1 u0_u9_u0_U53 (.ZN( u0_u9_u0_n169 ) , .A( u0_u9_u0_n91 ) );
  AOI211_X1 u0_u9_u0_U54 (.C1( u0_u9_u0_n118 ) , .A( u0_u9_u0_n123 ) , .B( u0_u9_u0_n96 ) , .C2( u0_u9_u0_n97 ) , .ZN( u0_u9_u0_n98 ) );
  NOR2_X1 u0_u9_u0_U55 (.A2( u0_u9_X_2 ) , .ZN( u0_u9_u0_n103 ) , .A1( u0_u9_u0_n164 ) );
  NOR2_X1 u0_u9_u0_U56 (.A2( u0_u9_X_4 ) , .A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n118 ) );
  NOR2_X1 u0_u9_u0_U57 (.A2( u0_u9_X_3 ) , .A1( u0_u9_X_6 ) , .ZN( u0_u9_u0_n94 ) );
  NOR2_X1 u0_u9_u0_U58 (.A2( u0_u9_X_6 ) , .ZN( u0_u9_u0_n100 ) , .A1( u0_u9_u0_n162 ) );
  NAND2_X1 u0_u9_u0_U59 (.A2( u0_u9_X_4 ) , .A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n144 ) );
  NOR2_X1 u0_u9_u0_U6 (.A1( u0_u9_u0_n108 ) , .ZN( u0_u9_u0_n123 ) , .A2( u0_u9_u0_n158 ) );
  NOR2_X1 u0_u9_u0_U60 (.A2( u0_u9_X_5 ) , .ZN( u0_u9_u0_n136 ) , .A1( u0_u9_u0_n159 ) );
  NAND2_X1 u0_u9_u0_U61 (.A1( u0_u9_X_5 ) , .ZN( u0_u9_u0_n138 ) , .A2( u0_u9_u0_n159 ) );
  AND2_X1 u0_u9_u0_U62 (.A2( u0_u9_X_3 ) , .A1( u0_u9_X_6 ) , .ZN( u0_u9_u0_n102 ) );
  AND2_X1 u0_u9_u0_U63 (.A1( u0_u9_X_6 ) , .A2( u0_u9_u0_n162 ) , .ZN( u0_u9_u0_n93 ) );
  INV_X1 u0_u9_u0_U64 (.A( u0_u9_X_4 ) , .ZN( u0_u9_u0_n159 ) );
  INV_X1 u0_u9_u0_U65 (.A( u0_u9_X_3 ) , .ZN( u0_u9_u0_n162 ) );
  INV_X1 u0_u9_u0_U66 (.A( u0_u9_X_2 ) , .ZN( u0_u9_u0_n163 ) );
  INV_X1 u0_u9_u0_U67 (.A( u0_u9_u0_n126 ) , .ZN( u0_u9_u0_n168 ) );
  AOI211_X1 u0_u9_u0_U68 (.B( u0_u9_u0_n133 ) , .A( u0_u9_u0_n134 ) , .C2( u0_u9_u0_n135 ) , .C1( u0_u9_u0_n136 ) , .ZN( u0_u9_u0_n137 ) );
  INV_X1 u0_u9_u0_U69 (.ZN( u0_u9_u0_n174 ) , .A( u0_u9_u0_n89 ) );
  OAI21_X1 u0_u9_u0_U7 (.B1( u0_u9_u0_n150 ) , .B2( u0_u9_u0_n158 ) , .A( u0_u9_u0_n172 ) , .ZN( u0_u9_u0_n89 ) );
  AOI211_X1 u0_u9_u0_U70 (.B( u0_u9_u0_n104 ) , .A( u0_u9_u0_n105 ) , .ZN( u0_u9_u0_n106 ) , .C2( u0_u9_u0_n113 ) , .C1( u0_u9_u0_n160 ) );
  OR4_X1 u0_u9_u0_U71 (.ZN( u0_out9_17 ) , .A4( u0_u9_u0_n122 ) , .A2( u0_u9_u0_n123 ) , .A1( u0_u9_u0_n124 ) , .A3( u0_u9_u0_n170 ) );
  AOI21_X1 u0_u9_u0_U72 (.B2( u0_u9_u0_n107 ) , .ZN( u0_u9_u0_n124 ) , .B1( u0_u9_u0_n128 ) , .A( u0_u9_u0_n161 ) );
  INV_X1 u0_u9_u0_U73 (.A( u0_u9_u0_n111 ) , .ZN( u0_u9_u0_n170 ) );
  OR4_X1 u0_u9_u0_U74 (.ZN( u0_out9_31 ) , .A4( u0_u9_u0_n155 ) , .A2( u0_u9_u0_n156 ) , .A1( u0_u9_u0_n157 ) , .A3( u0_u9_u0_n173 ) );
  AOI21_X1 u0_u9_u0_U75 (.A( u0_u9_u0_n138 ) , .B2( u0_u9_u0_n139 ) , .B1( u0_u9_u0_n140 ) , .ZN( u0_u9_u0_n157 ) );
  AOI21_X1 u0_u9_u0_U76 (.B2( u0_u9_u0_n141 ) , .B1( u0_u9_u0_n142 ) , .ZN( u0_u9_u0_n156 ) , .A( u0_u9_u0_n161 ) );
  AOI21_X1 u0_u9_u0_U77 (.B1( u0_u9_u0_n132 ) , .ZN( u0_u9_u0_n133 ) , .A( u0_u9_u0_n144 ) , .B2( u0_u9_u0_n166 ) );
  OAI22_X1 u0_u9_u0_U78 (.ZN( u0_u9_u0_n105 ) , .A2( u0_u9_u0_n132 ) , .B1( u0_u9_u0_n146 ) , .A1( u0_u9_u0_n147 ) , .B2( u0_u9_u0_n161 ) );
  NAND2_X1 u0_u9_u0_U79 (.ZN( u0_u9_u0_n110 ) , .A2( u0_u9_u0_n132 ) , .A1( u0_u9_u0_n145 ) );
  AND2_X1 u0_u9_u0_U8 (.A1( u0_u9_u0_n114 ) , .A2( u0_u9_u0_n121 ) , .ZN( u0_u9_u0_n146 ) );
  INV_X1 u0_u9_u0_U80 (.A( u0_u9_u0_n119 ) , .ZN( u0_u9_u0_n167 ) );
  NAND2_X1 u0_u9_u0_U81 (.ZN( u0_u9_u0_n148 ) , .A1( u0_u9_u0_n93 ) , .A2( u0_u9_u0_n95 ) );
  NAND2_X1 u0_u9_u0_U82 (.A1( u0_u9_u0_n100 ) , .ZN( u0_u9_u0_n129 ) , .A2( u0_u9_u0_n95 ) );
  NAND2_X1 u0_u9_u0_U83 (.A1( u0_u9_u0_n102 ) , .ZN( u0_u9_u0_n128 ) , .A2( u0_u9_u0_n95 ) );
  NOR2_X1 u0_u9_u0_U84 (.A2( u0_u9_X_1 ) , .A1( u0_u9_X_2 ) , .ZN( u0_u9_u0_n92 ) );
  NAND2_X1 u0_u9_u0_U85 (.ZN( u0_u9_u0_n142 ) , .A1( u0_u9_u0_n94 ) , .A2( u0_u9_u0_n95 ) );
  NOR2_X1 u0_u9_u0_U86 (.A2( u0_u9_X_1 ) , .ZN( u0_u9_u0_n101 ) , .A1( u0_u9_u0_n163 ) );
  INV_X1 u0_u9_u0_U87 (.A( u0_u9_X_1 ) , .ZN( u0_u9_u0_n164 ) );
  NAND3_X1 u0_u9_u0_U88 (.ZN( u0_out9_23 ) , .A3( u0_u9_u0_n137 ) , .A1( u0_u9_u0_n168 ) , .A2( u0_u9_u0_n171 ) );
  NAND3_X1 u0_u9_u0_U89 (.A3( u0_u9_u0_n127 ) , .A2( u0_u9_u0_n128 ) , .ZN( u0_u9_u0_n135 ) , .A1( u0_u9_u0_n150 ) );
  AND2_X1 u0_u9_u0_U9 (.A1( u0_u9_u0_n131 ) , .ZN( u0_u9_u0_n141 ) , .A2( u0_u9_u0_n150 ) );
  NAND3_X1 u0_u9_u0_U90 (.ZN( u0_u9_u0_n117 ) , .A3( u0_u9_u0_n132 ) , .A2( u0_u9_u0_n139 ) , .A1( u0_u9_u0_n148 ) );
  NAND3_X1 u0_u9_u0_U91 (.ZN( u0_u9_u0_n109 ) , .A2( u0_u9_u0_n114 ) , .A3( u0_u9_u0_n140 ) , .A1( u0_u9_u0_n149 ) );
  NAND3_X1 u0_u9_u0_U92 (.ZN( u0_out9_9 ) , .A3( u0_u9_u0_n106 ) , .A2( u0_u9_u0_n171 ) , .A1( u0_u9_u0_n174 ) );
  NAND3_X1 u0_u9_u0_U93 (.A2( u0_u9_u0_n128 ) , .A1( u0_u9_u0_n132 ) , .A3( u0_u9_u0_n146 ) , .ZN( u0_u9_u0_n97 ) );
  NAND2_X1 u0_uk_U1005 (.A1( u0_uk_K_r1_10 ) , .A2( u0_uk_n100 ) , .ZN( u0_uk_n841 ) );
  OAI22_X1 u0_uk_U102 (.ZN( u0_K7_5 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n384 ) , .B2( u0_uk_n401 ) );
  OAI21_X1 u0_uk_U1036 (.ZN( u0_K16_28 ) , .B1( u0_uk_n60 ) , .B2( u0_uk_n669 ) , .A( u0_uk_n905 ) );
  NAND2_X1 u0_uk_U1037 (.A1( u0_uk_K_r14_8 ) , .A2( u0_uk_n83 ) , .ZN( u0_uk_n905 ) );
  OAI21_X1 u0_uk_U1040 (.ZN( u0_K7_31 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n380 ) , .A( u0_uk_n772 ) );
  NAND2_X1 u0_uk_U1041 (.A1( u0_uk_K_r5_16 ) , .A2( u0_uk_n102 ) , .ZN( u0_uk_n772 ) );
  OAI21_X1 u0_uk_U1056 (.ZN( u0_K7_38 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n389 ) , .A( u0_uk_n767 ) );
  NAND2_X1 u0_uk_U1057 (.A1( u0_uk_K_r5_8 ) , .A2( u0_uk_n117 ) , .ZN( u0_uk_n767 ) );
  OAI21_X1 u0_uk_U1089 (.ZN( u0_K16_14 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n653 ) , .A( u0_uk_n908 ) );
  NAND2_X1 u0_uk_U1090 (.A1( u0_uk_K_r14_18 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n908 ) );
  INV_X1 u0_uk_U11 (.A( u0_uk_n231 ) , .ZN( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U110 (.ZN( u0_K12_41 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n144 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n153 ) );
  INV_X1 u0_uk_U1101 (.ZN( u0_K2_10 ) , .A( u0_uk_n868 ) );
  AOI22_X1 u0_uk_U1102 (.B2( u0_uk_K_r0_34 ) , .A2( u0_uk_K_r0_55 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n868 ) );
  INV_X1 u0_uk_U1109 (.ZN( u0_K11_8 ) , .A( u0_uk_n982 ) );
  AOI22_X1 u0_uk_U1110 (.B2( u0_uk_K_r9_12 ) , .A2( u0_uk_K_r9_18 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n982 ) );
  INV_X1 u0_uk_U1111 (.ZN( u0_K11_12 ) , .A( u0_uk_n1003 ) );
  AOI22_X1 u0_uk_U1112 (.B2( u0_uk_K_r9_25 ) , .A2( u0_uk_K_r9_6 ) , .ZN( u0_uk_n1003 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n207 ) );
  INV_X1 u0_uk_U1119 (.ZN( u0_K2_7 ) , .A( u0_uk_n855 ) );
  INV_X1 u0_uk_U1127 (.ZN( u0_K7_32 ) , .A( u0_uk_n771 ) );
  AOI22_X1 u0_uk_U1128 (.B2( u0_uk_K_r5_0 ) , .A2( u0_uk_K_r5_51 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n771 ) );
  INV_X1 u0_uk_U1131 (.ZN( u0_K12_42 ) , .A( u0_uk_n966 ) );
  AOI22_X1 u0_uk_U1132 (.B2( u0_uk_K_r10_28 ) , .A2( u0_uk_K_r10_9 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n966 ) );
  INV_X1 u0_uk_U1139 (.ZN( u0_K7_34 ) , .A( u0_uk_n770 ) );
  OAI22_X1 u0_uk_U119 (.ZN( u0_K7_47 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n388 ) , .A2( u0_uk_n402 ) );
  INV_X1 u0_uk_U133 (.ZN( u0_K12_15 ) , .A( u0_uk_n980 ) );
  AOI22_X1 u0_uk_U134 (.B2( u0_uk_K_r10_25 ) , .A2( u0_uk_K_r10_34 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n980 ) );
  INV_X1 u0_uk_U14 (.A( u0_uk_n222 ) , .ZN( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U142 (.ZN( u0_K2_15 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n597 ) , .A( u0_uk_n865 ) );
  NAND2_X1 u0_uk_U143 (.A1( u0_uk_K_r0_19 ) , .A2( u0_uk_n102 ) , .ZN( u0_uk_n865 ) );
  OAI22_X1 u0_uk_U145 (.ZN( u0_K16_15 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n645 ) , .B2( u0_uk_n652 ) );
  INV_X1 u0_uk_U16 (.ZN( u0_uk_n110 ) , .A( u0_uk_n222 ) );
  INV_X1 u0_uk_U17 (.ZN( u0_uk_n100 ) , .A( u0_uk_n214 ) );
  OAI21_X1 u0_uk_U175 (.ZN( u0_K16_30 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n632 ) , .A( u0_uk_n902 ) );
  NAND2_X1 u0_uk_U176 (.A1( u0_uk_K_r14_45 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n902 ) );
  OAI22_X1 u0_uk_U178 (.ZN( u0_K12_14 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n165 ) , .B2( u0_uk_n170 ) , .B1( u0_uk_n202 ) );
  INV_X1 u0_uk_U187 (.ZN( u0_K2_14 ) , .A( u0_uk_n866 ) );
  AOI22_X1 u0_uk_U188 (.B2( u0_uk_K_r0_11 ) , .A2( u0_uk_K_r0_32 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n866 ) );
  INV_X1 u0_uk_U198 (.ZN( u0_K3_24 ) , .A( u0_uk_n851 ) );
  AOI22_X1 u0_uk_U199 (.B2( u0_uk_K_r1_17 ) , .A2( u0_uk_K_r1_41 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n851 ) );
  INV_X1 u0_uk_U20 (.ZN( u0_uk_n109 ) , .A( u0_uk_n214 ) );
  INV_X1 u0_uk_U210 (.ZN( u0_K4_31 ) , .A( u0_uk_n826 ) );
  INV_X1 u0_uk_U218 (.ZN( u0_K11_31 ) , .A( u0_uk_n992 ) );
  AOI22_X1 u0_uk_U219 (.B2( u0_uk_K_r9_22 ) , .A2( u0_uk_K_r9_30 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n992 ) );
  INV_X1 u0_uk_U221 (.ZN( u0_K11_39 ) , .A( u0_uk_n988 ) );
  AOI22_X1 u0_uk_U222 (.B2( u0_uk_K_r9_30 ) , .A2( u0_uk_K_r9_7 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n988 ) );
  OAI22_X1 u0_uk_U229 (.ZN( u0_K3_31 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n549 ) , .B2( u0_uk_n555 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U25 (.ZN( u0_uk_n146 ) , .A( u0_uk_n148 ) );
  INV_X1 u0_uk_U26 (.ZN( u0_uk_n129 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U266 (.ZN( u0_K7_44 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n378 ) , .B2( u0_uk_n399 ) );
  OAI22_X1 u0_uk_U267 (.ZN( u0_K7_48 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n257 ) , .A2( u0_uk_n367 ) , .B2( u0_uk_n387 ) );
  BUF_X1 u0_uk_U27 (.Z( u0_uk_n163 ) , .A( u0_uk_n217 ) );
  OAI22_X1 u0_uk_U278 (.ZN( u0_K10_6 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n162 ) , .B2( u0_uk_n239 ) , .A2( u0_uk_n267 ) );
  BUF_X1 u0_uk_U28 (.Z( u0_uk_n147 ) , .A( u0_uk_n250 ) );
  OAI22_X1 u0_uk_U286 (.ZN( u0_K12_8 ) , .A2( u0_uk_n136 ) , .B2( u0_uk_n157 ) , .A1( u0_uk_n191 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U293 (.ZN( u0_K3_8 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n562 ) , .A2( u0_uk_n578 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U3 (.ZN( u0_uk_n142 ) , .A( u0_uk_n191 ) );
  BUF_X1 u0_uk_U31 (.Z( u0_uk_n155 ) , .A( u0_uk_n223 ) );
  BUF_X1 u0_uk_U32 (.Z( u0_uk_n148 ) , .A( u0_uk_n240 ) );
  BUF_X1 u0_uk_U33 (.Z( u0_uk_n191 ) , .A( u0_uk_n209 ) );
  OAI22_X1 u0_uk_U332 (.ZN( u0_K11_4 ) , .A1( u0_uk_n118 ) , .A2( u0_uk_n189 ) , .B2( u0_uk_n195 ) , .B1( u0_uk_n202 ) );
  INV_X1 u0_uk_U333 (.ZN( u0_K7_46 ) , .A( u0_uk_n765 ) );
  OAI22_X1 u0_uk_U339 (.ZN( u0_K10_4 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n227 ) , .B2( u0_uk_n246 ) , .B1( u0_uk_n92 ) );
  BUF_X1 u0_uk_U34 (.Z( u0_uk_n164 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U340 (.ZN( u0_K7_4 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n361 ) , .B2( u0_uk_n384 ) );
  OAI22_X1 u0_uk_U347 (.ZN( u0_K3_4 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n557 ) , .B2( u0_uk_n565 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U362 (.ZN( u0_K11_40 ) , .B2( u0_uk_n216 ) , .A2( u0_uk_n224 ) , .A1( u0_uk_n240 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U364 (.ZN( u0_K7_40 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n394 ) , .A2( u0_uk_n406 ) );
  OAI22_X1 u0_uk_U366 (.ZN( u0_K2_40 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n592 ) , .A2( u0_uk_n623 ) );
  BUF_X1 u0_uk_U38 (.Z( u0_uk_n203 ) , .A( u0_uk_n208 ) );
  OAI22_X1 u0_uk_U388 (.ZN( u0_K11_1 ) , .A2( u0_uk_n183 ) , .B2( u0_uk_n200 ) , .A1( u0_uk_n238 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U389 (.ZN( u0_K3_1 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n568 ) , .B2( u0_uk_n573 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U390 (.ZN( u0_K2_1 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n583 ) , .B2( u0_uk_n604 ) );
  OAI21_X1 u0_uk_U398 (.ZN( u0_K3_16 ) , .B1( u0_uk_n102 ) , .B2( u0_uk_n540 ) , .A( u0_uk_n853 ) );
  BUF_X1 u0_uk_U40 (.Z( u0_uk_n230 ) , .A( u0_uk_n257 ) );
  OAI22_X1 u0_uk_U408 (.ZN( u0_K11_9 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n195 ) , .B1( u0_uk_n203 ) , .B2( u0_uk_n225 ) );
  BUF_X1 u0_uk_U41 (.Z( u0_uk_n214 ) , .A( u0_uk_n257 ) );
  OAI21_X1 u0_uk_U422 (.ZN( u0_K3_9 ) , .B1( u0_uk_n209 ) , .B2( u0_uk_n563 ) , .A( u0_uk_n840 ) );
  NAND2_X1 u0_uk_U423 (.A1( u0_uk_K_r1_18 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n840 ) );
  OAI22_X1 u0_uk_U424 (.ZN( u0_K2_9 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n597 ) , .A2( u0_uk_n626 ) );
  BUF_X1 u0_uk_U43 (.Z( u0_uk_n220 ) , .A( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U430 (.ZN( u0_K16_16 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n644 ) , .B2( u0_uk_n651 ) );
  OAI22_X1 u0_uk_U431 (.ZN( u0_K2_16 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n596 ) , .B2( u0_uk_n614 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U436 (.ZN( u0_K11_33 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n199 ) , .B2( u0_uk_n205 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U447 (.ZN( u0_K7_33 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n374 ) , .B2( u0_uk_n394 ) );
  OAI22_X1 u0_uk_U449 (.ZN( u0_K4_33 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n148 ) , .A2( u0_uk_n532 ) , .B2( u0_uk_n539 ) );
  BUF_X1 u0_uk_U45 (.A( u0_uk_n238 ) , .Z( u0_uk_n240 ) );
  OAI22_X1 u0_uk_U450 (.ZN( u0_K3_33 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n549 ) , .B2( u0_uk_n566 ) );
  OAI22_X1 u0_uk_U456 (.ZN( u0_K12_37 ) , .A2( u0_uk_n139 ) , .B2( u0_uk_n179 ) , .A1( u0_uk_n238 ) , .B1( u0_uk_n92 ) );
  BUF_X1 u0_uk_U47 (.Z( u0_uk_n217 ) , .A( u0_uk_n240 ) );
  BUF_X1 u0_uk_U48 (.Z( u0_uk_n222 ) , .A( u0_uk_n250 ) );
  BUF_X1 u0_uk_U49 (.Z( u0_uk_n231 ) , .A( u0_uk_n250 ) );
  OAI22_X1 u0_uk_U490 (.ZN( u0_K11_2 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n181 ) , .B2( u0_uk_n215 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U491 (.ZN( u0_K3_2 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n552 ) , .B2( u0_uk_n557 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U492 (.ZN( u0_K2_2 ) , .A1( u0_uk_n164 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n583 ) , .B2( u0_uk_n615 ) );
  OAI21_X1 u0_uk_U520 (.ZN( u0_K12_12 ) , .B1( u0_uk_n109 ) , .B2( u0_uk_n169 ) , .A( u0_uk_n981 ) );
  BUF_X1 u0_uk_U53 (.A( u0_uk_n163 ) , .Z( u0_uk_n208 ) );
  OAI21_X1 u0_uk_U534 (.ZN( u0_K16_17 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n661 ) , .A( u0_uk_n907 ) );
  NAND2_X1 u0_uk_U535 (.A1( u0_uk_K_r14_10 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n907 ) );
  BUF_X1 u0_uk_U54 (.Z( u0_uk_n251 ) , .A( u0_uk_n257 ) );
  INV_X1 u0_uk_U540 (.ZN( u0_K12_17 ) , .A( u0_uk_n979 ) );
  AOI22_X1 u0_uk_U541 (.B2( u0_uk_K_r10_18 ) , .A2( u0_uk_K_r10_41 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n979 ) );
  OAI22_X1 u0_uk_U547 (.ZN( u0_K3_36 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n544 ) , .B2( u0_uk_n579 ) , .A1( u0_uk_n94 ) );
  BUF_X1 u0_uk_U55 (.A( u0_uk_n250 ) , .Z( u0_uk_n252 ) );
  INV_X1 u0_uk_U552 (.ZN( u0_K16_29 ) , .A( u0_uk_n904 ) );
  OAI22_X1 u0_uk_U555 (.ZN( u0_K12_38 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n153 ) , .B2( u0_uk_n180 ) );
  OAI22_X1 u0_uk_U556 (.ZN( u0_K11_38 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n203 ) , .A2( u0_uk_n210 ) , .B2( u0_uk_n218 ) );
  INV_X1 u0_uk_U558 (.ZN( u0_K7_36 ) , .A( u0_uk_n768 ) );
  AOI22_X1 u0_uk_U559 (.B2( u0_uk_K_r5_1 ) , .A2( u0_uk_K_r5_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n257 ) , .ZN( u0_uk_n768 ) );
  BUF_X1 u0_uk_U56 (.Z( u0_uk_n250 ) , .A( u0_uk_n257 ) );
  INV_X1 u0_uk_U560 (.ZN( u0_K11_36 ) , .A( u0_uk_n990 ) );
  OAI21_X1 u0_uk_U575 (.ZN( u0_K11_10 ) , .A( u0_uk_n1004 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n225 ) );
  OAI22_X1 u0_uk_U588 (.ZN( u0_K3_22 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n542 ) , .B2( u0_uk_n577 ) );
  INV_X1 u0_uk_U6 (.A( u0_uk_n231 ) , .ZN( u0_uk_n93 ) );
  INV_X1 u0_uk_U60 (.ZN( u0_K11_34 ) , .A( u0_uk_n991 ) );
  OAI22_X1 u0_uk_U604 (.ZN( u0_K11_35 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n185 ) , .B2( u0_uk_n193 ) , .B1( u0_uk_n222 ) );
  OAI21_X1 u0_uk_U606 (.ZN( u0_K7_35 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n406 ) , .A( u0_uk_n769 ) );
  NAND2_X1 u0_uk_U607 (.A1( u0_uk_K_r5_37 ) , .ZN( u0_uk_n769 ) , .A2( u0_uk_n92 ) );
  AOI22_X1 u0_uk_U61 (.B2( u0_uk_K_r9_45 ) , .A2( u0_uk_K_r9_49 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n991 ) );
  OAI22_X1 u0_uk_U627 (.ZN( u0_K11_11 ) , .A1( u0_uk_n145 ) , .A2( u0_uk_n206 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U634 (.ZN( u0_K3_11 ) , .A1( u0_uk_n11 ) , .B1( u0_uk_n242 ) , .B2( u0_uk_n573 ) , .A2( u0_uk_n578 ) );
  NAND2_X1 u0_uk_U636 (.A1( u0_uk_K_r0_25 ) , .A2( u0_uk_n109 ) , .ZN( u0_uk_n867 ) );
  OAI22_X1 u0_uk_U651 (.ZN( u0_K7_43 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n374 ) , .A2( u0_uk_n403 ) );
  OAI22_X1 u0_uk_U655 (.ZN( u0_K11_3 ) , .A2( u0_uk_n201 ) , .B2( u0_uk_n219 ) , .A1( u0_uk_n222 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U676 (.A1( u0_uk_K_r2_29 ) , .A2( u0_uk_n100 ) , .ZN( u0_uk_n823 ) );
  OAI21_X1 u0_uk_U682 (.ZN( u0_K11_7 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n197 ) , .A( u0_uk_n983 ) );
  NAND2_X1 u0_uk_U683 (.A1( u0_uk_K_r9_33 ) , .A2( u0_uk_n146 ) , .ZN( u0_uk_n983 ) );
  NAND2_X1 u0_uk_U693 (.A1( u0_uk_K_r0_22 ) , .ZN( u0_uk_n863 ) , .A2( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U694 (.ZN( u0_K16_25 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n240 ) , .A2( u0_uk_n642 ) , .B2( u0_uk_n649 ) );
  OAI22_X1 u0_uk_U70 (.ZN( u0_K4_34 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n208 ) , .A2( u0_uk_n506 ) , .B2( u0_uk_n522 ) );
  OAI21_X1 u0_uk_U714 (.ZN( u0_K10_2 ) , .A( u0_uk_n1015 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n266 ) );
  NAND2_X1 u0_uk_U715 (.A1( u0_uk_K_r8_41 ) , .ZN( u0_uk_n1015 ) , .A2( u0_uk_n220 ) );
  OAI22_X1 u0_uk_U716 (.ZN( u0_K4_32 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n508 ) , .A2( u0_uk_n532 ) );
  OAI22_X1 u0_uk_U719 (.ZN( u0_K11_32 ) , .A2( u0_uk_n198 ) , .A1( u0_uk_n208 ) , .B2( u0_uk_n218 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U722 (.ZN( u0_K3_32 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n545 ) , .B2( u0_uk_n580 ) );
  OAI22_X1 u0_uk_U729 (.ZN( u0_K11_42 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n186 ) , .B2( u0_uk_n194 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U735 (.ZN( u0_K2_42 ) , .A1( u0_uk_n188 ) , .A2( u0_uk_n584 ) , .B2( u0_uk_n592 ) , .B1( u0_uk_n83 ) );
  INV_X1 u0_uk_U736 (.ZN( u0_K7_42 ) , .A( u0_uk_n766 ) );
  OAI22_X1 u0_uk_U74 (.ZN( u0_K16_23 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n640 ) , .B2( u0_uk_n645 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U750 (.ZN( u0_K16_27 ) , .B1( u0_uk_n109 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n658 ) , .B2( u0_uk_n663 ) );
  OAI22_X1 u0_uk_U751 (.ZN( u0_K12_13 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n137 ) , .B2( u0_uk_n169 ) , .B1( u0_uk_n238 ) );
  OAI22_X1 u0_uk_U755 (.ZN( u0_K2_13 ) , .B1( u0_uk_n164 ) , .B2( u0_uk_n598 ) , .A2( u0_uk_n627 ) , .A1( u0_uk_n83 ) );
  OAI21_X1 u0_uk_U788 (.ZN( u0_K16_13 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n631 ) , .A( u0_uk_n909 ) );
  NAND2_X1 u0_uk_U789 (.A1( u0_uk_K_r14_46 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n909 ) );
  OAI21_X1 u0_uk_U800 (.ZN( u0_K7_1 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n396 ) , .A( u0_uk_n781 ) );
  NAND2_X1 u0_uk_U801 (.A1( u0_uk_K_r5_10 ) , .A2( u0_uk_n147 ) , .ZN( u0_uk_n781 ) );
  OAI22_X1 u0_uk_U814 (.ZN( u0_K2_18 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n588 ) , .B2( u0_uk_n619 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U821 (.ZN( u0_K3_20 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n562 ) , .B2( u0_uk_n568 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U822 (.ZN( u0_K16_20 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n629 ) , .B2( u0_uk_n636 ) );
  OAI21_X1 u0_uk_U84 (.ZN( u0_K11_41 ) , .B2( u0_uk_n186 ) , .B1( u0_uk_n203 ) , .A( u0_uk_n987 ) );
  OAI22_X1 u0_uk_U849 (.ZN( u0_K7_3 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n188 ) , .A2( u0_uk_n371 ) , .B2( u0_uk_n393 ) );
  NAND2_X1 u0_uk_U85 (.A1( u0_uk_K_r9_31 ) , .A2( u0_uk_n220 ) , .ZN( u0_uk_n987 ) );
  OAI21_X1 u0_uk_U858 (.ZN( u0_K3_3 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n540 ) , .A( u0_uk_n846 ) );
  NAND2_X1 u0_uk_U859 (.A1( u0_uk_K_r1_47 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n846 ) );
  INV_X1 u0_uk_U86 (.ZN( u0_K2_41 ) , .A( u0_uk_n858 ) );
  OAI21_X1 u0_uk_U864 (.ZN( u0_K10_1 ) , .A( u0_uk_n1021 ) , .B2( u0_uk_n258 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U869 (.ZN( u0_K10_5 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n246 ) , .B2( u0_uk_n263 ) , .B1( u0_uk_n94 ) );
  AOI22_X1 u0_uk_U87 (.B2( u0_uk_K_r0_28 ) , .A2( u0_uk_K_r0_49 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n858 ) );
  OAI22_X1 u0_uk_U881 (.ZN( u0_K12_10 ) , .B1( u0_uk_n142 ) , .A2( u0_uk_n149 ) , .B2( u0_uk_n170 ) , .A1( u0_uk_n191 ) );
  OAI22_X1 u0_uk_U882 (.ZN( u0_K12_11 ) , .B2( u0_uk_n149 ) , .A2( u0_uk_n175 ) , .A1( u0_uk_n182 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U894 (.ZN( u0_K10_3 ) , .A2( u0_uk_n235 ) , .A1( u0_uk_n238 ) , .B2( u0_uk_n255 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U9 (.A( u0_uk_n147 ) , .ZN( u0_uk_n17 ) );
  OAI22_X1 u0_uk_U90 (.ZN( u0_K7_41 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n372 ) , .A2( u0_uk_n402 ) );
  OAI22_X1 u0_uk_U903 (.ZN( u0_K3_21 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n542 ) , .B2( u0_uk_n567 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U908 (.ZN( u0_K16_21 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n654 ) , .B2( u0_uk_n661 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U915 (.ZN( u0_K3_13 ) , .A1( u0_uk_n191 ) , .A2( u0_uk_n564 ) , .B2( u0_uk_n569 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U916 (.ZN( u0_K4_36 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n208 ) , .A2( u0_uk_n507 ) , .B2( u0_uk_n512 ) );
  OAI22_X1 u0_uk_U917 (.ZN( u0_K2_17 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n611 ) , .A2( u0_uk_n627 ) );
  INV_X1 u0_uk_U92 (.ZN( u0_K11_5 ) , .A( u0_uk_n984 ) );
  OAI22_X1 u0_uk_U922 (.ZN( u0_K7_39 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n365 ) , .B2( u0_uk_n372 ) );
  OAI22_X1 u0_uk_U928 (.ZN( u0_K2_39 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n607 ) , .A2( u0_uk_n622 ) , .B1( u0_uk_n83 ) );
  AOI22_X1 u0_uk_U93 (.B2( u0_uk_K_r9_19 ) , .A2( u0_uk_K_r9_25 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n984 ) );
  OAI22_X1 u0_uk_U932 (.ZN( u0_K12_16 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n165 ) , .A2( u0_uk_n177 ) );
  OAI22_X1 u0_uk_U935 (.ZN( u0_K11_6 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n183 ) , .B2( u0_uk_n189 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U939 (.ZN( u0_K12_18 ) , .A1( u0_uk_n100 ) , .B2( u0_uk_n137 ) , .B1( u0_uk_n163 ) , .A2( u0_uk_n175 ) );
  OAI22_X1 u0_uk_U968 (.ZN( u0_K2_38 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n593 ) , .B2( u0_uk_n612 ) );
  OAI22_X1 u0_uk_U969 (.ZN( u0_K7_37 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n365 ) , .B2( u0_uk_n389 ) );
  OAI22_X1 u0_uk_U970 (.ZN( u0_K2_37 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n594 ) , .A2( u0_uk_n621 ) );
  OAI22_X1 u0_uk_U976 (.ZN( u0_K7_45 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n213 ) , .A2( u0_uk_n381 ) , .B2( u0_uk_n398 ) );
  OAI22_X1 u0_uk_U980 (.ZN( u0_K2_3 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n604 ) , .B2( u0_uk_n619 ) );
  OAI22_X1 u0_uk_U982 (.ZN( u0_K3_6 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n571 ) , .A2( u0_uk_n576 ) );
  OAI22_X1 u0_uk_U985 (.ZN( u0_K3_7 ) , .B1( u0_uk_n238 ) , .A2( u0_uk_n547 ) , .B2( u0_uk_n565 ) , .A1( u0_uk_n99 ) );
  NAND2_X1 u0_uk_U995 (.A1( u0_uk_K_r5_5 ) , .ZN( u0_uk_n778 ) , .A2( u0_uk_n93 ) );
  OAI21_X1 u0_uk_U998 (.ZN( u0_K3_35 ) , .B2( u0_uk_n580 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n847 ) );
  NAND2_X1 u0_uk_U999 (.A1( u0_uk_K_r1_7 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n847 ) );
  XOR2_X1 u1_U104 (.B( u1_L12_24 ) , .Z( u1_N439 ) , .A( u1_out13_24 ) );
  XOR2_X1 u1_U105 (.B( u1_L12_23 ) , .Z( u1_N438 ) , .A( u1_out13_23 ) );
  XOR2_X1 u1_U111 (.B( u1_L12_17 ) , .Z( u1_N432 ) , .A( u1_out13_17 ) );
  XOR2_X1 u1_U112 (.B( u1_L12_16 ) , .Z( u1_N431 ) , .A( u1_out13_16 ) );
  XOR2_X1 u1_U120 (.B( u1_L12_9 ) , .Z( u1_N424 ) , .A( u1_out13_9 ) );
  XOR2_X1 u1_U123 (.B( u1_L12_6 ) , .Z( u1_N421 ) , .A( u1_out13_6 ) );
  XOR2_X1 u1_U125 (.B( u1_L0_11 ) , .Z( u1_N42 ) , .A( u1_out1_11 ) );
  XOR2_X1 u1_U132 (.B( u1_L11_30 ) , .Z( u1_N413 ) , .A( u1_out12_30 ) );
  XOR2_X1 u1_U133 (.B( u1_L11_29 ) , .Z( u1_N412 ) , .A( u1_out12_29 ) );
  XOR2_X1 u1_U134 (.B( u1_L11_28 ) , .Z( u1_N411 ) , .A( u1_out12_28 ) );
  XOR2_X1 u1_U139 (.B( u1_L11_24 ) , .Z( u1_N407 ) , .A( u1_out12_24 ) );
  XOR2_X1 u1_U144 (.B( u1_L11_19 ) , .Z( u1_N402 ) , .A( u1_out12_19 ) );
  XOR2_X1 u1_U145 (.B( u1_L11_18 ) , .Z( u1_N401 ) , .A( u1_out12_18 ) );
  XOR2_X1 u1_U149 (.B( u1_L11_16 ) , .Z( u1_N399 ) , .A( u1_out12_16 ) );
  XOR2_X1 u1_U15 (.B( u1_L1_25 ) , .Z( u1_N88 ) , .A( u1_out2_25 ) );
  XOR2_X1 u1_U152 (.B( u1_L11_13 ) , .Z( u1_N396 ) , .A( u1_out12_13 ) );
  XOR2_X1 u1_U154 (.B( u1_L11_11 ) , .Z( u1_N394 ) , .A( u1_out12_11 ) );
  XOR2_X1 u1_U160 (.B( u1_L11_6 ) , .Z( u1_N389 ) , .A( u1_out12_6 ) );
  XOR2_X1 u1_U162 (.B( u1_L11_4 ) , .Z( u1_N387 ) , .A( u1_out12_4 ) );
  XOR2_X1 u1_U164 (.B( u1_L11_2 ) , .Z( u1_N385 ) , .A( u1_out12_2 ) );
  XOR2_X1 u1_U17 (.B( u1_L1_23 ) , .Z( u1_N86 ) , .A( u1_out2_23 ) );
  XOR2_X1 u1_U203 (.B( u1_L0_4 ) , .Z( u1_N35 ) , .A( u1_out1_4 ) );
  XOR2_X1 u1_U23 (.B( u1_L1_17 ) , .Z( u1_N80 ) , .A( u1_out2_17 ) );
  XOR2_X1 u1_U27 (.B( u1_L1_14 ) , .Z( u1_N77 ) , .A( u1_out2_14 ) );
  XOR2_X1 u1_U3 (.B( u1_L2_4 ) , .Z( u1_N99 ) , .A( u1_out3_4 ) );
  XOR2_X1 u1_U311 (.B( u1_L6_29 ) , .Z( u1_N252 ) , .A( u1_out7_29 ) );
  XOR2_X1 u1_U32 (.B( u1_L1_9 ) , .Z( u1_N72 ) , .A( u1_out2_9 ) );
  XOR2_X1 u1_U322 (.B( u1_L6_19 ) , .Z( u1_N242 ) , .A( u1_out7_19 ) );
  XOR2_X1 u1_U33 (.B( u1_L1_8 ) , .Z( u1_N71 ) , .A( u1_out2_8 ) );
  XOR2_X1 u1_U331 (.B( u1_L6_11 ) , .Z( u1_N234 ) , .A( u1_out7_11 ) );
  XOR2_X1 u1_U339 (.B( u1_L6_4 ) , .Z( u1_N227 ) , .A( u1_out7_4 ) );
  XOR2_X1 u1_U384 (.B( u1_L4_28 ) , .Z( u1_N187 ) , .A( u1_out5_28 ) );
  XOR2_X1 u1_U39 (.B( u1_L1_3 ) , .Z( u1_N66 ) , .A( u1_out2_3 ) );
  XOR2_X1 u1_U395 (.B( u1_L4_18 ) , .Z( u1_N177 ) , .A( u1_out5_18 ) );
  XOR2_X1 u1_U4 (.B( u1_L2_3 ) , .Z( u1_N98 ) , .A( u1_out3_3 ) );
  XOR2_X1 u1_U400 (.B( u1_L4_13 ) , .Z( u1_N172 ) , .A( u1_out5_13 ) );
  XOR2_X1 u1_U412 (.B( u1_L4_2 ) , .Z( u1_N161 ) , .A( u1_out5_2 ) );
  XOR2_X1 u1_U45 (.B( u1_L0_29 ) , .Z( u1_N60 ) , .A( u1_out1_29 ) );
  XOR2_X1 u1_U452 (.B( u1_L2_30 ) , .Z( u1_N125 ) , .A( u1_out3_30 ) );
  XOR2_X1 u1_U453 (.B( u1_L2_29 ) , .Z( u1_N124 ) , .A( u1_out3_29 ) );
  XOR2_X1 u1_U455 (.B( u1_L2_27 ) , .Z( u1_N122 ) , .A( u1_out3_27 ) );
  XOR2_X1 u1_U457 (.B( u1_L2_25 ) , .Z( u1_N120 ) , .A( u1_out3_25 ) );
  XOR2_X1 u1_U459 (.B( u1_L2_24 ) , .Z( u1_N119 ) , .A( u1_out3_24 ) );
  XOR2_X1 u1_U462 (.B( u1_L2_21 ) , .Z( u1_N116 ) , .A( u1_out3_21 ) );
  XOR2_X1 u1_U464 (.B( u1_L2_19 ) , .Z( u1_N114 ) , .A( u1_out3_19 ) );
  XOR2_X1 u1_U467 (.B( u1_L2_16 ) , .Z( u1_N111 ) , .A( u1_out3_16 ) );
  XOR2_X1 u1_U468 (.B( u1_L2_15 ) , .Z( u1_N110 ) , .A( u1_out3_15 ) );
  XOR2_X1 u1_U470 (.B( u1_L2_14 ) , .Z( u1_N109 ) , .A( u1_out3_14 ) );
  XOR2_X1 u1_U473 (.B( u1_L2_11 ) , .Z( u1_N106 ) , .A( u1_out3_11 ) );
  XOR2_X1 u1_U476 (.B( u1_L2_8 ) , .Z( u1_N103 ) , .A( u1_out3_8 ) );
  XOR2_X1 u1_U478 (.B( u1_L2_6 ) , .Z( u1_N101 ) , .A( u1_out3_6 ) );
  XOR2_X1 u1_U479 (.B( u1_L2_5 ) , .Z( u1_N100 ) , .A( u1_out3_5 ) );
  XOR2_X1 u1_U487 (.Z( u1_FP_5 ) , .B( u1_L14_5 ) , .A( u1_out15_5 ) );
  XOR2_X1 u1_U496 (.Z( u1_FP_27 ) , .B( u1_L14_27 ) , .A( u1_out15_27 ) );
  XOR2_X1 u1_U502 (.Z( u1_FP_21 ) , .B( u1_L14_21 ) , .A( u1_out15_21 ) );
  XOR2_X1 u1_U509 (.Z( u1_FP_15 ) , .B( u1_L14_15 ) , .A( u1_out15_15 ) );
  XOR2_X1 u1_U56 (.B( u1_L0_19 ) , .Z( u1_N50 ) , .A( u1_out1_19 ) );
  XOR2_X1 u1_U64 (.B( u1_L13_28 ) , .Z( u1_N475 ) , .A( u1_out14_28 ) );
  XOR2_X1 u1_U75 (.B( u1_L13_18 ) , .Z( u1_N465 ) , .A( u1_out14_18 ) );
  XOR2_X1 u1_U8 (.B( u1_L1_31 ) , .Z( u1_N94 ) , .A( u1_out2_31 ) );
  XOR2_X1 u1_U80 (.B( u1_L13_13 ) , .Z( u1_N460 ) , .A( u1_out14_13 ) );
  XOR2_X1 u1_U93 (.B( u1_L13_2 ) , .Z( u1_N449 ) , .A( u1_out14_2 ) );
  XOR2_X1 u1_U96 (.B( u1_L12_31 ) , .Z( u1_N446 ) , .A( u1_out13_31 ) );
  XOR2_X1 u1_U97 (.B( u1_L12_30 ) , .Z( u1_N445 ) , .A( u1_out13_30 ) );
  XOR2_X1 u1_u12_U1 (.B( u1_K13_9 ) , .A( u1_R11_6 ) , .Z( u1_u12_X_9 ) );
  XOR2_X1 u1_u12_U22 (.B( u1_K13_34 ) , .A( u1_R11_23 ) , .Z( u1_u12_X_34 ) );
  XOR2_X1 u1_u12_U23 (.B( u1_K13_33 ) , .A( u1_R11_22 ) , .Z( u1_u12_X_33 ) );
  XOR2_X1 u1_u12_U42 (.B( u1_K13_16 ) , .A( u1_R11_11 ) , .Z( u1_u12_X_16 ) );
  XOR2_X1 u1_u12_U43 (.B( u1_K13_15 ) , .A( u1_R11_10 ) , .Z( u1_u12_X_15 ) );
  XOR2_X1 u1_u12_U45 (.B( u1_K13_13 ) , .A( u1_R11_8 ) , .Z( u1_u12_X_13 ) );
  XOR2_X1 u1_u12_U47 (.B( u1_K13_11 ) , .A( u1_R11_8 ) , .Z( u1_u12_X_11 ) );
  XOR2_X1 u1_u12_U48 (.B( u1_K13_10 ) , .A( u1_R11_7 ) , .Z( u1_u12_X_10 ) );
  NOR2_X1 u1_u12_u1_U10 (.A1( u1_u12_u1_n112 ) , .A2( u1_u12_u1_n116 ) , .ZN( u1_u12_u1_n118 ) );
  NAND3_X1 u1_u12_u1_U100 (.ZN( u1_u12_u1_n113 ) , .A1( u1_u12_u1_n120 ) , .A3( u1_u12_u1_n133 ) , .A2( u1_u12_u1_n155 ) );
  OAI21_X1 u1_u12_u1_U11 (.ZN( u1_u12_u1_n101 ) , .B1( u1_u12_u1_n141 ) , .A( u1_u12_u1_n146 ) , .B2( u1_u12_u1_n183 ) );
  AOI21_X1 u1_u12_u1_U12 (.B2( u1_u12_u1_n155 ) , .B1( u1_u12_u1_n156 ) , .ZN( u1_u12_u1_n157 ) , .A( u1_u12_u1_n174 ) );
  NAND2_X1 u1_u12_u1_U13 (.ZN( u1_u12_u1_n140 ) , .A2( u1_u12_u1_n150 ) , .A1( u1_u12_u1_n155 ) );
  NAND2_X1 u1_u12_u1_U14 (.A1( u1_u12_u1_n131 ) , .ZN( u1_u12_u1_n147 ) , .A2( u1_u12_u1_n153 ) );
  INV_X1 u1_u12_u1_U15 (.A( u1_u12_u1_n139 ) , .ZN( u1_u12_u1_n174 ) );
  OR4_X1 u1_u12_u1_U16 (.A4( u1_u12_u1_n106 ) , .A3( u1_u12_u1_n107 ) , .ZN( u1_u12_u1_n108 ) , .A1( u1_u12_u1_n117 ) , .A2( u1_u12_u1_n184 ) );
  AOI21_X1 u1_u12_u1_U17 (.ZN( u1_u12_u1_n106 ) , .A( u1_u12_u1_n112 ) , .B1( u1_u12_u1_n154 ) , .B2( u1_u12_u1_n156 ) );
  INV_X1 u1_u12_u1_U18 (.A( u1_u12_u1_n101 ) , .ZN( u1_u12_u1_n184 ) );
  AOI21_X1 u1_u12_u1_U19 (.ZN( u1_u12_u1_n107 ) , .B1( u1_u12_u1_n134 ) , .B2( u1_u12_u1_n149 ) , .A( u1_u12_u1_n174 ) );
  INV_X1 u1_u12_u1_U20 (.A( u1_u12_u1_n112 ) , .ZN( u1_u12_u1_n171 ) );
  NAND2_X1 u1_u12_u1_U21 (.ZN( u1_u12_u1_n141 ) , .A1( u1_u12_u1_n153 ) , .A2( u1_u12_u1_n156 ) );
  AND2_X1 u1_u12_u1_U22 (.A1( u1_u12_u1_n123 ) , .ZN( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n161 ) );
  NAND2_X1 u1_u12_u1_U23 (.A2( u1_u12_u1_n115 ) , .A1( u1_u12_u1_n116 ) , .ZN( u1_u12_u1_n148 ) );
  NAND2_X1 u1_u12_u1_U24 (.A2( u1_u12_u1_n133 ) , .A1( u1_u12_u1_n135 ) , .ZN( u1_u12_u1_n159 ) );
  NAND2_X1 u1_u12_u1_U25 (.A2( u1_u12_u1_n115 ) , .A1( u1_u12_u1_n120 ) , .ZN( u1_u12_u1_n132 ) );
  INV_X1 u1_u12_u1_U26 (.A( u1_u12_u1_n154 ) , .ZN( u1_u12_u1_n178 ) );
  INV_X1 u1_u12_u1_U27 (.A( u1_u12_u1_n151 ) , .ZN( u1_u12_u1_n183 ) );
  AND2_X1 u1_u12_u1_U28 (.A1( u1_u12_u1_n129 ) , .A2( u1_u12_u1_n133 ) , .ZN( u1_u12_u1_n149 ) );
  INV_X1 u1_u12_u1_U29 (.A( u1_u12_u1_n131 ) , .ZN( u1_u12_u1_n180 ) );
  INV_X1 u1_u12_u1_U3 (.A( u1_u12_u1_n159 ) , .ZN( u1_u12_u1_n182 ) );
  AOI221_X1 u1_u12_u1_U30 (.B1( u1_u12_u1_n140 ) , .ZN( u1_u12_u1_n167 ) , .B2( u1_u12_u1_n172 ) , .C2( u1_u12_u1_n175 ) , .C1( u1_u12_u1_n178 ) , .A( u1_u12_u1_n188 ) );
  INV_X1 u1_u12_u1_U31 (.ZN( u1_u12_u1_n188 ) , .A( u1_u12_u1_n97 ) );
  AOI211_X1 u1_u12_u1_U32 (.A( u1_u12_u1_n118 ) , .C1( u1_u12_u1_n132 ) , .C2( u1_u12_u1_n139 ) , .B( u1_u12_u1_n96 ) , .ZN( u1_u12_u1_n97 ) );
  AOI21_X1 u1_u12_u1_U33 (.B2( u1_u12_u1_n121 ) , .B1( u1_u12_u1_n135 ) , .A( u1_u12_u1_n152 ) , .ZN( u1_u12_u1_n96 ) );
  OAI221_X1 u1_u12_u1_U34 (.A( u1_u12_u1_n119 ) , .C2( u1_u12_u1_n129 ) , .ZN( u1_u12_u1_n138 ) , .B2( u1_u12_u1_n152 ) , .C1( u1_u12_u1_n174 ) , .B1( u1_u12_u1_n187 ) );
  INV_X1 u1_u12_u1_U35 (.A( u1_u12_u1_n148 ) , .ZN( u1_u12_u1_n187 ) );
  AOI211_X1 u1_u12_u1_U36 (.B( u1_u12_u1_n117 ) , .A( u1_u12_u1_n118 ) , .ZN( u1_u12_u1_n119 ) , .C2( u1_u12_u1_n146 ) , .C1( u1_u12_u1_n159 ) );
  NOR2_X1 u1_u12_u1_U37 (.A1( u1_u12_u1_n168 ) , .A2( u1_u12_u1_n176 ) , .ZN( u1_u12_u1_n98 ) );
  AOI211_X1 u1_u12_u1_U38 (.B( u1_u12_u1_n162 ) , .A( u1_u12_u1_n163 ) , .C2( u1_u12_u1_n164 ) , .ZN( u1_u12_u1_n165 ) , .C1( u1_u12_u1_n171 ) );
  AOI21_X1 u1_u12_u1_U39 (.A( u1_u12_u1_n160 ) , .B2( u1_u12_u1_n161 ) , .ZN( u1_u12_u1_n162 ) , .B1( u1_u12_u1_n182 ) );
  AOI221_X1 u1_u12_u1_U4 (.A( u1_u12_u1_n138 ) , .C2( u1_u12_u1_n139 ) , .C1( u1_u12_u1_n140 ) , .B2( u1_u12_u1_n141 ) , .ZN( u1_u12_u1_n142 ) , .B1( u1_u12_u1_n175 ) );
  OR2_X1 u1_u12_u1_U40 (.A2( u1_u12_u1_n157 ) , .A1( u1_u12_u1_n158 ) , .ZN( u1_u12_u1_n163 ) );
  NAND2_X1 u1_u12_u1_U41 (.A1( u1_u12_u1_n128 ) , .ZN( u1_u12_u1_n146 ) , .A2( u1_u12_u1_n160 ) );
  NAND2_X1 u1_u12_u1_U42 (.A2( u1_u12_u1_n112 ) , .ZN( u1_u12_u1_n139 ) , .A1( u1_u12_u1_n152 ) );
  NAND2_X1 u1_u12_u1_U43 (.A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n156 ) , .A2( u1_u12_u1_n99 ) );
  NOR2_X1 u1_u12_u1_U44 (.ZN( u1_u12_u1_n117 ) , .A1( u1_u12_u1_n121 ) , .A2( u1_u12_u1_n160 ) );
  OAI21_X1 u1_u12_u1_U45 (.B2( u1_u12_u1_n123 ) , .ZN( u1_u12_u1_n145 ) , .B1( u1_u12_u1_n160 ) , .A( u1_u12_u1_n185 ) );
  INV_X1 u1_u12_u1_U46 (.A( u1_u12_u1_n122 ) , .ZN( u1_u12_u1_n185 ) );
  AOI21_X1 u1_u12_u1_U47 (.B2( u1_u12_u1_n120 ) , .B1( u1_u12_u1_n121 ) , .ZN( u1_u12_u1_n122 ) , .A( u1_u12_u1_n128 ) );
  AOI21_X1 u1_u12_u1_U48 (.A( u1_u12_u1_n128 ) , .B2( u1_u12_u1_n129 ) , .ZN( u1_u12_u1_n130 ) , .B1( u1_u12_u1_n150 ) );
  NAND2_X1 u1_u12_u1_U49 (.ZN( u1_u12_u1_n112 ) , .A1( u1_u12_u1_n169 ) , .A2( u1_u12_u1_n170 ) );
  AOI211_X1 u1_u12_u1_U5 (.ZN( u1_u12_u1_n124 ) , .A( u1_u12_u1_n138 ) , .C2( u1_u12_u1_n139 ) , .B( u1_u12_u1_n145 ) , .C1( u1_u12_u1_n147 ) );
  NAND2_X1 u1_u12_u1_U50 (.ZN( u1_u12_u1_n129 ) , .A2( u1_u12_u1_n95 ) , .A1( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U51 (.A1( u1_u12_u1_n102 ) , .ZN( u1_u12_u1_n154 ) , .A2( u1_u12_u1_n99 ) );
  NAND2_X1 u1_u12_u1_U52 (.A2( u1_u12_u1_n100 ) , .ZN( u1_u12_u1_n135 ) , .A1( u1_u12_u1_n99 ) );
  AOI21_X1 u1_u12_u1_U53 (.A( u1_u12_u1_n152 ) , .B2( u1_u12_u1_n153 ) , .B1( u1_u12_u1_n154 ) , .ZN( u1_u12_u1_n158 ) );
  INV_X1 u1_u12_u1_U54 (.A( u1_u12_u1_n160 ) , .ZN( u1_u12_u1_n175 ) );
  NAND2_X1 u1_u12_u1_U55 (.A1( u1_u12_u1_n100 ) , .ZN( u1_u12_u1_n116 ) , .A2( u1_u12_u1_n95 ) );
  NAND2_X1 u1_u12_u1_U56 (.A1( u1_u12_u1_n102 ) , .ZN( u1_u12_u1_n131 ) , .A2( u1_u12_u1_n95 ) );
  NAND2_X1 u1_u12_u1_U57 (.A2( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n121 ) , .A1( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U58 (.A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n153 ) , .A2( u1_u12_u1_n98 ) );
  NAND2_X1 u1_u12_u1_U59 (.A2( u1_u12_u1_n104 ) , .A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n133 ) );
  AOI22_X1 u1_u12_u1_U6 (.B2( u1_u12_u1_n113 ) , .A2( u1_u12_u1_n114 ) , .ZN( u1_u12_u1_n125 ) , .A1( u1_u12_u1_n171 ) , .B1( u1_u12_u1_n173 ) );
  NAND2_X1 u1_u12_u1_U60 (.ZN( u1_u12_u1_n150 ) , .A2( u1_u12_u1_n98 ) , .A1( u1_u12_u1_n99 ) );
  NAND2_X1 u1_u12_u1_U61 (.A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n155 ) , .A2( u1_u12_u1_n95 ) );
  OAI21_X1 u1_u12_u1_U62 (.ZN( u1_u12_u1_n109 ) , .B1( u1_u12_u1_n129 ) , .B2( u1_u12_u1_n160 ) , .A( u1_u12_u1_n167 ) );
  NAND2_X1 u1_u12_u1_U63 (.A2( u1_u12_u1_n100 ) , .A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n120 ) );
  NAND2_X1 u1_u12_u1_U64 (.A1( u1_u12_u1_n102 ) , .A2( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n115 ) );
  NAND2_X1 u1_u12_u1_U65 (.A2( u1_u12_u1_n100 ) , .A1( u1_u12_u1_n104 ) , .ZN( u1_u12_u1_n151 ) );
  NAND2_X1 u1_u12_u1_U66 (.A2( u1_u12_u1_n103 ) , .A1( u1_u12_u1_n105 ) , .ZN( u1_u12_u1_n161 ) );
  INV_X1 u1_u12_u1_U67 (.A( u1_u12_u1_n152 ) , .ZN( u1_u12_u1_n173 ) );
  INV_X1 u1_u12_u1_U68 (.A( u1_u12_u1_n128 ) , .ZN( u1_u12_u1_n172 ) );
  NAND2_X1 u1_u12_u1_U69 (.A2( u1_u12_u1_n102 ) , .A1( u1_u12_u1_n103 ) , .ZN( u1_u12_u1_n123 ) );
  NAND2_X1 u1_u12_u1_U7 (.ZN( u1_u12_u1_n114 ) , .A1( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n156 ) );
  NOR2_X1 u1_u12_u1_U70 (.A2( u1_u12_X_7 ) , .A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n95 ) );
  NOR2_X1 u1_u12_u1_U71 (.A1( u1_u12_X_12 ) , .A2( u1_u12_X_9 ) , .ZN( u1_u12_u1_n100 ) );
  NOR2_X1 u1_u12_u1_U72 (.A2( u1_u12_X_8 ) , .A1( u1_u12_u1_n177 ) , .ZN( u1_u12_u1_n99 ) );
  NOR2_X1 u1_u12_u1_U73 (.A2( u1_u12_X_12 ) , .ZN( u1_u12_u1_n102 ) , .A1( u1_u12_u1_n176 ) );
  NOR2_X1 u1_u12_u1_U74 (.A2( u1_u12_X_9 ) , .ZN( u1_u12_u1_n105 ) , .A1( u1_u12_u1_n168 ) );
  NAND2_X1 u1_u12_u1_U75 (.A1( u1_u12_X_10 ) , .ZN( u1_u12_u1_n160 ) , .A2( u1_u12_u1_n169 ) );
  NAND2_X1 u1_u12_u1_U76 (.A2( u1_u12_X_10 ) , .A1( u1_u12_X_11 ) , .ZN( u1_u12_u1_n152 ) );
  NAND2_X1 u1_u12_u1_U77 (.A1( u1_u12_X_11 ) , .ZN( u1_u12_u1_n128 ) , .A2( u1_u12_u1_n170 ) );
  AND2_X1 u1_u12_u1_U78 (.A2( u1_u12_X_7 ) , .A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n104 ) );
  AND2_X1 u1_u12_u1_U79 (.A1( u1_u12_X_8 ) , .ZN( u1_u12_u1_n103 ) , .A2( u1_u12_u1_n177 ) );
  AOI22_X1 u1_u12_u1_U8 (.B2( u1_u12_u1_n136 ) , .A2( u1_u12_u1_n137 ) , .ZN( u1_u12_u1_n143 ) , .A1( u1_u12_u1_n171 ) , .B1( u1_u12_u1_n173 ) );
  INV_X1 u1_u12_u1_U80 (.A( u1_u12_X_10 ) , .ZN( u1_u12_u1_n170 ) );
  INV_X1 u1_u12_u1_U81 (.A( u1_u12_X_9 ) , .ZN( u1_u12_u1_n176 ) );
  INV_X1 u1_u12_u1_U82 (.A( u1_u12_X_11 ) , .ZN( u1_u12_u1_n169 ) );
  INV_X1 u1_u12_u1_U83 (.A( u1_u12_X_12 ) , .ZN( u1_u12_u1_n168 ) );
  INV_X1 u1_u12_u1_U84 (.A( u1_u12_X_7 ) , .ZN( u1_u12_u1_n177 ) );
  NAND4_X1 u1_u12_u1_U85 (.ZN( u1_out12_28 ) , .A4( u1_u12_u1_n124 ) , .A3( u1_u12_u1_n125 ) , .A2( u1_u12_u1_n126 ) , .A1( u1_u12_u1_n127 ) );
  OAI21_X1 u1_u12_u1_U86 (.ZN( u1_u12_u1_n127 ) , .B2( u1_u12_u1_n139 ) , .B1( u1_u12_u1_n175 ) , .A( u1_u12_u1_n183 ) );
  OAI21_X1 u1_u12_u1_U87 (.ZN( u1_u12_u1_n126 ) , .B2( u1_u12_u1_n140 ) , .A( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n178 ) );
  NAND4_X1 u1_u12_u1_U88 (.ZN( u1_out12_18 ) , .A4( u1_u12_u1_n165 ) , .A3( u1_u12_u1_n166 ) , .A1( u1_u12_u1_n167 ) , .A2( u1_u12_u1_n186 ) );
  AOI22_X1 u1_u12_u1_U89 (.B2( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n147 ) , .A2( u1_u12_u1_n148 ) , .ZN( u1_u12_u1_n166 ) , .A1( u1_u12_u1_n172 ) );
  INV_X1 u1_u12_u1_U9 (.A( u1_u12_u1_n147 ) , .ZN( u1_u12_u1_n181 ) );
  INV_X1 u1_u12_u1_U90 (.A( u1_u12_u1_n145 ) , .ZN( u1_u12_u1_n186 ) );
  NAND4_X1 u1_u12_u1_U91 (.ZN( u1_out12_2 ) , .A4( u1_u12_u1_n142 ) , .A3( u1_u12_u1_n143 ) , .A2( u1_u12_u1_n144 ) , .A1( u1_u12_u1_n179 ) );
  OAI21_X1 u1_u12_u1_U92 (.B2( u1_u12_u1_n132 ) , .ZN( u1_u12_u1_n144 ) , .A( u1_u12_u1_n146 ) , .B1( u1_u12_u1_n180 ) );
  INV_X1 u1_u12_u1_U93 (.A( u1_u12_u1_n130 ) , .ZN( u1_u12_u1_n179 ) );
  OR4_X1 u1_u12_u1_U94 (.ZN( u1_out12_13 ) , .A4( u1_u12_u1_n108 ) , .A3( u1_u12_u1_n109 ) , .A2( u1_u12_u1_n110 ) , .A1( u1_u12_u1_n111 ) );
  AOI21_X1 u1_u12_u1_U95 (.ZN( u1_u12_u1_n111 ) , .A( u1_u12_u1_n128 ) , .B2( u1_u12_u1_n131 ) , .B1( u1_u12_u1_n135 ) );
  AOI21_X1 u1_u12_u1_U96 (.ZN( u1_u12_u1_n110 ) , .A( u1_u12_u1_n116 ) , .B1( u1_u12_u1_n152 ) , .B2( u1_u12_u1_n160 ) );
  NAND3_X1 u1_u12_u1_U97 (.A3( u1_u12_u1_n149 ) , .A2( u1_u12_u1_n150 ) , .A1( u1_u12_u1_n151 ) , .ZN( u1_u12_u1_n164 ) );
  NAND3_X1 u1_u12_u1_U98 (.A3( u1_u12_u1_n134 ) , .A2( u1_u12_u1_n135 ) , .ZN( u1_u12_u1_n136 ) , .A1( u1_u12_u1_n151 ) );
  NAND3_X1 u1_u12_u1_U99 (.A1( u1_u12_u1_n133 ) , .ZN( u1_u12_u1_n137 ) , .A2( u1_u12_u1_n154 ) , .A3( u1_u12_u1_n181 ) );
  OAI22_X1 u1_u12_u2_U10 (.B1( u1_u12_u2_n151 ) , .A2( u1_u12_u2_n152 ) , .A1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n160 ) , .B2( u1_u12_u2_n168 ) );
  NAND3_X1 u1_u12_u2_U100 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n98 ) );
  NOR3_X1 u1_u12_u2_U11 (.A1( u1_u12_u2_n150 ) , .ZN( u1_u12_u2_n151 ) , .A3( u1_u12_u2_n175 ) , .A2( u1_u12_u2_n188 ) );
  AOI21_X1 u1_u12_u2_U12 (.B2( u1_u12_u2_n123 ) , .ZN( u1_u12_u2_n125 ) , .A( u1_u12_u2_n171 ) , .B1( u1_u12_u2_n184 ) );
  INV_X1 u1_u12_u2_U13 (.A( u1_u12_u2_n150 ) , .ZN( u1_u12_u2_n184 ) );
  AOI21_X1 u1_u12_u2_U14 (.ZN( u1_u12_u2_n144 ) , .B2( u1_u12_u2_n155 ) , .A( u1_u12_u2_n172 ) , .B1( u1_u12_u2_n185 ) );
  AOI21_X1 u1_u12_u2_U15 (.B2( u1_u12_u2_n143 ) , .ZN( u1_u12_u2_n145 ) , .B1( u1_u12_u2_n152 ) , .A( u1_u12_u2_n171 ) );
  INV_X1 u1_u12_u2_U16 (.A( u1_u12_u2_n156 ) , .ZN( u1_u12_u2_n171 ) );
  INV_X1 u1_u12_u2_U17 (.A( u1_u12_u2_n120 ) , .ZN( u1_u12_u2_n188 ) );
  NAND2_X1 u1_u12_u2_U18 (.A2( u1_u12_u2_n122 ) , .ZN( u1_u12_u2_n150 ) , .A1( u1_u12_u2_n152 ) );
  INV_X1 u1_u12_u2_U19 (.A( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n170 ) );
  INV_X1 u1_u12_u2_U20 (.A( u1_u12_u2_n137 ) , .ZN( u1_u12_u2_n173 ) );
  NAND2_X1 u1_u12_u2_U21 (.A1( u1_u12_u2_n132 ) , .A2( u1_u12_u2_n139 ) , .ZN( u1_u12_u2_n157 ) );
  INV_X1 u1_u12_u2_U22 (.A( u1_u12_u2_n113 ) , .ZN( u1_u12_u2_n178 ) );
  INV_X1 u1_u12_u2_U23 (.A( u1_u12_u2_n139 ) , .ZN( u1_u12_u2_n175 ) );
  INV_X1 u1_u12_u2_U24 (.A( u1_u12_u2_n155 ) , .ZN( u1_u12_u2_n181 ) );
  INV_X1 u1_u12_u2_U25 (.A( u1_u12_u2_n119 ) , .ZN( u1_u12_u2_n177 ) );
  INV_X1 u1_u12_u2_U26 (.A( u1_u12_u2_n116 ) , .ZN( u1_u12_u2_n180 ) );
  INV_X1 u1_u12_u2_U27 (.A( u1_u12_u2_n131 ) , .ZN( u1_u12_u2_n179 ) );
  INV_X1 u1_u12_u2_U28 (.A( u1_u12_u2_n154 ) , .ZN( u1_u12_u2_n176 ) );
  NAND2_X1 u1_u12_u2_U29 (.A2( u1_u12_u2_n116 ) , .A1( u1_u12_u2_n117 ) , .ZN( u1_u12_u2_n118 ) );
  NOR2_X1 u1_u12_u2_U3 (.ZN( u1_u12_u2_n121 ) , .A2( u1_u12_u2_n177 ) , .A1( u1_u12_u2_n180 ) );
  INV_X1 u1_u12_u2_U30 (.A( u1_u12_u2_n132 ) , .ZN( u1_u12_u2_n182 ) );
  INV_X1 u1_u12_u2_U31 (.A( u1_u12_u2_n158 ) , .ZN( u1_u12_u2_n183 ) );
  OAI21_X1 u1_u12_u2_U32 (.A( u1_u12_u2_n156 ) , .B1( u1_u12_u2_n157 ) , .ZN( u1_u12_u2_n158 ) , .B2( u1_u12_u2_n179 ) );
  NOR2_X1 u1_u12_u2_U33 (.ZN( u1_u12_u2_n156 ) , .A1( u1_u12_u2_n166 ) , .A2( u1_u12_u2_n169 ) );
  NOR2_X1 u1_u12_u2_U34 (.A2( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n137 ) , .A1( u1_u12_u2_n140 ) );
  NOR2_X1 u1_u12_u2_U35 (.A2( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n153 ) , .A1( u1_u12_u2_n156 ) );
  AOI211_X1 u1_u12_u2_U36 (.ZN( u1_u12_u2_n130 ) , .C1( u1_u12_u2_n138 ) , .C2( u1_u12_u2_n179 ) , .B( u1_u12_u2_n96 ) , .A( u1_u12_u2_n97 ) );
  OAI22_X1 u1_u12_u2_U37 (.B1( u1_u12_u2_n133 ) , .A2( u1_u12_u2_n137 ) , .A1( u1_u12_u2_n152 ) , .B2( u1_u12_u2_n168 ) , .ZN( u1_u12_u2_n97 ) );
  OAI221_X1 u1_u12_u2_U38 (.B1( u1_u12_u2_n113 ) , .C1( u1_u12_u2_n132 ) , .A( u1_u12_u2_n149 ) , .B2( u1_u12_u2_n171 ) , .C2( u1_u12_u2_n172 ) , .ZN( u1_u12_u2_n96 ) );
  OAI221_X1 u1_u12_u2_U39 (.A( u1_u12_u2_n115 ) , .C2( u1_u12_u2_n123 ) , .B2( u1_u12_u2_n143 ) , .B1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n163 ) , .C1( u1_u12_u2_n168 ) );
  INV_X1 u1_u12_u2_U4 (.A( u1_u12_u2_n134 ) , .ZN( u1_u12_u2_n185 ) );
  OAI21_X1 u1_u12_u2_U40 (.A( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n115 ) , .B1( u1_u12_u2_n176 ) , .B2( u1_u12_u2_n178 ) );
  OAI221_X1 u1_u12_u2_U41 (.A( u1_u12_u2_n135 ) , .B2( u1_u12_u2_n136 ) , .B1( u1_u12_u2_n137 ) , .ZN( u1_u12_u2_n162 ) , .C2( u1_u12_u2_n167 ) , .C1( u1_u12_u2_n185 ) );
  AND3_X1 u1_u12_u2_U42 (.A3( u1_u12_u2_n131 ) , .A2( u1_u12_u2_n132 ) , .A1( u1_u12_u2_n133 ) , .ZN( u1_u12_u2_n136 ) );
  AOI22_X1 u1_u12_u2_U43 (.ZN( u1_u12_u2_n135 ) , .B1( u1_u12_u2_n140 ) , .A1( u1_u12_u2_n156 ) , .B2( u1_u12_u2_n180 ) , .A2( u1_u12_u2_n188 ) );
  AOI21_X1 u1_u12_u2_U44 (.ZN( u1_u12_u2_n149 ) , .B1( u1_u12_u2_n173 ) , .B2( u1_u12_u2_n188 ) , .A( u1_u12_u2_n95 ) );
  AND3_X1 u1_u12_u2_U45 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n156 ) , .ZN( u1_u12_u2_n95 ) );
  OAI21_X1 u1_u12_u2_U46 (.A( u1_u12_u2_n101 ) , .B2( u1_u12_u2_n121 ) , .B1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n164 ) );
  NAND2_X1 u1_u12_u2_U47 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n155 ) );
  NAND2_X1 u1_u12_u2_U48 (.A2( u1_u12_u2_n105 ) , .A1( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n143 ) );
  NAND2_X1 u1_u12_u2_U49 (.A1( u1_u12_u2_n104 ) , .A2( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n152 ) );
  NOR4_X1 u1_u12_u2_U5 (.A4( u1_u12_u2_n124 ) , .A3( u1_u12_u2_n125 ) , .A2( u1_u12_u2_n126 ) , .A1( u1_u12_u2_n127 ) , .ZN( u1_u12_u2_n128 ) );
  NAND2_X1 u1_u12_u2_U50 (.A1( u1_u12_u2_n100 ) , .A2( u1_u12_u2_n105 ) , .ZN( u1_u12_u2_n132 ) );
  INV_X1 u1_u12_u2_U51 (.A( u1_u12_u2_n140 ) , .ZN( u1_u12_u2_n168 ) );
  INV_X1 u1_u12_u2_U52 (.A( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n167 ) );
  OAI21_X1 u1_u12_u2_U53 (.A( u1_u12_u2_n141 ) , .B2( u1_u12_u2_n142 ) , .ZN( u1_u12_u2_n146 ) , .B1( u1_u12_u2_n153 ) );
  OAI21_X1 u1_u12_u2_U54 (.A( u1_u12_u2_n140 ) , .ZN( u1_u12_u2_n141 ) , .B1( u1_u12_u2_n176 ) , .B2( u1_u12_u2_n177 ) );
  NOR3_X1 u1_u12_u2_U55 (.ZN( u1_u12_u2_n142 ) , .A3( u1_u12_u2_n175 ) , .A2( u1_u12_u2_n178 ) , .A1( u1_u12_u2_n181 ) );
  NAND2_X1 u1_u12_u2_U56 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n113 ) );
  NAND2_X1 u1_u12_u2_U57 (.A1( u1_u12_u2_n106 ) , .A2( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n131 ) );
  NAND2_X1 u1_u12_u2_U58 (.A1( u1_u12_u2_n103 ) , .A2( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n139 ) );
  NAND2_X1 u1_u12_u2_U59 (.A1( u1_u12_u2_n103 ) , .A2( u1_u12_u2_n105 ) , .ZN( u1_u12_u2_n133 ) );
  AOI21_X1 u1_u12_u2_U6 (.B2( u1_u12_u2_n119 ) , .ZN( u1_u12_u2_n127 ) , .A( u1_u12_u2_n137 ) , .B1( u1_u12_u2_n155 ) );
  NAND2_X1 u1_u12_u2_U60 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n103 ) , .ZN( u1_u12_u2_n154 ) );
  NAND2_X1 u1_u12_u2_U61 (.A2( u1_u12_u2_n103 ) , .A1( u1_u12_u2_n104 ) , .ZN( u1_u12_u2_n119 ) );
  NAND2_X1 u1_u12_u2_U62 (.A2( u1_u12_u2_n107 ) , .A1( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n123 ) );
  NAND2_X1 u1_u12_u2_U63 (.A1( u1_u12_u2_n104 ) , .A2( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n122 ) );
  INV_X1 u1_u12_u2_U64 (.A( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n172 ) );
  NAND2_X1 u1_u12_u2_U65 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n102 ) , .ZN( u1_u12_u2_n116 ) );
  NAND2_X1 u1_u12_u2_U66 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n120 ) );
  NAND2_X1 u1_u12_u2_U67 (.A2( u1_u12_u2_n105 ) , .A1( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n117 ) );
  INV_X1 u1_u12_u2_U68 (.ZN( u1_u12_u2_n187 ) , .A( u1_u12_u2_n99 ) );
  OAI21_X1 u1_u12_u2_U69 (.B1( u1_u12_u2_n137 ) , .B2( u1_u12_u2_n143 ) , .A( u1_u12_u2_n98 ) , .ZN( u1_u12_u2_n99 ) );
  AOI21_X1 u1_u12_u2_U7 (.ZN( u1_u12_u2_n124 ) , .B1( u1_u12_u2_n131 ) , .B2( u1_u12_u2_n143 ) , .A( u1_u12_u2_n172 ) );
  NOR2_X1 u1_u12_u2_U70 (.A2( u1_u12_X_16 ) , .ZN( u1_u12_u2_n140 ) , .A1( u1_u12_u2_n166 ) );
  NOR2_X1 u1_u12_u2_U71 (.A2( u1_u12_X_13 ) , .A1( u1_u12_X_14 ) , .ZN( u1_u12_u2_n100 ) );
  NOR2_X1 u1_u12_u2_U72 (.A2( u1_u12_X_16 ) , .A1( u1_u12_X_17 ) , .ZN( u1_u12_u2_n138 ) );
  NOR2_X1 u1_u12_u2_U73 (.A2( u1_u12_X_15 ) , .A1( u1_u12_X_18 ) , .ZN( u1_u12_u2_n104 ) );
  NOR2_X1 u1_u12_u2_U74 (.A2( u1_u12_X_14 ) , .ZN( u1_u12_u2_n103 ) , .A1( u1_u12_u2_n174 ) );
  NOR2_X1 u1_u12_u2_U75 (.A2( u1_u12_X_15 ) , .ZN( u1_u12_u2_n102 ) , .A1( u1_u12_u2_n165 ) );
  NOR2_X1 u1_u12_u2_U76 (.A2( u1_u12_X_17 ) , .ZN( u1_u12_u2_n114 ) , .A1( u1_u12_u2_n169 ) );
  AND2_X1 u1_u12_u2_U77 (.A1( u1_u12_X_15 ) , .ZN( u1_u12_u2_n105 ) , .A2( u1_u12_u2_n165 ) );
  AND2_X1 u1_u12_u2_U78 (.A2( u1_u12_X_15 ) , .A1( u1_u12_X_18 ) , .ZN( u1_u12_u2_n107 ) );
  AND2_X1 u1_u12_u2_U79 (.A1( u1_u12_X_14 ) , .ZN( u1_u12_u2_n106 ) , .A2( u1_u12_u2_n174 ) );
  AOI21_X1 u1_u12_u2_U8 (.B2( u1_u12_u2_n120 ) , .B1( u1_u12_u2_n121 ) , .ZN( u1_u12_u2_n126 ) , .A( u1_u12_u2_n167 ) );
  AND2_X1 u1_u12_u2_U80 (.A1( u1_u12_X_13 ) , .A2( u1_u12_X_14 ) , .ZN( u1_u12_u2_n108 ) );
  INV_X1 u1_u12_u2_U81 (.A( u1_u12_X_16 ) , .ZN( u1_u12_u2_n169 ) );
  INV_X1 u1_u12_u2_U82 (.A( u1_u12_X_17 ) , .ZN( u1_u12_u2_n166 ) );
  INV_X1 u1_u12_u2_U83 (.A( u1_u12_X_13 ) , .ZN( u1_u12_u2_n174 ) );
  INV_X1 u1_u12_u2_U84 (.A( u1_u12_X_18 ) , .ZN( u1_u12_u2_n165 ) );
  NAND4_X1 u1_u12_u2_U85 (.ZN( u1_out12_30 ) , .A4( u1_u12_u2_n147 ) , .A3( u1_u12_u2_n148 ) , .A2( u1_u12_u2_n149 ) , .A1( u1_u12_u2_n187 ) );
  AOI21_X1 u1_u12_u2_U86 (.B2( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n148 ) , .A( u1_u12_u2_n162 ) , .B1( u1_u12_u2_n182 ) );
  NOR3_X1 u1_u12_u2_U87 (.A3( u1_u12_u2_n144 ) , .A2( u1_u12_u2_n145 ) , .A1( u1_u12_u2_n146 ) , .ZN( u1_u12_u2_n147 ) );
  NAND4_X1 u1_u12_u2_U88 (.ZN( u1_out12_24 ) , .A4( u1_u12_u2_n111 ) , .A3( u1_u12_u2_n112 ) , .A1( u1_u12_u2_n130 ) , .A2( u1_u12_u2_n187 ) );
  AOI221_X1 u1_u12_u2_U89 (.A( u1_u12_u2_n109 ) , .B1( u1_u12_u2_n110 ) , .ZN( u1_u12_u2_n111 ) , .C1( u1_u12_u2_n134 ) , .C2( u1_u12_u2_n170 ) , .B2( u1_u12_u2_n173 ) );
  OAI22_X1 u1_u12_u2_U9 (.ZN( u1_u12_u2_n109 ) , .A2( u1_u12_u2_n113 ) , .B2( u1_u12_u2_n133 ) , .B1( u1_u12_u2_n167 ) , .A1( u1_u12_u2_n168 ) );
  AOI21_X1 u1_u12_u2_U90 (.ZN( u1_u12_u2_n112 ) , .B2( u1_u12_u2_n156 ) , .A( u1_u12_u2_n164 ) , .B1( u1_u12_u2_n181 ) );
  NAND4_X1 u1_u12_u2_U91 (.ZN( u1_out12_16 ) , .A4( u1_u12_u2_n128 ) , .A3( u1_u12_u2_n129 ) , .A1( u1_u12_u2_n130 ) , .A2( u1_u12_u2_n186 ) );
  AOI22_X1 u1_u12_u2_U92 (.A2( u1_u12_u2_n118 ) , .ZN( u1_u12_u2_n129 ) , .A1( u1_u12_u2_n140 ) , .B1( u1_u12_u2_n157 ) , .B2( u1_u12_u2_n170 ) );
  INV_X1 u1_u12_u2_U93 (.A( u1_u12_u2_n163 ) , .ZN( u1_u12_u2_n186 ) );
  OR4_X1 u1_u12_u2_U94 (.ZN( u1_out12_6 ) , .A4( u1_u12_u2_n161 ) , .A3( u1_u12_u2_n162 ) , .A2( u1_u12_u2_n163 ) , .A1( u1_u12_u2_n164 ) );
  OR3_X1 u1_u12_u2_U95 (.A2( u1_u12_u2_n159 ) , .A1( u1_u12_u2_n160 ) , .ZN( u1_u12_u2_n161 ) , .A3( u1_u12_u2_n183 ) );
  AOI21_X1 u1_u12_u2_U96 (.B2( u1_u12_u2_n154 ) , .B1( u1_u12_u2_n155 ) , .ZN( u1_u12_u2_n159 ) , .A( u1_u12_u2_n167 ) );
  NAND3_X1 u1_u12_u2_U97 (.A2( u1_u12_u2_n117 ) , .A1( u1_u12_u2_n122 ) , .A3( u1_u12_u2_n123 ) , .ZN( u1_u12_u2_n134 ) );
  NAND3_X1 u1_u12_u2_U98 (.ZN( u1_u12_u2_n110 ) , .A2( u1_u12_u2_n131 ) , .A3( u1_u12_u2_n139 ) , .A1( u1_u12_u2_n154 ) );
  NAND3_X1 u1_u12_u2_U99 (.A2( u1_u12_u2_n100 ) , .ZN( u1_u12_u2_n101 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n114 ) );
  INV_X1 u1_u12_u5_U10 (.A( u1_u12_u5_n121 ) , .ZN( u1_u12_u5_n177 ) );
  NOR3_X1 u1_u12_u5_U100 (.A3( u1_u12_u5_n141 ) , .A1( u1_u12_u5_n142 ) , .ZN( u1_u12_u5_n143 ) , .A2( u1_u12_u5_n191 ) );
  NAND4_X1 u1_u12_u5_U101 (.ZN( u1_out12_4 ) , .A4( u1_u12_u5_n112 ) , .A2( u1_u12_u5_n113 ) , .A1( u1_u12_u5_n114 ) , .A3( u1_u12_u5_n195 ) );
  AOI211_X1 u1_u12_u5_U102 (.A( u1_u12_u5_n110 ) , .C1( u1_u12_u5_n111 ) , .ZN( u1_u12_u5_n112 ) , .B( u1_u12_u5_n118 ) , .C2( u1_u12_u5_n177 ) );
  AOI222_X1 u1_u12_u5_U103 (.ZN( u1_u12_u5_n113 ) , .A1( u1_u12_u5_n131 ) , .C1( u1_u12_u5_n148 ) , .B2( u1_u12_u5_n174 ) , .C2( u1_u12_u5_n178 ) , .A2( u1_u12_u5_n179 ) , .B1( u1_u12_u5_n99 ) );
  NAND3_X1 u1_u12_u5_U104 (.A2( u1_u12_u5_n154 ) , .A3( u1_u12_u5_n158 ) , .A1( u1_u12_u5_n161 ) , .ZN( u1_u12_u5_n99 ) );
  NOR2_X1 u1_u12_u5_U11 (.ZN( u1_u12_u5_n160 ) , .A2( u1_u12_u5_n173 ) , .A1( u1_u12_u5_n177 ) );
  INV_X1 u1_u12_u5_U12 (.A( u1_u12_u5_n150 ) , .ZN( u1_u12_u5_n174 ) );
  AOI21_X1 u1_u12_u5_U13 (.A( u1_u12_u5_n160 ) , .B2( u1_u12_u5_n161 ) , .ZN( u1_u12_u5_n162 ) , .B1( u1_u12_u5_n192 ) );
  INV_X1 u1_u12_u5_U14 (.A( u1_u12_u5_n159 ) , .ZN( u1_u12_u5_n192 ) );
  AOI21_X1 u1_u12_u5_U15 (.A( u1_u12_u5_n156 ) , .B2( u1_u12_u5_n157 ) , .B1( u1_u12_u5_n158 ) , .ZN( u1_u12_u5_n163 ) );
  AOI21_X1 u1_u12_u5_U16 (.B2( u1_u12_u5_n139 ) , .B1( u1_u12_u5_n140 ) , .ZN( u1_u12_u5_n141 ) , .A( u1_u12_u5_n150 ) );
  OAI21_X1 u1_u12_u5_U17 (.A( u1_u12_u5_n133 ) , .B2( u1_u12_u5_n134 ) , .B1( u1_u12_u5_n135 ) , .ZN( u1_u12_u5_n142 ) );
  OAI21_X1 u1_u12_u5_U18 (.ZN( u1_u12_u5_n133 ) , .B2( u1_u12_u5_n147 ) , .A( u1_u12_u5_n173 ) , .B1( u1_u12_u5_n188 ) );
  NAND2_X1 u1_u12_u5_U19 (.A2( u1_u12_u5_n119 ) , .A1( u1_u12_u5_n123 ) , .ZN( u1_u12_u5_n137 ) );
  INV_X1 u1_u12_u5_U20 (.A( u1_u12_u5_n155 ) , .ZN( u1_u12_u5_n194 ) );
  NAND2_X1 u1_u12_u5_U21 (.A1( u1_u12_u5_n121 ) , .ZN( u1_u12_u5_n132 ) , .A2( u1_u12_u5_n172 ) );
  NAND2_X1 u1_u12_u5_U22 (.A2( u1_u12_u5_n122 ) , .ZN( u1_u12_u5_n136 ) , .A1( u1_u12_u5_n154 ) );
  NAND2_X1 u1_u12_u5_U23 (.A2( u1_u12_u5_n119 ) , .A1( u1_u12_u5_n120 ) , .ZN( u1_u12_u5_n159 ) );
  INV_X1 u1_u12_u5_U24 (.A( u1_u12_u5_n156 ) , .ZN( u1_u12_u5_n175 ) );
  INV_X1 u1_u12_u5_U25 (.A( u1_u12_u5_n158 ) , .ZN( u1_u12_u5_n188 ) );
  INV_X1 u1_u12_u5_U26 (.A( u1_u12_u5_n152 ) , .ZN( u1_u12_u5_n179 ) );
  INV_X1 u1_u12_u5_U27 (.A( u1_u12_u5_n140 ) , .ZN( u1_u12_u5_n182 ) );
  INV_X1 u1_u12_u5_U28 (.A( u1_u12_u5_n151 ) , .ZN( u1_u12_u5_n183 ) );
  INV_X1 u1_u12_u5_U29 (.A( u1_u12_u5_n123 ) , .ZN( u1_u12_u5_n185 ) );
  NOR2_X1 u1_u12_u5_U3 (.ZN( u1_u12_u5_n134 ) , .A1( u1_u12_u5_n183 ) , .A2( u1_u12_u5_n190 ) );
  INV_X1 u1_u12_u5_U30 (.A( u1_u12_u5_n161 ) , .ZN( u1_u12_u5_n184 ) );
  INV_X1 u1_u12_u5_U31 (.A( u1_u12_u5_n139 ) , .ZN( u1_u12_u5_n189 ) );
  INV_X1 u1_u12_u5_U32 (.A( u1_u12_u5_n157 ) , .ZN( u1_u12_u5_n190 ) );
  INV_X1 u1_u12_u5_U33 (.A( u1_u12_u5_n120 ) , .ZN( u1_u12_u5_n193 ) );
  NAND2_X1 u1_u12_u5_U34 (.ZN( u1_u12_u5_n111 ) , .A1( u1_u12_u5_n140 ) , .A2( u1_u12_u5_n155 ) );
  NOR2_X1 u1_u12_u5_U35 (.ZN( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n170 ) , .A2( u1_u12_u5_n180 ) );
  INV_X1 u1_u12_u5_U36 (.A( u1_u12_u5_n117 ) , .ZN( u1_u12_u5_n196 ) );
  OAI221_X1 u1_u12_u5_U37 (.A( u1_u12_u5_n116 ) , .ZN( u1_u12_u5_n117 ) , .B2( u1_u12_u5_n119 ) , .C1( u1_u12_u5_n153 ) , .C2( u1_u12_u5_n158 ) , .B1( u1_u12_u5_n172 ) );
  AOI222_X1 u1_u12_u5_U38 (.ZN( u1_u12_u5_n116 ) , .B2( u1_u12_u5_n145 ) , .C1( u1_u12_u5_n148 ) , .A2( u1_u12_u5_n174 ) , .C2( u1_u12_u5_n177 ) , .B1( u1_u12_u5_n187 ) , .A1( u1_u12_u5_n193 ) );
  INV_X1 u1_u12_u5_U39 (.A( u1_u12_u5_n115 ) , .ZN( u1_u12_u5_n187 ) );
  INV_X1 u1_u12_u5_U4 (.A( u1_u12_u5_n138 ) , .ZN( u1_u12_u5_n191 ) );
  AOI22_X1 u1_u12_u5_U40 (.B2( u1_u12_u5_n131 ) , .A2( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n169 ) , .B1( u1_u12_u5_n174 ) , .A1( u1_u12_u5_n185 ) );
  NOR2_X1 u1_u12_u5_U41 (.A1( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n150 ) , .A2( u1_u12_u5_n173 ) );
  AOI21_X1 u1_u12_u5_U42 (.A( u1_u12_u5_n118 ) , .B2( u1_u12_u5_n145 ) , .ZN( u1_u12_u5_n168 ) , .B1( u1_u12_u5_n186 ) );
  INV_X1 u1_u12_u5_U43 (.A( u1_u12_u5_n122 ) , .ZN( u1_u12_u5_n186 ) );
  NOR2_X1 u1_u12_u5_U44 (.A1( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n152 ) , .A2( u1_u12_u5_n176 ) );
  NOR2_X1 u1_u12_u5_U45 (.A1( u1_u12_u5_n115 ) , .ZN( u1_u12_u5_n118 ) , .A2( u1_u12_u5_n153 ) );
  NOR2_X1 u1_u12_u5_U46 (.A2( u1_u12_u5_n145 ) , .ZN( u1_u12_u5_n156 ) , .A1( u1_u12_u5_n174 ) );
  NOR2_X1 u1_u12_u5_U47 (.ZN( u1_u12_u5_n121 ) , .A2( u1_u12_u5_n145 ) , .A1( u1_u12_u5_n176 ) );
  AOI22_X1 u1_u12_u5_U48 (.ZN( u1_u12_u5_n114 ) , .A2( u1_u12_u5_n137 ) , .A1( u1_u12_u5_n145 ) , .B2( u1_u12_u5_n175 ) , .B1( u1_u12_u5_n193 ) );
  OAI211_X1 u1_u12_u5_U49 (.B( u1_u12_u5_n124 ) , .A( u1_u12_u5_n125 ) , .C2( u1_u12_u5_n126 ) , .C1( u1_u12_u5_n127 ) , .ZN( u1_u12_u5_n128 ) );
  OAI21_X1 u1_u12_u5_U5 (.B2( u1_u12_u5_n136 ) , .B1( u1_u12_u5_n137 ) , .ZN( u1_u12_u5_n138 ) , .A( u1_u12_u5_n177 ) );
  NOR3_X1 u1_u12_u5_U50 (.ZN( u1_u12_u5_n127 ) , .A1( u1_u12_u5_n136 ) , .A3( u1_u12_u5_n148 ) , .A2( u1_u12_u5_n182 ) );
  OAI21_X1 u1_u12_u5_U51 (.ZN( u1_u12_u5_n124 ) , .A( u1_u12_u5_n177 ) , .B2( u1_u12_u5_n183 ) , .B1( u1_u12_u5_n189 ) );
  OAI21_X1 u1_u12_u5_U52 (.ZN( u1_u12_u5_n125 ) , .A( u1_u12_u5_n174 ) , .B2( u1_u12_u5_n185 ) , .B1( u1_u12_u5_n190 ) );
  AOI21_X1 u1_u12_u5_U53 (.A( u1_u12_u5_n153 ) , .B2( u1_u12_u5_n154 ) , .B1( u1_u12_u5_n155 ) , .ZN( u1_u12_u5_n164 ) );
  AOI21_X1 u1_u12_u5_U54 (.ZN( u1_u12_u5_n110 ) , .B1( u1_u12_u5_n122 ) , .B2( u1_u12_u5_n139 ) , .A( u1_u12_u5_n153 ) );
  INV_X1 u1_u12_u5_U55 (.A( u1_u12_u5_n153 ) , .ZN( u1_u12_u5_n176 ) );
  INV_X1 u1_u12_u5_U56 (.A( u1_u12_u5_n126 ) , .ZN( u1_u12_u5_n173 ) );
  AND2_X1 u1_u12_u5_U57 (.A2( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n107 ) , .ZN( u1_u12_u5_n147 ) );
  AND2_X1 u1_u12_u5_U58 (.A2( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n108 ) , .ZN( u1_u12_u5_n148 ) );
  NAND2_X1 u1_u12_u5_U59 (.A1( u1_u12_u5_n105 ) , .A2( u1_u12_u5_n106 ) , .ZN( u1_u12_u5_n158 ) );
  INV_X1 u1_u12_u5_U6 (.A( u1_u12_u5_n135 ) , .ZN( u1_u12_u5_n178 ) );
  NAND2_X1 u1_u12_u5_U60 (.A2( u1_u12_u5_n108 ) , .A1( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n139 ) );
  NAND2_X1 u1_u12_u5_U61 (.A1( u1_u12_u5_n106 ) , .A2( u1_u12_u5_n108 ) , .ZN( u1_u12_u5_n119 ) );
  NAND2_X1 u1_u12_u5_U62 (.A2( u1_u12_u5_n103 ) , .A1( u1_u12_u5_n105 ) , .ZN( u1_u12_u5_n140 ) );
  NAND2_X1 u1_u12_u5_U63 (.A2( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n105 ) , .ZN( u1_u12_u5_n155 ) );
  NAND2_X1 u1_u12_u5_U64 (.A2( u1_u12_u5_n106 ) , .A1( u1_u12_u5_n107 ) , .ZN( u1_u12_u5_n122 ) );
  NAND2_X1 u1_u12_u5_U65 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n106 ) , .ZN( u1_u12_u5_n115 ) );
  NAND2_X1 u1_u12_u5_U66 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n103 ) , .ZN( u1_u12_u5_n161 ) );
  NAND2_X1 u1_u12_u5_U67 (.A1( u1_u12_u5_n105 ) , .A2( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n154 ) );
  INV_X1 u1_u12_u5_U68 (.A( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n172 ) );
  NAND2_X1 u1_u12_u5_U69 (.A1( u1_u12_u5_n103 ) , .A2( u1_u12_u5_n108 ) , .ZN( u1_u12_u5_n123 ) );
  OAI22_X1 u1_u12_u5_U7 (.B2( u1_u12_u5_n149 ) , .B1( u1_u12_u5_n150 ) , .A2( u1_u12_u5_n151 ) , .A1( u1_u12_u5_n152 ) , .ZN( u1_u12_u5_n165 ) );
  NAND2_X1 u1_u12_u5_U70 (.A2( u1_u12_u5_n103 ) , .A1( u1_u12_u5_n107 ) , .ZN( u1_u12_u5_n151 ) );
  NAND2_X1 u1_u12_u5_U71 (.A2( u1_u12_u5_n107 ) , .A1( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n120 ) );
  NAND2_X1 u1_u12_u5_U72 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n109 ) , .ZN( u1_u12_u5_n157 ) );
  AND2_X1 u1_u12_u5_U73 (.A2( u1_u12_u5_n100 ) , .A1( u1_u12_u5_n104 ) , .ZN( u1_u12_u5_n131 ) );
  INV_X1 u1_u12_u5_U74 (.A( u1_u12_u5_n102 ) , .ZN( u1_u12_u5_n195 ) );
  OAI221_X1 u1_u12_u5_U75 (.A( u1_u12_u5_n101 ) , .ZN( u1_u12_u5_n102 ) , .C2( u1_u12_u5_n115 ) , .C1( u1_u12_u5_n126 ) , .B1( u1_u12_u5_n134 ) , .B2( u1_u12_u5_n160 ) );
  OAI21_X1 u1_u12_u5_U76 (.ZN( u1_u12_u5_n101 ) , .B1( u1_u12_u5_n137 ) , .A( u1_u12_u5_n146 ) , .B2( u1_u12_u5_n147 ) );
  NOR2_X1 u1_u12_u5_U77 (.A2( u1_u12_X_34 ) , .A1( u1_u12_X_35 ) , .ZN( u1_u12_u5_n145 ) );
  NOR2_X1 u1_u12_u5_U78 (.A2( u1_u12_X_34 ) , .ZN( u1_u12_u5_n146 ) , .A1( u1_u12_u5_n171 ) );
  NOR2_X1 u1_u12_u5_U79 (.A2( u1_u12_X_31 ) , .A1( u1_u12_X_32 ) , .ZN( u1_u12_u5_n103 ) );
  NOR3_X1 u1_u12_u5_U8 (.A2( u1_u12_u5_n147 ) , .A1( u1_u12_u5_n148 ) , .ZN( u1_u12_u5_n149 ) , .A3( u1_u12_u5_n194 ) );
  NOR2_X1 u1_u12_u5_U80 (.A2( u1_u12_X_36 ) , .ZN( u1_u12_u5_n105 ) , .A1( u1_u12_u5_n180 ) );
  NOR2_X1 u1_u12_u5_U81 (.A2( u1_u12_X_33 ) , .ZN( u1_u12_u5_n108 ) , .A1( u1_u12_u5_n170 ) );
  NOR2_X1 u1_u12_u5_U82 (.A2( u1_u12_X_33 ) , .A1( u1_u12_X_36 ) , .ZN( u1_u12_u5_n107 ) );
  NOR2_X1 u1_u12_u5_U83 (.A2( u1_u12_X_31 ) , .ZN( u1_u12_u5_n104 ) , .A1( u1_u12_u5_n181 ) );
  NAND2_X1 u1_u12_u5_U84 (.A2( u1_u12_X_34 ) , .A1( u1_u12_X_35 ) , .ZN( u1_u12_u5_n153 ) );
  NAND2_X1 u1_u12_u5_U85 (.A1( u1_u12_X_34 ) , .ZN( u1_u12_u5_n126 ) , .A2( u1_u12_u5_n171 ) );
  AND2_X1 u1_u12_u5_U86 (.A1( u1_u12_X_31 ) , .A2( u1_u12_X_32 ) , .ZN( u1_u12_u5_n106 ) );
  AND2_X1 u1_u12_u5_U87 (.A1( u1_u12_X_31 ) , .ZN( u1_u12_u5_n109 ) , .A2( u1_u12_u5_n181 ) );
  INV_X1 u1_u12_u5_U88 (.A( u1_u12_X_33 ) , .ZN( u1_u12_u5_n180 ) );
  INV_X1 u1_u12_u5_U89 (.A( u1_u12_X_35 ) , .ZN( u1_u12_u5_n171 ) );
  NOR2_X1 u1_u12_u5_U9 (.ZN( u1_u12_u5_n135 ) , .A1( u1_u12_u5_n173 ) , .A2( u1_u12_u5_n176 ) );
  INV_X1 u1_u12_u5_U90 (.A( u1_u12_X_36 ) , .ZN( u1_u12_u5_n170 ) );
  INV_X1 u1_u12_u5_U91 (.A( u1_u12_X_32 ) , .ZN( u1_u12_u5_n181 ) );
  NAND4_X1 u1_u12_u5_U92 (.ZN( u1_out12_29 ) , .A4( u1_u12_u5_n129 ) , .A3( u1_u12_u5_n130 ) , .A2( u1_u12_u5_n168 ) , .A1( u1_u12_u5_n196 ) );
  AOI221_X1 u1_u12_u5_U93 (.A( u1_u12_u5_n128 ) , .ZN( u1_u12_u5_n129 ) , .C2( u1_u12_u5_n132 ) , .B2( u1_u12_u5_n159 ) , .B1( u1_u12_u5_n176 ) , .C1( u1_u12_u5_n184 ) );
  AOI222_X1 u1_u12_u5_U94 (.ZN( u1_u12_u5_n130 ) , .A2( u1_u12_u5_n146 ) , .B1( u1_u12_u5_n147 ) , .C2( u1_u12_u5_n175 ) , .B2( u1_u12_u5_n179 ) , .A1( u1_u12_u5_n188 ) , .C1( u1_u12_u5_n194 ) );
  NAND4_X1 u1_u12_u5_U95 (.ZN( u1_out12_19 ) , .A4( u1_u12_u5_n166 ) , .A3( u1_u12_u5_n167 ) , .A2( u1_u12_u5_n168 ) , .A1( u1_u12_u5_n169 ) );
  AOI22_X1 u1_u12_u5_U96 (.B2( u1_u12_u5_n145 ) , .A2( u1_u12_u5_n146 ) , .ZN( u1_u12_u5_n167 ) , .B1( u1_u12_u5_n182 ) , .A1( u1_u12_u5_n189 ) );
  NOR4_X1 u1_u12_u5_U97 (.A4( u1_u12_u5_n162 ) , .A3( u1_u12_u5_n163 ) , .A2( u1_u12_u5_n164 ) , .A1( u1_u12_u5_n165 ) , .ZN( u1_u12_u5_n166 ) );
  NAND4_X1 u1_u12_u5_U98 (.ZN( u1_out12_11 ) , .A4( u1_u12_u5_n143 ) , .A3( u1_u12_u5_n144 ) , .A2( u1_u12_u5_n169 ) , .A1( u1_u12_u5_n196 ) );
  AOI22_X1 u1_u12_u5_U99 (.A2( u1_u12_u5_n132 ) , .ZN( u1_u12_u5_n144 ) , .B2( u1_u12_u5_n145 ) , .B1( u1_u12_u5_n184 ) , .A1( u1_u12_u5_n194 ) );
  XOR2_X1 u1_u13_U16 (.B( u1_K14_3 ) , .A( u1_R12_2 ) , .Z( u1_u13_X_3 ) );
  XOR2_X1 u1_u13_U42 (.B( u1_K14_16 ) , .A( u1_R12_11 ) , .Z( u1_u13_X_16 ) );
  XOR2_X1 u1_u13_U43 (.B( u1_K14_15 ) , .A( u1_R12_10 ) , .Z( u1_u13_X_15 ) );
  XOR2_X1 u1_u13_U6 (.B( u1_K14_4 ) , .A( u1_R12_3 ) , .Z( u1_u13_X_4 ) );
  AND3_X1 u1_u13_u0_U10 (.A2( u1_u13_u0_n112 ) , .ZN( u1_u13_u0_n127 ) , .A3( u1_u13_u0_n130 ) , .A1( u1_u13_u0_n148 ) );
  NAND2_X1 u1_u13_u0_U11 (.ZN( u1_u13_u0_n113 ) , .A1( u1_u13_u0_n139 ) , .A2( u1_u13_u0_n149 ) );
  AND2_X1 u1_u13_u0_U12 (.ZN( u1_u13_u0_n107 ) , .A1( u1_u13_u0_n130 ) , .A2( u1_u13_u0_n140 ) );
  AND2_X1 u1_u13_u0_U13 (.A2( u1_u13_u0_n129 ) , .A1( u1_u13_u0_n130 ) , .ZN( u1_u13_u0_n151 ) );
  AND2_X1 u1_u13_u0_U14 (.A1( u1_u13_u0_n108 ) , .A2( u1_u13_u0_n125 ) , .ZN( u1_u13_u0_n145 ) );
  INV_X1 u1_u13_u0_U15 (.A( u1_u13_u0_n143 ) , .ZN( u1_u13_u0_n173 ) );
  NOR2_X1 u1_u13_u0_U16 (.A2( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n147 ) , .A1( u1_u13_u0_n160 ) );
  INV_X1 u1_u13_u0_U17 (.ZN( u1_u13_u0_n172 ) , .A( u1_u13_u0_n88 ) );
  OAI222_X1 u1_u13_u0_U18 (.C1( u1_u13_u0_n108 ) , .A1( u1_u13_u0_n125 ) , .B2( u1_u13_u0_n128 ) , .B1( u1_u13_u0_n144 ) , .A2( u1_u13_u0_n158 ) , .C2( u1_u13_u0_n161 ) , .ZN( u1_u13_u0_n88 ) );
  NOR2_X1 u1_u13_u0_U19 (.A1( u1_u13_u0_n163 ) , .A2( u1_u13_u0_n164 ) , .ZN( u1_u13_u0_n95 ) );
  AOI21_X1 u1_u13_u0_U20 (.B1( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n132 ) , .A( u1_u13_u0_n165 ) , .B2( u1_u13_u0_n93 ) );
  INV_X1 u1_u13_u0_U21 (.A( u1_u13_u0_n142 ) , .ZN( u1_u13_u0_n165 ) );
  OAI221_X1 u1_u13_u0_U22 (.C1( u1_u13_u0_n121 ) , .ZN( u1_u13_u0_n122 ) , .B2( u1_u13_u0_n127 ) , .A( u1_u13_u0_n143 ) , .B1( u1_u13_u0_n144 ) , .C2( u1_u13_u0_n147 ) );
  OAI22_X1 u1_u13_u0_U23 (.B1( u1_u13_u0_n125 ) , .ZN( u1_u13_u0_n126 ) , .A1( u1_u13_u0_n138 ) , .A2( u1_u13_u0_n146 ) , .B2( u1_u13_u0_n147 ) );
  OAI22_X1 u1_u13_u0_U24 (.B1( u1_u13_u0_n131 ) , .A1( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n147 ) , .A2( u1_u13_u0_n90 ) , .ZN( u1_u13_u0_n91 ) );
  AND3_X1 u1_u13_u0_U25 (.A3( u1_u13_u0_n121 ) , .A2( u1_u13_u0_n125 ) , .A1( u1_u13_u0_n148 ) , .ZN( u1_u13_u0_n90 ) );
  INV_X1 u1_u13_u0_U26 (.A( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n161 ) );
  NOR2_X1 u1_u13_u0_U27 (.A1( u1_u13_u0_n120 ) , .ZN( u1_u13_u0_n143 ) , .A2( u1_u13_u0_n167 ) );
  OAI221_X1 u1_u13_u0_U28 (.C1( u1_u13_u0_n112 ) , .ZN( u1_u13_u0_n120 ) , .B1( u1_u13_u0_n138 ) , .B2( u1_u13_u0_n141 ) , .C2( u1_u13_u0_n147 ) , .A( u1_u13_u0_n172 ) );
  AOI211_X1 u1_u13_u0_U29 (.B( u1_u13_u0_n115 ) , .A( u1_u13_u0_n116 ) , .C2( u1_u13_u0_n117 ) , .C1( u1_u13_u0_n118 ) , .ZN( u1_u13_u0_n119 ) );
  INV_X1 u1_u13_u0_U3 (.A( u1_u13_u0_n113 ) , .ZN( u1_u13_u0_n166 ) );
  AOI22_X1 u1_u13_u0_U30 (.B2( u1_u13_u0_n109 ) , .A2( u1_u13_u0_n110 ) , .ZN( u1_u13_u0_n111 ) , .B1( u1_u13_u0_n118 ) , .A1( u1_u13_u0_n160 ) );
  INV_X1 u1_u13_u0_U31 (.A( u1_u13_u0_n118 ) , .ZN( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U32 (.ZN( u1_u13_u0_n104 ) , .B1( u1_u13_u0_n107 ) , .B2( u1_u13_u0_n141 ) , .A( u1_u13_u0_n144 ) );
  AOI21_X1 u1_u13_u0_U33 (.B1( u1_u13_u0_n127 ) , .B2( u1_u13_u0_n129 ) , .A( u1_u13_u0_n138 ) , .ZN( u1_u13_u0_n96 ) );
  AOI21_X1 u1_u13_u0_U34 (.ZN( u1_u13_u0_n116 ) , .B2( u1_u13_u0_n142 ) , .A( u1_u13_u0_n144 ) , .B1( u1_u13_u0_n166 ) );
  NAND2_X1 u1_u13_u0_U35 (.A1( u1_u13_u0_n100 ) , .A2( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n125 ) );
  NAND2_X1 u1_u13_u0_U36 (.A1( u1_u13_u0_n101 ) , .A2( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n150 ) );
  INV_X1 u1_u13_u0_U37 (.A( u1_u13_u0_n138 ) , .ZN( u1_u13_u0_n160 ) );
  NAND2_X1 u1_u13_u0_U38 (.A1( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n128 ) , .A2( u1_u13_u0_n95 ) );
  NAND2_X1 u1_u13_u0_U39 (.A1( u1_u13_u0_n100 ) , .ZN( u1_u13_u0_n129 ) , .A2( u1_u13_u0_n95 ) );
  AOI21_X1 u1_u13_u0_U4 (.B1( u1_u13_u0_n114 ) , .ZN( u1_u13_u0_n115 ) , .B2( u1_u13_u0_n129 ) , .A( u1_u13_u0_n161 ) );
  NAND2_X1 u1_u13_u0_U40 (.A2( u1_u13_u0_n100 ) , .ZN( u1_u13_u0_n131 ) , .A1( u1_u13_u0_n92 ) );
  NAND2_X1 u1_u13_u0_U41 (.A2( u1_u13_u0_n100 ) , .A1( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n139 ) );
  NAND2_X1 u1_u13_u0_U42 (.ZN( u1_u13_u0_n148 ) , .A1( u1_u13_u0_n93 ) , .A2( u1_u13_u0_n95 ) );
  NAND2_X1 u1_u13_u0_U43 (.A2( u1_u13_u0_n102 ) , .A1( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n149 ) );
  NAND2_X1 u1_u13_u0_U44 (.A2( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n114 ) , .A1( u1_u13_u0_n92 ) );
  NAND2_X1 u1_u13_u0_U45 (.A2( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n121 ) , .A1( u1_u13_u0_n93 ) );
  NAND2_X1 u1_u13_u0_U46 (.ZN( u1_u13_u0_n112 ) , .A2( u1_u13_u0_n92 ) , .A1( u1_u13_u0_n93 ) );
  OR3_X1 u1_u13_u0_U47 (.A3( u1_u13_u0_n152 ) , .A2( u1_u13_u0_n153 ) , .A1( u1_u13_u0_n154 ) , .ZN( u1_u13_u0_n155 ) );
  AOI21_X1 u1_u13_u0_U48 (.B2( u1_u13_u0_n150 ) , .B1( u1_u13_u0_n151 ) , .ZN( u1_u13_u0_n152 ) , .A( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U49 (.A( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n145 ) , .B1( u1_u13_u0_n146 ) , .ZN( u1_u13_u0_n154 ) );
  AOI21_X1 u1_u13_u0_U5 (.B2( u1_u13_u0_n131 ) , .ZN( u1_u13_u0_n134 ) , .B1( u1_u13_u0_n151 ) , .A( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U50 (.A( u1_u13_u0_n147 ) , .B2( u1_u13_u0_n148 ) , .B1( u1_u13_u0_n149 ) , .ZN( u1_u13_u0_n153 ) );
  INV_X1 u1_u13_u0_U51 (.ZN( u1_u13_u0_n171 ) , .A( u1_u13_u0_n99 ) );
  OAI211_X1 u1_u13_u0_U52 (.C2( u1_u13_u0_n140 ) , .C1( u1_u13_u0_n161 ) , .A( u1_u13_u0_n169 ) , .B( u1_u13_u0_n98 ) , .ZN( u1_u13_u0_n99 ) );
  AOI211_X1 u1_u13_u0_U53 (.C1( u1_u13_u0_n118 ) , .A( u1_u13_u0_n123 ) , .B( u1_u13_u0_n96 ) , .C2( u1_u13_u0_n97 ) , .ZN( u1_u13_u0_n98 ) );
  INV_X1 u1_u13_u0_U54 (.ZN( u1_u13_u0_n169 ) , .A( u1_u13_u0_n91 ) );
  NOR2_X1 u1_u13_u0_U55 (.A2( u1_u13_X_6 ) , .ZN( u1_u13_u0_n100 ) , .A1( u1_u13_u0_n162 ) );
  NOR2_X1 u1_u13_u0_U56 (.A2( u1_u13_X_4 ) , .A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n118 ) );
  NOR2_X1 u1_u13_u0_U57 (.A2( u1_u13_X_2 ) , .ZN( u1_u13_u0_n103 ) , .A1( u1_u13_u0_n164 ) );
  NOR2_X1 u1_u13_u0_U58 (.A2( u1_u13_X_1 ) , .A1( u1_u13_X_2 ) , .ZN( u1_u13_u0_n92 ) );
  NOR2_X1 u1_u13_u0_U59 (.A2( u1_u13_X_1 ) , .ZN( u1_u13_u0_n101 ) , .A1( u1_u13_u0_n163 ) );
  NOR2_X1 u1_u13_u0_U6 (.A1( u1_u13_u0_n108 ) , .ZN( u1_u13_u0_n123 ) , .A2( u1_u13_u0_n158 ) );
  NAND2_X1 u1_u13_u0_U60 (.A2( u1_u13_X_4 ) , .A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n144 ) );
  NOR2_X1 u1_u13_u0_U61 (.A2( u1_u13_X_5 ) , .ZN( u1_u13_u0_n136 ) , .A1( u1_u13_u0_n159 ) );
  NAND2_X1 u1_u13_u0_U62 (.A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n138 ) , .A2( u1_u13_u0_n159 ) );
  AND2_X1 u1_u13_u0_U63 (.A2( u1_u13_X_3 ) , .A1( u1_u13_X_6 ) , .ZN( u1_u13_u0_n102 ) );
  AND2_X1 u1_u13_u0_U64 (.A1( u1_u13_X_6 ) , .A2( u1_u13_u0_n162 ) , .ZN( u1_u13_u0_n93 ) );
  INV_X1 u1_u13_u0_U65 (.A( u1_u13_X_4 ) , .ZN( u1_u13_u0_n159 ) );
  INV_X1 u1_u13_u0_U66 (.A( u1_u13_X_1 ) , .ZN( u1_u13_u0_n164 ) );
  INV_X1 u1_u13_u0_U67 (.A( u1_u13_X_2 ) , .ZN( u1_u13_u0_n163 ) );
  INV_X1 u1_u13_u0_U68 (.A( u1_u13_u0_n126 ) , .ZN( u1_u13_u0_n168 ) );
  AOI211_X1 u1_u13_u0_U69 (.B( u1_u13_u0_n133 ) , .A( u1_u13_u0_n134 ) , .C2( u1_u13_u0_n135 ) , .C1( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n137 ) );
  OAI21_X1 u1_u13_u0_U7 (.B1( u1_u13_u0_n150 ) , .B2( u1_u13_u0_n158 ) , .A( u1_u13_u0_n172 ) , .ZN( u1_u13_u0_n89 ) );
  INV_X1 u1_u13_u0_U70 (.ZN( u1_u13_u0_n174 ) , .A( u1_u13_u0_n89 ) );
  AOI211_X1 u1_u13_u0_U71 (.B( u1_u13_u0_n104 ) , .A( u1_u13_u0_n105 ) , .ZN( u1_u13_u0_n106 ) , .C2( u1_u13_u0_n113 ) , .C1( u1_u13_u0_n160 ) );
  OR4_X1 u1_u13_u0_U72 (.ZN( u1_out13_17 ) , .A4( u1_u13_u0_n122 ) , .A2( u1_u13_u0_n123 ) , .A1( u1_u13_u0_n124 ) , .A3( u1_u13_u0_n170 ) );
  AOI21_X1 u1_u13_u0_U73 (.B2( u1_u13_u0_n107 ) , .ZN( u1_u13_u0_n124 ) , .B1( u1_u13_u0_n128 ) , .A( u1_u13_u0_n161 ) );
  INV_X1 u1_u13_u0_U74 (.A( u1_u13_u0_n111 ) , .ZN( u1_u13_u0_n170 ) );
  OR4_X1 u1_u13_u0_U75 (.ZN( u1_out13_31 ) , .A4( u1_u13_u0_n155 ) , .A2( u1_u13_u0_n156 ) , .A1( u1_u13_u0_n157 ) , .A3( u1_u13_u0_n173 ) );
  AOI21_X1 u1_u13_u0_U76 (.A( u1_u13_u0_n138 ) , .B2( u1_u13_u0_n139 ) , .B1( u1_u13_u0_n140 ) , .ZN( u1_u13_u0_n157 ) );
  AOI21_X1 u1_u13_u0_U77 (.B2( u1_u13_u0_n141 ) , .B1( u1_u13_u0_n142 ) , .ZN( u1_u13_u0_n156 ) , .A( u1_u13_u0_n161 ) );
  AOI21_X1 u1_u13_u0_U78 (.B1( u1_u13_u0_n132 ) , .ZN( u1_u13_u0_n133 ) , .A( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n166 ) );
  OAI22_X1 u1_u13_u0_U79 (.ZN( u1_u13_u0_n105 ) , .A2( u1_u13_u0_n132 ) , .B1( u1_u13_u0_n146 ) , .A1( u1_u13_u0_n147 ) , .B2( u1_u13_u0_n161 ) );
  AND2_X1 u1_u13_u0_U8 (.A1( u1_u13_u0_n114 ) , .A2( u1_u13_u0_n121 ) , .ZN( u1_u13_u0_n146 ) );
  NAND2_X1 u1_u13_u0_U80 (.ZN( u1_u13_u0_n110 ) , .A2( u1_u13_u0_n132 ) , .A1( u1_u13_u0_n145 ) );
  INV_X1 u1_u13_u0_U81 (.A( u1_u13_u0_n119 ) , .ZN( u1_u13_u0_n167 ) );
  NAND2_X1 u1_u13_u0_U82 (.A2( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n140 ) , .A1( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U83 (.A1( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n130 ) , .A2( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U84 (.ZN( u1_u13_u0_n108 ) , .A1( u1_u13_u0_n92 ) , .A2( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U85 (.ZN( u1_u13_u0_n142 ) , .A1( u1_u13_u0_n94 ) , .A2( u1_u13_u0_n95 ) );
  INV_X1 u1_u13_u0_U86 (.A( u1_u13_X_3 ) , .ZN( u1_u13_u0_n162 ) );
  NOR2_X1 u1_u13_u0_U87 (.A2( u1_u13_X_3 ) , .A1( u1_u13_X_6 ) , .ZN( u1_u13_u0_n94 ) );
  NAND3_X1 u1_u13_u0_U88 (.ZN( u1_out13_23 ) , .A3( u1_u13_u0_n137 ) , .A1( u1_u13_u0_n168 ) , .A2( u1_u13_u0_n171 ) );
  NAND3_X1 u1_u13_u0_U89 (.A3( u1_u13_u0_n127 ) , .A2( u1_u13_u0_n128 ) , .ZN( u1_u13_u0_n135 ) , .A1( u1_u13_u0_n150 ) );
  AND2_X1 u1_u13_u0_U9 (.A1( u1_u13_u0_n131 ) , .ZN( u1_u13_u0_n141 ) , .A2( u1_u13_u0_n150 ) );
  NAND3_X1 u1_u13_u0_U90 (.ZN( u1_u13_u0_n117 ) , .A3( u1_u13_u0_n132 ) , .A2( u1_u13_u0_n139 ) , .A1( u1_u13_u0_n148 ) );
  NAND3_X1 u1_u13_u0_U91 (.ZN( u1_u13_u0_n109 ) , .A2( u1_u13_u0_n114 ) , .A3( u1_u13_u0_n140 ) , .A1( u1_u13_u0_n149 ) );
  NAND3_X1 u1_u13_u0_U92 (.ZN( u1_out13_9 ) , .A3( u1_u13_u0_n106 ) , .A2( u1_u13_u0_n171 ) , .A1( u1_u13_u0_n174 ) );
  NAND3_X1 u1_u13_u0_U93 (.A2( u1_u13_u0_n128 ) , .A1( u1_u13_u0_n132 ) , .A3( u1_u13_u0_n146 ) , .ZN( u1_u13_u0_n97 ) );
  OAI22_X1 u1_u13_u2_U10 (.B1( u1_u13_u2_n151 ) , .A2( u1_u13_u2_n152 ) , .A1( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n160 ) , .B2( u1_u13_u2_n168 ) );
  NAND3_X1 u1_u13_u2_U100 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n104 ) , .A3( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n98 ) );
  NOR3_X1 u1_u13_u2_U11 (.A1( u1_u13_u2_n150 ) , .ZN( u1_u13_u2_n151 ) , .A3( u1_u13_u2_n175 ) , .A2( u1_u13_u2_n188 ) );
  AOI21_X1 u1_u13_u2_U12 (.B2( u1_u13_u2_n123 ) , .ZN( u1_u13_u2_n125 ) , .A( u1_u13_u2_n171 ) , .B1( u1_u13_u2_n184 ) );
  INV_X1 u1_u13_u2_U13 (.A( u1_u13_u2_n150 ) , .ZN( u1_u13_u2_n184 ) );
  AOI21_X1 u1_u13_u2_U14 (.ZN( u1_u13_u2_n144 ) , .B2( u1_u13_u2_n155 ) , .A( u1_u13_u2_n172 ) , .B1( u1_u13_u2_n185 ) );
  AOI21_X1 u1_u13_u2_U15 (.B2( u1_u13_u2_n143 ) , .ZN( u1_u13_u2_n145 ) , .B1( u1_u13_u2_n152 ) , .A( u1_u13_u2_n171 ) );
  INV_X1 u1_u13_u2_U16 (.A( u1_u13_u2_n156 ) , .ZN( u1_u13_u2_n171 ) );
  INV_X1 u1_u13_u2_U17 (.A( u1_u13_u2_n120 ) , .ZN( u1_u13_u2_n188 ) );
  NAND2_X1 u1_u13_u2_U18 (.A2( u1_u13_u2_n122 ) , .ZN( u1_u13_u2_n150 ) , .A1( u1_u13_u2_n152 ) );
  INV_X1 u1_u13_u2_U19 (.A( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n170 ) );
  INV_X1 u1_u13_u2_U20 (.A( u1_u13_u2_n137 ) , .ZN( u1_u13_u2_n173 ) );
  NAND2_X1 u1_u13_u2_U21 (.A1( u1_u13_u2_n132 ) , .A2( u1_u13_u2_n139 ) , .ZN( u1_u13_u2_n157 ) );
  INV_X1 u1_u13_u2_U22 (.A( u1_u13_u2_n113 ) , .ZN( u1_u13_u2_n178 ) );
  INV_X1 u1_u13_u2_U23 (.A( u1_u13_u2_n139 ) , .ZN( u1_u13_u2_n175 ) );
  INV_X1 u1_u13_u2_U24 (.A( u1_u13_u2_n155 ) , .ZN( u1_u13_u2_n181 ) );
  INV_X1 u1_u13_u2_U25 (.A( u1_u13_u2_n119 ) , .ZN( u1_u13_u2_n177 ) );
  INV_X1 u1_u13_u2_U26 (.A( u1_u13_u2_n116 ) , .ZN( u1_u13_u2_n180 ) );
  INV_X1 u1_u13_u2_U27 (.A( u1_u13_u2_n131 ) , .ZN( u1_u13_u2_n179 ) );
  INV_X1 u1_u13_u2_U28 (.A( u1_u13_u2_n154 ) , .ZN( u1_u13_u2_n176 ) );
  NAND2_X1 u1_u13_u2_U29 (.A2( u1_u13_u2_n116 ) , .A1( u1_u13_u2_n117 ) , .ZN( u1_u13_u2_n118 ) );
  NOR2_X1 u1_u13_u2_U3 (.ZN( u1_u13_u2_n121 ) , .A2( u1_u13_u2_n177 ) , .A1( u1_u13_u2_n180 ) );
  INV_X1 u1_u13_u2_U30 (.A( u1_u13_u2_n132 ) , .ZN( u1_u13_u2_n182 ) );
  INV_X1 u1_u13_u2_U31 (.A( u1_u13_u2_n158 ) , .ZN( u1_u13_u2_n183 ) );
  OAI21_X1 u1_u13_u2_U32 (.A( u1_u13_u2_n156 ) , .B1( u1_u13_u2_n157 ) , .ZN( u1_u13_u2_n158 ) , .B2( u1_u13_u2_n179 ) );
  NOR2_X1 u1_u13_u2_U33 (.ZN( u1_u13_u2_n156 ) , .A1( u1_u13_u2_n166 ) , .A2( u1_u13_u2_n169 ) );
  NOR2_X1 u1_u13_u2_U34 (.A2( u1_u13_u2_n114 ) , .ZN( u1_u13_u2_n137 ) , .A1( u1_u13_u2_n140 ) );
  NOR2_X1 u1_u13_u2_U35 (.A2( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n153 ) , .A1( u1_u13_u2_n156 ) );
  AOI211_X1 u1_u13_u2_U36 (.ZN( u1_u13_u2_n130 ) , .C1( u1_u13_u2_n138 ) , .C2( u1_u13_u2_n179 ) , .B( u1_u13_u2_n96 ) , .A( u1_u13_u2_n97 ) );
  OAI22_X1 u1_u13_u2_U37 (.B1( u1_u13_u2_n133 ) , .A2( u1_u13_u2_n137 ) , .A1( u1_u13_u2_n152 ) , .B2( u1_u13_u2_n168 ) , .ZN( u1_u13_u2_n97 ) );
  OAI221_X1 u1_u13_u2_U38 (.B1( u1_u13_u2_n113 ) , .C1( u1_u13_u2_n132 ) , .A( u1_u13_u2_n149 ) , .B2( u1_u13_u2_n171 ) , .C2( u1_u13_u2_n172 ) , .ZN( u1_u13_u2_n96 ) );
  OAI221_X1 u1_u13_u2_U39 (.A( u1_u13_u2_n115 ) , .C2( u1_u13_u2_n123 ) , .B2( u1_u13_u2_n143 ) , .B1( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n163 ) , .C1( u1_u13_u2_n168 ) );
  INV_X1 u1_u13_u2_U4 (.A( u1_u13_u2_n134 ) , .ZN( u1_u13_u2_n185 ) );
  OAI21_X1 u1_u13_u2_U40 (.A( u1_u13_u2_n114 ) , .ZN( u1_u13_u2_n115 ) , .B1( u1_u13_u2_n176 ) , .B2( u1_u13_u2_n178 ) );
  OAI221_X1 u1_u13_u2_U41 (.A( u1_u13_u2_n135 ) , .B2( u1_u13_u2_n136 ) , .B1( u1_u13_u2_n137 ) , .ZN( u1_u13_u2_n162 ) , .C2( u1_u13_u2_n167 ) , .C1( u1_u13_u2_n185 ) );
  AND3_X1 u1_u13_u2_U42 (.A3( u1_u13_u2_n131 ) , .A2( u1_u13_u2_n132 ) , .A1( u1_u13_u2_n133 ) , .ZN( u1_u13_u2_n136 ) );
  AOI22_X1 u1_u13_u2_U43 (.ZN( u1_u13_u2_n135 ) , .B1( u1_u13_u2_n140 ) , .A1( u1_u13_u2_n156 ) , .B2( u1_u13_u2_n180 ) , .A2( u1_u13_u2_n188 ) );
  AOI21_X1 u1_u13_u2_U44 (.ZN( u1_u13_u2_n149 ) , .B1( u1_u13_u2_n173 ) , .B2( u1_u13_u2_n188 ) , .A( u1_u13_u2_n95 ) );
  AND3_X1 u1_u13_u2_U45 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n104 ) , .A3( u1_u13_u2_n156 ) , .ZN( u1_u13_u2_n95 ) );
  OAI21_X1 u1_u13_u2_U46 (.A( u1_u13_u2_n101 ) , .B2( u1_u13_u2_n121 ) , .B1( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n164 ) );
  NAND2_X1 u1_u13_u2_U47 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n107 ) , .ZN( u1_u13_u2_n155 ) );
  NAND2_X1 u1_u13_u2_U48 (.A2( u1_u13_u2_n105 ) , .A1( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n143 ) );
  NAND2_X1 u1_u13_u2_U49 (.A1( u1_u13_u2_n104 ) , .A2( u1_u13_u2_n106 ) , .ZN( u1_u13_u2_n152 ) );
  NOR4_X1 u1_u13_u2_U5 (.A4( u1_u13_u2_n124 ) , .A3( u1_u13_u2_n125 ) , .A2( u1_u13_u2_n126 ) , .A1( u1_u13_u2_n127 ) , .ZN( u1_u13_u2_n128 ) );
  NAND2_X1 u1_u13_u2_U50 (.A1( u1_u13_u2_n100 ) , .A2( u1_u13_u2_n105 ) , .ZN( u1_u13_u2_n132 ) );
  INV_X1 u1_u13_u2_U51 (.A( u1_u13_u2_n140 ) , .ZN( u1_u13_u2_n168 ) );
  INV_X1 u1_u13_u2_U52 (.A( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n167 ) );
  OAI21_X1 u1_u13_u2_U53 (.A( u1_u13_u2_n141 ) , .B2( u1_u13_u2_n142 ) , .ZN( u1_u13_u2_n146 ) , .B1( u1_u13_u2_n153 ) );
  OAI21_X1 u1_u13_u2_U54 (.A( u1_u13_u2_n140 ) , .ZN( u1_u13_u2_n141 ) , .B1( u1_u13_u2_n176 ) , .B2( u1_u13_u2_n177 ) );
  NOR3_X1 u1_u13_u2_U55 (.ZN( u1_u13_u2_n142 ) , .A3( u1_u13_u2_n175 ) , .A2( u1_u13_u2_n178 ) , .A1( u1_u13_u2_n181 ) );
  NAND2_X1 u1_u13_u2_U56 (.A1( u1_u13_u2_n102 ) , .A2( u1_u13_u2_n106 ) , .ZN( u1_u13_u2_n113 ) );
  NAND2_X1 u1_u13_u2_U57 (.A1( u1_u13_u2_n106 ) , .A2( u1_u13_u2_n107 ) , .ZN( u1_u13_u2_n131 ) );
  NAND2_X1 u1_u13_u2_U58 (.A1( u1_u13_u2_n103 ) , .A2( u1_u13_u2_n107 ) , .ZN( u1_u13_u2_n139 ) );
  NAND2_X1 u1_u13_u2_U59 (.A1( u1_u13_u2_n103 ) , .A2( u1_u13_u2_n105 ) , .ZN( u1_u13_u2_n133 ) );
  AOI21_X1 u1_u13_u2_U6 (.B2( u1_u13_u2_n119 ) , .ZN( u1_u13_u2_n127 ) , .A( u1_u13_u2_n137 ) , .B1( u1_u13_u2_n155 ) );
  NAND2_X1 u1_u13_u2_U60 (.A1( u1_u13_u2_n102 ) , .A2( u1_u13_u2_n103 ) , .ZN( u1_u13_u2_n154 ) );
  NAND2_X1 u1_u13_u2_U61 (.A2( u1_u13_u2_n103 ) , .A1( u1_u13_u2_n104 ) , .ZN( u1_u13_u2_n119 ) );
  NAND2_X1 u1_u13_u2_U62 (.A2( u1_u13_u2_n107 ) , .A1( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n123 ) );
  NAND2_X1 u1_u13_u2_U63 (.A1( u1_u13_u2_n104 ) , .A2( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n122 ) );
  INV_X1 u1_u13_u2_U64 (.A( u1_u13_u2_n114 ) , .ZN( u1_u13_u2_n172 ) );
  NAND2_X1 u1_u13_u2_U65 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n102 ) , .ZN( u1_u13_u2_n116 ) );
  NAND2_X1 u1_u13_u2_U66 (.A1( u1_u13_u2_n102 ) , .A2( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n120 ) );
  NAND2_X1 u1_u13_u2_U67 (.A2( u1_u13_u2_n105 ) , .A1( u1_u13_u2_n106 ) , .ZN( u1_u13_u2_n117 ) );
  INV_X1 u1_u13_u2_U68 (.ZN( u1_u13_u2_n187 ) , .A( u1_u13_u2_n99 ) );
  OAI21_X1 u1_u13_u2_U69 (.B1( u1_u13_u2_n137 ) , .B2( u1_u13_u2_n143 ) , .A( u1_u13_u2_n98 ) , .ZN( u1_u13_u2_n99 ) );
  AOI21_X1 u1_u13_u2_U7 (.ZN( u1_u13_u2_n124 ) , .B1( u1_u13_u2_n131 ) , .B2( u1_u13_u2_n143 ) , .A( u1_u13_u2_n172 ) );
  NOR2_X1 u1_u13_u2_U70 (.A2( u1_u13_X_16 ) , .ZN( u1_u13_u2_n140 ) , .A1( u1_u13_u2_n166 ) );
  NOR2_X1 u1_u13_u2_U71 (.A2( u1_u13_X_13 ) , .A1( u1_u13_X_14 ) , .ZN( u1_u13_u2_n100 ) );
  NOR2_X1 u1_u13_u2_U72 (.A2( u1_u13_X_16 ) , .A1( u1_u13_X_17 ) , .ZN( u1_u13_u2_n138 ) );
  NOR2_X1 u1_u13_u2_U73 (.A2( u1_u13_X_15 ) , .A1( u1_u13_X_18 ) , .ZN( u1_u13_u2_n104 ) );
  NOR2_X1 u1_u13_u2_U74 (.A2( u1_u13_X_14 ) , .ZN( u1_u13_u2_n103 ) , .A1( u1_u13_u2_n174 ) );
  NOR2_X1 u1_u13_u2_U75 (.A2( u1_u13_X_15 ) , .ZN( u1_u13_u2_n102 ) , .A1( u1_u13_u2_n165 ) );
  NOR2_X1 u1_u13_u2_U76 (.A2( u1_u13_X_17 ) , .ZN( u1_u13_u2_n114 ) , .A1( u1_u13_u2_n169 ) );
  AND2_X1 u1_u13_u2_U77 (.A1( u1_u13_X_15 ) , .ZN( u1_u13_u2_n105 ) , .A2( u1_u13_u2_n165 ) );
  AND2_X1 u1_u13_u2_U78 (.A2( u1_u13_X_15 ) , .A1( u1_u13_X_18 ) , .ZN( u1_u13_u2_n107 ) );
  AND2_X1 u1_u13_u2_U79 (.A1( u1_u13_X_14 ) , .ZN( u1_u13_u2_n106 ) , .A2( u1_u13_u2_n174 ) );
  AOI21_X1 u1_u13_u2_U8 (.B2( u1_u13_u2_n120 ) , .B1( u1_u13_u2_n121 ) , .ZN( u1_u13_u2_n126 ) , .A( u1_u13_u2_n167 ) );
  AND2_X1 u1_u13_u2_U80 (.A1( u1_u13_X_13 ) , .A2( u1_u13_X_14 ) , .ZN( u1_u13_u2_n108 ) );
  INV_X1 u1_u13_u2_U81 (.A( u1_u13_X_16 ) , .ZN( u1_u13_u2_n169 ) );
  INV_X1 u1_u13_u2_U82 (.A( u1_u13_X_17 ) , .ZN( u1_u13_u2_n166 ) );
  INV_X1 u1_u13_u2_U83 (.A( u1_u13_X_13 ) , .ZN( u1_u13_u2_n174 ) );
  INV_X1 u1_u13_u2_U84 (.A( u1_u13_X_18 ) , .ZN( u1_u13_u2_n165 ) );
  NAND4_X1 u1_u13_u2_U85 (.ZN( u1_out13_30 ) , .A4( u1_u13_u2_n147 ) , .A3( u1_u13_u2_n148 ) , .A2( u1_u13_u2_n149 ) , .A1( u1_u13_u2_n187 ) );
  NOR3_X1 u1_u13_u2_U86 (.A3( u1_u13_u2_n144 ) , .A2( u1_u13_u2_n145 ) , .A1( u1_u13_u2_n146 ) , .ZN( u1_u13_u2_n147 ) );
  AOI21_X1 u1_u13_u2_U87 (.B2( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n148 ) , .A( u1_u13_u2_n162 ) , .B1( u1_u13_u2_n182 ) );
  NAND4_X1 u1_u13_u2_U88 (.ZN( u1_out13_24 ) , .A4( u1_u13_u2_n111 ) , .A3( u1_u13_u2_n112 ) , .A1( u1_u13_u2_n130 ) , .A2( u1_u13_u2_n187 ) );
  AOI221_X1 u1_u13_u2_U89 (.A( u1_u13_u2_n109 ) , .B1( u1_u13_u2_n110 ) , .ZN( u1_u13_u2_n111 ) , .C1( u1_u13_u2_n134 ) , .C2( u1_u13_u2_n170 ) , .B2( u1_u13_u2_n173 ) );
  OAI22_X1 u1_u13_u2_U9 (.ZN( u1_u13_u2_n109 ) , .A2( u1_u13_u2_n113 ) , .B2( u1_u13_u2_n133 ) , .B1( u1_u13_u2_n167 ) , .A1( u1_u13_u2_n168 ) );
  AOI21_X1 u1_u13_u2_U90 (.ZN( u1_u13_u2_n112 ) , .B2( u1_u13_u2_n156 ) , .A( u1_u13_u2_n164 ) , .B1( u1_u13_u2_n181 ) );
  NAND4_X1 u1_u13_u2_U91 (.ZN( u1_out13_16 ) , .A4( u1_u13_u2_n128 ) , .A3( u1_u13_u2_n129 ) , .A1( u1_u13_u2_n130 ) , .A2( u1_u13_u2_n186 ) );
  AOI22_X1 u1_u13_u2_U92 (.A2( u1_u13_u2_n118 ) , .ZN( u1_u13_u2_n129 ) , .A1( u1_u13_u2_n140 ) , .B1( u1_u13_u2_n157 ) , .B2( u1_u13_u2_n170 ) );
  INV_X1 u1_u13_u2_U93 (.A( u1_u13_u2_n163 ) , .ZN( u1_u13_u2_n186 ) );
  OR4_X1 u1_u13_u2_U94 (.ZN( u1_out13_6 ) , .A4( u1_u13_u2_n161 ) , .A3( u1_u13_u2_n162 ) , .A2( u1_u13_u2_n163 ) , .A1( u1_u13_u2_n164 ) );
  OR3_X1 u1_u13_u2_U95 (.A2( u1_u13_u2_n159 ) , .A1( u1_u13_u2_n160 ) , .ZN( u1_u13_u2_n161 ) , .A3( u1_u13_u2_n183 ) );
  AOI21_X1 u1_u13_u2_U96 (.B2( u1_u13_u2_n154 ) , .B1( u1_u13_u2_n155 ) , .ZN( u1_u13_u2_n159 ) , .A( u1_u13_u2_n167 ) );
  NAND3_X1 u1_u13_u2_U97 (.A2( u1_u13_u2_n117 ) , .A1( u1_u13_u2_n122 ) , .A3( u1_u13_u2_n123 ) , .ZN( u1_u13_u2_n134 ) );
  NAND3_X1 u1_u13_u2_U98 (.ZN( u1_u13_u2_n110 ) , .A2( u1_u13_u2_n131 ) , .A3( u1_u13_u2_n139 ) , .A1( u1_u13_u2_n154 ) );
  NAND3_X1 u1_u13_u2_U99 (.A2( u1_u13_u2_n100 ) , .ZN( u1_u13_u2_n101 ) , .A1( u1_u13_u2_n104 ) , .A3( u1_u13_u2_n114 ) );
  XOR2_X1 u1_u14_U1 (.B( u1_K15_9 ) , .A( u1_R13_6 ) , .Z( u1_u14_X_9 ) );
  XOR2_X1 u1_u14_U48 (.B( u1_K15_10 ) , .A( u1_R13_7 ) , .Z( u1_u14_X_10 ) );
  AOI21_X1 u1_u14_u1_U10 (.ZN( u1_u14_u1_n106 ) , .A( u1_u14_u1_n112 ) , .B1( u1_u14_u1_n154 ) , .B2( u1_u14_u1_n156 ) );
  NAND3_X1 u1_u14_u1_U100 (.ZN( u1_u14_u1_n113 ) , .A1( u1_u14_u1_n120 ) , .A3( u1_u14_u1_n133 ) , .A2( u1_u14_u1_n155 ) );
  INV_X1 u1_u14_u1_U11 (.A( u1_u14_u1_n101 ) , .ZN( u1_u14_u1_n184 ) );
  AOI21_X1 u1_u14_u1_U12 (.ZN( u1_u14_u1_n107 ) , .B1( u1_u14_u1_n134 ) , .B2( u1_u14_u1_n149 ) , .A( u1_u14_u1_n174 ) );
  NAND2_X1 u1_u14_u1_U13 (.ZN( u1_u14_u1_n140 ) , .A2( u1_u14_u1_n150 ) , .A1( u1_u14_u1_n155 ) );
  NAND2_X1 u1_u14_u1_U14 (.A1( u1_u14_u1_n131 ) , .ZN( u1_u14_u1_n147 ) , .A2( u1_u14_u1_n153 ) );
  AOI22_X1 u1_u14_u1_U15 (.B2( u1_u14_u1_n136 ) , .A2( u1_u14_u1_n137 ) , .ZN( u1_u14_u1_n143 ) , .A1( u1_u14_u1_n171 ) , .B1( u1_u14_u1_n173 ) );
  INV_X1 u1_u14_u1_U16 (.A( u1_u14_u1_n147 ) , .ZN( u1_u14_u1_n181 ) );
  INV_X1 u1_u14_u1_U17 (.A( u1_u14_u1_n139 ) , .ZN( u1_u14_u1_n174 ) );
  INV_X1 u1_u14_u1_U18 (.A( u1_u14_u1_n112 ) , .ZN( u1_u14_u1_n171 ) );
  NAND2_X1 u1_u14_u1_U19 (.ZN( u1_u14_u1_n141 ) , .A1( u1_u14_u1_n153 ) , .A2( u1_u14_u1_n156 ) );
  AND2_X1 u1_u14_u1_U20 (.A1( u1_u14_u1_n123 ) , .ZN( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n161 ) );
  NAND2_X1 u1_u14_u1_U21 (.A2( u1_u14_u1_n115 ) , .A1( u1_u14_u1_n116 ) , .ZN( u1_u14_u1_n148 ) );
  NAND2_X1 u1_u14_u1_U22 (.A2( u1_u14_u1_n133 ) , .A1( u1_u14_u1_n135 ) , .ZN( u1_u14_u1_n159 ) );
  NAND2_X1 u1_u14_u1_U23 (.A2( u1_u14_u1_n115 ) , .A1( u1_u14_u1_n120 ) , .ZN( u1_u14_u1_n132 ) );
  INV_X1 u1_u14_u1_U24 (.A( u1_u14_u1_n154 ) , .ZN( u1_u14_u1_n178 ) );
  AOI22_X1 u1_u14_u1_U25 (.B2( u1_u14_u1_n113 ) , .A2( u1_u14_u1_n114 ) , .ZN( u1_u14_u1_n125 ) , .A1( u1_u14_u1_n171 ) , .B1( u1_u14_u1_n173 ) );
  NAND2_X1 u1_u14_u1_U26 (.ZN( u1_u14_u1_n114 ) , .A1( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n156 ) );
  INV_X1 u1_u14_u1_U27 (.A( u1_u14_u1_n151 ) , .ZN( u1_u14_u1_n183 ) );
  AND2_X1 u1_u14_u1_U28 (.A1( u1_u14_u1_n129 ) , .A2( u1_u14_u1_n133 ) , .ZN( u1_u14_u1_n149 ) );
  INV_X1 u1_u14_u1_U29 (.A( u1_u14_u1_n131 ) , .ZN( u1_u14_u1_n180 ) );
  INV_X1 u1_u14_u1_U3 (.A( u1_u14_u1_n159 ) , .ZN( u1_u14_u1_n182 ) );
  AOI221_X1 u1_u14_u1_U30 (.B1( u1_u14_u1_n140 ) , .ZN( u1_u14_u1_n167 ) , .B2( u1_u14_u1_n172 ) , .C2( u1_u14_u1_n175 ) , .C1( u1_u14_u1_n178 ) , .A( u1_u14_u1_n188 ) );
  INV_X1 u1_u14_u1_U31 (.ZN( u1_u14_u1_n188 ) , .A( u1_u14_u1_n97 ) );
  AOI211_X1 u1_u14_u1_U32 (.A( u1_u14_u1_n118 ) , .C1( u1_u14_u1_n132 ) , .C2( u1_u14_u1_n139 ) , .B( u1_u14_u1_n96 ) , .ZN( u1_u14_u1_n97 ) );
  AOI21_X1 u1_u14_u1_U33 (.B2( u1_u14_u1_n121 ) , .B1( u1_u14_u1_n135 ) , .A( u1_u14_u1_n152 ) , .ZN( u1_u14_u1_n96 ) );
  OAI221_X1 u1_u14_u1_U34 (.A( u1_u14_u1_n119 ) , .C2( u1_u14_u1_n129 ) , .ZN( u1_u14_u1_n138 ) , .B2( u1_u14_u1_n152 ) , .C1( u1_u14_u1_n174 ) , .B1( u1_u14_u1_n187 ) );
  INV_X1 u1_u14_u1_U35 (.A( u1_u14_u1_n148 ) , .ZN( u1_u14_u1_n187 ) );
  AOI211_X1 u1_u14_u1_U36 (.B( u1_u14_u1_n117 ) , .A( u1_u14_u1_n118 ) , .ZN( u1_u14_u1_n119 ) , .C2( u1_u14_u1_n146 ) , .C1( u1_u14_u1_n159 ) );
  NOR2_X1 u1_u14_u1_U37 (.A1( u1_u14_u1_n168 ) , .A2( u1_u14_u1_n176 ) , .ZN( u1_u14_u1_n98 ) );
  AOI211_X1 u1_u14_u1_U38 (.B( u1_u14_u1_n162 ) , .A( u1_u14_u1_n163 ) , .C2( u1_u14_u1_n164 ) , .ZN( u1_u14_u1_n165 ) , .C1( u1_u14_u1_n171 ) );
  AOI21_X1 u1_u14_u1_U39 (.A( u1_u14_u1_n160 ) , .B2( u1_u14_u1_n161 ) , .ZN( u1_u14_u1_n162 ) , .B1( u1_u14_u1_n182 ) );
  AOI221_X1 u1_u14_u1_U4 (.A( u1_u14_u1_n138 ) , .C2( u1_u14_u1_n139 ) , .C1( u1_u14_u1_n140 ) , .B2( u1_u14_u1_n141 ) , .ZN( u1_u14_u1_n142 ) , .B1( u1_u14_u1_n175 ) );
  OR2_X1 u1_u14_u1_U40 (.A2( u1_u14_u1_n157 ) , .A1( u1_u14_u1_n158 ) , .ZN( u1_u14_u1_n163 ) );
  OAI21_X1 u1_u14_u1_U41 (.B2( u1_u14_u1_n123 ) , .ZN( u1_u14_u1_n145 ) , .B1( u1_u14_u1_n160 ) , .A( u1_u14_u1_n185 ) );
  INV_X1 u1_u14_u1_U42 (.A( u1_u14_u1_n122 ) , .ZN( u1_u14_u1_n185 ) );
  AOI21_X1 u1_u14_u1_U43 (.B2( u1_u14_u1_n120 ) , .B1( u1_u14_u1_n121 ) , .ZN( u1_u14_u1_n122 ) , .A( u1_u14_u1_n128 ) );
  NAND2_X1 u1_u14_u1_U44 (.A1( u1_u14_u1_n128 ) , .ZN( u1_u14_u1_n146 ) , .A2( u1_u14_u1_n160 ) );
  NAND2_X1 u1_u14_u1_U45 (.A2( u1_u14_u1_n112 ) , .ZN( u1_u14_u1_n139 ) , .A1( u1_u14_u1_n152 ) );
  NAND2_X1 u1_u14_u1_U46 (.A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n156 ) , .A2( u1_u14_u1_n99 ) );
  NOR2_X1 u1_u14_u1_U47 (.ZN( u1_u14_u1_n117 ) , .A1( u1_u14_u1_n121 ) , .A2( u1_u14_u1_n160 ) );
  AOI21_X1 u1_u14_u1_U48 (.A( u1_u14_u1_n128 ) , .B2( u1_u14_u1_n129 ) , .ZN( u1_u14_u1_n130 ) , .B1( u1_u14_u1_n150 ) );
  NAND2_X1 u1_u14_u1_U49 (.ZN( u1_u14_u1_n112 ) , .A1( u1_u14_u1_n169 ) , .A2( u1_u14_u1_n170 ) );
  AOI211_X1 u1_u14_u1_U5 (.ZN( u1_u14_u1_n124 ) , .A( u1_u14_u1_n138 ) , .C2( u1_u14_u1_n139 ) , .B( u1_u14_u1_n145 ) , .C1( u1_u14_u1_n147 ) );
  NAND2_X1 u1_u14_u1_U50 (.ZN( u1_u14_u1_n129 ) , .A2( u1_u14_u1_n95 ) , .A1( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U51 (.A1( u1_u14_u1_n102 ) , .ZN( u1_u14_u1_n154 ) , .A2( u1_u14_u1_n99 ) );
  NAND2_X1 u1_u14_u1_U52 (.A2( u1_u14_u1_n100 ) , .ZN( u1_u14_u1_n135 ) , .A1( u1_u14_u1_n99 ) );
  AOI21_X1 u1_u14_u1_U53 (.A( u1_u14_u1_n152 ) , .B2( u1_u14_u1_n153 ) , .B1( u1_u14_u1_n154 ) , .ZN( u1_u14_u1_n158 ) );
  INV_X1 u1_u14_u1_U54 (.A( u1_u14_u1_n160 ) , .ZN( u1_u14_u1_n175 ) );
  NAND2_X1 u1_u14_u1_U55 (.A1( u1_u14_u1_n100 ) , .ZN( u1_u14_u1_n116 ) , .A2( u1_u14_u1_n95 ) );
  NAND2_X1 u1_u14_u1_U56 (.A1( u1_u14_u1_n102 ) , .ZN( u1_u14_u1_n131 ) , .A2( u1_u14_u1_n95 ) );
  NAND2_X1 u1_u14_u1_U57 (.A2( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n121 ) , .A1( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U58 (.A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n153 ) , .A2( u1_u14_u1_n98 ) );
  NAND2_X1 u1_u14_u1_U59 (.A2( u1_u14_u1_n104 ) , .A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n133 ) );
  NOR2_X1 u1_u14_u1_U6 (.A1( u1_u14_u1_n112 ) , .A2( u1_u14_u1_n116 ) , .ZN( u1_u14_u1_n118 ) );
  NAND2_X1 u1_u14_u1_U60 (.ZN( u1_u14_u1_n150 ) , .A2( u1_u14_u1_n98 ) , .A1( u1_u14_u1_n99 ) );
  NAND2_X1 u1_u14_u1_U61 (.A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n155 ) , .A2( u1_u14_u1_n95 ) );
  OAI21_X1 u1_u14_u1_U62 (.ZN( u1_u14_u1_n109 ) , .B1( u1_u14_u1_n129 ) , .B2( u1_u14_u1_n160 ) , .A( u1_u14_u1_n167 ) );
  NAND2_X1 u1_u14_u1_U63 (.A2( u1_u14_u1_n100 ) , .A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n120 ) );
  NAND2_X1 u1_u14_u1_U64 (.A1( u1_u14_u1_n102 ) , .A2( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n115 ) );
  NAND2_X1 u1_u14_u1_U65 (.A2( u1_u14_u1_n100 ) , .A1( u1_u14_u1_n104 ) , .ZN( u1_u14_u1_n151 ) );
  NAND2_X1 u1_u14_u1_U66 (.A2( u1_u14_u1_n103 ) , .A1( u1_u14_u1_n105 ) , .ZN( u1_u14_u1_n161 ) );
  INV_X1 u1_u14_u1_U67 (.A( u1_u14_u1_n152 ) , .ZN( u1_u14_u1_n173 ) );
  INV_X1 u1_u14_u1_U68 (.A( u1_u14_u1_n128 ) , .ZN( u1_u14_u1_n172 ) );
  NAND2_X1 u1_u14_u1_U69 (.A2( u1_u14_u1_n102 ) , .A1( u1_u14_u1_n103 ) , .ZN( u1_u14_u1_n123 ) );
  OAI21_X1 u1_u14_u1_U7 (.ZN( u1_u14_u1_n101 ) , .B1( u1_u14_u1_n141 ) , .A( u1_u14_u1_n146 ) , .B2( u1_u14_u1_n183 ) );
  NOR2_X1 u1_u14_u1_U70 (.A2( u1_u14_X_7 ) , .A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n95 ) );
  NOR2_X1 u1_u14_u1_U71 (.A1( u1_u14_X_12 ) , .A2( u1_u14_X_9 ) , .ZN( u1_u14_u1_n100 ) );
  NOR2_X1 u1_u14_u1_U72 (.A2( u1_u14_X_8 ) , .A1( u1_u14_u1_n177 ) , .ZN( u1_u14_u1_n99 ) );
  NOR2_X1 u1_u14_u1_U73 (.A2( u1_u14_X_12 ) , .ZN( u1_u14_u1_n102 ) , .A1( u1_u14_u1_n176 ) );
  NOR2_X1 u1_u14_u1_U74 (.A2( u1_u14_X_9 ) , .ZN( u1_u14_u1_n105 ) , .A1( u1_u14_u1_n168 ) );
  NAND2_X1 u1_u14_u1_U75 (.A1( u1_u14_X_10 ) , .ZN( u1_u14_u1_n160 ) , .A2( u1_u14_u1_n169 ) );
  NAND2_X1 u1_u14_u1_U76 (.A2( u1_u14_X_10 ) , .A1( u1_u14_X_11 ) , .ZN( u1_u14_u1_n152 ) );
  NAND2_X1 u1_u14_u1_U77 (.A1( u1_u14_X_11 ) , .ZN( u1_u14_u1_n128 ) , .A2( u1_u14_u1_n170 ) );
  AND2_X1 u1_u14_u1_U78 (.A2( u1_u14_X_7 ) , .A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n104 ) );
  AND2_X1 u1_u14_u1_U79 (.A1( u1_u14_X_8 ) , .ZN( u1_u14_u1_n103 ) , .A2( u1_u14_u1_n177 ) );
  AOI21_X1 u1_u14_u1_U8 (.B2( u1_u14_u1_n155 ) , .B1( u1_u14_u1_n156 ) , .ZN( u1_u14_u1_n157 ) , .A( u1_u14_u1_n174 ) );
  INV_X1 u1_u14_u1_U80 (.A( u1_u14_X_10 ) , .ZN( u1_u14_u1_n170 ) );
  INV_X1 u1_u14_u1_U81 (.A( u1_u14_X_9 ) , .ZN( u1_u14_u1_n176 ) );
  INV_X1 u1_u14_u1_U82 (.A( u1_u14_X_11 ) , .ZN( u1_u14_u1_n169 ) );
  INV_X1 u1_u14_u1_U83 (.A( u1_u14_X_12 ) , .ZN( u1_u14_u1_n168 ) );
  INV_X1 u1_u14_u1_U84 (.A( u1_u14_X_7 ) , .ZN( u1_u14_u1_n177 ) );
  NAND4_X1 u1_u14_u1_U85 (.ZN( u1_out14_18 ) , .A4( u1_u14_u1_n165 ) , .A3( u1_u14_u1_n166 ) , .A1( u1_u14_u1_n167 ) , .A2( u1_u14_u1_n186 ) );
  AOI22_X1 u1_u14_u1_U86 (.B2( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n147 ) , .A2( u1_u14_u1_n148 ) , .ZN( u1_u14_u1_n166 ) , .A1( u1_u14_u1_n172 ) );
  INV_X1 u1_u14_u1_U87 (.A( u1_u14_u1_n145 ) , .ZN( u1_u14_u1_n186 ) );
  OR4_X1 u1_u14_u1_U88 (.ZN( u1_out14_13 ) , .A4( u1_u14_u1_n108 ) , .A3( u1_u14_u1_n109 ) , .A2( u1_u14_u1_n110 ) , .A1( u1_u14_u1_n111 ) );
  AOI21_X1 u1_u14_u1_U89 (.ZN( u1_u14_u1_n111 ) , .A( u1_u14_u1_n128 ) , .B2( u1_u14_u1_n131 ) , .B1( u1_u14_u1_n135 ) );
  OR4_X1 u1_u14_u1_U9 (.A4( u1_u14_u1_n106 ) , .A3( u1_u14_u1_n107 ) , .ZN( u1_u14_u1_n108 ) , .A1( u1_u14_u1_n117 ) , .A2( u1_u14_u1_n184 ) );
  AOI21_X1 u1_u14_u1_U90 (.ZN( u1_u14_u1_n110 ) , .A( u1_u14_u1_n116 ) , .B1( u1_u14_u1_n152 ) , .B2( u1_u14_u1_n160 ) );
  NAND4_X1 u1_u14_u1_U91 (.ZN( u1_out14_2 ) , .A4( u1_u14_u1_n142 ) , .A3( u1_u14_u1_n143 ) , .A2( u1_u14_u1_n144 ) , .A1( u1_u14_u1_n179 ) );
  OAI21_X1 u1_u14_u1_U92 (.B2( u1_u14_u1_n132 ) , .ZN( u1_u14_u1_n144 ) , .A( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n180 ) );
  INV_X1 u1_u14_u1_U93 (.A( u1_u14_u1_n130 ) , .ZN( u1_u14_u1_n179 ) );
  NAND4_X1 u1_u14_u1_U94 (.ZN( u1_out14_28 ) , .A4( u1_u14_u1_n124 ) , .A3( u1_u14_u1_n125 ) , .A2( u1_u14_u1_n126 ) , .A1( u1_u14_u1_n127 ) );
  OAI21_X1 u1_u14_u1_U95 (.ZN( u1_u14_u1_n127 ) , .B2( u1_u14_u1_n139 ) , .B1( u1_u14_u1_n175 ) , .A( u1_u14_u1_n183 ) );
  OAI21_X1 u1_u14_u1_U96 (.ZN( u1_u14_u1_n126 ) , .B2( u1_u14_u1_n140 ) , .A( u1_u14_u1_n146 ) , .B1( u1_u14_u1_n178 ) );
  NAND3_X1 u1_u14_u1_U97 (.A3( u1_u14_u1_n149 ) , .A2( u1_u14_u1_n150 ) , .A1( u1_u14_u1_n151 ) , .ZN( u1_u14_u1_n164 ) );
  NAND3_X1 u1_u14_u1_U98 (.A3( u1_u14_u1_n134 ) , .A2( u1_u14_u1_n135 ) , .ZN( u1_u14_u1_n136 ) , .A1( u1_u14_u1_n151 ) );
  NAND3_X1 u1_u14_u1_U99 (.A1( u1_u14_u1_n133 ) , .ZN( u1_u14_u1_n137 ) , .A2( u1_u14_u1_n154 ) , .A3( u1_u14_u1_n181 ) );
  XOR2_X1 u1_u15_U10 (.A( u1_FP_62 ) , .B( u1_K16_45 ) , .Z( u1_u15_X_45 ) );
  XOR2_X1 u1_u15_U9 (.A( u1_FP_63 ) , .B( u1_K16_46 ) , .Z( u1_u15_X_46 ) );
  OAI21_X1 u1_u15_u7_U10 (.A( u1_u15_u7_n161 ) , .B1( u1_u15_u7_n168 ) , .B2( u1_u15_u7_n173 ) , .ZN( u1_u15_u7_n91 ) );
  AOI211_X1 u1_u15_u7_U11 (.A( u1_u15_u7_n117 ) , .ZN( u1_u15_u7_n118 ) , .C2( u1_u15_u7_n126 ) , .C1( u1_u15_u7_n177 ) , .B( u1_u15_u7_n180 ) );
  OAI22_X1 u1_u15_u7_U12 (.B1( u1_u15_u7_n115 ) , .ZN( u1_u15_u7_n117 ) , .A2( u1_u15_u7_n133 ) , .A1( u1_u15_u7_n137 ) , .B2( u1_u15_u7_n162 ) );
  INV_X1 u1_u15_u7_U13 (.A( u1_u15_u7_n116 ) , .ZN( u1_u15_u7_n180 ) );
  NOR3_X1 u1_u15_u7_U14 (.ZN( u1_u15_u7_n115 ) , .A3( u1_u15_u7_n145 ) , .A2( u1_u15_u7_n168 ) , .A1( u1_u15_u7_n169 ) );
  OAI211_X1 u1_u15_u7_U15 (.B( u1_u15_u7_n122 ) , .A( u1_u15_u7_n123 ) , .C2( u1_u15_u7_n124 ) , .ZN( u1_u15_u7_n154 ) , .C1( u1_u15_u7_n162 ) );
  AOI222_X1 u1_u15_u7_U16 (.ZN( u1_u15_u7_n122 ) , .C2( u1_u15_u7_n126 ) , .C1( u1_u15_u7_n145 ) , .B1( u1_u15_u7_n161 ) , .A2( u1_u15_u7_n165 ) , .B2( u1_u15_u7_n170 ) , .A1( u1_u15_u7_n176 ) );
  INV_X1 u1_u15_u7_U17 (.A( u1_u15_u7_n133 ) , .ZN( u1_u15_u7_n176 ) );
  NOR3_X1 u1_u15_u7_U18 (.A2( u1_u15_u7_n134 ) , .A1( u1_u15_u7_n135 ) , .ZN( u1_u15_u7_n136 ) , .A3( u1_u15_u7_n171 ) );
  NOR2_X1 u1_u15_u7_U19 (.A1( u1_u15_u7_n130 ) , .A2( u1_u15_u7_n134 ) , .ZN( u1_u15_u7_n153 ) );
  INV_X1 u1_u15_u7_U20 (.A( u1_u15_u7_n101 ) , .ZN( u1_u15_u7_n165 ) );
  NOR2_X1 u1_u15_u7_U21 (.ZN( u1_u15_u7_n111 ) , .A2( u1_u15_u7_n134 ) , .A1( u1_u15_u7_n169 ) );
  AOI21_X1 u1_u15_u7_U22 (.ZN( u1_u15_u7_n104 ) , .B2( u1_u15_u7_n112 ) , .B1( u1_u15_u7_n127 ) , .A( u1_u15_u7_n164 ) );
  AOI21_X1 u1_u15_u7_U23 (.ZN( u1_u15_u7_n106 ) , .B1( u1_u15_u7_n133 ) , .B2( u1_u15_u7_n146 ) , .A( u1_u15_u7_n162 ) );
  AOI21_X1 u1_u15_u7_U24 (.A( u1_u15_u7_n101 ) , .ZN( u1_u15_u7_n107 ) , .B2( u1_u15_u7_n128 ) , .B1( u1_u15_u7_n175 ) );
  INV_X1 u1_u15_u7_U25 (.A( u1_u15_u7_n138 ) , .ZN( u1_u15_u7_n171 ) );
  INV_X1 u1_u15_u7_U26 (.A( u1_u15_u7_n131 ) , .ZN( u1_u15_u7_n177 ) );
  INV_X1 u1_u15_u7_U27 (.A( u1_u15_u7_n110 ) , .ZN( u1_u15_u7_n174 ) );
  NAND2_X1 u1_u15_u7_U28 (.A1( u1_u15_u7_n129 ) , .A2( u1_u15_u7_n132 ) , .ZN( u1_u15_u7_n149 ) );
  NAND2_X1 u1_u15_u7_U29 (.A1( u1_u15_u7_n113 ) , .A2( u1_u15_u7_n124 ) , .ZN( u1_u15_u7_n130 ) );
  INV_X1 u1_u15_u7_U3 (.A( u1_u15_u7_n111 ) , .ZN( u1_u15_u7_n170 ) );
  INV_X1 u1_u15_u7_U30 (.A( u1_u15_u7_n112 ) , .ZN( u1_u15_u7_n173 ) );
  INV_X1 u1_u15_u7_U31 (.A( u1_u15_u7_n128 ) , .ZN( u1_u15_u7_n168 ) );
  INV_X1 u1_u15_u7_U32 (.A( u1_u15_u7_n148 ) , .ZN( u1_u15_u7_n169 ) );
  INV_X1 u1_u15_u7_U33 (.A( u1_u15_u7_n127 ) , .ZN( u1_u15_u7_n179 ) );
  NOR2_X1 u1_u15_u7_U34 (.ZN( u1_u15_u7_n101 ) , .A2( u1_u15_u7_n150 ) , .A1( u1_u15_u7_n156 ) );
  AOI211_X1 u1_u15_u7_U35 (.B( u1_u15_u7_n154 ) , .A( u1_u15_u7_n155 ) , .C1( u1_u15_u7_n156 ) , .ZN( u1_u15_u7_n157 ) , .C2( u1_u15_u7_n172 ) );
  INV_X1 u1_u15_u7_U36 (.A( u1_u15_u7_n153 ) , .ZN( u1_u15_u7_n172 ) );
  AOI211_X1 u1_u15_u7_U37 (.B( u1_u15_u7_n139 ) , .A( u1_u15_u7_n140 ) , .C2( u1_u15_u7_n141 ) , .ZN( u1_u15_u7_n142 ) , .C1( u1_u15_u7_n156 ) );
  NAND4_X1 u1_u15_u7_U38 (.A3( u1_u15_u7_n127 ) , .A2( u1_u15_u7_n128 ) , .A1( u1_u15_u7_n129 ) , .ZN( u1_u15_u7_n141 ) , .A4( u1_u15_u7_n147 ) );
  AOI21_X1 u1_u15_u7_U39 (.A( u1_u15_u7_n137 ) , .B1( u1_u15_u7_n138 ) , .ZN( u1_u15_u7_n139 ) , .B2( u1_u15_u7_n146 ) );
  INV_X1 u1_u15_u7_U4 (.A( u1_u15_u7_n149 ) , .ZN( u1_u15_u7_n175 ) );
  OAI22_X1 u1_u15_u7_U40 (.B1( u1_u15_u7_n136 ) , .ZN( u1_u15_u7_n140 ) , .A1( u1_u15_u7_n153 ) , .B2( u1_u15_u7_n162 ) , .A2( u1_u15_u7_n164 ) );
  AOI21_X1 u1_u15_u7_U41 (.ZN( u1_u15_u7_n123 ) , .B1( u1_u15_u7_n165 ) , .B2( u1_u15_u7_n177 ) , .A( u1_u15_u7_n97 ) );
  AOI21_X1 u1_u15_u7_U42 (.B2( u1_u15_u7_n113 ) , .B1( u1_u15_u7_n124 ) , .A( u1_u15_u7_n125 ) , .ZN( u1_u15_u7_n97 ) );
  INV_X1 u1_u15_u7_U43 (.A( u1_u15_u7_n125 ) , .ZN( u1_u15_u7_n161 ) );
  INV_X1 u1_u15_u7_U44 (.A( u1_u15_u7_n152 ) , .ZN( u1_u15_u7_n162 ) );
  AOI22_X1 u1_u15_u7_U45 (.A2( u1_u15_u7_n114 ) , .ZN( u1_u15_u7_n119 ) , .B1( u1_u15_u7_n130 ) , .A1( u1_u15_u7_n156 ) , .B2( u1_u15_u7_n165 ) );
  NAND2_X1 u1_u15_u7_U46 (.A2( u1_u15_u7_n112 ) , .ZN( u1_u15_u7_n114 ) , .A1( u1_u15_u7_n175 ) );
  AOI22_X1 u1_u15_u7_U47 (.B2( u1_u15_u7_n149 ) , .B1( u1_u15_u7_n150 ) , .A2( u1_u15_u7_n151 ) , .A1( u1_u15_u7_n152 ) , .ZN( u1_u15_u7_n158 ) );
  AND2_X1 u1_u15_u7_U48 (.ZN( u1_u15_u7_n145 ) , .A2( u1_u15_u7_n98 ) , .A1( u1_u15_u7_n99 ) );
  NOR2_X1 u1_u15_u7_U49 (.ZN( u1_u15_u7_n137 ) , .A1( u1_u15_u7_n150 ) , .A2( u1_u15_u7_n161 ) );
  INV_X1 u1_u15_u7_U5 (.A( u1_u15_u7_n154 ) , .ZN( u1_u15_u7_n178 ) );
  AOI21_X1 u1_u15_u7_U50 (.ZN( u1_u15_u7_n105 ) , .B2( u1_u15_u7_n110 ) , .A( u1_u15_u7_n125 ) , .B1( u1_u15_u7_n147 ) );
  NAND2_X1 u1_u15_u7_U51 (.ZN( u1_u15_u7_n146 ) , .A1( u1_u15_u7_n95 ) , .A2( u1_u15_u7_n98 ) );
  NAND2_X1 u1_u15_u7_U52 (.A2( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n147 ) , .A1( u1_u15_u7_n93 ) );
  NAND2_X1 u1_u15_u7_U53 (.A1( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n127 ) , .A2( u1_u15_u7_n99 ) );
  OR2_X1 u1_u15_u7_U54 (.ZN( u1_u15_u7_n126 ) , .A2( u1_u15_u7_n152 ) , .A1( u1_u15_u7_n156 ) );
  NAND2_X1 u1_u15_u7_U55 (.A2( u1_u15_u7_n102 ) , .A1( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n133 ) );
  NAND2_X1 u1_u15_u7_U56 (.ZN( u1_u15_u7_n112 ) , .A2( u1_u15_u7_n96 ) , .A1( u1_u15_u7_n99 ) );
  NAND2_X1 u1_u15_u7_U57 (.A2( u1_u15_u7_n102 ) , .ZN( u1_u15_u7_n128 ) , .A1( u1_u15_u7_n98 ) );
  NAND2_X1 u1_u15_u7_U58 (.A1( u1_u15_u7_n100 ) , .ZN( u1_u15_u7_n113 ) , .A2( u1_u15_u7_n93 ) );
  NAND2_X1 u1_u15_u7_U59 (.A2( u1_u15_u7_n102 ) , .ZN( u1_u15_u7_n124 ) , .A1( u1_u15_u7_n96 ) );
  AOI211_X1 u1_u15_u7_U6 (.ZN( u1_u15_u7_n116 ) , .A( u1_u15_u7_n155 ) , .C1( u1_u15_u7_n161 ) , .C2( u1_u15_u7_n171 ) , .B( u1_u15_u7_n94 ) );
  NAND2_X1 u1_u15_u7_U60 (.ZN( u1_u15_u7_n110 ) , .A1( u1_u15_u7_n95 ) , .A2( u1_u15_u7_n96 ) );
  INV_X1 u1_u15_u7_U61 (.A( u1_u15_u7_n150 ) , .ZN( u1_u15_u7_n164 ) );
  AND2_X1 u1_u15_u7_U62 (.ZN( u1_u15_u7_n134 ) , .A1( u1_u15_u7_n93 ) , .A2( u1_u15_u7_n98 ) );
  NAND2_X1 u1_u15_u7_U63 (.A1( u1_u15_u7_n100 ) , .A2( u1_u15_u7_n102 ) , .ZN( u1_u15_u7_n129 ) );
  NAND2_X1 u1_u15_u7_U64 (.A2( u1_u15_u7_n103 ) , .ZN( u1_u15_u7_n131 ) , .A1( u1_u15_u7_n95 ) );
  NAND2_X1 u1_u15_u7_U65 (.A1( u1_u15_u7_n100 ) , .ZN( u1_u15_u7_n138 ) , .A2( u1_u15_u7_n99 ) );
  NAND2_X1 u1_u15_u7_U66 (.ZN( u1_u15_u7_n132 ) , .A1( u1_u15_u7_n93 ) , .A2( u1_u15_u7_n96 ) );
  NAND2_X1 u1_u15_u7_U67 (.A1( u1_u15_u7_n100 ) , .ZN( u1_u15_u7_n148 ) , .A2( u1_u15_u7_n95 ) );
  NOR2_X1 u1_u15_u7_U68 (.A2( u1_u15_X_47 ) , .ZN( u1_u15_u7_n150 ) , .A1( u1_u15_u7_n163 ) );
  NOR2_X1 u1_u15_u7_U69 (.A2( u1_u15_X_43 ) , .A1( u1_u15_X_44 ) , .ZN( u1_u15_u7_n103 ) );
  OAI222_X1 u1_u15_u7_U7 (.C2( u1_u15_u7_n101 ) , .B2( u1_u15_u7_n111 ) , .A1( u1_u15_u7_n113 ) , .C1( u1_u15_u7_n146 ) , .A2( u1_u15_u7_n162 ) , .B1( u1_u15_u7_n164 ) , .ZN( u1_u15_u7_n94 ) );
  NOR2_X1 u1_u15_u7_U70 (.A2( u1_u15_X_48 ) , .A1( u1_u15_u7_n166 ) , .ZN( u1_u15_u7_n95 ) );
  NOR2_X1 u1_u15_u7_U71 (.A2( u1_u15_X_45 ) , .A1( u1_u15_X_48 ) , .ZN( u1_u15_u7_n99 ) );
  NOR2_X1 u1_u15_u7_U72 (.A2( u1_u15_X_44 ) , .A1( u1_u15_u7_n167 ) , .ZN( u1_u15_u7_n98 ) );
  NOR2_X1 u1_u15_u7_U73 (.A2( u1_u15_X_46 ) , .A1( u1_u15_X_47 ) , .ZN( u1_u15_u7_n152 ) );
  AND2_X1 u1_u15_u7_U74 (.A1( u1_u15_X_47 ) , .ZN( u1_u15_u7_n156 ) , .A2( u1_u15_u7_n163 ) );
  NAND2_X1 u1_u15_u7_U75 (.A2( u1_u15_X_46 ) , .A1( u1_u15_X_47 ) , .ZN( u1_u15_u7_n125 ) );
  AND2_X1 u1_u15_u7_U76 (.A2( u1_u15_X_45 ) , .A1( u1_u15_X_48 ) , .ZN( u1_u15_u7_n102 ) );
  AND2_X1 u1_u15_u7_U77 (.A2( u1_u15_X_43 ) , .A1( u1_u15_X_44 ) , .ZN( u1_u15_u7_n96 ) );
  AND2_X1 u1_u15_u7_U78 (.A1( u1_u15_X_44 ) , .ZN( u1_u15_u7_n100 ) , .A2( u1_u15_u7_n167 ) );
  AND2_X1 u1_u15_u7_U79 (.A1( u1_u15_X_48 ) , .A2( u1_u15_u7_n166 ) , .ZN( u1_u15_u7_n93 ) );
  OAI221_X1 u1_u15_u7_U8 (.C1( u1_u15_u7_n101 ) , .C2( u1_u15_u7_n147 ) , .ZN( u1_u15_u7_n155 ) , .B2( u1_u15_u7_n162 ) , .A( u1_u15_u7_n91 ) , .B1( u1_u15_u7_n92 ) );
  INV_X1 u1_u15_u7_U80 (.A( u1_u15_X_46 ) , .ZN( u1_u15_u7_n163 ) );
  INV_X1 u1_u15_u7_U81 (.A( u1_u15_X_45 ) , .ZN( u1_u15_u7_n166 ) );
  INV_X1 u1_u15_u7_U82 (.A( u1_u15_X_43 ) , .ZN( u1_u15_u7_n167 ) );
  NAND4_X1 u1_u15_u7_U83 (.ZN( u1_out15_5 ) , .A4( u1_u15_u7_n108 ) , .A3( u1_u15_u7_n109 ) , .A1( u1_u15_u7_n116 ) , .A2( u1_u15_u7_n123 ) );
  AOI22_X1 u1_u15_u7_U84 (.ZN( u1_u15_u7_n109 ) , .A2( u1_u15_u7_n126 ) , .B2( u1_u15_u7_n145 ) , .B1( u1_u15_u7_n156 ) , .A1( u1_u15_u7_n171 ) );
  NOR4_X1 u1_u15_u7_U85 (.A4( u1_u15_u7_n104 ) , .A3( u1_u15_u7_n105 ) , .A2( u1_u15_u7_n106 ) , .A1( u1_u15_u7_n107 ) , .ZN( u1_u15_u7_n108 ) );
  NAND4_X1 u1_u15_u7_U86 (.ZN( u1_out15_27 ) , .A4( u1_u15_u7_n118 ) , .A3( u1_u15_u7_n119 ) , .A2( u1_u15_u7_n120 ) , .A1( u1_u15_u7_n121 ) );
  OAI21_X1 u1_u15_u7_U87 (.ZN( u1_u15_u7_n121 ) , .B2( u1_u15_u7_n145 ) , .A( u1_u15_u7_n150 ) , .B1( u1_u15_u7_n174 ) );
  OAI21_X1 u1_u15_u7_U88 (.ZN( u1_u15_u7_n120 ) , .A( u1_u15_u7_n161 ) , .B2( u1_u15_u7_n170 ) , .B1( u1_u15_u7_n179 ) );
  NAND4_X1 u1_u15_u7_U89 (.ZN( u1_out15_21 ) , .A4( u1_u15_u7_n157 ) , .A3( u1_u15_u7_n158 ) , .A2( u1_u15_u7_n159 ) , .A1( u1_u15_u7_n160 ) );
  AND3_X1 u1_u15_u7_U9 (.A3( u1_u15_u7_n110 ) , .A2( u1_u15_u7_n127 ) , .A1( u1_u15_u7_n132 ) , .ZN( u1_u15_u7_n92 ) );
  OAI21_X1 u1_u15_u7_U90 (.B1( u1_u15_u7_n145 ) , .ZN( u1_u15_u7_n160 ) , .A( u1_u15_u7_n161 ) , .B2( u1_u15_u7_n177 ) );
  OAI21_X1 u1_u15_u7_U91 (.ZN( u1_u15_u7_n159 ) , .A( u1_u15_u7_n165 ) , .B2( u1_u15_u7_n171 ) , .B1( u1_u15_u7_n174 ) );
  NAND4_X1 u1_u15_u7_U92 (.ZN( u1_out15_15 ) , .A4( u1_u15_u7_n142 ) , .A3( u1_u15_u7_n143 ) , .A2( u1_u15_u7_n144 ) , .A1( u1_u15_u7_n178 ) );
  OR2_X1 u1_u15_u7_U93 (.A2( u1_u15_u7_n125 ) , .A1( u1_u15_u7_n129 ) , .ZN( u1_u15_u7_n144 ) );
  AOI22_X1 u1_u15_u7_U94 (.A2( u1_u15_u7_n126 ) , .ZN( u1_u15_u7_n143 ) , .B2( u1_u15_u7_n165 ) , .B1( u1_u15_u7_n173 ) , .A1( u1_u15_u7_n174 ) );
  NAND3_X1 u1_u15_u7_U95 (.A3( u1_u15_u7_n146 ) , .A2( u1_u15_u7_n147 ) , .A1( u1_u15_u7_n148 ) , .ZN( u1_u15_u7_n151 ) );
  NAND3_X1 u1_u15_u7_U96 (.A3( u1_u15_u7_n131 ) , .A2( u1_u15_u7_n132 ) , .A1( u1_u15_u7_n133 ) , .ZN( u1_u15_u7_n135 ) );
  XOR2_X1 u1_u1_U22 (.B( u1_K2_34 ) , .A( u1_R0_23 ) , .Z( u1_u1_X_34 ) );
  XOR2_X1 u1_u1_U23 (.B( u1_K2_33 ) , .A( u1_R0_22 ) , .Z( u1_u1_X_33 ) );
  INV_X1 u1_u1_u5_U10 (.A( u1_u1_u5_n121 ) , .ZN( u1_u1_u5_n177 ) );
  NOR3_X1 u1_u1_u5_U100 (.A3( u1_u1_u5_n141 ) , .A1( u1_u1_u5_n142 ) , .ZN( u1_u1_u5_n143 ) , .A2( u1_u1_u5_n191 ) );
  NAND4_X1 u1_u1_u5_U101 (.ZN( u1_out1_4 ) , .A4( u1_u1_u5_n112 ) , .A2( u1_u1_u5_n113 ) , .A1( u1_u1_u5_n114 ) , .A3( u1_u1_u5_n195 ) );
  AOI211_X1 u1_u1_u5_U102 (.A( u1_u1_u5_n110 ) , .C1( u1_u1_u5_n111 ) , .ZN( u1_u1_u5_n112 ) , .B( u1_u1_u5_n118 ) , .C2( u1_u1_u5_n177 ) );
  AOI222_X1 u1_u1_u5_U103 (.ZN( u1_u1_u5_n113 ) , .A1( u1_u1_u5_n131 ) , .C1( u1_u1_u5_n148 ) , .B2( u1_u1_u5_n174 ) , .C2( u1_u1_u5_n178 ) , .A2( u1_u1_u5_n179 ) , .B1( u1_u1_u5_n99 ) );
  NAND3_X1 u1_u1_u5_U104 (.A2( u1_u1_u5_n154 ) , .A3( u1_u1_u5_n158 ) , .A1( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n99 ) );
  NOR2_X1 u1_u1_u5_U11 (.ZN( u1_u1_u5_n160 ) , .A2( u1_u1_u5_n173 ) , .A1( u1_u1_u5_n177 ) );
  INV_X1 u1_u1_u5_U12 (.A( u1_u1_u5_n150 ) , .ZN( u1_u1_u5_n174 ) );
  AOI21_X1 u1_u1_u5_U13 (.A( u1_u1_u5_n160 ) , .B2( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n162 ) , .B1( u1_u1_u5_n192 ) );
  INV_X1 u1_u1_u5_U14 (.A( u1_u1_u5_n159 ) , .ZN( u1_u1_u5_n192 ) );
  AOI21_X1 u1_u1_u5_U15 (.A( u1_u1_u5_n156 ) , .B2( u1_u1_u5_n157 ) , .B1( u1_u1_u5_n158 ) , .ZN( u1_u1_u5_n163 ) );
  AOI21_X1 u1_u1_u5_U16 (.B2( u1_u1_u5_n139 ) , .B1( u1_u1_u5_n140 ) , .ZN( u1_u1_u5_n141 ) , .A( u1_u1_u5_n150 ) );
  OAI21_X1 u1_u1_u5_U17 (.A( u1_u1_u5_n133 ) , .B2( u1_u1_u5_n134 ) , .B1( u1_u1_u5_n135 ) , .ZN( u1_u1_u5_n142 ) );
  OAI21_X1 u1_u1_u5_U18 (.ZN( u1_u1_u5_n133 ) , .B2( u1_u1_u5_n147 ) , .A( u1_u1_u5_n173 ) , .B1( u1_u1_u5_n188 ) );
  NAND2_X1 u1_u1_u5_U19 (.A2( u1_u1_u5_n119 ) , .A1( u1_u1_u5_n123 ) , .ZN( u1_u1_u5_n137 ) );
  INV_X1 u1_u1_u5_U20 (.A( u1_u1_u5_n155 ) , .ZN( u1_u1_u5_n194 ) );
  NAND2_X1 u1_u1_u5_U21 (.A1( u1_u1_u5_n121 ) , .ZN( u1_u1_u5_n132 ) , .A2( u1_u1_u5_n172 ) );
  NAND2_X1 u1_u1_u5_U22 (.A2( u1_u1_u5_n122 ) , .ZN( u1_u1_u5_n136 ) , .A1( u1_u1_u5_n154 ) );
  NAND2_X1 u1_u1_u5_U23 (.A2( u1_u1_u5_n119 ) , .A1( u1_u1_u5_n120 ) , .ZN( u1_u1_u5_n159 ) );
  INV_X1 u1_u1_u5_U24 (.A( u1_u1_u5_n156 ) , .ZN( u1_u1_u5_n175 ) );
  INV_X1 u1_u1_u5_U25 (.A( u1_u1_u5_n158 ) , .ZN( u1_u1_u5_n188 ) );
  INV_X1 u1_u1_u5_U26 (.A( u1_u1_u5_n152 ) , .ZN( u1_u1_u5_n179 ) );
  INV_X1 u1_u1_u5_U27 (.A( u1_u1_u5_n140 ) , .ZN( u1_u1_u5_n182 ) );
  INV_X1 u1_u1_u5_U28 (.A( u1_u1_u5_n151 ) , .ZN( u1_u1_u5_n183 ) );
  INV_X1 u1_u1_u5_U29 (.A( u1_u1_u5_n123 ) , .ZN( u1_u1_u5_n185 ) );
  NOR2_X1 u1_u1_u5_U3 (.ZN( u1_u1_u5_n134 ) , .A1( u1_u1_u5_n183 ) , .A2( u1_u1_u5_n190 ) );
  INV_X1 u1_u1_u5_U30 (.A( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n184 ) );
  INV_X1 u1_u1_u5_U31 (.A( u1_u1_u5_n139 ) , .ZN( u1_u1_u5_n189 ) );
  INV_X1 u1_u1_u5_U32 (.A( u1_u1_u5_n157 ) , .ZN( u1_u1_u5_n190 ) );
  INV_X1 u1_u1_u5_U33 (.A( u1_u1_u5_n120 ) , .ZN( u1_u1_u5_n193 ) );
  NAND2_X1 u1_u1_u5_U34 (.ZN( u1_u1_u5_n111 ) , .A1( u1_u1_u5_n140 ) , .A2( u1_u1_u5_n155 ) );
  INV_X1 u1_u1_u5_U35 (.A( u1_u1_u5_n117 ) , .ZN( u1_u1_u5_n196 ) );
  OAI221_X1 u1_u1_u5_U36 (.A( u1_u1_u5_n116 ) , .ZN( u1_u1_u5_n117 ) , .B2( u1_u1_u5_n119 ) , .C1( u1_u1_u5_n153 ) , .C2( u1_u1_u5_n158 ) , .B1( u1_u1_u5_n172 ) );
  AOI222_X1 u1_u1_u5_U37 (.ZN( u1_u1_u5_n116 ) , .B2( u1_u1_u5_n145 ) , .C1( u1_u1_u5_n148 ) , .A2( u1_u1_u5_n174 ) , .C2( u1_u1_u5_n177 ) , .B1( u1_u1_u5_n187 ) , .A1( u1_u1_u5_n193 ) );
  INV_X1 u1_u1_u5_U38 (.A( u1_u1_u5_n115 ) , .ZN( u1_u1_u5_n187 ) );
  NOR2_X1 u1_u1_u5_U39 (.ZN( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n170 ) , .A2( u1_u1_u5_n180 ) );
  INV_X1 u1_u1_u5_U4 (.A( u1_u1_u5_n138 ) , .ZN( u1_u1_u5_n191 ) );
  AOI22_X1 u1_u1_u5_U40 (.B2( u1_u1_u5_n131 ) , .A2( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n169 ) , .B1( u1_u1_u5_n174 ) , .A1( u1_u1_u5_n185 ) );
  NOR2_X1 u1_u1_u5_U41 (.A1( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n150 ) , .A2( u1_u1_u5_n173 ) );
  AOI21_X1 u1_u1_u5_U42 (.A( u1_u1_u5_n118 ) , .B2( u1_u1_u5_n145 ) , .ZN( u1_u1_u5_n168 ) , .B1( u1_u1_u5_n186 ) );
  INV_X1 u1_u1_u5_U43 (.A( u1_u1_u5_n122 ) , .ZN( u1_u1_u5_n186 ) );
  NOR2_X1 u1_u1_u5_U44 (.A1( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n152 ) , .A2( u1_u1_u5_n176 ) );
  NOR2_X1 u1_u1_u5_U45 (.A1( u1_u1_u5_n115 ) , .ZN( u1_u1_u5_n118 ) , .A2( u1_u1_u5_n153 ) );
  NOR2_X1 u1_u1_u5_U46 (.A2( u1_u1_u5_n145 ) , .ZN( u1_u1_u5_n156 ) , .A1( u1_u1_u5_n174 ) );
  NOR2_X1 u1_u1_u5_U47 (.ZN( u1_u1_u5_n121 ) , .A2( u1_u1_u5_n145 ) , .A1( u1_u1_u5_n176 ) );
  AOI22_X1 u1_u1_u5_U48 (.ZN( u1_u1_u5_n114 ) , .A2( u1_u1_u5_n137 ) , .A1( u1_u1_u5_n145 ) , .B2( u1_u1_u5_n175 ) , .B1( u1_u1_u5_n193 ) );
  OAI211_X1 u1_u1_u5_U49 (.B( u1_u1_u5_n124 ) , .A( u1_u1_u5_n125 ) , .C2( u1_u1_u5_n126 ) , .C1( u1_u1_u5_n127 ) , .ZN( u1_u1_u5_n128 ) );
  OAI21_X1 u1_u1_u5_U5 (.B2( u1_u1_u5_n136 ) , .B1( u1_u1_u5_n137 ) , .ZN( u1_u1_u5_n138 ) , .A( u1_u1_u5_n177 ) );
  OAI21_X1 u1_u1_u5_U50 (.ZN( u1_u1_u5_n124 ) , .A( u1_u1_u5_n177 ) , .B2( u1_u1_u5_n183 ) , .B1( u1_u1_u5_n189 ) );
  NOR3_X1 u1_u1_u5_U51 (.ZN( u1_u1_u5_n127 ) , .A1( u1_u1_u5_n136 ) , .A3( u1_u1_u5_n148 ) , .A2( u1_u1_u5_n182 ) );
  OAI21_X1 u1_u1_u5_U52 (.ZN( u1_u1_u5_n125 ) , .A( u1_u1_u5_n174 ) , .B2( u1_u1_u5_n185 ) , .B1( u1_u1_u5_n190 ) );
  AOI21_X1 u1_u1_u5_U53 (.A( u1_u1_u5_n153 ) , .B2( u1_u1_u5_n154 ) , .B1( u1_u1_u5_n155 ) , .ZN( u1_u1_u5_n164 ) );
  AOI21_X1 u1_u1_u5_U54 (.ZN( u1_u1_u5_n110 ) , .B1( u1_u1_u5_n122 ) , .B2( u1_u1_u5_n139 ) , .A( u1_u1_u5_n153 ) );
  INV_X1 u1_u1_u5_U55 (.A( u1_u1_u5_n153 ) , .ZN( u1_u1_u5_n176 ) );
  INV_X1 u1_u1_u5_U56 (.A( u1_u1_u5_n126 ) , .ZN( u1_u1_u5_n173 ) );
  AND2_X1 u1_u1_u5_U57 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n147 ) );
  AND2_X1 u1_u1_u5_U58 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n148 ) );
  NAND2_X1 u1_u1_u5_U59 (.A1( u1_u1_u5_n105 ) , .A2( u1_u1_u5_n106 ) , .ZN( u1_u1_u5_n158 ) );
  INV_X1 u1_u1_u5_U6 (.A( u1_u1_u5_n135 ) , .ZN( u1_u1_u5_n178 ) );
  NAND2_X1 u1_u1_u5_U60 (.A2( u1_u1_u5_n108 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n139 ) );
  NAND2_X1 u1_u1_u5_U61 (.A1( u1_u1_u5_n106 ) , .A2( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n119 ) );
  NAND2_X1 u1_u1_u5_U62 (.A2( u1_u1_u5_n103 ) , .A1( u1_u1_u5_n105 ) , .ZN( u1_u1_u5_n140 ) );
  NAND2_X1 u1_u1_u5_U63 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n105 ) , .ZN( u1_u1_u5_n155 ) );
  NAND2_X1 u1_u1_u5_U64 (.A2( u1_u1_u5_n106 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n122 ) );
  NAND2_X1 u1_u1_u5_U65 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n106 ) , .ZN( u1_u1_u5_n115 ) );
  NAND2_X1 u1_u1_u5_U66 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n103 ) , .ZN( u1_u1_u5_n161 ) );
  NAND2_X1 u1_u1_u5_U67 (.A1( u1_u1_u5_n105 ) , .A2( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n154 ) );
  INV_X1 u1_u1_u5_U68 (.A( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n172 ) );
  NAND2_X1 u1_u1_u5_U69 (.A1( u1_u1_u5_n103 ) , .A2( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n123 ) );
  OAI22_X1 u1_u1_u5_U7 (.B2( u1_u1_u5_n149 ) , .B1( u1_u1_u5_n150 ) , .A2( u1_u1_u5_n151 ) , .A1( u1_u1_u5_n152 ) , .ZN( u1_u1_u5_n165 ) );
  NAND2_X1 u1_u1_u5_U70 (.A2( u1_u1_u5_n103 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n151 ) );
  NAND2_X1 u1_u1_u5_U71 (.A2( u1_u1_u5_n107 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n120 ) );
  NAND2_X1 u1_u1_u5_U72 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n157 ) );
  AND2_X1 u1_u1_u5_U73 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n104 ) , .ZN( u1_u1_u5_n131 ) );
  INV_X1 u1_u1_u5_U74 (.A( u1_u1_u5_n102 ) , .ZN( u1_u1_u5_n195 ) );
  OAI221_X1 u1_u1_u5_U75 (.A( u1_u1_u5_n101 ) , .ZN( u1_u1_u5_n102 ) , .C2( u1_u1_u5_n115 ) , .C1( u1_u1_u5_n126 ) , .B1( u1_u1_u5_n134 ) , .B2( u1_u1_u5_n160 ) );
  OAI21_X1 u1_u1_u5_U76 (.ZN( u1_u1_u5_n101 ) , .B1( u1_u1_u5_n137 ) , .A( u1_u1_u5_n146 ) , .B2( u1_u1_u5_n147 ) );
  NOR2_X1 u1_u1_u5_U77 (.A2( u1_u1_X_34 ) , .A1( u1_u1_X_35 ) , .ZN( u1_u1_u5_n145 ) );
  NOR2_X1 u1_u1_u5_U78 (.A2( u1_u1_X_34 ) , .ZN( u1_u1_u5_n146 ) , .A1( u1_u1_u5_n171 ) );
  NOR2_X1 u1_u1_u5_U79 (.A2( u1_u1_X_31 ) , .A1( u1_u1_X_32 ) , .ZN( u1_u1_u5_n103 ) );
  NOR3_X1 u1_u1_u5_U8 (.A2( u1_u1_u5_n147 ) , .A1( u1_u1_u5_n148 ) , .ZN( u1_u1_u5_n149 ) , .A3( u1_u1_u5_n194 ) );
  NOR2_X1 u1_u1_u5_U80 (.A2( u1_u1_X_36 ) , .ZN( u1_u1_u5_n105 ) , .A1( u1_u1_u5_n180 ) );
  NOR2_X1 u1_u1_u5_U81 (.A2( u1_u1_X_33 ) , .ZN( u1_u1_u5_n108 ) , .A1( u1_u1_u5_n170 ) );
  NOR2_X1 u1_u1_u5_U82 (.A2( u1_u1_X_33 ) , .A1( u1_u1_X_36 ) , .ZN( u1_u1_u5_n107 ) );
  NOR2_X1 u1_u1_u5_U83 (.A2( u1_u1_X_31 ) , .ZN( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n181 ) );
  NAND2_X1 u1_u1_u5_U84 (.A2( u1_u1_X_34 ) , .A1( u1_u1_X_35 ) , .ZN( u1_u1_u5_n153 ) );
  NAND2_X1 u1_u1_u5_U85 (.A1( u1_u1_X_34 ) , .ZN( u1_u1_u5_n126 ) , .A2( u1_u1_u5_n171 ) );
  AND2_X1 u1_u1_u5_U86 (.A1( u1_u1_X_31 ) , .A2( u1_u1_X_32 ) , .ZN( u1_u1_u5_n106 ) );
  AND2_X1 u1_u1_u5_U87 (.A1( u1_u1_X_31 ) , .ZN( u1_u1_u5_n109 ) , .A2( u1_u1_u5_n181 ) );
  INV_X1 u1_u1_u5_U88 (.A( u1_u1_X_33 ) , .ZN( u1_u1_u5_n180 ) );
  INV_X1 u1_u1_u5_U89 (.A( u1_u1_X_35 ) , .ZN( u1_u1_u5_n171 ) );
  NOR2_X1 u1_u1_u5_U9 (.ZN( u1_u1_u5_n135 ) , .A1( u1_u1_u5_n173 ) , .A2( u1_u1_u5_n176 ) );
  INV_X1 u1_u1_u5_U90 (.A( u1_u1_X_36 ) , .ZN( u1_u1_u5_n170 ) );
  INV_X1 u1_u1_u5_U91 (.A( u1_u1_X_32 ) , .ZN( u1_u1_u5_n181 ) );
  NAND4_X1 u1_u1_u5_U92 (.ZN( u1_out1_29 ) , .A4( u1_u1_u5_n129 ) , .A3( u1_u1_u5_n130 ) , .A2( u1_u1_u5_n168 ) , .A1( u1_u1_u5_n196 ) );
  AOI221_X1 u1_u1_u5_U93 (.A( u1_u1_u5_n128 ) , .ZN( u1_u1_u5_n129 ) , .C2( u1_u1_u5_n132 ) , .B2( u1_u1_u5_n159 ) , .B1( u1_u1_u5_n176 ) , .C1( u1_u1_u5_n184 ) );
  AOI222_X1 u1_u1_u5_U94 (.ZN( u1_u1_u5_n130 ) , .A2( u1_u1_u5_n146 ) , .B1( u1_u1_u5_n147 ) , .C2( u1_u1_u5_n175 ) , .B2( u1_u1_u5_n179 ) , .A1( u1_u1_u5_n188 ) , .C1( u1_u1_u5_n194 ) );
  NAND4_X1 u1_u1_u5_U95 (.ZN( u1_out1_19 ) , .A4( u1_u1_u5_n166 ) , .A3( u1_u1_u5_n167 ) , .A2( u1_u1_u5_n168 ) , .A1( u1_u1_u5_n169 ) );
  AOI22_X1 u1_u1_u5_U96 (.B2( u1_u1_u5_n145 ) , .A2( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n167 ) , .B1( u1_u1_u5_n182 ) , .A1( u1_u1_u5_n189 ) );
  NOR4_X1 u1_u1_u5_U97 (.A4( u1_u1_u5_n162 ) , .A3( u1_u1_u5_n163 ) , .A2( u1_u1_u5_n164 ) , .A1( u1_u1_u5_n165 ) , .ZN( u1_u1_u5_n166 ) );
  NAND4_X1 u1_u1_u5_U98 (.ZN( u1_out1_11 ) , .A4( u1_u1_u5_n143 ) , .A3( u1_u1_u5_n144 ) , .A2( u1_u1_u5_n169 ) , .A1( u1_u1_u5_n196 ) );
  AOI22_X1 u1_u1_u5_U99 (.A2( u1_u1_u5_n132 ) , .ZN( u1_u1_u5_n144 ) , .B2( u1_u1_u5_n145 ) , .B1( u1_u1_u5_n184 ) , .A1( u1_u1_u5_n194 ) );
  XOR2_X1 u1_u2_U16 (.B( u1_K3_3 ) , .A( u1_R1_2 ) , .Z( u1_u2_X_3 ) );
  XOR2_X1 u1_u2_U29 (.B( u1_K3_28 ) , .A( u1_R1_19 ) , .Z( u1_u2_X_28 ) );
  XOR2_X1 u1_u2_U30 (.B( u1_K3_27 ) , .A( u1_R1_18 ) , .Z( u1_u2_X_27 ) );
  XOR2_X1 u1_u2_U6 (.B( u1_K3_4 ) , .A( u1_R1_3 ) , .Z( u1_u2_X_4 ) );
  AND3_X1 u1_u2_u0_U10 (.A2( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n127 ) , .A3( u1_u2_u0_n130 ) , .A1( u1_u2_u0_n148 ) );
  NAND2_X1 u1_u2_u0_U11 (.ZN( u1_u2_u0_n113 ) , .A1( u1_u2_u0_n139 ) , .A2( u1_u2_u0_n149 ) );
  AND2_X1 u1_u2_u0_U12 (.ZN( u1_u2_u0_n107 ) , .A1( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n140 ) );
  AND2_X1 u1_u2_u0_U13 (.A2( u1_u2_u0_n129 ) , .A1( u1_u2_u0_n130 ) , .ZN( u1_u2_u0_n151 ) );
  AND2_X1 u1_u2_u0_U14 (.A1( u1_u2_u0_n108 ) , .A2( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U15 (.A( u1_u2_u0_n143 ) , .ZN( u1_u2_u0_n173 ) );
  NOR2_X1 u1_u2_u0_U16 (.A2( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n147 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U17 (.ZN( u1_u2_u0_n172 ) , .A( u1_u2_u0_n88 ) );
  OAI222_X1 u1_u2_u0_U18 (.C1( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n125 ) , .B2( u1_u2_u0_n128 ) , .B1( u1_u2_u0_n144 ) , .A2( u1_u2_u0_n158 ) , .C2( u1_u2_u0_n161 ) , .ZN( u1_u2_u0_n88 ) );
  NOR2_X1 u1_u2_u0_U19 (.A1( u1_u2_u0_n163 ) , .A2( u1_u2_u0_n164 ) , .ZN( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U20 (.B1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n132 ) , .A( u1_u2_u0_n165 ) , .B2( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U21 (.A( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n165 ) );
  OAI221_X1 u1_u2_u0_U22 (.C1( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n122 ) , .B2( u1_u2_u0_n127 ) , .A( u1_u2_u0_n143 ) , .B1( u1_u2_u0_n144 ) , .C2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U23 (.B1( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n126 ) , .A1( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n146 ) , .B2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U24 (.B1( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n147 ) , .A2( u1_u2_u0_n90 ) , .ZN( u1_u2_u0_n91 ) );
  AND3_X1 u1_u2_u0_U25 (.A3( u1_u2_u0_n121 ) , .A2( u1_u2_u0_n125 ) , .A1( u1_u2_u0_n148 ) , .ZN( u1_u2_u0_n90 ) );
  INV_X1 u1_u2_u0_U26 (.A( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n161 ) );
  NOR2_X1 u1_u2_u0_U27 (.A1( u1_u2_u0_n120 ) , .ZN( u1_u2_u0_n143 ) , .A2( u1_u2_u0_n167 ) );
  OAI221_X1 u1_u2_u0_U28 (.C1( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n120 ) , .B1( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n141 ) , .C2( u1_u2_u0_n147 ) , .A( u1_u2_u0_n172 ) );
  AOI211_X1 u1_u2_u0_U29 (.B( u1_u2_u0_n115 ) , .A( u1_u2_u0_n116 ) , .C2( u1_u2_u0_n117 ) , .C1( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n119 ) );
  INV_X1 u1_u2_u0_U3 (.A( u1_u2_u0_n113 ) , .ZN( u1_u2_u0_n166 ) );
  AOI22_X1 u1_u2_u0_U30 (.B2( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n110 ) , .ZN( u1_u2_u0_n111 ) , .B1( u1_u2_u0_n118 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U31 (.A( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U32 (.ZN( u1_u2_u0_n104 ) , .B1( u1_u2_u0_n107 ) , .B2( u1_u2_u0_n141 ) , .A( u1_u2_u0_n144 ) );
  AOI21_X1 u1_u2_u0_U33 (.B1( u1_u2_u0_n127 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n96 ) );
  AOI21_X1 u1_u2_u0_U34 (.ZN( u1_u2_u0_n116 ) , .B2( u1_u2_u0_n142 ) , .A( u1_u2_u0_n144 ) , .B1( u1_u2_u0_n166 ) );
  NAND2_X1 u1_u2_u0_U35 (.A1( u1_u2_u0_n100 ) , .A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n125 ) );
  NAND2_X1 u1_u2_u0_U36 (.A1( u1_u2_u0_n101 ) , .A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n150 ) );
  INV_X1 u1_u2_u0_U37 (.A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n160 ) );
  NAND2_X1 u1_u2_u0_U38 (.A1( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n128 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U39 (.A1( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n129 ) , .A2( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U4 (.B1( u1_u2_u0_n114 ) , .ZN( u1_u2_u0_n115 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n161 ) );
  NAND2_X1 u1_u2_u0_U40 (.A2( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U41 (.A2( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n139 ) );
  NAND2_X1 u1_u2_u0_U42 (.ZN( u1_u2_u0_n148 ) , .A1( u1_u2_u0_n93 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U43 (.A2( u1_u2_u0_n102 ) , .A1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n149 ) );
  NAND2_X1 u1_u2_u0_U44 (.A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n114 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U45 (.A2( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n121 ) , .A1( u1_u2_u0_n93 ) );
  NAND2_X1 u1_u2_u0_U46 (.ZN( u1_u2_u0_n112 ) , .A2( u1_u2_u0_n92 ) , .A1( u1_u2_u0_n93 ) );
  OR3_X1 u1_u2_u0_U47 (.A3( u1_u2_u0_n152 ) , .A2( u1_u2_u0_n153 ) , .A1( u1_u2_u0_n154 ) , .ZN( u1_u2_u0_n155 ) );
  AOI21_X1 u1_u2_u0_U48 (.B2( u1_u2_u0_n150 ) , .B1( u1_u2_u0_n151 ) , .ZN( u1_u2_u0_n152 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U49 (.A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n145 ) , .B1( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n154 ) );
  AOI21_X1 u1_u2_u0_U5 (.B2( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n134 ) , .B1( u1_u2_u0_n151 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U50 (.A( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n148 ) , .B1( u1_u2_u0_n149 ) , .ZN( u1_u2_u0_n153 ) );
  INV_X1 u1_u2_u0_U51 (.ZN( u1_u2_u0_n171 ) , .A( u1_u2_u0_n99 ) );
  OAI211_X1 u1_u2_u0_U52 (.C2( u1_u2_u0_n140 ) , .C1( u1_u2_u0_n161 ) , .A( u1_u2_u0_n169 ) , .B( u1_u2_u0_n98 ) , .ZN( u1_u2_u0_n99 ) );
  AOI211_X1 u1_u2_u0_U53 (.C1( u1_u2_u0_n118 ) , .A( u1_u2_u0_n123 ) , .B( u1_u2_u0_n96 ) , .C2( u1_u2_u0_n97 ) , .ZN( u1_u2_u0_n98 ) );
  INV_X1 u1_u2_u0_U54 (.ZN( u1_u2_u0_n169 ) , .A( u1_u2_u0_n91 ) );
  NOR2_X1 u1_u2_u0_U55 (.A2( u1_u2_X_6 ) , .ZN( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U56 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n118 ) );
  NOR2_X1 u1_u2_u0_U57 (.A2( u1_u2_X_2 ) , .ZN( u1_u2_u0_n103 ) , .A1( u1_u2_u0_n164 ) );
  NOR2_X1 u1_u2_u0_U58 (.A2( u1_u2_X_1 ) , .A1( u1_u2_X_2 ) , .ZN( u1_u2_u0_n92 ) );
  NOR2_X1 u1_u2_u0_U59 (.A2( u1_u2_X_1 ) , .ZN( u1_u2_u0_n101 ) , .A1( u1_u2_u0_n163 ) );
  NOR2_X1 u1_u2_u0_U6 (.A1( u1_u2_u0_n108 ) , .ZN( u1_u2_u0_n123 ) , .A2( u1_u2_u0_n158 ) );
  NAND2_X1 u1_u2_u0_U60 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n144 ) );
  NOR2_X1 u1_u2_u0_U61 (.A2( u1_u2_X_5 ) , .ZN( u1_u2_u0_n136 ) , .A1( u1_u2_u0_n159 ) );
  NAND2_X1 u1_u2_u0_U62 (.A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n159 ) );
  AND2_X1 u1_u2_u0_U63 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n102 ) );
  AND2_X1 u1_u2_u0_U64 (.A1( u1_u2_X_6 ) , .A2( u1_u2_u0_n162 ) , .ZN( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U65 (.A( u1_u2_X_4 ) , .ZN( u1_u2_u0_n159 ) );
  INV_X1 u1_u2_u0_U66 (.A( u1_u2_X_1 ) , .ZN( u1_u2_u0_n164 ) );
  INV_X1 u1_u2_u0_U67 (.A( u1_u2_X_2 ) , .ZN( u1_u2_u0_n163 ) );
  INV_X1 u1_u2_u0_U68 (.ZN( u1_u2_u0_n174 ) , .A( u1_u2_u0_n89 ) );
  AOI211_X1 u1_u2_u0_U69 (.B( u1_u2_u0_n104 ) , .A( u1_u2_u0_n105 ) , .ZN( u1_u2_u0_n106 ) , .C2( u1_u2_u0_n113 ) , .C1( u1_u2_u0_n160 ) );
  OAI21_X1 u1_u2_u0_U7 (.B1( u1_u2_u0_n150 ) , .B2( u1_u2_u0_n158 ) , .A( u1_u2_u0_n172 ) , .ZN( u1_u2_u0_n89 ) );
  OR4_X1 u1_u2_u0_U70 (.ZN( u1_out2_17 ) , .A4( u1_u2_u0_n122 ) , .A2( u1_u2_u0_n123 ) , .A1( u1_u2_u0_n124 ) , .A3( u1_u2_u0_n170 ) );
  AOI21_X1 u1_u2_u0_U71 (.B2( u1_u2_u0_n107 ) , .ZN( u1_u2_u0_n124 ) , .B1( u1_u2_u0_n128 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U72 (.A( u1_u2_u0_n111 ) , .ZN( u1_u2_u0_n170 ) );
  OR4_X1 u1_u2_u0_U73 (.ZN( u1_out2_31 ) , .A4( u1_u2_u0_n155 ) , .A2( u1_u2_u0_n156 ) , .A1( u1_u2_u0_n157 ) , .A3( u1_u2_u0_n173 ) );
  AOI21_X1 u1_u2_u0_U74 (.A( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n139 ) , .B1( u1_u2_u0_n140 ) , .ZN( u1_u2_u0_n157 ) );
  AOI21_X1 u1_u2_u0_U75 (.B2( u1_u2_u0_n141 ) , .B1( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n156 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U76 (.A( u1_u2_u0_n126 ) , .ZN( u1_u2_u0_n168 ) );
  AOI211_X1 u1_u2_u0_U77 (.B( u1_u2_u0_n133 ) , .A( u1_u2_u0_n134 ) , .C2( u1_u2_u0_n135 ) , .C1( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n137 ) );
  AOI21_X1 u1_u2_u0_U78 (.B1( u1_u2_u0_n132 ) , .ZN( u1_u2_u0_n133 ) , .A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n166 ) );
  OAI22_X1 u1_u2_u0_U79 (.ZN( u1_u2_u0_n105 ) , .A2( u1_u2_u0_n132 ) , .B1( u1_u2_u0_n146 ) , .A1( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n161 ) );
  AND2_X1 u1_u2_u0_U8 (.A1( u1_u2_u0_n114 ) , .A2( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n146 ) );
  NAND2_X1 u1_u2_u0_U80 (.ZN( u1_u2_u0_n110 ) , .A2( u1_u2_u0_n132 ) , .A1( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U81 (.A( u1_u2_u0_n119 ) , .ZN( u1_u2_u0_n167 ) );
  NAND2_X1 u1_u2_u0_U82 (.A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U83 (.A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U84 (.ZN( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n92 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U85 (.ZN( u1_u2_u0_n142 ) , .A1( u1_u2_u0_n94 ) , .A2( u1_u2_u0_n95 ) );
  INV_X1 u1_u2_u0_U86 (.A( u1_u2_X_3 ) , .ZN( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U87 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n94 ) );
  NAND3_X1 u1_u2_u0_U88 (.ZN( u1_out2_23 ) , .A3( u1_u2_u0_n137 ) , .A1( u1_u2_u0_n168 ) , .A2( u1_u2_u0_n171 ) );
  NAND3_X1 u1_u2_u0_U89 (.A3( u1_u2_u0_n127 ) , .A2( u1_u2_u0_n128 ) , .ZN( u1_u2_u0_n135 ) , .A1( u1_u2_u0_n150 ) );
  AND2_X1 u1_u2_u0_U9 (.A1( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n141 ) , .A2( u1_u2_u0_n150 ) );
  NAND3_X1 u1_u2_u0_U90 (.ZN( u1_u2_u0_n117 ) , .A3( u1_u2_u0_n132 ) , .A2( u1_u2_u0_n139 ) , .A1( u1_u2_u0_n148 ) );
  NAND3_X1 u1_u2_u0_U91 (.ZN( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n114 ) , .A3( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n149 ) );
  NAND3_X1 u1_u2_u0_U92 (.ZN( u1_out2_9 ) , .A3( u1_u2_u0_n106 ) , .A2( u1_u2_u0_n171 ) , .A1( u1_u2_u0_n174 ) );
  NAND3_X1 u1_u2_u0_U93 (.A2( u1_u2_u0_n128 ) , .A1( u1_u2_u0_n132 ) , .A3( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n97 ) );
  OAI22_X1 u1_u2_u4_U10 (.B2( u1_u2_u4_n135 ) , .ZN( u1_u2_u4_n137 ) , .B1( u1_u2_u4_n153 ) , .A1( u1_u2_u4_n155 ) , .A2( u1_u2_u4_n171 ) );
  AND3_X1 u1_u2_u4_U11 (.A2( u1_u2_u4_n134 ) , .ZN( u1_u2_u4_n135 ) , .A3( u1_u2_u4_n145 ) , .A1( u1_u2_u4_n157 ) );
  NAND2_X1 u1_u2_u4_U12 (.ZN( u1_u2_u4_n132 ) , .A2( u1_u2_u4_n170 ) , .A1( u1_u2_u4_n173 ) );
  AOI21_X1 u1_u2_u4_U13 (.B2( u1_u2_u4_n160 ) , .B1( u1_u2_u4_n161 ) , .ZN( u1_u2_u4_n162 ) , .A( u1_u2_u4_n170 ) );
  AOI21_X1 u1_u2_u4_U14 (.ZN( u1_u2_u4_n107 ) , .B2( u1_u2_u4_n143 ) , .A( u1_u2_u4_n174 ) , .B1( u1_u2_u4_n184 ) );
  AOI21_X1 u1_u2_u4_U15 (.B2( u1_u2_u4_n158 ) , .B1( u1_u2_u4_n159 ) , .ZN( u1_u2_u4_n163 ) , .A( u1_u2_u4_n174 ) );
  AOI21_X1 u1_u2_u4_U16 (.A( u1_u2_u4_n153 ) , .B2( u1_u2_u4_n154 ) , .B1( u1_u2_u4_n155 ) , .ZN( u1_u2_u4_n165 ) );
  AOI21_X1 u1_u2_u4_U17 (.A( u1_u2_u4_n156 ) , .B2( u1_u2_u4_n157 ) , .ZN( u1_u2_u4_n164 ) , .B1( u1_u2_u4_n184 ) );
  INV_X1 u1_u2_u4_U18 (.A( u1_u2_u4_n138 ) , .ZN( u1_u2_u4_n170 ) );
  AND2_X1 u1_u2_u4_U19 (.A2( u1_u2_u4_n120 ) , .ZN( u1_u2_u4_n155 ) , .A1( u1_u2_u4_n160 ) );
  INV_X1 u1_u2_u4_U20 (.A( u1_u2_u4_n156 ) , .ZN( u1_u2_u4_n175 ) );
  NAND2_X1 u1_u2_u4_U21 (.A2( u1_u2_u4_n118 ) , .ZN( u1_u2_u4_n131 ) , .A1( u1_u2_u4_n147 ) );
  NAND2_X1 u1_u2_u4_U22 (.A1( u1_u2_u4_n119 ) , .A2( u1_u2_u4_n120 ) , .ZN( u1_u2_u4_n130 ) );
  NAND2_X1 u1_u2_u4_U23 (.ZN( u1_u2_u4_n117 ) , .A2( u1_u2_u4_n118 ) , .A1( u1_u2_u4_n148 ) );
  NAND2_X1 u1_u2_u4_U24 (.ZN( u1_u2_u4_n129 ) , .A1( u1_u2_u4_n134 ) , .A2( u1_u2_u4_n148 ) );
  AND3_X1 u1_u2_u4_U25 (.A1( u1_u2_u4_n119 ) , .A2( u1_u2_u4_n143 ) , .A3( u1_u2_u4_n154 ) , .ZN( u1_u2_u4_n161 ) );
  AND2_X1 u1_u2_u4_U26 (.A1( u1_u2_u4_n145 ) , .A2( u1_u2_u4_n147 ) , .ZN( u1_u2_u4_n159 ) );
  OR3_X1 u1_u2_u4_U27 (.A3( u1_u2_u4_n114 ) , .A2( u1_u2_u4_n115 ) , .A1( u1_u2_u4_n116 ) , .ZN( u1_u2_u4_n136 ) );
  AOI21_X1 u1_u2_u4_U28 (.A( u1_u2_u4_n113 ) , .ZN( u1_u2_u4_n116 ) , .B2( u1_u2_u4_n173 ) , .B1( u1_u2_u4_n174 ) );
  AOI21_X1 u1_u2_u4_U29 (.ZN( u1_u2_u4_n115 ) , .B2( u1_u2_u4_n145 ) , .B1( u1_u2_u4_n146 ) , .A( u1_u2_u4_n156 ) );
  NOR2_X1 u1_u2_u4_U3 (.ZN( u1_u2_u4_n121 ) , .A1( u1_u2_u4_n181 ) , .A2( u1_u2_u4_n182 ) );
  OAI22_X1 u1_u2_u4_U30 (.ZN( u1_u2_u4_n114 ) , .A2( u1_u2_u4_n121 ) , .B1( u1_u2_u4_n160 ) , .B2( u1_u2_u4_n170 ) , .A1( u1_u2_u4_n171 ) );
  INV_X1 u1_u2_u4_U31 (.A( u1_u2_u4_n158 ) , .ZN( u1_u2_u4_n182 ) );
  INV_X1 u1_u2_u4_U32 (.ZN( u1_u2_u4_n181 ) , .A( u1_u2_u4_n96 ) );
  INV_X1 u1_u2_u4_U33 (.A( u1_u2_u4_n144 ) , .ZN( u1_u2_u4_n179 ) );
  INV_X1 u1_u2_u4_U34 (.A( u1_u2_u4_n157 ) , .ZN( u1_u2_u4_n178 ) );
  NAND2_X1 u1_u2_u4_U35 (.A2( u1_u2_u4_n154 ) , .A1( u1_u2_u4_n96 ) , .ZN( u1_u2_u4_n97 ) );
  INV_X1 u1_u2_u4_U36 (.ZN( u1_u2_u4_n186 ) , .A( u1_u2_u4_n95 ) );
  OAI221_X1 u1_u2_u4_U37 (.C1( u1_u2_u4_n134 ) , .B1( u1_u2_u4_n158 ) , .B2( u1_u2_u4_n171 ) , .C2( u1_u2_u4_n173 ) , .A( u1_u2_u4_n94 ) , .ZN( u1_u2_u4_n95 ) );
  AOI222_X1 u1_u2_u4_U38 (.B2( u1_u2_u4_n132 ) , .A1( u1_u2_u4_n138 ) , .C2( u1_u2_u4_n175 ) , .A2( u1_u2_u4_n179 ) , .C1( u1_u2_u4_n181 ) , .B1( u1_u2_u4_n185 ) , .ZN( u1_u2_u4_n94 ) );
  INV_X1 u1_u2_u4_U39 (.A( u1_u2_u4_n113 ) , .ZN( u1_u2_u4_n185 ) );
  INV_X1 u1_u2_u4_U4 (.A( u1_u2_u4_n117 ) , .ZN( u1_u2_u4_n184 ) );
  INV_X1 u1_u2_u4_U40 (.A( u1_u2_u4_n143 ) , .ZN( u1_u2_u4_n183 ) );
  NOR2_X1 u1_u2_u4_U41 (.ZN( u1_u2_u4_n138 ) , .A1( u1_u2_u4_n168 ) , .A2( u1_u2_u4_n169 ) );
  NOR2_X1 u1_u2_u4_U42 (.A1( u1_u2_u4_n150 ) , .A2( u1_u2_u4_n152 ) , .ZN( u1_u2_u4_n153 ) );
  NOR2_X1 u1_u2_u4_U43 (.A2( u1_u2_u4_n128 ) , .A1( u1_u2_u4_n138 ) , .ZN( u1_u2_u4_n156 ) );
  AOI22_X1 u1_u2_u4_U44 (.B2( u1_u2_u4_n122 ) , .A1( u1_u2_u4_n123 ) , .ZN( u1_u2_u4_n124 ) , .B1( u1_u2_u4_n128 ) , .A2( u1_u2_u4_n172 ) );
  INV_X1 u1_u2_u4_U45 (.A( u1_u2_u4_n153 ) , .ZN( u1_u2_u4_n172 ) );
  NAND2_X1 u1_u2_u4_U46 (.A2( u1_u2_u4_n120 ) , .ZN( u1_u2_u4_n123 ) , .A1( u1_u2_u4_n161 ) );
  AOI22_X1 u1_u2_u4_U47 (.B2( u1_u2_u4_n132 ) , .A2( u1_u2_u4_n133 ) , .ZN( u1_u2_u4_n140 ) , .A1( u1_u2_u4_n150 ) , .B1( u1_u2_u4_n179 ) );
  NAND2_X1 u1_u2_u4_U48 (.ZN( u1_u2_u4_n133 ) , .A2( u1_u2_u4_n146 ) , .A1( u1_u2_u4_n154 ) );
  NAND2_X1 u1_u2_u4_U49 (.A1( u1_u2_u4_n103 ) , .ZN( u1_u2_u4_n154 ) , .A2( u1_u2_u4_n98 ) );
  NOR4_X1 u1_u2_u4_U5 (.A4( u1_u2_u4_n106 ) , .A3( u1_u2_u4_n107 ) , .A2( u1_u2_u4_n108 ) , .A1( u1_u2_u4_n109 ) , .ZN( u1_u2_u4_n110 ) );
  NAND2_X1 u1_u2_u4_U50 (.A1( u1_u2_u4_n101 ) , .ZN( u1_u2_u4_n158 ) , .A2( u1_u2_u4_n99 ) );
  AOI21_X1 u1_u2_u4_U51 (.ZN( u1_u2_u4_n127 ) , .A( u1_u2_u4_n136 ) , .B2( u1_u2_u4_n150 ) , .B1( u1_u2_u4_n180 ) );
  INV_X1 u1_u2_u4_U52 (.A( u1_u2_u4_n160 ) , .ZN( u1_u2_u4_n180 ) );
  NAND2_X1 u1_u2_u4_U53 (.A2( u1_u2_u4_n104 ) , .A1( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n146 ) );
  NAND2_X1 u1_u2_u4_U54 (.A2( u1_u2_u4_n101 ) , .A1( u1_u2_u4_n102 ) , .ZN( u1_u2_u4_n160 ) );
  NAND2_X1 u1_u2_u4_U55 (.ZN( u1_u2_u4_n134 ) , .A1( u1_u2_u4_n98 ) , .A2( u1_u2_u4_n99 ) );
  NAND2_X1 u1_u2_u4_U56 (.A1( u1_u2_u4_n103 ) , .A2( u1_u2_u4_n104 ) , .ZN( u1_u2_u4_n143 ) );
  NAND2_X1 u1_u2_u4_U57 (.A2( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n145 ) , .A1( u1_u2_u4_n98 ) );
  NAND2_X1 u1_u2_u4_U58 (.A1( u1_u2_u4_n100 ) , .A2( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n120 ) );
  NAND2_X1 u1_u2_u4_U59 (.A1( u1_u2_u4_n102 ) , .A2( u1_u2_u4_n104 ) , .ZN( u1_u2_u4_n148 ) );
  AOI21_X1 u1_u2_u4_U6 (.ZN( u1_u2_u4_n106 ) , .B2( u1_u2_u4_n146 ) , .B1( u1_u2_u4_n158 ) , .A( u1_u2_u4_n170 ) );
  NAND2_X1 u1_u2_u4_U60 (.A2( u1_u2_u4_n100 ) , .A1( u1_u2_u4_n103 ) , .ZN( u1_u2_u4_n157 ) );
  INV_X1 u1_u2_u4_U61 (.A( u1_u2_u4_n150 ) , .ZN( u1_u2_u4_n173 ) );
  INV_X1 u1_u2_u4_U62 (.A( u1_u2_u4_n152 ) , .ZN( u1_u2_u4_n171 ) );
  NAND2_X1 u1_u2_u4_U63 (.A1( u1_u2_u4_n100 ) , .ZN( u1_u2_u4_n118 ) , .A2( u1_u2_u4_n99 ) );
  NAND2_X1 u1_u2_u4_U64 (.A2( u1_u2_u4_n100 ) , .A1( u1_u2_u4_n102 ) , .ZN( u1_u2_u4_n144 ) );
  NAND2_X1 u1_u2_u4_U65 (.A2( u1_u2_u4_n101 ) , .A1( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n96 ) );
  INV_X1 u1_u2_u4_U66 (.A( u1_u2_u4_n128 ) , .ZN( u1_u2_u4_n174 ) );
  NAND2_X1 u1_u2_u4_U67 (.A2( u1_u2_u4_n102 ) , .ZN( u1_u2_u4_n119 ) , .A1( u1_u2_u4_n98 ) );
  NAND2_X1 u1_u2_u4_U68 (.A2( u1_u2_u4_n101 ) , .A1( u1_u2_u4_n103 ) , .ZN( u1_u2_u4_n147 ) );
  NAND2_X1 u1_u2_u4_U69 (.A2( u1_u2_u4_n104 ) , .ZN( u1_u2_u4_n113 ) , .A1( u1_u2_u4_n99 ) );
  AOI21_X1 u1_u2_u4_U7 (.ZN( u1_u2_u4_n108 ) , .B2( u1_u2_u4_n134 ) , .B1( u1_u2_u4_n155 ) , .A( u1_u2_u4_n156 ) );
  NOR2_X1 u1_u2_u4_U70 (.A2( u1_u2_X_28 ) , .ZN( u1_u2_u4_n150 ) , .A1( u1_u2_u4_n168 ) );
  NOR2_X1 u1_u2_u4_U71 (.A2( u1_u2_X_29 ) , .ZN( u1_u2_u4_n152 ) , .A1( u1_u2_u4_n169 ) );
  NOR2_X1 u1_u2_u4_U72 (.A2( u1_u2_X_30 ) , .ZN( u1_u2_u4_n105 ) , .A1( u1_u2_u4_n176 ) );
  NOR2_X1 u1_u2_u4_U73 (.A2( u1_u2_X_26 ) , .ZN( u1_u2_u4_n100 ) , .A1( u1_u2_u4_n177 ) );
  NOR2_X1 u1_u2_u4_U74 (.A2( u1_u2_X_28 ) , .A1( u1_u2_X_29 ) , .ZN( u1_u2_u4_n128 ) );
  NOR2_X1 u1_u2_u4_U75 (.A2( u1_u2_X_27 ) , .A1( u1_u2_X_30 ) , .ZN( u1_u2_u4_n102 ) );
  NOR2_X1 u1_u2_u4_U76 (.A2( u1_u2_X_25 ) , .A1( u1_u2_X_26 ) , .ZN( u1_u2_u4_n98 ) );
  AND2_X1 u1_u2_u4_U77 (.A2( u1_u2_X_25 ) , .A1( u1_u2_X_26 ) , .ZN( u1_u2_u4_n104 ) );
  AND2_X1 u1_u2_u4_U78 (.A1( u1_u2_X_30 ) , .A2( u1_u2_u4_n176 ) , .ZN( u1_u2_u4_n99 ) );
  AND2_X1 u1_u2_u4_U79 (.A1( u1_u2_X_26 ) , .ZN( u1_u2_u4_n101 ) , .A2( u1_u2_u4_n177 ) );
  AOI21_X1 u1_u2_u4_U8 (.ZN( u1_u2_u4_n109 ) , .A( u1_u2_u4_n153 ) , .B1( u1_u2_u4_n159 ) , .B2( u1_u2_u4_n184 ) );
  AND2_X1 u1_u2_u4_U80 (.A1( u1_u2_X_27 ) , .A2( u1_u2_X_30 ) , .ZN( u1_u2_u4_n103 ) );
  INV_X1 u1_u2_u4_U81 (.A( u1_u2_X_28 ) , .ZN( u1_u2_u4_n169 ) );
  INV_X1 u1_u2_u4_U82 (.A( u1_u2_X_29 ) , .ZN( u1_u2_u4_n168 ) );
  INV_X1 u1_u2_u4_U83 (.A( u1_u2_X_25 ) , .ZN( u1_u2_u4_n177 ) );
  INV_X1 u1_u2_u4_U84 (.A( u1_u2_X_27 ) , .ZN( u1_u2_u4_n176 ) );
  NAND4_X1 u1_u2_u4_U85 (.ZN( u1_out2_25 ) , .A4( u1_u2_u4_n139 ) , .A3( u1_u2_u4_n140 ) , .A2( u1_u2_u4_n141 ) , .A1( u1_u2_u4_n142 ) );
  OAI21_X1 u1_u2_u4_U86 (.A( u1_u2_u4_n128 ) , .B2( u1_u2_u4_n129 ) , .B1( u1_u2_u4_n130 ) , .ZN( u1_u2_u4_n142 ) );
  OAI21_X1 u1_u2_u4_U87 (.B2( u1_u2_u4_n131 ) , .ZN( u1_u2_u4_n141 ) , .A( u1_u2_u4_n175 ) , .B1( u1_u2_u4_n183 ) );
  NAND4_X1 u1_u2_u4_U88 (.ZN( u1_out2_14 ) , .A4( u1_u2_u4_n124 ) , .A3( u1_u2_u4_n125 ) , .A2( u1_u2_u4_n126 ) , .A1( u1_u2_u4_n127 ) );
  AOI22_X1 u1_u2_u4_U89 (.B2( u1_u2_u4_n117 ) , .ZN( u1_u2_u4_n126 ) , .A1( u1_u2_u4_n129 ) , .B1( u1_u2_u4_n152 ) , .A2( u1_u2_u4_n175 ) );
  AOI211_X1 u1_u2_u4_U9 (.B( u1_u2_u4_n136 ) , .A( u1_u2_u4_n137 ) , .C2( u1_u2_u4_n138 ) , .ZN( u1_u2_u4_n139 ) , .C1( u1_u2_u4_n182 ) );
  AOI22_X1 u1_u2_u4_U90 (.ZN( u1_u2_u4_n125 ) , .B2( u1_u2_u4_n131 ) , .A2( u1_u2_u4_n132 ) , .B1( u1_u2_u4_n138 ) , .A1( u1_u2_u4_n178 ) );
  NAND4_X1 u1_u2_u4_U91 (.ZN( u1_out2_8 ) , .A4( u1_u2_u4_n110 ) , .A3( u1_u2_u4_n111 ) , .A2( u1_u2_u4_n112 ) , .A1( u1_u2_u4_n186 ) );
  NAND2_X1 u1_u2_u4_U92 (.ZN( u1_u2_u4_n112 ) , .A2( u1_u2_u4_n130 ) , .A1( u1_u2_u4_n150 ) );
  AOI22_X1 u1_u2_u4_U93 (.ZN( u1_u2_u4_n111 ) , .B2( u1_u2_u4_n132 ) , .A1( u1_u2_u4_n152 ) , .B1( u1_u2_u4_n178 ) , .A2( u1_u2_u4_n97 ) );
  AOI22_X1 u1_u2_u4_U94 (.B2( u1_u2_u4_n149 ) , .B1( u1_u2_u4_n150 ) , .A2( u1_u2_u4_n151 ) , .A1( u1_u2_u4_n152 ) , .ZN( u1_u2_u4_n167 ) );
  NOR4_X1 u1_u2_u4_U95 (.A4( u1_u2_u4_n162 ) , .A3( u1_u2_u4_n163 ) , .A2( u1_u2_u4_n164 ) , .A1( u1_u2_u4_n165 ) , .ZN( u1_u2_u4_n166 ) );
  NAND3_X1 u1_u2_u4_U96 (.ZN( u1_out2_3 ) , .A3( u1_u2_u4_n166 ) , .A1( u1_u2_u4_n167 ) , .A2( u1_u2_u4_n186 ) );
  NAND3_X1 u1_u2_u4_U97 (.A3( u1_u2_u4_n146 ) , .A2( u1_u2_u4_n147 ) , .A1( u1_u2_u4_n148 ) , .ZN( u1_u2_u4_n149 ) );
  NAND3_X1 u1_u2_u4_U98 (.A3( u1_u2_u4_n143 ) , .A2( u1_u2_u4_n144 ) , .A1( u1_u2_u4_n145 ) , .ZN( u1_u2_u4_n151 ) );
  NAND3_X1 u1_u2_u4_U99 (.A3( u1_u2_u4_n121 ) , .ZN( u1_u2_u4_n122 ) , .A2( u1_u2_u4_n144 ) , .A1( u1_u2_u4_n154 ) );
  XOR2_X1 u1_u3_U10 (.B( u1_K4_45 ) , .A( u1_R2_30 ) , .Z( u1_u3_X_45 ) );
  XOR2_X1 u1_u3_U22 (.B( u1_K4_34 ) , .A( u1_R2_23 ) , .Z( u1_u3_X_34 ) );
  XOR2_X1 u1_u3_U23 (.B( u1_K4_33 ) , .A( u1_R2_22 ) , .Z( u1_u3_X_33 ) );
  XOR2_X1 u1_u3_U24 (.B( u1_K4_32 ) , .A( u1_R2_21 ) , .Z( u1_u3_X_32 ) );
  XOR2_X1 u1_u3_U25 (.B( u1_K4_31 ) , .A( u1_R2_20 ) , .Z( u1_u3_X_31 ) );
  XOR2_X1 u1_u3_U26 (.B( u1_K4_30 ) , .A( u1_R2_21 ) , .Z( u1_u3_X_30 ) );
  XOR2_X1 u1_u3_U28 (.B( u1_K4_29 ) , .A( u1_R2_20 ) , .Z( u1_u3_X_29 ) );
  XOR2_X1 u1_u3_U29 (.B( u1_K4_28 ) , .A( u1_R2_19 ) , .Z( u1_u3_X_28 ) );
  XOR2_X1 u1_u3_U30 (.B( u1_K4_27 ) , .A( u1_R2_18 ) , .Z( u1_u3_X_27 ) );
  XOR2_X1 u1_u3_U42 (.B( u1_K4_16 ) , .A( u1_R2_11 ) , .Z( u1_u3_X_16 ) );
  XOR2_X1 u1_u3_U43 (.B( u1_K4_15 ) , .A( u1_R2_10 ) , .Z( u1_u3_X_15 ) );
  XOR2_X1 u1_u3_U9 (.B( u1_K4_46 ) , .A( u1_R2_31 ) , .Z( u1_u3_X_46 ) );
  OAI22_X1 u1_u3_u2_U10 (.B1( u1_u3_u2_n151 ) , .A2( u1_u3_u2_n152 ) , .A1( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n160 ) , .B2( u1_u3_u2_n168 ) );
  NAND3_X1 u1_u3_u2_U100 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n104 ) , .A3( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n98 ) );
  NOR3_X1 u1_u3_u2_U11 (.A1( u1_u3_u2_n150 ) , .ZN( u1_u3_u2_n151 ) , .A3( u1_u3_u2_n175 ) , .A2( u1_u3_u2_n188 ) );
  AOI21_X1 u1_u3_u2_U12 (.B2( u1_u3_u2_n123 ) , .ZN( u1_u3_u2_n125 ) , .A( u1_u3_u2_n171 ) , .B1( u1_u3_u2_n184 ) );
  INV_X1 u1_u3_u2_U13 (.A( u1_u3_u2_n150 ) , .ZN( u1_u3_u2_n184 ) );
  AOI21_X1 u1_u3_u2_U14 (.ZN( u1_u3_u2_n144 ) , .B2( u1_u3_u2_n155 ) , .A( u1_u3_u2_n172 ) , .B1( u1_u3_u2_n185 ) );
  AOI21_X1 u1_u3_u2_U15 (.B2( u1_u3_u2_n143 ) , .ZN( u1_u3_u2_n145 ) , .B1( u1_u3_u2_n152 ) , .A( u1_u3_u2_n171 ) );
  INV_X1 u1_u3_u2_U16 (.A( u1_u3_u2_n156 ) , .ZN( u1_u3_u2_n171 ) );
  INV_X1 u1_u3_u2_U17 (.A( u1_u3_u2_n120 ) , .ZN( u1_u3_u2_n188 ) );
  NAND2_X1 u1_u3_u2_U18 (.A2( u1_u3_u2_n122 ) , .ZN( u1_u3_u2_n150 ) , .A1( u1_u3_u2_n152 ) );
  INV_X1 u1_u3_u2_U19 (.A( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n170 ) );
  INV_X1 u1_u3_u2_U20 (.A( u1_u3_u2_n137 ) , .ZN( u1_u3_u2_n173 ) );
  NAND2_X1 u1_u3_u2_U21 (.A1( u1_u3_u2_n132 ) , .A2( u1_u3_u2_n139 ) , .ZN( u1_u3_u2_n157 ) );
  INV_X1 u1_u3_u2_U22 (.A( u1_u3_u2_n113 ) , .ZN( u1_u3_u2_n178 ) );
  INV_X1 u1_u3_u2_U23 (.A( u1_u3_u2_n139 ) , .ZN( u1_u3_u2_n175 ) );
  INV_X1 u1_u3_u2_U24 (.A( u1_u3_u2_n155 ) , .ZN( u1_u3_u2_n181 ) );
  INV_X1 u1_u3_u2_U25 (.A( u1_u3_u2_n119 ) , .ZN( u1_u3_u2_n177 ) );
  INV_X1 u1_u3_u2_U26 (.A( u1_u3_u2_n116 ) , .ZN( u1_u3_u2_n180 ) );
  INV_X1 u1_u3_u2_U27 (.A( u1_u3_u2_n131 ) , .ZN( u1_u3_u2_n179 ) );
  INV_X1 u1_u3_u2_U28 (.A( u1_u3_u2_n154 ) , .ZN( u1_u3_u2_n176 ) );
  NAND2_X1 u1_u3_u2_U29 (.A2( u1_u3_u2_n116 ) , .A1( u1_u3_u2_n117 ) , .ZN( u1_u3_u2_n118 ) );
  NOR2_X1 u1_u3_u2_U3 (.ZN( u1_u3_u2_n121 ) , .A2( u1_u3_u2_n177 ) , .A1( u1_u3_u2_n180 ) );
  INV_X1 u1_u3_u2_U30 (.A( u1_u3_u2_n132 ) , .ZN( u1_u3_u2_n182 ) );
  INV_X1 u1_u3_u2_U31 (.A( u1_u3_u2_n158 ) , .ZN( u1_u3_u2_n183 ) );
  OAI21_X1 u1_u3_u2_U32 (.A( u1_u3_u2_n156 ) , .B1( u1_u3_u2_n157 ) , .ZN( u1_u3_u2_n158 ) , .B2( u1_u3_u2_n179 ) );
  NOR2_X1 u1_u3_u2_U33 (.ZN( u1_u3_u2_n156 ) , .A1( u1_u3_u2_n166 ) , .A2( u1_u3_u2_n169 ) );
  NOR2_X1 u1_u3_u2_U34 (.A2( u1_u3_u2_n114 ) , .ZN( u1_u3_u2_n137 ) , .A1( u1_u3_u2_n140 ) );
  NOR2_X1 u1_u3_u2_U35 (.A2( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n153 ) , .A1( u1_u3_u2_n156 ) );
  AOI211_X1 u1_u3_u2_U36 (.ZN( u1_u3_u2_n130 ) , .C1( u1_u3_u2_n138 ) , .C2( u1_u3_u2_n179 ) , .B( u1_u3_u2_n96 ) , .A( u1_u3_u2_n97 ) );
  OAI22_X1 u1_u3_u2_U37 (.B1( u1_u3_u2_n133 ) , .A2( u1_u3_u2_n137 ) , .A1( u1_u3_u2_n152 ) , .B2( u1_u3_u2_n168 ) , .ZN( u1_u3_u2_n97 ) );
  OAI221_X1 u1_u3_u2_U38 (.B1( u1_u3_u2_n113 ) , .C1( u1_u3_u2_n132 ) , .A( u1_u3_u2_n149 ) , .B2( u1_u3_u2_n171 ) , .C2( u1_u3_u2_n172 ) , .ZN( u1_u3_u2_n96 ) );
  OAI221_X1 u1_u3_u2_U39 (.A( u1_u3_u2_n115 ) , .C2( u1_u3_u2_n123 ) , .B2( u1_u3_u2_n143 ) , .B1( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n163 ) , .C1( u1_u3_u2_n168 ) );
  INV_X1 u1_u3_u2_U4 (.A( u1_u3_u2_n134 ) , .ZN( u1_u3_u2_n185 ) );
  OAI21_X1 u1_u3_u2_U40 (.A( u1_u3_u2_n114 ) , .ZN( u1_u3_u2_n115 ) , .B1( u1_u3_u2_n176 ) , .B2( u1_u3_u2_n178 ) );
  OAI221_X1 u1_u3_u2_U41 (.A( u1_u3_u2_n135 ) , .B2( u1_u3_u2_n136 ) , .B1( u1_u3_u2_n137 ) , .ZN( u1_u3_u2_n162 ) , .C2( u1_u3_u2_n167 ) , .C1( u1_u3_u2_n185 ) );
  AND3_X1 u1_u3_u2_U42 (.A3( u1_u3_u2_n131 ) , .A2( u1_u3_u2_n132 ) , .A1( u1_u3_u2_n133 ) , .ZN( u1_u3_u2_n136 ) );
  AOI22_X1 u1_u3_u2_U43 (.ZN( u1_u3_u2_n135 ) , .B1( u1_u3_u2_n140 ) , .A1( u1_u3_u2_n156 ) , .B2( u1_u3_u2_n180 ) , .A2( u1_u3_u2_n188 ) );
  AOI21_X1 u1_u3_u2_U44 (.ZN( u1_u3_u2_n149 ) , .B1( u1_u3_u2_n173 ) , .B2( u1_u3_u2_n188 ) , .A( u1_u3_u2_n95 ) );
  AND3_X1 u1_u3_u2_U45 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n104 ) , .A3( u1_u3_u2_n156 ) , .ZN( u1_u3_u2_n95 ) );
  OAI21_X1 u1_u3_u2_U46 (.A( u1_u3_u2_n101 ) , .B2( u1_u3_u2_n121 ) , .B1( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n164 ) );
  NAND2_X1 u1_u3_u2_U47 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n107 ) , .ZN( u1_u3_u2_n155 ) );
  NAND2_X1 u1_u3_u2_U48 (.A2( u1_u3_u2_n105 ) , .A1( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n143 ) );
  NAND2_X1 u1_u3_u2_U49 (.A1( u1_u3_u2_n104 ) , .A2( u1_u3_u2_n106 ) , .ZN( u1_u3_u2_n152 ) );
  NOR4_X1 u1_u3_u2_U5 (.A4( u1_u3_u2_n124 ) , .A3( u1_u3_u2_n125 ) , .A2( u1_u3_u2_n126 ) , .A1( u1_u3_u2_n127 ) , .ZN( u1_u3_u2_n128 ) );
  NAND2_X1 u1_u3_u2_U50 (.A1( u1_u3_u2_n100 ) , .A2( u1_u3_u2_n105 ) , .ZN( u1_u3_u2_n132 ) );
  INV_X1 u1_u3_u2_U51 (.A( u1_u3_u2_n140 ) , .ZN( u1_u3_u2_n168 ) );
  INV_X1 u1_u3_u2_U52 (.A( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n167 ) );
  OAI21_X1 u1_u3_u2_U53 (.A( u1_u3_u2_n141 ) , .B2( u1_u3_u2_n142 ) , .ZN( u1_u3_u2_n146 ) , .B1( u1_u3_u2_n153 ) );
  OAI21_X1 u1_u3_u2_U54 (.A( u1_u3_u2_n140 ) , .ZN( u1_u3_u2_n141 ) , .B1( u1_u3_u2_n176 ) , .B2( u1_u3_u2_n177 ) );
  NOR3_X1 u1_u3_u2_U55 (.ZN( u1_u3_u2_n142 ) , .A3( u1_u3_u2_n175 ) , .A2( u1_u3_u2_n178 ) , .A1( u1_u3_u2_n181 ) );
  INV_X1 u1_u3_u2_U56 (.ZN( u1_u3_u2_n187 ) , .A( u1_u3_u2_n99 ) );
  OAI21_X1 u1_u3_u2_U57 (.B1( u1_u3_u2_n137 ) , .B2( u1_u3_u2_n143 ) , .A( u1_u3_u2_n98 ) , .ZN( u1_u3_u2_n99 ) );
  NAND2_X1 u1_u3_u2_U58 (.A1( u1_u3_u2_n102 ) , .A2( u1_u3_u2_n106 ) , .ZN( u1_u3_u2_n113 ) );
  NAND2_X1 u1_u3_u2_U59 (.A1( u1_u3_u2_n106 ) , .A2( u1_u3_u2_n107 ) , .ZN( u1_u3_u2_n131 ) );
  AOI21_X1 u1_u3_u2_U6 (.B2( u1_u3_u2_n119 ) , .ZN( u1_u3_u2_n127 ) , .A( u1_u3_u2_n137 ) , .B1( u1_u3_u2_n155 ) );
  NAND2_X1 u1_u3_u2_U60 (.A1( u1_u3_u2_n103 ) , .A2( u1_u3_u2_n107 ) , .ZN( u1_u3_u2_n139 ) );
  NAND2_X1 u1_u3_u2_U61 (.A1( u1_u3_u2_n103 ) , .A2( u1_u3_u2_n105 ) , .ZN( u1_u3_u2_n133 ) );
  NAND2_X1 u1_u3_u2_U62 (.A1( u1_u3_u2_n102 ) , .A2( u1_u3_u2_n103 ) , .ZN( u1_u3_u2_n154 ) );
  NAND2_X1 u1_u3_u2_U63 (.A2( u1_u3_u2_n103 ) , .A1( u1_u3_u2_n104 ) , .ZN( u1_u3_u2_n119 ) );
  NAND2_X1 u1_u3_u2_U64 (.A2( u1_u3_u2_n107 ) , .A1( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n123 ) );
  NAND2_X1 u1_u3_u2_U65 (.A1( u1_u3_u2_n104 ) , .A2( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n122 ) );
  INV_X1 u1_u3_u2_U66 (.A( u1_u3_u2_n114 ) , .ZN( u1_u3_u2_n172 ) );
  NAND2_X1 u1_u3_u2_U67 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n102 ) , .ZN( u1_u3_u2_n116 ) );
  NAND2_X1 u1_u3_u2_U68 (.A1( u1_u3_u2_n102 ) , .A2( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n120 ) );
  NAND2_X1 u1_u3_u2_U69 (.A2( u1_u3_u2_n105 ) , .A1( u1_u3_u2_n106 ) , .ZN( u1_u3_u2_n117 ) );
  AOI21_X1 u1_u3_u2_U7 (.ZN( u1_u3_u2_n124 ) , .B1( u1_u3_u2_n131 ) , .B2( u1_u3_u2_n143 ) , .A( u1_u3_u2_n172 ) );
  NOR2_X1 u1_u3_u2_U70 (.A2( u1_u3_X_16 ) , .ZN( u1_u3_u2_n140 ) , .A1( u1_u3_u2_n166 ) );
  NOR2_X1 u1_u3_u2_U71 (.A2( u1_u3_X_13 ) , .A1( u1_u3_X_14 ) , .ZN( u1_u3_u2_n100 ) );
  NOR2_X1 u1_u3_u2_U72 (.A2( u1_u3_X_16 ) , .A1( u1_u3_X_17 ) , .ZN( u1_u3_u2_n138 ) );
  NOR2_X1 u1_u3_u2_U73 (.A2( u1_u3_X_15 ) , .A1( u1_u3_X_18 ) , .ZN( u1_u3_u2_n104 ) );
  NOR2_X1 u1_u3_u2_U74 (.A2( u1_u3_X_14 ) , .ZN( u1_u3_u2_n103 ) , .A1( u1_u3_u2_n174 ) );
  NOR2_X1 u1_u3_u2_U75 (.A2( u1_u3_X_15 ) , .ZN( u1_u3_u2_n102 ) , .A1( u1_u3_u2_n165 ) );
  NOR2_X1 u1_u3_u2_U76 (.A2( u1_u3_X_17 ) , .ZN( u1_u3_u2_n114 ) , .A1( u1_u3_u2_n169 ) );
  AND2_X1 u1_u3_u2_U77 (.A1( u1_u3_X_15 ) , .ZN( u1_u3_u2_n105 ) , .A2( u1_u3_u2_n165 ) );
  AND2_X1 u1_u3_u2_U78 (.A2( u1_u3_X_15 ) , .A1( u1_u3_X_18 ) , .ZN( u1_u3_u2_n107 ) );
  AND2_X1 u1_u3_u2_U79 (.A1( u1_u3_X_14 ) , .ZN( u1_u3_u2_n106 ) , .A2( u1_u3_u2_n174 ) );
  AOI21_X1 u1_u3_u2_U8 (.B2( u1_u3_u2_n120 ) , .B1( u1_u3_u2_n121 ) , .ZN( u1_u3_u2_n126 ) , .A( u1_u3_u2_n167 ) );
  AND2_X1 u1_u3_u2_U80 (.A1( u1_u3_X_13 ) , .A2( u1_u3_X_14 ) , .ZN( u1_u3_u2_n108 ) );
  INV_X1 u1_u3_u2_U81 (.A( u1_u3_X_16 ) , .ZN( u1_u3_u2_n169 ) );
  INV_X1 u1_u3_u2_U82 (.A( u1_u3_X_17 ) , .ZN( u1_u3_u2_n166 ) );
  INV_X1 u1_u3_u2_U83 (.A( u1_u3_X_13 ) , .ZN( u1_u3_u2_n174 ) );
  INV_X1 u1_u3_u2_U84 (.A( u1_u3_X_18 ) , .ZN( u1_u3_u2_n165 ) );
  NAND4_X1 u1_u3_u2_U85 (.ZN( u1_out3_30 ) , .A4( u1_u3_u2_n147 ) , .A3( u1_u3_u2_n148 ) , .A2( u1_u3_u2_n149 ) , .A1( u1_u3_u2_n187 ) );
  AOI21_X1 u1_u3_u2_U86 (.B2( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n148 ) , .A( u1_u3_u2_n162 ) , .B1( u1_u3_u2_n182 ) );
  NOR3_X1 u1_u3_u2_U87 (.A3( u1_u3_u2_n144 ) , .A2( u1_u3_u2_n145 ) , .A1( u1_u3_u2_n146 ) , .ZN( u1_u3_u2_n147 ) );
  NAND4_X1 u1_u3_u2_U88 (.ZN( u1_out3_24 ) , .A4( u1_u3_u2_n111 ) , .A3( u1_u3_u2_n112 ) , .A1( u1_u3_u2_n130 ) , .A2( u1_u3_u2_n187 ) );
  AOI221_X1 u1_u3_u2_U89 (.A( u1_u3_u2_n109 ) , .B1( u1_u3_u2_n110 ) , .ZN( u1_u3_u2_n111 ) , .C1( u1_u3_u2_n134 ) , .C2( u1_u3_u2_n170 ) , .B2( u1_u3_u2_n173 ) );
  OAI22_X1 u1_u3_u2_U9 (.ZN( u1_u3_u2_n109 ) , .A2( u1_u3_u2_n113 ) , .B2( u1_u3_u2_n133 ) , .B1( u1_u3_u2_n167 ) , .A1( u1_u3_u2_n168 ) );
  AOI21_X1 u1_u3_u2_U90 (.ZN( u1_u3_u2_n112 ) , .B2( u1_u3_u2_n156 ) , .A( u1_u3_u2_n164 ) , .B1( u1_u3_u2_n181 ) );
  NAND4_X1 u1_u3_u2_U91 (.ZN( u1_out3_16 ) , .A4( u1_u3_u2_n128 ) , .A3( u1_u3_u2_n129 ) , .A1( u1_u3_u2_n130 ) , .A2( u1_u3_u2_n186 ) );
  AOI22_X1 u1_u3_u2_U92 (.A2( u1_u3_u2_n118 ) , .ZN( u1_u3_u2_n129 ) , .A1( u1_u3_u2_n140 ) , .B1( u1_u3_u2_n157 ) , .B2( u1_u3_u2_n170 ) );
  INV_X1 u1_u3_u2_U93 (.A( u1_u3_u2_n163 ) , .ZN( u1_u3_u2_n186 ) );
  OR4_X1 u1_u3_u2_U94 (.ZN( u1_out3_6 ) , .A4( u1_u3_u2_n161 ) , .A3( u1_u3_u2_n162 ) , .A2( u1_u3_u2_n163 ) , .A1( u1_u3_u2_n164 ) );
  OR3_X1 u1_u3_u2_U95 (.A2( u1_u3_u2_n159 ) , .A1( u1_u3_u2_n160 ) , .ZN( u1_u3_u2_n161 ) , .A3( u1_u3_u2_n183 ) );
  AOI21_X1 u1_u3_u2_U96 (.B2( u1_u3_u2_n154 ) , .B1( u1_u3_u2_n155 ) , .ZN( u1_u3_u2_n159 ) , .A( u1_u3_u2_n167 ) );
  NAND3_X1 u1_u3_u2_U97 (.A2( u1_u3_u2_n117 ) , .A1( u1_u3_u2_n122 ) , .A3( u1_u3_u2_n123 ) , .ZN( u1_u3_u2_n134 ) );
  NAND3_X1 u1_u3_u2_U98 (.ZN( u1_u3_u2_n110 ) , .A2( u1_u3_u2_n131 ) , .A3( u1_u3_u2_n139 ) , .A1( u1_u3_u2_n154 ) );
  NAND3_X1 u1_u3_u2_U99 (.A2( u1_u3_u2_n100 ) , .ZN( u1_u3_u2_n101 ) , .A1( u1_u3_u2_n104 ) , .A3( u1_u3_u2_n114 ) );
  OAI22_X1 u1_u3_u4_U10 (.B2( u1_u3_u4_n135 ) , .ZN( u1_u3_u4_n137 ) , .B1( u1_u3_u4_n153 ) , .A1( u1_u3_u4_n155 ) , .A2( u1_u3_u4_n171 ) );
  AND3_X1 u1_u3_u4_U11 (.A2( u1_u3_u4_n134 ) , .ZN( u1_u3_u4_n135 ) , .A3( u1_u3_u4_n145 ) , .A1( u1_u3_u4_n157 ) );
  NAND2_X1 u1_u3_u4_U12 (.ZN( u1_u3_u4_n132 ) , .A2( u1_u3_u4_n170 ) , .A1( u1_u3_u4_n173 ) );
  AOI21_X1 u1_u3_u4_U13 (.B2( u1_u3_u4_n160 ) , .B1( u1_u3_u4_n161 ) , .ZN( u1_u3_u4_n162 ) , .A( u1_u3_u4_n170 ) );
  AOI21_X1 u1_u3_u4_U14 (.ZN( u1_u3_u4_n107 ) , .B2( u1_u3_u4_n143 ) , .A( u1_u3_u4_n174 ) , .B1( u1_u3_u4_n184 ) );
  AOI21_X1 u1_u3_u4_U15 (.B2( u1_u3_u4_n158 ) , .B1( u1_u3_u4_n159 ) , .ZN( u1_u3_u4_n163 ) , .A( u1_u3_u4_n174 ) );
  AOI21_X1 u1_u3_u4_U16 (.A( u1_u3_u4_n153 ) , .B2( u1_u3_u4_n154 ) , .B1( u1_u3_u4_n155 ) , .ZN( u1_u3_u4_n165 ) );
  AOI21_X1 u1_u3_u4_U17 (.A( u1_u3_u4_n156 ) , .B2( u1_u3_u4_n157 ) , .ZN( u1_u3_u4_n164 ) , .B1( u1_u3_u4_n184 ) );
  INV_X1 u1_u3_u4_U18 (.A( u1_u3_u4_n138 ) , .ZN( u1_u3_u4_n170 ) );
  AND2_X1 u1_u3_u4_U19 (.A2( u1_u3_u4_n120 ) , .ZN( u1_u3_u4_n155 ) , .A1( u1_u3_u4_n160 ) );
  INV_X1 u1_u3_u4_U20 (.A( u1_u3_u4_n156 ) , .ZN( u1_u3_u4_n175 ) );
  NAND2_X1 u1_u3_u4_U21 (.A2( u1_u3_u4_n118 ) , .ZN( u1_u3_u4_n131 ) , .A1( u1_u3_u4_n147 ) );
  NAND2_X1 u1_u3_u4_U22 (.A1( u1_u3_u4_n119 ) , .A2( u1_u3_u4_n120 ) , .ZN( u1_u3_u4_n130 ) );
  NAND2_X1 u1_u3_u4_U23 (.ZN( u1_u3_u4_n117 ) , .A2( u1_u3_u4_n118 ) , .A1( u1_u3_u4_n148 ) );
  NAND2_X1 u1_u3_u4_U24 (.ZN( u1_u3_u4_n129 ) , .A1( u1_u3_u4_n134 ) , .A2( u1_u3_u4_n148 ) );
  AND3_X1 u1_u3_u4_U25 (.A1( u1_u3_u4_n119 ) , .A2( u1_u3_u4_n143 ) , .A3( u1_u3_u4_n154 ) , .ZN( u1_u3_u4_n161 ) );
  AND2_X1 u1_u3_u4_U26 (.A1( u1_u3_u4_n145 ) , .A2( u1_u3_u4_n147 ) , .ZN( u1_u3_u4_n159 ) );
  OR3_X1 u1_u3_u4_U27 (.A3( u1_u3_u4_n114 ) , .A2( u1_u3_u4_n115 ) , .A1( u1_u3_u4_n116 ) , .ZN( u1_u3_u4_n136 ) );
  AOI21_X1 u1_u3_u4_U28 (.A( u1_u3_u4_n113 ) , .ZN( u1_u3_u4_n116 ) , .B2( u1_u3_u4_n173 ) , .B1( u1_u3_u4_n174 ) );
  AOI21_X1 u1_u3_u4_U29 (.ZN( u1_u3_u4_n115 ) , .B2( u1_u3_u4_n145 ) , .B1( u1_u3_u4_n146 ) , .A( u1_u3_u4_n156 ) );
  NOR2_X1 u1_u3_u4_U3 (.ZN( u1_u3_u4_n121 ) , .A1( u1_u3_u4_n181 ) , .A2( u1_u3_u4_n182 ) );
  OAI22_X1 u1_u3_u4_U30 (.ZN( u1_u3_u4_n114 ) , .A2( u1_u3_u4_n121 ) , .B1( u1_u3_u4_n160 ) , .B2( u1_u3_u4_n170 ) , .A1( u1_u3_u4_n171 ) );
  INV_X1 u1_u3_u4_U31 (.A( u1_u3_u4_n158 ) , .ZN( u1_u3_u4_n182 ) );
  INV_X1 u1_u3_u4_U32 (.ZN( u1_u3_u4_n181 ) , .A( u1_u3_u4_n96 ) );
  INV_X1 u1_u3_u4_U33 (.A( u1_u3_u4_n144 ) , .ZN( u1_u3_u4_n179 ) );
  INV_X1 u1_u3_u4_U34 (.A( u1_u3_u4_n157 ) , .ZN( u1_u3_u4_n178 ) );
  NAND2_X1 u1_u3_u4_U35 (.A2( u1_u3_u4_n154 ) , .A1( u1_u3_u4_n96 ) , .ZN( u1_u3_u4_n97 ) );
  INV_X1 u1_u3_u4_U36 (.ZN( u1_u3_u4_n186 ) , .A( u1_u3_u4_n95 ) );
  OAI221_X1 u1_u3_u4_U37 (.C1( u1_u3_u4_n134 ) , .B1( u1_u3_u4_n158 ) , .B2( u1_u3_u4_n171 ) , .C2( u1_u3_u4_n173 ) , .A( u1_u3_u4_n94 ) , .ZN( u1_u3_u4_n95 ) );
  AOI222_X1 u1_u3_u4_U38 (.B2( u1_u3_u4_n132 ) , .A1( u1_u3_u4_n138 ) , .C2( u1_u3_u4_n175 ) , .A2( u1_u3_u4_n179 ) , .C1( u1_u3_u4_n181 ) , .B1( u1_u3_u4_n185 ) , .ZN( u1_u3_u4_n94 ) );
  INV_X1 u1_u3_u4_U39 (.A( u1_u3_u4_n113 ) , .ZN( u1_u3_u4_n185 ) );
  INV_X1 u1_u3_u4_U4 (.A( u1_u3_u4_n117 ) , .ZN( u1_u3_u4_n184 ) );
  INV_X1 u1_u3_u4_U40 (.A( u1_u3_u4_n143 ) , .ZN( u1_u3_u4_n183 ) );
  NOR2_X1 u1_u3_u4_U41 (.ZN( u1_u3_u4_n138 ) , .A1( u1_u3_u4_n168 ) , .A2( u1_u3_u4_n169 ) );
  NOR2_X1 u1_u3_u4_U42 (.A1( u1_u3_u4_n150 ) , .A2( u1_u3_u4_n152 ) , .ZN( u1_u3_u4_n153 ) );
  NOR2_X1 u1_u3_u4_U43 (.A2( u1_u3_u4_n128 ) , .A1( u1_u3_u4_n138 ) , .ZN( u1_u3_u4_n156 ) );
  AOI22_X1 u1_u3_u4_U44 (.B2( u1_u3_u4_n122 ) , .A1( u1_u3_u4_n123 ) , .ZN( u1_u3_u4_n124 ) , .B1( u1_u3_u4_n128 ) , .A2( u1_u3_u4_n172 ) );
  INV_X1 u1_u3_u4_U45 (.A( u1_u3_u4_n153 ) , .ZN( u1_u3_u4_n172 ) );
  NAND2_X1 u1_u3_u4_U46 (.A2( u1_u3_u4_n120 ) , .ZN( u1_u3_u4_n123 ) , .A1( u1_u3_u4_n161 ) );
  AOI22_X1 u1_u3_u4_U47 (.B2( u1_u3_u4_n132 ) , .A2( u1_u3_u4_n133 ) , .ZN( u1_u3_u4_n140 ) , .A1( u1_u3_u4_n150 ) , .B1( u1_u3_u4_n179 ) );
  NAND2_X1 u1_u3_u4_U48 (.ZN( u1_u3_u4_n133 ) , .A2( u1_u3_u4_n146 ) , .A1( u1_u3_u4_n154 ) );
  NAND2_X1 u1_u3_u4_U49 (.A1( u1_u3_u4_n103 ) , .ZN( u1_u3_u4_n154 ) , .A2( u1_u3_u4_n98 ) );
  NOR4_X1 u1_u3_u4_U5 (.A4( u1_u3_u4_n106 ) , .A3( u1_u3_u4_n107 ) , .A2( u1_u3_u4_n108 ) , .A1( u1_u3_u4_n109 ) , .ZN( u1_u3_u4_n110 ) );
  NAND2_X1 u1_u3_u4_U50 (.A1( u1_u3_u4_n101 ) , .ZN( u1_u3_u4_n158 ) , .A2( u1_u3_u4_n99 ) );
  AOI21_X1 u1_u3_u4_U51 (.ZN( u1_u3_u4_n127 ) , .A( u1_u3_u4_n136 ) , .B2( u1_u3_u4_n150 ) , .B1( u1_u3_u4_n180 ) );
  INV_X1 u1_u3_u4_U52 (.A( u1_u3_u4_n160 ) , .ZN( u1_u3_u4_n180 ) );
  NAND2_X1 u1_u3_u4_U53 (.A2( u1_u3_u4_n104 ) , .A1( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n146 ) );
  NAND2_X1 u1_u3_u4_U54 (.A2( u1_u3_u4_n101 ) , .A1( u1_u3_u4_n102 ) , .ZN( u1_u3_u4_n160 ) );
  NAND2_X1 u1_u3_u4_U55 (.ZN( u1_u3_u4_n134 ) , .A1( u1_u3_u4_n98 ) , .A2( u1_u3_u4_n99 ) );
  NAND2_X1 u1_u3_u4_U56 (.A1( u1_u3_u4_n103 ) , .A2( u1_u3_u4_n104 ) , .ZN( u1_u3_u4_n143 ) );
  NAND2_X1 u1_u3_u4_U57 (.A2( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n145 ) , .A1( u1_u3_u4_n98 ) );
  NAND2_X1 u1_u3_u4_U58 (.A1( u1_u3_u4_n100 ) , .A2( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n120 ) );
  NAND2_X1 u1_u3_u4_U59 (.A1( u1_u3_u4_n102 ) , .A2( u1_u3_u4_n104 ) , .ZN( u1_u3_u4_n148 ) );
  AOI21_X1 u1_u3_u4_U6 (.ZN( u1_u3_u4_n106 ) , .B2( u1_u3_u4_n146 ) , .B1( u1_u3_u4_n158 ) , .A( u1_u3_u4_n170 ) );
  NAND2_X1 u1_u3_u4_U60 (.A2( u1_u3_u4_n100 ) , .A1( u1_u3_u4_n103 ) , .ZN( u1_u3_u4_n157 ) );
  INV_X1 u1_u3_u4_U61 (.A( u1_u3_u4_n150 ) , .ZN( u1_u3_u4_n173 ) );
  INV_X1 u1_u3_u4_U62 (.A( u1_u3_u4_n152 ) , .ZN( u1_u3_u4_n171 ) );
  NAND2_X1 u1_u3_u4_U63 (.A1( u1_u3_u4_n100 ) , .ZN( u1_u3_u4_n118 ) , .A2( u1_u3_u4_n99 ) );
  NAND2_X1 u1_u3_u4_U64 (.A2( u1_u3_u4_n100 ) , .A1( u1_u3_u4_n102 ) , .ZN( u1_u3_u4_n144 ) );
  NAND2_X1 u1_u3_u4_U65 (.A2( u1_u3_u4_n101 ) , .A1( u1_u3_u4_n105 ) , .ZN( u1_u3_u4_n96 ) );
  INV_X1 u1_u3_u4_U66 (.A( u1_u3_u4_n128 ) , .ZN( u1_u3_u4_n174 ) );
  NAND2_X1 u1_u3_u4_U67 (.A2( u1_u3_u4_n102 ) , .ZN( u1_u3_u4_n119 ) , .A1( u1_u3_u4_n98 ) );
  NAND2_X1 u1_u3_u4_U68 (.A2( u1_u3_u4_n101 ) , .A1( u1_u3_u4_n103 ) , .ZN( u1_u3_u4_n147 ) );
  NAND2_X1 u1_u3_u4_U69 (.A2( u1_u3_u4_n104 ) , .ZN( u1_u3_u4_n113 ) , .A1( u1_u3_u4_n99 ) );
  AOI21_X1 u1_u3_u4_U7 (.ZN( u1_u3_u4_n109 ) , .A( u1_u3_u4_n153 ) , .B1( u1_u3_u4_n159 ) , .B2( u1_u3_u4_n184 ) );
  NOR2_X1 u1_u3_u4_U70 (.A2( u1_u3_X_28 ) , .ZN( u1_u3_u4_n150 ) , .A1( u1_u3_u4_n168 ) );
  NOR2_X1 u1_u3_u4_U71 (.A2( u1_u3_X_29 ) , .ZN( u1_u3_u4_n152 ) , .A1( u1_u3_u4_n169 ) );
  NOR2_X1 u1_u3_u4_U72 (.A2( u1_u3_X_30 ) , .ZN( u1_u3_u4_n105 ) , .A1( u1_u3_u4_n176 ) );
  NOR2_X1 u1_u3_u4_U73 (.A2( u1_u3_X_26 ) , .ZN( u1_u3_u4_n100 ) , .A1( u1_u3_u4_n177 ) );
  NOR2_X1 u1_u3_u4_U74 (.A2( u1_u3_X_28 ) , .A1( u1_u3_X_29 ) , .ZN( u1_u3_u4_n128 ) );
  NOR2_X1 u1_u3_u4_U75 (.A2( u1_u3_X_27 ) , .A1( u1_u3_X_30 ) , .ZN( u1_u3_u4_n102 ) );
  NOR2_X1 u1_u3_u4_U76 (.A2( u1_u3_X_25 ) , .A1( u1_u3_X_26 ) , .ZN( u1_u3_u4_n98 ) );
  AND2_X1 u1_u3_u4_U77 (.A2( u1_u3_X_25 ) , .A1( u1_u3_X_26 ) , .ZN( u1_u3_u4_n104 ) );
  AND2_X1 u1_u3_u4_U78 (.A1( u1_u3_X_30 ) , .A2( u1_u3_u4_n176 ) , .ZN( u1_u3_u4_n99 ) );
  AND2_X1 u1_u3_u4_U79 (.A1( u1_u3_X_26 ) , .ZN( u1_u3_u4_n101 ) , .A2( u1_u3_u4_n177 ) );
  AOI21_X1 u1_u3_u4_U8 (.ZN( u1_u3_u4_n108 ) , .B2( u1_u3_u4_n134 ) , .B1( u1_u3_u4_n155 ) , .A( u1_u3_u4_n156 ) );
  AND2_X1 u1_u3_u4_U80 (.A1( u1_u3_X_27 ) , .A2( u1_u3_X_30 ) , .ZN( u1_u3_u4_n103 ) );
  INV_X1 u1_u3_u4_U81 (.A( u1_u3_X_28 ) , .ZN( u1_u3_u4_n169 ) );
  INV_X1 u1_u3_u4_U82 (.A( u1_u3_X_29 ) , .ZN( u1_u3_u4_n168 ) );
  INV_X1 u1_u3_u4_U83 (.A( u1_u3_X_25 ) , .ZN( u1_u3_u4_n177 ) );
  INV_X1 u1_u3_u4_U84 (.A( u1_u3_X_27 ) , .ZN( u1_u3_u4_n176 ) );
  NAND4_X1 u1_u3_u4_U85 (.ZN( u1_out3_25 ) , .A4( u1_u3_u4_n139 ) , .A3( u1_u3_u4_n140 ) , .A2( u1_u3_u4_n141 ) , .A1( u1_u3_u4_n142 ) );
  OAI21_X1 u1_u3_u4_U86 (.A( u1_u3_u4_n128 ) , .B2( u1_u3_u4_n129 ) , .B1( u1_u3_u4_n130 ) , .ZN( u1_u3_u4_n142 ) );
  OAI21_X1 u1_u3_u4_U87 (.B2( u1_u3_u4_n131 ) , .ZN( u1_u3_u4_n141 ) , .A( u1_u3_u4_n175 ) , .B1( u1_u3_u4_n183 ) );
  NAND4_X1 u1_u3_u4_U88 (.ZN( u1_out3_14 ) , .A4( u1_u3_u4_n124 ) , .A3( u1_u3_u4_n125 ) , .A2( u1_u3_u4_n126 ) , .A1( u1_u3_u4_n127 ) );
  AOI22_X1 u1_u3_u4_U89 (.B2( u1_u3_u4_n117 ) , .ZN( u1_u3_u4_n126 ) , .A1( u1_u3_u4_n129 ) , .B1( u1_u3_u4_n152 ) , .A2( u1_u3_u4_n175 ) );
  AOI211_X1 u1_u3_u4_U9 (.B( u1_u3_u4_n136 ) , .A( u1_u3_u4_n137 ) , .C2( u1_u3_u4_n138 ) , .ZN( u1_u3_u4_n139 ) , .C1( u1_u3_u4_n182 ) );
  AOI22_X1 u1_u3_u4_U90 (.ZN( u1_u3_u4_n125 ) , .B2( u1_u3_u4_n131 ) , .A2( u1_u3_u4_n132 ) , .B1( u1_u3_u4_n138 ) , .A1( u1_u3_u4_n178 ) );
  NAND4_X1 u1_u3_u4_U91 (.ZN( u1_out3_8 ) , .A4( u1_u3_u4_n110 ) , .A3( u1_u3_u4_n111 ) , .A2( u1_u3_u4_n112 ) , .A1( u1_u3_u4_n186 ) );
  NAND2_X1 u1_u3_u4_U92 (.ZN( u1_u3_u4_n112 ) , .A2( u1_u3_u4_n130 ) , .A1( u1_u3_u4_n150 ) );
  AOI22_X1 u1_u3_u4_U93 (.ZN( u1_u3_u4_n111 ) , .B2( u1_u3_u4_n132 ) , .A1( u1_u3_u4_n152 ) , .B1( u1_u3_u4_n178 ) , .A2( u1_u3_u4_n97 ) );
  AOI22_X1 u1_u3_u4_U94 (.B2( u1_u3_u4_n149 ) , .B1( u1_u3_u4_n150 ) , .A2( u1_u3_u4_n151 ) , .A1( u1_u3_u4_n152 ) , .ZN( u1_u3_u4_n167 ) );
  NOR4_X1 u1_u3_u4_U95 (.A4( u1_u3_u4_n162 ) , .A3( u1_u3_u4_n163 ) , .A2( u1_u3_u4_n164 ) , .A1( u1_u3_u4_n165 ) , .ZN( u1_u3_u4_n166 ) );
  NAND3_X1 u1_u3_u4_U96 (.ZN( u1_out3_3 ) , .A3( u1_u3_u4_n166 ) , .A1( u1_u3_u4_n167 ) , .A2( u1_u3_u4_n186 ) );
  NAND3_X1 u1_u3_u4_U97 (.A3( u1_u3_u4_n146 ) , .A2( u1_u3_u4_n147 ) , .A1( u1_u3_u4_n148 ) , .ZN( u1_u3_u4_n149 ) );
  NAND3_X1 u1_u3_u4_U98 (.A3( u1_u3_u4_n143 ) , .A2( u1_u3_u4_n144 ) , .A1( u1_u3_u4_n145 ) , .ZN( u1_u3_u4_n151 ) );
  NAND3_X1 u1_u3_u4_U99 (.A3( u1_u3_u4_n121 ) , .ZN( u1_u3_u4_n122 ) , .A2( u1_u3_u4_n144 ) , .A1( u1_u3_u4_n154 ) );
  INV_X1 u1_u3_u5_U10 (.A( u1_u3_u5_n121 ) , .ZN( u1_u3_u5_n177 ) );
  NOR3_X1 u1_u3_u5_U100 (.A3( u1_u3_u5_n141 ) , .A1( u1_u3_u5_n142 ) , .ZN( u1_u3_u5_n143 ) , .A2( u1_u3_u5_n191 ) );
  NAND4_X1 u1_u3_u5_U101 (.ZN( u1_out3_4 ) , .A4( u1_u3_u5_n112 ) , .A2( u1_u3_u5_n113 ) , .A1( u1_u3_u5_n114 ) , .A3( u1_u3_u5_n195 ) );
  AOI211_X1 u1_u3_u5_U102 (.A( u1_u3_u5_n110 ) , .C1( u1_u3_u5_n111 ) , .ZN( u1_u3_u5_n112 ) , .B( u1_u3_u5_n118 ) , .C2( u1_u3_u5_n177 ) );
  AOI222_X1 u1_u3_u5_U103 (.ZN( u1_u3_u5_n113 ) , .A1( u1_u3_u5_n131 ) , .C1( u1_u3_u5_n148 ) , .B2( u1_u3_u5_n174 ) , .C2( u1_u3_u5_n178 ) , .A2( u1_u3_u5_n179 ) , .B1( u1_u3_u5_n99 ) );
  NAND3_X1 u1_u3_u5_U104 (.A2( u1_u3_u5_n154 ) , .A3( u1_u3_u5_n158 ) , .A1( u1_u3_u5_n161 ) , .ZN( u1_u3_u5_n99 ) );
  NOR2_X1 u1_u3_u5_U11 (.ZN( u1_u3_u5_n160 ) , .A2( u1_u3_u5_n173 ) , .A1( u1_u3_u5_n177 ) );
  INV_X1 u1_u3_u5_U12 (.A( u1_u3_u5_n150 ) , .ZN( u1_u3_u5_n174 ) );
  AOI21_X1 u1_u3_u5_U13 (.A( u1_u3_u5_n160 ) , .B2( u1_u3_u5_n161 ) , .ZN( u1_u3_u5_n162 ) , .B1( u1_u3_u5_n192 ) );
  INV_X1 u1_u3_u5_U14 (.A( u1_u3_u5_n159 ) , .ZN( u1_u3_u5_n192 ) );
  AOI21_X1 u1_u3_u5_U15 (.A( u1_u3_u5_n156 ) , .B2( u1_u3_u5_n157 ) , .B1( u1_u3_u5_n158 ) , .ZN( u1_u3_u5_n163 ) );
  AOI21_X1 u1_u3_u5_U16 (.B2( u1_u3_u5_n139 ) , .B1( u1_u3_u5_n140 ) , .ZN( u1_u3_u5_n141 ) , .A( u1_u3_u5_n150 ) );
  OAI21_X1 u1_u3_u5_U17 (.A( u1_u3_u5_n133 ) , .B2( u1_u3_u5_n134 ) , .B1( u1_u3_u5_n135 ) , .ZN( u1_u3_u5_n142 ) );
  OAI21_X1 u1_u3_u5_U18 (.ZN( u1_u3_u5_n133 ) , .B2( u1_u3_u5_n147 ) , .A( u1_u3_u5_n173 ) , .B1( u1_u3_u5_n188 ) );
  NAND2_X1 u1_u3_u5_U19 (.A2( u1_u3_u5_n119 ) , .A1( u1_u3_u5_n123 ) , .ZN( u1_u3_u5_n137 ) );
  INV_X1 u1_u3_u5_U20 (.A( u1_u3_u5_n155 ) , .ZN( u1_u3_u5_n194 ) );
  NAND2_X1 u1_u3_u5_U21 (.A1( u1_u3_u5_n121 ) , .ZN( u1_u3_u5_n132 ) , .A2( u1_u3_u5_n172 ) );
  NAND2_X1 u1_u3_u5_U22 (.A2( u1_u3_u5_n122 ) , .ZN( u1_u3_u5_n136 ) , .A1( u1_u3_u5_n154 ) );
  NAND2_X1 u1_u3_u5_U23 (.A2( u1_u3_u5_n119 ) , .A1( u1_u3_u5_n120 ) , .ZN( u1_u3_u5_n159 ) );
  INV_X1 u1_u3_u5_U24 (.A( u1_u3_u5_n156 ) , .ZN( u1_u3_u5_n175 ) );
  INV_X1 u1_u3_u5_U25 (.A( u1_u3_u5_n158 ) , .ZN( u1_u3_u5_n188 ) );
  INV_X1 u1_u3_u5_U26 (.A( u1_u3_u5_n152 ) , .ZN( u1_u3_u5_n179 ) );
  INV_X1 u1_u3_u5_U27 (.A( u1_u3_u5_n140 ) , .ZN( u1_u3_u5_n182 ) );
  INV_X1 u1_u3_u5_U28 (.A( u1_u3_u5_n151 ) , .ZN( u1_u3_u5_n183 ) );
  INV_X1 u1_u3_u5_U29 (.A( u1_u3_u5_n123 ) , .ZN( u1_u3_u5_n185 ) );
  NOR2_X1 u1_u3_u5_U3 (.ZN( u1_u3_u5_n134 ) , .A1( u1_u3_u5_n183 ) , .A2( u1_u3_u5_n190 ) );
  INV_X1 u1_u3_u5_U30 (.A( u1_u3_u5_n161 ) , .ZN( u1_u3_u5_n184 ) );
  INV_X1 u1_u3_u5_U31 (.A( u1_u3_u5_n139 ) , .ZN( u1_u3_u5_n189 ) );
  INV_X1 u1_u3_u5_U32 (.A( u1_u3_u5_n157 ) , .ZN( u1_u3_u5_n190 ) );
  INV_X1 u1_u3_u5_U33 (.A( u1_u3_u5_n120 ) , .ZN( u1_u3_u5_n193 ) );
  NAND2_X1 u1_u3_u5_U34 (.ZN( u1_u3_u5_n111 ) , .A1( u1_u3_u5_n140 ) , .A2( u1_u3_u5_n155 ) );
  INV_X1 u1_u3_u5_U35 (.A( u1_u3_u5_n117 ) , .ZN( u1_u3_u5_n196 ) );
  OAI221_X1 u1_u3_u5_U36 (.A( u1_u3_u5_n116 ) , .ZN( u1_u3_u5_n117 ) , .B2( u1_u3_u5_n119 ) , .C1( u1_u3_u5_n153 ) , .C2( u1_u3_u5_n158 ) , .B1( u1_u3_u5_n172 ) );
  AOI222_X1 u1_u3_u5_U37 (.ZN( u1_u3_u5_n116 ) , .B2( u1_u3_u5_n145 ) , .C1( u1_u3_u5_n148 ) , .A2( u1_u3_u5_n174 ) , .C2( u1_u3_u5_n177 ) , .B1( u1_u3_u5_n187 ) , .A1( u1_u3_u5_n193 ) );
  INV_X1 u1_u3_u5_U38 (.A( u1_u3_u5_n115 ) , .ZN( u1_u3_u5_n187 ) );
  NOR2_X1 u1_u3_u5_U39 (.ZN( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n170 ) , .A2( u1_u3_u5_n180 ) );
  INV_X1 u1_u3_u5_U4 (.A( u1_u3_u5_n138 ) , .ZN( u1_u3_u5_n191 ) );
  AOI22_X1 u1_u3_u5_U40 (.B2( u1_u3_u5_n131 ) , .A2( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n169 ) , .B1( u1_u3_u5_n174 ) , .A1( u1_u3_u5_n185 ) );
  NOR2_X1 u1_u3_u5_U41 (.A1( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n150 ) , .A2( u1_u3_u5_n173 ) );
  AOI21_X1 u1_u3_u5_U42 (.A( u1_u3_u5_n118 ) , .B2( u1_u3_u5_n145 ) , .ZN( u1_u3_u5_n168 ) , .B1( u1_u3_u5_n186 ) );
  INV_X1 u1_u3_u5_U43 (.A( u1_u3_u5_n122 ) , .ZN( u1_u3_u5_n186 ) );
  NOR2_X1 u1_u3_u5_U44 (.A1( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n152 ) , .A2( u1_u3_u5_n176 ) );
  NOR2_X1 u1_u3_u5_U45 (.A1( u1_u3_u5_n115 ) , .ZN( u1_u3_u5_n118 ) , .A2( u1_u3_u5_n153 ) );
  NOR2_X1 u1_u3_u5_U46 (.A2( u1_u3_u5_n145 ) , .ZN( u1_u3_u5_n156 ) , .A1( u1_u3_u5_n174 ) );
  NOR2_X1 u1_u3_u5_U47 (.ZN( u1_u3_u5_n121 ) , .A2( u1_u3_u5_n145 ) , .A1( u1_u3_u5_n176 ) );
  AOI22_X1 u1_u3_u5_U48 (.ZN( u1_u3_u5_n114 ) , .A2( u1_u3_u5_n137 ) , .A1( u1_u3_u5_n145 ) , .B2( u1_u3_u5_n175 ) , .B1( u1_u3_u5_n193 ) );
  OAI211_X1 u1_u3_u5_U49 (.B( u1_u3_u5_n124 ) , .A( u1_u3_u5_n125 ) , .C2( u1_u3_u5_n126 ) , .C1( u1_u3_u5_n127 ) , .ZN( u1_u3_u5_n128 ) );
  OAI21_X1 u1_u3_u5_U5 (.B2( u1_u3_u5_n136 ) , .B1( u1_u3_u5_n137 ) , .ZN( u1_u3_u5_n138 ) , .A( u1_u3_u5_n177 ) );
  NOR3_X1 u1_u3_u5_U50 (.ZN( u1_u3_u5_n127 ) , .A1( u1_u3_u5_n136 ) , .A3( u1_u3_u5_n148 ) , .A2( u1_u3_u5_n182 ) );
  OAI21_X1 u1_u3_u5_U51 (.ZN( u1_u3_u5_n124 ) , .A( u1_u3_u5_n177 ) , .B2( u1_u3_u5_n183 ) , .B1( u1_u3_u5_n189 ) );
  OAI21_X1 u1_u3_u5_U52 (.ZN( u1_u3_u5_n125 ) , .A( u1_u3_u5_n174 ) , .B2( u1_u3_u5_n185 ) , .B1( u1_u3_u5_n190 ) );
  AOI21_X1 u1_u3_u5_U53 (.A( u1_u3_u5_n153 ) , .B2( u1_u3_u5_n154 ) , .B1( u1_u3_u5_n155 ) , .ZN( u1_u3_u5_n164 ) );
  AOI21_X1 u1_u3_u5_U54 (.ZN( u1_u3_u5_n110 ) , .B1( u1_u3_u5_n122 ) , .B2( u1_u3_u5_n139 ) , .A( u1_u3_u5_n153 ) );
  INV_X1 u1_u3_u5_U55 (.A( u1_u3_u5_n153 ) , .ZN( u1_u3_u5_n176 ) );
  INV_X1 u1_u3_u5_U56 (.A( u1_u3_u5_n126 ) , .ZN( u1_u3_u5_n173 ) );
  AND2_X1 u1_u3_u5_U57 (.A2( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n107 ) , .ZN( u1_u3_u5_n147 ) );
  AND2_X1 u1_u3_u5_U58 (.A2( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n108 ) , .ZN( u1_u3_u5_n148 ) );
  NAND2_X1 u1_u3_u5_U59 (.A1( u1_u3_u5_n105 ) , .A2( u1_u3_u5_n106 ) , .ZN( u1_u3_u5_n158 ) );
  INV_X1 u1_u3_u5_U6 (.A( u1_u3_u5_n135 ) , .ZN( u1_u3_u5_n178 ) );
  NAND2_X1 u1_u3_u5_U60 (.A2( u1_u3_u5_n108 ) , .A1( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n139 ) );
  NAND2_X1 u1_u3_u5_U61 (.A1( u1_u3_u5_n106 ) , .A2( u1_u3_u5_n108 ) , .ZN( u1_u3_u5_n119 ) );
  NAND2_X1 u1_u3_u5_U62 (.A2( u1_u3_u5_n103 ) , .A1( u1_u3_u5_n105 ) , .ZN( u1_u3_u5_n140 ) );
  NAND2_X1 u1_u3_u5_U63 (.A2( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n105 ) , .ZN( u1_u3_u5_n155 ) );
  NAND2_X1 u1_u3_u5_U64 (.A2( u1_u3_u5_n106 ) , .A1( u1_u3_u5_n107 ) , .ZN( u1_u3_u5_n122 ) );
  NAND2_X1 u1_u3_u5_U65 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n106 ) , .ZN( u1_u3_u5_n115 ) );
  NAND2_X1 u1_u3_u5_U66 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n103 ) , .ZN( u1_u3_u5_n161 ) );
  NAND2_X1 u1_u3_u5_U67 (.A1( u1_u3_u5_n105 ) , .A2( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n154 ) );
  INV_X1 u1_u3_u5_U68 (.A( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n172 ) );
  NAND2_X1 u1_u3_u5_U69 (.A1( u1_u3_u5_n103 ) , .A2( u1_u3_u5_n108 ) , .ZN( u1_u3_u5_n123 ) );
  OAI22_X1 u1_u3_u5_U7 (.B2( u1_u3_u5_n149 ) , .B1( u1_u3_u5_n150 ) , .A2( u1_u3_u5_n151 ) , .A1( u1_u3_u5_n152 ) , .ZN( u1_u3_u5_n165 ) );
  NAND2_X1 u1_u3_u5_U70 (.A2( u1_u3_u5_n103 ) , .A1( u1_u3_u5_n107 ) , .ZN( u1_u3_u5_n151 ) );
  NAND2_X1 u1_u3_u5_U71 (.A2( u1_u3_u5_n107 ) , .A1( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n120 ) );
  NAND2_X1 u1_u3_u5_U72 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n109 ) , .ZN( u1_u3_u5_n157 ) );
  AND2_X1 u1_u3_u5_U73 (.A2( u1_u3_u5_n100 ) , .A1( u1_u3_u5_n104 ) , .ZN( u1_u3_u5_n131 ) );
  INV_X1 u1_u3_u5_U74 (.A( u1_u3_u5_n102 ) , .ZN( u1_u3_u5_n195 ) );
  OAI221_X1 u1_u3_u5_U75 (.A( u1_u3_u5_n101 ) , .ZN( u1_u3_u5_n102 ) , .C2( u1_u3_u5_n115 ) , .C1( u1_u3_u5_n126 ) , .B1( u1_u3_u5_n134 ) , .B2( u1_u3_u5_n160 ) );
  OAI21_X1 u1_u3_u5_U76 (.ZN( u1_u3_u5_n101 ) , .B1( u1_u3_u5_n137 ) , .A( u1_u3_u5_n146 ) , .B2( u1_u3_u5_n147 ) );
  NOR2_X1 u1_u3_u5_U77 (.A2( u1_u3_X_34 ) , .A1( u1_u3_X_35 ) , .ZN( u1_u3_u5_n145 ) );
  NOR2_X1 u1_u3_u5_U78 (.A2( u1_u3_X_34 ) , .ZN( u1_u3_u5_n146 ) , .A1( u1_u3_u5_n171 ) );
  NOR2_X1 u1_u3_u5_U79 (.A2( u1_u3_X_31 ) , .A1( u1_u3_X_32 ) , .ZN( u1_u3_u5_n103 ) );
  NOR3_X1 u1_u3_u5_U8 (.A2( u1_u3_u5_n147 ) , .A1( u1_u3_u5_n148 ) , .ZN( u1_u3_u5_n149 ) , .A3( u1_u3_u5_n194 ) );
  NOR2_X1 u1_u3_u5_U80 (.A2( u1_u3_X_36 ) , .ZN( u1_u3_u5_n105 ) , .A1( u1_u3_u5_n180 ) );
  NOR2_X1 u1_u3_u5_U81 (.A2( u1_u3_X_33 ) , .ZN( u1_u3_u5_n108 ) , .A1( u1_u3_u5_n170 ) );
  NOR2_X1 u1_u3_u5_U82 (.A2( u1_u3_X_33 ) , .A1( u1_u3_X_36 ) , .ZN( u1_u3_u5_n107 ) );
  NOR2_X1 u1_u3_u5_U83 (.A2( u1_u3_X_31 ) , .ZN( u1_u3_u5_n104 ) , .A1( u1_u3_u5_n181 ) );
  NAND2_X1 u1_u3_u5_U84 (.A2( u1_u3_X_34 ) , .A1( u1_u3_X_35 ) , .ZN( u1_u3_u5_n153 ) );
  NAND2_X1 u1_u3_u5_U85 (.A1( u1_u3_X_34 ) , .ZN( u1_u3_u5_n126 ) , .A2( u1_u3_u5_n171 ) );
  AND2_X1 u1_u3_u5_U86 (.A1( u1_u3_X_31 ) , .A2( u1_u3_X_32 ) , .ZN( u1_u3_u5_n106 ) );
  AND2_X1 u1_u3_u5_U87 (.A1( u1_u3_X_31 ) , .ZN( u1_u3_u5_n109 ) , .A2( u1_u3_u5_n181 ) );
  INV_X1 u1_u3_u5_U88 (.A( u1_u3_X_33 ) , .ZN( u1_u3_u5_n180 ) );
  INV_X1 u1_u3_u5_U89 (.A( u1_u3_X_35 ) , .ZN( u1_u3_u5_n171 ) );
  NOR2_X1 u1_u3_u5_U9 (.ZN( u1_u3_u5_n135 ) , .A1( u1_u3_u5_n173 ) , .A2( u1_u3_u5_n176 ) );
  INV_X1 u1_u3_u5_U90 (.A( u1_u3_X_36 ) , .ZN( u1_u3_u5_n170 ) );
  INV_X1 u1_u3_u5_U91 (.A( u1_u3_X_32 ) , .ZN( u1_u3_u5_n181 ) );
  NAND4_X1 u1_u3_u5_U92 (.ZN( u1_out3_29 ) , .A4( u1_u3_u5_n129 ) , .A3( u1_u3_u5_n130 ) , .A2( u1_u3_u5_n168 ) , .A1( u1_u3_u5_n196 ) );
  AOI221_X1 u1_u3_u5_U93 (.A( u1_u3_u5_n128 ) , .ZN( u1_u3_u5_n129 ) , .C2( u1_u3_u5_n132 ) , .B2( u1_u3_u5_n159 ) , .B1( u1_u3_u5_n176 ) , .C1( u1_u3_u5_n184 ) );
  AOI222_X1 u1_u3_u5_U94 (.ZN( u1_u3_u5_n130 ) , .A2( u1_u3_u5_n146 ) , .B1( u1_u3_u5_n147 ) , .C2( u1_u3_u5_n175 ) , .B2( u1_u3_u5_n179 ) , .A1( u1_u3_u5_n188 ) , .C1( u1_u3_u5_n194 ) );
  NAND4_X1 u1_u3_u5_U95 (.ZN( u1_out3_19 ) , .A4( u1_u3_u5_n166 ) , .A3( u1_u3_u5_n167 ) , .A2( u1_u3_u5_n168 ) , .A1( u1_u3_u5_n169 ) );
  AOI22_X1 u1_u3_u5_U96 (.B2( u1_u3_u5_n145 ) , .A2( u1_u3_u5_n146 ) , .ZN( u1_u3_u5_n167 ) , .B1( u1_u3_u5_n182 ) , .A1( u1_u3_u5_n189 ) );
  NOR4_X1 u1_u3_u5_U97 (.A4( u1_u3_u5_n162 ) , .A3( u1_u3_u5_n163 ) , .A2( u1_u3_u5_n164 ) , .A1( u1_u3_u5_n165 ) , .ZN( u1_u3_u5_n166 ) );
  NAND4_X1 u1_u3_u5_U98 (.ZN( u1_out3_11 ) , .A4( u1_u3_u5_n143 ) , .A3( u1_u3_u5_n144 ) , .A2( u1_u3_u5_n169 ) , .A1( u1_u3_u5_n196 ) );
  AOI22_X1 u1_u3_u5_U99 (.A2( u1_u3_u5_n132 ) , .ZN( u1_u3_u5_n144 ) , .B2( u1_u3_u5_n145 ) , .B1( u1_u3_u5_n184 ) , .A1( u1_u3_u5_n194 ) );
  AND3_X1 u1_u3_u7_U10 (.A3( u1_u3_u7_n110 ) , .A2( u1_u3_u7_n127 ) , .A1( u1_u3_u7_n132 ) , .ZN( u1_u3_u7_n92 ) );
  OAI21_X1 u1_u3_u7_U11 (.A( u1_u3_u7_n161 ) , .B1( u1_u3_u7_n168 ) , .B2( u1_u3_u7_n173 ) , .ZN( u1_u3_u7_n91 ) );
  AOI211_X1 u1_u3_u7_U12 (.A( u1_u3_u7_n117 ) , .ZN( u1_u3_u7_n118 ) , .C2( u1_u3_u7_n126 ) , .C1( u1_u3_u7_n177 ) , .B( u1_u3_u7_n180 ) );
  OAI22_X1 u1_u3_u7_U13 (.B1( u1_u3_u7_n115 ) , .ZN( u1_u3_u7_n117 ) , .A2( u1_u3_u7_n133 ) , .A1( u1_u3_u7_n137 ) , .B2( u1_u3_u7_n162 ) );
  INV_X1 u1_u3_u7_U14 (.A( u1_u3_u7_n116 ) , .ZN( u1_u3_u7_n180 ) );
  NOR3_X1 u1_u3_u7_U15 (.ZN( u1_u3_u7_n115 ) , .A3( u1_u3_u7_n145 ) , .A2( u1_u3_u7_n168 ) , .A1( u1_u3_u7_n169 ) );
  OAI211_X1 u1_u3_u7_U16 (.B( u1_u3_u7_n122 ) , .A( u1_u3_u7_n123 ) , .C2( u1_u3_u7_n124 ) , .ZN( u1_u3_u7_n154 ) , .C1( u1_u3_u7_n162 ) );
  AOI222_X1 u1_u3_u7_U17 (.ZN( u1_u3_u7_n122 ) , .C2( u1_u3_u7_n126 ) , .C1( u1_u3_u7_n145 ) , .B1( u1_u3_u7_n161 ) , .A2( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n170 ) , .A1( u1_u3_u7_n176 ) );
  INV_X1 u1_u3_u7_U18 (.A( u1_u3_u7_n133 ) , .ZN( u1_u3_u7_n176 ) );
  NOR3_X1 u1_u3_u7_U19 (.A2( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n135 ) , .ZN( u1_u3_u7_n136 ) , .A3( u1_u3_u7_n171 ) );
  NOR2_X1 u1_u3_u7_U20 (.A1( u1_u3_u7_n130 ) , .A2( u1_u3_u7_n134 ) , .ZN( u1_u3_u7_n153 ) );
  INV_X1 u1_u3_u7_U21 (.A( u1_u3_u7_n101 ) , .ZN( u1_u3_u7_n165 ) );
  NOR2_X1 u1_u3_u7_U22 (.ZN( u1_u3_u7_n111 ) , .A2( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n169 ) );
  AOI21_X1 u1_u3_u7_U23 (.ZN( u1_u3_u7_n104 ) , .B2( u1_u3_u7_n112 ) , .B1( u1_u3_u7_n127 ) , .A( u1_u3_u7_n164 ) );
  AOI21_X1 u1_u3_u7_U24 (.ZN( u1_u3_u7_n106 ) , .B1( u1_u3_u7_n133 ) , .B2( u1_u3_u7_n146 ) , .A( u1_u3_u7_n162 ) );
  AOI21_X1 u1_u3_u7_U25 (.A( u1_u3_u7_n101 ) , .ZN( u1_u3_u7_n107 ) , .B2( u1_u3_u7_n128 ) , .B1( u1_u3_u7_n175 ) );
  INV_X1 u1_u3_u7_U26 (.A( u1_u3_u7_n138 ) , .ZN( u1_u3_u7_n171 ) );
  INV_X1 u1_u3_u7_U27 (.A( u1_u3_u7_n131 ) , .ZN( u1_u3_u7_n177 ) );
  INV_X1 u1_u3_u7_U28 (.A( u1_u3_u7_n110 ) , .ZN( u1_u3_u7_n174 ) );
  NAND2_X1 u1_u3_u7_U29 (.A1( u1_u3_u7_n129 ) , .A2( u1_u3_u7_n132 ) , .ZN( u1_u3_u7_n149 ) );
  OAI21_X1 u1_u3_u7_U3 (.ZN( u1_u3_u7_n159 ) , .A( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n171 ) , .B1( u1_u3_u7_n174 ) );
  NAND2_X1 u1_u3_u7_U30 (.A1( u1_u3_u7_n113 ) , .A2( u1_u3_u7_n124 ) , .ZN( u1_u3_u7_n130 ) );
  INV_X1 u1_u3_u7_U31 (.A( u1_u3_u7_n112 ) , .ZN( u1_u3_u7_n173 ) );
  INV_X1 u1_u3_u7_U32 (.A( u1_u3_u7_n128 ) , .ZN( u1_u3_u7_n168 ) );
  INV_X1 u1_u3_u7_U33 (.A( u1_u3_u7_n148 ) , .ZN( u1_u3_u7_n169 ) );
  INV_X1 u1_u3_u7_U34 (.A( u1_u3_u7_n127 ) , .ZN( u1_u3_u7_n179 ) );
  NOR2_X1 u1_u3_u7_U35 (.ZN( u1_u3_u7_n101 ) , .A2( u1_u3_u7_n150 ) , .A1( u1_u3_u7_n156 ) );
  AOI211_X1 u1_u3_u7_U36 (.B( u1_u3_u7_n154 ) , .A( u1_u3_u7_n155 ) , .C1( u1_u3_u7_n156 ) , .ZN( u1_u3_u7_n157 ) , .C2( u1_u3_u7_n172 ) );
  INV_X1 u1_u3_u7_U37 (.A( u1_u3_u7_n153 ) , .ZN( u1_u3_u7_n172 ) );
  AOI211_X1 u1_u3_u7_U38 (.B( u1_u3_u7_n139 ) , .A( u1_u3_u7_n140 ) , .C2( u1_u3_u7_n141 ) , .ZN( u1_u3_u7_n142 ) , .C1( u1_u3_u7_n156 ) );
  NAND4_X1 u1_u3_u7_U39 (.A3( u1_u3_u7_n127 ) , .A2( u1_u3_u7_n128 ) , .A1( u1_u3_u7_n129 ) , .ZN( u1_u3_u7_n141 ) , .A4( u1_u3_u7_n147 ) );
  INV_X1 u1_u3_u7_U4 (.A( u1_u3_u7_n111 ) , .ZN( u1_u3_u7_n170 ) );
  AOI21_X1 u1_u3_u7_U40 (.A( u1_u3_u7_n137 ) , .B1( u1_u3_u7_n138 ) , .ZN( u1_u3_u7_n139 ) , .B2( u1_u3_u7_n146 ) );
  OAI22_X1 u1_u3_u7_U41 (.B1( u1_u3_u7_n136 ) , .ZN( u1_u3_u7_n140 ) , .A1( u1_u3_u7_n153 ) , .B2( u1_u3_u7_n162 ) , .A2( u1_u3_u7_n164 ) );
  AOI21_X1 u1_u3_u7_U42 (.ZN( u1_u3_u7_n123 ) , .B1( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n177 ) , .A( u1_u3_u7_n97 ) );
  AOI21_X1 u1_u3_u7_U43 (.B2( u1_u3_u7_n113 ) , .B1( u1_u3_u7_n124 ) , .A( u1_u3_u7_n125 ) , .ZN( u1_u3_u7_n97 ) );
  INV_X1 u1_u3_u7_U44 (.A( u1_u3_u7_n125 ) , .ZN( u1_u3_u7_n161 ) );
  INV_X1 u1_u3_u7_U45 (.A( u1_u3_u7_n152 ) , .ZN( u1_u3_u7_n162 ) );
  AOI22_X1 u1_u3_u7_U46 (.A2( u1_u3_u7_n114 ) , .ZN( u1_u3_u7_n119 ) , .B1( u1_u3_u7_n130 ) , .A1( u1_u3_u7_n156 ) , .B2( u1_u3_u7_n165 ) );
  NAND2_X1 u1_u3_u7_U47 (.A2( u1_u3_u7_n112 ) , .ZN( u1_u3_u7_n114 ) , .A1( u1_u3_u7_n175 ) );
  AND2_X1 u1_u3_u7_U48 (.ZN( u1_u3_u7_n145 ) , .A2( u1_u3_u7_n98 ) , .A1( u1_u3_u7_n99 ) );
  NOR2_X1 u1_u3_u7_U49 (.ZN( u1_u3_u7_n137 ) , .A1( u1_u3_u7_n150 ) , .A2( u1_u3_u7_n161 ) );
  INV_X1 u1_u3_u7_U5 (.A( u1_u3_u7_n149 ) , .ZN( u1_u3_u7_n175 ) );
  AOI21_X1 u1_u3_u7_U50 (.ZN( u1_u3_u7_n105 ) , .B2( u1_u3_u7_n110 ) , .A( u1_u3_u7_n125 ) , .B1( u1_u3_u7_n147 ) );
  NAND2_X1 u1_u3_u7_U51 (.ZN( u1_u3_u7_n146 ) , .A1( u1_u3_u7_n95 ) , .A2( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U52 (.A2( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n147 ) , .A1( u1_u3_u7_n93 ) );
  NAND2_X1 u1_u3_u7_U53 (.A1( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n127 ) , .A2( u1_u3_u7_n99 ) );
  OR2_X1 u1_u3_u7_U54 (.ZN( u1_u3_u7_n126 ) , .A2( u1_u3_u7_n152 ) , .A1( u1_u3_u7_n156 ) );
  NAND2_X1 u1_u3_u7_U55 (.A2( u1_u3_u7_n102 ) , .A1( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n133 ) );
  NAND2_X1 u1_u3_u7_U56 (.ZN( u1_u3_u7_n112 ) , .A2( u1_u3_u7_n96 ) , .A1( u1_u3_u7_n99 ) );
  NAND2_X1 u1_u3_u7_U57 (.A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n128 ) , .A1( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U58 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n113 ) , .A2( u1_u3_u7_n93 ) );
  NAND2_X1 u1_u3_u7_U59 (.A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n124 ) , .A1( u1_u3_u7_n96 ) );
  INV_X1 u1_u3_u7_U6 (.A( u1_u3_u7_n154 ) , .ZN( u1_u3_u7_n178 ) );
  NAND2_X1 u1_u3_u7_U60 (.ZN( u1_u3_u7_n110 ) , .A1( u1_u3_u7_n95 ) , .A2( u1_u3_u7_n96 ) );
  INV_X1 u1_u3_u7_U61 (.A( u1_u3_u7_n150 ) , .ZN( u1_u3_u7_n164 ) );
  AND2_X1 u1_u3_u7_U62 (.ZN( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n93 ) , .A2( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U63 (.A1( u1_u3_u7_n100 ) , .A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n129 ) );
  NAND2_X1 u1_u3_u7_U64 (.A2( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n131 ) , .A1( u1_u3_u7_n95 ) );
  NAND2_X1 u1_u3_u7_U65 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n138 ) , .A2( u1_u3_u7_n99 ) );
  NAND2_X1 u1_u3_u7_U66 (.ZN( u1_u3_u7_n132 ) , .A1( u1_u3_u7_n93 ) , .A2( u1_u3_u7_n96 ) );
  NAND2_X1 u1_u3_u7_U67 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n148 ) , .A2( u1_u3_u7_n95 ) );
  NOR2_X1 u1_u3_u7_U68 (.A2( u1_u3_X_47 ) , .ZN( u1_u3_u7_n150 ) , .A1( u1_u3_u7_n163 ) );
  NOR2_X1 u1_u3_u7_U69 (.A2( u1_u3_X_43 ) , .A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n103 ) );
  AOI211_X1 u1_u3_u7_U7 (.ZN( u1_u3_u7_n116 ) , .A( u1_u3_u7_n155 ) , .C1( u1_u3_u7_n161 ) , .C2( u1_u3_u7_n171 ) , .B( u1_u3_u7_n94 ) );
  NOR2_X1 u1_u3_u7_U70 (.A2( u1_u3_X_48 ) , .A1( u1_u3_u7_n166 ) , .ZN( u1_u3_u7_n95 ) );
  NOR2_X1 u1_u3_u7_U71 (.A2( u1_u3_X_45 ) , .A1( u1_u3_X_48 ) , .ZN( u1_u3_u7_n99 ) );
  NOR2_X1 u1_u3_u7_U72 (.A2( u1_u3_X_44 ) , .A1( u1_u3_u7_n167 ) , .ZN( u1_u3_u7_n98 ) );
  NOR2_X1 u1_u3_u7_U73 (.A2( u1_u3_X_46 ) , .A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n152 ) );
  AND2_X1 u1_u3_u7_U74 (.A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n156 ) , .A2( u1_u3_u7_n163 ) );
  NAND2_X1 u1_u3_u7_U75 (.A2( u1_u3_X_46 ) , .A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n125 ) );
  AND2_X1 u1_u3_u7_U76 (.A2( u1_u3_X_45 ) , .A1( u1_u3_X_48 ) , .ZN( u1_u3_u7_n102 ) );
  AND2_X1 u1_u3_u7_U77 (.A2( u1_u3_X_43 ) , .A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n96 ) );
  AND2_X1 u1_u3_u7_U78 (.A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n100 ) , .A2( u1_u3_u7_n167 ) );
  AND2_X1 u1_u3_u7_U79 (.A1( u1_u3_X_48 ) , .A2( u1_u3_u7_n166 ) , .ZN( u1_u3_u7_n93 ) );
  OAI222_X1 u1_u3_u7_U8 (.C2( u1_u3_u7_n101 ) , .B2( u1_u3_u7_n111 ) , .A1( u1_u3_u7_n113 ) , .C1( u1_u3_u7_n146 ) , .A2( u1_u3_u7_n162 ) , .B1( u1_u3_u7_n164 ) , .ZN( u1_u3_u7_n94 ) );
  INV_X1 u1_u3_u7_U80 (.A( u1_u3_X_46 ) , .ZN( u1_u3_u7_n163 ) );
  INV_X1 u1_u3_u7_U81 (.A( u1_u3_X_43 ) , .ZN( u1_u3_u7_n167 ) );
  INV_X1 u1_u3_u7_U82 (.A( u1_u3_X_45 ) , .ZN( u1_u3_u7_n166 ) );
  NAND4_X1 u1_u3_u7_U83 (.ZN( u1_out3_5 ) , .A4( u1_u3_u7_n108 ) , .A3( u1_u3_u7_n109 ) , .A1( u1_u3_u7_n116 ) , .A2( u1_u3_u7_n123 ) );
  AOI22_X1 u1_u3_u7_U84 (.ZN( u1_u3_u7_n109 ) , .A2( u1_u3_u7_n126 ) , .B2( u1_u3_u7_n145 ) , .B1( u1_u3_u7_n156 ) , .A1( u1_u3_u7_n171 ) );
  NOR4_X1 u1_u3_u7_U85 (.A4( u1_u3_u7_n104 ) , .A3( u1_u3_u7_n105 ) , .A2( u1_u3_u7_n106 ) , .A1( u1_u3_u7_n107 ) , .ZN( u1_u3_u7_n108 ) );
  NAND4_X1 u1_u3_u7_U86 (.ZN( u1_out3_27 ) , .A4( u1_u3_u7_n118 ) , .A3( u1_u3_u7_n119 ) , .A2( u1_u3_u7_n120 ) , .A1( u1_u3_u7_n121 ) );
  OAI21_X1 u1_u3_u7_U87 (.ZN( u1_u3_u7_n121 ) , .B2( u1_u3_u7_n145 ) , .A( u1_u3_u7_n150 ) , .B1( u1_u3_u7_n174 ) );
  OAI21_X1 u1_u3_u7_U88 (.ZN( u1_u3_u7_n120 ) , .A( u1_u3_u7_n161 ) , .B2( u1_u3_u7_n170 ) , .B1( u1_u3_u7_n179 ) );
  NAND4_X1 u1_u3_u7_U89 (.ZN( u1_out3_21 ) , .A4( u1_u3_u7_n157 ) , .A3( u1_u3_u7_n158 ) , .A2( u1_u3_u7_n159 ) , .A1( u1_u3_u7_n160 ) );
  OAI221_X1 u1_u3_u7_U9 (.C1( u1_u3_u7_n101 ) , .C2( u1_u3_u7_n147 ) , .ZN( u1_u3_u7_n155 ) , .B2( u1_u3_u7_n162 ) , .A( u1_u3_u7_n91 ) , .B1( u1_u3_u7_n92 ) );
  OAI21_X1 u1_u3_u7_U90 (.B1( u1_u3_u7_n145 ) , .ZN( u1_u3_u7_n160 ) , .A( u1_u3_u7_n161 ) , .B2( u1_u3_u7_n177 ) );
  AOI22_X1 u1_u3_u7_U91 (.B2( u1_u3_u7_n149 ) , .B1( u1_u3_u7_n150 ) , .A2( u1_u3_u7_n151 ) , .A1( u1_u3_u7_n152 ) , .ZN( u1_u3_u7_n158 ) );
  NAND4_X1 u1_u3_u7_U92 (.ZN( u1_out3_15 ) , .A4( u1_u3_u7_n142 ) , .A3( u1_u3_u7_n143 ) , .A2( u1_u3_u7_n144 ) , .A1( u1_u3_u7_n178 ) );
  OR2_X1 u1_u3_u7_U93 (.A2( u1_u3_u7_n125 ) , .A1( u1_u3_u7_n129 ) , .ZN( u1_u3_u7_n144 ) );
  AOI22_X1 u1_u3_u7_U94 (.A2( u1_u3_u7_n126 ) , .ZN( u1_u3_u7_n143 ) , .B2( u1_u3_u7_n165 ) , .B1( u1_u3_u7_n173 ) , .A1( u1_u3_u7_n174 ) );
  NAND3_X1 u1_u3_u7_U95 (.A3( u1_u3_u7_n146 ) , .A2( u1_u3_u7_n147 ) , .A1( u1_u3_u7_n148 ) , .ZN( u1_u3_u7_n151 ) );
  NAND3_X1 u1_u3_u7_U96 (.A3( u1_u3_u7_n131 ) , .A2( u1_u3_u7_n132 ) , .A1( u1_u3_u7_n133 ) , .ZN( u1_u3_u7_n135 ) );
  XOR2_X1 u1_u5_U1 (.B( u1_K6_9 ) , .A( u1_R4_6 ) , .Z( u1_u5_X_9 ) );
  XOR2_X1 u1_u5_U48 (.B( u1_K6_10 ) , .A( u1_R4_7 ) , .Z( u1_u5_X_10 ) );
  AOI21_X1 u1_u5_u1_U10 (.B2( u1_u5_u1_n155 ) , .B1( u1_u5_u1_n156 ) , .ZN( u1_u5_u1_n157 ) , .A( u1_u5_u1_n174 ) );
  NAND3_X1 u1_u5_u1_U100 (.ZN( u1_u5_u1_n113 ) , .A1( u1_u5_u1_n120 ) , .A3( u1_u5_u1_n133 ) , .A2( u1_u5_u1_n155 ) );
  NAND2_X1 u1_u5_u1_U11 (.ZN( u1_u5_u1_n140 ) , .A2( u1_u5_u1_n150 ) , .A1( u1_u5_u1_n155 ) );
  NAND2_X1 u1_u5_u1_U12 (.A1( u1_u5_u1_n131 ) , .ZN( u1_u5_u1_n147 ) , .A2( u1_u5_u1_n153 ) );
  INV_X1 u1_u5_u1_U13 (.A( u1_u5_u1_n139 ) , .ZN( u1_u5_u1_n174 ) );
  OR4_X1 u1_u5_u1_U14 (.A4( u1_u5_u1_n106 ) , .A3( u1_u5_u1_n107 ) , .ZN( u1_u5_u1_n108 ) , .A1( u1_u5_u1_n117 ) , .A2( u1_u5_u1_n184 ) );
  AOI21_X1 u1_u5_u1_U15 (.ZN( u1_u5_u1_n106 ) , .A( u1_u5_u1_n112 ) , .B1( u1_u5_u1_n154 ) , .B2( u1_u5_u1_n156 ) );
  INV_X1 u1_u5_u1_U16 (.A( u1_u5_u1_n101 ) , .ZN( u1_u5_u1_n184 ) );
  AOI21_X1 u1_u5_u1_U17 (.ZN( u1_u5_u1_n107 ) , .B1( u1_u5_u1_n134 ) , .B2( u1_u5_u1_n149 ) , .A( u1_u5_u1_n174 ) );
  INV_X1 u1_u5_u1_U18 (.A( u1_u5_u1_n112 ) , .ZN( u1_u5_u1_n171 ) );
  NAND2_X1 u1_u5_u1_U19 (.ZN( u1_u5_u1_n141 ) , .A1( u1_u5_u1_n153 ) , .A2( u1_u5_u1_n156 ) );
  AND2_X1 u1_u5_u1_U20 (.A1( u1_u5_u1_n123 ) , .ZN( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n161 ) );
  NAND2_X1 u1_u5_u1_U21 (.A2( u1_u5_u1_n115 ) , .A1( u1_u5_u1_n116 ) , .ZN( u1_u5_u1_n148 ) );
  NAND2_X1 u1_u5_u1_U22 (.A2( u1_u5_u1_n133 ) , .A1( u1_u5_u1_n135 ) , .ZN( u1_u5_u1_n159 ) );
  NAND2_X1 u1_u5_u1_U23 (.A2( u1_u5_u1_n115 ) , .A1( u1_u5_u1_n120 ) , .ZN( u1_u5_u1_n132 ) );
  INV_X1 u1_u5_u1_U24 (.A( u1_u5_u1_n154 ) , .ZN( u1_u5_u1_n178 ) );
  AOI22_X1 u1_u5_u1_U25 (.B2( u1_u5_u1_n113 ) , .A2( u1_u5_u1_n114 ) , .ZN( u1_u5_u1_n125 ) , .A1( u1_u5_u1_n171 ) , .B1( u1_u5_u1_n173 ) );
  NAND2_X1 u1_u5_u1_U26 (.ZN( u1_u5_u1_n114 ) , .A1( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n156 ) );
  INV_X1 u1_u5_u1_U27 (.A( u1_u5_u1_n151 ) , .ZN( u1_u5_u1_n183 ) );
  AND2_X1 u1_u5_u1_U28 (.A1( u1_u5_u1_n129 ) , .A2( u1_u5_u1_n133 ) , .ZN( u1_u5_u1_n149 ) );
  INV_X1 u1_u5_u1_U29 (.A( u1_u5_u1_n131 ) , .ZN( u1_u5_u1_n180 ) );
  INV_X1 u1_u5_u1_U3 (.A( u1_u5_u1_n159 ) , .ZN( u1_u5_u1_n182 ) );
  OAI221_X1 u1_u5_u1_U30 (.A( u1_u5_u1_n119 ) , .C2( u1_u5_u1_n129 ) , .ZN( u1_u5_u1_n138 ) , .B2( u1_u5_u1_n152 ) , .C1( u1_u5_u1_n174 ) , .B1( u1_u5_u1_n187 ) );
  INV_X1 u1_u5_u1_U31 (.A( u1_u5_u1_n148 ) , .ZN( u1_u5_u1_n187 ) );
  AOI211_X1 u1_u5_u1_U32 (.B( u1_u5_u1_n117 ) , .A( u1_u5_u1_n118 ) , .ZN( u1_u5_u1_n119 ) , .C2( u1_u5_u1_n146 ) , .C1( u1_u5_u1_n159 ) );
  NOR2_X1 u1_u5_u1_U33 (.A1( u1_u5_u1_n168 ) , .A2( u1_u5_u1_n176 ) , .ZN( u1_u5_u1_n98 ) );
  AOI211_X1 u1_u5_u1_U34 (.B( u1_u5_u1_n162 ) , .A( u1_u5_u1_n163 ) , .C2( u1_u5_u1_n164 ) , .ZN( u1_u5_u1_n165 ) , .C1( u1_u5_u1_n171 ) );
  AOI21_X1 u1_u5_u1_U35 (.A( u1_u5_u1_n160 ) , .B2( u1_u5_u1_n161 ) , .ZN( u1_u5_u1_n162 ) , .B1( u1_u5_u1_n182 ) );
  OR2_X1 u1_u5_u1_U36 (.A2( u1_u5_u1_n157 ) , .A1( u1_u5_u1_n158 ) , .ZN( u1_u5_u1_n163 ) );
  OAI21_X1 u1_u5_u1_U37 (.B2( u1_u5_u1_n123 ) , .ZN( u1_u5_u1_n145 ) , .B1( u1_u5_u1_n160 ) , .A( u1_u5_u1_n185 ) );
  INV_X1 u1_u5_u1_U38 (.A( u1_u5_u1_n122 ) , .ZN( u1_u5_u1_n185 ) );
  AOI21_X1 u1_u5_u1_U39 (.B2( u1_u5_u1_n120 ) , .B1( u1_u5_u1_n121 ) , .ZN( u1_u5_u1_n122 ) , .A( u1_u5_u1_n128 ) );
  AOI221_X1 u1_u5_u1_U4 (.A( u1_u5_u1_n138 ) , .C2( u1_u5_u1_n139 ) , .C1( u1_u5_u1_n140 ) , .B2( u1_u5_u1_n141 ) , .ZN( u1_u5_u1_n142 ) , .B1( u1_u5_u1_n175 ) );
  NAND2_X1 u1_u5_u1_U40 (.A1( u1_u5_u1_n128 ) , .ZN( u1_u5_u1_n146 ) , .A2( u1_u5_u1_n160 ) );
  NAND2_X1 u1_u5_u1_U41 (.A2( u1_u5_u1_n112 ) , .ZN( u1_u5_u1_n139 ) , .A1( u1_u5_u1_n152 ) );
  NAND2_X1 u1_u5_u1_U42 (.A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n156 ) , .A2( u1_u5_u1_n99 ) );
  AOI221_X1 u1_u5_u1_U43 (.B1( u1_u5_u1_n140 ) , .ZN( u1_u5_u1_n167 ) , .B2( u1_u5_u1_n172 ) , .C2( u1_u5_u1_n175 ) , .C1( u1_u5_u1_n178 ) , .A( u1_u5_u1_n188 ) );
  INV_X1 u1_u5_u1_U44 (.ZN( u1_u5_u1_n188 ) , .A( u1_u5_u1_n97 ) );
  AOI211_X1 u1_u5_u1_U45 (.A( u1_u5_u1_n118 ) , .C1( u1_u5_u1_n132 ) , .C2( u1_u5_u1_n139 ) , .B( u1_u5_u1_n96 ) , .ZN( u1_u5_u1_n97 ) );
  AOI21_X1 u1_u5_u1_U46 (.B2( u1_u5_u1_n121 ) , .B1( u1_u5_u1_n135 ) , .A( u1_u5_u1_n152 ) , .ZN( u1_u5_u1_n96 ) );
  NOR2_X1 u1_u5_u1_U47 (.ZN( u1_u5_u1_n117 ) , .A1( u1_u5_u1_n121 ) , .A2( u1_u5_u1_n160 ) );
  AOI21_X1 u1_u5_u1_U48 (.A( u1_u5_u1_n128 ) , .B2( u1_u5_u1_n129 ) , .ZN( u1_u5_u1_n130 ) , .B1( u1_u5_u1_n150 ) );
  NAND2_X1 u1_u5_u1_U49 (.ZN( u1_u5_u1_n112 ) , .A1( u1_u5_u1_n169 ) , .A2( u1_u5_u1_n170 ) );
  AOI211_X1 u1_u5_u1_U5 (.ZN( u1_u5_u1_n124 ) , .A( u1_u5_u1_n138 ) , .C2( u1_u5_u1_n139 ) , .B( u1_u5_u1_n145 ) , .C1( u1_u5_u1_n147 ) );
  NAND2_X1 u1_u5_u1_U50 (.ZN( u1_u5_u1_n129 ) , .A2( u1_u5_u1_n95 ) , .A1( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U51 (.A1( u1_u5_u1_n102 ) , .ZN( u1_u5_u1_n154 ) , .A2( u1_u5_u1_n99 ) );
  NAND2_X1 u1_u5_u1_U52 (.A2( u1_u5_u1_n100 ) , .ZN( u1_u5_u1_n135 ) , .A1( u1_u5_u1_n99 ) );
  AOI21_X1 u1_u5_u1_U53 (.A( u1_u5_u1_n152 ) , .B2( u1_u5_u1_n153 ) , .B1( u1_u5_u1_n154 ) , .ZN( u1_u5_u1_n158 ) );
  INV_X1 u1_u5_u1_U54 (.A( u1_u5_u1_n160 ) , .ZN( u1_u5_u1_n175 ) );
  NAND2_X1 u1_u5_u1_U55 (.A1( u1_u5_u1_n100 ) , .ZN( u1_u5_u1_n116 ) , .A2( u1_u5_u1_n95 ) );
  NAND2_X1 u1_u5_u1_U56 (.A1( u1_u5_u1_n102 ) , .ZN( u1_u5_u1_n131 ) , .A2( u1_u5_u1_n95 ) );
  NAND2_X1 u1_u5_u1_U57 (.A2( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n121 ) , .A1( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U58 (.A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n153 ) , .A2( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U59 (.A2( u1_u5_u1_n104 ) , .A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n133 ) );
  AOI22_X1 u1_u5_u1_U6 (.B2( u1_u5_u1_n136 ) , .A2( u1_u5_u1_n137 ) , .ZN( u1_u5_u1_n143 ) , .A1( u1_u5_u1_n171 ) , .B1( u1_u5_u1_n173 ) );
  NAND2_X1 u1_u5_u1_U60 (.ZN( u1_u5_u1_n150 ) , .A2( u1_u5_u1_n98 ) , .A1( u1_u5_u1_n99 ) );
  NAND2_X1 u1_u5_u1_U61 (.A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n155 ) , .A2( u1_u5_u1_n95 ) );
  OAI21_X1 u1_u5_u1_U62 (.ZN( u1_u5_u1_n109 ) , .B1( u1_u5_u1_n129 ) , .B2( u1_u5_u1_n160 ) , .A( u1_u5_u1_n167 ) );
  NAND2_X1 u1_u5_u1_U63 (.A2( u1_u5_u1_n100 ) , .A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n120 ) );
  NAND2_X1 u1_u5_u1_U64 (.A1( u1_u5_u1_n102 ) , .A2( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n115 ) );
  NAND2_X1 u1_u5_u1_U65 (.A2( u1_u5_u1_n100 ) , .A1( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n151 ) );
  NAND2_X1 u1_u5_u1_U66 (.A2( u1_u5_u1_n103 ) , .A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n161 ) );
  INV_X1 u1_u5_u1_U67 (.A( u1_u5_u1_n152 ) , .ZN( u1_u5_u1_n173 ) );
  INV_X1 u1_u5_u1_U68 (.A( u1_u5_u1_n128 ) , .ZN( u1_u5_u1_n172 ) );
  NAND2_X1 u1_u5_u1_U69 (.A2( u1_u5_u1_n102 ) , .A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n123 ) );
  INV_X1 u1_u5_u1_U7 (.A( u1_u5_u1_n147 ) , .ZN( u1_u5_u1_n181 ) );
  NOR2_X1 u1_u5_u1_U70 (.A2( u1_u5_X_7 ) , .A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n95 ) );
  NOR2_X1 u1_u5_u1_U71 (.A1( u1_u5_X_12 ) , .A2( u1_u5_X_9 ) , .ZN( u1_u5_u1_n100 ) );
  NOR2_X1 u1_u5_u1_U72 (.A2( u1_u5_X_8 ) , .A1( u1_u5_u1_n177 ) , .ZN( u1_u5_u1_n99 ) );
  NOR2_X1 u1_u5_u1_U73 (.A2( u1_u5_X_12 ) , .ZN( u1_u5_u1_n102 ) , .A1( u1_u5_u1_n176 ) );
  NOR2_X1 u1_u5_u1_U74 (.A2( u1_u5_X_9 ) , .ZN( u1_u5_u1_n105 ) , .A1( u1_u5_u1_n168 ) );
  NAND2_X1 u1_u5_u1_U75 (.A1( u1_u5_X_10 ) , .ZN( u1_u5_u1_n160 ) , .A2( u1_u5_u1_n169 ) );
  NAND2_X1 u1_u5_u1_U76 (.A2( u1_u5_X_10 ) , .A1( u1_u5_X_11 ) , .ZN( u1_u5_u1_n152 ) );
  NAND2_X1 u1_u5_u1_U77 (.A1( u1_u5_X_11 ) , .ZN( u1_u5_u1_n128 ) , .A2( u1_u5_u1_n170 ) );
  AND2_X1 u1_u5_u1_U78 (.A2( u1_u5_X_7 ) , .A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n104 ) );
  AND2_X1 u1_u5_u1_U79 (.A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n103 ) , .A2( u1_u5_u1_n177 ) );
  NOR2_X1 u1_u5_u1_U8 (.A1( u1_u5_u1_n112 ) , .A2( u1_u5_u1_n116 ) , .ZN( u1_u5_u1_n118 ) );
  INV_X1 u1_u5_u1_U80 (.A( u1_u5_X_10 ) , .ZN( u1_u5_u1_n170 ) );
  INV_X1 u1_u5_u1_U81 (.A( u1_u5_X_9 ) , .ZN( u1_u5_u1_n176 ) );
  INV_X1 u1_u5_u1_U82 (.A( u1_u5_X_11 ) , .ZN( u1_u5_u1_n169 ) );
  INV_X1 u1_u5_u1_U83 (.A( u1_u5_X_12 ) , .ZN( u1_u5_u1_n168 ) );
  INV_X1 u1_u5_u1_U84 (.A( u1_u5_X_7 ) , .ZN( u1_u5_u1_n177 ) );
  NAND4_X1 u1_u5_u1_U85 (.ZN( u1_out5_18 ) , .A4( u1_u5_u1_n165 ) , .A3( u1_u5_u1_n166 ) , .A1( u1_u5_u1_n167 ) , .A2( u1_u5_u1_n186 ) );
  AOI22_X1 u1_u5_u1_U86 (.B2( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n147 ) , .A2( u1_u5_u1_n148 ) , .ZN( u1_u5_u1_n166 ) , .A1( u1_u5_u1_n172 ) );
  INV_X1 u1_u5_u1_U87 (.A( u1_u5_u1_n145 ) , .ZN( u1_u5_u1_n186 ) );
  OR4_X1 u1_u5_u1_U88 (.ZN( u1_out5_13 ) , .A4( u1_u5_u1_n108 ) , .A3( u1_u5_u1_n109 ) , .A2( u1_u5_u1_n110 ) , .A1( u1_u5_u1_n111 ) );
  AOI21_X1 u1_u5_u1_U89 (.ZN( u1_u5_u1_n110 ) , .A( u1_u5_u1_n116 ) , .B1( u1_u5_u1_n152 ) , .B2( u1_u5_u1_n160 ) );
  OAI21_X1 u1_u5_u1_U9 (.ZN( u1_u5_u1_n101 ) , .B1( u1_u5_u1_n141 ) , .A( u1_u5_u1_n146 ) , .B2( u1_u5_u1_n183 ) );
  AOI21_X1 u1_u5_u1_U90 (.ZN( u1_u5_u1_n111 ) , .A( u1_u5_u1_n128 ) , .B2( u1_u5_u1_n131 ) , .B1( u1_u5_u1_n135 ) );
  NAND4_X1 u1_u5_u1_U91 (.ZN( u1_out5_2 ) , .A4( u1_u5_u1_n142 ) , .A3( u1_u5_u1_n143 ) , .A2( u1_u5_u1_n144 ) , .A1( u1_u5_u1_n179 ) );
  OAI21_X1 u1_u5_u1_U92 (.B2( u1_u5_u1_n132 ) , .ZN( u1_u5_u1_n144 ) , .A( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n180 ) );
  INV_X1 u1_u5_u1_U93 (.A( u1_u5_u1_n130 ) , .ZN( u1_u5_u1_n179 ) );
  NAND4_X1 u1_u5_u1_U94 (.ZN( u1_out5_28 ) , .A4( u1_u5_u1_n124 ) , .A3( u1_u5_u1_n125 ) , .A2( u1_u5_u1_n126 ) , .A1( u1_u5_u1_n127 ) );
  OAI21_X1 u1_u5_u1_U95 (.ZN( u1_u5_u1_n127 ) , .B2( u1_u5_u1_n139 ) , .B1( u1_u5_u1_n175 ) , .A( u1_u5_u1_n183 ) );
  OAI21_X1 u1_u5_u1_U96 (.ZN( u1_u5_u1_n126 ) , .B2( u1_u5_u1_n140 ) , .A( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n178 ) );
  NAND3_X1 u1_u5_u1_U97 (.A3( u1_u5_u1_n149 ) , .A2( u1_u5_u1_n150 ) , .A1( u1_u5_u1_n151 ) , .ZN( u1_u5_u1_n164 ) );
  NAND3_X1 u1_u5_u1_U98 (.A3( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n135 ) , .ZN( u1_u5_u1_n136 ) , .A1( u1_u5_u1_n151 ) );
  NAND3_X1 u1_u5_u1_U99 (.A1( u1_u5_u1_n133 ) , .ZN( u1_u5_u1_n137 ) , .A2( u1_u5_u1_n154 ) , .A3( u1_u5_u1_n181 ) );
  XOR2_X1 u1_u7_U22 (.B( u1_K8_34 ) , .A( u1_R6_23 ) , .Z( u1_u7_X_34 ) );
  XOR2_X1 u1_u7_U23 (.B( u1_K8_33 ) , .A( u1_R6_22 ) , .Z( u1_u7_X_33 ) );
  INV_X1 u1_u7_u5_U10 (.A( u1_u7_u5_n121 ) , .ZN( u1_u7_u5_n177 ) );
  NOR3_X1 u1_u7_u5_U100 (.A3( u1_u7_u5_n141 ) , .A1( u1_u7_u5_n142 ) , .ZN( u1_u7_u5_n143 ) , .A2( u1_u7_u5_n191 ) );
  NAND4_X1 u1_u7_u5_U101 (.ZN( u1_out7_4 ) , .A4( u1_u7_u5_n112 ) , .A2( u1_u7_u5_n113 ) , .A1( u1_u7_u5_n114 ) , .A3( u1_u7_u5_n195 ) );
  AOI211_X1 u1_u7_u5_U102 (.A( u1_u7_u5_n110 ) , .C1( u1_u7_u5_n111 ) , .ZN( u1_u7_u5_n112 ) , .B( u1_u7_u5_n118 ) , .C2( u1_u7_u5_n177 ) );
  AOI222_X1 u1_u7_u5_U103 (.ZN( u1_u7_u5_n113 ) , .A1( u1_u7_u5_n131 ) , .C1( u1_u7_u5_n148 ) , .B2( u1_u7_u5_n174 ) , .C2( u1_u7_u5_n178 ) , .A2( u1_u7_u5_n179 ) , .B1( u1_u7_u5_n99 ) );
  NAND3_X1 u1_u7_u5_U104 (.A2( u1_u7_u5_n154 ) , .A3( u1_u7_u5_n158 ) , .A1( u1_u7_u5_n161 ) , .ZN( u1_u7_u5_n99 ) );
  NOR2_X1 u1_u7_u5_U11 (.ZN( u1_u7_u5_n160 ) , .A2( u1_u7_u5_n173 ) , .A1( u1_u7_u5_n177 ) );
  INV_X1 u1_u7_u5_U12 (.A( u1_u7_u5_n150 ) , .ZN( u1_u7_u5_n174 ) );
  AOI21_X1 u1_u7_u5_U13 (.A( u1_u7_u5_n160 ) , .B2( u1_u7_u5_n161 ) , .ZN( u1_u7_u5_n162 ) , .B1( u1_u7_u5_n192 ) );
  INV_X1 u1_u7_u5_U14 (.A( u1_u7_u5_n159 ) , .ZN( u1_u7_u5_n192 ) );
  AOI21_X1 u1_u7_u5_U15 (.A( u1_u7_u5_n156 ) , .B2( u1_u7_u5_n157 ) , .B1( u1_u7_u5_n158 ) , .ZN( u1_u7_u5_n163 ) );
  AOI21_X1 u1_u7_u5_U16 (.B2( u1_u7_u5_n139 ) , .B1( u1_u7_u5_n140 ) , .ZN( u1_u7_u5_n141 ) , .A( u1_u7_u5_n150 ) );
  OAI21_X1 u1_u7_u5_U17 (.A( u1_u7_u5_n133 ) , .B2( u1_u7_u5_n134 ) , .B1( u1_u7_u5_n135 ) , .ZN( u1_u7_u5_n142 ) );
  OAI21_X1 u1_u7_u5_U18 (.ZN( u1_u7_u5_n133 ) , .B2( u1_u7_u5_n147 ) , .A( u1_u7_u5_n173 ) , .B1( u1_u7_u5_n188 ) );
  NAND2_X1 u1_u7_u5_U19 (.A2( u1_u7_u5_n119 ) , .A1( u1_u7_u5_n123 ) , .ZN( u1_u7_u5_n137 ) );
  INV_X1 u1_u7_u5_U20 (.A( u1_u7_u5_n155 ) , .ZN( u1_u7_u5_n194 ) );
  NAND2_X1 u1_u7_u5_U21 (.A1( u1_u7_u5_n121 ) , .ZN( u1_u7_u5_n132 ) , .A2( u1_u7_u5_n172 ) );
  NAND2_X1 u1_u7_u5_U22 (.A2( u1_u7_u5_n122 ) , .ZN( u1_u7_u5_n136 ) , .A1( u1_u7_u5_n154 ) );
  NAND2_X1 u1_u7_u5_U23 (.A2( u1_u7_u5_n119 ) , .A1( u1_u7_u5_n120 ) , .ZN( u1_u7_u5_n159 ) );
  INV_X1 u1_u7_u5_U24 (.A( u1_u7_u5_n156 ) , .ZN( u1_u7_u5_n175 ) );
  INV_X1 u1_u7_u5_U25 (.A( u1_u7_u5_n158 ) , .ZN( u1_u7_u5_n188 ) );
  INV_X1 u1_u7_u5_U26 (.A( u1_u7_u5_n152 ) , .ZN( u1_u7_u5_n179 ) );
  INV_X1 u1_u7_u5_U27 (.A( u1_u7_u5_n140 ) , .ZN( u1_u7_u5_n182 ) );
  INV_X1 u1_u7_u5_U28 (.A( u1_u7_u5_n151 ) , .ZN( u1_u7_u5_n183 ) );
  INV_X1 u1_u7_u5_U29 (.A( u1_u7_u5_n123 ) , .ZN( u1_u7_u5_n185 ) );
  NOR2_X1 u1_u7_u5_U3 (.ZN( u1_u7_u5_n134 ) , .A1( u1_u7_u5_n183 ) , .A2( u1_u7_u5_n190 ) );
  INV_X1 u1_u7_u5_U30 (.A( u1_u7_u5_n161 ) , .ZN( u1_u7_u5_n184 ) );
  INV_X1 u1_u7_u5_U31 (.A( u1_u7_u5_n139 ) , .ZN( u1_u7_u5_n189 ) );
  INV_X1 u1_u7_u5_U32 (.A( u1_u7_u5_n157 ) , .ZN( u1_u7_u5_n190 ) );
  INV_X1 u1_u7_u5_U33 (.A( u1_u7_u5_n120 ) , .ZN( u1_u7_u5_n193 ) );
  NAND2_X1 u1_u7_u5_U34 (.ZN( u1_u7_u5_n111 ) , .A1( u1_u7_u5_n140 ) , .A2( u1_u7_u5_n155 ) );
  NOR2_X1 u1_u7_u5_U35 (.ZN( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n170 ) , .A2( u1_u7_u5_n180 ) );
  INV_X1 u1_u7_u5_U36 (.A( u1_u7_u5_n117 ) , .ZN( u1_u7_u5_n196 ) );
  OAI221_X1 u1_u7_u5_U37 (.A( u1_u7_u5_n116 ) , .ZN( u1_u7_u5_n117 ) , .B2( u1_u7_u5_n119 ) , .C1( u1_u7_u5_n153 ) , .C2( u1_u7_u5_n158 ) , .B1( u1_u7_u5_n172 ) );
  AOI222_X1 u1_u7_u5_U38 (.ZN( u1_u7_u5_n116 ) , .B2( u1_u7_u5_n145 ) , .C1( u1_u7_u5_n148 ) , .A2( u1_u7_u5_n174 ) , .C2( u1_u7_u5_n177 ) , .B1( u1_u7_u5_n187 ) , .A1( u1_u7_u5_n193 ) );
  INV_X1 u1_u7_u5_U39 (.A( u1_u7_u5_n115 ) , .ZN( u1_u7_u5_n187 ) );
  INV_X1 u1_u7_u5_U4 (.A( u1_u7_u5_n138 ) , .ZN( u1_u7_u5_n191 ) );
  AOI22_X1 u1_u7_u5_U40 (.B2( u1_u7_u5_n131 ) , .A2( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n169 ) , .B1( u1_u7_u5_n174 ) , .A1( u1_u7_u5_n185 ) );
  NOR2_X1 u1_u7_u5_U41 (.A1( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n150 ) , .A2( u1_u7_u5_n173 ) );
  AOI21_X1 u1_u7_u5_U42 (.A( u1_u7_u5_n118 ) , .B2( u1_u7_u5_n145 ) , .ZN( u1_u7_u5_n168 ) , .B1( u1_u7_u5_n186 ) );
  INV_X1 u1_u7_u5_U43 (.A( u1_u7_u5_n122 ) , .ZN( u1_u7_u5_n186 ) );
  NOR2_X1 u1_u7_u5_U44 (.A1( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n152 ) , .A2( u1_u7_u5_n176 ) );
  NOR2_X1 u1_u7_u5_U45 (.A1( u1_u7_u5_n115 ) , .ZN( u1_u7_u5_n118 ) , .A2( u1_u7_u5_n153 ) );
  NOR2_X1 u1_u7_u5_U46 (.A2( u1_u7_u5_n145 ) , .ZN( u1_u7_u5_n156 ) , .A1( u1_u7_u5_n174 ) );
  NOR2_X1 u1_u7_u5_U47 (.ZN( u1_u7_u5_n121 ) , .A2( u1_u7_u5_n145 ) , .A1( u1_u7_u5_n176 ) );
  AOI22_X1 u1_u7_u5_U48 (.ZN( u1_u7_u5_n114 ) , .A2( u1_u7_u5_n137 ) , .A1( u1_u7_u5_n145 ) , .B2( u1_u7_u5_n175 ) , .B1( u1_u7_u5_n193 ) );
  OAI211_X1 u1_u7_u5_U49 (.B( u1_u7_u5_n124 ) , .A( u1_u7_u5_n125 ) , .C2( u1_u7_u5_n126 ) , .C1( u1_u7_u5_n127 ) , .ZN( u1_u7_u5_n128 ) );
  OAI21_X1 u1_u7_u5_U5 (.B2( u1_u7_u5_n136 ) , .B1( u1_u7_u5_n137 ) , .ZN( u1_u7_u5_n138 ) , .A( u1_u7_u5_n177 ) );
  NOR3_X1 u1_u7_u5_U50 (.ZN( u1_u7_u5_n127 ) , .A1( u1_u7_u5_n136 ) , .A3( u1_u7_u5_n148 ) , .A2( u1_u7_u5_n182 ) );
  OAI21_X1 u1_u7_u5_U51 (.ZN( u1_u7_u5_n124 ) , .A( u1_u7_u5_n177 ) , .B2( u1_u7_u5_n183 ) , .B1( u1_u7_u5_n189 ) );
  OAI21_X1 u1_u7_u5_U52 (.ZN( u1_u7_u5_n125 ) , .A( u1_u7_u5_n174 ) , .B2( u1_u7_u5_n185 ) , .B1( u1_u7_u5_n190 ) );
  AOI21_X1 u1_u7_u5_U53 (.A( u1_u7_u5_n153 ) , .B2( u1_u7_u5_n154 ) , .B1( u1_u7_u5_n155 ) , .ZN( u1_u7_u5_n164 ) );
  AOI21_X1 u1_u7_u5_U54 (.ZN( u1_u7_u5_n110 ) , .B1( u1_u7_u5_n122 ) , .B2( u1_u7_u5_n139 ) , .A( u1_u7_u5_n153 ) );
  INV_X1 u1_u7_u5_U55 (.A( u1_u7_u5_n153 ) , .ZN( u1_u7_u5_n176 ) );
  INV_X1 u1_u7_u5_U56 (.A( u1_u7_u5_n126 ) , .ZN( u1_u7_u5_n173 ) );
  AND2_X1 u1_u7_u5_U57 (.A2( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n107 ) , .ZN( u1_u7_u5_n147 ) );
  AND2_X1 u1_u7_u5_U58 (.A2( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n108 ) , .ZN( u1_u7_u5_n148 ) );
  NAND2_X1 u1_u7_u5_U59 (.A1( u1_u7_u5_n105 ) , .A2( u1_u7_u5_n106 ) , .ZN( u1_u7_u5_n158 ) );
  INV_X1 u1_u7_u5_U6 (.A( u1_u7_u5_n135 ) , .ZN( u1_u7_u5_n178 ) );
  NAND2_X1 u1_u7_u5_U60 (.A2( u1_u7_u5_n108 ) , .A1( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n139 ) );
  NAND2_X1 u1_u7_u5_U61 (.A1( u1_u7_u5_n106 ) , .A2( u1_u7_u5_n108 ) , .ZN( u1_u7_u5_n119 ) );
  NAND2_X1 u1_u7_u5_U62 (.A2( u1_u7_u5_n103 ) , .A1( u1_u7_u5_n105 ) , .ZN( u1_u7_u5_n140 ) );
  NAND2_X1 u1_u7_u5_U63 (.A2( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n105 ) , .ZN( u1_u7_u5_n155 ) );
  NAND2_X1 u1_u7_u5_U64 (.A2( u1_u7_u5_n106 ) , .A1( u1_u7_u5_n107 ) , .ZN( u1_u7_u5_n122 ) );
  NAND2_X1 u1_u7_u5_U65 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n106 ) , .ZN( u1_u7_u5_n115 ) );
  NAND2_X1 u1_u7_u5_U66 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n103 ) , .ZN( u1_u7_u5_n161 ) );
  NAND2_X1 u1_u7_u5_U67 (.A1( u1_u7_u5_n105 ) , .A2( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n154 ) );
  INV_X1 u1_u7_u5_U68 (.A( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n172 ) );
  NAND2_X1 u1_u7_u5_U69 (.A1( u1_u7_u5_n103 ) , .A2( u1_u7_u5_n108 ) , .ZN( u1_u7_u5_n123 ) );
  OAI22_X1 u1_u7_u5_U7 (.B2( u1_u7_u5_n149 ) , .B1( u1_u7_u5_n150 ) , .A2( u1_u7_u5_n151 ) , .A1( u1_u7_u5_n152 ) , .ZN( u1_u7_u5_n165 ) );
  NAND2_X1 u1_u7_u5_U70 (.A2( u1_u7_u5_n103 ) , .A1( u1_u7_u5_n107 ) , .ZN( u1_u7_u5_n151 ) );
  NAND2_X1 u1_u7_u5_U71 (.A2( u1_u7_u5_n107 ) , .A1( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n120 ) );
  NAND2_X1 u1_u7_u5_U72 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n157 ) );
  AND2_X1 u1_u7_u5_U73 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n104 ) , .ZN( u1_u7_u5_n131 ) );
  INV_X1 u1_u7_u5_U74 (.A( u1_u7_u5_n102 ) , .ZN( u1_u7_u5_n195 ) );
  OAI221_X1 u1_u7_u5_U75 (.A( u1_u7_u5_n101 ) , .ZN( u1_u7_u5_n102 ) , .C2( u1_u7_u5_n115 ) , .C1( u1_u7_u5_n126 ) , .B1( u1_u7_u5_n134 ) , .B2( u1_u7_u5_n160 ) );
  OAI21_X1 u1_u7_u5_U76 (.ZN( u1_u7_u5_n101 ) , .B1( u1_u7_u5_n137 ) , .A( u1_u7_u5_n146 ) , .B2( u1_u7_u5_n147 ) );
  NOR2_X1 u1_u7_u5_U77 (.A2( u1_u7_X_34 ) , .A1( u1_u7_X_35 ) , .ZN( u1_u7_u5_n145 ) );
  NOR2_X1 u1_u7_u5_U78 (.A2( u1_u7_X_34 ) , .ZN( u1_u7_u5_n146 ) , .A1( u1_u7_u5_n171 ) );
  NOR2_X1 u1_u7_u5_U79 (.A2( u1_u7_X_31 ) , .A1( u1_u7_X_32 ) , .ZN( u1_u7_u5_n103 ) );
  NOR3_X1 u1_u7_u5_U8 (.A2( u1_u7_u5_n147 ) , .A1( u1_u7_u5_n148 ) , .ZN( u1_u7_u5_n149 ) , .A3( u1_u7_u5_n194 ) );
  NOR2_X1 u1_u7_u5_U80 (.A2( u1_u7_X_36 ) , .ZN( u1_u7_u5_n105 ) , .A1( u1_u7_u5_n180 ) );
  NOR2_X1 u1_u7_u5_U81 (.A2( u1_u7_X_33 ) , .ZN( u1_u7_u5_n108 ) , .A1( u1_u7_u5_n170 ) );
  NOR2_X1 u1_u7_u5_U82 (.A2( u1_u7_X_33 ) , .A1( u1_u7_X_36 ) , .ZN( u1_u7_u5_n107 ) );
  NOR2_X1 u1_u7_u5_U83 (.A2( u1_u7_X_31 ) , .ZN( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n181 ) );
  NAND2_X1 u1_u7_u5_U84 (.A2( u1_u7_X_34 ) , .A1( u1_u7_X_35 ) , .ZN( u1_u7_u5_n153 ) );
  NAND2_X1 u1_u7_u5_U85 (.A1( u1_u7_X_34 ) , .ZN( u1_u7_u5_n126 ) , .A2( u1_u7_u5_n171 ) );
  AND2_X1 u1_u7_u5_U86 (.A1( u1_u7_X_31 ) , .A2( u1_u7_X_32 ) , .ZN( u1_u7_u5_n106 ) );
  AND2_X1 u1_u7_u5_U87 (.A1( u1_u7_X_31 ) , .ZN( u1_u7_u5_n109 ) , .A2( u1_u7_u5_n181 ) );
  INV_X1 u1_u7_u5_U88 (.A( u1_u7_X_33 ) , .ZN( u1_u7_u5_n180 ) );
  INV_X1 u1_u7_u5_U89 (.A( u1_u7_X_35 ) , .ZN( u1_u7_u5_n171 ) );
  NOR2_X1 u1_u7_u5_U9 (.ZN( u1_u7_u5_n135 ) , .A1( u1_u7_u5_n173 ) , .A2( u1_u7_u5_n176 ) );
  INV_X1 u1_u7_u5_U90 (.A( u1_u7_X_36 ) , .ZN( u1_u7_u5_n170 ) );
  INV_X1 u1_u7_u5_U91 (.A( u1_u7_X_32 ) , .ZN( u1_u7_u5_n181 ) );
  NAND4_X1 u1_u7_u5_U92 (.ZN( u1_out7_29 ) , .A4( u1_u7_u5_n129 ) , .A3( u1_u7_u5_n130 ) , .A2( u1_u7_u5_n168 ) , .A1( u1_u7_u5_n196 ) );
  AOI221_X1 u1_u7_u5_U93 (.A( u1_u7_u5_n128 ) , .ZN( u1_u7_u5_n129 ) , .C2( u1_u7_u5_n132 ) , .B2( u1_u7_u5_n159 ) , .B1( u1_u7_u5_n176 ) , .C1( u1_u7_u5_n184 ) );
  AOI222_X1 u1_u7_u5_U94 (.ZN( u1_u7_u5_n130 ) , .A2( u1_u7_u5_n146 ) , .B1( u1_u7_u5_n147 ) , .C2( u1_u7_u5_n175 ) , .B2( u1_u7_u5_n179 ) , .A1( u1_u7_u5_n188 ) , .C1( u1_u7_u5_n194 ) );
  NAND4_X1 u1_u7_u5_U95 (.ZN( u1_out7_19 ) , .A4( u1_u7_u5_n166 ) , .A3( u1_u7_u5_n167 ) , .A2( u1_u7_u5_n168 ) , .A1( u1_u7_u5_n169 ) );
  AOI22_X1 u1_u7_u5_U96 (.B2( u1_u7_u5_n145 ) , .A2( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n167 ) , .B1( u1_u7_u5_n182 ) , .A1( u1_u7_u5_n189 ) );
  NOR4_X1 u1_u7_u5_U97 (.A4( u1_u7_u5_n162 ) , .A3( u1_u7_u5_n163 ) , .A2( u1_u7_u5_n164 ) , .A1( u1_u7_u5_n165 ) , .ZN( u1_u7_u5_n166 ) );
  NAND4_X1 u1_u7_u5_U98 (.ZN( u1_out7_11 ) , .A4( u1_u7_u5_n143 ) , .A3( u1_u7_u5_n144 ) , .A2( u1_u7_u5_n169 ) , .A1( u1_u7_u5_n196 ) );
  AOI22_X1 u1_u7_u5_U99 (.A2( u1_u7_u5_n132 ) , .ZN( u1_u7_u5_n144 ) , .B2( u1_u7_u5_n145 ) , .B1( u1_u7_u5_n184 ) , .A1( u1_u7_u5_n194 ) );
  INV_X1 u1_uk_U1117 (.ZN( u1_K13_10 ) , .A( u1_uk_n671 ) );
  INV_X1 u1_uk_U141 (.ZN( u1_K13_15 ) , .A( u1_uk_n678 ) );
  INV_X1 u1_uk_U218 (.ZN( u1_K4_31 ) , .A( u1_uk_n1063 ) );
  INV_X1 u1_uk_U449 (.ZN( u1_K6_9 ) , .A( u1_uk_n1104 ) );
  INV_X1 u1_uk_U501 (.ZN( u1_K4_29 ) , .A( u1_uk_n1060 ) );
  INV_X1 u1_uk_U590 (.ZN( u1_K6_10 ) , .A( u1_uk_n1088 ) );
  INV_X1 u1_uk_U642 (.ZN( u1_K13_11 ) , .A( u1_uk_n672 ) );
  INV_X1 u1_uk_U71 (.ZN( u1_K8_34 ) , .A( u1_uk_n1137 ) );
  INV_X1 u1_uk_U781 (.ZN( u1_K13_13 ) , .A( u1_uk_n677 ) );
  XOR2_X1 u2_U309 (.B( u2_L6_31 ) , .Z( u2_N254 ) , .A( u2_out7_31 ) );
  XOR2_X1 u2_U318 (.B( u2_L6_23 ) , .Z( u2_N246 ) , .A( u2_out7_23 ) );
  XOR2_X1 u2_U324 (.B( u2_L6_17 ) , .Z( u2_N240 ) , .A( u2_out7_17 ) );
  XOR2_X1 u2_U333 (.B( u2_L6_9 ) , .Z( u2_N232 ) , .A( u2_out7_9 ) );
  XOR2_X1 u2_U382 (.B( u2_L4_30 ) , .Z( u2_N189 ) , .A( u2_out5_30 ) );
  XOR2_X1 u2_U388 (.B( u2_L4_24 ) , .Z( u2_N183 ) , .A( u2_out5_24 ) );
  XOR2_X1 u2_U397 (.B( u2_L4_16 ) , .Z( u2_N175 ) , .A( u2_out5_16 ) );
  XOR2_X1 u2_U408 (.B( u2_L4_6 ) , .Z( u2_N165 ) , .A( u2_out5_6 ) );
  XOR2_X1 u2_u5_U40 (.B( u2_K6_18 ) , .A( u2_R4_13 ) , .Z( u2_u5_X_18 ) );
  XOR2_X1 u2_u5_U41 (.B( u2_K6_17 ) , .A( u2_R4_12 ) , .Z( u2_u5_X_17 ) );
  XOR2_X1 u2_u5_U42 (.B( u2_K6_16 ) , .A( u2_R4_11 ) , .Z( u2_u5_X_16 ) );
  XOR2_X1 u2_u5_U43 (.B( u2_K6_15 ) , .A( u2_R4_10 ) , .Z( u2_u5_X_15 ) );
  XOR2_X1 u2_u5_U44 (.B( u2_K6_14 ) , .A( u2_R4_9 ) , .Z( u2_u5_X_14 ) );
  XOR2_X1 u2_u5_U45 (.B( u2_K6_13 ) , .A( u2_R4_8 ) , .Z( u2_u5_X_13 ) );
  OAI22_X1 u2_u5_u2_U10 (.ZN( u2_u5_u2_n109 ) , .A2( u2_u5_u2_n113 ) , .B2( u2_u5_u2_n133 ) , .B1( u2_u5_u2_n167 ) , .A1( u2_u5_u2_n168 ) );
  NAND3_X1 u2_u5_u2_U100 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n98 ) );
  OAI22_X1 u2_u5_u2_U11 (.B1( u2_u5_u2_n151 ) , .A2( u2_u5_u2_n152 ) , .A1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n160 ) , .B2( u2_u5_u2_n168 ) );
  NOR3_X1 u2_u5_u2_U12 (.A1( u2_u5_u2_n150 ) , .ZN( u2_u5_u2_n151 ) , .A3( u2_u5_u2_n175 ) , .A2( u2_u5_u2_n188 ) );
  AOI21_X1 u2_u5_u2_U13 (.ZN( u2_u5_u2_n144 ) , .B2( u2_u5_u2_n155 ) , .A( u2_u5_u2_n172 ) , .B1( u2_u5_u2_n185 ) );
  AOI21_X1 u2_u5_u2_U14 (.B2( u2_u5_u2_n143 ) , .ZN( u2_u5_u2_n145 ) , .B1( u2_u5_u2_n152 ) , .A( u2_u5_u2_n171 ) );
  AOI21_X1 u2_u5_u2_U15 (.B2( u2_u5_u2_n120 ) , .B1( u2_u5_u2_n121 ) , .ZN( u2_u5_u2_n126 ) , .A( u2_u5_u2_n167 ) );
  INV_X1 u2_u5_u2_U16 (.A( u2_u5_u2_n156 ) , .ZN( u2_u5_u2_n171 ) );
  INV_X1 u2_u5_u2_U17 (.A( u2_u5_u2_n120 ) , .ZN( u2_u5_u2_n188 ) );
  NAND2_X1 u2_u5_u2_U18 (.A2( u2_u5_u2_n122 ) , .ZN( u2_u5_u2_n150 ) , .A1( u2_u5_u2_n152 ) );
  INV_X1 u2_u5_u2_U19 (.A( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n170 ) );
  INV_X1 u2_u5_u2_U20 (.A( u2_u5_u2_n137 ) , .ZN( u2_u5_u2_n173 ) );
  NAND2_X1 u2_u5_u2_U21 (.A1( u2_u5_u2_n132 ) , .A2( u2_u5_u2_n139 ) , .ZN( u2_u5_u2_n157 ) );
  INV_X1 u2_u5_u2_U22 (.A( u2_u5_u2_n113 ) , .ZN( u2_u5_u2_n178 ) );
  INV_X1 u2_u5_u2_U23 (.A( u2_u5_u2_n139 ) , .ZN( u2_u5_u2_n175 ) );
  INV_X1 u2_u5_u2_U24 (.A( u2_u5_u2_n155 ) , .ZN( u2_u5_u2_n181 ) );
  INV_X1 u2_u5_u2_U25 (.A( u2_u5_u2_n119 ) , .ZN( u2_u5_u2_n177 ) );
  INV_X1 u2_u5_u2_U26 (.A( u2_u5_u2_n116 ) , .ZN( u2_u5_u2_n180 ) );
  INV_X1 u2_u5_u2_U27 (.A( u2_u5_u2_n131 ) , .ZN( u2_u5_u2_n179 ) );
  INV_X1 u2_u5_u2_U28 (.A( u2_u5_u2_n154 ) , .ZN( u2_u5_u2_n176 ) );
  NAND2_X1 u2_u5_u2_U29 (.A2( u2_u5_u2_n116 ) , .A1( u2_u5_u2_n117 ) , .ZN( u2_u5_u2_n118 ) );
  NOR2_X1 u2_u5_u2_U3 (.ZN( u2_u5_u2_n121 ) , .A2( u2_u5_u2_n177 ) , .A1( u2_u5_u2_n180 ) );
  INV_X1 u2_u5_u2_U30 (.A( u2_u5_u2_n132 ) , .ZN( u2_u5_u2_n182 ) );
  INV_X1 u2_u5_u2_U31 (.A( u2_u5_u2_n158 ) , .ZN( u2_u5_u2_n183 ) );
  OAI21_X1 u2_u5_u2_U32 (.A( u2_u5_u2_n156 ) , .B1( u2_u5_u2_n157 ) , .ZN( u2_u5_u2_n158 ) , .B2( u2_u5_u2_n179 ) );
  NOR2_X1 u2_u5_u2_U33 (.ZN( u2_u5_u2_n156 ) , .A1( u2_u5_u2_n166 ) , .A2( u2_u5_u2_n169 ) );
  NOR2_X1 u2_u5_u2_U34 (.A2( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n137 ) , .A1( u2_u5_u2_n140 ) );
  NOR2_X1 u2_u5_u2_U35 (.A2( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n153 ) , .A1( u2_u5_u2_n156 ) );
  AOI211_X1 u2_u5_u2_U36 (.ZN( u2_u5_u2_n130 ) , .C1( u2_u5_u2_n138 ) , .C2( u2_u5_u2_n179 ) , .B( u2_u5_u2_n96 ) , .A( u2_u5_u2_n97 ) );
  OAI22_X1 u2_u5_u2_U37 (.B1( u2_u5_u2_n133 ) , .A2( u2_u5_u2_n137 ) , .A1( u2_u5_u2_n152 ) , .B2( u2_u5_u2_n168 ) , .ZN( u2_u5_u2_n97 ) );
  OAI221_X1 u2_u5_u2_U38 (.B1( u2_u5_u2_n113 ) , .C1( u2_u5_u2_n132 ) , .A( u2_u5_u2_n149 ) , .B2( u2_u5_u2_n171 ) , .C2( u2_u5_u2_n172 ) , .ZN( u2_u5_u2_n96 ) );
  OAI221_X1 u2_u5_u2_U39 (.A( u2_u5_u2_n115 ) , .C2( u2_u5_u2_n123 ) , .B2( u2_u5_u2_n143 ) , .B1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n163 ) , .C1( u2_u5_u2_n168 ) );
  INV_X1 u2_u5_u2_U4 (.A( u2_u5_u2_n134 ) , .ZN( u2_u5_u2_n185 ) );
  OAI21_X1 u2_u5_u2_U40 (.A( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n115 ) , .B1( u2_u5_u2_n176 ) , .B2( u2_u5_u2_n178 ) );
  OAI221_X1 u2_u5_u2_U41 (.A( u2_u5_u2_n135 ) , .B2( u2_u5_u2_n136 ) , .B1( u2_u5_u2_n137 ) , .ZN( u2_u5_u2_n162 ) , .C2( u2_u5_u2_n167 ) , .C1( u2_u5_u2_n185 ) );
  AND3_X1 u2_u5_u2_U42 (.A3( u2_u5_u2_n131 ) , .A2( u2_u5_u2_n132 ) , .A1( u2_u5_u2_n133 ) , .ZN( u2_u5_u2_n136 ) );
  AOI22_X1 u2_u5_u2_U43 (.ZN( u2_u5_u2_n135 ) , .B1( u2_u5_u2_n140 ) , .A1( u2_u5_u2_n156 ) , .B2( u2_u5_u2_n180 ) , .A2( u2_u5_u2_n188 ) );
  AOI21_X1 u2_u5_u2_U44 (.ZN( u2_u5_u2_n149 ) , .B1( u2_u5_u2_n173 ) , .B2( u2_u5_u2_n188 ) , .A( u2_u5_u2_n95 ) );
  AND3_X1 u2_u5_u2_U45 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n156 ) , .ZN( u2_u5_u2_n95 ) );
  OAI21_X1 u2_u5_u2_U46 (.A( u2_u5_u2_n141 ) , .B2( u2_u5_u2_n142 ) , .ZN( u2_u5_u2_n146 ) , .B1( u2_u5_u2_n153 ) );
  OAI21_X1 u2_u5_u2_U47 (.A( u2_u5_u2_n140 ) , .ZN( u2_u5_u2_n141 ) , .B1( u2_u5_u2_n176 ) , .B2( u2_u5_u2_n177 ) );
  NOR3_X1 u2_u5_u2_U48 (.ZN( u2_u5_u2_n142 ) , .A3( u2_u5_u2_n175 ) , .A2( u2_u5_u2_n178 ) , .A1( u2_u5_u2_n181 ) );
  OAI21_X1 u2_u5_u2_U49 (.A( u2_u5_u2_n101 ) , .B2( u2_u5_u2_n121 ) , .B1( u2_u5_u2_n153 ) , .ZN( u2_u5_u2_n164 ) );
  INV_X1 u2_u5_u2_U5 (.A( u2_u5_u2_n150 ) , .ZN( u2_u5_u2_n184 ) );
  NAND2_X1 u2_u5_u2_U50 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n155 ) );
  NAND2_X1 u2_u5_u2_U51 (.A2( u2_u5_u2_n105 ) , .A1( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n143 ) );
  NAND2_X1 u2_u5_u2_U52 (.A1( u2_u5_u2_n104 ) , .A2( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n152 ) );
  NAND2_X1 u2_u5_u2_U53 (.A1( u2_u5_u2_n100 ) , .A2( u2_u5_u2_n105 ) , .ZN( u2_u5_u2_n132 ) );
  INV_X1 u2_u5_u2_U54 (.A( u2_u5_u2_n140 ) , .ZN( u2_u5_u2_n168 ) );
  INV_X1 u2_u5_u2_U55 (.A( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n167 ) );
  NAND2_X1 u2_u5_u2_U56 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n113 ) );
  NAND2_X1 u2_u5_u2_U57 (.A1( u2_u5_u2_n106 ) , .A2( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n131 ) );
  NAND2_X1 u2_u5_u2_U58 (.A1( u2_u5_u2_n103 ) , .A2( u2_u5_u2_n107 ) , .ZN( u2_u5_u2_n139 ) );
  NAND2_X1 u2_u5_u2_U59 (.A1( u2_u5_u2_n103 ) , .A2( u2_u5_u2_n105 ) , .ZN( u2_u5_u2_n133 ) );
  NOR4_X1 u2_u5_u2_U6 (.A4( u2_u5_u2_n124 ) , .A3( u2_u5_u2_n125 ) , .A2( u2_u5_u2_n126 ) , .A1( u2_u5_u2_n127 ) , .ZN( u2_u5_u2_n128 ) );
  NAND2_X1 u2_u5_u2_U60 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n103 ) , .ZN( u2_u5_u2_n154 ) );
  NAND2_X1 u2_u5_u2_U61 (.A2( u2_u5_u2_n103 ) , .A1( u2_u5_u2_n104 ) , .ZN( u2_u5_u2_n119 ) );
  NAND2_X1 u2_u5_u2_U62 (.A2( u2_u5_u2_n107 ) , .A1( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n123 ) );
  NAND2_X1 u2_u5_u2_U63 (.A1( u2_u5_u2_n104 ) , .A2( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n122 ) );
  INV_X1 u2_u5_u2_U64 (.A( u2_u5_u2_n114 ) , .ZN( u2_u5_u2_n172 ) );
  NAND2_X1 u2_u5_u2_U65 (.A2( u2_u5_u2_n100 ) , .A1( u2_u5_u2_n102 ) , .ZN( u2_u5_u2_n116 ) );
  NAND2_X1 u2_u5_u2_U66 (.A1( u2_u5_u2_n102 ) , .A2( u2_u5_u2_n108 ) , .ZN( u2_u5_u2_n120 ) );
  NAND2_X1 u2_u5_u2_U67 (.A2( u2_u5_u2_n105 ) , .A1( u2_u5_u2_n106 ) , .ZN( u2_u5_u2_n117 ) );
  INV_X1 u2_u5_u2_U68 (.ZN( u2_u5_u2_n187 ) , .A( u2_u5_u2_n99 ) );
  OAI21_X1 u2_u5_u2_U69 (.B1( u2_u5_u2_n137 ) , .B2( u2_u5_u2_n143 ) , .A( u2_u5_u2_n98 ) , .ZN( u2_u5_u2_n99 ) );
  AOI21_X1 u2_u5_u2_U7 (.B2( u2_u5_u2_n119 ) , .ZN( u2_u5_u2_n127 ) , .A( u2_u5_u2_n137 ) , .B1( u2_u5_u2_n155 ) );
  NOR2_X1 u2_u5_u2_U70 (.A2( u2_u5_X_16 ) , .ZN( u2_u5_u2_n140 ) , .A1( u2_u5_u2_n166 ) );
  NOR2_X1 u2_u5_u2_U71 (.A2( u2_u5_X_13 ) , .A1( u2_u5_X_14 ) , .ZN( u2_u5_u2_n100 ) );
  NOR2_X1 u2_u5_u2_U72 (.A2( u2_u5_X_16 ) , .A1( u2_u5_X_17 ) , .ZN( u2_u5_u2_n138 ) );
  NOR2_X1 u2_u5_u2_U73 (.A2( u2_u5_X_15 ) , .A1( u2_u5_X_18 ) , .ZN( u2_u5_u2_n104 ) );
  NOR2_X1 u2_u5_u2_U74 (.A2( u2_u5_X_14 ) , .ZN( u2_u5_u2_n103 ) , .A1( u2_u5_u2_n174 ) );
  NOR2_X1 u2_u5_u2_U75 (.A2( u2_u5_X_15 ) , .ZN( u2_u5_u2_n102 ) , .A1( u2_u5_u2_n165 ) );
  NOR2_X1 u2_u5_u2_U76 (.A2( u2_u5_X_17 ) , .ZN( u2_u5_u2_n114 ) , .A1( u2_u5_u2_n169 ) );
  AND2_X1 u2_u5_u2_U77 (.A1( u2_u5_X_15 ) , .ZN( u2_u5_u2_n105 ) , .A2( u2_u5_u2_n165 ) );
  AND2_X1 u2_u5_u2_U78 (.A2( u2_u5_X_15 ) , .A1( u2_u5_X_18 ) , .ZN( u2_u5_u2_n107 ) );
  AND2_X1 u2_u5_u2_U79 (.A1( u2_u5_X_14 ) , .ZN( u2_u5_u2_n106 ) , .A2( u2_u5_u2_n174 ) );
  AOI21_X1 u2_u5_u2_U8 (.ZN( u2_u5_u2_n124 ) , .B1( u2_u5_u2_n131 ) , .B2( u2_u5_u2_n143 ) , .A( u2_u5_u2_n172 ) );
  AND2_X1 u2_u5_u2_U80 (.A1( u2_u5_X_13 ) , .A2( u2_u5_X_14 ) , .ZN( u2_u5_u2_n108 ) );
  INV_X1 u2_u5_u2_U81 (.A( u2_u5_X_16 ) , .ZN( u2_u5_u2_n169 ) );
  INV_X1 u2_u5_u2_U82 (.A( u2_u5_X_17 ) , .ZN( u2_u5_u2_n166 ) );
  INV_X1 u2_u5_u2_U83 (.A( u2_u5_X_13 ) , .ZN( u2_u5_u2_n174 ) );
  INV_X1 u2_u5_u2_U84 (.A( u2_u5_X_18 ) , .ZN( u2_u5_u2_n165 ) );
  NAND4_X1 u2_u5_u2_U85 (.ZN( u2_out5_24 ) , .A4( u2_u5_u2_n111 ) , .A3( u2_u5_u2_n112 ) , .A1( u2_u5_u2_n130 ) , .A2( u2_u5_u2_n187 ) );
  AOI221_X1 u2_u5_u2_U86 (.A( u2_u5_u2_n109 ) , .B1( u2_u5_u2_n110 ) , .ZN( u2_u5_u2_n111 ) , .C1( u2_u5_u2_n134 ) , .C2( u2_u5_u2_n170 ) , .B2( u2_u5_u2_n173 ) );
  AOI21_X1 u2_u5_u2_U87 (.ZN( u2_u5_u2_n112 ) , .B2( u2_u5_u2_n156 ) , .A( u2_u5_u2_n164 ) , .B1( u2_u5_u2_n181 ) );
  NAND4_X1 u2_u5_u2_U88 (.ZN( u2_out5_16 ) , .A4( u2_u5_u2_n128 ) , .A3( u2_u5_u2_n129 ) , .A1( u2_u5_u2_n130 ) , .A2( u2_u5_u2_n186 ) );
  AOI22_X1 u2_u5_u2_U89 (.A2( u2_u5_u2_n118 ) , .ZN( u2_u5_u2_n129 ) , .A1( u2_u5_u2_n140 ) , .B1( u2_u5_u2_n157 ) , .B2( u2_u5_u2_n170 ) );
  AOI21_X1 u2_u5_u2_U9 (.B2( u2_u5_u2_n123 ) , .ZN( u2_u5_u2_n125 ) , .A( u2_u5_u2_n171 ) , .B1( u2_u5_u2_n184 ) );
  INV_X1 u2_u5_u2_U90 (.A( u2_u5_u2_n163 ) , .ZN( u2_u5_u2_n186 ) );
  NAND4_X1 u2_u5_u2_U91 (.ZN( u2_out5_30 ) , .A4( u2_u5_u2_n147 ) , .A3( u2_u5_u2_n148 ) , .A2( u2_u5_u2_n149 ) , .A1( u2_u5_u2_n187 ) );
  NOR3_X1 u2_u5_u2_U92 (.A3( u2_u5_u2_n144 ) , .A2( u2_u5_u2_n145 ) , .A1( u2_u5_u2_n146 ) , .ZN( u2_u5_u2_n147 ) );
  AOI21_X1 u2_u5_u2_U93 (.B2( u2_u5_u2_n138 ) , .ZN( u2_u5_u2_n148 ) , .A( u2_u5_u2_n162 ) , .B1( u2_u5_u2_n182 ) );
  OR4_X1 u2_u5_u2_U94 (.ZN( u2_out5_6 ) , .A4( u2_u5_u2_n161 ) , .A3( u2_u5_u2_n162 ) , .A2( u2_u5_u2_n163 ) , .A1( u2_u5_u2_n164 ) );
  OR3_X1 u2_u5_u2_U95 (.A2( u2_u5_u2_n159 ) , .A1( u2_u5_u2_n160 ) , .ZN( u2_u5_u2_n161 ) , .A3( u2_u5_u2_n183 ) );
  AOI21_X1 u2_u5_u2_U96 (.B2( u2_u5_u2_n154 ) , .B1( u2_u5_u2_n155 ) , .ZN( u2_u5_u2_n159 ) , .A( u2_u5_u2_n167 ) );
  NAND3_X1 u2_u5_u2_U97 (.A2( u2_u5_u2_n117 ) , .A1( u2_u5_u2_n122 ) , .A3( u2_u5_u2_n123 ) , .ZN( u2_u5_u2_n134 ) );
  NAND3_X1 u2_u5_u2_U98 (.ZN( u2_u5_u2_n110 ) , .A2( u2_u5_u2_n131 ) , .A3( u2_u5_u2_n139 ) , .A1( u2_u5_u2_n154 ) );
  NAND3_X1 u2_u5_u2_U99 (.A2( u2_u5_u2_n100 ) , .ZN( u2_u5_u2_n101 ) , .A1( u2_u5_u2_n104 ) , .A3( u2_u5_u2_n114 ) );
  XOR2_X1 u2_u7_U16 (.B( u2_K8_3 ) , .A( u2_R6_2 ) , .Z( u2_u7_X_3 ) );
  XOR2_X1 u2_u7_U27 (.B( u2_K8_2 ) , .A( u2_R6_1 ) , .Z( u2_u7_X_2 ) );
  XOR2_X1 u2_u7_U38 (.B( u2_K8_1 ) , .A( u2_R6_32 ) , .Z( u2_u7_X_1 ) );
  XOR2_X1 u2_u7_U4 (.B( u2_K8_6 ) , .A( u2_R6_5 ) , .Z( u2_u7_X_6 ) );
  XOR2_X1 u2_u7_U5 (.B( u2_K8_5 ) , .A( u2_R6_4 ) , .Z( u2_u7_X_5 ) );
  XOR2_X1 u2_u7_U6 (.B( u2_K8_4 ) , .A( u2_R6_3 ) , .Z( u2_u7_X_4 ) );
  AND3_X1 u2_u7_u0_U10 (.A2( u2_u7_u0_n112 ) , .ZN( u2_u7_u0_n127 ) , .A3( u2_u7_u0_n130 ) , .A1( u2_u7_u0_n148 ) );
  NAND2_X1 u2_u7_u0_U11 (.ZN( u2_u7_u0_n113 ) , .A1( u2_u7_u0_n139 ) , .A2( u2_u7_u0_n149 ) );
  AND2_X1 u2_u7_u0_U12 (.ZN( u2_u7_u0_n107 ) , .A1( u2_u7_u0_n130 ) , .A2( u2_u7_u0_n140 ) );
  AND2_X1 u2_u7_u0_U13 (.A2( u2_u7_u0_n129 ) , .A1( u2_u7_u0_n130 ) , .ZN( u2_u7_u0_n151 ) );
  AND2_X1 u2_u7_u0_U14 (.A1( u2_u7_u0_n108 ) , .A2( u2_u7_u0_n125 ) , .ZN( u2_u7_u0_n145 ) );
  INV_X1 u2_u7_u0_U15 (.A( u2_u7_u0_n143 ) , .ZN( u2_u7_u0_n173 ) );
  NOR2_X1 u2_u7_u0_U16 (.A2( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n147 ) , .A1( u2_u7_u0_n160 ) );
  INV_X1 u2_u7_u0_U17 (.ZN( u2_u7_u0_n172 ) , .A( u2_u7_u0_n88 ) );
  OAI222_X1 u2_u7_u0_U18 (.C1( u2_u7_u0_n108 ) , .A1( u2_u7_u0_n125 ) , .B2( u2_u7_u0_n128 ) , .B1( u2_u7_u0_n144 ) , .A2( u2_u7_u0_n158 ) , .C2( u2_u7_u0_n161 ) , .ZN( u2_u7_u0_n88 ) );
  NOR2_X1 u2_u7_u0_U19 (.A1( u2_u7_u0_n163 ) , .A2( u2_u7_u0_n164 ) , .ZN( u2_u7_u0_n95 ) );
  OAI22_X1 u2_u7_u0_U20 (.B1( u2_u7_u0_n125 ) , .ZN( u2_u7_u0_n126 ) , .A1( u2_u7_u0_n138 ) , .A2( u2_u7_u0_n146 ) , .B2( u2_u7_u0_n147 ) );
  OAI22_X1 u2_u7_u0_U21 (.B1( u2_u7_u0_n131 ) , .A1( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n147 ) , .A2( u2_u7_u0_n90 ) , .ZN( u2_u7_u0_n91 ) );
  AND3_X1 u2_u7_u0_U22 (.A3( u2_u7_u0_n121 ) , .A2( u2_u7_u0_n125 ) , .A1( u2_u7_u0_n148 ) , .ZN( u2_u7_u0_n90 ) );
  INV_X1 u2_u7_u0_U23 (.A( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n161 ) );
  AOI22_X1 u2_u7_u0_U24 (.B2( u2_u7_u0_n109 ) , .A2( u2_u7_u0_n110 ) , .ZN( u2_u7_u0_n111 ) , .B1( u2_u7_u0_n118 ) , .A1( u2_u7_u0_n160 ) );
  INV_X1 u2_u7_u0_U25 (.A( u2_u7_u0_n118 ) , .ZN( u2_u7_u0_n158 ) );
  AOI21_X1 u2_u7_u0_U26 (.ZN( u2_u7_u0_n104 ) , .B1( u2_u7_u0_n107 ) , .B2( u2_u7_u0_n141 ) , .A( u2_u7_u0_n144 ) );
  AOI21_X1 u2_u7_u0_U27 (.B1( u2_u7_u0_n127 ) , .B2( u2_u7_u0_n129 ) , .A( u2_u7_u0_n138 ) , .ZN( u2_u7_u0_n96 ) );
  AOI21_X1 u2_u7_u0_U28 (.ZN( u2_u7_u0_n116 ) , .B2( u2_u7_u0_n142 ) , .A( u2_u7_u0_n144 ) , .B1( u2_u7_u0_n166 ) );
  INV_X1 u2_u7_u0_U29 (.ZN( u2_u7_u0_n171 ) , .A( u2_u7_u0_n99 ) );
  INV_X1 u2_u7_u0_U3 (.A( u2_u7_u0_n113 ) , .ZN( u2_u7_u0_n166 ) );
  OAI211_X1 u2_u7_u0_U30 (.C2( u2_u7_u0_n140 ) , .C1( u2_u7_u0_n161 ) , .A( u2_u7_u0_n169 ) , .B( u2_u7_u0_n98 ) , .ZN( u2_u7_u0_n99 ) );
  INV_X1 u2_u7_u0_U31 (.ZN( u2_u7_u0_n169 ) , .A( u2_u7_u0_n91 ) );
  AOI211_X1 u2_u7_u0_U32 (.C1( u2_u7_u0_n118 ) , .A( u2_u7_u0_n123 ) , .B( u2_u7_u0_n96 ) , .C2( u2_u7_u0_n97 ) , .ZN( u2_u7_u0_n98 ) );
  NOR2_X1 u2_u7_u0_U33 (.A1( u2_u7_u0_n120 ) , .ZN( u2_u7_u0_n143 ) , .A2( u2_u7_u0_n167 ) );
  OAI221_X1 u2_u7_u0_U34 (.C1( u2_u7_u0_n112 ) , .ZN( u2_u7_u0_n120 ) , .B1( u2_u7_u0_n138 ) , .B2( u2_u7_u0_n141 ) , .C2( u2_u7_u0_n147 ) , .A( u2_u7_u0_n172 ) );
  AOI211_X1 u2_u7_u0_U35 (.B( u2_u7_u0_n115 ) , .A( u2_u7_u0_n116 ) , .C2( u2_u7_u0_n117 ) , .C1( u2_u7_u0_n118 ) , .ZN( u2_u7_u0_n119 ) );
  NAND2_X1 u2_u7_u0_U36 (.A1( u2_u7_u0_n101 ) , .A2( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n150 ) );
  INV_X1 u2_u7_u0_U37 (.A( u2_u7_u0_n138 ) , .ZN( u2_u7_u0_n160 ) );
  NAND2_X1 u2_u7_u0_U38 (.A1( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n128 ) , .A2( u2_u7_u0_n95 ) );
  NAND2_X1 u2_u7_u0_U39 (.ZN( u2_u7_u0_n148 ) , .A1( u2_u7_u0_n93 ) , .A2( u2_u7_u0_n95 ) );
  AOI21_X1 u2_u7_u0_U4 (.B1( u2_u7_u0_n114 ) , .ZN( u2_u7_u0_n115 ) , .B2( u2_u7_u0_n129 ) , .A( u2_u7_u0_n161 ) );
  NAND2_X1 u2_u7_u0_U40 (.A2( u2_u7_u0_n102 ) , .A1( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n149 ) );
  NAND2_X1 u2_u7_u0_U41 (.A2( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n114 ) , .A1( u2_u7_u0_n92 ) );
  NAND2_X1 u2_u7_u0_U42 (.A2( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n121 ) , .A1( u2_u7_u0_n93 ) );
  NAND2_X1 u2_u7_u0_U43 (.ZN( u2_u7_u0_n112 ) , .A2( u2_u7_u0_n92 ) , .A1( u2_u7_u0_n93 ) );
  AOI21_X1 u2_u7_u0_U44 (.B1( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n132 ) , .A( u2_u7_u0_n165 ) , .B2( u2_u7_u0_n93 ) );
  INV_X1 u2_u7_u0_U45 (.A( u2_u7_u0_n142 ) , .ZN( u2_u7_u0_n165 ) );
  OR3_X1 u2_u7_u0_U46 (.A3( u2_u7_u0_n152 ) , .A2( u2_u7_u0_n153 ) , .A1( u2_u7_u0_n154 ) , .ZN( u2_u7_u0_n155 ) );
  AOI21_X1 u2_u7_u0_U47 (.A( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n145 ) , .B1( u2_u7_u0_n146 ) , .ZN( u2_u7_u0_n154 ) );
  AOI21_X1 u2_u7_u0_U48 (.B2( u2_u7_u0_n150 ) , .B1( u2_u7_u0_n151 ) , .ZN( u2_u7_u0_n152 ) , .A( u2_u7_u0_n158 ) );
  AOI21_X1 u2_u7_u0_U49 (.A( u2_u7_u0_n147 ) , .B2( u2_u7_u0_n148 ) , .B1( u2_u7_u0_n149 ) , .ZN( u2_u7_u0_n153 ) );
  AOI21_X1 u2_u7_u0_U5 (.B2( u2_u7_u0_n131 ) , .ZN( u2_u7_u0_n134 ) , .B1( u2_u7_u0_n151 ) , .A( u2_u7_u0_n158 ) );
  NOR2_X1 u2_u7_u0_U50 (.A2( u2_u7_X_4 ) , .A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n118 ) );
  NAND2_X1 u2_u7_u0_U51 (.A2( u2_u7_X_4 ) , .A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n144 ) );
  NOR2_X1 u2_u7_u0_U52 (.A2( u2_u7_X_1 ) , .A1( u2_u7_X_2 ) , .ZN( u2_u7_u0_n92 ) );
  NOR2_X1 u2_u7_u0_U53 (.A2( u2_u7_X_1 ) , .ZN( u2_u7_u0_n101 ) , .A1( u2_u7_u0_n163 ) );
  NOR2_X1 u2_u7_u0_U54 (.A2( u2_u7_X_2 ) , .ZN( u2_u7_u0_n103 ) , .A1( u2_u7_u0_n164 ) );
  NOR2_X1 u2_u7_u0_U55 (.A2( u2_u7_X_5 ) , .ZN( u2_u7_u0_n136 ) , .A1( u2_u7_u0_n159 ) );
  NAND2_X1 u2_u7_u0_U56 (.A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n138 ) , .A2( u2_u7_u0_n159 ) );
  AND2_X1 u2_u7_u0_U57 (.A2( u2_u7_X_3 ) , .A1( u2_u7_X_6 ) , .ZN( u2_u7_u0_n102 ) );
  AND2_X1 u2_u7_u0_U58 (.A1( u2_u7_X_6 ) , .A2( u2_u7_u0_n162 ) , .ZN( u2_u7_u0_n93 ) );
  INV_X1 u2_u7_u0_U59 (.A( u2_u7_X_4 ) , .ZN( u2_u7_u0_n159 ) );
  NOR2_X1 u2_u7_u0_U6 (.A1( u2_u7_u0_n108 ) , .ZN( u2_u7_u0_n123 ) , .A2( u2_u7_u0_n158 ) );
  INV_X1 u2_u7_u0_U60 (.A( u2_u7_X_1 ) , .ZN( u2_u7_u0_n164 ) );
  INV_X1 u2_u7_u0_U61 (.A( u2_u7_X_2 ) , .ZN( u2_u7_u0_n163 ) );
  INV_X1 u2_u7_u0_U62 (.A( u2_u7_u0_n126 ) , .ZN( u2_u7_u0_n168 ) );
  AOI211_X1 u2_u7_u0_U63 (.B( u2_u7_u0_n133 ) , .A( u2_u7_u0_n134 ) , .C2( u2_u7_u0_n135 ) , .C1( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n137 ) );
  OR4_X1 u2_u7_u0_U64 (.ZN( u2_out7_17 ) , .A4( u2_u7_u0_n122 ) , .A2( u2_u7_u0_n123 ) , .A1( u2_u7_u0_n124 ) , .A3( u2_u7_u0_n170 ) );
  AOI21_X1 u2_u7_u0_U65 (.B2( u2_u7_u0_n107 ) , .ZN( u2_u7_u0_n124 ) , .B1( u2_u7_u0_n128 ) , .A( u2_u7_u0_n161 ) );
  INV_X1 u2_u7_u0_U66 (.A( u2_u7_u0_n111 ) , .ZN( u2_u7_u0_n170 ) );
  OR4_X1 u2_u7_u0_U67 (.ZN( u2_out7_31 ) , .A4( u2_u7_u0_n155 ) , .A2( u2_u7_u0_n156 ) , .A1( u2_u7_u0_n157 ) , .A3( u2_u7_u0_n173 ) );
  AOI21_X1 u2_u7_u0_U68 (.A( u2_u7_u0_n138 ) , .B2( u2_u7_u0_n139 ) , .B1( u2_u7_u0_n140 ) , .ZN( u2_u7_u0_n157 ) );
  AOI21_X1 u2_u7_u0_U69 (.B2( u2_u7_u0_n141 ) , .B1( u2_u7_u0_n142 ) , .ZN( u2_u7_u0_n156 ) , .A( u2_u7_u0_n161 ) );
  OAI21_X1 u2_u7_u0_U7 (.B1( u2_u7_u0_n150 ) , .B2( u2_u7_u0_n158 ) , .A( u2_u7_u0_n172 ) , .ZN( u2_u7_u0_n89 ) );
  INV_X1 u2_u7_u0_U70 (.ZN( u2_u7_u0_n174 ) , .A( u2_u7_u0_n89 ) );
  AOI211_X1 u2_u7_u0_U71 (.B( u2_u7_u0_n104 ) , .A( u2_u7_u0_n105 ) , .ZN( u2_u7_u0_n106 ) , .C2( u2_u7_u0_n113 ) , .C1( u2_u7_u0_n160 ) );
  NAND2_X1 u2_u7_u0_U72 (.A2( u2_u7_u0_n100 ) , .A1( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n139 ) );
  NAND2_X1 u2_u7_u0_U73 (.A1( u2_u7_u0_n100 ) , .A2( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n125 ) );
  NAND2_X1 u2_u7_u0_U74 (.A1( u2_u7_u0_n100 ) , .ZN( u2_u7_u0_n129 ) , .A2( u2_u7_u0_n95 ) );
  NAND2_X1 u2_u7_u0_U75 (.A2( u2_u7_u0_n100 ) , .ZN( u2_u7_u0_n131 ) , .A1( u2_u7_u0_n92 ) );
  OAI221_X1 u2_u7_u0_U76 (.C1( u2_u7_u0_n121 ) , .ZN( u2_u7_u0_n122 ) , .B2( u2_u7_u0_n127 ) , .A( u2_u7_u0_n143 ) , .B1( u2_u7_u0_n144 ) , .C2( u2_u7_u0_n147 ) );
  NOR2_X1 u2_u7_u0_U77 (.A2( u2_u7_X_6 ) , .ZN( u2_u7_u0_n100 ) , .A1( u2_u7_u0_n162 ) );
  AOI21_X1 u2_u7_u0_U78 (.B1( u2_u7_u0_n132 ) , .ZN( u2_u7_u0_n133 ) , .A( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n166 ) );
  OAI22_X1 u2_u7_u0_U79 (.ZN( u2_u7_u0_n105 ) , .A2( u2_u7_u0_n132 ) , .B1( u2_u7_u0_n146 ) , .A1( u2_u7_u0_n147 ) , .B2( u2_u7_u0_n161 ) );
  AND2_X1 u2_u7_u0_U8 (.A1( u2_u7_u0_n114 ) , .A2( u2_u7_u0_n121 ) , .ZN( u2_u7_u0_n146 ) );
  NAND2_X1 u2_u7_u0_U80 (.ZN( u2_u7_u0_n110 ) , .A2( u2_u7_u0_n132 ) , .A1( u2_u7_u0_n145 ) );
  INV_X1 u2_u7_u0_U81 (.A( u2_u7_u0_n119 ) , .ZN( u2_u7_u0_n167 ) );
  NAND2_X1 u2_u7_u0_U82 (.A2( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n140 ) , .A1( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U83 (.A1( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n130 ) , .A2( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U84 (.ZN( u2_u7_u0_n108 ) , .A1( u2_u7_u0_n92 ) , .A2( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U85 (.ZN( u2_u7_u0_n142 ) , .A1( u2_u7_u0_n94 ) , .A2( u2_u7_u0_n95 ) );
  INV_X1 u2_u7_u0_U86 (.A( u2_u7_X_3 ) , .ZN( u2_u7_u0_n162 ) );
  NOR2_X1 u2_u7_u0_U87 (.A2( u2_u7_X_3 ) , .A1( u2_u7_X_6 ) , .ZN( u2_u7_u0_n94 ) );
  NAND3_X1 u2_u7_u0_U88 (.ZN( u2_out7_23 ) , .A3( u2_u7_u0_n137 ) , .A1( u2_u7_u0_n168 ) , .A2( u2_u7_u0_n171 ) );
  NAND3_X1 u2_u7_u0_U89 (.A3( u2_u7_u0_n127 ) , .A2( u2_u7_u0_n128 ) , .ZN( u2_u7_u0_n135 ) , .A1( u2_u7_u0_n150 ) );
  AND2_X1 u2_u7_u0_U9 (.A1( u2_u7_u0_n131 ) , .ZN( u2_u7_u0_n141 ) , .A2( u2_u7_u0_n150 ) );
  NAND3_X1 u2_u7_u0_U90 (.ZN( u2_u7_u0_n117 ) , .A3( u2_u7_u0_n132 ) , .A2( u2_u7_u0_n139 ) , .A1( u2_u7_u0_n148 ) );
  NAND3_X1 u2_u7_u0_U91 (.ZN( u2_u7_u0_n109 ) , .A2( u2_u7_u0_n114 ) , .A3( u2_u7_u0_n140 ) , .A1( u2_u7_u0_n149 ) );
  NAND3_X1 u2_u7_u0_U92 (.ZN( u2_out7_9 ) , .A3( u2_u7_u0_n106 ) , .A2( u2_u7_u0_n171 ) , .A1( u2_u7_u0_n174 ) );
  NAND3_X1 u2_u7_u0_U93 (.A2( u2_u7_u0_n128 ) , .A1( u2_u7_u0_n132 ) , .A3( u2_u7_u0_n146 ) , .ZN( u2_u7_u0_n97 ) );
  INV_X1 u2_uk_U1088 (.ZN( u2_K8_3 ) , .A( u2_uk_n1110 ) );
  AOI22_X1 u2_uk_U1089 (.B2( u2_uk_K_r6_10 ) , .A2( u2_uk_K_r6_3 ) , .ZN( u2_uk_n1110 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n162 ) );
  OAI21_X1 u2_uk_U499 (.ZN( u2_K8_2 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1105 ) , .B2( u2_uk_n1515 ) );
  INV_X1 u2_uk_U546 (.ZN( u2_K6_17 ) , .A( u2_uk_n1059 ) );
  AOI22_X1 u2_uk_U547 (.B2( u2_uk_K_r4_4 ) , .A2( u2_uk_K_r4_55 ) , .ZN( u2_uk_n1059 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n147 ) );
  INV_X1 u2_uk_U822 (.ZN( u2_K6_18 ) , .A( u2_uk_n1060 ) );
  AOI22_X1 u2_uk_U823 (.B2( u2_uk_K_r4_11 ) , .A2( u2_uk_K_r4_17 ) , .A1( u2_uk_n100 ) , .ZN( u2_uk_n1060 ) , .B1( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U828 (.ZN( u2_K8_6 ) , .B2( u2_uk_n1514 ) , .A2( u2_uk_n1519 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U870 (.ZN( u2_K8_1 ) , .A2( u2_uk_n1502 ) , .B2( u2_uk_n1518 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n27 ) );
  OAI21_X1 u2_uk_U989 (.ZN( u2_K8_4 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1116 ) , .B2( u2_uk_n1507 ) );
endmodule

