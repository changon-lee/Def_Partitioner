module des_des_die_4 ( u0_L13_11, u0_L13_19, u0_L13_29, u0_L13_4, u0_L1_12, u0_L1_15, u0_L1_21, u0_L1_22, u0_L1_27, 
       u0_L1_32, u0_L1_5, u0_L1_7, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, 
       u0_R1_1, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_30, u0_R1_31, 
       u0_R1_32, u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_22, u0_uk_K_r5_13, u0_uk_n110, u0_uk_n118, u0_uk_n128, 
       u0_uk_n13, u0_uk_n148, u0_uk_n155, u0_uk_n164, u0_uk_n18, u0_uk_n187, u0_uk_n202, u0_uk_n208, u0_uk_n209, 
       u0_uk_n230, u0_uk_n27, u0_uk_n28, u0_uk_n31, u0_uk_n32, u0_uk_n33, u0_uk_n4, u0_uk_n45, u0_uk_n546, 
       u0_uk_n550, u0_uk_n553, u0_uk_n554, u0_uk_n558, u0_uk_n560, u0_uk_n561, u0_uk_n566, u0_uk_n570, u0_uk_n574, 
       u0_uk_n575, u0_uk_n581, u0_uk_n83, u0_uk_n917, u0_uk_n918, u0_uk_n92, u1_FP_33, u1_FP_34, u1_FP_35, 
       u1_FP_36, u1_FP_37, u1_FP_38, u1_FP_39, u1_FP_40, u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_46, 
       u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_64, u1_L10_11, u1_L10_12, u1_L10_15, u1_L10_19, u1_L10_21, 
       u1_L10_22, u1_L10_27, u1_L10_29, u1_L10_32, u1_L10_4, u1_L10_5, u1_L10_7, u1_L12_13, u1_L12_16, 
       u1_L12_17, u1_L12_18, u1_L12_2, u1_L12_23, u1_L12_24, u1_L12_28, u1_L12_30, u1_L12_31, u1_L12_6, 
       u1_L12_9, u1_L14_1, u1_L14_10, u1_L14_13, u1_L14_17, u1_L14_18, u1_L14_2, u1_L14_20, u1_L14_23, 
       u1_L14_26, u1_L14_28, u1_L14_31, u1_L14_9, u1_L2_1, u1_L2_10, u1_L2_15, u1_L2_16, u1_L2_17, 
       u1_L2_20, u1_L2_21, u1_L2_23, u1_L2_24, u1_L2_26, u1_L2_27, u1_L2_30, u1_L2_31, u1_L2_5, 
       u1_L2_6, u1_L2_9, u1_L6_15, u1_L6_21, u1_L6_27, u1_L6_5, u1_L8_11, u1_L8_12, u1_L8_19, 
       u1_L8_22, u1_L8_29, u1_L8_32, u1_L8_4, u1_L8_7, u1_R10_1, u1_R10_20, u1_R10_21, u1_R10_22, 
       u1_R10_23, u1_R10_24, u1_R10_25, u1_R10_26, u1_R10_27, u1_R10_28, u1_R10_29, u1_R10_30, u1_R10_31, 
       u1_R10_32, u1_R12_1, u1_R12_10, u1_R12_11, u1_R12_12, u1_R12_13, u1_R12_2, u1_R12_3, u1_R12_32, 
       u1_R12_4, u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R2_1, u1_R2_10, u1_R2_11, 
       u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_2, u1_R2_28, u1_R2_29, 
       u1_R2_3, u1_R2_30, u1_R2_31, u1_R2_32, u1_R2_4, u1_R2_5, u1_R2_8, u1_R2_9, u1_R6_1, 
       u1_R6_28, u1_R6_29, u1_R6_30, u1_R6_31, u1_R6_32, u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_23, 
       u1_R8_24, u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_23, 
       u1_uk_K_r10_28, u1_uk_K_r10_37, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r12_10, 
       u1_uk_K_r12_18, u1_uk_K_r12_47, u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_3, u1_uk_K_r14_39, u1_uk_K_r2_13, u1_uk_K_r2_18, u1_uk_K_r2_20, 
       u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_29, u1_uk_K_r2_33, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, 
       u1_uk_K_r2_47, u1_uk_K_r2_53, u1_uk_K_r2_55, u1_uk_K_r6_0, u1_uk_K_r6_21, u1_uk_K_r6_28, u1_uk_K_r6_37, u1_uk_K_r8_16, u1_uk_K_r8_2, 
       u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_28, u1_uk_K_r8_37, u1_uk_K_r8_42, u1_uk_K_r8_44, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, 
       u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n110, u1_uk_n118, u1_uk_n1220, u1_uk_n1221, 
       u1_uk_n1224, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1242, 
       u1_uk_n1243, u1_uk_n1244, u1_uk_n1248, u1_uk_n1249, u1_uk_n1251, u1_uk_n1252, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, 
       u1_uk_n128, u1_uk_n129, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1357, 
       u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1363, u1_uk_n1365, u1_uk_n1367, u1_uk_n1369, u1_uk_n1371, u1_uk_n1374, 
       u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1393, u1_uk_n141, 
       u1_uk_n142, u1_uk_n145, u1_uk_n146, u1_uk_n147, u1_uk_n1528, u1_uk_n1534, u1_uk_n1541, u1_uk_n155, u1_uk_n1561, 
       u1_uk_n1562, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n161, u1_uk_n1618, u1_uk_n1619, u1_uk_n162, u1_uk_n1624, 
       u1_uk_n163, u1_uk_n1644, u1_uk_n1645, u1_uk_n1652, u1_uk_n17, u1_uk_n1708, u1_uk_n1709, u1_uk_n1714, u1_uk_n1715, 
       u1_uk_n1717, u1_uk_n1720, u1_uk_n1721, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, 
       u1_uk_n1744, u1_uk_n1748, u1_uk_n1749, u1_uk_n1801, u1_uk_n1803, u1_uk_n1804, u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, 
       u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n182, u1_uk_n1824, 
       u1_uk_n1826, u1_uk_n1831, u1_uk_n1834, u1_uk_n1835, u1_uk_n1841, u1_uk_n1842, u1_uk_n187, u1_uk_n188, u1_uk_n191, 
       u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, u1_uk_n209, u1_uk_n213, u1_uk_n214, u1_uk_n217, u1_uk_n220, 
       u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, 
       u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, 
       u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n63, u1_uk_n94, u1_uk_n99, u2_FP_52, u2_FP_53, 
       u2_FP_54, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_K16_31, 
       u2_K16_42, u2_K7_26, u2_K7_31, u2_K7_33, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_45, 
       u2_K7_48, u2_L14_11, u2_L14_12, u2_L14_19, u2_L14_22, u2_L14_29, u2_L14_32, u2_L14_4, u2_L14_7, 
       u2_L5_11, u2_L5_12, u2_L5_14, u2_L5_15, u2_L5_19, u2_L5_21, u2_L5_22, u2_L5_25, u2_L5_27, 
       u2_L5_29, u2_L5_3, u2_L5_32, u2_L5_4, u2_L5_5, u2_L5_7, u2_L5_8, u2_R5_1, u2_R5_16, 
       u2_R5_17, u2_R5_18, u2_R5_19, u2_R5_20, u2_R5_21, u2_R5_22, u2_R5_23, u2_R5_24, u2_R5_25, 
       u2_R5_26, u2_R5_27, u2_R5_28, u2_R5_29, u2_R5_30, u2_R5_31, u2_R5_32, u2_key_r_50, u2_uk_K_r14_15, 
       u2_uk_K_r14_2, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_21, u2_uk_K_r5_23, u2_uk_K_r5_31, u2_uk_K_r5_43, 
       u2_uk_K_r5_51, u2_uk_K_r5_7, u2_uk_n10, u2_uk_n1089, u2_uk_n1093, u2_uk_n1094, u2_uk_n11, u2_uk_n117, u2_uk_n118, 
       u2_uk_n1188, u2_uk_n1201, u2_uk_n1203, u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1215, u2_uk_n1217, u2_uk_n1220, 
       u2_uk_n1225, u2_uk_n1226, u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n1452, u2_uk_n1456, u2_uk_n1459, 
       u2_uk_n1460, u2_uk_n1464, u2_uk_n147, u2_uk_n1470, u2_uk_n1471, u2_uk_n1480, u2_uk_n1486, u2_uk_n1490, u2_uk_n1491, 
       u2_uk_n1493, u2_uk_n161, u2_uk_n164, u2_uk_n182, u2_uk_n202, u2_uk_n208, u2_uk_n213, u2_uk_n217, u2_uk_n223, 
       u2_uk_n231, u2_uk_n238, u2_uk_n94, u2_uk_n961, u0_N451, u0_N458, u0_N466, u0_N476, u0_N68, u0_N70, u0_N75, u0_N78, u0_N84, 
        u0_N85, u0_N90, u0_N95, u0_uk_n191, u0_uk_n63, u0_uk_n777, u1_FP_1, u1_FP_10, u1_FP_13, 
        u1_FP_17, u1_FP_18, u1_FP_2, u1_FP_20, u1_FP_23, u1_FP_26, u1_FP_28, u1_FP_31, u1_FP_9, 
        u1_N100, u1_N101, u1_N104, u1_N105, u1_N110, u1_N111, u1_N112, u1_N115, u1_N116, 
        u1_N118, u1_N119, u1_N121, u1_N122, u1_N125, u1_N126, u1_N228, u1_N238, u1_N244, 
        u1_N250, u1_N291, u1_N294, u1_N298, u1_N299, u1_N306, u1_N309, u1_N316, u1_N319, 
        u1_N355, u1_N356, u1_N358, u1_N362, u1_N363, u1_N366, u1_N370, u1_N372, u1_N373, 
        u1_N378, u1_N380, u1_N383, u1_N417, u1_N421, u1_N424, u1_N428, u1_N431, u1_N432, 
        u1_N433, u1_N438, u1_N439, u1_N443, u1_N445, u1_N446, u1_N96, u1_uk_n117, u1_uk_n83, 
        u2_FP_11, u2_FP_12, u2_FP_19, u2_FP_22, u2_FP_29, u2_FP_32, u2_FP_4, u2_FP_7, u2_N194, 
        u2_N195, u2_N196, u2_N198, u2_N199, u2_N202, u2_N203, u2_N205, u2_N206, u2_N210, 
        u2_N212, u2_N213, u2_N216, u2_N218, u2_N220, u2_N223, u2_uk_n31, u2_uk_n983 );
  input u0_L13_11, u0_L13_19, u0_L13_29, u0_L13_4, u0_L1_12, u0_L1_15, u0_L1_21, u0_L1_22, u0_L1_27, 
        u0_L1_32, u0_L1_5, u0_L1_7, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, u0_R13_24, u0_R13_25, 
        u0_R1_1, u0_R1_24, u0_R1_25, u0_R1_26, u0_R1_27, u0_R1_28, u0_R1_29, u0_R1_30, u0_R1_31, 
        u0_R1_32, u0_uk_K_r1_15, u0_uk_K_r1_16, u0_uk_K_r1_21, u0_uk_K_r1_22, u0_uk_K_r5_13, u0_uk_n110, u0_uk_n118, u0_uk_n128, 
        u0_uk_n13, u0_uk_n148, u0_uk_n155, u0_uk_n164, u0_uk_n18, u0_uk_n187, u0_uk_n202, u0_uk_n208, u0_uk_n209, 
        u0_uk_n230, u0_uk_n27, u0_uk_n28, u0_uk_n31, u0_uk_n32, u0_uk_n33, u0_uk_n4, u0_uk_n45, u0_uk_n546, 
        u0_uk_n550, u0_uk_n553, u0_uk_n554, u0_uk_n558, u0_uk_n560, u0_uk_n561, u0_uk_n566, u0_uk_n570, u0_uk_n574, 
        u0_uk_n575, u0_uk_n581, u0_uk_n83, u0_uk_n917, u0_uk_n918, u0_uk_n92, u1_FP_33, u1_FP_34, u1_FP_35, 
        u1_FP_36, u1_FP_37, u1_FP_38, u1_FP_39, u1_FP_40, u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_46, 
        u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_64, u1_L10_11, u1_L10_12, u1_L10_15, u1_L10_19, u1_L10_21, 
        u1_L10_22, u1_L10_27, u1_L10_29, u1_L10_32, u1_L10_4, u1_L10_5, u1_L10_7, u1_L12_13, u1_L12_16, 
        u1_L12_17, u1_L12_18, u1_L12_2, u1_L12_23, u1_L12_24, u1_L12_28, u1_L12_30, u1_L12_31, u1_L12_6, 
        u1_L12_9, u1_L14_1, u1_L14_10, u1_L14_13, u1_L14_17, u1_L14_18, u1_L14_2, u1_L14_20, u1_L14_23, 
        u1_L14_26, u1_L14_28, u1_L14_31, u1_L14_9, u1_L2_1, u1_L2_10, u1_L2_15, u1_L2_16, u1_L2_17, 
        u1_L2_20, u1_L2_21, u1_L2_23, u1_L2_24, u1_L2_26, u1_L2_27, u1_L2_30, u1_L2_31, u1_L2_5, 
        u1_L2_6, u1_L2_9, u1_L6_15, u1_L6_21, u1_L6_27, u1_L6_5, u1_L8_11, u1_L8_12, u1_L8_19, 
        u1_L8_22, u1_L8_29, u1_L8_32, u1_L8_4, u1_L8_7, u1_R10_1, u1_R10_20, u1_R10_21, u1_R10_22, 
        u1_R10_23, u1_R10_24, u1_R10_25, u1_R10_26, u1_R10_27, u1_R10_28, u1_R10_29, u1_R10_30, u1_R10_31, 
        u1_R10_32, u1_R12_1, u1_R12_10, u1_R12_11, u1_R12_12, u1_R12_13, u1_R12_2, u1_R12_3, u1_R12_32, 
        u1_R12_4, u1_R12_5, u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R2_1, u1_R2_10, u1_R2_11, 
        u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, u1_R2_17, u1_R2_2, u1_R2_28, u1_R2_29, 
        u1_R2_3, u1_R2_30, u1_R2_31, u1_R2_32, u1_R2_4, u1_R2_5, u1_R2_8, u1_R2_9, u1_R6_1, 
        u1_R6_28, u1_R6_29, u1_R6_30, u1_R6_31, u1_R6_32, u1_R8_20, u1_R8_21, u1_R8_22, u1_R8_23, 
        u1_R8_24, u1_R8_25, u1_R8_26, u1_R8_27, u1_R8_28, u1_R8_29, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_23, 
        u1_uk_K_r10_28, u1_uk_K_r10_37, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r12_10, 
        u1_uk_K_r12_18, u1_uk_K_r12_47, u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_3, u1_uk_K_r14_39, u1_uk_K_r2_13, u1_uk_K_r2_18, u1_uk_K_r2_20, 
        u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_29, u1_uk_K_r2_33, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, 
        u1_uk_K_r2_47, u1_uk_K_r2_53, u1_uk_K_r2_55, u1_uk_K_r6_0, u1_uk_K_r6_21, u1_uk_K_r6_28, u1_uk_K_r6_37, u1_uk_K_r8_16, u1_uk_K_r8_2, 
        u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_28, u1_uk_K_r8_37, u1_uk_K_r8_42, u1_uk_K_r8_44, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, 
        u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n110, u1_uk_n118, u1_uk_n1220, u1_uk_n1221, 
        u1_uk_n1224, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1242, 
        u1_uk_n1243, u1_uk_n1244, u1_uk_n1248, u1_uk_n1249, u1_uk_n1251, u1_uk_n1252, u1_uk_n1257, u1_uk_n1258, u1_uk_n1259, 
        u1_uk_n128, u1_uk_n129, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1357, 
        u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1363, u1_uk_n1365, u1_uk_n1367, u1_uk_n1369, u1_uk_n1371, u1_uk_n1374, 
        u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1393, u1_uk_n141, 
        u1_uk_n142, u1_uk_n145, u1_uk_n146, u1_uk_n147, u1_uk_n1528, u1_uk_n1534, u1_uk_n1541, u1_uk_n155, u1_uk_n1561, 
        u1_uk_n1562, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n161, u1_uk_n1618, u1_uk_n1619, u1_uk_n162, u1_uk_n1624, 
        u1_uk_n163, u1_uk_n1644, u1_uk_n1645, u1_uk_n1652, u1_uk_n17, u1_uk_n1708, u1_uk_n1709, u1_uk_n1714, u1_uk_n1715, 
        u1_uk_n1717, u1_uk_n1720, u1_uk_n1721, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, 
        u1_uk_n1744, u1_uk_n1748, u1_uk_n1749, u1_uk_n1801, u1_uk_n1803, u1_uk_n1804, u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, 
        u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1816, u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n182, u1_uk_n1824, 
        u1_uk_n1826, u1_uk_n1831, u1_uk_n1834, u1_uk_n1835, u1_uk_n1841, u1_uk_n1842, u1_uk_n187, u1_uk_n188, u1_uk_n191, 
        u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, u1_uk_n209, u1_uk_n213, u1_uk_n214, u1_uk_n217, u1_uk_n220, 
        u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, 
        u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, 
        u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n60, u1_uk_n63, u1_uk_n94, u1_uk_n99, u2_FP_52, u2_FP_53, 
        u2_FP_54, u2_FP_55, u2_FP_56, u2_FP_57, u2_FP_58, u2_FP_59, u2_FP_60, u2_FP_61, u2_K16_31, 
        u2_K16_42, u2_K7_26, u2_K7_31, u2_K7_33, u2_K7_35, u2_K7_37, u2_K7_38, u2_K7_43, u2_K7_45, 
        u2_K7_48, u2_L14_11, u2_L14_12, u2_L14_19, u2_L14_22, u2_L14_29, u2_L14_32, u2_L14_4, u2_L14_7, 
        u2_L5_11, u2_L5_12, u2_L5_14, u2_L5_15, u2_L5_19, u2_L5_21, u2_L5_22, u2_L5_25, u2_L5_27, 
        u2_L5_29, u2_L5_3, u2_L5_32, u2_L5_4, u2_L5_5, u2_L5_7, u2_L5_8, u2_R5_1, u2_R5_16, 
        u2_R5_17, u2_R5_18, u2_R5_19, u2_R5_20, u2_R5_21, u2_R5_22, u2_R5_23, u2_R5_24, u2_R5_25, 
        u2_R5_26, u2_R5_27, u2_R5_28, u2_R5_29, u2_R5_30, u2_R5_31, u2_R5_32, u2_key_r_50, u2_uk_K_r14_15, 
        u2_uk_K_r14_2, u2_uk_K_r14_50, u2_uk_K_r14_9, u2_uk_K_r5_0, u2_uk_K_r5_1, u2_uk_K_r5_21, u2_uk_K_r5_23, u2_uk_K_r5_31, u2_uk_K_r5_43, 
        u2_uk_K_r5_51, u2_uk_K_r5_7, u2_uk_n10, u2_uk_n1089, u2_uk_n1093, u2_uk_n1094, u2_uk_n11, u2_uk_n117, u2_uk_n118, 
        u2_uk_n1188, u2_uk_n1201, u2_uk_n1203, u2_uk_n1208, u2_uk_n1209, u2_uk_n1210, u2_uk_n1215, u2_uk_n1217, u2_uk_n1220, 
        u2_uk_n1225, u2_uk_n1226, u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n1452, u2_uk_n1456, u2_uk_n1459, 
        u2_uk_n1460, u2_uk_n1464, u2_uk_n147, u2_uk_n1470, u2_uk_n1471, u2_uk_n1480, u2_uk_n1486, u2_uk_n1490, u2_uk_n1491, 
        u2_uk_n1493, u2_uk_n161, u2_uk_n164, u2_uk_n182, u2_uk_n202, u2_uk_n208, u2_uk_n213, u2_uk_n217, u2_uk_n223, 
        u2_uk_n231, u2_uk_n238, u2_uk_n94, u2_uk_n961;
  output u0_N451, u0_N458, u0_N466, u0_N476, u0_N68, u0_N70, u0_N75, u0_N78, u0_N84, 
        u0_N85, u0_N90, u0_N95, u0_uk_n191, u0_uk_n63, u0_uk_n777, u1_FP_1, u1_FP_10, u1_FP_13, 
        u1_FP_17, u1_FP_18, u1_FP_2, u1_FP_20, u1_FP_23, u1_FP_26, u1_FP_28, u1_FP_31, u1_FP_9, 
        u1_N100, u1_N101, u1_N104, u1_N105, u1_N110, u1_N111, u1_N112, u1_N115, u1_N116, 
        u1_N118, u1_N119, u1_N121, u1_N122, u1_N125, u1_N126, u1_N228, u1_N238, u1_N244, 
        u1_N250, u1_N291, u1_N294, u1_N298, u1_N299, u1_N306, u1_N309, u1_N316, u1_N319, 
        u1_N355, u1_N356, u1_N358, u1_N362, u1_N363, u1_N366, u1_N370, u1_N372, u1_N373, 
        u1_N378, u1_N380, u1_N383, u1_N417, u1_N421, u1_N424, u1_N428, u1_N431, u1_N432, 
        u1_N433, u1_N438, u1_N439, u1_N443, u1_N445, u1_N446, u1_N96, u1_uk_n117, u1_uk_n83, 
        u2_FP_11, u2_FP_12, u2_FP_19, u2_FP_22, u2_FP_29, u2_FP_32, u2_FP_4, u2_FP_7, u2_N194, 
        u2_N195, u2_N196, u2_N198, u2_N199, u2_N202, u2_N203, u2_N205, u2_N206, u2_N210, 
        u2_N212, u2_N213, u2_N216, u2_N218, u2_N220, u2_N223, u2_uk_n31, u2_uk_n983;
  wire u0_K15_31, u0_K15_32, u0_K15_33, u0_K15_34, u0_K15_35, u0_K15_36, u0_K3_37, u0_K3_38, u0_K3_39, 
       u0_K3_40, u0_K3_41, u0_K3_42, u0_K3_43, u0_K3_44, u0_K3_45, u0_K3_46, u0_K3_47, u0_K3_48, 
       u0_out14_11, u0_out14_19, u0_out14_29, u0_out14_4, u0_out2_12, u0_out2_15, u0_out2_21, u0_out2_22, u0_out2_27, 
       u0_out2_32, u0_out2_5, u0_out2_7, u0_u14_X_31, u0_u14_X_32, u0_u14_X_33, u0_u14_X_34, u0_u14_X_35, u0_u14_X_36, 
       u0_u14_u5_n100, u0_u14_u5_n101, u0_u14_u5_n102, u0_u14_u5_n103, u0_u14_u5_n104, u0_u14_u5_n105, u0_u14_u5_n106, u0_u14_u5_n107, u0_u14_u5_n108, 
       u0_u14_u5_n109, u0_u14_u5_n110, u0_u14_u5_n111, u0_u14_u5_n112, u0_u14_u5_n113, u0_u14_u5_n114, u0_u14_u5_n115, u0_u14_u5_n116, u0_u14_u5_n117, 
       u0_u14_u5_n118, u0_u14_u5_n119, u0_u14_u5_n120, u0_u14_u5_n121, u0_u14_u5_n122, u0_u14_u5_n123, u0_u14_u5_n124, u0_u14_u5_n125, u0_u14_u5_n126, 
       u0_u14_u5_n127, u0_u14_u5_n128, u0_u14_u5_n129, u0_u14_u5_n130, u0_u14_u5_n131, u0_u14_u5_n132, u0_u14_u5_n133, u0_u14_u5_n134, u0_u14_u5_n135, 
       u0_u14_u5_n136, u0_u14_u5_n137, u0_u14_u5_n138, u0_u14_u5_n139, u0_u14_u5_n140, u0_u14_u5_n141, u0_u14_u5_n142, u0_u14_u5_n143, u0_u14_u5_n144, 
       u0_u14_u5_n145, u0_u14_u5_n146, u0_u14_u5_n147, u0_u14_u5_n148, u0_u14_u5_n149, u0_u14_u5_n150, u0_u14_u5_n151, u0_u14_u5_n152, u0_u14_u5_n153, 
       u0_u14_u5_n154, u0_u14_u5_n155, u0_u14_u5_n156, u0_u14_u5_n157, u0_u14_u5_n158, u0_u14_u5_n159, u0_u14_u5_n160, u0_u14_u5_n161, u0_u14_u5_n162, 
       u0_u14_u5_n163, u0_u14_u5_n164, u0_u14_u5_n165, u0_u14_u5_n166, u0_u14_u5_n167, u0_u14_u5_n168, u0_u14_u5_n169, u0_u14_u5_n170, u0_u14_u5_n171, 
       u0_u14_u5_n172, u0_u14_u5_n173, u0_u14_u5_n174, u0_u14_u5_n175, u0_u14_u5_n176, u0_u14_u5_n177, u0_u14_u5_n178, u0_u14_u5_n179, u0_u14_u5_n180, 
       u0_u14_u5_n181, u0_u14_u5_n182, u0_u14_u5_n183, u0_u14_u5_n184, u0_u14_u5_n185, u0_u14_u5_n186, u0_u14_u5_n187, u0_u14_u5_n188, u0_u14_u5_n189, 
       u0_u14_u5_n190, u0_u14_u5_n191, u0_u14_u5_n192, u0_u14_u5_n193, u0_u14_u5_n194, u0_u14_u5_n195, u0_u14_u5_n196, u0_u14_u5_n99, u0_u2_X_37, 
       u0_u2_X_38, u0_u2_X_39, u0_u2_X_40, u0_u2_X_41, u0_u2_X_42, u0_u2_X_43, u0_u2_X_44, u0_u2_X_45, u0_u2_X_46, 
       u0_u2_X_47, u0_u2_X_48, u0_u2_u6_n100, u0_u2_u6_n101, u0_u2_u6_n102, u0_u2_u6_n103, u0_u2_u6_n104, u0_u2_u6_n105, u0_u2_u6_n106, 
       u0_u2_u6_n107, u0_u2_u6_n108, u0_u2_u6_n109, u0_u2_u6_n110, u0_u2_u6_n111, u0_u2_u6_n112, u0_u2_u6_n113, u0_u2_u6_n114, u0_u2_u6_n115, 
       u0_u2_u6_n116, u0_u2_u6_n117, u0_u2_u6_n118, u0_u2_u6_n119, u0_u2_u6_n120, u0_u2_u6_n121, u0_u2_u6_n122, u0_u2_u6_n123, u0_u2_u6_n124, 
       u0_u2_u6_n125, u0_u2_u6_n126, u0_u2_u6_n127, u0_u2_u6_n128, u0_u2_u6_n129, u0_u2_u6_n130, u0_u2_u6_n131, u0_u2_u6_n132, u0_u2_u6_n133, 
       u0_u2_u6_n134, u0_u2_u6_n135, u0_u2_u6_n136, u0_u2_u6_n137, u0_u2_u6_n138, u0_u2_u6_n139, u0_u2_u6_n140, u0_u2_u6_n141, u0_u2_u6_n142, 
       u0_u2_u6_n143, u0_u2_u6_n144, u0_u2_u6_n145, u0_u2_u6_n146, u0_u2_u6_n147, u0_u2_u6_n148, u0_u2_u6_n149, u0_u2_u6_n150, u0_u2_u6_n151, 
       u0_u2_u6_n152, u0_u2_u6_n153, u0_u2_u6_n154, u0_u2_u6_n155, u0_u2_u6_n156, u0_u2_u6_n157, u0_u2_u6_n158, u0_u2_u6_n159, u0_u2_u6_n160, 
       u0_u2_u6_n161, u0_u2_u6_n162, u0_u2_u6_n163, u0_u2_u6_n164, u0_u2_u6_n165, u0_u2_u6_n166, u0_u2_u6_n167, u0_u2_u6_n168, u0_u2_u6_n169, 
       u0_u2_u6_n170, u0_u2_u6_n171, u0_u2_u6_n172, u0_u2_u6_n173, u0_u2_u6_n174, u0_u2_u6_n88, u0_u2_u6_n89, u0_u2_u6_n90, u0_u2_u6_n91, 
       u0_u2_u6_n92, u0_u2_u6_n93, u0_u2_u6_n94, u0_u2_u6_n95, u0_u2_u6_n96, u0_u2_u6_n97, u0_u2_u6_n98, u0_u2_u6_n99, u0_u2_u7_n100, 
       u0_u2_u7_n101, u0_u2_u7_n102, u0_u2_u7_n103, u0_u2_u7_n104, u0_u2_u7_n105, u0_u2_u7_n106, u0_u2_u7_n107, u0_u2_u7_n108, u0_u2_u7_n109, 
       u0_u2_u7_n110, u0_u2_u7_n111, u0_u2_u7_n112, u0_u2_u7_n113, u0_u2_u7_n114, u0_u2_u7_n115, u0_u2_u7_n116, u0_u2_u7_n117, u0_u2_u7_n118, 
       u0_u2_u7_n119, u0_u2_u7_n120, u0_u2_u7_n121, u0_u2_u7_n122, u0_u2_u7_n123, u0_u2_u7_n124, u0_u2_u7_n125, u0_u2_u7_n126, u0_u2_u7_n127, 
       u0_u2_u7_n128, u0_u2_u7_n129, u0_u2_u7_n130, u0_u2_u7_n131, u0_u2_u7_n132, u0_u2_u7_n133, u0_u2_u7_n134, u0_u2_u7_n135, u0_u2_u7_n136, 
       u0_u2_u7_n137, u0_u2_u7_n138, u0_u2_u7_n139, u0_u2_u7_n140, u0_u2_u7_n141, u0_u2_u7_n142, u0_u2_u7_n143, u0_u2_u7_n144, u0_u2_u7_n145, 
       u0_u2_u7_n146, u0_u2_u7_n147, u0_u2_u7_n148, u0_u2_u7_n149, u0_u2_u7_n150, u0_u2_u7_n151, u0_u2_u7_n152, u0_u2_u7_n153, u0_u2_u7_n154, 
       u0_u2_u7_n155, u0_u2_u7_n156, u0_u2_u7_n157, u0_u2_u7_n158, u0_u2_u7_n159, u0_u2_u7_n160, u0_u2_u7_n161, u0_u2_u7_n162, u0_u2_u7_n163, 
       u0_u2_u7_n164, u0_u2_u7_n165, u0_u2_u7_n166, u0_u2_u7_n167, u0_u2_u7_n168, u0_u2_u7_n169, u0_u2_u7_n170, u0_u2_u7_n171, u0_u2_u7_n172, 
       u0_u2_u7_n173, u0_u2_u7_n174, u0_u2_u7_n175, u0_u2_u7_n176, u0_u2_u7_n177, u0_u2_u7_n178, u0_u2_u7_n179, u0_u2_u7_n180, u0_u2_u7_n91, 
       u0_u2_u7_n92, u0_u2_u7_n93, u0_u2_u7_n94, u0_u2_u7_n95, u0_u2_u7_n96, u0_u2_u7_n97, u0_u2_u7_n98, u0_u2_u7_n99, u0_uk_n842, 
       u0_uk_n843, u0_uk_n844, u0_uk_n845, u1_K10_31, u1_K10_32, u1_K10_33, u1_K10_34, u1_K10_35, u1_K10_36, 
       u1_K10_37, u1_K10_38, u1_K10_39, u1_K10_40, u1_K10_41, u1_K10_42, u1_K12_31, u1_K12_32, u1_K12_33, 
       u1_K12_34, u1_K12_35, u1_K12_36, u1_K12_37, u1_K12_38, u1_K12_39, u1_K12_40, u1_K12_41, u1_K12_42, 
       u1_K12_43, u1_K12_44, u1_K12_45, u1_K12_46, u1_K12_47, u1_K12_48, u1_K14_1, u1_K14_10, u1_K14_11, 
       u1_K14_12, u1_K14_13, u1_K14_14, u1_K14_15, u1_K14_16, u1_K14_17, u1_K14_18, u1_K14_2, u1_K14_3, 
       u1_K14_4, u1_K14_5, u1_K14_6, u1_K14_7, u1_K14_8, u1_K14_9, u1_K16_1, u1_K16_10, u1_K16_11, 
       u1_K16_12, u1_K16_19, u1_K16_2, u1_K16_20, u1_K16_21, u1_K16_22, u1_K16_23, u1_K16_24, u1_K16_3, 
       u1_K16_4, u1_K16_5, u1_K16_6, u1_K16_7, u1_K16_8, u1_K16_9, u1_K4_1, u1_K4_13, u1_K4_14, 
       u1_K4_15, u1_K4_16, u1_K4_17, u1_K4_18, u1_K4_19, u1_K4_2, u1_K4_20, u1_K4_21, u1_K4_22, 
       u1_K4_23, u1_K4_24, u1_K4_3, u1_K4_4, u1_K4_43, u1_K4_44, u1_K4_45, u1_K4_46, u1_K4_47, 
       u1_K4_48, u1_K4_5, u1_K4_6, u1_K8_43, u1_K8_44, u1_K8_45, u1_K8_46, u1_K8_47, u1_K8_48, 
       u1_out11_11, u1_out11_12, u1_out11_15, u1_out11_19, u1_out11_21, u1_out11_22, u1_out11_27, u1_out11_29, u1_out11_32, 
       u1_out11_4, u1_out11_5, u1_out11_7, u1_out13_13, u1_out13_16, u1_out13_17, u1_out13_18, u1_out13_2, u1_out13_23, 
       u1_out13_24, u1_out13_28, u1_out13_30, u1_out13_31, u1_out13_6, u1_out13_9, u1_out15_1, u1_out15_10, u1_out15_13, 
       u1_out15_17, u1_out15_18, u1_out15_2, u1_out15_20, u1_out15_23, u1_out15_26, u1_out15_28, u1_out15_31, u1_out15_9, 
       u1_out3_1, u1_out3_10, u1_out3_15, u1_out3_16, u1_out3_17, u1_out3_20, u1_out3_21, u1_out3_23, u1_out3_24, 
       u1_out3_26, u1_out3_27, u1_out3_30, u1_out3_31, u1_out3_5, u1_out3_6, u1_out3_9, u1_out7_15, u1_out7_21, 
       u1_out7_27, u1_out7_5, u1_out9_11, u1_out9_12, u1_out9_19, u1_out9_22, u1_out9_29, u1_out9_32, u1_out9_4, 
       u1_out9_7, u1_u11_X_31, u1_u11_X_32, u1_u11_X_33, u1_u11_X_34, u1_u11_X_35, u1_u11_X_36, u1_u11_X_37, u1_u11_X_38, 
       u1_u11_X_39, u1_u11_X_40, u1_u11_X_41, u1_u11_X_42, u1_u11_X_43, u1_u11_X_44, u1_u11_X_45, u1_u11_X_46, u1_u11_X_47, 
       u1_u11_X_48, u1_u11_u5_n100, u1_u11_u5_n101, u1_u11_u5_n102, u1_u11_u5_n103, u1_u11_u5_n104, u1_u11_u5_n105, u1_u11_u5_n106, u1_u11_u5_n107, 
       u1_u11_u5_n108, u1_u11_u5_n109, u1_u11_u5_n110, u1_u11_u5_n111, u1_u11_u5_n112, u1_u11_u5_n113, u1_u11_u5_n114, u1_u11_u5_n115, u1_u11_u5_n116, 
       u1_u11_u5_n117, u1_u11_u5_n118, u1_u11_u5_n119, u1_u11_u5_n120, u1_u11_u5_n121, u1_u11_u5_n122, u1_u11_u5_n123, u1_u11_u5_n124, u1_u11_u5_n125, 
       u1_u11_u5_n126, u1_u11_u5_n127, u1_u11_u5_n128, u1_u11_u5_n129, u1_u11_u5_n130, u1_u11_u5_n131, u1_u11_u5_n132, u1_u11_u5_n133, u1_u11_u5_n134, 
       u1_u11_u5_n135, u1_u11_u5_n136, u1_u11_u5_n137, u1_u11_u5_n138, u1_u11_u5_n139, u1_u11_u5_n140, u1_u11_u5_n141, u1_u11_u5_n142, u1_u11_u5_n143, 
       u1_u11_u5_n144, u1_u11_u5_n145, u1_u11_u5_n146, u1_u11_u5_n147, u1_u11_u5_n148, u1_u11_u5_n149, u1_u11_u5_n150, u1_u11_u5_n151, u1_u11_u5_n152, 
       u1_u11_u5_n153, u1_u11_u5_n154, u1_u11_u5_n155, u1_u11_u5_n156, u1_u11_u5_n157, u1_u11_u5_n158, u1_u11_u5_n159, u1_u11_u5_n160, u1_u11_u5_n161, 
       u1_u11_u5_n162, u1_u11_u5_n163, u1_u11_u5_n164, u1_u11_u5_n165, u1_u11_u5_n166, u1_u11_u5_n167, u1_u11_u5_n168, u1_u11_u5_n169, u1_u11_u5_n170, 
       u1_u11_u5_n171, u1_u11_u5_n172, u1_u11_u5_n173, u1_u11_u5_n174, u1_u11_u5_n175, u1_u11_u5_n176, u1_u11_u5_n177, u1_u11_u5_n178, u1_u11_u5_n179, 
       u1_u11_u5_n180, u1_u11_u5_n181, u1_u11_u5_n182, u1_u11_u5_n183, u1_u11_u5_n184, u1_u11_u5_n185, u1_u11_u5_n186, u1_u11_u5_n187, u1_u11_u5_n188, 
       u1_u11_u5_n189, u1_u11_u5_n190, u1_u11_u5_n191, u1_u11_u5_n192, u1_u11_u5_n193, u1_u11_u5_n194, u1_u11_u5_n195, u1_u11_u5_n196, u1_u11_u5_n99, 
       u1_u11_u6_n100, u1_u11_u6_n101, u1_u11_u6_n102, u1_u11_u6_n103, u1_u11_u6_n104, u1_u11_u6_n105, u1_u11_u6_n106, u1_u11_u6_n107, u1_u11_u6_n108, 
       u1_u11_u6_n109, u1_u11_u6_n110, u1_u11_u6_n111, u1_u11_u6_n112, u1_u11_u6_n113, u1_u11_u6_n114, u1_u11_u6_n115, u1_u11_u6_n116, u1_u11_u6_n117, 
       u1_u11_u6_n118, u1_u11_u6_n119, u1_u11_u6_n120, u1_u11_u6_n121, u1_u11_u6_n122, u1_u11_u6_n123, u1_u11_u6_n124, u1_u11_u6_n125, u1_u11_u6_n126, 
       u1_u11_u6_n127, u1_u11_u6_n128, u1_u11_u6_n129, u1_u11_u6_n130, u1_u11_u6_n131, u1_u11_u6_n132, u1_u11_u6_n133, u1_u11_u6_n134, u1_u11_u6_n135, 
       u1_u11_u6_n136, u1_u11_u6_n137, u1_u11_u6_n138, u1_u11_u6_n139, u1_u11_u6_n140, u1_u11_u6_n141, u1_u11_u6_n142, u1_u11_u6_n143, u1_u11_u6_n144, 
       u1_u11_u6_n145, u1_u11_u6_n146, u1_u11_u6_n147, u1_u11_u6_n148, u1_u11_u6_n149, u1_u11_u6_n150, u1_u11_u6_n151, u1_u11_u6_n152, u1_u11_u6_n153, 
       u1_u11_u6_n154, u1_u11_u6_n155, u1_u11_u6_n156, u1_u11_u6_n157, u1_u11_u6_n158, u1_u11_u6_n159, u1_u11_u6_n160, u1_u11_u6_n161, u1_u11_u6_n162, 
       u1_u11_u6_n163, u1_u11_u6_n164, u1_u11_u6_n165, u1_u11_u6_n166, u1_u11_u6_n167, u1_u11_u6_n168, u1_u11_u6_n169, u1_u11_u6_n170, u1_u11_u6_n171, 
       u1_u11_u6_n172, u1_u11_u6_n173, u1_u11_u6_n174, u1_u11_u6_n88, u1_u11_u6_n89, u1_u11_u6_n90, u1_u11_u6_n91, u1_u11_u6_n92, u1_u11_u6_n93, 
       u1_u11_u6_n94, u1_u11_u6_n95, u1_u11_u6_n96, u1_u11_u6_n97, u1_u11_u6_n98, u1_u11_u6_n99, u1_u11_u7_n100, u1_u11_u7_n101, u1_u11_u7_n102, 
       u1_u11_u7_n103, u1_u11_u7_n104, u1_u11_u7_n105, u1_u11_u7_n106, u1_u11_u7_n107, u1_u11_u7_n108, u1_u11_u7_n109, u1_u11_u7_n110, u1_u11_u7_n111, 
       u1_u11_u7_n112, u1_u11_u7_n113, u1_u11_u7_n114, u1_u11_u7_n115, u1_u11_u7_n116, u1_u11_u7_n117, u1_u11_u7_n118, u1_u11_u7_n119, u1_u11_u7_n120, 
       u1_u11_u7_n121, u1_u11_u7_n122, u1_u11_u7_n123, u1_u11_u7_n124, u1_u11_u7_n125, u1_u11_u7_n126, u1_u11_u7_n127, u1_u11_u7_n128, u1_u11_u7_n129, 
       u1_u11_u7_n130, u1_u11_u7_n131, u1_u11_u7_n132, u1_u11_u7_n133, u1_u11_u7_n134, u1_u11_u7_n135, u1_u11_u7_n136, u1_u11_u7_n137, u1_u11_u7_n138, 
       u1_u11_u7_n139, u1_u11_u7_n140, u1_u11_u7_n141, u1_u11_u7_n142, u1_u11_u7_n143, u1_u11_u7_n144, u1_u11_u7_n145, u1_u11_u7_n146, u1_u11_u7_n147, 
       u1_u11_u7_n148, u1_u11_u7_n149, u1_u11_u7_n150, u1_u11_u7_n151, u1_u11_u7_n152, u1_u11_u7_n153, u1_u11_u7_n154, u1_u11_u7_n155, u1_u11_u7_n156, 
       u1_u11_u7_n157, u1_u11_u7_n158, u1_u11_u7_n159, u1_u11_u7_n160, u1_u11_u7_n161, u1_u11_u7_n162, u1_u11_u7_n163, u1_u11_u7_n164, u1_u11_u7_n165, 
       u1_u11_u7_n166, u1_u11_u7_n167, u1_u11_u7_n168, u1_u11_u7_n169, u1_u11_u7_n170, u1_u11_u7_n171, u1_u11_u7_n172, u1_u11_u7_n173, u1_u11_u7_n174, 
       u1_u11_u7_n175, u1_u11_u7_n176, u1_u11_u7_n177, u1_u11_u7_n178, u1_u11_u7_n179, u1_u11_u7_n180, u1_u11_u7_n91, u1_u11_u7_n92, u1_u11_u7_n93, 
       u1_u11_u7_n94, u1_u11_u7_n95, u1_u11_u7_n96, u1_u11_u7_n97, u1_u11_u7_n98, u1_u11_u7_n99, u1_u13_X_1, u1_u13_X_10, u1_u13_X_11, 
       u1_u13_X_12, u1_u13_X_13, u1_u13_X_14, u1_u13_X_15, u1_u13_X_16, u1_u13_X_17, u1_u13_X_18, u1_u13_X_2, u1_u13_X_3, 
       u1_u13_X_4, u1_u13_X_5, u1_u13_X_6, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, u1_u13_u0_n100, u1_u13_u0_n101, u1_u13_u0_n102, 
       u1_u13_u0_n103, u1_u13_u0_n104, u1_u13_u0_n105, u1_u13_u0_n106, u1_u13_u0_n107, u1_u13_u0_n108, u1_u13_u0_n109, u1_u13_u0_n110, u1_u13_u0_n111, 
       u1_u13_u0_n112, u1_u13_u0_n113, u1_u13_u0_n114, u1_u13_u0_n115, u1_u13_u0_n116, u1_u13_u0_n117, u1_u13_u0_n118, u1_u13_u0_n119, u1_u13_u0_n120, 
       u1_u13_u0_n121, u1_u13_u0_n122, u1_u13_u0_n123, u1_u13_u0_n124, u1_u13_u0_n125, u1_u13_u0_n126, u1_u13_u0_n127, u1_u13_u0_n128, u1_u13_u0_n129, 
       u1_u13_u0_n130, u1_u13_u0_n131, u1_u13_u0_n132, u1_u13_u0_n133, u1_u13_u0_n134, u1_u13_u0_n135, u1_u13_u0_n136, u1_u13_u0_n137, u1_u13_u0_n138, 
       u1_u13_u0_n139, u1_u13_u0_n140, u1_u13_u0_n141, u1_u13_u0_n142, u1_u13_u0_n143, u1_u13_u0_n144, u1_u13_u0_n145, u1_u13_u0_n146, u1_u13_u0_n147, 
       u1_u13_u0_n148, u1_u13_u0_n149, u1_u13_u0_n150, u1_u13_u0_n151, u1_u13_u0_n152, u1_u13_u0_n153, u1_u13_u0_n154, u1_u13_u0_n155, u1_u13_u0_n156, 
       u1_u13_u0_n157, u1_u13_u0_n158, u1_u13_u0_n159, u1_u13_u0_n160, u1_u13_u0_n161, u1_u13_u0_n162, u1_u13_u0_n163, u1_u13_u0_n164, u1_u13_u0_n165, 
       u1_u13_u0_n166, u1_u13_u0_n167, u1_u13_u0_n168, u1_u13_u0_n169, u1_u13_u0_n170, u1_u13_u0_n171, u1_u13_u0_n172, u1_u13_u0_n173, u1_u13_u0_n174, 
       u1_u13_u0_n88, u1_u13_u0_n89, u1_u13_u0_n90, u1_u13_u0_n91, u1_u13_u0_n92, u1_u13_u0_n93, u1_u13_u0_n94, u1_u13_u0_n95, u1_u13_u0_n96, 
       u1_u13_u0_n97, u1_u13_u0_n98, u1_u13_u0_n99, u1_u13_u1_n100, u1_u13_u1_n101, u1_u13_u1_n102, u1_u13_u1_n103, u1_u13_u1_n104, u1_u13_u1_n105, 
       u1_u13_u1_n106, u1_u13_u1_n107, u1_u13_u1_n108, u1_u13_u1_n109, u1_u13_u1_n110, u1_u13_u1_n111, u1_u13_u1_n112, u1_u13_u1_n113, u1_u13_u1_n114, 
       u1_u13_u1_n115, u1_u13_u1_n116, u1_u13_u1_n117, u1_u13_u1_n118, u1_u13_u1_n119, u1_u13_u1_n120, u1_u13_u1_n121, u1_u13_u1_n122, u1_u13_u1_n123, 
       u1_u13_u1_n124, u1_u13_u1_n125, u1_u13_u1_n126, u1_u13_u1_n127, u1_u13_u1_n128, u1_u13_u1_n129, u1_u13_u1_n130, u1_u13_u1_n131, u1_u13_u1_n132, 
       u1_u13_u1_n133, u1_u13_u1_n134, u1_u13_u1_n135, u1_u13_u1_n136, u1_u13_u1_n137, u1_u13_u1_n138, u1_u13_u1_n139, u1_u13_u1_n140, u1_u13_u1_n141, 
       u1_u13_u1_n142, u1_u13_u1_n143, u1_u13_u1_n144, u1_u13_u1_n145, u1_u13_u1_n146, u1_u13_u1_n147, u1_u13_u1_n148, u1_u13_u1_n149, u1_u13_u1_n150, 
       u1_u13_u1_n151, u1_u13_u1_n152, u1_u13_u1_n153, u1_u13_u1_n154, u1_u13_u1_n155, u1_u13_u1_n156, u1_u13_u1_n157, u1_u13_u1_n158, u1_u13_u1_n159, 
       u1_u13_u1_n160, u1_u13_u1_n161, u1_u13_u1_n162, u1_u13_u1_n163, u1_u13_u1_n164, u1_u13_u1_n165, u1_u13_u1_n166, u1_u13_u1_n167, u1_u13_u1_n168, 
       u1_u13_u1_n169, u1_u13_u1_n170, u1_u13_u1_n171, u1_u13_u1_n172, u1_u13_u1_n173, u1_u13_u1_n174, u1_u13_u1_n175, u1_u13_u1_n176, u1_u13_u1_n177, 
       u1_u13_u1_n178, u1_u13_u1_n179, u1_u13_u1_n180, u1_u13_u1_n181, u1_u13_u1_n182, u1_u13_u1_n183, u1_u13_u1_n184, u1_u13_u1_n185, u1_u13_u1_n186, 
       u1_u13_u1_n187, u1_u13_u1_n188, u1_u13_u1_n95, u1_u13_u1_n96, u1_u13_u1_n97, u1_u13_u1_n98, u1_u13_u1_n99, u1_u13_u2_n100, u1_u13_u2_n101, 
       u1_u13_u2_n102, u1_u13_u2_n103, u1_u13_u2_n104, u1_u13_u2_n105, u1_u13_u2_n106, u1_u13_u2_n107, u1_u13_u2_n108, u1_u13_u2_n109, u1_u13_u2_n110, 
       u1_u13_u2_n111, u1_u13_u2_n112, u1_u13_u2_n113, u1_u13_u2_n114, u1_u13_u2_n115, u1_u13_u2_n116, u1_u13_u2_n117, u1_u13_u2_n118, u1_u13_u2_n119, 
       u1_u13_u2_n120, u1_u13_u2_n121, u1_u13_u2_n122, u1_u13_u2_n123, u1_u13_u2_n124, u1_u13_u2_n125, u1_u13_u2_n126, u1_u13_u2_n127, u1_u13_u2_n128, 
       u1_u13_u2_n129, u1_u13_u2_n130, u1_u13_u2_n131, u1_u13_u2_n132, u1_u13_u2_n133, u1_u13_u2_n134, u1_u13_u2_n135, u1_u13_u2_n136, u1_u13_u2_n137, 
       u1_u13_u2_n138, u1_u13_u2_n139, u1_u13_u2_n140, u1_u13_u2_n141, u1_u13_u2_n142, u1_u13_u2_n143, u1_u13_u2_n144, u1_u13_u2_n145, u1_u13_u2_n146, 
       u1_u13_u2_n147, u1_u13_u2_n148, u1_u13_u2_n149, u1_u13_u2_n150, u1_u13_u2_n151, u1_u13_u2_n152, u1_u13_u2_n153, u1_u13_u2_n154, u1_u13_u2_n155, 
       u1_u13_u2_n156, u1_u13_u2_n157, u1_u13_u2_n158, u1_u13_u2_n159, u1_u13_u2_n160, u1_u13_u2_n161, u1_u13_u2_n162, u1_u13_u2_n163, u1_u13_u2_n164, 
       u1_u13_u2_n165, u1_u13_u2_n166, u1_u13_u2_n167, u1_u13_u2_n168, u1_u13_u2_n169, u1_u13_u2_n170, u1_u13_u2_n171, u1_u13_u2_n172, u1_u13_u2_n173, 
       u1_u13_u2_n174, u1_u13_u2_n175, u1_u13_u2_n176, u1_u13_u2_n177, u1_u13_u2_n178, u1_u13_u2_n179, u1_u13_u2_n180, u1_u13_u2_n181, u1_u13_u2_n182, 
       u1_u13_u2_n183, u1_u13_u2_n184, u1_u13_u2_n185, u1_u13_u2_n186, u1_u13_u2_n187, u1_u13_u2_n188, u1_u13_u2_n95, u1_u13_u2_n96, u1_u13_u2_n97, 
       u1_u13_u2_n98, u1_u13_u2_n99, u1_u15_X_1, u1_u15_X_10, u1_u15_X_11, u1_u15_X_12, u1_u15_X_19, u1_u15_X_2, u1_u15_X_20, 
       u1_u15_X_21, u1_u15_X_22, u1_u15_X_23, u1_u15_X_24, u1_u15_X_3, u1_u15_X_4, u1_u15_X_5, u1_u15_X_6, u1_u15_X_7, 
       u1_u15_X_8, u1_u15_X_9, u1_u15_u0_n100, u1_u15_u0_n101, u1_u15_u0_n102, u1_u15_u0_n103, u1_u15_u0_n104, u1_u15_u0_n105, u1_u15_u0_n106, 
       u1_u15_u0_n107, u1_u15_u0_n108, u1_u15_u0_n109, u1_u15_u0_n110, u1_u15_u0_n111, u1_u15_u0_n112, u1_u15_u0_n113, u1_u15_u0_n114, u1_u15_u0_n115, 
       u1_u15_u0_n116, u1_u15_u0_n117, u1_u15_u0_n118, u1_u15_u0_n119, u1_u15_u0_n120, u1_u15_u0_n121, u1_u15_u0_n122, u1_u15_u0_n123, u1_u15_u0_n124, 
       u1_u15_u0_n125, u1_u15_u0_n126, u1_u15_u0_n127, u1_u15_u0_n128, u1_u15_u0_n129, u1_u15_u0_n130, u1_u15_u0_n131, u1_u15_u0_n132, u1_u15_u0_n133, 
       u1_u15_u0_n134, u1_u15_u0_n135, u1_u15_u0_n136, u1_u15_u0_n137, u1_u15_u0_n138, u1_u15_u0_n139, u1_u15_u0_n140, u1_u15_u0_n141, u1_u15_u0_n142, 
       u1_u15_u0_n143, u1_u15_u0_n144, u1_u15_u0_n145, u1_u15_u0_n146, u1_u15_u0_n147, u1_u15_u0_n148, u1_u15_u0_n149, u1_u15_u0_n150, u1_u15_u0_n151, 
       u1_u15_u0_n152, u1_u15_u0_n153, u1_u15_u0_n154, u1_u15_u0_n155, u1_u15_u0_n156, u1_u15_u0_n157, u1_u15_u0_n158, u1_u15_u0_n159, u1_u15_u0_n160, 
       u1_u15_u0_n161, u1_u15_u0_n162, u1_u15_u0_n163, u1_u15_u0_n164, u1_u15_u0_n165, u1_u15_u0_n166, u1_u15_u0_n167, u1_u15_u0_n168, u1_u15_u0_n169, 
       u1_u15_u0_n170, u1_u15_u0_n171, u1_u15_u0_n172, u1_u15_u0_n173, u1_u15_u0_n174, u1_u15_u0_n88, u1_u15_u0_n89, u1_u15_u0_n90, u1_u15_u0_n91, 
       u1_u15_u0_n92, u1_u15_u0_n93, u1_u15_u0_n94, u1_u15_u0_n95, u1_u15_u0_n96, u1_u15_u0_n97, u1_u15_u0_n98, u1_u15_u0_n99, u1_u15_u1_n100, 
       u1_u15_u1_n101, u1_u15_u1_n102, u1_u15_u1_n103, u1_u15_u1_n104, u1_u15_u1_n105, u1_u15_u1_n106, u1_u15_u1_n107, u1_u15_u1_n108, u1_u15_u1_n109, 
       u1_u15_u1_n110, u1_u15_u1_n111, u1_u15_u1_n112, u1_u15_u1_n113, u1_u15_u1_n114, u1_u15_u1_n115, u1_u15_u1_n116, u1_u15_u1_n117, u1_u15_u1_n118, 
       u1_u15_u1_n119, u1_u15_u1_n120, u1_u15_u1_n121, u1_u15_u1_n122, u1_u15_u1_n123, u1_u15_u1_n124, u1_u15_u1_n125, u1_u15_u1_n126, u1_u15_u1_n127, 
       u1_u15_u1_n128, u1_u15_u1_n129, u1_u15_u1_n130, u1_u15_u1_n131, u1_u15_u1_n132, u1_u15_u1_n133, u1_u15_u1_n134, u1_u15_u1_n135, u1_u15_u1_n136, 
       u1_u15_u1_n137, u1_u15_u1_n138, u1_u15_u1_n139, u1_u15_u1_n140, u1_u15_u1_n141, u1_u15_u1_n142, u1_u15_u1_n143, u1_u15_u1_n144, u1_u15_u1_n145, 
       u1_u15_u1_n146, u1_u15_u1_n147, u1_u15_u1_n148, u1_u15_u1_n149, u1_u15_u1_n150, u1_u15_u1_n151, u1_u15_u1_n152, u1_u15_u1_n153, u1_u15_u1_n154, 
       u1_u15_u1_n155, u1_u15_u1_n156, u1_u15_u1_n157, u1_u15_u1_n158, u1_u15_u1_n159, u1_u15_u1_n160, u1_u15_u1_n161, u1_u15_u1_n162, u1_u15_u1_n163, 
       u1_u15_u1_n164, u1_u15_u1_n165, u1_u15_u1_n166, u1_u15_u1_n167, u1_u15_u1_n168, u1_u15_u1_n169, u1_u15_u1_n170, u1_u15_u1_n171, u1_u15_u1_n172, 
       u1_u15_u1_n173, u1_u15_u1_n174, u1_u15_u1_n175, u1_u15_u1_n176, u1_u15_u1_n177, u1_u15_u1_n178, u1_u15_u1_n179, u1_u15_u1_n180, u1_u15_u1_n181, 
       u1_u15_u1_n182, u1_u15_u1_n183, u1_u15_u1_n184, u1_u15_u1_n185, u1_u15_u1_n186, u1_u15_u1_n187, u1_u15_u1_n188, u1_u15_u1_n95, u1_u15_u1_n96, 
       u1_u15_u1_n97, u1_u15_u1_n98, u1_u15_u1_n99, u1_u15_u3_n100, u1_u15_u3_n101, u1_u15_u3_n102, u1_u15_u3_n103, u1_u15_u3_n104, u1_u15_u3_n105, 
       u1_u15_u3_n106, u1_u15_u3_n107, u1_u15_u3_n108, u1_u15_u3_n109, u1_u15_u3_n110, u1_u15_u3_n111, u1_u15_u3_n112, u1_u15_u3_n113, u1_u15_u3_n114, 
       u1_u15_u3_n115, u1_u15_u3_n116, u1_u15_u3_n117, u1_u15_u3_n118, u1_u15_u3_n119, u1_u15_u3_n120, u1_u15_u3_n121, u1_u15_u3_n122, u1_u15_u3_n123, 
       u1_u15_u3_n124, u1_u15_u3_n125, u1_u15_u3_n126, u1_u15_u3_n127, u1_u15_u3_n128, u1_u15_u3_n129, u1_u15_u3_n130, u1_u15_u3_n131, u1_u15_u3_n132, 
       u1_u15_u3_n133, u1_u15_u3_n134, u1_u15_u3_n135, u1_u15_u3_n136, u1_u15_u3_n137, u1_u15_u3_n138, u1_u15_u3_n139, u1_u15_u3_n140, u1_u15_u3_n141, 
       u1_u15_u3_n142, u1_u15_u3_n143, u1_u15_u3_n144, u1_u15_u3_n145, u1_u15_u3_n146, u1_u15_u3_n147, u1_u15_u3_n148, u1_u15_u3_n149, u1_u15_u3_n150, 
       u1_u15_u3_n151, u1_u15_u3_n152, u1_u15_u3_n153, u1_u15_u3_n154, u1_u15_u3_n155, u1_u15_u3_n156, u1_u15_u3_n157, u1_u15_u3_n158, u1_u15_u3_n159, 
       u1_u15_u3_n160, u1_u15_u3_n161, u1_u15_u3_n162, u1_u15_u3_n163, u1_u15_u3_n164, u1_u15_u3_n165, u1_u15_u3_n166, u1_u15_u3_n167, u1_u15_u3_n168, 
       u1_u15_u3_n169, u1_u15_u3_n170, u1_u15_u3_n171, u1_u15_u3_n172, u1_u15_u3_n173, u1_u15_u3_n174, u1_u15_u3_n175, u1_u15_u3_n176, u1_u15_u3_n177, 
       u1_u15_u3_n178, u1_u15_u3_n179, u1_u15_u3_n180, u1_u15_u3_n181, u1_u15_u3_n182, u1_u15_u3_n183, u1_u15_u3_n184, u1_u15_u3_n185, u1_u15_u3_n186, 
       u1_u15_u3_n94, u1_u15_u3_n95, u1_u15_u3_n96, u1_u15_u3_n97, u1_u15_u3_n98, u1_u15_u3_n99, u1_u3_X_1, u1_u3_X_13, u1_u3_X_14, 
       u1_u3_X_15, u1_u3_X_16, u1_u3_X_17, u1_u3_X_18, u1_u3_X_19, u1_u3_X_2, u1_u3_X_20, u1_u3_X_21, u1_u3_X_22, 
       u1_u3_X_23, u1_u3_X_24, u1_u3_X_3, u1_u3_X_4, u1_u3_X_43, u1_u3_X_44, u1_u3_X_45, u1_u3_X_46, u1_u3_X_47, 
       u1_u3_X_48, u1_u3_X_5, u1_u3_X_6, u1_u3_u0_n100, u1_u3_u0_n101, u1_u3_u0_n102, u1_u3_u0_n103, u1_u3_u0_n104, u1_u3_u0_n105, 
       u1_u3_u0_n106, u1_u3_u0_n107, u1_u3_u0_n108, u1_u3_u0_n109, u1_u3_u0_n110, u1_u3_u0_n111, u1_u3_u0_n112, u1_u3_u0_n113, u1_u3_u0_n114, 
       u1_u3_u0_n115, u1_u3_u0_n116, u1_u3_u0_n117, u1_u3_u0_n118, u1_u3_u0_n119, u1_u3_u0_n120, u1_u3_u0_n121, u1_u3_u0_n122, u1_u3_u0_n123, 
       u1_u3_u0_n124, u1_u3_u0_n125, u1_u3_u0_n126, u1_u3_u0_n127, u1_u3_u0_n128, u1_u3_u0_n129, u1_u3_u0_n130, u1_u3_u0_n131, u1_u3_u0_n132, 
       u1_u3_u0_n133, u1_u3_u0_n134, u1_u3_u0_n135, u1_u3_u0_n136, u1_u3_u0_n137, u1_u3_u0_n138, u1_u3_u0_n139, u1_u3_u0_n140, u1_u3_u0_n141, 
       u1_u3_u0_n142, u1_u3_u0_n143, u1_u3_u0_n144, u1_u3_u0_n145, u1_u3_u0_n146, u1_u3_u0_n147, u1_u3_u0_n148, u1_u3_u0_n149, u1_u3_u0_n150, 
       u1_u3_u0_n151, u1_u3_u0_n152, u1_u3_u0_n153, u1_u3_u0_n154, u1_u3_u0_n155, u1_u3_u0_n156, u1_u3_u0_n157, u1_u3_u0_n158, u1_u3_u0_n159, 
       u1_u3_u0_n160, u1_u3_u0_n161, u1_u3_u0_n162, u1_u3_u0_n163, u1_u3_u0_n164, u1_u3_u0_n165, u1_u3_u0_n166, u1_u3_u0_n167, u1_u3_u0_n168, 
       u1_u3_u0_n169, u1_u3_u0_n170, u1_u3_u0_n171, u1_u3_u0_n172, u1_u3_u0_n173, u1_u3_u0_n174, u1_u3_u0_n88, u1_u3_u0_n89, u1_u3_u0_n90, 
       u1_u3_u0_n91, u1_u3_u0_n92, u1_u3_u0_n93, u1_u3_u0_n94, u1_u3_u0_n95, u1_u3_u0_n96, u1_u3_u0_n97, u1_u3_u0_n98, u1_u3_u0_n99, 
       u1_u3_u2_n100, u1_u3_u2_n101, u1_u3_u2_n102, u1_u3_u2_n103, u1_u3_u2_n104, u1_u3_u2_n105, u1_u3_u2_n106, u1_u3_u2_n107, u1_u3_u2_n108, 
       u1_u3_u2_n109, u1_u3_u2_n110, u1_u3_u2_n111, u1_u3_u2_n112, u1_u3_u2_n113, u1_u3_u2_n114, u1_u3_u2_n115, u1_u3_u2_n116, u1_u3_u2_n117, 
       u1_u3_u2_n118, u1_u3_u2_n119, u1_u3_u2_n120, u1_u3_u2_n121, u1_u3_u2_n122, u1_u3_u2_n123, u1_u3_u2_n124, u1_u3_u2_n125, u1_u3_u2_n126, 
       u1_u3_u2_n127, u1_u3_u2_n128, u1_u3_u2_n129, u1_u3_u2_n130, u1_u3_u2_n131, u1_u3_u2_n132, u1_u3_u2_n133, u1_u3_u2_n134, u1_u3_u2_n135, 
       u1_u3_u2_n136, u1_u3_u2_n137, u1_u3_u2_n138, u1_u3_u2_n139, u1_u3_u2_n140, u1_u3_u2_n141, u1_u3_u2_n142, u1_u3_u2_n143, u1_u3_u2_n144, 
       u1_u3_u2_n145, u1_u3_u2_n146, u1_u3_u2_n147, u1_u3_u2_n148, u1_u3_u2_n149, u1_u3_u2_n150, u1_u3_u2_n151, u1_u3_u2_n152, u1_u3_u2_n153, 
       u1_u3_u2_n154, u1_u3_u2_n155, u1_u3_u2_n156, u1_u3_u2_n157, u1_u3_u2_n158, u1_u3_u2_n159, u1_u3_u2_n160, u1_u3_u2_n161, u1_u3_u2_n162, 
       u1_u3_u2_n163, u1_u3_u2_n164, u1_u3_u2_n165, u1_u3_u2_n166, u1_u3_u2_n167, u1_u3_u2_n168, u1_u3_u2_n169, u1_u3_u2_n170, u1_u3_u2_n171, 
       u1_u3_u2_n172, u1_u3_u2_n173, u1_u3_u2_n174, u1_u3_u2_n175, u1_u3_u2_n176, u1_u3_u2_n177, u1_u3_u2_n178, u1_u3_u2_n179, u1_u3_u2_n180, 
       u1_u3_u2_n181, u1_u3_u2_n182, u1_u3_u2_n183, u1_u3_u2_n184, u1_u3_u2_n185, u1_u3_u2_n186, u1_u3_u2_n187, u1_u3_u2_n188, u1_u3_u2_n95, 
       u1_u3_u2_n96, u1_u3_u2_n97, u1_u3_u2_n98, u1_u3_u2_n99, u1_u3_u3_n100, u1_u3_u3_n101, u1_u3_u3_n102, u1_u3_u3_n103, u1_u3_u3_n104, 
       u1_u3_u3_n105, u1_u3_u3_n106, u1_u3_u3_n107, u1_u3_u3_n108, u1_u3_u3_n109, u1_u3_u3_n110, u1_u3_u3_n111, u1_u3_u3_n112, u1_u3_u3_n113, 
       u1_u3_u3_n114, u1_u3_u3_n115, u1_u3_u3_n116, u1_u3_u3_n117, u1_u3_u3_n118, u1_u3_u3_n119, u1_u3_u3_n120, u1_u3_u3_n121, u1_u3_u3_n122, 
       u1_u3_u3_n123, u1_u3_u3_n124, u1_u3_u3_n125, u1_u3_u3_n126, u1_u3_u3_n127, u1_u3_u3_n128, u1_u3_u3_n129, u1_u3_u3_n130, u1_u3_u3_n131, 
       u1_u3_u3_n132, u1_u3_u3_n133, u1_u3_u3_n134, u1_u3_u3_n135, u1_u3_u3_n136, u1_u3_u3_n137, u1_u3_u3_n138, u1_u3_u3_n139, u1_u3_u3_n140, 
       u1_u3_u3_n141, u1_u3_u3_n142, u1_u3_u3_n143, u1_u3_u3_n144, u1_u3_u3_n145, u1_u3_u3_n146, u1_u3_u3_n147, u1_u3_u3_n148, u1_u3_u3_n149, 
       u1_u3_u3_n150, u1_u3_u3_n151, u1_u3_u3_n152, u1_u3_u3_n153, u1_u3_u3_n154, u1_u3_u3_n155, u1_u3_u3_n156, u1_u3_u3_n157, u1_u3_u3_n158, 
       u1_u3_u3_n159, u1_u3_u3_n160, u1_u3_u3_n161, u1_u3_u3_n162, u1_u3_u3_n163, u1_u3_u3_n164, u1_u3_u3_n165, u1_u3_u3_n166, u1_u3_u3_n167, 
       u1_u3_u3_n168, u1_u3_u3_n169, u1_u3_u3_n170, u1_u3_u3_n171, u1_u3_u3_n172, u1_u3_u3_n173, u1_u3_u3_n174, u1_u3_u3_n175, u1_u3_u3_n176, 
       u1_u3_u3_n177, u1_u3_u3_n178, u1_u3_u3_n179, u1_u3_u3_n180, u1_u3_u3_n181, u1_u3_u3_n182, u1_u3_u3_n183, u1_u3_u3_n184, u1_u3_u3_n185, 
       u1_u3_u3_n186, u1_u3_u3_n94, u1_u3_u3_n95, u1_u3_u3_n96, u1_u3_u3_n97, u1_u3_u3_n98, u1_u3_u3_n99, u1_u3_u7_n100, u1_u3_u7_n101, 
       u1_u3_u7_n102, u1_u3_u7_n103, u1_u3_u7_n104, u1_u3_u7_n105, u1_u3_u7_n106, u1_u3_u7_n107, u1_u3_u7_n108, u1_u3_u7_n109, u1_u3_u7_n110, 
       u1_u3_u7_n111, u1_u3_u7_n112, u1_u3_u7_n113, u1_u3_u7_n114, u1_u3_u7_n115, u1_u3_u7_n116, u1_u3_u7_n117, u1_u3_u7_n118, u1_u3_u7_n119, 
       u1_u3_u7_n120, u1_u3_u7_n121, u1_u3_u7_n122, u1_u3_u7_n123, u1_u3_u7_n124, u1_u3_u7_n125, u1_u3_u7_n126, u1_u3_u7_n127, u1_u3_u7_n128, 
       u1_u3_u7_n129, u1_u3_u7_n130, u1_u3_u7_n131, u1_u3_u7_n132, u1_u3_u7_n133, u1_u3_u7_n134, u1_u3_u7_n135, u1_u3_u7_n136, u1_u3_u7_n137, 
       u1_u3_u7_n138, u1_u3_u7_n139, u1_u3_u7_n140, u1_u3_u7_n141, u1_u3_u7_n142, u1_u3_u7_n143, u1_u3_u7_n144, u1_u3_u7_n145, u1_u3_u7_n146, 
       u1_u3_u7_n147, u1_u3_u7_n148, u1_u3_u7_n149, u1_u3_u7_n150, u1_u3_u7_n151, u1_u3_u7_n152, u1_u3_u7_n153, u1_u3_u7_n154, u1_u3_u7_n155, 
       u1_u3_u7_n156, u1_u3_u7_n157, u1_u3_u7_n158, u1_u3_u7_n159, u1_u3_u7_n160, u1_u3_u7_n161, u1_u3_u7_n162, u1_u3_u7_n163, u1_u3_u7_n164, 
       u1_u3_u7_n165, u1_u3_u7_n166, u1_u3_u7_n167, u1_u3_u7_n168, u1_u3_u7_n169, u1_u3_u7_n170, u1_u3_u7_n171, u1_u3_u7_n172, u1_u3_u7_n173, 
       u1_u3_u7_n174, u1_u3_u7_n175, u1_u3_u7_n176, u1_u3_u7_n177, u1_u3_u7_n178, u1_u3_u7_n179, u1_u3_u7_n180, u1_u3_u7_n91, u1_u3_u7_n92, 
       u1_u3_u7_n93, u1_u3_u7_n94, u1_u3_u7_n95, u1_u3_u7_n96, u1_u3_u7_n97, u1_u3_u7_n98, u1_u3_u7_n99, u1_u7_X_43, u1_u7_X_44, 
       u1_u7_X_45, u1_u7_X_46, u1_u7_X_47, u1_u7_X_48, u1_u7_u7_n100, u1_u7_u7_n101, u1_u7_u7_n102, u1_u7_u7_n103, u1_u7_u7_n104, 
       u1_u7_u7_n105, u1_u7_u7_n106, u1_u7_u7_n107, u1_u7_u7_n108, u1_u7_u7_n109, u1_u7_u7_n110, u1_u7_u7_n111, u1_u7_u7_n112, u1_u7_u7_n113, 
       u1_u7_u7_n114, u1_u7_u7_n115, u1_u7_u7_n116, u1_u7_u7_n117, u1_u7_u7_n118, u1_u7_u7_n119, u1_u7_u7_n120, u1_u7_u7_n121, u1_u7_u7_n122, 
       u1_u7_u7_n123, u1_u7_u7_n124, u1_u7_u7_n125, u1_u7_u7_n126, u1_u7_u7_n127, u1_u7_u7_n128, u1_u7_u7_n129, u1_u7_u7_n130, u1_u7_u7_n131, 
       u1_u7_u7_n132, u1_u7_u7_n133, u1_u7_u7_n134, u1_u7_u7_n135, u1_u7_u7_n136, u1_u7_u7_n137, u1_u7_u7_n138, u1_u7_u7_n139, u1_u7_u7_n140, 
       u1_u7_u7_n141, u1_u7_u7_n142, u1_u7_u7_n143, u1_u7_u7_n144, u1_u7_u7_n145, u1_u7_u7_n146, u1_u7_u7_n147, u1_u7_u7_n148, u1_u7_u7_n149, 
       u1_u7_u7_n150, u1_u7_u7_n151, u1_u7_u7_n152, u1_u7_u7_n153, u1_u7_u7_n154, u1_u7_u7_n155, u1_u7_u7_n156, u1_u7_u7_n157, u1_u7_u7_n158, 
       u1_u7_u7_n159, u1_u7_u7_n160, u1_u7_u7_n161, u1_u7_u7_n162, u1_u7_u7_n163, u1_u7_u7_n164, u1_u7_u7_n165, u1_u7_u7_n166, u1_u7_u7_n167, 
       u1_u7_u7_n168, u1_u7_u7_n169, u1_u7_u7_n170, u1_u7_u7_n171, u1_u7_u7_n172, u1_u7_u7_n173, u1_u7_u7_n174, u1_u7_u7_n175, u1_u7_u7_n176, 
       u1_u7_u7_n177, u1_u7_u7_n178, u1_u7_u7_n179, u1_u7_u7_n180, u1_u7_u7_n91, u1_u7_u7_n92, u1_u7_u7_n93, u1_u7_u7_n94, u1_u7_u7_n95, 
       u1_u7_u7_n96, u1_u7_u7_n97, u1_u7_u7_n98, u1_u7_u7_n99, u1_u9_X_31, u1_u9_X_32, u1_u9_X_33, u1_u9_X_34, u1_u9_X_35, 
       u1_u9_X_36, u1_u9_X_37, u1_u9_X_38, u1_u9_X_39, u1_u9_X_40, u1_u9_X_41, u1_u9_X_42, u1_u9_u5_n100, u1_u9_u5_n101, 
       u1_u9_u5_n102, u1_u9_u5_n103, u1_u9_u5_n104, u1_u9_u5_n105, u1_u9_u5_n106, u1_u9_u5_n107, u1_u9_u5_n108, u1_u9_u5_n109, u1_u9_u5_n110, 
       u1_u9_u5_n111, u1_u9_u5_n112, u1_u9_u5_n113, u1_u9_u5_n114, u1_u9_u5_n115, u1_u9_u5_n116, u1_u9_u5_n117, u1_u9_u5_n118, u1_u9_u5_n119, 
       u1_u9_u5_n120, u1_u9_u5_n121, u1_u9_u5_n122, u1_u9_u5_n123, u1_u9_u5_n124, u1_u9_u5_n125, u1_u9_u5_n126, u1_u9_u5_n127, u1_u9_u5_n128, 
       u1_u9_u5_n129, u1_u9_u5_n130, u1_u9_u5_n131, u1_u9_u5_n132, u1_u9_u5_n133, u1_u9_u5_n134, u1_u9_u5_n135, u1_u9_u5_n136, u1_u9_u5_n137, 
       u1_u9_u5_n138, u1_u9_u5_n139, u1_u9_u5_n140, u1_u9_u5_n141, u1_u9_u5_n142, u1_u9_u5_n143, u1_u9_u5_n144, u1_u9_u5_n145, u1_u9_u5_n146, 
       u1_u9_u5_n147, u1_u9_u5_n148, u1_u9_u5_n149, u1_u9_u5_n150, u1_u9_u5_n151, u1_u9_u5_n152, u1_u9_u5_n153, u1_u9_u5_n154, u1_u9_u5_n155, 
       u1_u9_u5_n156, u1_u9_u5_n157, u1_u9_u5_n158, u1_u9_u5_n159, u1_u9_u5_n160, u1_u9_u5_n161, u1_u9_u5_n162, u1_u9_u5_n163, u1_u9_u5_n164, 
       u1_u9_u5_n165, u1_u9_u5_n166, u1_u9_u5_n167, u1_u9_u5_n168, u1_u9_u5_n169, u1_u9_u5_n170, u1_u9_u5_n171, u1_u9_u5_n172, u1_u9_u5_n173, 
       u1_u9_u5_n174, u1_u9_u5_n175, u1_u9_u5_n176, u1_u9_u5_n177, u1_u9_u5_n178, u1_u9_u5_n179, u1_u9_u5_n180, u1_u9_u5_n181, u1_u9_u5_n182, 
       u1_u9_u5_n183, u1_u9_u5_n184, u1_u9_u5_n185, u1_u9_u5_n186, u1_u9_u5_n187, u1_u9_u5_n188, u1_u9_u5_n189, u1_u9_u5_n190, u1_u9_u5_n191, 
       u1_u9_u5_n192, u1_u9_u5_n193, u1_u9_u5_n194, u1_u9_u5_n195, u1_u9_u5_n196, u1_u9_u5_n99, u1_u9_u6_n100, u1_u9_u6_n101, u1_u9_u6_n102, 
       u1_u9_u6_n103, u1_u9_u6_n104, u1_u9_u6_n105, u1_u9_u6_n106, u1_u9_u6_n107, u1_u9_u6_n108, u1_u9_u6_n109, u1_u9_u6_n110, u1_u9_u6_n111, 
       u1_u9_u6_n112, u1_u9_u6_n113, u1_u9_u6_n114, u1_u9_u6_n115, u1_u9_u6_n116, u1_u9_u6_n117, u1_u9_u6_n118, u1_u9_u6_n119, u1_u9_u6_n120, 
       u1_u9_u6_n121, u1_u9_u6_n122, u1_u9_u6_n123, u1_u9_u6_n124, u1_u9_u6_n125, u1_u9_u6_n126, u1_u9_u6_n127, u1_u9_u6_n128, u1_u9_u6_n129, 
       u1_u9_u6_n130, u1_u9_u6_n131, u1_u9_u6_n132, u1_u9_u6_n133, u1_u9_u6_n134, u1_u9_u6_n135, u1_u9_u6_n136, u1_u9_u6_n137, u1_u9_u6_n138, 
       u1_u9_u6_n139, u1_u9_u6_n140, u1_u9_u6_n141, u1_u9_u6_n142, u1_u9_u6_n143, u1_u9_u6_n144, u1_u9_u6_n145, u1_u9_u6_n146, u1_u9_u6_n147, 
       u1_u9_u6_n148, u1_u9_u6_n149, u1_u9_u6_n150, u1_u9_u6_n151, u1_u9_u6_n152, u1_u9_u6_n153, u1_u9_u6_n154, u1_u9_u6_n155, u1_u9_u6_n156, 
       u1_u9_u6_n157, u1_u9_u6_n158, u1_u9_u6_n159, u1_u9_u6_n160, u1_u9_u6_n161, u1_u9_u6_n162, u1_u9_u6_n163, u1_u9_u6_n164, u1_u9_u6_n165, 
       u1_u9_u6_n166, u1_u9_u6_n167, u1_u9_u6_n168, u1_u9_u6_n169, u1_u9_u6_n170, u1_u9_u6_n171, u1_u9_u6_n172, u1_u9_u6_n173, u1_u9_u6_n174, 
       u1_u9_u6_n88, u1_u9_u6_n89, u1_u9_u6_n90, u1_u9_u6_n91, u1_u9_u6_n92, u1_u9_u6_n93, u1_u9_u6_n94, u1_u9_u6_n95, u1_u9_u6_n96, 
       u1_u9_u6_n97, u1_u9_u6_n98, u1_u9_u6_n99, u1_uk_n1051, u1_uk_n1052, u1_uk_n1053, u1_uk_n1054, u1_uk_n1055, u1_uk_n1056, 
       u1_uk_n1061, u1_uk_n1065, u1_uk_n1066, u1_uk_n1067, u1_uk_n1068, u1_uk_n1069, u1_uk_n1143, u1_uk_n1144, u1_uk_n1145, 
       u1_uk_n342, u1_uk_n346, u1_uk_n349, u1_uk_n353, u1_uk_n363, u1_uk_n366, u1_uk_n369, u1_uk_n373, u1_uk_n375, 
       u1_uk_n551, u1_uk_n582, u1_uk_n586, u1_uk_n587, u1_uk_n590, u1_uk_n603, u1_uk_n605, u1_uk_n608, u1_uk_n634, 
       u1_uk_n957, u1_uk_n962, u1_uk_n963, u1_uk_n978, u1_uk_n979, u1_uk_n986, u1_uk_n995, u2_K16_32, u2_K16_33, 
       u2_K16_34, u2_K16_35, u2_K16_36, u2_K16_37, u2_K16_38, u2_K16_39, u2_K16_40, u2_K16_41, u2_K7_25, 
       u2_K7_27, u2_K7_28, u2_K7_29, u2_K7_30, u2_K7_32, u2_K7_34, u2_K7_36, u2_K7_39, u2_K7_40, 
       u2_K7_41, u2_K7_42, u2_K7_44, u2_K7_46, u2_K7_47, u2_out15_11, u2_out15_12, u2_out15_19, u2_out15_22, 
       u2_out15_29, u2_out15_32, u2_out15_4, u2_out15_7, u2_out6_11, u2_out6_12, u2_out6_14, u2_out6_15, u2_out6_19, 
       u2_out6_21, u2_out6_22, u2_out6_25, u2_out6_27, u2_out6_29, u2_out6_3, u2_out6_32, u2_out6_4, u2_out6_5, 
       u2_out6_7, u2_out6_8, u2_u15_X_31, u2_u15_X_32, u2_u15_X_33, u2_u15_X_34, u2_u15_X_35, u2_u15_X_36, u2_u15_X_37, 
       u2_u15_X_38, u2_u15_X_39, u2_u15_X_40, u2_u15_X_41, u2_u15_X_42, u2_u15_u5_n100, u2_u15_u5_n101, u2_u15_u5_n102, u2_u15_u5_n103, 
       u2_u15_u5_n104, u2_u15_u5_n105, u2_u15_u5_n106, u2_u15_u5_n107, u2_u15_u5_n108, u2_u15_u5_n109, u2_u15_u5_n110, u2_u15_u5_n111, u2_u15_u5_n112, 
       u2_u15_u5_n113, u2_u15_u5_n114, u2_u15_u5_n115, u2_u15_u5_n116, u2_u15_u5_n117, u2_u15_u5_n118, u2_u15_u5_n119, u2_u15_u5_n120, u2_u15_u5_n121, 
       u2_u15_u5_n122, u2_u15_u5_n123, u2_u15_u5_n124, u2_u15_u5_n125, u2_u15_u5_n126, u2_u15_u5_n127, u2_u15_u5_n128, u2_u15_u5_n129, u2_u15_u5_n130, 
       u2_u15_u5_n131, u2_u15_u5_n132, u2_u15_u5_n133, u2_u15_u5_n134, u2_u15_u5_n135, u2_u15_u5_n136, u2_u15_u5_n137, u2_u15_u5_n138, u2_u15_u5_n139, 
       u2_u15_u5_n140, u2_u15_u5_n141, u2_u15_u5_n142, u2_u15_u5_n143, u2_u15_u5_n144, u2_u15_u5_n145, u2_u15_u5_n146, u2_u15_u5_n147, u2_u15_u5_n148, 
       u2_u15_u5_n149, u2_u15_u5_n150, u2_u15_u5_n151, u2_u15_u5_n152, u2_u15_u5_n153, u2_u15_u5_n154, u2_u15_u5_n155, u2_u15_u5_n156, u2_u15_u5_n157, 
       u2_u15_u5_n158, u2_u15_u5_n159, u2_u15_u5_n160, u2_u15_u5_n161, u2_u15_u5_n162, u2_u15_u5_n163, u2_u15_u5_n164, u2_u15_u5_n165, u2_u15_u5_n166, 
       u2_u15_u5_n167, u2_u15_u5_n168, u2_u15_u5_n169, u2_u15_u5_n170, u2_u15_u5_n171, u2_u15_u5_n172, u2_u15_u5_n173, u2_u15_u5_n174, u2_u15_u5_n175, 
       u2_u15_u5_n176, u2_u15_u5_n177, u2_u15_u5_n178, u2_u15_u5_n179, u2_u15_u5_n180, u2_u15_u5_n181, u2_u15_u5_n182, u2_u15_u5_n183, u2_u15_u5_n184, 
       u2_u15_u5_n185, u2_u15_u5_n186, u2_u15_u5_n187, u2_u15_u5_n188, u2_u15_u5_n189, u2_u15_u5_n190, u2_u15_u5_n191, u2_u15_u5_n192, u2_u15_u5_n193, 
       u2_u15_u5_n194, u2_u15_u5_n195, u2_u15_u5_n196, u2_u15_u5_n99, u2_u15_u6_n100, u2_u15_u6_n101, u2_u15_u6_n102, u2_u15_u6_n103, u2_u15_u6_n104, 
       u2_u15_u6_n105, u2_u15_u6_n106, u2_u15_u6_n107, u2_u15_u6_n108, u2_u15_u6_n109, u2_u15_u6_n110, u2_u15_u6_n111, u2_u15_u6_n112, u2_u15_u6_n113, 
       u2_u15_u6_n114, u2_u15_u6_n115, u2_u15_u6_n116, u2_u15_u6_n117, u2_u15_u6_n118, u2_u15_u6_n119, u2_u15_u6_n120, u2_u15_u6_n121, u2_u15_u6_n122, 
       u2_u15_u6_n123, u2_u15_u6_n124, u2_u15_u6_n125, u2_u15_u6_n126, u2_u15_u6_n127, u2_u15_u6_n128, u2_u15_u6_n129, u2_u15_u6_n130, u2_u15_u6_n131, 
       u2_u15_u6_n132, u2_u15_u6_n133, u2_u15_u6_n134, u2_u15_u6_n135, u2_u15_u6_n136, u2_u15_u6_n137, u2_u15_u6_n138, u2_u15_u6_n139, u2_u15_u6_n140, 
       u2_u15_u6_n141, u2_u15_u6_n142, u2_u15_u6_n143, u2_u15_u6_n144, u2_u15_u6_n145, u2_u15_u6_n146, u2_u15_u6_n147, u2_u15_u6_n148, u2_u15_u6_n149, 
       u2_u15_u6_n150, u2_u15_u6_n151, u2_u15_u6_n152, u2_u15_u6_n153, u2_u15_u6_n154, u2_u15_u6_n155, u2_u15_u6_n156, u2_u15_u6_n157, u2_u15_u6_n158, 
       u2_u15_u6_n159, u2_u15_u6_n160, u2_u15_u6_n161, u2_u15_u6_n162, u2_u15_u6_n163, u2_u15_u6_n164, u2_u15_u6_n165, u2_u15_u6_n166, u2_u15_u6_n167, 
       u2_u15_u6_n168, u2_u15_u6_n169, u2_u15_u6_n170, u2_u15_u6_n171, u2_u15_u6_n172, u2_u15_u6_n173, u2_u15_u6_n174, u2_u15_u6_n88, u2_u15_u6_n89, 
       u2_u15_u6_n90, u2_u15_u6_n91, u2_u15_u6_n92, u2_u15_u6_n93, u2_u15_u6_n94, u2_u15_u6_n95, u2_u15_u6_n96, u2_u15_u6_n97, u2_u15_u6_n98, 
       u2_u15_u6_n99, u2_u6_X_25, u2_u6_X_26, u2_u6_X_27, u2_u6_X_28, u2_u6_X_29, u2_u6_X_30, u2_u6_X_31, u2_u6_X_32, 
       u2_u6_X_33, u2_u6_X_34, u2_u6_X_35, u2_u6_X_36, u2_u6_X_37, u2_u6_X_38, u2_u6_X_39, u2_u6_X_40, u2_u6_X_41, 
       u2_u6_X_42, u2_u6_X_43, u2_u6_X_44, u2_u6_X_45, u2_u6_X_46, u2_u6_X_47, u2_u6_X_48, u2_u6_u4_n100, u2_u6_u4_n101, 
       u2_u6_u4_n102, u2_u6_u4_n103, u2_u6_u4_n104, u2_u6_u4_n105, u2_u6_u4_n106, u2_u6_u4_n107, u2_u6_u4_n108, u2_u6_u4_n109, u2_u6_u4_n110, 
       u2_u6_u4_n111, u2_u6_u4_n112, u2_u6_u4_n113, u2_u6_u4_n114, u2_u6_u4_n115, u2_u6_u4_n116, u2_u6_u4_n117, u2_u6_u4_n118, u2_u6_u4_n119, 
       u2_u6_u4_n120, u2_u6_u4_n121, u2_u6_u4_n122, u2_u6_u4_n123, u2_u6_u4_n124, u2_u6_u4_n125, u2_u6_u4_n126, u2_u6_u4_n127, u2_u6_u4_n128, 
       u2_u6_u4_n129, u2_u6_u4_n130, u2_u6_u4_n131, u2_u6_u4_n132, u2_u6_u4_n133, u2_u6_u4_n134, u2_u6_u4_n135, u2_u6_u4_n136, u2_u6_u4_n137, 
       u2_u6_u4_n138, u2_u6_u4_n139, u2_u6_u4_n140, u2_u6_u4_n141, u2_u6_u4_n142, u2_u6_u4_n143, u2_u6_u4_n144, u2_u6_u4_n145, u2_u6_u4_n146, 
       u2_u6_u4_n147, u2_u6_u4_n148, u2_u6_u4_n149, u2_u6_u4_n150, u2_u6_u4_n151, u2_u6_u4_n152, u2_u6_u4_n153, u2_u6_u4_n154, u2_u6_u4_n155, 
       u2_u6_u4_n156, u2_u6_u4_n157, u2_u6_u4_n158, u2_u6_u4_n159, u2_u6_u4_n160, u2_u6_u4_n161, u2_u6_u4_n162, u2_u6_u4_n163, u2_u6_u4_n164, 
       u2_u6_u4_n165, u2_u6_u4_n166, u2_u6_u4_n167, u2_u6_u4_n168, u2_u6_u4_n169, u2_u6_u4_n170, u2_u6_u4_n171, u2_u6_u4_n172, u2_u6_u4_n173, 
       u2_u6_u4_n174, u2_u6_u4_n175, u2_u6_u4_n176, u2_u6_u4_n177, u2_u6_u4_n178, u2_u6_u4_n179, u2_u6_u4_n180, u2_u6_u4_n181, u2_u6_u4_n182, 
       u2_u6_u4_n183, u2_u6_u4_n184, u2_u6_u4_n185, u2_u6_u4_n186, u2_u6_u4_n94, u2_u6_u4_n95, u2_u6_u4_n96, u2_u6_u4_n97, u2_u6_u4_n98, 
       u2_u6_u4_n99, u2_u6_u5_n100, u2_u6_u5_n101, u2_u6_u5_n102, u2_u6_u5_n103, u2_u6_u5_n104, u2_u6_u5_n105, u2_u6_u5_n106, u2_u6_u5_n107, 
       u2_u6_u5_n108, u2_u6_u5_n109, u2_u6_u5_n110, u2_u6_u5_n111, u2_u6_u5_n112, u2_u6_u5_n113, u2_u6_u5_n114, u2_u6_u5_n115, u2_u6_u5_n116, 
       u2_u6_u5_n117, u2_u6_u5_n118, u2_u6_u5_n119, u2_u6_u5_n120, u2_u6_u5_n121, u2_u6_u5_n122, u2_u6_u5_n123, u2_u6_u5_n124, u2_u6_u5_n125, 
       u2_u6_u5_n126, u2_u6_u5_n127, u2_u6_u5_n128, u2_u6_u5_n129, u2_u6_u5_n130, u2_u6_u5_n131, u2_u6_u5_n132, u2_u6_u5_n133, u2_u6_u5_n134, 
       u2_u6_u5_n135, u2_u6_u5_n136, u2_u6_u5_n137, u2_u6_u5_n138, u2_u6_u5_n139, u2_u6_u5_n140, u2_u6_u5_n141, u2_u6_u5_n142, u2_u6_u5_n143, 
       u2_u6_u5_n144, u2_u6_u5_n145, u2_u6_u5_n146, u2_u6_u5_n147, u2_u6_u5_n148, u2_u6_u5_n149, u2_u6_u5_n150, u2_u6_u5_n151, u2_u6_u5_n152, 
       u2_u6_u5_n153, u2_u6_u5_n154, u2_u6_u5_n155, u2_u6_u5_n156, u2_u6_u5_n157, u2_u6_u5_n158, u2_u6_u5_n159, u2_u6_u5_n160, u2_u6_u5_n161, 
       u2_u6_u5_n162, u2_u6_u5_n163, u2_u6_u5_n164, u2_u6_u5_n165, u2_u6_u5_n166, u2_u6_u5_n167, u2_u6_u5_n168, u2_u6_u5_n169, u2_u6_u5_n170, 
       u2_u6_u5_n171, u2_u6_u5_n172, u2_u6_u5_n173, u2_u6_u5_n174, u2_u6_u5_n175, u2_u6_u5_n176, u2_u6_u5_n177, u2_u6_u5_n178, u2_u6_u5_n179, 
       u2_u6_u5_n180, u2_u6_u5_n181, u2_u6_u5_n182, u2_u6_u5_n183, u2_u6_u5_n184, u2_u6_u5_n185, u2_u6_u5_n186, u2_u6_u5_n187, u2_u6_u5_n188, 
       u2_u6_u5_n189, u2_u6_u5_n190, u2_u6_u5_n191, u2_u6_u5_n192, u2_u6_u5_n193, u2_u6_u5_n194, u2_u6_u5_n195, u2_u6_u5_n196, u2_u6_u5_n99, 
       u2_u6_u6_n100, u2_u6_u6_n101, u2_u6_u6_n102, u2_u6_u6_n103, u2_u6_u6_n104, u2_u6_u6_n105, u2_u6_u6_n106, u2_u6_u6_n107, u2_u6_u6_n108, 
       u2_u6_u6_n109, u2_u6_u6_n110, u2_u6_u6_n111, u2_u6_u6_n112, u2_u6_u6_n113, u2_u6_u6_n114, u2_u6_u6_n115, u2_u6_u6_n116, u2_u6_u6_n117, 
       u2_u6_u6_n118, u2_u6_u6_n119, u2_u6_u6_n120, u2_u6_u6_n121, u2_u6_u6_n122, u2_u6_u6_n123, u2_u6_u6_n124, u2_u6_u6_n125, u2_u6_u6_n126, 
       u2_u6_u6_n127, u2_u6_u6_n128, u2_u6_u6_n129, u2_u6_u6_n130, u2_u6_u6_n131, u2_u6_u6_n132, u2_u6_u6_n133, u2_u6_u6_n134, u2_u6_u6_n135, 
       u2_u6_u6_n136, u2_u6_u6_n137, u2_u6_u6_n138, u2_u6_u6_n139, u2_u6_u6_n140, u2_u6_u6_n141, u2_u6_u6_n142, u2_u6_u6_n143, u2_u6_u6_n144, 
       u2_u6_u6_n145, u2_u6_u6_n146, u2_u6_u6_n147, u2_u6_u6_n148, u2_u6_u6_n149, u2_u6_u6_n150, u2_u6_u6_n151, u2_u6_u6_n152, u2_u6_u6_n153, 
       u2_u6_u6_n154, u2_u6_u6_n155, u2_u6_u6_n156, u2_u6_u6_n157, u2_u6_u6_n158, u2_u6_u6_n159, u2_u6_u6_n160, u2_u6_u6_n161, u2_u6_u6_n162, 
       u2_u6_u6_n163, u2_u6_u6_n164, u2_u6_u6_n165, u2_u6_u6_n166, u2_u6_u6_n167, u2_u6_u6_n168, u2_u6_u6_n169, u2_u6_u6_n170, u2_u6_u6_n171, 
       u2_u6_u6_n172, u2_u6_u6_n173, u2_u6_u6_n174, u2_u6_u6_n88, u2_u6_u6_n89, u2_u6_u6_n90, u2_u6_u6_n91, u2_u6_u6_n92, u2_u6_u6_n93, 
       u2_u6_u6_n94, u2_u6_u6_n95, u2_u6_u6_n96, u2_u6_u6_n97, u2_u6_u6_n98, u2_u6_u6_n99, u2_u6_u7_n100, u2_u6_u7_n101, u2_u6_u7_n102, 
       u2_u6_u7_n103, u2_u6_u7_n104, u2_u6_u7_n105, u2_u6_u7_n106, u2_u6_u7_n107, u2_u6_u7_n108, u2_u6_u7_n109, u2_u6_u7_n110, u2_u6_u7_n111, 
       u2_u6_u7_n112, u2_u6_u7_n113, u2_u6_u7_n114, u2_u6_u7_n115, u2_u6_u7_n116, u2_u6_u7_n117, u2_u6_u7_n118, u2_u6_u7_n119, u2_u6_u7_n120, 
       u2_u6_u7_n121, u2_u6_u7_n122, u2_u6_u7_n123, u2_u6_u7_n124, u2_u6_u7_n125, u2_u6_u7_n126, u2_u6_u7_n127, u2_u6_u7_n128, u2_u6_u7_n129, 
       u2_u6_u7_n130, u2_u6_u7_n131, u2_u6_u7_n132, u2_u6_u7_n133, u2_u6_u7_n134, u2_u6_u7_n135, u2_u6_u7_n136, u2_u6_u7_n137, u2_u6_u7_n138, 
       u2_u6_u7_n139, u2_u6_u7_n140, u2_u6_u7_n141, u2_u6_u7_n142, u2_u6_u7_n143, u2_u6_u7_n144, u2_u6_u7_n145, u2_u6_u7_n146, u2_u6_u7_n147, 
       u2_u6_u7_n148, u2_u6_u7_n149, u2_u6_u7_n150, u2_u6_u7_n151, u2_u6_u7_n152, u2_u6_u7_n153, u2_u6_u7_n154, u2_u6_u7_n155, u2_u6_u7_n156, 
       u2_u6_u7_n157, u2_u6_u7_n158, u2_u6_u7_n159, u2_u6_u7_n160, u2_u6_u7_n161, u2_u6_u7_n162, u2_u6_u7_n163, u2_u6_u7_n164, u2_u6_u7_n165, 
       u2_u6_u7_n166, u2_u6_u7_n167, u2_u6_u7_n168, u2_u6_u7_n169, u2_u6_u7_n170, u2_u6_u7_n171, u2_u6_u7_n172, u2_u6_u7_n173, u2_u6_u7_n174, 
       u2_u6_u7_n175, u2_u6_u7_n176, u2_u6_u7_n177, u2_u6_u7_n178, u2_u6_u7_n179, u2_u6_u7_n180, u2_u6_u7_n91, u2_u6_u7_n92, u2_u6_u7_n93, 
       u2_u6_u7_n94, u2_u6_u7_n95, u2_u6_u7_n96, u2_u6_u7_n97, u2_u6_u7_n98, u2_u6_u7_n99, u2_uk_n1084, u2_uk_n1085, u2_uk_n1088, 
       u2_uk_n1091, u2_uk_n958, u2_uk_n959,  u2_uk_n960;
  XOR2_X1 u0_U12 (.B( u0_L1_27 ) , .Z( u0_N90 ) , .A( u0_out2_27 ) );
  XOR2_X1 u0_U18 (.B( u0_L1_22 ) , .Z( u0_N85 ) , .A( u0_out2_22 ) );
  XOR2_X1 u0_U19 (.B( u0_L1_21 ) , .Z( u0_N84 ) , .A( u0_out2_21 ) );
  XOR2_X1 u0_U26 (.B( u0_L1_15 ) , .Z( u0_N78 ) , .A( u0_out2_15 ) );
  XOR2_X1 u0_U29 (.B( u0_L1_12 ) , .Z( u0_N75 ) , .A( u0_out2_12 ) );
  XOR2_X1 u0_U34 (.B( u0_L1_7 ) , .Z( u0_N70 ) , .A( u0_out2_7 ) );
  XOR2_X1 u0_U37 (.B( u0_L1_5 ) , .Z( u0_N68 ) , .A( u0_out2_5 ) );
  XOR2_X1 u0_U63 (.B( u0_L13_29 ) , .Z( u0_N476 ) , .A( u0_out14_29 ) );
  XOR2_X1 u0_U7 (.B( u0_L1_32 ) , .Z( u0_N95 ) , .A( u0_out2_32 ) );
  XOR2_X1 u0_U74 (.B( u0_L13_19 ) , .Z( u0_N466 ) , .A( u0_out14_19 ) );
  XOR2_X1 u0_U83 (.B( u0_L13_11 ) , .Z( u0_N458 ) , .A( u0_out14_11 ) );
  XOR2_X1 u0_U90 (.B( u0_L13_4 ) , .Z( u0_N451 ) , .A( u0_out14_4 ) );
  XOR2_X1 u0_u14_U20 (.B( u0_K15_36 ) , .A( u0_R13_25 ) , .Z( u0_u14_X_36 ) );
  XOR2_X1 u0_u14_U21 (.B( u0_K15_35 ) , .A( u0_R13_24 ) , .Z( u0_u14_X_35 ) );
  XOR2_X1 u0_u14_U22 (.B( u0_K15_34 ) , .A( u0_R13_23 ) , .Z( u0_u14_X_34 ) );
  XOR2_X1 u0_u14_U23 (.B( u0_K15_33 ) , .A( u0_R13_22 ) , .Z( u0_u14_X_33 ) );
  XOR2_X1 u0_u14_U24 (.B( u0_K15_32 ) , .A( u0_R13_21 ) , .Z( u0_u14_X_32 ) );
  XOR2_X1 u0_u14_U25 (.B( u0_K15_31 ) , .A( u0_R13_20 ) , .Z( u0_u14_X_31 ) );
  INV_X1 u0_u14_u5_U10 (.A( u0_u14_u5_n121 ) , .ZN( u0_u14_u5_n177 ) );
  NOR3_X1 u0_u14_u5_U100 (.A3( u0_u14_u5_n141 ) , .A1( u0_u14_u5_n142 ) , .ZN( u0_u14_u5_n143 ) , .A2( u0_u14_u5_n191 ) );
  NAND4_X1 u0_u14_u5_U101 (.ZN( u0_out14_4 ) , .A4( u0_u14_u5_n112 ) , .A2( u0_u14_u5_n113 ) , .A1( u0_u14_u5_n114 ) , .A3( u0_u14_u5_n195 ) );
  AOI211_X1 u0_u14_u5_U102 (.A( u0_u14_u5_n110 ) , .C1( u0_u14_u5_n111 ) , .ZN( u0_u14_u5_n112 ) , .B( u0_u14_u5_n118 ) , .C2( u0_u14_u5_n177 ) );
  AOI222_X1 u0_u14_u5_U103 (.ZN( u0_u14_u5_n113 ) , .A1( u0_u14_u5_n131 ) , .C1( u0_u14_u5_n148 ) , .B2( u0_u14_u5_n174 ) , .C2( u0_u14_u5_n178 ) , .A2( u0_u14_u5_n179 ) , .B1( u0_u14_u5_n99 ) );
  NAND3_X1 u0_u14_u5_U104 (.A2( u0_u14_u5_n154 ) , .A3( u0_u14_u5_n158 ) , .A1( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n99 ) );
  NOR2_X1 u0_u14_u5_U11 (.ZN( u0_u14_u5_n160 ) , .A2( u0_u14_u5_n173 ) , .A1( u0_u14_u5_n177 ) );
  INV_X1 u0_u14_u5_U12 (.A( u0_u14_u5_n150 ) , .ZN( u0_u14_u5_n174 ) );
  AOI21_X1 u0_u14_u5_U13 (.A( u0_u14_u5_n160 ) , .B2( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n162 ) , .B1( u0_u14_u5_n192 ) );
  INV_X1 u0_u14_u5_U14 (.A( u0_u14_u5_n159 ) , .ZN( u0_u14_u5_n192 ) );
  AOI21_X1 u0_u14_u5_U15 (.A( u0_u14_u5_n156 ) , .B2( u0_u14_u5_n157 ) , .B1( u0_u14_u5_n158 ) , .ZN( u0_u14_u5_n163 ) );
  AOI21_X1 u0_u14_u5_U16 (.B2( u0_u14_u5_n139 ) , .B1( u0_u14_u5_n140 ) , .ZN( u0_u14_u5_n141 ) , .A( u0_u14_u5_n150 ) );
  OAI21_X1 u0_u14_u5_U17 (.A( u0_u14_u5_n133 ) , .B2( u0_u14_u5_n134 ) , .B1( u0_u14_u5_n135 ) , .ZN( u0_u14_u5_n142 ) );
  OAI21_X1 u0_u14_u5_U18 (.ZN( u0_u14_u5_n133 ) , .B2( u0_u14_u5_n147 ) , .A( u0_u14_u5_n173 ) , .B1( u0_u14_u5_n188 ) );
  NAND2_X1 u0_u14_u5_U19 (.A2( u0_u14_u5_n119 ) , .A1( u0_u14_u5_n123 ) , .ZN( u0_u14_u5_n137 ) );
  INV_X1 u0_u14_u5_U20 (.A( u0_u14_u5_n155 ) , .ZN( u0_u14_u5_n194 ) );
  NAND2_X1 u0_u14_u5_U21 (.A1( u0_u14_u5_n121 ) , .ZN( u0_u14_u5_n132 ) , .A2( u0_u14_u5_n172 ) );
  NAND2_X1 u0_u14_u5_U22 (.A2( u0_u14_u5_n122 ) , .ZN( u0_u14_u5_n136 ) , .A1( u0_u14_u5_n154 ) );
  NAND2_X1 u0_u14_u5_U23 (.A2( u0_u14_u5_n119 ) , .A1( u0_u14_u5_n120 ) , .ZN( u0_u14_u5_n159 ) );
  INV_X1 u0_u14_u5_U24 (.A( u0_u14_u5_n156 ) , .ZN( u0_u14_u5_n175 ) );
  INV_X1 u0_u14_u5_U25 (.A( u0_u14_u5_n158 ) , .ZN( u0_u14_u5_n188 ) );
  INV_X1 u0_u14_u5_U26 (.A( u0_u14_u5_n152 ) , .ZN( u0_u14_u5_n179 ) );
  INV_X1 u0_u14_u5_U27 (.A( u0_u14_u5_n140 ) , .ZN( u0_u14_u5_n182 ) );
  INV_X1 u0_u14_u5_U28 (.A( u0_u14_u5_n151 ) , .ZN( u0_u14_u5_n183 ) );
  INV_X1 u0_u14_u5_U29 (.A( u0_u14_u5_n123 ) , .ZN( u0_u14_u5_n185 ) );
  NOR2_X1 u0_u14_u5_U3 (.ZN( u0_u14_u5_n134 ) , .A1( u0_u14_u5_n183 ) , .A2( u0_u14_u5_n190 ) );
  INV_X1 u0_u14_u5_U30 (.A( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n184 ) );
  INV_X1 u0_u14_u5_U31 (.A( u0_u14_u5_n139 ) , .ZN( u0_u14_u5_n189 ) );
  INV_X1 u0_u14_u5_U32 (.A( u0_u14_u5_n157 ) , .ZN( u0_u14_u5_n190 ) );
  INV_X1 u0_u14_u5_U33 (.A( u0_u14_u5_n120 ) , .ZN( u0_u14_u5_n193 ) );
  NAND2_X1 u0_u14_u5_U34 (.ZN( u0_u14_u5_n111 ) , .A1( u0_u14_u5_n140 ) , .A2( u0_u14_u5_n155 ) );
  INV_X1 u0_u14_u5_U35 (.A( u0_u14_u5_n117 ) , .ZN( u0_u14_u5_n196 ) );
  OAI221_X1 u0_u14_u5_U36 (.A( u0_u14_u5_n116 ) , .ZN( u0_u14_u5_n117 ) , .B2( u0_u14_u5_n119 ) , .C1( u0_u14_u5_n153 ) , .C2( u0_u14_u5_n158 ) , .B1( u0_u14_u5_n172 ) );
  AOI222_X1 u0_u14_u5_U37 (.ZN( u0_u14_u5_n116 ) , .B2( u0_u14_u5_n145 ) , .C1( u0_u14_u5_n148 ) , .A2( u0_u14_u5_n174 ) , .C2( u0_u14_u5_n177 ) , .B1( u0_u14_u5_n187 ) , .A1( u0_u14_u5_n193 ) );
  INV_X1 u0_u14_u5_U38 (.A( u0_u14_u5_n115 ) , .ZN( u0_u14_u5_n187 ) );
  NOR2_X1 u0_u14_u5_U39 (.ZN( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n170 ) , .A2( u0_u14_u5_n180 ) );
  INV_X1 u0_u14_u5_U4 (.A( u0_u14_u5_n138 ) , .ZN( u0_u14_u5_n191 ) );
  AOI22_X1 u0_u14_u5_U40 (.B2( u0_u14_u5_n131 ) , .A2( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n169 ) , .B1( u0_u14_u5_n174 ) , .A1( u0_u14_u5_n185 ) );
  NOR2_X1 u0_u14_u5_U41 (.A1( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n150 ) , .A2( u0_u14_u5_n173 ) );
  AOI21_X1 u0_u14_u5_U42 (.A( u0_u14_u5_n118 ) , .B2( u0_u14_u5_n145 ) , .ZN( u0_u14_u5_n168 ) , .B1( u0_u14_u5_n186 ) );
  INV_X1 u0_u14_u5_U43 (.A( u0_u14_u5_n122 ) , .ZN( u0_u14_u5_n186 ) );
  NOR2_X1 u0_u14_u5_U44 (.A1( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n152 ) , .A2( u0_u14_u5_n176 ) );
  NOR2_X1 u0_u14_u5_U45 (.A1( u0_u14_u5_n115 ) , .ZN( u0_u14_u5_n118 ) , .A2( u0_u14_u5_n153 ) );
  NOR2_X1 u0_u14_u5_U46 (.A2( u0_u14_u5_n145 ) , .ZN( u0_u14_u5_n156 ) , .A1( u0_u14_u5_n174 ) );
  NOR2_X1 u0_u14_u5_U47 (.ZN( u0_u14_u5_n121 ) , .A2( u0_u14_u5_n145 ) , .A1( u0_u14_u5_n176 ) );
  AOI22_X1 u0_u14_u5_U48 (.ZN( u0_u14_u5_n114 ) , .A2( u0_u14_u5_n137 ) , .A1( u0_u14_u5_n145 ) , .B2( u0_u14_u5_n175 ) , .B1( u0_u14_u5_n193 ) );
  OAI211_X1 u0_u14_u5_U49 (.B( u0_u14_u5_n124 ) , .A( u0_u14_u5_n125 ) , .C2( u0_u14_u5_n126 ) , .C1( u0_u14_u5_n127 ) , .ZN( u0_u14_u5_n128 ) );
  OAI21_X1 u0_u14_u5_U5 (.B2( u0_u14_u5_n136 ) , .B1( u0_u14_u5_n137 ) , .ZN( u0_u14_u5_n138 ) , .A( u0_u14_u5_n177 ) );
  NOR3_X1 u0_u14_u5_U50 (.ZN( u0_u14_u5_n127 ) , .A1( u0_u14_u5_n136 ) , .A3( u0_u14_u5_n148 ) , .A2( u0_u14_u5_n182 ) );
  OAI21_X1 u0_u14_u5_U51 (.ZN( u0_u14_u5_n124 ) , .A( u0_u14_u5_n177 ) , .B2( u0_u14_u5_n183 ) , .B1( u0_u14_u5_n189 ) );
  OAI21_X1 u0_u14_u5_U52 (.ZN( u0_u14_u5_n125 ) , .A( u0_u14_u5_n174 ) , .B2( u0_u14_u5_n185 ) , .B1( u0_u14_u5_n190 ) );
  AOI21_X1 u0_u14_u5_U53 (.A( u0_u14_u5_n153 ) , .B2( u0_u14_u5_n154 ) , .B1( u0_u14_u5_n155 ) , .ZN( u0_u14_u5_n164 ) );
  AOI21_X1 u0_u14_u5_U54 (.ZN( u0_u14_u5_n110 ) , .B1( u0_u14_u5_n122 ) , .B2( u0_u14_u5_n139 ) , .A( u0_u14_u5_n153 ) );
  INV_X1 u0_u14_u5_U55 (.A( u0_u14_u5_n153 ) , .ZN( u0_u14_u5_n176 ) );
  INV_X1 u0_u14_u5_U56 (.A( u0_u14_u5_n126 ) , .ZN( u0_u14_u5_n173 ) );
  AND2_X1 u0_u14_u5_U57 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n147 ) );
  AND2_X1 u0_u14_u5_U58 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n148 ) );
  NAND2_X1 u0_u14_u5_U59 (.A1( u0_u14_u5_n105 ) , .A2( u0_u14_u5_n106 ) , .ZN( u0_u14_u5_n158 ) );
  INV_X1 u0_u14_u5_U6 (.A( u0_u14_u5_n135 ) , .ZN( u0_u14_u5_n178 ) );
  NAND2_X1 u0_u14_u5_U60 (.A2( u0_u14_u5_n108 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n139 ) );
  NAND2_X1 u0_u14_u5_U61 (.A1( u0_u14_u5_n106 ) , .A2( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n119 ) );
  NAND2_X1 u0_u14_u5_U62 (.A2( u0_u14_u5_n103 ) , .A1( u0_u14_u5_n105 ) , .ZN( u0_u14_u5_n140 ) );
  NAND2_X1 u0_u14_u5_U63 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n105 ) , .ZN( u0_u14_u5_n155 ) );
  NAND2_X1 u0_u14_u5_U64 (.A2( u0_u14_u5_n106 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n122 ) );
  NAND2_X1 u0_u14_u5_U65 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n106 ) , .ZN( u0_u14_u5_n115 ) );
  NAND2_X1 u0_u14_u5_U66 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n103 ) , .ZN( u0_u14_u5_n161 ) );
  NAND2_X1 u0_u14_u5_U67 (.A1( u0_u14_u5_n105 ) , .A2( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n154 ) );
  INV_X1 u0_u14_u5_U68 (.A( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n172 ) );
  NAND2_X1 u0_u14_u5_U69 (.A1( u0_u14_u5_n103 ) , .A2( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n123 ) );
  OAI22_X1 u0_u14_u5_U7 (.B2( u0_u14_u5_n149 ) , .B1( u0_u14_u5_n150 ) , .A2( u0_u14_u5_n151 ) , .A1( u0_u14_u5_n152 ) , .ZN( u0_u14_u5_n165 ) );
  NAND2_X1 u0_u14_u5_U70 (.A2( u0_u14_u5_n103 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n151 ) );
  NAND2_X1 u0_u14_u5_U71 (.A2( u0_u14_u5_n107 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n120 ) );
  NAND2_X1 u0_u14_u5_U72 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n157 ) );
  AND2_X1 u0_u14_u5_U73 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n104 ) , .ZN( u0_u14_u5_n131 ) );
  INV_X1 u0_u14_u5_U74 (.A( u0_u14_u5_n102 ) , .ZN( u0_u14_u5_n195 ) );
  OAI221_X1 u0_u14_u5_U75 (.A( u0_u14_u5_n101 ) , .ZN( u0_u14_u5_n102 ) , .C2( u0_u14_u5_n115 ) , .C1( u0_u14_u5_n126 ) , .B1( u0_u14_u5_n134 ) , .B2( u0_u14_u5_n160 ) );
  OAI21_X1 u0_u14_u5_U76 (.ZN( u0_u14_u5_n101 ) , .B1( u0_u14_u5_n137 ) , .A( u0_u14_u5_n146 ) , .B2( u0_u14_u5_n147 ) );
  NOR2_X1 u0_u14_u5_U77 (.A2( u0_u14_X_34 ) , .A1( u0_u14_X_35 ) , .ZN( u0_u14_u5_n145 ) );
  NOR2_X1 u0_u14_u5_U78 (.A2( u0_u14_X_34 ) , .ZN( u0_u14_u5_n146 ) , .A1( u0_u14_u5_n171 ) );
  NOR2_X1 u0_u14_u5_U79 (.A2( u0_u14_X_31 ) , .A1( u0_u14_X_32 ) , .ZN( u0_u14_u5_n103 ) );
  NOR3_X1 u0_u14_u5_U8 (.A2( u0_u14_u5_n147 ) , .A1( u0_u14_u5_n148 ) , .ZN( u0_u14_u5_n149 ) , .A3( u0_u14_u5_n194 ) );
  NOR2_X1 u0_u14_u5_U80 (.A2( u0_u14_X_36 ) , .ZN( u0_u14_u5_n105 ) , .A1( u0_u14_u5_n180 ) );
  NOR2_X1 u0_u14_u5_U81 (.A2( u0_u14_X_33 ) , .ZN( u0_u14_u5_n108 ) , .A1( u0_u14_u5_n170 ) );
  NOR2_X1 u0_u14_u5_U82 (.A2( u0_u14_X_33 ) , .A1( u0_u14_X_36 ) , .ZN( u0_u14_u5_n107 ) );
  NOR2_X1 u0_u14_u5_U83 (.A2( u0_u14_X_31 ) , .ZN( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n181 ) );
  NAND2_X1 u0_u14_u5_U84 (.A2( u0_u14_X_34 ) , .A1( u0_u14_X_35 ) , .ZN( u0_u14_u5_n153 ) );
  NAND2_X1 u0_u14_u5_U85 (.A1( u0_u14_X_34 ) , .ZN( u0_u14_u5_n126 ) , .A2( u0_u14_u5_n171 ) );
  AND2_X1 u0_u14_u5_U86 (.A1( u0_u14_X_31 ) , .A2( u0_u14_X_32 ) , .ZN( u0_u14_u5_n106 ) );
  AND2_X1 u0_u14_u5_U87 (.A1( u0_u14_X_31 ) , .ZN( u0_u14_u5_n109 ) , .A2( u0_u14_u5_n181 ) );
  INV_X1 u0_u14_u5_U88 (.A( u0_u14_X_33 ) , .ZN( u0_u14_u5_n180 ) );
  INV_X1 u0_u14_u5_U89 (.A( u0_u14_X_35 ) , .ZN( u0_u14_u5_n171 ) );
  NOR2_X1 u0_u14_u5_U9 (.ZN( u0_u14_u5_n135 ) , .A1( u0_u14_u5_n173 ) , .A2( u0_u14_u5_n176 ) );
  INV_X1 u0_u14_u5_U90 (.A( u0_u14_X_36 ) , .ZN( u0_u14_u5_n170 ) );
  INV_X1 u0_u14_u5_U91 (.A( u0_u14_X_32 ) , .ZN( u0_u14_u5_n181 ) );
  NAND4_X1 u0_u14_u5_U92 (.ZN( u0_out14_29 ) , .A4( u0_u14_u5_n129 ) , .A3( u0_u14_u5_n130 ) , .A2( u0_u14_u5_n168 ) , .A1( u0_u14_u5_n196 ) );
  AOI221_X1 u0_u14_u5_U93 (.A( u0_u14_u5_n128 ) , .ZN( u0_u14_u5_n129 ) , .C2( u0_u14_u5_n132 ) , .B2( u0_u14_u5_n159 ) , .B1( u0_u14_u5_n176 ) , .C1( u0_u14_u5_n184 ) );
  AOI222_X1 u0_u14_u5_U94 (.ZN( u0_u14_u5_n130 ) , .A2( u0_u14_u5_n146 ) , .B1( u0_u14_u5_n147 ) , .C2( u0_u14_u5_n175 ) , .B2( u0_u14_u5_n179 ) , .A1( u0_u14_u5_n188 ) , .C1( u0_u14_u5_n194 ) );
  NAND4_X1 u0_u14_u5_U95 (.ZN( u0_out14_19 ) , .A4( u0_u14_u5_n166 ) , .A3( u0_u14_u5_n167 ) , .A2( u0_u14_u5_n168 ) , .A1( u0_u14_u5_n169 ) );
  AOI22_X1 u0_u14_u5_U96 (.B2( u0_u14_u5_n145 ) , .A2( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n167 ) , .B1( u0_u14_u5_n182 ) , .A1( u0_u14_u5_n189 ) );
  NOR4_X1 u0_u14_u5_U97 (.A4( u0_u14_u5_n162 ) , .A3( u0_u14_u5_n163 ) , .A2( u0_u14_u5_n164 ) , .A1( u0_u14_u5_n165 ) , .ZN( u0_u14_u5_n166 ) );
  NAND4_X1 u0_u14_u5_U98 (.ZN( u0_out14_11 ) , .A4( u0_u14_u5_n143 ) , .A3( u0_u14_u5_n144 ) , .A2( u0_u14_u5_n169 ) , .A1( u0_u14_u5_n196 ) );
  AOI22_X1 u0_u14_u5_U99 (.A2( u0_u14_u5_n132 ) , .ZN( u0_u14_u5_n144 ) , .B2( u0_u14_u5_n145 ) , .B1( u0_u14_u5_n184 ) , .A1( u0_u14_u5_n194 ) );
  XOR2_X1 u0_u2_U10 (.B( u0_K3_45 ) , .A( u0_R1_30 ) , .Z( u0_u2_X_45 ) );
  XOR2_X1 u0_u2_U11 (.B( u0_K3_44 ) , .A( u0_R1_29 ) , .Z( u0_u2_X_44 ) );
  XOR2_X1 u0_u2_U12 (.B( u0_K3_43 ) , .A( u0_R1_28 ) , .Z( u0_u2_X_43 ) );
  XOR2_X1 u0_u2_U13 (.B( u0_K3_42 ) , .A( u0_R1_29 ) , .Z( u0_u2_X_42 ) );
  XOR2_X1 u0_u2_U14 (.B( u0_K3_41 ) , .A( u0_R1_28 ) , .Z( u0_u2_X_41 ) );
  XOR2_X1 u0_u2_U15 (.B( u0_K3_40 ) , .A( u0_R1_27 ) , .Z( u0_u2_X_40 ) );
  XOR2_X1 u0_u2_U17 (.B( u0_K3_39 ) , .A( u0_R1_26 ) , .Z( u0_u2_X_39 ) );
  XOR2_X1 u0_u2_U18 (.B( u0_K3_38 ) , .A( u0_R1_25 ) , .Z( u0_u2_X_38 ) );
  XOR2_X1 u0_u2_U19 (.B( u0_K3_37 ) , .A( u0_R1_24 ) , .Z( u0_u2_X_37 ) );
  XOR2_X1 u0_u2_U7 (.B( u0_K3_48 ) , .A( u0_R1_1 ) , .Z( u0_u2_X_48 ) );
  XOR2_X1 u0_u2_U8 (.B( u0_K3_47 ) , .A( u0_R1_32 ) , .Z( u0_u2_X_47 ) );
  XOR2_X1 u0_u2_U9 (.B( u0_K3_46 ) , .A( u0_R1_31 ) , .Z( u0_u2_X_46 ) );
  OAI21_X1 u0_u2_u6_U10 (.A( u0_u2_u6_n159 ) , .B1( u0_u2_u6_n169 ) , .B2( u0_u2_u6_n173 ) , .ZN( u0_u2_u6_n90 ) );
  INV_X1 u0_u2_u6_U11 (.ZN( u0_u2_u6_n172 ) , .A( u0_u2_u6_n88 ) );
  AOI22_X1 u0_u2_u6_U12 (.A2( u0_u2_u6_n151 ) , .B2( u0_u2_u6_n161 ) , .A1( u0_u2_u6_n167 ) , .B1( u0_u2_u6_n170 ) , .ZN( u0_u2_u6_n89 ) );
  AOI21_X1 u0_u2_u6_U13 (.ZN( u0_u2_u6_n106 ) , .A( u0_u2_u6_n142 ) , .B2( u0_u2_u6_n159 ) , .B1( u0_u2_u6_n164 ) );
  INV_X1 u0_u2_u6_U14 (.A( u0_u2_u6_n155 ) , .ZN( u0_u2_u6_n161 ) );
  INV_X1 u0_u2_u6_U15 (.A( u0_u2_u6_n128 ) , .ZN( u0_u2_u6_n164 ) );
  NAND2_X1 u0_u2_u6_U16 (.ZN( u0_u2_u6_n110 ) , .A1( u0_u2_u6_n122 ) , .A2( u0_u2_u6_n129 ) );
  NAND2_X1 u0_u2_u6_U17 (.ZN( u0_u2_u6_n124 ) , .A2( u0_u2_u6_n146 ) , .A1( u0_u2_u6_n148 ) );
  INV_X1 u0_u2_u6_U18 (.A( u0_u2_u6_n132 ) , .ZN( u0_u2_u6_n171 ) );
  AND2_X1 u0_u2_u6_U19 (.A1( u0_u2_u6_n100 ) , .ZN( u0_u2_u6_n130 ) , .A2( u0_u2_u6_n147 ) );
  INV_X1 u0_u2_u6_U20 (.A( u0_u2_u6_n127 ) , .ZN( u0_u2_u6_n173 ) );
  INV_X1 u0_u2_u6_U21 (.A( u0_u2_u6_n121 ) , .ZN( u0_u2_u6_n167 ) );
  INV_X1 u0_u2_u6_U22 (.A( u0_u2_u6_n100 ) , .ZN( u0_u2_u6_n169 ) );
  INV_X1 u0_u2_u6_U23 (.A( u0_u2_u6_n123 ) , .ZN( u0_u2_u6_n170 ) );
  INV_X1 u0_u2_u6_U24 (.A( u0_u2_u6_n113 ) , .ZN( u0_u2_u6_n168 ) );
  AND2_X1 u0_u2_u6_U25 (.A1( u0_u2_u6_n107 ) , .A2( u0_u2_u6_n119 ) , .ZN( u0_u2_u6_n133 ) );
  AND2_X1 u0_u2_u6_U26 (.A2( u0_u2_u6_n121 ) , .A1( u0_u2_u6_n122 ) , .ZN( u0_u2_u6_n131 ) );
  AND3_X1 u0_u2_u6_U27 (.ZN( u0_u2_u6_n120 ) , .A2( u0_u2_u6_n127 ) , .A1( u0_u2_u6_n132 ) , .A3( u0_u2_u6_n145 ) );
  INV_X1 u0_u2_u6_U28 (.A( u0_u2_u6_n146 ) , .ZN( u0_u2_u6_n163 ) );
  AOI222_X1 u0_u2_u6_U29 (.ZN( u0_u2_u6_n114 ) , .A1( u0_u2_u6_n118 ) , .A2( u0_u2_u6_n126 ) , .B2( u0_u2_u6_n151 ) , .C2( u0_u2_u6_n159 ) , .C1( u0_u2_u6_n168 ) , .B1( u0_u2_u6_n169 ) );
  INV_X1 u0_u2_u6_U3 (.A( u0_u2_u6_n110 ) , .ZN( u0_u2_u6_n166 ) );
  NOR2_X1 u0_u2_u6_U30 (.A1( u0_u2_u6_n162 ) , .A2( u0_u2_u6_n165 ) , .ZN( u0_u2_u6_n98 ) );
  NAND2_X1 u0_u2_u6_U31 (.A1( u0_u2_u6_n144 ) , .ZN( u0_u2_u6_n151 ) , .A2( u0_u2_u6_n158 ) );
  NAND2_X1 u0_u2_u6_U32 (.ZN( u0_u2_u6_n132 ) , .A1( u0_u2_u6_n91 ) , .A2( u0_u2_u6_n97 ) );
  AOI22_X1 u0_u2_u6_U33 (.B2( u0_u2_u6_n110 ) , .B1( u0_u2_u6_n111 ) , .A1( u0_u2_u6_n112 ) , .ZN( u0_u2_u6_n115 ) , .A2( u0_u2_u6_n161 ) );
  NAND4_X1 u0_u2_u6_U34 (.A3( u0_u2_u6_n109 ) , .ZN( u0_u2_u6_n112 ) , .A4( u0_u2_u6_n132 ) , .A2( u0_u2_u6_n147 ) , .A1( u0_u2_u6_n166 ) );
  NOR2_X1 u0_u2_u6_U35 (.ZN( u0_u2_u6_n109 ) , .A1( u0_u2_u6_n170 ) , .A2( u0_u2_u6_n173 ) );
  NOR2_X1 u0_u2_u6_U36 (.A2( u0_u2_u6_n126 ) , .ZN( u0_u2_u6_n155 ) , .A1( u0_u2_u6_n160 ) );
  NAND2_X1 u0_u2_u6_U37 (.ZN( u0_u2_u6_n146 ) , .A2( u0_u2_u6_n94 ) , .A1( u0_u2_u6_n99 ) );
  AOI21_X1 u0_u2_u6_U38 (.A( u0_u2_u6_n144 ) , .B2( u0_u2_u6_n145 ) , .B1( u0_u2_u6_n146 ) , .ZN( u0_u2_u6_n150 ) );
  INV_X1 u0_u2_u6_U39 (.A( u0_u2_u6_n111 ) , .ZN( u0_u2_u6_n158 ) );
  INV_X1 u0_u2_u6_U4 (.A( u0_u2_u6_n142 ) , .ZN( u0_u2_u6_n174 ) );
  NAND2_X1 u0_u2_u6_U40 (.ZN( u0_u2_u6_n127 ) , .A1( u0_u2_u6_n91 ) , .A2( u0_u2_u6_n92 ) );
  NAND2_X1 u0_u2_u6_U41 (.ZN( u0_u2_u6_n129 ) , .A2( u0_u2_u6_n95 ) , .A1( u0_u2_u6_n96 ) );
  INV_X1 u0_u2_u6_U42 (.A( u0_u2_u6_n144 ) , .ZN( u0_u2_u6_n159 ) );
  NAND2_X1 u0_u2_u6_U43 (.ZN( u0_u2_u6_n145 ) , .A2( u0_u2_u6_n97 ) , .A1( u0_u2_u6_n98 ) );
  NAND2_X1 u0_u2_u6_U44 (.ZN( u0_u2_u6_n148 ) , .A2( u0_u2_u6_n92 ) , .A1( u0_u2_u6_n94 ) );
  NAND2_X1 u0_u2_u6_U45 (.ZN( u0_u2_u6_n108 ) , .A2( u0_u2_u6_n139 ) , .A1( u0_u2_u6_n144 ) );
  NAND2_X1 u0_u2_u6_U46 (.ZN( u0_u2_u6_n121 ) , .A2( u0_u2_u6_n95 ) , .A1( u0_u2_u6_n97 ) );
  NAND2_X1 u0_u2_u6_U47 (.ZN( u0_u2_u6_n107 ) , .A2( u0_u2_u6_n92 ) , .A1( u0_u2_u6_n95 ) );
  AND2_X1 u0_u2_u6_U48 (.ZN( u0_u2_u6_n118 ) , .A2( u0_u2_u6_n91 ) , .A1( u0_u2_u6_n99 ) );
  NAND2_X1 u0_u2_u6_U49 (.ZN( u0_u2_u6_n147 ) , .A2( u0_u2_u6_n98 ) , .A1( u0_u2_u6_n99 ) );
  NAND2_X1 u0_u2_u6_U5 (.A2( u0_u2_u6_n143 ) , .ZN( u0_u2_u6_n152 ) , .A1( u0_u2_u6_n166 ) );
  NAND2_X1 u0_u2_u6_U50 (.ZN( u0_u2_u6_n128 ) , .A1( u0_u2_u6_n94 ) , .A2( u0_u2_u6_n96 ) );
  AOI211_X1 u0_u2_u6_U51 (.B( u0_u2_u6_n134 ) , .A( u0_u2_u6_n135 ) , .C1( u0_u2_u6_n136 ) , .ZN( u0_u2_u6_n137 ) , .C2( u0_u2_u6_n151 ) );
  AOI21_X1 u0_u2_u6_U52 (.B2( u0_u2_u6_n132 ) , .B1( u0_u2_u6_n133 ) , .ZN( u0_u2_u6_n134 ) , .A( u0_u2_u6_n158 ) );
  AOI21_X1 u0_u2_u6_U53 (.B1( u0_u2_u6_n131 ) , .ZN( u0_u2_u6_n135 ) , .A( u0_u2_u6_n144 ) , .B2( u0_u2_u6_n146 ) );
  NAND4_X1 u0_u2_u6_U54 (.A4( u0_u2_u6_n127 ) , .A3( u0_u2_u6_n128 ) , .A2( u0_u2_u6_n129 ) , .A1( u0_u2_u6_n130 ) , .ZN( u0_u2_u6_n136 ) );
  NAND2_X1 u0_u2_u6_U55 (.ZN( u0_u2_u6_n119 ) , .A2( u0_u2_u6_n95 ) , .A1( u0_u2_u6_n99 ) );
  NAND2_X1 u0_u2_u6_U56 (.ZN( u0_u2_u6_n123 ) , .A2( u0_u2_u6_n91 ) , .A1( u0_u2_u6_n96 ) );
  NAND2_X1 u0_u2_u6_U57 (.ZN( u0_u2_u6_n100 ) , .A2( u0_u2_u6_n92 ) , .A1( u0_u2_u6_n98 ) );
  NAND2_X1 u0_u2_u6_U58 (.ZN( u0_u2_u6_n122 ) , .A1( u0_u2_u6_n94 ) , .A2( u0_u2_u6_n97 ) );
  INV_X1 u0_u2_u6_U59 (.A( u0_u2_u6_n139 ) , .ZN( u0_u2_u6_n160 ) );
  AOI22_X1 u0_u2_u6_U6 (.B2( u0_u2_u6_n101 ) , .A1( u0_u2_u6_n102 ) , .ZN( u0_u2_u6_n103 ) , .B1( u0_u2_u6_n160 ) , .A2( u0_u2_u6_n161 ) );
  NAND2_X1 u0_u2_u6_U60 (.ZN( u0_u2_u6_n113 ) , .A1( u0_u2_u6_n96 ) , .A2( u0_u2_u6_n98 ) );
  NOR2_X1 u0_u2_u6_U61 (.A2( u0_u2_X_40 ) , .A1( u0_u2_X_41 ) , .ZN( u0_u2_u6_n126 ) );
  NOR2_X1 u0_u2_u6_U62 (.A2( u0_u2_X_39 ) , .A1( u0_u2_X_42 ) , .ZN( u0_u2_u6_n92 ) );
  NOR2_X1 u0_u2_u6_U63 (.A2( u0_u2_X_39 ) , .A1( u0_u2_u6_n156 ) , .ZN( u0_u2_u6_n97 ) );
  NOR2_X1 u0_u2_u6_U64 (.A2( u0_u2_X_38 ) , .A1( u0_u2_u6_n165 ) , .ZN( u0_u2_u6_n95 ) );
  NOR2_X1 u0_u2_u6_U65 (.A2( u0_u2_X_41 ) , .ZN( u0_u2_u6_n111 ) , .A1( u0_u2_u6_n157 ) );
  NOR2_X1 u0_u2_u6_U66 (.A2( u0_u2_X_37 ) , .A1( u0_u2_u6_n162 ) , .ZN( u0_u2_u6_n94 ) );
  NOR2_X1 u0_u2_u6_U67 (.A2( u0_u2_X_37 ) , .A1( u0_u2_X_38 ) , .ZN( u0_u2_u6_n91 ) );
  NAND2_X1 u0_u2_u6_U68 (.A1( u0_u2_X_41 ) , .ZN( u0_u2_u6_n144 ) , .A2( u0_u2_u6_n157 ) );
  NAND2_X1 u0_u2_u6_U69 (.A2( u0_u2_X_40 ) , .A1( u0_u2_X_41 ) , .ZN( u0_u2_u6_n139 ) );
  NOR2_X1 u0_u2_u6_U7 (.A1( u0_u2_u6_n118 ) , .ZN( u0_u2_u6_n143 ) , .A2( u0_u2_u6_n168 ) );
  AND2_X1 u0_u2_u6_U70 (.A1( u0_u2_X_39 ) , .A2( u0_u2_u6_n156 ) , .ZN( u0_u2_u6_n96 ) );
  AND2_X1 u0_u2_u6_U71 (.A1( u0_u2_X_39 ) , .A2( u0_u2_X_42 ) , .ZN( u0_u2_u6_n99 ) );
  INV_X1 u0_u2_u6_U72 (.A( u0_u2_X_40 ) , .ZN( u0_u2_u6_n157 ) );
  INV_X1 u0_u2_u6_U73 (.A( u0_u2_X_37 ) , .ZN( u0_u2_u6_n165 ) );
  INV_X1 u0_u2_u6_U74 (.A( u0_u2_X_38 ) , .ZN( u0_u2_u6_n162 ) );
  INV_X1 u0_u2_u6_U75 (.A( u0_u2_X_42 ) , .ZN( u0_u2_u6_n156 ) );
  NAND4_X1 u0_u2_u6_U76 (.ZN( u0_out2_32 ) , .A4( u0_u2_u6_n103 ) , .A3( u0_u2_u6_n104 ) , .A2( u0_u2_u6_n105 ) , .A1( u0_u2_u6_n106 ) );
  AOI22_X1 u0_u2_u6_U77 (.ZN( u0_u2_u6_n105 ) , .A2( u0_u2_u6_n108 ) , .A1( u0_u2_u6_n118 ) , .B2( u0_u2_u6_n126 ) , .B1( u0_u2_u6_n171 ) );
  AOI22_X1 u0_u2_u6_U78 (.ZN( u0_u2_u6_n104 ) , .A1( u0_u2_u6_n111 ) , .B1( u0_u2_u6_n124 ) , .B2( u0_u2_u6_n151 ) , .A2( u0_u2_u6_n93 ) );
  NAND4_X1 u0_u2_u6_U79 (.ZN( u0_out2_12 ) , .A4( u0_u2_u6_n114 ) , .A3( u0_u2_u6_n115 ) , .A2( u0_u2_u6_n116 ) , .A1( u0_u2_u6_n117 ) );
  AOI21_X1 u0_u2_u6_U8 (.B1( u0_u2_u6_n107 ) , .B2( u0_u2_u6_n132 ) , .A( u0_u2_u6_n158 ) , .ZN( u0_u2_u6_n88 ) );
  OAI22_X1 u0_u2_u6_U80 (.B2( u0_u2_u6_n111 ) , .ZN( u0_u2_u6_n116 ) , .B1( u0_u2_u6_n126 ) , .A2( u0_u2_u6_n164 ) , .A1( u0_u2_u6_n167 ) );
  OAI21_X1 u0_u2_u6_U81 (.A( u0_u2_u6_n108 ) , .ZN( u0_u2_u6_n117 ) , .B2( u0_u2_u6_n141 ) , .B1( u0_u2_u6_n163 ) );
  OAI211_X1 u0_u2_u6_U82 (.ZN( u0_out2_7 ) , .B( u0_u2_u6_n153 ) , .C2( u0_u2_u6_n154 ) , .C1( u0_u2_u6_n155 ) , .A( u0_u2_u6_n174 ) );
  NOR3_X1 u0_u2_u6_U83 (.A1( u0_u2_u6_n141 ) , .ZN( u0_u2_u6_n154 ) , .A3( u0_u2_u6_n164 ) , .A2( u0_u2_u6_n171 ) );
  AOI211_X1 u0_u2_u6_U84 (.B( u0_u2_u6_n149 ) , .A( u0_u2_u6_n150 ) , .C2( u0_u2_u6_n151 ) , .C1( u0_u2_u6_n152 ) , .ZN( u0_u2_u6_n153 ) );
  OAI211_X1 u0_u2_u6_U85 (.ZN( u0_out2_22 ) , .B( u0_u2_u6_n137 ) , .A( u0_u2_u6_n138 ) , .C2( u0_u2_u6_n139 ) , .C1( u0_u2_u6_n140 ) );
  AOI22_X1 u0_u2_u6_U86 (.B1( u0_u2_u6_n124 ) , .A2( u0_u2_u6_n125 ) , .A1( u0_u2_u6_n126 ) , .ZN( u0_u2_u6_n138 ) , .B2( u0_u2_u6_n161 ) );
  AND4_X1 u0_u2_u6_U87 (.A3( u0_u2_u6_n119 ) , .A1( u0_u2_u6_n120 ) , .A4( u0_u2_u6_n129 ) , .ZN( u0_u2_u6_n140 ) , .A2( u0_u2_u6_n143 ) );
  NAND3_X1 u0_u2_u6_U88 (.A2( u0_u2_u6_n123 ) , .ZN( u0_u2_u6_n125 ) , .A1( u0_u2_u6_n130 ) , .A3( u0_u2_u6_n131 ) );
  NAND3_X1 u0_u2_u6_U89 (.A3( u0_u2_u6_n133 ) , .ZN( u0_u2_u6_n141 ) , .A1( u0_u2_u6_n145 ) , .A2( u0_u2_u6_n148 ) );
  AOI21_X1 u0_u2_u6_U9 (.B2( u0_u2_u6_n147 ) , .B1( u0_u2_u6_n148 ) , .ZN( u0_u2_u6_n149 ) , .A( u0_u2_u6_n158 ) );
  NAND3_X1 u0_u2_u6_U90 (.ZN( u0_u2_u6_n101 ) , .A3( u0_u2_u6_n107 ) , .A2( u0_u2_u6_n121 ) , .A1( u0_u2_u6_n127 ) );
  NAND3_X1 u0_u2_u6_U91 (.ZN( u0_u2_u6_n102 ) , .A3( u0_u2_u6_n130 ) , .A2( u0_u2_u6_n145 ) , .A1( u0_u2_u6_n166 ) );
  NAND3_X1 u0_u2_u6_U92 (.A3( u0_u2_u6_n113 ) , .A1( u0_u2_u6_n119 ) , .A2( u0_u2_u6_n123 ) , .ZN( u0_u2_u6_n93 ) );
  NAND3_X1 u0_u2_u6_U93 (.ZN( u0_u2_u6_n142 ) , .A2( u0_u2_u6_n172 ) , .A3( u0_u2_u6_n89 ) , .A1( u0_u2_u6_n90 ) );
  AND3_X1 u0_u2_u7_U10 (.A3( u0_u2_u7_n110 ) , .A2( u0_u2_u7_n127 ) , .A1( u0_u2_u7_n132 ) , .ZN( u0_u2_u7_n92 ) );
  OAI21_X1 u0_u2_u7_U11 (.A( u0_u2_u7_n161 ) , .B1( u0_u2_u7_n168 ) , .B2( u0_u2_u7_n173 ) , .ZN( u0_u2_u7_n91 ) );
  AOI211_X1 u0_u2_u7_U12 (.A( u0_u2_u7_n117 ) , .ZN( u0_u2_u7_n118 ) , .C2( u0_u2_u7_n126 ) , .C1( u0_u2_u7_n177 ) , .B( u0_u2_u7_n180 ) );
  OAI22_X1 u0_u2_u7_U13 (.B1( u0_u2_u7_n115 ) , .ZN( u0_u2_u7_n117 ) , .A2( u0_u2_u7_n133 ) , .A1( u0_u2_u7_n137 ) , .B2( u0_u2_u7_n162 ) );
  INV_X1 u0_u2_u7_U14 (.A( u0_u2_u7_n116 ) , .ZN( u0_u2_u7_n180 ) );
  NOR3_X1 u0_u2_u7_U15 (.ZN( u0_u2_u7_n115 ) , .A3( u0_u2_u7_n145 ) , .A2( u0_u2_u7_n168 ) , .A1( u0_u2_u7_n169 ) );
  OAI211_X1 u0_u2_u7_U16 (.B( u0_u2_u7_n122 ) , .A( u0_u2_u7_n123 ) , .C2( u0_u2_u7_n124 ) , .ZN( u0_u2_u7_n154 ) , .C1( u0_u2_u7_n162 ) );
  AOI222_X1 u0_u2_u7_U17 (.ZN( u0_u2_u7_n122 ) , .C2( u0_u2_u7_n126 ) , .C1( u0_u2_u7_n145 ) , .B1( u0_u2_u7_n161 ) , .A2( u0_u2_u7_n165 ) , .B2( u0_u2_u7_n170 ) , .A1( u0_u2_u7_n176 ) );
  INV_X1 u0_u2_u7_U18 (.A( u0_u2_u7_n133 ) , .ZN( u0_u2_u7_n176 ) );
  NOR3_X1 u0_u2_u7_U19 (.A2( u0_u2_u7_n134 ) , .A1( u0_u2_u7_n135 ) , .ZN( u0_u2_u7_n136 ) , .A3( u0_u2_u7_n171 ) );
  NOR2_X1 u0_u2_u7_U20 (.A1( u0_u2_u7_n130 ) , .A2( u0_u2_u7_n134 ) , .ZN( u0_u2_u7_n153 ) );
  INV_X1 u0_u2_u7_U21 (.A( u0_u2_u7_n101 ) , .ZN( u0_u2_u7_n165 ) );
  NOR2_X1 u0_u2_u7_U22 (.ZN( u0_u2_u7_n111 ) , .A2( u0_u2_u7_n134 ) , .A1( u0_u2_u7_n169 ) );
  AOI21_X1 u0_u2_u7_U23 (.ZN( u0_u2_u7_n104 ) , .B2( u0_u2_u7_n112 ) , .B1( u0_u2_u7_n127 ) , .A( u0_u2_u7_n164 ) );
  AOI21_X1 u0_u2_u7_U24 (.ZN( u0_u2_u7_n106 ) , .B1( u0_u2_u7_n133 ) , .B2( u0_u2_u7_n146 ) , .A( u0_u2_u7_n162 ) );
  AOI21_X1 u0_u2_u7_U25 (.A( u0_u2_u7_n101 ) , .ZN( u0_u2_u7_n107 ) , .B2( u0_u2_u7_n128 ) , .B1( u0_u2_u7_n175 ) );
  INV_X1 u0_u2_u7_U26 (.A( u0_u2_u7_n138 ) , .ZN( u0_u2_u7_n171 ) );
  INV_X1 u0_u2_u7_U27 (.A( u0_u2_u7_n131 ) , .ZN( u0_u2_u7_n177 ) );
  INV_X1 u0_u2_u7_U28 (.A( u0_u2_u7_n110 ) , .ZN( u0_u2_u7_n174 ) );
  NAND2_X1 u0_u2_u7_U29 (.A1( u0_u2_u7_n129 ) , .A2( u0_u2_u7_n132 ) , .ZN( u0_u2_u7_n149 ) );
  OAI21_X1 u0_u2_u7_U3 (.ZN( u0_u2_u7_n159 ) , .A( u0_u2_u7_n165 ) , .B2( u0_u2_u7_n171 ) , .B1( u0_u2_u7_n174 ) );
  NAND2_X1 u0_u2_u7_U30 (.A1( u0_u2_u7_n113 ) , .A2( u0_u2_u7_n124 ) , .ZN( u0_u2_u7_n130 ) );
  INV_X1 u0_u2_u7_U31 (.A( u0_u2_u7_n112 ) , .ZN( u0_u2_u7_n173 ) );
  INV_X1 u0_u2_u7_U32 (.A( u0_u2_u7_n128 ) , .ZN( u0_u2_u7_n168 ) );
  INV_X1 u0_u2_u7_U33 (.A( u0_u2_u7_n148 ) , .ZN( u0_u2_u7_n169 ) );
  INV_X1 u0_u2_u7_U34 (.A( u0_u2_u7_n127 ) , .ZN( u0_u2_u7_n179 ) );
  NOR2_X1 u0_u2_u7_U35 (.ZN( u0_u2_u7_n101 ) , .A2( u0_u2_u7_n150 ) , .A1( u0_u2_u7_n156 ) );
  AOI211_X1 u0_u2_u7_U36 (.B( u0_u2_u7_n154 ) , .A( u0_u2_u7_n155 ) , .C1( u0_u2_u7_n156 ) , .ZN( u0_u2_u7_n157 ) , .C2( u0_u2_u7_n172 ) );
  INV_X1 u0_u2_u7_U37 (.A( u0_u2_u7_n153 ) , .ZN( u0_u2_u7_n172 ) );
  AOI211_X1 u0_u2_u7_U38 (.B( u0_u2_u7_n139 ) , .A( u0_u2_u7_n140 ) , .C2( u0_u2_u7_n141 ) , .ZN( u0_u2_u7_n142 ) , .C1( u0_u2_u7_n156 ) );
  NAND4_X1 u0_u2_u7_U39 (.A3( u0_u2_u7_n127 ) , .A2( u0_u2_u7_n128 ) , .A1( u0_u2_u7_n129 ) , .ZN( u0_u2_u7_n141 ) , .A4( u0_u2_u7_n147 ) );
  INV_X1 u0_u2_u7_U4 (.A( u0_u2_u7_n111 ) , .ZN( u0_u2_u7_n170 ) );
  AOI21_X1 u0_u2_u7_U40 (.A( u0_u2_u7_n137 ) , .B1( u0_u2_u7_n138 ) , .ZN( u0_u2_u7_n139 ) , .B2( u0_u2_u7_n146 ) );
  OAI22_X1 u0_u2_u7_U41 (.B1( u0_u2_u7_n136 ) , .ZN( u0_u2_u7_n140 ) , .A1( u0_u2_u7_n153 ) , .B2( u0_u2_u7_n162 ) , .A2( u0_u2_u7_n164 ) );
  AOI21_X1 u0_u2_u7_U42 (.ZN( u0_u2_u7_n123 ) , .B1( u0_u2_u7_n165 ) , .B2( u0_u2_u7_n177 ) , .A( u0_u2_u7_n97 ) );
  AOI21_X1 u0_u2_u7_U43 (.B2( u0_u2_u7_n113 ) , .B1( u0_u2_u7_n124 ) , .A( u0_u2_u7_n125 ) , .ZN( u0_u2_u7_n97 ) );
  INV_X1 u0_u2_u7_U44 (.A( u0_u2_u7_n125 ) , .ZN( u0_u2_u7_n161 ) );
  INV_X1 u0_u2_u7_U45 (.A( u0_u2_u7_n152 ) , .ZN( u0_u2_u7_n162 ) );
  AOI22_X1 u0_u2_u7_U46 (.A2( u0_u2_u7_n114 ) , .ZN( u0_u2_u7_n119 ) , .B1( u0_u2_u7_n130 ) , .A1( u0_u2_u7_n156 ) , .B2( u0_u2_u7_n165 ) );
  NAND2_X1 u0_u2_u7_U47 (.A2( u0_u2_u7_n112 ) , .ZN( u0_u2_u7_n114 ) , .A1( u0_u2_u7_n175 ) );
  AND2_X1 u0_u2_u7_U48 (.ZN( u0_u2_u7_n145 ) , .A2( u0_u2_u7_n98 ) , .A1( u0_u2_u7_n99 ) );
  NOR2_X1 u0_u2_u7_U49 (.ZN( u0_u2_u7_n137 ) , .A1( u0_u2_u7_n150 ) , .A2( u0_u2_u7_n161 ) );
  INV_X1 u0_u2_u7_U5 (.A( u0_u2_u7_n149 ) , .ZN( u0_u2_u7_n175 ) );
  AOI21_X1 u0_u2_u7_U50 (.ZN( u0_u2_u7_n105 ) , .B2( u0_u2_u7_n110 ) , .A( u0_u2_u7_n125 ) , .B1( u0_u2_u7_n147 ) );
  NAND2_X1 u0_u2_u7_U51 (.ZN( u0_u2_u7_n146 ) , .A1( u0_u2_u7_n95 ) , .A2( u0_u2_u7_n98 ) );
  NAND2_X1 u0_u2_u7_U52 (.A2( u0_u2_u7_n103 ) , .ZN( u0_u2_u7_n147 ) , .A1( u0_u2_u7_n93 ) );
  NAND2_X1 u0_u2_u7_U53 (.A1( u0_u2_u7_n103 ) , .ZN( u0_u2_u7_n127 ) , .A2( u0_u2_u7_n99 ) );
  OR2_X1 u0_u2_u7_U54 (.ZN( u0_u2_u7_n126 ) , .A2( u0_u2_u7_n152 ) , .A1( u0_u2_u7_n156 ) );
  NAND2_X1 u0_u2_u7_U55 (.A2( u0_u2_u7_n102 ) , .A1( u0_u2_u7_n103 ) , .ZN( u0_u2_u7_n133 ) );
  NAND2_X1 u0_u2_u7_U56 (.ZN( u0_u2_u7_n112 ) , .A2( u0_u2_u7_n96 ) , .A1( u0_u2_u7_n99 ) );
  NAND2_X1 u0_u2_u7_U57 (.A2( u0_u2_u7_n102 ) , .ZN( u0_u2_u7_n128 ) , .A1( u0_u2_u7_n98 ) );
  NAND2_X1 u0_u2_u7_U58 (.A1( u0_u2_u7_n100 ) , .ZN( u0_u2_u7_n113 ) , .A2( u0_u2_u7_n93 ) );
  NAND2_X1 u0_u2_u7_U59 (.A2( u0_u2_u7_n102 ) , .ZN( u0_u2_u7_n124 ) , .A1( u0_u2_u7_n96 ) );
  INV_X1 u0_u2_u7_U6 (.A( u0_u2_u7_n154 ) , .ZN( u0_u2_u7_n178 ) );
  NAND2_X1 u0_u2_u7_U60 (.ZN( u0_u2_u7_n110 ) , .A1( u0_u2_u7_n95 ) , .A2( u0_u2_u7_n96 ) );
  INV_X1 u0_u2_u7_U61 (.A( u0_u2_u7_n150 ) , .ZN( u0_u2_u7_n164 ) );
  AND2_X1 u0_u2_u7_U62 (.ZN( u0_u2_u7_n134 ) , .A1( u0_u2_u7_n93 ) , .A2( u0_u2_u7_n98 ) );
  NAND2_X1 u0_u2_u7_U63 (.A1( u0_u2_u7_n100 ) , .A2( u0_u2_u7_n102 ) , .ZN( u0_u2_u7_n129 ) );
  NAND2_X1 u0_u2_u7_U64 (.A2( u0_u2_u7_n103 ) , .ZN( u0_u2_u7_n131 ) , .A1( u0_u2_u7_n95 ) );
  NAND2_X1 u0_u2_u7_U65 (.A1( u0_u2_u7_n100 ) , .ZN( u0_u2_u7_n138 ) , .A2( u0_u2_u7_n99 ) );
  NAND2_X1 u0_u2_u7_U66 (.ZN( u0_u2_u7_n132 ) , .A1( u0_u2_u7_n93 ) , .A2( u0_u2_u7_n96 ) );
  NAND2_X1 u0_u2_u7_U67 (.A1( u0_u2_u7_n100 ) , .ZN( u0_u2_u7_n148 ) , .A2( u0_u2_u7_n95 ) );
  NOR2_X1 u0_u2_u7_U68 (.A2( u0_u2_X_47 ) , .ZN( u0_u2_u7_n150 ) , .A1( u0_u2_u7_n163 ) );
  NOR2_X1 u0_u2_u7_U69 (.A2( u0_u2_X_43 ) , .A1( u0_u2_X_44 ) , .ZN( u0_u2_u7_n103 ) );
  AOI211_X1 u0_u2_u7_U7 (.ZN( u0_u2_u7_n116 ) , .A( u0_u2_u7_n155 ) , .C1( u0_u2_u7_n161 ) , .C2( u0_u2_u7_n171 ) , .B( u0_u2_u7_n94 ) );
  NOR2_X1 u0_u2_u7_U70 (.A2( u0_u2_X_48 ) , .A1( u0_u2_u7_n166 ) , .ZN( u0_u2_u7_n95 ) );
  NOR2_X1 u0_u2_u7_U71 (.A2( u0_u2_X_45 ) , .A1( u0_u2_X_48 ) , .ZN( u0_u2_u7_n99 ) );
  NOR2_X1 u0_u2_u7_U72 (.A2( u0_u2_X_44 ) , .A1( u0_u2_u7_n167 ) , .ZN( u0_u2_u7_n98 ) );
  NOR2_X1 u0_u2_u7_U73 (.A2( u0_u2_X_46 ) , .A1( u0_u2_X_47 ) , .ZN( u0_u2_u7_n152 ) );
  AND2_X1 u0_u2_u7_U74 (.A1( u0_u2_X_47 ) , .ZN( u0_u2_u7_n156 ) , .A2( u0_u2_u7_n163 ) );
  NAND2_X1 u0_u2_u7_U75 (.A2( u0_u2_X_46 ) , .A1( u0_u2_X_47 ) , .ZN( u0_u2_u7_n125 ) );
  AND2_X1 u0_u2_u7_U76 (.A2( u0_u2_X_45 ) , .A1( u0_u2_X_48 ) , .ZN( u0_u2_u7_n102 ) );
  AND2_X1 u0_u2_u7_U77 (.A2( u0_u2_X_43 ) , .A1( u0_u2_X_44 ) , .ZN( u0_u2_u7_n96 ) );
  AND2_X1 u0_u2_u7_U78 (.A1( u0_u2_X_44 ) , .ZN( u0_u2_u7_n100 ) , .A2( u0_u2_u7_n167 ) );
  AND2_X1 u0_u2_u7_U79 (.A1( u0_u2_X_48 ) , .A2( u0_u2_u7_n166 ) , .ZN( u0_u2_u7_n93 ) );
  OAI222_X1 u0_u2_u7_U8 (.C2( u0_u2_u7_n101 ) , .B2( u0_u2_u7_n111 ) , .A1( u0_u2_u7_n113 ) , .C1( u0_u2_u7_n146 ) , .A2( u0_u2_u7_n162 ) , .B1( u0_u2_u7_n164 ) , .ZN( u0_u2_u7_n94 ) );
  INV_X1 u0_u2_u7_U80 (.A( u0_u2_X_46 ) , .ZN( u0_u2_u7_n163 ) );
  INV_X1 u0_u2_u7_U81 (.A( u0_u2_X_43 ) , .ZN( u0_u2_u7_n167 ) );
  INV_X1 u0_u2_u7_U82 (.A( u0_u2_X_45 ) , .ZN( u0_u2_u7_n166 ) );
  NAND4_X1 u0_u2_u7_U83 (.ZN( u0_out2_5 ) , .A4( u0_u2_u7_n108 ) , .A3( u0_u2_u7_n109 ) , .A1( u0_u2_u7_n116 ) , .A2( u0_u2_u7_n123 ) );
  AOI22_X1 u0_u2_u7_U84 (.ZN( u0_u2_u7_n109 ) , .A2( u0_u2_u7_n126 ) , .B2( u0_u2_u7_n145 ) , .B1( u0_u2_u7_n156 ) , .A1( u0_u2_u7_n171 ) );
  NOR4_X1 u0_u2_u7_U85 (.A4( u0_u2_u7_n104 ) , .A3( u0_u2_u7_n105 ) , .A2( u0_u2_u7_n106 ) , .A1( u0_u2_u7_n107 ) , .ZN( u0_u2_u7_n108 ) );
  NAND4_X1 u0_u2_u7_U86 (.ZN( u0_out2_27 ) , .A4( u0_u2_u7_n118 ) , .A3( u0_u2_u7_n119 ) , .A2( u0_u2_u7_n120 ) , .A1( u0_u2_u7_n121 ) );
  OAI21_X1 u0_u2_u7_U87 (.ZN( u0_u2_u7_n121 ) , .B2( u0_u2_u7_n145 ) , .A( u0_u2_u7_n150 ) , .B1( u0_u2_u7_n174 ) );
  OAI21_X1 u0_u2_u7_U88 (.ZN( u0_u2_u7_n120 ) , .A( u0_u2_u7_n161 ) , .B2( u0_u2_u7_n170 ) , .B1( u0_u2_u7_n179 ) );
  NAND4_X1 u0_u2_u7_U89 (.ZN( u0_out2_21 ) , .A4( u0_u2_u7_n157 ) , .A3( u0_u2_u7_n158 ) , .A2( u0_u2_u7_n159 ) , .A1( u0_u2_u7_n160 ) );
  OAI221_X1 u0_u2_u7_U9 (.C1( u0_u2_u7_n101 ) , .C2( u0_u2_u7_n147 ) , .ZN( u0_u2_u7_n155 ) , .B2( u0_u2_u7_n162 ) , .A( u0_u2_u7_n91 ) , .B1( u0_u2_u7_n92 ) );
  OAI21_X1 u0_u2_u7_U90 (.B1( u0_u2_u7_n145 ) , .ZN( u0_u2_u7_n160 ) , .A( u0_u2_u7_n161 ) , .B2( u0_u2_u7_n177 ) );
  AOI22_X1 u0_u2_u7_U91 (.B2( u0_u2_u7_n149 ) , .B1( u0_u2_u7_n150 ) , .A2( u0_u2_u7_n151 ) , .A1( u0_u2_u7_n152 ) , .ZN( u0_u2_u7_n158 ) );
  NAND4_X1 u0_u2_u7_U92 (.ZN( u0_out2_15 ) , .A4( u0_u2_u7_n142 ) , .A3( u0_u2_u7_n143 ) , .A2( u0_u2_u7_n144 ) , .A1( u0_u2_u7_n178 ) );
  OR2_X1 u0_u2_u7_U93 (.A2( u0_u2_u7_n125 ) , .A1( u0_u2_u7_n129 ) , .ZN( u0_u2_u7_n144 ) );
  AOI22_X1 u0_u2_u7_U94 (.A2( u0_u2_u7_n126 ) , .ZN( u0_u2_u7_n143 ) , .B2( u0_u2_u7_n165 ) , .B1( u0_u2_u7_n173 ) , .A1( u0_u2_u7_n174 ) );
  NAND3_X1 u0_u2_u7_U95 (.A3( u0_u2_u7_n146 ) , .A2( u0_u2_u7_n147 ) , .A1( u0_u2_u7_n148 ) , .ZN( u0_u2_u7_n151 ) );
  NAND3_X1 u0_u2_u7_U96 (.A3( u0_u2_u7_n131 ) , .A2( u0_u2_u7_n132 ) , .A1( u0_u2_u7_n133 ) , .ZN( u0_u2_u7_n135 ) );
  OAI21_X1 u0_uk_U1006 (.ZN( u0_K3_45 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n553 ) , .A( u0_uk_n843 ) );
  NAND2_X1 u0_uk_U1007 (.A1( u0_uk_K_r1_16 ) , .A2( u0_uk_n110 ) , .ZN( u0_uk_n843 ) );
  OAI21_X1 u0_uk_U1050 (.ZN( u0_K15_32 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n33 ) , .A( u0_uk_n918 ) );
  OAI21_X1 u0_uk_U1091 (.ZN( u0_K3_40 ) , .B1( u0_uk_n209 ) , .B2( u0_uk_n558 ) , .A( u0_uk_n845 ) );
  NAND2_X1 u0_uk_U1092 (.A1( u0_uk_K_r1_21 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n845 ) );
  OAI22_X1 u0_uk_U111 (.ZN( u0_K3_41 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n570 ) , .A2( u0_uk_n575 ) );
  OAI22_X1 u0_uk_U230 (.ZN( u0_K15_31 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n28 ) , .B2( u0_uk_n45 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U273 (.ZN( u0_K3_44 ) , .B2( u0_uk_n574 ) , .B1( u0_uk_n83 ) , .A( u0_uk_n844 ) );
  NAND2_X1 u0_uk_U274 (.A1( u0_uk_K_r1_15 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n844 ) );
  OAI22_X1 u0_uk_U275 (.ZN( u0_K3_48 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n546 ) , .B2( u0_uk_n581 ) );
  OAI21_X1 u0_uk_U327 (.ZN( u0_K3_46 ) , .B1( u0_uk_n209 ) , .B2( u0_uk_n561 ) , .A( u0_uk_n842 ) );
  NAND2_X1 u0_uk_U328 (.A1( u0_uk_K_r1_22 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n842 ) );
  BUF_X1 u0_uk_U33 (.Z( u0_uk_n191 ) , .A( u0_uk_n209 ) );
  OAI21_X1 u0_uk_U367 (.ZN( u0_K15_33 ) , .B2( u0_uk_n18 ) , .B1( u0_uk_n83 ) , .A( u0_uk_n917 ) );
  OAI22_X1 u0_uk_U468 (.ZN( u0_K3_37 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n560 ) , .B2( u0_uk_n566 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U544 (.ZN( u0_K15_36 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n18 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n32 ) );
  OAI22_X1 u0_uk_U611 (.ZN( u0_K15_35 ) , .A2( u0_uk_n13 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n28 ) );
  OAI22_X1 u0_uk_U64 (.ZN( u0_K15_34 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n32 ) , .A2( u0_uk_n4 ) );
  OAI22_X1 u0_uk_U652 (.ZN( u0_K3_43 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n550 ) , .B2( u0_uk_n554 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U734 (.ZN( u0_K3_42 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n554 ) , .B2( u0_uk_n581 ) , .B1( u0_uk_n63 ) );
  INV_X1 u0_uk_U8 (.A( u0_uk_n148 ) , .ZN( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U878 (.ZN( u0_K3_47 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n553 ) , .B2( u0_uk_n561 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U926 (.ZN( u0_K3_38 ) , .A1( u0_uk_n191 ) , .B2( u0_uk_n558 ) , .A2( u0_uk_n574 ) , .B1( u0_uk_n63 ) );
  OAI22_X1 u0_uk_U927 (.ZN( u0_K3_39 ) , .A1( u0_uk_n209 ) , .A2( u0_uk_n546 ) , .B2( u0_uk_n550 ) , .B1( u0_uk_n63 ) );
  NAND2_X1 u0_uk_U997 (.A1( u0_uk_K_r5_13 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n777 ) );
  XOR2_X1 u1_U104 (.B( u1_L12_24 ) , .Z( u1_N439 ) , .A( u1_out13_24 ) );
  XOR2_X1 u1_U105 (.B( u1_L12_23 ) , .Z( u1_N438 ) , .A( u1_out13_23 ) );
  XOR2_X1 u1_U110 (.B( u1_L12_18 ) , .Z( u1_N433 ) , .A( u1_out13_18 ) );
  XOR2_X1 u1_U111 (.B( u1_L12_17 ) , .Z( u1_N432 ) , .A( u1_out13_17 ) );
  XOR2_X1 u1_U112 (.B( u1_L12_16 ) , .Z( u1_N431 ) , .A( u1_out13_16 ) );
  XOR2_X1 u1_U116 (.B( u1_L12_13 ) , .Z( u1_N428 ) , .A( u1_out13_13 ) );
  XOR2_X1 u1_U120 (.B( u1_L12_9 ) , .Z( u1_N424 ) , .A( u1_out13_9 ) );
  XOR2_X1 u1_U123 (.B( u1_L12_6 ) , .Z( u1_N421 ) , .A( u1_out13_6 ) );
  XOR2_X1 u1_U128 (.B( u1_L12_2 ) , .Z( u1_N417 ) , .A( u1_out13_2 ) );
  XOR2_X1 u1_U166 (.B( u1_L10_32 ) , .Z( u1_N383 ) , .A( u1_out11_32 ) );
  XOR2_X1 u1_U169 (.B( u1_L10_29 ) , .Z( u1_N380 ) , .A( u1_out11_29 ) );
  XOR2_X1 u1_U172 (.B( u1_L10_27 ) , .Z( u1_N378 ) , .A( u1_out11_27 ) );
  XOR2_X1 u1_U177 (.B( u1_L10_22 ) , .Z( u1_N373 ) , .A( u1_out11_22 ) );
  XOR2_X1 u1_U178 (.B( u1_L10_21 ) , .Z( u1_N372 ) , .A( u1_out11_21 ) );
  XOR2_X1 u1_U180 (.B( u1_L10_19 ) , .Z( u1_N370 ) , .A( u1_out11_19 ) );
  XOR2_X1 u1_U185 (.B( u1_L10_15 ) , .Z( u1_N366 ) , .A( u1_out11_15 ) );
  XOR2_X1 u1_U188 (.B( u1_L10_12 ) , .Z( u1_N363 ) , .A( u1_out11_12 ) );
  XOR2_X1 u1_U189 (.B( u1_L10_11 ) , .Z( u1_N362 ) , .A( u1_out11_11 ) );
  XOR2_X1 u1_U194 (.B( u1_L10_7 ) , .Z( u1_N358 ) , .A( u1_out11_7 ) );
  XOR2_X1 u1_U196 (.B( u1_L10_5 ) , .Z( u1_N356 ) , .A( u1_out11_5 ) );
  XOR2_X1 u1_U197 (.B( u1_L10_4 ) , .Z( u1_N355 ) , .A( u1_out11_4 ) );
  XOR2_X1 u1_U237 (.B( u1_L8_32 ) , .Z( u1_N319 ) , .A( u1_out9_32 ) );
  XOR2_X1 u1_U240 (.B( u1_L8_29 ) , .Z( u1_N316 ) , .A( u1_out9_29 ) );
  XOR2_X1 u1_U248 (.B( u1_L8_22 ) , .Z( u1_N309 ) , .A( u1_out9_22 ) );
  XOR2_X1 u1_U251 (.B( u1_L8_19 ) , .Z( u1_N306 ) , .A( u1_out9_19 ) );
  XOR2_X1 u1_U260 (.B( u1_L8_12 ) , .Z( u1_N299 ) , .A( u1_out9_12 ) );
  XOR2_X1 u1_U261 (.B( u1_L8_11 ) , .Z( u1_N298 ) , .A( u1_out9_11 ) );
  XOR2_X1 u1_U265 (.B( u1_L8_7 ) , .Z( u1_N294 ) , .A( u1_out9_7 ) );
  XOR2_X1 u1_U268 (.B( u1_L8_4 ) , .Z( u1_N291 ) , .A( u1_out9_4 ) );
  XOR2_X1 u1_U313 (.B( u1_L6_27 ) , .Z( u1_N250 ) , .A( u1_out7_27 ) );
  XOR2_X1 u1_U320 (.B( u1_L6_21 ) , .Z( u1_N244 ) , .A( u1_out7_21 ) );
  XOR2_X1 u1_U327 (.B( u1_L6_15 ) , .Z( u1_N238 ) , .A( u1_out7_15 ) );
  XOR2_X1 u1_U338 (.B( u1_L6_5 ) , .Z( u1_N228 ) , .A( u1_out7_5 ) );
  XOR2_X1 u1_U451 (.B( u1_L2_31 ) , .Z( u1_N126 ) , .A( u1_out3_31 ) );
  XOR2_X1 u1_U452 (.B( u1_L2_30 ) , .Z( u1_N125 ) , .A( u1_out3_30 ) );
  XOR2_X1 u1_U455 (.B( u1_L2_27 ) , .Z( u1_N122 ) , .A( u1_out3_27 ) );
  XOR2_X1 u1_U456 (.B( u1_L2_26 ) , .Z( u1_N121 ) , .A( u1_out3_26 ) );
  XOR2_X1 u1_U459 (.B( u1_L2_24 ) , .Z( u1_N119 ) , .A( u1_out3_24 ) );
  XOR2_X1 u1_U460 (.B( u1_L2_23 ) , .Z( u1_N118 ) , .A( u1_out3_23 ) );
  XOR2_X1 u1_U462 (.B( u1_L2_21 ) , .Z( u1_N116 ) , .A( u1_out3_21 ) );
  XOR2_X1 u1_U463 (.B( u1_L2_20 ) , .Z( u1_N115 ) , .A( u1_out3_20 ) );
  XOR2_X1 u1_U466 (.B( u1_L2_17 ) , .Z( u1_N112 ) , .A( u1_out3_17 ) );
  XOR2_X1 u1_U467 (.B( u1_L2_16 ) , .Z( u1_N111 ) , .A( u1_out3_16 ) );
  XOR2_X1 u1_U468 (.B( u1_L2_15 ) , .Z( u1_N110 ) , .A( u1_out3_15 ) );
  XOR2_X1 u1_U474 (.B( u1_L2_10 ) , .Z( u1_N105 ) , .A( u1_out3_10 ) );
  XOR2_X1 u1_U475 (.B( u1_L2_9 ) , .Z( u1_N104 ) , .A( u1_out3_9 ) );
  XOR2_X1 u1_U478 (.B( u1_L2_6 ) , .Z( u1_N101 ) , .A( u1_out3_6 ) );
  XOR2_X1 u1_U479 (.B( u1_L2_5 ) , .Z( u1_N100 ) , .A( u1_out3_5 ) );
  XOR2_X1 u1_U483 (.Z( u1_FP_9 ) , .B( u1_L14_9 ) , .A( u1_out15_9 ) );
  XOR2_X1 u1_U491 (.Z( u1_FP_31 ) , .B( u1_L14_31 ) , .A( u1_out15_31 ) );
  XOR2_X1 u1_U493 (.Z( u1_FP_2 ) , .B( u1_L14_2 ) , .A( u1_out15_2 ) );
  XOR2_X1 u1_U495 (.Z( u1_FP_28 ) , .B( u1_L14_28 ) , .A( u1_out15_28 ) );
  XOR2_X1 u1_U497 (.Z( u1_FP_26 ) , .B( u1_L14_26 ) , .A( u1_out15_26 ) );
  XOR2_X1 u1_U500 (.Z( u1_FP_23 ) , .B( u1_L14_23 ) , .A( u1_out15_23 ) );
  XOR2_X1 u1_U503 (.Z( u1_FP_20 ) , .B( u1_L14_20 ) , .A( u1_out15_20 ) );
  XOR2_X1 u1_U504 (.Z( u1_FP_1 ) , .B( u1_L14_1 ) , .A( u1_out15_1 ) );
  XOR2_X1 u1_U506 (.Z( u1_FP_18 ) , .B( u1_L14_18 ) , .A( u1_out15_18 ) );
  XOR2_X1 u1_U507 (.Z( u1_FP_17 ) , .B( u1_L14_17 ) , .A( u1_out15_17 ) );
  XOR2_X1 u1_U511 (.Z( u1_FP_13 ) , .B( u1_L14_13 ) , .A( u1_out15_13 ) );
  XOR2_X1 u1_U514 (.Z( u1_FP_10 ) , .B( u1_L14_10 ) , .A( u1_out15_10 ) );
  XOR2_X1 u1_U6 (.B( u1_L2_1 ) , .Z( u1_N96 ) , .A( u1_out3_1 ) );
  XOR2_X1 u1_U96 (.B( u1_L12_31 ) , .Z( u1_N446 ) , .A( u1_out13_31 ) );
  XOR2_X1 u1_U97 (.B( u1_L12_30 ) , .Z( u1_N445 ) , .A( u1_out13_30 ) );
  XOR2_X1 u1_U99 (.B( u1_L12_28 ) , .Z( u1_N443 ) , .A( u1_out13_28 ) );
  XOR2_X1 u1_u11_U10 (.B( u1_K12_45 ) , .A( u1_R10_30 ) , .Z( u1_u11_X_45 ) );
  XOR2_X1 u1_u11_U11 (.B( u1_K12_44 ) , .A( u1_R10_29 ) , .Z( u1_u11_X_44 ) );
  XOR2_X1 u1_u11_U12 (.B( u1_K12_43 ) , .A( u1_R10_28 ) , .Z( u1_u11_X_43 ) );
  XOR2_X1 u1_u11_U13 (.B( u1_K12_42 ) , .A( u1_R10_29 ) , .Z( u1_u11_X_42 ) );
  XOR2_X1 u1_u11_U14 (.B( u1_K12_41 ) , .A( u1_R10_28 ) , .Z( u1_u11_X_41 ) );
  XOR2_X1 u1_u11_U15 (.B( u1_K12_40 ) , .A( u1_R10_27 ) , .Z( u1_u11_X_40 ) );
  XOR2_X1 u1_u11_U17 (.B( u1_K12_39 ) , .A( u1_R10_26 ) , .Z( u1_u11_X_39 ) );
  XOR2_X1 u1_u11_U18 (.B( u1_K12_38 ) , .A( u1_R10_25 ) , .Z( u1_u11_X_38 ) );
  XOR2_X1 u1_u11_U19 (.B( u1_K12_37 ) , .A( u1_R10_24 ) , .Z( u1_u11_X_37 ) );
  XOR2_X1 u1_u11_U20 (.B( u1_K12_36 ) , .A( u1_R10_25 ) , .Z( u1_u11_X_36 ) );
  XOR2_X1 u1_u11_U21 (.B( u1_K12_35 ) , .A( u1_R10_24 ) , .Z( u1_u11_X_35 ) );
  XOR2_X1 u1_u11_U22 (.B( u1_K12_34 ) , .A( u1_R10_23 ) , .Z( u1_u11_X_34 ) );
  XOR2_X1 u1_u11_U23 (.B( u1_K12_33 ) , .A( u1_R10_22 ) , .Z( u1_u11_X_33 ) );
  XOR2_X1 u1_u11_U24 (.B( u1_K12_32 ) , .A( u1_R10_21 ) , .Z( u1_u11_X_32 ) );
  XOR2_X1 u1_u11_U25 (.B( u1_K12_31 ) , .A( u1_R10_20 ) , .Z( u1_u11_X_31 ) );
  XOR2_X1 u1_u11_U7 (.B( u1_K12_48 ) , .A( u1_R10_1 ) , .Z( u1_u11_X_48 ) );
  XOR2_X1 u1_u11_U8 (.B( u1_K12_47 ) , .A( u1_R10_32 ) , .Z( u1_u11_X_47 ) );
  XOR2_X1 u1_u11_U9 (.B( u1_K12_46 ) , .A( u1_R10_31 ) , .Z( u1_u11_X_46 ) );
  INV_X1 u1_u11_u5_U10 (.A( u1_u11_u5_n121 ) , .ZN( u1_u11_u5_n177 ) );
  NOR3_X1 u1_u11_u5_U100 (.A3( u1_u11_u5_n141 ) , .A1( u1_u11_u5_n142 ) , .ZN( u1_u11_u5_n143 ) , .A2( u1_u11_u5_n191 ) );
  NAND4_X1 u1_u11_u5_U101 (.ZN( u1_out11_4 ) , .A4( u1_u11_u5_n112 ) , .A2( u1_u11_u5_n113 ) , .A1( u1_u11_u5_n114 ) , .A3( u1_u11_u5_n195 ) );
  AOI211_X1 u1_u11_u5_U102 (.A( u1_u11_u5_n110 ) , .C1( u1_u11_u5_n111 ) , .ZN( u1_u11_u5_n112 ) , .B( u1_u11_u5_n118 ) , .C2( u1_u11_u5_n177 ) );
  AOI222_X1 u1_u11_u5_U103 (.ZN( u1_u11_u5_n113 ) , .A1( u1_u11_u5_n131 ) , .C1( u1_u11_u5_n148 ) , .B2( u1_u11_u5_n174 ) , .C2( u1_u11_u5_n178 ) , .A2( u1_u11_u5_n179 ) , .B1( u1_u11_u5_n99 ) );
  NAND3_X1 u1_u11_u5_U104 (.A2( u1_u11_u5_n154 ) , .A3( u1_u11_u5_n158 ) , .A1( u1_u11_u5_n161 ) , .ZN( u1_u11_u5_n99 ) );
  NOR2_X1 u1_u11_u5_U11 (.ZN( u1_u11_u5_n160 ) , .A2( u1_u11_u5_n173 ) , .A1( u1_u11_u5_n177 ) );
  INV_X1 u1_u11_u5_U12 (.A( u1_u11_u5_n150 ) , .ZN( u1_u11_u5_n174 ) );
  AOI21_X1 u1_u11_u5_U13 (.A( u1_u11_u5_n160 ) , .B2( u1_u11_u5_n161 ) , .ZN( u1_u11_u5_n162 ) , .B1( u1_u11_u5_n192 ) );
  INV_X1 u1_u11_u5_U14 (.A( u1_u11_u5_n159 ) , .ZN( u1_u11_u5_n192 ) );
  AOI21_X1 u1_u11_u5_U15 (.A( u1_u11_u5_n156 ) , .B2( u1_u11_u5_n157 ) , .B1( u1_u11_u5_n158 ) , .ZN( u1_u11_u5_n163 ) );
  AOI21_X1 u1_u11_u5_U16 (.B2( u1_u11_u5_n139 ) , .B1( u1_u11_u5_n140 ) , .ZN( u1_u11_u5_n141 ) , .A( u1_u11_u5_n150 ) );
  OAI21_X1 u1_u11_u5_U17 (.A( u1_u11_u5_n133 ) , .B2( u1_u11_u5_n134 ) , .B1( u1_u11_u5_n135 ) , .ZN( u1_u11_u5_n142 ) );
  OAI21_X1 u1_u11_u5_U18 (.ZN( u1_u11_u5_n133 ) , .B2( u1_u11_u5_n147 ) , .A( u1_u11_u5_n173 ) , .B1( u1_u11_u5_n188 ) );
  NAND2_X1 u1_u11_u5_U19 (.A2( u1_u11_u5_n119 ) , .A1( u1_u11_u5_n123 ) , .ZN( u1_u11_u5_n137 ) );
  INV_X1 u1_u11_u5_U20 (.A( u1_u11_u5_n155 ) , .ZN( u1_u11_u5_n194 ) );
  NAND2_X1 u1_u11_u5_U21 (.A1( u1_u11_u5_n121 ) , .ZN( u1_u11_u5_n132 ) , .A2( u1_u11_u5_n172 ) );
  NAND2_X1 u1_u11_u5_U22 (.A2( u1_u11_u5_n122 ) , .ZN( u1_u11_u5_n136 ) , .A1( u1_u11_u5_n154 ) );
  NAND2_X1 u1_u11_u5_U23 (.A2( u1_u11_u5_n119 ) , .A1( u1_u11_u5_n120 ) , .ZN( u1_u11_u5_n159 ) );
  INV_X1 u1_u11_u5_U24 (.A( u1_u11_u5_n156 ) , .ZN( u1_u11_u5_n175 ) );
  INV_X1 u1_u11_u5_U25 (.A( u1_u11_u5_n158 ) , .ZN( u1_u11_u5_n188 ) );
  INV_X1 u1_u11_u5_U26 (.A( u1_u11_u5_n152 ) , .ZN( u1_u11_u5_n179 ) );
  INV_X1 u1_u11_u5_U27 (.A( u1_u11_u5_n140 ) , .ZN( u1_u11_u5_n182 ) );
  INV_X1 u1_u11_u5_U28 (.A( u1_u11_u5_n151 ) , .ZN( u1_u11_u5_n183 ) );
  INV_X1 u1_u11_u5_U29 (.A( u1_u11_u5_n123 ) , .ZN( u1_u11_u5_n185 ) );
  NOR2_X1 u1_u11_u5_U3 (.ZN( u1_u11_u5_n134 ) , .A1( u1_u11_u5_n183 ) , .A2( u1_u11_u5_n190 ) );
  INV_X1 u1_u11_u5_U30 (.A( u1_u11_u5_n161 ) , .ZN( u1_u11_u5_n184 ) );
  INV_X1 u1_u11_u5_U31 (.A( u1_u11_u5_n139 ) , .ZN( u1_u11_u5_n189 ) );
  INV_X1 u1_u11_u5_U32 (.A( u1_u11_u5_n157 ) , .ZN( u1_u11_u5_n190 ) );
  INV_X1 u1_u11_u5_U33 (.A( u1_u11_u5_n120 ) , .ZN( u1_u11_u5_n193 ) );
  NAND2_X1 u1_u11_u5_U34 (.ZN( u1_u11_u5_n111 ) , .A1( u1_u11_u5_n140 ) , .A2( u1_u11_u5_n155 ) );
  NOR2_X1 u1_u11_u5_U35 (.ZN( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n170 ) , .A2( u1_u11_u5_n180 ) );
  INV_X1 u1_u11_u5_U36 (.A( u1_u11_u5_n117 ) , .ZN( u1_u11_u5_n196 ) );
  OAI221_X1 u1_u11_u5_U37 (.A( u1_u11_u5_n116 ) , .ZN( u1_u11_u5_n117 ) , .B2( u1_u11_u5_n119 ) , .C1( u1_u11_u5_n153 ) , .C2( u1_u11_u5_n158 ) , .B1( u1_u11_u5_n172 ) );
  AOI222_X1 u1_u11_u5_U38 (.ZN( u1_u11_u5_n116 ) , .B2( u1_u11_u5_n145 ) , .C1( u1_u11_u5_n148 ) , .A2( u1_u11_u5_n174 ) , .C2( u1_u11_u5_n177 ) , .B1( u1_u11_u5_n187 ) , .A1( u1_u11_u5_n193 ) );
  INV_X1 u1_u11_u5_U39 (.A( u1_u11_u5_n115 ) , .ZN( u1_u11_u5_n187 ) );
  INV_X1 u1_u11_u5_U4 (.A( u1_u11_u5_n138 ) , .ZN( u1_u11_u5_n191 ) );
  AOI22_X1 u1_u11_u5_U40 (.B2( u1_u11_u5_n131 ) , .A2( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n169 ) , .B1( u1_u11_u5_n174 ) , .A1( u1_u11_u5_n185 ) );
  NOR2_X1 u1_u11_u5_U41 (.A1( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n150 ) , .A2( u1_u11_u5_n173 ) );
  AOI21_X1 u1_u11_u5_U42 (.A( u1_u11_u5_n118 ) , .B2( u1_u11_u5_n145 ) , .ZN( u1_u11_u5_n168 ) , .B1( u1_u11_u5_n186 ) );
  INV_X1 u1_u11_u5_U43 (.A( u1_u11_u5_n122 ) , .ZN( u1_u11_u5_n186 ) );
  NOR2_X1 u1_u11_u5_U44 (.A1( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n152 ) , .A2( u1_u11_u5_n176 ) );
  NOR2_X1 u1_u11_u5_U45 (.A1( u1_u11_u5_n115 ) , .ZN( u1_u11_u5_n118 ) , .A2( u1_u11_u5_n153 ) );
  NOR2_X1 u1_u11_u5_U46 (.A2( u1_u11_u5_n145 ) , .ZN( u1_u11_u5_n156 ) , .A1( u1_u11_u5_n174 ) );
  NOR2_X1 u1_u11_u5_U47 (.ZN( u1_u11_u5_n121 ) , .A2( u1_u11_u5_n145 ) , .A1( u1_u11_u5_n176 ) );
  AOI22_X1 u1_u11_u5_U48 (.ZN( u1_u11_u5_n114 ) , .A2( u1_u11_u5_n137 ) , .A1( u1_u11_u5_n145 ) , .B2( u1_u11_u5_n175 ) , .B1( u1_u11_u5_n193 ) );
  OAI211_X1 u1_u11_u5_U49 (.B( u1_u11_u5_n124 ) , .A( u1_u11_u5_n125 ) , .C2( u1_u11_u5_n126 ) , .C1( u1_u11_u5_n127 ) , .ZN( u1_u11_u5_n128 ) );
  OAI21_X1 u1_u11_u5_U5 (.B2( u1_u11_u5_n136 ) , .B1( u1_u11_u5_n137 ) , .ZN( u1_u11_u5_n138 ) , .A( u1_u11_u5_n177 ) );
  OAI21_X1 u1_u11_u5_U50 (.ZN( u1_u11_u5_n124 ) , .A( u1_u11_u5_n177 ) , .B2( u1_u11_u5_n183 ) , .B1( u1_u11_u5_n189 ) );
  NOR3_X1 u1_u11_u5_U51 (.ZN( u1_u11_u5_n127 ) , .A1( u1_u11_u5_n136 ) , .A3( u1_u11_u5_n148 ) , .A2( u1_u11_u5_n182 ) );
  OAI21_X1 u1_u11_u5_U52 (.ZN( u1_u11_u5_n125 ) , .A( u1_u11_u5_n174 ) , .B2( u1_u11_u5_n185 ) , .B1( u1_u11_u5_n190 ) );
  AOI21_X1 u1_u11_u5_U53 (.A( u1_u11_u5_n153 ) , .B2( u1_u11_u5_n154 ) , .B1( u1_u11_u5_n155 ) , .ZN( u1_u11_u5_n164 ) );
  AOI21_X1 u1_u11_u5_U54 (.ZN( u1_u11_u5_n110 ) , .B1( u1_u11_u5_n122 ) , .B2( u1_u11_u5_n139 ) , .A( u1_u11_u5_n153 ) );
  INV_X1 u1_u11_u5_U55 (.A( u1_u11_u5_n153 ) , .ZN( u1_u11_u5_n176 ) );
  INV_X1 u1_u11_u5_U56 (.A( u1_u11_u5_n126 ) , .ZN( u1_u11_u5_n173 ) );
  AND2_X1 u1_u11_u5_U57 (.A2( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n107 ) , .ZN( u1_u11_u5_n147 ) );
  AND2_X1 u1_u11_u5_U58 (.A2( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n108 ) , .ZN( u1_u11_u5_n148 ) );
  NAND2_X1 u1_u11_u5_U59 (.A1( u1_u11_u5_n105 ) , .A2( u1_u11_u5_n106 ) , .ZN( u1_u11_u5_n158 ) );
  INV_X1 u1_u11_u5_U6 (.A( u1_u11_u5_n135 ) , .ZN( u1_u11_u5_n178 ) );
  NAND2_X1 u1_u11_u5_U60 (.A2( u1_u11_u5_n108 ) , .A1( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n139 ) );
  NAND2_X1 u1_u11_u5_U61 (.A1( u1_u11_u5_n106 ) , .A2( u1_u11_u5_n108 ) , .ZN( u1_u11_u5_n119 ) );
  NAND2_X1 u1_u11_u5_U62 (.A2( u1_u11_u5_n103 ) , .A1( u1_u11_u5_n105 ) , .ZN( u1_u11_u5_n140 ) );
  NAND2_X1 u1_u11_u5_U63 (.A2( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n105 ) , .ZN( u1_u11_u5_n155 ) );
  NAND2_X1 u1_u11_u5_U64 (.A2( u1_u11_u5_n106 ) , .A1( u1_u11_u5_n107 ) , .ZN( u1_u11_u5_n122 ) );
  NAND2_X1 u1_u11_u5_U65 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n106 ) , .ZN( u1_u11_u5_n115 ) );
  NAND2_X1 u1_u11_u5_U66 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n103 ) , .ZN( u1_u11_u5_n161 ) );
  NAND2_X1 u1_u11_u5_U67 (.A1( u1_u11_u5_n105 ) , .A2( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n154 ) );
  INV_X1 u1_u11_u5_U68 (.A( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n172 ) );
  NAND2_X1 u1_u11_u5_U69 (.A1( u1_u11_u5_n103 ) , .A2( u1_u11_u5_n108 ) , .ZN( u1_u11_u5_n123 ) );
  OAI22_X1 u1_u11_u5_U7 (.B2( u1_u11_u5_n149 ) , .B1( u1_u11_u5_n150 ) , .A2( u1_u11_u5_n151 ) , .A1( u1_u11_u5_n152 ) , .ZN( u1_u11_u5_n165 ) );
  NAND2_X1 u1_u11_u5_U70 (.A2( u1_u11_u5_n103 ) , .A1( u1_u11_u5_n107 ) , .ZN( u1_u11_u5_n151 ) );
  NAND2_X1 u1_u11_u5_U71 (.A2( u1_u11_u5_n107 ) , .A1( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n120 ) );
  NAND2_X1 u1_u11_u5_U72 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n157 ) );
  AND2_X1 u1_u11_u5_U73 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n104 ) , .ZN( u1_u11_u5_n131 ) );
  INV_X1 u1_u11_u5_U74 (.A( u1_u11_u5_n102 ) , .ZN( u1_u11_u5_n195 ) );
  OAI221_X1 u1_u11_u5_U75 (.A( u1_u11_u5_n101 ) , .ZN( u1_u11_u5_n102 ) , .C2( u1_u11_u5_n115 ) , .C1( u1_u11_u5_n126 ) , .B1( u1_u11_u5_n134 ) , .B2( u1_u11_u5_n160 ) );
  OAI21_X1 u1_u11_u5_U76 (.ZN( u1_u11_u5_n101 ) , .B1( u1_u11_u5_n137 ) , .A( u1_u11_u5_n146 ) , .B2( u1_u11_u5_n147 ) );
  NOR2_X1 u1_u11_u5_U77 (.A2( u1_u11_X_34 ) , .A1( u1_u11_X_35 ) , .ZN( u1_u11_u5_n145 ) );
  NOR2_X1 u1_u11_u5_U78 (.A2( u1_u11_X_34 ) , .ZN( u1_u11_u5_n146 ) , .A1( u1_u11_u5_n171 ) );
  NOR2_X1 u1_u11_u5_U79 (.A2( u1_u11_X_31 ) , .A1( u1_u11_X_32 ) , .ZN( u1_u11_u5_n103 ) );
  NOR3_X1 u1_u11_u5_U8 (.A2( u1_u11_u5_n147 ) , .A1( u1_u11_u5_n148 ) , .ZN( u1_u11_u5_n149 ) , .A3( u1_u11_u5_n194 ) );
  NOR2_X1 u1_u11_u5_U80 (.A2( u1_u11_X_36 ) , .ZN( u1_u11_u5_n105 ) , .A1( u1_u11_u5_n180 ) );
  NOR2_X1 u1_u11_u5_U81 (.A2( u1_u11_X_33 ) , .ZN( u1_u11_u5_n108 ) , .A1( u1_u11_u5_n170 ) );
  NOR2_X1 u1_u11_u5_U82 (.A2( u1_u11_X_33 ) , .A1( u1_u11_X_36 ) , .ZN( u1_u11_u5_n107 ) );
  NOR2_X1 u1_u11_u5_U83 (.A2( u1_u11_X_31 ) , .ZN( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n181 ) );
  NAND2_X1 u1_u11_u5_U84 (.A2( u1_u11_X_34 ) , .A1( u1_u11_X_35 ) , .ZN( u1_u11_u5_n153 ) );
  NAND2_X1 u1_u11_u5_U85 (.A1( u1_u11_X_34 ) , .ZN( u1_u11_u5_n126 ) , .A2( u1_u11_u5_n171 ) );
  AND2_X1 u1_u11_u5_U86 (.A1( u1_u11_X_31 ) , .A2( u1_u11_X_32 ) , .ZN( u1_u11_u5_n106 ) );
  AND2_X1 u1_u11_u5_U87 (.A1( u1_u11_X_31 ) , .ZN( u1_u11_u5_n109 ) , .A2( u1_u11_u5_n181 ) );
  INV_X1 u1_u11_u5_U88 (.A( u1_u11_X_33 ) , .ZN( u1_u11_u5_n180 ) );
  INV_X1 u1_u11_u5_U89 (.A( u1_u11_X_35 ) , .ZN( u1_u11_u5_n171 ) );
  NOR2_X1 u1_u11_u5_U9 (.ZN( u1_u11_u5_n135 ) , .A1( u1_u11_u5_n173 ) , .A2( u1_u11_u5_n176 ) );
  INV_X1 u1_u11_u5_U90 (.A( u1_u11_X_36 ) , .ZN( u1_u11_u5_n170 ) );
  INV_X1 u1_u11_u5_U91 (.A( u1_u11_X_32 ) , .ZN( u1_u11_u5_n181 ) );
  NAND4_X1 u1_u11_u5_U92 (.ZN( u1_out11_29 ) , .A4( u1_u11_u5_n129 ) , .A3( u1_u11_u5_n130 ) , .A2( u1_u11_u5_n168 ) , .A1( u1_u11_u5_n196 ) );
  AOI221_X1 u1_u11_u5_U93 (.A( u1_u11_u5_n128 ) , .ZN( u1_u11_u5_n129 ) , .C2( u1_u11_u5_n132 ) , .B2( u1_u11_u5_n159 ) , .B1( u1_u11_u5_n176 ) , .C1( u1_u11_u5_n184 ) );
  AOI222_X1 u1_u11_u5_U94 (.ZN( u1_u11_u5_n130 ) , .A2( u1_u11_u5_n146 ) , .B1( u1_u11_u5_n147 ) , .C2( u1_u11_u5_n175 ) , .B2( u1_u11_u5_n179 ) , .A1( u1_u11_u5_n188 ) , .C1( u1_u11_u5_n194 ) );
  NAND4_X1 u1_u11_u5_U95 (.ZN( u1_out11_19 ) , .A4( u1_u11_u5_n166 ) , .A3( u1_u11_u5_n167 ) , .A2( u1_u11_u5_n168 ) , .A1( u1_u11_u5_n169 ) );
  AOI22_X1 u1_u11_u5_U96 (.B2( u1_u11_u5_n145 ) , .A2( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n167 ) , .B1( u1_u11_u5_n182 ) , .A1( u1_u11_u5_n189 ) );
  NOR4_X1 u1_u11_u5_U97 (.A4( u1_u11_u5_n162 ) , .A3( u1_u11_u5_n163 ) , .A2( u1_u11_u5_n164 ) , .A1( u1_u11_u5_n165 ) , .ZN( u1_u11_u5_n166 ) );
  NAND4_X1 u1_u11_u5_U98 (.ZN( u1_out11_11 ) , .A4( u1_u11_u5_n143 ) , .A3( u1_u11_u5_n144 ) , .A2( u1_u11_u5_n169 ) , .A1( u1_u11_u5_n196 ) );
  AOI22_X1 u1_u11_u5_U99 (.A2( u1_u11_u5_n132 ) , .ZN( u1_u11_u5_n144 ) , .B2( u1_u11_u5_n145 ) , .B1( u1_u11_u5_n184 ) , .A1( u1_u11_u5_n194 ) );
  OAI21_X1 u1_u11_u6_U10 (.A( u1_u11_u6_n159 ) , .B1( u1_u11_u6_n169 ) , .B2( u1_u11_u6_n173 ) , .ZN( u1_u11_u6_n90 ) );
  INV_X1 u1_u11_u6_U11 (.ZN( u1_u11_u6_n172 ) , .A( u1_u11_u6_n88 ) );
  AOI22_X1 u1_u11_u6_U12 (.A2( u1_u11_u6_n151 ) , .B2( u1_u11_u6_n161 ) , .A1( u1_u11_u6_n167 ) , .B1( u1_u11_u6_n170 ) , .ZN( u1_u11_u6_n89 ) );
  AOI21_X1 u1_u11_u6_U13 (.ZN( u1_u11_u6_n106 ) , .A( u1_u11_u6_n142 ) , .B2( u1_u11_u6_n159 ) , .B1( u1_u11_u6_n164 ) );
  INV_X1 u1_u11_u6_U14 (.A( u1_u11_u6_n155 ) , .ZN( u1_u11_u6_n161 ) );
  INV_X1 u1_u11_u6_U15 (.A( u1_u11_u6_n128 ) , .ZN( u1_u11_u6_n164 ) );
  NAND2_X1 u1_u11_u6_U16 (.ZN( u1_u11_u6_n110 ) , .A1( u1_u11_u6_n122 ) , .A2( u1_u11_u6_n129 ) );
  NAND2_X1 u1_u11_u6_U17 (.ZN( u1_u11_u6_n124 ) , .A2( u1_u11_u6_n146 ) , .A1( u1_u11_u6_n148 ) );
  INV_X1 u1_u11_u6_U18 (.A( u1_u11_u6_n132 ) , .ZN( u1_u11_u6_n171 ) );
  AND2_X1 u1_u11_u6_U19 (.A1( u1_u11_u6_n100 ) , .ZN( u1_u11_u6_n130 ) , .A2( u1_u11_u6_n147 ) );
  INV_X1 u1_u11_u6_U20 (.A( u1_u11_u6_n127 ) , .ZN( u1_u11_u6_n173 ) );
  INV_X1 u1_u11_u6_U21 (.A( u1_u11_u6_n121 ) , .ZN( u1_u11_u6_n167 ) );
  INV_X1 u1_u11_u6_U22 (.A( u1_u11_u6_n100 ) , .ZN( u1_u11_u6_n169 ) );
  INV_X1 u1_u11_u6_U23 (.A( u1_u11_u6_n123 ) , .ZN( u1_u11_u6_n170 ) );
  INV_X1 u1_u11_u6_U24 (.A( u1_u11_u6_n113 ) , .ZN( u1_u11_u6_n168 ) );
  AND2_X1 u1_u11_u6_U25 (.A1( u1_u11_u6_n107 ) , .A2( u1_u11_u6_n119 ) , .ZN( u1_u11_u6_n133 ) );
  AND2_X1 u1_u11_u6_U26 (.A2( u1_u11_u6_n121 ) , .A1( u1_u11_u6_n122 ) , .ZN( u1_u11_u6_n131 ) );
  AND3_X1 u1_u11_u6_U27 (.ZN( u1_u11_u6_n120 ) , .A2( u1_u11_u6_n127 ) , .A1( u1_u11_u6_n132 ) , .A3( u1_u11_u6_n145 ) );
  INV_X1 u1_u11_u6_U28 (.A( u1_u11_u6_n146 ) , .ZN( u1_u11_u6_n163 ) );
  AOI222_X1 u1_u11_u6_U29 (.ZN( u1_u11_u6_n114 ) , .A1( u1_u11_u6_n118 ) , .A2( u1_u11_u6_n126 ) , .B2( u1_u11_u6_n151 ) , .C2( u1_u11_u6_n159 ) , .C1( u1_u11_u6_n168 ) , .B1( u1_u11_u6_n169 ) );
  INV_X1 u1_u11_u6_U3 (.A( u1_u11_u6_n110 ) , .ZN( u1_u11_u6_n166 ) );
  NOR2_X1 u1_u11_u6_U30 (.A1( u1_u11_u6_n162 ) , .A2( u1_u11_u6_n165 ) , .ZN( u1_u11_u6_n98 ) );
  NAND2_X1 u1_u11_u6_U31 (.A1( u1_u11_u6_n144 ) , .ZN( u1_u11_u6_n151 ) , .A2( u1_u11_u6_n158 ) );
  NAND2_X1 u1_u11_u6_U32 (.ZN( u1_u11_u6_n132 ) , .A1( u1_u11_u6_n91 ) , .A2( u1_u11_u6_n97 ) );
  AOI22_X1 u1_u11_u6_U33 (.B2( u1_u11_u6_n110 ) , .B1( u1_u11_u6_n111 ) , .A1( u1_u11_u6_n112 ) , .ZN( u1_u11_u6_n115 ) , .A2( u1_u11_u6_n161 ) );
  NAND4_X1 u1_u11_u6_U34 (.A3( u1_u11_u6_n109 ) , .ZN( u1_u11_u6_n112 ) , .A4( u1_u11_u6_n132 ) , .A2( u1_u11_u6_n147 ) , .A1( u1_u11_u6_n166 ) );
  NOR2_X1 u1_u11_u6_U35 (.ZN( u1_u11_u6_n109 ) , .A1( u1_u11_u6_n170 ) , .A2( u1_u11_u6_n173 ) );
  NOR2_X1 u1_u11_u6_U36 (.A2( u1_u11_u6_n126 ) , .ZN( u1_u11_u6_n155 ) , .A1( u1_u11_u6_n160 ) );
  NAND2_X1 u1_u11_u6_U37 (.ZN( u1_u11_u6_n146 ) , .A2( u1_u11_u6_n94 ) , .A1( u1_u11_u6_n99 ) );
  AOI21_X1 u1_u11_u6_U38 (.A( u1_u11_u6_n144 ) , .B2( u1_u11_u6_n145 ) , .B1( u1_u11_u6_n146 ) , .ZN( u1_u11_u6_n150 ) );
  AOI211_X1 u1_u11_u6_U39 (.B( u1_u11_u6_n134 ) , .A( u1_u11_u6_n135 ) , .C1( u1_u11_u6_n136 ) , .ZN( u1_u11_u6_n137 ) , .C2( u1_u11_u6_n151 ) );
  INV_X1 u1_u11_u6_U4 (.A( u1_u11_u6_n142 ) , .ZN( u1_u11_u6_n174 ) );
  NAND4_X1 u1_u11_u6_U40 (.A4( u1_u11_u6_n127 ) , .A3( u1_u11_u6_n128 ) , .A2( u1_u11_u6_n129 ) , .A1( u1_u11_u6_n130 ) , .ZN( u1_u11_u6_n136 ) );
  AOI21_X1 u1_u11_u6_U41 (.B2( u1_u11_u6_n132 ) , .B1( u1_u11_u6_n133 ) , .ZN( u1_u11_u6_n134 ) , .A( u1_u11_u6_n158 ) );
  AOI21_X1 u1_u11_u6_U42 (.B1( u1_u11_u6_n131 ) , .ZN( u1_u11_u6_n135 ) , .A( u1_u11_u6_n144 ) , .B2( u1_u11_u6_n146 ) );
  INV_X1 u1_u11_u6_U43 (.A( u1_u11_u6_n111 ) , .ZN( u1_u11_u6_n158 ) );
  NAND2_X1 u1_u11_u6_U44 (.ZN( u1_u11_u6_n127 ) , .A1( u1_u11_u6_n91 ) , .A2( u1_u11_u6_n92 ) );
  NAND2_X1 u1_u11_u6_U45 (.ZN( u1_u11_u6_n129 ) , .A2( u1_u11_u6_n95 ) , .A1( u1_u11_u6_n96 ) );
  INV_X1 u1_u11_u6_U46 (.A( u1_u11_u6_n144 ) , .ZN( u1_u11_u6_n159 ) );
  NAND2_X1 u1_u11_u6_U47 (.ZN( u1_u11_u6_n145 ) , .A2( u1_u11_u6_n97 ) , .A1( u1_u11_u6_n98 ) );
  NAND2_X1 u1_u11_u6_U48 (.ZN( u1_u11_u6_n148 ) , .A2( u1_u11_u6_n92 ) , .A1( u1_u11_u6_n94 ) );
  NAND2_X1 u1_u11_u6_U49 (.ZN( u1_u11_u6_n108 ) , .A2( u1_u11_u6_n139 ) , .A1( u1_u11_u6_n144 ) );
  NAND2_X1 u1_u11_u6_U5 (.A2( u1_u11_u6_n143 ) , .ZN( u1_u11_u6_n152 ) , .A1( u1_u11_u6_n166 ) );
  NAND2_X1 u1_u11_u6_U50 (.ZN( u1_u11_u6_n121 ) , .A2( u1_u11_u6_n95 ) , .A1( u1_u11_u6_n97 ) );
  NAND2_X1 u1_u11_u6_U51 (.ZN( u1_u11_u6_n107 ) , .A2( u1_u11_u6_n92 ) , .A1( u1_u11_u6_n95 ) );
  AND2_X1 u1_u11_u6_U52 (.ZN( u1_u11_u6_n118 ) , .A2( u1_u11_u6_n91 ) , .A1( u1_u11_u6_n99 ) );
  NAND2_X1 u1_u11_u6_U53 (.ZN( u1_u11_u6_n147 ) , .A2( u1_u11_u6_n98 ) , .A1( u1_u11_u6_n99 ) );
  NAND2_X1 u1_u11_u6_U54 (.ZN( u1_u11_u6_n128 ) , .A1( u1_u11_u6_n94 ) , .A2( u1_u11_u6_n96 ) );
  NAND2_X1 u1_u11_u6_U55 (.ZN( u1_u11_u6_n119 ) , .A2( u1_u11_u6_n95 ) , .A1( u1_u11_u6_n99 ) );
  NAND2_X1 u1_u11_u6_U56 (.ZN( u1_u11_u6_n123 ) , .A2( u1_u11_u6_n91 ) , .A1( u1_u11_u6_n96 ) );
  NAND2_X1 u1_u11_u6_U57 (.ZN( u1_u11_u6_n100 ) , .A2( u1_u11_u6_n92 ) , .A1( u1_u11_u6_n98 ) );
  NAND2_X1 u1_u11_u6_U58 (.ZN( u1_u11_u6_n122 ) , .A1( u1_u11_u6_n94 ) , .A2( u1_u11_u6_n97 ) );
  INV_X1 u1_u11_u6_U59 (.A( u1_u11_u6_n139 ) , .ZN( u1_u11_u6_n160 ) );
  AOI22_X1 u1_u11_u6_U6 (.B2( u1_u11_u6_n101 ) , .A1( u1_u11_u6_n102 ) , .ZN( u1_u11_u6_n103 ) , .B1( u1_u11_u6_n160 ) , .A2( u1_u11_u6_n161 ) );
  NAND2_X1 u1_u11_u6_U60 (.ZN( u1_u11_u6_n113 ) , .A1( u1_u11_u6_n96 ) , .A2( u1_u11_u6_n98 ) );
  NOR2_X1 u1_u11_u6_U61 (.A2( u1_u11_X_40 ) , .A1( u1_u11_X_41 ) , .ZN( u1_u11_u6_n126 ) );
  NOR2_X1 u1_u11_u6_U62 (.A2( u1_u11_X_39 ) , .A1( u1_u11_X_42 ) , .ZN( u1_u11_u6_n92 ) );
  NOR2_X1 u1_u11_u6_U63 (.A2( u1_u11_X_39 ) , .A1( u1_u11_u6_n156 ) , .ZN( u1_u11_u6_n97 ) );
  NOR2_X1 u1_u11_u6_U64 (.A2( u1_u11_X_38 ) , .A1( u1_u11_u6_n165 ) , .ZN( u1_u11_u6_n95 ) );
  NOR2_X1 u1_u11_u6_U65 (.A2( u1_u11_X_41 ) , .ZN( u1_u11_u6_n111 ) , .A1( u1_u11_u6_n157 ) );
  NOR2_X1 u1_u11_u6_U66 (.A2( u1_u11_X_37 ) , .A1( u1_u11_u6_n162 ) , .ZN( u1_u11_u6_n94 ) );
  NOR2_X1 u1_u11_u6_U67 (.A2( u1_u11_X_37 ) , .A1( u1_u11_X_38 ) , .ZN( u1_u11_u6_n91 ) );
  NAND2_X1 u1_u11_u6_U68 (.A1( u1_u11_X_41 ) , .ZN( u1_u11_u6_n144 ) , .A2( u1_u11_u6_n157 ) );
  NAND2_X1 u1_u11_u6_U69 (.A2( u1_u11_X_40 ) , .A1( u1_u11_X_41 ) , .ZN( u1_u11_u6_n139 ) );
  NOR2_X1 u1_u11_u6_U7 (.A1( u1_u11_u6_n118 ) , .ZN( u1_u11_u6_n143 ) , .A2( u1_u11_u6_n168 ) );
  AND2_X1 u1_u11_u6_U70 (.A1( u1_u11_X_39 ) , .A2( u1_u11_u6_n156 ) , .ZN( u1_u11_u6_n96 ) );
  AND2_X1 u1_u11_u6_U71 (.A1( u1_u11_X_39 ) , .A2( u1_u11_X_42 ) , .ZN( u1_u11_u6_n99 ) );
  INV_X1 u1_u11_u6_U72 (.A( u1_u11_X_40 ) , .ZN( u1_u11_u6_n157 ) );
  INV_X1 u1_u11_u6_U73 (.A( u1_u11_X_37 ) , .ZN( u1_u11_u6_n165 ) );
  INV_X1 u1_u11_u6_U74 (.A( u1_u11_X_38 ) , .ZN( u1_u11_u6_n162 ) );
  INV_X1 u1_u11_u6_U75 (.A( u1_u11_X_42 ) , .ZN( u1_u11_u6_n156 ) );
  NAND4_X1 u1_u11_u6_U76 (.ZN( u1_out11_32 ) , .A4( u1_u11_u6_n103 ) , .A3( u1_u11_u6_n104 ) , .A2( u1_u11_u6_n105 ) , .A1( u1_u11_u6_n106 ) );
  AOI22_X1 u1_u11_u6_U77 (.ZN( u1_u11_u6_n105 ) , .A2( u1_u11_u6_n108 ) , .A1( u1_u11_u6_n118 ) , .B2( u1_u11_u6_n126 ) , .B1( u1_u11_u6_n171 ) );
  AOI22_X1 u1_u11_u6_U78 (.ZN( u1_u11_u6_n104 ) , .A1( u1_u11_u6_n111 ) , .B1( u1_u11_u6_n124 ) , .B2( u1_u11_u6_n151 ) , .A2( u1_u11_u6_n93 ) );
  NAND4_X1 u1_u11_u6_U79 (.ZN( u1_out11_12 ) , .A4( u1_u11_u6_n114 ) , .A3( u1_u11_u6_n115 ) , .A2( u1_u11_u6_n116 ) , .A1( u1_u11_u6_n117 ) );
  AOI21_X1 u1_u11_u6_U8 (.B1( u1_u11_u6_n107 ) , .B2( u1_u11_u6_n132 ) , .A( u1_u11_u6_n158 ) , .ZN( u1_u11_u6_n88 ) );
  OAI22_X1 u1_u11_u6_U80 (.B2( u1_u11_u6_n111 ) , .ZN( u1_u11_u6_n116 ) , .B1( u1_u11_u6_n126 ) , .A2( u1_u11_u6_n164 ) , .A1( u1_u11_u6_n167 ) );
  OAI21_X1 u1_u11_u6_U81 (.A( u1_u11_u6_n108 ) , .ZN( u1_u11_u6_n117 ) , .B2( u1_u11_u6_n141 ) , .B1( u1_u11_u6_n163 ) );
  OAI211_X1 u1_u11_u6_U82 (.ZN( u1_out11_7 ) , .B( u1_u11_u6_n153 ) , .C2( u1_u11_u6_n154 ) , .C1( u1_u11_u6_n155 ) , .A( u1_u11_u6_n174 ) );
  NOR3_X1 u1_u11_u6_U83 (.A1( u1_u11_u6_n141 ) , .ZN( u1_u11_u6_n154 ) , .A3( u1_u11_u6_n164 ) , .A2( u1_u11_u6_n171 ) );
  AOI211_X1 u1_u11_u6_U84 (.B( u1_u11_u6_n149 ) , .A( u1_u11_u6_n150 ) , .C2( u1_u11_u6_n151 ) , .C1( u1_u11_u6_n152 ) , .ZN( u1_u11_u6_n153 ) );
  OAI211_X1 u1_u11_u6_U85 (.ZN( u1_out11_22 ) , .B( u1_u11_u6_n137 ) , .A( u1_u11_u6_n138 ) , .C2( u1_u11_u6_n139 ) , .C1( u1_u11_u6_n140 ) );
  AOI22_X1 u1_u11_u6_U86 (.B1( u1_u11_u6_n124 ) , .A2( u1_u11_u6_n125 ) , .A1( u1_u11_u6_n126 ) , .ZN( u1_u11_u6_n138 ) , .B2( u1_u11_u6_n161 ) );
  AND4_X1 u1_u11_u6_U87 (.A3( u1_u11_u6_n119 ) , .A1( u1_u11_u6_n120 ) , .A4( u1_u11_u6_n129 ) , .ZN( u1_u11_u6_n140 ) , .A2( u1_u11_u6_n143 ) );
  NAND3_X1 u1_u11_u6_U88 (.A2( u1_u11_u6_n123 ) , .ZN( u1_u11_u6_n125 ) , .A1( u1_u11_u6_n130 ) , .A3( u1_u11_u6_n131 ) );
  NAND3_X1 u1_u11_u6_U89 (.A3( u1_u11_u6_n133 ) , .ZN( u1_u11_u6_n141 ) , .A1( u1_u11_u6_n145 ) , .A2( u1_u11_u6_n148 ) );
  AOI21_X1 u1_u11_u6_U9 (.B2( u1_u11_u6_n147 ) , .B1( u1_u11_u6_n148 ) , .ZN( u1_u11_u6_n149 ) , .A( u1_u11_u6_n158 ) );
  NAND3_X1 u1_u11_u6_U90 (.ZN( u1_u11_u6_n101 ) , .A3( u1_u11_u6_n107 ) , .A2( u1_u11_u6_n121 ) , .A1( u1_u11_u6_n127 ) );
  NAND3_X1 u1_u11_u6_U91 (.ZN( u1_u11_u6_n102 ) , .A3( u1_u11_u6_n130 ) , .A2( u1_u11_u6_n145 ) , .A1( u1_u11_u6_n166 ) );
  NAND3_X1 u1_u11_u6_U92 (.A3( u1_u11_u6_n113 ) , .A1( u1_u11_u6_n119 ) , .A2( u1_u11_u6_n123 ) , .ZN( u1_u11_u6_n93 ) );
  NAND3_X1 u1_u11_u6_U93 (.ZN( u1_u11_u6_n142 ) , .A2( u1_u11_u6_n172 ) , .A3( u1_u11_u6_n89 ) , .A1( u1_u11_u6_n90 ) );
  AND3_X1 u1_u11_u7_U10 (.A3( u1_u11_u7_n110 ) , .A2( u1_u11_u7_n127 ) , .A1( u1_u11_u7_n132 ) , .ZN( u1_u11_u7_n92 ) );
  OAI21_X1 u1_u11_u7_U11 (.A( u1_u11_u7_n161 ) , .B1( u1_u11_u7_n168 ) , .B2( u1_u11_u7_n173 ) , .ZN( u1_u11_u7_n91 ) );
  AOI211_X1 u1_u11_u7_U12 (.A( u1_u11_u7_n117 ) , .ZN( u1_u11_u7_n118 ) , .C2( u1_u11_u7_n126 ) , .C1( u1_u11_u7_n177 ) , .B( u1_u11_u7_n180 ) );
  OAI22_X1 u1_u11_u7_U13 (.B1( u1_u11_u7_n115 ) , .ZN( u1_u11_u7_n117 ) , .A2( u1_u11_u7_n133 ) , .A1( u1_u11_u7_n137 ) , .B2( u1_u11_u7_n162 ) );
  INV_X1 u1_u11_u7_U14 (.A( u1_u11_u7_n116 ) , .ZN( u1_u11_u7_n180 ) );
  NOR3_X1 u1_u11_u7_U15 (.ZN( u1_u11_u7_n115 ) , .A3( u1_u11_u7_n145 ) , .A2( u1_u11_u7_n168 ) , .A1( u1_u11_u7_n169 ) );
  OAI211_X1 u1_u11_u7_U16 (.B( u1_u11_u7_n122 ) , .A( u1_u11_u7_n123 ) , .C2( u1_u11_u7_n124 ) , .ZN( u1_u11_u7_n154 ) , .C1( u1_u11_u7_n162 ) );
  AOI222_X1 u1_u11_u7_U17 (.ZN( u1_u11_u7_n122 ) , .C2( u1_u11_u7_n126 ) , .C1( u1_u11_u7_n145 ) , .B1( u1_u11_u7_n161 ) , .A2( u1_u11_u7_n165 ) , .B2( u1_u11_u7_n170 ) , .A1( u1_u11_u7_n176 ) );
  INV_X1 u1_u11_u7_U18 (.A( u1_u11_u7_n133 ) , .ZN( u1_u11_u7_n176 ) );
  NOR3_X1 u1_u11_u7_U19 (.A2( u1_u11_u7_n134 ) , .A1( u1_u11_u7_n135 ) , .ZN( u1_u11_u7_n136 ) , .A3( u1_u11_u7_n171 ) );
  NOR2_X1 u1_u11_u7_U20 (.A1( u1_u11_u7_n130 ) , .A2( u1_u11_u7_n134 ) , .ZN( u1_u11_u7_n153 ) );
  INV_X1 u1_u11_u7_U21 (.A( u1_u11_u7_n101 ) , .ZN( u1_u11_u7_n165 ) );
  NOR2_X1 u1_u11_u7_U22 (.ZN( u1_u11_u7_n111 ) , .A2( u1_u11_u7_n134 ) , .A1( u1_u11_u7_n169 ) );
  AOI21_X1 u1_u11_u7_U23 (.ZN( u1_u11_u7_n104 ) , .B2( u1_u11_u7_n112 ) , .B1( u1_u11_u7_n127 ) , .A( u1_u11_u7_n164 ) );
  AOI21_X1 u1_u11_u7_U24 (.ZN( u1_u11_u7_n106 ) , .B1( u1_u11_u7_n133 ) , .B2( u1_u11_u7_n146 ) , .A( u1_u11_u7_n162 ) );
  AOI21_X1 u1_u11_u7_U25 (.A( u1_u11_u7_n101 ) , .ZN( u1_u11_u7_n107 ) , .B2( u1_u11_u7_n128 ) , .B1( u1_u11_u7_n175 ) );
  INV_X1 u1_u11_u7_U26 (.A( u1_u11_u7_n138 ) , .ZN( u1_u11_u7_n171 ) );
  INV_X1 u1_u11_u7_U27 (.A( u1_u11_u7_n131 ) , .ZN( u1_u11_u7_n177 ) );
  INV_X1 u1_u11_u7_U28 (.A( u1_u11_u7_n110 ) , .ZN( u1_u11_u7_n174 ) );
  NAND2_X1 u1_u11_u7_U29 (.A1( u1_u11_u7_n129 ) , .A2( u1_u11_u7_n132 ) , .ZN( u1_u11_u7_n149 ) );
  OAI21_X1 u1_u11_u7_U3 (.ZN( u1_u11_u7_n159 ) , .A( u1_u11_u7_n165 ) , .B2( u1_u11_u7_n171 ) , .B1( u1_u11_u7_n174 ) );
  NAND2_X1 u1_u11_u7_U30 (.A1( u1_u11_u7_n113 ) , .A2( u1_u11_u7_n124 ) , .ZN( u1_u11_u7_n130 ) );
  INV_X1 u1_u11_u7_U31 (.A( u1_u11_u7_n112 ) , .ZN( u1_u11_u7_n173 ) );
  INV_X1 u1_u11_u7_U32 (.A( u1_u11_u7_n128 ) , .ZN( u1_u11_u7_n168 ) );
  INV_X1 u1_u11_u7_U33 (.A( u1_u11_u7_n148 ) , .ZN( u1_u11_u7_n169 ) );
  INV_X1 u1_u11_u7_U34 (.A( u1_u11_u7_n127 ) , .ZN( u1_u11_u7_n179 ) );
  NOR2_X1 u1_u11_u7_U35 (.ZN( u1_u11_u7_n101 ) , .A2( u1_u11_u7_n150 ) , .A1( u1_u11_u7_n156 ) );
  AOI211_X1 u1_u11_u7_U36 (.B( u1_u11_u7_n154 ) , .A( u1_u11_u7_n155 ) , .C1( u1_u11_u7_n156 ) , .ZN( u1_u11_u7_n157 ) , .C2( u1_u11_u7_n172 ) );
  INV_X1 u1_u11_u7_U37 (.A( u1_u11_u7_n153 ) , .ZN( u1_u11_u7_n172 ) );
  AOI211_X1 u1_u11_u7_U38 (.B( u1_u11_u7_n139 ) , .A( u1_u11_u7_n140 ) , .C2( u1_u11_u7_n141 ) , .ZN( u1_u11_u7_n142 ) , .C1( u1_u11_u7_n156 ) );
  AOI21_X1 u1_u11_u7_U39 (.A( u1_u11_u7_n137 ) , .B1( u1_u11_u7_n138 ) , .ZN( u1_u11_u7_n139 ) , .B2( u1_u11_u7_n146 ) );
  INV_X1 u1_u11_u7_U4 (.A( u1_u11_u7_n111 ) , .ZN( u1_u11_u7_n170 ) );
  NAND4_X1 u1_u11_u7_U40 (.A3( u1_u11_u7_n127 ) , .A2( u1_u11_u7_n128 ) , .A1( u1_u11_u7_n129 ) , .ZN( u1_u11_u7_n141 ) , .A4( u1_u11_u7_n147 ) );
  OAI22_X1 u1_u11_u7_U41 (.B1( u1_u11_u7_n136 ) , .ZN( u1_u11_u7_n140 ) , .A1( u1_u11_u7_n153 ) , .B2( u1_u11_u7_n162 ) , .A2( u1_u11_u7_n164 ) );
  AOI21_X1 u1_u11_u7_U42 (.ZN( u1_u11_u7_n123 ) , .B1( u1_u11_u7_n165 ) , .B2( u1_u11_u7_n177 ) , .A( u1_u11_u7_n97 ) );
  AOI21_X1 u1_u11_u7_U43 (.B2( u1_u11_u7_n113 ) , .B1( u1_u11_u7_n124 ) , .A( u1_u11_u7_n125 ) , .ZN( u1_u11_u7_n97 ) );
  INV_X1 u1_u11_u7_U44 (.A( u1_u11_u7_n125 ) , .ZN( u1_u11_u7_n161 ) );
  INV_X1 u1_u11_u7_U45 (.A( u1_u11_u7_n152 ) , .ZN( u1_u11_u7_n162 ) );
  AOI22_X1 u1_u11_u7_U46 (.A2( u1_u11_u7_n114 ) , .ZN( u1_u11_u7_n119 ) , .B1( u1_u11_u7_n130 ) , .A1( u1_u11_u7_n156 ) , .B2( u1_u11_u7_n165 ) );
  NAND2_X1 u1_u11_u7_U47 (.A2( u1_u11_u7_n112 ) , .ZN( u1_u11_u7_n114 ) , .A1( u1_u11_u7_n175 ) );
  AND2_X1 u1_u11_u7_U48 (.ZN( u1_u11_u7_n145 ) , .A2( u1_u11_u7_n98 ) , .A1( u1_u11_u7_n99 ) );
  NOR2_X1 u1_u11_u7_U49 (.ZN( u1_u11_u7_n137 ) , .A1( u1_u11_u7_n150 ) , .A2( u1_u11_u7_n161 ) );
  INV_X1 u1_u11_u7_U5 (.A( u1_u11_u7_n149 ) , .ZN( u1_u11_u7_n175 ) );
  AOI21_X1 u1_u11_u7_U50 (.ZN( u1_u11_u7_n105 ) , .B2( u1_u11_u7_n110 ) , .A( u1_u11_u7_n125 ) , .B1( u1_u11_u7_n147 ) );
  NAND2_X1 u1_u11_u7_U51 (.ZN( u1_u11_u7_n146 ) , .A1( u1_u11_u7_n95 ) , .A2( u1_u11_u7_n98 ) );
  NAND2_X1 u1_u11_u7_U52 (.A2( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n147 ) , .A1( u1_u11_u7_n93 ) );
  NAND2_X1 u1_u11_u7_U53 (.A1( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n127 ) , .A2( u1_u11_u7_n99 ) );
  OR2_X1 u1_u11_u7_U54 (.ZN( u1_u11_u7_n126 ) , .A2( u1_u11_u7_n152 ) , .A1( u1_u11_u7_n156 ) );
  NAND2_X1 u1_u11_u7_U55 (.A2( u1_u11_u7_n102 ) , .A1( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n133 ) );
  NAND2_X1 u1_u11_u7_U56 (.ZN( u1_u11_u7_n112 ) , .A2( u1_u11_u7_n96 ) , .A1( u1_u11_u7_n99 ) );
  NAND2_X1 u1_u11_u7_U57 (.A2( u1_u11_u7_n102 ) , .ZN( u1_u11_u7_n128 ) , .A1( u1_u11_u7_n98 ) );
  NAND2_X1 u1_u11_u7_U58 (.A1( u1_u11_u7_n100 ) , .ZN( u1_u11_u7_n113 ) , .A2( u1_u11_u7_n93 ) );
  NAND2_X1 u1_u11_u7_U59 (.A2( u1_u11_u7_n102 ) , .ZN( u1_u11_u7_n124 ) , .A1( u1_u11_u7_n96 ) );
  INV_X1 u1_u11_u7_U6 (.A( u1_u11_u7_n154 ) , .ZN( u1_u11_u7_n178 ) );
  NAND2_X1 u1_u11_u7_U60 (.ZN( u1_u11_u7_n110 ) , .A1( u1_u11_u7_n95 ) , .A2( u1_u11_u7_n96 ) );
  INV_X1 u1_u11_u7_U61 (.A( u1_u11_u7_n150 ) , .ZN( u1_u11_u7_n164 ) );
  AND2_X1 u1_u11_u7_U62 (.ZN( u1_u11_u7_n134 ) , .A1( u1_u11_u7_n93 ) , .A2( u1_u11_u7_n98 ) );
  NAND2_X1 u1_u11_u7_U63 (.A1( u1_u11_u7_n100 ) , .A2( u1_u11_u7_n102 ) , .ZN( u1_u11_u7_n129 ) );
  NAND2_X1 u1_u11_u7_U64 (.A2( u1_u11_u7_n103 ) , .ZN( u1_u11_u7_n131 ) , .A1( u1_u11_u7_n95 ) );
  NAND2_X1 u1_u11_u7_U65 (.A1( u1_u11_u7_n100 ) , .ZN( u1_u11_u7_n138 ) , .A2( u1_u11_u7_n99 ) );
  NAND2_X1 u1_u11_u7_U66 (.ZN( u1_u11_u7_n132 ) , .A1( u1_u11_u7_n93 ) , .A2( u1_u11_u7_n96 ) );
  NAND2_X1 u1_u11_u7_U67 (.A1( u1_u11_u7_n100 ) , .ZN( u1_u11_u7_n148 ) , .A2( u1_u11_u7_n95 ) );
  NOR2_X1 u1_u11_u7_U68 (.A2( u1_u11_X_47 ) , .ZN( u1_u11_u7_n150 ) , .A1( u1_u11_u7_n163 ) );
  NOR2_X1 u1_u11_u7_U69 (.A2( u1_u11_X_43 ) , .A1( u1_u11_X_44 ) , .ZN( u1_u11_u7_n103 ) );
  AOI211_X1 u1_u11_u7_U7 (.ZN( u1_u11_u7_n116 ) , .A( u1_u11_u7_n155 ) , .C1( u1_u11_u7_n161 ) , .C2( u1_u11_u7_n171 ) , .B( u1_u11_u7_n94 ) );
  NOR2_X1 u1_u11_u7_U70 (.A2( u1_u11_X_48 ) , .A1( u1_u11_u7_n166 ) , .ZN( u1_u11_u7_n95 ) );
  NOR2_X1 u1_u11_u7_U71 (.A2( u1_u11_X_45 ) , .A1( u1_u11_X_48 ) , .ZN( u1_u11_u7_n99 ) );
  NOR2_X1 u1_u11_u7_U72 (.A2( u1_u11_X_44 ) , .A1( u1_u11_u7_n167 ) , .ZN( u1_u11_u7_n98 ) );
  NOR2_X1 u1_u11_u7_U73 (.A2( u1_u11_X_46 ) , .A1( u1_u11_X_47 ) , .ZN( u1_u11_u7_n152 ) );
  AND2_X1 u1_u11_u7_U74 (.A1( u1_u11_X_47 ) , .ZN( u1_u11_u7_n156 ) , .A2( u1_u11_u7_n163 ) );
  NAND2_X1 u1_u11_u7_U75 (.A2( u1_u11_X_46 ) , .A1( u1_u11_X_47 ) , .ZN( u1_u11_u7_n125 ) );
  AND2_X1 u1_u11_u7_U76 (.A2( u1_u11_X_45 ) , .A1( u1_u11_X_48 ) , .ZN( u1_u11_u7_n102 ) );
  AND2_X1 u1_u11_u7_U77 (.A2( u1_u11_X_43 ) , .A1( u1_u11_X_44 ) , .ZN( u1_u11_u7_n96 ) );
  AND2_X1 u1_u11_u7_U78 (.A1( u1_u11_X_44 ) , .ZN( u1_u11_u7_n100 ) , .A2( u1_u11_u7_n167 ) );
  AND2_X1 u1_u11_u7_U79 (.A1( u1_u11_X_48 ) , .A2( u1_u11_u7_n166 ) , .ZN( u1_u11_u7_n93 ) );
  OAI222_X1 u1_u11_u7_U8 (.C2( u1_u11_u7_n101 ) , .B2( u1_u11_u7_n111 ) , .A1( u1_u11_u7_n113 ) , .C1( u1_u11_u7_n146 ) , .A2( u1_u11_u7_n162 ) , .B1( u1_u11_u7_n164 ) , .ZN( u1_u11_u7_n94 ) );
  INV_X1 u1_u11_u7_U80 (.A( u1_u11_X_46 ) , .ZN( u1_u11_u7_n163 ) );
  INV_X1 u1_u11_u7_U81 (.A( u1_u11_X_43 ) , .ZN( u1_u11_u7_n167 ) );
  INV_X1 u1_u11_u7_U82 (.A( u1_u11_X_45 ) , .ZN( u1_u11_u7_n166 ) );
  NAND4_X1 u1_u11_u7_U83 (.ZN( u1_out11_5 ) , .A4( u1_u11_u7_n108 ) , .A3( u1_u11_u7_n109 ) , .A1( u1_u11_u7_n116 ) , .A2( u1_u11_u7_n123 ) );
  AOI22_X1 u1_u11_u7_U84 (.ZN( u1_u11_u7_n109 ) , .A2( u1_u11_u7_n126 ) , .B2( u1_u11_u7_n145 ) , .B1( u1_u11_u7_n156 ) , .A1( u1_u11_u7_n171 ) );
  NOR4_X1 u1_u11_u7_U85 (.A4( u1_u11_u7_n104 ) , .A3( u1_u11_u7_n105 ) , .A2( u1_u11_u7_n106 ) , .A1( u1_u11_u7_n107 ) , .ZN( u1_u11_u7_n108 ) );
  NAND4_X1 u1_u11_u7_U86 (.ZN( u1_out11_27 ) , .A4( u1_u11_u7_n118 ) , .A3( u1_u11_u7_n119 ) , .A2( u1_u11_u7_n120 ) , .A1( u1_u11_u7_n121 ) );
  OAI21_X1 u1_u11_u7_U87 (.ZN( u1_u11_u7_n121 ) , .B2( u1_u11_u7_n145 ) , .A( u1_u11_u7_n150 ) , .B1( u1_u11_u7_n174 ) );
  OAI21_X1 u1_u11_u7_U88 (.ZN( u1_u11_u7_n120 ) , .A( u1_u11_u7_n161 ) , .B2( u1_u11_u7_n170 ) , .B1( u1_u11_u7_n179 ) );
  NAND4_X1 u1_u11_u7_U89 (.ZN( u1_out11_21 ) , .A4( u1_u11_u7_n157 ) , .A3( u1_u11_u7_n158 ) , .A2( u1_u11_u7_n159 ) , .A1( u1_u11_u7_n160 ) );
  OAI221_X1 u1_u11_u7_U9 (.C1( u1_u11_u7_n101 ) , .C2( u1_u11_u7_n147 ) , .ZN( u1_u11_u7_n155 ) , .B2( u1_u11_u7_n162 ) , .A( u1_u11_u7_n91 ) , .B1( u1_u11_u7_n92 ) );
  OAI21_X1 u1_u11_u7_U90 (.B1( u1_u11_u7_n145 ) , .ZN( u1_u11_u7_n160 ) , .A( u1_u11_u7_n161 ) , .B2( u1_u11_u7_n177 ) );
  AOI22_X1 u1_u11_u7_U91 (.B2( u1_u11_u7_n149 ) , .B1( u1_u11_u7_n150 ) , .A2( u1_u11_u7_n151 ) , .A1( u1_u11_u7_n152 ) , .ZN( u1_u11_u7_n158 ) );
  NAND4_X1 u1_u11_u7_U92 (.ZN( u1_out11_15 ) , .A4( u1_u11_u7_n142 ) , .A3( u1_u11_u7_n143 ) , .A2( u1_u11_u7_n144 ) , .A1( u1_u11_u7_n178 ) );
  OR2_X1 u1_u11_u7_U93 (.A2( u1_u11_u7_n125 ) , .A1( u1_u11_u7_n129 ) , .ZN( u1_u11_u7_n144 ) );
  AOI22_X1 u1_u11_u7_U94 (.A2( u1_u11_u7_n126 ) , .ZN( u1_u11_u7_n143 ) , .B2( u1_u11_u7_n165 ) , .B1( u1_u11_u7_n173 ) , .A1( u1_u11_u7_n174 ) );
  NAND3_X1 u1_u11_u7_U95 (.A3( u1_u11_u7_n146 ) , .A2( u1_u11_u7_n147 ) , .A1( u1_u11_u7_n148 ) , .ZN( u1_u11_u7_n151 ) );
  NAND3_X1 u1_u11_u7_U96 (.A3( u1_u11_u7_n131 ) , .A2( u1_u11_u7_n132 ) , .A1( u1_u11_u7_n133 ) , .ZN( u1_u11_u7_n135 ) );
  XOR2_X1 u1_u13_U1 (.B( u1_K14_9 ) , .A( u1_R12_6 ) , .Z( u1_u13_X_9 ) );
  XOR2_X1 u1_u13_U16 (.B( u1_K14_3 ) , .A( u1_R12_2 ) , .Z( u1_u13_X_3 ) );
  XOR2_X1 u1_u13_U2 (.B( u1_K14_8 ) , .A( u1_R12_5 ) , .Z( u1_u13_X_8 ) );
  XOR2_X1 u1_u13_U27 (.B( u1_K14_2 ) , .A( u1_R12_1 ) , .Z( u1_u13_X_2 ) );
  XOR2_X1 u1_u13_U3 (.B( u1_K14_7 ) , .A( u1_R12_4 ) , .Z( u1_u13_X_7 ) );
  XOR2_X1 u1_u13_U38 (.B( u1_K14_1 ) , .A( u1_R12_32 ) , .Z( u1_u13_X_1 ) );
  XOR2_X1 u1_u13_U4 (.B( u1_K14_6 ) , .A( u1_R12_5 ) , .Z( u1_u13_X_6 ) );
  XOR2_X1 u1_u13_U40 (.B( u1_K14_18 ) , .A( u1_R12_13 ) , .Z( u1_u13_X_18 ) );
  XOR2_X1 u1_u13_U41 (.B( u1_K14_17 ) , .A( u1_R12_12 ) , .Z( u1_u13_X_17 ) );
  XOR2_X1 u1_u13_U42 (.B( u1_K14_16 ) , .A( u1_R12_11 ) , .Z( u1_u13_X_16 ) );
  XOR2_X1 u1_u13_U43 (.B( u1_K14_15 ) , .A( u1_R12_10 ) , .Z( u1_u13_X_15 ) );
  XOR2_X1 u1_u13_U44 (.B( u1_K14_14 ) , .A( u1_R12_9 ) , .Z( u1_u13_X_14 ) );
  XOR2_X1 u1_u13_U45 (.B( u1_K14_13 ) , .A( u1_R12_8 ) , .Z( u1_u13_X_13 ) );
  XOR2_X1 u1_u13_U46 (.B( u1_K14_12 ) , .A( u1_R12_9 ) , .Z( u1_u13_X_12 ) );
  XOR2_X1 u1_u13_U47 (.B( u1_K14_11 ) , .A( u1_R12_8 ) , .Z( u1_u13_X_11 ) );
  XOR2_X1 u1_u13_U48 (.B( u1_K14_10 ) , .A( u1_R12_7 ) , .Z( u1_u13_X_10 ) );
  XOR2_X1 u1_u13_U5 (.B( u1_K14_5 ) , .A( u1_R12_4 ) , .Z( u1_u13_X_5 ) );
  XOR2_X1 u1_u13_U6 (.B( u1_K14_4 ) , .A( u1_R12_3 ) , .Z( u1_u13_X_4 ) );
  AND3_X1 u1_u13_u0_U10 (.A2( u1_u13_u0_n112 ) , .ZN( u1_u13_u0_n127 ) , .A3( u1_u13_u0_n130 ) , .A1( u1_u13_u0_n148 ) );
  NAND2_X1 u1_u13_u0_U11 (.ZN( u1_u13_u0_n113 ) , .A1( u1_u13_u0_n139 ) , .A2( u1_u13_u0_n149 ) );
  AND2_X1 u1_u13_u0_U12 (.ZN( u1_u13_u0_n107 ) , .A1( u1_u13_u0_n130 ) , .A2( u1_u13_u0_n140 ) );
  AND2_X1 u1_u13_u0_U13 (.A2( u1_u13_u0_n129 ) , .A1( u1_u13_u0_n130 ) , .ZN( u1_u13_u0_n151 ) );
  AND2_X1 u1_u13_u0_U14 (.A1( u1_u13_u0_n108 ) , .A2( u1_u13_u0_n125 ) , .ZN( u1_u13_u0_n145 ) );
  INV_X1 u1_u13_u0_U15 (.A( u1_u13_u0_n143 ) , .ZN( u1_u13_u0_n173 ) );
  NOR2_X1 u1_u13_u0_U16 (.A2( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n147 ) , .A1( u1_u13_u0_n160 ) );
  INV_X1 u1_u13_u0_U17 (.ZN( u1_u13_u0_n172 ) , .A( u1_u13_u0_n88 ) );
  OAI222_X1 u1_u13_u0_U18 (.C1( u1_u13_u0_n108 ) , .A1( u1_u13_u0_n125 ) , .B2( u1_u13_u0_n128 ) , .B1( u1_u13_u0_n144 ) , .A2( u1_u13_u0_n158 ) , .C2( u1_u13_u0_n161 ) , .ZN( u1_u13_u0_n88 ) );
  NOR2_X1 u1_u13_u0_U19 (.A1( u1_u13_u0_n163 ) , .A2( u1_u13_u0_n164 ) , .ZN( u1_u13_u0_n95 ) );
  AOI21_X1 u1_u13_u0_U20 (.B1( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n132 ) , .A( u1_u13_u0_n165 ) , .B2( u1_u13_u0_n93 ) );
  INV_X1 u1_u13_u0_U21 (.A( u1_u13_u0_n142 ) , .ZN( u1_u13_u0_n165 ) );
  OAI221_X1 u1_u13_u0_U22 (.C1( u1_u13_u0_n121 ) , .ZN( u1_u13_u0_n122 ) , .B2( u1_u13_u0_n127 ) , .A( u1_u13_u0_n143 ) , .B1( u1_u13_u0_n144 ) , .C2( u1_u13_u0_n147 ) );
  OAI22_X1 u1_u13_u0_U23 (.B1( u1_u13_u0_n125 ) , .ZN( u1_u13_u0_n126 ) , .A1( u1_u13_u0_n138 ) , .A2( u1_u13_u0_n146 ) , .B2( u1_u13_u0_n147 ) );
  OAI22_X1 u1_u13_u0_U24 (.B1( u1_u13_u0_n131 ) , .A1( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n147 ) , .A2( u1_u13_u0_n90 ) , .ZN( u1_u13_u0_n91 ) );
  AND3_X1 u1_u13_u0_U25 (.A3( u1_u13_u0_n121 ) , .A2( u1_u13_u0_n125 ) , .A1( u1_u13_u0_n148 ) , .ZN( u1_u13_u0_n90 ) );
  INV_X1 u1_u13_u0_U26 (.A( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n161 ) );
  NOR2_X1 u1_u13_u0_U27 (.A1( u1_u13_u0_n120 ) , .ZN( u1_u13_u0_n143 ) , .A2( u1_u13_u0_n167 ) );
  OAI221_X1 u1_u13_u0_U28 (.C1( u1_u13_u0_n112 ) , .ZN( u1_u13_u0_n120 ) , .B1( u1_u13_u0_n138 ) , .B2( u1_u13_u0_n141 ) , .C2( u1_u13_u0_n147 ) , .A( u1_u13_u0_n172 ) );
  AOI211_X1 u1_u13_u0_U29 (.B( u1_u13_u0_n115 ) , .A( u1_u13_u0_n116 ) , .C2( u1_u13_u0_n117 ) , .C1( u1_u13_u0_n118 ) , .ZN( u1_u13_u0_n119 ) );
  INV_X1 u1_u13_u0_U3 (.A( u1_u13_u0_n113 ) , .ZN( u1_u13_u0_n166 ) );
  AOI22_X1 u1_u13_u0_U30 (.B2( u1_u13_u0_n109 ) , .A2( u1_u13_u0_n110 ) , .ZN( u1_u13_u0_n111 ) , .B1( u1_u13_u0_n118 ) , .A1( u1_u13_u0_n160 ) );
  INV_X1 u1_u13_u0_U31 (.A( u1_u13_u0_n118 ) , .ZN( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U32 (.ZN( u1_u13_u0_n104 ) , .B1( u1_u13_u0_n107 ) , .B2( u1_u13_u0_n141 ) , .A( u1_u13_u0_n144 ) );
  AOI21_X1 u1_u13_u0_U33 (.B1( u1_u13_u0_n127 ) , .B2( u1_u13_u0_n129 ) , .A( u1_u13_u0_n138 ) , .ZN( u1_u13_u0_n96 ) );
  AOI21_X1 u1_u13_u0_U34 (.ZN( u1_u13_u0_n116 ) , .B2( u1_u13_u0_n142 ) , .A( u1_u13_u0_n144 ) , .B1( u1_u13_u0_n166 ) );
  NAND2_X1 u1_u13_u0_U35 (.A1( u1_u13_u0_n100 ) , .A2( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n125 ) );
  NAND2_X1 u1_u13_u0_U36 (.A1( u1_u13_u0_n101 ) , .A2( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n150 ) );
  INV_X1 u1_u13_u0_U37 (.A( u1_u13_u0_n138 ) , .ZN( u1_u13_u0_n160 ) );
  NAND2_X1 u1_u13_u0_U38 (.A1( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n128 ) , .A2( u1_u13_u0_n95 ) );
  NAND2_X1 u1_u13_u0_U39 (.A1( u1_u13_u0_n100 ) , .ZN( u1_u13_u0_n129 ) , .A2( u1_u13_u0_n95 ) );
  AOI21_X1 u1_u13_u0_U4 (.B1( u1_u13_u0_n114 ) , .ZN( u1_u13_u0_n115 ) , .B2( u1_u13_u0_n129 ) , .A( u1_u13_u0_n161 ) );
  NAND2_X1 u1_u13_u0_U40 (.A2( u1_u13_u0_n100 ) , .ZN( u1_u13_u0_n131 ) , .A1( u1_u13_u0_n92 ) );
  NAND2_X1 u1_u13_u0_U41 (.A2( u1_u13_u0_n100 ) , .A1( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n139 ) );
  NAND2_X1 u1_u13_u0_U42 (.ZN( u1_u13_u0_n148 ) , .A1( u1_u13_u0_n93 ) , .A2( u1_u13_u0_n95 ) );
  NAND2_X1 u1_u13_u0_U43 (.A2( u1_u13_u0_n102 ) , .A1( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n149 ) );
  NAND2_X1 u1_u13_u0_U44 (.A2( u1_u13_u0_n102 ) , .ZN( u1_u13_u0_n114 ) , .A1( u1_u13_u0_n92 ) );
  NAND2_X1 u1_u13_u0_U45 (.A2( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n121 ) , .A1( u1_u13_u0_n93 ) );
  NAND2_X1 u1_u13_u0_U46 (.ZN( u1_u13_u0_n112 ) , .A2( u1_u13_u0_n92 ) , .A1( u1_u13_u0_n93 ) );
  OR3_X1 u1_u13_u0_U47 (.A3( u1_u13_u0_n152 ) , .A2( u1_u13_u0_n153 ) , .A1( u1_u13_u0_n154 ) , .ZN( u1_u13_u0_n155 ) );
  AOI21_X1 u1_u13_u0_U48 (.B2( u1_u13_u0_n150 ) , .B1( u1_u13_u0_n151 ) , .ZN( u1_u13_u0_n152 ) , .A( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U49 (.A( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n145 ) , .B1( u1_u13_u0_n146 ) , .ZN( u1_u13_u0_n154 ) );
  AOI21_X1 u1_u13_u0_U5 (.B2( u1_u13_u0_n131 ) , .ZN( u1_u13_u0_n134 ) , .B1( u1_u13_u0_n151 ) , .A( u1_u13_u0_n158 ) );
  AOI21_X1 u1_u13_u0_U50 (.A( u1_u13_u0_n147 ) , .B2( u1_u13_u0_n148 ) , .B1( u1_u13_u0_n149 ) , .ZN( u1_u13_u0_n153 ) );
  INV_X1 u1_u13_u0_U51 (.ZN( u1_u13_u0_n171 ) , .A( u1_u13_u0_n99 ) );
  OAI211_X1 u1_u13_u0_U52 (.C2( u1_u13_u0_n140 ) , .C1( u1_u13_u0_n161 ) , .A( u1_u13_u0_n169 ) , .B( u1_u13_u0_n98 ) , .ZN( u1_u13_u0_n99 ) );
  AOI211_X1 u1_u13_u0_U53 (.C1( u1_u13_u0_n118 ) , .A( u1_u13_u0_n123 ) , .B( u1_u13_u0_n96 ) , .C2( u1_u13_u0_n97 ) , .ZN( u1_u13_u0_n98 ) );
  INV_X1 u1_u13_u0_U54 (.ZN( u1_u13_u0_n169 ) , .A( u1_u13_u0_n91 ) );
  NOR2_X1 u1_u13_u0_U55 (.A2( u1_u13_X_6 ) , .ZN( u1_u13_u0_n100 ) , .A1( u1_u13_u0_n162 ) );
  NOR2_X1 u1_u13_u0_U56 (.A2( u1_u13_X_4 ) , .A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n118 ) );
  NOR2_X1 u1_u13_u0_U57 (.A2( u1_u13_X_2 ) , .ZN( u1_u13_u0_n103 ) , .A1( u1_u13_u0_n164 ) );
  NOR2_X1 u1_u13_u0_U58 (.A2( u1_u13_X_1 ) , .A1( u1_u13_X_2 ) , .ZN( u1_u13_u0_n92 ) );
  NOR2_X1 u1_u13_u0_U59 (.A2( u1_u13_X_1 ) , .ZN( u1_u13_u0_n101 ) , .A1( u1_u13_u0_n163 ) );
  NOR2_X1 u1_u13_u0_U6 (.A1( u1_u13_u0_n108 ) , .ZN( u1_u13_u0_n123 ) , .A2( u1_u13_u0_n158 ) );
  NAND2_X1 u1_u13_u0_U60 (.A2( u1_u13_X_4 ) , .A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n144 ) );
  NOR2_X1 u1_u13_u0_U61 (.A2( u1_u13_X_5 ) , .ZN( u1_u13_u0_n136 ) , .A1( u1_u13_u0_n159 ) );
  NAND2_X1 u1_u13_u0_U62 (.A1( u1_u13_X_5 ) , .ZN( u1_u13_u0_n138 ) , .A2( u1_u13_u0_n159 ) );
  AND2_X1 u1_u13_u0_U63 (.A2( u1_u13_X_3 ) , .A1( u1_u13_X_6 ) , .ZN( u1_u13_u0_n102 ) );
  AND2_X1 u1_u13_u0_U64 (.A1( u1_u13_X_6 ) , .A2( u1_u13_u0_n162 ) , .ZN( u1_u13_u0_n93 ) );
  INV_X1 u1_u13_u0_U65 (.A( u1_u13_X_4 ) , .ZN( u1_u13_u0_n159 ) );
  INV_X1 u1_u13_u0_U66 (.A( u1_u13_X_1 ) , .ZN( u1_u13_u0_n164 ) );
  INV_X1 u1_u13_u0_U67 (.A( u1_u13_X_2 ) , .ZN( u1_u13_u0_n163 ) );
  INV_X1 u1_u13_u0_U68 (.A( u1_u13_u0_n126 ) , .ZN( u1_u13_u0_n168 ) );
  AOI211_X1 u1_u13_u0_U69 (.B( u1_u13_u0_n133 ) , .A( u1_u13_u0_n134 ) , .C2( u1_u13_u0_n135 ) , .C1( u1_u13_u0_n136 ) , .ZN( u1_u13_u0_n137 ) );
  OAI21_X1 u1_u13_u0_U7 (.B1( u1_u13_u0_n150 ) , .B2( u1_u13_u0_n158 ) , .A( u1_u13_u0_n172 ) , .ZN( u1_u13_u0_n89 ) );
  INV_X1 u1_u13_u0_U70 (.ZN( u1_u13_u0_n174 ) , .A( u1_u13_u0_n89 ) );
  AOI211_X1 u1_u13_u0_U71 (.B( u1_u13_u0_n104 ) , .A( u1_u13_u0_n105 ) , .ZN( u1_u13_u0_n106 ) , .C2( u1_u13_u0_n113 ) , .C1( u1_u13_u0_n160 ) );
  OR4_X1 u1_u13_u0_U72 (.ZN( u1_out13_17 ) , .A4( u1_u13_u0_n122 ) , .A2( u1_u13_u0_n123 ) , .A1( u1_u13_u0_n124 ) , .A3( u1_u13_u0_n170 ) );
  AOI21_X1 u1_u13_u0_U73 (.B2( u1_u13_u0_n107 ) , .ZN( u1_u13_u0_n124 ) , .B1( u1_u13_u0_n128 ) , .A( u1_u13_u0_n161 ) );
  INV_X1 u1_u13_u0_U74 (.A( u1_u13_u0_n111 ) , .ZN( u1_u13_u0_n170 ) );
  OR4_X1 u1_u13_u0_U75 (.ZN( u1_out13_31 ) , .A4( u1_u13_u0_n155 ) , .A2( u1_u13_u0_n156 ) , .A1( u1_u13_u0_n157 ) , .A3( u1_u13_u0_n173 ) );
  AOI21_X1 u1_u13_u0_U76 (.A( u1_u13_u0_n138 ) , .B2( u1_u13_u0_n139 ) , .B1( u1_u13_u0_n140 ) , .ZN( u1_u13_u0_n157 ) );
  AOI21_X1 u1_u13_u0_U77 (.B2( u1_u13_u0_n141 ) , .B1( u1_u13_u0_n142 ) , .ZN( u1_u13_u0_n156 ) , .A( u1_u13_u0_n161 ) );
  AOI21_X1 u1_u13_u0_U78 (.B1( u1_u13_u0_n132 ) , .ZN( u1_u13_u0_n133 ) , .A( u1_u13_u0_n144 ) , .B2( u1_u13_u0_n166 ) );
  OAI22_X1 u1_u13_u0_U79 (.ZN( u1_u13_u0_n105 ) , .A2( u1_u13_u0_n132 ) , .B1( u1_u13_u0_n146 ) , .A1( u1_u13_u0_n147 ) , .B2( u1_u13_u0_n161 ) );
  AND2_X1 u1_u13_u0_U8 (.A1( u1_u13_u0_n114 ) , .A2( u1_u13_u0_n121 ) , .ZN( u1_u13_u0_n146 ) );
  NAND2_X1 u1_u13_u0_U80 (.ZN( u1_u13_u0_n110 ) , .A2( u1_u13_u0_n132 ) , .A1( u1_u13_u0_n145 ) );
  INV_X1 u1_u13_u0_U81 (.A( u1_u13_u0_n119 ) , .ZN( u1_u13_u0_n167 ) );
  NAND2_X1 u1_u13_u0_U82 (.A2( u1_u13_u0_n103 ) , .ZN( u1_u13_u0_n140 ) , .A1( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U83 (.A1( u1_u13_u0_n101 ) , .ZN( u1_u13_u0_n130 ) , .A2( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U84 (.ZN( u1_u13_u0_n108 ) , .A1( u1_u13_u0_n92 ) , .A2( u1_u13_u0_n94 ) );
  NAND2_X1 u1_u13_u0_U85 (.ZN( u1_u13_u0_n142 ) , .A1( u1_u13_u0_n94 ) , .A2( u1_u13_u0_n95 ) );
  INV_X1 u1_u13_u0_U86 (.A( u1_u13_X_3 ) , .ZN( u1_u13_u0_n162 ) );
  NOR2_X1 u1_u13_u0_U87 (.A2( u1_u13_X_3 ) , .A1( u1_u13_X_6 ) , .ZN( u1_u13_u0_n94 ) );
  NAND3_X1 u1_u13_u0_U88 (.ZN( u1_out13_23 ) , .A3( u1_u13_u0_n137 ) , .A1( u1_u13_u0_n168 ) , .A2( u1_u13_u0_n171 ) );
  NAND3_X1 u1_u13_u0_U89 (.A3( u1_u13_u0_n127 ) , .A2( u1_u13_u0_n128 ) , .ZN( u1_u13_u0_n135 ) , .A1( u1_u13_u0_n150 ) );
  AND2_X1 u1_u13_u0_U9 (.A1( u1_u13_u0_n131 ) , .ZN( u1_u13_u0_n141 ) , .A2( u1_u13_u0_n150 ) );
  NAND3_X1 u1_u13_u0_U90 (.ZN( u1_u13_u0_n117 ) , .A3( u1_u13_u0_n132 ) , .A2( u1_u13_u0_n139 ) , .A1( u1_u13_u0_n148 ) );
  NAND3_X1 u1_u13_u0_U91 (.ZN( u1_u13_u0_n109 ) , .A2( u1_u13_u0_n114 ) , .A3( u1_u13_u0_n140 ) , .A1( u1_u13_u0_n149 ) );
  NAND3_X1 u1_u13_u0_U92 (.ZN( u1_out13_9 ) , .A3( u1_u13_u0_n106 ) , .A2( u1_u13_u0_n171 ) , .A1( u1_u13_u0_n174 ) );
  NAND3_X1 u1_u13_u0_U93 (.A2( u1_u13_u0_n128 ) , .A1( u1_u13_u0_n132 ) , .A3( u1_u13_u0_n146 ) , .ZN( u1_u13_u0_n97 ) );
  NAND2_X1 u1_u13_u1_U10 (.A1( u1_u13_u1_n131 ) , .ZN( u1_u13_u1_n147 ) , .A2( u1_u13_u1_n153 ) );
  NAND3_X1 u1_u13_u1_U100 (.ZN( u1_u13_u1_n113 ) , .A1( u1_u13_u1_n120 ) , .A3( u1_u13_u1_n133 ) , .A2( u1_u13_u1_n155 ) );
  AOI22_X1 u1_u13_u1_U11 (.B2( u1_u13_u1_n136 ) , .A2( u1_u13_u1_n137 ) , .ZN( u1_u13_u1_n143 ) , .A1( u1_u13_u1_n171 ) , .B1( u1_u13_u1_n173 ) );
  INV_X1 u1_u13_u1_U12 (.A( u1_u13_u1_n147 ) , .ZN( u1_u13_u1_n181 ) );
  INV_X1 u1_u13_u1_U13 (.A( u1_u13_u1_n139 ) , .ZN( u1_u13_u1_n174 ) );
  OR4_X1 u1_u13_u1_U14 (.A4( u1_u13_u1_n106 ) , .A3( u1_u13_u1_n107 ) , .ZN( u1_u13_u1_n108 ) , .A1( u1_u13_u1_n117 ) , .A2( u1_u13_u1_n184 ) );
  AOI21_X1 u1_u13_u1_U15 (.ZN( u1_u13_u1_n106 ) , .A( u1_u13_u1_n112 ) , .B1( u1_u13_u1_n154 ) , .B2( u1_u13_u1_n156 ) );
  AOI21_X1 u1_u13_u1_U16 (.ZN( u1_u13_u1_n107 ) , .B1( u1_u13_u1_n134 ) , .B2( u1_u13_u1_n149 ) , .A( u1_u13_u1_n174 ) );
  INV_X1 u1_u13_u1_U17 (.A( u1_u13_u1_n101 ) , .ZN( u1_u13_u1_n184 ) );
  INV_X1 u1_u13_u1_U18 (.A( u1_u13_u1_n112 ) , .ZN( u1_u13_u1_n171 ) );
  NAND2_X1 u1_u13_u1_U19 (.ZN( u1_u13_u1_n141 ) , .A1( u1_u13_u1_n153 ) , .A2( u1_u13_u1_n156 ) );
  AND2_X1 u1_u13_u1_U20 (.A1( u1_u13_u1_n123 ) , .ZN( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n161 ) );
  NAND2_X1 u1_u13_u1_U21 (.A2( u1_u13_u1_n115 ) , .A1( u1_u13_u1_n116 ) , .ZN( u1_u13_u1_n148 ) );
  NAND2_X1 u1_u13_u1_U22 (.A2( u1_u13_u1_n133 ) , .A1( u1_u13_u1_n135 ) , .ZN( u1_u13_u1_n159 ) );
  NAND2_X1 u1_u13_u1_U23 (.A2( u1_u13_u1_n115 ) , .A1( u1_u13_u1_n120 ) , .ZN( u1_u13_u1_n132 ) );
  INV_X1 u1_u13_u1_U24 (.A( u1_u13_u1_n154 ) , .ZN( u1_u13_u1_n178 ) );
  AOI22_X1 u1_u13_u1_U25 (.B2( u1_u13_u1_n113 ) , .A2( u1_u13_u1_n114 ) , .ZN( u1_u13_u1_n125 ) , .A1( u1_u13_u1_n171 ) , .B1( u1_u13_u1_n173 ) );
  NAND2_X1 u1_u13_u1_U26 (.ZN( u1_u13_u1_n114 ) , .A1( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n156 ) );
  INV_X1 u1_u13_u1_U27 (.A( u1_u13_u1_n151 ) , .ZN( u1_u13_u1_n183 ) );
  AND2_X1 u1_u13_u1_U28 (.A1( u1_u13_u1_n129 ) , .A2( u1_u13_u1_n133 ) , .ZN( u1_u13_u1_n149 ) );
  INV_X1 u1_u13_u1_U29 (.A( u1_u13_u1_n131 ) , .ZN( u1_u13_u1_n180 ) );
  INV_X1 u1_u13_u1_U3 (.A( u1_u13_u1_n159 ) , .ZN( u1_u13_u1_n182 ) );
  OAI221_X1 u1_u13_u1_U30 (.A( u1_u13_u1_n119 ) , .C2( u1_u13_u1_n129 ) , .ZN( u1_u13_u1_n138 ) , .B2( u1_u13_u1_n152 ) , .C1( u1_u13_u1_n174 ) , .B1( u1_u13_u1_n187 ) );
  INV_X1 u1_u13_u1_U31 (.A( u1_u13_u1_n148 ) , .ZN( u1_u13_u1_n187 ) );
  AOI211_X1 u1_u13_u1_U32 (.B( u1_u13_u1_n117 ) , .A( u1_u13_u1_n118 ) , .ZN( u1_u13_u1_n119 ) , .C2( u1_u13_u1_n146 ) , .C1( u1_u13_u1_n159 ) );
  NOR2_X1 u1_u13_u1_U33 (.A1( u1_u13_u1_n168 ) , .A2( u1_u13_u1_n176 ) , .ZN( u1_u13_u1_n98 ) );
  AOI211_X1 u1_u13_u1_U34 (.B( u1_u13_u1_n162 ) , .A( u1_u13_u1_n163 ) , .C2( u1_u13_u1_n164 ) , .ZN( u1_u13_u1_n165 ) , .C1( u1_u13_u1_n171 ) );
  AOI21_X1 u1_u13_u1_U35 (.A( u1_u13_u1_n160 ) , .B2( u1_u13_u1_n161 ) , .ZN( u1_u13_u1_n162 ) , .B1( u1_u13_u1_n182 ) );
  OR2_X1 u1_u13_u1_U36 (.A2( u1_u13_u1_n157 ) , .A1( u1_u13_u1_n158 ) , .ZN( u1_u13_u1_n163 ) );
  OAI21_X1 u1_u13_u1_U37 (.B2( u1_u13_u1_n123 ) , .ZN( u1_u13_u1_n145 ) , .B1( u1_u13_u1_n160 ) , .A( u1_u13_u1_n185 ) );
  INV_X1 u1_u13_u1_U38 (.A( u1_u13_u1_n122 ) , .ZN( u1_u13_u1_n185 ) );
  AOI21_X1 u1_u13_u1_U39 (.B2( u1_u13_u1_n120 ) , .B1( u1_u13_u1_n121 ) , .ZN( u1_u13_u1_n122 ) , .A( u1_u13_u1_n128 ) );
  AOI221_X1 u1_u13_u1_U4 (.A( u1_u13_u1_n138 ) , .C2( u1_u13_u1_n139 ) , .C1( u1_u13_u1_n140 ) , .B2( u1_u13_u1_n141 ) , .ZN( u1_u13_u1_n142 ) , .B1( u1_u13_u1_n175 ) );
  NAND2_X1 u1_u13_u1_U40 (.A1( u1_u13_u1_n128 ) , .ZN( u1_u13_u1_n146 ) , .A2( u1_u13_u1_n160 ) );
  NAND2_X1 u1_u13_u1_U41 (.A2( u1_u13_u1_n112 ) , .ZN( u1_u13_u1_n139 ) , .A1( u1_u13_u1_n152 ) );
  NAND2_X1 u1_u13_u1_U42 (.A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n156 ) , .A2( u1_u13_u1_n99 ) );
  AOI221_X1 u1_u13_u1_U43 (.B1( u1_u13_u1_n140 ) , .ZN( u1_u13_u1_n167 ) , .B2( u1_u13_u1_n172 ) , .C2( u1_u13_u1_n175 ) , .C1( u1_u13_u1_n178 ) , .A( u1_u13_u1_n188 ) );
  INV_X1 u1_u13_u1_U44 (.ZN( u1_u13_u1_n188 ) , .A( u1_u13_u1_n97 ) );
  AOI211_X1 u1_u13_u1_U45 (.A( u1_u13_u1_n118 ) , .C1( u1_u13_u1_n132 ) , .C2( u1_u13_u1_n139 ) , .B( u1_u13_u1_n96 ) , .ZN( u1_u13_u1_n97 ) );
  AOI21_X1 u1_u13_u1_U46 (.B2( u1_u13_u1_n121 ) , .B1( u1_u13_u1_n135 ) , .A( u1_u13_u1_n152 ) , .ZN( u1_u13_u1_n96 ) );
  NOR2_X1 u1_u13_u1_U47 (.ZN( u1_u13_u1_n117 ) , .A1( u1_u13_u1_n121 ) , .A2( u1_u13_u1_n160 ) );
  AOI21_X1 u1_u13_u1_U48 (.A( u1_u13_u1_n128 ) , .B2( u1_u13_u1_n129 ) , .ZN( u1_u13_u1_n130 ) , .B1( u1_u13_u1_n150 ) );
  NAND2_X1 u1_u13_u1_U49 (.ZN( u1_u13_u1_n112 ) , .A1( u1_u13_u1_n169 ) , .A2( u1_u13_u1_n170 ) );
  AOI211_X1 u1_u13_u1_U5 (.ZN( u1_u13_u1_n124 ) , .A( u1_u13_u1_n138 ) , .C2( u1_u13_u1_n139 ) , .B( u1_u13_u1_n145 ) , .C1( u1_u13_u1_n147 ) );
  NAND2_X1 u1_u13_u1_U50 (.ZN( u1_u13_u1_n129 ) , .A2( u1_u13_u1_n95 ) , .A1( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U51 (.A1( u1_u13_u1_n102 ) , .ZN( u1_u13_u1_n154 ) , .A2( u1_u13_u1_n99 ) );
  NAND2_X1 u1_u13_u1_U52 (.A2( u1_u13_u1_n100 ) , .ZN( u1_u13_u1_n135 ) , .A1( u1_u13_u1_n99 ) );
  AOI21_X1 u1_u13_u1_U53 (.A( u1_u13_u1_n152 ) , .B2( u1_u13_u1_n153 ) , .B1( u1_u13_u1_n154 ) , .ZN( u1_u13_u1_n158 ) );
  INV_X1 u1_u13_u1_U54 (.A( u1_u13_u1_n160 ) , .ZN( u1_u13_u1_n175 ) );
  NAND2_X1 u1_u13_u1_U55 (.A1( u1_u13_u1_n100 ) , .ZN( u1_u13_u1_n116 ) , .A2( u1_u13_u1_n95 ) );
  NAND2_X1 u1_u13_u1_U56 (.A1( u1_u13_u1_n102 ) , .ZN( u1_u13_u1_n131 ) , .A2( u1_u13_u1_n95 ) );
  NAND2_X1 u1_u13_u1_U57 (.A2( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n121 ) , .A1( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U58 (.A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n153 ) , .A2( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U59 (.A2( u1_u13_u1_n104 ) , .A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n133 ) );
  NOR2_X1 u1_u13_u1_U6 (.A1( u1_u13_u1_n112 ) , .A2( u1_u13_u1_n116 ) , .ZN( u1_u13_u1_n118 ) );
  NAND2_X1 u1_u13_u1_U60 (.ZN( u1_u13_u1_n150 ) , .A2( u1_u13_u1_n98 ) , .A1( u1_u13_u1_n99 ) );
  NAND2_X1 u1_u13_u1_U61 (.A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n155 ) , .A2( u1_u13_u1_n95 ) );
  OAI21_X1 u1_u13_u1_U62 (.ZN( u1_u13_u1_n109 ) , .B1( u1_u13_u1_n129 ) , .B2( u1_u13_u1_n160 ) , .A( u1_u13_u1_n167 ) );
  NAND2_X1 u1_u13_u1_U63 (.A2( u1_u13_u1_n100 ) , .A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n120 ) );
  NAND2_X1 u1_u13_u1_U64 (.A1( u1_u13_u1_n102 ) , .A2( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n115 ) );
  NAND2_X1 u1_u13_u1_U65 (.A2( u1_u13_u1_n100 ) , .A1( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n151 ) );
  NAND2_X1 u1_u13_u1_U66 (.A2( u1_u13_u1_n103 ) , .A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n161 ) );
  INV_X1 u1_u13_u1_U67 (.A( u1_u13_u1_n152 ) , .ZN( u1_u13_u1_n173 ) );
  INV_X1 u1_u13_u1_U68 (.A( u1_u13_u1_n128 ) , .ZN( u1_u13_u1_n172 ) );
  NAND2_X1 u1_u13_u1_U69 (.A2( u1_u13_u1_n102 ) , .A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n123 ) );
  OAI21_X1 u1_u13_u1_U7 (.ZN( u1_u13_u1_n101 ) , .B1( u1_u13_u1_n141 ) , .A( u1_u13_u1_n146 ) , .B2( u1_u13_u1_n183 ) );
  NOR2_X1 u1_u13_u1_U70 (.A2( u1_u13_X_7 ) , .A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n95 ) );
  NOR2_X1 u1_u13_u1_U71 (.A1( u1_u13_X_12 ) , .A2( u1_u13_X_9 ) , .ZN( u1_u13_u1_n100 ) );
  NOR2_X1 u1_u13_u1_U72 (.A2( u1_u13_X_8 ) , .A1( u1_u13_u1_n177 ) , .ZN( u1_u13_u1_n99 ) );
  NOR2_X1 u1_u13_u1_U73 (.A2( u1_u13_X_12 ) , .ZN( u1_u13_u1_n102 ) , .A1( u1_u13_u1_n176 ) );
  NOR2_X1 u1_u13_u1_U74 (.A2( u1_u13_X_9 ) , .ZN( u1_u13_u1_n105 ) , .A1( u1_u13_u1_n168 ) );
  NAND2_X1 u1_u13_u1_U75 (.A1( u1_u13_X_10 ) , .ZN( u1_u13_u1_n160 ) , .A2( u1_u13_u1_n169 ) );
  NAND2_X1 u1_u13_u1_U76 (.A2( u1_u13_X_10 ) , .A1( u1_u13_X_11 ) , .ZN( u1_u13_u1_n152 ) );
  NAND2_X1 u1_u13_u1_U77 (.A1( u1_u13_X_11 ) , .ZN( u1_u13_u1_n128 ) , .A2( u1_u13_u1_n170 ) );
  AND2_X1 u1_u13_u1_U78 (.A2( u1_u13_X_7 ) , .A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n104 ) );
  AND2_X1 u1_u13_u1_U79 (.A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n103 ) , .A2( u1_u13_u1_n177 ) );
  AOI21_X1 u1_u13_u1_U8 (.B2( u1_u13_u1_n155 ) , .B1( u1_u13_u1_n156 ) , .ZN( u1_u13_u1_n157 ) , .A( u1_u13_u1_n174 ) );
  INV_X1 u1_u13_u1_U80 (.A( u1_u13_X_10 ) , .ZN( u1_u13_u1_n170 ) );
  INV_X1 u1_u13_u1_U81 (.A( u1_u13_X_9 ) , .ZN( u1_u13_u1_n176 ) );
  INV_X1 u1_u13_u1_U82 (.A( u1_u13_X_11 ) , .ZN( u1_u13_u1_n169 ) );
  INV_X1 u1_u13_u1_U83 (.A( u1_u13_X_12 ) , .ZN( u1_u13_u1_n168 ) );
  INV_X1 u1_u13_u1_U84 (.A( u1_u13_X_7 ) , .ZN( u1_u13_u1_n177 ) );
  NAND4_X1 u1_u13_u1_U85 (.ZN( u1_out13_18 ) , .A4( u1_u13_u1_n165 ) , .A3( u1_u13_u1_n166 ) , .A1( u1_u13_u1_n167 ) , .A2( u1_u13_u1_n186 ) );
  AOI22_X1 u1_u13_u1_U86 (.B2( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n147 ) , .A2( u1_u13_u1_n148 ) , .ZN( u1_u13_u1_n166 ) , .A1( u1_u13_u1_n172 ) );
  INV_X1 u1_u13_u1_U87 (.A( u1_u13_u1_n145 ) , .ZN( u1_u13_u1_n186 ) );
  NAND4_X1 u1_u13_u1_U88 (.ZN( u1_out13_2 ) , .A4( u1_u13_u1_n142 ) , .A3( u1_u13_u1_n143 ) , .A2( u1_u13_u1_n144 ) , .A1( u1_u13_u1_n179 ) );
  OAI21_X1 u1_u13_u1_U89 (.B2( u1_u13_u1_n132 ) , .ZN( u1_u13_u1_n144 ) , .A( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n180 ) );
  NAND2_X1 u1_u13_u1_U9 (.ZN( u1_u13_u1_n140 ) , .A2( u1_u13_u1_n150 ) , .A1( u1_u13_u1_n155 ) );
  INV_X1 u1_u13_u1_U90 (.A( u1_u13_u1_n130 ) , .ZN( u1_u13_u1_n179 ) );
  NAND4_X1 u1_u13_u1_U91 (.ZN( u1_out13_28 ) , .A4( u1_u13_u1_n124 ) , .A3( u1_u13_u1_n125 ) , .A2( u1_u13_u1_n126 ) , .A1( u1_u13_u1_n127 ) );
  OAI21_X1 u1_u13_u1_U92 (.ZN( u1_u13_u1_n127 ) , .B2( u1_u13_u1_n139 ) , .B1( u1_u13_u1_n175 ) , .A( u1_u13_u1_n183 ) );
  OAI21_X1 u1_u13_u1_U93 (.ZN( u1_u13_u1_n126 ) , .B2( u1_u13_u1_n140 ) , .A( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n178 ) );
  OR4_X1 u1_u13_u1_U94 (.ZN( u1_out13_13 ) , .A4( u1_u13_u1_n108 ) , .A3( u1_u13_u1_n109 ) , .A2( u1_u13_u1_n110 ) , .A1( u1_u13_u1_n111 ) );
  AOI21_X1 u1_u13_u1_U95 (.ZN( u1_u13_u1_n111 ) , .A( u1_u13_u1_n128 ) , .B2( u1_u13_u1_n131 ) , .B1( u1_u13_u1_n135 ) );
  AOI21_X1 u1_u13_u1_U96 (.ZN( u1_u13_u1_n110 ) , .A( u1_u13_u1_n116 ) , .B1( u1_u13_u1_n152 ) , .B2( u1_u13_u1_n160 ) );
  NAND3_X1 u1_u13_u1_U97 (.A3( u1_u13_u1_n149 ) , .A2( u1_u13_u1_n150 ) , .A1( u1_u13_u1_n151 ) , .ZN( u1_u13_u1_n164 ) );
  NAND3_X1 u1_u13_u1_U98 (.A3( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n135 ) , .ZN( u1_u13_u1_n136 ) , .A1( u1_u13_u1_n151 ) );
  NAND3_X1 u1_u13_u1_U99 (.A1( u1_u13_u1_n133 ) , .ZN( u1_u13_u1_n137 ) , .A2( u1_u13_u1_n154 ) , .A3( u1_u13_u1_n181 ) );
  OAI22_X1 u1_u13_u2_U10 (.B1( u1_u13_u2_n151 ) , .A2( u1_u13_u2_n152 ) , .A1( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n160 ) , .B2( u1_u13_u2_n168 ) );
  NAND3_X1 u1_u13_u2_U100 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n104 ) , .A3( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n98 ) );
  NOR3_X1 u1_u13_u2_U11 (.A1( u1_u13_u2_n150 ) , .ZN( u1_u13_u2_n151 ) , .A3( u1_u13_u2_n175 ) , .A2( u1_u13_u2_n188 ) );
  AOI21_X1 u1_u13_u2_U12 (.B2( u1_u13_u2_n123 ) , .ZN( u1_u13_u2_n125 ) , .A( u1_u13_u2_n171 ) , .B1( u1_u13_u2_n184 ) );
  INV_X1 u1_u13_u2_U13 (.A( u1_u13_u2_n150 ) , .ZN( u1_u13_u2_n184 ) );
  AOI21_X1 u1_u13_u2_U14 (.ZN( u1_u13_u2_n144 ) , .B2( u1_u13_u2_n155 ) , .A( u1_u13_u2_n172 ) , .B1( u1_u13_u2_n185 ) );
  AOI21_X1 u1_u13_u2_U15 (.B2( u1_u13_u2_n143 ) , .ZN( u1_u13_u2_n145 ) , .B1( u1_u13_u2_n152 ) , .A( u1_u13_u2_n171 ) );
  INV_X1 u1_u13_u2_U16 (.A( u1_u13_u2_n156 ) , .ZN( u1_u13_u2_n171 ) );
  INV_X1 u1_u13_u2_U17 (.A( u1_u13_u2_n120 ) , .ZN( u1_u13_u2_n188 ) );
  NAND2_X1 u1_u13_u2_U18 (.A2( u1_u13_u2_n122 ) , .ZN( u1_u13_u2_n150 ) , .A1( u1_u13_u2_n152 ) );
  INV_X1 u1_u13_u2_U19 (.A( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n170 ) );
  INV_X1 u1_u13_u2_U20 (.A( u1_u13_u2_n137 ) , .ZN( u1_u13_u2_n173 ) );
  NAND2_X1 u1_u13_u2_U21 (.A1( u1_u13_u2_n132 ) , .A2( u1_u13_u2_n139 ) , .ZN( u1_u13_u2_n157 ) );
  INV_X1 u1_u13_u2_U22 (.A( u1_u13_u2_n113 ) , .ZN( u1_u13_u2_n178 ) );
  INV_X1 u1_u13_u2_U23 (.A( u1_u13_u2_n139 ) , .ZN( u1_u13_u2_n175 ) );
  INV_X1 u1_u13_u2_U24 (.A( u1_u13_u2_n155 ) , .ZN( u1_u13_u2_n181 ) );
  INV_X1 u1_u13_u2_U25 (.A( u1_u13_u2_n119 ) , .ZN( u1_u13_u2_n177 ) );
  INV_X1 u1_u13_u2_U26 (.A( u1_u13_u2_n116 ) , .ZN( u1_u13_u2_n180 ) );
  INV_X1 u1_u13_u2_U27 (.A( u1_u13_u2_n131 ) , .ZN( u1_u13_u2_n179 ) );
  INV_X1 u1_u13_u2_U28 (.A( u1_u13_u2_n154 ) , .ZN( u1_u13_u2_n176 ) );
  NAND2_X1 u1_u13_u2_U29 (.A2( u1_u13_u2_n116 ) , .A1( u1_u13_u2_n117 ) , .ZN( u1_u13_u2_n118 ) );
  NOR2_X1 u1_u13_u2_U3 (.ZN( u1_u13_u2_n121 ) , .A2( u1_u13_u2_n177 ) , .A1( u1_u13_u2_n180 ) );
  INV_X1 u1_u13_u2_U30 (.A( u1_u13_u2_n132 ) , .ZN( u1_u13_u2_n182 ) );
  INV_X1 u1_u13_u2_U31 (.A( u1_u13_u2_n158 ) , .ZN( u1_u13_u2_n183 ) );
  OAI21_X1 u1_u13_u2_U32 (.A( u1_u13_u2_n156 ) , .B1( u1_u13_u2_n157 ) , .ZN( u1_u13_u2_n158 ) , .B2( u1_u13_u2_n179 ) );
  NOR2_X1 u1_u13_u2_U33 (.ZN( u1_u13_u2_n156 ) , .A1( u1_u13_u2_n166 ) , .A2( u1_u13_u2_n169 ) );
  NOR2_X1 u1_u13_u2_U34 (.A2( u1_u13_u2_n114 ) , .ZN( u1_u13_u2_n137 ) , .A1( u1_u13_u2_n140 ) );
  NOR2_X1 u1_u13_u2_U35 (.A2( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n153 ) , .A1( u1_u13_u2_n156 ) );
  AOI211_X1 u1_u13_u2_U36 (.ZN( u1_u13_u2_n130 ) , .C1( u1_u13_u2_n138 ) , .C2( u1_u13_u2_n179 ) , .B( u1_u13_u2_n96 ) , .A( u1_u13_u2_n97 ) );
  OAI22_X1 u1_u13_u2_U37 (.B1( u1_u13_u2_n133 ) , .A2( u1_u13_u2_n137 ) , .A1( u1_u13_u2_n152 ) , .B2( u1_u13_u2_n168 ) , .ZN( u1_u13_u2_n97 ) );
  OAI221_X1 u1_u13_u2_U38 (.B1( u1_u13_u2_n113 ) , .C1( u1_u13_u2_n132 ) , .A( u1_u13_u2_n149 ) , .B2( u1_u13_u2_n171 ) , .C2( u1_u13_u2_n172 ) , .ZN( u1_u13_u2_n96 ) );
  OAI221_X1 u1_u13_u2_U39 (.A( u1_u13_u2_n115 ) , .C2( u1_u13_u2_n123 ) , .B2( u1_u13_u2_n143 ) , .B1( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n163 ) , .C1( u1_u13_u2_n168 ) );
  INV_X1 u1_u13_u2_U4 (.A( u1_u13_u2_n134 ) , .ZN( u1_u13_u2_n185 ) );
  OAI21_X1 u1_u13_u2_U40 (.A( u1_u13_u2_n114 ) , .ZN( u1_u13_u2_n115 ) , .B1( u1_u13_u2_n176 ) , .B2( u1_u13_u2_n178 ) );
  OAI221_X1 u1_u13_u2_U41 (.A( u1_u13_u2_n135 ) , .B2( u1_u13_u2_n136 ) , .B1( u1_u13_u2_n137 ) , .ZN( u1_u13_u2_n162 ) , .C2( u1_u13_u2_n167 ) , .C1( u1_u13_u2_n185 ) );
  AND3_X1 u1_u13_u2_U42 (.A3( u1_u13_u2_n131 ) , .A2( u1_u13_u2_n132 ) , .A1( u1_u13_u2_n133 ) , .ZN( u1_u13_u2_n136 ) );
  AOI22_X1 u1_u13_u2_U43 (.ZN( u1_u13_u2_n135 ) , .B1( u1_u13_u2_n140 ) , .A1( u1_u13_u2_n156 ) , .B2( u1_u13_u2_n180 ) , .A2( u1_u13_u2_n188 ) );
  AOI21_X1 u1_u13_u2_U44 (.ZN( u1_u13_u2_n149 ) , .B1( u1_u13_u2_n173 ) , .B2( u1_u13_u2_n188 ) , .A( u1_u13_u2_n95 ) );
  AND3_X1 u1_u13_u2_U45 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n104 ) , .A3( u1_u13_u2_n156 ) , .ZN( u1_u13_u2_n95 ) );
  OAI21_X1 u1_u13_u2_U46 (.A( u1_u13_u2_n101 ) , .B2( u1_u13_u2_n121 ) , .B1( u1_u13_u2_n153 ) , .ZN( u1_u13_u2_n164 ) );
  NAND2_X1 u1_u13_u2_U47 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n107 ) , .ZN( u1_u13_u2_n155 ) );
  NAND2_X1 u1_u13_u2_U48 (.A2( u1_u13_u2_n105 ) , .A1( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n143 ) );
  NAND2_X1 u1_u13_u2_U49 (.A1( u1_u13_u2_n104 ) , .A2( u1_u13_u2_n106 ) , .ZN( u1_u13_u2_n152 ) );
  NOR4_X1 u1_u13_u2_U5 (.A4( u1_u13_u2_n124 ) , .A3( u1_u13_u2_n125 ) , .A2( u1_u13_u2_n126 ) , .A1( u1_u13_u2_n127 ) , .ZN( u1_u13_u2_n128 ) );
  NAND2_X1 u1_u13_u2_U50 (.A1( u1_u13_u2_n100 ) , .A2( u1_u13_u2_n105 ) , .ZN( u1_u13_u2_n132 ) );
  INV_X1 u1_u13_u2_U51 (.A( u1_u13_u2_n140 ) , .ZN( u1_u13_u2_n168 ) );
  INV_X1 u1_u13_u2_U52 (.A( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n167 ) );
  OAI21_X1 u1_u13_u2_U53 (.A( u1_u13_u2_n141 ) , .B2( u1_u13_u2_n142 ) , .ZN( u1_u13_u2_n146 ) , .B1( u1_u13_u2_n153 ) );
  OAI21_X1 u1_u13_u2_U54 (.A( u1_u13_u2_n140 ) , .ZN( u1_u13_u2_n141 ) , .B1( u1_u13_u2_n176 ) , .B2( u1_u13_u2_n177 ) );
  NOR3_X1 u1_u13_u2_U55 (.ZN( u1_u13_u2_n142 ) , .A3( u1_u13_u2_n175 ) , .A2( u1_u13_u2_n178 ) , .A1( u1_u13_u2_n181 ) );
  NAND2_X1 u1_u13_u2_U56 (.A1( u1_u13_u2_n102 ) , .A2( u1_u13_u2_n106 ) , .ZN( u1_u13_u2_n113 ) );
  NAND2_X1 u1_u13_u2_U57 (.A1( u1_u13_u2_n106 ) , .A2( u1_u13_u2_n107 ) , .ZN( u1_u13_u2_n131 ) );
  NAND2_X1 u1_u13_u2_U58 (.A1( u1_u13_u2_n103 ) , .A2( u1_u13_u2_n107 ) , .ZN( u1_u13_u2_n139 ) );
  NAND2_X1 u1_u13_u2_U59 (.A1( u1_u13_u2_n103 ) , .A2( u1_u13_u2_n105 ) , .ZN( u1_u13_u2_n133 ) );
  AOI21_X1 u1_u13_u2_U6 (.B2( u1_u13_u2_n119 ) , .ZN( u1_u13_u2_n127 ) , .A( u1_u13_u2_n137 ) , .B1( u1_u13_u2_n155 ) );
  NAND2_X1 u1_u13_u2_U60 (.A1( u1_u13_u2_n102 ) , .A2( u1_u13_u2_n103 ) , .ZN( u1_u13_u2_n154 ) );
  NAND2_X1 u1_u13_u2_U61 (.A2( u1_u13_u2_n103 ) , .A1( u1_u13_u2_n104 ) , .ZN( u1_u13_u2_n119 ) );
  NAND2_X1 u1_u13_u2_U62 (.A2( u1_u13_u2_n107 ) , .A1( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n123 ) );
  NAND2_X1 u1_u13_u2_U63 (.A1( u1_u13_u2_n104 ) , .A2( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n122 ) );
  INV_X1 u1_u13_u2_U64 (.A( u1_u13_u2_n114 ) , .ZN( u1_u13_u2_n172 ) );
  NAND2_X1 u1_u13_u2_U65 (.A2( u1_u13_u2_n100 ) , .A1( u1_u13_u2_n102 ) , .ZN( u1_u13_u2_n116 ) );
  NAND2_X1 u1_u13_u2_U66 (.A1( u1_u13_u2_n102 ) , .A2( u1_u13_u2_n108 ) , .ZN( u1_u13_u2_n120 ) );
  NAND2_X1 u1_u13_u2_U67 (.A2( u1_u13_u2_n105 ) , .A1( u1_u13_u2_n106 ) , .ZN( u1_u13_u2_n117 ) );
  INV_X1 u1_u13_u2_U68 (.ZN( u1_u13_u2_n187 ) , .A( u1_u13_u2_n99 ) );
  OAI21_X1 u1_u13_u2_U69 (.B1( u1_u13_u2_n137 ) , .B2( u1_u13_u2_n143 ) , .A( u1_u13_u2_n98 ) , .ZN( u1_u13_u2_n99 ) );
  AOI21_X1 u1_u13_u2_U7 (.ZN( u1_u13_u2_n124 ) , .B1( u1_u13_u2_n131 ) , .B2( u1_u13_u2_n143 ) , .A( u1_u13_u2_n172 ) );
  NOR2_X1 u1_u13_u2_U70 (.A2( u1_u13_X_16 ) , .ZN( u1_u13_u2_n140 ) , .A1( u1_u13_u2_n166 ) );
  NOR2_X1 u1_u13_u2_U71 (.A2( u1_u13_X_13 ) , .A1( u1_u13_X_14 ) , .ZN( u1_u13_u2_n100 ) );
  NOR2_X1 u1_u13_u2_U72 (.A2( u1_u13_X_16 ) , .A1( u1_u13_X_17 ) , .ZN( u1_u13_u2_n138 ) );
  NOR2_X1 u1_u13_u2_U73 (.A2( u1_u13_X_15 ) , .A1( u1_u13_X_18 ) , .ZN( u1_u13_u2_n104 ) );
  NOR2_X1 u1_u13_u2_U74 (.A2( u1_u13_X_14 ) , .ZN( u1_u13_u2_n103 ) , .A1( u1_u13_u2_n174 ) );
  NOR2_X1 u1_u13_u2_U75 (.A2( u1_u13_X_15 ) , .ZN( u1_u13_u2_n102 ) , .A1( u1_u13_u2_n165 ) );
  NOR2_X1 u1_u13_u2_U76 (.A2( u1_u13_X_17 ) , .ZN( u1_u13_u2_n114 ) , .A1( u1_u13_u2_n169 ) );
  AND2_X1 u1_u13_u2_U77 (.A1( u1_u13_X_15 ) , .ZN( u1_u13_u2_n105 ) , .A2( u1_u13_u2_n165 ) );
  AND2_X1 u1_u13_u2_U78 (.A2( u1_u13_X_15 ) , .A1( u1_u13_X_18 ) , .ZN( u1_u13_u2_n107 ) );
  AND2_X1 u1_u13_u2_U79 (.A1( u1_u13_X_14 ) , .ZN( u1_u13_u2_n106 ) , .A2( u1_u13_u2_n174 ) );
  AOI21_X1 u1_u13_u2_U8 (.B2( u1_u13_u2_n120 ) , .B1( u1_u13_u2_n121 ) , .ZN( u1_u13_u2_n126 ) , .A( u1_u13_u2_n167 ) );
  AND2_X1 u1_u13_u2_U80 (.A1( u1_u13_X_13 ) , .A2( u1_u13_X_14 ) , .ZN( u1_u13_u2_n108 ) );
  INV_X1 u1_u13_u2_U81 (.A( u1_u13_X_16 ) , .ZN( u1_u13_u2_n169 ) );
  INV_X1 u1_u13_u2_U82 (.A( u1_u13_X_17 ) , .ZN( u1_u13_u2_n166 ) );
  INV_X1 u1_u13_u2_U83 (.A( u1_u13_X_13 ) , .ZN( u1_u13_u2_n174 ) );
  INV_X1 u1_u13_u2_U84 (.A( u1_u13_X_18 ) , .ZN( u1_u13_u2_n165 ) );
  NAND4_X1 u1_u13_u2_U85 (.ZN( u1_out13_30 ) , .A4( u1_u13_u2_n147 ) , .A3( u1_u13_u2_n148 ) , .A2( u1_u13_u2_n149 ) , .A1( u1_u13_u2_n187 ) );
  NOR3_X1 u1_u13_u2_U86 (.A3( u1_u13_u2_n144 ) , .A2( u1_u13_u2_n145 ) , .A1( u1_u13_u2_n146 ) , .ZN( u1_u13_u2_n147 ) );
  AOI21_X1 u1_u13_u2_U87 (.B2( u1_u13_u2_n138 ) , .ZN( u1_u13_u2_n148 ) , .A( u1_u13_u2_n162 ) , .B1( u1_u13_u2_n182 ) );
  NAND4_X1 u1_u13_u2_U88 (.ZN( u1_out13_24 ) , .A4( u1_u13_u2_n111 ) , .A3( u1_u13_u2_n112 ) , .A1( u1_u13_u2_n130 ) , .A2( u1_u13_u2_n187 ) );
  AOI221_X1 u1_u13_u2_U89 (.A( u1_u13_u2_n109 ) , .B1( u1_u13_u2_n110 ) , .ZN( u1_u13_u2_n111 ) , .C1( u1_u13_u2_n134 ) , .C2( u1_u13_u2_n170 ) , .B2( u1_u13_u2_n173 ) );
  OAI22_X1 u1_u13_u2_U9 (.ZN( u1_u13_u2_n109 ) , .A2( u1_u13_u2_n113 ) , .B2( u1_u13_u2_n133 ) , .B1( u1_u13_u2_n167 ) , .A1( u1_u13_u2_n168 ) );
  AOI21_X1 u1_u13_u2_U90 (.ZN( u1_u13_u2_n112 ) , .B2( u1_u13_u2_n156 ) , .A( u1_u13_u2_n164 ) , .B1( u1_u13_u2_n181 ) );
  NAND4_X1 u1_u13_u2_U91 (.ZN( u1_out13_16 ) , .A4( u1_u13_u2_n128 ) , .A3( u1_u13_u2_n129 ) , .A1( u1_u13_u2_n130 ) , .A2( u1_u13_u2_n186 ) );
  AOI22_X1 u1_u13_u2_U92 (.A2( u1_u13_u2_n118 ) , .ZN( u1_u13_u2_n129 ) , .A1( u1_u13_u2_n140 ) , .B1( u1_u13_u2_n157 ) , .B2( u1_u13_u2_n170 ) );
  INV_X1 u1_u13_u2_U93 (.A( u1_u13_u2_n163 ) , .ZN( u1_u13_u2_n186 ) );
  OR4_X1 u1_u13_u2_U94 (.ZN( u1_out13_6 ) , .A4( u1_u13_u2_n161 ) , .A3( u1_u13_u2_n162 ) , .A2( u1_u13_u2_n163 ) , .A1( u1_u13_u2_n164 ) );
  OR3_X1 u1_u13_u2_U95 (.A2( u1_u13_u2_n159 ) , .A1( u1_u13_u2_n160 ) , .ZN( u1_u13_u2_n161 ) , .A3( u1_u13_u2_n183 ) );
  AOI21_X1 u1_u13_u2_U96 (.B2( u1_u13_u2_n154 ) , .B1( u1_u13_u2_n155 ) , .ZN( u1_u13_u2_n159 ) , .A( u1_u13_u2_n167 ) );
  NAND3_X1 u1_u13_u2_U97 (.A2( u1_u13_u2_n117 ) , .A1( u1_u13_u2_n122 ) , .A3( u1_u13_u2_n123 ) , .ZN( u1_u13_u2_n134 ) );
  NAND3_X1 u1_u13_u2_U98 (.ZN( u1_u13_u2_n110 ) , .A2( u1_u13_u2_n131 ) , .A3( u1_u13_u2_n139 ) , .A1( u1_u13_u2_n154 ) );
  NAND3_X1 u1_u13_u2_U99 (.A2( u1_u13_u2_n100 ) , .ZN( u1_u13_u2_n101 ) , .A1( u1_u13_u2_n104 ) , .A3( u1_u13_u2_n114 ) );
  XOR2_X1 u1_u15_U1 (.A( u1_FP_38 ) , .B( u1_K16_9 ) , .Z( u1_u15_X_9 ) );
  XOR2_X1 u1_u15_U16 (.A( u1_FP_34 ) , .B( u1_K16_3 ) , .Z( u1_u15_X_3 ) );
  XOR2_X1 u1_u15_U2 (.A( u1_FP_37 ) , .B( u1_K16_8 ) , .Z( u1_u15_X_8 ) );
  XOR2_X1 u1_u15_U27 (.A( u1_FP_33 ) , .B( u1_K16_2 ) , .Z( u1_u15_X_2 ) );
  XOR2_X1 u1_u15_U3 (.A( u1_FP_36 ) , .B( u1_K16_7 ) , .Z( u1_u15_X_7 ) );
  XOR2_X1 u1_u15_U33 (.A( u1_FP_49 ) , .B( u1_K16_24 ) , .Z( u1_u15_X_24 ) );
  XOR2_X1 u1_u15_U34 (.A( u1_FP_48 ) , .B( u1_K16_23 ) , .Z( u1_u15_X_23 ) );
  XOR2_X1 u1_u15_U35 (.A( u1_FP_47 ) , .B( u1_K16_22 ) , .Z( u1_u15_X_22 ) );
  XOR2_X1 u1_u15_U36 (.A( u1_FP_46 ) , .B( u1_K16_21 ) , .Z( u1_u15_X_21 ) );
  XOR2_X1 u1_u15_U37 (.A( u1_FP_45 ) , .B( u1_K16_20 ) , .Z( u1_u15_X_20 ) );
  XOR2_X1 u1_u15_U38 (.A( u1_FP_64 ) , .B( u1_K16_1 ) , .Z( u1_u15_X_1 ) );
  XOR2_X1 u1_u15_U39 (.A( u1_FP_44 ) , .B( u1_K16_19 ) , .Z( u1_u15_X_19 ) );
  XOR2_X1 u1_u15_U4 (.A( u1_FP_37 ) , .B( u1_K16_6 ) , .Z( u1_u15_X_6 ) );
  XOR2_X1 u1_u15_U46 (.A( u1_FP_41 ) , .B( u1_K16_12 ) , .Z( u1_u15_X_12 ) );
  XOR2_X1 u1_u15_U47 (.A( u1_FP_40 ) , .B( u1_K16_11 ) , .Z( u1_u15_X_11 ) );
  XOR2_X1 u1_u15_U48 (.A( u1_FP_39 ) , .B( u1_K16_10 ) , .Z( u1_u15_X_10 ) );
  XOR2_X1 u1_u15_U5 (.A( u1_FP_36 ) , .B( u1_K16_5 ) , .Z( u1_u15_X_5 ) );
  XOR2_X1 u1_u15_U6 (.A( u1_FP_35 ) , .B( u1_K16_4 ) , .Z( u1_u15_X_4 ) );
  AND3_X1 u1_u15_u0_U10 (.A2( u1_u15_u0_n112 ) , .ZN( u1_u15_u0_n127 ) , .A3( u1_u15_u0_n130 ) , .A1( u1_u15_u0_n148 ) );
  NAND2_X1 u1_u15_u0_U11 (.ZN( u1_u15_u0_n113 ) , .A1( u1_u15_u0_n139 ) , .A2( u1_u15_u0_n149 ) );
  AND2_X1 u1_u15_u0_U12 (.ZN( u1_u15_u0_n107 ) , .A1( u1_u15_u0_n130 ) , .A2( u1_u15_u0_n140 ) );
  AND2_X1 u1_u15_u0_U13 (.A2( u1_u15_u0_n129 ) , .A1( u1_u15_u0_n130 ) , .ZN( u1_u15_u0_n151 ) );
  AND2_X1 u1_u15_u0_U14 (.A1( u1_u15_u0_n108 ) , .A2( u1_u15_u0_n125 ) , .ZN( u1_u15_u0_n145 ) );
  INV_X1 u1_u15_u0_U15 (.A( u1_u15_u0_n143 ) , .ZN( u1_u15_u0_n173 ) );
  NOR2_X1 u1_u15_u0_U16 (.A2( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n147 ) , .A1( u1_u15_u0_n160 ) );
  AOI21_X1 u1_u15_u0_U17 (.B1( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n132 ) , .A( u1_u15_u0_n165 ) , .B2( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U18 (.A( u1_u15_u0_n142 ) , .ZN( u1_u15_u0_n165 ) );
  OAI221_X1 u1_u15_u0_U19 (.C1( u1_u15_u0_n121 ) , .ZN( u1_u15_u0_n122 ) , .B2( u1_u15_u0_n127 ) , .A( u1_u15_u0_n143 ) , .B1( u1_u15_u0_n144 ) , .C2( u1_u15_u0_n147 ) );
  OAI22_X1 u1_u15_u0_U20 (.B1( u1_u15_u0_n131 ) , .A1( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n147 ) , .A2( u1_u15_u0_n90 ) , .ZN( u1_u15_u0_n91 ) );
  AND3_X1 u1_u15_u0_U21 (.A3( u1_u15_u0_n121 ) , .A2( u1_u15_u0_n125 ) , .A1( u1_u15_u0_n148 ) , .ZN( u1_u15_u0_n90 ) );
  OAI22_X1 u1_u15_u0_U22 (.B1( u1_u15_u0_n125 ) , .ZN( u1_u15_u0_n126 ) , .A1( u1_u15_u0_n138 ) , .A2( u1_u15_u0_n146 ) , .B2( u1_u15_u0_n147 ) );
  NOR2_X1 u1_u15_u0_U23 (.A1( u1_u15_u0_n163 ) , .A2( u1_u15_u0_n164 ) , .ZN( u1_u15_u0_n95 ) );
  INV_X1 u1_u15_u0_U24 (.A( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n161 ) );
  NOR2_X1 u1_u15_u0_U25 (.A1( u1_u15_u0_n120 ) , .ZN( u1_u15_u0_n143 ) , .A2( u1_u15_u0_n167 ) );
  OAI221_X1 u1_u15_u0_U26 (.C1( u1_u15_u0_n112 ) , .ZN( u1_u15_u0_n120 ) , .B1( u1_u15_u0_n138 ) , .B2( u1_u15_u0_n141 ) , .C2( u1_u15_u0_n147 ) , .A( u1_u15_u0_n172 ) );
  AOI211_X1 u1_u15_u0_U27 (.B( u1_u15_u0_n115 ) , .A( u1_u15_u0_n116 ) , .C2( u1_u15_u0_n117 ) , .C1( u1_u15_u0_n118 ) , .ZN( u1_u15_u0_n119 ) );
  AOI22_X1 u1_u15_u0_U28 (.B2( u1_u15_u0_n109 ) , .A2( u1_u15_u0_n110 ) , .ZN( u1_u15_u0_n111 ) , .B1( u1_u15_u0_n118 ) , .A1( u1_u15_u0_n160 ) );
  NAND2_X1 u1_u15_u0_U29 (.A2( u1_u15_u0_n102 ) , .A1( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n149 ) );
  INV_X1 u1_u15_u0_U3 (.A( u1_u15_u0_n113 ) , .ZN( u1_u15_u0_n166 ) );
  INV_X1 u1_u15_u0_U30 (.A( u1_u15_u0_n118 ) , .ZN( u1_u15_u0_n158 ) );
  NAND2_X1 u1_u15_u0_U31 (.A2( u1_u15_u0_n100 ) , .ZN( u1_u15_u0_n131 ) , .A1( u1_u15_u0_n92 ) );
  NAND2_X1 u1_u15_u0_U32 (.ZN( u1_u15_u0_n108 ) , .A1( u1_u15_u0_n92 ) , .A2( u1_u15_u0_n94 ) );
  AOI21_X1 u1_u15_u0_U33 (.ZN( u1_u15_u0_n104 ) , .B1( u1_u15_u0_n107 ) , .B2( u1_u15_u0_n141 ) , .A( u1_u15_u0_n144 ) );
  AOI21_X1 u1_u15_u0_U34 (.B1( u1_u15_u0_n127 ) , .B2( u1_u15_u0_n129 ) , .A( u1_u15_u0_n138 ) , .ZN( u1_u15_u0_n96 ) );
  NAND2_X1 u1_u15_u0_U35 (.A2( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n114 ) , .A1( u1_u15_u0_n92 ) );
  AOI21_X1 u1_u15_u0_U36 (.ZN( u1_u15_u0_n116 ) , .B2( u1_u15_u0_n142 ) , .A( u1_u15_u0_n144 ) , .B1( u1_u15_u0_n166 ) );
  NAND2_X1 u1_u15_u0_U37 (.A2( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n140 ) , .A1( u1_u15_u0_n94 ) );
  NAND2_X1 u1_u15_u0_U38 (.A1( u1_u15_u0_n100 ) , .A2( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n125 ) );
  NAND2_X1 u1_u15_u0_U39 (.A1( u1_u15_u0_n101 ) , .A2( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n150 ) );
  AOI21_X1 u1_u15_u0_U4 (.B1( u1_u15_u0_n114 ) , .ZN( u1_u15_u0_n115 ) , .B2( u1_u15_u0_n129 ) , .A( u1_u15_u0_n161 ) );
  INV_X1 u1_u15_u0_U40 (.A( u1_u15_u0_n138 ) , .ZN( u1_u15_u0_n160 ) );
  NAND2_X1 u1_u15_u0_U41 (.A2( u1_u15_u0_n100 ) , .A1( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n139 ) );
  NAND2_X1 u1_u15_u0_U42 (.ZN( u1_u15_u0_n112 ) , .A2( u1_u15_u0_n92 ) , .A1( u1_u15_u0_n93 ) );
  NAND2_X1 u1_u15_u0_U43 (.A1( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n130 ) , .A2( u1_u15_u0_n94 ) );
  NAND2_X1 u1_u15_u0_U44 (.A2( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n121 ) , .A1( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U45 (.ZN( u1_u15_u0_n172 ) , .A( u1_u15_u0_n88 ) );
  OAI222_X1 u1_u15_u0_U46 (.C1( u1_u15_u0_n108 ) , .A1( u1_u15_u0_n125 ) , .B2( u1_u15_u0_n128 ) , .B1( u1_u15_u0_n144 ) , .A2( u1_u15_u0_n158 ) , .C2( u1_u15_u0_n161 ) , .ZN( u1_u15_u0_n88 ) );
  OR3_X1 u1_u15_u0_U47 (.A3( u1_u15_u0_n152 ) , .A2( u1_u15_u0_n153 ) , .A1( u1_u15_u0_n154 ) , .ZN( u1_u15_u0_n155 ) );
  AOI21_X1 u1_u15_u0_U48 (.B2( u1_u15_u0_n150 ) , .B1( u1_u15_u0_n151 ) , .ZN( u1_u15_u0_n152 ) , .A( u1_u15_u0_n158 ) );
  AOI21_X1 u1_u15_u0_U49 (.A( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n145 ) , .B1( u1_u15_u0_n146 ) , .ZN( u1_u15_u0_n154 ) );
  AOI21_X1 u1_u15_u0_U5 (.B2( u1_u15_u0_n131 ) , .ZN( u1_u15_u0_n134 ) , .B1( u1_u15_u0_n151 ) , .A( u1_u15_u0_n158 ) );
  AOI21_X1 u1_u15_u0_U50 (.A( u1_u15_u0_n147 ) , .B2( u1_u15_u0_n148 ) , .B1( u1_u15_u0_n149 ) , .ZN( u1_u15_u0_n153 ) );
  INV_X1 u1_u15_u0_U51 (.ZN( u1_u15_u0_n171 ) , .A( u1_u15_u0_n99 ) );
  OAI211_X1 u1_u15_u0_U52 (.C2( u1_u15_u0_n140 ) , .C1( u1_u15_u0_n161 ) , .A( u1_u15_u0_n169 ) , .B( u1_u15_u0_n98 ) , .ZN( u1_u15_u0_n99 ) );
  AOI211_X1 u1_u15_u0_U53 (.C1( u1_u15_u0_n118 ) , .A( u1_u15_u0_n123 ) , .B( u1_u15_u0_n96 ) , .C2( u1_u15_u0_n97 ) , .ZN( u1_u15_u0_n98 ) );
  INV_X1 u1_u15_u0_U54 (.ZN( u1_u15_u0_n169 ) , .A( u1_u15_u0_n91 ) );
  NOR2_X1 u1_u15_u0_U55 (.A2( u1_u15_X_4 ) , .A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n118 ) );
  NOR2_X1 u1_u15_u0_U56 (.A2( u1_u15_X_1 ) , .ZN( u1_u15_u0_n101 ) , .A1( u1_u15_u0_n163 ) );
  NOR2_X1 u1_u15_u0_U57 (.A2( u1_u15_X_3 ) , .A1( u1_u15_X_6 ) , .ZN( u1_u15_u0_n94 ) );
  NOR2_X1 u1_u15_u0_U58 (.A2( u1_u15_X_6 ) , .ZN( u1_u15_u0_n100 ) , .A1( u1_u15_u0_n162 ) );
  NAND2_X1 u1_u15_u0_U59 (.A2( u1_u15_X_4 ) , .A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n144 ) );
  NOR2_X1 u1_u15_u0_U6 (.A1( u1_u15_u0_n108 ) , .ZN( u1_u15_u0_n123 ) , .A2( u1_u15_u0_n158 ) );
  NOR2_X1 u1_u15_u0_U60 (.A2( u1_u15_X_5 ) , .ZN( u1_u15_u0_n136 ) , .A1( u1_u15_u0_n159 ) );
  NAND2_X1 u1_u15_u0_U61 (.A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n138 ) , .A2( u1_u15_u0_n159 ) );
  AND2_X1 u1_u15_u0_U62 (.A2( u1_u15_X_3 ) , .A1( u1_u15_X_6 ) , .ZN( u1_u15_u0_n102 ) );
  AND2_X1 u1_u15_u0_U63 (.A1( u1_u15_X_6 ) , .A2( u1_u15_u0_n162 ) , .ZN( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U64 (.A( u1_u15_X_4 ) , .ZN( u1_u15_u0_n159 ) );
  INV_X1 u1_u15_u0_U65 (.A( u1_u15_X_1 ) , .ZN( u1_u15_u0_n164 ) );
  INV_X1 u1_u15_u0_U66 (.A( u1_u15_X_3 ) , .ZN( u1_u15_u0_n162 ) );
  INV_X1 u1_u15_u0_U67 (.A( u1_u15_u0_n126 ) , .ZN( u1_u15_u0_n168 ) );
  AOI211_X1 u1_u15_u0_U68 (.B( u1_u15_u0_n133 ) , .A( u1_u15_u0_n134 ) , .C2( u1_u15_u0_n135 ) , .C1( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n137 ) );
  INV_X1 u1_u15_u0_U69 (.ZN( u1_u15_u0_n174 ) , .A( u1_u15_u0_n89 ) );
  OAI21_X1 u1_u15_u0_U7 (.B1( u1_u15_u0_n150 ) , .B2( u1_u15_u0_n158 ) , .A( u1_u15_u0_n172 ) , .ZN( u1_u15_u0_n89 ) );
  AOI211_X1 u1_u15_u0_U70 (.B( u1_u15_u0_n104 ) , .A( u1_u15_u0_n105 ) , .ZN( u1_u15_u0_n106 ) , .C2( u1_u15_u0_n113 ) , .C1( u1_u15_u0_n160 ) );
  OR4_X1 u1_u15_u0_U71 (.ZN( u1_out15_17 ) , .A4( u1_u15_u0_n122 ) , .A2( u1_u15_u0_n123 ) , .A1( u1_u15_u0_n124 ) , .A3( u1_u15_u0_n170 ) );
  AOI21_X1 u1_u15_u0_U72 (.B2( u1_u15_u0_n107 ) , .ZN( u1_u15_u0_n124 ) , .B1( u1_u15_u0_n128 ) , .A( u1_u15_u0_n161 ) );
  INV_X1 u1_u15_u0_U73 (.A( u1_u15_u0_n111 ) , .ZN( u1_u15_u0_n170 ) );
  OR4_X1 u1_u15_u0_U74 (.ZN( u1_out15_31 ) , .A4( u1_u15_u0_n155 ) , .A2( u1_u15_u0_n156 ) , .A1( u1_u15_u0_n157 ) , .A3( u1_u15_u0_n173 ) );
  AOI21_X1 u1_u15_u0_U75 (.A( u1_u15_u0_n138 ) , .B2( u1_u15_u0_n139 ) , .B1( u1_u15_u0_n140 ) , .ZN( u1_u15_u0_n157 ) );
  AOI21_X1 u1_u15_u0_U76 (.B2( u1_u15_u0_n141 ) , .B1( u1_u15_u0_n142 ) , .ZN( u1_u15_u0_n156 ) , .A( u1_u15_u0_n161 ) );
  AOI21_X1 u1_u15_u0_U77 (.B1( u1_u15_u0_n132 ) , .ZN( u1_u15_u0_n133 ) , .A( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n166 ) );
  OAI22_X1 u1_u15_u0_U78 (.ZN( u1_u15_u0_n105 ) , .A2( u1_u15_u0_n132 ) , .B1( u1_u15_u0_n146 ) , .A1( u1_u15_u0_n147 ) , .B2( u1_u15_u0_n161 ) );
  NAND2_X1 u1_u15_u0_U79 (.ZN( u1_u15_u0_n110 ) , .A2( u1_u15_u0_n132 ) , .A1( u1_u15_u0_n145 ) );
  AND2_X1 u1_u15_u0_U8 (.A1( u1_u15_u0_n114 ) , .A2( u1_u15_u0_n121 ) , .ZN( u1_u15_u0_n146 ) );
  INV_X1 u1_u15_u0_U80 (.A( u1_u15_u0_n119 ) , .ZN( u1_u15_u0_n167 ) );
  NAND2_X1 u1_u15_u0_U81 (.ZN( u1_u15_u0_n148 ) , .A1( u1_u15_u0_n93 ) , .A2( u1_u15_u0_n95 ) );
  NAND2_X1 u1_u15_u0_U82 (.A1( u1_u15_u0_n100 ) , .ZN( u1_u15_u0_n129 ) , .A2( u1_u15_u0_n95 ) );
  NAND2_X1 u1_u15_u0_U83 (.A1( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n128 ) , .A2( u1_u15_u0_n95 ) );
  NOR2_X1 u1_u15_u0_U84 (.A2( u1_u15_X_1 ) , .A1( u1_u15_X_2 ) , .ZN( u1_u15_u0_n92 ) );
  NAND2_X1 u1_u15_u0_U85 (.ZN( u1_u15_u0_n142 ) , .A1( u1_u15_u0_n94 ) , .A2( u1_u15_u0_n95 ) );
  NOR2_X1 u1_u15_u0_U86 (.A2( u1_u15_X_2 ) , .ZN( u1_u15_u0_n103 ) , .A1( u1_u15_u0_n164 ) );
  INV_X1 u1_u15_u0_U87 (.A( u1_u15_X_2 ) , .ZN( u1_u15_u0_n163 ) );
  NAND3_X1 u1_u15_u0_U88 (.ZN( u1_out15_23 ) , .A3( u1_u15_u0_n137 ) , .A1( u1_u15_u0_n168 ) , .A2( u1_u15_u0_n171 ) );
  NAND3_X1 u1_u15_u0_U89 (.A3( u1_u15_u0_n127 ) , .A2( u1_u15_u0_n128 ) , .ZN( u1_u15_u0_n135 ) , .A1( u1_u15_u0_n150 ) );
  AND2_X1 u1_u15_u0_U9 (.A1( u1_u15_u0_n131 ) , .ZN( u1_u15_u0_n141 ) , .A2( u1_u15_u0_n150 ) );
  NAND3_X1 u1_u15_u0_U90 (.ZN( u1_u15_u0_n117 ) , .A3( u1_u15_u0_n132 ) , .A2( u1_u15_u0_n139 ) , .A1( u1_u15_u0_n148 ) );
  NAND3_X1 u1_u15_u0_U91 (.ZN( u1_u15_u0_n109 ) , .A2( u1_u15_u0_n114 ) , .A3( u1_u15_u0_n140 ) , .A1( u1_u15_u0_n149 ) );
  NAND3_X1 u1_u15_u0_U92 (.ZN( u1_out15_9 ) , .A3( u1_u15_u0_n106 ) , .A2( u1_u15_u0_n171 ) , .A1( u1_u15_u0_n174 ) );
  NAND3_X1 u1_u15_u0_U93 (.A2( u1_u15_u0_n128 ) , .A1( u1_u15_u0_n132 ) , .A3( u1_u15_u0_n146 ) , .ZN( u1_u15_u0_n97 ) );
  AOI21_X1 u1_u15_u1_U10 (.B2( u1_u15_u1_n155 ) , .B1( u1_u15_u1_n156 ) , .ZN( u1_u15_u1_n157 ) , .A( u1_u15_u1_n174 ) );
  NAND3_X1 u1_u15_u1_U100 (.ZN( u1_u15_u1_n113 ) , .A1( u1_u15_u1_n120 ) , .A3( u1_u15_u1_n133 ) , .A2( u1_u15_u1_n155 ) );
  NAND2_X1 u1_u15_u1_U11 (.ZN( u1_u15_u1_n140 ) , .A2( u1_u15_u1_n150 ) , .A1( u1_u15_u1_n155 ) );
  NAND2_X1 u1_u15_u1_U12 (.A1( u1_u15_u1_n131 ) , .ZN( u1_u15_u1_n147 ) , .A2( u1_u15_u1_n153 ) );
  INV_X1 u1_u15_u1_U13 (.A( u1_u15_u1_n139 ) , .ZN( u1_u15_u1_n174 ) );
  OR4_X1 u1_u15_u1_U14 (.A4( u1_u15_u1_n106 ) , .A3( u1_u15_u1_n107 ) , .ZN( u1_u15_u1_n108 ) , .A1( u1_u15_u1_n117 ) , .A2( u1_u15_u1_n184 ) );
  AOI21_X1 u1_u15_u1_U15 (.ZN( u1_u15_u1_n106 ) , .A( u1_u15_u1_n112 ) , .B1( u1_u15_u1_n154 ) , .B2( u1_u15_u1_n156 ) );
  AOI21_X1 u1_u15_u1_U16 (.ZN( u1_u15_u1_n107 ) , .B1( u1_u15_u1_n134 ) , .B2( u1_u15_u1_n149 ) , .A( u1_u15_u1_n174 ) );
  INV_X1 u1_u15_u1_U17 (.A( u1_u15_u1_n101 ) , .ZN( u1_u15_u1_n184 ) );
  INV_X1 u1_u15_u1_U18 (.A( u1_u15_u1_n112 ) , .ZN( u1_u15_u1_n171 ) );
  NAND2_X1 u1_u15_u1_U19 (.ZN( u1_u15_u1_n141 ) , .A1( u1_u15_u1_n153 ) , .A2( u1_u15_u1_n156 ) );
  AND2_X1 u1_u15_u1_U20 (.A1( u1_u15_u1_n123 ) , .ZN( u1_u15_u1_n134 ) , .A2( u1_u15_u1_n161 ) );
  NAND2_X1 u1_u15_u1_U21 (.A2( u1_u15_u1_n115 ) , .A1( u1_u15_u1_n116 ) , .ZN( u1_u15_u1_n148 ) );
  NAND2_X1 u1_u15_u1_U22 (.A2( u1_u15_u1_n133 ) , .A1( u1_u15_u1_n135 ) , .ZN( u1_u15_u1_n159 ) );
  NAND2_X1 u1_u15_u1_U23 (.A2( u1_u15_u1_n115 ) , .A1( u1_u15_u1_n120 ) , .ZN( u1_u15_u1_n132 ) );
  INV_X1 u1_u15_u1_U24 (.A( u1_u15_u1_n154 ) , .ZN( u1_u15_u1_n178 ) );
  AOI22_X1 u1_u15_u1_U25 (.B2( u1_u15_u1_n113 ) , .A2( u1_u15_u1_n114 ) , .ZN( u1_u15_u1_n125 ) , .A1( u1_u15_u1_n171 ) , .B1( u1_u15_u1_n173 ) );
  NAND2_X1 u1_u15_u1_U26 (.ZN( u1_u15_u1_n114 ) , .A1( u1_u15_u1_n134 ) , .A2( u1_u15_u1_n156 ) );
  INV_X1 u1_u15_u1_U27 (.A( u1_u15_u1_n151 ) , .ZN( u1_u15_u1_n183 ) );
  AND2_X1 u1_u15_u1_U28 (.A1( u1_u15_u1_n129 ) , .A2( u1_u15_u1_n133 ) , .ZN( u1_u15_u1_n149 ) );
  INV_X1 u1_u15_u1_U29 (.A( u1_u15_u1_n131 ) , .ZN( u1_u15_u1_n180 ) );
  INV_X1 u1_u15_u1_U3 (.A( u1_u15_u1_n159 ) , .ZN( u1_u15_u1_n182 ) );
  OAI221_X1 u1_u15_u1_U30 (.A( u1_u15_u1_n119 ) , .C2( u1_u15_u1_n129 ) , .ZN( u1_u15_u1_n138 ) , .B2( u1_u15_u1_n152 ) , .C1( u1_u15_u1_n174 ) , .B1( u1_u15_u1_n187 ) );
  INV_X1 u1_u15_u1_U31 (.A( u1_u15_u1_n148 ) , .ZN( u1_u15_u1_n187 ) );
  AOI211_X1 u1_u15_u1_U32 (.B( u1_u15_u1_n117 ) , .A( u1_u15_u1_n118 ) , .ZN( u1_u15_u1_n119 ) , .C2( u1_u15_u1_n146 ) , .C1( u1_u15_u1_n159 ) );
  NOR2_X1 u1_u15_u1_U33 (.A1( u1_u15_u1_n168 ) , .A2( u1_u15_u1_n176 ) , .ZN( u1_u15_u1_n98 ) );
  AOI211_X1 u1_u15_u1_U34 (.B( u1_u15_u1_n162 ) , .A( u1_u15_u1_n163 ) , .C2( u1_u15_u1_n164 ) , .ZN( u1_u15_u1_n165 ) , .C1( u1_u15_u1_n171 ) );
  AOI21_X1 u1_u15_u1_U35 (.A( u1_u15_u1_n160 ) , .B2( u1_u15_u1_n161 ) , .ZN( u1_u15_u1_n162 ) , .B1( u1_u15_u1_n182 ) );
  OR2_X1 u1_u15_u1_U36 (.A2( u1_u15_u1_n157 ) , .A1( u1_u15_u1_n158 ) , .ZN( u1_u15_u1_n163 ) );
  NAND2_X1 u1_u15_u1_U37 (.A1( u1_u15_u1_n128 ) , .ZN( u1_u15_u1_n146 ) , .A2( u1_u15_u1_n160 ) );
  NAND2_X1 u1_u15_u1_U38 (.A2( u1_u15_u1_n112 ) , .ZN( u1_u15_u1_n139 ) , .A1( u1_u15_u1_n152 ) );
  NAND2_X1 u1_u15_u1_U39 (.A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n156 ) , .A2( u1_u15_u1_n99 ) );
  AOI221_X1 u1_u15_u1_U4 (.A( u1_u15_u1_n138 ) , .C2( u1_u15_u1_n139 ) , .C1( u1_u15_u1_n140 ) , .B2( u1_u15_u1_n141 ) , .ZN( u1_u15_u1_n142 ) , .B1( u1_u15_u1_n175 ) );
  AOI221_X1 u1_u15_u1_U40 (.B1( u1_u15_u1_n140 ) , .ZN( u1_u15_u1_n167 ) , .B2( u1_u15_u1_n172 ) , .C2( u1_u15_u1_n175 ) , .C1( u1_u15_u1_n178 ) , .A( u1_u15_u1_n188 ) );
  INV_X1 u1_u15_u1_U41 (.ZN( u1_u15_u1_n188 ) , .A( u1_u15_u1_n97 ) );
  AOI211_X1 u1_u15_u1_U42 (.A( u1_u15_u1_n118 ) , .C1( u1_u15_u1_n132 ) , .C2( u1_u15_u1_n139 ) , .B( u1_u15_u1_n96 ) , .ZN( u1_u15_u1_n97 ) );
  AOI21_X1 u1_u15_u1_U43 (.B2( u1_u15_u1_n121 ) , .B1( u1_u15_u1_n135 ) , .A( u1_u15_u1_n152 ) , .ZN( u1_u15_u1_n96 ) );
  NOR2_X1 u1_u15_u1_U44 (.ZN( u1_u15_u1_n117 ) , .A1( u1_u15_u1_n121 ) , .A2( u1_u15_u1_n160 ) );
  AOI21_X1 u1_u15_u1_U45 (.A( u1_u15_u1_n128 ) , .B2( u1_u15_u1_n129 ) , .ZN( u1_u15_u1_n130 ) , .B1( u1_u15_u1_n150 ) );
  OAI21_X1 u1_u15_u1_U46 (.B2( u1_u15_u1_n123 ) , .ZN( u1_u15_u1_n145 ) , .B1( u1_u15_u1_n160 ) , .A( u1_u15_u1_n185 ) );
  INV_X1 u1_u15_u1_U47 (.A( u1_u15_u1_n122 ) , .ZN( u1_u15_u1_n185 ) );
  AOI21_X1 u1_u15_u1_U48 (.B2( u1_u15_u1_n120 ) , .B1( u1_u15_u1_n121 ) , .ZN( u1_u15_u1_n122 ) , .A( u1_u15_u1_n128 ) );
  NAND2_X1 u1_u15_u1_U49 (.ZN( u1_u15_u1_n112 ) , .A1( u1_u15_u1_n169 ) , .A2( u1_u15_u1_n170 ) );
  AOI211_X1 u1_u15_u1_U5 (.ZN( u1_u15_u1_n124 ) , .A( u1_u15_u1_n138 ) , .C2( u1_u15_u1_n139 ) , .B( u1_u15_u1_n145 ) , .C1( u1_u15_u1_n147 ) );
  NAND2_X1 u1_u15_u1_U50 (.ZN( u1_u15_u1_n129 ) , .A2( u1_u15_u1_n95 ) , .A1( u1_u15_u1_n98 ) );
  NAND2_X1 u1_u15_u1_U51 (.A1( u1_u15_u1_n102 ) , .ZN( u1_u15_u1_n154 ) , .A2( u1_u15_u1_n99 ) );
  NAND2_X1 u1_u15_u1_U52 (.A2( u1_u15_u1_n100 ) , .ZN( u1_u15_u1_n135 ) , .A1( u1_u15_u1_n99 ) );
  AOI21_X1 u1_u15_u1_U53 (.A( u1_u15_u1_n152 ) , .B2( u1_u15_u1_n153 ) , .B1( u1_u15_u1_n154 ) , .ZN( u1_u15_u1_n158 ) );
  INV_X1 u1_u15_u1_U54 (.A( u1_u15_u1_n160 ) , .ZN( u1_u15_u1_n175 ) );
  NAND2_X1 u1_u15_u1_U55 (.A1( u1_u15_u1_n100 ) , .ZN( u1_u15_u1_n116 ) , .A2( u1_u15_u1_n95 ) );
  NAND2_X1 u1_u15_u1_U56 (.A1( u1_u15_u1_n102 ) , .ZN( u1_u15_u1_n131 ) , .A2( u1_u15_u1_n95 ) );
  NAND2_X1 u1_u15_u1_U57 (.A2( u1_u15_u1_n104 ) , .ZN( u1_u15_u1_n121 ) , .A1( u1_u15_u1_n98 ) );
  NAND2_X1 u1_u15_u1_U58 (.A1( u1_u15_u1_n103 ) , .ZN( u1_u15_u1_n153 ) , .A2( u1_u15_u1_n98 ) );
  NAND2_X1 u1_u15_u1_U59 (.A2( u1_u15_u1_n104 ) , .A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n133 ) );
  AOI22_X1 u1_u15_u1_U6 (.B2( u1_u15_u1_n136 ) , .A2( u1_u15_u1_n137 ) , .ZN( u1_u15_u1_n143 ) , .A1( u1_u15_u1_n171 ) , .B1( u1_u15_u1_n173 ) );
  NAND2_X1 u1_u15_u1_U60 (.ZN( u1_u15_u1_n150 ) , .A2( u1_u15_u1_n98 ) , .A1( u1_u15_u1_n99 ) );
  NAND2_X1 u1_u15_u1_U61 (.A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n155 ) , .A2( u1_u15_u1_n95 ) );
  OAI21_X1 u1_u15_u1_U62 (.ZN( u1_u15_u1_n109 ) , .B1( u1_u15_u1_n129 ) , .B2( u1_u15_u1_n160 ) , .A( u1_u15_u1_n167 ) );
  NAND2_X1 u1_u15_u1_U63 (.A2( u1_u15_u1_n100 ) , .A1( u1_u15_u1_n103 ) , .ZN( u1_u15_u1_n120 ) );
  NAND2_X1 u1_u15_u1_U64 (.A1( u1_u15_u1_n102 ) , .A2( u1_u15_u1_n104 ) , .ZN( u1_u15_u1_n115 ) );
  NAND2_X1 u1_u15_u1_U65 (.A2( u1_u15_u1_n100 ) , .A1( u1_u15_u1_n104 ) , .ZN( u1_u15_u1_n151 ) );
  NAND2_X1 u1_u15_u1_U66 (.A2( u1_u15_u1_n103 ) , .A1( u1_u15_u1_n105 ) , .ZN( u1_u15_u1_n161 ) );
  INV_X1 u1_u15_u1_U67 (.A( u1_u15_u1_n152 ) , .ZN( u1_u15_u1_n173 ) );
  INV_X1 u1_u15_u1_U68 (.A( u1_u15_u1_n128 ) , .ZN( u1_u15_u1_n172 ) );
  NAND2_X1 u1_u15_u1_U69 (.A2( u1_u15_u1_n102 ) , .A1( u1_u15_u1_n103 ) , .ZN( u1_u15_u1_n123 ) );
  INV_X1 u1_u15_u1_U7 (.A( u1_u15_u1_n147 ) , .ZN( u1_u15_u1_n181 ) );
  NOR2_X1 u1_u15_u1_U70 (.A2( u1_u15_X_7 ) , .A1( u1_u15_X_8 ) , .ZN( u1_u15_u1_n95 ) );
  NOR2_X1 u1_u15_u1_U71 (.A1( u1_u15_X_12 ) , .A2( u1_u15_X_9 ) , .ZN( u1_u15_u1_n100 ) );
  NOR2_X1 u1_u15_u1_U72 (.A2( u1_u15_X_8 ) , .A1( u1_u15_u1_n177 ) , .ZN( u1_u15_u1_n99 ) );
  NOR2_X1 u1_u15_u1_U73 (.A2( u1_u15_X_12 ) , .ZN( u1_u15_u1_n102 ) , .A1( u1_u15_u1_n176 ) );
  NOR2_X1 u1_u15_u1_U74 (.A2( u1_u15_X_9 ) , .ZN( u1_u15_u1_n105 ) , .A1( u1_u15_u1_n168 ) );
  NAND2_X1 u1_u15_u1_U75 (.A1( u1_u15_X_10 ) , .ZN( u1_u15_u1_n160 ) , .A2( u1_u15_u1_n169 ) );
  NAND2_X1 u1_u15_u1_U76 (.A2( u1_u15_X_10 ) , .A1( u1_u15_X_11 ) , .ZN( u1_u15_u1_n152 ) );
  NAND2_X1 u1_u15_u1_U77 (.A1( u1_u15_X_11 ) , .ZN( u1_u15_u1_n128 ) , .A2( u1_u15_u1_n170 ) );
  AND2_X1 u1_u15_u1_U78 (.A2( u1_u15_X_7 ) , .A1( u1_u15_X_8 ) , .ZN( u1_u15_u1_n104 ) );
  AND2_X1 u1_u15_u1_U79 (.A1( u1_u15_X_8 ) , .ZN( u1_u15_u1_n103 ) , .A2( u1_u15_u1_n177 ) );
  NOR2_X1 u1_u15_u1_U8 (.A1( u1_u15_u1_n112 ) , .A2( u1_u15_u1_n116 ) , .ZN( u1_u15_u1_n118 ) );
  INV_X1 u1_u15_u1_U80 (.A( u1_u15_X_10 ) , .ZN( u1_u15_u1_n170 ) );
  INV_X1 u1_u15_u1_U81 (.A( u1_u15_X_9 ) , .ZN( u1_u15_u1_n176 ) );
  INV_X1 u1_u15_u1_U82 (.A( u1_u15_X_11 ) , .ZN( u1_u15_u1_n169 ) );
  INV_X1 u1_u15_u1_U83 (.A( u1_u15_X_12 ) , .ZN( u1_u15_u1_n168 ) );
  INV_X1 u1_u15_u1_U84 (.A( u1_u15_X_7 ) , .ZN( u1_u15_u1_n177 ) );
  NAND4_X1 u1_u15_u1_U85 (.ZN( u1_out15_18 ) , .A4( u1_u15_u1_n165 ) , .A3( u1_u15_u1_n166 ) , .A1( u1_u15_u1_n167 ) , .A2( u1_u15_u1_n186 ) );
  AOI22_X1 u1_u15_u1_U86 (.B2( u1_u15_u1_n146 ) , .B1( u1_u15_u1_n147 ) , .A2( u1_u15_u1_n148 ) , .ZN( u1_u15_u1_n166 ) , .A1( u1_u15_u1_n172 ) );
  INV_X1 u1_u15_u1_U87 (.A( u1_u15_u1_n145 ) , .ZN( u1_u15_u1_n186 ) );
  NAND4_X1 u1_u15_u1_U88 (.ZN( u1_out15_2 ) , .A4( u1_u15_u1_n142 ) , .A3( u1_u15_u1_n143 ) , .A2( u1_u15_u1_n144 ) , .A1( u1_u15_u1_n179 ) );
  OAI21_X1 u1_u15_u1_U89 (.B2( u1_u15_u1_n132 ) , .ZN( u1_u15_u1_n144 ) , .A( u1_u15_u1_n146 ) , .B1( u1_u15_u1_n180 ) );
  OAI21_X1 u1_u15_u1_U9 (.ZN( u1_u15_u1_n101 ) , .B1( u1_u15_u1_n141 ) , .A( u1_u15_u1_n146 ) , .B2( u1_u15_u1_n183 ) );
  INV_X1 u1_u15_u1_U90 (.A( u1_u15_u1_n130 ) , .ZN( u1_u15_u1_n179 ) );
  NAND4_X1 u1_u15_u1_U91 (.ZN( u1_out15_28 ) , .A4( u1_u15_u1_n124 ) , .A3( u1_u15_u1_n125 ) , .A2( u1_u15_u1_n126 ) , .A1( u1_u15_u1_n127 ) );
  OAI21_X1 u1_u15_u1_U92 (.ZN( u1_u15_u1_n127 ) , .B2( u1_u15_u1_n139 ) , .B1( u1_u15_u1_n175 ) , .A( u1_u15_u1_n183 ) );
  OAI21_X1 u1_u15_u1_U93 (.ZN( u1_u15_u1_n126 ) , .B2( u1_u15_u1_n140 ) , .A( u1_u15_u1_n146 ) , .B1( u1_u15_u1_n178 ) );
  OR4_X1 u1_u15_u1_U94 (.ZN( u1_out15_13 ) , .A4( u1_u15_u1_n108 ) , .A3( u1_u15_u1_n109 ) , .A2( u1_u15_u1_n110 ) , .A1( u1_u15_u1_n111 ) );
  AOI21_X1 u1_u15_u1_U95 (.ZN( u1_u15_u1_n111 ) , .A( u1_u15_u1_n128 ) , .B2( u1_u15_u1_n131 ) , .B1( u1_u15_u1_n135 ) );
  AOI21_X1 u1_u15_u1_U96 (.ZN( u1_u15_u1_n110 ) , .A( u1_u15_u1_n116 ) , .B1( u1_u15_u1_n152 ) , .B2( u1_u15_u1_n160 ) );
  NAND3_X1 u1_u15_u1_U97 (.A3( u1_u15_u1_n149 ) , .A2( u1_u15_u1_n150 ) , .A1( u1_u15_u1_n151 ) , .ZN( u1_u15_u1_n164 ) );
  NAND3_X1 u1_u15_u1_U98 (.A3( u1_u15_u1_n134 ) , .A2( u1_u15_u1_n135 ) , .ZN( u1_u15_u1_n136 ) , .A1( u1_u15_u1_n151 ) );
  NAND3_X1 u1_u15_u1_U99 (.A1( u1_u15_u1_n133 ) , .ZN( u1_u15_u1_n137 ) , .A2( u1_u15_u1_n154 ) , .A3( u1_u15_u1_n181 ) );
  OAI22_X1 u1_u15_u3_U10 (.B1( u1_u15_u3_n113 ) , .A2( u1_u15_u3_n135 ) , .A1( u1_u15_u3_n150 ) , .B2( u1_u15_u3_n164 ) , .ZN( u1_u15_u3_n98 ) );
  OAI211_X1 u1_u15_u3_U11 (.B( u1_u15_u3_n106 ) , .ZN( u1_u15_u3_n119 ) , .C2( u1_u15_u3_n128 ) , .C1( u1_u15_u3_n167 ) , .A( u1_u15_u3_n181 ) );
  AOI221_X1 u1_u15_u3_U12 (.C1( u1_u15_u3_n105 ) , .ZN( u1_u15_u3_n106 ) , .A( u1_u15_u3_n131 ) , .B2( u1_u15_u3_n132 ) , .C2( u1_u15_u3_n133 ) , .B1( u1_u15_u3_n169 ) );
  INV_X1 u1_u15_u3_U13 (.ZN( u1_u15_u3_n181 ) , .A( u1_u15_u3_n98 ) );
  NAND2_X1 u1_u15_u3_U14 (.ZN( u1_u15_u3_n105 ) , .A2( u1_u15_u3_n130 ) , .A1( u1_u15_u3_n155 ) );
  AOI22_X1 u1_u15_u3_U15 (.B1( u1_u15_u3_n115 ) , .A2( u1_u15_u3_n116 ) , .ZN( u1_u15_u3_n123 ) , .B2( u1_u15_u3_n133 ) , .A1( u1_u15_u3_n169 ) );
  NAND2_X1 u1_u15_u3_U16 (.ZN( u1_u15_u3_n116 ) , .A2( u1_u15_u3_n151 ) , .A1( u1_u15_u3_n182 ) );
  NOR2_X1 u1_u15_u3_U17 (.ZN( u1_u15_u3_n126 ) , .A2( u1_u15_u3_n150 ) , .A1( u1_u15_u3_n164 ) );
  AOI21_X1 u1_u15_u3_U18 (.ZN( u1_u15_u3_n112 ) , .B2( u1_u15_u3_n146 ) , .B1( u1_u15_u3_n155 ) , .A( u1_u15_u3_n167 ) );
  NAND2_X1 u1_u15_u3_U19 (.A1( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n142 ) , .A2( u1_u15_u3_n164 ) );
  NAND2_X1 u1_u15_u3_U20 (.ZN( u1_u15_u3_n132 ) , .A2( u1_u15_u3_n152 ) , .A1( u1_u15_u3_n156 ) );
  AND2_X1 u1_u15_u3_U21 (.A2( u1_u15_u3_n113 ) , .A1( u1_u15_u3_n114 ) , .ZN( u1_u15_u3_n151 ) );
  INV_X1 u1_u15_u3_U22 (.A( u1_u15_u3_n133 ) , .ZN( u1_u15_u3_n165 ) );
  INV_X1 u1_u15_u3_U23 (.A( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n170 ) );
  NAND2_X1 u1_u15_u3_U24 (.A1( u1_u15_u3_n107 ) , .A2( u1_u15_u3_n108 ) , .ZN( u1_u15_u3_n140 ) );
  NAND2_X1 u1_u15_u3_U25 (.ZN( u1_u15_u3_n117 ) , .A1( u1_u15_u3_n124 ) , .A2( u1_u15_u3_n148 ) );
  NAND2_X1 u1_u15_u3_U26 (.ZN( u1_u15_u3_n143 ) , .A1( u1_u15_u3_n165 ) , .A2( u1_u15_u3_n167 ) );
  INV_X1 u1_u15_u3_U27 (.A( u1_u15_u3_n130 ) , .ZN( u1_u15_u3_n177 ) );
  INV_X1 u1_u15_u3_U28 (.A( u1_u15_u3_n128 ) , .ZN( u1_u15_u3_n176 ) );
  INV_X1 u1_u15_u3_U29 (.A( u1_u15_u3_n155 ) , .ZN( u1_u15_u3_n174 ) );
  INV_X1 u1_u15_u3_U3 (.A( u1_u15_u3_n129 ) , .ZN( u1_u15_u3_n183 ) );
  INV_X1 u1_u15_u3_U30 (.A( u1_u15_u3_n139 ) , .ZN( u1_u15_u3_n185 ) );
  NOR2_X1 u1_u15_u3_U31 (.ZN( u1_u15_u3_n135 ) , .A2( u1_u15_u3_n141 ) , .A1( u1_u15_u3_n169 ) );
  OAI222_X1 u1_u15_u3_U32 (.C2( u1_u15_u3_n107 ) , .A2( u1_u15_u3_n108 ) , .B1( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n138 ) , .B2( u1_u15_u3_n146 ) , .C1( u1_u15_u3_n154 ) , .A1( u1_u15_u3_n164 ) );
  NOR4_X1 u1_u15_u3_U33 (.A4( u1_u15_u3_n157 ) , .A3( u1_u15_u3_n158 ) , .A2( u1_u15_u3_n159 ) , .A1( u1_u15_u3_n160 ) , .ZN( u1_u15_u3_n161 ) );
  AOI21_X1 u1_u15_u3_U34 (.B2( u1_u15_u3_n152 ) , .B1( u1_u15_u3_n153 ) , .ZN( u1_u15_u3_n158 ) , .A( u1_u15_u3_n164 ) );
  AOI21_X1 u1_u15_u3_U35 (.A( u1_u15_u3_n154 ) , .B2( u1_u15_u3_n155 ) , .B1( u1_u15_u3_n156 ) , .ZN( u1_u15_u3_n157 ) );
  AOI21_X1 u1_u15_u3_U36 (.A( u1_u15_u3_n149 ) , .B2( u1_u15_u3_n150 ) , .B1( u1_u15_u3_n151 ) , .ZN( u1_u15_u3_n159 ) );
  AOI211_X1 u1_u15_u3_U37 (.ZN( u1_u15_u3_n109 ) , .A( u1_u15_u3_n119 ) , .C2( u1_u15_u3_n129 ) , .B( u1_u15_u3_n138 ) , .C1( u1_u15_u3_n141 ) );
  AOI211_X1 u1_u15_u3_U38 (.B( u1_u15_u3_n119 ) , .A( u1_u15_u3_n120 ) , .C2( u1_u15_u3_n121 ) , .ZN( u1_u15_u3_n122 ) , .C1( u1_u15_u3_n179 ) );
  INV_X1 u1_u15_u3_U39 (.A( u1_u15_u3_n156 ) , .ZN( u1_u15_u3_n179 ) );
  INV_X1 u1_u15_u3_U4 (.A( u1_u15_u3_n140 ) , .ZN( u1_u15_u3_n182 ) );
  OAI22_X1 u1_u15_u3_U40 (.B1( u1_u15_u3_n118 ) , .ZN( u1_u15_u3_n120 ) , .A1( u1_u15_u3_n135 ) , .B2( u1_u15_u3_n154 ) , .A2( u1_u15_u3_n178 ) );
  AND3_X1 u1_u15_u3_U41 (.ZN( u1_u15_u3_n118 ) , .A2( u1_u15_u3_n124 ) , .A1( u1_u15_u3_n144 ) , .A3( u1_u15_u3_n152 ) );
  INV_X1 u1_u15_u3_U42 (.A( u1_u15_u3_n121 ) , .ZN( u1_u15_u3_n164 ) );
  NAND2_X1 u1_u15_u3_U43 (.ZN( u1_u15_u3_n133 ) , .A1( u1_u15_u3_n154 ) , .A2( u1_u15_u3_n164 ) );
  OAI211_X1 u1_u15_u3_U44 (.B( u1_u15_u3_n127 ) , .ZN( u1_u15_u3_n139 ) , .C1( u1_u15_u3_n150 ) , .C2( u1_u15_u3_n154 ) , .A( u1_u15_u3_n184 ) );
  INV_X1 u1_u15_u3_U45 (.A( u1_u15_u3_n125 ) , .ZN( u1_u15_u3_n184 ) );
  AOI221_X1 u1_u15_u3_U46 (.A( u1_u15_u3_n126 ) , .ZN( u1_u15_u3_n127 ) , .C2( u1_u15_u3_n132 ) , .C1( u1_u15_u3_n169 ) , .B2( u1_u15_u3_n170 ) , .B1( u1_u15_u3_n174 ) );
  OAI22_X1 u1_u15_u3_U47 (.A1( u1_u15_u3_n124 ) , .ZN( u1_u15_u3_n125 ) , .B2( u1_u15_u3_n145 ) , .A2( u1_u15_u3_n165 ) , .B1( u1_u15_u3_n167 ) );
  NOR2_X1 u1_u15_u3_U48 (.A1( u1_u15_u3_n113 ) , .ZN( u1_u15_u3_n131 ) , .A2( u1_u15_u3_n154 ) );
  NAND2_X1 u1_u15_u3_U49 (.A1( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n150 ) , .A2( u1_u15_u3_n99 ) );
  INV_X1 u1_u15_u3_U5 (.A( u1_u15_u3_n117 ) , .ZN( u1_u15_u3_n178 ) );
  NAND2_X1 u1_u15_u3_U50 (.A2( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n155 ) , .A1( u1_u15_u3_n97 ) );
  INV_X1 u1_u15_u3_U51 (.A( u1_u15_u3_n141 ) , .ZN( u1_u15_u3_n167 ) );
  AOI21_X1 u1_u15_u3_U52 (.B2( u1_u15_u3_n114 ) , .B1( u1_u15_u3_n146 ) , .A( u1_u15_u3_n154 ) , .ZN( u1_u15_u3_n94 ) );
  AOI21_X1 u1_u15_u3_U53 (.ZN( u1_u15_u3_n110 ) , .B2( u1_u15_u3_n142 ) , .B1( u1_u15_u3_n186 ) , .A( u1_u15_u3_n95 ) );
  INV_X1 u1_u15_u3_U54 (.A( u1_u15_u3_n145 ) , .ZN( u1_u15_u3_n186 ) );
  AOI21_X1 u1_u15_u3_U55 (.B1( u1_u15_u3_n124 ) , .A( u1_u15_u3_n149 ) , .B2( u1_u15_u3_n155 ) , .ZN( u1_u15_u3_n95 ) );
  INV_X1 u1_u15_u3_U56 (.A( u1_u15_u3_n149 ) , .ZN( u1_u15_u3_n169 ) );
  NAND2_X1 u1_u15_u3_U57 (.ZN( u1_u15_u3_n124 ) , .A1( u1_u15_u3_n96 ) , .A2( u1_u15_u3_n97 ) );
  NAND2_X1 u1_u15_u3_U58 (.A2( u1_u15_u3_n100 ) , .ZN( u1_u15_u3_n146 ) , .A1( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U59 (.A1( u1_u15_u3_n101 ) , .ZN( u1_u15_u3_n145 ) , .A2( u1_u15_u3_n99 ) );
  AOI221_X1 u1_u15_u3_U6 (.A( u1_u15_u3_n131 ) , .C2( u1_u15_u3_n132 ) , .C1( u1_u15_u3_n133 ) , .ZN( u1_u15_u3_n134 ) , .B1( u1_u15_u3_n143 ) , .B2( u1_u15_u3_n177 ) );
  NAND2_X1 u1_u15_u3_U60 (.A1( u1_u15_u3_n100 ) , .ZN( u1_u15_u3_n156 ) , .A2( u1_u15_u3_n99 ) );
  NAND2_X1 u1_u15_u3_U61 (.A2( u1_u15_u3_n101 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n148 ) );
  NAND2_X1 u1_u15_u3_U62 (.A1( u1_u15_u3_n100 ) , .A2( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n128 ) );
  NAND2_X1 u1_u15_u3_U63 (.A2( u1_u15_u3_n101 ) , .A1( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n152 ) );
  NAND2_X1 u1_u15_u3_U64 (.A2( u1_u15_u3_n101 ) , .ZN( u1_u15_u3_n114 ) , .A1( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U65 (.ZN( u1_u15_u3_n107 ) , .A1( u1_u15_u3_n97 ) , .A2( u1_u15_u3_n99 ) );
  NAND2_X1 u1_u15_u3_U66 (.A2( u1_u15_u3_n100 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n113 ) );
  NAND2_X1 u1_u15_u3_U67 (.A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n153 ) , .A2( u1_u15_u3_n97 ) );
  NAND2_X1 u1_u15_u3_U68 (.A2( u1_u15_u3_n103 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n130 ) );
  NAND2_X1 u1_u15_u3_U69 (.A2( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n144 ) , .A1( u1_u15_u3_n96 ) );
  OAI22_X1 u1_u15_u3_U7 (.B2( u1_u15_u3_n147 ) , .A2( u1_u15_u3_n148 ) , .ZN( u1_u15_u3_n160 ) , .B1( u1_u15_u3_n165 ) , .A1( u1_u15_u3_n168 ) );
  NAND2_X1 u1_u15_u3_U70 (.A1( u1_u15_u3_n102 ) , .A2( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n108 ) );
  NOR2_X1 u1_u15_u3_U71 (.A2( u1_u15_X_19 ) , .A1( u1_u15_X_20 ) , .ZN( u1_u15_u3_n99 ) );
  NOR2_X1 u1_u15_u3_U72 (.A2( u1_u15_X_21 ) , .A1( u1_u15_X_24 ) , .ZN( u1_u15_u3_n103 ) );
  NOR2_X1 u1_u15_u3_U73 (.A2( u1_u15_X_24 ) , .A1( u1_u15_u3_n171 ) , .ZN( u1_u15_u3_n97 ) );
  NOR2_X1 u1_u15_u3_U74 (.A2( u1_u15_X_23 ) , .ZN( u1_u15_u3_n141 ) , .A1( u1_u15_u3_n166 ) );
  NOR2_X1 u1_u15_u3_U75 (.A2( u1_u15_X_19 ) , .A1( u1_u15_u3_n172 ) , .ZN( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U76 (.A1( u1_u15_X_22 ) , .A2( u1_u15_X_23 ) , .ZN( u1_u15_u3_n154 ) );
  NAND2_X1 u1_u15_u3_U77 (.A1( u1_u15_X_23 ) , .ZN( u1_u15_u3_n149 ) , .A2( u1_u15_u3_n166 ) );
  NOR2_X1 u1_u15_u3_U78 (.A2( u1_u15_X_22 ) , .A1( u1_u15_X_23 ) , .ZN( u1_u15_u3_n121 ) );
  AND2_X1 u1_u15_u3_U79 (.A1( u1_u15_X_24 ) , .ZN( u1_u15_u3_n101 ) , .A2( u1_u15_u3_n171 ) );
  AND3_X1 u1_u15_u3_U8 (.A3( u1_u15_u3_n144 ) , .A2( u1_u15_u3_n145 ) , .A1( u1_u15_u3_n146 ) , .ZN( u1_u15_u3_n147 ) );
  AND2_X1 u1_u15_u3_U80 (.A1( u1_u15_X_19 ) , .ZN( u1_u15_u3_n102 ) , .A2( u1_u15_u3_n172 ) );
  AND2_X1 u1_u15_u3_U81 (.A1( u1_u15_X_21 ) , .A2( u1_u15_X_24 ) , .ZN( u1_u15_u3_n100 ) );
  AND2_X1 u1_u15_u3_U82 (.A2( u1_u15_X_19 ) , .A1( u1_u15_X_20 ) , .ZN( u1_u15_u3_n104 ) );
  INV_X1 u1_u15_u3_U83 (.A( u1_u15_X_22 ) , .ZN( u1_u15_u3_n166 ) );
  INV_X1 u1_u15_u3_U84 (.A( u1_u15_X_21 ) , .ZN( u1_u15_u3_n171 ) );
  INV_X1 u1_u15_u3_U85 (.A( u1_u15_X_20 ) , .ZN( u1_u15_u3_n172 ) );
  OR4_X1 u1_u15_u3_U86 (.ZN( u1_out15_10 ) , .A4( u1_u15_u3_n136 ) , .A3( u1_u15_u3_n137 ) , .A1( u1_u15_u3_n138 ) , .A2( u1_u15_u3_n139 ) );
  OAI222_X1 u1_u15_u3_U87 (.C1( u1_u15_u3_n128 ) , .ZN( u1_u15_u3_n137 ) , .B1( u1_u15_u3_n148 ) , .A2( u1_u15_u3_n150 ) , .B2( u1_u15_u3_n154 ) , .C2( u1_u15_u3_n164 ) , .A1( u1_u15_u3_n167 ) );
  OAI221_X1 u1_u15_u3_U88 (.A( u1_u15_u3_n134 ) , .B2( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n136 ) , .C1( u1_u15_u3_n149 ) , .B1( u1_u15_u3_n151 ) , .C2( u1_u15_u3_n183 ) );
  NAND4_X1 u1_u15_u3_U89 (.ZN( u1_out15_1 ) , .A4( u1_u15_u3_n161 ) , .A3( u1_u15_u3_n162 ) , .A2( u1_u15_u3_n163 ) , .A1( u1_u15_u3_n185 ) );
  INV_X1 u1_u15_u3_U9 (.A( u1_u15_u3_n143 ) , .ZN( u1_u15_u3_n168 ) );
  NAND2_X1 u1_u15_u3_U90 (.ZN( u1_u15_u3_n163 ) , .A2( u1_u15_u3_n170 ) , .A1( u1_u15_u3_n176 ) );
  AOI22_X1 u1_u15_u3_U91 (.B2( u1_u15_u3_n140 ) , .B1( u1_u15_u3_n141 ) , .A2( u1_u15_u3_n142 ) , .ZN( u1_u15_u3_n162 ) , .A1( u1_u15_u3_n177 ) );
  NAND4_X1 u1_u15_u3_U92 (.ZN( u1_out15_26 ) , .A4( u1_u15_u3_n109 ) , .A3( u1_u15_u3_n110 ) , .A2( u1_u15_u3_n111 ) , .A1( u1_u15_u3_n173 ) );
  INV_X1 u1_u15_u3_U93 (.ZN( u1_u15_u3_n173 ) , .A( u1_u15_u3_n94 ) );
  OAI21_X1 u1_u15_u3_U94 (.ZN( u1_u15_u3_n111 ) , .B2( u1_u15_u3_n117 ) , .A( u1_u15_u3_n133 ) , .B1( u1_u15_u3_n176 ) );
  NAND4_X1 u1_u15_u3_U95 (.ZN( u1_out15_20 ) , .A4( u1_u15_u3_n122 ) , .A3( u1_u15_u3_n123 ) , .A1( u1_u15_u3_n175 ) , .A2( u1_u15_u3_n180 ) );
  INV_X1 u1_u15_u3_U96 (.A( u1_u15_u3_n126 ) , .ZN( u1_u15_u3_n180 ) );
  INV_X1 u1_u15_u3_U97 (.A( u1_u15_u3_n112 ) , .ZN( u1_u15_u3_n175 ) );
  NAND3_X1 u1_u15_u3_U98 (.A1( u1_u15_u3_n114 ) , .ZN( u1_u15_u3_n115 ) , .A2( u1_u15_u3_n145 ) , .A3( u1_u15_u3_n153 ) );
  NAND3_X1 u1_u15_u3_U99 (.ZN( u1_u15_u3_n129 ) , .A2( u1_u15_u3_n144 ) , .A1( u1_u15_u3_n153 ) , .A3( u1_u15_u3_n182 ) );
  XOR2_X1 u1_u3_U10 (.B( u1_K4_45 ) , .A( u1_R2_30 ) , .Z( u1_u3_X_45 ) );
  XOR2_X1 u1_u3_U11 (.B( u1_K4_44 ) , .A( u1_R2_29 ) , .Z( u1_u3_X_44 ) );
  XOR2_X1 u1_u3_U12 (.B( u1_K4_43 ) , .A( u1_R2_28 ) , .Z( u1_u3_X_43 ) );
  XOR2_X1 u1_u3_U16 (.B( u1_K4_3 ) , .A( u1_R2_2 ) , .Z( u1_u3_X_3 ) );
  XOR2_X1 u1_u3_U27 (.B( u1_K4_2 ) , .A( u1_R2_1 ) , .Z( u1_u3_X_2 ) );
  XOR2_X1 u1_u3_U33 (.B( u1_K4_24 ) , .A( u1_R2_17 ) , .Z( u1_u3_X_24 ) );
  XOR2_X1 u1_u3_U34 (.B( u1_K4_23 ) , .A( u1_R2_16 ) , .Z( u1_u3_X_23 ) );
  XOR2_X1 u1_u3_U35 (.B( u1_K4_22 ) , .A( u1_R2_15 ) , .Z( u1_u3_X_22 ) );
  XOR2_X1 u1_u3_U36 (.B( u1_K4_21 ) , .A( u1_R2_14 ) , .Z( u1_u3_X_21 ) );
  XOR2_X1 u1_u3_U37 (.B( u1_K4_20 ) , .A( u1_R2_13 ) , .Z( u1_u3_X_20 ) );
  XOR2_X1 u1_u3_U38 (.B( u1_K4_1 ) , .A( u1_R2_32 ) , .Z( u1_u3_X_1 ) );
  XOR2_X1 u1_u3_U39 (.B( u1_K4_19 ) , .A( u1_R2_12 ) , .Z( u1_u3_X_19 ) );
  XOR2_X1 u1_u3_U4 (.B( u1_K4_6 ) , .A( u1_R2_5 ) , .Z( u1_u3_X_6 ) );
  XOR2_X1 u1_u3_U40 (.B( u1_K4_18 ) , .A( u1_R2_13 ) , .Z( u1_u3_X_18 ) );
  XOR2_X1 u1_u3_U41 (.B( u1_K4_17 ) , .A( u1_R2_12 ) , .Z( u1_u3_X_17 ) );
  XOR2_X1 u1_u3_U42 (.B( u1_K4_16 ) , .A( u1_R2_11 ) , .Z( u1_u3_X_16 ) );
  XOR2_X1 u1_u3_U43 (.B( u1_K4_15 ) , .A( u1_R2_10 ) , .Z( u1_u3_X_15 ) );
  XOR2_X1 u1_u3_U44 (.B( u1_K4_14 ) , .A( u1_R2_9 ) , .Z( u1_u3_X_14 ) );
  XOR2_X1 u1_u3_U45 (.B( u1_K4_13 ) , .A( u1_R2_8 ) , .Z( u1_u3_X_13 ) );
  XOR2_X1 u1_u3_U5 (.B( u1_K4_5 ) , .A( u1_R2_4 ) , .Z( u1_u3_X_5 ) );
  XOR2_X1 u1_u3_U6 (.B( u1_K4_4 ) , .A( u1_R2_3 ) , .Z( u1_u3_X_4 ) );
  XOR2_X1 u1_u3_U7 (.B( u1_K4_48 ) , .A( u1_R2_1 ) , .Z( u1_u3_X_48 ) );
  XOR2_X1 u1_u3_U8 (.B( u1_K4_47 ) , .A( u1_R2_32 ) , .Z( u1_u3_X_47 ) );
  XOR2_X1 u1_u3_U9 (.B( u1_K4_46 ) , .A( u1_R2_31 ) , .Z( u1_u3_X_46 ) );
  AND2_X1 u1_u3_u0_U10 (.A1( u1_u3_u0_n131 ) , .ZN( u1_u3_u0_n141 ) , .A2( u1_u3_u0_n150 ) );
  AND3_X1 u1_u3_u0_U11 (.A2( u1_u3_u0_n112 ) , .ZN( u1_u3_u0_n127 ) , .A3( u1_u3_u0_n130 ) , .A1( u1_u3_u0_n148 ) );
  AND2_X1 u1_u3_u0_U12 (.ZN( u1_u3_u0_n107 ) , .A1( u1_u3_u0_n130 ) , .A2( u1_u3_u0_n140 ) );
  AND2_X1 u1_u3_u0_U13 (.A2( u1_u3_u0_n129 ) , .A1( u1_u3_u0_n130 ) , .ZN( u1_u3_u0_n151 ) );
  AND2_X1 u1_u3_u0_U14 (.A1( u1_u3_u0_n108 ) , .A2( u1_u3_u0_n125 ) , .ZN( u1_u3_u0_n145 ) );
  INV_X1 u1_u3_u0_U15 (.A( u1_u3_u0_n143 ) , .ZN( u1_u3_u0_n173 ) );
  NOR2_X1 u1_u3_u0_U16 (.A2( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n147 ) , .A1( u1_u3_u0_n160 ) );
  AOI21_X1 u1_u3_u0_U17 (.B1( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n132 ) , .A( u1_u3_u0_n165 ) , .B2( u1_u3_u0_n93 ) );
  OAI22_X1 u1_u3_u0_U18 (.B1( u1_u3_u0_n131 ) , .A1( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n147 ) , .A2( u1_u3_u0_n90 ) , .ZN( u1_u3_u0_n91 ) );
  AND3_X1 u1_u3_u0_U19 (.A3( u1_u3_u0_n121 ) , .A2( u1_u3_u0_n125 ) , .A1( u1_u3_u0_n148 ) , .ZN( u1_u3_u0_n90 ) );
  OAI22_X1 u1_u3_u0_U20 (.B1( u1_u3_u0_n125 ) , .ZN( u1_u3_u0_n126 ) , .A1( u1_u3_u0_n138 ) , .A2( u1_u3_u0_n146 ) , .B2( u1_u3_u0_n147 ) );
  NOR2_X1 u1_u3_u0_U21 (.A1( u1_u3_u0_n163 ) , .A2( u1_u3_u0_n164 ) , .ZN( u1_u3_u0_n95 ) );
  AOI22_X1 u1_u3_u0_U22 (.B2( u1_u3_u0_n109 ) , .A2( u1_u3_u0_n110 ) , .ZN( u1_u3_u0_n111 ) , .B1( u1_u3_u0_n118 ) , .A1( u1_u3_u0_n160 ) );
  NAND2_X1 u1_u3_u0_U23 (.A2( u1_u3_u0_n102 ) , .A1( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n149 ) );
  INV_X1 u1_u3_u0_U24 (.A( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n161 ) );
  INV_X1 u1_u3_u0_U25 (.A( u1_u3_u0_n118 ) , .ZN( u1_u3_u0_n158 ) );
  NAND2_X1 u1_u3_u0_U26 (.A2( u1_u3_u0_n100 ) , .ZN( u1_u3_u0_n131 ) , .A1( u1_u3_u0_n92 ) );
  NAND2_X1 u1_u3_u0_U27 (.ZN( u1_u3_u0_n108 ) , .A1( u1_u3_u0_n92 ) , .A2( u1_u3_u0_n94 ) );
  AOI21_X1 u1_u3_u0_U28 (.ZN( u1_u3_u0_n104 ) , .B1( u1_u3_u0_n107 ) , .B2( u1_u3_u0_n141 ) , .A( u1_u3_u0_n144 ) );
  AOI21_X1 u1_u3_u0_U29 (.B1( u1_u3_u0_n127 ) , .B2( u1_u3_u0_n129 ) , .A( u1_u3_u0_n138 ) , .ZN( u1_u3_u0_n96 ) );
  INV_X1 u1_u3_u0_U3 (.A( u1_u3_u0_n113 ) , .ZN( u1_u3_u0_n166 ) );
  NAND2_X1 u1_u3_u0_U30 (.A2( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n114 ) , .A1( u1_u3_u0_n92 ) );
  NOR2_X1 u1_u3_u0_U31 (.A1( u1_u3_u0_n120 ) , .ZN( u1_u3_u0_n143 ) , .A2( u1_u3_u0_n167 ) );
  OAI221_X1 u1_u3_u0_U32 (.C1( u1_u3_u0_n112 ) , .ZN( u1_u3_u0_n120 ) , .B1( u1_u3_u0_n138 ) , .B2( u1_u3_u0_n141 ) , .C2( u1_u3_u0_n147 ) , .A( u1_u3_u0_n172 ) );
  AOI211_X1 u1_u3_u0_U33 (.B( u1_u3_u0_n115 ) , .A( u1_u3_u0_n116 ) , .C2( u1_u3_u0_n117 ) , .C1( u1_u3_u0_n118 ) , .ZN( u1_u3_u0_n119 ) );
  NAND2_X1 u1_u3_u0_U34 (.A2( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n140 ) , .A1( u1_u3_u0_n94 ) );
  NAND2_X1 u1_u3_u0_U35 (.A1( u1_u3_u0_n100 ) , .A2( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n125 ) );
  NAND2_X1 u1_u3_u0_U36 (.A1( u1_u3_u0_n101 ) , .A2( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n150 ) );
  INV_X1 u1_u3_u0_U37 (.A( u1_u3_u0_n138 ) , .ZN( u1_u3_u0_n160 ) );
  NAND2_X1 u1_u3_u0_U38 (.A2( u1_u3_u0_n100 ) , .A1( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n139 ) );
  NAND2_X1 u1_u3_u0_U39 (.ZN( u1_u3_u0_n112 ) , .A2( u1_u3_u0_n92 ) , .A1( u1_u3_u0_n93 ) );
  AOI21_X1 u1_u3_u0_U4 (.B1( u1_u3_u0_n114 ) , .ZN( u1_u3_u0_n115 ) , .B2( u1_u3_u0_n129 ) , .A( u1_u3_u0_n161 ) );
  NAND2_X1 u1_u3_u0_U40 (.A1( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n130 ) , .A2( u1_u3_u0_n94 ) );
  INV_X1 u1_u3_u0_U41 (.ZN( u1_u3_u0_n172 ) , .A( u1_u3_u0_n88 ) );
  OAI222_X1 u1_u3_u0_U42 (.C1( u1_u3_u0_n108 ) , .A1( u1_u3_u0_n125 ) , .B2( u1_u3_u0_n128 ) , .B1( u1_u3_u0_n144 ) , .A2( u1_u3_u0_n158 ) , .C2( u1_u3_u0_n161 ) , .ZN( u1_u3_u0_n88 ) );
  NAND2_X1 u1_u3_u0_U43 (.A2( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n121 ) , .A1( u1_u3_u0_n93 ) );
  OR3_X1 u1_u3_u0_U44 (.A3( u1_u3_u0_n152 ) , .A2( u1_u3_u0_n153 ) , .A1( u1_u3_u0_n154 ) , .ZN( u1_u3_u0_n155 ) );
  AOI21_X1 u1_u3_u0_U45 (.A( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n145 ) , .B1( u1_u3_u0_n146 ) , .ZN( u1_u3_u0_n154 ) );
  AOI21_X1 u1_u3_u0_U46 (.B2( u1_u3_u0_n150 ) , .B1( u1_u3_u0_n151 ) , .ZN( u1_u3_u0_n152 ) , .A( u1_u3_u0_n158 ) );
  AOI21_X1 u1_u3_u0_U47 (.A( u1_u3_u0_n147 ) , .B2( u1_u3_u0_n148 ) , .B1( u1_u3_u0_n149 ) , .ZN( u1_u3_u0_n153 ) );
  INV_X1 u1_u3_u0_U48 (.ZN( u1_u3_u0_n171 ) , .A( u1_u3_u0_n99 ) );
  OAI211_X1 u1_u3_u0_U49 (.C2( u1_u3_u0_n140 ) , .C1( u1_u3_u0_n161 ) , .A( u1_u3_u0_n169 ) , .B( u1_u3_u0_n98 ) , .ZN( u1_u3_u0_n99 ) );
  AOI21_X1 u1_u3_u0_U5 (.B2( u1_u3_u0_n131 ) , .ZN( u1_u3_u0_n134 ) , .B1( u1_u3_u0_n151 ) , .A( u1_u3_u0_n158 ) );
  AOI211_X1 u1_u3_u0_U50 (.C1( u1_u3_u0_n118 ) , .A( u1_u3_u0_n123 ) , .B( u1_u3_u0_n96 ) , .C2( u1_u3_u0_n97 ) , .ZN( u1_u3_u0_n98 ) );
  INV_X1 u1_u3_u0_U51 (.ZN( u1_u3_u0_n169 ) , .A( u1_u3_u0_n91 ) );
  NOR2_X1 u1_u3_u0_U52 (.A2( u1_u3_X_4 ) , .A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n118 ) );
  NOR2_X1 u1_u3_u0_U53 (.A2( u1_u3_X_1 ) , .ZN( u1_u3_u0_n101 ) , .A1( u1_u3_u0_n163 ) );
  NOR2_X1 u1_u3_u0_U54 (.A2( u1_u3_X_3 ) , .A1( u1_u3_X_6 ) , .ZN( u1_u3_u0_n94 ) );
  NOR2_X1 u1_u3_u0_U55 (.A2( u1_u3_X_6 ) , .ZN( u1_u3_u0_n100 ) , .A1( u1_u3_u0_n162 ) );
  NAND2_X1 u1_u3_u0_U56 (.A2( u1_u3_X_4 ) , .A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n144 ) );
  NOR2_X1 u1_u3_u0_U57 (.A2( u1_u3_X_5 ) , .ZN( u1_u3_u0_n136 ) , .A1( u1_u3_u0_n159 ) );
  NAND2_X1 u1_u3_u0_U58 (.A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n138 ) , .A2( u1_u3_u0_n159 ) );
  AND2_X1 u1_u3_u0_U59 (.A2( u1_u3_X_3 ) , .A1( u1_u3_X_6 ) , .ZN( u1_u3_u0_n102 ) );
  NOR2_X1 u1_u3_u0_U6 (.A1( u1_u3_u0_n108 ) , .ZN( u1_u3_u0_n123 ) , .A2( u1_u3_u0_n158 ) );
  AND2_X1 u1_u3_u0_U60 (.A1( u1_u3_X_6 ) , .A2( u1_u3_u0_n162 ) , .ZN( u1_u3_u0_n93 ) );
  INV_X1 u1_u3_u0_U61 (.A( u1_u3_X_4 ) , .ZN( u1_u3_u0_n159 ) );
  INV_X1 u1_u3_u0_U62 (.A( u1_u3_X_1 ) , .ZN( u1_u3_u0_n164 ) );
  INV_X1 u1_u3_u0_U63 (.A( u1_u3_X_3 ) , .ZN( u1_u3_u0_n162 ) );
  INV_X1 u1_u3_u0_U64 (.A( u1_u3_u0_n126 ) , .ZN( u1_u3_u0_n168 ) );
  AOI211_X1 u1_u3_u0_U65 (.B( u1_u3_u0_n133 ) , .A( u1_u3_u0_n134 ) , .C2( u1_u3_u0_n135 ) , .C1( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n137 ) );
  OR4_X1 u1_u3_u0_U66 (.ZN( u1_out3_17 ) , .A4( u1_u3_u0_n122 ) , .A2( u1_u3_u0_n123 ) , .A1( u1_u3_u0_n124 ) , .A3( u1_u3_u0_n170 ) );
  AOI21_X1 u1_u3_u0_U67 (.B2( u1_u3_u0_n107 ) , .ZN( u1_u3_u0_n124 ) , .B1( u1_u3_u0_n128 ) , .A( u1_u3_u0_n161 ) );
  INV_X1 u1_u3_u0_U68 (.A( u1_u3_u0_n111 ) , .ZN( u1_u3_u0_n170 ) );
  OR4_X1 u1_u3_u0_U69 (.ZN( u1_out3_31 ) , .A4( u1_u3_u0_n155 ) , .A2( u1_u3_u0_n156 ) , .A1( u1_u3_u0_n157 ) , .A3( u1_u3_u0_n173 ) );
  OAI21_X1 u1_u3_u0_U7 (.B1( u1_u3_u0_n150 ) , .B2( u1_u3_u0_n158 ) , .A( u1_u3_u0_n172 ) , .ZN( u1_u3_u0_n89 ) );
  AOI21_X1 u1_u3_u0_U70 (.A( u1_u3_u0_n138 ) , .B2( u1_u3_u0_n139 ) , .B1( u1_u3_u0_n140 ) , .ZN( u1_u3_u0_n157 ) );
  INV_X1 u1_u3_u0_U71 (.ZN( u1_u3_u0_n174 ) , .A( u1_u3_u0_n89 ) );
  AOI211_X1 u1_u3_u0_U72 (.B( u1_u3_u0_n104 ) , .A( u1_u3_u0_n105 ) , .ZN( u1_u3_u0_n106 ) , .C2( u1_u3_u0_n113 ) , .C1( u1_u3_u0_n160 ) );
  AOI21_X1 u1_u3_u0_U73 (.B2( u1_u3_u0_n141 ) , .B1( u1_u3_u0_n142 ) , .ZN( u1_u3_u0_n156 ) , .A( u1_u3_u0_n161 ) );
  AOI21_X1 u1_u3_u0_U74 (.ZN( u1_u3_u0_n116 ) , .B2( u1_u3_u0_n142 ) , .A( u1_u3_u0_n144 ) , .B1( u1_u3_u0_n166 ) );
  INV_X1 u1_u3_u0_U75 (.A( u1_u3_u0_n142 ) , .ZN( u1_u3_u0_n165 ) );
  NOR2_X1 u1_u3_u0_U76 (.A2( u1_u3_X_1 ) , .A1( u1_u3_X_2 ) , .ZN( u1_u3_u0_n92 ) );
  NOR2_X1 u1_u3_u0_U77 (.A2( u1_u3_X_2 ) , .ZN( u1_u3_u0_n103 ) , .A1( u1_u3_u0_n164 ) );
  INV_X1 u1_u3_u0_U78 (.A( u1_u3_X_2 ) , .ZN( u1_u3_u0_n163 ) );
  OAI221_X1 u1_u3_u0_U79 (.C1( u1_u3_u0_n121 ) , .ZN( u1_u3_u0_n122 ) , .B2( u1_u3_u0_n127 ) , .A( u1_u3_u0_n143 ) , .B1( u1_u3_u0_n144 ) , .C2( u1_u3_u0_n147 ) );
  AND2_X1 u1_u3_u0_U8 (.A1( u1_u3_u0_n114 ) , .A2( u1_u3_u0_n121 ) , .ZN( u1_u3_u0_n146 ) );
  AOI21_X1 u1_u3_u0_U80 (.B1( u1_u3_u0_n132 ) , .ZN( u1_u3_u0_n133 ) , .A( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n166 ) );
  OAI22_X1 u1_u3_u0_U81 (.ZN( u1_u3_u0_n105 ) , .A2( u1_u3_u0_n132 ) , .B1( u1_u3_u0_n146 ) , .A1( u1_u3_u0_n147 ) , .B2( u1_u3_u0_n161 ) );
  NAND2_X1 u1_u3_u0_U82 (.ZN( u1_u3_u0_n110 ) , .A2( u1_u3_u0_n132 ) , .A1( u1_u3_u0_n145 ) );
  INV_X1 u1_u3_u0_U83 (.A( u1_u3_u0_n119 ) , .ZN( u1_u3_u0_n167 ) );
  NAND2_X1 u1_u3_u0_U84 (.ZN( u1_u3_u0_n148 ) , .A1( u1_u3_u0_n93 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U85 (.A1( u1_u3_u0_n100 ) , .ZN( u1_u3_u0_n129 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U86 (.A1( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n128 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U87 (.ZN( u1_u3_u0_n142 ) , .A1( u1_u3_u0_n94 ) , .A2( u1_u3_u0_n95 ) );
  NAND3_X1 u1_u3_u0_U88 (.ZN( u1_out3_23 ) , .A3( u1_u3_u0_n137 ) , .A1( u1_u3_u0_n168 ) , .A2( u1_u3_u0_n171 ) );
  NAND3_X1 u1_u3_u0_U89 (.A3( u1_u3_u0_n127 ) , .A2( u1_u3_u0_n128 ) , .ZN( u1_u3_u0_n135 ) , .A1( u1_u3_u0_n150 ) );
  NAND2_X1 u1_u3_u0_U9 (.ZN( u1_u3_u0_n113 ) , .A1( u1_u3_u0_n139 ) , .A2( u1_u3_u0_n149 ) );
  NAND3_X1 u1_u3_u0_U90 (.ZN( u1_u3_u0_n117 ) , .A3( u1_u3_u0_n132 ) , .A2( u1_u3_u0_n139 ) , .A1( u1_u3_u0_n148 ) );
  NAND3_X1 u1_u3_u0_U91 (.ZN( u1_u3_u0_n109 ) , .A2( u1_u3_u0_n114 ) , .A3( u1_u3_u0_n140 ) , .A1( u1_u3_u0_n149 ) );
  NAND3_X1 u1_u3_u0_U92 (.ZN( u1_out3_9 ) , .A3( u1_u3_u0_n106 ) , .A2( u1_u3_u0_n171 ) , .A1( u1_u3_u0_n174 ) );
  NAND3_X1 u1_u3_u0_U93 (.A2( u1_u3_u0_n128 ) , .A1( u1_u3_u0_n132 ) , .A3( u1_u3_u0_n146 ) , .ZN( u1_u3_u0_n97 ) );
  OAI22_X1 u1_u3_u2_U10 (.B1( u1_u3_u2_n151 ) , .A2( u1_u3_u2_n152 ) , .A1( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n160 ) , .B2( u1_u3_u2_n168 ) );
  NAND3_X1 u1_u3_u2_U100 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n104 ) , .A3( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n98 ) );
  NOR3_X1 u1_u3_u2_U11 (.A1( u1_u3_u2_n150 ) , .ZN( u1_u3_u2_n151 ) , .A3( u1_u3_u2_n175 ) , .A2( u1_u3_u2_n188 ) );
  AOI21_X1 u1_u3_u2_U12 (.B2( u1_u3_u2_n123 ) , .ZN( u1_u3_u2_n125 ) , .A( u1_u3_u2_n171 ) , .B1( u1_u3_u2_n184 ) );
  INV_X1 u1_u3_u2_U13 (.A( u1_u3_u2_n150 ) , .ZN( u1_u3_u2_n184 ) );
  AOI21_X1 u1_u3_u2_U14 (.ZN( u1_u3_u2_n144 ) , .B2( u1_u3_u2_n155 ) , .A( u1_u3_u2_n172 ) , .B1( u1_u3_u2_n185 ) );
  AOI21_X1 u1_u3_u2_U15 (.B2( u1_u3_u2_n143 ) , .ZN( u1_u3_u2_n145 ) , .B1( u1_u3_u2_n152 ) , .A( u1_u3_u2_n171 ) );
  INV_X1 u1_u3_u2_U16 (.A( u1_u3_u2_n156 ) , .ZN( u1_u3_u2_n171 ) );
  INV_X1 u1_u3_u2_U17 (.A( u1_u3_u2_n120 ) , .ZN( u1_u3_u2_n188 ) );
  NAND2_X1 u1_u3_u2_U18 (.A2( u1_u3_u2_n122 ) , .ZN( u1_u3_u2_n150 ) , .A1( u1_u3_u2_n152 ) );
  INV_X1 u1_u3_u2_U19 (.A( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n170 ) );
  INV_X1 u1_u3_u2_U20 (.A( u1_u3_u2_n137 ) , .ZN( u1_u3_u2_n173 ) );
  NAND2_X1 u1_u3_u2_U21 (.A1( u1_u3_u2_n132 ) , .A2( u1_u3_u2_n139 ) , .ZN( u1_u3_u2_n157 ) );
  INV_X1 u1_u3_u2_U22 (.A( u1_u3_u2_n113 ) , .ZN( u1_u3_u2_n178 ) );
  INV_X1 u1_u3_u2_U23 (.A( u1_u3_u2_n139 ) , .ZN( u1_u3_u2_n175 ) );
  INV_X1 u1_u3_u2_U24 (.A( u1_u3_u2_n155 ) , .ZN( u1_u3_u2_n181 ) );
  INV_X1 u1_u3_u2_U25 (.A( u1_u3_u2_n119 ) , .ZN( u1_u3_u2_n177 ) );
  INV_X1 u1_u3_u2_U26 (.A( u1_u3_u2_n116 ) , .ZN( u1_u3_u2_n180 ) );
  INV_X1 u1_u3_u2_U27 (.A( u1_u3_u2_n131 ) , .ZN( u1_u3_u2_n179 ) );
  INV_X1 u1_u3_u2_U28 (.A( u1_u3_u2_n154 ) , .ZN( u1_u3_u2_n176 ) );
  NAND2_X1 u1_u3_u2_U29 (.A2( u1_u3_u2_n116 ) , .A1( u1_u3_u2_n117 ) , .ZN( u1_u3_u2_n118 ) );
  NOR2_X1 u1_u3_u2_U3 (.ZN( u1_u3_u2_n121 ) , .A2( u1_u3_u2_n177 ) , .A1( u1_u3_u2_n180 ) );
  INV_X1 u1_u3_u2_U30 (.A( u1_u3_u2_n132 ) , .ZN( u1_u3_u2_n182 ) );
  INV_X1 u1_u3_u2_U31 (.A( u1_u3_u2_n158 ) , .ZN( u1_u3_u2_n183 ) );
  OAI21_X1 u1_u3_u2_U32 (.A( u1_u3_u2_n156 ) , .B1( u1_u3_u2_n157 ) , .ZN( u1_u3_u2_n158 ) , .B2( u1_u3_u2_n179 ) );
  NOR2_X1 u1_u3_u2_U33 (.ZN( u1_u3_u2_n156 ) , .A1( u1_u3_u2_n166 ) , .A2( u1_u3_u2_n169 ) );
  NOR2_X1 u1_u3_u2_U34 (.A2( u1_u3_u2_n114 ) , .ZN( u1_u3_u2_n137 ) , .A1( u1_u3_u2_n140 ) );
  NOR2_X1 u1_u3_u2_U35 (.A2( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n153 ) , .A1( u1_u3_u2_n156 ) );
  AOI211_X1 u1_u3_u2_U36 (.ZN( u1_u3_u2_n130 ) , .C1( u1_u3_u2_n138 ) , .C2( u1_u3_u2_n179 ) , .B( u1_u3_u2_n96 ) , .A( u1_u3_u2_n97 ) );
  OAI22_X1 u1_u3_u2_U37 (.B1( u1_u3_u2_n133 ) , .A2( u1_u3_u2_n137 ) , .A1( u1_u3_u2_n152 ) , .B2( u1_u3_u2_n168 ) , .ZN( u1_u3_u2_n97 ) );
  OAI221_X1 u1_u3_u2_U38 (.B1( u1_u3_u2_n113 ) , .C1( u1_u3_u2_n132 ) , .A( u1_u3_u2_n149 ) , .B2( u1_u3_u2_n171 ) , .C2( u1_u3_u2_n172 ) , .ZN( u1_u3_u2_n96 ) );
  OAI221_X1 u1_u3_u2_U39 (.A( u1_u3_u2_n115 ) , .C2( u1_u3_u2_n123 ) , .B2( u1_u3_u2_n143 ) , .B1( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n163 ) , .C1( u1_u3_u2_n168 ) );
  INV_X1 u1_u3_u2_U4 (.A( u1_u3_u2_n134 ) , .ZN( u1_u3_u2_n185 ) );
  OAI21_X1 u1_u3_u2_U40 (.A( u1_u3_u2_n114 ) , .ZN( u1_u3_u2_n115 ) , .B1( u1_u3_u2_n176 ) , .B2( u1_u3_u2_n178 ) );
  OAI221_X1 u1_u3_u2_U41 (.A( u1_u3_u2_n135 ) , .B2( u1_u3_u2_n136 ) , .B1( u1_u3_u2_n137 ) , .ZN( u1_u3_u2_n162 ) , .C2( u1_u3_u2_n167 ) , .C1( u1_u3_u2_n185 ) );
  AND3_X1 u1_u3_u2_U42 (.A3( u1_u3_u2_n131 ) , .A2( u1_u3_u2_n132 ) , .A1( u1_u3_u2_n133 ) , .ZN( u1_u3_u2_n136 ) );
  AOI22_X1 u1_u3_u2_U43 (.ZN( u1_u3_u2_n135 ) , .B1( u1_u3_u2_n140 ) , .A1( u1_u3_u2_n156 ) , .B2( u1_u3_u2_n180 ) , .A2( u1_u3_u2_n188 ) );
  AOI21_X1 u1_u3_u2_U44 (.ZN( u1_u3_u2_n149 ) , .B1( u1_u3_u2_n173 ) , .B2( u1_u3_u2_n188 ) , .A( u1_u3_u2_n95 ) );
  AND3_X1 u1_u3_u2_U45 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n104 ) , .A3( u1_u3_u2_n156 ) , .ZN( u1_u3_u2_n95 ) );
  OAI21_X1 u1_u3_u2_U46 (.A( u1_u3_u2_n101 ) , .B2( u1_u3_u2_n121 ) , .B1( u1_u3_u2_n153 ) , .ZN( u1_u3_u2_n164 ) );
  NAND2_X1 u1_u3_u2_U47 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n107 ) , .ZN( u1_u3_u2_n155 ) );
  NAND2_X1 u1_u3_u2_U48 (.A2( u1_u3_u2_n105 ) , .A1( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n143 ) );
  NAND2_X1 u1_u3_u2_U49 (.A1( u1_u3_u2_n104 ) , .A2( u1_u3_u2_n106 ) , .ZN( u1_u3_u2_n152 ) );
  NOR4_X1 u1_u3_u2_U5 (.A4( u1_u3_u2_n124 ) , .A3( u1_u3_u2_n125 ) , .A2( u1_u3_u2_n126 ) , .A1( u1_u3_u2_n127 ) , .ZN( u1_u3_u2_n128 ) );
  NAND2_X1 u1_u3_u2_U50 (.A1( u1_u3_u2_n100 ) , .A2( u1_u3_u2_n105 ) , .ZN( u1_u3_u2_n132 ) );
  INV_X1 u1_u3_u2_U51 (.A( u1_u3_u2_n140 ) , .ZN( u1_u3_u2_n168 ) );
  INV_X1 u1_u3_u2_U52 (.A( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n167 ) );
  OAI21_X1 u1_u3_u2_U53 (.A( u1_u3_u2_n141 ) , .B2( u1_u3_u2_n142 ) , .ZN( u1_u3_u2_n146 ) , .B1( u1_u3_u2_n153 ) );
  OAI21_X1 u1_u3_u2_U54 (.A( u1_u3_u2_n140 ) , .ZN( u1_u3_u2_n141 ) , .B1( u1_u3_u2_n176 ) , .B2( u1_u3_u2_n177 ) );
  NOR3_X1 u1_u3_u2_U55 (.ZN( u1_u3_u2_n142 ) , .A3( u1_u3_u2_n175 ) , .A2( u1_u3_u2_n178 ) , .A1( u1_u3_u2_n181 ) );
  INV_X1 u1_u3_u2_U56 (.ZN( u1_u3_u2_n187 ) , .A( u1_u3_u2_n99 ) );
  OAI21_X1 u1_u3_u2_U57 (.B1( u1_u3_u2_n137 ) , .B2( u1_u3_u2_n143 ) , .A( u1_u3_u2_n98 ) , .ZN( u1_u3_u2_n99 ) );
  NAND2_X1 u1_u3_u2_U58 (.A1( u1_u3_u2_n102 ) , .A2( u1_u3_u2_n106 ) , .ZN( u1_u3_u2_n113 ) );
  NAND2_X1 u1_u3_u2_U59 (.A1( u1_u3_u2_n106 ) , .A2( u1_u3_u2_n107 ) , .ZN( u1_u3_u2_n131 ) );
  AOI21_X1 u1_u3_u2_U6 (.B2( u1_u3_u2_n119 ) , .ZN( u1_u3_u2_n127 ) , .A( u1_u3_u2_n137 ) , .B1( u1_u3_u2_n155 ) );
  NAND2_X1 u1_u3_u2_U60 (.A1( u1_u3_u2_n103 ) , .A2( u1_u3_u2_n107 ) , .ZN( u1_u3_u2_n139 ) );
  NAND2_X1 u1_u3_u2_U61 (.A1( u1_u3_u2_n103 ) , .A2( u1_u3_u2_n105 ) , .ZN( u1_u3_u2_n133 ) );
  NAND2_X1 u1_u3_u2_U62 (.A1( u1_u3_u2_n102 ) , .A2( u1_u3_u2_n103 ) , .ZN( u1_u3_u2_n154 ) );
  NAND2_X1 u1_u3_u2_U63 (.A2( u1_u3_u2_n103 ) , .A1( u1_u3_u2_n104 ) , .ZN( u1_u3_u2_n119 ) );
  NAND2_X1 u1_u3_u2_U64 (.A2( u1_u3_u2_n107 ) , .A1( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n123 ) );
  NAND2_X1 u1_u3_u2_U65 (.A1( u1_u3_u2_n104 ) , .A2( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n122 ) );
  INV_X1 u1_u3_u2_U66 (.A( u1_u3_u2_n114 ) , .ZN( u1_u3_u2_n172 ) );
  NAND2_X1 u1_u3_u2_U67 (.A2( u1_u3_u2_n100 ) , .A1( u1_u3_u2_n102 ) , .ZN( u1_u3_u2_n116 ) );
  NAND2_X1 u1_u3_u2_U68 (.A1( u1_u3_u2_n102 ) , .A2( u1_u3_u2_n108 ) , .ZN( u1_u3_u2_n120 ) );
  NAND2_X1 u1_u3_u2_U69 (.A2( u1_u3_u2_n105 ) , .A1( u1_u3_u2_n106 ) , .ZN( u1_u3_u2_n117 ) );
  AOI21_X1 u1_u3_u2_U7 (.ZN( u1_u3_u2_n124 ) , .B1( u1_u3_u2_n131 ) , .B2( u1_u3_u2_n143 ) , .A( u1_u3_u2_n172 ) );
  NOR2_X1 u1_u3_u2_U70 (.A2( u1_u3_X_16 ) , .ZN( u1_u3_u2_n140 ) , .A1( u1_u3_u2_n166 ) );
  NOR2_X1 u1_u3_u2_U71 (.A2( u1_u3_X_13 ) , .A1( u1_u3_X_14 ) , .ZN( u1_u3_u2_n100 ) );
  NOR2_X1 u1_u3_u2_U72 (.A2( u1_u3_X_16 ) , .A1( u1_u3_X_17 ) , .ZN( u1_u3_u2_n138 ) );
  NOR2_X1 u1_u3_u2_U73 (.A2( u1_u3_X_15 ) , .A1( u1_u3_X_18 ) , .ZN( u1_u3_u2_n104 ) );
  NOR2_X1 u1_u3_u2_U74 (.A2( u1_u3_X_14 ) , .ZN( u1_u3_u2_n103 ) , .A1( u1_u3_u2_n174 ) );
  NOR2_X1 u1_u3_u2_U75 (.A2( u1_u3_X_15 ) , .ZN( u1_u3_u2_n102 ) , .A1( u1_u3_u2_n165 ) );
  NOR2_X1 u1_u3_u2_U76 (.A2( u1_u3_X_17 ) , .ZN( u1_u3_u2_n114 ) , .A1( u1_u3_u2_n169 ) );
  AND2_X1 u1_u3_u2_U77 (.A1( u1_u3_X_15 ) , .ZN( u1_u3_u2_n105 ) , .A2( u1_u3_u2_n165 ) );
  AND2_X1 u1_u3_u2_U78 (.A2( u1_u3_X_15 ) , .A1( u1_u3_X_18 ) , .ZN( u1_u3_u2_n107 ) );
  AND2_X1 u1_u3_u2_U79 (.A1( u1_u3_X_14 ) , .ZN( u1_u3_u2_n106 ) , .A2( u1_u3_u2_n174 ) );
  AOI21_X1 u1_u3_u2_U8 (.B2( u1_u3_u2_n120 ) , .B1( u1_u3_u2_n121 ) , .ZN( u1_u3_u2_n126 ) , .A( u1_u3_u2_n167 ) );
  AND2_X1 u1_u3_u2_U80 (.A1( u1_u3_X_13 ) , .A2( u1_u3_X_14 ) , .ZN( u1_u3_u2_n108 ) );
  INV_X1 u1_u3_u2_U81 (.A( u1_u3_X_16 ) , .ZN( u1_u3_u2_n169 ) );
  INV_X1 u1_u3_u2_U82 (.A( u1_u3_X_17 ) , .ZN( u1_u3_u2_n166 ) );
  INV_X1 u1_u3_u2_U83 (.A( u1_u3_X_13 ) , .ZN( u1_u3_u2_n174 ) );
  INV_X1 u1_u3_u2_U84 (.A( u1_u3_X_18 ) , .ZN( u1_u3_u2_n165 ) );
  NAND4_X1 u1_u3_u2_U85 (.ZN( u1_out3_30 ) , .A4( u1_u3_u2_n147 ) , .A3( u1_u3_u2_n148 ) , .A2( u1_u3_u2_n149 ) , .A1( u1_u3_u2_n187 ) );
  AOI21_X1 u1_u3_u2_U86 (.B2( u1_u3_u2_n138 ) , .ZN( u1_u3_u2_n148 ) , .A( u1_u3_u2_n162 ) , .B1( u1_u3_u2_n182 ) );
  NOR3_X1 u1_u3_u2_U87 (.A3( u1_u3_u2_n144 ) , .A2( u1_u3_u2_n145 ) , .A1( u1_u3_u2_n146 ) , .ZN( u1_u3_u2_n147 ) );
  NAND4_X1 u1_u3_u2_U88 (.ZN( u1_out3_24 ) , .A4( u1_u3_u2_n111 ) , .A3( u1_u3_u2_n112 ) , .A1( u1_u3_u2_n130 ) , .A2( u1_u3_u2_n187 ) );
  AOI221_X1 u1_u3_u2_U89 (.A( u1_u3_u2_n109 ) , .B1( u1_u3_u2_n110 ) , .ZN( u1_u3_u2_n111 ) , .C1( u1_u3_u2_n134 ) , .C2( u1_u3_u2_n170 ) , .B2( u1_u3_u2_n173 ) );
  OAI22_X1 u1_u3_u2_U9 (.ZN( u1_u3_u2_n109 ) , .A2( u1_u3_u2_n113 ) , .B2( u1_u3_u2_n133 ) , .B1( u1_u3_u2_n167 ) , .A1( u1_u3_u2_n168 ) );
  AOI21_X1 u1_u3_u2_U90 (.ZN( u1_u3_u2_n112 ) , .B2( u1_u3_u2_n156 ) , .A( u1_u3_u2_n164 ) , .B1( u1_u3_u2_n181 ) );
  NAND4_X1 u1_u3_u2_U91 (.ZN( u1_out3_16 ) , .A4( u1_u3_u2_n128 ) , .A3( u1_u3_u2_n129 ) , .A1( u1_u3_u2_n130 ) , .A2( u1_u3_u2_n186 ) );
  AOI22_X1 u1_u3_u2_U92 (.A2( u1_u3_u2_n118 ) , .ZN( u1_u3_u2_n129 ) , .A1( u1_u3_u2_n140 ) , .B1( u1_u3_u2_n157 ) , .B2( u1_u3_u2_n170 ) );
  INV_X1 u1_u3_u2_U93 (.A( u1_u3_u2_n163 ) , .ZN( u1_u3_u2_n186 ) );
  OR4_X1 u1_u3_u2_U94 (.ZN( u1_out3_6 ) , .A4( u1_u3_u2_n161 ) , .A3( u1_u3_u2_n162 ) , .A2( u1_u3_u2_n163 ) , .A1( u1_u3_u2_n164 ) );
  OR3_X1 u1_u3_u2_U95 (.A2( u1_u3_u2_n159 ) , .A1( u1_u3_u2_n160 ) , .ZN( u1_u3_u2_n161 ) , .A3( u1_u3_u2_n183 ) );
  AOI21_X1 u1_u3_u2_U96 (.B2( u1_u3_u2_n154 ) , .B1( u1_u3_u2_n155 ) , .ZN( u1_u3_u2_n159 ) , .A( u1_u3_u2_n167 ) );
  NAND3_X1 u1_u3_u2_U97 (.A2( u1_u3_u2_n117 ) , .A1( u1_u3_u2_n122 ) , .A3( u1_u3_u2_n123 ) , .ZN( u1_u3_u2_n134 ) );
  NAND3_X1 u1_u3_u2_U98 (.ZN( u1_u3_u2_n110 ) , .A2( u1_u3_u2_n131 ) , .A3( u1_u3_u2_n139 ) , .A1( u1_u3_u2_n154 ) );
  NAND3_X1 u1_u3_u2_U99 (.A2( u1_u3_u2_n100 ) , .ZN( u1_u3_u2_n101 ) , .A1( u1_u3_u2_n104 ) , .A3( u1_u3_u2_n114 ) );
  OAI22_X1 u1_u3_u3_U10 (.B1( u1_u3_u3_n113 ) , .A2( u1_u3_u3_n135 ) , .A1( u1_u3_u3_n150 ) , .B2( u1_u3_u3_n164 ) , .ZN( u1_u3_u3_n98 ) );
  OAI211_X1 u1_u3_u3_U11 (.B( u1_u3_u3_n106 ) , .ZN( u1_u3_u3_n119 ) , .C2( u1_u3_u3_n128 ) , .C1( u1_u3_u3_n167 ) , .A( u1_u3_u3_n181 ) );
  AOI221_X1 u1_u3_u3_U12 (.C1( u1_u3_u3_n105 ) , .ZN( u1_u3_u3_n106 ) , .A( u1_u3_u3_n131 ) , .B2( u1_u3_u3_n132 ) , .C2( u1_u3_u3_n133 ) , .B1( u1_u3_u3_n169 ) );
  INV_X1 u1_u3_u3_U13 (.ZN( u1_u3_u3_n181 ) , .A( u1_u3_u3_n98 ) );
  NAND2_X1 u1_u3_u3_U14 (.ZN( u1_u3_u3_n105 ) , .A2( u1_u3_u3_n130 ) , .A1( u1_u3_u3_n155 ) );
  AOI22_X1 u1_u3_u3_U15 (.B1( u1_u3_u3_n115 ) , .A2( u1_u3_u3_n116 ) , .ZN( u1_u3_u3_n123 ) , .B2( u1_u3_u3_n133 ) , .A1( u1_u3_u3_n169 ) );
  NAND2_X1 u1_u3_u3_U16 (.ZN( u1_u3_u3_n116 ) , .A2( u1_u3_u3_n151 ) , .A1( u1_u3_u3_n182 ) );
  NOR2_X1 u1_u3_u3_U17 (.ZN( u1_u3_u3_n126 ) , .A2( u1_u3_u3_n150 ) , .A1( u1_u3_u3_n164 ) );
  AOI21_X1 u1_u3_u3_U18 (.ZN( u1_u3_u3_n112 ) , .B2( u1_u3_u3_n146 ) , .B1( u1_u3_u3_n155 ) , .A( u1_u3_u3_n167 ) );
  NAND2_X1 u1_u3_u3_U19 (.A1( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n142 ) , .A2( u1_u3_u3_n164 ) );
  NAND2_X1 u1_u3_u3_U20 (.ZN( u1_u3_u3_n132 ) , .A2( u1_u3_u3_n152 ) , .A1( u1_u3_u3_n156 ) );
  INV_X1 u1_u3_u3_U21 (.A( u1_u3_u3_n133 ) , .ZN( u1_u3_u3_n165 ) );
  NAND2_X1 u1_u3_u3_U22 (.ZN( u1_u3_u3_n143 ) , .A1( u1_u3_u3_n165 ) , .A2( u1_u3_u3_n167 ) );
  AND2_X1 u1_u3_u3_U23 (.A2( u1_u3_u3_n113 ) , .A1( u1_u3_u3_n114 ) , .ZN( u1_u3_u3_n151 ) );
  INV_X1 u1_u3_u3_U24 (.A( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n170 ) );
  NAND2_X1 u1_u3_u3_U25 (.A1( u1_u3_u3_n107 ) , .A2( u1_u3_u3_n108 ) , .ZN( u1_u3_u3_n140 ) );
  NAND2_X1 u1_u3_u3_U26 (.ZN( u1_u3_u3_n117 ) , .A1( u1_u3_u3_n124 ) , .A2( u1_u3_u3_n148 ) );
  INV_X1 u1_u3_u3_U27 (.A( u1_u3_u3_n130 ) , .ZN( u1_u3_u3_n177 ) );
  INV_X1 u1_u3_u3_U28 (.A( u1_u3_u3_n128 ) , .ZN( u1_u3_u3_n176 ) );
  INV_X1 u1_u3_u3_U29 (.A( u1_u3_u3_n155 ) , .ZN( u1_u3_u3_n174 ) );
  INV_X1 u1_u3_u3_U3 (.A( u1_u3_u3_n140 ) , .ZN( u1_u3_u3_n182 ) );
  INV_X1 u1_u3_u3_U30 (.A( u1_u3_u3_n139 ) , .ZN( u1_u3_u3_n185 ) );
  NOR2_X1 u1_u3_u3_U31 (.ZN( u1_u3_u3_n135 ) , .A2( u1_u3_u3_n141 ) , .A1( u1_u3_u3_n169 ) );
  INV_X1 u1_u3_u3_U32 (.A( u1_u3_u3_n156 ) , .ZN( u1_u3_u3_n179 ) );
  OAI22_X1 u1_u3_u3_U33 (.B1( u1_u3_u3_n118 ) , .ZN( u1_u3_u3_n120 ) , .A1( u1_u3_u3_n135 ) , .B2( u1_u3_u3_n154 ) , .A2( u1_u3_u3_n178 ) );
  AND3_X1 u1_u3_u3_U34 (.ZN( u1_u3_u3_n118 ) , .A2( u1_u3_u3_n124 ) , .A1( u1_u3_u3_n144 ) , .A3( u1_u3_u3_n152 ) );
  OAI222_X1 u1_u3_u3_U35 (.C2( u1_u3_u3_n107 ) , .A2( u1_u3_u3_n108 ) , .B1( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n138 ) , .B2( u1_u3_u3_n146 ) , .C1( u1_u3_u3_n154 ) , .A1( u1_u3_u3_n164 ) );
  NOR4_X1 u1_u3_u3_U36 (.A4( u1_u3_u3_n157 ) , .A3( u1_u3_u3_n158 ) , .A2( u1_u3_u3_n159 ) , .A1( u1_u3_u3_n160 ) , .ZN( u1_u3_u3_n161 ) );
  AOI21_X1 u1_u3_u3_U37 (.B2( u1_u3_u3_n152 ) , .B1( u1_u3_u3_n153 ) , .ZN( u1_u3_u3_n158 ) , .A( u1_u3_u3_n164 ) );
  AOI21_X1 u1_u3_u3_U38 (.A( u1_u3_u3_n149 ) , .B2( u1_u3_u3_n150 ) , .B1( u1_u3_u3_n151 ) , .ZN( u1_u3_u3_n159 ) );
  AOI21_X1 u1_u3_u3_U39 (.A( u1_u3_u3_n154 ) , .B2( u1_u3_u3_n155 ) , .B1( u1_u3_u3_n156 ) , .ZN( u1_u3_u3_n157 ) );
  INV_X1 u1_u3_u3_U4 (.A( u1_u3_u3_n129 ) , .ZN( u1_u3_u3_n183 ) );
  AOI211_X1 u1_u3_u3_U40 (.ZN( u1_u3_u3_n109 ) , .A( u1_u3_u3_n119 ) , .C2( u1_u3_u3_n129 ) , .B( u1_u3_u3_n138 ) , .C1( u1_u3_u3_n141 ) );
  INV_X1 u1_u3_u3_U41 (.A( u1_u3_u3_n121 ) , .ZN( u1_u3_u3_n164 ) );
  NAND2_X1 u1_u3_u3_U42 (.ZN( u1_u3_u3_n133 ) , .A1( u1_u3_u3_n154 ) , .A2( u1_u3_u3_n164 ) );
  OAI211_X1 u1_u3_u3_U43 (.B( u1_u3_u3_n127 ) , .ZN( u1_u3_u3_n139 ) , .C1( u1_u3_u3_n150 ) , .C2( u1_u3_u3_n154 ) , .A( u1_u3_u3_n184 ) );
  INV_X1 u1_u3_u3_U44 (.A( u1_u3_u3_n125 ) , .ZN( u1_u3_u3_n184 ) );
  AOI221_X1 u1_u3_u3_U45 (.A( u1_u3_u3_n126 ) , .ZN( u1_u3_u3_n127 ) , .C2( u1_u3_u3_n132 ) , .C1( u1_u3_u3_n169 ) , .B2( u1_u3_u3_n170 ) , .B1( u1_u3_u3_n174 ) );
  OAI22_X1 u1_u3_u3_U46 (.A1( u1_u3_u3_n124 ) , .ZN( u1_u3_u3_n125 ) , .B2( u1_u3_u3_n145 ) , .A2( u1_u3_u3_n165 ) , .B1( u1_u3_u3_n167 ) );
  NOR2_X1 u1_u3_u3_U47 (.A1( u1_u3_u3_n113 ) , .ZN( u1_u3_u3_n131 ) , .A2( u1_u3_u3_n154 ) );
  NAND2_X1 u1_u3_u3_U48 (.A1( u1_u3_u3_n103 ) , .ZN( u1_u3_u3_n150 ) , .A2( u1_u3_u3_n99 ) );
  NAND2_X1 u1_u3_u3_U49 (.A2( u1_u3_u3_n102 ) , .ZN( u1_u3_u3_n155 ) , .A1( u1_u3_u3_n97 ) );
  INV_X1 u1_u3_u3_U5 (.A( u1_u3_u3_n117 ) , .ZN( u1_u3_u3_n178 ) );
  INV_X1 u1_u3_u3_U50 (.A( u1_u3_u3_n141 ) , .ZN( u1_u3_u3_n167 ) );
  AOI21_X1 u1_u3_u3_U51 (.B2( u1_u3_u3_n114 ) , .B1( u1_u3_u3_n146 ) , .A( u1_u3_u3_n154 ) , .ZN( u1_u3_u3_n94 ) );
  AOI21_X1 u1_u3_u3_U52 (.ZN( u1_u3_u3_n110 ) , .B2( u1_u3_u3_n142 ) , .B1( u1_u3_u3_n186 ) , .A( u1_u3_u3_n95 ) );
  INV_X1 u1_u3_u3_U53 (.A( u1_u3_u3_n145 ) , .ZN( u1_u3_u3_n186 ) );
  AOI21_X1 u1_u3_u3_U54 (.B1( u1_u3_u3_n124 ) , .A( u1_u3_u3_n149 ) , .B2( u1_u3_u3_n155 ) , .ZN( u1_u3_u3_n95 ) );
  INV_X1 u1_u3_u3_U55 (.A( u1_u3_u3_n149 ) , .ZN( u1_u3_u3_n169 ) );
  NAND2_X1 u1_u3_u3_U56 (.ZN( u1_u3_u3_n124 ) , .A1( u1_u3_u3_n96 ) , .A2( u1_u3_u3_n97 ) );
  NAND2_X1 u1_u3_u3_U57 (.A2( u1_u3_u3_n100 ) , .ZN( u1_u3_u3_n146 ) , .A1( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U58 (.A1( u1_u3_u3_n101 ) , .ZN( u1_u3_u3_n145 ) , .A2( u1_u3_u3_n99 ) );
  NAND2_X1 u1_u3_u3_U59 (.A1( u1_u3_u3_n100 ) , .ZN( u1_u3_u3_n156 ) , .A2( u1_u3_u3_n99 ) );
  AOI221_X1 u1_u3_u3_U6 (.A( u1_u3_u3_n131 ) , .C2( u1_u3_u3_n132 ) , .C1( u1_u3_u3_n133 ) , .ZN( u1_u3_u3_n134 ) , .B1( u1_u3_u3_n143 ) , .B2( u1_u3_u3_n177 ) );
  NAND2_X1 u1_u3_u3_U60 (.A2( u1_u3_u3_n101 ) , .A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n148 ) );
  NAND2_X1 u1_u3_u3_U61 (.A1( u1_u3_u3_n100 ) , .A2( u1_u3_u3_n102 ) , .ZN( u1_u3_u3_n128 ) );
  NAND2_X1 u1_u3_u3_U62 (.A2( u1_u3_u3_n101 ) , .A1( u1_u3_u3_n102 ) , .ZN( u1_u3_u3_n152 ) );
  NAND2_X1 u1_u3_u3_U63 (.A2( u1_u3_u3_n101 ) , .ZN( u1_u3_u3_n114 ) , .A1( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U64 (.ZN( u1_u3_u3_n107 ) , .A1( u1_u3_u3_n97 ) , .A2( u1_u3_u3_n99 ) );
  NAND2_X1 u1_u3_u3_U65 (.A2( u1_u3_u3_n100 ) , .A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n113 ) );
  NAND2_X1 u1_u3_u3_U66 (.A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n153 ) , .A2( u1_u3_u3_n97 ) );
  NAND2_X1 u1_u3_u3_U67 (.A2( u1_u3_u3_n103 ) , .A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n130 ) );
  NAND2_X1 u1_u3_u3_U68 (.A2( u1_u3_u3_n103 ) , .ZN( u1_u3_u3_n144 ) , .A1( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U69 (.A1( u1_u3_u3_n102 ) , .A2( u1_u3_u3_n103 ) , .ZN( u1_u3_u3_n108 ) );
  OAI22_X1 u1_u3_u3_U7 (.B2( u1_u3_u3_n147 ) , .A2( u1_u3_u3_n148 ) , .ZN( u1_u3_u3_n160 ) , .B1( u1_u3_u3_n165 ) , .A1( u1_u3_u3_n168 ) );
  NOR2_X1 u1_u3_u3_U70 (.A2( u1_u3_X_19 ) , .A1( u1_u3_X_20 ) , .ZN( u1_u3_u3_n99 ) );
  NOR2_X1 u1_u3_u3_U71 (.A2( u1_u3_X_21 ) , .A1( u1_u3_X_24 ) , .ZN( u1_u3_u3_n103 ) );
  NOR2_X1 u1_u3_u3_U72 (.A2( u1_u3_X_24 ) , .A1( u1_u3_u3_n171 ) , .ZN( u1_u3_u3_n97 ) );
  NOR2_X1 u1_u3_u3_U73 (.A2( u1_u3_X_19 ) , .A1( u1_u3_u3_n172 ) , .ZN( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U74 (.A1( u1_u3_X_22 ) , .A2( u1_u3_X_23 ) , .ZN( u1_u3_u3_n154 ) );
  AND2_X1 u1_u3_u3_U75 (.A1( u1_u3_X_24 ) , .ZN( u1_u3_u3_n101 ) , .A2( u1_u3_u3_n171 ) );
  AND2_X1 u1_u3_u3_U76 (.A1( u1_u3_X_19 ) , .ZN( u1_u3_u3_n102 ) , .A2( u1_u3_u3_n172 ) );
  AND2_X1 u1_u3_u3_U77 (.A1( u1_u3_X_21 ) , .A2( u1_u3_X_24 ) , .ZN( u1_u3_u3_n100 ) );
  AND2_X1 u1_u3_u3_U78 (.A2( u1_u3_X_19 ) , .A1( u1_u3_X_20 ) , .ZN( u1_u3_u3_n104 ) );
  INV_X1 u1_u3_u3_U79 (.A( u1_u3_X_21 ) , .ZN( u1_u3_u3_n171 ) );
  AND3_X1 u1_u3_u3_U8 (.A3( u1_u3_u3_n144 ) , .A2( u1_u3_u3_n145 ) , .A1( u1_u3_u3_n146 ) , .ZN( u1_u3_u3_n147 ) );
  INV_X1 u1_u3_u3_U80 (.A( u1_u3_X_20 ) , .ZN( u1_u3_u3_n172 ) );
  INV_X1 u1_u3_u3_U81 (.A( u1_u3_X_22 ) , .ZN( u1_u3_u3_n166 ) );
  NAND4_X1 u1_u3_u3_U82 (.ZN( u1_out3_26 ) , .A4( u1_u3_u3_n109 ) , .A3( u1_u3_u3_n110 ) , .A2( u1_u3_u3_n111 ) , .A1( u1_u3_u3_n173 ) );
  INV_X1 u1_u3_u3_U83 (.ZN( u1_u3_u3_n173 ) , .A( u1_u3_u3_n94 ) );
  OAI21_X1 u1_u3_u3_U84 (.ZN( u1_u3_u3_n111 ) , .B2( u1_u3_u3_n117 ) , .A( u1_u3_u3_n133 ) , .B1( u1_u3_u3_n176 ) );
  NAND4_X1 u1_u3_u3_U85 (.ZN( u1_out3_1 ) , .A4( u1_u3_u3_n161 ) , .A3( u1_u3_u3_n162 ) , .A2( u1_u3_u3_n163 ) , .A1( u1_u3_u3_n185 ) );
  NAND2_X1 u1_u3_u3_U86 (.ZN( u1_u3_u3_n163 ) , .A2( u1_u3_u3_n170 ) , .A1( u1_u3_u3_n176 ) );
  AOI22_X1 u1_u3_u3_U87 (.B2( u1_u3_u3_n140 ) , .B1( u1_u3_u3_n141 ) , .A2( u1_u3_u3_n142 ) , .ZN( u1_u3_u3_n162 ) , .A1( u1_u3_u3_n177 ) );
  NAND4_X1 u1_u3_u3_U88 (.ZN( u1_out3_20 ) , .A4( u1_u3_u3_n122 ) , .A3( u1_u3_u3_n123 ) , .A1( u1_u3_u3_n175 ) , .A2( u1_u3_u3_n180 ) );
  INV_X1 u1_u3_u3_U89 (.A( u1_u3_u3_n126 ) , .ZN( u1_u3_u3_n180 ) );
  INV_X1 u1_u3_u3_U9 (.A( u1_u3_u3_n143 ) , .ZN( u1_u3_u3_n168 ) );
  INV_X1 u1_u3_u3_U90 (.A( u1_u3_u3_n112 ) , .ZN( u1_u3_u3_n175 ) );
  OR4_X1 u1_u3_u3_U91 (.ZN( u1_out3_10 ) , .A4( u1_u3_u3_n136 ) , .A3( u1_u3_u3_n137 ) , .A1( u1_u3_u3_n138 ) , .A2( u1_u3_u3_n139 ) );
  OAI222_X1 u1_u3_u3_U92 (.C1( u1_u3_u3_n128 ) , .ZN( u1_u3_u3_n137 ) , .B1( u1_u3_u3_n148 ) , .A2( u1_u3_u3_n150 ) , .B2( u1_u3_u3_n154 ) , .C2( u1_u3_u3_n164 ) , .A1( u1_u3_u3_n167 ) );
  AOI211_X1 u1_u3_u3_U93 (.B( u1_u3_u3_n119 ) , .A( u1_u3_u3_n120 ) , .C2( u1_u3_u3_n121 ) , .ZN( u1_u3_u3_n122 ) , .C1( u1_u3_u3_n179 ) );
  OAI221_X1 u1_u3_u3_U94 (.A( u1_u3_u3_n134 ) , .B2( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n136 ) , .C1( u1_u3_u3_n149 ) , .B1( u1_u3_u3_n151 ) , .C2( u1_u3_u3_n183 ) );
  NOR2_X1 u1_u3_u3_U95 (.A2( u1_u3_X_23 ) , .ZN( u1_u3_u3_n141 ) , .A1( u1_u3_u3_n166 ) );
  NAND2_X1 u1_u3_u3_U96 (.A1( u1_u3_X_23 ) , .ZN( u1_u3_u3_n149 ) , .A2( u1_u3_u3_n166 ) );
  NOR2_X1 u1_u3_u3_U97 (.A2( u1_u3_X_22 ) , .A1( u1_u3_X_23 ) , .ZN( u1_u3_u3_n121 ) );
  NAND3_X1 u1_u3_u3_U98 (.A1( u1_u3_u3_n114 ) , .ZN( u1_u3_u3_n115 ) , .A2( u1_u3_u3_n145 ) , .A3( u1_u3_u3_n153 ) );
  NAND3_X1 u1_u3_u3_U99 (.ZN( u1_u3_u3_n129 ) , .A2( u1_u3_u3_n144 ) , .A1( u1_u3_u3_n153 ) , .A3( u1_u3_u3_n182 ) );
  AND3_X1 u1_u3_u7_U10 (.A3( u1_u3_u7_n110 ) , .A2( u1_u3_u7_n127 ) , .A1( u1_u3_u7_n132 ) , .ZN( u1_u3_u7_n92 ) );
  OAI21_X1 u1_u3_u7_U11 (.A( u1_u3_u7_n161 ) , .B1( u1_u3_u7_n168 ) , .B2( u1_u3_u7_n173 ) , .ZN( u1_u3_u7_n91 ) );
  AOI211_X1 u1_u3_u7_U12 (.A( u1_u3_u7_n117 ) , .ZN( u1_u3_u7_n118 ) , .C2( u1_u3_u7_n126 ) , .C1( u1_u3_u7_n177 ) , .B( u1_u3_u7_n180 ) );
  OAI22_X1 u1_u3_u7_U13 (.B1( u1_u3_u7_n115 ) , .ZN( u1_u3_u7_n117 ) , .A2( u1_u3_u7_n133 ) , .A1( u1_u3_u7_n137 ) , .B2( u1_u3_u7_n162 ) );
  INV_X1 u1_u3_u7_U14 (.A( u1_u3_u7_n116 ) , .ZN( u1_u3_u7_n180 ) );
  NOR3_X1 u1_u3_u7_U15 (.ZN( u1_u3_u7_n115 ) , .A3( u1_u3_u7_n145 ) , .A2( u1_u3_u7_n168 ) , .A1( u1_u3_u7_n169 ) );
  OAI211_X1 u1_u3_u7_U16 (.B( u1_u3_u7_n122 ) , .A( u1_u3_u7_n123 ) , .C2( u1_u3_u7_n124 ) , .ZN( u1_u3_u7_n154 ) , .C1( u1_u3_u7_n162 ) );
  AOI222_X1 u1_u3_u7_U17 (.ZN( u1_u3_u7_n122 ) , .C2( u1_u3_u7_n126 ) , .C1( u1_u3_u7_n145 ) , .B1( u1_u3_u7_n161 ) , .A2( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n170 ) , .A1( u1_u3_u7_n176 ) );
  INV_X1 u1_u3_u7_U18 (.A( u1_u3_u7_n133 ) , .ZN( u1_u3_u7_n176 ) );
  NOR3_X1 u1_u3_u7_U19 (.A2( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n135 ) , .ZN( u1_u3_u7_n136 ) , .A3( u1_u3_u7_n171 ) );
  NOR2_X1 u1_u3_u7_U20 (.A1( u1_u3_u7_n130 ) , .A2( u1_u3_u7_n134 ) , .ZN( u1_u3_u7_n153 ) );
  INV_X1 u1_u3_u7_U21 (.A( u1_u3_u7_n101 ) , .ZN( u1_u3_u7_n165 ) );
  NOR2_X1 u1_u3_u7_U22 (.ZN( u1_u3_u7_n111 ) , .A2( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n169 ) );
  AOI21_X1 u1_u3_u7_U23 (.ZN( u1_u3_u7_n104 ) , .B2( u1_u3_u7_n112 ) , .B1( u1_u3_u7_n127 ) , .A( u1_u3_u7_n164 ) );
  AOI21_X1 u1_u3_u7_U24 (.ZN( u1_u3_u7_n106 ) , .B1( u1_u3_u7_n133 ) , .B2( u1_u3_u7_n146 ) , .A( u1_u3_u7_n162 ) );
  AOI21_X1 u1_u3_u7_U25 (.A( u1_u3_u7_n101 ) , .ZN( u1_u3_u7_n107 ) , .B2( u1_u3_u7_n128 ) , .B1( u1_u3_u7_n175 ) );
  INV_X1 u1_u3_u7_U26 (.A( u1_u3_u7_n138 ) , .ZN( u1_u3_u7_n171 ) );
  INV_X1 u1_u3_u7_U27 (.A( u1_u3_u7_n131 ) , .ZN( u1_u3_u7_n177 ) );
  INV_X1 u1_u3_u7_U28 (.A( u1_u3_u7_n110 ) , .ZN( u1_u3_u7_n174 ) );
  NAND2_X1 u1_u3_u7_U29 (.A1( u1_u3_u7_n129 ) , .A2( u1_u3_u7_n132 ) , .ZN( u1_u3_u7_n149 ) );
  OAI21_X1 u1_u3_u7_U3 (.ZN( u1_u3_u7_n159 ) , .A( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n171 ) , .B1( u1_u3_u7_n174 ) );
  NAND2_X1 u1_u3_u7_U30 (.A1( u1_u3_u7_n113 ) , .A2( u1_u3_u7_n124 ) , .ZN( u1_u3_u7_n130 ) );
  INV_X1 u1_u3_u7_U31 (.A( u1_u3_u7_n112 ) , .ZN( u1_u3_u7_n173 ) );
  INV_X1 u1_u3_u7_U32 (.A( u1_u3_u7_n128 ) , .ZN( u1_u3_u7_n168 ) );
  INV_X1 u1_u3_u7_U33 (.A( u1_u3_u7_n148 ) , .ZN( u1_u3_u7_n169 ) );
  INV_X1 u1_u3_u7_U34 (.A( u1_u3_u7_n127 ) , .ZN( u1_u3_u7_n179 ) );
  NOR2_X1 u1_u3_u7_U35 (.ZN( u1_u3_u7_n101 ) , .A2( u1_u3_u7_n150 ) , .A1( u1_u3_u7_n156 ) );
  AOI211_X1 u1_u3_u7_U36 (.B( u1_u3_u7_n154 ) , .A( u1_u3_u7_n155 ) , .C1( u1_u3_u7_n156 ) , .ZN( u1_u3_u7_n157 ) , .C2( u1_u3_u7_n172 ) );
  INV_X1 u1_u3_u7_U37 (.A( u1_u3_u7_n153 ) , .ZN( u1_u3_u7_n172 ) );
  AOI211_X1 u1_u3_u7_U38 (.B( u1_u3_u7_n139 ) , .A( u1_u3_u7_n140 ) , .C2( u1_u3_u7_n141 ) , .ZN( u1_u3_u7_n142 ) , .C1( u1_u3_u7_n156 ) );
  NAND4_X1 u1_u3_u7_U39 (.A3( u1_u3_u7_n127 ) , .A2( u1_u3_u7_n128 ) , .A1( u1_u3_u7_n129 ) , .ZN( u1_u3_u7_n141 ) , .A4( u1_u3_u7_n147 ) );
  INV_X1 u1_u3_u7_U4 (.A( u1_u3_u7_n111 ) , .ZN( u1_u3_u7_n170 ) );
  AOI21_X1 u1_u3_u7_U40 (.A( u1_u3_u7_n137 ) , .B1( u1_u3_u7_n138 ) , .ZN( u1_u3_u7_n139 ) , .B2( u1_u3_u7_n146 ) );
  OAI22_X1 u1_u3_u7_U41 (.B1( u1_u3_u7_n136 ) , .ZN( u1_u3_u7_n140 ) , .A1( u1_u3_u7_n153 ) , .B2( u1_u3_u7_n162 ) , .A2( u1_u3_u7_n164 ) );
  AOI21_X1 u1_u3_u7_U42 (.ZN( u1_u3_u7_n123 ) , .B1( u1_u3_u7_n165 ) , .B2( u1_u3_u7_n177 ) , .A( u1_u3_u7_n97 ) );
  AOI21_X1 u1_u3_u7_U43 (.B2( u1_u3_u7_n113 ) , .B1( u1_u3_u7_n124 ) , .A( u1_u3_u7_n125 ) , .ZN( u1_u3_u7_n97 ) );
  INV_X1 u1_u3_u7_U44 (.A( u1_u3_u7_n125 ) , .ZN( u1_u3_u7_n161 ) );
  INV_X1 u1_u3_u7_U45 (.A( u1_u3_u7_n152 ) , .ZN( u1_u3_u7_n162 ) );
  AOI22_X1 u1_u3_u7_U46 (.A2( u1_u3_u7_n114 ) , .ZN( u1_u3_u7_n119 ) , .B1( u1_u3_u7_n130 ) , .A1( u1_u3_u7_n156 ) , .B2( u1_u3_u7_n165 ) );
  NAND2_X1 u1_u3_u7_U47 (.A2( u1_u3_u7_n112 ) , .ZN( u1_u3_u7_n114 ) , .A1( u1_u3_u7_n175 ) );
  AND2_X1 u1_u3_u7_U48 (.ZN( u1_u3_u7_n145 ) , .A2( u1_u3_u7_n98 ) , .A1( u1_u3_u7_n99 ) );
  NOR2_X1 u1_u3_u7_U49 (.ZN( u1_u3_u7_n137 ) , .A1( u1_u3_u7_n150 ) , .A2( u1_u3_u7_n161 ) );
  INV_X1 u1_u3_u7_U5 (.A( u1_u3_u7_n149 ) , .ZN( u1_u3_u7_n175 ) );
  AOI21_X1 u1_u3_u7_U50 (.ZN( u1_u3_u7_n105 ) , .B2( u1_u3_u7_n110 ) , .A( u1_u3_u7_n125 ) , .B1( u1_u3_u7_n147 ) );
  NAND2_X1 u1_u3_u7_U51 (.ZN( u1_u3_u7_n146 ) , .A1( u1_u3_u7_n95 ) , .A2( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U52 (.A2( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n147 ) , .A1( u1_u3_u7_n93 ) );
  NAND2_X1 u1_u3_u7_U53 (.A1( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n127 ) , .A2( u1_u3_u7_n99 ) );
  OR2_X1 u1_u3_u7_U54 (.ZN( u1_u3_u7_n126 ) , .A2( u1_u3_u7_n152 ) , .A1( u1_u3_u7_n156 ) );
  NAND2_X1 u1_u3_u7_U55 (.A2( u1_u3_u7_n102 ) , .A1( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n133 ) );
  NAND2_X1 u1_u3_u7_U56 (.ZN( u1_u3_u7_n112 ) , .A2( u1_u3_u7_n96 ) , .A1( u1_u3_u7_n99 ) );
  NAND2_X1 u1_u3_u7_U57 (.A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n128 ) , .A1( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U58 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n113 ) , .A2( u1_u3_u7_n93 ) );
  NAND2_X1 u1_u3_u7_U59 (.A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n124 ) , .A1( u1_u3_u7_n96 ) );
  INV_X1 u1_u3_u7_U6 (.A( u1_u3_u7_n154 ) , .ZN( u1_u3_u7_n178 ) );
  NAND2_X1 u1_u3_u7_U60 (.ZN( u1_u3_u7_n110 ) , .A1( u1_u3_u7_n95 ) , .A2( u1_u3_u7_n96 ) );
  INV_X1 u1_u3_u7_U61 (.A( u1_u3_u7_n150 ) , .ZN( u1_u3_u7_n164 ) );
  AND2_X1 u1_u3_u7_U62 (.ZN( u1_u3_u7_n134 ) , .A1( u1_u3_u7_n93 ) , .A2( u1_u3_u7_n98 ) );
  NAND2_X1 u1_u3_u7_U63 (.A1( u1_u3_u7_n100 ) , .A2( u1_u3_u7_n102 ) , .ZN( u1_u3_u7_n129 ) );
  NAND2_X1 u1_u3_u7_U64 (.A2( u1_u3_u7_n103 ) , .ZN( u1_u3_u7_n131 ) , .A1( u1_u3_u7_n95 ) );
  NAND2_X1 u1_u3_u7_U65 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n138 ) , .A2( u1_u3_u7_n99 ) );
  NAND2_X1 u1_u3_u7_U66 (.ZN( u1_u3_u7_n132 ) , .A1( u1_u3_u7_n93 ) , .A2( u1_u3_u7_n96 ) );
  NAND2_X1 u1_u3_u7_U67 (.A1( u1_u3_u7_n100 ) , .ZN( u1_u3_u7_n148 ) , .A2( u1_u3_u7_n95 ) );
  NOR2_X1 u1_u3_u7_U68 (.A2( u1_u3_X_47 ) , .ZN( u1_u3_u7_n150 ) , .A1( u1_u3_u7_n163 ) );
  NOR2_X1 u1_u3_u7_U69 (.A2( u1_u3_X_43 ) , .A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n103 ) );
  AOI211_X1 u1_u3_u7_U7 (.ZN( u1_u3_u7_n116 ) , .A( u1_u3_u7_n155 ) , .C1( u1_u3_u7_n161 ) , .C2( u1_u3_u7_n171 ) , .B( u1_u3_u7_n94 ) );
  NOR2_X1 u1_u3_u7_U70 (.A2( u1_u3_X_48 ) , .A1( u1_u3_u7_n166 ) , .ZN( u1_u3_u7_n95 ) );
  NOR2_X1 u1_u3_u7_U71 (.A2( u1_u3_X_45 ) , .A1( u1_u3_X_48 ) , .ZN( u1_u3_u7_n99 ) );
  NOR2_X1 u1_u3_u7_U72 (.A2( u1_u3_X_44 ) , .A1( u1_u3_u7_n167 ) , .ZN( u1_u3_u7_n98 ) );
  NOR2_X1 u1_u3_u7_U73 (.A2( u1_u3_X_46 ) , .A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n152 ) );
  AND2_X1 u1_u3_u7_U74 (.A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n156 ) , .A2( u1_u3_u7_n163 ) );
  NAND2_X1 u1_u3_u7_U75 (.A2( u1_u3_X_46 ) , .A1( u1_u3_X_47 ) , .ZN( u1_u3_u7_n125 ) );
  AND2_X1 u1_u3_u7_U76 (.A2( u1_u3_X_45 ) , .A1( u1_u3_X_48 ) , .ZN( u1_u3_u7_n102 ) );
  AND2_X1 u1_u3_u7_U77 (.A2( u1_u3_X_43 ) , .A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n96 ) );
  AND2_X1 u1_u3_u7_U78 (.A1( u1_u3_X_44 ) , .ZN( u1_u3_u7_n100 ) , .A2( u1_u3_u7_n167 ) );
  AND2_X1 u1_u3_u7_U79 (.A1( u1_u3_X_48 ) , .A2( u1_u3_u7_n166 ) , .ZN( u1_u3_u7_n93 ) );
  OAI222_X1 u1_u3_u7_U8 (.C2( u1_u3_u7_n101 ) , .B2( u1_u3_u7_n111 ) , .A1( u1_u3_u7_n113 ) , .C1( u1_u3_u7_n146 ) , .A2( u1_u3_u7_n162 ) , .B1( u1_u3_u7_n164 ) , .ZN( u1_u3_u7_n94 ) );
  INV_X1 u1_u3_u7_U80 (.A( u1_u3_X_46 ) , .ZN( u1_u3_u7_n163 ) );
  INV_X1 u1_u3_u7_U81 (.A( u1_u3_X_43 ) , .ZN( u1_u3_u7_n167 ) );
  INV_X1 u1_u3_u7_U82 (.A( u1_u3_X_45 ) , .ZN( u1_u3_u7_n166 ) );
  NAND4_X1 u1_u3_u7_U83 (.ZN( u1_out3_5 ) , .A4( u1_u3_u7_n108 ) , .A3( u1_u3_u7_n109 ) , .A1( u1_u3_u7_n116 ) , .A2( u1_u3_u7_n123 ) );
  AOI22_X1 u1_u3_u7_U84 (.ZN( u1_u3_u7_n109 ) , .A2( u1_u3_u7_n126 ) , .B2( u1_u3_u7_n145 ) , .B1( u1_u3_u7_n156 ) , .A1( u1_u3_u7_n171 ) );
  NOR4_X1 u1_u3_u7_U85 (.A4( u1_u3_u7_n104 ) , .A3( u1_u3_u7_n105 ) , .A2( u1_u3_u7_n106 ) , .A1( u1_u3_u7_n107 ) , .ZN( u1_u3_u7_n108 ) );
  NAND4_X1 u1_u3_u7_U86 (.ZN( u1_out3_27 ) , .A4( u1_u3_u7_n118 ) , .A3( u1_u3_u7_n119 ) , .A2( u1_u3_u7_n120 ) , .A1( u1_u3_u7_n121 ) );
  OAI21_X1 u1_u3_u7_U87 (.ZN( u1_u3_u7_n121 ) , .B2( u1_u3_u7_n145 ) , .A( u1_u3_u7_n150 ) , .B1( u1_u3_u7_n174 ) );
  OAI21_X1 u1_u3_u7_U88 (.ZN( u1_u3_u7_n120 ) , .A( u1_u3_u7_n161 ) , .B2( u1_u3_u7_n170 ) , .B1( u1_u3_u7_n179 ) );
  NAND4_X1 u1_u3_u7_U89 (.ZN( u1_out3_21 ) , .A4( u1_u3_u7_n157 ) , .A3( u1_u3_u7_n158 ) , .A2( u1_u3_u7_n159 ) , .A1( u1_u3_u7_n160 ) );
  OAI221_X1 u1_u3_u7_U9 (.C1( u1_u3_u7_n101 ) , .C2( u1_u3_u7_n147 ) , .ZN( u1_u3_u7_n155 ) , .B2( u1_u3_u7_n162 ) , .A( u1_u3_u7_n91 ) , .B1( u1_u3_u7_n92 ) );
  OAI21_X1 u1_u3_u7_U90 (.B1( u1_u3_u7_n145 ) , .ZN( u1_u3_u7_n160 ) , .A( u1_u3_u7_n161 ) , .B2( u1_u3_u7_n177 ) );
  AOI22_X1 u1_u3_u7_U91 (.B2( u1_u3_u7_n149 ) , .B1( u1_u3_u7_n150 ) , .A2( u1_u3_u7_n151 ) , .A1( u1_u3_u7_n152 ) , .ZN( u1_u3_u7_n158 ) );
  NAND4_X1 u1_u3_u7_U92 (.ZN( u1_out3_15 ) , .A4( u1_u3_u7_n142 ) , .A3( u1_u3_u7_n143 ) , .A2( u1_u3_u7_n144 ) , .A1( u1_u3_u7_n178 ) );
  OR2_X1 u1_u3_u7_U93 (.A2( u1_u3_u7_n125 ) , .A1( u1_u3_u7_n129 ) , .ZN( u1_u3_u7_n144 ) );
  AOI22_X1 u1_u3_u7_U94 (.A2( u1_u3_u7_n126 ) , .ZN( u1_u3_u7_n143 ) , .B2( u1_u3_u7_n165 ) , .B1( u1_u3_u7_n173 ) , .A1( u1_u3_u7_n174 ) );
  NAND3_X1 u1_u3_u7_U95 (.A3( u1_u3_u7_n146 ) , .A2( u1_u3_u7_n147 ) , .A1( u1_u3_u7_n148 ) , .ZN( u1_u3_u7_n151 ) );
  NAND3_X1 u1_u3_u7_U96 (.A3( u1_u3_u7_n131 ) , .A2( u1_u3_u7_n132 ) , .A1( u1_u3_u7_n133 ) , .ZN( u1_u3_u7_n135 ) );
  XOR2_X1 u1_u7_U10 (.B( u1_K8_45 ) , .A( u1_R6_30 ) , .Z( u1_u7_X_45 ) );
  XOR2_X1 u1_u7_U11 (.B( u1_K8_44 ) , .A( u1_R6_29 ) , .Z( u1_u7_X_44 ) );
  XOR2_X1 u1_u7_U12 (.B( u1_K8_43 ) , .A( u1_R6_28 ) , .Z( u1_u7_X_43 ) );
  XOR2_X1 u1_u7_U7 (.B( u1_K8_48 ) , .A( u1_R6_1 ) , .Z( u1_u7_X_48 ) );
  XOR2_X1 u1_u7_U8 (.B( u1_K8_47 ) , .A( u1_R6_32 ) , .Z( u1_u7_X_47 ) );
  XOR2_X1 u1_u7_U9 (.B( u1_K8_46 ) , .A( u1_R6_31 ) , .Z( u1_u7_X_46 ) );
  OAI221_X1 u1_u7_u7_U10 (.C1( u1_u7_u7_n101 ) , .C2( u1_u7_u7_n147 ) , .ZN( u1_u7_u7_n155 ) , .B2( u1_u7_u7_n162 ) , .A( u1_u7_u7_n91 ) , .B1( u1_u7_u7_n92 ) );
  AND3_X1 u1_u7_u7_U11 (.A3( u1_u7_u7_n110 ) , .A2( u1_u7_u7_n127 ) , .A1( u1_u7_u7_n132 ) , .ZN( u1_u7_u7_n92 ) );
  OAI21_X1 u1_u7_u7_U12 (.A( u1_u7_u7_n161 ) , .B1( u1_u7_u7_n168 ) , .B2( u1_u7_u7_n173 ) , .ZN( u1_u7_u7_n91 ) );
  AOI211_X1 u1_u7_u7_U13 (.A( u1_u7_u7_n117 ) , .ZN( u1_u7_u7_n118 ) , .C2( u1_u7_u7_n126 ) , .C1( u1_u7_u7_n177 ) , .B( u1_u7_u7_n180 ) );
  OAI22_X1 u1_u7_u7_U14 (.B1( u1_u7_u7_n115 ) , .ZN( u1_u7_u7_n117 ) , .A2( u1_u7_u7_n133 ) , .A1( u1_u7_u7_n137 ) , .B2( u1_u7_u7_n162 ) );
  INV_X1 u1_u7_u7_U15 (.A( u1_u7_u7_n116 ) , .ZN( u1_u7_u7_n180 ) );
  NOR3_X1 u1_u7_u7_U16 (.ZN( u1_u7_u7_n115 ) , .A3( u1_u7_u7_n145 ) , .A2( u1_u7_u7_n168 ) , .A1( u1_u7_u7_n169 ) );
  NOR3_X1 u1_u7_u7_U17 (.A2( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n135 ) , .ZN( u1_u7_u7_n136 ) , .A3( u1_u7_u7_n171 ) );
  NOR2_X1 u1_u7_u7_U18 (.A1( u1_u7_u7_n130 ) , .A2( u1_u7_u7_n134 ) , .ZN( u1_u7_u7_n153 ) );
  NOR2_X1 u1_u7_u7_U19 (.ZN( u1_u7_u7_n111 ) , .A2( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n169 ) );
  AOI21_X1 u1_u7_u7_U20 (.ZN( u1_u7_u7_n104 ) , .B2( u1_u7_u7_n112 ) , .B1( u1_u7_u7_n127 ) , .A( u1_u7_u7_n164 ) );
  AOI21_X1 u1_u7_u7_U21 (.ZN( u1_u7_u7_n106 ) , .B1( u1_u7_u7_n133 ) , .B2( u1_u7_u7_n146 ) , .A( u1_u7_u7_n162 ) );
  AOI21_X1 u1_u7_u7_U22 (.A( u1_u7_u7_n101 ) , .ZN( u1_u7_u7_n107 ) , .B2( u1_u7_u7_n128 ) , .B1( u1_u7_u7_n175 ) );
  INV_X1 u1_u7_u7_U23 (.A( u1_u7_u7_n101 ) , .ZN( u1_u7_u7_n165 ) );
  INV_X1 u1_u7_u7_U24 (.A( u1_u7_u7_n138 ) , .ZN( u1_u7_u7_n171 ) );
  INV_X1 u1_u7_u7_U25 (.A( u1_u7_u7_n131 ) , .ZN( u1_u7_u7_n177 ) );
  INV_X1 u1_u7_u7_U26 (.A( u1_u7_u7_n110 ) , .ZN( u1_u7_u7_n174 ) );
  NAND2_X1 u1_u7_u7_U27 (.A1( u1_u7_u7_n129 ) , .A2( u1_u7_u7_n132 ) , .ZN( u1_u7_u7_n149 ) );
  NAND2_X1 u1_u7_u7_U28 (.A1( u1_u7_u7_n113 ) , .A2( u1_u7_u7_n124 ) , .ZN( u1_u7_u7_n130 ) );
  INV_X1 u1_u7_u7_U29 (.A( u1_u7_u7_n128 ) , .ZN( u1_u7_u7_n168 ) );
  OAI21_X1 u1_u7_u7_U3 (.ZN( u1_u7_u7_n159 ) , .A( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n171 ) , .B1( u1_u7_u7_n174 ) );
  INV_X1 u1_u7_u7_U30 (.A( u1_u7_u7_n148 ) , .ZN( u1_u7_u7_n169 ) );
  INV_X1 u1_u7_u7_U31 (.A( u1_u7_u7_n112 ) , .ZN( u1_u7_u7_n173 ) );
  INV_X1 u1_u7_u7_U32 (.A( u1_u7_u7_n127 ) , .ZN( u1_u7_u7_n179 ) );
  NOR2_X1 u1_u7_u7_U33 (.ZN( u1_u7_u7_n101 ) , .A2( u1_u7_u7_n150 ) , .A1( u1_u7_u7_n156 ) );
  AOI211_X1 u1_u7_u7_U34 (.B( u1_u7_u7_n154 ) , .A( u1_u7_u7_n155 ) , .C1( u1_u7_u7_n156 ) , .ZN( u1_u7_u7_n157 ) , .C2( u1_u7_u7_n172 ) );
  INV_X1 u1_u7_u7_U35 (.A( u1_u7_u7_n153 ) , .ZN( u1_u7_u7_n172 ) );
  AOI211_X1 u1_u7_u7_U36 (.B( u1_u7_u7_n139 ) , .A( u1_u7_u7_n140 ) , .C2( u1_u7_u7_n141 ) , .ZN( u1_u7_u7_n142 ) , .C1( u1_u7_u7_n156 ) );
  NAND4_X1 u1_u7_u7_U37 (.A3( u1_u7_u7_n127 ) , .A2( u1_u7_u7_n128 ) , .A1( u1_u7_u7_n129 ) , .ZN( u1_u7_u7_n141 ) , .A4( u1_u7_u7_n147 ) );
  AOI21_X1 u1_u7_u7_U38 (.A( u1_u7_u7_n137 ) , .B1( u1_u7_u7_n138 ) , .ZN( u1_u7_u7_n139 ) , .B2( u1_u7_u7_n146 ) );
  OAI22_X1 u1_u7_u7_U39 (.B1( u1_u7_u7_n136 ) , .ZN( u1_u7_u7_n140 ) , .A1( u1_u7_u7_n153 ) , .B2( u1_u7_u7_n162 ) , .A2( u1_u7_u7_n164 ) );
  INV_X1 u1_u7_u7_U4 (.A( u1_u7_u7_n149 ) , .ZN( u1_u7_u7_n175 ) );
  INV_X1 u1_u7_u7_U40 (.A( u1_u7_u7_n125 ) , .ZN( u1_u7_u7_n161 ) );
  AOI21_X1 u1_u7_u7_U41 (.ZN( u1_u7_u7_n123 ) , .B1( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n177 ) , .A( u1_u7_u7_n97 ) );
  AOI21_X1 u1_u7_u7_U42 (.B2( u1_u7_u7_n113 ) , .B1( u1_u7_u7_n124 ) , .A( u1_u7_u7_n125 ) , .ZN( u1_u7_u7_n97 ) );
  INV_X1 u1_u7_u7_U43 (.A( u1_u7_u7_n152 ) , .ZN( u1_u7_u7_n162 ) );
  AOI22_X1 u1_u7_u7_U44 (.A2( u1_u7_u7_n114 ) , .ZN( u1_u7_u7_n119 ) , .B1( u1_u7_u7_n130 ) , .A1( u1_u7_u7_n156 ) , .B2( u1_u7_u7_n165 ) );
  NAND2_X1 u1_u7_u7_U45 (.A2( u1_u7_u7_n112 ) , .ZN( u1_u7_u7_n114 ) , .A1( u1_u7_u7_n175 ) );
  NOR2_X1 u1_u7_u7_U46 (.ZN( u1_u7_u7_n137 ) , .A1( u1_u7_u7_n150 ) , .A2( u1_u7_u7_n161 ) );
  AND2_X1 u1_u7_u7_U47 (.ZN( u1_u7_u7_n145 ) , .A2( u1_u7_u7_n98 ) , .A1( u1_u7_u7_n99 ) );
  AOI21_X1 u1_u7_u7_U48 (.ZN( u1_u7_u7_n105 ) , .B2( u1_u7_u7_n110 ) , .A( u1_u7_u7_n125 ) , .B1( u1_u7_u7_n147 ) );
  NAND2_X1 u1_u7_u7_U49 (.ZN( u1_u7_u7_n146 ) , .A1( u1_u7_u7_n95 ) , .A2( u1_u7_u7_n98 ) );
  INV_X1 u1_u7_u7_U5 (.A( u1_u7_u7_n154 ) , .ZN( u1_u7_u7_n178 ) );
  NAND2_X1 u1_u7_u7_U50 (.A2( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n147 ) , .A1( u1_u7_u7_n93 ) );
  NAND2_X1 u1_u7_u7_U51 (.A1( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n127 ) , .A2( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U52 (.A2( u1_u7_u7_n102 ) , .A1( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n133 ) );
  OR2_X1 u1_u7_u7_U53 (.ZN( u1_u7_u7_n126 ) , .A2( u1_u7_u7_n152 ) , .A1( u1_u7_u7_n156 ) );
  NAND2_X1 u1_u7_u7_U54 (.ZN( u1_u7_u7_n112 ) , .A2( u1_u7_u7_n96 ) , .A1( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U55 (.A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n128 ) , .A1( u1_u7_u7_n98 ) );
  INV_X1 u1_u7_u7_U56 (.A( u1_u7_u7_n150 ) , .ZN( u1_u7_u7_n164 ) );
  AND2_X1 u1_u7_u7_U57 (.ZN( u1_u7_u7_n134 ) , .A1( u1_u7_u7_n93 ) , .A2( u1_u7_u7_n98 ) );
  NAND2_X1 u1_u7_u7_U58 (.ZN( u1_u7_u7_n110 ) , .A1( u1_u7_u7_n95 ) , .A2( u1_u7_u7_n96 ) );
  NAND2_X1 u1_u7_u7_U59 (.A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n124 ) , .A1( u1_u7_u7_n96 ) );
  INV_X1 u1_u7_u7_U6 (.A( u1_u7_u7_n111 ) , .ZN( u1_u7_u7_n170 ) );
  NAND2_X1 u1_u7_u7_U60 (.ZN( u1_u7_u7_n132 ) , .A1( u1_u7_u7_n93 ) , .A2( u1_u7_u7_n96 ) );
  NAND2_X1 u1_u7_u7_U61 (.A2( u1_u7_u7_n103 ) , .ZN( u1_u7_u7_n131 ) , .A1( u1_u7_u7_n95 ) );
  NOR2_X1 u1_u7_u7_U62 (.A2( u1_u7_X_47 ) , .ZN( u1_u7_u7_n150 ) , .A1( u1_u7_u7_n163 ) );
  NOR2_X1 u1_u7_u7_U63 (.A2( u1_u7_X_43 ) , .A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n103 ) );
  NOR2_X1 u1_u7_u7_U64 (.A2( u1_u7_X_48 ) , .A1( u1_u7_u7_n166 ) , .ZN( u1_u7_u7_n95 ) );
  NOR2_X1 u1_u7_u7_U65 (.A2( u1_u7_X_44 ) , .A1( u1_u7_u7_n167 ) , .ZN( u1_u7_u7_n98 ) );
  NOR2_X1 u1_u7_u7_U66 (.A2( u1_u7_X_45 ) , .A1( u1_u7_X_48 ) , .ZN( u1_u7_u7_n99 ) );
  NOR2_X1 u1_u7_u7_U67 (.A2( u1_u7_X_46 ) , .A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n152 ) );
  AND2_X1 u1_u7_u7_U68 (.A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n156 ) , .A2( u1_u7_u7_n163 ) );
  NAND2_X1 u1_u7_u7_U69 (.A2( u1_u7_X_46 ) , .A1( u1_u7_X_47 ) , .ZN( u1_u7_u7_n125 ) );
  AOI211_X1 u1_u7_u7_U7 (.ZN( u1_u7_u7_n116 ) , .A( u1_u7_u7_n155 ) , .C1( u1_u7_u7_n161 ) , .C2( u1_u7_u7_n171 ) , .B( u1_u7_u7_n94 ) );
  AND2_X1 u1_u7_u7_U70 (.A2( u1_u7_X_43 ) , .A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n96 ) );
  AND2_X1 u1_u7_u7_U71 (.A2( u1_u7_X_45 ) , .A1( u1_u7_X_48 ) , .ZN( u1_u7_u7_n102 ) );
  AND2_X1 u1_u7_u7_U72 (.A1( u1_u7_X_48 ) , .A2( u1_u7_u7_n166 ) , .ZN( u1_u7_u7_n93 ) );
  INV_X1 u1_u7_u7_U73 (.A( u1_u7_X_46 ) , .ZN( u1_u7_u7_n163 ) );
  AND2_X1 u1_u7_u7_U74 (.A1( u1_u7_X_44 ) , .ZN( u1_u7_u7_n100 ) , .A2( u1_u7_u7_n167 ) );
  INV_X1 u1_u7_u7_U75 (.A( u1_u7_X_45 ) , .ZN( u1_u7_u7_n166 ) );
  INV_X1 u1_u7_u7_U76 (.A( u1_u7_X_43 ) , .ZN( u1_u7_u7_n167 ) );
  NAND4_X1 u1_u7_u7_U77 (.ZN( u1_out7_5 ) , .A4( u1_u7_u7_n108 ) , .A3( u1_u7_u7_n109 ) , .A1( u1_u7_u7_n116 ) , .A2( u1_u7_u7_n123 ) );
  AOI22_X1 u1_u7_u7_U78 (.ZN( u1_u7_u7_n109 ) , .A2( u1_u7_u7_n126 ) , .B2( u1_u7_u7_n145 ) , .B1( u1_u7_u7_n156 ) , .A1( u1_u7_u7_n171 ) );
  NOR4_X1 u1_u7_u7_U79 (.A4( u1_u7_u7_n104 ) , .A3( u1_u7_u7_n105 ) , .A2( u1_u7_u7_n106 ) , .A1( u1_u7_u7_n107 ) , .ZN( u1_u7_u7_n108 ) );
  OAI222_X1 u1_u7_u7_U8 (.C2( u1_u7_u7_n101 ) , .B2( u1_u7_u7_n111 ) , .A1( u1_u7_u7_n113 ) , .C1( u1_u7_u7_n146 ) , .A2( u1_u7_u7_n162 ) , .B1( u1_u7_u7_n164 ) , .ZN( u1_u7_u7_n94 ) );
  NAND4_X1 u1_u7_u7_U80 (.ZN( u1_out7_27 ) , .A4( u1_u7_u7_n118 ) , .A3( u1_u7_u7_n119 ) , .A2( u1_u7_u7_n120 ) , .A1( u1_u7_u7_n121 ) );
  OAI21_X1 u1_u7_u7_U81 (.ZN( u1_u7_u7_n121 ) , .B2( u1_u7_u7_n145 ) , .A( u1_u7_u7_n150 ) , .B1( u1_u7_u7_n174 ) );
  OAI21_X1 u1_u7_u7_U82 (.ZN( u1_u7_u7_n120 ) , .A( u1_u7_u7_n161 ) , .B2( u1_u7_u7_n170 ) , .B1( u1_u7_u7_n179 ) );
  NAND4_X1 u1_u7_u7_U83 (.ZN( u1_out7_21 ) , .A4( u1_u7_u7_n157 ) , .A3( u1_u7_u7_n158 ) , .A2( u1_u7_u7_n159 ) , .A1( u1_u7_u7_n160 ) );
  OAI21_X1 u1_u7_u7_U84 (.B1( u1_u7_u7_n145 ) , .ZN( u1_u7_u7_n160 ) , .A( u1_u7_u7_n161 ) , .B2( u1_u7_u7_n177 ) );
  AOI22_X1 u1_u7_u7_U85 (.B2( u1_u7_u7_n149 ) , .B1( u1_u7_u7_n150 ) , .A2( u1_u7_u7_n151 ) , .A1( u1_u7_u7_n152 ) , .ZN( u1_u7_u7_n158 ) );
  NAND4_X1 u1_u7_u7_U86 (.ZN( u1_out7_15 ) , .A4( u1_u7_u7_n142 ) , .A3( u1_u7_u7_n143 ) , .A2( u1_u7_u7_n144 ) , .A1( u1_u7_u7_n178 ) );
  OR2_X1 u1_u7_u7_U87 (.A2( u1_u7_u7_n125 ) , .A1( u1_u7_u7_n129 ) , .ZN( u1_u7_u7_n144 ) );
  AOI22_X1 u1_u7_u7_U88 (.A2( u1_u7_u7_n126 ) , .ZN( u1_u7_u7_n143 ) , .B2( u1_u7_u7_n165 ) , .B1( u1_u7_u7_n173 ) , .A1( u1_u7_u7_n174 ) );
  NAND2_X1 u1_u7_u7_U89 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n148 ) , .A2( u1_u7_u7_n95 ) );
  INV_X1 u1_u7_u7_U9 (.A( u1_u7_u7_n133 ) , .ZN( u1_u7_u7_n176 ) );
  NAND2_X1 u1_u7_u7_U90 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n113 ) , .A2( u1_u7_u7_n93 ) );
  NAND2_X1 u1_u7_u7_U91 (.A1( u1_u7_u7_n100 ) , .ZN( u1_u7_u7_n138 ) , .A2( u1_u7_u7_n99 ) );
  NAND2_X1 u1_u7_u7_U92 (.A1( u1_u7_u7_n100 ) , .A2( u1_u7_u7_n102 ) , .ZN( u1_u7_u7_n129 ) );
  OAI211_X1 u1_u7_u7_U93 (.B( u1_u7_u7_n122 ) , .A( u1_u7_u7_n123 ) , .C2( u1_u7_u7_n124 ) , .ZN( u1_u7_u7_n154 ) , .C1( u1_u7_u7_n162 ) );
  AOI222_X1 u1_u7_u7_U94 (.ZN( u1_u7_u7_n122 ) , .C2( u1_u7_u7_n126 ) , .C1( u1_u7_u7_n145 ) , .B1( u1_u7_u7_n161 ) , .A2( u1_u7_u7_n165 ) , .B2( u1_u7_u7_n170 ) , .A1( u1_u7_u7_n176 ) );
  NAND3_X1 u1_u7_u7_U95 (.A3( u1_u7_u7_n146 ) , .A2( u1_u7_u7_n147 ) , .A1( u1_u7_u7_n148 ) , .ZN( u1_u7_u7_n151 ) );
  NAND3_X1 u1_u7_u7_U96 (.A3( u1_u7_u7_n131 ) , .A2( u1_u7_u7_n132 ) , .A1( u1_u7_u7_n133 ) , .ZN( u1_u7_u7_n135 ) );
  XOR2_X1 u1_u9_U13 (.B( u1_K10_42 ) , .A( u1_R8_29 ) , .Z( u1_u9_X_42 ) );
  XOR2_X1 u1_u9_U14 (.B( u1_K10_41 ) , .A( u1_R8_28 ) , .Z( u1_u9_X_41 ) );
  XOR2_X1 u1_u9_U15 (.B( u1_K10_40 ) , .A( u1_R8_27 ) , .Z( u1_u9_X_40 ) );
  XOR2_X1 u1_u9_U17 (.B( u1_K10_39 ) , .A( u1_R8_26 ) , .Z( u1_u9_X_39 ) );
  XOR2_X1 u1_u9_U18 (.B( u1_K10_38 ) , .A( u1_R8_25 ) , .Z( u1_u9_X_38 ) );
  XOR2_X1 u1_u9_U19 (.B( u1_K10_37 ) , .A( u1_R8_24 ) , .Z( u1_u9_X_37 ) );
  XOR2_X1 u1_u9_U20 (.B( u1_K10_36 ) , .A( u1_R8_25 ) , .Z( u1_u9_X_36 ) );
  XOR2_X1 u1_u9_U21 (.B( u1_K10_35 ) , .A( u1_R8_24 ) , .Z( u1_u9_X_35 ) );
  XOR2_X1 u1_u9_U22 (.B( u1_K10_34 ) , .A( u1_R8_23 ) , .Z( u1_u9_X_34 ) );
  XOR2_X1 u1_u9_U23 (.B( u1_K10_33 ) , .A( u1_R8_22 ) , .Z( u1_u9_X_33 ) );
  XOR2_X1 u1_u9_U24 (.B( u1_K10_32 ) , .A( u1_R8_21 ) , .Z( u1_u9_X_32 ) );
  XOR2_X1 u1_u9_U25 (.B( u1_K10_31 ) , .A( u1_R8_20 ) , .Z( u1_u9_X_31 ) );
  NOR2_X1 u1_u9_u5_U10 (.ZN( u1_u9_u5_n135 ) , .A1( u1_u9_u5_n173 ) , .A2( u1_u9_u5_n176 ) );
  NOR3_X1 u1_u9_u5_U100 (.A3( u1_u9_u5_n141 ) , .A1( u1_u9_u5_n142 ) , .ZN( u1_u9_u5_n143 ) , .A2( u1_u9_u5_n191 ) );
  NAND4_X1 u1_u9_u5_U101 (.ZN( u1_out9_4 ) , .A4( u1_u9_u5_n112 ) , .A2( u1_u9_u5_n113 ) , .A1( u1_u9_u5_n114 ) , .A3( u1_u9_u5_n195 ) );
  AOI211_X1 u1_u9_u5_U102 (.A( u1_u9_u5_n110 ) , .C1( u1_u9_u5_n111 ) , .ZN( u1_u9_u5_n112 ) , .B( u1_u9_u5_n118 ) , .C2( u1_u9_u5_n177 ) );
  INV_X1 u1_u9_u5_U103 (.A( u1_u9_u5_n102 ) , .ZN( u1_u9_u5_n195 ) );
  NAND3_X1 u1_u9_u5_U104 (.A2( u1_u9_u5_n154 ) , .A3( u1_u9_u5_n158 ) , .A1( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n99 ) );
  INV_X1 u1_u9_u5_U11 (.A( u1_u9_u5_n121 ) , .ZN( u1_u9_u5_n177 ) );
  NOR2_X1 u1_u9_u5_U12 (.ZN( u1_u9_u5_n160 ) , .A2( u1_u9_u5_n173 ) , .A1( u1_u9_u5_n177 ) );
  INV_X1 u1_u9_u5_U13 (.A( u1_u9_u5_n150 ) , .ZN( u1_u9_u5_n174 ) );
  AOI21_X1 u1_u9_u5_U14 (.A( u1_u9_u5_n160 ) , .B2( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n162 ) , .B1( u1_u9_u5_n192 ) );
  INV_X1 u1_u9_u5_U15 (.A( u1_u9_u5_n159 ) , .ZN( u1_u9_u5_n192 ) );
  AOI21_X1 u1_u9_u5_U16 (.A( u1_u9_u5_n156 ) , .B2( u1_u9_u5_n157 ) , .B1( u1_u9_u5_n158 ) , .ZN( u1_u9_u5_n163 ) );
  AOI21_X1 u1_u9_u5_U17 (.B2( u1_u9_u5_n139 ) , .B1( u1_u9_u5_n140 ) , .ZN( u1_u9_u5_n141 ) , .A( u1_u9_u5_n150 ) );
  OAI21_X1 u1_u9_u5_U18 (.A( u1_u9_u5_n133 ) , .B2( u1_u9_u5_n134 ) , .B1( u1_u9_u5_n135 ) , .ZN( u1_u9_u5_n142 ) );
  OAI21_X1 u1_u9_u5_U19 (.ZN( u1_u9_u5_n133 ) , .B2( u1_u9_u5_n147 ) , .A( u1_u9_u5_n173 ) , .B1( u1_u9_u5_n188 ) );
  NAND2_X1 u1_u9_u5_U20 (.A2( u1_u9_u5_n119 ) , .A1( u1_u9_u5_n123 ) , .ZN( u1_u9_u5_n137 ) );
  INV_X1 u1_u9_u5_U21 (.A( u1_u9_u5_n155 ) , .ZN( u1_u9_u5_n194 ) );
  NAND2_X1 u1_u9_u5_U22 (.A1( u1_u9_u5_n121 ) , .ZN( u1_u9_u5_n132 ) , .A2( u1_u9_u5_n172 ) );
  NAND2_X1 u1_u9_u5_U23 (.A2( u1_u9_u5_n122 ) , .ZN( u1_u9_u5_n136 ) , .A1( u1_u9_u5_n154 ) );
  NAND2_X1 u1_u9_u5_U24 (.A2( u1_u9_u5_n119 ) , .A1( u1_u9_u5_n120 ) , .ZN( u1_u9_u5_n159 ) );
  INV_X1 u1_u9_u5_U25 (.A( u1_u9_u5_n156 ) , .ZN( u1_u9_u5_n175 ) );
  INV_X1 u1_u9_u5_U26 (.A( u1_u9_u5_n158 ) , .ZN( u1_u9_u5_n188 ) );
  INV_X1 u1_u9_u5_U27 (.A( u1_u9_u5_n152 ) , .ZN( u1_u9_u5_n179 ) );
  INV_X1 u1_u9_u5_U28 (.A( u1_u9_u5_n140 ) , .ZN( u1_u9_u5_n182 ) );
  INV_X1 u1_u9_u5_U29 (.A( u1_u9_u5_n151 ) , .ZN( u1_u9_u5_n183 ) );
  NOR2_X1 u1_u9_u5_U3 (.ZN( u1_u9_u5_n134 ) , .A1( u1_u9_u5_n183 ) , .A2( u1_u9_u5_n190 ) );
  INV_X1 u1_u9_u5_U30 (.A( u1_u9_u5_n123 ) , .ZN( u1_u9_u5_n185 ) );
  INV_X1 u1_u9_u5_U31 (.A( u1_u9_u5_n161 ) , .ZN( u1_u9_u5_n184 ) );
  INV_X1 u1_u9_u5_U32 (.A( u1_u9_u5_n139 ) , .ZN( u1_u9_u5_n189 ) );
  INV_X1 u1_u9_u5_U33 (.A( u1_u9_u5_n157 ) , .ZN( u1_u9_u5_n190 ) );
  INV_X1 u1_u9_u5_U34 (.A( u1_u9_u5_n120 ) , .ZN( u1_u9_u5_n193 ) );
  NAND2_X1 u1_u9_u5_U35 (.ZN( u1_u9_u5_n111 ) , .A1( u1_u9_u5_n140 ) , .A2( u1_u9_u5_n155 ) );
  NOR2_X1 u1_u9_u5_U36 (.ZN( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n170 ) , .A2( u1_u9_u5_n180 ) );
  INV_X1 u1_u9_u5_U37 (.A( u1_u9_u5_n117 ) , .ZN( u1_u9_u5_n196 ) );
  OAI221_X1 u1_u9_u5_U38 (.A( u1_u9_u5_n116 ) , .ZN( u1_u9_u5_n117 ) , .B2( u1_u9_u5_n119 ) , .C1( u1_u9_u5_n153 ) , .C2( u1_u9_u5_n158 ) , .B1( u1_u9_u5_n172 ) );
  AOI222_X1 u1_u9_u5_U39 (.ZN( u1_u9_u5_n116 ) , .B2( u1_u9_u5_n145 ) , .C1( u1_u9_u5_n148 ) , .A2( u1_u9_u5_n174 ) , .C2( u1_u9_u5_n177 ) , .B1( u1_u9_u5_n187 ) , .A1( u1_u9_u5_n193 ) );
  INV_X1 u1_u9_u5_U4 (.A( u1_u9_u5_n138 ) , .ZN( u1_u9_u5_n191 ) );
  INV_X1 u1_u9_u5_U40 (.A( u1_u9_u5_n115 ) , .ZN( u1_u9_u5_n187 ) );
  OAI221_X1 u1_u9_u5_U41 (.A( u1_u9_u5_n101 ) , .ZN( u1_u9_u5_n102 ) , .C2( u1_u9_u5_n115 ) , .C1( u1_u9_u5_n126 ) , .B1( u1_u9_u5_n134 ) , .B2( u1_u9_u5_n160 ) );
  OAI21_X1 u1_u9_u5_U42 (.ZN( u1_u9_u5_n101 ) , .B1( u1_u9_u5_n137 ) , .A( u1_u9_u5_n146 ) , .B2( u1_u9_u5_n147 ) );
  AOI22_X1 u1_u9_u5_U43 (.B2( u1_u9_u5_n131 ) , .A2( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n169 ) , .B1( u1_u9_u5_n174 ) , .A1( u1_u9_u5_n185 ) );
  NOR2_X1 u1_u9_u5_U44 (.A1( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n150 ) , .A2( u1_u9_u5_n173 ) );
  AOI21_X1 u1_u9_u5_U45 (.A( u1_u9_u5_n118 ) , .B2( u1_u9_u5_n145 ) , .ZN( u1_u9_u5_n168 ) , .B1( u1_u9_u5_n186 ) );
  INV_X1 u1_u9_u5_U46 (.A( u1_u9_u5_n122 ) , .ZN( u1_u9_u5_n186 ) );
  NOR2_X1 u1_u9_u5_U47 (.A1( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n152 ) , .A2( u1_u9_u5_n176 ) );
  NOR2_X1 u1_u9_u5_U48 (.A1( u1_u9_u5_n115 ) , .ZN( u1_u9_u5_n118 ) , .A2( u1_u9_u5_n153 ) );
  NOR2_X1 u1_u9_u5_U49 (.A2( u1_u9_u5_n145 ) , .ZN( u1_u9_u5_n156 ) , .A1( u1_u9_u5_n174 ) );
  OAI21_X1 u1_u9_u5_U5 (.B2( u1_u9_u5_n136 ) , .B1( u1_u9_u5_n137 ) , .ZN( u1_u9_u5_n138 ) , .A( u1_u9_u5_n177 ) );
  NOR2_X1 u1_u9_u5_U50 (.ZN( u1_u9_u5_n121 ) , .A2( u1_u9_u5_n145 ) , .A1( u1_u9_u5_n176 ) );
  AOI22_X1 u1_u9_u5_U51 (.ZN( u1_u9_u5_n114 ) , .A2( u1_u9_u5_n137 ) , .A1( u1_u9_u5_n145 ) , .B2( u1_u9_u5_n175 ) , .B1( u1_u9_u5_n193 ) );
  OAI211_X1 u1_u9_u5_U52 (.B( u1_u9_u5_n124 ) , .A( u1_u9_u5_n125 ) , .C2( u1_u9_u5_n126 ) , .C1( u1_u9_u5_n127 ) , .ZN( u1_u9_u5_n128 ) );
  NOR3_X1 u1_u9_u5_U53 (.ZN( u1_u9_u5_n127 ) , .A1( u1_u9_u5_n136 ) , .A3( u1_u9_u5_n148 ) , .A2( u1_u9_u5_n182 ) );
  OAI21_X1 u1_u9_u5_U54 (.ZN( u1_u9_u5_n124 ) , .A( u1_u9_u5_n177 ) , .B2( u1_u9_u5_n183 ) , .B1( u1_u9_u5_n189 ) );
  OAI21_X1 u1_u9_u5_U55 (.ZN( u1_u9_u5_n125 ) , .A( u1_u9_u5_n174 ) , .B2( u1_u9_u5_n185 ) , .B1( u1_u9_u5_n190 ) );
  AOI21_X1 u1_u9_u5_U56 (.A( u1_u9_u5_n153 ) , .B2( u1_u9_u5_n154 ) , .B1( u1_u9_u5_n155 ) , .ZN( u1_u9_u5_n164 ) );
  AOI21_X1 u1_u9_u5_U57 (.ZN( u1_u9_u5_n110 ) , .B1( u1_u9_u5_n122 ) , .B2( u1_u9_u5_n139 ) , .A( u1_u9_u5_n153 ) );
  INV_X1 u1_u9_u5_U58 (.A( u1_u9_u5_n153 ) , .ZN( u1_u9_u5_n176 ) );
  INV_X1 u1_u9_u5_U59 (.A( u1_u9_u5_n126 ) , .ZN( u1_u9_u5_n173 ) );
  AOI222_X1 u1_u9_u5_U6 (.ZN( u1_u9_u5_n113 ) , .A1( u1_u9_u5_n131 ) , .C1( u1_u9_u5_n148 ) , .B2( u1_u9_u5_n174 ) , .C2( u1_u9_u5_n178 ) , .A2( u1_u9_u5_n179 ) , .B1( u1_u9_u5_n99 ) );
  AND2_X1 u1_u9_u5_U60 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n147 ) );
  AND2_X1 u1_u9_u5_U61 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n148 ) );
  NAND2_X1 u1_u9_u5_U62 (.A1( u1_u9_u5_n105 ) , .A2( u1_u9_u5_n106 ) , .ZN( u1_u9_u5_n158 ) );
  NAND2_X1 u1_u9_u5_U63 (.A2( u1_u9_u5_n108 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n139 ) );
  NAND2_X1 u1_u9_u5_U64 (.A1( u1_u9_u5_n106 ) , .A2( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n119 ) );
  NAND2_X1 u1_u9_u5_U65 (.A2( u1_u9_u5_n103 ) , .A1( u1_u9_u5_n105 ) , .ZN( u1_u9_u5_n140 ) );
  NAND2_X1 u1_u9_u5_U66 (.A2( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n105 ) , .ZN( u1_u9_u5_n155 ) );
  NAND2_X1 u1_u9_u5_U67 (.A2( u1_u9_u5_n106 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n122 ) );
  NAND2_X1 u1_u9_u5_U68 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n106 ) , .ZN( u1_u9_u5_n115 ) );
  NAND2_X1 u1_u9_u5_U69 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n103 ) , .ZN( u1_u9_u5_n161 ) );
  INV_X1 u1_u9_u5_U7 (.A( u1_u9_u5_n135 ) , .ZN( u1_u9_u5_n178 ) );
  NAND2_X1 u1_u9_u5_U70 (.A1( u1_u9_u5_n105 ) , .A2( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n154 ) );
  INV_X1 u1_u9_u5_U71 (.A( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n172 ) );
  NAND2_X1 u1_u9_u5_U72 (.A1( u1_u9_u5_n103 ) , .A2( u1_u9_u5_n108 ) , .ZN( u1_u9_u5_n123 ) );
  NAND2_X1 u1_u9_u5_U73 (.A2( u1_u9_u5_n103 ) , .A1( u1_u9_u5_n107 ) , .ZN( u1_u9_u5_n151 ) );
  NAND2_X1 u1_u9_u5_U74 (.A2( u1_u9_u5_n107 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n120 ) );
  NAND2_X1 u1_u9_u5_U75 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n109 ) , .ZN( u1_u9_u5_n157 ) );
  AND2_X1 u1_u9_u5_U76 (.A2( u1_u9_u5_n100 ) , .A1( u1_u9_u5_n104 ) , .ZN( u1_u9_u5_n131 ) );
  NOR2_X1 u1_u9_u5_U77 (.A2( u1_u9_X_34 ) , .A1( u1_u9_X_35 ) , .ZN( u1_u9_u5_n145 ) );
  NOR2_X1 u1_u9_u5_U78 (.A2( u1_u9_X_34 ) , .ZN( u1_u9_u5_n146 ) , .A1( u1_u9_u5_n171 ) );
  NOR2_X1 u1_u9_u5_U79 (.A2( u1_u9_X_31 ) , .A1( u1_u9_X_32 ) , .ZN( u1_u9_u5_n103 ) );
  OAI22_X1 u1_u9_u5_U8 (.B2( u1_u9_u5_n149 ) , .B1( u1_u9_u5_n150 ) , .A2( u1_u9_u5_n151 ) , .A1( u1_u9_u5_n152 ) , .ZN( u1_u9_u5_n165 ) );
  NOR2_X1 u1_u9_u5_U80 (.A2( u1_u9_X_36 ) , .ZN( u1_u9_u5_n105 ) , .A1( u1_u9_u5_n180 ) );
  NOR2_X1 u1_u9_u5_U81 (.A2( u1_u9_X_33 ) , .ZN( u1_u9_u5_n108 ) , .A1( u1_u9_u5_n170 ) );
  NOR2_X1 u1_u9_u5_U82 (.A2( u1_u9_X_33 ) , .A1( u1_u9_X_36 ) , .ZN( u1_u9_u5_n107 ) );
  NOR2_X1 u1_u9_u5_U83 (.A2( u1_u9_X_31 ) , .ZN( u1_u9_u5_n104 ) , .A1( u1_u9_u5_n181 ) );
  NAND2_X1 u1_u9_u5_U84 (.A2( u1_u9_X_34 ) , .A1( u1_u9_X_35 ) , .ZN( u1_u9_u5_n153 ) );
  NAND2_X1 u1_u9_u5_U85 (.A1( u1_u9_X_34 ) , .ZN( u1_u9_u5_n126 ) , .A2( u1_u9_u5_n171 ) );
  AND2_X1 u1_u9_u5_U86 (.A1( u1_u9_X_31 ) , .A2( u1_u9_X_32 ) , .ZN( u1_u9_u5_n106 ) );
  AND2_X1 u1_u9_u5_U87 (.A1( u1_u9_X_31 ) , .ZN( u1_u9_u5_n109 ) , .A2( u1_u9_u5_n181 ) );
  INV_X1 u1_u9_u5_U88 (.A( u1_u9_X_33 ) , .ZN( u1_u9_u5_n180 ) );
  INV_X1 u1_u9_u5_U89 (.A( u1_u9_X_35 ) , .ZN( u1_u9_u5_n171 ) );
  NOR3_X1 u1_u9_u5_U9 (.A2( u1_u9_u5_n147 ) , .A1( u1_u9_u5_n148 ) , .ZN( u1_u9_u5_n149 ) , .A3( u1_u9_u5_n194 ) );
  INV_X1 u1_u9_u5_U90 (.A( u1_u9_X_36 ) , .ZN( u1_u9_u5_n170 ) );
  INV_X1 u1_u9_u5_U91 (.A( u1_u9_X_32 ) , .ZN( u1_u9_u5_n181 ) );
  NAND4_X1 u1_u9_u5_U92 (.ZN( u1_out9_29 ) , .A4( u1_u9_u5_n129 ) , .A3( u1_u9_u5_n130 ) , .A2( u1_u9_u5_n168 ) , .A1( u1_u9_u5_n196 ) );
  AOI221_X1 u1_u9_u5_U93 (.A( u1_u9_u5_n128 ) , .ZN( u1_u9_u5_n129 ) , .C2( u1_u9_u5_n132 ) , .B2( u1_u9_u5_n159 ) , .B1( u1_u9_u5_n176 ) , .C1( u1_u9_u5_n184 ) );
  AOI222_X1 u1_u9_u5_U94 (.ZN( u1_u9_u5_n130 ) , .A2( u1_u9_u5_n146 ) , .B1( u1_u9_u5_n147 ) , .C2( u1_u9_u5_n175 ) , .B2( u1_u9_u5_n179 ) , .A1( u1_u9_u5_n188 ) , .C1( u1_u9_u5_n194 ) );
  NAND4_X1 u1_u9_u5_U95 (.ZN( u1_out9_19 ) , .A4( u1_u9_u5_n166 ) , .A3( u1_u9_u5_n167 ) , .A2( u1_u9_u5_n168 ) , .A1( u1_u9_u5_n169 ) );
  AOI22_X1 u1_u9_u5_U96 (.B2( u1_u9_u5_n145 ) , .A2( u1_u9_u5_n146 ) , .ZN( u1_u9_u5_n167 ) , .B1( u1_u9_u5_n182 ) , .A1( u1_u9_u5_n189 ) );
  NOR4_X1 u1_u9_u5_U97 (.A4( u1_u9_u5_n162 ) , .A3( u1_u9_u5_n163 ) , .A2( u1_u9_u5_n164 ) , .A1( u1_u9_u5_n165 ) , .ZN( u1_u9_u5_n166 ) );
  NAND4_X1 u1_u9_u5_U98 (.ZN( u1_out9_11 ) , .A4( u1_u9_u5_n143 ) , .A3( u1_u9_u5_n144 ) , .A2( u1_u9_u5_n169 ) , .A1( u1_u9_u5_n196 ) );
  AOI22_X1 u1_u9_u5_U99 (.A2( u1_u9_u5_n132 ) , .ZN( u1_u9_u5_n144 ) , .B2( u1_u9_u5_n145 ) , .B1( u1_u9_u5_n184 ) , .A1( u1_u9_u5_n194 ) );
  AOI22_X1 u1_u9_u6_U10 (.A2( u1_u9_u6_n151 ) , .B2( u1_u9_u6_n161 ) , .A1( u1_u9_u6_n167 ) , .B1( u1_u9_u6_n170 ) , .ZN( u1_u9_u6_n89 ) );
  AOI21_X1 u1_u9_u6_U11 (.B1( u1_u9_u6_n107 ) , .B2( u1_u9_u6_n132 ) , .A( u1_u9_u6_n158 ) , .ZN( u1_u9_u6_n88 ) );
  AOI21_X1 u1_u9_u6_U12 (.B2( u1_u9_u6_n147 ) , .B1( u1_u9_u6_n148 ) , .ZN( u1_u9_u6_n149 ) , .A( u1_u9_u6_n158 ) );
  AOI21_X1 u1_u9_u6_U13 (.ZN( u1_u9_u6_n106 ) , .A( u1_u9_u6_n142 ) , .B2( u1_u9_u6_n159 ) , .B1( u1_u9_u6_n164 ) );
  INV_X1 u1_u9_u6_U14 (.A( u1_u9_u6_n155 ) , .ZN( u1_u9_u6_n161 ) );
  INV_X1 u1_u9_u6_U15 (.A( u1_u9_u6_n128 ) , .ZN( u1_u9_u6_n164 ) );
  NAND2_X1 u1_u9_u6_U16 (.ZN( u1_u9_u6_n110 ) , .A1( u1_u9_u6_n122 ) , .A2( u1_u9_u6_n129 ) );
  NAND2_X1 u1_u9_u6_U17 (.ZN( u1_u9_u6_n124 ) , .A2( u1_u9_u6_n146 ) , .A1( u1_u9_u6_n148 ) );
  INV_X1 u1_u9_u6_U18 (.A( u1_u9_u6_n132 ) , .ZN( u1_u9_u6_n171 ) );
  AND2_X1 u1_u9_u6_U19 (.A1( u1_u9_u6_n100 ) , .ZN( u1_u9_u6_n130 ) , .A2( u1_u9_u6_n147 ) );
  INV_X1 u1_u9_u6_U20 (.A( u1_u9_u6_n127 ) , .ZN( u1_u9_u6_n173 ) );
  INV_X1 u1_u9_u6_U21 (.A( u1_u9_u6_n121 ) , .ZN( u1_u9_u6_n167 ) );
  INV_X1 u1_u9_u6_U22 (.A( u1_u9_u6_n100 ) , .ZN( u1_u9_u6_n169 ) );
  INV_X1 u1_u9_u6_U23 (.A( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n170 ) );
  INV_X1 u1_u9_u6_U24 (.A( u1_u9_u6_n113 ) , .ZN( u1_u9_u6_n168 ) );
  AND2_X1 u1_u9_u6_U25 (.A1( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n119 ) , .ZN( u1_u9_u6_n133 ) );
  AND2_X1 u1_u9_u6_U26 (.A2( u1_u9_u6_n121 ) , .A1( u1_u9_u6_n122 ) , .ZN( u1_u9_u6_n131 ) );
  AND3_X1 u1_u9_u6_U27 (.ZN( u1_u9_u6_n120 ) , .A2( u1_u9_u6_n127 ) , .A1( u1_u9_u6_n132 ) , .A3( u1_u9_u6_n145 ) );
  INV_X1 u1_u9_u6_U28 (.A( u1_u9_u6_n146 ) , .ZN( u1_u9_u6_n163 ) );
  AOI222_X1 u1_u9_u6_U29 (.ZN( u1_u9_u6_n114 ) , .A1( u1_u9_u6_n118 ) , .A2( u1_u9_u6_n126 ) , .B2( u1_u9_u6_n151 ) , .C2( u1_u9_u6_n159 ) , .C1( u1_u9_u6_n168 ) , .B1( u1_u9_u6_n169 ) );
  INV_X1 u1_u9_u6_U3 (.A( u1_u9_u6_n110 ) , .ZN( u1_u9_u6_n166 ) );
  NOR2_X1 u1_u9_u6_U30 (.A1( u1_u9_u6_n162 ) , .A2( u1_u9_u6_n165 ) , .ZN( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U31 (.A1( u1_u9_u6_n144 ) , .ZN( u1_u9_u6_n151 ) , .A2( u1_u9_u6_n158 ) );
  NAND2_X1 u1_u9_u6_U32 (.ZN( u1_u9_u6_n132 ) , .A1( u1_u9_u6_n91 ) , .A2( u1_u9_u6_n97 ) );
  AOI22_X1 u1_u9_u6_U33 (.B2( u1_u9_u6_n110 ) , .B1( u1_u9_u6_n111 ) , .A1( u1_u9_u6_n112 ) , .ZN( u1_u9_u6_n115 ) , .A2( u1_u9_u6_n161 ) );
  NAND4_X1 u1_u9_u6_U34 (.A3( u1_u9_u6_n109 ) , .ZN( u1_u9_u6_n112 ) , .A4( u1_u9_u6_n132 ) , .A2( u1_u9_u6_n147 ) , .A1( u1_u9_u6_n166 ) );
  NOR2_X1 u1_u9_u6_U35 (.ZN( u1_u9_u6_n109 ) , .A1( u1_u9_u6_n170 ) , .A2( u1_u9_u6_n173 ) );
  NOR2_X1 u1_u9_u6_U36 (.A2( u1_u9_u6_n126 ) , .ZN( u1_u9_u6_n155 ) , .A1( u1_u9_u6_n160 ) );
  NAND2_X1 u1_u9_u6_U37 (.ZN( u1_u9_u6_n146 ) , .A2( u1_u9_u6_n94 ) , .A1( u1_u9_u6_n99 ) );
  AOI21_X1 u1_u9_u6_U38 (.A( u1_u9_u6_n144 ) , .B2( u1_u9_u6_n145 ) , .B1( u1_u9_u6_n146 ) , .ZN( u1_u9_u6_n150 ) );
  AOI211_X1 u1_u9_u6_U39 (.B( u1_u9_u6_n134 ) , .A( u1_u9_u6_n135 ) , .C1( u1_u9_u6_n136 ) , .ZN( u1_u9_u6_n137 ) , .C2( u1_u9_u6_n151 ) );
  INV_X1 u1_u9_u6_U4 (.A( u1_u9_u6_n142 ) , .ZN( u1_u9_u6_n174 ) );
  NAND4_X1 u1_u9_u6_U40 (.A4( u1_u9_u6_n127 ) , .A3( u1_u9_u6_n128 ) , .A2( u1_u9_u6_n129 ) , .A1( u1_u9_u6_n130 ) , .ZN( u1_u9_u6_n136 ) );
  AOI21_X1 u1_u9_u6_U41 (.B2( u1_u9_u6_n132 ) , .B1( u1_u9_u6_n133 ) , .ZN( u1_u9_u6_n134 ) , .A( u1_u9_u6_n158 ) );
  AOI21_X1 u1_u9_u6_U42 (.B1( u1_u9_u6_n131 ) , .ZN( u1_u9_u6_n135 ) , .A( u1_u9_u6_n144 ) , .B2( u1_u9_u6_n146 ) );
  INV_X1 u1_u9_u6_U43 (.A( u1_u9_u6_n111 ) , .ZN( u1_u9_u6_n158 ) );
  NAND2_X1 u1_u9_u6_U44 (.ZN( u1_u9_u6_n127 ) , .A1( u1_u9_u6_n91 ) , .A2( u1_u9_u6_n92 ) );
  NAND2_X1 u1_u9_u6_U45 (.ZN( u1_u9_u6_n129 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n96 ) );
  INV_X1 u1_u9_u6_U46 (.A( u1_u9_u6_n144 ) , .ZN( u1_u9_u6_n159 ) );
  NAND2_X1 u1_u9_u6_U47 (.ZN( u1_u9_u6_n145 ) , .A2( u1_u9_u6_n97 ) , .A1( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U48 (.ZN( u1_u9_u6_n148 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n94 ) );
  NAND2_X1 u1_u9_u6_U49 (.ZN( u1_u9_u6_n108 ) , .A2( u1_u9_u6_n139 ) , .A1( u1_u9_u6_n144 ) );
  NAND2_X1 u1_u9_u6_U5 (.A2( u1_u9_u6_n143 ) , .ZN( u1_u9_u6_n152 ) , .A1( u1_u9_u6_n166 ) );
  NAND2_X1 u1_u9_u6_U50 (.ZN( u1_u9_u6_n121 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n97 ) );
  NAND2_X1 u1_u9_u6_U51 (.ZN( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n95 ) );
  AND2_X1 u1_u9_u6_U52 (.ZN( u1_u9_u6_n118 ) , .A2( u1_u9_u6_n91 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U53 (.ZN( u1_u9_u6_n147 ) , .A2( u1_u9_u6_n98 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U54 (.ZN( u1_u9_u6_n128 ) , .A1( u1_u9_u6_n94 ) , .A2( u1_u9_u6_n96 ) );
  NAND2_X1 u1_u9_u6_U55 (.ZN( u1_u9_u6_n119 ) , .A2( u1_u9_u6_n95 ) , .A1( u1_u9_u6_n99 ) );
  NAND2_X1 u1_u9_u6_U56 (.ZN( u1_u9_u6_n123 ) , .A2( u1_u9_u6_n91 ) , .A1( u1_u9_u6_n96 ) );
  NAND2_X1 u1_u9_u6_U57 (.ZN( u1_u9_u6_n100 ) , .A2( u1_u9_u6_n92 ) , .A1( u1_u9_u6_n98 ) );
  NAND2_X1 u1_u9_u6_U58 (.ZN( u1_u9_u6_n122 ) , .A1( u1_u9_u6_n94 ) , .A2( u1_u9_u6_n97 ) );
  INV_X1 u1_u9_u6_U59 (.A( u1_u9_u6_n139 ) , .ZN( u1_u9_u6_n160 ) );
  AOI22_X1 u1_u9_u6_U6 (.B2( u1_u9_u6_n101 ) , .A1( u1_u9_u6_n102 ) , .ZN( u1_u9_u6_n103 ) , .B1( u1_u9_u6_n160 ) , .A2( u1_u9_u6_n161 ) );
  NAND2_X1 u1_u9_u6_U60 (.ZN( u1_u9_u6_n113 ) , .A1( u1_u9_u6_n96 ) , .A2( u1_u9_u6_n98 ) );
  NOR2_X1 u1_u9_u6_U61 (.A2( u1_u9_X_40 ) , .A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n126 ) );
  NOR2_X1 u1_u9_u6_U62 (.A2( u1_u9_X_39 ) , .A1( u1_u9_X_42 ) , .ZN( u1_u9_u6_n92 ) );
  NOR2_X1 u1_u9_u6_U63 (.A2( u1_u9_X_39 ) , .A1( u1_u9_u6_n156 ) , .ZN( u1_u9_u6_n97 ) );
  NOR2_X1 u1_u9_u6_U64 (.A2( u1_u9_X_38 ) , .A1( u1_u9_u6_n165 ) , .ZN( u1_u9_u6_n95 ) );
  NOR2_X1 u1_u9_u6_U65 (.A2( u1_u9_X_41 ) , .ZN( u1_u9_u6_n111 ) , .A1( u1_u9_u6_n157 ) );
  NOR2_X1 u1_u9_u6_U66 (.A2( u1_u9_X_37 ) , .A1( u1_u9_u6_n162 ) , .ZN( u1_u9_u6_n94 ) );
  NOR2_X1 u1_u9_u6_U67 (.A2( u1_u9_X_37 ) , .A1( u1_u9_X_38 ) , .ZN( u1_u9_u6_n91 ) );
  NAND2_X1 u1_u9_u6_U68 (.A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n144 ) , .A2( u1_u9_u6_n157 ) );
  NAND2_X1 u1_u9_u6_U69 (.A2( u1_u9_X_40 ) , .A1( u1_u9_X_41 ) , .ZN( u1_u9_u6_n139 ) );
  NOR2_X1 u1_u9_u6_U7 (.A1( u1_u9_u6_n118 ) , .ZN( u1_u9_u6_n143 ) , .A2( u1_u9_u6_n168 ) );
  AND2_X1 u1_u9_u6_U70 (.A1( u1_u9_X_39 ) , .A2( u1_u9_u6_n156 ) , .ZN( u1_u9_u6_n96 ) );
  AND2_X1 u1_u9_u6_U71 (.A1( u1_u9_X_39 ) , .A2( u1_u9_X_42 ) , .ZN( u1_u9_u6_n99 ) );
  INV_X1 u1_u9_u6_U72 (.A( u1_u9_X_40 ) , .ZN( u1_u9_u6_n157 ) );
  INV_X1 u1_u9_u6_U73 (.A( u1_u9_X_37 ) , .ZN( u1_u9_u6_n165 ) );
  INV_X1 u1_u9_u6_U74 (.A( u1_u9_X_38 ) , .ZN( u1_u9_u6_n162 ) );
  INV_X1 u1_u9_u6_U75 (.A( u1_u9_X_42 ) , .ZN( u1_u9_u6_n156 ) );
  NAND4_X1 u1_u9_u6_U76 (.ZN( u1_out9_12 ) , .A4( u1_u9_u6_n114 ) , .A3( u1_u9_u6_n115 ) , .A2( u1_u9_u6_n116 ) , .A1( u1_u9_u6_n117 ) );
  OAI22_X1 u1_u9_u6_U77 (.B2( u1_u9_u6_n111 ) , .ZN( u1_u9_u6_n116 ) , .B1( u1_u9_u6_n126 ) , .A2( u1_u9_u6_n164 ) , .A1( u1_u9_u6_n167 ) );
  OAI21_X1 u1_u9_u6_U78 (.A( u1_u9_u6_n108 ) , .ZN( u1_u9_u6_n117 ) , .B2( u1_u9_u6_n141 ) , .B1( u1_u9_u6_n163 ) );
  NAND4_X1 u1_u9_u6_U79 (.ZN( u1_out9_32 ) , .A4( u1_u9_u6_n103 ) , .A3( u1_u9_u6_n104 ) , .A2( u1_u9_u6_n105 ) , .A1( u1_u9_u6_n106 ) );
  OAI21_X1 u1_u9_u6_U8 (.A( u1_u9_u6_n159 ) , .B1( u1_u9_u6_n169 ) , .B2( u1_u9_u6_n173 ) , .ZN( u1_u9_u6_n90 ) );
  AOI22_X1 u1_u9_u6_U80 (.ZN( u1_u9_u6_n105 ) , .A2( u1_u9_u6_n108 ) , .A1( u1_u9_u6_n118 ) , .B2( u1_u9_u6_n126 ) , .B1( u1_u9_u6_n171 ) );
  AOI22_X1 u1_u9_u6_U81 (.ZN( u1_u9_u6_n104 ) , .A1( u1_u9_u6_n111 ) , .B1( u1_u9_u6_n124 ) , .B2( u1_u9_u6_n151 ) , .A2( u1_u9_u6_n93 ) );
  OAI211_X1 u1_u9_u6_U82 (.ZN( u1_out9_7 ) , .B( u1_u9_u6_n153 ) , .C2( u1_u9_u6_n154 ) , .C1( u1_u9_u6_n155 ) , .A( u1_u9_u6_n174 ) );
  NOR3_X1 u1_u9_u6_U83 (.A1( u1_u9_u6_n141 ) , .ZN( u1_u9_u6_n154 ) , .A3( u1_u9_u6_n164 ) , .A2( u1_u9_u6_n171 ) );
  AOI211_X1 u1_u9_u6_U84 (.B( u1_u9_u6_n149 ) , .A( u1_u9_u6_n150 ) , .C2( u1_u9_u6_n151 ) , .C1( u1_u9_u6_n152 ) , .ZN( u1_u9_u6_n153 ) );
  OAI211_X1 u1_u9_u6_U85 (.ZN( u1_out9_22 ) , .B( u1_u9_u6_n137 ) , .A( u1_u9_u6_n138 ) , .C2( u1_u9_u6_n139 ) , .C1( u1_u9_u6_n140 ) );
  AOI22_X1 u1_u9_u6_U86 (.B1( u1_u9_u6_n124 ) , .A2( u1_u9_u6_n125 ) , .A1( u1_u9_u6_n126 ) , .ZN( u1_u9_u6_n138 ) , .B2( u1_u9_u6_n161 ) );
  AND4_X1 u1_u9_u6_U87 (.A3( u1_u9_u6_n119 ) , .A1( u1_u9_u6_n120 ) , .A4( u1_u9_u6_n129 ) , .ZN( u1_u9_u6_n140 ) , .A2( u1_u9_u6_n143 ) );
  NAND3_X1 u1_u9_u6_U88 (.A2( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n125 ) , .A1( u1_u9_u6_n130 ) , .A3( u1_u9_u6_n131 ) );
  NAND3_X1 u1_u9_u6_U89 (.A3( u1_u9_u6_n133 ) , .ZN( u1_u9_u6_n141 ) , .A1( u1_u9_u6_n145 ) , .A2( u1_u9_u6_n148 ) );
  INV_X1 u1_u9_u6_U9 (.ZN( u1_u9_u6_n172 ) , .A( u1_u9_u6_n88 ) );
  NAND3_X1 u1_u9_u6_U90 (.ZN( u1_u9_u6_n101 ) , .A3( u1_u9_u6_n107 ) , .A2( u1_u9_u6_n121 ) , .A1( u1_u9_u6_n127 ) );
  NAND3_X1 u1_u9_u6_U91 (.ZN( u1_u9_u6_n102 ) , .A3( u1_u9_u6_n130 ) , .A2( u1_u9_u6_n145 ) , .A1( u1_u9_u6_n166 ) );
  NAND3_X1 u1_u9_u6_U92 (.A3( u1_u9_u6_n113 ) , .A1( u1_u9_u6_n119 ) , .A2( u1_u9_u6_n123 ) , .ZN( u1_u9_u6_n93 ) );
  NAND3_X1 u1_u9_u6_U93 (.ZN( u1_u9_u6_n142 ) , .A2( u1_u9_u6_n172 ) , .A3( u1_u9_u6_n89 ) , .A1( u1_u9_u6_n90 ) );
  INV_X1 u1_uk_U10 (.A( u1_uk_n209 ) , .ZN( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1006 (.ZN( u1_K16_4 ) , .B2( u1_uk_n1257 ) , .B1( u1_uk_n99 ) , .A( u1_uk_n995 ) );
  NAND2_X1 u1_uk_U1007 (.A1( u1_uk_K_r14_3 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n995 ) );
  OAI21_X1 u1_uk_U1012 (.ZN( u1_K4_5 ) , .A( u1_uk_n1068 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1386 ) );
  NAND2_X1 u1_uk_U1013 (.A1( u1_uk_K_r2_53 ) , .ZN( u1_uk_n1068 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1036 (.ZN( u1_K8_46 ) , .A( u1_uk_n1145 ) , .B2( u1_uk_n1562 ) , .B1( u1_uk_n188 ) );
  NAND2_X1 u1_uk_U1037 (.A1( u1_uk_K_r6_37 ) , .ZN( u1_uk_n1145 ) , .A2( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U1040 (.ZN( u1_K12_36 ) , .B2( u1_uk_n1728 ) , .A( u1_uk_n587 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1041 (.A1( u1_uk_K_r10_52 ) , .A2( u1_uk_n110 ) , .ZN( u1_uk_n587 ) );
  OAI21_X1 u1_uk_U1060 (.ZN( u1_K12_40 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1729 ) , .A( u1_uk_n603 ) );
  NAND2_X1 u1_uk_U1061 (.A1( u1_uk_K_r10_49 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n603 ) );
  OAI21_X1 u1_uk_U1064 (.ZN( u1_K10_32 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1618 ) , .A( u1_uk_n346 ) );
  NAND2_X1 u1_uk_U1065 (.A1( u1_uk_K_r8_51 ) , .A2( u1_uk_n142 ) , .ZN( u1_uk_n346 ) );
  OAI22_X1 u1_uk_U108 (.ZN( u1_K16_5 ) , .A2( u1_uk_n1221 ) , .B2( u1_uk_n1224 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n294 ) );
  OAI21_X1 u1_uk_U110 (.ZN( u1_K14_5 ) , .B2( u1_uk_n1826 ) , .B1( u1_uk_n250 ) , .A( u1_uk_n962 ) );
  NAND2_X1 u1_uk_U111 (.A1( u1_uk_K_r12_10 ) , .A2( u1_uk_n298 ) , .ZN( u1_uk_n962 ) );
  INV_X1 u1_uk_U1141 (.ZN( u1_K12_32 ) , .A( u1_uk_n582 ) );
  AOI22_X1 u1_uk_U1142 (.B2( u1_uk_K_r10_23 ) , .A2( u1_uk_K_r10_28 ) , .B1( u1_uk_n10 ) , .A1( u1_uk_n294 ) , .ZN( u1_uk_n582 ) );
  INV_X1 u1_uk_U1147 (.ZN( u1_K4_20 ) , .A( u1_uk_n1054 ) );
  AOI22_X1 u1_uk_U1148 (.B2( u1_uk_K_r2_13 ) , .A2( u1_uk_K_r2_33 ) , .ZN( u1_uk_n1054 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n207 ) );
  INV_X1 u1_uk_U1171 (.ZN( u1_K4_2 ) , .A( u1_uk_n1061 ) );
  OAI22_X1 u1_uk_U119 (.ZN( u1_K10_41 ) , .A2( u1_uk_n1624 ) , .B2( u1_uk_n1652 ) , .A1( u1_uk_n223 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U121 (.ZN( u1_K12_41 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1735 ) , .A2( u1_uk_n1744 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U125 (.ZN( u1_K12_47 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1709 ) , .A2( u1_uk_n1736 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U129 (.ZN( u1_K8_47 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1561 ) , .A2( u1_uk_n1567 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U134 (.ZN( u1_K4_47 ) , .B2( u1_uk_n1380 ) , .A2( u1_uk_n1389 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U138 (.ZN( u1_K4_15 ) , .B2( u1_uk_n1358 ) , .A2( u1_uk_n1386 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U166 (.ZN( u1_K4_19 ) , .B2( u1_uk_n1365 ) , .A2( u1_uk_n1377 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U171 (.ZN( u1_K14_15 ) , .A1( u1_uk_n146 ) , .A2( u1_uk_n1803 ) , .B2( u1_uk_n1841 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U205 (.ZN( u1_K4_24 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1352 ) , .A2( u1_uk_n1393 ) , .B1( u1_uk_n213 ) );
  OAI21_X1 u1_uk_U224 (.ZN( u1_K12_31 ) , .B2( u1_uk_n1715 ) , .B1( u1_uk_n207 ) , .A( u1_uk_n551 ) );
  NAND2_X1 u1_uk_U225 (.A1( u1_uk_K_r10_44 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n551 ) );
  INV_X1 u1_uk_U23 (.ZN( u1_uk_n117 ) , .A( u1_uk_n277 ) );
  INV_X1 u1_uk_U231 (.ZN( u1_K10_39 ) , .A( u1_uk_n373 ) );
  AOI22_X1 u1_uk_U232 (.B2( u1_uk_K_r8_44 ) , .A2( u1_uk_K_r8_52 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n209 ) , .ZN( u1_uk_n373 ) );
  OAI21_X1 u1_uk_U234 (.ZN( u1_K10_31 ) , .B2( u1_uk_n1645 ) , .B1( u1_uk_n298 ) , .A( u1_uk_n342 ) );
  NAND2_X1 u1_uk_U235 (.A1( u1_uk_K_r8_16 ) , .A2( u1_uk_n277 ) , .ZN( u1_uk_n342 ) );
  OAI21_X1 u1_uk_U249 (.ZN( u1_K12_39 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1720 ) , .A( u1_uk_n590 ) );
  NAND2_X1 u1_uk_U250 (.A1( u1_uk_K_r10_16 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n590 ) );
  OAI21_X1 u1_uk_U254 (.ZN( u1_K8_44 ) , .A( u1_uk_n1144 ) , .B1( u1_uk_n141 ) , .B2( u1_uk_n1568 ) );
  NAND2_X1 u1_uk_U255 (.A1( u1_uk_K_r6_0 ) , .ZN( u1_uk_n1144 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U256 (.ZN( u1_K8_48 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1534 ) , .B2( u1_uk_n1541 ) , .B1( u1_uk_n220 ) );
  INV_X1 u1_uk_U270 (.ZN( u1_K12_44 ) , .A( u1_uk_n608 ) );
  AOI22_X1 u1_uk_U271 (.B2( u1_uk_K_r10_37 ) , .A2( u1_uk_K_r10_42 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n271 ) , .ZN( u1_uk_n608 ) );
  OAI22_X1 u1_uk_U272 (.ZN( u1_K12_48 ) , .B2( u1_uk_n1721 ) , .A2( u1_uk_n1730 ) , .B1( u1_uk_n207 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U282 (.ZN( u1_K4_44 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1350 ) , .A2( u1_uk_n1367 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U287 (.ZN( u1_K16_6 ) , .B2( u1_uk_n1244 ) , .A2( u1_uk_n1249 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U295 (.ZN( u1_K4_6 ) , .A( u1_uk_n1069 ) , .B2( u1_uk_n1365 ) , .B1( u1_uk_n83 ) );
  NAND2_X1 u1_uk_U296 (.A1( u1_uk_K_r2_24 ) , .ZN( u1_uk_n1069 ) , .A2( u1_uk_n145 ) );
  OAI22_X1 u1_uk_U314 (.ZN( u1_K16_8 ) , .A2( u1_uk_n1221 ) , .B2( u1_uk_n1234 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U338 (.ZN( u1_K12_46 ) , .B2( u1_uk_n1708 ) , .A2( u1_uk_n1748 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U339 (.ZN( u1_K4_46 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1360 ) , .A2( u1_uk_n1374 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U347 (.ZN( u1_K14_4 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1816 ) , .A2( u1_uk_n1824 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U353 (.ZN( u1_K4_4 ) , .A( u1_uk_n1067 ) );
  AOI22_X1 u1_uk_U354 (.B2( u1_uk_K_r2_13 ) , .A2( u1_uk_K_r2_18 ) , .ZN( u1_uk_n1067 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U371 (.ZN( u1_K10_40 ) , .A( u1_uk_n375 ) );
  AOI22_X1 u1_uk_U372 (.A2( u1_uk_K_r8_2 ) , .B2( u1_uk_K_r8_22 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n250 ) , .ZN( u1_uk_n375 ) );
  OAI22_X1 u1_uk_U396 (.ZN( u1_K14_1 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1808 ) , .A2( u1_uk_n1813 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U412 (.ZN( u1_K4_16 ) , .B2( u1_uk_n1359 ) , .A2( u1_uk_n1363 ) , .B1( u1_uk_n145 ) , .A1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U418 (.ZN( u1_K14_9 ) , .B2( u1_uk_n1818 ) , .B1( u1_uk_n83 ) , .A( u1_uk_n963 ) );
  NAND2_X1 u1_uk_U419 (.A1( u1_uk_K_r12_18 ) , .ZN( u1_uk_n963 ) , .A2( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U429 (.ZN( u1_K16_9 ) , .B2( u1_uk_n1251 ) , .A2( u1_uk_n1258 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U430 (.ZN( u1_K12_33 ) , .B2( u1_uk_n1748 ) , .A( u1_uk_n586 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U431 (.A1( u1_uk_K_r10_14 ) , .A2( u1_uk_n117 ) , .ZN( u1_uk_n586 ) );
  INV_X1 u1_uk_U441 (.ZN( u1_K10_37 ) , .A( u1_uk_n366 ) );
  AOI22_X1 u1_uk_U442 (.B2( u1_uk_K_r8_28 ) , .A2( u1_uk_K_r8_52 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n208 ) , .ZN( u1_uk_n366 ) );
  INV_X1 u1_uk_U463 (.ZN( u1_K10_33 ) , .A( u1_uk_n349 ) );
  AOI22_X1 u1_uk_U464 (.B2( u1_uk_K_r8_22 ) , .A2( u1_uk_K_r8_42 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n297 ) , .ZN( u1_uk_n349 ) );
  OAI22_X1 u1_uk_U472 (.ZN( u1_K12_37 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1709 ) , .A2( u1_uk_n1749 ) , .A1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U481 (.ZN( u1_K10_36 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1619 ) , .A( u1_uk_n363 ) );
  NAND2_X1 u1_uk_U482 (.A1( u1_uk_K_r8_21 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n363 ) );
  OAI22_X1 u1_uk_U505 (.ZN( u1_K14_2 ) , .A1( u1_uk_n182 ) , .B2( u1_uk_n1824 ) , .A2( u1_uk_n1831 ) , .B1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U526 (.ZN( u1_K4_17 ) , .A( u1_uk_n1051 ) , .B2( u1_uk_n1369 ) , .B1( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U527 (.A1( u1_uk_K_r2_27 ) , .ZN( u1_uk_n1051 ) , .A2( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U530 (.ZN( u1_K14_12 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1831 ) , .A2( u1_uk_n1835 ) , .B1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U546 (.ZN( u1_K16_12 ) , .B2( u1_uk_n1228 ) , .B1( u1_uk_n223 ) , .A( u1_uk_n979 ) );
  NAND2_X1 u1_uk_U547 (.A1( u1_uk_K_r14_12 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n979 ) );
  OAI22_X1 u1_uk_U552 (.ZN( u1_K14_17 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1810 ) , .A2( u1_uk_n1834 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U563 (.ZN( u1_K12_38 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1708 ) , .A2( u1_uk_n1735 ) , .B1( u1_uk_n209 ) );
  INV_X1 u1_uk_U574 (.ZN( u1_K10_38 ) , .A( u1_uk_n369 ) );
  AOI22_X1 u1_uk_U575 (.B2( u1_uk_K_r8_28 ) , .A2( u1_uk_K_r8_8 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n369 ) );
  OAI22_X1 u1_uk_U579 (.ZN( u1_K16_10 ) , .B2( u1_uk_n1249 ) , .A2( u1_uk_n1252 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U582 (.ZN( u1_K14_10 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1809 ) , .A2( u1_uk_n1814 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U596 (.ZN( u1_K16_22 ) , .B2( u1_uk_n1235 ) , .A2( u1_uk_n1242 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U619 (.ZN( u1_K12_35 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1728 ) , .A2( u1_uk_n1737 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U622 (.ZN( u1_K10_35 ) , .A( u1_uk_n353 ) );
  AOI22_X1 u1_uk_U623 (.B2( u1_uk_K_r8_2 ) , .A2( u1_uk_K_r8_37 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n252 ) , .ZN( u1_uk_n353 ) );
  OAI21_X1 u1_uk_U633 (.ZN( u1_K16_11 ) , .B2( u1_uk_n1242 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n978 ) );
  NAND2_X1 u1_uk_U634 (.A1( u1_uk_K_r14_39 ) , .A2( u1_uk_n94 ) , .ZN( u1_uk_n978 ) );
  OAI22_X1 u1_uk_U637 (.ZN( u1_K14_11 ) , .A2( u1_uk_n1801 ) , .B2( u1_uk_n1808 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n99 ) );
  INV_X1 u1_uk_U650 (.ZN( u1_K4_23 ) , .A( u1_uk_n1056 ) );
  AOI22_X1 u1_uk_U651 (.B2( u1_uk_K_r2_18 ) , .A2( u1_uk_K_r2_55 ) , .ZN( u1_uk_n1056 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n251 ) );
  OAI21_X1 u1_uk_U656 (.ZN( u1_K4_43 ) , .A( u1_uk_n1066 ) , .B2( u1_uk_n1389 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U657 (.A1( u1_uk_K_r2_29 ) , .ZN( u1_uk_n1066 ) , .A2( u1_uk_n128 ) );
  OAI21_X1 u1_uk_U673 (.ZN( u1_K12_45 ) , .B2( u1_uk_n1714 ) , .B1( u1_uk_n191 ) , .A( u1_uk_n634 ) );
  NAND2_X1 u1_uk_U674 (.A1( u1_uk_K_r10_43 ) , .A2( u1_uk_n214 ) , .ZN( u1_uk_n634 ) );
  INV_X1 u1_uk_U698 (.ZN( u1_K8_43 ) , .A( u1_uk_n1143 ) );
  AOI22_X1 u1_uk_U699 (.B2( u1_uk_K_r6_21 ) , .A2( u1_uk_K_r6_28 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1143 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U700 (.ZN( u1_K16_3 ) , .B2( u1_uk_n1228 ) , .A2( u1_uk_n1236 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U702 (.ZN( u1_K16_7 ) , .B2( u1_uk_n1229 ) , .A2( u1_uk_n1237 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U707 (.ZN( u1_K4_3 ) , .A( u1_uk_n1065 ) );
  AOI22_X1 u1_uk_U708 (.A2( u1_uk_K_r2_4 ) , .B2( u1_uk_K_r2_41 ) , .ZN( u1_uk_n1065 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U736 (.ZN( u1_K10_42 ) , .B2( u1_uk_n1619 ) , .A1( u1_uk_n162 ) , .A2( u1_uk_n1645 ) , .B1( u1_uk_n291 ) );
  INV_X1 u1_uk_U740 (.ZN( u1_K12_42 ) , .A( u1_uk_n605 ) );
  AOI22_X1 u1_uk_U741 (.B2( u1_uk_K_r10_28 ) , .A2( u1_uk_K_r10_9 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n294 ) , .ZN( u1_uk_n605 ) );
  OAI22_X1 u1_uk_U773 (.ZN( u1_K4_21 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1371 ) , .A2( u1_uk_n1377 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U775 (.ZN( u1_K14_13 ) , .B2( u1_uk_n1812 ) , .A2( u1_uk_n1817 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U778 (.ZN( u1_K4_13 ) , .A2( u1_uk_n1354 ) , .B2( u1_uk_n1358 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U78 (.ZN( u1_K12_34 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1715 ) , .B2( u1_uk_n1730 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U802 (.ZN( u1_K16_1 ) , .B2( u1_uk_n1248 ) , .A2( u1_uk_n1251 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U808 (.ZN( u1_K4_1 ) , .A( u1_uk_n1053 ) , .B2( u1_uk_n1353 ) , .B1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U809 (.A1( u1_uk_K_r2_25 ) , .ZN( u1_uk_n1053 ) , .A2( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U810 (.ZN( u1_K4_18 ) , .A( u1_uk_n1052 ) , .B2( u1_uk_n1378 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U811 (.A1( u1_uk_K_r2_20 ) , .ZN( u1_uk_n1052 ) , .A2( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U828 (.ZN( u1_K16_20 ) , .B2( u1_uk_n1252 ) , .A2( u1_uk_n1259 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U841 (.ZN( u1_K4_22 ) , .A( u1_uk_n1055 ) , .B2( u1_uk_n1357 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U842 (.A1( u1_uk_K_r2_47 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n1055 ) );
  OAI22_X1 u1_uk_U85 (.ZN( u1_K16_23 ) , .B2( u1_uk_n1243 ) , .A2( u1_uk_n1248 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI21_X1 u1_uk_U853 (.ZN( u1_K14_3 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1842 ) , .A( u1_uk_n957 ) );
  NAND2_X1 u1_uk_U854 (.A1( u1_uk_K_r12_47 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n957 ) );
  OAI21_X1 u1_uk_U857 (.ZN( u1_K16_2 ) , .B2( u1_uk_n1220 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n986 ) );
  NAND2_X1 u1_uk_U858 (.A1( u1_uk_K_r14_11 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n986 ) );
  AOI22_X1 u1_uk_U860 (.B2( u1_uk_K_r2_26 ) , .A2( u1_uk_K_r2_46 ) , .ZN( u1_uk_n1061 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U887 (.ZN( u1_K12_43 ) , .B2( u1_uk_n1717 ) , .A2( u1_uk_n1737 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U891 (.ZN( u1_K14_6 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1803 ) , .B2( u1_uk_n1810 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U898 (.ZN( u1_K14_7 ) , .B2( u1_uk_n1816 ) , .A2( u1_uk_n1835 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U907 (.ZN( u1_K16_21 ) , .B2( u1_uk_n1227 ) , .A2( u1_uk_n1234 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U909 (.ZN( u1_K16_24 ) , .B2( u1_uk_n1224 ) , .A2( u1_uk_n1229 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U913 (.ZN( u1_K4_14 ) , .B1( u1_uk_n110 ) , .B2( u1_uk_n1352 ) , .A2( u1_uk_n1378 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U937 (.ZN( u1_K14_8 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1801 ) , .B2( u1_uk_n1819 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U942 (.ZN( u1_K14_14 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1834 ) , .A2( u1_uk_n1841 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U948 (.ZN( u1_K10_34 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1618 ) , .A2( u1_uk_n1644 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U953 (.ZN( u1_K4_48 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1355 ) , .B2( u1_uk_n1383 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U959 (.ZN( u1_K14_18 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1818 ) , .A2( u1_uk_n1826 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U961 (.ZN( u1_K16_19 ) , .B2( u1_uk_n1220 ) , .A2( u1_uk_n1258 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U964 (.ZN( u1_K14_16 ) , .A1( u1_uk_n142 ) , .A2( u1_uk_n1804 ) , .B2( u1_uk_n1842 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U974 (.ZN( u1_K8_45 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1528 ) , .A2( u1_uk_n1566 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U978 (.ZN( u1_K4_45 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1351 ) , .A2( u1_uk_n1390 ) , .B1( u1_uk_n242 ) );
  XOR2_X1 u2_U343 (.B( u2_L5_32 ) , .Z( u2_N223 ) , .A( u2_out6_32 ) );
  XOR2_X1 u2_U346 (.B( u2_L5_29 ) , .Z( u2_N220 ) , .A( u2_out6_29 ) );
  XOR2_X1 u2_U349 (.B( u2_L5_27 ) , .Z( u2_N218 ) , .A( u2_out6_27 ) );
  XOR2_X1 u2_U351 (.B( u2_L5_25 ) , .Z( u2_N216 ) , .A( u2_out6_25 ) );
  XOR2_X1 u2_U354 (.B( u2_L5_22 ) , .Z( u2_N213 ) , .A( u2_out6_22 ) );
  XOR2_X1 u2_U355 (.B( u2_L5_21 ) , .Z( u2_N212 ) , .A( u2_out6_21 ) );
  XOR2_X1 u2_U357 (.B( u2_L5_19 ) , .Z( u2_N210 ) , .A( u2_out6_19 ) );
  XOR2_X1 u2_U362 (.B( u2_L5_15 ) , .Z( u2_N206 ) , .A( u2_out6_15 ) );
  XOR2_X1 u2_U363 (.B( u2_L5_14 ) , .Z( u2_N205 ) , .A( u2_out6_14 ) );
  XOR2_X1 u2_U365 (.B( u2_L5_12 ) , .Z( u2_N203 ) , .A( u2_out6_12 ) );
  XOR2_X1 u2_U366 (.B( u2_L5_11 ) , .Z( u2_N202 ) , .A( u2_out6_11 ) );
  XOR2_X1 u2_U371 (.B( u2_L5_8 ) , .Z( u2_N199 ) , .A( u2_out6_8 ) );
  XOR2_X1 u2_U372 (.B( u2_L5_7 ) , .Z( u2_N198 ) , .A( u2_out6_7 ) );
  XOR2_X1 u2_U374 (.B( u2_L5_5 ) , .Z( u2_N196 ) , .A( u2_out6_5 ) );
  XOR2_X1 u2_U375 (.B( u2_L5_4 ) , .Z( u2_N195 ) , .A( u2_out6_4 ) );
  XOR2_X1 u2_U376 (.B( u2_L5_3 ) , .Z( u2_N194 ) , .A( u2_out6_3 ) );
  XOR2_X1 u2_U485 (.Z( u2_FP_7 ) , .B( u2_L14_7 ) , .A( u2_out15_7 ) );
  XOR2_X1 u2_U488 (.Z( u2_FP_4 ) , .B( u2_L14_4 ) , .A( u2_out15_4 ) );
  XOR2_X1 u2_U490 (.Z( u2_FP_32 ) , .B( u2_L14_32 ) , .A( u2_out15_32 ) );
  XOR2_X1 u2_U494 (.Z( u2_FP_29 ) , .B( u2_L14_29 ) , .A( u2_out15_29 ) );
  XOR2_X1 u2_U501 (.Z( u2_FP_22 ) , .B( u2_L14_22 ) , .A( u2_out15_22 ) );
  XOR2_X1 u2_U505 (.Z( u2_FP_19 ) , .B( u2_L14_19 ) , .A( u2_out15_19 ) );
  XOR2_X1 u2_U512 (.Z( u2_FP_12 ) , .B( u2_L14_12 ) , .A( u2_out15_12 ) );
  XOR2_X1 u2_U513 (.Z( u2_FP_11 ) , .B( u2_L14_11 ) , .A( u2_out15_11 ) );
  XOR2_X1 u2_u15_U13 (.A( u2_FP_61 ) , .B( u2_K16_42 ) , .Z( u2_u15_X_42 ) );
  XOR2_X1 u2_u15_U14 (.A( u2_FP_60 ) , .B( u2_K16_41 ) , .Z( u2_u15_X_41 ) );
  XOR2_X1 u2_u15_U15 (.A( u2_FP_59 ) , .B( u2_K16_40 ) , .Z( u2_u15_X_40 ) );
  XOR2_X1 u2_u15_U17 (.A( u2_FP_58 ) , .B( u2_K16_39 ) , .Z( u2_u15_X_39 ) );
  XOR2_X1 u2_u15_U18 (.A( u2_FP_57 ) , .B( u2_K16_38 ) , .Z( u2_u15_X_38 ) );
  XOR2_X1 u2_u15_U19 (.A( u2_FP_56 ) , .B( u2_K16_37 ) , .Z( u2_u15_X_37 ) );
  XOR2_X1 u2_u15_U20 (.A( u2_FP_57 ) , .B( u2_K16_36 ) , .Z( u2_u15_X_36 ) );
  XOR2_X1 u2_u15_U21 (.A( u2_FP_56 ) , .B( u2_K16_35 ) , .Z( u2_u15_X_35 ) );
  XOR2_X1 u2_u15_U22 (.A( u2_FP_55 ) , .B( u2_K16_34 ) , .Z( u2_u15_X_34 ) );
  XOR2_X1 u2_u15_U23 (.A( u2_FP_54 ) , .B( u2_K16_33 ) , .Z( u2_u15_X_33 ) );
  XOR2_X1 u2_u15_U24 (.A( u2_FP_53 ) , .B( u2_K16_32 ) , .Z( u2_u15_X_32 ) );
  XOR2_X1 u2_u15_U25 (.A( u2_FP_52 ) , .B( u2_K16_31 ) , .Z( u2_u15_X_31 ) );
  INV_X1 u2_u15_u5_U10 (.A( u2_u15_u5_n121 ) , .ZN( u2_u15_u5_n177 ) );
  AOI222_X1 u2_u15_u5_U100 (.ZN( u2_u15_u5_n113 ) , .A1( u2_u15_u5_n131 ) , .C1( u2_u15_u5_n148 ) , .B2( u2_u15_u5_n174 ) , .C2( u2_u15_u5_n178 ) , .A2( u2_u15_u5_n179 ) , .B1( u2_u15_u5_n99 ) );
  NAND4_X1 u2_u15_u5_U101 (.ZN( u2_out15_29 ) , .A4( u2_u15_u5_n129 ) , .A3( u2_u15_u5_n130 ) , .A2( u2_u15_u5_n168 ) , .A1( u2_u15_u5_n196 ) );
  AOI221_X1 u2_u15_u5_U102 (.A( u2_u15_u5_n128 ) , .ZN( u2_u15_u5_n129 ) , .C2( u2_u15_u5_n132 ) , .B2( u2_u15_u5_n159 ) , .B1( u2_u15_u5_n176 ) , .C1( u2_u15_u5_n184 ) );
  AOI222_X1 u2_u15_u5_U103 (.ZN( u2_u15_u5_n130 ) , .A2( u2_u15_u5_n146 ) , .B1( u2_u15_u5_n147 ) , .C2( u2_u15_u5_n175 ) , .B2( u2_u15_u5_n179 ) , .A1( u2_u15_u5_n188 ) , .C1( u2_u15_u5_n194 ) );
  NAND3_X1 u2_u15_u5_U104 (.A2( u2_u15_u5_n154 ) , .A3( u2_u15_u5_n158 ) , .A1( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n99 ) );
  NOR2_X1 u2_u15_u5_U11 (.ZN( u2_u15_u5_n160 ) , .A2( u2_u15_u5_n173 ) , .A1( u2_u15_u5_n177 ) );
  INV_X1 u2_u15_u5_U12 (.A( u2_u15_u5_n150 ) , .ZN( u2_u15_u5_n174 ) );
  AOI21_X1 u2_u15_u5_U13 (.A( u2_u15_u5_n160 ) , .B2( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n162 ) , .B1( u2_u15_u5_n192 ) );
  INV_X1 u2_u15_u5_U14 (.A( u2_u15_u5_n159 ) , .ZN( u2_u15_u5_n192 ) );
  AOI21_X1 u2_u15_u5_U15 (.A( u2_u15_u5_n156 ) , .B2( u2_u15_u5_n157 ) , .B1( u2_u15_u5_n158 ) , .ZN( u2_u15_u5_n163 ) );
  AOI21_X1 u2_u15_u5_U16 (.B2( u2_u15_u5_n139 ) , .B1( u2_u15_u5_n140 ) , .ZN( u2_u15_u5_n141 ) , .A( u2_u15_u5_n150 ) );
  OAI21_X1 u2_u15_u5_U17 (.A( u2_u15_u5_n133 ) , .B2( u2_u15_u5_n134 ) , .B1( u2_u15_u5_n135 ) , .ZN( u2_u15_u5_n142 ) );
  OAI21_X1 u2_u15_u5_U18 (.ZN( u2_u15_u5_n133 ) , .B2( u2_u15_u5_n147 ) , .A( u2_u15_u5_n173 ) , .B1( u2_u15_u5_n188 ) );
  NAND2_X1 u2_u15_u5_U19 (.A2( u2_u15_u5_n119 ) , .A1( u2_u15_u5_n123 ) , .ZN( u2_u15_u5_n137 ) );
  INV_X1 u2_u15_u5_U20 (.A( u2_u15_u5_n155 ) , .ZN( u2_u15_u5_n194 ) );
  NAND2_X1 u2_u15_u5_U21 (.A1( u2_u15_u5_n121 ) , .ZN( u2_u15_u5_n132 ) , .A2( u2_u15_u5_n172 ) );
  NAND2_X1 u2_u15_u5_U22 (.A2( u2_u15_u5_n122 ) , .ZN( u2_u15_u5_n136 ) , .A1( u2_u15_u5_n154 ) );
  NAND2_X1 u2_u15_u5_U23 (.A2( u2_u15_u5_n119 ) , .A1( u2_u15_u5_n120 ) , .ZN( u2_u15_u5_n159 ) );
  INV_X1 u2_u15_u5_U24 (.A( u2_u15_u5_n156 ) , .ZN( u2_u15_u5_n175 ) );
  INV_X1 u2_u15_u5_U25 (.A( u2_u15_u5_n158 ) , .ZN( u2_u15_u5_n188 ) );
  INV_X1 u2_u15_u5_U26 (.A( u2_u15_u5_n152 ) , .ZN( u2_u15_u5_n179 ) );
  INV_X1 u2_u15_u5_U27 (.A( u2_u15_u5_n140 ) , .ZN( u2_u15_u5_n182 ) );
  INV_X1 u2_u15_u5_U28 (.A( u2_u15_u5_n151 ) , .ZN( u2_u15_u5_n183 ) );
  INV_X1 u2_u15_u5_U29 (.A( u2_u15_u5_n123 ) , .ZN( u2_u15_u5_n185 ) );
  NOR2_X1 u2_u15_u5_U3 (.ZN( u2_u15_u5_n134 ) , .A1( u2_u15_u5_n183 ) , .A2( u2_u15_u5_n190 ) );
  INV_X1 u2_u15_u5_U30 (.A( u2_u15_u5_n161 ) , .ZN( u2_u15_u5_n184 ) );
  INV_X1 u2_u15_u5_U31 (.A( u2_u15_u5_n139 ) , .ZN( u2_u15_u5_n189 ) );
  INV_X1 u2_u15_u5_U32 (.A( u2_u15_u5_n157 ) , .ZN( u2_u15_u5_n190 ) );
  INV_X1 u2_u15_u5_U33 (.A( u2_u15_u5_n120 ) , .ZN( u2_u15_u5_n193 ) );
  NAND2_X1 u2_u15_u5_U34 (.ZN( u2_u15_u5_n111 ) , .A1( u2_u15_u5_n140 ) , .A2( u2_u15_u5_n155 ) );
  NOR2_X1 u2_u15_u5_U35 (.ZN( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n170 ) , .A2( u2_u15_u5_n180 ) );
  INV_X1 u2_u15_u5_U36 (.A( u2_u15_u5_n117 ) , .ZN( u2_u15_u5_n196 ) );
  OAI221_X1 u2_u15_u5_U37 (.A( u2_u15_u5_n116 ) , .ZN( u2_u15_u5_n117 ) , .B2( u2_u15_u5_n119 ) , .C1( u2_u15_u5_n153 ) , .C2( u2_u15_u5_n158 ) , .B1( u2_u15_u5_n172 ) );
  AOI222_X1 u2_u15_u5_U38 (.ZN( u2_u15_u5_n116 ) , .B2( u2_u15_u5_n145 ) , .C1( u2_u15_u5_n148 ) , .A2( u2_u15_u5_n174 ) , .C2( u2_u15_u5_n177 ) , .B1( u2_u15_u5_n187 ) , .A1( u2_u15_u5_n193 ) );
  INV_X1 u2_u15_u5_U39 (.A( u2_u15_u5_n115 ) , .ZN( u2_u15_u5_n187 ) );
  INV_X1 u2_u15_u5_U4 (.A( u2_u15_u5_n138 ) , .ZN( u2_u15_u5_n191 ) );
  AOI22_X1 u2_u15_u5_U40 (.B2( u2_u15_u5_n131 ) , .A2( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n169 ) , .B1( u2_u15_u5_n174 ) , .A1( u2_u15_u5_n185 ) );
  NOR2_X1 u2_u15_u5_U41 (.A1( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n150 ) , .A2( u2_u15_u5_n173 ) );
  AOI21_X1 u2_u15_u5_U42 (.A( u2_u15_u5_n118 ) , .B2( u2_u15_u5_n145 ) , .ZN( u2_u15_u5_n168 ) , .B1( u2_u15_u5_n186 ) );
  INV_X1 u2_u15_u5_U43 (.A( u2_u15_u5_n122 ) , .ZN( u2_u15_u5_n186 ) );
  NOR2_X1 u2_u15_u5_U44 (.A1( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n152 ) , .A2( u2_u15_u5_n176 ) );
  NOR2_X1 u2_u15_u5_U45 (.A1( u2_u15_u5_n115 ) , .ZN( u2_u15_u5_n118 ) , .A2( u2_u15_u5_n153 ) );
  NOR2_X1 u2_u15_u5_U46 (.A2( u2_u15_u5_n145 ) , .ZN( u2_u15_u5_n156 ) , .A1( u2_u15_u5_n174 ) );
  NOR2_X1 u2_u15_u5_U47 (.ZN( u2_u15_u5_n121 ) , .A2( u2_u15_u5_n145 ) , .A1( u2_u15_u5_n176 ) );
  AOI22_X1 u2_u15_u5_U48 (.ZN( u2_u15_u5_n114 ) , .A2( u2_u15_u5_n137 ) , .A1( u2_u15_u5_n145 ) , .B2( u2_u15_u5_n175 ) , .B1( u2_u15_u5_n193 ) );
  OAI211_X1 u2_u15_u5_U49 (.B( u2_u15_u5_n124 ) , .A( u2_u15_u5_n125 ) , .C2( u2_u15_u5_n126 ) , .C1( u2_u15_u5_n127 ) , .ZN( u2_u15_u5_n128 ) );
  OAI21_X1 u2_u15_u5_U5 (.B2( u2_u15_u5_n136 ) , .B1( u2_u15_u5_n137 ) , .ZN( u2_u15_u5_n138 ) , .A( u2_u15_u5_n177 ) );
  NOR3_X1 u2_u15_u5_U50 (.ZN( u2_u15_u5_n127 ) , .A1( u2_u15_u5_n136 ) , .A3( u2_u15_u5_n148 ) , .A2( u2_u15_u5_n182 ) );
  OAI21_X1 u2_u15_u5_U51 (.ZN( u2_u15_u5_n124 ) , .A( u2_u15_u5_n177 ) , .B2( u2_u15_u5_n183 ) , .B1( u2_u15_u5_n189 ) );
  OAI21_X1 u2_u15_u5_U52 (.ZN( u2_u15_u5_n125 ) , .A( u2_u15_u5_n174 ) , .B2( u2_u15_u5_n185 ) , .B1( u2_u15_u5_n190 ) );
  AOI21_X1 u2_u15_u5_U53 (.A( u2_u15_u5_n153 ) , .B2( u2_u15_u5_n154 ) , .B1( u2_u15_u5_n155 ) , .ZN( u2_u15_u5_n164 ) );
  AOI21_X1 u2_u15_u5_U54 (.ZN( u2_u15_u5_n110 ) , .B1( u2_u15_u5_n122 ) , .B2( u2_u15_u5_n139 ) , .A( u2_u15_u5_n153 ) );
  INV_X1 u2_u15_u5_U55 (.A( u2_u15_u5_n153 ) , .ZN( u2_u15_u5_n176 ) );
  INV_X1 u2_u15_u5_U56 (.A( u2_u15_u5_n126 ) , .ZN( u2_u15_u5_n173 ) );
  AND2_X1 u2_u15_u5_U57 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n147 ) );
  AND2_X1 u2_u15_u5_U58 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n148 ) );
  NAND2_X1 u2_u15_u5_U59 (.A1( u2_u15_u5_n105 ) , .A2( u2_u15_u5_n106 ) , .ZN( u2_u15_u5_n158 ) );
  INV_X1 u2_u15_u5_U6 (.A( u2_u15_u5_n135 ) , .ZN( u2_u15_u5_n178 ) );
  NAND2_X1 u2_u15_u5_U60 (.A2( u2_u15_u5_n108 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n139 ) );
  NAND2_X1 u2_u15_u5_U61 (.A1( u2_u15_u5_n106 ) , .A2( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n119 ) );
  NAND2_X1 u2_u15_u5_U62 (.A2( u2_u15_u5_n103 ) , .A1( u2_u15_u5_n105 ) , .ZN( u2_u15_u5_n140 ) );
  NAND2_X1 u2_u15_u5_U63 (.A2( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n105 ) , .ZN( u2_u15_u5_n155 ) );
  NAND2_X1 u2_u15_u5_U64 (.A2( u2_u15_u5_n106 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n122 ) );
  NAND2_X1 u2_u15_u5_U65 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n106 ) , .ZN( u2_u15_u5_n115 ) );
  NAND2_X1 u2_u15_u5_U66 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n103 ) , .ZN( u2_u15_u5_n161 ) );
  NAND2_X1 u2_u15_u5_U67 (.A1( u2_u15_u5_n105 ) , .A2( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n154 ) );
  INV_X1 u2_u15_u5_U68 (.A( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n172 ) );
  NAND2_X1 u2_u15_u5_U69 (.A1( u2_u15_u5_n103 ) , .A2( u2_u15_u5_n108 ) , .ZN( u2_u15_u5_n123 ) );
  OAI22_X1 u2_u15_u5_U7 (.B2( u2_u15_u5_n149 ) , .B1( u2_u15_u5_n150 ) , .A2( u2_u15_u5_n151 ) , .A1( u2_u15_u5_n152 ) , .ZN( u2_u15_u5_n165 ) );
  NAND2_X1 u2_u15_u5_U70 (.A2( u2_u15_u5_n103 ) , .A1( u2_u15_u5_n107 ) , .ZN( u2_u15_u5_n151 ) );
  NAND2_X1 u2_u15_u5_U71 (.A2( u2_u15_u5_n107 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n120 ) );
  NAND2_X1 u2_u15_u5_U72 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n109 ) , .ZN( u2_u15_u5_n157 ) );
  AND2_X1 u2_u15_u5_U73 (.A2( u2_u15_u5_n100 ) , .A1( u2_u15_u5_n104 ) , .ZN( u2_u15_u5_n131 ) );
  INV_X1 u2_u15_u5_U74 (.A( u2_u15_u5_n102 ) , .ZN( u2_u15_u5_n195 ) );
  OAI221_X1 u2_u15_u5_U75 (.A( u2_u15_u5_n101 ) , .ZN( u2_u15_u5_n102 ) , .C2( u2_u15_u5_n115 ) , .C1( u2_u15_u5_n126 ) , .B1( u2_u15_u5_n134 ) , .B2( u2_u15_u5_n160 ) );
  OAI21_X1 u2_u15_u5_U76 (.ZN( u2_u15_u5_n101 ) , .B1( u2_u15_u5_n137 ) , .A( u2_u15_u5_n146 ) , .B2( u2_u15_u5_n147 ) );
  NOR2_X1 u2_u15_u5_U77 (.A2( u2_u15_X_34 ) , .A1( u2_u15_X_35 ) , .ZN( u2_u15_u5_n145 ) );
  NOR2_X1 u2_u15_u5_U78 (.A2( u2_u15_X_34 ) , .ZN( u2_u15_u5_n146 ) , .A1( u2_u15_u5_n171 ) );
  NOR2_X1 u2_u15_u5_U79 (.A2( u2_u15_X_31 ) , .A1( u2_u15_X_32 ) , .ZN( u2_u15_u5_n103 ) );
  NOR3_X1 u2_u15_u5_U8 (.A2( u2_u15_u5_n147 ) , .A1( u2_u15_u5_n148 ) , .ZN( u2_u15_u5_n149 ) , .A3( u2_u15_u5_n194 ) );
  NOR2_X1 u2_u15_u5_U80 (.A2( u2_u15_X_36 ) , .ZN( u2_u15_u5_n105 ) , .A1( u2_u15_u5_n180 ) );
  NOR2_X1 u2_u15_u5_U81 (.A2( u2_u15_X_33 ) , .ZN( u2_u15_u5_n108 ) , .A1( u2_u15_u5_n170 ) );
  NOR2_X1 u2_u15_u5_U82 (.A2( u2_u15_X_33 ) , .A1( u2_u15_X_36 ) , .ZN( u2_u15_u5_n107 ) );
  NOR2_X1 u2_u15_u5_U83 (.A2( u2_u15_X_31 ) , .ZN( u2_u15_u5_n104 ) , .A1( u2_u15_u5_n181 ) );
  NAND2_X1 u2_u15_u5_U84 (.A2( u2_u15_X_34 ) , .A1( u2_u15_X_35 ) , .ZN( u2_u15_u5_n153 ) );
  NAND2_X1 u2_u15_u5_U85 (.A1( u2_u15_X_34 ) , .ZN( u2_u15_u5_n126 ) , .A2( u2_u15_u5_n171 ) );
  AND2_X1 u2_u15_u5_U86 (.A1( u2_u15_X_31 ) , .A2( u2_u15_X_32 ) , .ZN( u2_u15_u5_n106 ) );
  AND2_X1 u2_u15_u5_U87 (.A1( u2_u15_X_31 ) , .ZN( u2_u15_u5_n109 ) , .A2( u2_u15_u5_n181 ) );
  INV_X1 u2_u15_u5_U88 (.A( u2_u15_X_33 ) , .ZN( u2_u15_u5_n180 ) );
  INV_X1 u2_u15_u5_U89 (.A( u2_u15_X_35 ) , .ZN( u2_u15_u5_n171 ) );
  NOR2_X1 u2_u15_u5_U9 (.ZN( u2_u15_u5_n135 ) , .A1( u2_u15_u5_n173 ) , .A2( u2_u15_u5_n176 ) );
  INV_X1 u2_u15_u5_U90 (.A( u2_u15_X_36 ) , .ZN( u2_u15_u5_n170 ) );
  INV_X1 u2_u15_u5_U91 (.A( u2_u15_X_32 ) , .ZN( u2_u15_u5_n181 ) );
  NAND4_X1 u2_u15_u5_U92 (.ZN( u2_out15_19 ) , .A4( u2_u15_u5_n166 ) , .A3( u2_u15_u5_n167 ) , .A2( u2_u15_u5_n168 ) , .A1( u2_u15_u5_n169 ) );
  AOI22_X1 u2_u15_u5_U93 (.B2( u2_u15_u5_n145 ) , .A2( u2_u15_u5_n146 ) , .ZN( u2_u15_u5_n167 ) , .B1( u2_u15_u5_n182 ) , .A1( u2_u15_u5_n189 ) );
  NOR4_X1 u2_u15_u5_U94 (.A4( u2_u15_u5_n162 ) , .A3( u2_u15_u5_n163 ) , .A2( u2_u15_u5_n164 ) , .A1( u2_u15_u5_n165 ) , .ZN( u2_u15_u5_n166 ) );
  NAND4_X1 u2_u15_u5_U95 (.ZN( u2_out15_11 ) , .A4( u2_u15_u5_n143 ) , .A3( u2_u15_u5_n144 ) , .A2( u2_u15_u5_n169 ) , .A1( u2_u15_u5_n196 ) );
  AOI22_X1 u2_u15_u5_U96 (.A2( u2_u15_u5_n132 ) , .ZN( u2_u15_u5_n144 ) , .B2( u2_u15_u5_n145 ) , .B1( u2_u15_u5_n184 ) , .A1( u2_u15_u5_n194 ) );
  NOR3_X1 u2_u15_u5_U97 (.A3( u2_u15_u5_n141 ) , .A1( u2_u15_u5_n142 ) , .ZN( u2_u15_u5_n143 ) , .A2( u2_u15_u5_n191 ) );
  NAND4_X1 u2_u15_u5_U98 (.ZN( u2_out15_4 ) , .A4( u2_u15_u5_n112 ) , .A2( u2_u15_u5_n113 ) , .A1( u2_u15_u5_n114 ) , .A3( u2_u15_u5_n195 ) );
  AOI211_X1 u2_u15_u5_U99 (.A( u2_u15_u5_n110 ) , .C1( u2_u15_u5_n111 ) , .ZN( u2_u15_u5_n112 ) , .B( u2_u15_u5_n118 ) , .C2( u2_u15_u5_n177 ) );
  INV_X1 u2_u15_u6_U10 (.ZN( u2_u15_u6_n172 ) , .A( u2_u15_u6_n88 ) );
  OAI21_X1 u2_u15_u6_U11 (.A( u2_u15_u6_n159 ) , .B1( u2_u15_u6_n169 ) , .B2( u2_u15_u6_n173 ) , .ZN( u2_u15_u6_n90 ) );
  AOI22_X1 u2_u15_u6_U12 (.A2( u2_u15_u6_n151 ) , .B2( u2_u15_u6_n161 ) , .A1( u2_u15_u6_n167 ) , .B1( u2_u15_u6_n170 ) , .ZN( u2_u15_u6_n89 ) );
  AOI21_X1 u2_u15_u6_U13 (.ZN( u2_u15_u6_n106 ) , .A( u2_u15_u6_n142 ) , .B2( u2_u15_u6_n159 ) , .B1( u2_u15_u6_n164 ) );
  INV_X1 u2_u15_u6_U14 (.A( u2_u15_u6_n155 ) , .ZN( u2_u15_u6_n161 ) );
  INV_X1 u2_u15_u6_U15 (.A( u2_u15_u6_n128 ) , .ZN( u2_u15_u6_n164 ) );
  NAND2_X1 u2_u15_u6_U16 (.ZN( u2_u15_u6_n110 ) , .A1( u2_u15_u6_n122 ) , .A2( u2_u15_u6_n129 ) );
  NAND2_X1 u2_u15_u6_U17 (.ZN( u2_u15_u6_n124 ) , .A2( u2_u15_u6_n146 ) , .A1( u2_u15_u6_n148 ) );
  INV_X1 u2_u15_u6_U18 (.A( u2_u15_u6_n132 ) , .ZN( u2_u15_u6_n171 ) );
  AND2_X1 u2_u15_u6_U19 (.A1( u2_u15_u6_n100 ) , .ZN( u2_u15_u6_n130 ) , .A2( u2_u15_u6_n147 ) );
  INV_X1 u2_u15_u6_U20 (.A( u2_u15_u6_n127 ) , .ZN( u2_u15_u6_n173 ) );
  INV_X1 u2_u15_u6_U21 (.A( u2_u15_u6_n121 ) , .ZN( u2_u15_u6_n167 ) );
  INV_X1 u2_u15_u6_U22 (.A( u2_u15_u6_n100 ) , .ZN( u2_u15_u6_n169 ) );
  INV_X1 u2_u15_u6_U23 (.A( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n170 ) );
  INV_X1 u2_u15_u6_U24 (.A( u2_u15_u6_n113 ) , .ZN( u2_u15_u6_n168 ) );
  AND2_X1 u2_u15_u6_U25 (.A1( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n119 ) , .ZN( u2_u15_u6_n133 ) );
  AND2_X1 u2_u15_u6_U26 (.A2( u2_u15_u6_n121 ) , .A1( u2_u15_u6_n122 ) , .ZN( u2_u15_u6_n131 ) );
  AND3_X1 u2_u15_u6_U27 (.ZN( u2_u15_u6_n120 ) , .A2( u2_u15_u6_n127 ) , .A1( u2_u15_u6_n132 ) , .A3( u2_u15_u6_n145 ) );
  INV_X1 u2_u15_u6_U28 (.A( u2_u15_u6_n146 ) , .ZN( u2_u15_u6_n163 ) );
  AOI222_X1 u2_u15_u6_U29 (.ZN( u2_u15_u6_n114 ) , .A1( u2_u15_u6_n118 ) , .A2( u2_u15_u6_n126 ) , .B2( u2_u15_u6_n151 ) , .C2( u2_u15_u6_n159 ) , .C1( u2_u15_u6_n168 ) , .B1( u2_u15_u6_n169 ) );
  INV_X1 u2_u15_u6_U3 (.A( u2_u15_u6_n110 ) , .ZN( u2_u15_u6_n166 ) );
  NOR2_X1 u2_u15_u6_U30 (.A1( u2_u15_u6_n162 ) , .A2( u2_u15_u6_n165 ) , .ZN( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U31 (.A1( u2_u15_u6_n144 ) , .ZN( u2_u15_u6_n151 ) , .A2( u2_u15_u6_n158 ) );
  NAND2_X1 u2_u15_u6_U32 (.ZN( u2_u15_u6_n132 ) , .A1( u2_u15_u6_n91 ) , .A2( u2_u15_u6_n97 ) );
  AOI22_X1 u2_u15_u6_U33 (.B2( u2_u15_u6_n110 ) , .B1( u2_u15_u6_n111 ) , .A1( u2_u15_u6_n112 ) , .ZN( u2_u15_u6_n115 ) , .A2( u2_u15_u6_n161 ) );
  NAND4_X1 u2_u15_u6_U34 (.A3( u2_u15_u6_n109 ) , .ZN( u2_u15_u6_n112 ) , .A4( u2_u15_u6_n132 ) , .A2( u2_u15_u6_n147 ) , .A1( u2_u15_u6_n166 ) );
  NOR2_X1 u2_u15_u6_U35 (.ZN( u2_u15_u6_n109 ) , .A1( u2_u15_u6_n170 ) , .A2( u2_u15_u6_n173 ) );
  NOR2_X1 u2_u15_u6_U36 (.A2( u2_u15_u6_n126 ) , .ZN( u2_u15_u6_n155 ) , .A1( u2_u15_u6_n160 ) );
  NAND2_X1 u2_u15_u6_U37 (.ZN( u2_u15_u6_n146 ) , .A2( u2_u15_u6_n94 ) , .A1( u2_u15_u6_n99 ) );
  AOI21_X1 u2_u15_u6_U38 (.A( u2_u15_u6_n144 ) , .B2( u2_u15_u6_n145 ) , .B1( u2_u15_u6_n146 ) , .ZN( u2_u15_u6_n150 ) );
  AOI211_X1 u2_u15_u6_U39 (.B( u2_u15_u6_n134 ) , .A( u2_u15_u6_n135 ) , .C1( u2_u15_u6_n136 ) , .ZN( u2_u15_u6_n137 ) , .C2( u2_u15_u6_n151 ) );
  INV_X1 u2_u15_u6_U4 (.A( u2_u15_u6_n142 ) , .ZN( u2_u15_u6_n174 ) );
  NAND4_X1 u2_u15_u6_U40 (.A4( u2_u15_u6_n127 ) , .A3( u2_u15_u6_n128 ) , .A2( u2_u15_u6_n129 ) , .A1( u2_u15_u6_n130 ) , .ZN( u2_u15_u6_n136 ) );
  AOI21_X1 u2_u15_u6_U41 (.B2( u2_u15_u6_n132 ) , .B1( u2_u15_u6_n133 ) , .ZN( u2_u15_u6_n134 ) , .A( u2_u15_u6_n158 ) );
  AOI21_X1 u2_u15_u6_U42 (.B1( u2_u15_u6_n131 ) , .ZN( u2_u15_u6_n135 ) , .A( u2_u15_u6_n144 ) , .B2( u2_u15_u6_n146 ) );
  INV_X1 u2_u15_u6_U43 (.A( u2_u15_u6_n111 ) , .ZN( u2_u15_u6_n158 ) );
  NAND2_X1 u2_u15_u6_U44 (.ZN( u2_u15_u6_n127 ) , .A1( u2_u15_u6_n91 ) , .A2( u2_u15_u6_n92 ) );
  NAND2_X1 u2_u15_u6_U45 (.ZN( u2_u15_u6_n129 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n96 ) );
  INV_X1 u2_u15_u6_U46 (.A( u2_u15_u6_n144 ) , .ZN( u2_u15_u6_n159 ) );
  NAND2_X1 u2_u15_u6_U47 (.ZN( u2_u15_u6_n145 ) , .A2( u2_u15_u6_n97 ) , .A1( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U48 (.ZN( u2_u15_u6_n148 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n94 ) );
  NAND2_X1 u2_u15_u6_U49 (.ZN( u2_u15_u6_n108 ) , .A2( u2_u15_u6_n139 ) , .A1( u2_u15_u6_n144 ) );
  NAND2_X1 u2_u15_u6_U5 (.A2( u2_u15_u6_n143 ) , .ZN( u2_u15_u6_n152 ) , .A1( u2_u15_u6_n166 ) );
  NAND2_X1 u2_u15_u6_U50 (.ZN( u2_u15_u6_n121 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n97 ) );
  NAND2_X1 u2_u15_u6_U51 (.ZN( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n95 ) );
  AND2_X1 u2_u15_u6_U52 (.ZN( u2_u15_u6_n118 ) , .A2( u2_u15_u6_n91 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U53 (.ZN( u2_u15_u6_n147 ) , .A2( u2_u15_u6_n98 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U54 (.ZN( u2_u15_u6_n128 ) , .A1( u2_u15_u6_n94 ) , .A2( u2_u15_u6_n96 ) );
  NAND2_X1 u2_u15_u6_U55 (.ZN( u2_u15_u6_n119 ) , .A2( u2_u15_u6_n95 ) , .A1( u2_u15_u6_n99 ) );
  NAND2_X1 u2_u15_u6_U56 (.ZN( u2_u15_u6_n123 ) , .A2( u2_u15_u6_n91 ) , .A1( u2_u15_u6_n96 ) );
  NAND2_X1 u2_u15_u6_U57 (.ZN( u2_u15_u6_n100 ) , .A2( u2_u15_u6_n92 ) , .A1( u2_u15_u6_n98 ) );
  NAND2_X1 u2_u15_u6_U58 (.ZN( u2_u15_u6_n122 ) , .A1( u2_u15_u6_n94 ) , .A2( u2_u15_u6_n97 ) );
  INV_X1 u2_u15_u6_U59 (.A( u2_u15_u6_n139 ) , .ZN( u2_u15_u6_n160 ) );
  AOI22_X1 u2_u15_u6_U6 (.B2( u2_u15_u6_n101 ) , .A1( u2_u15_u6_n102 ) , .ZN( u2_u15_u6_n103 ) , .B1( u2_u15_u6_n160 ) , .A2( u2_u15_u6_n161 ) );
  NAND2_X1 u2_u15_u6_U60 (.ZN( u2_u15_u6_n113 ) , .A1( u2_u15_u6_n96 ) , .A2( u2_u15_u6_n98 ) );
  NOR2_X1 u2_u15_u6_U61 (.A2( u2_u15_X_40 ) , .A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n126 ) );
  NOR2_X1 u2_u15_u6_U62 (.A2( u2_u15_X_39 ) , .A1( u2_u15_X_42 ) , .ZN( u2_u15_u6_n92 ) );
  NOR2_X1 u2_u15_u6_U63 (.A2( u2_u15_X_39 ) , .A1( u2_u15_u6_n156 ) , .ZN( u2_u15_u6_n97 ) );
  NOR2_X1 u2_u15_u6_U64 (.A2( u2_u15_X_38 ) , .A1( u2_u15_u6_n165 ) , .ZN( u2_u15_u6_n95 ) );
  NOR2_X1 u2_u15_u6_U65 (.A2( u2_u15_X_41 ) , .ZN( u2_u15_u6_n111 ) , .A1( u2_u15_u6_n157 ) );
  NOR2_X1 u2_u15_u6_U66 (.A2( u2_u15_X_37 ) , .A1( u2_u15_u6_n162 ) , .ZN( u2_u15_u6_n94 ) );
  NOR2_X1 u2_u15_u6_U67 (.A2( u2_u15_X_37 ) , .A1( u2_u15_X_38 ) , .ZN( u2_u15_u6_n91 ) );
  NAND2_X1 u2_u15_u6_U68 (.A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n144 ) , .A2( u2_u15_u6_n157 ) );
  NAND2_X1 u2_u15_u6_U69 (.A2( u2_u15_X_40 ) , .A1( u2_u15_X_41 ) , .ZN( u2_u15_u6_n139 ) );
  NOR2_X1 u2_u15_u6_U7 (.A1( u2_u15_u6_n118 ) , .ZN( u2_u15_u6_n143 ) , .A2( u2_u15_u6_n168 ) );
  AND2_X1 u2_u15_u6_U70 (.A1( u2_u15_X_39 ) , .A2( u2_u15_u6_n156 ) , .ZN( u2_u15_u6_n96 ) );
  AND2_X1 u2_u15_u6_U71 (.A1( u2_u15_X_39 ) , .A2( u2_u15_X_42 ) , .ZN( u2_u15_u6_n99 ) );
  INV_X1 u2_u15_u6_U72 (.A( u2_u15_X_40 ) , .ZN( u2_u15_u6_n157 ) );
  INV_X1 u2_u15_u6_U73 (.A( u2_u15_X_37 ) , .ZN( u2_u15_u6_n165 ) );
  INV_X1 u2_u15_u6_U74 (.A( u2_u15_X_38 ) , .ZN( u2_u15_u6_n162 ) );
  INV_X1 u2_u15_u6_U75 (.A( u2_u15_X_42 ) , .ZN( u2_u15_u6_n156 ) );
  NAND4_X1 u2_u15_u6_U76 (.ZN( u2_out15_12 ) , .A4( u2_u15_u6_n114 ) , .A3( u2_u15_u6_n115 ) , .A2( u2_u15_u6_n116 ) , .A1( u2_u15_u6_n117 ) );
  OAI22_X1 u2_u15_u6_U77 (.B2( u2_u15_u6_n111 ) , .ZN( u2_u15_u6_n116 ) , .B1( u2_u15_u6_n126 ) , .A2( u2_u15_u6_n164 ) , .A1( u2_u15_u6_n167 ) );
  OAI21_X1 u2_u15_u6_U78 (.A( u2_u15_u6_n108 ) , .ZN( u2_u15_u6_n117 ) , .B2( u2_u15_u6_n141 ) , .B1( u2_u15_u6_n163 ) );
  NAND4_X1 u2_u15_u6_U79 (.ZN( u2_out15_32 ) , .A4( u2_u15_u6_n103 ) , .A3( u2_u15_u6_n104 ) , .A2( u2_u15_u6_n105 ) , .A1( u2_u15_u6_n106 ) );
  AOI21_X1 u2_u15_u6_U8 (.B1( u2_u15_u6_n107 ) , .B2( u2_u15_u6_n132 ) , .A( u2_u15_u6_n158 ) , .ZN( u2_u15_u6_n88 ) );
  AOI22_X1 u2_u15_u6_U80 (.ZN( u2_u15_u6_n105 ) , .A2( u2_u15_u6_n108 ) , .A1( u2_u15_u6_n118 ) , .B2( u2_u15_u6_n126 ) , .B1( u2_u15_u6_n171 ) );
  AOI22_X1 u2_u15_u6_U81 (.ZN( u2_u15_u6_n104 ) , .A1( u2_u15_u6_n111 ) , .B1( u2_u15_u6_n124 ) , .B2( u2_u15_u6_n151 ) , .A2( u2_u15_u6_n93 ) );
  OAI211_X1 u2_u15_u6_U82 (.ZN( u2_out15_22 ) , .B( u2_u15_u6_n137 ) , .A( u2_u15_u6_n138 ) , .C2( u2_u15_u6_n139 ) , .C1( u2_u15_u6_n140 ) );
  AOI22_X1 u2_u15_u6_U83 (.B1( u2_u15_u6_n124 ) , .A2( u2_u15_u6_n125 ) , .A1( u2_u15_u6_n126 ) , .ZN( u2_u15_u6_n138 ) , .B2( u2_u15_u6_n161 ) );
  AND4_X1 u2_u15_u6_U84 (.A3( u2_u15_u6_n119 ) , .A1( u2_u15_u6_n120 ) , .A4( u2_u15_u6_n129 ) , .ZN( u2_u15_u6_n140 ) , .A2( u2_u15_u6_n143 ) );
  OAI211_X1 u2_u15_u6_U85 (.ZN( u2_out15_7 ) , .B( u2_u15_u6_n153 ) , .C2( u2_u15_u6_n154 ) , .C1( u2_u15_u6_n155 ) , .A( u2_u15_u6_n174 ) );
  NOR3_X1 u2_u15_u6_U86 (.A1( u2_u15_u6_n141 ) , .ZN( u2_u15_u6_n154 ) , .A3( u2_u15_u6_n164 ) , .A2( u2_u15_u6_n171 ) );
  AOI211_X1 u2_u15_u6_U87 (.B( u2_u15_u6_n149 ) , .A( u2_u15_u6_n150 ) , .C2( u2_u15_u6_n151 ) , .C1( u2_u15_u6_n152 ) , .ZN( u2_u15_u6_n153 ) );
  NAND3_X1 u2_u15_u6_U88 (.A2( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n125 ) , .A1( u2_u15_u6_n130 ) , .A3( u2_u15_u6_n131 ) );
  NAND3_X1 u2_u15_u6_U89 (.A3( u2_u15_u6_n133 ) , .ZN( u2_u15_u6_n141 ) , .A1( u2_u15_u6_n145 ) , .A2( u2_u15_u6_n148 ) );
  AOI21_X1 u2_u15_u6_U9 (.B2( u2_u15_u6_n147 ) , .B1( u2_u15_u6_n148 ) , .ZN( u2_u15_u6_n149 ) , .A( u2_u15_u6_n158 ) );
  NAND3_X1 u2_u15_u6_U90 (.ZN( u2_u15_u6_n101 ) , .A3( u2_u15_u6_n107 ) , .A2( u2_u15_u6_n121 ) , .A1( u2_u15_u6_n127 ) );
  NAND3_X1 u2_u15_u6_U91 (.ZN( u2_u15_u6_n102 ) , .A3( u2_u15_u6_n130 ) , .A2( u2_u15_u6_n145 ) , .A1( u2_u15_u6_n166 ) );
  NAND3_X1 u2_u15_u6_U92 (.A3( u2_u15_u6_n113 ) , .A1( u2_u15_u6_n119 ) , .A2( u2_u15_u6_n123 ) , .ZN( u2_u15_u6_n93 ) );
  NAND3_X1 u2_u15_u6_U93 (.ZN( u2_u15_u6_n142 ) , .A2( u2_u15_u6_n172 ) , .A3( u2_u15_u6_n89 ) , .A1( u2_u15_u6_n90 ) );
  XOR2_X1 u2_u6_U10 (.B( u2_K7_45 ) , .A( u2_R5_30 ) , .Z( u2_u6_X_45 ) );
  XOR2_X1 u2_u6_U11 (.B( u2_K7_44 ) , .A( u2_R5_29 ) , .Z( u2_u6_X_44 ) );
  XOR2_X1 u2_u6_U12 (.B( u2_K7_43 ) , .A( u2_R5_28 ) , .Z( u2_u6_X_43 ) );
  XOR2_X1 u2_u6_U13 (.B( u2_K7_42 ) , .A( u2_R5_29 ) , .Z( u2_u6_X_42 ) );
  XOR2_X1 u2_u6_U14 (.B( u2_K7_41 ) , .A( u2_R5_28 ) , .Z( u2_u6_X_41 ) );
  XOR2_X1 u2_u6_U15 (.B( u2_K7_40 ) , .A( u2_R5_27 ) , .Z( u2_u6_X_40 ) );
  XOR2_X1 u2_u6_U17 (.B( u2_K7_39 ) , .A( u2_R5_26 ) , .Z( u2_u6_X_39 ) );
  XOR2_X1 u2_u6_U18 (.B( u2_K7_38 ) , .A( u2_R5_25 ) , .Z( u2_u6_X_38 ) );
  XOR2_X1 u2_u6_U19 (.B( u2_K7_37 ) , .A( u2_R5_24 ) , .Z( u2_u6_X_37 ) );
  XOR2_X1 u2_u6_U20 (.B( u2_K7_36 ) , .A( u2_R5_25 ) , .Z( u2_u6_X_36 ) );
  XOR2_X1 u2_u6_U21 (.B( u2_K7_35 ) , .A( u2_R5_24 ) , .Z( u2_u6_X_35 ) );
  XOR2_X1 u2_u6_U22 (.B( u2_K7_34 ) , .A( u2_R5_23 ) , .Z( u2_u6_X_34 ) );
  XOR2_X1 u2_u6_U23 (.B( u2_K7_33 ) , .A( u2_R5_22 ) , .Z( u2_u6_X_33 ) );
  XOR2_X1 u2_u6_U24 (.B( u2_K7_32 ) , .A( u2_R5_21 ) , .Z( u2_u6_X_32 ) );
  XOR2_X1 u2_u6_U25 (.B( u2_K7_31 ) , .A( u2_R5_20 ) , .Z( u2_u6_X_31 ) );
  XOR2_X1 u2_u6_U26 (.B( u2_K7_30 ) , .A( u2_R5_21 ) , .Z( u2_u6_X_30 ) );
  XOR2_X1 u2_u6_U28 (.B( u2_K7_29 ) , .A( u2_R5_20 ) , .Z( u2_u6_X_29 ) );
  XOR2_X1 u2_u6_U29 (.B( u2_K7_28 ) , .A( u2_R5_19 ) , .Z( u2_u6_X_28 ) );
  XOR2_X1 u2_u6_U30 (.B( u2_K7_27 ) , .A( u2_R5_18 ) , .Z( u2_u6_X_27 ) );
  XOR2_X1 u2_u6_U31 (.B( u2_K7_26 ) , .A( u2_R5_17 ) , .Z( u2_u6_X_26 ) );
  XOR2_X1 u2_u6_U32 (.B( u2_K7_25 ) , .A( u2_R5_16 ) , .Z( u2_u6_X_25 ) );
  XOR2_X1 u2_u6_U7 (.B( u2_K7_48 ) , .A( u2_R5_1 ) , .Z( u2_u6_X_48 ) );
  XOR2_X1 u2_u6_U8 (.B( u2_K7_47 ) , .A( u2_R5_32 ) , .Z( u2_u6_X_47 ) );
  XOR2_X1 u2_u6_U9 (.B( u2_K7_46 ) , .A( u2_R5_31 ) , .Z( u2_u6_X_46 ) );
  OAI22_X1 u2_u6_u4_U10 (.B2( u2_u6_u4_n135 ) , .ZN( u2_u6_u4_n137 ) , .B1( u2_u6_u4_n153 ) , .A1( u2_u6_u4_n155 ) , .A2( u2_u6_u4_n171 ) );
  AND3_X1 u2_u6_u4_U11 (.A2( u2_u6_u4_n134 ) , .ZN( u2_u6_u4_n135 ) , .A3( u2_u6_u4_n145 ) , .A1( u2_u6_u4_n157 ) );
  NAND2_X1 u2_u6_u4_U12 (.ZN( u2_u6_u4_n132 ) , .A2( u2_u6_u4_n170 ) , .A1( u2_u6_u4_n173 ) );
  AOI21_X1 u2_u6_u4_U13 (.B2( u2_u6_u4_n160 ) , .B1( u2_u6_u4_n161 ) , .ZN( u2_u6_u4_n162 ) , .A( u2_u6_u4_n170 ) );
  AOI21_X1 u2_u6_u4_U14 (.ZN( u2_u6_u4_n107 ) , .B2( u2_u6_u4_n143 ) , .A( u2_u6_u4_n174 ) , .B1( u2_u6_u4_n184 ) );
  AOI21_X1 u2_u6_u4_U15 (.B2( u2_u6_u4_n158 ) , .B1( u2_u6_u4_n159 ) , .ZN( u2_u6_u4_n163 ) , .A( u2_u6_u4_n174 ) );
  AOI21_X1 u2_u6_u4_U16 (.A( u2_u6_u4_n153 ) , .B2( u2_u6_u4_n154 ) , .B1( u2_u6_u4_n155 ) , .ZN( u2_u6_u4_n165 ) );
  AOI21_X1 u2_u6_u4_U17 (.A( u2_u6_u4_n156 ) , .B2( u2_u6_u4_n157 ) , .ZN( u2_u6_u4_n164 ) , .B1( u2_u6_u4_n184 ) );
  INV_X1 u2_u6_u4_U18 (.A( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n170 ) );
  AND2_X1 u2_u6_u4_U19 (.A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n155 ) , .A1( u2_u6_u4_n160 ) );
  INV_X1 u2_u6_u4_U20 (.A( u2_u6_u4_n156 ) , .ZN( u2_u6_u4_n175 ) );
  NAND2_X1 u2_u6_u4_U21 (.A2( u2_u6_u4_n118 ) , .ZN( u2_u6_u4_n131 ) , .A1( u2_u6_u4_n147 ) );
  NAND2_X1 u2_u6_u4_U22 (.A1( u2_u6_u4_n119 ) , .A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n130 ) );
  NAND2_X1 u2_u6_u4_U23 (.ZN( u2_u6_u4_n117 ) , .A2( u2_u6_u4_n118 ) , .A1( u2_u6_u4_n148 ) );
  NAND2_X1 u2_u6_u4_U24 (.ZN( u2_u6_u4_n129 ) , .A1( u2_u6_u4_n134 ) , .A2( u2_u6_u4_n148 ) );
  AND3_X1 u2_u6_u4_U25 (.A1( u2_u6_u4_n119 ) , .A2( u2_u6_u4_n143 ) , .A3( u2_u6_u4_n154 ) , .ZN( u2_u6_u4_n161 ) );
  AND2_X1 u2_u6_u4_U26 (.A1( u2_u6_u4_n145 ) , .A2( u2_u6_u4_n147 ) , .ZN( u2_u6_u4_n159 ) );
  OR3_X1 u2_u6_u4_U27 (.A3( u2_u6_u4_n114 ) , .A2( u2_u6_u4_n115 ) , .A1( u2_u6_u4_n116 ) , .ZN( u2_u6_u4_n136 ) );
  AOI21_X1 u2_u6_u4_U28 (.A( u2_u6_u4_n113 ) , .ZN( u2_u6_u4_n116 ) , .B2( u2_u6_u4_n173 ) , .B1( u2_u6_u4_n174 ) );
  AOI21_X1 u2_u6_u4_U29 (.ZN( u2_u6_u4_n115 ) , .B2( u2_u6_u4_n145 ) , .B1( u2_u6_u4_n146 ) , .A( u2_u6_u4_n156 ) );
  NOR2_X1 u2_u6_u4_U3 (.ZN( u2_u6_u4_n121 ) , .A1( u2_u6_u4_n181 ) , .A2( u2_u6_u4_n182 ) );
  OAI22_X1 u2_u6_u4_U30 (.ZN( u2_u6_u4_n114 ) , .A2( u2_u6_u4_n121 ) , .B1( u2_u6_u4_n160 ) , .B2( u2_u6_u4_n170 ) , .A1( u2_u6_u4_n171 ) );
  INV_X1 u2_u6_u4_U31 (.A( u2_u6_u4_n158 ) , .ZN( u2_u6_u4_n182 ) );
  INV_X1 u2_u6_u4_U32 (.ZN( u2_u6_u4_n181 ) , .A( u2_u6_u4_n96 ) );
  INV_X1 u2_u6_u4_U33 (.A( u2_u6_u4_n144 ) , .ZN( u2_u6_u4_n179 ) );
  INV_X1 u2_u6_u4_U34 (.A( u2_u6_u4_n157 ) , .ZN( u2_u6_u4_n178 ) );
  NAND2_X1 u2_u6_u4_U35 (.A2( u2_u6_u4_n154 ) , .A1( u2_u6_u4_n96 ) , .ZN( u2_u6_u4_n97 ) );
  INV_X1 u2_u6_u4_U36 (.ZN( u2_u6_u4_n186 ) , .A( u2_u6_u4_n95 ) );
  OAI221_X1 u2_u6_u4_U37 (.C1( u2_u6_u4_n134 ) , .B1( u2_u6_u4_n158 ) , .B2( u2_u6_u4_n171 ) , .C2( u2_u6_u4_n173 ) , .A( u2_u6_u4_n94 ) , .ZN( u2_u6_u4_n95 ) );
  AOI222_X1 u2_u6_u4_U38 (.B2( u2_u6_u4_n132 ) , .A1( u2_u6_u4_n138 ) , .C2( u2_u6_u4_n175 ) , .A2( u2_u6_u4_n179 ) , .C1( u2_u6_u4_n181 ) , .B1( u2_u6_u4_n185 ) , .ZN( u2_u6_u4_n94 ) );
  INV_X1 u2_u6_u4_U39 (.A( u2_u6_u4_n113 ) , .ZN( u2_u6_u4_n185 ) );
  INV_X1 u2_u6_u4_U4 (.A( u2_u6_u4_n117 ) , .ZN( u2_u6_u4_n184 ) );
  INV_X1 u2_u6_u4_U40 (.A( u2_u6_u4_n143 ) , .ZN( u2_u6_u4_n183 ) );
  NOR2_X1 u2_u6_u4_U41 (.ZN( u2_u6_u4_n138 ) , .A1( u2_u6_u4_n168 ) , .A2( u2_u6_u4_n169 ) );
  NOR2_X1 u2_u6_u4_U42 (.A1( u2_u6_u4_n150 ) , .A2( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n153 ) );
  NOR2_X1 u2_u6_u4_U43 (.A2( u2_u6_u4_n128 ) , .A1( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n156 ) );
  AOI22_X1 u2_u6_u4_U44 (.B2( u2_u6_u4_n122 ) , .A1( u2_u6_u4_n123 ) , .ZN( u2_u6_u4_n124 ) , .B1( u2_u6_u4_n128 ) , .A2( u2_u6_u4_n172 ) );
  INV_X1 u2_u6_u4_U45 (.A( u2_u6_u4_n153 ) , .ZN( u2_u6_u4_n172 ) );
  NAND2_X1 u2_u6_u4_U46 (.A2( u2_u6_u4_n120 ) , .ZN( u2_u6_u4_n123 ) , .A1( u2_u6_u4_n161 ) );
  AOI22_X1 u2_u6_u4_U47 (.B2( u2_u6_u4_n132 ) , .A2( u2_u6_u4_n133 ) , .ZN( u2_u6_u4_n140 ) , .A1( u2_u6_u4_n150 ) , .B1( u2_u6_u4_n179 ) );
  NAND2_X1 u2_u6_u4_U48 (.ZN( u2_u6_u4_n133 ) , .A2( u2_u6_u4_n146 ) , .A1( u2_u6_u4_n154 ) );
  NAND2_X1 u2_u6_u4_U49 (.A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n154 ) , .A2( u2_u6_u4_n98 ) );
  NOR4_X1 u2_u6_u4_U5 (.A4( u2_u6_u4_n106 ) , .A3( u2_u6_u4_n107 ) , .A2( u2_u6_u4_n108 ) , .A1( u2_u6_u4_n109 ) , .ZN( u2_u6_u4_n110 ) );
  NAND2_X1 u2_u6_u4_U50 (.A1( u2_u6_u4_n101 ) , .ZN( u2_u6_u4_n158 ) , .A2( u2_u6_u4_n99 ) );
  AOI21_X1 u2_u6_u4_U51 (.ZN( u2_u6_u4_n127 ) , .A( u2_u6_u4_n136 ) , .B2( u2_u6_u4_n150 ) , .B1( u2_u6_u4_n180 ) );
  INV_X1 u2_u6_u4_U52 (.A( u2_u6_u4_n160 ) , .ZN( u2_u6_u4_n180 ) );
  NAND2_X1 u2_u6_u4_U53 (.A2( u2_u6_u4_n104 ) , .A1( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n146 ) );
  NAND2_X1 u2_u6_u4_U54 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n160 ) );
  NAND2_X1 u2_u6_u4_U55 (.ZN( u2_u6_u4_n134 ) , .A1( u2_u6_u4_n98 ) , .A2( u2_u6_u4_n99 ) );
  NAND2_X1 u2_u6_u4_U56 (.A1( u2_u6_u4_n103 ) , .A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n143 ) );
  NAND2_X1 u2_u6_u4_U57 (.A2( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n145 ) , .A1( u2_u6_u4_n98 ) );
  NAND2_X1 u2_u6_u4_U58 (.A1( u2_u6_u4_n100 ) , .A2( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n120 ) );
  NAND2_X1 u2_u6_u4_U59 (.A1( u2_u6_u4_n102 ) , .A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n148 ) );
  AOI21_X1 u2_u6_u4_U6 (.ZN( u2_u6_u4_n106 ) , .B2( u2_u6_u4_n146 ) , .B1( u2_u6_u4_n158 ) , .A( u2_u6_u4_n170 ) );
  NAND2_X1 u2_u6_u4_U60 (.A2( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n157 ) );
  INV_X1 u2_u6_u4_U61 (.A( u2_u6_u4_n150 ) , .ZN( u2_u6_u4_n173 ) );
  INV_X1 u2_u6_u4_U62 (.A( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n171 ) );
  NAND2_X1 u2_u6_u4_U63 (.A1( u2_u6_u4_n100 ) , .ZN( u2_u6_u4_n118 ) , .A2( u2_u6_u4_n99 ) );
  NAND2_X1 u2_u6_u4_U64 (.A2( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n144 ) );
  NAND2_X1 u2_u6_u4_U65 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n105 ) , .ZN( u2_u6_u4_n96 ) );
  INV_X1 u2_u6_u4_U66 (.A( u2_u6_u4_n128 ) , .ZN( u2_u6_u4_n174 ) );
  NAND2_X1 u2_u6_u4_U67 (.A2( u2_u6_u4_n102 ) , .ZN( u2_u6_u4_n119 ) , .A1( u2_u6_u4_n98 ) );
  NAND2_X1 u2_u6_u4_U68 (.A2( u2_u6_u4_n101 ) , .A1( u2_u6_u4_n103 ) , .ZN( u2_u6_u4_n147 ) );
  NAND2_X1 u2_u6_u4_U69 (.A2( u2_u6_u4_n104 ) , .ZN( u2_u6_u4_n113 ) , .A1( u2_u6_u4_n99 ) );
  AOI21_X1 u2_u6_u4_U7 (.ZN( u2_u6_u4_n108 ) , .B2( u2_u6_u4_n134 ) , .B1( u2_u6_u4_n155 ) , .A( u2_u6_u4_n156 ) );
  NOR2_X1 u2_u6_u4_U70 (.A2( u2_u6_X_28 ) , .ZN( u2_u6_u4_n150 ) , .A1( u2_u6_u4_n168 ) );
  NOR2_X1 u2_u6_u4_U71 (.A2( u2_u6_X_29 ) , .ZN( u2_u6_u4_n152 ) , .A1( u2_u6_u4_n169 ) );
  NOR2_X1 u2_u6_u4_U72 (.A2( u2_u6_X_30 ) , .ZN( u2_u6_u4_n105 ) , .A1( u2_u6_u4_n176 ) );
  NOR2_X1 u2_u6_u4_U73 (.A2( u2_u6_X_26 ) , .ZN( u2_u6_u4_n100 ) , .A1( u2_u6_u4_n177 ) );
  NOR2_X1 u2_u6_u4_U74 (.A2( u2_u6_X_28 ) , .A1( u2_u6_X_29 ) , .ZN( u2_u6_u4_n128 ) );
  NOR2_X1 u2_u6_u4_U75 (.A2( u2_u6_X_27 ) , .A1( u2_u6_X_30 ) , .ZN( u2_u6_u4_n102 ) );
  NOR2_X1 u2_u6_u4_U76 (.A2( u2_u6_X_25 ) , .A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n98 ) );
  AND2_X1 u2_u6_u4_U77 (.A2( u2_u6_X_25 ) , .A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n104 ) );
  AND2_X1 u2_u6_u4_U78 (.A1( u2_u6_X_30 ) , .A2( u2_u6_u4_n176 ) , .ZN( u2_u6_u4_n99 ) );
  AND2_X1 u2_u6_u4_U79 (.A1( u2_u6_X_26 ) , .ZN( u2_u6_u4_n101 ) , .A2( u2_u6_u4_n177 ) );
  AOI21_X1 u2_u6_u4_U8 (.ZN( u2_u6_u4_n109 ) , .A( u2_u6_u4_n153 ) , .B1( u2_u6_u4_n159 ) , .B2( u2_u6_u4_n184 ) );
  AND2_X1 u2_u6_u4_U80 (.A1( u2_u6_X_27 ) , .A2( u2_u6_X_30 ) , .ZN( u2_u6_u4_n103 ) );
  INV_X1 u2_u6_u4_U81 (.A( u2_u6_X_28 ) , .ZN( u2_u6_u4_n169 ) );
  INV_X1 u2_u6_u4_U82 (.A( u2_u6_X_29 ) , .ZN( u2_u6_u4_n168 ) );
  INV_X1 u2_u6_u4_U83 (.A( u2_u6_X_25 ) , .ZN( u2_u6_u4_n177 ) );
  INV_X1 u2_u6_u4_U84 (.A( u2_u6_X_27 ) , .ZN( u2_u6_u4_n176 ) );
  NAND4_X1 u2_u6_u4_U85 (.ZN( u2_out6_25 ) , .A4( u2_u6_u4_n139 ) , .A3( u2_u6_u4_n140 ) , .A2( u2_u6_u4_n141 ) , .A1( u2_u6_u4_n142 ) );
  OAI21_X1 u2_u6_u4_U86 (.B2( u2_u6_u4_n131 ) , .ZN( u2_u6_u4_n141 ) , .A( u2_u6_u4_n175 ) , .B1( u2_u6_u4_n183 ) );
  OAI21_X1 u2_u6_u4_U87 (.A( u2_u6_u4_n128 ) , .B2( u2_u6_u4_n129 ) , .B1( u2_u6_u4_n130 ) , .ZN( u2_u6_u4_n142 ) );
  NAND4_X1 u2_u6_u4_U88 (.ZN( u2_out6_14 ) , .A4( u2_u6_u4_n124 ) , .A3( u2_u6_u4_n125 ) , .A2( u2_u6_u4_n126 ) , .A1( u2_u6_u4_n127 ) );
  AOI22_X1 u2_u6_u4_U89 (.B2( u2_u6_u4_n117 ) , .ZN( u2_u6_u4_n126 ) , .A1( u2_u6_u4_n129 ) , .B1( u2_u6_u4_n152 ) , .A2( u2_u6_u4_n175 ) );
  AOI211_X1 u2_u6_u4_U9 (.B( u2_u6_u4_n136 ) , .A( u2_u6_u4_n137 ) , .C2( u2_u6_u4_n138 ) , .ZN( u2_u6_u4_n139 ) , .C1( u2_u6_u4_n182 ) );
  AOI22_X1 u2_u6_u4_U90 (.ZN( u2_u6_u4_n125 ) , .B2( u2_u6_u4_n131 ) , .A2( u2_u6_u4_n132 ) , .B1( u2_u6_u4_n138 ) , .A1( u2_u6_u4_n178 ) );
  NAND4_X1 u2_u6_u4_U91 (.ZN( u2_out6_8 ) , .A4( u2_u6_u4_n110 ) , .A3( u2_u6_u4_n111 ) , .A2( u2_u6_u4_n112 ) , .A1( u2_u6_u4_n186 ) );
  NAND2_X1 u2_u6_u4_U92 (.ZN( u2_u6_u4_n112 ) , .A2( u2_u6_u4_n130 ) , .A1( u2_u6_u4_n150 ) );
  AOI22_X1 u2_u6_u4_U93 (.ZN( u2_u6_u4_n111 ) , .B2( u2_u6_u4_n132 ) , .A1( u2_u6_u4_n152 ) , .B1( u2_u6_u4_n178 ) , .A2( u2_u6_u4_n97 ) );
  AOI22_X1 u2_u6_u4_U94 (.B2( u2_u6_u4_n149 ) , .B1( u2_u6_u4_n150 ) , .A2( u2_u6_u4_n151 ) , .A1( u2_u6_u4_n152 ) , .ZN( u2_u6_u4_n167 ) );
  NOR4_X1 u2_u6_u4_U95 (.A4( u2_u6_u4_n162 ) , .A3( u2_u6_u4_n163 ) , .A2( u2_u6_u4_n164 ) , .A1( u2_u6_u4_n165 ) , .ZN( u2_u6_u4_n166 ) );
  NAND3_X1 u2_u6_u4_U96 (.ZN( u2_out6_3 ) , .A3( u2_u6_u4_n166 ) , .A1( u2_u6_u4_n167 ) , .A2( u2_u6_u4_n186 ) );
  NAND3_X1 u2_u6_u4_U97 (.A3( u2_u6_u4_n146 ) , .A2( u2_u6_u4_n147 ) , .A1( u2_u6_u4_n148 ) , .ZN( u2_u6_u4_n149 ) );
  NAND3_X1 u2_u6_u4_U98 (.A3( u2_u6_u4_n143 ) , .A2( u2_u6_u4_n144 ) , .A1( u2_u6_u4_n145 ) , .ZN( u2_u6_u4_n151 ) );
  NAND3_X1 u2_u6_u4_U99 (.A3( u2_u6_u4_n121 ) , .ZN( u2_u6_u4_n122 ) , .A2( u2_u6_u4_n144 ) , .A1( u2_u6_u4_n154 ) );
  INV_X1 u2_u6_u5_U10 (.A( u2_u6_u5_n121 ) , .ZN( u2_u6_u5_n177 ) );
  NOR3_X1 u2_u6_u5_U100 (.A3( u2_u6_u5_n141 ) , .A1( u2_u6_u5_n142 ) , .ZN( u2_u6_u5_n143 ) , .A2( u2_u6_u5_n191 ) );
  NAND4_X1 u2_u6_u5_U101 (.ZN( u2_out6_4 ) , .A4( u2_u6_u5_n112 ) , .A2( u2_u6_u5_n113 ) , .A1( u2_u6_u5_n114 ) , .A3( u2_u6_u5_n195 ) );
  AOI211_X1 u2_u6_u5_U102 (.A( u2_u6_u5_n110 ) , .C1( u2_u6_u5_n111 ) , .ZN( u2_u6_u5_n112 ) , .B( u2_u6_u5_n118 ) , .C2( u2_u6_u5_n177 ) );
  AOI222_X1 u2_u6_u5_U103 (.ZN( u2_u6_u5_n113 ) , .A1( u2_u6_u5_n131 ) , .C1( u2_u6_u5_n148 ) , .B2( u2_u6_u5_n174 ) , .C2( u2_u6_u5_n178 ) , .A2( u2_u6_u5_n179 ) , .B1( u2_u6_u5_n99 ) );
  NAND3_X1 u2_u6_u5_U104 (.A2( u2_u6_u5_n154 ) , .A3( u2_u6_u5_n158 ) , .A1( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n99 ) );
  NOR2_X1 u2_u6_u5_U11 (.ZN( u2_u6_u5_n160 ) , .A2( u2_u6_u5_n173 ) , .A1( u2_u6_u5_n177 ) );
  INV_X1 u2_u6_u5_U12 (.A( u2_u6_u5_n150 ) , .ZN( u2_u6_u5_n174 ) );
  AOI21_X1 u2_u6_u5_U13 (.A( u2_u6_u5_n160 ) , .B2( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n162 ) , .B1( u2_u6_u5_n192 ) );
  INV_X1 u2_u6_u5_U14 (.A( u2_u6_u5_n159 ) , .ZN( u2_u6_u5_n192 ) );
  AOI21_X1 u2_u6_u5_U15 (.A( u2_u6_u5_n156 ) , .B2( u2_u6_u5_n157 ) , .B1( u2_u6_u5_n158 ) , .ZN( u2_u6_u5_n163 ) );
  AOI21_X1 u2_u6_u5_U16 (.B2( u2_u6_u5_n139 ) , .B1( u2_u6_u5_n140 ) , .ZN( u2_u6_u5_n141 ) , .A( u2_u6_u5_n150 ) );
  OAI21_X1 u2_u6_u5_U17 (.A( u2_u6_u5_n133 ) , .B2( u2_u6_u5_n134 ) , .B1( u2_u6_u5_n135 ) , .ZN( u2_u6_u5_n142 ) );
  OAI21_X1 u2_u6_u5_U18 (.ZN( u2_u6_u5_n133 ) , .B2( u2_u6_u5_n147 ) , .A( u2_u6_u5_n173 ) , .B1( u2_u6_u5_n188 ) );
  NAND2_X1 u2_u6_u5_U19 (.A2( u2_u6_u5_n119 ) , .A1( u2_u6_u5_n123 ) , .ZN( u2_u6_u5_n137 ) );
  INV_X1 u2_u6_u5_U20 (.A( u2_u6_u5_n155 ) , .ZN( u2_u6_u5_n194 ) );
  NAND2_X1 u2_u6_u5_U21 (.A1( u2_u6_u5_n121 ) , .ZN( u2_u6_u5_n132 ) , .A2( u2_u6_u5_n172 ) );
  NAND2_X1 u2_u6_u5_U22 (.A2( u2_u6_u5_n122 ) , .ZN( u2_u6_u5_n136 ) , .A1( u2_u6_u5_n154 ) );
  NAND2_X1 u2_u6_u5_U23 (.A2( u2_u6_u5_n119 ) , .A1( u2_u6_u5_n120 ) , .ZN( u2_u6_u5_n159 ) );
  INV_X1 u2_u6_u5_U24 (.A( u2_u6_u5_n156 ) , .ZN( u2_u6_u5_n175 ) );
  INV_X1 u2_u6_u5_U25 (.A( u2_u6_u5_n158 ) , .ZN( u2_u6_u5_n188 ) );
  INV_X1 u2_u6_u5_U26 (.A( u2_u6_u5_n152 ) , .ZN( u2_u6_u5_n179 ) );
  INV_X1 u2_u6_u5_U27 (.A( u2_u6_u5_n140 ) , .ZN( u2_u6_u5_n182 ) );
  INV_X1 u2_u6_u5_U28 (.A( u2_u6_u5_n151 ) , .ZN( u2_u6_u5_n183 ) );
  INV_X1 u2_u6_u5_U29 (.A( u2_u6_u5_n123 ) , .ZN( u2_u6_u5_n185 ) );
  NOR2_X1 u2_u6_u5_U3 (.ZN( u2_u6_u5_n134 ) , .A1( u2_u6_u5_n183 ) , .A2( u2_u6_u5_n190 ) );
  INV_X1 u2_u6_u5_U30 (.A( u2_u6_u5_n161 ) , .ZN( u2_u6_u5_n184 ) );
  INV_X1 u2_u6_u5_U31 (.A( u2_u6_u5_n139 ) , .ZN( u2_u6_u5_n189 ) );
  INV_X1 u2_u6_u5_U32 (.A( u2_u6_u5_n157 ) , .ZN( u2_u6_u5_n190 ) );
  INV_X1 u2_u6_u5_U33 (.A( u2_u6_u5_n120 ) , .ZN( u2_u6_u5_n193 ) );
  NAND2_X1 u2_u6_u5_U34 (.ZN( u2_u6_u5_n111 ) , .A1( u2_u6_u5_n140 ) , .A2( u2_u6_u5_n155 ) );
  INV_X1 u2_u6_u5_U35 (.A( u2_u6_u5_n117 ) , .ZN( u2_u6_u5_n196 ) );
  OAI221_X1 u2_u6_u5_U36 (.A( u2_u6_u5_n116 ) , .ZN( u2_u6_u5_n117 ) , .B2( u2_u6_u5_n119 ) , .C1( u2_u6_u5_n153 ) , .C2( u2_u6_u5_n158 ) , .B1( u2_u6_u5_n172 ) );
  AOI222_X1 u2_u6_u5_U37 (.ZN( u2_u6_u5_n116 ) , .B2( u2_u6_u5_n145 ) , .C1( u2_u6_u5_n148 ) , .A2( u2_u6_u5_n174 ) , .C2( u2_u6_u5_n177 ) , .B1( u2_u6_u5_n187 ) , .A1( u2_u6_u5_n193 ) );
  INV_X1 u2_u6_u5_U38 (.A( u2_u6_u5_n115 ) , .ZN( u2_u6_u5_n187 ) );
  NOR2_X1 u2_u6_u5_U39 (.ZN( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n170 ) , .A2( u2_u6_u5_n180 ) );
  INV_X1 u2_u6_u5_U4 (.A( u2_u6_u5_n138 ) , .ZN( u2_u6_u5_n191 ) );
  AOI22_X1 u2_u6_u5_U40 (.B2( u2_u6_u5_n131 ) , .A2( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n169 ) , .B1( u2_u6_u5_n174 ) , .A1( u2_u6_u5_n185 ) );
  NOR2_X1 u2_u6_u5_U41 (.A1( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n150 ) , .A2( u2_u6_u5_n173 ) );
  AOI21_X1 u2_u6_u5_U42 (.A( u2_u6_u5_n118 ) , .B2( u2_u6_u5_n145 ) , .ZN( u2_u6_u5_n168 ) , .B1( u2_u6_u5_n186 ) );
  INV_X1 u2_u6_u5_U43 (.A( u2_u6_u5_n122 ) , .ZN( u2_u6_u5_n186 ) );
  NOR2_X1 u2_u6_u5_U44 (.A1( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n152 ) , .A2( u2_u6_u5_n176 ) );
  NOR2_X1 u2_u6_u5_U45 (.A1( u2_u6_u5_n115 ) , .ZN( u2_u6_u5_n118 ) , .A2( u2_u6_u5_n153 ) );
  NOR2_X1 u2_u6_u5_U46 (.A2( u2_u6_u5_n145 ) , .ZN( u2_u6_u5_n156 ) , .A1( u2_u6_u5_n174 ) );
  NOR2_X1 u2_u6_u5_U47 (.ZN( u2_u6_u5_n121 ) , .A2( u2_u6_u5_n145 ) , .A1( u2_u6_u5_n176 ) );
  AOI22_X1 u2_u6_u5_U48 (.ZN( u2_u6_u5_n114 ) , .A2( u2_u6_u5_n137 ) , .A1( u2_u6_u5_n145 ) , .B2( u2_u6_u5_n175 ) , .B1( u2_u6_u5_n193 ) );
  OAI211_X1 u2_u6_u5_U49 (.B( u2_u6_u5_n124 ) , .A( u2_u6_u5_n125 ) , .C2( u2_u6_u5_n126 ) , .C1( u2_u6_u5_n127 ) , .ZN( u2_u6_u5_n128 ) );
  OAI21_X1 u2_u6_u5_U5 (.B2( u2_u6_u5_n136 ) , .B1( u2_u6_u5_n137 ) , .ZN( u2_u6_u5_n138 ) , .A( u2_u6_u5_n177 ) );
  NOR3_X1 u2_u6_u5_U50 (.ZN( u2_u6_u5_n127 ) , .A1( u2_u6_u5_n136 ) , .A3( u2_u6_u5_n148 ) , .A2( u2_u6_u5_n182 ) );
  OAI21_X1 u2_u6_u5_U51 (.ZN( u2_u6_u5_n124 ) , .A( u2_u6_u5_n177 ) , .B2( u2_u6_u5_n183 ) , .B1( u2_u6_u5_n189 ) );
  OAI21_X1 u2_u6_u5_U52 (.ZN( u2_u6_u5_n125 ) , .A( u2_u6_u5_n174 ) , .B2( u2_u6_u5_n185 ) , .B1( u2_u6_u5_n190 ) );
  AOI21_X1 u2_u6_u5_U53 (.A( u2_u6_u5_n153 ) , .B2( u2_u6_u5_n154 ) , .B1( u2_u6_u5_n155 ) , .ZN( u2_u6_u5_n164 ) );
  AOI21_X1 u2_u6_u5_U54 (.ZN( u2_u6_u5_n110 ) , .B1( u2_u6_u5_n122 ) , .B2( u2_u6_u5_n139 ) , .A( u2_u6_u5_n153 ) );
  INV_X1 u2_u6_u5_U55 (.A( u2_u6_u5_n153 ) , .ZN( u2_u6_u5_n176 ) );
  INV_X1 u2_u6_u5_U56 (.A( u2_u6_u5_n126 ) , .ZN( u2_u6_u5_n173 ) );
  AND2_X1 u2_u6_u5_U57 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n147 ) );
  AND2_X1 u2_u6_u5_U58 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n148 ) );
  NAND2_X1 u2_u6_u5_U59 (.A1( u2_u6_u5_n105 ) , .A2( u2_u6_u5_n106 ) , .ZN( u2_u6_u5_n158 ) );
  INV_X1 u2_u6_u5_U6 (.A( u2_u6_u5_n135 ) , .ZN( u2_u6_u5_n178 ) );
  NAND2_X1 u2_u6_u5_U60 (.A2( u2_u6_u5_n108 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n139 ) );
  NAND2_X1 u2_u6_u5_U61 (.A1( u2_u6_u5_n106 ) , .A2( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n119 ) );
  NAND2_X1 u2_u6_u5_U62 (.A2( u2_u6_u5_n103 ) , .A1( u2_u6_u5_n105 ) , .ZN( u2_u6_u5_n140 ) );
  NAND2_X1 u2_u6_u5_U63 (.A2( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n105 ) , .ZN( u2_u6_u5_n155 ) );
  NAND2_X1 u2_u6_u5_U64 (.A2( u2_u6_u5_n106 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n122 ) );
  NAND2_X1 u2_u6_u5_U65 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n106 ) , .ZN( u2_u6_u5_n115 ) );
  NAND2_X1 u2_u6_u5_U66 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n103 ) , .ZN( u2_u6_u5_n161 ) );
  NAND2_X1 u2_u6_u5_U67 (.A1( u2_u6_u5_n105 ) , .A2( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n154 ) );
  INV_X1 u2_u6_u5_U68 (.A( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n172 ) );
  NAND2_X1 u2_u6_u5_U69 (.A1( u2_u6_u5_n103 ) , .A2( u2_u6_u5_n108 ) , .ZN( u2_u6_u5_n123 ) );
  OAI22_X1 u2_u6_u5_U7 (.B2( u2_u6_u5_n149 ) , .B1( u2_u6_u5_n150 ) , .A2( u2_u6_u5_n151 ) , .A1( u2_u6_u5_n152 ) , .ZN( u2_u6_u5_n165 ) );
  NAND2_X1 u2_u6_u5_U70 (.A2( u2_u6_u5_n103 ) , .A1( u2_u6_u5_n107 ) , .ZN( u2_u6_u5_n151 ) );
  NAND2_X1 u2_u6_u5_U71 (.A2( u2_u6_u5_n107 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n120 ) );
  NAND2_X1 u2_u6_u5_U72 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n109 ) , .ZN( u2_u6_u5_n157 ) );
  AND2_X1 u2_u6_u5_U73 (.A2( u2_u6_u5_n100 ) , .A1( u2_u6_u5_n104 ) , .ZN( u2_u6_u5_n131 ) );
  INV_X1 u2_u6_u5_U74 (.A( u2_u6_u5_n102 ) , .ZN( u2_u6_u5_n195 ) );
  OAI221_X1 u2_u6_u5_U75 (.A( u2_u6_u5_n101 ) , .ZN( u2_u6_u5_n102 ) , .C2( u2_u6_u5_n115 ) , .C1( u2_u6_u5_n126 ) , .B1( u2_u6_u5_n134 ) , .B2( u2_u6_u5_n160 ) );
  OAI21_X1 u2_u6_u5_U76 (.ZN( u2_u6_u5_n101 ) , .B1( u2_u6_u5_n137 ) , .A( u2_u6_u5_n146 ) , .B2( u2_u6_u5_n147 ) );
  NOR2_X1 u2_u6_u5_U77 (.A2( u2_u6_X_34 ) , .A1( u2_u6_X_35 ) , .ZN( u2_u6_u5_n145 ) );
  NOR2_X1 u2_u6_u5_U78 (.A2( u2_u6_X_34 ) , .ZN( u2_u6_u5_n146 ) , .A1( u2_u6_u5_n171 ) );
  NOR2_X1 u2_u6_u5_U79 (.A2( u2_u6_X_31 ) , .A1( u2_u6_X_32 ) , .ZN( u2_u6_u5_n103 ) );
  NOR3_X1 u2_u6_u5_U8 (.A2( u2_u6_u5_n147 ) , .A1( u2_u6_u5_n148 ) , .ZN( u2_u6_u5_n149 ) , .A3( u2_u6_u5_n194 ) );
  NOR2_X1 u2_u6_u5_U80 (.A2( u2_u6_X_36 ) , .ZN( u2_u6_u5_n105 ) , .A1( u2_u6_u5_n180 ) );
  NOR2_X1 u2_u6_u5_U81 (.A2( u2_u6_X_33 ) , .ZN( u2_u6_u5_n108 ) , .A1( u2_u6_u5_n170 ) );
  NOR2_X1 u2_u6_u5_U82 (.A2( u2_u6_X_33 ) , .A1( u2_u6_X_36 ) , .ZN( u2_u6_u5_n107 ) );
  NOR2_X1 u2_u6_u5_U83 (.A2( u2_u6_X_31 ) , .ZN( u2_u6_u5_n104 ) , .A1( u2_u6_u5_n181 ) );
  NAND2_X1 u2_u6_u5_U84 (.A2( u2_u6_X_34 ) , .A1( u2_u6_X_35 ) , .ZN( u2_u6_u5_n153 ) );
  NAND2_X1 u2_u6_u5_U85 (.A1( u2_u6_X_34 ) , .ZN( u2_u6_u5_n126 ) , .A2( u2_u6_u5_n171 ) );
  AND2_X1 u2_u6_u5_U86 (.A1( u2_u6_X_31 ) , .A2( u2_u6_X_32 ) , .ZN( u2_u6_u5_n106 ) );
  AND2_X1 u2_u6_u5_U87 (.A1( u2_u6_X_31 ) , .ZN( u2_u6_u5_n109 ) , .A2( u2_u6_u5_n181 ) );
  INV_X1 u2_u6_u5_U88 (.A( u2_u6_X_33 ) , .ZN( u2_u6_u5_n180 ) );
  INV_X1 u2_u6_u5_U89 (.A( u2_u6_X_35 ) , .ZN( u2_u6_u5_n171 ) );
  NOR2_X1 u2_u6_u5_U9 (.ZN( u2_u6_u5_n135 ) , .A1( u2_u6_u5_n173 ) , .A2( u2_u6_u5_n176 ) );
  INV_X1 u2_u6_u5_U90 (.A( u2_u6_X_36 ) , .ZN( u2_u6_u5_n170 ) );
  INV_X1 u2_u6_u5_U91 (.A( u2_u6_X_32 ) , .ZN( u2_u6_u5_n181 ) );
  NAND4_X1 u2_u6_u5_U92 (.ZN( u2_out6_29 ) , .A4( u2_u6_u5_n129 ) , .A3( u2_u6_u5_n130 ) , .A2( u2_u6_u5_n168 ) , .A1( u2_u6_u5_n196 ) );
  AOI221_X1 u2_u6_u5_U93 (.A( u2_u6_u5_n128 ) , .ZN( u2_u6_u5_n129 ) , .C2( u2_u6_u5_n132 ) , .B2( u2_u6_u5_n159 ) , .B1( u2_u6_u5_n176 ) , .C1( u2_u6_u5_n184 ) );
  AOI222_X1 u2_u6_u5_U94 (.ZN( u2_u6_u5_n130 ) , .A2( u2_u6_u5_n146 ) , .B1( u2_u6_u5_n147 ) , .C2( u2_u6_u5_n175 ) , .B2( u2_u6_u5_n179 ) , .A1( u2_u6_u5_n188 ) , .C1( u2_u6_u5_n194 ) );
  NAND4_X1 u2_u6_u5_U95 (.ZN( u2_out6_19 ) , .A4( u2_u6_u5_n166 ) , .A3( u2_u6_u5_n167 ) , .A2( u2_u6_u5_n168 ) , .A1( u2_u6_u5_n169 ) );
  AOI22_X1 u2_u6_u5_U96 (.B2( u2_u6_u5_n145 ) , .A2( u2_u6_u5_n146 ) , .ZN( u2_u6_u5_n167 ) , .B1( u2_u6_u5_n182 ) , .A1( u2_u6_u5_n189 ) );
  NOR4_X1 u2_u6_u5_U97 (.A4( u2_u6_u5_n162 ) , .A3( u2_u6_u5_n163 ) , .A2( u2_u6_u5_n164 ) , .A1( u2_u6_u5_n165 ) , .ZN( u2_u6_u5_n166 ) );
  NAND4_X1 u2_u6_u5_U98 (.ZN( u2_out6_11 ) , .A4( u2_u6_u5_n143 ) , .A3( u2_u6_u5_n144 ) , .A2( u2_u6_u5_n169 ) , .A1( u2_u6_u5_n196 ) );
  AOI22_X1 u2_u6_u5_U99 (.A2( u2_u6_u5_n132 ) , .ZN( u2_u6_u5_n144 ) , .B2( u2_u6_u5_n145 ) , .B1( u2_u6_u5_n184 ) , .A1( u2_u6_u5_n194 ) );
  AOI21_X1 u2_u6_u6_U10 (.ZN( u2_u6_u6_n106 ) , .A( u2_u6_u6_n142 ) , .B2( u2_u6_u6_n159 ) , .B1( u2_u6_u6_n164 ) );
  INV_X1 u2_u6_u6_U11 (.A( u2_u6_u6_n155 ) , .ZN( u2_u6_u6_n161 ) );
  INV_X1 u2_u6_u6_U12 (.A( u2_u6_u6_n128 ) , .ZN( u2_u6_u6_n164 ) );
  NAND2_X1 u2_u6_u6_U13 (.ZN( u2_u6_u6_n110 ) , .A1( u2_u6_u6_n122 ) , .A2( u2_u6_u6_n129 ) );
  NAND2_X1 u2_u6_u6_U14 (.ZN( u2_u6_u6_n124 ) , .A2( u2_u6_u6_n146 ) , .A1( u2_u6_u6_n148 ) );
  INV_X1 u2_u6_u6_U15 (.A( u2_u6_u6_n132 ) , .ZN( u2_u6_u6_n171 ) );
  AND2_X1 u2_u6_u6_U16 (.A1( u2_u6_u6_n100 ) , .ZN( u2_u6_u6_n130 ) , .A2( u2_u6_u6_n147 ) );
  INV_X1 u2_u6_u6_U17 (.A( u2_u6_u6_n127 ) , .ZN( u2_u6_u6_n173 ) );
  INV_X1 u2_u6_u6_U18 (.A( u2_u6_u6_n121 ) , .ZN( u2_u6_u6_n167 ) );
  INV_X1 u2_u6_u6_U19 (.A( u2_u6_u6_n100 ) , .ZN( u2_u6_u6_n169 ) );
  INV_X1 u2_u6_u6_U20 (.A( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n170 ) );
  INV_X1 u2_u6_u6_U21 (.A( u2_u6_u6_n113 ) , .ZN( u2_u6_u6_n168 ) );
  AND2_X1 u2_u6_u6_U22 (.A1( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n119 ) , .ZN( u2_u6_u6_n133 ) );
  AND2_X1 u2_u6_u6_U23 (.A2( u2_u6_u6_n121 ) , .A1( u2_u6_u6_n122 ) , .ZN( u2_u6_u6_n131 ) );
  AND3_X1 u2_u6_u6_U24 (.ZN( u2_u6_u6_n120 ) , .A2( u2_u6_u6_n127 ) , .A1( u2_u6_u6_n132 ) , .A3( u2_u6_u6_n145 ) );
  INV_X1 u2_u6_u6_U25 (.A( u2_u6_u6_n146 ) , .ZN( u2_u6_u6_n163 ) );
  AOI222_X1 u2_u6_u6_U26 (.ZN( u2_u6_u6_n114 ) , .A1( u2_u6_u6_n118 ) , .A2( u2_u6_u6_n126 ) , .B2( u2_u6_u6_n151 ) , .C2( u2_u6_u6_n159 ) , .C1( u2_u6_u6_n168 ) , .B1( u2_u6_u6_n169 ) );
  NOR2_X1 u2_u6_u6_U27 (.A1( u2_u6_u6_n162 ) , .A2( u2_u6_u6_n165 ) , .ZN( u2_u6_u6_n98 ) );
  AOI211_X1 u2_u6_u6_U28 (.B( u2_u6_u6_n149 ) , .A( u2_u6_u6_n150 ) , .C2( u2_u6_u6_n151 ) , .C1( u2_u6_u6_n152 ) , .ZN( u2_u6_u6_n153 ) );
  AOI21_X1 u2_u6_u6_U29 (.B2( u2_u6_u6_n147 ) , .B1( u2_u6_u6_n148 ) , .ZN( u2_u6_u6_n149 ) , .A( u2_u6_u6_n158 ) );
  INV_X1 u2_u6_u6_U3 (.A( u2_u6_u6_n110 ) , .ZN( u2_u6_u6_n166 ) );
  AOI21_X1 u2_u6_u6_U30 (.A( u2_u6_u6_n144 ) , .B2( u2_u6_u6_n145 ) , .B1( u2_u6_u6_n146 ) , .ZN( u2_u6_u6_n150 ) );
  NAND2_X1 u2_u6_u6_U31 (.A2( u2_u6_u6_n143 ) , .ZN( u2_u6_u6_n152 ) , .A1( u2_u6_u6_n166 ) );
  NAND2_X1 u2_u6_u6_U32 (.A1( u2_u6_u6_n144 ) , .ZN( u2_u6_u6_n151 ) , .A2( u2_u6_u6_n158 ) );
  NAND2_X1 u2_u6_u6_U33 (.ZN( u2_u6_u6_n132 ) , .A1( u2_u6_u6_n91 ) , .A2( u2_u6_u6_n97 ) );
  AOI22_X1 u2_u6_u6_U34 (.B2( u2_u6_u6_n110 ) , .B1( u2_u6_u6_n111 ) , .A1( u2_u6_u6_n112 ) , .ZN( u2_u6_u6_n115 ) , .A2( u2_u6_u6_n161 ) );
  NAND4_X1 u2_u6_u6_U35 (.A3( u2_u6_u6_n109 ) , .ZN( u2_u6_u6_n112 ) , .A4( u2_u6_u6_n132 ) , .A2( u2_u6_u6_n147 ) , .A1( u2_u6_u6_n166 ) );
  NOR2_X1 u2_u6_u6_U36 (.ZN( u2_u6_u6_n109 ) , .A1( u2_u6_u6_n170 ) , .A2( u2_u6_u6_n173 ) );
  NOR2_X1 u2_u6_u6_U37 (.A2( u2_u6_u6_n126 ) , .ZN( u2_u6_u6_n155 ) , .A1( u2_u6_u6_n160 ) );
  NAND2_X1 u2_u6_u6_U38 (.ZN( u2_u6_u6_n146 ) , .A2( u2_u6_u6_n94 ) , .A1( u2_u6_u6_n99 ) );
  AOI211_X1 u2_u6_u6_U39 (.B( u2_u6_u6_n134 ) , .A( u2_u6_u6_n135 ) , .C1( u2_u6_u6_n136 ) , .ZN( u2_u6_u6_n137 ) , .C2( u2_u6_u6_n151 ) );
  AOI22_X1 u2_u6_u6_U4 (.B2( u2_u6_u6_n101 ) , .A1( u2_u6_u6_n102 ) , .ZN( u2_u6_u6_n103 ) , .B1( u2_u6_u6_n160 ) , .A2( u2_u6_u6_n161 ) );
  NAND4_X1 u2_u6_u6_U40 (.A4( u2_u6_u6_n127 ) , .A3( u2_u6_u6_n128 ) , .A2( u2_u6_u6_n129 ) , .A1( u2_u6_u6_n130 ) , .ZN( u2_u6_u6_n136 ) );
  AOI21_X1 u2_u6_u6_U41 (.B2( u2_u6_u6_n132 ) , .B1( u2_u6_u6_n133 ) , .ZN( u2_u6_u6_n134 ) , .A( u2_u6_u6_n158 ) );
  AOI21_X1 u2_u6_u6_U42 (.B1( u2_u6_u6_n131 ) , .ZN( u2_u6_u6_n135 ) , .A( u2_u6_u6_n144 ) , .B2( u2_u6_u6_n146 ) );
  INV_X1 u2_u6_u6_U43 (.A( u2_u6_u6_n111 ) , .ZN( u2_u6_u6_n158 ) );
  NAND2_X1 u2_u6_u6_U44 (.ZN( u2_u6_u6_n127 ) , .A1( u2_u6_u6_n91 ) , .A2( u2_u6_u6_n92 ) );
  NAND2_X1 u2_u6_u6_U45 (.ZN( u2_u6_u6_n129 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n96 ) );
  INV_X1 u2_u6_u6_U46 (.A( u2_u6_u6_n144 ) , .ZN( u2_u6_u6_n159 ) );
  NAND2_X1 u2_u6_u6_U47 (.ZN( u2_u6_u6_n145 ) , .A2( u2_u6_u6_n97 ) , .A1( u2_u6_u6_n98 ) );
  NAND2_X1 u2_u6_u6_U48 (.ZN( u2_u6_u6_n148 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n94 ) );
  NAND2_X1 u2_u6_u6_U49 (.ZN( u2_u6_u6_n108 ) , .A2( u2_u6_u6_n139 ) , .A1( u2_u6_u6_n144 ) );
  NOR2_X1 u2_u6_u6_U5 (.A1( u2_u6_u6_n118 ) , .ZN( u2_u6_u6_n143 ) , .A2( u2_u6_u6_n168 ) );
  NAND2_X1 u2_u6_u6_U50 (.ZN( u2_u6_u6_n121 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n97 ) );
  NAND2_X1 u2_u6_u6_U51 (.ZN( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n95 ) );
  AND2_X1 u2_u6_u6_U52 (.ZN( u2_u6_u6_n118 ) , .A2( u2_u6_u6_n91 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U53 (.ZN( u2_u6_u6_n147 ) , .A2( u2_u6_u6_n98 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U54 (.ZN( u2_u6_u6_n128 ) , .A1( u2_u6_u6_n94 ) , .A2( u2_u6_u6_n96 ) );
  NAND2_X1 u2_u6_u6_U55 (.ZN( u2_u6_u6_n119 ) , .A2( u2_u6_u6_n95 ) , .A1( u2_u6_u6_n99 ) );
  NAND2_X1 u2_u6_u6_U56 (.ZN( u2_u6_u6_n123 ) , .A2( u2_u6_u6_n91 ) , .A1( u2_u6_u6_n96 ) );
  NAND2_X1 u2_u6_u6_U57 (.ZN( u2_u6_u6_n100 ) , .A2( u2_u6_u6_n92 ) , .A1( u2_u6_u6_n98 ) );
  NAND2_X1 u2_u6_u6_U58 (.ZN( u2_u6_u6_n122 ) , .A1( u2_u6_u6_n94 ) , .A2( u2_u6_u6_n97 ) );
  INV_X1 u2_u6_u6_U59 (.A( u2_u6_u6_n139 ) , .ZN( u2_u6_u6_n160 ) );
  AOI21_X1 u2_u6_u6_U6 (.B1( u2_u6_u6_n107 ) , .B2( u2_u6_u6_n132 ) , .A( u2_u6_u6_n158 ) , .ZN( u2_u6_u6_n88 ) );
  NAND2_X1 u2_u6_u6_U60 (.ZN( u2_u6_u6_n113 ) , .A1( u2_u6_u6_n96 ) , .A2( u2_u6_u6_n98 ) );
  NOR2_X1 u2_u6_u6_U61 (.A2( u2_u6_X_40 ) , .A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n126 ) );
  NOR2_X1 u2_u6_u6_U62 (.A2( u2_u6_X_39 ) , .A1( u2_u6_X_42 ) , .ZN( u2_u6_u6_n92 ) );
  NOR2_X1 u2_u6_u6_U63 (.A2( u2_u6_X_39 ) , .A1( u2_u6_u6_n156 ) , .ZN( u2_u6_u6_n97 ) );
  NOR2_X1 u2_u6_u6_U64 (.A2( u2_u6_X_38 ) , .A1( u2_u6_u6_n165 ) , .ZN( u2_u6_u6_n95 ) );
  NOR2_X1 u2_u6_u6_U65 (.A2( u2_u6_X_41 ) , .ZN( u2_u6_u6_n111 ) , .A1( u2_u6_u6_n157 ) );
  NOR2_X1 u2_u6_u6_U66 (.A2( u2_u6_X_37 ) , .A1( u2_u6_u6_n162 ) , .ZN( u2_u6_u6_n94 ) );
  NOR2_X1 u2_u6_u6_U67 (.A2( u2_u6_X_37 ) , .A1( u2_u6_X_38 ) , .ZN( u2_u6_u6_n91 ) );
  NAND2_X1 u2_u6_u6_U68 (.A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n144 ) , .A2( u2_u6_u6_n157 ) );
  NAND2_X1 u2_u6_u6_U69 (.A2( u2_u6_X_40 ) , .A1( u2_u6_X_41 ) , .ZN( u2_u6_u6_n139 ) );
  OAI21_X1 u2_u6_u6_U7 (.A( u2_u6_u6_n159 ) , .B1( u2_u6_u6_n169 ) , .B2( u2_u6_u6_n173 ) , .ZN( u2_u6_u6_n90 ) );
  AND2_X1 u2_u6_u6_U70 (.A1( u2_u6_X_39 ) , .A2( u2_u6_u6_n156 ) , .ZN( u2_u6_u6_n96 ) );
  AND2_X1 u2_u6_u6_U71 (.A1( u2_u6_X_39 ) , .A2( u2_u6_X_42 ) , .ZN( u2_u6_u6_n99 ) );
  INV_X1 u2_u6_u6_U72 (.A( u2_u6_X_40 ) , .ZN( u2_u6_u6_n157 ) );
  INV_X1 u2_u6_u6_U73 (.A( u2_u6_X_37 ) , .ZN( u2_u6_u6_n165 ) );
  INV_X1 u2_u6_u6_U74 (.A( u2_u6_X_38 ) , .ZN( u2_u6_u6_n162 ) );
  INV_X1 u2_u6_u6_U75 (.A( u2_u6_X_42 ) , .ZN( u2_u6_u6_n156 ) );
  NAND4_X1 u2_u6_u6_U76 (.ZN( u2_out6_32 ) , .A4( u2_u6_u6_n103 ) , .A3( u2_u6_u6_n104 ) , .A2( u2_u6_u6_n105 ) , .A1( u2_u6_u6_n106 ) );
  AOI22_X1 u2_u6_u6_U77 (.ZN( u2_u6_u6_n104 ) , .A1( u2_u6_u6_n111 ) , .B1( u2_u6_u6_n124 ) , .B2( u2_u6_u6_n151 ) , .A2( u2_u6_u6_n93 ) );
  AOI22_X1 u2_u6_u6_U78 (.ZN( u2_u6_u6_n105 ) , .A2( u2_u6_u6_n108 ) , .A1( u2_u6_u6_n118 ) , .B2( u2_u6_u6_n126 ) , .B1( u2_u6_u6_n171 ) );
  NAND4_X1 u2_u6_u6_U79 (.ZN( u2_out6_12 ) , .A4( u2_u6_u6_n114 ) , .A3( u2_u6_u6_n115 ) , .A2( u2_u6_u6_n116 ) , .A1( u2_u6_u6_n117 ) );
  INV_X1 u2_u6_u6_U8 (.ZN( u2_u6_u6_n172 ) , .A( u2_u6_u6_n88 ) );
  OAI22_X1 u2_u6_u6_U80 (.B2( u2_u6_u6_n111 ) , .ZN( u2_u6_u6_n116 ) , .B1( u2_u6_u6_n126 ) , .A2( u2_u6_u6_n164 ) , .A1( u2_u6_u6_n167 ) );
  OAI21_X1 u2_u6_u6_U81 (.A( u2_u6_u6_n108 ) , .ZN( u2_u6_u6_n117 ) , .B2( u2_u6_u6_n141 ) , .B1( u2_u6_u6_n163 ) );
  OAI211_X1 u2_u6_u6_U82 (.ZN( u2_out6_22 ) , .B( u2_u6_u6_n137 ) , .A( u2_u6_u6_n138 ) , .C2( u2_u6_u6_n139 ) , .C1( u2_u6_u6_n140 ) );
  AOI22_X1 u2_u6_u6_U83 (.B1( u2_u6_u6_n124 ) , .A2( u2_u6_u6_n125 ) , .A1( u2_u6_u6_n126 ) , .ZN( u2_u6_u6_n138 ) , .B2( u2_u6_u6_n161 ) );
  AND4_X1 u2_u6_u6_U84 (.A3( u2_u6_u6_n119 ) , .A1( u2_u6_u6_n120 ) , .A4( u2_u6_u6_n129 ) , .ZN( u2_u6_u6_n140 ) , .A2( u2_u6_u6_n143 ) );
  OAI211_X1 u2_u6_u6_U85 (.ZN( u2_out6_7 ) , .B( u2_u6_u6_n153 ) , .C2( u2_u6_u6_n154 ) , .C1( u2_u6_u6_n155 ) , .A( u2_u6_u6_n174 ) );
  NOR3_X1 u2_u6_u6_U86 (.A1( u2_u6_u6_n141 ) , .ZN( u2_u6_u6_n154 ) , .A3( u2_u6_u6_n164 ) , .A2( u2_u6_u6_n171 ) );
  INV_X1 u2_u6_u6_U87 (.A( u2_u6_u6_n142 ) , .ZN( u2_u6_u6_n174 ) );
  NAND3_X1 u2_u6_u6_U88 (.A2( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n125 ) , .A1( u2_u6_u6_n130 ) , .A3( u2_u6_u6_n131 ) );
  NAND3_X1 u2_u6_u6_U89 (.A3( u2_u6_u6_n133 ) , .ZN( u2_u6_u6_n141 ) , .A1( u2_u6_u6_n145 ) , .A2( u2_u6_u6_n148 ) );
  AOI22_X1 u2_u6_u6_U9 (.A2( u2_u6_u6_n151 ) , .B2( u2_u6_u6_n161 ) , .A1( u2_u6_u6_n167 ) , .B1( u2_u6_u6_n170 ) , .ZN( u2_u6_u6_n89 ) );
  NAND3_X1 u2_u6_u6_U90 (.ZN( u2_u6_u6_n101 ) , .A3( u2_u6_u6_n107 ) , .A2( u2_u6_u6_n121 ) , .A1( u2_u6_u6_n127 ) );
  NAND3_X1 u2_u6_u6_U91 (.ZN( u2_u6_u6_n102 ) , .A3( u2_u6_u6_n130 ) , .A2( u2_u6_u6_n145 ) , .A1( u2_u6_u6_n166 ) );
  NAND3_X1 u2_u6_u6_U92 (.A3( u2_u6_u6_n113 ) , .A1( u2_u6_u6_n119 ) , .A2( u2_u6_u6_n123 ) , .ZN( u2_u6_u6_n93 ) );
  NAND3_X1 u2_u6_u6_U93 (.ZN( u2_u6_u6_n142 ) , .A2( u2_u6_u6_n172 ) , .A3( u2_u6_u6_n89 ) , .A1( u2_u6_u6_n90 ) );
  AND3_X1 u2_u6_u7_U10 (.A3( u2_u6_u7_n110 ) , .A2( u2_u6_u7_n127 ) , .A1( u2_u6_u7_n132 ) , .ZN( u2_u6_u7_n92 ) );
  OAI21_X1 u2_u6_u7_U11 (.A( u2_u6_u7_n161 ) , .B1( u2_u6_u7_n168 ) , .B2( u2_u6_u7_n173 ) , .ZN( u2_u6_u7_n91 ) );
  AOI211_X1 u2_u6_u7_U12 (.A( u2_u6_u7_n117 ) , .ZN( u2_u6_u7_n118 ) , .C2( u2_u6_u7_n126 ) , .C1( u2_u6_u7_n177 ) , .B( u2_u6_u7_n180 ) );
  OAI22_X1 u2_u6_u7_U13 (.B1( u2_u6_u7_n115 ) , .ZN( u2_u6_u7_n117 ) , .A2( u2_u6_u7_n133 ) , .A1( u2_u6_u7_n137 ) , .B2( u2_u6_u7_n162 ) );
  INV_X1 u2_u6_u7_U14 (.A( u2_u6_u7_n116 ) , .ZN( u2_u6_u7_n180 ) );
  NOR3_X1 u2_u6_u7_U15 (.ZN( u2_u6_u7_n115 ) , .A3( u2_u6_u7_n145 ) , .A2( u2_u6_u7_n168 ) , .A1( u2_u6_u7_n169 ) );
  OAI211_X1 u2_u6_u7_U16 (.B( u2_u6_u7_n122 ) , .A( u2_u6_u7_n123 ) , .C2( u2_u6_u7_n124 ) , .ZN( u2_u6_u7_n154 ) , .C1( u2_u6_u7_n162 ) );
  AOI222_X1 u2_u6_u7_U17 (.ZN( u2_u6_u7_n122 ) , .C2( u2_u6_u7_n126 ) , .C1( u2_u6_u7_n145 ) , .B1( u2_u6_u7_n161 ) , .A2( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n170 ) , .A1( u2_u6_u7_n176 ) );
  INV_X1 u2_u6_u7_U18 (.A( u2_u6_u7_n133 ) , .ZN( u2_u6_u7_n176 ) );
  NOR3_X1 u2_u6_u7_U19 (.A2( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n135 ) , .ZN( u2_u6_u7_n136 ) , .A3( u2_u6_u7_n171 ) );
  NOR2_X1 u2_u6_u7_U20 (.A1( u2_u6_u7_n130 ) , .A2( u2_u6_u7_n134 ) , .ZN( u2_u6_u7_n153 ) );
  INV_X1 u2_u6_u7_U21 (.A( u2_u6_u7_n101 ) , .ZN( u2_u6_u7_n165 ) );
  NOR2_X1 u2_u6_u7_U22 (.ZN( u2_u6_u7_n111 ) , .A2( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n169 ) );
  AOI21_X1 u2_u6_u7_U23 (.ZN( u2_u6_u7_n104 ) , .B2( u2_u6_u7_n112 ) , .B1( u2_u6_u7_n127 ) , .A( u2_u6_u7_n164 ) );
  AOI21_X1 u2_u6_u7_U24 (.ZN( u2_u6_u7_n106 ) , .B1( u2_u6_u7_n133 ) , .B2( u2_u6_u7_n146 ) , .A( u2_u6_u7_n162 ) );
  AOI21_X1 u2_u6_u7_U25 (.A( u2_u6_u7_n101 ) , .ZN( u2_u6_u7_n107 ) , .B2( u2_u6_u7_n128 ) , .B1( u2_u6_u7_n175 ) );
  INV_X1 u2_u6_u7_U26 (.A( u2_u6_u7_n138 ) , .ZN( u2_u6_u7_n171 ) );
  INV_X1 u2_u6_u7_U27 (.A( u2_u6_u7_n131 ) , .ZN( u2_u6_u7_n177 ) );
  INV_X1 u2_u6_u7_U28 (.A( u2_u6_u7_n110 ) , .ZN( u2_u6_u7_n174 ) );
  NAND2_X1 u2_u6_u7_U29 (.A1( u2_u6_u7_n129 ) , .A2( u2_u6_u7_n132 ) , .ZN( u2_u6_u7_n149 ) );
  OAI21_X1 u2_u6_u7_U3 (.ZN( u2_u6_u7_n159 ) , .A( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n171 ) , .B1( u2_u6_u7_n174 ) );
  NAND2_X1 u2_u6_u7_U30 (.A1( u2_u6_u7_n113 ) , .A2( u2_u6_u7_n124 ) , .ZN( u2_u6_u7_n130 ) );
  INV_X1 u2_u6_u7_U31 (.A( u2_u6_u7_n112 ) , .ZN( u2_u6_u7_n173 ) );
  INV_X1 u2_u6_u7_U32 (.A( u2_u6_u7_n128 ) , .ZN( u2_u6_u7_n168 ) );
  INV_X1 u2_u6_u7_U33 (.A( u2_u6_u7_n148 ) , .ZN( u2_u6_u7_n169 ) );
  INV_X1 u2_u6_u7_U34 (.A( u2_u6_u7_n127 ) , .ZN( u2_u6_u7_n179 ) );
  NOR2_X1 u2_u6_u7_U35 (.ZN( u2_u6_u7_n101 ) , .A2( u2_u6_u7_n150 ) , .A1( u2_u6_u7_n156 ) );
  AOI211_X1 u2_u6_u7_U36 (.B( u2_u6_u7_n154 ) , .A( u2_u6_u7_n155 ) , .C1( u2_u6_u7_n156 ) , .ZN( u2_u6_u7_n157 ) , .C2( u2_u6_u7_n172 ) );
  INV_X1 u2_u6_u7_U37 (.A( u2_u6_u7_n153 ) , .ZN( u2_u6_u7_n172 ) );
  AOI211_X1 u2_u6_u7_U38 (.B( u2_u6_u7_n139 ) , .A( u2_u6_u7_n140 ) , .C2( u2_u6_u7_n141 ) , .ZN( u2_u6_u7_n142 ) , .C1( u2_u6_u7_n156 ) );
  NAND4_X1 u2_u6_u7_U39 (.A3( u2_u6_u7_n127 ) , .A2( u2_u6_u7_n128 ) , .A1( u2_u6_u7_n129 ) , .ZN( u2_u6_u7_n141 ) , .A4( u2_u6_u7_n147 ) );
  INV_X1 u2_u6_u7_U4 (.A( u2_u6_u7_n111 ) , .ZN( u2_u6_u7_n170 ) );
  AOI21_X1 u2_u6_u7_U40 (.A( u2_u6_u7_n137 ) , .B1( u2_u6_u7_n138 ) , .ZN( u2_u6_u7_n139 ) , .B2( u2_u6_u7_n146 ) );
  OAI22_X1 u2_u6_u7_U41 (.B1( u2_u6_u7_n136 ) , .ZN( u2_u6_u7_n140 ) , .A1( u2_u6_u7_n153 ) , .B2( u2_u6_u7_n162 ) , .A2( u2_u6_u7_n164 ) );
  AOI21_X1 u2_u6_u7_U42 (.ZN( u2_u6_u7_n123 ) , .B1( u2_u6_u7_n165 ) , .B2( u2_u6_u7_n177 ) , .A( u2_u6_u7_n97 ) );
  AOI21_X1 u2_u6_u7_U43 (.B2( u2_u6_u7_n113 ) , .B1( u2_u6_u7_n124 ) , .A( u2_u6_u7_n125 ) , .ZN( u2_u6_u7_n97 ) );
  INV_X1 u2_u6_u7_U44 (.A( u2_u6_u7_n125 ) , .ZN( u2_u6_u7_n161 ) );
  INV_X1 u2_u6_u7_U45 (.A( u2_u6_u7_n152 ) , .ZN( u2_u6_u7_n162 ) );
  AOI22_X1 u2_u6_u7_U46 (.A2( u2_u6_u7_n114 ) , .ZN( u2_u6_u7_n119 ) , .B1( u2_u6_u7_n130 ) , .A1( u2_u6_u7_n156 ) , .B2( u2_u6_u7_n165 ) );
  NAND2_X1 u2_u6_u7_U47 (.A2( u2_u6_u7_n112 ) , .ZN( u2_u6_u7_n114 ) , .A1( u2_u6_u7_n175 ) );
  AND2_X1 u2_u6_u7_U48 (.ZN( u2_u6_u7_n145 ) , .A2( u2_u6_u7_n98 ) , .A1( u2_u6_u7_n99 ) );
  NOR2_X1 u2_u6_u7_U49 (.ZN( u2_u6_u7_n137 ) , .A1( u2_u6_u7_n150 ) , .A2( u2_u6_u7_n161 ) );
  INV_X1 u2_u6_u7_U5 (.A( u2_u6_u7_n149 ) , .ZN( u2_u6_u7_n175 ) );
  AOI21_X1 u2_u6_u7_U50 (.ZN( u2_u6_u7_n105 ) , .B2( u2_u6_u7_n110 ) , .A( u2_u6_u7_n125 ) , .B1( u2_u6_u7_n147 ) );
  NAND2_X1 u2_u6_u7_U51 (.ZN( u2_u6_u7_n146 ) , .A1( u2_u6_u7_n95 ) , .A2( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U52 (.A2( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n147 ) , .A1( u2_u6_u7_n93 ) );
  NAND2_X1 u2_u6_u7_U53 (.A1( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n127 ) , .A2( u2_u6_u7_n99 ) );
  OR2_X1 u2_u6_u7_U54 (.ZN( u2_u6_u7_n126 ) , .A2( u2_u6_u7_n152 ) , .A1( u2_u6_u7_n156 ) );
  NAND2_X1 u2_u6_u7_U55 (.A2( u2_u6_u7_n102 ) , .A1( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n133 ) );
  NAND2_X1 u2_u6_u7_U56 (.ZN( u2_u6_u7_n112 ) , .A2( u2_u6_u7_n96 ) , .A1( u2_u6_u7_n99 ) );
  NAND2_X1 u2_u6_u7_U57 (.A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n128 ) , .A1( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U58 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n113 ) , .A2( u2_u6_u7_n93 ) );
  NAND2_X1 u2_u6_u7_U59 (.A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n124 ) , .A1( u2_u6_u7_n96 ) );
  INV_X1 u2_u6_u7_U6 (.A( u2_u6_u7_n154 ) , .ZN( u2_u6_u7_n178 ) );
  NAND2_X1 u2_u6_u7_U60 (.ZN( u2_u6_u7_n110 ) , .A1( u2_u6_u7_n95 ) , .A2( u2_u6_u7_n96 ) );
  INV_X1 u2_u6_u7_U61 (.A( u2_u6_u7_n150 ) , .ZN( u2_u6_u7_n164 ) );
  AND2_X1 u2_u6_u7_U62 (.ZN( u2_u6_u7_n134 ) , .A1( u2_u6_u7_n93 ) , .A2( u2_u6_u7_n98 ) );
  NAND2_X1 u2_u6_u7_U63 (.A1( u2_u6_u7_n100 ) , .A2( u2_u6_u7_n102 ) , .ZN( u2_u6_u7_n129 ) );
  NAND2_X1 u2_u6_u7_U64 (.A2( u2_u6_u7_n103 ) , .ZN( u2_u6_u7_n131 ) , .A1( u2_u6_u7_n95 ) );
  NAND2_X1 u2_u6_u7_U65 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n138 ) , .A2( u2_u6_u7_n99 ) );
  NAND2_X1 u2_u6_u7_U66 (.ZN( u2_u6_u7_n132 ) , .A1( u2_u6_u7_n93 ) , .A2( u2_u6_u7_n96 ) );
  NAND2_X1 u2_u6_u7_U67 (.A1( u2_u6_u7_n100 ) , .ZN( u2_u6_u7_n148 ) , .A2( u2_u6_u7_n95 ) );
  NOR2_X1 u2_u6_u7_U68 (.A2( u2_u6_X_47 ) , .ZN( u2_u6_u7_n150 ) , .A1( u2_u6_u7_n163 ) );
  NOR2_X1 u2_u6_u7_U69 (.A2( u2_u6_X_43 ) , .A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n103 ) );
  AOI211_X1 u2_u6_u7_U7 (.ZN( u2_u6_u7_n116 ) , .A( u2_u6_u7_n155 ) , .C1( u2_u6_u7_n161 ) , .C2( u2_u6_u7_n171 ) , .B( u2_u6_u7_n94 ) );
  NOR2_X1 u2_u6_u7_U70 (.A2( u2_u6_X_48 ) , .A1( u2_u6_u7_n166 ) , .ZN( u2_u6_u7_n95 ) );
  NOR2_X1 u2_u6_u7_U71 (.A2( u2_u6_X_45 ) , .A1( u2_u6_X_48 ) , .ZN( u2_u6_u7_n99 ) );
  NOR2_X1 u2_u6_u7_U72 (.A2( u2_u6_X_44 ) , .A1( u2_u6_u7_n167 ) , .ZN( u2_u6_u7_n98 ) );
  NOR2_X1 u2_u6_u7_U73 (.A2( u2_u6_X_46 ) , .A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n152 ) );
  AND2_X1 u2_u6_u7_U74 (.A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n156 ) , .A2( u2_u6_u7_n163 ) );
  NAND2_X1 u2_u6_u7_U75 (.A2( u2_u6_X_46 ) , .A1( u2_u6_X_47 ) , .ZN( u2_u6_u7_n125 ) );
  AND2_X1 u2_u6_u7_U76 (.A2( u2_u6_X_45 ) , .A1( u2_u6_X_48 ) , .ZN( u2_u6_u7_n102 ) );
  AND2_X1 u2_u6_u7_U77 (.A2( u2_u6_X_43 ) , .A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n96 ) );
  AND2_X1 u2_u6_u7_U78 (.A1( u2_u6_X_44 ) , .ZN( u2_u6_u7_n100 ) , .A2( u2_u6_u7_n167 ) );
  AND2_X1 u2_u6_u7_U79 (.A1( u2_u6_X_48 ) , .A2( u2_u6_u7_n166 ) , .ZN( u2_u6_u7_n93 ) );
  OAI222_X1 u2_u6_u7_U8 (.C2( u2_u6_u7_n101 ) , .B2( u2_u6_u7_n111 ) , .A1( u2_u6_u7_n113 ) , .C1( u2_u6_u7_n146 ) , .A2( u2_u6_u7_n162 ) , .B1( u2_u6_u7_n164 ) , .ZN( u2_u6_u7_n94 ) );
  INV_X1 u2_u6_u7_U80 (.A( u2_u6_X_46 ) , .ZN( u2_u6_u7_n163 ) );
  INV_X1 u2_u6_u7_U81 (.A( u2_u6_X_43 ) , .ZN( u2_u6_u7_n167 ) );
  INV_X1 u2_u6_u7_U82 (.A( u2_u6_X_45 ) , .ZN( u2_u6_u7_n166 ) );
  NAND4_X1 u2_u6_u7_U83 (.ZN( u2_out6_5 ) , .A4( u2_u6_u7_n108 ) , .A3( u2_u6_u7_n109 ) , .A1( u2_u6_u7_n116 ) , .A2( u2_u6_u7_n123 ) );
  AOI22_X1 u2_u6_u7_U84 (.ZN( u2_u6_u7_n109 ) , .A2( u2_u6_u7_n126 ) , .B2( u2_u6_u7_n145 ) , .B1( u2_u6_u7_n156 ) , .A1( u2_u6_u7_n171 ) );
  NOR4_X1 u2_u6_u7_U85 (.A4( u2_u6_u7_n104 ) , .A3( u2_u6_u7_n105 ) , .A2( u2_u6_u7_n106 ) , .A1( u2_u6_u7_n107 ) , .ZN( u2_u6_u7_n108 ) );
  NAND4_X1 u2_u6_u7_U86 (.ZN( u2_out6_27 ) , .A4( u2_u6_u7_n118 ) , .A3( u2_u6_u7_n119 ) , .A2( u2_u6_u7_n120 ) , .A1( u2_u6_u7_n121 ) );
  OAI21_X1 u2_u6_u7_U87 (.ZN( u2_u6_u7_n121 ) , .B2( u2_u6_u7_n145 ) , .A( u2_u6_u7_n150 ) , .B1( u2_u6_u7_n174 ) );
  OAI21_X1 u2_u6_u7_U88 (.ZN( u2_u6_u7_n120 ) , .A( u2_u6_u7_n161 ) , .B2( u2_u6_u7_n170 ) , .B1( u2_u6_u7_n179 ) );
  NAND4_X1 u2_u6_u7_U89 (.ZN( u2_out6_21 ) , .A4( u2_u6_u7_n157 ) , .A3( u2_u6_u7_n158 ) , .A2( u2_u6_u7_n159 ) , .A1( u2_u6_u7_n160 ) );
  OAI221_X1 u2_u6_u7_U9 (.C1( u2_u6_u7_n101 ) , .C2( u2_u6_u7_n147 ) , .ZN( u2_u6_u7_n155 ) , .B2( u2_u6_u7_n162 ) , .A( u2_u6_u7_n91 ) , .B1( u2_u6_u7_n92 ) );
  OAI21_X1 u2_u6_u7_U90 (.B1( u2_u6_u7_n145 ) , .ZN( u2_u6_u7_n160 ) , .A( u2_u6_u7_n161 ) , .B2( u2_u6_u7_n177 ) );
  AOI22_X1 u2_u6_u7_U91 (.B2( u2_u6_u7_n149 ) , .B1( u2_u6_u7_n150 ) , .A2( u2_u6_u7_n151 ) , .A1( u2_u6_u7_n152 ) , .ZN( u2_u6_u7_n158 ) );
  NAND4_X1 u2_u6_u7_U92 (.ZN( u2_out6_15 ) , .A4( u2_u6_u7_n142 ) , .A3( u2_u6_u7_n143 ) , .A2( u2_u6_u7_n144 ) , .A1( u2_u6_u7_n178 ) );
  OR2_X1 u2_u6_u7_U93 (.A2( u2_u6_u7_n125 ) , .A1( u2_u6_u7_n129 ) , .ZN( u2_u6_u7_n144 ) );
  AOI22_X1 u2_u6_u7_U94 (.A2( u2_u6_u7_n126 ) , .ZN( u2_u6_u7_n143 ) , .B2( u2_u6_u7_n165 ) , .B1( u2_u6_u7_n173 ) , .A1( u2_u6_u7_n174 ) );
  NAND3_X1 u2_u6_u7_U95 (.A3( u2_u6_u7_n146 ) , .A2( u2_u6_u7_n147 ) , .A1( u2_u6_u7_n148 ) , .ZN( u2_u6_u7_n151 ) );
  NAND3_X1 u2_u6_u7_U96 (.A3( u2_u6_u7_n131 ) , .A2( u2_u6_u7_n132 ) , .A1( u2_u6_u7_n133 ) , .ZN( u2_u6_u7_n135 ) );
  NAND2_X1 u2_uk_U1008 (.A1( u2_key_r_50 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n983 ) );
  OAI21_X1 u2_uk_U1074 (.ZN( u2_K16_39 ) , .B2( u2_uk_n1201 ) , .B1( u2_uk_n202 ) , .A( u2_uk_n960 ) );
  NAND2_X1 u2_uk_U1075 (.A1( u2_uk_K_r14_15 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n960 ) );
  INV_X1 u2_uk_U1120 (.ZN( u2_K7_32 ) , .A( u2_uk_n1088 ) );
  AOI22_X1 u2_uk_U1121 (.B2( u2_uk_K_r5_0 ) , .A2( u2_uk_K_r5_51 ) , .ZN( u2_uk_n1088 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U117 (.ZN( u2_K7_47 ) , .A2( u2_uk_n1456 ) , .B2( u2_uk_n1470 ) , .A1( u2_uk_n164 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U267 (.ZN( u2_K7_44 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1459 ) , .A2( u2_uk_n1480 ) );
  INV_X1 u2_uk_U348 (.ZN( u2_K7_46 ) , .A( u2_uk_n1094 ) );
  OAI22_X1 u2_uk_U354 (.ZN( u2_K16_40 ) , .B2( u2_uk_n1188 ) , .A2( u2_uk_n1226 ) , .B1( u2_uk_n238 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U359 (.ZN( u2_K7_40 ) , .A2( u2_uk_n1452 ) , .B2( u2_uk_n1464 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U380 (.ZN( u2_K7_28 ) , .B2( u2_uk_n1471 ) , .A2( u2_uk_n1480 ) , .A1( u2_uk_n223 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U441 (.ZN( u2_K16_37 ) , .A( u2_uk_n959 ) );
  AOI22_X1 u2_uk_U442 (.B2( u2_uk_K_r14_2 ) , .A2( u2_uk_K_r14_50 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n959 ) );
  OAI22_X1 u2_uk_U452 (.ZN( u2_K16_33 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1220 ) , .A2( u2_uk_n1225 ) , .A1( u2_uk_n129 ) );
  OAI22_X1 u2_uk_U493 (.ZN( u2_K7_29 ) , .B2( u2_uk_n1459 ) , .A2( u2_uk_n1490 ) , .A1( u2_uk_n238 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U52 (.ZN( u2_K16_34 ) , .A( u2_uk_n958 ) );
  AOI22_X1 u2_uk_U53 (.B2( u2_uk_K_r14_2 ) , .A2( u2_uk_K_r14_9 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n238 ) , .ZN( u2_uk_n958 ) );
  INV_X1 u2_uk_U557 (.ZN( u2_K7_36 ) , .A( u2_uk_n1091 ) );
  AOI22_X1 u2_uk_U558 (.B2( u2_uk_K_r5_1 ) , .A2( u2_uk_K_r5_21 ) , .ZN( u2_uk_n1091 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n202 ) );
  OAI22_X1 u2_uk_U563 (.ZN( u2_K16_36 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1203 ) , .A2( u2_uk_n1210 ) , .A1( u2_uk_n129 ) );
  INV_X1 u2_uk_U58 (.ZN( u2_K7_34 ) , .A( u2_uk_n1089 ) );
  OAI22_X1 u2_uk_U604 (.ZN( u2_K16_35 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1208 ) , .A2( u2_uk_n1215 ) , .A1( u2_uk_n129 ) );
  INV_X1 u2_uk_U701 (.ZN( u2_K7_25 ) , .A( u2_uk_n1084 ) );
  AOI22_X1 u2_uk_U702 (.B2( u2_uk_K_r5_31 ) , .A2( u2_uk_K_r5_7 ) , .A1( u2_uk_n10 ) , .ZN( u2_uk_n1084 ) , .B1( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U714 (.ZN( u2_K16_32 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1201 ) , .A2( u2_uk_n1209 ) , .A1( u2_uk_n202 ) );
  INV_X1 u2_uk_U737 (.ZN( u2_K7_42 ) , .A( u2_uk_n1093 ) );
  INV_X1 u2_uk_U789 (.ZN( u2_K7_27 ) , .A( u2_uk_n1085 ) );
  AOI22_X1 u2_uk_U790 (.B2( u2_uk_K_r5_23 ) , .A2( u2_uk_K_r5_43 ) , .ZN( u2_uk_n1085 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n141 ) );
  OAI21_X1 u2_uk_U80 (.ZN( u2_K16_41 ) , .B2( u2_uk_n1215 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n961 ) );
  OAI22_X1 u2_uk_U888 (.ZN( u2_K7_30 ) , .B2( u2_uk_n1460 ) , .A2( u2_uk_n1491 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U897 (.ZN( u2_K16_38 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1210 ) , .A2( u2_uk_n1217 ) , .A1( u2_uk_n161 ) );
  OAI22_X1 u2_uk_U899 (.ZN( u2_K7_39 ) , .B2( u2_uk_n1486 ) , .A2( u2_uk_n1493 ) , .A1( u2_uk_n161 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U9 (.A( u2_uk_n129 ) , .ZN( u2_uk_n31 ) );
  OAI22_X1 u2_uk_U90 (.ZN( u2_K7_41 ) , .A1( u2_uk_n118 ) , .A2( u2_uk_n1456 ) , .B2( u2_uk_n1486 ) , .B1( u2_uk_n208 ) );
endmodule

