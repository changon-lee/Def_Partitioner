module aes_aes_die_19 ( sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7 );
  input sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7;
  output sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7;
  wire us23_n438, us23_n439, us23_n440, us23_n441, us23_n442, us23_n443, us23_n444, us23_n445, us23_n446, 
       us23_n447, us23_n448, us23_n449, us23_n450, us23_n451, us23_n452, us23_n453, us23_n454, us23_n455, 
       us23_n456, us23_n457, us23_n458, us23_n459, us23_n460, us23_n461, us23_n462, us23_n463, us23_n464, 
       us23_n465, us23_n466, us23_n467, us23_n468, us23_n469, us23_n470, us23_n471, us23_n472, us23_n473, 
       us23_n474, us23_n475, us23_n476, us23_n477, us23_n478, us23_n479, us23_n480, us23_n481, us23_n482, 
       us23_n483, us23_n484, us23_n485, us23_n486, us23_n487, us23_n488, us23_n489, us23_n490, us23_n491, 
       us23_n492, us23_n493, us23_n494, us23_n495, us23_n496, us23_n497, us23_n498, us23_n499, us23_n500, 
       us23_n501, us23_n502, us23_n503, us23_n504, us23_n505, us23_n506, us23_n507, us23_n508, us23_n509, 
       us23_n510, us23_n511, us23_n512, us23_n513, us23_n514, us23_n515, us23_n516, us23_n517, us23_n518, 
       us23_n519, us23_n520, us23_n521, us23_n522, us23_n523, us23_n524, us23_n525, us23_n526, us23_n527, 
       us23_n528, us23_n529, us23_n530, us23_n531, us23_n532, us23_n533, us23_n534, us23_n535, us23_n536, 
       us23_n537, us23_n538, us23_n539, us23_n540, us23_n541, us23_n542, us23_n543, us23_n544, us23_n545, 
       us23_n546, us23_n547, us23_n548, us23_n549, us23_n550, us23_n551, us23_n552, us23_n553, us23_n554, 
       us23_n555, us23_n556, us23_n557, us23_n558, us23_n559, us23_n560, us23_n561, us23_n562, us23_n563, 
       us23_n564, us23_n565, us23_n566, us23_n567, us23_n568, us23_n569, us23_n570, us23_n571, us23_n572, 
       us23_n573, us23_n574, us23_n575, us23_n576, us23_n577, us23_n578, us23_n579, us23_n580, us23_n581, 
       us23_n582, us23_n583, us23_n584, us23_n585, us23_n586, us23_n587, us23_n588, us23_n589, us23_n590, 
       us23_n591, us23_n592, us23_n593, us23_n594, us23_n595, us23_n596, us23_n597, us23_n598, us23_n599, 
       us23_n600, us23_n601, us23_n602, us23_n603, us23_n604, us23_n605, us23_n606, us23_n607, us23_n608, 
       us23_n609, us23_n610, us23_n611, us23_n612, us23_n613, us23_n614, us23_n615, us23_n616, us23_n617, 
       us23_n618, us23_n619, us23_n620, us23_n621, us23_n622, us23_n623, us23_n624, us23_n625, us23_n626, 
       us23_n627, us23_n628, us23_n629, us23_n630, us23_n631, us23_n632, us23_n633, us23_n634, us23_n635, 
       us23_n636, us23_n637, us23_n638, us23_n639, us23_n640, us23_n641, us23_n642, us23_n643, us23_n644, 
       us23_n645, us23_n646, us23_n647, us23_n648, us23_n649, us23_n650, us23_n651, us23_n652, us23_n653, 
       us23_n654, us23_n655, us23_n656, us23_n657, us23_n658, us23_n659, us23_n660, us23_n661, us23_n662, 
       us23_n663, us23_n664, us23_n665, us23_n666, us23_n667, us23_n668, us23_n669, us23_n670, us23_n671, 
       us23_n672, us23_n673, us23_n674, us23_n675, us23_n676, us23_n677, us23_n678, us23_n679, us23_n680, 
       us23_n681, us23_n682, us23_n683, us23_n684, us23_n685, us23_n686, us23_n687, us23_n688, us23_n689, 
       us23_n690, us23_n691, us23_n692, us23_n693, us23_n694, us23_n695, us23_n696, us23_n697, us23_n698, 
       us23_n699, us23_n700, us23_n701, us23_n702, us23_n703, us23_n704, us23_n705, us23_n706, us23_n707, 
       us23_n708, us23_n709, us23_n710, us23_n711, us23_n712, us23_n713, us23_n714, us23_n715, us23_n716, 
       us23_n717, us23_n718, us23_n719, us23_n720, us23_n721, us23_n722, us23_n723, us23_n724, us23_n725, 
       us23_n726, us23_n727, us23_n728, us23_n729, us23_n730, us23_n731, us23_n732, us23_n733, us23_n734, 
       us23_n735, us23_n736, us23_n737, us23_n738, us23_n739, us23_n740, us23_n741, us23_n742, us23_n743, 
       us23_n744, us23_n745, us23_n746, us23_n747, us23_n748, us23_n749, us23_n750, us23_n751, us23_n752, 
       us23_n753, us23_n754, us23_n755, us23_n756, us23_n757, us23_n758, us23_n759, us23_n760, us23_n761, 
       us23_n762, us23_n763, us23_n764, us23_n765, us23_n766, us23_n767, us23_n768, us23_n769, us23_n770, 
       us23_n771, us23_n772, us23_n773, us23_n774, us23_n775, us23_n776, us23_n777, us23_n778, us23_n779, 
       us23_n780, us23_n781, us23_n782, us23_n783, us23_n784, us23_n785, us23_n786, us23_n787, us23_n788, 
       us23_n789, us23_n790, us23_n791, us23_n792, us23_n793, us23_n794, us23_n795, us23_n796, us23_n797, 
       us23_n798, us23_n799, us23_n800, us23_n801, us23_n802, us23_n803, us23_n804, us23_n805, us23_n806, 
       us23_n807, us23_n808, us23_n809, us23_n810, us23_n811, us23_n812, us23_n813, us23_n814, us23_n815, 
       us23_n816, us23_n817, us23_n818, us23_n819, us23_n820, us23_n821, us23_n822, us23_n823, us23_n824, 
       us23_n825, us23_n826, us23_n827, us23_n828, us23_n829, us23_n830, us23_n831, us23_n832, us23_n833, 
       us23_n834, us23_n835, us23_n836, us23_n837, us23_n838, us23_n839, us23_n840, us23_n841, us23_n842, 
       us23_n843, us23_n844, us23_n845, us23_n846, us23_n847, us23_n848, us23_n849, us23_n850, us23_n851, 
       us23_n852, us23_n853, us23_n854, us23_n855, us23_n856, us23_n857, us23_n858, us23_n859, us23_n860, 
       us23_n861, us23_n862, us23_n863, us23_n864, us23_n865, us23_n866, us23_n867, us23_n868, us23_n869, 
       us23_n870, us23_n871, us23_n872, us23_n873, us23_n874,  us23_n875;
  INV_X1 us23_U10 (.A( us23_n679 ) , .ZN( us23_n839 ) );
  NOR4_X1 us23_U100 (.A4( us23_n483 ) , .ZN( us23_n486 ) , .A1( us23_n565 ) , .A2( us23_n580 ) , .A3( us23_n601 ) );
  NOR4_X1 us23_U101 (.ZN( us23_n485 ) , .A1( us23_n506 ) , .A2( us23_n518 ) , .A4( us23_n545 ) , .A3( us23_n610 ) );
  NOR4_X1 us23_U102 (.ZN( us23_n484 ) , .A2( us23_n532 ) , .A1( us23_n557 ) , .A3( us23_n630 ) , .A4( us23_n717 ) );
  NAND4_X1 us23_U103 (.A4( us23_n690 ) , .A3( us23_n691 ) , .A1( us23_n692 ) , .ZN( us23_n775 ) , .A2( us23_n871 ) );
  AOI221_X1 us23_U104 (.A( us23_n680 ) , .ZN( us23_n691 ) , .B2( us23_n839 ) , .C1( us23_n841 ) , .C2( us23_n861 ) , .B1( us23_n864 ) );
  INV_X1 us23_U105 (.A( us23_n678 ) , .ZN( us23_n871 ) );
  NOR4_X1 us23_U106 (.A4( us23_n686 ) , .A3( us23_n687 ) , .A2( us23_n688 ) , .A1( us23_n689 ) , .ZN( us23_n690 ) );
  NAND4_X1 us23_U107 (.A4( us23_n559 ) , .A3( us23_n560 ) , .A2( us23_n561 ) , .A1( us23_n562 ) , .ZN( us23_n606 ) );
  NOR4_X1 us23_U108 (.ZN( us23_n560 ) , .A1( us23_n652 ) , .A3( us23_n660 ) , .A4( us23_n684 ) , .A2( us23_n767 ) );
  NOR4_X1 us23_U109 (.A4( us23_n551 ) , .A3( us23_n552 ) , .A2( us23_n553 ) , .A1( us23_n554 ) , .ZN( us23_n561 ) );
  NOR4_X1 us23_U11 (.A4( us23_n444 ) , .A3( us23_n445 ) , .A2( us23_n515 ) , .A1( us23_n540 ) , .ZN( us23_n705 ) );
  NOR4_X1 us23_U110 (.A4( us23_n555 ) , .A3( us23_n556 ) , .A2( us23_n557 ) , .A1( us23_n558 ) , .ZN( us23_n559 ) );
  NAND4_X1 us23_U111 (.A4( us23_n718 ) , .A3( us23_n719 ) , .A2( us23_n720 ) , .ZN( us23_n740 ) , .A1( us23_n856 ) );
  INV_X1 us23_U112 (.A( us23_n708 ) , .ZN( us23_n856 ) );
  AOI221_X1 us23_U113 (.A( us23_n709 ) , .ZN( us23_n720 ) , .C2( us23_n843 ) , .B2( us23_n844 ) , .C1( us23_n860 ) , .B1( us23_n861 ) );
  NOR4_X1 us23_U114 (.A4( us23_n714 ) , .A3( us23_n715 ) , .A2( us23_n716 ) , .A1( us23_n717 ) , .ZN( us23_n718 ) );
  NAND4_X1 us23_U115 (.A4( us23_n472 ) , .A3( us23_n473 ) , .A2( us23_n474 ) , .A1( us23_n475 ) , .ZN( us23_n677 ) );
  NOR4_X1 us23_U116 (.A4( us23_n469 ) , .ZN( us23_n475 ) , .A3( us23_n555 ) , .A1( us23_n734 ) , .A2( us23_n754 ) );
  NOR4_X1 us23_U117 (.ZN( us23_n474 ) , .A1( us23_n530 ) , .A3( us23_n567 ) , .A4( us23_n599 ) , .A2( us23_n641 ) );
  NOR4_X1 us23_U118 (.ZN( us23_n473 ) , .A1( us23_n505 ) , .A3( us23_n543 ) , .A2( us23_n582 ) , .A4( us23_n715 ) );
  NOR2_X1 us23_U119 (.ZN( us23_n732 ) , .A2( us23_n831 ) , .A1( us23_n844 ) );
  OR3_X1 us23_U12 (.ZN( us23_n445 ) , .A1( us23_n527 ) , .A3( us23_n576 ) , .A2( us23_n874 ) );
  NOR2_X1 us23_U120 (.ZN( us23_n788 ) , .A2( us23_n861 ) , .A1( us23_n867 ) );
  NAND4_X1 us23_U121 (.A4( us23_n572 ) , .A3( us23_n573 ) , .A1( us23_n574 ) , .ZN( us23_n722 ) , .A2( us23_n873 ) );
  NOR4_X1 us23_U122 (.A4( us23_n568 ) , .A3( us23_n569 ) , .A2( us23_n570 ) , .A1( us23_n571 ) , .ZN( us23_n572 ) );
  AOI221_X1 us23_U123 (.A( us23_n563 ) , .C2( us23_n564 ) , .ZN( us23_n573 ) , .B2( us23_n844 ) , .B1( us23_n851 ) , .C1( us23_n852 ) );
  INV_X1 us23_U124 (.A( us23_n606 ) , .ZN( us23_n873 ) );
  NAND4_X1 us23_U125 (.A4( us23_n492 ) , .A3( us23_n493 ) , .A1( us23_n494 ) , .ZN( us23_n801 ) , .A2( us23_n866 ) );
  AOI221_X1 us23_U126 (.A( us23_n488 ) , .ZN( us23_n493 ) , .B2( us23_n835 ) , .C2( us23_n840 ) , .C1( us23_n850 ) , .B1( us23_n859 ) );
  INV_X1 us23_U127 (.A( us23_n777 ) , .ZN( us23_n866 ) );
  NOR2_X1 us23_U128 (.ZN( us23_n494 ) , .A1( us23_n677 ) , .A2( us23_n693 ) );
  NOR2_X1 us23_U129 (.ZN( us23_n747 ) , .A1( us23_n860 ) , .A2( us23_n861 ) );
  OR4_X1 us23_U13 (.A4( us23_n441 ) , .A2( us23_n442 ) , .A1( us23_n443 ) , .ZN( us23_n444 ) , .A3( us23_n552 ) );
  AOI222_X1 us23_U130 (.ZN( us23_n512 ) , .C1( us23_n831 ) , .B2( us23_n836 ) , .A2( us23_n842 ) , .C2( us23_n861 ) , .B1( us23_n862 ) , .A1( us23_n865 ) );
  NOR4_X1 us23_U131 (.A4( us23_n508 ) , .A2( us23_n509 ) , .A1( us23_n510 ) , .ZN( us23_n511 ) , .A3( us23_n669 ) );
  INV_X1 us23_U132 (.A( us23_n504 ) , .ZN( us23_n870 ) );
  INV_X1 us23_U133 (.A( us23_n761 ) , .ZN( us23_n829 ) );
  NOR2_X1 us23_U134 (.ZN( us23_n646 ) , .A1( us23_n853 ) , .A2( us23_n867 ) );
  OR4_X1 us23_U135 (.A4( us23_n579 ) , .A3( us23_n580 ) , .A2( us23_n581 ) , .A1( us23_n582 ) , .ZN( us23_n583 ) );
  OR4_X1 us23_U136 (.A4( us23_n681 ) , .A3( us23_n682 ) , .A2( us23_n683 ) , .A1( us23_n684 ) , .ZN( us23_n689 ) );
  OR4_X1 us23_U137 (.A4( us23_n565 ) , .A3( us23_n566 ) , .A2( us23_n567 ) , .ZN( us23_n571 ) , .A1( us23_n664 ) );
  OR4_X1 us23_U138 (.A4( us23_n517 ) , .A2( us23_n518 ) , .A1( us23_n519 ) , .ZN( us23_n521 ) , .A3( us23_n820 ) );
  OR4_X1 us23_U139 (.ZN( us23_n465 ) , .A4( us23_n517 ) , .A3( us23_n528 ) , .A2( us23_n577 ) , .A1( us23_n711 ) );
  INV_X1 us23_U14 (.A( us23_n612 ) , .ZN( us23_n874 ) );
  NAND2_X1 us23_U140 (.ZN( us23_n612 ) , .A2( us23_n836 ) , .A1( us23_n872 ) );
  OR3_X1 us23_U141 (.A3( us23_n505 ) , .A2( us23_n506 ) , .A1( us23_n507 ) , .ZN( us23_n510 ) );
  AOI221_X1 us23_U142 (.A( us23_n712 ) , .B2( us23_n713 ) , .ZN( us23_n719 ) , .C1( us23_n831 ) , .B1( us23_n838 ) , .C2( us23_n862 ) );
  OR2_X1 us23_U143 (.A2( us23_n710 ) , .A1( us23_n711 ) , .ZN( us23_n712 ) );
  INV_X1 us23_U144 (.A( us23_n462 ) , .ZN( us23_n863 ) );
  OAI21_X1 us23_U145 (.ZN( us23_n462 ) , .B1( us23_n808 ) , .A( us23_n833 ) , .B2( us23_n850 ) );
  INV_X1 us23_U146 (.A( us23_n753 ) , .ZN( us23_n868 ) );
  OAI21_X1 us23_U147 (.B1( us23_n752 ) , .ZN( us23_n753 ) , .A( us23_n844 ) , .B2( us23_n867 ) );
  INV_X1 us23_U148 (.A( us23_n671 ) , .ZN( us23_n858 ) );
  AOI21_X1 us23_U149 (.A( us23_n669 ) , .B1( us23_n670 ) , .ZN( us23_n671 ) , .B2( us23_n855 ) );
  INV_X1 us23_U15 (.A( us23_n748 ) , .ZN( us23_n862 ) );
  AOI222_X1 us23_U150 (.ZN( us23_n659 ) , .A2( us23_n838 ) , .B1( us23_n840 ) , .C2( us23_n844 ) , .A1( us23_n859 ) , .C1( us23_n862 ) , .B2( us23_n869 ) );
  INV_X1 us23_U151 (.A( us23_n646 ) , .ZN( us23_n869 ) );
  OAI222_X1 us23_U152 (.B2( us23_n707 ) , .ZN( us23_n708 ) , .C2( us23_n723 ) , .B1( us23_n746 ) , .A1( us23_n805 ) , .C1( us23_n813 ) , .A2( us23_n814 ) );
  OAI222_X1 us23_U153 (.A2( us23_n668 ) , .ZN( us23_n673 ) , .B1( us23_n746 ) , .B2( us23_n783 ) , .C2( us23_n787 ) , .C1( us23_n814 ) , .A1( us23_n816 ) );
  NAND2_X1 us23_U154 (.A1( us23_n446 ) , .A2( us23_n464 ) , .ZN( us23_n748 ) );
  NOR4_X1 us23_U155 (.A2( us23_n490 ) , .A1( us23_n491 ) , .ZN( us23_n492 ) , .A3( us23_n579 ) , .A4( us23_n611 ) );
  OR4_X1 us23_U156 (.ZN( us23_n491 ) , .A4( us23_n533 ) , .A2( us23_n546 ) , .A1( us23_n558 ) , .A3( us23_n631 ) );
  OAI22_X1 us23_U157 (.B1( us23_n489 ) , .ZN( us23_n490 ) , .A1( us23_n685 ) , .A2( us23_n762 ) , .B2( us23_n816 ) );
  NOR3_X1 us23_U158 (.ZN( us23_n489 ) , .A1( us23_n781 ) , .A2( us23_n849 ) , .A3( us23_n862 ) );
  AOI22_X1 us23_U159 (.ZN( us23_n695 ) , .A1( us23_n829 ) , .B2( us23_n842 ) , .A2( us23_n864 ) , .B1( us23_n867 ) );
  AOI222_X1 us23_U16 (.ZN( us23_n604 ) , .B2( us23_n670 ) , .B1( us23_n752 ) , .C2( us23_n830 ) , .A1( us23_n832 ) , .A2( us23_n861 ) , .C1( us23_n862 ) );
  AOI21_X1 us23_U160 (.ZN( us23_n638 ) , .B2( us23_n748 ) , .A( us23_n787 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U161 (.ZN( us23_n639 ) , .B2( us23_n746 ) , .A( us23_n791 ) , .B1( us23_n802 ) );
  AOI21_X1 us23_U162 (.ZN( us23_n640 ) , .B1( us23_n679 ) , .A( us23_n790 ) , .B2( us23_n816 ) );
  INV_X1 us23_U163 (.A( us23_n729 ) , .ZN( us23_n838 ) );
  AOI221_X1 us23_U164 (.A( us23_n763 ) , .ZN( us23_n773 ) , .C2( us23_n809 ) , .B2( us23_n834 ) , .C1( us23_n854 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U165 (.B2( us23_n762 ) , .ZN( us23_n763 ) , .A( us23_n787 ) , .B1( us23_n791 ) );
  INV_X1 us23_U166 (.A( us23_n760 ) , .ZN( us23_n834 ) );
  AOI221_X1 us23_U167 (.A( us23_n449 ) , .ZN( us23_n458 ) , .C2( us23_n752 ) , .B1( us23_n831 ) , .C1( us23_n841 ) , .B2( us23_n860 ) );
  AOI21_X1 us23_U168 (.ZN( us23_n449 ) , .B2( us23_n791 ) , .A( us23_n802 ) , .B1( us23_n814 ) );
  AOI221_X1 us23_U169 (.A( us23_n482 ) , .ZN( us23_n487 ) , .B1( us23_n830 ) , .C2( us23_n843 ) , .C1( us23_n851 ) , .B2( us23_n861 ) );
  AOI222_X1 us23_U17 (.ZN( us23_n562 ) , .B1( us23_n829 ) , .C1( us23_n840 ) , .A2( us23_n842 ) , .A1( us23_n853 ) , .B2( us23_n862 ) , .C2( us23_n872 ) );
  OAI22_X1 us23_U170 (.ZN( us23_n482 ) , .A1( us23_n707 ) , .B2( us23_n784 ) , .A2( us23_n805 ) , .B1( us23_n811 ) );
  INV_X1 us23_U171 (.A( us23_n789 ) , .ZN( us23_n831 ) );
  NAND2_X1 us23_U172 (.A1( us23_n450 ) , .A2( us23_n452 ) , .ZN( us23_n761 ) );
  INV_X1 us23_U173 (.A( us23_n783 ) , .ZN( us23_n860 ) );
  INV_X1 us23_U174 (.A( us23_n785 ) , .ZN( us23_n861 ) );
  INV_X1 us23_U175 (.A( us23_n815 ) , .ZN( us23_n830 ) );
  OAI22_X1 us23_U176 (.ZN( us23_n709 ) , .A2( us23_n727 ) , .B2( us23_n728 ) , .A1( us23_n743 ) , .B1( us23_n812 ) );
  OAI22_X1 us23_U177 (.ZN( us23_n623 ) , .B1( us23_n668 ) , .B2( us23_n746 ) , .A1( us23_n814 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U178 (.ZN( us23_n587 ) , .A2( us23_n746 ) , .B2( us23_n761 ) , .A1( us23_n762 ) , .B1( us23_n783 ) );
  INV_X1 us23_U179 (.A( us23_n743 ) , .ZN( us23_n836 ) );
  NOR4_X1 us23_U18 (.ZN( us23_n472 ) , .A2( us23_n520 ) , .A4( us23_n593 ) , .A1( us23_n608 ) , .A3( us23_n628 ) );
  INV_X1 us23_U180 (.A( us23_n787 ) , .ZN( us23_n844 ) );
  OAI22_X1 us23_U181 (.A1( us23_n723 ) , .ZN( us23_n725 ) , .B2( us23_n749 ) , .B1( us23_n811 ) , .A2( us23_n815 ) );
  OAI22_X1 us23_U182 (.B2( us23_n778 ) , .B1( us23_n779 ) , .ZN( us23_n780 ) , .A2( us23_n813 ) , .A1( us23_n814 ) );
  OAI22_X1 us23_U183 (.ZN( us23_n680 ) , .A1( us23_n698 ) , .A2( us23_n729 ) , .B2( us23_n783 ) , .B1( us23_n816 ) );
  OAI22_X1 us23_U184 (.B2( us23_n749 ) , .B1( us23_n750 ) , .A1( us23_n751 ) , .ZN( us23_n755 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U185 (.ZN( us23_n750 ) , .A2( us23_n851 ) , .A1( us23_n859 ) );
  NOR3_X1 us23_U186 (.ZN( us23_n751 ) , .A2( us23_n852 ) , .A1( us23_n862 ) , .A3( us23_n864 ) );
  OAI22_X1 us23_U187 (.B2( us23_n743 ) , .ZN( us23_n745 ) , .A2( us23_n761 ) , .B1( us23_n779 ) , .A1( us23_n791 ) );
  INV_X1 us23_U188 (.A( us23_n802 ) , .ZN( us23_n842 ) );
  INV_X1 us23_U189 (.A( us23_n813 ) , .ZN( us23_n832 ) );
  NOR4_X1 us23_U19 (.A4( us23_n531 ) , .A3( us23_n532 ) , .A2( us23_n533 ) , .ZN( us23_n534 ) , .A1( us23_n819 ) );
  INV_X1 us23_U190 (.A( us23_n804 ) , .ZN( us23_n859 ) );
  OAI22_X1 us23_U191 (.B2( us23_n802 ) , .B1( us23_n803 ) , .A2( us23_n804 ) , .A1( us23_n805 ) , .ZN( us23_n807 ) );
  OAI22_X1 us23_U192 (.ZN( us23_n495 ) , .A2( us23_n743 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U193 (.ZN( us23_n488 ) , .A1( us23_n723 ) , .B2( us23_n727 ) , .B1( us23_n729 ) , .A2( us23_n778 ) );
  INV_X1 us23_U194 (.A( us23_n668 ) , .ZN( us23_n864 ) );
  OAI22_X1 us23_U195 (.ZN( us23_n694 ) , .A2( us23_n729 ) , .A1( us23_n779 ) , .B1( us23_n790 ) , .B2( us23_n816 ) );
  OAI22_X1 us23_U196 (.ZN( us23_n636 ) , .A1( us23_n698 ) , .B2( us23_n727 ) , .A2( us23_n761 ) , .B1( us23_n815 ) );
  NOR2_X1 us23_U197 (.A1( us23_n696 ) , .ZN( us23_n769 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U198 (.ZN( us23_n714 ) , .A1( us23_n804 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U199 (.ZN( us23_n717 ) , .A2( us23_n723 ) , .A1( us23_n743 ) );
  NOR4_X1 us23_U20 (.ZN( us23_n478 ) , .A1( us23_n519 ) , .A4( us23_n556 ) , .A3( us23_n581 ) , .A2( us23_n629 ) );
  NOR2_X1 us23_U200 (.ZN( us23_n545 ) , .A2( us23_n779 ) , .A1( us23_n813 ) );
  INV_X1 us23_U201 (.A( us23_n749 ) , .ZN( us23_n841 ) );
  NOR2_X1 us23_U202 (.ZN( us23_n651 ) , .A1( us23_n668 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U203 (.ZN( us23_n531 ) , .A2( us23_n748 ) , .A1( us23_n749 ) );
  NOR2_X1 us23_U204 (.ZN( us23_n576 ) , .A2( us23_n698 ) , .A1( us23_n813 ) );
  NOR2_X1 us23_U205 (.ZN( us23_n599 ) , .A2( us23_n696 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U206 (.A1( us23_n668 ) , .ZN( us23_n672 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U207 (.ZN( us23_n601 ) , .A1( us23_n668 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U208 (.A1( us23_n668 ) , .ZN( us23_n687 ) , .A2( us23_n815 ) );
  NOR2_X1 us23_U209 (.ZN( us23_n628 ) , .A2( us23_n727 ) , .A1( us23_n784 ) );
  NOR4_X1 us23_U21 (.A4( us23_n540 ) , .A3( us23_n541 ) , .A2( us23_n542 ) , .ZN( us23_n549 ) , .A1( us23_n687 ) );
  NOR2_X1 us23_U210 (.ZN( us23_n614 ) , .A1( us23_n784 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U211 (.A2( us23_n743 ) , .ZN( us23_n754 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U212 (.A1( us23_n668 ) , .ZN( us23_n765 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U213 (.ZN( us23_n734 ) , .A2( us23_n802 ) , .A1( us23_n804 ) );
  NOR2_X1 us23_U214 (.A1( us23_n698 ) , .ZN( us23_n767 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U215 (.A2( us23_n743 ) , .ZN( us23_n768 ) , .A1( us23_n811 ) );
  NOR2_X1 us23_U216 (.ZN( us23_n530 ) , .A2( us23_n779 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U217 (.ZN( us23_n526 ) , .A1( us23_n668 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U218 (.ZN( us23_n540 ) , .A2( us23_n696 ) , .A1( us23_n698 ) );
  NOR2_X1 us23_U219 (.ZN( us23_n598 ) , .A2( us23_n790 ) , .A1( us23_n815 ) );
  NOR2_X1 us23_U22 (.ZN( us23_n679 ) , .A2( us23_n833 ) , .A1( us23_n838 ) );
  NOR2_X1 us23_U220 (.ZN( us23_n627 ) , .A2( us23_n668 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U221 (.ZN( us23_n600 ) , .A2( us23_n779 ) , .A1( us23_n802 ) );
  INV_X1 us23_U222 (.A( us23_n746 ) , .ZN( us23_n833 ) );
  NOR2_X1 us23_U223 (.ZN( us23_n610 ) , .A2( us23_n779 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U224 (.ZN( us23_n527 ) , .A2( us23_n723 ) , .A1( us23_n802 ) );
  NOR2_X1 us23_U225 (.ZN( us23_n609 ) , .A1( us23_n783 ) , .A2( us23_n815 ) );
  INV_X1 us23_U226 (.A( us23_n791 ) , .ZN( us23_n850 ) );
  NOR2_X1 us23_U227 (.ZN( us23_n650 ) , .A1( us23_n783 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U228 (.A2( us23_n707 ) , .A1( us23_n749 ) , .ZN( us23_n770 ) );
  NOR2_X1 us23_U229 (.ZN( us23_n666 ) , .A1( us23_n749 ) , .A2( us23_n814 ) );
  AOI222_X1 us23_U23 (.ZN( us23_n468 ) , .B1( us23_n831 ) , .A1( us23_n838 ) , .C1( us23_n841 ) , .C2( us23_n850 ) , .A2( us23_n854 ) , .B2( us23_n864 ) );
  NOR2_X1 us23_U230 (.ZN( us23_n554 ) , .A1( us23_n749 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U231 (.ZN( us23_n507 ) , .A2( us23_n779 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U232 (.ZN( us23_n542 ) , .A2( us23_n707 ) , .A1( us23_n784 ) );
  NOR2_X1 us23_U233 (.ZN( us23_n663 ) , .A1( us23_n784 ) , .A2( us23_n790 ) );
  OAI22_X1 us23_U234 (.B1( us23_n439 ) , .ZN( us23_n443 ) , .A2( us23_n727 ) , .A1( us23_n743 ) , .B2( us23_n748 ) );
  NOR3_X1 us23_U235 (.ZN( us23_n439 ) , .A2( us23_n835 ) , .A3( us23_n836 ) , .A1( us23_n845 ) );
  NOR2_X1 us23_U236 (.A2( us23_n696 ) , .ZN( us23_n715 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U237 (.ZN( us23_n506 ) , .A1( us23_n811 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U238 (.ZN( us23_n593 ) , .A2( us23_n696 ) , .A1( us23_n727 ) );
  NOR2_X1 us23_U239 (.ZN( us23_n661 ) , .A2( us23_n696 ) , .A1( us23_n728 ) );
  NOR4_X1 us23_U24 (.A1( us23_n465 ) , .ZN( us23_n466 ) , .A4( us23_n541 ) , .A2( us23_n553 ) , .A3( us23_n613 ) );
  NOR2_X1 us23_U240 (.ZN( us23_n556 ) , .A1( us23_n791 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U241 (.ZN( us23_n544 ) , .A1( us23_n748 ) , .A2( us23_n813 ) );
  NOR2_X1 us23_U242 (.ZN( us23_n555 ) , .A1( us23_n761 ) , .A2( us23_n804 ) );
  NOR2_X1 us23_U243 (.ZN( us23_n529 ) , .A2( us23_n743 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U244 (.A2( us23_n696 ) , .A1( us23_n779 ) , .ZN( us23_n819 ) );
  NOR2_X1 us23_U245 (.ZN( us23_n508 ) , .A1( us23_n728 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U246 (.ZN( us23_n665 ) , .A1( us23_n727 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U247 (.ZN( us23_n543 ) , .A2( us23_n784 ) , .A1( us23_n791 ) );
  NOR2_X1 us23_U248 (.A1( us23_n748 ) , .ZN( us23_n766 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U249 (.ZN( us23_n613 ) , .A1( us23_n761 ) , .A2( us23_n811 ) );
  AOI221_X1 us23_U25 (.ZN( us23_n467 ) , .C2( us23_n713 ) , .B2( us23_n830 ) , .C1( us23_n844 ) , .B1( us23_n859 ) , .A( us23_n863 ) );
  NOR2_X1 us23_U250 (.ZN( us23_n515 ) , .A1( us23_n707 ) , .A2( us23_n743 ) );
  NOR2_X1 us23_U251 (.ZN( us23_n630 ) , .A1( us23_n723 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U252 (.ZN( us23_n569 ) , .A1( us23_n727 ) , .A2( us23_n805 ) );
  NOR2_X1 us23_U253 (.ZN( us23_n557 ) , .A1( us23_n707 ) , .A2( us23_n815 ) );
  INV_X1 us23_U254 (.A( us23_n762 ) , .ZN( us23_n865 ) );
  NOR2_X1 us23_U255 (.ZN( us23_n653 ) , .A1( us23_n727 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U256 (.ZN( us23_n516 ) , .A1( us23_n707 ) , .A2( us23_n802 ) );
  NOR2_X1 us23_U257 (.ZN( us23_n520 ) , .A1( us23_n789 ) , .A2( us23_n811 ) );
  NOR2_X1 us23_U258 (.ZN( us23_n662 ) , .A1( us23_n728 ) , .A2( us23_n784 ) );
  NOR2_X1 us23_U259 (.ZN( us23_n654 ) , .A1( us23_n789 ) , .A2( us23_n814 ) );
  NOR4_X1 us23_U26 (.A4( us23_n664 ) , .A3( us23_n665 ) , .A2( us23_n666 ) , .A1( us23_n667 ) , .ZN( us23_n675 ) );
  NOR2_X1 us23_U260 (.ZN( us23_n629 ) , .A1( us23_n746 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U261 (.ZN( us23_n667 ) , .A2( us23_n707 ) , .A1( us23_n789 ) );
  NOR2_X1 us23_U262 (.ZN( us23_n669 ) , .A1( us23_n789 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U263 (.ZN( us23_n570 ) , .B2( us23_n696 ) , .B1( us23_n805 ) , .A( us23_n811 ) );
  NOR2_X1 us23_U264 (.ZN( us23_n541 ) , .A1( us23_n761 ) , .A2( us23_n790 ) );
  NOR2_X1 us23_U265 (.ZN( us23_n655 ) , .A1( us23_n746 ) , .A2( us23_n779 ) );
  INV_X1 us23_U266 (.A( us23_n805 ) , .ZN( us23_n840 ) );
  NOR2_X1 us23_U267 (.ZN( us23_n608 ) , .A2( us23_n723 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U268 (.A( us23_n814 ) , .B2( us23_n815 ) , .B1( us23_n816 ) , .ZN( us23_n817 ) );
  AOI21_X1 us23_U269 (.ZN( us23_n625 ) , .B2( us23_n668 ) , .A( us23_n789 ) , .B1( us23_n790 ) );
  NOR4_X1 us23_U27 (.A4( us23_n660 ) , .A3( us23_n661 ) , .A2( us23_n662 ) , .A1( us23_n663 ) , .ZN( us23_n676 ) );
  NOR2_X1 us23_U270 (.ZN( us23_n660 ) , .A1( us23_n728 ) , .A2( us23_n789 ) );
  INV_X1 us23_U271 (.A( us23_n811 ) , .ZN( us23_n853 ) );
  NOR2_X1 us23_U272 (.ZN( us23_n578 ) , .A2( us23_n707 ) , .A1( us23_n729 ) );
  NOR2_X1 us23_U273 (.ZN( us23_n532 ) , .A2( us23_n723 ) , .A1( us23_n729 ) );
  AOI21_X1 us23_U274 (.ZN( us23_n498 ) , .B1( us23_n679 ) , .A( us23_n811 ) , .B2( us23_n815 ) );
  AOI21_X1 us23_U275 (.ZN( us23_n551 ) , .B1( us23_n668 ) , .A( us23_n696 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U276 (.ZN( us23_n581 ) , .A1( us23_n743 ) , .A2( us23_n814 ) );
  NOR2_X1 us23_U277 (.A2( us23_n707 ) , .A1( us23_n761 ) , .ZN( us23_n793 ) );
  AOI21_X1 us23_U278 (.B1( us23_n624 ) , .ZN( us23_n626 ) , .A( us23_n762 ) , .B2( us23_n813 ) );
  AOI21_X1 us23_U279 (.ZN( us23_n514 ) , .A( us23_n728 ) , .B1( us23_n749 ) , .B2( us23_n802 ) );
  NOR4_X1 us23_U28 (.A3( us23_n672 ) , .A1( us23_n673 ) , .ZN( us23_n674 ) , .A4( us23_n714 ) , .A2( us23_n858 ) );
  AOI21_X1 us23_U280 (.A( us23_n811 ) , .B2( us23_n812 ) , .B1( us23_n813 ) , .ZN( us23_n818 ) );
  AOI21_X1 us23_U281 (.ZN( us23_n477 ) , .B2( us23_n696 ) , .A( us23_n748 ) , .B1( us23_n778 ) );
  AOI21_X1 us23_U282 (.ZN( us23_n509 ) , .B2( us23_n668 ) , .A( us23_n729 ) , .B1( us23_n814 ) );
  NOR2_X1 us23_U283 (.ZN( us23_n505 ) , .A2( us23_n727 ) , .A1( us23_n761 ) );
  AOI21_X1 us23_U284 (.ZN( us23_n591 ) , .B1( us23_n727 ) , .B2( us23_n783 ) , .A( us23_n789 ) );
  NOR2_X1 us23_U285 (.ZN( us23_n518 ) , .A2( us23_n698 ) , .A1( us23_n815 ) );
  AOI21_X1 us23_U286 (.ZN( us23_n592 ) , .B1( us23_n749 ) , .A( us23_n791 ) , .B2( us23_n812 ) );
  AOI21_X1 us23_U287 (.ZN( us23_n649 ) , .A( us23_n778 ) , .B1( us23_n791 ) , .B2( us23_n804 ) );
  NOR2_X1 us23_U288 (.ZN( us23_n580 ) , .A1( us23_n668 ) , .A2( us23_n787 ) );
  NOR2_X1 us23_U289 (.ZN( us23_n519 ) , .A2( us23_n707 ) , .A1( us23_n813 ) );
  NOR4_X1 us23_U29 (.A4( us23_n513 ) , .A3( us23_n514 ) , .A2( us23_n515 ) , .A1( us23_n516 ) , .ZN( us23_n523 ) );
  AOI21_X1 us23_U290 (.ZN( us23_n476 ) , .A( us23_n668 ) , .B1( us23_n749 ) , .B2( us23_n805 ) );
  NOR2_X1 us23_U291 (.ZN( us23_n558 ) , .A2( us23_n790 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U292 (.ZN( us23_n647 ) , .A( us23_n761 ) , .B2( us23_n783 ) , .B1( us23_n791 ) );
  AOI21_X1 us23_U293 (.ZN( us23_n622 ) , .B1( us23_n698 ) , .A( us23_n778 ) , .B2( us23_n783 ) );
  AOI21_X1 us23_U294 (.ZN( us23_n588 ) , .B2( us23_n698 ) , .B1( us23_n814 ) , .A( us23_n816 ) );
  NOR2_X1 us23_U295 (.ZN( us23_n552 ) , .A2( us23_n743 ) , .A1( us23_n783 ) );
  NOR2_X1 us23_U296 (.ZN( us23_n682 ) , .A2( us23_n698 ) , .A1( us23_n802 ) );
  AOI21_X1 us23_U297 (.B1( us23_n698 ) , .ZN( us23_n699 ) , .A( us23_n731 ) , .B2( us23_n762 ) );
  AOI21_X1 us23_U298 (.ZN( us23_n590 ) , .B2( us23_n762 ) , .A( us23_n784 ) , .B1( us23_n811 ) );
  AOI21_X1 us23_U299 (.ZN( us23_n538 ) , .B2( us23_n811 ) , .A( us23_n813 ) , .B1( us23_n814 ) );
  NOR3_X1 us23_U3 (.ZN( us23_n597 ) , .A1( us23_n607 ) , .A3( us23_n722 ) , .A2( us23_n741 ) );
  AOI222_X1 us23_U30 (.ZN( us23_n524 ) , .A1( us23_n833 ) , .B2( us23_n836 ) , .C1( us23_n843 ) , .C2( us23_n849 ) , .A2( us23_n851 ) , .B1( us23_n865 ) );
  AOI21_X1 us23_U300 (.ZN( us23_n539 ) , .A( us23_n762 ) , .B2( us23_n778 ) , .B1( us23_n816 ) );
  NOR2_X1 us23_U301 (.ZN( us23_n546 ) , .A1( us23_n698 ) , .A2( us23_n743 ) );
  INV_X1 us23_U302 (.A( us23_n812 ) , .ZN( us23_n835 ) );
  INV_X1 us23_U303 (.A( us23_n727 ) , .ZN( us23_n851 ) );
  AOI21_X1 us23_U304 (.ZN( us23_n648 ) , .B1( us23_n728 ) , .B2( us23_n762 ) , .A( us23_n812 ) );
  INV_X1 us23_U305 (.A( us23_n790 ) , .ZN( us23_n872 ) );
  OAI221_X1 us23_U306 (.A( us23_n726 ) , .C2( us23_n727 ) , .B2( us23_n728 ) , .B1( us23_n729 ) , .ZN( us23_n736 ) , .C1( us23_n816 ) );
  AOI22_X1 us23_U307 (.ZN( us23_n726 ) , .B1( us23_n831 ) , .A2( us23_n837 ) , .A1( us23_n862 ) , .B2( us23_n865 ) );
  AOI21_X1 us23_U308 (.ZN( us23_n497 ) , .A( us23_n723 ) , .B2( us23_n761 ) , .B1( us23_n813 ) );
  NOR2_X1 us23_U309 (.ZN( us23_n565 ) , .A2( us23_n696 ) , .A1( us23_n762 ) );
  NOR4_X1 us23_U31 (.A3( us23_n520 ) , .A1( us23_n521 ) , .ZN( us23_n522 ) , .A2( us23_n672 ) , .A4( us23_n768 ) );
  INV_X1 us23_U310 (.A( us23_n698 ) , .ZN( us23_n852 ) );
  AOI21_X1 us23_U311 (.ZN( us23_n568 ) , .B1( us23_n749 ) , .B2( us23_n761 ) , .A( us23_n779 ) );
  AOI21_X1 us23_U312 (.ZN( us23_n513 ) , .A( us23_n778 ) , .B2( us23_n791 ) , .B1( us23_n811 ) );
  NOR2_X1 us23_U313 (.ZN( us23_n579 ) , .A2( us23_n696 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U314 (.ZN( us23_n684 ) , .A1( us23_n728 ) , .A2( us23_n815 ) );
  AOI21_X1 us23_U315 (.ZN( us23_n563 ) , .B1( us23_n723 ) , .A( us23_n778 ) , .B2( us23_n790 ) );
  AOI21_X1 us23_U316 (.ZN( us23_n496 ) , .A( us23_n778 ) , .B2( us23_n790 ) , .B1( us23_n803 ) );
  INV_X1 us23_U317 (.A( us23_n728 ) , .ZN( us23_n867 ) );
  NOR2_X1 us23_U318 (.ZN( us23_n664 ) , .A1( us23_n779 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U319 (.ZN( us23_n631 ) , .A2( us23_n696 ) , .A1( us23_n723 ) );
  AOI221_X1 us23_U32 (.A( us23_n780 ) , .ZN( us23_n797 ) , .C2( us23_n836 ) , .B2( us23_n837 ) , .B1( us23_n864 ) , .C1( us23_n865 ) );
  NOR2_X1 us23_U320 (.ZN( us23_n528 ) , .A1( us23_n707 ) , .A2( us23_n778 ) );
  NOR2_X1 us23_U321 (.ZN( us23_n577 ) , .A1( us23_n707 ) , .A2( us23_n812 ) );
  AOI21_X1 us23_U322 (.A( us23_n789 ) , .B2( us23_n790 ) , .B1( us23_n791 ) , .ZN( us23_n792 ) );
  AOI21_X1 us23_U323 (.ZN( us23_n688 ) , .B2( us23_n748 ) , .B1( us23_n762 ) , .A( us23_n805 ) );
  NOR2_X1 us23_U324 (.ZN( us23_n683 ) , .A1( us23_n790 ) , .A2( us23_n812 ) );
  NOR2_X1 us23_U325 (.ZN( us23_n566 ) , .A1( us23_n746 ) , .A2( us23_n804 ) );
  NAND2_X1 us23_U326 (.ZN( us23_n752 ) , .A1( us23_n762 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U327 (.A( us23_n732 ) , .ZN( us23_n733 ) , .B2( us23_n779 ) , .B1( us23_n791 ) );
  NOR2_X1 us23_U328 (.A2( us23_n812 ) , .A1( us23_n814 ) , .ZN( us23_n820 ) );
  NOR2_X1 us23_U329 (.ZN( us23_n710 ) , .A1( us23_n761 ) , .A2( us23_n762 ) );
  NOR4_X1 us23_U33 (.A4( us23_n792 ) , .A3( us23_n793 ) , .A2( us23_n794 ) , .A1( us23_n795 ) , .ZN( us23_n796 ) );
  NOR2_X1 us23_U330 (.ZN( us23_n641 ) , .A2( us23_n787 ) , .A1( us23_n790 ) );
  NOR2_X1 us23_U331 (.ZN( us23_n582 ) , .A1( us23_n791 ) , .A2( us23_n816 ) );
  NOR2_X1 us23_U332 (.ZN( us23_n681 ) , .A2( us23_n707 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U333 (.ZN( us23_n533 ) , .A1( us23_n723 ) , .A2( us23_n787 ) );
  AOI21_X1 us23_U334 (.B1( us23_n685 ) , .ZN( us23_n686 ) , .A( us23_n727 ) , .B2( us23_n760 ) );
  INV_X1 us23_U335 (.A( us23_n696 ) , .ZN( us23_n837 ) );
  INV_X1 us23_U336 (.A( us23_n814 ) , .ZN( us23_n854 ) );
  NOR2_X1 us23_U337 (.ZN( us23_n567 ) , .A1( us23_n728 ) , .A2( us23_n761 ) );
  AOI21_X1 us23_U338 (.ZN( us23_n441 ) , .A( us23_n698 ) , .B1( us23_n732 ) , .B2( us23_n749 ) );
  OAI21_X1 us23_U339 (.A( us23_n730 ) , .B1( us23_n731 ) , .ZN( us23_n735 ) , .B2( us23_n804 ) );
  NOR4_X1 us23_U34 (.A4( us23_n775 ) , .A3( us23_n776 ) , .A1( us23_n777 ) , .ZN( us23_n798 ) , .A2( us23_n800 ) );
  OAI21_X1 us23_U340 (.ZN( us23_n730 ) , .A( us23_n832 ) , .B2( us23_n851 ) , .B1( us23_n872 ) );
  OAI21_X1 us23_U341 (.A( us23_n697 ) , .ZN( us23_n701 ) , .B2( us23_n749 ) , .B1( us23_n803 ) );
  OAI21_X1 us23_U342 (.ZN( us23_n697 ) , .B2( us23_n832 ) , .B1( us23_n837 ) , .A( us23_n859 ) );
  OAI21_X1 us23_U343 (.A( us23_n612 ) , .ZN( us23_n615 ) , .B1( us23_n624 ) , .B2( us23_n783 ) );
  INV_X1 us23_U344 (.A( us23_n779 ) , .ZN( us23_n849 ) );
  AOI22_X1 us23_U345 (.A2( us23_n781 ) , .ZN( us23_n782 ) , .B2( us23_n830 ) , .A1( us23_n833 ) , .B1( us23_n862 ) );
  NAND2_X1 us23_U346 (.ZN( us23_n670 ) , .A1( us23_n805 ) , .A2( us23_n815 ) );
  OAI21_X1 us23_U347 (.A( us23_n786 ) , .B2( us23_n787 ) , .B1( us23_n788 ) , .ZN( us23_n794 ) );
  OAI21_X1 us23_U348 (.ZN( us23_n786 ) , .A( us23_n838 ) , .B1( us23_n862 ) , .B2( us23_n872 ) );
  NAND2_X1 us23_U349 (.A1( us23_n728 ) , .A2( us23_n783 ) , .ZN( us23_n810 ) );
  NOR4_X1 us23_U35 (.A4( us23_n733 ) , .A3( us23_n734 ) , .A2( us23_n735 ) , .A1( us23_n736 ) , .ZN( us23_n737 ) );
  NOR2_X1 us23_U350 (.ZN( us23_n483 ) , .A1( us23_n787 ) , .A2( us23_n804 ) );
  AOI21_X1 us23_U351 (.ZN( us23_n442 ) , .B1( us23_n788 ) , .B2( us23_n790 ) , .A( us23_n813 ) );
  NAND2_X1 us23_U352 (.A2( us23_n761 ) , .A1( us23_n805 ) , .ZN( us23_n809 ) );
  NOR2_X1 us23_U353 (.ZN( us23_n469 ) , .A2( us23_n778 ) , .A1( us23_n814 ) );
  NAND2_X1 us23_U354 (.A1( us23_n698 ) , .A2( us23_n728 ) , .ZN( us23_n781 ) );
  NOR2_X1 us23_U355 (.ZN( us23_n711 ) , .A2( us23_n723 ) , .A1( us23_n789 ) );
  INV_X1 us23_U356 (.A( us23_n784 ) , .ZN( us23_n845 ) );
  NOR2_X1 us23_U357 (.ZN( us23_n525 ) , .A1( us23_n723 ) , .A2( us23_n749 ) );
  NOR2_X1 us23_U358 (.ZN( us23_n517 ) , .A1( us23_n707 ) , .A2( us23_n787 ) );
  INV_X1 us23_U359 (.A( us23_n816 ) , .ZN( us23_n843 ) );
  AOI211_X1 us23_U36 (.B( us23_n724 ) , .A( us23_n725 ) , .ZN( us23_n738 ) , .C1( us23_n842 ) , .C2( us23_n854 ) );
  NAND2_X1 us23_U360 (.ZN( us23_n713 ) , .A1( us23_n727 ) , .A2( us23_n779 ) );
  INV_X1 us23_U361 (.A( us23_n723 ) , .ZN( us23_n855 ) );
  AND2_X1 us23_U362 (.ZN( us23_n731 ) , .A1( us23_n778 ) , .A2( us23_n784 ) );
  NAND2_X1 us23_U363 (.A2( us23_n460 ) , .A1( us23_n470 ) , .ZN( us23_n696 ) );
  NAND2_X1 us23_U364 (.A1( us23_n451 ) , .A2( us23_n464 ) , .ZN( us23_n668 ) );
  NAND2_X1 us23_U365 (.A1( us23_n450 ) , .A2( us23_n470 ) , .ZN( us23_n815 ) );
  NAND2_X1 us23_U366 (.A1( us23_n452 ) , .A2( us23_n460 ) , .ZN( us23_n743 ) );
  NAND2_X1 us23_U367 (.A1( us23_n454 ) , .A2( us23_n470 ) , .ZN( us23_n802 ) );
  NAND2_X1 us23_U368 (.A1( us23_n450 ) , .A2( us23_n453 ) , .ZN( us23_n813 ) );
  NAND2_X1 us23_U369 (.A1( us23_n454 ) , .A2( us23_n461 ) , .ZN( us23_n749 ) );
  NOR3_X1 us23_U37 (.A3( us23_n721 ) , .A1( us23_n722 ) , .ZN( us23_n739 ) , .A2( us23_n740 ) );
  NAND2_X1 us23_U370 (.A1( us23_n446 ) , .A2( us23_n448 ) , .ZN( us23_n804 ) );
  NAND2_X1 us23_U371 (.A1( us23_n453 ) , .A2( us23_n460 ) , .ZN( us23_n812 ) );
  NAND2_X1 us23_U372 (.A2( us23_n440 ) , .A1( us23_n446 ) , .ZN( us23_n783 ) );
  NAND2_X1 us23_U373 (.A2( us23_n453 ) , .A1( us23_n471 ) , .ZN( us23_n778 ) );
  NAND2_X1 us23_U374 (.A2( us23_n452 ) , .A1( us23_n454 ) , .ZN( us23_n805 ) );
  NAND2_X1 us23_U375 (.A1( us23_n452 ) , .A2( us23_n471 ) , .ZN( us23_n784 ) );
  NAND2_X1 us23_U376 (.A1( us23_n440 ) , .A2( us23_n459 ) , .ZN( us23_n698 ) );
  NAND2_X1 us23_U377 (.A2( us23_n463 ) , .A1( us23_n464 ) , .ZN( us23_n811 ) );
  NAND2_X1 us23_U378 (.A2( us23_n448 ) , .A1( us23_n451 ) , .ZN( us23_n762 ) );
  NAND2_X1 us23_U379 (.A1( us23_n461 ) , .A2( us23_n471 ) , .ZN( us23_n787 ) );
  NOR4_X1 us23_U38 (.A3( us23_n754 ) , .A2( us23_n755 ) , .A1( us23_n756 ) , .ZN( us23_n757 ) , .A4( us23_n868 ) );
  NAND2_X1 us23_U380 (.A2( us23_n460 ) , .A1( us23_n461 ) , .ZN( us23_n746 ) );
  NOR2_X1 us23_U381 (.ZN( us23_n464 ) , .A2( us23_n846 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U382 (.ZN( us23_n452 ) , .A1( us23_n825 ) , .A2( us23_n826 ) );
  NAND2_X1 us23_U383 (.A1( us23_n450 ) , .A2( us23_n461 ) , .ZN( us23_n789 ) );
  NOR2_X1 us23_U384 (.ZN( us23_n450 ) , .A1( us23_n827 ) , .A2( us23_n828 ) );
  NAND2_X2 us23_U385 (.A2( us23_n447 ) , .A1( us23_n463 ) , .ZN( us23_n814 ) );
  NAND2_X1 us23_U386 (.A2( us23_n453 ) , .A1( us23_n454 ) , .ZN( us23_n729 ) );
  NAND2_X2 us23_U387 (.A2( us23_n440 ) , .A1( us23_n451 ) , .ZN( us23_n790 ) );
  NAND2_X2 us23_U388 (.A1( us23_n448 ) , .A2( us23_n459 ) , .ZN( us23_n791 ) );
  NAND2_X2 us23_U389 (.A1( us23_n448 ) , .A2( us23_n463 ) , .ZN( us23_n723 ) );
  AOI211_X1 us23_U39 (.B( us23_n744 ) , .A( us23_n745 ) , .ZN( us23_n758 ) , .C1( us23_n831 ) , .C2( us23_n852 ) );
  NAND2_X2 us23_U390 (.A1( us23_n440 ) , .A2( us23_n463 ) , .ZN( us23_n707 ) );
  NAND2_X2 us23_U391 (.A2( us23_n470 ) , .A1( us23_n471 ) , .ZN( us23_n816 ) );
  NAND2_X2 us23_U392 (.A2( us23_n459 ) , .A1( us23_n464 ) , .ZN( us23_n779 ) );
  NOR2_X1 us23_U393 (.ZN( us23_n446 ) , .A2( us23_n848 ) , .A1( us23_n857 ) );
  NAND2_X1 us23_U394 (.A1( us23_n446 ) , .A2( us23_n447 ) , .ZN( us23_n785 ) );
  NAND2_X1 us23_U395 (.A2( us23_n447 ) , .A1( us23_n459 ) , .ZN( us23_n727 ) );
  NAND2_X1 us23_U396 (.A2( us23_n447 ) , .A1( us23_n451 ) , .ZN( us23_n728 ) );
  NOR2_X1 us23_U397 (.A2( sa23_5 ) , .ZN( us23_n447 ) , .A1( us23_n846 ) );
  NOR2_X1 us23_U398 (.A2( sa23_7 ) , .ZN( us23_n459 ) , .A1( us23_n848 ) );
  NOR2_X1 us23_U399 (.A2( sa23_6 ) , .A1( sa23_7 ) , .ZN( us23_n463 ) );
  NOR3_X1 us23_U4 (.A3( us23_n799 ) , .A2( us23_n800 ) , .A1( us23_n801 ) , .ZN( us23_n824 ) );
  NOR3_X1 us23_U40 (.A3( us23_n740 ) , .A2( us23_n741 ) , .A1( us23_n742 ) , .ZN( us23_n759 ) );
  NOR2_X1 us23_U400 (.A2( sa23_4 ) , .ZN( us23_n448 ) , .A1( us23_n847 ) );
  NOR2_X1 us23_U401 (.A2( sa23_4 ) , .A1( sa23_5 ) , .ZN( us23_n440 ) );
  NOR2_X1 us23_U402 (.A2( sa23_6 ) , .ZN( us23_n451 ) , .A1( us23_n857 ) );
  NOR2_X1 us23_U403 (.A2( sa23_1 ) , .ZN( us23_n470 ) , .A1( us23_n825 ) );
  NOR2_X1 us23_U404 (.A2( sa23_2 ) , .A1( sa23_3 ) , .ZN( us23_n471 ) );
  NOR2_X1 us23_U405 (.A2( sa23_2 ) , .ZN( us23_n460 ) , .A1( us23_n828 ) );
  NOR2_X1 us23_U406 (.A2( sa23_0 ) , .ZN( us23_n453 ) , .A1( us23_n826 ) );
  NOR2_X1 us23_U407 (.A2( sa23_0 ) , .A1( sa23_1 ) , .ZN( us23_n461 ) );
  NOR2_X1 us23_U408 (.A2( sa23_3 ) , .ZN( us23_n454 ) , .A1( us23_n827 ) );
  INV_X1 us23_U409 (.A( sa23_6 ) , .ZN( us23_n848 ) );
  NAND4_X1 us23_U41 (.ZN( sa21_sr_3 ) , .A4( us23_n703 ) , .A3( us23_n704 ) , .A2( us23_n705 ) , .A1( us23_n706 ) );
  INV_X1 us23_U410 (.A( sa23_4 ) , .ZN( us23_n846 ) );
  INV_X1 us23_U411 (.A( sa23_1 ) , .ZN( us23_n826 ) );
  INV_X1 us23_U412 (.A( sa23_3 ) , .ZN( us23_n828 ) );
  INV_X1 us23_U413 (.A( sa23_2 ) , .ZN( us23_n827 ) );
  INV_X1 us23_U414 (.A( sa23_0 ) , .ZN( us23_n825 ) );
  INV_X1 us23_U415 (.A( sa23_7 ) , .ZN( us23_n857 ) );
  INV_X1 us23_U416 (.A( sa23_5 ) , .ZN( us23_n847 ) );
  OAI221_X1 us23_U417 (.A( us23_n782 ) , .C2( us23_n783 ) , .B2( us23_n784 ) , .B1( us23_n785 ) , .ZN( us23_n795 ) , .C1( us23_n812 ) );
  OAI222_X1 us23_U418 (.B2( us23_n746 ) , .B1( us23_n747 ) , .A2( us23_n748 ) , .ZN( us23_n756 ) , .C2( us23_n804 ) , .C1( us23_n813 ) , .A1( us23_n816 ) );
  AOI21_X1 us23_U419 (.ZN( us23_n499 ) , .A( us23_n696 ) , .B1( us23_n707 ) , .B2( us23_n785 ) );
  NOR4_X1 us23_U42 (.A4( us23_n699 ) , .A3( us23_n700 ) , .A2( us23_n701 ) , .A1( us23_n702 ) , .ZN( us23_n703 ) );
  OAI221_X1 us23_U420 (.A( us23_n695 ) , .ZN( us23_n702 ) , .C2( us23_n783 ) , .C1( us23_n784 ) , .B1( us23_n785 ) , .B2( us23_n805 ) );
  OAI22_X1 us23_U421 (.ZN( us23_n589 ) , .B1( us23_n729 ) , .B2( us23_n748 ) , .A2( us23_n785 ) , .A1( us23_n802 ) );
  OAI222_X1 us23_U422 (.ZN( us23_n504 ) , .C2( us23_n624 ) , .B2( us23_n646 ) , .B1( us23_n746 ) , .A2( us23_n747 ) , .C1( us23_n804 ) , .A1( us23_n805 ) );
  NOR2_X1 us23_U423 (.ZN( us23_n611 ) , .A1( us23_n778 ) , .A2( us23_n785 ) );
  OAI222_X1 us23_U424 (.ZN( us23_n616 ) , .B1( us23_n696 ) , .C1( us23_n723 ) , .C2( us23_n746 ) , .B2( us23_n785 ) , .A2( us23_n791 ) , .A1( us23_n815 ) );
  NAND2_X1 us23_U425 (.A2( us23_n748 ) , .A1( us23_n785 ) , .ZN( us23_n808 ) );
  AOI21_X1 us23_U426 (.ZN( us23_n575 ) , .B2( us23_n723 ) , .B1( us23_n747 ) , .A( us23_n784 ) );
  NOR2_X1 us23_U427 (.ZN( us23_n716 ) , .A2( us23_n743 ) , .A1( us23_n785 ) );
  NOR2_X1 us23_U428 (.ZN( us23_n652 ) , .A1( us23_n761 ) , .A2( us23_n785 ) );
  NOR2_X1 us23_U429 (.ZN( us23_n553 ) , .A1( us23_n785 ) , .A2( us23_n812 ) );
  AOI211_X1 us23_U43 (.B( us23_n693 ) , .A( us23_n694 ) , .ZN( us23_n704 ) , .C2( us23_n830 ) , .C1( us23_n850 ) );
  NOR2_X1 us23_U430 (.ZN( us23_n700 ) , .A2( us23_n785 ) , .A1( us23_n816 ) );
  NOR2_X1 us23_U431 (.A1( us23_n729 ) , .ZN( us23_n764 ) , .A2( us23_n785 ) );
  NAND2_X1 us23_U432 (.ZN( sa21_sr_2 ) , .A1( us23_n438 ) , .A2( us23_n644 ) );
  NOR3_X1 us23_U433 (.A2( us23_n606 ) , .A1( us23_n607 ) , .ZN( us23_n645 ) , .A3( us23_n721 ) );
  AOI222_X1 us23_U434 (.B2( us23_n637 ) , .ZN( us23_n643 ) , .B1( us23_n840 ) , .A1( us23_n841 ) , .C2( us23_n845 ) , .C1( us23_n862 ) , .A2( us23_n864 ) );
  NOR4_X1 us23_U435 (.A4( us23_n638 ) , .A3( us23_n639 ) , .A2( us23_n640 ) , .A1( us23_n641 ) , .ZN( us23_n642 ) );
  AOI211_X1 us23_U436 (.A( us23_n636 ) , .ZN( us23_n644 ) , .B( us23_n742 ) , .C2( us23_n838 ) , .C1( us23_n853 ) );
  NAND3_X1 us23_U437 (.ZN( sa21_sr_6 ) , .A3( us23_n796 ) , .A2( us23_n797 ) , .A1( us23_n798 ) );
  NAND3_X1 us23_U438 (.ZN( sa21_sr_5 ) , .A3( us23_n757 ) , .A2( us23_n758 ) , .A1( us23_n759 ) );
  NAND3_X1 us23_U439 (.ZN( sa21_sr_4 ) , .A3( us23_n737 ) , .A2( us23_n738 ) , .A1( us23_n739 ) );
  NOR2_X1 us23_U44 (.ZN( us23_n706 ) , .A2( us23_n775 ) , .A1( us23_n799 ) );
  NAND3_X1 us23_U440 (.A3( us23_n674 ) , .A2( us23_n675 ) , .A1( us23_n676 ) , .ZN( us23_n806 ) );
  NAND3_X1 us23_U441 (.ZN( us23_n637 ) , .A3( us23_n707 ) , .A2( us23_n723 ) , .A1( us23_n791 ) );
  NAND3_X1 us23_U442 (.A3( us23_n617 ) , .A2( us23_n618 ) , .A1( us23_n619 ) , .ZN( us23_n724 ) );
  NAND3_X1 us23_U443 (.A3( us23_n584 ) , .A2( us23_n585 ) , .A1( us23_n586 ) , .ZN( us23_n620 ) );
  NAND3_X1 us23_U444 (.ZN( us23_n564 ) , .A3( us23_n679 ) , .A2( us23_n749 ) , .A1( us23_n784 ) );
  NAND3_X1 us23_U445 (.A3( us23_n522 ) , .A2( us23_n523 ) , .A1( us23_n524 ) , .ZN( us23_n741 ) );
  NAND3_X1 us23_U446 (.A3( us23_n511 ) , .A1( us23_n512 ) , .ZN( us23_n607 ) , .A2( us23_n870 ) );
  NAND3_X1 us23_U447 (.A3( us23_n466 ) , .A2( us23_n467 ) , .A1( us23_n468 ) , .ZN( us23_n776 ) );
  NAND4_X1 us23_U448 (.A4( us23_n632 ) , .A3( us23_n633 ) , .A2( us23_n634 ) , .A1( us23_n635 ) , .ZN( us23_n742 ) );
  NOR2_X1 us23_U45 (.ZN( us23_n803 ) , .A1( us23_n853 ) , .A2( us23_n860 ) );
  NAND4_X1 us23_U46 (.ZN( sa21_sr_7 ) , .A4( us23_n821 ) , .A3( us23_n822 ) , .A2( us23_n823 ) , .A1( us23_n824 ) );
  AOI222_X1 us23_U47 (.C2( us23_n808 ) , .B2( us23_n809 ) , .A2( us23_n810 ) , .ZN( us23_n822 ) , .C1( us23_n831 ) , .A1( us23_n838 ) , .B1( us23_n852 ) );
  NOR4_X1 us23_U48 (.A4( us23_n817 ) , .A3( us23_n818 ) , .A2( us23_n819 ) , .A1( us23_n820 ) , .ZN( us23_n821 ) );
  AOI211_X1 us23_U49 (.B( us23_n806 ) , .A( us23_n807 ) , .ZN( us23_n823 ) , .C1( us23_n841 ) , .C2( us23_n849 ) );
  NOR3_X1 us23_U5 (.ZN( us23_n503 ) , .A2( us23_n678 ) , .A3( us23_n776 ) , .A1( us23_n875 ) );
  NAND4_X1 us23_U50 (.ZN( sa21_sr_0 ) , .A4( us23_n500 ) , .A3( us23_n501 ) , .A2( us23_n502 ) , .A1( us23_n503 ) );
  NOR4_X1 us23_U51 (.A4( us23_n497 ) , .A3( us23_n498 ) , .A2( us23_n499 ) , .ZN( us23_n500 ) , .A1( us23_n526 ) );
  AOI221_X1 us23_U52 (.A( us23_n496 ) , .ZN( us23_n501 ) , .B2( us23_n842 ) , .C1( us23_n845 ) , .C2( us23_n859 ) , .B1( us23_n861 ) );
  AOI211_X1 us23_U53 (.A( us23_n495 ) , .ZN( us23_n502 ) , .B( us23_n801 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  AND3_X1 us23_U54 (.ZN( us23_n438 ) , .A2( us23_n642 ) , .A3( us23_n643 ) , .A1( us23_n645 ) );
  NAND4_X1 us23_U55 (.ZN( sa21_sr_1 ) , .A4( us23_n594 ) , .A3( us23_n595 ) , .A2( us23_n596 ) , .A1( us23_n597 ) );
  NOR4_X1 us23_U56 (.A4( us23_n590 ) , .A3( us23_n591 ) , .A2( us23_n592 ) , .A1( us23_n593 ) , .ZN( us23_n594 ) );
  AOI211_X1 us23_U57 (.B( us23_n588 ) , .A( us23_n589 ) , .ZN( us23_n595 ) , .C2( us23_n810 ) , .C1( us23_n832 ) );
  AOI211_X1 us23_U58 (.A( us23_n587 ) , .ZN( us23_n596 ) , .B( us23_n620 ) , .C1( us23_n844 ) , .C2( us23_n854 ) );
  NOR2_X1 us23_U59 (.ZN( us23_n624 ) , .A2( us23_n835 ) , .A1( us23_n838 ) );
  INV_X1 us23_U6 (.A( us23_n705 ) , .ZN( us23_n875 ) );
  NOR4_X1 us23_U60 (.A4( us23_n628 ) , .A3( us23_n629 ) , .A2( us23_n630 ) , .A1( us23_n631 ) , .ZN( us23_n632 ) );
  AOI211_X1 us23_U61 (.B( us23_n622 ) , .A( us23_n623 ) , .ZN( us23_n634 ) , .C2( us23_n835 ) , .C1( us23_n862 ) );
  NOR4_X1 us23_U62 (.A4( us23_n625 ) , .A3( us23_n626 ) , .A2( us23_n627 ) , .ZN( us23_n633 ) , .A1( us23_n663 ) );
  NAND4_X1 us23_U63 (.A4( us23_n656 ) , .A3( us23_n657 ) , .A2( us23_n658 ) , .A1( us23_n659 ) , .ZN( us23_n799 ) );
  NOR3_X1 us23_U64 (.A3( us23_n650 ) , .A2( us23_n651 ) , .A1( us23_n652 ) , .ZN( us23_n657 ) );
  NOR3_X1 us23_U65 (.A3( us23_n647 ) , .A2( us23_n648 ) , .A1( us23_n649 ) , .ZN( us23_n658 ) );
  NOR3_X1 us23_U66 (.A3( us23_n653 ) , .A2( us23_n654 ) , .A1( us23_n655 ) , .ZN( us23_n656 ) );
  NAND4_X1 us23_U67 (.A4( us23_n771 ) , .A3( us23_n772 ) , .A2( us23_n773 ) , .A1( us23_n774 ) , .ZN( us23_n800 ) );
  NOR3_X1 us23_U68 (.A3( us23_n764 ) , .A2( us23_n765 ) , .A1( us23_n766 ) , .ZN( us23_n772 ) );
  NOR4_X1 us23_U69 (.A4( us23_n767 ) , .A3( us23_n768 ) , .A2( us23_n769 ) , .A1( us23_n770 ) , .ZN( us23_n771 ) );
  NOR3_X1 us23_U7 (.A3( us23_n620 ) , .A2( us23_n621 ) , .ZN( us23_n635 ) , .A1( us23_n724 ) );
  AOI222_X1 us23_U70 (.ZN( us23_n774 ) , .A1( us23_n829 ) , .C1( us23_n833 ) , .B2( us23_n840 ) , .A2( us23_n849 ) , .B1( us23_n860 ) , .C2( us23_n872 ) );
  NOR4_X1 us23_U71 (.A4( us23_n576 ) , .A3( us23_n577 ) , .A2( us23_n578 ) , .ZN( us23_n585 ) , .A1( us23_n682 ) );
  NOR4_X1 us23_U72 (.A1( us23_n583 ) , .ZN( us23_n584 ) , .A3( us23_n651 ) , .A2( us23_n661 ) , .A4( us23_n766 ) );
  AOI221_X1 us23_U73 (.A( us23_n575 ) , .ZN( us23_n586 ) , .B2( us23_n830 ) , .C2( us23_n842 ) , .B1( us23_n853 ) , .C1( us23_n860 ) );
  NOR2_X1 us23_U74 (.ZN( us23_n760 ) , .A1( us23_n832 ) , .A2( us23_n833 ) );
  NAND4_X1 us23_U75 (.A4( us23_n455 ) , .A3( us23_n456 ) , .A2( us23_n457 ) , .A1( us23_n458 ) , .ZN( us23_n678 ) );
  NOR3_X1 us23_U76 (.ZN( us23_n456 ) , .A3( us23_n529 ) , .A1( us23_n554 ) , .A2( us23_n569 ) );
  NOR4_X1 us23_U77 (.ZN( us23_n457 ) , .A2( us23_n508 ) , .A1( us23_n598 ) , .A4( us23_n627 ) , .A3( us23_n710 ) );
  NOR4_X1 us23_U78 (.ZN( us23_n455 ) , .A2( us23_n516 ) , .A1( us23_n542 ) , .A3( us23_n578 ) , .A4( us23_n614 ) );
  NAND4_X1 us23_U79 (.A4( us23_n602 ) , .A3( us23_n603 ) , .A2( us23_n604 ) , .A1( us23_n605 ) , .ZN( us23_n721 ) );
  NOR2_X1 us23_U8 (.ZN( us23_n574 ) , .A1( us23_n621 ) , .A2( us23_n744 ) );
  NOR3_X1 us23_U80 (.A1( us23_n598 ) , .ZN( us23_n603 ) , .A3( us23_n662 ) , .A2( us23_n769 ) );
  NOR4_X1 us23_U81 (.A3( us23_n599 ) , .A2( us23_n600 ) , .A1( us23_n601 ) , .ZN( us23_n602 ) , .A4( us23_n654 ) );
  AOI222_X1 us23_U82 (.ZN( us23_n605 ) , .A1( us23_n829 ) , .C2( us23_n836 ) , .B1( us23_n841 ) , .A2( us23_n855 ) , .B2( us23_n860 ) , .C1( us23_n867 ) );
  NAND4_X1 us23_U83 (.A4( us23_n534 ) , .A3( us23_n535 ) , .A2( us23_n536 ) , .A1( us23_n537 ) , .ZN( us23_n621 ) );
  NOR4_X1 us23_U84 (.A4( us23_n525 ) , .A2( us23_n526 ) , .A1( us23_n527 ) , .ZN( us23_n537 ) , .A3( us23_n700 ) );
  NOR4_X1 us23_U85 (.A1( us23_n530 ) , .ZN( us23_n535 ) , .A2( us23_n653 ) , .A4( us23_n667 ) , .A3( us23_n764 ) );
  NOR4_X1 us23_U86 (.A4( us23_n528 ) , .A3( us23_n529 ) , .ZN( us23_n536 ) , .A2( us23_n683 ) , .A1( us23_n793 ) );
  NOR2_X1 us23_U87 (.ZN( us23_n685 ) , .A1( us23_n830 ) , .A2( us23_n831 ) );
  NAND4_X1 us23_U88 (.A4( us23_n547 ) , .A3( us23_n548 ) , .A2( us23_n549 ) , .A1( us23_n550 ) , .ZN( us23_n744 ) );
  NOR3_X1 us23_U89 (.ZN( us23_n548 ) , .A2( us23_n650 ) , .A1( us23_n666 ) , .A3( us23_n770 ) );
  NOR2_X1 us23_U9 (.A1( us23_n677 ) , .ZN( us23_n692 ) , .A2( us23_n806 ) );
  AOI211_X1 us23_U90 (.B( us23_n538 ) , .A( us23_n539 ) , .ZN( us23_n550 ) , .C2( us23_n838 ) , .C1( us23_n850 ) );
  NOR4_X1 us23_U91 (.A4( us23_n543 ) , .A3( us23_n544 ) , .A2( us23_n545 ) , .A1( us23_n546 ) , .ZN( us23_n547 ) );
  NAND4_X1 us23_U92 (.A4( us23_n478 ) , .A3( us23_n479 ) , .A2( us23_n480 ) , .A1( us23_n481 ) , .ZN( us23_n693 ) );
  NOR3_X1 us23_U93 (.ZN( us23_n479 ) , .A2( us23_n507 ) , .A3( us23_n600 ) , .A1( us23_n609 ) );
  AOI211_X1 us23_U94 (.B( us23_n476 ) , .A( us23_n477 ) , .ZN( us23_n481 ) , .C2( us23_n832 ) , .C1( us23_n860 ) );
  NOR4_X1 us23_U95 (.ZN( us23_n480 ) , .A3( us23_n531 ) , .A4( us23_n544 ) , .A2( us23_n566 ) , .A1( us23_n716 ) );
  NOR4_X1 us23_U96 (.ZN( us23_n619 ) , .A1( us23_n655 ) , .A3( us23_n665 ) , .A4( us23_n681 ) , .A2( us23_n765 ) );
  NOR4_X1 us23_U97 (.A4( us23_n608 ) , .A3( us23_n609 ) , .A2( us23_n610 ) , .A1( us23_n611 ) , .ZN( us23_n618 ) );
  NOR4_X1 us23_U98 (.A4( us23_n613 ) , .A3( us23_n614 ) , .A2( us23_n615 ) , .A1( us23_n616 ) , .ZN( us23_n617 ) );
  NAND4_X1 us23_U99 (.A4( us23_n484 ) , .A3( us23_n485 ) , .A2( us23_n486 ) , .A1( us23_n487 ) , .ZN( us23_n777 ) );
endmodule

