module des_des_die_14 ( u0_L12_11, u0_L12_19, u0_L12_29, u0_L12_4, u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, 
       u0_R12_25, u0_uk_K_r12_1, u0_uk_K_r12_30, u0_uk_K_r12_36, u0_uk_K_r12_7, u0_uk_n117, u0_uk_n141, u0_uk_n164, u0_uk_n220, 
       u0_uk_n230, u0_uk_n240, u0_uk_n251, u0_uk_n50, u0_uk_n51, u0_uk_n55, u0_uk_n61, u0_uk_n73, u0_uk_n88, 
       u0_uk_n89, u0_uk_n93, u0_uk_n94, u1_L0_11, u1_L0_19, u1_L0_29, u1_L0_4, u1_L10_1, u1_L10_10, 
       u1_L10_16, u1_L10_20, u1_L10_24, u1_L10_26, u1_L10_30, u1_L10_6, u1_L1_11, u1_L1_14, u1_L1_19, 
       u1_L1_25, u1_L1_29, u1_L1_3, u1_L1_4, u1_L1_8, u1_L3_12, u1_L3_22, u1_L3_32, u1_L3_7, 
       u1_L4_13, u1_L4_15, u1_L4_18, u1_L4_2, u1_L4_21, u1_L4_27, u1_L4_28, u1_L4_5, u1_R0_20, 
       u1_R0_21, u1_R0_22, u1_R0_23, u1_R0_24, u1_R0_25, u1_R10_10, u1_R10_11, u1_R10_12, u1_R10_13, 
       u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_8, u1_R10_9, u1_R1_16, u1_R1_17, u1_R1_18, 
       u1_R1_19, u1_R1_20, u1_R1_21, u1_R1_22, u1_R1_23, u1_R1_24, u1_R1_25, u1_R3_24, u1_R3_25, 
       u1_R3_26, u1_R3_27, u1_R3_28, u1_R3_29, u1_R4_1, u1_R4_28, u1_R4_29, u1_R4_30, u1_R4_31, 
       u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, u1_R4_7, u1_R4_8, u1_R4_9, u1_uk_K_r0_15, u1_uk_K_r0_31, 
       u1_uk_K_r0_36, u1_uk_K_r10_18, u1_uk_K_r10_25, u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_41, u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r1_36, 
       u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_7, u1_uk_K_r3_16, u1_uk_K_r3_9, u1_uk_K_r4_18, u1_uk_K_r4_23, u1_uk_K_r4_3, u1_uk_K_r4_33, 
       u1_uk_K_r4_41, u1_uk_K_r4_54, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n110, u1_uk_n118, 
       u1_uk_n1260, u1_uk_n1272, u1_uk_n1275, u1_uk_n1288, u1_uk_n129, u1_uk_n1293, u1_uk_n1303, u1_uk_n1308, u1_uk_n1309, 
       u1_uk_n1313, u1_uk_n1318, u1_uk_n1322, u1_uk_n1328, u1_uk_n1329, u1_uk_n1333, u1_uk_n1339, u1_uk_n1343, u1_uk_n1344, 
       u1_uk_n1345, u1_uk_n1394, u1_uk_n1395, u1_uk_n1406, u1_uk_n141, u1_uk_n1412, u1_uk_n1413, u1_uk_n1418, u1_uk_n142, 
       u1_uk_n1426, u1_uk_n1430, u1_uk_n1433, u1_uk_n1438, u1_uk_n1440, u1_uk_n1443, u1_uk_n1446, u1_uk_n1449, u1_uk_n145, 
       u1_uk_n1453, u1_uk_n1454, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n146, u1_uk_n1463, u1_uk_n1465, 
       u1_uk_n147, u1_uk_n1470, u1_uk_n1471, u1_uk_n1476, u1_uk_n1477, u1_uk_n161, u1_uk_n162, u1_uk_n163, u1_uk_n164, 
       u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, u1_uk_n1716, u1_uk_n1718, u1_uk_n1719, u1_uk_n1722, u1_uk_n1723, u1_uk_n1732, 
       u1_uk_n1745, u1_uk_n1750, u1_uk_n1751, u1_uk_n182, u1_uk_n188, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, 
       u1_uk_n208, u1_uk_n209, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n231, u1_uk_n238, u1_uk_n240, 
       u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n286, 
       u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n93, u1_uk_n94, u1_uk_n99, u2_K12_20, u2_K12_22, 
       u2_K12_24, u2_K9_45, u2_L10_1, u2_L10_10, u2_L10_16, u2_L10_20, u2_L10_24, u2_L10_26, u2_L10_30, 
       u2_L10_6, u2_L7_15, u2_L7_21, u2_L7_27, u2_L7_5, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, 
       u2_R10_14, u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_8, u2_R10_9, u2_R7_1, u2_R7_28, u2_R7_29, 
       u2_R7_30, u2_R7_31, u2_R7_32, u2_uk_K_r10_25, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_41, u2_uk_K_r1_7, u2_uk_K_r7_0, 
       u2_uk_K_r7_37, u2_uk_n10, u2_uk_n102, u2_uk_n109, u2_uk_n1140, u2_uk_n117, u2_uk_n128, u2_uk_n155, u2_uk_n1558, 
       u2_uk_n1565, u2_uk_n1576, u2_uk_n1577, u2_uk_n1583, u2_uk_n1585, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, 
       u2_uk_n1689, u2_uk_n1693, u2_uk_n1720, u2_uk_n1721, u2_uk_n203, u2_uk_n209, u2_uk_n214, u2_uk_n220, u2_uk_n222, 
       u2_uk_n231, u2_uk_n415, u2_uk_n443, u2_uk_n92, u0_N419, u0_N426, u0_N434, u0_N444, u1_N134, u1_N139, u1_N149, u1_N159, u1_N161, 
        u1_N164, u1_N172, u1_N174, u1_N177, u1_N180, u1_N186, u1_N187, u1_N35, u1_N352, 
        u1_N357, u1_N361, u1_N367, u1_N371, u1_N375, u1_N377, u1_N381, u1_N42, u1_N50, 
        u1_N60, u1_N66, u1_N67, u1_N71, u1_N74, u1_N77, u1_N82, u1_N88, u1_N92, 
        u2_N260, u2_N270, u2_N276, u2_N282, u2_N352, u2_N357, u2_N361, u2_N367, u2_N371, 
        u2_N375, u2_N377, u2_N381, u2_uk_n1012 );
  input u0_L12_11, u0_L12_19, u0_L12_29, u0_L12_4, u0_R12_20, u0_R12_21, u0_R12_22, u0_R12_23, u0_R12_24, 
        u0_R12_25, u0_uk_K_r12_1, u0_uk_K_r12_30, u0_uk_K_r12_36, u0_uk_K_r12_7, u0_uk_n117, u0_uk_n141, u0_uk_n164, u0_uk_n220, 
        u0_uk_n230, u0_uk_n240, u0_uk_n251, u0_uk_n50, u0_uk_n51, u0_uk_n55, u0_uk_n61, u0_uk_n73, u0_uk_n88, 
        u0_uk_n89, u0_uk_n93, u0_uk_n94, u1_L0_11, u1_L0_19, u1_L0_29, u1_L0_4, u1_L10_1, u1_L10_10, 
        u1_L10_16, u1_L10_20, u1_L10_24, u1_L10_26, u1_L10_30, u1_L10_6, u1_L1_11, u1_L1_14, u1_L1_19, 
        u1_L1_25, u1_L1_29, u1_L1_3, u1_L1_4, u1_L1_8, u1_L3_12, u1_L3_22, u1_L3_32, u1_L3_7, 
        u1_L4_13, u1_L4_15, u1_L4_18, u1_L4_2, u1_L4_21, u1_L4_27, u1_L4_28, u1_L4_5, u1_R0_20, 
        u1_R0_21, u1_R0_22, u1_R0_23, u1_R0_24, u1_R0_25, u1_R10_10, u1_R10_11, u1_R10_12, u1_R10_13, 
        u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_8, u1_R10_9, u1_R1_16, u1_R1_17, u1_R1_18, 
        u1_R1_19, u1_R1_20, u1_R1_21, u1_R1_22, u1_R1_23, u1_R1_24, u1_R1_25, u1_R3_24, u1_R3_25, 
        u1_R3_26, u1_R3_27, u1_R3_28, u1_R3_29, u1_R4_1, u1_R4_28, u1_R4_29, u1_R4_30, u1_R4_31, 
        u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_6, u1_R4_7, u1_R4_8, u1_R4_9, u1_uk_K_r0_15, u1_uk_K_r0_31, 
        u1_uk_K_r0_36, u1_uk_K_r10_18, u1_uk_K_r10_25, u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_41, u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r1_36, 
        u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_7, u1_uk_K_r3_16, u1_uk_K_r3_9, u1_uk_K_r4_18, u1_uk_K_r4_23, u1_uk_K_r4_3, u1_uk_K_r4_33, 
        u1_uk_K_r4_41, u1_uk_K_r4_54, u1_uk_n10, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n11, u1_uk_n110, u1_uk_n118, 
        u1_uk_n1260, u1_uk_n1272, u1_uk_n1275, u1_uk_n1288, u1_uk_n129, u1_uk_n1293, u1_uk_n1303, u1_uk_n1308, u1_uk_n1309, 
        u1_uk_n1313, u1_uk_n1318, u1_uk_n1322, u1_uk_n1328, u1_uk_n1329, u1_uk_n1333, u1_uk_n1339, u1_uk_n1343, u1_uk_n1344, 
        u1_uk_n1345, u1_uk_n1394, u1_uk_n1395, u1_uk_n1406, u1_uk_n141, u1_uk_n1412, u1_uk_n1413, u1_uk_n1418, u1_uk_n142, 
        u1_uk_n1426, u1_uk_n1430, u1_uk_n1433, u1_uk_n1438, u1_uk_n1440, u1_uk_n1443, u1_uk_n1446, u1_uk_n1449, u1_uk_n145, 
        u1_uk_n1453, u1_uk_n1454, u1_uk_n1456, u1_uk_n1457, u1_uk_n1458, u1_uk_n1459, u1_uk_n146, u1_uk_n1463, u1_uk_n1465, 
        u1_uk_n147, u1_uk_n1470, u1_uk_n1471, u1_uk_n1476, u1_uk_n1477, u1_uk_n161, u1_uk_n162, u1_uk_n163, u1_uk_n164, 
        u1_uk_n1711, u1_uk_n1712, u1_uk_n1713, u1_uk_n1716, u1_uk_n1718, u1_uk_n1719, u1_uk_n1722, u1_uk_n1723, u1_uk_n1732, 
        u1_uk_n1745, u1_uk_n1750, u1_uk_n1751, u1_uk_n182, u1_uk_n188, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, 
        u1_uk_n208, u1_uk_n209, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n231, u1_uk_n238, u1_uk_n240, 
        u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n286, 
        u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n31, u1_uk_n93, u1_uk_n94, u1_uk_n99, u2_K12_20, u2_K12_22, 
        u2_K12_24, u2_K9_45, u2_L10_1, u2_L10_10, u2_L10_16, u2_L10_20, u2_L10_24, u2_L10_26, u2_L10_30, 
        u2_L10_6, u2_L7_15, u2_L7_21, u2_L7_27, u2_L7_5, u2_R10_10, u2_R10_11, u2_R10_12, u2_R10_13, 
        u2_R10_14, u2_R10_15, u2_R10_16, u2_R10_17, u2_R10_8, u2_R10_9, u2_R7_1, u2_R7_28, u2_R7_29, 
        u2_R7_30, u2_R7_31, u2_R7_32, u2_uk_K_r10_25, u2_uk_K_r10_32, u2_uk_K_r10_34, u2_uk_K_r10_41, u2_uk_K_r1_7, u2_uk_K_r7_0, 
        u2_uk_K_r7_37, u2_uk_n10, u2_uk_n102, u2_uk_n109, u2_uk_n1140, u2_uk_n117, u2_uk_n128, u2_uk_n155, u2_uk_n1558, 
        u2_uk_n1565, u2_uk_n1576, u2_uk_n1577, u2_uk_n1583, u2_uk_n1585, u2_uk_n1681, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, 
        u2_uk_n1689, u2_uk_n1693, u2_uk_n1720, u2_uk_n1721, u2_uk_n203, u2_uk_n209, u2_uk_n214, u2_uk_n220, u2_uk_n222, 
        u2_uk_n231, u2_uk_n415, u2_uk_n443, u2_uk_n92;
  output u0_N419, u0_N426, u0_N434, u0_N444, u1_N134, u1_N139, u1_N149, u1_N159, u1_N161, 
        u1_N164, u1_N172, u1_N174, u1_N177, u1_N180, u1_N186, u1_N187, u1_N35, u1_N352, 
        u1_N357, u1_N361, u1_N367, u1_N371, u1_N375, u1_N377, u1_N381, u1_N42, u1_N50, 
        u1_N60, u1_N66, u1_N67, u1_N71, u1_N74, u1_N77, u1_N82, u1_N88, u1_N92, 
        u2_N260, u2_N270, u2_N276, u2_N282, u2_N352, u2_N357, u2_N361, u2_N367, u2_N371, 
        u2_N375, u2_N377, u2_N381, u2_uk_n1012;
  wire u0_K14_31, u0_K14_32, u0_K14_33, u0_K14_34, u0_K14_35, u0_K14_36, u0_out13_11, u0_out13_19, u0_out13_29, 
       u0_out13_4, u0_u13_X_31, u0_u13_X_32, u0_u13_X_33, u0_u13_X_34, u0_u13_X_35, u0_u13_X_36, u0_u13_u5_n100, u0_u13_u5_n101, 
       u0_u13_u5_n102, u0_u13_u5_n103, u0_u13_u5_n104, u0_u13_u5_n105, u0_u13_u5_n106, u0_u13_u5_n107, u0_u13_u5_n108, u0_u13_u5_n109, u0_u13_u5_n110, 
       u0_u13_u5_n111, u0_u13_u5_n112, u0_u13_u5_n113, u0_u13_u5_n114, u0_u13_u5_n115, u0_u13_u5_n116, u0_u13_u5_n117, u0_u13_u5_n118, u0_u13_u5_n119, 
       u0_u13_u5_n120, u0_u13_u5_n121, u0_u13_u5_n122, u0_u13_u5_n123, u0_u13_u5_n124, u0_u13_u5_n125, u0_u13_u5_n126, u0_u13_u5_n127, u0_u13_u5_n128, 
       u0_u13_u5_n129, u0_u13_u5_n130, u0_u13_u5_n131, u0_u13_u5_n132, u0_u13_u5_n133, u0_u13_u5_n134, u0_u13_u5_n135, u0_u13_u5_n136, u0_u13_u5_n137, 
       u0_u13_u5_n138, u0_u13_u5_n139, u0_u13_u5_n140, u0_u13_u5_n141, u0_u13_u5_n142, u0_u13_u5_n143, u0_u13_u5_n144, u0_u13_u5_n145, u0_u13_u5_n146, 
       u0_u13_u5_n147, u0_u13_u5_n148, u0_u13_u5_n149, u0_u13_u5_n150, u0_u13_u5_n151, u0_u13_u5_n152, u0_u13_u5_n153, u0_u13_u5_n154, u0_u13_u5_n155, 
       u0_u13_u5_n156, u0_u13_u5_n157, u0_u13_u5_n158, u0_u13_u5_n159, u0_u13_u5_n160, u0_u13_u5_n161, u0_u13_u5_n162, u0_u13_u5_n163, u0_u13_u5_n164, 
       u0_u13_u5_n165, u0_u13_u5_n166, u0_u13_u5_n167, u0_u13_u5_n168, u0_u13_u5_n169, u0_u13_u5_n170, u0_u13_u5_n171, u0_u13_u5_n172, u0_u13_u5_n173, 
       u0_u13_u5_n174, u0_u13_u5_n175, u0_u13_u5_n176, u0_u13_u5_n177, u0_u13_u5_n178, u0_u13_u5_n179, u0_u13_u5_n180, u0_u13_u5_n181, u0_u13_u5_n182, 
       u0_u13_u5_n183, u0_u13_u5_n184, u0_u13_u5_n185, u0_u13_u5_n186, u0_u13_u5_n187, u0_u13_u5_n188, u0_u13_u5_n189, u0_u13_u5_n190, u0_u13_u5_n191, 
       u0_u13_u5_n192, u0_u13_u5_n193, u0_u13_u5_n194, u0_u13_u5_n195, u0_u13_u5_n196, u0_u13_u5_n99, u0_uk_n933, u0_uk_n934, u1_K12_13, 
       u1_K12_14, u1_K12_15, u1_K12_16, u1_K12_17, u1_K12_18, u1_K12_19, u1_K12_20, u1_K12_21, u1_K12_22, 
       u1_K12_23, u1_K12_24, u1_K2_31, u1_K2_32, u1_K2_33, u1_K2_34, u1_K2_35, u1_K2_36, u1_K3_25, 
       u1_K3_26, u1_K3_27, u1_K3_28, u1_K3_29, u1_K3_30, u1_K3_31, u1_K3_32, u1_K3_33, u1_K3_34, 
       u1_K3_35, u1_K3_36, u1_K5_37, u1_K5_38, u1_K5_39, u1_K5_40, u1_K5_41, u1_K5_42, u1_K6_10, 
       u1_K6_11, u1_K6_12, u1_K6_43, u1_K6_44, u1_K6_45, u1_K6_46, u1_K6_47, u1_K6_48, u1_K6_7, 
       u1_K6_8, u1_K6_9, u1_out11_1, u1_out11_10, u1_out11_16, u1_out11_20, u1_out11_24, u1_out11_26, u1_out11_30, 
       u1_out11_6, u1_out1_11, u1_out1_19, u1_out1_29, u1_out1_4, u1_out2_11, u1_out2_14, u1_out2_19, u1_out2_25, 
       u1_out2_29, u1_out2_3, u1_out2_4, u1_out2_8, u1_out4_12, u1_out4_22, u1_out4_32, u1_out4_7, u1_out5_13, 
       u1_out5_15, u1_out5_18, u1_out5_2, u1_out5_21, u1_out5_27, u1_out5_28, u1_out5_5, u1_u11_X_13, u1_u11_X_14, 
       u1_u11_X_15, u1_u11_X_16, u1_u11_X_17, u1_u11_X_18, u1_u11_X_19, u1_u11_X_20, u1_u11_X_21, u1_u11_X_22, u1_u11_X_23, 
       u1_u11_X_24, u1_u11_u2_n100, u1_u11_u2_n101, u1_u11_u2_n102, u1_u11_u2_n103, u1_u11_u2_n104, u1_u11_u2_n105, u1_u11_u2_n106, u1_u11_u2_n107, 
       u1_u11_u2_n108, u1_u11_u2_n109, u1_u11_u2_n110, u1_u11_u2_n111, u1_u11_u2_n112, u1_u11_u2_n113, u1_u11_u2_n114, u1_u11_u2_n115, u1_u11_u2_n116, 
       u1_u11_u2_n117, u1_u11_u2_n118, u1_u11_u2_n119, u1_u11_u2_n120, u1_u11_u2_n121, u1_u11_u2_n122, u1_u11_u2_n123, u1_u11_u2_n124, u1_u11_u2_n125, 
       u1_u11_u2_n126, u1_u11_u2_n127, u1_u11_u2_n128, u1_u11_u2_n129, u1_u11_u2_n130, u1_u11_u2_n131, u1_u11_u2_n132, u1_u11_u2_n133, u1_u11_u2_n134, 
       u1_u11_u2_n135, u1_u11_u2_n136, u1_u11_u2_n137, u1_u11_u2_n138, u1_u11_u2_n139, u1_u11_u2_n140, u1_u11_u2_n141, u1_u11_u2_n142, u1_u11_u2_n143, 
       u1_u11_u2_n144, u1_u11_u2_n145, u1_u11_u2_n146, u1_u11_u2_n147, u1_u11_u2_n148, u1_u11_u2_n149, u1_u11_u2_n150, u1_u11_u2_n151, u1_u11_u2_n152, 
       u1_u11_u2_n153, u1_u11_u2_n154, u1_u11_u2_n155, u1_u11_u2_n156, u1_u11_u2_n157, u1_u11_u2_n158, u1_u11_u2_n159, u1_u11_u2_n160, u1_u11_u2_n161, 
       u1_u11_u2_n162, u1_u11_u2_n163, u1_u11_u2_n164, u1_u11_u2_n165, u1_u11_u2_n166, u1_u11_u2_n167, u1_u11_u2_n168, u1_u11_u2_n169, u1_u11_u2_n170, 
       u1_u11_u2_n171, u1_u11_u2_n172, u1_u11_u2_n173, u1_u11_u2_n174, u1_u11_u2_n175, u1_u11_u2_n176, u1_u11_u2_n177, u1_u11_u2_n178, u1_u11_u2_n179, 
       u1_u11_u2_n180, u1_u11_u2_n181, u1_u11_u2_n182, u1_u11_u2_n183, u1_u11_u2_n184, u1_u11_u2_n185, u1_u11_u2_n186, u1_u11_u2_n187, u1_u11_u2_n188, 
       u1_u11_u2_n95, u1_u11_u2_n96, u1_u11_u2_n97, u1_u11_u2_n98, u1_u11_u2_n99, u1_u11_u3_n100, u1_u11_u3_n101, u1_u11_u3_n102, u1_u11_u3_n103, 
       u1_u11_u3_n104, u1_u11_u3_n105, u1_u11_u3_n106, u1_u11_u3_n107, u1_u11_u3_n108, u1_u11_u3_n109, u1_u11_u3_n110, u1_u11_u3_n111, u1_u11_u3_n112, 
       u1_u11_u3_n113, u1_u11_u3_n114, u1_u11_u3_n115, u1_u11_u3_n116, u1_u11_u3_n117, u1_u11_u3_n118, u1_u11_u3_n119, u1_u11_u3_n120, u1_u11_u3_n121, 
       u1_u11_u3_n122, u1_u11_u3_n123, u1_u11_u3_n124, u1_u11_u3_n125, u1_u11_u3_n126, u1_u11_u3_n127, u1_u11_u3_n128, u1_u11_u3_n129, u1_u11_u3_n130, 
       u1_u11_u3_n131, u1_u11_u3_n132, u1_u11_u3_n133, u1_u11_u3_n134, u1_u11_u3_n135, u1_u11_u3_n136, u1_u11_u3_n137, u1_u11_u3_n138, u1_u11_u3_n139, 
       u1_u11_u3_n140, u1_u11_u3_n141, u1_u11_u3_n142, u1_u11_u3_n143, u1_u11_u3_n144, u1_u11_u3_n145, u1_u11_u3_n146, u1_u11_u3_n147, u1_u11_u3_n148, 
       u1_u11_u3_n149, u1_u11_u3_n150, u1_u11_u3_n151, u1_u11_u3_n152, u1_u11_u3_n153, u1_u11_u3_n154, u1_u11_u3_n155, u1_u11_u3_n156, u1_u11_u3_n157, 
       u1_u11_u3_n158, u1_u11_u3_n159, u1_u11_u3_n160, u1_u11_u3_n161, u1_u11_u3_n162, u1_u11_u3_n163, u1_u11_u3_n164, u1_u11_u3_n165, u1_u11_u3_n166, 
       u1_u11_u3_n167, u1_u11_u3_n168, u1_u11_u3_n169, u1_u11_u3_n170, u1_u11_u3_n171, u1_u11_u3_n172, u1_u11_u3_n173, u1_u11_u3_n174, u1_u11_u3_n175, 
       u1_u11_u3_n176, u1_u11_u3_n177, u1_u11_u3_n178, u1_u11_u3_n179, u1_u11_u3_n180, u1_u11_u3_n181, u1_u11_u3_n182, u1_u11_u3_n183, u1_u11_u3_n184, 
       u1_u11_u3_n185, u1_u11_u3_n186, u1_u11_u3_n94, u1_u11_u3_n95, u1_u11_u3_n96, u1_u11_u3_n97, u1_u11_u3_n98, u1_u11_u3_n99, u1_u1_X_31, 
       u1_u1_X_32, u1_u1_X_33, u1_u1_X_34, u1_u1_X_35, u1_u1_X_36, u1_u1_u5_n100, u1_u1_u5_n101, u1_u1_u5_n102, u1_u1_u5_n103, 
       u1_u1_u5_n104, u1_u1_u5_n105, u1_u1_u5_n106, u1_u1_u5_n107, u1_u1_u5_n108, u1_u1_u5_n109, u1_u1_u5_n110, u1_u1_u5_n111, u1_u1_u5_n112, 
       u1_u1_u5_n113, u1_u1_u5_n114, u1_u1_u5_n115, u1_u1_u5_n116, u1_u1_u5_n117, u1_u1_u5_n118, u1_u1_u5_n119, u1_u1_u5_n120, u1_u1_u5_n121, 
       u1_u1_u5_n122, u1_u1_u5_n123, u1_u1_u5_n124, u1_u1_u5_n125, u1_u1_u5_n126, u1_u1_u5_n127, u1_u1_u5_n128, u1_u1_u5_n129, u1_u1_u5_n130, 
       u1_u1_u5_n131, u1_u1_u5_n132, u1_u1_u5_n133, u1_u1_u5_n134, u1_u1_u5_n135, u1_u1_u5_n136, u1_u1_u5_n137, u1_u1_u5_n138, u1_u1_u5_n139, 
       u1_u1_u5_n140, u1_u1_u5_n141, u1_u1_u5_n142, u1_u1_u5_n143, u1_u1_u5_n144, u1_u1_u5_n145, u1_u1_u5_n146, u1_u1_u5_n147, u1_u1_u5_n148, 
       u1_u1_u5_n149, u1_u1_u5_n150, u1_u1_u5_n151, u1_u1_u5_n152, u1_u1_u5_n153, u1_u1_u5_n154, u1_u1_u5_n155, u1_u1_u5_n156, u1_u1_u5_n157, 
       u1_u1_u5_n158, u1_u1_u5_n159, u1_u1_u5_n160, u1_u1_u5_n161, u1_u1_u5_n162, u1_u1_u5_n163, u1_u1_u5_n164, u1_u1_u5_n165, u1_u1_u5_n166, 
       u1_u1_u5_n167, u1_u1_u5_n168, u1_u1_u5_n169, u1_u1_u5_n170, u1_u1_u5_n171, u1_u1_u5_n172, u1_u1_u5_n173, u1_u1_u5_n174, u1_u1_u5_n175, 
       u1_u1_u5_n176, u1_u1_u5_n177, u1_u1_u5_n178, u1_u1_u5_n179, u1_u1_u5_n180, u1_u1_u5_n181, u1_u1_u5_n182, u1_u1_u5_n183, u1_u1_u5_n184, 
       u1_u1_u5_n185, u1_u1_u5_n186, u1_u1_u5_n187, u1_u1_u5_n188, u1_u1_u5_n189, u1_u1_u5_n190, u1_u1_u5_n191, u1_u1_u5_n192, u1_u1_u5_n193, 
       u1_u1_u5_n194, u1_u1_u5_n195, u1_u1_u5_n196, u1_u1_u5_n99, u1_u2_X_25, u1_u2_X_26, u1_u2_X_27, u1_u2_X_28, u1_u2_X_29, 
       u1_u2_X_30, u1_u2_X_31, u1_u2_X_32, u1_u2_X_33, u1_u2_X_34, u1_u2_X_35, u1_u2_X_36, u1_u2_u4_n100, u1_u2_u4_n101, 
       u1_u2_u4_n102, u1_u2_u4_n103, u1_u2_u4_n104, u1_u2_u4_n105, u1_u2_u4_n106, u1_u2_u4_n107, u1_u2_u4_n108, u1_u2_u4_n109, u1_u2_u4_n110, 
       u1_u2_u4_n111, u1_u2_u4_n112, u1_u2_u4_n113, u1_u2_u4_n114, u1_u2_u4_n115, u1_u2_u4_n116, u1_u2_u4_n117, u1_u2_u4_n118, u1_u2_u4_n119, 
       u1_u2_u4_n120, u1_u2_u4_n121, u1_u2_u4_n122, u1_u2_u4_n123, u1_u2_u4_n124, u1_u2_u4_n125, u1_u2_u4_n126, u1_u2_u4_n127, u1_u2_u4_n128, 
       u1_u2_u4_n129, u1_u2_u4_n130, u1_u2_u4_n131, u1_u2_u4_n132, u1_u2_u4_n133, u1_u2_u4_n134, u1_u2_u4_n135, u1_u2_u4_n136, u1_u2_u4_n137, 
       u1_u2_u4_n138, u1_u2_u4_n139, u1_u2_u4_n140, u1_u2_u4_n141, u1_u2_u4_n142, u1_u2_u4_n143, u1_u2_u4_n144, u1_u2_u4_n145, u1_u2_u4_n146, 
       u1_u2_u4_n147, u1_u2_u4_n148, u1_u2_u4_n149, u1_u2_u4_n150, u1_u2_u4_n151, u1_u2_u4_n152, u1_u2_u4_n153, u1_u2_u4_n154, u1_u2_u4_n155, 
       u1_u2_u4_n156, u1_u2_u4_n157, u1_u2_u4_n158, u1_u2_u4_n159, u1_u2_u4_n160, u1_u2_u4_n161, u1_u2_u4_n162, u1_u2_u4_n163, u1_u2_u4_n164, 
       u1_u2_u4_n165, u1_u2_u4_n166, u1_u2_u4_n167, u1_u2_u4_n168, u1_u2_u4_n169, u1_u2_u4_n170, u1_u2_u4_n171, u1_u2_u4_n172, u1_u2_u4_n173, 
       u1_u2_u4_n174, u1_u2_u4_n175, u1_u2_u4_n176, u1_u2_u4_n177, u1_u2_u4_n178, u1_u2_u4_n179, u1_u2_u4_n180, u1_u2_u4_n181, u1_u2_u4_n182, 
       u1_u2_u4_n183, u1_u2_u4_n184, u1_u2_u4_n185, u1_u2_u4_n186, u1_u2_u4_n94, u1_u2_u4_n95, u1_u2_u4_n96, u1_u2_u4_n97, u1_u2_u4_n98, 
       u1_u2_u4_n99, u1_u2_u5_n100, u1_u2_u5_n101, u1_u2_u5_n102, u1_u2_u5_n103, u1_u2_u5_n104, u1_u2_u5_n105, u1_u2_u5_n106, u1_u2_u5_n107, 
       u1_u2_u5_n108, u1_u2_u5_n109, u1_u2_u5_n110, u1_u2_u5_n111, u1_u2_u5_n112, u1_u2_u5_n113, u1_u2_u5_n114, u1_u2_u5_n115, u1_u2_u5_n116, 
       u1_u2_u5_n117, u1_u2_u5_n118, u1_u2_u5_n119, u1_u2_u5_n120, u1_u2_u5_n121, u1_u2_u5_n122, u1_u2_u5_n123, u1_u2_u5_n124, u1_u2_u5_n125, 
       u1_u2_u5_n126, u1_u2_u5_n127, u1_u2_u5_n128, u1_u2_u5_n129, u1_u2_u5_n130, u1_u2_u5_n131, u1_u2_u5_n132, u1_u2_u5_n133, u1_u2_u5_n134, 
       u1_u2_u5_n135, u1_u2_u5_n136, u1_u2_u5_n137, u1_u2_u5_n138, u1_u2_u5_n139, u1_u2_u5_n140, u1_u2_u5_n141, u1_u2_u5_n142, u1_u2_u5_n143, 
       u1_u2_u5_n144, u1_u2_u5_n145, u1_u2_u5_n146, u1_u2_u5_n147, u1_u2_u5_n148, u1_u2_u5_n149, u1_u2_u5_n150, u1_u2_u5_n151, u1_u2_u5_n152, 
       u1_u2_u5_n153, u1_u2_u5_n154, u1_u2_u5_n155, u1_u2_u5_n156, u1_u2_u5_n157, u1_u2_u5_n158, u1_u2_u5_n159, u1_u2_u5_n160, u1_u2_u5_n161, 
       u1_u2_u5_n162, u1_u2_u5_n163, u1_u2_u5_n164, u1_u2_u5_n165, u1_u2_u5_n166, u1_u2_u5_n167, u1_u2_u5_n168, u1_u2_u5_n169, u1_u2_u5_n170, 
       u1_u2_u5_n171, u1_u2_u5_n172, u1_u2_u5_n173, u1_u2_u5_n174, u1_u2_u5_n175, u1_u2_u5_n176, u1_u2_u5_n177, u1_u2_u5_n178, u1_u2_u5_n179, 
       u1_u2_u5_n180, u1_u2_u5_n181, u1_u2_u5_n182, u1_u2_u5_n183, u1_u2_u5_n184, u1_u2_u5_n185, u1_u2_u5_n186, u1_u2_u5_n187, u1_u2_u5_n188, 
       u1_u2_u5_n189, u1_u2_u5_n190, u1_u2_u5_n191, u1_u2_u5_n192, u1_u2_u5_n193, u1_u2_u5_n194, u1_u2_u5_n195, u1_u2_u5_n196, u1_u2_u5_n99, 
       u1_u4_X_37, u1_u4_X_38, u1_u4_X_39, u1_u4_X_40, u1_u4_X_41, u1_u4_X_42, u1_u4_u6_n100, u1_u4_u6_n101, u1_u4_u6_n102, 
       u1_u4_u6_n103, u1_u4_u6_n104, u1_u4_u6_n105, u1_u4_u6_n106, u1_u4_u6_n107, u1_u4_u6_n108, u1_u4_u6_n109, u1_u4_u6_n110, u1_u4_u6_n111, 
       u1_u4_u6_n112, u1_u4_u6_n113, u1_u4_u6_n114, u1_u4_u6_n115, u1_u4_u6_n116, u1_u4_u6_n117, u1_u4_u6_n118, u1_u4_u6_n119, u1_u4_u6_n120, 
       u1_u4_u6_n121, u1_u4_u6_n122, u1_u4_u6_n123, u1_u4_u6_n124, u1_u4_u6_n125, u1_u4_u6_n126, u1_u4_u6_n127, u1_u4_u6_n128, u1_u4_u6_n129, 
       u1_u4_u6_n130, u1_u4_u6_n131, u1_u4_u6_n132, u1_u4_u6_n133, u1_u4_u6_n134, u1_u4_u6_n135, u1_u4_u6_n136, u1_u4_u6_n137, u1_u4_u6_n138, 
       u1_u4_u6_n139, u1_u4_u6_n140, u1_u4_u6_n141, u1_u4_u6_n142, u1_u4_u6_n143, u1_u4_u6_n144, u1_u4_u6_n145, u1_u4_u6_n146, u1_u4_u6_n147, 
       u1_u4_u6_n148, u1_u4_u6_n149, u1_u4_u6_n150, u1_u4_u6_n151, u1_u4_u6_n152, u1_u4_u6_n153, u1_u4_u6_n154, u1_u4_u6_n155, u1_u4_u6_n156, 
       u1_u4_u6_n157, u1_u4_u6_n158, u1_u4_u6_n159, u1_u4_u6_n160, u1_u4_u6_n161, u1_u4_u6_n162, u1_u4_u6_n163, u1_u4_u6_n164, u1_u4_u6_n165, 
       u1_u4_u6_n166, u1_u4_u6_n167, u1_u4_u6_n168, u1_u4_u6_n169, u1_u4_u6_n170, u1_u4_u6_n171, u1_u4_u6_n172, u1_u4_u6_n173, u1_u4_u6_n174, 
       u1_u4_u6_n88, u1_u4_u6_n89, u1_u4_u6_n90, u1_u4_u6_n91, u1_u4_u6_n92, u1_u4_u6_n93, u1_u4_u6_n94, u1_u4_u6_n95, u1_u4_u6_n96, 
       u1_u4_u6_n97, u1_u4_u6_n98, u1_u4_u6_n99, u1_u5_X_10, u1_u5_X_11, u1_u5_X_12, u1_u5_X_43, u1_u5_X_44, u1_u5_X_45, 
       u1_u5_X_46, u1_u5_X_47, u1_u5_X_48, u1_u5_X_7, u1_u5_X_8, u1_u5_X_9, u1_u5_u1_n100, u1_u5_u1_n101, u1_u5_u1_n102, 
       u1_u5_u1_n103, u1_u5_u1_n104, u1_u5_u1_n105, u1_u5_u1_n106, u1_u5_u1_n107, u1_u5_u1_n108, u1_u5_u1_n109, u1_u5_u1_n110, u1_u5_u1_n111, 
       u1_u5_u1_n112, u1_u5_u1_n113, u1_u5_u1_n114, u1_u5_u1_n115, u1_u5_u1_n116, u1_u5_u1_n117, u1_u5_u1_n118, u1_u5_u1_n119, u1_u5_u1_n120, 
       u1_u5_u1_n121, u1_u5_u1_n122, u1_u5_u1_n123, u1_u5_u1_n124, u1_u5_u1_n125, u1_u5_u1_n126, u1_u5_u1_n127, u1_u5_u1_n128, u1_u5_u1_n129, 
       u1_u5_u1_n130, u1_u5_u1_n131, u1_u5_u1_n132, u1_u5_u1_n133, u1_u5_u1_n134, u1_u5_u1_n135, u1_u5_u1_n136, u1_u5_u1_n137, u1_u5_u1_n138, 
       u1_u5_u1_n139, u1_u5_u1_n140, u1_u5_u1_n141, u1_u5_u1_n142, u1_u5_u1_n143, u1_u5_u1_n144, u1_u5_u1_n145, u1_u5_u1_n146, u1_u5_u1_n147, 
       u1_u5_u1_n148, u1_u5_u1_n149, u1_u5_u1_n150, u1_u5_u1_n151, u1_u5_u1_n152, u1_u5_u1_n153, u1_u5_u1_n154, u1_u5_u1_n155, u1_u5_u1_n156, 
       u1_u5_u1_n157, u1_u5_u1_n158, u1_u5_u1_n159, u1_u5_u1_n160, u1_u5_u1_n161, u1_u5_u1_n162, u1_u5_u1_n163, u1_u5_u1_n164, u1_u5_u1_n165, 
       u1_u5_u1_n166, u1_u5_u1_n167, u1_u5_u1_n168, u1_u5_u1_n169, u1_u5_u1_n170, u1_u5_u1_n171, u1_u5_u1_n172, u1_u5_u1_n173, u1_u5_u1_n174, 
       u1_u5_u1_n175, u1_u5_u1_n176, u1_u5_u1_n177, u1_u5_u1_n178, u1_u5_u1_n179, u1_u5_u1_n180, u1_u5_u1_n181, u1_u5_u1_n182, u1_u5_u1_n183, 
       u1_u5_u1_n184, u1_u5_u1_n185, u1_u5_u1_n186, u1_u5_u1_n187, u1_u5_u1_n188, u1_u5_u1_n95, u1_u5_u1_n96, u1_u5_u1_n97, u1_u5_u1_n98, 
       u1_u5_u1_n99, u1_u5_u7_n100, u1_u5_u7_n101, u1_u5_u7_n102, u1_u5_u7_n103, u1_u5_u7_n104, u1_u5_u7_n105, u1_u5_u7_n106, u1_u5_u7_n107, 
       u1_u5_u7_n108, u1_u5_u7_n109, u1_u5_u7_n110, u1_u5_u7_n111, u1_u5_u7_n112, u1_u5_u7_n113, u1_u5_u7_n114, u1_u5_u7_n115, u1_u5_u7_n116, 
       u1_u5_u7_n117, u1_u5_u7_n118, u1_u5_u7_n119, u1_u5_u7_n120, u1_u5_u7_n121, u1_u5_u7_n122, u1_u5_u7_n123, u1_u5_u7_n124, u1_u5_u7_n125, 
       u1_u5_u7_n126, u1_u5_u7_n127, u1_u5_u7_n128, u1_u5_u7_n129, u1_u5_u7_n130, u1_u5_u7_n131, u1_u5_u7_n132, u1_u5_u7_n133, u1_u5_u7_n134, 
       u1_u5_u7_n135, u1_u5_u7_n136, u1_u5_u7_n137, u1_u5_u7_n138, u1_u5_u7_n139, u1_u5_u7_n140, u1_u5_u7_n141, u1_u5_u7_n142, u1_u5_u7_n143, 
       u1_u5_u7_n144, u1_u5_u7_n145, u1_u5_u7_n146, u1_u5_u7_n147, u1_u5_u7_n148, u1_u5_u7_n149, u1_u5_u7_n150, u1_u5_u7_n151, u1_u5_u7_n152, 
       u1_u5_u7_n153, u1_u5_u7_n154, u1_u5_u7_n155, u1_u5_u7_n156, u1_u5_u7_n157, u1_u5_u7_n158, u1_u5_u7_n159, u1_u5_u7_n160, u1_u5_u7_n161, 
       u1_u5_u7_n162, u1_u5_u7_n163, u1_u5_u7_n164, u1_u5_u7_n165, u1_u5_u7_n166, u1_u5_u7_n167, u1_u5_u7_n168, u1_u5_u7_n169, u1_u5_u7_n170, 
       u1_u5_u7_n171, u1_u5_u7_n172, u1_u5_u7_n173, u1_u5_u7_n174, u1_u5_u7_n175, u1_u5_u7_n176, u1_u5_u7_n177, u1_u5_u7_n178, u1_u5_u7_n179, 
       u1_u5_u7_n180, u1_u5_u7_n91, u1_u5_u7_n92, u1_u5_u7_n93, u1_u5_u7_n94, u1_u5_u7_n95, u1_u5_u7_n96, u1_u5_u7_n97, u1_u5_u7_n98, 
       u1_u5_u7_n99, u1_uk_n1029, u1_uk_n1030, u1_uk_n1039, u1_uk_n1040, u1_uk_n1041, u1_uk_n1042, u1_uk_n1081, u1_uk_n1082, 
       u1_uk_n1088, u1_uk_n1100, u1_uk_n1102, u1_uk_n1103, u1_uk_n1104, u1_uk_n504, u1_uk_n509, u1_uk_n518, u1_uk_n520, 
       u1_uk_n524, u2_K12_13, u2_K12_14, u2_K12_15, u2_K12_16, u2_K12_17, u2_K12_18, u2_K12_19, u2_K12_21, 
       u2_K12_23, u2_K9_43, u2_K9_44, u2_K9_46, u2_K9_47, u2_K9_48, u2_out11_1, u2_out11_10, u2_out11_16, 
       u2_out11_20, u2_out11_24, u2_out11_26, u2_out11_30, u2_out11_6, u2_out8_15, u2_out8_21, u2_out8_27, u2_out8_5, 
       u2_u11_X_13, u2_u11_X_14, u2_u11_X_15, u2_u11_X_16, u2_u11_X_17, u2_u11_X_18, u2_u11_X_19, u2_u11_X_20, u2_u11_X_21, 
       u2_u11_X_22, u2_u11_X_23, u2_u11_X_24, u2_u11_u2_n100, u2_u11_u2_n101, u2_u11_u2_n102, u2_u11_u2_n103, u2_u11_u2_n104, u2_u11_u2_n105, 
       u2_u11_u2_n106, u2_u11_u2_n107, u2_u11_u2_n108, u2_u11_u2_n109, u2_u11_u2_n110, u2_u11_u2_n111, u2_u11_u2_n112, u2_u11_u2_n113, u2_u11_u2_n114, 
       u2_u11_u2_n115, u2_u11_u2_n116, u2_u11_u2_n117, u2_u11_u2_n118, u2_u11_u2_n119, u2_u11_u2_n120, u2_u11_u2_n121, u2_u11_u2_n122, u2_u11_u2_n123, 
       u2_u11_u2_n124, u2_u11_u2_n125, u2_u11_u2_n126, u2_u11_u2_n127, u2_u11_u2_n128, u2_u11_u2_n129, u2_u11_u2_n130, u2_u11_u2_n131, u2_u11_u2_n132, 
       u2_u11_u2_n133, u2_u11_u2_n134, u2_u11_u2_n135, u2_u11_u2_n136, u2_u11_u2_n137, u2_u11_u2_n138, u2_u11_u2_n139, u2_u11_u2_n140, u2_u11_u2_n141, 
       u2_u11_u2_n142, u2_u11_u2_n143, u2_u11_u2_n144, u2_u11_u2_n145, u2_u11_u2_n146, u2_u11_u2_n147, u2_u11_u2_n148, u2_u11_u2_n149, u2_u11_u2_n150, 
       u2_u11_u2_n151, u2_u11_u2_n152, u2_u11_u2_n153, u2_u11_u2_n154, u2_u11_u2_n155, u2_u11_u2_n156, u2_u11_u2_n157, u2_u11_u2_n158, u2_u11_u2_n159, 
       u2_u11_u2_n160, u2_u11_u2_n161, u2_u11_u2_n162, u2_u11_u2_n163, u2_u11_u2_n164, u2_u11_u2_n165, u2_u11_u2_n166, u2_u11_u2_n167, u2_u11_u2_n168, 
       u2_u11_u2_n169, u2_u11_u2_n170, u2_u11_u2_n171, u2_u11_u2_n172, u2_u11_u2_n173, u2_u11_u2_n174, u2_u11_u2_n175, u2_u11_u2_n176, u2_u11_u2_n177, 
       u2_u11_u2_n178, u2_u11_u2_n179, u2_u11_u2_n180, u2_u11_u2_n181, u2_u11_u2_n182, u2_u11_u2_n183, u2_u11_u2_n184, u2_u11_u2_n185, u2_u11_u2_n186, 
       u2_u11_u2_n187, u2_u11_u2_n188, u2_u11_u2_n95, u2_u11_u2_n96, u2_u11_u2_n97, u2_u11_u2_n98, u2_u11_u2_n99, u2_u11_u3_n100, u2_u11_u3_n101, 
       u2_u11_u3_n102, u2_u11_u3_n103, u2_u11_u3_n104, u2_u11_u3_n105, u2_u11_u3_n106, u2_u11_u3_n107, u2_u11_u3_n108, u2_u11_u3_n109, u2_u11_u3_n110, 
       u2_u11_u3_n111, u2_u11_u3_n112, u2_u11_u3_n113, u2_u11_u3_n114, u2_u11_u3_n115, u2_u11_u3_n116, u2_u11_u3_n117, u2_u11_u3_n118, u2_u11_u3_n119, 
       u2_u11_u3_n120, u2_u11_u3_n121, u2_u11_u3_n122, u2_u11_u3_n123, u2_u11_u3_n124, u2_u11_u3_n125, u2_u11_u3_n126, u2_u11_u3_n127, u2_u11_u3_n128, 
       u2_u11_u3_n129, u2_u11_u3_n130, u2_u11_u3_n131, u2_u11_u3_n132, u2_u11_u3_n133, u2_u11_u3_n134, u2_u11_u3_n135, u2_u11_u3_n136, u2_u11_u3_n137, 
       u2_u11_u3_n138, u2_u11_u3_n139, u2_u11_u3_n140, u2_u11_u3_n141, u2_u11_u3_n142, u2_u11_u3_n143, u2_u11_u3_n144, u2_u11_u3_n145, u2_u11_u3_n146, 
       u2_u11_u3_n147, u2_u11_u3_n148, u2_u11_u3_n149, u2_u11_u3_n150, u2_u11_u3_n151, u2_u11_u3_n152, u2_u11_u3_n153, u2_u11_u3_n154, u2_u11_u3_n155, 
       u2_u11_u3_n156, u2_u11_u3_n157, u2_u11_u3_n158, u2_u11_u3_n159, u2_u11_u3_n160, u2_u11_u3_n161, u2_u11_u3_n162, u2_u11_u3_n163, u2_u11_u3_n164, 
       u2_u11_u3_n165, u2_u11_u3_n166, u2_u11_u3_n167, u2_u11_u3_n168, u2_u11_u3_n169, u2_u11_u3_n170, u2_u11_u3_n171, u2_u11_u3_n172, u2_u11_u3_n173, 
       u2_u11_u3_n174, u2_u11_u3_n175, u2_u11_u3_n176, u2_u11_u3_n177, u2_u11_u3_n178, u2_u11_u3_n179, u2_u11_u3_n180, u2_u11_u3_n181, u2_u11_u3_n182, 
       u2_u11_u3_n183, u2_u11_u3_n184, u2_u11_u3_n185, u2_u11_u3_n186, u2_u11_u3_n94, u2_u11_u3_n95, u2_u11_u3_n96, u2_u11_u3_n97, u2_u11_u3_n98, 
       u2_u11_u3_n99, u2_u8_X_43, u2_u8_X_44, u2_u8_X_45, u2_u8_X_46, u2_u8_X_47, u2_u8_X_48, u2_u8_u7_n100, u2_u8_u7_n101, 
       u2_u8_u7_n102, u2_u8_u7_n103, u2_u8_u7_n104, u2_u8_u7_n105, u2_u8_u7_n106, u2_u8_u7_n107, u2_u8_u7_n108, u2_u8_u7_n109, u2_u8_u7_n110, 
       u2_u8_u7_n111, u2_u8_u7_n112, u2_u8_u7_n113, u2_u8_u7_n114, u2_u8_u7_n115, u2_u8_u7_n116, u2_u8_u7_n117, u2_u8_u7_n118, u2_u8_u7_n119, 
       u2_u8_u7_n120, u2_u8_u7_n121, u2_u8_u7_n122, u2_u8_u7_n123, u2_u8_u7_n124, u2_u8_u7_n125, u2_u8_u7_n126, u2_u8_u7_n127, u2_u8_u7_n128, 
       u2_u8_u7_n129, u2_u8_u7_n130, u2_u8_u7_n131, u2_u8_u7_n132, u2_u8_u7_n133, u2_u8_u7_n134, u2_u8_u7_n135, u2_u8_u7_n136, u2_u8_u7_n137, 
       u2_u8_u7_n138, u2_u8_u7_n139, u2_u8_u7_n140, u2_u8_u7_n141, u2_u8_u7_n142, u2_u8_u7_n143, u2_u8_u7_n144, u2_u8_u7_n145, u2_u8_u7_n146, 
       u2_u8_u7_n147, u2_u8_u7_n148, u2_u8_u7_n149, u2_u8_u7_n150, u2_u8_u7_n151, u2_u8_u7_n152, u2_u8_u7_n153, u2_u8_u7_n154, u2_u8_u7_n155, 
       u2_u8_u7_n156, u2_u8_u7_n157, u2_u8_u7_n158, u2_u8_u7_n159, u2_u8_u7_n160, u2_u8_u7_n161, u2_u8_u7_n162, u2_u8_u7_n163, u2_u8_u7_n164, 
       u2_u8_u7_n165, u2_u8_u7_n166, u2_u8_u7_n167, u2_u8_u7_n168, u2_u8_u7_n169, u2_u8_u7_n170, u2_u8_u7_n171, u2_u8_u7_n172, u2_u8_u7_n173, 
       u2_u8_u7_n174, u2_u8_u7_n175, u2_u8_u7_n176, u2_u8_u7_n177, u2_u8_u7_n178, u2_u8_u7_n179, u2_u8_u7_n180, u2_u8_u7_n91, u2_u8_u7_n92, 
       u2_u8_u7_n93, u2_u8_u7_n94, u2_u8_u7_n95, u2_u8_u7_n96, u2_u8_u7_n97, u2_u8_u7_n98, u2_u8_u7_n99, u2_uk_n1138, u2_uk_n1139, 
       u2_uk_n409,  u2_uk_n454;
  XOR2_X1 u0_U109 (.B( u0_L12_19 ) , .Z( u0_N434 ) , .A( u0_out13_19 ) );
  XOR2_X1 u0_U118 (.B( u0_L12_11 ) , .Z( u0_N426 ) , .A( u0_out13_11 ) );
  XOR2_X1 u0_U126 (.B( u0_L12_4 ) , .Z( u0_N419 ) , .A( u0_out13_4 ) );
  XOR2_X1 u0_U98 (.B( u0_L12_29 ) , .Z( u0_N444 ) , .A( u0_out13_29 ) );
  XOR2_X1 u0_u13_U20 (.B( u0_K14_36 ) , .A( u0_R12_25 ) , .Z( u0_u13_X_36 ) );
  XOR2_X1 u0_u13_U21 (.B( u0_K14_35 ) , .A( u0_R12_24 ) , .Z( u0_u13_X_35 ) );
  XOR2_X1 u0_u13_U22 (.B( u0_K14_34 ) , .A( u0_R12_23 ) , .Z( u0_u13_X_34 ) );
  XOR2_X1 u0_u13_U23 (.B( u0_K14_33 ) , .A( u0_R12_22 ) , .Z( u0_u13_X_33 ) );
  XOR2_X1 u0_u13_U24 (.B( u0_K14_32 ) , .A( u0_R12_21 ) , .Z( u0_u13_X_32 ) );
  XOR2_X1 u0_u13_U25 (.B( u0_K14_31 ) , .A( u0_R12_20 ) , .Z( u0_u13_X_31 ) );
  INV_X1 u0_u13_u5_U10 (.A( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U100 (.A3( u0_u13_u5_n141 ) , .A1( u0_u13_u5_n142 ) , .ZN( u0_u13_u5_n143 ) , .A2( u0_u13_u5_n191 ) );
  NAND4_X1 u0_u13_u5_U101 (.ZN( u0_out13_4 ) , .A4( u0_u13_u5_n112 ) , .A2( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n114 ) , .A3( u0_u13_u5_n195 ) );
  AOI211_X1 u0_u13_u5_U102 (.A( u0_u13_u5_n110 ) , .C1( u0_u13_u5_n111 ) , .ZN( u0_u13_u5_n112 ) , .B( u0_u13_u5_n118 ) , .C2( u0_u13_u5_n177 ) );
  AOI222_X1 u0_u13_u5_U103 (.ZN( u0_u13_u5_n113 ) , .A1( u0_u13_u5_n131 ) , .C1( u0_u13_u5_n148 ) , .B2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n178 ) , .A2( u0_u13_u5_n179 ) , .B1( u0_u13_u5_n99 ) );
  NAND3_X1 u0_u13_u5_U104 (.A2( u0_u13_u5_n154 ) , .A3( u0_u13_u5_n158 ) , .A1( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n99 ) );
  NOR2_X1 u0_u13_u5_U11 (.ZN( u0_u13_u5_n160 ) , .A2( u0_u13_u5_n173 ) , .A1( u0_u13_u5_n177 ) );
  INV_X1 u0_u13_u5_U12 (.A( u0_u13_u5_n150 ) , .ZN( u0_u13_u5_n174 ) );
  AOI21_X1 u0_u13_u5_U13 (.A( u0_u13_u5_n160 ) , .B2( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n162 ) , .B1( u0_u13_u5_n192 ) );
  INV_X1 u0_u13_u5_U14 (.A( u0_u13_u5_n159 ) , .ZN( u0_u13_u5_n192 ) );
  AOI21_X1 u0_u13_u5_U15 (.A( u0_u13_u5_n156 ) , .B2( u0_u13_u5_n157 ) , .B1( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n163 ) );
  AOI21_X1 u0_u13_u5_U16 (.B2( u0_u13_u5_n139 ) , .B1( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n141 ) , .A( u0_u13_u5_n150 ) );
  OAI21_X1 u0_u13_u5_U17 (.A( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n134 ) , .B1( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n142 ) );
  OAI21_X1 u0_u13_u5_U18 (.ZN( u0_u13_u5_n133 ) , .B2( u0_u13_u5_n147 ) , .A( u0_u13_u5_n173 ) , .B1( u0_u13_u5_n188 ) );
  NAND2_X1 u0_u13_u5_U19 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n137 ) );
  INV_X1 u0_u13_u5_U20 (.A( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n194 ) );
  NAND2_X1 u0_u13_u5_U21 (.A1( u0_u13_u5_n121 ) , .ZN( u0_u13_u5_n132 ) , .A2( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U22 (.A2( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n136 ) , .A1( u0_u13_u5_n154 ) );
  NAND2_X1 u0_u13_u5_U23 (.A2( u0_u13_u5_n119 ) , .A1( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n159 ) );
  INV_X1 u0_u13_u5_U24 (.A( u0_u13_u5_n156 ) , .ZN( u0_u13_u5_n175 ) );
  INV_X1 u0_u13_u5_U25 (.A( u0_u13_u5_n158 ) , .ZN( u0_u13_u5_n188 ) );
  INV_X1 u0_u13_u5_U26 (.A( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n179 ) );
  INV_X1 u0_u13_u5_U27 (.A( u0_u13_u5_n140 ) , .ZN( u0_u13_u5_n182 ) );
  INV_X1 u0_u13_u5_U28 (.A( u0_u13_u5_n151 ) , .ZN( u0_u13_u5_n183 ) );
  INV_X1 u0_u13_u5_U29 (.A( u0_u13_u5_n123 ) , .ZN( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U3 (.ZN( u0_u13_u5_n134 ) , .A1( u0_u13_u5_n183 ) , .A2( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U30 (.A( u0_u13_u5_n161 ) , .ZN( u0_u13_u5_n184 ) );
  INV_X1 u0_u13_u5_U31 (.A( u0_u13_u5_n139 ) , .ZN( u0_u13_u5_n189 ) );
  INV_X1 u0_u13_u5_U32 (.A( u0_u13_u5_n157 ) , .ZN( u0_u13_u5_n190 ) );
  INV_X1 u0_u13_u5_U33 (.A( u0_u13_u5_n120 ) , .ZN( u0_u13_u5_n193 ) );
  NAND2_X1 u0_u13_u5_U34 (.ZN( u0_u13_u5_n111 ) , .A1( u0_u13_u5_n140 ) , .A2( u0_u13_u5_n155 ) );
  INV_X1 u0_u13_u5_U35 (.A( u0_u13_u5_n117 ) , .ZN( u0_u13_u5_n196 ) );
  OAI221_X1 u0_u13_u5_U36 (.A( u0_u13_u5_n116 ) , .ZN( u0_u13_u5_n117 ) , .B2( u0_u13_u5_n119 ) , .C1( u0_u13_u5_n153 ) , .C2( u0_u13_u5_n158 ) , .B1( u0_u13_u5_n172 ) );
  AOI222_X1 u0_u13_u5_U37 (.ZN( u0_u13_u5_n116 ) , .B2( u0_u13_u5_n145 ) , .C1( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n174 ) , .C2( u0_u13_u5_n177 ) , .B1( u0_u13_u5_n187 ) , .A1( u0_u13_u5_n193 ) );
  INV_X1 u0_u13_u5_U38 (.A( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n187 ) );
  NOR2_X1 u0_u13_u5_U39 (.ZN( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n170 ) , .A2( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U4 (.A( u0_u13_u5_n138 ) , .ZN( u0_u13_u5_n191 ) );
  AOI22_X1 u0_u13_u5_U40 (.B2( u0_u13_u5_n131 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n169 ) , .B1( u0_u13_u5_n174 ) , .A1( u0_u13_u5_n185 ) );
  NOR2_X1 u0_u13_u5_U41 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n173 ) );
  AOI21_X1 u0_u13_u5_U42 (.A( u0_u13_u5_n118 ) , .B2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n168 ) , .B1( u0_u13_u5_n186 ) );
  INV_X1 u0_u13_u5_U43 (.A( u0_u13_u5_n122 ) , .ZN( u0_u13_u5_n186 ) );
  NOR2_X1 u0_u13_u5_U44 (.A1( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n152 ) , .A2( u0_u13_u5_n176 ) );
  NOR2_X1 u0_u13_u5_U45 (.A1( u0_u13_u5_n115 ) , .ZN( u0_u13_u5_n118 ) , .A2( u0_u13_u5_n153 ) );
  NOR2_X1 u0_u13_u5_U46 (.A2( u0_u13_u5_n145 ) , .ZN( u0_u13_u5_n156 ) , .A1( u0_u13_u5_n174 ) );
  NOR2_X1 u0_u13_u5_U47 (.ZN( u0_u13_u5_n121 ) , .A2( u0_u13_u5_n145 ) , .A1( u0_u13_u5_n176 ) );
  AOI22_X1 u0_u13_u5_U48 (.ZN( u0_u13_u5_n114 ) , .A2( u0_u13_u5_n137 ) , .A1( u0_u13_u5_n145 ) , .B2( u0_u13_u5_n175 ) , .B1( u0_u13_u5_n193 ) );
  OAI211_X1 u0_u13_u5_U49 (.B( u0_u13_u5_n124 ) , .A( u0_u13_u5_n125 ) , .C2( u0_u13_u5_n126 ) , .C1( u0_u13_u5_n127 ) , .ZN( u0_u13_u5_n128 ) );
  OAI21_X1 u0_u13_u5_U5 (.B2( u0_u13_u5_n136 ) , .B1( u0_u13_u5_n137 ) , .ZN( u0_u13_u5_n138 ) , .A( u0_u13_u5_n177 ) );
  NOR3_X1 u0_u13_u5_U50 (.ZN( u0_u13_u5_n127 ) , .A1( u0_u13_u5_n136 ) , .A3( u0_u13_u5_n148 ) , .A2( u0_u13_u5_n182 ) );
  OAI21_X1 u0_u13_u5_U51 (.ZN( u0_u13_u5_n124 ) , .A( u0_u13_u5_n177 ) , .B2( u0_u13_u5_n183 ) , .B1( u0_u13_u5_n189 ) );
  OAI21_X1 u0_u13_u5_U52 (.ZN( u0_u13_u5_n125 ) , .A( u0_u13_u5_n174 ) , .B2( u0_u13_u5_n185 ) , .B1( u0_u13_u5_n190 ) );
  AOI21_X1 u0_u13_u5_U53 (.A( u0_u13_u5_n153 ) , .B2( u0_u13_u5_n154 ) , .B1( u0_u13_u5_n155 ) , .ZN( u0_u13_u5_n164 ) );
  AOI21_X1 u0_u13_u5_U54 (.ZN( u0_u13_u5_n110 ) , .B1( u0_u13_u5_n122 ) , .B2( u0_u13_u5_n139 ) , .A( u0_u13_u5_n153 ) );
  INV_X1 u0_u13_u5_U55 (.A( u0_u13_u5_n153 ) , .ZN( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U56 (.A( u0_u13_u5_n126 ) , .ZN( u0_u13_u5_n173 ) );
  AND2_X1 u0_u13_u5_U57 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n147 ) );
  AND2_X1 u0_u13_u5_U58 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n148 ) );
  NAND2_X1 u0_u13_u5_U59 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n158 ) );
  INV_X1 u0_u13_u5_U6 (.A( u0_u13_u5_n135 ) , .ZN( u0_u13_u5_n178 ) );
  NAND2_X1 u0_u13_u5_U60 (.A2( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n139 ) );
  NAND2_X1 u0_u13_u5_U61 (.A1( u0_u13_u5_n106 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n119 ) );
  NAND2_X1 u0_u13_u5_U62 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n140 ) );
  NAND2_X1 u0_u13_u5_U63 (.A2( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n105 ) , .ZN( u0_u13_u5_n155 ) );
  NAND2_X1 u0_u13_u5_U64 (.A2( u0_u13_u5_n106 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n122 ) );
  NAND2_X1 u0_u13_u5_U65 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n106 ) , .ZN( u0_u13_u5_n115 ) );
  NAND2_X1 u0_u13_u5_U66 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n103 ) , .ZN( u0_u13_u5_n161 ) );
  NAND2_X1 u0_u13_u5_U67 (.A1( u0_u13_u5_n105 ) , .A2( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n154 ) );
  INV_X1 u0_u13_u5_U68 (.A( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n172 ) );
  NAND2_X1 u0_u13_u5_U69 (.A1( u0_u13_u5_n103 ) , .A2( u0_u13_u5_n108 ) , .ZN( u0_u13_u5_n123 ) );
  OAI22_X1 u0_u13_u5_U7 (.B2( u0_u13_u5_n149 ) , .B1( u0_u13_u5_n150 ) , .A2( u0_u13_u5_n151 ) , .A1( u0_u13_u5_n152 ) , .ZN( u0_u13_u5_n165 ) );
  NAND2_X1 u0_u13_u5_U70 (.A2( u0_u13_u5_n103 ) , .A1( u0_u13_u5_n107 ) , .ZN( u0_u13_u5_n151 ) );
  NAND2_X1 u0_u13_u5_U71 (.A2( u0_u13_u5_n107 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n120 ) );
  NAND2_X1 u0_u13_u5_U72 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n109 ) , .ZN( u0_u13_u5_n157 ) );
  AND2_X1 u0_u13_u5_U73 (.A2( u0_u13_u5_n100 ) , .A1( u0_u13_u5_n104 ) , .ZN( u0_u13_u5_n131 ) );
  INV_X1 u0_u13_u5_U74 (.A( u0_u13_u5_n102 ) , .ZN( u0_u13_u5_n195 ) );
  OAI221_X1 u0_u13_u5_U75 (.A( u0_u13_u5_n101 ) , .ZN( u0_u13_u5_n102 ) , .C2( u0_u13_u5_n115 ) , .C1( u0_u13_u5_n126 ) , .B1( u0_u13_u5_n134 ) , .B2( u0_u13_u5_n160 ) );
  OAI21_X1 u0_u13_u5_U76 (.ZN( u0_u13_u5_n101 ) , .B1( u0_u13_u5_n137 ) , .A( u0_u13_u5_n146 ) , .B2( u0_u13_u5_n147 ) );
  NOR2_X1 u0_u13_u5_U77 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n145 ) );
  NOR2_X1 u0_u13_u5_U78 (.A2( u0_u13_X_34 ) , .ZN( u0_u13_u5_n146 ) , .A1( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U79 (.A2( u0_u13_X_31 ) , .A1( u0_u13_X_32 ) , .ZN( u0_u13_u5_n103 ) );
  NOR3_X1 u0_u13_u5_U8 (.A2( u0_u13_u5_n147 ) , .A1( u0_u13_u5_n148 ) , .ZN( u0_u13_u5_n149 ) , .A3( u0_u13_u5_n194 ) );
  NOR2_X1 u0_u13_u5_U80 (.A2( u0_u13_X_36 ) , .ZN( u0_u13_u5_n105 ) , .A1( u0_u13_u5_n180 ) );
  NOR2_X1 u0_u13_u5_U81 (.A2( u0_u13_X_33 ) , .ZN( u0_u13_u5_n108 ) , .A1( u0_u13_u5_n170 ) );
  NOR2_X1 u0_u13_u5_U82 (.A2( u0_u13_X_33 ) , .A1( u0_u13_X_36 ) , .ZN( u0_u13_u5_n107 ) );
  NOR2_X1 u0_u13_u5_U83 (.A2( u0_u13_X_31 ) , .ZN( u0_u13_u5_n104 ) , .A1( u0_u13_u5_n181 ) );
  NAND2_X1 u0_u13_u5_U84 (.A2( u0_u13_X_34 ) , .A1( u0_u13_X_35 ) , .ZN( u0_u13_u5_n153 ) );
  NAND2_X1 u0_u13_u5_U85 (.A1( u0_u13_X_34 ) , .ZN( u0_u13_u5_n126 ) , .A2( u0_u13_u5_n171 ) );
  AND2_X1 u0_u13_u5_U86 (.A1( u0_u13_X_31 ) , .A2( u0_u13_X_32 ) , .ZN( u0_u13_u5_n106 ) );
  AND2_X1 u0_u13_u5_U87 (.A1( u0_u13_X_31 ) , .ZN( u0_u13_u5_n109 ) , .A2( u0_u13_u5_n181 ) );
  INV_X1 u0_u13_u5_U88 (.A( u0_u13_X_33 ) , .ZN( u0_u13_u5_n180 ) );
  INV_X1 u0_u13_u5_U89 (.A( u0_u13_X_35 ) , .ZN( u0_u13_u5_n171 ) );
  NOR2_X1 u0_u13_u5_U9 (.ZN( u0_u13_u5_n135 ) , .A1( u0_u13_u5_n173 ) , .A2( u0_u13_u5_n176 ) );
  INV_X1 u0_u13_u5_U90 (.A( u0_u13_X_36 ) , .ZN( u0_u13_u5_n170 ) );
  INV_X1 u0_u13_u5_U91 (.A( u0_u13_X_32 ) , .ZN( u0_u13_u5_n181 ) );
  NAND4_X1 u0_u13_u5_U92 (.ZN( u0_out13_29 ) , .A4( u0_u13_u5_n129 ) , .A3( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n196 ) );
  AOI221_X1 u0_u13_u5_U93 (.A( u0_u13_u5_n128 ) , .ZN( u0_u13_u5_n129 ) , .C2( u0_u13_u5_n132 ) , .B2( u0_u13_u5_n159 ) , .B1( u0_u13_u5_n176 ) , .C1( u0_u13_u5_n184 ) );
  AOI222_X1 u0_u13_u5_U94 (.ZN( u0_u13_u5_n130 ) , .A2( u0_u13_u5_n146 ) , .B1( u0_u13_u5_n147 ) , .C2( u0_u13_u5_n175 ) , .B2( u0_u13_u5_n179 ) , .A1( u0_u13_u5_n188 ) , .C1( u0_u13_u5_n194 ) );
  NAND4_X1 u0_u13_u5_U95 (.ZN( u0_out13_19 ) , .A4( u0_u13_u5_n166 ) , .A3( u0_u13_u5_n167 ) , .A2( u0_u13_u5_n168 ) , .A1( u0_u13_u5_n169 ) );
  AOI22_X1 u0_u13_u5_U96 (.B2( u0_u13_u5_n145 ) , .A2( u0_u13_u5_n146 ) , .ZN( u0_u13_u5_n167 ) , .B1( u0_u13_u5_n182 ) , .A1( u0_u13_u5_n189 ) );
  NOR4_X1 u0_u13_u5_U97 (.A4( u0_u13_u5_n162 ) , .A3( u0_u13_u5_n163 ) , .A2( u0_u13_u5_n164 ) , .A1( u0_u13_u5_n165 ) , .ZN( u0_u13_u5_n166 ) );
  NAND4_X1 u0_u13_u5_U98 (.ZN( u0_out13_11 ) , .A4( u0_u13_u5_n143 ) , .A3( u0_u13_u5_n144 ) , .A2( u0_u13_u5_n169 ) , .A1( u0_u13_u5_n196 ) );
  AOI22_X1 u0_u13_u5_U99 (.A2( u0_u13_u5_n132 ) , .ZN( u0_u13_u5_n144 ) , .B2( u0_u13_u5_n145 ) , .B1( u0_u13_u5_n184 ) , .A1( u0_u13_u5_n194 ) );
  OAI22_X1 u0_uk_U234 (.ZN( u0_K14_31 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n240 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n61 ) );
  OAI22_X1 u0_uk_U444 (.ZN( u0_K14_33 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n55 ) , .B2( u0_uk_n73 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U545 (.ZN( u0_K14_36 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n50 ) , .B2( u0_uk_n88 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U612 (.ZN( u0_K14_35 ) , .A( u0_uk_n933 ) );
  AOI22_X1 u0_uk_U613 (.B2( u0_uk_K_r12_1 ) , .A2( u0_uk_K_r12_7 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n933 ) );
  INV_X1 u0_uk_U65 (.ZN( u0_K14_34 ) , .A( u0_uk_n934 ) );
  AOI22_X1 u0_uk_U66 (.B2( u0_uk_K_r12_30 ) , .A2( u0_uk_K_r12_36 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n934 ) );
  OAI22_X1 u0_uk_U724 (.ZN( u0_K14_32 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n51 ) , .B2( u0_uk_n89 ) , .B1( u0_uk_n94 ) );
  XOR2_X1 u1_U10 (.B( u1_L1_29 ) , .Z( u1_N92 ) , .A( u1_out2_29 ) );
  XOR2_X1 u1_U125 (.B( u1_L0_11 ) , .Z( u1_N42 ) , .A( u1_out1_11 ) );
  XOR2_X1 u1_U15 (.B( u1_L1_25 ) , .Z( u1_N88 ) , .A( u1_out2_25 ) );
  XOR2_X1 u1_U168 (.B( u1_L10_30 ) , .Z( u1_N381 ) , .A( u1_out11_30 ) );
  XOR2_X1 u1_U173 (.B( u1_L10_26 ) , .Z( u1_N377 ) , .A( u1_out11_26 ) );
  XOR2_X1 u1_U175 (.B( u1_L10_24 ) , .Z( u1_N375 ) , .A( u1_out11_24 ) );
  XOR2_X1 u1_U179 (.B( u1_L10_20 ) , .Z( u1_N371 ) , .A( u1_out11_20 ) );
  XOR2_X1 u1_U184 (.B( u1_L10_16 ) , .Z( u1_N367 ) , .A( u1_out11_16 ) );
  XOR2_X1 u1_U190 (.B( u1_L10_10 ) , .Z( u1_N361 ) , .A( u1_out11_10 ) );
  XOR2_X1 u1_U195 (.B( u1_L10_6 ) , .Z( u1_N357 ) , .A( u1_out11_6 ) );
  XOR2_X1 u1_U200 (.B( u1_L10_1 ) , .Z( u1_N352 ) , .A( u1_out11_1 ) );
  XOR2_X1 u1_U203 (.B( u1_L0_4 ) , .Z( u1_N35 ) , .A( u1_out1_4 ) );
  XOR2_X1 u1_U21 (.B( u1_L1_19 ) , .Z( u1_N82 ) , .A( u1_out2_19 ) );
  XOR2_X1 u1_U27 (.B( u1_L1_14 ) , .Z( u1_N77 ) , .A( u1_out2_14 ) );
  XOR2_X1 u1_U30 (.B( u1_L1_11 ) , .Z( u1_N74 ) , .A( u1_out2_11 ) );
  XOR2_X1 u1_U33 (.B( u1_L1_8 ) , .Z( u1_N71 ) , .A( u1_out2_8 ) );
  XOR2_X1 u1_U38 (.B( u1_L1_4 ) , .Z( u1_N67 ) , .A( u1_out2_4 ) );
  XOR2_X1 u1_U384 (.B( u1_L4_28 ) , .Z( u1_N187 ) , .A( u1_out5_28 ) );
  XOR2_X1 u1_U385 (.B( u1_L4_27 ) , .Z( u1_N186 ) , .A( u1_out5_27 ) );
  XOR2_X1 u1_U39 (.B( u1_L1_3 ) , .Z( u1_N66 ) , .A( u1_out2_3 ) );
  XOR2_X1 u1_U391 (.B( u1_L4_21 ) , .Z( u1_N180 ) , .A( u1_out5_21 ) );
  XOR2_X1 u1_U395 (.B( u1_L4_18 ) , .Z( u1_N177 ) , .A( u1_out5_18 ) );
  XOR2_X1 u1_U398 (.B( u1_L4_15 ) , .Z( u1_N174 ) , .A( u1_out5_15 ) );
  XOR2_X1 u1_U400 (.B( u1_L4_13 ) , .Z( u1_N172 ) , .A( u1_out5_13 ) );
  XOR2_X1 u1_U409 (.B( u1_L4_5 ) , .Z( u1_N164 ) , .A( u1_out5_5 ) );
  XOR2_X1 u1_U412 (.B( u1_L4_2 ) , .Z( u1_N161 ) , .A( u1_out5_2 ) );
  XOR2_X1 u1_U415 (.B( u1_L3_32 ) , .Z( u1_N159 ) , .A( u1_out4_32 ) );
  XOR2_X1 u1_U426 (.B( u1_L3_22 ) , .Z( u1_N149 ) , .A( u1_out4_22 ) );
  XOR2_X1 u1_U437 (.B( u1_L3_12 ) , .Z( u1_N139 ) , .A( u1_out4_12 ) );
  XOR2_X1 u1_U442 (.B( u1_L3_7 ) , .Z( u1_N134 ) , .A( u1_out4_7 ) );
  XOR2_X1 u1_U45 (.B( u1_L0_29 ) , .Z( u1_N60 ) , .A( u1_out1_29 ) );
  XOR2_X1 u1_U56 (.B( u1_L0_19 ) , .Z( u1_N50 ) , .A( u1_out1_19 ) );
  XOR2_X1 u1_u11_U33 (.B( u1_K12_24 ) , .A( u1_R10_17 ) , .Z( u1_u11_X_24 ) );
  XOR2_X1 u1_u11_U34 (.B( u1_K12_23 ) , .A( u1_R10_16 ) , .Z( u1_u11_X_23 ) );
  XOR2_X1 u1_u11_U35 (.B( u1_K12_22 ) , .A( u1_R10_15 ) , .Z( u1_u11_X_22 ) );
  XOR2_X1 u1_u11_U36 (.B( u1_K12_21 ) , .A( u1_R10_14 ) , .Z( u1_u11_X_21 ) );
  XOR2_X1 u1_u11_U37 (.B( u1_K12_20 ) , .A( u1_R10_13 ) , .Z( u1_u11_X_20 ) );
  XOR2_X1 u1_u11_U39 (.B( u1_K12_19 ) , .A( u1_R10_12 ) , .Z( u1_u11_X_19 ) );
  XOR2_X1 u1_u11_U40 (.B( u1_K12_18 ) , .A( u1_R10_13 ) , .Z( u1_u11_X_18 ) );
  XOR2_X1 u1_u11_U41 (.B( u1_K12_17 ) , .A( u1_R10_12 ) , .Z( u1_u11_X_17 ) );
  XOR2_X1 u1_u11_U42 (.B( u1_K12_16 ) , .A( u1_R10_11 ) , .Z( u1_u11_X_16 ) );
  XOR2_X1 u1_u11_U43 (.B( u1_K12_15 ) , .A( u1_R10_10 ) , .Z( u1_u11_X_15 ) );
  XOR2_X1 u1_u11_U44 (.B( u1_K12_14 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_14 ) );
  XOR2_X1 u1_u11_U45 (.B( u1_K12_13 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_13 ) );
  OAI22_X1 u1_u11_u2_U10 (.ZN( u1_u11_u2_n109 ) , .A2( u1_u11_u2_n113 ) , .B2( u1_u11_u2_n133 ) , .B1( u1_u11_u2_n167 ) , .A1( u1_u11_u2_n168 ) );
  NAND3_X1 u1_u11_u2_U100 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n98 ) );
  OAI22_X1 u1_u11_u2_U11 (.B1( u1_u11_u2_n151 ) , .A2( u1_u11_u2_n152 ) , .A1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n160 ) , .B2( u1_u11_u2_n168 ) );
  NOR3_X1 u1_u11_u2_U12 (.A1( u1_u11_u2_n150 ) , .ZN( u1_u11_u2_n151 ) , .A3( u1_u11_u2_n175 ) , .A2( u1_u11_u2_n188 ) );
  AOI21_X1 u1_u11_u2_U13 (.ZN( u1_u11_u2_n144 ) , .B2( u1_u11_u2_n155 ) , .A( u1_u11_u2_n172 ) , .B1( u1_u11_u2_n185 ) );
  AOI21_X1 u1_u11_u2_U14 (.B2( u1_u11_u2_n143 ) , .ZN( u1_u11_u2_n145 ) , .B1( u1_u11_u2_n152 ) , .A( u1_u11_u2_n171 ) );
  AOI21_X1 u1_u11_u2_U15 (.B2( u1_u11_u2_n120 ) , .B1( u1_u11_u2_n121 ) , .ZN( u1_u11_u2_n126 ) , .A( u1_u11_u2_n167 ) );
  INV_X1 u1_u11_u2_U16 (.A( u1_u11_u2_n156 ) , .ZN( u1_u11_u2_n171 ) );
  INV_X1 u1_u11_u2_U17 (.A( u1_u11_u2_n120 ) , .ZN( u1_u11_u2_n188 ) );
  NAND2_X1 u1_u11_u2_U18 (.A2( u1_u11_u2_n122 ) , .ZN( u1_u11_u2_n150 ) , .A1( u1_u11_u2_n152 ) );
  INV_X1 u1_u11_u2_U19 (.A( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n170 ) );
  INV_X1 u1_u11_u2_U20 (.A( u1_u11_u2_n137 ) , .ZN( u1_u11_u2_n173 ) );
  NAND2_X1 u1_u11_u2_U21 (.A1( u1_u11_u2_n132 ) , .A2( u1_u11_u2_n139 ) , .ZN( u1_u11_u2_n157 ) );
  INV_X1 u1_u11_u2_U22 (.A( u1_u11_u2_n113 ) , .ZN( u1_u11_u2_n178 ) );
  INV_X1 u1_u11_u2_U23 (.A( u1_u11_u2_n139 ) , .ZN( u1_u11_u2_n175 ) );
  INV_X1 u1_u11_u2_U24 (.A( u1_u11_u2_n155 ) , .ZN( u1_u11_u2_n181 ) );
  INV_X1 u1_u11_u2_U25 (.A( u1_u11_u2_n119 ) , .ZN( u1_u11_u2_n177 ) );
  INV_X1 u1_u11_u2_U26 (.A( u1_u11_u2_n116 ) , .ZN( u1_u11_u2_n180 ) );
  INV_X1 u1_u11_u2_U27 (.A( u1_u11_u2_n131 ) , .ZN( u1_u11_u2_n179 ) );
  INV_X1 u1_u11_u2_U28 (.A( u1_u11_u2_n154 ) , .ZN( u1_u11_u2_n176 ) );
  NAND2_X1 u1_u11_u2_U29 (.A2( u1_u11_u2_n116 ) , .A1( u1_u11_u2_n117 ) , .ZN( u1_u11_u2_n118 ) );
  NOR2_X1 u1_u11_u2_U3 (.ZN( u1_u11_u2_n121 ) , .A2( u1_u11_u2_n177 ) , .A1( u1_u11_u2_n180 ) );
  INV_X1 u1_u11_u2_U30 (.A( u1_u11_u2_n132 ) , .ZN( u1_u11_u2_n182 ) );
  INV_X1 u1_u11_u2_U31 (.A( u1_u11_u2_n158 ) , .ZN( u1_u11_u2_n183 ) );
  OAI21_X1 u1_u11_u2_U32 (.A( u1_u11_u2_n156 ) , .B1( u1_u11_u2_n157 ) , .ZN( u1_u11_u2_n158 ) , .B2( u1_u11_u2_n179 ) );
  NOR2_X1 u1_u11_u2_U33 (.ZN( u1_u11_u2_n156 ) , .A1( u1_u11_u2_n166 ) , .A2( u1_u11_u2_n169 ) );
  NOR2_X1 u1_u11_u2_U34 (.A2( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n137 ) , .A1( u1_u11_u2_n140 ) );
  NOR2_X1 u1_u11_u2_U35 (.A2( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n153 ) , .A1( u1_u11_u2_n156 ) );
  AOI211_X1 u1_u11_u2_U36 (.ZN( u1_u11_u2_n130 ) , .C1( u1_u11_u2_n138 ) , .C2( u1_u11_u2_n179 ) , .B( u1_u11_u2_n96 ) , .A( u1_u11_u2_n97 ) );
  OAI22_X1 u1_u11_u2_U37 (.B1( u1_u11_u2_n133 ) , .A2( u1_u11_u2_n137 ) , .A1( u1_u11_u2_n152 ) , .B2( u1_u11_u2_n168 ) , .ZN( u1_u11_u2_n97 ) );
  OAI221_X1 u1_u11_u2_U38 (.B1( u1_u11_u2_n113 ) , .C1( u1_u11_u2_n132 ) , .A( u1_u11_u2_n149 ) , .B2( u1_u11_u2_n171 ) , .C2( u1_u11_u2_n172 ) , .ZN( u1_u11_u2_n96 ) );
  OAI221_X1 u1_u11_u2_U39 (.A( u1_u11_u2_n115 ) , .C2( u1_u11_u2_n123 ) , .B2( u1_u11_u2_n143 ) , .B1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n163 ) , .C1( u1_u11_u2_n168 ) );
  INV_X1 u1_u11_u2_U4 (.A( u1_u11_u2_n134 ) , .ZN( u1_u11_u2_n185 ) );
  OAI21_X1 u1_u11_u2_U40 (.A( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n115 ) , .B1( u1_u11_u2_n176 ) , .B2( u1_u11_u2_n178 ) );
  OAI221_X1 u1_u11_u2_U41 (.A( u1_u11_u2_n135 ) , .B2( u1_u11_u2_n136 ) , .B1( u1_u11_u2_n137 ) , .ZN( u1_u11_u2_n162 ) , .C2( u1_u11_u2_n167 ) , .C1( u1_u11_u2_n185 ) );
  AND3_X1 u1_u11_u2_U42 (.A3( u1_u11_u2_n131 ) , .A2( u1_u11_u2_n132 ) , .A1( u1_u11_u2_n133 ) , .ZN( u1_u11_u2_n136 ) );
  AOI22_X1 u1_u11_u2_U43 (.ZN( u1_u11_u2_n135 ) , .B1( u1_u11_u2_n140 ) , .A1( u1_u11_u2_n156 ) , .B2( u1_u11_u2_n180 ) , .A2( u1_u11_u2_n188 ) );
  AOI21_X1 u1_u11_u2_U44 (.ZN( u1_u11_u2_n149 ) , .B1( u1_u11_u2_n173 ) , .B2( u1_u11_u2_n188 ) , .A( u1_u11_u2_n95 ) );
  AND3_X1 u1_u11_u2_U45 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n156 ) , .ZN( u1_u11_u2_n95 ) );
  OAI21_X1 u1_u11_u2_U46 (.A( u1_u11_u2_n101 ) , .B2( u1_u11_u2_n121 ) , .B1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n164 ) );
  NAND2_X1 u1_u11_u2_U47 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n155 ) );
  NAND2_X1 u1_u11_u2_U48 (.A2( u1_u11_u2_n105 ) , .A1( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n143 ) );
  NAND2_X1 u1_u11_u2_U49 (.A1( u1_u11_u2_n104 ) , .A2( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n152 ) );
  INV_X1 u1_u11_u2_U5 (.A( u1_u11_u2_n150 ) , .ZN( u1_u11_u2_n184 ) );
  NAND2_X1 u1_u11_u2_U50 (.A1( u1_u11_u2_n100 ) , .A2( u1_u11_u2_n105 ) , .ZN( u1_u11_u2_n132 ) );
  INV_X1 u1_u11_u2_U51 (.A( u1_u11_u2_n140 ) , .ZN( u1_u11_u2_n168 ) );
  INV_X1 u1_u11_u2_U52 (.A( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n167 ) );
  OAI21_X1 u1_u11_u2_U53 (.A( u1_u11_u2_n141 ) , .B2( u1_u11_u2_n142 ) , .ZN( u1_u11_u2_n146 ) , .B1( u1_u11_u2_n153 ) );
  OAI21_X1 u1_u11_u2_U54 (.A( u1_u11_u2_n140 ) , .ZN( u1_u11_u2_n141 ) , .B1( u1_u11_u2_n176 ) , .B2( u1_u11_u2_n177 ) );
  NOR3_X1 u1_u11_u2_U55 (.ZN( u1_u11_u2_n142 ) , .A3( u1_u11_u2_n175 ) , .A2( u1_u11_u2_n178 ) , .A1( u1_u11_u2_n181 ) );
  INV_X1 u1_u11_u2_U56 (.ZN( u1_u11_u2_n187 ) , .A( u1_u11_u2_n99 ) );
  OAI21_X1 u1_u11_u2_U57 (.B1( u1_u11_u2_n137 ) , .B2( u1_u11_u2_n143 ) , .A( u1_u11_u2_n98 ) , .ZN( u1_u11_u2_n99 ) );
  NAND2_X1 u1_u11_u2_U58 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n113 ) );
  NAND2_X1 u1_u11_u2_U59 (.A1( u1_u11_u2_n106 ) , .A2( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n131 ) );
  NOR4_X1 u1_u11_u2_U6 (.A4( u1_u11_u2_n124 ) , .A3( u1_u11_u2_n125 ) , .A2( u1_u11_u2_n126 ) , .A1( u1_u11_u2_n127 ) , .ZN( u1_u11_u2_n128 ) );
  NAND2_X1 u1_u11_u2_U60 (.A1( u1_u11_u2_n103 ) , .A2( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n139 ) );
  NAND2_X1 u1_u11_u2_U61 (.A1( u1_u11_u2_n103 ) , .A2( u1_u11_u2_n105 ) , .ZN( u1_u11_u2_n133 ) );
  NAND2_X1 u1_u11_u2_U62 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n103 ) , .ZN( u1_u11_u2_n154 ) );
  NAND2_X1 u1_u11_u2_U63 (.A2( u1_u11_u2_n103 ) , .A1( u1_u11_u2_n104 ) , .ZN( u1_u11_u2_n119 ) );
  NAND2_X1 u1_u11_u2_U64 (.A2( u1_u11_u2_n107 ) , .A1( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n123 ) );
  NAND2_X1 u1_u11_u2_U65 (.A1( u1_u11_u2_n104 ) , .A2( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n122 ) );
  INV_X1 u1_u11_u2_U66 (.A( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n172 ) );
  NAND2_X1 u1_u11_u2_U67 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n102 ) , .ZN( u1_u11_u2_n116 ) );
  NAND2_X1 u1_u11_u2_U68 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n120 ) );
  NAND2_X1 u1_u11_u2_U69 (.A2( u1_u11_u2_n105 ) , .A1( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n117 ) );
  AOI21_X1 u1_u11_u2_U7 (.ZN( u1_u11_u2_n124 ) , .B1( u1_u11_u2_n131 ) , .B2( u1_u11_u2_n143 ) , .A( u1_u11_u2_n172 ) );
  NOR2_X1 u1_u11_u2_U70 (.A2( u1_u11_X_16 ) , .ZN( u1_u11_u2_n140 ) , .A1( u1_u11_u2_n166 ) );
  NOR2_X1 u1_u11_u2_U71 (.A2( u1_u11_X_13 ) , .A1( u1_u11_X_14 ) , .ZN( u1_u11_u2_n100 ) );
  NOR2_X1 u1_u11_u2_U72 (.A2( u1_u11_X_16 ) , .A1( u1_u11_X_17 ) , .ZN( u1_u11_u2_n138 ) );
  NOR2_X1 u1_u11_u2_U73 (.A2( u1_u11_X_15 ) , .A1( u1_u11_X_18 ) , .ZN( u1_u11_u2_n104 ) );
  NOR2_X1 u1_u11_u2_U74 (.A2( u1_u11_X_14 ) , .ZN( u1_u11_u2_n103 ) , .A1( u1_u11_u2_n174 ) );
  NOR2_X1 u1_u11_u2_U75 (.A2( u1_u11_X_15 ) , .ZN( u1_u11_u2_n102 ) , .A1( u1_u11_u2_n165 ) );
  NOR2_X1 u1_u11_u2_U76 (.A2( u1_u11_X_17 ) , .ZN( u1_u11_u2_n114 ) , .A1( u1_u11_u2_n169 ) );
  AND2_X1 u1_u11_u2_U77 (.A1( u1_u11_X_15 ) , .ZN( u1_u11_u2_n105 ) , .A2( u1_u11_u2_n165 ) );
  AND2_X1 u1_u11_u2_U78 (.A2( u1_u11_X_15 ) , .A1( u1_u11_X_18 ) , .ZN( u1_u11_u2_n107 ) );
  AND2_X1 u1_u11_u2_U79 (.A1( u1_u11_X_14 ) , .ZN( u1_u11_u2_n106 ) , .A2( u1_u11_u2_n174 ) );
  AOI21_X1 u1_u11_u2_U8 (.B2( u1_u11_u2_n119 ) , .ZN( u1_u11_u2_n127 ) , .A( u1_u11_u2_n137 ) , .B1( u1_u11_u2_n155 ) );
  AND2_X1 u1_u11_u2_U80 (.A1( u1_u11_X_13 ) , .A2( u1_u11_X_14 ) , .ZN( u1_u11_u2_n108 ) );
  INV_X1 u1_u11_u2_U81 (.A( u1_u11_X_16 ) , .ZN( u1_u11_u2_n169 ) );
  INV_X1 u1_u11_u2_U82 (.A( u1_u11_X_17 ) , .ZN( u1_u11_u2_n166 ) );
  INV_X1 u1_u11_u2_U83 (.A( u1_u11_X_13 ) , .ZN( u1_u11_u2_n174 ) );
  INV_X1 u1_u11_u2_U84 (.A( u1_u11_X_18 ) , .ZN( u1_u11_u2_n165 ) );
  NAND4_X1 u1_u11_u2_U85 (.ZN( u1_out11_30 ) , .A4( u1_u11_u2_n147 ) , .A3( u1_u11_u2_n148 ) , .A2( u1_u11_u2_n149 ) , .A1( u1_u11_u2_n187 ) );
  NOR3_X1 u1_u11_u2_U86 (.A3( u1_u11_u2_n144 ) , .A2( u1_u11_u2_n145 ) , .A1( u1_u11_u2_n146 ) , .ZN( u1_u11_u2_n147 ) );
  AOI21_X1 u1_u11_u2_U87 (.B2( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n148 ) , .A( u1_u11_u2_n162 ) , .B1( u1_u11_u2_n182 ) );
  NAND4_X1 u1_u11_u2_U88 (.ZN( u1_out11_24 ) , .A4( u1_u11_u2_n111 ) , .A3( u1_u11_u2_n112 ) , .A1( u1_u11_u2_n130 ) , .A2( u1_u11_u2_n187 ) );
  AOI221_X1 u1_u11_u2_U89 (.A( u1_u11_u2_n109 ) , .B1( u1_u11_u2_n110 ) , .ZN( u1_u11_u2_n111 ) , .C1( u1_u11_u2_n134 ) , .C2( u1_u11_u2_n170 ) , .B2( u1_u11_u2_n173 ) );
  AOI21_X1 u1_u11_u2_U9 (.B2( u1_u11_u2_n123 ) , .ZN( u1_u11_u2_n125 ) , .A( u1_u11_u2_n171 ) , .B1( u1_u11_u2_n184 ) );
  AOI21_X1 u1_u11_u2_U90 (.ZN( u1_u11_u2_n112 ) , .B2( u1_u11_u2_n156 ) , .A( u1_u11_u2_n164 ) , .B1( u1_u11_u2_n181 ) );
  NAND4_X1 u1_u11_u2_U91 (.ZN( u1_out11_16 ) , .A4( u1_u11_u2_n128 ) , .A3( u1_u11_u2_n129 ) , .A1( u1_u11_u2_n130 ) , .A2( u1_u11_u2_n186 ) );
  AOI22_X1 u1_u11_u2_U92 (.A2( u1_u11_u2_n118 ) , .ZN( u1_u11_u2_n129 ) , .A1( u1_u11_u2_n140 ) , .B1( u1_u11_u2_n157 ) , .B2( u1_u11_u2_n170 ) );
  INV_X1 u1_u11_u2_U93 (.A( u1_u11_u2_n163 ) , .ZN( u1_u11_u2_n186 ) );
  OR4_X1 u1_u11_u2_U94 (.ZN( u1_out11_6 ) , .A4( u1_u11_u2_n161 ) , .A3( u1_u11_u2_n162 ) , .A2( u1_u11_u2_n163 ) , .A1( u1_u11_u2_n164 ) );
  OR3_X1 u1_u11_u2_U95 (.A2( u1_u11_u2_n159 ) , .A1( u1_u11_u2_n160 ) , .ZN( u1_u11_u2_n161 ) , .A3( u1_u11_u2_n183 ) );
  AOI21_X1 u1_u11_u2_U96 (.B2( u1_u11_u2_n154 ) , .B1( u1_u11_u2_n155 ) , .ZN( u1_u11_u2_n159 ) , .A( u1_u11_u2_n167 ) );
  NAND3_X1 u1_u11_u2_U97 (.A2( u1_u11_u2_n117 ) , .A1( u1_u11_u2_n122 ) , .A3( u1_u11_u2_n123 ) , .ZN( u1_u11_u2_n134 ) );
  NAND3_X1 u1_u11_u2_U98 (.ZN( u1_u11_u2_n110 ) , .A2( u1_u11_u2_n131 ) , .A3( u1_u11_u2_n139 ) , .A1( u1_u11_u2_n154 ) );
  NAND3_X1 u1_u11_u2_U99 (.A2( u1_u11_u2_n100 ) , .ZN( u1_u11_u2_n101 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n114 ) );
  OAI211_X1 u1_u11_u3_U10 (.B( u1_u11_u3_n106 ) , .ZN( u1_u11_u3_n119 ) , .C2( u1_u11_u3_n128 ) , .C1( u1_u11_u3_n167 ) , .A( u1_u11_u3_n181 ) );
  INV_X1 u1_u11_u3_U11 (.ZN( u1_u11_u3_n181 ) , .A( u1_u11_u3_n98 ) );
  AOI221_X1 u1_u11_u3_U12 (.C1( u1_u11_u3_n105 ) , .ZN( u1_u11_u3_n106 ) , .A( u1_u11_u3_n131 ) , .B2( u1_u11_u3_n132 ) , .C2( u1_u11_u3_n133 ) , .B1( u1_u11_u3_n169 ) );
  OAI22_X1 u1_u11_u3_U13 (.B1( u1_u11_u3_n113 ) , .A2( u1_u11_u3_n135 ) , .A1( u1_u11_u3_n150 ) , .B2( u1_u11_u3_n164 ) , .ZN( u1_u11_u3_n98 ) );
  AOI22_X1 u1_u11_u3_U14 (.B1( u1_u11_u3_n115 ) , .A2( u1_u11_u3_n116 ) , .ZN( u1_u11_u3_n123 ) , .B2( u1_u11_u3_n133 ) , .A1( u1_u11_u3_n169 ) );
  NAND2_X1 u1_u11_u3_U15 (.ZN( u1_u11_u3_n116 ) , .A2( u1_u11_u3_n151 ) , .A1( u1_u11_u3_n182 ) );
  NOR2_X1 u1_u11_u3_U16 (.ZN( u1_u11_u3_n126 ) , .A2( u1_u11_u3_n150 ) , .A1( u1_u11_u3_n164 ) );
  AOI21_X1 u1_u11_u3_U17 (.ZN( u1_u11_u3_n112 ) , .B2( u1_u11_u3_n146 ) , .B1( u1_u11_u3_n155 ) , .A( u1_u11_u3_n167 ) );
  NAND2_X1 u1_u11_u3_U18 (.A1( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n142 ) , .A2( u1_u11_u3_n164 ) );
  NAND2_X1 u1_u11_u3_U19 (.ZN( u1_u11_u3_n132 ) , .A2( u1_u11_u3_n152 ) , .A1( u1_u11_u3_n156 ) );
  INV_X1 u1_u11_u3_U20 (.A( u1_u11_u3_n133 ) , .ZN( u1_u11_u3_n165 ) );
  AND2_X1 u1_u11_u3_U21 (.A2( u1_u11_u3_n113 ) , .A1( u1_u11_u3_n114 ) , .ZN( u1_u11_u3_n151 ) );
  INV_X1 u1_u11_u3_U22 (.A( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n170 ) );
  NAND2_X1 u1_u11_u3_U23 (.A1( u1_u11_u3_n107 ) , .A2( u1_u11_u3_n108 ) , .ZN( u1_u11_u3_n140 ) );
  NAND2_X1 u1_u11_u3_U24 (.ZN( u1_u11_u3_n117 ) , .A1( u1_u11_u3_n124 ) , .A2( u1_u11_u3_n148 ) );
  NAND2_X1 u1_u11_u3_U25 (.ZN( u1_u11_u3_n143 ) , .A1( u1_u11_u3_n165 ) , .A2( u1_u11_u3_n167 ) );
  INV_X1 u1_u11_u3_U26 (.A( u1_u11_u3_n130 ) , .ZN( u1_u11_u3_n177 ) );
  INV_X1 u1_u11_u3_U27 (.A( u1_u11_u3_n128 ) , .ZN( u1_u11_u3_n176 ) );
  NAND2_X1 u1_u11_u3_U28 (.ZN( u1_u11_u3_n105 ) , .A2( u1_u11_u3_n130 ) , .A1( u1_u11_u3_n155 ) );
  INV_X1 u1_u11_u3_U29 (.A( u1_u11_u3_n155 ) , .ZN( u1_u11_u3_n174 ) );
  INV_X1 u1_u11_u3_U3 (.A( u1_u11_u3_n140 ) , .ZN( u1_u11_u3_n182 ) );
  INV_X1 u1_u11_u3_U30 (.A( u1_u11_u3_n139 ) , .ZN( u1_u11_u3_n185 ) );
  NOR2_X1 u1_u11_u3_U31 (.ZN( u1_u11_u3_n135 ) , .A2( u1_u11_u3_n141 ) , .A1( u1_u11_u3_n169 ) );
  OAI222_X1 u1_u11_u3_U32 (.C2( u1_u11_u3_n107 ) , .A2( u1_u11_u3_n108 ) , .B1( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n138 ) , .B2( u1_u11_u3_n146 ) , .C1( u1_u11_u3_n154 ) , .A1( u1_u11_u3_n164 ) );
  NOR4_X1 u1_u11_u3_U33 (.A4( u1_u11_u3_n157 ) , .A3( u1_u11_u3_n158 ) , .A2( u1_u11_u3_n159 ) , .A1( u1_u11_u3_n160 ) , .ZN( u1_u11_u3_n161 ) );
  AOI21_X1 u1_u11_u3_U34 (.B2( u1_u11_u3_n152 ) , .B1( u1_u11_u3_n153 ) , .ZN( u1_u11_u3_n158 ) , .A( u1_u11_u3_n164 ) );
  AOI21_X1 u1_u11_u3_U35 (.A( u1_u11_u3_n154 ) , .B2( u1_u11_u3_n155 ) , .B1( u1_u11_u3_n156 ) , .ZN( u1_u11_u3_n157 ) );
  AOI21_X1 u1_u11_u3_U36 (.A( u1_u11_u3_n149 ) , .B2( u1_u11_u3_n150 ) , .B1( u1_u11_u3_n151 ) , .ZN( u1_u11_u3_n159 ) );
  AOI211_X1 u1_u11_u3_U37 (.ZN( u1_u11_u3_n109 ) , .A( u1_u11_u3_n119 ) , .C2( u1_u11_u3_n129 ) , .B( u1_u11_u3_n138 ) , .C1( u1_u11_u3_n141 ) );
  AOI211_X1 u1_u11_u3_U38 (.B( u1_u11_u3_n119 ) , .A( u1_u11_u3_n120 ) , .C2( u1_u11_u3_n121 ) , .ZN( u1_u11_u3_n122 ) , .C1( u1_u11_u3_n179 ) );
  INV_X1 u1_u11_u3_U39 (.A( u1_u11_u3_n156 ) , .ZN( u1_u11_u3_n179 ) );
  INV_X1 u1_u11_u3_U4 (.A( u1_u11_u3_n129 ) , .ZN( u1_u11_u3_n183 ) );
  OAI22_X1 u1_u11_u3_U40 (.B1( u1_u11_u3_n118 ) , .ZN( u1_u11_u3_n120 ) , .A1( u1_u11_u3_n135 ) , .B2( u1_u11_u3_n154 ) , .A2( u1_u11_u3_n178 ) );
  AND3_X1 u1_u11_u3_U41 (.ZN( u1_u11_u3_n118 ) , .A2( u1_u11_u3_n124 ) , .A1( u1_u11_u3_n144 ) , .A3( u1_u11_u3_n152 ) );
  INV_X1 u1_u11_u3_U42 (.A( u1_u11_u3_n121 ) , .ZN( u1_u11_u3_n164 ) );
  NAND2_X1 u1_u11_u3_U43 (.ZN( u1_u11_u3_n133 ) , .A1( u1_u11_u3_n154 ) , .A2( u1_u11_u3_n164 ) );
  NOR2_X1 u1_u11_u3_U44 (.A1( u1_u11_u3_n113 ) , .ZN( u1_u11_u3_n131 ) , .A2( u1_u11_u3_n154 ) );
  NAND2_X1 u1_u11_u3_U45 (.A1( u1_u11_u3_n103 ) , .ZN( u1_u11_u3_n150 ) , .A2( u1_u11_u3_n99 ) );
  NAND2_X1 u1_u11_u3_U46 (.A2( u1_u11_u3_n102 ) , .ZN( u1_u11_u3_n155 ) , .A1( u1_u11_u3_n97 ) );
  OAI211_X1 u1_u11_u3_U47 (.B( u1_u11_u3_n127 ) , .ZN( u1_u11_u3_n139 ) , .C1( u1_u11_u3_n150 ) , .C2( u1_u11_u3_n154 ) , .A( u1_u11_u3_n184 ) );
  INV_X1 u1_u11_u3_U48 (.A( u1_u11_u3_n125 ) , .ZN( u1_u11_u3_n184 ) );
  AOI221_X1 u1_u11_u3_U49 (.A( u1_u11_u3_n126 ) , .ZN( u1_u11_u3_n127 ) , .C2( u1_u11_u3_n132 ) , .C1( u1_u11_u3_n169 ) , .B2( u1_u11_u3_n170 ) , .B1( u1_u11_u3_n174 ) );
  INV_X1 u1_u11_u3_U5 (.A( u1_u11_u3_n117 ) , .ZN( u1_u11_u3_n178 ) );
  OAI22_X1 u1_u11_u3_U50 (.A1( u1_u11_u3_n124 ) , .ZN( u1_u11_u3_n125 ) , .B2( u1_u11_u3_n145 ) , .A2( u1_u11_u3_n165 ) , .B1( u1_u11_u3_n167 ) );
  INV_X1 u1_u11_u3_U51 (.A( u1_u11_u3_n141 ) , .ZN( u1_u11_u3_n167 ) );
  AOI21_X1 u1_u11_u3_U52 (.B2( u1_u11_u3_n114 ) , .B1( u1_u11_u3_n146 ) , .A( u1_u11_u3_n154 ) , .ZN( u1_u11_u3_n94 ) );
  AOI21_X1 u1_u11_u3_U53 (.ZN( u1_u11_u3_n110 ) , .B2( u1_u11_u3_n142 ) , .B1( u1_u11_u3_n186 ) , .A( u1_u11_u3_n95 ) );
  INV_X1 u1_u11_u3_U54 (.A( u1_u11_u3_n145 ) , .ZN( u1_u11_u3_n186 ) );
  AOI21_X1 u1_u11_u3_U55 (.B1( u1_u11_u3_n124 ) , .A( u1_u11_u3_n149 ) , .B2( u1_u11_u3_n155 ) , .ZN( u1_u11_u3_n95 ) );
  INV_X1 u1_u11_u3_U56 (.A( u1_u11_u3_n149 ) , .ZN( u1_u11_u3_n169 ) );
  NAND2_X1 u1_u11_u3_U57 (.ZN( u1_u11_u3_n124 ) , .A1( u1_u11_u3_n96 ) , .A2( u1_u11_u3_n97 ) );
  NAND2_X1 u1_u11_u3_U58 (.A2( u1_u11_u3_n100 ) , .ZN( u1_u11_u3_n146 ) , .A1( u1_u11_u3_n96 ) );
  NAND2_X1 u1_u11_u3_U59 (.A1( u1_u11_u3_n101 ) , .ZN( u1_u11_u3_n145 ) , .A2( u1_u11_u3_n99 ) );
  AOI221_X1 u1_u11_u3_U6 (.A( u1_u11_u3_n131 ) , .C2( u1_u11_u3_n132 ) , .C1( u1_u11_u3_n133 ) , .ZN( u1_u11_u3_n134 ) , .B1( u1_u11_u3_n143 ) , .B2( u1_u11_u3_n177 ) );
  NAND2_X1 u1_u11_u3_U60 (.A1( u1_u11_u3_n100 ) , .ZN( u1_u11_u3_n156 ) , .A2( u1_u11_u3_n99 ) );
  NAND2_X1 u1_u11_u3_U61 (.A2( u1_u11_u3_n101 ) , .A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n148 ) );
  NAND2_X1 u1_u11_u3_U62 (.A1( u1_u11_u3_n100 ) , .A2( u1_u11_u3_n102 ) , .ZN( u1_u11_u3_n128 ) );
  NAND2_X1 u1_u11_u3_U63 (.A2( u1_u11_u3_n101 ) , .A1( u1_u11_u3_n102 ) , .ZN( u1_u11_u3_n152 ) );
  NAND2_X1 u1_u11_u3_U64 (.A2( u1_u11_u3_n101 ) , .ZN( u1_u11_u3_n114 ) , .A1( u1_u11_u3_n96 ) );
  NAND2_X1 u1_u11_u3_U65 (.ZN( u1_u11_u3_n107 ) , .A1( u1_u11_u3_n97 ) , .A2( u1_u11_u3_n99 ) );
  NAND2_X1 u1_u11_u3_U66 (.A2( u1_u11_u3_n100 ) , .A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n113 ) );
  NAND2_X1 u1_u11_u3_U67 (.A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n153 ) , .A2( u1_u11_u3_n97 ) );
  NAND2_X1 u1_u11_u3_U68 (.A2( u1_u11_u3_n103 ) , .A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n130 ) );
  NAND2_X1 u1_u11_u3_U69 (.A2( u1_u11_u3_n103 ) , .ZN( u1_u11_u3_n144 ) , .A1( u1_u11_u3_n96 ) );
  OAI22_X1 u1_u11_u3_U7 (.B2( u1_u11_u3_n147 ) , .A2( u1_u11_u3_n148 ) , .ZN( u1_u11_u3_n160 ) , .B1( u1_u11_u3_n165 ) , .A1( u1_u11_u3_n168 ) );
  NAND2_X1 u1_u11_u3_U70 (.A1( u1_u11_u3_n102 ) , .A2( u1_u11_u3_n103 ) , .ZN( u1_u11_u3_n108 ) );
  NOR2_X1 u1_u11_u3_U71 (.A2( u1_u11_X_19 ) , .A1( u1_u11_X_20 ) , .ZN( u1_u11_u3_n99 ) );
  NOR2_X1 u1_u11_u3_U72 (.A2( u1_u11_X_21 ) , .A1( u1_u11_X_24 ) , .ZN( u1_u11_u3_n103 ) );
  NOR2_X1 u1_u11_u3_U73 (.A2( u1_u11_X_24 ) , .A1( u1_u11_u3_n171 ) , .ZN( u1_u11_u3_n97 ) );
  NOR2_X1 u1_u11_u3_U74 (.A2( u1_u11_X_23 ) , .ZN( u1_u11_u3_n141 ) , .A1( u1_u11_u3_n166 ) );
  NOR2_X1 u1_u11_u3_U75 (.A2( u1_u11_X_19 ) , .A1( u1_u11_u3_n172 ) , .ZN( u1_u11_u3_n96 ) );
  NAND2_X1 u1_u11_u3_U76 (.A1( u1_u11_X_22 ) , .A2( u1_u11_X_23 ) , .ZN( u1_u11_u3_n154 ) );
  NAND2_X1 u1_u11_u3_U77 (.A1( u1_u11_X_23 ) , .ZN( u1_u11_u3_n149 ) , .A2( u1_u11_u3_n166 ) );
  NOR2_X1 u1_u11_u3_U78 (.A2( u1_u11_X_22 ) , .A1( u1_u11_X_23 ) , .ZN( u1_u11_u3_n121 ) );
  AND2_X1 u1_u11_u3_U79 (.A1( u1_u11_X_24 ) , .ZN( u1_u11_u3_n101 ) , .A2( u1_u11_u3_n171 ) );
  AND3_X1 u1_u11_u3_U8 (.A3( u1_u11_u3_n144 ) , .A2( u1_u11_u3_n145 ) , .A1( u1_u11_u3_n146 ) , .ZN( u1_u11_u3_n147 ) );
  AND2_X1 u1_u11_u3_U80 (.A1( u1_u11_X_19 ) , .ZN( u1_u11_u3_n102 ) , .A2( u1_u11_u3_n172 ) );
  AND2_X1 u1_u11_u3_U81 (.A1( u1_u11_X_21 ) , .A2( u1_u11_X_24 ) , .ZN( u1_u11_u3_n100 ) );
  AND2_X1 u1_u11_u3_U82 (.A2( u1_u11_X_19 ) , .A1( u1_u11_X_20 ) , .ZN( u1_u11_u3_n104 ) );
  INV_X1 u1_u11_u3_U83 (.A( u1_u11_X_22 ) , .ZN( u1_u11_u3_n166 ) );
  INV_X1 u1_u11_u3_U84 (.A( u1_u11_X_21 ) , .ZN( u1_u11_u3_n171 ) );
  INV_X1 u1_u11_u3_U85 (.A( u1_u11_X_20 ) , .ZN( u1_u11_u3_n172 ) );
  NAND4_X1 u1_u11_u3_U86 (.ZN( u1_out11_26 ) , .A4( u1_u11_u3_n109 ) , .A3( u1_u11_u3_n110 ) , .A2( u1_u11_u3_n111 ) , .A1( u1_u11_u3_n173 ) );
  INV_X1 u1_u11_u3_U87 (.ZN( u1_u11_u3_n173 ) , .A( u1_u11_u3_n94 ) );
  OAI21_X1 u1_u11_u3_U88 (.ZN( u1_u11_u3_n111 ) , .B2( u1_u11_u3_n117 ) , .A( u1_u11_u3_n133 ) , .B1( u1_u11_u3_n176 ) );
  NAND4_X1 u1_u11_u3_U89 (.ZN( u1_out11_20 ) , .A4( u1_u11_u3_n122 ) , .A3( u1_u11_u3_n123 ) , .A1( u1_u11_u3_n175 ) , .A2( u1_u11_u3_n180 ) );
  INV_X1 u1_u11_u3_U9 (.A( u1_u11_u3_n143 ) , .ZN( u1_u11_u3_n168 ) );
  INV_X1 u1_u11_u3_U90 (.A( u1_u11_u3_n126 ) , .ZN( u1_u11_u3_n180 ) );
  INV_X1 u1_u11_u3_U91 (.A( u1_u11_u3_n112 ) , .ZN( u1_u11_u3_n175 ) );
  OAI222_X1 u1_u11_u3_U92 (.C1( u1_u11_u3_n128 ) , .ZN( u1_u11_u3_n137 ) , .B1( u1_u11_u3_n148 ) , .A2( u1_u11_u3_n150 ) , .B2( u1_u11_u3_n154 ) , .C2( u1_u11_u3_n164 ) , .A1( u1_u11_u3_n167 ) );
  NAND4_X1 u1_u11_u3_U93 (.ZN( u1_out11_1 ) , .A4( u1_u11_u3_n161 ) , .A3( u1_u11_u3_n162 ) , .A2( u1_u11_u3_n163 ) , .A1( u1_u11_u3_n185 ) );
  NAND2_X1 u1_u11_u3_U94 (.ZN( u1_u11_u3_n163 ) , .A2( u1_u11_u3_n170 ) , .A1( u1_u11_u3_n176 ) );
  AOI22_X1 u1_u11_u3_U95 (.B2( u1_u11_u3_n140 ) , .B1( u1_u11_u3_n141 ) , .A2( u1_u11_u3_n142 ) , .ZN( u1_u11_u3_n162 ) , .A1( u1_u11_u3_n177 ) );
  OR4_X1 u1_u11_u3_U96 (.ZN( u1_out11_10 ) , .A4( u1_u11_u3_n136 ) , .A3( u1_u11_u3_n137 ) , .A1( u1_u11_u3_n138 ) , .A2( u1_u11_u3_n139 ) );
  OAI221_X1 u1_u11_u3_U97 (.A( u1_u11_u3_n134 ) , .B2( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n136 ) , .C1( u1_u11_u3_n149 ) , .B1( u1_u11_u3_n151 ) , .C2( u1_u11_u3_n183 ) );
  NAND3_X1 u1_u11_u3_U98 (.A1( u1_u11_u3_n114 ) , .ZN( u1_u11_u3_n115 ) , .A2( u1_u11_u3_n145 ) , .A3( u1_u11_u3_n153 ) );
  NAND3_X1 u1_u11_u3_U99 (.ZN( u1_u11_u3_n129 ) , .A2( u1_u11_u3_n144 ) , .A1( u1_u11_u3_n153 ) , .A3( u1_u11_u3_n182 ) );
  XOR2_X1 u1_u1_U20 (.B( u1_K2_36 ) , .A( u1_R0_25 ) , .Z( u1_u1_X_36 ) );
  XOR2_X1 u1_u1_U21 (.B( u1_K2_35 ) , .A( u1_R0_24 ) , .Z( u1_u1_X_35 ) );
  XOR2_X1 u1_u1_U22 (.B( u1_K2_34 ) , .A( u1_R0_23 ) , .Z( u1_u1_X_34 ) );
  XOR2_X1 u1_u1_U23 (.B( u1_K2_33 ) , .A( u1_R0_22 ) , .Z( u1_u1_X_33 ) );
  XOR2_X1 u1_u1_U24 (.B( u1_K2_32 ) , .A( u1_R0_21 ) , .Z( u1_u1_X_32 ) );
  XOR2_X1 u1_u1_U25 (.B( u1_K2_31 ) , .A( u1_R0_20 ) , .Z( u1_u1_X_31 ) );
  INV_X1 u1_u1_u5_U10 (.A( u1_u1_u5_n121 ) , .ZN( u1_u1_u5_n177 ) );
  NOR3_X1 u1_u1_u5_U100 (.A3( u1_u1_u5_n141 ) , .A1( u1_u1_u5_n142 ) , .ZN( u1_u1_u5_n143 ) , .A2( u1_u1_u5_n191 ) );
  NAND4_X1 u1_u1_u5_U101 (.ZN( u1_out1_4 ) , .A4( u1_u1_u5_n112 ) , .A2( u1_u1_u5_n113 ) , .A1( u1_u1_u5_n114 ) , .A3( u1_u1_u5_n195 ) );
  AOI211_X1 u1_u1_u5_U102 (.A( u1_u1_u5_n110 ) , .C1( u1_u1_u5_n111 ) , .ZN( u1_u1_u5_n112 ) , .B( u1_u1_u5_n118 ) , .C2( u1_u1_u5_n177 ) );
  AOI222_X1 u1_u1_u5_U103 (.ZN( u1_u1_u5_n113 ) , .A1( u1_u1_u5_n131 ) , .C1( u1_u1_u5_n148 ) , .B2( u1_u1_u5_n174 ) , .C2( u1_u1_u5_n178 ) , .A2( u1_u1_u5_n179 ) , .B1( u1_u1_u5_n99 ) );
  NAND3_X1 u1_u1_u5_U104 (.A2( u1_u1_u5_n154 ) , .A3( u1_u1_u5_n158 ) , .A1( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n99 ) );
  NOR2_X1 u1_u1_u5_U11 (.ZN( u1_u1_u5_n160 ) , .A2( u1_u1_u5_n173 ) , .A1( u1_u1_u5_n177 ) );
  INV_X1 u1_u1_u5_U12 (.A( u1_u1_u5_n150 ) , .ZN( u1_u1_u5_n174 ) );
  AOI21_X1 u1_u1_u5_U13 (.A( u1_u1_u5_n160 ) , .B2( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n162 ) , .B1( u1_u1_u5_n192 ) );
  INV_X1 u1_u1_u5_U14 (.A( u1_u1_u5_n159 ) , .ZN( u1_u1_u5_n192 ) );
  AOI21_X1 u1_u1_u5_U15 (.A( u1_u1_u5_n156 ) , .B2( u1_u1_u5_n157 ) , .B1( u1_u1_u5_n158 ) , .ZN( u1_u1_u5_n163 ) );
  AOI21_X1 u1_u1_u5_U16 (.B2( u1_u1_u5_n139 ) , .B1( u1_u1_u5_n140 ) , .ZN( u1_u1_u5_n141 ) , .A( u1_u1_u5_n150 ) );
  OAI21_X1 u1_u1_u5_U17 (.A( u1_u1_u5_n133 ) , .B2( u1_u1_u5_n134 ) , .B1( u1_u1_u5_n135 ) , .ZN( u1_u1_u5_n142 ) );
  OAI21_X1 u1_u1_u5_U18 (.ZN( u1_u1_u5_n133 ) , .B2( u1_u1_u5_n147 ) , .A( u1_u1_u5_n173 ) , .B1( u1_u1_u5_n188 ) );
  NAND2_X1 u1_u1_u5_U19 (.A2( u1_u1_u5_n119 ) , .A1( u1_u1_u5_n123 ) , .ZN( u1_u1_u5_n137 ) );
  INV_X1 u1_u1_u5_U20 (.A( u1_u1_u5_n155 ) , .ZN( u1_u1_u5_n194 ) );
  NAND2_X1 u1_u1_u5_U21 (.A1( u1_u1_u5_n121 ) , .ZN( u1_u1_u5_n132 ) , .A2( u1_u1_u5_n172 ) );
  NAND2_X1 u1_u1_u5_U22 (.A2( u1_u1_u5_n122 ) , .ZN( u1_u1_u5_n136 ) , .A1( u1_u1_u5_n154 ) );
  NAND2_X1 u1_u1_u5_U23 (.A2( u1_u1_u5_n119 ) , .A1( u1_u1_u5_n120 ) , .ZN( u1_u1_u5_n159 ) );
  INV_X1 u1_u1_u5_U24 (.A( u1_u1_u5_n156 ) , .ZN( u1_u1_u5_n175 ) );
  INV_X1 u1_u1_u5_U25 (.A( u1_u1_u5_n158 ) , .ZN( u1_u1_u5_n188 ) );
  INV_X1 u1_u1_u5_U26 (.A( u1_u1_u5_n152 ) , .ZN( u1_u1_u5_n179 ) );
  INV_X1 u1_u1_u5_U27 (.A( u1_u1_u5_n140 ) , .ZN( u1_u1_u5_n182 ) );
  INV_X1 u1_u1_u5_U28 (.A( u1_u1_u5_n151 ) , .ZN( u1_u1_u5_n183 ) );
  INV_X1 u1_u1_u5_U29 (.A( u1_u1_u5_n123 ) , .ZN( u1_u1_u5_n185 ) );
  NOR2_X1 u1_u1_u5_U3 (.ZN( u1_u1_u5_n134 ) , .A1( u1_u1_u5_n183 ) , .A2( u1_u1_u5_n190 ) );
  INV_X1 u1_u1_u5_U30 (.A( u1_u1_u5_n161 ) , .ZN( u1_u1_u5_n184 ) );
  INV_X1 u1_u1_u5_U31 (.A( u1_u1_u5_n139 ) , .ZN( u1_u1_u5_n189 ) );
  INV_X1 u1_u1_u5_U32 (.A( u1_u1_u5_n157 ) , .ZN( u1_u1_u5_n190 ) );
  INV_X1 u1_u1_u5_U33 (.A( u1_u1_u5_n120 ) , .ZN( u1_u1_u5_n193 ) );
  NAND2_X1 u1_u1_u5_U34 (.ZN( u1_u1_u5_n111 ) , .A1( u1_u1_u5_n140 ) , .A2( u1_u1_u5_n155 ) );
  INV_X1 u1_u1_u5_U35 (.A( u1_u1_u5_n117 ) , .ZN( u1_u1_u5_n196 ) );
  OAI221_X1 u1_u1_u5_U36 (.A( u1_u1_u5_n116 ) , .ZN( u1_u1_u5_n117 ) , .B2( u1_u1_u5_n119 ) , .C1( u1_u1_u5_n153 ) , .C2( u1_u1_u5_n158 ) , .B1( u1_u1_u5_n172 ) );
  AOI222_X1 u1_u1_u5_U37 (.ZN( u1_u1_u5_n116 ) , .B2( u1_u1_u5_n145 ) , .C1( u1_u1_u5_n148 ) , .A2( u1_u1_u5_n174 ) , .C2( u1_u1_u5_n177 ) , .B1( u1_u1_u5_n187 ) , .A1( u1_u1_u5_n193 ) );
  INV_X1 u1_u1_u5_U38 (.A( u1_u1_u5_n115 ) , .ZN( u1_u1_u5_n187 ) );
  NOR2_X1 u1_u1_u5_U39 (.ZN( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n170 ) , .A2( u1_u1_u5_n180 ) );
  INV_X1 u1_u1_u5_U4 (.A( u1_u1_u5_n138 ) , .ZN( u1_u1_u5_n191 ) );
  AOI22_X1 u1_u1_u5_U40 (.B2( u1_u1_u5_n131 ) , .A2( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n169 ) , .B1( u1_u1_u5_n174 ) , .A1( u1_u1_u5_n185 ) );
  NOR2_X1 u1_u1_u5_U41 (.A1( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n150 ) , .A2( u1_u1_u5_n173 ) );
  AOI21_X1 u1_u1_u5_U42 (.A( u1_u1_u5_n118 ) , .B2( u1_u1_u5_n145 ) , .ZN( u1_u1_u5_n168 ) , .B1( u1_u1_u5_n186 ) );
  INV_X1 u1_u1_u5_U43 (.A( u1_u1_u5_n122 ) , .ZN( u1_u1_u5_n186 ) );
  NOR2_X1 u1_u1_u5_U44 (.A1( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n152 ) , .A2( u1_u1_u5_n176 ) );
  NOR2_X1 u1_u1_u5_U45 (.A1( u1_u1_u5_n115 ) , .ZN( u1_u1_u5_n118 ) , .A2( u1_u1_u5_n153 ) );
  NOR2_X1 u1_u1_u5_U46 (.A2( u1_u1_u5_n145 ) , .ZN( u1_u1_u5_n156 ) , .A1( u1_u1_u5_n174 ) );
  NOR2_X1 u1_u1_u5_U47 (.ZN( u1_u1_u5_n121 ) , .A2( u1_u1_u5_n145 ) , .A1( u1_u1_u5_n176 ) );
  AOI22_X1 u1_u1_u5_U48 (.ZN( u1_u1_u5_n114 ) , .A2( u1_u1_u5_n137 ) , .A1( u1_u1_u5_n145 ) , .B2( u1_u1_u5_n175 ) , .B1( u1_u1_u5_n193 ) );
  OAI211_X1 u1_u1_u5_U49 (.B( u1_u1_u5_n124 ) , .A( u1_u1_u5_n125 ) , .C2( u1_u1_u5_n126 ) , .C1( u1_u1_u5_n127 ) , .ZN( u1_u1_u5_n128 ) );
  OAI21_X1 u1_u1_u5_U5 (.B2( u1_u1_u5_n136 ) , .B1( u1_u1_u5_n137 ) , .ZN( u1_u1_u5_n138 ) , .A( u1_u1_u5_n177 ) );
  OAI21_X1 u1_u1_u5_U50 (.ZN( u1_u1_u5_n124 ) , .A( u1_u1_u5_n177 ) , .B2( u1_u1_u5_n183 ) , .B1( u1_u1_u5_n189 ) );
  NOR3_X1 u1_u1_u5_U51 (.ZN( u1_u1_u5_n127 ) , .A1( u1_u1_u5_n136 ) , .A3( u1_u1_u5_n148 ) , .A2( u1_u1_u5_n182 ) );
  OAI21_X1 u1_u1_u5_U52 (.ZN( u1_u1_u5_n125 ) , .A( u1_u1_u5_n174 ) , .B2( u1_u1_u5_n185 ) , .B1( u1_u1_u5_n190 ) );
  AOI21_X1 u1_u1_u5_U53 (.A( u1_u1_u5_n153 ) , .B2( u1_u1_u5_n154 ) , .B1( u1_u1_u5_n155 ) , .ZN( u1_u1_u5_n164 ) );
  AOI21_X1 u1_u1_u5_U54 (.ZN( u1_u1_u5_n110 ) , .B1( u1_u1_u5_n122 ) , .B2( u1_u1_u5_n139 ) , .A( u1_u1_u5_n153 ) );
  INV_X1 u1_u1_u5_U55 (.A( u1_u1_u5_n153 ) , .ZN( u1_u1_u5_n176 ) );
  INV_X1 u1_u1_u5_U56 (.A( u1_u1_u5_n126 ) , .ZN( u1_u1_u5_n173 ) );
  AND2_X1 u1_u1_u5_U57 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n147 ) );
  AND2_X1 u1_u1_u5_U58 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n148 ) );
  NAND2_X1 u1_u1_u5_U59 (.A1( u1_u1_u5_n105 ) , .A2( u1_u1_u5_n106 ) , .ZN( u1_u1_u5_n158 ) );
  INV_X1 u1_u1_u5_U6 (.A( u1_u1_u5_n135 ) , .ZN( u1_u1_u5_n178 ) );
  NAND2_X1 u1_u1_u5_U60 (.A2( u1_u1_u5_n108 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n139 ) );
  NAND2_X1 u1_u1_u5_U61 (.A1( u1_u1_u5_n106 ) , .A2( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n119 ) );
  NAND2_X1 u1_u1_u5_U62 (.A2( u1_u1_u5_n103 ) , .A1( u1_u1_u5_n105 ) , .ZN( u1_u1_u5_n140 ) );
  NAND2_X1 u1_u1_u5_U63 (.A2( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n105 ) , .ZN( u1_u1_u5_n155 ) );
  NAND2_X1 u1_u1_u5_U64 (.A2( u1_u1_u5_n106 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n122 ) );
  NAND2_X1 u1_u1_u5_U65 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n106 ) , .ZN( u1_u1_u5_n115 ) );
  NAND2_X1 u1_u1_u5_U66 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n103 ) , .ZN( u1_u1_u5_n161 ) );
  NAND2_X1 u1_u1_u5_U67 (.A1( u1_u1_u5_n105 ) , .A2( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n154 ) );
  INV_X1 u1_u1_u5_U68 (.A( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n172 ) );
  NAND2_X1 u1_u1_u5_U69 (.A1( u1_u1_u5_n103 ) , .A2( u1_u1_u5_n108 ) , .ZN( u1_u1_u5_n123 ) );
  OAI22_X1 u1_u1_u5_U7 (.B2( u1_u1_u5_n149 ) , .B1( u1_u1_u5_n150 ) , .A2( u1_u1_u5_n151 ) , .A1( u1_u1_u5_n152 ) , .ZN( u1_u1_u5_n165 ) );
  NAND2_X1 u1_u1_u5_U70 (.A2( u1_u1_u5_n103 ) , .A1( u1_u1_u5_n107 ) , .ZN( u1_u1_u5_n151 ) );
  NAND2_X1 u1_u1_u5_U71 (.A2( u1_u1_u5_n107 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n120 ) );
  NAND2_X1 u1_u1_u5_U72 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n109 ) , .ZN( u1_u1_u5_n157 ) );
  AND2_X1 u1_u1_u5_U73 (.A2( u1_u1_u5_n100 ) , .A1( u1_u1_u5_n104 ) , .ZN( u1_u1_u5_n131 ) );
  INV_X1 u1_u1_u5_U74 (.A( u1_u1_u5_n102 ) , .ZN( u1_u1_u5_n195 ) );
  OAI221_X1 u1_u1_u5_U75 (.A( u1_u1_u5_n101 ) , .ZN( u1_u1_u5_n102 ) , .C2( u1_u1_u5_n115 ) , .C1( u1_u1_u5_n126 ) , .B1( u1_u1_u5_n134 ) , .B2( u1_u1_u5_n160 ) );
  OAI21_X1 u1_u1_u5_U76 (.ZN( u1_u1_u5_n101 ) , .B1( u1_u1_u5_n137 ) , .A( u1_u1_u5_n146 ) , .B2( u1_u1_u5_n147 ) );
  NOR2_X1 u1_u1_u5_U77 (.A2( u1_u1_X_34 ) , .A1( u1_u1_X_35 ) , .ZN( u1_u1_u5_n145 ) );
  NOR2_X1 u1_u1_u5_U78 (.A2( u1_u1_X_34 ) , .ZN( u1_u1_u5_n146 ) , .A1( u1_u1_u5_n171 ) );
  NOR2_X1 u1_u1_u5_U79 (.A2( u1_u1_X_31 ) , .A1( u1_u1_X_32 ) , .ZN( u1_u1_u5_n103 ) );
  NOR3_X1 u1_u1_u5_U8 (.A2( u1_u1_u5_n147 ) , .A1( u1_u1_u5_n148 ) , .ZN( u1_u1_u5_n149 ) , .A3( u1_u1_u5_n194 ) );
  NOR2_X1 u1_u1_u5_U80 (.A2( u1_u1_X_36 ) , .ZN( u1_u1_u5_n105 ) , .A1( u1_u1_u5_n180 ) );
  NOR2_X1 u1_u1_u5_U81 (.A2( u1_u1_X_33 ) , .ZN( u1_u1_u5_n108 ) , .A1( u1_u1_u5_n170 ) );
  NOR2_X1 u1_u1_u5_U82 (.A2( u1_u1_X_33 ) , .A1( u1_u1_X_36 ) , .ZN( u1_u1_u5_n107 ) );
  NOR2_X1 u1_u1_u5_U83 (.A2( u1_u1_X_31 ) , .ZN( u1_u1_u5_n104 ) , .A1( u1_u1_u5_n181 ) );
  NAND2_X1 u1_u1_u5_U84 (.A2( u1_u1_X_34 ) , .A1( u1_u1_X_35 ) , .ZN( u1_u1_u5_n153 ) );
  NAND2_X1 u1_u1_u5_U85 (.A1( u1_u1_X_34 ) , .ZN( u1_u1_u5_n126 ) , .A2( u1_u1_u5_n171 ) );
  AND2_X1 u1_u1_u5_U86 (.A1( u1_u1_X_31 ) , .A2( u1_u1_X_32 ) , .ZN( u1_u1_u5_n106 ) );
  AND2_X1 u1_u1_u5_U87 (.A1( u1_u1_X_31 ) , .ZN( u1_u1_u5_n109 ) , .A2( u1_u1_u5_n181 ) );
  INV_X1 u1_u1_u5_U88 (.A( u1_u1_X_33 ) , .ZN( u1_u1_u5_n180 ) );
  INV_X1 u1_u1_u5_U89 (.A( u1_u1_X_35 ) , .ZN( u1_u1_u5_n171 ) );
  NOR2_X1 u1_u1_u5_U9 (.ZN( u1_u1_u5_n135 ) , .A1( u1_u1_u5_n173 ) , .A2( u1_u1_u5_n176 ) );
  INV_X1 u1_u1_u5_U90 (.A( u1_u1_X_36 ) , .ZN( u1_u1_u5_n170 ) );
  INV_X1 u1_u1_u5_U91 (.A( u1_u1_X_32 ) , .ZN( u1_u1_u5_n181 ) );
  NAND4_X1 u1_u1_u5_U92 (.ZN( u1_out1_29 ) , .A4( u1_u1_u5_n129 ) , .A3( u1_u1_u5_n130 ) , .A2( u1_u1_u5_n168 ) , .A1( u1_u1_u5_n196 ) );
  AOI221_X1 u1_u1_u5_U93 (.A( u1_u1_u5_n128 ) , .ZN( u1_u1_u5_n129 ) , .C2( u1_u1_u5_n132 ) , .B2( u1_u1_u5_n159 ) , .B1( u1_u1_u5_n176 ) , .C1( u1_u1_u5_n184 ) );
  AOI222_X1 u1_u1_u5_U94 (.ZN( u1_u1_u5_n130 ) , .A2( u1_u1_u5_n146 ) , .B1( u1_u1_u5_n147 ) , .C2( u1_u1_u5_n175 ) , .B2( u1_u1_u5_n179 ) , .A1( u1_u1_u5_n188 ) , .C1( u1_u1_u5_n194 ) );
  NAND4_X1 u1_u1_u5_U95 (.ZN( u1_out1_19 ) , .A4( u1_u1_u5_n166 ) , .A3( u1_u1_u5_n167 ) , .A2( u1_u1_u5_n168 ) , .A1( u1_u1_u5_n169 ) );
  AOI22_X1 u1_u1_u5_U96 (.B2( u1_u1_u5_n145 ) , .A2( u1_u1_u5_n146 ) , .ZN( u1_u1_u5_n167 ) , .B1( u1_u1_u5_n182 ) , .A1( u1_u1_u5_n189 ) );
  NOR4_X1 u1_u1_u5_U97 (.A4( u1_u1_u5_n162 ) , .A3( u1_u1_u5_n163 ) , .A2( u1_u1_u5_n164 ) , .A1( u1_u1_u5_n165 ) , .ZN( u1_u1_u5_n166 ) );
  NAND4_X1 u1_u1_u5_U98 (.ZN( u1_out1_11 ) , .A4( u1_u1_u5_n143 ) , .A3( u1_u1_u5_n144 ) , .A2( u1_u1_u5_n169 ) , .A1( u1_u1_u5_n196 ) );
  AOI22_X1 u1_u1_u5_U99 (.A2( u1_u1_u5_n132 ) , .ZN( u1_u1_u5_n144 ) , .B2( u1_u1_u5_n145 ) , .B1( u1_u1_u5_n184 ) , .A1( u1_u1_u5_n194 ) );
  XOR2_X1 u1_u2_U20 (.B( u1_K3_36 ) , .A( u1_R1_25 ) , .Z( u1_u2_X_36 ) );
  XOR2_X1 u1_u2_U21 (.B( u1_K3_35 ) , .A( u1_R1_24 ) , .Z( u1_u2_X_35 ) );
  XOR2_X1 u1_u2_U22 (.B( u1_K3_34 ) , .A( u1_R1_23 ) , .Z( u1_u2_X_34 ) );
  XOR2_X1 u1_u2_U23 (.B( u1_K3_33 ) , .A( u1_R1_22 ) , .Z( u1_u2_X_33 ) );
  XOR2_X1 u1_u2_U24 (.B( u1_K3_32 ) , .A( u1_R1_21 ) , .Z( u1_u2_X_32 ) );
  XOR2_X1 u1_u2_U25 (.B( u1_K3_31 ) , .A( u1_R1_20 ) , .Z( u1_u2_X_31 ) );
  XOR2_X1 u1_u2_U26 (.B( u1_K3_30 ) , .A( u1_R1_21 ) , .Z( u1_u2_X_30 ) );
  XOR2_X1 u1_u2_U28 (.B( u1_K3_29 ) , .A( u1_R1_20 ) , .Z( u1_u2_X_29 ) );
  XOR2_X1 u1_u2_U29 (.B( u1_K3_28 ) , .A( u1_R1_19 ) , .Z( u1_u2_X_28 ) );
  XOR2_X1 u1_u2_U30 (.B( u1_K3_27 ) , .A( u1_R1_18 ) , .Z( u1_u2_X_27 ) );
  XOR2_X1 u1_u2_U31 (.B( u1_K3_26 ) , .A( u1_R1_17 ) , .Z( u1_u2_X_26 ) );
  XOR2_X1 u1_u2_U32 (.B( u1_K3_25 ) , .A( u1_R1_16 ) , .Z( u1_u2_X_25 ) );
  OAI22_X1 u1_u2_u4_U10 (.B2( u1_u2_u4_n135 ) , .ZN( u1_u2_u4_n137 ) , .B1( u1_u2_u4_n153 ) , .A1( u1_u2_u4_n155 ) , .A2( u1_u2_u4_n171 ) );
  AND3_X1 u1_u2_u4_U11 (.A2( u1_u2_u4_n134 ) , .ZN( u1_u2_u4_n135 ) , .A3( u1_u2_u4_n145 ) , .A1( u1_u2_u4_n157 ) );
  NAND2_X1 u1_u2_u4_U12 (.ZN( u1_u2_u4_n132 ) , .A2( u1_u2_u4_n170 ) , .A1( u1_u2_u4_n173 ) );
  AOI21_X1 u1_u2_u4_U13 (.B2( u1_u2_u4_n160 ) , .B1( u1_u2_u4_n161 ) , .ZN( u1_u2_u4_n162 ) , .A( u1_u2_u4_n170 ) );
  AOI21_X1 u1_u2_u4_U14 (.ZN( u1_u2_u4_n107 ) , .B2( u1_u2_u4_n143 ) , .A( u1_u2_u4_n174 ) , .B1( u1_u2_u4_n184 ) );
  AOI21_X1 u1_u2_u4_U15 (.B2( u1_u2_u4_n158 ) , .B1( u1_u2_u4_n159 ) , .ZN( u1_u2_u4_n163 ) , .A( u1_u2_u4_n174 ) );
  AOI21_X1 u1_u2_u4_U16 (.A( u1_u2_u4_n153 ) , .B2( u1_u2_u4_n154 ) , .B1( u1_u2_u4_n155 ) , .ZN( u1_u2_u4_n165 ) );
  AOI21_X1 u1_u2_u4_U17 (.A( u1_u2_u4_n156 ) , .B2( u1_u2_u4_n157 ) , .ZN( u1_u2_u4_n164 ) , .B1( u1_u2_u4_n184 ) );
  INV_X1 u1_u2_u4_U18 (.A( u1_u2_u4_n138 ) , .ZN( u1_u2_u4_n170 ) );
  AND2_X1 u1_u2_u4_U19 (.A2( u1_u2_u4_n120 ) , .ZN( u1_u2_u4_n155 ) , .A1( u1_u2_u4_n160 ) );
  INV_X1 u1_u2_u4_U20 (.A( u1_u2_u4_n156 ) , .ZN( u1_u2_u4_n175 ) );
  NAND2_X1 u1_u2_u4_U21 (.A2( u1_u2_u4_n118 ) , .ZN( u1_u2_u4_n131 ) , .A1( u1_u2_u4_n147 ) );
  NAND2_X1 u1_u2_u4_U22 (.A1( u1_u2_u4_n119 ) , .A2( u1_u2_u4_n120 ) , .ZN( u1_u2_u4_n130 ) );
  NAND2_X1 u1_u2_u4_U23 (.ZN( u1_u2_u4_n117 ) , .A2( u1_u2_u4_n118 ) , .A1( u1_u2_u4_n148 ) );
  NAND2_X1 u1_u2_u4_U24 (.ZN( u1_u2_u4_n129 ) , .A1( u1_u2_u4_n134 ) , .A2( u1_u2_u4_n148 ) );
  AND3_X1 u1_u2_u4_U25 (.A1( u1_u2_u4_n119 ) , .A2( u1_u2_u4_n143 ) , .A3( u1_u2_u4_n154 ) , .ZN( u1_u2_u4_n161 ) );
  AND2_X1 u1_u2_u4_U26 (.A1( u1_u2_u4_n145 ) , .A2( u1_u2_u4_n147 ) , .ZN( u1_u2_u4_n159 ) );
  OR3_X1 u1_u2_u4_U27 (.A3( u1_u2_u4_n114 ) , .A2( u1_u2_u4_n115 ) , .A1( u1_u2_u4_n116 ) , .ZN( u1_u2_u4_n136 ) );
  AOI21_X1 u1_u2_u4_U28 (.A( u1_u2_u4_n113 ) , .ZN( u1_u2_u4_n116 ) , .B2( u1_u2_u4_n173 ) , .B1( u1_u2_u4_n174 ) );
  AOI21_X1 u1_u2_u4_U29 (.ZN( u1_u2_u4_n115 ) , .B2( u1_u2_u4_n145 ) , .B1( u1_u2_u4_n146 ) , .A( u1_u2_u4_n156 ) );
  NOR2_X1 u1_u2_u4_U3 (.ZN( u1_u2_u4_n121 ) , .A1( u1_u2_u4_n181 ) , .A2( u1_u2_u4_n182 ) );
  OAI22_X1 u1_u2_u4_U30 (.ZN( u1_u2_u4_n114 ) , .A2( u1_u2_u4_n121 ) , .B1( u1_u2_u4_n160 ) , .B2( u1_u2_u4_n170 ) , .A1( u1_u2_u4_n171 ) );
  INV_X1 u1_u2_u4_U31 (.A( u1_u2_u4_n158 ) , .ZN( u1_u2_u4_n182 ) );
  INV_X1 u1_u2_u4_U32 (.ZN( u1_u2_u4_n181 ) , .A( u1_u2_u4_n96 ) );
  INV_X1 u1_u2_u4_U33 (.A( u1_u2_u4_n144 ) , .ZN( u1_u2_u4_n179 ) );
  INV_X1 u1_u2_u4_U34 (.A( u1_u2_u4_n157 ) , .ZN( u1_u2_u4_n178 ) );
  NAND2_X1 u1_u2_u4_U35 (.A2( u1_u2_u4_n154 ) , .A1( u1_u2_u4_n96 ) , .ZN( u1_u2_u4_n97 ) );
  INV_X1 u1_u2_u4_U36 (.ZN( u1_u2_u4_n186 ) , .A( u1_u2_u4_n95 ) );
  OAI221_X1 u1_u2_u4_U37 (.C1( u1_u2_u4_n134 ) , .B1( u1_u2_u4_n158 ) , .B2( u1_u2_u4_n171 ) , .C2( u1_u2_u4_n173 ) , .A( u1_u2_u4_n94 ) , .ZN( u1_u2_u4_n95 ) );
  AOI222_X1 u1_u2_u4_U38 (.B2( u1_u2_u4_n132 ) , .A1( u1_u2_u4_n138 ) , .C2( u1_u2_u4_n175 ) , .A2( u1_u2_u4_n179 ) , .C1( u1_u2_u4_n181 ) , .B1( u1_u2_u4_n185 ) , .ZN( u1_u2_u4_n94 ) );
  INV_X1 u1_u2_u4_U39 (.A( u1_u2_u4_n113 ) , .ZN( u1_u2_u4_n185 ) );
  INV_X1 u1_u2_u4_U4 (.A( u1_u2_u4_n117 ) , .ZN( u1_u2_u4_n184 ) );
  INV_X1 u1_u2_u4_U40 (.A( u1_u2_u4_n143 ) , .ZN( u1_u2_u4_n183 ) );
  NOR2_X1 u1_u2_u4_U41 (.ZN( u1_u2_u4_n138 ) , .A1( u1_u2_u4_n168 ) , .A2( u1_u2_u4_n169 ) );
  NOR2_X1 u1_u2_u4_U42 (.A1( u1_u2_u4_n150 ) , .A2( u1_u2_u4_n152 ) , .ZN( u1_u2_u4_n153 ) );
  NOR2_X1 u1_u2_u4_U43 (.A2( u1_u2_u4_n128 ) , .A1( u1_u2_u4_n138 ) , .ZN( u1_u2_u4_n156 ) );
  AOI22_X1 u1_u2_u4_U44 (.B2( u1_u2_u4_n122 ) , .A1( u1_u2_u4_n123 ) , .ZN( u1_u2_u4_n124 ) , .B1( u1_u2_u4_n128 ) , .A2( u1_u2_u4_n172 ) );
  INV_X1 u1_u2_u4_U45 (.A( u1_u2_u4_n153 ) , .ZN( u1_u2_u4_n172 ) );
  NAND2_X1 u1_u2_u4_U46 (.A2( u1_u2_u4_n120 ) , .ZN( u1_u2_u4_n123 ) , .A1( u1_u2_u4_n161 ) );
  AOI22_X1 u1_u2_u4_U47 (.B2( u1_u2_u4_n132 ) , .A2( u1_u2_u4_n133 ) , .ZN( u1_u2_u4_n140 ) , .A1( u1_u2_u4_n150 ) , .B1( u1_u2_u4_n179 ) );
  NAND2_X1 u1_u2_u4_U48 (.ZN( u1_u2_u4_n133 ) , .A2( u1_u2_u4_n146 ) , .A1( u1_u2_u4_n154 ) );
  NAND2_X1 u1_u2_u4_U49 (.A1( u1_u2_u4_n103 ) , .ZN( u1_u2_u4_n154 ) , .A2( u1_u2_u4_n98 ) );
  NOR4_X1 u1_u2_u4_U5 (.A4( u1_u2_u4_n106 ) , .A3( u1_u2_u4_n107 ) , .A2( u1_u2_u4_n108 ) , .A1( u1_u2_u4_n109 ) , .ZN( u1_u2_u4_n110 ) );
  NAND2_X1 u1_u2_u4_U50 (.A1( u1_u2_u4_n101 ) , .ZN( u1_u2_u4_n158 ) , .A2( u1_u2_u4_n99 ) );
  AOI21_X1 u1_u2_u4_U51 (.ZN( u1_u2_u4_n127 ) , .A( u1_u2_u4_n136 ) , .B2( u1_u2_u4_n150 ) , .B1( u1_u2_u4_n180 ) );
  INV_X1 u1_u2_u4_U52 (.A( u1_u2_u4_n160 ) , .ZN( u1_u2_u4_n180 ) );
  NAND2_X1 u1_u2_u4_U53 (.A2( u1_u2_u4_n104 ) , .A1( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n146 ) );
  NAND2_X1 u1_u2_u4_U54 (.A2( u1_u2_u4_n101 ) , .A1( u1_u2_u4_n102 ) , .ZN( u1_u2_u4_n160 ) );
  NAND2_X1 u1_u2_u4_U55 (.ZN( u1_u2_u4_n134 ) , .A1( u1_u2_u4_n98 ) , .A2( u1_u2_u4_n99 ) );
  NAND2_X1 u1_u2_u4_U56 (.A1( u1_u2_u4_n103 ) , .A2( u1_u2_u4_n104 ) , .ZN( u1_u2_u4_n143 ) );
  NAND2_X1 u1_u2_u4_U57 (.A2( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n145 ) , .A1( u1_u2_u4_n98 ) );
  NAND2_X1 u1_u2_u4_U58 (.A1( u1_u2_u4_n100 ) , .A2( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n120 ) );
  NAND2_X1 u1_u2_u4_U59 (.A1( u1_u2_u4_n102 ) , .A2( u1_u2_u4_n104 ) , .ZN( u1_u2_u4_n148 ) );
  AOI21_X1 u1_u2_u4_U6 (.ZN( u1_u2_u4_n106 ) , .B2( u1_u2_u4_n146 ) , .B1( u1_u2_u4_n158 ) , .A( u1_u2_u4_n170 ) );
  NAND2_X1 u1_u2_u4_U60 (.A2( u1_u2_u4_n100 ) , .A1( u1_u2_u4_n103 ) , .ZN( u1_u2_u4_n157 ) );
  INV_X1 u1_u2_u4_U61 (.A( u1_u2_u4_n150 ) , .ZN( u1_u2_u4_n173 ) );
  INV_X1 u1_u2_u4_U62 (.A( u1_u2_u4_n152 ) , .ZN( u1_u2_u4_n171 ) );
  NAND2_X1 u1_u2_u4_U63 (.A1( u1_u2_u4_n100 ) , .ZN( u1_u2_u4_n118 ) , .A2( u1_u2_u4_n99 ) );
  NAND2_X1 u1_u2_u4_U64 (.A2( u1_u2_u4_n100 ) , .A1( u1_u2_u4_n102 ) , .ZN( u1_u2_u4_n144 ) );
  NAND2_X1 u1_u2_u4_U65 (.A2( u1_u2_u4_n101 ) , .A1( u1_u2_u4_n105 ) , .ZN( u1_u2_u4_n96 ) );
  INV_X1 u1_u2_u4_U66 (.A( u1_u2_u4_n128 ) , .ZN( u1_u2_u4_n174 ) );
  NAND2_X1 u1_u2_u4_U67 (.A2( u1_u2_u4_n102 ) , .ZN( u1_u2_u4_n119 ) , .A1( u1_u2_u4_n98 ) );
  NAND2_X1 u1_u2_u4_U68 (.A2( u1_u2_u4_n101 ) , .A1( u1_u2_u4_n103 ) , .ZN( u1_u2_u4_n147 ) );
  NAND2_X1 u1_u2_u4_U69 (.A2( u1_u2_u4_n104 ) , .ZN( u1_u2_u4_n113 ) , .A1( u1_u2_u4_n99 ) );
  AOI21_X1 u1_u2_u4_U7 (.ZN( u1_u2_u4_n108 ) , .B2( u1_u2_u4_n134 ) , .B1( u1_u2_u4_n155 ) , .A( u1_u2_u4_n156 ) );
  NOR2_X1 u1_u2_u4_U70 (.A2( u1_u2_X_28 ) , .ZN( u1_u2_u4_n150 ) , .A1( u1_u2_u4_n168 ) );
  NOR2_X1 u1_u2_u4_U71 (.A2( u1_u2_X_29 ) , .ZN( u1_u2_u4_n152 ) , .A1( u1_u2_u4_n169 ) );
  NOR2_X1 u1_u2_u4_U72 (.A2( u1_u2_X_30 ) , .ZN( u1_u2_u4_n105 ) , .A1( u1_u2_u4_n176 ) );
  NOR2_X1 u1_u2_u4_U73 (.A2( u1_u2_X_26 ) , .ZN( u1_u2_u4_n100 ) , .A1( u1_u2_u4_n177 ) );
  NOR2_X1 u1_u2_u4_U74 (.A2( u1_u2_X_28 ) , .A1( u1_u2_X_29 ) , .ZN( u1_u2_u4_n128 ) );
  NOR2_X1 u1_u2_u4_U75 (.A2( u1_u2_X_27 ) , .A1( u1_u2_X_30 ) , .ZN( u1_u2_u4_n102 ) );
  NOR2_X1 u1_u2_u4_U76 (.A2( u1_u2_X_25 ) , .A1( u1_u2_X_26 ) , .ZN( u1_u2_u4_n98 ) );
  AND2_X1 u1_u2_u4_U77 (.A2( u1_u2_X_25 ) , .A1( u1_u2_X_26 ) , .ZN( u1_u2_u4_n104 ) );
  AND2_X1 u1_u2_u4_U78 (.A1( u1_u2_X_30 ) , .A2( u1_u2_u4_n176 ) , .ZN( u1_u2_u4_n99 ) );
  AND2_X1 u1_u2_u4_U79 (.A1( u1_u2_X_26 ) , .ZN( u1_u2_u4_n101 ) , .A2( u1_u2_u4_n177 ) );
  AOI21_X1 u1_u2_u4_U8 (.ZN( u1_u2_u4_n109 ) , .A( u1_u2_u4_n153 ) , .B1( u1_u2_u4_n159 ) , .B2( u1_u2_u4_n184 ) );
  AND2_X1 u1_u2_u4_U80 (.A1( u1_u2_X_27 ) , .A2( u1_u2_X_30 ) , .ZN( u1_u2_u4_n103 ) );
  INV_X1 u1_u2_u4_U81 (.A( u1_u2_X_28 ) , .ZN( u1_u2_u4_n169 ) );
  INV_X1 u1_u2_u4_U82 (.A( u1_u2_X_29 ) , .ZN( u1_u2_u4_n168 ) );
  INV_X1 u1_u2_u4_U83 (.A( u1_u2_X_25 ) , .ZN( u1_u2_u4_n177 ) );
  INV_X1 u1_u2_u4_U84 (.A( u1_u2_X_27 ) , .ZN( u1_u2_u4_n176 ) );
  NAND4_X1 u1_u2_u4_U85 (.ZN( u1_out2_25 ) , .A4( u1_u2_u4_n139 ) , .A3( u1_u2_u4_n140 ) , .A2( u1_u2_u4_n141 ) , .A1( u1_u2_u4_n142 ) );
  OAI21_X1 u1_u2_u4_U86 (.A( u1_u2_u4_n128 ) , .B2( u1_u2_u4_n129 ) , .B1( u1_u2_u4_n130 ) , .ZN( u1_u2_u4_n142 ) );
  OAI21_X1 u1_u2_u4_U87 (.B2( u1_u2_u4_n131 ) , .ZN( u1_u2_u4_n141 ) , .A( u1_u2_u4_n175 ) , .B1( u1_u2_u4_n183 ) );
  NAND4_X1 u1_u2_u4_U88 (.ZN( u1_out2_14 ) , .A4( u1_u2_u4_n124 ) , .A3( u1_u2_u4_n125 ) , .A2( u1_u2_u4_n126 ) , .A1( u1_u2_u4_n127 ) );
  AOI22_X1 u1_u2_u4_U89 (.B2( u1_u2_u4_n117 ) , .ZN( u1_u2_u4_n126 ) , .A1( u1_u2_u4_n129 ) , .B1( u1_u2_u4_n152 ) , .A2( u1_u2_u4_n175 ) );
  AOI211_X1 u1_u2_u4_U9 (.B( u1_u2_u4_n136 ) , .A( u1_u2_u4_n137 ) , .C2( u1_u2_u4_n138 ) , .ZN( u1_u2_u4_n139 ) , .C1( u1_u2_u4_n182 ) );
  AOI22_X1 u1_u2_u4_U90 (.ZN( u1_u2_u4_n125 ) , .B2( u1_u2_u4_n131 ) , .A2( u1_u2_u4_n132 ) , .B1( u1_u2_u4_n138 ) , .A1( u1_u2_u4_n178 ) );
  NAND4_X1 u1_u2_u4_U91 (.ZN( u1_out2_8 ) , .A4( u1_u2_u4_n110 ) , .A3( u1_u2_u4_n111 ) , .A2( u1_u2_u4_n112 ) , .A1( u1_u2_u4_n186 ) );
  NAND2_X1 u1_u2_u4_U92 (.ZN( u1_u2_u4_n112 ) , .A2( u1_u2_u4_n130 ) , .A1( u1_u2_u4_n150 ) );
  AOI22_X1 u1_u2_u4_U93 (.ZN( u1_u2_u4_n111 ) , .B2( u1_u2_u4_n132 ) , .A1( u1_u2_u4_n152 ) , .B1( u1_u2_u4_n178 ) , .A2( u1_u2_u4_n97 ) );
  AOI22_X1 u1_u2_u4_U94 (.B2( u1_u2_u4_n149 ) , .B1( u1_u2_u4_n150 ) , .A2( u1_u2_u4_n151 ) , .A1( u1_u2_u4_n152 ) , .ZN( u1_u2_u4_n167 ) );
  NOR4_X1 u1_u2_u4_U95 (.A4( u1_u2_u4_n162 ) , .A3( u1_u2_u4_n163 ) , .A2( u1_u2_u4_n164 ) , .A1( u1_u2_u4_n165 ) , .ZN( u1_u2_u4_n166 ) );
  NAND3_X1 u1_u2_u4_U96 (.ZN( u1_out2_3 ) , .A3( u1_u2_u4_n166 ) , .A1( u1_u2_u4_n167 ) , .A2( u1_u2_u4_n186 ) );
  NAND3_X1 u1_u2_u4_U97 (.A3( u1_u2_u4_n146 ) , .A2( u1_u2_u4_n147 ) , .A1( u1_u2_u4_n148 ) , .ZN( u1_u2_u4_n149 ) );
  NAND3_X1 u1_u2_u4_U98 (.A3( u1_u2_u4_n143 ) , .A2( u1_u2_u4_n144 ) , .A1( u1_u2_u4_n145 ) , .ZN( u1_u2_u4_n151 ) );
  NAND3_X1 u1_u2_u4_U99 (.A3( u1_u2_u4_n121 ) , .ZN( u1_u2_u4_n122 ) , .A2( u1_u2_u4_n144 ) , .A1( u1_u2_u4_n154 ) );
  INV_X1 u1_u2_u5_U10 (.A( u1_u2_u5_n121 ) , .ZN( u1_u2_u5_n177 ) );
  NOR3_X1 u1_u2_u5_U100 (.A3( u1_u2_u5_n141 ) , .A1( u1_u2_u5_n142 ) , .ZN( u1_u2_u5_n143 ) , .A2( u1_u2_u5_n191 ) );
  NAND4_X1 u1_u2_u5_U101 (.ZN( u1_out2_4 ) , .A4( u1_u2_u5_n112 ) , .A2( u1_u2_u5_n113 ) , .A1( u1_u2_u5_n114 ) , .A3( u1_u2_u5_n195 ) );
  AOI211_X1 u1_u2_u5_U102 (.A( u1_u2_u5_n110 ) , .C1( u1_u2_u5_n111 ) , .ZN( u1_u2_u5_n112 ) , .B( u1_u2_u5_n118 ) , .C2( u1_u2_u5_n177 ) );
  AOI222_X1 u1_u2_u5_U103 (.ZN( u1_u2_u5_n113 ) , .A1( u1_u2_u5_n131 ) , .C1( u1_u2_u5_n148 ) , .B2( u1_u2_u5_n174 ) , .C2( u1_u2_u5_n178 ) , .A2( u1_u2_u5_n179 ) , .B1( u1_u2_u5_n99 ) );
  NAND3_X1 u1_u2_u5_U104 (.A2( u1_u2_u5_n154 ) , .A3( u1_u2_u5_n158 ) , .A1( u1_u2_u5_n161 ) , .ZN( u1_u2_u5_n99 ) );
  NOR2_X1 u1_u2_u5_U11 (.ZN( u1_u2_u5_n160 ) , .A2( u1_u2_u5_n173 ) , .A1( u1_u2_u5_n177 ) );
  INV_X1 u1_u2_u5_U12 (.A( u1_u2_u5_n150 ) , .ZN( u1_u2_u5_n174 ) );
  AOI21_X1 u1_u2_u5_U13 (.A( u1_u2_u5_n160 ) , .B2( u1_u2_u5_n161 ) , .ZN( u1_u2_u5_n162 ) , .B1( u1_u2_u5_n192 ) );
  INV_X1 u1_u2_u5_U14 (.A( u1_u2_u5_n159 ) , .ZN( u1_u2_u5_n192 ) );
  AOI21_X1 u1_u2_u5_U15 (.A( u1_u2_u5_n156 ) , .B2( u1_u2_u5_n157 ) , .B1( u1_u2_u5_n158 ) , .ZN( u1_u2_u5_n163 ) );
  AOI21_X1 u1_u2_u5_U16 (.B2( u1_u2_u5_n139 ) , .B1( u1_u2_u5_n140 ) , .ZN( u1_u2_u5_n141 ) , .A( u1_u2_u5_n150 ) );
  OAI21_X1 u1_u2_u5_U17 (.A( u1_u2_u5_n133 ) , .B2( u1_u2_u5_n134 ) , .B1( u1_u2_u5_n135 ) , .ZN( u1_u2_u5_n142 ) );
  OAI21_X1 u1_u2_u5_U18 (.ZN( u1_u2_u5_n133 ) , .B2( u1_u2_u5_n147 ) , .A( u1_u2_u5_n173 ) , .B1( u1_u2_u5_n188 ) );
  NAND2_X1 u1_u2_u5_U19 (.A2( u1_u2_u5_n119 ) , .A1( u1_u2_u5_n123 ) , .ZN( u1_u2_u5_n137 ) );
  INV_X1 u1_u2_u5_U20 (.A( u1_u2_u5_n155 ) , .ZN( u1_u2_u5_n194 ) );
  NAND2_X1 u1_u2_u5_U21 (.A1( u1_u2_u5_n121 ) , .ZN( u1_u2_u5_n132 ) , .A2( u1_u2_u5_n172 ) );
  NAND2_X1 u1_u2_u5_U22 (.A2( u1_u2_u5_n122 ) , .ZN( u1_u2_u5_n136 ) , .A1( u1_u2_u5_n154 ) );
  NAND2_X1 u1_u2_u5_U23 (.A2( u1_u2_u5_n119 ) , .A1( u1_u2_u5_n120 ) , .ZN( u1_u2_u5_n159 ) );
  INV_X1 u1_u2_u5_U24 (.A( u1_u2_u5_n156 ) , .ZN( u1_u2_u5_n175 ) );
  INV_X1 u1_u2_u5_U25 (.A( u1_u2_u5_n158 ) , .ZN( u1_u2_u5_n188 ) );
  INV_X1 u1_u2_u5_U26 (.A( u1_u2_u5_n152 ) , .ZN( u1_u2_u5_n179 ) );
  INV_X1 u1_u2_u5_U27 (.A( u1_u2_u5_n140 ) , .ZN( u1_u2_u5_n182 ) );
  INV_X1 u1_u2_u5_U28 (.A( u1_u2_u5_n151 ) , .ZN( u1_u2_u5_n183 ) );
  INV_X1 u1_u2_u5_U29 (.A( u1_u2_u5_n123 ) , .ZN( u1_u2_u5_n185 ) );
  NOR2_X1 u1_u2_u5_U3 (.ZN( u1_u2_u5_n134 ) , .A1( u1_u2_u5_n183 ) , .A2( u1_u2_u5_n190 ) );
  INV_X1 u1_u2_u5_U30 (.A( u1_u2_u5_n161 ) , .ZN( u1_u2_u5_n184 ) );
  INV_X1 u1_u2_u5_U31 (.A( u1_u2_u5_n139 ) , .ZN( u1_u2_u5_n189 ) );
  INV_X1 u1_u2_u5_U32 (.A( u1_u2_u5_n157 ) , .ZN( u1_u2_u5_n190 ) );
  INV_X1 u1_u2_u5_U33 (.A( u1_u2_u5_n120 ) , .ZN( u1_u2_u5_n193 ) );
  NAND2_X1 u1_u2_u5_U34 (.ZN( u1_u2_u5_n111 ) , .A1( u1_u2_u5_n140 ) , .A2( u1_u2_u5_n155 ) );
  INV_X1 u1_u2_u5_U35 (.A( u1_u2_u5_n117 ) , .ZN( u1_u2_u5_n196 ) );
  OAI221_X1 u1_u2_u5_U36 (.A( u1_u2_u5_n116 ) , .ZN( u1_u2_u5_n117 ) , .B2( u1_u2_u5_n119 ) , .C1( u1_u2_u5_n153 ) , .C2( u1_u2_u5_n158 ) , .B1( u1_u2_u5_n172 ) );
  AOI222_X1 u1_u2_u5_U37 (.ZN( u1_u2_u5_n116 ) , .B2( u1_u2_u5_n145 ) , .C1( u1_u2_u5_n148 ) , .A2( u1_u2_u5_n174 ) , .C2( u1_u2_u5_n177 ) , .B1( u1_u2_u5_n187 ) , .A1( u1_u2_u5_n193 ) );
  INV_X1 u1_u2_u5_U38 (.A( u1_u2_u5_n115 ) , .ZN( u1_u2_u5_n187 ) );
  NOR2_X1 u1_u2_u5_U39 (.ZN( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n170 ) , .A2( u1_u2_u5_n180 ) );
  INV_X1 u1_u2_u5_U4 (.A( u1_u2_u5_n138 ) , .ZN( u1_u2_u5_n191 ) );
  AOI22_X1 u1_u2_u5_U40 (.B2( u1_u2_u5_n131 ) , .A2( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n169 ) , .B1( u1_u2_u5_n174 ) , .A1( u1_u2_u5_n185 ) );
  NOR2_X1 u1_u2_u5_U41 (.A1( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n150 ) , .A2( u1_u2_u5_n173 ) );
  AOI21_X1 u1_u2_u5_U42 (.A( u1_u2_u5_n118 ) , .B2( u1_u2_u5_n145 ) , .ZN( u1_u2_u5_n168 ) , .B1( u1_u2_u5_n186 ) );
  INV_X1 u1_u2_u5_U43 (.A( u1_u2_u5_n122 ) , .ZN( u1_u2_u5_n186 ) );
  NOR2_X1 u1_u2_u5_U44 (.A1( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n152 ) , .A2( u1_u2_u5_n176 ) );
  NOR2_X1 u1_u2_u5_U45 (.A1( u1_u2_u5_n115 ) , .ZN( u1_u2_u5_n118 ) , .A2( u1_u2_u5_n153 ) );
  NOR2_X1 u1_u2_u5_U46 (.A2( u1_u2_u5_n145 ) , .ZN( u1_u2_u5_n156 ) , .A1( u1_u2_u5_n174 ) );
  NOR2_X1 u1_u2_u5_U47 (.ZN( u1_u2_u5_n121 ) , .A2( u1_u2_u5_n145 ) , .A1( u1_u2_u5_n176 ) );
  AOI22_X1 u1_u2_u5_U48 (.ZN( u1_u2_u5_n114 ) , .A2( u1_u2_u5_n137 ) , .A1( u1_u2_u5_n145 ) , .B2( u1_u2_u5_n175 ) , .B1( u1_u2_u5_n193 ) );
  OAI211_X1 u1_u2_u5_U49 (.B( u1_u2_u5_n124 ) , .A( u1_u2_u5_n125 ) , .C2( u1_u2_u5_n126 ) , .C1( u1_u2_u5_n127 ) , .ZN( u1_u2_u5_n128 ) );
  OAI21_X1 u1_u2_u5_U5 (.B2( u1_u2_u5_n136 ) , .B1( u1_u2_u5_n137 ) , .ZN( u1_u2_u5_n138 ) , .A( u1_u2_u5_n177 ) );
  NOR3_X1 u1_u2_u5_U50 (.ZN( u1_u2_u5_n127 ) , .A1( u1_u2_u5_n136 ) , .A3( u1_u2_u5_n148 ) , .A2( u1_u2_u5_n182 ) );
  OAI21_X1 u1_u2_u5_U51 (.ZN( u1_u2_u5_n124 ) , .A( u1_u2_u5_n177 ) , .B2( u1_u2_u5_n183 ) , .B1( u1_u2_u5_n189 ) );
  OAI21_X1 u1_u2_u5_U52 (.ZN( u1_u2_u5_n125 ) , .A( u1_u2_u5_n174 ) , .B2( u1_u2_u5_n185 ) , .B1( u1_u2_u5_n190 ) );
  AOI21_X1 u1_u2_u5_U53 (.A( u1_u2_u5_n153 ) , .B2( u1_u2_u5_n154 ) , .B1( u1_u2_u5_n155 ) , .ZN( u1_u2_u5_n164 ) );
  AOI21_X1 u1_u2_u5_U54 (.ZN( u1_u2_u5_n110 ) , .B1( u1_u2_u5_n122 ) , .B2( u1_u2_u5_n139 ) , .A( u1_u2_u5_n153 ) );
  INV_X1 u1_u2_u5_U55 (.A( u1_u2_u5_n153 ) , .ZN( u1_u2_u5_n176 ) );
  INV_X1 u1_u2_u5_U56 (.A( u1_u2_u5_n126 ) , .ZN( u1_u2_u5_n173 ) );
  AND2_X1 u1_u2_u5_U57 (.A2( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n107 ) , .ZN( u1_u2_u5_n147 ) );
  AND2_X1 u1_u2_u5_U58 (.A2( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n108 ) , .ZN( u1_u2_u5_n148 ) );
  NAND2_X1 u1_u2_u5_U59 (.A1( u1_u2_u5_n105 ) , .A2( u1_u2_u5_n106 ) , .ZN( u1_u2_u5_n158 ) );
  INV_X1 u1_u2_u5_U6 (.A( u1_u2_u5_n135 ) , .ZN( u1_u2_u5_n178 ) );
  NAND2_X1 u1_u2_u5_U60 (.A2( u1_u2_u5_n108 ) , .A1( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n139 ) );
  NAND2_X1 u1_u2_u5_U61 (.A1( u1_u2_u5_n106 ) , .A2( u1_u2_u5_n108 ) , .ZN( u1_u2_u5_n119 ) );
  NAND2_X1 u1_u2_u5_U62 (.A2( u1_u2_u5_n103 ) , .A1( u1_u2_u5_n105 ) , .ZN( u1_u2_u5_n140 ) );
  NAND2_X1 u1_u2_u5_U63 (.A2( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n105 ) , .ZN( u1_u2_u5_n155 ) );
  NAND2_X1 u1_u2_u5_U64 (.A2( u1_u2_u5_n106 ) , .A1( u1_u2_u5_n107 ) , .ZN( u1_u2_u5_n122 ) );
  NAND2_X1 u1_u2_u5_U65 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n106 ) , .ZN( u1_u2_u5_n115 ) );
  NAND2_X1 u1_u2_u5_U66 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n103 ) , .ZN( u1_u2_u5_n161 ) );
  NAND2_X1 u1_u2_u5_U67 (.A1( u1_u2_u5_n105 ) , .A2( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n154 ) );
  INV_X1 u1_u2_u5_U68 (.A( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n172 ) );
  NAND2_X1 u1_u2_u5_U69 (.A1( u1_u2_u5_n103 ) , .A2( u1_u2_u5_n108 ) , .ZN( u1_u2_u5_n123 ) );
  OAI22_X1 u1_u2_u5_U7 (.B2( u1_u2_u5_n149 ) , .B1( u1_u2_u5_n150 ) , .A2( u1_u2_u5_n151 ) , .A1( u1_u2_u5_n152 ) , .ZN( u1_u2_u5_n165 ) );
  NAND2_X1 u1_u2_u5_U70 (.A2( u1_u2_u5_n103 ) , .A1( u1_u2_u5_n107 ) , .ZN( u1_u2_u5_n151 ) );
  NAND2_X1 u1_u2_u5_U71 (.A2( u1_u2_u5_n107 ) , .A1( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n120 ) );
  NAND2_X1 u1_u2_u5_U72 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n157 ) );
  AND2_X1 u1_u2_u5_U73 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n104 ) , .ZN( u1_u2_u5_n131 ) );
  INV_X1 u1_u2_u5_U74 (.A( u1_u2_u5_n102 ) , .ZN( u1_u2_u5_n195 ) );
  OAI221_X1 u1_u2_u5_U75 (.A( u1_u2_u5_n101 ) , .ZN( u1_u2_u5_n102 ) , .C2( u1_u2_u5_n115 ) , .C1( u1_u2_u5_n126 ) , .B1( u1_u2_u5_n134 ) , .B2( u1_u2_u5_n160 ) );
  OAI21_X1 u1_u2_u5_U76 (.ZN( u1_u2_u5_n101 ) , .B1( u1_u2_u5_n137 ) , .A( u1_u2_u5_n146 ) , .B2( u1_u2_u5_n147 ) );
  NOR2_X1 u1_u2_u5_U77 (.A2( u1_u2_X_34 ) , .A1( u1_u2_X_35 ) , .ZN( u1_u2_u5_n145 ) );
  NOR2_X1 u1_u2_u5_U78 (.A2( u1_u2_X_34 ) , .ZN( u1_u2_u5_n146 ) , .A1( u1_u2_u5_n171 ) );
  NOR2_X1 u1_u2_u5_U79 (.A2( u1_u2_X_31 ) , .A1( u1_u2_X_32 ) , .ZN( u1_u2_u5_n103 ) );
  NOR3_X1 u1_u2_u5_U8 (.A2( u1_u2_u5_n147 ) , .A1( u1_u2_u5_n148 ) , .ZN( u1_u2_u5_n149 ) , .A3( u1_u2_u5_n194 ) );
  NOR2_X1 u1_u2_u5_U80 (.A2( u1_u2_X_36 ) , .ZN( u1_u2_u5_n105 ) , .A1( u1_u2_u5_n180 ) );
  NOR2_X1 u1_u2_u5_U81 (.A2( u1_u2_X_33 ) , .ZN( u1_u2_u5_n108 ) , .A1( u1_u2_u5_n170 ) );
  NOR2_X1 u1_u2_u5_U82 (.A2( u1_u2_X_33 ) , .A1( u1_u2_X_36 ) , .ZN( u1_u2_u5_n107 ) );
  NOR2_X1 u1_u2_u5_U83 (.A2( u1_u2_X_31 ) , .ZN( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n181 ) );
  NAND2_X1 u1_u2_u5_U84 (.A2( u1_u2_X_34 ) , .A1( u1_u2_X_35 ) , .ZN( u1_u2_u5_n153 ) );
  NAND2_X1 u1_u2_u5_U85 (.A1( u1_u2_X_34 ) , .ZN( u1_u2_u5_n126 ) , .A2( u1_u2_u5_n171 ) );
  AND2_X1 u1_u2_u5_U86 (.A1( u1_u2_X_31 ) , .A2( u1_u2_X_32 ) , .ZN( u1_u2_u5_n106 ) );
  AND2_X1 u1_u2_u5_U87 (.A1( u1_u2_X_31 ) , .ZN( u1_u2_u5_n109 ) , .A2( u1_u2_u5_n181 ) );
  INV_X1 u1_u2_u5_U88 (.A( u1_u2_X_33 ) , .ZN( u1_u2_u5_n180 ) );
  INV_X1 u1_u2_u5_U89 (.A( u1_u2_X_35 ) , .ZN( u1_u2_u5_n171 ) );
  NOR2_X1 u1_u2_u5_U9 (.ZN( u1_u2_u5_n135 ) , .A1( u1_u2_u5_n173 ) , .A2( u1_u2_u5_n176 ) );
  INV_X1 u1_u2_u5_U90 (.A( u1_u2_X_36 ) , .ZN( u1_u2_u5_n170 ) );
  INV_X1 u1_u2_u5_U91 (.A( u1_u2_X_32 ) , .ZN( u1_u2_u5_n181 ) );
  NAND4_X1 u1_u2_u5_U92 (.ZN( u1_out2_29 ) , .A4( u1_u2_u5_n129 ) , .A3( u1_u2_u5_n130 ) , .A2( u1_u2_u5_n168 ) , .A1( u1_u2_u5_n196 ) );
  AOI221_X1 u1_u2_u5_U93 (.A( u1_u2_u5_n128 ) , .ZN( u1_u2_u5_n129 ) , .C2( u1_u2_u5_n132 ) , .B2( u1_u2_u5_n159 ) , .B1( u1_u2_u5_n176 ) , .C1( u1_u2_u5_n184 ) );
  AOI222_X1 u1_u2_u5_U94 (.ZN( u1_u2_u5_n130 ) , .A2( u1_u2_u5_n146 ) , .B1( u1_u2_u5_n147 ) , .C2( u1_u2_u5_n175 ) , .B2( u1_u2_u5_n179 ) , .A1( u1_u2_u5_n188 ) , .C1( u1_u2_u5_n194 ) );
  NAND4_X1 u1_u2_u5_U95 (.ZN( u1_out2_19 ) , .A4( u1_u2_u5_n166 ) , .A3( u1_u2_u5_n167 ) , .A2( u1_u2_u5_n168 ) , .A1( u1_u2_u5_n169 ) );
  AOI22_X1 u1_u2_u5_U96 (.B2( u1_u2_u5_n145 ) , .A2( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n167 ) , .B1( u1_u2_u5_n182 ) , .A1( u1_u2_u5_n189 ) );
  NOR4_X1 u1_u2_u5_U97 (.A4( u1_u2_u5_n162 ) , .A3( u1_u2_u5_n163 ) , .A2( u1_u2_u5_n164 ) , .A1( u1_u2_u5_n165 ) , .ZN( u1_u2_u5_n166 ) );
  NAND4_X1 u1_u2_u5_U98 (.ZN( u1_out2_11 ) , .A4( u1_u2_u5_n143 ) , .A3( u1_u2_u5_n144 ) , .A2( u1_u2_u5_n169 ) , .A1( u1_u2_u5_n196 ) );
  AOI22_X1 u1_u2_u5_U99 (.A2( u1_u2_u5_n132 ) , .ZN( u1_u2_u5_n144 ) , .B2( u1_u2_u5_n145 ) , .B1( u1_u2_u5_n184 ) , .A1( u1_u2_u5_n194 ) );
  XOR2_X1 u1_u4_U13 (.B( u1_K5_42 ) , .A( u1_R3_29 ) , .Z( u1_u4_X_42 ) );
  XOR2_X1 u1_u4_U14 (.B( u1_K5_41 ) , .A( u1_R3_28 ) , .Z( u1_u4_X_41 ) );
  XOR2_X1 u1_u4_U15 (.B( u1_K5_40 ) , .A( u1_R3_27 ) , .Z( u1_u4_X_40 ) );
  XOR2_X1 u1_u4_U17 (.B( u1_K5_39 ) , .A( u1_R3_26 ) , .Z( u1_u4_X_39 ) );
  XOR2_X1 u1_u4_U18 (.B( u1_K5_38 ) , .A( u1_R3_25 ) , .Z( u1_u4_X_38 ) );
  XOR2_X1 u1_u4_U19 (.B( u1_K5_37 ) , .A( u1_R3_24 ) , .Z( u1_u4_X_37 ) );
  AOI22_X1 u1_u4_u6_U10 (.A2( u1_u4_u6_n151 ) , .B2( u1_u4_u6_n161 ) , .A1( u1_u4_u6_n167 ) , .B1( u1_u4_u6_n170 ) , .ZN( u1_u4_u6_n89 ) );
  AOI21_X1 u1_u4_u6_U11 (.B1( u1_u4_u6_n107 ) , .B2( u1_u4_u6_n132 ) , .A( u1_u4_u6_n158 ) , .ZN( u1_u4_u6_n88 ) );
  AOI21_X1 u1_u4_u6_U12 (.B2( u1_u4_u6_n147 ) , .B1( u1_u4_u6_n148 ) , .ZN( u1_u4_u6_n149 ) , .A( u1_u4_u6_n158 ) );
  AOI21_X1 u1_u4_u6_U13 (.ZN( u1_u4_u6_n106 ) , .A( u1_u4_u6_n142 ) , .B2( u1_u4_u6_n159 ) , .B1( u1_u4_u6_n164 ) );
  INV_X1 u1_u4_u6_U14 (.A( u1_u4_u6_n155 ) , .ZN( u1_u4_u6_n161 ) );
  INV_X1 u1_u4_u6_U15 (.A( u1_u4_u6_n128 ) , .ZN( u1_u4_u6_n164 ) );
  NAND2_X1 u1_u4_u6_U16 (.ZN( u1_u4_u6_n110 ) , .A1( u1_u4_u6_n122 ) , .A2( u1_u4_u6_n129 ) );
  NAND2_X1 u1_u4_u6_U17 (.ZN( u1_u4_u6_n124 ) , .A2( u1_u4_u6_n146 ) , .A1( u1_u4_u6_n148 ) );
  INV_X1 u1_u4_u6_U18 (.A( u1_u4_u6_n132 ) , .ZN( u1_u4_u6_n171 ) );
  AND2_X1 u1_u4_u6_U19 (.A1( u1_u4_u6_n100 ) , .ZN( u1_u4_u6_n130 ) , .A2( u1_u4_u6_n147 ) );
  INV_X1 u1_u4_u6_U20 (.A( u1_u4_u6_n127 ) , .ZN( u1_u4_u6_n173 ) );
  INV_X1 u1_u4_u6_U21 (.A( u1_u4_u6_n121 ) , .ZN( u1_u4_u6_n167 ) );
  INV_X1 u1_u4_u6_U22 (.A( u1_u4_u6_n100 ) , .ZN( u1_u4_u6_n169 ) );
  INV_X1 u1_u4_u6_U23 (.A( u1_u4_u6_n123 ) , .ZN( u1_u4_u6_n170 ) );
  INV_X1 u1_u4_u6_U24 (.A( u1_u4_u6_n113 ) , .ZN( u1_u4_u6_n168 ) );
  AND2_X1 u1_u4_u6_U25 (.A1( u1_u4_u6_n107 ) , .A2( u1_u4_u6_n119 ) , .ZN( u1_u4_u6_n133 ) );
  AND2_X1 u1_u4_u6_U26 (.A2( u1_u4_u6_n121 ) , .A1( u1_u4_u6_n122 ) , .ZN( u1_u4_u6_n131 ) );
  AND3_X1 u1_u4_u6_U27 (.ZN( u1_u4_u6_n120 ) , .A2( u1_u4_u6_n127 ) , .A1( u1_u4_u6_n132 ) , .A3( u1_u4_u6_n145 ) );
  INV_X1 u1_u4_u6_U28 (.A( u1_u4_u6_n146 ) , .ZN( u1_u4_u6_n163 ) );
  AOI222_X1 u1_u4_u6_U29 (.ZN( u1_u4_u6_n114 ) , .A1( u1_u4_u6_n118 ) , .A2( u1_u4_u6_n126 ) , .B2( u1_u4_u6_n151 ) , .C2( u1_u4_u6_n159 ) , .C1( u1_u4_u6_n168 ) , .B1( u1_u4_u6_n169 ) );
  INV_X1 u1_u4_u6_U3 (.A( u1_u4_u6_n110 ) , .ZN( u1_u4_u6_n166 ) );
  NOR2_X1 u1_u4_u6_U30 (.A1( u1_u4_u6_n162 ) , .A2( u1_u4_u6_n165 ) , .ZN( u1_u4_u6_n98 ) );
  NAND2_X1 u1_u4_u6_U31 (.A1( u1_u4_u6_n144 ) , .ZN( u1_u4_u6_n151 ) , .A2( u1_u4_u6_n158 ) );
  NAND2_X1 u1_u4_u6_U32 (.ZN( u1_u4_u6_n132 ) , .A1( u1_u4_u6_n91 ) , .A2( u1_u4_u6_n97 ) );
  AOI22_X1 u1_u4_u6_U33 (.B2( u1_u4_u6_n110 ) , .B1( u1_u4_u6_n111 ) , .A1( u1_u4_u6_n112 ) , .ZN( u1_u4_u6_n115 ) , .A2( u1_u4_u6_n161 ) );
  NAND4_X1 u1_u4_u6_U34 (.A3( u1_u4_u6_n109 ) , .ZN( u1_u4_u6_n112 ) , .A4( u1_u4_u6_n132 ) , .A2( u1_u4_u6_n147 ) , .A1( u1_u4_u6_n166 ) );
  NOR2_X1 u1_u4_u6_U35 (.ZN( u1_u4_u6_n109 ) , .A1( u1_u4_u6_n170 ) , .A2( u1_u4_u6_n173 ) );
  NOR2_X1 u1_u4_u6_U36 (.A2( u1_u4_u6_n126 ) , .ZN( u1_u4_u6_n155 ) , .A1( u1_u4_u6_n160 ) );
  NAND2_X1 u1_u4_u6_U37 (.ZN( u1_u4_u6_n146 ) , .A2( u1_u4_u6_n94 ) , .A1( u1_u4_u6_n99 ) );
  AOI21_X1 u1_u4_u6_U38 (.A( u1_u4_u6_n144 ) , .B2( u1_u4_u6_n145 ) , .B1( u1_u4_u6_n146 ) , .ZN( u1_u4_u6_n150 ) );
  AOI211_X1 u1_u4_u6_U39 (.B( u1_u4_u6_n134 ) , .A( u1_u4_u6_n135 ) , .C1( u1_u4_u6_n136 ) , .ZN( u1_u4_u6_n137 ) , .C2( u1_u4_u6_n151 ) );
  INV_X1 u1_u4_u6_U4 (.A( u1_u4_u6_n142 ) , .ZN( u1_u4_u6_n174 ) );
  NAND4_X1 u1_u4_u6_U40 (.A4( u1_u4_u6_n127 ) , .A3( u1_u4_u6_n128 ) , .A2( u1_u4_u6_n129 ) , .A1( u1_u4_u6_n130 ) , .ZN( u1_u4_u6_n136 ) );
  AOI21_X1 u1_u4_u6_U41 (.B2( u1_u4_u6_n132 ) , .B1( u1_u4_u6_n133 ) , .ZN( u1_u4_u6_n134 ) , .A( u1_u4_u6_n158 ) );
  AOI21_X1 u1_u4_u6_U42 (.B1( u1_u4_u6_n131 ) , .ZN( u1_u4_u6_n135 ) , .A( u1_u4_u6_n144 ) , .B2( u1_u4_u6_n146 ) );
  INV_X1 u1_u4_u6_U43 (.A( u1_u4_u6_n111 ) , .ZN( u1_u4_u6_n158 ) );
  NAND2_X1 u1_u4_u6_U44 (.ZN( u1_u4_u6_n127 ) , .A1( u1_u4_u6_n91 ) , .A2( u1_u4_u6_n92 ) );
  NAND2_X1 u1_u4_u6_U45 (.ZN( u1_u4_u6_n129 ) , .A2( u1_u4_u6_n95 ) , .A1( u1_u4_u6_n96 ) );
  INV_X1 u1_u4_u6_U46 (.A( u1_u4_u6_n144 ) , .ZN( u1_u4_u6_n159 ) );
  NAND2_X1 u1_u4_u6_U47 (.ZN( u1_u4_u6_n145 ) , .A2( u1_u4_u6_n97 ) , .A1( u1_u4_u6_n98 ) );
  NAND2_X1 u1_u4_u6_U48 (.ZN( u1_u4_u6_n148 ) , .A2( u1_u4_u6_n92 ) , .A1( u1_u4_u6_n94 ) );
  NAND2_X1 u1_u4_u6_U49 (.ZN( u1_u4_u6_n108 ) , .A2( u1_u4_u6_n139 ) , .A1( u1_u4_u6_n144 ) );
  NAND2_X1 u1_u4_u6_U5 (.A2( u1_u4_u6_n143 ) , .ZN( u1_u4_u6_n152 ) , .A1( u1_u4_u6_n166 ) );
  NAND2_X1 u1_u4_u6_U50 (.ZN( u1_u4_u6_n121 ) , .A2( u1_u4_u6_n95 ) , .A1( u1_u4_u6_n97 ) );
  NAND2_X1 u1_u4_u6_U51 (.ZN( u1_u4_u6_n107 ) , .A2( u1_u4_u6_n92 ) , .A1( u1_u4_u6_n95 ) );
  AND2_X1 u1_u4_u6_U52 (.ZN( u1_u4_u6_n118 ) , .A2( u1_u4_u6_n91 ) , .A1( u1_u4_u6_n99 ) );
  NAND2_X1 u1_u4_u6_U53 (.ZN( u1_u4_u6_n147 ) , .A2( u1_u4_u6_n98 ) , .A1( u1_u4_u6_n99 ) );
  NAND2_X1 u1_u4_u6_U54 (.ZN( u1_u4_u6_n128 ) , .A1( u1_u4_u6_n94 ) , .A2( u1_u4_u6_n96 ) );
  NAND2_X1 u1_u4_u6_U55 (.ZN( u1_u4_u6_n119 ) , .A2( u1_u4_u6_n95 ) , .A1( u1_u4_u6_n99 ) );
  NAND2_X1 u1_u4_u6_U56 (.ZN( u1_u4_u6_n123 ) , .A2( u1_u4_u6_n91 ) , .A1( u1_u4_u6_n96 ) );
  NAND2_X1 u1_u4_u6_U57 (.ZN( u1_u4_u6_n100 ) , .A2( u1_u4_u6_n92 ) , .A1( u1_u4_u6_n98 ) );
  NAND2_X1 u1_u4_u6_U58 (.ZN( u1_u4_u6_n122 ) , .A1( u1_u4_u6_n94 ) , .A2( u1_u4_u6_n97 ) );
  INV_X1 u1_u4_u6_U59 (.A( u1_u4_u6_n139 ) , .ZN( u1_u4_u6_n160 ) );
  AOI22_X1 u1_u4_u6_U6 (.B2( u1_u4_u6_n101 ) , .A1( u1_u4_u6_n102 ) , .ZN( u1_u4_u6_n103 ) , .B1( u1_u4_u6_n160 ) , .A2( u1_u4_u6_n161 ) );
  NAND2_X1 u1_u4_u6_U60 (.ZN( u1_u4_u6_n113 ) , .A1( u1_u4_u6_n96 ) , .A2( u1_u4_u6_n98 ) );
  NOR2_X1 u1_u4_u6_U61 (.A2( u1_u4_X_40 ) , .A1( u1_u4_X_41 ) , .ZN( u1_u4_u6_n126 ) );
  NOR2_X1 u1_u4_u6_U62 (.A2( u1_u4_X_39 ) , .A1( u1_u4_X_42 ) , .ZN( u1_u4_u6_n92 ) );
  NOR2_X1 u1_u4_u6_U63 (.A2( u1_u4_X_39 ) , .A1( u1_u4_u6_n156 ) , .ZN( u1_u4_u6_n97 ) );
  NOR2_X1 u1_u4_u6_U64 (.A2( u1_u4_X_38 ) , .A1( u1_u4_u6_n165 ) , .ZN( u1_u4_u6_n95 ) );
  NOR2_X1 u1_u4_u6_U65 (.A2( u1_u4_X_41 ) , .ZN( u1_u4_u6_n111 ) , .A1( u1_u4_u6_n157 ) );
  NOR2_X1 u1_u4_u6_U66 (.A2( u1_u4_X_37 ) , .A1( u1_u4_u6_n162 ) , .ZN( u1_u4_u6_n94 ) );
  NOR2_X1 u1_u4_u6_U67 (.A2( u1_u4_X_37 ) , .A1( u1_u4_X_38 ) , .ZN( u1_u4_u6_n91 ) );
  NAND2_X1 u1_u4_u6_U68 (.A1( u1_u4_X_41 ) , .ZN( u1_u4_u6_n144 ) , .A2( u1_u4_u6_n157 ) );
  NAND2_X1 u1_u4_u6_U69 (.A2( u1_u4_X_40 ) , .A1( u1_u4_X_41 ) , .ZN( u1_u4_u6_n139 ) );
  NOR2_X1 u1_u4_u6_U7 (.A1( u1_u4_u6_n118 ) , .ZN( u1_u4_u6_n143 ) , .A2( u1_u4_u6_n168 ) );
  AND2_X1 u1_u4_u6_U70 (.A1( u1_u4_X_39 ) , .A2( u1_u4_u6_n156 ) , .ZN( u1_u4_u6_n96 ) );
  AND2_X1 u1_u4_u6_U71 (.A1( u1_u4_X_39 ) , .A2( u1_u4_X_42 ) , .ZN( u1_u4_u6_n99 ) );
  INV_X1 u1_u4_u6_U72 (.A( u1_u4_X_40 ) , .ZN( u1_u4_u6_n157 ) );
  INV_X1 u1_u4_u6_U73 (.A( u1_u4_X_37 ) , .ZN( u1_u4_u6_n165 ) );
  INV_X1 u1_u4_u6_U74 (.A( u1_u4_X_38 ) , .ZN( u1_u4_u6_n162 ) );
  INV_X1 u1_u4_u6_U75 (.A( u1_u4_X_42 ) , .ZN( u1_u4_u6_n156 ) );
  NAND4_X1 u1_u4_u6_U76 (.ZN( u1_out4_32 ) , .A4( u1_u4_u6_n103 ) , .A3( u1_u4_u6_n104 ) , .A2( u1_u4_u6_n105 ) , .A1( u1_u4_u6_n106 ) );
  AOI22_X1 u1_u4_u6_U77 (.ZN( u1_u4_u6_n105 ) , .A2( u1_u4_u6_n108 ) , .A1( u1_u4_u6_n118 ) , .B2( u1_u4_u6_n126 ) , .B1( u1_u4_u6_n171 ) );
  AOI22_X1 u1_u4_u6_U78 (.ZN( u1_u4_u6_n104 ) , .A1( u1_u4_u6_n111 ) , .B1( u1_u4_u6_n124 ) , .B2( u1_u4_u6_n151 ) , .A2( u1_u4_u6_n93 ) );
  NAND4_X1 u1_u4_u6_U79 (.ZN( u1_out4_12 ) , .A4( u1_u4_u6_n114 ) , .A3( u1_u4_u6_n115 ) , .A2( u1_u4_u6_n116 ) , .A1( u1_u4_u6_n117 ) );
  INV_X1 u1_u4_u6_U8 (.ZN( u1_u4_u6_n172 ) , .A( u1_u4_u6_n88 ) );
  OAI22_X1 u1_u4_u6_U80 (.B2( u1_u4_u6_n111 ) , .ZN( u1_u4_u6_n116 ) , .B1( u1_u4_u6_n126 ) , .A2( u1_u4_u6_n164 ) , .A1( u1_u4_u6_n167 ) );
  OAI21_X1 u1_u4_u6_U81 (.A( u1_u4_u6_n108 ) , .ZN( u1_u4_u6_n117 ) , .B2( u1_u4_u6_n141 ) , .B1( u1_u4_u6_n163 ) );
  OAI211_X1 u1_u4_u6_U82 (.ZN( u1_out4_22 ) , .B( u1_u4_u6_n137 ) , .A( u1_u4_u6_n138 ) , .C2( u1_u4_u6_n139 ) , .C1( u1_u4_u6_n140 ) );
  AOI22_X1 u1_u4_u6_U83 (.B1( u1_u4_u6_n124 ) , .A2( u1_u4_u6_n125 ) , .A1( u1_u4_u6_n126 ) , .ZN( u1_u4_u6_n138 ) , .B2( u1_u4_u6_n161 ) );
  AND4_X1 u1_u4_u6_U84 (.A3( u1_u4_u6_n119 ) , .A1( u1_u4_u6_n120 ) , .A4( u1_u4_u6_n129 ) , .ZN( u1_u4_u6_n140 ) , .A2( u1_u4_u6_n143 ) );
  OAI211_X1 u1_u4_u6_U85 (.ZN( u1_out4_7 ) , .B( u1_u4_u6_n153 ) , .C2( u1_u4_u6_n154 ) , .C1( u1_u4_u6_n155 ) , .A( u1_u4_u6_n174 ) );
  NOR3_X1 u1_u4_u6_U86 (.A1( u1_u4_u6_n141 ) , .ZN( u1_u4_u6_n154 ) , .A3( u1_u4_u6_n164 ) , .A2( u1_u4_u6_n171 ) );
  AOI211_X1 u1_u4_u6_U87 (.B( u1_u4_u6_n149 ) , .A( u1_u4_u6_n150 ) , .C2( u1_u4_u6_n151 ) , .C1( u1_u4_u6_n152 ) , .ZN( u1_u4_u6_n153 ) );
  NAND3_X1 u1_u4_u6_U88 (.A2( u1_u4_u6_n123 ) , .ZN( u1_u4_u6_n125 ) , .A1( u1_u4_u6_n130 ) , .A3( u1_u4_u6_n131 ) );
  NAND3_X1 u1_u4_u6_U89 (.A3( u1_u4_u6_n133 ) , .ZN( u1_u4_u6_n141 ) , .A1( u1_u4_u6_n145 ) , .A2( u1_u4_u6_n148 ) );
  OAI21_X1 u1_u4_u6_U9 (.A( u1_u4_u6_n159 ) , .B1( u1_u4_u6_n169 ) , .B2( u1_u4_u6_n173 ) , .ZN( u1_u4_u6_n90 ) );
  NAND3_X1 u1_u4_u6_U90 (.ZN( u1_u4_u6_n101 ) , .A3( u1_u4_u6_n107 ) , .A2( u1_u4_u6_n121 ) , .A1( u1_u4_u6_n127 ) );
  NAND3_X1 u1_u4_u6_U91 (.ZN( u1_u4_u6_n102 ) , .A3( u1_u4_u6_n130 ) , .A2( u1_u4_u6_n145 ) , .A1( u1_u4_u6_n166 ) );
  NAND3_X1 u1_u4_u6_U92 (.A3( u1_u4_u6_n113 ) , .A1( u1_u4_u6_n119 ) , .A2( u1_u4_u6_n123 ) , .ZN( u1_u4_u6_n93 ) );
  NAND3_X1 u1_u4_u6_U93 (.ZN( u1_u4_u6_n142 ) , .A2( u1_u4_u6_n172 ) , .A3( u1_u4_u6_n89 ) , .A1( u1_u4_u6_n90 ) );
  XOR2_X1 u1_u5_U1 (.B( u1_K6_9 ) , .A( u1_R4_6 ) , .Z( u1_u5_X_9 ) );
  XOR2_X1 u1_u5_U10 (.B( u1_K6_45 ) , .A( u1_R4_30 ) , .Z( u1_u5_X_45 ) );
  XOR2_X1 u1_u5_U11 (.B( u1_K6_44 ) , .A( u1_R4_29 ) , .Z( u1_u5_X_44 ) );
  XOR2_X1 u1_u5_U12 (.B( u1_K6_43 ) , .A( u1_R4_28 ) , .Z( u1_u5_X_43 ) );
  XOR2_X1 u1_u5_U2 (.B( u1_K6_8 ) , .A( u1_R4_5 ) , .Z( u1_u5_X_8 ) );
  XOR2_X1 u1_u5_U3 (.B( u1_K6_7 ) , .A( u1_R4_4 ) , .Z( u1_u5_X_7 ) );
  XOR2_X1 u1_u5_U46 (.B( u1_K6_12 ) , .A( u1_R4_9 ) , .Z( u1_u5_X_12 ) );
  XOR2_X1 u1_u5_U47 (.B( u1_K6_11 ) , .A( u1_R4_8 ) , .Z( u1_u5_X_11 ) );
  XOR2_X1 u1_u5_U48 (.B( u1_K6_10 ) , .A( u1_R4_7 ) , .Z( u1_u5_X_10 ) );
  XOR2_X1 u1_u5_U7 (.B( u1_K6_48 ) , .A( u1_R4_1 ) , .Z( u1_u5_X_48 ) );
  XOR2_X1 u1_u5_U8 (.B( u1_K6_47 ) , .A( u1_R4_32 ) , .Z( u1_u5_X_47 ) );
  XOR2_X1 u1_u5_U9 (.B( u1_K6_46 ) , .A( u1_R4_31 ) , .Z( u1_u5_X_46 ) );
  AOI21_X1 u1_u5_u1_U10 (.B2( u1_u5_u1_n155 ) , .B1( u1_u5_u1_n156 ) , .ZN( u1_u5_u1_n157 ) , .A( u1_u5_u1_n174 ) );
  NAND3_X1 u1_u5_u1_U100 (.ZN( u1_u5_u1_n113 ) , .A1( u1_u5_u1_n120 ) , .A3( u1_u5_u1_n133 ) , .A2( u1_u5_u1_n155 ) );
  NAND2_X1 u1_u5_u1_U11 (.ZN( u1_u5_u1_n140 ) , .A2( u1_u5_u1_n150 ) , .A1( u1_u5_u1_n155 ) );
  NAND2_X1 u1_u5_u1_U12 (.A1( u1_u5_u1_n131 ) , .ZN( u1_u5_u1_n147 ) , .A2( u1_u5_u1_n153 ) );
  INV_X1 u1_u5_u1_U13 (.A( u1_u5_u1_n139 ) , .ZN( u1_u5_u1_n174 ) );
  OR4_X1 u1_u5_u1_U14 (.A4( u1_u5_u1_n106 ) , .A3( u1_u5_u1_n107 ) , .ZN( u1_u5_u1_n108 ) , .A1( u1_u5_u1_n117 ) , .A2( u1_u5_u1_n184 ) );
  AOI21_X1 u1_u5_u1_U15 (.ZN( u1_u5_u1_n106 ) , .A( u1_u5_u1_n112 ) , .B1( u1_u5_u1_n154 ) , .B2( u1_u5_u1_n156 ) );
  INV_X1 u1_u5_u1_U16 (.A( u1_u5_u1_n101 ) , .ZN( u1_u5_u1_n184 ) );
  AOI21_X1 u1_u5_u1_U17 (.ZN( u1_u5_u1_n107 ) , .B1( u1_u5_u1_n134 ) , .B2( u1_u5_u1_n149 ) , .A( u1_u5_u1_n174 ) );
  INV_X1 u1_u5_u1_U18 (.A( u1_u5_u1_n112 ) , .ZN( u1_u5_u1_n171 ) );
  NAND2_X1 u1_u5_u1_U19 (.ZN( u1_u5_u1_n141 ) , .A1( u1_u5_u1_n153 ) , .A2( u1_u5_u1_n156 ) );
  AND2_X1 u1_u5_u1_U20 (.A1( u1_u5_u1_n123 ) , .ZN( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n161 ) );
  NAND2_X1 u1_u5_u1_U21 (.A2( u1_u5_u1_n115 ) , .A1( u1_u5_u1_n116 ) , .ZN( u1_u5_u1_n148 ) );
  NAND2_X1 u1_u5_u1_U22 (.A2( u1_u5_u1_n133 ) , .A1( u1_u5_u1_n135 ) , .ZN( u1_u5_u1_n159 ) );
  NAND2_X1 u1_u5_u1_U23 (.A2( u1_u5_u1_n115 ) , .A1( u1_u5_u1_n120 ) , .ZN( u1_u5_u1_n132 ) );
  INV_X1 u1_u5_u1_U24 (.A( u1_u5_u1_n154 ) , .ZN( u1_u5_u1_n178 ) );
  AOI22_X1 u1_u5_u1_U25 (.B2( u1_u5_u1_n113 ) , .A2( u1_u5_u1_n114 ) , .ZN( u1_u5_u1_n125 ) , .A1( u1_u5_u1_n171 ) , .B1( u1_u5_u1_n173 ) );
  NAND2_X1 u1_u5_u1_U26 (.ZN( u1_u5_u1_n114 ) , .A1( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n156 ) );
  INV_X1 u1_u5_u1_U27 (.A( u1_u5_u1_n151 ) , .ZN( u1_u5_u1_n183 ) );
  AND2_X1 u1_u5_u1_U28 (.A1( u1_u5_u1_n129 ) , .A2( u1_u5_u1_n133 ) , .ZN( u1_u5_u1_n149 ) );
  INV_X1 u1_u5_u1_U29 (.A( u1_u5_u1_n131 ) , .ZN( u1_u5_u1_n180 ) );
  INV_X1 u1_u5_u1_U3 (.A( u1_u5_u1_n159 ) , .ZN( u1_u5_u1_n182 ) );
  OAI221_X1 u1_u5_u1_U30 (.A( u1_u5_u1_n119 ) , .C2( u1_u5_u1_n129 ) , .ZN( u1_u5_u1_n138 ) , .B2( u1_u5_u1_n152 ) , .C1( u1_u5_u1_n174 ) , .B1( u1_u5_u1_n187 ) );
  INV_X1 u1_u5_u1_U31 (.A( u1_u5_u1_n148 ) , .ZN( u1_u5_u1_n187 ) );
  AOI211_X1 u1_u5_u1_U32 (.B( u1_u5_u1_n117 ) , .A( u1_u5_u1_n118 ) , .ZN( u1_u5_u1_n119 ) , .C2( u1_u5_u1_n146 ) , .C1( u1_u5_u1_n159 ) );
  NOR2_X1 u1_u5_u1_U33 (.A1( u1_u5_u1_n168 ) , .A2( u1_u5_u1_n176 ) , .ZN( u1_u5_u1_n98 ) );
  AOI211_X1 u1_u5_u1_U34 (.B( u1_u5_u1_n162 ) , .A( u1_u5_u1_n163 ) , .C2( u1_u5_u1_n164 ) , .ZN( u1_u5_u1_n165 ) , .C1( u1_u5_u1_n171 ) );
  AOI21_X1 u1_u5_u1_U35 (.A( u1_u5_u1_n160 ) , .B2( u1_u5_u1_n161 ) , .ZN( u1_u5_u1_n162 ) , .B1( u1_u5_u1_n182 ) );
  OR2_X1 u1_u5_u1_U36 (.A2( u1_u5_u1_n157 ) , .A1( u1_u5_u1_n158 ) , .ZN( u1_u5_u1_n163 ) );
  OAI21_X1 u1_u5_u1_U37 (.B2( u1_u5_u1_n123 ) , .ZN( u1_u5_u1_n145 ) , .B1( u1_u5_u1_n160 ) , .A( u1_u5_u1_n185 ) );
  INV_X1 u1_u5_u1_U38 (.A( u1_u5_u1_n122 ) , .ZN( u1_u5_u1_n185 ) );
  AOI21_X1 u1_u5_u1_U39 (.B2( u1_u5_u1_n120 ) , .B1( u1_u5_u1_n121 ) , .ZN( u1_u5_u1_n122 ) , .A( u1_u5_u1_n128 ) );
  AOI221_X1 u1_u5_u1_U4 (.A( u1_u5_u1_n138 ) , .C2( u1_u5_u1_n139 ) , .C1( u1_u5_u1_n140 ) , .B2( u1_u5_u1_n141 ) , .ZN( u1_u5_u1_n142 ) , .B1( u1_u5_u1_n175 ) );
  NAND2_X1 u1_u5_u1_U40 (.A1( u1_u5_u1_n128 ) , .ZN( u1_u5_u1_n146 ) , .A2( u1_u5_u1_n160 ) );
  NAND2_X1 u1_u5_u1_U41 (.A2( u1_u5_u1_n112 ) , .ZN( u1_u5_u1_n139 ) , .A1( u1_u5_u1_n152 ) );
  NAND2_X1 u1_u5_u1_U42 (.A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n156 ) , .A2( u1_u5_u1_n99 ) );
  AOI221_X1 u1_u5_u1_U43 (.B1( u1_u5_u1_n140 ) , .ZN( u1_u5_u1_n167 ) , .B2( u1_u5_u1_n172 ) , .C2( u1_u5_u1_n175 ) , .C1( u1_u5_u1_n178 ) , .A( u1_u5_u1_n188 ) );
  INV_X1 u1_u5_u1_U44 (.ZN( u1_u5_u1_n188 ) , .A( u1_u5_u1_n97 ) );
  AOI211_X1 u1_u5_u1_U45 (.A( u1_u5_u1_n118 ) , .C1( u1_u5_u1_n132 ) , .C2( u1_u5_u1_n139 ) , .B( u1_u5_u1_n96 ) , .ZN( u1_u5_u1_n97 ) );
  AOI21_X1 u1_u5_u1_U46 (.B2( u1_u5_u1_n121 ) , .B1( u1_u5_u1_n135 ) , .A( u1_u5_u1_n152 ) , .ZN( u1_u5_u1_n96 ) );
  NOR2_X1 u1_u5_u1_U47 (.ZN( u1_u5_u1_n117 ) , .A1( u1_u5_u1_n121 ) , .A2( u1_u5_u1_n160 ) );
  AOI21_X1 u1_u5_u1_U48 (.A( u1_u5_u1_n128 ) , .B2( u1_u5_u1_n129 ) , .ZN( u1_u5_u1_n130 ) , .B1( u1_u5_u1_n150 ) );
  NAND2_X1 u1_u5_u1_U49 (.ZN( u1_u5_u1_n112 ) , .A1( u1_u5_u1_n169 ) , .A2( u1_u5_u1_n170 ) );
  AOI211_X1 u1_u5_u1_U5 (.ZN( u1_u5_u1_n124 ) , .A( u1_u5_u1_n138 ) , .C2( u1_u5_u1_n139 ) , .B( u1_u5_u1_n145 ) , .C1( u1_u5_u1_n147 ) );
  NAND2_X1 u1_u5_u1_U50 (.ZN( u1_u5_u1_n129 ) , .A2( u1_u5_u1_n95 ) , .A1( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U51 (.A1( u1_u5_u1_n102 ) , .ZN( u1_u5_u1_n154 ) , .A2( u1_u5_u1_n99 ) );
  NAND2_X1 u1_u5_u1_U52 (.A2( u1_u5_u1_n100 ) , .ZN( u1_u5_u1_n135 ) , .A1( u1_u5_u1_n99 ) );
  AOI21_X1 u1_u5_u1_U53 (.A( u1_u5_u1_n152 ) , .B2( u1_u5_u1_n153 ) , .B1( u1_u5_u1_n154 ) , .ZN( u1_u5_u1_n158 ) );
  INV_X1 u1_u5_u1_U54 (.A( u1_u5_u1_n160 ) , .ZN( u1_u5_u1_n175 ) );
  NAND2_X1 u1_u5_u1_U55 (.A1( u1_u5_u1_n100 ) , .ZN( u1_u5_u1_n116 ) , .A2( u1_u5_u1_n95 ) );
  NAND2_X1 u1_u5_u1_U56 (.A1( u1_u5_u1_n102 ) , .ZN( u1_u5_u1_n131 ) , .A2( u1_u5_u1_n95 ) );
  NAND2_X1 u1_u5_u1_U57 (.A2( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n121 ) , .A1( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U58 (.A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n153 ) , .A2( u1_u5_u1_n98 ) );
  NAND2_X1 u1_u5_u1_U59 (.A2( u1_u5_u1_n104 ) , .A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n133 ) );
  AOI22_X1 u1_u5_u1_U6 (.B2( u1_u5_u1_n136 ) , .A2( u1_u5_u1_n137 ) , .ZN( u1_u5_u1_n143 ) , .A1( u1_u5_u1_n171 ) , .B1( u1_u5_u1_n173 ) );
  NAND2_X1 u1_u5_u1_U60 (.ZN( u1_u5_u1_n150 ) , .A2( u1_u5_u1_n98 ) , .A1( u1_u5_u1_n99 ) );
  NAND2_X1 u1_u5_u1_U61 (.A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n155 ) , .A2( u1_u5_u1_n95 ) );
  OAI21_X1 u1_u5_u1_U62 (.ZN( u1_u5_u1_n109 ) , .B1( u1_u5_u1_n129 ) , .B2( u1_u5_u1_n160 ) , .A( u1_u5_u1_n167 ) );
  NAND2_X1 u1_u5_u1_U63 (.A2( u1_u5_u1_n100 ) , .A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n120 ) );
  NAND2_X1 u1_u5_u1_U64 (.A1( u1_u5_u1_n102 ) , .A2( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n115 ) );
  NAND2_X1 u1_u5_u1_U65 (.A2( u1_u5_u1_n100 ) , .A1( u1_u5_u1_n104 ) , .ZN( u1_u5_u1_n151 ) );
  NAND2_X1 u1_u5_u1_U66 (.A2( u1_u5_u1_n103 ) , .A1( u1_u5_u1_n105 ) , .ZN( u1_u5_u1_n161 ) );
  INV_X1 u1_u5_u1_U67 (.A( u1_u5_u1_n152 ) , .ZN( u1_u5_u1_n173 ) );
  INV_X1 u1_u5_u1_U68 (.A( u1_u5_u1_n128 ) , .ZN( u1_u5_u1_n172 ) );
  NAND2_X1 u1_u5_u1_U69 (.A2( u1_u5_u1_n102 ) , .A1( u1_u5_u1_n103 ) , .ZN( u1_u5_u1_n123 ) );
  INV_X1 u1_u5_u1_U7 (.A( u1_u5_u1_n147 ) , .ZN( u1_u5_u1_n181 ) );
  NOR2_X1 u1_u5_u1_U70 (.A2( u1_u5_X_7 ) , .A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n95 ) );
  NOR2_X1 u1_u5_u1_U71 (.A1( u1_u5_X_12 ) , .A2( u1_u5_X_9 ) , .ZN( u1_u5_u1_n100 ) );
  NOR2_X1 u1_u5_u1_U72 (.A2( u1_u5_X_8 ) , .A1( u1_u5_u1_n177 ) , .ZN( u1_u5_u1_n99 ) );
  NOR2_X1 u1_u5_u1_U73 (.A2( u1_u5_X_12 ) , .ZN( u1_u5_u1_n102 ) , .A1( u1_u5_u1_n176 ) );
  NOR2_X1 u1_u5_u1_U74 (.A2( u1_u5_X_9 ) , .ZN( u1_u5_u1_n105 ) , .A1( u1_u5_u1_n168 ) );
  NAND2_X1 u1_u5_u1_U75 (.A1( u1_u5_X_10 ) , .ZN( u1_u5_u1_n160 ) , .A2( u1_u5_u1_n169 ) );
  NAND2_X1 u1_u5_u1_U76 (.A2( u1_u5_X_10 ) , .A1( u1_u5_X_11 ) , .ZN( u1_u5_u1_n152 ) );
  NAND2_X1 u1_u5_u1_U77 (.A1( u1_u5_X_11 ) , .ZN( u1_u5_u1_n128 ) , .A2( u1_u5_u1_n170 ) );
  AND2_X1 u1_u5_u1_U78 (.A2( u1_u5_X_7 ) , .A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n104 ) );
  AND2_X1 u1_u5_u1_U79 (.A1( u1_u5_X_8 ) , .ZN( u1_u5_u1_n103 ) , .A2( u1_u5_u1_n177 ) );
  NOR2_X1 u1_u5_u1_U8 (.A1( u1_u5_u1_n112 ) , .A2( u1_u5_u1_n116 ) , .ZN( u1_u5_u1_n118 ) );
  INV_X1 u1_u5_u1_U80 (.A( u1_u5_X_10 ) , .ZN( u1_u5_u1_n170 ) );
  INV_X1 u1_u5_u1_U81 (.A( u1_u5_X_9 ) , .ZN( u1_u5_u1_n176 ) );
  INV_X1 u1_u5_u1_U82 (.A( u1_u5_X_11 ) , .ZN( u1_u5_u1_n169 ) );
  INV_X1 u1_u5_u1_U83 (.A( u1_u5_X_12 ) , .ZN( u1_u5_u1_n168 ) );
  INV_X1 u1_u5_u1_U84 (.A( u1_u5_X_7 ) , .ZN( u1_u5_u1_n177 ) );
  NAND4_X1 u1_u5_u1_U85 (.ZN( u1_out5_18 ) , .A4( u1_u5_u1_n165 ) , .A3( u1_u5_u1_n166 ) , .A1( u1_u5_u1_n167 ) , .A2( u1_u5_u1_n186 ) );
  AOI22_X1 u1_u5_u1_U86 (.B2( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n147 ) , .A2( u1_u5_u1_n148 ) , .ZN( u1_u5_u1_n166 ) , .A1( u1_u5_u1_n172 ) );
  INV_X1 u1_u5_u1_U87 (.A( u1_u5_u1_n145 ) , .ZN( u1_u5_u1_n186 ) );
  OR4_X1 u1_u5_u1_U88 (.ZN( u1_out5_13 ) , .A4( u1_u5_u1_n108 ) , .A3( u1_u5_u1_n109 ) , .A2( u1_u5_u1_n110 ) , .A1( u1_u5_u1_n111 ) );
  AOI21_X1 u1_u5_u1_U89 (.ZN( u1_u5_u1_n110 ) , .A( u1_u5_u1_n116 ) , .B1( u1_u5_u1_n152 ) , .B2( u1_u5_u1_n160 ) );
  OAI21_X1 u1_u5_u1_U9 (.ZN( u1_u5_u1_n101 ) , .B1( u1_u5_u1_n141 ) , .A( u1_u5_u1_n146 ) , .B2( u1_u5_u1_n183 ) );
  AOI21_X1 u1_u5_u1_U90 (.ZN( u1_u5_u1_n111 ) , .A( u1_u5_u1_n128 ) , .B2( u1_u5_u1_n131 ) , .B1( u1_u5_u1_n135 ) );
  NAND4_X1 u1_u5_u1_U91 (.ZN( u1_out5_2 ) , .A4( u1_u5_u1_n142 ) , .A3( u1_u5_u1_n143 ) , .A2( u1_u5_u1_n144 ) , .A1( u1_u5_u1_n179 ) );
  OAI21_X1 u1_u5_u1_U92 (.B2( u1_u5_u1_n132 ) , .ZN( u1_u5_u1_n144 ) , .A( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n180 ) );
  INV_X1 u1_u5_u1_U93 (.A( u1_u5_u1_n130 ) , .ZN( u1_u5_u1_n179 ) );
  NAND4_X1 u1_u5_u1_U94 (.ZN( u1_out5_28 ) , .A4( u1_u5_u1_n124 ) , .A3( u1_u5_u1_n125 ) , .A2( u1_u5_u1_n126 ) , .A1( u1_u5_u1_n127 ) );
  OAI21_X1 u1_u5_u1_U95 (.ZN( u1_u5_u1_n127 ) , .B2( u1_u5_u1_n139 ) , .B1( u1_u5_u1_n175 ) , .A( u1_u5_u1_n183 ) );
  OAI21_X1 u1_u5_u1_U96 (.ZN( u1_u5_u1_n126 ) , .B2( u1_u5_u1_n140 ) , .A( u1_u5_u1_n146 ) , .B1( u1_u5_u1_n178 ) );
  NAND3_X1 u1_u5_u1_U97 (.A3( u1_u5_u1_n149 ) , .A2( u1_u5_u1_n150 ) , .A1( u1_u5_u1_n151 ) , .ZN( u1_u5_u1_n164 ) );
  NAND3_X1 u1_u5_u1_U98 (.A3( u1_u5_u1_n134 ) , .A2( u1_u5_u1_n135 ) , .ZN( u1_u5_u1_n136 ) , .A1( u1_u5_u1_n151 ) );
  NAND3_X1 u1_u5_u1_U99 (.A1( u1_u5_u1_n133 ) , .ZN( u1_u5_u1_n137 ) , .A2( u1_u5_u1_n154 ) , .A3( u1_u5_u1_n181 ) );
  AND3_X1 u1_u5_u7_U10 (.A3( u1_u5_u7_n110 ) , .A2( u1_u5_u7_n127 ) , .A1( u1_u5_u7_n132 ) , .ZN( u1_u5_u7_n92 ) );
  OAI21_X1 u1_u5_u7_U11 (.A( u1_u5_u7_n161 ) , .B1( u1_u5_u7_n168 ) , .B2( u1_u5_u7_n173 ) , .ZN( u1_u5_u7_n91 ) );
  AOI211_X1 u1_u5_u7_U12 (.A( u1_u5_u7_n117 ) , .ZN( u1_u5_u7_n118 ) , .C2( u1_u5_u7_n126 ) , .C1( u1_u5_u7_n177 ) , .B( u1_u5_u7_n180 ) );
  OAI22_X1 u1_u5_u7_U13 (.B1( u1_u5_u7_n115 ) , .ZN( u1_u5_u7_n117 ) , .A2( u1_u5_u7_n133 ) , .A1( u1_u5_u7_n137 ) , .B2( u1_u5_u7_n162 ) );
  INV_X1 u1_u5_u7_U14 (.A( u1_u5_u7_n116 ) , .ZN( u1_u5_u7_n180 ) );
  NOR3_X1 u1_u5_u7_U15 (.ZN( u1_u5_u7_n115 ) , .A3( u1_u5_u7_n145 ) , .A2( u1_u5_u7_n168 ) , .A1( u1_u5_u7_n169 ) );
  OAI211_X1 u1_u5_u7_U16 (.B( u1_u5_u7_n122 ) , .A( u1_u5_u7_n123 ) , .C2( u1_u5_u7_n124 ) , .ZN( u1_u5_u7_n154 ) , .C1( u1_u5_u7_n162 ) );
  AOI222_X1 u1_u5_u7_U17 (.ZN( u1_u5_u7_n122 ) , .C2( u1_u5_u7_n126 ) , .C1( u1_u5_u7_n145 ) , .B1( u1_u5_u7_n161 ) , .A2( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n170 ) , .A1( u1_u5_u7_n176 ) );
  INV_X1 u1_u5_u7_U18 (.A( u1_u5_u7_n133 ) , .ZN( u1_u5_u7_n176 ) );
  NOR3_X1 u1_u5_u7_U19 (.A2( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n135 ) , .ZN( u1_u5_u7_n136 ) , .A3( u1_u5_u7_n171 ) );
  NOR2_X1 u1_u5_u7_U20 (.A1( u1_u5_u7_n130 ) , .A2( u1_u5_u7_n134 ) , .ZN( u1_u5_u7_n153 ) );
  INV_X1 u1_u5_u7_U21 (.A( u1_u5_u7_n101 ) , .ZN( u1_u5_u7_n165 ) );
  NOR2_X1 u1_u5_u7_U22 (.ZN( u1_u5_u7_n111 ) , .A2( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n169 ) );
  AOI21_X1 u1_u5_u7_U23 (.ZN( u1_u5_u7_n104 ) , .B2( u1_u5_u7_n112 ) , .B1( u1_u5_u7_n127 ) , .A( u1_u5_u7_n164 ) );
  AOI21_X1 u1_u5_u7_U24 (.ZN( u1_u5_u7_n106 ) , .B1( u1_u5_u7_n133 ) , .B2( u1_u5_u7_n146 ) , .A( u1_u5_u7_n162 ) );
  AOI21_X1 u1_u5_u7_U25 (.A( u1_u5_u7_n101 ) , .ZN( u1_u5_u7_n107 ) , .B2( u1_u5_u7_n128 ) , .B1( u1_u5_u7_n175 ) );
  INV_X1 u1_u5_u7_U26 (.A( u1_u5_u7_n138 ) , .ZN( u1_u5_u7_n171 ) );
  INV_X1 u1_u5_u7_U27 (.A( u1_u5_u7_n131 ) , .ZN( u1_u5_u7_n177 ) );
  INV_X1 u1_u5_u7_U28 (.A( u1_u5_u7_n110 ) , .ZN( u1_u5_u7_n174 ) );
  NAND2_X1 u1_u5_u7_U29 (.A1( u1_u5_u7_n129 ) , .A2( u1_u5_u7_n132 ) , .ZN( u1_u5_u7_n149 ) );
  OAI21_X1 u1_u5_u7_U3 (.ZN( u1_u5_u7_n159 ) , .A( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n171 ) , .B1( u1_u5_u7_n174 ) );
  NAND2_X1 u1_u5_u7_U30 (.A1( u1_u5_u7_n113 ) , .A2( u1_u5_u7_n124 ) , .ZN( u1_u5_u7_n130 ) );
  INV_X1 u1_u5_u7_U31 (.A( u1_u5_u7_n112 ) , .ZN( u1_u5_u7_n173 ) );
  INV_X1 u1_u5_u7_U32 (.A( u1_u5_u7_n128 ) , .ZN( u1_u5_u7_n168 ) );
  INV_X1 u1_u5_u7_U33 (.A( u1_u5_u7_n148 ) , .ZN( u1_u5_u7_n169 ) );
  INV_X1 u1_u5_u7_U34 (.A( u1_u5_u7_n127 ) , .ZN( u1_u5_u7_n179 ) );
  NOR2_X1 u1_u5_u7_U35 (.ZN( u1_u5_u7_n101 ) , .A2( u1_u5_u7_n150 ) , .A1( u1_u5_u7_n156 ) );
  AOI211_X1 u1_u5_u7_U36 (.B( u1_u5_u7_n154 ) , .A( u1_u5_u7_n155 ) , .C1( u1_u5_u7_n156 ) , .ZN( u1_u5_u7_n157 ) , .C2( u1_u5_u7_n172 ) );
  INV_X1 u1_u5_u7_U37 (.A( u1_u5_u7_n153 ) , .ZN( u1_u5_u7_n172 ) );
  AOI211_X1 u1_u5_u7_U38 (.B( u1_u5_u7_n139 ) , .A( u1_u5_u7_n140 ) , .C2( u1_u5_u7_n141 ) , .ZN( u1_u5_u7_n142 ) , .C1( u1_u5_u7_n156 ) );
  NAND4_X1 u1_u5_u7_U39 (.A3( u1_u5_u7_n127 ) , .A2( u1_u5_u7_n128 ) , .A1( u1_u5_u7_n129 ) , .ZN( u1_u5_u7_n141 ) , .A4( u1_u5_u7_n147 ) );
  INV_X1 u1_u5_u7_U4 (.A( u1_u5_u7_n111 ) , .ZN( u1_u5_u7_n170 ) );
  AOI21_X1 u1_u5_u7_U40 (.A( u1_u5_u7_n137 ) , .B1( u1_u5_u7_n138 ) , .ZN( u1_u5_u7_n139 ) , .B2( u1_u5_u7_n146 ) );
  OAI22_X1 u1_u5_u7_U41 (.B1( u1_u5_u7_n136 ) , .ZN( u1_u5_u7_n140 ) , .A1( u1_u5_u7_n153 ) , .B2( u1_u5_u7_n162 ) , .A2( u1_u5_u7_n164 ) );
  AOI21_X1 u1_u5_u7_U42 (.ZN( u1_u5_u7_n123 ) , .B1( u1_u5_u7_n165 ) , .B2( u1_u5_u7_n177 ) , .A( u1_u5_u7_n97 ) );
  AOI21_X1 u1_u5_u7_U43 (.B2( u1_u5_u7_n113 ) , .B1( u1_u5_u7_n124 ) , .A( u1_u5_u7_n125 ) , .ZN( u1_u5_u7_n97 ) );
  INV_X1 u1_u5_u7_U44 (.A( u1_u5_u7_n125 ) , .ZN( u1_u5_u7_n161 ) );
  INV_X1 u1_u5_u7_U45 (.A( u1_u5_u7_n152 ) , .ZN( u1_u5_u7_n162 ) );
  AOI22_X1 u1_u5_u7_U46 (.A2( u1_u5_u7_n114 ) , .ZN( u1_u5_u7_n119 ) , .B1( u1_u5_u7_n130 ) , .A1( u1_u5_u7_n156 ) , .B2( u1_u5_u7_n165 ) );
  NAND2_X1 u1_u5_u7_U47 (.A2( u1_u5_u7_n112 ) , .ZN( u1_u5_u7_n114 ) , .A1( u1_u5_u7_n175 ) );
  AND2_X1 u1_u5_u7_U48 (.ZN( u1_u5_u7_n145 ) , .A2( u1_u5_u7_n98 ) , .A1( u1_u5_u7_n99 ) );
  NOR2_X1 u1_u5_u7_U49 (.ZN( u1_u5_u7_n137 ) , .A1( u1_u5_u7_n150 ) , .A2( u1_u5_u7_n161 ) );
  INV_X1 u1_u5_u7_U5 (.A( u1_u5_u7_n149 ) , .ZN( u1_u5_u7_n175 ) );
  AOI21_X1 u1_u5_u7_U50 (.ZN( u1_u5_u7_n105 ) , .B2( u1_u5_u7_n110 ) , .A( u1_u5_u7_n125 ) , .B1( u1_u5_u7_n147 ) );
  NAND2_X1 u1_u5_u7_U51 (.ZN( u1_u5_u7_n146 ) , .A1( u1_u5_u7_n95 ) , .A2( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U52 (.A2( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n147 ) , .A1( u1_u5_u7_n93 ) );
  NAND2_X1 u1_u5_u7_U53 (.A1( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n127 ) , .A2( u1_u5_u7_n99 ) );
  OR2_X1 u1_u5_u7_U54 (.ZN( u1_u5_u7_n126 ) , .A2( u1_u5_u7_n152 ) , .A1( u1_u5_u7_n156 ) );
  NAND2_X1 u1_u5_u7_U55 (.A2( u1_u5_u7_n102 ) , .A1( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n133 ) );
  NAND2_X1 u1_u5_u7_U56 (.ZN( u1_u5_u7_n112 ) , .A2( u1_u5_u7_n96 ) , .A1( u1_u5_u7_n99 ) );
  NAND2_X1 u1_u5_u7_U57 (.A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n128 ) , .A1( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U58 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n113 ) , .A2( u1_u5_u7_n93 ) );
  NAND2_X1 u1_u5_u7_U59 (.A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n124 ) , .A1( u1_u5_u7_n96 ) );
  INV_X1 u1_u5_u7_U6 (.A( u1_u5_u7_n154 ) , .ZN( u1_u5_u7_n178 ) );
  NAND2_X1 u1_u5_u7_U60 (.ZN( u1_u5_u7_n110 ) , .A1( u1_u5_u7_n95 ) , .A2( u1_u5_u7_n96 ) );
  INV_X1 u1_u5_u7_U61 (.A( u1_u5_u7_n150 ) , .ZN( u1_u5_u7_n164 ) );
  AND2_X1 u1_u5_u7_U62 (.ZN( u1_u5_u7_n134 ) , .A1( u1_u5_u7_n93 ) , .A2( u1_u5_u7_n98 ) );
  NAND2_X1 u1_u5_u7_U63 (.A1( u1_u5_u7_n100 ) , .A2( u1_u5_u7_n102 ) , .ZN( u1_u5_u7_n129 ) );
  NAND2_X1 u1_u5_u7_U64 (.A2( u1_u5_u7_n103 ) , .ZN( u1_u5_u7_n131 ) , .A1( u1_u5_u7_n95 ) );
  NAND2_X1 u1_u5_u7_U65 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n138 ) , .A2( u1_u5_u7_n99 ) );
  NAND2_X1 u1_u5_u7_U66 (.ZN( u1_u5_u7_n132 ) , .A1( u1_u5_u7_n93 ) , .A2( u1_u5_u7_n96 ) );
  NAND2_X1 u1_u5_u7_U67 (.A1( u1_u5_u7_n100 ) , .ZN( u1_u5_u7_n148 ) , .A2( u1_u5_u7_n95 ) );
  NOR2_X1 u1_u5_u7_U68 (.A2( u1_u5_X_47 ) , .ZN( u1_u5_u7_n150 ) , .A1( u1_u5_u7_n163 ) );
  NOR2_X1 u1_u5_u7_U69 (.A2( u1_u5_X_43 ) , .A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n103 ) );
  AOI211_X1 u1_u5_u7_U7 (.ZN( u1_u5_u7_n116 ) , .A( u1_u5_u7_n155 ) , .C1( u1_u5_u7_n161 ) , .C2( u1_u5_u7_n171 ) , .B( u1_u5_u7_n94 ) );
  NOR2_X1 u1_u5_u7_U70 (.A2( u1_u5_X_48 ) , .A1( u1_u5_u7_n166 ) , .ZN( u1_u5_u7_n95 ) );
  NOR2_X1 u1_u5_u7_U71 (.A2( u1_u5_X_45 ) , .A1( u1_u5_X_48 ) , .ZN( u1_u5_u7_n99 ) );
  NOR2_X1 u1_u5_u7_U72 (.A2( u1_u5_X_44 ) , .A1( u1_u5_u7_n167 ) , .ZN( u1_u5_u7_n98 ) );
  NOR2_X1 u1_u5_u7_U73 (.A2( u1_u5_X_46 ) , .A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n152 ) );
  AND2_X1 u1_u5_u7_U74 (.A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n156 ) , .A2( u1_u5_u7_n163 ) );
  NAND2_X1 u1_u5_u7_U75 (.A2( u1_u5_X_46 ) , .A1( u1_u5_X_47 ) , .ZN( u1_u5_u7_n125 ) );
  AND2_X1 u1_u5_u7_U76 (.A2( u1_u5_X_45 ) , .A1( u1_u5_X_48 ) , .ZN( u1_u5_u7_n102 ) );
  AND2_X1 u1_u5_u7_U77 (.A2( u1_u5_X_43 ) , .A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n96 ) );
  AND2_X1 u1_u5_u7_U78 (.A1( u1_u5_X_44 ) , .ZN( u1_u5_u7_n100 ) , .A2( u1_u5_u7_n167 ) );
  AND2_X1 u1_u5_u7_U79 (.A1( u1_u5_X_48 ) , .A2( u1_u5_u7_n166 ) , .ZN( u1_u5_u7_n93 ) );
  OAI222_X1 u1_u5_u7_U8 (.C2( u1_u5_u7_n101 ) , .B2( u1_u5_u7_n111 ) , .A1( u1_u5_u7_n113 ) , .C1( u1_u5_u7_n146 ) , .A2( u1_u5_u7_n162 ) , .B1( u1_u5_u7_n164 ) , .ZN( u1_u5_u7_n94 ) );
  INV_X1 u1_u5_u7_U80 (.A( u1_u5_X_46 ) , .ZN( u1_u5_u7_n163 ) );
  INV_X1 u1_u5_u7_U81 (.A( u1_u5_X_43 ) , .ZN( u1_u5_u7_n167 ) );
  INV_X1 u1_u5_u7_U82 (.A( u1_u5_X_45 ) , .ZN( u1_u5_u7_n166 ) );
  NAND4_X1 u1_u5_u7_U83 (.ZN( u1_out5_5 ) , .A4( u1_u5_u7_n108 ) , .A3( u1_u5_u7_n109 ) , .A1( u1_u5_u7_n116 ) , .A2( u1_u5_u7_n123 ) );
  AOI22_X1 u1_u5_u7_U84 (.ZN( u1_u5_u7_n109 ) , .A2( u1_u5_u7_n126 ) , .B2( u1_u5_u7_n145 ) , .B1( u1_u5_u7_n156 ) , .A1( u1_u5_u7_n171 ) );
  NOR4_X1 u1_u5_u7_U85 (.A4( u1_u5_u7_n104 ) , .A3( u1_u5_u7_n105 ) , .A2( u1_u5_u7_n106 ) , .A1( u1_u5_u7_n107 ) , .ZN( u1_u5_u7_n108 ) );
  NAND4_X1 u1_u5_u7_U86 (.ZN( u1_out5_27 ) , .A4( u1_u5_u7_n118 ) , .A3( u1_u5_u7_n119 ) , .A2( u1_u5_u7_n120 ) , .A1( u1_u5_u7_n121 ) );
  OAI21_X1 u1_u5_u7_U87 (.ZN( u1_u5_u7_n121 ) , .B2( u1_u5_u7_n145 ) , .A( u1_u5_u7_n150 ) , .B1( u1_u5_u7_n174 ) );
  OAI21_X1 u1_u5_u7_U88 (.ZN( u1_u5_u7_n120 ) , .A( u1_u5_u7_n161 ) , .B2( u1_u5_u7_n170 ) , .B1( u1_u5_u7_n179 ) );
  NAND4_X1 u1_u5_u7_U89 (.ZN( u1_out5_21 ) , .A4( u1_u5_u7_n157 ) , .A3( u1_u5_u7_n158 ) , .A2( u1_u5_u7_n159 ) , .A1( u1_u5_u7_n160 ) );
  OAI221_X1 u1_u5_u7_U9 (.C1( u1_u5_u7_n101 ) , .C2( u1_u5_u7_n147 ) , .ZN( u1_u5_u7_n155 ) , .B2( u1_u5_u7_n162 ) , .A( u1_u5_u7_n91 ) , .B1( u1_u5_u7_n92 ) );
  OAI21_X1 u1_u5_u7_U90 (.B1( u1_u5_u7_n145 ) , .ZN( u1_u5_u7_n160 ) , .A( u1_u5_u7_n161 ) , .B2( u1_u5_u7_n177 ) );
  AOI22_X1 u1_u5_u7_U91 (.B2( u1_u5_u7_n149 ) , .B1( u1_u5_u7_n150 ) , .A2( u1_u5_u7_n151 ) , .A1( u1_u5_u7_n152 ) , .ZN( u1_u5_u7_n158 ) );
  NAND4_X1 u1_u5_u7_U92 (.ZN( u1_out5_15 ) , .A4( u1_u5_u7_n142 ) , .A3( u1_u5_u7_n143 ) , .A2( u1_u5_u7_n144 ) , .A1( u1_u5_u7_n178 ) );
  OR2_X1 u1_u5_u7_U93 (.A2( u1_u5_u7_n125 ) , .A1( u1_u5_u7_n129 ) , .ZN( u1_u5_u7_n144 ) );
  AOI22_X1 u1_u5_u7_U94 (.A2( u1_u5_u7_n126 ) , .ZN( u1_u5_u7_n143 ) , .B2( u1_u5_u7_n165 ) , .B1( u1_u5_u7_n173 ) , .A1( u1_u5_u7_n174 ) );
  NAND3_X1 u1_u5_u7_U95 (.A3( u1_u5_u7_n146 ) , .A2( u1_u5_u7_n147 ) , .A1( u1_u5_u7_n148 ) , .ZN( u1_u5_u7_n151 ) );
  NAND3_X1 u1_u5_u7_U96 (.A3( u1_u5_u7_n131 ) , .A2( u1_u5_u7_n132 ) , .A1( u1_u5_u7_n133 ) , .ZN( u1_u5_u7_n135 ) );
  OAI21_X1 u1_uk_U1002 (.ZN( u1_K3_35 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1042 ) , .B2( u1_uk_n1308 ) );
  NAND2_X1 u1_uk_U1003 (.A1( u1_uk_K_r1_7 ) , .ZN( u1_uk_n1042 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U1074 (.ZN( u1_K5_42 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1082 ) , .B2( u1_uk_n1412 ) );
  NAND2_X1 u1_uk_U1075 (.A1( u1_uk_K_r3_9 ) , .ZN( u1_uk_n1082 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1115 (.ZN( u1_K5_39 ) , .A( u1_uk_n1081 ) , .B2( u1_uk_n1406 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U1116 (.A1( u1_uk_K_r3_16 ) , .ZN( u1_uk_n1081 ) , .A2( u1_uk_n242 ) );
  INV_X1 u1_uk_U1143 (.ZN( u1_K2_32 ) , .A( u1_uk_n1029 ) );
  AOI22_X1 u1_uk_U1144 (.B2( u1_uk_K_r0_15 ) , .A2( u1_uk_K_r0_36 ) , .ZN( u1_uk_n1029 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U131 (.ZN( u1_K6_47 ) , .A( u1_uk_n1100 ) , .B1( u1_uk_n142 ) , .B2( u1_uk_n1449 ) );
  NAND2_X1 u1_uk_U132 (.A1( u1_uk_K_r4_23 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1100 ) );
  INV_X1 u1_uk_U144 (.ZN( u1_K12_15 ) , .A( u1_uk_n504 ) );
  AOI22_X1 u1_uk_U145 (.B2( u1_uk_K_r10_25 ) , .A2( u1_uk_K_r10_34 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n252 ) , .ZN( u1_uk_n504 ) );
  OAI22_X1 u1_uk_U180 (.ZN( u1_K12_24 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1716 ) , .A2( u1_uk_n1745 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U189 (.ZN( u1_K12_14 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1718 ) , .A2( u1_uk_n1723 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U228 (.ZN( u1_K2_31 ) , .B2( u1_uk_n1260 ) , .A2( u1_uk_n1275 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U237 (.ZN( u1_K3_31 ) , .B2( u1_uk_n1333 ) , .A2( u1_uk_n1339 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U280 (.ZN( u1_K6_44 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1458 ) , .A2( u1_uk_n1476 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U281 (.ZN( u1_K6_48 ) , .B2( u1_uk_n1463 ) , .A2( u1_uk_n1470 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U291 (.ZN( u1_K6_8 ) , .A( u1_uk_n1103 ) , .B2( u1_uk_n1446 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U292 (.A1( u1_uk_K_r4_18 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1103 ) );
  OAI22_X1 u1_uk_U334 (.ZN( u1_K3_26 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1329 ) , .A2( u1_uk_n1345 ) , .B1( u1_uk_n202 ) );
  OAI21_X1 u1_uk_U380 (.ZN( u1_K2_33 ) , .A( u1_uk_n1030 ) , .B2( u1_uk_n1288 ) , .B1( u1_uk_n223 ) );
  NAND2_X1 u1_uk_U381 (.A1( u1_uk_K_r0_31 ) , .ZN( u1_uk_n1030 ) , .A2( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U387 (.ZN( u1_K3_28 ) , .B2( u1_uk_n1328 ) , .A2( u1_uk_n1333 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U439 (.ZN( u1_K5_37 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1395 ) , .A2( u1_uk_n1433 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U449 (.ZN( u1_K6_9 ) , .A( u1_uk_n1104 ) );
  AOI22_X1 u1_uk_U450 (.B2( u1_uk_K_r4_3 ) , .A2( u1_uk_K_r4_41 ) , .ZN( u1_uk_n1104 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U460 (.ZN( u1_K3_33 ) , .B2( u1_uk_n1322 ) , .A2( u1_uk_n1339 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n203 ) );
  OAI21_X1 u1_uk_U488 (.ZN( u1_K3_29 ) , .A( u1_uk_n1040 ) , .B2( u1_uk_n1343 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U489 (.A1( u1_uk_K_r1_44 ) , .ZN( u1_uk_n1040 ) , .A2( u1_uk_n294 ) );
  INV_X1 u1_uk_U534 (.ZN( u1_K12_17 ) , .A( u1_uk_n509 ) );
  AOI22_X1 u1_uk_U535 (.B2( u1_uk_K_r10_18 ) , .A2( u1_uk_K_r10_41 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n257 ) , .ZN( u1_uk_n509 ) );
  OAI22_X1 u1_uk_U559 (.ZN( u1_K3_36 ) , .B2( u1_uk_n1309 ) , .A2( u1_uk_n1344 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U560 (.ZN( u1_K2_36 ) , .B2( u1_uk_n1272 ) , .A2( u1_uk_n1288 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U578 (.ZN( u1_K5_38 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1394 ) , .A2( u1_uk_n1418 ) , .A1( u1_uk_n286 ) );
  INV_X1 u1_uk_U590 (.ZN( u1_K6_10 ) , .A( u1_uk_n1088 ) );
  AOI22_X1 u1_uk_U591 (.B2( u1_uk_K_r4_3 ) , .A2( u1_uk_K_r4_54 ) , .ZN( u1_uk_n1088 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U597 (.ZN( u1_K12_22 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1722 ) , .A2( u1_uk_n1732 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U630 (.ZN( u1_K2_35 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1275 ) , .A2( u1_uk_n1293 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U648 (.ZN( u1_K6_11 ) , .B2( u1_uk_n1453 ) , .A2( u1_uk_n1457 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U682 (.ZN( u1_K6_7 ) , .A( u1_uk_n1102 ) , .B2( u1_uk_n1465 ) , .B1( u1_uk_n222 ) );
  NAND2_X1 u1_uk_U683 (.A1( u1_uk_K_r4_33 ) , .ZN( u1_uk_n1102 ) , .A2( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U728 (.ZN( u1_K3_32 ) , .B2( u1_uk_n1308 ) , .A2( u1_uk_n1343 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U755 (.ZN( u1_K12_13 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1719 ) , .A2( u1_uk_n1751 ) , .B1( u1_uk_n286 ) );
  INV_X1 u1_uk_U779 (.ZN( u1_K12_21 ) , .A( u1_uk_n520 ) );
  AOI22_X1 u1_uk_U780 (.B2( u1_uk_K_r10_25 ) , .A2( u1_uk_K_r10_48 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n250 ) , .ZN( u1_uk_n520 ) );
  OAI21_X1 u1_uk_U794 (.ZN( u1_K3_27 ) , .A( u1_uk_n1039 ) , .B2( u1_uk_n1345 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U795 (.A1( u1_uk_K_r1_42 ) , .ZN( u1_uk_n1039 ) , .A2( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U82 (.ZN( u1_K3_34 ) , .B1( u1_uk_n100 ) , .A( u1_uk_n1041 ) , .B2( u1_uk_n1329 ) );
  OAI21_X1 u1_uk_U826 (.ZN( u1_K12_20 ) , .B1( u1_uk_n162 ) , .B2( u1_uk_n1722 ) , .A( u1_uk_n518 ) );
  NAND2_X1 u1_uk_U827 (.A1( u1_uk_K_r10_47 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n518 ) );
  NAND2_X1 u1_uk_U83 (.A1( u1_uk_K_r1_36 ) , .ZN( u1_uk_n1041 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U84 (.ZN( u1_K2_34 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1272 ) , .A2( u1_uk_n1303 ) , .A1( u1_uk_n217 ) );
  INV_X1 u1_uk_U86 (.ZN( u1_K12_23 ) , .A( u1_uk_n524 ) );
  OAI22_X1 u1_uk_U869 (.ZN( u1_K5_41 ) , .B2( u1_uk_n1418 ) , .A2( u1_uk_n1426 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U87 (.B2( u1_uk_K_r10_32 ) , .A2( u1_uk_K_r10_41 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n238 ) , .ZN( u1_uk_n524 ) );
  OAI22_X1 u1_uk_U888 (.ZN( u1_K6_45 ) , .B2( u1_uk_n1454 ) , .A2( u1_uk_n1459 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U889 (.ZN( u1_K3_30 ) , .B2( u1_uk_n1318 ) , .A2( u1_uk_n1344 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U895 (.ZN( u1_K6_12 ) , .A2( u1_uk_n1440 ) , .B2( u1_uk_n1456 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U918 (.ZN( u1_K3_25 ) , .B2( u1_uk_n1309 ) , .A2( u1_uk_n1313 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U931 (.ZN( u1_K12_16 ) , .A2( u1_uk_n1711 ) , .B2( u1_uk_n1723 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U938 (.ZN( u1_K12_18 ) , .A1( u1_uk_n164 ) , .A2( u1_uk_n1713 ) , .B2( u1_uk_n1751 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U950 (.ZN( u1_K6_46 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1443 ) , .B2( u1_uk_n1471 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U960 (.ZN( u1_K12_19 ) , .A1( u1_uk_n110 ) , .A2( u1_uk_n1712 ) , .B2( u1_uk_n1750 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U972 (.ZN( u1_K5_40 ) , .B2( u1_uk_n1413 ) , .A2( u1_uk_n1430 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U977 (.ZN( u1_K6_43 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1438 ) , .A2( u1_uk_n1477 ) , .B1( u1_uk_n203 ) );
  XOR2_X1 u2_U168 (.B( u2_L10_30 ) , .Z( u2_N381 ) , .A( u2_out11_30 ) );
  XOR2_X1 u2_U173 (.B( u2_L10_26 ) , .Z( u2_N377 ) , .A( u2_out11_26 ) );
  XOR2_X1 u2_U175 (.B( u2_L10_24 ) , .Z( u2_N375 ) , .A( u2_out11_24 ) );
  XOR2_X1 u2_U179 (.B( u2_L10_20 ) , .Z( u2_N371 ) , .A( u2_out11_20 ) );
  XOR2_X1 u2_U184 (.B( u2_L10_16 ) , .Z( u2_N367 ) , .A( u2_out11_16 ) );
  XOR2_X1 u2_U190 (.B( u2_L10_10 ) , .Z( u2_N361 ) , .A( u2_out11_10 ) );
  XOR2_X1 u2_U195 (.B( u2_L10_6 ) , .Z( u2_N357 ) , .A( u2_out11_6 ) );
  XOR2_X1 u2_U200 (.B( u2_L10_1 ) , .Z( u2_N352 ) , .A( u2_out11_1 ) );
  XOR2_X1 u2_U278 (.B( u2_L7_27 ) , .Z( u2_N282 ) , .A( u2_out8_27 ) );
  XOR2_X1 u2_U285 (.B( u2_L7_21 ) , .Z( u2_N276 ) , .A( u2_out8_21 ) );
  XOR2_X1 u2_U291 (.B( u2_L7_15 ) , .Z( u2_N270 ) , .A( u2_out8_15 ) );
  XOR2_X1 u2_U302 (.B( u2_L7_5 ) , .Z( u2_N260 ) , .A( u2_out8_5 ) );
  XOR2_X1 u2_u11_U33 (.B( u2_K12_24 ) , .A( u2_R10_17 ) , .Z( u2_u11_X_24 ) );
  XOR2_X1 u2_u11_U34 (.B( u2_K12_23 ) , .A( u2_R10_16 ) , .Z( u2_u11_X_23 ) );
  XOR2_X1 u2_u11_U35 (.B( u2_K12_22 ) , .A( u2_R10_15 ) , .Z( u2_u11_X_22 ) );
  XOR2_X1 u2_u11_U36 (.B( u2_K12_21 ) , .A( u2_R10_14 ) , .Z( u2_u11_X_21 ) );
  XOR2_X1 u2_u11_U37 (.B( u2_K12_20 ) , .A( u2_R10_13 ) , .Z( u2_u11_X_20 ) );
  XOR2_X1 u2_u11_U39 (.B( u2_K12_19 ) , .A( u2_R10_12 ) , .Z( u2_u11_X_19 ) );
  XOR2_X1 u2_u11_U40 (.B( u2_K12_18 ) , .A( u2_R10_13 ) , .Z( u2_u11_X_18 ) );
  XOR2_X1 u2_u11_U41 (.B( u2_K12_17 ) , .A( u2_R10_12 ) , .Z( u2_u11_X_17 ) );
  XOR2_X1 u2_u11_U42 (.B( u2_K12_16 ) , .A( u2_R10_11 ) , .Z( u2_u11_X_16 ) );
  XOR2_X1 u2_u11_U43 (.B( u2_K12_15 ) , .A( u2_R10_10 ) , .Z( u2_u11_X_15 ) );
  XOR2_X1 u2_u11_U44 (.B( u2_K12_14 ) , .A( u2_R10_9 ) , .Z( u2_u11_X_14 ) );
  XOR2_X1 u2_u11_U45 (.B( u2_K12_13 ) , .A( u2_R10_8 ) , .Z( u2_u11_X_13 ) );
  OAI22_X1 u2_u11_u2_U10 (.ZN( u2_u11_u2_n109 ) , .A2( u2_u11_u2_n113 ) , .B2( u2_u11_u2_n133 ) , .B1( u2_u11_u2_n167 ) , .A1( u2_u11_u2_n168 ) );
  NAND3_X1 u2_u11_u2_U100 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n98 ) );
  OAI22_X1 u2_u11_u2_U11 (.B1( u2_u11_u2_n151 ) , .A2( u2_u11_u2_n152 ) , .A1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n160 ) , .B2( u2_u11_u2_n168 ) );
  NOR3_X1 u2_u11_u2_U12 (.A1( u2_u11_u2_n150 ) , .ZN( u2_u11_u2_n151 ) , .A3( u2_u11_u2_n175 ) , .A2( u2_u11_u2_n188 ) );
  AOI21_X1 u2_u11_u2_U13 (.ZN( u2_u11_u2_n144 ) , .B2( u2_u11_u2_n155 ) , .A( u2_u11_u2_n172 ) , .B1( u2_u11_u2_n185 ) );
  AOI21_X1 u2_u11_u2_U14 (.B2( u2_u11_u2_n143 ) , .ZN( u2_u11_u2_n145 ) , .B1( u2_u11_u2_n152 ) , .A( u2_u11_u2_n171 ) );
  AOI21_X1 u2_u11_u2_U15 (.B2( u2_u11_u2_n120 ) , .B1( u2_u11_u2_n121 ) , .ZN( u2_u11_u2_n126 ) , .A( u2_u11_u2_n167 ) );
  INV_X1 u2_u11_u2_U16 (.A( u2_u11_u2_n156 ) , .ZN( u2_u11_u2_n171 ) );
  INV_X1 u2_u11_u2_U17 (.A( u2_u11_u2_n120 ) , .ZN( u2_u11_u2_n188 ) );
  NAND2_X1 u2_u11_u2_U18 (.A2( u2_u11_u2_n122 ) , .ZN( u2_u11_u2_n150 ) , .A1( u2_u11_u2_n152 ) );
  INV_X1 u2_u11_u2_U19 (.A( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n170 ) );
  INV_X1 u2_u11_u2_U20 (.A( u2_u11_u2_n137 ) , .ZN( u2_u11_u2_n173 ) );
  NAND2_X1 u2_u11_u2_U21 (.A1( u2_u11_u2_n132 ) , .A2( u2_u11_u2_n139 ) , .ZN( u2_u11_u2_n157 ) );
  INV_X1 u2_u11_u2_U22 (.A( u2_u11_u2_n113 ) , .ZN( u2_u11_u2_n178 ) );
  INV_X1 u2_u11_u2_U23 (.A( u2_u11_u2_n139 ) , .ZN( u2_u11_u2_n175 ) );
  INV_X1 u2_u11_u2_U24 (.A( u2_u11_u2_n155 ) , .ZN( u2_u11_u2_n181 ) );
  INV_X1 u2_u11_u2_U25 (.A( u2_u11_u2_n119 ) , .ZN( u2_u11_u2_n177 ) );
  INV_X1 u2_u11_u2_U26 (.A( u2_u11_u2_n116 ) , .ZN( u2_u11_u2_n180 ) );
  INV_X1 u2_u11_u2_U27 (.A( u2_u11_u2_n131 ) , .ZN( u2_u11_u2_n179 ) );
  INV_X1 u2_u11_u2_U28 (.A( u2_u11_u2_n154 ) , .ZN( u2_u11_u2_n176 ) );
  NAND2_X1 u2_u11_u2_U29 (.A2( u2_u11_u2_n116 ) , .A1( u2_u11_u2_n117 ) , .ZN( u2_u11_u2_n118 ) );
  NOR2_X1 u2_u11_u2_U3 (.ZN( u2_u11_u2_n121 ) , .A2( u2_u11_u2_n177 ) , .A1( u2_u11_u2_n180 ) );
  INV_X1 u2_u11_u2_U30 (.A( u2_u11_u2_n132 ) , .ZN( u2_u11_u2_n182 ) );
  INV_X1 u2_u11_u2_U31 (.A( u2_u11_u2_n158 ) , .ZN( u2_u11_u2_n183 ) );
  OAI21_X1 u2_u11_u2_U32 (.A( u2_u11_u2_n156 ) , .B1( u2_u11_u2_n157 ) , .ZN( u2_u11_u2_n158 ) , .B2( u2_u11_u2_n179 ) );
  NOR2_X1 u2_u11_u2_U33 (.ZN( u2_u11_u2_n156 ) , .A1( u2_u11_u2_n166 ) , .A2( u2_u11_u2_n169 ) );
  NOR2_X1 u2_u11_u2_U34 (.A2( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n137 ) , .A1( u2_u11_u2_n140 ) );
  NOR2_X1 u2_u11_u2_U35 (.A2( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n153 ) , .A1( u2_u11_u2_n156 ) );
  AOI211_X1 u2_u11_u2_U36 (.ZN( u2_u11_u2_n130 ) , .C1( u2_u11_u2_n138 ) , .C2( u2_u11_u2_n179 ) , .B( u2_u11_u2_n96 ) , .A( u2_u11_u2_n97 ) );
  OAI22_X1 u2_u11_u2_U37 (.B1( u2_u11_u2_n133 ) , .A2( u2_u11_u2_n137 ) , .A1( u2_u11_u2_n152 ) , .B2( u2_u11_u2_n168 ) , .ZN( u2_u11_u2_n97 ) );
  OAI221_X1 u2_u11_u2_U38 (.B1( u2_u11_u2_n113 ) , .C1( u2_u11_u2_n132 ) , .A( u2_u11_u2_n149 ) , .B2( u2_u11_u2_n171 ) , .C2( u2_u11_u2_n172 ) , .ZN( u2_u11_u2_n96 ) );
  OAI221_X1 u2_u11_u2_U39 (.A( u2_u11_u2_n115 ) , .C2( u2_u11_u2_n123 ) , .B2( u2_u11_u2_n143 ) , .B1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n163 ) , .C1( u2_u11_u2_n168 ) );
  INV_X1 u2_u11_u2_U4 (.A( u2_u11_u2_n134 ) , .ZN( u2_u11_u2_n185 ) );
  OAI21_X1 u2_u11_u2_U40 (.A( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n115 ) , .B1( u2_u11_u2_n176 ) , .B2( u2_u11_u2_n178 ) );
  OAI221_X1 u2_u11_u2_U41 (.A( u2_u11_u2_n135 ) , .B2( u2_u11_u2_n136 ) , .B1( u2_u11_u2_n137 ) , .ZN( u2_u11_u2_n162 ) , .C2( u2_u11_u2_n167 ) , .C1( u2_u11_u2_n185 ) );
  AND3_X1 u2_u11_u2_U42 (.A3( u2_u11_u2_n131 ) , .A2( u2_u11_u2_n132 ) , .A1( u2_u11_u2_n133 ) , .ZN( u2_u11_u2_n136 ) );
  AOI22_X1 u2_u11_u2_U43 (.ZN( u2_u11_u2_n135 ) , .B1( u2_u11_u2_n140 ) , .A1( u2_u11_u2_n156 ) , .B2( u2_u11_u2_n180 ) , .A2( u2_u11_u2_n188 ) );
  AOI21_X1 u2_u11_u2_U44 (.ZN( u2_u11_u2_n149 ) , .B1( u2_u11_u2_n173 ) , .B2( u2_u11_u2_n188 ) , .A( u2_u11_u2_n95 ) );
  AND3_X1 u2_u11_u2_U45 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n156 ) , .ZN( u2_u11_u2_n95 ) );
  OAI21_X1 u2_u11_u2_U46 (.A( u2_u11_u2_n101 ) , .B2( u2_u11_u2_n121 ) , .B1( u2_u11_u2_n153 ) , .ZN( u2_u11_u2_n164 ) );
  NAND2_X1 u2_u11_u2_U47 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n155 ) );
  NAND2_X1 u2_u11_u2_U48 (.A2( u2_u11_u2_n105 ) , .A1( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n143 ) );
  NAND2_X1 u2_u11_u2_U49 (.A1( u2_u11_u2_n104 ) , .A2( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n152 ) );
  INV_X1 u2_u11_u2_U5 (.A( u2_u11_u2_n150 ) , .ZN( u2_u11_u2_n184 ) );
  NAND2_X1 u2_u11_u2_U50 (.A1( u2_u11_u2_n100 ) , .A2( u2_u11_u2_n105 ) , .ZN( u2_u11_u2_n132 ) );
  INV_X1 u2_u11_u2_U51 (.A( u2_u11_u2_n140 ) , .ZN( u2_u11_u2_n168 ) );
  INV_X1 u2_u11_u2_U52 (.A( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n167 ) );
  OAI21_X1 u2_u11_u2_U53 (.A( u2_u11_u2_n141 ) , .B2( u2_u11_u2_n142 ) , .ZN( u2_u11_u2_n146 ) , .B1( u2_u11_u2_n153 ) );
  OAI21_X1 u2_u11_u2_U54 (.A( u2_u11_u2_n140 ) , .ZN( u2_u11_u2_n141 ) , .B1( u2_u11_u2_n176 ) , .B2( u2_u11_u2_n177 ) );
  NOR3_X1 u2_u11_u2_U55 (.ZN( u2_u11_u2_n142 ) , .A3( u2_u11_u2_n175 ) , .A2( u2_u11_u2_n178 ) , .A1( u2_u11_u2_n181 ) );
  NAND2_X1 u2_u11_u2_U56 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n113 ) );
  NAND2_X1 u2_u11_u2_U57 (.A1( u2_u11_u2_n106 ) , .A2( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n131 ) );
  NAND2_X1 u2_u11_u2_U58 (.A1( u2_u11_u2_n103 ) , .A2( u2_u11_u2_n107 ) , .ZN( u2_u11_u2_n139 ) );
  NAND2_X1 u2_u11_u2_U59 (.A1( u2_u11_u2_n103 ) , .A2( u2_u11_u2_n105 ) , .ZN( u2_u11_u2_n133 ) );
  NOR4_X1 u2_u11_u2_U6 (.A4( u2_u11_u2_n124 ) , .A3( u2_u11_u2_n125 ) , .A2( u2_u11_u2_n126 ) , .A1( u2_u11_u2_n127 ) , .ZN( u2_u11_u2_n128 ) );
  NAND2_X1 u2_u11_u2_U60 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n103 ) , .ZN( u2_u11_u2_n154 ) );
  NAND2_X1 u2_u11_u2_U61 (.A2( u2_u11_u2_n103 ) , .A1( u2_u11_u2_n104 ) , .ZN( u2_u11_u2_n119 ) );
  NAND2_X1 u2_u11_u2_U62 (.A2( u2_u11_u2_n107 ) , .A1( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n123 ) );
  NAND2_X1 u2_u11_u2_U63 (.A1( u2_u11_u2_n104 ) , .A2( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n122 ) );
  INV_X1 u2_u11_u2_U64 (.A( u2_u11_u2_n114 ) , .ZN( u2_u11_u2_n172 ) );
  NAND2_X1 u2_u11_u2_U65 (.A2( u2_u11_u2_n100 ) , .A1( u2_u11_u2_n102 ) , .ZN( u2_u11_u2_n116 ) );
  NAND2_X1 u2_u11_u2_U66 (.A1( u2_u11_u2_n102 ) , .A2( u2_u11_u2_n108 ) , .ZN( u2_u11_u2_n120 ) );
  NAND2_X1 u2_u11_u2_U67 (.A2( u2_u11_u2_n105 ) , .A1( u2_u11_u2_n106 ) , .ZN( u2_u11_u2_n117 ) );
  INV_X1 u2_u11_u2_U68 (.ZN( u2_u11_u2_n187 ) , .A( u2_u11_u2_n99 ) );
  OAI21_X1 u2_u11_u2_U69 (.B1( u2_u11_u2_n137 ) , .B2( u2_u11_u2_n143 ) , .A( u2_u11_u2_n98 ) , .ZN( u2_u11_u2_n99 ) );
  AOI21_X1 u2_u11_u2_U7 (.ZN( u2_u11_u2_n124 ) , .B1( u2_u11_u2_n131 ) , .B2( u2_u11_u2_n143 ) , .A( u2_u11_u2_n172 ) );
  NOR2_X1 u2_u11_u2_U70 (.A2( u2_u11_X_16 ) , .ZN( u2_u11_u2_n140 ) , .A1( u2_u11_u2_n166 ) );
  NOR2_X1 u2_u11_u2_U71 (.A2( u2_u11_X_13 ) , .A1( u2_u11_X_14 ) , .ZN( u2_u11_u2_n100 ) );
  NOR2_X1 u2_u11_u2_U72 (.A2( u2_u11_X_16 ) , .A1( u2_u11_X_17 ) , .ZN( u2_u11_u2_n138 ) );
  NOR2_X1 u2_u11_u2_U73 (.A2( u2_u11_X_15 ) , .A1( u2_u11_X_18 ) , .ZN( u2_u11_u2_n104 ) );
  NOR2_X1 u2_u11_u2_U74 (.A2( u2_u11_X_14 ) , .ZN( u2_u11_u2_n103 ) , .A1( u2_u11_u2_n174 ) );
  NOR2_X1 u2_u11_u2_U75 (.A2( u2_u11_X_15 ) , .ZN( u2_u11_u2_n102 ) , .A1( u2_u11_u2_n165 ) );
  NOR2_X1 u2_u11_u2_U76 (.A2( u2_u11_X_17 ) , .ZN( u2_u11_u2_n114 ) , .A1( u2_u11_u2_n169 ) );
  AND2_X1 u2_u11_u2_U77 (.A1( u2_u11_X_15 ) , .ZN( u2_u11_u2_n105 ) , .A2( u2_u11_u2_n165 ) );
  AND2_X1 u2_u11_u2_U78 (.A2( u2_u11_X_15 ) , .A1( u2_u11_X_18 ) , .ZN( u2_u11_u2_n107 ) );
  AND2_X1 u2_u11_u2_U79 (.A1( u2_u11_X_14 ) , .ZN( u2_u11_u2_n106 ) , .A2( u2_u11_u2_n174 ) );
  AOI21_X1 u2_u11_u2_U8 (.B2( u2_u11_u2_n119 ) , .ZN( u2_u11_u2_n127 ) , .A( u2_u11_u2_n137 ) , .B1( u2_u11_u2_n155 ) );
  AND2_X1 u2_u11_u2_U80 (.A1( u2_u11_X_13 ) , .A2( u2_u11_X_14 ) , .ZN( u2_u11_u2_n108 ) );
  INV_X1 u2_u11_u2_U81 (.A( u2_u11_X_16 ) , .ZN( u2_u11_u2_n169 ) );
  INV_X1 u2_u11_u2_U82 (.A( u2_u11_X_17 ) , .ZN( u2_u11_u2_n166 ) );
  INV_X1 u2_u11_u2_U83 (.A( u2_u11_X_13 ) , .ZN( u2_u11_u2_n174 ) );
  INV_X1 u2_u11_u2_U84 (.A( u2_u11_X_18 ) , .ZN( u2_u11_u2_n165 ) );
  NAND4_X1 u2_u11_u2_U85 (.ZN( u2_out11_30 ) , .A4( u2_u11_u2_n147 ) , .A3( u2_u11_u2_n148 ) , .A2( u2_u11_u2_n149 ) , .A1( u2_u11_u2_n187 ) );
  NOR3_X1 u2_u11_u2_U86 (.A3( u2_u11_u2_n144 ) , .A2( u2_u11_u2_n145 ) , .A1( u2_u11_u2_n146 ) , .ZN( u2_u11_u2_n147 ) );
  AOI21_X1 u2_u11_u2_U87 (.B2( u2_u11_u2_n138 ) , .ZN( u2_u11_u2_n148 ) , .A( u2_u11_u2_n162 ) , .B1( u2_u11_u2_n182 ) );
  NAND4_X1 u2_u11_u2_U88 (.ZN( u2_out11_24 ) , .A4( u2_u11_u2_n111 ) , .A3( u2_u11_u2_n112 ) , .A1( u2_u11_u2_n130 ) , .A2( u2_u11_u2_n187 ) );
  AOI221_X1 u2_u11_u2_U89 (.A( u2_u11_u2_n109 ) , .B1( u2_u11_u2_n110 ) , .ZN( u2_u11_u2_n111 ) , .C1( u2_u11_u2_n134 ) , .C2( u2_u11_u2_n170 ) , .B2( u2_u11_u2_n173 ) );
  AOI21_X1 u2_u11_u2_U9 (.B2( u2_u11_u2_n123 ) , .ZN( u2_u11_u2_n125 ) , .A( u2_u11_u2_n171 ) , .B1( u2_u11_u2_n184 ) );
  AOI21_X1 u2_u11_u2_U90 (.ZN( u2_u11_u2_n112 ) , .B2( u2_u11_u2_n156 ) , .A( u2_u11_u2_n164 ) , .B1( u2_u11_u2_n181 ) );
  NAND4_X1 u2_u11_u2_U91 (.ZN( u2_out11_16 ) , .A4( u2_u11_u2_n128 ) , .A3( u2_u11_u2_n129 ) , .A1( u2_u11_u2_n130 ) , .A2( u2_u11_u2_n186 ) );
  AOI22_X1 u2_u11_u2_U92 (.A2( u2_u11_u2_n118 ) , .ZN( u2_u11_u2_n129 ) , .A1( u2_u11_u2_n140 ) , .B1( u2_u11_u2_n157 ) , .B2( u2_u11_u2_n170 ) );
  INV_X1 u2_u11_u2_U93 (.A( u2_u11_u2_n163 ) , .ZN( u2_u11_u2_n186 ) );
  OR4_X1 u2_u11_u2_U94 (.ZN( u2_out11_6 ) , .A4( u2_u11_u2_n161 ) , .A3( u2_u11_u2_n162 ) , .A2( u2_u11_u2_n163 ) , .A1( u2_u11_u2_n164 ) );
  OR3_X1 u2_u11_u2_U95 (.A2( u2_u11_u2_n159 ) , .A1( u2_u11_u2_n160 ) , .ZN( u2_u11_u2_n161 ) , .A3( u2_u11_u2_n183 ) );
  AOI21_X1 u2_u11_u2_U96 (.B2( u2_u11_u2_n154 ) , .B1( u2_u11_u2_n155 ) , .ZN( u2_u11_u2_n159 ) , .A( u2_u11_u2_n167 ) );
  NAND3_X1 u2_u11_u2_U97 (.A2( u2_u11_u2_n117 ) , .A1( u2_u11_u2_n122 ) , .A3( u2_u11_u2_n123 ) , .ZN( u2_u11_u2_n134 ) );
  NAND3_X1 u2_u11_u2_U98 (.ZN( u2_u11_u2_n110 ) , .A2( u2_u11_u2_n131 ) , .A3( u2_u11_u2_n139 ) , .A1( u2_u11_u2_n154 ) );
  NAND3_X1 u2_u11_u2_U99 (.A2( u2_u11_u2_n100 ) , .ZN( u2_u11_u2_n101 ) , .A1( u2_u11_u2_n104 ) , .A3( u2_u11_u2_n114 ) );
  OAI211_X1 u2_u11_u3_U10 (.B( u2_u11_u3_n106 ) , .ZN( u2_u11_u3_n119 ) , .C2( u2_u11_u3_n128 ) , .C1( u2_u11_u3_n167 ) , .A( u2_u11_u3_n181 ) );
  INV_X1 u2_u11_u3_U11 (.ZN( u2_u11_u3_n181 ) , .A( u2_u11_u3_n98 ) );
  AOI221_X1 u2_u11_u3_U12 (.C1( u2_u11_u3_n105 ) , .ZN( u2_u11_u3_n106 ) , .A( u2_u11_u3_n131 ) , .B2( u2_u11_u3_n132 ) , .C2( u2_u11_u3_n133 ) , .B1( u2_u11_u3_n169 ) );
  OAI22_X1 u2_u11_u3_U13 (.B1( u2_u11_u3_n113 ) , .A2( u2_u11_u3_n135 ) , .A1( u2_u11_u3_n150 ) , .B2( u2_u11_u3_n164 ) , .ZN( u2_u11_u3_n98 ) );
  AOI22_X1 u2_u11_u3_U14 (.B1( u2_u11_u3_n115 ) , .A2( u2_u11_u3_n116 ) , .ZN( u2_u11_u3_n123 ) , .B2( u2_u11_u3_n133 ) , .A1( u2_u11_u3_n169 ) );
  NAND2_X1 u2_u11_u3_U15 (.ZN( u2_u11_u3_n116 ) , .A2( u2_u11_u3_n151 ) , .A1( u2_u11_u3_n182 ) );
  NOR2_X1 u2_u11_u3_U16 (.ZN( u2_u11_u3_n126 ) , .A2( u2_u11_u3_n150 ) , .A1( u2_u11_u3_n164 ) );
  AOI21_X1 u2_u11_u3_U17 (.ZN( u2_u11_u3_n112 ) , .B2( u2_u11_u3_n146 ) , .B1( u2_u11_u3_n155 ) , .A( u2_u11_u3_n167 ) );
  NAND2_X1 u2_u11_u3_U18 (.A1( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n142 ) , .A2( u2_u11_u3_n164 ) );
  NAND2_X1 u2_u11_u3_U19 (.ZN( u2_u11_u3_n132 ) , .A2( u2_u11_u3_n152 ) , .A1( u2_u11_u3_n156 ) );
  INV_X1 u2_u11_u3_U20 (.A( u2_u11_u3_n133 ) , .ZN( u2_u11_u3_n165 ) );
  AND2_X1 u2_u11_u3_U21 (.A2( u2_u11_u3_n113 ) , .A1( u2_u11_u3_n114 ) , .ZN( u2_u11_u3_n151 ) );
  INV_X1 u2_u11_u3_U22 (.A( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n170 ) );
  NAND2_X1 u2_u11_u3_U23 (.A1( u2_u11_u3_n107 ) , .A2( u2_u11_u3_n108 ) , .ZN( u2_u11_u3_n140 ) );
  NAND2_X1 u2_u11_u3_U24 (.ZN( u2_u11_u3_n117 ) , .A1( u2_u11_u3_n124 ) , .A2( u2_u11_u3_n148 ) );
  NAND2_X1 u2_u11_u3_U25 (.ZN( u2_u11_u3_n143 ) , .A1( u2_u11_u3_n165 ) , .A2( u2_u11_u3_n167 ) );
  INV_X1 u2_u11_u3_U26 (.A( u2_u11_u3_n130 ) , .ZN( u2_u11_u3_n177 ) );
  INV_X1 u2_u11_u3_U27 (.A( u2_u11_u3_n128 ) , .ZN( u2_u11_u3_n176 ) );
  NAND2_X1 u2_u11_u3_U28 (.ZN( u2_u11_u3_n105 ) , .A2( u2_u11_u3_n130 ) , .A1( u2_u11_u3_n155 ) );
  INV_X1 u2_u11_u3_U29 (.A( u2_u11_u3_n155 ) , .ZN( u2_u11_u3_n174 ) );
  INV_X1 u2_u11_u3_U3 (.A( u2_u11_u3_n140 ) , .ZN( u2_u11_u3_n182 ) );
  INV_X1 u2_u11_u3_U30 (.A( u2_u11_u3_n139 ) , .ZN( u2_u11_u3_n185 ) );
  NOR2_X1 u2_u11_u3_U31 (.ZN( u2_u11_u3_n135 ) , .A2( u2_u11_u3_n141 ) , .A1( u2_u11_u3_n169 ) );
  OAI222_X1 u2_u11_u3_U32 (.C2( u2_u11_u3_n107 ) , .A2( u2_u11_u3_n108 ) , .B1( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n138 ) , .B2( u2_u11_u3_n146 ) , .C1( u2_u11_u3_n154 ) , .A1( u2_u11_u3_n164 ) );
  NOR4_X1 u2_u11_u3_U33 (.A4( u2_u11_u3_n157 ) , .A3( u2_u11_u3_n158 ) , .A2( u2_u11_u3_n159 ) , .A1( u2_u11_u3_n160 ) , .ZN( u2_u11_u3_n161 ) );
  AOI21_X1 u2_u11_u3_U34 (.B2( u2_u11_u3_n152 ) , .B1( u2_u11_u3_n153 ) , .ZN( u2_u11_u3_n158 ) , .A( u2_u11_u3_n164 ) );
  AOI21_X1 u2_u11_u3_U35 (.A( u2_u11_u3_n154 ) , .B2( u2_u11_u3_n155 ) , .B1( u2_u11_u3_n156 ) , .ZN( u2_u11_u3_n157 ) );
  AOI21_X1 u2_u11_u3_U36 (.A( u2_u11_u3_n149 ) , .B2( u2_u11_u3_n150 ) , .B1( u2_u11_u3_n151 ) , .ZN( u2_u11_u3_n159 ) );
  AOI211_X1 u2_u11_u3_U37 (.ZN( u2_u11_u3_n109 ) , .A( u2_u11_u3_n119 ) , .C2( u2_u11_u3_n129 ) , .B( u2_u11_u3_n138 ) , .C1( u2_u11_u3_n141 ) );
  AOI211_X1 u2_u11_u3_U38 (.B( u2_u11_u3_n119 ) , .A( u2_u11_u3_n120 ) , .C2( u2_u11_u3_n121 ) , .ZN( u2_u11_u3_n122 ) , .C1( u2_u11_u3_n179 ) );
  INV_X1 u2_u11_u3_U39 (.A( u2_u11_u3_n156 ) , .ZN( u2_u11_u3_n179 ) );
  INV_X1 u2_u11_u3_U4 (.A( u2_u11_u3_n129 ) , .ZN( u2_u11_u3_n183 ) );
  OAI22_X1 u2_u11_u3_U40 (.B1( u2_u11_u3_n118 ) , .ZN( u2_u11_u3_n120 ) , .A1( u2_u11_u3_n135 ) , .B2( u2_u11_u3_n154 ) , .A2( u2_u11_u3_n178 ) );
  AND3_X1 u2_u11_u3_U41 (.ZN( u2_u11_u3_n118 ) , .A2( u2_u11_u3_n124 ) , .A1( u2_u11_u3_n144 ) , .A3( u2_u11_u3_n152 ) );
  INV_X1 u2_u11_u3_U42 (.A( u2_u11_u3_n121 ) , .ZN( u2_u11_u3_n164 ) );
  NAND2_X1 u2_u11_u3_U43 (.ZN( u2_u11_u3_n133 ) , .A1( u2_u11_u3_n154 ) , .A2( u2_u11_u3_n164 ) );
  NOR2_X1 u2_u11_u3_U44 (.A1( u2_u11_u3_n113 ) , .ZN( u2_u11_u3_n131 ) , .A2( u2_u11_u3_n154 ) );
  NAND2_X1 u2_u11_u3_U45 (.A1( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n150 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U46 (.A2( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n155 ) , .A1( u2_u11_u3_n97 ) );
  OAI211_X1 u2_u11_u3_U47 (.B( u2_u11_u3_n127 ) , .ZN( u2_u11_u3_n139 ) , .C1( u2_u11_u3_n150 ) , .C2( u2_u11_u3_n154 ) , .A( u2_u11_u3_n184 ) );
  INV_X1 u2_u11_u3_U48 (.A( u2_u11_u3_n125 ) , .ZN( u2_u11_u3_n184 ) );
  AOI221_X1 u2_u11_u3_U49 (.A( u2_u11_u3_n126 ) , .ZN( u2_u11_u3_n127 ) , .C2( u2_u11_u3_n132 ) , .C1( u2_u11_u3_n169 ) , .B2( u2_u11_u3_n170 ) , .B1( u2_u11_u3_n174 ) );
  INV_X1 u2_u11_u3_U5 (.A( u2_u11_u3_n117 ) , .ZN( u2_u11_u3_n178 ) );
  OAI22_X1 u2_u11_u3_U50 (.A1( u2_u11_u3_n124 ) , .ZN( u2_u11_u3_n125 ) , .B2( u2_u11_u3_n145 ) , .A2( u2_u11_u3_n165 ) , .B1( u2_u11_u3_n167 ) );
  INV_X1 u2_u11_u3_U51 (.A( u2_u11_u3_n141 ) , .ZN( u2_u11_u3_n167 ) );
  AOI21_X1 u2_u11_u3_U52 (.B2( u2_u11_u3_n114 ) , .B1( u2_u11_u3_n146 ) , .A( u2_u11_u3_n154 ) , .ZN( u2_u11_u3_n94 ) );
  AOI21_X1 u2_u11_u3_U53 (.ZN( u2_u11_u3_n110 ) , .B2( u2_u11_u3_n142 ) , .B1( u2_u11_u3_n186 ) , .A( u2_u11_u3_n95 ) );
  INV_X1 u2_u11_u3_U54 (.A( u2_u11_u3_n145 ) , .ZN( u2_u11_u3_n186 ) );
  AOI21_X1 u2_u11_u3_U55 (.B1( u2_u11_u3_n124 ) , .A( u2_u11_u3_n149 ) , .B2( u2_u11_u3_n155 ) , .ZN( u2_u11_u3_n95 ) );
  INV_X1 u2_u11_u3_U56 (.A( u2_u11_u3_n149 ) , .ZN( u2_u11_u3_n169 ) );
  NAND2_X1 u2_u11_u3_U57 (.ZN( u2_u11_u3_n124 ) , .A1( u2_u11_u3_n96 ) , .A2( u2_u11_u3_n97 ) );
  NAND2_X1 u2_u11_u3_U58 (.A2( u2_u11_u3_n100 ) , .ZN( u2_u11_u3_n146 ) , .A1( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U59 (.A1( u2_u11_u3_n101 ) , .ZN( u2_u11_u3_n145 ) , .A2( u2_u11_u3_n99 ) );
  AOI221_X1 u2_u11_u3_U6 (.A( u2_u11_u3_n131 ) , .C2( u2_u11_u3_n132 ) , .C1( u2_u11_u3_n133 ) , .ZN( u2_u11_u3_n134 ) , .B1( u2_u11_u3_n143 ) , .B2( u2_u11_u3_n177 ) );
  NAND2_X1 u2_u11_u3_U60 (.A1( u2_u11_u3_n100 ) , .ZN( u2_u11_u3_n156 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U61 (.A2( u2_u11_u3_n101 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n148 ) );
  NAND2_X1 u2_u11_u3_U62 (.A1( u2_u11_u3_n100 ) , .A2( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n128 ) );
  NAND2_X1 u2_u11_u3_U63 (.A2( u2_u11_u3_n101 ) , .A1( u2_u11_u3_n102 ) , .ZN( u2_u11_u3_n152 ) );
  NAND2_X1 u2_u11_u3_U64 (.A2( u2_u11_u3_n101 ) , .ZN( u2_u11_u3_n114 ) , .A1( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U65 (.ZN( u2_u11_u3_n107 ) , .A1( u2_u11_u3_n97 ) , .A2( u2_u11_u3_n99 ) );
  NAND2_X1 u2_u11_u3_U66 (.A2( u2_u11_u3_n100 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n113 ) );
  NAND2_X1 u2_u11_u3_U67 (.A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n153 ) , .A2( u2_u11_u3_n97 ) );
  NAND2_X1 u2_u11_u3_U68 (.A2( u2_u11_u3_n103 ) , .A1( u2_u11_u3_n104 ) , .ZN( u2_u11_u3_n130 ) );
  NAND2_X1 u2_u11_u3_U69 (.A2( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n144 ) , .A1( u2_u11_u3_n96 ) );
  OAI22_X1 u2_u11_u3_U7 (.B2( u2_u11_u3_n147 ) , .A2( u2_u11_u3_n148 ) , .ZN( u2_u11_u3_n160 ) , .B1( u2_u11_u3_n165 ) , .A1( u2_u11_u3_n168 ) );
  NAND2_X1 u2_u11_u3_U70 (.A1( u2_u11_u3_n102 ) , .A2( u2_u11_u3_n103 ) , .ZN( u2_u11_u3_n108 ) );
  NOR2_X1 u2_u11_u3_U71 (.A2( u2_u11_X_19 ) , .A1( u2_u11_X_20 ) , .ZN( u2_u11_u3_n99 ) );
  NOR2_X1 u2_u11_u3_U72 (.A2( u2_u11_X_21 ) , .A1( u2_u11_X_24 ) , .ZN( u2_u11_u3_n103 ) );
  NOR2_X1 u2_u11_u3_U73 (.A2( u2_u11_X_24 ) , .A1( u2_u11_u3_n171 ) , .ZN( u2_u11_u3_n97 ) );
  NOR2_X1 u2_u11_u3_U74 (.A2( u2_u11_X_23 ) , .ZN( u2_u11_u3_n141 ) , .A1( u2_u11_u3_n166 ) );
  NOR2_X1 u2_u11_u3_U75 (.A2( u2_u11_X_19 ) , .A1( u2_u11_u3_n172 ) , .ZN( u2_u11_u3_n96 ) );
  NAND2_X1 u2_u11_u3_U76 (.A1( u2_u11_X_22 ) , .A2( u2_u11_X_23 ) , .ZN( u2_u11_u3_n154 ) );
  NAND2_X1 u2_u11_u3_U77 (.A1( u2_u11_X_23 ) , .ZN( u2_u11_u3_n149 ) , .A2( u2_u11_u3_n166 ) );
  NOR2_X1 u2_u11_u3_U78 (.A2( u2_u11_X_22 ) , .A1( u2_u11_X_23 ) , .ZN( u2_u11_u3_n121 ) );
  AND2_X1 u2_u11_u3_U79 (.A1( u2_u11_X_24 ) , .ZN( u2_u11_u3_n101 ) , .A2( u2_u11_u3_n171 ) );
  AND3_X1 u2_u11_u3_U8 (.A3( u2_u11_u3_n144 ) , .A2( u2_u11_u3_n145 ) , .A1( u2_u11_u3_n146 ) , .ZN( u2_u11_u3_n147 ) );
  AND2_X1 u2_u11_u3_U80 (.A1( u2_u11_X_19 ) , .ZN( u2_u11_u3_n102 ) , .A2( u2_u11_u3_n172 ) );
  AND2_X1 u2_u11_u3_U81 (.A1( u2_u11_X_21 ) , .A2( u2_u11_X_24 ) , .ZN( u2_u11_u3_n100 ) );
  AND2_X1 u2_u11_u3_U82 (.A2( u2_u11_X_19 ) , .A1( u2_u11_X_20 ) , .ZN( u2_u11_u3_n104 ) );
  INV_X1 u2_u11_u3_U83 (.A( u2_u11_X_22 ) , .ZN( u2_u11_u3_n166 ) );
  INV_X1 u2_u11_u3_U84 (.A( u2_u11_X_21 ) , .ZN( u2_u11_u3_n171 ) );
  INV_X1 u2_u11_u3_U85 (.A( u2_u11_X_20 ) , .ZN( u2_u11_u3_n172 ) );
  NAND4_X1 u2_u11_u3_U86 (.ZN( u2_out11_26 ) , .A4( u2_u11_u3_n109 ) , .A3( u2_u11_u3_n110 ) , .A2( u2_u11_u3_n111 ) , .A1( u2_u11_u3_n173 ) );
  INV_X1 u2_u11_u3_U87 (.ZN( u2_u11_u3_n173 ) , .A( u2_u11_u3_n94 ) );
  OAI21_X1 u2_u11_u3_U88 (.ZN( u2_u11_u3_n111 ) , .B2( u2_u11_u3_n117 ) , .A( u2_u11_u3_n133 ) , .B1( u2_u11_u3_n176 ) );
  NAND4_X1 u2_u11_u3_U89 (.ZN( u2_out11_20 ) , .A4( u2_u11_u3_n122 ) , .A3( u2_u11_u3_n123 ) , .A1( u2_u11_u3_n175 ) , .A2( u2_u11_u3_n180 ) );
  INV_X1 u2_u11_u3_U9 (.A( u2_u11_u3_n143 ) , .ZN( u2_u11_u3_n168 ) );
  INV_X1 u2_u11_u3_U90 (.A( u2_u11_u3_n126 ) , .ZN( u2_u11_u3_n180 ) );
  INV_X1 u2_u11_u3_U91 (.A( u2_u11_u3_n112 ) , .ZN( u2_u11_u3_n175 ) );
  NAND4_X1 u2_u11_u3_U92 (.ZN( u2_out11_1 ) , .A4( u2_u11_u3_n161 ) , .A3( u2_u11_u3_n162 ) , .A2( u2_u11_u3_n163 ) , .A1( u2_u11_u3_n185 ) );
  NAND2_X1 u2_u11_u3_U93 (.ZN( u2_u11_u3_n163 ) , .A2( u2_u11_u3_n170 ) , .A1( u2_u11_u3_n176 ) );
  AOI22_X1 u2_u11_u3_U94 (.B2( u2_u11_u3_n140 ) , .B1( u2_u11_u3_n141 ) , .A2( u2_u11_u3_n142 ) , .ZN( u2_u11_u3_n162 ) , .A1( u2_u11_u3_n177 ) );
  OAI222_X1 u2_u11_u3_U95 (.C1( u2_u11_u3_n128 ) , .ZN( u2_u11_u3_n137 ) , .B1( u2_u11_u3_n148 ) , .A2( u2_u11_u3_n150 ) , .B2( u2_u11_u3_n154 ) , .C2( u2_u11_u3_n164 ) , .A1( u2_u11_u3_n167 ) );
  OR4_X1 u2_u11_u3_U96 (.ZN( u2_out11_10 ) , .A4( u2_u11_u3_n136 ) , .A3( u2_u11_u3_n137 ) , .A1( u2_u11_u3_n138 ) , .A2( u2_u11_u3_n139 ) );
  OAI221_X1 u2_u11_u3_U97 (.A( u2_u11_u3_n134 ) , .B2( u2_u11_u3_n135 ) , .ZN( u2_u11_u3_n136 ) , .C1( u2_u11_u3_n149 ) , .B1( u2_u11_u3_n151 ) , .C2( u2_u11_u3_n183 ) );
  NAND3_X1 u2_u11_u3_U98 (.A1( u2_u11_u3_n114 ) , .ZN( u2_u11_u3_n115 ) , .A2( u2_u11_u3_n145 ) , .A3( u2_u11_u3_n153 ) );
  NAND3_X1 u2_u11_u3_U99 (.ZN( u2_u11_u3_n129 ) , .A2( u2_u11_u3_n144 ) , .A1( u2_u11_u3_n153 ) , .A3( u2_u11_u3_n182 ) );
  XOR2_X1 u2_u8_U10 (.B( u2_K9_45 ) , .A( u2_R7_30 ) , .Z( u2_u8_X_45 ) );
  XOR2_X1 u2_u8_U11 (.B( u2_K9_44 ) , .A( u2_R7_29 ) , .Z( u2_u8_X_44 ) );
  XOR2_X1 u2_u8_U12 (.B( u2_K9_43 ) , .A( u2_R7_28 ) , .Z( u2_u8_X_43 ) );
  XOR2_X1 u2_u8_U7 (.B( u2_K9_48 ) , .A( u2_R7_1 ) , .Z( u2_u8_X_48 ) );
  XOR2_X1 u2_u8_U8 (.B( u2_K9_47 ) , .A( u2_R7_32 ) , .Z( u2_u8_X_47 ) );
  XOR2_X1 u2_u8_U9 (.B( u2_K9_46 ) , .A( u2_R7_31 ) , .Z( u2_u8_X_46 ) );
  AND3_X1 u2_u8_u7_U10 (.A3( u2_u8_u7_n110 ) , .A2( u2_u8_u7_n127 ) , .A1( u2_u8_u7_n132 ) , .ZN( u2_u8_u7_n92 ) );
  OAI21_X1 u2_u8_u7_U11 (.A( u2_u8_u7_n161 ) , .B1( u2_u8_u7_n168 ) , .B2( u2_u8_u7_n173 ) , .ZN( u2_u8_u7_n91 ) );
  AOI211_X1 u2_u8_u7_U12 (.A( u2_u8_u7_n117 ) , .ZN( u2_u8_u7_n118 ) , .C2( u2_u8_u7_n126 ) , .C1( u2_u8_u7_n177 ) , .B( u2_u8_u7_n180 ) );
  OAI22_X1 u2_u8_u7_U13 (.B1( u2_u8_u7_n115 ) , .ZN( u2_u8_u7_n117 ) , .A2( u2_u8_u7_n133 ) , .A1( u2_u8_u7_n137 ) , .B2( u2_u8_u7_n162 ) );
  INV_X1 u2_u8_u7_U14 (.A( u2_u8_u7_n116 ) , .ZN( u2_u8_u7_n180 ) );
  NOR3_X1 u2_u8_u7_U15 (.ZN( u2_u8_u7_n115 ) , .A3( u2_u8_u7_n145 ) , .A2( u2_u8_u7_n168 ) , .A1( u2_u8_u7_n169 ) );
  OAI211_X1 u2_u8_u7_U16 (.B( u2_u8_u7_n122 ) , .A( u2_u8_u7_n123 ) , .C2( u2_u8_u7_n124 ) , .ZN( u2_u8_u7_n154 ) , .C1( u2_u8_u7_n162 ) );
  AOI222_X1 u2_u8_u7_U17 (.ZN( u2_u8_u7_n122 ) , .C2( u2_u8_u7_n126 ) , .C1( u2_u8_u7_n145 ) , .B1( u2_u8_u7_n161 ) , .A2( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n170 ) , .A1( u2_u8_u7_n176 ) );
  INV_X1 u2_u8_u7_U18 (.A( u2_u8_u7_n133 ) , .ZN( u2_u8_u7_n176 ) );
  NOR3_X1 u2_u8_u7_U19 (.A2( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n135 ) , .ZN( u2_u8_u7_n136 ) , .A3( u2_u8_u7_n171 ) );
  NOR2_X1 u2_u8_u7_U20 (.A1( u2_u8_u7_n130 ) , .A2( u2_u8_u7_n134 ) , .ZN( u2_u8_u7_n153 ) );
  INV_X1 u2_u8_u7_U21 (.A( u2_u8_u7_n101 ) , .ZN( u2_u8_u7_n165 ) );
  NOR2_X1 u2_u8_u7_U22 (.ZN( u2_u8_u7_n111 ) , .A2( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n169 ) );
  AOI21_X1 u2_u8_u7_U23 (.ZN( u2_u8_u7_n104 ) , .B2( u2_u8_u7_n112 ) , .B1( u2_u8_u7_n127 ) , .A( u2_u8_u7_n164 ) );
  AOI21_X1 u2_u8_u7_U24 (.ZN( u2_u8_u7_n106 ) , .B1( u2_u8_u7_n133 ) , .B2( u2_u8_u7_n146 ) , .A( u2_u8_u7_n162 ) );
  AOI21_X1 u2_u8_u7_U25 (.A( u2_u8_u7_n101 ) , .ZN( u2_u8_u7_n107 ) , .B2( u2_u8_u7_n128 ) , .B1( u2_u8_u7_n175 ) );
  INV_X1 u2_u8_u7_U26 (.A( u2_u8_u7_n138 ) , .ZN( u2_u8_u7_n171 ) );
  INV_X1 u2_u8_u7_U27 (.A( u2_u8_u7_n131 ) , .ZN( u2_u8_u7_n177 ) );
  INV_X1 u2_u8_u7_U28 (.A( u2_u8_u7_n110 ) , .ZN( u2_u8_u7_n174 ) );
  NAND2_X1 u2_u8_u7_U29 (.A1( u2_u8_u7_n129 ) , .A2( u2_u8_u7_n132 ) , .ZN( u2_u8_u7_n149 ) );
  OAI21_X1 u2_u8_u7_U3 (.ZN( u2_u8_u7_n159 ) , .A( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n171 ) , .B1( u2_u8_u7_n174 ) );
  NAND2_X1 u2_u8_u7_U30 (.A1( u2_u8_u7_n113 ) , .A2( u2_u8_u7_n124 ) , .ZN( u2_u8_u7_n130 ) );
  INV_X1 u2_u8_u7_U31 (.A( u2_u8_u7_n112 ) , .ZN( u2_u8_u7_n173 ) );
  INV_X1 u2_u8_u7_U32 (.A( u2_u8_u7_n128 ) , .ZN( u2_u8_u7_n168 ) );
  INV_X1 u2_u8_u7_U33 (.A( u2_u8_u7_n148 ) , .ZN( u2_u8_u7_n169 ) );
  INV_X1 u2_u8_u7_U34 (.A( u2_u8_u7_n127 ) , .ZN( u2_u8_u7_n179 ) );
  NOR2_X1 u2_u8_u7_U35 (.ZN( u2_u8_u7_n101 ) , .A2( u2_u8_u7_n150 ) , .A1( u2_u8_u7_n156 ) );
  AOI211_X1 u2_u8_u7_U36 (.B( u2_u8_u7_n154 ) , .A( u2_u8_u7_n155 ) , .C1( u2_u8_u7_n156 ) , .ZN( u2_u8_u7_n157 ) , .C2( u2_u8_u7_n172 ) );
  INV_X1 u2_u8_u7_U37 (.A( u2_u8_u7_n153 ) , .ZN( u2_u8_u7_n172 ) );
  AOI211_X1 u2_u8_u7_U38 (.B( u2_u8_u7_n139 ) , .A( u2_u8_u7_n140 ) , .C2( u2_u8_u7_n141 ) , .ZN( u2_u8_u7_n142 ) , .C1( u2_u8_u7_n156 ) );
  NAND4_X1 u2_u8_u7_U39 (.A3( u2_u8_u7_n127 ) , .A2( u2_u8_u7_n128 ) , .A1( u2_u8_u7_n129 ) , .ZN( u2_u8_u7_n141 ) , .A4( u2_u8_u7_n147 ) );
  INV_X1 u2_u8_u7_U4 (.A( u2_u8_u7_n111 ) , .ZN( u2_u8_u7_n170 ) );
  AOI21_X1 u2_u8_u7_U40 (.A( u2_u8_u7_n137 ) , .B1( u2_u8_u7_n138 ) , .ZN( u2_u8_u7_n139 ) , .B2( u2_u8_u7_n146 ) );
  OAI22_X1 u2_u8_u7_U41 (.B1( u2_u8_u7_n136 ) , .ZN( u2_u8_u7_n140 ) , .A1( u2_u8_u7_n153 ) , .B2( u2_u8_u7_n162 ) , .A2( u2_u8_u7_n164 ) );
  AOI21_X1 u2_u8_u7_U42 (.ZN( u2_u8_u7_n123 ) , .B1( u2_u8_u7_n165 ) , .B2( u2_u8_u7_n177 ) , .A( u2_u8_u7_n97 ) );
  AOI21_X1 u2_u8_u7_U43 (.B2( u2_u8_u7_n113 ) , .B1( u2_u8_u7_n124 ) , .A( u2_u8_u7_n125 ) , .ZN( u2_u8_u7_n97 ) );
  INV_X1 u2_u8_u7_U44 (.A( u2_u8_u7_n125 ) , .ZN( u2_u8_u7_n161 ) );
  INV_X1 u2_u8_u7_U45 (.A( u2_u8_u7_n152 ) , .ZN( u2_u8_u7_n162 ) );
  AOI22_X1 u2_u8_u7_U46 (.A2( u2_u8_u7_n114 ) , .ZN( u2_u8_u7_n119 ) , .B1( u2_u8_u7_n130 ) , .A1( u2_u8_u7_n156 ) , .B2( u2_u8_u7_n165 ) );
  NAND2_X1 u2_u8_u7_U47 (.A2( u2_u8_u7_n112 ) , .ZN( u2_u8_u7_n114 ) , .A1( u2_u8_u7_n175 ) );
  AND2_X1 u2_u8_u7_U48 (.ZN( u2_u8_u7_n145 ) , .A2( u2_u8_u7_n98 ) , .A1( u2_u8_u7_n99 ) );
  NOR2_X1 u2_u8_u7_U49 (.ZN( u2_u8_u7_n137 ) , .A1( u2_u8_u7_n150 ) , .A2( u2_u8_u7_n161 ) );
  INV_X1 u2_u8_u7_U5 (.A( u2_u8_u7_n149 ) , .ZN( u2_u8_u7_n175 ) );
  AOI21_X1 u2_u8_u7_U50 (.ZN( u2_u8_u7_n105 ) , .B2( u2_u8_u7_n110 ) , .A( u2_u8_u7_n125 ) , .B1( u2_u8_u7_n147 ) );
  NAND2_X1 u2_u8_u7_U51 (.ZN( u2_u8_u7_n146 ) , .A1( u2_u8_u7_n95 ) , .A2( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U52 (.A2( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n147 ) , .A1( u2_u8_u7_n93 ) );
  NAND2_X1 u2_u8_u7_U53 (.A1( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n127 ) , .A2( u2_u8_u7_n99 ) );
  OR2_X1 u2_u8_u7_U54 (.ZN( u2_u8_u7_n126 ) , .A2( u2_u8_u7_n152 ) , .A1( u2_u8_u7_n156 ) );
  NAND2_X1 u2_u8_u7_U55 (.A2( u2_u8_u7_n102 ) , .A1( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n133 ) );
  NAND2_X1 u2_u8_u7_U56 (.ZN( u2_u8_u7_n112 ) , .A2( u2_u8_u7_n96 ) , .A1( u2_u8_u7_n99 ) );
  NAND2_X1 u2_u8_u7_U57 (.A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n128 ) , .A1( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U58 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n113 ) , .A2( u2_u8_u7_n93 ) );
  NAND2_X1 u2_u8_u7_U59 (.A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n124 ) , .A1( u2_u8_u7_n96 ) );
  INV_X1 u2_u8_u7_U6 (.A( u2_u8_u7_n154 ) , .ZN( u2_u8_u7_n178 ) );
  NAND2_X1 u2_u8_u7_U60 (.ZN( u2_u8_u7_n110 ) , .A1( u2_u8_u7_n95 ) , .A2( u2_u8_u7_n96 ) );
  INV_X1 u2_u8_u7_U61 (.A( u2_u8_u7_n150 ) , .ZN( u2_u8_u7_n164 ) );
  AND2_X1 u2_u8_u7_U62 (.ZN( u2_u8_u7_n134 ) , .A1( u2_u8_u7_n93 ) , .A2( u2_u8_u7_n98 ) );
  NAND2_X1 u2_u8_u7_U63 (.A1( u2_u8_u7_n100 ) , .A2( u2_u8_u7_n102 ) , .ZN( u2_u8_u7_n129 ) );
  NAND2_X1 u2_u8_u7_U64 (.A2( u2_u8_u7_n103 ) , .ZN( u2_u8_u7_n131 ) , .A1( u2_u8_u7_n95 ) );
  NAND2_X1 u2_u8_u7_U65 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n138 ) , .A2( u2_u8_u7_n99 ) );
  NAND2_X1 u2_u8_u7_U66 (.ZN( u2_u8_u7_n132 ) , .A1( u2_u8_u7_n93 ) , .A2( u2_u8_u7_n96 ) );
  NAND2_X1 u2_u8_u7_U67 (.A1( u2_u8_u7_n100 ) , .ZN( u2_u8_u7_n148 ) , .A2( u2_u8_u7_n95 ) );
  NOR2_X1 u2_u8_u7_U68 (.A2( u2_u8_X_47 ) , .ZN( u2_u8_u7_n150 ) , .A1( u2_u8_u7_n163 ) );
  NOR2_X1 u2_u8_u7_U69 (.A2( u2_u8_X_43 ) , .A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n103 ) );
  AOI211_X1 u2_u8_u7_U7 (.ZN( u2_u8_u7_n116 ) , .A( u2_u8_u7_n155 ) , .C1( u2_u8_u7_n161 ) , .C2( u2_u8_u7_n171 ) , .B( u2_u8_u7_n94 ) );
  NOR2_X1 u2_u8_u7_U70 (.A2( u2_u8_X_48 ) , .A1( u2_u8_u7_n166 ) , .ZN( u2_u8_u7_n95 ) );
  NOR2_X1 u2_u8_u7_U71 (.A2( u2_u8_X_45 ) , .A1( u2_u8_X_48 ) , .ZN( u2_u8_u7_n99 ) );
  NOR2_X1 u2_u8_u7_U72 (.A2( u2_u8_X_44 ) , .A1( u2_u8_u7_n167 ) , .ZN( u2_u8_u7_n98 ) );
  NOR2_X1 u2_u8_u7_U73 (.A2( u2_u8_X_46 ) , .A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n152 ) );
  AND2_X1 u2_u8_u7_U74 (.A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n156 ) , .A2( u2_u8_u7_n163 ) );
  NAND2_X1 u2_u8_u7_U75 (.A2( u2_u8_X_46 ) , .A1( u2_u8_X_47 ) , .ZN( u2_u8_u7_n125 ) );
  AND2_X1 u2_u8_u7_U76 (.A2( u2_u8_X_45 ) , .A1( u2_u8_X_48 ) , .ZN( u2_u8_u7_n102 ) );
  AND2_X1 u2_u8_u7_U77 (.A2( u2_u8_X_43 ) , .A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n96 ) );
  AND2_X1 u2_u8_u7_U78 (.A1( u2_u8_X_44 ) , .ZN( u2_u8_u7_n100 ) , .A2( u2_u8_u7_n167 ) );
  AND2_X1 u2_u8_u7_U79 (.A1( u2_u8_X_48 ) , .A2( u2_u8_u7_n166 ) , .ZN( u2_u8_u7_n93 ) );
  OAI222_X1 u2_u8_u7_U8 (.C2( u2_u8_u7_n101 ) , .B2( u2_u8_u7_n111 ) , .A1( u2_u8_u7_n113 ) , .C1( u2_u8_u7_n146 ) , .A2( u2_u8_u7_n162 ) , .B1( u2_u8_u7_n164 ) , .ZN( u2_u8_u7_n94 ) );
  INV_X1 u2_u8_u7_U80 (.A( u2_u8_X_46 ) , .ZN( u2_u8_u7_n163 ) );
  INV_X1 u2_u8_u7_U81 (.A( u2_u8_X_43 ) , .ZN( u2_u8_u7_n167 ) );
  INV_X1 u2_u8_u7_U82 (.A( u2_u8_X_45 ) , .ZN( u2_u8_u7_n166 ) );
  NAND4_X1 u2_u8_u7_U83 (.ZN( u2_out8_27 ) , .A4( u2_u8_u7_n118 ) , .A3( u2_u8_u7_n119 ) , .A2( u2_u8_u7_n120 ) , .A1( u2_u8_u7_n121 ) );
  OAI21_X1 u2_u8_u7_U84 (.ZN( u2_u8_u7_n121 ) , .B2( u2_u8_u7_n145 ) , .A( u2_u8_u7_n150 ) , .B1( u2_u8_u7_n174 ) );
  OAI21_X1 u2_u8_u7_U85 (.ZN( u2_u8_u7_n120 ) , .A( u2_u8_u7_n161 ) , .B2( u2_u8_u7_n170 ) , .B1( u2_u8_u7_n179 ) );
  NAND4_X1 u2_u8_u7_U86 (.ZN( u2_out8_21 ) , .A4( u2_u8_u7_n157 ) , .A3( u2_u8_u7_n158 ) , .A2( u2_u8_u7_n159 ) , .A1( u2_u8_u7_n160 ) );
  OAI21_X1 u2_u8_u7_U87 (.B1( u2_u8_u7_n145 ) , .ZN( u2_u8_u7_n160 ) , .A( u2_u8_u7_n161 ) , .B2( u2_u8_u7_n177 ) );
  AOI22_X1 u2_u8_u7_U88 (.B2( u2_u8_u7_n149 ) , .B1( u2_u8_u7_n150 ) , .A2( u2_u8_u7_n151 ) , .A1( u2_u8_u7_n152 ) , .ZN( u2_u8_u7_n158 ) );
  NAND4_X1 u2_u8_u7_U89 (.ZN( u2_out8_15 ) , .A4( u2_u8_u7_n142 ) , .A3( u2_u8_u7_n143 ) , .A2( u2_u8_u7_n144 ) , .A1( u2_u8_u7_n178 ) );
  OAI221_X1 u2_u8_u7_U9 (.C1( u2_u8_u7_n101 ) , .C2( u2_u8_u7_n147 ) , .ZN( u2_u8_u7_n155 ) , .B2( u2_u8_u7_n162 ) , .A( u2_u8_u7_n91 ) , .B1( u2_u8_u7_n92 ) );
  OR2_X1 u2_u8_u7_U90 (.A2( u2_u8_u7_n125 ) , .A1( u2_u8_u7_n129 ) , .ZN( u2_u8_u7_n144 ) );
  AOI22_X1 u2_u8_u7_U91 (.A2( u2_u8_u7_n126 ) , .ZN( u2_u8_u7_n143 ) , .B2( u2_u8_u7_n165 ) , .B1( u2_u8_u7_n173 ) , .A1( u2_u8_u7_n174 ) );
  NAND4_X1 u2_u8_u7_U92 (.ZN( u2_out8_5 ) , .A4( u2_u8_u7_n108 ) , .A3( u2_u8_u7_n109 ) , .A1( u2_u8_u7_n116 ) , .A2( u2_u8_u7_n123 ) );
  AOI22_X1 u2_u8_u7_U93 (.ZN( u2_u8_u7_n109 ) , .A2( u2_u8_u7_n126 ) , .B2( u2_u8_u7_n145 ) , .B1( u2_u8_u7_n156 ) , .A1( u2_u8_u7_n171 ) );
  NOR4_X1 u2_u8_u7_U94 (.A4( u2_u8_u7_n104 ) , .A3( u2_u8_u7_n105 ) , .A2( u2_u8_u7_n106 ) , .A1( u2_u8_u7_n107 ) , .ZN( u2_u8_u7_n108 ) );
  NAND3_X1 u2_u8_u7_U95 (.A3( u2_u8_u7_n146 ) , .A2( u2_u8_u7_n147 ) , .A1( u2_u8_u7_n148 ) , .ZN( u2_u8_u7_n151 ) );
  NAND3_X1 u2_u8_u7_U96 (.A3( u2_u8_u7_n131 ) , .A2( u2_u8_u7_n132 ) , .A1( u2_u8_u7_n133 ) , .ZN( u2_u8_u7_n135 ) );
  OAI21_X1 u2_uk_U1013 (.ZN( u2_K9_44 ) , .A( u2_uk_n1138 ) , .B2( u2_uk_n1585 ) , .B1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U1014 (.A1( u2_uk_K_r7_0 ) , .ZN( u2_uk_n1138 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1106 (.ZN( u2_K12_23 ) , .A( u2_uk_n454 ) );
  AOI22_X1 u2_uk_U1107 (.B2( u2_uk_K_r10_32 ) , .A2( u2_uk_K_r10_41 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n454 ) );
  INV_X1 u2_uk_U131 (.ZN( u2_K12_15 ) , .A( u2_uk_n409 ) );
  AOI22_X1 u2_uk_U132 (.B2( u2_uk_K_r10_25 ) , .A2( u2_uk_K_r10_34 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n222 ) , .ZN( u2_uk_n409 ) );
  OAI22_X1 u2_uk_U176 (.ZN( u2_K12_14 ) , .B2( u2_uk_n1688 ) , .A2( u2_uk_n1693 ) , .B1( u2_uk_n214 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U262 (.ZN( u2_K9_48 ) , .A( u2_uk_n1140 ) );
  OAI21_X1 u2_uk_U336 (.ZN( u2_K9_46 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1139 ) , .B2( u2_uk_n1577 ) );
  NAND2_X1 u2_uk_U337 (.A1( u2_uk_K_r7_37 ) , .A2( u2_uk_n10 ) , .ZN( u2_uk_n1139 ) );
  INV_X1 u2_uk_U542 (.ZN( u2_K12_17 ) , .A( u2_uk_n415 ) );
  OAI22_X1 u2_uk_U652 (.ZN( u2_K9_43 ) , .A1( u2_uk_n102 ) , .B2( u2_uk_n1558 ) , .A2( u2_uk_n1565 ) , .B1( u2_uk_n214 ) );
  OAI22_X1 u2_uk_U748 (.ZN( u2_K12_13 ) , .B2( u2_uk_n1689 ) , .A2( u2_uk_n1721 ) , .B1( u2_uk_n209 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U770 (.ZN( u2_K12_21 ) , .A( u2_uk_n443 ) );
  OAI22_X1 u2_uk_U909 (.ZN( u2_K9_47 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1576 ) , .A2( u2_uk_n1583 ) , .B1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U910 (.ZN( u2_K12_16 ) , .A2( u2_uk_n1681 ) , .B2( u2_uk_n1693 ) , .B1( u2_uk_n209 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U916 (.ZN( u2_K12_18 ) , .A2( u2_uk_n1683 ) , .B2( u2_uk_n1721 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U938 (.ZN( u2_K12_19 ) , .A1( u2_uk_n128 ) , .A2( u2_uk_n1682 ) , .B2( u2_uk_n1720 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U982 (.A1( u2_uk_K_r1_7 ) , .ZN( u2_uk_n1012 ) , .A2( u2_uk_n92 ) );
endmodule

