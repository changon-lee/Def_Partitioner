module des_des_die_4 ( u0_FP_33, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, 
       u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, 
       u0_K10_19, u0_K10_20, u0_K13_30, u0_K15_18, u0_K16_38, u0_K2_44, u0_K2_45, u0_K2_46, u0_K2_47, 
       u0_K2_48, u0_K6_27, u0_K6_41, u0_K7_22, u0_K7_23, u0_K9_14, u0_K9_15, u0_K9_4, u0_K9_45, 
       u0_K9_6, u0_L0_15, u0_L0_21, u0_L0_27, u0_L0_5, u0_L11_14, u0_L11_25, u0_L11_3, u0_L11_8, 
       u0_L13_1, u0_L13_10, u0_L13_11, u0_L13_13, u0_L13_16, u0_L13_18, u0_L13_19, u0_L13_2, u0_L13_20, 
       u0_L13_24, u0_L13_26, u0_L13_28, u0_L13_29, u0_L13_30, u0_L13_4, u0_L13_6, u0_L14_11, u0_L14_12, 
       u0_L14_15, u0_L14_19, u0_L14_21, u0_L14_22, u0_L14_27, u0_L14_29, u0_L14_32, u0_L14_4, u0_L14_5, 
       u0_L14_7, u0_L4_12, u0_L4_14, u0_L4_22, u0_L4_25, u0_L4_3, u0_L4_32, u0_L4_7, u0_L4_8, 
       u0_L5_1, u0_L5_10, u0_L5_14, u0_L5_20, u0_L5_25, u0_L5_26, u0_L5_3, u0_L5_8, u0_L7_1, 
       u0_L7_10, u0_L7_13, u0_L7_14, u0_L7_15, u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_2, u0_L7_20, 
       u0_L7_21, u0_L7_23, u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_28, u0_L7_3, u0_L7_30, 
       u0_L7_31, u0_L7_5, u0_L7_6, u0_L7_8, u0_L7_9, u0_L8_1, u0_L8_10, u0_L8_13, u0_L8_16, 
       u0_L8_18, u0_L8_2, u0_L8_20, u0_L8_24, u0_L8_26, u0_L8_28, u0_L8_30, u0_L8_6, u0_L9_14, 
       u0_L9_25, u0_L9_3, u0_L9_8, u0_R0_1, u0_R0_28, u0_R0_29, u0_R0_30, u0_R0_31, u0_R0_32, 
       u0_R11_16, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_20, u0_R11_21, u0_R13_10, u0_R13_11, u0_R13_12, 
       u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_17, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, 
       u0_R13_24, u0_R13_25, u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_8, u0_R13_9, u0_R4_16, 
       u0_R4_17, u0_R4_18, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_24, u0_R4_25, u0_R4_26, u0_R4_27, 
       u0_R4_28, u0_R4_29, u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_15, u0_R5_16, u0_R5_17, u0_R5_18, 
       u0_R5_19, u0_R5_20, u0_R5_21, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, u0_R7_13, u0_R7_14, 
       u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_20, u0_R7_21, u0_R7_28, 
       u0_R7_29, u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, 
       u0_R7_8, u0_R7_9, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, 
       u0_R8_17, u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_R9_16, u0_R9_17, 
       u0_R9_18, u0_R9_19, u0_R9_20, u0_R9_21, u0_uk_K_r0_2, u0_uk_K_r11_21, u0_uk_K_r12_18, u0_uk_K_r13_13, u0_uk_K_r13_17, 
       u0_uk_K_r13_19, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_4, u0_uk_K_r13_55, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_2, u0_uk_K_r14_3, 
       u0_uk_K_r14_43, u0_uk_K_r14_5, u0_uk_K_r14_50, u0_uk_K_r14_9, u0_uk_K_r4_0, u0_uk_K_r4_31, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r5_18, 
       u0_uk_K_r5_19, u0_uk_K_r5_23, u0_uk_K_r5_40, u0_uk_K_r5_43, u0_uk_K_r6_51, u0_uk_K_r6_55, u0_uk_K_r7_0, u0_uk_K_r7_13, u0_uk_K_r7_2, 
       u0_uk_K_r7_20, u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_48, u0_uk_K_r7_55, 
       u0_uk_K_r7_6, u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_17, u0_uk_K_r8_27, u0_uk_K_r8_32, u0_uk_K_r8_40, u0_uk_K_r9_0, u0_uk_K_r9_1, 
       u0_uk_K_r9_35, u0_uk_K_r9_9, u0_uk_n10, u0_uk_n100, u0_uk_n1019, u0_uk_n102, u0_uk_n1020, u0_uk_n1024, u0_uk_n105, 
       u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n111, u0_uk_n113, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n123, 
       u0_uk_n129, u0_uk_n13, u0_uk_n134, u0_uk_n14, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, 
       u0_uk_n15, u0_uk_n155, u0_uk_n16, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n18, 
       u0_uk_n182, u0_uk_n184, u0_uk_n19, u0_uk_n191, u0_uk_n192, u0_uk_n193, u0_uk_n198, u0_uk_n202, u0_uk_n203, 
       u0_uk_n204, u0_uk_n207, u0_uk_n208, u0_uk_n211, u0_uk_n213, u0_uk_n214, u0_uk_n216, u0_uk_n217, u0_uk_n220, 
       u0_uk_n222, u0_uk_n223, u0_uk_n224, u0_uk_n228, u0_uk_n229, u0_uk_n230, u0_uk_n231, u0_uk_n234, u0_uk_n238, 
       u0_uk_n24, u0_uk_n240, u0_uk_n242, u0_uk_n245, u0_uk_n25, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n253, 
       u0_uk_n254, u0_uk_n257, u0_uk_n259, u0_uk_n26, u0_uk_n262, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n27, 
       u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, u0_uk_n278, u0_uk_n28, u0_uk_n280, u0_uk_n281, u0_uk_n282, 
       u0_uk_n285, u0_uk_n288, u0_uk_n289, u0_uk_n29, u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n30, u0_uk_n300, 
       u0_uk_n303, u0_uk_n304, u0_uk_n309, u0_uk_n31, u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, u0_uk_n32, 
       u0_uk_n33, u0_uk_n35, u0_uk_n362, u0_uk_n367, u0_uk_n368, u0_uk_n37, u0_uk_n378, u0_uk_n38, u0_uk_n383, 
       u0_uk_n387, u0_uk_n388, u0_uk_n393, u0_uk_n398, u0_uk_n399, u0_uk_n4, u0_uk_n411, u0_uk_n413, u0_uk_n418, 
       u0_uk_n419, u0_uk_n42, u0_uk_n420, u0_uk_n428, u0_uk_n43, u0_uk_n433, u0_uk_n434, u0_uk_n438, u0_uk_n44, 
       u0_uk_n440, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n45, u0_uk_n450, u0_uk_n60, u0_uk_n612, u0_uk_n63, 
       u0_uk_n632, u0_uk_n633, u0_uk_n635, u0_uk_n638, u0_uk_n641, u0_uk_n642, u0_uk_n643, u0_uk_n647, u0_uk_n648, 
       u0_uk_n649, u0_uk_n650, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n663, u0_uk_n666, u0_uk_n669, u0_uk_n670, 
       u0_uk_n7, u0_uk_n719, u0_uk_n720, u0_uk_n728, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, 
       u0_uk_n740, u0_uk_n775, u0_uk_n780, u0_uk_n8, u0_uk_n83, u0_uk_n897, u0_uk_n898, u0_uk_n917, u0_uk_n918, 
       u0_uk_n93, u0_uk_n94, u0_uk_n948, u0_uk_n98, u1_FP_34, u1_FP_35, u1_K10_27, u1_K10_28, u1_K11_10, 
       u1_K11_27, u1_K11_28, u1_K11_29, u1_K11_3, u1_K11_32, u1_K11_33, u1_K11_4, u1_K11_6, u1_K11_7, 
       u1_K11_9, u1_K12_33, u1_K12_34, u1_K13_39, u1_K13_40, u1_K14_33, u1_K15_27, u1_K15_28, u1_K16_3, 
       u1_K16_4, u1_K1_15, u1_K1_16, u1_K3_15, u1_K3_16, u1_K3_33, u1_K3_34, u1_K5_10, u1_K5_21, 
       u1_K5_3, u1_K5_4, u1_K5_5, u1_K5_7, u1_K5_9, u1_K7_28, u1_K7_3, u1_K7_39, u1_K7_4, 
       u1_K7_40, u1_K8_21, u1_K8_22, u1_K9_34, u1_L10_11, u1_L10_19, u1_L10_29, u1_L10_4, u1_L11_12, 
       u1_L11_22, u1_L11_32, u1_L11_7, u1_L12_11, u1_L12_19, u1_L12_29, u1_L12_4, u1_L13_14, u1_L13_25, 
       u1_L13_3, u1_L13_8, u1_L14_17, u1_L14_23, u1_L14_31, u1_L14_9, u1_L1_11, u1_L1_16, u1_L1_19, 
       u1_L1_24, u1_L1_29, u1_L1_30, u1_L1_4, u1_L1_6, u1_L2_17, u1_L2_23, u1_L2_31, u1_L2_9, 
       u1_L3_1, u1_L3_10, u1_L3_13, u1_L3_17, u1_L3_18, u1_L3_2, u1_L3_20, u1_L3_23, u1_L3_26, 
       u1_L3_28, u1_L3_31, u1_L3_9, u1_L5_12, u1_L5_14, u1_L5_17, u1_L5_22, u1_L5_23, u1_L5_25, 
       u1_L5_3, u1_L5_31, u1_L5_32, u1_L5_7, u1_L5_8, u1_L5_9, u1_L6_1, u1_L6_10, u1_L6_20, 
       u1_L6_26, u1_L7_11, u1_L7_19, u1_L7_29, u1_L7_4, u1_L8_14, u1_L8_25, u1_L8_3, u1_L8_8, 
       u1_L9_11, u1_L9_13, u1_L9_14, u1_L9_17, u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_23, u1_L9_25, 
       u1_L9_28, u1_L9_29, u1_L9_3, u1_L9_31, u1_L9_4, u1_L9_8, u1_L9_9, u1_R10_22, u1_R10_23, 
       u1_R11_26, u1_R11_27, u1_R12_22, u1_R12_23, u1_R13_18, u1_R13_19, u1_R1_10, u1_R1_11, u1_R1_22, 
       u1_R1_23, u1_R2_2, u1_R2_3, u1_R3_14, u1_R3_15, u1_R3_2, u1_R3_3, u1_R3_4, u1_R3_6, 
       u1_R3_7, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_26, u1_R5_27, u1_R5_3, u1_R6_14, u1_R6_15, 
       u1_R7_22, u1_R7_23, u1_R8_18, u1_R8_19, u1_R9_18, u1_R9_19, u1_R9_2, u1_R9_20, u1_R9_21, 
       u1_R9_22, u1_R9_23, u1_R9_3, u1_R9_4, u1_R9_5, u1_R9_6, u1_R9_7, u1_desIn_r_13, u1_desIn_r_21, 
       u1_desIn_r_40, u1_desIn_r_46, u1_desIn_r_58, u1_desIn_r_60, u1_u0_X_13, u1_u0_X_14, u1_u0_X_17, u1_u0_X_18, u1_u10_X_1, 
       u1_u10_X_11, u1_u10_X_12, u1_u10_X_2, u1_u10_X_25, u1_u10_X_26, u1_u10_X_35, u1_u10_X_36, u1_u11_X_31, u1_u11_X_32, 
       u1_u11_X_35, u1_u11_X_36, u1_u12_X_37, u1_u12_X_38, u1_u12_X_41, u1_u12_X_42, u1_u13_X_31, u1_u13_X_32, u1_u13_X_35, 
       u1_u13_X_36, u1_u14_X_25, u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u15_X_1, u1_u15_X_2, u1_u15_X_5, u1_u15_X_6, 
       u1_u2_X_13, u1_u2_X_14, u1_u2_X_17, u1_u2_X_18, u1_u2_X_31, u1_u2_X_32, u1_u2_X_35, u1_u2_X_36, u1_u3_X_1, 
       u1_u3_X_2, u1_u3_X_5, u1_u3_X_6, u1_u4_X_1, u1_u4_X_11, u1_u4_X_12, u1_u4_X_19, u1_u4_X_2, u1_u4_X_20, 
       u1_u4_X_23, u1_u4_X_24, u1_u4_X_6, u1_u4_X_8, u1_u6_X_1, u1_u6_X_2, u1_u6_X_25, u1_u6_X_26, u1_u6_X_29, 
       u1_u6_X_30, u1_u6_X_37, u1_u6_X_38, u1_u6_X_41, u1_u6_X_42, u1_u6_X_5, u1_u6_X_6, u1_u7_X_19, u1_u7_X_20, 
       u1_u7_X_23, u1_u7_X_24, u1_u8_X_31, u1_u8_X_32, u1_u8_X_35, u1_u8_X_36, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, 
       u1_u9_X_30, u1_uk_n1065, u1_uk_n1067, u1_uk_n1074, u1_uk_n1115, u1_uk_n1162, u1_uk_n421, u1_uk_n437, u1_uk_n443, 
       u1_uk_n496, u1_uk_n501, u1_uk_n955, u2_K8_24, u2_L6_1, u2_L6_10, u2_L6_20, u2_L6_26, u2_R6_12, 
       u2_R6_13, u2_R6_14, u2_R6_15, u2_R6_16, u2_R6_17, u2_uk_n1508, u2_uk_n1513, u2_uk_n1515, u2_uk_n1518, 
       u2_uk_n1521, u2_uk_n1522, u2_uk_n1527, u2_uk_n1528, u2_uk_n1529, u2_uk_n1535, u2_uk_n202, u2_uk_n213, u2_uk_n220, 
       u2_uk_n27, u0_FP_11, u0_FP_12, u0_FP_15, u0_FP_19, u0_FP_21, u0_FP_22, u0_FP_27, u0_FP_29, u0_FP_32, 
        u0_FP_4, u0_FP_5, u0_FP_7, u0_N162, u0_N166, u0_N167, u0_N171, u0_N173, u0_N181, 
        u0_N184, u0_N191, u0_N192, u0_N194, u0_N199, u0_N201, u0_N205, u0_N211, u0_N216, 
        u0_N217, u0_N256, u0_N257, u0_N258, u0_N260, u0_N261, u0_N263, u0_N264, u0_N265, 
        u0_N268, u0_N269, u0_N270, u0_N271, u0_N272, u0_N273, u0_N275, u0_N276, u0_N278, 
        u0_N279, u0_N280, u0_N281, u0_N282, u0_N283, u0_N285, u0_N286, u0_N288, u0_N289, 
        u0_N293, u0_N297, u0_N300, u0_N303, u0_N305, u0_N307, u0_N311, u0_N313, u0_N315, 
        u0_N317, u0_N322, u0_N327, u0_N333, u0_N344, u0_N36, u0_N386, u0_N391, u0_N397, 
        u0_N408, u0_N448, u0_N449, u0_N451, u0_N453, u0_N457, u0_N458, u0_N46, u0_N460, 
        u0_N463, u0_N465, u0_N466, u0_N467, u0_N471, u0_N473, u0_N475, u0_N476, u0_N477, 
        u0_N52, u0_N58, u0_uk_n128, u0_uk_n187, u0_uk_n188, u0_uk_n756, u0_uk_n762, u0_uk_n790, u0_uk_n894, 
        u0_uk_n906, u0_uk_n92, u0_uk_n926, u0_uk_n99, u1_FP_17, u1_FP_23, u1_FP_31, u1_FP_9, u1_N104, 
        u1_N112, u1_N118, u1_N126, u1_N128, u1_N129, u1_N136, u1_N137, u1_N140, u1_N144, 
        u1_N145, u1_N147, u1_N15, u1_N150, u1_N153, u1_N155, u1_N158, u1_N194, u1_N198, 
        u1_N199, u1_N200, u1_N203, u1_N205, u1_N208, u1_N213, u1_N214, u1_N216, u1_N222, 
        u1_N223, u1_N224, u1_N23, u1_N233, u1_N243, u1_N249, u1_N259, u1_N266, u1_N274, 
        u1_N284, u1_N29, u1_N290, u1_N295, u1_N301, u1_N312, u1_N321, u1_N322, u1_N323, 
        u1_N327, u1_N328, u1_N330, u1_N332, u1_N333, u1_N336, u1_N337, u1_N338, u1_N342, 
        u1_N344, u1_N347, u1_N348, u1_N350, u1_N355, u1_N362, u1_N370, u1_N380, u1_N390, 
        u1_N395, u1_N405, u1_N415, u1_N419, u1_N426, u1_N434, u1_N444, u1_N450, u1_N455, 
        u1_N461, u1_N472, u1_N5, u1_N67, u1_N69, u1_N74, u1_N79, u1_N82, u1_N87, 
        u1_N92, u1_N93, u2_N224, u2_N233, u2_N243, u2_N249 );
  input u0_FP_33, u0_FP_52, u0_FP_53, u0_FP_54, u0_FP_55, u0_FP_56, u0_FP_57, u0_FP_58, u0_FP_59, 
        u0_FP_60, u0_FP_61, u0_FP_62, u0_FP_63, u0_FP_64, u0_K10_10, u0_K10_13, u0_K10_14, u0_K10_18, 
        u0_K10_19, u0_K10_20, u0_K13_30, u0_K15_18, u0_K16_38, u0_K2_44, u0_K2_45, u0_K2_46, u0_K2_47, 
        u0_K2_48, u0_K6_27, u0_K6_41, u0_K7_22, u0_K7_23, u0_K9_14, u0_K9_15, u0_K9_4, u0_K9_45, 
        u0_K9_6, u0_L0_15, u0_L0_21, u0_L0_27, u0_L0_5, u0_L11_14, u0_L11_25, u0_L11_3, u0_L11_8, 
        u0_L13_1, u0_L13_10, u0_L13_11, u0_L13_13, u0_L13_16, u0_L13_18, u0_L13_19, u0_L13_2, u0_L13_20, 
        u0_L13_24, u0_L13_26, u0_L13_28, u0_L13_29, u0_L13_30, u0_L13_4, u0_L13_6, u0_L14_11, u0_L14_12, 
        u0_L14_15, u0_L14_19, u0_L14_21, u0_L14_22, u0_L14_27, u0_L14_29, u0_L14_32, u0_L14_4, u0_L14_5, 
        u0_L14_7, u0_L4_12, u0_L4_14, u0_L4_22, u0_L4_25, u0_L4_3, u0_L4_32, u0_L4_7, u0_L4_8, 
        u0_L5_1, u0_L5_10, u0_L5_14, u0_L5_20, u0_L5_25, u0_L5_26, u0_L5_3, u0_L5_8, u0_L7_1, 
        u0_L7_10, u0_L7_13, u0_L7_14, u0_L7_15, u0_L7_16, u0_L7_17, u0_L7_18, u0_L7_2, u0_L7_20, 
        u0_L7_21, u0_L7_23, u0_L7_24, u0_L7_25, u0_L7_26, u0_L7_27, u0_L7_28, u0_L7_3, u0_L7_30, 
        u0_L7_31, u0_L7_5, u0_L7_6, u0_L7_8, u0_L7_9, u0_L8_1, u0_L8_10, u0_L8_13, u0_L8_16, 
        u0_L8_18, u0_L8_2, u0_L8_20, u0_L8_24, u0_L8_26, u0_L8_28, u0_L8_30, u0_L8_6, u0_L9_14, 
        u0_L9_25, u0_L9_3, u0_L9_8, u0_R0_1, u0_R0_28, u0_R0_29, u0_R0_30, u0_R0_31, u0_R0_32, 
        u0_R11_16, u0_R11_17, u0_R11_18, u0_R11_19, u0_R11_20, u0_R11_21, u0_R13_10, u0_R13_11, u0_R13_12, 
        u0_R13_13, u0_R13_14, u0_R13_15, u0_R13_16, u0_R13_17, u0_R13_20, u0_R13_21, u0_R13_22, u0_R13_23, 
        u0_R13_24, u0_R13_25, u0_R13_4, u0_R13_5, u0_R13_6, u0_R13_7, u0_R13_8, u0_R13_9, u0_R4_16, 
        u0_R4_17, u0_R4_18, u0_R4_19, u0_R4_20, u0_R4_21, u0_R4_24, u0_R4_25, u0_R4_26, u0_R4_27, 
        u0_R4_28, u0_R4_29, u0_R5_12, u0_R5_13, u0_R5_14, u0_R5_15, u0_R5_16, u0_R5_17, u0_R5_18, 
        u0_R5_19, u0_R5_20, u0_R5_21, u0_R7_1, u0_R7_10, u0_R7_11, u0_R7_12, u0_R7_13, u0_R7_14, 
        u0_R7_15, u0_R7_16, u0_R7_17, u0_R7_18, u0_R7_19, u0_R7_2, u0_R7_20, u0_R7_21, u0_R7_28, 
        u0_R7_29, u0_R7_3, u0_R7_30, u0_R7_31, u0_R7_32, u0_R7_4, u0_R7_5, u0_R7_6, u0_R7_7, 
        u0_R7_8, u0_R7_9, u0_R8_10, u0_R8_11, u0_R8_12, u0_R8_13, u0_R8_14, u0_R8_15, u0_R8_16, 
        u0_R8_17, u0_R8_4, u0_R8_5, u0_R8_6, u0_R8_7, u0_R8_8, u0_R8_9, u0_R9_16, u0_R9_17, 
        u0_R9_18, u0_R9_19, u0_R9_20, u0_R9_21, u0_uk_K_r0_2, u0_uk_K_r11_21, u0_uk_K_r12_18, u0_uk_K_r13_13, u0_uk_K_r13_17, 
        u0_uk_K_r13_19, u0_uk_K_r13_25, u0_uk_K_r13_32, u0_uk_K_r13_4, u0_uk_K_r13_55, u0_uk_K_r14_15, u0_uk_K_r14_16, u0_uk_K_r14_2, u0_uk_K_r14_3, 
        u0_uk_K_r14_43, u0_uk_K_r14_5, u0_uk_K_r14_50, u0_uk_K_r14_9, u0_uk_K_r4_0, u0_uk_K_r4_31, u0_uk_K_r4_35, u0_uk_K_r4_38, u0_uk_K_r5_18, 
        u0_uk_K_r5_19, u0_uk_K_r5_23, u0_uk_K_r5_40, u0_uk_K_r5_43, u0_uk_K_r6_51, u0_uk_K_r6_55, u0_uk_K_r7_0, u0_uk_K_r7_13, u0_uk_K_r7_2, 
        u0_uk_K_r7_20, u0_uk_K_r7_24, u0_uk_K_r7_25, u0_uk_K_r7_26, u0_uk_K_r7_27, u0_uk_K_r7_32, u0_uk_K_r7_39, u0_uk_K_r7_48, u0_uk_K_r7_55, 
        u0_uk_K_r7_6, u0_uk_K_r7_9, u0_uk_K_r8_13, u0_uk_K_r8_17, u0_uk_K_r8_27, u0_uk_K_r8_32, u0_uk_K_r8_40, u0_uk_K_r9_0, u0_uk_K_r9_1, 
        u0_uk_K_r9_35, u0_uk_K_r9_9, u0_uk_n10, u0_uk_n100, u0_uk_n1019, u0_uk_n102, u0_uk_n1020, u0_uk_n1024, u0_uk_n105, 
        u0_uk_n109, u0_uk_n11, u0_uk_n110, u0_uk_n111, u0_uk_n113, u0_uk_n116, u0_uk_n117, u0_uk_n118, u0_uk_n123, 
        u0_uk_n129, u0_uk_n13, u0_uk_n134, u0_uk_n14, u0_uk_n141, u0_uk_n142, u0_uk_n145, u0_uk_n146, u0_uk_n147, 
        u0_uk_n15, u0_uk_n155, u0_uk_n16, u0_uk_n161, u0_uk_n162, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n18, 
        u0_uk_n182, u0_uk_n184, u0_uk_n19, u0_uk_n191, u0_uk_n192, u0_uk_n193, u0_uk_n198, u0_uk_n202, u0_uk_n203, 
        u0_uk_n204, u0_uk_n207, u0_uk_n208, u0_uk_n211, u0_uk_n213, u0_uk_n214, u0_uk_n216, u0_uk_n217, u0_uk_n220, 
        u0_uk_n222, u0_uk_n223, u0_uk_n224, u0_uk_n228, u0_uk_n229, u0_uk_n230, u0_uk_n231, u0_uk_n234, u0_uk_n238, 
        u0_uk_n24, u0_uk_n240, u0_uk_n242, u0_uk_n245, u0_uk_n25, u0_uk_n250, u0_uk_n251, u0_uk_n252, u0_uk_n253, 
        u0_uk_n254, u0_uk_n257, u0_uk_n259, u0_uk_n26, u0_uk_n262, u0_uk_n266, u0_uk_n267, u0_uk_n268, u0_uk_n27, 
        u0_uk_n272, u0_uk_n273, u0_uk_n274, u0_uk_n275, u0_uk_n278, u0_uk_n28, u0_uk_n280, u0_uk_n281, u0_uk_n282, 
        u0_uk_n285, u0_uk_n288, u0_uk_n289, u0_uk_n29, u0_uk_n290, u0_uk_n293, u0_uk_n296, u0_uk_n30, u0_uk_n300, 
        u0_uk_n303, u0_uk_n304, u0_uk_n309, u0_uk_n31, u0_uk_n310, u0_uk_n311, u0_uk_n314, u0_uk_n315, u0_uk_n32, 
        u0_uk_n33, u0_uk_n35, u0_uk_n362, u0_uk_n367, u0_uk_n368, u0_uk_n37, u0_uk_n378, u0_uk_n38, u0_uk_n383, 
        u0_uk_n387, u0_uk_n388, u0_uk_n393, u0_uk_n398, u0_uk_n399, u0_uk_n4, u0_uk_n411, u0_uk_n413, u0_uk_n418, 
        u0_uk_n419, u0_uk_n42, u0_uk_n420, u0_uk_n428, u0_uk_n43, u0_uk_n433, u0_uk_n434, u0_uk_n438, u0_uk_n44, 
        u0_uk_n440, u0_uk_n445, u0_uk_n446, u0_uk_n447, u0_uk_n45, u0_uk_n450, u0_uk_n60, u0_uk_n612, u0_uk_n63, 
        u0_uk_n632, u0_uk_n633, u0_uk_n635, u0_uk_n638, u0_uk_n641, u0_uk_n642, u0_uk_n643, u0_uk_n647, u0_uk_n648, 
        u0_uk_n649, u0_uk_n650, u0_uk_n655, u0_uk_n657, u0_uk_n658, u0_uk_n663, u0_uk_n666, u0_uk_n669, u0_uk_n670, 
        u0_uk_n7, u0_uk_n719, u0_uk_n720, u0_uk_n728, u0_uk_n731, u0_uk_n732, u0_uk_n735, u0_uk_n736, u0_uk_n739, 
        u0_uk_n740, u0_uk_n775, u0_uk_n780, u0_uk_n8, u0_uk_n83, u0_uk_n897, u0_uk_n898, u0_uk_n917, u0_uk_n918, 
        u0_uk_n93, u0_uk_n94, u0_uk_n948, u0_uk_n98, u1_FP_34, u1_FP_35, u1_K10_27, u1_K10_28, u1_K11_10, 
        u1_K11_27, u1_K11_28, u1_K11_29, u1_K11_3, u1_K11_32, u1_K11_33, u1_K11_4, u1_K11_6, u1_K11_7, 
        u1_K11_9, u1_K12_33, u1_K12_34, u1_K13_39, u1_K13_40, u1_K14_33, u1_K15_27, u1_K15_28, u1_K16_3, 
        u1_K16_4, u1_K1_15, u1_K1_16, u1_K3_15, u1_K3_16, u1_K3_33, u1_K3_34, u1_K5_10, u1_K5_21, 
        u1_K5_3, u1_K5_4, u1_K5_5, u1_K5_7, u1_K5_9, u1_K7_28, u1_K7_3, u1_K7_39, u1_K7_4, 
        u1_K7_40, u1_K8_21, u1_K8_22, u1_K9_34, u1_L10_11, u1_L10_19, u1_L10_29, u1_L10_4, u1_L11_12, 
        u1_L11_22, u1_L11_32, u1_L11_7, u1_L12_11, u1_L12_19, u1_L12_29, u1_L12_4, u1_L13_14, u1_L13_25, 
        u1_L13_3, u1_L13_8, u1_L14_17, u1_L14_23, u1_L14_31, u1_L14_9, u1_L1_11, u1_L1_16, u1_L1_19, 
        u1_L1_24, u1_L1_29, u1_L1_30, u1_L1_4, u1_L1_6, u1_L2_17, u1_L2_23, u1_L2_31, u1_L2_9, 
        u1_L3_1, u1_L3_10, u1_L3_13, u1_L3_17, u1_L3_18, u1_L3_2, u1_L3_20, u1_L3_23, u1_L3_26, 
        u1_L3_28, u1_L3_31, u1_L3_9, u1_L5_12, u1_L5_14, u1_L5_17, u1_L5_22, u1_L5_23, u1_L5_25, 
        u1_L5_3, u1_L5_31, u1_L5_32, u1_L5_7, u1_L5_8, u1_L5_9, u1_L6_1, u1_L6_10, u1_L6_20, 
        u1_L6_26, u1_L7_11, u1_L7_19, u1_L7_29, u1_L7_4, u1_L8_14, u1_L8_25, u1_L8_3, u1_L8_8, 
        u1_L9_11, u1_L9_13, u1_L9_14, u1_L9_17, u1_L9_18, u1_L9_19, u1_L9_2, u1_L9_23, u1_L9_25, 
        u1_L9_28, u1_L9_29, u1_L9_3, u1_L9_31, u1_L9_4, u1_L9_8, u1_L9_9, u1_R10_22, u1_R10_23, 
        u1_R11_26, u1_R11_27, u1_R12_22, u1_R12_23, u1_R13_18, u1_R13_19, u1_R1_10, u1_R1_11, u1_R1_22, 
        u1_R1_23, u1_R2_2, u1_R2_3, u1_R3_14, u1_R3_15, u1_R3_2, u1_R3_3, u1_R3_4, u1_R3_6, 
        u1_R3_7, u1_R5_18, u1_R5_19, u1_R5_2, u1_R5_26, u1_R5_27, u1_R5_3, u1_R6_14, u1_R6_15, 
        u1_R7_22, u1_R7_23, u1_R8_18, u1_R8_19, u1_R9_18, u1_R9_19, u1_R9_2, u1_R9_20, u1_R9_21, 
        u1_R9_22, u1_R9_23, u1_R9_3, u1_R9_4, u1_R9_5, u1_R9_6, u1_R9_7, u1_desIn_r_13, u1_desIn_r_21, 
        u1_desIn_r_40, u1_desIn_r_46, u1_desIn_r_58, u1_desIn_r_60, u1_u0_X_13, u1_u0_X_14, u1_u0_X_17, u1_u0_X_18, u1_u10_X_1, 
        u1_u10_X_11, u1_u10_X_12, u1_u10_X_2, u1_u10_X_25, u1_u10_X_26, u1_u10_X_35, u1_u10_X_36, u1_u11_X_31, u1_u11_X_32, 
        u1_u11_X_35, u1_u11_X_36, u1_u12_X_37, u1_u12_X_38, u1_u12_X_41, u1_u12_X_42, u1_u13_X_31, u1_u13_X_32, u1_u13_X_35, 
        u1_u13_X_36, u1_u14_X_25, u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u15_X_1, u1_u15_X_2, u1_u15_X_5, u1_u15_X_6, 
        u1_u2_X_13, u1_u2_X_14, u1_u2_X_17, u1_u2_X_18, u1_u2_X_31, u1_u2_X_32, u1_u2_X_35, u1_u2_X_36, u1_u3_X_1, 
        u1_u3_X_2, u1_u3_X_5, u1_u3_X_6, u1_u4_X_1, u1_u4_X_11, u1_u4_X_12, u1_u4_X_19, u1_u4_X_2, u1_u4_X_20, 
        u1_u4_X_23, u1_u4_X_24, u1_u4_X_6, u1_u4_X_8, u1_u6_X_1, u1_u6_X_2, u1_u6_X_25, u1_u6_X_26, u1_u6_X_29, 
        u1_u6_X_30, u1_u6_X_37, u1_u6_X_38, u1_u6_X_41, u1_u6_X_42, u1_u6_X_5, u1_u6_X_6, u1_u7_X_19, u1_u7_X_20, 
        u1_u7_X_23, u1_u7_X_24, u1_u8_X_31, u1_u8_X_32, u1_u8_X_35, u1_u8_X_36, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, 
        u1_u9_X_30, u1_uk_n1065, u1_uk_n1067, u1_uk_n1074, u1_uk_n1115, u1_uk_n1162, u1_uk_n421, u1_uk_n437, u1_uk_n443, 
        u1_uk_n496, u1_uk_n501, u1_uk_n955, u2_K8_24, u2_L6_1, u2_L6_10, u2_L6_20, u2_L6_26, u2_R6_12, 
        u2_R6_13, u2_R6_14, u2_R6_15, u2_R6_16, u2_R6_17, u2_uk_n1508, u2_uk_n1513, u2_uk_n1515, u2_uk_n1518, 
        u2_uk_n1521, u2_uk_n1522, u2_uk_n1527, u2_uk_n1528, u2_uk_n1529, u2_uk_n1535, u2_uk_n202, u2_uk_n213, u2_uk_n220, 
        u2_uk_n27;
  output u0_FP_11, u0_FP_12, u0_FP_15, u0_FP_19, u0_FP_21, u0_FP_22, u0_FP_27, u0_FP_29, u0_FP_32, 
        u0_FP_4, u0_FP_5, u0_FP_7, u0_N162, u0_N166, u0_N167, u0_N171, u0_N173, u0_N181, 
        u0_N184, u0_N191, u0_N192, u0_N194, u0_N199, u0_N201, u0_N205, u0_N211, u0_N216, 
        u0_N217, u0_N256, u0_N257, u0_N258, u0_N260, u0_N261, u0_N263, u0_N264, u0_N265, 
        u0_N268, u0_N269, u0_N270, u0_N271, u0_N272, u0_N273, u0_N275, u0_N276, u0_N278, 
        u0_N279, u0_N280, u0_N281, u0_N282, u0_N283, u0_N285, u0_N286, u0_N288, u0_N289, 
        u0_N293, u0_N297, u0_N300, u0_N303, u0_N305, u0_N307, u0_N311, u0_N313, u0_N315, 
        u0_N317, u0_N322, u0_N327, u0_N333, u0_N344, u0_N36, u0_N386, u0_N391, u0_N397, 
        u0_N408, u0_N448, u0_N449, u0_N451, u0_N453, u0_N457, u0_N458, u0_N46, u0_N460, 
        u0_N463, u0_N465, u0_N466, u0_N467, u0_N471, u0_N473, u0_N475, u0_N476, u0_N477, 
        u0_N52, u0_N58, u0_uk_n128, u0_uk_n187, u0_uk_n188, u0_uk_n756, u0_uk_n762, u0_uk_n790, u0_uk_n894, 
        u0_uk_n906, u0_uk_n92, u0_uk_n926, u0_uk_n99, u1_FP_17, u1_FP_23, u1_FP_31, u1_FP_9, u1_N104, 
        u1_N112, u1_N118, u1_N126, u1_N128, u1_N129, u1_N136, u1_N137, u1_N140, u1_N144, 
        u1_N145, u1_N147, u1_N15, u1_N150, u1_N153, u1_N155, u1_N158, u1_N194, u1_N198, 
        u1_N199, u1_N200, u1_N203, u1_N205, u1_N208, u1_N213, u1_N214, u1_N216, u1_N222, 
        u1_N223, u1_N224, u1_N23, u1_N233, u1_N243, u1_N249, u1_N259, u1_N266, u1_N274, 
        u1_N284, u1_N29, u1_N290, u1_N295, u1_N301, u1_N312, u1_N321, u1_N322, u1_N323, 
        u1_N327, u1_N328, u1_N330, u1_N332, u1_N333, u1_N336, u1_N337, u1_N338, u1_N342, 
        u1_N344, u1_N347, u1_N348, u1_N350, u1_N355, u1_N362, u1_N370, u1_N380, u1_N390, 
        u1_N395, u1_N405, u1_N415, u1_N419, u1_N426, u1_N434, u1_N444, u1_N450, u1_N455, 
        u1_N461, u1_N472, u1_N5, u1_N67, u1_N69, u1_N74, u1_N79, u1_N82, u1_N87, 
        u1_N92, u1_N93, u2_N224, u2_N233, u2_N243, u2_N249;
  wire u0_K10_11, u0_K10_12, u0_K10_15, u0_K10_16, u0_K10_17, u0_K10_21, u0_K10_22, u0_K10_23, u0_K10_24, 
       u0_K10_7, u0_K10_8, u0_K10_9, u0_K11_25, u0_K11_26, u0_K11_27, u0_K11_28, u0_K11_29, u0_K11_30, 
       u0_K13_25, u0_K13_26, u0_K13_27, u0_K13_28, u0_K13_29, u0_K15_10, u0_K15_11, u0_K15_12, u0_K15_13, 
       u0_K15_14, u0_K15_15, u0_K15_16, u0_K15_17, u0_K15_19, u0_K15_20, u0_K15_21, u0_K15_22, u0_K15_23, 
       u0_K15_24, u0_K15_31, u0_K15_32, u0_K15_33, u0_K15_34, u0_K15_35, u0_K15_36, u0_K15_7, u0_K15_8, 
       u0_K15_9, u0_K16_31, u0_K16_32, u0_K16_33, u0_K16_34, u0_K16_35, u0_K16_36, u0_K16_37, u0_K16_39, 
       u0_K16_40, u0_K16_41, u0_K16_42, u0_K16_43, u0_K16_44, u0_K16_45, u0_K16_46, u0_K16_47, u0_K16_48, 
       u0_K2_43, u0_K6_25, u0_K6_26, u0_K6_28, u0_K6_29, u0_K6_30, u0_K6_37, u0_K6_38, u0_K6_39, 
       u0_K6_40, u0_K6_42, u0_K7_19, u0_K7_20, u0_K7_21, u0_K7_24, u0_K7_25, u0_K7_26, u0_K7_27, 
       u0_K7_28, u0_K7_29, u0_K7_30, u0_K9_1, u0_K9_10, u0_K9_11, u0_K9_12, u0_K9_13, u0_K9_16, 
       u0_K9_17, u0_K9_18, u0_K9_19, u0_K9_2, u0_K9_20, u0_K9_21, u0_K9_22, u0_K9_23, u0_K9_24, 
       u0_K9_25, u0_K9_26, u0_K9_27, u0_K9_28, u0_K9_29, u0_K9_3, u0_K9_30, u0_K9_43, u0_K9_44, 
       u0_K9_46, u0_K9_47, u0_K9_48, u0_K9_5, u0_K9_7, u0_K9_8, u0_K9_9, u0_out10_14, u0_out10_25, 
       u0_out10_3, u0_out10_8, u0_out12_14, u0_out12_25, u0_out12_3, u0_out12_8, u0_out14_1, u0_out14_10, u0_out14_11, 
       u0_out14_13, u0_out14_16, u0_out14_18, u0_out14_19, u0_out14_2, u0_out14_20, u0_out14_24, u0_out14_26, u0_out14_28, 
       u0_out14_29, u0_out14_30, u0_out14_4, u0_out14_6, u0_out15_11, u0_out15_12, u0_out15_15, u0_out15_19, u0_out15_21, 
       u0_out15_22, u0_out15_27, u0_out15_29, u0_out15_32, u0_out15_4, u0_out15_5, u0_out15_7, u0_out1_15, u0_out1_21, 
       u0_out1_27, u0_out1_5, u0_out5_12, u0_out5_14, u0_out5_22, u0_out5_25, u0_out5_3, u0_out5_32, u0_out5_7, 
       u0_out5_8, u0_out6_1, u0_out6_10, u0_out6_14, u0_out6_20, u0_out6_25, u0_out6_26, u0_out6_3, u0_out6_8, 
       u0_out8_1, u0_out8_10, u0_out8_13, u0_out8_14, u0_out8_15, u0_out8_16, u0_out8_17, u0_out8_18, u0_out8_2, 
       u0_out8_20, u0_out8_21, u0_out8_23, u0_out8_24, u0_out8_25, u0_out8_26, u0_out8_27, u0_out8_28, u0_out8_3, 
       u0_out8_30, u0_out8_31, u0_out8_5, u0_out8_6, u0_out8_8, u0_out8_9, u0_out9_1, u0_out9_10, u0_out9_13, 
       u0_out9_16, u0_out9_18, u0_out9_2, u0_out9_20, u0_out9_24, u0_out9_26, u0_out9_28, u0_out9_30, u0_out9_6, 
       u0_u10_X_25, u0_u10_X_26, u0_u10_X_27, u0_u10_X_28, u0_u10_X_29, u0_u10_X_30, u0_u10_u4_n100, u0_u10_u4_n101, u0_u10_u4_n102, 
       u0_u10_u4_n103, u0_u10_u4_n104, u0_u10_u4_n105, u0_u10_u4_n106, u0_u10_u4_n107, u0_u10_u4_n108, u0_u10_u4_n109, u0_u10_u4_n110, u0_u10_u4_n111, 
       u0_u10_u4_n112, u0_u10_u4_n113, u0_u10_u4_n114, u0_u10_u4_n115, u0_u10_u4_n116, u0_u10_u4_n117, u0_u10_u4_n118, u0_u10_u4_n119, u0_u10_u4_n120, 
       u0_u10_u4_n121, u0_u10_u4_n122, u0_u10_u4_n123, u0_u10_u4_n124, u0_u10_u4_n125, u0_u10_u4_n126, u0_u10_u4_n127, u0_u10_u4_n128, u0_u10_u4_n129, 
       u0_u10_u4_n130, u0_u10_u4_n131, u0_u10_u4_n132, u0_u10_u4_n133, u0_u10_u4_n134, u0_u10_u4_n135, u0_u10_u4_n136, u0_u10_u4_n137, u0_u10_u4_n138, 
       u0_u10_u4_n139, u0_u10_u4_n140, u0_u10_u4_n141, u0_u10_u4_n142, u0_u10_u4_n143, u0_u10_u4_n144, u0_u10_u4_n145, u0_u10_u4_n146, u0_u10_u4_n147, 
       u0_u10_u4_n148, u0_u10_u4_n149, u0_u10_u4_n150, u0_u10_u4_n151, u0_u10_u4_n152, u0_u10_u4_n153, u0_u10_u4_n154, u0_u10_u4_n155, u0_u10_u4_n156, 
       u0_u10_u4_n157, u0_u10_u4_n158, u0_u10_u4_n159, u0_u10_u4_n160, u0_u10_u4_n161, u0_u10_u4_n162, u0_u10_u4_n163, u0_u10_u4_n164, u0_u10_u4_n165, 
       u0_u10_u4_n166, u0_u10_u4_n167, u0_u10_u4_n168, u0_u10_u4_n169, u0_u10_u4_n170, u0_u10_u4_n171, u0_u10_u4_n172, u0_u10_u4_n173, u0_u10_u4_n174, 
       u0_u10_u4_n175, u0_u10_u4_n176, u0_u10_u4_n177, u0_u10_u4_n178, u0_u10_u4_n179, u0_u10_u4_n180, u0_u10_u4_n181, u0_u10_u4_n182, u0_u10_u4_n183, 
       u0_u10_u4_n184, u0_u10_u4_n185, u0_u10_u4_n186, u0_u10_u4_n94, u0_u10_u4_n95, u0_u10_u4_n96, u0_u10_u4_n97, u0_u10_u4_n98, u0_u10_u4_n99, 
       u0_u12_X_25, u0_u12_X_26, u0_u12_X_27, u0_u12_X_28, u0_u12_X_29, u0_u12_X_30, u0_u12_u4_n100, u0_u12_u4_n101, u0_u12_u4_n102, 
       u0_u12_u4_n103, u0_u12_u4_n104, u0_u12_u4_n105, u0_u12_u4_n106, u0_u12_u4_n107, u0_u12_u4_n108, u0_u12_u4_n109, u0_u12_u4_n110, u0_u12_u4_n111, 
       u0_u12_u4_n112, u0_u12_u4_n113, u0_u12_u4_n114, u0_u12_u4_n115, u0_u12_u4_n116, u0_u12_u4_n117, u0_u12_u4_n118, u0_u12_u4_n119, u0_u12_u4_n120, 
       u0_u12_u4_n121, u0_u12_u4_n122, u0_u12_u4_n123, u0_u12_u4_n124, u0_u12_u4_n125, u0_u12_u4_n126, u0_u12_u4_n127, u0_u12_u4_n128, u0_u12_u4_n129, 
       u0_u12_u4_n130, u0_u12_u4_n131, u0_u12_u4_n132, u0_u12_u4_n133, u0_u12_u4_n134, u0_u12_u4_n135, u0_u12_u4_n136, u0_u12_u4_n137, u0_u12_u4_n138, 
       u0_u12_u4_n139, u0_u12_u4_n140, u0_u12_u4_n141, u0_u12_u4_n142, u0_u12_u4_n143, u0_u12_u4_n144, u0_u12_u4_n145, u0_u12_u4_n146, u0_u12_u4_n147, 
       u0_u12_u4_n148, u0_u12_u4_n149, u0_u12_u4_n150, u0_u12_u4_n151, u0_u12_u4_n152, u0_u12_u4_n153, u0_u12_u4_n154, u0_u12_u4_n155, u0_u12_u4_n156, 
       u0_u12_u4_n157, u0_u12_u4_n158, u0_u12_u4_n159, u0_u12_u4_n160, u0_u12_u4_n161, u0_u12_u4_n162, u0_u12_u4_n163, u0_u12_u4_n164, u0_u12_u4_n165, 
       u0_u12_u4_n166, u0_u12_u4_n167, u0_u12_u4_n168, u0_u12_u4_n169, u0_u12_u4_n170, u0_u12_u4_n171, u0_u12_u4_n172, u0_u12_u4_n173, u0_u12_u4_n174, 
       u0_u12_u4_n175, u0_u12_u4_n176, u0_u12_u4_n177, u0_u12_u4_n178, u0_u12_u4_n179, u0_u12_u4_n180, u0_u12_u4_n181, u0_u12_u4_n182, u0_u12_u4_n183, 
       u0_u12_u4_n184, u0_u12_u4_n185, u0_u12_u4_n186, u0_u12_u4_n94, u0_u12_u4_n95, u0_u12_u4_n96, u0_u12_u4_n97, u0_u12_u4_n98, u0_u12_u4_n99, 
       u0_u14_X_10, u0_u14_X_11, u0_u14_X_12, u0_u14_X_13, u0_u14_X_14, u0_u14_X_15, u0_u14_X_16, u0_u14_X_17, u0_u14_X_18, 
       u0_u14_X_19, u0_u14_X_20, u0_u14_X_21, u0_u14_X_22, u0_u14_X_23, u0_u14_X_24, u0_u14_X_31, u0_u14_X_32, u0_u14_X_33, 
       u0_u14_X_34, u0_u14_X_35, u0_u14_X_36, u0_u14_X_7, u0_u14_X_8, u0_u14_X_9, u0_u14_u1_n100, u0_u14_u1_n101, u0_u14_u1_n102, 
       u0_u14_u1_n103, u0_u14_u1_n104, u0_u14_u1_n105, u0_u14_u1_n106, u0_u14_u1_n107, u0_u14_u1_n108, u0_u14_u1_n109, u0_u14_u1_n110, u0_u14_u1_n111, 
       u0_u14_u1_n112, u0_u14_u1_n113, u0_u14_u1_n114, u0_u14_u1_n115, u0_u14_u1_n116, u0_u14_u1_n117, u0_u14_u1_n118, u0_u14_u1_n119, u0_u14_u1_n120, 
       u0_u14_u1_n121, u0_u14_u1_n122, u0_u14_u1_n123, u0_u14_u1_n124, u0_u14_u1_n125, u0_u14_u1_n126, u0_u14_u1_n127, u0_u14_u1_n128, u0_u14_u1_n129, 
       u0_u14_u1_n130, u0_u14_u1_n131, u0_u14_u1_n132, u0_u14_u1_n133, u0_u14_u1_n134, u0_u14_u1_n135, u0_u14_u1_n136, u0_u14_u1_n137, u0_u14_u1_n138, 
       u0_u14_u1_n139, u0_u14_u1_n140, u0_u14_u1_n141, u0_u14_u1_n142, u0_u14_u1_n143, u0_u14_u1_n144, u0_u14_u1_n145, u0_u14_u1_n146, u0_u14_u1_n147, 
       u0_u14_u1_n148, u0_u14_u1_n149, u0_u14_u1_n150, u0_u14_u1_n151, u0_u14_u1_n152, u0_u14_u1_n153, u0_u14_u1_n154, u0_u14_u1_n155, u0_u14_u1_n156, 
       u0_u14_u1_n157, u0_u14_u1_n158, u0_u14_u1_n159, u0_u14_u1_n160, u0_u14_u1_n161, u0_u14_u1_n162, u0_u14_u1_n163, u0_u14_u1_n164, u0_u14_u1_n165, 
       u0_u14_u1_n166, u0_u14_u1_n167, u0_u14_u1_n168, u0_u14_u1_n169, u0_u14_u1_n170, u0_u14_u1_n171, u0_u14_u1_n172, u0_u14_u1_n173, u0_u14_u1_n174, 
       u0_u14_u1_n175, u0_u14_u1_n176, u0_u14_u1_n177, u0_u14_u1_n178, u0_u14_u1_n179, u0_u14_u1_n180, u0_u14_u1_n181, u0_u14_u1_n182, u0_u14_u1_n183, 
       u0_u14_u1_n184, u0_u14_u1_n185, u0_u14_u1_n186, u0_u14_u1_n187, u0_u14_u1_n188, u0_u14_u1_n95, u0_u14_u1_n96, u0_u14_u1_n97, u0_u14_u1_n98, 
       u0_u14_u1_n99, u0_u14_u2_n100, u0_u14_u2_n101, u0_u14_u2_n102, u0_u14_u2_n103, u0_u14_u2_n104, u0_u14_u2_n105, u0_u14_u2_n106, u0_u14_u2_n107, 
       u0_u14_u2_n108, u0_u14_u2_n109, u0_u14_u2_n110, u0_u14_u2_n111, u0_u14_u2_n112, u0_u14_u2_n113, u0_u14_u2_n114, u0_u14_u2_n115, u0_u14_u2_n116, 
       u0_u14_u2_n117, u0_u14_u2_n118, u0_u14_u2_n119, u0_u14_u2_n120, u0_u14_u2_n121, u0_u14_u2_n122, u0_u14_u2_n123, u0_u14_u2_n124, u0_u14_u2_n125, 
       u0_u14_u2_n126, u0_u14_u2_n127, u0_u14_u2_n128, u0_u14_u2_n129, u0_u14_u2_n130, u0_u14_u2_n131, u0_u14_u2_n132, u0_u14_u2_n133, u0_u14_u2_n134, 
       u0_u14_u2_n135, u0_u14_u2_n136, u0_u14_u2_n137, u0_u14_u2_n138, u0_u14_u2_n139, u0_u14_u2_n140, u0_u14_u2_n141, u0_u14_u2_n142, u0_u14_u2_n143, 
       u0_u14_u2_n144, u0_u14_u2_n145, u0_u14_u2_n146, u0_u14_u2_n147, u0_u14_u2_n148, u0_u14_u2_n149, u0_u14_u2_n150, u0_u14_u2_n151, u0_u14_u2_n152, 
       u0_u14_u2_n153, u0_u14_u2_n154, u0_u14_u2_n155, u0_u14_u2_n156, u0_u14_u2_n157, u0_u14_u2_n158, u0_u14_u2_n159, u0_u14_u2_n160, u0_u14_u2_n161, 
       u0_u14_u2_n162, u0_u14_u2_n163, u0_u14_u2_n164, u0_u14_u2_n165, u0_u14_u2_n166, u0_u14_u2_n167, u0_u14_u2_n168, u0_u14_u2_n169, u0_u14_u2_n170, 
       u0_u14_u2_n171, u0_u14_u2_n172, u0_u14_u2_n173, u0_u14_u2_n174, u0_u14_u2_n175, u0_u14_u2_n176, u0_u14_u2_n177, u0_u14_u2_n178, u0_u14_u2_n179, 
       u0_u14_u2_n180, u0_u14_u2_n181, u0_u14_u2_n182, u0_u14_u2_n183, u0_u14_u2_n184, u0_u14_u2_n185, u0_u14_u2_n186, u0_u14_u2_n187, u0_u14_u2_n188, 
       u0_u14_u2_n95, u0_u14_u2_n96, u0_u14_u2_n97, u0_u14_u2_n98, u0_u14_u2_n99, u0_u14_u3_n100, u0_u14_u3_n101, u0_u14_u3_n102, u0_u14_u3_n103, 
       u0_u14_u3_n104, u0_u14_u3_n105, u0_u14_u3_n106, u0_u14_u3_n107, u0_u14_u3_n108, u0_u14_u3_n109, u0_u14_u3_n110, u0_u14_u3_n111, u0_u14_u3_n112, 
       u0_u14_u3_n113, u0_u14_u3_n114, u0_u14_u3_n115, u0_u14_u3_n116, u0_u14_u3_n117, u0_u14_u3_n118, u0_u14_u3_n119, u0_u14_u3_n120, u0_u14_u3_n121, 
       u0_u14_u3_n122, u0_u14_u3_n123, u0_u14_u3_n124, u0_u14_u3_n125, u0_u14_u3_n126, u0_u14_u3_n127, u0_u14_u3_n128, u0_u14_u3_n129, u0_u14_u3_n130, 
       u0_u14_u3_n131, u0_u14_u3_n132, u0_u14_u3_n133, u0_u14_u3_n134, u0_u14_u3_n135, u0_u14_u3_n136, u0_u14_u3_n137, u0_u14_u3_n138, u0_u14_u3_n139, 
       u0_u14_u3_n140, u0_u14_u3_n141, u0_u14_u3_n142, u0_u14_u3_n143, u0_u14_u3_n144, u0_u14_u3_n145, u0_u14_u3_n146, u0_u14_u3_n147, u0_u14_u3_n148, 
       u0_u14_u3_n149, u0_u14_u3_n150, u0_u14_u3_n151, u0_u14_u3_n152, u0_u14_u3_n153, u0_u14_u3_n154, u0_u14_u3_n155, u0_u14_u3_n156, u0_u14_u3_n157, 
       u0_u14_u3_n158, u0_u14_u3_n159, u0_u14_u3_n160, u0_u14_u3_n161, u0_u14_u3_n162, u0_u14_u3_n163, u0_u14_u3_n164, u0_u14_u3_n165, u0_u14_u3_n166, 
       u0_u14_u3_n167, u0_u14_u3_n168, u0_u14_u3_n169, u0_u14_u3_n170, u0_u14_u3_n171, u0_u14_u3_n172, u0_u14_u3_n173, u0_u14_u3_n174, u0_u14_u3_n175, 
       u0_u14_u3_n176, u0_u14_u3_n177, u0_u14_u3_n178, u0_u14_u3_n179, u0_u14_u3_n180, u0_u14_u3_n181, u0_u14_u3_n182, u0_u14_u3_n183, u0_u14_u3_n184, 
       u0_u14_u3_n185, u0_u14_u3_n186, u0_u14_u3_n94, u0_u14_u3_n95, u0_u14_u3_n96, u0_u14_u3_n97, u0_u14_u3_n98, u0_u14_u3_n99, u0_u14_u5_n100, 
       u0_u14_u5_n101, u0_u14_u5_n102, u0_u14_u5_n103, u0_u14_u5_n104, u0_u14_u5_n105, u0_u14_u5_n106, u0_u14_u5_n107, u0_u14_u5_n108, u0_u14_u5_n109, 
       u0_u14_u5_n110, u0_u14_u5_n111, u0_u14_u5_n112, u0_u14_u5_n113, u0_u14_u5_n114, u0_u14_u5_n115, u0_u14_u5_n116, u0_u14_u5_n117, u0_u14_u5_n118, 
       u0_u14_u5_n119, u0_u14_u5_n120, u0_u14_u5_n121, u0_u14_u5_n122, u0_u14_u5_n123, u0_u14_u5_n124, u0_u14_u5_n125, u0_u14_u5_n126, u0_u14_u5_n127, 
       u0_u14_u5_n128, u0_u14_u5_n129, u0_u14_u5_n130, u0_u14_u5_n131, u0_u14_u5_n132, u0_u14_u5_n133, u0_u14_u5_n134, u0_u14_u5_n135, u0_u14_u5_n136, 
       u0_u14_u5_n137, u0_u14_u5_n138, u0_u14_u5_n139, u0_u14_u5_n140, u0_u14_u5_n141, u0_u14_u5_n142, u0_u14_u5_n143, u0_u14_u5_n144, u0_u14_u5_n145, 
       u0_u14_u5_n146, u0_u14_u5_n147, u0_u14_u5_n148, u0_u14_u5_n149, u0_u14_u5_n150, u0_u14_u5_n151, u0_u14_u5_n152, u0_u14_u5_n153, u0_u14_u5_n154, 
       u0_u14_u5_n155, u0_u14_u5_n156, u0_u14_u5_n157, u0_u14_u5_n158, u0_u14_u5_n159, u0_u14_u5_n160, u0_u14_u5_n161, u0_u14_u5_n162, u0_u14_u5_n163, 
       u0_u14_u5_n164, u0_u14_u5_n165, u0_u14_u5_n166, u0_u14_u5_n167, u0_u14_u5_n168, u0_u14_u5_n169, u0_u14_u5_n170, u0_u14_u5_n171, u0_u14_u5_n172, 
       u0_u14_u5_n173, u0_u14_u5_n174, u0_u14_u5_n175, u0_u14_u5_n176, u0_u14_u5_n177, u0_u14_u5_n178, u0_u14_u5_n179, u0_u14_u5_n180, u0_u14_u5_n181, 
       u0_u14_u5_n182, u0_u14_u5_n183, u0_u14_u5_n184, u0_u14_u5_n185, u0_u14_u5_n186, u0_u14_u5_n187, u0_u14_u5_n188, u0_u14_u5_n189, u0_u14_u5_n190, 
       u0_u14_u5_n191, u0_u14_u5_n192, u0_u14_u5_n193, u0_u14_u5_n194, u0_u14_u5_n195, u0_u14_u5_n196, u0_u14_u5_n99, u0_u15_X_31, u0_u15_X_32, 
       u0_u15_X_33, u0_u15_X_34, u0_u15_X_35, u0_u15_X_36, u0_u15_X_37, u0_u15_X_38, u0_u15_X_39, u0_u15_X_40, u0_u15_X_41, 
       u0_u15_X_42, u0_u15_X_43, u0_u15_X_44, u0_u15_X_45, u0_u15_X_46, u0_u15_X_47, u0_u15_X_48, u0_u15_u5_n100, u0_u15_u5_n101, 
       u0_u15_u5_n102, u0_u15_u5_n103, u0_u15_u5_n104, u0_u15_u5_n105, u0_u15_u5_n106, u0_u15_u5_n107, u0_u15_u5_n108, u0_u15_u5_n109, u0_u15_u5_n110, 
       u0_u15_u5_n111, u0_u15_u5_n112, u0_u15_u5_n113, u0_u15_u5_n114, u0_u15_u5_n115, u0_u15_u5_n116, u0_u15_u5_n117, u0_u15_u5_n118, u0_u15_u5_n119, 
       u0_u15_u5_n120, u0_u15_u5_n121, u0_u15_u5_n122, u0_u15_u5_n123, u0_u15_u5_n124, u0_u15_u5_n125, u0_u15_u5_n126, u0_u15_u5_n127, u0_u15_u5_n128, 
       u0_u15_u5_n129, u0_u15_u5_n130, u0_u15_u5_n131, u0_u15_u5_n132, u0_u15_u5_n133, u0_u15_u5_n134, u0_u15_u5_n135, u0_u15_u5_n136, u0_u15_u5_n137, 
       u0_u15_u5_n138, u0_u15_u5_n139, u0_u15_u5_n140, u0_u15_u5_n141, u0_u15_u5_n142, u0_u15_u5_n143, u0_u15_u5_n144, u0_u15_u5_n145, u0_u15_u5_n146, 
       u0_u15_u5_n147, u0_u15_u5_n148, u0_u15_u5_n149, u0_u15_u5_n150, u0_u15_u5_n151, u0_u15_u5_n152, u0_u15_u5_n153, u0_u15_u5_n154, u0_u15_u5_n155, 
       u0_u15_u5_n156, u0_u15_u5_n157, u0_u15_u5_n158, u0_u15_u5_n159, u0_u15_u5_n160, u0_u15_u5_n161, u0_u15_u5_n162, u0_u15_u5_n163, u0_u15_u5_n164, 
       u0_u15_u5_n165, u0_u15_u5_n166, u0_u15_u5_n167, u0_u15_u5_n168, u0_u15_u5_n169, u0_u15_u5_n170, u0_u15_u5_n171, u0_u15_u5_n172, u0_u15_u5_n173, 
       u0_u15_u5_n174, u0_u15_u5_n175, u0_u15_u5_n176, u0_u15_u5_n177, u0_u15_u5_n178, u0_u15_u5_n179, u0_u15_u5_n180, u0_u15_u5_n181, u0_u15_u5_n182, 
       u0_u15_u5_n183, u0_u15_u5_n184, u0_u15_u5_n185, u0_u15_u5_n186, u0_u15_u5_n187, u0_u15_u5_n188, u0_u15_u5_n189, u0_u15_u5_n190, u0_u15_u5_n191, 
       u0_u15_u5_n192, u0_u15_u5_n193, u0_u15_u5_n194, u0_u15_u5_n195, u0_u15_u5_n196, u0_u15_u5_n99, u0_u15_u6_n100, u0_u15_u6_n101, u0_u15_u6_n102, 
       u0_u15_u6_n103, u0_u15_u6_n104, u0_u15_u6_n105, u0_u15_u6_n106, u0_u15_u6_n107, u0_u15_u6_n108, u0_u15_u6_n109, u0_u15_u6_n110, u0_u15_u6_n111, 
       u0_u15_u6_n112, u0_u15_u6_n113, u0_u15_u6_n114, u0_u15_u6_n115, u0_u15_u6_n116, u0_u15_u6_n117, u0_u15_u6_n118, u0_u15_u6_n119, u0_u15_u6_n120, 
       u0_u15_u6_n121, u0_u15_u6_n122, u0_u15_u6_n123, u0_u15_u6_n124, u0_u15_u6_n125, u0_u15_u6_n126, u0_u15_u6_n127, u0_u15_u6_n128, u0_u15_u6_n129, 
       u0_u15_u6_n130, u0_u15_u6_n131, u0_u15_u6_n132, u0_u15_u6_n133, u0_u15_u6_n134, u0_u15_u6_n135, u0_u15_u6_n136, u0_u15_u6_n137, u0_u15_u6_n138, 
       u0_u15_u6_n139, u0_u15_u6_n140, u0_u15_u6_n141, u0_u15_u6_n142, u0_u15_u6_n143, u0_u15_u6_n144, u0_u15_u6_n145, u0_u15_u6_n146, u0_u15_u6_n147, 
       u0_u15_u6_n148, u0_u15_u6_n149, u0_u15_u6_n150, u0_u15_u6_n151, u0_u15_u6_n152, u0_u15_u6_n153, u0_u15_u6_n154, u0_u15_u6_n155, u0_u15_u6_n156, 
       u0_u15_u6_n157, u0_u15_u6_n158, u0_u15_u6_n159, u0_u15_u6_n160, u0_u15_u6_n161, u0_u15_u6_n162, u0_u15_u6_n163, u0_u15_u6_n164, u0_u15_u6_n165, 
       u0_u15_u6_n166, u0_u15_u6_n167, u0_u15_u6_n168, u0_u15_u6_n169, u0_u15_u6_n170, u0_u15_u6_n171, u0_u15_u6_n172, u0_u15_u6_n173, u0_u15_u6_n174, 
       u0_u15_u6_n88, u0_u15_u6_n89, u0_u15_u6_n90, u0_u15_u6_n91, u0_u15_u6_n92, u0_u15_u6_n93, u0_u15_u6_n94, u0_u15_u6_n95, u0_u15_u6_n96, 
       u0_u15_u6_n97, u0_u15_u6_n98, u0_u15_u6_n99, u0_u15_u7_n100, u0_u15_u7_n101, u0_u15_u7_n102, u0_u15_u7_n103, u0_u15_u7_n104, u0_u15_u7_n105, 
       u0_u15_u7_n106, u0_u15_u7_n107, u0_u15_u7_n108, u0_u15_u7_n109, u0_u15_u7_n110, u0_u15_u7_n111, u0_u15_u7_n112, u0_u15_u7_n113, u0_u15_u7_n114, 
       u0_u15_u7_n115, u0_u15_u7_n116, u0_u15_u7_n117, u0_u15_u7_n118, u0_u15_u7_n119, u0_u15_u7_n120, u0_u15_u7_n121, u0_u15_u7_n122, u0_u15_u7_n123, 
       u0_u15_u7_n124, u0_u15_u7_n125, u0_u15_u7_n126, u0_u15_u7_n127, u0_u15_u7_n128, u0_u15_u7_n129, u0_u15_u7_n130, u0_u15_u7_n131, u0_u15_u7_n132, 
       u0_u15_u7_n133, u0_u15_u7_n134, u0_u15_u7_n135, u0_u15_u7_n136, u0_u15_u7_n137, u0_u15_u7_n138, u0_u15_u7_n139, u0_u15_u7_n140, u0_u15_u7_n141, 
       u0_u15_u7_n142, u0_u15_u7_n143, u0_u15_u7_n144, u0_u15_u7_n145, u0_u15_u7_n146, u0_u15_u7_n147, u0_u15_u7_n148, u0_u15_u7_n149, u0_u15_u7_n150, 
       u0_u15_u7_n151, u0_u15_u7_n152, u0_u15_u7_n153, u0_u15_u7_n154, u0_u15_u7_n155, u0_u15_u7_n156, u0_u15_u7_n157, u0_u15_u7_n158, u0_u15_u7_n159, 
       u0_u15_u7_n160, u0_u15_u7_n161, u0_u15_u7_n162, u0_u15_u7_n163, u0_u15_u7_n164, u0_u15_u7_n165, u0_u15_u7_n166, u0_u15_u7_n167, u0_u15_u7_n168, 
       u0_u15_u7_n169, u0_u15_u7_n170, u0_u15_u7_n171, u0_u15_u7_n172, u0_u15_u7_n173, u0_u15_u7_n174, u0_u15_u7_n175, u0_u15_u7_n176, u0_u15_u7_n177, 
       u0_u15_u7_n178, u0_u15_u7_n179, u0_u15_u7_n180, u0_u15_u7_n91, u0_u15_u7_n92, u0_u15_u7_n93, u0_u15_u7_n94, u0_u15_u7_n95, u0_u15_u7_n96, 
       u0_u15_u7_n97, u0_u15_u7_n98, u0_u15_u7_n99, u0_u1_X_43, u0_u1_X_44, u0_u1_X_45, u0_u1_X_46, u0_u1_X_47, u0_u1_X_48, 
       u0_u1_u7_n100, u0_u1_u7_n101, u0_u1_u7_n102, u0_u1_u7_n103, u0_u1_u7_n104, u0_u1_u7_n105, u0_u1_u7_n106, u0_u1_u7_n107, u0_u1_u7_n108, 
       u0_u1_u7_n109, u0_u1_u7_n110, u0_u1_u7_n111, u0_u1_u7_n112, u0_u1_u7_n113, u0_u1_u7_n114, u0_u1_u7_n115, u0_u1_u7_n116, u0_u1_u7_n117, 
       u0_u1_u7_n118, u0_u1_u7_n119, u0_u1_u7_n120, u0_u1_u7_n121, u0_u1_u7_n122, u0_u1_u7_n123, u0_u1_u7_n124, u0_u1_u7_n125, u0_u1_u7_n126, 
       u0_u1_u7_n127, u0_u1_u7_n128, u0_u1_u7_n129, u0_u1_u7_n130, u0_u1_u7_n131, u0_u1_u7_n132, u0_u1_u7_n133, u0_u1_u7_n134, u0_u1_u7_n135, 
       u0_u1_u7_n136, u0_u1_u7_n137, u0_u1_u7_n138, u0_u1_u7_n139, u0_u1_u7_n140, u0_u1_u7_n141, u0_u1_u7_n142, u0_u1_u7_n143, u0_u1_u7_n144, 
       u0_u1_u7_n145, u0_u1_u7_n146, u0_u1_u7_n147, u0_u1_u7_n148, u0_u1_u7_n149, u0_u1_u7_n150, u0_u1_u7_n151, u0_u1_u7_n152, u0_u1_u7_n153, 
       u0_u1_u7_n154, u0_u1_u7_n155, u0_u1_u7_n156, u0_u1_u7_n157, u0_u1_u7_n158, u0_u1_u7_n159, u0_u1_u7_n160, u0_u1_u7_n161, u0_u1_u7_n162, 
       u0_u1_u7_n163, u0_u1_u7_n164, u0_u1_u7_n165, u0_u1_u7_n166, u0_u1_u7_n167, u0_u1_u7_n168, u0_u1_u7_n169, u0_u1_u7_n170, u0_u1_u7_n171, 
       u0_u1_u7_n172, u0_u1_u7_n173, u0_u1_u7_n174, u0_u1_u7_n175, u0_u1_u7_n176, u0_u1_u7_n177, u0_u1_u7_n178, u0_u1_u7_n179, u0_u1_u7_n180, 
       u0_u1_u7_n91, u0_u1_u7_n92, u0_u1_u7_n93, u0_u1_u7_n94, u0_u1_u7_n95, u0_u1_u7_n96, u0_u1_u7_n97, u0_u1_u7_n98, u0_u1_u7_n99, 
       u0_u5_X_25, u0_u5_X_26, u0_u5_X_27, u0_u5_X_28, u0_u5_X_29, u0_u5_X_30, u0_u5_X_37, u0_u5_X_38, u0_u5_X_39, 
       u0_u5_X_40, u0_u5_X_41, u0_u5_X_42, u0_u5_u4_n100, u0_u5_u4_n101, u0_u5_u4_n102, u0_u5_u4_n103, u0_u5_u4_n104, u0_u5_u4_n105, 
       u0_u5_u4_n106, u0_u5_u4_n107, u0_u5_u4_n108, u0_u5_u4_n109, u0_u5_u4_n110, u0_u5_u4_n111, u0_u5_u4_n112, u0_u5_u4_n113, u0_u5_u4_n114, 
       u0_u5_u4_n115, u0_u5_u4_n116, u0_u5_u4_n117, u0_u5_u4_n118, u0_u5_u4_n119, u0_u5_u4_n120, u0_u5_u4_n121, u0_u5_u4_n122, u0_u5_u4_n123, 
       u0_u5_u4_n124, u0_u5_u4_n125, u0_u5_u4_n126, u0_u5_u4_n127, u0_u5_u4_n128, u0_u5_u4_n129, u0_u5_u4_n130, u0_u5_u4_n131, u0_u5_u4_n132, 
       u0_u5_u4_n133, u0_u5_u4_n134, u0_u5_u4_n135, u0_u5_u4_n136, u0_u5_u4_n137, u0_u5_u4_n138, u0_u5_u4_n139, u0_u5_u4_n140, u0_u5_u4_n141, 
       u0_u5_u4_n142, u0_u5_u4_n143, u0_u5_u4_n144, u0_u5_u4_n145, u0_u5_u4_n146, u0_u5_u4_n147, u0_u5_u4_n148, u0_u5_u4_n149, u0_u5_u4_n150, 
       u0_u5_u4_n151, u0_u5_u4_n152, u0_u5_u4_n153, u0_u5_u4_n154, u0_u5_u4_n155, u0_u5_u4_n156, u0_u5_u4_n157, u0_u5_u4_n158, u0_u5_u4_n159, 
       u0_u5_u4_n160, u0_u5_u4_n161, u0_u5_u4_n162, u0_u5_u4_n163, u0_u5_u4_n164, u0_u5_u4_n165, u0_u5_u4_n166, u0_u5_u4_n167, u0_u5_u4_n168, 
       u0_u5_u4_n169, u0_u5_u4_n170, u0_u5_u4_n171, u0_u5_u4_n172, u0_u5_u4_n173, u0_u5_u4_n174, u0_u5_u4_n175, u0_u5_u4_n176, u0_u5_u4_n177, 
       u0_u5_u4_n178, u0_u5_u4_n179, u0_u5_u4_n180, u0_u5_u4_n181, u0_u5_u4_n182, u0_u5_u4_n183, u0_u5_u4_n184, u0_u5_u4_n185, u0_u5_u4_n186, 
       u0_u5_u4_n94, u0_u5_u4_n95, u0_u5_u4_n96, u0_u5_u4_n97, u0_u5_u4_n98, u0_u5_u4_n99, u0_u5_u6_n100, u0_u5_u6_n101, u0_u5_u6_n102, 
       u0_u5_u6_n103, u0_u5_u6_n104, u0_u5_u6_n105, u0_u5_u6_n106, u0_u5_u6_n107, u0_u5_u6_n108, u0_u5_u6_n109, u0_u5_u6_n110, u0_u5_u6_n111, 
       u0_u5_u6_n112, u0_u5_u6_n113, u0_u5_u6_n114, u0_u5_u6_n115, u0_u5_u6_n116, u0_u5_u6_n117, u0_u5_u6_n118, u0_u5_u6_n119, u0_u5_u6_n120, 
       u0_u5_u6_n121, u0_u5_u6_n122, u0_u5_u6_n123, u0_u5_u6_n124, u0_u5_u6_n125, u0_u5_u6_n126, u0_u5_u6_n127, u0_u5_u6_n128, u0_u5_u6_n129, 
       u0_u5_u6_n130, u0_u5_u6_n131, u0_u5_u6_n132, u0_u5_u6_n133, u0_u5_u6_n134, u0_u5_u6_n135, u0_u5_u6_n136, u0_u5_u6_n137, u0_u5_u6_n138, 
       u0_u5_u6_n139, u0_u5_u6_n140, u0_u5_u6_n141, u0_u5_u6_n142, u0_u5_u6_n143, u0_u5_u6_n144, u0_u5_u6_n145, u0_u5_u6_n146, u0_u5_u6_n147, 
       u0_u5_u6_n148, u0_u5_u6_n149, u0_u5_u6_n150, u0_u5_u6_n151, u0_u5_u6_n152, u0_u5_u6_n153, u0_u5_u6_n154, u0_u5_u6_n155, u0_u5_u6_n156, 
       u0_u5_u6_n157, u0_u5_u6_n158, u0_u5_u6_n159, u0_u5_u6_n160, u0_u5_u6_n161, u0_u5_u6_n162, u0_u5_u6_n163, u0_u5_u6_n164, u0_u5_u6_n165, 
       u0_u5_u6_n166, u0_u5_u6_n167, u0_u5_u6_n168, u0_u5_u6_n169, u0_u5_u6_n170, u0_u5_u6_n171, u0_u5_u6_n172, u0_u5_u6_n173, u0_u5_u6_n174, 
       u0_u5_u6_n88, u0_u5_u6_n89, u0_u5_u6_n90, u0_u5_u6_n91, u0_u5_u6_n92, u0_u5_u6_n93, u0_u5_u6_n94, u0_u5_u6_n95, u0_u5_u6_n96, 
       u0_u5_u6_n97, u0_u5_u6_n98, u0_u5_u6_n99, u0_u6_X_19, u0_u6_X_20, u0_u6_X_21, u0_u6_X_22, u0_u6_X_23, u0_u6_X_24, 
       u0_u6_X_25, u0_u6_X_26, u0_u6_X_27, u0_u6_X_28, u0_u6_X_29, u0_u6_X_30, u0_u6_u3_n100, u0_u6_u3_n101, u0_u6_u3_n102, 
       u0_u6_u3_n103, u0_u6_u3_n104, u0_u6_u3_n105, u0_u6_u3_n106, u0_u6_u3_n107, u0_u6_u3_n108, u0_u6_u3_n109, u0_u6_u3_n110, u0_u6_u3_n111, 
       u0_u6_u3_n112, u0_u6_u3_n113, u0_u6_u3_n114, u0_u6_u3_n115, u0_u6_u3_n116, u0_u6_u3_n117, u0_u6_u3_n118, u0_u6_u3_n119, u0_u6_u3_n120, 
       u0_u6_u3_n121, u0_u6_u3_n122, u0_u6_u3_n123, u0_u6_u3_n124, u0_u6_u3_n125, u0_u6_u3_n126, u0_u6_u3_n127, u0_u6_u3_n128, u0_u6_u3_n129, 
       u0_u6_u3_n130, u0_u6_u3_n131, u0_u6_u3_n132, u0_u6_u3_n133, u0_u6_u3_n134, u0_u6_u3_n135, u0_u6_u3_n136, u0_u6_u3_n137, u0_u6_u3_n138, 
       u0_u6_u3_n139, u0_u6_u3_n140, u0_u6_u3_n141, u0_u6_u3_n142, u0_u6_u3_n143, u0_u6_u3_n144, u0_u6_u3_n145, u0_u6_u3_n146, u0_u6_u3_n147, 
       u0_u6_u3_n148, u0_u6_u3_n149, u0_u6_u3_n150, u0_u6_u3_n151, u0_u6_u3_n152, u0_u6_u3_n153, u0_u6_u3_n154, u0_u6_u3_n155, u0_u6_u3_n156, 
       u0_u6_u3_n157, u0_u6_u3_n158, u0_u6_u3_n159, u0_u6_u3_n160, u0_u6_u3_n161, u0_u6_u3_n162, u0_u6_u3_n163, u0_u6_u3_n164, u0_u6_u3_n165, 
       u0_u6_u3_n166, u0_u6_u3_n167, u0_u6_u3_n168, u0_u6_u3_n169, u0_u6_u3_n170, u0_u6_u3_n171, u0_u6_u3_n172, u0_u6_u3_n173, u0_u6_u3_n174, 
       u0_u6_u3_n175, u0_u6_u3_n176, u0_u6_u3_n177, u0_u6_u3_n178, u0_u6_u3_n179, u0_u6_u3_n180, u0_u6_u3_n181, u0_u6_u3_n182, u0_u6_u3_n183, 
       u0_u6_u3_n184, u0_u6_u3_n185, u0_u6_u3_n186, u0_u6_u3_n94, u0_u6_u3_n95, u0_u6_u3_n96, u0_u6_u3_n97, u0_u6_u3_n98, u0_u6_u3_n99, 
       u0_u6_u4_n100, u0_u6_u4_n101, u0_u6_u4_n102, u0_u6_u4_n103, u0_u6_u4_n104, u0_u6_u4_n105, u0_u6_u4_n106, u0_u6_u4_n107, u0_u6_u4_n108, 
       u0_u6_u4_n109, u0_u6_u4_n110, u0_u6_u4_n111, u0_u6_u4_n112, u0_u6_u4_n113, u0_u6_u4_n114, u0_u6_u4_n115, u0_u6_u4_n116, u0_u6_u4_n117, 
       u0_u6_u4_n118, u0_u6_u4_n119, u0_u6_u4_n120, u0_u6_u4_n121, u0_u6_u4_n122, u0_u6_u4_n123, u0_u6_u4_n124, u0_u6_u4_n125, u0_u6_u4_n126, 
       u0_u6_u4_n127, u0_u6_u4_n128, u0_u6_u4_n129, u0_u6_u4_n130, u0_u6_u4_n131, u0_u6_u4_n132, u0_u6_u4_n133, u0_u6_u4_n134, u0_u6_u4_n135, 
       u0_u6_u4_n136, u0_u6_u4_n137, u0_u6_u4_n138, u0_u6_u4_n139, u0_u6_u4_n140, u0_u6_u4_n141, u0_u6_u4_n142, u0_u6_u4_n143, u0_u6_u4_n144, 
       u0_u6_u4_n145, u0_u6_u4_n146, u0_u6_u4_n147, u0_u6_u4_n148, u0_u6_u4_n149, u0_u6_u4_n150, u0_u6_u4_n151, u0_u6_u4_n152, u0_u6_u4_n153, 
       u0_u6_u4_n154, u0_u6_u4_n155, u0_u6_u4_n156, u0_u6_u4_n157, u0_u6_u4_n158, u0_u6_u4_n159, u0_u6_u4_n160, u0_u6_u4_n161, u0_u6_u4_n162, 
       u0_u6_u4_n163, u0_u6_u4_n164, u0_u6_u4_n165, u0_u6_u4_n166, u0_u6_u4_n167, u0_u6_u4_n168, u0_u6_u4_n169, u0_u6_u4_n170, u0_u6_u4_n171, 
       u0_u6_u4_n172, u0_u6_u4_n173, u0_u6_u4_n174, u0_u6_u4_n175, u0_u6_u4_n176, u0_u6_u4_n177, u0_u6_u4_n178, u0_u6_u4_n179, u0_u6_u4_n180, 
       u0_u6_u4_n181, u0_u6_u4_n182, u0_u6_u4_n183, u0_u6_u4_n184, u0_u6_u4_n185, u0_u6_u4_n186, u0_u6_u4_n94, u0_u6_u4_n95, u0_u6_u4_n96, 
       u0_u6_u4_n97, u0_u6_u4_n98, u0_u6_u4_n99, u0_u8_X_1, u0_u8_X_10, u0_u8_X_11, u0_u8_X_12, u0_u8_X_13, u0_u8_X_14, 
       u0_u8_X_15, u0_u8_X_16, u0_u8_X_17, u0_u8_X_18, u0_u8_X_19, u0_u8_X_2, u0_u8_X_20, u0_u8_X_21, u0_u8_X_22, 
       u0_u8_X_23, u0_u8_X_24, u0_u8_X_25, u0_u8_X_26, u0_u8_X_27, u0_u8_X_28, u0_u8_X_29, u0_u8_X_3, u0_u8_X_30, 
       u0_u8_X_4, u0_u8_X_43, u0_u8_X_44, u0_u8_X_45, u0_u8_X_46, u0_u8_X_47, u0_u8_X_48, u0_u8_X_5, u0_u8_X_6, 
       u0_u8_X_7, u0_u8_X_8, u0_u8_X_9, u0_u8_u0_n100, u0_u8_u0_n101, u0_u8_u0_n102, u0_u8_u0_n103, u0_u8_u0_n104, u0_u8_u0_n105, 
       u0_u8_u0_n106, u0_u8_u0_n107, u0_u8_u0_n108, u0_u8_u0_n109, u0_u8_u0_n110, u0_u8_u0_n111, u0_u8_u0_n112, u0_u8_u0_n113, u0_u8_u0_n114, 
       u0_u8_u0_n115, u0_u8_u0_n116, u0_u8_u0_n117, u0_u8_u0_n118, u0_u8_u0_n119, u0_u8_u0_n120, u0_u8_u0_n121, u0_u8_u0_n122, u0_u8_u0_n123, 
       u0_u8_u0_n124, u0_u8_u0_n125, u0_u8_u0_n126, u0_u8_u0_n127, u0_u8_u0_n128, u0_u8_u0_n129, u0_u8_u0_n130, u0_u8_u0_n131, u0_u8_u0_n132, 
       u0_u8_u0_n133, u0_u8_u0_n134, u0_u8_u0_n135, u0_u8_u0_n136, u0_u8_u0_n137, u0_u8_u0_n138, u0_u8_u0_n139, u0_u8_u0_n140, u0_u8_u0_n141, 
       u0_u8_u0_n142, u0_u8_u0_n143, u0_u8_u0_n144, u0_u8_u0_n145, u0_u8_u0_n146, u0_u8_u0_n147, u0_u8_u0_n148, u0_u8_u0_n149, u0_u8_u0_n150, 
       u0_u8_u0_n151, u0_u8_u0_n152, u0_u8_u0_n153, u0_u8_u0_n154, u0_u8_u0_n155, u0_u8_u0_n156, u0_u8_u0_n157, u0_u8_u0_n158, u0_u8_u0_n159, 
       u0_u8_u0_n160, u0_u8_u0_n161, u0_u8_u0_n162, u0_u8_u0_n163, u0_u8_u0_n164, u0_u8_u0_n165, u0_u8_u0_n166, u0_u8_u0_n167, u0_u8_u0_n168, 
       u0_u8_u0_n169, u0_u8_u0_n170, u0_u8_u0_n171, u0_u8_u0_n172, u0_u8_u0_n173, u0_u8_u0_n174, u0_u8_u0_n88, u0_u8_u0_n89, u0_u8_u0_n90, 
       u0_u8_u0_n91, u0_u8_u0_n92, u0_u8_u0_n93, u0_u8_u0_n94, u0_u8_u0_n95, u0_u8_u0_n96, u0_u8_u0_n97, u0_u8_u0_n98, u0_u8_u0_n99, 
       u0_u8_u1_n100, u0_u8_u1_n101, u0_u8_u1_n102, u0_u8_u1_n103, u0_u8_u1_n104, u0_u8_u1_n105, u0_u8_u1_n106, u0_u8_u1_n107, u0_u8_u1_n108, 
       u0_u8_u1_n109, u0_u8_u1_n110, u0_u8_u1_n111, u0_u8_u1_n112, u0_u8_u1_n113, u0_u8_u1_n114, u0_u8_u1_n115, u0_u8_u1_n116, u0_u8_u1_n117, 
       u0_u8_u1_n118, u0_u8_u1_n119, u0_u8_u1_n120, u0_u8_u1_n121, u0_u8_u1_n122, u0_u8_u1_n123, u0_u8_u1_n124, u0_u8_u1_n125, u0_u8_u1_n126, 
       u0_u8_u1_n127, u0_u8_u1_n128, u0_u8_u1_n129, u0_u8_u1_n130, u0_u8_u1_n131, u0_u8_u1_n132, u0_u8_u1_n133, u0_u8_u1_n134, u0_u8_u1_n135, 
       u0_u8_u1_n136, u0_u8_u1_n137, u0_u8_u1_n138, u0_u8_u1_n139, u0_u8_u1_n140, u0_u8_u1_n141, u0_u8_u1_n142, u0_u8_u1_n143, u0_u8_u1_n144, 
       u0_u8_u1_n145, u0_u8_u1_n146, u0_u8_u1_n147, u0_u8_u1_n148, u0_u8_u1_n149, u0_u8_u1_n150, u0_u8_u1_n151, u0_u8_u1_n152, u0_u8_u1_n153, 
       u0_u8_u1_n154, u0_u8_u1_n155, u0_u8_u1_n156, u0_u8_u1_n157, u0_u8_u1_n158, u0_u8_u1_n159, u0_u8_u1_n160, u0_u8_u1_n161, u0_u8_u1_n162, 
       u0_u8_u1_n163, u0_u8_u1_n164, u0_u8_u1_n165, u0_u8_u1_n166, u0_u8_u1_n167, u0_u8_u1_n168, u0_u8_u1_n169, u0_u8_u1_n170, u0_u8_u1_n171, 
       u0_u8_u1_n172, u0_u8_u1_n173, u0_u8_u1_n174, u0_u8_u1_n175, u0_u8_u1_n176, u0_u8_u1_n177, u0_u8_u1_n178, u0_u8_u1_n179, u0_u8_u1_n180, 
       u0_u8_u1_n181, u0_u8_u1_n182, u0_u8_u1_n183, u0_u8_u1_n184, u0_u8_u1_n185, u0_u8_u1_n186, u0_u8_u1_n187, u0_u8_u1_n188, u0_u8_u1_n95, 
       u0_u8_u1_n96, u0_u8_u1_n97, u0_u8_u1_n98, u0_u8_u1_n99, u0_u8_u2_n100, u0_u8_u2_n101, u0_u8_u2_n102, u0_u8_u2_n103, u0_u8_u2_n104, 
       u0_u8_u2_n105, u0_u8_u2_n106, u0_u8_u2_n107, u0_u8_u2_n108, u0_u8_u2_n109, u0_u8_u2_n110, u0_u8_u2_n111, u0_u8_u2_n112, u0_u8_u2_n113, 
       u0_u8_u2_n114, u0_u8_u2_n115, u0_u8_u2_n116, u0_u8_u2_n117, u0_u8_u2_n118, u0_u8_u2_n119, u0_u8_u2_n120, u0_u8_u2_n121, u0_u8_u2_n122, 
       u0_u8_u2_n123, u0_u8_u2_n124, u0_u8_u2_n125, u0_u8_u2_n126, u0_u8_u2_n127, u0_u8_u2_n128, u0_u8_u2_n129, u0_u8_u2_n130, u0_u8_u2_n131, 
       u0_u8_u2_n132, u0_u8_u2_n133, u0_u8_u2_n134, u0_u8_u2_n135, u0_u8_u2_n136, u0_u8_u2_n137, u0_u8_u2_n138, u0_u8_u2_n139, u0_u8_u2_n140, 
       u0_u8_u2_n141, u0_u8_u2_n142, u0_u8_u2_n143, u0_u8_u2_n144, u0_u8_u2_n145, u0_u8_u2_n146, u0_u8_u2_n147, u0_u8_u2_n148, u0_u8_u2_n149, 
       u0_u8_u2_n150, u0_u8_u2_n151, u0_u8_u2_n152, u0_u8_u2_n153, u0_u8_u2_n154, u0_u8_u2_n155, u0_u8_u2_n156, u0_u8_u2_n157, u0_u8_u2_n158, 
       u0_u8_u2_n159, u0_u8_u2_n160, u0_u8_u2_n161, u0_u8_u2_n162, u0_u8_u2_n163, u0_u8_u2_n164, u0_u8_u2_n165, u0_u8_u2_n166, u0_u8_u2_n167, 
       u0_u8_u2_n168, u0_u8_u2_n169, u0_u8_u2_n170, u0_u8_u2_n171, u0_u8_u2_n172, u0_u8_u2_n173, u0_u8_u2_n174, u0_u8_u2_n175, u0_u8_u2_n176, 
       u0_u8_u2_n177, u0_u8_u2_n178, u0_u8_u2_n179, u0_u8_u2_n180, u0_u8_u2_n181, u0_u8_u2_n182, u0_u8_u2_n183, u0_u8_u2_n184, u0_u8_u2_n185, 
       u0_u8_u2_n186, u0_u8_u2_n187, u0_u8_u2_n188, u0_u8_u2_n95, u0_u8_u2_n96, u0_u8_u2_n97, u0_u8_u2_n98, u0_u8_u2_n99, u0_u8_u3_n100, 
       u0_u8_u3_n101, u0_u8_u3_n102, u0_u8_u3_n103, u0_u8_u3_n104, u0_u8_u3_n105, u0_u8_u3_n106, u0_u8_u3_n107, u0_u8_u3_n108, u0_u8_u3_n109, 
       u0_u8_u3_n110, u0_u8_u3_n111, u0_u8_u3_n112, u0_u8_u3_n113, u0_u8_u3_n114, u0_u8_u3_n115, u0_u8_u3_n116, u0_u8_u3_n117, u0_u8_u3_n118, 
       u0_u8_u3_n119, u0_u8_u3_n120, u0_u8_u3_n121, u0_u8_u3_n122, u0_u8_u3_n123, u0_u8_u3_n124, u0_u8_u3_n125, u0_u8_u3_n126, u0_u8_u3_n127, 
       u0_u8_u3_n128, u0_u8_u3_n129, u0_u8_u3_n130, u0_u8_u3_n131, u0_u8_u3_n132, u0_u8_u3_n133, u0_u8_u3_n134, u0_u8_u3_n135, u0_u8_u3_n136, 
       u0_u8_u3_n137, u0_u8_u3_n138, u0_u8_u3_n139, u0_u8_u3_n140, u0_u8_u3_n141, u0_u8_u3_n142, u0_u8_u3_n143, u0_u8_u3_n144, u0_u8_u3_n145, 
       u0_u8_u3_n146, u0_u8_u3_n147, u0_u8_u3_n148, u0_u8_u3_n149, u0_u8_u3_n150, u0_u8_u3_n151, u0_u8_u3_n152, u0_u8_u3_n153, u0_u8_u3_n154, 
       u0_u8_u3_n155, u0_u8_u3_n156, u0_u8_u3_n157, u0_u8_u3_n158, u0_u8_u3_n159, u0_u8_u3_n160, u0_u8_u3_n161, u0_u8_u3_n162, u0_u8_u3_n163, 
       u0_u8_u3_n164, u0_u8_u3_n165, u0_u8_u3_n166, u0_u8_u3_n167, u0_u8_u3_n168, u0_u8_u3_n169, u0_u8_u3_n170, u0_u8_u3_n171, u0_u8_u3_n172, 
       u0_u8_u3_n173, u0_u8_u3_n174, u0_u8_u3_n175, u0_u8_u3_n176, u0_u8_u3_n177, u0_u8_u3_n178, u0_u8_u3_n179, u0_u8_u3_n180, u0_u8_u3_n181, 
       u0_u8_u3_n182, u0_u8_u3_n183, u0_u8_u3_n184, u0_u8_u3_n185, u0_u8_u3_n186, u0_u8_u3_n94, u0_u8_u3_n95, u0_u8_u3_n96, u0_u8_u3_n97, 
       u0_u8_u3_n98, u0_u8_u3_n99, u0_u8_u4_n100, u0_u8_u4_n101, u0_u8_u4_n102, u0_u8_u4_n103, u0_u8_u4_n104, u0_u8_u4_n105, u0_u8_u4_n106, 
       u0_u8_u4_n107, u0_u8_u4_n108, u0_u8_u4_n109, u0_u8_u4_n110, u0_u8_u4_n111, u0_u8_u4_n112, u0_u8_u4_n113, u0_u8_u4_n114, u0_u8_u4_n115, 
       u0_u8_u4_n116, u0_u8_u4_n117, u0_u8_u4_n118, u0_u8_u4_n119, u0_u8_u4_n120, u0_u8_u4_n121, u0_u8_u4_n122, u0_u8_u4_n123, u0_u8_u4_n124, 
       u0_u8_u4_n125, u0_u8_u4_n126, u0_u8_u4_n127, u0_u8_u4_n128, u0_u8_u4_n129, u0_u8_u4_n130, u0_u8_u4_n131, u0_u8_u4_n132, u0_u8_u4_n133, 
       u0_u8_u4_n134, u0_u8_u4_n135, u0_u8_u4_n136, u0_u8_u4_n137, u0_u8_u4_n138, u0_u8_u4_n139, u0_u8_u4_n140, u0_u8_u4_n141, u0_u8_u4_n142, 
       u0_u8_u4_n143, u0_u8_u4_n144, u0_u8_u4_n145, u0_u8_u4_n146, u0_u8_u4_n147, u0_u8_u4_n148, u0_u8_u4_n149, u0_u8_u4_n150, u0_u8_u4_n151, 
       u0_u8_u4_n152, u0_u8_u4_n153, u0_u8_u4_n154, u0_u8_u4_n155, u0_u8_u4_n156, u0_u8_u4_n157, u0_u8_u4_n158, u0_u8_u4_n159, u0_u8_u4_n160, 
       u0_u8_u4_n161, u0_u8_u4_n162, u0_u8_u4_n163, u0_u8_u4_n164, u0_u8_u4_n165, u0_u8_u4_n166, u0_u8_u4_n167, u0_u8_u4_n168, u0_u8_u4_n169, 
       u0_u8_u4_n170, u0_u8_u4_n171, u0_u8_u4_n172, u0_u8_u4_n173, u0_u8_u4_n174, u0_u8_u4_n175, u0_u8_u4_n176, u0_u8_u4_n177, u0_u8_u4_n178, 
       u0_u8_u4_n179, u0_u8_u4_n180, u0_u8_u4_n181, u0_u8_u4_n182, u0_u8_u4_n183, u0_u8_u4_n184, u0_u8_u4_n185, u0_u8_u4_n186, u0_u8_u4_n94, 
       u0_u8_u4_n95, u0_u8_u4_n96, u0_u8_u4_n97, u0_u8_u4_n98, u0_u8_u4_n99, u0_u8_u7_n100, u0_u8_u7_n101, u0_u8_u7_n102, u0_u8_u7_n103, 
       u0_u8_u7_n104, u0_u8_u7_n105, u0_u8_u7_n106, u0_u8_u7_n107, u0_u8_u7_n108, u0_u8_u7_n109, u0_u8_u7_n110, u0_u8_u7_n111, u0_u8_u7_n112, 
       u0_u8_u7_n113, u0_u8_u7_n114, u0_u8_u7_n115, u0_u8_u7_n116, u0_u8_u7_n117, u0_u8_u7_n118, u0_u8_u7_n119, u0_u8_u7_n120, u0_u8_u7_n121, 
       u0_u8_u7_n122, u0_u8_u7_n123, u0_u8_u7_n124, u0_u8_u7_n125, u0_u8_u7_n126, u0_u8_u7_n127, u0_u8_u7_n128, u0_u8_u7_n129, u0_u8_u7_n130, 
       u0_u8_u7_n131, u0_u8_u7_n132, u0_u8_u7_n133, u0_u8_u7_n134, u0_u8_u7_n135, u0_u8_u7_n136, u0_u8_u7_n137, u0_u8_u7_n138, u0_u8_u7_n139, 
       u0_u8_u7_n140, u0_u8_u7_n141, u0_u8_u7_n142, u0_u8_u7_n143, u0_u8_u7_n144, u0_u8_u7_n145, u0_u8_u7_n146, u0_u8_u7_n147, u0_u8_u7_n148, 
       u0_u8_u7_n149, u0_u8_u7_n150, u0_u8_u7_n151, u0_u8_u7_n152, u0_u8_u7_n153, u0_u8_u7_n154, u0_u8_u7_n155, u0_u8_u7_n156, u0_u8_u7_n157, 
       u0_u8_u7_n158, u0_u8_u7_n159, u0_u8_u7_n160, u0_u8_u7_n161, u0_u8_u7_n162, u0_u8_u7_n163, u0_u8_u7_n164, u0_u8_u7_n165, u0_u8_u7_n166, 
       u0_u8_u7_n167, u0_u8_u7_n168, u0_u8_u7_n169, u0_u8_u7_n170, u0_u8_u7_n171, u0_u8_u7_n172, u0_u8_u7_n173, u0_u8_u7_n174, u0_u8_u7_n175, 
       u0_u8_u7_n176, u0_u8_u7_n177, u0_u8_u7_n178, u0_u8_u7_n179, u0_u8_u7_n180, u0_u8_u7_n91, u0_u8_u7_n92, u0_u8_u7_n93, u0_u8_u7_n94, 
       u0_u8_u7_n95, u0_u8_u7_n96, u0_u8_u7_n97, u0_u8_u7_n98, u0_u8_u7_n99, u0_u9_X_10, u0_u9_X_11, u0_u9_X_12, u0_u9_X_13, 
       u0_u9_X_14, u0_u9_X_15, u0_u9_X_16, u0_u9_X_17, u0_u9_X_18, u0_u9_X_19, u0_u9_X_20, u0_u9_X_21, u0_u9_X_22, 
       u0_u9_X_23, u0_u9_X_24, u0_u9_X_7, u0_u9_X_8, u0_u9_X_9, u0_u9_u1_n100, u0_u9_u1_n101, u0_u9_u1_n102, u0_u9_u1_n103, 
       u0_u9_u1_n104, u0_u9_u1_n105, u0_u9_u1_n106, u0_u9_u1_n107, u0_u9_u1_n108, u0_u9_u1_n109, u0_u9_u1_n110, u0_u9_u1_n111, u0_u9_u1_n112, 
       u0_u9_u1_n113, u0_u9_u1_n114, u0_u9_u1_n115, u0_u9_u1_n116, u0_u9_u1_n117, u0_u9_u1_n118, u0_u9_u1_n119, u0_u9_u1_n120, u0_u9_u1_n121, 
       u0_u9_u1_n122, u0_u9_u1_n123, u0_u9_u1_n124, u0_u9_u1_n125, u0_u9_u1_n126, u0_u9_u1_n127, u0_u9_u1_n128, u0_u9_u1_n129, u0_u9_u1_n130, 
       u0_u9_u1_n131, u0_u9_u1_n132, u0_u9_u1_n133, u0_u9_u1_n134, u0_u9_u1_n135, u0_u9_u1_n136, u0_u9_u1_n137, u0_u9_u1_n138, u0_u9_u1_n139, 
       u0_u9_u1_n140, u0_u9_u1_n141, u0_u9_u1_n142, u0_u9_u1_n143, u0_u9_u1_n144, u0_u9_u1_n145, u0_u9_u1_n146, u0_u9_u1_n147, u0_u9_u1_n148, 
       u0_u9_u1_n149, u0_u9_u1_n150, u0_u9_u1_n151, u0_u9_u1_n152, u0_u9_u1_n153, u0_u9_u1_n154, u0_u9_u1_n155, u0_u9_u1_n156, u0_u9_u1_n157, 
       u0_u9_u1_n158, u0_u9_u1_n159, u0_u9_u1_n160, u0_u9_u1_n161, u0_u9_u1_n162, u0_u9_u1_n163, u0_u9_u1_n164, u0_u9_u1_n165, u0_u9_u1_n166, 
       u0_u9_u1_n167, u0_u9_u1_n168, u0_u9_u1_n169, u0_u9_u1_n170, u0_u9_u1_n171, u0_u9_u1_n172, u0_u9_u1_n173, u0_u9_u1_n174, u0_u9_u1_n175, 
       u0_u9_u1_n176, u0_u9_u1_n177, u0_u9_u1_n178, u0_u9_u1_n179, u0_u9_u1_n180, u0_u9_u1_n181, u0_u9_u1_n182, u0_u9_u1_n183, u0_u9_u1_n184, 
       u0_u9_u1_n185, u0_u9_u1_n186, u0_u9_u1_n187, u0_u9_u1_n188, u0_u9_u1_n95, u0_u9_u1_n96, u0_u9_u1_n97, u0_u9_u1_n98, u0_u9_u1_n99, 
       u0_u9_u2_n100, u0_u9_u2_n101, u0_u9_u2_n102, u0_u9_u2_n103, u0_u9_u2_n104, u0_u9_u2_n105, u0_u9_u2_n106, u0_u9_u2_n107, u0_u9_u2_n108, 
       u0_u9_u2_n109, u0_u9_u2_n110, u0_u9_u2_n111, u0_u9_u2_n112, u0_u9_u2_n113, u0_u9_u2_n114, u0_u9_u2_n115, u0_u9_u2_n116, u0_u9_u2_n117, 
       u0_u9_u2_n118, u0_u9_u2_n119, u0_u9_u2_n120, u0_u9_u2_n121, u0_u9_u2_n122, u0_u9_u2_n123, u0_u9_u2_n124, u0_u9_u2_n125, u0_u9_u2_n126, 
       u0_u9_u2_n127, u0_u9_u2_n128, u0_u9_u2_n129, u0_u9_u2_n130, u0_u9_u2_n131, u0_u9_u2_n132, u0_u9_u2_n133, u0_u9_u2_n134, u0_u9_u2_n135, 
       u0_u9_u2_n136, u0_u9_u2_n137, u0_u9_u2_n138, u0_u9_u2_n139, u0_u9_u2_n140, u0_u9_u2_n141, u0_u9_u2_n142, u0_u9_u2_n143, u0_u9_u2_n144, 
       u0_u9_u2_n145, u0_u9_u2_n146, u0_u9_u2_n147, u0_u9_u2_n148, u0_u9_u2_n149, u0_u9_u2_n150, u0_u9_u2_n151, u0_u9_u2_n152, u0_u9_u2_n153, 
       u0_u9_u2_n154, u0_u9_u2_n155, u0_u9_u2_n156, u0_u9_u2_n157, u0_u9_u2_n158, u0_u9_u2_n159, u0_u9_u2_n160, u0_u9_u2_n161, u0_u9_u2_n162, 
       u0_u9_u2_n163, u0_u9_u2_n164, u0_u9_u2_n165, u0_u9_u2_n166, u0_u9_u2_n167, u0_u9_u2_n168, u0_u9_u2_n169, u0_u9_u2_n170, u0_u9_u2_n171, 
       u0_u9_u2_n172, u0_u9_u2_n173, u0_u9_u2_n174, u0_u9_u2_n175, u0_u9_u2_n176, u0_u9_u2_n177, u0_u9_u2_n178, u0_u9_u2_n179, u0_u9_u2_n180, 
       u0_u9_u2_n181, u0_u9_u2_n182, u0_u9_u2_n183, u0_u9_u2_n184, u0_u9_u2_n185, u0_u9_u2_n186, u0_u9_u2_n187, u0_u9_u2_n188, u0_u9_u2_n95, 
       u0_u9_u2_n96, u0_u9_u2_n97, u0_u9_u2_n98, u0_u9_u2_n99, u0_u9_u3_n100, u0_u9_u3_n101, u0_u9_u3_n102, u0_u9_u3_n103, u0_u9_u3_n104, 
       u0_u9_u3_n105, u0_u9_u3_n106, u0_u9_u3_n107, u0_u9_u3_n108, u0_u9_u3_n109, u0_u9_u3_n110, u0_u9_u3_n111, u0_u9_u3_n112, u0_u9_u3_n113, 
       u0_u9_u3_n114, u0_u9_u3_n115, u0_u9_u3_n116, u0_u9_u3_n117, u0_u9_u3_n118, u0_u9_u3_n119, u0_u9_u3_n120, u0_u9_u3_n121, u0_u9_u3_n122, 
       u0_u9_u3_n123, u0_u9_u3_n124, u0_u9_u3_n125, u0_u9_u3_n126, u0_u9_u3_n127, u0_u9_u3_n128, u0_u9_u3_n129, u0_u9_u3_n130, u0_u9_u3_n131, 
       u0_u9_u3_n132, u0_u9_u3_n133, u0_u9_u3_n134, u0_u9_u3_n135, u0_u9_u3_n136, u0_u9_u3_n137, u0_u9_u3_n138, u0_u9_u3_n139, u0_u9_u3_n140, 
       u0_u9_u3_n141, u0_u9_u3_n142, u0_u9_u3_n143, u0_u9_u3_n144, u0_u9_u3_n145, u0_u9_u3_n146, u0_u9_u3_n147, u0_u9_u3_n148, u0_u9_u3_n149, 
       u0_u9_u3_n150, u0_u9_u3_n151, u0_u9_u3_n152, u0_u9_u3_n153, u0_u9_u3_n154, u0_u9_u3_n155, u0_u9_u3_n156, u0_u9_u3_n157, u0_u9_u3_n158, 
       u0_u9_u3_n159, u0_u9_u3_n160, u0_u9_u3_n161, u0_u9_u3_n162, u0_u9_u3_n163, u0_u9_u3_n164, u0_u9_u3_n165, u0_u9_u3_n166, u0_u9_u3_n167, 
       u0_u9_u3_n168, u0_u9_u3_n169, u0_u9_u3_n170, u0_u9_u3_n171, u0_u9_u3_n172, u0_u9_u3_n173, u0_u9_u3_n174, u0_u9_u3_n175, u0_u9_u3_n176, 
       u0_u9_u3_n177, u0_u9_u3_n178, u0_u9_u3_n179, u0_u9_u3_n180, u0_u9_u3_n181, u0_u9_u3_n182, u0_u9_u3_n183, u0_u9_u3_n184, u0_u9_u3_n185, 
       u0_u9_u3_n186, u0_u9_u3_n94, u0_u9_u3_n95, u0_u9_u3_n96, u0_u9_u3_n97, u0_u9_u3_n98, u0_u9_u3_n99, u0_uk_n1005, u0_uk_n1017, 
       u0_uk_n1018, u0_uk_n1022, u0_uk_n718, u0_uk_n721, u0_uk_n729, u0_uk_n730, u0_uk_n733, u0_uk_n734, u0_uk_n737, 
       u0_uk_n741, u0_uk_n742, u0_uk_n774, u0_uk_n776, u0_uk_n779, u0_uk_n791, u0_uk_n794, u0_uk_n795, u0_uk_n857, 
       u0_uk_n895, u0_uk_n896, u0_uk_n899, u0_uk_n900, u0_uk_n901, u0_uk_n912, u0_uk_n913, u0_uk_n922, u0_uk_n923, 
       u0_uk_n924, u0_uk_n925, u0_uk_n947, u0_uk_n993, u0_uk_n994, u0_uk_n995, u1_K11_30, u1_K11_31, u1_K11_34, 
       u1_K11_5, u1_K11_8, u1_K14_34, u1_K4_3, u1_K4_4, u1_K5_22, u1_K7_27, u1_K9_33, u1_out0_16, 
       u1_out0_24, u1_out0_30, u1_out0_6, u1_out10_11, u1_out10_13, u1_out10_14, u1_out10_17, u1_out10_18, u1_out10_19, 
       u1_out10_2, u1_out10_23, u1_out10_25, u1_out10_28, u1_out10_29, u1_out10_3, u1_out10_31, u1_out10_4, u1_out10_8, 
       u1_out10_9, u1_out11_11, u1_out11_19, u1_out11_29, u1_out11_4, u1_out12_12, u1_out12_22, u1_out12_32, u1_out12_7, 
       u1_out13_11, u1_out13_19, u1_out13_29, u1_out13_4, u1_out14_14, u1_out14_25, u1_out14_3, u1_out14_8, u1_out15_17, 
       u1_out15_23, u1_out15_31, u1_out15_9, u1_out2_11, u1_out2_16, u1_out2_19, u1_out2_24, u1_out2_29, u1_out2_30, 
       u1_out2_4, u1_out2_6, u1_out3_17, u1_out3_23, u1_out3_31, u1_out3_9, u1_out4_1, u1_out4_10, u1_out4_13, 
       u1_out4_17, u1_out4_18, u1_out4_2, u1_out4_20, u1_out4_23, u1_out4_26, u1_out4_28, u1_out4_31, u1_out4_9, 
       u1_out6_12, u1_out6_14, u1_out6_17, u1_out6_22, u1_out6_23, u1_out6_25, u1_out6_3, u1_out6_31, u1_out6_32, 
       u1_out6_7, u1_out6_8, u1_out6_9, u1_out7_1, u1_out7_10, u1_out7_20, u1_out7_26, u1_out8_11, u1_out8_19, 
       u1_out8_29, u1_out8_4, u1_out9_14, u1_out9_25, u1_out9_3, u1_out9_8, u1_u0_X_15, u1_u0_X_16, u1_u0_u2_n100, 
       u1_u0_u2_n101, u1_u0_u2_n102, u1_u0_u2_n103, u1_u0_u2_n104, u1_u0_u2_n105, u1_u0_u2_n106, u1_u0_u2_n107, u1_u0_u2_n108, u1_u0_u2_n109, 
       u1_u0_u2_n110, u1_u0_u2_n111, u1_u0_u2_n112, u1_u0_u2_n113, u1_u0_u2_n114, u1_u0_u2_n115, u1_u0_u2_n116, u1_u0_u2_n117, u1_u0_u2_n118, 
       u1_u0_u2_n119, u1_u0_u2_n120, u1_u0_u2_n121, u1_u0_u2_n122, u1_u0_u2_n123, u1_u0_u2_n124, u1_u0_u2_n125, u1_u0_u2_n126, u1_u0_u2_n127, 
       u1_u0_u2_n128, u1_u0_u2_n129, u1_u0_u2_n130, u1_u0_u2_n131, u1_u0_u2_n132, u1_u0_u2_n133, u1_u0_u2_n134, u1_u0_u2_n135, u1_u0_u2_n136, 
       u1_u0_u2_n137, u1_u0_u2_n138, u1_u0_u2_n139, u1_u0_u2_n140, u1_u0_u2_n141, u1_u0_u2_n142, u1_u0_u2_n143, u1_u0_u2_n144, u1_u0_u2_n145, 
       u1_u0_u2_n146, u1_u0_u2_n147, u1_u0_u2_n148, u1_u0_u2_n149, u1_u0_u2_n150, u1_u0_u2_n151, u1_u0_u2_n152, u1_u0_u2_n153, u1_u0_u2_n154, 
       u1_u0_u2_n155, u1_u0_u2_n156, u1_u0_u2_n157, u1_u0_u2_n158, u1_u0_u2_n159, u1_u0_u2_n160, u1_u0_u2_n161, u1_u0_u2_n162, u1_u0_u2_n163, 
       u1_u0_u2_n164, u1_u0_u2_n165, u1_u0_u2_n166, u1_u0_u2_n167, u1_u0_u2_n168, u1_u0_u2_n169, u1_u0_u2_n170, u1_u0_u2_n171, u1_u0_u2_n172, 
       u1_u0_u2_n173, u1_u0_u2_n174, u1_u0_u2_n175, u1_u0_u2_n176, u1_u0_u2_n177, u1_u0_u2_n178, u1_u0_u2_n179, u1_u0_u2_n180, u1_u0_u2_n181, 
       u1_u0_u2_n182, u1_u0_u2_n183, u1_u0_u2_n184, u1_u0_u2_n185, u1_u0_u2_n186, u1_u0_u2_n187, u1_u0_u2_n188, u1_u0_u2_n95, u1_u0_u2_n96, 
       u1_u0_u2_n97, u1_u0_u2_n98, u1_u0_u2_n99, u1_u10_X_10, u1_u10_X_27, u1_u10_X_28, u1_u10_X_29, u1_u10_X_3, u1_u10_X_30, 
       u1_u10_X_31, u1_u10_X_32, u1_u10_X_33, u1_u10_X_34, u1_u10_X_4, u1_u10_X_5, u1_u10_X_6, u1_u10_X_7, u1_u10_X_8, 
       u1_u10_X_9, u1_u10_u0_n100, u1_u10_u0_n101, u1_u10_u0_n102, u1_u10_u0_n103, u1_u10_u0_n104, u1_u10_u0_n105, u1_u10_u0_n106, u1_u10_u0_n107, 
       u1_u10_u0_n108, u1_u10_u0_n109, u1_u10_u0_n110, u1_u10_u0_n111, u1_u10_u0_n112, u1_u10_u0_n113, u1_u10_u0_n114, u1_u10_u0_n115, u1_u10_u0_n116, 
       u1_u10_u0_n117, u1_u10_u0_n118, u1_u10_u0_n119, u1_u10_u0_n120, u1_u10_u0_n121, u1_u10_u0_n122, u1_u10_u0_n123, u1_u10_u0_n124, u1_u10_u0_n125, 
       u1_u10_u0_n126, u1_u10_u0_n127, u1_u10_u0_n128, u1_u10_u0_n129, u1_u10_u0_n130, u1_u10_u0_n131, u1_u10_u0_n132, u1_u10_u0_n133, u1_u10_u0_n134, 
       u1_u10_u0_n135, u1_u10_u0_n136, u1_u10_u0_n137, u1_u10_u0_n138, u1_u10_u0_n139, u1_u10_u0_n140, u1_u10_u0_n141, u1_u10_u0_n142, u1_u10_u0_n143, 
       u1_u10_u0_n144, u1_u10_u0_n145, u1_u10_u0_n146, u1_u10_u0_n147, u1_u10_u0_n148, u1_u10_u0_n149, u1_u10_u0_n150, u1_u10_u0_n151, u1_u10_u0_n152, 
       u1_u10_u0_n153, u1_u10_u0_n154, u1_u10_u0_n155, u1_u10_u0_n156, u1_u10_u0_n157, u1_u10_u0_n158, u1_u10_u0_n159, u1_u10_u0_n160, u1_u10_u0_n161, 
       u1_u10_u0_n162, u1_u10_u0_n163, u1_u10_u0_n164, u1_u10_u0_n165, u1_u10_u0_n166, u1_u10_u0_n167, u1_u10_u0_n168, u1_u10_u0_n169, u1_u10_u0_n170, 
       u1_u10_u0_n171, u1_u10_u0_n172, u1_u10_u0_n173, u1_u10_u0_n174, u1_u10_u0_n88, u1_u10_u0_n89, u1_u10_u0_n90, u1_u10_u0_n91, u1_u10_u0_n92, 
       u1_u10_u0_n93, u1_u10_u0_n94, u1_u10_u0_n95, u1_u10_u0_n96, u1_u10_u0_n97, u1_u10_u0_n98, u1_u10_u0_n99, u1_u10_u1_n100, u1_u10_u1_n101, 
       u1_u10_u1_n102, u1_u10_u1_n103, u1_u10_u1_n104, u1_u10_u1_n105, u1_u10_u1_n106, u1_u10_u1_n107, u1_u10_u1_n108, u1_u10_u1_n109, u1_u10_u1_n110, 
       u1_u10_u1_n111, u1_u10_u1_n112, u1_u10_u1_n113, u1_u10_u1_n114, u1_u10_u1_n115, u1_u10_u1_n116, u1_u10_u1_n117, u1_u10_u1_n118, u1_u10_u1_n119, 
       u1_u10_u1_n120, u1_u10_u1_n121, u1_u10_u1_n122, u1_u10_u1_n123, u1_u10_u1_n124, u1_u10_u1_n125, u1_u10_u1_n126, u1_u10_u1_n127, u1_u10_u1_n128, 
       u1_u10_u1_n129, u1_u10_u1_n130, u1_u10_u1_n131, u1_u10_u1_n132, u1_u10_u1_n133, u1_u10_u1_n134, u1_u10_u1_n135, u1_u10_u1_n136, u1_u10_u1_n137, 
       u1_u10_u1_n138, u1_u10_u1_n139, u1_u10_u1_n140, u1_u10_u1_n141, u1_u10_u1_n142, u1_u10_u1_n143, u1_u10_u1_n144, u1_u10_u1_n145, u1_u10_u1_n146, 
       u1_u10_u1_n147, u1_u10_u1_n148, u1_u10_u1_n149, u1_u10_u1_n150, u1_u10_u1_n151, u1_u10_u1_n152, u1_u10_u1_n153, u1_u10_u1_n154, u1_u10_u1_n155, 
       u1_u10_u1_n156, u1_u10_u1_n157, u1_u10_u1_n158, u1_u10_u1_n159, u1_u10_u1_n160, u1_u10_u1_n161, u1_u10_u1_n162, u1_u10_u1_n163, u1_u10_u1_n164, 
       u1_u10_u1_n165, u1_u10_u1_n166, u1_u10_u1_n167, u1_u10_u1_n168, u1_u10_u1_n169, u1_u10_u1_n170, u1_u10_u1_n171, u1_u10_u1_n172, u1_u10_u1_n173, 
       u1_u10_u1_n174, u1_u10_u1_n175, u1_u10_u1_n176, u1_u10_u1_n177, u1_u10_u1_n178, u1_u10_u1_n179, u1_u10_u1_n180, u1_u10_u1_n181, u1_u10_u1_n182, 
       u1_u10_u1_n183, u1_u10_u1_n184, u1_u10_u1_n185, u1_u10_u1_n186, u1_u10_u1_n187, u1_u10_u1_n188, u1_u10_u1_n95, u1_u10_u1_n96, u1_u10_u1_n97, 
       u1_u10_u1_n98, u1_u10_u1_n99, u1_u10_u4_n100, u1_u10_u4_n101, u1_u10_u4_n102, u1_u10_u4_n103, u1_u10_u4_n104, u1_u10_u4_n105, u1_u10_u4_n106, 
       u1_u10_u4_n107, u1_u10_u4_n108, u1_u10_u4_n109, u1_u10_u4_n110, u1_u10_u4_n111, u1_u10_u4_n112, u1_u10_u4_n113, u1_u10_u4_n114, u1_u10_u4_n115, 
       u1_u10_u4_n116, u1_u10_u4_n117, u1_u10_u4_n118, u1_u10_u4_n119, u1_u10_u4_n120, u1_u10_u4_n121, u1_u10_u4_n122, u1_u10_u4_n123, u1_u10_u4_n124, 
       u1_u10_u4_n125, u1_u10_u4_n126, u1_u10_u4_n127, u1_u10_u4_n128, u1_u10_u4_n129, u1_u10_u4_n130, u1_u10_u4_n131, u1_u10_u4_n132, u1_u10_u4_n133, 
       u1_u10_u4_n134, u1_u10_u4_n135, u1_u10_u4_n136, u1_u10_u4_n137, u1_u10_u4_n138, u1_u10_u4_n139, u1_u10_u4_n140, u1_u10_u4_n141, u1_u10_u4_n142, 
       u1_u10_u4_n143, u1_u10_u4_n144, u1_u10_u4_n145, u1_u10_u4_n146, u1_u10_u4_n147, u1_u10_u4_n148, u1_u10_u4_n149, u1_u10_u4_n150, u1_u10_u4_n151, 
       u1_u10_u4_n152, u1_u10_u4_n153, u1_u10_u4_n154, u1_u10_u4_n155, u1_u10_u4_n156, u1_u10_u4_n157, u1_u10_u4_n158, u1_u10_u4_n159, u1_u10_u4_n160, 
       u1_u10_u4_n161, u1_u10_u4_n162, u1_u10_u4_n163, u1_u10_u4_n164, u1_u10_u4_n165, u1_u10_u4_n166, u1_u10_u4_n167, u1_u10_u4_n168, u1_u10_u4_n169, 
       u1_u10_u4_n170, u1_u10_u4_n171, u1_u10_u4_n172, u1_u10_u4_n173, u1_u10_u4_n174, u1_u10_u4_n175, u1_u10_u4_n176, u1_u10_u4_n177, u1_u10_u4_n178, 
       u1_u10_u4_n179, u1_u10_u4_n180, u1_u10_u4_n181, u1_u10_u4_n182, u1_u10_u4_n183, u1_u10_u4_n184, u1_u10_u4_n185, u1_u10_u4_n186, u1_u10_u4_n94, 
       u1_u10_u4_n95, u1_u10_u4_n96, u1_u10_u4_n97, u1_u10_u4_n98, u1_u10_u4_n99, u1_u10_u5_n100, u1_u10_u5_n101, u1_u10_u5_n102, u1_u10_u5_n103, 
       u1_u10_u5_n104, u1_u10_u5_n105, u1_u10_u5_n106, u1_u10_u5_n107, u1_u10_u5_n108, u1_u10_u5_n109, u1_u10_u5_n110, u1_u10_u5_n111, u1_u10_u5_n112, 
       u1_u10_u5_n113, u1_u10_u5_n114, u1_u10_u5_n115, u1_u10_u5_n116, u1_u10_u5_n117, u1_u10_u5_n118, u1_u10_u5_n119, u1_u10_u5_n120, u1_u10_u5_n121, 
       u1_u10_u5_n122, u1_u10_u5_n123, u1_u10_u5_n124, u1_u10_u5_n125, u1_u10_u5_n126, u1_u10_u5_n127, u1_u10_u5_n128, u1_u10_u5_n129, u1_u10_u5_n130, 
       u1_u10_u5_n131, u1_u10_u5_n132, u1_u10_u5_n133, u1_u10_u5_n134, u1_u10_u5_n135, u1_u10_u5_n136, u1_u10_u5_n137, u1_u10_u5_n138, u1_u10_u5_n139, 
       u1_u10_u5_n140, u1_u10_u5_n141, u1_u10_u5_n142, u1_u10_u5_n143, u1_u10_u5_n144, u1_u10_u5_n145, u1_u10_u5_n146, u1_u10_u5_n147, u1_u10_u5_n148, 
       u1_u10_u5_n149, u1_u10_u5_n150, u1_u10_u5_n151, u1_u10_u5_n152, u1_u10_u5_n153, u1_u10_u5_n154, u1_u10_u5_n155, u1_u10_u5_n156, u1_u10_u5_n157, 
       u1_u10_u5_n158, u1_u10_u5_n159, u1_u10_u5_n160, u1_u10_u5_n161, u1_u10_u5_n162, u1_u10_u5_n163, u1_u10_u5_n164, u1_u10_u5_n165, u1_u10_u5_n166, 
       u1_u10_u5_n167, u1_u10_u5_n168, u1_u10_u5_n169, u1_u10_u5_n170, u1_u10_u5_n171, u1_u10_u5_n172, u1_u10_u5_n173, u1_u10_u5_n174, u1_u10_u5_n175, 
       u1_u10_u5_n176, u1_u10_u5_n177, u1_u10_u5_n178, u1_u10_u5_n179, u1_u10_u5_n180, u1_u10_u5_n181, u1_u10_u5_n182, u1_u10_u5_n183, u1_u10_u5_n184, 
       u1_u10_u5_n185, u1_u10_u5_n186, u1_u10_u5_n187, u1_u10_u5_n188, u1_u10_u5_n189, u1_u10_u5_n190, u1_u10_u5_n191, u1_u10_u5_n192, u1_u10_u5_n193, 
       u1_u10_u5_n194, u1_u10_u5_n195, u1_u10_u5_n196, u1_u10_u5_n99, u1_u11_X_33, u1_u11_X_34, u1_u11_u5_n100, u1_u11_u5_n101, u1_u11_u5_n102, 
       u1_u11_u5_n103, u1_u11_u5_n104, u1_u11_u5_n105, u1_u11_u5_n106, u1_u11_u5_n107, u1_u11_u5_n108, u1_u11_u5_n109, u1_u11_u5_n110, u1_u11_u5_n111, 
       u1_u11_u5_n112, u1_u11_u5_n113, u1_u11_u5_n114, u1_u11_u5_n115, u1_u11_u5_n116, u1_u11_u5_n117, u1_u11_u5_n118, u1_u11_u5_n119, u1_u11_u5_n120, 
       u1_u11_u5_n121, u1_u11_u5_n122, u1_u11_u5_n123, u1_u11_u5_n124, u1_u11_u5_n125, u1_u11_u5_n126, u1_u11_u5_n127, u1_u11_u5_n128, u1_u11_u5_n129, 
       u1_u11_u5_n130, u1_u11_u5_n131, u1_u11_u5_n132, u1_u11_u5_n133, u1_u11_u5_n134, u1_u11_u5_n135, u1_u11_u5_n136, u1_u11_u5_n137, u1_u11_u5_n138, 
       u1_u11_u5_n139, u1_u11_u5_n140, u1_u11_u5_n141, u1_u11_u5_n142, u1_u11_u5_n143, u1_u11_u5_n144, u1_u11_u5_n145, u1_u11_u5_n146, u1_u11_u5_n147, 
       u1_u11_u5_n148, u1_u11_u5_n149, u1_u11_u5_n150, u1_u11_u5_n151, u1_u11_u5_n152, u1_u11_u5_n153, u1_u11_u5_n154, u1_u11_u5_n155, u1_u11_u5_n156, 
       u1_u11_u5_n157, u1_u11_u5_n158, u1_u11_u5_n159, u1_u11_u5_n160, u1_u11_u5_n161, u1_u11_u5_n162, u1_u11_u5_n163, u1_u11_u5_n164, u1_u11_u5_n165, 
       u1_u11_u5_n166, u1_u11_u5_n167, u1_u11_u5_n168, u1_u11_u5_n169, u1_u11_u5_n170, u1_u11_u5_n171, u1_u11_u5_n172, u1_u11_u5_n173, u1_u11_u5_n174, 
       u1_u11_u5_n175, u1_u11_u5_n176, u1_u11_u5_n177, u1_u11_u5_n178, u1_u11_u5_n179, u1_u11_u5_n180, u1_u11_u5_n181, u1_u11_u5_n182, u1_u11_u5_n183, 
       u1_u11_u5_n184, u1_u11_u5_n185, u1_u11_u5_n186, u1_u11_u5_n187, u1_u11_u5_n188, u1_u11_u5_n189, u1_u11_u5_n190, u1_u11_u5_n191, u1_u11_u5_n192, 
       u1_u11_u5_n193, u1_u11_u5_n194, u1_u11_u5_n195, u1_u11_u5_n196, u1_u11_u5_n99, u1_u12_X_39, u1_u12_X_40, u1_u12_u6_n100, u1_u12_u6_n101, 
       u1_u12_u6_n102, u1_u12_u6_n103, u1_u12_u6_n104, u1_u12_u6_n105, u1_u12_u6_n106, u1_u12_u6_n107, u1_u12_u6_n108, u1_u12_u6_n109, u1_u12_u6_n110, 
       u1_u12_u6_n111, u1_u12_u6_n112, u1_u12_u6_n113, u1_u12_u6_n114, u1_u12_u6_n115, u1_u12_u6_n116, u1_u12_u6_n117, u1_u12_u6_n118, u1_u12_u6_n119, 
       u1_u12_u6_n120, u1_u12_u6_n121, u1_u12_u6_n122, u1_u12_u6_n123, u1_u12_u6_n124, u1_u12_u6_n125, u1_u12_u6_n126, u1_u12_u6_n127, u1_u12_u6_n128, 
       u1_u12_u6_n129, u1_u12_u6_n130, u1_u12_u6_n131, u1_u12_u6_n132, u1_u12_u6_n133, u1_u12_u6_n134, u1_u12_u6_n135, u1_u12_u6_n136, u1_u12_u6_n137, 
       u1_u12_u6_n138, u1_u12_u6_n139, u1_u12_u6_n140, u1_u12_u6_n141, u1_u12_u6_n142, u1_u12_u6_n143, u1_u12_u6_n144, u1_u12_u6_n145, u1_u12_u6_n146, 
       u1_u12_u6_n147, u1_u12_u6_n148, u1_u12_u6_n149, u1_u12_u6_n150, u1_u12_u6_n151, u1_u12_u6_n152, u1_u12_u6_n153, u1_u12_u6_n154, u1_u12_u6_n155, 
       u1_u12_u6_n156, u1_u12_u6_n157, u1_u12_u6_n158, u1_u12_u6_n159, u1_u12_u6_n160, u1_u12_u6_n161, u1_u12_u6_n162, u1_u12_u6_n163, u1_u12_u6_n164, 
       u1_u12_u6_n165, u1_u12_u6_n166, u1_u12_u6_n167, u1_u12_u6_n168, u1_u12_u6_n169, u1_u12_u6_n170, u1_u12_u6_n171, u1_u12_u6_n172, u1_u12_u6_n173, 
       u1_u12_u6_n174, u1_u12_u6_n88, u1_u12_u6_n89, u1_u12_u6_n90, u1_u12_u6_n91, u1_u12_u6_n92, u1_u12_u6_n93, u1_u12_u6_n94, u1_u12_u6_n95, 
       u1_u12_u6_n96, u1_u12_u6_n97, u1_u12_u6_n98, u1_u12_u6_n99, u1_u13_X_33, u1_u13_X_34, u1_u13_u5_n100, u1_u13_u5_n101, u1_u13_u5_n102, 
       u1_u13_u5_n103, u1_u13_u5_n104, u1_u13_u5_n105, u1_u13_u5_n106, u1_u13_u5_n107, u1_u13_u5_n108, u1_u13_u5_n109, u1_u13_u5_n110, u1_u13_u5_n111, 
       u1_u13_u5_n112, u1_u13_u5_n113, u1_u13_u5_n114, u1_u13_u5_n115, u1_u13_u5_n116, u1_u13_u5_n117, u1_u13_u5_n118, u1_u13_u5_n119, u1_u13_u5_n120, 
       u1_u13_u5_n121, u1_u13_u5_n122, u1_u13_u5_n123, u1_u13_u5_n124, u1_u13_u5_n125, u1_u13_u5_n126, u1_u13_u5_n127, u1_u13_u5_n128, u1_u13_u5_n129, 
       u1_u13_u5_n130, u1_u13_u5_n131, u1_u13_u5_n132, u1_u13_u5_n133, u1_u13_u5_n134, u1_u13_u5_n135, u1_u13_u5_n136, u1_u13_u5_n137, u1_u13_u5_n138, 
       u1_u13_u5_n139, u1_u13_u5_n140, u1_u13_u5_n141, u1_u13_u5_n142, u1_u13_u5_n143, u1_u13_u5_n144, u1_u13_u5_n145, u1_u13_u5_n146, u1_u13_u5_n147, 
       u1_u13_u5_n148, u1_u13_u5_n149, u1_u13_u5_n150, u1_u13_u5_n151, u1_u13_u5_n152, u1_u13_u5_n153, u1_u13_u5_n154, u1_u13_u5_n155, u1_u13_u5_n156, 
       u1_u13_u5_n157, u1_u13_u5_n158, u1_u13_u5_n159, u1_u13_u5_n160, u1_u13_u5_n161, u1_u13_u5_n162, u1_u13_u5_n163, u1_u13_u5_n164, u1_u13_u5_n165, 
       u1_u13_u5_n166, u1_u13_u5_n167, u1_u13_u5_n168, u1_u13_u5_n169, u1_u13_u5_n170, u1_u13_u5_n171, u1_u13_u5_n172, u1_u13_u5_n173, u1_u13_u5_n174, 
       u1_u13_u5_n175, u1_u13_u5_n176, u1_u13_u5_n177, u1_u13_u5_n178, u1_u13_u5_n179, u1_u13_u5_n180, u1_u13_u5_n181, u1_u13_u5_n182, u1_u13_u5_n183, 
       u1_u13_u5_n184, u1_u13_u5_n185, u1_u13_u5_n186, u1_u13_u5_n187, u1_u13_u5_n188, u1_u13_u5_n189, u1_u13_u5_n190, u1_u13_u5_n191, u1_u13_u5_n192, 
       u1_u13_u5_n193, u1_u13_u5_n194, u1_u13_u5_n195, u1_u13_u5_n196, u1_u13_u5_n99, u1_u14_X_27, u1_u14_X_28, u1_u14_u4_n100, u1_u14_u4_n101, 
       u1_u14_u4_n102, u1_u14_u4_n103, u1_u14_u4_n104, u1_u14_u4_n105, u1_u14_u4_n106, u1_u14_u4_n107, u1_u14_u4_n108, u1_u14_u4_n109, u1_u14_u4_n110, 
       u1_u14_u4_n111, u1_u14_u4_n112, u1_u14_u4_n113, u1_u14_u4_n114, u1_u14_u4_n115, u1_u14_u4_n116, u1_u14_u4_n117, u1_u14_u4_n118, u1_u14_u4_n119, 
       u1_u14_u4_n120, u1_u14_u4_n121, u1_u14_u4_n122, u1_u14_u4_n123, u1_u14_u4_n124, u1_u14_u4_n125, u1_u14_u4_n126, u1_u14_u4_n127, u1_u14_u4_n128, 
       u1_u14_u4_n129, u1_u14_u4_n130, u1_u14_u4_n131, u1_u14_u4_n132, u1_u14_u4_n133, u1_u14_u4_n134, u1_u14_u4_n135, u1_u14_u4_n136, u1_u14_u4_n137, 
       u1_u14_u4_n138, u1_u14_u4_n139, u1_u14_u4_n140, u1_u14_u4_n141, u1_u14_u4_n142, u1_u14_u4_n143, u1_u14_u4_n144, u1_u14_u4_n145, u1_u14_u4_n146, 
       u1_u14_u4_n147, u1_u14_u4_n148, u1_u14_u4_n149, u1_u14_u4_n150, u1_u14_u4_n151, u1_u14_u4_n152, u1_u14_u4_n153, u1_u14_u4_n154, u1_u14_u4_n155, 
       u1_u14_u4_n156, u1_u14_u4_n157, u1_u14_u4_n158, u1_u14_u4_n159, u1_u14_u4_n160, u1_u14_u4_n161, u1_u14_u4_n162, u1_u14_u4_n163, u1_u14_u4_n164, 
       u1_u14_u4_n165, u1_u14_u4_n166, u1_u14_u4_n167, u1_u14_u4_n168, u1_u14_u4_n169, u1_u14_u4_n170, u1_u14_u4_n171, u1_u14_u4_n172, u1_u14_u4_n173, 
       u1_u14_u4_n174, u1_u14_u4_n175, u1_u14_u4_n176, u1_u14_u4_n177, u1_u14_u4_n178, u1_u14_u4_n179, u1_u14_u4_n180, u1_u14_u4_n181, u1_u14_u4_n182, 
       u1_u14_u4_n183, u1_u14_u4_n184, u1_u14_u4_n185, u1_u14_u4_n186, u1_u14_u4_n94, u1_u14_u4_n95, u1_u14_u4_n96, u1_u14_u4_n97, u1_u14_u4_n98, 
       u1_u14_u4_n99, u1_u15_X_3, u1_u15_X_4, u1_u15_u0_n100, u1_u15_u0_n101, u1_u15_u0_n102, u1_u15_u0_n103, u1_u15_u0_n104, u1_u15_u0_n105, 
       u1_u15_u0_n106, u1_u15_u0_n107, u1_u15_u0_n108, u1_u15_u0_n109, u1_u15_u0_n110, u1_u15_u0_n111, u1_u15_u0_n112, u1_u15_u0_n113, u1_u15_u0_n114, 
       u1_u15_u0_n115, u1_u15_u0_n116, u1_u15_u0_n117, u1_u15_u0_n118, u1_u15_u0_n119, u1_u15_u0_n120, u1_u15_u0_n121, u1_u15_u0_n122, u1_u15_u0_n123, 
       u1_u15_u0_n124, u1_u15_u0_n125, u1_u15_u0_n126, u1_u15_u0_n127, u1_u15_u0_n128, u1_u15_u0_n129, u1_u15_u0_n130, u1_u15_u0_n131, u1_u15_u0_n132, 
       u1_u15_u0_n133, u1_u15_u0_n134, u1_u15_u0_n135, u1_u15_u0_n136, u1_u15_u0_n137, u1_u15_u0_n138, u1_u15_u0_n139, u1_u15_u0_n140, u1_u15_u0_n141, 
       u1_u15_u0_n142, u1_u15_u0_n143, u1_u15_u0_n144, u1_u15_u0_n145, u1_u15_u0_n146, u1_u15_u0_n147, u1_u15_u0_n148, u1_u15_u0_n149, u1_u15_u0_n150, 
       u1_u15_u0_n151, u1_u15_u0_n152, u1_u15_u0_n153, u1_u15_u0_n154, u1_u15_u0_n155, u1_u15_u0_n156, u1_u15_u0_n157, u1_u15_u0_n158, u1_u15_u0_n159, 
       u1_u15_u0_n160, u1_u15_u0_n161, u1_u15_u0_n162, u1_u15_u0_n163, u1_u15_u0_n164, u1_u15_u0_n165, u1_u15_u0_n166, u1_u15_u0_n167, u1_u15_u0_n168, 
       u1_u15_u0_n169, u1_u15_u0_n170, u1_u15_u0_n171, u1_u15_u0_n172, u1_u15_u0_n173, u1_u15_u0_n174, u1_u15_u0_n88, u1_u15_u0_n89, u1_u15_u0_n90, 
       u1_u15_u0_n91, u1_u15_u0_n92, u1_u15_u0_n93, u1_u15_u0_n94, u1_u15_u0_n95, u1_u15_u0_n96, u1_u15_u0_n97, u1_u15_u0_n98, u1_u15_u0_n99, 
       u1_u2_X_15, u1_u2_X_16, u1_u2_X_33, u1_u2_X_34, u1_u2_u2_n100, u1_u2_u2_n101, u1_u2_u2_n102, u1_u2_u2_n103, u1_u2_u2_n104, 
       u1_u2_u2_n105, u1_u2_u2_n106, u1_u2_u2_n107, u1_u2_u2_n108, u1_u2_u2_n109, u1_u2_u2_n110, u1_u2_u2_n111, u1_u2_u2_n112, u1_u2_u2_n113, 
       u1_u2_u2_n114, u1_u2_u2_n115, u1_u2_u2_n116, u1_u2_u2_n117, u1_u2_u2_n118, u1_u2_u2_n119, u1_u2_u2_n120, u1_u2_u2_n121, u1_u2_u2_n122, 
       u1_u2_u2_n123, u1_u2_u2_n124, u1_u2_u2_n125, u1_u2_u2_n126, u1_u2_u2_n127, u1_u2_u2_n128, u1_u2_u2_n129, u1_u2_u2_n130, u1_u2_u2_n131, 
       u1_u2_u2_n132, u1_u2_u2_n133, u1_u2_u2_n134, u1_u2_u2_n135, u1_u2_u2_n136, u1_u2_u2_n137, u1_u2_u2_n138, u1_u2_u2_n139, u1_u2_u2_n140, 
       u1_u2_u2_n141, u1_u2_u2_n142, u1_u2_u2_n143, u1_u2_u2_n144, u1_u2_u2_n145, u1_u2_u2_n146, u1_u2_u2_n147, u1_u2_u2_n148, u1_u2_u2_n149, 
       u1_u2_u2_n150, u1_u2_u2_n151, u1_u2_u2_n152, u1_u2_u2_n153, u1_u2_u2_n154, u1_u2_u2_n155, u1_u2_u2_n156, u1_u2_u2_n157, u1_u2_u2_n158, 
       u1_u2_u2_n159, u1_u2_u2_n160, u1_u2_u2_n161, u1_u2_u2_n162, u1_u2_u2_n163, u1_u2_u2_n164, u1_u2_u2_n165, u1_u2_u2_n166, u1_u2_u2_n167, 
       u1_u2_u2_n168, u1_u2_u2_n169, u1_u2_u2_n170, u1_u2_u2_n171, u1_u2_u2_n172, u1_u2_u2_n173, u1_u2_u2_n174, u1_u2_u2_n175, u1_u2_u2_n176, 
       u1_u2_u2_n177, u1_u2_u2_n178, u1_u2_u2_n179, u1_u2_u2_n180, u1_u2_u2_n181, u1_u2_u2_n182, u1_u2_u2_n183, u1_u2_u2_n184, u1_u2_u2_n185, 
       u1_u2_u2_n186, u1_u2_u2_n187, u1_u2_u2_n188, u1_u2_u2_n95, u1_u2_u2_n96, u1_u2_u2_n97, u1_u2_u2_n98, u1_u2_u2_n99, u1_u2_u5_n100, 
       u1_u2_u5_n101, u1_u2_u5_n102, u1_u2_u5_n103, u1_u2_u5_n104, u1_u2_u5_n105, u1_u2_u5_n106, u1_u2_u5_n107, u1_u2_u5_n108, u1_u2_u5_n109, 
       u1_u2_u5_n110, u1_u2_u5_n111, u1_u2_u5_n112, u1_u2_u5_n113, u1_u2_u5_n114, u1_u2_u5_n115, u1_u2_u5_n116, u1_u2_u5_n117, u1_u2_u5_n118, 
       u1_u2_u5_n119, u1_u2_u5_n120, u1_u2_u5_n121, u1_u2_u5_n122, u1_u2_u5_n123, u1_u2_u5_n124, u1_u2_u5_n125, u1_u2_u5_n126, u1_u2_u5_n127, 
       u1_u2_u5_n128, u1_u2_u5_n129, u1_u2_u5_n130, u1_u2_u5_n131, u1_u2_u5_n132, u1_u2_u5_n133, u1_u2_u5_n134, u1_u2_u5_n135, u1_u2_u5_n136, 
       u1_u2_u5_n137, u1_u2_u5_n138, u1_u2_u5_n139, u1_u2_u5_n140, u1_u2_u5_n141, u1_u2_u5_n142, u1_u2_u5_n143, u1_u2_u5_n144, u1_u2_u5_n145, 
       u1_u2_u5_n146, u1_u2_u5_n147, u1_u2_u5_n148, u1_u2_u5_n149, u1_u2_u5_n150, u1_u2_u5_n151, u1_u2_u5_n152, u1_u2_u5_n153, u1_u2_u5_n154, 
       u1_u2_u5_n155, u1_u2_u5_n156, u1_u2_u5_n157, u1_u2_u5_n158, u1_u2_u5_n159, u1_u2_u5_n160, u1_u2_u5_n161, u1_u2_u5_n162, u1_u2_u5_n163, 
       u1_u2_u5_n164, u1_u2_u5_n165, u1_u2_u5_n166, u1_u2_u5_n167, u1_u2_u5_n168, u1_u2_u5_n169, u1_u2_u5_n170, u1_u2_u5_n171, u1_u2_u5_n172, 
       u1_u2_u5_n173, u1_u2_u5_n174, u1_u2_u5_n175, u1_u2_u5_n176, u1_u2_u5_n177, u1_u2_u5_n178, u1_u2_u5_n179, u1_u2_u5_n180, u1_u2_u5_n181, 
       u1_u2_u5_n182, u1_u2_u5_n183, u1_u2_u5_n184, u1_u2_u5_n185, u1_u2_u5_n186, u1_u2_u5_n187, u1_u2_u5_n188, u1_u2_u5_n189, u1_u2_u5_n190, 
       u1_u2_u5_n191, u1_u2_u5_n192, u1_u2_u5_n193, u1_u2_u5_n194, u1_u2_u5_n195, u1_u2_u5_n196, u1_u2_u5_n99, u1_u3_X_3, u1_u3_X_4, 
       u1_u3_u0_n100, u1_u3_u0_n101, u1_u3_u0_n102, u1_u3_u0_n103, u1_u3_u0_n104, u1_u3_u0_n105, u1_u3_u0_n106, u1_u3_u0_n107, u1_u3_u0_n108, 
       u1_u3_u0_n109, u1_u3_u0_n110, u1_u3_u0_n111, u1_u3_u0_n112, u1_u3_u0_n113, u1_u3_u0_n114, u1_u3_u0_n115, u1_u3_u0_n116, u1_u3_u0_n117, 
       u1_u3_u0_n118, u1_u3_u0_n119, u1_u3_u0_n120, u1_u3_u0_n121, u1_u3_u0_n122, u1_u3_u0_n123, u1_u3_u0_n124, u1_u3_u0_n125, u1_u3_u0_n126, 
       u1_u3_u0_n127, u1_u3_u0_n128, u1_u3_u0_n129, u1_u3_u0_n130, u1_u3_u0_n131, u1_u3_u0_n132, u1_u3_u0_n133, u1_u3_u0_n134, u1_u3_u0_n135, 
       u1_u3_u0_n136, u1_u3_u0_n137, u1_u3_u0_n138, u1_u3_u0_n139, u1_u3_u0_n140, u1_u3_u0_n141, u1_u3_u0_n142, u1_u3_u0_n143, u1_u3_u0_n144, 
       u1_u3_u0_n145, u1_u3_u0_n146, u1_u3_u0_n147, u1_u3_u0_n148, u1_u3_u0_n149, u1_u3_u0_n150, u1_u3_u0_n151, u1_u3_u0_n152, u1_u3_u0_n153, 
       u1_u3_u0_n154, u1_u3_u0_n155, u1_u3_u0_n156, u1_u3_u0_n157, u1_u3_u0_n158, u1_u3_u0_n159, u1_u3_u0_n160, u1_u3_u0_n161, u1_u3_u0_n162, 
       u1_u3_u0_n163, u1_u3_u0_n164, u1_u3_u0_n165, u1_u3_u0_n166, u1_u3_u0_n167, u1_u3_u0_n168, u1_u3_u0_n169, u1_u3_u0_n170, u1_u3_u0_n171, 
       u1_u3_u0_n172, u1_u3_u0_n173, u1_u3_u0_n174, u1_u3_u0_n88, u1_u3_u0_n89, u1_u3_u0_n90, u1_u3_u0_n91, u1_u3_u0_n92, u1_u3_u0_n93, 
       u1_u3_u0_n94, u1_u3_u0_n95, u1_u3_u0_n96, u1_u3_u0_n97, u1_u3_u0_n98, u1_u3_u0_n99, u1_u4_X_10, u1_u4_X_21, u1_u4_X_22, 
       u1_u4_X_3, u1_u4_X_4, u1_u4_X_5, u1_u4_X_7, u1_u4_X_9, u1_u4_u0_n100, u1_u4_u0_n101, u1_u4_u0_n102, u1_u4_u0_n103, 
       u1_u4_u0_n104, u1_u4_u0_n105, u1_u4_u0_n106, u1_u4_u0_n107, u1_u4_u0_n108, u1_u4_u0_n109, u1_u4_u0_n110, u1_u4_u0_n111, u1_u4_u0_n112, 
       u1_u4_u0_n113, u1_u4_u0_n114, u1_u4_u0_n115, u1_u4_u0_n116, u1_u4_u0_n117, u1_u4_u0_n118, u1_u4_u0_n119, u1_u4_u0_n120, u1_u4_u0_n121, 
       u1_u4_u0_n122, u1_u4_u0_n123, u1_u4_u0_n124, u1_u4_u0_n125, u1_u4_u0_n126, u1_u4_u0_n127, u1_u4_u0_n128, u1_u4_u0_n129, u1_u4_u0_n130, 
       u1_u4_u0_n131, u1_u4_u0_n132, u1_u4_u0_n133, u1_u4_u0_n134, u1_u4_u0_n135, u1_u4_u0_n136, u1_u4_u0_n137, u1_u4_u0_n138, u1_u4_u0_n139, 
       u1_u4_u0_n140, u1_u4_u0_n141, u1_u4_u0_n142, u1_u4_u0_n143, u1_u4_u0_n144, u1_u4_u0_n145, u1_u4_u0_n146, u1_u4_u0_n147, u1_u4_u0_n148, 
       u1_u4_u0_n149, u1_u4_u0_n150, u1_u4_u0_n151, u1_u4_u0_n152, u1_u4_u0_n153, u1_u4_u0_n154, u1_u4_u0_n155, u1_u4_u0_n156, u1_u4_u0_n157, 
       u1_u4_u0_n158, u1_u4_u0_n159, u1_u4_u0_n160, u1_u4_u0_n161, u1_u4_u0_n162, u1_u4_u0_n163, u1_u4_u0_n164, u1_u4_u0_n165, u1_u4_u0_n166, 
       u1_u4_u0_n167, u1_u4_u0_n168, u1_u4_u0_n169, u1_u4_u0_n170, u1_u4_u0_n171, u1_u4_u0_n172, u1_u4_u0_n173, u1_u4_u0_n174, u1_u4_u0_n88, 
       u1_u4_u0_n89, u1_u4_u0_n90, u1_u4_u0_n91, u1_u4_u0_n92, u1_u4_u0_n93, u1_u4_u0_n94, u1_u4_u0_n95, u1_u4_u0_n96, u1_u4_u0_n97, 
       u1_u4_u0_n98, u1_u4_u0_n99, u1_u4_u1_n100, u1_u4_u1_n101, u1_u4_u1_n102, u1_u4_u1_n103, u1_u4_u1_n104, u1_u4_u1_n105, u1_u4_u1_n106, 
       u1_u4_u1_n107, u1_u4_u1_n108, u1_u4_u1_n109, u1_u4_u1_n110, u1_u4_u1_n111, u1_u4_u1_n112, u1_u4_u1_n113, u1_u4_u1_n114, u1_u4_u1_n115, 
       u1_u4_u1_n116, u1_u4_u1_n117, u1_u4_u1_n118, u1_u4_u1_n119, u1_u4_u1_n120, u1_u4_u1_n121, u1_u4_u1_n122, u1_u4_u1_n123, u1_u4_u1_n124, 
       u1_u4_u1_n125, u1_u4_u1_n126, u1_u4_u1_n127, u1_u4_u1_n128, u1_u4_u1_n129, u1_u4_u1_n130, u1_u4_u1_n131, u1_u4_u1_n132, u1_u4_u1_n133, 
       u1_u4_u1_n134, u1_u4_u1_n135, u1_u4_u1_n136, u1_u4_u1_n137, u1_u4_u1_n138, u1_u4_u1_n139, u1_u4_u1_n140, u1_u4_u1_n141, u1_u4_u1_n142, 
       u1_u4_u1_n143, u1_u4_u1_n144, u1_u4_u1_n145, u1_u4_u1_n146, u1_u4_u1_n147, u1_u4_u1_n148, u1_u4_u1_n149, u1_u4_u1_n150, u1_u4_u1_n151, 
       u1_u4_u1_n152, u1_u4_u1_n153, u1_u4_u1_n154, u1_u4_u1_n155, u1_u4_u1_n156, u1_u4_u1_n157, u1_u4_u1_n158, u1_u4_u1_n159, u1_u4_u1_n160, 
       u1_u4_u1_n161, u1_u4_u1_n162, u1_u4_u1_n163, u1_u4_u1_n164, u1_u4_u1_n165, u1_u4_u1_n166, u1_u4_u1_n167, u1_u4_u1_n168, u1_u4_u1_n169, 
       u1_u4_u1_n170, u1_u4_u1_n171, u1_u4_u1_n172, u1_u4_u1_n173, u1_u4_u1_n174, u1_u4_u1_n175, u1_u4_u1_n176, u1_u4_u1_n177, u1_u4_u1_n178, 
       u1_u4_u1_n179, u1_u4_u1_n180, u1_u4_u1_n181, u1_u4_u1_n182, u1_u4_u1_n183, u1_u4_u1_n184, u1_u4_u1_n185, u1_u4_u1_n186, u1_u4_u1_n187, 
       u1_u4_u1_n188, u1_u4_u1_n95, u1_u4_u1_n96, u1_u4_u1_n97, u1_u4_u1_n98, u1_u4_u1_n99, u1_u4_u3_n100, u1_u4_u3_n101, u1_u4_u3_n102, 
       u1_u4_u3_n103, u1_u4_u3_n104, u1_u4_u3_n105, u1_u4_u3_n106, u1_u4_u3_n107, u1_u4_u3_n108, u1_u4_u3_n109, u1_u4_u3_n110, u1_u4_u3_n111, 
       u1_u4_u3_n112, u1_u4_u3_n113, u1_u4_u3_n114, u1_u4_u3_n115, u1_u4_u3_n116, u1_u4_u3_n117, u1_u4_u3_n118, u1_u4_u3_n119, u1_u4_u3_n120, 
       u1_u4_u3_n121, u1_u4_u3_n122, u1_u4_u3_n123, u1_u4_u3_n124, u1_u4_u3_n125, u1_u4_u3_n126, u1_u4_u3_n127, u1_u4_u3_n128, u1_u4_u3_n129, 
       u1_u4_u3_n130, u1_u4_u3_n131, u1_u4_u3_n132, u1_u4_u3_n133, u1_u4_u3_n134, u1_u4_u3_n135, u1_u4_u3_n136, u1_u4_u3_n137, u1_u4_u3_n138, 
       u1_u4_u3_n139, u1_u4_u3_n140, u1_u4_u3_n141, u1_u4_u3_n142, u1_u4_u3_n143, u1_u4_u3_n144, u1_u4_u3_n145, u1_u4_u3_n146, u1_u4_u3_n147, 
       u1_u4_u3_n148, u1_u4_u3_n149, u1_u4_u3_n150, u1_u4_u3_n151, u1_u4_u3_n152, u1_u4_u3_n153, u1_u4_u3_n154, u1_u4_u3_n155, u1_u4_u3_n156, 
       u1_u4_u3_n157, u1_u4_u3_n158, u1_u4_u3_n159, u1_u4_u3_n160, u1_u4_u3_n161, u1_u4_u3_n162, u1_u4_u3_n163, u1_u4_u3_n164, u1_u4_u3_n165, 
       u1_u4_u3_n166, u1_u4_u3_n167, u1_u4_u3_n168, u1_u4_u3_n169, u1_u4_u3_n170, u1_u4_u3_n171, u1_u4_u3_n172, u1_u4_u3_n173, u1_u4_u3_n174, 
       u1_u4_u3_n175, u1_u4_u3_n176, u1_u4_u3_n177, u1_u4_u3_n178, u1_u4_u3_n179, u1_u4_u3_n180, u1_u4_u3_n181, u1_u4_u3_n182, u1_u4_u3_n183, 
       u1_u4_u3_n184, u1_u4_u3_n185, u1_u4_u3_n186, u1_u4_u3_n94, u1_u4_u3_n95, u1_u4_u3_n96, u1_u4_u3_n97, u1_u4_u3_n98, u1_u4_u3_n99, 
       u1_u6_X_27, u1_u6_X_28, u1_u6_X_3, u1_u6_X_39, u1_u6_X_4, u1_u6_X_40, u1_u6_u0_n100, u1_u6_u0_n101, u1_u6_u0_n102, 
       u1_u6_u0_n103, u1_u6_u0_n104, u1_u6_u0_n105, u1_u6_u0_n106, u1_u6_u0_n107, u1_u6_u0_n108, u1_u6_u0_n109, u1_u6_u0_n110, u1_u6_u0_n111, 
       u1_u6_u0_n112, u1_u6_u0_n113, u1_u6_u0_n114, u1_u6_u0_n115, u1_u6_u0_n116, u1_u6_u0_n117, u1_u6_u0_n118, u1_u6_u0_n119, u1_u6_u0_n120, 
       u1_u6_u0_n121, u1_u6_u0_n122, u1_u6_u0_n123, u1_u6_u0_n124, u1_u6_u0_n125, u1_u6_u0_n126, u1_u6_u0_n127, u1_u6_u0_n128, u1_u6_u0_n129, 
       u1_u6_u0_n130, u1_u6_u0_n131, u1_u6_u0_n132, u1_u6_u0_n133, u1_u6_u0_n134, u1_u6_u0_n135, u1_u6_u0_n136, u1_u6_u0_n137, u1_u6_u0_n138, 
       u1_u6_u0_n139, u1_u6_u0_n140, u1_u6_u0_n141, u1_u6_u0_n142, u1_u6_u0_n143, u1_u6_u0_n144, u1_u6_u0_n145, u1_u6_u0_n146, u1_u6_u0_n147, 
       u1_u6_u0_n148, u1_u6_u0_n149, u1_u6_u0_n150, u1_u6_u0_n151, u1_u6_u0_n152, u1_u6_u0_n153, u1_u6_u0_n154, u1_u6_u0_n155, u1_u6_u0_n156, 
       u1_u6_u0_n157, u1_u6_u0_n158, u1_u6_u0_n159, u1_u6_u0_n160, u1_u6_u0_n161, u1_u6_u0_n162, u1_u6_u0_n163, u1_u6_u0_n164, u1_u6_u0_n165, 
       u1_u6_u0_n166, u1_u6_u0_n167, u1_u6_u0_n168, u1_u6_u0_n169, u1_u6_u0_n170, u1_u6_u0_n171, u1_u6_u0_n172, u1_u6_u0_n173, u1_u6_u0_n174, 
       u1_u6_u0_n88, u1_u6_u0_n89, u1_u6_u0_n90, u1_u6_u0_n91, u1_u6_u0_n92, u1_u6_u0_n93, u1_u6_u0_n94, u1_u6_u0_n95, u1_u6_u0_n96, 
       u1_u6_u0_n97, u1_u6_u0_n98, u1_u6_u0_n99, u1_u6_u4_n100, u1_u6_u4_n101, u1_u6_u4_n102, u1_u6_u4_n103, u1_u6_u4_n104, u1_u6_u4_n105, 
       u1_u6_u4_n106, u1_u6_u4_n107, u1_u6_u4_n108, u1_u6_u4_n109, u1_u6_u4_n110, u1_u6_u4_n111, u1_u6_u4_n112, u1_u6_u4_n113, u1_u6_u4_n114, 
       u1_u6_u4_n115, u1_u6_u4_n116, u1_u6_u4_n117, u1_u6_u4_n118, u1_u6_u4_n119, u1_u6_u4_n120, u1_u6_u4_n121, u1_u6_u4_n122, u1_u6_u4_n123, 
       u1_u6_u4_n124, u1_u6_u4_n125, u1_u6_u4_n126, u1_u6_u4_n127, u1_u6_u4_n128, u1_u6_u4_n129, u1_u6_u4_n130, u1_u6_u4_n131, u1_u6_u4_n132, 
       u1_u6_u4_n133, u1_u6_u4_n134, u1_u6_u4_n135, u1_u6_u4_n136, u1_u6_u4_n137, u1_u6_u4_n138, u1_u6_u4_n139, u1_u6_u4_n140, u1_u6_u4_n141, 
       u1_u6_u4_n142, u1_u6_u4_n143, u1_u6_u4_n144, u1_u6_u4_n145, u1_u6_u4_n146, u1_u6_u4_n147, u1_u6_u4_n148, u1_u6_u4_n149, u1_u6_u4_n150, 
       u1_u6_u4_n151, u1_u6_u4_n152, u1_u6_u4_n153, u1_u6_u4_n154, u1_u6_u4_n155, u1_u6_u4_n156, u1_u6_u4_n157, u1_u6_u4_n158, u1_u6_u4_n159, 
       u1_u6_u4_n160, u1_u6_u4_n161, u1_u6_u4_n162, u1_u6_u4_n163, u1_u6_u4_n164, u1_u6_u4_n165, u1_u6_u4_n166, u1_u6_u4_n167, u1_u6_u4_n168, 
       u1_u6_u4_n169, u1_u6_u4_n170, u1_u6_u4_n171, u1_u6_u4_n172, u1_u6_u4_n173, u1_u6_u4_n174, u1_u6_u4_n175, u1_u6_u4_n176, u1_u6_u4_n177, 
       u1_u6_u4_n178, u1_u6_u4_n179, u1_u6_u4_n180, u1_u6_u4_n181, u1_u6_u4_n182, u1_u6_u4_n183, u1_u6_u4_n184, u1_u6_u4_n185, u1_u6_u4_n186, 
       u1_u6_u4_n94, u1_u6_u4_n95, u1_u6_u4_n96, u1_u6_u4_n97, u1_u6_u4_n98, u1_u6_u4_n99, u1_u6_u6_n100, u1_u6_u6_n101, u1_u6_u6_n102, 
       u1_u6_u6_n103, u1_u6_u6_n104, u1_u6_u6_n105, u1_u6_u6_n106, u1_u6_u6_n107, u1_u6_u6_n108, u1_u6_u6_n109, u1_u6_u6_n110, u1_u6_u6_n111, 
       u1_u6_u6_n112, u1_u6_u6_n113, u1_u6_u6_n114, u1_u6_u6_n115, u1_u6_u6_n116, u1_u6_u6_n117, u1_u6_u6_n118, u1_u6_u6_n119, u1_u6_u6_n120, 
       u1_u6_u6_n121, u1_u6_u6_n122, u1_u6_u6_n123, u1_u6_u6_n124, u1_u6_u6_n125, u1_u6_u6_n126, u1_u6_u6_n127, u1_u6_u6_n128, u1_u6_u6_n129, 
       u1_u6_u6_n130, u1_u6_u6_n131, u1_u6_u6_n132, u1_u6_u6_n133, u1_u6_u6_n134, u1_u6_u6_n135, u1_u6_u6_n136, u1_u6_u6_n137, u1_u6_u6_n138, 
       u1_u6_u6_n139, u1_u6_u6_n140, u1_u6_u6_n141, u1_u6_u6_n142, u1_u6_u6_n143, u1_u6_u6_n144, u1_u6_u6_n145, u1_u6_u6_n146, u1_u6_u6_n147, 
       u1_u6_u6_n148, u1_u6_u6_n149, u1_u6_u6_n150, u1_u6_u6_n151, u1_u6_u6_n152, u1_u6_u6_n153, u1_u6_u6_n154, u1_u6_u6_n155, u1_u6_u6_n156, 
       u1_u6_u6_n157, u1_u6_u6_n158, u1_u6_u6_n159, u1_u6_u6_n160, u1_u6_u6_n161, u1_u6_u6_n162, u1_u6_u6_n163, u1_u6_u6_n164, u1_u6_u6_n165, 
       u1_u6_u6_n166, u1_u6_u6_n167, u1_u6_u6_n168, u1_u6_u6_n169, u1_u6_u6_n170, u1_u6_u6_n171, u1_u6_u6_n172, u1_u6_u6_n173, u1_u6_u6_n174, 
       u1_u6_u6_n88, u1_u6_u6_n89, u1_u6_u6_n90, u1_u6_u6_n91, u1_u6_u6_n92, u1_u6_u6_n93, u1_u6_u6_n94, u1_u6_u6_n95, u1_u6_u6_n96, 
       u1_u6_u6_n97, u1_u6_u6_n98, u1_u6_u6_n99, u1_u7_X_21, u1_u7_X_22, u1_u7_u3_n100, u1_u7_u3_n101, u1_u7_u3_n102, u1_u7_u3_n103, 
       u1_u7_u3_n104, u1_u7_u3_n105, u1_u7_u3_n106, u1_u7_u3_n107, u1_u7_u3_n108, u1_u7_u3_n109, u1_u7_u3_n110, u1_u7_u3_n111, u1_u7_u3_n112, 
       u1_u7_u3_n113, u1_u7_u3_n114, u1_u7_u3_n115, u1_u7_u3_n116, u1_u7_u3_n117, u1_u7_u3_n118, u1_u7_u3_n119, u1_u7_u3_n120, u1_u7_u3_n121, 
       u1_u7_u3_n122, u1_u7_u3_n123, u1_u7_u3_n124, u1_u7_u3_n125, u1_u7_u3_n126, u1_u7_u3_n127, u1_u7_u3_n128, u1_u7_u3_n129, u1_u7_u3_n130, 
       u1_u7_u3_n131, u1_u7_u3_n132, u1_u7_u3_n133, u1_u7_u3_n134, u1_u7_u3_n135, u1_u7_u3_n136, u1_u7_u3_n137, u1_u7_u3_n138, u1_u7_u3_n139, 
       u1_u7_u3_n140, u1_u7_u3_n141, u1_u7_u3_n142, u1_u7_u3_n143, u1_u7_u3_n144, u1_u7_u3_n145, u1_u7_u3_n146, u1_u7_u3_n147, u1_u7_u3_n148, 
       u1_u7_u3_n149, u1_u7_u3_n150, u1_u7_u3_n151, u1_u7_u3_n152, u1_u7_u3_n153, u1_u7_u3_n154, u1_u7_u3_n155, u1_u7_u3_n156, u1_u7_u3_n157, 
       u1_u7_u3_n158, u1_u7_u3_n159, u1_u7_u3_n160, u1_u7_u3_n161, u1_u7_u3_n162, u1_u7_u3_n163, u1_u7_u3_n164, u1_u7_u3_n165, u1_u7_u3_n166, 
       u1_u7_u3_n167, u1_u7_u3_n168, u1_u7_u3_n169, u1_u7_u3_n170, u1_u7_u3_n171, u1_u7_u3_n172, u1_u7_u3_n173, u1_u7_u3_n174, u1_u7_u3_n175, 
       u1_u7_u3_n176, u1_u7_u3_n177, u1_u7_u3_n178, u1_u7_u3_n179, u1_u7_u3_n180, u1_u7_u3_n181, u1_u7_u3_n182, u1_u7_u3_n183, u1_u7_u3_n184, 
       u1_u7_u3_n185, u1_u7_u3_n186, u1_u7_u3_n94, u1_u7_u3_n95, u1_u7_u3_n96, u1_u7_u3_n97, u1_u7_u3_n98, u1_u7_u3_n99, u1_u8_X_33, 
       u1_u8_X_34, u1_u8_u5_n100, u1_u8_u5_n101, u1_u8_u5_n102, u1_u8_u5_n103, u1_u8_u5_n104, u1_u8_u5_n105, u1_u8_u5_n106, u1_u8_u5_n107, 
       u1_u8_u5_n108, u1_u8_u5_n109, u1_u8_u5_n110, u1_u8_u5_n111, u1_u8_u5_n112, u1_u8_u5_n113, u1_u8_u5_n114, u1_u8_u5_n115, u1_u8_u5_n116, 
       u1_u8_u5_n117, u1_u8_u5_n118, u1_u8_u5_n119, u1_u8_u5_n120, u1_u8_u5_n121, u1_u8_u5_n122, u1_u8_u5_n123, u1_u8_u5_n124, u1_u8_u5_n125, 
       u1_u8_u5_n126, u1_u8_u5_n127, u1_u8_u5_n128, u1_u8_u5_n129, u1_u8_u5_n130, u1_u8_u5_n131, u1_u8_u5_n132, u1_u8_u5_n133, u1_u8_u5_n134, 
       u1_u8_u5_n135, u1_u8_u5_n136, u1_u8_u5_n137, u1_u8_u5_n138, u1_u8_u5_n139, u1_u8_u5_n140, u1_u8_u5_n141, u1_u8_u5_n142, u1_u8_u5_n143, 
       u1_u8_u5_n144, u1_u8_u5_n145, u1_u8_u5_n146, u1_u8_u5_n147, u1_u8_u5_n148, u1_u8_u5_n149, u1_u8_u5_n150, u1_u8_u5_n151, u1_u8_u5_n152, 
       u1_u8_u5_n153, u1_u8_u5_n154, u1_u8_u5_n155, u1_u8_u5_n156, u1_u8_u5_n157, u1_u8_u5_n158, u1_u8_u5_n159, u1_u8_u5_n160, u1_u8_u5_n161, 
       u1_u8_u5_n162, u1_u8_u5_n163, u1_u8_u5_n164, u1_u8_u5_n165, u1_u8_u5_n166, u1_u8_u5_n167, u1_u8_u5_n168, u1_u8_u5_n169, u1_u8_u5_n170, 
       u1_u8_u5_n171, u1_u8_u5_n172, u1_u8_u5_n173, u1_u8_u5_n174, u1_u8_u5_n175, u1_u8_u5_n176, u1_u8_u5_n177, u1_u8_u5_n178, u1_u8_u5_n179, 
       u1_u8_u5_n180, u1_u8_u5_n181, u1_u8_u5_n182, u1_u8_u5_n183, u1_u8_u5_n184, u1_u8_u5_n185, u1_u8_u5_n186, u1_u8_u5_n187, u1_u8_u5_n188, 
       u1_u8_u5_n189, u1_u8_u5_n190, u1_u8_u5_n191, u1_u8_u5_n192, u1_u8_u5_n193, u1_u8_u5_n194, u1_u8_u5_n195, u1_u8_u5_n196, u1_u8_u5_n99, 
       u1_u9_X_27, u1_u9_X_28, u1_u9_u4_n100, u1_u9_u4_n101, u1_u9_u4_n102, u1_u9_u4_n103, u1_u9_u4_n104, u1_u9_u4_n105, u1_u9_u4_n106, 
       u1_u9_u4_n107, u1_u9_u4_n108, u1_u9_u4_n109, u1_u9_u4_n110, u1_u9_u4_n111, u1_u9_u4_n112, u1_u9_u4_n113, u1_u9_u4_n114, u1_u9_u4_n115, 
       u1_u9_u4_n116, u1_u9_u4_n117, u1_u9_u4_n118, u1_u9_u4_n119, u1_u9_u4_n120, u1_u9_u4_n121, u1_u9_u4_n122, u1_u9_u4_n123, u1_u9_u4_n124, 
       u1_u9_u4_n125, u1_u9_u4_n126, u1_u9_u4_n127, u1_u9_u4_n128, u1_u9_u4_n129, u1_u9_u4_n130, u1_u9_u4_n131, u1_u9_u4_n132, u1_u9_u4_n133, 
       u1_u9_u4_n134, u1_u9_u4_n135, u1_u9_u4_n136, u1_u9_u4_n137, u1_u9_u4_n138, u1_u9_u4_n139, u1_u9_u4_n140, u1_u9_u4_n141, u1_u9_u4_n142, 
       u1_u9_u4_n143, u1_u9_u4_n144, u1_u9_u4_n145, u1_u9_u4_n146, u1_u9_u4_n147, u1_u9_u4_n148, u1_u9_u4_n149, u1_u9_u4_n150, u1_u9_u4_n151, 
       u1_u9_u4_n152, u1_u9_u4_n153, u1_u9_u4_n154, u1_u9_u4_n155, u1_u9_u4_n156, u1_u9_u4_n157, u1_u9_u4_n158, u1_u9_u4_n159, u1_u9_u4_n160, 
       u1_u9_u4_n161, u1_u9_u4_n162, u1_u9_u4_n163, u1_u9_u4_n164, u1_u9_u4_n165, u1_u9_u4_n166, u1_u9_u4_n167, u1_u9_u4_n168, u1_u9_u4_n169, 
       u1_u9_u4_n170, u1_u9_u4_n171, u1_u9_u4_n172, u1_u9_u4_n173, u1_u9_u4_n174, u1_u9_u4_n175, u1_u9_u4_n176, u1_u9_u4_n177, u1_u9_u4_n178, 
       u1_u9_u4_n179, u1_u9_u4_n180, u1_u9_u4_n181, u1_u9_u4_n182, u1_u9_u4_n183, u1_u9_u4_n184, u1_u9_u4_n185, u1_u9_u4_n186, u1_u9_u4_n94, 
       u1_u9_u4_n95, u1_u9_u4_n96, u1_u9_u4_n97, u1_u9_u4_n98, u1_u9_u4_n99, u2_K8_19, u2_K8_20, u2_K8_21, u2_K8_22, 
       u2_K8_23, u2_out7_1, u2_out7_10, u2_out7_20, u2_out7_26, u2_u7_X_19, u2_u7_X_20, u2_u7_X_21, u2_u7_X_22, 
       u2_u7_X_23, u2_u7_X_24, u2_u7_u3_n100, u2_u7_u3_n101, u2_u7_u3_n102, u2_u7_u3_n103, u2_u7_u3_n104, u2_u7_u3_n105, u2_u7_u3_n106, 
       u2_u7_u3_n107, u2_u7_u3_n108, u2_u7_u3_n109, u2_u7_u3_n110, u2_u7_u3_n111, u2_u7_u3_n112, u2_u7_u3_n113, u2_u7_u3_n114, u2_u7_u3_n115, 
       u2_u7_u3_n116, u2_u7_u3_n117, u2_u7_u3_n118, u2_u7_u3_n119, u2_u7_u3_n120, u2_u7_u3_n121, u2_u7_u3_n122, u2_u7_u3_n123, u2_u7_u3_n124, 
       u2_u7_u3_n125, u2_u7_u3_n126, u2_u7_u3_n127, u2_u7_u3_n128, u2_u7_u3_n129, u2_u7_u3_n130, u2_u7_u3_n131, u2_u7_u3_n132, u2_u7_u3_n133, 
       u2_u7_u3_n134, u2_u7_u3_n135, u2_u7_u3_n136, u2_u7_u3_n137, u2_u7_u3_n138, u2_u7_u3_n139, u2_u7_u3_n140, u2_u7_u3_n141, u2_u7_u3_n142, 
       u2_u7_u3_n143, u2_u7_u3_n144, u2_u7_u3_n145, u2_u7_u3_n146, u2_u7_u3_n147, u2_u7_u3_n148, u2_u7_u3_n149, u2_u7_u3_n150, u2_u7_u3_n151, 
       u2_u7_u3_n152, u2_u7_u3_n153, u2_u7_u3_n154, u2_u7_u3_n155, u2_u7_u3_n156, u2_u7_u3_n157, u2_u7_u3_n158, u2_u7_u3_n159, u2_u7_u3_n160, 
       u2_u7_u3_n161, u2_u7_u3_n162, u2_u7_u3_n163, u2_u7_u3_n164, u2_u7_u3_n165, u2_u7_u3_n166, u2_u7_u3_n167, u2_u7_u3_n168, u2_u7_u3_n169, 
       u2_u7_u3_n170, u2_u7_u3_n171, u2_u7_u3_n172, u2_u7_u3_n173, u2_u7_u3_n174, u2_u7_u3_n175, u2_u7_u3_n176, u2_u7_u3_n177, u2_u7_u3_n178, 
       u2_u7_u3_n179, u2_u7_u3_n180, u2_u7_u3_n181, u2_u7_u3_n182, u2_u7_u3_n183, u2_u7_u3_n184, u2_u7_u3_n185, u2_u7_u3_n186, u2_u7_u3_n94, 
       u2_u7_u3_n95, u2_u7_u3_n96, u2_u7_u3_n97, u2_u7_u3_n98,  u2_u7_u3_n99;
  XOR2_X1 u0_U138 (.B( u0_L11_25 ) , .Z( u0_N408 ) , .A( u0_out12_25 ) );
  XOR2_X1 u0_U151 (.B( u0_L11_14 ) , .Z( u0_N397 ) , .A( u0_out12_14 ) );
  XOR2_X1 u0_U157 (.B( u0_L11_8 ) , .Z( u0_N391 ) , .A( u0_out12_8 ) );
  XOR2_X1 u0_U163 (.B( u0_L11_3 ) , .Z( u0_N386 ) , .A( u0_out12_3 ) );
  XOR2_X1 u0_U192 (.B( u0_L0_5 ) , .Z( u0_N36 ) , .A( u0_out1_5 ) );
  XOR2_X1 u0_U209 (.B( u0_L9_25 ) , .Z( u0_N344 ) , .A( u0_out10_25 ) );
  XOR2_X1 u0_U221 (.B( u0_L9_14 ) , .Z( u0_N333 ) , .A( u0_out10_14 ) );
  XOR2_X1 u0_U228 (.B( u0_L9_8 ) , .Z( u0_N327 ) , .A( u0_out10_8 ) );
  XOR2_X1 u0_U233 (.B( u0_L9_3 ) , .Z( u0_N322 ) , .A( u0_out10_3 ) );
  XOR2_X1 u0_U239 (.B( u0_L8_30 ) , .Z( u0_N317 ) , .A( u0_out9_30 ) );
  XOR2_X1 u0_U241 (.B( u0_L8_28 ) , .Z( u0_N315 ) , .A( u0_out9_28 ) );
  XOR2_X1 u0_U243 (.B( u0_L8_26 ) , .Z( u0_N313 ) , .A( u0_out9_26 ) );
  XOR2_X1 u0_U245 (.B( u0_L8_24 ) , .Z( u0_N311 ) , .A( u0_out9_24 ) );
  XOR2_X1 u0_U250 (.B( u0_L8_20 ) , .Z( u0_N307 ) , .A( u0_out9_20 ) );
  XOR2_X1 u0_U252 (.B( u0_L8_18 ) , .Z( u0_N305 ) , .A( u0_out9_18 ) );
  XOR2_X1 u0_U254 (.B( u0_L8_16 ) , .Z( u0_N303 ) , .A( u0_out9_16 ) );
  XOR2_X1 u0_U257 (.B( u0_L8_13 ) , .Z( u0_N300 ) , .A( u0_out9_13 ) );
  XOR2_X1 u0_U262 (.B( u0_L8_10 ) , .Z( u0_N297 ) , .A( u0_out9_10 ) );
  XOR2_X1 u0_U266 (.B( u0_L8_6 ) , .Z( u0_N293 ) , .A( u0_out9_6 ) );
  XOR2_X1 u0_U271 (.B( u0_L8_2 ) , .Z( u0_N289 ) , .A( u0_out9_2 ) );
  XOR2_X1 u0_U272 (.B( u0_L8_1 ) , .Z( u0_N288 ) , .A( u0_out9_1 ) );
  XOR2_X1 u0_U274 (.B( u0_L7_31 ) , .Z( u0_N286 ) , .A( u0_out8_31 ) );
  XOR2_X1 u0_U275 (.B( u0_L7_30 ) , .Z( u0_N285 ) , .A( u0_out8_30 ) );
  XOR2_X1 u0_U277 (.B( u0_L7_28 ) , .Z( u0_N283 ) , .A( u0_out8_28 ) );
  XOR2_X1 u0_U278 (.B( u0_L7_27 ) , .Z( u0_N282 ) , .A( u0_out8_27 ) );
  XOR2_X1 u0_U279 (.B( u0_L7_26 ) , .Z( u0_N281 ) , .A( u0_out8_26 ) );
  XOR2_X1 u0_U280 (.B( u0_L7_25 ) , .Z( u0_N280 ) , .A( u0_out8_25 ) );
  XOR2_X1 u0_U282 (.B( u0_L7_24 ) , .Z( u0_N279 ) , .A( u0_out8_24 ) );
  XOR2_X1 u0_U283 (.B( u0_L7_23 ) , .Z( u0_N278 ) , .A( u0_out8_23 ) );
  XOR2_X1 u0_U285 (.B( u0_L7_21 ) , .Z( u0_N276 ) , .A( u0_out8_21 ) );
  XOR2_X1 u0_U286 (.B( u0_L7_20 ) , .Z( u0_N275 ) , .A( u0_out8_20 ) );
  XOR2_X1 u0_U288 (.B( u0_L7_18 ) , .Z( u0_N273 ) , .A( u0_out8_18 ) );
  XOR2_X1 u0_U289 (.B( u0_L7_17 ) , .Z( u0_N272 ) , .A( u0_out8_17 ) );
  XOR2_X1 u0_U290 (.B( u0_L7_16 ) , .Z( u0_N271 ) , .A( u0_out8_16 ) );
  XOR2_X1 u0_U291 (.B( u0_L7_15 ) , .Z( u0_N270 ) , .A( u0_out8_15 ) );
  XOR2_X1 u0_U293 (.B( u0_L7_14 ) , .Z( u0_N269 ) , .A( u0_out8_14 ) );
  XOR2_X1 u0_U294 (.B( u0_L7_13 ) , .Z( u0_N268 ) , .A( u0_out8_13 ) );
  XOR2_X1 u0_U297 (.B( u0_L7_10 ) , .Z( u0_N265 ) , .A( u0_out8_10 ) );
  XOR2_X1 u0_U298 (.B( u0_L7_9 ) , .Z( u0_N264 ) , .A( u0_out8_9 ) );
  XOR2_X1 u0_U299 (.B( u0_L7_8 ) , .Z( u0_N263 ) , .A( u0_out8_8 ) );
  XOR2_X1 u0_U301 (.B( u0_L7_6 ) , .Z( u0_N261 ) , .A( u0_out8_6 ) );
  XOR2_X1 u0_U302 (.B( u0_L7_5 ) , .Z( u0_N260 ) , .A( u0_out8_5 ) );
  XOR2_X1 u0_U305 (.B( u0_L7_3 ) , .Z( u0_N258 ) , .A( u0_out8_3 ) );
  XOR2_X1 u0_U306 (.B( u0_L7_2 ) , .Z( u0_N257 ) , .A( u0_out8_2 ) );
  XOR2_X1 u0_U307 (.B( u0_L7_1 ) , .Z( u0_N256 ) , .A( u0_out8_1 ) );
  XOR2_X1 u0_U350 (.B( u0_L5_26 ) , .Z( u0_N217 ) , .A( u0_out6_26 ) );
  XOR2_X1 u0_U351 (.B( u0_L5_25 ) , .Z( u0_N216 ) , .A( u0_out6_25 ) );
  XOR2_X1 u0_U356 (.B( u0_L5_20 ) , .Z( u0_N211 ) , .A( u0_out6_20 ) );
  XOR2_X1 u0_U363 (.B( u0_L5_14 ) , .Z( u0_N205 ) , .A( u0_out6_14 ) );
  XOR2_X1 u0_U367 (.B( u0_L5_10 ) , .Z( u0_N201 ) , .A( u0_out6_10 ) );
  XOR2_X1 u0_U371 (.B( u0_L5_8 ) , .Z( u0_N199 ) , .A( u0_out6_8 ) );
  XOR2_X1 u0_U376 (.B( u0_L5_3 ) , .Z( u0_N194 ) , .A( u0_out6_3 ) );
  XOR2_X1 u0_U378 (.B( u0_L5_1 ) , .Z( u0_N192 ) , .A( u0_out6_1 ) );
  XOR2_X1 u0_U379 (.B( u0_L4_32 ) , .Z( u0_N191 ) , .A( u0_out5_32 ) );
  XOR2_X1 u0_U387 (.B( u0_L4_25 ) , .Z( u0_N184 ) , .A( u0_out5_25 ) );
  XOR2_X1 u0_U390 (.B( u0_L4_22 ) , .Z( u0_N181 ) , .A( u0_out5_22 ) );
  XOR2_X1 u0_U399 (.B( u0_L4_14 ) , .Z( u0_N173 ) , .A( u0_out5_14 ) );
  XOR2_X1 u0_U401 (.B( u0_L4_12 ) , .Z( u0_N171 ) , .A( u0_out5_12 ) );
  XOR2_X1 u0_U406 (.B( u0_L4_8 ) , .Z( u0_N167 ) , .A( u0_out5_8 ) );
  XOR2_X1 u0_U407 (.B( u0_L4_7 ) , .Z( u0_N166 ) , .A( u0_out5_7 ) );
  XOR2_X1 u0_U411 (.B( u0_L4_3 ) , .Z( u0_N162 ) , .A( u0_out5_3 ) );
  XOR2_X1 u0_U48 (.B( u0_L0_27 ) , .Z( u0_N58 ) , .A( u0_out1_27 ) );
  XOR2_X1 u0_U485 (.Z( u0_FP_7 ) , .B( u0_L14_7 ) , .A( u0_out15_7 ) );
  XOR2_X1 u0_U487 (.Z( u0_FP_5 ) , .B( u0_L14_5 ) , .A( u0_out15_5 ) );
  XOR2_X1 u0_U488 (.Z( u0_FP_4 ) , .B( u0_L14_4 ) , .A( u0_out15_4 ) );
  XOR2_X1 u0_U490 (.Z( u0_FP_32 ) , .B( u0_L14_32 ) , .A( u0_out15_32 ) );
  XOR2_X1 u0_U494 (.Z( u0_FP_29 ) , .B( u0_L14_29 ) , .A( u0_out15_29 ) );
  XOR2_X1 u0_U496 (.Z( u0_FP_27 ) , .B( u0_L14_27 ) , .A( u0_out15_27 ) );
  XOR2_X1 u0_U501 (.Z( u0_FP_22 ) , .B( u0_L14_22 ) , .A( u0_out15_22 ) );
  XOR2_X1 u0_U502 (.Z( u0_FP_21 ) , .B( u0_L14_21 ) , .A( u0_out15_21 ) );
  XOR2_X1 u0_U505 (.Z( u0_FP_19 ) , .B( u0_L14_19 ) , .A( u0_out15_19 ) );
  XOR2_X1 u0_U509 (.Z( u0_FP_15 ) , .B( u0_L14_15 ) , .A( u0_out15_15 ) );
  XOR2_X1 u0_U512 (.Z( u0_FP_12 ) , .B( u0_L14_12 ) , .A( u0_out15_12 ) );
  XOR2_X1 u0_U513 (.Z( u0_FP_11 ) , .B( u0_L14_11 ) , .A( u0_out15_11 ) );
  XOR2_X1 u0_U54 (.B( u0_L0_21 ) , .Z( u0_N52 ) , .A( u0_out1_21 ) );
  XOR2_X1 u0_U62 (.B( u0_L13_30 ) , .Z( u0_N477 ) , .A( u0_out14_30 ) );
  XOR2_X1 u0_U63 (.B( u0_L13_29 ) , .Z( u0_N476 ) , .A( u0_out14_29 ) );
  XOR2_X1 u0_U64 (.B( u0_L13_28 ) , .Z( u0_N475 ) , .A( u0_out14_28 ) );
  XOR2_X1 u0_U66 (.B( u0_L13_26 ) , .Z( u0_N473 ) , .A( u0_out14_26 ) );
  XOR2_X1 u0_U68 (.B( u0_L13_24 ) , .Z( u0_N471 ) , .A( u0_out14_24 ) );
  XOR2_X1 u0_U73 (.B( u0_L13_20 ) , .Z( u0_N467 ) , .A( u0_out14_20 ) );
  XOR2_X1 u0_U74 (.B( u0_L13_19 ) , .Z( u0_N466 ) , .A( u0_out14_19 ) );
  XOR2_X1 u0_U75 (.B( u0_L13_18 ) , .Z( u0_N465 ) , .A( u0_out14_18 ) );
  XOR2_X1 u0_U77 (.B( u0_L13_16 ) , .Z( u0_N463 ) , .A( u0_out14_16 ) );
  XOR2_X1 u0_U80 (.B( u0_L13_13 ) , .Z( u0_N460 ) , .A( u0_out14_13 ) );
  XOR2_X1 u0_U81 (.B( u0_L0_15 ) , .Z( u0_N46 ) , .A( u0_out1_15 ) );
  XOR2_X1 u0_U83 (.B( u0_L13_11 ) , .Z( u0_N458 ) , .A( u0_out14_11 ) );
  XOR2_X1 u0_U84 (.B( u0_L13_10 ) , .Z( u0_N457 ) , .A( u0_out14_10 ) );
  XOR2_X1 u0_U88 (.B( u0_L13_6 ) , .Z( u0_N453 ) , .A( u0_out14_6 ) );
  XOR2_X1 u0_U90 (.B( u0_L13_4 ) , .Z( u0_N451 ) , .A( u0_out14_4 ) );
  XOR2_X1 u0_U93 (.B( u0_L13_2 ) , .Z( u0_N449 ) , .A( u0_out14_2 ) );
  XOR2_X1 u0_U94 (.B( u0_L13_1 ) , .Z( u0_N448 ) , .A( u0_out14_1 ) );
  XOR2_X1 u0_u10_U26 (.B( u0_K11_30 ) , .A( u0_R9_21 ) , .Z( u0_u10_X_30 ) );
  XOR2_X1 u0_u10_U28 (.B( u0_K11_29 ) , .A( u0_R9_20 ) , .Z( u0_u10_X_29 ) );
  XOR2_X1 u0_u10_U29 (.B( u0_K11_28 ) , .A( u0_R9_19 ) , .Z( u0_u10_X_28 ) );
  XOR2_X1 u0_u10_U30 (.B( u0_K11_27 ) , .A( u0_R9_18 ) , .Z( u0_u10_X_27 ) );
  XOR2_X1 u0_u10_U31 (.B( u0_K11_26 ) , .A( u0_R9_17 ) , .Z( u0_u10_X_26 ) );
  XOR2_X1 u0_u10_U32 (.B( u0_K11_25 ) , .A( u0_R9_16 ) , .Z( u0_u10_X_25 ) );
  AOI21_X1 u0_u10_u4_U10 (.ZN( u0_u10_u4_n106 ) , .B2( u0_u10_u4_n146 ) , .B1( u0_u10_u4_n158 ) , .A( u0_u10_u4_n170 ) );
  AOI21_X1 u0_u10_u4_U11 (.ZN( u0_u10_u4_n108 ) , .B2( u0_u10_u4_n134 ) , .B1( u0_u10_u4_n155 ) , .A( u0_u10_u4_n156 ) );
  AOI21_X1 u0_u10_u4_U12 (.ZN( u0_u10_u4_n109 ) , .A( u0_u10_u4_n153 ) , .B1( u0_u10_u4_n159 ) , .B2( u0_u10_u4_n184 ) );
  AOI211_X1 u0_u10_u4_U13 (.B( u0_u10_u4_n136 ) , .A( u0_u10_u4_n137 ) , .C2( u0_u10_u4_n138 ) , .ZN( u0_u10_u4_n139 ) , .C1( u0_u10_u4_n182 ) );
  OAI22_X1 u0_u10_u4_U14 (.B2( u0_u10_u4_n135 ) , .ZN( u0_u10_u4_n137 ) , .B1( u0_u10_u4_n153 ) , .A1( u0_u10_u4_n155 ) , .A2( u0_u10_u4_n171 ) );
  AND3_X1 u0_u10_u4_U15 (.A2( u0_u10_u4_n134 ) , .ZN( u0_u10_u4_n135 ) , .A3( u0_u10_u4_n145 ) , .A1( u0_u10_u4_n157 ) );
  NAND2_X1 u0_u10_u4_U16 (.ZN( u0_u10_u4_n132 ) , .A2( u0_u10_u4_n170 ) , .A1( u0_u10_u4_n173 ) );
  AOI21_X1 u0_u10_u4_U17 (.B2( u0_u10_u4_n160 ) , .B1( u0_u10_u4_n161 ) , .ZN( u0_u10_u4_n162 ) , .A( u0_u10_u4_n170 ) );
  AOI21_X1 u0_u10_u4_U18 (.ZN( u0_u10_u4_n107 ) , .B2( u0_u10_u4_n143 ) , .A( u0_u10_u4_n174 ) , .B1( u0_u10_u4_n184 ) );
  AOI21_X1 u0_u10_u4_U19 (.B2( u0_u10_u4_n158 ) , .B1( u0_u10_u4_n159 ) , .ZN( u0_u10_u4_n163 ) , .A( u0_u10_u4_n174 ) );
  AOI21_X1 u0_u10_u4_U20 (.A( u0_u10_u4_n153 ) , .B2( u0_u10_u4_n154 ) , .B1( u0_u10_u4_n155 ) , .ZN( u0_u10_u4_n165 ) );
  AOI21_X1 u0_u10_u4_U21 (.A( u0_u10_u4_n156 ) , .B2( u0_u10_u4_n157 ) , .ZN( u0_u10_u4_n164 ) , .B1( u0_u10_u4_n184 ) );
  INV_X1 u0_u10_u4_U22 (.A( u0_u10_u4_n138 ) , .ZN( u0_u10_u4_n170 ) );
  AND2_X1 u0_u10_u4_U23 (.A2( u0_u10_u4_n120 ) , .ZN( u0_u10_u4_n155 ) , .A1( u0_u10_u4_n160 ) );
  INV_X1 u0_u10_u4_U24 (.A( u0_u10_u4_n156 ) , .ZN( u0_u10_u4_n175 ) );
  NAND2_X1 u0_u10_u4_U25 (.A2( u0_u10_u4_n118 ) , .ZN( u0_u10_u4_n131 ) , .A1( u0_u10_u4_n147 ) );
  NAND2_X1 u0_u10_u4_U26 (.A1( u0_u10_u4_n119 ) , .A2( u0_u10_u4_n120 ) , .ZN( u0_u10_u4_n130 ) );
  NAND2_X1 u0_u10_u4_U27 (.ZN( u0_u10_u4_n117 ) , .A2( u0_u10_u4_n118 ) , .A1( u0_u10_u4_n148 ) );
  NAND2_X1 u0_u10_u4_U28 (.ZN( u0_u10_u4_n129 ) , .A1( u0_u10_u4_n134 ) , .A2( u0_u10_u4_n148 ) );
  AND3_X1 u0_u10_u4_U29 (.A1( u0_u10_u4_n119 ) , .A2( u0_u10_u4_n143 ) , .A3( u0_u10_u4_n154 ) , .ZN( u0_u10_u4_n161 ) );
  NOR2_X1 u0_u10_u4_U3 (.ZN( u0_u10_u4_n121 ) , .A1( u0_u10_u4_n181 ) , .A2( u0_u10_u4_n182 ) );
  AND2_X1 u0_u10_u4_U30 (.A1( u0_u10_u4_n145 ) , .A2( u0_u10_u4_n147 ) , .ZN( u0_u10_u4_n159 ) );
  OR3_X1 u0_u10_u4_U31 (.A3( u0_u10_u4_n114 ) , .A2( u0_u10_u4_n115 ) , .A1( u0_u10_u4_n116 ) , .ZN( u0_u10_u4_n136 ) );
  AOI21_X1 u0_u10_u4_U32 (.A( u0_u10_u4_n113 ) , .ZN( u0_u10_u4_n116 ) , .B2( u0_u10_u4_n173 ) , .B1( u0_u10_u4_n174 ) );
  AOI21_X1 u0_u10_u4_U33 (.ZN( u0_u10_u4_n115 ) , .B2( u0_u10_u4_n145 ) , .B1( u0_u10_u4_n146 ) , .A( u0_u10_u4_n156 ) );
  OAI22_X1 u0_u10_u4_U34 (.ZN( u0_u10_u4_n114 ) , .A2( u0_u10_u4_n121 ) , .B1( u0_u10_u4_n160 ) , .B2( u0_u10_u4_n170 ) , .A1( u0_u10_u4_n171 ) );
  INV_X1 u0_u10_u4_U35 (.A( u0_u10_u4_n158 ) , .ZN( u0_u10_u4_n182 ) );
  INV_X1 u0_u10_u4_U36 (.ZN( u0_u10_u4_n181 ) , .A( u0_u10_u4_n96 ) );
  INV_X1 u0_u10_u4_U37 (.A( u0_u10_u4_n144 ) , .ZN( u0_u10_u4_n179 ) );
  INV_X1 u0_u10_u4_U38 (.A( u0_u10_u4_n157 ) , .ZN( u0_u10_u4_n178 ) );
  NAND2_X1 u0_u10_u4_U39 (.A2( u0_u10_u4_n154 ) , .A1( u0_u10_u4_n96 ) , .ZN( u0_u10_u4_n97 ) );
  INV_X1 u0_u10_u4_U4 (.A( u0_u10_u4_n117 ) , .ZN( u0_u10_u4_n184 ) );
  INV_X1 u0_u10_u4_U40 (.A( u0_u10_u4_n143 ) , .ZN( u0_u10_u4_n183 ) );
  NOR2_X1 u0_u10_u4_U41 (.ZN( u0_u10_u4_n138 ) , .A1( u0_u10_u4_n168 ) , .A2( u0_u10_u4_n169 ) );
  NOR2_X1 u0_u10_u4_U42 (.A1( u0_u10_u4_n150 ) , .A2( u0_u10_u4_n152 ) , .ZN( u0_u10_u4_n153 ) );
  NOR2_X1 u0_u10_u4_U43 (.A2( u0_u10_u4_n128 ) , .A1( u0_u10_u4_n138 ) , .ZN( u0_u10_u4_n156 ) );
  AOI22_X1 u0_u10_u4_U44 (.B2( u0_u10_u4_n122 ) , .A1( u0_u10_u4_n123 ) , .ZN( u0_u10_u4_n124 ) , .B1( u0_u10_u4_n128 ) , .A2( u0_u10_u4_n172 ) );
  INV_X1 u0_u10_u4_U45 (.A( u0_u10_u4_n153 ) , .ZN( u0_u10_u4_n172 ) );
  NAND2_X1 u0_u10_u4_U46 (.A2( u0_u10_u4_n120 ) , .ZN( u0_u10_u4_n123 ) , .A1( u0_u10_u4_n161 ) );
  AOI22_X1 u0_u10_u4_U47 (.B2( u0_u10_u4_n132 ) , .A2( u0_u10_u4_n133 ) , .ZN( u0_u10_u4_n140 ) , .A1( u0_u10_u4_n150 ) , .B1( u0_u10_u4_n179 ) );
  NAND2_X1 u0_u10_u4_U48 (.ZN( u0_u10_u4_n133 ) , .A2( u0_u10_u4_n146 ) , .A1( u0_u10_u4_n154 ) );
  NAND2_X1 u0_u10_u4_U49 (.A1( u0_u10_u4_n103 ) , .ZN( u0_u10_u4_n154 ) , .A2( u0_u10_u4_n98 ) );
  INV_X1 u0_u10_u4_U5 (.ZN( u0_u10_u4_n186 ) , .A( u0_u10_u4_n95 ) );
  NAND2_X1 u0_u10_u4_U50 (.A1( u0_u10_u4_n101 ) , .ZN( u0_u10_u4_n158 ) , .A2( u0_u10_u4_n99 ) );
  AOI21_X1 u0_u10_u4_U51 (.ZN( u0_u10_u4_n127 ) , .A( u0_u10_u4_n136 ) , .B2( u0_u10_u4_n150 ) , .B1( u0_u10_u4_n180 ) );
  INV_X1 u0_u10_u4_U52 (.A( u0_u10_u4_n160 ) , .ZN( u0_u10_u4_n180 ) );
  NAND2_X1 u0_u10_u4_U53 (.A2( u0_u10_u4_n104 ) , .A1( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n146 ) );
  NAND2_X1 u0_u10_u4_U54 (.A2( u0_u10_u4_n101 ) , .A1( u0_u10_u4_n102 ) , .ZN( u0_u10_u4_n160 ) );
  NAND2_X1 u0_u10_u4_U55 (.ZN( u0_u10_u4_n134 ) , .A1( u0_u10_u4_n98 ) , .A2( u0_u10_u4_n99 ) );
  NAND2_X1 u0_u10_u4_U56 (.A1( u0_u10_u4_n103 ) , .A2( u0_u10_u4_n104 ) , .ZN( u0_u10_u4_n143 ) );
  NAND2_X1 u0_u10_u4_U57 (.A2( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n145 ) , .A1( u0_u10_u4_n98 ) );
  NAND2_X1 u0_u10_u4_U58 (.A1( u0_u10_u4_n100 ) , .A2( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n120 ) );
  NAND2_X1 u0_u10_u4_U59 (.A1( u0_u10_u4_n102 ) , .A2( u0_u10_u4_n104 ) , .ZN( u0_u10_u4_n148 ) );
  OAI221_X1 u0_u10_u4_U6 (.C1( u0_u10_u4_n134 ) , .B1( u0_u10_u4_n158 ) , .B2( u0_u10_u4_n171 ) , .C2( u0_u10_u4_n173 ) , .A( u0_u10_u4_n94 ) , .ZN( u0_u10_u4_n95 ) );
  NAND2_X1 u0_u10_u4_U60 (.A2( u0_u10_u4_n100 ) , .A1( u0_u10_u4_n103 ) , .ZN( u0_u10_u4_n157 ) );
  INV_X1 u0_u10_u4_U61 (.A( u0_u10_u4_n150 ) , .ZN( u0_u10_u4_n173 ) );
  INV_X1 u0_u10_u4_U62 (.A( u0_u10_u4_n152 ) , .ZN( u0_u10_u4_n171 ) );
  NAND2_X1 u0_u10_u4_U63 (.A1( u0_u10_u4_n100 ) , .ZN( u0_u10_u4_n118 ) , .A2( u0_u10_u4_n99 ) );
  NAND2_X1 u0_u10_u4_U64 (.A2( u0_u10_u4_n100 ) , .A1( u0_u10_u4_n102 ) , .ZN( u0_u10_u4_n144 ) );
  NAND2_X1 u0_u10_u4_U65 (.A2( u0_u10_u4_n101 ) , .A1( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n96 ) );
  INV_X1 u0_u10_u4_U66 (.A( u0_u10_u4_n128 ) , .ZN( u0_u10_u4_n174 ) );
  NAND2_X1 u0_u10_u4_U67 (.A2( u0_u10_u4_n102 ) , .ZN( u0_u10_u4_n119 ) , .A1( u0_u10_u4_n98 ) );
  NAND2_X1 u0_u10_u4_U68 (.A2( u0_u10_u4_n101 ) , .A1( u0_u10_u4_n103 ) , .ZN( u0_u10_u4_n147 ) );
  NAND2_X1 u0_u10_u4_U69 (.A2( u0_u10_u4_n104 ) , .ZN( u0_u10_u4_n113 ) , .A1( u0_u10_u4_n99 ) );
  AOI222_X1 u0_u10_u4_U7 (.B2( u0_u10_u4_n132 ) , .A1( u0_u10_u4_n138 ) , .C2( u0_u10_u4_n175 ) , .A2( u0_u10_u4_n179 ) , .C1( u0_u10_u4_n181 ) , .B1( u0_u10_u4_n185 ) , .ZN( u0_u10_u4_n94 ) );
  NOR2_X1 u0_u10_u4_U70 (.A2( u0_u10_X_28 ) , .ZN( u0_u10_u4_n150 ) , .A1( u0_u10_u4_n168 ) );
  NOR2_X1 u0_u10_u4_U71 (.A2( u0_u10_X_29 ) , .ZN( u0_u10_u4_n152 ) , .A1( u0_u10_u4_n169 ) );
  NOR2_X1 u0_u10_u4_U72 (.A2( u0_u10_X_30 ) , .ZN( u0_u10_u4_n105 ) , .A1( u0_u10_u4_n176 ) );
  NOR2_X1 u0_u10_u4_U73 (.A2( u0_u10_X_26 ) , .ZN( u0_u10_u4_n100 ) , .A1( u0_u10_u4_n177 ) );
  NOR2_X1 u0_u10_u4_U74 (.A2( u0_u10_X_28 ) , .A1( u0_u10_X_29 ) , .ZN( u0_u10_u4_n128 ) );
  NOR2_X1 u0_u10_u4_U75 (.A2( u0_u10_X_27 ) , .A1( u0_u10_X_30 ) , .ZN( u0_u10_u4_n102 ) );
  NOR2_X1 u0_u10_u4_U76 (.A2( u0_u10_X_25 ) , .A1( u0_u10_X_26 ) , .ZN( u0_u10_u4_n98 ) );
  AND2_X1 u0_u10_u4_U77 (.A2( u0_u10_X_25 ) , .A1( u0_u10_X_26 ) , .ZN( u0_u10_u4_n104 ) );
  AND2_X1 u0_u10_u4_U78 (.A1( u0_u10_X_30 ) , .A2( u0_u10_u4_n176 ) , .ZN( u0_u10_u4_n99 ) );
  AND2_X1 u0_u10_u4_U79 (.A1( u0_u10_X_26 ) , .ZN( u0_u10_u4_n101 ) , .A2( u0_u10_u4_n177 ) );
  INV_X1 u0_u10_u4_U8 (.A( u0_u10_u4_n113 ) , .ZN( u0_u10_u4_n185 ) );
  AND2_X1 u0_u10_u4_U80 (.A1( u0_u10_X_27 ) , .A2( u0_u10_X_30 ) , .ZN( u0_u10_u4_n103 ) );
  INV_X1 u0_u10_u4_U81 (.A( u0_u10_X_28 ) , .ZN( u0_u10_u4_n169 ) );
  INV_X1 u0_u10_u4_U82 (.A( u0_u10_X_29 ) , .ZN( u0_u10_u4_n168 ) );
  INV_X1 u0_u10_u4_U83 (.A( u0_u10_X_25 ) , .ZN( u0_u10_u4_n177 ) );
  INV_X1 u0_u10_u4_U84 (.A( u0_u10_X_27 ) , .ZN( u0_u10_u4_n176 ) );
  NAND4_X1 u0_u10_u4_U85 (.ZN( u0_out10_25 ) , .A4( u0_u10_u4_n139 ) , .A3( u0_u10_u4_n140 ) , .A2( u0_u10_u4_n141 ) , .A1( u0_u10_u4_n142 ) );
  OAI21_X1 u0_u10_u4_U86 (.A( u0_u10_u4_n128 ) , .B2( u0_u10_u4_n129 ) , .B1( u0_u10_u4_n130 ) , .ZN( u0_u10_u4_n142 ) );
  OAI21_X1 u0_u10_u4_U87 (.B2( u0_u10_u4_n131 ) , .ZN( u0_u10_u4_n141 ) , .A( u0_u10_u4_n175 ) , .B1( u0_u10_u4_n183 ) );
  NAND4_X1 u0_u10_u4_U88 (.ZN( u0_out10_14 ) , .A4( u0_u10_u4_n124 ) , .A3( u0_u10_u4_n125 ) , .A2( u0_u10_u4_n126 ) , .A1( u0_u10_u4_n127 ) );
  AOI22_X1 u0_u10_u4_U89 (.B2( u0_u10_u4_n117 ) , .ZN( u0_u10_u4_n126 ) , .A1( u0_u10_u4_n129 ) , .B1( u0_u10_u4_n152 ) , .A2( u0_u10_u4_n175 ) );
  NOR4_X1 u0_u10_u4_U9 (.A4( u0_u10_u4_n106 ) , .A3( u0_u10_u4_n107 ) , .A2( u0_u10_u4_n108 ) , .A1( u0_u10_u4_n109 ) , .ZN( u0_u10_u4_n110 ) );
  AOI22_X1 u0_u10_u4_U90 (.ZN( u0_u10_u4_n125 ) , .B2( u0_u10_u4_n131 ) , .A2( u0_u10_u4_n132 ) , .B1( u0_u10_u4_n138 ) , .A1( u0_u10_u4_n178 ) );
  NAND4_X1 u0_u10_u4_U91 (.ZN( u0_out10_8 ) , .A4( u0_u10_u4_n110 ) , .A3( u0_u10_u4_n111 ) , .A2( u0_u10_u4_n112 ) , .A1( u0_u10_u4_n186 ) );
  NAND2_X1 u0_u10_u4_U92 (.ZN( u0_u10_u4_n112 ) , .A2( u0_u10_u4_n130 ) , .A1( u0_u10_u4_n150 ) );
  AOI22_X1 u0_u10_u4_U93 (.ZN( u0_u10_u4_n111 ) , .B2( u0_u10_u4_n132 ) , .A1( u0_u10_u4_n152 ) , .B1( u0_u10_u4_n178 ) , .A2( u0_u10_u4_n97 ) );
  AOI22_X1 u0_u10_u4_U94 (.B2( u0_u10_u4_n149 ) , .B1( u0_u10_u4_n150 ) , .A2( u0_u10_u4_n151 ) , .A1( u0_u10_u4_n152 ) , .ZN( u0_u10_u4_n167 ) );
  NOR4_X1 u0_u10_u4_U95 (.A4( u0_u10_u4_n162 ) , .A3( u0_u10_u4_n163 ) , .A2( u0_u10_u4_n164 ) , .A1( u0_u10_u4_n165 ) , .ZN( u0_u10_u4_n166 ) );
  NAND3_X1 u0_u10_u4_U96 (.ZN( u0_out10_3 ) , .A3( u0_u10_u4_n166 ) , .A1( u0_u10_u4_n167 ) , .A2( u0_u10_u4_n186 ) );
  NAND3_X1 u0_u10_u4_U97 (.A3( u0_u10_u4_n146 ) , .A2( u0_u10_u4_n147 ) , .A1( u0_u10_u4_n148 ) , .ZN( u0_u10_u4_n149 ) );
  NAND3_X1 u0_u10_u4_U98 (.A3( u0_u10_u4_n143 ) , .A2( u0_u10_u4_n144 ) , .A1( u0_u10_u4_n145 ) , .ZN( u0_u10_u4_n151 ) );
  NAND3_X1 u0_u10_u4_U99 (.A3( u0_u10_u4_n121 ) , .ZN( u0_u10_u4_n122 ) , .A2( u0_u10_u4_n144 ) , .A1( u0_u10_u4_n154 ) );
  XOR2_X1 u0_u12_U26 (.B( u0_K13_30 ) , .A( u0_R11_21 ) , .Z( u0_u12_X_30 ) );
  XOR2_X1 u0_u12_U28 (.B( u0_K13_29 ) , .A( u0_R11_20 ) , .Z( u0_u12_X_29 ) );
  XOR2_X1 u0_u12_U29 (.B( u0_K13_28 ) , .A( u0_R11_19 ) , .Z( u0_u12_X_28 ) );
  XOR2_X1 u0_u12_U30 (.B( u0_K13_27 ) , .A( u0_R11_18 ) , .Z( u0_u12_X_27 ) );
  XOR2_X1 u0_u12_U31 (.B( u0_K13_26 ) , .A( u0_R11_17 ) , .Z( u0_u12_X_26 ) );
  XOR2_X1 u0_u12_U32 (.B( u0_K13_25 ) , .A( u0_R11_16 ) , .Z( u0_u12_X_25 ) );
  OAI22_X1 u0_u12_u4_U10 (.B2( u0_u12_u4_n135 ) , .ZN( u0_u12_u4_n137 ) , .B1( u0_u12_u4_n153 ) , .A1( u0_u12_u4_n155 ) , .A2( u0_u12_u4_n171 ) );
  AND3_X1 u0_u12_u4_U11 (.A2( u0_u12_u4_n134 ) , .ZN( u0_u12_u4_n135 ) , .A3( u0_u12_u4_n145 ) , .A1( u0_u12_u4_n157 ) );
  NAND2_X1 u0_u12_u4_U12 (.ZN( u0_u12_u4_n132 ) , .A2( u0_u12_u4_n170 ) , .A1( u0_u12_u4_n173 ) );
  AOI21_X1 u0_u12_u4_U13 (.B2( u0_u12_u4_n160 ) , .B1( u0_u12_u4_n161 ) , .ZN( u0_u12_u4_n162 ) , .A( u0_u12_u4_n170 ) );
  AOI21_X1 u0_u12_u4_U14 (.ZN( u0_u12_u4_n107 ) , .B2( u0_u12_u4_n143 ) , .A( u0_u12_u4_n174 ) , .B1( u0_u12_u4_n184 ) );
  AOI21_X1 u0_u12_u4_U15 (.B2( u0_u12_u4_n158 ) , .B1( u0_u12_u4_n159 ) , .ZN( u0_u12_u4_n163 ) , .A( u0_u12_u4_n174 ) );
  AOI21_X1 u0_u12_u4_U16 (.A( u0_u12_u4_n153 ) , .B2( u0_u12_u4_n154 ) , .B1( u0_u12_u4_n155 ) , .ZN( u0_u12_u4_n165 ) );
  AOI21_X1 u0_u12_u4_U17 (.A( u0_u12_u4_n156 ) , .B2( u0_u12_u4_n157 ) , .ZN( u0_u12_u4_n164 ) , .B1( u0_u12_u4_n184 ) );
  INV_X1 u0_u12_u4_U18 (.A( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n170 ) );
  AND2_X1 u0_u12_u4_U19 (.A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n155 ) , .A1( u0_u12_u4_n160 ) );
  INV_X1 u0_u12_u4_U20 (.A( u0_u12_u4_n156 ) , .ZN( u0_u12_u4_n175 ) );
  NAND2_X1 u0_u12_u4_U21 (.A2( u0_u12_u4_n118 ) , .ZN( u0_u12_u4_n131 ) , .A1( u0_u12_u4_n147 ) );
  NAND2_X1 u0_u12_u4_U22 (.A1( u0_u12_u4_n119 ) , .A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n130 ) );
  NAND2_X1 u0_u12_u4_U23 (.ZN( u0_u12_u4_n117 ) , .A2( u0_u12_u4_n118 ) , .A1( u0_u12_u4_n148 ) );
  NAND2_X1 u0_u12_u4_U24 (.ZN( u0_u12_u4_n129 ) , .A1( u0_u12_u4_n134 ) , .A2( u0_u12_u4_n148 ) );
  AND3_X1 u0_u12_u4_U25 (.A1( u0_u12_u4_n119 ) , .A2( u0_u12_u4_n143 ) , .A3( u0_u12_u4_n154 ) , .ZN( u0_u12_u4_n161 ) );
  AND2_X1 u0_u12_u4_U26 (.A1( u0_u12_u4_n145 ) , .A2( u0_u12_u4_n147 ) , .ZN( u0_u12_u4_n159 ) );
  OR3_X1 u0_u12_u4_U27 (.A3( u0_u12_u4_n114 ) , .A2( u0_u12_u4_n115 ) , .A1( u0_u12_u4_n116 ) , .ZN( u0_u12_u4_n136 ) );
  AOI21_X1 u0_u12_u4_U28 (.A( u0_u12_u4_n113 ) , .ZN( u0_u12_u4_n116 ) , .B2( u0_u12_u4_n173 ) , .B1( u0_u12_u4_n174 ) );
  AOI21_X1 u0_u12_u4_U29 (.ZN( u0_u12_u4_n115 ) , .B2( u0_u12_u4_n145 ) , .B1( u0_u12_u4_n146 ) , .A( u0_u12_u4_n156 ) );
  NOR2_X1 u0_u12_u4_U3 (.ZN( u0_u12_u4_n121 ) , .A1( u0_u12_u4_n181 ) , .A2( u0_u12_u4_n182 ) );
  OAI22_X1 u0_u12_u4_U30 (.ZN( u0_u12_u4_n114 ) , .A2( u0_u12_u4_n121 ) , .B1( u0_u12_u4_n160 ) , .B2( u0_u12_u4_n170 ) , .A1( u0_u12_u4_n171 ) );
  INV_X1 u0_u12_u4_U31 (.A( u0_u12_u4_n158 ) , .ZN( u0_u12_u4_n182 ) );
  INV_X1 u0_u12_u4_U32 (.ZN( u0_u12_u4_n181 ) , .A( u0_u12_u4_n96 ) );
  INV_X1 u0_u12_u4_U33 (.A( u0_u12_u4_n144 ) , .ZN( u0_u12_u4_n179 ) );
  INV_X1 u0_u12_u4_U34 (.A( u0_u12_u4_n157 ) , .ZN( u0_u12_u4_n178 ) );
  NAND2_X1 u0_u12_u4_U35 (.A2( u0_u12_u4_n154 ) , .A1( u0_u12_u4_n96 ) , .ZN( u0_u12_u4_n97 ) );
  INV_X1 u0_u12_u4_U36 (.ZN( u0_u12_u4_n186 ) , .A( u0_u12_u4_n95 ) );
  OAI221_X1 u0_u12_u4_U37 (.C1( u0_u12_u4_n134 ) , .B1( u0_u12_u4_n158 ) , .B2( u0_u12_u4_n171 ) , .C2( u0_u12_u4_n173 ) , .A( u0_u12_u4_n94 ) , .ZN( u0_u12_u4_n95 ) );
  AOI222_X1 u0_u12_u4_U38 (.B2( u0_u12_u4_n132 ) , .A1( u0_u12_u4_n138 ) , .C2( u0_u12_u4_n175 ) , .A2( u0_u12_u4_n179 ) , .C1( u0_u12_u4_n181 ) , .B1( u0_u12_u4_n185 ) , .ZN( u0_u12_u4_n94 ) );
  INV_X1 u0_u12_u4_U39 (.A( u0_u12_u4_n113 ) , .ZN( u0_u12_u4_n185 ) );
  INV_X1 u0_u12_u4_U4 (.A( u0_u12_u4_n117 ) , .ZN( u0_u12_u4_n184 ) );
  INV_X1 u0_u12_u4_U40 (.A( u0_u12_u4_n143 ) , .ZN( u0_u12_u4_n183 ) );
  NOR2_X1 u0_u12_u4_U41 (.ZN( u0_u12_u4_n138 ) , .A1( u0_u12_u4_n168 ) , .A2( u0_u12_u4_n169 ) );
  NOR2_X1 u0_u12_u4_U42 (.A1( u0_u12_u4_n150 ) , .A2( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n153 ) );
  NOR2_X1 u0_u12_u4_U43 (.A2( u0_u12_u4_n128 ) , .A1( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n156 ) );
  AOI22_X1 u0_u12_u4_U44 (.B2( u0_u12_u4_n122 ) , .A1( u0_u12_u4_n123 ) , .ZN( u0_u12_u4_n124 ) , .B1( u0_u12_u4_n128 ) , .A2( u0_u12_u4_n172 ) );
  INV_X1 u0_u12_u4_U45 (.A( u0_u12_u4_n153 ) , .ZN( u0_u12_u4_n172 ) );
  NAND2_X1 u0_u12_u4_U46 (.A2( u0_u12_u4_n120 ) , .ZN( u0_u12_u4_n123 ) , .A1( u0_u12_u4_n161 ) );
  AOI22_X1 u0_u12_u4_U47 (.B2( u0_u12_u4_n132 ) , .A2( u0_u12_u4_n133 ) , .ZN( u0_u12_u4_n140 ) , .A1( u0_u12_u4_n150 ) , .B1( u0_u12_u4_n179 ) );
  NAND2_X1 u0_u12_u4_U48 (.ZN( u0_u12_u4_n133 ) , .A2( u0_u12_u4_n146 ) , .A1( u0_u12_u4_n154 ) );
  NAND2_X1 u0_u12_u4_U49 (.A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n154 ) , .A2( u0_u12_u4_n98 ) );
  NOR4_X1 u0_u12_u4_U5 (.A4( u0_u12_u4_n106 ) , .A3( u0_u12_u4_n107 ) , .A2( u0_u12_u4_n108 ) , .A1( u0_u12_u4_n109 ) , .ZN( u0_u12_u4_n110 ) );
  NAND2_X1 u0_u12_u4_U50 (.A1( u0_u12_u4_n101 ) , .ZN( u0_u12_u4_n158 ) , .A2( u0_u12_u4_n99 ) );
  AOI21_X1 u0_u12_u4_U51 (.ZN( u0_u12_u4_n127 ) , .A( u0_u12_u4_n136 ) , .B2( u0_u12_u4_n150 ) , .B1( u0_u12_u4_n180 ) );
  INV_X1 u0_u12_u4_U52 (.A( u0_u12_u4_n160 ) , .ZN( u0_u12_u4_n180 ) );
  NAND2_X1 u0_u12_u4_U53 (.A2( u0_u12_u4_n104 ) , .A1( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n146 ) );
  NAND2_X1 u0_u12_u4_U54 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n160 ) );
  NAND2_X1 u0_u12_u4_U55 (.ZN( u0_u12_u4_n134 ) , .A1( u0_u12_u4_n98 ) , .A2( u0_u12_u4_n99 ) );
  NAND2_X1 u0_u12_u4_U56 (.A1( u0_u12_u4_n103 ) , .A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n143 ) );
  NAND2_X1 u0_u12_u4_U57 (.A2( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n145 ) , .A1( u0_u12_u4_n98 ) );
  NAND2_X1 u0_u12_u4_U58 (.A1( u0_u12_u4_n100 ) , .A2( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n120 ) );
  NAND2_X1 u0_u12_u4_U59 (.A1( u0_u12_u4_n102 ) , .A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n148 ) );
  AOI21_X1 u0_u12_u4_U6 (.ZN( u0_u12_u4_n106 ) , .B2( u0_u12_u4_n146 ) , .B1( u0_u12_u4_n158 ) , .A( u0_u12_u4_n170 ) );
  NAND2_X1 u0_u12_u4_U60 (.A2( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n157 ) );
  INV_X1 u0_u12_u4_U61 (.A( u0_u12_u4_n150 ) , .ZN( u0_u12_u4_n173 ) );
  INV_X1 u0_u12_u4_U62 (.A( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n171 ) );
  NAND2_X1 u0_u12_u4_U63 (.A1( u0_u12_u4_n100 ) , .ZN( u0_u12_u4_n118 ) , .A2( u0_u12_u4_n99 ) );
  NAND2_X1 u0_u12_u4_U64 (.A2( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n144 ) );
  NAND2_X1 u0_u12_u4_U65 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n105 ) , .ZN( u0_u12_u4_n96 ) );
  INV_X1 u0_u12_u4_U66 (.A( u0_u12_u4_n128 ) , .ZN( u0_u12_u4_n174 ) );
  NAND2_X1 u0_u12_u4_U67 (.A2( u0_u12_u4_n102 ) , .ZN( u0_u12_u4_n119 ) , .A1( u0_u12_u4_n98 ) );
  NAND2_X1 u0_u12_u4_U68 (.A2( u0_u12_u4_n101 ) , .A1( u0_u12_u4_n103 ) , .ZN( u0_u12_u4_n147 ) );
  NAND2_X1 u0_u12_u4_U69 (.A2( u0_u12_u4_n104 ) , .ZN( u0_u12_u4_n113 ) , .A1( u0_u12_u4_n99 ) );
  AOI21_X1 u0_u12_u4_U7 (.ZN( u0_u12_u4_n108 ) , .B2( u0_u12_u4_n134 ) , .B1( u0_u12_u4_n155 ) , .A( u0_u12_u4_n156 ) );
  NOR2_X1 u0_u12_u4_U70 (.A2( u0_u12_X_28 ) , .ZN( u0_u12_u4_n150 ) , .A1( u0_u12_u4_n168 ) );
  NOR2_X1 u0_u12_u4_U71 (.A2( u0_u12_X_29 ) , .ZN( u0_u12_u4_n152 ) , .A1( u0_u12_u4_n169 ) );
  NOR2_X1 u0_u12_u4_U72 (.A2( u0_u12_X_30 ) , .ZN( u0_u12_u4_n105 ) , .A1( u0_u12_u4_n176 ) );
  NOR2_X1 u0_u12_u4_U73 (.A2( u0_u12_X_26 ) , .ZN( u0_u12_u4_n100 ) , .A1( u0_u12_u4_n177 ) );
  NOR2_X1 u0_u12_u4_U74 (.A2( u0_u12_X_28 ) , .A1( u0_u12_X_29 ) , .ZN( u0_u12_u4_n128 ) );
  NOR2_X1 u0_u12_u4_U75 (.A2( u0_u12_X_27 ) , .A1( u0_u12_X_30 ) , .ZN( u0_u12_u4_n102 ) );
  NOR2_X1 u0_u12_u4_U76 (.A2( u0_u12_X_25 ) , .A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n98 ) );
  AND2_X1 u0_u12_u4_U77 (.A2( u0_u12_X_25 ) , .A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n104 ) );
  AND2_X1 u0_u12_u4_U78 (.A1( u0_u12_X_30 ) , .A2( u0_u12_u4_n176 ) , .ZN( u0_u12_u4_n99 ) );
  AND2_X1 u0_u12_u4_U79 (.A1( u0_u12_X_26 ) , .ZN( u0_u12_u4_n101 ) , .A2( u0_u12_u4_n177 ) );
  AOI21_X1 u0_u12_u4_U8 (.ZN( u0_u12_u4_n109 ) , .A( u0_u12_u4_n153 ) , .B1( u0_u12_u4_n159 ) , .B2( u0_u12_u4_n184 ) );
  AND2_X1 u0_u12_u4_U80 (.A1( u0_u12_X_27 ) , .A2( u0_u12_X_30 ) , .ZN( u0_u12_u4_n103 ) );
  INV_X1 u0_u12_u4_U81 (.A( u0_u12_X_28 ) , .ZN( u0_u12_u4_n169 ) );
  INV_X1 u0_u12_u4_U82 (.A( u0_u12_X_29 ) , .ZN( u0_u12_u4_n168 ) );
  INV_X1 u0_u12_u4_U83 (.A( u0_u12_X_25 ) , .ZN( u0_u12_u4_n177 ) );
  INV_X1 u0_u12_u4_U84 (.A( u0_u12_X_27 ) , .ZN( u0_u12_u4_n176 ) );
  NAND4_X1 u0_u12_u4_U85 (.ZN( u0_out12_25 ) , .A4( u0_u12_u4_n139 ) , .A3( u0_u12_u4_n140 ) , .A2( u0_u12_u4_n141 ) , .A1( u0_u12_u4_n142 ) );
  OAI21_X1 u0_u12_u4_U86 (.A( u0_u12_u4_n128 ) , .B2( u0_u12_u4_n129 ) , .B1( u0_u12_u4_n130 ) , .ZN( u0_u12_u4_n142 ) );
  OAI21_X1 u0_u12_u4_U87 (.B2( u0_u12_u4_n131 ) , .ZN( u0_u12_u4_n141 ) , .A( u0_u12_u4_n175 ) , .B1( u0_u12_u4_n183 ) );
  NAND4_X1 u0_u12_u4_U88 (.ZN( u0_out12_14 ) , .A4( u0_u12_u4_n124 ) , .A3( u0_u12_u4_n125 ) , .A2( u0_u12_u4_n126 ) , .A1( u0_u12_u4_n127 ) );
  AOI22_X1 u0_u12_u4_U89 (.B2( u0_u12_u4_n117 ) , .ZN( u0_u12_u4_n126 ) , .A1( u0_u12_u4_n129 ) , .B1( u0_u12_u4_n152 ) , .A2( u0_u12_u4_n175 ) );
  AOI211_X1 u0_u12_u4_U9 (.B( u0_u12_u4_n136 ) , .A( u0_u12_u4_n137 ) , .C2( u0_u12_u4_n138 ) , .ZN( u0_u12_u4_n139 ) , .C1( u0_u12_u4_n182 ) );
  AOI22_X1 u0_u12_u4_U90 (.ZN( u0_u12_u4_n125 ) , .B2( u0_u12_u4_n131 ) , .A2( u0_u12_u4_n132 ) , .B1( u0_u12_u4_n138 ) , .A1( u0_u12_u4_n178 ) );
  NAND4_X1 u0_u12_u4_U91 (.ZN( u0_out12_8 ) , .A4( u0_u12_u4_n110 ) , .A3( u0_u12_u4_n111 ) , .A2( u0_u12_u4_n112 ) , .A1( u0_u12_u4_n186 ) );
  NAND2_X1 u0_u12_u4_U92 (.ZN( u0_u12_u4_n112 ) , .A2( u0_u12_u4_n130 ) , .A1( u0_u12_u4_n150 ) );
  AOI22_X1 u0_u12_u4_U93 (.ZN( u0_u12_u4_n111 ) , .B2( u0_u12_u4_n132 ) , .A1( u0_u12_u4_n152 ) , .B1( u0_u12_u4_n178 ) , .A2( u0_u12_u4_n97 ) );
  AOI22_X1 u0_u12_u4_U94 (.B2( u0_u12_u4_n149 ) , .B1( u0_u12_u4_n150 ) , .A2( u0_u12_u4_n151 ) , .A1( u0_u12_u4_n152 ) , .ZN( u0_u12_u4_n167 ) );
  NOR4_X1 u0_u12_u4_U95 (.A4( u0_u12_u4_n162 ) , .A3( u0_u12_u4_n163 ) , .A2( u0_u12_u4_n164 ) , .A1( u0_u12_u4_n165 ) , .ZN( u0_u12_u4_n166 ) );
  NAND3_X1 u0_u12_u4_U96 (.ZN( u0_out12_3 ) , .A3( u0_u12_u4_n166 ) , .A1( u0_u12_u4_n167 ) , .A2( u0_u12_u4_n186 ) );
  NAND3_X1 u0_u12_u4_U97 (.A3( u0_u12_u4_n146 ) , .A2( u0_u12_u4_n147 ) , .A1( u0_u12_u4_n148 ) , .ZN( u0_u12_u4_n149 ) );
  NAND3_X1 u0_u12_u4_U98 (.A3( u0_u12_u4_n143 ) , .A2( u0_u12_u4_n144 ) , .A1( u0_u12_u4_n145 ) , .ZN( u0_u12_u4_n151 ) );
  NAND3_X1 u0_u12_u4_U99 (.A3( u0_u12_u4_n121 ) , .ZN( u0_u12_u4_n122 ) , .A2( u0_u12_u4_n144 ) , .A1( u0_u12_u4_n154 ) );
  XOR2_X1 u0_u14_U1 (.B( u0_K15_9 ) , .A( u0_R13_6 ) , .Z( u0_u14_X_9 ) );
  XOR2_X1 u0_u14_U2 (.B( u0_K15_8 ) , .A( u0_R13_5 ) , .Z( u0_u14_X_8 ) );
  XOR2_X1 u0_u14_U20 (.B( u0_K15_36 ) , .A( u0_R13_25 ) , .Z( u0_u14_X_36 ) );
  XOR2_X1 u0_u14_U21 (.B( u0_K15_35 ) , .A( u0_R13_24 ) , .Z( u0_u14_X_35 ) );
  XOR2_X1 u0_u14_U22 (.B( u0_K15_34 ) , .A( u0_R13_23 ) , .Z( u0_u14_X_34 ) );
  XOR2_X1 u0_u14_U23 (.B( u0_K15_33 ) , .A( u0_R13_22 ) , .Z( u0_u14_X_33 ) );
  XOR2_X1 u0_u14_U24 (.B( u0_K15_32 ) , .A( u0_R13_21 ) , .Z( u0_u14_X_32 ) );
  XOR2_X1 u0_u14_U25 (.B( u0_K15_31 ) , .A( u0_R13_20 ) , .Z( u0_u14_X_31 ) );
  XOR2_X1 u0_u14_U3 (.B( u0_K15_7 ) , .A( u0_R13_4 ) , .Z( u0_u14_X_7 ) );
  XOR2_X1 u0_u14_U33 (.B( u0_K15_24 ) , .A( u0_R13_17 ) , .Z( u0_u14_X_24 ) );
  XOR2_X1 u0_u14_U34 (.B( u0_K15_23 ) , .A( u0_R13_16 ) , .Z( u0_u14_X_23 ) );
  XOR2_X1 u0_u14_U35 (.B( u0_K15_22 ) , .A( u0_R13_15 ) , .Z( u0_u14_X_22 ) );
  XOR2_X1 u0_u14_U36 (.B( u0_K15_21 ) , .A( u0_R13_14 ) , .Z( u0_u14_X_21 ) );
  XOR2_X1 u0_u14_U37 (.B( u0_K15_20 ) , .A( u0_R13_13 ) , .Z( u0_u14_X_20 ) );
  XOR2_X1 u0_u14_U39 (.B( u0_K15_19 ) , .A( u0_R13_12 ) , .Z( u0_u14_X_19 ) );
  XOR2_X1 u0_u14_U40 (.B( u0_K15_18 ) , .A( u0_R13_13 ) , .Z( u0_u14_X_18 ) );
  XOR2_X1 u0_u14_U41 (.B( u0_K15_17 ) , .A( u0_R13_12 ) , .Z( u0_u14_X_17 ) );
  XOR2_X1 u0_u14_U42 (.B( u0_K15_16 ) , .A( u0_R13_11 ) , .Z( u0_u14_X_16 ) );
  XOR2_X1 u0_u14_U43 (.B( u0_K15_15 ) , .A( u0_R13_10 ) , .Z( u0_u14_X_15 ) );
  XOR2_X1 u0_u14_U44 (.B( u0_K15_14 ) , .A( u0_R13_9 ) , .Z( u0_u14_X_14 ) );
  XOR2_X1 u0_u14_U45 (.B( u0_K15_13 ) , .A( u0_R13_8 ) , .Z( u0_u14_X_13 ) );
  XOR2_X1 u0_u14_U46 (.B( u0_K15_12 ) , .A( u0_R13_9 ) , .Z( u0_u14_X_12 ) );
  XOR2_X1 u0_u14_U47 (.B( u0_K15_11 ) , .A( u0_R13_8 ) , .Z( u0_u14_X_11 ) );
  XOR2_X1 u0_u14_U48 (.B( u0_K15_10 ) , .A( u0_R13_7 ) , .Z( u0_u14_X_10 ) );
  AOI21_X1 u0_u14_u1_U10 (.ZN( u0_u14_u1_n106 ) , .A( u0_u14_u1_n112 ) , .B1( u0_u14_u1_n154 ) , .B2( u0_u14_u1_n156 ) );
  NAND3_X1 u0_u14_u1_U100 (.ZN( u0_u14_u1_n113 ) , .A1( u0_u14_u1_n120 ) , .A3( u0_u14_u1_n133 ) , .A2( u0_u14_u1_n155 ) );
  INV_X1 u0_u14_u1_U11 (.A( u0_u14_u1_n101 ) , .ZN( u0_u14_u1_n184 ) );
  AOI21_X1 u0_u14_u1_U12 (.ZN( u0_u14_u1_n107 ) , .B1( u0_u14_u1_n134 ) , .B2( u0_u14_u1_n149 ) , .A( u0_u14_u1_n174 ) );
  NAND2_X1 u0_u14_u1_U13 (.ZN( u0_u14_u1_n140 ) , .A2( u0_u14_u1_n150 ) , .A1( u0_u14_u1_n155 ) );
  NAND2_X1 u0_u14_u1_U14 (.A1( u0_u14_u1_n131 ) , .ZN( u0_u14_u1_n147 ) , .A2( u0_u14_u1_n153 ) );
  AOI22_X1 u0_u14_u1_U15 (.B2( u0_u14_u1_n136 ) , .A2( u0_u14_u1_n137 ) , .ZN( u0_u14_u1_n143 ) , .A1( u0_u14_u1_n171 ) , .B1( u0_u14_u1_n173 ) );
  INV_X1 u0_u14_u1_U16 (.A( u0_u14_u1_n147 ) , .ZN( u0_u14_u1_n181 ) );
  INV_X1 u0_u14_u1_U17 (.A( u0_u14_u1_n139 ) , .ZN( u0_u14_u1_n174 ) );
  INV_X1 u0_u14_u1_U18 (.A( u0_u14_u1_n112 ) , .ZN( u0_u14_u1_n171 ) );
  NAND2_X1 u0_u14_u1_U19 (.ZN( u0_u14_u1_n141 ) , .A1( u0_u14_u1_n153 ) , .A2( u0_u14_u1_n156 ) );
  AND2_X1 u0_u14_u1_U20 (.A1( u0_u14_u1_n123 ) , .ZN( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n161 ) );
  NAND2_X1 u0_u14_u1_U21 (.A2( u0_u14_u1_n115 ) , .A1( u0_u14_u1_n116 ) , .ZN( u0_u14_u1_n148 ) );
  NAND2_X1 u0_u14_u1_U22 (.A2( u0_u14_u1_n133 ) , .A1( u0_u14_u1_n135 ) , .ZN( u0_u14_u1_n159 ) );
  NAND2_X1 u0_u14_u1_U23 (.A2( u0_u14_u1_n115 ) , .A1( u0_u14_u1_n120 ) , .ZN( u0_u14_u1_n132 ) );
  INV_X1 u0_u14_u1_U24 (.A( u0_u14_u1_n154 ) , .ZN( u0_u14_u1_n178 ) );
  AOI22_X1 u0_u14_u1_U25 (.B2( u0_u14_u1_n113 ) , .A2( u0_u14_u1_n114 ) , .ZN( u0_u14_u1_n125 ) , .A1( u0_u14_u1_n171 ) , .B1( u0_u14_u1_n173 ) );
  NAND2_X1 u0_u14_u1_U26 (.ZN( u0_u14_u1_n114 ) , .A1( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n156 ) );
  INV_X1 u0_u14_u1_U27 (.A( u0_u14_u1_n151 ) , .ZN( u0_u14_u1_n183 ) );
  AND2_X1 u0_u14_u1_U28 (.A1( u0_u14_u1_n129 ) , .A2( u0_u14_u1_n133 ) , .ZN( u0_u14_u1_n149 ) );
  INV_X1 u0_u14_u1_U29 (.A( u0_u14_u1_n131 ) , .ZN( u0_u14_u1_n180 ) );
  INV_X1 u0_u14_u1_U3 (.A( u0_u14_u1_n159 ) , .ZN( u0_u14_u1_n182 ) );
  AOI221_X1 u0_u14_u1_U30 (.B1( u0_u14_u1_n140 ) , .ZN( u0_u14_u1_n167 ) , .B2( u0_u14_u1_n172 ) , .C2( u0_u14_u1_n175 ) , .C1( u0_u14_u1_n178 ) , .A( u0_u14_u1_n188 ) );
  INV_X1 u0_u14_u1_U31 (.ZN( u0_u14_u1_n188 ) , .A( u0_u14_u1_n97 ) );
  AOI211_X1 u0_u14_u1_U32 (.A( u0_u14_u1_n118 ) , .C1( u0_u14_u1_n132 ) , .C2( u0_u14_u1_n139 ) , .B( u0_u14_u1_n96 ) , .ZN( u0_u14_u1_n97 ) );
  AOI21_X1 u0_u14_u1_U33 (.B2( u0_u14_u1_n121 ) , .B1( u0_u14_u1_n135 ) , .A( u0_u14_u1_n152 ) , .ZN( u0_u14_u1_n96 ) );
  OAI221_X1 u0_u14_u1_U34 (.A( u0_u14_u1_n119 ) , .C2( u0_u14_u1_n129 ) , .ZN( u0_u14_u1_n138 ) , .B2( u0_u14_u1_n152 ) , .C1( u0_u14_u1_n174 ) , .B1( u0_u14_u1_n187 ) );
  INV_X1 u0_u14_u1_U35 (.A( u0_u14_u1_n148 ) , .ZN( u0_u14_u1_n187 ) );
  AOI211_X1 u0_u14_u1_U36 (.B( u0_u14_u1_n117 ) , .A( u0_u14_u1_n118 ) , .ZN( u0_u14_u1_n119 ) , .C2( u0_u14_u1_n146 ) , .C1( u0_u14_u1_n159 ) );
  NOR2_X1 u0_u14_u1_U37 (.A1( u0_u14_u1_n168 ) , .A2( u0_u14_u1_n176 ) , .ZN( u0_u14_u1_n98 ) );
  AOI211_X1 u0_u14_u1_U38 (.B( u0_u14_u1_n162 ) , .A( u0_u14_u1_n163 ) , .C2( u0_u14_u1_n164 ) , .ZN( u0_u14_u1_n165 ) , .C1( u0_u14_u1_n171 ) );
  AOI21_X1 u0_u14_u1_U39 (.A( u0_u14_u1_n160 ) , .B2( u0_u14_u1_n161 ) , .ZN( u0_u14_u1_n162 ) , .B1( u0_u14_u1_n182 ) );
  AOI221_X1 u0_u14_u1_U4 (.A( u0_u14_u1_n138 ) , .C2( u0_u14_u1_n139 ) , .C1( u0_u14_u1_n140 ) , .B2( u0_u14_u1_n141 ) , .ZN( u0_u14_u1_n142 ) , .B1( u0_u14_u1_n175 ) );
  OR2_X1 u0_u14_u1_U40 (.A2( u0_u14_u1_n157 ) , .A1( u0_u14_u1_n158 ) , .ZN( u0_u14_u1_n163 ) );
  OAI21_X1 u0_u14_u1_U41 (.B2( u0_u14_u1_n123 ) , .ZN( u0_u14_u1_n145 ) , .B1( u0_u14_u1_n160 ) , .A( u0_u14_u1_n185 ) );
  INV_X1 u0_u14_u1_U42 (.A( u0_u14_u1_n122 ) , .ZN( u0_u14_u1_n185 ) );
  AOI21_X1 u0_u14_u1_U43 (.B2( u0_u14_u1_n120 ) , .B1( u0_u14_u1_n121 ) , .ZN( u0_u14_u1_n122 ) , .A( u0_u14_u1_n128 ) );
  NAND2_X1 u0_u14_u1_U44 (.A1( u0_u14_u1_n128 ) , .ZN( u0_u14_u1_n146 ) , .A2( u0_u14_u1_n160 ) );
  NAND2_X1 u0_u14_u1_U45 (.A2( u0_u14_u1_n112 ) , .ZN( u0_u14_u1_n139 ) , .A1( u0_u14_u1_n152 ) );
  NAND2_X1 u0_u14_u1_U46 (.A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n156 ) , .A2( u0_u14_u1_n99 ) );
  NOR2_X1 u0_u14_u1_U47 (.ZN( u0_u14_u1_n117 ) , .A1( u0_u14_u1_n121 ) , .A2( u0_u14_u1_n160 ) );
  AOI21_X1 u0_u14_u1_U48 (.A( u0_u14_u1_n128 ) , .B2( u0_u14_u1_n129 ) , .ZN( u0_u14_u1_n130 ) , .B1( u0_u14_u1_n150 ) );
  NAND2_X1 u0_u14_u1_U49 (.ZN( u0_u14_u1_n112 ) , .A1( u0_u14_u1_n169 ) , .A2( u0_u14_u1_n170 ) );
  AOI211_X1 u0_u14_u1_U5 (.ZN( u0_u14_u1_n124 ) , .A( u0_u14_u1_n138 ) , .C2( u0_u14_u1_n139 ) , .B( u0_u14_u1_n145 ) , .C1( u0_u14_u1_n147 ) );
  NAND2_X1 u0_u14_u1_U50 (.ZN( u0_u14_u1_n129 ) , .A2( u0_u14_u1_n95 ) , .A1( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U51 (.A1( u0_u14_u1_n102 ) , .ZN( u0_u14_u1_n154 ) , .A2( u0_u14_u1_n99 ) );
  NAND2_X1 u0_u14_u1_U52 (.A2( u0_u14_u1_n100 ) , .ZN( u0_u14_u1_n135 ) , .A1( u0_u14_u1_n99 ) );
  AOI21_X1 u0_u14_u1_U53 (.A( u0_u14_u1_n152 ) , .B2( u0_u14_u1_n153 ) , .B1( u0_u14_u1_n154 ) , .ZN( u0_u14_u1_n158 ) );
  INV_X1 u0_u14_u1_U54 (.A( u0_u14_u1_n160 ) , .ZN( u0_u14_u1_n175 ) );
  NAND2_X1 u0_u14_u1_U55 (.A1( u0_u14_u1_n100 ) , .ZN( u0_u14_u1_n116 ) , .A2( u0_u14_u1_n95 ) );
  NAND2_X1 u0_u14_u1_U56 (.A1( u0_u14_u1_n102 ) , .ZN( u0_u14_u1_n131 ) , .A2( u0_u14_u1_n95 ) );
  NAND2_X1 u0_u14_u1_U57 (.A2( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n121 ) , .A1( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U58 (.A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n153 ) , .A2( u0_u14_u1_n98 ) );
  NAND2_X1 u0_u14_u1_U59 (.A2( u0_u14_u1_n104 ) , .A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n133 ) );
  NOR2_X1 u0_u14_u1_U6 (.A1( u0_u14_u1_n112 ) , .A2( u0_u14_u1_n116 ) , .ZN( u0_u14_u1_n118 ) );
  NAND2_X1 u0_u14_u1_U60 (.ZN( u0_u14_u1_n150 ) , .A2( u0_u14_u1_n98 ) , .A1( u0_u14_u1_n99 ) );
  NAND2_X1 u0_u14_u1_U61 (.A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n155 ) , .A2( u0_u14_u1_n95 ) );
  OAI21_X1 u0_u14_u1_U62 (.ZN( u0_u14_u1_n109 ) , .B1( u0_u14_u1_n129 ) , .B2( u0_u14_u1_n160 ) , .A( u0_u14_u1_n167 ) );
  NAND2_X1 u0_u14_u1_U63 (.A2( u0_u14_u1_n100 ) , .A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n120 ) );
  NAND2_X1 u0_u14_u1_U64 (.A1( u0_u14_u1_n102 ) , .A2( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n115 ) );
  NAND2_X1 u0_u14_u1_U65 (.A2( u0_u14_u1_n100 ) , .A1( u0_u14_u1_n104 ) , .ZN( u0_u14_u1_n151 ) );
  NAND2_X1 u0_u14_u1_U66 (.A2( u0_u14_u1_n103 ) , .A1( u0_u14_u1_n105 ) , .ZN( u0_u14_u1_n161 ) );
  INV_X1 u0_u14_u1_U67 (.A( u0_u14_u1_n152 ) , .ZN( u0_u14_u1_n173 ) );
  INV_X1 u0_u14_u1_U68 (.A( u0_u14_u1_n128 ) , .ZN( u0_u14_u1_n172 ) );
  NAND2_X1 u0_u14_u1_U69 (.A2( u0_u14_u1_n102 ) , .A1( u0_u14_u1_n103 ) , .ZN( u0_u14_u1_n123 ) );
  OAI21_X1 u0_u14_u1_U7 (.ZN( u0_u14_u1_n101 ) , .B1( u0_u14_u1_n141 ) , .A( u0_u14_u1_n146 ) , .B2( u0_u14_u1_n183 ) );
  NOR2_X1 u0_u14_u1_U70 (.A2( u0_u14_X_7 ) , .A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n95 ) );
  NOR2_X1 u0_u14_u1_U71 (.A1( u0_u14_X_12 ) , .A2( u0_u14_X_9 ) , .ZN( u0_u14_u1_n100 ) );
  NOR2_X1 u0_u14_u1_U72 (.A2( u0_u14_X_8 ) , .A1( u0_u14_u1_n177 ) , .ZN( u0_u14_u1_n99 ) );
  NOR2_X1 u0_u14_u1_U73 (.A2( u0_u14_X_12 ) , .ZN( u0_u14_u1_n102 ) , .A1( u0_u14_u1_n176 ) );
  NOR2_X1 u0_u14_u1_U74 (.A2( u0_u14_X_9 ) , .ZN( u0_u14_u1_n105 ) , .A1( u0_u14_u1_n168 ) );
  NAND2_X1 u0_u14_u1_U75 (.A1( u0_u14_X_10 ) , .ZN( u0_u14_u1_n160 ) , .A2( u0_u14_u1_n169 ) );
  NAND2_X1 u0_u14_u1_U76 (.A2( u0_u14_X_10 ) , .A1( u0_u14_X_11 ) , .ZN( u0_u14_u1_n152 ) );
  NAND2_X1 u0_u14_u1_U77 (.A1( u0_u14_X_11 ) , .ZN( u0_u14_u1_n128 ) , .A2( u0_u14_u1_n170 ) );
  AND2_X1 u0_u14_u1_U78 (.A2( u0_u14_X_7 ) , .A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n104 ) );
  AND2_X1 u0_u14_u1_U79 (.A1( u0_u14_X_8 ) , .ZN( u0_u14_u1_n103 ) , .A2( u0_u14_u1_n177 ) );
  AOI21_X1 u0_u14_u1_U8 (.B2( u0_u14_u1_n155 ) , .B1( u0_u14_u1_n156 ) , .ZN( u0_u14_u1_n157 ) , .A( u0_u14_u1_n174 ) );
  INV_X1 u0_u14_u1_U80 (.A( u0_u14_X_10 ) , .ZN( u0_u14_u1_n170 ) );
  INV_X1 u0_u14_u1_U81 (.A( u0_u14_X_9 ) , .ZN( u0_u14_u1_n176 ) );
  INV_X1 u0_u14_u1_U82 (.A( u0_u14_X_11 ) , .ZN( u0_u14_u1_n169 ) );
  INV_X1 u0_u14_u1_U83 (.A( u0_u14_X_12 ) , .ZN( u0_u14_u1_n168 ) );
  INV_X1 u0_u14_u1_U84 (.A( u0_u14_X_7 ) , .ZN( u0_u14_u1_n177 ) );
  NAND4_X1 u0_u14_u1_U85 (.ZN( u0_out14_28 ) , .A4( u0_u14_u1_n124 ) , .A3( u0_u14_u1_n125 ) , .A2( u0_u14_u1_n126 ) , .A1( u0_u14_u1_n127 ) );
  OAI21_X1 u0_u14_u1_U86 (.ZN( u0_u14_u1_n127 ) , .B2( u0_u14_u1_n139 ) , .B1( u0_u14_u1_n175 ) , .A( u0_u14_u1_n183 ) );
  OAI21_X1 u0_u14_u1_U87 (.ZN( u0_u14_u1_n126 ) , .B2( u0_u14_u1_n140 ) , .A( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n178 ) );
  NAND4_X1 u0_u14_u1_U88 (.ZN( u0_out14_18 ) , .A4( u0_u14_u1_n165 ) , .A3( u0_u14_u1_n166 ) , .A1( u0_u14_u1_n167 ) , .A2( u0_u14_u1_n186 ) );
  AOI22_X1 u0_u14_u1_U89 (.B2( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n147 ) , .A2( u0_u14_u1_n148 ) , .ZN( u0_u14_u1_n166 ) , .A1( u0_u14_u1_n172 ) );
  OR4_X1 u0_u14_u1_U9 (.A4( u0_u14_u1_n106 ) , .A3( u0_u14_u1_n107 ) , .ZN( u0_u14_u1_n108 ) , .A1( u0_u14_u1_n117 ) , .A2( u0_u14_u1_n184 ) );
  INV_X1 u0_u14_u1_U90 (.A( u0_u14_u1_n145 ) , .ZN( u0_u14_u1_n186 ) );
  NAND4_X1 u0_u14_u1_U91 (.ZN( u0_out14_2 ) , .A4( u0_u14_u1_n142 ) , .A3( u0_u14_u1_n143 ) , .A2( u0_u14_u1_n144 ) , .A1( u0_u14_u1_n179 ) );
  OAI21_X1 u0_u14_u1_U92 (.B2( u0_u14_u1_n132 ) , .ZN( u0_u14_u1_n144 ) , .A( u0_u14_u1_n146 ) , .B1( u0_u14_u1_n180 ) );
  INV_X1 u0_u14_u1_U93 (.A( u0_u14_u1_n130 ) , .ZN( u0_u14_u1_n179 ) );
  OR4_X1 u0_u14_u1_U94 (.ZN( u0_out14_13 ) , .A4( u0_u14_u1_n108 ) , .A3( u0_u14_u1_n109 ) , .A2( u0_u14_u1_n110 ) , .A1( u0_u14_u1_n111 ) );
  AOI21_X1 u0_u14_u1_U95 (.ZN( u0_u14_u1_n111 ) , .A( u0_u14_u1_n128 ) , .B2( u0_u14_u1_n131 ) , .B1( u0_u14_u1_n135 ) );
  AOI21_X1 u0_u14_u1_U96 (.ZN( u0_u14_u1_n110 ) , .A( u0_u14_u1_n116 ) , .B1( u0_u14_u1_n152 ) , .B2( u0_u14_u1_n160 ) );
  NAND3_X1 u0_u14_u1_U97 (.A3( u0_u14_u1_n149 ) , .A2( u0_u14_u1_n150 ) , .A1( u0_u14_u1_n151 ) , .ZN( u0_u14_u1_n164 ) );
  NAND3_X1 u0_u14_u1_U98 (.A3( u0_u14_u1_n134 ) , .A2( u0_u14_u1_n135 ) , .ZN( u0_u14_u1_n136 ) , .A1( u0_u14_u1_n151 ) );
  NAND3_X1 u0_u14_u1_U99 (.A1( u0_u14_u1_n133 ) , .ZN( u0_u14_u1_n137 ) , .A2( u0_u14_u1_n154 ) , .A3( u0_u14_u1_n181 ) );
  OAI22_X1 u0_u14_u2_U10 (.ZN( u0_u14_u2_n109 ) , .A2( u0_u14_u2_n113 ) , .B2( u0_u14_u2_n133 ) , .B1( u0_u14_u2_n167 ) , .A1( u0_u14_u2_n168 ) );
  NAND3_X1 u0_u14_u2_U100 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n98 ) );
  OAI22_X1 u0_u14_u2_U11 (.B1( u0_u14_u2_n151 ) , .A2( u0_u14_u2_n152 ) , .A1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n160 ) , .B2( u0_u14_u2_n168 ) );
  NOR3_X1 u0_u14_u2_U12 (.A1( u0_u14_u2_n150 ) , .ZN( u0_u14_u2_n151 ) , .A3( u0_u14_u2_n175 ) , .A2( u0_u14_u2_n188 ) );
  AOI21_X1 u0_u14_u2_U13 (.ZN( u0_u14_u2_n144 ) , .B2( u0_u14_u2_n155 ) , .A( u0_u14_u2_n172 ) , .B1( u0_u14_u2_n185 ) );
  AOI21_X1 u0_u14_u2_U14 (.B2( u0_u14_u2_n143 ) , .ZN( u0_u14_u2_n145 ) , .B1( u0_u14_u2_n152 ) , .A( u0_u14_u2_n171 ) );
  AOI21_X1 u0_u14_u2_U15 (.B2( u0_u14_u2_n120 ) , .B1( u0_u14_u2_n121 ) , .ZN( u0_u14_u2_n126 ) , .A( u0_u14_u2_n167 ) );
  INV_X1 u0_u14_u2_U16 (.A( u0_u14_u2_n156 ) , .ZN( u0_u14_u2_n171 ) );
  INV_X1 u0_u14_u2_U17 (.A( u0_u14_u2_n120 ) , .ZN( u0_u14_u2_n188 ) );
  NAND2_X1 u0_u14_u2_U18 (.A2( u0_u14_u2_n122 ) , .ZN( u0_u14_u2_n150 ) , .A1( u0_u14_u2_n152 ) );
  INV_X1 u0_u14_u2_U19 (.A( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n170 ) );
  INV_X1 u0_u14_u2_U20 (.A( u0_u14_u2_n137 ) , .ZN( u0_u14_u2_n173 ) );
  NAND2_X1 u0_u14_u2_U21 (.A1( u0_u14_u2_n132 ) , .A2( u0_u14_u2_n139 ) , .ZN( u0_u14_u2_n157 ) );
  INV_X1 u0_u14_u2_U22 (.A( u0_u14_u2_n113 ) , .ZN( u0_u14_u2_n178 ) );
  INV_X1 u0_u14_u2_U23 (.A( u0_u14_u2_n139 ) , .ZN( u0_u14_u2_n175 ) );
  INV_X1 u0_u14_u2_U24 (.A( u0_u14_u2_n155 ) , .ZN( u0_u14_u2_n181 ) );
  INV_X1 u0_u14_u2_U25 (.A( u0_u14_u2_n119 ) , .ZN( u0_u14_u2_n177 ) );
  INV_X1 u0_u14_u2_U26 (.A( u0_u14_u2_n116 ) , .ZN( u0_u14_u2_n180 ) );
  INV_X1 u0_u14_u2_U27 (.A( u0_u14_u2_n131 ) , .ZN( u0_u14_u2_n179 ) );
  INV_X1 u0_u14_u2_U28 (.A( u0_u14_u2_n154 ) , .ZN( u0_u14_u2_n176 ) );
  NAND2_X1 u0_u14_u2_U29 (.A2( u0_u14_u2_n116 ) , .A1( u0_u14_u2_n117 ) , .ZN( u0_u14_u2_n118 ) );
  NOR2_X1 u0_u14_u2_U3 (.ZN( u0_u14_u2_n121 ) , .A2( u0_u14_u2_n177 ) , .A1( u0_u14_u2_n180 ) );
  INV_X1 u0_u14_u2_U30 (.A( u0_u14_u2_n132 ) , .ZN( u0_u14_u2_n182 ) );
  INV_X1 u0_u14_u2_U31 (.A( u0_u14_u2_n158 ) , .ZN( u0_u14_u2_n183 ) );
  OAI21_X1 u0_u14_u2_U32 (.A( u0_u14_u2_n156 ) , .B1( u0_u14_u2_n157 ) , .ZN( u0_u14_u2_n158 ) , .B2( u0_u14_u2_n179 ) );
  NOR2_X1 u0_u14_u2_U33 (.ZN( u0_u14_u2_n156 ) , .A1( u0_u14_u2_n166 ) , .A2( u0_u14_u2_n169 ) );
  NOR2_X1 u0_u14_u2_U34 (.A2( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n137 ) , .A1( u0_u14_u2_n140 ) );
  NOR2_X1 u0_u14_u2_U35 (.A2( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n153 ) , .A1( u0_u14_u2_n156 ) );
  AOI211_X1 u0_u14_u2_U36 (.ZN( u0_u14_u2_n130 ) , .C1( u0_u14_u2_n138 ) , .C2( u0_u14_u2_n179 ) , .B( u0_u14_u2_n96 ) , .A( u0_u14_u2_n97 ) );
  OAI22_X1 u0_u14_u2_U37 (.B1( u0_u14_u2_n133 ) , .A2( u0_u14_u2_n137 ) , .A1( u0_u14_u2_n152 ) , .B2( u0_u14_u2_n168 ) , .ZN( u0_u14_u2_n97 ) );
  OAI221_X1 u0_u14_u2_U38 (.B1( u0_u14_u2_n113 ) , .C1( u0_u14_u2_n132 ) , .A( u0_u14_u2_n149 ) , .B2( u0_u14_u2_n171 ) , .C2( u0_u14_u2_n172 ) , .ZN( u0_u14_u2_n96 ) );
  OAI221_X1 u0_u14_u2_U39 (.A( u0_u14_u2_n115 ) , .C2( u0_u14_u2_n123 ) , .B2( u0_u14_u2_n143 ) , .B1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n163 ) , .C1( u0_u14_u2_n168 ) );
  INV_X1 u0_u14_u2_U4 (.A( u0_u14_u2_n134 ) , .ZN( u0_u14_u2_n185 ) );
  OAI21_X1 u0_u14_u2_U40 (.A( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n115 ) , .B1( u0_u14_u2_n176 ) , .B2( u0_u14_u2_n178 ) );
  OAI221_X1 u0_u14_u2_U41 (.A( u0_u14_u2_n135 ) , .B2( u0_u14_u2_n136 ) , .B1( u0_u14_u2_n137 ) , .ZN( u0_u14_u2_n162 ) , .C2( u0_u14_u2_n167 ) , .C1( u0_u14_u2_n185 ) );
  AND3_X1 u0_u14_u2_U42 (.A3( u0_u14_u2_n131 ) , .A2( u0_u14_u2_n132 ) , .A1( u0_u14_u2_n133 ) , .ZN( u0_u14_u2_n136 ) );
  AOI22_X1 u0_u14_u2_U43 (.ZN( u0_u14_u2_n135 ) , .B1( u0_u14_u2_n140 ) , .A1( u0_u14_u2_n156 ) , .B2( u0_u14_u2_n180 ) , .A2( u0_u14_u2_n188 ) );
  AOI21_X1 u0_u14_u2_U44 (.ZN( u0_u14_u2_n149 ) , .B1( u0_u14_u2_n173 ) , .B2( u0_u14_u2_n188 ) , .A( u0_u14_u2_n95 ) );
  AND3_X1 u0_u14_u2_U45 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n156 ) , .ZN( u0_u14_u2_n95 ) );
  OAI21_X1 u0_u14_u2_U46 (.A( u0_u14_u2_n141 ) , .B2( u0_u14_u2_n142 ) , .ZN( u0_u14_u2_n146 ) , .B1( u0_u14_u2_n153 ) );
  OAI21_X1 u0_u14_u2_U47 (.A( u0_u14_u2_n140 ) , .ZN( u0_u14_u2_n141 ) , .B1( u0_u14_u2_n176 ) , .B2( u0_u14_u2_n177 ) );
  NOR3_X1 u0_u14_u2_U48 (.ZN( u0_u14_u2_n142 ) , .A3( u0_u14_u2_n175 ) , .A2( u0_u14_u2_n178 ) , .A1( u0_u14_u2_n181 ) );
  OAI21_X1 u0_u14_u2_U49 (.A( u0_u14_u2_n101 ) , .B2( u0_u14_u2_n121 ) , .B1( u0_u14_u2_n153 ) , .ZN( u0_u14_u2_n164 ) );
  INV_X1 u0_u14_u2_U5 (.A( u0_u14_u2_n150 ) , .ZN( u0_u14_u2_n184 ) );
  NAND2_X1 u0_u14_u2_U50 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n155 ) );
  NAND2_X1 u0_u14_u2_U51 (.A2( u0_u14_u2_n105 ) , .A1( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n143 ) );
  NAND2_X1 u0_u14_u2_U52 (.A1( u0_u14_u2_n104 ) , .A2( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n152 ) );
  NAND2_X1 u0_u14_u2_U53 (.A1( u0_u14_u2_n100 ) , .A2( u0_u14_u2_n105 ) , .ZN( u0_u14_u2_n132 ) );
  INV_X1 u0_u14_u2_U54 (.A( u0_u14_u2_n140 ) , .ZN( u0_u14_u2_n168 ) );
  INV_X1 u0_u14_u2_U55 (.A( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n167 ) );
  INV_X1 u0_u14_u2_U56 (.ZN( u0_u14_u2_n187 ) , .A( u0_u14_u2_n99 ) );
  OAI21_X1 u0_u14_u2_U57 (.B1( u0_u14_u2_n137 ) , .B2( u0_u14_u2_n143 ) , .A( u0_u14_u2_n98 ) , .ZN( u0_u14_u2_n99 ) );
  NAND2_X1 u0_u14_u2_U58 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n113 ) );
  NAND2_X1 u0_u14_u2_U59 (.A1( u0_u14_u2_n106 ) , .A2( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n131 ) );
  NOR4_X1 u0_u14_u2_U6 (.A4( u0_u14_u2_n124 ) , .A3( u0_u14_u2_n125 ) , .A2( u0_u14_u2_n126 ) , .A1( u0_u14_u2_n127 ) , .ZN( u0_u14_u2_n128 ) );
  NAND2_X1 u0_u14_u2_U60 (.A1( u0_u14_u2_n103 ) , .A2( u0_u14_u2_n107 ) , .ZN( u0_u14_u2_n139 ) );
  NAND2_X1 u0_u14_u2_U61 (.A1( u0_u14_u2_n103 ) , .A2( u0_u14_u2_n105 ) , .ZN( u0_u14_u2_n133 ) );
  NAND2_X1 u0_u14_u2_U62 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n103 ) , .ZN( u0_u14_u2_n154 ) );
  NAND2_X1 u0_u14_u2_U63 (.A2( u0_u14_u2_n103 ) , .A1( u0_u14_u2_n104 ) , .ZN( u0_u14_u2_n119 ) );
  NAND2_X1 u0_u14_u2_U64 (.A2( u0_u14_u2_n107 ) , .A1( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n123 ) );
  NAND2_X1 u0_u14_u2_U65 (.A1( u0_u14_u2_n104 ) , .A2( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n122 ) );
  INV_X1 u0_u14_u2_U66 (.A( u0_u14_u2_n114 ) , .ZN( u0_u14_u2_n172 ) );
  NAND2_X1 u0_u14_u2_U67 (.A2( u0_u14_u2_n100 ) , .A1( u0_u14_u2_n102 ) , .ZN( u0_u14_u2_n116 ) );
  NAND2_X1 u0_u14_u2_U68 (.A1( u0_u14_u2_n102 ) , .A2( u0_u14_u2_n108 ) , .ZN( u0_u14_u2_n120 ) );
  NAND2_X1 u0_u14_u2_U69 (.A2( u0_u14_u2_n105 ) , .A1( u0_u14_u2_n106 ) , .ZN( u0_u14_u2_n117 ) );
  AOI21_X1 u0_u14_u2_U7 (.B2( u0_u14_u2_n119 ) , .ZN( u0_u14_u2_n127 ) , .A( u0_u14_u2_n137 ) , .B1( u0_u14_u2_n155 ) );
  NOR2_X1 u0_u14_u2_U70 (.A2( u0_u14_X_16 ) , .ZN( u0_u14_u2_n140 ) , .A1( u0_u14_u2_n166 ) );
  NOR2_X1 u0_u14_u2_U71 (.A2( u0_u14_X_13 ) , .A1( u0_u14_X_14 ) , .ZN( u0_u14_u2_n100 ) );
  NOR2_X1 u0_u14_u2_U72 (.A2( u0_u14_X_16 ) , .A1( u0_u14_X_17 ) , .ZN( u0_u14_u2_n138 ) );
  NOR2_X1 u0_u14_u2_U73 (.A2( u0_u14_X_15 ) , .A1( u0_u14_X_18 ) , .ZN( u0_u14_u2_n104 ) );
  NOR2_X1 u0_u14_u2_U74 (.A2( u0_u14_X_14 ) , .ZN( u0_u14_u2_n103 ) , .A1( u0_u14_u2_n174 ) );
  NOR2_X1 u0_u14_u2_U75 (.A2( u0_u14_X_15 ) , .ZN( u0_u14_u2_n102 ) , .A1( u0_u14_u2_n165 ) );
  NOR2_X1 u0_u14_u2_U76 (.A2( u0_u14_X_17 ) , .ZN( u0_u14_u2_n114 ) , .A1( u0_u14_u2_n169 ) );
  AND2_X1 u0_u14_u2_U77 (.A1( u0_u14_X_15 ) , .ZN( u0_u14_u2_n105 ) , .A2( u0_u14_u2_n165 ) );
  AND2_X1 u0_u14_u2_U78 (.A2( u0_u14_X_15 ) , .A1( u0_u14_X_18 ) , .ZN( u0_u14_u2_n107 ) );
  AND2_X1 u0_u14_u2_U79 (.A1( u0_u14_X_14 ) , .ZN( u0_u14_u2_n106 ) , .A2( u0_u14_u2_n174 ) );
  AOI21_X1 u0_u14_u2_U8 (.ZN( u0_u14_u2_n124 ) , .B1( u0_u14_u2_n131 ) , .B2( u0_u14_u2_n143 ) , .A( u0_u14_u2_n172 ) );
  AND2_X1 u0_u14_u2_U80 (.A1( u0_u14_X_13 ) , .A2( u0_u14_X_14 ) , .ZN( u0_u14_u2_n108 ) );
  INV_X1 u0_u14_u2_U81 (.A( u0_u14_X_16 ) , .ZN( u0_u14_u2_n169 ) );
  INV_X1 u0_u14_u2_U82 (.A( u0_u14_X_17 ) , .ZN( u0_u14_u2_n166 ) );
  INV_X1 u0_u14_u2_U83 (.A( u0_u14_X_13 ) , .ZN( u0_u14_u2_n174 ) );
  INV_X1 u0_u14_u2_U84 (.A( u0_u14_X_18 ) , .ZN( u0_u14_u2_n165 ) );
  NAND4_X1 u0_u14_u2_U85 (.ZN( u0_out14_30 ) , .A4( u0_u14_u2_n147 ) , .A3( u0_u14_u2_n148 ) , .A2( u0_u14_u2_n149 ) , .A1( u0_u14_u2_n187 ) );
  NOR3_X1 u0_u14_u2_U86 (.A3( u0_u14_u2_n144 ) , .A2( u0_u14_u2_n145 ) , .A1( u0_u14_u2_n146 ) , .ZN( u0_u14_u2_n147 ) );
  AOI21_X1 u0_u14_u2_U87 (.B2( u0_u14_u2_n138 ) , .ZN( u0_u14_u2_n148 ) , .A( u0_u14_u2_n162 ) , .B1( u0_u14_u2_n182 ) );
  NAND4_X1 u0_u14_u2_U88 (.ZN( u0_out14_24 ) , .A4( u0_u14_u2_n111 ) , .A3( u0_u14_u2_n112 ) , .A1( u0_u14_u2_n130 ) , .A2( u0_u14_u2_n187 ) );
  AOI221_X1 u0_u14_u2_U89 (.A( u0_u14_u2_n109 ) , .B1( u0_u14_u2_n110 ) , .ZN( u0_u14_u2_n111 ) , .C1( u0_u14_u2_n134 ) , .C2( u0_u14_u2_n170 ) , .B2( u0_u14_u2_n173 ) );
  AOI21_X1 u0_u14_u2_U9 (.B2( u0_u14_u2_n123 ) , .ZN( u0_u14_u2_n125 ) , .A( u0_u14_u2_n171 ) , .B1( u0_u14_u2_n184 ) );
  AOI21_X1 u0_u14_u2_U90 (.ZN( u0_u14_u2_n112 ) , .B2( u0_u14_u2_n156 ) , .A( u0_u14_u2_n164 ) , .B1( u0_u14_u2_n181 ) );
  NAND4_X1 u0_u14_u2_U91 (.ZN( u0_out14_16 ) , .A4( u0_u14_u2_n128 ) , .A3( u0_u14_u2_n129 ) , .A1( u0_u14_u2_n130 ) , .A2( u0_u14_u2_n186 ) );
  AOI22_X1 u0_u14_u2_U92 (.A2( u0_u14_u2_n118 ) , .ZN( u0_u14_u2_n129 ) , .A1( u0_u14_u2_n140 ) , .B1( u0_u14_u2_n157 ) , .B2( u0_u14_u2_n170 ) );
  INV_X1 u0_u14_u2_U93 (.A( u0_u14_u2_n163 ) , .ZN( u0_u14_u2_n186 ) );
  OR4_X1 u0_u14_u2_U94 (.ZN( u0_out14_6 ) , .A4( u0_u14_u2_n161 ) , .A3( u0_u14_u2_n162 ) , .A2( u0_u14_u2_n163 ) , .A1( u0_u14_u2_n164 ) );
  OR3_X1 u0_u14_u2_U95 (.A2( u0_u14_u2_n159 ) , .A1( u0_u14_u2_n160 ) , .ZN( u0_u14_u2_n161 ) , .A3( u0_u14_u2_n183 ) );
  AOI21_X1 u0_u14_u2_U96 (.B2( u0_u14_u2_n154 ) , .B1( u0_u14_u2_n155 ) , .ZN( u0_u14_u2_n159 ) , .A( u0_u14_u2_n167 ) );
  NAND3_X1 u0_u14_u2_U97 (.A2( u0_u14_u2_n117 ) , .A1( u0_u14_u2_n122 ) , .A3( u0_u14_u2_n123 ) , .ZN( u0_u14_u2_n134 ) );
  NAND3_X1 u0_u14_u2_U98 (.ZN( u0_u14_u2_n110 ) , .A2( u0_u14_u2_n131 ) , .A3( u0_u14_u2_n139 ) , .A1( u0_u14_u2_n154 ) );
  NAND3_X1 u0_u14_u2_U99 (.A2( u0_u14_u2_n100 ) , .ZN( u0_u14_u2_n101 ) , .A1( u0_u14_u2_n104 ) , .A3( u0_u14_u2_n114 ) );
  OAI22_X1 u0_u14_u3_U10 (.B1( u0_u14_u3_n113 ) , .A2( u0_u14_u3_n135 ) , .A1( u0_u14_u3_n150 ) , .B2( u0_u14_u3_n164 ) , .ZN( u0_u14_u3_n98 ) );
  OAI211_X1 u0_u14_u3_U11 (.B( u0_u14_u3_n106 ) , .ZN( u0_u14_u3_n119 ) , .C2( u0_u14_u3_n128 ) , .C1( u0_u14_u3_n167 ) , .A( u0_u14_u3_n181 ) );
  AOI221_X1 u0_u14_u3_U12 (.C1( u0_u14_u3_n105 ) , .ZN( u0_u14_u3_n106 ) , .A( u0_u14_u3_n131 ) , .B2( u0_u14_u3_n132 ) , .C2( u0_u14_u3_n133 ) , .B1( u0_u14_u3_n169 ) );
  INV_X1 u0_u14_u3_U13 (.ZN( u0_u14_u3_n181 ) , .A( u0_u14_u3_n98 ) );
  NAND2_X1 u0_u14_u3_U14 (.ZN( u0_u14_u3_n105 ) , .A2( u0_u14_u3_n130 ) , .A1( u0_u14_u3_n155 ) );
  AOI22_X1 u0_u14_u3_U15 (.B1( u0_u14_u3_n115 ) , .A2( u0_u14_u3_n116 ) , .ZN( u0_u14_u3_n123 ) , .B2( u0_u14_u3_n133 ) , .A1( u0_u14_u3_n169 ) );
  NAND2_X1 u0_u14_u3_U16 (.ZN( u0_u14_u3_n116 ) , .A2( u0_u14_u3_n151 ) , .A1( u0_u14_u3_n182 ) );
  NOR2_X1 u0_u14_u3_U17 (.ZN( u0_u14_u3_n126 ) , .A2( u0_u14_u3_n150 ) , .A1( u0_u14_u3_n164 ) );
  AOI21_X1 u0_u14_u3_U18 (.ZN( u0_u14_u3_n112 ) , .B2( u0_u14_u3_n146 ) , .B1( u0_u14_u3_n155 ) , .A( u0_u14_u3_n167 ) );
  NAND2_X1 u0_u14_u3_U19 (.A1( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n142 ) , .A2( u0_u14_u3_n164 ) );
  NAND2_X1 u0_u14_u3_U20 (.ZN( u0_u14_u3_n132 ) , .A2( u0_u14_u3_n152 ) , .A1( u0_u14_u3_n156 ) );
  AND2_X1 u0_u14_u3_U21 (.A2( u0_u14_u3_n113 ) , .A1( u0_u14_u3_n114 ) , .ZN( u0_u14_u3_n151 ) );
  INV_X1 u0_u14_u3_U22 (.A( u0_u14_u3_n133 ) , .ZN( u0_u14_u3_n165 ) );
  INV_X1 u0_u14_u3_U23 (.A( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n170 ) );
  NAND2_X1 u0_u14_u3_U24 (.A1( u0_u14_u3_n107 ) , .A2( u0_u14_u3_n108 ) , .ZN( u0_u14_u3_n140 ) );
  NAND2_X1 u0_u14_u3_U25 (.ZN( u0_u14_u3_n117 ) , .A1( u0_u14_u3_n124 ) , .A2( u0_u14_u3_n148 ) );
  NAND2_X1 u0_u14_u3_U26 (.ZN( u0_u14_u3_n143 ) , .A1( u0_u14_u3_n165 ) , .A2( u0_u14_u3_n167 ) );
  INV_X1 u0_u14_u3_U27 (.A( u0_u14_u3_n130 ) , .ZN( u0_u14_u3_n177 ) );
  INV_X1 u0_u14_u3_U28 (.A( u0_u14_u3_n128 ) , .ZN( u0_u14_u3_n176 ) );
  INV_X1 u0_u14_u3_U29 (.A( u0_u14_u3_n155 ) , .ZN( u0_u14_u3_n174 ) );
  INV_X1 u0_u14_u3_U3 (.A( u0_u14_u3_n129 ) , .ZN( u0_u14_u3_n183 ) );
  INV_X1 u0_u14_u3_U30 (.A( u0_u14_u3_n139 ) , .ZN( u0_u14_u3_n185 ) );
  NOR2_X1 u0_u14_u3_U31 (.ZN( u0_u14_u3_n135 ) , .A2( u0_u14_u3_n141 ) , .A1( u0_u14_u3_n169 ) );
  OAI222_X1 u0_u14_u3_U32 (.C2( u0_u14_u3_n107 ) , .A2( u0_u14_u3_n108 ) , .B1( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n138 ) , .B2( u0_u14_u3_n146 ) , .C1( u0_u14_u3_n154 ) , .A1( u0_u14_u3_n164 ) );
  NOR4_X1 u0_u14_u3_U33 (.A4( u0_u14_u3_n157 ) , .A3( u0_u14_u3_n158 ) , .A2( u0_u14_u3_n159 ) , .A1( u0_u14_u3_n160 ) , .ZN( u0_u14_u3_n161 ) );
  AOI21_X1 u0_u14_u3_U34 (.B2( u0_u14_u3_n152 ) , .B1( u0_u14_u3_n153 ) , .ZN( u0_u14_u3_n158 ) , .A( u0_u14_u3_n164 ) );
  AOI21_X1 u0_u14_u3_U35 (.A( u0_u14_u3_n154 ) , .B2( u0_u14_u3_n155 ) , .B1( u0_u14_u3_n156 ) , .ZN( u0_u14_u3_n157 ) );
  AOI21_X1 u0_u14_u3_U36 (.A( u0_u14_u3_n149 ) , .B2( u0_u14_u3_n150 ) , .B1( u0_u14_u3_n151 ) , .ZN( u0_u14_u3_n159 ) );
  AOI211_X1 u0_u14_u3_U37 (.ZN( u0_u14_u3_n109 ) , .A( u0_u14_u3_n119 ) , .C2( u0_u14_u3_n129 ) , .B( u0_u14_u3_n138 ) , .C1( u0_u14_u3_n141 ) );
  AOI211_X1 u0_u14_u3_U38 (.B( u0_u14_u3_n119 ) , .A( u0_u14_u3_n120 ) , .C2( u0_u14_u3_n121 ) , .ZN( u0_u14_u3_n122 ) , .C1( u0_u14_u3_n179 ) );
  INV_X1 u0_u14_u3_U39 (.A( u0_u14_u3_n156 ) , .ZN( u0_u14_u3_n179 ) );
  INV_X1 u0_u14_u3_U4 (.A( u0_u14_u3_n140 ) , .ZN( u0_u14_u3_n182 ) );
  OAI22_X1 u0_u14_u3_U40 (.B1( u0_u14_u3_n118 ) , .ZN( u0_u14_u3_n120 ) , .A1( u0_u14_u3_n135 ) , .B2( u0_u14_u3_n154 ) , .A2( u0_u14_u3_n178 ) );
  AND3_X1 u0_u14_u3_U41 (.ZN( u0_u14_u3_n118 ) , .A2( u0_u14_u3_n124 ) , .A1( u0_u14_u3_n144 ) , .A3( u0_u14_u3_n152 ) );
  INV_X1 u0_u14_u3_U42 (.A( u0_u14_u3_n121 ) , .ZN( u0_u14_u3_n164 ) );
  NAND2_X1 u0_u14_u3_U43 (.ZN( u0_u14_u3_n133 ) , .A1( u0_u14_u3_n154 ) , .A2( u0_u14_u3_n164 ) );
  OAI211_X1 u0_u14_u3_U44 (.B( u0_u14_u3_n127 ) , .ZN( u0_u14_u3_n139 ) , .C1( u0_u14_u3_n150 ) , .C2( u0_u14_u3_n154 ) , .A( u0_u14_u3_n184 ) );
  INV_X1 u0_u14_u3_U45 (.A( u0_u14_u3_n125 ) , .ZN( u0_u14_u3_n184 ) );
  AOI221_X1 u0_u14_u3_U46 (.A( u0_u14_u3_n126 ) , .ZN( u0_u14_u3_n127 ) , .C2( u0_u14_u3_n132 ) , .C1( u0_u14_u3_n169 ) , .B2( u0_u14_u3_n170 ) , .B1( u0_u14_u3_n174 ) );
  OAI22_X1 u0_u14_u3_U47 (.A1( u0_u14_u3_n124 ) , .ZN( u0_u14_u3_n125 ) , .B2( u0_u14_u3_n145 ) , .A2( u0_u14_u3_n165 ) , .B1( u0_u14_u3_n167 ) );
  NOR2_X1 u0_u14_u3_U48 (.A1( u0_u14_u3_n113 ) , .ZN( u0_u14_u3_n131 ) , .A2( u0_u14_u3_n154 ) );
  NAND2_X1 u0_u14_u3_U49 (.A1( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n150 ) , .A2( u0_u14_u3_n99 ) );
  INV_X1 u0_u14_u3_U5 (.A( u0_u14_u3_n117 ) , .ZN( u0_u14_u3_n178 ) );
  NAND2_X1 u0_u14_u3_U50 (.A2( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n155 ) , .A1( u0_u14_u3_n97 ) );
  INV_X1 u0_u14_u3_U51 (.A( u0_u14_u3_n141 ) , .ZN( u0_u14_u3_n167 ) );
  AOI21_X1 u0_u14_u3_U52 (.B2( u0_u14_u3_n114 ) , .B1( u0_u14_u3_n146 ) , .A( u0_u14_u3_n154 ) , .ZN( u0_u14_u3_n94 ) );
  AOI21_X1 u0_u14_u3_U53 (.ZN( u0_u14_u3_n110 ) , .B2( u0_u14_u3_n142 ) , .B1( u0_u14_u3_n186 ) , .A( u0_u14_u3_n95 ) );
  INV_X1 u0_u14_u3_U54 (.A( u0_u14_u3_n145 ) , .ZN( u0_u14_u3_n186 ) );
  AOI21_X1 u0_u14_u3_U55 (.B1( u0_u14_u3_n124 ) , .A( u0_u14_u3_n149 ) , .B2( u0_u14_u3_n155 ) , .ZN( u0_u14_u3_n95 ) );
  INV_X1 u0_u14_u3_U56 (.A( u0_u14_u3_n149 ) , .ZN( u0_u14_u3_n169 ) );
  NAND2_X1 u0_u14_u3_U57 (.ZN( u0_u14_u3_n124 ) , .A1( u0_u14_u3_n96 ) , .A2( u0_u14_u3_n97 ) );
  NAND2_X1 u0_u14_u3_U58 (.A2( u0_u14_u3_n100 ) , .ZN( u0_u14_u3_n146 ) , .A1( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U59 (.A1( u0_u14_u3_n101 ) , .ZN( u0_u14_u3_n145 ) , .A2( u0_u14_u3_n99 ) );
  AOI221_X1 u0_u14_u3_U6 (.A( u0_u14_u3_n131 ) , .C2( u0_u14_u3_n132 ) , .C1( u0_u14_u3_n133 ) , .ZN( u0_u14_u3_n134 ) , .B1( u0_u14_u3_n143 ) , .B2( u0_u14_u3_n177 ) );
  NAND2_X1 u0_u14_u3_U60 (.A1( u0_u14_u3_n100 ) , .ZN( u0_u14_u3_n156 ) , .A2( u0_u14_u3_n99 ) );
  NAND2_X1 u0_u14_u3_U61 (.A2( u0_u14_u3_n101 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n148 ) );
  NAND2_X1 u0_u14_u3_U62 (.A1( u0_u14_u3_n100 ) , .A2( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n128 ) );
  NAND2_X1 u0_u14_u3_U63 (.A2( u0_u14_u3_n101 ) , .A1( u0_u14_u3_n102 ) , .ZN( u0_u14_u3_n152 ) );
  NAND2_X1 u0_u14_u3_U64 (.A2( u0_u14_u3_n101 ) , .ZN( u0_u14_u3_n114 ) , .A1( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U65 (.ZN( u0_u14_u3_n107 ) , .A1( u0_u14_u3_n97 ) , .A2( u0_u14_u3_n99 ) );
  NAND2_X1 u0_u14_u3_U66 (.A2( u0_u14_u3_n100 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n113 ) );
  NAND2_X1 u0_u14_u3_U67 (.A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n153 ) , .A2( u0_u14_u3_n97 ) );
  NAND2_X1 u0_u14_u3_U68 (.A2( u0_u14_u3_n103 ) , .A1( u0_u14_u3_n104 ) , .ZN( u0_u14_u3_n130 ) );
  NAND2_X1 u0_u14_u3_U69 (.A2( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n144 ) , .A1( u0_u14_u3_n96 ) );
  OAI22_X1 u0_u14_u3_U7 (.B2( u0_u14_u3_n147 ) , .A2( u0_u14_u3_n148 ) , .ZN( u0_u14_u3_n160 ) , .B1( u0_u14_u3_n165 ) , .A1( u0_u14_u3_n168 ) );
  NAND2_X1 u0_u14_u3_U70 (.A1( u0_u14_u3_n102 ) , .A2( u0_u14_u3_n103 ) , .ZN( u0_u14_u3_n108 ) );
  NOR2_X1 u0_u14_u3_U71 (.A2( u0_u14_X_19 ) , .A1( u0_u14_X_20 ) , .ZN( u0_u14_u3_n99 ) );
  NOR2_X1 u0_u14_u3_U72 (.A2( u0_u14_X_21 ) , .A1( u0_u14_X_24 ) , .ZN( u0_u14_u3_n103 ) );
  NOR2_X1 u0_u14_u3_U73 (.A2( u0_u14_X_24 ) , .A1( u0_u14_u3_n171 ) , .ZN( u0_u14_u3_n97 ) );
  NOR2_X1 u0_u14_u3_U74 (.A2( u0_u14_X_23 ) , .ZN( u0_u14_u3_n141 ) , .A1( u0_u14_u3_n166 ) );
  NOR2_X1 u0_u14_u3_U75 (.A2( u0_u14_X_19 ) , .A1( u0_u14_u3_n172 ) , .ZN( u0_u14_u3_n96 ) );
  NAND2_X1 u0_u14_u3_U76 (.A1( u0_u14_X_22 ) , .A2( u0_u14_X_23 ) , .ZN( u0_u14_u3_n154 ) );
  NAND2_X1 u0_u14_u3_U77 (.A1( u0_u14_X_23 ) , .ZN( u0_u14_u3_n149 ) , .A2( u0_u14_u3_n166 ) );
  NOR2_X1 u0_u14_u3_U78 (.A2( u0_u14_X_22 ) , .A1( u0_u14_X_23 ) , .ZN( u0_u14_u3_n121 ) );
  AND2_X1 u0_u14_u3_U79 (.A1( u0_u14_X_24 ) , .ZN( u0_u14_u3_n101 ) , .A2( u0_u14_u3_n171 ) );
  AND3_X1 u0_u14_u3_U8 (.A3( u0_u14_u3_n144 ) , .A2( u0_u14_u3_n145 ) , .A1( u0_u14_u3_n146 ) , .ZN( u0_u14_u3_n147 ) );
  AND2_X1 u0_u14_u3_U80 (.A1( u0_u14_X_19 ) , .ZN( u0_u14_u3_n102 ) , .A2( u0_u14_u3_n172 ) );
  AND2_X1 u0_u14_u3_U81 (.A1( u0_u14_X_21 ) , .A2( u0_u14_X_24 ) , .ZN( u0_u14_u3_n100 ) );
  AND2_X1 u0_u14_u3_U82 (.A2( u0_u14_X_19 ) , .A1( u0_u14_X_20 ) , .ZN( u0_u14_u3_n104 ) );
  INV_X1 u0_u14_u3_U83 (.A( u0_u14_X_22 ) , .ZN( u0_u14_u3_n166 ) );
  INV_X1 u0_u14_u3_U84 (.A( u0_u14_X_21 ) , .ZN( u0_u14_u3_n171 ) );
  INV_X1 u0_u14_u3_U85 (.A( u0_u14_X_20 ) , .ZN( u0_u14_u3_n172 ) );
  NAND4_X1 u0_u14_u3_U86 (.ZN( u0_out14_26 ) , .A4( u0_u14_u3_n109 ) , .A3( u0_u14_u3_n110 ) , .A2( u0_u14_u3_n111 ) , .A1( u0_u14_u3_n173 ) );
  INV_X1 u0_u14_u3_U87 (.ZN( u0_u14_u3_n173 ) , .A( u0_u14_u3_n94 ) );
  OAI21_X1 u0_u14_u3_U88 (.ZN( u0_u14_u3_n111 ) , .B2( u0_u14_u3_n117 ) , .A( u0_u14_u3_n133 ) , .B1( u0_u14_u3_n176 ) );
  NAND4_X1 u0_u14_u3_U89 (.ZN( u0_out14_20 ) , .A4( u0_u14_u3_n122 ) , .A3( u0_u14_u3_n123 ) , .A1( u0_u14_u3_n175 ) , .A2( u0_u14_u3_n180 ) );
  INV_X1 u0_u14_u3_U9 (.A( u0_u14_u3_n143 ) , .ZN( u0_u14_u3_n168 ) );
  INV_X1 u0_u14_u3_U90 (.A( u0_u14_u3_n126 ) , .ZN( u0_u14_u3_n180 ) );
  INV_X1 u0_u14_u3_U91 (.A( u0_u14_u3_n112 ) , .ZN( u0_u14_u3_n175 ) );
  NAND4_X1 u0_u14_u3_U92 (.ZN( u0_out14_1 ) , .A4( u0_u14_u3_n161 ) , .A3( u0_u14_u3_n162 ) , .A2( u0_u14_u3_n163 ) , .A1( u0_u14_u3_n185 ) );
  NAND2_X1 u0_u14_u3_U93 (.ZN( u0_u14_u3_n163 ) , .A2( u0_u14_u3_n170 ) , .A1( u0_u14_u3_n176 ) );
  AOI22_X1 u0_u14_u3_U94 (.B2( u0_u14_u3_n140 ) , .B1( u0_u14_u3_n141 ) , .A2( u0_u14_u3_n142 ) , .ZN( u0_u14_u3_n162 ) , .A1( u0_u14_u3_n177 ) );
  OR4_X1 u0_u14_u3_U95 (.ZN( u0_out14_10 ) , .A4( u0_u14_u3_n136 ) , .A3( u0_u14_u3_n137 ) , .A1( u0_u14_u3_n138 ) , .A2( u0_u14_u3_n139 ) );
  OAI222_X1 u0_u14_u3_U96 (.C1( u0_u14_u3_n128 ) , .ZN( u0_u14_u3_n137 ) , .B1( u0_u14_u3_n148 ) , .A2( u0_u14_u3_n150 ) , .B2( u0_u14_u3_n154 ) , .C2( u0_u14_u3_n164 ) , .A1( u0_u14_u3_n167 ) );
  OAI221_X1 u0_u14_u3_U97 (.A( u0_u14_u3_n134 ) , .B2( u0_u14_u3_n135 ) , .ZN( u0_u14_u3_n136 ) , .C1( u0_u14_u3_n149 ) , .B1( u0_u14_u3_n151 ) , .C2( u0_u14_u3_n183 ) );
  NAND3_X1 u0_u14_u3_U98 (.A1( u0_u14_u3_n114 ) , .ZN( u0_u14_u3_n115 ) , .A2( u0_u14_u3_n145 ) , .A3( u0_u14_u3_n153 ) );
  NAND3_X1 u0_u14_u3_U99 (.ZN( u0_u14_u3_n129 ) , .A2( u0_u14_u3_n144 ) , .A1( u0_u14_u3_n153 ) , .A3( u0_u14_u3_n182 ) );
  INV_X1 u0_u14_u5_U10 (.A( u0_u14_u5_n121 ) , .ZN( u0_u14_u5_n177 ) );
  NOR3_X1 u0_u14_u5_U100 (.A3( u0_u14_u5_n141 ) , .A1( u0_u14_u5_n142 ) , .ZN( u0_u14_u5_n143 ) , .A2( u0_u14_u5_n191 ) );
  NAND4_X1 u0_u14_u5_U101 (.ZN( u0_out14_4 ) , .A4( u0_u14_u5_n112 ) , .A2( u0_u14_u5_n113 ) , .A1( u0_u14_u5_n114 ) , .A3( u0_u14_u5_n195 ) );
  AOI211_X1 u0_u14_u5_U102 (.A( u0_u14_u5_n110 ) , .C1( u0_u14_u5_n111 ) , .ZN( u0_u14_u5_n112 ) , .B( u0_u14_u5_n118 ) , .C2( u0_u14_u5_n177 ) );
  AOI222_X1 u0_u14_u5_U103 (.ZN( u0_u14_u5_n113 ) , .A1( u0_u14_u5_n131 ) , .C1( u0_u14_u5_n148 ) , .B2( u0_u14_u5_n174 ) , .C2( u0_u14_u5_n178 ) , .A2( u0_u14_u5_n179 ) , .B1( u0_u14_u5_n99 ) );
  NAND3_X1 u0_u14_u5_U104 (.A2( u0_u14_u5_n154 ) , .A3( u0_u14_u5_n158 ) , .A1( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n99 ) );
  NOR2_X1 u0_u14_u5_U11 (.ZN( u0_u14_u5_n160 ) , .A2( u0_u14_u5_n173 ) , .A1( u0_u14_u5_n177 ) );
  INV_X1 u0_u14_u5_U12 (.A( u0_u14_u5_n150 ) , .ZN( u0_u14_u5_n174 ) );
  AOI21_X1 u0_u14_u5_U13 (.A( u0_u14_u5_n160 ) , .B2( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n162 ) , .B1( u0_u14_u5_n192 ) );
  INV_X1 u0_u14_u5_U14 (.A( u0_u14_u5_n159 ) , .ZN( u0_u14_u5_n192 ) );
  AOI21_X1 u0_u14_u5_U15 (.A( u0_u14_u5_n156 ) , .B2( u0_u14_u5_n157 ) , .B1( u0_u14_u5_n158 ) , .ZN( u0_u14_u5_n163 ) );
  AOI21_X1 u0_u14_u5_U16 (.B2( u0_u14_u5_n139 ) , .B1( u0_u14_u5_n140 ) , .ZN( u0_u14_u5_n141 ) , .A( u0_u14_u5_n150 ) );
  OAI21_X1 u0_u14_u5_U17 (.A( u0_u14_u5_n133 ) , .B2( u0_u14_u5_n134 ) , .B1( u0_u14_u5_n135 ) , .ZN( u0_u14_u5_n142 ) );
  OAI21_X1 u0_u14_u5_U18 (.ZN( u0_u14_u5_n133 ) , .B2( u0_u14_u5_n147 ) , .A( u0_u14_u5_n173 ) , .B1( u0_u14_u5_n188 ) );
  NAND2_X1 u0_u14_u5_U19 (.A2( u0_u14_u5_n119 ) , .A1( u0_u14_u5_n123 ) , .ZN( u0_u14_u5_n137 ) );
  INV_X1 u0_u14_u5_U20 (.A( u0_u14_u5_n155 ) , .ZN( u0_u14_u5_n194 ) );
  NAND2_X1 u0_u14_u5_U21 (.A1( u0_u14_u5_n121 ) , .ZN( u0_u14_u5_n132 ) , .A2( u0_u14_u5_n172 ) );
  NAND2_X1 u0_u14_u5_U22 (.A2( u0_u14_u5_n122 ) , .ZN( u0_u14_u5_n136 ) , .A1( u0_u14_u5_n154 ) );
  NAND2_X1 u0_u14_u5_U23 (.A2( u0_u14_u5_n119 ) , .A1( u0_u14_u5_n120 ) , .ZN( u0_u14_u5_n159 ) );
  INV_X1 u0_u14_u5_U24 (.A( u0_u14_u5_n156 ) , .ZN( u0_u14_u5_n175 ) );
  INV_X1 u0_u14_u5_U25 (.A( u0_u14_u5_n158 ) , .ZN( u0_u14_u5_n188 ) );
  INV_X1 u0_u14_u5_U26 (.A( u0_u14_u5_n152 ) , .ZN( u0_u14_u5_n179 ) );
  INV_X1 u0_u14_u5_U27 (.A( u0_u14_u5_n140 ) , .ZN( u0_u14_u5_n182 ) );
  INV_X1 u0_u14_u5_U28 (.A( u0_u14_u5_n151 ) , .ZN( u0_u14_u5_n183 ) );
  INV_X1 u0_u14_u5_U29 (.A( u0_u14_u5_n123 ) , .ZN( u0_u14_u5_n185 ) );
  NOR2_X1 u0_u14_u5_U3 (.ZN( u0_u14_u5_n134 ) , .A1( u0_u14_u5_n183 ) , .A2( u0_u14_u5_n190 ) );
  INV_X1 u0_u14_u5_U30 (.A( u0_u14_u5_n161 ) , .ZN( u0_u14_u5_n184 ) );
  INV_X1 u0_u14_u5_U31 (.A( u0_u14_u5_n139 ) , .ZN( u0_u14_u5_n189 ) );
  INV_X1 u0_u14_u5_U32 (.A( u0_u14_u5_n157 ) , .ZN( u0_u14_u5_n190 ) );
  INV_X1 u0_u14_u5_U33 (.A( u0_u14_u5_n120 ) , .ZN( u0_u14_u5_n193 ) );
  NAND2_X1 u0_u14_u5_U34 (.ZN( u0_u14_u5_n111 ) , .A1( u0_u14_u5_n140 ) , .A2( u0_u14_u5_n155 ) );
  INV_X1 u0_u14_u5_U35 (.A( u0_u14_u5_n117 ) , .ZN( u0_u14_u5_n196 ) );
  OAI221_X1 u0_u14_u5_U36 (.A( u0_u14_u5_n116 ) , .ZN( u0_u14_u5_n117 ) , .B2( u0_u14_u5_n119 ) , .C1( u0_u14_u5_n153 ) , .C2( u0_u14_u5_n158 ) , .B1( u0_u14_u5_n172 ) );
  AOI222_X1 u0_u14_u5_U37 (.ZN( u0_u14_u5_n116 ) , .B2( u0_u14_u5_n145 ) , .C1( u0_u14_u5_n148 ) , .A2( u0_u14_u5_n174 ) , .C2( u0_u14_u5_n177 ) , .B1( u0_u14_u5_n187 ) , .A1( u0_u14_u5_n193 ) );
  INV_X1 u0_u14_u5_U38 (.A( u0_u14_u5_n115 ) , .ZN( u0_u14_u5_n187 ) );
  NOR2_X1 u0_u14_u5_U39 (.ZN( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n170 ) , .A2( u0_u14_u5_n180 ) );
  INV_X1 u0_u14_u5_U4 (.A( u0_u14_u5_n138 ) , .ZN( u0_u14_u5_n191 ) );
  AOI22_X1 u0_u14_u5_U40 (.B2( u0_u14_u5_n131 ) , .A2( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n169 ) , .B1( u0_u14_u5_n174 ) , .A1( u0_u14_u5_n185 ) );
  NOR2_X1 u0_u14_u5_U41 (.A1( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n150 ) , .A2( u0_u14_u5_n173 ) );
  AOI21_X1 u0_u14_u5_U42 (.A( u0_u14_u5_n118 ) , .B2( u0_u14_u5_n145 ) , .ZN( u0_u14_u5_n168 ) , .B1( u0_u14_u5_n186 ) );
  INV_X1 u0_u14_u5_U43 (.A( u0_u14_u5_n122 ) , .ZN( u0_u14_u5_n186 ) );
  NOR2_X1 u0_u14_u5_U44 (.A1( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n152 ) , .A2( u0_u14_u5_n176 ) );
  NOR2_X1 u0_u14_u5_U45 (.A1( u0_u14_u5_n115 ) , .ZN( u0_u14_u5_n118 ) , .A2( u0_u14_u5_n153 ) );
  NOR2_X1 u0_u14_u5_U46 (.A2( u0_u14_u5_n145 ) , .ZN( u0_u14_u5_n156 ) , .A1( u0_u14_u5_n174 ) );
  NOR2_X1 u0_u14_u5_U47 (.ZN( u0_u14_u5_n121 ) , .A2( u0_u14_u5_n145 ) , .A1( u0_u14_u5_n176 ) );
  AOI22_X1 u0_u14_u5_U48 (.ZN( u0_u14_u5_n114 ) , .A2( u0_u14_u5_n137 ) , .A1( u0_u14_u5_n145 ) , .B2( u0_u14_u5_n175 ) , .B1( u0_u14_u5_n193 ) );
  OAI211_X1 u0_u14_u5_U49 (.B( u0_u14_u5_n124 ) , .A( u0_u14_u5_n125 ) , .C2( u0_u14_u5_n126 ) , .C1( u0_u14_u5_n127 ) , .ZN( u0_u14_u5_n128 ) );
  OAI21_X1 u0_u14_u5_U5 (.B2( u0_u14_u5_n136 ) , .B1( u0_u14_u5_n137 ) , .ZN( u0_u14_u5_n138 ) , .A( u0_u14_u5_n177 ) );
  NOR3_X1 u0_u14_u5_U50 (.ZN( u0_u14_u5_n127 ) , .A1( u0_u14_u5_n136 ) , .A3( u0_u14_u5_n148 ) , .A2( u0_u14_u5_n182 ) );
  OAI21_X1 u0_u14_u5_U51 (.ZN( u0_u14_u5_n124 ) , .A( u0_u14_u5_n177 ) , .B2( u0_u14_u5_n183 ) , .B1( u0_u14_u5_n189 ) );
  OAI21_X1 u0_u14_u5_U52 (.ZN( u0_u14_u5_n125 ) , .A( u0_u14_u5_n174 ) , .B2( u0_u14_u5_n185 ) , .B1( u0_u14_u5_n190 ) );
  AOI21_X1 u0_u14_u5_U53 (.A( u0_u14_u5_n153 ) , .B2( u0_u14_u5_n154 ) , .B1( u0_u14_u5_n155 ) , .ZN( u0_u14_u5_n164 ) );
  AOI21_X1 u0_u14_u5_U54 (.ZN( u0_u14_u5_n110 ) , .B1( u0_u14_u5_n122 ) , .B2( u0_u14_u5_n139 ) , .A( u0_u14_u5_n153 ) );
  INV_X1 u0_u14_u5_U55 (.A( u0_u14_u5_n153 ) , .ZN( u0_u14_u5_n176 ) );
  INV_X1 u0_u14_u5_U56 (.A( u0_u14_u5_n126 ) , .ZN( u0_u14_u5_n173 ) );
  AND2_X1 u0_u14_u5_U57 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n147 ) );
  AND2_X1 u0_u14_u5_U58 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n148 ) );
  NAND2_X1 u0_u14_u5_U59 (.A1( u0_u14_u5_n105 ) , .A2( u0_u14_u5_n106 ) , .ZN( u0_u14_u5_n158 ) );
  INV_X1 u0_u14_u5_U6 (.A( u0_u14_u5_n135 ) , .ZN( u0_u14_u5_n178 ) );
  NAND2_X1 u0_u14_u5_U60 (.A2( u0_u14_u5_n108 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n139 ) );
  NAND2_X1 u0_u14_u5_U61 (.A1( u0_u14_u5_n106 ) , .A2( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n119 ) );
  NAND2_X1 u0_u14_u5_U62 (.A2( u0_u14_u5_n103 ) , .A1( u0_u14_u5_n105 ) , .ZN( u0_u14_u5_n140 ) );
  NAND2_X1 u0_u14_u5_U63 (.A2( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n105 ) , .ZN( u0_u14_u5_n155 ) );
  NAND2_X1 u0_u14_u5_U64 (.A2( u0_u14_u5_n106 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n122 ) );
  NAND2_X1 u0_u14_u5_U65 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n106 ) , .ZN( u0_u14_u5_n115 ) );
  NAND2_X1 u0_u14_u5_U66 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n103 ) , .ZN( u0_u14_u5_n161 ) );
  NAND2_X1 u0_u14_u5_U67 (.A1( u0_u14_u5_n105 ) , .A2( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n154 ) );
  INV_X1 u0_u14_u5_U68 (.A( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n172 ) );
  NAND2_X1 u0_u14_u5_U69 (.A1( u0_u14_u5_n103 ) , .A2( u0_u14_u5_n108 ) , .ZN( u0_u14_u5_n123 ) );
  OAI22_X1 u0_u14_u5_U7 (.B2( u0_u14_u5_n149 ) , .B1( u0_u14_u5_n150 ) , .A2( u0_u14_u5_n151 ) , .A1( u0_u14_u5_n152 ) , .ZN( u0_u14_u5_n165 ) );
  NAND2_X1 u0_u14_u5_U70 (.A2( u0_u14_u5_n103 ) , .A1( u0_u14_u5_n107 ) , .ZN( u0_u14_u5_n151 ) );
  NAND2_X1 u0_u14_u5_U71 (.A2( u0_u14_u5_n107 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n120 ) );
  NAND2_X1 u0_u14_u5_U72 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n109 ) , .ZN( u0_u14_u5_n157 ) );
  AND2_X1 u0_u14_u5_U73 (.A2( u0_u14_u5_n100 ) , .A1( u0_u14_u5_n104 ) , .ZN( u0_u14_u5_n131 ) );
  INV_X1 u0_u14_u5_U74 (.A( u0_u14_u5_n102 ) , .ZN( u0_u14_u5_n195 ) );
  OAI221_X1 u0_u14_u5_U75 (.A( u0_u14_u5_n101 ) , .ZN( u0_u14_u5_n102 ) , .C2( u0_u14_u5_n115 ) , .C1( u0_u14_u5_n126 ) , .B1( u0_u14_u5_n134 ) , .B2( u0_u14_u5_n160 ) );
  OAI21_X1 u0_u14_u5_U76 (.ZN( u0_u14_u5_n101 ) , .B1( u0_u14_u5_n137 ) , .A( u0_u14_u5_n146 ) , .B2( u0_u14_u5_n147 ) );
  NOR2_X1 u0_u14_u5_U77 (.A2( u0_u14_X_34 ) , .A1( u0_u14_X_35 ) , .ZN( u0_u14_u5_n145 ) );
  NOR2_X1 u0_u14_u5_U78 (.A2( u0_u14_X_34 ) , .ZN( u0_u14_u5_n146 ) , .A1( u0_u14_u5_n171 ) );
  NOR2_X1 u0_u14_u5_U79 (.A2( u0_u14_X_31 ) , .A1( u0_u14_X_32 ) , .ZN( u0_u14_u5_n103 ) );
  NOR3_X1 u0_u14_u5_U8 (.A2( u0_u14_u5_n147 ) , .A1( u0_u14_u5_n148 ) , .ZN( u0_u14_u5_n149 ) , .A3( u0_u14_u5_n194 ) );
  NOR2_X1 u0_u14_u5_U80 (.A2( u0_u14_X_36 ) , .ZN( u0_u14_u5_n105 ) , .A1( u0_u14_u5_n180 ) );
  NOR2_X1 u0_u14_u5_U81 (.A2( u0_u14_X_33 ) , .ZN( u0_u14_u5_n108 ) , .A1( u0_u14_u5_n170 ) );
  NOR2_X1 u0_u14_u5_U82 (.A2( u0_u14_X_33 ) , .A1( u0_u14_X_36 ) , .ZN( u0_u14_u5_n107 ) );
  NOR2_X1 u0_u14_u5_U83 (.A2( u0_u14_X_31 ) , .ZN( u0_u14_u5_n104 ) , .A1( u0_u14_u5_n181 ) );
  NAND2_X1 u0_u14_u5_U84 (.A2( u0_u14_X_34 ) , .A1( u0_u14_X_35 ) , .ZN( u0_u14_u5_n153 ) );
  NAND2_X1 u0_u14_u5_U85 (.A1( u0_u14_X_34 ) , .ZN( u0_u14_u5_n126 ) , .A2( u0_u14_u5_n171 ) );
  AND2_X1 u0_u14_u5_U86 (.A1( u0_u14_X_31 ) , .A2( u0_u14_X_32 ) , .ZN( u0_u14_u5_n106 ) );
  AND2_X1 u0_u14_u5_U87 (.A1( u0_u14_X_31 ) , .ZN( u0_u14_u5_n109 ) , .A2( u0_u14_u5_n181 ) );
  INV_X1 u0_u14_u5_U88 (.A( u0_u14_X_33 ) , .ZN( u0_u14_u5_n180 ) );
  INV_X1 u0_u14_u5_U89 (.A( u0_u14_X_35 ) , .ZN( u0_u14_u5_n171 ) );
  NOR2_X1 u0_u14_u5_U9 (.ZN( u0_u14_u5_n135 ) , .A1( u0_u14_u5_n173 ) , .A2( u0_u14_u5_n176 ) );
  INV_X1 u0_u14_u5_U90 (.A( u0_u14_X_36 ) , .ZN( u0_u14_u5_n170 ) );
  INV_X1 u0_u14_u5_U91 (.A( u0_u14_X_32 ) , .ZN( u0_u14_u5_n181 ) );
  NAND4_X1 u0_u14_u5_U92 (.ZN( u0_out14_29 ) , .A4( u0_u14_u5_n129 ) , .A3( u0_u14_u5_n130 ) , .A2( u0_u14_u5_n168 ) , .A1( u0_u14_u5_n196 ) );
  AOI221_X1 u0_u14_u5_U93 (.A( u0_u14_u5_n128 ) , .ZN( u0_u14_u5_n129 ) , .C2( u0_u14_u5_n132 ) , .B2( u0_u14_u5_n159 ) , .B1( u0_u14_u5_n176 ) , .C1( u0_u14_u5_n184 ) );
  AOI222_X1 u0_u14_u5_U94 (.ZN( u0_u14_u5_n130 ) , .A2( u0_u14_u5_n146 ) , .B1( u0_u14_u5_n147 ) , .C2( u0_u14_u5_n175 ) , .B2( u0_u14_u5_n179 ) , .A1( u0_u14_u5_n188 ) , .C1( u0_u14_u5_n194 ) );
  NAND4_X1 u0_u14_u5_U95 (.ZN( u0_out14_19 ) , .A4( u0_u14_u5_n166 ) , .A3( u0_u14_u5_n167 ) , .A2( u0_u14_u5_n168 ) , .A1( u0_u14_u5_n169 ) );
  AOI22_X1 u0_u14_u5_U96 (.B2( u0_u14_u5_n145 ) , .A2( u0_u14_u5_n146 ) , .ZN( u0_u14_u5_n167 ) , .B1( u0_u14_u5_n182 ) , .A1( u0_u14_u5_n189 ) );
  NOR4_X1 u0_u14_u5_U97 (.A4( u0_u14_u5_n162 ) , .A3( u0_u14_u5_n163 ) , .A2( u0_u14_u5_n164 ) , .A1( u0_u14_u5_n165 ) , .ZN( u0_u14_u5_n166 ) );
  NAND4_X1 u0_u14_u5_U98 (.ZN( u0_out14_11 ) , .A4( u0_u14_u5_n143 ) , .A3( u0_u14_u5_n144 ) , .A2( u0_u14_u5_n169 ) , .A1( u0_u14_u5_n196 ) );
  AOI22_X1 u0_u14_u5_U99 (.A2( u0_u14_u5_n132 ) , .ZN( u0_u14_u5_n144 ) , .B2( u0_u14_u5_n145 ) , .B1( u0_u14_u5_n184 ) , .A1( u0_u14_u5_n194 ) );
  XOR2_X1 u0_u15_U10 (.A( u0_FP_62 ) , .B( u0_K16_45 ) , .Z( u0_u15_X_45 ) );
  XOR2_X1 u0_u15_U11 (.A( u0_FP_61 ) , .B( u0_K16_44 ) , .Z( u0_u15_X_44 ) );
  XOR2_X1 u0_u15_U12 (.A( u0_FP_60 ) , .B( u0_K16_43 ) , .Z( u0_u15_X_43 ) );
  XOR2_X1 u0_u15_U13 (.A( u0_FP_61 ) , .B( u0_K16_42 ) , .Z( u0_u15_X_42 ) );
  XOR2_X1 u0_u15_U14 (.A( u0_FP_60 ) , .B( u0_K16_41 ) , .Z( u0_u15_X_41 ) );
  XOR2_X1 u0_u15_U15 (.A( u0_FP_59 ) , .B( u0_K16_40 ) , .Z( u0_u15_X_40 ) );
  XOR2_X1 u0_u15_U17 (.A( u0_FP_58 ) , .B( u0_K16_39 ) , .Z( u0_u15_X_39 ) );
  XOR2_X1 u0_u15_U18 (.A( u0_FP_57 ) , .B( u0_K16_38 ) , .Z( u0_u15_X_38 ) );
  XOR2_X1 u0_u15_U19 (.A( u0_FP_56 ) , .B( u0_K16_37 ) , .Z( u0_u15_X_37 ) );
  XOR2_X1 u0_u15_U20 (.A( u0_FP_57 ) , .B( u0_K16_36 ) , .Z( u0_u15_X_36 ) );
  XOR2_X1 u0_u15_U21 (.A( u0_FP_56 ) , .B( u0_K16_35 ) , .Z( u0_u15_X_35 ) );
  XOR2_X1 u0_u15_U22 (.A( u0_FP_55 ) , .B( u0_K16_34 ) , .Z( u0_u15_X_34 ) );
  XOR2_X1 u0_u15_U23 (.A( u0_FP_54 ) , .B( u0_K16_33 ) , .Z( u0_u15_X_33 ) );
  XOR2_X1 u0_u15_U24 (.A( u0_FP_53 ) , .B( u0_K16_32 ) , .Z( u0_u15_X_32 ) );
  XOR2_X1 u0_u15_U25 (.A( u0_FP_52 ) , .B( u0_K16_31 ) , .Z( u0_u15_X_31 ) );
  XOR2_X1 u0_u15_U7 (.A( u0_FP_33 ) , .B( u0_K16_48 ) , .Z( u0_u15_X_48 ) );
  XOR2_X1 u0_u15_U8 (.A( u0_FP_64 ) , .B( u0_K16_47 ) , .Z( u0_u15_X_47 ) );
  XOR2_X1 u0_u15_U9 (.A( u0_FP_63 ) , .B( u0_K16_46 ) , .Z( u0_u15_X_46 ) );
  INV_X1 u0_u15_u5_U10 (.A( u0_u15_u5_n121 ) , .ZN( u0_u15_u5_n177 ) );
  AOI222_X1 u0_u15_u5_U100 (.ZN( u0_u15_u5_n113 ) , .A1( u0_u15_u5_n131 ) , .C1( u0_u15_u5_n148 ) , .B2( u0_u15_u5_n174 ) , .C2( u0_u15_u5_n178 ) , .A2( u0_u15_u5_n179 ) , .B1( u0_u15_u5_n99 ) );
  NAND4_X1 u0_u15_u5_U101 (.ZN( u0_out15_29 ) , .A4( u0_u15_u5_n129 ) , .A3( u0_u15_u5_n130 ) , .A2( u0_u15_u5_n168 ) , .A1( u0_u15_u5_n196 ) );
  AOI221_X1 u0_u15_u5_U102 (.A( u0_u15_u5_n128 ) , .ZN( u0_u15_u5_n129 ) , .C2( u0_u15_u5_n132 ) , .B2( u0_u15_u5_n159 ) , .B1( u0_u15_u5_n176 ) , .C1( u0_u15_u5_n184 ) );
  AOI222_X1 u0_u15_u5_U103 (.ZN( u0_u15_u5_n130 ) , .A2( u0_u15_u5_n146 ) , .B1( u0_u15_u5_n147 ) , .C2( u0_u15_u5_n175 ) , .B2( u0_u15_u5_n179 ) , .A1( u0_u15_u5_n188 ) , .C1( u0_u15_u5_n194 ) );
  NAND3_X1 u0_u15_u5_U104 (.A2( u0_u15_u5_n154 ) , .A3( u0_u15_u5_n158 ) , .A1( u0_u15_u5_n161 ) , .ZN( u0_u15_u5_n99 ) );
  NOR2_X1 u0_u15_u5_U11 (.ZN( u0_u15_u5_n160 ) , .A2( u0_u15_u5_n173 ) , .A1( u0_u15_u5_n177 ) );
  INV_X1 u0_u15_u5_U12 (.A( u0_u15_u5_n150 ) , .ZN( u0_u15_u5_n174 ) );
  AOI21_X1 u0_u15_u5_U13 (.A( u0_u15_u5_n160 ) , .B2( u0_u15_u5_n161 ) , .ZN( u0_u15_u5_n162 ) , .B1( u0_u15_u5_n192 ) );
  INV_X1 u0_u15_u5_U14 (.A( u0_u15_u5_n159 ) , .ZN( u0_u15_u5_n192 ) );
  AOI21_X1 u0_u15_u5_U15 (.A( u0_u15_u5_n156 ) , .B2( u0_u15_u5_n157 ) , .B1( u0_u15_u5_n158 ) , .ZN( u0_u15_u5_n163 ) );
  AOI21_X1 u0_u15_u5_U16 (.B2( u0_u15_u5_n139 ) , .B1( u0_u15_u5_n140 ) , .ZN( u0_u15_u5_n141 ) , .A( u0_u15_u5_n150 ) );
  OAI21_X1 u0_u15_u5_U17 (.A( u0_u15_u5_n133 ) , .B2( u0_u15_u5_n134 ) , .B1( u0_u15_u5_n135 ) , .ZN( u0_u15_u5_n142 ) );
  OAI21_X1 u0_u15_u5_U18 (.ZN( u0_u15_u5_n133 ) , .B2( u0_u15_u5_n147 ) , .A( u0_u15_u5_n173 ) , .B1( u0_u15_u5_n188 ) );
  NAND2_X1 u0_u15_u5_U19 (.A2( u0_u15_u5_n119 ) , .A1( u0_u15_u5_n123 ) , .ZN( u0_u15_u5_n137 ) );
  INV_X1 u0_u15_u5_U20 (.A( u0_u15_u5_n155 ) , .ZN( u0_u15_u5_n194 ) );
  NAND2_X1 u0_u15_u5_U21 (.A1( u0_u15_u5_n121 ) , .ZN( u0_u15_u5_n132 ) , .A2( u0_u15_u5_n172 ) );
  NAND2_X1 u0_u15_u5_U22 (.A2( u0_u15_u5_n122 ) , .ZN( u0_u15_u5_n136 ) , .A1( u0_u15_u5_n154 ) );
  NAND2_X1 u0_u15_u5_U23 (.A2( u0_u15_u5_n119 ) , .A1( u0_u15_u5_n120 ) , .ZN( u0_u15_u5_n159 ) );
  INV_X1 u0_u15_u5_U24 (.A( u0_u15_u5_n156 ) , .ZN( u0_u15_u5_n175 ) );
  INV_X1 u0_u15_u5_U25 (.A( u0_u15_u5_n158 ) , .ZN( u0_u15_u5_n188 ) );
  INV_X1 u0_u15_u5_U26 (.A( u0_u15_u5_n152 ) , .ZN( u0_u15_u5_n179 ) );
  INV_X1 u0_u15_u5_U27 (.A( u0_u15_u5_n140 ) , .ZN( u0_u15_u5_n182 ) );
  INV_X1 u0_u15_u5_U28 (.A( u0_u15_u5_n151 ) , .ZN( u0_u15_u5_n183 ) );
  INV_X1 u0_u15_u5_U29 (.A( u0_u15_u5_n123 ) , .ZN( u0_u15_u5_n185 ) );
  NOR2_X1 u0_u15_u5_U3 (.ZN( u0_u15_u5_n134 ) , .A1( u0_u15_u5_n183 ) , .A2( u0_u15_u5_n190 ) );
  INV_X1 u0_u15_u5_U30 (.A( u0_u15_u5_n161 ) , .ZN( u0_u15_u5_n184 ) );
  INV_X1 u0_u15_u5_U31 (.A( u0_u15_u5_n139 ) , .ZN( u0_u15_u5_n189 ) );
  INV_X1 u0_u15_u5_U32 (.A( u0_u15_u5_n157 ) , .ZN( u0_u15_u5_n190 ) );
  INV_X1 u0_u15_u5_U33 (.A( u0_u15_u5_n120 ) , .ZN( u0_u15_u5_n193 ) );
  NAND2_X1 u0_u15_u5_U34 (.ZN( u0_u15_u5_n111 ) , .A1( u0_u15_u5_n140 ) , .A2( u0_u15_u5_n155 ) );
  NOR2_X1 u0_u15_u5_U35 (.ZN( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n170 ) , .A2( u0_u15_u5_n180 ) );
  INV_X1 u0_u15_u5_U36 (.A( u0_u15_u5_n117 ) , .ZN( u0_u15_u5_n196 ) );
  OAI221_X1 u0_u15_u5_U37 (.A( u0_u15_u5_n116 ) , .ZN( u0_u15_u5_n117 ) , .B2( u0_u15_u5_n119 ) , .C1( u0_u15_u5_n153 ) , .C2( u0_u15_u5_n158 ) , .B1( u0_u15_u5_n172 ) );
  AOI222_X1 u0_u15_u5_U38 (.ZN( u0_u15_u5_n116 ) , .B2( u0_u15_u5_n145 ) , .C1( u0_u15_u5_n148 ) , .A2( u0_u15_u5_n174 ) , .C2( u0_u15_u5_n177 ) , .B1( u0_u15_u5_n187 ) , .A1( u0_u15_u5_n193 ) );
  INV_X1 u0_u15_u5_U39 (.A( u0_u15_u5_n115 ) , .ZN( u0_u15_u5_n187 ) );
  INV_X1 u0_u15_u5_U4 (.A( u0_u15_u5_n138 ) , .ZN( u0_u15_u5_n191 ) );
  AOI22_X1 u0_u15_u5_U40 (.B2( u0_u15_u5_n131 ) , .A2( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n169 ) , .B1( u0_u15_u5_n174 ) , .A1( u0_u15_u5_n185 ) );
  NOR2_X1 u0_u15_u5_U41 (.A1( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n150 ) , .A2( u0_u15_u5_n173 ) );
  AOI21_X1 u0_u15_u5_U42 (.A( u0_u15_u5_n118 ) , .B2( u0_u15_u5_n145 ) , .ZN( u0_u15_u5_n168 ) , .B1( u0_u15_u5_n186 ) );
  INV_X1 u0_u15_u5_U43 (.A( u0_u15_u5_n122 ) , .ZN( u0_u15_u5_n186 ) );
  NOR2_X1 u0_u15_u5_U44 (.A1( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n152 ) , .A2( u0_u15_u5_n176 ) );
  NOR2_X1 u0_u15_u5_U45 (.A1( u0_u15_u5_n115 ) , .ZN( u0_u15_u5_n118 ) , .A2( u0_u15_u5_n153 ) );
  NOR2_X1 u0_u15_u5_U46 (.A2( u0_u15_u5_n145 ) , .ZN( u0_u15_u5_n156 ) , .A1( u0_u15_u5_n174 ) );
  NOR2_X1 u0_u15_u5_U47 (.ZN( u0_u15_u5_n121 ) , .A2( u0_u15_u5_n145 ) , .A1( u0_u15_u5_n176 ) );
  AOI22_X1 u0_u15_u5_U48 (.ZN( u0_u15_u5_n114 ) , .A2( u0_u15_u5_n137 ) , .A1( u0_u15_u5_n145 ) , .B2( u0_u15_u5_n175 ) , .B1( u0_u15_u5_n193 ) );
  OAI211_X1 u0_u15_u5_U49 (.B( u0_u15_u5_n124 ) , .A( u0_u15_u5_n125 ) , .C2( u0_u15_u5_n126 ) , .C1( u0_u15_u5_n127 ) , .ZN( u0_u15_u5_n128 ) );
  OAI21_X1 u0_u15_u5_U5 (.B2( u0_u15_u5_n136 ) , .B1( u0_u15_u5_n137 ) , .ZN( u0_u15_u5_n138 ) , .A( u0_u15_u5_n177 ) );
  NOR3_X1 u0_u15_u5_U50 (.ZN( u0_u15_u5_n127 ) , .A1( u0_u15_u5_n136 ) , .A3( u0_u15_u5_n148 ) , .A2( u0_u15_u5_n182 ) );
  OAI21_X1 u0_u15_u5_U51 (.ZN( u0_u15_u5_n124 ) , .A( u0_u15_u5_n177 ) , .B2( u0_u15_u5_n183 ) , .B1( u0_u15_u5_n189 ) );
  OAI21_X1 u0_u15_u5_U52 (.ZN( u0_u15_u5_n125 ) , .A( u0_u15_u5_n174 ) , .B2( u0_u15_u5_n185 ) , .B1( u0_u15_u5_n190 ) );
  AOI21_X1 u0_u15_u5_U53 (.A( u0_u15_u5_n153 ) , .B2( u0_u15_u5_n154 ) , .B1( u0_u15_u5_n155 ) , .ZN( u0_u15_u5_n164 ) );
  AOI21_X1 u0_u15_u5_U54 (.ZN( u0_u15_u5_n110 ) , .B1( u0_u15_u5_n122 ) , .B2( u0_u15_u5_n139 ) , .A( u0_u15_u5_n153 ) );
  INV_X1 u0_u15_u5_U55 (.A( u0_u15_u5_n153 ) , .ZN( u0_u15_u5_n176 ) );
  INV_X1 u0_u15_u5_U56 (.A( u0_u15_u5_n126 ) , .ZN( u0_u15_u5_n173 ) );
  AND2_X1 u0_u15_u5_U57 (.A2( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n107 ) , .ZN( u0_u15_u5_n147 ) );
  AND2_X1 u0_u15_u5_U58 (.A2( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n108 ) , .ZN( u0_u15_u5_n148 ) );
  NAND2_X1 u0_u15_u5_U59 (.A1( u0_u15_u5_n105 ) , .A2( u0_u15_u5_n106 ) , .ZN( u0_u15_u5_n158 ) );
  INV_X1 u0_u15_u5_U6 (.A( u0_u15_u5_n135 ) , .ZN( u0_u15_u5_n178 ) );
  NAND2_X1 u0_u15_u5_U60 (.A2( u0_u15_u5_n108 ) , .A1( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n139 ) );
  NAND2_X1 u0_u15_u5_U61 (.A1( u0_u15_u5_n106 ) , .A2( u0_u15_u5_n108 ) , .ZN( u0_u15_u5_n119 ) );
  NAND2_X1 u0_u15_u5_U62 (.A2( u0_u15_u5_n103 ) , .A1( u0_u15_u5_n105 ) , .ZN( u0_u15_u5_n140 ) );
  NAND2_X1 u0_u15_u5_U63 (.A2( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n105 ) , .ZN( u0_u15_u5_n155 ) );
  NAND2_X1 u0_u15_u5_U64 (.A2( u0_u15_u5_n106 ) , .A1( u0_u15_u5_n107 ) , .ZN( u0_u15_u5_n122 ) );
  NAND2_X1 u0_u15_u5_U65 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n106 ) , .ZN( u0_u15_u5_n115 ) );
  NAND2_X1 u0_u15_u5_U66 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n103 ) , .ZN( u0_u15_u5_n161 ) );
  NAND2_X1 u0_u15_u5_U67 (.A1( u0_u15_u5_n105 ) , .A2( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n154 ) );
  INV_X1 u0_u15_u5_U68 (.A( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n172 ) );
  NAND2_X1 u0_u15_u5_U69 (.A1( u0_u15_u5_n103 ) , .A2( u0_u15_u5_n108 ) , .ZN( u0_u15_u5_n123 ) );
  OAI22_X1 u0_u15_u5_U7 (.B2( u0_u15_u5_n149 ) , .B1( u0_u15_u5_n150 ) , .A2( u0_u15_u5_n151 ) , .A1( u0_u15_u5_n152 ) , .ZN( u0_u15_u5_n165 ) );
  NAND2_X1 u0_u15_u5_U70 (.A2( u0_u15_u5_n103 ) , .A1( u0_u15_u5_n107 ) , .ZN( u0_u15_u5_n151 ) );
  NAND2_X1 u0_u15_u5_U71 (.A2( u0_u15_u5_n107 ) , .A1( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n120 ) );
  NAND2_X1 u0_u15_u5_U72 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n109 ) , .ZN( u0_u15_u5_n157 ) );
  AND2_X1 u0_u15_u5_U73 (.A2( u0_u15_u5_n100 ) , .A1( u0_u15_u5_n104 ) , .ZN( u0_u15_u5_n131 ) );
  INV_X1 u0_u15_u5_U74 (.A( u0_u15_u5_n102 ) , .ZN( u0_u15_u5_n195 ) );
  OAI221_X1 u0_u15_u5_U75 (.A( u0_u15_u5_n101 ) , .ZN( u0_u15_u5_n102 ) , .C2( u0_u15_u5_n115 ) , .C1( u0_u15_u5_n126 ) , .B1( u0_u15_u5_n134 ) , .B2( u0_u15_u5_n160 ) );
  OAI21_X1 u0_u15_u5_U76 (.ZN( u0_u15_u5_n101 ) , .B1( u0_u15_u5_n137 ) , .A( u0_u15_u5_n146 ) , .B2( u0_u15_u5_n147 ) );
  NOR2_X1 u0_u15_u5_U77 (.A2( u0_u15_X_34 ) , .A1( u0_u15_X_35 ) , .ZN( u0_u15_u5_n145 ) );
  NOR2_X1 u0_u15_u5_U78 (.A2( u0_u15_X_34 ) , .ZN( u0_u15_u5_n146 ) , .A1( u0_u15_u5_n171 ) );
  NOR2_X1 u0_u15_u5_U79 (.A2( u0_u15_X_31 ) , .A1( u0_u15_X_32 ) , .ZN( u0_u15_u5_n103 ) );
  NOR3_X1 u0_u15_u5_U8 (.A2( u0_u15_u5_n147 ) , .A1( u0_u15_u5_n148 ) , .ZN( u0_u15_u5_n149 ) , .A3( u0_u15_u5_n194 ) );
  NOR2_X1 u0_u15_u5_U80 (.A2( u0_u15_X_36 ) , .ZN( u0_u15_u5_n105 ) , .A1( u0_u15_u5_n180 ) );
  NOR2_X1 u0_u15_u5_U81 (.A2( u0_u15_X_33 ) , .ZN( u0_u15_u5_n108 ) , .A1( u0_u15_u5_n170 ) );
  NOR2_X1 u0_u15_u5_U82 (.A2( u0_u15_X_33 ) , .A1( u0_u15_X_36 ) , .ZN( u0_u15_u5_n107 ) );
  NOR2_X1 u0_u15_u5_U83 (.A2( u0_u15_X_31 ) , .ZN( u0_u15_u5_n104 ) , .A1( u0_u15_u5_n181 ) );
  NAND2_X1 u0_u15_u5_U84 (.A2( u0_u15_X_34 ) , .A1( u0_u15_X_35 ) , .ZN( u0_u15_u5_n153 ) );
  NAND2_X1 u0_u15_u5_U85 (.A1( u0_u15_X_34 ) , .ZN( u0_u15_u5_n126 ) , .A2( u0_u15_u5_n171 ) );
  AND2_X1 u0_u15_u5_U86 (.A1( u0_u15_X_31 ) , .A2( u0_u15_X_32 ) , .ZN( u0_u15_u5_n106 ) );
  AND2_X1 u0_u15_u5_U87 (.A1( u0_u15_X_31 ) , .ZN( u0_u15_u5_n109 ) , .A2( u0_u15_u5_n181 ) );
  INV_X1 u0_u15_u5_U88 (.A( u0_u15_X_33 ) , .ZN( u0_u15_u5_n180 ) );
  INV_X1 u0_u15_u5_U89 (.A( u0_u15_X_35 ) , .ZN( u0_u15_u5_n171 ) );
  NOR2_X1 u0_u15_u5_U9 (.ZN( u0_u15_u5_n135 ) , .A1( u0_u15_u5_n173 ) , .A2( u0_u15_u5_n176 ) );
  INV_X1 u0_u15_u5_U90 (.A( u0_u15_X_36 ) , .ZN( u0_u15_u5_n170 ) );
  INV_X1 u0_u15_u5_U91 (.A( u0_u15_X_32 ) , .ZN( u0_u15_u5_n181 ) );
  NAND4_X1 u0_u15_u5_U92 (.ZN( u0_out15_19 ) , .A4( u0_u15_u5_n166 ) , .A3( u0_u15_u5_n167 ) , .A2( u0_u15_u5_n168 ) , .A1( u0_u15_u5_n169 ) );
  AOI22_X1 u0_u15_u5_U93 (.B2( u0_u15_u5_n145 ) , .A2( u0_u15_u5_n146 ) , .ZN( u0_u15_u5_n167 ) , .B1( u0_u15_u5_n182 ) , .A1( u0_u15_u5_n189 ) );
  NOR4_X1 u0_u15_u5_U94 (.A4( u0_u15_u5_n162 ) , .A3( u0_u15_u5_n163 ) , .A2( u0_u15_u5_n164 ) , .A1( u0_u15_u5_n165 ) , .ZN( u0_u15_u5_n166 ) );
  NAND4_X1 u0_u15_u5_U95 (.ZN( u0_out15_11 ) , .A4( u0_u15_u5_n143 ) , .A3( u0_u15_u5_n144 ) , .A2( u0_u15_u5_n169 ) , .A1( u0_u15_u5_n196 ) );
  AOI22_X1 u0_u15_u5_U96 (.A2( u0_u15_u5_n132 ) , .ZN( u0_u15_u5_n144 ) , .B2( u0_u15_u5_n145 ) , .B1( u0_u15_u5_n184 ) , .A1( u0_u15_u5_n194 ) );
  NOR3_X1 u0_u15_u5_U97 (.A3( u0_u15_u5_n141 ) , .A1( u0_u15_u5_n142 ) , .ZN( u0_u15_u5_n143 ) , .A2( u0_u15_u5_n191 ) );
  NAND4_X1 u0_u15_u5_U98 (.ZN( u0_out15_4 ) , .A4( u0_u15_u5_n112 ) , .A2( u0_u15_u5_n113 ) , .A1( u0_u15_u5_n114 ) , .A3( u0_u15_u5_n195 ) );
  AOI211_X1 u0_u15_u5_U99 (.A( u0_u15_u5_n110 ) , .C1( u0_u15_u5_n111 ) , .ZN( u0_u15_u5_n112 ) , .B( u0_u15_u5_n118 ) , .C2( u0_u15_u5_n177 ) );
  INV_X1 u0_u15_u6_U10 (.ZN( u0_u15_u6_n172 ) , .A( u0_u15_u6_n88 ) );
  OAI21_X1 u0_u15_u6_U11 (.A( u0_u15_u6_n159 ) , .B1( u0_u15_u6_n169 ) , .B2( u0_u15_u6_n173 ) , .ZN( u0_u15_u6_n90 ) );
  AOI22_X1 u0_u15_u6_U12 (.A2( u0_u15_u6_n151 ) , .B2( u0_u15_u6_n161 ) , .A1( u0_u15_u6_n167 ) , .B1( u0_u15_u6_n170 ) , .ZN( u0_u15_u6_n89 ) );
  AOI21_X1 u0_u15_u6_U13 (.ZN( u0_u15_u6_n106 ) , .A( u0_u15_u6_n142 ) , .B2( u0_u15_u6_n159 ) , .B1( u0_u15_u6_n164 ) );
  INV_X1 u0_u15_u6_U14 (.A( u0_u15_u6_n155 ) , .ZN( u0_u15_u6_n161 ) );
  INV_X1 u0_u15_u6_U15 (.A( u0_u15_u6_n128 ) , .ZN( u0_u15_u6_n164 ) );
  NAND2_X1 u0_u15_u6_U16 (.ZN( u0_u15_u6_n110 ) , .A1( u0_u15_u6_n122 ) , .A2( u0_u15_u6_n129 ) );
  NAND2_X1 u0_u15_u6_U17 (.ZN( u0_u15_u6_n124 ) , .A2( u0_u15_u6_n146 ) , .A1( u0_u15_u6_n148 ) );
  INV_X1 u0_u15_u6_U18 (.A( u0_u15_u6_n132 ) , .ZN( u0_u15_u6_n171 ) );
  AND2_X1 u0_u15_u6_U19 (.A1( u0_u15_u6_n100 ) , .ZN( u0_u15_u6_n130 ) , .A2( u0_u15_u6_n147 ) );
  INV_X1 u0_u15_u6_U20 (.A( u0_u15_u6_n127 ) , .ZN( u0_u15_u6_n173 ) );
  INV_X1 u0_u15_u6_U21 (.A( u0_u15_u6_n121 ) , .ZN( u0_u15_u6_n167 ) );
  INV_X1 u0_u15_u6_U22 (.A( u0_u15_u6_n100 ) , .ZN( u0_u15_u6_n169 ) );
  INV_X1 u0_u15_u6_U23 (.A( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n170 ) );
  INV_X1 u0_u15_u6_U24 (.A( u0_u15_u6_n113 ) , .ZN( u0_u15_u6_n168 ) );
  AND2_X1 u0_u15_u6_U25 (.A1( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n119 ) , .ZN( u0_u15_u6_n133 ) );
  AND2_X1 u0_u15_u6_U26 (.A2( u0_u15_u6_n121 ) , .A1( u0_u15_u6_n122 ) , .ZN( u0_u15_u6_n131 ) );
  AND3_X1 u0_u15_u6_U27 (.ZN( u0_u15_u6_n120 ) , .A2( u0_u15_u6_n127 ) , .A1( u0_u15_u6_n132 ) , .A3( u0_u15_u6_n145 ) );
  INV_X1 u0_u15_u6_U28 (.A( u0_u15_u6_n146 ) , .ZN( u0_u15_u6_n163 ) );
  AOI222_X1 u0_u15_u6_U29 (.ZN( u0_u15_u6_n114 ) , .A1( u0_u15_u6_n118 ) , .A2( u0_u15_u6_n126 ) , .B2( u0_u15_u6_n151 ) , .C2( u0_u15_u6_n159 ) , .C1( u0_u15_u6_n168 ) , .B1( u0_u15_u6_n169 ) );
  INV_X1 u0_u15_u6_U3 (.A( u0_u15_u6_n110 ) , .ZN( u0_u15_u6_n166 ) );
  NOR2_X1 u0_u15_u6_U30 (.A1( u0_u15_u6_n162 ) , .A2( u0_u15_u6_n165 ) , .ZN( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U31 (.A1( u0_u15_u6_n144 ) , .ZN( u0_u15_u6_n151 ) , .A2( u0_u15_u6_n158 ) );
  NAND2_X1 u0_u15_u6_U32 (.ZN( u0_u15_u6_n132 ) , .A1( u0_u15_u6_n91 ) , .A2( u0_u15_u6_n97 ) );
  AOI22_X1 u0_u15_u6_U33 (.B2( u0_u15_u6_n110 ) , .B1( u0_u15_u6_n111 ) , .A1( u0_u15_u6_n112 ) , .ZN( u0_u15_u6_n115 ) , .A2( u0_u15_u6_n161 ) );
  NAND4_X1 u0_u15_u6_U34 (.A3( u0_u15_u6_n109 ) , .ZN( u0_u15_u6_n112 ) , .A4( u0_u15_u6_n132 ) , .A2( u0_u15_u6_n147 ) , .A1( u0_u15_u6_n166 ) );
  NOR2_X1 u0_u15_u6_U35 (.ZN( u0_u15_u6_n109 ) , .A1( u0_u15_u6_n170 ) , .A2( u0_u15_u6_n173 ) );
  NOR2_X1 u0_u15_u6_U36 (.A2( u0_u15_u6_n126 ) , .ZN( u0_u15_u6_n155 ) , .A1( u0_u15_u6_n160 ) );
  NAND2_X1 u0_u15_u6_U37 (.ZN( u0_u15_u6_n146 ) , .A2( u0_u15_u6_n94 ) , .A1( u0_u15_u6_n99 ) );
  AOI21_X1 u0_u15_u6_U38 (.A( u0_u15_u6_n144 ) , .B2( u0_u15_u6_n145 ) , .B1( u0_u15_u6_n146 ) , .ZN( u0_u15_u6_n150 ) );
  AOI211_X1 u0_u15_u6_U39 (.B( u0_u15_u6_n134 ) , .A( u0_u15_u6_n135 ) , .C1( u0_u15_u6_n136 ) , .ZN( u0_u15_u6_n137 ) , .C2( u0_u15_u6_n151 ) );
  INV_X1 u0_u15_u6_U4 (.A( u0_u15_u6_n142 ) , .ZN( u0_u15_u6_n174 ) );
  NAND4_X1 u0_u15_u6_U40 (.A4( u0_u15_u6_n127 ) , .A3( u0_u15_u6_n128 ) , .A2( u0_u15_u6_n129 ) , .A1( u0_u15_u6_n130 ) , .ZN( u0_u15_u6_n136 ) );
  AOI21_X1 u0_u15_u6_U41 (.B2( u0_u15_u6_n132 ) , .B1( u0_u15_u6_n133 ) , .ZN( u0_u15_u6_n134 ) , .A( u0_u15_u6_n158 ) );
  AOI21_X1 u0_u15_u6_U42 (.B1( u0_u15_u6_n131 ) , .ZN( u0_u15_u6_n135 ) , .A( u0_u15_u6_n144 ) , .B2( u0_u15_u6_n146 ) );
  INV_X1 u0_u15_u6_U43 (.A( u0_u15_u6_n111 ) , .ZN( u0_u15_u6_n158 ) );
  NAND2_X1 u0_u15_u6_U44 (.ZN( u0_u15_u6_n127 ) , .A1( u0_u15_u6_n91 ) , .A2( u0_u15_u6_n92 ) );
  NAND2_X1 u0_u15_u6_U45 (.ZN( u0_u15_u6_n129 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n96 ) );
  INV_X1 u0_u15_u6_U46 (.A( u0_u15_u6_n144 ) , .ZN( u0_u15_u6_n159 ) );
  NAND2_X1 u0_u15_u6_U47 (.ZN( u0_u15_u6_n145 ) , .A2( u0_u15_u6_n97 ) , .A1( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U48 (.ZN( u0_u15_u6_n148 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n94 ) );
  NAND2_X1 u0_u15_u6_U49 (.ZN( u0_u15_u6_n108 ) , .A2( u0_u15_u6_n139 ) , .A1( u0_u15_u6_n144 ) );
  NAND2_X1 u0_u15_u6_U5 (.A2( u0_u15_u6_n143 ) , .ZN( u0_u15_u6_n152 ) , .A1( u0_u15_u6_n166 ) );
  NAND2_X1 u0_u15_u6_U50 (.ZN( u0_u15_u6_n121 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n97 ) );
  NAND2_X1 u0_u15_u6_U51 (.ZN( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n95 ) );
  AND2_X1 u0_u15_u6_U52 (.ZN( u0_u15_u6_n118 ) , .A2( u0_u15_u6_n91 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U53 (.ZN( u0_u15_u6_n147 ) , .A2( u0_u15_u6_n98 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U54 (.ZN( u0_u15_u6_n128 ) , .A1( u0_u15_u6_n94 ) , .A2( u0_u15_u6_n96 ) );
  NAND2_X1 u0_u15_u6_U55 (.ZN( u0_u15_u6_n119 ) , .A2( u0_u15_u6_n95 ) , .A1( u0_u15_u6_n99 ) );
  NAND2_X1 u0_u15_u6_U56 (.ZN( u0_u15_u6_n123 ) , .A2( u0_u15_u6_n91 ) , .A1( u0_u15_u6_n96 ) );
  NAND2_X1 u0_u15_u6_U57 (.ZN( u0_u15_u6_n100 ) , .A2( u0_u15_u6_n92 ) , .A1( u0_u15_u6_n98 ) );
  NAND2_X1 u0_u15_u6_U58 (.ZN( u0_u15_u6_n122 ) , .A1( u0_u15_u6_n94 ) , .A2( u0_u15_u6_n97 ) );
  INV_X1 u0_u15_u6_U59 (.A( u0_u15_u6_n139 ) , .ZN( u0_u15_u6_n160 ) );
  AOI22_X1 u0_u15_u6_U6 (.B2( u0_u15_u6_n101 ) , .A1( u0_u15_u6_n102 ) , .ZN( u0_u15_u6_n103 ) , .B1( u0_u15_u6_n160 ) , .A2( u0_u15_u6_n161 ) );
  NAND2_X1 u0_u15_u6_U60 (.ZN( u0_u15_u6_n113 ) , .A1( u0_u15_u6_n96 ) , .A2( u0_u15_u6_n98 ) );
  NOR2_X1 u0_u15_u6_U61 (.A2( u0_u15_X_40 ) , .A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n126 ) );
  NOR2_X1 u0_u15_u6_U62 (.A2( u0_u15_X_39 ) , .A1( u0_u15_X_42 ) , .ZN( u0_u15_u6_n92 ) );
  NOR2_X1 u0_u15_u6_U63 (.A2( u0_u15_X_39 ) , .A1( u0_u15_u6_n156 ) , .ZN( u0_u15_u6_n97 ) );
  NOR2_X1 u0_u15_u6_U64 (.A2( u0_u15_X_38 ) , .A1( u0_u15_u6_n165 ) , .ZN( u0_u15_u6_n95 ) );
  NOR2_X1 u0_u15_u6_U65 (.A2( u0_u15_X_41 ) , .ZN( u0_u15_u6_n111 ) , .A1( u0_u15_u6_n157 ) );
  NOR2_X1 u0_u15_u6_U66 (.A2( u0_u15_X_37 ) , .A1( u0_u15_u6_n162 ) , .ZN( u0_u15_u6_n94 ) );
  NOR2_X1 u0_u15_u6_U67 (.A2( u0_u15_X_37 ) , .A1( u0_u15_X_38 ) , .ZN( u0_u15_u6_n91 ) );
  NAND2_X1 u0_u15_u6_U68 (.A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n144 ) , .A2( u0_u15_u6_n157 ) );
  NAND2_X1 u0_u15_u6_U69 (.A2( u0_u15_X_40 ) , .A1( u0_u15_X_41 ) , .ZN( u0_u15_u6_n139 ) );
  NOR2_X1 u0_u15_u6_U7 (.A1( u0_u15_u6_n118 ) , .ZN( u0_u15_u6_n143 ) , .A2( u0_u15_u6_n168 ) );
  AND2_X1 u0_u15_u6_U70 (.A1( u0_u15_X_39 ) , .A2( u0_u15_u6_n156 ) , .ZN( u0_u15_u6_n96 ) );
  AND2_X1 u0_u15_u6_U71 (.A1( u0_u15_X_39 ) , .A2( u0_u15_X_42 ) , .ZN( u0_u15_u6_n99 ) );
  INV_X1 u0_u15_u6_U72 (.A( u0_u15_X_40 ) , .ZN( u0_u15_u6_n157 ) );
  INV_X1 u0_u15_u6_U73 (.A( u0_u15_X_37 ) , .ZN( u0_u15_u6_n165 ) );
  INV_X1 u0_u15_u6_U74 (.A( u0_u15_X_38 ) , .ZN( u0_u15_u6_n162 ) );
  INV_X1 u0_u15_u6_U75 (.A( u0_u15_X_42 ) , .ZN( u0_u15_u6_n156 ) );
  NAND4_X1 u0_u15_u6_U76 (.ZN( u0_out15_12 ) , .A4( u0_u15_u6_n114 ) , .A3( u0_u15_u6_n115 ) , .A2( u0_u15_u6_n116 ) , .A1( u0_u15_u6_n117 ) );
  OAI22_X1 u0_u15_u6_U77 (.B2( u0_u15_u6_n111 ) , .ZN( u0_u15_u6_n116 ) , .B1( u0_u15_u6_n126 ) , .A2( u0_u15_u6_n164 ) , .A1( u0_u15_u6_n167 ) );
  OAI21_X1 u0_u15_u6_U78 (.A( u0_u15_u6_n108 ) , .ZN( u0_u15_u6_n117 ) , .B2( u0_u15_u6_n141 ) , .B1( u0_u15_u6_n163 ) );
  NAND4_X1 u0_u15_u6_U79 (.ZN( u0_out15_32 ) , .A4( u0_u15_u6_n103 ) , .A3( u0_u15_u6_n104 ) , .A2( u0_u15_u6_n105 ) , .A1( u0_u15_u6_n106 ) );
  AOI21_X1 u0_u15_u6_U8 (.B1( u0_u15_u6_n107 ) , .B2( u0_u15_u6_n132 ) , .A( u0_u15_u6_n158 ) , .ZN( u0_u15_u6_n88 ) );
  AOI22_X1 u0_u15_u6_U80 (.ZN( u0_u15_u6_n105 ) , .A2( u0_u15_u6_n108 ) , .A1( u0_u15_u6_n118 ) , .B2( u0_u15_u6_n126 ) , .B1( u0_u15_u6_n171 ) );
  AOI22_X1 u0_u15_u6_U81 (.ZN( u0_u15_u6_n104 ) , .A1( u0_u15_u6_n111 ) , .B1( u0_u15_u6_n124 ) , .B2( u0_u15_u6_n151 ) , .A2( u0_u15_u6_n93 ) );
  OAI211_X1 u0_u15_u6_U82 (.ZN( u0_out15_22 ) , .B( u0_u15_u6_n137 ) , .A( u0_u15_u6_n138 ) , .C2( u0_u15_u6_n139 ) , .C1( u0_u15_u6_n140 ) );
  AOI22_X1 u0_u15_u6_U83 (.B1( u0_u15_u6_n124 ) , .A2( u0_u15_u6_n125 ) , .A1( u0_u15_u6_n126 ) , .ZN( u0_u15_u6_n138 ) , .B2( u0_u15_u6_n161 ) );
  AND4_X1 u0_u15_u6_U84 (.A3( u0_u15_u6_n119 ) , .A1( u0_u15_u6_n120 ) , .A4( u0_u15_u6_n129 ) , .ZN( u0_u15_u6_n140 ) , .A2( u0_u15_u6_n143 ) );
  OAI211_X1 u0_u15_u6_U85 (.ZN( u0_out15_7 ) , .B( u0_u15_u6_n153 ) , .C2( u0_u15_u6_n154 ) , .C1( u0_u15_u6_n155 ) , .A( u0_u15_u6_n174 ) );
  NOR3_X1 u0_u15_u6_U86 (.A1( u0_u15_u6_n141 ) , .ZN( u0_u15_u6_n154 ) , .A3( u0_u15_u6_n164 ) , .A2( u0_u15_u6_n171 ) );
  AOI211_X1 u0_u15_u6_U87 (.B( u0_u15_u6_n149 ) , .A( u0_u15_u6_n150 ) , .C2( u0_u15_u6_n151 ) , .C1( u0_u15_u6_n152 ) , .ZN( u0_u15_u6_n153 ) );
  NAND3_X1 u0_u15_u6_U88 (.A2( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n125 ) , .A1( u0_u15_u6_n130 ) , .A3( u0_u15_u6_n131 ) );
  NAND3_X1 u0_u15_u6_U89 (.A3( u0_u15_u6_n133 ) , .ZN( u0_u15_u6_n141 ) , .A1( u0_u15_u6_n145 ) , .A2( u0_u15_u6_n148 ) );
  AOI21_X1 u0_u15_u6_U9 (.B2( u0_u15_u6_n147 ) , .B1( u0_u15_u6_n148 ) , .ZN( u0_u15_u6_n149 ) , .A( u0_u15_u6_n158 ) );
  NAND3_X1 u0_u15_u6_U90 (.ZN( u0_u15_u6_n101 ) , .A3( u0_u15_u6_n107 ) , .A2( u0_u15_u6_n121 ) , .A1( u0_u15_u6_n127 ) );
  NAND3_X1 u0_u15_u6_U91 (.ZN( u0_u15_u6_n102 ) , .A3( u0_u15_u6_n130 ) , .A2( u0_u15_u6_n145 ) , .A1( u0_u15_u6_n166 ) );
  NAND3_X1 u0_u15_u6_U92 (.A3( u0_u15_u6_n113 ) , .A1( u0_u15_u6_n119 ) , .A2( u0_u15_u6_n123 ) , .ZN( u0_u15_u6_n93 ) );
  NAND3_X1 u0_u15_u6_U93 (.ZN( u0_u15_u6_n142 ) , .A2( u0_u15_u6_n172 ) , .A3( u0_u15_u6_n89 ) , .A1( u0_u15_u6_n90 ) );
  OAI21_X1 u0_u15_u7_U10 (.A( u0_u15_u7_n161 ) , .B1( u0_u15_u7_n168 ) , .B2( u0_u15_u7_n173 ) , .ZN( u0_u15_u7_n91 ) );
  AOI211_X1 u0_u15_u7_U11 (.A( u0_u15_u7_n117 ) , .ZN( u0_u15_u7_n118 ) , .C2( u0_u15_u7_n126 ) , .C1( u0_u15_u7_n177 ) , .B( u0_u15_u7_n180 ) );
  OAI22_X1 u0_u15_u7_U12 (.B1( u0_u15_u7_n115 ) , .ZN( u0_u15_u7_n117 ) , .A2( u0_u15_u7_n133 ) , .A1( u0_u15_u7_n137 ) , .B2( u0_u15_u7_n162 ) );
  INV_X1 u0_u15_u7_U13 (.A( u0_u15_u7_n116 ) , .ZN( u0_u15_u7_n180 ) );
  NOR3_X1 u0_u15_u7_U14 (.ZN( u0_u15_u7_n115 ) , .A3( u0_u15_u7_n145 ) , .A2( u0_u15_u7_n168 ) , .A1( u0_u15_u7_n169 ) );
  OAI211_X1 u0_u15_u7_U15 (.B( u0_u15_u7_n122 ) , .A( u0_u15_u7_n123 ) , .C2( u0_u15_u7_n124 ) , .ZN( u0_u15_u7_n154 ) , .C1( u0_u15_u7_n162 ) );
  AOI222_X1 u0_u15_u7_U16 (.ZN( u0_u15_u7_n122 ) , .C2( u0_u15_u7_n126 ) , .C1( u0_u15_u7_n145 ) , .B1( u0_u15_u7_n161 ) , .A2( u0_u15_u7_n165 ) , .B2( u0_u15_u7_n170 ) , .A1( u0_u15_u7_n176 ) );
  INV_X1 u0_u15_u7_U17 (.A( u0_u15_u7_n133 ) , .ZN( u0_u15_u7_n176 ) );
  NOR3_X1 u0_u15_u7_U18 (.A2( u0_u15_u7_n134 ) , .A1( u0_u15_u7_n135 ) , .ZN( u0_u15_u7_n136 ) , .A3( u0_u15_u7_n171 ) );
  NOR2_X1 u0_u15_u7_U19 (.A1( u0_u15_u7_n130 ) , .A2( u0_u15_u7_n134 ) , .ZN( u0_u15_u7_n153 ) );
  INV_X1 u0_u15_u7_U20 (.A( u0_u15_u7_n101 ) , .ZN( u0_u15_u7_n165 ) );
  NOR2_X1 u0_u15_u7_U21 (.ZN( u0_u15_u7_n111 ) , .A2( u0_u15_u7_n134 ) , .A1( u0_u15_u7_n169 ) );
  AOI21_X1 u0_u15_u7_U22 (.ZN( u0_u15_u7_n104 ) , .B2( u0_u15_u7_n112 ) , .B1( u0_u15_u7_n127 ) , .A( u0_u15_u7_n164 ) );
  AOI21_X1 u0_u15_u7_U23 (.ZN( u0_u15_u7_n106 ) , .B1( u0_u15_u7_n133 ) , .B2( u0_u15_u7_n146 ) , .A( u0_u15_u7_n162 ) );
  AOI21_X1 u0_u15_u7_U24 (.A( u0_u15_u7_n101 ) , .ZN( u0_u15_u7_n107 ) , .B2( u0_u15_u7_n128 ) , .B1( u0_u15_u7_n175 ) );
  INV_X1 u0_u15_u7_U25 (.A( u0_u15_u7_n138 ) , .ZN( u0_u15_u7_n171 ) );
  INV_X1 u0_u15_u7_U26 (.A( u0_u15_u7_n131 ) , .ZN( u0_u15_u7_n177 ) );
  INV_X1 u0_u15_u7_U27 (.A( u0_u15_u7_n110 ) , .ZN( u0_u15_u7_n174 ) );
  NAND2_X1 u0_u15_u7_U28 (.A1( u0_u15_u7_n129 ) , .A2( u0_u15_u7_n132 ) , .ZN( u0_u15_u7_n149 ) );
  NAND2_X1 u0_u15_u7_U29 (.A1( u0_u15_u7_n113 ) , .A2( u0_u15_u7_n124 ) , .ZN( u0_u15_u7_n130 ) );
  INV_X1 u0_u15_u7_U3 (.A( u0_u15_u7_n111 ) , .ZN( u0_u15_u7_n170 ) );
  INV_X1 u0_u15_u7_U30 (.A( u0_u15_u7_n112 ) , .ZN( u0_u15_u7_n173 ) );
  INV_X1 u0_u15_u7_U31 (.A( u0_u15_u7_n128 ) , .ZN( u0_u15_u7_n168 ) );
  INV_X1 u0_u15_u7_U32 (.A( u0_u15_u7_n148 ) , .ZN( u0_u15_u7_n169 ) );
  INV_X1 u0_u15_u7_U33 (.A( u0_u15_u7_n127 ) , .ZN( u0_u15_u7_n179 ) );
  NOR2_X1 u0_u15_u7_U34 (.ZN( u0_u15_u7_n101 ) , .A2( u0_u15_u7_n150 ) , .A1( u0_u15_u7_n156 ) );
  AOI211_X1 u0_u15_u7_U35 (.B( u0_u15_u7_n154 ) , .A( u0_u15_u7_n155 ) , .C1( u0_u15_u7_n156 ) , .ZN( u0_u15_u7_n157 ) , .C2( u0_u15_u7_n172 ) );
  INV_X1 u0_u15_u7_U36 (.A( u0_u15_u7_n153 ) , .ZN( u0_u15_u7_n172 ) );
  AOI211_X1 u0_u15_u7_U37 (.B( u0_u15_u7_n139 ) , .A( u0_u15_u7_n140 ) , .C2( u0_u15_u7_n141 ) , .ZN( u0_u15_u7_n142 ) , .C1( u0_u15_u7_n156 ) );
  NAND4_X1 u0_u15_u7_U38 (.A3( u0_u15_u7_n127 ) , .A2( u0_u15_u7_n128 ) , .A1( u0_u15_u7_n129 ) , .ZN( u0_u15_u7_n141 ) , .A4( u0_u15_u7_n147 ) );
  AOI21_X1 u0_u15_u7_U39 (.A( u0_u15_u7_n137 ) , .B1( u0_u15_u7_n138 ) , .ZN( u0_u15_u7_n139 ) , .B2( u0_u15_u7_n146 ) );
  INV_X1 u0_u15_u7_U4 (.A( u0_u15_u7_n149 ) , .ZN( u0_u15_u7_n175 ) );
  OAI22_X1 u0_u15_u7_U40 (.B1( u0_u15_u7_n136 ) , .ZN( u0_u15_u7_n140 ) , .A1( u0_u15_u7_n153 ) , .B2( u0_u15_u7_n162 ) , .A2( u0_u15_u7_n164 ) );
  AOI21_X1 u0_u15_u7_U41 (.ZN( u0_u15_u7_n123 ) , .B1( u0_u15_u7_n165 ) , .B2( u0_u15_u7_n177 ) , .A( u0_u15_u7_n97 ) );
  AOI21_X1 u0_u15_u7_U42 (.B2( u0_u15_u7_n113 ) , .B1( u0_u15_u7_n124 ) , .A( u0_u15_u7_n125 ) , .ZN( u0_u15_u7_n97 ) );
  INV_X1 u0_u15_u7_U43 (.A( u0_u15_u7_n125 ) , .ZN( u0_u15_u7_n161 ) );
  INV_X1 u0_u15_u7_U44 (.A( u0_u15_u7_n152 ) , .ZN( u0_u15_u7_n162 ) );
  AOI22_X1 u0_u15_u7_U45 (.A2( u0_u15_u7_n114 ) , .ZN( u0_u15_u7_n119 ) , .B1( u0_u15_u7_n130 ) , .A1( u0_u15_u7_n156 ) , .B2( u0_u15_u7_n165 ) );
  NAND2_X1 u0_u15_u7_U46 (.A2( u0_u15_u7_n112 ) , .ZN( u0_u15_u7_n114 ) , .A1( u0_u15_u7_n175 ) );
  AOI22_X1 u0_u15_u7_U47 (.B2( u0_u15_u7_n149 ) , .B1( u0_u15_u7_n150 ) , .A2( u0_u15_u7_n151 ) , .A1( u0_u15_u7_n152 ) , .ZN( u0_u15_u7_n158 ) );
  AND2_X1 u0_u15_u7_U48 (.ZN( u0_u15_u7_n145 ) , .A2( u0_u15_u7_n98 ) , .A1( u0_u15_u7_n99 ) );
  NOR2_X1 u0_u15_u7_U49 (.ZN( u0_u15_u7_n137 ) , .A1( u0_u15_u7_n150 ) , .A2( u0_u15_u7_n161 ) );
  INV_X1 u0_u15_u7_U5 (.A( u0_u15_u7_n154 ) , .ZN( u0_u15_u7_n178 ) );
  AOI21_X1 u0_u15_u7_U50 (.ZN( u0_u15_u7_n105 ) , .B2( u0_u15_u7_n110 ) , .A( u0_u15_u7_n125 ) , .B1( u0_u15_u7_n147 ) );
  NAND2_X1 u0_u15_u7_U51 (.ZN( u0_u15_u7_n146 ) , .A1( u0_u15_u7_n95 ) , .A2( u0_u15_u7_n98 ) );
  NAND2_X1 u0_u15_u7_U52 (.A2( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n147 ) , .A1( u0_u15_u7_n93 ) );
  NAND2_X1 u0_u15_u7_U53 (.A1( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n127 ) , .A2( u0_u15_u7_n99 ) );
  OR2_X1 u0_u15_u7_U54 (.ZN( u0_u15_u7_n126 ) , .A2( u0_u15_u7_n152 ) , .A1( u0_u15_u7_n156 ) );
  NAND2_X1 u0_u15_u7_U55 (.A2( u0_u15_u7_n102 ) , .A1( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n133 ) );
  NAND2_X1 u0_u15_u7_U56 (.ZN( u0_u15_u7_n112 ) , .A2( u0_u15_u7_n96 ) , .A1( u0_u15_u7_n99 ) );
  NAND2_X1 u0_u15_u7_U57 (.A2( u0_u15_u7_n102 ) , .ZN( u0_u15_u7_n128 ) , .A1( u0_u15_u7_n98 ) );
  NAND2_X1 u0_u15_u7_U58 (.A1( u0_u15_u7_n100 ) , .ZN( u0_u15_u7_n113 ) , .A2( u0_u15_u7_n93 ) );
  NAND2_X1 u0_u15_u7_U59 (.A2( u0_u15_u7_n102 ) , .ZN( u0_u15_u7_n124 ) , .A1( u0_u15_u7_n96 ) );
  AOI211_X1 u0_u15_u7_U6 (.ZN( u0_u15_u7_n116 ) , .A( u0_u15_u7_n155 ) , .C1( u0_u15_u7_n161 ) , .C2( u0_u15_u7_n171 ) , .B( u0_u15_u7_n94 ) );
  NAND2_X1 u0_u15_u7_U60 (.ZN( u0_u15_u7_n110 ) , .A1( u0_u15_u7_n95 ) , .A2( u0_u15_u7_n96 ) );
  INV_X1 u0_u15_u7_U61 (.A( u0_u15_u7_n150 ) , .ZN( u0_u15_u7_n164 ) );
  AND2_X1 u0_u15_u7_U62 (.ZN( u0_u15_u7_n134 ) , .A1( u0_u15_u7_n93 ) , .A2( u0_u15_u7_n98 ) );
  NAND2_X1 u0_u15_u7_U63 (.A1( u0_u15_u7_n100 ) , .A2( u0_u15_u7_n102 ) , .ZN( u0_u15_u7_n129 ) );
  NAND2_X1 u0_u15_u7_U64 (.A2( u0_u15_u7_n103 ) , .ZN( u0_u15_u7_n131 ) , .A1( u0_u15_u7_n95 ) );
  NAND2_X1 u0_u15_u7_U65 (.A1( u0_u15_u7_n100 ) , .ZN( u0_u15_u7_n138 ) , .A2( u0_u15_u7_n99 ) );
  NAND2_X1 u0_u15_u7_U66 (.ZN( u0_u15_u7_n132 ) , .A1( u0_u15_u7_n93 ) , .A2( u0_u15_u7_n96 ) );
  NAND2_X1 u0_u15_u7_U67 (.A1( u0_u15_u7_n100 ) , .ZN( u0_u15_u7_n148 ) , .A2( u0_u15_u7_n95 ) );
  NOR2_X1 u0_u15_u7_U68 (.A2( u0_u15_X_47 ) , .ZN( u0_u15_u7_n150 ) , .A1( u0_u15_u7_n163 ) );
  NOR2_X1 u0_u15_u7_U69 (.A2( u0_u15_X_43 ) , .A1( u0_u15_X_44 ) , .ZN( u0_u15_u7_n103 ) );
  OAI222_X1 u0_u15_u7_U7 (.C2( u0_u15_u7_n101 ) , .B2( u0_u15_u7_n111 ) , .A1( u0_u15_u7_n113 ) , .C1( u0_u15_u7_n146 ) , .A2( u0_u15_u7_n162 ) , .B1( u0_u15_u7_n164 ) , .ZN( u0_u15_u7_n94 ) );
  NOR2_X1 u0_u15_u7_U70 (.A2( u0_u15_X_48 ) , .A1( u0_u15_u7_n166 ) , .ZN( u0_u15_u7_n95 ) );
  NOR2_X1 u0_u15_u7_U71 (.A2( u0_u15_X_45 ) , .A1( u0_u15_X_48 ) , .ZN( u0_u15_u7_n99 ) );
  NOR2_X1 u0_u15_u7_U72 (.A2( u0_u15_X_44 ) , .A1( u0_u15_u7_n167 ) , .ZN( u0_u15_u7_n98 ) );
  NOR2_X1 u0_u15_u7_U73 (.A2( u0_u15_X_46 ) , .A1( u0_u15_X_47 ) , .ZN( u0_u15_u7_n152 ) );
  AND2_X1 u0_u15_u7_U74 (.A1( u0_u15_X_47 ) , .ZN( u0_u15_u7_n156 ) , .A2( u0_u15_u7_n163 ) );
  NAND2_X1 u0_u15_u7_U75 (.A2( u0_u15_X_46 ) , .A1( u0_u15_X_47 ) , .ZN( u0_u15_u7_n125 ) );
  AND2_X1 u0_u15_u7_U76 (.A2( u0_u15_X_45 ) , .A1( u0_u15_X_48 ) , .ZN( u0_u15_u7_n102 ) );
  AND2_X1 u0_u15_u7_U77 (.A2( u0_u15_X_43 ) , .A1( u0_u15_X_44 ) , .ZN( u0_u15_u7_n96 ) );
  AND2_X1 u0_u15_u7_U78 (.A1( u0_u15_X_44 ) , .ZN( u0_u15_u7_n100 ) , .A2( u0_u15_u7_n167 ) );
  AND2_X1 u0_u15_u7_U79 (.A1( u0_u15_X_48 ) , .A2( u0_u15_u7_n166 ) , .ZN( u0_u15_u7_n93 ) );
  OAI221_X1 u0_u15_u7_U8 (.C1( u0_u15_u7_n101 ) , .C2( u0_u15_u7_n147 ) , .ZN( u0_u15_u7_n155 ) , .B2( u0_u15_u7_n162 ) , .A( u0_u15_u7_n91 ) , .B1( u0_u15_u7_n92 ) );
  INV_X1 u0_u15_u7_U80 (.A( u0_u15_X_46 ) , .ZN( u0_u15_u7_n163 ) );
  INV_X1 u0_u15_u7_U81 (.A( u0_u15_X_45 ) , .ZN( u0_u15_u7_n166 ) );
  INV_X1 u0_u15_u7_U82 (.A( u0_u15_X_43 ) , .ZN( u0_u15_u7_n167 ) );
  NAND4_X1 u0_u15_u7_U83 (.ZN( u0_out15_5 ) , .A4( u0_u15_u7_n108 ) , .A3( u0_u15_u7_n109 ) , .A1( u0_u15_u7_n116 ) , .A2( u0_u15_u7_n123 ) );
  AOI22_X1 u0_u15_u7_U84 (.ZN( u0_u15_u7_n109 ) , .A2( u0_u15_u7_n126 ) , .B2( u0_u15_u7_n145 ) , .B1( u0_u15_u7_n156 ) , .A1( u0_u15_u7_n171 ) );
  NOR4_X1 u0_u15_u7_U85 (.A4( u0_u15_u7_n104 ) , .A3( u0_u15_u7_n105 ) , .A2( u0_u15_u7_n106 ) , .A1( u0_u15_u7_n107 ) , .ZN( u0_u15_u7_n108 ) );
  NAND4_X1 u0_u15_u7_U86 (.ZN( u0_out15_21 ) , .A4( u0_u15_u7_n157 ) , .A3( u0_u15_u7_n158 ) , .A2( u0_u15_u7_n159 ) , .A1( u0_u15_u7_n160 ) );
  OAI21_X1 u0_u15_u7_U87 (.B1( u0_u15_u7_n145 ) , .ZN( u0_u15_u7_n160 ) , .A( u0_u15_u7_n161 ) , .B2( u0_u15_u7_n177 ) );
  OAI21_X1 u0_u15_u7_U88 (.ZN( u0_u15_u7_n159 ) , .A( u0_u15_u7_n165 ) , .B2( u0_u15_u7_n171 ) , .B1( u0_u15_u7_n174 ) );
  NAND4_X1 u0_u15_u7_U89 (.ZN( u0_out15_15 ) , .A4( u0_u15_u7_n142 ) , .A3( u0_u15_u7_n143 ) , .A2( u0_u15_u7_n144 ) , .A1( u0_u15_u7_n178 ) );
  AND3_X1 u0_u15_u7_U9 (.A3( u0_u15_u7_n110 ) , .A2( u0_u15_u7_n127 ) , .A1( u0_u15_u7_n132 ) , .ZN( u0_u15_u7_n92 ) );
  OR2_X1 u0_u15_u7_U90 (.A2( u0_u15_u7_n125 ) , .A1( u0_u15_u7_n129 ) , .ZN( u0_u15_u7_n144 ) );
  AOI22_X1 u0_u15_u7_U91 (.A2( u0_u15_u7_n126 ) , .ZN( u0_u15_u7_n143 ) , .B2( u0_u15_u7_n165 ) , .B1( u0_u15_u7_n173 ) , .A1( u0_u15_u7_n174 ) );
  NAND4_X1 u0_u15_u7_U92 (.ZN( u0_out15_27 ) , .A4( u0_u15_u7_n118 ) , .A3( u0_u15_u7_n119 ) , .A2( u0_u15_u7_n120 ) , .A1( u0_u15_u7_n121 ) );
  OAI21_X1 u0_u15_u7_U93 (.ZN( u0_u15_u7_n121 ) , .B2( u0_u15_u7_n145 ) , .A( u0_u15_u7_n150 ) , .B1( u0_u15_u7_n174 ) );
  OAI21_X1 u0_u15_u7_U94 (.ZN( u0_u15_u7_n120 ) , .A( u0_u15_u7_n161 ) , .B2( u0_u15_u7_n170 ) , .B1( u0_u15_u7_n179 ) );
  NAND3_X1 u0_u15_u7_U95 (.A3( u0_u15_u7_n146 ) , .A2( u0_u15_u7_n147 ) , .A1( u0_u15_u7_n148 ) , .ZN( u0_u15_u7_n151 ) );
  NAND3_X1 u0_u15_u7_U96 (.A3( u0_u15_u7_n131 ) , .A2( u0_u15_u7_n132 ) , .A1( u0_u15_u7_n133 ) , .ZN( u0_u15_u7_n135 ) );
  XOR2_X1 u0_u1_U10 (.B( u0_K2_45 ) , .A( u0_R0_30 ) , .Z( u0_u1_X_45 ) );
  XOR2_X1 u0_u1_U11 (.B( u0_K2_44 ) , .A( u0_R0_29 ) , .Z( u0_u1_X_44 ) );
  XOR2_X1 u0_u1_U12 (.B( u0_K2_43 ) , .A( u0_R0_28 ) , .Z( u0_u1_X_43 ) );
  XOR2_X1 u0_u1_U7 (.B( u0_K2_48 ) , .A( u0_R0_1 ) , .Z( u0_u1_X_48 ) );
  XOR2_X1 u0_u1_U8 (.B( u0_K2_47 ) , .A( u0_R0_32 ) , .Z( u0_u1_X_47 ) );
  XOR2_X1 u0_u1_U9 (.B( u0_K2_46 ) , .A( u0_R0_31 ) , .Z( u0_u1_X_46 ) );
  AND3_X1 u0_u1_u7_U10 (.A3( u0_u1_u7_n110 ) , .A2( u0_u1_u7_n127 ) , .A1( u0_u1_u7_n132 ) , .ZN( u0_u1_u7_n92 ) );
  OAI21_X1 u0_u1_u7_U11 (.A( u0_u1_u7_n161 ) , .B1( u0_u1_u7_n168 ) , .B2( u0_u1_u7_n173 ) , .ZN( u0_u1_u7_n91 ) );
  AOI211_X1 u0_u1_u7_U12 (.A( u0_u1_u7_n117 ) , .ZN( u0_u1_u7_n118 ) , .C2( u0_u1_u7_n126 ) , .C1( u0_u1_u7_n177 ) , .B( u0_u1_u7_n180 ) );
  OAI22_X1 u0_u1_u7_U13 (.B1( u0_u1_u7_n115 ) , .ZN( u0_u1_u7_n117 ) , .A2( u0_u1_u7_n133 ) , .A1( u0_u1_u7_n137 ) , .B2( u0_u1_u7_n162 ) );
  INV_X1 u0_u1_u7_U14 (.A( u0_u1_u7_n116 ) , .ZN( u0_u1_u7_n180 ) );
  NOR3_X1 u0_u1_u7_U15 (.ZN( u0_u1_u7_n115 ) , .A3( u0_u1_u7_n145 ) , .A2( u0_u1_u7_n168 ) , .A1( u0_u1_u7_n169 ) );
  OAI211_X1 u0_u1_u7_U16 (.B( u0_u1_u7_n122 ) , .A( u0_u1_u7_n123 ) , .C2( u0_u1_u7_n124 ) , .ZN( u0_u1_u7_n154 ) , .C1( u0_u1_u7_n162 ) );
  AOI222_X1 u0_u1_u7_U17 (.ZN( u0_u1_u7_n122 ) , .C2( u0_u1_u7_n126 ) , .C1( u0_u1_u7_n145 ) , .B1( u0_u1_u7_n161 ) , .A2( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n170 ) , .A1( u0_u1_u7_n176 ) );
  INV_X1 u0_u1_u7_U18 (.A( u0_u1_u7_n133 ) , .ZN( u0_u1_u7_n176 ) );
  NOR3_X1 u0_u1_u7_U19 (.A2( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n135 ) , .ZN( u0_u1_u7_n136 ) , .A3( u0_u1_u7_n171 ) );
  NOR2_X1 u0_u1_u7_U20 (.A1( u0_u1_u7_n130 ) , .A2( u0_u1_u7_n134 ) , .ZN( u0_u1_u7_n153 ) );
  INV_X1 u0_u1_u7_U21 (.A( u0_u1_u7_n101 ) , .ZN( u0_u1_u7_n165 ) );
  NOR2_X1 u0_u1_u7_U22 (.ZN( u0_u1_u7_n111 ) , .A2( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n169 ) );
  AOI21_X1 u0_u1_u7_U23 (.ZN( u0_u1_u7_n104 ) , .B2( u0_u1_u7_n112 ) , .B1( u0_u1_u7_n127 ) , .A( u0_u1_u7_n164 ) );
  AOI21_X1 u0_u1_u7_U24 (.ZN( u0_u1_u7_n106 ) , .B1( u0_u1_u7_n133 ) , .B2( u0_u1_u7_n146 ) , .A( u0_u1_u7_n162 ) );
  AOI21_X1 u0_u1_u7_U25 (.A( u0_u1_u7_n101 ) , .ZN( u0_u1_u7_n107 ) , .B2( u0_u1_u7_n128 ) , .B1( u0_u1_u7_n175 ) );
  INV_X1 u0_u1_u7_U26 (.A( u0_u1_u7_n138 ) , .ZN( u0_u1_u7_n171 ) );
  INV_X1 u0_u1_u7_U27 (.A( u0_u1_u7_n131 ) , .ZN( u0_u1_u7_n177 ) );
  INV_X1 u0_u1_u7_U28 (.A( u0_u1_u7_n110 ) , .ZN( u0_u1_u7_n174 ) );
  NAND2_X1 u0_u1_u7_U29 (.A1( u0_u1_u7_n129 ) , .A2( u0_u1_u7_n132 ) , .ZN( u0_u1_u7_n149 ) );
  OAI21_X1 u0_u1_u7_U3 (.ZN( u0_u1_u7_n159 ) , .A( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n171 ) , .B1( u0_u1_u7_n174 ) );
  NAND2_X1 u0_u1_u7_U30 (.A1( u0_u1_u7_n113 ) , .A2( u0_u1_u7_n124 ) , .ZN( u0_u1_u7_n130 ) );
  INV_X1 u0_u1_u7_U31 (.A( u0_u1_u7_n112 ) , .ZN( u0_u1_u7_n173 ) );
  INV_X1 u0_u1_u7_U32 (.A( u0_u1_u7_n128 ) , .ZN( u0_u1_u7_n168 ) );
  INV_X1 u0_u1_u7_U33 (.A( u0_u1_u7_n148 ) , .ZN( u0_u1_u7_n169 ) );
  INV_X1 u0_u1_u7_U34 (.A( u0_u1_u7_n127 ) , .ZN( u0_u1_u7_n179 ) );
  NOR2_X1 u0_u1_u7_U35 (.ZN( u0_u1_u7_n101 ) , .A2( u0_u1_u7_n150 ) , .A1( u0_u1_u7_n156 ) );
  AOI211_X1 u0_u1_u7_U36 (.B( u0_u1_u7_n154 ) , .A( u0_u1_u7_n155 ) , .C1( u0_u1_u7_n156 ) , .ZN( u0_u1_u7_n157 ) , .C2( u0_u1_u7_n172 ) );
  INV_X1 u0_u1_u7_U37 (.A( u0_u1_u7_n153 ) , .ZN( u0_u1_u7_n172 ) );
  AOI211_X1 u0_u1_u7_U38 (.B( u0_u1_u7_n139 ) , .A( u0_u1_u7_n140 ) , .C2( u0_u1_u7_n141 ) , .ZN( u0_u1_u7_n142 ) , .C1( u0_u1_u7_n156 ) );
  NAND4_X1 u0_u1_u7_U39 (.A3( u0_u1_u7_n127 ) , .A2( u0_u1_u7_n128 ) , .A1( u0_u1_u7_n129 ) , .ZN( u0_u1_u7_n141 ) , .A4( u0_u1_u7_n147 ) );
  INV_X1 u0_u1_u7_U4 (.A( u0_u1_u7_n111 ) , .ZN( u0_u1_u7_n170 ) );
  AOI21_X1 u0_u1_u7_U40 (.A( u0_u1_u7_n137 ) , .B1( u0_u1_u7_n138 ) , .ZN( u0_u1_u7_n139 ) , .B2( u0_u1_u7_n146 ) );
  OAI22_X1 u0_u1_u7_U41 (.B1( u0_u1_u7_n136 ) , .ZN( u0_u1_u7_n140 ) , .A1( u0_u1_u7_n153 ) , .B2( u0_u1_u7_n162 ) , .A2( u0_u1_u7_n164 ) );
  AOI21_X1 u0_u1_u7_U42 (.ZN( u0_u1_u7_n123 ) , .B1( u0_u1_u7_n165 ) , .B2( u0_u1_u7_n177 ) , .A( u0_u1_u7_n97 ) );
  AOI21_X1 u0_u1_u7_U43 (.B2( u0_u1_u7_n113 ) , .B1( u0_u1_u7_n124 ) , .A( u0_u1_u7_n125 ) , .ZN( u0_u1_u7_n97 ) );
  INV_X1 u0_u1_u7_U44 (.A( u0_u1_u7_n125 ) , .ZN( u0_u1_u7_n161 ) );
  INV_X1 u0_u1_u7_U45 (.A( u0_u1_u7_n152 ) , .ZN( u0_u1_u7_n162 ) );
  AOI22_X1 u0_u1_u7_U46 (.A2( u0_u1_u7_n114 ) , .ZN( u0_u1_u7_n119 ) , .B1( u0_u1_u7_n130 ) , .A1( u0_u1_u7_n156 ) , .B2( u0_u1_u7_n165 ) );
  NAND2_X1 u0_u1_u7_U47 (.A2( u0_u1_u7_n112 ) , .ZN( u0_u1_u7_n114 ) , .A1( u0_u1_u7_n175 ) );
  AND2_X1 u0_u1_u7_U48 (.ZN( u0_u1_u7_n145 ) , .A2( u0_u1_u7_n98 ) , .A1( u0_u1_u7_n99 ) );
  NOR2_X1 u0_u1_u7_U49 (.ZN( u0_u1_u7_n137 ) , .A1( u0_u1_u7_n150 ) , .A2( u0_u1_u7_n161 ) );
  INV_X1 u0_u1_u7_U5 (.A( u0_u1_u7_n149 ) , .ZN( u0_u1_u7_n175 ) );
  AOI21_X1 u0_u1_u7_U50 (.ZN( u0_u1_u7_n105 ) , .B2( u0_u1_u7_n110 ) , .A( u0_u1_u7_n125 ) , .B1( u0_u1_u7_n147 ) );
  NAND2_X1 u0_u1_u7_U51 (.ZN( u0_u1_u7_n146 ) , .A1( u0_u1_u7_n95 ) , .A2( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U52 (.A2( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n147 ) , .A1( u0_u1_u7_n93 ) );
  NAND2_X1 u0_u1_u7_U53 (.A1( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n127 ) , .A2( u0_u1_u7_n99 ) );
  OR2_X1 u0_u1_u7_U54 (.ZN( u0_u1_u7_n126 ) , .A2( u0_u1_u7_n152 ) , .A1( u0_u1_u7_n156 ) );
  NAND2_X1 u0_u1_u7_U55 (.A2( u0_u1_u7_n102 ) , .A1( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n133 ) );
  NAND2_X1 u0_u1_u7_U56 (.ZN( u0_u1_u7_n112 ) , .A2( u0_u1_u7_n96 ) , .A1( u0_u1_u7_n99 ) );
  NAND2_X1 u0_u1_u7_U57 (.A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n128 ) , .A1( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U58 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n113 ) , .A2( u0_u1_u7_n93 ) );
  NAND2_X1 u0_u1_u7_U59 (.A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n124 ) , .A1( u0_u1_u7_n96 ) );
  INV_X1 u0_u1_u7_U6 (.A( u0_u1_u7_n154 ) , .ZN( u0_u1_u7_n178 ) );
  NAND2_X1 u0_u1_u7_U60 (.ZN( u0_u1_u7_n110 ) , .A1( u0_u1_u7_n95 ) , .A2( u0_u1_u7_n96 ) );
  INV_X1 u0_u1_u7_U61 (.A( u0_u1_u7_n150 ) , .ZN( u0_u1_u7_n164 ) );
  AND2_X1 u0_u1_u7_U62 (.ZN( u0_u1_u7_n134 ) , .A1( u0_u1_u7_n93 ) , .A2( u0_u1_u7_n98 ) );
  NAND2_X1 u0_u1_u7_U63 (.A1( u0_u1_u7_n100 ) , .A2( u0_u1_u7_n102 ) , .ZN( u0_u1_u7_n129 ) );
  NAND2_X1 u0_u1_u7_U64 (.A2( u0_u1_u7_n103 ) , .ZN( u0_u1_u7_n131 ) , .A1( u0_u1_u7_n95 ) );
  NAND2_X1 u0_u1_u7_U65 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n138 ) , .A2( u0_u1_u7_n99 ) );
  NAND2_X1 u0_u1_u7_U66 (.ZN( u0_u1_u7_n132 ) , .A1( u0_u1_u7_n93 ) , .A2( u0_u1_u7_n96 ) );
  NAND2_X1 u0_u1_u7_U67 (.A1( u0_u1_u7_n100 ) , .ZN( u0_u1_u7_n148 ) , .A2( u0_u1_u7_n95 ) );
  NOR2_X1 u0_u1_u7_U68 (.A2( u0_u1_X_47 ) , .ZN( u0_u1_u7_n150 ) , .A1( u0_u1_u7_n163 ) );
  NOR2_X1 u0_u1_u7_U69 (.A2( u0_u1_X_43 ) , .A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n103 ) );
  AOI211_X1 u0_u1_u7_U7 (.ZN( u0_u1_u7_n116 ) , .A( u0_u1_u7_n155 ) , .C1( u0_u1_u7_n161 ) , .C2( u0_u1_u7_n171 ) , .B( u0_u1_u7_n94 ) );
  NOR2_X1 u0_u1_u7_U70 (.A2( u0_u1_X_48 ) , .A1( u0_u1_u7_n166 ) , .ZN( u0_u1_u7_n95 ) );
  NOR2_X1 u0_u1_u7_U71 (.A2( u0_u1_X_45 ) , .A1( u0_u1_X_48 ) , .ZN( u0_u1_u7_n99 ) );
  NOR2_X1 u0_u1_u7_U72 (.A2( u0_u1_X_44 ) , .A1( u0_u1_u7_n167 ) , .ZN( u0_u1_u7_n98 ) );
  NOR2_X1 u0_u1_u7_U73 (.A2( u0_u1_X_46 ) , .A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n152 ) );
  AND2_X1 u0_u1_u7_U74 (.A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n156 ) , .A2( u0_u1_u7_n163 ) );
  NAND2_X1 u0_u1_u7_U75 (.A2( u0_u1_X_46 ) , .A1( u0_u1_X_47 ) , .ZN( u0_u1_u7_n125 ) );
  AND2_X1 u0_u1_u7_U76 (.A2( u0_u1_X_45 ) , .A1( u0_u1_X_48 ) , .ZN( u0_u1_u7_n102 ) );
  AND2_X1 u0_u1_u7_U77 (.A2( u0_u1_X_43 ) , .A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n96 ) );
  AND2_X1 u0_u1_u7_U78 (.A1( u0_u1_X_44 ) , .ZN( u0_u1_u7_n100 ) , .A2( u0_u1_u7_n167 ) );
  AND2_X1 u0_u1_u7_U79 (.A1( u0_u1_X_48 ) , .A2( u0_u1_u7_n166 ) , .ZN( u0_u1_u7_n93 ) );
  OAI222_X1 u0_u1_u7_U8 (.C2( u0_u1_u7_n101 ) , .B2( u0_u1_u7_n111 ) , .A1( u0_u1_u7_n113 ) , .C1( u0_u1_u7_n146 ) , .A2( u0_u1_u7_n162 ) , .B1( u0_u1_u7_n164 ) , .ZN( u0_u1_u7_n94 ) );
  INV_X1 u0_u1_u7_U80 (.A( u0_u1_X_46 ) , .ZN( u0_u1_u7_n163 ) );
  INV_X1 u0_u1_u7_U81 (.A( u0_u1_X_43 ) , .ZN( u0_u1_u7_n167 ) );
  INV_X1 u0_u1_u7_U82 (.A( u0_u1_X_45 ) , .ZN( u0_u1_u7_n166 ) );
  NAND4_X1 u0_u1_u7_U83 (.ZN( u0_out1_27 ) , .A4( u0_u1_u7_n118 ) , .A3( u0_u1_u7_n119 ) , .A2( u0_u1_u7_n120 ) , .A1( u0_u1_u7_n121 ) );
  OAI21_X1 u0_u1_u7_U84 (.ZN( u0_u1_u7_n121 ) , .B2( u0_u1_u7_n145 ) , .A( u0_u1_u7_n150 ) , .B1( u0_u1_u7_n174 ) );
  OAI21_X1 u0_u1_u7_U85 (.ZN( u0_u1_u7_n120 ) , .A( u0_u1_u7_n161 ) , .B2( u0_u1_u7_n170 ) , .B1( u0_u1_u7_n179 ) );
  NAND4_X1 u0_u1_u7_U86 (.ZN( u0_out1_15 ) , .A4( u0_u1_u7_n142 ) , .A3( u0_u1_u7_n143 ) , .A2( u0_u1_u7_n144 ) , .A1( u0_u1_u7_n178 ) );
  OR2_X1 u0_u1_u7_U87 (.A2( u0_u1_u7_n125 ) , .A1( u0_u1_u7_n129 ) , .ZN( u0_u1_u7_n144 ) );
  AOI22_X1 u0_u1_u7_U88 (.A2( u0_u1_u7_n126 ) , .ZN( u0_u1_u7_n143 ) , .B2( u0_u1_u7_n165 ) , .B1( u0_u1_u7_n173 ) , .A1( u0_u1_u7_n174 ) );
  NAND4_X1 u0_u1_u7_U89 (.ZN( u0_out1_5 ) , .A4( u0_u1_u7_n108 ) , .A3( u0_u1_u7_n109 ) , .A1( u0_u1_u7_n116 ) , .A2( u0_u1_u7_n123 ) );
  OAI221_X1 u0_u1_u7_U9 (.C1( u0_u1_u7_n101 ) , .C2( u0_u1_u7_n147 ) , .ZN( u0_u1_u7_n155 ) , .B2( u0_u1_u7_n162 ) , .A( u0_u1_u7_n91 ) , .B1( u0_u1_u7_n92 ) );
  AOI22_X1 u0_u1_u7_U90 (.ZN( u0_u1_u7_n109 ) , .A2( u0_u1_u7_n126 ) , .B2( u0_u1_u7_n145 ) , .B1( u0_u1_u7_n156 ) , .A1( u0_u1_u7_n171 ) );
  NOR4_X1 u0_u1_u7_U91 (.A4( u0_u1_u7_n104 ) , .A3( u0_u1_u7_n105 ) , .A2( u0_u1_u7_n106 ) , .A1( u0_u1_u7_n107 ) , .ZN( u0_u1_u7_n108 ) );
  NAND4_X1 u0_u1_u7_U92 (.ZN( u0_out1_21 ) , .A4( u0_u1_u7_n157 ) , .A3( u0_u1_u7_n158 ) , .A2( u0_u1_u7_n159 ) , .A1( u0_u1_u7_n160 ) );
  OAI21_X1 u0_u1_u7_U93 (.B1( u0_u1_u7_n145 ) , .ZN( u0_u1_u7_n160 ) , .A( u0_u1_u7_n161 ) , .B2( u0_u1_u7_n177 ) );
  AOI22_X1 u0_u1_u7_U94 (.B2( u0_u1_u7_n149 ) , .B1( u0_u1_u7_n150 ) , .A2( u0_u1_u7_n151 ) , .A1( u0_u1_u7_n152 ) , .ZN( u0_u1_u7_n158 ) );
  NAND3_X1 u0_u1_u7_U95 (.A3( u0_u1_u7_n146 ) , .A2( u0_u1_u7_n147 ) , .A1( u0_u1_u7_n148 ) , .ZN( u0_u1_u7_n151 ) );
  NAND3_X1 u0_u1_u7_U96 (.A3( u0_u1_u7_n131 ) , .A2( u0_u1_u7_n132 ) , .A1( u0_u1_u7_n133 ) , .ZN( u0_u1_u7_n135 ) );
  XOR2_X1 u0_u5_U13 (.B( u0_K6_42 ) , .A( u0_R4_29 ) , .Z( u0_u5_X_42 ) );
  XOR2_X1 u0_u5_U14 (.B( u0_K6_41 ) , .A( u0_R4_28 ) , .Z( u0_u5_X_41 ) );
  XOR2_X1 u0_u5_U15 (.B( u0_K6_40 ) , .A( u0_R4_27 ) , .Z( u0_u5_X_40 ) );
  XOR2_X1 u0_u5_U17 (.B( u0_K6_39 ) , .A( u0_R4_26 ) , .Z( u0_u5_X_39 ) );
  XOR2_X1 u0_u5_U18 (.B( u0_K6_38 ) , .A( u0_R4_25 ) , .Z( u0_u5_X_38 ) );
  XOR2_X1 u0_u5_U19 (.B( u0_K6_37 ) , .A( u0_R4_24 ) , .Z( u0_u5_X_37 ) );
  XOR2_X1 u0_u5_U26 (.B( u0_K6_30 ) , .A( u0_R4_21 ) , .Z( u0_u5_X_30 ) );
  XOR2_X1 u0_u5_U28 (.B( u0_K6_29 ) , .A( u0_R4_20 ) , .Z( u0_u5_X_29 ) );
  XOR2_X1 u0_u5_U29 (.B( u0_K6_28 ) , .A( u0_R4_19 ) , .Z( u0_u5_X_28 ) );
  XOR2_X1 u0_u5_U30 (.B( u0_K6_27 ) , .A( u0_R4_18 ) , .Z( u0_u5_X_27 ) );
  XOR2_X1 u0_u5_U31 (.B( u0_K6_26 ) , .A( u0_R4_17 ) , .Z( u0_u5_X_26 ) );
  XOR2_X1 u0_u5_U32 (.B( u0_K6_25 ) , .A( u0_R4_16 ) , .Z( u0_u5_X_25 ) );
  OAI22_X1 u0_u5_u4_U10 (.B2( u0_u5_u4_n135 ) , .ZN( u0_u5_u4_n137 ) , .B1( u0_u5_u4_n153 ) , .A1( u0_u5_u4_n155 ) , .A2( u0_u5_u4_n171 ) );
  AND3_X1 u0_u5_u4_U11 (.A2( u0_u5_u4_n134 ) , .ZN( u0_u5_u4_n135 ) , .A3( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n157 ) );
  NAND2_X1 u0_u5_u4_U12 (.ZN( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n173 ) );
  AOI21_X1 u0_u5_u4_U13 (.B2( u0_u5_u4_n160 ) , .B1( u0_u5_u4_n161 ) , .ZN( u0_u5_u4_n162 ) , .A( u0_u5_u4_n170 ) );
  AOI21_X1 u0_u5_u4_U14 (.ZN( u0_u5_u4_n107 ) , .B2( u0_u5_u4_n143 ) , .A( u0_u5_u4_n174 ) , .B1( u0_u5_u4_n184 ) );
  AOI21_X1 u0_u5_u4_U15 (.B2( u0_u5_u4_n158 ) , .B1( u0_u5_u4_n159 ) , .ZN( u0_u5_u4_n163 ) , .A( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U16 (.A( u0_u5_u4_n153 ) , .B2( u0_u5_u4_n154 ) , .B1( u0_u5_u4_n155 ) , .ZN( u0_u5_u4_n165 ) );
  AOI21_X1 u0_u5_u4_U17 (.A( u0_u5_u4_n156 ) , .B2( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n164 ) , .B1( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U18 (.A( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n170 ) );
  AND2_X1 u0_u5_u4_U19 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n155 ) , .A1( u0_u5_u4_n160 ) );
  INV_X1 u0_u5_u4_U20 (.A( u0_u5_u4_n156 ) , .ZN( u0_u5_u4_n175 ) );
  NAND2_X1 u0_u5_u4_U21 (.A2( u0_u5_u4_n118 ) , .ZN( u0_u5_u4_n131 ) , .A1( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U22 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n130 ) );
  NAND2_X1 u0_u5_u4_U23 (.ZN( u0_u5_u4_n117 ) , .A2( u0_u5_u4_n118 ) , .A1( u0_u5_u4_n148 ) );
  NAND2_X1 u0_u5_u4_U24 (.ZN( u0_u5_u4_n129 ) , .A1( u0_u5_u4_n134 ) , .A2( u0_u5_u4_n148 ) );
  AND3_X1 u0_u5_u4_U25 (.A1( u0_u5_u4_n119 ) , .A2( u0_u5_u4_n143 ) , .A3( u0_u5_u4_n154 ) , .ZN( u0_u5_u4_n161 ) );
  AND2_X1 u0_u5_u4_U26 (.A1( u0_u5_u4_n145 ) , .A2( u0_u5_u4_n147 ) , .ZN( u0_u5_u4_n159 ) );
  OR3_X1 u0_u5_u4_U27 (.A3( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n115 ) , .A1( u0_u5_u4_n116 ) , .ZN( u0_u5_u4_n136 ) );
  AOI21_X1 u0_u5_u4_U28 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n116 ) , .B2( u0_u5_u4_n173 ) , .B1( u0_u5_u4_n174 ) );
  AOI21_X1 u0_u5_u4_U29 (.ZN( u0_u5_u4_n115 ) , .B2( u0_u5_u4_n145 ) , .B1( u0_u5_u4_n146 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U3 (.ZN( u0_u5_u4_n121 ) , .A1( u0_u5_u4_n181 ) , .A2( u0_u5_u4_n182 ) );
  OAI22_X1 u0_u5_u4_U30 (.ZN( u0_u5_u4_n114 ) , .A2( u0_u5_u4_n121 ) , .B1( u0_u5_u4_n160 ) , .B2( u0_u5_u4_n170 ) , .A1( u0_u5_u4_n171 ) );
  INV_X1 u0_u5_u4_U31 (.A( u0_u5_u4_n158 ) , .ZN( u0_u5_u4_n182 ) );
  INV_X1 u0_u5_u4_U32 (.ZN( u0_u5_u4_n181 ) , .A( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U33 (.A( u0_u5_u4_n144 ) , .ZN( u0_u5_u4_n179 ) );
  INV_X1 u0_u5_u4_U34 (.A( u0_u5_u4_n157 ) , .ZN( u0_u5_u4_n178 ) );
  NAND2_X1 u0_u5_u4_U35 (.A2( u0_u5_u4_n154 ) , .A1( u0_u5_u4_n96 ) , .ZN( u0_u5_u4_n97 ) );
  INV_X1 u0_u5_u4_U36 (.ZN( u0_u5_u4_n186 ) , .A( u0_u5_u4_n95 ) );
  OAI221_X1 u0_u5_u4_U37 (.C1( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n158 ) , .B2( u0_u5_u4_n171 ) , .C2( u0_u5_u4_n173 ) , .A( u0_u5_u4_n94 ) , .ZN( u0_u5_u4_n95 ) );
  AOI222_X1 u0_u5_u4_U38 (.B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n138 ) , .C2( u0_u5_u4_n175 ) , .A2( u0_u5_u4_n179 ) , .C1( u0_u5_u4_n181 ) , .B1( u0_u5_u4_n185 ) , .ZN( u0_u5_u4_n94 ) );
  INV_X1 u0_u5_u4_U39 (.A( u0_u5_u4_n113 ) , .ZN( u0_u5_u4_n185 ) );
  INV_X1 u0_u5_u4_U4 (.A( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n184 ) );
  INV_X1 u0_u5_u4_U40 (.A( u0_u5_u4_n143 ) , .ZN( u0_u5_u4_n183 ) );
  NOR2_X1 u0_u5_u4_U41 (.ZN( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n168 ) , .A2( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U42 (.A1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n153 ) );
  NOR2_X1 u0_u5_u4_U43 (.A2( u0_u5_u4_n128 ) , .A1( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n156 ) );
  AOI22_X1 u0_u5_u4_U44 (.B2( u0_u5_u4_n122 ) , .A1( u0_u5_u4_n123 ) , .ZN( u0_u5_u4_n124 ) , .B1( u0_u5_u4_n128 ) , .A2( u0_u5_u4_n172 ) );
  INV_X1 u0_u5_u4_U45 (.A( u0_u5_u4_n153 ) , .ZN( u0_u5_u4_n172 ) );
  NAND2_X1 u0_u5_u4_U46 (.A2( u0_u5_u4_n120 ) , .ZN( u0_u5_u4_n123 ) , .A1( u0_u5_u4_n161 ) );
  AOI22_X1 u0_u5_u4_U47 (.B2( u0_u5_u4_n132 ) , .A2( u0_u5_u4_n133 ) , .ZN( u0_u5_u4_n140 ) , .A1( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n179 ) );
  NAND2_X1 u0_u5_u4_U48 (.ZN( u0_u5_u4_n133 ) , .A2( u0_u5_u4_n146 ) , .A1( u0_u5_u4_n154 ) );
  NAND2_X1 u0_u5_u4_U49 (.A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n154 ) , .A2( u0_u5_u4_n98 ) );
  NOR4_X1 u0_u5_u4_U5 (.A4( u0_u5_u4_n106 ) , .A3( u0_u5_u4_n107 ) , .A2( u0_u5_u4_n108 ) , .A1( u0_u5_u4_n109 ) , .ZN( u0_u5_u4_n110 ) );
  NAND2_X1 u0_u5_u4_U50 (.A1( u0_u5_u4_n101 ) , .ZN( u0_u5_u4_n158 ) , .A2( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U51 (.ZN( u0_u5_u4_n127 ) , .A( u0_u5_u4_n136 ) , .B2( u0_u5_u4_n150 ) , .B1( u0_u5_u4_n180 ) );
  INV_X1 u0_u5_u4_U52 (.A( u0_u5_u4_n160 ) , .ZN( u0_u5_u4_n180 ) );
  NAND2_X1 u0_u5_u4_U53 (.A2( u0_u5_u4_n104 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n146 ) );
  NAND2_X1 u0_u5_u4_U54 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n160 ) );
  NAND2_X1 u0_u5_u4_U55 (.ZN( u0_u5_u4_n134 ) , .A1( u0_u5_u4_n98 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U56 (.A1( u0_u5_u4_n103 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n143 ) );
  NAND2_X1 u0_u5_u4_U57 (.A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n145 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U58 (.A1( u0_u5_u4_n100 ) , .A2( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n120 ) );
  NAND2_X1 u0_u5_u4_U59 (.A1( u0_u5_u4_n102 ) , .A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n148 ) );
  AOI21_X1 u0_u5_u4_U6 (.ZN( u0_u5_u4_n106 ) , .B2( u0_u5_u4_n146 ) , .B1( u0_u5_u4_n158 ) , .A( u0_u5_u4_n170 ) );
  NAND2_X1 u0_u5_u4_U60 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n157 ) );
  INV_X1 u0_u5_u4_U61 (.A( u0_u5_u4_n150 ) , .ZN( u0_u5_u4_n173 ) );
  INV_X1 u0_u5_u4_U62 (.A( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n171 ) );
  NAND2_X1 u0_u5_u4_U63 (.A1( u0_u5_u4_n100 ) , .ZN( u0_u5_u4_n118 ) , .A2( u0_u5_u4_n99 ) );
  NAND2_X1 u0_u5_u4_U64 (.A2( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n144 ) );
  NAND2_X1 u0_u5_u4_U65 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n105 ) , .ZN( u0_u5_u4_n96 ) );
  INV_X1 u0_u5_u4_U66 (.A( u0_u5_u4_n128 ) , .ZN( u0_u5_u4_n174 ) );
  NAND2_X1 u0_u5_u4_U67 (.A2( u0_u5_u4_n102 ) , .ZN( u0_u5_u4_n119 ) , .A1( u0_u5_u4_n98 ) );
  NAND2_X1 u0_u5_u4_U68 (.A2( u0_u5_u4_n101 ) , .A1( u0_u5_u4_n103 ) , .ZN( u0_u5_u4_n147 ) );
  NAND2_X1 u0_u5_u4_U69 (.A2( u0_u5_u4_n104 ) , .ZN( u0_u5_u4_n113 ) , .A1( u0_u5_u4_n99 ) );
  AOI21_X1 u0_u5_u4_U7 (.ZN( u0_u5_u4_n108 ) , .B2( u0_u5_u4_n134 ) , .B1( u0_u5_u4_n155 ) , .A( u0_u5_u4_n156 ) );
  NOR2_X1 u0_u5_u4_U70 (.A2( u0_u5_X_28 ) , .ZN( u0_u5_u4_n150 ) , .A1( u0_u5_u4_n168 ) );
  NOR2_X1 u0_u5_u4_U71 (.A2( u0_u5_X_29 ) , .ZN( u0_u5_u4_n152 ) , .A1( u0_u5_u4_n169 ) );
  NOR2_X1 u0_u5_u4_U72 (.A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n105 ) , .A1( u0_u5_u4_n176 ) );
  NOR2_X1 u0_u5_u4_U73 (.A2( u0_u5_X_26 ) , .ZN( u0_u5_u4_n100 ) , .A1( u0_u5_u4_n177 ) );
  NOR2_X1 u0_u5_u4_U74 (.A2( u0_u5_X_28 ) , .A1( u0_u5_X_29 ) , .ZN( u0_u5_u4_n128 ) );
  NOR2_X1 u0_u5_u4_U75 (.A2( u0_u5_X_27 ) , .A1( u0_u5_X_30 ) , .ZN( u0_u5_u4_n102 ) );
  NOR2_X1 u0_u5_u4_U76 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n98 ) );
  AND2_X1 u0_u5_u4_U77 (.A2( u0_u5_X_25 ) , .A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n104 ) );
  AND2_X1 u0_u5_u4_U78 (.A1( u0_u5_X_30 ) , .A2( u0_u5_u4_n176 ) , .ZN( u0_u5_u4_n99 ) );
  AND2_X1 u0_u5_u4_U79 (.A1( u0_u5_X_26 ) , .ZN( u0_u5_u4_n101 ) , .A2( u0_u5_u4_n177 ) );
  AOI21_X1 u0_u5_u4_U8 (.ZN( u0_u5_u4_n109 ) , .A( u0_u5_u4_n153 ) , .B1( u0_u5_u4_n159 ) , .B2( u0_u5_u4_n184 ) );
  AND2_X1 u0_u5_u4_U80 (.A1( u0_u5_X_27 ) , .A2( u0_u5_X_30 ) , .ZN( u0_u5_u4_n103 ) );
  INV_X1 u0_u5_u4_U81 (.A( u0_u5_X_28 ) , .ZN( u0_u5_u4_n169 ) );
  INV_X1 u0_u5_u4_U82 (.A( u0_u5_X_29 ) , .ZN( u0_u5_u4_n168 ) );
  INV_X1 u0_u5_u4_U83 (.A( u0_u5_X_25 ) , .ZN( u0_u5_u4_n177 ) );
  INV_X1 u0_u5_u4_U84 (.A( u0_u5_X_27 ) , .ZN( u0_u5_u4_n176 ) );
  NAND4_X1 u0_u5_u4_U85 (.ZN( u0_out5_25 ) , .A4( u0_u5_u4_n139 ) , .A3( u0_u5_u4_n140 ) , .A2( u0_u5_u4_n141 ) , .A1( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U86 (.A( u0_u5_u4_n128 ) , .B2( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n130 ) , .ZN( u0_u5_u4_n142 ) );
  OAI21_X1 u0_u5_u4_U87 (.B2( u0_u5_u4_n131 ) , .ZN( u0_u5_u4_n141 ) , .A( u0_u5_u4_n175 ) , .B1( u0_u5_u4_n183 ) );
  NAND4_X1 u0_u5_u4_U88 (.ZN( u0_out5_14 ) , .A4( u0_u5_u4_n124 ) , .A3( u0_u5_u4_n125 ) , .A2( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n127 ) );
  AOI22_X1 u0_u5_u4_U89 (.B2( u0_u5_u4_n117 ) , .ZN( u0_u5_u4_n126 ) , .A1( u0_u5_u4_n129 ) , .B1( u0_u5_u4_n152 ) , .A2( u0_u5_u4_n175 ) );
  AOI211_X1 u0_u5_u4_U9 (.B( u0_u5_u4_n136 ) , .A( u0_u5_u4_n137 ) , .C2( u0_u5_u4_n138 ) , .ZN( u0_u5_u4_n139 ) , .C1( u0_u5_u4_n182 ) );
  AOI22_X1 u0_u5_u4_U90 (.ZN( u0_u5_u4_n125 ) , .B2( u0_u5_u4_n131 ) , .A2( u0_u5_u4_n132 ) , .B1( u0_u5_u4_n138 ) , .A1( u0_u5_u4_n178 ) );
  NAND4_X1 u0_u5_u4_U91 (.ZN( u0_out5_8 ) , .A4( u0_u5_u4_n110 ) , .A3( u0_u5_u4_n111 ) , .A2( u0_u5_u4_n112 ) , .A1( u0_u5_u4_n186 ) );
  NAND2_X1 u0_u5_u4_U92 (.ZN( u0_u5_u4_n112 ) , .A2( u0_u5_u4_n130 ) , .A1( u0_u5_u4_n150 ) );
  AOI22_X1 u0_u5_u4_U93 (.ZN( u0_u5_u4_n111 ) , .B2( u0_u5_u4_n132 ) , .A1( u0_u5_u4_n152 ) , .B1( u0_u5_u4_n178 ) , .A2( u0_u5_u4_n97 ) );
  AOI22_X1 u0_u5_u4_U94 (.B2( u0_u5_u4_n149 ) , .B1( u0_u5_u4_n150 ) , .A2( u0_u5_u4_n151 ) , .A1( u0_u5_u4_n152 ) , .ZN( u0_u5_u4_n167 ) );
  NOR4_X1 u0_u5_u4_U95 (.A4( u0_u5_u4_n162 ) , .A3( u0_u5_u4_n163 ) , .A2( u0_u5_u4_n164 ) , .A1( u0_u5_u4_n165 ) , .ZN( u0_u5_u4_n166 ) );
  NAND3_X1 u0_u5_u4_U96 (.ZN( u0_out5_3 ) , .A3( u0_u5_u4_n166 ) , .A1( u0_u5_u4_n167 ) , .A2( u0_u5_u4_n186 ) );
  NAND3_X1 u0_u5_u4_U97 (.A3( u0_u5_u4_n146 ) , .A2( u0_u5_u4_n147 ) , .A1( u0_u5_u4_n148 ) , .ZN( u0_u5_u4_n149 ) );
  NAND3_X1 u0_u5_u4_U98 (.A3( u0_u5_u4_n143 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n145 ) , .ZN( u0_u5_u4_n151 ) );
  NAND3_X1 u0_u5_u4_U99 (.A3( u0_u5_u4_n121 ) , .ZN( u0_u5_u4_n122 ) , .A2( u0_u5_u4_n144 ) , .A1( u0_u5_u4_n154 ) );
  OAI21_X1 u0_u5_u6_U10 (.A( u0_u5_u6_n159 ) , .B1( u0_u5_u6_n169 ) , .B2( u0_u5_u6_n173 ) , .ZN( u0_u5_u6_n90 ) );
  INV_X1 u0_u5_u6_U11 (.ZN( u0_u5_u6_n172 ) , .A( u0_u5_u6_n88 ) );
  AOI22_X1 u0_u5_u6_U12 (.A2( u0_u5_u6_n151 ) , .B2( u0_u5_u6_n161 ) , .A1( u0_u5_u6_n167 ) , .B1( u0_u5_u6_n170 ) , .ZN( u0_u5_u6_n89 ) );
  AOI21_X1 u0_u5_u6_U13 (.ZN( u0_u5_u6_n106 ) , .A( u0_u5_u6_n142 ) , .B2( u0_u5_u6_n159 ) , .B1( u0_u5_u6_n164 ) );
  INV_X1 u0_u5_u6_U14 (.A( u0_u5_u6_n155 ) , .ZN( u0_u5_u6_n161 ) );
  INV_X1 u0_u5_u6_U15 (.A( u0_u5_u6_n128 ) , .ZN( u0_u5_u6_n164 ) );
  NAND2_X1 u0_u5_u6_U16 (.ZN( u0_u5_u6_n110 ) , .A1( u0_u5_u6_n122 ) , .A2( u0_u5_u6_n129 ) );
  NAND2_X1 u0_u5_u6_U17 (.ZN( u0_u5_u6_n124 ) , .A2( u0_u5_u6_n146 ) , .A1( u0_u5_u6_n148 ) );
  INV_X1 u0_u5_u6_U18 (.A( u0_u5_u6_n132 ) , .ZN( u0_u5_u6_n171 ) );
  AND2_X1 u0_u5_u6_U19 (.A1( u0_u5_u6_n100 ) , .ZN( u0_u5_u6_n130 ) , .A2( u0_u5_u6_n147 ) );
  INV_X1 u0_u5_u6_U20 (.A( u0_u5_u6_n127 ) , .ZN( u0_u5_u6_n173 ) );
  INV_X1 u0_u5_u6_U21 (.A( u0_u5_u6_n121 ) , .ZN( u0_u5_u6_n167 ) );
  INV_X1 u0_u5_u6_U22 (.A( u0_u5_u6_n100 ) , .ZN( u0_u5_u6_n169 ) );
  INV_X1 u0_u5_u6_U23 (.A( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n170 ) );
  INV_X1 u0_u5_u6_U24 (.A( u0_u5_u6_n113 ) , .ZN( u0_u5_u6_n168 ) );
  AND2_X1 u0_u5_u6_U25 (.A1( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n119 ) , .ZN( u0_u5_u6_n133 ) );
  AND2_X1 u0_u5_u6_U26 (.A2( u0_u5_u6_n121 ) , .A1( u0_u5_u6_n122 ) , .ZN( u0_u5_u6_n131 ) );
  AND3_X1 u0_u5_u6_U27 (.ZN( u0_u5_u6_n120 ) , .A2( u0_u5_u6_n127 ) , .A1( u0_u5_u6_n132 ) , .A3( u0_u5_u6_n145 ) );
  INV_X1 u0_u5_u6_U28 (.A( u0_u5_u6_n146 ) , .ZN( u0_u5_u6_n163 ) );
  AOI222_X1 u0_u5_u6_U29 (.ZN( u0_u5_u6_n114 ) , .A1( u0_u5_u6_n118 ) , .A2( u0_u5_u6_n126 ) , .B2( u0_u5_u6_n151 ) , .C2( u0_u5_u6_n159 ) , .C1( u0_u5_u6_n168 ) , .B1( u0_u5_u6_n169 ) );
  INV_X1 u0_u5_u6_U3 (.A( u0_u5_u6_n110 ) , .ZN( u0_u5_u6_n166 ) );
  NOR2_X1 u0_u5_u6_U30 (.A1( u0_u5_u6_n162 ) , .A2( u0_u5_u6_n165 ) , .ZN( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U31 (.A1( u0_u5_u6_n144 ) , .ZN( u0_u5_u6_n151 ) , .A2( u0_u5_u6_n158 ) );
  NAND2_X1 u0_u5_u6_U32 (.ZN( u0_u5_u6_n132 ) , .A1( u0_u5_u6_n91 ) , .A2( u0_u5_u6_n97 ) );
  NOR2_X1 u0_u5_u6_U33 (.A2( u0_u5_u6_n126 ) , .ZN( u0_u5_u6_n155 ) , .A1( u0_u5_u6_n160 ) );
  NAND2_X1 u0_u5_u6_U34 (.ZN( u0_u5_u6_n146 ) , .A2( u0_u5_u6_n94 ) , .A1( u0_u5_u6_n99 ) );
  AOI21_X1 u0_u5_u6_U35 (.A( u0_u5_u6_n144 ) , .B2( u0_u5_u6_n145 ) , .B1( u0_u5_u6_n146 ) , .ZN( u0_u5_u6_n150 ) );
  INV_X1 u0_u5_u6_U36 (.A( u0_u5_u6_n111 ) , .ZN( u0_u5_u6_n158 ) );
  NAND2_X1 u0_u5_u6_U37 (.ZN( u0_u5_u6_n127 ) , .A1( u0_u5_u6_n91 ) , .A2( u0_u5_u6_n92 ) );
  NAND2_X1 u0_u5_u6_U38 (.ZN( u0_u5_u6_n129 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n96 ) );
  INV_X1 u0_u5_u6_U39 (.A( u0_u5_u6_n144 ) , .ZN( u0_u5_u6_n159 ) );
  INV_X1 u0_u5_u6_U4 (.A( u0_u5_u6_n142 ) , .ZN( u0_u5_u6_n174 ) );
  NAND2_X1 u0_u5_u6_U40 (.ZN( u0_u5_u6_n145 ) , .A2( u0_u5_u6_n97 ) , .A1( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U41 (.ZN( u0_u5_u6_n148 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n94 ) );
  NAND2_X1 u0_u5_u6_U42 (.ZN( u0_u5_u6_n108 ) , .A2( u0_u5_u6_n139 ) , .A1( u0_u5_u6_n144 ) );
  NAND2_X1 u0_u5_u6_U43 (.ZN( u0_u5_u6_n121 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n97 ) );
  NAND2_X1 u0_u5_u6_U44 (.ZN( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n95 ) );
  AND2_X1 u0_u5_u6_U45 (.ZN( u0_u5_u6_n118 ) , .A2( u0_u5_u6_n91 ) , .A1( u0_u5_u6_n99 ) );
  AOI22_X1 u0_u5_u6_U46 (.B2( u0_u5_u6_n110 ) , .B1( u0_u5_u6_n111 ) , .A1( u0_u5_u6_n112 ) , .ZN( u0_u5_u6_n115 ) , .A2( u0_u5_u6_n161 ) );
  NAND4_X1 u0_u5_u6_U47 (.A3( u0_u5_u6_n109 ) , .ZN( u0_u5_u6_n112 ) , .A4( u0_u5_u6_n132 ) , .A2( u0_u5_u6_n147 ) , .A1( u0_u5_u6_n166 ) );
  NOR2_X1 u0_u5_u6_U48 (.ZN( u0_u5_u6_n109 ) , .A1( u0_u5_u6_n170 ) , .A2( u0_u5_u6_n173 ) );
  NAND2_X1 u0_u5_u6_U49 (.ZN( u0_u5_u6_n147 ) , .A2( u0_u5_u6_n98 ) , .A1( u0_u5_u6_n99 ) );
  NAND2_X1 u0_u5_u6_U5 (.A2( u0_u5_u6_n143 ) , .ZN( u0_u5_u6_n152 ) , .A1( u0_u5_u6_n166 ) );
  NAND2_X1 u0_u5_u6_U50 (.ZN( u0_u5_u6_n128 ) , .A1( u0_u5_u6_n94 ) , .A2( u0_u5_u6_n96 ) );
  AOI211_X1 u0_u5_u6_U51 (.B( u0_u5_u6_n134 ) , .A( u0_u5_u6_n135 ) , .C1( u0_u5_u6_n136 ) , .ZN( u0_u5_u6_n137 ) , .C2( u0_u5_u6_n151 ) );
  AOI21_X1 u0_u5_u6_U52 (.B2( u0_u5_u6_n132 ) , .B1( u0_u5_u6_n133 ) , .ZN( u0_u5_u6_n134 ) , .A( u0_u5_u6_n158 ) );
  AOI21_X1 u0_u5_u6_U53 (.B1( u0_u5_u6_n131 ) , .ZN( u0_u5_u6_n135 ) , .A( u0_u5_u6_n144 ) , .B2( u0_u5_u6_n146 ) );
  NAND4_X1 u0_u5_u6_U54 (.A4( u0_u5_u6_n127 ) , .A3( u0_u5_u6_n128 ) , .A2( u0_u5_u6_n129 ) , .A1( u0_u5_u6_n130 ) , .ZN( u0_u5_u6_n136 ) );
  NAND2_X1 u0_u5_u6_U55 (.ZN( u0_u5_u6_n119 ) , .A2( u0_u5_u6_n95 ) , .A1( u0_u5_u6_n99 ) );
  NAND2_X1 u0_u5_u6_U56 (.ZN( u0_u5_u6_n123 ) , .A2( u0_u5_u6_n91 ) , .A1( u0_u5_u6_n96 ) );
  NAND2_X1 u0_u5_u6_U57 (.ZN( u0_u5_u6_n100 ) , .A2( u0_u5_u6_n92 ) , .A1( u0_u5_u6_n98 ) );
  NAND2_X1 u0_u5_u6_U58 (.ZN( u0_u5_u6_n122 ) , .A1( u0_u5_u6_n94 ) , .A2( u0_u5_u6_n97 ) );
  INV_X1 u0_u5_u6_U59 (.A( u0_u5_u6_n139 ) , .ZN( u0_u5_u6_n160 ) );
  AOI22_X1 u0_u5_u6_U6 (.B2( u0_u5_u6_n101 ) , .A1( u0_u5_u6_n102 ) , .ZN( u0_u5_u6_n103 ) , .B1( u0_u5_u6_n160 ) , .A2( u0_u5_u6_n161 ) );
  NAND2_X1 u0_u5_u6_U60 (.ZN( u0_u5_u6_n113 ) , .A1( u0_u5_u6_n96 ) , .A2( u0_u5_u6_n98 ) );
  NOR2_X1 u0_u5_u6_U61 (.A2( u0_u5_X_40 ) , .A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n126 ) );
  NOR2_X1 u0_u5_u6_U62 (.A2( u0_u5_X_39 ) , .A1( u0_u5_X_42 ) , .ZN( u0_u5_u6_n92 ) );
  NOR2_X1 u0_u5_u6_U63 (.A2( u0_u5_X_39 ) , .A1( u0_u5_u6_n156 ) , .ZN( u0_u5_u6_n97 ) );
  NOR2_X1 u0_u5_u6_U64 (.A2( u0_u5_X_38 ) , .A1( u0_u5_u6_n165 ) , .ZN( u0_u5_u6_n95 ) );
  NOR2_X1 u0_u5_u6_U65 (.A2( u0_u5_X_41 ) , .ZN( u0_u5_u6_n111 ) , .A1( u0_u5_u6_n157 ) );
  NOR2_X1 u0_u5_u6_U66 (.A2( u0_u5_X_37 ) , .A1( u0_u5_u6_n162 ) , .ZN( u0_u5_u6_n94 ) );
  NOR2_X1 u0_u5_u6_U67 (.A2( u0_u5_X_37 ) , .A1( u0_u5_X_38 ) , .ZN( u0_u5_u6_n91 ) );
  NAND2_X1 u0_u5_u6_U68 (.A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n144 ) , .A2( u0_u5_u6_n157 ) );
  NAND2_X1 u0_u5_u6_U69 (.A2( u0_u5_X_40 ) , .A1( u0_u5_X_41 ) , .ZN( u0_u5_u6_n139 ) );
  NOR2_X1 u0_u5_u6_U7 (.A1( u0_u5_u6_n118 ) , .ZN( u0_u5_u6_n143 ) , .A2( u0_u5_u6_n168 ) );
  AND2_X1 u0_u5_u6_U70 (.A1( u0_u5_X_39 ) , .A2( u0_u5_u6_n156 ) , .ZN( u0_u5_u6_n96 ) );
  AND2_X1 u0_u5_u6_U71 (.A1( u0_u5_X_39 ) , .A2( u0_u5_X_42 ) , .ZN( u0_u5_u6_n99 ) );
  INV_X1 u0_u5_u6_U72 (.A( u0_u5_X_40 ) , .ZN( u0_u5_u6_n157 ) );
  INV_X1 u0_u5_u6_U73 (.A( u0_u5_X_37 ) , .ZN( u0_u5_u6_n165 ) );
  INV_X1 u0_u5_u6_U74 (.A( u0_u5_X_38 ) , .ZN( u0_u5_u6_n162 ) );
  INV_X1 u0_u5_u6_U75 (.A( u0_u5_X_42 ) , .ZN( u0_u5_u6_n156 ) );
  NAND4_X1 u0_u5_u6_U76 (.ZN( u0_out5_32 ) , .A4( u0_u5_u6_n103 ) , .A3( u0_u5_u6_n104 ) , .A2( u0_u5_u6_n105 ) , .A1( u0_u5_u6_n106 ) );
  AOI22_X1 u0_u5_u6_U77 (.ZN( u0_u5_u6_n105 ) , .A2( u0_u5_u6_n108 ) , .A1( u0_u5_u6_n118 ) , .B2( u0_u5_u6_n126 ) , .B1( u0_u5_u6_n171 ) );
  AOI22_X1 u0_u5_u6_U78 (.ZN( u0_u5_u6_n104 ) , .A1( u0_u5_u6_n111 ) , .B1( u0_u5_u6_n124 ) , .B2( u0_u5_u6_n151 ) , .A2( u0_u5_u6_n93 ) );
  NAND4_X1 u0_u5_u6_U79 (.ZN( u0_out5_12 ) , .A4( u0_u5_u6_n114 ) , .A3( u0_u5_u6_n115 ) , .A2( u0_u5_u6_n116 ) , .A1( u0_u5_u6_n117 ) );
  AOI21_X1 u0_u5_u6_U8 (.B1( u0_u5_u6_n107 ) , .B2( u0_u5_u6_n132 ) , .A( u0_u5_u6_n158 ) , .ZN( u0_u5_u6_n88 ) );
  OAI22_X1 u0_u5_u6_U80 (.B2( u0_u5_u6_n111 ) , .ZN( u0_u5_u6_n116 ) , .B1( u0_u5_u6_n126 ) , .A2( u0_u5_u6_n164 ) , .A1( u0_u5_u6_n167 ) );
  OAI21_X1 u0_u5_u6_U81 (.A( u0_u5_u6_n108 ) , .ZN( u0_u5_u6_n117 ) , .B2( u0_u5_u6_n141 ) , .B1( u0_u5_u6_n163 ) );
  OAI211_X1 u0_u5_u6_U82 (.ZN( u0_out5_22 ) , .B( u0_u5_u6_n137 ) , .A( u0_u5_u6_n138 ) , .C2( u0_u5_u6_n139 ) , .C1( u0_u5_u6_n140 ) );
  AOI22_X1 u0_u5_u6_U83 (.B1( u0_u5_u6_n124 ) , .A2( u0_u5_u6_n125 ) , .A1( u0_u5_u6_n126 ) , .ZN( u0_u5_u6_n138 ) , .B2( u0_u5_u6_n161 ) );
  AND4_X1 u0_u5_u6_U84 (.A3( u0_u5_u6_n119 ) , .A1( u0_u5_u6_n120 ) , .A4( u0_u5_u6_n129 ) , .ZN( u0_u5_u6_n140 ) , .A2( u0_u5_u6_n143 ) );
  OAI211_X1 u0_u5_u6_U85 (.ZN( u0_out5_7 ) , .B( u0_u5_u6_n153 ) , .C2( u0_u5_u6_n154 ) , .C1( u0_u5_u6_n155 ) , .A( u0_u5_u6_n174 ) );
  NOR3_X1 u0_u5_u6_U86 (.A1( u0_u5_u6_n141 ) , .ZN( u0_u5_u6_n154 ) , .A3( u0_u5_u6_n164 ) , .A2( u0_u5_u6_n171 ) );
  AOI211_X1 u0_u5_u6_U87 (.B( u0_u5_u6_n149 ) , .A( u0_u5_u6_n150 ) , .C2( u0_u5_u6_n151 ) , .C1( u0_u5_u6_n152 ) , .ZN( u0_u5_u6_n153 ) );
  NAND3_X1 u0_u5_u6_U88 (.A2( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n125 ) , .A1( u0_u5_u6_n130 ) , .A3( u0_u5_u6_n131 ) );
  NAND3_X1 u0_u5_u6_U89 (.A3( u0_u5_u6_n133 ) , .ZN( u0_u5_u6_n141 ) , .A1( u0_u5_u6_n145 ) , .A2( u0_u5_u6_n148 ) );
  AOI21_X1 u0_u5_u6_U9 (.B2( u0_u5_u6_n147 ) , .B1( u0_u5_u6_n148 ) , .ZN( u0_u5_u6_n149 ) , .A( u0_u5_u6_n158 ) );
  NAND3_X1 u0_u5_u6_U90 (.ZN( u0_u5_u6_n101 ) , .A3( u0_u5_u6_n107 ) , .A2( u0_u5_u6_n121 ) , .A1( u0_u5_u6_n127 ) );
  NAND3_X1 u0_u5_u6_U91 (.ZN( u0_u5_u6_n102 ) , .A3( u0_u5_u6_n130 ) , .A2( u0_u5_u6_n145 ) , .A1( u0_u5_u6_n166 ) );
  NAND3_X1 u0_u5_u6_U92 (.A3( u0_u5_u6_n113 ) , .A1( u0_u5_u6_n119 ) , .A2( u0_u5_u6_n123 ) , .ZN( u0_u5_u6_n93 ) );
  NAND3_X1 u0_u5_u6_U93 (.ZN( u0_u5_u6_n142 ) , .A2( u0_u5_u6_n172 ) , .A3( u0_u5_u6_n89 ) , .A1( u0_u5_u6_n90 ) );
  XOR2_X1 u0_u6_U26 (.B( u0_K7_30 ) , .A( u0_R5_21 ) , .Z( u0_u6_X_30 ) );
  XOR2_X1 u0_u6_U28 (.B( u0_K7_29 ) , .A( u0_R5_20 ) , .Z( u0_u6_X_29 ) );
  XOR2_X1 u0_u6_U29 (.B( u0_K7_28 ) , .A( u0_R5_19 ) , .Z( u0_u6_X_28 ) );
  XOR2_X1 u0_u6_U30 (.B( u0_K7_27 ) , .A( u0_R5_18 ) , .Z( u0_u6_X_27 ) );
  XOR2_X1 u0_u6_U31 (.B( u0_K7_26 ) , .A( u0_R5_17 ) , .Z( u0_u6_X_26 ) );
  XOR2_X1 u0_u6_U32 (.B( u0_K7_25 ) , .A( u0_R5_16 ) , .Z( u0_u6_X_25 ) );
  XOR2_X1 u0_u6_U33 (.B( u0_K7_24 ) , .A( u0_R5_17 ) , .Z( u0_u6_X_24 ) );
  XOR2_X1 u0_u6_U34 (.B( u0_K7_23 ) , .A( u0_R5_16 ) , .Z( u0_u6_X_23 ) );
  XOR2_X1 u0_u6_U35 (.B( u0_K7_22 ) , .A( u0_R5_15 ) , .Z( u0_u6_X_22 ) );
  XOR2_X1 u0_u6_U36 (.B( u0_K7_21 ) , .A( u0_R5_14 ) , .Z( u0_u6_X_21 ) );
  XOR2_X1 u0_u6_U37 (.B( u0_K7_20 ) , .A( u0_R5_13 ) , .Z( u0_u6_X_20 ) );
  XOR2_X1 u0_u6_U39 (.B( u0_K7_19 ) , .A( u0_R5_12 ) , .Z( u0_u6_X_19 ) );
  OAI22_X1 u0_u6_u3_U10 (.B1( u0_u6_u3_n113 ) , .A2( u0_u6_u3_n135 ) , .A1( u0_u6_u3_n150 ) , .B2( u0_u6_u3_n164 ) , .ZN( u0_u6_u3_n98 ) );
  OAI211_X1 u0_u6_u3_U11 (.B( u0_u6_u3_n106 ) , .ZN( u0_u6_u3_n119 ) , .C2( u0_u6_u3_n128 ) , .C1( u0_u6_u3_n167 ) , .A( u0_u6_u3_n181 ) );
  AOI221_X1 u0_u6_u3_U12 (.C1( u0_u6_u3_n105 ) , .ZN( u0_u6_u3_n106 ) , .A( u0_u6_u3_n131 ) , .B2( u0_u6_u3_n132 ) , .C2( u0_u6_u3_n133 ) , .B1( u0_u6_u3_n169 ) );
  INV_X1 u0_u6_u3_U13 (.ZN( u0_u6_u3_n181 ) , .A( u0_u6_u3_n98 ) );
  NAND2_X1 u0_u6_u3_U14 (.ZN( u0_u6_u3_n105 ) , .A2( u0_u6_u3_n130 ) , .A1( u0_u6_u3_n155 ) );
  NOR2_X1 u0_u6_u3_U15 (.ZN( u0_u6_u3_n126 ) , .A2( u0_u6_u3_n150 ) , .A1( u0_u6_u3_n164 ) );
  AOI21_X1 u0_u6_u3_U16 (.ZN( u0_u6_u3_n112 ) , .B2( u0_u6_u3_n146 ) , .B1( u0_u6_u3_n155 ) , .A( u0_u6_u3_n167 ) );
  NAND2_X1 u0_u6_u3_U17 (.A1( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n142 ) , .A2( u0_u6_u3_n164 ) );
  NAND2_X1 u0_u6_u3_U18 (.ZN( u0_u6_u3_n132 ) , .A2( u0_u6_u3_n152 ) , .A1( u0_u6_u3_n156 ) );
  AND2_X1 u0_u6_u3_U19 (.A2( u0_u6_u3_n113 ) , .A1( u0_u6_u3_n114 ) , .ZN( u0_u6_u3_n151 ) );
  INV_X1 u0_u6_u3_U20 (.A( u0_u6_u3_n133 ) , .ZN( u0_u6_u3_n165 ) );
  INV_X1 u0_u6_u3_U21 (.A( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n170 ) );
  NAND2_X1 u0_u6_u3_U22 (.A1( u0_u6_u3_n107 ) , .A2( u0_u6_u3_n108 ) , .ZN( u0_u6_u3_n140 ) );
  NAND2_X1 u0_u6_u3_U23 (.ZN( u0_u6_u3_n117 ) , .A1( u0_u6_u3_n124 ) , .A2( u0_u6_u3_n148 ) );
  NAND2_X1 u0_u6_u3_U24 (.ZN( u0_u6_u3_n143 ) , .A1( u0_u6_u3_n165 ) , .A2( u0_u6_u3_n167 ) );
  INV_X1 u0_u6_u3_U25 (.A( u0_u6_u3_n130 ) , .ZN( u0_u6_u3_n177 ) );
  INV_X1 u0_u6_u3_U26 (.A( u0_u6_u3_n128 ) , .ZN( u0_u6_u3_n176 ) );
  INV_X1 u0_u6_u3_U27 (.A( u0_u6_u3_n155 ) , .ZN( u0_u6_u3_n174 ) );
  AOI22_X1 u0_u6_u3_U28 (.B1( u0_u6_u3_n115 ) , .A2( u0_u6_u3_n116 ) , .ZN( u0_u6_u3_n123 ) , .B2( u0_u6_u3_n133 ) , .A1( u0_u6_u3_n169 ) );
  NAND2_X1 u0_u6_u3_U29 (.ZN( u0_u6_u3_n116 ) , .A2( u0_u6_u3_n151 ) , .A1( u0_u6_u3_n182 ) );
  INV_X1 u0_u6_u3_U3 (.A( u0_u6_u3_n129 ) , .ZN( u0_u6_u3_n183 ) );
  INV_X1 u0_u6_u3_U30 (.A( u0_u6_u3_n139 ) , .ZN( u0_u6_u3_n185 ) );
  NOR2_X1 u0_u6_u3_U31 (.ZN( u0_u6_u3_n135 ) , .A2( u0_u6_u3_n141 ) , .A1( u0_u6_u3_n169 ) );
  OAI222_X1 u0_u6_u3_U32 (.C2( u0_u6_u3_n107 ) , .A2( u0_u6_u3_n108 ) , .B1( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n138 ) , .B2( u0_u6_u3_n146 ) , .C1( u0_u6_u3_n154 ) , .A1( u0_u6_u3_n164 ) );
  NOR4_X1 u0_u6_u3_U33 (.A4( u0_u6_u3_n157 ) , .A3( u0_u6_u3_n158 ) , .A2( u0_u6_u3_n159 ) , .A1( u0_u6_u3_n160 ) , .ZN( u0_u6_u3_n161 ) );
  AOI21_X1 u0_u6_u3_U34 (.B2( u0_u6_u3_n152 ) , .B1( u0_u6_u3_n153 ) , .ZN( u0_u6_u3_n158 ) , .A( u0_u6_u3_n164 ) );
  AOI21_X1 u0_u6_u3_U35 (.A( u0_u6_u3_n154 ) , .B2( u0_u6_u3_n155 ) , .B1( u0_u6_u3_n156 ) , .ZN( u0_u6_u3_n157 ) );
  AOI21_X1 u0_u6_u3_U36 (.A( u0_u6_u3_n149 ) , .B2( u0_u6_u3_n150 ) , .B1( u0_u6_u3_n151 ) , .ZN( u0_u6_u3_n159 ) );
  AOI211_X1 u0_u6_u3_U37 (.ZN( u0_u6_u3_n109 ) , .A( u0_u6_u3_n119 ) , .C2( u0_u6_u3_n129 ) , .B( u0_u6_u3_n138 ) , .C1( u0_u6_u3_n141 ) );
  AOI211_X1 u0_u6_u3_U38 (.B( u0_u6_u3_n119 ) , .A( u0_u6_u3_n120 ) , .C2( u0_u6_u3_n121 ) , .ZN( u0_u6_u3_n122 ) , .C1( u0_u6_u3_n179 ) );
  INV_X1 u0_u6_u3_U39 (.A( u0_u6_u3_n156 ) , .ZN( u0_u6_u3_n179 ) );
  INV_X1 u0_u6_u3_U4 (.A( u0_u6_u3_n140 ) , .ZN( u0_u6_u3_n182 ) );
  OAI22_X1 u0_u6_u3_U40 (.B1( u0_u6_u3_n118 ) , .ZN( u0_u6_u3_n120 ) , .A1( u0_u6_u3_n135 ) , .B2( u0_u6_u3_n154 ) , .A2( u0_u6_u3_n178 ) );
  AND3_X1 u0_u6_u3_U41 (.ZN( u0_u6_u3_n118 ) , .A2( u0_u6_u3_n124 ) , .A1( u0_u6_u3_n144 ) , .A3( u0_u6_u3_n152 ) );
  INV_X1 u0_u6_u3_U42 (.A( u0_u6_u3_n121 ) , .ZN( u0_u6_u3_n164 ) );
  NAND2_X1 u0_u6_u3_U43 (.ZN( u0_u6_u3_n133 ) , .A1( u0_u6_u3_n154 ) , .A2( u0_u6_u3_n164 ) );
  OAI211_X1 u0_u6_u3_U44 (.B( u0_u6_u3_n127 ) , .ZN( u0_u6_u3_n139 ) , .C1( u0_u6_u3_n150 ) , .C2( u0_u6_u3_n154 ) , .A( u0_u6_u3_n184 ) );
  INV_X1 u0_u6_u3_U45 (.A( u0_u6_u3_n125 ) , .ZN( u0_u6_u3_n184 ) );
  AOI221_X1 u0_u6_u3_U46 (.A( u0_u6_u3_n126 ) , .ZN( u0_u6_u3_n127 ) , .C2( u0_u6_u3_n132 ) , .C1( u0_u6_u3_n169 ) , .B2( u0_u6_u3_n170 ) , .B1( u0_u6_u3_n174 ) );
  OAI22_X1 u0_u6_u3_U47 (.A1( u0_u6_u3_n124 ) , .ZN( u0_u6_u3_n125 ) , .B2( u0_u6_u3_n145 ) , .A2( u0_u6_u3_n165 ) , .B1( u0_u6_u3_n167 ) );
  NOR2_X1 u0_u6_u3_U48 (.A1( u0_u6_u3_n113 ) , .ZN( u0_u6_u3_n131 ) , .A2( u0_u6_u3_n154 ) );
  NAND2_X1 u0_u6_u3_U49 (.A1( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n150 ) , .A2( u0_u6_u3_n99 ) );
  INV_X1 u0_u6_u3_U5 (.A( u0_u6_u3_n117 ) , .ZN( u0_u6_u3_n178 ) );
  NAND2_X1 u0_u6_u3_U50 (.A2( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n155 ) , .A1( u0_u6_u3_n97 ) );
  INV_X1 u0_u6_u3_U51 (.A( u0_u6_u3_n141 ) , .ZN( u0_u6_u3_n167 ) );
  AOI21_X1 u0_u6_u3_U52 (.B2( u0_u6_u3_n114 ) , .B1( u0_u6_u3_n146 ) , .A( u0_u6_u3_n154 ) , .ZN( u0_u6_u3_n94 ) );
  AOI21_X1 u0_u6_u3_U53 (.ZN( u0_u6_u3_n110 ) , .B2( u0_u6_u3_n142 ) , .B1( u0_u6_u3_n186 ) , .A( u0_u6_u3_n95 ) );
  INV_X1 u0_u6_u3_U54 (.A( u0_u6_u3_n145 ) , .ZN( u0_u6_u3_n186 ) );
  AOI21_X1 u0_u6_u3_U55 (.B1( u0_u6_u3_n124 ) , .A( u0_u6_u3_n149 ) , .B2( u0_u6_u3_n155 ) , .ZN( u0_u6_u3_n95 ) );
  INV_X1 u0_u6_u3_U56 (.A( u0_u6_u3_n149 ) , .ZN( u0_u6_u3_n169 ) );
  NAND2_X1 u0_u6_u3_U57 (.ZN( u0_u6_u3_n124 ) , .A1( u0_u6_u3_n96 ) , .A2( u0_u6_u3_n97 ) );
  NAND2_X1 u0_u6_u3_U58 (.A2( u0_u6_u3_n100 ) , .ZN( u0_u6_u3_n146 ) , .A1( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U59 (.A1( u0_u6_u3_n101 ) , .ZN( u0_u6_u3_n145 ) , .A2( u0_u6_u3_n99 ) );
  AOI221_X1 u0_u6_u3_U6 (.A( u0_u6_u3_n131 ) , .C2( u0_u6_u3_n132 ) , .C1( u0_u6_u3_n133 ) , .ZN( u0_u6_u3_n134 ) , .B1( u0_u6_u3_n143 ) , .B2( u0_u6_u3_n177 ) );
  NAND2_X1 u0_u6_u3_U60 (.A1( u0_u6_u3_n100 ) , .ZN( u0_u6_u3_n156 ) , .A2( u0_u6_u3_n99 ) );
  NAND2_X1 u0_u6_u3_U61 (.A2( u0_u6_u3_n101 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n148 ) );
  NAND2_X1 u0_u6_u3_U62 (.A1( u0_u6_u3_n100 ) , .A2( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n128 ) );
  NAND2_X1 u0_u6_u3_U63 (.A2( u0_u6_u3_n101 ) , .A1( u0_u6_u3_n102 ) , .ZN( u0_u6_u3_n152 ) );
  NAND2_X1 u0_u6_u3_U64 (.A2( u0_u6_u3_n101 ) , .ZN( u0_u6_u3_n114 ) , .A1( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U65 (.ZN( u0_u6_u3_n107 ) , .A1( u0_u6_u3_n97 ) , .A2( u0_u6_u3_n99 ) );
  NAND2_X1 u0_u6_u3_U66 (.A2( u0_u6_u3_n100 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n113 ) );
  NAND2_X1 u0_u6_u3_U67 (.A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n153 ) , .A2( u0_u6_u3_n97 ) );
  NAND2_X1 u0_u6_u3_U68 (.A2( u0_u6_u3_n103 ) , .A1( u0_u6_u3_n104 ) , .ZN( u0_u6_u3_n130 ) );
  NAND2_X1 u0_u6_u3_U69 (.A2( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n144 ) , .A1( u0_u6_u3_n96 ) );
  OAI22_X1 u0_u6_u3_U7 (.B2( u0_u6_u3_n147 ) , .A2( u0_u6_u3_n148 ) , .ZN( u0_u6_u3_n160 ) , .B1( u0_u6_u3_n165 ) , .A1( u0_u6_u3_n168 ) );
  NAND2_X1 u0_u6_u3_U70 (.A1( u0_u6_u3_n102 ) , .A2( u0_u6_u3_n103 ) , .ZN( u0_u6_u3_n108 ) );
  NOR2_X1 u0_u6_u3_U71 (.A2( u0_u6_X_19 ) , .A1( u0_u6_X_20 ) , .ZN( u0_u6_u3_n99 ) );
  NOR2_X1 u0_u6_u3_U72 (.A2( u0_u6_X_21 ) , .A1( u0_u6_X_24 ) , .ZN( u0_u6_u3_n103 ) );
  NOR2_X1 u0_u6_u3_U73 (.A2( u0_u6_X_24 ) , .A1( u0_u6_u3_n171 ) , .ZN( u0_u6_u3_n97 ) );
  NOR2_X1 u0_u6_u3_U74 (.A2( u0_u6_X_23 ) , .ZN( u0_u6_u3_n141 ) , .A1( u0_u6_u3_n166 ) );
  NOR2_X1 u0_u6_u3_U75 (.A2( u0_u6_X_19 ) , .A1( u0_u6_u3_n172 ) , .ZN( u0_u6_u3_n96 ) );
  NAND2_X1 u0_u6_u3_U76 (.A1( u0_u6_X_22 ) , .A2( u0_u6_X_23 ) , .ZN( u0_u6_u3_n154 ) );
  NAND2_X1 u0_u6_u3_U77 (.A1( u0_u6_X_23 ) , .ZN( u0_u6_u3_n149 ) , .A2( u0_u6_u3_n166 ) );
  NOR2_X1 u0_u6_u3_U78 (.A2( u0_u6_X_22 ) , .A1( u0_u6_X_23 ) , .ZN( u0_u6_u3_n121 ) );
  AND2_X1 u0_u6_u3_U79 (.A1( u0_u6_X_24 ) , .ZN( u0_u6_u3_n101 ) , .A2( u0_u6_u3_n171 ) );
  AND3_X1 u0_u6_u3_U8 (.A3( u0_u6_u3_n144 ) , .A2( u0_u6_u3_n145 ) , .A1( u0_u6_u3_n146 ) , .ZN( u0_u6_u3_n147 ) );
  AND2_X1 u0_u6_u3_U80 (.A1( u0_u6_X_19 ) , .ZN( u0_u6_u3_n102 ) , .A2( u0_u6_u3_n172 ) );
  AND2_X1 u0_u6_u3_U81 (.A1( u0_u6_X_21 ) , .A2( u0_u6_X_24 ) , .ZN( u0_u6_u3_n100 ) );
  AND2_X1 u0_u6_u3_U82 (.A2( u0_u6_X_19 ) , .A1( u0_u6_X_20 ) , .ZN( u0_u6_u3_n104 ) );
  INV_X1 u0_u6_u3_U83 (.A( u0_u6_X_22 ) , .ZN( u0_u6_u3_n166 ) );
  INV_X1 u0_u6_u3_U84 (.A( u0_u6_X_21 ) , .ZN( u0_u6_u3_n171 ) );
  INV_X1 u0_u6_u3_U85 (.A( u0_u6_X_20 ) , .ZN( u0_u6_u3_n172 ) );
  NAND4_X1 u0_u6_u3_U86 (.ZN( u0_out6_26 ) , .A4( u0_u6_u3_n109 ) , .A3( u0_u6_u3_n110 ) , .A2( u0_u6_u3_n111 ) , .A1( u0_u6_u3_n173 ) );
  INV_X1 u0_u6_u3_U87 (.ZN( u0_u6_u3_n173 ) , .A( u0_u6_u3_n94 ) );
  OAI21_X1 u0_u6_u3_U88 (.ZN( u0_u6_u3_n111 ) , .B2( u0_u6_u3_n117 ) , .A( u0_u6_u3_n133 ) , .B1( u0_u6_u3_n176 ) );
  NAND4_X1 u0_u6_u3_U89 (.ZN( u0_out6_20 ) , .A4( u0_u6_u3_n122 ) , .A3( u0_u6_u3_n123 ) , .A1( u0_u6_u3_n175 ) , .A2( u0_u6_u3_n180 ) );
  INV_X1 u0_u6_u3_U9 (.A( u0_u6_u3_n143 ) , .ZN( u0_u6_u3_n168 ) );
  INV_X1 u0_u6_u3_U90 (.A( u0_u6_u3_n126 ) , .ZN( u0_u6_u3_n180 ) );
  INV_X1 u0_u6_u3_U91 (.A( u0_u6_u3_n112 ) , .ZN( u0_u6_u3_n175 ) );
  NAND4_X1 u0_u6_u3_U92 (.ZN( u0_out6_1 ) , .A4( u0_u6_u3_n161 ) , .A3( u0_u6_u3_n162 ) , .A2( u0_u6_u3_n163 ) , .A1( u0_u6_u3_n185 ) );
  NAND2_X1 u0_u6_u3_U93 (.ZN( u0_u6_u3_n163 ) , .A2( u0_u6_u3_n170 ) , .A1( u0_u6_u3_n176 ) );
  AOI22_X1 u0_u6_u3_U94 (.B2( u0_u6_u3_n140 ) , .B1( u0_u6_u3_n141 ) , .A2( u0_u6_u3_n142 ) , .ZN( u0_u6_u3_n162 ) , .A1( u0_u6_u3_n177 ) );
  OR4_X1 u0_u6_u3_U95 (.ZN( u0_out6_10 ) , .A4( u0_u6_u3_n136 ) , .A3( u0_u6_u3_n137 ) , .A1( u0_u6_u3_n138 ) , .A2( u0_u6_u3_n139 ) );
  OAI222_X1 u0_u6_u3_U96 (.C1( u0_u6_u3_n128 ) , .ZN( u0_u6_u3_n137 ) , .B1( u0_u6_u3_n148 ) , .A2( u0_u6_u3_n150 ) , .B2( u0_u6_u3_n154 ) , .C2( u0_u6_u3_n164 ) , .A1( u0_u6_u3_n167 ) );
  OAI221_X1 u0_u6_u3_U97 (.A( u0_u6_u3_n134 ) , .B2( u0_u6_u3_n135 ) , .ZN( u0_u6_u3_n136 ) , .C1( u0_u6_u3_n149 ) , .B1( u0_u6_u3_n151 ) , .C2( u0_u6_u3_n183 ) );
  NAND3_X1 u0_u6_u3_U98 (.A1( u0_u6_u3_n114 ) , .ZN( u0_u6_u3_n115 ) , .A2( u0_u6_u3_n145 ) , .A3( u0_u6_u3_n153 ) );
  NAND3_X1 u0_u6_u3_U99 (.ZN( u0_u6_u3_n129 ) , .A2( u0_u6_u3_n144 ) , .A1( u0_u6_u3_n153 ) , .A3( u0_u6_u3_n182 ) );
  OAI22_X1 u0_u6_u4_U10 (.B2( u0_u6_u4_n135 ) , .ZN( u0_u6_u4_n137 ) , .B1( u0_u6_u4_n153 ) , .A1( u0_u6_u4_n155 ) , .A2( u0_u6_u4_n171 ) );
  AND3_X1 u0_u6_u4_U11 (.A2( u0_u6_u4_n134 ) , .ZN( u0_u6_u4_n135 ) , .A3( u0_u6_u4_n145 ) , .A1( u0_u6_u4_n157 ) );
  NAND2_X1 u0_u6_u4_U12 (.ZN( u0_u6_u4_n132 ) , .A2( u0_u6_u4_n170 ) , .A1( u0_u6_u4_n173 ) );
  AOI21_X1 u0_u6_u4_U13 (.B2( u0_u6_u4_n160 ) , .B1( u0_u6_u4_n161 ) , .ZN( u0_u6_u4_n162 ) , .A( u0_u6_u4_n170 ) );
  AOI21_X1 u0_u6_u4_U14 (.ZN( u0_u6_u4_n107 ) , .B2( u0_u6_u4_n143 ) , .A( u0_u6_u4_n174 ) , .B1( u0_u6_u4_n184 ) );
  AOI21_X1 u0_u6_u4_U15 (.B2( u0_u6_u4_n158 ) , .B1( u0_u6_u4_n159 ) , .ZN( u0_u6_u4_n163 ) , .A( u0_u6_u4_n174 ) );
  AOI21_X1 u0_u6_u4_U16 (.A( u0_u6_u4_n153 ) , .B2( u0_u6_u4_n154 ) , .B1( u0_u6_u4_n155 ) , .ZN( u0_u6_u4_n165 ) );
  AOI21_X1 u0_u6_u4_U17 (.A( u0_u6_u4_n156 ) , .B2( u0_u6_u4_n157 ) , .ZN( u0_u6_u4_n164 ) , .B1( u0_u6_u4_n184 ) );
  INV_X1 u0_u6_u4_U18 (.A( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n170 ) );
  AND2_X1 u0_u6_u4_U19 (.A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n155 ) , .A1( u0_u6_u4_n160 ) );
  INV_X1 u0_u6_u4_U20 (.A( u0_u6_u4_n156 ) , .ZN( u0_u6_u4_n175 ) );
  NAND2_X1 u0_u6_u4_U21 (.A2( u0_u6_u4_n118 ) , .ZN( u0_u6_u4_n131 ) , .A1( u0_u6_u4_n147 ) );
  NAND2_X1 u0_u6_u4_U22 (.A1( u0_u6_u4_n119 ) , .A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n130 ) );
  NAND2_X1 u0_u6_u4_U23 (.ZN( u0_u6_u4_n117 ) , .A2( u0_u6_u4_n118 ) , .A1( u0_u6_u4_n148 ) );
  NAND2_X1 u0_u6_u4_U24 (.ZN( u0_u6_u4_n129 ) , .A1( u0_u6_u4_n134 ) , .A2( u0_u6_u4_n148 ) );
  AND3_X1 u0_u6_u4_U25 (.A1( u0_u6_u4_n119 ) , .A2( u0_u6_u4_n143 ) , .A3( u0_u6_u4_n154 ) , .ZN( u0_u6_u4_n161 ) );
  AND2_X1 u0_u6_u4_U26 (.A1( u0_u6_u4_n145 ) , .A2( u0_u6_u4_n147 ) , .ZN( u0_u6_u4_n159 ) );
  OR3_X1 u0_u6_u4_U27 (.A3( u0_u6_u4_n114 ) , .A2( u0_u6_u4_n115 ) , .A1( u0_u6_u4_n116 ) , .ZN( u0_u6_u4_n136 ) );
  AOI21_X1 u0_u6_u4_U28 (.A( u0_u6_u4_n113 ) , .ZN( u0_u6_u4_n116 ) , .B2( u0_u6_u4_n173 ) , .B1( u0_u6_u4_n174 ) );
  AOI21_X1 u0_u6_u4_U29 (.ZN( u0_u6_u4_n115 ) , .B2( u0_u6_u4_n145 ) , .B1( u0_u6_u4_n146 ) , .A( u0_u6_u4_n156 ) );
  NOR2_X1 u0_u6_u4_U3 (.ZN( u0_u6_u4_n121 ) , .A1( u0_u6_u4_n181 ) , .A2( u0_u6_u4_n182 ) );
  OAI22_X1 u0_u6_u4_U30 (.ZN( u0_u6_u4_n114 ) , .A2( u0_u6_u4_n121 ) , .B1( u0_u6_u4_n160 ) , .B2( u0_u6_u4_n170 ) , .A1( u0_u6_u4_n171 ) );
  INV_X1 u0_u6_u4_U31 (.A( u0_u6_u4_n158 ) , .ZN( u0_u6_u4_n182 ) );
  INV_X1 u0_u6_u4_U32 (.ZN( u0_u6_u4_n181 ) , .A( u0_u6_u4_n96 ) );
  INV_X1 u0_u6_u4_U33 (.A( u0_u6_u4_n144 ) , .ZN( u0_u6_u4_n179 ) );
  INV_X1 u0_u6_u4_U34 (.A( u0_u6_u4_n157 ) , .ZN( u0_u6_u4_n178 ) );
  NAND2_X1 u0_u6_u4_U35 (.A2( u0_u6_u4_n154 ) , .A1( u0_u6_u4_n96 ) , .ZN( u0_u6_u4_n97 ) );
  INV_X1 u0_u6_u4_U36 (.ZN( u0_u6_u4_n186 ) , .A( u0_u6_u4_n95 ) );
  OAI221_X1 u0_u6_u4_U37 (.C1( u0_u6_u4_n134 ) , .B1( u0_u6_u4_n158 ) , .B2( u0_u6_u4_n171 ) , .C2( u0_u6_u4_n173 ) , .A( u0_u6_u4_n94 ) , .ZN( u0_u6_u4_n95 ) );
  AOI222_X1 u0_u6_u4_U38 (.B2( u0_u6_u4_n132 ) , .A1( u0_u6_u4_n138 ) , .C2( u0_u6_u4_n175 ) , .A2( u0_u6_u4_n179 ) , .C1( u0_u6_u4_n181 ) , .B1( u0_u6_u4_n185 ) , .ZN( u0_u6_u4_n94 ) );
  INV_X1 u0_u6_u4_U39 (.A( u0_u6_u4_n113 ) , .ZN( u0_u6_u4_n185 ) );
  INV_X1 u0_u6_u4_U4 (.A( u0_u6_u4_n117 ) , .ZN( u0_u6_u4_n184 ) );
  INV_X1 u0_u6_u4_U40 (.A( u0_u6_u4_n143 ) , .ZN( u0_u6_u4_n183 ) );
  NOR2_X1 u0_u6_u4_U41 (.ZN( u0_u6_u4_n138 ) , .A1( u0_u6_u4_n168 ) , .A2( u0_u6_u4_n169 ) );
  NOR2_X1 u0_u6_u4_U42 (.A1( u0_u6_u4_n150 ) , .A2( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n153 ) );
  NOR2_X1 u0_u6_u4_U43 (.A2( u0_u6_u4_n128 ) , .A1( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n156 ) );
  AOI22_X1 u0_u6_u4_U44 (.B2( u0_u6_u4_n122 ) , .A1( u0_u6_u4_n123 ) , .ZN( u0_u6_u4_n124 ) , .B1( u0_u6_u4_n128 ) , .A2( u0_u6_u4_n172 ) );
  INV_X1 u0_u6_u4_U45 (.A( u0_u6_u4_n153 ) , .ZN( u0_u6_u4_n172 ) );
  NAND2_X1 u0_u6_u4_U46 (.A2( u0_u6_u4_n120 ) , .ZN( u0_u6_u4_n123 ) , .A1( u0_u6_u4_n161 ) );
  AOI22_X1 u0_u6_u4_U47 (.B2( u0_u6_u4_n132 ) , .A2( u0_u6_u4_n133 ) , .ZN( u0_u6_u4_n140 ) , .A1( u0_u6_u4_n150 ) , .B1( u0_u6_u4_n179 ) );
  NAND2_X1 u0_u6_u4_U48 (.ZN( u0_u6_u4_n133 ) , .A2( u0_u6_u4_n146 ) , .A1( u0_u6_u4_n154 ) );
  NAND2_X1 u0_u6_u4_U49 (.A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n154 ) , .A2( u0_u6_u4_n98 ) );
  NOR4_X1 u0_u6_u4_U5 (.A4( u0_u6_u4_n106 ) , .A3( u0_u6_u4_n107 ) , .A2( u0_u6_u4_n108 ) , .A1( u0_u6_u4_n109 ) , .ZN( u0_u6_u4_n110 ) );
  NAND2_X1 u0_u6_u4_U50 (.A1( u0_u6_u4_n101 ) , .ZN( u0_u6_u4_n158 ) , .A2( u0_u6_u4_n99 ) );
  AOI21_X1 u0_u6_u4_U51 (.ZN( u0_u6_u4_n127 ) , .A( u0_u6_u4_n136 ) , .B2( u0_u6_u4_n150 ) , .B1( u0_u6_u4_n180 ) );
  INV_X1 u0_u6_u4_U52 (.A( u0_u6_u4_n160 ) , .ZN( u0_u6_u4_n180 ) );
  NAND2_X1 u0_u6_u4_U53 (.A2( u0_u6_u4_n104 ) , .A1( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n146 ) );
  NAND2_X1 u0_u6_u4_U54 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n160 ) );
  NAND2_X1 u0_u6_u4_U55 (.ZN( u0_u6_u4_n134 ) , .A1( u0_u6_u4_n98 ) , .A2( u0_u6_u4_n99 ) );
  NAND2_X1 u0_u6_u4_U56 (.A1( u0_u6_u4_n103 ) , .A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n143 ) );
  NAND2_X1 u0_u6_u4_U57 (.A2( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n145 ) , .A1( u0_u6_u4_n98 ) );
  NAND2_X1 u0_u6_u4_U58 (.A1( u0_u6_u4_n100 ) , .A2( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n120 ) );
  NAND2_X1 u0_u6_u4_U59 (.A1( u0_u6_u4_n102 ) , .A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n148 ) );
  AOI21_X1 u0_u6_u4_U6 (.ZN( u0_u6_u4_n106 ) , .B2( u0_u6_u4_n146 ) , .B1( u0_u6_u4_n158 ) , .A( u0_u6_u4_n170 ) );
  NAND2_X1 u0_u6_u4_U60 (.A2( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n157 ) );
  INV_X1 u0_u6_u4_U61 (.A( u0_u6_u4_n150 ) , .ZN( u0_u6_u4_n173 ) );
  INV_X1 u0_u6_u4_U62 (.A( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n171 ) );
  NAND2_X1 u0_u6_u4_U63 (.A1( u0_u6_u4_n100 ) , .ZN( u0_u6_u4_n118 ) , .A2( u0_u6_u4_n99 ) );
  NAND2_X1 u0_u6_u4_U64 (.A2( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n144 ) );
  NAND2_X1 u0_u6_u4_U65 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n105 ) , .ZN( u0_u6_u4_n96 ) );
  INV_X1 u0_u6_u4_U66 (.A( u0_u6_u4_n128 ) , .ZN( u0_u6_u4_n174 ) );
  NAND2_X1 u0_u6_u4_U67 (.A2( u0_u6_u4_n102 ) , .ZN( u0_u6_u4_n119 ) , .A1( u0_u6_u4_n98 ) );
  NAND2_X1 u0_u6_u4_U68 (.A2( u0_u6_u4_n101 ) , .A1( u0_u6_u4_n103 ) , .ZN( u0_u6_u4_n147 ) );
  NAND2_X1 u0_u6_u4_U69 (.A2( u0_u6_u4_n104 ) , .ZN( u0_u6_u4_n113 ) , .A1( u0_u6_u4_n99 ) );
  AOI21_X1 u0_u6_u4_U7 (.ZN( u0_u6_u4_n108 ) , .B2( u0_u6_u4_n134 ) , .B1( u0_u6_u4_n155 ) , .A( u0_u6_u4_n156 ) );
  NOR2_X1 u0_u6_u4_U70 (.A2( u0_u6_X_28 ) , .ZN( u0_u6_u4_n150 ) , .A1( u0_u6_u4_n168 ) );
  NOR2_X1 u0_u6_u4_U71 (.A2( u0_u6_X_29 ) , .ZN( u0_u6_u4_n152 ) , .A1( u0_u6_u4_n169 ) );
  NOR2_X1 u0_u6_u4_U72 (.A2( u0_u6_X_30 ) , .ZN( u0_u6_u4_n105 ) , .A1( u0_u6_u4_n176 ) );
  NOR2_X1 u0_u6_u4_U73 (.A2( u0_u6_X_26 ) , .ZN( u0_u6_u4_n100 ) , .A1( u0_u6_u4_n177 ) );
  NOR2_X1 u0_u6_u4_U74 (.A2( u0_u6_X_28 ) , .A1( u0_u6_X_29 ) , .ZN( u0_u6_u4_n128 ) );
  NOR2_X1 u0_u6_u4_U75 (.A2( u0_u6_X_27 ) , .A1( u0_u6_X_30 ) , .ZN( u0_u6_u4_n102 ) );
  NOR2_X1 u0_u6_u4_U76 (.A2( u0_u6_X_25 ) , .A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n98 ) );
  AND2_X1 u0_u6_u4_U77 (.A2( u0_u6_X_25 ) , .A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n104 ) );
  AND2_X1 u0_u6_u4_U78 (.A1( u0_u6_X_30 ) , .A2( u0_u6_u4_n176 ) , .ZN( u0_u6_u4_n99 ) );
  AND2_X1 u0_u6_u4_U79 (.A1( u0_u6_X_26 ) , .ZN( u0_u6_u4_n101 ) , .A2( u0_u6_u4_n177 ) );
  AOI21_X1 u0_u6_u4_U8 (.ZN( u0_u6_u4_n109 ) , .A( u0_u6_u4_n153 ) , .B1( u0_u6_u4_n159 ) , .B2( u0_u6_u4_n184 ) );
  AND2_X1 u0_u6_u4_U80 (.A1( u0_u6_X_27 ) , .A2( u0_u6_X_30 ) , .ZN( u0_u6_u4_n103 ) );
  INV_X1 u0_u6_u4_U81 (.A( u0_u6_X_28 ) , .ZN( u0_u6_u4_n169 ) );
  INV_X1 u0_u6_u4_U82 (.A( u0_u6_X_29 ) , .ZN( u0_u6_u4_n168 ) );
  INV_X1 u0_u6_u4_U83 (.A( u0_u6_X_25 ) , .ZN( u0_u6_u4_n177 ) );
  INV_X1 u0_u6_u4_U84 (.A( u0_u6_X_27 ) , .ZN( u0_u6_u4_n176 ) );
  NAND4_X1 u0_u6_u4_U85 (.ZN( u0_out6_25 ) , .A4( u0_u6_u4_n139 ) , .A3( u0_u6_u4_n140 ) , .A2( u0_u6_u4_n141 ) , .A1( u0_u6_u4_n142 ) );
  OAI21_X1 u0_u6_u4_U86 (.B2( u0_u6_u4_n131 ) , .ZN( u0_u6_u4_n141 ) , .A( u0_u6_u4_n175 ) , .B1( u0_u6_u4_n183 ) );
  OAI21_X1 u0_u6_u4_U87 (.A( u0_u6_u4_n128 ) , .B2( u0_u6_u4_n129 ) , .B1( u0_u6_u4_n130 ) , .ZN( u0_u6_u4_n142 ) );
  NAND4_X1 u0_u6_u4_U88 (.ZN( u0_out6_14 ) , .A4( u0_u6_u4_n124 ) , .A3( u0_u6_u4_n125 ) , .A2( u0_u6_u4_n126 ) , .A1( u0_u6_u4_n127 ) );
  AOI22_X1 u0_u6_u4_U89 (.B2( u0_u6_u4_n117 ) , .ZN( u0_u6_u4_n126 ) , .A1( u0_u6_u4_n129 ) , .B1( u0_u6_u4_n152 ) , .A2( u0_u6_u4_n175 ) );
  AOI211_X1 u0_u6_u4_U9 (.B( u0_u6_u4_n136 ) , .A( u0_u6_u4_n137 ) , .C2( u0_u6_u4_n138 ) , .ZN( u0_u6_u4_n139 ) , .C1( u0_u6_u4_n182 ) );
  AOI22_X1 u0_u6_u4_U90 (.ZN( u0_u6_u4_n125 ) , .B2( u0_u6_u4_n131 ) , .A2( u0_u6_u4_n132 ) , .B1( u0_u6_u4_n138 ) , .A1( u0_u6_u4_n178 ) );
  NAND4_X1 u0_u6_u4_U91 (.ZN( u0_out6_8 ) , .A4( u0_u6_u4_n110 ) , .A3( u0_u6_u4_n111 ) , .A2( u0_u6_u4_n112 ) , .A1( u0_u6_u4_n186 ) );
  NAND2_X1 u0_u6_u4_U92 (.ZN( u0_u6_u4_n112 ) , .A2( u0_u6_u4_n130 ) , .A1( u0_u6_u4_n150 ) );
  AOI22_X1 u0_u6_u4_U93 (.ZN( u0_u6_u4_n111 ) , .B2( u0_u6_u4_n132 ) , .A1( u0_u6_u4_n152 ) , .B1( u0_u6_u4_n178 ) , .A2( u0_u6_u4_n97 ) );
  AOI22_X1 u0_u6_u4_U94 (.B2( u0_u6_u4_n149 ) , .B1( u0_u6_u4_n150 ) , .A2( u0_u6_u4_n151 ) , .A1( u0_u6_u4_n152 ) , .ZN( u0_u6_u4_n167 ) );
  NOR4_X1 u0_u6_u4_U95 (.A4( u0_u6_u4_n162 ) , .A3( u0_u6_u4_n163 ) , .A2( u0_u6_u4_n164 ) , .A1( u0_u6_u4_n165 ) , .ZN( u0_u6_u4_n166 ) );
  NAND3_X1 u0_u6_u4_U96 (.ZN( u0_out6_3 ) , .A3( u0_u6_u4_n166 ) , .A1( u0_u6_u4_n167 ) , .A2( u0_u6_u4_n186 ) );
  NAND3_X1 u0_u6_u4_U97 (.A3( u0_u6_u4_n146 ) , .A2( u0_u6_u4_n147 ) , .A1( u0_u6_u4_n148 ) , .ZN( u0_u6_u4_n149 ) );
  NAND3_X1 u0_u6_u4_U98 (.A3( u0_u6_u4_n143 ) , .A2( u0_u6_u4_n144 ) , .A1( u0_u6_u4_n145 ) , .ZN( u0_u6_u4_n151 ) );
  NAND3_X1 u0_u6_u4_U99 (.A3( u0_u6_u4_n121 ) , .ZN( u0_u6_u4_n122 ) , .A2( u0_u6_u4_n144 ) , .A1( u0_u6_u4_n154 ) );
  XOR2_X1 u0_u8_U1 (.B( u0_K9_9 ) , .A( u0_R7_6 ) , .Z( u0_u8_X_9 ) );
  XOR2_X1 u0_u8_U10 (.B( u0_K9_45 ) , .A( u0_R7_30 ) , .Z( u0_u8_X_45 ) );
  XOR2_X1 u0_u8_U11 (.B( u0_K9_44 ) , .A( u0_R7_29 ) , .Z( u0_u8_X_44 ) );
  XOR2_X1 u0_u8_U12 (.B( u0_K9_43 ) , .A( u0_R7_28 ) , .Z( u0_u8_X_43 ) );
  XOR2_X1 u0_u8_U16 (.B( u0_K9_3 ) , .A( u0_R7_2 ) , .Z( u0_u8_X_3 ) );
  XOR2_X1 u0_u8_U2 (.B( u0_K9_8 ) , .A( u0_R7_5 ) , .Z( u0_u8_X_8 ) );
  XOR2_X1 u0_u8_U26 (.B( u0_K9_30 ) , .A( u0_R7_21 ) , .Z( u0_u8_X_30 ) );
  XOR2_X1 u0_u8_U27 (.B( u0_K9_2 ) , .A( u0_R7_1 ) , .Z( u0_u8_X_2 ) );
  XOR2_X1 u0_u8_U28 (.B( u0_K9_29 ) , .A( u0_R7_20 ) , .Z( u0_u8_X_29 ) );
  XOR2_X1 u0_u8_U29 (.B( u0_K9_28 ) , .A( u0_R7_19 ) , .Z( u0_u8_X_28 ) );
  XOR2_X1 u0_u8_U3 (.B( u0_K9_7 ) , .A( u0_R7_4 ) , .Z( u0_u8_X_7 ) );
  XOR2_X1 u0_u8_U30 (.B( u0_K9_27 ) , .A( u0_R7_18 ) , .Z( u0_u8_X_27 ) );
  XOR2_X1 u0_u8_U31 (.B( u0_K9_26 ) , .A( u0_R7_17 ) , .Z( u0_u8_X_26 ) );
  XOR2_X1 u0_u8_U32 (.B( u0_K9_25 ) , .A( u0_R7_16 ) , .Z( u0_u8_X_25 ) );
  XOR2_X1 u0_u8_U33 (.B( u0_K9_24 ) , .A( u0_R7_17 ) , .Z( u0_u8_X_24 ) );
  XOR2_X1 u0_u8_U34 (.B( u0_K9_23 ) , .A( u0_R7_16 ) , .Z( u0_u8_X_23 ) );
  XOR2_X1 u0_u8_U35 (.B( u0_K9_22 ) , .A( u0_R7_15 ) , .Z( u0_u8_X_22 ) );
  XOR2_X1 u0_u8_U36 (.B( u0_K9_21 ) , .A( u0_R7_14 ) , .Z( u0_u8_X_21 ) );
  XOR2_X1 u0_u8_U37 (.B( u0_K9_20 ) , .A( u0_R7_13 ) , .Z( u0_u8_X_20 ) );
  XOR2_X1 u0_u8_U38 (.B( u0_K9_1 ) , .A( u0_R7_32 ) , .Z( u0_u8_X_1 ) );
  XOR2_X1 u0_u8_U39 (.B( u0_K9_19 ) , .A( u0_R7_12 ) , .Z( u0_u8_X_19 ) );
  XOR2_X1 u0_u8_U4 (.B( u0_K9_6 ) , .A( u0_R7_5 ) , .Z( u0_u8_X_6 ) );
  XOR2_X1 u0_u8_U40 (.B( u0_K9_18 ) , .A( u0_R7_13 ) , .Z( u0_u8_X_18 ) );
  XOR2_X1 u0_u8_U41 (.B( u0_K9_17 ) , .A( u0_R7_12 ) , .Z( u0_u8_X_17 ) );
  XOR2_X1 u0_u8_U42 (.B( u0_K9_16 ) , .A( u0_R7_11 ) , .Z( u0_u8_X_16 ) );
  XOR2_X1 u0_u8_U43 (.B( u0_K9_15 ) , .A( u0_R7_10 ) , .Z( u0_u8_X_15 ) );
  XOR2_X1 u0_u8_U44 (.B( u0_K9_14 ) , .A( u0_R7_9 ) , .Z( u0_u8_X_14 ) );
  XOR2_X1 u0_u8_U45 (.B( u0_K9_13 ) , .A( u0_R7_8 ) , .Z( u0_u8_X_13 ) );
  XOR2_X1 u0_u8_U46 (.B( u0_K9_12 ) , .A( u0_R7_9 ) , .Z( u0_u8_X_12 ) );
  XOR2_X1 u0_u8_U47 (.B( u0_K9_11 ) , .A( u0_R7_8 ) , .Z( u0_u8_X_11 ) );
  XOR2_X1 u0_u8_U48 (.B( u0_K9_10 ) , .A( u0_R7_7 ) , .Z( u0_u8_X_10 ) );
  XOR2_X1 u0_u8_U5 (.B( u0_K9_5 ) , .A( u0_R7_4 ) , .Z( u0_u8_X_5 ) );
  XOR2_X1 u0_u8_U6 (.B( u0_K9_4 ) , .A( u0_R7_3 ) , .Z( u0_u8_X_4 ) );
  XOR2_X1 u0_u8_U7 (.B( u0_K9_48 ) , .A( u0_R7_1 ) , .Z( u0_u8_X_48 ) );
  XOR2_X1 u0_u8_U8 (.B( u0_K9_47 ) , .A( u0_R7_32 ) , .Z( u0_u8_X_47 ) );
  XOR2_X1 u0_u8_U9 (.B( u0_K9_46 ) , .A( u0_R7_31 ) , .Z( u0_u8_X_46 ) );
  AND3_X1 u0_u8_u0_U10 (.A2( u0_u8_u0_n112 ) , .ZN( u0_u8_u0_n127 ) , .A3( u0_u8_u0_n130 ) , .A1( u0_u8_u0_n148 ) );
  NAND2_X1 u0_u8_u0_U11 (.ZN( u0_u8_u0_n113 ) , .A1( u0_u8_u0_n139 ) , .A2( u0_u8_u0_n149 ) );
  AND2_X1 u0_u8_u0_U12 (.ZN( u0_u8_u0_n107 ) , .A1( u0_u8_u0_n130 ) , .A2( u0_u8_u0_n140 ) );
  AND2_X1 u0_u8_u0_U13 (.A2( u0_u8_u0_n129 ) , .A1( u0_u8_u0_n130 ) , .ZN( u0_u8_u0_n151 ) );
  AND2_X1 u0_u8_u0_U14 (.A1( u0_u8_u0_n108 ) , .A2( u0_u8_u0_n125 ) , .ZN( u0_u8_u0_n145 ) );
  INV_X1 u0_u8_u0_U15 (.A( u0_u8_u0_n143 ) , .ZN( u0_u8_u0_n173 ) );
  NOR2_X1 u0_u8_u0_U16 (.A2( u0_u8_u0_n136 ) , .ZN( u0_u8_u0_n147 ) , .A1( u0_u8_u0_n160 ) );
  AOI21_X1 u0_u8_u0_U17 (.B1( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n132 ) , .A( u0_u8_u0_n165 ) , .B2( u0_u8_u0_n93 ) );
  INV_X1 u0_u8_u0_U18 (.A( u0_u8_u0_n142 ) , .ZN( u0_u8_u0_n165 ) );
  OAI22_X1 u0_u8_u0_U19 (.B1( u0_u8_u0_n125 ) , .ZN( u0_u8_u0_n126 ) , .A1( u0_u8_u0_n138 ) , .A2( u0_u8_u0_n146 ) , .B2( u0_u8_u0_n147 ) );
  OAI22_X1 u0_u8_u0_U20 (.B1( u0_u8_u0_n131 ) , .A1( u0_u8_u0_n144 ) , .B2( u0_u8_u0_n147 ) , .A2( u0_u8_u0_n90 ) , .ZN( u0_u8_u0_n91 ) );
  AND3_X1 u0_u8_u0_U21 (.A3( u0_u8_u0_n121 ) , .A2( u0_u8_u0_n125 ) , .A1( u0_u8_u0_n148 ) , .ZN( u0_u8_u0_n90 ) );
  INV_X1 u0_u8_u0_U22 (.A( u0_u8_u0_n136 ) , .ZN( u0_u8_u0_n161 ) );
  AOI22_X1 u0_u8_u0_U23 (.B2( u0_u8_u0_n109 ) , .A2( u0_u8_u0_n110 ) , .ZN( u0_u8_u0_n111 ) , .B1( u0_u8_u0_n118 ) , .A1( u0_u8_u0_n160 ) );
  INV_X1 u0_u8_u0_U24 (.A( u0_u8_u0_n118 ) , .ZN( u0_u8_u0_n158 ) );
  AOI21_X1 u0_u8_u0_U25 (.ZN( u0_u8_u0_n104 ) , .B1( u0_u8_u0_n107 ) , .B2( u0_u8_u0_n141 ) , .A( u0_u8_u0_n144 ) );
  AOI21_X1 u0_u8_u0_U26 (.B1( u0_u8_u0_n127 ) , .B2( u0_u8_u0_n129 ) , .A( u0_u8_u0_n138 ) , .ZN( u0_u8_u0_n96 ) );
  AOI21_X1 u0_u8_u0_U27 (.ZN( u0_u8_u0_n116 ) , .B2( u0_u8_u0_n142 ) , .A( u0_u8_u0_n144 ) , .B1( u0_u8_u0_n166 ) );
  NOR2_X1 u0_u8_u0_U28 (.A1( u0_u8_u0_n120 ) , .ZN( u0_u8_u0_n143 ) , .A2( u0_u8_u0_n167 ) );
  OAI221_X1 u0_u8_u0_U29 (.C1( u0_u8_u0_n112 ) , .ZN( u0_u8_u0_n120 ) , .B1( u0_u8_u0_n138 ) , .B2( u0_u8_u0_n141 ) , .C2( u0_u8_u0_n147 ) , .A( u0_u8_u0_n172 ) );
  INV_X1 u0_u8_u0_U3 (.A( u0_u8_u0_n113 ) , .ZN( u0_u8_u0_n166 ) );
  AOI211_X1 u0_u8_u0_U30 (.B( u0_u8_u0_n115 ) , .A( u0_u8_u0_n116 ) , .C2( u0_u8_u0_n117 ) , .C1( u0_u8_u0_n118 ) , .ZN( u0_u8_u0_n119 ) );
  NAND2_X1 u0_u8_u0_U31 (.A1( u0_u8_u0_n100 ) , .A2( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n125 ) );
  NAND2_X1 u0_u8_u0_U32 (.A2( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n140 ) , .A1( u0_u8_u0_n94 ) );
  NAND2_X1 u0_u8_u0_U33 (.A1( u0_u8_u0_n101 ) , .A2( u0_u8_u0_n102 ) , .ZN( u0_u8_u0_n150 ) );
  INV_X1 u0_u8_u0_U34 (.A( u0_u8_u0_n138 ) , .ZN( u0_u8_u0_n160 ) );
  NAND2_X1 u0_u8_u0_U35 (.A2( u0_u8_u0_n102 ) , .A1( u0_u8_u0_n103 ) , .ZN( u0_u8_u0_n149 ) );
  NAND2_X1 u0_u8_u0_U36 (.A2( u0_u8_u0_n100 ) , .A1( u0_u8_u0_n101 ) , .ZN( u0_u8_u0_n139 ) );
  NAND2_X1 u0_u8_u0_U37 (.A2( u0_u8_u0_n100 ) , .ZN( u0_u8_u0_n131 ) , .A1( u0_u8_u0_n92 ) );
  NAND2_X1 u0_u8_u0_U38 (.ZN( u0_u8_u0_n108 ) , .A1( u0_u8_u0_n92 ) , .A2( u0_u8_u0_n94 ) );
  NAND2_X1 u0_u8_u0_U39 (.A2( u0_u8_u0_n102 ) , .ZN( u0_u8_u0_n114 ) , .A1( u0_u8_u0_n92 ) );
  AOI21_X1 u0_u8_u0_U4 (.B1( u0_u8_u0_n114 ) , .ZN( u0_u8_u0_n115 ) , .B2( u0_u8_u0_n129 ) , .A( u0_u8_u0_n161 ) );
  NAND2_X1 u0_u8_u0_U40 (.A1( u0_u8_u0_n101 ) , .ZN( u0_u8_u0_n130 ) , .A2( u0_u8_u0_n94 ) );
  NAND2_X1 u0_u8_u0_U41 (.A2( u0_u8_u0_n101 ) , .ZN( u0_u8_u0_n121 ) , .A1( u0_u8_u0_n93 ) );
  INV_X1 u0_u8_u0_U42 (.ZN( u0_u8_u0_n172 ) , .A( u0_u8_u0_n88 ) );
  OAI222_X1 u0_u8_u0_U43 (.C1( u0_u8_u0_n108 ) , .A1( u0_u8_u0_n125 ) , .B2( u0_u8_u0_n128 ) , .B1( u0_u8_u0_n144 ) , .A2( u0_u8_u0_n158 ) , .C2( u0_u8_u0_n161 ) , .ZN( u0_u8_u0_n88 ) );
  NAND2_X1 u0_u8_u0_U44 (.ZN( u0_u8_u0_n112 ) , .A2( u0_u8_u0_n92 ) , .A1( u0_u8_u0_n93 ) );
  OR3_X1 u0_u8_u0_U45 (.A3( u0_u8_u0_n152 ) , .A2( u0_u8_u0_n153 ) , .A1( u0_u8_u0_n154 ) , .ZN( u0_u8_u0_n155 ) );
  AOI21_X1 u0_u8_u0_U46 (.A( u0_u8_u0_n144 ) , .B2( u0_u8_u0_n145 ) , .B1( u0_u8_u0_n146 ) , .ZN( u0_u8_u0_n154 ) );
  AOI21_X1 u0_u8_u0_U47 (.B2( u0_u8_u0_n150 ) , .B1( u0_u8_u0_n151 ) , .ZN( u0_u8_u0_n152 ) , .A( u0_u8_u0_n158 ) );
  AOI21_X1 u0_u8_u0_U48 (.A( u0_u8_u0_n147 ) , .B2( u0_u8_u0_n148 ) , .B1( u0_u8_u0_n149 ) , .ZN( u0_u8_u0_n153 ) );
  INV_X1 u0_u8_u0_U49 (.ZN( u0_u8_u0_n171 ) , .A( u0_u8_u0_n99 ) );
  AOI21_X1 u0_u8_u0_U5 (.B2( u0_u8_u0_n131 ) , .ZN( u0_u8_u0_n134 ) , .B1( u0_u8_u0_n151 ) , .A( u0_u8_u0_n158 ) );
  OAI211_X1 u0_u8_u0_U50 (.C2( u0_u8_u0_n140 ) , .C1( u0_u8_u0_n161 ) , .A( u0_u8_u0_n169 ) , .B( u0_u8_u0_n98 ) , .ZN( u0_u8_u0_n99 ) );
  INV_X1 u0_u8_u0_U51 (.ZN( u0_u8_u0_n169 ) , .A( u0_u8_u0_n91 ) );
  AOI211_X1 u0_u8_u0_U52 (.C1( u0_u8_u0_n118 ) , .A( u0_u8_u0_n123 ) , .B( u0_u8_u0_n96 ) , .C2( u0_u8_u0_n97 ) , .ZN( u0_u8_u0_n98 ) );
  NOR2_X1 u0_u8_u0_U53 (.A2( u0_u8_X_2 ) , .ZN( u0_u8_u0_n103 ) , .A1( u0_u8_u0_n164 ) );
  NOR2_X1 u0_u8_u0_U54 (.A2( u0_u8_X_4 ) , .A1( u0_u8_X_5 ) , .ZN( u0_u8_u0_n118 ) );
  NOR2_X1 u0_u8_u0_U55 (.A2( u0_u8_X_1 ) , .A1( u0_u8_X_2 ) , .ZN( u0_u8_u0_n92 ) );
  NOR2_X1 u0_u8_u0_U56 (.A2( u0_u8_X_1 ) , .ZN( u0_u8_u0_n101 ) , .A1( u0_u8_u0_n163 ) );
  NOR2_X1 u0_u8_u0_U57 (.A2( u0_u8_X_3 ) , .A1( u0_u8_X_6 ) , .ZN( u0_u8_u0_n94 ) );
  NOR2_X1 u0_u8_u0_U58 (.A2( u0_u8_X_6 ) , .ZN( u0_u8_u0_n100 ) , .A1( u0_u8_u0_n162 ) );
  NAND2_X1 u0_u8_u0_U59 (.A2( u0_u8_X_4 ) , .A1( u0_u8_X_5 ) , .ZN( u0_u8_u0_n144 ) );
  NOR2_X1 u0_u8_u0_U6 (.A1( u0_u8_u0_n108 ) , .ZN( u0_u8_u0_n123 ) , .A2( u0_u8_u0_n158 ) );
  NOR2_X1 u0_u8_u0_U60 (.A2( u0_u8_X_5 ) , .ZN( u0_u8_u0_n136 ) , .A1( u0_u8_u0_n159 ) );
  NAND2_X1 u0_u8_u0_U61 (.A1( u0_u8_X_5 ) , .ZN( u0_u8_u0_n138 ) , .A2( u0_u8_u0_n159 ) );
  AND2_X1 u0_u8_u0_U62 (.A2( u0_u8_X_3 ) , .A1( u0_u8_X_6 ) , .ZN( u0_u8_u0_n102 ) );
  AND2_X1 u0_u8_u0_U63 (.A1( u0_u8_X_6 ) , .A2( u0_u8_u0_n162 ) , .ZN( u0_u8_u0_n93 ) );
  INV_X1 u0_u8_u0_U64 (.A( u0_u8_X_4 ) , .ZN( u0_u8_u0_n159 ) );
  INV_X1 u0_u8_u0_U65 (.A( u0_u8_X_2 ) , .ZN( u0_u8_u0_n163 ) );
  INV_X1 u0_u8_u0_U66 (.A( u0_u8_X_3 ) , .ZN( u0_u8_u0_n162 ) );
  INV_X1 u0_u8_u0_U67 (.A( u0_u8_u0_n126 ) , .ZN( u0_u8_u0_n168 ) );
  AOI211_X1 u0_u8_u0_U68 (.B( u0_u8_u0_n133 ) , .A( u0_u8_u0_n134 ) , .C2( u0_u8_u0_n135 ) , .C1( u0_u8_u0_n136 ) , .ZN( u0_u8_u0_n137 ) );
  OR4_X1 u0_u8_u0_U69 (.ZN( u0_out8_17 ) , .A4( u0_u8_u0_n122 ) , .A2( u0_u8_u0_n123 ) , .A1( u0_u8_u0_n124 ) , .A3( u0_u8_u0_n170 ) );
  OAI21_X1 u0_u8_u0_U7 (.B1( u0_u8_u0_n150 ) , .B2( u0_u8_u0_n158 ) , .A( u0_u8_u0_n172 ) , .ZN( u0_u8_u0_n89 ) );
  AOI21_X1 u0_u8_u0_U70 (.B2( u0_u8_u0_n107 ) , .ZN( u0_u8_u0_n124 ) , .B1( u0_u8_u0_n128 ) , .A( u0_u8_u0_n161 ) );
  INV_X1 u0_u8_u0_U71 (.A( u0_u8_u0_n111 ) , .ZN( u0_u8_u0_n170 ) );
  OR4_X1 u0_u8_u0_U72 (.ZN( u0_out8_31 ) , .A4( u0_u8_u0_n155 ) , .A2( u0_u8_u0_n156 ) , .A1( u0_u8_u0_n157 ) , .A3( u0_u8_u0_n173 ) );
  AOI21_X1 u0_u8_u0_U73 (.A( u0_u8_u0_n138 ) , .B2( u0_u8_u0_n139 ) , .B1( u0_u8_u0_n140 ) , .ZN( u0_u8_u0_n157 ) );
  AOI21_X1 u0_u8_u0_U74 (.B2( u0_u8_u0_n141 ) , .B1( u0_u8_u0_n142 ) , .ZN( u0_u8_u0_n156 ) , .A( u0_u8_u0_n161 ) );
  INV_X1 u0_u8_u0_U75 (.ZN( u0_u8_u0_n174 ) , .A( u0_u8_u0_n89 ) );
  AOI211_X1 u0_u8_u0_U76 (.B( u0_u8_u0_n104 ) , .A( u0_u8_u0_n105 ) , .ZN( u0_u8_u0_n106 ) , .C2( u0_u8_u0_n113 ) , .C1( u0_u8_u0_n160 ) );
  INV_X1 u0_u8_u0_U77 (.A( u0_u8_X_1 ) , .ZN( u0_u8_u0_n164 ) );
  NOR2_X1 u0_u8_u0_U78 (.A1( u0_u8_u0_n163 ) , .A2( u0_u8_u0_n164 ) , .ZN( u0_u8_u0_n95 ) );
  OAI221_X1 u0_u8_u0_U79 (.C1( u0_u8_u0_n121 ) , .ZN( u0_u8_u0_n122 ) , .B2( u0_u8_u0_n127 ) , .A( u0_u8_u0_n143 ) , .B1( u0_u8_u0_n144 ) , .C2( u0_u8_u0_n147 ) );
  AND2_X1 u0_u8_u0_U8 (.A1( u0_u8_u0_n114 ) , .A2( u0_u8_u0_n121 ) , .ZN( u0_u8_u0_n146 ) );
  AOI21_X1 u0_u8_u0_U80 (.B1( u0_u8_u0_n132 ) , .ZN( u0_u8_u0_n133 ) , .A( u0_u8_u0_n144 ) , .B2( u0_u8_u0_n166 ) );
  OAI22_X1 u0_u8_u0_U81 (.ZN( u0_u8_u0_n105 ) , .A2( u0_u8_u0_n132 ) , .B1( u0_u8_u0_n146 ) , .A1( u0_u8_u0_n147 ) , .B2( u0_u8_u0_n161 ) );
  NAND2_X1 u0_u8_u0_U82 (.ZN( u0_u8_u0_n110 ) , .A2( u0_u8_u0_n132 ) , .A1( u0_u8_u0_n145 ) );
  INV_X1 u0_u8_u0_U83 (.A( u0_u8_u0_n119 ) , .ZN( u0_u8_u0_n167 ) );
  NAND2_X1 u0_u8_u0_U84 (.ZN( u0_u8_u0_n148 ) , .A1( u0_u8_u0_n93 ) , .A2( u0_u8_u0_n95 ) );
  NAND2_X1 u0_u8_u0_U85 (.A1( u0_u8_u0_n100 ) , .ZN( u0_u8_u0_n129 ) , .A2( u0_u8_u0_n95 ) );
  NAND2_X1 u0_u8_u0_U86 (.A1( u0_u8_u0_n102 ) , .ZN( u0_u8_u0_n128 ) , .A2( u0_u8_u0_n95 ) );
  NAND2_X1 u0_u8_u0_U87 (.ZN( u0_u8_u0_n142 ) , .A1( u0_u8_u0_n94 ) , .A2( u0_u8_u0_n95 ) );
  NAND3_X1 u0_u8_u0_U88 (.ZN( u0_out8_23 ) , .A3( u0_u8_u0_n137 ) , .A1( u0_u8_u0_n168 ) , .A2( u0_u8_u0_n171 ) );
  NAND3_X1 u0_u8_u0_U89 (.A3( u0_u8_u0_n127 ) , .A2( u0_u8_u0_n128 ) , .ZN( u0_u8_u0_n135 ) , .A1( u0_u8_u0_n150 ) );
  AND2_X1 u0_u8_u0_U9 (.A1( u0_u8_u0_n131 ) , .ZN( u0_u8_u0_n141 ) , .A2( u0_u8_u0_n150 ) );
  NAND3_X1 u0_u8_u0_U90 (.ZN( u0_u8_u0_n117 ) , .A3( u0_u8_u0_n132 ) , .A2( u0_u8_u0_n139 ) , .A1( u0_u8_u0_n148 ) );
  NAND3_X1 u0_u8_u0_U91 (.ZN( u0_u8_u0_n109 ) , .A2( u0_u8_u0_n114 ) , .A3( u0_u8_u0_n140 ) , .A1( u0_u8_u0_n149 ) );
  NAND3_X1 u0_u8_u0_U92 (.ZN( u0_out8_9 ) , .A3( u0_u8_u0_n106 ) , .A2( u0_u8_u0_n171 ) , .A1( u0_u8_u0_n174 ) );
  NAND3_X1 u0_u8_u0_U93 (.A2( u0_u8_u0_n128 ) , .A1( u0_u8_u0_n132 ) , .A3( u0_u8_u0_n146 ) , .ZN( u0_u8_u0_n97 ) );
  AOI21_X1 u0_u8_u1_U10 (.B2( u0_u8_u1_n155 ) , .B1( u0_u8_u1_n156 ) , .ZN( u0_u8_u1_n157 ) , .A( u0_u8_u1_n174 ) );
  NAND3_X1 u0_u8_u1_U100 (.ZN( u0_u8_u1_n113 ) , .A1( u0_u8_u1_n120 ) , .A3( u0_u8_u1_n133 ) , .A2( u0_u8_u1_n155 ) );
  NAND2_X1 u0_u8_u1_U11 (.ZN( u0_u8_u1_n140 ) , .A2( u0_u8_u1_n150 ) , .A1( u0_u8_u1_n155 ) );
  NAND2_X1 u0_u8_u1_U12 (.A1( u0_u8_u1_n131 ) , .ZN( u0_u8_u1_n147 ) , .A2( u0_u8_u1_n153 ) );
  AOI22_X1 u0_u8_u1_U13 (.B2( u0_u8_u1_n136 ) , .A2( u0_u8_u1_n137 ) , .ZN( u0_u8_u1_n143 ) , .A1( u0_u8_u1_n171 ) , .B1( u0_u8_u1_n173 ) );
  INV_X1 u0_u8_u1_U14 (.A( u0_u8_u1_n147 ) , .ZN( u0_u8_u1_n181 ) );
  INV_X1 u0_u8_u1_U15 (.A( u0_u8_u1_n139 ) , .ZN( u0_u8_u1_n174 ) );
  OR4_X1 u0_u8_u1_U16 (.A4( u0_u8_u1_n106 ) , .A3( u0_u8_u1_n107 ) , .ZN( u0_u8_u1_n108 ) , .A1( u0_u8_u1_n117 ) , .A2( u0_u8_u1_n184 ) );
  AOI21_X1 u0_u8_u1_U17 (.ZN( u0_u8_u1_n106 ) , .A( u0_u8_u1_n112 ) , .B1( u0_u8_u1_n154 ) , .B2( u0_u8_u1_n156 ) );
  AOI21_X1 u0_u8_u1_U18 (.ZN( u0_u8_u1_n107 ) , .B1( u0_u8_u1_n134 ) , .B2( u0_u8_u1_n149 ) , .A( u0_u8_u1_n174 ) );
  INV_X1 u0_u8_u1_U19 (.A( u0_u8_u1_n101 ) , .ZN( u0_u8_u1_n184 ) );
  INV_X1 u0_u8_u1_U20 (.A( u0_u8_u1_n112 ) , .ZN( u0_u8_u1_n171 ) );
  NAND2_X1 u0_u8_u1_U21 (.ZN( u0_u8_u1_n141 ) , .A1( u0_u8_u1_n153 ) , .A2( u0_u8_u1_n156 ) );
  AND2_X1 u0_u8_u1_U22 (.A1( u0_u8_u1_n123 ) , .ZN( u0_u8_u1_n134 ) , .A2( u0_u8_u1_n161 ) );
  NAND2_X1 u0_u8_u1_U23 (.A2( u0_u8_u1_n115 ) , .A1( u0_u8_u1_n116 ) , .ZN( u0_u8_u1_n148 ) );
  NAND2_X1 u0_u8_u1_U24 (.A2( u0_u8_u1_n133 ) , .A1( u0_u8_u1_n135 ) , .ZN( u0_u8_u1_n159 ) );
  NAND2_X1 u0_u8_u1_U25 (.A2( u0_u8_u1_n115 ) , .A1( u0_u8_u1_n120 ) , .ZN( u0_u8_u1_n132 ) );
  INV_X1 u0_u8_u1_U26 (.A( u0_u8_u1_n154 ) , .ZN( u0_u8_u1_n178 ) );
  INV_X1 u0_u8_u1_U27 (.A( u0_u8_u1_n151 ) , .ZN( u0_u8_u1_n183 ) );
  AND2_X1 u0_u8_u1_U28 (.A1( u0_u8_u1_n129 ) , .A2( u0_u8_u1_n133 ) , .ZN( u0_u8_u1_n149 ) );
  INV_X1 u0_u8_u1_U29 (.A( u0_u8_u1_n131 ) , .ZN( u0_u8_u1_n180 ) );
  INV_X1 u0_u8_u1_U3 (.A( u0_u8_u1_n159 ) , .ZN( u0_u8_u1_n182 ) );
  AOI221_X1 u0_u8_u1_U30 (.B1( u0_u8_u1_n140 ) , .ZN( u0_u8_u1_n167 ) , .B2( u0_u8_u1_n172 ) , .C2( u0_u8_u1_n175 ) , .C1( u0_u8_u1_n178 ) , .A( u0_u8_u1_n188 ) );
  INV_X1 u0_u8_u1_U31 (.ZN( u0_u8_u1_n188 ) , .A( u0_u8_u1_n97 ) );
  AOI211_X1 u0_u8_u1_U32 (.A( u0_u8_u1_n118 ) , .C1( u0_u8_u1_n132 ) , .C2( u0_u8_u1_n139 ) , .B( u0_u8_u1_n96 ) , .ZN( u0_u8_u1_n97 ) );
  AOI21_X1 u0_u8_u1_U33 (.B2( u0_u8_u1_n121 ) , .B1( u0_u8_u1_n135 ) , .A( u0_u8_u1_n152 ) , .ZN( u0_u8_u1_n96 ) );
  OAI221_X1 u0_u8_u1_U34 (.A( u0_u8_u1_n119 ) , .C2( u0_u8_u1_n129 ) , .ZN( u0_u8_u1_n138 ) , .B2( u0_u8_u1_n152 ) , .C1( u0_u8_u1_n174 ) , .B1( u0_u8_u1_n187 ) );
  INV_X1 u0_u8_u1_U35 (.A( u0_u8_u1_n148 ) , .ZN( u0_u8_u1_n187 ) );
  AOI211_X1 u0_u8_u1_U36 (.B( u0_u8_u1_n117 ) , .A( u0_u8_u1_n118 ) , .ZN( u0_u8_u1_n119 ) , .C2( u0_u8_u1_n146 ) , .C1( u0_u8_u1_n159 ) );
  NOR2_X1 u0_u8_u1_U37 (.A1( u0_u8_u1_n168 ) , .A2( u0_u8_u1_n176 ) , .ZN( u0_u8_u1_n98 ) );
  AOI211_X1 u0_u8_u1_U38 (.B( u0_u8_u1_n162 ) , .A( u0_u8_u1_n163 ) , .C2( u0_u8_u1_n164 ) , .ZN( u0_u8_u1_n165 ) , .C1( u0_u8_u1_n171 ) );
  AOI21_X1 u0_u8_u1_U39 (.A( u0_u8_u1_n160 ) , .B2( u0_u8_u1_n161 ) , .ZN( u0_u8_u1_n162 ) , .B1( u0_u8_u1_n182 ) );
  AOI221_X1 u0_u8_u1_U4 (.A( u0_u8_u1_n138 ) , .C2( u0_u8_u1_n139 ) , .C1( u0_u8_u1_n140 ) , .B2( u0_u8_u1_n141 ) , .ZN( u0_u8_u1_n142 ) , .B1( u0_u8_u1_n175 ) );
  OR2_X1 u0_u8_u1_U40 (.A2( u0_u8_u1_n157 ) , .A1( u0_u8_u1_n158 ) , .ZN( u0_u8_u1_n163 ) );
  NAND2_X1 u0_u8_u1_U41 (.A1( u0_u8_u1_n128 ) , .ZN( u0_u8_u1_n146 ) , .A2( u0_u8_u1_n160 ) );
  NAND2_X1 u0_u8_u1_U42 (.A2( u0_u8_u1_n112 ) , .ZN( u0_u8_u1_n139 ) , .A1( u0_u8_u1_n152 ) );
  NAND2_X1 u0_u8_u1_U43 (.A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n156 ) , .A2( u0_u8_u1_n99 ) );
  NOR2_X1 u0_u8_u1_U44 (.ZN( u0_u8_u1_n117 ) , .A1( u0_u8_u1_n121 ) , .A2( u0_u8_u1_n160 ) );
  OAI21_X1 u0_u8_u1_U45 (.B2( u0_u8_u1_n123 ) , .ZN( u0_u8_u1_n145 ) , .B1( u0_u8_u1_n160 ) , .A( u0_u8_u1_n185 ) );
  INV_X1 u0_u8_u1_U46 (.A( u0_u8_u1_n122 ) , .ZN( u0_u8_u1_n185 ) );
  AOI21_X1 u0_u8_u1_U47 (.B2( u0_u8_u1_n120 ) , .B1( u0_u8_u1_n121 ) , .ZN( u0_u8_u1_n122 ) , .A( u0_u8_u1_n128 ) );
  AOI21_X1 u0_u8_u1_U48 (.A( u0_u8_u1_n128 ) , .B2( u0_u8_u1_n129 ) , .ZN( u0_u8_u1_n130 ) , .B1( u0_u8_u1_n150 ) );
  NAND2_X1 u0_u8_u1_U49 (.ZN( u0_u8_u1_n112 ) , .A1( u0_u8_u1_n169 ) , .A2( u0_u8_u1_n170 ) );
  AOI211_X1 u0_u8_u1_U5 (.ZN( u0_u8_u1_n124 ) , .A( u0_u8_u1_n138 ) , .C2( u0_u8_u1_n139 ) , .B( u0_u8_u1_n145 ) , .C1( u0_u8_u1_n147 ) );
  NAND2_X1 u0_u8_u1_U50 (.ZN( u0_u8_u1_n129 ) , .A2( u0_u8_u1_n95 ) , .A1( u0_u8_u1_n98 ) );
  NAND2_X1 u0_u8_u1_U51 (.A1( u0_u8_u1_n102 ) , .ZN( u0_u8_u1_n154 ) , .A2( u0_u8_u1_n99 ) );
  NAND2_X1 u0_u8_u1_U52 (.A2( u0_u8_u1_n100 ) , .ZN( u0_u8_u1_n135 ) , .A1( u0_u8_u1_n99 ) );
  AOI21_X1 u0_u8_u1_U53 (.A( u0_u8_u1_n152 ) , .B2( u0_u8_u1_n153 ) , .B1( u0_u8_u1_n154 ) , .ZN( u0_u8_u1_n158 ) );
  INV_X1 u0_u8_u1_U54 (.A( u0_u8_u1_n160 ) , .ZN( u0_u8_u1_n175 ) );
  NAND2_X1 u0_u8_u1_U55 (.A1( u0_u8_u1_n100 ) , .ZN( u0_u8_u1_n116 ) , .A2( u0_u8_u1_n95 ) );
  NAND2_X1 u0_u8_u1_U56 (.A1( u0_u8_u1_n102 ) , .ZN( u0_u8_u1_n131 ) , .A2( u0_u8_u1_n95 ) );
  NAND2_X1 u0_u8_u1_U57 (.A2( u0_u8_u1_n104 ) , .ZN( u0_u8_u1_n121 ) , .A1( u0_u8_u1_n98 ) );
  NAND2_X1 u0_u8_u1_U58 (.A1( u0_u8_u1_n103 ) , .ZN( u0_u8_u1_n153 ) , .A2( u0_u8_u1_n98 ) );
  NAND2_X1 u0_u8_u1_U59 (.A2( u0_u8_u1_n104 ) , .A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n133 ) );
  AOI22_X1 u0_u8_u1_U6 (.B2( u0_u8_u1_n113 ) , .A2( u0_u8_u1_n114 ) , .ZN( u0_u8_u1_n125 ) , .A1( u0_u8_u1_n171 ) , .B1( u0_u8_u1_n173 ) );
  NAND2_X1 u0_u8_u1_U60 (.ZN( u0_u8_u1_n150 ) , .A2( u0_u8_u1_n98 ) , .A1( u0_u8_u1_n99 ) );
  NAND2_X1 u0_u8_u1_U61 (.A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n155 ) , .A2( u0_u8_u1_n95 ) );
  OAI21_X1 u0_u8_u1_U62 (.ZN( u0_u8_u1_n109 ) , .B1( u0_u8_u1_n129 ) , .B2( u0_u8_u1_n160 ) , .A( u0_u8_u1_n167 ) );
  NAND2_X1 u0_u8_u1_U63 (.A2( u0_u8_u1_n100 ) , .A1( u0_u8_u1_n103 ) , .ZN( u0_u8_u1_n120 ) );
  NAND2_X1 u0_u8_u1_U64 (.A1( u0_u8_u1_n102 ) , .A2( u0_u8_u1_n104 ) , .ZN( u0_u8_u1_n115 ) );
  NAND2_X1 u0_u8_u1_U65 (.A2( u0_u8_u1_n100 ) , .A1( u0_u8_u1_n104 ) , .ZN( u0_u8_u1_n151 ) );
  NAND2_X1 u0_u8_u1_U66 (.A2( u0_u8_u1_n103 ) , .A1( u0_u8_u1_n105 ) , .ZN( u0_u8_u1_n161 ) );
  INV_X1 u0_u8_u1_U67 (.A( u0_u8_u1_n152 ) , .ZN( u0_u8_u1_n173 ) );
  INV_X1 u0_u8_u1_U68 (.A( u0_u8_u1_n128 ) , .ZN( u0_u8_u1_n172 ) );
  NAND2_X1 u0_u8_u1_U69 (.A2( u0_u8_u1_n102 ) , .A1( u0_u8_u1_n103 ) , .ZN( u0_u8_u1_n123 ) );
  NAND2_X1 u0_u8_u1_U7 (.ZN( u0_u8_u1_n114 ) , .A1( u0_u8_u1_n134 ) , .A2( u0_u8_u1_n156 ) );
  NOR2_X1 u0_u8_u1_U70 (.A2( u0_u8_X_7 ) , .A1( u0_u8_X_8 ) , .ZN( u0_u8_u1_n95 ) );
  NOR2_X1 u0_u8_u1_U71 (.A1( u0_u8_X_12 ) , .A2( u0_u8_X_9 ) , .ZN( u0_u8_u1_n100 ) );
  NOR2_X1 u0_u8_u1_U72 (.A2( u0_u8_X_8 ) , .A1( u0_u8_u1_n177 ) , .ZN( u0_u8_u1_n99 ) );
  NOR2_X1 u0_u8_u1_U73 (.A2( u0_u8_X_12 ) , .ZN( u0_u8_u1_n102 ) , .A1( u0_u8_u1_n176 ) );
  NOR2_X1 u0_u8_u1_U74 (.A2( u0_u8_X_9 ) , .ZN( u0_u8_u1_n105 ) , .A1( u0_u8_u1_n168 ) );
  NAND2_X1 u0_u8_u1_U75 (.A1( u0_u8_X_10 ) , .ZN( u0_u8_u1_n160 ) , .A2( u0_u8_u1_n169 ) );
  NAND2_X1 u0_u8_u1_U76 (.A2( u0_u8_X_10 ) , .A1( u0_u8_X_11 ) , .ZN( u0_u8_u1_n152 ) );
  NAND2_X1 u0_u8_u1_U77 (.A1( u0_u8_X_11 ) , .ZN( u0_u8_u1_n128 ) , .A2( u0_u8_u1_n170 ) );
  AND2_X1 u0_u8_u1_U78 (.A2( u0_u8_X_7 ) , .A1( u0_u8_X_8 ) , .ZN( u0_u8_u1_n104 ) );
  AND2_X1 u0_u8_u1_U79 (.A1( u0_u8_X_8 ) , .ZN( u0_u8_u1_n103 ) , .A2( u0_u8_u1_n177 ) );
  NOR2_X1 u0_u8_u1_U8 (.A1( u0_u8_u1_n112 ) , .A2( u0_u8_u1_n116 ) , .ZN( u0_u8_u1_n118 ) );
  INV_X1 u0_u8_u1_U80 (.A( u0_u8_X_10 ) , .ZN( u0_u8_u1_n170 ) );
  INV_X1 u0_u8_u1_U81 (.A( u0_u8_X_9 ) , .ZN( u0_u8_u1_n176 ) );
  INV_X1 u0_u8_u1_U82 (.A( u0_u8_X_11 ) , .ZN( u0_u8_u1_n169 ) );
  INV_X1 u0_u8_u1_U83 (.A( u0_u8_X_12 ) , .ZN( u0_u8_u1_n168 ) );
  INV_X1 u0_u8_u1_U84 (.A( u0_u8_X_7 ) , .ZN( u0_u8_u1_n177 ) );
  NAND4_X1 u0_u8_u1_U85 (.ZN( u0_out8_28 ) , .A4( u0_u8_u1_n124 ) , .A3( u0_u8_u1_n125 ) , .A2( u0_u8_u1_n126 ) , .A1( u0_u8_u1_n127 ) );
  OAI21_X1 u0_u8_u1_U86 (.ZN( u0_u8_u1_n127 ) , .B2( u0_u8_u1_n139 ) , .B1( u0_u8_u1_n175 ) , .A( u0_u8_u1_n183 ) );
  OAI21_X1 u0_u8_u1_U87 (.ZN( u0_u8_u1_n126 ) , .B2( u0_u8_u1_n140 ) , .A( u0_u8_u1_n146 ) , .B1( u0_u8_u1_n178 ) );
  NAND4_X1 u0_u8_u1_U88 (.ZN( u0_out8_18 ) , .A4( u0_u8_u1_n165 ) , .A3( u0_u8_u1_n166 ) , .A1( u0_u8_u1_n167 ) , .A2( u0_u8_u1_n186 ) );
  AOI22_X1 u0_u8_u1_U89 (.B2( u0_u8_u1_n146 ) , .B1( u0_u8_u1_n147 ) , .A2( u0_u8_u1_n148 ) , .ZN( u0_u8_u1_n166 ) , .A1( u0_u8_u1_n172 ) );
  OAI21_X1 u0_u8_u1_U9 (.ZN( u0_u8_u1_n101 ) , .B1( u0_u8_u1_n141 ) , .A( u0_u8_u1_n146 ) , .B2( u0_u8_u1_n183 ) );
  INV_X1 u0_u8_u1_U90 (.A( u0_u8_u1_n145 ) , .ZN( u0_u8_u1_n186 ) );
  NAND4_X1 u0_u8_u1_U91 (.ZN( u0_out8_2 ) , .A4( u0_u8_u1_n142 ) , .A3( u0_u8_u1_n143 ) , .A2( u0_u8_u1_n144 ) , .A1( u0_u8_u1_n179 ) );
  OAI21_X1 u0_u8_u1_U92 (.B2( u0_u8_u1_n132 ) , .ZN( u0_u8_u1_n144 ) , .A( u0_u8_u1_n146 ) , .B1( u0_u8_u1_n180 ) );
  INV_X1 u0_u8_u1_U93 (.A( u0_u8_u1_n130 ) , .ZN( u0_u8_u1_n179 ) );
  OR4_X1 u0_u8_u1_U94 (.ZN( u0_out8_13 ) , .A4( u0_u8_u1_n108 ) , .A3( u0_u8_u1_n109 ) , .A2( u0_u8_u1_n110 ) , .A1( u0_u8_u1_n111 ) );
  AOI21_X1 u0_u8_u1_U95 (.ZN( u0_u8_u1_n111 ) , .A( u0_u8_u1_n128 ) , .B2( u0_u8_u1_n131 ) , .B1( u0_u8_u1_n135 ) );
  AOI21_X1 u0_u8_u1_U96 (.ZN( u0_u8_u1_n110 ) , .A( u0_u8_u1_n116 ) , .B1( u0_u8_u1_n152 ) , .B2( u0_u8_u1_n160 ) );
  NAND3_X1 u0_u8_u1_U97 (.A3( u0_u8_u1_n149 ) , .A2( u0_u8_u1_n150 ) , .A1( u0_u8_u1_n151 ) , .ZN( u0_u8_u1_n164 ) );
  NAND3_X1 u0_u8_u1_U98 (.A3( u0_u8_u1_n134 ) , .A2( u0_u8_u1_n135 ) , .ZN( u0_u8_u1_n136 ) , .A1( u0_u8_u1_n151 ) );
  NAND3_X1 u0_u8_u1_U99 (.A1( u0_u8_u1_n133 ) , .ZN( u0_u8_u1_n137 ) , .A2( u0_u8_u1_n154 ) , .A3( u0_u8_u1_n181 ) );
  OAI22_X1 u0_u8_u2_U10 (.B1( u0_u8_u2_n151 ) , .A2( u0_u8_u2_n152 ) , .A1( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n160 ) , .B2( u0_u8_u2_n168 ) );
  NAND3_X1 u0_u8_u2_U100 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n104 ) , .A3( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n98 ) );
  NOR3_X1 u0_u8_u2_U11 (.A1( u0_u8_u2_n150 ) , .ZN( u0_u8_u2_n151 ) , .A3( u0_u8_u2_n175 ) , .A2( u0_u8_u2_n188 ) );
  AOI21_X1 u0_u8_u2_U12 (.B2( u0_u8_u2_n123 ) , .ZN( u0_u8_u2_n125 ) , .A( u0_u8_u2_n171 ) , .B1( u0_u8_u2_n184 ) );
  INV_X1 u0_u8_u2_U13 (.A( u0_u8_u2_n150 ) , .ZN( u0_u8_u2_n184 ) );
  AOI21_X1 u0_u8_u2_U14 (.ZN( u0_u8_u2_n144 ) , .B2( u0_u8_u2_n155 ) , .A( u0_u8_u2_n172 ) , .B1( u0_u8_u2_n185 ) );
  AOI21_X1 u0_u8_u2_U15 (.B2( u0_u8_u2_n143 ) , .ZN( u0_u8_u2_n145 ) , .B1( u0_u8_u2_n152 ) , .A( u0_u8_u2_n171 ) );
  INV_X1 u0_u8_u2_U16 (.A( u0_u8_u2_n156 ) , .ZN( u0_u8_u2_n171 ) );
  INV_X1 u0_u8_u2_U17 (.A( u0_u8_u2_n120 ) , .ZN( u0_u8_u2_n188 ) );
  NAND2_X1 u0_u8_u2_U18 (.A2( u0_u8_u2_n122 ) , .ZN( u0_u8_u2_n150 ) , .A1( u0_u8_u2_n152 ) );
  INV_X1 u0_u8_u2_U19 (.A( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n170 ) );
  INV_X1 u0_u8_u2_U20 (.A( u0_u8_u2_n137 ) , .ZN( u0_u8_u2_n173 ) );
  NAND2_X1 u0_u8_u2_U21 (.A1( u0_u8_u2_n132 ) , .A2( u0_u8_u2_n139 ) , .ZN( u0_u8_u2_n157 ) );
  INV_X1 u0_u8_u2_U22 (.A( u0_u8_u2_n113 ) , .ZN( u0_u8_u2_n178 ) );
  INV_X1 u0_u8_u2_U23 (.A( u0_u8_u2_n139 ) , .ZN( u0_u8_u2_n175 ) );
  INV_X1 u0_u8_u2_U24 (.A( u0_u8_u2_n155 ) , .ZN( u0_u8_u2_n181 ) );
  INV_X1 u0_u8_u2_U25 (.A( u0_u8_u2_n119 ) , .ZN( u0_u8_u2_n177 ) );
  INV_X1 u0_u8_u2_U26 (.A( u0_u8_u2_n116 ) , .ZN( u0_u8_u2_n180 ) );
  INV_X1 u0_u8_u2_U27 (.A( u0_u8_u2_n131 ) , .ZN( u0_u8_u2_n179 ) );
  INV_X1 u0_u8_u2_U28 (.A( u0_u8_u2_n154 ) , .ZN( u0_u8_u2_n176 ) );
  NAND2_X1 u0_u8_u2_U29 (.A2( u0_u8_u2_n116 ) , .A1( u0_u8_u2_n117 ) , .ZN( u0_u8_u2_n118 ) );
  NOR2_X1 u0_u8_u2_U3 (.ZN( u0_u8_u2_n121 ) , .A2( u0_u8_u2_n177 ) , .A1( u0_u8_u2_n180 ) );
  INV_X1 u0_u8_u2_U30 (.A( u0_u8_u2_n132 ) , .ZN( u0_u8_u2_n182 ) );
  INV_X1 u0_u8_u2_U31 (.A( u0_u8_u2_n158 ) , .ZN( u0_u8_u2_n183 ) );
  OAI21_X1 u0_u8_u2_U32 (.A( u0_u8_u2_n156 ) , .B1( u0_u8_u2_n157 ) , .ZN( u0_u8_u2_n158 ) , .B2( u0_u8_u2_n179 ) );
  NOR2_X1 u0_u8_u2_U33 (.ZN( u0_u8_u2_n156 ) , .A1( u0_u8_u2_n166 ) , .A2( u0_u8_u2_n169 ) );
  NOR2_X1 u0_u8_u2_U34 (.A2( u0_u8_u2_n114 ) , .ZN( u0_u8_u2_n137 ) , .A1( u0_u8_u2_n140 ) );
  NOR2_X1 u0_u8_u2_U35 (.A2( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n153 ) , .A1( u0_u8_u2_n156 ) );
  AOI211_X1 u0_u8_u2_U36 (.ZN( u0_u8_u2_n130 ) , .C1( u0_u8_u2_n138 ) , .C2( u0_u8_u2_n179 ) , .B( u0_u8_u2_n96 ) , .A( u0_u8_u2_n97 ) );
  OAI22_X1 u0_u8_u2_U37 (.B1( u0_u8_u2_n133 ) , .A2( u0_u8_u2_n137 ) , .A1( u0_u8_u2_n152 ) , .B2( u0_u8_u2_n168 ) , .ZN( u0_u8_u2_n97 ) );
  OAI221_X1 u0_u8_u2_U38 (.B1( u0_u8_u2_n113 ) , .C1( u0_u8_u2_n132 ) , .A( u0_u8_u2_n149 ) , .B2( u0_u8_u2_n171 ) , .C2( u0_u8_u2_n172 ) , .ZN( u0_u8_u2_n96 ) );
  OAI221_X1 u0_u8_u2_U39 (.A( u0_u8_u2_n115 ) , .C2( u0_u8_u2_n123 ) , .B2( u0_u8_u2_n143 ) , .B1( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n163 ) , .C1( u0_u8_u2_n168 ) );
  INV_X1 u0_u8_u2_U4 (.A( u0_u8_u2_n134 ) , .ZN( u0_u8_u2_n185 ) );
  OAI21_X1 u0_u8_u2_U40 (.A( u0_u8_u2_n114 ) , .ZN( u0_u8_u2_n115 ) , .B1( u0_u8_u2_n176 ) , .B2( u0_u8_u2_n178 ) );
  OAI221_X1 u0_u8_u2_U41 (.A( u0_u8_u2_n135 ) , .B2( u0_u8_u2_n136 ) , .B1( u0_u8_u2_n137 ) , .ZN( u0_u8_u2_n162 ) , .C2( u0_u8_u2_n167 ) , .C1( u0_u8_u2_n185 ) );
  AND3_X1 u0_u8_u2_U42 (.A3( u0_u8_u2_n131 ) , .A2( u0_u8_u2_n132 ) , .A1( u0_u8_u2_n133 ) , .ZN( u0_u8_u2_n136 ) );
  AOI22_X1 u0_u8_u2_U43 (.ZN( u0_u8_u2_n135 ) , .B1( u0_u8_u2_n140 ) , .A1( u0_u8_u2_n156 ) , .B2( u0_u8_u2_n180 ) , .A2( u0_u8_u2_n188 ) );
  AOI21_X1 u0_u8_u2_U44 (.ZN( u0_u8_u2_n149 ) , .B1( u0_u8_u2_n173 ) , .B2( u0_u8_u2_n188 ) , .A( u0_u8_u2_n95 ) );
  AND3_X1 u0_u8_u2_U45 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n104 ) , .A3( u0_u8_u2_n156 ) , .ZN( u0_u8_u2_n95 ) );
  OAI21_X1 u0_u8_u2_U46 (.A( u0_u8_u2_n141 ) , .B2( u0_u8_u2_n142 ) , .ZN( u0_u8_u2_n146 ) , .B1( u0_u8_u2_n153 ) );
  OAI21_X1 u0_u8_u2_U47 (.A( u0_u8_u2_n140 ) , .ZN( u0_u8_u2_n141 ) , .B1( u0_u8_u2_n176 ) , .B2( u0_u8_u2_n177 ) );
  NOR3_X1 u0_u8_u2_U48 (.ZN( u0_u8_u2_n142 ) , .A3( u0_u8_u2_n175 ) , .A2( u0_u8_u2_n178 ) , .A1( u0_u8_u2_n181 ) );
  OAI21_X1 u0_u8_u2_U49 (.A( u0_u8_u2_n101 ) , .B2( u0_u8_u2_n121 ) , .B1( u0_u8_u2_n153 ) , .ZN( u0_u8_u2_n164 ) );
  NOR4_X1 u0_u8_u2_U5 (.A4( u0_u8_u2_n124 ) , .A3( u0_u8_u2_n125 ) , .A2( u0_u8_u2_n126 ) , .A1( u0_u8_u2_n127 ) , .ZN( u0_u8_u2_n128 ) );
  NAND2_X1 u0_u8_u2_U50 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n107 ) , .ZN( u0_u8_u2_n155 ) );
  NAND2_X1 u0_u8_u2_U51 (.A2( u0_u8_u2_n105 ) , .A1( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n143 ) );
  NAND2_X1 u0_u8_u2_U52 (.A1( u0_u8_u2_n104 ) , .A2( u0_u8_u2_n106 ) , .ZN( u0_u8_u2_n152 ) );
  NAND2_X1 u0_u8_u2_U53 (.A1( u0_u8_u2_n100 ) , .A2( u0_u8_u2_n105 ) , .ZN( u0_u8_u2_n132 ) );
  INV_X1 u0_u8_u2_U54 (.A( u0_u8_u2_n140 ) , .ZN( u0_u8_u2_n168 ) );
  INV_X1 u0_u8_u2_U55 (.A( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n167 ) );
  NAND2_X1 u0_u8_u2_U56 (.A1( u0_u8_u2_n102 ) , .A2( u0_u8_u2_n106 ) , .ZN( u0_u8_u2_n113 ) );
  NAND2_X1 u0_u8_u2_U57 (.A1( u0_u8_u2_n106 ) , .A2( u0_u8_u2_n107 ) , .ZN( u0_u8_u2_n131 ) );
  NAND2_X1 u0_u8_u2_U58 (.A1( u0_u8_u2_n103 ) , .A2( u0_u8_u2_n107 ) , .ZN( u0_u8_u2_n139 ) );
  NAND2_X1 u0_u8_u2_U59 (.A1( u0_u8_u2_n103 ) , .A2( u0_u8_u2_n105 ) , .ZN( u0_u8_u2_n133 ) );
  AOI21_X1 u0_u8_u2_U6 (.B2( u0_u8_u2_n119 ) , .ZN( u0_u8_u2_n127 ) , .A( u0_u8_u2_n137 ) , .B1( u0_u8_u2_n155 ) );
  NAND2_X1 u0_u8_u2_U60 (.A1( u0_u8_u2_n102 ) , .A2( u0_u8_u2_n103 ) , .ZN( u0_u8_u2_n154 ) );
  NAND2_X1 u0_u8_u2_U61 (.A2( u0_u8_u2_n103 ) , .A1( u0_u8_u2_n104 ) , .ZN( u0_u8_u2_n119 ) );
  NAND2_X1 u0_u8_u2_U62 (.A2( u0_u8_u2_n107 ) , .A1( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n123 ) );
  NAND2_X1 u0_u8_u2_U63 (.A1( u0_u8_u2_n104 ) , .A2( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n122 ) );
  INV_X1 u0_u8_u2_U64 (.A( u0_u8_u2_n114 ) , .ZN( u0_u8_u2_n172 ) );
  NAND2_X1 u0_u8_u2_U65 (.A2( u0_u8_u2_n100 ) , .A1( u0_u8_u2_n102 ) , .ZN( u0_u8_u2_n116 ) );
  NAND2_X1 u0_u8_u2_U66 (.A1( u0_u8_u2_n102 ) , .A2( u0_u8_u2_n108 ) , .ZN( u0_u8_u2_n120 ) );
  NAND2_X1 u0_u8_u2_U67 (.A2( u0_u8_u2_n105 ) , .A1( u0_u8_u2_n106 ) , .ZN( u0_u8_u2_n117 ) );
  INV_X1 u0_u8_u2_U68 (.ZN( u0_u8_u2_n187 ) , .A( u0_u8_u2_n99 ) );
  OAI21_X1 u0_u8_u2_U69 (.B1( u0_u8_u2_n137 ) , .B2( u0_u8_u2_n143 ) , .A( u0_u8_u2_n98 ) , .ZN( u0_u8_u2_n99 ) );
  AOI21_X1 u0_u8_u2_U7 (.ZN( u0_u8_u2_n124 ) , .B1( u0_u8_u2_n131 ) , .B2( u0_u8_u2_n143 ) , .A( u0_u8_u2_n172 ) );
  NOR2_X1 u0_u8_u2_U70 (.A2( u0_u8_X_16 ) , .ZN( u0_u8_u2_n140 ) , .A1( u0_u8_u2_n166 ) );
  NOR2_X1 u0_u8_u2_U71 (.A2( u0_u8_X_13 ) , .A1( u0_u8_X_14 ) , .ZN( u0_u8_u2_n100 ) );
  NOR2_X1 u0_u8_u2_U72 (.A2( u0_u8_X_16 ) , .A1( u0_u8_X_17 ) , .ZN( u0_u8_u2_n138 ) );
  NOR2_X1 u0_u8_u2_U73 (.A2( u0_u8_X_15 ) , .A1( u0_u8_X_18 ) , .ZN( u0_u8_u2_n104 ) );
  NOR2_X1 u0_u8_u2_U74 (.A2( u0_u8_X_14 ) , .ZN( u0_u8_u2_n103 ) , .A1( u0_u8_u2_n174 ) );
  NOR2_X1 u0_u8_u2_U75 (.A2( u0_u8_X_15 ) , .ZN( u0_u8_u2_n102 ) , .A1( u0_u8_u2_n165 ) );
  NOR2_X1 u0_u8_u2_U76 (.A2( u0_u8_X_17 ) , .ZN( u0_u8_u2_n114 ) , .A1( u0_u8_u2_n169 ) );
  AND2_X1 u0_u8_u2_U77 (.A1( u0_u8_X_15 ) , .ZN( u0_u8_u2_n105 ) , .A2( u0_u8_u2_n165 ) );
  AND2_X1 u0_u8_u2_U78 (.A2( u0_u8_X_15 ) , .A1( u0_u8_X_18 ) , .ZN( u0_u8_u2_n107 ) );
  AND2_X1 u0_u8_u2_U79 (.A1( u0_u8_X_14 ) , .ZN( u0_u8_u2_n106 ) , .A2( u0_u8_u2_n174 ) );
  AOI21_X1 u0_u8_u2_U8 (.B2( u0_u8_u2_n120 ) , .B1( u0_u8_u2_n121 ) , .ZN( u0_u8_u2_n126 ) , .A( u0_u8_u2_n167 ) );
  AND2_X1 u0_u8_u2_U80 (.A1( u0_u8_X_13 ) , .A2( u0_u8_X_14 ) , .ZN( u0_u8_u2_n108 ) );
  INV_X1 u0_u8_u2_U81 (.A( u0_u8_X_16 ) , .ZN( u0_u8_u2_n169 ) );
  INV_X1 u0_u8_u2_U82 (.A( u0_u8_X_17 ) , .ZN( u0_u8_u2_n166 ) );
  INV_X1 u0_u8_u2_U83 (.A( u0_u8_X_13 ) , .ZN( u0_u8_u2_n174 ) );
  INV_X1 u0_u8_u2_U84 (.A( u0_u8_X_18 ) , .ZN( u0_u8_u2_n165 ) );
  NAND4_X1 u0_u8_u2_U85 (.ZN( u0_out8_30 ) , .A4( u0_u8_u2_n147 ) , .A3( u0_u8_u2_n148 ) , .A2( u0_u8_u2_n149 ) , .A1( u0_u8_u2_n187 ) );
  NOR3_X1 u0_u8_u2_U86 (.A3( u0_u8_u2_n144 ) , .A2( u0_u8_u2_n145 ) , .A1( u0_u8_u2_n146 ) , .ZN( u0_u8_u2_n147 ) );
  AOI21_X1 u0_u8_u2_U87 (.B2( u0_u8_u2_n138 ) , .ZN( u0_u8_u2_n148 ) , .A( u0_u8_u2_n162 ) , .B1( u0_u8_u2_n182 ) );
  NAND4_X1 u0_u8_u2_U88 (.ZN( u0_out8_24 ) , .A4( u0_u8_u2_n111 ) , .A3( u0_u8_u2_n112 ) , .A1( u0_u8_u2_n130 ) , .A2( u0_u8_u2_n187 ) );
  AOI221_X1 u0_u8_u2_U89 (.A( u0_u8_u2_n109 ) , .B1( u0_u8_u2_n110 ) , .ZN( u0_u8_u2_n111 ) , .C1( u0_u8_u2_n134 ) , .C2( u0_u8_u2_n170 ) , .B2( u0_u8_u2_n173 ) );
  OAI22_X1 u0_u8_u2_U9 (.ZN( u0_u8_u2_n109 ) , .A2( u0_u8_u2_n113 ) , .B2( u0_u8_u2_n133 ) , .B1( u0_u8_u2_n167 ) , .A1( u0_u8_u2_n168 ) );
  AOI21_X1 u0_u8_u2_U90 (.ZN( u0_u8_u2_n112 ) , .B2( u0_u8_u2_n156 ) , .A( u0_u8_u2_n164 ) , .B1( u0_u8_u2_n181 ) );
  NAND4_X1 u0_u8_u2_U91 (.ZN( u0_out8_16 ) , .A4( u0_u8_u2_n128 ) , .A3( u0_u8_u2_n129 ) , .A1( u0_u8_u2_n130 ) , .A2( u0_u8_u2_n186 ) );
  AOI22_X1 u0_u8_u2_U92 (.A2( u0_u8_u2_n118 ) , .ZN( u0_u8_u2_n129 ) , .A1( u0_u8_u2_n140 ) , .B1( u0_u8_u2_n157 ) , .B2( u0_u8_u2_n170 ) );
  INV_X1 u0_u8_u2_U93 (.A( u0_u8_u2_n163 ) , .ZN( u0_u8_u2_n186 ) );
  OR4_X1 u0_u8_u2_U94 (.ZN( u0_out8_6 ) , .A4( u0_u8_u2_n161 ) , .A3( u0_u8_u2_n162 ) , .A2( u0_u8_u2_n163 ) , .A1( u0_u8_u2_n164 ) );
  OR3_X1 u0_u8_u2_U95 (.A2( u0_u8_u2_n159 ) , .A1( u0_u8_u2_n160 ) , .ZN( u0_u8_u2_n161 ) , .A3( u0_u8_u2_n183 ) );
  AOI21_X1 u0_u8_u2_U96 (.B2( u0_u8_u2_n154 ) , .B1( u0_u8_u2_n155 ) , .ZN( u0_u8_u2_n159 ) , .A( u0_u8_u2_n167 ) );
  NAND3_X1 u0_u8_u2_U97 (.A2( u0_u8_u2_n117 ) , .A1( u0_u8_u2_n122 ) , .A3( u0_u8_u2_n123 ) , .ZN( u0_u8_u2_n134 ) );
  NAND3_X1 u0_u8_u2_U98 (.ZN( u0_u8_u2_n110 ) , .A2( u0_u8_u2_n131 ) , .A3( u0_u8_u2_n139 ) , .A1( u0_u8_u2_n154 ) );
  NAND3_X1 u0_u8_u2_U99 (.A2( u0_u8_u2_n100 ) , .ZN( u0_u8_u2_n101 ) , .A1( u0_u8_u2_n104 ) , .A3( u0_u8_u2_n114 ) );
  OAI22_X1 u0_u8_u3_U10 (.B1( u0_u8_u3_n113 ) , .A2( u0_u8_u3_n135 ) , .A1( u0_u8_u3_n150 ) , .B2( u0_u8_u3_n164 ) , .ZN( u0_u8_u3_n98 ) );
  OAI211_X1 u0_u8_u3_U11 (.B( u0_u8_u3_n106 ) , .ZN( u0_u8_u3_n119 ) , .C2( u0_u8_u3_n128 ) , .C1( u0_u8_u3_n167 ) , .A( u0_u8_u3_n181 ) );
  AOI221_X1 u0_u8_u3_U12 (.C1( u0_u8_u3_n105 ) , .ZN( u0_u8_u3_n106 ) , .A( u0_u8_u3_n131 ) , .B2( u0_u8_u3_n132 ) , .C2( u0_u8_u3_n133 ) , .B1( u0_u8_u3_n169 ) );
  INV_X1 u0_u8_u3_U13 (.ZN( u0_u8_u3_n181 ) , .A( u0_u8_u3_n98 ) );
  NAND2_X1 u0_u8_u3_U14 (.ZN( u0_u8_u3_n105 ) , .A2( u0_u8_u3_n130 ) , .A1( u0_u8_u3_n155 ) );
  AOI22_X1 u0_u8_u3_U15 (.B1( u0_u8_u3_n115 ) , .A2( u0_u8_u3_n116 ) , .ZN( u0_u8_u3_n123 ) , .B2( u0_u8_u3_n133 ) , .A1( u0_u8_u3_n169 ) );
  NAND2_X1 u0_u8_u3_U16 (.ZN( u0_u8_u3_n116 ) , .A2( u0_u8_u3_n151 ) , .A1( u0_u8_u3_n182 ) );
  NOR2_X1 u0_u8_u3_U17 (.ZN( u0_u8_u3_n126 ) , .A2( u0_u8_u3_n150 ) , .A1( u0_u8_u3_n164 ) );
  AOI21_X1 u0_u8_u3_U18 (.ZN( u0_u8_u3_n112 ) , .B2( u0_u8_u3_n146 ) , .B1( u0_u8_u3_n155 ) , .A( u0_u8_u3_n167 ) );
  NAND2_X1 u0_u8_u3_U19 (.A1( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n142 ) , .A2( u0_u8_u3_n164 ) );
  NAND2_X1 u0_u8_u3_U20 (.ZN( u0_u8_u3_n132 ) , .A2( u0_u8_u3_n152 ) , .A1( u0_u8_u3_n156 ) );
  AND2_X1 u0_u8_u3_U21 (.A2( u0_u8_u3_n113 ) , .A1( u0_u8_u3_n114 ) , .ZN( u0_u8_u3_n151 ) );
  INV_X1 u0_u8_u3_U22 (.A( u0_u8_u3_n133 ) , .ZN( u0_u8_u3_n165 ) );
  INV_X1 u0_u8_u3_U23 (.A( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n170 ) );
  NAND2_X1 u0_u8_u3_U24 (.A1( u0_u8_u3_n107 ) , .A2( u0_u8_u3_n108 ) , .ZN( u0_u8_u3_n140 ) );
  NAND2_X1 u0_u8_u3_U25 (.ZN( u0_u8_u3_n117 ) , .A1( u0_u8_u3_n124 ) , .A2( u0_u8_u3_n148 ) );
  NAND2_X1 u0_u8_u3_U26 (.ZN( u0_u8_u3_n143 ) , .A1( u0_u8_u3_n165 ) , .A2( u0_u8_u3_n167 ) );
  INV_X1 u0_u8_u3_U27 (.A( u0_u8_u3_n130 ) , .ZN( u0_u8_u3_n177 ) );
  INV_X1 u0_u8_u3_U28 (.A( u0_u8_u3_n128 ) , .ZN( u0_u8_u3_n176 ) );
  INV_X1 u0_u8_u3_U29 (.A( u0_u8_u3_n155 ) , .ZN( u0_u8_u3_n174 ) );
  INV_X1 u0_u8_u3_U3 (.A( u0_u8_u3_n129 ) , .ZN( u0_u8_u3_n183 ) );
  INV_X1 u0_u8_u3_U30 (.A( u0_u8_u3_n139 ) , .ZN( u0_u8_u3_n185 ) );
  NOR2_X1 u0_u8_u3_U31 (.ZN( u0_u8_u3_n135 ) , .A2( u0_u8_u3_n141 ) , .A1( u0_u8_u3_n169 ) );
  OAI222_X1 u0_u8_u3_U32 (.C2( u0_u8_u3_n107 ) , .A2( u0_u8_u3_n108 ) , .B1( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n138 ) , .B2( u0_u8_u3_n146 ) , .C1( u0_u8_u3_n154 ) , .A1( u0_u8_u3_n164 ) );
  NOR4_X1 u0_u8_u3_U33 (.A4( u0_u8_u3_n157 ) , .A3( u0_u8_u3_n158 ) , .A2( u0_u8_u3_n159 ) , .A1( u0_u8_u3_n160 ) , .ZN( u0_u8_u3_n161 ) );
  AOI21_X1 u0_u8_u3_U34 (.B2( u0_u8_u3_n152 ) , .B1( u0_u8_u3_n153 ) , .ZN( u0_u8_u3_n158 ) , .A( u0_u8_u3_n164 ) );
  AOI21_X1 u0_u8_u3_U35 (.A( u0_u8_u3_n149 ) , .B2( u0_u8_u3_n150 ) , .B1( u0_u8_u3_n151 ) , .ZN( u0_u8_u3_n159 ) );
  AOI21_X1 u0_u8_u3_U36 (.A( u0_u8_u3_n154 ) , .B2( u0_u8_u3_n155 ) , .B1( u0_u8_u3_n156 ) , .ZN( u0_u8_u3_n157 ) );
  AOI211_X1 u0_u8_u3_U37 (.ZN( u0_u8_u3_n109 ) , .A( u0_u8_u3_n119 ) , .C2( u0_u8_u3_n129 ) , .B( u0_u8_u3_n138 ) , .C1( u0_u8_u3_n141 ) );
  AOI211_X1 u0_u8_u3_U38 (.B( u0_u8_u3_n119 ) , .A( u0_u8_u3_n120 ) , .C2( u0_u8_u3_n121 ) , .ZN( u0_u8_u3_n122 ) , .C1( u0_u8_u3_n179 ) );
  INV_X1 u0_u8_u3_U39 (.A( u0_u8_u3_n156 ) , .ZN( u0_u8_u3_n179 ) );
  INV_X1 u0_u8_u3_U4 (.A( u0_u8_u3_n140 ) , .ZN( u0_u8_u3_n182 ) );
  OAI22_X1 u0_u8_u3_U40 (.B1( u0_u8_u3_n118 ) , .ZN( u0_u8_u3_n120 ) , .A1( u0_u8_u3_n135 ) , .B2( u0_u8_u3_n154 ) , .A2( u0_u8_u3_n178 ) );
  AND3_X1 u0_u8_u3_U41 (.ZN( u0_u8_u3_n118 ) , .A2( u0_u8_u3_n124 ) , .A1( u0_u8_u3_n144 ) , .A3( u0_u8_u3_n152 ) );
  INV_X1 u0_u8_u3_U42 (.A( u0_u8_u3_n121 ) , .ZN( u0_u8_u3_n164 ) );
  NAND2_X1 u0_u8_u3_U43 (.ZN( u0_u8_u3_n133 ) , .A1( u0_u8_u3_n154 ) , .A2( u0_u8_u3_n164 ) );
  OAI211_X1 u0_u8_u3_U44 (.B( u0_u8_u3_n127 ) , .ZN( u0_u8_u3_n139 ) , .C1( u0_u8_u3_n150 ) , .C2( u0_u8_u3_n154 ) , .A( u0_u8_u3_n184 ) );
  INV_X1 u0_u8_u3_U45 (.A( u0_u8_u3_n125 ) , .ZN( u0_u8_u3_n184 ) );
  AOI221_X1 u0_u8_u3_U46 (.A( u0_u8_u3_n126 ) , .ZN( u0_u8_u3_n127 ) , .C2( u0_u8_u3_n132 ) , .C1( u0_u8_u3_n169 ) , .B2( u0_u8_u3_n170 ) , .B1( u0_u8_u3_n174 ) );
  OAI22_X1 u0_u8_u3_U47 (.A1( u0_u8_u3_n124 ) , .ZN( u0_u8_u3_n125 ) , .B2( u0_u8_u3_n145 ) , .A2( u0_u8_u3_n165 ) , .B1( u0_u8_u3_n167 ) );
  NOR2_X1 u0_u8_u3_U48 (.A1( u0_u8_u3_n113 ) , .ZN( u0_u8_u3_n131 ) , .A2( u0_u8_u3_n154 ) );
  NAND2_X1 u0_u8_u3_U49 (.A1( u0_u8_u3_n103 ) , .ZN( u0_u8_u3_n150 ) , .A2( u0_u8_u3_n99 ) );
  INV_X1 u0_u8_u3_U5 (.A( u0_u8_u3_n117 ) , .ZN( u0_u8_u3_n178 ) );
  NAND2_X1 u0_u8_u3_U50 (.A2( u0_u8_u3_n102 ) , .ZN( u0_u8_u3_n155 ) , .A1( u0_u8_u3_n97 ) );
  INV_X1 u0_u8_u3_U51 (.A( u0_u8_u3_n141 ) , .ZN( u0_u8_u3_n167 ) );
  AOI21_X1 u0_u8_u3_U52 (.B2( u0_u8_u3_n114 ) , .B1( u0_u8_u3_n146 ) , .A( u0_u8_u3_n154 ) , .ZN( u0_u8_u3_n94 ) );
  AOI21_X1 u0_u8_u3_U53 (.ZN( u0_u8_u3_n110 ) , .B2( u0_u8_u3_n142 ) , .B1( u0_u8_u3_n186 ) , .A( u0_u8_u3_n95 ) );
  INV_X1 u0_u8_u3_U54 (.A( u0_u8_u3_n145 ) , .ZN( u0_u8_u3_n186 ) );
  AOI21_X1 u0_u8_u3_U55 (.B1( u0_u8_u3_n124 ) , .A( u0_u8_u3_n149 ) , .B2( u0_u8_u3_n155 ) , .ZN( u0_u8_u3_n95 ) );
  INV_X1 u0_u8_u3_U56 (.A( u0_u8_u3_n149 ) , .ZN( u0_u8_u3_n169 ) );
  NAND2_X1 u0_u8_u3_U57 (.ZN( u0_u8_u3_n124 ) , .A1( u0_u8_u3_n96 ) , .A2( u0_u8_u3_n97 ) );
  NAND2_X1 u0_u8_u3_U58 (.A2( u0_u8_u3_n100 ) , .ZN( u0_u8_u3_n146 ) , .A1( u0_u8_u3_n96 ) );
  NAND2_X1 u0_u8_u3_U59 (.A1( u0_u8_u3_n101 ) , .ZN( u0_u8_u3_n145 ) , .A2( u0_u8_u3_n99 ) );
  AOI221_X1 u0_u8_u3_U6 (.A( u0_u8_u3_n131 ) , .C2( u0_u8_u3_n132 ) , .C1( u0_u8_u3_n133 ) , .ZN( u0_u8_u3_n134 ) , .B1( u0_u8_u3_n143 ) , .B2( u0_u8_u3_n177 ) );
  NAND2_X1 u0_u8_u3_U60 (.A1( u0_u8_u3_n100 ) , .ZN( u0_u8_u3_n156 ) , .A2( u0_u8_u3_n99 ) );
  NAND2_X1 u0_u8_u3_U61 (.A2( u0_u8_u3_n101 ) , .A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n148 ) );
  NAND2_X1 u0_u8_u3_U62 (.A1( u0_u8_u3_n100 ) , .A2( u0_u8_u3_n102 ) , .ZN( u0_u8_u3_n128 ) );
  NAND2_X1 u0_u8_u3_U63 (.A2( u0_u8_u3_n101 ) , .A1( u0_u8_u3_n102 ) , .ZN( u0_u8_u3_n152 ) );
  NAND2_X1 u0_u8_u3_U64 (.A2( u0_u8_u3_n101 ) , .ZN( u0_u8_u3_n114 ) , .A1( u0_u8_u3_n96 ) );
  NAND2_X1 u0_u8_u3_U65 (.ZN( u0_u8_u3_n107 ) , .A1( u0_u8_u3_n97 ) , .A2( u0_u8_u3_n99 ) );
  NAND2_X1 u0_u8_u3_U66 (.A2( u0_u8_u3_n100 ) , .A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n113 ) );
  NAND2_X1 u0_u8_u3_U67 (.A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n153 ) , .A2( u0_u8_u3_n97 ) );
  NAND2_X1 u0_u8_u3_U68 (.A2( u0_u8_u3_n103 ) , .A1( u0_u8_u3_n104 ) , .ZN( u0_u8_u3_n130 ) );
  NAND2_X1 u0_u8_u3_U69 (.A2( u0_u8_u3_n103 ) , .ZN( u0_u8_u3_n144 ) , .A1( u0_u8_u3_n96 ) );
  OAI22_X1 u0_u8_u3_U7 (.B2( u0_u8_u3_n147 ) , .A2( u0_u8_u3_n148 ) , .ZN( u0_u8_u3_n160 ) , .B1( u0_u8_u3_n165 ) , .A1( u0_u8_u3_n168 ) );
  NAND2_X1 u0_u8_u3_U70 (.A1( u0_u8_u3_n102 ) , .A2( u0_u8_u3_n103 ) , .ZN( u0_u8_u3_n108 ) );
  NOR2_X1 u0_u8_u3_U71 (.A2( u0_u8_X_19 ) , .A1( u0_u8_X_20 ) , .ZN( u0_u8_u3_n99 ) );
  NOR2_X1 u0_u8_u3_U72 (.A2( u0_u8_X_21 ) , .A1( u0_u8_X_24 ) , .ZN( u0_u8_u3_n103 ) );
  NOR2_X1 u0_u8_u3_U73 (.A2( u0_u8_X_24 ) , .A1( u0_u8_u3_n171 ) , .ZN( u0_u8_u3_n97 ) );
  NOR2_X1 u0_u8_u3_U74 (.A2( u0_u8_X_23 ) , .ZN( u0_u8_u3_n141 ) , .A1( u0_u8_u3_n166 ) );
  NOR2_X1 u0_u8_u3_U75 (.A2( u0_u8_X_19 ) , .A1( u0_u8_u3_n172 ) , .ZN( u0_u8_u3_n96 ) );
  NAND2_X1 u0_u8_u3_U76 (.A1( u0_u8_X_22 ) , .A2( u0_u8_X_23 ) , .ZN( u0_u8_u3_n154 ) );
  NAND2_X1 u0_u8_u3_U77 (.A1( u0_u8_X_23 ) , .ZN( u0_u8_u3_n149 ) , .A2( u0_u8_u3_n166 ) );
  NOR2_X1 u0_u8_u3_U78 (.A2( u0_u8_X_22 ) , .A1( u0_u8_X_23 ) , .ZN( u0_u8_u3_n121 ) );
  AND2_X1 u0_u8_u3_U79 (.A1( u0_u8_X_24 ) , .ZN( u0_u8_u3_n101 ) , .A2( u0_u8_u3_n171 ) );
  AND3_X1 u0_u8_u3_U8 (.A3( u0_u8_u3_n144 ) , .A2( u0_u8_u3_n145 ) , .A1( u0_u8_u3_n146 ) , .ZN( u0_u8_u3_n147 ) );
  AND2_X1 u0_u8_u3_U80 (.A1( u0_u8_X_19 ) , .ZN( u0_u8_u3_n102 ) , .A2( u0_u8_u3_n172 ) );
  AND2_X1 u0_u8_u3_U81 (.A1( u0_u8_X_21 ) , .A2( u0_u8_X_24 ) , .ZN( u0_u8_u3_n100 ) );
  AND2_X1 u0_u8_u3_U82 (.A2( u0_u8_X_19 ) , .A1( u0_u8_X_20 ) , .ZN( u0_u8_u3_n104 ) );
  INV_X1 u0_u8_u3_U83 (.A( u0_u8_X_22 ) , .ZN( u0_u8_u3_n166 ) );
  INV_X1 u0_u8_u3_U84 (.A( u0_u8_X_21 ) , .ZN( u0_u8_u3_n171 ) );
  INV_X1 u0_u8_u3_U85 (.A( u0_u8_X_20 ) , .ZN( u0_u8_u3_n172 ) );
  OR4_X1 u0_u8_u3_U86 (.ZN( u0_out8_10 ) , .A4( u0_u8_u3_n136 ) , .A3( u0_u8_u3_n137 ) , .A1( u0_u8_u3_n138 ) , .A2( u0_u8_u3_n139 ) );
  OAI222_X1 u0_u8_u3_U87 (.C1( u0_u8_u3_n128 ) , .ZN( u0_u8_u3_n137 ) , .B1( u0_u8_u3_n148 ) , .A2( u0_u8_u3_n150 ) , .B2( u0_u8_u3_n154 ) , .C2( u0_u8_u3_n164 ) , .A1( u0_u8_u3_n167 ) );
  OAI221_X1 u0_u8_u3_U88 (.A( u0_u8_u3_n134 ) , .B2( u0_u8_u3_n135 ) , .ZN( u0_u8_u3_n136 ) , .C1( u0_u8_u3_n149 ) , .B1( u0_u8_u3_n151 ) , .C2( u0_u8_u3_n183 ) );
  NAND4_X1 u0_u8_u3_U89 (.ZN( u0_out8_26 ) , .A4( u0_u8_u3_n109 ) , .A3( u0_u8_u3_n110 ) , .A2( u0_u8_u3_n111 ) , .A1( u0_u8_u3_n173 ) );
  INV_X1 u0_u8_u3_U9 (.A( u0_u8_u3_n143 ) , .ZN( u0_u8_u3_n168 ) );
  INV_X1 u0_u8_u3_U90 (.ZN( u0_u8_u3_n173 ) , .A( u0_u8_u3_n94 ) );
  OAI21_X1 u0_u8_u3_U91 (.ZN( u0_u8_u3_n111 ) , .B2( u0_u8_u3_n117 ) , .A( u0_u8_u3_n133 ) , .B1( u0_u8_u3_n176 ) );
  NAND4_X1 u0_u8_u3_U92 (.ZN( u0_out8_20 ) , .A4( u0_u8_u3_n122 ) , .A3( u0_u8_u3_n123 ) , .A1( u0_u8_u3_n175 ) , .A2( u0_u8_u3_n180 ) );
  INV_X1 u0_u8_u3_U93 (.A( u0_u8_u3_n126 ) , .ZN( u0_u8_u3_n180 ) );
  INV_X1 u0_u8_u3_U94 (.A( u0_u8_u3_n112 ) , .ZN( u0_u8_u3_n175 ) );
  NAND4_X1 u0_u8_u3_U95 (.ZN( u0_out8_1 ) , .A4( u0_u8_u3_n161 ) , .A3( u0_u8_u3_n162 ) , .A2( u0_u8_u3_n163 ) , .A1( u0_u8_u3_n185 ) );
  NAND2_X1 u0_u8_u3_U96 (.ZN( u0_u8_u3_n163 ) , .A2( u0_u8_u3_n170 ) , .A1( u0_u8_u3_n176 ) );
  AOI22_X1 u0_u8_u3_U97 (.B2( u0_u8_u3_n140 ) , .B1( u0_u8_u3_n141 ) , .A2( u0_u8_u3_n142 ) , .ZN( u0_u8_u3_n162 ) , .A1( u0_u8_u3_n177 ) );
  NAND3_X1 u0_u8_u3_U98 (.A1( u0_u8_u3_n114 ) , .ZN( u0_u8_u3_n115 ) , .A2( u0_u8_u3_n145 ) , .A3( u0_u8_u3_n153 ) );
  NAND3_X1 u0_u8_u3_U99 (.ZN( u0_u8_u3_n129 ) , .A2( u0_u8_u3_n144 ) , .A1( u0_u8_u3_n153 ) , .A3( u0_u8_u3_n182 ) );
  OAI22_X1 u0_u8_u4_U10 (.B2( u0_u8_u4_n135 ) , .ZN( u0_u8_u4_n137 ) , .B1( u0_u8_u4_n153 ) , .A1( u0_u8_u4_n155 ) , .A2( u0_u8_u4_n171 ) );
  AND3_X1 u0_u8_u4_U11 (.A2( u0_u8_u4_n134 ) , .ZN( u0_u8_u4_n135 ) , .A3( u0_u8_u4_n145 ) , .A1( u0_u8_u4_n157 ) );
  NAND2_X1 u0_u8_u4_U12 (.ZN( u0_u8_u4_n132 ) , .A2( u0_u8_u4_n170 ) , .A1( u0_u8_u4_n173 ) );
  AOI21_X1 u0_u8_u4_U13 (.B2( u0_u8_u4_n160 ) , .B1( u0_u8_u4_n161 ) , .ZN( u0_u8_u4_n162 ) , .A( u0_u8_u4_n170 ) );
  AOI21_X1 u0_u8_u4_U14 (.ZN( u0_u8_u4_n107 ) , .B2( u0_u8_u4_n143 ) , .A( u0_u8_u4_n174 ) , .B1( u0_u8_u4_n184 ) );
  AOI21_X1 u0_u8_u4_U15 (.B2( u0_u8_u4_n158 ) , .B1( u0_u8_u4_n159 ) , .ZN( u0_u8_u4_n163 ) , .A( u0_u8_u4_n174 ) );
  AOI21_X1 u0_u8_u4_U16 (.A( u0_u8_u4_n153 ) , .B2( u0_u8_u4_n154 ) , .B1( u0_u8_u4_n155 ) , .ZN( u0_u8_u4_n165 ) );
  AOI21_X1 u0_u8_u4_U17 (.A( u0_u8_u4_n156 ) , .B2( u0_u8_u4_n157 ) , .ZN( u0_u8_u4_n164 ) , .B1( u0_u8_u4_n184 ) );
  INV_X1 u0_u8_u4_U18 (.A( u0_u8_u4_n138 ) , .ZN( u0_u8_u4_n170 ) );
  AND2_X1 u0_u8_u4_U19 (.A2( u0_u8_u4_n120 ) , .ZN( u0_u8_u4_n155 ) , .A1( u0_u8_u4_n160 ) );
  INV_X1 u0_u8_u4_U20 (.A( u0_u8_u4_n156 ) , .ZN( u0_u8_u4_n175 ) );
  NAND2_X1 u0_u8_u4_U21 (.A2( u0_u8_u4_n118 ) , .ZN( u0_u8_u4_n131 ) , .A1( u0_u8_u4_n147 ) );
  NAND2_X1 u0_u8_u4_U22 (.A1( u0_u8_u4_n119 ) , .A2( u0_u8_u4_n120 ) , .ZN( u0_u8_u4_n130 ) );
  NAND2_X1 u0_u8_u4_U23 (.ZN( u0_u8_u4_n117 ) , .A2( u0_u8_u4_n118 ) , .A1( u0_u8_u4_n148 ) );
  NAND2_X1 u0_u8_u4_U24 (.ZN( u0_u8_u4_n129 ) , .A1( u0_u8_u4_n134 ) , .A2( u0_u8_u4_n148 ) );
  AND3_X1 u0_u8_u4_U25 (.A1( u0_u8_u4_n119 ) , .A2( u0_u8_u4_n143 ) , .A3( u0_u8_u4_n154 ) , .ZN( u0_u8_u4_n161 ) );
  AND2_X1 u0_u8_u4_U26 (.A1( u0_u8_u4_n145 ) , .A2( u0_u8_u4_n147 ) , .ZN( u0_u8_u4_n159 ) );
  OR3_X1 u0_u8_u4_U27 (.A3( u0_u8_u4_n114 ) , .A2( u0_u8_u4_n115 ) , .A1( u0_u8_u4_n116 ) , .ZN( u0_u8_u4_n136 ) );
  AOI21_X1 u0_u8_u4_U28 (.A( u0_u8_u4_n113 ) , .ZN( u0_u8_u4_n116 ) , .B2( u0_u8_u4_n173 ) , .B1( u0_u8_u4_n174 ) );
  AOI21_X1 u0_u8_u4_U29 (.ZN( u0_u8_u4_n115 ) , .B2( u0_u8_u4_n145 ) , .B1( u0_u8_u4_n146 ) , .A( u0_u8_u4_n156 ) );
  NOR2_X1 u0_u8_u4_U3 (.ZN( u0_u8_u4_n121 ) , .A1( u0_u8_u4_n181 ) , .A2( u0_u8_u4_n182 ) );
  OAI22_X1 u0_u8_u4_U30 (.ZN( u0_u8_u4_n114 ) , .A2( u0_u8_u4_n121 ) , .B1( u0_u8_u4_n160 ) , .B2( u0_u8_u4_n170 ) , .A1( u0_u8_u4_n171 ) );
  INV_X1 u0_u8_u4_U31 (.A( u0_u8_u4_n158 ) , .ZN( u0_u8_u4_n182 ) );
  INV_X1 u0_u8_u4_U32 (.ZN( u0_u8_u4_n181 ) , .A( u0_u8_u4_n96 ) );
  INV_X1 u0_u8_u4_U33 (.A( u0_u8_u4_n144 ) , .ZN( u0_u8_u4_n179 ) );
  INV_X1 u0_u8_u4_U34 (.A( u0_u8_u4_n157 ) , .ZN( u0_u8_u4_n178 ) );
  NAND2_X1 u0_u8_u4_U35 (.A2( u0_u8_u4_n154 ) , .A1( u0_u8_u4_n96 ) , .ZN( u0_u8_u4_n97 ) );
  INV_X1 u0_u8_u4_U36 (.ZN( u0_u8_u4_n186 ) , .A( u0_u8_u4_n95 ) );
  OAI221_X1 u0_u8_u4_U37 (.C1( u0_u8_u4_n134 ) , .B1( u0_u8_u4_n158 ) , .B2( u0_u8_u4_n171 ) , .C2( u0_u8_u4_n173 ) , .A( u0_u8_u4_n94 ) , .ZN( u0_u8_u4_n95 ) );
  AOI222_X1 u0_u8_u4_U38 (.B2( u0_u8_u4_n132 ) , .A1( u0_u8_u4_n138 ) , .C2( u0_u8_u4_n175 ) , .A2( u0_u8_u4_n179 ) , .C1( u0_u8_u4_n181 ) , .B1( u0_u8_u4_n185 ) , .ZN( u0_u8_u4_n94 ) );
  INV_X1 u0_u8_u4_U39 (.A( u0_u8_u4_n113 ) , .ZN( u0_u8_u4_n185 ) );
  INV_X1 u0_u8_u4_U4 (.A( u0_u8_u4_n117 ) , .ZN( u0_u8_u4_n184 ) );
  INV_X1 u0_u8_u4_U40 (.A( u0_u8_u4_n143 ) , .ZN( u0_u8_u4_n183 ) );
  NOR2_X1 u0_u8_u4_U41 (.ZN( u0_u8_u4_n138 ) , .A1( u0_u8_u4_n168 ) , .A2( u0_u8_u4_n169 ) );
  NOR2_X1 u0_u8_u4_U42 (.A1( u0_u8_u4_n150 ) , .A2( u0_u8_u4_n152 ) , .ZN( u0_u8_u4_n153 ) );
  NOR2_X1 u0_u8_u4_U43 (.A2( u0_u8_u4_n128 ) , .A1( u0_u8_u4_n138 ) , .ZN( u0_u8_u4_n156 ) );
  AOI22_X1 u0_u8_u4_U44 (.B2( u0_u8_u4_n122 ) , .A1( u0_u8_u4_n123 ) , .ZN( u0_u8_u4_n124 ) , .B1( u0_u8_u4_n128 ) , .A2( u0_u8_u4_n172 ) );
  INV_X1 u0_u8_u4_U45 (.A( u0_u8_u4_n153 ) , .ZN( u0_u8_u4_n172 ) );
  NAND2_X1 u0_u8_u4_U46 (.A2( u0_u8_u4_n120 ) , .ZN( u0_u8_u4_n123 ) , .A1( u0_u8_u4_n161 ) );
  AOI22_X1 u0_u8_u4_U47 (.B2( u0_u8_u4_n132 ) , .A2( u0_u8_u4_n133 ) , .ZN( u0_u8_u4_n140 ) , .A1( u0_u8_u4_n150 ) , .B1( u0_u8_u4_n179 ) );
  NAND2_X1 u0_u8_u4_U48 (.ZN( u0_u8_u4_n133 ) , .A2( u0_u8_u4_n146 ) , .A1( u0_u8_u4_n154 ) );
  NAND2_X1 u0_u8_u4_U49 (.A1( u0_u8_u4_n103 ) , .ZN( u0_u8_u4_n154 ) , .A2( u0_u8_u4_n98 ) );
  NOR4_X1 u0_u8_u4_U5 (.A4( u0_u8_u4_n106 ) , .A3( u0_u8_u4_n107 ) , .A2( u0_u8_u4_n108 ) , .A1( u0_u8_u4_n109 ) , .ZN( u0_u8_u4_n110 ) );
  NAND2_X1 u0_u8_u4_U50 (.A1( u0_u8_u4_n101 ) , .ZN( u0_u8_u4_n158 ) , .A2( u0_u8_u4_n99 ) );
  AOI21_X1 u0_u8_u4_U51 (.ZN( u0_u8_u4_n127 ) , .A( u0_u8_u4_n136 ) , .B2( u0_u8_u4_n150 ) , .B1( u0_u8_u4_n180 ) );
  INV_X1 u0_u8_u4_U52 (.A( u0_u8_u4_n160 ) , .ZN( u0_u8_u4_n180 ) );
  NAND2_X1 u0_u8_u4_U53 (.A2( u0_u8_u4_n104 ) , .A1( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n146 ) );
  NAND2_X1 u0_u8_u4_U54 (.A2( u0_u8_u4_n101 ) , .A1( u0_u8_u4_n102 ) , .ZN( u0_u8_u4_n160 ) );
  NAND2_X1 u0_u8_u4_U55 (.ZN( u0_u8_u4_n134 ) , .A1( u0_u8_u4_n98 ) , .A2( u0_u8_u4_n99 ) );
  NAND2_X1 u0_u8_u4_U56 (.A1( u0_u8_u4_n103 ) , .A2( u0_u8_u4_n104 ) , .ZN( u0_u8_u4_n143 ) );
  NAND2_X1 u0_u8_u4_U57 (.A2( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n145 ) , .A1( u0_u8_u4_n98 ) );
  NAND2_X1 u0_u8_u4_U58 (.A1( u0_u8_u4_n100 ) , .A2( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n120 ) );
  NAND2_X1 u0_u8_u4_U59 (.A1( u0_u8_u4_n102 ) , .A2( u0_u8_u4_n104 ) , .ZN( u0_u8_u4_n148 ) );
  AOI21_X1 u0_u8_u4_U6 (.ZN( u0_u8_u4_n106 ) , .B2( u0_u8_u4_n146 ) , .B1( u0_u8_u4_n158 ) , .A( u0_u8_u4_n170 ) );
  NAND2_X1 u0_u8_u4_U60 (.A2( u0_u8_u4_n100 ) , .A1( u0_u8_u4_n103 ) , .ZN( u0_u8_u4_n157 ) );
  INV_X1 u0_u8_u4_U61 (.A( u0_u8_u4_n150 ) , .ZN( u0_u8_u4_n173 ) );
  INV_X1 u0_u8_u4_U62 (.A( u0_u8_u4_n152 ) , .ZN( u0_u8_u4_n171 ) );
  NAND2_X1 u0_u8_u4_U63 (.A1( u0_u8_u4_n100 ) , .ZN( u0_u8_u4_n118 ) , .A2( u0_u8_u4_n99 ) );
  NAND2_X1 u0_u8_u4_U64 (.A2( u0_u8_u4_n100 ) , .A1( u0_u8_u4_n102 ) , .ZN( u0_u8_u4_n144 ) );
  NAND2_X1 u0_u8_u4_U65 (.A2( u0_u8_u4_n101 ) , .A1( u0_u8_u4_n105 ) , .ZN( u0_u8_u4_n96 ) );
  INV_X1 u0_u8_u4_U66 (.A( u0_u8_u4_n128 ) , .ZN( u0_u8_u4_n174 ) );
  NAND2_X1 u0_u8_u4_U67 (.A2( u0_u8_u4_n102 ) , .ZN( u0_u8_u4_n119 ) , .A1( u0_u8_u4_n98 ) );
  NAND2_X1 u0_u8_u4_U68 (.A2( u0_u8_u4_n101 ) , .A1( u0_u8_u4_n103 ) , .ZN( u0_u8_u4_n147 ) );
  NAND2_X1 u0_u8_u4_U69 (.A2( u0_u8_u4_n104 ) , .ZN( u0_u8_u4_n113 ) , .A1( u0_u8_u4_n99 ) );
  AOI21_X1 u0_u8_u4_U7 (.ZN( u0_u8_u4_n108 ) , .B2( u0_u8_u4_n134 ) , .B1( u0_u8_u4_n155 ) , .A( u0_u8_u4_n156 ) );
  NOR2_X1 u0_u8_u4_U70 (.A2( u0_u8_X_28 ) , .ZN( u0_u8_u4_n150 ) , .A1( u0_u8_u4_n168 ) );
  NOR2_X1 u0_u8_u4_U71 (.A2( u0_u8_X_29 ) , .ZN( u0_u8_u4_n152 ) , .A1( u0_u8_u4_n169 ) );
  NOR2_X1 u0_u8_u4_U72 (.A2( u0_u8_X_30 ) , .ZN( u0_u8_u4_n105 ) , .A1( u0_u8_u4_n176 ) );
  NOR2_X1 u0_u8_u4_U73 (.A2( u0_u8_X_26 ) , .ZN( u0_u8_u4_n100 ) , .A1( u0_u8_u4_n177 ) );
  NOR2_X1 u0_u8_u4_U74 (.A2( u0_u8_X_28 ) , .A1( u0_u8_X_29 ) , .ZN( u0_u8_u4_n128 ) );
  NOR2_X1 u0_u8_u4_U75 (.A2( u0_u8_X_27 ) , .A1( u0_u8_X_30 ) , .ZN( u0_u8_u4_n102 ) );
  NOR2_X1 u0_u8_u4_U76 (.A2( u0_u8_X_25 ) , .A1( u0_u8_X_26 ) , .ZN( u0_u8_u4_n98 ) );
  AND2_X1 u0_u8_u4_U77 (.A2( u0_u8_X_25 ) , .A1( u0_u8_X_26 ) , .ZN( u0_u8_u4_n104 ) );
  AND2_X1 u0_u8_u4_U78 (.A1( u0_u8_X_30 ) , .A2( u0_u8_u4_n176 ) , .ZN( u0_u8_u4_n99 ) );
  AND2_X1 u0_u8_u4_U79 (.A1( u0_u8_X_26 ) , .ZN( u0_u8_u4_n101 ) , .A2( u0_u8_u4_n177 ) );
  AOI21_X1 u0_u8_u4_U8 (.ZN( u0_u8_u4_n109 ) , .A( u0_u8_u4_n153 ) , .B1( u0_u8_u4_n159 ) , .B2( u0_u8_u4_n184 ) );
  AND2_X1 u0_u8_u4_U80 (.A1( u0_u8_X_27 ) , .A2( u0_u8_X_30 ) , .ZN( u0_u8_u4_n103 ) );
  INV_X1 u0_u8_u4_U81 (.A( u0_u8_X_28 ) , .ZN( u0_u8_u4_n169 ) );
  INV_X1 u0_u8_u4_U82 (.A( u0_u8_X_29 ) , .ZN( u0_u8_u4_n168 ) );
  INV_X1 u0_u8_u4_U83 (.A( u0_u8_X_25 ) , .ZN( u0_u8_u4_n177 ) );
  INV_X1 u0_u8_u4_U84 (.A( u0_u8_X_27 ) , .ZN( u0_u8_u4_n176 ) );
  NAND4_X1 u0_u8_u4_U85 (.ZN( u0_out8_25 ) , .A4( u0_u8_u4_n139 ) , .A3( u0_u8_u4_n140 ) , .A2( u0_u8_u4_n141 ) , .A1( u0_u8_u4_n142 ) );
  OAI21_X1 u0_u8_u4_U86 (.B2( u0_u8_u4_n131 ) , .ZN( u0_u8_u4_n141 ) , .A( u0_u8_u4_n175 ) , .B1( u0_u8_u4_n183 ) );
  OAI21_X1 u0_u8_u4_U87 (.A( u0_u8_u4_n128 ) , .B2( u0_u8_u4_n129 ) , .B1( u0_u8_u4_n130 ) , .ZN( u0_u8_u4_n142 ) );
  NAND4_X1 u0_u8_u4_U88 (.ZN( u0_out8_14 ) , .A4( u0_u8_u4_n124 ) , .A3( u0_u8_u4_n125 ) , .A2( u0_u8_u4_n126 ) , .A1( u0_u8_u4_n127 ) );
  AOI22_X1 u0_u8_u4_U89 (.B2( u0_u8_u4_n117 ) , .ZN( u0_u8_u4_n126 ) , .A1( u0_u8_u4_n129 ) , .B1( u0_u8_u4_n152 ) , .A2( u0_u8_u4_n175 ) );
  AOI211_X1 u0_u8_u4_U9 (.B( u0_u8_u4_n136 ) , .A( u0_u8_u4_n137 ) , .C2( u0_u8_u4_n138 ) , .ZN( u0_u8_u4_n139 ) , .C1( u0_u8_u4_n182 ) );
  AOI22_X1 u0_u8_u4_U90 (.ZN( u0_u8_u4_n125 ) , .B2( u0_u8_u4_n131 ) , .A2( u0_u8_u4_n132 ) , .B1( u0_u8_u4_n138 ) , .A1( u0_u8_u4_n178 ) );
  NAND4_X1 u0_u8_u4_U91 (.ZN( u0_out8_8 ) , .A4( u0_u8_u4_n110 ) , .A3( u0_u8_u4_n111 ) , .A2( u0_u8_u4_n112 ) , .A1( u0_u8_u4_n186 ) );
  NAND2_X1 u0_u8_u4_U92 (.ZN( u0_u8_u4_n112 ) , .A2( u0_u8_u4_n130 ) , .A1( u0_u8_u4_n150 ) );
  AOI22_X1 u0_u8_u4_U93 (.ZN( u0_u8_u4_n111 ) , .B2( u0_u8_u4_n132 ) , .A1( u0_u8_u4_n152 ) , .B1( u0_u8_u4_n178 ) , .A2( u0_u8_u4_n97 ) );
  AOI22_X1 u0_u8_u4_U94 (.B2( u0_u8_u4_n149 ) , .B1( u0_u8_u4_n150 ) , .A2( u0_u8_u4_n151 ) , .A1( u0_u8_u4_n152 ) , .ZN( u0_u8_u4_n167 ) );
  NOR4_X1 u0_u8_u4_U95 (.A4( u0_u8_u4_n162 ) , .A3( u0_u8_u4_n163 ) , .A2( u0_u8_u4_n164 ) , .A1( u0_u8_u4_n165 ) , .ZN( u0_u8_u4_n166 ) );
  NAND3_X1 u0_u8_u4_U96 (.ZN( u0_out8_3 ) , .A3( u0_u8_u4_n166 ) , .A1( u0_u8_u4_n167 ) , .A2( u0_u8_u4_n186 ) );
  NAND3_X1 u0_u8_u4_U97 (.A3( u0_u8_u4_n146 ) , .A2( u0_u8_u4_n147 ) , .A1( u0_u8_u4_n148 ) , .ZN( u0_u8_u4_n149 ) );
  NAND3_X1 u0_u8_u4_U98 (.A3( u0_u8_u4_n143 ) , .A2( u0_u8_u4_n144 ) , .A1( u0_u8_u4_n145 ) , .ZN( u0_u8_u4_n151 ) );
  NAND3_X1 u0_u8_u4_U99 (.A3( u0_u8_u4_n121 ) , .ZN( u0_u8_u4_n122 ) , .A2( u0_u8_u4_n144 ) , .A1( u0_u8_u4_n154 ) );
  AND3_X1 u0_u8_u7_U10 (.A3( u0_u8_u7_n110 ) , .A2( u0_u8_u7_n127 ) , .A1( u0_u8_u7_n132 ) , .ZN( u0_u8_u7_n92 ) );
  OAI21_X1 u0_u8_u7_U11 (.A( u0_u8_u7_n161 ) , .B1( u0_u8_u7_n168 ) , .B2( u0_u8_u7_n173 ) , .ZN( u0_u8_u7_n91 ) );
  AOI211_X1 u0_u8_u7_U12 (.A( u0_u8_u7_n117 ) , .ZN( u0_u8_u7_n118 ) , .C2( u0_u8_u7_n126 ) , .C1( u0_u8_u7_n177 ) , .B( u0_u8_u7_n180 ) );
  OAI22_X1 u0_u8_u7_U13 (.B1( u0_u8_u7_n115 ) , .ZN( u0_u8_u7_n117 ) , .A2( u0_u8_u7_n133 ) , .A1( u0_u8_u7_n137 ) , .B2( u0_u8_u7_n162 ) );
  INV_X1 u0_u8_u7_U14 (.A( u0_u8_u7_n116 ) , .ZN( u0_u8_u7_n180 ) );
  NOR3_X1 u0_u8_u7_U15 (.ZN( u0_u8_u7_n115 ) , .A3( u0_u8_u7_n145 ) , .A2( u0_u8_u7_n168 ) , .A1( u0_u8_u7_n169 ) );
  OAI211_X1 u0_u8_u7_U16 (.B( u0_u8_u7_n122 ) , .A( u0_u8_u7_n123 ) , .C2( u0_u8_u7_n124 ) , .ZN( u0_u8_u7_n154 ) , .C1( u0_u8_u7_n162 ) );
  AOI222_X1 u0_u8_u7_U17 (.ZN( u0_u8_u7_n122 ) , .C2( u0_u8_u7_n126 ) , .C1( u0_u8_u7_n145 ) , .B1( u0_u8_u7_n161 ) , .A2( u0_u8_u7_n165 ) , .B2( u0_u8_u7_n170 ) , .A1( u0_u8_u7_n176 ) );
  INV_X1 u0_u8_u7_U18 (.A( u0_u8_u7_n133 ) , .ZN( u0_u8_u7_n176 ) );
  NOR3_X1 u0_u8_u7_U19 (.A2( u0_u8_u7_n134 ) , .A1( u0_u8_u7_n135 ) , .ZN( u0_u8_u7_n136 ) , .A3( u0_u8_u7_n171 ) );
  NOR2_X1 u0_u8_u7_U20 (.A1( u0_u8_u7_n130 ) , .A2( u0_u8_u7_n134 ) , .ZN( u0_u8_u7_n153 ) );
  INV_X1 u0_u8_u7_U21 (.A( u0_u8_u7_n101 ) , .ZN( u0_u8_u7_n165 ) );
  NOR2_X1 u0_u8_u7_U22 (.ZN( u0_u8_u7_n111 ) , .A2( u0_u8_u7_n134 ) , .A1( u0_u8_u7_n169 ) );
  AOI21_X1 u0_u8_u7_U23 (.ZN( u0_u8_u7_n104 ) , .B2( u0_u8_u7_n112 ) , .B1( u0_u8_u7_n127 ) , .A( u0_u8_u7_n164 ) );
  AOI21_X1 u0_u8_u7_U24 (.ZN( u0_u8_u7_n106 ) , .B1( u0_u8_u7_n133 ) , .B2( u0_u8_u7_n146 ) , .A( u0_u8_u7_n162 ) );
  AOI21_X1 u0_u8_u7_U25 (.A( u0_u8_u7_n101 ) , .ZN( u0_u8_u7_n107 ) , .B2( u0_u8_u7_n128 ) , .B1( u0_u8_u7_n175 ) );
  INV_X1 u0_u8_u7_U26 (.A( u0_u8_u7_n138 ) , .ZN( u0_u8_u7_n171 ) );
  INV_X1 u0_u8_u7_U27 (.A( u0_u8_u7_n131 ) , .ZN( u0_u8_u7_n177 ) );
  INV_X1 u0_u8_u7_U28 (.A( u0_u8_u7_n110 ) , .ZN( u0_u8_u7_n174 ) );
  NAND2_X1 u0_u8_u7_U29 (.A1( u0_u8_u7_n129 ) , .A2( u0_u8_u7_n132 ) , .ZN( u0_u8_u7_n149 ) );
  OAI21_X1 u0_u8_u7_U3 (.ZN( u0_u8_u7_n159 ) , .A( u0_u8_u7_n165 ) , .B2( u0_u8_u7_n171 ) , .B1( u0_u8_u7_n174 ) );
  NAND2_X1 u0_u8_u7_U30 (.A1( u0_u8_u7_n113 ) , .A2( u0_u8_u7_n124 ) , .ZN( u0_u8_u7_n130 ) );
  INV_X1 u0_u8_u7_U31 (.A( u0_u8_u7_n112 ) , .ZN( u0_u8_u7_n173 ) );
  INV_X1 u0_u8_u7_U32 (.A( u0_u8_u7_n128 ) , .ZN( u0_u8_u7_n168 ) );
  INV_X1 u0_u8_u7_U33 (.A( u0_u8_u7_n148 ) , .ZN( u0_u8_u7_n169 ) );
  INV_X1 u0_u8_u7_U34 (.A( u0_u8_u7_n127 ) , .ZN( u0_u8_u7_n179 ) );
  NOR2_X1 u0_u8_u7_U35 (.ZN( u0_u8_u7_n101 ) , .A2( u0_u8_u7_n150 ) , .A1( u0_u8_u7_n156 ) );
  AOI211_X1 u0_u8_u7_U36 (.B( u0_u8_u7_n154 ) , .A( u0_u8_u7_n155 ) , .C1( u0_u8_u7_n156 ) , .ZN( u0_u8_u7_n157 ) , .C2( u0_u8_u7_n172 ) );
  INV_X1 u0_u8_u7_U37 (.A( u0_u8_u7_n153 ) , .ZN( u0_u8_u7_n172 ) );
  AOI211_X1 u0_u8_u7_U38 (.B( u0_u8_u7_n139 ) , .A( u0_u8_u7_n140 ) , .C2( u0_u8_u7_n141 ) , .ZN( u0_u8_u7_n142 ) , .C1( u0_u8_u7_n156 ) );
  NAND4_X1 u0_u8_u7_U39 (.A3( u0_u8_u7_n127 ) , .A2( u0_u8_u7_n128 ) , .A1( u0_u8_u7_n129 ) , .ZN( u0_u8_u7_n141 ) , .A4( u0_u8_u7_n147 ) );
  INV_X1 u0_u8_u7_U4 (.A( u0_u8_u7_n111 ) , .ZN( u0_u8_u7_n170 ) );
  AOI21_X1 u0_u8_u7_U40 (.A( u0_u8_u7_n137 ) , .B1( u0_u8_u7_n138 ) , .ZN( u0_u8_u7_n139 ) , .B2( u0_u8_u7_n146 ) );
  OAI22_X1 u0_u8_u7_U41 (.B1( u0_u8_u7_n136 ) , .ZN( u0_u8_u7_n140 ) , .A1( u0_u8_u7_n153 ) , .B2( u0_u8_u7_n162 ) , .A2( u0_u8_u7_n164 ) );
  AOI21_X1 u0_u8_u7_U42 (.ZN( u0_u8_u7_n123 ) , .B1( u0_u8_u7_n165 ) , .B2( u0_u8_u7_n177 ) , .A( u0_u8_u7_n97 ) );
  AOI21_X1 u0_u8_u7_U43 (.B2( u0_u8_u7_n113 ) , .B1( u0_u8_u7_n124 ) , .A( u0_u8_u7_n125 ) , .ZN( u0_u8_u7_n97 ) );
  INV_X1 u0_u8_u7_U44 (.A( u0_u8_u7_n125 ) , .ZN( u0_u8_u7_n161 ) );
  INV_X1 u0_u8_u7_U45 (.A( u0_u8_u7_n152 ) , .ZN( u0_u8_u7_n162 ) );
  AOI22_X1 u0_u8_u7_U46 (.A2( u0_u8_u7_n114 ) , .ZN( u0_u8_u7_n119 ) , .B1( u0_u8_u7_n130 ) , .A1( u0_u8_u7_n156 ) , .B2( u0_u8_u7_n165 ) );
  NAND2_X1 u0_u8_u7_U47 (.A2( u0_u8_u7_n112 ) , .ZN( u0_u8_u7_n114 ) , .A1( u0_u8_u7_n175 ) );
  AND2_X1 u0_u8_u7_U48 (.ZN( u0_u8_u7_n145 ) , .A2( u0_u8_u7_n98 ) , .A1( u0_u8_u7_n99 ) );
  NOR2_X1 u0_u8_u7_U49 (.ZN( u0_u8_u7_n137 ) , .A1( u0_u8_u7_n150 ) , .A2( u0_u8_u7_n161 ) );
  INV_X1 u0_u8_u7_U5 (.A( u0_u8_u7_n149 ) , .ZN( u0_u8_u7_n175 ) );
  AOI21_X1 u0_u8_u7_U50 (.ZN( u0_u8_u7_n105 ) , .B2( u0_u8_u7_n110 ) , .A( u0_u8_u7_n125 ) , .B1( u0_u8_u7_n147 ) );
  NAND2_X1 u0_u8_u7_U51 (.ZN( u0_u8_u7_n146 ) , .A1( u0_u8_u7_n95 ) , .A2( u0_u8_u7_n98 ) );
  NAND2_X1 u0_u8_u7_U52 (.A2( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n147 ) , .A1( u0_u8_u7_n93 ) );
  NAND2_X1 u0_u8_u7_U53 (.A1( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n127 ) , .A2( u0_u8_u7_n99 ) );
  OR2_X1 u0_u8_u7_U54 (.ZN( u0_u8_u7_n126 ) , .A2( u0_u8_u7_n152 ) , .A1( u0_u8_u7_n156 ) );
  NAND2_X1 u0_u8_u7_U55 (.A2( u0_u8_u7_n102 ) , .A1( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n133 ) );
  NAND2_X1 u0_u8_u7_U56 (.ZN( u0_u8_u7_n112 ) , .A2( u0_u8_u7_n96 ) , .A1( u0_u8_u7_n99 ) );
  NAND2_X1 u0_u8_u7_U57 (.A2( u0_u8_u7_n102 ) , .ZN( u0_u8_u7_n128 ) , .A1( u0_u8_u7_n98 ) );
  NAND2_X1 u0_u8_u7_U58 (.A1( u0_u8_u7_n100 ) , .ZN( u0_u8_u7_n113 ) , .A2( u0_u8_u7_n93 ) );
  NAND2_X1 u0_u8_u7_U59 (.A2( u0_u8_u7_n102 ) , .ZN( u0_u8_u7_n124 ) , .A1( u0_u8_u7_n96 ) );
  INV_X1 u0_u8_u7_U6 (.A( u0_u8_u7_n154 ) , .ZN( u0_u8_u7_n178 ) );
  NAND2_X1 u0_u8_u7_U60 (.ZN( u0_u8_u7_n110 ) , .A1( u0_u8_u7_n95 ) , .A2( u0_u8_u7_n96 ) );
  INV_X1 u0_u8_u7_U61 (.A( u0_u8_u7_n150 ) , .ZN( u0_u8_u7_n164 ) );
  AND2_X1 u0_u8_u7_U62 (.ZN( u0_u8_u7_n134 ) , .A1( u0_u8_u7_n93 ) , .A2( u0_u8_u7_n98 ) );
  NAND2_X1 u0_u8_u7_U63 (.A1( u0_u8_u7_n100 ) , .A2( u0_u8_u7_n102 ) , .ZN( u0_u8_u7_n129 ) );
  NAND2_X1 u0_u8_u7_U64 (.A2( u0_u8_u7_n103 ) , .ZN( u0_u8_u7_n131 ) , .A1( u0_u8_u7_n95 ) );
  NAND2_X1 u0_u8_u7_U65 (.A1( u0_u8_u7_n100 ) , .ZN( u0_u8_u7_n138 ) , .A2( u0_u8_u7_n99 ) );
  NAND2_X1 u0_u8_u7_U66 (.ZN( u0_u8_u7_n132 ) , .A1( u0_u8_u7_n93 ) , .A2( u0_u8_u7_n96 ) );
  NAND2_X1 u0_u8_u7_U67 (.A1( u0_u8_u7_n100 ) , .ZN( u0_u8_u7_n148 ) , .A2( u0_u8_u7_n95 ) );
  NOR2_X1 u0_u8_u7_U68 (.A2( u0_u8_X_47 ) , .ZN( u0_u8_u7_n150 ) , .A1( u0_u8_u7_n163 ) );
  NOR2_X1 u0_u8_u7_U69 (.A2( u0_u8_X_43 ) , .A1( u0_u8_X_44 ) , .ZN( u0_u8_u7_n103 ) );
  AOI211_X1 u0_u8_u7_U7 (.ZN( u0_u8_u7_n116 ) , .A( u0_u8_u7_n155 ) , .C1( u0_u8_u7_n161 ) , .C2( u0_u8_u7_n171 ) , .B( u0_u8_u7_n94 ) );
  NOR2_X1 u0_u8_u7_U70 (.A2( u0_u8_X_48 ) , .A1( u0_u8_u7_n166 ) , .ZN( u0_u8_u7_n95 ) );
  NOR2_X1 u0_u8_u7_U71 (.A2( u0_u8_X_45 ) , .A1( u0_u8_X_48 ) , .ZN( u0_u8_u7_n99 ) );
  NOR2_X1 u0_u8_u7_U72 (.A2( u0_u8_X_44 ) , .A1( u0_u8_u7_n167 ) , .ZN( u0_u8_u7_n98 ) );
  NOR2_X1 u0_u8_u7_U73 (.A2( u0_u8_X_46 ) , .A1( u0_u8_X_47 ) , .ZN( u0_u8_u7_n152 ) );
  AND2_X1 u0_u8_u7_U74 (.A1( u0_u8_X_47 ) , .ZN( u0_u8_u7_n156 ) , .A2( u0_u8_u7_n163 ) );
  NAND2_X1 u0_u8_u7_U75 (.A2( u0_u8_X_46 ) , .A1( u0_u8_X_47 ) , .ZN( u0_u8_u7_n125 ) );
  AND2_X1 u0_u8_u7_U76 (.A2( u0_u8_X_45 ) , .A1( u0_u8_X_48 ) , .ZN( u0_u8_u7_n102 ) );
  AND2_X1 u0_u8_u7_U77 (.A2( u0_u8_X_43 ) , .A1( u0_u8_X_44 ) , .ZN( u0_u8_u7_n96 ) );
  AND2_X1 u0_u8_u7_U78 (.A1( u0_u8_X_44 ) , .ZN( u0_u8_u7_n100 ) , .A2( u0_u8_u7_n167 ) );
  AND2_X1 u0_u8_u7_U79 (.A1( u0_u8_X_48 ) , .A2( u0_u8_u7_n166 ) , .ZN( u0_u8_u7_n93 ) );
  OAI222_X1 u0_u8_u7_U8 (.C2( u0_u8_u7_n101 ) , .B2( u0_u8_u7_n111 ) , .A1( u0_u8_u7_n113 ) , .C1( u0_u8_u7_n146 ) , .A2( u0_u8_u7_n162 ) , .B1( u0_u8_u7_n164 ) , .ZN( u0_u8_u7_n94 ) );
  INV_X1 u0_u8_u7_U80 (.A( u0_u8_X_46 ) , .ZN( u0_u8_u7_n163 ) );
  INV_X1 u0_u8_u7_U81 (.A( u0_u8_X_43 ) , .ZN( u0_u8_u7_n167 ) );
  INV_X1 u0_u8_u7_U82 (.A( u0_u8_X_45 ) , .ZN( u0_u8_u7_n166 ) );
  NAND4_X1 u0_u8_u7_U83 (.ZN( u0_out8_27 ) , .A4( u0_u8_u7_n118 ) , .A3( u0_u8_u7_n119 ) , .A2( u0_u8_u7_n120 ) , .A1( u0_u8_u7_n121 ) );
  OAI21_X1 u0_u8_u7_U84 (.ZN( u0_u8_u7_n121 ) , .B2( u0_u8_u7_n145 ) , .A( u0_u8_u7_n150 ) , .B1( u0_u8_u7_n174 ) );
  OAI21_X1 u0_u8_u7_U85 (.ZN( u0_u8_u7_n120 ) , .A( u0_u8_u7_n161 ) , .B2( u0_u8_u7_n170 ) , .B1( u0_u8_u7_n179 ) );
  NAND4_X1 u0_u8_u7_U86 (.ZN( u0_out8_15 ) , .A4( u0_u8_u7_n142 ) , .A3( u0_u8_u7_n143 ) , .A2( u0_u8_u7_n144 ) , .A1( u0_u8_u7_n178 ) );
  OR2_X1 u0_u8_u7_U87 (.A2( u0_u8_u7_n125 ) , .A1( u0_u8_u7_n129 ) , .ZN( u0_u8_u7_n144 ) );
  AOI22_X1 u0_u8_u7_U88 (.A2( u0_u8_u7_n126 ) , .ZN( u0_u8_u7_n143 ) , .B2( u0_u8_u7_n165 ) , .B1( u0_u8_u7_n173 ) , .A1( u0_u8_u7_n174 ) );
  NAND4_X1 u0_u8_u7_U89 (.ZN( u0_out8_5 ) , .A4( u0_u8_u7_n108 ) , .A3( u0_u8_u7_n109 ) , .A1( u0_u8_u7_n116 ) , .A2( u0_u8_u7_n123 ) );
  OAI221_X1 u0_u8_u7_U9 (.C1( u0_u8_u7_n101 ) , .C2( u0_u8_u7_n147 ) , .ZN( u0_u8_u7_n155 ) , .B2( u0_u8_u7_n162 ) , .A( u0_u8_u7_n91 ) , .B1( u0_u8_u7_n92 ) );
  AOI22_X1 u0_u8_u7_U90 (.ZN( u0_u8_u7_n109 ) , .A2( u0_u8_u7_n126 ) , .B2( u0_u8_u7_n145 ) , .B1( u0_u8_u7_n156 ) , .A1( u0_u8_u7_n171 ) );
  NOR4_X1 u0_u8_u7_U91 (.A4( u0_u8_u7_n104 ) , .A3( u0_u8_u7_n105 ) , .A2( u0_u8_u7_n106 ) , .A1( u0_u8_u7_n107 ) , .ZN( u0_u8_u7_n108 ) );
  NAND4_X1 u0_u8_u7_U92 (.ZN( u0_out8_21 ) , .A4( u0_u8_u7_n157 ) , .A3( u0_u8_u7_n158 ) , .A2( u0_u8_u7_n159 ) , .A1( u0_u8_u7_n160 ) );
  OAI21_X1 u0_u8_u7_U93 (.B1( u0_u8_u7_n145 ) , .ZN( u0_u8_u7_n160 ) , .A( u0_u8_u7_n161 ) , .B2( u0_u8_u7_n177 ) );
  AOI22_X1 u0_u8_u7_U94 (.B2( u0_u8_u7_n149 ) , .B1( u0_u8_u7_n150 ) , .A2( u0_u8_u7_n151 ) , .A1( u0_u8_u7_n152 ) , .ZN( u0_u8_u7_n158 ) );
  NAND3_X1 u0_u8_u7_U95 (.A3( u0_u8_u7_n146 ) , .A2( u0_u8_u7_n147 ) , .A1( u0_u8_u7_n148 ) , .ZN( u0_u8_u7_n151 ) );
  NAND3_X1 u0_u8_u7_U96 (.A3( u0_u8_u7_n131 ) , .A2( u0_u8_u7_n132 ) , .A1( u0_u8_u7_n133 ) , .ZN( u0_u8_u7_n135 ) );
  XOR2_X1 u0_u9_U1 (.B( u0_K10_9 ) , .A( u0_R8_6 ) , .Z( u0_u9_X_9 ) );
  XOR2_X1 u0_u9_U2 (.B( u0_K10_8 ) , .A( u0_R8_5 ) , .Z( u0_u9_X_8 ) );
  XOR2_X1 u0_u9_U3 (.B( u0_K10_7 ) , .A( u0_R8_4 ) , .Z( u0_u9_X_7 ) );
  XOR2_X1 u0_u9_U33 (.B( u0_K10_24 ) , .A( u0_R8_17 ) , .Z( u0_u9_X_24 ) );
  XOR2_X1 u0_u9_U34 (.B( u0_K10_23 ) , .A( u0_R8_16 ) , .Z( u0_u9_X_23 ) );
  XOR2_X1 u0_u9_U35 (.B( u0_K10_22 ) , .A( u0_R8_15 ) , .Z( u0_u9_X_22 ) );
  XOR2_X1 u0_u9_U36 (.B( u0_K10_21 ) , .A( u0_R8_14 ) , .Z( u0_u9_X_21 ) );
  XOR2_X1 u0_u9_U37 (.B( u0_K10_20 ) , .A( u0_R8_13 ) , .Z( u0_u9_X_20 ) );
  XOR2_X1 u0_u9_U39 (.B( u0_K10_19 ) , .A( u0_R8_12 ) , .Z( u0_u9_X_19 ) );
  XOR2_X1 u0_u9_U40 (.B( u0_K10_18 ) , .A( u0_R8_13 ) , .Z( u0_u9_X_18 ) );
  XOR2_X1 u0_u9_U41 (.B( u0_K10_17 ) , .A( u0_R8_12 ) , .Z( u0_u9_X_17 ) );
  XOR2_X1 u0_u9_U42 (.B( u0_K10_16 ) , .A( u0_R8_11 ) , .Z( u0_u9_X_16 ) );
  XOR2_X1 u0_u9_U43 (.B( u0_K10_15 ) , .A( u0_R8_10 ) , .Z( u0_u9_X_15 ) );
  XOR2_X1 u0_u9_U44 (.B( u0_K10_14 ) , .A( u0_R8_9 ) , .Z( u0_u9_X_14 ) );
  XOR2_X1 u0_u9_U45 (.B( u0_K10_13 ) , .A( u0_R8_8 ) , .Z( u0_u9_X_13 ) );
  XOR2_X1 u0_u9_U46 (.B( u0_K10_12 ) , .A( u0_R8_9 ) , .Z( u0_u9_X_12 ) );
  XOR2_X1 u0_u9_U47 (.B( u0_K10_11 ) , .A( u0_R8_8 ) , .Z( u0_u9_X_11 ) );
  XOR2_X1 u0_u9_U48 (.B( u0_K10_10 ) , .A( u0_R8_7 ) , .Z( u0_u9_X_10 ) );
  NOR2_X1 u0_u9_u1_U10 (.A1( u0_u9_u1_n112 ) , .A2( u0_u9_u1_n116 ) , .ZN( u0_u9_u1_n118 ) );
  NAND3_X1 u0_u9_u1_U100 (.ZN( u0_u9_u1_n113 ) , .A1( u0_u9_u1_n120 ) , .A3( u0_u9_u1_n133 ) , .A2( u0_u9_u1_n155 ) );
  OAI21_X1 u0_u9_u1_U11 (.ZN( u0_u9_u1_n101 ) , .B1( u0_u9_u1_n141 ) , .A( u0_u9_u1_n146 ) , .B2( u0_u9_u1_n183 ) );
  AOI21_X1 u0_u9_u1_U12 (.B2( u0_u9_u1_n155 ) , .B1( u0_u9_u1_n156 ) , .ZN( u0_u9_u1_n157 ) , .A( u0_u9_u1_n174 ) );
  NAND2_X1 u0_u9_u1_U13 (.ZN( u0_u9_u1_n140 ) , .A2( u0_u9_u1_n150 ) , .A1( u0_u9_u1_n155 ) );
  NAND2_X1 u0_u9_u1_U14 (.A1( u0_u9_u1_n131 ) , .ZN( u0_u9_u1_n147 ) , .A2( u0_u9_u1_n153 ) );
  INV_X1 u0_u9_u1_U15 (.A( u0_u9_u1_n139 ) , .ZN( u0_u9_u1_n174 ) );
  OR4_X1 u0_u9_u1_U16 (.A4( u0_u9_u1_n106 ) , .A3( u0_u9_u1_n107 ) , .ZN( u0_u9_u1_n108 ) , .A1( u0_u9_u1_n117 ) , .A2( u0_u9_u1_n184 ) );
  AOI21_X1 u0_u9_u1_U17 (.ZN( u0_u9_u1_n106 ) , .A( u0_u9_u1_n112 ) , .B1( u0_u9_u1_n154 ) , .B2( u0_u9_u1_n156 ) );
  AOI21_X1 u0_u9_u1_U18 (.ZN( u0_u9_u1_n107 ) , .B1( u0_u9_u1_n134 ) , .B2( u0_u9_u1_n149 ) , .A( u0_u9_u1_n174 ) );
  INV_X1 u0_u9_u1_U19 (.A( u0_u9_u1_n101 ) , .ZN( u0_u9_u1_n184 ) );
  INV_X1 u0_u9_u1_U20 (.A( u0_u9_u1_n112 ) , .ZN( u0_u9_u1_n171 ) );
  NAND2_X1 u0_u9_u1_U21 (.ZN( u0_u9_u1_n141 ) , .A1( u0_u9_u1_n153 ) , .A2( u0_u9_u1_n156 ) );
  AND2_X1 u0_u9_u1_U22 (.A1( u0_u9_u1_n123 ) , .ZN( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n161 ) );
  NAND2_X1 u0_u9_u1_U23 (.A2( u0_u9_u1_n115 ) , .A1( u0_u9_u1_n116 ) , .ZN( u0_u9_u1_n148 ) );
  NAND2_X1 u0_u9_u1_U24 (.A2( u0_u9_u1_n133 ) , .A1( u0_u9_u1_n135 ) , .ZN( u0_u9_u1_n159 ) );
  NAND2_X1 u0_u9_u1_U25 (.A2( u0_u9_u1_n115 ) , .A1( u0_u9_u1_n120 ) , .ZN( u0_u9_u1_n132 ) );
  INV_X1 u0_u9_u1_U26 (.A( u0_u9_u1_n154 ) , .ZN( u0_u9_u1_n178 ) );
  INV_X1 u0_u9_u1_U27 (.A( u0_u9_u1_n151 ) , .ZN( u0_u9_u1_n183 ) );
  AND2_X1 u0_u9_u1_U28 (.A1( u0_u9_u1_n129 ) , .A2( u0_u9_u1_n133 ) , .ZN( u0_u9_u1_n149 ) );
  INV_X1 u0_u9_u1_U29 (.A( u0_u9_u1_n131 ) , .ZN( u0_u9_u1_n180 ) );
  INV_X1 u0_u9_u1_U3 (.A( u0_u9_u1_n159 ) , .ZN( u0_u9_u1_n182 ) );
  OAI221_X1 u0_u9_u1_U30 (.A( u0_u9_u1_n119 ) , .C2( u0_u9_u1_n129 ) , .ZN( u0_u9_u1_n138 ) , .B2( u0_u9_u1_n152 ) , .C1( u0_u9_u1_n174 ) , .B1( u0_u9_u1_n187 ) );
  INV_X1 u0_u9_u1_U31 (.A( u0_u9_u1_n148 ) , .ZN( u0_u9_u1_n187 ) );
  AOI211_X1 u0_u9_u1_U32 (.B( u0_u9_u1_n117 ) , .A( u0_u9_u1_n118 ) , .ZN( u0_u9_u1_n119 ) , .C2( u0_u9_u1_n146 ) , .C1( u0_u9_u1_n159 ) );
  NOR2_X1 u0_u9_u1_U33 (.A1( u0_u9_u1_n168 ) , .A2( u0_u9_u1_n176 ) , .ZN( u0_u9_u1_n98 ) );
  AOI211_X1 u0_u9_u1_U34 (.B( u0_u9_u1_n162 ) , .A( u0_u9_u1_n163 ) , .C2( u0_u9_u1_n164 ) , .ZN( u0_u9_u1_n165 ) , .C1( u0_u9_u1_n171 ) );
  AOI21_X1 u0_u9_u1_U35 (.A( u0_u9_u1_n160 ) , .B2( u0_u9_u1_n161 ) , .ZN( u0_u9_u1_n162 ) , .B1( u0_u9_u1_n182 ) );
  OR2_X1 u0_u9_u1_U36 (.A2( u0_u9_u1_n157 ) , .A1( u0_u9_u1_n158 ) , .ZN( u0_u9_u1_n163 ) );
  NAND2_X1 u0_u9_u1_U37 (.A1( u0_u9_u1_n128 ) , .ZN( u0_u9_u1_n146 ) , .A2( u0_u9_u1_n160 ) );
  NAND2_X1 u0_u9_u1_U38 (.A2( u0_u9_u1_n112 ) , .ZN( u0_u9_u1_n139 ) , .A1( u0_u9_u1_n152 ) );
  NAND2_X1 u0_u9_u1_U39 (.A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n156 ) , .A2( u0_u9_u1_n99 ) );
  AOI221_X1 u0_u9_u1_U4 (.A( u0_u9_u1_n138 ) , .C2( u0_u9_u1_n139 ) , .C1( u0_u9_u1_n140 ) , .B2( u0_u9_u1_n141 ) , .ZN( u0_u9_u1_n142 ) , .B1( u0_u9_u1_n175 ) );
  AOI221_X1 u0_u9_u1_U40 (.B1( u0_u9_u1_n140 ) , .ZN( u0_u9_u1_n167 ) , .B2( u0_u9_u1_n172 ) , .C2( u0_u9_u1_n175 ) , .C1( u0_u9_u1_n178 ) , .A( u0_u9_u1_n188 ) );
  INV_X1 u0_u9_u1_U41 (.ZN( u0_u9_u1_n188 ) , .A( u0_u9_u1_n97 ) );
  AOI211_X1 u0_u9_u1_U42 (.A( u0_u9_u1_n118 ) , .C1( u0_u9_u1_n132 ) , .C2( u0_u9_u1_n139 ) , .B( u0_u9_u1_n96 ) , .ZN( u0_u9_u1_n97 ) );
  AOI21_X1 u0_u9_u1_U43 (.B2( u0_u9_u1_n121 ) , .B1( u0_u9_u1_n135 ) , .A( u0_u9_u1_n152 ) , .ZN( u0_u9_u1_n96 ) );
  NOR2_X1 u0_u9_u1_U44 (.ZN( u0_u9_u1_n117 ) , .A1( u0_u9_u1_n121 ) , .A2( u0_u9_u1_n160 ) );
  OAI21_X1 u0_u9_u1_U45 (.B2( u0_u9_u1_n123 ) , .ZN( u0_u9_u1_n145 ) , .B1( u0_u9_u1_n160 ) , .A( u0_u9_u1_n185 ) );
  INV_X1 u0_u9_u1_U46 (.A( u0_u9_u1_n122 ) , .ZN( u0_u9_u1_n185 ) );
  AOI21_X1 u0_u9_u1_U47 (.B2( u0_u9_u1_n120 ) , .B1( u0_u9_u1_n121 ) , .ZN( u0_u9_u1_n122 ) , .A( u0_u9_u1_n128 ) );
  AOI21_X1 u0_u9_u1_U48 (.A( u0_u9_u1_n128 ) , .B2( u0_u9_u1_n129 ) , .ZN( u0_u9_u1_n130 ) , .B1( u0_u9_u1_n150 ) );
  NAND2_X1 u0_u9_u1_U49 (.ZN( u0_u9_u1_n112 ) , .A1( u0_u9_u1_n169 ) , .A2( u0_u9_u1_n170 ) );
  AOI211_X1 u0_u9_u1_U5 (.ZN( u0_u9_u1_n124 ) , .A( u0_u9_u1_n138 ) , .C2( u0_u9_u1_n139 ) , .B( u0_u9_u1_n145 ) , .C1( u0_u9_u1_n147 ) );
  NAND2_X1 u0_u9_u1_U50 (.ZN( u0_u9_u1_n129 ) , .A2( u0_u9_u1_n95 ) , .A1( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U51 (.A1( u0_u9_u1_n102 ) , .ZN( u0_u9_u1_n154 ) , .A2( u0_u9_u1_n99 ) );
  NAND2_X1 u0_u9_u1_U52 (.A2( u0_u9_u1_n100 ) , .ZN( u0_u9_u1_n135 ) , .A1( u0_u9_u1_n99 ) );
  AOI21_X1 u0_u9_u1_U53 (.A( u0_u9_u1_n152 ) , .B2( u0_u9_u1_n153 ) , .B1( u0_u9_u1_n154 ) , .ZN( u0_u9_u1_n158 ) );
  INV_X1 u0_u9_u1_U54 (.A( u0_u9_u1_n160 ) , .ZN( u0_u9_u1_n175 ) );
  NAND2_X1 u0_u9_u1_U55 (.A1( u0_u9_u1_n100 ) , .ZN( u0_u9_u1_n116 ) , .A2( u0_u9_u1_n95 ) );
  NAND2_X1 u0_u9_u1_U56 (.A1( u0_u9_u1_n102 ) , .ZN( u0_u9_u1_n131 ) , .A2( u0_u9_u1_n95 ) );
  NAND2_X1 u0_u9_u1_U57 (.A2( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n121 ) , .A1( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U58 (.A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n153 ) , .A2( u0_u9_u1_n98 ) );
  NAND2_X1 u0_u9_u1_U59 (.A2( u0_u9_u1_n104 ) , .A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n133 ) );
  AOI22_X1 u0_u9_u1_U6 (.B2( u0_u9_u1_n136 ) , .A2( u0_u9_u1_n137 ) , .ZN( u0_u9_u1_n143 ) , .A1( u0_u9_u1_n171 ) , .B1( u0_u9_u1_n173 ) );
  NAND2_X1 u0_u9_u1_U60 (.ZN( u0_u9_u1_n150 ) , .A2( u0_u9_u1_n98 ) , .A1( u0_u9_u1_n99 ) );
  NAND2_X1 u0_u9_u1_U61 (.A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n155 ) , .A2( u0_u9_u1_n95 ) );
  OAI21_X1 u0_u9_u1_U62 (.ZN( u0_u9_u1_n109 ) , .B1( u0_u9_u1_n129 ) , .B2( u0_u9_u1_n160 ) , .A( u0_u9_u1_n167 ) );
  NAND2_X1 u0_u9_u1_U63 (.A2( u0_u9_u1_n100 ) , .A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n120 ) );
  NAND2_X1 u0_u9_u1_U64 (.A1( u0_u9_u1_n102 ) , .A2( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n115 ) );
  NAND2_X1 u0_u9_u1_U65 (.A2( u0_u9_u1_n100 ) , .A1( u0_u9_u1_n104 ) , .ZN( u0_u9_u1_n151 ) );
  NAND2_X1 u0_u9_u1_U66 (.A2( u0_u9_u1_n103 ) , .A1( u0_u9_u1_n105 ) , .ZN( u0_u9_u1_n161 ) );
  INV_X1 u0_u9_u1_U67 (.A( u0_u9_u1_n152 ) , .ZN( u0_u9_u1_n173 ) );
  INV_X1 u0_u9_u1_U68 (.A( u0_u9_u1_n128 ) , .ZN( u0_u9_u1_n172 ) );
  NAND2_X1 u0_u9_u1_U69 (.A2( u0_u9_u1_n102 ) , .A1( u0_u9_u1_n103 ) , .ZN( u0_u9_u1_n123 ) );
  INV_X1 u0_u9_u1_U7 (.A( u0_u9_u1_n147 ) , .ZN( u0_u9_u1_n181 ) );
  NOR2_X1 u0_u9_u1_U70 (.A2( u0_u9_X_7 ) , .A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n95 ) );
  NOR2_X1 u0_u9_u1_U71 (.A1( u0_u9_X_12 ) , .A2( u0_u9_X_9 ) , .ZN( u0_u9_u1_n100 ) );
  NOR2_X1 u0_u9_u1_U72 (.A2( u0_u9_X_8 ) , .A1( u0_u9_u1_n177 ) , .ZN( u0_u9_u1_n99 ) );
  NOR2_X1 u0_u9_u1_U73 (.A2( u0_u9_X_12 ) , .ZN( u0_u9_u1_n102 ) , .A1( u0_u9_u1_n176 ) );
  NOR2_X1 u0_u9_u1_U74 (.A2( u0_u9_X_9 ) , .ZN( u0_u9_u1_n105 ) , .A1( u0_u9_u1_n168 ) );
  NAND2_X1 u0_u9_u1_U75 (.A1( u0_u9_X_10 ) , .ZN( u0_u9_u1_n160 ) , .A2( u0_u9_u1_n169 ) );
  NAND2_X1 u0_u9_u1_U76 (.A2( u0_u9_X_10 ) , .A1( u0_u9_X_11 ) , .ZN( u0_u9_u1_n152 ) );
  NAND2_X1 u0_u9_u1_U77 (.A1( u0_u9_X_11 ) , .ZN( u0_u9_u1_n128 ) , .A2( u0_u9_u1_n170 ) );
  AND2_X1 u0_u9_u1_U78 (.A2( u0_u9_X_7 ) , .A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n104 ) );
  AND2_X1 u0_u9_u1_U79 (.A1( u0_u9_X_8 ) , .ZN( u0_u9_u1_n103 ) , .A2( u0_u9_u1_n177 ) );
  AOI22_X1 u0_u9_u1_U8 (.B2( u0_u9_u1_n113 ) , .A2( u0_u9_u1_n114 ) , .ZN( u0_u9_u1_n125 ) , .A1( u0_u9_u1_n171 ) , .B1( u0_u9_u1_n173 ) );
  INV_X1 u0_u9_u1_U80 (.A( u0_u9_X_10 ) , .ZN( u0_u9_u1_n170 ) );
  INV_X1 u0_u9_u1_U81 (.A( u0_u9_X_9 ) , .ZN( u0_u9_u1_n176 ) );
  INV_X1 u0_u9_u1_U82 (.A( u0_u9_X_11 ) , .ZN( u0_u9_u1_n169 ) );
  INV_X1 u0_u9_u1_U83 (.A( u0_u9_X_12 ) , .ZN( u0_u9_u1_n168 ) );
  INV_X1 u0_u9_u1_U84 (.A( u0_u9_X_7 ) , .ZN( u0_u9_u1_n177 ) );
  NAND4_X1 u0_u9_u1_U85 (.ZN( u0_out9_28 ) , .A4( u0_u9_u1_n124 ) , .A3( u0_u9_u1_n125 ) , .A2( u0_u9_u1_n126 ) , .A1( u0_u9_u1_n127 ) );
  OAI21_X1 u0_u9_u1_U86 (.ZN( u0_u9_u1_n127 ) , .B2( u0_u9_u1_n139 ) , .B1( u0_u9_u1_n175 ) , .A( u0_u9_u1_n183 ) );
  OAI21_X1 u0_u9_u1_U87 (.ZN( u0_u9_u1_n126 ) , .B2( u0_u9_u1_n140 ) , .A( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n178 ) );
  NAND4_X1 u0_u9_u1_U88 (.ZN( u0_out9_18 ) , .A4( u0_u9_u1_n165 ) , .A3( u0_u9_u1_n166 ) , .A1( u0_u9_u1_n167 ) , .A2( u0_u9_u1_n186 ) );
  AOI22_X1 u0_u9_u1_U89 (.B2( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n147 ) , .A2( u0_u9_u1_n148 ) , .ZN( u0_u9_u1_n166 ) , .A1( u0_u9_u1_n172 ) );
  NAND2_X1 u0_u9_u1_U9 (.ZN( u0_u9_u1_n114 ) , .A1( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n156 ) );
  INV_X1 u0_u9_u1_U90 (.A( u0_u9_u1_n145 ) , .ZN( u0_u9_u1_n186 ) );
  NAND4_X1 u0_u9_u1_U91 (.ZN( u0_out9_2 ) , .A4( u0_u9_u1_n142 ) , .A3( u0_u9_u1_n143 ) , .A2( u0_u9_u1_n144 ) , .A1( u0_u9_u1_n179 ) );
  OAI21_X1 u0_u9_u1_U92 (.B2( u0_u9_u1_n132 ) , .ZN( u0_u9_u1_n144 ) , .A( u0_u9_u1_n146 ) , .B1( u0_u9_u1_n180 ) );
  INV_X1 u0_u9_u1_U93 (.A( u0_u9_u1_n130 ) , .ZN( u0_u9_u1_n179 ) );
  OR4_X1 u0_u9_u1_U94 (.ZN( u0_out9_13 ) , .A4( u0_u9_u1_n108 ) , .A3( u0_u9_u1_n109 ) , .A2( u0_u9_u1_n110 ) , .A1( u0_u9_u1_n111 ) );
  AOI21_X1 u0_u9_u1_U95 (.ZN( u0_u9_u1_n110 ) , .A( u0_u9_u1_n116 ) , .B1( u0_u9_u1_n152 ) , .B2( u0_u9_u1_n160 ) );
  AOI21_X1 u0_u9_u1_U96 (.ZN( u0_u9_u1_n111 ) , .A( u0_u9_u1_n128 ) , .B2( u0_u9_u1_n131 ) , .B1( u0_u9_u1_n135 ) );
  NAND3_X1 u0_u9_u1_U97 (.A3( u0_u9_u1_n149 ) , .A2( u0_u9_u1_n150 ) , .A1( u0_u9_u1_n151 ) , .ZN( u0_u9_u1_n164 ) );
  NAND3_X1 u0_u9_u1_U98 (.A3( u0_u9_u1_n134 ) , .A2( u0_u9_u1_n135 ) , .ZN( u0_u9_u1_n136 ) , .A1( u0_u9_u1_n151 ) );
  NAND3_X1 u0_u9_u1_U99 (.A1( u0_u9_u1_n133 ) , .ZN( u0_u9_u1_n137 ) , .A2( u0_u9_u1_n154 ) , .A3( u0_u9_u1_n181 ) );
  OAI22_X1 u0_u9_u2_U10 (.B1( u0_u9_u2_n151 ) , .A2( u0_u9_u2_n152 ) , .A1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n160 ) , .B2( u0_u9_u2_n168 ) );
  NAND3_X1 u0_u9_u2_U100 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n98 ) );
  NOR3_X1 u0_u9_u2_U11 (.A1( u0_u9_u2_n150 ) , .ZN( u0_u9_u2_n151 ) , .A3( u0_u9_u2_n175 ) , .A2( u0_u9_u2_n188 ) );
  AOI21_X1 u0_u9_u2_U12 (.B2( u0_u9_u2_n123 ) , .ZN( u0_u9_u2_n125 ) , .A( u0_u9_u2_n171 ) , .B1( u0_u9_u2_n184 ) );
  INV_X1 u0_u9_u2_U13 (.A( u0_u9_u2_n150 ) , .ZN( u0_u9_u2_n184 ) );
  AOI21_X1 u0_u9_u2_U14 (.ZN( u0_u9_u2_n144 ) , .B2( u0_u9_u2_n155 ) , .A( u0_u9_u2_n172 ) , .B1( u0_u9_u2_n185 ) );
  AOI21_X1 u0_u9_u2_U15 (.B2( u0_u9_u2_n143 ) , .ZN( u0_u9_u2_n145 ) , .B1( u0_u9_u2_n152 ) , .A( u0_u9_u2_n171 ) );
  INV_X1 u0_u9_u2_U16 (.A( u0_u9_u2_n156 ) , .ZN( u0_u9_u2_n171 ) );
  INV_X1 u0_u9_u2_U17 (.A( u0_u9_u2_n120 ) , .ZN( u0_u9_u2_n188 ) );
  NAND2_X1 u0_u9_u2_U18 (.A2( u0_u9_u2_n122 ) , .ZN( u0_u9_u2_n150 ) , .A1( u0_u9_u2_n152 ) );
  INV_X1 u0_u9_u2_U19 (.A( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n170 ) );
  INV_X1 u0_u9_u2_U20 (.A( u0_u9_u2_n137 ) , .ZN( u0_u9_u2_n173 ) );
  NAND2_X1 u0_u9_u2_U21 (.A1( u0_u9_u2_n132 ) , .A2( u0_u9_u2_n139 ) , .ZN( u0_u9_u2_n157 ) );
  INV_X1 u0_u9_u2_U22 (.A( u0_u9_u2_n113 ) , .ZN( u0_u9_u2_n178 ) );
  INV_X1 u0_u9_u2_U23 (.A( u0_u9_u2_n139 ) , .ZN( u0_u9_u2_n175 ) );
  INV_X1 u0_u9_u2_U24 (.A( u0_u9_u2_n155 ) , .ZN( u0_u9_u2_n181 ) );
  INV_X1 u0_u9_u2_U25 (.A( u0_u9_u2_n119 ) , .ZN( u0_u9_u2_n177 ) );
  INV_X1 u0_u9_u2_U26 (.A( u0_u9_u2_n116 ) , .ZN( u0_u9_u2_n180 ) );
  INV_X1 u0_u9_u2_U27 (.A( u0_u9_u2_n131 ) , .ZN( u0_u9_u2_n179 ) );
  INV_X1 u0_u9_u2_U28 (.A( u0_u9_u2_n154 ) , .ZN( u0_u9_u2_n176 ) );
  NAND2_X1 u0_u9_u2_U29 (.A2( u0_u9_u2_n116 ) , .A1( u0_u9_u2_n117 ) , .ZN( u0_u9_u2_n118 ) );
  NOR2_X1 u0_u9_u2_U3 (.ZN( u0_u9_u2_n121 ) , .A2( u0_u9_u2_n177 ) , .A1( u0_u9_u2_n180 ) );
  INV_X1 u0_u9_u2_U30 (.A( u0_u9_u2_n132 ) , .ZN( u0_u9_u2_n182 ) );
  INV_X1 u0_u9_u2_U31 (.A( u0_u9_u2_n158 ) , .ZN( u0_u9_u2_n183 ) );
  OAI21_X1 u0_u9_u2_U32 (.A( u0_u9_u2_n156 ) , .B1( u0_u9_u2_n157 ) , .ZN( u0_u9_u2_n158 ) , .B2( u0_u9_u2_n179 ) );
  NOR2_X1 u0_u9_u2_U33 (.ZN( u0_u9_u2_n156 ) , .A1( u0_u9_u2_n166 ) , .A2( u0_u9_u2_n169 ) );
  NOR2_X1 u0_u9_u2_U34 (.A2( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n137 ) , .A1( u0_u9_u2_n140 ) );
  NOR2_X1 u0_u9_u2_U35 (.A2( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n153 ) , .A1( u0_u9_u2_n156 ) );
  AOI211_X1 u0_u9_u2_U36 (.ZN( u0_u9_u2_n130 ) , .C1( u0_u9_u2_n138 ) , .C2( u0_u9_u2_n179 ) , .B( u0_u9_u2_n96 ) , .A( u0_u9_u2_n97 ) );
  OAI22_X1 u0_u9_u2_U37 (.B1( u0_u9_u2_n133 ) , .A2( u0_u9_u2_n137 ) , .A1( u0_u9_u2_n152 ) , .B2( u0_u9_u2_n168 ) , .ZN( u0_u9_u2_n97 ) );
  OAI221_X1 u0_u9_u2_U38 (.B1( u0_u9_u2_n113 ) , .C1( u0_u9_u2_n132 ) , .A( u0_u9_u2_n149 ) , .B2( u0_u9_u2_n171 ) , .C2( u0_u9_u2_n172 ) , .ZN( u0_u9_u2_n96 ) );
  OAI221_X1 u0_u9_u2_U39 (.A( u0_u9_u2_n115 ) , .C2( u0_u9_u2_n123 ) , .B2( u0_u9_u2_n143 ) , .B1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n163 ) , .C1( u0_u9_u2_n168 ) );
  INV_X1 u0_u9_u2_U4 (.A( u0_u9_u2_n134 ) , .ZN( u0_u9_u2_n185 ) );
  OAI21_X1 u0_u9_u2_U40 (.A( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n115 ) , .B1( u0_u9_u2_n176 ) , .B2( u0_u9_u2_n178 ) );
  OAI221_X1 u0_u9_u2_U41 (.A( u0_u9_u2_n135 ) , .B2( u0_u9_u2_n136 ) , .B1( u0_u9_u2_n137 ) , .ZN( u0_u9_u2_n162 ) , .C2( u0_u9_u2_n167 ) , .C1( u0_u9_u2_n185 ) );
  AND3_X1 u0_u9_u2_U42 (.A3( u0_u9_u2_n131 ) , .A2( u0_u9_u2_n132 ) , .A1( u0_u9_u2_n133 ) , .ZN( u0_u9_u2_n136 ) );
  AOI22_X1 u0_u9_u2_U43 (.ZN( u0_u9_u2_n135 ) , .B1( u0_u9_u2_n140 ) , .A1( u0_u9_u2_n156 ) , .B2( u0_u9_u2_n180 ) , .A2( u0_u9_u2_n188 ) );
  AOI21_X1 u0_u9_u2_U44 (.ZN( u0_u9_u2_n149 ) , .B1( u0_u9_u2_n173 ) , .B2( u0_u9_u2_n188 ) , .A( u0_u9_u2_n95 ) );
  AND3_X1 u0_u9_u2_U45 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n156 ) , .ZN( u0_u9_u2_n95 ) );
  OAI21_X1 u0_u9_u2_U46 (.A( u0_u9_u2_n141 ) , .B2( u0_u9_u2_n142 ) , .ZN( u0_u9_u2_n146 ) , .B1( u0_u9_u2_n153 ) );
  OAI21_X1 u0_u9_u2_U47 (.A( u0_u9_u2_n140 ) , .ZN( u0_u9_u2_n141 ) , .B1( u0_u9_u2_n176 ) , .B2( u0_u9_u2_n177 ) );
  NOR3_X1 u0_u9_u2_U48 (.ZN( u0_u9_u2_n142 ) , .A3( u0_u9_u2_n175 ) , .A2( u0_u9_u2_n178 ) , .A1( u0_u9_u2_n181 ) );
  OAI21_X1 u0_u9_u2_U49 (.A( u0_u9_u2_n101 ) , .B2( u0_u9_u2_n121 ) , .B1( u0_u9_u2_n153 ) , .ZN( u0_u9_u2_n164 ) );
  NOR4_X1 u0_u9_u2_U5 (.A4( u0_u9_u2_n124 ) , .A3( u0_u9_u2_n125 ) , .A2( u0_u9_u2_n126 ) , .A1( u0_u9_u2_n127 ) , .ZN( u0_u9_u2_n128 ) );
  NAND2_X1 u0_u9_u2_U50 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n155 ) );
  NAND2_X1 u0_u9_u2_U51 (.A2( u0_u9_u2_n105 ) , .A1( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n143 ) );
  NAND2_X1 u0_u9_u2_U52 (.A1( u0_u9_u2_n104 ) , .A2( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n152 ) );
  NAND2_X1 u0_u9_u2_U53 (.A1( u0_u9_u2_n100 ) , .A2( u0_u9_u2_n105 ) , .ZN( u0_u9_u2_n132 ) );
  INV_X1 u0_u9_u2_U54 (.A( u0_u9_u2_n140 ) , .ZN( u0_u9_u2_n168 ) );
  INV_X1 u0_u9_u2_U55 (.A( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n167 ) );
  NAND2_X1 u0_u9_u2_U56 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n113 ) );
  NAND2_X1 u0_u9_u2_U57 (.A1( u0_u9_u2_n106 ) , .A2( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n131 ) );
  NAND2_X1 u0_u9_u2_U58 (.A1( u0_u9_u2_n103 ) , .A2( u0_u9_u2_n107 ) , .ZN( u0_u9_u2_n139 ) );
  NAND2_X1 u0_u9_u2_U59 (.A1( u0_u9_u2_n103 ) , .A2( u0_u9_u2_n105 ) , .ZN( u0_u9_u2_n133 ) );
  AOI21_X1 u0_u9_u2_U6 (.B2( u0_u9_u2_n119 ) , .ZN( u0_u9_u2_n127 ) , .A( u0_u9_u2_n137 ) , .B1( u0_u9_u2_n155 ) );
  NAND2_X1 u0_u9_u2_U60 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n103 ) , .ZN( u0_u9_u2_n154 ) );
  NAND2_X1 u0_u9_u2_U61 (.A2( u0_u9_u2_n103 ) , .A1( u0_u9_u2_n104 ) , .ZN( u0_u9_u2_n119 ) );
  NAND2_X1 u0_u9_u2_U62 (.A2( u0_u9_u2_n107 ) , .A1( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n123 ) );
  NAND2_X1 u0_u9_u2_U63 (.A1( u0_u9_u2_n104 ) , .A2( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n122 ) );
  INV_X1 u0_u9_u2_U64 (.A( u0_u9_u2_n114 ) , .ZN( u0_u9_u2_n172 ) );
  NAND2_X1 u0_u9_u2_U65 (.A2( u0_u9_u2_n100 ) , .A1( u0_u9_u2_n102 ) , .ZN( u0_u9_u2_n116 ) );
  NAND2_X1 u0_u9_u2_U66 (.A1( u0_u9_u2_n102 ) , .A2( u0_u9_u2_n108 ) , .ZN( u0_u9_u2_n120 ) );
  NAND2_X1 u0_u9_u2_U67 (.A2( u0_u9_u2_n105 ) , .A1( u0_u9_u2_n106 ) , .ZN( u0_u9_u2_n117 ) );
  INV_X1 u0_u9_u2_U68 (.ZN( u0_u9_u2_n187 ) , .A( u0_u9_u2_n99 ) );
  OAI21_X1 u0_u9_u2_U69 (.B1( u0_u9_u2_n137 ) , .B2( u0_u9_u2_n143 ) , .A( u0_u9_u2_n98 ) , .ZN( u0_u9_u2_n99 ) );
  AOI21_X1 u0_u9_u2_U7 (.ZN( u0_u9_u2_n124 ) , .B1( u0_u9_u2_n131 ) , .B2( u0_u9_u2_n143 ) , .A( u0_u9_u2_n172 ) );
  NOR2_X1 u0_u9_u2_U70 (.A2( u0_u9_X_16 ) , .ZN( u0_u9_u2_n140 ) , .A1( u0_u9_u2_n166 ) );
  NOR2_X1 u0_u9_u2_U71 (.A2( u0_u9_X_13 ) , .A1( u0_u9_X_14 ) , .ZN( u0_u9_u2_n100 ) );
  NOR2_X1 u0_u9_u2_U72 (.A2( u0_u9_X_16 ) , .A1( u0_u9_X_17 ) , .ZN( u0_u9_u2_n138 ) );
  NOR2_X1 u0_u9_u2_U73 (.A2( u0_u9_X_15 ) , .A1( u0_u9_X_18 ) , .ZN( u0_u9_u2_n104 ) );
  NOR2_X1 u0_u9_u2_U74 (.A2( u0_u9_X_14 ) , .ZN( u0_u9_u2_n103 ) , .A1( u0_u9_u2_n174 ) );
  NOR2_X1 u0_u9_u2_U75 (.A2( u0_u9_X_15 ) , .ZN( u0_u9_u2_n102 ) , .A1( u0_u9_u2_n165 ) );
  NOR2_X1 u0_u9_u2_U76 (.A2( u0_u9_X_17 ) , .ZN( u0_u9_u2_n114 ) , .A1( u0_u9_u2_n169 ) );
  AND2_X1 u0_u9_u2_U77 (.A1( u0_u9_X_15 ) , .ZN( u0_u9_u2_n105 ) , .A2( u0_u9_u2_n165 ) );
  AND2_X1 u0_u9_u2_U78 (.A2( u0_u9_X_15 ) , .A1( u0_u9_X_18 ) , .ZN( u0_u9_u2_n107 ) );
  AND2_X1 u0_u9_u2_U79 (.A1( u0_u9_X_14 ) , .ZN( u0_u9_u2_n106 ) , .A2( u0_u9_u2_n174 ) );
  AOI21_X1 u0_u9_u2_U8 (.B2( u0_u9_u2_n120 ) , .B1( u0_u9_u2_n121 ) , .ZN( u0_u9_u2_n126 ) , .A( u0_u9_u2_n167 ) );
  AND2_X1 u0_u9_u2_U80 (.A1( u0_u9_X_13 ) , .A2( u0_u9_X_14 ) , .ZN( u0_u9_u2_n108 ) );
  INV_X1 u0_u9_u2_U81 (.A( u0_u9_X_16 ) , .ZN( u0_u9_u2_n169 ) );
  INV_X1 u0_u9_u2_U82 (.A( u0_u9_X_17 ) , .ZN( u0_u9_u2_n166 ) );
  INV_X1 u0_u9_u2_U83 (.A( u0_u9_X_13 ) , .ZN( u0_u9_u2_n174 ) );
  INV_X1 u0_u9_u2_U84 (.A( u0_u9_X_18 ) , .ZN( u0_u9_u2_n165 ) );
  NAND4_X1 u0_u9_u2_U85 (.ZN( u0_out9_30 ) , .A4( u0_u9_u2_n147 ) , .A3( u0_u9_u2_n148 ) , .A2( u0_u9_u2_n149 ) , .A1( u0_u9_u2_n187 ) );
  AOI21_X1 u0_u9_u2_U86 (.B2( u0_u9_u2_n138 ) , .ZN( u0_u9_u2_n148 ) , .A( u0_u9_u2_n162 ) , .B1( u0_u9_u2_n182 ) );
  NOR3_X1 u0_u9_u2_U87 (.A3( u0_u9_u2_n144 ) , .A2( u0_u9_u2_n145 ) , .A1( u0_u9_u2_n146 ) , .ZN( u0_u9_u2_n147 ) );
  NAND4_X1 u0_u9_u2_U88 (.ZN( u0_out9_24 ) , .A4( u0_u9_u2_n111 ) , .A3( u0_u9_u2_n112 ) , .A1( u0_u9_u2_n130 ) , .A2( u0_u9_u2_n187 ) );
  AOI221_X1 u0_u9_u2_U89 (.A( u0_u9_u2_n109 ) , .B1( u0_u9_u2_n110 ) , .ZN( u0_u9_u2_n111 ) , .C1( u0_u9_u2_n134 ) , .C2( u0_u9_u2_n170 ) , .B2( u0_u9_u2_n173 ) );
  OAI22_X1 u0_u9_u2_U9 (.ZN( u0_u9_u2_n109 ) , .A2( u0_u9_u2_n113 ) , .B2( u0_u9_u2_n133 ) , .B1( u0_u9_u2_n167 ) , .A1( u0_u9_u2_n168 ) );
  AOI21_X1 u0_u9_u2_U90 (.ZN( u0_u9_u2_n112 ) , .B2( u0_u9_u2_n156 ) , .A( u0_u9_u2_n164 ) , .B1( u0_u9_u2_n181 ) );
  NAND4_X1 u0_u9_u2_U91 (.ZN( u0_out9_16 ) , .A4( u0_u9_u2_n128 ) , .A3( u0_u9_u2_n129 ) , .A1( u0_u9_u2_n130 ) , .A2( u0_u9_u2_n186 ) );
  AOI22_X1 u0_u9_u2_U92 (.A2( u0_u9_u2_n118 ) , .ZN( u0_u9_u2_n129 ) , .A1( u0_u9_u2_n140 ) , .B1( u0_u9_u2_n157 ) , .B2( u0_u9_u2_n170 ) );
  INV_X1 u0_u9_u2_U93 (.A( u0_u9_u2_n163 ) , .ZN( u0_u9_u2_n186 ) );
  OR4_X1 u0_u9_u2_U94 (.ZN( u0_out9_6 ) , .A4( u0_u9_u2_n161 ) , .A3( u0_u9_u2_n162 ) , .A2( u0_u9_u2_n163 ) , .A1( u0_u9_u2_n164 ) );
  OR3_X1 u0_u9_u2_U95 (.A2( u0_u9_u2_n159 ) , .A1( u0_u9_u2_n160 ) , .ZN( u0_u9_u2_n161 ) , .A3( u0_u9_u2_n183 ) );
  AOI21_X1 u0_u9_u2_U96 (.B2( u0_u9_u2_n154 ) , .B1( u0_u9_u2_n155 ) , .ZN( u0_u9_u2_n159 ) , .A( u0_u9_u2_n167 ) );
  NAND3_X1 u0_u9_u2_U97 (.A2( u0_u9_u2_n117 ) , .A1( u0_u9_u2_n122 ) , .A3( u0_u9_u2_n123 ) , .ZN( u0_u9_u2_n134 ) );
  NAND3_X1 u0_u9_u2_U98 (.ZN( u0_u9_u2_n110 ) , .A2( u0_u9_u2_n131 ) , .A3( u0_u9_u2_n139 ) , .A1( u0_u9_u2_n154 ) );
  NAND3_X1 u0_u9_u2_U99 (.A2( u0_u9_u2_n100 ) , .ZN( u0_u9_u2_n101 ) , .A1( u0_u9_u2_n104 ) , .A3( u0_u9_u2_n114 ) );
  OAI22_X1 u0_u9_u3_U10 (.B1( u0_u9_u3_n113 ) , .A2( u0_u9_u3_n135 ) , .A1( u0_u9_u3_n150 ) , .B2( u0_u9_u3_n164 ) , .ZN( u0_u9_u3_n98 ) );
  OAI211_X1 u0_u9_u3_U11 (.B( u0_u9_u3_n106 ) , .ZN( u0_u9_u3_n119 ) , .C2( u0_u9_u3_n128 ) , .C1( u0_u9_u3_n167 ) , .A( u0_u9_u3_n181 ) );
  AOI221_X1 u0_u9_u3_U12 (.C1( u0_u9_u3_n105 ) , .ZN( u0_u9_u3_n106 ) , .A( u0_u9_u3_n131 ) , .B2( u0_u9_u3_n132 ) , .C2( u0_u9_u3_n133 ) , .B1( u0_u9_u3_n169 ) );
  INV_X1 u0_u9_u3_U13 (.ZN( u0_u9_u3_n181 ) , .A( u0_u9_u3_n98 ) );
  NAND2_X1 u0_u9_u3_U14 (.ZN( u0_u9_u3_n105 ) , .A2( u0_u9_u3_n130 ) , .A1( u0_u9_u3_n155 ) );
  AOI22_X1 u0_u9_u3_U15 (.B1( u0_u9_u3_n115 ) , .A2( u0_u9_u3_n116 ) , .ZN( u0_u9_u3_n123 ) , .B2( u0_u9_u3_n133 ) , .A1( u0_u9_u3_n169 ) );
  NAND2_X1 u0_u9_u3_U16 (.ZN( u0_u9_u3_n116 ) , .A2( u0_u9_u3_n151 ) , .A1( u0_u9_u3_n182 ) );
  NOR2_X1 u0_u9_u3_U17 (.ZN( u0_u9_u3_n126 ) , .A2( u0_u9_u3_n150 ) , .A1( u0_u9_u3_n164 ) );
  AOI21_X1 u0_u9_u3_U18 (.ZN( u0_u9_u3_n112 ) , .B2( u0_u9_u3_n146 ) , .B1( u0_u9_u3_n155 ) , .A( u0_u9_u3_n167 ) );
  NAND2_X1 u0_u9_u3_U19 (.A1( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n142 ) , .A2( u0_u9_u3_n164 ) );
  NAND2_X1 u0_u9_u3_U20 (.ZN( u0_u9_u3_n132 ) , .A2( u0_u9_u3_n152 ) , .A1( u0_u9_u3_n156 ) );
  AND2_X1 u0_u9_u3_U21 (.A2( u0_u9_u3_n113 ) , .A1( u0_u9_u3_n114 ) , .ZN( u0_u9_u3_n151 ) );
  INV_X1 u0_u9_u3_U22 (.A( u0_u9_u3_n133 ) , .ZN( u0_u9_u3_n165 ) );
  INV_X1 u0_u9_u3_U23 (.A( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n170 ) );
  NAND2_X1 u0_u9_u3_U24 (.A1( u0_u9_u3_n107 ) , .A2( u0_u9_u3_n108 ) , .ZN( u0_u9_u3_n140 ) );
  NAND2_X1 u0_u9_u3_U25 (.ZN( u0_u9_u3_n117 ) , .A1( u0_u9_u3_n124 ) , .A2( u0_u9_u3_n148 ) );
  NAND2_X1 u0_u9_u3_U26 (.ZN( u0_u9_u3_n143 ) , .A1( u0_u9_u3_n165 ) , .A2( u0_u9_u3_n167 ) );
  INV_X1 u0_u9_u3_U27 (.A( u0_u9_u3_n130 ) , .ZN( u0_u9_u3_n177 ) );
  INV_X1 u0_u9_u3_U28 (.A( u0_u9_u3_n128 ) , .ZN( u0_u9_u3_n176 ) );
  INV_X1 u0_u9_u3_U29 (.A( u0_u9_u3_n155 ) , .ZN( u0_u9_u3_n174 ) );
  INV_X1 u0_u9_u3_U3 (.A( u0_u9_u3_n129 ) , .ZN( u0_u9_u3_n183 ) );
  INV_X1 u0_u9_u3_U30 (.A( u0_u9_u3_n139 ) , .ZN( u0_u9_u3_n185 ) );
  NOR2_X1 u0_u9_u3_U31 (.ZN( u0_u9_u3_n135 ) , .A2( u0_u9_u3_n141 ) , .A1( u0_u9_u3_n169 ) );
  OAI222_X1 u0_u9_u3_U32 (.C2( u0_u9_u3_n107 ) , .A2( u0_u9_u3_n108 ) , .B1( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n138 ) , .B2( u0_u9_u3_n146 ) , .C1( u0_u9_u3_n154 ) , .A1( u0_u9_u3_n164 ) );
  NOR4_X1 u0_u9_u3_U33 (.A4( u0_u9_u3_n157 ) , .A3( u0_u9_u3_n158 ) , .A2( u0_u9_u3_n159 ) , .A1( u0_u9_u3_n160 ) , .ZN( u0_u9_u3_n161 ) );
  AOI21_X1 u0_u9_u3_U34 (.B2( u0_u9_u3_n152 ) , .B1( u0_u9_u3_n153 ) , .ZN( u0_u9_u3_n158 ) , .A( u0_u9_u3_n164 ) );
  AOI21_X1 u0_u9_u3_U35 (.A( u0_u9_u3_n154 ) , .B2( u0_u9_u3_n155 ) , .B1( u0_u9_u3_n156 ) , .ZN( u0_u9_u3_n157 ) );
  AOI21_X1 u0_u9_u3_U36 (.A( u0_u9_u3_n149 ) , .B2( u0_u9_u3_n150 ) , .B1( u0_u9_u3_n151 ) , .ZN( u0_u9_u3_n159 ) );
  AOI211_X1 u0_u9_u3_U37 (.ZN( u0_u9_u3_n109 ) , .A( u0_u9_u3_n119 ) , .C2( u0_u9_u3_n129 ) , .B( u0_u9_u3_n138 ) , .C1( u0_u9_u3_n141 ) );
  AOI211_X1 u0_u9_u3_U38 (.B( u0_u9_u3_n119 ) , .A( u0_u9_u3_n120 ) , .C2( u0_u9_u3_n121 ) , .ZN( u0_u9_u3_n122 ) , .C1( u0_u9_u3_n179 ) );
  INV_X1 u0_u9_u3_U39 (.A( u0_u9_u3_n156 ) , .ZN( u0_u9_u3_n179 ) );
  INV_X1 u0_u9_u3_U4 (.A( u0_u9_u3_n140 ) , .ZN( u0_u9_u3_n182 ) );
  OAI22_X1 u0_u9_u3_U40 (.B1( u0_u9_u3_n118 ) , .ZN( u0_u9_u3_n120 ) , .A1( u0_u9_u3_n135 ) , .B2( u0_u9_u3_n154 ) , .A2( u0_u9_u3_n178 ) );
  AND3_X1 u0_u9_u3_U41 (.ZN( u0_u9_u3_n118 ) , .A2( u0_u9_u3_n124 ) , .A1( u0_u9_u3_n144 ) , .A3( u0_u9_u3_n152 ) );
  INV_X1 u0_u9_u3_U42 (.A( u0_u9_u3_n121 ) , .ZN( u0_u9_u3_n164 ) );
  NAND2_X1 u0_u9_u3_U43 (.ZN( u0_u9_u3_n133 ) , .A1( u0_u9_u3_n154 ) , .A2( u0_u9_u3_n164 ) );
  OAI211_X1 u0_u9_u3_U44 (.B( u0_u9_u3_n127 ) , .ZN( u0_u9_u3_n139 ) , .C1( u0_u9_u3_n150 ) , .C2( u0_u9_u3_n154 ) , .A( u0_u9_u3_n184 ) );
  INV_X1 u0_u9_u3_U45 (.A( u0_u9_u3_n125 ) , .ZN( u0_u9_u3_n184 ) );
  AOI221_X1 u0_u9_u3_U46 (.A( u0_u9_u3_n126 ) , .ZN( u0_u9_u3_n127 ) , .C2( u0_u9_u3_n132 ) , .C1( u0_u9_u3_n169 ) , .B2( u0_u9_u3_n170 ) , .B1( u0_u9_u3_n174 ) );
  OAI22_X1 u0_u9_u3_U47 (.A1( u0_u9_u3_n124 ) , .ZN( u0_u9_u3_n125 ) , .B2( u0_u9_u3_n145 ) , .A2( u0_u9_u3_n165 ) , .B1( u0_u9_u3_n167 ) );
  NOR2_X1 u0_u9_u3_U48 (.A1( u0_u9_u3_n113 ) , .ZN( u0_u9_u3_n131 ) , .A2( u0_u9_u3_n154 ) );
  NAND2_X1 u0_u9_u3_U49 (.A1( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n150 ) , .A2( u0_u9_u3_n99 ) );
  INV_X1 u0_u9_u3_U5 (.A( u0_u9_u3_n117 ) , .ZN( u0_u9_u3_n178 ) );
  NAND2_X1 u0_u9_u3_U50 (.A2( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n155 ) , .A1( u0_u9_u3_n97 ) );
  INV_X1 u0_u9_u3_U51 (.A( u0_u9_u3_n141 ) , .ZN( u0_u9_u3_n167 ) );
  AOI21_X1 u0_u9_u3_U52 (.B2( u0_u9_u3_n114 ) , .B1( u0_u9_u3_n146 ) , .A( u0_u9_u3_n154 ) , .ZN( u0_u9_u3_n94 ) );
  AOI21_X1 u0_u9_u3_U53 (.ZN( u0_u9_u3_n110 ) , .B2( u0_u9_u3_n142 ) , .B1( u0_u9_u3_n186 ) , .A( u0_u9_u3_n95 ) );
  INV_X1 u0_u9_u3_U54 (.A( u0_u9_u3_n145 ) , .ZN( u0_u9_u3_n186 ) );
  AOI21_X1 u0_u9_u3_U55 (.B1( u0_u9_u3_n124 ) , .A( u0_u9_u3_n149 ) , .B2( u0_u9_u3_n155 ) , .ZN( u0_u9_u3_n95 ) );
  INV_X1 u0_u9_u3_U56 (.A( u0_u9_u3_n149 ) , .ZN( u0_u9_u3_n169 ) );
  NAND2_X1 u0_u9_u3_U57 (.ZN( u0_u9_u3_n124 ) , .A1( u0_u9_u3_n96 ) , .A2( u0_u9_u3_n97 ) );
  NAND2_X1 u0_u9_u3_U58 (.A2( u0_u9_u3_n100 ) , .ZN( u0_u9_u3_n146 ) , .A1( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U59 (.A1( u0_u9_u3_n101 ) , .ZN( u0_u9_u3_n145 ) , .A2( u0_u9_u3_n99 ) );
  AOI221_X1 u0_u9_u3_U6 (.A( u0_u9_u3_n131 ) , .C2( u0_u9_u3_n132 ) , .C1( u0_u9_u3_n133 ) , .ZN( u0_u9_u3_n134 ) , .B1( u0_u9_u3_n143 ) , .B2( u0_u9_u3_n177 ) );
  NAND2_X1 u0_u9_u3_U60 (.A1( u0_u9_u3_n100 ) , .ZN( u0_u9_u3_n156 ) , .A2( u0_u9_u3_n99 ) );
  NAND2_X1 u0_u9_u3_U61 (.A2( u0_u9_u3_n101 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n148 ) );
  NAND2_X1 u0_u9_u3_U62 (.A1( u0_u9_u3_n100 ) , .A2( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n128 ) );
  NAND2_X1 u0_u9_u3_U63 (.A2( u0_u9_u3_n101 ) , .A1( u0_u9_u3_n102 ) , .ZN( u0_u9_u3_n152 ) );
  NAND2_X1 u0_u9_u3_U64 (.A2( u0_u9_u3_n101 ) , .ZN( u0_u9_u3_n114 ) , .A1( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U65 (.ZN( u0_u9_u3_n107 ) , .A1( u0_u9_u3_n97 ) , .A2( u0_u9_u3_n99 ) );
  NAND2_X1 u0_u9_u3_U66 (.A2( u0_u9_u3_n100 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n113 ) );
  NAND2_X1 u0_u9_u3_U67 (.A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n153 ) , .A2( u0_u9_u3_n97 ) );
  NAND2_X1 u0_u9_u3_U68 (.A2( u0_u9_u3_n103 ) , .A1( u0_u9_u3_n104 ) , .ZN( u0_u9_u3_n130 ) );
  NAND2_X1 u0_u9_u3_U69 (.A2( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n144 ) , .A1( u0_u9_u3_n96 ) );
  OAI22_X1 u0_u9_u3_U7 (.B2( u0_u9_u3_n147 ) , .A2( u0_u9_u3_n148 ) , .ZN( u0_u9_u3_n160 ) , .B1( u0_u9_u3_n165 ) , .A1( u0_u9_u3_n168 ) );
  NAND2_X1 u0_u9_u3_U70 (.A1( u0_u9_u3_n102 ) , .A2( u0_u9_u3_n103 ) , .ZN( u0_u9_u3_n108 ) );
  NOR2_X1 u0_u9_u3_U71 (.A2( u0_u9_X_19 ) , .A1( u0_u9_X_20 ) , .ZN( u0_u9_u3_n99 ) );
  NOR2_X1 u0_u9_u3_U72 (.A2( u0_u9_X_21 ) , .A1( u0_u9_X_24 ) , .ZN( u0_u9_u3_n103 ) );
  NOR2_X1 u0_u9_u3_U73 (.A2( u0_u9_X_24 ) , .A1( u0_u9_u3_n171 ) , .ZN( u0_u9_u3_n97 ) );
  NOR2_X1 u0_u9_u3_U74 (.A2( u0_u9_X_23 ) , .ZN( u0_u9_u3_n141 ) , .A1( u0_u9_u3_n166 ) );
  NOR2_X1 u0_u9_u3_U75 (.A2( u0_u9_X_19 ) , .A1( u0_u9_u3_n172 ) , .ZN( u0_u9_u3_n96 ) );
  NAND2_X1 u0_u9_u3_U76 (.A1( u0_u9_X_22 ) , .A2( u0_u9_X_23 ) , .ZN( u0_u9_u3_n154 ) );
  NAND2_X1 u0_u9_u3_U77 (.A1( u0_u9_X_23 ) , .ZN( u0_u9_u3_n149 ) , .A2( u0_u9_u3_n166 ) );
  NOR2_X1 u0_u9_u3_U78 (.A2( u0_u9_X_22 ) , .A1( u0_u9_X_23 ) , .ZN( u0_u9_u3_n121 ) );
  AND2_X1 u0_u9_u3_U79 (.A1( u0_u9_X_24 ) , .ZN( u0_u9_u3_n101 ) , .A2( u0_u9_u3_n171 ) );
  AND3_X1 u0_u9_u3_U8 (.A3( u0_u9_u3_n144 ) , .A2( u0_u9_u3_n145 ) , .A1( u0_u9_u3_n146 ) , .ZN( u0_u9_u3_n147 ) );
  AND2_X1 u0_u9_u3_U80 (.A1( u0_u9_X_19 ) , .ZN( u0_u9_u3_n102 ) , .A2( u0_u9_u3_n172 ) );
  AND2_X1 u0_u9_u3_U81 (.A1( u0_u9_X_21 ) , .A2( u0_u9_X_24 ) , .ZN( u0_u9_u3_n100 ) );
  AND2_X1 u0_u9_u3_U82 (.A2( u0_u9_X_19 ) , .A1( u0_u9_X_20 ) , .ZN( u0_u9_u3_n104 ) );
  INV_X1 u0_u9_u3_U83 (.A( u0_u9_X_22 ) , .ZN( u0_u9_u3_n166 ) );
  INV_X1 u0_u9_u3_U84 (.A( u0_u9_X_21 ) , .ZN( u0_u9_u3_n171 ) );
  INV_X1 u0_u9_u3_U85 (.A( u0_u9_X_20 ) , .ZN( u0_u9_u3_n172 ) );
  OR4_X1 u0_u9_u3_U86 (.ZN( u0_out9_10 ) , .A4( u0_u9_u3_n136 ) , .A3( u0_u9_u3_n137 ) , .A1( u0_u9_u3_n138 ) , .A2( u0_u9_u3_n139 ) );
  OAI222_X1 u0_u9_u3_U87 (.C1( u0_u9_u3_n128 ) , .ZN( u0_u9_u3_n137 ) , .B1( u0_u9_u3_n148 ) , .A2( u0_u9_u3_n150 ) , .B2( u0_u9_u3_n154 ) , .C2( u0_u9_u3_n164 ) , .A1( u0_u9_u3_n167 ) );
  OAI221_X1 u0_u9_u3_U88 (.A( u0_u9_u3_n134 ) , .B2( u0_u9_u3_n135 ) , .ZN( u0_u9_u3_n136 ) , .C1( u0_u9_u3_n149 ) , .B1( u0_u9_u3_n151 ) , .C2( u0_u9_u3_n183 ) );
  NAND4_X1 u0_u9_u3_U89 (.ZN( u0_out9_26 ) , .A4( u0_u9_u3_n109 ) , .A3( u0_u9_u3_n110 ) , .A2( u0_u9_u3_n111 ) , .A1( u0_u9_u3_n173 ) );
  INV_X1 u0_u9_u3_U9 (.A( u0_u9_u3_n143 ) , .ZN( u0_u9_u3_n168 ) );
  INV_X1 u0_u9_u3_U90 (.ZN( u0_u9_u3_n173 ) , .A( u0_u9_u3_n94 ) );
  OAI21_X1 u0_u9_u3_U91 (.ZN( u0_u9_u3_n111 ) , .B2( u0_u9_u3_n117 ) , .A( u0_u9_u3_n133 ) , .B1( u0_u9_u3_n176 ) );
  NAND4_X1 u0_u9_u3_U92 (.ZN( u0_out9_20 ) , .A4( u0_u9_u3_n122 ) , .A3( u0_u9_u3_n123 ) , .A1( u0_u9_u3_n175 ) , .A2( u0_u9_u3_n180 ) );
  INV_X1 u0_u9_u3_U93 (.A( u0_u9_u3_n126 ) , .ZN( u0_u9_u3_n180 ) );
  INV_X1 u0_u9_u3_U94 (.A( u0_u9_u3_n112 ) , .ZN( u0_u9_u3_n175 ) );
  NAND4_X1 u0_u9_u3_U95 (.ZN( u0_out9_1 ) , .A4( u0_u9_u3_n161 ) , .A3( u0_u9_u3_n162 ) , .A2( u0_u9_u3_n163 ) , .A1( u0_u9_u3_n185 ) );
  NAND2_X1 u0_u9_u3_U96 (.ZN( u0_u9_u3_n163 ) , .A2( u0_u9_u3_n170 ) , .A1( u0_u9_u3_n176 ) );
  AOI22_X1 u0_u9_u3_U97 (.B2( u0_u9_u3_n140 ) , .B1( u0_u9_u3_n141 ) , .A2( u0_u9_u3_n142 ) , .ZN( u0_u9_u3_n162 ) , .A1( u0_u9_u3_n177 ) );
  NAND3_X1 u0_u9_u3_U98 (.A1( u0_u9_u3_n114 ) , .ZN( u0_u9_u3_n115 ) , .A2( u0_u9_u3_n145 ) , .A3( u0_u9_u3_n153 ) );
  NAND3_X1 u0_u9_u3_U99 (.ZN( u0_u9_u3_n129 ) , .A2( u0_u9_u3_n144 ) , .A1( u0_u9_u3_n153 ) , .A3( u0_u9_u3_n182 ) );
  OAI22_X1 u0_uk_U101 (.ZN( u0_K9_5 ) , .A1( u0_uk_n142 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n272 ) , .B2( u0_uk_n278 ) );
  OAI21_X1 u0_uk_U1012 (.ZN( u0_K10_21 ) , .A( u0_uk_n1020 ) , .B2( u0_uk_n228 ) , .B1( u0_uk_n31 ) );
  OAI21_X1 u0_uk_U1022 (.ZN( u0_K9_44 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n273 ) , .A( u0_uk_n721 ) );
  NAND2_X1 u0_uk_U1023 (.A1( u0_uk_K_r7_0 ) , .A2( u0_uk_n217 ) , .ZN( u0_uk_n721 ) );
  OAI21_X1 u0_uk_U1030 (.ZN( u0_K16_41 ) , .B1( u0_uk_n142 ) , .B2( u0_uk_n643 ) , .A( u0_uk_n898 ) );
  NAND2_X1 u0_uk_U1035 (.A1( u0_uk_K_r4_31 ) , .ZN( u0_uk_n790 ) , .A2( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U1039 (.A1( u0_uk_K_r6_51 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n756 ) );
  OAI21_X1 u0_uk_U1044 (.ZN( u0_K15_14 ) , .B2( u0_uk_n37 ) , .B1( u0_uk_n92 ) , .A( u0_uk_n923 ) );
  NAND2_X1 u0_uk_U1045 (.A1( u0_uk_K_r13_32 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n923 ) );
  OAI21_X1 u0_uk_U1050 (.ZN( u0_K15_32 ) , .B1( u0_uk_n31 ) , .B2( u0_uk_n33 ) , .A( u0_uk_n918 ) );
  OAI21_X1 u0_uk_U1052 (.ZN( u0_K16_42 ) , .B2( u0_uk_n647 ) , .A( u0_uk_n897 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U1085 (.ZN( u0_K13_28 ) , .B2( u0_uk_n105 ) , .B1( u0_uk_n252 ) , .A( u0_uk_n947 ) );
  NAND2_X1 u0_uk_U1086 (.A1( u0_uk_K_r11_21 ) , .A2( u0_uk_n214 ) , .ZN( u0_uk_n947 ) );
  OAI21_X1 u0_uk_U1093 (.ZN( u0_K16_39 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n657 ) , .A( u0_uk_n899 ) );
  NAND2_X1 u0_uk_U1094 (.A1( u0_uk_K_r14_15 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n899 ) );
  OAI22_X1 u0_uk_U112 (.ZN( u0_K16_47 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n666 ) , .B2( u0_uk_n670 ) );
  INV_X1 u0_uk_U1141 (.ZN( u0_K10_12 ) , .A( u0_uk_n1024 ) );
  AOI22_X1 u0_uk_U1153 (.B2( u0_uk_K_r7_24 ) , .A2( u0_uk_K_r7_6 ) , .B1( u0_uk_n10 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n734 ) );
  INV_X1 u0_uk_U1154 (.ZN( u0_K9_1 ) , .A( u0_uk_n734 ) );
  AOI22_X1 u0_uk_U1162 (.B2( u0_uk_K_r7_20 ) , .A2( u0_uk_K_r7_27 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n729 ) );
  INV_X1 u0_uk_U1163 (.ZN( u0_K9_2 ) , .A( u0_uk_n729 ) );
  INV_X1 u0_uk_U12 (.A( u0_uk_n187 ) , .ZN( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U146 (.ZN( u0_K10_15 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n229 ) , .A2( u0_uk_n266 ) , .A1( u0_uk_n94 ) );
  OAI21_X1 u0_uk_U147 (.ZN( u0_K15_15 ) , .B2( u0_uk_n15 ) , .B1( u0_uk_n163 ) , .A( u0_uk_n922 ) );
  NAND2_X1 u0_uk_U148 (.A1( u0_uk_K_r13_19 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n922 ) );
  INV_X1 u0_uk_U15 (.A( u0_uk_n155 ) , .ZN( u0_uk_n99 ) );
  INV_X1 u0_uk_U153 (.ZN( u0_K9_19 ) , .A( u0_uk_n735 ) );
  OAI22_X1 u0_uk_U155 (.ZN( u0_K7_19 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n383 ) , .B2( u0_uk_n393 ) );
  OAI21_X1 u0_uk_U182 (.ZN( u0_K10_24 ) , .A( u0_uk_n1017 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n259 ) );
  NAND2_X1 u0_uk_U183 (.A1( u0_uk_K_r8_40 ) , .ZN( u0_uk_n1017 ) , .A2( u0_uk_n11 ) );
  INV_X1 u0_uk_U190 (.ZN( u0_K11_30 ) , .A( u0_uk_n993 ) );
  AOI22_X1 u0_uk_U191 (.B2( u0_uk_K_r9_1 ) , .A2( u0_uk_K_r9_9 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n163 ) , .ZN( u0_uk_n993 ) );
  INV_X1 u0_uk_U195 (.ZN( u0_K7_24 ) , .A( u0_uk_n776 ) );
  AOI22_X1 u0_uk_U196 (.B2( u0_uk_K_r5_18 ) , .A2( u0_uk_K_r5_40 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n162 ) , .ZN( u0_uk_n776 ) );
  OAI22_X1 u0_uk_U200 (.ZN( u0_K15_24 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n24 ) , .A2( u0_uk_n42 ) );
  OAI21_X1 u0_uk_U203 (.ZN( u0_K9_30 ) , .B2( u0_uk_n288 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n728 ) );
  OAI22_X1 u0_uk_U214 (.ZN( u0_K16_31 ) , .B1( u0_uk_n155 ) , .B2( u0_uk_n663 ) , .A2( u0_uk_n666 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U22 (.ZN( u0_uk_n128 ) , .A( u0_uk_n214 ) );
  OAI22_X1 u0_uk_U230 (.ZN( u0_K15_31 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n28 ) , .B2( u0_uk_n45 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U241 (.ZN( u0_K16_48 ) , .B1( u0_uk_n102 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n650 ) , .B2( u0_uk_n658 ) );
  OAI21_X1 u0_uk_U242 (.ZN( u0_K16_44 ) , .B1( u0_uk_n110 ) , .B2( u0_uk_n642 ) , .A( u0_uk_n895 ) );
  NAND2_X1 u0_uk_U243 (.A1( u0_uk_K_r14_43 ) , .ZN( u0_uk_n895 ) , .A2( u0_uk_n99 ) );
  INV_X1 u0_uk_U264 (.ZN( u0_K9_48 ) , .A( u0_uk_n719 ) );
  INV_X1 u0_uk_U284 (.ZN( u0_K15_8 ) , .A( u0_uk_n913 ) );
  AOI22_X1 u0_uk_U285 (.B2( u0_uk_K_r13_13 ) , .A2( u0_uk_K_r13_17 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n230 ) , .ZN( u0_uk_n913 ) );
  OAI22_X1 u0_uk_U296 (.ZN( u0_K7_26 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n230 ) , .A2( u0_uk_n368 ) , .B2( u0_uk_n388 ) );
  INV_X1 u0_uk_U300 (.ZN( u0_K9_26 ) , .A( u0_uk_n731 ) );
  OAI21_X1 u0_uk_U306 (.ZN( u0_K6_26 ) , .B1( u0_uk_n217 ) , .B2( u0_uk_n419 ) , .A( u0_uk_n795 ) );
  NAND2_X1 u0_uk_U307 (.A1( u0_uk_K_r4_35 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n795 ) );
  OAI21_X1 u0_uk_U308 (.ZN( u0_K11_26 ) , .B2( u0_uk_n193 ) , .B1( u0_uk_n93 ) , .A( u0_uk_n995 ) );
  NAND2_X1 u0_uk_U309 (.A1( u0_uk_K_r9_35 ) , .A2( u0_uk_n92 ) , .ZN( u0_uk_n995 ) );
  OAI21_X1 u0_uk_U310 (.ZN( u0_K13_26 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n123 ) , .A( u0_uk_n948 ) );
  OAI21_X1 u0_uk_U323 (.ZN( u0_K9_46 ) , .B1( u0_uk_n11 ) , .B2( u0_uk_n281 ) , .A( u0_uk_n720 ) );
  NAND2_X1 u0_uk_U336 (.A1( u0_uk_K_r14_3 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n894 ) );
  BUF_X1 u0_uk_U35 (.A( u0_uk_n155 ) , .Z( u0_uk_n187 ) );
  OAI22_X1 u0_uk_U351 (.ZN( u0_K16_40 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n632 ) , .B2( u0_uk_n670 ) );
  OAI22_X1 u0_uk_U352 (.ZN( u0_K6_40 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .B2( u0_uk_n438 ) , .A2( u0_uk_n446 ) );
  BUF_X1 u0_uk_U36 (.Z( u0_uk_n188 ) , .A( u0_uk_n230 ) );
  OAI21_X1 u0_uk_U367 (.ZN( u0_K15_33 ) , .B2( u0_uk_n18 ) , .B1( u0_uk_n83 ) , .A( u0_uk_n917 ) );
  OAI22_X1 u0_uk_U374 (.ZN( u0_K11_28 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n184 ) , .B2( u0_uk_n216 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U375 (.ZN( u0_K6_28 ) , .A1( u0_uk_n251 ) , .A2( u0_uk_n411 ) , .B2( u0_uk_n438 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U384 (.ZN( u0_K9_28 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n274 ) , .B2( u0_uk_n281 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U385 (.ZN( u0_K7_28 ) , .A1( u0_uk_n223 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n378 ) , .B2( u0_uk_n387 ) );
  OAI21_X1 u0_uk_U393 (.ZN( u0_K10_16 ) , .A( u0_uk_n1022 ) , .B2( u0_uk_n228 ) , .B1( u0_uk_n250 ) );
  NAND2_X1 u0_uk_U394 (.A1( u0_uk_K_r8_32 ) , .ZN( u0_uk_n1022 ) , .A2( u0_uk_n251 ) );
  OAI22_X1 u0_uk_U395 (.ZN( u0_K9_16 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n231 ) , .A2( u0_uk_n303 ) , .B2( u0_uk_n310 ) );
  OAI21_X1 u0_uk_U402 (.ZN( u0_K15_9 ) , .B2( u0_uk_n15 ) , .A( u0_uk_n912 ) , .B1( u0_uk_n93 ) );
  NAND2_X1 u0_uk_U403 (.A1( u0_uk_K_r13_4 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n912 ) );
  NAND2_X1 u0_uk_U405 (.A1( u0_uk_K_r12_18 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n926 ) );
  INV_X1 u0_uk_U416 (.ZN( u0_K10_9 ) , .A( u0_uk_n1005 ) );
  AOI22_X1 u0_uk_U417 (.B2( u0_uk_K_r8_17 ) , .A2( u0_uk_K_r8_27 ) , .ZN( u0_uk_n1005 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n220 ) );
  INV_X1 u0_uk_U418 (.ZN( u0_K9_9 ) , .A( u0_uk_n718 ) );
  AOI22_X1 u0_uk_U419 (.B2( u0_uk_K_r7_13 ) , .A1( u0_uk_K_r7_6 ) , .A2( u0_uk_n128 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n718 ) );
  OAI22_X1 u0_uk_U434 (.ZN( u0_K15_16 ) , .A2( u0_uk_n14 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n29 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U443 (.ZN( u0_K16_33 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n633 ) , .B2( u0_uk_n638 ) );
  INV_X1 u0_uk_U452 (.ZN( u0_K16_37 ) , .A( u0_uk_n900 ) );
  AOI22_X1 u0_uk_U453 (.B2( u0_uk_K_r14_2 ) , .A2( u0_uk_K_r14_50 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n900 ) );
  OAI21_X1 u0_uk_U461 (.ZN( u0_K6_37 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n420 ) , .A( u0_uk_n791 ) );
  NAND2_X1 u0_uk_U462 (.A1( u0_uk_K_r4_38 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n791 ) );
  OAI22_X1 u0_uk_U474 (.ZN( u0_K13_29 ) , .A2( u0_uk_n113 ) , .B2( u0_uk_n116 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n161 ) );
  OAI21_X1 u0_uk_U475 (.ZN( u0_K11_29 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n224 ) , .A( u0_uk_n994 ) );
  NAND2_X1 u0_uk_U476 (.A1( u0_uk_K_r9_0 ) , .A2( u0_uk_n60 ) , .ZN( u0_uk_n994 ) );
  OAI21_X1 u0_uk_U477 (.ZN( u0_K6_29 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n446 ) , .A( u0_uk_n794 ) );
  NAND2_X1 u0_uk_U478 (.A1( u0_uk_K_r4_0 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n794 ) );
  OAI22_X1 u0_uk_U484 (.ZN( u0_K9_29 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n289 ) , .B2( u0_uk_n293 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U486 (.ZN( u0_K7_29 ) , .A1( u0_uk_n162 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n368 ) , .B2( u0_uk_n399 ) );
  OAI21_X1 u0_uk_U497 (.ZN( u0_K9_12 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n315 ) , .A( u0_uk_n740 ) );
  OAI22_X1 u0_uk_U503 (.ZN( u0_K10_17 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n234 ) , .B2( u0_uk_n262 ) , .A1( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U504 (.ZN( u0_K9_17 ) , .B2( u0_uk_n290 ) , .A( u0_uk_n737 ) , .B1( u0_uk_n99 ) );
  NAND2_X1 u0_uk_U505 (.A1( u0_uk_K_r7_26 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n737 ) );
  OAI22_X1 u0_uk_U518 (.ZN( u0_K15_12 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n231 ) , .B2( u0_uk_n25 ) , .A2( u0_uk_n43 ) );
  OAI22_X1 u0_uk_U537 (.ZN( u0_K15_17 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n220 ) , .B2( u0_uk_n26 ) , .A2( u0_uk_n44 ) );
  OAI22_X1 u0_uk_U544 (.ZN( u0_K15_36 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n18 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n32 ) );
  OAI22_X1 u0_uk_U554 (.ZN( u0_K16_36 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n63 ) , .A2( u0_uk_n648 ) , .B2( u0_uk_n655 ) );
  OAI22_X1 u0_uk_U567 (.ZN( u0_K6_38 ) , .A1( u0_uk_n213 ) , .A2( u0_uk_n433 ) , .B2( u0_uk_n440 ) , .B1( u0_uk_n60 ) );
  OAI21_X1 u0_uk_U572 (.ZN( u0_K15_10 ) , .B1( u0_uk_n128 ) , .B2( u0_uk_n19 ) , .A( u0_uk_n925 ) );
  NAND2_X1 u0_uk_U573 (.A1( u0_uk_K_r13_55 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n925 ) );
  INV_X1 u0_uk_U579 (.ZN( u0_K9_10 ) , .A( u0_uk_n742 ) );
  INV_X1 u0_uk_U58 (.ZN( u0_K16_34 ) , .A( u0_uk_n901 ) );
  AOI22_X1 u0_uk_U580 (.B2( u0_uk_K_r7_25 ) , .A2( u0_uk_K_r7_32 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n242 ) , .ZN( u0_uk_n742 ) );
  AOI22_X1 u0_uk_U59 (.B2( u0_uk_K_r14_2 ) , .A2( u0_uk_K_r14_9 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n202 ) , .ZN( u0_uk_n901 ) );
  INV_X1 u0_uk_U594 (.ZN( u0_K10_22 ) , .A( u0_uk_n1019 ) );
  INV_X1 u0_uk_U596 (.ZN( u0_K9_22 ) , .A( u0_uk_n732 ) );
  OAI22_X1 u0_uk_U603 (.ZN( u0_K16_35 ) , .B1( u0_uk_n100 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n643 ) , .B2( u0_uk_n650 ) );
  OAI22_X1 u0_uk_U611 (.ZN( u0_K15_35 ) , .A2( u0_uk_n13 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n28 ) );
  OAI21_X1 u0_uk_U624 (.ZN( u0_K15_11 ) , .B1( u0_uk_n163 ) , .B2( u0_uk_n8 ) , .A( u0_uk_n924 ) );
  NAND2_X1 u0_uk_U625 (.A1( u0_uk_K_r13_25 ) , .A2( u0_uk_n251 ) , .ZN( u0_uk_n924 ) );
  OAI22_X1 u0_uk_U630 (.ZN( u0_K10_11 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n245 ) , .B2( u0_uk_n262 ) , .B1( u0_uk_n83 ) );
  NAND2_X1 u0_uk_U632 (.A1( u0_uk_K_r6_55 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n762 ) );
  INV_X1 u0_uk_U637 (.ZN( u0_K9_11 ) , .A( u0_uk_n741 ) );
  AOI22_X1 u0_uk_U638 (.B2( u0_uk_K_r7_48 ) , .A2( u0_uk_K_r7_55 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n741 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U64 (.ZN( u0_K15_34 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n32 ) , .A2( u0_uk_n4 ) );
  OAI22_X1 u0_uk_U647 (.ZN( u0_K16_45 ) , .B1( u0_uk_n110 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n638 ) , .B2( u0_uk_n641 ) );
  OAI21_X1 u0_uk_U653 (.ZN( u0_K2_43 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n612 ) , .A( u0_uk_n857 ) );
  NAND2_X1 u0_uk_U654 (.A1( u0_uk_K_r0_2 ) , .A2( u0_uk_n63 ) , .ZN( u0_uk_n857 ) );
  OAI22_X1 u0_uk_U657 (.ZN( u0_K9_25 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n273 ) , .B2( u0_uk_n280 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U658 (.ZN( u0_K16_43 ) , .A( u0_uk_n896 ) );
  AOI22_X1 u0_uk_U659 (.B2( u0_uk_K_r14_16 ) , .A2( u0_uk_K_r14_9 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n191 ) , .ZN( u0_uk_n896 ) );
  OAI22_X1 u0_uk_U671 (.ZN( u0_K9_43 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n155 ) , .A2( u0_uk_n293 ) , .B2( u0_uk_n300 ) );
  OAI22_X1 u0_uk_U678 (.ZN( u0_K10_7 ) , .A1( u0_uk_n223 ) , .A2( u0_uk_n234 ) , .B2( u0_uk_n254 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U679 (.ZN( u0_K15_7 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n19 ) , .B2( u0_uk_n35 ) );
  OAI22_X1 u0_uk_U688 (.ZN( u0_K11_25 ) , .A2( u0_uk_n192 ) , .B2( u0_uk_n211 ) , .A1( u0_uk_n242 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U689 (.ZN( u0_K13_25 ) , .A1( u0_uk_n118 ) , .B2( u0_uk_n123 ) , .B1( u0_uk_n242 ) , .A2( u0_uk_n98 ) );
  INV_X1 u0_uk_U708 (.ZN( u0_K7_25 ) , .A( u0_uk_n775 ) );
  OAI22_X1 u0_uk_U717 (.ZN( u0_K16_32 ) , .B1( u0_uk_n118 ) , .A1( u0_uk_n155 ) , .A2( u0_uk_n649 ) , .B2( u0_uk_n657 ) );
  OAI21_X1 u0_uk_U757 (.ZN( u0_K9_13 ) , .B2( u0_uk_n309 ) , .B1( u0_uk_n63 ) , .A( u0_uk_n739 ) );
  OAI22_X1 u0_uk_U759 (.ZN( u0_K11_27 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n198 ) , .B2( u0_uk_n204 ) );
  OAI22_X1 u0_uk_U760 (.ZN( u0_K13_27 ) , .A2( u0_uk_n111 ) , .B2( u0_uk_n134 ) , .B1( u0_uk_n238 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U764 (.ZN( u0_K9_21 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n285 ) , .B2( u0_uk_n290 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U768 (.ZN( u0_K15_21 ) , .A1( u0_uk_n164 ) , .B2( u0_uk_n38 ) , .A2( u0_uk_n42 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U77 (.ZN( u0_K10_23 ) , .A( u0_uk_n1018 ) , .B1( u0_uk_n147 ) , .B2( u0_uk_n268 ) );
  NAND2_X1 u0_uk_U78 (.A1( u0_uk_K_r8_13 ) , .ZN( u0_uk_n1018 ) , .A2( u0_uk_n252 ) );
  OAI21_X1 u0_uk_U790 (.ZN( u0_K7_21 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n362 ) , .A( u0_uk_n779 ) );
  NAND2_X1 u0_uk_U791 (.A1( u0_uk_K_r5_19 ) , .A2( u0_uk_n252 ) , .ZN( u0_uk_n779 ) );
  INV_X1 u0_uk_U792 (.ZN( u0_K7_27 ) , .A( u0_uk_n774 ) );
  AOI22_X1 u0_uk_U793 (.B2( u0_uk_K_r5_23 ) , .A2( u0_uk_K_r5_43 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n223 ) , .ZN( u0_uk_n774 ) );
  INV_X1 u0_uk_U796 (.ZN( u0_K9_27 ) , .A( u0_uk_n730 ) );
  AOI22_X1 u0_uk_U797 (.B2( u0_uk_K_r7_2 ) , .A2( u0_uk_K_r7_9 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n730 ) , .B1( u0_uk_n94 ) );
  NAND2_X1 u0_uk_U816 (.A1( u0_uk_K_r14_5 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n906 ) );
  OAI22_X1 u0_uk_U823 (.ZN( u0_K15_20 ) , .B2( u0_uk_n14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n43 ) , .B1( u0_uk_n92 ) );
  INV_X1 u0_uk_U825 (.ZN( u0_K9_18 ) , .A( u0_uk_n736 ) );
  INV_X1 u0_uk_U831 (.ZN( u0_K9_20 ) , .A( u0_uk_n733 ) );
  AOI22_X1 u0_uk_U832 (.B2( u0_uk_K_r7_32 ) , .A2( u0_uk_K_r7_39 ) , .B1( u0_uk_n10 ) , .A1( u0_uk_n240 ) , .ZN( u0_uk_n733 ) );
  INV_X1 u0_uk_U833 (.ZN( u0_K7_20 ) , .A( u0_uk_n780 ) );
  OAI22_X1 u0_uk_U871 (.ZN( u0_K15_22 ) , .A2( u0_uk_n16 ) , .A1( u0_uk_n188 ) , .B2( u0_uk_n30 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U873 (.ZN( u0_K15_23 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n25 ) , .A2( u0_uk_n7 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U895 (.ZN( u0_K9_3 ) , .A1( u0_uk_n161 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n311 ) , .A2( u0_uk_n315 ) );
  OAI22_X1 u0_uk_U896 (.ZN( u0_K9_7 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n310 ) , .A2( u0_uk_n314 ) );
  OAI22_X1 u0_uk_U902 (.ZN( u0_K15_13 ) , .B2( u0_uk_n16 ) , .A1( u0_uk_n230 ) , .A2( u0_uk_n44 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U904 (.ZN( u0_K9_24 ) , .A1( u0_uk_n257 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n272 ) , .B2( u0_uk_n314 ) );
  OAI22_X1 u0_uk_U911 (.ZN( u0_K7_30 ) , .A1( u0_uk_n213 ) , .B1( u0_uk_n31 ) , .A2( u0_uk_n367 ) , .B2( u0_uk_n398 ) );
  OAI22_X1 u0_uk_U918 (.ZN( u0_K6_30 ) , .A1( u0_uk_n203 ) , .A2( u0_uk_n445 ) , .B2( u0_uk_n450 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U923 (.ZN( u0_K6_42 ) , .A1( u0_uk_n161 ) , .A2( u0_uk_n413 ) , .B2( u0_uk_n420 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U924 (.ZN( u0_K6_39 ) , .A1( u0_uk_n162 ) , .B2( u0_uk_n428 ) , .A2( u0_uk_n447 ) , .B1( u0_uk_n60 ) );
  OAI22_X1 u0_uk_U930 (.ZN( u0_K9_23 ) , .B1( u0_uk_n162 ) , .A2( u0_uk_n296 ) , .B2( u0_uk_n304 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U931 (.ZN( u0_K9_47 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n187 ) , .A2( u0_uk_n275 ) , .B2( u0_uk_n282 ) );
  OAI22_X1 u0_uk_U937 (.ZN( u0_K9_8 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n147 ) , .A2( u0_uk_n278 ) , .B2( u0_uk_n285 ) );
  OAI22_X1 u0_uk_U945 (.ZN( u0_K16_46 ) , .A1( u0_uk_n117 ) , .B1( u0_uk_n223 ) , .A2( u0_uk_n635 ) , .B2( u0_uk_n669 ) );
  OAI22_X1 u0_uk_U956 (.ZN( u0_K10_8 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n182 ) , .B2( u0_uk_n253 ) , .A2( u0_uk_n267 ) );
  OAI22_X1 u0_uk_U962 (.ZN( u0_K15_19 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n37 ) , .A2( u0_uk_n7 ) );
  OAI22_X1 u0_uk_U988 (.ZN( u0_K6_25 ) , .A1( u0_uk_n102 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n418 ) , .B2( u0_uk_n434 ) );
  XOR2_X1 u1_U10 (.B( u1_L1_29 ) , .Z( u1_N92 ) , .A( u1_out2_29 ) );
  XOR2_X1 u1_U109 (.B( u1_L12_19 ) , .Z( u1_N434 ) , .A( u1_out13_19 ) );
  XOR2_X1 u1_U118 (.B( u1_L12_11 ) , .Z( u1_N426 ) , .A( u1_out13_11 ) );
  XOR2_X1 u1_U126 (.B( u1_L12_4 ) , .Z( u1_N419 ) , .A( u1_out13_4 ) );
  XOR2_X1 u1_U130 (.B( u1_L11_32 ) , .Z( u1_N415 ) , .A( u1_out12_32 ) );
  XOR2_X1 u1_U141 (.B( u1_L11_22 ) , .Z( u1_N405 ) , .A( u1_out12_22 ) );
  XOR2_X1 u1_U153 (.B( u1_L11_12 ) , .Z( u1_N395 ) , .A( u1_out12_12 ) );
  XOR2_X1 u1_U158 (.B( u1_L11_7 ) , .Z( u1_N390 ) , .A( u1_out12_7 ) );
  XOR2_X1 u1_U16 (.B( u1_L1_24 ) , .Z( u1_N87 ) , .A( u1_out2_24 ) );
  XOR2_X1 u1_U169 (.B( u1_L10_29 ) , .Z( u1_N380 ) , .A( u1_out11_29 ) );
  XOR2_X1 u1_U180 (.B( u1_L10_19 ) , .Z( u1_N370 ) , .A( u1_out11_19 ) );
  XOR2_X1 u1_U189 (.B( u1_L10_11 ) , .Z( u1_N362 ) , .A( u1_out11_11 ) );
  XOR2_X1 u1_U197 (.B( u1_L10_4 ) , .Z( u1_N355 ) , .A( u1_out11_4 ) );
  XOR2_X1 u1_U202 (.B( u1_L9_31 ) , .Z( u1_N350 ) , .A( u1_out10_31 ) );
  XOR2_X1 u1_U205 (.B( u1_L9_29 ) , .Z( u1_N348 ) , .A( u1_out10_29 ) );
  XOR2_X1 u1_U206 (.B( u1_L9_28 ) , .Z( u1_N347 ) , .A( u1_out10_28 ) );
  XOR2_X1 u1_U209 (.B( u1_L9_25 ) , .Z( u1_N344 ) , .A( u1_out10_25 ) );
  XOR2_X1 u1_U21 (.B( u1_L1_19 ) , .Z( u1_N82 ) , .A( u1_out2_19 ) );
  XOR2_X1 u1_U211 (.B( u1_L9_23 ) , .Z( u1_N342 ) , .A( u1_out10_23 ) );
  XOR2_X1 u1_U216 (.B( u1_L9_19 ) , .Z( u1_N338 ) , .A( u1_out10_19 ) );
  XOR2_X1 u1_U217 (.B( u1_L9_18 ) , .Z( u1_N337 ) , .A( u1_out10_18 ) );
  XOR2_X1 u1_U218 (.B( u1_L9_17 ) , .Z( u1_N336 ) , .A( u1_out10_17 ) );
  XOR2_X1 u1_U221 (.B( u1_L9_14 ) , .Z( u1_N333 ) , .A( u1_out10_14 ) );
  XOR2_X1 u1_U222 (.B( u1_L9_13 ) , .Z( u1_N332 ) , .A( u1_out10_13 ) );
  XOR2_X1 u1_U224 (.B( u1_L9_11 ) , .Z( u1_N330 ) , .A( u1_out10_11 ) );
  XOR2_X1 u1_U227 (.B( u1_L9_9 ) , .Z( u1_N328 ) , .A( u1_out10_9 ) );
  XOR2_X1 u1_U228 (.B( u1_L9_8 ) , .Z( u1_N327 ) , .A( u1_out10_8 ) );
  XOR2_X1 u1_U232 (.B( u1_L9_4 ) , .Z( u1_N323 ) , .A( u1_out10_4 ) );
  XOR2_X1 u1_U233 (.B( u1_L9_3 ) , .Z( u1_N322 ) , .A( u1_out10_3 ) );
  XOR2_X1 u1_U234 (.B( u1_L9_2 ) , .Z( u1_N321 ) , .A( u1_out10_2 ) );
  XOR2_X1 u1_U244 (.B( u1_L8_25 ) , .Z( u1_N312 ) , .A( u1_out9_25 ) );
  XOR2_X1 u1_U25 (.B( u1_L1_16 ) , .Z( u1_N79 ) , .A( u1_out2_16 ) );
  XOR2_X1 u1_U256 (.B( u1_L8_14 ) , .Z( u1_N301 ) , .A( u1_out9_14 ) );
  XOR2_X1 u1_U264 (.B( u1_L8_8 ) , .Z( u1_N295 ) , .A( u1_out9_8 ) );
  XOR2_X1 u1_U269 (.B( u1_L8_3 ) , .Z( u1_N290 ) , .A( u1_out9_3 ) );
  XOR2_X1 u1_U270 (.Z( u1_N29 ) , .B( u1_desIn_r_40 ) , .A( u1_out0_30 ) );
  XOR2_X1 u1_U276 (.B( u1_L7_29 ) , .Z( u1_N284 ) , .A( u1_out8_29 ) );
  XOR2_X1 u1_U287 (.B( u1_L7_19 ) , .Z( u1_N274 ) , .A( u1_out8_19 ) );
  XOR2_X1 u1_U296 (.B( u1_L7_11 ) , .Z( u1_N266 ) , .A( u1_out8_11 ) );
  XOR2_X1 u1_U30 (.B( u1_L1_11 ) , .Z( u1_N74 ) , .A( u1_out2_11 ) );
  XOR2_X1 u1_U304 (.B( u1_L7_4 ) , .Z( u1_N259 ) , .A( u1_out8_4 ) );
  XOR2_X1 u1_U315 (.B( u1_L6_26 ) , .Z( u1_N249 ) , .A( u1_out7_26 ) );
  XOR2_X1 u1_U321 (.B( u1_L6_20 ) , .Z( u1_N243 ) , .A( u1_out7_20 ) );
  XOR2_X1 u1_U332 (.B( u1_L6_10 ) , .Z( u1_N233 ) , .A( u1_out7_10 ) );
  XOR2_X1 u1_U336 (.Z( u1_N23 ) , .B( u1_desIn_r_58 ) , .A( u1_out0_24 ) );
  XOR2_X1 u1_U342 (.B( u1_L6_1 ) , .Z( u1_N224 ) , .A( u1_out7_1 ) );
  XOR2_X1 u1_U343 (.B( u1_L5_32 ) , .Z( u1_N223 ) , .A( u1_out6_32 ) );
  XOR2_X1 u1_U344 (.B( u1_L5_31 ) , .Z( u1_N222 ) , .A( u1_out6_31 ) );
  XOR2_X1 u1_U351 (.B( u1_L5_25 ) , .Z( u1_N216 ) , .A( u1_out6_25 ) );
  XOR2_X1 u1_U353 (.B( u1_L5_23 ) , .Z( u1_N214 ) , .A( u1_out6_23 ) );
  XOR2_X1 u1_U354 (.B( u1_L5_22 ) , .Z( u1_N213 ) , .A( u1_out6_22 ) );
  XOR2_X1 u1_U36 (.B( u1_L1_6 ) , .Z( u1_N69 ) , .A( u1_out2_6 ) );
  XOR2_X1 u1_U360 (.B( u1_L5_17 ) , .Z( u1_N208 ) , .A( u1_out6_17 ) );
  XOR2_X1 u1_U363 (.B( u1_L5_14 ) , .Z( u1_N205 ) , .A( u1_out6_14 ) );
  XOR2_X1 u1_U365 (.B( u1_L5_12 ) , .Z( u1_N203 ) , .A( u1_out6_12 ) );
  XOR2_X1 u1_U368 (.B( u1_L5_9 ) , .Z( u1_N200 ) , .A( u1_out6_9 ) );
  XOR2_X1 u1_U371 (.B( u1_L5_8 ) , .Z( u1_N199 ) , .A( u1_out6_8 ) );
  XOR2_X1 u1_U372 (.B( u1_L5_7 ) , .Z( u1_N198 ) , .A( u1_out6_7 ) );
  XOR2_X1 u1_U376 (.B( u1_L5_3 ) , .Z( u1_N194 ) , .A( u1_out6_3 ) );
  XOR2_X1 u1_U38 (.B( u1_L1_4 ) , .Z( u1_N67 ) , .A( u1_out2_4 ) );
  XOR2_X1 u1_U416 (.B( u1_L3_31 ) , .Z( u1_N158 ) , .A( u1_out4_31 ) );
  XOR2_X1 u1_U419 (.B( u1_L3_28 ) , .Z( u1_N155 ) , .A( u1_out4_28 ) );
  XOR2_X1 u1_U421 (.B( u1_L3_26 ) , .Z( u1_N153 ) , .A( u1_out4_26 ) );
  XOR2_X1 u1_U424 (.B( u1_L3_23 ) , .Z( u1_N150 ) , .A( u1_out4_23 ) );
  XOR2_X1 u1_U425 (.Z( u1_N15 ) , .B( u1_desIn_r_60 ) , .A( u1_out0_16 ) );
  XOR2_X1 u1_U428 (.B( u1_L3_20 ) , .Z( u1_N147 ) , .A( u1_out4_20 ) );
  XOR2_X1 u1_U430 (.B( u1_L3_18 ) , .Z( u1_N145 ) , .A( u1_out4_18 ) );
  XOR2_X1 u1_U431 (.B( u1_L3_17 ) , .Z( u1_N144 ) , .A( u1_out4_17 ) );
  XOR2_X1 u1_U435 (.B( u1_L3_13 ) , .Z( u1_N140 ) , .A( u1_out4_13 ) );
  XOR2_X1 u1_U439 (.B( u1_L3_10 ) , .Z( u1_N137 ) , .A( u1_out4_10 ) );
  XOR2_X1 u1_U440 (.B( u1_L3_9 ) , .Z( u1_N136 ) , .A( u1_out4_9 ) );
  XOR2_X1 u1_U448 (.B( u1_L3_2 ) , .Z( u1_N129 ) , .A( u1_out4_2 ) );
  XOR2_X1 u1_U449 (.B( u1_L3_1 ) , .Z( u1_N128 ) , .A( u1_out4_1 ) );
  XOR2_X1 u1_U451 (.B( u1_L2_31 ) , .Z( u1_N126 ) , .A( u1_out3_31 ) );
  XOR2_X1 u1_U460 (.B( u1_L2_23 ) , .Z( u1_N118 ) , .A( u1_out3_23 ) );
  XOR2_X1 u1_U466 (.B( u1_L2_17 ) , .Z( u1_N112 ) , .A( u1_out3_17 ) );
  XOR2_X1 u1_U475 (.B( u1_L2_9 ) , .Z( u1_N104 ) , .A( u1_out3_9 ) );
  XOR2_X1 u1_U483 (.Z( u1_FP_9 ) , .B( u1_L14_9 ) , .A( u1_out15_9 ) );
  XOR2_X1 u1_U491 (.Z( u1_FP_31 ) , .B( u1_L14_31 ) , .A( u1_out15_31 ) );
  XOR2_X1 u1_U500 (.Z( u1_FP_23 ) , .B( u1_L14_23 ) , .A( u1_out15_23 ) );
  XOR2_X1 u1_U507 (.Z( u1_FP_17 ) , .B( u1_L14_17 ) , .A( u1_out15_17 ) );
  XOR2_X1 u1_U57 (.Z( u1_N5 ) , .B( u1_desIn_r_46 ) , .A( u1_out0_6 ) );
  XOR2_X1 u1_U67 (.B( u1_L13_25 ) , .Z( u1_N472 ) , .A( u1_out14_25 ) );
  XOR2_X1 u1_U79 (.B( u1_L13_14 ) , .Z( u1_N461 ) , .A( u1_out14_14 ) );
  XOR2_X1 u1_U86 (.B( u1_L13_8 ) , .Z( u1_N455 ) , .A( u1_out14_8 ) );
  XOR2_X1 u1_U9 (.B( u1_L1_30 ) , .Z( u1_N93 ) , .A( u1_out2_30 ) );
  XOR2_X1 u1_U91 (.B( u1_L13_3 ) , .Z( u1_N450 ) , .A( u1_out14_3 ) );
  XOR2_X1 u1_U98 (.B( u1_L12_29 ) , .Z( u1_N444 ) , .A( u1_out13_29 ) );
  XOR2_X1 u1_u0_U42 (.B( u1_K1_16 ) , .A( u1_desIn_r_21 ) , .Z( u1_u0_X_16 ) );
  XOR2_X1 u1_u0_U43 (.B( u1_K1_15 ) , .A( u1_desIn_r_13 ) , .Z( u1_u0_X_15 ) );
  OAI22_X1 u1_u0_u2_U10 (.B1( u1_u0_u2_n151 ) , .A2( u1_u0_u2_n152 ) , .A1( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n160 ) , .B2( u1_u0_u2_n168 ) );
  NAND3_X1 u1_u0_u2_U100 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n104 ) , .A3( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n98 ) );
  NOR3_X1 u1_u0_u2_U11 (.A1( u1_u0_u2_n150 ) , .ZN( u1_u0_u2_n151 ) , .A3( u1_u0_u2_n175 ) , .A2( u1_u0_u2_n188 ) );
  AOI21_X1 u1_u0_u2_U12 (.B2( u1_u0_u2_n123 ) , .ZN( u1_u0_u2_n125 ) , .A( u1_u0_u2_n171 ) , .B1( u1_u0_u2_n184 ) );
  INV_X1 u1_u0_u2_U13 (.A( u1_u0_u2_n150 ) , .ZN( u1_u0_u2_n184 ) );
  AOI21_X1 u1_u0_u2_U14 (.ZN( u1_u0_u2_n144 ) , .B2( u1_u0_u2_n155 ) , .A( u1_u0_u2_n172 ) , .B1( u1_u0_u2_n185 ) );
  AOI21_X1 u1_u0_u2_U15 (.B2( u1_u0_u2_n143 ) , .ZN( u1_u0_u2_n145 ) , .B1( u1_u0_u2_n152 ) , .A( u1_u0_u2_n171 ) );
  INV_X1 u1_u0_u2_U16 (.A( u1_u0_u2_n156 ) , .ZN( u1_u0_u2_n171 ) );
  INV_X1 u1_u0_u2_U17 (.A( u1_u0_u2_n120 ) , .ZN( u1_u0_u2_n188 ) );
  NAND2_X1 u1_u0_u2_U18 (.A2( u1_u0_u2_n122 ) , .ZN( u1_u0_u2_n150 ) , .A1( u1_u0_u2_n152 ) );
  INV_X1 u1_u0_u2_U19 (.A( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n170 ) );
  INV_X1 u1_u0_u2_U20 (.A( u1_u0_u2_n137 ) , .ZN( u1_u0_u2_n173 ) );
  NAND2_X1 u1_u0_u2_U21 (.A1( u1_u0_u2_n132 ) , .A2( u1_u0_u2_n139 ) , .ZN( u1_u0_u2_n157 ) );
  INV_X1 u1_u0_u2_U22 (.A( u1_u0_u2_n113 ) , .ZN( u1_u0_u2_n178 ) );
  INV_X1 u1_u0_u2_U23 (.A( u1_u0_u2_n139 ) , .ZN( u1_u0_u2_n175 ) );
  INV_X1 u1_u0_u2_U24 (.A( u1_u0_u2_n155 ) , .ZN( u1_u0_u2_n181 ) );
  INV_X1 u1_u0_u2_U25 (.A( u1_u0_u2_n119 ) , .ZN( u1_u0_u2_n177 ) );
  INV_X1 u1_u0_u2_U26 (.A( u1_u0_u2_n116 ) , .ZN( u1_u0_u2_n180 ) );
  INV_X1 u1_u0_u2_U27 (.A( u1_u0_u2_n131 ) , .ZN( u1_u0_u2_n179 ) );
  INV_X1 u1_u0_u2_U28 (.A( u1_u0_u2_n154 ) , .ZN( u1_u0_u2_n176 ) );
  NAND2_X1 u1_u0_u2_U29 (.A2( u1_u0_u2_n116 ) , .A1( u1_u0_u2_n117 ) , .ZN( u1_u0_u2_n118 ) );
  NOR2_X1 u1_u0_u2_U3 (.ZN( u1_u0_u2_n121 ) , .A2( u1_u0_u2_n177 ) , .A1( u1_u0_u2_n180 ) );
  INV_X1 u1_u0_u2_U30 (.A( u1_u0_u2_n132 ) , .ZN( u1_u0_u2_n182 ) );
  INV_X1 u1_u0_u2_U31 (.A( u1_u0_u2_n158 ) , .ZN( u1_u0_u2_n183 ) );
  OAI21_X1 u1_u0_u2_U32 (.A( u1_u0_u2_n156 ) , .B1( u1_u0_u2_n157 ) , .ZN( u1_u0_u2_n158 ) , .B2( u1_u0_u2_n179 ) );
  NOR2_X1 u1_u0_u2_U33 (.ZN( u1_u0_u2_n156 ) , .A1( u1_u0_u2_n166 ) , .A2( u1_u0_u2_n169 ) );
  NOR2_X1 u1_u0_u2_U34 (.A2( u1_u0_u2_n114 ) , .ZN( u1_u0_u2_n137 ) , .A1( u1_u0_u2_n140 ) );
  NOR2_X1 u1_u0_u2_U35 (.A2( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n153 ) , .A1( u1_u0_u2_n156 ) );
  AOI211_X1 u1_u0_u2_U36 (.ZN( u1_u0_u2_n130 ) , .C1( u1_u0_u2_n138 ) , .C2( u1_u0_u2_n179 ) , .B( u1_u0_u2_n96 ) , .A( u1_u0_u2_n97 ) );
  OAI22_X1 u1_u0_u2_U37 (.B1( u1_u0_u2_n133 ) , .A2( u1_u0_u2_n137 ) , .A1( u1_u0_u2_n152 ) , .B2( u1_u0_u2_n168 ) , .ZN( u1_u0_u2_n97 ) );
  OAI221_X1 u1_u0_u2_U38 (.B1( u1_u0_u2_n113 ) , .C1( u1_u0_u2_n132 ) , .A( u1_u0_u2_n149 ) , .B2( u1_u0_u2_n171 ) , .C2( u1_u0_u2_n172 ) , .ZN( u1_u0_u2_n96 ) );
  OAI221_X1 u1_u0_u2_U39 (.A( u1_u0_u2_n115 ) , .C2( u1_u0_u2_n123 ) , .B2( u1_u0_u2_n143 ) , .B1( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n163 ) , .C1( u1_u0_u2_n168 ) );
  INV_X1 u1_u0_u2_U4 (.A( u1_u0_u2_n134 ) , .ZN( u1_u0_u2_n185 ) );
  OAI21_X1 u1_u0_u2_U40 (.A( u1_u0_u2_n114 ) , .ZN( u1_u0_u2_n115 ) , .B1( u1_u0_u2_n176 ) , .B2( u1_u0_u2_n178 ) );
  OAI221_X1 u1_u0_u2_U41 (.A( u1_u0_u2_n135 ) , .B2( u1_u0_u2_n136 ) , .B1( u1_u0_u2_n137 ) , .ZN( u1_u0_u2_n162 ) , .C2( u1_u0_u2_n167 ) , .C1( u1_u0_u2_n185 ) );
  AND3_X1 u1_u0_u2_U42 (.A3( u1_u0_u2_n131 ) , .A2( u1_u0_u2_n132 ) , .A1( u1_u0_u2_n133 ) , .ZN( u1_u0_u2_n136 ) );
  AOI22_X1 u1_u0_u2_U43 (.ZN( u1_u0_u2_n135 ) , .B1( u1_u0_u2_n140 ) , .A1( u1_u0_u2_n156 ) , .B2( u1_u0_u2_n180 ) , .A2( u1_u0_u2_n188 ) );
  AOI21_X1 u1_u0_u2_U44 (.ZN( u1_u0_u2_n149 ) , .B1( u1_u0_u2_n173 ) , .B2( u1_u0_u2_n188 ) , .A( u1_u0_u2_n95 ) );
  AND3_X1 u1_u0_u2_U45 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n104 ) , .A3( u1_u0_u2_n156 ) , .ZN( u1_u0_u2_n95 ) );
  OAI21_X1 u1_u0_u2_U46 (.A( u1_u0_u2_n101 ) , .B2( u1_u0_u2_n121 ) , .B1( u1_u0_u2_n153 ) , .ZN( u1_u0_u2_n164 ) );
  NAND2_X1 u1_u0_u2_U47 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n107 ) , .ZN( u1_u0_u2_n155 ) );
  NAND2_X1 u1_u0_u2_U48 (.A2( u1_u0_u2_n105 ) , .A1( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n143 ) );
  NAND2_X1 u1_u0_u2_U49 (.A1( u1_u0_u2_n104 ) , .A2( u1_u0_u2_n106 ) , .ZN( u1_u0_u2_n152 ) );
  NOR4_X1 u1_u0_u2_U5 (.A4( u1_u0_u2_n124 ) , .A3( u1_u0_u2_n125 ) , .A2( u1_u0_u2_n126 ) , .A1( u1_u0_u2_n127 ) , .ZN( u1_u0_u2_n128 ) );
  NAND2_X1 u1_u0_u2_U50 (.A1( u1_u0_u2_n100 ) , .A2( u1_u0_u2_n105 ) , .ZN( u1_u0_u2_n132 ) );
  INV_X1 u1_u0_u2_U51 (.A( u1_u0_u2_n140 ) , .ZN( u1_u0_u2_n168 ) );
  INV_X1 u1_u0_u2_U52 (.A( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n167 ) );
  OAI21_X1 u1_u0_u2_U53 (.A( u1_u0_u2_n141 ) , .B2( u1_u0_u2_n142 ) , .ZN( u1_u0_u2_n146 ) , .B1( u1_u0_u2_n153 ) );
  OAI21_X1 u1_u0_u2_U54 (.A( u1_u0_u2_n140 ) , .ZN( u1_u0_u2_n141 ) , .B1( u1_u0_u2_n176 ) , .B2( u1_u0_u2_n177 ) );
  NOR3_X1 u1_u0_u2_U55 (.ZN( u1_u0_u2_n142 ) , .A3( u1_u0_u2_n175 ) , .A2( u1_u0_u2_n178 ) , .A1( u1_u0_u2_n181 ) );
  NAND2_X1 u1_u0_u2_U56 (.A1( u1_u0_u2_n102 ) , .A2( u1_u0_u2_n106 ) , .ZN( u1_u0_u2_n113 ) );
  NAND2_X1 u1_u0_u2_U57 (.A1( u1_u0_u2_n106 ) , .A2( u1_u0_u2_n107 ) , .ZN( u1_u0_u2_n131 ) );
  NAND2_X1 u1_u0_u2_U58 (.A1( u1_u0_u2_n103 ) , .A2( u1_u0_u2_n107 ) , .ZN( u1_u0_u2_n139 ) );
  NAND2_X1 u1_u0_u2_U59 (.A1( u1_u0_u2_n103 ) , .A2( u1_u0_u2_n105 ) , .ZN( u1_u0_u2_n133 ) );
  AOI21_X1 u1_u0_u2_U6 (.B2( u1_u0_u2_n119 ) , .ZN( u1_u0_u2_n127 ) , .A( u1_u0_u2_n137 ) , .B1( u1_u0_u2_n155 ) );
  NAND2_X1 u1_u0_u2_U60 (.A1( u1_u0_u2_n102 ) , .A2( u1_u0_u2_n103 ) , .ZN( u1_u0_u2_n154 ) );
  NAND2_X1 u1_u0_u2_U61 (.A2( u1_u0_u2_n103 ) , .A1( u1_u0_u2_n104 ) , .ZN( u1_u0_u2_n119 ) );
  NAND2_X1 u1_u0_u2_U62 (.A2( u1_u0_u2_n107 ) , .A1( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n123 ) );
  NAND2_X1 u1_u0_u2_U63 (.A1( u1_u0_u2_n104 ) , .A2( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n122 ) );
  INV_X1 u1_u0_u2_U64 (.A( u1_u0_u2_n114 ) , .ZN( u1_u0_u2_n172 ) );
  NAND2_X1 u1_u0_u2_U65 (.A2( u1_u0_u2_n100 ) , .A1( u1_u0_u2_n102 ) , .ZN( u1_u0_u2_n116 ) );
  NAND2_X1 u1_u0_u2_U66 (.A1( u1_u0_u2_n102 ) , .A2( u1_u0_u2_n108 ) , .ZN( u1_u0_u2_n120 ) );
  NAND2_X1 u1_u0_u2_U67 (.A2( u1_u0_u2_n105 ) , .A1( u1_u0_u2_n106 ) , .ZN( u1_u0_u2_n117 ) );
  INV_X1 u1_u0_u2_U68 (.ZN( u1_u0_u2_n187 ) , .A( u1_u0_u2_n99 ) );
  OAI21_X1 u1_u0_u2_U69 (.B1( u1_u0_u2_n137 ) , .B2( u1_u0_u2_n143 ) , .A( u1_u0_u2_n98 ) , .ZN( u1_u0_u2_n99 ) );
  AOI21_X1 u1_u0_u2_U7 (.ZN( u1_u0_u2_n124 ) , .B1( u1_u0_u2_n131 ) , .B2( u1_u0_u2_n143 ) , .A( u1_u0_u2_n172 ) );
  NOR2_X1 u1_u0_u2_U70 (.A2( u1_u0_X_16 ) , .ZN( u1_u0_u2_n140 ) , .A1( u1_u0_u2_n166 ) );
  NOR2_X1 u1_u0_u2_U71 (.A2( u1_u0_X_13 ) , .A1( u1_u0_X_14 ) , .ZN( u1_u0_u2_n100 ) );
  NOR2_X1 u1_u0_u2_U72 (.A2( u1_u0_X_16 ) , .A1( u1_u0_X_17 ) , .ZN( u1_u0_u2_n138 ) );
  NOR2_X1 u1_u0_u2_U73 (.A2( u1_u0_X_15 ) , .A1( u1_u0_X_18 ) , .ZN( u1_u0_u2_n104 ) );
  NOR2_X1 u1_u0_u2_U74 (.A2( u1_u0_X_14 ) , .ZN( u1_u0_u2_n103 ) , .A1( u1_u0_u2_n174 ) );
  NOR2_X1 u1_u0_u2_U75 (.A2( u1_u0_X_15 ) , .ZN( u1_u0_u2_n102 ) , .A1( u1_u0_u2_n165 ) );
  NOR2_X1 u1_u0_u2_U76 (.A2( u1_u0_X_17 ) , .ZN( u1_u0_u2_n114 ) , .A1( u1_u0_u2_n169 ) );
  AND2_X1 u1_u0_u2_U77 (.A1( u1_u0_X_15 ) , .ZN( u1_u0_u2_n105 ) , .A2( u1_u0_u2_n165 ) );
  AND2_X1 u1_u0_u2_U78 (.A2( u1_u0_X_15 ) , .A1( u1_u0_X_18 ) , .ZN( u1_u0_u2_n107 ) );
  AND2_X1 u1_u0_u2_U79 (.A1( u1_u0_X_14 ) , .ZN( u1_u0_u2_n106 ) , .A2( u1_u0_u2_n174 ) );
  AOI21_X1 u1_u0_u2_U8 (.B2( u1_u0_u2_n120 ) , .B1( u1_u0_u2_n121 ) , .ZN( u1_u0_u2_n126 ) , .A( u1_u0_u2_n167 ) );
  AND2_X1 u1_u0_u2_U80 (.A1( u1_u0_X_13 ) , .A2( u1_u0_X_14 ) , .ZN( u1_u0_u2_n108 ) );
  INV_X1 u1_u0_u2_U81 (.A( u1_u0_X_16 ) , .ZN( u1_u0_u2_n169 ) );
  INV_X1 u1_u0_u2_U82 (.A( u1_u0_X_17 ) , .ZN( u1_u0_u2_n166 ) );
  INV_X1 u1_u0_u2_U83 (.A( u1_u0_X_13 ) , .ZN( u1_u0_u2_n174 ) );
  INV_X1 u1_u0_u2_U84 (.A( u1_u0_X_18 ) , .ZN( u1_u0_u2_n165 ) );
  NAND4_X1 u1_u0_u2_U85 (.ZN( u1_out0_30 ) , .A4( u1_u0_u2_n147 ) , .A3( u1_u0_u2_n148 ) , .A2( u1_u0_u2_n149 ) , .A1( u1_u0_u2_n187 ) );
  NOR3_X1 u1_u0_u2_U86 (.A3( u1_u0_u2_n144 ) , .A2( u1_u0_u2_n145 ) , .A1( u1_u0_u2_n146 ) , .ZN( u1_u0_u2_n147 ) );
  AOI21_X1 u1_u0_u2_U87 (.B2( u1_u0_u2_n138 ) , .ZN( u1_u0_u2_n148 ) , .A( u1_u0_u2_n162 ) , .B1( u1_u0_u2_n182 ) );
  NAND4_X1 u1_u0_u2_U88 (.ZN( u1_out0_24 ) , .A4( u1_u0_u2_n111 ) , .A3( u1_u0_u2_n112 ) , .A1( u1_u0_u2_n130 ) , .A2( u1_u0_u2_n187 ) );
  AOI221_X1 u1_u0_u2_U89 (.A( u1_u0_u2_n109 ) , .B1( u1_u0_u2_n110 ) , .ZN( u1_u0_u2_n111 ) , .C1( u1_u0_u2_n134 ) , .C2( u1_u0_u2_n170 ) , .B2( u1_u0_u2_n173 ) );
  OAI22_X1 u1_u0_u2_U9 (.ZN( u1_u0_u2_n109 ) , .A2( u1_u0_u2_n113 ) , .B2( u1_u0_u2_n133 ) , .B1( u1_u0_u2_n167 ) , .A1( u1_u0_u2_n168 ) );
  AOI21_X1 u1_u0_u2_U90 (.ZN( u1_u0_u2_n112 ) , .B2( u1_u0_u2_n156 ) , .A( u1_u0_u2_n164 ) , .B1( u1_u0_u2_n181 ) );
  NAND4_X1 u1_u0_u2_U91 (.ZN( u1_out0_16 ) , .A4( u1_u0_u2_n128 ) , .A3( u1_u0_u2_n129 ) , .A1( u1_u0_u2_n130 ) , .A2( u1_u0_u2_n186 ) );
  AOI22_X1 u1_u0_u2_U92 (.A2( u1_u0_u2_n118 ) , .ZN( u1_u0_u2_n129 ) , .A1( u1_u0_u2_n140 ) , .B1( u1_u0_u2_n157 ) , .B2( u1_u0_u2_n170 ) );
  INV_X1 u1_u0_u2_U93 (.A( u1_u0_u2_n163 ) , .ZN( u1_u0_u2_n186 ) );
  OR4_X1 u1_u0_u2_U94 (.ZN( u1_out0_6 ) , .A4( u1_u0_u2_n161 ) , .A3( u1_u0_u2_n162 ) , .A2( u1_u0_u2_n163 ) , .A1( u1_u0_u2_n164 ) );
  OR3_X1 u1_u0_u2_U95 (.A2( u1_u0_u2_n159 ) , .A1( u1_u0_u2_n160 ) , .ZN( u1_u0_u2_n161 ) , .A3( u1_u0_u2_n183 ) );
  AOI21_X1 u1_u0_u2_U96 (.B2( u1_u0_u2_n154 ) , .B1( u1_u0_u2_n155 ) , .ZN( u1_u0_u2_n159 ) , .A( u1_u0_u2_n167 ) );
  NAND3_X1 u1_u0_u2_U97 (.A2( u1_u0_u2_n117 ) , .A1( u1_u0_u2_n122 ) , .A3( u1_u0_u2_n123 ) , .ZN( u1_u0_u2_n134 ) );
  NAND3_X1 u1_u0_u2_U98 (.ZN( u1_u0_u2_n110 ) , .A2( u1_u0_u2_n131 ) , .A3( u1_u0_u2_n139 ) , .A1( u1_u0_u2_n154 ) );
  NAND3_X1 u1_u0_u2_U99 (.A2( u1_u0_u2_n100 ) , .ZN( u1_u0_u2_n101 ) , .A1( u1_u0_u2_n104 ) , .A3( u1_u0_u2_n114 ) );
  XOR2_X1 u1_u10_U1 (.B( u1_K11_9 ) , .A( u1_R9_6 ) , .Z( u1_u10_X_9 ) );
  XOR2_X1 u1_u10_U16 (.B( u1_K11_3 ) , .A( u1_R9_2 ) , .Z( u1_u10_X_3 ) );
  XOR2_X1 u1_u10_U2 (.B( u1_K11_8 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_8 ) );
  XOR2_X1 u1_u10_U22 (.B( u1_K11_34 ) , .A( u1_R9_23 ) , .Z( u1_u10_X_34 ) );
  XOR2_X1 u1_u10_U23 (.B( u1_K11_33 ) , .A( u1_R9_22 ) , .Z( u1_u10_X_33 ) );
  XOR2_X1 u1_u10_U24 (.B( u1_K11_32 ) , .A( u1_R9_21 ) , .Z( u1_u10_X_32 ) );
  XOR2_X1 u1_u10_U25 (.B( u1_K11_31 ) , .A( u1_R9_20 ) , .Z( u1_u10_X_31 ) );
  XOR2_X1 u1_u10_U26 (.B( u1_K11_30 ) , .A( u1_R9_21 ) , .Z( u1_u10_X_30 ) );
  XOR2_X1 u1_u10_U28 (.B( u1_K11_29 ) , .A( u1_R9_20 ) , .Z( u1_u10_X_29 ) );
  XOR2_X1 u1_u10_U29 (.B( u1_K11_28 ) , .A( u1_R9_19 ) , .Z( u1_u10_X_28 ) );
  XOR2_X1 u1_u10_U3 (.B( u1_K11_7 ) , .A( u1_R9_4 ) , .Z( u1_u10_X_7 ) );
  XOR2_X1 u1_u10_U30 (.B( u1_K11_27 ) , .A( u1_R9_18 ) , .Z( u1_u10_X_27 ) );
  XOR2_X1 u1_u10_U4 (.B( u1_K11_6 ) , .A( u1_R9_5 ) , .Z( u1_u10_X_6 ) );
  XOR2_X1 u1_u10_U48 (.B( u1_K11_10 ) , .A( u1_R9_7 ) , .Z( u1_u10_X_10 ) );
  XOR2_X1 u1_u10_U5 (.B( u1_K11_5 ) , .A( u1_R9_4 ) , .Z( u1_u10_X_5 ) );
  XOR2_X1 u1_u10_U6 (.B( u1_K11_4 ) , .A( u1_R9_3 ) , .Z( u1_u10_X_4 ) );
  AND3_X1 u1_u10_u0_U10 (.A2( u1_u10_u0_n112 ) , .ZN( u1_u10_u0_n127 ) , .A3( u1_u10_u0_n130 ) , .A1( u1_u10_u0_n148 ) );
  NAND2_X1 u1_u10_u0_U11 (.ZN( u1_u10_u0_n113 ) , .A1( u1_u10_u0_n139 ) , .A2( u1_u10_u0_n149 ) );
  AND2_X1 u1_u10_u0_U12 (.ZN( u1_u10_u0_n107 ) , .A1( u1_u10_u0_n130 ) , .A2( u1_u10_u0_n140 ) );
  AND2_X1 u1_u10_u0_U13 (.A2( u1_u10_u0_n129 ) , .A1( u1_u10_u0_n130 ) , .ZN( u1_u10_u0_n151 ) );
  AND2_X1 u1_u10_u0_U14 (.A1( u1_u10_u0_n108 ) , .A2( u1_u10_u0_n125 ) , .ZN( u1_u10_u0_n145 ) );
  INV_X1 u1_u10_u0_U15 (.A( u1_u10_u0_n143 ) , .ZN( u1_u10_u0_n173 ) );
  NOR2_X1 u1_u10_u0_U16 (.A2( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n147 ) , .A1( u1_u10_u0_n160 ) );
  NOR2_X1 u1_u10_u0_U17 (.A1( u1_u10_u0_n163 ) , .A2( u1_u10_u0_n164 ) , .ZN( u1_u10_u0_n95 ) );
  AOI21_X1 u1_u10_u0_U18 (.B1( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n132 ) , .A( u1_u10_u0_n165 ) , .B2( u1_u10_u0_n93 ) );
  INV_X1 u1_u10_u0_U19 (.A( u1_u10_u0_n142 ) , .ZN( u1_u10_u0_n165 ) );
  OAI221_X1 u1_u10_u0_U20 (.C1( u1_u10_u0_n121 ) , .ZN( u1_u10_u0_n122 ) , .B2( u1_u10_u0_n127 ) , .A( u1_u10_u0_n143 ) , .B1( u1_u10_u0_n144 ) , .C2( u1_u10_u0_n147 ) );
  OAI22_X1 u1_u10_u0_U21 (.B1( u1_u10_u0_n125 ) , .ZN( u1_u10_u0_n126 ) , .A1( u1_u10_u0_n138 ) , .A2( u1_u10_u0_n146 ) , .B2( u1_u10_u0_n147 ) );
  OAI22_X1 u1_u10_u0_U22 (.B1( u1_u10_u0_n131 ) , .A1( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n147 ) , .A2( u1_u10_u0_n90 ) , .ZN( u1_u10_u0_n91 ) );
  AND3_X1 u1_u10_u0_U23 (.A3( u1_u10_u0_n121 ) , .A2( u1_u10_u0_n125 ) , .A1( u1_u10_u0_n148 ) , .ZN( u1_u10_u0_n90 ) );
  INV_X1 u1_u10_u0_U24 (.A( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n161 ) );
  NOR2_X1 u1_u10_u0_U25 (.A1( u1_u10_u0_n120 ) , .ZN( u1_u10_u0_n143 ) , .A2( u1_u10_u0_n167 ) );
  OAI221_X1 u1_u10_u0_U26 (.C1( u1_u10_u0_n112 ) , .ZN( u1_u10_u0_n120 ) , .B1( u1_u10_u0_n138 ) , .B2( u1_u10_u0_n141 ) , .C2( u1_u10_u0_n147 ) , .A( u1_u10_u0_n172 ) );
  AOI22_X1 u1_u10_u0_U27 (.B2( u1_u10_u0_n109 ) , .A2( u1_u10_u0_n110 ) , .ZN( u1_u10_u0_n111 ) , .B1( u1_u10_u0_n118 ) , .A1( u1_u10_u0_n160 ) );
  INV_X1 u1_u10_u0_U28 (.A( u1_u10_u0_n118 ) , .ZN( u1_u10_u0_n158 ) );
  AOI21_X1 u1_u10_u0_U29 (.B1( u1_u10_u0_n132 ) , .ZN( u1_u10_u0_n133 ) , .A( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n166 ) );
  INV_X1 u1_u10_u0_U3 (.A( u1_u10_u0_n113 ) , .ZN( u1_u10_u0_n166 ) );
  AOI21_X1 u1_u10_u0_U30 (.ZN( u1_u10_u0_n104 ) , .B1( u1_u10_u0_n107 ) , .B2( u1_u10_u0_n141 ) , .A( u1_u10_u0_n144 ) );
  AOI21_X1 u1_u10_u0_U31 (.B1( u1_u10_u0_n127 ) , .B2( u1_u10_u0_n129 ) , .A( u1_u10_u0_n138 ) , .ZN( u1_u10_u0_n96 ) );
  AOI21_X1 u1_u10_u0_U32 (.ZN( u1_u10_u0_n116 ) , .B2( u1_u10_u0_n142 ) , .A( u1_u10_u0_n144 ) , .B1( u1_u10_u0_n166 ) );
  NAND2_X1 u1_u10_u0_U33 (.A1( u1_u10_u0_n100 ) , .A2( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n125 ) );
  NAND2_X1 u1_u10_u0_U34 (.A2( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n140 ) , .A1( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U35 (.A1( u1_u10_u0_n101 ) , .A2( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n150 ) );
  INV_X1 u1_u10_u0_U36 (.A( u1_u10_u0_n138 ) , .ZN( u1_u10_u0_n160 ) );
  NAND2_X1 u1_u10_u0_U37 (.ZN( u1_u10_u0_n142 ) , .A1( u1_u10_u0_n94 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U38 (.A1( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n128 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U39 (.A2( u1_u10_u0_n102 ) , .A1( u1_u10_u0_n103 ) , .ZN( u1_u10_u0_n149 ) );
  AOI21_X1 u1_u10_u0_U4 (.B2( u1_u10_u0_n131 ) , .ZN( u1_u10_u0_n134 ) , .B1( u1_u10_u0_n151 ) , .A( u1_u10_u0_n158 ) );
  NAND2_X1 u1_u10_u0_U40 (.A1( u1_u10_u0_n100 ) , .ZN( u1_u10_u0_n129 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U41 (.A2( u1_u10_u0_n100 ) , .A1( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n139 ) );
  NAND2_X1 u1_u10_u0_U42 (.A2( u1_u10_u0_n100 ) , .ZN( u1_u10_u0_n131 ) , .A1( u1_u10_u0_n92 ) );
  NAND2_X1 u1_u10_u0_U43 (.ZN( u1_u10_u0_n108 ) , .A1( u1_u10_u0_n92 ) , .A2( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U44 (.ZN( u1_u10_u0_n148 ) , .A1( u1_u10_u0_n93 ) , .A2( u1_u10_u0_n95 ) );
  NAND2_X1 u1_u10_u0_U45 (.A2( u1_u10_u0_n102 ) , .ZN( u1_u10_u0_n114 ) , .A1( u1_u10_u0_n92 ) );
  NAND2_X1 u1_u10_u0_U46 (.A1( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n130 ) , .A2( u1_u10_u0_n94 ) );
  NAND2_X1 u1_u10_u0_U47 (.A2( u1_u10_u0_n101 ) , .ZN( u1_u10_u0_n121 ) , .A1( u1_u10_u0_n93 ) );
  INV_X1 u1_u10_u0_U48 (.ZN( u1_u10_u0_n172 ) , .A( u1_u10_u0_n88 ) );
  OAI222_X1 u1_u10_u0_U49 (.C1( u1_u10_u0_n108 ) , .A1( u1_u10_u0_n125 ) , .B2( u1_u10_u0_n128 ) , .B1( u1_u10_u0_n144 ) , .A2( u1_u10_u0_n158 ) , .C2( u1_u10_u0_n161 ) , .ZN( u1_u10_u0_n88 ) );
  NOR2_X1 u1_u10_u0_U5 (.A1( u1_u10_u0_n108 ) , .ZN( u1_u10_u0_n123 ) , .A2( u1_u10_u0_n158 ) );
  NAND2_X1 u1_u10_u0_U50 (.ZN( u1_u10_u0_n112 ) , .A2( u1_u10_u0_n92 ) , .A1( u1_u10_u0_n93 ) );
  OR3_X1 u1_u10_u0_U51 (.A3( u1_u10_u0_n152 ) , .A2( u1_u10_u0_n153 ) , .A1( u1_u10_u0_n154 ) , .ZN( u1_u10_u0_n155 ) );
  AOI21_X1 u1_u10_u0_U52 (.A( u1_u10_u0_n144 ) , .B2( u1_u10_u0_n145 ) , .B1( u1_u10_u0_n146 ) , .ZN( u1_u10_u0_n154 ) );
  AOI21_X1 u1_u10_u0_U53 (.B2( u1_u10_u0_n150 ) , .B1( u1_u10_u0_n151 ) , .ZN( u1_u10_u0_n152 ) , .A( u1_u10_u0_n158 ) );
  AOI21_X1 u1_u10_u0_U54 (.A( u1_u10_u0_n147 ) , .B2( u1_u10_u0_n148 ) , .B1( u1_u10_u0_n149 ) , .ZN( u1_u10_u0_n153 ) );
  INV_X1 u1_u10_u0_U55 (.ZN( u1_u10_u0_n171 ) , .A( u1_u10_u0_n99 ) );
  OAI211_X1 u1_u10_u0_U56 (.C2( u1_u10_u0_n140 ) , .C1( u1_u10_u0_n161 ) , .A( u1_u10_u0_n169 ) , .B( u1_u10_u0_n98 ) , .ZN( u1_u10_u0_n99 ) );
  INV_X1 u1_u10_u0_U57 (.ZN( u1_u10_u0_n169 ) , .A( u1_u10_u0_n91 ) );
  AOI211_X1 u1_u10_u0_U58 (.C1( u1_u10_u0_n118 ) , .A( u1_u10_u0_n123 ) , .B( u1_u10_u0_n96 ) , .C2( u1_u10_u0_n97 ) , .ZN( u1_u10_u0_n98 ) );
  NOR2_X1 u1_u10_u0_U59 (.A2( u1_u10_X_2 ) , .ZN( u1_u10_u0_n103 ) , .A1( u1_u10_u0_n164 ) );
  OAI21_X1 u1_u10_u0_U6 (.B1( u1_u10_u0_n150 ) , .B2( u1_u10_u0_n158 ) , .A( u1_u10_u0_n172 ) , .ZN( u1_u10_u0_n89 ) );
  NOR2_X1 u1_u10_u0_U60 (.A2( u1_u10_X_3 ) , .A1( u1_u10_X_6 ) , .ZN( u1_u10_u0_n94 ) );
  NOR2_X1 u1_u10_u0_U61 (.A2( u1_u10_X_6 ) , .ZN( u1_u10_u0_n100 ) , .A1( u1_u10_u0_n162 ) );
  NOR2_X1 u1_u10_u0_U62 (.A2( u1_u10_X_1 ) , .A1( u1_u10_X_2 ) , .ZN( u1_u10_u0_n92 ) );
  NOR2_X1 u1_u10_u0_U63 (.A2( u1_u10_X_1 ) , .ZN( u1_u10_u0_n101 ) , .A1( u1_u10_u0_n163 ) );
  NOR2_X1 u1_u10_u0_U64 (.A2( u1_u10_X_4 ) , .A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n118 ) );
  NAND2_X1 u1_u10_u0_U65 (.A2( u1_u10_X_4 ) , .A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n144 ) );
  NOR2_X1 u1_u10_u0_U66 (.A2( u1_u10_X_5 ) , .ZN( u1_u10_u0_n136 ) , .A1( u1_u10_u0_n159 ) );
  NAND2_X1 u1_u10_u0_U67 (.A1( u1_u10_X_5 ) , .ZN( u1_u10_u0_n138 ) , .A2( u1_u10_u0_n159 ) );
  AND2_X1 u1_u10_u0_U68 (.A2( u1_u10_X_3 ) , .A1( u1_u10_X_6 ) , .ZN( u1_u10_u0_n102 ) );
  AND2_X1 u1_u10_u0_U69 (.A1( u1_u10_X_6 ) , .A2( u1_u10_u0_n162 ) , .ZN( u1_u10_u0_n93 ) );
  AOI21_X1 u1_u10_u0_U7 (.B1( u1_u10_u0_n114 ) , .ZN( u1_u10_u0_n115 ) , .B2( u1_u10_u0_n129 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U70 (.A( u1_u10_X_4 ) , .ZN( u1_u10_u0_n159 ) );
  INV_X1 u1_u10_u0_U71 (.A( u1_u10_X_1 ) , .ZN( u1_u10_u0_n164 ) );
  INV_X1 u1_u10_u0_U72 (.A( u1_u10_X_2 ) , .ZN( u1_u10_u0_n163 ) );
  INV_X1 u1_u10_u0_U73 (.A( u1_u10_X_3 ) , .ZN( u1_u10_u0_n162 ) );
  INV_X1 u1_u10_u0_U74 (.ZN( u1_u10_u0_n174 ) , .A( u1_u10_u0_n89 ) );
  AOI211_X1 u1_u10_u0_U75 (.B( u1_u10_u0_n104 ) , .A( u1_u10_u0_n105 ) , .ZN( u1_u10_u0_n106 ) , .C2( u1_u10_u0_n113 ) , .C1( u1_u10_u0_n160 ) );
  OR4_X1 u1_u10_u0_U76 (.ZN( u1_out10_17 ) , .A4( u1_u10_u0_n122 ) , .A2( u1_u10_u0_n123 ) , .A1( u1_u10_u0_n124 ) , .A3( u1_u10_u0_n170 ) );
  AOI21_X1 u1_u10_u0_U77 (.B2( u1_u10_u0_n107 ) , .ZN( u1_u10_u0_n124 ) , .B1( u1_u10_u0_n128 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U78 (.A( u1_u10_u0_n111 ) , .ZN( u1_u10_u0_n170 ) );
  OR4_X1 u1_u10_u0_U79 (.ZN( u1_out10_31 ) , .A4( u1_u10_u0_n155 ) , .A2( u1_u10_u0_n156 ) , .A1( u1_u10_u0_n157 ) , .A3( u1_u10_u0_n173 ) );
  AND2_X1 u1_u10_u0_U8 (.A1( u1_u10_u0_n114 ) , .A2( u1_u10_u0_n121 ) , .ZN( u1_u10_u0_n146 ) );
  AOI21_X1 u1_u10_u0_U80 (.A( u1_u10_u0_n138 ) , .B2( u1_u10_u0_n139 ) , .B1( u1_u10_u0_n140 ) , .ZN( u1_u10_u0_n157 ) );
  AOI21_X1 u1_u10_u0_U81 (.B2( u1_u10_u0_n141 ) , .B1( u1_u10_u0_n142 ) , .ZN( u1_u10_u0_n156 ) , .A( u1_u10_u0_n161 ) );
  INV_X1 u1_u10_u0_U82 (.A( u1_u10_u0_n126 ) , .ZN( u1_u10_u0_n168 ) );
  AOI211_X1 u1_u10_u0_U83 (.B( u1_u10_u0_n133 ) , .A( u1_u10_u0_n134 ) , .C2( u1_u10_u0_n135 ) , .C1( u1_u10_u0_n136 ) , .ZN( u1_u10_u0_n137 ) );
  AOI211_X1 u1_u10_u0_U84 (.B( u1_u10_u0_n115 ) , .A( u1_u10_u0_n116 ) , .C2( u1_u10_u0_n117 ) , .C1( u1_u10_u0_n118 ) , .ZN( u1_u10_u0_n119 ) );
  INV_X1 u1_u10_u0_U85 (.A( u1_u10_u0_n119 ) , .ZN( u1_u10_u0_n167 ) );
  NAND2_X1 u1_u10_u0_U86 (.ZN( u1_u10_u0_n110 ) , .A2( u1_u10_u0_n132 ) , .A1( u1_u10_u0_n145 ) );
  OAI22_X1 u1_u10_u0_U87 (.ZN( u1_u10_u0_n105 ) , .A2( u1_u10_u0_n132 ) , .B1( u1_u10_u0_n146 ) , .A1( u1_u10_u0_n147 ) , .B2( u1_u10_u0_n161 ) );
  NAND3_X1 u1_u10_u0_U88 (.ZN( u1_out10_23 ) , .A3( u1_u10_u0_n137 ) , .A1( u1_u10_u0_n168 ) , .A2( u1_u10_u0_n171 ) );
  NAND3_X1 u1_u10_u0_U89 (.A3( u1_u10_u0_n127 ) , .A2( u1_u10_u0_n128 ) , .ZN( u1_u10_u0_n135 ) , .A1( u1_u10_u0_n150 ) );
  AND2_X1 u1_u10_u0_U9 (.A1( u1_u10_u0_n131 ) , .ZN( u1_u10_u0_n141 ) , .A2( u1_u10_u0_n150 ) );
  NAND3_X1 u1_u10_u0_U90 (.ZN( u1_u10_u0_n117 ) , .A3( u1_u10_u0_n132 ) , .A2( u1_u10_u0_n139 ) , .A1( u1_u10_u0_n148 ) );
  NAND3_X1 u1_u10_u0_U91 (.ZN( u1_u10_u0_n109 ) , .A2( u1_u10_u0_n114 ) , .A3( u1_u10_u0_n140 ) , .A1( u1_u10_u0_n149 ) );
  NAND3_X1 u1_u10_u0_U92 (.ZN( u1_out10_9 ) , .A3( u1_u10_u0_n106 ) , .A2( u1_u10_u0_n171 ) , .A1( u1_u10_u0_n174 ) );
  NAND3_X1 u1_u10_u0_U93 (.A2( u1_u10_u0_n128 ) , .A1( u1_u10_u0_n132 ) , .A3( u1_u10_u0_n146 ) , .ZN( u1_u10_u0_n97 ) );
  AOI21_X1 u1_u10_u1_U10 (.B2( u1_u10_u1_n155 ) , .B1( u1_u10_u1_n156 ) , .ZN( u1_u10_u1_n157 ) , .A( u1_u10_u1_n174 ) );
  NAND3_X1 u1_u10_u1_U100 (.ZN( u1_u10_u1_n113 ) , .A1( u1_u10_u1_n120 ) , .A3( u1_u10_u1_n133 ) , .A2( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U11 (.ZN( u1_u10_u1_n140 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n155 ) );
  NAND2_X1 u1_u10_u1_U12 (.A1( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n153 ) );
  AOI22_X1 u1_u10_u1_U13 (.B2( u1_u10_u1_n136 ) , .A2( u1_u10_u1_n137 ) , .ZN( u1_u10_u1_n143 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U14 (.A( u1_u10_u1_n147 ) , .ZN( u1_u10_u1_n181 ) );
  INV_X1 u1_u10_u1_U15 (.A( u1_u10_u1_n139 ) , .ZN( u1_u10_u1_n174 ) );
  OR4_X1 u1_u10_u1_U16 (.A4( u1_u10_u1_n106 ) , .A3( u1_u10_u1_n107 ) , .ZN( u1_u10_u1_n108 ) , .A1( u1_u10_u1_n117 ) , .A2( u1_u10_u1_n184 ) );
  AOI21_X1 u1_u10_u1_U17 (.ZN( u1_u10_u1_n106 ) , .A( u1_u10_u1_n112 ) , .B1( u1_u10_u1_n154 ) , .B2( u1_u10_u1_n156 ) );
  AOI21_X1 u1_u10_u1_U18 (.ZN( u1_u10_u1_n107 ) , .B1( u1_u10_u1_n134 ) , .B2( u1_u10_u1_n149 ) , .A( u1_u10_u1_n174 ) );
  INV_X1 u1_u10_u1_U19 (.A( u1_u10_u1_n101 ) , .ZN( u1_u10_u1_n184 ) );
  INV_X1 u1_u10_u1_U20 (.A( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n171 ) );
  NAND2_X1 u1_u10_u1_U21 (.ZN( u1_u10_u1_n141 ) , .A1( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n156 ) );
  AND2_X1 u1_u10_u1_U22 (.A1( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n161 ) );
  NAND2_X1 u1_u10_u1_U23 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n148 ) );
  NAND2_X1 u1_u10_u1_U24 (.A2( u1_u10_u1_n133 ) , .A1( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n159 ) );
  NAND2_X1 u1_u10_u1_U25 (.A2( u1_u10_u1_n115 ) , .A1( u1_u10_u1_n120 ) , .ZN( u1_u10_u1_n132 ) );
  INV_X1 u1_u10_u1_U26 (.A( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n178 ) );
  INV_X1 u1_u10_u1_U27 (.A( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n183 ) );
  AND2_X1 u1_u10_u1_U28 (.A1( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n149 ) );
  INV_X1 u1_u10_u1_U29 (.A( u1_u10_u1_n131 ) , .ZN( u1_u10_u1_n180 ) );
  INV_X1 u1_u10_u1_U3 (.A( u1_u10_u1_n159 ) , .ZN( u1_u10_u1_n182 ) );
  OAI221_X1 u1_u10_u1_U30 (.A( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n138 ) , .B2( u1_u10_u1_n152 ) , .C1( u1_u10_u1_n174 ) , .B1( u1_u10_u1_n187 ) );
  INV_X1 u1_u10_u1_U31 (.A( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n187 ) );
  AOI211_X1 u1_u10_u1_U32 (.B( u1_u10_u1_n117 ) , .A( u1_u10_u1_n118 ) , .ZN( u1_u10_u1_n119 ) , .C2( u1_u10_u1_n146 ) , .C1( u1_u10_u1_n159 ) );
  NOR2_X1 u1_u10_u1_U33 (.A1( u1_u10_u1_n168 ) , .A2( u1_u10_u1_n176 ) , .ZN( u1_u10_u1_n98 ) );
  AOI211_X1 u1_u10_u1_U34 (.B( u1_u10_u1_n162 ) , .A( u1_u10_u1_n163 ) , .C2( u1_u10_u1_n164 ) , .ZN( u1_u10_u1_n165 ) , .C1( u1_u10_u1_n171 ) );
  AOI21_X1 u1_u10_u1_U35 (.A( u1_u10_u1_n160 ) , .B2( u1_u10_u1_n161 ) , .ZN( u1_u10_u1_n162 ) , .B1( u1_u10_u1_n182 ) );
  OR2_X1 u1_u10_u1_U36 (.A2( u1_u10_u1_n157 ) , .A1( u1_u10_u1_n158 ) , .ZN( u1_u10_u1_n163 ) );
  OAI21_X1 u1_u10_u1_U37 (.B2( u1_u10_u1_n123 ) , .ZN( u1_u10_u1_n145 ) , .B1( u1_u10_u1_n160 ) , .A( u1_u10_u1_n185 ) );
  INV_X1 u1_u10_u1_U38 (.A( u1_u10_u1_n122 ) , .ZN( u1_u10_u1_n185 ) );
  AOI21_X1 u1_u10_u1_U39 (.B2( u1_u10_u1_n120 ) , .B1( u1_u10_u1_n121 ) , .ZN( u1_u10_u1_n122 ) , .A( u1_u10_u1_n128 ) );
  AOI221_X1 u1_u10_u1_U4 (.A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .C1( u1_u10_u1_n140 ) , .B2( u1_u10_u1_n141 ) , .ZN( u1_u10_u1_n142 ) , .B1( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U40 (.A1( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n146 ) , .A2( u1_u10_u1_n160 ) );
  NAND2_X1 u1_u10_u1_U41 (.A2( u1_u10_u1_n112 ) , .ZN( u1_u10_u1_n139 ) , .A1( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U42 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n156 ) , .A2( u1_u10_u1_n99 ) );
  AOI221_X1 u1_u10_u1_U43 (.B1( u1_u10_u1_n140 ) , .ZN( u1_u10_u1_n167 ) , .B2( u1_u10_u1_n172 ) , .C2( u1_u10_u1_n175 ) , .C1( u1_u10_u1_n178 ) , .A( u1_u10_u1_n188 ) );
  INV_X1 u1_u10_u1_U44 (.ZN( u1_u10_u1_n188 ) , .A( u1_u10_u1_n97 ) );
  AOI211_X1 u1_u10_u1_U45 (.A( u1_u10_u1_n118 ) , .C1( u1_u10_u1_n132 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n96 ) , .ZN( u1_u10_u1_n97 ) );
  AOI21_X1 u1_u10_u1_U46 (.B2( u1_u10_u1_n121 ) , .B1( u1_u10_u1_n135 ) , .A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n96 ) );
  NOR2_X1 u1_u10_u1_U47 (.ZN( u1_u10_u1_n117 ) , .A1( u1_u10_u1_n121 ) , .A2( u1_u10_u1_n160 ) );
  AOI21_X1 u1_u10_u1_U48 (.A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n129 ) , .ZN( u1_u10_u1_n130 ) , .B1( u1_u10_u1_n150 ) );
  NAND2_X1 u1_u10_u1_U49 (.ZN( u1_u10_u1_n112 ) , .A1( u1_u10_u1_n169 ) , .A2( u1_u10_u1_n170 ) );
  AOI211_X1 u1_u10_u1_U5 (.ZN( u1_u10_u1_n124 ) , .A( u1_u10_u1_n138 ) , .C2( u1_u10_u1_n139 ) , .B( u1_u10_u1_n145 ) , .C1( u1_u10_u1_n147 ) );
  NAND2_X1 u1_u10_u1_U50 (.ZN( u1_u10_u1_n129 ) , .A2( u1_u10_u1_n95 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U51 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n154 ) , .A2( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U52 (.A2( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n135 ) , .A1( u1_u10_u1_n99 ) );
  AOI21_X1 u1_u10_u1_U53 (.A( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n153 ) , .B1( u1_u10_u1_n154 ) , .ZN( u1_u10_u1_n158 ) );
  INV_X1 u1_u10_u1_U54 (.A( u1_u10_u1_n160 ) , .ZN( u1_u10_u1_n175 ) );
  NAND2_X1 u1_u10_u1_U55 (.A1( u1_u10_u1_n100 ) , .ZN( u1_u10_u1_n116 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U56 (.A1( u1_u10_u1_n102 ) , .ZN( u1_u10_u1_n131 ) , .A2( u1_u10_u1_n95 ) );
  NAND2_X1 u1_u10_u1_U57 (.A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n121 ) , .A1( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U58 (.A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n153 ) , .A2( u1_u10_u1_n98 ) );
  NAND2_X1 u1_u10_u1_U59 (.A2( u1_u10_u1_n104 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n133 ) );
  AOI22_X1 u1_u10_u1_U6 (.B2( u1_u10_u1_n113 ) , .A2( u1_u10_u1_n114 ) , .ZN( u1_u10_u1_n125 ) , .A1( u1_u10_u1_n171 ) , .B1( u1_u10_u1_n173 ) );
  NAND2_X1 u1_u10_u1_U60 (.ZN( u1_u10_u1_n150 ) , .A2( u1_u10_u1_n98 ) , .A1( u1_u10_u1_n99 ) );
  NAND2_X1 u1_u10_u1_U61 (.A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n155 ) , .A2( u1_u10_u1_n95 ) );
  OAI21_X1 u1_u10_u1_U62 (.ZN( u1_u10_u1_n109 ) , .B1( u1_u10_u1_n129 ) , .B2( u1_u10_u1_n160 ) , .A( u1_u10_u1_n167 ) );
  NAND2_X1 u1_u10_u1_U63 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n120 ) );
  NAND2_X1 u1_u10_u1_U64 (.A1( u1_u10_u1_n102 ) , .A2( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n115 ) );
  NAND2_X1 u1_u10_u1_U65 (.A2( u1_u10_u1_n100 ) , .A1( u1_u10_u1_n104 ) , .ZN( u1_u10_u1_n151 ) );
  NAND2_X1 u1_u10_u1_U66 (.A2( u1_u10_u1_n103 ) , .A1( u1_u10_u1_n105 ) , .ZN( u1_u10_u1_n161 ) );
  INV_X1 u1_u10_u1_U67 (.A( u1_u10_u1_n152 ) , .ZN( u1_u10_u1_n173 ) );
  INV_X1 u1_u10_u1_U68 (.A( u1_u10_u1_n128 ) , .ZN( u1_u10_u1_n172 ) );
  NAND2_X1 u1_u10_u1_U69 (.A2( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n103 ) , .ZN( u1_u10_u1_n123 ) );
  NAND2_X1 u1_u10_u1_U7 (.ZN( u1_u10_u1_n114 ) , .A1( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n156 ) );
  NOR2_X1 u1_u10_u1_U70 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n95 ) );
  NOR2_X1 u1_u10_u1_U71 (.A1( u1_u10_X_12 ) , .A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n100 ) );
  NOR2_X1 u1_u10_u1_U72 (.A2( u1_u10_X_8 ) , .A1( u1_u10_u1_n177 ) , .ZN( u1_u10_u1_n99 ) );
  NOR2_X1 u1_u10_u1_U73 (.A2( u1_u10_X_12 ) , .ZN( u1_u10_u1_n102 ) , .A1( u1_u10_u1_n176 ) );
  NOR2_X1 u1_u10_u1_U74 (.A2( u1_u10_X_9 ) , .ZN( u1_u10_u1_n105 ) , .A1( u1_u10_u1_n168 ) );
  NAND2_X1 u1_u10_u1_U75 (.A1( u1_u10_X_10 ) , .ZN( u1_u10_u1_n160 ) , .A2( u1_u10_u1_n169 ) );
  NAND2_X1 u1_u10_u1_U76 (.A2( u1_u10_X_10 ) , .A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n152 ) );
  NAND2_X1 u1_u10_u1_U77 (.A1( u1_u10_X_11 ) , .ZN( u1_u10_u1_n128 ) , .A2( u1_u10_u1_n170 ) );
  AND2_X1 u1_u10_u1_U78 (.A2( u1_u10_X_7 ) , .A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n104 ) );
  AND2_X1 u1_u10_u1_U79 (.A1( u1_u10_X_8 ) , .ZN( u1_u10_u1_n103 ) , .A2( u1_u10_u1_n177 ) );
  NOR2_X1 u1_u10_u1_U8 (.A1( u1_u10_u1_n112 ) , .A2( u1_u10_u1_n116 ) , .ZN( u1_u10_u1_n118 ) );
  INV_X1 u1_u10_u1_U80 (.A( u1_u10_X_10 ) , .ZN( u1_u10_u1_n170 ) );
  INV_X1 u1_u10_u1_U81 (.A( u1_u10_X_9 ) , .ZN( u1_u10_u1_n176 ) );
  INV_X1 u1_u10_u1_U82 (.A( u1_u10_X_11 ) , .ZN( u1_u10_u1_n169 ) );
  INV_X1 u1_u10_u1_U83 (.A( u1_u10_X_12 ) , .ZN( u1_u10_u1_n168 ) );
  INV_X1 u1_u10_u1_U84 (.A( u1_u10_X_7 ) , .ZN( u1_u10_u1_n177 ) );
  NAND4_X1 u1_u10_u1_U85 (.ZN( u1_out10_18 ) , .A4( u1_u10_u1_n165 ) , .A3( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n167 ) , .A2( u1_u10_u1_n186 ) );
  AOI22_X1 u1_u10_u1_U86 (.B2( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n147 ) , .A2( u1_u10_u1_n148 ) , .ZN( u1_u10_u1_n166 ) , .A1( u1_u10_u1_n172 ) );
  INV_X1 u1_u10_u1_U87 (.A( u1_u10_u1_n145 ) , .ZN( u1_u10_u1_n186 ) );
  NAND4_X1 u1_u10_u1_U88 (.ZN( u1_out10_2 ) , .A4( u1_u10_u1_n142 ) , .A3( u1_u10_u1_n143 ) , .A2( u1_u10_u1_n144 ) , .A1( u1_u10_u1_n179 ) );
  OAI21_X1 u1_u10_u1_U89 (.B2( u1_u10_u1_n132 ) , .ZN( u1_u10_u1_n144 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n180 ) );
  OAI21_X1 u1_u10_u1_U9 (.ZN( u1_u10_u1_n101 ) , .B1( u1_u10_u1_n141 ) , .A( u1_u10_u1_n146 ) , .B2( u1_u10_u1_n183 ) );
  INV_X1 u1_u10_u1_U90 (.A( u1_u10_u1_n130 ) , .ZN( u1_u10_u1_n179 ) );
  OR4_X1 u1_u10_u1_U91 (.ZN( u1_out10_13 ) , .A4( u1_u10_u1_n108 ) , .A3( u1_u10_u1_n109 ) , .A2( u1_u10_u1_n110 ) , .A1( u1_u10_u1_n111 ) );
  AOI21_X1 u1_u10_u1_U92 (.ZN( u1_u10_u1_n111 ) , .A( u1_u10_u1_n128 ) , .B2( u1_u10_u1_n131 ) , .B1( u1_u10_u1_n135 ) );
  AOI21_X1 u1_u10_u1_U93 (.ZN( u1_u10_u1_n110 ) , .A( u1_u10_u1_n116 ) , .B1( u1_u10_u1_n152 ) , .B2( u1_u10_u1_n160 ) );
  NAND4_X1 u1_u10_u1_U94 (.ZN( u1_out10_28 ) , .A4( u1_u10_u1_n124 ) , .A3( u1_u10_u1_n125 ) , .A2( u1_u10_u1_n126 ) , .A1( u1_u10_u1_n127 ) );
  OAI21_X1 u1_u10_u1_U95 (.ZN( u1_u10_u1_n127 ) , .B2( u1_u10_u1_n139 ) , .B1( u1_u10_u1_n175 ) , .A( u1_u10_u1_n183 ) );
  OAI21_X1 u1_u10_u1_U96 (.ZN( u1_u10_u1_n126 ) , .B2( u1_u10_u1_n140 ) , .A( u1_u10_u1_n146 ) , .B1( u1_u10_u1_n178 ) );
  NAND3_X1 u1_u10_u1_U97 (.A3( u1_u10_u1_n149 ) , .A2( u1_u10_u1_n150 ) , .A1( u1_u10_u1_n151 ) , .ZN( u1_u10_u1_n164 ) );
  NAND3_X1 u1_u10_u1_U98 (.A3( u1_u10_u1_n134 ) , .A2( u1_u10_u1_n135 ) , .ZN( u1_u10_u1_n136 ) , .A1( u1_u10_u1_n151 ) );
  NAND3_X1 u1_u10_u1_U99 (.A1( u1_u10_u1_n133 ) , .ZN( u1_u10_u1_n137 ) , .A2( u1_u10_u1_n154 ) , .A3( u1_u10_u1_n181 ) );
  OAI22_X1 u1_u10_u4_U10 (.B2( u1_u10_u4_n135 ) , .ZN( u1_u10_u4_n137 ) , .B1( u1_u10_u4_n153 ) , .A1( u1_u10_u4_n155 ) , .A2( u1_u10_u4_n171 ) );
  AND3_X1 u1_u10_u4_U11 (.A2( u1_u10_u4_n134 ) , .ZN( u1_u10_u4_n135 ) , .A3( u1_u10_u4_n145 ) , .A1( u1_u10_u4_n157 ) );
  NAND2_X1 u1_u10_u4_U12 (.ZN( u1_u10_u4_n132 ) , .A2( u1_u10_u4_n170 ) , .A1( u1_u10_u4_n173 ) );
  AOI21_X1 u1_u10_u4_U13 (.B2( u1_u10_u4_n160 ) , .B1( u1_u10_u4_n161 ) , .ZN( u1_u10_u4_n162 ) , .A( u1_u10_u4_n170 ) );
  AOI21_X1 u1_u10_u4_U14 (.ZN( u1_u10_u4_n107 ) , .B2( u1_u10_u4_n143 ) , .A( u1_u10_u4_n174 ) , .B1( u1_u10_u4_n184 ) );
  AOI21_X1 u1_u10_u4_U15 (.B2( u1_u10_u4_n158 ) , .B1( u1_u10_u4_n159 ) , .ZN( u1_u10_u4_n163 ) , .A( u1_u10_u4_n174 ) );
  AOI21_X1 u1_u10_u4_U16 (.A( u1_u10_u4_n153 ) , .B2( u1_u10_u4_n154 ) , .B1( u1_u10_u4_n155 ) , .ZN( u1_u10_u4_n165 ) );
  AOI21_X1 u1_u10_u4_U17 (.A( u1_u10_u4_n156 ) , .B2( u1_u10_u4_n157 ) , .ZN( u1_u10_u4_n164 ) , .B1( u1_u10_u4_n184 ) );
  INV_X1 u1_u10_u4_U18 (.A( u1_u10_u4_n138 ) , .ZN( u1_u10_u4_n170 ) );
  AND2_X1 u1_u10_u4_U19 (.A2( u1_u10_u4_n120 ) , .ZN( u1_u10_u4_n155 ) , .A1( u1_u10_u4_n160 ) );
  INV_X1 u1_u10_u4_U20 (.A( u1_u10_u4_n156 ) , .ZN( u1_u10_u4_n175 ) );
  NAND2_X1 u1_u10_u4_U21 (.A2( u1_u10_u4_n118 ) , .ZN( u1_u10_u4_n131 ) , .A1( u1_u10_u4_n147 ) );
  NAND2_X1 u1_u10_u4_U22 (.A1( u1_u10_u4_n119 ) , .A2( u1_u10_u4_n120 ) , .ZN( u1_u10_u4_n130 ) );
  NAND2_X1 u1_u10_u4_U23 (.ZN( u1_u10_u4_n117 ) , .A2( u1_u10_u4_n118 ) , .A1( u1_u10_u4_n148 ) );
  NAND2_X1 u1_u10_u4_U24 (.ZN( u1_u10_u4_n129 ) , .A1( u1_u10_u4_n134 ) , .A2( u1_u10_u4_n148 ) );
  AND3_X1 u1_u10_u4_U25 (.A1( u1_u10_u4_n119 ) , .A2( u1_u10_u4_n143 ) , .A3( u1_u10_u4_n154 ) , .ZN( u1_u10_u4_n161 ) );
  AND2_X1 u1_u10_u4_U26 (.A1( u1_u10_u4_n145 ) , .A2( u1_u10_u4_n147 ) , .ZN( u1_u10_u4_n159 ) );
  OR3_X1 u1_u10_u4_U27 (.A3( u1_u10_u4_n114 ) , .A2( u1_u10_u4_n115 ) , .A1( u1_u10_u4_n116 ) , .ZN( u1_u10_u4_n136 ) );
  AOI21_X1 u1_u10_u4_U28 (.A( u1_u10_u4_n113 ) , .ZN( u1_u10_u4_n116 ) , .B2( u1_u10_u4_n173 ) , .B1( u1_u10_u4_n174 ) );
  AOI21_X1 u1_u10_u4_U29 (.ZN( u1_u10_u4_n115 ) , .B2( u1_u10_u4_n145 ) , .B1( u1_u10_u4_n146 ) , .A( u1_u10_u4_n156 ) );
  NOR2_X1 u1_u10_u4_U3 (.ZN( u1_u10_u4_n121 ) , .A1( u1_u10_u4_n181 ) , .A2( u1_u10_u4_n182 ) );
  OAI22_X1 u1_u10_u4_U30 (.ZN( u1_u10_u4_n114 ) , .A2( u1_u10_u4_n121 ) , .B1( u1_u10_u4_n160 ) , .B2( u1_u10_u4_n170 ) , .A1( u1_u10_u4_n171 ) );
  INV_X1 u1_u10_u4_U31 (.A( u1_u10_u4_n158 ) , .ZN( u1_u10_u4_n182 ) );
  INV_X1 u1_u10_u4_U32 (.ZN( u1_u10_u4_n181 ) , .A( u1_u10_u4_n96 ) );
  INV_X1 u1_u10_u4_U33 (.A( u1_u10_u4_n144 ) , .ZN( u1_u10_u4_n179 ) );
  INV_X1 u1_u10_u4_U34 (.A( u1_u10_u4_n157 ) , .ZN( u1_u10_u4_n178 ) );
  NAND2_X1 u1_u10_u4_U35 (.A2( u1_u10_u4_n154 ) , .A1( u1_u10_u4_n96 ) , .ZN( u1_u10_u4_n97 ) );
  INV_X1 u1_u10_u4_U36 (.ZN( u1_u10_u4_n186 ) , .A( u1_u10_u4_n95 ) );
  OAI221_X1 u1_u10_u4_U37 (.C1( u1_u10_u4_n134 ) , .B1( u1_u10_u4_n158 ) , .B2( u1_u10_u4_n171 ) , .C2( u1_u10_u4_n173 ) , .A( u1_u10_u4_n94 ) , .ZN( u1_u10_u4_n95 ) );
  AOI222_X1 u1_u10_u4_U38 (.B2( u1_u10_u4_n132 ) , .A1( u1_u10_u4_n138 ) , .C2( u1_u10_u4_n175 ) , .A2( u1_u10_u4_n179 ) , .C1( u1_u10_u4_n181 ) , .B1( u1_u10_u4_n185 ) , .ZN( u1_u10_u4_n94 ) );
  INV_X1 u1_u10_u4_U39 (.A( u1_u10_u4_n113 ) , .ZN( u1_u10_u4_n185 ) );
  INV_X1 u1_u10_u4_U4 (.A( u1_u10_u4_n117 ) , .ZN( u1_u10_u4_n184 ) );
  INV_X1 u1_u10_u4_U40 (.A( u1_u10_u4_n143 ) , .ZN( u1_u10_u4_n183 ) );
  NOR2_X1 u1_u10_u4_U41 (.ZN( u1_u10_u4_n138 ) , .A1( u1_u10_u4_n168 ) , .A2( u1_u10_u4_n169 ) );
  NOR2_X1 u1_u10_u4_U42 (.A1( u1_u10_u4_n150 ) , .A2( u1_u10_u4_n152 ) , .ZN( u1_u10_u4_n153 ) );
  NOR2_X1 u1_u10_u4_U43 (.A2( u1_u10_u4_n128 ) , .A1( u1_u10_u4_n138 ) , .ZN( u1_u10_u4_n156 ) );
  AOI22_X1 u1_u10_u4_U44 (.B2( u1_u10_u4_n122 ) , .A1( u1_u10_u4_n123 ) , .ZN( u1_u10_u4_n124 ) , .B1( u1_u10_u4_n128 ) , .A2( u1_u10_u4_n172 ) );
  INV_X1 u1_u10_u4_U45 (.A( u1_u10_u4_n153 ) , .ZN( u1_u10_u4_n172 ) );
  NAND2_X1 u1_u10_u4_U46 (.A2( u1_u10_u4_n120 ) , .ZN( u1_u10_u4_n123 ) , .A1( u1_u10_u4_n161 ) );
  AOI22_X1 u1_u10_u4_U47 (.B2( u1_u10_u4_n132 ) , .A2( u1_u10_u4_n133 ) , .ZN( u1_u10_u4_n140 ) , .A1( u1_u10_u4_n150 ) , .B1( u1_u10_u4_n179 ) );
  NAND2_X1 u1_u10_u4_U48 (.ZN( u1_u10_u4_n133 ) , .A2( u1_u10_u4_n146 ) , .A1( u1_u10_u4_n154 ) );
  NAND2_X1 u1_u10_u4_U49 (.A1( u1_u10_u4_n103 ) , .ZN( u1_u10_u4_n154 ) , .A2( u1_u10_u4_n98 ) );
  NOR4_X1 u1_u10_u4_U5 (.A4( u1_u10_u4_n106 ) , .A3( u1_u10_u4_n107 ) , .A2( u1_u10_u4_n108 ) , .A1( u1_u10_u4_n109 ) , .ZN( u1_u10_u4_n110 ) );
  NAND2_X1 u1_u10_u4_U50 (.A1( u1_u10_u4_n101 ) , .ZN( u1_u10_u4_n158 ) , .A2( u1_u10_u4_n99 ) );
  AOI21_X1 u1_u10_u4_U51 (.ZN( u1_u10_u4_n127 ) , .A( u1_u10_u4_n136 ) , .B2( u1_u10_u4_n150 ) , .B1( u1_u10_u4_n180 ) );
  INV_X1 u1_u10_u4_U52 (.A( u1_u10_u4_n160 ) , .ZN( u1_u10_u4_n180 ) );
  NAND2_X1 u1_u10_u4_U53 (.A2( u1_u10_u4_n104 ) , .A1( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n146 ) );
  NAND2_X1 u1_u10_u4_U54 (.A2( u1_u10_u4_n101 ) , .A1( u1_u10_u4_n102 ) , .ZN( u1_u10_u4_n160 ) );
  NAND2_X1 u1_u10_u4_U55 (.ZN( u1_u10_u4_n134 ) , .A1( u1_u10_u4_n98 ) , .A2( u1_u10_u4_n99 ) );
  NAND2_X1 u1_u10_u4_U56 (.A1( u1_u10_u4_n103 ) , .A2( u1_u10_u4_n104 ) , .ZN( u1_u10_u4_n143 ) );
  NAND2_X1 u1_u10_u4_U57 (.A2( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n145 ) , .A1( u1_u10_u4_n98 ) );
  NAND2_X1 u1_u10_u4_U58 (.A1( u1_u10_u4_n100 ) , .A2( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n120 ) );
  NAND2_X1 u1_u10_u4_U59 (.A1( u1_u10_u4_n102 ) , .A2( u1_u10_u4_n104 ) , .ZN( u1_u10_u4_n148 ) );
  AOI21_X1 u1_u10_u4_U6 (.ZN( u1_u10_u4_n106 ) , .B2( u1_u10_u4_n146 ) , .B1( u1_u10_u4_n158 ) , .A( u1_u10_u4_n170 ) );
  NAND2_X1 u1_u10_u4_U60 (.A2( u1_u10_u4_n100 ) , .A1( u1_u10_u4_n103 ) , .ZN( u1_u10_u4_n157 ) );
  INV_X1 u1_u10_u4_U61 (.A( u1_u10_u4_n150 ) , .ZN( u1_u10_u4_n173 ) );
  INV_X1 u1_u10_u4_U62 (.A( u1_u10_u4_n152 ) , .ZN( u1_u10_u4_n171 ) );
  NAND2_X1 u1_u10_u4_U63 (.A1( u1_u10_u4_n100 ) , .ZN( u1_u10_u4_n118 ) , .A2( u1_u10_u4_n99 ) );
  NAND2_X1 u1_u10_u4_U64 (.A2( u1_u10_u4_n100 ) , .A1( u1_u10_u4_n102 ) , .ZN( u1_u10_u4_n144 ) );
  NAND2_X1 u1_u10_u4_U65 (.A2( u1_u10_u4_n101 ) , .A1( u1_u10_u4_n105 ) , .ZN( u1_u10_u4_n96 ) );
  INV_X1 u1_u10_u4_U66 (.A( u1_u10_u4_n128 ) , .ZN( u1_u10_u4_n174 ) );
  NAND2_X1 u1_u10_u4_U67 (.A2( u1_u10_u4_n102 ) , .ZN( u1_u10_u4_n119 ) , .A1( u1_u10_u4_n98 ) );
  NAND2_X1 u1_u10_u4_U68 (.A2( u1_u10_u4_n101 ) , .A1( u1_u10_u4_n103 ) , .ZN( u1_u10_u4_n147 ) );
  NAND2_X1 u1_u10_u4_U69 (.A2( u1_u10_u4_n104 ) , .ZN( u1_u10_u4_n113 ) , .A1( u1_u10_u4_n99 ) );
  AOI21_X1 u1_u10_u4_U7 (.ZN( u1_u10_u4_n108 ) , .B2( u1_u10_u4_n134 ) , .B1( u1_u10_u4_n155 ) , .A( u1_u10_u4_n156 ) );
  NOR2_X1 u1_u10_u4_U70 (.A2( u1_u10_X_28 ) , .ZN( u1_u10_u4_n150 ) , .A1( u1_u10_u4_n168 ) );
  NOR2_X1 u1_u10_u4_U71 (.A2( u1_u10_X_29 ) , .ZN( u1_u10_u4_n152 ) , .A1( u1_u10_u4_n169 ) );
  NOR2_X1 u1_u10_u4_U72 (.A2( u1_u10_X_30 ) , .ZN( u1_u10_u4_n105 ) , .A1( u1_u10_u4_n176 ) );
  NOR2_X1 u1_u10_u4_U73 (.A2( u1_u10_X_26 ) , .ZN( u1_u10_u4_n100 ) , .A1( u1_u10_u4_n177 ) );
  NOR2_X1 u1_u10_u4_U74 (.A2( u1_u10_X_28 ) , .A1( u1_u10_X_29 ) , .ZN( u1_u10_u4_n128 ) );
  NOR2_X1 u1_u10_u4_U75 (.A2( u1_u10_X_27 ) , .A1( u1_u10_X_30 ) , .ZN( u1_u10_u4_n102 ) );
  NOR2_X1 u1_u10_u4_U76 (.A2( u1_u10_X_25 ) , .A1( u1_u10_X_26 ) , .ZN( u1_u10_u4_n98 ) );
  AND2_X1 u1_u10_u4_U77 (.A2( u1_u10_X_25 ) , .A1( u1_u10_X_26 ) , .ZN( u1_u10_u4_n104 ) );
  AND2_X1 u1_u10_u4_U78 (.A1( u1_u10_X_30 ) , .A2( u1_u10_u4_n176 ) , .ZN( u1_u10_u4_n99 ) );
  AND2_X1 u1_u10_u4_U79 (.A1( u1_u10_X_26 ) , .ZN( u1_u10_u4_n101 ) , .A2( u1_u10_u4_n177 ) );
  AOI21_X1 u1_u10_u4_U8 (.ZN( u1_u10_u4_n109 ) , .A( u1_u10_u4_n153 ) , .B1( u1_u10_u4_n159 ) , .B2( u1_u10_u4_n184 ) );
  AND2_X1 u1_u10_u4_U80 (.A1( u1_u10_X_27 ) , .A2( u1_u10_X_30 ) , .ZN( u1_u10_u4_n103 ) );
  INV_X1 u1_u10_u4_U81 (.A( u1_u10_X_28 ) , .ZN( u1_u10_u4_n169 ) );
  INV_X1 u1_u10_u4_U82 (.A( u1_u10_X_29 ) , .ZN( u1_u10_u4_n168 ) );
  INV_X1 u1_u10_u4_U83 (.A( u1_u10_X_25 ) , .ZN( u1_u10_u4_n177 ) );
  INV_X1 u1_u10_u4_U84 (.A( u1_u10_X_27 ) , .ZN( u1_u10_u4_n176 ) );
  NAND4_X1 u1_u10_u4_U85 (.ZN( u1_out10_25 ) , .A4( u1_u10_u4_n139 ) , .A3( u1_u10_u4_n140 ) , .A2( u1_u10_u4_n141 ) , .A1( u1_u10_u4_n142 ) );
  OAI21_X1 u1_u10_u4_U86 (.A( u1_u10_u4_n128 ) , .B2( u1_u10_u4_n129 ) , .B1( u1_u10_u4_n130 ) , .ZN( u1_u10_u4_n142 ) );
  OAI21_X1 u1_u10_u4_U87 (.B2( u1_u10_u4_n131 ) , .ZN( u1_u10_u4_n141 ) , .A( u1_u10_u4_n175 ) , .B1( u1_u10_u4_n183 ) );
  NAND4_X1 u1_u10_u4_U88 (.ZN( u1_out10_14 ) , .A4( u1_u10_u4_n124 ) , .A3( u1_u10_u4_n125 ) , .A2( u1_u10_u4_n126 ) , .A1( u1_u10_u4_n127 ) );
  AOI22_X1 u1_u10_u4_U89 (.B2( u1_u10_u4_n117 ) , .ZN( u1_u10_u4_n126 ) , .A1( u1_u10_u4_n129 ) , .B1( u1_u10_u4_n152 ) , .A2( u1_u10_u4_n175 ) );
  AOI211_X1 u1_u10_u4_U9 (.B( u1_u10_u4_n136 ) , .A( u1_u10_u4_n137 ) , .C2( u1_u10_u4_n138 ) , .ZN( u1_u10_u4_n139 ) , .C1( u1_u10_u4_n182 ) );
  AOI22_X1 u1_u10_u4_U90 (.ZN( u1_u10_u4_n125 ) , .B2( u1_u10_u4_n131 ) , .A2( u1_u10_u4_n132 ) , .B1( u1_u10_u4_n138 ) , .A1( u1_u10_u4_n178 ) );
  NAND4_X1 u1_u10_u4_U91 (.ZN( u1_out10_8 ) , .A4( u1_u10_u4_n110 ) , .A3( u1_u10_u4_n111 ) , .A2( u1_u10_u4_n112 ) , .A1( u1_u10_u4_n186 ) );
  NAND2_X1 u1_u10_u4_U92 (.ZN( u1_u10_u4_n112 ) , .A2( u1_u10_u4_n130 ) , .A1( u1_u10_u4_n150 ) );
  AOI22_X1 u1_u10_u4_U93 (.ZN( u1_u10_u4_n111 ) , .B2( u1_u10_u4_n132 ) , .A1( u1_u10_u4_n152 ) , .B1( u1_u10_u4_n178 ) , .A2( u1_u10_u4_n97 ) );
  AOI22_X1 u1_u10_u4_U94 (.B2( u1_u10_u4_n149 ) , .B1( u1_u10_u4_n150 ) , .A2( u1_u10_u4_n151 ) , .A1( u1_u10_u4_n152 ) , .ZN( u1_u10_u4_n167 ) );
  NOR4_X1 u1_u10_u4_U95 (.A4( u1_u10_u4_n162 ) , .A3( u1_u10_u4_n163 ) , .A2( u1_u10_u4_n164 ) , .A1( u1_u10_u4_n165 ) , .ZN( u1_u10_u4_n166 ) );
  NAND3_X1 u1_u10_u4_U96 (.ZN( u1_out10_3 ) , .A3( u1_u10_u4_n166 ) , .A1( u1_u10_u4_n167 ) , .A2( u1_u10_u4_n186 ) );
  NAND3_X1 u1_u10_u4_U97 (.A3( u1_u10_u4_n146 ) , .A2( u1_u10_u4_n147 ) , .A1( u1_u10_u4_n148 ) , .ZN( u1_u10_u4_n149 ) );
  NAND3_X1 u1_u10_u4_U98 (.A3( u1_u10_u4_n143 ) , .A2( u1_u10_u4_n144 ) , .A1( u1_u10_u4_n145 ) , .ZN( u1_u10_u4_n151 ) );
  NAND3_X1 u1_u10_u4_U99 (.A3( u1_u10_u4_n121 ) , .ZN( u1_u10_u4_n122 ) , .A2( u1_u10_u4_n144 ) , .A1( u1_u10_u4_n154 ) );
  INV_X1 u1_u10_u5_U10 (.A( u1_u10_u5_n121 ) , .ZN( u1_u10_u5_n177 ) );
  NOR3_X1 u1_u10_u5_U100 (.A3( u1_u10_u5_n141 ) , .A1( u1_u10_u5_n142 ) , .ZN( u1_u10_u5_n143 ) , .A2( u1_u10_u5_n191 ) );
  NAND4_X1 u1_u10_u5_U101 (.ZN( u1_out10_4 ) , .A4( u1_u10_u5_n112 ) , .A2( u1_u10_u5_n113 ) , .A1( u1_u10_u5_n114 ) , .A3( u1_u10_u5_n195 ) );
  AOI211_X1 u1_u10_u5_U102 (.A( u1_u10_u5_n110 ) , .C1( u1_u10_u5_n111 ) , .ZN( u1_u10_u5_n112 ) , .B( u1_u10_u5_n118 ) , .C2( u1_u10_u5_n177 ) );
  AOI222_X1 u1_u10_u5_U103 (.ZN( u1_u10_u5_n113 ) , .A1( u1_u10_u5_n131 ) , .C1( u1_u10_u5_n148 ) , .B2( u1_u10_u5_n174 ) , .C2( u1_u10_u5_n178 ) , .A2( u1_u10_u5_n179 ) , .B1( u1_u10_u5_n99 ) );
  NAND3_X1 u1_u10_u5_U104 (.A2( u1_u10_u5_n154 ) , .A3( u1_u10_u5_n158 ) , .A1( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n99 ) );
  NOR2_X1 u1_u10_u5_U11 (.ZN( u1_u10_u5_n160 ) , .A2( u1_u10_u5_n173 ) , .A1( u1_u10_u5_n177 ) );
  INV_X1 u1_u10_u5_U12 (.A( u1_u10_u5_n150 ) , .ZN( u1_u10_u5_n174 ) );
  AOI21_X1 u1_u10_u5_U13 (.A( u1_u10_u5_n160 ) , .B2( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n162 ) , .B1( u1_u10_u5_n192 ) );
  INV_X1 u1_u10_u5_U14 (.A( u1_u10_u5_n159 ) , .ZN( u1_u10_u5_n192 ) );
  AOI21_X1 u1_u10_u5_U15 (.A( u1_u10_u5_n156 ) , .B2( u1_u10_u5_n157 ) , .B1( u1_u10_u5_n158 ) , .ZN( u1_u10_u5_n163 ) );
  AOI21_X1 u1_u10_u5_U16 (.B2( u1_u10_u5_n139 ) , .B1( u1_u10_u5_n140 ) , .ZN( u1_u10_u5_n141 ) , .A( u1_u10_u5_n150 ) );
  OAI21_X1 u1_u10_u5_U17 (.A( u1_u10_u5_n133 ) , .B2( u1_u10_u5_n134 ) , .B1( u1_u10_u5_n135 ) , .ZN( u1_u10_u5_n142 ) );
  OAI21_X1 u1_u10_u5_U18 (.ZN( u1_u10_u5_n133 ) , .B2( u1_u10_u5_n147 ) , .A( u1_u10_u5_n173 ) , .B1( u1_u10_u5_n188 ) );
  NAND2_X1 u1_u10_u5_U19 (.A2( u1_u10_u5_n119 ) , .A1( u1_u10_u5_n123 ) , .ZN( u1_u10_u5_n137 ) );
  INV_X1 u1_u10_u5_U20 (.A( u1_u10_u5_n155 ) , .ZN( u1_u10_u5_n194 ) );
  NAND2_X1 u1_u10_u5_U21 (.A1( u1_u10_u5_n121 ) , .ZN( u1_u10_u5_n132 ) , .A2( u1_u10_u5_n172 ) );
  NAND2_X1 u1_u10_u5_U22 (.A2( u1_u10_u5_n122 ) , .ZN( u1_u10_u5_n136 ) , .A1( u1_u10_u5_n154 ) );
  NAND2_X1 u1_u10_u5_U23 (.A2( u1_u10_u5_n119 ) , .A1( u1_u10_u5_n120 ) , .ZN( u1_u10_u5_n159 ) );
  INV_X1 u1_u10_u5_U24 (.A( u1_u10_u5_n156 ) , .ZN( u1_u10_u5_n175 ) );
  INV_X1 u1_u10_u5_U25 (.A( u1_u10_u5_n158 ) , .ZN( u1_u10_u5_n188 ) );
  INV_X1 u1_u10_u5_U26 (.A( u1_u10_u5_n152 ) , .ZN( u1_u10_u5_n179 ) );
  INV_X1 u1_u10_u5_U27 (.A( u1_u10_u5_n140 ) , .ZN( u1_u10_u5_n182 ) );
  INV_X1 u1_u10_u5_U28 (.A( u1_u10_u5_n151 ) , .ZN( u1_u10_u5_n183 ) );
  INV_X1 u1_u10_u5_U29 (.A( u1_u10_u5_n123 ) , .ZN( u1_u10_u5_n185 ) );
  NOR2_X1 u1_u10_u5_U3 (.ZN( u1_u10_u5_n134 ) , .A1( u1_u10_u5_n183 ) , .A2( u1_u10_u5_n190 ) );
  INV_X1 u1_u10_u5_U30 (.A( u1_u10_u5_n161 ) , .ZN( u1_u10_u5_n184 ) );
  INV_X1 u1_u10_u5_U31 (.A( u1_u10_u5_n139 ) , .ZN( u1_u10_u5_n189 ) );
  INV_X1 u1_u10_u5_U32 (.A( u1_u10_u5_n157 ) , .ZN( u1_u10_u5_n190 ) );
  INV_X1 u1_u10_u5_U33 (.A( u1_u10_u5_n120 ) , .ZN( u1_u10_u5_n193 ) );
  NAND2_X1 u1_u10_u5_U34 (.ZN( u1_u10_u5_n111 ) , .A1( u1_u10_u5_n140 ) , .A2( u1_u10_u5_n155 ) );
  INV_X1 u1_u10_u5_U35 (.A( u1_u10_u5_n117 ) , .ZN( u1_u10_u5_n196 ) );
  OAI221_X1 u1_u10_u5_U36 (.A( u1_u10_u5_n116 ) , .ZN( u1_u10_u5_n117 ) , .B2( u1_u10_u5_n119 ) , .C1( u1_u10_u5_n153 ) , .C2( u1_u10_u5_n158 ) , .B1( u1_u10_u5_n172 ) );
  AOI222_X1 u1_u10_u5_U37 (.ZN( u1_u10_u5_n116 ) , .B2( u1_u10_u5_n145 ) , .C1( u1_u10_u5_n148 ) , .A2( u1_u10_u5_n174 ) , .C2( u1_u10_u5_n177 ) , .B1( u1_u10_u5_n187 ) , .A1( u1_u10_u5_n193 ) );
  INV_X1 u1_u10_u5_U38 (.A( u1_u10_u5_n115 ) , .ZN( u1_u10_u5_n187 ) );
  NOR2_X1 u1_u10_u5_U39 (.ZN( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n170 ) , .A2( u1_u10_u5_n180 ) );
  INV_X1 u1_u10_u5_U4 (.A( u1_u10_u5_n138 ) , .ZN( u1_u10_u5_n191 ) );
  AOI22_X1 u1_u10_u5_U40 (.B2( u1_u10_u5_n131 ) , .A2( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n169 ) , .B1( u1_u10_u5_n174 ) , .A1( u1_u10_u5_n185 ) );
  NOR2_X1 u1_u10_u5_U41 (.A1( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n150 ) , .A2( u1_u10_u5_n173 ) );
  AOI21_X1 u1_u10_u5_U42 (.A( u1_u10_u5_n118 ) , .B2( u1_u10_u5_n145 ) , .ZN( u1_u10_u5_n168 ) , .B1( u1_u10_u5_n186 ) );
  INV_X1 u1_u10_u5_U43 (.A( u1_u10_u5_n122 ) , .ZN( u1_u10_u5_n186 ) );
  NOR2_X1 u1_u10_u5_U44 (.A1( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n152 ) , .A2( u1_u10_u5_n176 ) );
  NOR2_X1 u1_u10_u5_U45 (.A1( u1_u10_u5_n115 ) , .ZN( u1_u10_u5_n118 ) , .A2( u1_u10_u5_n153 ) );
  NOR2_X1 u1_u10_u5_U46 (.A2( u1_u10_u5_n145 ) , .ZN( u1_u10_u5_n156 ) , .A1( u1_u10_u5_n174 ) );
  NOR2_X1 u1_u10_u5_U47 (.ZN( u1_u10_u5_n121 ) , .A2( u1_u10_u5_n145 ) , .A1( u1_u10_u5_n176 ) );
  AOI22_X1 u1_u10_u5_U48 (.ZN( u1_u10_u5_n114 ) , .A2( u1_u10_u5_n137 ) , .A1( u1_u10_u5_n145 ) , .B2( u1_u10_u5_n175 ) , .B1( u1_u10_u5_n193 ) );
  OAI211_X1 u1_u10_u5_U49 (.B( u1_u10_u5_n124 ) , .A( u1_u10_u5_n125 ) , .C2( u1_u10_u5_n126 ) , .C1( u1_u10_u5_n127 ) , .ZN( u1_u10_u5_n128 ) );
  OAI21_X1 u1_u10_u5_U5 (.B2( u1_u10_u5_n136 ) , .B1( u1_u10_u5_n137 ) , .ZN( u1_u10_u5_n138 ) , .A( u1_u10_u5_n177 ) );
  NOR3_X1 u1_u10_u5_U50 (.ZN( u1_u10_u5_n127 ) , .A1( u1_u10_u5_n136 ) , .A3( u1_u10_u5_n148 ) , .A2( u1_u10_u5_n182 ) );
  OAI21_X1 u1_u10_u5_U51 (.ZN( u1_u10_u5_n124 ) , .A( u1_u10_u5_n177 ) , .B2( u1_u10_u5_n183 ) , .B1( u1_u10_u5_n189 ) );
  OAI21_X1 u1_u10_u5_U52 (.ZN( u1_u10_u5_n125 ) , .A( u1_u10_u5_n174 ) , .B2( u1_u10_u5_n185 ) , .B1( u1_u10_u5_n190 ) );
  AOI21_X1 u1_u10_u5_U53 (.A( u1_u10_u5_n153 ) , .B2( u1_u10_u5_n154 ) , .B1( u1_u10_u5_n155 ) , .ZN( u1_u10_u5_n164 ) );
  AOI21_X1 u1_u10_u5_U54 (.ZN( u1_u10_u5_n110 ) , .B1( u1_u10_u5_n122 ) , .B2( u1_u10_u5_n139 ) , .A( u1_u10_u5_n153 ) );
  INV_X1 u1_u10_u5_U55 (.A( u1_u10_u5_n153 ) , .ZN( u1_u10_u5_n176 ) );
  INV_X1 u1_u10_u5_U56 (.A( u1_u10_u5_n126 ) , .ZN( u1_u10_u5_n173 ) );
  AND2_X1 u1_u10_u5_U57 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n147 ) );
  AND2_X1 u1_u10_u5_U58 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n148 ) );
  NAND2_X1 u1_u10_u5_U59 (.A1( u1_u10_u5_n105 ) , .A2( u1_u10_u5_n106 ) , .ZN( u1_u10_u5_n158 ) );
  INV_X1 u1_u10_u5_U6 (.A( u1_u10_u5_n135 ) , .ZN( u1_u10_u5_n178 ) );
  NAND2_X1 u1_u10_u5_U60 (.A2( u1_u10_u5_n108 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n139 ) );
  NAND2_X1 u1_u10_u5_U61 (.A1( u1_u10_u5_n106 ) , .A2( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n119 ) );
  NAND2_X1 u1_u10_u5_U62 (.A2( u1_u10_u5_n103 ) , .A1( u1_u10_u5_n105 ) , .ZN( u1_u10_u5_n140 ) );
  NAND2_X1 u1_u10_u5_U63 (.A2( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n105 ) , .ZN( u1_u10_u5_n155 ) );
  NAND2_X1 u1_u10_u5_U64 (.A2( u1_u10_u5_n106 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n122 ) );
  NAND2_X1 u1_u10_u5_U65 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n106 ) , .ZN( u1_u10_u5_n115 ) );
  NAND2_X1 u1_u10_u5_U66 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n103 ) , .ZN( u1_u10_u5_n161 ) );
  NAND2_X1 u1_u10_u5_U67 (.A1( u1_u10_u5_n105 ) , .A2( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n154 ) );
  INV_X1 u1_u10_u5_U68 (.A( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n172 ) );
  NAND2_X1 u1_u10_u5_U69 (.A1( u1_u10_u5_n103 ) , .A2( u1_u10_u5_n108 ) , .ZN( u1_u10_u5_n123 ) );
  OAI22_X1 u1_u10_u5_U7 (.B2( u1_u10_u5_n149 ) , .B1( u1_u10_u5_n150 ) , .A2( u1_u10_u5_n151 ) , .A1( u1_u10_u5_n152 ) , .ZN( u1_u10_u5_n165 ) );
  NAND2_X1 u1_u10_u5_U70 (.A2( u1_u10_u5_n103 ) , .A1( u1_u10_u5_n107 ) , .ZN( u1_u10_u5_n151 ) );
  NAND2_X1 u1_u10_u5_U71 (.A2( u1_u10_u5_n107 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n120 ) );
  NAND2_X1 u1_u10_u5_U72 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n109 ) , .ZN( u1_u10_u5_n157 ) );
  AND2_X1 u1_u10_u5_U73 (.A2( u1_u10_u5_n100 ) , .A1( u1_u10_u5_n104 ) , .ZN( u1_u10_u5_n131 ) );
  INV_X1 u1_u10_u5_U74 (.A( u1_u10_u5_n102 ) , .ZN( u1_u10_u5_n195 ) );
  OAI221_X1 u1_u10_u5_U75 (.A( u1_u10_u5_n101 ) , .ZN( u1_u10_u5_n102 ) , .C2( u1_u10_u5_n115 ) , .C1( u1_u10_u5_n126 ) , .B1( u1_u10_u5_n134 ) , .B2( u1_u10_u5_n160 ) );
  OAI21_X1 u1_u10_u5_U76 (.ZN( u1_u10_u5_n101 ) , .B1( u1_u10_u5_n137 ) , .A( u1_u10_u5_n146 ) , .B2( u1_u10_u5_n147 ) );
  NOR2_X1 u1_u10_u5_U77 (.A2( u1_u10_X_34 ) , .A1( u1_u10_X_35 ) , .ZN( u1_u10_u5_n145 ) );
  NOR2_X1 u1_u10_u5_U78 (.A2( u1_u10_X_34 ) , .ZN( u1_u10_u5_n146 ) , .A1( u1_u10_u5_n171 ) );
  NOR2_X1 u1_u10_u5_U79 (.A2( u1_u10_X_31 ) , .A1( u1_u10_X_32 ) , .ZN( u1_u10_u5_n103 ) );
  NOR3_X1 u1_u10_u5_U8 (.A2( u1_u10_u5_n147 ) , .A1( u1_u10_u5_n148 ) , .ZN( u1_u10_u5_n149 ) , .A3( u1_u10_u5_n194 ) );
  NOR2_X1 u1_u10_u5_U80 (.A2( u1_u10_X_36 ) , .ZN( u1_u10_u5_n105 ) , .A1( u1_u10_u5_n180 ) );
  NOR2_X1 u1_u10_u5_U81 (.A2( u1_u10_X_33 ) , .ZN( u1_u10_u5_n108 ) , .A1( u1_u10_u5_n170 ) );
  NOR2_X1 u1_u10_u5_U82 (.A2( u1_u10_X_33 ) , .A1( u1_u10_X_36 ) , .ZN( u1_u10_u5_n107 ) );
  NOR2_X1 u1_u10_u5_U83 (.A2( u1_u10_X_31 ) , .ZN( u1_u10_u5_n104 ) , .A1( u1_u10_u5_n181 ) );
  NAND2_X1 u1_u10_u5_U84 (.A2( u1_u10_X_34 ) , .A1( u1_u10_X_35 ) , .ZN( u1_u10_u5_n153 ) );
  NAND2_X1 u1_u10_u5_U85 (.A1( u1_u10_X_34 ) , .ZN( u1_u10_u5_n126 ) , .A2( u1_u10_u5_n171 ) );
  AND2_X1 u1_u10_u5_U86 (.A1( u1_u10_X_31 ) , .A2( u1_u10_X_32 ) , .ZN( u1_u10_u5_n106 ) );
  AND2_X1 u1_u10_u5_U87 (.A1( u1_u10_X_31 ) , .ZN( u1_u10_u5_n109 ) , .A2( u1_u10_u5_n181 ) );
  INV_X1 u1_u10_u5_U88 (.A( u1_u10_X_33 ) , .ZN( u1_u10_u5_n180 ) );
  INV_X1 u1_u10_u5_U89 (.A( u1_u10_X_35 ) , .ZN( u1_u10_u5_n171 ) );
  NOR2_X1 u1_u10_u5_U9 (.ZN( u1_u10_u5_n135 ) , .A1( u1_u10_u5_n173 ) , .A2( u1_u10_u5_n176 ) );
  INV_X1 u1_u10_u5_U90 (.A( u1_u10_X_36 ) , .ZN( u1_u10_u5_n170 ) );
  INV_X1 u1_u10_u5_U91 (.A( u1_u10_X_32 ) , .ZN( u1_u10_u5_n181 ) );
  NAND4_X1 u1_u10_u5_U92 (.ZN( u1_out10_29 ) , .A4( u1_u10_u5_n129 ) , .A3( u1_u10_u5_n130 ) , .A2( u1_u10_u5_n168 ) , .A1( u1_u10_u5_n196 ) );
  AOI221_X1 u1_u10_u5_U93 (.A( u1_u10_u5_n128 ) , .ZN( u1_u10_u5_n129 ) , .C2( u1_u10_u5_n132 ) , .B2( u1_u10_u5_n159 ) , .B1( u1_u10_u5_n176 ) , .C1( u1_u10_u5_n184 ) );
  AOI222_X1 u1_u10_u5_U94 (.ZN( u1_u10_u5_n130 ) , .A2( u1_u10_u5_n146 ) , .B1( u1_u10_u5_n147 ) , .C2( u1_u10_u5_n175 ) , .B2( u1_u10_u5_n179 ) , .A1( u1_u10_u5_n188 ) , .C1( u1_u10_u5_n194 ) );
  NAND4_X1 u1_u10_u5_U95 (.ZN( u1_out10_19 ) , .A4( u1_u10_u5_n166 ) , .A3( u1_u10_u5_n167 ) , .A2( u1_u10_u5_n168 ) , .A1( u1_u10_u5_n169 ) );
  AOI22_X1 u1_u10_u5_U96 (.B2( u1_u10_u5_n145 ) , .A2( u1_u10_u5_n146 ) , .ZN( u1_u10_u5_n167 ) , .B1( u1_u10_u5_n182 ) , .A1( u1_u10_u5_n189 ) );
  NOR4_X1 u1_u10_u5_U97 (.A4( u1_u10_u5_n162 ) , .A3( u1_u10_u5_n163 ) , .A2( u1_u10_u5_n164 ) , .A1( u1_u10_u5_n165 ) , .ZN( u1_u10_u5_n166 ) );
  NAND4_X1 u1_u10_u5_U98 (.ZN( u1_out10_11 ) , .A4( u1_u10_u5_n143 ) , .A3( u1_u10_u5_n144 ) , .A2( u1_u10_u5_n169 ) , .A1( u1_u10_u5_n196 ) );
  AOI22_X1 u1_u10_u5_U99 (.A2( u1_u10_u5_n132 ) , .ZN( u1_u10_u5_n144 ) , .B2( u1_u10_u5_n145 ) , .B1( u1_u10_u5_n184 ) , .A1( u1_u10_u5_n194 ) );
  XOR2_X1 u1_u11_U22 (.B( u1_K12_34 ) , .A( u1_R10_23 ) , .Z( u1_u11_X_34 ) );
  XOR2_X1 u1_u11_U23 (.B( u1_K12_33 ) , .A( u1_R10_22 ) , .Z( u1_u11_X_33 ) );
  INV_X1 u1_u11_u5_U10 (.A( u1_u11_u5_n121 ) , .ZN( u1_u11_u5_n177 ) );
  NOR3_X1 u1_u11_u5_U100 (.A3( u1_u11_u5_n141 ) , .A1( u1_u11_u5_n142 ) , .ZN( u1_u11_u5_n143 ) , .A2( u1_u11_u5_n191 ) );
  NAND4_X1 u1_u11_u5_U101 (.ZN( u1_out11_4 ) , .A4( u1_u11_u5_n112 ) , .A2( u1_u11_u5_n113 ) , .A1( u1_u11_u5_n114 ) , .A3( u1_u11_u5_n195 ) );
  AOI211_X1 u1_u11_u5_U102 (.A( u1_u11_u5_n110 ) , .C1( u1_u11_u5_n111 ) , .ZN( u1_u11_u5_n112 ) , .B( u1_u11_u5_n118 ) , .C2( u1_u11_u5_n177 ) );
  AOI222_X1 u1_u11_u5_U103 (.ZN( u1_u11_u5_n113 ) , .A1( u1_u11_u5_n131 ) , .C1( u1_u11_u5_n148 ) , .B2( u1_u11_u5_n174 ) , .C2( u1_u11_u5_n178 ) , .A2( u1_u11_u5_n179 ) , .B1( u1_u11_u5_n99 ) );
  NAND3_X1 u1_u11_u5_U104 (.A2( u1_u11_u5_n154 ) , .A3( u1_u11_u5_n158 ) , .A1( u1_u11_u5_n161 ) , .ZN( u1_u11_u5_n99 ) );
  NOR2_X1 u1_u11_u5_U11 (.ZN( u1_u11_u5_n160 ) , .A2( u1_u11_u5_n173 ) , .A1( u1_u11_u5_n177 ) );
  INV_X1 u1_u11_u5_U12 (.A( u1_u11_u5_n150 ) , .ZN( u1_u11_u5_n174 ) );
  AOI21_X1 u1_u11_u5_U13 (.A( u1_u11_u5_n160 ) , .B2( u1_u11_u5_n161 ) , .ZN( u1_u11_u5_n162 ) , .B1( u1_u11_u5_n192 ) );
  INV_X1 u1_u11_u5_U14 (.A( u1_u11_u5_n159 ) , .ZN( u1_u11_u5_n192 ) );
  AOI21_X1 u1_u11_u5_U15 (.A( u1_u11_u5_n156 ) , .B2( u1_u11_u5_n157 ) , .B1( u1_u11_u5_n158 ) , .ZN( u1_u11_u5_n163 ) );
  AOI21_X1 u1_u11_u5_U16 (.B2( u1_u11_u5_n139 ) , .B1( u1_u11_u5_n140 ) , .ZN( u1_u11_u5_n141 ) , .A( u1_u11_u5_n150 ) );
  OAI21_X1 u1_u11_u5_U17 (.A( u1_u11_u5_n133 ) , .B2( u1_u11_u5_n134 ) , .B1( u1_u11_u5_n135 ) , .ZN( u1_u11_u5_n142 ) );
  OAI21_X1 u1_u11_u5_U18 (.ZN( u1_u11_u5_n133 ) , .B2( u1_u11_u5_n147 ) , .A( u1_u11_u5_n173 ) , .B1( u1_u11_u5_n188 ) );
  NAND2_X1 u1_u11_u5_U19 (.A2( u1_u11_u5_n119 ) , .A1( u1_u11_u5_n123 ) , .ZN( u1_u11_u5_n137 ) );
  INV_X1 u1_u11_u5_U20 (.A( u1_u11_u5_n155 ) , .ZN( u1_u11_u5_n194 ) );
  NAND2_X1 u1_u11_u5_U21 (.A1( u1_u11_u5_n121 ) , .ZN( u1_u11_u5_n132 ) , .A2( u1_u11_u5_n172 ) );
  NAND2_X1 u1_u11_u5_U22 (.A2( u1_u11_u5_n122 ) , .ZN( u1_u11_u5_n136 ) , .A1( u1_u11_u5_n154 ) );
  NAND2_X1 u1_u11_u5_U23 (.A2( u1_u11_u5_n119 ) , .A1( u1_u11_u5_n120 ) , .ZN( u1_u11_u5_n159 ) );
  INV_X1 u1_u11_u5_U24 (.A( u1_u11_u5_n156 ) , .ZN( u1_u11_u5_n175 ) );
  INV_X1 u1_u11_u5_U25 (.A( u1_u11_u5_n158 ) , .ZN( u1_u11_u5_n188 ) );
  INV_X1 u1_u11_u5_U26 (.A( u1_u11_u5_n152 ) , .ZN( u1_u11_u5_n179 ) );
  INV_X1 u1_u11_u5_U27 (.A( u1_u11_u5_n140 ) , .ZN( u1_u11_u5_n182 ) );
  INV_X1 u1_u11_u5_U28 (.A( u1_u11_u5_n151 ) , .ZN( u1_u11_u5_n183 ) );
  INV_X1 u1_u11_u5_U29 (.A( u1_u11_u5_n123 ) , .ZN( u1_u11_u5_n185 ) );
  NOR2_X1 u1_u11_u5_U3 (.ZN( u1_u11_u5_n134 ) , .A1( u1_u11_u5_n183 ) , .A2( u1_u11_u5_n190 ) );
  INV_X1 u1_u11_u5_U30 (.A( u1_u11_u5_n161 ) , .ZN( u1_u11_u5_n184 ) );
  INV_X1 u1_u11_u5_U31 (.A( u1_u11_u5_n139 ) , .ZN( u1_u11_u5_n189 ) );
  INV_X1 u1_u11_u5_U32 (.A( u1_u11_u5_n157 ) , .ZN( u1_u11_u5_n190 ) );
  INV_X1 u1_u11_u5_U33 (.A( u1_u11_u5_n120 ) , .ZN( u1_u11_u5_n193 ) );
  NAND2_X1 u1_u11_u5_U34 (.ZN( u1_u11_u5_n111 ) , .A1( u1_u11_u5_n140 ) , .A2( u1_u11_u5_n155 ) );
  NOR2_X1 u1_u11_u5_U35 (.ZN( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n170 ) , .A2( u1_u11_u5_n180 ) );
  INV_X1 u1_u11_u5_U36 (.A( u1_u11_u5_n117 ) , .ZN( u1_u11_u5_n196 ) );
  OAI221_X1 u1_u11_u5_U37 (.A( u1_u11_u5_n116 ) , .ZN( u1_u11_u5_n117 ) , .B2( u1_u11_u5_n119 ) , .C1( u1_u11_u5_n153 ) , .C2( u1_u11_u5_n158 ) , .B1( u1_u11_u5_n172 ) );
  AOI222_X1 u1_u11_u5_U38 (.ZN( u1_u11_u5_n116 ) , .B2( u1_u11_u5_n145 ) , .C1( u1_u11_u5_n148 ) , .A2( u1_u11_u5_n174 ) , .C2( u1_u11_u5_n177 ) , .B1( u1_u11_u5_n187 ) , .A1( u1_u11_u5_n193 ) );
  INV_X1 u1_u11_u5_U39 (.A( u1_u11_u5_n115 ) , .ZN( u1_u11_u5_n187 ) );
  INV_X1 u1_u11_u5_U4 (.A( u1_u11_u5_n138 ) , .ZN( u1_u11_u5_n191 ) );
  AOI22_X1 u1_u11_u5_U40 (.B2( u1_u11_u5_n131 ) , .A2( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n169 ) , .B1( u1_u11_u5_n174 ) , .A1( u1_u11_u5_n185 ) );
  NOR2_X1 u1_u11_u5_U41 (.A1( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n150 ) , .A2( u1_u11_u5_n173 ) );
  AOI21_X1 u1_u11_u5_U42 (.A( u1_u11_u5_n118 ) , .B2( u1_u11_u5_n145 ) , .ZN( u1_u11_u5_n168 ) , .B1( u1_u11_u5_n186 ) );
  INV_X1 u1_u11_u5_U43 (.A( u1_u11_u5_n122 ) , .ZN( u1_u11_u5_n186 ) );
  NOR2_X1 u1_u11_u5_U44 (.A1( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n152 ) , .A2( u1_u11_u5_n176 ) );
  NOR2_X1 u1_u11_u5_U45 (.A1( u1_u11_u5_n115 ) , .ZN( u1_u11_u5_n118 ) , .A2( u1_u11_u5_n153 ) );
  NOR2_X1 u1_u11_u5_U46 (.A2( u1_u11_u5_n145 ) , .ZN( u1_u11_u5_n156 ) , .A1( u1_u11_u5_n174 ) );
  NOR2_X1 u1_u11_u5_U47 (.ZN( u1_u11_u5_n121 ) , .A2( u1_u11_u5_n145 ) , .A1( u1_u11_u5_n176 ) );
  AOI22_X1 u1_u11_u5_U48 (.ZN( u1_u11_u5_n114 ) , .A2( u1_u11_u5_n137 ) , .A1( u1_u11_u5_n145 ) , .B2( u1_u11_u5_n175 ) , .B1( u1_u11_u5_n193 ) );
  OAI211_X1 u1_u11_u5_U49 (.B( u1_u11_u5_n124 ) , .A( u1_u11_u5_n125 ) , .C2( u1_u11_u5_n126 ) , .C1( u1_u11_u5_n127 ) , .ZN( u1_u11_u5_n128 ) );
  OAI21_X1 u1_u11_u5_U5 (.B2( u1_u11_u5_n136 ) , .B1( u1_u11_u5_n137 ) , .ZN( u1_u11_u5_n138 ) , .A( u1_u11_u5_n177 ) );
  OAI21_X1 u1_u11_u5_U50 (.ZN( u1_u11_u5_n124 ) , .A( u1_u11_u5_n177 ) , .B2( u1_u11_u5_n183 ) , .B1( u1_u11_u5_n189 ) );
  NOR3_X1 u1_u11_u5_U51 (.ZN( u1_u11_u5_n127 ) , .A1( u1_u11_u5_n136 ) , .A3( u1_u11_u5_n148 ) , .A2( u1_u11_u5_n182 ) );
  OAI21_X1 u1_u11_u5_U52 (.ZN( u1_u11_u5_n125 ) , .A( u1_u11_u5_n174 ) , .B2( u1_u11_u5_n185 ) , .B1( u1_u11_u5_n190 ) );
  AOI21_X1 u1_u11_u5_U53 (.A( u1_u11_u5_n153 ) , .B2( u1_u11_u5_n154 ) , .B1( u1_u11_u5_n155 ) , .ZN( u1_u11_u5_n164 ) );
  AOI21_X1 u1_u11_u5_U54 (.ZN( u1_u11_u5_n110 ) , .B1( u1_u11_u5_n122 ) , .B2( u1_u11_u5_n139 ) , .A( u1_u11_u5_n153 ) );
  INV_X1 u1_u11_u5_U55 (.A( u1_u11_u5_n153 ) , .ZN( u1_u11_u5_n176 ) );
  INV_X1 u1_u11_u5_U56 (.A( u1_u11_u5_n126 ) , .ZN( u1_u11_u5_n173 ) );
  AND2_X1 u1_u11_u5_U57 (.A2( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n107 ) , .ZN( u1_u11_u5_n147 ) );
  AND2_X1 u1_u11_u5_U58 (.A2( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n108 ) , .ZN( u1_u11_u5_n148 ) );
  NAND2_X1 u1_u11_u5_U59 (.A1( u1_u11_u5_n105 ) , .A2( u1_u11_u5_n106 ) , .ZN( u1_u11_u5_n158 ) );
  INV_X1 u1_u11_u5_U6 (.A( u1_u11_u5_n135 ) , .ZN( u1_u11_u5_n178 ) );
  NAND2_X1 u1_u11_u5_U60 (.A2( u1_u11_u5_n108 ) , .A1( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n139 ) );
  NAND2_X1 u1_u11_u5_U61 (.A1( u1_u11_u5_n106 ) , .A2( u1_u11_u5_n108 ) , .ZN( u1_u11_u5_n119 ) );
  NAND2_X1 u1_u11_u5_U62 (.A2( u1_u11_u5_n103 ) , .A1( u1_u11_u5_n105 ) , .ZN( u1_u11_u5_n140 ) );
  NAND2_X1 u1_u11_u5_U63 (.A2( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n105 ) , .ZN( u1_u11_u5_n155 ) );
  NAND2_X1 u1_u11_u5_U64 (.A2( u1_u11_u5_n106 ) , .A1( u1_u11_u5_n107 ) , .ZN( u1_u11_u5_n122 ) );
  NAND2_X1 u1_u11_u5_U65 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n106 ) , .ZN( u1_u11_u5_n115 ) );
  NAND2_X1 u1_u11_u5_U66 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n103 ) , .ZN( u1_u11_u5_n161 ) );
  NAND2_X1 u1_u11_u5_U67 (.A1( u1_u11_u5_n105 ) , .A2( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n154 ) );
  INV_X1 u1_u11_u5_U68 (.A( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n172 ) );
  NAND2_X1 u1_u11_u5_U69 (.A1( u1_u11_u5_n103 ) , .A2( u1_u11_u5_n108 ) , .ZN( u1_u11_u5_n123 ) );
  OAI22_X1 u1_u11_u5_U7 (.B2( u1_u11_u5_n149 ) , .B1( u1_u11_u5_n150 ) , .A2( u1_u11_u5_n151 ) , .A1( u1_u11_u5_n152 ) , .ZN( u1_u11_u5_n165 ) );
  NAND2_X1 u1_u11_u5_U70 (.A2( u1_u11_u5_n103 ) , .A1( u1_u11_u5_n107 ) , .ZN( u1_u11_u5_n151 ) );
  NAND2_X1 u1_u11_u5_U71 (.A2( u1_u11_u5_n107 ) , .A1( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n120 ) );
  NAND2_X1 u1_u11_u5_U72 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n109 ) , .ZN( u1_u11_u5_n157 ) );
  AND2_X1 u1_u11_u5_U73 (.A2( u1_u11_u5_n100 ) , .A1( u1_u11_u5_n104 ) , .ZN( u1_u11_u5_n131 ) );
  INV_X1 u1_u11_u5_U74 (.A( u1_u11_u5_n102 ) , .ZN( u1_u11_u5_n195 ) );
  OAI221_X1 u1_u11_u5_U75 (.A( u1_u11_u5_n101 ) , .ZN( u1_u11_u5_n102 ) , .C2( u1_u11_u5_n115 ) , .C1( u1_u11_u5_n126 ) , .B1( u1_u11_u5_n134 ) , .B2( u1_u11_u5_n160 ) );
  OAI21_X1 u1_u11_u5_U76 (.ZN( u1_u11_u5_n101 ) , .B1( u1_u11_u5_n137 ) , .A( u1_u11_u5_n146 ) , .B2( u1_u11_u5_n147 ) );
  NOR2_X1 u1_u11_u5_U77 (.A2( u1_u11_X_34 ) , .A1( u1_u11_X_35 ) , .ZN( u1_u11_u5_n145 ) );
  NOR2_X1 u1_u11_u5_U78 (.A2( u1_u11_X_34 ) , .ZN( u1_u11_u5_n146 ) , .A1( u1_u11_u5_n171 ) );
  NOR2_X1 u1_u11_u5_U79 (.A2( u1_u11_X_31 ) , .A1( u1_u11_X_32 ) , .ZN( u1_u11_u5_n103 ) );
  NOR3_X1 u1_u11_u5_U8 (.A2( u1_u11_u5_n147 ) , .A1( u1_u11_u5_n148 ) , .ZN( u1_u11_u5_n149 ) , .A3( u1_u11_u5_n194 ) );
  NOR2_X1 u1_u11_u5_U80 (.A2( u1_u11_X_36 ) , .ZN( u1_u11_u5_n105 ) , .A1( u1_u11_u5_n180 ) );
  NOR2_X1 u1_u11_u5_U81 (.A2( u1_u11_X_33 ) , .ZN( u1_u11_u5_n108 ) , .A1( u1_u11_u5_n170 ) );
  NOR2_X1 u1_u11_u5_U82 (.A2( u1_u11_X_33 ) , .A1( u1_u11_X_36 ) , .ZN( u1_u11_u5_n107 ) );
  NOR2_X1 u1_u11_u5_U83 (.A2( u1_u11_X_31 ) , .ZN( u1_u11_u5_n104 ) , .A1( u1_u11_u5_n181 ) );
  NAND2_X1 u1_u11_u5_U84 (.A2( u1_u11_X_34 ) , .A1( u1_u11_X_35 ) , .ZN( u1_u11_u5_n153 ) );
  NAND2_X1 u1_u11_u5_U85 (.A1( u1_u11_X_34 ) , .ZN( u1_u11_u5_n126 ) , .A2( u1_u11_u5_n171 ) );
  AND2_X1 u1_u11_u5_U86 (.A1( u1_u11_X_31 ) , .A2( u1_u11_X_32 ) , .ZN( u1_u11_u5_n106 ) );
  AND2_X1 u1_u11_u5_U87 (.A1( u1_u11_X_31 ) , .ZN( u1_u11_u5_n109 ) , .A2( u1_u11_u5_n181 ) );
  INV_X1 u1_u11_u5_U88 (.A( u1_u11_X_33 ) , .ZN( u1_u11_u5_n180 ) );
  INV_X1 u1_u11_u5_U89 (.A( u1_u11_X_35 ) , .ZN( u1_u11_u5_n171 ) );
  NOR2_X1 u1_u11_u5_U9 (.ZN( u1_u11_u5_n135 ) , .A1( u1_u11_u5_n173 ) , .A2( u1_u11_u5_n176 ) );
  INV_X1 u1_u11_u5_U90 (.A( u1_u11_X_36 ) , .ZN( u1_u11_u5_n170 ) );
  INV_X1 u1_u11_u5_U91 (.A( u1_u11_X_32 ) , .ZN( u1_u11_u5_n181 ) );
  NAND4_X1 u1_u11_u5_U92 (.ZN( u1_out11_29 ) , .A4( u1_u11_u5_n129 ) , .A3( u1_u11_u5_n130 ) , .A2( u1_u11_u5_n168 ) , .A1( u1_u11_u5_n196 ) );
  AOI221_X1 u1_u11_u5_U93 (.A( u1_u11_u5_n128 ) , .ZN( u1_u11_u5_n129 ) , .C2( u1_u11_u5_n132 ) , .B2( u1_u11_u5_n159 ) , .B1( u1_u11_u5_n176 ) , .C1( u1_u11_u5_n184 ) );
  AOI222_X1 u1_u11_u5_U94 (.ZN( u1_u11_u5_n130 ) , .A2( u1_u11_u5_n146 ) , .B1( u1_u11_u5_n147 ) , .C2( u1_u11_u5_n175 ) , .B2( u1_u11_u5_n179 ) , .A1( u1_u11_u5_n188 ) , .C1( u1_u11_u5_n194 ) );
  NAND4_X1 u1_u11_u5_U95 (.ZN( u1_out11_19 ) , .A4( u1_u11_u5_n166 ) , .A3( u1_u11_u5_n167 ) , .A2( u1_u11_u5_n168 ) , .A1( u1_u11_u5_n169 ) );
  AOI22_X1 u1_u11_u5_U96 (.B2( u1_u11_u5_n145 ) , .A2( u1_u11_u5_n146 ) , .ZN( u1_u11_u5_n167 ) , .B1( u1_u11_u5_n182 ) , .A1( u1_u11_u5_n189 ) );
  NOR4_X1 u1_u11_u5_U97 (.A4( u1_u11_u5_n162 ) , .A3( u1_u11_u5_n163 ) , .A2( u1_u11_u5_n164 ) , .A1( u1_u11_u5_n165 ) , .ZN( u1_u11_u5_n166 ) );
  NAND4_X1 u1_u11_u5_U98 (.ZN( u1_out11_11 ) , .A4( u1_u11_u5_n143 ) , .A3( u1_u11_u5_n144 ) , .A2( u1_u11_u5_n169 ) , .A1( u1_u11_u5_n196 ) );
  AOI22_X1 u1_u11_u5_U99 (.A2( u1_u11_u5_n132 ) , .ZN( u1_u11_u5_n144 ) , .B2( u1_u11_u5_n145 ) , .B1( u1_u11_u5_n184 ) , .A1( u1_u11_u5_n194 ) );
  XOR2_X1 u1_u12_U15 (.B( u1_K13_40 ) , .A( u1_R11_27 ) , .Z( u1_u12_X_40 ) );
  XOR2_X1 u1_u12_U17 (.B( u1_K13_39 ) , .A( u1_R11_26 ) , .Z( u1_u12_X_39 ) );
  AOI22_X1 u1_u12_u6_U10 (.A2( u1_u12_u6_n151 ) , .B2( u1_u12_u6_n161 ) , .A1( u1_u12_u6_n167 ) , .B1( u1_u12_u6_n170 ) , .ZN( u1_u12_u6_n89 ) );
  AOI21_X1 u1_u12_u6_U11 (.B1( u1_u12_u6_n107 ) , .B2( u1_u12_u6_n132 ) , .A( u1_u12_u6_n158 ) , .ZN( u1_u12_u6_n88 ) );
  AOI21_X1 u1_u12_u6_U12 (.B2( u1_u12_u6_n147 ) , .B1( u1_u12_u6_n148 ) , .ZN( u1_u12_u6_n149 ) , .A( u1_u12_u6_n158 ) );
  AOI21_X1 u1_u12_u6_U13 (.ZN( u1_u12_u6_n106 ) , .A( u1_u12_u6_n142 ) , .B2( u1_u12_u6_n159 ) , .B1( u1_u12_u6_n164 ) );
  INV_X1 u1_u12_u6_U14 (.A( u1_u12_u6_n155 ) , .ZN( u1_u12_u6_n161 ) );
  INV_X1 u1_u12_u6_U15 (.A( u1_u12_u6_n128 ) , .ZN( u1_u12_u6_n164 ) );
  NAND2_X1 u1_u12_u6_U16 (.ZN( u1_u12_u6_n110 ) , .A1( u1_u12_u6_n122 ) , .A2( u1_u12_u6_n129 ) );
  NAND2_X1 u1_u12_u6_U17 (.ZN( u1_u12_u6_n124 ) , .A2( u1_u12_u6_n146 ) , .A1( u1_u12_u6_n148 ) );
  INV_X1 u1_u12_u6_U18 (.A( u1_u12_u6_n132 ) , .ZN( u1_u12_u6_n171 ) );
  AND2_X1 u1_u12_u6_U19 (.A1( u1_u12_u6_n100 ) , .ZN( u1_u12_u6_n130 ) , .A2( u1_u12_u6_n147 ) );
  INV_X1 u1_u12_u6_U20 (.A( u1_u12_u6_n127 ) , .ZN( u1_u12_u6_n173 ) );
  INV_X1 u1_u12_u6_U21 (.A( u1_u12_u6_n121 ) , .ZN( u1_u12_u6_n167 ) );
  INV_X1 u1_u12_u6_U22 (.A( u1_u12_u6_n100 ) , .ZN( u1_u12_u6_n169 ) );
  INV_X1 u1_u12_u6_U23 (.A( u1_u12_u6_n123 ) , .ZN( u1_u12_u6_n170 ) );
  INV_X1 u1_u12_u6_U24 (.A( u1_u12_u6_n113 ) , .ZN( u1_u12_u6_n168 ) );
  AND2_X1 u1_u12_u6_U25 (.A1( u1_u12_u6_n107 ) , .A2( u1_u12_u6_n119 ) , .ZN( u1_u12_u6_n133 ) );
  AND2_X1 u1_u12_u6_U26 (.A2( u1_u12_u6_n121 ) , .A1( u1_u12_u6_n122 ) , .ZN( u1_u12_u6_n131 ) );
  AND3_X1 u1_u12_u6_U27 (.ZN( u1_u12_u6_n120 ) , .A2( u1_u12_u6_n127 ) , .A1( u1_u12_u6_n132 ) , .A3( u1_u12_u6_n145 ) );
  INV_X1 u1_u12_u6_U28 (.A( u1_u12_u6_n146 ) , .ZN( u1_u12_u6_n163 ) );
  AOI222_X1 u1_u12_u6_U29 (.ZN( u1_u12_u6_n114 ) , .A1( u1_u12_u6_n118 ) , .A2( u1_u12_u6_n126 ) , .B2( u1_u12_u6_n151 ) , .C2( u1_u12_u6_n159 ) , .C1( u1_u12_u6_n168 ) , .B1( u1_u12_u6_n169 ) );
  INV_X1 u1_u12_u6_U3 (.A( u1_u12_u6_n110 ) , .ZN( u1_u12_u6_n166 ) );
  NOR2_X1 u1_u12_u6_U30 (.A1( u1_u12_u6_n162 ) , .A2( u1_u12_u6_n165 ) , .ZN( u1_u12_u6_n98 ) );
  AOI211_X1 u1_u12_u6_U31 (.B( u1_u12_u6_n134 ) , .A( u1_u12_u6_n135 ) , .C1( u1_u12_u6_n136 ) , .ZN( u1_u12_u6_n137 ) , .C2( u1_u12_u6_n151 ) );
  AOI21_X1 u1_u12_u6_U32 (.B2( u1_u12_u6_n132 ) , .B1( u1_u12_u6_n133 ) , .ZN( u1_u12_u6_n134 ) , .A( u1_u12_u6_n158 ) );
  AOI21_X1 u1_u12_u6_U33 (.B1( u1_u12_u6_n131 ) , .ZN( u1_u12_u6_n135 ) , .A( u1_u12_u6_n144 ) , .B2( u1_u12_u6_n146 ) );
  NAND4_X1 u1_u12_u6_U34 (.A4( u1_u12_u6_n127 ) , .A3( u1_u12_u6_n128 ) , .A2( u1_u12_u6_n129 ) , .A1( u1_u12_u6_n130 ) , .ZN( u1_u12_u6_n136 ) );
  NAND2_X1 u1_u12_u6_U35 (.A1( u1_u12_u6_n144 ) , .ZN( u1_u12_u6_n151 ) , .A2( u1_u12_u6_n158 ) );
  NAND2_X1 u1_u12_u6_U36 (.ZN( u1_u12_u6_n132 ) , .A1( u1_u12_u6_n91 ) , .A2( u1_u12_u6_n97 ) );
  AOI22_X1 u1_u12_u6_U37 (.B2( u1_u12_u6_n110 ) , .B1( u1_u12_u6_n111 ) , .A1( u1_u12_u6_n112 ) , .ZN( u1_u12_u6_n115 ) , .A2( u1_u12_u6_n161 ) );
  NAND4_X1 u1_u12_u6_U38 (.A3( u1_u12_u6_n109 ) , .ZN( u1_u12_u6_n112 ) , .A4( u1_u12_u6_n132 ) , .A2( u1_u12_u6_n147 ) , .A1( u1_u12_u6_n166 ) );
  NOR2_X1 u1_u12_u6_U39 (.ZN( u1_u12_u6_n109 ) , .A1( u1_u12_u6_n170 ) , .A2( u1_u12_u6_n173 ) );
  INV_X1 u1_u12_u6_U4 (.A( u1_u12_u6_n142 ) , .ZN( u1_u12_u6_n174 ) );
  NOR2_X1 u1_u12_u6_U40 (.A2( u1_u12_u6_n126 ) , .ZN( u1_u12_u6_n155 ) , .A1( u1_u12_u6_n160 ) );
  NAND2_X1 u1_u12_u6_U41 (.ZN( u1_u12_u6_n146 ) , .A2( u1_u12_u6_n94 ) , .A1( u1_u12_u6_n99 ) );
  AOI21_X1 u1_u12_u6_U42 (.A( u1_u12_u6_n144 ) , .B2( u1_u12_u6_n145 ) , .B1( u1_u12_u6_n146 ) , .ZN( u1_u12_u6_n150 ) );
  INV_X1 u1_u12_u6_U43 (.A( u1_u12_u6_n111 ) , .ZN( u1_u12_u6_n158 ) );
  NAND2_X1 u1_u12_u6_U44 (.ZN( u1_u12_u6_n127 ) , .A1( u1_u12_u6_n91 ) , .A2( u1_u12_u6_n92 ) );
  NAND2_X1 u1_u12_u6_U45 (.ZN( u1_u12_u6_n129 ) , .A2( u1_u12_u6_n95 ) , .A1( u1_u12_u6_n96 ) );
  INV_X1 u1_u12_u6_U46 (.A( u1_u12_u6_n144 ) , .ZN( u1_u12_u6_n159 ) );
  NAND2_X1 u1_u12_u6_U47 (.ZN( u1_u12_u6_n145 ) , .A2( u1_u12_u6_n97 ) , .A1( u1_u12_u6_n98 ) );
  NAND2_X1 u1_u12_u6_U48 (.ZN( u1_u12_u6_n148 ) , .A2( u1_u12_u6_n92 ) , .A1( u1_u12_u6_n94 ) );
  NAND2_X1 u1_u12_u6_U49 (.ZN( u1_u12_u6_n108 ) , .A2( u1_u12_u6_n139 ) , .A1( u1_u12_u6_n144 ) );
  NAND2_X1 u1_u12_u6_U5 (.A2( u1_u12_u6_n143 ) , .ZN( u1_u12_u6_n152 ) , .A1( u1_u12_u6_n166 ) );
  NAND2_X1 u1_u12_u6_U50 (.ZN( u1_u12_u6_n121 ) , .A2( u1_u12_u6_n95 ) , .A1( u1_u12_u6_n97 ) );
  NAND2_X1 u1_u12_u6_U51 (.ZN( u1_u12_u6_n107 ) , .A2( u1_u12_u6_n92 ) , .A1( u1_u12_u6_n95 ) );
  AND2_X1 u1_u12_u6_U52 (.ZN( u1_u12_u6_n118 ) , .A2( u1_u12_u6_n91 ) , .A1( u1_u12_u6_n99 ) );
  NAND2_X1 u1_u12_u6_U53 (.ZN( u1_u12_u6_n147 ) , .A2( u1_u12_u6_n98 ) , .A1( u1_u12_u6_n99 ) );
  NAND2_X1 u1_u12_u6_U54 (.ZN( u1_u12_u6_n128 ) , .A1( u1_u12_u6_n94 ) , .A2( u1_u12_u6_n96 ) );
  NAND2_X1 u1_u12_u6_U55 (.ZN( u1_u12_u6_n119 ) , .A2( u1_u12_u6_n95 ) , .A1( u1_u12_u6_n99 ) );
  NAND2_X1 u1_u12_u6_U56 (.ZN( u1_u12_u6_n123 ) , .A2( u1_u12_u6_n91 ) , .A1( u1_u12_u6_n96 ) );
  NAND2_X1 u1_u12_u6_U57 (.ZN( u1_u12_u6_n100 ) , .A2( u1_u12_u6_n92 ) , .A1( u1_u12_u6_n98 ) );
  NAND2_X1 u1_u12_u6_U58 (.ZN( u1_u12_u6_n122 ) , .A1( u1_u12_u6_n94 ) , .A2( u1_u12_u6_n97 ) );
  INV_X1 u1_u12_u6_U59 (.A( u1_u12_u6_n139 ) , .ZN( u1_u12_u6_n160 ) );
  AOI22_X1 u1_u12_u6_U6 (.B2( u1_u12_u6_n101 ) , .A1( u1_u12_u6_n102 ) , .ZN( u1_u12_u6_n103 ) , .B1( u1_u12_u6_n160 ) , .A2( u1_u12_u6_n161 ) );
  NAND2_X1 u1_u12_u6_U60 (.ZN( u1_u12_u6_n113 ) , .A1( u1_u12_u6_n96 ) , .A2( u1_u12_u6_n98 ) );
  NOR2_X1 u1_u12_u6_U61 (.A2( u1_u12_X_40 ) , .A1( u1_u12_X_41 ) , .ZN( u1_u12_u6_n126 ) );
  NOR2_X1 u1_u12_u6_U62 (.A2( u1_u12_X_39 ) , .A1( u1_u12_X_42 ) , .ZN( u1_u12_u6_n92 ) );
  NOR2_X1 u1_u12_u6_U63 (.A2( u1_u12_X_39 ) , .A1( u1_u12_u6_n156 ) , .ZN( u1_u12_u6_n97 ) );
  NOR2_X1 u1_u12_u6_U64 (.A2( u1_u12_X_38 ) , .A1( u1_u12_u6_n165 ) , .ZN( u1_u12_u6_n95 ) );
  NOR2_X1 u1_u12_u6_U65 (.A2( u1_u12_X_41 ) , .ZN( u1_u12_u6_n111 ) , .A1( u1_u12_u6_n157 ) );
  NOR2_X1 u1_u12_u6_U66 (.A2( u1_u12_X_37 ) , .A1( u1_u12_u6_n162 ) , .ZN( u1_u12_u6_n94 ) );
  NOR2_X1 u1_u12_u6_U67 (.A2( u1_u12_X_37 ) , .A1( u1_u12_X_38 ) , .ZN( u1_u12_u6_n91 ) );
  NAND2_X1 u1_u12_u6_U68 (.A1( u1_u12_X_41 ) , .ZN( u1_u12_u6_n144 ) , .A2( u1_u12_u6_n157 ) );
  NAND2_X1 u1_u12_u6_U69 (.A2( u1_u12_X_40 ) , .A1( u1_u12_X_41 ) , .ZN( u1_u12_u6_n139 ) );
  NOR2_X1 u1_u12_u6_U7 (.A1( u1_u12_u6_n118 ) , .ZN( u1_u12_u6_n143 ) , .A2( u1_u12_u6_n168 ) );
  AND2_X1 u1_u12_u6_U70 (.A1( u1_u12_X_39 ) , .A2( u1_u12_u6_n156 ) , .ZN( u1_u12_u6_n96 ) );
  AND2_X1 u1_u12_u6_U71 (.A1( u1_u12_X_39 ) , .A2( u1_u12_X_42 ) , .ZN( u1_u12_u6_n99 ) );
  INV_X1 u1_u12_u6_U72 (.A( u1_u12_X_40 ) , .ZN( u1_u12_u6_n157 ) );
  INV_X1 u1_u12_u6_U73 (.A( u1_u12_X_37 ) , .ZN( u1_u12_u6_n165 ) );
  INV_X1 u1_u12_u6_U74 (.A( u1_u12_X_38 ) , .ZN( u1_u12_u6_n162 ) );
  INV_X1 u1_u12_u6_U75 (.A( u1_u12_X_42 ) , .ZN( u1_u12_u6_n156 ) );
  NAND4_X1 u1_u12_u6_U76 (.ZN( u1_out12_32 ) , .A4( u1_u12_u6_n103 ) , .A3( u1_u12_u6_n104 ) , .A2( u1_u12_u6_n105 ) , .A1( u1_u12_u6_n106 ) );
  AOI22_X1 u1_u12_u6_U77 (.ZN( u1_u12_u6_n105 ) , .A2( u1_u12_u6_n108 ) , .A1( u1_u12_u6_n118 ) , .B2( u1_u12_u6_n126 ) , .B1( u1_u12_u6_n171 ) );
  AOI22_X1 u1_u12_u6_U78 (.ZN( u1_u12_u6_n104 ) , .A1( u1_u12_u6_n111 ) , .B1( u1_u12_u6_n124 ) , .B2( u1_u12_u6_n151 ) , .A2( u1_u12_u6_n93 ) );
  NAND4_X1 u1_u12_u6_U79 (.ZN( u1_out12_12 ) , .A4( u1_u12_u6_n114 ) , .A3( u1_u12_u6_n115 ) , .A2( u1_u12_u6_n116 ) , .A1( u1_u12_u6_n117 ) );
  INV_X1 u1_u12_u6_U8 (.ZN( u1_u12_u6_n172 ) , .A( u1_u12_u6_n88 ) );
  OAI22_X1 u1_u12_u6_U80 (.B2( u1_u12_u6_n111 ) , .ZN( u1_u12_u6_n116 ) , .B1( u1_u12_u6_n126 ) , .A2( u1_u12_u6_n164 ) , .A1( u1_u12_u6_n167 ) );
  OAI21_X1 u1_u12_u6_U81 (.A( u1_u12_u6_n108 ) , .ZN( u1_u12_u6_n117 ) , .B2( u1_u12_u6_n141 ) , .B1( u1_u12_u6_n163 ) );
  OAI211_X1 u1_u12_u6_U82 (.ZN( u1_out12_22 ) , .B( u1_u12_u6_n137 ) , .A( u1_u12_u6_n138 ) , .C2( u1_u12_u6_n139 ) , .C1( u1_u12_u6_n140 ) );
  AOI22_X1 u1_u12_u6_U83 (.B1( u1_u12_u6_n124 ) , .A2( u1_u12_u6_n125 ) , .A1( u1_u12_u6_n126 ) , .ZN( u1_u12_u6_n138 ) , .B2( u1_u12_u6_n161 ) );
  AND4_X1 u1_u12_u6_U84 (.A3( u1_u12_u6_n119 ) , .A1( u1_u12_u6_n120 ) , .A4( u1_u12_u6_n129 ) , .ZN( u1_u12_u6_n140 ) , .A2( u1_u12_u6_n143 ) );
  OAI211_X1 u1_u12_u6_U85 (.ZN( u1_out12_7 ) , .B( u1_u12_u6_n153 ) , .C2( u1_u12_u6_n154 ) , .C1( u1_u12_u6_n155 ) , .A( u1_u12_u6_n174 ) );
  NOR3_X1 u1_u12_u6_U86 (.A1( u1_u12_u6_n141 ) , .ZN( u1_u12_u6_n154 ) , .A3( u1_u12_u6_n164 ) , .A2( u1_u12_u6_n171 ) );
  AOI211_X1 u1_u12_u6_U87 (.B( u1_u12_u6_n149 ) , .A( u1_u12_u6_n150 ) , .C2( u1_u12_u6_n151 ) , .C1( u1_u12_u6_n152 ) , .ZN( u1_u12_u6_n153 ) );
  NAND3_X1 u1_u12_u6_U88 (.A2( u1_u12_u6_n123 ) , .ZN( u1_u12_u6_n125 ) , .A1( u1_u12_u6_n130 ) , .A3( u1_u12_u6_n131 ) );
  NAND3_X1 u1_u12_u6_U89 (.A3( u1_u12_u6_n133 ) , .ZN( u1_u12_u6_n141 ) , .A1( u1_u12_u6_n145 ) , .A2( u1_u12_u6_n148 ) );
  OAI21_X1 u1_u12_u6_U9 (.A( u1_u12_u6_n159 ) , .B1( u1_u12_u6_n169 ) , .B2( u1_u12_u6_n173 ) , .ZN( u1_u12_u6_n90 ) );
  NAND3_X1 u1_u12_u6_U90 (.ZN( u1_u12_u6_n101 ) , .A3( u1_u12_u6_n107 ) , .A2( u1_u12_u6_n121 ) , .A1( u1_u12_u6_n127 ) );
  NAND3_X1 u1_u12_u6_U91 (.ZN( u1_u12_u6_n102 ) , .A3( u1_u12_u6_n130 ) , .A2( u1_u12_u6_n145 ) , .A1( u1_u12_u6_n166 ) );
  NAND3_X1 u1_u12_u6_U92 (.A3( u1_u12_u6_n113 ) , .A1( u1_u12_u6_n119 ) , .A2( u1_u12_u6_n123 ) , .ZN( u1_u12_u6_n93 ) );
  NAND3_X1 u1_u12_u6_U93 (.ZN( u1_u12_u6_n142 ) , .A2( u1_u12_u6_n172 ) , .A3( u1_u12_u6_n89 ) , .A1( u1_u12_u6_n90 ) );
  XOR2_X1 u1_u13_U22 (.B( u1_K14_34 ) , .A( u1_R12_23 ) , .Z( u1_u13_X_34 ) );
  XOR2_X1 u1_u13_U23 (.B( u1_K14_33 ) , .A( u1_R12_22 ) , .Z( u1_u13_X_33 ) );
  INV_X1 u1_u13_u5_U10 (.A( u1_u13_u5_n121 ) , .ZN( u1_u13_u5_n177 ) );
  AOI222_X1 u1_u13_u5_U100 (.ZN( u1_u13_u5_n113 ) , .A1( u1_u13_u5_n131 ) , .C1( u1_u13_u5_n148 ) , .B2( u1_u13_u5_n174 ) , .C2( u1_u13_u5_n178 ) , .A2( u1_u13_u5_n179 ) , .B1( u1_u13_u5_n99 ) );
  NAND4_X1 u1_u13_u5_U101 (.ZN( u1_out13_11 ) , .A4( u1_u13_u5_n143 ) , .A3( u1_u13_u5_n144 ) , .A2( u1_u13_u5_n169 ) , .A1( u1_u13_u5_n196 ) );
  AOI22_X1 u1_u13_u5_U102 (.A2( u1_u13_u5_n132 ) , .ZN( u1_u13_u5_n144 ) , .B2( u1_u13_u5_n145 ) , .B1( u1_u13_u5_n184 ) , .A1( u1_u13_u5_n194 ) );
  NOR3_X1 u1_u13_u5_U103 (.A3( u1_u13_u5_n141 ) , .A1( u1_u13_u5_n142 ) , .ZN( u1_u13_u5_n143 ) , .A2( u1_u13_u5_n191 ) );
  NAND3_X1 u1_u13_u5_U104 (.A2( u1_u13_u5_n154 ) , .A3( u1_u13_u5_n158 ) , .A1( u1_u13_u5_n161 ) , .ZN( u1_u13_u5_n99 ) );
  NOR2_X1 u1_u13_u5_U11 (.ZN( u1_u13_u5_n160 ) , .A2( u1_u13_u5_n173 ) , .A1( u1_u13_u5_n177 ) );
  INV_X1 u1_u13_u5_U12 (.A( u1_u13_u5_n150 ) , .ZN( u1_u13_u5_n174 ) );
  AOI21_X1 u1_u13_u5_U13 (.A( u1_u13_u5_n160 ) , .B2( u1_u13_u5_n161 ) , .ZN( u1_u13_u5_n162 ) , .B1( u1_u13_u5_n192 ) );
  INV_X1 u1_u13_u5_U14 (.A( u1_u13_u5_n159 ) , .ZN( u1_u13_u5_n192 ) );
  AOI21_X1 u1_u13_u5_U15 (.A( u1_u13_u5_n156 ) , .B2( u1_u13_u5_n157 ) , .B1( u1_u13_u5_n158 ) , .ZN( u1_u13_u5_n163 ) );
  AOI21_X1 u1_u13_u5_U16 (.B2( u1_u13_u5_n139 ) , .B1( u1_u13_u5_n140 ) , .ZN( u1_u13_u5_n141 ) , .A( u1_u13_u5_n150 ) );
  OAI21_X1 u1_u13_u5_U17 (.A( u1_u13_u5_n133 ) , .B2( u1_u13_u5_n134 ) , .B1( u1_u13_u5_n135 ) , .ZN( u1_u13_u5_n142 ) );
  OAI21_X1 u1_u13_u5_U18 (.ZN( u1_u13_u5_n133 ) , .B2( u1_u13_u5_n147 ) , .A( u1_u13_u5_n173 ) , .B1( u1_u13_u5_n188 ) );
  NAND2_X1 u1_u13_u5_U19 (.A2( u1_u13_u5_n119 ) , .A1( u1_u13_u5_n123 ) , .ZN( u1_u13_u5_n137 ) );
  INV_X1 u1_u13_u5_U20 (.A( u1_u13_u5_n155 ) , .ZN( u1_u13_u5_n194 ) );
  NAND2_X1 u1_u13_u5_U21 (.A1( u1_u13_u5_n121 ) , .ZN( u1_u13_u5_n132 ) , .A2( u1_u13_u5_n172 ) );
  NAND2_X1 u1_u13_u5_U22 (.A2( u1_u13_u5_n122 ) , .ZN( u1_u13_u5_n136 ) , .A1( u1_u13_u5_n154 ) );
  NAND2_X1 u1_u13_u5_U23 (.A2( u1_u13_u5_n119 ) , .A1( u1_u13_u5_n120 ) , .ZN( u1_u13_u5_n159 ) );
  INV_X1 u1_u13_u5_U24 (.A( u1_u13_u5_n156 ) , .ZN( u1_u13_u5_n175 ) );
  INV_X1 u1_u13_u5_U25 (.A( u1_u13_u5_n158 ) , .ZN( u1_u13_u5_n188 ) );
  INV_X1 u1_u13_u5_U26 (.A( u1_u13_u5_n152 ) , .ZN( u1_u13_u5_n179 ) );
  INV_X1 u1_u13_u5_U27 (.A( u1_u13_u5_n140 ) , .ZN( u1_u13_u5_n182 ) );
  INV_X1 u1_u13_u5_U28 (.A( u1_u13_u5_n151 ) , .ZN( u1_u13_u5_n183 ) );
  INV_X1 u1_u13_u5_U29 (.A( u1_u13_u5_n123 ) , .ZN( u1_u13_u5_n185 ) );
  NOR2_X1 u1_u13_u5_U3 (.ZN( u1_u13_u5_n134 ) , .A1( u1_u13_u5_n183 ) , .A2( u1_u13_u5_n190 ) );
  INV_X1 u1_u13_u5_U30 (.A( u1_u13_u5_n161 ) , .ZN( u1_u13_u5_n184 ) );
  INV_X1 u1_u13_u5_U31 (.A( u1_u13_u5_n139 ) , .ZN( u1_u13_u5_n189 ) );
  INV_X1 u1_u13_u5_U32 (.A( u1_u13_u5_n157 ) , .ZN( u1_u13_u5_n190 ) );
  INV_X1 u1_u13_u5_U33 (.A( u1_u13_u5_n120 ) , .ZN( u1_u13_u5_n193 ) );
  NAND2_X1 u1_u13_u5_U34 (.ZN( u1_u13_u5_n111 ) , .A1( u1_u13_u5_n140 ) , .A2( u1_u13_u5_n155 ) );
  INV_X1 u1_u13_u5_U35 (.A( u1_u13_u5_n117 ) , .ZN( u1_u13_u5_n196 ) );
  OAI221_X1 u1_u13_u5_U36 (.A( u1_u13_u5_n116 ) , .ZN( u1_u13_u5_n117 ) , .B2( u1_u13_u5_n119 ) , .C1( u1_u13_u5_n153 ) , .C2( u1_u13_u5_n158 ) , .B1( u1_u13_u5_n172 ) );
  AOI222_X1 u1_u13_u5_U37 (.ZN( u1_u13_u5_n116 ) , .B2( u1_u13_u5_n145 ) , .C1( u1_u13_u5_n148 ) , .A2( u1_u13_u5_n174 ) , .C2( u1_u13_u5_n177 ) , .B1( u1_u13_u5_n187 ) , .A1( u1_u13_u5_n193 ) );
  INV_X1 u1_u13_u5_U38 (.A( u1_u13_u5_n115 ) , .ZN( u1_u13_u5_n187 ) );
  NOR2_X1 u1_u13_u5_U39 (.ZN( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n170 ) , .A2( u1_u13_u5_n180 ) );
  INV_X1 u1_u13_u5_U4 (.A( u1_u13_u5_n138 ) , .ZN( u1_u13_u5_n191 ) );
  AOI22_X1 u1_u13_u5_U40 (.B2( u1_u13_u5_n131 ) , .A2( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n169 ) , .B1( u1_u13_u5_n174 ) , .A1( u1_u13_u5_n185 ) );
  NOR2_X1 u1_u13_u5_U41 (.A1( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n150 ) , .A2( u1_u13_u5_n173 ) );
  AOI21_X1 u1_u13_u5_U42 (.A( u1_u13_u5_n118 ) , .B2( u1_u13_u5_n145 ) , .ZN( u1_u13_u5_n168 ) , .B1( u1_u13_u5_n186 ) );
  INV_X1 u1_u13_u5_U43 (.A( u1_u13_u5_n122 ) , .ZN( u1_u13_u5_n186 ) );
  NOR2_X1 u1_u13_u5_U44 (.A1( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n152 ) , .A2( u1_u13_u5_n176 ) );
  NOR2_X1 u1_u13_u5_U45 (.A1( u1_u13_u5_n115 ) , .ZN( u1_u13_u5_n118 ) , .A2( u1_u13_u5_n153 ) );
  NOR2_X1 u1_u13_u5_U46 (.A2( u1_u13_u5_n145 ) , .ZN( u1_u13_u5_n156 ) , .A1( u1_u13_u5_n174 ) );
  NOR2_X1 u1_u13_u5_U47 (.ZN( u1_u13_u5_n121 ) , .A2( u1_u13_u5_n145 ) , .A1( u1_u13_u5_n176 ) );
  AOI22_X1 u1_u13_u5_U48 (.ZN( u1_u13_u5_n114 ) , .A2( u1_u13_u5_n137 ) , .A1( u1_u13_u5_n145 ) , .B2( u1_u13_u5_n175 ) , .B1( u1_u13_u5_n193 ) );
  OAI211_X1 u1_u13_u5_U49 (.B( u1_u13_u5_n124 ) , .A( u1_u13_u5_n125 ) , .C2( u1_u13_u5_n126 ) , .C1( u1_u13_u5_n127 ) , .ZN( u1_u13_u5_n128 ) );
  OAI21_X1 u1_u13_u5_U5 (.B2( u1_u13_u5_n136 ) , .B1( u1_u13_u5_n137 ) , .ZN( u1_u13_u5_n138 ) , .A( u1_u13_u5_n177 ) );
  NOR3_X1 u1_u13_u5_U50 (.ZN( u1_u13_u5_n127 ) , .A1( u1_u13_u5_n136 ) , .A3( u1_u13_u5_n148 ) , .A2( u1_u13_u5_n182 ) );
  OAI21_X1 u1_u13_u5_U51 (.ZN( u1_u13_u5_n124 ) , .A( u1_u13_u5_n177 ) , .B2( u1_u13_u5_n183 ) , .B1( u1_u13_u5_n189 ) );
  OAI21_X1 u1_u13_u5_U52 (.ZN( u1_u13_u5_n125 ) , .A( u1_u13_u5_n174 ) , .B2( u1_u13_u5_n185 ) , .B1( u1_u13_u5_n190 ) );
  AOI21_X1 u1_u13_u5_U53 (.A( u1_u13_u5_n153 ) , .B2( u1_u13_u5_n154 ) , .B1( u1_u13_u5_n155 ) , .ZN( u1_u13_u5_n164 ) );
  AOI21_X1 u1_u13_u5_U54 (.ZN( u1_u13_u5_n110 ) , .B1( u1_u13_u5_n122 ) , .B2( u1_u13_u5_n139 ) , .A( u1_u13_u5_n153 ) );
  INV_X1 u1_u13_u5_U55 (.A( u1_u13_u5_n153 ) , .ZN( u1_u13_u5_n176 ) );
  INV_X1 u1_u13_u5_U56 (.A( u1_u13_u5_n126 ) , .ZN( u1_u13_u5_n173 ) );
  AND2_X1 u1_u13_u5_U57 (.A2( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n107 ) , .ZN( u1_u13_u5_n147 ) );
  AND2_X1 u1_u13_u5_U58 (.A2( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n108 ) , .ZN( u1_u13_u5_n148 ) );
  NAND2_X1 u1_u13_u5_U59 (.A1( u1_u13_u5_n105 ) , .A2( u1_u13_u5_n106 ) , .ZN( u1_u13_u5_n158 ) );
  INV_X1 u1_u13_u5_U6 (.A( u1_u13_u5_n135 ) , .ZN( u1_u13_u5_n178 ) );
  NAND2_X1 u1_u13_u5_U60 (.A2( u1_u13_u5_n108 ) , .A1( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n139 ) );
  NAND2_X1 u1_u13_u5_U61 (.A1( u1_u13_u5_n106 ) , .A2( u1_u13_u5_n108 ) , .ZN( u1_u13_u5_n119 ) );
  NAND2_X1 u1_u13_u5_U62 (.A2( u1_u13_u5_n103 ) , .A1( u1_u13_u5_n105 ) , .ZN( u1_u13_u5_n140 ) );
  NAND2_X1 u1_u13_u5_U63 (.A2( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n105 ) , .ZN( u1_u13_u5_n155 ) );
  NAND2_X1 u1_u13_u5_U64 (.A2( u1_u13_u5_n106 ) , .A1( u1_u13_u5_n107 ) , .ZN( u1_u13_u5_n122 ) );
  NAND2_X1 u1_u13_u5_U65 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n106 ) , .ZN( u1_u13_u5_n115 ) );
  NAND2_X1 u1_u13_u5_U66 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n103 ) , .ZN( u1_u13_u5_n161 ) );
  NAND2_X1 u1_u13_u5_U67 (.A1( u1_u13_u5_n105 ) , .A2( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n154 ) );
  INV_X1 u1_u13_u5_U68 (.A( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n172 ) );
  NAND2_X1 u1_u13_u5_U69 (.A1( u1_u13_u5_n103 ) , .A2( u1_u13_u5_n108 ) , .ZN( u1_u13_u5_n123 ) );
  OAI22_X1 u1_u13_u5_U7 (.B2( u1_u13_u5_n149 ) , .B1( u1_u13_u5_n150 ) , .A2( u1_u13_u5_n151 ) , .A1( u1_u13_u5_n152 ) , .ZN( u1_u13_u5_n165 ) );
  NAND2_X1 u1_u13_u5_U70 (.A2( u1_u13_u5_n103 ) , .A1( u1_u13_u5_n107 ) , .ZN( u1_u13_u5_n151 ) );
  NAND2_X1 u1_u13_u5_U71 (.A2( u1_u13_u5_n107 ) , .A1( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n120 ) );
  NAND2_X1 u1_u13_u5_U72 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n157 ) );
  AND2_X1 u1_u13_u5_U73 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n104 ) , .ZN( u1_u13_u5_n131 ) );
  INV_X1 u1_u13_u5_U74 (.A( u1_u13_u5_n102 ) , .ZN( u1_u13_u5_n195 ) );
  OAI221_X1 u1_u13_u5_U75 (.A( u1_u13_u5_n101 ) , .ZN( u1_u13_u5_n102 ) , .C2( u1_u13_u5_n115 ) , .C1( u1_u13_u5_n126 ) , .B1( u1_u13_u5_n134 ) , .B2( u1_u13_u5_n160 ) );
  OAI21_X1 u1_u13_u5_U76 (.ZN( u1_u13_u5_n101 ) , .B1( u1_u13_u5_n137 ) , .A( u1_u13_u5_n146 ) , .B2( u1_u13_u5_n147 ) );
  NOR2_X1 u1_u13_u5_U77 (.A2( u1_u13_X_34 ) , .A1( u1_u13_X_35 ) , .ZN( u1_u13_u5_n145 ) );
  NOR2_X1 u1_u13_u5_U78 (.A2( u1_u13_X_34 ) , .ZN( u1_u13_u5_n146 ) , .A1( u1_u13_u5_n171 ) );
  NOR2_X1 u1_u13_u5_U79 (.A2( u1_u13_X_31 ) , .A1( u1_u13_X_32 ) , .ZN( u1_u13_u5_n103 ) );
  NOR3_X1 u1_u13_u5_U8 (.A2( u1_u13_u5_n147 ) , .A1( u1_u13_u5_n148 ) , .ZN( u1_u13_u5_n149 ) , .A3( u1_u13_u5_n194 ) );
  NOR2_X1 u1_u13_u5_U80 (.A2( u1_u13_X_36 ) , .ZN( u1_u13_u5_n105 ) , .A1( u1_u13_u5_n180 ) );
  NOR2_X1 u1_u13_u5_U81 (.A2( u1_u13_X_33 ) , .ZN( u1_u13_u5_n108 ) , .A1( u1_u13_u5_n170 ) );
  NOR2_X1 u1_u13_u5_U82 (.A2( u1_u13_X_33 ) , .A1( u1_u13_X_36 ) , .ZN( u1_u13_u5_n107 ) );
  NOR2_X1 u1_u13_u5_U83 (.A2( u1_u13_X_31 ) , .ZN( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n181 ) );
  NAND2_X1 u1_u13_u5_U84 (.A2( u1_u13_X_34 ) , .A1( u1_u13_X_35 ) , .ZN( u1_u13_u5_n153 ) );
  NAND2_X1 u1_u13_u5_U85 (.A1( u1_u13_X_34 ) , .ZN( u1_u13_u5_n126 ) , .A2( u1_u13_u5_n171 ) );
  AND2_X1 u1_u13_u5_U86 (.A1( u1_u13_X_31 ) , .A2( u1_u13_X_32 ) , .ZN( u1_u13_u5_n106 ) );
  AND2_X1 u1_u13_u5_U87 (.A1( u1_u13_X_31 ) , .ZN( u1_u13_u5_n109 ) , .A2( u1_u13_u5_n181 ) );
  INV_X1 u1_u13_u5_U88 (.A( u1_u13_X_33 ) , .ZN( u1_u13_u5_n180 ) );
  INV_X1 u1_u13_u5_U89 (.A( u1_u13_X_35 ) , .ZN( u1_u13_u5_n171 ) );
  NOR2_X1 u1_u13_u5_U9 (.ZN( u1_u13_u5_n135 ) , .A1( u1_u13_u5_n173 ) , .A2( u1_u13_u5_n176 ) );
  INV_X1 u1_u13_u5_U90 (.A( u1_u13_X_36 ) , .ZN( u1_u13_u5_n170 ) );
  INV_X1 u1_u13_u5_U91 (.A( u1_u13_X_32 ) , .ZN( u1_u13_u5_n181 ) );
  NAND4_X1 u1_u13_u5_U92 (.ZN( u1_out13_29 ) , .A4( u1_u13_u5_n129 ) , .A3( u1_u13_u5_n130 ) , .A2( u1_u13_u5_n168 ) , .A1( u1_u13_u5_n196 ) );
  AOI221_X1 u1_u13_u5_U93 (.A( u1_u13_u5_n128 ) , .ZN( u1_u13_u5_n129 ) , .C2( u1_u13_u5_n132 ) , .B2( u1_u13_u5_n159 ) , .B1( u1_u13_u5_n176 ) , .C1( u1_u13_u5_n184 ) );
  AOI222_X1 u1_u13_u5_U94 (.ZN( u1_u13_u5_n130 ) , .A2( u1_u13_u5_n146 ) , .B1( u1_u13_u5_n147 ) , .C2( u1_u13_u5_n175 ) , .B2( u1_u13_u5_n179 ) , .A1( u1_u13_u5_n188 ) , .C1( u1_u13_u5_n194 ) );
  NAND4_X1 u1_u13_u5_U95 (.ZN( u1_out13_19 ) , .A4( u1_u13_u5_n166 ) , .A3( u1_u13_u5_n167 ) , .A2( u1_u13_u5_n168 ) , .A1( u1_u13_u5_n169 ) );
  AOI22_X1 u1_u13_u5_U96 (.B2( u1_u13_u5_n145 ) , .A2( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n167 ) , .B1( u1_u13_u5_n182 ) , .A1( u1_u13_u5_n189 ) );
  NOR4_X1 u1_u13_u5_U97 (.A4( u1_u13_u5_n162 ) , .A3( u1_u13_u5_n163 ) , .A2( u1_u13_u5_n164 ) , .A1( u1_u13_u5_n165 ) , .ZN( u1_u13_u5_n166 ) );
  NAND4_X1 u1_u13_u5_U98 (.ZN( u1_out13_4 ) , .A4( u1_u13_u5_n112 ) , .A2( u1_u13_u5_n113 ) , .A1( u1_u13_u5_n114 ) , .A3( u1_u13_u5_n195 ) );
  AOI211_X1 u1_u13_u5_U99 (.A( u1_u13_u5_n110 ) , .C1( u1_u13_u5_n111 ) , .ZN( u1_u13_u5_n112 ) , .B( u1_u13_u5_n118 ) , .C2( u1_u13_u5_n177 ) );
  XOR2_X1 u1_u14_U29 (.B( u1_K15_28 ) , .A( u1_R13_19 ) , .Z( u1_u14_X_28 ) );
  XOR2_X1 u1_u14_U30 (.B( u1_K15_27 ) , .A( u1_R13_18 ) , .Z( u1_u14_X_27 ) );
  OAI22_X1 u1_u14_u4_U10 (.B2( u1_u14_u4_n135 ) , .ZN( u1_u14_u4_n137 ) , .B1( u1_u14_u4_n153 ) , .A1( u1_u14_u4_n155 ) , .A2( u1_u14_u4_n171 ) );
  AND3_X1 u1_u14_u4_U11 (.A2( u1_u14_u4_n134 ) , .ZN( u1_u14_u4_n135 ) , .A3( u1_u14_u4_n145 ) , .A1( u1_u14_u4_n157 ) );
  NAND2_X1 u1_u14_u4_U12 (.ZN( u1_u14_u4_n132 ) , .A2( u1_u14_u4_n170 ) , .A1( u1_u14_u4_n173 ) );
  AOI21_X1 u1_u14_u4_U13 (.B2( u1_u14_u4_n160 ) , .B1( u1_u14_u4_n161 ) , .ZN( u1_u14_u4_n162 ) , .A( u1_u14_u4_n170 ) );
  AOI21_X1 u1_u14_u4_U14 (.ZN( u1_u14_u4_n107 ) , .B2( u1_u14_u4_n143 ) , .A( u1_u14_u4_n174 ) , .B1( u1_u14_u4_n184 ) );
  AOI21_X1 u1_u14_u4_U15 (.B2( u1_u14_u4_n158 ) , .B1( u1_u14_u4_n159 ) , .ZN( u1_u14_u4_n163 ) , .A( u1_u14_u4_n174 ) );
  AOI21_X1 u1_u14_u4_U16 (.A( u1_u14_u4_n153 ) , .B2( u1_u14_u4_n154 ) , .B1( u1_u14_u4_n155 ) , .ZN( u1_u14_u4_n165 ) );
  AOI21_X1 u1_u14_u4_U17 (.A( u1_u14_u4_n156 ) , .B2( u1_u14_u4_n157 ) , .ZN( u1_u14_u4_n164 ) , .B1( u1_u14_u4_n184 ) );
  INV_X1 u1_u14_u4_U18 (.A( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n170 ) );
  AND2_X1 u1_u14_u4_U19 (.A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n155 ) , .A1( u1_u14_u4_n160 ) );
  INV_X1 u1_u14_u4_U20 (.A( u1_u14_u4_n156 ) , .ZN( u1_u14_u4_n175 ) );
  NAND2_X1 u1_u14_u4_U21 (.A2( u1_u14_u4_n118 ) , .ZN( u1_u14_u4_n131 ) , .A1( u1_u14_u4_n147 ) );
  NAND2_X1 u1_u14_u4_U22 (.A1( u1_u14_u4_n119 ) , .A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n130 ) );
  NAND2_X1 u1_u14_u4_U23 (.ZN( u1_u14_u4_n117 ) , .A2( u1_u14_u4_n118 ) , .A1( u1_u14_u4_n148 ) );
  NAND2_X1 u1_u14_u4_U24 (.ZN( u1_u14_u4_n129 ) , .A1( u1_u14_u4_n134 ) , .A2( u1_u14_u4_n148 ) );
  AND3_X1 u1_u14_u4_U25 (.A1( u1_u14_u4_n119 ) , .A2( u1_u14_u4_n143 ) , .A3( u1_u14_u4_n154 ) , .ZN( u1_u14_u4_n161 ) );
  AND2_X1 u1_u14_u4_U26 (.A1( u1_u14_u4_n145 ) , .A2( u1_u14_u4_n147 ) , .ZN( u1_u14_u4_n159 ) );
  OR3_X1 u1_u14_u4_U27 (.A3( u1_u14_u4_n114 ) , .A2( u1_u14_u4_n115 ) , .A1( u1_u14_u4_n116 ) , .ZN( u1_u14_u4_n136 ) );
  AOI21_X1 u1_u14_u4_U28 (.A( u1_u14_u4_n113 ) , .ZN( u1_u14_u4_n116 ) , .B2( u1_u14_u4_n173 ) , .B1( u1_u14_u4_n174 ) );
  AOI21_X1 u1_u14_u4_U29 (.ZN( u1_u14_u4_n115 ) , .B2( u1_u14_u4_n145 ) , .B1( u1_u14_u4_n146 ) , .A( u1_u14_u4_n156 ) );
  NOR2_X1 u1_u14_u4_U3 (.ZN( u1_u14_u4_n121 ) , .A1( u1_u14_u4_n181 ) , .A2( u1_u14_u4_n182 ) );
  OAI22_X1 u1_u14_u4_U30 (.ZN( u1_u14_u4_n114 ) , .A2( u1_u14_u4_n121 ) , .B1( u1_u14_u4_n160 ) , .B2( u1_u14_u4_n170 ) , .A1( u1_u14_u4_n171 ) );
  INV_X1 u1_u14_u4_U31 (.A( u1_u14_u4_n158 ) , .ZN( u1_u14_u4_n182 ) );
  INV_X1 u1_u14_u4_U32 (.ZN( u1_u14_u4_n181 ) , .A( u1_u14_u4_n96 ) );
  INV_X1 u1_u14_u4_U33 (.A( u1_u14_u4_n144 ) , .ZN( u1_u14_u4_n179 ) );
  INV_X1 u1_u14_u4_U34 (.A( u1_u14_u4_n157 ) , .ZN( u1_u14_u4_n178 ) );
  NAND2_X1 u1_u14_u4_U35 (.A2( u1_u14_u4_n154 ) , .A1( u1_u14_u4_n96 ) , .ZN( u1_u14_u4_n97 ) );
  INV_X1 u1_u14_u4_U36 (.ZN( u1_u14_u4_n186 ) , .A( u1_u14_u4_n95 ) );
  OAI221_X1 u1_u14_u4_U37 (.C1( u1_u14_u4_n134 ) , .B1( u1_u14_u4_n158 ) , .B2( u1_u14_u4_n171 ) , .C2( u1_u14_u4_n173 ) , .A( u1_u14_u4_n94 ) , .ZN( u1_u14_u4_n95 ) );
  AOI222_X1 u1_u14_u4_U38 (.B2( u1_u14_u4_n132 ) , .A1( u1_u14_u4_n138 ) , .C2( u1_u14_u4_n175 ) , .A2( u1_u14_u4_n179 ) , .C1( u1_u14_u4_n181 ) , .B1( u1_u14_u4_n185 ) , .ZN( u1_u14_u4_n94 ) );
  INV_X1 u1_u14_u4_U39 (.A( u1_u14_u4_n113 ) , .ZN( u1_u14_u4_n185 ) );
  INV_X1 u1_u14_u4_U4 (.A( u1_u14_u4_n117 ) , .ZN( u1_u14_u4_n184 ) );
  INV_X1 u1_u14_u4_U40 (.A( u1_u14_u4_n143 ) , .ZN( u1_u14_u4_n183 ) );
  NOR2_X1 u1_u14_u4_U41 (.ZN( u1_u14_u4_n138 ) , .A1( u1_u14_u4_n168 ) , .A2( u1_u14_u4_n169 ) );
  NOR2_X1 u1_u14_u4_U42 (.A1( u1_u14_u4_n150 ) , .A2( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n153 ) );
  NOR2_X1 u1_u14_u4_U43 (.A2( u1_u14_u4_n128 ) , .A1( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n156 ) );
  AOI22_X1 u1_u14_u4_U44 (.B2( u1_u14_u4_n122 ) , .A1( u1_u14_u4_n123 ) , .ZN( u1_u14_u4_n124 ) , .B1( u1_u14_u4_n128 ) , .A2( u1_u14_u4_n172 ) );
  INV_X1 u1_u14_u4_U45 (.A( u1_u14_u4_n153 ) , .ZN( u1_u14_u4_n172 ) );
  NAND2_X1 u1_u14_u4_U46 (.A2( u1_u14_u4_n120 ) , .ZN( u1_u14_u4_n123 ) , .A1( u1_u14_u4_n161 ) );
  AOI22_X1 u1_u14_u4_U47 (.B2( u1_u14_u4_n132 ) , .A2( u1_u14_u4_n133 ) , .ZN( u1_u14_u4_n140 ) , .A1( u1_u14_u4_n150 ) , .B1( u1_u14_u4_n179 ) );
  NAND2_X1 u1_u14_u4_U48 (.ZN( u1_u14_u4_n133 ) , .A2( u1_u14_u4_n146 ) , .A1( u1_u14_u4_n154 ) );
  NAND2_X1 u1_u14_u4_U49 (.A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n154 ) , .A2( u1_u14_u4_n98 ) );
  NOR4_X1 u1_u14_u4_U5 (.A4( u1_u14_u4_n106 ) , .A3( u1_u14_u4_n107 ) , .A2( u1_u14_u4_n108 ) , .A1( u1_u14_u4_n109 ) , .ZN( u1_u14_u4_n110 ) );
  NAND2_X1 u1_u14_u4_U50 (.A1( u1_u14_u4_n101 ) , .ZN( u1_u14_u4_n158 ) , .A2( u1_u14_u4_n99 ) );
  AOI21_X1 u1_u14_u4_U51 (.ZN( u1_u14_u4_n127 ) , .A( u1_u14_u4_n136 ) , .B2( u1_u14_u4_n150 ) , .B1( u1_u14_u4_n180 ) );
  INV_X1 u1_u14_u4_U52 (.A( u1_u14_u4_n160 ) , .ZN( u1_u14_u4_n180 ) );
  NAND2_X1 u1_u14_u4_U53 (.A2( u1_u14_u4_n104 ) , .A1( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n146 ) );
  NAND2_X1 u1_u14_u4_U54 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n160 ) );
  NAND2_X1 u1_u14_u4_U55 (.ZN( u1_u14_u4_n134 ) , .A1( u1_u14_u4_n98 ) , .A2( u1_u14_u4_n99 ) );
  NAND2_X1 u1_u14_u4_U56 (.A1( u1_u14_u4_n103 ) , .A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n143 ) );
  NAND2_X1 u1_u14_u4_U57 (.A2( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n145 ) , .A1( u1_u14_u4_n98 ) );
  NAND2_X1 u1_u14_u4_U58 (.A1( u1_u14_u4_n100 ) , .A2( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n120 ) );
  NAND2_X1 u1_u14_u4_U59 (.A1( u1_u14_u4_n102 ) , .A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n148 ) );
  AOI21_X1 u1_u14_u4_U6 (.ZN( u1_u14_u4_n106 ) , .B2( u1_u14_u4_n146 ) , .B1( u1_u14_u4_n158 ) , .A( u1_u14_u4_n170 ) );
  NAND2_X1 u1_u14_u4_U60 (.A2( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n157 ) );
  INV_X1 u1_u14_u4_U61 (.A( u1_u14_u4_n150 ) , .ZN( u1_u14_u4_n173 ) );
  INV_X1 u1_u14_u4_U62 (.A( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n171 ) );
  NAND2_X1 u1_u14_u4_U63 (.A1( u1_u14_u4_n100 ) , .ZN( u1_u14_u4_n118 ) , .A2( u1_u14_u4_n99 ) );
  NAND2_X1 u1_u14_u4_U64 (.A2( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n144 ) );
  NAND2_X1 u1_u14_u4_U65 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n105 ) , .ZN( u1_u14_u4_n96 ) );
  INV_X1 u1_u14_u4_U66 (.A( u1_u14_u4_n128 ) , .ZN( u1_u14_u4_n174 ) );
  NAND2_X1 u1_u14_u4_U67 (.A2( u1_u14_u4_n102 ) , .ZN( u1_u14_u4_n119 ) , .A1( u1_u14_u4_n98 ) );
  NAND2_X1 u1_u14_u4_U68 (.A2( u1_u14_u4_n101 ) , .A1( u1_u14_u4_n103 ) , .ZN( u1_u14_u4_n147 ) );
  NAND2_X1 u1_u14_u4_U69 (.A2( u1_u14_u4_n104 ) , .ZN( u1_u14_u4_n113 ) , .A1( u1_u14_u4_n99 ) );
  AOI21_X1 u1_u14_u4_U7 (.ZN( u1_u14_u4_n108 ) , .B2( u1_u14_u4_n134 ) , .B1( u1_u14_u4_n155 ) , .A( u1_u14_u4_n156 ) );
  NOR2_X1 u1_u14_u4_U70 (.A2( u1_u14_X_28 ) , .ZN( u1_u14_u4_n150 ) , .A1( u1_u14_u4_n168 ) );
  NOR2_X1 u1_u14_u4_U71 (.A2( u1_u14_X_29 ) , .ZN( u1_u14_u4_n152 ) , .A1( u1_u14_u4_n169 ) );
  NOR2_X1 u1_u14_u4_U72 (.A2( u1_u14_X_30 ) , .ZN( u1_u14_u4_n105 ) , .A1( u1_u14_u4_n176 ) );
  NOR2_X1 u1_u14_u4_U73 (.A2( u1_u14_X_26 ) , .ZN( u1_u14_u4_n100 ) , .A1( u1_u14_u4_n177 ) );
  NOR2_X1 u1_u14_u4_U74 (.A2( u1_u14_X_28 ) , .A1( u1_u14_X_29 ) , .ZN( u1_u14_u4_n128 ) );
  NOR2_X1 u1_u14_u4_U75 (.A2( u1_u14_X_27 ) , .A1( u1_u14_X_30 ) , .ZN( u1_u14_u4_n102 ) );
  NOR2_X1 u1_u14_u4_U76 (.A2( u1_u14_X_25 ) , .A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n98 ) );
  AND2_X1 u1_u14_u4_U77 (.A2( u1_u14_X_25 ) , .A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n104 ) );
  AND2_X1 u1_u14_u4_U78 (.A1( u1_u14_X_30 ) , .A2( u1_u14_u4_n176 ) , .ZN( u1_u14_u4_n99 ) );
  AND2_X1 u1_u14_u4_U79 (.A1( u1_u14_X_26 ) , .ZN( u1_u14_u4_n101 ) , .A2( u1_u14_u4_n177 ) );
  AOI21_X1 u1_u14_u4_U8 (.ZN( u1_u14_u4_n109 ) , .A( u1_u14_u4_n153 ) , .B1( u1_u14_u4_n159 ) , .B2( u1_u14_u4_n184 ) );
  AND2_X1 u1_u14_u4_U80 (.A1( u1_u14_X_27 ) , .A2( u1_u14_X_30 ) , .ZN( u1_u14_u4_n103 ) );
  INV_X1 u1_u14_u4_U81 (.A( u1_u14_X_28 ) , .ZN( u1_u14_u4_n169 ) );
  INV_X1 u1_u14_u4_U82 (.A( u1_u14_X_29 ) , .ZN( u1_u14_u4_n168 ) );
  INV_X1 u1_u14_u4_U83 (.A( u1_u14_X_25 ) , .ZN( u1_u14_u4_n177 ) );
  INV_X1 u1_u14_u4_U84 (.A( u1_u14_X_27 ) , .ZN( u1_u14_u4_n176 ) );
  NAND4_X1 u1_u14_u4_U85 (.ZN( u1_out14_25 ) , .A4( u1_u14_u4_n139 ) , .A3( u1_u14_u4_n140 ) , .A2( u1_u14_u4_n141 ) , .A1( u1_u14_u4_n142 ) );
  OAI21_X1 u1_u14_u4_U86 (.A( u1_u14_u4_n128 ) , .B2( u1_u14_u4_n129 ) , .B1( u1_u14_u4_n130 ) , .ZN( u1_u14_u4_n142 ) );
  OAI21_X1 u1_u14_u4_U87 (.B2( u1_u14_u4_n131 ) , .ZN( u1_u14_u4_n141 ) , .A( u1_u14_u4_n175 ) , .B1( u1_u14_u4_n183 ) );
  NAND4_X1 u1_u14_u4_U88 (.ZN( u1_out14_14 ) , .A4( u1_u14_u4_n124 ) , .A3( u1_u14_u4_n125 ) , .A2( u1_u14_u4_n126 ) , .A1( u1_u14_u4_n127 ) );
  AOI22_X1 u1_u14_u4_U89 (.B2( u1_u14_u4_n117 ) , .ZN( u1_u14_u4_n126 ) , .A1( u1_u14_u4_n129 ) , .B1( u1_u14_u4_n152 ) , .A2( u1_u14_u4_n175 ) );
  AOI211_X1 u1_u14_u4_U9 (.B( u1_u14_u4_n136 ) , .A( u1_u14_u4_n137 ) , .C2( u1_u14_u4_n138 ) , .ZN( u1_u14_u4_n139 ) , .C1( u1_u14_u4_n182 ) );
  AOI22_X1 u1_u14_u4_U90 (.ZN( u1_u14_u4_n125 ) , .B2( u1_u14_u4_n131 ) , .A2( u1_u14_u4_n132 ) , .B1( u1_u14_u4_n138 ) , .A1( u1_u14_u4_n178 ) );
  NAND4_X1 u1_u14_u4_U91 (.ZN( u1_out14_8 ) , .A4( u1_u14_u4_n110 ) , .A3( u1_u14_u4_n111 ) , .A2( u1_u14_u4_n112 ) , .A1( u1_u14_u4_n186 ) );
  NAND2_X1 u1_u14_u4_U92 (.ZN( u1_u14_u4_n112 ) , .A2( u1_u14_u4_n130 ) , .A1( u1_u14_u4_n150 ) );
  AOI22_X1 u1_u14_u4_U93 (.ZN( u1_u14_u4_n111 ) , .B2( u1_u14_u4_n132 ) , .A1( u1_u14_u4_n152 ) , .B1( u1_u14_u4_n178 ) , .A2( u1_u14_u4_n97 ) );
  AOI22_X1 u1_u14_u4_U94 (.B2( u1_u14_u4_n149 ) , .B1( u1_u14_u4_n150 ) , .A2( u1_u14_u4_n151 ) , .A1( u1_u14_u4_n152 ) , .ZN( u1_u14_u4_n167 ) );
  NOR4_X1 u1_u14_u4_U95 (.A4( u1_u14_u4_n162 ) , .A3( u1_u14_u4_n163 ) , .A2( u1_u14_u4_n164 ) , .A1( u1_u14_u4_n165 ) , .ZN( u1_u14_u4_n166 ) );
  NAND3_X1 u1_u14_u4_U96 (.ZN( u1_out14_3 ) , .A3( u1_u14_u4_n166 ) , .A1( u1_u14_u4_n167 ) , .A2( u1_u14_u4_n186 ) );
  NAND3_X1 u1_u14_u4_U97 (.A3( u1_u14_u4_n146 ) , .A2( u1_u14_u4_n147 ) , .A1( u1_u14_u4_n148 ) , .ZN( u1_u14_u4_n149 ) );
  NAND3_X1 u1_u14_u4_U98 (.A3( u1_u14_u4_n143 ) , .A2( u1_u14_u4_n144 ) , .A1( u1_u14_u4_n145 ) , .ZN( u1_u14_u4_n151 ) );
  NAND3_X1 u1_u14_u4_U99 (.A3( u1_u14_u4_n121 ) , .ZN( u1_u14_u4_n122 ) , .A2( u1_u14_u4_n144 ) , .A1( u1_u14_u4_n154 ) );
  XOR2_X1 u1_u15_U16 (.A( u1_FP_34 ) , .B( u1_K16_3 ) , .Z( u1_u15_X_3 ) );
  XOR2_X1 u1_u15_U6 (.A( u1_FP_35 ) , .B( u1_K16_4 ) , .Z( u1_u15_X_4 ) );
  AND3_X1 u1_u15_u0_U10 (.A2( u1_u15_u0_n112 ) , .ZN( u1_u15_u0_n127 ) , .A3( u1_u15_u0_n130 ) , .A1( u1_u15_u0_n148 ) );
  NAND2_X1 u1_u15_u0_U11 (.ZN( u1_u15_u0_n113 ) , .A1( u1_u15_u0_n139 ) , .A2( u1_u15_u0_n149 ) );
  AND2_X1 u1_u15_u0_U12 (.ZN( u1_u15_u0_n107 ) , .A1( u1_u15_u0_n130 ) , .A2( u1_u15_u0_n140 ) );
  AND2_X1 u1_u15_u0_U13 (.A2( u1_u15_u0_n129 ) , .A1( u1_u15_u0_n130 ) , .ZN( u1_u15_u0_n151 ) );
  AND2_X1 u1_u15_u0_U14 (.A1( u1_u15_u0_n108 ) , .A2( u1_u15_u0_n125 ) , .ZN( u1_u15_u0_n145 ) );
  INV_X1 u1_u15_u0_U15 (.A( u1_u15_u0_n143 ) , .ZN( u1_u15_u0_n173 ) );
  NOR2_X1 u1_u15_u0_U16 (.A2( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n147 ) , .A1( u1_u15_u0_n160 ) );
  AOI21_X1 u1_u15_u0_U17 (.B1( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n132 ) , .A( u1_u15_u0_n165 ) , .B2( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U18 (.A( u1_u15_u0_n142 ) , .ZN( u1_u15_u0_n165 ) );
  OAI221_X1 u1_u15_u0_U19 (.C1( u1_u15_u0_n121 ) , .ZN( u1_u15_u0_n122 ) , .B2( u1_u15_u0_n127 ) , .A( u1_u15_u0_n143 ) , .B1( u1_u15_u0_n144 ) , .C2( u1_u15_u0_n147 ) );
  OAI22_X1 u1_u15_u0_U20 (.B1( u1_u15_u0_n131 ) , .A1( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n147 ) , .A2( u1_u15_u0_n90 ) , .ZN( u1_u15_u0_n91 ) );
  AND3_X1 u1_u15_u0_U21 (.A3( u1_u15_u0_n121 ) , .A2( u1_u15_u0_n125 ) , .A1( u1_u15_u0_n148 ) , .ZN( u1_u15_u0_n90 ) );
  OAI22_X1 u1_u15_u0_U22 (.B1( u1_u15_u0_n125 ) , .ZN( u1_u15_u0_n126 ) , .A1( u1_u15_u0_n138 ) , .A2( u1_u15_u0_n146 ) , .B2( u1_u15_u0_n147 ) );
  NOR2_X1 u1_u15_u0_U23 (.A1( u1_u15_u0_n163 ) , .A2( u1_u15_u0_n164 ) , .ZN( u1_u15_u0_n95 ) );
  INV_X1 u1_u15_u0_U24 (.A( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n161 ) );
  NOR2_X1 u1_u15_u0_U25 (.A1( u1_u15_u0_n120 ) , .ZN( u1_u15_u0_n143 ) , .A2( u1_u15_u0_n167 ) );
  OAI221_X1 u1_u15_u0_U26 (.C1( u1_u15_u0_n112 ) , .ZN( u1_u15_u0_n120 ) , .B1( u1_u15_u0_n138 ) , .B2( u1_u15_u0_n141 ) , .C2( u1_u15_u0_n147 ) , .A( u1_u15_u0_n172 ) );
  AOI211_X1 u1_u15_u0_U27 (.B( u1_u15_u0_n115 ) , .A( u1_u15_u0_n116 ) , .C2( u1_u15_u0_n117 ) , .C1( u1_u15_u0_n118 ) , .ZN( u1_u15_u0_n119 ) );
  AOI22_X1 u1_u15_u0_U28 (.B2( u1_u15_u0_n109 ) , .A2( u1_u15_u0_n110 ) , .ZN( u1_u15_u0_n111 ) , .B1( u1_u15_u0_n118 ) , .A1( u1_u15_u0_n160 ) );
  NAND2_X1 u1_u15_u0_U29 (.A2( u1_u15_u0_n102 ) , .A1( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n149 ) );
  INV_X1 u1_u15_u0_U3 (.A( u1_u15_u0_n113 ) , .ZN( u1_u15_u0_n166 ) );
  INV_X1 u1_u15_u0_U30 (.A( u1_u15_u0_n118 ) , .ZN( u1_u15_u0_n158 ) );
  NAND2_X1 u1_u15_u0_U31 (.A2( u1_u15_u0_n100 ) , .ZN( u1_u15_u0_n131 ) , .A1( u1_u15_u0_n92 ) );
  NAND2_X1 u1_u15_u0_U32 (.ZN( u1_u15_u0_n108 ) , .A1( u1_u15_u0_n92 ) , .A2( u1_u15_u0_n94 ) );
  AOI21_X1 u1_u15_u0_U33 (.ZN( u1_u15_u0_n104 ) , .B1( u1_u15_u0_n107 ) , .B2( u1_u15_u0_n141 ) , .A( u1_u15_u0_n144 ) );
  AOI21_X1 u1_u15_u0_U34 (.B1( u1_u15_u0_n127 ) , .B2( u1_u15_u0_n129 ) , .A( u1_u15_u0_n138 ) , .ZN( u1_u15_u0_n96 ) );
  NAND2_X1 u1_u15_u0_U35 (.A2( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n114 ) , .A1( u1_u15_u0_n92 ) );
  AOI21_X1 u1_u15_u0_U36 (.ZN( u1_u15_u0_n116 ) , .B2( u1_u15_u0_n142 ) , .A( u1_u15_u0_n144 ) , .B1( u1_u15_u0_n166 ) );
  NAND2_X1 u1_u15_u0_U37 (.A2( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n140 ) , .A1( u1_u15_u0_n94 ) );
  NAND2_X1 u1_u15_u0_U38 (.A1( u1_u15_u0_n100 ) , .A2( u1_u15_u0_n103 ) , .ZN( u1_u15_u0_n125 ) );
  NAND2_X1 u1_u15_u0_U39 (.A1( u1_u15_u0_n101 ) , .A2( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n150 ) );
  AOI21_X1 u1_u15_u0_U4 (.B1( u1_u15_u0_n114 ) , .ZN( u1_u15_u0_n115 ) , .B2( u1_u15_u0_n129 ) , .A( u1_u15_u0_n161 ) );
  INV_X1 u1_u15_u0_U40 (.A( u1_u15_u0_n138 ) , .ZN( u1_u15_u0_n160 ) );
  NAND2_X1 u1_u15_u0_U41 (.A2( u1_u15_u0_n100 ) , .A1( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n139 ) );
  NAND2_X1 u1_u15_u0_U42 (.ZN( u1_u15_u0_n112 ) , .A2( u1_u15_u0_n92 ) , .A1( u1_u15_u0_n93 ) );
  NAND2_X1 u1_u15_u0_U43 (.A1( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n130 ) , .A2( u1_u15_u0_n94 ) );
  NAND2_X1 u1_u15_u0_U44 (.A2( u1_u15_u0_n101 ) , .ZN( u1_u15_u0_n121 ) , .A1( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U45 (.ZN( u1_u15_u0_n172 ) , .A( u1_u15_u0_n88 ) );
  OAI222_X1 u1_u15_u0_U46 (.C1( u1_u15_u0_n108 ) , .A1( u1_u15_u0_n125 ) , .B2( u1_u15_u0_n128 ) , .B1( u1_u15_u0_n144 ) , .A2( u1_u15_u0_n158 ) , .C2( u1_u15_u0_n161 ) , .ZN( u1_u15_u0_n88 ) );
  OR3_X1 u1_u15_u0_U47 (.A3( u1_u15_u0_n152 ) , .A2( u1_u15_u0_n153 ) , .A1( u1_u15_u0_n154 ) , .ZN( u1_u15_u0_n155 ) );
  AOI21_X1 u1_u15_u0_U48 (.B2( u1_u15_u0_n150 ) , .B1( u1_u15_u0_n151 ) , .ZN( u1_u15_u0_n152 ) , .A( u1_u15_u0_n158 ) );
  AOI21_X1 u1_u15_u0_U49 (.A( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n145 ) , .B1( u1_u15_u0_n146 ) , .ZN( u1_u15_u0_n154 ) );
  AOI21_X1 u1_u15_u0_U5 (.B2( u1_u15_u0_n131 ) , .ZN( u1_u15_u0_n134 ) , .B1( u1_u15_u0_n151 ) , .A( u1_u15_u0_n158 ) );
  AOI21_X1 u1_u15_u0_U50 (.A( u1_u15_u0_n147 ) , .B2( u1_u15_u0_n148 ) , .B1( u1_u15_u0_n149 ) , .ZN( u1_u15_u0_n153 ) );
  INV_X1 u1_u15_u0_U51 (.ZN( u1_u15_u0_n171 ) , .A( u1_u15_u0_n99 ) );
  OAI211_X1 u1_u15_u0_U52 (.C2( u1_u15_u0_n140 ) , .C1( u1_u15_u0_n161 ) , .A( u1_u15_u0_n169 ) , .B( u1_u15_u0_n98 ) , .ZN( u1_u15_u0_n99 ) );
  AOI211_X1 u1_u15_u0_U53 (.C1( u1_u15_u0_n118 ) , .A( u1_u15_u0_n123 ) , .B( u1_u15_u0_n96 ) , .C2( u1_u15_u0_n97 ) , .ZN( u1_u15_u0_n98 ) );
  INV_X1 u1_u15_u0_U54 (.ZN( u1_u15_u0_n169 ) , .A( u1_u15_u0_n91 ) );
  NOR2_X1 u1_u15_u0_U55 (.A2( u1_u15_X_4 ) , .A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n118 ) );
  NOR2_X1 u1_u15_u0_U56 (.A2( u1_u15_X_1 ) , .ZN( u1_u15_u0_n101 ) , .A1( u1_u15_u0_n163 ) );
  NOR2_X1 u1_u15_u0_U57 (.A2( u1_u15_X_3 ) , .A1( u1_u15_X_6 ) , .ZN( u1_u15_u0_n94 ) );
  NOR2_X1 u1_u15_u0_U58 (.A2( u1_u15_X_6 ) , .ZN( u1_u15_u0_n100 ) , .A1( u1_u15_u0_n162 ) );
  NAND2_X1 u1_u15_u0_U59 (.A2( u1_u15_X_4 ) , .A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n144 ) );
  NOR2_X1 u1_u15_u0_U6 (.A1( u1_u15_u0_n108 ) , .ZN( u1_u15_u0_n123 ) , .A2( u1_u15_u0_n158 ) );
  NOR2_X1 u1_u15_u0_U60 (.A2( u1_u15_X_5 ) , .ZN( u1_u15_u0_n136 ) , .A1( u1_u15_u0_n159 ) );
  NAND2_X1 u1_u15_u0_U61 (.A1( u1_u15_X_5 ) , .ZN( u1_u15_u0_n138 ) , .A2( u1_u15_u0_n159 ) );
  AND2_X1 u1_u15_u0_U62 (.A2( u1_u15_X_3 ) , .A1( u1_u15_X_6 ) , .ZN( u1_u15_u0_n102 ) );
  AND2_X1 u1_u15_u0_U63 (.A1( u1_u15_X_6 ) , .A2( u1_u15_u0_n162 ) , .ZN( u1_u15_u0_n93 ) );
  INV_X1 u1_u15_u0_U64 (.A( u1_u15_X_4 ) , .ZN( u1_u15_u0_n159 ) );
  INV_X1 u1_u15_u0_U65 (.A( u1_u15_X_1 ) , .ZN( u1_u15_u0_n164 ) );
  INV_X1 u1_u15_u0_U66 (.A( u1_u15_X_3 ) , .ZN( u1_u15_u0_n162 ) );
  INV_X1 u1_u15_u0_U67 (.A( u1_u15_u0_n126 ) , .ZN( u1_u15_u0_n168 ) );
  AOI211_X1 u1_u15_u0_U68 (.B( u1_u15_u0_n133 ) , .A( u1_u15_u0_n134 ) , .C2( u1_u15_u0_n135 ) , .C1( u1_u15_u0_n136 ) , .ZN( u1_u15_u0_n137 ) );
  INV_X1 u1_u15_u0_U69 (.ZN( u1_u15_u0_n174 ) , .A( u1_u15_u0_n89 ) );
  OAI21_X1 u1_u15_u0_U7 (.B1( u1_u15_u0_n150 ) , .B2( u1_u15_u0_n158 ) , .A( u1_u15_u0_n172 ) , .ZN( u1_u15_u0_n89 ) );
  AOI211_X1 u1_u15_u0_U70 (.B( u1_u15_u0_n104 ) , .A( u1_u15_u0_n105 ) , .ZN( u1_u15_u0_n106 ) , .C2( u1_u15_u0_n113 ) , .C1( u1_u15_u0_n160 ) );
  OR4_X1 u1_u15_u0_U71 (.ZN( u1_out15_17 ) , .A4( u1_u15_u0_n122 ) , .A2( u1_u15_u0_n123 ) , .A1( u1_u15_u0_n124 ) , .A3( u1_u15_u0_n170 ) );
  AOI21_X1 u1_u15_u0_U72 (.B2( u1_u15_u0_n107 ) , .ZN( u1_u15_u0_n124 ) , .B1( u1_u15_u0_n128 ) , .A( u1_u15_u0_n161 ) );
  INV_X1 u1_u15_u0_U73 (.A( u1_u15_u0_n111 ) , .ZN( u1_u15_u0_n170 ) );
  OR4_X1 u1_u15_u0_U74 (.ZN( u1_out15_31 ) , .A4( u1_u15_u0_n155 ) , .A2( u1_u15_u0_n156 ) , .A1( u1_u15_u0_n157 ) , .A3( u1_u15_u0_n173 ) );
  AOI21_X1 u1_u15_u0_U75 (.A( u1_u15_u0_n138 ) , .B2( u1_u15_u0_n139 ) , .B1( u1_u15_u0_n140 ) , .ZN( u1_u15_u0_n157 ) );
  AOI21_X1 u1_u15_u0_U76 (.B2( u1_u15_u0_n141 ) , .B1( u1_u15_u0_n142 ) , .ZN( u1_u15_u0_n156 ) , .A( u1_u15_u0_n161 ) );
  AOI21_X1 u1_u15_u0_U77 (.B1( u1_u15_u0_n132 ) , .ZN( u1_u15_u0_n133 ) , .A( u1_u15_u0_n144 ) , .B2( u1_u15_u0_n166 ) );
  OAI22_X1 u1_u15_u0_U78 (.ZN( u1_u15_u0_n105 ) , .A2( u1_u15_u0_n132 ) , .B1( u1_u15_u0_n146 ) , .A1( u1_u15_u0_n147 ) , .B2( u1_u15_u0_n161 ) );
  NAND2_X1 u1_u15_u0_U79 (.ZN( u1_u15_u0_n110 ) , .A2( u1_u15_u0_n132 ) , .A1( u1_u15_u0_n145 ) );
  AND2_X1 u1_u15_u0_U8 (.A1( u1_u15_u0_n114 ) , .A2( u1_u15_u0_n121 ) , .ZN( u1_u15_u0_n146 ) );
  INV_X1 u1_u15_u0_U80 (.A( u1_u15_u0_n119 ) , .ZN( u1_u15_u0_n167 ) );
  NAND2_X1 u1_u15_u0_U81 (.ZN( u1_u15_u0_n148 ) , .A1( u1_u15_u0_n93 ) , .A2( u1_u15_u0_n95 ) );
  NAND2_X1 u1_u15_u0_U82 (.A1( u1_u15_u0_n100 ) , .ZN( u1_u15_u0_n129 ) , .A2( u1_u15_u0_n95 ) );
  NAND2_X1 u1_u15_u0_U83 (.A1( u1_u15_u0_n102 ) , .ZN( u1_u15_u0_n128 ) , .A2( u1_u15_u0_n95 ) );
  NOR2_X1 u1_u15_u0_U84 (.A2( u1_u15_X_1 ) , .A1( u1_u15_X_2 ) , .ZN( u1_u15_u0_n92 ) );
  NAND2_X1 u1_u15_u0_U85 (.ZN( u1_u15_u0_n142 ) , .A1( u1_u15_u0_n94 ) , .A2( u1_u15_u0_n95 ) );
  NOR2_X1 u1_u15_u0_U86 (.A2( u1_u15_X_2 ) , .ZN( u1_u15_u0_n103 ) , .A1( u1_u15_u0_n164 ) );
  INV_X1 u1_u15_u0_U87 (.A( u1_u15_X_2 ) , .ZN( u1_u15_u0_n163 ) );
  NAND3_X1 u1_u15_u0_U88 (.ZN( u1_out15_23 ) , .A3( u1_u15_u0_n137 ) , .A1( u1_u15_u0_n168 ) , .A2( u1_u15_u0_n171 ) );
  NAND3_X1 u1_u15_u0_U89 (.A3( u1_u15_u0_n127 ) , .A2( u1_u15_u0_n128 ) , .ZN( u1_u15_u0_n135 ) , .A1( u1_u15_u0_n150 ) );
  AND2_X1 u1_u15_u0_U9 (.A1( u1_u15_u0_n131 ) , .ZN( u1_u15_u0_n141 ) , .A2( u1_u15_u0_n150 ) );
  NAND3_X1 u1_u15_u0_U90 (.ZN( u1_u15_u0_n117 ) , .A3( u1_u15_u0_n132 ) , .A2( u1_u15_u0_n139 ) , .A1( u1_u15_u0_n148 ) );
  NAND3_X1 u1_u15_u0_U91 (.ZN( u1_u15_u0_n109 ) , .A2( u1_u15_u0_n114 ) , .A3( u1_u15_u0_n140 ) , .A1( u1_u15_u0_n149 ) );
  NAND3_X1 u1_u15_u0_U92 (.ZN( u1_out15_9 ) , .A3( u1_u15_u0_n106 ) , .A2( u1_u15_u0_n171 ) , .A1( u1_u15_u0_n174 ) );
  NAND3_X1 u1_u15_u0_U93 (.A2( u1_u15_u0_n128 ) , .A1( u1_u15_u0_n132 ) , .A3( u1_u15_u0_n146 ) , .ZN( u1_u15_u0_n97 ) );
  XOR2_X1 u1_u2_U22 (.B( u1_K3_34 ) , .A( u1_R1_23 ) , .Z( u1_u2_X_34 ) );
  XOR2_X1 u1_u2_U23 (.B( u1_K3_33 ) , .A( u1_R1_22 ) , .Z( u1_u2_X_33 ) );
  XOR2_X1 u1_u2_U42 (.B( u1_K3_16 ) , .A( u1_R1_11 ) , .Z( u1_u2_X_16 ) );
  XOR2_X1 u1_u2_U43 (.B( u1_K3_15 ) , .A( u1_R1_10 ) , .Z( u1_u2_X_15 ) );
  OAI22_X1 u1_u2_u2_U10 (.B1( u1_u2_u2_n151 ) , .A2( u1_u2_u2_n152 ) , .A1( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n160 ) , .B2( u1_u2_u2_n168 ) );
  NAND3_X1 u1_u2_u2_U100 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n104 ) , .A3( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n98 ) );
  NOR3_X1 u1_u2_u2_U11 (.A1( u1_u2_u2_n150 ) , .ZN( u1_u2_u2_n151 ) , .A3( u1_u2_u2_n175 ) , .A2( u1_u2_u2_n188 ) );
  AOI21_X1 u1_u2_u2_U12 (.B2( u1_u2_u2_n123 ) , .ZN( u1_u2_u2_n125 ) , .A( u1_u2_u2_n171 ) , .B1( u1_u2_u2_n184 ) );
  INV_X1 u1_u2_u2_U13 (.A( u1_u2_u2_n150 ) , .ZN( u1_u2_u2_n184 ) );
  AOI21_X1 u1_u2_u2_U14 (.ZN( u1_u2_u2_n144 ) , .B2( u1_u2_u2_n155 ) , .A( u1_u2_u2_n172 ) , .B1( u1_u2_u2_n185 ) );
  AOI21_X1 u1_u2_u2_U15 (.B2( u1_u2_u2_n143 ) , .ZN( u1_u2_u2_n145 ) , .B1( u1_u2_u2_n152 ) , .A( u1_u2_u2_n171 ) );
  INV_X1 u1_u2_u2_U16 (.A( u1_u2_u2_n156 ) , .ZN( u1_u2_u2_n171 ) );
  INV_X1 u1_u2_u2_U17 (.A( u1_u2_u2_n120 ) , .ZN( u1_u2_u2_n188 ) );
  NAND2_X1 u1_u2_u2_U18 (.A2( u1_u2_u2_n122 ) , .ZN( u1_u2_u2_n150 ) , .A1( u1_u2_u2_n152 ) );
  INV_X1 u1_u2_u2_U19 (.A( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n170 ) );
  INV_X1 u1_u2_u2_U20 (.A( u1_u2_u2_n137 ) , .ZN( u1_u2_u2_n173 ) );
  NAND2_X1 u1_u2_u2_U21 (.A1( u1_u2_u2_n132 ) , .A2( u1_u2_u2_n139 ) , .ZN( u1_u2_u2_n157 ) );
  INV_X1 u1_u2_u2_U22 (.A( u1_u2_u2_n113 ) , .ZN( u1_u2_u2_n178 ) );
  INV_X1 u1_u2_u2_U23 (.A( u1_u2_u2_n139 ) , .ZN( u1_u2_u2_n175 ) );
  INV_X1 u1_u2_u2_U24 (.A( u1_u2_u2_n155 ) , .ZN( u1_u2_u2_n181 ) );
  INV_X1 u1_u2_u2_U25 (.A( u1_u2_u2_n119 ) , .ZN( u1_u2_u2_n177 ) );
  INV_X1 u1_u2_u2_U26 (.A( u1_u2_u2_n116 ) , .ZN( u1_u2_u2_n180 ) );
  INV_X1 u1_u2_u2_U27 (.A( u1_u2_u2_n131 ) , .ZN( u1_u2_u2_n179 ) );
  INV_X1 u1_u2_u2_U28 (.A( u1_u2_u2_n154 ) , .ZN( u1_u2_u2_n176 ) );
  NAND2_X1 u1_u2_u2_U29 (.A2( u1_u2_u2_n116 ) , .A1( u1_u2_u2_n117 ) , .ZN( u1_u2_u2_n118 ) );
  NOR2_X1 u1_u2_u2_U3 (.ZN( u1_u2_u2_n121 ) , .A2( u1_u2_u2_n177 ) , .A1( u1_u2_u2_n180 ) );
  INV_X1 u1_u2_u2_U30 (.A( u1_u2_u2_n132 ) , .ZN( u1_u2_u2_n182 ) );
  INV_X1 u1_u2_u2_U31 (.A( u1_u2_u2_n158 ) , .ZN( u1_u2_u2_n183 ) );
  OAI21_X1 u1_u2_u2_U32 (.A( u1_u2_u2_n156 ) , .B1( u1_u2_u2_n157 ) , .ZN( u1_u2_u2_n158 ) , .B2( u1_u2_u2_n179 ) );
  NOR2_X1 u1_u2_u2_U33 (.ZN( u1_u2_u2_n156 ) , .A1( u1_u2_u2_n166 ) , .A2( u1_u2_u2_n169 ) );
  NOR2_X1 u1_u2_u2_U34 (.A2( u1_u2_u2_n114 ) , .ZN( u1_u2_u2_n137 ) , .A1( u1_u2_u2_n140 ) );
  NOR2_X1 u1_u2_u2_U35 (.A2( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n153 ) , .A1( u1_u2_u2_n156 ) );
  AOI211_X1 u1_u2_u2_U36 (.ZN( u1_u2_u2_n130 ) , .C1( u1_u2_u2_n138 ) , .C2( u1_u2_u2_n179 ) , .B( u1_u2_u2_n96 ) , .A( u1_u2_u2_n97 ) );
  OAI22_X1 u1_u2_u2_U37 (.B1( u1_u2_u2_n133 ) , .A2( u1_u2_u2_n137 ) , .A1( u1_u2_u2_n152 ) , .B2( u1_u2_u2_n168 ) , .ZN( u1_u2_u2_n97 ) );
  OAI221_X1 u1_u2_u2_U38 (.B1( u1_u2_u2_n113 ) , .C1( u1_u2_u2_n132 ) , .A( u1_u2_u2_n149 ) , .B2( u1_u2_u2_n171 ) , .C2( u1_u2_u2_n172 ) , .ZN( u1_u2_u2_n96 ) );
  OAI221_X1 u1_u2_u2_U39 (.A( u1_u2_u2_n115 ) , .C2( u1_u2_u2_n123 ) , .B2( u1_u2_u2_n143 ) , .B1( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n163 ) , .C1( u1_u2_u2_n168 ) );
  INV_X1 u1_u2_u2_U4 (.A( u1_u2_u2_n134 ) , .ZN( u1_u2_u2_n185 ) );
  OAI21_X1 u1_u2_u2_U40 (.A( u1_u2_u2_n114 ) , .ZN( u1_u2_u2_n115 ) , .B1( u1_u2_u2_n176 ) , .B2( u1_u2_u2_n178 ) );
  OAI221_X1 u1_u2_u2_U41 (.A( u1_u2_u2_n135 ) , .B2( u1_u2_u2_n136 ) , .B1( u1_u2_u2_n137 ) , .ZN( u1_u2_u2_n162 ) , .C2( u1_u2_u2_n167 ) , .C1( u1_u2_u2_n185 ) );
  AND3_X1 u1_u2_u2_U42 (.A3( u1_u2_u2_n131 ) , .A2( u1_u2_u2_n132 ) , .A1( u1_u2_u2_n133 ) , .ZN( u1_u2_u2_n136 ) );
  AOI22_X1 u1_u2_u2_U43 (.ZN( u1_u2_u2_n135 ) , .B1( u1_u2_u2_n140 ) , .A1( u1_u2_u2_n156 ) , .B2( u1_u2_u2_n180 ) , .A2( u1_u2_u2_n188 ) );
  AOI21_X1 u1_u2_u2_U44 (.ZN( u1_u2_u2_n149 ) , .B1( u1_u2_u2_n173 ) , .B2( u1_u2_u2_n188 ) , .A( u1_u2_u2_n95 ) );
  AND3_X1 u1_u2_u2_U45 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n104 ) , .A3( u1_u2_u2_n156 ) , .ZN( u1_u2_u2_n95 ) );
  OAI21_X1 u1_u2_u2_U46 (.A( u1_u2_u2_n101 ) , .B2( u1_u2_u2_n121 ) , .B1( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n164 ) );
  NAND2_X1 u1_u2_u2_U47 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n107 ) , .ZN( u1_u2_u2_n155 ) );
  NAND2_X1 u1_u2_u2_U48 (.A2( u1_u2_u2_n105 ) , .A1( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n143 ) );
  NAND2_X1 u1_u2_u2_U49 (.A1( u1_u2_u2_n104 ) , .A2( u1_u2_u2_n106 ) , .ZN( u1_u2_u2_n152 ) );
  NOR4_X1 u1_u2_u2_U5 (.A4( u1_u2_u2_n124 ) , .A3( u1_u2_u2_n125 ) , .A2( u1_u2_u2_n126 ) , .A1( u1_u2_u2_n127 ) , .ZN( u1_u2_u2_n128 ) );
  NAND2_X1 u1_u2_u2_U50 (.A1( u1_u2_u2_n100 ) , .A2( u1_u2_u2_n105 ) , .ZN( u1_u2_u2_n132 ) );
  INV_X1 u1_u2_u2_U51 (.A( u1_u2_u2_n140 ) , .ZN( u1_u2_u2_n168 ) );
  INV_X1 u1_u2_u2_U52 (.A( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n167 ) );
  OAI21_X1 u1_u2_u2_U53 (.A( u1_u2_u2_n141 ) , .B2( u1_u2_u2_n142 ) , .ZN( u1_u2_u2_n146 ) , .B1( u1_u2_u2_n153 ) );
  OAI21_X1 u1_u2_u2_U54 (.A( u1_u2_u2_n140 ) , .ZN( u1_u2_u2_n141 ) , .B1( u1_u2_u2_n176 ) , .B2( u1_u2_u2_n177 ) );
  NOR3_X1 u1_u2_u2_U55 (.ZN( u1_u2_u2_n142 ) , .A3( u1_u2_u2_n175 ) , .A2( u1_u2_u2_n178 ) , .A1( u1_u2_u2_n181 ) );
  NAND2_X1 u1_u2_u2_U56 (.A1( u1_u2_u2_n102 ) , .A2( u1_u2_u2_n106 ) , .ZN( u1_u2_u2_n113 ) );
  NAND2_X1 u1_u2_u2_U57 (.A1( u1_u2_u2_n106 ) , .A2( u1_u2_u2_n107 ) , .ZN( u1_u2_u2_n131 ) );
  NAND2_X1 u1_u2_u2_U58 (.A1( u1_u2_u2_n103 ) , .A2( u1_u2_u2_n107 ) , .ZN( u1_u2_u2_n139 ) );
  NAND2_X1 u1_u2_u2_U59 (.A1( u1_u2_u2_n103 ) , .A2( u1_u2_u2_n105 ) , .ZN( u1_u2_u2_n133 ) );
  AOI21_X1 u1_u2_u2_U6 (.B2( u1_u2_u2_n119 ) , .ZN( u1_u2_u2_n127 ) , .A( u1_u2_u2_n137 ) , .B1( u1_u2_u2_n155 ) );
  NAND2_X1 u1_u2_u2_U60 (.A1( u1_u2_u2_n102 ) , .A2( u1_u2_u2_n103 ) , .ZN( u1_u2_u2_n154 ) );
  NAND2_X1 u1_u2_u2_U61 (.A2( u1_u2_u2_n103 ) , .A1( u1_u2_u2_n104 ) , .ZN( u1_u2_u2_n119 ) );
  NAND2_X1 u1_u2_u2_U62 (.A2( u1_u2_u2_n107 ) , .A1( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n123 ) );
  NAND2_X1 u1_u2_u2_U63 (.A1( u1_u2_u2_n104 ) , .A2( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n122 ) );
  INV_X1 u1_u2_u2_U64 (.A( u1_u2_u2_n114 ) , .ZN( u1_u2_u2_n172 ) );
  NAND2_X1 u1_u2_u2_U65 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n102 ) , .ZN( u1_u2_u2_n116 ) );
  NAND2_X1 u1_u2_u2_U66 (.A1( u1_u2_u2_n102 ) , .A2( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n120 ) );
  NAND2_X1 u1_u2_u2_U67 (.A2( u1_u2_u2_n105 ) , .A1( u1_u2_u2_n106 ) , .ZN( u1_u2_u2_n117 ) );
  INV_X1 u1_u2_u2_U68 (.ZN( u1_u2_u2_n187 ) , .A( u1_u2_u2_n99 ) );
  OAI21_X1 u1_u2_u2_U69 (.B1( u1_u2_u2_n137 ) , .B2( u1_u2_u2_n143 ) , .A( u1_u2_u2_n98 ) , .ZN( u1_u2_u2_n99 ) );
  AOI21_X1 u1_u2_u2_U7 (.ZN( u1_u2_u2_n124 ) , .B1( u1_u2_u2_n131 ) , .B2( u1_u2_u2_n143 ) , .A( u1_u2_u2_n172 ) );
  NOR2_X1 u1_u2_u2_U70 (.A2( u1_u2_X_16 ) , .ZN( u1_u2_u2_n140 ) , .A1( u1_u2_u2_n166 ) );
  NOR2_X1 u1_u2_u2_U71 (.A2( u1_u2_X_13 ) , .A1( u1_u2_X_14 ) , .ZN( u1_u2_u2_n100 ) );
  NOR2_X1 u1_u2_u2_U72 (.A2( u1_u2_X_16 ) , .A1( u1_u2_X_17 ) , .ZN( u1_u2_u2_n138 ) );
  NOR2_X1 u1_u2_u2_U73 (.A2( u1_u2_X_15 ) , .A1( u1_u2_X_18 ) , .ZN( u1_u2_u2_n104 ) );
  NOR2_X1 u1_u2_u2_U74 (.A2( u1_u2_X_14 ) , .ZN( u1_u2_u2_n103 ) , .A1( u1_u2_u2_n174 ) );
  NOR2_X1 u1_u2_u2_U75 (.A2( u1_u2_X_15 ) , .ZN( u1_u2_u2_n102 ) , .A1( u1_u2_u2_n165 ) );
  NOR2_X1 u1_u2_u2_U76 (.A2( u1_u2_X_17 ) , .ZN( u1_u2_u2_n114 ) , .A1( u1_u2_u2_n169 ) );
  AND2_X1 u1_u2_u2_U77 (.A1( u1_u2_X_15 ) , .ZN( u1_u2_u2_n105 ) , .A2( u1_u2_u2_n165 ) );
  AND2_X1 u1_u2_u2_U78 (.A2( u1_u2_X_15 ) , .A1( u1_u2_X_18 ) , .ZN( u1_u2_u2_n107 ) );
  AND2_X1 u1_u2_u2_U79 (.A1( u1_u2_X_14 ) , .ZN( u1_u2_u2_n106 ) , .A2( u1_u2_u2_n174 ) );
  AOI21_X1 u1_u2_u2_U8 (.B2( u1_u2_u2_n120 ) , .B1( u1_u2_u2_n121 ) , .ZN( u1_u2_u2_n126 ) , .A( u1_u2_u2_n167 ) );
  AND2_X1 u1_u2_u2_U80 (.A1( u1_u2_X_13 ) , .A2( u1_u2_X_14 ) , .ZN( u1_u2_u2_n108 ) );
  INV_X1 u1_u2_u2_U81 (.A( u1_u2_X_16 ) , .ZN( u1_u2_u2_n169 ) );
  INV_X1 u1_u2_u2_U82 (.A( u1_u2_X_17 ) , .ZN( u1_u2_u2_n166 ) );
  INV_X1 u1_u2_u2_U83 (.A( u1_u2_X_13 ) , .ZN( u1_u2_u2_n174 ) );
  INV_X1 u1_u2_u2_U84 (.A( u1_u2_X_18 ) , .ZN( u1_u2_u2_n165 ) );
  NAND4_X1 u1_u2_u2_U85 (.ZN( u1_out2_24 ) , .A4( u1_u2_u2_n111 ) , .A3( u1_u2_u2_n112 ) , .A1( u1_u2_u2_n130 ) , .A2( u1_u2_u2_n187 ) );
  AOI21_X1 u1_u2_u2_U86 (.ZN( u1_u2_u2_n112 ) , .B2( u1_u2_u2_n156 ) , .A( u1_u2_u2_n164 ) , .B1( u1_u2_u2_n181 ) );
  AOI221_X1 u1_u2_u2_U87 (.A( u1_u2_u2_n109 ) , .B1( u1_u2_u2_n110 ) , .ZN( u1_u2_u2_n111 ) , .C1( u1_u2_u2_n134 ) , .C2( u1_u2_u2_n170 ) , .B2( u1_u2_u2_n173 ) );
  NAND4_X1 u1_u2_u2_U88 (.ZN( u1_out2_16 ) , .A4( u1_u2_u2_n128 ) , .A3( u1_u2_u2_n129 ) , .A1( u1_u2_u2_n130 ) , .A2( u1_u2_u2_n186 ) );
  AOI22_X1 u1_u2_u2_U89 (.A2( u1_u2_u2_n118 ) , .ZN( u1_u2_u2_n129 ) , .A1( u1_u2_u2_n140 ) , .B1( u1_u2_u2_n157 ) , .B2( u1_u2_u2_n170 ) );
  OAI22_X1 u1_u2_u2_U9 (.ZN( u1_u2_u2_n109 ) , .A2( u1_u2_u2_n113 ) , .B2( u1_u2_u2_n133 ) , .B1( u1_u2_u2_n167 ) , .A1( u1_u2_u2_n168 ) );
  INV_X1 u1_u2_u2_U90 (.A( u1_u2_u2_n163 ) , .ZN( u1_u2_u2_n186 ) );
  NAND4_X1 u1_u2_u2_U91 (.ZN( u1_out2_30 ) , .A4( u1_u2_u2_n147 ) , .A3( u1_u2_u2_n148 ) , .A2( u1_u2_u2_n149 ) , .A1( u1_u2_u2_n187 ) );
  NOR3_X1 u1_u2_u2_U92 (.A3( u1_u2_u2_n144 ) , .A2( u1_u2_u2_n145 ) , .A1( u1_u2_u2_n146 ) , .ZN( u1_u2_u2_n147 ) );
  AOI21_X1 u1_u2_u2_U93 (.B2( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n148 ) , .A( u1_u2_u2_n162 ) , .B1( u1_u2_u2_n182 ) );
  OR4_X1 u1_u2_u2_U94 (.ZN( u1_out2_6 ) , .A4( u1_u2_u2_n161 ) , .A3( u1_u2_u2_n162 ) , .A2( u1_u2_u2_n163 ) , .A1( u1_u2_u2_n164 ) );
  OR3_X1 u1_u2_u2_U95 (.A2( u1_u2_u2_n159 ) , .A1( u1_u2_u2_n160 ) , .ZN( u1_u2_u2_n161 ) , .A3( u1_u2_u2_n183 ) );
  AOI21_X1 u1_u2_u2_U96 (.B2( u1_u2_u2_n154 ) , .B1( u1_u2_u2_n155 ) , .ZN( u1_u2_u2_n159 ) , .A( u1_u2_u2_n167 ) );
  NAND3_X1 u1_u2_u2_U97 (.A2( u1_u2_u2_n117 ) , .A1( u1_u2_u2_n122 ) , .A3( u1_u2_u2_n123 ) , .ZN( u1_u2_u2_n134 ) );
  NAND3_X1 u1_u2_u2_U98 (.ZN( u1_u2_u2_n110 ) , .A2( u1_u2_u2_n131 ) , .A3( u1_u2_u2_n139 ) , .A1( u1_u2_u2_n154 ) );
  NAND3_X1 u1_u2_u2_U99 (.A2( u1_u2_u2_n100 ) , .ZN( u1_u2_u2_n101 ) , .A1( u1_u2_u2_n104 ) , .A3( u1_u2_u2_n114 ) );
  INV_X1 u1_u2_u5_U10 (.A( u1_u2_u5_n121 ) , .ZN( u1_u2_u5_n177 ) );
  NOR3_X1 u1_u2_u5_U100 (.A3( u1_u2_u5_n141 ) , .A1( u1_u2_u5_n142 ) , .ZN( u1_u2_u5_n143 ) , .A2( u1_u2_u5_n191 ) );
  NAND4_X1 u1_u2_u5_U101 (.ZN( u1_out2_4 ) , .A4( u1_u2_u5_n112 ) , .A2( u1_u2_u5_n113 ) , .A1( u1_u2_u5_n114 ) , .A3( u1_u2_u5_n195 ) );
  AOI211_X1 u1_u2_u5_U102 (.A( u1_u2_u5_n110 ) , .C1( u1_u2_u5_n111 ) , .ZN( u1_u2_u5_n112 ) , .B( u1_u2_u5_n118 ) , .C2( u1_u2_u5_n177 ) );
  AOI222_X1 u1_u2_u5_U103 (.ZN( u1_u2_u5_n113 ) , .A1( u1_u2_u5_n131 ) , .C1( u1_u2_u5_n148 ) , .B2( u1_u2_u5_n174 ) , .C2( u1_u2_u5_n178 ) , .A2( u1_u2_u5_n179 ) , .B1( u1_u2_u5_n99 ) );
  NAND3_X1 u1_u2_u5_U104 (.A2( u1_u2_u5_n154 ) , .A3( u1_u2_u5_n158 ) , .A1( u1_u2_u5_n161 ) , .ZN( u1_u2_u5_n99 ) );
  NOR2_X1 u1_u2_u5_U11 (.ZN( u1_u2_u5_n160 ) , .A2( u1_u2_u5_n173 ) , .A1( u1_u2_u5_n177 ) );
  INV_X1 u1_u2_u5_U12 (.A( u1_u2_u5_n150 ) , .ZN( u1_u2_u5_n174 ) );
  AOI21_X1 u1_u2_u5_U13 (.A( u1_u2_u5_n160 ) , .B2( u1_u2_u5_n161 ) , .ZN( u1_u2_u5_n162 ) , .B1( u1_u2_u5_n192 ) );
  INV_X1 u1_u2_u5_U14 (.A( u1_u2_u5_n159 ) , .ZN( u1_u2_u5_n192 ) );
  AOI21_X1 u1_u2_u5_U15 (.A( u1_u2_u5_n156 ) , .B2( u1_u2_u5_n157 ) , .B1( u1_u2_u5_n158 ) , .ZN( u1_u2_u5_n163 ) );
  AOI21_X1 u1_u2_u5_U16 (.B2( u1_u2_u5_n139 ) , .B1( u1_u2_u5_n140 ) , .ZN( u1_u2_u5_n141 ) , .A( u1_u2_u5_n150 ) );
  OAI21_X1 u1_u2_u5_U17 (.A( u1_u2_u5_n133 ) , .B2( u1_u2_u5_n134 ) , .B1( u1_u2_u5_n135 ) , .ZN( u1_u2_u5_n142 ) );
  OAI21_X1 u1_u2_u5_U18 (.ZN( u1_u2_u5_n133 ) , .B2( u1_u2_u5_n147 ) , .A( u1_u2_u5_n173 ) , .B1( u1_u2_u5_n188 ) );
  NAND2_X1 u1_u2_u5_U19 (.A2( u1_u2_u5_n119 ) , .A1( u1_u2_u5_n123 ) , .ZN( u1_u2_u5_n137 ) );
  INV_X1 u1_u2_u5_U20 (.A( u1_u2_u5_n155 ) , .ZN( u1_u2_u5_n194 ) );
  NAND2_X1 u1_u2_u5_U21 (.A1( u1_u2_u5_n121 ) , .ZN( u1_u2_u5_n132 ) , .A2( u1_u2_u5_n172 ) );
  NAND2_X1 u1_u2_u5_U22 (.A2( u1_u2_u5_n122 ) , .ZN( u1_u2_u5_n136 ) , .A1( u1_u2_u5_n154 ) );
  NAND2_X1 u1_u2_u5_U23 (.A2( u1_u2_u5_n119 ) , .A1( u1_u2_u5_n120 ) , .ZN( u1_u2_u5_n159 ) );
  INV_X1 u1_u2_u5_U24 (.A( u1_u2_u5_n156 ) , .ZN( u1_u2_u5_n175 ) );
  INV_X1 u1_u2_u5_U25 (.A( u1_u2_u5_n158 ) , .ZN( u1_u2_u5_n188 ) );
  INV_X1 u1_u2_u5_U26 (.A( u1_u2_u5_n152 ) , .ZN( u1_u2_u5_n179 ) );
  INV_X1 u1_u2_u5_U27 (.A( u1_u2_u5_n140 ) , .ZN( u1_u2_u5_n182 ) );
  INV_X1 u1_u2_u5_U28 (.A( u1_u2_u5_n151 ) , .ZN( u1_u2_u5_n183 ) );
  INV_X1 u1_u2_u5_U29 (.A( u1_u2_u5_n123 ) , .ZN( u1_u2_u5_n185 ) );
  NOR2_X1 u1_u2_u5_U3 (.ZN( u1_u2_u5_n134 ) , .A1( u1_u2_u5_n183 ) , .A2( u1_u2_u5_n190 ) );
  INV_X1 u1_u2_u5_U30 (.A( u1_u2_u5_n161 ) , .ZN( u1_u2_u5_n184 ) );
  INV_X1 u1_u2_u5_U31 (.A( u1_u2_u5_n139 ) , .ZN( u1_u2_u5_n189 ) );
  INV_X1 u1_u2_u5_U32 (.A( u1_u2_u5_n157 ) , .ZN( u1_u2_u5_n190 ) );
  INV_X1 u1_u2_u5_U33 (.A( u1_u2_u5_n120 ) , .ZN( u1_u2_u5_n193 ) );
  NAND2_X1 u1_u2_u5_U34 (.ZN( u1_u2_u5_n111 ) , .A1( u1_u2_u5_n140 ) , .A2( u1_u2_u5_n155 ) );
  INV_X1 u1_u2_u5_U35 (.A( u1_u2_u5_n117 ) , .ZN( u1_u2_u5_n196 ) );
  OAI221_X1 u1_u2_u5_U36 (.A( u1_u2_u5_n116 ) , .ZN( u1_u2_u5_n117 ) , .B2( u1_u2_u5_n119 ) , .C1( u1_u2_u5_n153 ) , .C2( u1_u2_u5_n158 ) , .B1( u1_u2_u5_n172 ) );
  AOI222_X1 u1_u2_u5_U37 (.ZN( u1_u2_u5_n116 ) , .B2( u1_u2_u5_n145 ) , .C1( u1_u2_u5_n148 ) , .A2( u1_u2_u5_n174 ) , .C2( u1_u2_u5_n177 ) , .B1( u1_u2_u5_n187 ) , .A1( u1_u2_u5_n193 ) );
  INV_X1 u1_u2_u5_U38 (.A( u1_u2_u5_n115 ) , .ZN( u1_u2_u5_n187 ) );
  NOR2_X1 u1_u2_u5_U39 (.ZN( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n170 ) , .A2( u1_u2_u5_n180 ) );
  INV_X1 u1_u2_u5_U4 (.A( u1_u2_u5_n138 ) , .ZN( u1_u2_u5_n191 ) );
  AOI22_X1 u1_u2_u5_U40 (.B2( u1_u2_u5_n131 ) , .A2( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n169 ) , .B1( u1_u2_u5_n174 ) , .A1( u1_u2_u5_n185 ) );
  NOR2_X1 u1_u2_u5_U41 (.A1( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n150 ) , .A2( u1_u2_u5_n173 ) );
  AOI21_X1 u1_u2_u5_U42 (.A( u1_u2_u5_n118 ) , .B2( u1_u2_u5_n145 ) , .ZN( u1_u2_u5_n168 ) , .B1( u1_u2_u5_n186 ) );
  INV_X1 u1_u2_u5_U43 (.A( u1_u2_u5_n122 ) , .ZN( u1_u2_u5_n186 ) );
  NOR2_X1 u1_u2_u5_U44 (.A1( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n152 ) , .A2( u1_u2_u5_n176 ) );
  NOR2_X1 u1_u2_u5_U45 (.A1( u1_u2_u5_n115 ) , .ZN( u1_u2_u5_n118 ) , .A2( u1_u2_u5_n153 ) );
  NOR2_X1 u1_u2_u5_U46 (.A2( u1_u2_u5_n145 ) , .ZN( u1_u2_u5_n156 ) , .A1( u1_u2_u5_n174 ) );
  NOR2_X1 u1_u2_u5_U47 (.ZN( u1_u2_u5_n121 ) , .A2( u1_u2_u5_n145 ) , .A1( u1_u2_u5_n176 ) );
  AOI22_X1 u1_u2_u5_U48 (.ZN( u1_u2_u5_n114 ) , .A2( u1_u2_u5_n137 ) , .A1( u1_u2_u5_n145 ) , .B2( u1_u2_u5_n175 ) , .B1( u1_u2_u5_n193 ) );
  OAI211_X1 u1_u2_u5_U49 (.B( u1_u2_u5_n124 ) , .A( u1_u2_u5_n125 ) , .C2( u1_u2_u5_n126 ) , .C1( u1_u2_u5_n127 ) , .ZN( u1_u2_u5_n128 ) );
  OAI21_X1 u1_u2_u5_U5 (.B2( u1_u2_u5_n136 ) , .B1( u1_u2_u5_n137 ) , .ZN( u1_u2_u5_n138 ) , .A( u1_u2_u5_n177 ) );
  NOR3_X1 u1_u2_u5_U50 (.ZN( u1_u2_u5_n127 ) , .A1( u1_u2_u5_n136 ) , .A3( u1_u2_u5_n148 ) , .A2( u1_u2_u5_n182 ) );
  OAI21_X1 u1_u2_u5_U51 (.ZN( u1_u2_u5_n124 ) , .A( u1_u2_u5_n177 ) , .B2( u1_u2_u5_n183 ) , .B1( u1_u2_u5_n189 ) );
  OAI21_X1 u1_u2_u5_U52 (.ZN( u1_u2_u5_n125 ) , .A( u1_u2_u5_n174 ) , .B2( u1_u2_u5_n185 ) , .B1( u1_u2_u5_n190 ) );
  AOI21_X1 u1_u2_u5_U53 (.A( u1_u2_u5_n153 ) , .B2( u1_u2_u5_n154 ) , .B1( u1_u2_u5_n155 ) , .ZN( u1_u2_u5_n164 ) );
  AOI21_X1 u1_u2_u5_U54 (.ZN( u1_u2_u5_n110 ) , .B1( u1_u2_u5_n122 ) , .B2( u1_u2_u5_n139 ) , .A( u1_u2_u5_n153 ) );
  INV_X1 u1_u2_u5_U55 (.A( u1_u2_u5_n153 ) , .ZN( u1_u2_u5_n176 ) );
  INV_X1 u1_u2_u5_U56 (.A( u1_u2_u5_n126 ) , .ZN( u1_u2_u5_n173 ) );
  AND2_X1 u1_u2_u5_U57 (.A2( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n107 ) , .ZN( u1_u2_u5_n147 ) );
  AND2_X1 u1_u2_u5_U58 (.A2( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n108 ) , .ZN( u1_u2_u5_n148 ) );
  NAND2_X1 u1_u2_u5_U59 (.A1( u1_u2_u5_n105 ) , .A2( u1_u2_u5_n106 ) , .ZN( u1_u2_u5_n158 ) );
  INV_X1 u1_u2_u5_U6 (.A( u1_u2_u5_n135 ) , .ZN( u1_u2_u5_n178 ) );
  NAND2_X1 u1_u2_u5_U60 (.A2( u1_u2_u5_n108 ) , .A1( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n139 ) );
  NAND2_X1 u1_u2_u5_U61 (.A1( u1_u2_u5_n106 ) , .A2( u1_u2_u5_n108 ) , .ZN( u1_u2_u5_n119 ) );
  NAND2_X1 u1_u2_u5_U62 (.A2( u1_u2_u5_n103 ) , .A1( u1_u2_u5_n105 ) , .ZN( u1_u2_u5_n140 ) );
  NAND2_X1 u1_u2_u5_U63 (.A2( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n105 ) , .ZN( u1_u2_u5_n155 ) );
  NAND2_X1 u1_u2_u5_U64 (.A2( u1_u2_u5_n106 ) , .A1( u1_u2_u5_n107 ) , .ZN( u1_u2_u5_n122 ) );
  NAND2_X1 u1_u2_u5_U65 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n106 ) , .ZN( u1_u2_u5_n115 ) );
  NAND2_X1 u1_u2_u5_U66 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n103 ) , .ZN( u1_u2_u5_n161 ) );
  NAND2_X1 u1_u2_u5_U67 (.A1( u1_u2_u5_n105 ) , .A2( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n154 ) );
  INV_X1 u1_u2_u5_U68 (.A( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n172 ) );
  NAND2_X1 u1_u2_u5_U69 (.A1( u1_u2_u5_n103 ) , .A2( u1_u2_u5_n108 ) , .ZN( u1_u2_u5_n123 ) );
  OAI22_X1 u1_u2_u5_U7 (.B2( u1_u2_u5_n149 ) , .B1( u1_u2_u5_n150 ) , .A2( u1_u2_u5_n151 ) , .A1( u1_u2_u5_n152 ) , .ZN( u1_u2_u5_n165 ) );
  NAND2_X1 u1_u2_u5_U70 (.A2( u1_u2_u5_n103 ) , .A1( u1_u2_u5_n107 ) , .ZN( u1_u2_u5_n151 ) );
  NAND2_X1 u1_u2_u5_U71 (.A2( u1_u2_u5_n107 ) , .A1( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n120 ) );
  NAND2_X1 u1_u2_u5_U72 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n109 ) , .ZN( u1_u2_u5_n157 ) );
  AND2_X1 u1_u2_u5_U73 (.A2( u1_u2_u5_n100 ) , .A1( u1_u2_u5_n104 ) , .ZN( u1_u2_u5_n131 ) );
  INV_X1 u1_u2_u5_U74 (.A( u1_u2_u5_n102 ) , .ZN( u1_u2_u5_n195 ) );
  OAI221_X1 u1_u2_u5_U75 (.A( u1_u2_u5_n101 ) , .ZN( u1_u2_u5_n102 ) , .C2( u1_u2_u5_n115 ) , .C1( u1_u2_u5_n126 ) , .B1( u1_u2_u5_n134 ) , .B2( u1_u2_u5_n160 ) );
  OAI21_X1 u1_u2_u5_U76 (.ZN( u1_u2_u5_n101 ) , .B1( u1_u2_u5_n137 ) , .A( u1_u2_u5_n146 ) , .B2( u1_u2_u5_n147 ) );
  NOR2_X1 u1_u2_u5_U77 (.A2( u1_u2_X_34 ) , .A1( u1_u2_X_35 ) , .ZN( u1_u2_u5_n145 ) );
  NOR2_X1 u1_u2_u5_U78 (.A2( u1_u2_X_34 ) , .ZN( u1_u2_u5_n146 ) , .A1( u1_u2_u5_n171 ) );
  NOR2_X1 u1_u2_u5_U79 (.A2( u1_u2_X_31 ) , .A1( u1_u2_X_32 ) , .ZN( u1_u2_u5_n103 ) );
  NOR3_X1 u1_u2_u5_U8 (.A2( u1_u2_u5_n147 ) , .A1( u1_u2_u5_n148 ) , .ZN( u1_u2_u5_n149 ) , .A3( u1_u2_u5_n194 ) );
  NOR2_X1 u1_u2_u5_U80 (.A2( u1_u2_X_36 ) , .ZN( u1_u2_u5_n105 ) , .A1( u1_u2_u5_n180 ) );
  NOR2_X1 u1_u2_u5_U81 (.A2( u1_u2_X_33 ) , .ZN( u1_u2_u5_n108 ) , .A1( u1_u2_u5_n170 ) );
  NOR2_X1 u1_u2_u5_U82 (.A2( u1_u2_X_33 ) , .A1( u1_u2_X_36 ) , .ZN( u1_u2_u5_n107 ) );
  NOR2_X1 u1_u2_u5_U83 (.A2( u1_u2_X_31 ) , .ZN( u1_u2_u5_n104 ) , .A1( u1_u2_u5_n181 ) );
  NAND2_X1 u1_u2_u5_U84 (.A2( u1_u2_X_34 ) , .A1( u1_u2_X_35 ) , .ZN( u1_u2_u5_n153 ) );
  NAND2_X1 u1_u2_u5_U85 (.A1( u1_u2_X_34 ) , .ZN( u1_u2_u5_n126 ) , .A2( u1_u2_u5_n171 ) );
  AND2_X1 u1_u2_u5_U86 (.A1( u1_u2_X_31 ) , .A2( u1_u2_X_32 ) , .ZN( u1_u2_u5_n106 ) );
  AND2_X1 u1_u2_u5_U87 (.A1( u1_u2_X_31 ) , .ZN( u1_u2_u5_n109 ) , .A2( u1_u2_u5_n181 ) );
  INV_X1 u1_u2_u5_U88 (.A( u1_u2_X_33 ) , .ZN( u1_u2_u5_n180 ) );
  INV_X1 u1_u2_u5_U89 (.A( u1_u2_X_35 ) , .ZN( u1_u2_u5_n171 ) );
  NOR2_X1 u1_u2_u5_U9 (.ZN( u1_u2_u5_n135 ) , .A1( u1_u2_u5_n173 ) , .A2( u1_u2_u5_n176 ) );
  INV_X1 u1_u2_u5_U90 (.A( u1_u2_X_36 ) , .ZN( u1_u2_u5_n170 ) );
  INV_X1 u1_u2_u5_U91 (.A( u1_u2_X_32 ) , .ZN( u1_u2_u5_n181 ) );
  NAND4_X1 u1_u2_u5_U92 (.ZN( u1_out2_29 ) , .A4( u1_u2_u5_n129 ) , .A3( u1_u2_u5_n130 ) , .A2( u1_u2_u5_n168 ) , .A1( u1_u2_u5_n196 ) );
  AOI221_X1 u1_u2_u5_U93 (.A( u1_u2_u5_n128 ) , .ZN( u1_u2_u5_n129 ) , .C2( u1_u2_u5_n132 ) , .B2( u1_u2_u5_n159 ) , .B1( u1_u2_u5_n176 ) , .C1( u1_u2_u5_n184 ) );
  AOI222_X1 u1_u2_u5_U94 (.ZN( u1_u2_u5_n130 ) , .A2( u1_u2_u5_n146 ) , .B1( u1_u2_u5_n147 ) , .C2( u1_u2_u5_n175 ) , .B2( u1_u2_u5_n179 ) , .A1( u1_u2_u5_n188 ) , .C1( u1_u2_u5_n194 ) );
  NAND4_X1 u1_u2_u5_U95 (.ZN( u1_out2_19 ) , .A4( u1_u2_u5_n166 ) , .A3( u1_u2_u5_n167 ) , .A2( u1_u2_u5_n168 ) , .A1( u1_u2_u5_n169 ) );
  AOI22_X1 u1_u2_u5_U96 (.B2( u1_u2_u5_n145 ) , .A2( u1_u2_u5_n146 ) , .ZN( u1_u2_u5_n167 ) , .B1( u1_u2_u5_n182 ) , .A1( u1_u2_u5_n189 ) );
  NOR4_X1 u1_u2_u5_U97 (.A4( u1_u2_u5_n162 ) , .A3( u1_u2_u5_n163 ) , .A2( u1_u2_u5_n164 ) , .A1( u1_u2_u5_n165 ) , .ZN( u1_u2_u5_n166 ) );
  NAND4_X1 u1_u2_u5_U98 (.ZN( u1_out2_11 ) , .A4( u1_u2_u5_n143 ) , .A3( u1_u2_u5_n144 ) , .A2( u1_u2_u5_n169 ) , .A1( u1_u2_u5_n196 ) );
  AOI22_X1 u1_u2_u5_U99 (.A2( u1_u2_u5_n132 ) , .ZN( u1_u2_u5_n144 ) , .B2( u1_u2_u5_n145 ) , .B1( u1_u2_u5_n184 ) , .A1( u1_u2_u5_n194 ) );
  XOR2_X1 u1_u3_U16 (.B( u1_K4_3 ) , .A( u1_R2_2 ) , .Z( u1_u3_X_3 ) );
  XOR2_X1 u1_u3_U6 (.B( u1_K4_4 ) , .A( u1_R2_3 ) , .Z( u1_u3_X_4 ) );
  AND2_X1 u1_u3_u0_U10 (.A1( u1_u3_u0_n131 ) , .ZN( u1_u3_u0_n141 ) , .A2( u1_u3_u0_n150 ) );
  AND3_X1 u1_u3_u0_U11 (.A2( u1_u3_u0_n112 ) , .ZN( u1_u3_u0_n127 ) , .A3( u1_u3_u0_n130 ) , .A1( u1_u3_u0_n148 ) );
  AND2_X1 u1_u3_u0_U12 (.ZN( u1_u3_u0_n107 ) , .A1( u1_u3_u0_n130 ) , .A2( u1_u3_u0_n140 ) );
  AND2_X1 u1_u3_u0_U13 (.A2( u1_u3_u0_n129 ) , .A1( u1_u3_u0_n130 ) , .ZN( u1_u3_u0_n151 ) );
  AND2_X1 u1_u3_u0_U14 (.A1( u1_u3_u0_n108 ) , .A2( u1_u3_u0_n125 ) , .ZN( u1_u3_u0_n145 ) );
  INV_X1 u1_u3_u0_U15 (.A( u1_u3_u0_n143 ) , .ZN( u1_u3_u0_n173 ) );
  NOR2_X1 u1_u3_u0_U16 (.A2( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n147 ) , .A1( u1_u3_u0_n160 ) );
  AOI21_X1 u1_u3_u0_U17 (.B1( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n132 ) , .A( u1_u3_u0_n165 ) , .B2( u1_u3_u0_n93 ) );
  OAI22_X1 u1_u3_u0_U18 (.B1( u1_u3_u0_n131 ) , .A1( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n147 ) , .A2( u1_u3_u0_n90 ) , .ZN( u1_u3_u0_n91 ) );
  AND3_X1 u1_u3_u0_U19 (.A3( u1_u3_u0_n121 ) , .A2( u1_u3_u0_n125 ) , .A1( u1_u3_u0_n148 ) , .ZN( u1_u3_u0_n90 ) );
  OAI22_X1 u1_u3_u0_U20 (.B1( u1_u3_u0_n125 ) , .ZN( u1_u3_u0_n126 ) , .A1( u1_u3_u0_n138 ) , .A2( u1_u3_u0_n146 ) , .B2( u1_u3_u0_n147 ) );
  NOR2_X1 u1_u3_u0_U21 (.A1( u1_u3_u0_n163 ) , .A2( u1_u3_u0_n164 ) , .ZN( u1_u3_u0_n95 ) );
  AOI22_X1 u1_u3_u0_U22 (.B2( u1_u3_u0_n109 ) , .A2( u1_u3_u0_n110 ) , .ZN( u1_u3_u0_n111 ) , .B1( u1_u3_u0_n118 ) , .A1( u1_u3_u0_n160 ) );
  NAND2_X1 u1_u3_u0_U23 (.A2( u1_u3_u0_n102 ) , .A1( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n149 ) );
  INV_X1 u1_u3_u0_U24 (.A( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n161 ) );
  INV_X1 u1_u3_u0_U25 (.A( u1_u3_u0_n118 ) , .ZN( u1_u3_u0_n158 ) );
  NAND2_X1 u1_u3_u0_U26 (.A2( u1_u3_u0_n100 ) , .ZN( u1_u3_u0_n131 ) , .A1( u1_u3_u0_n92 ) );
  NAND2_X1 u1_u3_u0_U27 (.ZN( u1_u3_u0_n108 ) , .A1( u1_u3_u0_n92 ) , .A2( u1_u3_u0_n94 ) );
  AOI21_X1 u1_u3_u0_U28 (.ZN( u1_u3_u0_n104 ) , .B1( u1_u3_u0_n107 ) , .B2( u1_u3_u0_n141 ) , .A( u1_u3_u0_n144 ) );
  AOI21_X1 u1_u3_u0_U29 (.B1( u1_u3_u0_n127 ) , .B2( u1_u3_u0_n129 ) , .A( u1_u3_u0_n138 ) , .ZN( u1_u3_u0_n96 ) );
  INV_X1 u1_u3_u0_U3 (.A( u1_u3_u0_n113 ) , .ZN( u1_u3_u0_n166 ) );
  NAND2_X1 u1_u3_u0_U30 (.A2( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n114 ) , .A1( u1_u3_u0_n92 ) );
  NOR2_X1 u1_u3_u0_U31 (.A1( u1_u3_u0_n120 ) , .ZN( u1_u3_u0_n143 ) , .A2( u1_u3_u0_n167 ) );
  OAI221_X1 u1_u3_u0_U32 (.C1( u1_u3_u0_n112 ) , .ZN( u1_u3_u0_n120 ) , .B1( u1_u3_u0_n138 ) , .B2( u1_u3_u0_n141 ) , .C2( u1_u3_u0_n147 ) , .A( u1_u3_u0_n172 ) );
  AOI211_X1 u1_u3_u0_U33 (.B( u1_u3_u0_n115 ) , .A( u1_u3_u0_n116 ) , .C2( u1_u3_u0_n117 ) , .C1( u1_u3_u0_n118 ) , .ZN( u1_u3_u0_n119 ) );
  NAND2_X1 u1_u3_u0_U34 (.A2( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n140 ) , .A1( u1_u3_u0_n94 ) );
  NAND2_X1 u1_u3_u0_U35 (.A1( u1_u3_u0_n100 ) , .A2( u1_u3_u0_n103 ) , .ZN( u1_u3_u0_n125 ) );
  NAND2_X1 u1_u3_u0_U36 (.A1( u1_u3_u0_n101 ) , .A2( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n150 ) );
  INV_X1 u1_u3_u0_U37 (.A( u1_u3_u0_n138 ) , .ZN( u1_u3_u0_n160 ) );
  NAND2_X1 u1_u3_u0_U38 (.A2( u1_u3_u0_n100 ) , .A1( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n139 ) );
  NAND2_X1 u1_u3_u0_U39 (.ZN( u1_u3_u0_n112 ) , .A2( u1_u3_u0_n92 ) , .A1( u1_u3_u0_n93 ) );
  AOI21_X1 u1_u3_u0_U4 (.B1( u1_u3_u0_n114 ) , .ZN( u1_u3_u0_n115 ) , .B2( u1_u3_u0_n129 ) , .A( u1_u3_u0_n161 ) );
  NAND2_X1 u1_u3_u0_U40 (.A1( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n130 ) , .A2( u1_u3_u0_n94 ) );
  INV_X1 u1_u3_u0_U41 (.ZN( u1_u3_u0_n172 ) , .A( u1_u3_u0_n88 ) );
  OAI222_X1 u1_u3_u0_U42 (.C1( u1_u3_u0_n108 ) , .A1( u1_u3_u0_n125 ) , .B2( u1_u3_u0_n128 ) , .B1( u1_u3_u0_n144 ) , .A2( u1_u3_u0_n158 ) , .C2( u1_u3_u0_n161 ) , .ZN( u1_u3_u0_n88 ) );
  NAND2_X1 u1_u3_u0_U43 (.A2( u1_u3_u0_n101 ) , .ZN( u1_u3_u0_n121 ) , .A1( u1_u3_u0_n93 ) );
  OR3_X1 u1_u3_u0_U44 (.A3( u1_u3_u0_n152 ) , .A2( u1_u3_u0_n153 ) , .A1( u1_u3_u0_n154 ) , .ZN( u1_u3_u0_n155 ) );
  AOI21_X1 u1_u3_u0_U45 (.A( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n145 ) , .B1( u1_u3_u0_n146 ) , .ZN( u1_u3_u0_n154 ) );
  AOI21_X1 u1_u3_u0_U46 (.B2( u1_u3_u0_n150 ) , .B1( u1_u3_u0_n151 ) , .ZN( u1_u3_u0_n152 ) , .A( u1_u3_u0_n158 ) );
  AOI21_X1 u1_u3_u0_U47 (.A( u1_u3_u0_n147 ) , .B2( u1_u3_u0_n148 ) , .B1( u1_u3_u0_n149 ) , .ZN( u1_u3_u0_n153 ) );
  INV_X1 u1_u3_u0_U48 (.ZN( u1_u3_u0_n171 ) , .A( u1_u3_u0_n99 ) );
  OAI211_X1 u1_u3_u0_U49 (.C2( u1_u3_u0_n140 ) , .C1( u1_u3_u0_n161 ) , .A( u1_u3_u0_n169 ) , .B( u1_u3_u0_n98 ) , .ZN( u1_u3_u0_n99 ) );
  AOI21_X1 u1_u3_u0_U5 (.B2( u1_u3_u0_n131 ) , .ZN( u1_u3_u0_n134 ) , .B1( u1_u3_u0_n151 ) , .A( u1_u3_u0_n158 ) );
  AOI211_X1 u1_u3_u0_U50 (.C1( u1_u3_u0_n118 ) , .A( u1_u3_u0_n123 ) , .B( u1_u3_u0_n96 ) , .C2( u1_u3_u0_n97 ) , .ZN( u1_u3_u0_n98 ) );
  INV_X1 u1_u3_u0_U51 (.ZN( u1_u3_u0_n169 ) , .A( u1_u3_u0_n91 ) );
  NOR2_X1 u1_u3_u0_U52 (.A2( u1_u3_X_4 ) , .A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n118 ) );
  NOR2_X1 u1_u3_u0_U53 (.A2( u1_u3_X_1 ) , .ZN( u1_u3_u0_n101 ) , .A1( u1_u3_u0_n163 ) );
  NOR2_X1 u1_u3_u0_U54 (.A2( u1_u3_X_3 ) , .A1( u1_u3_X_6 ) , .ZN( u1_u3_u0_n94 ) );
  NOR2_X1 u1_u3_u0_U55 (.A2( u1_u3_X_6 ) , .ZN( u1_u3_u0_n100 ) , .A1( u1_u3_u0_n162 ) );
  NAND2_X1 u1_u3_u0_U56 (.A2( u1_u3_X_4 ) , .A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n144 ) );
  NOR2_X1 u1_u3_u0_U57 (.A2( u1_u3_X_5 ) , .ZN( u1_u3_u0_n136 ) , .A1( u1_u3_u0_n159 ) );
  NAND2_X1 u1_u3_u0_U58 (.A1( u1_u3_X_5 ) , .ZN( u1_u3_u0_n138 ) , .A2( u1_u3_u0_n159 ) );
  AND2_X1 u1_u3_u0_U59 (.A2( u1_u3_X_3 ) , .A1( u1_u3_X_6 ) , .ZN( u1_u3_u0_n102 ) );
  NOR2_X1 u1_u3_u0_U6 (.A1( u1_u3_u0_n108 ) , .ZN( u1_u3_u0_n123 ) , .A2( u1_u3_u0_n158 ) );
  AND2_X1 u1_u3_u0_U60 (.A1( u1_u3_X_6 ) , .A2( u1_u3_u0_n162 ) , .ZN( u1_u3_u0_n93 ) );
  INV_X1 u1_u3_u0_U61 (.A( u1_u3_X_4 ) , .ZN( u1_u3_u0_n159 ) );
  INV_X1 u1_u3_u0_U62 (.A( u1_u3_X_1 ) , .ZN( u1_u3_u0_n164 ) );
  INV_X1 u1_u3_u0_U63 (.A( u1_u3_X_3 ) , .ZN( u1_u3_u0_n162 ) );
  INV_X1 u1_u3_u0_U64 (.A( u1_u3_u0_n126 ) , .ZN( u1_u3_u0_n168 ) );
  AOI211_X1 u1_u3_u0_U65 (.B( u1_u3_u0_n133 ) , .A( u1_u3_u0_n134 ) , .C2( u1_u3_u0_n135 ) , .C1( u1_u3_u0_n136 ) , .ZN( u1_u3_u0_n137 ) );
  OR4_X1 u1_u3_u0_U66 (.ZN( u1_out3_17 ) , .A4( u1_u3_u0_n122 ) , .A2( u1_u3_u0_n123 ) , .A1( u1_u3_u0_n124 ) , .A3( u1_u3_u0_n170 ) );
  AOI21_X1 u1_u3_u0_U67 (.B2( u1_u3_u0_n107 ) , .ZN( u1_u3_u0_n124 ) , .B1( u1_u3_u0_n128 ) , .A( u1_u3_u0_n161 ) );
  INV_X1 u1_u3_u0_U68 (.A( u1_u3_u0_n111 ) , .ZN( u1_u3_u0_n170 ) );
  OR4_X1 u1_u3_u0_U69 (.ZN( u1_out3_31 ) , .A4( u1_u3_u0_n155 ) , .A2( u1_u3_u0_n156 ) , .A1( u1_u3_u0_n157 ) , .A3( u1_u3_u0_n173 ) );
  OAI21_X1 u1_u3_u0_U7 (.B1( u1_u3_u0_n150 ) , .B2( u1_u3_u0_n158 ) , .A( u1_u3_u0_n172 ) , .ZN( u1_u3_u0_n89 ) );
  AOI21_X1 u1_u3_u0_U70 (.A( u1_u3_u0_n138 ) , .B2( u1_u3_u0_n139 ) , .B1( u1_u3_u0_n140 ) , .ZN( u1_u3_u0_n157 ) );
  INV_X1 u1_u3_u0_U71 (.ZN( u1_u3_u0_n174 ) , .A( u1_u3_u0_n89 ) );
  AOI211_X1 u1_u3_u0_U72 (.B( u1_u3_u0_n104 ) , .A( u1_u3_u0_n105 ) , .ZN( u1_u3_u0_n106 ) , .C2( u1_u3_u0_n113 ) , .C1( u1_u3_u0_n160 ) );
  AOI21_X1 u1_u3_u0_U73 (.B2( u1_u3_u0_n141 ) , .B1( u1_u3_u0_n142 ) , .ZN( u1_u3_u0_n156 ) , .A( u1_u3_u0_n161 ) );
  AOI21_X1 u1_u3_u0_U74 (.ZN( u1_u3_u0_n116 ) , .B2( u1_u3_u0_n142 ) , .A( u1_u3_u0_n144 ) , .B1( u1_u3_u0_n166 ) );
  INV_X1 u1_u3_u0_U75 (.A( u1_u3_u0_n142 ) , .ZN( u1_u3_u0_n165 ) );
  NOR2_X1 u1_u3_u0_U76 (.A2( u1_u3_X_1 ) , .A1( u1_u3_X_2 ) , .ZN( u1_u3_u0_n92 ) );
  NOR2_X1 u1_u3_u0_U77 (.A2( u1_u3_X_2 ) , .ZN( u1_u3_u0_n103 ) , .A1( u1_u3_u0_n164 ) );
  INV_X1 u1_u3_u0_U78 (.A( u1_u3_X_2 ) , .ZN( u1_u3_u0_n163 ) );
  OAI221_X1 u1_u3_u0_U79 (.C1( u1_u3_u0_n121 ) , .ZN( u1_u3_u0_n122 ) , .B2( u1_u3_u0_n127 ) , .A( u1_u3_u0_n143 ) , .B1( u1_u3_u0_n144 ) , .C2( u1_u3_u0_n147 ) );
  AND2_X1 u1_u3_u0_U8 (.A1( u1_u3_u0_n114 ) , .A2( u1_u3_u0_n121 ) , .ZN( u1_u3_u0_n146 ) );
  AOI21_X1 u1_u3_u0_U80 (.B1( u1_u3_u0_n132 ) , .ZN( u1_u3_u0_n133 ) , .A( u1_u3_u0_n144 ) , .B2( u1_u3_u0_n166 ) );
  OAI22_X1 u1_u3_u0_U81 (.ZN( u1_u3_u0_n105 ) , .A2( u1_u3_u0_n132 ) , .B1( u1_u3_u0_n146 ) , .A1( u1_u3_u0_n147 ) , .B2( u1_u3_u0_n161 ) );
  NAND2_X1 u1_u3_u0_U82 (.ZN( u1_u3_u0_n110 ) , .A2( u1_u3_u0_n132 ) , .A1( u1_u3_u0_n145 ) );
  INV_X1 u1_u3_u0_U83 (.A( u1_u3_u0_n119 ) , .ZN( u1_u3_u0_n167 ) );
  NAND2_X1 u1_u3_u0_U84 (.ZN( u1_u3_u0_n148 ) , .A1( u1_u3_u0_n93 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U85 (.A1( u1_u3_u0_n100 ) , .ZN( u1_u3_u0_n129 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U86 (.A1( u1_u3_u0_n102 ) , .ZN( u1_u3_u0_n128 ) , .A2( u1_u3_u0_n95 ) );
  NAND2_X1 u1_u3_u0_U87 (.ZN( u1_u3_u0_n142 ) , .A1( u1_u3_u0_n94 ) , .A2( u1_u3_u0_n95 ) );
  NAND3_X1 u1_u3_u0_U88 (.ZN( u1_out3_23 ) , .A3( u1_u3_u0_n137 ) , .A1( u1_u3_u0_n168 ) , .A2( u1_u3_u0_n171 ) );
  NAND3_X1 u1_u3_u0_U89 (.A3( u1_u3_u0_n127 ) , .A2( u1_u3_u0_n128 ) , .ZN( u1_u3_u0_n135 ) , .A1( u1_u3_u0_n150 ) );
  NAND2_X1 u1_u3_u0_U9 (.ZN( u1_u3_u0_n113 ) , .A1( u1_u3_u0_n139 ) , .A2( u1_u3_u0_n149 ) );
  NAND3_X1 u1_u3_u0_U90 (.ZN( u1_u3_u0_n117 ) , .A3( u1_u3_u0_n132 ) , .A2( u1_u3_u0_n139 ) , .A1( u1_u3_u0_n148 ) );
  NAND3_X1 u1_u3_u0_U91 (.ZN( u1_u3_u0_n109 ) , .A2( u1_u3_u0_n114 ) , .A3( u1_u3_u0_n140 ) , .A1( u1_u3_u0_n149 ) );
  NAND3_X1 u1_u3_u0_U92 (.ZN( u1_out3_9 ) , .A3( u1_u3_u0_n106 ) , .A2( u1_u3_u0_n171 ) , .A1( u1_u3_u0_n174 ) );
  NAND3_X1 u1_u3_u0_U93 (.A2( u1_u3_u0_n128 ) , .A1( u1_u3_u0_n132 ) , .A3( u1_u3_u0_n146 ) , .ZN( u1_u3_u0_n97 ) );
  XOR2_X1 u1_u4_U1 (.B( u1_K5_9 ) , .A( u1_R3_6 ) , .Z( u1_u4_X_9 ) );
  XOR2_X1 u1_u4_U16 (.B( u1_K5_3 ) , .A( u1_R3_2 ) , .Z( u1_u4_X_3 ) );
  XOR2_X1 u1_u4_U3 (.B( u1_K5_7 ) , .A( u1_R3_4 ) , .Z( u1_u4_X_7 ) );
  XOR2_X1 u1_u4_U35 (.B( u1_K5_22 ) , .A( u1_R3_15 ) , .Z( u1_u4_X_22 ) );
  XOR2_X1 u1_u4_U36 (.B( u1_K5_21 ) , .A( u1_R3_14 ) , .Z( u1_u4_X_21 ) );
  XOR2_X1 u1_u4_U48 (.B( u1_K5_10 ) , .A( u1_R3_7 ) , .Z( u1_u4_X_10 ) );
  XOR2_X1 u1_u4_U5 (.B( u1_K5_5 ) , .A( u1_R3_4 ) , .Z( u1_u4_X_5 ) );
  XOR2_X1 u1_u4_U6 (.B( u1_K5_4 ) , .A( u1_R3_3 ) , .Z( u1_u4_X_4 ) );
  AND3_X1 u1_u4_u0_U10 (.A2( u1_u4_u0_n112 ) , .ZN( u1_u4_u0_n127 ) , .A3( u1_u4_u0_n130 ) , .A1( u1_u4_u0_n148 ) );
  NAND2_X1 u1_u4_u0_U11 (.ZN( u1_u4_u0_n113 ) , .A1( u1_u4_u0_n139 ) , .A2( u1_u4_u0_n149 ) );
  AND2_X1 u1_u4_u0_U12 (.ZN( u1_u4_u0_n107 ) , .A1( u1_u4_u0_n130 ) , .A2( u1_u4_u0_n140 ) );
  AND2_X1 u1_u4_u0_U13 (.A2( u1_u4_u0_n129 ) , .A1( u1_u4_u0_n130 ) , .ZN( u1_u4_u0_n151 ) );
  AND2_X1 u1_u4_u0_U14 (.A1( u1_u4_u0_n108 ) , .A2( u1_u4_u0_n125 ) , .ZN( u1_u4_u0_n145 ) );
  INV_X1 u1_u4_u0_U15 (.A( u1_u4_u0_n143 ) , .ZN( u1_u4_u0_n173 ) );
  NOR2_X1 u1_u4_u0_U16 (.A2( u1_u4_u0_n136 ) , .ZN( u1_u4_u0_n147 ) , .A1( u1_u4_u0_n160 ) );
  NOR2_X1 u1_u4_u0_U17 (.A1( u1_u4_u0_n163 ) , .A2( u1_u4_u0_n164 ) , .ZN( u1_u4_u0_n95 ) );
  AOI21_X1 u1_u4_u0_U18 (.B1( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n132 ) , .A( u1_u4_u0_n165 ) , .B2( u1_u4_u0_n93 ) );
  INV_X1 u1_u4_u0_U19 (.A( u1_u4_u0_n142 ) , .ZN( u1_u4_u0_n165 ) );
  OAI221_X1 u1_u4_u0_U20 (.C1( u1_u4_u0_n112 ) , .ZN( u1_u4_u0_n120 ) , .B1( u1_u4_u0_n138 ) , .B2( u1_u4_u0_n141 ) , .C2( u1_u4_u0_n147 ) , .A( u1_u4_u0_n172 ) );
  AOI211_X1 u1_u4_u0_U21 (.B( u1_u4_u0_n115 ) , .A( u1_u4_u0_n116 ) , .C2( u1_u4_u0_n117 ) , .C1( u1_u4_u0_n118 ) , .ZN( u1_u4_u0_n119 ) );
  OAI22_X1 u1_u4_u0_U22 (.B1( u1_u4_u0_n125 ) , .ZN( u1_u4_u0_n126 ) , .A1( u1_u4_u0_n138 ) , .A2( u1_u4_u0_n146 ) , .B2( u1_u4_u0_n147 ) );
  OAI22_X1 u1_u4_u0_U23 (.B1( u1_u4_u0_n131 ) , .A1( u1_u4_u0_n144 ) , .B2( u1_u4_u0_n147 ) , .A2( u1_u4_u0_n90 ) , .ZN( u1_u4_u0_n91 ) );
  AND3_X1 u1_u4_u0_U24 (.A3( u1_u4_u0_n121 ) , .A2( u1_u4_u0_n125 ) , .A1( u1_u4_u0_n148 ) , .ZN( u1_u4_u0_n90 ) );
  INV_X1 u1_u4_u0_U25 (.A( u1_u4_u0_n136 ) , .ZN( u1_u4_u0_n161 ) );
  AOI22_X1 u1_u4_u0_U26 (.B2( u1_u4_u0_n109 ) , .A2( u1_u4_u0_n110 ) , .ZN( u1_u4_u0_n111 ) , .B1( u1_u4_u0_n118 ) , .A1( u1_u4_u0_n160 ) );
  INV_X1 u1_u4_u0_U27 (.A( u1_u4_u0_n118 ) , .ZN( u1_u4_u0_n158 ) );
  AOI21_X1 u1_u4_u0_U28 (.ZN( u1_u4_u0_n104 ) , .B1( u1_u4_u0_n107 ) , .B2( u1_u4_u0_n141 ) , .A( u1_u4_u0_n144 ) );
  AOI21_X1 u1_u4_u0_U29 (.B1( u1_u4_u0_n127 ) , .B2( u1_u4_u0_n129 ) , .A( u1_u4_u0_n138 ) , .ZN( u1_u4_u0_n96 ) );
  INV_X1 u1_u4_u0_U3 (.A( u1_u4_u0_n113 ) , .ZN( u1_u4_u0_n166 ) );
  AOI21_X1 u1_u4_u0_U30 (.ZN( u1_u4_u0_n116 ) , .B2( u1_u4_u0_n142 ) , .A( u1_u4_u0_n144 ) , .B1( u1_u4_u0_n166 ) );
  NAND2_X1 u1_u4_u0_U31 (.A1( u1_u4_u0_n100 ) , .A2( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n125 ) );
  NAND2_X1 u1_u4_u0_U32 (.A1( u1_u4_u0_n101 ) , .A2( u1_u4_u0_n102 ) , .ZN( u1_u4_u0_n150 ) );
  INV_X1 u1_u4_u0_U33 (.A( u1_u4_u0_n138 ) , .ZN( u1_u4_u0_n160 ) );
  NAND2_X1 u1_u4_u0_U34 (.A1( u1_u4_u0_n102 ) , .ZN( u1_u4_u0_n128 ) , .A2( u1_u4_u0_n95 ) );
  NAND2_X1 u1_u4_u0_U35 (.A1( u1_u4_u0_n100 ) , .ZN( u1_u4_u0_n129 ) , .A2( u1_u4_u0_n95 ) );
  NAND2_X1 u1_u4_u0_U36 (.A2( u1_u4_u0_n100 ) , .ZN( u1_u4_u0_n131 ) , .A1( u1_u4_u0_n92 ) );
  NAND2_X1 u1_u4_u0_U37 (.A2( u1_u4_u0_n100 ) , .A1( u1_u4_u0_n101 ) , .ZN( u1_u4_u0_n139 ) );
  NAND2_X1 u1_u4_u0_U38 (.ZN( u1_u4_u0_n148 ) , .A1( u1_u4_u0_n93 ) , .A2( u1_u4_u0_n95 ) );
  NAND2_X1 u1_u4_u0_U39 (.A2( u1_u4_u0_n102 ) , .A1( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n149 ) );
  AOI21_X1 u1_u4_u0_U4 (.B1( u1_u4_u0_n114 ) , .ZN( u1_u4_u0_n115 ) , .B2( u1_u4_u0_n129 ) , .A( u1_u4_u0_n161 ) );
  NAND2_X1 u1_u4_u0_U40 (.A2( u1_u4_u0_n102 ) , .ZN( u1_u4_u0_n114 ) , .A1( u1_u4_u0_n92 ) );
  NAND2_X1 u1_u4_u0_U41 (.A2( u1_u4_u0_n101 ) , .ZN( u1_u4_u0_n121 ) , .A1( u1_u4_u0_n93 ) );
  INV_X1 u1_u4_u0_U42 (.ZN( u1_u4_u0_n172 ) , .A( u1_u4_u0_n88 ) );
  OAI222_X1 u1_u4_u0_U43 (.C1( u1_u4_u0_n108 ) , .A1( u1_u4_u0_n125 ) , .B2( u1_u4_u0_n128 ) , .B1( u1_u4_u0_n144 ) , .A2( u1_u4_u0_n158 ) , .C2( u1_u4_u0_n161 ) , .ZN( u1_u4_u0_n88 ) );
  NAND2_X1 u1_u4_u0_U44 (.ZN( u1_u4_u0_n112 ) , .A2( u1_u4_u0_n92 ) , .A1( u1_u4_u0_n93 ) );
  OR3_X1 u1_u4_u0_U45 (.A3( u1_u4_u0_n152 ) , .A2( u1_u4_u0_n153 ) , .A1( u1_u4_u0_n154 ) , .ZN( u1_u4_u0_n155 ) );
  AOI21_X1 u1_u4_u0_U46 (.A( u1_u4_u0_n144 ) , .B2( u1_u4_u0_n145 ) , .B1( u1_u4_u0_n146 ) , .ZN( u1_u4_u0_n154 ) );
  AOI21_X1 u1_u4_u0_U47 (.B2( u1_u4_u0_n150 ) , .B1( u1_u4_u0_n151 ) , .ZN( u1_u4_u0_n152 ) , .A( u1_u4_u0_n158 ) );
  AOI21_X1 u1_u4_u0_U48 (.A( u1_u4_u0_n147 ) , .B2( u1_u4_u0_n148 ) , .B1( u1_u4_u0_n149 ) , .ZN( u1_u4_u0_n153 ) );
  INV_X1 u1_u4_u0_U49 (.ZN( u1_u4_u0_n171 ) , .A( u1_u4_u0_n99 ) );
  AOI21_X1 u1_u4_u0_U5 (.B2( u1_u4_u0_n131 ) , .ZN( u1_u4_u0_n134 ) , .B1( u1_u4_u0_n151 ) , .A( u1_u4_u0_n158 ) );
  OAI211_X1 u1_u4_u0_U50 (.C2( u1_u4_u0_n140 ) , .C1( u1_u4_u0_n161 ) , .A( u1_u4_u0_n169 ) , .B( u1_u4_u0_n98 ) , .ZN( u1_u4_u0_n99 ) );
  INV_X1 u1_u4_u0_U51 (.ZN( u1_u4_u0_n169 ) , .A( u1_u4_u0_n91 ) );
  AOI211_X1 u1_u4_u0_U52 (.C1( u1_u4_u0_n118 ) , .A( u1_u4_u0_n123 ) , .B( u1_u4_u0_n96 ) , .C2( u1_u4_u0_n97 ) , .ZN( u1_u4_u0_n98 ) );
  NOR2_X1 u1_u4_u0_U53 (.A2( u1_u4_X_6 ) , .ZN( u1_u4_u0_n100 ) , .A1( u1_u4_u0_n162 ) );
  NOR2_X1 u1_u4_u0_U54 (.A2( u1_u4_X_4 ) , .A1( u1_u4_X_5 ) , .ZN( u1_u4_u0_n118 ) );
  NOR2_X1 u1_u4_u0_U55 (.A2( u1_u4_X_2 ) , .ZN( u1_u4_u0_n103 ) , .A1( u1_u4_u0_n164 ) );
  NOR2_X1 u1_u4_u0_U56 (.A2( u1_u4_X_1 ) , .A1( u1_u4_X_2 ) , .ZN( u1_u4_u0_n92 ) );
  NOR2_X1 u1_u4_u0_U57 (.A2( u1_u4_X_1 ) , .ZN( u1_u4_u0_n101 ) , .A1( u1_u4_u0_n163 ) );
  NAND2_X1 u1_u4_u0_U58 (.A2( u1_u4_X_4 ) , .A1( u1_u4_X_5 ) , .ZN( u1_u4_u0_n144 ) );
  NOR2_X1 u1_u4_u0_U59 (.A2( u1_u4_X_5 ) , .ZN( u1_u4_u0_n136 ) , .A1( u1_u4_u0_n159 ) );
  NOR2_X1 u1_u4_u0_U6 (.A1( u1_u4_u0_n108 ) , .ZN( u1_u4_u0_n123 ) , .A2( u1_u4_u0_n158 ) );
  NAND2_X1 u1_u4_u0_U60 (.A1( u1_u4_X_5 ) , .ZN( u1_u4_u0_n138 ) , .A2( u1_u4_u0_n159 ) );
  NOR2_X1 u1_u4_u0_U61 (.A2( u1_u4_X_3 ) , .A1( u1_u4_X_6 ) , .ZN( u1_u4_u0_n94 ) );
  AND2_X1 u1_u4_u0_U62 (.A2( u1_u4_X_3 ) , .A1( u1_u4_X_6 ) , .ZN( u1_u4_u0_n102 ) );
  AND2_X1 u1_u4_u0_U63 (.A1( u1_u4_X_6 ) , .A2( u1_u4_u0_n162 ) , .ZN( u1_u4_u0_n93 ) );
  INV_X1 u1_u4_u0_U64 (.A( u1_u4_X_4 ) , .ZN( u1_u4_u0_n159 ) );
  INV_X1 u1_u4_u0_U65 (.A( u1_u4_X_1 ) , .ZN( u1_u4_u0_n164 ) );
  INV_X1 u1_u4_u0_U66 (.A( u1_u4_X_2 ) , .ZN( u1_u4_u0_n163 ) );
  INV_X1 u1_u4_u0_U67 (.A( u1_u4_X_3 ) , .ZN( u1_u4_u0_n162 ) );
  INV_X1 u1_u4_u0_U68 (.A( u1_u4_u0_n126 ) , .ZN( u1_u4_u0_n168 ) );
  AOI211_X1 u1_u4_u0_U69 (.B( u1_u4_u0_n133 ) , .A( u1_u4_u0_n134 ) , .C2( u1_u4_u0_n135 ) , .C1( u1_u4_u0_n136 ) , .ZN( u1_u4_u0_n137 ) );
  OAI21_X1 u1_u4_u0_U7 (.B1( u1_u4_u0_n150 ) , .B2( u1_u4_u0_n158 ) , .A( u1_u4_u0_n172 ) , .ZN( u1_u4_u0_n89 ) );
  AOI21_X1 u1_u4_u0_U70 (.B2( u1_u4_u0_n107 ) , .ZN( u1_u4_u0_n124 ) , .B1( u1_u4_u0_n128 ) , .A( u1_u4_u0_n161 ) );
  INV_X1 u1_u4_u0_U71 (.A( u1_u4_u0_n111 ) , .ZN( u1_u4_u0_n170 ) );
  OR4_X1 u1_u4_u0_U72 (.ZN( u1_out4_31 ) , .A4( u1_u4_u0_n155 ) , .A2( u1_u4_u0_n156 ) , .A1( u1_u4_u0_n157 ) , .A3( u1_u4_u0_n173 ) );
  AOI21_X1 u1_u4_u0_U73 (.A( u1_u4_u0_n138 ) , .B2( u1_u4_u0_n139 ) , .B1( u1_u4_u0_n140 ) , .ZN( u1_u4_u0_n157 ) );
  AOI21_X1 u1_u4_u0_U74 (.B2( u1_u4_u0_n141 ) , .B1( u1_u4_u0_n142 ) , .ZN( u1_u4_u0_n156 ) , .A( u1_u4_u0_n161 ) );
  INV_X1 u1_u4_u0_U75 (.ZN( u1_u4_u0_n174 ) , .A( u1_u4_u0_n89 ) );
  AOI211_X1 u1_u4_u0_U76 (.B( u1_u4_u0_n104 ) , .A( u1_u4_u0_n105 ) , .ZN( u1_u4_u0_n106 ) , .C2( u1_u4_u0_n113 ) , .C1( u1_u4_u0_n160 ) );
  OR4_X1 u1_u4_u0_U77 (.ZN( u1_out4_17 ) , .A4( u1_u4_u0_n122 ) , .A2( u1_u4_u0_n123 ) , .A1( u1_u4_u0_n124 ) , .A3( u1_u4_u0_n170 ) );
  OAI221_X1 u1_u4_u0_U78 (.C1( u1_u4_u0_n121 ) , .ZN( u1_u4_u0_n122 ) , .B2( u1_u4_u0_n127 ) , .A( u1_u4_u0_n143 ) , .B1( u1_u4_u0_n144 ) , .C2( u1_u4_u0_n147 ) );
  NOR2_X1 u1_u4_u0_U79 (.A1( u1_u4_u0_n120 ) , .ZN( u1_u4_u0_n143 ) , .A2( u1_u4_u0_n167 ) );
  AND2_X1 u1_u4_u0_U8 (.A1( u1_u4_u0_n114 ) , .A2( u1_u4_u0_n121 ) , .ZN( u1_u4_u0_n146 ) );
  AOI21_X1 u1_u4_u0_U80 (.B1( u1_u4_u0_n132 ) , .ZN( u1_u4_u0_n133 ) , .A( u1_u4_u0_n144 ) , .B2( u1_u4_u0_n166 ) );
  OAI22_X1 u1_u4_u0_U81 (.ZN( u1_u4_u0_n105 ) , .A2( u1_u4_u0_n132 ) , .B1( u1_u4_u0_n146 ) , .A1( u1_u4_u0_n147 ) , .B2( u1_u4_u0_n161 ) );
  NAND2_X1 u1_u4_u0_U82 (.ZN( u1_u4_u0_n110 ) , .A2( u1_u4_u0_n132 ) , .A1( u1_u4_u0_n145 ) );
  INV_X1 u1_u4_u0_U83 (.A( u1_u4_u0_n119 ) , .ZN( u1_u4_u0_n167 ) );
  NAND2_X1 u1_u4_u0_U84 (.A2( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n140 ) , .A1( u1_u4_u0_n94 ) );
  NAND2_X1 u1_u4_u0_U85 (.A1( u1_u4_u0_n101 ) , .ZN( u1_u4_u0_n130 ) , .A2( u1_u4_u0_n94 ) );
  NAND2_X1 u1_u4_u0_U86 (.ZN( u1_u4_u0_n108 ) , .A1( u1_u4_u0_n92 ) , .A2( u1_u4_u0_n94 ) );
  NAND2_X1 u1_u4_u0_U87 (.ZN( u1_u4_u0_n142 ) , .A1( u1_u4_u0_n94 ) , .A2( u1_u4_u0_n95 ) );
  NAND3_X1 u1_u4_u0_U88 (.ZN( u1_out4_23 ) , .A3( u1_u4_u0_n137 ) , .A1( u1_u4_u0_n168 ) , .A2( u1_u4_u0_n171 ) );
  NAND3_X1 u1_u4_u0_U89 (.A3( u1_u4_u0_n127 ) , .A2( u1_u4_u0_n128 ) , .ZN( u1_u4_u0_n135 ) , .A1( u1_u4_u0_n150 ) );
  AND2_X1 u1_u4_u0_U9 (.A1( u1_u4_u0_n131 ) , .ZN( u1_u4_u0_n141 ) , .A2( u1_u4_u0_n150 ) );
  NAND3_X1 u1_u4_u0_U90 (.ZN( u1_u4_u0_n117 ) , .A3( u1_u4_u0_n132 ) , .A2( u1_u4_u0_n139 ) , .A1( u1_u4_u0_n148 ) );
  NAND3_X1 u1_u4_u0_U91 (.ZN( u1_u4_u0_n109 ) , .A2( u1_u4_u0_n114 ) , .A3( u1_u4_u0_n140 ) , .A1( u1_u4_u0_n149 ) );
  NAND3_X1 u1_u4_u0_U92 (.ZN( u1_out4_9 ) , .A3( u1_u4_u0_n106 ) , .A2( u1_u4_u0_n171 ) , .A1( u1_u4_u0_n174 ) );
  NAND3_X1 u1_u4_u0_U93 (.A2( u1_u4_u0_n128 ) , .A1( u1_u4_u0_n132 ) , .A3( u1_u4_u0_n146 ) , .ZN( u1_u4_u0_n97 ) );
  NOR2_X1 u1_u4_u1_U10 (.A1( u1_u4_u1_n112 ) , .A2( u1_u4_u1_n116 ) , .ZN( u1_u4_u1_n118 ) );
  NAND3_X1 u1_u4_u1_U100 (.ZN( u1_u4_u1_n113 ) , .A1( u1_u4_u1_n120 ) , .A3( u1_u4_u1_n133 ) , .A2( u1_u4_u1_n155 ) );
  OAI21_X1 u1_u4_u1_U11 (.ZN( u1_u4_u1_n101 ) , .B1( u1_u4_u1_n141 ) , .A( u1_u4_u1_n146 ) , .B2( u1_u4_u1_n183 ) );
  AOI21_X1 u1_u4_u1_U12 (.B2( u1_u4_u1_n155 ) , .B1( u1_u4_u1_n156 ) , .ZN( u1_u4_u1_n157 ) , .A( u1_u4_u1_n174 ) );
  NAND2_X1 u1_u4_u1_U13 (.ZN( u1_u4_u1_n140 ) , .A2( u1_u4_u1_n150 ) , .A1( u1_u4_u1_n155 ) );
  NAND2_X1 u1_u4_u1_U14 (.A1( u1_u4_u1_n131 ) , .ZN( u1_u4_u1_n147 ) , .A2( u1_u4_u1_n153 ) );
  INV_X1 u1_u4_u1_U15 (.A( u1_u4_u1_n139 ) , .ZN( u1_u4_u1_n174 ) );
  OR4_X1 u1_u4_u1_U16 (.A4( u1_u4_u1_n106 ) , .A3( u1_u4_u1_n107 ) , .ZN( u1_u4_u1_n108 ) , .A1( u1_u4_u1_n117 ) , .A2( u1_u4_u1_n184 ) );
  AOI21_X1 u1_u4_u1_U17 (.ZN( u1_u4_u1_n106 ) , .A( u1_u4_u1_n112 ) , .B1( u1_u4_u1_n154 ) , .B2( u1_u4_u1_n156 ) );
  AOI21_X1 u1_u4_u1_U18 (.ZN( u1_u4_u1_n107 ) , .B1( u1_u4_u1_n134 ) , .B2( u1_u4_u1_n149 ) , .A( u1_u4_u1_n174 ) );
  INV_X1 u1_u4_u1_U19 (.A( u1_u4_u1_n101 ) , .ZN( u1_u4_u1_n184 ) );
  INV_X1 u1_u4_u1_U20 (.A( u1_u4_u1_n112 ) , .ZN( u1_u4_u1_n171 ) );
  NAND2_X1 u1_u4_u1_U21 (.ZN( u1_u4_u1_n141 ) , .A1( u1_u4_u1_n153 ) , .A2( u1_u4_u1_n156 ) );
  AND2_X1 u1_u4_u1_U22 (.A1( u1_u4_u1_n123 ) , .ZN( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n161 ) );
  NAND2_X1 u1_u4_u1_U23 (.A2( u1_u4_u1_n115 ) , .A1( u1_u4_u1_n116 ) , .ZN( u1_u4_u1_n148 ) );
  NAND2_X1 u1_u4_u1_U24 (.A2( u1_u4_u1_n133 ) , .A1( u1_u4_u1_n135 ) , .ZN( u1_u4_u1_n159 ) );
  NAND2_X1 u1_u4_u1_U25 (.A2( u1_u4_u1_n115 ) , .A1( u1_u4_u1_n120 ) , .ZN( u1_u4_u1_n132 ) );
  INV_X1 u1_u4_u1_U26 (.A( u1_u4_u1_n154 ) , .ZN( u1_u4_u1_n178 ) );
  INV_X1 u1_u4_u1_U27 (.A( u1_u4_u1_n151 ) , .ZN( u1_u4_u1_n183 ) );
  AND2_X1 u1_u4_u1_U28 (.A1( u1_u4_u1_n129 ) , .A2( u1_u4_u1_n133 ) , .ZN( u1_u4_u1_n149 ) );
  INV_X1 u1_u4_u1_U29 (.A( u1_u4_u1_n131 ) , .ZN( u1_u4_u1_n180 ) );
  INV_X1 u1_u4_u1_U3 (.A( u1_u4_u1_n159 ) , .ZN( u1_u4_u1_n182 ) );
  OAI221_X1 u1_u4_u1_U30 (.A( u1_u4_u1_n119 ) , .C2( u1_u4_u1_n129 ) , .ZN( u1_u4_u1_n138 ) , .B2( u1_u4_u1_n152 ) , .C1( u1_u4_u1_n174 ) , .B1( u1_u4_u1_n187 ) );
  INV_X1 u1_u4_u1_U31 (.A( u1_u4_u1_n148 ) , .ZN( u1_u4_u1_n187 ) );
  AOI211_X1 u1_u4_u1_U32 (.B( u1_u4_u1_n117 ) , .A( u1_u4_u1_n118 ) , .ZN( u1_u4_u1_n119 ) , .C2( u1_u4_u1_n146 ) , .C1( u1_u4_u1_n159 ) );
  NOR2_X1 u1_u4_u1_U33 (.A1( u1_u4_u1_n168 ) , .A2( u1_u4_u1_n176 ) , .ZN( u1_u4_u1_n98 ) );
  AOI211_X1 u1_u4_u1_U34 (.B( u1_u4_u1_n162 ) , .A( u1_u4_u1_n163 ) , .C2( u1_u4_u1_n164 ) , .ZN( u1_u4_u1_n165 ) , .C1( u1_u4_u1_n171 ) );
  AOI21_X1 u1_u4_u1_U35 (.A( u1_u4_u1_n160 ) , .B2( u1_u4_u1_n161 ) , .ZN( u1_u4_u1_n162 ) , .B1( u1_u4_u1_n182 ) );
  OR2_X1 u1_u4_u1_U36 (.A2( u1_u4_u1_n157 ) , .A1( u1_u4_u1_n158 ) , .ZN( u1_u4_u1_n163 ) );
  NAND2_X1 u1_u4_u1_U37 (.A1( u1_u4_u1_n128 ) , .ZN( u1_u4_u1_n146 ) , .A2( u1_u4_u1_n160 ) );
  NAND2_X1 u1_u4_u1_U38 (.A2( u1_u4_u1_n112 ) , .ZN( u1_u4_u1_n139 ) , .A1( u1_u4_u1_n152 ) );
  NAND2_X1 u1_u4_u1_U39 (.A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n156 ) , .A2( u1_u4_u1_n99 ) );
  AOI221_X1 u1_u4_u1_U4 (.A( u1_u4_u1_n138 ) , .C2( u1_u4_u1_n139 ) , .C1( u1_u4_u1_n140 ) , .B2( u1_u4_u1_n141 ) , .ZN( u1_u4_u1_n142 ) , .B1( u1_u4_u1_n175 ) );
  AOI221_X1 u1_u4_u1_U40 (.B1( u1_u4_u1_n140 ) , .ZN( u1_u4_u1_n167 ) , .B2( u1_u4_u1_n172 ) , .C2( u1_u4_u1_n175 ) , .C1( u1_u4_u1_n178 ) , .A( u1_u4_u1_n188 ) );
  INV_X1 u1_u4_u1_U41 (.ZN( u1_u4_u1_n188 ) , .A( u1_u4_u1_n97 ) );
  AOI211_X1 u1_u4_u1_U42 (.A( u1_u4_u1_n118 ) , .C1( u1_u4_u1_n132 ) , .C2( u1_u4_u1_n139 ) , .B( u1_u4_u1_n96 ) , .ZN( u1_u4_u1_n97 ) );
  AOI21_X1 u1_u4_u1_U43 (.B2( u1_u4_u1_n121 ) , .B1( u1_u4_u1_n135 ) , .A( u1_u4_u1_n152 ) , .ZN( u1_u4_u1_n96 ) );
  NOR2_X1 u1_u4_u1_U44 (.ZN( u1_u4_u1_n117 ) , .A1( u1_u4_u1_n121 ) , .A2( u1_u4_u1_n160 ) );
  OAI21_X1 u1_u4_u1_U45 (.B2( u1_u4_u1_n123 ) , .ZN( u1_u4_u1_n145 ) , .B1( u1_u4_u1_n160 ) , .A( u1_u4_u1_n185 ) );
  INV_X1 u1_u4_u1_U46 (.A( u1_u4_u1_n122 ) , .ZN( u1_u4_u1_n185 ) );
  AOI21_X1 u1_u4_u1_U47 (.B2( u1_u4_u1_n120 ) , .B1( u1_u4_u1_n121 ) , .ZN( u1_u4_u1_n122 ) , .A( u1_u4_u1_n128 ) );
  AOI21_X1 u1_u4_u1_U48 (.A( u1_u4_u1_n128 ) , .B2( u1_u4_u1_n129 ) , .ZN( u1_u4_u1_n130 ) , .B1( u1_u4_u1_n150 ) );
  NAND2_X1 u1_u4_u1_U49 (.ZN( u1_u4_u1_n112 ) , .A1( u1_u4_u1_n169 ) , .A2( u1_u4_u1_n170 ) );
  AOI211_X1 u1_u4_u1_U5 (.ZN( u1_u4_u1_n124 ) , .A( u1_u4_u1_n138 ) , .C2( u1_u4_u1_n139 ) , .B( u1_u4_u1_n145 ) , .C1( u1_u4_u1_n147 ) );
  NAND2_X1 u1_u4_u1_U50 (.ZN( u1_u4_u1_n129 ) , .A2( u1_u4_u1_n95 ) , .A1( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U51 (.A1( u1_u4_u1_n102 ) , .ZN( u1_u4_u1_n154 ) , .A2( u1_u4_u1_n99 ) );
  NAND2_X1 u1_u4_u1_U52 (.A2( u1_u4_u1_n100 ) , .ZN( u1_u4_u1_n135 ) , .A1( u1_u4_u1_n99 ) );
  AOI21_X1 u1_u4_u1_U53 (.A( u1_u4_u1_n152 ) , .B2( u1_u4_u1_n153 ) , .B1( u1_u4_u1_n154 ) , .ZN( u1_u4_u1_n158 ) );
  INV_X1 u1_u4_u1_U54 (.A( u1_u4_u1_n160 ) , .ZN( u1_u4_u1_n175 ) );
  NAND2_X1 u1_u4_u1_U55 (.A1( u1_u4_u1_n100 ) , .ZN( u1_u4_u1_n116 ) , .A2( u1_u4_u1_n95 ) );
  NAND2_X1 u1_u4_u1_U56 (.A1( u1_u4_u1_n102 ) , .ZN( u1_u4_u1_n131 ) , .A2( u1_u4_u1_n95 ) );
  NAND2_X1 u1_u4_u1_U57 (.A2( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n121 ) , .A1( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U58 (.A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n153 ) , .A2( u1_u4_u1_n98 ) );
  NAND2_X1 u1_u4_u1_U59 (.A2( u1_u4_u1_n104 ) , .A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n133 ) );
  AOI22_X1 u1_u4_u1_U6 (.B2( u1_u4_u1_n113 ) , .A2( u1_u4_u1_n114 ) , .ZN( u1_u4_u1_n125 ) , .A1( u1_u4_u1_n171 ) , .B1( u1_u4_u1_n173 ) );
  NAND2_X1 u1_u4_u1_U60 (.ZN( u1_u4_u1_n150 ) , .A2( u1_u4_u1_n98 ) , .A1( u1_u4_u1_n99 ) );
  NAND2_X1 u1_u4_u1_U61 (.A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n155 ) , .A2( u1_u4_u1_n95 ) );
  OAI21_X1 u1_u4_u1_U62 (.ZN( u1_u4_u1_n109 ) , .B1( u1_u4_u1_n129 ) , .B2( u1_u4_u1_n160 ) , .A( u1_u4_u1_n167 ) );
  NAND2_X1 u1_u4_u1_U63 (.A2( u1_u4_u1_n100 ) , .A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n120 ) );
  NAND2_X1 u1_u4_u1_U64 (.A1( u1_u4_u1_n102 ) , .A2( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n115 ) );
  NAND2_X1 u1_u4_u1_U65 (.A2( u1_u4_u1_n100 ) , .A1( u1_u4_u1_n104 ) , .ZN( u1_u4_u1_n151 ) );
  NAND2_X1 u1_u4_u1_U66 (.A2( u1_u4_u1_n103 ) , .A1( u1_u4_u1_n105 ) , .ZN( u1_u4_u1_n161 ) );
  INV_X1 u1_u4_u1_U67 (.A( u1_u4_u1_n152 ) , .ZN( u1_u4_u1_n173 ) );
  INV_X1 u1_u4_u1_U68 (.A( u1_u4_u1_n128 ) , .ZN( u1_u4_u1_n172 ) );
  NAND2_X1 u1_u4_u1_U69 (.A2( u1_u4_u1_n102 ) , .A1( u1_u4_u1_n103 ) , .ZN( u1_u4_u1_n123 ) );
  NAND2_X1 u1_u4_u1_U7 (.ZN( u1_u4_u1_n114 ) , .A1( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n156 ) );
  NOR2_X1 u1_u4_u1_U70 (.A2( u1_u4_X_7 ) , .A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n95 ) );
  NOR2_X1 u1_u4_u1_U71 (.A1( u1_u4_X_12 ) , .A2( u1_u4_X_9 ) , .ZN( u1_u4_u1_n100 ) );
  NOR2_X1 u1_u4_u1_U72 (.A2( u1_u4_X_8 ) , .A1( u1_u4_u1_n177 ) , .ZN( u1_u4_u1_n99 ) );
  NOR2_X1 u1_u4_u1_U73 (.A2( u1_u4_X_12 ) , .ZN( u1_u4_u1_n102 ) , .A1( u1_u4_u1_n176 ) );
  NOR2_X1 u1_u4_u1_U74 (.A2( u1_u4_X_9 ) , .ZN( u1_u4_u1_n105 ) , .A1( u1_u4_u1_n168 ) );
  NAND2_X1 u1_u4_u1_U75 (.A1( u1_u4_X_10 ) , .ZN( u1_u4_u1_n160 ) , .A2( u1_u4_u1_n169 ) );
  NAND2_X1 u1_u4_u1_U76 (.A2( u1_u4_X_10 ) , .A1( u1_u4_X_11 ) , .ZN( u1_u4_u1_n152 ) );
  NAND2_X1 u1_u4_u1_U77 (.A1( u1_u4_X_11 ) , .ZN( u1_u4_u1_n128 ) , .A2( u1_u4_u1_n170 ) );
  AND2_X1 u1_u4_u1_U78 (.A2( u1_u4_X_7 ) , .A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n104 ) );
  AND2_X1 u1_u4_u1_U79 (.A1( u1_u4_X_8 ) , .ZN( u1_u4_u1_n103 ) , .A2( u1_u4_u1_n177 ) );
  AOI22_X1 u1_u4_u1_U8 (.B2( u1_u4_u1_n136 ) , .A2( u1_u4_u1_n137 ) , .ZN( u1_u4_u1_n143 ) , .A1( u1_u4_u1_n171 ) , .B1( u1_u4_u1_n173 ) );
  INV_X1 u1_u4_u1_U80 (.A( u1_u4_X_10 ) , .ZN( u1_u4_u1_n170 ) );
  INV_X1 u1_u4_u1_U81 (.A( u1_u4_X_9 ) , .ZN( u1_u4_u1_n176 ) );
  INV_X1 u1_u4_u1_U82 (.A( u1_u4_X_11 ) , .ZN( u1_u4_u1_n169 ) );
  INV_X1 u1_u4_u1_U83 (.A( u1_u4_X_12 ) , .ZN( u1_u4_u1_n168 ) );
  INV_X1 u1_u4_u1_U84 (.A( u1_u4_X_7 ) , .ZN( u1_u4_u1_n177 ) );
  NAND4_X1 u1_u4_u1_U85 (.ZN( u1_out4_18 ) , .A4( u1_u4_u1_n165 ) , .A3( u1_u4_u1_n166 ) , .A1( u1_u4_u1_n167 ) , .A2( u1_u4_u1_n186 ) );
  AOI22_X1 u1_u4_u1_U86 (.B2( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n147 ) , .A2( u1_u4_u1_n148 ) , .ZN( u1_u4_u1_n166 ) , .A1( u1_u4_u1_n172 ) );
  INV_X1 u1_u4_u1_U87 (.A( u1_u4_u1_n145 ) , .ZN( u1_u4_u1_n186 ) );
  NAND4_X1 u1_u4_u1_U88 (.ZN( u1_out4_2 ) , .A4( u1_u4_u1_n142 ) , .A3( u1_u4_u1_n143 ) , .A2( u1_u4_u1_n144 ) , .A1( u1_u4_u1_n179 ) );
  OAI21_X1 u1_u4_u1_U89 (.B2( u1_u4_u1_n132 ) , .ZN( u1_u4_u1_n144 ) , .A( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n180 ) );
  INV_X1 u1_u4_u1_U9 (.A( u1_u4_u1_n147 ) , .ZN( u1_u4_u1_n181 ) );
  INV_X1 u1_u4_u1_U90 (.A( u1_u4_u1_n130 ) , .ZN( u1_u4_u1_n179 ) );
  NAND4_X1 u1_u4_u1_U91 (.ZN( u1_out4_28 ) , .A4( u1_u4_u1_n124 ) , .A3( u1_u4_u1_n125 ) , .A2( u1_u4_u1_n126 ) , .A1( u1_u4_u1_n127 ) );
  OAI21_X1 u1_u4_u1_U92 (.ZN( u1_u4_u1_n127 ) , .B2( u1_u4_u1_n139 ) , .B1( u1_u4_u1_n175 ) , .A( u1_u4_u1_n183 ) );
  OAI21_X1 u1_u4_u1_U93 (.ZN( u1_u4_u1_n126 ) , .B2( u1_u4_u1_n140 ) , .A( u1_u4_u1_n146 ) , .B1( u1_u4_u1_n178 ) );
  OR4_X1 u1_u4_u1_U94 (.ZN( u1_out4_13 ) , .A4( u1_u4_u1_n108 ) , .A3( u1_u4_u1_n109 ) , .A2( u1_u4_u1_n110 ) , .A1( u1_u4_u1_n111 ) );
  AOI21_X1 u1_u4_u1_U95 (.ZN( u1_u4_u1_n111 ) , .A( u1_u4_u1_n128 ) , .B2( u1_u4_u1_n131 ) , .B1( u1_u4_u1_n135 ) );
  AOI21_X1 u1_u4_u1_U96 (.ZN( u1_u4_u1_n110 ) , .A( u1_u4_u1_n116 ) , .B1( u1_u4_u1_n152 ) , .B2( u1_u4_u1_n160 ) );
  NAND3_X1 u1_u4_u1_U97 (.A3( u1_u4_u1_n149 ) , .A2( u1_u4_u1_n150 ) , .A1( u1_u4_u1_n151 ) , .ZN( u1_u4_u1_n164 ) );
  NAND3_X1 u1_u4_u1_U98 (.A3( u1_u4_u1_n134 ) , .A2( u1_u4_u1_n135 ) , .ZN( u1_u4_u1_n136 ) , .A1( u1_u4_u1_n151 ) );
  NAND3_X1 u1_u4_u1_U99 (.A1( u1_u4_u1_n133 ) , .ZN( u1_u4_u1_n137 ) , .A2( u1_u4_u1_n154 ) , .A3( u1_u4_u1_n181 ) );
  OAI22_X1 u1_u4_u3_U10 (.B1( u1_u4_u3_n113 ) , .A2( u1_u4_u3_n135 ) , .A1( u1_u4_u3_n150 ) , .B2( u1_u4_u3_n164 ) , .ZN( u1_u4_u3_n98 ) );
  OAI211_X1 u1_u4_u3_U11 (.B( u1_u4_u3_n106 ) , .ZN( u1_u4_u3_n119 ) , .C2( u1_u4_u3_n128 ) , .C1( u1_u4_u3_n167 ) , .A( u1_u4_u3_n181 ) );
  AOI221_X1 u1_u4_u3_U12 (.C1( u1_u4_u3_n105 ) , .ZN( u1_u4_u3_n106 ) , .A( u1_u4_u3_n131 ) , .B2( u1_u4_u3_n132 ) , .C2( u1_u4_u3_n133 ) , .B1( u1_u4_u3_n169 ) );
  INV_X1 u1_u4_u3_U13 (.ZN( u1_u4_u3_n181 ) , .A( u1_u4_u3_n98 ) );
  NAND2_X1 u1_u4_u3_U14 (.ZN( u1_u4_u3_n105 ) , .A2( u1_u4_u3_n130 ) , .A1( u1_u4_u3_n155 ) );
  AOI22_X1 u1_u4_u3_U15 (.B1( u1_u4_u3_n115 ) , .A2( u1_u4_u3_n116 ) , .ZN( u1_u4_u3_n123 ) , .B2( u1_u4_u3_n133 ) , .A1( u1_u4_u3_n169 ) );
  NAND2_X1 u1_u4_u3_U16 (.ZN( u1_u4_u3_n116 ) , .A2( u1_u4_u3_n151 ) , .A1( u1_u4_u3_n182 ) );
  NOR2_X1 u1_u4_u3_U17 (.ZN( u1_u4_u3_n126 ) , .A2( u1_u4_u3_n150 ) , .A1( u1_u4_u3_n164 ) );
  AOI21_X1 u1_u4_u3_U18 (.ZN( u1_u4_u3_n112 ) , .B2( u1_u4_u3_n146 ) , .B1( u1_u4_u3_n155 ) , .A( u1_u4_u3_n167 ) );
  NAND2_X1 u1_u4_u3_U19 (.A1( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n142 ) , .A2( u1_u4_u3_n164 ) );
  NAND2_X1 u1_u4_u3_U20 (.ZN( u1_u4_u3_n132 ) , .A2( u1_u4_u3_n152 ) , .A1( u1_u4_u3_n156 ) );
  AND2_X1 u1_u4_u3_U21 (.A2( u1_u4_u3_n113 ) , .A1( u1_u4_u3_n114 ) , .ZN( u1_u4_u3_n151 ) );
  INV_X1 u1_u4_u3_U22 (.A( u1_u4_u3_n133 ) , .ZN( u1_u4_u3_n165 ) );
  INV_X1 u1_u4_u3_U23 (.A( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n170 ) );
  NAND2_X1 u1_u4_u3_U24 (.A1( u1_u4_u3_n107 ) , .A2( u1_u4_u3_n108 ) , .ZN( u1_u4_u3_n140 ) );
  NAND2_X1 u1_u4_u3_U25 (.ZN( u1_u4_u3_n117 ) , .A1( u1_u4_u3_n124 ) , .A2( u1_u4_u3_n148 ) );
  NAND2_X1 u1_u4_u3_U26 (.ZN( u1_u4_u3_n143 ) , .A1( u1_u4_u3_n165 ) , .A2( u1_u4_u3_n167 ) );
  INV_X1 u1_u4_u3_U27 (.A( u1_u4_u3_n130 ) , .ZN( u1_u4_u3_n177 ) );
  INV_X1 u1_u4_u3_U28 (.A( u1_u4_u3_n128 ) , .ZN( u1_u4_u3_n176 ) );
  INV_X1 u1_u4_u3_U29 (.A( u1_u4_u3_n155 ) , .ZN( u1_u4_u3_n174 ) );
  INV_X1 u1_u4_u3_U3 (.A( u1_u4_u3_n129 ) , .ZN( u1_u4_u3_n183 ) );
  INV_X1 u1_u4_u3_U30 (.A( u1_u4_u3_n139 ) , .ZN( u1_u4_u3_n185 ) );
  NOR2_X1 u1_u4_u3_U31 (.ZN( u1_u4_u3_n135 ) , .A2( u1_u4_u3_n141 ) , .A1( u1_u4_u3_n169 ) );
  OAI222_X1 u1_u4_u3_U32 (.C2( u1_u4_u3_n107 ) , .A2( u1_u4_u3_n108 ) , .B1( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n138 ) , .B2( u1_u4_u3_n146 ) , .C1( u1_u4_u3_n154 ) , .A1( u1_u4_u3_n164 ) );
  NOR4_X1 u1_u4_u3_U33 (.A4( u1_u4_u3_n157 ) , .A3( u1_u4_u3_n158 ) , .A2( u1_u4_u3_n159 ) , .A1( u1_u4_u3_n160 ) , .ZN( u1_u4_u3_n161 ) );
  AOI21_X1 u1_u4_u3_U34 (.B2( u1_u4_u3_n152 ) , .B1( u1_u4_u3_n153 ) , .ZN( u1_u4_u3_n158 ) , .A( u1_u4_u3_n164 ) );
  AOI21_X1 u1_u4_u3_U35 (.A( u1_u4_u3_n149 ) , .B2( u1_u4_u3_n150 ) , .B1( u1_u4_u3_n151 ) , .ZN( u1_u4_u3_n159 ) );
  AOI21_X1 u1_u4_u3_U36 (.A( u1_u4_u3_n154 ) , .B2( u1_u4_u3_n155 ) , .B1( u1_u4_u3_n156 ) , .ZN( u1_u4_u3_n157 ) );
  AOI211_X1 u1_u4_u3_U37 (.ZN( u1_u4_u3_n109 ) , .A( u1_u4_u3_n119 ) , .C2( u1_u4_u3_n129 ) , .B( u1_u4_u3_n138 ) , .C1( u1_u4_u3_n141 ) );
  AOI211_X1 u1_u4_u3_U38 (.B( u1_u4_u3_n119 ) , .A( u1_u4_u3_n120 ) , .C2( u1_u4_u3_n121 ) , .ZN( u1_u4_u3_n122 ) , .C1( u1_u4_u3_n179 ) );
  INV_X1 u1_u4_u3_U39 (.A( u1_u4_u3_n156 ) , .ZN( u1_u4_u3_n179 ) );
  INV_X1 u1_u4_u3_U4 (.A( u1_u4_u3_n140 ) , .ZN( u1_u4_u3_n182 ) );
  OAI22_X1 u1_u4_u3_U40 (.B1( u1_u4_u3_n118 ) , .ZN( u1_u4_u3_n120 ) , .A1( u1_u4_u3_n135 ) , .B2( u1_u4_u3_n154 ) , .A2( u1_u4_u3_n178 ) );
  AND3_X1 u1_u4_u3_U41 (.ZN( u1_u4_u3_n118 ) , .A2( u1_u4_u3_n124 ) , .A1( u1_u4_u3_n144 ) , .A3( u1_u4_u3_n152 ) );
  INV_X1 u1_u4_u3_U42 (.A( u1_u4_u3_n121 ) , .ZN( u1_u4_u3_n164 ) );
  NAND2_X1 u1_u4_u3_U43 (.ZN( u1_u4_u3_n133 ) , .A1( u1_u4_u3_n154 ) , .A2( u1_u4_u3_n164 ) );
  OAI211_X1 u1_u4_u3_U44 (.B( u1_u4_u3_n127 ) , .ZN( u1_u4_u3_n139 ) , .C1( u1_u4_u3_n150 ) , .C2( u1_u4_u3_n154 ) , .A( u1_u4_u3_n184 ) );
  INV_X1 u1_u4_u3_U45 (.A( u1_u4_u3_n125 ) , .ZN( u1_u4_u3_n184 ) );
  AOI221_X1 u1_u4_u3_U46 (.A( u1_u4_u3_n126 ) , .ZN( u1_u4_u3_n127 ) , .C2( u1_u4_u3_n132 ) , .C1( u1_u4_u3_n169 ) , .B2( u1_u4_u3_n170 ) , .B1( u1_u4_u3_n174 ) );
  OAI22_X1 u1_u4_u3_U47 (.A1( u1_u4_u3_n124 ) , .ZN( u1_u4_u3_n125 ) , .B2( u1_u4_u3_n145 ) , .A2( u1_u4_u3_n165 ) , .B1( u1_u4_u3_n167 ) );
  NOR2_X1 u1_u4_u3_U48 (.A1( u1_u4_u3_n113 ) , .ZN( u1_u4_u3_n131 ) , .A2( u1_u4_u3_n154 ) );
  NAND2_X1 u1_u4_u3_U49 (.A1( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n150 ) , .A2( u1_u4_u3_n99 ) );
  INV_X1 u1_u4_u3_U5 (.A( u1_u4_u3_n117 ) , .ZN( u1_u4_u3_n178 ) );
  NAND2_X1 u1_u4_u3_U50 (.A2( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n155 ) , .A1( u1_u4_u3_n97 ) );
  INV_X1 u1_u4_u3_U51 (.A( u1_u4_u3_n141 ) , .ZN( u1_u4_u3_n167 ) );
  AOI21_X1 u1_u4_u3_U52 (.B2( u1_u4_u3_n114 ) , .B1( u1_u4_u3_n146 ) , .A( u1_u4_u3_n154 ) , .ZN( u1_u4_u3_n94 ) );
  AOI21_X1 u1_u4_u3_U53 (.ZN( u1_u4_u3_n110 ) , .B2( u1_u4_u3_n142 ) , .B1( u1_u4_u3_n186 ) , .A( u1_u4_u3_n95 ) );
  INV_X1 u1_u4_u3_U54 (.A( u1_u4_u3_n145 ) , .ZN( u1_u4_u3_n186 ) );
  AOI21_X1 u1_u4_u3_U55 (.B1( u1_u4_u3_n124 ) , .A( u1_u4_u3_n149 ) , .B2( u1_u4_u3_n155 ) , .ZN( u1_u4_u3_n95 ) );
  INV_X1 u1_u4_u3_U56 (.A( u1_u4_u3_n149 ) , .ZN( u1_u4_u3_n169 ) );
  NAND2_X1 u1_u4_u3_U57 (.ZN( u1_u4_u3_n124 ) , .A1( u1_u4_u3_n96 ) , .A2( u1_u4_u3_n97 ) );
  NAND2_X1 u1_u4_u3_U58 (.A2( u1_u4_u3_n100 ) , .ZN( u1_u4_u3_n146 ) , .A1( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U59 (.A1( u1_u4_u3_n101 ) , .ZN( u1_u4_u3_n145 ) , .A2( u1_u4_u3_n99 ) );
  AOI221_X1 u1_u4_u3_U6 (.A( u1_u4_u3_n131 ) , .C2( u1_u4_u3_n132 ) , .C1( u1_u4_u3_n133 ) , .ZN( u1_u4_u3_n134 ) , .B1( u1_u4_u3_n143 ) , .B2( u1_u4_u3_n177 ) );
  NAND2_X1 u1_u4_u3_U60 (.A1( u1_u4_u3_n100 ) , .ZN( u1_u4_u3_n156 ) , .A2( u1_u4_u3_n99 ) );
  NAND2_X1 u1_u4_u3_U61 (.A2( u1_u4_u3_n101 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n148 ) );
  NAND2_X1 u1_u4_u3_U62 (.A1( u1_u4_u3_n100 ) , .A2( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n128 ) );
  NAND2_X1 u1_u4_u3_U63 (.A2( u1_u4_u3_n101 ) , .A1( u1_u4_u3_n102 ) , .ZN( u1_u4_u3_n152 ) );
  NAND2_X1 u1_u4_u3_U64 (.A2( u1_u4_u3_n101 ) , .ZN( u1_u4_u3_n114 ) , .A1( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U65 (.ZN( u1_u4_u3_n107 ) , .A1( u1_u4_u3_n97 ) , .A2( u1_u4_u3_n99 ) );
  NAND2_X1 u1_u4_u3_U66 (.A2( u1_u4_u3_n100 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n113 ) );
  NAND2_X1 u1_u4_u3_U67 (.A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n153 ) , .A2( u1_u4_u3_n97 ) );
  NAND2_X1 u1_u4_u3_U68 (.A2( u1_u4_u3_n103 ) , .A1( u1_u4_u3_n104 ) , .ZN( u1_u4_u3_n130 ) );
  NAND2_X1 u1_u4_u3_U69 (.A2( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n144 ) , .A1( u1_u4_u3_n96 ) );
  OAI22_X1 u1_u4_u3_U7 (.B2( u1_u4_u3_n147 ) , .A2( u1_u4_u3_n148 ) , .ZN( u1_u4_u3_n160 ) , .B1( u1_u4_u3_n165 ) , .A1( u1_u4_u3_n168 ) );
  NAND2_X1 u1_u4_u3_U70 (.A1( u1_u4_u3_n102 ) , .A2( u1_u4_u3_n103 ) , .ZN( u1_u4_u3_n108 ) );
  NOR2_X1 u1_u4_u3_U71 (.A2( u1_u4_X_19 ) , .A1( u1_u4_X_20 ) , .ZN( u1_u4_u3_n99 ) );
  NOR2_X1 u1_u4_u3_U72 (.A2( u1_u4_X_21 ) , .A1( u1_u4_X_24 ) , .ZN( u1_u4_u3_n103 ) );
  NOR2_X1 u1_u4_u3_U73 (.A2( u1_u4_X_24 ) , .A1( u1_u4_u3_n171 ) , .ZN( u1_u4_u3_n97 ) );
  NOR2_X1 u1_u4_u3_U74 (.A2( u1_u4_X_23 ) , .ZN( u1_u4_u3_n141 ) , .A1( u1_u4_u3_n166 ) );
  NOR2_X1 u1_u4_u3_U75 (.A2( u1_u4_X_19 ) , .A1( u1_u4_u3_n172 ) , .ZN( u1_u4_u3_n96 ) );
  NAND2_X1 u1_u4_u3_U76 (.A1( u1_u4_X_22 ) , .A2( u1_u4_X_23 ) , .ZN( u1_u4_u3_n154 ) );
  NAND2_X1 u1_u4_u3_U77 (.A1( u1_u4_X_23 ) , .ZN( u1_u4_u3_n149 ) , .A2( u1_u4_u3_n166 ) );
  NOR2_X1 u1_u4_u3_U78 (.A2( u1_u4_X_22 ) , .A1( u1_u4_X_23 ) , .ZN( u1_u4_u3_n121 ) );
  AND2_X1 u1_u4_u3_U79 (.A1( u1_u4_X_24 ) , .ZN( u1_u4_u3_n101 ) , .A2( u1_u4_u3_n171 ) );
  AND3_X1 u1_u4_u3_U8 (.A3( u1_u4_u3_n144 ) , .A2( u1_u4_u3_n145 ) , .A1( u1_u4_u3_n146 ) , .ZN( u1_u4_u3_n147 ) );
  AND2_X1 u1_u4_u3_U80 (.A1( u1_u4_X_19 ) , .ZN( u1_u4_u3_n102 ) , .A2( u1_u4_u3_n172 ) );
  AND2_X1 u1_u4_u3_U81 (.A1( u1_u4_X_21 ) , .A2( u1_u4_X_24 ) , .ZN( u1_u4_u3_n100 ) );
  AND2_X1 u1_u4_u3_U82 (.A2( u1_u4_X_19 ) , .A1( u1_u4_X_20 ) , .ZN( u1_u4_u3_n104 ) );
  INV_X1 u1_u4_u3_U83 (.A( u1_u4_X_22 ) , .ZN( u1_u4_u3_n166 ) );
  INV_X1 u1_u4_u3_U84 (.A( u1_u4_X_21 ) , .ZN( u1_u4_u3_n171 ) );
  INV_X1 u1_u4_u3_U85 (.A( u1_u4_X_20 ) , .ZN( u1_u4_u3_n172 ) );
  NAND4_X1 u1_u4_u3_U86 (.ZN( u1_out4_26 ) , .A4( u1_u4_u3_n109 ) , .A3( u1_u4_u3_n110 ) , .A2( u1_u4_u3_n111 ) , .A1( u1_u4_u3_n173 ) );
  INV_X1 u1_u4_u3_U87 (.ZN( u1_u4_u3_n173 ) , .A( u1_u4_u3_n94 ) );
  OAI21_X1 u1_u4_u3_U88 (.ZN( u1_u4_u3_n111 ) , .B2( u1_u4_u3_n117 ) , .A( u1_u4_u3_n133 ) , .B1( u1_u4_u3_n176 ) );
  NAND4_X1 u1_u4_u3_U89 (.ZN( u1_out4_20 ) , .A4( u1_u4_u3_n122 ) , .A3( u1_u4_u3_n123 ) , .A1( u1_u4_u3_n175 ) , .A2( u1_u4_u3_n180 ) );
  INV_X1 u1_u4_u3_U9 (.A( u1_u4_u3_n143 ) , .ZN( u1_u4_u3_n168 ) );
  INV_X1 u1_u4_u3_U90 (.A( u1_u4_u3_n126 ) , .ZN( u1_u4_u3_n180 ) );
  INV_X1 u1_u4_u3_U91 (.A( u1_u4_u3_n112 ) , .ZN( u1_u4_u3_n175 ) );
  NAND4_X1 u1_u4_u3_U92 (.ZN( u1_out4_1 ) , .A4( u1_u4_u3_n161 ) , .A3( u1_u4_u3_n162 ) , .A2( u1_u4_u3_n163 ) , .A1( u1_u4_u3_n185 ) );
  NAND2_X1 u1_u4_u3_U93 (.ZN( u1_u4_u3_n163 ) , .A2( u1_u4_u3_n170 ) , .A1( u1_u4_u3_n176 ) );
  AOI22_X1 u1_u4_u3_U94 (.B2( u1_u4_u3_n140 ) , .B1( u1_u4_u3_n141 ) , .A2( u1_u4_u3_n142 ) , .ZN( u1_u4_u3_n162 ) , .A1( u1_u4_u3_n177 ) );
  OR4_X1 u1_u4_u3_U95 (.ZN( u1_out4_10 ) , .A4( u1_u4_u3_n136 ) , .A3( u1_u4_u3_n137 ) , .A1( u1_u4_u3_n138 ) , .A2( u1_u4_u3_n139 ) );
  OAI222_X1 u1_u4_u3_U96 (.C1( u1_u4_u3_n128 ) , .ZN( u1_u4_u3_n137 ) , .B1( u1_u4_u3_n148 ) , .A2( u1_u4_u3_n150 ) , .B2( u1_u4_u3_n154 ) , .C2( u1_u4_u3_n164 ) , .A1( u1_u4_u3_n167 ) );
  OAI221_X1 u1_u4_u3_U97 (.A( u1_u4_u3_n134 ) , .B2( u1_u4_u3_n135 ) , .ZN( u1_u4_u3_n136 ) , .C1( u1_u4_u3_n149 ) , .B1( u1_u4_u3_n151 ) , .C2( u1_u4_u3_n183 ) );
  NAND3_X1 u1_u4_u3_U98 (.A1( u1_u4_u3_n114 ) , .ZN( u1_u4_u3_n115 ) , .A2( u1_u4_u3_n145 ) , .A3( u1_u4_u3_n153 ) );
  NAND3_X1 u1_u4_u3_U99 (.ZN( u1_u4_u3_n129 ) , .A2( u1_u4_u3_n144 ) , .A1( u1_u4_u3_n153 ) , .A3( u1_u4_u3_n182 ) );
  XOR2_X1 u1_u6_U15 (.B( u1_K7_40 ) , .A( u1_R5_27 ) , .Z( u1_u6_X_40 ) );
  XOR2_X1 u1_u6_U16 (.B( u1_K7_3 ) , .A( u1_R5_2 ) , .Z( u1_u6_X_3 ) );
  XOR2_X1 u1_u6_U17 (.B( u1_K7_39 ) , .A( u1_R5_26 ) , .Z( u1_u6_X_39 ) );
  XOR2_X1 u1_u6_U29 (.B( u1_K7_28 ) , .A( u1_R5_19 ) , .Z( u1_u6_X_28 ) );
  XOR2_X1 u1_u6_U30 (.B( u1_K7_27 ) , .A( u1_R5_18 ) , .Z( u1_u6_X_27 ) );
  XOR2_X1 u1_u6_U6 (.B( u1_K7_4 ) , .A( u1_R5_3 ) , .Z( u1_u6_X_4 ) );
  AND3_X1 u1_u6_u0_U10 (.A2( u1_u6_u0_n112 ) , .ZN( u1_u6_u0_n127 ) , .A3( u1_u6_u0_n130 ) , .A1( u1_u6_u0_n148 ) );
  NAND2_X1 u1_u6_u0_U11 (.ZN( u1_u6_u0_n113 ) , .A1( u1_u6_u0_n139 ) , .A2( u1_u6_u0_n149 ) );
  AND2_X1 u1_u6_u0_U12 (.ZN( u1_u6_u0_n107 ) , .A1( u1_u6_u0_n130 ) , .A2( u1_u6_u0_n140 ) );
  AND2_X1 u1_u6_u0_U13 (.A2( u1_u6_u0_n129 ) , .A1( u1_u6_u0_n130 ) , .ZN( u1_u6_u0_n151 ) );
  AND2_X1 u1_u6_u0_U14 (.A1( u1_u6_u0_n108 ) , .A2( u1_u6_u0_n125 ) , .ZN( u1_u6_u0_n145 ) );
  INV_X1 u1_u6_u0_U15 (.A( u1_u6_u0_n143 ) , .ZN( u1_u6_u0_n173 ) );
  NOR2_X1 u1_u6_u0_U16 (.A2( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n147 ) , .A1( u1_u6_u0_n160 ) );
  NOR2_X1 u1_u6_u0_U17 (.A1( u1_u6_u0_n163 ) , .A2( u1_u6_u0_n164 ) , .ZN( u1_u6_u0_n95 ) );
  AOI21_X1 u1_u6_u0_U18 (.B1( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n132 ) , .A( u1_u6_u0_n165 ) , .B2( u1_u6_u0_n93 ) );
  INV_X1 u1_u6_u0_U19 (.A( u1_u6_u0_n142 ) , .ZN( u1_u6_u0_n165 ) );
  OAI221_X1 u1_u6_u0_U20 (.C1( u1_u6_u0_n112 ) , .ZN( u1_u6_u0_n120 ) , .B1( u1_u6_u0_n138 ) , .B2( u1_u6_u0_n141 ) , .C2( u1_u6_u0_n147 ) , .A( u1_u6_u0_n172 ) );
  AOI211_X1 u1_u6_u0_U21 (.B( u1_u6_u0_n115 ) , .A( u1_u6_u0_n116 ) , .C2( u1_u6_u0_n117 ) , .C1( u1_u6_u0_n118 ) , .ZN( u1_u6_u0_n119 ) );
  OAI22_X1 u1_u6_u0_U22 (.B1( u1_u6_u0_n125 ) , .ZN( u1_u6_u0_n126 ) , .A1( u1_u6_u0_n138 ) , .A2( u1_u6_u0_n146 ) , .B2( u1_u6_u0_n147 ) );
  OAI22_X1 u1_u6_u0_U23 (.B1( u1_u6_u0_n131 ) , .A1( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n147 ) , .A2( u1_u6_u0_n90 ) , .ZN( u1_u6_u0_n91 ) );
  AND3_X1 u1_u6_u0_U24 (.A3( u1_u6_u0_n121 ) , .A2( u1_u6_u0_n125 ) , .A1( u1_u6_u0_n148 ) , .ZN( u1_u6_u0_n90 ) );
  NAND2_X1 u1_u6_u0_U25 (.A1( u1_u6_u0_n100 ) , .A2( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n125 ) );
  INV_X1 u1_u6_u0_U26 (.A( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n161 ) );
  AOI22_X1 u1_u6_u0_U27 (.B2( u1_u6_u0_n109 ) , .A2( u1_u6_u0_n110 ) , .ZN( u1_u6_u0_n111 ) , .B1( u1_u6_u0_n118 ) , .A1( u1_u6_u0_n160 ) );
  NAND2_X1 u1_u6_u0_U28 (.A1( u1_u6_u0_n100 ) , .ZN( u1_u6_u0_n129 ) , .A2( u1_u6_u0_n95 ) );
  INV_X1 u1_u6_u0_U29 (.A( u1_u6_u0_n118 ) , .ZN( u1_u6_u0_n158 ) );
  INV_X1 u1_u6_u0_U3 (.A( u1_u6_u0_n113 ) , .ZN( u1_u6_u0_n166 ) );
  AOI21_X1 u1_u6_u0_U30 (.ZN( u1_u6_u0_n104 ) , .B1( u1_u6_u0_n107 ) , .B2( u1_u6_u0_n141 ) , .A( u1_u6_u0_n144 ) );
  AOI21_X1 u1_u6_u0_U31 (.B1( u1_u6_u0_n127 ) , .B2( u1_u6_u0_n129 ) , .A( u1_u6_u0_n138 ) , .ZN( u1_u6_u0_n96 ) );
  AOI21_X1 u1_u6_u0_U32 (.ZN( u1_u6_u0_n116 ) , .B2( u1_u6_u0_n142 ) , .A( u1_u6_u0_n144 ) , .B1( u1_u6_u0_n166 ) );
  NAND2_X1 u1_u6_u0_U33 (.A2( u1_u6_u0_n100 ) , .A1( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n139 ) );
  NAND2_X1 u1_u6_u0_U34 (.A2( u1_u6_u0_n100 ) , .ZN( u1_u6_u0_n131 ) , .A1( u1_u6_u0_n92 ) );
  NAND2_X1 u1_u6_u0_U35 (.A1( u1_u6_u0_n101 ) , .A2( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n150 ) );
  INV_X1 u1_u6_u0_U36 (.A( u1_u6_u0_n138 ) , .ZN( u1_u6_u0_n160 ) );
  NAND2_X1 u1_u6_u0_U37 (.A1( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n128 ) , .A2( u1_u6_u0_n95 ) );
  NAND2_X1 u1_u6_u0_U38 (.ZN( u1_u6_u0_n148 ) , .A1( u1_u6_u0_n93 ) , .A2( u1_u6_u0_n95 ) );
  NAND2_X1 u1_u6_u0_U39 (.A2( u1_u6_u0_n102 ) , .A1( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n149 ) );
  AOI21_X1 u1_u6_u0_U4 (.B1( u1_u6_u0_n114 ) , .ZN( u1_u6_u0_n115 ) , .B2( u1_u6_u0_n129 ) , .A( u1_u6_u0_n161 ) );
  NAND2_X1 u1_u6_u0_U40 (.A2( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n114 ) , .A1( u1_u6_u0_n92 ) );
  NAND2_X1 u1_u6_u0_U41 (.A2( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n121 ) , .A1( u1_u6_u0_n93 ) );
  NAND2_X1 u1_u6_u0_U42 (.ZN( u1_u6_u0_n112 ) , .A2( u1_u6_u0_n92 ) , .A1( u1_u6_u0_n93 ) );
  INV_X1 u1_u6_u0_U43 (.ZN( u1_u6_u0_n172 ) , .A( u1_u6_u0_n88 ) );
  OAI222_X1 u1_u6_u0_U44 (.C1( u1_u6_u0_n108 ) , .A1( u1_u6_u0_n125 ) , .B2( u1_u6_u0_n128 ) , .B1( u1_u6_u0_n144 ) , .A2( u1_u6_u0_n158 ) , .C2( u1_u6_u0_n161 ) , .ZN( u1_u6_u0_n88 ) );
  OR3_X1 u1_u6_u0_U45 (.A3( u1_u6_u0_n152 ) , .A2( u1_u6_u0_n153 ) , .A1( u1_u6_u0_n154 ) , .ZN( u1_u6_u0_n155 ) );
  AOI21_X1 u1_u6_u0_U46 (.A( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n145 ) , .B1( u1_u6_u0_n146 ) , .ZN( u1_u6_u0_n154 ) );
  AOI21_X1 u1_u6_u0_U47 (.B2( u1_u6_u0_n150 ) , .B1( u1_u6_u0_n151 ) , .ZN( u1_u6_u0_n152 ) , .A( u1_u6_u0_n158 ) );
  AOI21_X1 u1_u6_u0_U48 (.A( u1_u6_u0_n147 ) , .B2( u1_u6_u0_n148 ) , .B1( u1_u6_u0_n149 ) , .ZN( u1_u6_u0_n153 ) );
  INV_X1 u1_u6_u0_U49 (.ZN( u1_u6_u0_n171 ) , .A( u1_u6_u0_n99 ) );
  AOI21_X1 u1_u6_u0_U5 (.B2( u1_u6_u0_n131 ) , .ZN( u1_u6_u0_n134 ) , .B1( u1_u6_u0_n151 ) , .A( u1_u6_u0_n158 ) );
  OAI211_X1 u1_u6_u0_U50 (.C2( u1_u6_u0_n140 ) , .C1( u1_u6_u0_n161 ) , .A( u1_u6_u0_n169 ) , .B( u1_u6_u0_n98 ) , .ZN( u1_u6_u0_n99 ) );
  INV_X1 u1_u6_u0_U51 (.ZN( u1_u6_u0_n169 ) , .A( u1_u6_u0_n91 ) );
  AOI211_X1 u1_u6_u0_U52 (.C1( u1_u6_u0_n118 ) , .A( u1_u6_u0_n123 ) , .B( u1_u6_u0_n96 ) , .C2( u1_u6_u0_n97 ) , .ZN( u1_u6_u0_n98 ) );
  NOR2_X1 u1_u6_u0_U53 (.A2( u1_u6_X_4 ) , .A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n118 ) );
  NOR2_X1 u1_u6_u0_U54 (.A2( u1_u6_X_2 ) , .ZN( u1_u6_u0_n103 ) , .A1( u1_u6_u0_n164 ) );
  NOR2_X1 u1_u6_u0_U55 (.A2( u1_u6_X_1 ) , .A1( u1_u6_X_2 ) , .ZN( u1_u6_u0_n92 ) );
  NOR2_X1 u1_u6_u0_U56 (.A2( u1_u6_X_1 ) , .ZN( u1_u6_u0_n101 ) , .A1( u1_u6_u0_n163 ) );
  NAND2_X1 u1_u6_u0_U57 (.A2( u1_u6_X_4 ) , .A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n144 ) );
  NOR2_X1 u1_u6_u0_U58 (.A2( u1_u6_X_5 ) , .ZN( u1_u6_u0_n136 ) , .A1( u1_u6_u0_n159 ) );
  NAND2_X1 u1_u6_u0_U59 (.A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n138 ) , .A2( u1_u6_u0_n159 ) );
  NOR2_X1 u1_u6_u0_U6 (.A1( u1_u6_u0_n108 ) , .ZN( u1_u6_u0_n123 ) , .A2( u1_u6_u0_n158 ) );
  AND2_X1 u1_u6_u0_U60 (.A2( u1_u6_X_3 ) , .A1( u1_u6_X_6 ) , .ZN( u1_u6_u0_n102 ) );
  INV_X1 u1_u6_u0_U61 (.A( u1_u6_X_4 ) , .ZN( u1_u6_u0_n159 ) );
  INV_X1 u1_u6_u0_U62 (.A( u1_u6_X_1 ) , .ZN( u1_u6_u0_n164 ) );
  INV_X1 u1_u6_u0_U63 (.A( u1_u6_X_2 ) , .ZN( u1_u6_u0_n163 ) );
  INV_X1 u1_u6_u0_U64 (.A( u1_u6_X_3 ) , .ZN( u1_u6_u0_n162 ) );
  INV_X1 u1_u6_u0_U65 (.A( u1_u6_u0_n126 ) , .ZN( u1_u6_u0_n168 ) );
  AOI211_X1 u1_u6_u0_U66 (.B( u1_u6_u0_n133 ) , .A( u1_u6_u0_n134 ) , .C2( u1_u6_u0_n135 ) , .C1( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n137 ) );
  OR4_X1 u1_u6_u0_U67 (.ZN( u1_out6_17 ) , .A4( u1_u6_u0_n122 ) , .A2( u1_u6_u0_n123 ) , .A1( u1_u6_u0_n124 ) , .A3( u1_u6_u0_n170 ) );
  AOI21_X1 u1_u6_u0_U68 (.B2( u1_u6_u0_n107 ) , .ZN( u1_u6_u0_n124 ) , .B1( u1_u6_u0_n128 ) , .A( u1_u6_u0_n161 ) );
  INV_X1 u1_u6_u0_U69 (.A( u1_u6_u0_n111 ) , .ZN( u1_u6_u0_n170 ) );
  OAI21_X1 u1_u6_u0_U7 (.B1( u1_u6_u0_n150 ) , .B2( u1_u6_u0_n158 ) , .A( u1_u6_u0_n172 ) , .ZN( u1_u6_u0_n89 ) );
  OR4_X1 u1_u6_u0_U70 (.ZN( u1_out6_31 ) , .A4( u1_u6_u0_n155 ) , .A2( u1_u6_u0_n156 ) , .A1( u1_u6_u0_n157 ) , .A3( u1_u6_u0_n173 ) );
  AOI21_X1 u1_u6_u0_U71 (.A( u1_u6_u0_n138 ) , .B2( u1_u6_u0_n139 ) , .B1( u1_u6_u0_n140 ) , .ZN( u1_u6_u0_n157 ) );
  AOI21_X1 u1_u6_u0_U72 (.B2( u1_u6_u0_n141 ) , .B1( u1_u6_u0_n142 ) , .ZN( u1_u6_u0_n156 ) , .A( u1_u6_u0_n161 ) );
  INV_X1 u1_u6_u0_U73 (.ZN( u1_u6_u0_n174 ) , .A( u1_u6_u0_n89 ) );
  AOI211_X1 u1_u6_u0_U74 (.B( u1_u6_u0_n104 ) , .A( u1_u6_u0_n105 ) , .ZN( u1_u6_u0_n106 ) , .C2( u1_u6_u0_n113 ) , .C1( u1_u6_u0_n160 ) );
  OAI221_X1 u1_u6_u0_U75 (.C1( u1_u6_u0_n121 ) , .ZN( u1_u6_u0_n122 ) , .B2( u1_u6_u0_n127 ) , .A( u1_u6_u0_n143 ) , .B1( u1_u6_u0_n144 ) , .C2( u1_u6_u0_n147 ) );
  NOR2_X1 u1_u6_u0_U76 (.A1( u1_u6_u0_n120 ) , .ZN( u1_u6_u0_n143 ) , .A2( u1_u6_u0_n167 ) );
  AOI21_X1 u1_u6_u0_U77 (.B1( u1_u6_u0_n132 ) , .ZN( u1_u6_u0_n133 ) , .A( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n166 ) );
  OAI22_X1 u1_u6_u0_U78 (.ZN( u1_u6_u0_n105 ) , .A2( u1_u6_u0_n132 ) , .B1( u1_u6_u0_n146 ) , .A1( u1_u6_u0_n147 ) , .B2( u1_u6_u0_n161 ) );
  NAND2_X1 u1_u6_u0_U79 (.ZN( u1_u6_u0_n110 ) , .A2( u1_u6_u0_n132 ) , .A1( u1_u6_u0_n145 ) );
  AND2_X1 u1_u6_u0_U8 (.A1( u1_u6_u0_n114 ) , .A2( u1_u6_u0_n121 ) , .ZN( u1_u6_u0_n146 ) );
  INV_X1 u1_u6_u0_U80 (.A( u1_u6_u0_n119 ) , .ZN( u1_u6_u0_n167 ) );
  NAND2_X1 u1_u6_u0_U81 (.A2( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n140 ) , .A1( u1_u6_u0_n94 ) );
  NAND2_X1 u1_u6_u0_U82 (.A1( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n130 ) , .A2( u1_u6_u0_n94 ) );
  NAND2_X1 u1_u6_u0_U83 (.ZN( u1_u6_u0_n108 ) , .A1( u1_u6_u0_n92 ) , .A2( u1_u6_u0_n94 ) );
  AND2_X1 u1_u6_u0_U84 (.A1( u1_u6_X_6 ) , .A2( u1_u6_u0_n162 ) , .ZN( u1_u6_u0_n93 ) );
  NAND2_X1 u1_u6_u0_U85 (.ZN( u1_u6_u0_n142 ) , .A1( u1_u6_u0_n94 ) , .A2( u1_u6_u0_n95 ) );
  NOR2_X1 u1_u6_u0_U86 (.A2( u1_u6_X_6 ) , .ZN( u1_u6_u0_n100 ) , .A1( u1_u6_u0_n162 ) );
  NOR2_X1 u1_u6_u0_U87 (.A2( u1_u6_X_3 ) , .A1( u1_u6_X_6 ) , .ZN( u1_u6_u0_n94 ) );
  NAND3_X1 u1_u6_u0_U88 (.ZN( u1_out6_23 ) , .A3( u1_u6_u0_n137 ) , .A1( u1_u6_u0_n168 ) , .A2( u1_u6_u0_n171 ) );
  NAND3_X1 u1_u6_u0_U89 (.A3( u1_u6_u0_n127 ) , .A2( u1_u6_u0_n128 ) , .ZN( u1_u6_u0_n135 ) , .A1( u1_u6_u0_n150 ) );
  AND2_X1 u1_u6_u0_U9 (.A1( u1_u6_u0_n131 ) , .ZN( u1_u6_u0_n141 ) , .A2( u1_u6_u0_n150 ) );
  NAND3_X1 u1_u6_u0_U90 (.ZN( u1_u6_u0_n117 ) , .A3( u1_u6_u0_n132 ) , .A2( u1_u6_u0_n139 ) , .A1( u1_u6_u0_n148 ) );
  NAND3_X1 u1_u6_u0_U91 (.ZN( u1_u6_u0_n109 ) , .A2( u1_u6_u0_n114 ) , .A3( u1_u6_u0_n140 ) , .A1( u1_u6_u0_n149 ) );
  NAND3_X1 u1_u6_u0_U92 (.ZN( u1_out6_9 ) , .A3( u1_u6_u0_n106 ) , .A2( u1_u6_u0_n171 ) , .A1( u1_u6_u0_n174 ) );
  NAND3_X1 u1_u6_u0_U93 (.A2( u1_u6_u0_n128 ) , .A1( u1_u6_u0_n132 ) , .A3( u1_u6_u0_n146 ) , .ZN( u1_u6_u0_n97 ) );
  OAI22_X1 u1_u6_u4_U10 (.B2( u1_u6_u4_n135 ) , .ZN( u1_u6_u4_n137 ) , .B1( u1_u6_u4_n153 ) , .A1( u1_u6_u4_n155 ) , .A2( u1_u6_u4_n171 ) );
  AND3_X1 u1_u6_u4_U11 (.A2( u1_u6_u4_n134 ) , .ZN( u1_u6_u4_n135 ) , .A3( u1_u6_u4_n145 ) , .A1( u1_u6_u4_n157 ) );
  NAND2_X1 u1_u6_u4_U12 (.ZN( u1_u6_u4_n132 ) , .A2( u1_u6_u4_n170 ) , .A1( u1_u6_u4_n173 ) );
  AOI21_X1 u1_u6_u4_U13 (.B2( u1_u6_u4_n160 ) , .B1( u1_u6_u4_n161 ) , .ZN( u1_u6_u4_n162 ) , .A( u1_u6_u4_n170 ) );
  AOI21_X1 u1_u6_u4_U14 (.ZN( u1_u6_u4_n107 ) , .B2( u1_u6_u4_n143 ) , .A( u1_u6_u4_n174 ) , .B1( u1_u6_u4_n184 ) );
  AOI21_X1 u1_u6_u4_U15 (.B2( u1_u6_u4_n158 ) , .B1( u1_u6_u4_n159 ) , .ZN( u1_u6_u4_n163 ) , .A( u1_u6_u4_n174 ) );
  AOI21_X1 u1_u6_u4_U16 (.A( u1_u6_u4_n153 ) , .B2( u1_u6_u4_n154 ) , .B1( u1_u6_u4_n155 ) , .ZN( u1_u6_u4_n165 ) );
  AOI21_X1 u1_u6_u4_U17 (.A( u1_u6_u4_n156 ) , .B2( u1_u6_u4_n157 ) , .ZN( u1_u6_u4_n164 ) , .B1( u1_u6_u4_n184 ) );
  INV_X1 u1_u6_u4_U18 (.A( u1_u6_u4_n138 ) , .ZN( u1_u6_u4_n170 ) );
  AND2_X1 u1_u6_u4_U19 (.A2( u1_u6_u4_n120 ) , .ZN( u1_u6_u4_n155 ) , .A1( u1_u6_u4_n160 ) );
  INV_X1 u1_u6_u4_U20 (.A( u1_u6_u4_n156 ) , .ZN( u1_u6_u4_n175 ) );
  NAND2_X1 u1_u6_u4_U21 (.A2( u1_u6_u4_n118 ) , .ZN( u1_u6_u4_n131 ) , .A1( u1_u6_u4_n147 ) );
  NAND2_X1 u1_u6_u4_U22 (.A1( u1_u6_u4_n119 ) , .A2( u1_u6_u4_n120 ) , .ZN( u1_u6_u4_n130 ) );
  NAND2_X1 u1_u6_u4_U23 (.ZN( u1_u6_u4_n117 ) , .A2( u1_u6_u4_n118 ) , .A1( u1_u6_u4_n148 ) );
  NAND2_X1 u1_u6_u4_U24 (.ZN( u1_u6_u4_n129 ) , .A1( u1_u6_u4_n134 ) , .A2( u1_u6_u4_n148 ) );
  AND3_X1 u1_u6_u4_U25 (.A1( u1_u6_u4_n119 ) , .A2( u1_u6_u4_n143 ) , .A3( u1_u6_u4_n154 ) , .ZN( u1_u6_u4_n161 ) );
  AND2_X1 u1_u6_u4_U26 (.A1( u1_u6_u4_n145 ) , .A2( u1_u6_u4_n147 ) , .ZN( u1_u6_u4_n159 ) );
  OR3_X1 u1_u6_u4_U27 (.A3( u1_u6_u4_n114 ) , .A2( u1_u6_u4_n115 ) , .A1( u1_u6_u4_n116 ) , .ZN( u1_u6_u4_n136 ) );
  AOI21_X1 u1_u6_u4_U28 (.A( u1_u6_u4_n113 ) , .ZN( u1_u6_u4_n116 ) , .B2( u1_u6_u4_n173 ) , .B1( u1_u6_u4_n174 ) );
  AOI21_X1 u1_u6_u4_U29 (.ZN( u1_u6_u4_n115 ) , .B2( u1_u6_u4_n145 ) , .B1( u1_u6_u4_n146 ) , .A( u1_u6_u4_n156 ) );
  NOR2_X1 u1_u6_u4_U3 (.ZN( u1_u6_u4_n121 ) , .A1( u1_u6_u4_n181 ) , .A2( u1_u6_u4_n182 ) );
  OAI22_X1 u1_u6_u4_U30 (.ZN( u1_u6_u4_n114 ) , .A2( u1_u6_u4_n121 ) , .B1( u1_u6_u4_n160 ) , .B2( u1_u6_u4_n170 ) , .A1( u1_u6_u4_n171 ) );
  INV_X1 u1_u6_u4_U31 (.A( u1_u6_u4_n158 ) , .ZN( u1_u6_u4_n182 ) );
  INV_X1 u1_u6_u4_U32 (.ZN( u1_u6_u4_n181 ) , .A( u1_u6_u4_n96 ) );
  INV_X1 u1_u6_u4_U33 (.A( u1_u6_u4_n144 ) , .ZN( u1_u6_u4_n179 ) );
  INV_X1 u1_u6_u4_U34 (.A( u1_u6_u4_n157 ) , .ZN( u1_u6_u4_n178 ) );
  NAND2_X1 u1_u6_u4_U35 (.A2( u1_u6_u4_n154 ) , .A1( u1_u6_u4_n96 ) , .ZN( u1_u6_u4_n97 ) );
  INV_X1 u1_u6_u4_U36 (.ZN( u1_u6_u4_n186 ) , .A( u1_u6_u4_n95 ) );
  OAI221_X1 u1_u6_u4_U37 (.C1( u1_u6_u4_n134 ) , .B1( u1_u6_u4_n158 ) , .B2( u1_u6_u4_n171 ) , .C2( u1_u6_u4_n173 ) , .A( u1_u6_u4_n94 ) , .ZN( u1_u6_u4_n95 ) );
  AOI222_X1 u1_u6_u4_U38 (.B2( u1_u6_u4_n132 ) , .A1( u1_u6_u4_n138 ) , .C2( u1_u6_u4_n175 ) , .A2( u1_u6_u4_n179 ) , .C1( u1_u6_u4_n181 ) , .B1( u1_u6_u4_n185 ) , .ZN( u1_u6_u4_n94 ) );
  INV_X1 u1_u6_u4_U39 (.A( u1_u6_u4_n113 ) , .ZN( u1_u6_u4_n185 ) );
  INV_X1 u1_u6_u4_U4 (.A( u1_u6_u4_n117 ) , .ZN( u1_u6_u4_n184 ) );
  INV_X1 u1_u6_u4_U40 (.A( u1_u6_u4_n143 ) , .ZN( u1_u6_u4_n183 ) );
  NOR2_X1 u1_u6_u4_U41 (.ZN( u1_u6_u4_n138 ) , .A1( u1_u6_u4_n168 ) , .A2( u1_u6_u4_n169 ) );
  NOR2_X1 u1_u6_u4_U42 (.A1( u1_u6_u4_n150 ) , .A2( u1_u6_u4_n152 ) , .ZN( u1_u6_u4_n153 ) );
  NOR2_X1 u1_u6_u4_U43 (.A2( u1_u6_u4_n128 ) , .A1( u1_u6_u4_n138 ) , .ZN( u1_u6_u4_n156 ) );
  AOI22_X1 u1_u6_u4_U44 (.B2( u1_u6_u4_n122 ) , .A1( u1_u6_u4_n123 ) , .ZN( u1_u6_u4_n124 ) , .B1( u1_u6_u4_n128 ) , .A2( u1_u6_u4_n172 ) );
  INV_X1 u1_u6_u4_U45 (.A( u1_u6_u4_n153 ) , .ZN( u1_u6_u4_n172 ) );
  NAND2_X1 u1_u6_u4_U46 (.A2( u1_u6_u4_n120 ) , .ZN( u1_u6_u4_n123 ) , .A1( u1_u6_u4_n161 ) );
  AOI22_X1 u1_u6_u4_U47 (.B2( u1_u6_u4_n132 ) , .A2( u1_u6_u4_n133 ) , .ZN( u1_u6_u4_n140 ) , .A1( u1_u6_u4_n150 ) , .B1( u1_u6_u4_n179 ) );
  NAND2_X1 u1_u6_u4_U48 (.ZN( u1_u6_u4_n133 ) , .A2( u1_u6_u4_n146 ) , .A1( u1_u6_u4_n154 ) );
  NAND2_X1 u1_u6_u4_U49 (.A1( u1_u6_u4_n103 ) , .ZN( u1_u6_u4_n154 ) , .A2( u1_u6_u4_n98 ) );
  NOR4_X1 u1_u6_u4_U5 (.A4( u1_u6_u4_n106 ) , .A3( u1_u6_u4_n107 ) , .A2( u1_u6_u4_n108 ) , .A1( u1_u6_u4_n109 ) , .ZN( u1_u6_u4_n110 ) );
  NAND2_X1 u1_u6_u4_U50 (.A1( u1_u6_u4_n101 ) , .ZN( u1_u6_u4_n158 ) , .A2( u1_u6_u4_n99 ) );
  AOI21_X1 u1_u6_u4_U51 (.ZN( u1_u6_u4_n127 ) , .A( u1_u6_u4_n136 ) , .B2( u1_u6_u4_n150 ) , .B1( u1_u6_u4_n180 ) );
  INV_X1 u1_u6_u4_U52 (.A( u1_u6_u4_n160 ) , .ZN( u1_u6_u4_n180 ) );
  NAND2_X1 u1_u6_u4_U53 (.A2( u1_u6_u4_n104 ) , .A1( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n146 ) );
  NAND2_X1 u1_u6_u4_U54 (.A2( u1_u6_u4_n101 ) , .A1( u1_u6_u4_n102 ) , .ZN( u1_u6_u4_n160 ) );
  NAND2_X1 u1_u6_u4_U55 (.ZN( u1_u6_u4_n134 ) , .A1( u1_u6_u4_n98 ) , .A2( u1_u6_u4_n99 ) );
  NAND2_X1 u1_u6_u4_U56 (.A1( u1_u6_u4_n103 ) , .A2( u1_u6_u4_n104 ) , .ZN( u1_u6_u4_n143 ) );
  NAND2_X1 u1_u6_u4_U57 (.A2( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n145 ) , .A1( u1_u6_u4_n98 ) );
  NAND2_X1 u1_u6_u4_U58 (.A1( u1_u6_u4_n100 ) , .A2( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n120 ) );
  NAND2_X1 u1_u6_u4_U59 (.A1( u1_u6_u4_n102 ) , .A2( u1_u6_u4_n104 ) , .ZN( u1_u6_u4_n148 ) );
  AOI21_X1 u1_u6_u4_U6 (.ZN( u1_u6_u4_n106 ) , .B2( u1_u6_u4_n146 ) , .B1( u1_u6_u4_n158 ) , .A( u1_u6_u4_n170 ) );
  NAND2_X1 u1_u6_u4_U60 (.A2( u1_u6_u4_n100 ) , .A1( u1_u6_u4_n103 ) , .ZN( u1_u6_u4_n157 ) );
  INV_X1 u1_u6_u4_U61 (.A( u1_u6_u4_n150 ) , .ZN( u1_u6_u4_n173 ) );
  INV_X1 u1_u6_u4_U62 (.A( u1_u6_u4_n152 ) , .ZN( u1_u6_u4_n171 ) );
  NAND2_X1 u1_u6_u4_U63 (.A1( u1_u6_u4_n100 ) , .ZN( u1_u6_u4_n118 ) , .A2( u1_u6_u4_n99 ) );
  NAND2_X1 u1_u6_u4_U64 (.A2( u1_u6_u4_n100 ) , .A1( u1_u6_u4_n102 ) , .ZN( u1_u6_u4_n144 ) );
  NAND2_X1 u1_u6_u4_U65 (.A2( u1_u6_u4_n101 ) , .A1( u1_u6_u4_n105 ) , .ZN( u1_u6_u4_n96 ) );
  INV_X1 u1_u6_u4_U66 (.A( u1_u6_u4_n128 ) , .ZN( u1_u6_u4_n174 ) );
  NAND2_X1 u1_u6_u4_U67 (.A2( u1_u6_u4_n102 ) , .ZN( u1_u6_u4_n119 ) , .A1( u1_u6_u4_n98 ) );
  NAND2_X1 u1_u6_u4_U68 (.A2( u1_u6_u4_n101 ) , .A1( u1_u6_u4_n103 ) , .ZN( u1_u6_u4_n147 ) );
  NAND2_X1 u1_u6_u4_U69 (.A2( u1_u6_u4_n104 ) , .ZN( u1_u6_u4_n113 ) , .A1( u1_u6_u4_n99 ) );
  AOI21_X1 u1_u6_u4_U7 (.ZN( u1_u6_u4_n108 ) , .B2( u1_u6_u4_n134 ) , .B1( u1_u6_u4_n155 ) , .A( u1_u6_u4_n156 ) );
  NOR2_X1 u1_u6_u4_U70 (.A2( u1_u6_X_28 ) , .ZN( u1_u6_u4_n150 ) , .A1( u1_u6_u4_n168 ) );
  NOR2_X1 u1_u6_u4_U71 (.A2( u1_u6_X_29 ) , .ZN( u1_u6_u4_n152 ) , .A1( u1_u6_u4_n169 ) );
  NOR2_X1 u1_u6_u4_U72 (.A2( u1_u6_X_30 ) , .ZN( u1_u6_u4_n105 ) , .A1( u1_u6_u4_n176 ) );
  NOR2_X1 u1_u6_u4_U73 (.A2( u1_u6_X_26 ) , .ZN( u1_u6_u4_n100 ) , .A1( u1_u6_u4_n177 ) );
  NOR2_X1 u1_u6_u4_U74 (.A2( u1_u6_X_28 ) , .A1( u1_u6_X_29 ) , .ZN( u1_u6_u4_n128 ) );
  NOR2_X1 u1_u6_u4_U75 (.A2( u1_u6_X_27 ) , .A1( u1_u6_X_30 ) , .ZN( u1_u6_u4_n102 ) );
  NOR2_X1 u1_u6_u4_U76 (.A2( u1_u6_X_25 ) , .A1( u1_u6_X_26 ) , .ZN( u1_u6_u4_n98 ) );
  AND2_X1 u1_u6_u4_U77 (.A2( u1_u6_X_25 ) , .A1( u1_u6_X_26 ) , .ZN( u1_u6_u4_n104 ) );
  AND2_X1 u1_u6_u4_U78 (.A1( u1_u6_X_30 ) , .A2( u1_u6_u4_n176 ) , .ZN( u1_u6_u4_n99 ) );
  AND2_X1 u1_u6_u4_U79 (.A1( u1_u6_X_26 ) , .ZN( u1_u6_u4_n101 ) , .A2( u1_u6_u4_n177 ) );
  AOI21_X1 u1_u6_u4_U8 (.ZN( u1_u6_u4_n109 ) , .A( u1_u6_u4_n153 ) , .B1( u1_u6_u4_n159 ) , .B2( u1_u6_u4_n184 ) );
  AND2_X1 u1_u6_u4_U80 (.A1( u1_u6_X_27 ) , .A2( u1_u6_X_30 ) , .ZN( u1_u6_u4_n103 ) );
  INV_X1 u1_u6_u4_U81 (.A( u1_u6_X_28 ) , .ZN( u1_u6_u4_n169 ) );
  INV_X1 u1_u6_u4_U82 (.A( u1_u6_X_29 ) , .ZN( u1_u6_u4_n168 ) );
  INV_X1 u1_u6_u4_U83 (.A( u1_u6_X_25 ) , .ZN( u1_u6_u4_n177 ) );
  INV_X1 u1_u6_u4_U84 (.A( u1_u6_X_27 ) , .ZN( u1_u6_u4_n176 ) );
  NAND4_X1 u1_u6_u4_U85 (.ZN( u1_out6_8 ) , .A4( u1_u6_u4_n110 ) , .A3( u1_u6_u4_n111 ) , .A2( u1_u6_u4_n112 ) , .A1( u1_u6_u4_n186 ) );
  NAND2_X1 u1_u6_u4_U86 (.ZN( u1_u6_u4_n112 ) , .A2( u1_u6_u4_n130 ) , .A1( u1_u6_u4_n150 ) );
  AOI22_X1 u1_u6_u4_U87 (.ZN( u1_u6_u4_n111 ) , .B2( u1_u6_u4_n132 ) , .A1( u1_u6_u4_n152 ) , .B1( u1_u6_u4_n178 ) , .A2( u1_u6_u4_n97 ) );
  NAND4_X1 u1_u6_u4_U88 (.ZN( u1_out6_25 ) , .A4( u1_u6_u4_n139 ) , .A3( u1_u6_u4_n140 ) , .A2( u1_u6_u4_n141 ) , .A1( u1_u6_u4_n142 ) );
  OAI21_X1 u1_u6_u4_U89 (.B2( u1_u6_u4_n131 ) , .ZN( u1_u6_u4_n141 ) , .A( u1_u6_u4_n175 ) , .B1( u1_u6_u4_n183 ) );
  AOI211_X1 u1_u6_u4_U9 (.B( u1_u6_u4_n136 ) , .A( u1_u6_u4_n137 ) , .C2( u1_u6_u4_n138 ) , .ZN( u1_u6_u4_n139 ) , .C1( u1_u6_u4_n182 ) );
  OAI21_X1 u1_u6_u4_U90 (.A( u1_u6_u4_n128 ) , .B2( u1_u6_u4_n129 ) , .B1( u1_u6_u4_n130 ) , .ZN( u1_u6_u4_n142 ) );
  NAND4_X1 u1_u6_u4_U91 (.ZN( u1_out6_14 ) , .A4( u1_u6_u4_n124 ) , .A3( u1_u6_u4_n125 ) , .A2( u1_u6_u4_n126 ) , .A1( u1_u6_u4_n127 ) );
  AOI22_X1 u1_u6_u4_U92 (.B2( u1_u6_u4_n117 ) , .ZN( u1_u6_u4_n126 ) , .A1( u1_u6_u4_n129 ) , .B1( u1_u6_u4_n152 ) , .A2( u1_u6_u4_n175 ) );
  AOI22_X1 u1_u6_u4_U93 (.ZN( u1_u6_u4_n125 ) , .B2( u1_u6_u4_n131 ) , .A2( u1_u6_u4_n132 ) , .B1( u1_u6_u4_n138 ) , .A1( u1_u6_u4_n178 ) );
  AOI22_X1 u1_u6_u4_U94 (.B2( u1_u6_u4_n149 ) , .B1( u1_u6_u4_n150 ) , .A2( u1_u6_u4_n151 ) , .A1( u1_u6_u4_n152 ) , .ZN( u1_u6_u4_n167 ) );
  NOR4_X1 u1_u6_u4_U95 (.A4( u1_u6_u4_n162 ) , .A3( u1_u6_u4_n163 ) , .A2( u1_u6_u4_n164 ) , .A1( u1_u6_u4_n165 ) , .ZN( u1_u6_u4_n166 ) );
  NAND3_X1 u1_u6_u4_U96 (.ZN( u1_out6_3 ) , .A3( u1_u6_u4_n166 ) , .A1( u1_u6_u4_n167 ) , .A2( u1_u6_u4_n186 ) );
  NAND3_X1 u1_u6_u4_U97 (.A3( u1_u6_u4_n146 ) , .A2( u1_u6_u4_n147 ) , .A1( u1_u6_u4_n148 ) , .ZN( u1_u6_u4_n149 ) );
  NAND3_X1 u1_u6_u4_U98 (.A3( u1_u6_u4_n143 ) , .A2( u1_u6_u4_n144 ) , .A1( u1_u6_u4_n145 ) , .ZN( u1_u6_u4_n151 ) );
  NAND3_X1 u1_u6_u4_U99 (.A3( u1_u6_u4_n121 ) , .ZN( u1_u6_u4_n122 ) , .A2( u1_u6_u4_n144 ) , .A1( u1_u6_u4_n154 ) );
  AOI21_X1 u1_u6_u6_U10 (.ZN( u1_u6_u6_n106 ) , .A( u1_u6_u6_n142 ) , .B2( u1_u6_u6_n159 ) , .B1( u1_u6_u6_n164 ) );
  INV_X1 u1_u6_u6_U11 (.A( u1_u6_u6_n155 ) , .ZN( u1_u6_u6_n161 ) );
  INV_X1 u1_u6_u6_U12 (.A( u1_u6_u6_n128 ) , .ZN( u1_u6_u6_n164 ) );
  NAND2_X1 u1_u6_u6_U13 (.ZN( u1_u6_u6_n110 ) , .A1( u1_u6_u6_n122 ) , .A2( u1_u6_u6_n129 ) );
  NAND2_X1 u1_u6_u6_U14 (.ZN( u1_u6_u6_n124 ) , .A2( u1_u6_u6_n146 ) , .A1( u1_u6_u6_n148 ) );
  INV_X1 u1_u6_u6_U15 (.A( u1_u6_u6_n132 ) , .ZN( u1_u6_u6_n171 ) );
  AND2_X1 u1_u6_u6_U16 (.A1( u1_u6_u6_n100 ) , .ZN( u1_u6_u6_n130 ) , .A2( u1_u6_u6_n147 ) );
  INV_X1 u1_u6_u6_U17 (.A( u1_u6_u6_n127 ) , .ZN( u1_u6_u6_n173 ) );
  INV_X1 u1_u6_u6_U18 (.A( u1_u6_u6_n121 ) , .ZN( u1_u6_u6_n167 ) );
  INV_X1 u1_u6_u6_U19 (.A( u1_u6_u6_n100 ) , .ZN( u1_u6_u6_n169 ) );
  INV_X1 u1_u6_u6_U20 (.A( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n170 ) );
  INV_X1 u1_u6_u6_U21 (.A( u1_u6_u6_n113 ) , .ZN( u1_u6_u6_n168 ) );
  AND2_X1 u1_u6_u6_U22 (.A1( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n119 ) , .ZN( u1_u6_u6_n133 ) );
  AND2_X1 u1_u6_u6_U23 (.A2( u1_u6_u6_n121 ) , .A1( u1_u6_u6_n122 ) , .ZN( u1_u6_u6_n131 ) );
  AND3_X1 u1_u6_u6_U24 (.ZN( u1_u6_u6_n120 ) , .A2( u1_u6_u6_n127 ) , .A1( u1_u6_u6_n132 ) , .A3( u1_u6_u6_n145 ) );
  INV_X1 u1_u6_u6_U25 (.A( u1_u6_u6_n146 ) , .ZN( u1_u6_u6_n163 ) );
  AOI222_X1 u1_u6_u6_U26 (.ZN( u1_u6_u6_n114 ) , .A1( u1_u6_u6_n118 ) , .A2( u1_u6_u6_n126 ) , .B2( u1_u6_u6_n151 ) , .C2( u1_u6_u6_n159 ) , .C1( u1_u6_u6_n168 ) , .B1( u1_u6_u6_n169 ) );
  NOR2_X1 u1_u6_u6_U27 (.A1( u1_u6_u6_n162 ) , .A2( u1_u6_u6_n165 ) , .ZN( u1_u6_u6_n98 ) );
  AOI211_X1 u1_u6_u6_U28 (.B( u1_u6_u6_n149 ) , .A( u1_u6_u6_n150 ) , .C2( u1_u6_u6_n151 ) , .C1( u1_u6_u6_n152 ) , .ZN( u1_u6_u6_n153 ) );
  AOI21_X1 u1_u6_u6_U29 (.B2( u1_u6_u6_n147 ) , .B1( u1_u6_u6_n148 ) , .ZN( u1_u6_u6_n149 ) , .A( u1_u6_u6_n158 ) );
  INV_X1 u1_u6_u6_U3 (.A( u1_u6_u6_n110 ) , .ZN( u1_u6_u6_n166 ) );
  AOI21_X1 u1_u6_u6_U30 (.A( u1_u6_u6_n144 ) , .B2( u1_u6_u6_n145 ) , .B1( u1_u6_u6_n146 ) , .ZN( u1_u6_u6_n150 ) );
  NAND2_X1 u1_u6_u6_U31 (.A2( u1_u6_u6_n143 ) , .ZN( u1_u6_u6_n152 ) , .A1( u1_u6_u6_n166 ) );
  NAND2_X1 u1_u6_u6_U32 (.A1( u1_u6_u6_n144 ) , .ZN( u1_u6_u6_n151 ) , .A2( u1_u6_u6_n158 ) );
  NAND2_X1 u1_u6_u6_U33 (.ZN( u1_u6_u6_n132 ) , .A1( u1_u6_u6_n91 ) , .A2( u1_u6_u6_n97 ) );
  AOI22_X1 u1_u6_u6_U34 (.B2( u1_u6_u6_n110 ) , .B1( u1_u6_u6_n111 ) , .A1( u1_u6_u6_n112 ) , .ZN( u1_u6_u6_n115 ) , .A2( u1_u6_u6_n161 ) );
  NAND4_X1 u1_u6_u6_U35 (.A3( u1_u6_u6_n109 ) , .ZN( u1_u6_u6_n112 ) , .A4( u1_u6_u6_n132 ) , .A2( u1_u6_u6_n147 ) , .A1( u1_u6_u6_n166 ) );
  NOR2_X1 u1_u6_u6_U36 (.ZN( u1_u6_u6_n109 ) , .A1( u1_u6_u6_n170 ) , .A2( u1_u6_u6_n173 ) );
  NOR2_X1 u1_u6_u6_U37 (.A2( u1_u6_u6_n126 ) , .ZN( u1_u6_u6_n155 ) , .A1( u1_u6_u6_n160 ) );
  NAND2_X1 u1_u6_u6_U38 (.ZN( u1_u6_u6_n146 ) , .A2( u1_u6_u6_n94 ) , .A1( u1_u6_u6_n99 ) );
  AOI211_X1 u1_u6_u6_U39 (.B( u1_u6_u6_n134 ) , .A( u1_u6_u6_n135 ) , .C1( u1_u6_u6_n136 ) , .ZN( u1_u6_u6_n137 ) , .C2( u1_u6_u6_n151 ) );
  AOI22_X1 u1_u6_u6_U4 (.B2( u1_u6_u6_n101 ) , .A1( u1_u6_u6_n102 ) , .ZN( u1_u6_u6_n103 ) , .B1( u1_u6_u6_n160 ) , .A2( u1_u6_u6_n161 ) );
  NAND4_X1 u1_u6_u6_U40 (.A4( u1_u6_u6_n127 ) , .A3( u1_u6_u6_n128 ) , .A2( u1_u6_u6_n129 ) , .A1( u1_u6_u6_n130 ) , .ZN( u1_u6_u6_n136 ) );
  AOI21_X1 u1_u6_u6_U41 (.B2( u1_u6_u6_n132 ) , .B1( u1_u6_u6_n133 ) , .ZN( u1_u6_u6_n134 ) , .A( u1_u6_u6_n158 ) );
  AOI21_X1 u1_u6_u6_U42 (.B1( u1_u6_u6_n131 ) , .ZN( u1_u6_u6_n135 ) , .A( u1_u6_u6_n144 ) , .B2( u1_u6_u6_n146 ) );
  INV_X1 u1_u6_u6_U43 (.A( u1_u6_u6_n111 ) , .ZN( u1_u6_u6_n158 ) );
  NAND2_X1 u1_u6_u6_U44 (.ZN( u1_u6_u6_n127 ) , .A1( u1_u6_u6_n91 ) , .A2( u1_u6_u6_n92 ) );
  NAND2_X1 u1_u6_u6_U45 (.ZN( u1_u6_u6_n129 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n96 ) );
  INV_X1 u1_u6_u6_U46 (.A( u1_u6_u6_n144 ) , .ZN( u1_u6_u6_n159 ) );
  NAND2_X1 u1_u6_u6_U47 (.ZN( u1_u6_u6_n145 ) , .A2( u1_u6_u6_n97 ) , .A1( u1_u6_u6_n98 ) );
  NAND2_X1 u1_u6_u6_U48 (.ZN( u1_u6_u6_n148 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n94 ) );
  NAND2_X1 u1_u6_u6_U49 (.ZN( u1_u6_u6_n108 ) , .A2( u1_u6_u6_n139 ) , .A1( u1_u6_u6_n144 ) );
  NOR2_X1 u1_u6_u6_U5 (.A1( u1_u6_u6_n118 ) , .ZN( u1_u6_u6_n143 ) , .A2( u1_u6_u6_n168 ) );
  NAND2_X1 u1_u6_u6_U50 (.ZN( u1_u6_u6_n121 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n97 ) );
  NAND2_X1 u1_u6_u6_U51 (.ZN( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n95 ) );
  AND2_X1 u1_u6_u6_U52 (.ZN( u1_u6_u6_n118 ) , .A2( u1_u6_u6_n91 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U53 (.ZN( u1_u6_u6_n147 ) , .A2( u1_u6_u6_n98 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U54 (.ZN( u1_u6_u6_n128 ) , .A1( u1_u6_u6_n94 ) , .A2( u1_u6_u6_n96 ) );
  NAND2_X1 u1_u6_u6_U55 (.ZN( u1_u6_u6_n119 ) , .A2( u1_u6_u6_n95 ) , .A1( u1_u6_u6_n99 ) );
  NAND2_X1 u1_u6_u6_U56 (.ZN( u1_u6_u6_n123 ) , .A2( u1_u6_u6_n91 ) , .A1( u1_u6_u6_n96 ) );
  NAND2_X1 u1_u6_u6_U57 (.ZN( u1_u6_u6_n100 ) , .A2( u1_u6_u6_n92 ) , .A1( u1_u6_u6_n98 ) );
  NAND2_X1 u1_u6_u6_U58 (.ZN( u1_u6_u6_n122 ) , .A1( u1_u6_u6_n94 ) , .A2( u1_u6_u6_n97 ) );
  INV_X1 u1_u6_u6_U59 (.A( u1_u6_u6_n139 ) , .ZN( u1_u6_u6_n160 ) );
  AOI21_X1 u1_u6_u6_U6 (.B1( u1_u6_u6_n107 ) , .B2( u1_u6_u6_n132 ) , .A( u1_u6_u6_n158 ) , .ZN( u1_u6_u6_n88 ) );
  NAND2_X1 u1_u6_u6_U60 (.ZN( u1_u6_u6_n113 ) , .A1( u1_u6_u6_n96 ) , .A2( u1_u6_u6_n98 ) );
  NOR2_X1 u1_u6_u6_U61 (.A2( u1_u6_X_40 ) , .A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n126 ) );
  NOR2_X1 u1_u6_u6_U62 (.A2( u1_u6_X_39 ) , .A1( u1_u6_X_42 ) , .ZN( u1_u6_u6_n92 ) );
  NOR2_X1 u1_u6_u6_U63 (.A2( u1_u6_X_39 ) , .A1( u1_u6_u6_n156 ) , .ZN( u1_u6_u6_n97 ) );
  NOR2_X1 u1_u6_u6_U64 (.A2( u1_u6_X_38 ) , .A1( u1_u6_u6_n165 ) , .ZN( u1_u6_u6_n95 ) );
  NOR2_X1 u1_u6_u6_U65 (.A2( u1_u6_X_41 ) , .ZN( u1_u6_u6_n111 ) , .A1( u1_u6_u6_n157 ) );
  NOR2_X1 u1_u6_u6_U66 (.A2( u1_u6_X_37 ) , .A1( u1_u6_u6_n162 ) , .ZN( u1_u6_u6_n94 ) );
  NOR2_X1 u1_u6_u6_U67 (.A2( u1_u6_X_37 ) , .A1( u1_u6_X_38 ) , .ZN( u1_u6_u6_n91 ) );
  NAND2_X1 u1_u6_u6_U68 (.A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n144 ) , .A2( u1_u6_u6_n157 ) );
  NAND2_X1 u1_u6_u6_U69 (.A2( u1_u6_X_40 ) , .A1( u1_u6_X_41 ) , .ZN( u1_u6_u6_n139 ) );
  OAI21_X1 u1_u6_u6_U7 (.A( u1_u6_u6_n159 ) , .B1( u1_u6_u6_n169 ) , .B2( u1_u6_u6_n173 ) , .ZN( u1_u6_u6_n90 ) );
  AND2_X1 u1_u6_u6_U70 (.A1( u1_u6_X_39 ) , .A2( u1_u6_u6_n156 ) , .ZN( u1_u6_u6_n96 ) );
  AND2_X1 u1_u6_u6_U71 (.A1( u1_u6_X_39 ) , .A2( u1_u6_X_42 ) , .ZN( u1_u6_u6_n99 ) );
  INV_X1 u1_u6_u6_U72 (.A( u1_u6_X_40 ) , .ZN( u1_u6_u6_n157 ) );
  INV_X1 u1_u6_u6_U73 (.A( u1_u6_X_37 ) , .ZN( u1_u6_u6_n165 ) );
  INV_X1 u1_u6_u6_U74 (.A( u1_u6_X_38 ) , .ZN( u1_u6_u6_n162 ) );
  INV_X1 u1_u6_u6_U75 (.A( u1_u6_X_42 ) , .ZN( u1_u6_u6_n156 ) );
  NAND4_X1 u1_u6_u6_U76 (.ZN( u1_out6_12 ) , .A4( u1_u6_u6_n114 ) , .A3( u1_u6_u6_n115 ) , .A2( u1_u6_u6_n116 ) , .A1( u1_u6_u6_n117 ) );
  OAI22_X1 u1_u6_u6_U77 (.B2( u1_u6_u6_n111 ) , .ZN( u1_u6_u6_n116 ) , .B1( u1_u6_u6_n126 ) , .A2( u1_u6_u6_n164 ) , .A1( u1_u6_u6_n167 ) );
  OAI21_X1 u1_u6_u6_U78 (.A( u1_u6_u6_n108 ) , .ZN( u1_u6_u6_n117 ) , .B2( u1_u6_u6_n141 ) , .B1( u1_u6_u6_n163 ) );
  NAND4_X1 u1_u6_u6_U79 (.ZN( u1_out6_32 ) , .A4( u1_u6_u6_n103 ) , .A3( u1_u6_u6_n104 ) , .A2( u1_u6_u6_n105 ) , .A1( u1_u6_u6_n106 ) );
  INV_X1 u1_u6_u6_U8 (.ZN( u1_u6_u6_n172 ) , .A( u1_u6_u6_n88 ) );
  AOI22_X1 u1_u6_u6_U80 (.ZN( u1_u6_u6_n104 ) , .A1( u1_u6_u6_n111 ) , .B1( u1_u6_u6_n124 ) , .B2( u1_u6_u6_n151 ) , .A2( u1_u6_u6_n93 ) );
  AOI22_X1 u1_u6_u6_U81 (.ZN( u1_u6_u6_n105 ) , .A2( u1_u6_u6_n108 ) , .A1( u1_u6_u6_n118 ) , .B2( u1_u6_u6_n126 ) , .B1( u1_u6_u6_n171 ) );
  OAI211_X1 u1_u6_u6_U82 (.ZN( u1_out6_22 ) , .B( u1_u6_u6_n137 ) , .A( u1_u6_u6_n138 ) , .C2( u1_u6_u6_n139 ) , .C1( u1_u6_u6_n140 ) );
  AOI22_X1 u1_u6_u6_U83 (.B1( u1_u6_u6_n124 ) , .A2( u1_u6_u6_n125 ) , .A1( u1_u6_u6_n126 ) , .ZN( u1_u6_u6_n138 ) , .B2( u1_u6_u6_n161 ) );
  AND4_X1 u1_u6_u6_U84 (.A3( u1_u6_u6_n119 ) , .A1( u1_u6_u6_n120 ) , .A4( u1_u6_u6_n129 ) , .ZN( u1_u6_u6_n140 ) , .A2( u1_u6_u6_n143 ) );
  OAI211_X1 u1_u6_u6_U85 (.ZN( u1_out6_7 ) , .B( u1_u6_u6_n153 ) , .C2( u1_u6_u6_n154 ) , .C1( u1_u6_u6_n155 ) , .A( u1_u6_u6_n174 ) );
  NOR3_X1 u1_u6_u6_U86 (.A1( u1_u6_u6_n141 ) , .ZN( u1_u6_u6_n154 ) , .A3( u1_u6_u6_n164 ) , .A2( u1_u6_u6_n171 ) );
  INV_X1 u1_u6_u6_U87 (.A( u1_u6_u6_n142 ) , .ZN( u1_u6_u6_n174 ) );
  NAND3_X1 u1_u6_u6_U88 (.A2( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n125 ) , .A1( u1_u6_u6_n130 ) , .A3( u1_u6_u6_n131 ) );
  NAND3_X1 u1_u6_u6_U89 (.A3( u1_u6_u6_n133 ) , .ZN( u1_u6_u6_n141 ) , .A1( u1_u6_u6_n145 ) , .A2( u1_u6_u6_n148 ) );
  AOI22_X1 u1_u6_u6_U9 (.A2( u1_u6_u6_n151 ) , .B2( u1_u6_u6_n161 ) , .A1( u1_u6_u6_n167 ) , .B1( u1_u6_u6_n170 ) , .ZN( u1_u6_u6_n89 ) );
  NAND3_X1 u1_u6_u6_U90 (.ZN( u1_u6_u6_n101 ) , .A3( u1_u6_u6_n107 ) , .A2( u1_u6_u6_n121 ) , .A1( u1_u6_u6_n127 ) );
  NAND3_X1 u1_u6_u6_U91 (.ZN( u1_u6_u6_n102 ) , .A3( u1_u6_u6_n130 ) , .A2( u1_u6_u6_n145 ) , .A1( u1_u6_u6_n166 ) );
  NAND3_X1 u1_u6_u6_U92 (.A3( u1_u6_u6_n113 ) , .A1( u1_u6_u6_n119 ) , .A2( u1_u6_u6_n123 ) , .ZN( u1_u6_u6_n93 ) );
  NAND3_X1 u1_u6_u6_U93 (.ZN( u1_u6_u6_n142 ) , .A2( u1_u6_u6_n172 ) , .A3( u1_u6_u6_n89 ) , .A1( u1_u6_u6_n90 ) );
  XOR2_X1 u1_u7_U35 (.B( u1_K8_22 ) , .A( u1_R6_15 ) , .Z( u1_u7_X_22 ) );
  XOR2_X1 u1_u7_U36 (.B( u1_K8_21 ) , .A( u1_R6_14 ) , .Z( u1_u7_X_21 ) );
  OAI22_X1 u1_u7_u3_U10 (.B1( u1_u7_u3_n113 ) , .A2( u1_u7_u3_n135 ) , .A1( u1_u7_u3_n150 ) , .B2( u1_u7_u3_n164 ) , .ZN( u1_u7_u3_n98 ) );
  OAI211_X1 u1_u7_u3_U11 (.B( u1_u7_u3_n106 ) , .ZN( u1_u7_u3_n119 ) , .C2( u1_u7_u3_n128 ) , .C1( u1_u7_u3_n167 ) , .A( u1_u7_u3_n181 ) );
  AOI221_X1 u1_u7_u3_U12 (.C1( u1_u7_u3_n105 ) , .ZN( u1_u7_u3_n106 ) , .A( u1_u7_u3_n131 ) , .B2( u1_u7_u3_n132 ) , .C2( u1_u7_u3_n133 ) , .B1( u1_u7_u3_n169 ) );
  INV_X1 u1_u7_u3_U13 (.ZN( u1_u7_u3_n181 ) , .A( u1_u7_u3_n98 ) );
  NAND2_X1 u1_u7_u3_U14 (.ZN( u1_u7_u3_n105 ) , .A2( u1_u7_u3_n130 ) , .A1( u1_u7_u3_n155 ) );
  AOI22_X1 u1_u7_u3_U15 (.B1( u1_u7_u3_n115 ) , .A2( u1_u7_u3_n116 ) , .ZN( u1_u7_u3_n123 ) , .B2( u1_u7_u3_n133 ) , .A1( u1_u7_u3_n169 ) );
  NAND2_X1 u1_u7_u3_U16 (.ZN( u1_u7_u3_n116 ) , .A2( u1_u7_u3_n151 ) , .A1( u1_u7_u3_n182 ) );
  NOR2_X1 u1_u7_u3_U17 (.ZN( u1_u7_u3_n126 ) , .A2( u1_u7_u3_n150 ) , .A1( u1_u7_u3_n164 ) );
  AOI21_X1 u1_u7_u3_U18 (.ZN( u1_u7_u3_n112 ) , .B2( u1_u7_u3_n146 ) , .B1( u1_u7_u3_n155 ) , .A( u1_u7_u3_n167 ) );
  NAND2_X1 u1_u7_u3_U19 (.A1( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n142 ) , .A2( u1_u7_u3_n164 ) );
  NAND2_X1 u1_u7_u3_U20 (.ZN( u1_u7_u3_n132 ) , .A2( u1_u7_u3_n152 ) , .A1( u1_u7_u3_n156 ) );
  AND2_X1 u1_u7_u3_U21 (.A2( u1_u7_u3_n113 ) , .A1( u1_u7_u3_n114 ) , .ZN( u1_u7_u3_n151 ) );
  INV_X1 u1_u7_u3_U22 (.A( u1_u7_u3_n133 ) , .ZN( u1_u7_u3_n165 ) );
  INV_X1 u1_u7_u3_U23 (.A( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n170 ) );
  NAND2_X1 u1_u7_u3_U24 (.A1( u1_u7_u3_n107 ) , .A2( u1_u7_u3_n108 ) , .ZN( u1_u7_u3_n140 ) );
  NAND2_X1 u1_u7_u3_U25 (.ZN( u1_u7_u3_n117 ) , .A1( u1_u7_u3_n124 ) , .A2( u1_u7_u3_n148 ) );
  NAND2_X1 u1_u7_u3_U26 (.ZN( u1_u7_u3_n143 ) , .A1( u1_u7_u3_n165 ) , .A2( u1_u7_u3_n167 ) );
  INV_X1 u1_u7_u3_U27 (.A( u1_u7_u3_n130 ) , .ZN( u1_u7_u3_n177 ) );
  INV_X1 u1_u7_u3_U28 (.A( u1_u7_u3_n128 ) , .ZN( u1_u7_u3_n176 ) );
  INV_X1 u1_u7_u3_U29 (.A( u1_u7_u3_n155 ) , .ZN( u1_u7_u3_n174 ) );
  INV_X1 u1_u7_u3_U3 (.A( u1_u7_u3_n129 ) , .ZN( u1_u7_u3_n183 ) );
  INV_X1 u1_u7_u3_U30 (.A( u1_u7_u3_n139 ) , .ZN( u1_u7_u3_n185 ) );
  NOR2_X1 u1_u7_u3_U31 (.ZN( u1_u7_u3_n135 ) , .A2( u1_u7_u3_n141 ) , .A1( u1_u7_u3_n169 ) );
  OAI222_X1 u1_u7_u3_U32 (.C2( u1_u7_u3_n107 ) , .A2( u1_u7_u3_n108 ) , .B1( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n138 ) , .B2( u1_u7_u3_n146 ) , .C1( u1_u7_u3_n154 ) , .A1( u1_u7_u3_n164 ) );
  NOR4_X1 u1_u7_u3_U33 (.A4( u1_u7_u3_n157 ) , .A3( u1_u7_u3_n158 ) , .A2( u1_u7_u3_n159 ) , .A1( u1_u7_u3_n160 ) , .ZN( u1_u7_u3_n161 ) );
  AOI21_X1 u1_u7_u3_U34 (.B2( u1_u7_u3_n152 ) , .B1( u1_u7_u3_n153 ) , .ZN( u1_u7_u3_n158 ) , .A( u1_u7_u3_n164 ) );
  AOI21_X1 u1_u7_u3_U35 (.A( u1_u7_u3_n154 ) , .B2( u1_u7_u3_n155 ) , .B1( u1_u7_u3_n156 ) , .ZN( u1_u7_u3_n157 ) );
  AOI21_X1 u1_u7_u3_U36 (.A( u1_u7_u3_n149 ) , .B2( u1_u7_u3_n150 ) , .B1( u1_u7_u3_n151 ) , .ZN( u1_u7_u3_n159 ) );
  AOI211_X1 u1_u7_u3_U37 (.ZN( u1_u7_u3_n109 ) , .A( u1_u7_u3_n119 ) , .C2( u1_u7_u3_n129 ) , .B( u1_u7_u3_n138 ) , .C1( u1_u7_u3_n141 ) );
  AOI211_X1 u1_u7_u3_U38 (.B( u1_u7_u3_n119 ) , .A( u1_u7_u3_n120 ) , .C2( u1_u7_u3_n121 ) , .ZN( u1_u7_u3_n122 ) , .C1( u1_u7_u3_n179 ) );
  INV_X1 u1_u7_u3_U39 (.A( u1_u7_u3_n156 ) , .ZN( u1_u7_u3_n179 ) );
  INV_X1 u1_u7_u3_U4 (.A( u1_u7_u3_n140 ) , .ZN( u1_u7_u3_n182 ) );
  OAI22_X1 u1_u7_u3_U40 (.B1( u1_u7_u3_n118 ) , .ZN( u1_u7_u3_n120 ) , .A1( u1_u7_u3_n135 ) , .B2( u1_u7_u3_n154 ) , .A2( u1_u7_u3_n178 ) );
  AND3_X1 u1_u7_u3_U41 (.ZN( u1_u7_u3_n118 ) , .A2( u1_u7_u3_n124 ) , .A1( u1_u7_u3_n144 ) , .A3( u1_u7_u3_n152 ) );
  INV_X1 u1_u7_u3_U42 (.A( u1_u7_u3_n121 ) , .ZN( u1_u7_u3_n164 ) );
  NAND2_X1 u1_u7_u3_U43 (.ZN( u1_u7_u3_n133 ) , .A1( u1_u7_u3_n154 ) , .A2( u1_u7_u3_n164 ) );
  OAI211_X1 u1_u7_u3_U44 (.B( u1_u7_u3_n127 ) , .ZN( u1_u7_u3_n139 ) , .C1( u1_u7_u3_n150 ) , .C2( u1_u7_u3_n154 ) , .A( u1_u7_u3_n184 ) );
  INV_X1 u1_u7_u3_U45 (.A( u1_u7_u3_n125 ) , .ZN( u1_u7_u3_n184 ) );
  AOI221_X1 u1_u7_u3_U46 (.A( u1_u7_u3_n126 ) , .ZN( u1_u7_u3_n127 ) , .C2( u1_u7_u3_n132 ) , .C1( u1_u7_u3_n169 ) , .B2( u1_u7_u3_n170 ) , .B1( u1_u7_u3_n174 ) );
  OAI22_X1 u1_u7_u3_U47 (.A1( u1_u7_u3_n124 ) , .ZN( u1_u7_u3_n125 ) , .B2( u1_u7_u3_n145 ) , .A2( u1_u7_u3_n165 ) , .B1( u1_u7_u3_n167 ) );
  NOR2_X1 u1_u7_u3_U48 (.A1( u1_u7_u3_n113 ) , .ZN( u1_u7_u3_n131 ) , .A2( u1_u7_u3_n154 ) );
  NAND2_X1 u1_u7_u3_U49 (.A1( u1_u7_u3_n103 ) , .ZN( u1_u7_u3_n150 ) , .A2( u1_u7_u3_n99 ) );
  INV_X1 u1_u7_u3_U5 (.A( u1_u7_u3_n117 ) , .ZN( u1_u7_u3_n178 ) );
  NAND2_X1 u1_u7_u3_U50 (.A2( u1_u7_u3_n102 ) , .ZN( u1_u7_u3_n155 ) , .A1( u1_u7_u3_n97 ) );
  INV_X1 u1_u7_u3_U51 (.A( u1_u7_u3_n141 ) , .ZN( u1_u7_u3_n167 ) );
  AOI21_X1 u1_u7_u3_U52 (.B2( u1_u7_u3_n114 ) , .B1( u1_u7_u3_n146 ) , .A( u1_u7_u3_n154 ) , .ZN( u1_u7_u3_n94 ) );
  AOI21_X1 u1_u7_u3_U53 (.ZN( u1_u7_u3_n110 ) , .B2( u1_u7_u3_n142 ) , .B1( u1_u7_u3_n186 ) , .A( u1_u7_u3_n95 ) );
  INV_X1 u1_u7_u3_U54 (.A( u1_u7_u3_n145 ) , .ZN( u1_u7_u3_n186 ) );
  AOI21_X1 u1_u7_u3_U55 (.B1( u1_u7_u3_n124 ) , .A( u1_u7_u3_n149 ) , .B2( u1_u7_u3_n155 ) , .ZN( u1_u7_u3_n95 ) );
  INV_X1 u1_u7_u3_U56 (.A( u1_u7_u3_n149 ) , .ZN( u1_u7_u3_n169 ) );
  NAND2_X1 u1_u7_u3_U57 (.ZN( u1_u7_u3_n124 ) , .A1( u1_u7_u3_n96 ) , .A2( u1_u7_u3_n97 ) );
  NAND2_X1 u1_u7_u3_U58 (.A2( u1_u7_u3_n100 ) , .ZN( u1_u7_u3_n146 ) , .A1( u1_u7_u3_n96 ) );
  NAND2_X1 u1_u7_u3_U59 (.A1( u1_u7_u3_n101 ) , .ZN( u1_u7_u3_n145 ) , .A2( u1_u7_u3_n99 ) );
  AOI221_X1 u1_u7_u3_U6 (.A( u1_u7_u3_n131 ) , .C2( u1_u7_u3_n132 ) , .C1( u1_u7_u3_n133 ) , .ZN( u1_u7_u3_n134 ) , .B1( u1_u7_u3_n143 ) , .B2( u1_u7_u3_n177 ) );
  NAND2_X1 u1_u7_u3_U60 (.A1( u1_u7_u3_n100 ) , .ZN( u1_u7_u3_n156 ) , .A2( u1_u7_u3_n99 ) );
  NAND2_X1 u1_u7_u3_U61 (.A2( u1_u7_u3_n101 ) , .A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n148 ) );
  NAND2_X1 u1_u7_u3_U62 (.A1( u1_u7_u3_n100 ) , .A2( u1_u7_u3_n102 ) , .ZN( u1_u7_u3_n128 ) );
  NAND2_X1 u1_u7_u3_U63 (.A2( u1_u7_u3_n101 ) , .A1( u1_u7_u3_n102 ) , .ZN( u1_u7_u3_n152 ) );
  NAND2_X1 u1_u7_u3_U64 (.A2( u1_u7_u3_n101 ) , .ZN( u1_u7_u3_n114 ) , .A1( u1_u7_u3_n96 ) );
  NAND2_X1 u1_u7_u3_U65 (.ZN( u1_u7_u3_n107 ) , .A1( u1_u7_u3_n97 ) , .A2( u1_u7_u3_n99 ) );
  NAND2_X1 u1_u7_u3_U66 (.A2( u1_u7_u3_n100 ) , .A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n113 ) );
  NAND2_X1 u1_u7_u3_U67 (.A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n153 ) , .A2( u1_u7_u3_n97 ) );
  NAND2_X1 u1_u7_u3_U68 (.A2( u1_u7_u3_n103 ) , .A1( u1_u7_u3_n104 ) , .ZN( u1_u7_u3_n130 ) );
  NAND2_X1 u1_u7_u3_U69 (.A2( u1_u7_u3_n103 ) , .ZN( u1_u7_u3_n144 ) , .A1( u1_u7_u3_n96 ) );
  OAI22_X1 u1_u7_u3_U7 (.B2( u1_u7_u3_n147 ) , .A2( u1_u7_u3_n148 ) , .ZN( u1_u7_u3_n160 ) , .B1( u1_u7_u3_n165 ) , .A1( u1_u7_u3_n168 ) );
  NAND2_X1 u1_u7_u3_U70 (.A1( u1_u7_u3_n102 ) , .A2( u1_u7_u3_n103 ) , .ZN( u1_u7_u3_n108 ) );
  NOR2_X1 u1_u7_u3_U71 (.A2( u1_u7_X_19 ) , .A1( u1_u7_X_20 ) , .ZN( u1_u7_u3_n99 ) );
  NOR2_X1 u1_u7_u3_U72 (.A2( u1_u7_X_21 ) , .A1( u1_u7_X_24 ) , .ZN( u1_u7_u3_n103 ) );
  NOR2_X1 u1_u7_u3_U73 (.A2( u1_u7_X_24 ) , .A1( u1_u7_u3_n171 ) , .ZN( u1_u7_u3_n97 ) );
  NOR2_X1 u1_u7_u3_U74 (.A2( u1_u7_X_23 ) , .ZN( u1_u7_u3_n141 ) , .A1( u1_u7_u3_n166 ) );
  NOR2_X1 u1_u7_u3_U75 (.A2( u1_u7_X_19 ) , .A1( u1_u7_u3_n172 ) , .ZN( u1_u7_u3_n96 ) );
  NAND2_X1 u1_u7_u3_U76 (.A1( u1_u7_X_22 ) , .A2( u1_u7_X_23 ) , .ZN( u1_u7_u3_n154 ) );
  NAND2_X1 u1_u7_u3_U77 (.A1( u1_u7_X_23 ) , .ZN( u1_u7_u3_n149 ) , .A2( u1_u7_u3_n166 ) );
  NOR2_X1 u1_u7_u3_U78 (.A2( u1_u7_X_22 ) , .A1( u1_u7_X_23 ) , .ZN( u1_u7_u3_n121 ) );
  AND2_X1 u1_u7_u3_U79 (.A1( u1_u7_X_24 ) , .ZN( u1_u7_u3_n101 ) , .A2( u1_u7_u3_n171 ) );
  AND3_X1 u1_u7_u3_U8 (.A3( u1_u7_u3_n144 ) , .A2( u1_u7_u3_n145 ) , .A1( u1_u7_u3_n146 ) , .ZN( u1_u7_u3_n147 ) );
  AND2_X1 u1_u7_u3_U80 (.A1( u1_u7_X_19 ) , .ZN( u1_u7_u3_n102 ) , .A2( u1_u7_u3_n172 ) );
  AND2_X1 u1_u7_u3_U81 (.A1( u1_u7_X_21 ) , .A2( u1_u7_X_24 ) , .ZN( u1_u7_u3_n100 ) );
  AND2_X1 u1_u7_u3_U82 (.A2( u1_u7_X_19 ) , .A1( u1_u7_X_20 ) , .ZN( u1_u7_u3_n104 ) );
  INV_X1 u1_u7_u3_U83 (.A( u1_u7_X_22 ) , .ZN( u1_u7_u3_n166 ) );
  INV_X1 u1_u7_u3_U84 (.A( u1_u7_X_21 ) , .ZN( u1_u7_u3_n171 ) );
  INV_X1 u1_u7_u3_U85 (.A( u1_u7_X_20 ) , .ZN( u1_u7_u3_n172 ) );
  OR4_X1 u1_u7_u3_U86 (.ZN( u1_out7_10 ) , .A4( u1_u7_u3_n136 ) , .A3( u1_u7_u3_n137 ) , .A1( u1_u7_u3_n138 ) , .A2( u1_u7_u3_n139 ) );
  OAI222_X1 u1_u7_u3_U87 (.C1( u1_u7_u3_n128 ) , .ZN( u1_u7_u3_n137 ) , .B1( u1_u7_u3_n148 ) , .A2( u1_u7_u3_n150 ) , .B2( u1_u7_u3_n154 ) , .C2( u1_u7_u3_n164 ) , .A1( u1_u7_u3_n167 ) );
  OAI221_X1 u1_u7_u3_U88 (.A( u1_u7_u3_n134 ) , .B2( u1_u7_u3_n135 ) , .ZN( u1_u7_u3_n136 ) , .C1( u1_u7_u3_n149 ) , .B1( u1_u7_u3_n151 ) , .C2( u1_u7_u3_n183 ) );
  NAND4_X1 u1_u7_u3_U89 (.ZN( u1_out7_26 ) , .A4( u1_u7_u3_n109 ) , .A3( u1_u7_u3_n110 ) , .A2( u1_u7_u3_n111 ) , .A1( u1_u7_u3_n173 ) );
  INV_X1 u1_u7_u3_U9 (.A( u1_u7_u3_n143 ) , .ZN( u1_u7_u3_n168 ) );
  INV_X1 u1_u7_u3_U90 (.ZN( u1_u7_u3_n173 ) , .A( u1_u7_u3_n94 ) );
  OAI21_X1 u1_u7_u3_U91 (.ZN( u1_u7_u3_n111 ) , .B2( u1_u7_u3_n117 ) , .A( u1_u7_u3_n133 ) , .B1( u1_u7_u3_n176 ) );
  NAND4_X1 u1_u7_u3_U92 (.ZN( u1_out7_20 ) , .A4( u1_u7_u3_n122 ) , .A3( u1_u7_u3_n123 ) , .A1( u1_u7_u3_n175 ) , .A2( u1_u7_u3_n180 ) );
  INV_X1 u1_u7_u3_U93 (.A( u1_u7_u3_n126 ) , .ZN( u1_u7_u3_n180 ) );
  INV_X1 u1_u7_u3_U94 (.A( u1_u7_u3_n112 ) , .ZN( u1_u7_u3_n175 ) );
  NAND4_X1 u1_u7_u3_U95 (.ZN( u1_out7_1 ) , .A4( u1_u7_u3_n161 ) , .A3( u1_u7_u3_n162 ) , .A2( u1_u7_u3_n163 ) , .A1( u1_u7_u3_n185 ) );
  NAND2_X1 u1_u7_u3_U96 (.ZN( u1_u7_u3_n163 ) , .A2( u1_u7_u3_n170 ) , .A1( u1_u7_u3_n176 ) );
  AOI22_X1 u1_u7_u3_U97 (.B2( u1_u7_u3_n140 ) , .B1( u1_u7_u3_n141 ) , .A2( u1_u7_u3_n142 ) , .ZN( u1_u7_u3_n162 ) , .A1( u1_u7_u3_n177 ) );
  NAND3_X1 u1_u7_u3_U98 (.A1( u1_u7_u3_n114 ) , .ZN( u1_u7_u3_n115 ) , .A2( u1_u7_u3_n145 ) , .A3( u1_u7_u3_n153 ) );
  NAND3_X1 u1_u7_u3_U99 (.ZN( u1_u7_u3_n129 ) , .A2( u1_u7_u3_n144 ) , .A1( u1_u7_u3_n153 ) , .A3( u1_u7_u3_n182 ) );
  XOR2_X1 u1_u8_U22 (.B( u1_K9_34 ) , .A( u1_R7_23 ) , .Z( u1_u8_X_34 ) );
  XOR2_X1 u1_u8_U23 (.B( u1_K9_33 ) , .A( u1_R7_22 ) , .Z( u1_u8_X_33 ) );
  NOR2_X1 u1_u8_u5_U10 (.ZN( u1_u8_u5_n135 ) , .A1( u1_u8_u5_n173 ) , .A2( u1_u8_u5_n176 ) );
  NOR3_X1 u1_u8_u5_U100 (.A3( u1_u8_u5_n141 ) , .A1( u1_u8_u5_n142 ) , .ZN( u1_u8_u5_n143 ) , .A2( u1_u8_u5_n191 ) );
  NAND4_X1 u1_u8_u5_U101 (.ZN( u1_out8_4 ) , .A4( u1_u8_u5_n112 ) , .A2( u1_u8_u5_n113 ) , .A1( u1_u8_u5_n114 ) , .A3( u1_u8_u5_n195 ) );
  AOI211_X1 u1_u8_u5_U102 (.A( u1_u8_u5_n110 ) , .C1( u1_u8_u5_n111 ) , .ZN( u1_u8_u5_n112 ) , .B( u1_u8_u5_n118 ) , .C2( u1_u8_u5_n177 ) );
  INV_X1 u1_u8_u5_U103 (.A( u1_u8_u5_n102 ) , .ZN( u1_u8_u5_n195 ) );
  NAND3_X1 u1_u8_u5_U104 (.A2( u1_u8_u5_n154 ) , .A3( u1_u8_u5_n158 ) , .A1( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n99 ) );
  INV_X1 u1_u8_u5_U11 (.A( u1_u8_u5_n121 ) , .ZN( u1_u8_u5_n177 ) );
  NOR2_X1 u1_u8_u5_U12 (.ZN( u1_u8_u5_n160 ) , .A2( u1_u8_u5_n173 ) , .A1( u1_u8_u5_n177 ) );
  INV_X1 u1_u8_u5_U13 (.A( u1_u8_u5_n150 ) , .ZN( u1_u8_u5_n174 ) );
  AOI21_X1 u1_u8_u5_U14 (.A( u1_u8_u5_n160 ) , .B2( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n162 ) , .B1( u1_u8_u5_n192 ) );
  INV_X1 u1_u8_u5_U15 (.A( u1_u8_u5_n159 ) , .ZN( u1_u8_u5_n192 ) );
  AOI21_X1 u1_u8_u5_U16 (.A( u1_u8_u5_n156 ) , .B2( u1_u8_u5_n157 ) , .B1( u1_u8_u5_n158 ) , .ZN( u1_u8_u5_n163 ) );
  AOI21_X1 u1_u8_u5_U17 (.B2( u1_u8_u5_n139 ) , .B1( u1_u8_u5_n140 ) , .ZN( u1_u8_u5_n141 ) , .A( u1_u8_u5_n150 ) );
  OAI21_X1 u1_u8_u5_U18 (.A( u1_u8_u5_n133 ) , .B2( u1_u8_u5_n134 ) , .B1( u1_u8_u5_n135 ) , .ZN( u1_u8_u5_n142 ) );
  OAI21_X1 u1_u8_u5_U19 (.ZN( u1_u8_u5_n133 ) , .B2( u1_u8_u5_n147 ) , .A( u1_u8_u5_n173 ) , .B1( u1_u8_u5_n188 ) );
  NAND2_X1 u1_u8_u5_U20 (.A2( u1_u8_u5_n119 ) , .A1( u1_u8_u5_n123 ) , .ZN( u1_u8_u5_n137 ) );
  INV_X1 u1_u8_u5_U21 (.A( u1_u8_u5_n155 ) , .ZN( u1_u8_u5_n194 ) );
  NAND2_X1 u1_u8_u5_U22 (.A1( u1_u8_u5_n121 ) , .ZN( u1_u8_u5_n132 ) , .A2( u1_u8_u5_n172 ) );
  NAND2_X1 u1_u8_u5_U23 (.A2( u1_u8_u5_n122 ) , .ZN( u1_u8_u5_n136 ) , .A1( u1_u8_u5_n154 ) );
  NAND2_X1 u1_u8_u5_U24 (.A2( u1_u8_u5_n119 ) , .A1( u1_u8_u5_n120 ) , .ZN( u1_u8_u5_n159 ) );
  INV_X1 u1_u8_u5_U25 (.A( u1_u8_u5_n156 ) , .ZN( u1_u8_u5_n175 ) );
  INV_X1 u1_u8_u5_U26 (.A( u1_u8_u5_n158 ) , .ZN( u1_u8_u5_n188 ) );
  INV_X1 u1_u8_u5_U27 (.A( u1_u8_u5_n152 ) , .ZN( u1_u8_u5_n179 ) );
  INV_X1 u1_u8_u5_U28 (.A( u1_u8_u5_n140 ) , .ZN( u1_u8_u5_n182 ) );
  INV_X1 u1_u8_u5_U29 (.A( u1_u8_u5_n151 ) , .ZN( u1_u8_u5_n183 ) );
  NOR2_X1 u1_u8_u5_U3 (.ZN( u1_u8_u5_n134 ) , .A1( u1_u8_u5_n183 ) , .A2( u1_u8_u5_n190 ) );
  INV_X1 u1_u8_u5_U30 (.A( u1_u8_u5_n123 ) , .ZN( u1_u8_u5_n185 ) );
  INV_X1 u1_u8_u5_U31 (.A( u1_u8_u5_n161 ) , .ZN( u1_u8_u5_n184 ) );
  INV_X1 u1_u8_u5_U32 (.A( u1_u8_u5_n139 ) , .ZN( u1_u8_u5_n189 ) );
  INV_X1 u1_u8_u5_U33 (.A( u1_u8_u5_n157 ) , .ZN( u1_u8_u5_n190 ) );
  INV_X1 u1_u8_u5_U34 (.A( u1_u8_u5_n120 ) , .ZN( u1_u8_u5_n193 ) );
  NAND2_X1 u1_u8_u5_U35 (.ZN( u1_u8_u5_n111 ) , .A1( u1_u8_u5_n140 ) , .A2( u1_u8_u5_n155 ) );
  INV_X1 u1_u8_u5_U36 (.A( u1_u8_u5_n117 ) , .ZN( u1_u8_u5_n196 ) );
  OAI221_X1 u1_u8_u5_U37 (.A( u1_u8_u5_n116 ) , .ZN( u1_u8_u5_n117 ) , .B2( u1_u8_u5_n119 ) , .C1( u1_u8_u5_n153 ) , .C2( u1_u8_u5_n158 ) , .B1( u1_u8_u5_n172 ) );
  AOI222_X1 u1_u8_u5_U38 (.ZN( u1_u8_u5_n116 ) , .B2( u1_u8_u5_n145 ) , .C1( u1_u8_u5_n148 ) , .A2( u1_u8_u5_n174 ) , .C2( u1_u8_u5_n177 ) , .B1( u1_u8_u5_n187 ) , .A1( u1_u8_u5_n193 ) );
  INV_X1 u1_u8_u5_U39 (.A( u1_u8_u5_n115 ) , .ZN( u1_u8_u5_n187 ) );
  INV_X1 u1_u8_u5_U4 (.A( u1_u8_u5_n138 ) , .ZN( u1_u8_u5_n191 ) );
  NOR2_X1 u1_u8_u5_U40 (.ZN( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n170 ) , .A2( u1_u8_u5_n180 ) );
  OAI221_X1 u1_u8_u5_U41 (.A( u1_u8_u5_n101 ) , .ZN( u1_u8_u5_n102 ) , .C2( u1_u8_u5_n115 ) , .C1( u1_u8_u5_n126 ) , .B1( u1_u8_u5_n134 ) , .B2( u1_u8_u5_n160 ) );
  OAI21_X1 u1_u8_u5_U42 (.ZN( u1_u8_u5_n101 ) , .B1( u1_u8_u5_n137 ) , .A( u1_u8_u5_n146 ) , .B2( u1_u8_u5_n147 ) );
  AOI22_X1 u1_u8_u5_U43 (.B2( u1_u8_u5_n131 ) , .A2( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n169 ) , .B1( u1_u8_u5_n174 ) , .A1( u1_u8_u5_n185 ) );
  NOR2_X1 u1_u8_u5_U44 (.A1( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n150 ) , .A2( u1_u8_u5_n173 ) );
  AOI21_X1 u1_u8_u5_U45 (.A( u1_u8_u5_n118 ) , .B2( u1_u8_u5_n145 ) , .ZN( u1_u8_u5_n168 ) , .B1( u1_u8_u5_n186 ) );
  INV_X1 u1_u8_u5_U46 (.A( u1_u8_u5_n122 ) , .ZN( u1_u8_u5_n186 ) );
  NOR2_X1 u1_u8_u5_U47 (.A1( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n152 ) , .A2( u1_u8_u5_n176 ) );
  NOR2_X1 u1_u8_u5_U48 (.A1( u1_u8_u5_n115 ) , .ZN( u1_u8_u5_n118 ) , .A2( u1_u8_u5_n153 ) );
  NOR2_X1 u1_u8_u5_U49 (.A2( u1_u8_u5_n145 ) , .ZN( u1_u8_u5_n156 ) , .A1( u1_u8_u5_n174 ) );
  OAI21_X1 u1_u8_u5_U5 (.B2( u1_u8_u5_n136 ) , .B1( u1_u8_u5_n137 ) , .ZN( u1_u8_u5_n138 ) , .A( u1_u8_u5_n177 ) );
  NOR2_X1 u1_u8_u5_U50 (.ZN( u1_u8_u5_n121 ) , .A2( u1_u8_u5_n145 ) , .A1( u1_u8_u5_n176 ) );
  AOI22_X1 u1_u8_u5_U51 (.ZN( u1_u8_u5_n114 ) , .A2( u1_u8_u5_n137 ) , .A1( u1_u8_u5_n145 ) , .B2( u1_u8_u5_n175 ) , .B1( u1_u8_u5_n193 ) );
  OAI211_X1 u1_u8_u5_U52 (.B( u1_u8_u5_n124 ) , .A( u1_u8_u5_n125 ) , .C2( u1_u8_u5_n126 ) , .C1( u1_u8_u5_n127 ) , .ZN( u1_u8_u5_n128 ) );
  NOR3_X1 u1_u8_u5_U53 (.ZN( u1_u8_u5_n127 ) , .A1( u1_u8_u5_n136 ) , .A3( u1_u8_u5_n148 ) , .A2( u1_u8_u5_n182 ) );
  OAI21_X1 u1_u8_u5_U54 (.ZN( u1_u8_u5_n124 ) , .A( u1_u8_u5_n177 ) , .B2( u1_u8_u5_n183 ) , .B1( u1_u8_u5_n189 ) );
  OAI21_X1 u1_u8_u5_U55 (.ZN( u1_u8_u5_n125 ) , .A( u1_u8_u5_n174 ) , .B2( u1_u8_u5_n185 ) , .B1( u1_u8_u5_n190 ) );
  AOI21_X1 u1_u8_u5_U56 (.A( u1_u8_u5_n153 ) , .B2( u1_u8_u5_n154 ) , .B1( u1_u8_u5_n155 ) , .ZN( u1_u8_u5_n164 ) );
  AOI21_X1 u1_u8_u5_U57 (.ZN( u1_u8_u5_n110 ) , .B1( u1_u8_u5_n122 ) , .B2( u1_u8_u5_n139 ) , .A( u1_u8_u5_n153 ) );
  INV_X1 u1_u8_u5_U58 (.A( u1_u8_u5_n153 ) , .ZN( u1_u8_u5_n176 ) );
  INV_X1 u1_u8_u5_U59 (.A( u1_u8_u5_n126 ) , .ZN( u1_u8_u5_n173 ) );
  AOI222_X1 u1_u8_u5_U6 (.ZN( u1_u8_u5_n113 ) , .A1( u1_u8_u5_n131 ) , .C1( u1_u8_u5_n148 ) , .B2( u1_u8_u5_n174 ) , .C2( u1_u8_u5_n178 ) , .A2( u1_u8_u5_n179 ) , .B1( u1_u8_u5_n99 ) );
  AND2_X1 u1_u8_u5_U60 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n147 ) );
  AND2_X1 u1_u8_u5_U61 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n148 ) );
  NAND2_X1 u1_u8_u5_U62 (.A1( u1_u8_u5_n105 ) , .A2( u1_u8_u5_n106 ) , .ZN( u1_u8_u5_n158 ) );
  NAND2_X1 u1_u8_u5_U63 (.A2( u1_u8_u5_n108 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n139 ) );
  NAND2_X1 u1_u8_u5_U64 (.A1( u1_u8_u5_n106 ) , .A2( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n119 ) );
  NAND2_X1 u1_u8_u5_U65 (.A2( u1_u8_u5_n103 ) , .A1( u1_u8_u5_n105 ) , .ZN( u1_u8_u5_n140 ) );
  NAND2_X1 u1_u8_u5_U66 (.A2( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n105 ) , .ZN( u1_u8_u5_n155 ) );
  NAND2_X1 u1_u8_u5_U67 (.A2( u1_u8_u5_n106 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n122 ) );
  NAND2_X1 u1_u8_u5_U68 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n106 ) , .ZN( u1_u8_u5_n115 ) );
  NAND2_X1 u1_u8_u5_U69 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n103 ) , .ZN( u1_u8_u5_n161 ) );
  INV_X1 u1_u8_u5_U7 (.A( u1_u8_u5_n135 ) , .ZN( u1_u8_u5_n178 ) );
  NAND2_X1 u1_u8_u5_U70 (.A1( u1_u8_u5_n105 ) , .A2( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n154 ) );
  INV_X1 u1_u8_u5_U71 (.A( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n172 ) );
  NAND2_X1 u1_u8_u5_U72 (.A1( u1_u8_u5_n103 ) , .A2( u1_u8_u5_n108 ) , .ZN( u1_u8_u5_n123 ) );
  NAND2_X1 u1_u8_u5_U73 (.A2( u1_u8_u5_n103 ) , .A1( u1_u8_u5_n107 ) , .ZN( u1_u8_u5_n151 ) );
  NAND2_X1 u1_u8_u5_U74 (.A2( u1_u8_u5_n107 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n120 ) );
  NAND2_X1 u1_u8_u5_U75 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n109 ) , .ZN( u1_u8_u5_n157 ) );
  AND2_X1 u1_u8_u5_U76 (.A2( u1_u8_u5_n100 ) , .A1( u1_u8_u5_n104 ) , .ZN( u1_u8_u5_n131 ) );
  NOR2_X1 u1_u8_u5_U77 (.A2( u1_u8_X_34 ) , .A1( u1_u8_X_35 ) , .ZN( u1_u8_u5_n145 ) );
  NOR2_X1 u1_u8_u5_U78 (.A2( u1_u8_X_34 ) , .ZN( u1_u8_u5_n146 ) , .A1( u1_u8_u5_n171 ) );
  NOR2_X1 u1_u8_u5_U79 (.A2( u1_u8_X_31 ) , .A1( u1_u8_X_32 ) , .ZN( u1_u8_u5_n103 ) );
  OAI22_X1 u1_u8_u5_U8 (.B2( u1_u8_u5_n149 ) , .B1( u1_u8_u5_n150 ) , .A2( u1_u8_u5_n151 ) , .A1( u1_u8_u5_n152 ) , .ZN( u1_u8_u5_n165 ) );
  NOR2_X1 u1_u8_u5_U80 (.A2( u1_u8_X_36 ) , .ZN( u1_u8_u5_n105 ) , .A1( u1_u8_u5_n180 ) );
  NOR2_X1 u1_u8_u5_U81 (.A2( u1_u8_X_33 ) , .ZN( u1_u8_u5_n108 ) , .A1( u1_u8_u5_n170 ) );
  NOR2_X1 u1_u8_u5_U82 (.A2( u1_u8_X_33 ) , .A1( u1_u8_X_36 ) , .ZN( u1_u8_u5_n107 ) );
  NOR2_X1 u1_u8_u5_U83 (.A2( u1_u8_X_31 ) , .ZN( u1_u8_u5_n104 ) , .A1( u1_u8_u5_n181 ) );
  NAND2_X1 u1_u8_u5_U84 (.A2( u1_u8_X_34 ) , .A1( u1_u8_X_35 ) , .ZN( u1_u8_u5_n153 ) );
  NAND2_X1 u1_u8_u5_U85 (.A1( u1_u8_X_34 ) , .ZN( u1_u8_u5_n126 ) , .A2( u1_u8_u5_n171 ) );
  AND2_X1 u1_u8_u5_U86 (.A1( u1_u8_X_31 ) , .A2( u1_u8_X_32 ) , .ZN( u1_u8_u5_n106 ) );
  AND2_X1 u1_u8_u5_U87 (.A1( u1_u8_X_31 ) , .ZN( u1_u8_u5_n109 ) , .A2( u1_u8_u5_n181 ) );
  INV_X1 u1_u8_u5_U88 (.A( u1_u8_X_33 ) , .ZN( u1_u8_u5_n180 ) );
  INV_X1 u1_u8_u5_U89 (.A( u1_u8_X_35 ) , .ZN( u1_u8_u5_n171 ) );
  NOR3_X1 u1_u8_u5_U9 (.A2( u1_u8_u5_n147 ) , .A1( u1_u8_u5_n148 ) , .ZN( u1_u8_u5_n149 ) , .A3( u1_u8_u5_n194 ) );
  INV_X1 u1_u8_u5_U90 (.A( u1_u8_X_36 ) , .ZN( u1_u8_u5_n170 ) );
  INV_X1 u1_u8_u5_U91 (.A( u1_u8_X_32 ) , .ZN( u1_u8_u5_n181 ) );
  NAND4_X1 u1_u8_u5_U92 (.ZN( u1_out8_29 ) , .A4( u1_u8_u5_n129 ) , .A3( u1_u8_u5_n130 ) , .A2( u1_u8_u5_n168 ) , .A1( u1_u8_u5_n196 ) );
  AOI221_X1 u1_u8_u5_U93 (.A( u1_u8_u5_n128 ) , .ZN( u1_u8_u5_n129 ) , .C2( u1_u8_u5_n132 ) , .B2( u1_u8_u5_n159 ) , .B1( u1_u8_u5_n176 ) , .C1( u1_u8_u5_n184 ) );
  AOI222_X1 u1_u8_u5_U94 (.ZN( u1_u8_u5_n130 ) , .A2( u1_u8_u5_n146 ) , .B1( u1_u8_u5_n147 ) , .C2( u1_u8_u5_n175 ) , .B2( u1_u8_u5_n179 ) , .A1( u1_u8_u5_n188 ) , .C1( u1_u8_u5_n194 ) );
  NAND4_X1 u1_u8_u5_U95 (.ZN( u1_out8_19 ) , .A4( u1_u8_u5_n166 ) , .A3( u1_u8_u5_n167 ) , .A2( u1_u8_u5_n168 ) , .A1( u1_u8_u5_n169 ) );
  AOI22_X1 u1_u8_u5_U96 (.B2( u1_u8_u5_n145 ) , .A2( u1_u8_u5_n146 ) , .ZN( u1_u8_u5_n167 ) , .B1( u1_u8_u5_n182 ) , .A1( u1_u8_u5_n189 ) );
  NOR4_X1 u1_u8_u5_U97 (.A4( u1_u8_u5_n162 ) , .A3( u1_u8_u5_n163 ) , .A2( u1_u8_u5_n164 ) , .A1( u1_u8_u5_n165 ) , .ZN( u1_u8_u5_n166 ) );
  NAND4_X1 u1_u8_u5_U98 (.ZN( u1_out8_11 ) , .A4( u1_u8_u5_n143 ) , .A3( u1_u8_u5_n144 ) , .A2( u1_u8_u5_n169 ) , .A1( u1_u8_u5_n196 ) );
  AOI22_X1 u1_u8_u5_U99 (.A2( u1_u8_u5_n132 ) , .ZN( u1_u8_u5_n144 ) , .B2( u1_u8_u5_n145 ) , .B1( u1_u8_u5_n184 ) , .A1( u1_u8_u5_n194 ) );
  XOR2_X1 u1_u9_U29 (.B( u1_K10_28 ) , .A( u1_R8_19 ) , .Z( u1_u9_X_28 ) );
  XOR2_X1 u1_u9_U30 (.B( u1_K10_27 ) , .A( u1_R8_18 ) , .Z( u1_u9_X_27 ) );
  OAI22_X1 u1_u9_u4_U10 (.B2( u1_u9_u4_n135 ) , .ZN( u1_u9_u4_n137 ) , .B1( u1_u9_u4_n153 ) , .A1( u1_u9_u4_n155 ) , .A2( u1_u9_u4_n171 ) );
  AND3_X1 u1_u9_u4_U11 (.A2( u1_u9_u4_n134 ) , .ZN( u1_u9_u4_n135 ) , .A3( u1_u9_u4_n145 ) , .A1( u1_u9_u4_n157 ) );
  NAND2_X1 u1_u9_u4_U12 (.ZN( u1_u9_u4_n132 ) , .A2( u1_u9_u4_n170 ) , .A1( u1_u9_u4_n173 ) );
  AOI21_X1 u1_u9_u4_U13 (.B2( u1_u9_u4_n160 ) , .B1( u1_u9_u4_n161 ) , .ZN( u1_u9_u4_n162 ) , .A( u1_u9_u4_n170 ) );
  AOI21_X1 u1_u9_u4_U14 (.ZN( u1_u9_u4_n107 ) , .B2( u1_u9_u4_n143 ) , .A( u1_u9_u4_n174 ) , .B1( u1_u9_u4_n184 ) );
  AOI21_X1 u1_u9_u4_U15 (.B2( u1_u9_u4_n158 ) , .B1( u1_u9_u4_n159 ) , .ZN( u1_u9_u4_n163 ) , .A( u1_u9_u4_n174 ) );
  AOI21_X1 u1_u9_u4_U16 (.A( u1_u9_u4_n153 ) , .B2( u1_u9_u4_n154 ) , .B1( u1_u9_u4_n155 ) , .ZN( u1_u9_u4_n165 ) );
  AOI21_X1 u1_u9_u4_U17 (.A( u1_u9_u4_n156 ) , .B2( u1_u9_u4_n157 ) , .ZN( u1_u9_u4_n164 ) , .B1( u1_u9_u4_n184 ) );
  INV_X1 u1_u9_u4_U18 (.A( u1_u9_u4_n138 ) , .ZN( u1_u9_u4_n170 ) );
  AND2_X1 u1_u9_u4_U19 (.A2( u1_u9_u4_n120 ) , .ZN( u1_u9_u4_n155 ) , .A1( u1_u9_u4_n160 ) );
  INV_X1 u1_u9_u4_U20 (.A( u1_u9_u4_n156 ) , .ZN( u1_u9_u4_n175 ) );
  NAND2_X1 u1_u9_u4_U21 (.A2( u1_u9_u4_n118 ) , .ZN( u1_u9_u4_n131 ) , .A1( u1_u9_u4_n147 ) );
  NAND2_X1 u1_u9_u4_U22 (.A1( u1_u9_u4_n119 ) , .A2( u1_u9_u4_n120 ) , .ZN( u1_u9_u4_n130 ) );
  NAND2_X1 u1_u9_u4_U23 (.ZN( u1_u9_u4_n117 ) , .A2( u1_u9_u4_n118 ) , .A1( u1_u9_u4_n148 ) );
  NAND2_X1 u1_u9_u4_U24 (.ZN( u1_u9_u4_n129 ) , .A1( u1_u9_u4_n134 ) , .A2( u1_u9_u4_n148 ) );
  AND3_X1 u1_u9_u4_U25 (.A1( u1_u9_u4_n119 ) , .A2( u1_u9_u4_n143 ) , .A3( u1_u9_u4_n154 ) , .ZN( u1_u9_u4_n161 ) );
  AND2_X1 u1_u9_u4_U26 (.A1( u1_u9_u4_n145 ) , .A2( u1_u9_u4_n147 ) , .ZN( u1_u9_u4_n159 ) );
  OR3_X1 u1_u9_u4_U27 (.A3( u1_u9_u4_n114 ) , .A2( u1_u9_u4_n115 ) , .A1( u1_u9_u4_n116 ) , .ZN( u1_u9_u4_n136 ) );
  AOI21_X1 u1_u9_u4_U28 (.A( u1_u9_u4_n113 ) , .ZN( u1_u9_u4_n116 ) , .B2( u1_u9_u4_n173 ) , .B1( u1_u9_u4_n174 ) );
  AOI21_X1 u1_u9_u4_U29 (.ZN( u1_u9_u4_n115 ) , .B2( u1_u9_u4_n145 ) , .B1( u1_u9_u4_n146 ) , .A( u1_u9_u4_n156 ) );
  NOR2_X1 u1_u9_u4_U3 (.ZN( u1_u9_u4_n121 ) , .A1( u1_u9_u4_n181 ) , .A2( u1_u9_u4_n182 ) );
  OAI22_X1 u1_u9_u4_U30 (.ZN( u1_u9_u4_n114 ) , .A2( u1_u9_u4_n121 ) , .B1( u1_u9_u4_n160 ) , .B2( u1_u9_u4_n170 ) , .A1( u1_u9_u4_n171 ) );
  INV_X1 u1_u9_u4_U31 (.A( u1_u9_u4_n158 ) , .ZN( u1_u9_u4_n182 ) );
  INV_X1 u1_u9_u4_U32 (.ZN( u1_u9_u4_n181 ) , .A( u1_u9_u4_n96 ) );
  INV_X1 u1_u9_u4_U33 (.A( u1_u9_u4_n144 ) , .ZN( u1_u9_u4_n179 ) );
  INV_X1 u1_u9_u4_U34 (.A( u1_u9_u4_n157 ) , .ZN( u1_u9_u4_n178 ) );
  NAND2_X1 u1_u9_u4_U35 (.A2( u1_u9_u4_n154 ) , .A1( u1_u9_u4_n96 ) , .ZN( u1_u9_u4_n97 ) );
  INV_X1 u1_u9_u4_U36 (.ZN( u1_u9_u4_n186 ) , .A( u1_u9_u4_n95 ) );
  OAI221_X1 u1_u9_u4_U37 (.C1( u1_u9_u4_n134 ) , .B1( u1_u9_u4_n158 ) , .B2( u1_u9_u4_n171 ) , .C2( u1_u9_u4_n173 ) , .A( u1_u9_u4_n94 ) , .ZN( u1_u9_u4_n95 ) );
  AOI222_X1 u1_u9_u4_U38 (.B2( u1_u9_u4_n132 ) , .A1( u1_u9_u4_n138 ) , .C2( u1_u9_u4_n175 ) , .A2( u1_u9_u4_n179 ) , .C1( u1_u9_u4_n181 ) , .B1( u1_u9_u4_n185 ) , .ZN( u1_u9_u4_n94 ) );
  INV_X1 u1_u9_u4_U39 (.A( u1_u9_u4_n113 ) , .ZN( u1_u9_u4_n185 ) );
  INV_X1 u1_u9_u4_U4 (.A( u1_u9_u4_n117 ) , .ZN( u1_u9_u4_n184 ) );
  INV_X1 u1_u9_u4_U40 (.A( u1_u9_u4_n143 ) , .ZN( u1_u9_u4_n183 ) );
  NOR2_X1 u1_u9_u4_U41 (.ZN( u1_u9_u4_n138 ) , .A1( u1_u9_u4_n168 ) , .A2( u1_u9_u4_n169 ) );
  NOR2_X1 u1_u9_u4_U42 (.A1( u1_u9_u4_n150 ) , .A2( u1_u9_u4_n152 ) , .ZN( u1_u9_u4_n153 ) );
  NOR2_X1 u1_u9_u4_U43 (.A2( u1_u9_u4_n128 ) , .A1( u1_u9_u4_n138 ) , .ZN( u1_u9_u4_n156 ) );
  AOI22_X1 u1_u9_u4_U44 (.B2( u1_u9_u4_n122 ) , .A1( u1_u9_u4_n123 ) , .ZN( u1_u9_u4_n124 ) , .B1( u1_u9_u4_n128 ) , .A2( u1_u9_u4_n172 ) );
  INV_X1 u1_u9_u4_U45 (.A( u1_u9_u4_n153 ) , .ZN( u1_u9_u4_n172 ) );
  NAND2_X1 u1_u9_u4_U46 (.A2( u1_u9_u4_n120 ) , .ZN( u1_u9_u4_n123 ) , .A1( u1_u9_u4_n161 ) );
  AOI22_X1 u1_u9_u4_U47 (.B2( u1_u9_u4_n132 ) , .A2( u1_u9_u4_n133 ) , .ZN( u1_u9_u4_n140 ) , .A1( u1_u9_u4_n150 ) , .B1( u1_u9_u4_n179 ) );
  NAND2_X1 u1_u9_u4_U48 (.ZN( u1_u9_u4_n133 ) , .A2( u1_u9_u4_n146 ) , .A1( u1_u9_u4_n154 ) );
  NAND2_X1 u1_u9_u4_U49 (.A1( u1_u9_u4_n103 ) , .ZN( u1_u9_u4_n154 ) , .A2( u1_u9_u4_n98 ) );
  NOR4_X1 u1_u9_u4_U5 (.A4( u1_u9_u4_n106 ) , .A3( u1_u9_u4_n107 ) , .A2( u1_u9_u4_n108 ) , .A1( u1_u9_u4_n109 ) , .ZN( u1_u9_u4_n110 ) );
  NAND2_X1 u1_u9_u4_U50 (.A1( u1_u9_u4_n101 ) , .ZN( u1_u9_u4_n158 ) , .A2( u1_u9_u4_n99 ) );
  AOI21_X1 u1_u9_u4_U51 (.ZN( u1_u9_u4_n127 ) , .A( u1_u9_u4_n136 ) , .B2( u1_u9_u4_n150 ) , .B1( u1_u9_u4_n180 ) );
  INV_X1 u1_u9_u4_U52 (.A( u1_u9_u4_n160 ) , .ZN( u1_u9_u4_n180 ) );
  NAND2_X1 u1_u9_u4_U53 (.A2( u1_u9_u4_n104 ) , .A1( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n146 ) );
  NAND2_X1 u1_u9_u4_U54 (.A2( u1_u9_u4_n101 ) , .A1( u1_u9_u4_n102 ) , .ZN( u1_u9_u4_n160 ) );
  NAND2_X1 u1_u9_u4_U55 (.ZN( u1_u9_u4_n134 ) , .A1( u1_u9_u4_n98 ) , .A2( u1_u9_u4_n99 ) );
  NAND2_X1 u1_u9_u4_U56 (.A1( u1_u9_u4_n103 ) , .A2( u1_u9_u4_n104 ) , .ZN( u1_u9_u4_n143 ) );
  NAND2_X1 u1_u9_u4_U57 (.A2( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n145 ) , .A1( u1_u9_u4_n98 ) );
  NAND2_X1 u1_u9_u4_U58 (.A1( u1_u9_u4_n100 ) , .A2( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n120 ) );
  NAND2_X1 u1_u9_u4_U59 (.A1( u1_u9_u4_n102 ) , .A2( u1_u9_u4_n104 ) , .ZN( u1_u9_u4_n148 ) );
  AOI21_X1 u1_u9_u4_U6 (.ZN( u1_u9_u4_n106 ) , .B2( u1_u9_u4_n146 ) , .B1( u1_u9_u4_n158 ) , .A( u1_u9_u4_n170 ) );
  NAND2_X1 u1_u9_u4_U60 (.A2( u1_u9_u4_n100 ) , .A1( u1_u9_u4_n103 ) , .ZN( u1_u9_u4_n157 ) );
  INV_X1 u1_u9_u4_U61 (.A( u1_u9_u4_n150 ) , .ZN( u1_u9_u4_n173 ) );
  INV_X1 u1_u9_u4_U62 (.A( u1_u9_u4_n152 ) , .ZN( u1_u9_u4_n171 ) );
  NAND2_X1 u1_u9_u4_U63 (.A1( u1_u9_u4_n100 ) , .ZN( u1_u9_u4_n118 ) , .A2( u1_u9_u4_n99 ) );
  NAND2_X1 u1_u9_u4_U64 (.A2( u1_u9_u4_n100 ) , .A1( u1_u9_u4_n102 ) , .ZN( u1_u9_u4_n144 ) );
  NAND2_X1 u1_u9_u4_U65 (.A2( u1_u9_u4_n101 ) , .A1( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n96 ) );
  INV_X1 u1_u9_u4_U66 (.A( u1_u9_u4_n128 ) , .ZN( u1_u9_u4_n174 ) );
  NAND2_X1 u1_u9_u4_U67 (.A2( u1_u9_u4_n102 ) , .ZN( u1_u9_u4_n119 ) , .A1( u1_u9_u4_n98 ) );
  NAND2_X1 u1_u9_u4_U68 (.A2( u1_u9_u4_n101 ) , .A1( u1_u9_u4_n103 ) , .ZN( u1_u9_u4_n147 ) );
  NAND2_X1 u1_u9_u4_U69 (.A2( u1_u9_u4_n104 ) , .ZN( u1_u9_u4_n113 ) , .A1( u1_u9_u4_n99 ) );
  AOI21_X1 u1_u9_u4_U7 (.ZN( u1_u9_u4_n108 ) , .B2( u1_u9_u4_n134 ) , .B1( u1_u9_u4_n155 ) , .A( u1_u9_u4_n156 ) );
  NOR2_X1 u1_u9_u4_U70 (.A2( u1_u9_X_28 ) , .ZN( u1_u9_u4_n150 ) , .A1( u1_u9_u4_n168 ) );
  NOR2_X1 u1_u9_u4_U71 (.A2( u1_u9_X_29 ) , .ZN( u1_u9_u4_n152 ) , .A1( u1_u9_u4_n169 ) );
  NOR2_X1 u1_u9_u4_U72 (.A2( u1_u9_X_30 ) , .ZN( u1_u9_u4_n105 ) , .A1( u1_u9_u4_n176 ) );
  NOR2_X1 u1_u9_u4_U73 (.A2( u1_u9_X_26 ) , .ZN( u1_u9_u4_n100 ) , .A1( u1_u9_u4_n177 ) );
  NOR2_X1 u1_u9_u4_U74 (.A2( u1_u9_X_28 ) , .A1( u1_u9_X_29 ) , .ZN( u1_u9_u4_n128 ) );
  NOR2_X1 u1_u9_u4_U75 (.A2( u1_u9_X_27 ) , .A1( u1_u9_X_30 ) , .ZN( u1_u9_u4_n102 ) );
  NOR2_X1 u1_u9_u4_U76 (.A2( u1_u9_X_25 ) , .A1( u1_u9_X_26 ) , .ZN( u1_u9_u4_n98 ) );
  AND2_X1 u1_u9_u4_U77 (.A2( u1_u9_X_25 ) , .A1( u1_u9_X_26 ) , .ZN( u1_u9_u4_n104 ) );
  AND2_X1 u1_u9_u4_U78 (.A1( u1_u9_X_30 ) , .A2( u1_u9_u4_n176 ) , .ZN( u1_u9_u4_n99 ) );
  AND2_X1 u1_u9_u4_U79 (.A1( u1_u9_X_26 ) , .ZN( u1_u9_u4_n101 ) , .A2( u1_u9_u4_n177 ) );
  AOI21_X1 u1_u9_u4_U8 (.ZN( u1_u9_u4_n109 ) , .A( u1_u9_u4_n153 ) , .B1( u1_u9_u4_n159 ) , .B2( u1_u9_u4_n184 ) );
  AND2_X1 u1_u9_u4_U80 (.A1( u1_u9_X_27 ) , .A2( u1_u9_X_30 ) , .ZN( u1_u9_u4_n103 ) );
  INV_X1 u1_u9_u4_U81 (.A( u1_u9_X_28 ) , .ZN( u1_u9_u4_n169 ) );
  INV_X1 u1_u9_u4_U82 (.A( u1_u9_X_29 ) , .ZN( u1_u9_u4_n168 ) );
  INV_X1 u1_u9_u4_U83 (.A( u1_u9_X_25 ) , .ZN( u1_u9_u4_n177 ) );
  INV_X1 u1_u9_u4_U84 (.A( u1_u9_X_27 ) , .ZN( u1_u9_u4_n176 ) );
  NAND4_X1 u1_u9_u4_U85 (.ZN( u1_out9_25 ) , .A4( u1_u9_u4_n139 ) , .A3( u1_u9_u4_n140 ) , .A2( u1_u9_u4_n141 ) , .A1( u1_u9_u4_n142 ) );
  OAI21_X1 u1_u9_u4_U86 (.A( u1_u9_u4_n128 ) , .B2( u1_u9_u4_n129 ) , .B1( u1_u9_u4_n130 ) , .ZN( u1_u9_u4_n142 ) );
  OAI21_X1 u1_u9_u4_U87 (.B2( u1_u9_u4_n131 ) , .ZN( u1_u9_u4_n141 ) , .A( u1_u9_u4_n175 ) , .B1( u1_u9_u4_n183 ) );
  NAND4_X1 u1_u9_u4_U88 (.ZN( u1_out9_14 ) , .A4( u1_u9_u4_n124 ) , .A3( u1_u9_u4_n125 ) , .A2( u1_u9_u4_n126 ) , .A1( u1_u9_u4_n127 ) );
  AOI22_X1 u1_u9_u4_U89 (.B2( u1_u9_u4_n117 ) , .ZN( u1_u9_u4_n126 ) , .A1( u1_u9_u4_n129 ) , .B1( u1_u9_u4_n152 ) , .A2( u1_u9_u4_n175 ) );
  AOI211_X1 u1_u9_u4_U9 (.B( u1_u9_u4_n136 ) , .A( u1_u9_u4_n137 ) , .C2( u1_u9_u4_n138 ) , .ZN( u1_u9_u4_n139 ) , .C1( u1_u9_u4_n182 ) );
  AOI22_X1 u1_u9_u4_U90 (.ZN( u1_u9_u4_n125 ) , .B2( u1_u9_u4_n131 ) , .A2( u1_u9_u4_n132 ) , .B1( u1_u9_u4_n138 ) , .A1( u1_u9_u4_n178 ) );
  NAND4_X1 u1_u9_u4_U91 (.ZN( u1_out9_8 ) , .A4( u1_u9_u4_n110 ) , .A3( u1_u9_u4_n111 ) , .A2( u1_u9_u4_n112 ) , .A1( u1_u9_u4_n186 ) );
  NAND2_X1 u1_u9_u4_U92 (.ZN( u1_u9_u4_n112 ) , .A2( u1_u9_u4_n130 ) , .A1( u1_u9_u4_n150 ) );
  AOI22_X1 u1_u9_u4_U93 (.ZN( u1_u9_u4_n111 ) , .B2( u1_u9_u4_n132 ) , .A1( u1_u9_u4_n152 ) , .B1( u1_u9_u4_n178 ) , .A2( u1_u9_u4_n97 ) );
  AOI22_X1 u1_u9_u4_U94 (.B2( u1_u9_u4_n149 ) , .B1( u1_u9_u4_n150 ) , .A2( u1_u9_u4_n151 ) , .A1( u1_u9_u4_n152 ) , .ZN( u1_u9_u4_n167 ) );
  NOR4_X1 u1_u9_u4_U95 (.A4( u1_u9_u4_n162 ) , .A3( u1_u9_u4_n163 ) , .A2( u1_u9_u4_n164 ) , .A1( u1_u9_u4_n165 ) , .ZN( u1_u9_u4_n166 ) );
  NAND3_X1 u1_u9_u4_U96 (.ZN( u1_out9_3 ) , .A3( u1_u9_u4_n166 ) , .A1( u1_u9_u4_n167 ) , .A2( u1_u9_u4_n186 ) );
  NAND3_X1 u1_u9_u4_U97 (.A3( u1_u9_u4_n146 ) , .A2( u1_u9_u4_n147 ) , .A1( u1_u9_u4_n148 ) , .ZN( u1_u9_u4_n149 ) );
  NAND3_X1 u1_u9_u4_U98 (.A3( u1_u9_u4_n143 ) , .A2( u1_u9_u4_n144 ) , .A1( u1_u9_u4_n145 ) , .ZN( u1_u9_u4_n151 ) );
  NAND3_X1 u1_u9_u4_U99 (.A3( u1_u9_u4_n121 ) , .ZN( u1_u9_u4_n122 ) , .A2( u1_u9_u4_n144 ) , .A1( u1_u9_u4_n154 ) );
  INV_X1 u1_uk_U105 (.ZN( u1_K11_5 ) , .A( u1_uk_n496 ) );
  INV_X1 u1_uk_U1129 (.ZN( u1_K11_8 ) , .A( u1_uk_n501 ) );
  INV_X1 u1_uk_U1139 (.ZN( u1_K11_30 ) , .A( u1_uk_n421 ) );
  INV_X1 u1_uk_U226 (.ZN( u1_K11_31 ) , .A( u1_uk_n437 ) );
  INV_X1 u1_uk_U353 (.ZN( u1_K4_4 ) , .A( u1_uk_n1067 ) );
  INV_X1 u1_uk_U461 (.ZN( u1_K9_33 ) , .A( u1_uk_n1162 ) );
  INV_X1 u1_uk_U608 (.ZN( u1_K5_22 ) , .A( u1_uk_n1074 ) );
  INV_X1 u1_uk_U69 (.ZN( u1_K11_34 ) , .A( u1_uk_n443 ) );
  INV_X1 u1_uk_U707 (.ZN( u1_K4_3 ) , .A( u1_uk_n1065 ) );
  INV_X1 u1_uk_U76 (.ZN( u1_K14_34 ) , .A( u1_uk_n955 ) );
  INV_X1 u1_uk_U796 (.ZN( u1_K7_27 ) , .A( u1_uk_n1115 ) );
  XOR2_X1 u2_U315 (.B( u2_L6_26 ) , .Z( u2_N249 ) , .A( u2_out7_26 ) );
  XOR2_X1 u2_U321 (.B( u2_L6_20 ) , .Z( u2_N243 ) , .A( u2_out7_20 ) );
  XOR2_X1 u2_U332 (.B( u2_L6_10 ) , .Z( u2_N233 ) , .A( u2_out7_10 ) );
  XOR2_X1 u2_U342 (.B( u2_L6_1 ) , .Z( u2_N224 ) , .A( u2_out7_1 ) );
  XOR2_X1 u2_u7_U33 (.B( u2_K8_24 ) , .A( u2_R6_17 ) , .Z( u2_u7_X_24 ) );
  XOR2_X1 u2_u7_U34 (.B( u2_K8_23 ) , .A( u2_R6_16 ) , .Z( u2_u7_X_23 ) );
  XOR2_X1 u2_u7_U35 (.B( u2_K8_22 ) , .A( u2_R6_15 ) , .Z( u2_u7_X_22 ) );
  XOR2_X1 u2_u7_U36 (.B( u2_K8_21 ) , .A( u2_R6_14 ) , .Z( u2_u7_X_21 ) );
  XOR2_X1 u2_u7_U37 (.B( u2_K8_20 ) , .A( u2_R6_13 ) , .Z( u2_u7_X_20 ) );
  XOR2_X1 u2_u7_U39 (.B( u2_K8_19 ) , .A( u2_R6_12 ) , .Z( u2_u7_X_19 ) );
  OAI22_X1 u2_u7_u3_U10 (.B1( u2_u7_u3_n113 ) , .A2( u2_u7_u3_n135 ) , .A1( u2_u7_u3_n150 ) , .B2( u2_u7_u3_n164 ) , .ZN( u2_u7_u3_n98 ) );
  OAI211_X1 u2_u7_u3_U11 (.B( u2_u7_u3_n106 ) , .ZN( u2_u7_u3_n119 ) , .C2( u2_u7_u3_n128 ) , .C1( u2_u7_u3_n167 ) , .A( u2_u7_u3_n181 ) );
  AOI221_X1 u2_u7_u3_U12 (.C1( u2_u7_u3_n105 ) , .ZN( u2_u7_u3_n106 ) , .A( u2_u7_u3_n131 ) , .B2( u2_u7_u3_n132 ) , .C2( u2_u7_u3_n133 ) , .B1( u2_u7_u3_n169 ) );
  INV_X1 u2_u7_u3_U13 (.ZN( u2_u7_u3_n181 ) , .A( u2_u7_u3_n98 ) );
  NAND2_X1 u2_u7_u3_U14 (.ZN( u2_u7_u3_n105 ) , .A2( u2_u7_u3_n130 ) , .A1( u2_u7_u3_n155 ) );
  AOI22_X1 u2_u7_u3_U15 (.B1( u2_u7_u3_n115 ) , .A2( u2_u7_u3_n116 ) , .ZN( u2_u7_u3_n123 ) , .B2( u2_u7_u3_n133 ) , .A1( u2_u7_u3_n169 ) );
  NAND2_X1 u2_u7_u3_U16 (.ZN( u2_u7_u3_n116 ) , .A2( u2_u7_u3_n151 ) , .A1( u2_u7_u3_n182 ) );
  NOR2_X1 u2_u7_u3_U17 (.ZN( u2_u7_u3_n126 ) , .A2( u2_u7_u3_n150 ) , .A1( u2_u7_u3_n164 ) );
  AOI21_X1 u2_u7_u3_U18 (.ZN( u2_u7_u3_n112 ) , .B2( u2_u7_u3_n146 ) , .B1( u2_u7_u3_n155 ) , .A( u2_u7_u3_n167 ) );
  NAND2_X1 u2_u7_u3_U19 (.A1( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n142 ) , .A2( u2_u7_u3_n164 ) );
  NAND2_X1 u2_u7_u3_U20 (.ZN( u2_u7_u3_n132 ) , .A2( u2_u7_u3_n152 ) , .A1( u2_u7_u3_n156 ) );
  AND2_X1 u2_u7_u3_U21 (.A2( u2_u7_u3_n113 ) , .A1( u2_u7_u3_n114 ) , .ZN( u2_u7_u3_n151 ) );
  INV_X1 u2_u7_u3_U22 (.A( u2_u7_u3_n133 ) , .ZN( u2_u7_u3_n165 ) );
  INV_X1 u2_u7_u3_U23 (.A( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n170 ) );
  NAND2_X1 u2_u7_u3_U24 (.A1( u2_u7_u3_n107 ) , .A2( u2_u7_u3_n108 ) , .ZN( u2_u7_u3_n140 ) );
  NAND2_X1 u2_u7_u3_U25 (.ZN( u2_u7_u3_n117 ) , .A1( u2_u7_u3_n124 ) , .A2( u2_u7_u3_n148 ) );
  NAND2_X1 u2_u7_u3_U26 (.ZN( u2_u7_u3_n143 ) , .A1( u2_u7_u3_n165 ) , .A2( u2_u7_u3_n167 ) );
  INV_X1 u2_u7_u3_U27 (.A( u2_u7_u3_n130 ) , .ZN( u2_u7_u3_n177 ) );
  INV_X1 u2_u7_u3_U28 (.A( u2_u7_u3_n128 ) , .ZN( u2_u7_u3_n176 ) );
  INV_X1 u2_u7_u3_U29 (.A( u2_u7_u3_n155 ) , .ZN( u2_u7_u3_n174 ) );
  INV_X1 u2_u7_u3_U3 (.A( u2_u7_u3_n129 ) , .ZN( u2_u7_u3_n183 ) );
  INV_X1 u2_u7_u3_U30 (.A( u2_u7_u3_n139 ) , .ZN( u2_u7_u3_n185 ) );
  NOR2_X1 u2_u7_u3_U31 (.ZN( u2_u7_u3_n135 ) , .A2( u2_u7_u3_n141 ) , .A1( u2_u7_u3_n169 ) );
  OAI222_X1 u2_u7_u3_U32 (.C2( u2_u7_u3_n107 ) , .A2( u2_u7_u3_n108 ) , .B1( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n138 ) , .B2( u2_u7_u3_n146 ) , .C1( u2_u7_u3_n154 ) , .A1( u2_u7_u3_n164 ) );
  NOR4_X1 u2_u7_u3_U33 (.A4( u2_u7_u3_n157 ) , .A3( u2_u7_u3_n158 ) , .A2( u2_u7_u3_n159 ) , .A1( u2_u7_u3_n160 ) , .ZN( u2_u7_u3_n161 ) );
  AOI21_X1 u2_u7_u3_U34 (.B2( u2_u7_u3_n152 ) , .B1( u2_u7_u3_n153 ) , .ZN( u2_u7_u3_n158 ) , .A( u2_u7_u3_n164 ) );
  AOI21_X1 u2_u7_u3_U35 (.A( u2_u7_u3_n154 ) , .B2( u2_u7_u3_n155 ) , .B1( u2_u7_u3_n156 ) , .ZN( u2_u7_u3_n157 ) );
  AOI21_X1 u2_u7_u3_U36 (.A( u2_u7_u3_n149 ) , .B2( u2_u7_u3_n150 ) , .B1( u2_u7_u3_n151 ) , .ZN( u2_u7_u3_n159 ) );
  AOI211_X1 u2_u7_u3_U37 (.ZN( u2_u7_u3_n109 ) , .A( u2_u7_u3_n119 ) , .C2( u2_u7_u3_n129 ) , .B( u2_u7_u3_n138 ) , .C1( u2_u7_u3_n141 ) );
  AOI211_X1 u2_u7_u3_U38 (.B( u2_u7_u3_n119 ) , .A( u2_u7_u3_n120 ) , .C2( u2_u7_u3_n121 ) , .ZN( u2_u7_u3_n122 ) , .C1( u2_u7_u3_n179 ) );
  INV_X1 u2_u7_u3_U39 (.A( u2_u7_u3_n156 ) , .ZN( u2_u7_u3_n179 ) );
  INV_X1 u2_u7_u3_U4 (.A( u2_u7_u3_n140 ) , .ZN( u2_u7_u3_n182 ) );
  OAI22_X1 u2_u7_u3_U40 (.B1( u2_u7_u3_n118 ) , .ZN( u2_u7_u3_n120 ) , .A1( u2_u7_u3_n135 ) , .B2( u2_u7_u3_n154 ) , .A2( u2_u7_u3_n178 ) );
  AND3_X1 u2_u7_u3_U41 (.ZN( u2_u7_u3_n118 ) , .A2( u2_u7_u3_n124 ) , .A1( u2_u7_u3_n144 ) , .A3( u2_u7_u3_n152 ) );
  INV_X1 u2_u7_u3_U42 (.A( u2_u7_u3_n121 ) , .ZN( u2_u7_u3_n164 ) );
  NAND2_X1 u2_u7_u3_U43 (.ZN( u2_u7_u3_n133 ) , .A1( u2_u7_u3_n154 ) , .A2( u2_u7_u3_n164 ) );
  OAI211_X1 u2_u7_u3_U44 (.B( u2_u7_u3_n127 ) , .ZN( u2_u7_u3_n139 ) , .C1( u2_u7_u3_n150 ) , .C2( u2_u7_u3_n154 ) , .A( u2_u7_u3_n184 ) );
  INV_X1 u2_u7_u3_U45 (.A( u2_u7_u3_n125 ) , .ZN( u2_u7_u3_n184 ) );
  AOI221_X1 u2_u7_u3_U46 (.A( u2_u7_u3_n126 ) , .ZN( u2_u7_u3_n127 ) , .C2( u2_u7_u3_n132 ) , .C1( u2_u7_u3_n169 ) , .B2( u2_u7_u3_n170 ) , .B1( u2_u7_u3_n174 ) );
  OAI22_X1 u2_u7_u3_U47 (.A1( u2_u7_u3_n124 ) , .ZN( u2_u7_u3_n125 ) , .B2( u2_u7_u3_n145 ) , .A2( u2_u7_u3_n165 ) , .B1( u2_u7_u3_n167 ) );
  NOR2_X1 u2_u7_u3_U48 (.A1( u2_u7_u3_n113 ) , .ZN( u2_u7_u3_n131 ) , .A2( u2_u7_u3_n154 ) );
  NAND2_X1 u2_u7_u3_U49 (.A1( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n150 ) , .A2( u2_u7_u3_n99 ) );
  INV_X1 u2_u7_u3_U5 (.A( u2_u7_u3_n117 ) , .ZN( u2_u7_u3_n178 ) );
  NAND2_X1 u2_u7_u3_U50 (.A2( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n155 ) , .A1( u2_u7_u3_n97 ) );
  INV_X1 u2_u7_u3_U51 (.A( u2_u7_u3_n141 ) , .ZN( u2_u7_u3_n167 ) );
  AOI21_X1 u2_u7_u3_U52 (.B2( u2_u7_u3_n114 ) , .B1( u2_u7_u3_n146 ) , .A( u2_u7_u3_n154 ) , .ZN( u2_u7_u3_n94 ) );
  AOI21_X1 u2_u7_u3_U53 (.ZN( u2_u7_u3_n110 ) , .B2( u2_u7_u3_n142 ) , .B1( u2_u7_u3_n186 ) , .A( u2_u7_u3_n95 ) );
  INV_X1 u2_u7_u3_U54 (.A( u2_u7_u3_n145 ) , .ZN( u2_u7_u3_n186 ) );
  AOI21_X1 u2_u7_u3_U55 (.B1( u2_u7_u3_n124 ) , .A( u2_u7_u3_n149 ) , .B2( u2_u7_u3_n155 ) , .ZN( u2_u7_u3_n95 ) );
  INV_X1 u2_u7_u3_U56 (.A( u2_u7_u3_n149 ) , .ZN( u2_u7_u3_n169 ) );
  NAND2_X1 u2_u7_u3_U57 (.ZN( u2_u7_u3_n124 ) , .A1( u2_u7_u3_n96 ) , .A2( u2_u7_u3_n97 ) );
  NAND2_X1 u2_u7_u3_U58 (.A2( u2_u7_u3_n100 ) , .ZN( u2_u7_u3_n146 ) , .A1( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U59 (.A1( u2_u7_u3_n101 ) , .ZN( u2_u7_u3_n145 ) , .A2( u2_u7_u3_n99 ) );
  AOI221_X1 u2_u7_u3_U6 (.A( u2_u7_u3_n131 ) , .C2( u2_u7_u3_n132 ) , .C1( u2_u7_u3_n133 ) , .ZN( u2_u7_u3_n134 ) , .B1( u2_u7_u3_n143 ) , .B2( u2_u7_u3_n177 ) );
  NAND2_X1 u2_u7_u3_U60 (.A1( u2_u7_u3_n100 ) , .ZN( u2_u7_u3_n156 ) , .A2( u2_u7_u3_n99 ) );
  NAND2_X1 u2_u7_u3_U61 (.A2( u2_u7_u3_n101 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n148 ) );
  NAND2_X1 u2_u7_u3_U62 (.A1( u2_u7_u3_n100 ) , .A2( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n128 ) );
  NAND2_X1 u2_u7_u3_U63 (.A2( u2_u7_u3_n101 ) , .A1( u2_u7_u3_n102 ) , .ZN( u2_u7_u3_n152 ) );
  NAND2_X1 u2_u7_u3_U64 (.A2( u2_u7_u3_n101 ) , .ZN( u2_u7_u3_n114 ) , .A1( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U65 (.ZN( u2_u7_u3_n107 ) , .A1( u2_u7_u3_n97 ) , .A2( u2_u7_u3_n99 ) );
  NAND2_X1 u2_u7_u3_U66 (.A2( u2_u7_u3_n100 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n113 ) );
  NAND2_X1 u2_u7_u3_U67 (.A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n153 ) , .A2( u2_u7_u3_n97 ) );
  NAND2_X1 u2_u7_u3_U68 (.A2( u2_u7_u3_n103 ) , .A1( u2_u7_u3_n104 ) , .ZN( u2_u7_u3_n130 ) );
  NAND2_X1 u2_u7_u3_U69 (.A2( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n144 ) , .A1( u2_u7_u3_n96 ) );
  OAI22_X1 u2_u7_u3_U7 (.B2( u2_u7_u3_n147 ) , .A2( u2_u7_u3_n148 ) , .ZN( u2_u7_u3_n160 ) , .B1( u2_u7_u3_n165 ) , .A1( u2_u7_u3_n168 ) );
  NAND2_X1 u2_u7_u3_U70 (.A1( u2_u7_u3_n102 ) , .A2( u2_u7_u3_n103 ) , .ZN( u2_u7_u3_n108 ) );
  NOR2_X1 u2_u7_u3_U71 (.A2( u2_u7_X_19 ) , .A1( u2_u7_X_20 ) , .ZN( u2_u7_u3_n99 ) );
  NOR2_X1 u2_u7_u3_U72 (.A2( u2_u7_X_21 ) , .A1( u2_u7_X_24 ) , .ZN( u2_u7_u3_n103 ) );
  NOR2_X1 u2_u7_u3_U73 (.A2( u2_u7_X_24 ) , .A1( u2_u7_u3_n171 ) , .ZN( u2_u7_u3_n97 ) );
  NOR2_X1 u2_u7_u3_U74 (.A2( u2_u7_X_23 ) , .ZN( u2_u7_u3_n141 ) , .A1( u2_u7_u3_n166 ) );
  NOR2_X1 u2_u7_u3_U75 (.A2( u2_u7_X_19 ) , .A1( u2_u7_u3_n172 ) , .ZN( u2_u7_u3_n96 ) );
  NAND2_X1 u2_u7_u3_U76 (.A1( u2_u7_X_22 ) , .A2( u2_u7_X_23 ) , .ZN( u2_u7_u3_n154 ) );
  NAND2_X1 u2_u7_u3_U77 (.A1( u2_u7_X_23 ) , .ZN( u2_u7_u3_n149 ) , .A2( u2_u7_u3_n166 ) );
  NOR2_X1 u2_u7_u3_U78 (.A2( u2_u7_X_22 ) , .A1( u2_u7_X_23 ) , .ZN( u2_u7_u3_n121 ) );
  AND2_X1 u2_u7_u3_U79 (.A1( u2_u7_X_24 ) , .ZN( u2_u7_u3_n101 ) , .A2( u2_u7_u3_n171 ) );
  AND3_X1 u2_u7_u3_U8 (.A3( u2_u7_u3_n144 ) , .A2( u2_u7_u3_n145 ) , .A1( u2_u7_u3_n146 ) , .ZN( u2_u7_u3_n147 ) );
  AND2_X1 u2_u7_u3_U80 (.A1( u2_u7_X_19 ) , .ZN( u2_u7_u3_n102 ) , .A2( u2_u7_u3_n172 ) );
  AND2_X1 u2_u7_u3_U81 (.A1( u2_u7_X_21 ) , .A2( u2_u7_X_24 ) , .ZN( u2_u7_u3_n100 ) );
  AND2_X1 u2_u7_u3_U82 (.A2( u2_u7_X_19 ) , .A1( u2_u7_X_20 ) , .ZN( u2_u7_u3_n104 ) );
  INV_X1 u2_u7_u3_U83 (.A( u2_u7_X_22 ) , .ZN( u2_u7_u3_n166 ) );
  INV_X1 u2_u7_u3_U84 (.A( u2_u7_X_21 ) , .ZN( u2_u7_u3_n171 ) );
  INV_X1 u2_u7_u3_U85 (.A( u2_u7_X_20 ) , .ZN( u2_u7_u3_n172 ) );
  OR4_X1 u2_u7_u3_U86 (.ZN( u2_out7_10 ) , .A4( u2_u7_u3_n136 ) , .A3( u2_u7_u3_n137 ) , .A1( u2_u7_u3_n138 ) , .A2( u2_u7_u3_n139 ) );
  OAI222_X1 u2_u7_u3_U87 (.C1( u2_u7_u3_n128 ) , .ZN( u2_u7_u3_n137 ) , .B1( u2_u7_u3_n148 ) , .A2( u2_u7_u3_n150 ) , .B2( u2_u7_u3_n154 ) , .C2( u2_u7_u3_n164 ) , .A1( u2_u7_u3_n167 ) );
  OAI221_X1 u2_u7_u3_U88 (.A( u2_u7_u3_n134 ) , .B2( u2_u7_u3_n135 ) , .ZN( u2_u7_u3_n136 ) , .C1( u2_u7_u3_n149 ) , .B1( u2_u7_u3_n151 ) , .C2( u2_u7_u3_n183 ) );
  NAND4_X1 u2_u7_u3_U89 (.ZN( u2_out7_26 ) , .A4( u2_u7_u3_n109 ) , .A3( u2_u7_u3_n110 ) , .A2( u2_u7_u3_n111 ) , .A1( u2_u7_u3_n173 ) );
  INV_X1 u2_u7_u3_U9 (.A( u2_u7_u3_n143 ) , .ZN( u2_u7_u3_n168 ) );
  INV_X1 u2_u7_u3_U90 (.ZN( u2_u7_u3_n173 ) , .A( u2_u7_u3_n94 ) );
  OAI21_X1 u2_u7_u3_U91 (.ZN( u2_u7_u3_n111 ) , .B2( u2_u7_u3_n117 ) , .A( u2_u7_u3_n133 ) , .B1( u2_u7_u3_n176 ) );
  NAND4_X1 u2_u7_u3_U92 (.ZN( u2_out7_20 ) , .A4( u2_u7_u3_n122 ) , .A3( u2_u7_u3_n123 ) , .A1( u2_u7_u3_n175 ) , .A2( u2_u7_u3_n180 ) );
  INV_X1 u2_u7_u3_U93 (.A( u2_u7_u3_n126 ) , .ZN( u2_u7_u3_n180 ) );
  INV_X1 u2_u7_u3_U94 (.A( u2_u7_u3_n112 ) , .ZN( u2_u7_u3_n175 ) );
  NAND4_X1 u2_u7_u3_U95 (.ZN( u2_out7_1 ) , .A4( u2_u7_u3_n161 ) , .A3( u2_u7_u3_n162 ) , .A2( u2_u7_u3_n163 ) , .A1( u2_u7_u3_n185 ) );
  NAND2_X1 u2_u7_u3_U96 (.ZN( u2_u7_u3_n163 ) , .A2( u2_u7_u3_n170 ) , .A1( u2_u7_u3_n176 ) );
  AOI22_X1 u2_u7_u3_U97 (.B2( u2_u7_u3_n140 ) , .B1( u2_u7_u3_n141 ) , .A2( u2_u7_u3_n142 ) , .ZN( u2_u7_u3_n162 ) , .A1( u2_u7_u3_n177 ) );
  NAND3_X1 u2_u7_u3_U98 (.A1( u2_u7_u3_n114 ) , .ZN( u2_u7_u3_n115 ) , .A2( u2_u7_u3_n145 ) , .A3( u2_u7_u3_n153 ) );
  NAND3_X1 u2_u7_u3_U99 (.ZN( u2_u7_u3_n129 ) , .A2( u2_u7_u3_n144 ) , .A1( u2_u7_u3_n153 ) , .A3( u2_u7_u3_n182 ) );
  OAI22_X1 u2_uk_U159 (.ZN( u2_K8_19 ) , .B2( u2_uk_n1508 ) , .A2( u2_uk_n1515 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U597 (.ZN( u2_K8_22 ) , .B2( u2_uk_n1529 ) , .A2( u2_uk_n1535 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U75 (.ZN( u2_K8_23 ) , .B2( u2_uk_n1513 ) , .A2( u2_uk_n1518 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U819 (.ZN( u2_K8_20 ) , .B2( u2_uk_n1521 ) , .A2( u2_uk_n1527 ) , .A1( u2_uk_n220 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U886 (.ZN( u2_K8_21 ) , .B2( u2_uk_n1522 ) , .A2( u2_uk_n1528 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
endmodule

