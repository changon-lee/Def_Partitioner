module des_des_die_7 ( n116, u0_K11_21, u0_K15_47, u0_K4_24, u0_K4_6, u0_K5_26, u0_K5_28, u0_L13_12, u0_L13_14, 
       u0_L13_15, u0_L13_17, u0_L13_21, u0_L13_22, u0_L13_23, u0_L13_25, u0_L13_27, u0_L13_3, u0_L13_31, 
       u0_L13_32, u0_L13_5, u0_L13_7, u0_L13_8, u0_L13_9, u0_L2_1, u0_L2_10, u0_L2_13, u0_L2_16, 
       u0_L2_17, u0_L2_18, u0_L2_2, u0_L2_20, u0_L2_23, u0_L2_24, u0_L2_26, u0_L2_28, u0_L2_30, 
       u0_L2_31, u0_L2_6, u0_L2_9, u0_L3_14, u0_L3_25, u0_L3_3, u0_L3_8, u0_L9_1, u0_L9_10, 
       u0_L9_16, u0_L9_20, u0_L9_24, u0_L9_26, u0_L9_30, u0_L9_6, u0_R13_1, u0_R13_16, u0_R13_17, 
       u0_R13_18, u0_R13_19, u0_R13_2, u0_R13_20, u0_R13_21, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, 
       u0_R13_28, u0_R13_29, u0_R13_3, u0_R13_30, u0_R13_31, u0_R13_32, u0_R13_4, u0_R13_5, u0_R2_1, 
       u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_2, 
       u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_16, 
       u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_20, u0_R3_21, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, 
       u0_R9_14, u0_R9_15, u0_R9_16, u0_R9_17, u0_R9_8, u0_R9_9, u0_key_r_18, u0_key_r_33, u0_key_r_44, 
       u0_uk_K_r0_52, u0_uk_K_r13_0, u0_uk_K_r13_2, u0_uk_K_r13_22, u0_uk_K_r13_23, u0_uk_K_r13_35, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r2_13, 
       u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, 
       u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_35, u0_uk_K_r9_10, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_27, u0_uk_K_r9_38, u0_uk_K_r9_48, 
       u0_uk_K_r9_5, u0_uk_n1, u0_uk_n10, u0_uk_n100, u0_uk_n1001, u0_uk_n1002, u0_uk_n109, u0_uk_n110, u0_uk_n117, 
       u0_uk_n118, u0_uk_n12, u0_uk_n128, u0_uk_n129, u0_uk_n13, u0_uk_n141, u0_uk_n142, u0_uk_n146, u0_uk_n147, 
       u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, 
       u0_uk_n190, u0_uk_n196, u0_uk_n197, u0_uk_n20, u0_uk_n200, u0_uk_n201, u0_uk_n202, u0_uk_n203, u0_uk_n206, 
       u0_uk_n207, u0_uk_n208, u0_uk_n21, u0_uk_n212, u0_uk_n214, u0_uk_n215, u0_uk_n217, u0_uk_n22, u0_uk_n220, 
       u0_uk_n221, u0_uk_n222, u0_uk_n23, u0_uk_n230, u0_uk_n238, u0_uk_n24, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
       u0_uk_n251, u0_uk_n252, u0_uk_n26, u0_uk_n27, u0_uk_n29, u0_uk_n3, u0_uk_n30, u0_uk_n31, u0_uk_n33, 
       u0_uk_n34, u0_uk_n36, u0_uk_n38, u0_uk_n39, u0_uk_n4, u0_uk_n40, u0_uk_n41, u0_uk_n462, u0_uk_n463, 
       u0_uk_n475, u0_uk_n480, u0_uk_n481, u0_uk_n497, u0_uk_n5, u0_uk_n502, u0_uk_n510, u0_uk_n511, u0_uk_n517, 
       u0_uk_n519, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n534, u0_uk_n535, u0_uk_n536, 
       u0_uk_n6, u0_uk_n60, u0_uk_n8, u0_uk_n813, u0_uk_n83, u0_uk_n834, u0_uk_n839, u0_uk_n9, u0_uk_n916, 
       u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u0_uk_n999, u1_FP_33, u1_FP_36, u1_FP_37, u1_FP_40, 
       u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_46, u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, 
       u1_FP_52, u1_FP_53, u1_FP_56, u1_FP_57, u1_FP_60, u1_FP_61, u1_FP_64, u1_L0_1, u1_L0_10, 
       u1_L0_12, u1_L0_14, u1_L0_15, u1_L0_16, u1_L0_17, u1_L0_20, u1_L0_21, u1_L0_22, u1_L0_23, 
       u1_L0_24, u1_L0_25, u1_L0_26, u1_L0_27, u1_L0_3, u1_L0_30, u1_L0_31, u1_L0_32, u1_L0_5, 
       u1_L0_6, u1_L0_7, u1_L0_8, u1_L0_9, u1_L10_1, u1_L10_10, u1_L10_13, u1_L10_14, u1_L10_16, 
       u1_L10_18, u1_L10_2, u1_L10_20, u1_L10_24, u1_L10_25, u1_L10_26, u1_L10_28, u1_L10_3, u1_L10_30, 
       u1_L10_6, u1_L10_8, u1_L11_1, u1_L11_10, u1_L11_14, u1_L11_17, u1_L11_20, u1_L11_23, u1_L11_25, 
       u1_L11_26, u1_L11_3, u1_L11_31, u1_L11_8, u1_L11_9, u1_L12_12, u1_L12_13, u1_L12_14, u1_L12_15, 
       u1_L12_18, u1_L12_2, u1_L12_21, u1_L12_22, u1_L12_25, u1_L12_27, u1_L12_28, u1_L12_3, u1_L12_32, 
       u1_L12_5, u1_L12_7, u1_L12_8, u1_L13_11, u1_L13_12, u1_L13_15, u1_L13_16, u1_L13_19, u1_L13_21, 
       u1_L13_22, u1_L13_24, u1_L13_27, u1_L13_29, u1_L13_30, u1_L13_32, u1_L13_4, u1_L13_5, u1_L13_6, 
       u1_L13_7, u1_L14_1, u1_L14_10, u1_L14_14, u1_L14_20, u1_L14_25, u1_L14_26, u1_L14_3, u1_L14_8, 
       u1_L1_1, u1_L1_10, u1_L1_15, u1_L1_20, u1_L1_21, u1_L1_26, u1_L1_27, u1_L1_5, u1_L2_1, 
       u1_L2_10, u1_L2_20, u1_L2_26, u1_L3_11, u1_L3_15, u1_L3_19, u1_L3_21, u1_L3_27, u1_L3_29, 
       u1_L3_4, u1_L3_5, u1_L4_1, u1_L4_10, u1_L4_12, u1_L4_16, u1_L4_17, u1_L4_20, u1_L4_22, 
       u1_L4_23, u1_L4_24, u1_L4_26, u1_L4_30, u1_L4_31, u1_L4_32, u1_L4_6, u1_L4_7, u1_L4_9, 
       u1_L5_1, u1_L5_10, u1_L5_16, u1_L5_20, u1_L5_24, u1_L5_26, u1_L5_30, u1_L5_6, u1_L6_12, 
       u1_L6_13, u1_L6_14, u1_L6_16, u1_L6_17, u1_L6_18, u1_L6_2, u1_L6_22, u1_L6_23, u1_L6_24, 
       u1_L6_25, u1_L6_28, u1_L6_3, u1_L6_30, u1_L6_31, u1_L6_32, u1_L6_6, u1_L6_7, u1_L6_8, 
       u1_L6_9, u1_L7_1, u1_L7_10, u1_L7_12, u1_L7_13, u1_L7_15, u1_L7_16, u1_L7_18, u1_L7_2, 
       u1_L7_20, u1_L7_21, u1_L7_22, u1_L7_24, u1_L7_26, u1_L7_27, u1_L7_28, u1_L7_30, u1_L7_32, 
       u1_L7_5, u1_L7_6, u1_L7_7, u1_L8_15, u1_L8_17, u1_L8_21, u1_L8_23, u1_L8_27, u1_L8_31, 
       u1_L8_5, u1_L8_9, u1_L9_12, u1_L9_22, u1_L9_32, u1_L9_7, u1_R0_1, u1_R0_10, u1_R0_11, 
       u1_R0_12, u1_R0_13, u1_R0_14, u1_R0_15, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_2, 
       u1_R0_20, u1_R0_21, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, u1_R0_3, 
       u1_R0_30, u1_R0_31, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_8, u1_R0_9, u1_R10_1, u1_R10_10, 
       u1_R10_11, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_18, u1_R10_19, 
       u1_R10_20, u1_R10_21, u1_R10_24, u1_R10_25, u1_R10_28, u1_R10_29, u1_R10_32, u1_R10_4, u1_R10_5, 
       u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_1, u1_R11_12, u1_R11_13, u1_R11_14, u1_R11_15, 
       u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_20, u1_R11_21, u1_R11_24, u1_R11_25, 
       u1_R11_28, u1_R11_29, u1_R11_3, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_9, u1_R12_1, u1_R12_12, 
       u1_R12_13, u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, u1_R12_20, u1_R12_21, u1_R12_24, u1_R12_25, 
       u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_29, u1_R12_30, u1_R12_31, u1_R12_32, u1_R12_4, u1_R12_5, 
       u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_1, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, 
       u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, 
       u1_R13_27, u1_R13_28, u1_R13_29, u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_4, u1_R13_5, u1_R13_8, 
       u1_R13_9, u1_R1_1, u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, u1_R1_17, u1_R1_20, 
       u1_R1_21, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_30, u1_R1_31, u1_R1_32, u1_R1_4, 
       u1_R1_5, u1_R1_8, u1_R1_9, u1_R2_1, u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, 
       u1_R2_17, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_32, u1_R2_4, u1_R2_5, u1_R2_8, 
       u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_16, u1_R3_17, u1_R3_20, u1_R3_21, u1_R3_22, 
       u1_R3_23, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_30, u1_R3_31, u1_R3_32, u1_R3_5, 
       u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_10, u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, 
       u1_R4_16, u1_R4_17, u1_R4_2, u1_R4_21, u1_R4_24, u1_R4_25, u1_R4_26, u1_R4_27, u1_R4_28, 
       u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_10, 
       u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_14, u1_R5_15, u1_R5_16, u1_R5_17, u1_R5_20, u1_R5_21, 
       u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_8, u1_R5_9, 
       u1_R6_1, u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_16, u1_R6_17, u1_R6_18, u1_R6_19, 
       u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, 
       u1_R6_3, u1_R6_32, u1_R6_4, u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, 
       u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_20, 
       u1_R7_21, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, u1_R7_29, u1_R7_30, u1_R7_31, 
       u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_16, 
       u1_R8_17, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_30, u1_R8_31, 
       u1_R8_32, u1_R8_4, u1_R8_5, u1_R9_1, u1_R9_16, u1_R9_17, u1_R9_24, u1_R9_25, u1_R9_26, 
       u1_R9_27, u1_R9_28, u1_R9_29, u1_R9_32, u1_R9_8, u1_R9_9, u1_desIn_r_1, u1_desIn_r_10, u1_desIn_r_12, 
       u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_16, u1_desIn_r_17, u1_desIn_r_2, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_25, u1_desIn_r_26, 
       u1_desIn_r_28, u1_desIn_r_29, u1_desIn_r_3, u1_desIn_r_31, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_36, u1_desIn_r_37, 
       u1_desIn_r_38, u1_desIn_r_39, u1_desIn_r_4, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_45, u1_desIn_r_47, u1_desIn_r_48, u1_desIn_r_49, 
       u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_52, u1_desIn_r_53, u1_desIn_r_54, u1_desIn_r_55, u1_desIn_r_56, u1_desIn_r_57, u1_desIn_r_59, 
       u1_desIn_r_6, u1_desIn_r_61, u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_8, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, 
       u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, 
       u1_key_r_2, u1_key_r_20, u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, 
       u1_key_r_28, u1_key_r_29, u1_key_r_3, u1_key_r_30, u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, 
       u1_key_r_36, u1_key_r_37, u1_key_r_38, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, 
       u1_key_r_44, u1_key_r_45, u1_key_r_46, u1_key_r_47, u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, 
       u1_key_r_52, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_11, 
       u1_uk_K_r0_13, u1_uk_K_r0_15, u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, u1_uk_K_r0_31, 
       u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, u1_uk_K_r10_10, 
       u1_uk_K_r10_11, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, u1_uk_K_r10_28, 
       u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, 
       u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, u1_uk_K_r11_19, 
       u1_uk_K_r11_20, u1_uk_K_r11_21, u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_33, 
       u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, u1_uk_K_r11_54, 
       u1_uk_K_r11_6, u1_uk_K_r11_7, u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, u1_uk_K_r12_21, 
       u1_uk_K_r12_22, u1_uk_K_r12_25, u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_47, 
       u1_uk_K_r12_7, u1_uk_K_r13_0, u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_25, 
       u1_uk_K_r13_31, u1_uk_K_r13_32, u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, u1_uk_K_r14_10, 
       u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, 
       u1_uk_K_r14_39, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, 
       u1_uk_K_r1_10, u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, u1_uk_K_r1_36, 
       u1_uk_K_r1_41, u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, u1_uk_K_r2_18, 
       u1_uk_K_r2_20, u1_uk_K_r2_21, u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_31, 
       u1_uk_K_r2_33, u1_uk_K_r2_36, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r2_53, 
       u1_uk_K_r2_55, u1_uk_K_r2_6, u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, u1_uk_K_r3_19, 
       u1_uk_K_r3_24, u1_uk_K_r3_29, u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, u1_uk_K_r3_44, 
       u1_uk_K_r3_47, u1_uk_K_r3_51, u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_23, 
       u1_uk_K_r4_27, u1_uk_K_r4_3, u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, u1_uk_K_r4_47, 
       u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_13, 
       u1_uk_K_r5_16, u1_uk_K_r5_17, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, 
       u1_uk_K_r5_35, u1_uk_K_r5_36, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, u1_uk_K_r5_48, 
       u1_uk_K_r5_5, u1_uk_K_r5_51, u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, u1_uk_K_r6_17, 
       u1_uk_K_r6_19, u1_uk_K_r6_21, u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, 
       u1_uk_K_r6_31, u1_uk_K_r6_34, u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r6_7, 
       u1_uk_K_r7_0, u1_uk_K_r7_1, u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, u1_uk_K_r7_23, 
       u1_uk_K_r7_24, u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, u1_uk_K_r7_34, 
       u1_uk_K_r7_37, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, 
       u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, u1_uk_K_r8_2, 
       u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, u1_uk_K_r8_41, 
       u1_uk_K_r8_42, u1_uk_K_r8_43, u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, u1_uk_K_r9_0, 
       u1_uk_K_r9_1, u1_uk_K_r9_10, u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_23, 
       u1_uk_K_r9_25, u1_uk_K_r9_27, u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, u1_uk_K_r9_45, 
       u1_uk_K_r9_48, u1_uk_K_r9_49, u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, u1_uk_n1218, 
       u1_uk_n1219, u1_uk_n1220, u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, 
       u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, 
       u1_uk_n1240, u1_uk_n1241, u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, 
       u1_uk_n1249, u1_uk_n1250, u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, 
       u1_uk_n1259, u1_uk_n1260, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, 
       u1_uk_n1268, u1_uk_n1269, u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, 
       u1_uk_n1277, u1_uk_n1278, u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, 
       u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, 
       u1_uk_n1300, u1_uk_n1303, u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, 
       u1_uk_n1312, u1_uk_n1313, u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, 
       u1_uk_n1321, u1_uk_n1322, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, 
       u1_uk_n1330, u1_uk_n1331, u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, 
       u1_uk_n1340, u1_uk_n1341, u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, 
       u1_uk_n1349, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, 
       u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, 
       u1_uk_n1371, u1_uk_n1372, u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, 
       u1_uk_n1382, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, 
       u1_uk_n1396, u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, 
       u1_uk_n1405, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, 
       u1_uk_n1414, u1_uk_n1415, u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, 
       u1_uk_n1426, u1_uk_n1427, u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, 
       u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, 
       u1_uk_n1448, u1_uk_n1449, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, 
       u1_uk_n1458, u1_uk_n1459, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, 
       u1_uk_n1468, u1_uk_n1469, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, 
       u1_uk_n1478, u1_uk_n1482, u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, 
       u1_uk_n1490, u1_uk_n1491, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, 
       u1_uk_n1501, u1_uk_n1504, u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, 
       u1_uk_n1518, u1_uk_n1520, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, 
       u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, 
       u1_uk_n1541, u1_uk_n1543, u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, 
       u1_uk_n1554, u1_uk_n1555, u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, 
       u1_uk_n1563, u1_uk_n1564, u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, 
       u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, 
       u1_uk_n1588, u1_uk_n1592, u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, 
       u1_uk_n1604, u1_uk_n1605, u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, 
       u1_uk_n1615, u1_uk_n1616, u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, 
       u1_uk_n1625, u1_uk_n1626, u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, 
       u1_uk_n1635, u1_uk_n1639, u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, 
       u1_uk_n1649, u1_uk_n1651, u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, 
       u1_uk_n1661, u1_uk_n1662, u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, 
       u1_uk_n1676, u1_uk_n1677, u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, 
       u1_uk_n1690, u1_uk_n1691, u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, 
       u1_uk_n1702, u1_uk_n1703, u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, 
       u1_uk_n1712, u1_uk_n1713, u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, 
       u1_uk_n1721, u1_uk_n1722, u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, 
       u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, 
       u1_uk_n1750, u1_uk_n1751, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, 
       u1_uk_n1761, u1_uk_n1762, u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, 
       u1_uk_n1772, u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, 
       u1_uk_n1783, u1_uk_n1784, u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, 
       u1_uk_n1798, u1_uk_n1799, u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, 
       u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, 
       u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, 
       u1_uk_n1827, u1_uk_n1829, u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, 
       u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, 
       u1_uk_n1846, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, 
       u1_uk_n1855, u1_uk_n1856, u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, 
       u1_uk_n1866, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, 
       u1_uk_n1876, u1_uk_n1879, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, 
       u1_uk_n1887, u2_K11_11, u2_K11_21, u2_K11_29, u2_K11_4, u2_K11_6, u2_K11_7, u2_K11_9, u2_K13_37, 
       u2_K13_40, u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, u2_K14_10, u2_K14_11, u2_K14_12, 
       u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_21, u2_K14_3, u2_K14_39, u2_K14_42, 
       u2_K14_6, u2_K14_8, u2_K2_34, u2_K2_35, u2_K2_36, u2_L0_11, u2_L0_19, u2_L0_29, u2_L0_4, 
       u2_L11_12, u2_L11_15, u2_L11_21, u2_L11_22, u2_L11_27, u2_L11_32, u2_L11_5, u2_L11_7, u2_L12_1, 
       u2_L12_10, u2_L12_12, u2_L12_13, u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_2, u2_L12_20, 
       u2_L12_21, u2_L12_22, u2_L12_23, u2_L12_24, u2_L12_26, u2_L12_27, u2_L12_28, u2_L12_30, u2_L12_31, 
       u2_L12_32, u2_L12_5, u2_L12_6, u2_L12_7, u2_L12_9, u2_L9_1, u2_L9_10, u2_L9_13, u2_L9_14, 
       u2_L9_17, u2_L9_18, u2_L9_2, u2_L9_20, u2_L9_23, u2_L9_25, u2_L9_26, u2_L9_28, u2_L9_3, 
       u2_L9_31, u2_L9_8, u2_L9_9, u2_R0_20, u2_R0_21, u2_R0_22, u2_R0_23, u2_R0_24, u2_R0_25, 
       u2_R11_1, u2_R11_24, u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_30, u2_R11_31, 
       u2_R11_32, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_14, u2_R12_15, u2_R12_16, 
       u2_R12_17, u2_R12_2, u2_R12_24, u2_R12_25, u2_R12_26, u2_R12_27, u2_R12_28, u2_R12_29, u2_R12_3, 
       u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, 
       u2_R9_1, u2_R9_12, u2_R9_13, u2_R9_14, u2_R9_15, u2_R9_16, u2_R9_17, u2_R9_18, u2_R9_19, 
       u2_R9_2, u2_R9_20, u2_R9_21, u2_R9_3, u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_6, u2_R9_7, 
       u2_R9_8, u2_R9_9, u2_key_r_1, u2_key_r_13, u2_key_r_54, u2_key_r_8, u2_uk_K_r0_15, u2_uk_K_r0_31, u2_uk_K_r0_36, 
       u2_uk_K_r11_29, u2_uk_K_r12_10, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_33, u2_uk_K_r12_41, u2_uk_K_r9_1, u2_uk_K_r9_10, 
       u2_uk_K_r9_12, u2_uk_K_r9_13, u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_25, u2_uk_K_r9_27, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_K_r9_54, 
       u2_uk_K_r9_9, u2_uk_n100, u2_uk_n102, u2_uk_n110, u2_uk_n117, u2_uk_n118, u2_uk_n1230, u2_uk_n1245, u2_uk_n1258, 
       u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
       u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n1633, u2_uk_n1639, u2_uk_n164, u2_uk_n1642, u2_uk_n1643, u2_uk_n1647, 
       u2_uk_n1652, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, u2_uk_n1660, u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1674, 
       u2_uk_n1675, u2_uk_n1677, u2_uk_n17, u2_uk_n1723, u2_uk_n1725, u2_uk_n1738, u2_uk_n1744, u2_uk_n1755, u2_uk_n1761, 
       u2_uk_n1762, u2_uk_n1768, u2_uk_n1772, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1779, u2_uk_n1781, 
       u2_uk_n1782, u2_uk_n1783, u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, u2_uk_n1791, u2_uk_n1793, 
       u2_uk_n1794, u2_uk_n1796, u2_uk_n1799, u2_uk_n1800, u2_uk_n1801, u2_uk_n1802, u2_uk_n1805, u2_uk_n1806, u2_uk_n1810, 
       u2_uk_n1811, u2_uk_n187, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n220, u2_uk_n222, 
       u2_uk_n223, u2_uk_n230, u2_uk_n238, u2_uk_n31, u2_uk_n313, u2_uk_n363, u2_uk_n63, u2_uk_n677, u2_uk_n702, 
       u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n931, u2_uk_n933, u2_uk_n94, u2_uk_n99, u0_N101, u0_N104, u0_N105, u0_N108, u0_N111, u0_N112, u0_N113, u0_N115, u0_N118, 
        u0_N119, u0_N121, u0_N123, u0_N125, u0_N126, u0_N130, u0_N135, u0_N141, u0_N152, 
        u0_N320, u0_N325, u0_N329, u0_N335, u0_N339, u0_N343, u0_N345, u0_N349, u0_N450, 
        u0_N452, u0_N454, u0_N455, u0_N456, u0_N459, u0_N461, u0_N462, u0_N464, u0_N468, 
        u0_N469, u0_N470, u0_N472, u0_N474, u0_N478, u0_N479, u0_N96, u0_N97, u0_uk_n680, 
        u0_uk_n691, u0_uk_n856, u0_uk_n889, u0_uk_n989, u0_uk_n998, u1_FP_1, u1_FP_10, u1_FP_14, u1_FP_20, 
        u1_FP_25, u1_FP_26, u1_FP_3, u1_FP_8, u1_K10_10, u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_15, 
        u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_27, u1_K10_28, u1_K10_34, 
        u1_K10_36, u1_K11_10, u1_K11_15, u1_K11_16, u1_K11_18, u1_K11_21, u1_K11_27, u1_K11_28, u1_K11_29, 
        u1_K11_3, u1_K11_32, u1_K11_33, u1_K11_4, u1_K11_45, u1_K11_6, u1_K11_7, u1_K11_9, u1_K12_33, 
        u1_K12_34, u1_K12_39, u1_K12_40, u1_K12_45, u1_K12_46, u1_K13_16, u1_K13_33, u1_K13_34, u1_K13_39, 
        u1_K13_40, u1_K13_45, u1_K13_46, u1_K13_9, u1_K14_15, u1_K14_16, u1_K14_21, u1_K14_22, u1_K14_3, 
        u1_K14_33, u1_K14_4, u1_K15_10, u1_K15_21, u1_K15_22, u1_K15_27, u1_K15_28, u1_K15_3, u1_K15_4, 
        u1_K15_9, u1_K16_10, u1_K16_15, u1_K16_16, u1_K16_3, u1_K16_33, u1_K16_39, u1_K16_4, u1_K16_40, 
        u1_K16_45, u1_K16_46, u1_K16_9, u1_K1_15, u1_K1_16, u1_K1_28, u1_K1_29, u1_K1_31, u1_K1_34, 
        u1_K2_33, u1_K2_34, u1_K2_9, u1_K3_10, u1_K3_15, u1_K3_16, u1_K3_27, u1_K3_28, u1_K3_3, 
        u1_K3_33, u1_K3_34, u1_K3_39, u1_K3_4, u1_K3_40, u1_K3_9, u1_K4_15, u1_K4_16, u1_K4_27, 
        u1_K4_28, u1_K4_30, u1_K4_32, u1_K4_33, u1_K4_34, u1_K4_39, u1_K4_40, u1_K4_45, u1_K4_46, 
        u1_K4_9, u1_K5_10, u1_K5_15, u1_K5_16, u1_K5_21, u1_K5_28, u1_K5_3, u1_K5_39, u1_K5_4, 
        u1_K5_40, u1_K5_5, u1_K5_7, u1_K5_9, u1_K6_27, u1_K6_28, u1_K6_29, u1_K6_31, u1_K6_33, 
        u1_K6_34, u1_K6_45, u1_K6_46, u1_K7_10, u1_K7_28, u1_K7_3, u1_K7_33, u1_K7_39, u1_K7_4, 
        u1_K7_40, u1_K7_45, u1_K7_9, u1_K8_21, u1_K8_22, u1_K8_33, u1_K8_45, u1_K8_46, u1_K9_28, 
        u1_K9_3, u1_K9_34, u1_K9_4, u1_N0, u1_N1, u1_N105, u1_N11, u1_N115, u1_N12, 
        u1_N121, u1_N131, u1_N132, u1_N138, u1_N14, u1_N142, u1_N146, u1_N148, u1_N154, 
        u1_N156, u1_N16, u1_N160, u1_N165, u1_N166, u1_N168, u1_N169, u1_N17, u1_N171, 
        u1_N175, u1_N176, u1_N179, u1_N181, u1_N182, u1_N183, u1_N185, u1_N189, u1_N19, 
        u1_N190, u1_N191, u1_N192, u1_N197, u1_N20, u1_N201, u1_N207, u1_N21, u1_N211, 
        u1_N215, u1_N217, u1_N22, u1_N221, u1_N225, u1_N226, u1_N229, u1_N230, u1_N231, 
        u1_N232, u1_N235, u1_N236, u1_N237, u1_N239, u1_N240, u1_N241, u1_N245, u1_N246, 
        u1_N247, u1_N248, u1_N25, u1_N251, u1_N253, u1_N254, u1_N255, u1_N256, u1_N257, 
        u1_N26, u1_N260, u1_N261, u1_N262, u1_N265, u1_N267, u1_N268, u1_N27, u1_N270, 
        u1_N271, u1_N273, u1_N275, u1_N276, u1_N277, u1_N279, u1_N281, u1_N282, u1_N283, 
        u1_N285, u1_N287, u1_N292, u1_N296, u1_N30, u1_N302, u1_N304, u1_N308, u1_N31, 
        u1_N310, u1_N314, u1_N318, u1_N32, u1_N326, u1_N331, u1_N34, u1_N341, u1_N351, 
        u1_N352, u1_N353, u1_N354, u1_N357, u1_N359, u1_N36, u1_N361, u1_N364, u1_N365, 
        u1_N367, u1_N369, u1_N37, u1_N371, u1_N375, u1_N376, u1_N377, u1_N379, u1_N38, 
        u1_N381, u1_N384, u1_N386, u1_N39, u1_N391, u1_N392, u1_N393, u1_N397, u1_N4, 
        u1_N40, u1_N400, u1_N403, u1_N406, u1_N408, u1_N409, u1_N41, u1_N414, u1_N417, 
        u1_N418, u1_N420, u1_N422, u1_N423, u1_N427, u1_N428, u1_N429, u1_N43, u1_N430, 
        u1_N433, u1_N436, u1_N437, u1_N440, u1_N442, u1_N443, u1_N447, u1_N45, u1_N451, 
        u1_N452, u1_N453, u1_N454, u1_N458, u1_N459, u1_N46, u1_N462, u1_N463, u1_N466, 
        u1_N468, u1_N469, u1_N47, u1_N471, u1_N474, u1_N476, u1_N477, u1_N479, u1_N48, 
        u1_N51, u1_N52, u1_N53, u1_N54, u1_N55, u1_N56, u1_N57, u1_N58, u1_N6, 
        u1_N61, u1_N62, u1_N63, u1_N64, u1_N68, u1_N73, u1_N78, u1_N8, u1_N83, 
        u1_N84, u1_N89, u1_N9, u1_N90, u1_N96, u1_u0_X_13, u1_u0_X_14, u1_u0_X_17, u1_u0_X_18, 
        u1_u0_X_25, u1_u0_X_26, u1_u0_X_30, u1_u0_X_32, u1_u0_X_35, u1_u0_X_36, u1_u10_X_1, u1_u10_X_11, u1_u10_X_12, 
        u1_u10_X_13, u1_u10_X_14, u1_u10_X_2, u1_u10_X_23, u1_u10_X_24, u1_u10_X_25, u1_u10_X_26, u1_u10_X_35, u1_u10_X_36, 
        u1_u10_X_43, u1_u10_X_44, u1_u10_X_47, u1_u10_X_48, u1_u11_X_1, u1_u11_X_2, u1_u11_X_31, u1_u11_X_32, u1_u11_X_35, 
        u1_u11_X_36, u1_u11_X_37, u1_u11_X_38, u1_u11_X_41, u1_u11_X_42, u1_u11_X_43, u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, 
        u1_u11_X_5, u1_u11_X_6, u1_u12_X_12, u1_u12_X_14, u1_u12_X_17, u1_u12_X_18, u1_u12_X_31, u1_u12_X_32, u1_u12_X_35, 
        u1_u12_X_36, u1_u12_X_37, u1_u12_X_38, u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_47, u1_u12_X_48, 
        u1_u12_X_7, u1_u12_X_8, u1_u13_X_1, u1_u13_X_13, u1_u13_X_14, u1_u13_X_17, u1_u13_X_18, u1_u13_X_19, u1_u13_X_2, 
        u1_u13_X_20, u1_u13_X_23, u1_u13_X_24, u1_u13_X_31, u1_u13_X_32, u1_u13_X_35, u1_u13_X_36, u1_u13_X_5, u1_u13_X_6, 
        u1_u14_X_1, u1_u14_X_11, u1_u14_X_12, u1_u14_X_19, u1_u14_X_2, u1_u14_X_20, u1_u14_X_23, u1_u14_X_24, u1_u14_X_25, 
        u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u14_X_5, u1_u14_X_6, u1_u14_X_7, u1_u14_X_8, u1_u15_X_1, u1_u15_X_11, 
        u1_u15_X_12, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_2, u1_u15_X_31, u1_u15_X_32, u1_u15_X_35, 
        u1_u15_X_36, u1_u15_X_37, u1_u15_X_38, u1_u15_X_41, u1_u15_X_42, u1_u15_X_43, u1_u15_X_44, u1_u15_X_47, u1_u15_X_48, 
        u1_u15_X_5, u1_u15_X_6, u1_u15_X_7, u1_u15_X_8, u1_u1_X_11, u1_u1_X_12, u1_u1_X_31, u1_u1_X_32, u1_u1_X_35, 
        u1_u1_X_36, u1_u1_X_7, u1_u1_X_8, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_13, u1_u2_X_14, u1_u2_X_17, 
        u1_u2_X_18, u1_u2_X_2, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, u1_u2_X_31, u1_u2_X_32, u1_u2_X_35, 
        u1_u2_X_36, u1_u2_X_37, u1_u2_X_38, u1_u2_X_41, u1_u2_X_42, u1_u2_X_5, u1_u2_X_6, u1_u2_X_7, u1_u2_X_8, 
        u1_u3_X_1, u1_u3_X_11, u1_u3_X_12, u1_u3_X_13, u1_u3_X_14, u1_u3_X_17, u1_u3_X_18, u1_u3_X_2, u1_u3_X_25, 
        u1_u3_X_26, u1_u3_X_35, u1_u3_X_36, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, u1_u3_X_42, u1_u3_X_43, u1_u3_X_44, 
        u1_u3_X_47, u1_u3_X_48, u1_u3_X_5, u1_u3_X_6, u1_u3_X_7, u1_u3_X_8, u1_u4_X_1, u1_u4_X_11, u1_u4_X_12, 
        u1_u4_X_13, u1_u4_X_14, u1_u4_X_17, u1_u4_X_18, u1_u4_X_19, u1_u4_X_2, u1_u4_X_20, u1_u4_X_23, u1_u4_X_24, 
        u1_u4_X_25, u1_u4_X_26, u1_u4_X_29, u1_u4_X_30, u1_u4_X_37, u1_u4_X_38, u1_u4_X_41, u1_u4_X_42, u1_u4_X_6, 
        u1_u4_X_8, u1_u5_X_11, u1_u5_X_12, u1_u5_X_25, u1_u5_X_26, u1_u5_X_30, u1_u5_X_32, u1_u5_X_35, u1_u5_X_36, 
        u1_u5_X_43, u1_u5_X_44, u1_u5_X_47, u1_u5_X_48, u1_u5_X_7, u1_u5_X_8, u1_u6_X_1, u1_u6_X_11, u1_u6_X_12, 
        u1_u6_X_2, u1_u6_X_25, u1_u6_X_26, u1_u6_X_29, u1_u6_X_30, u1_u6_X_31, u1_u6_X_32, u1_u6_X_35, u1_u6_X_36, 
        u1_u6_X_37, u1_u6_X_38, u1_u6_X_41, u1_u6_X_42, u1_u6_X_43, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, u1_u6_X_5, 
        u1_u6_X_6, u1_u6_X_7, u1_u6_X_8, u1_u7_X_19, u1_u7_X_20, u1_u7_X_23, u1_u7_X_24, u1_u7_X_31, u1_u7_X_32, 
        u1_u7_X_35, u1_u7_X_36, u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_1, u1_u8_X_2, u1_u8_X_25, 
        u1_u8_X_26, u1_u8_X_29, u1_u8_X_30, u1_u8_X_31, u1_u8_X_32, u1_u8_X_35, u1_u8_X_36, u1_u8_X_5, u1_u8_X_6, 
        u1_u9_X_23, u1_u9_X_24, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, u1_u9_X_30, u1_u9_X_31, u1_u9_X_32, u1_u9_X_41, 
        u1_u9_X_42, u1_u9_X_7, u1_u9_X_8, u1_uk_n1007, u1_uk_n1011, u1_uk_n1021, u1_uk_n1050, u1_uk_n1060, u1_uk_n1063, 
        u1_uk_n1065, u1_uk_n1067, u1_uk_n1074, u1_uk_n1076, u1_uk_n1088, u1_uk_n1104, u1_uk_n1115, u1_uk_n1119, u1_uk_n1124, 
        u1_uk_n1137, u1_uk_n1159, u1_uk_n1162, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, 
        u1_uk_n373, u1_uk_n375, u1_uk_n376, u1_uk_n385, u1_uk_n386, u1_uk_n391, u1_uk_n407, u1_uk_n421, u1_uk_n437, 
        u1_uk_n443, u1_uk_n468, u1_uk_n496, u1_uk_n501, u1_uk_n601, u1_uk_n656, u1_uk_n671, u1_uk_n672, u1_uk_n677, 
        u1_uk_n678, u1_uk_n955, u1_uk_n988, u2_N320, u2_N321, u2_N322, u2_N327, u2_N328, u2_N329, 
        u2_N332, u2_N333, u2_N336, u2_N337, u2_N339, u2_N342, u2_N344, u2_N345, u2_N347, 
        u2_N35, u2_N350, u2_N388, u2_N390, u2_N395, u2_N398, u2_N404, u2_N405, u2_N410, 
        u2_N415, u2_N416, u2_N417, u2_N42, u2_N420, u2_N421, u2_N422, u2_N424, u2_N425, 
        u2_N427, u2_N428, u2_N430, u2_N431, u2_N432, u2_N433, u2_N435, u2_N436, u2_N437, 
        u2_N438, u2_N439, u2_N441, u2_N442, u2_N443, u2_N445, u2_N446, u2_N447, u2_N50, 
        u2_N60, u2_uk_n1143, u2_uk_n1148, u2_uk_n1150, u2_uk_n1185 );
  input n116, u0_K11_21, u0_K15_47, u0_K4_24, u0_K4_6, u0_K5_26, u0_K5_28, u0_L13_12, u0_L13_14, 
        u0_L13_15, u0_L13_17, u0_L13_21, u0_L13_22, u0_L13_23, u0_L13_25, u0_L13_27, u0_L13_3, u0_L13_31, 
        u0_L13_32, u0_L13_5, u0_L13_7, u0_L13_8, u0_L13_9, u0_L2_1, u0_L2_10, u0_L2_13, u0_L2_16, 
        u0_L2_17, u0_L2_18, u0_L2_2, u0_L2_20, u0_L2_23, u0_L2_24, u0_L2_26, u0_L2_28, u0_L2_30, 
        u0_L2_31, u0_L2_6, u0_L2_9, u0_L3_14, u0_L3_25, u0_L3_3, u0_L3_8, u0_L9_1, u0_L9_10, 
        u0_L9_16, u0_L9_20, u0_L9_24, u0_L9_26, u0_L9_30, u0_L9_6, u0_R13_1, u0_R13_16, u0_R13_17, 
        u0_R13_18, u0_R13_19, u0_R13_2, u0_R13_20, u0_R13_21, u0_R13_24, u0_R13_25, u0_R13_26, u0_R13_27, 
        u0_R13_28, u0_R13_29, u0_R13_3, u0_R13_30, u0_R13_31, u0_R13_32, u0_R13_4, u0_R13_5, u0_R2_1, 
        u0_R2_10, u0_R2_11, u0_R2_12, u0_R2_13, u0_R2_14, u0_R2_15, u0_R2_16, u0_R2_17, u0_R2_2, 
        u0_R2_3, u0_R2_32, u0_R2_4, u0_R2_5, u0_R2_6, u0_R2_7, u0_R2_8, u0_R2_9, u0_R3_16, 
        u0_R3_17, u0_R3_18, u0_R3_19, u0_R3_20, u0_R3_21, u0_R9_10, u0_R9_11, u0_R9_12, u0_R9_13, 
        u0_R9_14, u0_R9_15, u0_R9_16, u0_R9_17, u0_R9_8, u0_R9_9, u0_key_r_18, u0_key_r_33, u0_key_r_44, 
        u0_uk_K_r0_52, u0_uk_K_r13_0, u0_uk_K_r13_2, u0_uk_K_r13_22, u0_uk_K_r13_23, u0_uk_K_r13_35, u0_uk_K_r13_38, u0_uk_K_r13_44, u0_uk_K_r2_13, 
        u0_uk_K_r2_18, u0_uk_K_r2_20, u0_uk_K_r2_25, u0_uk_K_r2_26, u0_uk_K_r2_27, u0_uk_K_r2_33, u0_uk_K_r2_4, u0_uk_K_r2_41, u0_uk_K_r2_46, 
        u0_uk_K_r2_53, u0_uk_K_r2_55, u0_uk_K_r3_35, u0_uk_K_r9_10, u0_uk_K_r9_13, u0_uk_K_r9_19, u0_uk_K_r9_27, u0_uk_K_r9_38, u0_uk_K_r9_48, 
        u0_uk_K_r9_5, u0_uk_n1, u0_uk_n10, u0_uk_n100, u0_uk_n1001, u0_uk_n1002, u0_uk_n109, u0_uk_n110, u0_uk_n117, 
        u0_uk_n118, u0_uk_n12, u0_uk_n128, u0_uk_n129, u0_uk_n13, u0_uk_n141, u0_uk_n142, u0_uk_n146, u0_uk_n147, 
        u0_uk_n148, u0_uk_n155, u0_uk_n161, u0_uk_n163, u0_uk_n164, u0_uk_n17, u0_uk_n182, u0_uk_n187, u0_uk_n188, 
        u0_uk_n190, u0_uk_n196, u0_uk_n197, u0_uk_n20, u0_uk_n200, u0_uk_n201, u0_uk_n202, u0_uk_n203, u0_uk_n206, 
        u0_uk_n207, u0_uk_n208, u0_uk_n21, u0_uk_n212, u0_uk_n214, u0_uk_n215, u0_uk_n217, u0_uk_n22, u0_uk_n220, 
        u0_uk_n221, u0_uk_n222, u0_uk_n23, u0_uk_n230, u0_uk_n238, u0_uk_n24, u0_uk_n240, u0_uk_n242, u0_uk_n250, 
        u0_uk_n251, u0_uk_n252, u0_uk_n26, u0_uk_n27, u0_uk_n29, u0_uk_n3, u0_uk_n30, u0_uk_n31, u0_uk_n33, 
        u0_uk_n34, u0_uk_n36, u0_uk_n38, u0_uk_n39, u0_uk_n4, u0_uk_n40, u0_uk_n41, u0_uk_n462, u0_uk_n463, 
        u0_uk_n475, u0_uk_n480, u0_uk_n481, u0_uk_n497, u0_uk_n5, u0_uk_n502, u0_uk_n510, u0_uk_n511, u0_uk_n517, 
        u0_uk_n519, u0_uk_n523, u0_uk_n525, u0_uk_n529, u0_uk_n530, u0_uk_n531, u0_uk_n534, u0_uk_n535, u0_uk_n536, 
        u0_uk_n6, u0_uk_n60, u0_uk_n8, u0_uk_n813, u0_uk_n83, u0_uk_n834, u0_uk_n839, u0_uk_n9, u0_uk_n916, 
        u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n99, u0_uk_n999, u1_FP_33, u1_FP_36, u1_FP_37, u1_FP_40, 
        u1_FP_41, u1_FP_44, u1_FP_45, u1_FP_46, u1_FP_47, u1_FP_48, u1_FP_49, u1_FP_50, u1_FP_51, 
        u1_FP_52, u1_FP_53, u1_FP_56, u1_FP_57, u1_FP_60, u1_FP_61, u1_FP_64, u1_L0_1, u1_L0_10, 
        u1_L0_12, u1_L0_14, u1_L0_15, u1_L0_16, u1_L0_17, u1_L0_20, u1_L0_21, u1_L0_22, u1_L0_23, 
        u1_L0_24, u1_L0_25, u1_L0_26, u1_L0_27, u1_L0_3, u1_L0_30, u1_L0_31, u1_L0_32, u1_L0_5, 
        u1_L0_6, u1_L0_7, u1_L0_8, u1_L0_9, u1_L10_1, u1_L10_10, u1_L10_13, u1_L10_14, u1_L10_16, 
        u1_L10_18, u1_L10_2, u1_L10_20, u1_L10_24, u1_L10_25, u1_L10_26, u1_L10_28, u1_L10_3, u1_L10_30, 
        u1_L10_6, u1_L10_8, u1_L11_1, u1_L11_10, u1_L11_14, u1_L11_17, u1_L11_20, u1_L11_23, u1_L11_25, 
        u1_L11_26, u1_L11_3, u1_L11_31, u1_L11_8, u1_L11_9, u1_L12_12, u1_L12_13, u1_L12_14, u1_L12_15, 
        u1_L12_18, u1_L12_2, u1_L12_21, u1_L12_22, u1_L12_25, u1_L12_27, u1_L12_28, u1_L12_3, u1_L12_32, 
        u1_L12_5, u1_L12_7, u1_L12_8, u1_L13_11, u1_L13_12, u1_L13_15, u1_L13_16, u1_L13_19, u1_L13_21, 
        u1_L13_22, u1_L13_24, u1_L13_27, u1_L13_29, u1_L13_30, u1_L13_32, u1_L13_4, u1_L13_5, u1_L13_6, 
        u1_L13_7, u1_L14_1, u1_L14_10, u1_L14_14, u1_L14_20, u1_L14_25, u1_L14_26, u1_L14_3, u1_L14_8, 
        u1_L1_1, u1_L1_10, u1_L1_15, u1_L1_20, u1_L1_21, u1_L1_26, u1_L1_27, u1_L1_5, u1_L2_1, 
        u1_L2_10, u1_L2_20, u1_L2_26, u1_L3_11, u1_L3_15, u1_L3_19, u1_L3_21, u1_L3_27, u1_L3_29, 
        u1_L3_4, u1_L3_5, u1_L4_1, u1_L4_10, u1_L4_12, u1_L4_16, u1_L4_17, u1_L4_20, u1_L4_22, 
        u1_L4_23, u1_L4_24, u1_L4_26, u1_L4_30, u1_L4_31, u1_L4_32, u1_L4_6, u1_L4_7, u1_L4_9, 
        u1_L5_1, u1_L5_10, u1_L5_16, u1_L5_20, u1_L5_24, u1_L5_26, u1_L5_30, u1_L5_6, u1_L6_12, 
        u1_L6_13, u1_L6_14, u1_L6_16, u1_L6_17, u1_L6_18, u1_L6_2, u1_L6_22, u1_L6_23, u1_L6_24, 
        u1_L6_25, u1_L6_28, u1_L6_3, u1_L6_30, u1_L6_31, u1_L6_32, u1_L6_6, u1_L6_7, u1_L6_8, 
        u1_L6_9, u1_L7_1, u1_L7_10, u1_L7_12, u1_L7_13, u1_L7_15, u1_L7_16, u1_L7_18, u1_L7_2, 
        u1_L7_20, u1_L7_21, u1_L7_22, u1_L7_24, u1_L7_26, u1_L7_27, u1_L7_28, u1_L7_30, u1_L7_32, 
        u1_L7_5, u1_L7_6, u1_L7_7, u1_L8_15, u1_L8_17, u1_L8_21, u1_L8_23, u1_L8_27, u1_L8_31, 
        u1_L8_5, u1_L8_9, u1_L9_12, u1_L9_22, u1_L9_32, u1_L9_7, u1_R0_1, u1_R0_10, u1_R0_11, 
        u1_R0_12, u1_R0_13, u1_R0_14, u1_R0_15, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_2, 
        u1_R0_20, u1_R0_21, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, u1_R0_3, 
        u1_R0_30, u1_R0_31, u1_R0_32, u1_R0_4, u1_R0_5, u1_R0_8, u1_R0_9, u1_R10_1, u1_R10_10, 
        u1_R10_11, u1_R10_12, u1_R10_13, u1_R10_14, u1_R10_15, u1_R10_16, u1_R10_17, u1_R10_18, u1_R10_19, 
        u1_R10_20, u1_R10_21, u1_R10_24, u1_R10_25, u1_R10_28, u1_R10_29, u1_R10_32, u1_R10_4, u1_R10_5, 
        u1_R10_6, u1_R10_7, u1_R10_8, u1_R10_9, u1_R11_1, u1_R11_12, u1_R11_13, u1_R11_14, u1_R11_15, 
        u1_R11_16, u1_R11_17, u1_R11_18, u1_R11_19, u1_R11_2, u1_R11_20, u1_R11_21, u1_R11_24, u1_R11_25, 
        u1_R11_28, u1_R11_29, u1_R11_3, u1_R11_32, u1_R11_4, u1_R11_5, u1_R11_9, u1_R12_1, u1_R12_12, 
        u1_R12_13, u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, u1_R12_20, u1_R12_21, u1_R12_24, u1_R12_25, 
        u1_R12_26, u1_R12_27, u1_R12_28, u1_R12_29, u1_R12_30, u1_R12_31, u1_R12_32, u1_R12_4, u1_R12_5, 
        u1_R12_6, u1_R12_7, u1_R12_8, u1_R12_9, u1_R13_1, u1_R13_10, u1_R13_11, u1_R13_12, u1_R13_13, 
        u1_R13_16, u1_R13_17, u1_R13_20, u1_R13_21, u1_R13_22, u1_R13_23, u1_R13_24, u1_R13_25, u1_R13_26, 
        u1_R13_27, u1_R13_28, u1_R13_29, u1_R13_30, u1_R13_31, u1_R13_32, u1_R13_4, u1_R13_5, u1_R13_8, 
        u1_R13_9, u1_R1_1, u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, u1_R1_17, u1_R1_20, 
        u1_R1_21, u1_R1_24, u1_R1_25, u1_R1_28, u1_R1_29, u1_R1_30, u1_R1_31, u1_R1_32, u1_R1_4, 
        u1_R1_5, u1_R1_8, u1_R1_9, u1_R2_1, u1_R2_12, u1_R2_13, u1_R2_14, u1_R2_15, u1_R2_16, 
        u1_R2_17, u1_R2_24, u1_R2_25, u1_R2_28, u1_R2_29, u1_R2_32, u1_R2_4, u1_R2_5, u1_R2_8, 
        u1_R2_9, u1_R3_1, u1_R3_12, u1_R3_13, u1_R3_16, u1_R3_17, u1_R3_20, u1_R3_21, u1_R3_22, 
        u1_R3_23, u1_R3_24, u1_R3_25, u1_R3_28, u1_R3_29, u1_R3_30, u1_R3_31, u1_R3_32, u1_R3_5, 
        u1_R3_8, u1_R3_9, u1_R4_1, u1_R4_10, u1_R4_11, u1_R4_12, u1_R4_13, u1_R4_14, u1_R4_15, 
        u1_R4_16, u1_R4_17, u1_R4_2, u1_R4_21, u1_R4_24, u1_R4_25, u1_R4_26, u1_R4_27, u1_R4_28, 
        u1_R4_29, u1_R4_3, u1_R4_32, u1_R4_4, u1_R4_5, u1_R4_8, u1_R4_9, u1_R5_1, u1_R5_10, 
        u1_R5_11, u1_R5_12, u1_R5_13, u1_R5_14, u1_R5_15, u1_R5_16, u1_R5_17, u1_R5_20, u1_R5_21, 
        u1_R5_24, u1_R5_25, u1_R5_28, u1_R5_29, u1_R5_32, u1_R5_4, u1_R5_5, u1_R5_8, u1_R5_9, 
        u1_R6_1, u1_R6_10, u1_R6_11, u1_R6_12, u1_R6_13, u1_R6_16, u1_R6_17, u1_R6_18, u1_R6_19, 
        u1_R6_2, u1_R6_20, u1_R6_21, u1_R6_24, u1_R6_25, u1_R6_26, u1_R6_27, u1_R6_28, u1_R6_29, 
        u1_R6_3, u1_R6_32, u1_R6_4, u1_R6_5, u1_R6_6, u1_R6_7, u1_R6_8, u1_R6_9, u1_R7_1, 
        u1_R7_10, u1_R7_11, u1_R7_12, u1_R7_13, u1_R7_14, u1_R7_15, u1_R7_16, u1_R7_17, u1_R7_20, 
        u1_R7_21, u1_R7_24, u1_R7_25, u1_R7_26, u1_R7_27, u1_R7_28, u1_R7_29, u1_R7_30, u1_R7_31, 
        u1_R7_32, u1_R7_4, u1_R7_5, u1_R7_6, u1_R7_7, u1_R7_8, u1_R7_9, u1_R8_1, u1_R8_16, 
        u1_R8_17, u1_R8_2, u1_R8_20, u1_R8_21, u1_R8_28, u1_R8_29, u1_R8_3, u1_R8_30, u1_R8_31, 
        u1_R8_32, u1_R8_4, u1_R8_5, u1_R9_1, u1_R9_16, u1_R9_17, u1_R9_24, u1_R9_25, u1_R9_26, 
        u1_R9_27, u1_R9_28, u1_R9_29, u1_R9_32, u1_R9_8, u1_R9_9, u1_desIn_r_1, u1_desIn_r_10, u1_desIn_r_12, 
        u1_desIn_r_14, u1_desIn_r_15, u1_desIn_r_16, u1_desIn_r_17, u1_desIn_r_2, u1_desIn_r_23, u1_desIn_r_24, u1_desIn_r_25, u1_desIn_r_26, 
        u1_desIn_r_28, u1_desIn_r_29, u1_desIn_r_3, u1_desIn_r_31, u1_desIn_r_33, u1_desIn_r_34, u1_desIn_r_35, u1_desIn_r_36, u1_desIn_r_37, 
        u1_desIn_r_38, u1_desIn_r_39, u1_desIn_r_4, u1_desIn_r_41, u1_desIn_r_42, u1_desIn_r_45, u1_desIn_r_47, u1_desIn_r_48, u1_desIn_r_49, 
        u1_desIn_r_5, u1_desIn_r_50, u1_desIn_r_52, u1_desIn_r_53, u1_desIn_r_54, u1_desIn_r_55, u1_desIn_r_56, u1_desIn_r_57, u1_desIn_r_59, 
        u1_desIn_r_6, u1_desIn_r_61, u1_desIn_r_63, u1_desIn_r_7, u1_desIn_r_8, u1_desIn_r_9, u1_key_r_0, u1_key_r_1, u1_key_r_10, 
        u1_key_r_11, u1_key_r_12, u1_key_r_13, u1_key_r_14, u1_key_r_15, u1_key_r_16, u1_key_r_17, u1_key_r_18, u1_key_r_19, 
        u1_key_r_2, u1_key_r_20, u1_key_r_21, u1_key_r_22, u1_key_r_23, u1_key_r_24, u1_key_r_25, u1_key_r_26, u1_key_r_27, 
        u1_key_r_28, u1_key_r_29, u1_key_r_3, u1_key_r_30, u1_key_r_31, u1_key_r_32, u1_key_r_33, u1_key_r_34, u1_key_r_35, 
        u1_key_r_36, u1_key_r_37, u1_key_r_38, u1_key_r_39, u1_key_r_4, u1_key_r_40, u1_key_r_41, u1_key_r_42, u1_key_r_43, 
        u1_key_r_44, u1_key_r_45, u1_key_r_46, u1_key_r_47, u1_key_r_48, u1_key_r_49, u1_key_r_5, u1_key_r_50, u1_key_r_51, 
        u1_key_r_52, u1_key_r_53, u1_key_r_54, u1_key_r_55, u1_key_r_6, u1_key_r_7, u1_key_r_8, u1_key_r_9, u1_uk_K_r0_11, 
        u1_uk_K_r0_13, u1_uk_K_r0_15, u1_uk_K_r0_17, u1_uk_K_r0_19, u1_uk_K_r0_2, u1_uk_K_r0_22, u1_uk_K_r0_25, u1_uk_K_r0_28, u1_uk_K_r0_31, 
        u1_uk_K_r0_32, u1_uk_K_r0_34, u1_uk_K_r0_36, u1_uk_K_r0_47, u1_uk_K_r0_49, u1_uk_K_r0_52, u1_uk_K_r0_55, u1_uk_K_r0_7, u1_uk_K_r10_10, 
        u1_uk_K_r10_11, u1_uk_K_r10_14, u1_uk_K_r10_16, u1_uk_K_r10_18, u1_uk_K_r10_19, u1_uk_K_r10_23, u1_uk_K_r10_25, u1_uk_K_r10_27, u1_uk_K_r10_28, 
        u1_uk_K_r10_32, u1_uk_K_r10_34, u1_uk_K_r10_37, u1_uk_K_r10_39, u1_uk_K_r10_4, u1_uk_K_r10_41, u1_uk_K_r10_42, u1_uk_K_r10_43, u1_uk_K_r10_44, 
        u1_uk_K_r10_47, u1_uk_K_r10_48, u1_uk_K_r10_49, u1_uk_K_r10_52, u1_uk_K_r10_9, u1_uk_K_r11_10, u1_uk_K_r11_11, u1_uk_K_r11_17, u1_uk_K_r11_19, 
        u1_uk_K_r11_20, u1_uk_K_r11_21, u1_uk_K_r11_24, u1_uk_K_r11_25, u1_uk_K_r11_26, u1_uk_K_r11_27, u1_uk_K_r11_28, u1_uk_K_r11_29, u1_uk_K_r11_33, 
        u1_uk_K_r11_34, u1_uk_K_r11_39, u1_uk_K_r11_4, u1_uk_K_r11_46, u1_uk_K_r11_47, u1_uk_K_r11_48, u1_uk_K_r11_5, u1_uk_K_r11_53, u1_uk_K_r11_54, 
        u1_uk_K_r11_6, u1_uk_K_r11_7, u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_10, u1_uk_K_r12_15, u1_uk_K_r12_16, u1_uk_K_r12_18, u1_uk_K_r12_21, 
        u1_uk_K_r12_22, u1_uk_K_r12_25, u1_uk_K_r12_30, u1_uk_K_r12_33, u1_uk_K_r12_36, u1_uk_K_r12_41, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_47, 
        u1_uk_K_r12_7, u1_uk_K_r13_0, u1_uk_K_r13_13, u1_uk_K_r13_17, u1_uk_K_r13_19, u1_uk_K_r13_2, u1_uk_K_r13_22, u1_uk_K_r13_23, u1_uk_K_r13_25, 
        u1_uk_K_r13_31, u1_uk_K_r13_32, u1_uk_K_r13_35, u1_uk_K_r13_36, u1_uk_K_r13_38, u1_uk_K_r13_4, u1_uk_K_r13_44, u1_uk_K_r13_55, u1_uk_K_r14_10, 
        u1_uk_K_r14_11, u1_uk_K_r14_12, u1_uk_K_r14_15, u1_uk_K_r14_16, u1_uk_K_r14_18, u1_uk_K_r14_2, u1_uk_K_r14_23, u1_uk_K_r14_3, u1_uk_K_r14_38, 
        u1_uk_K_r14_39, u1_uk_K_r14_42, u1_uk_K_r14_43, u1_uk_K_r14_45, u1_uk_K_r14_46, u1_uk_K_r14_5, u1_uk_K_r14_50, u1_uk_K_r14_8, u1_uk_K_r14_9, 
        u1_uk_K_r1_10, u1_uk_K_r1_15, u1_uk_K_r1_16, u1_uk_K_r1_17, u1_uk_K_r1_18, u1_uk_K_r1_21, u1_uk_K_r1_22, u1_uk_K_r1_33, u1_uk_K_r1_36, 
        u1_uk_K_r1_41, u1_uk_K_r1_42, u1_uk_K_r1_44, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r1_7, u1_uk_K_r2_13, u1_uk_K_r2_16, u1_uk_K_r2_18, 
        u1_uk_K_r2_20, u1_uk_K_r2_21, u1_uk_K_r2_24, u1_uk_K_r2_25, u1_uk_K_r2_26, u1_uk_K_r2_27, u1_uk_K_r2_28, u1_uk_K_r2_29, u1_uk_K_r2_31, 
        u1_uk_K_r2_33, u1_uk_K_r2_36, u1_uk_K_r2_4, u1_uk_K_r2_41, u1_uk_K_r2_46, u1_uk_K_r2_47, u1_uk_K_r2_49, u1_uk_K_r2_50, u1_uk_K_r2_53, 
        u1_uk_K_r2_55, u1_uk_K_r2_6, u1_uk_K_r2_7, u1_uk_K_r3_10, u1_uk_K_r3_11, u1_uk_K_r3_14, u1_uk_K_r3_15, u1_uk_K_r3_16, u1_uk_K_r3_19, 
        u1_uk_K_r3_24, u1_uk_K_r3_29, u1_uk_K_r3_33, u1_uk_K_r3_34, u1_uk_K_r3_35, u1_uk_K_r3_38, u1_uk_K_r3_4, u1_uk_K_r3_43, u1_uk_K_r3_44, 
        u1_uk_K_r3_47, u1_uk_K_r3_51, u1_uk_K_r3_52, u1_uk_K_r3_9, u1_uk_K_r4_0, u1_uk_K_r4_11, u1_uk_K_r4_17, u1_uk_K_r4_18, u1_uk_K_r4_23, 
        u1_uk_K_r4_27, u1_uk_K_r4_3, u1_uk_K_r4_31, u1_uk_K_r4_33, u1_uk_K_r4_35, u1_uk_K_r4_38, u1_uk_K_r4_4, u1_uk_K_r4_41, u1_uk_K_r4_47, 
        u1_uk_K_r4_48, u1_uk_K_r4_49, u1_uk_K_r4_5, u1_uk_K_r4_54, u1_uk_K_r4_55, u1_uk_K_r5_0, u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_13, 
        u1_uk_K_r5_16, u1_uk_K_r5_17, u1_uk_K_r5_18, u1_uk_K_r5_19, u1_uk_K_r5_21, u1_uk_K_r5_23, u1_uk_K_r5_26, u1_uk_K_r5_31, u1_uk_K_r5_32, 
        u1_uk_K_r5_35, u1_uk_K_r5_36, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_40, u1_uk_K_r5_41, u1_uk_K_r5_43, u1_uk_K_r5_48, 
        u1_uk_K_r5_5, u1_uk_K_r5_51, u1_uk_K_r5_53, u1_uk_K_r5_7, u1_uk_K_r5_8, u1_uk_K_r6_0, u1_uk_K_r6_10, u1_uk_K_r6_14, u1_uk_K_r6_17, 
        u1_uk_K_r6_19, u1_uk_K_r6_21, u1_uk_K_r6_22, u1_uk_K_r6_26, u1_uk_K_r6_27, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_3, u1_uk_K_r6_30, 
        u1_uk_K_r6_31, u1_uk_K_r6_34, u1_uk_K_r6_35, u1_uk_K_r6_37, u1_uk_K_r6_46, u1_uk_K_r6_51, u1_uk_K_r6_53, u1_uk_K_r6_55, u1_uk_K_r6_7, 
        u1_uk_K_r7_0, u1_uk_K_r7_1, u1_uk_K_r7_13, u1_uk_K_r7_15, u1_uk_K_r7_16, u1_uk_K_r7_2, u1_uk_K_r7_20, u1_uk_K_r7_22, u1_uk_K_r7_23, 
        u1_uk_K_r7_24, u1_uk_K_r7_25, u1_uk_K_r7_26, u1_uk_K_r7_27, u1_uk_K_r7_29, u1_uk_K_r7_30, u1_uk_K_r7_31, u1_uk_K_r7_32, u1_uk_K_r7_34, 
        u1_uk_K_r7_37, u1_uk_K_r7_39, u1_uk_K_r7_41, u1_uk_K_r7_46, u1_uk_K_r7_48, u1_uk_K_r7_5, u1_uk_K_r7_53, u1_uk_K_r7_55, u1_uk_K_r7_6, 
        u1_uk_K_r7_7, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_10, u1_uk_K_r8_13, u1_uk_K_r8_16, u1_uk_K_r8_17, u1_uk_K_r8_19, u1_uk_K_r8_2, 
        u1_uk_K_r8_21, u1_uk_K_r8_22, u1_uk_K_r8_27, u1_uk_K_r8_28, u1_uk_K_r8_32, u1_uk_K_r8_37, u1_uk_K_r8_39, u1_uk_K_r8_40, u1_uk_K_r8_41, 
        u1_uk_K_r8_42, u1_uk_K_r8_43, u1_uk_K_r8_44, u1_uk_K_r8_48, u1_uk_K_r8_5, u1_uk_K_r8_51, u1_uk_K_r8_52, u1_uk_K_r8_8, u1_uk_K_r9_0, 
        u1_uk_K_r9_1, u1_uk_K_r9_10, u1_uk_K_r9_12, u1_uk_K_r9_13, u1_uk_K_r9_15, u1_uk_K_r9_18, u1_uk_K_r9_19, u1_uk_K_r9_22, u1_uk_K_r9_23, 
        u1_uk_K_r9_25, u1_uk_K_r9_27, u1_uk_K_r9_30, u1_uk_K_r9_31, u1_uk_K_r9_33, u1_uk_K_r9_35, u1_uk_K_r9_38, u1_uk_K_r9_4, u1_uk_K_r9_45, 
        u1_uk_K_r9_48, u1_uk_K_r9_49, u1_uk_K_r9_5, u1_uk_K_r9_54, u1_uk_K_r9_55, u1_uk_K_r9_6, u1_uk_K_r9_7, u1_uk_K_r9_9, u1_uk_n1218, 
        u1_uk_n1219, u1_uk_n1220, u1_uk_n1221, u1_uk_n1222, u1_uk_n1224, u1_uk_n1225, u1_uk_n1227, u1_uk_n1228, u1_uk_n1229, 
        u1_uk_n1230, u1_uk_n1231, u1_uk_n1233, u1_uk_n1234, u1_uk_n1235, u1_uk_n1236, u1_uk_n1237, u1_uk_n1238, u1_uk_n1239, 
        u1_uk_n1240, u1_uk_n1241, u1_uk_n1242, u1_uk_n1243, u1_uk_n1244, u1_uk_n1245, u1_uk_n1246, u1_uk_n1247, u1_uk_n1248, 
        u1_uk_n1249, u1_uk_n1250, u1_uk_n1251, u1_uk_n1252, u1_uk_n1253, u1_uk_n1255, u1_uk_n1256, u1_uk_n1257, u1_uk_n1258, 
        u1_uk_n1259, u1_uk_n1260, u1_uk_n1261, u1_uk_n1262, u1_uk_n1263, u1_uk_n1264, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, 
        u1_uk_n1268, u1_uk_n1269, u1_uk_n1270, u1_uk_n1271, u1_uk_n1272, u1_uk_n1273, u1_uk_n1274, u1_uk_n1275, u1_uk_n1276, 
        u1_uk_n1277, u1_uk_n1278, u1_uk_n1279, u1_uk_n1281, u1_uk_n1282, u1_uk_n1284, u1_uk_n1286, u1_uk_n1288, u1_uk_n1289, 
        u1_uk_n1290, u1_uk_n1291, u1_uk_n1292, u1_uk_n1293, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1297, u1_uk_n1299, 
        u1_uk_n1300, u1_uk_n1303, u1_uk_n1304, u1_uk_n1305, u1_uk_n1307, u1_uk_n1308, u1_uk_n1309, u1_uk_n1310, u1_uk_n1311, 
        u1_uk_n1312, u1_uk_n1313, u1_uk_n1314, u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1318, u1_uk_n1319, u1_uk_n1320, 
        u1_uk_n1321, u1_uk_n1322, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, u1_uk_n1326, u1_uk_n1327, u1_uk_n1328, u1_uk_n1329, 
        u1_uk_n1330, u1_uk_n1331, u1_uk_n1332, u1_uk_n1333, u1_uk_n1334, u1_uk_n1335, u1_uk_n1336, u1_uk_n1338, u1_uk_n1339, 
        u1_uk_n1340, u1_uk_n1341, u1_uk_n1342, u1_uk_n1343, u1_uk_n1344, u1_uk_n1345, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, 
        u1_uk_n1349, u1_uk_n1350, u1_uk_n1351, u1_uk_n1352, u1_uk_n1353, u1_uk_n1354, u1_uk_n1355, u1_uk_n1356, u1_uk_n1357, 
        u1_uk_n1358, u1_uk_n1359, u1_uk_n1360, u1_uk_n1361, u1_uk_n1363, u1_uk_n1365, u1_uk_n1366, u1_uk_n1367, u1_uk_n1369, 
        u1_uk_n1371, u1_uk_n1372, u1_uk_n1374, u1_uk_n1375, u1_uk_n1376, u1_uk_n1377, u1_uk_n1378, u1_uk_n1380, u1_uk_n1381, 
        u1_uk_n1382, u1_uk_n1383, u1_uk_n1386, u1_uk_n1389, u1_uk_n1390, u1_uk_n1391, u1_uk_n1393, u1_uk_n1394, u1_uk_n1395, 
        u1_uk_n1396, u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1400, u1_uk_n1401, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, 
        u1_uk_n1405, u1_uk_n1406, u1_uk_n1407, u1_uk_n1408, u1_uk_n1409, u1_uk_n1410, u1_uk_n1411, u1_uk_n1412, u1_uk_n1413, 
        u1_uk_n1414, u1_uk_n1415, u1_uk_n1417, u1_uk_n1418, u1_uk_n1419, u1_uk_n1422, u1_uk_n1423, u1_uk_n1424, u1_uk_n1425, 
        u1_uk_n1426, u1_uk_n1427, u1_uk_n1429, u1_uk_n1430, u1_uk_n1431, u1_uk_n1433, u1_uk_n1435, u1_uk_n1436, u1_uk_n1437, 
        u1_uk_n1438, u1_uk_n1439, u1_uk_n1440, u1_uk_n1441, u1_uk_n1442, u1_uk_n1443, u1_uk_n1444, u1_uk_n1446, u1_uk_n1447, 
        u1_uk_n1448, u1_uk_n1449, u1_uk_n1450, u1_uk_n1452, u1_uk_n1453, u1_uk_n1454, u1_uk_n1455, u1_uk_n1456, u1_uk_n1457, 
        u1_uk_n1458, u1_uk_n1459, u1_uk_n1460, u1_uk_n1461, u1_uk_n1462, u1_uk_n1463, u1_uk_n1464, u1_uk_n1465, u1_uk_n1466, 
        u1_uk_n1468, u1_uk_n1469, u1_uk_n1470, u1_uk_n1471, u1_uk_n1472, u1_uk_n1474, u1_uk_n1475, u1_uk_n1476, u1_uk_n1477, 
        u1_uk_n1478, u1_uk_n1482, u1_uk_n1483, u1_uk_n1484, u1_uk_n1485, u1_uk_n1486, u1_uk_n1487, u1_uk_n1488, u1_uk_n1489, 
        u1_uk_n1490, u1_uk_n1491, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1496, u1_uk_n1498, u1_uk_n1499, u1_uk_n1500, 
        u1_uk_n1501, u1_uk_n1504, u1_uk_n1505, u1_uk_n1507, u1_uk_n1508, u1_uk_n1510, u1_uk_n1514, u1_uk_n1516, u1_uk_n1517, 
        u1_uk_n1518, u1_uk_n1520, u1_uk_n1521, u1_uk_n1523, u1_uk_n1524, u1_uk_n1526, u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, 
        u1_uk_n1530, u1_uk_n1531, u1_uk_n1532, u1_uk_n1533, u1_uk_n1534, u1_uk_n1536, u1_uk_n1537, u1_uk_n1538, u1_uk_n1540, 
        u1_uk_n1541, u1_uk_n1543, u1_uk_n1544, u1_uk_n1545, u1_uk_n1547, u1_uk_n1548, u1_uk_n1549, u1_uk_n1551, u1_uk_n1552, 
        u1_uk_n1554, u1_uk_n1555, u1_uk_n1556, u1_uk_n1557, u1_uk_n1558, u1_uk_n1559, u1_uk_n1560, u1_uk_n1561, u1_uk_n1562, 
        u1_uk_n1563, u1_uk_n1564, u1_uk_n1565, u1_uk_n1566, u1_uk_n1567, u1_uk_n1568, u1_uk_n1570, u1_uk_n1571, u1_uk_n1572, 
        u1_uk_n1573, u1_uk_n1574, u1_uk_n1577, u1_uk_n1578, u1_uk_n1579, u1_uk_n1581, u1_uk_n1584, u1_uk_n1585, u1_uk_n1586, 
        u1_uk_n1588, u1_uk_n1592, u1_uk_n1593, u1_uk_n1595, u1_uk_n1598, u1_uk_n1599, u1_uk_n1600, u1_uk_n1601, u1_uk_n1603, 
        u1_uk_n1604, u1_uk_n1605, u1_uk_n1606, u1_uk_n1607, u1_uk_n1608, u1_uk_n1610, u1_uk_n1612, u1_uk_n1613, u1_uk_n1614, 
        u1_uk_n1615, u1_uk_n1616, u1_uk_n1618, u1_uk_n1619, u1_uk_n1620, u1_uk_n1621, u1_uk_n1622, u1_uk_n1623, u1_uk_n1624, 
        u1_uk_n1625, u1_uk_n1626, u1_uk_n1627, u1_uk_n1628, u1_uk_n1629, u1_uk_n1630, u1_uk_n1632, u1_uk_n1633, u1_uk_n1634, 
        u1_uk_n1635, u1_uk_n1639, u1_uk_n1640, u1_uk_n1641, u1_uk_n1642, u1_uk_n1643, u1_uk_n1644, u1_uk_n1645, u1_uk_n1647, 
        u1_uk_n1649, u1_uk_n1651, u1_uk_n1652, u1_uk_n1653, u1_uk_n1654, u1_uk_n1655, u1_uk_n1656, u1_uk_n1659, u1_uk_n1660, 
        u1_uk_n1661, u1_uk_n1662, u1_uk_n1663, u1_uk_n1664, u1_uk_n1667, u1_uk_n1669, u1_uk_n1670, u1_uk_n1672, u1_uk_n1673, 
        u1_uk_n1676, u1_uk_n1677, u1_uk_n1678, u1_uk_n1682, u1_uk_n1683, u1_uk_n1684, u1_uk_n1687, u1_uk_n1688, u1_uk_n1689, 
        u1_uk_n1690, u1_uk_n1691, u1_uk_n1692, u1_uk_n1693, u1_uk_n1694, u1_uk_n1695, u1_uk_n1696, u1_uk_n1698, u1_uk_n1699, 
        u1_uk_n1702, u1_uk_n1703, u1_uk_n1704, u1_uk_n1705, u1_uk_n1707, u1_uk_n1708, u1_uk_n1709, u1_uk_n1710, u1_uk_n1711, 
        u1_uk_n1712, u1_uk_n1713, u1_uk_n1714, u1_uk_n1715, u1_uk_n1716, u1_uk_n1717, u1_uk_n1718, u1_uk_n1719, u1_uk_n1720, 
        u1_uk_n1721, u1_uk_n1722, u1_uk_n1723, u1_uk_n1728, u1_uk_n1729, u1_uk_n1730, u1_uk_n1731, u1_uk_n1732, u1_uk_n1734, 
        u1_uk_n1735, u1_uk_n1736, u1_uk_n1737, u1_uk_n1738, u1_uk_n1739, u1_uk_n1744, u1_uk_n1745, u1_uk_n1748, u1_uk_n1749, 
        u1_uk_n1750, u1_uk_n1751, u1_uk_n1752, u1_uk_n1753, u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1757, u1_uk_n1758, 
        u1_uk_n1761, u1_uk_n1762, u1_uk_n1763, u1_uk_n1764, u1_uk_n1765, u1_uk_n1766, u1_uk_n1767, u1_uk_n1768, u1_uk_n1769, 
        u1_uk_n1772, u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1777, u1_uk_n1780, u1_uk_n1781, u1_uk_n1782, 
        u1_uk_n1783, u1_uk_n1784, u1_uk_n1785, u1_uk_n1787, u1_uk_n1790, u1_uk_n1791, u1_uk_n1792, u1_uk_n1793, u1_uk_n1797, 
        u1_uk_n1798, u1_uk_n1799, u1_uk_n1800, u1_uk_n1801, u1_uk_n1802, u1_uk_n1803, u1_uk_n1804, u1_uk_n1806, u1_uk_n1807, 
        u1_uk_n1808, u1_uk_n1809, u1_uk_n1810, u1_uk_n1811, u1_uk_n1812, u1_uk_n1813, u1_uk_n1814, u1_uk_n1815, u1_uk_n1816, 
        u1_uk_n1817, u1_uk_n1818, u1_uk_n1819, u1_uk_n1820, u1_uk_n1821, u1_uk_n1822, u1_uk_n1823, u1_uk_n1824, u1_uk_n1826, 
        u1_uk_n1827, u1_uk_n1829, u1_uk_n1830, u1_uk_n1831, u1_uk_n1832, u1_uk_n1833, u1_uk_n1834, u1_uk_n1835, u1_uk_n1836, 
        u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n1840, u1_uk_n1841, u1_uk_n1842, u1_uk_n1843, u1_uk_n1844, u1_uk_n1845, 
        u1_uk_n1846, u1_uk_n1847, u1_uk_n1848, u1_uk_n1849, u1_uk_n1850, u1_uk_n1851, u1_uk_n1852, u1_uk_n1853, u1_uk_n1854, 
        u1_uk_n1855, u1_uk_n1856, u1_uk_n1858, u1_uk_n1859, u1_uk_n1860, u1_uk_n1862, u1_uk_n1863, u1_uk_n1864, u1_uk_n1865, 
        u1_uk_n1866, u1_uk_n1867, u1_uk_n1868, u1_uk_n1869, u1_uk_n1870, u1_uk_n1872, u1_uk_n1873, u1_uk_n1874, u1_uk_n1875, 
        u1_uk_n1876, u1_uk_n1879, u1_uk_n1880, u1_uk_n1881, u1_uk_n1882, u1_uk_n1883, u1_uk_n1884, u1_uk_n1885, u1_uk_n1886, 
        u1_uk_n1887, u2_K11_11, u2_K11_21, u2_K11_29, u2_K11_4, u2_K11_6, u2_K11_7, u2_K11_9, u2_K13_37, 
        u2_K13_40, u2_K13_42, u2_K13_44, u2_K13_45, u2_K13_46, u2_K13_47, u2_K14_10, u2_K14_11, u2_K14_12, 
        u2_K14_13, u2_K14_14, u2_K14_16, u2_K14_17, u2_K14_18, u2_K14_21, u2_K14_3, u2_K14_39, u2_K14_42, 
        u2_K14_6, u2_K14_8, u2_K2_34, u2_K2_35, u2_K2_36, u2_L0_11, u2_L0_19, u2_L0_29, u2_L0_4, 
        u2_L11_12, u2_L11_15, u2_L11_21, u2_L11_22, u2_L11_27, u2_L11_32, u2_L11_5, u2_L11_7, u2_L12_1, 
        u2_L12_10, u2_L12_12, u2_L12_13, u2_L12_15, u2_L12_16, u2_L12_17, u2_L12_18, u2_L12_2, u2_L12_20, 
        u2_L12_21, u2_L12_22, u2_L12_23, u2_L12_24, u2_L12_26, u2_L12_27, u2_L12_28, u2_L12_30, u2_L12_31, 
        u2_L12_32, u2_L12_5, u2_L12_6, u2_L12_7, u2_L12_9, u2_L9_1, u2_L9_10, u2_L9_13, u2_L9_14, 
        u2_L9_17, u2_L9_18, u2_L9_2, u2_L9_20, u2_L9_23, u2_L9_25, u2_L9_26, u2_L9_28, u2_L9_3, 
        u2_L9_31, u2_L9_8, u2_L9_9, u2_R0_20, u2_R0_21, u2_R0_22, u2_R0_23, u2_R0_24, u2_R0_25, 
        u2_R11_1, u2_R11_24, u2_R11_25, u2_R11_26, u2_R11_27, u2_R11_28, u2_R11_29, u2_R11_30, u2_R11_31, 
        u2_R11_32, u2_R12_1, u2_R12_10, u2_R12_11, u2_R12_12, u2_R12_13, u2_R12_14, u2_R12_15, u2_R12_16, 
        u2_R12_17, u2_R12_2, u2_R12_24, u2_R12_25, u2_R12_26, u2_R12_27, u2_R12_28, u2_R12_29, u2_R12_3, 
        u2_R12_30, u2_R12_31, u2_R12_32, u2_R12_4, u2_R12_5, u2_R12_6, u2_R12_7, u2_R12_8, u2_R12_9, 
        u2_R9_1, u2_R9_12, u2_R9_13, u2_R9_14, u2_R9_15, u2_R9_16, u2_R9_17, u2_R9_18, u2_R9_19, 
        u2_R9_2, u2_R9_20, u2_R9_21, u2_R9_3, u2_R9_32, u2_R9_4, u2_R9_5, u2_R9_6, u2_R9_7, 
        u2_R9_8, u2_R9_9, u2_key_r_1, u2_key_r_13, u2_key_r_54, u2_key_r_8, u2_uk_K_r0_15, u2_uk_K_r0_31, u2_uk_K_r0_36, 
        u2_uk_K_r11_29, u2_uk_K_r12_10, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r12_25, u2_uk_K_r12_33, u2_uk_K_r12_41, u2_uk_K_r9_1, u2_uk_K_r9_10, 
        u2_uk_K_r9_12, u2_uk_K_r9_13, u2_uk_K_r9_18, u2_uk_K_r9_19, u2_uk_K_r9_25, u2_uk_K_r9_27, u2_uk_K_r9_4, u2_uk_K_r9_48, u2_uk_K_r9_54, 
        u2_uk_K_r9_9, u2_uk_n100, u2_uk_n102, u2_uk_n110, u2_uk_n117, u2_uk_n118, u2_uk_n1230, u2_uk_n1245, u2_uk_n1258, 
        u2_uk_n128, u2_uk_n129, u2_uk_n141, u2_uk_n142, u2_uk_n145, u2_uk_n146, u2_uk_n147, u2_uk_n148, u2_uk_n155, 
        u2_uk_n161, u2_uk_n162, u2_uk_n163, u2_uk_n1633, u2_uk_n1639, u2_uk_n164, u2_uk_n1642, u2_uk_n1643, u2_uk_n1647, 
        u2_uk_n1652, u2_uk_n1654, u2_uk_n1657, u2_uk_n1658, u2_uk_n1660, u2_uk_n1665, u2_uk_n1666, u2_uk_n1668, u2_uk_n1674, 
        u2_uk_n1675, u2_uk_n1677, u2_uk_n17, u2_uk_n1723, u2_uk_n1725, u2_uk_n1738, u2_uk_n1744, u2_uk_n1755, u2_uk_n1761, 
        u2_uk_n1762, u2_uk_n1768, u2_uk_n1772, u2_uk_n1773, u2_uk_n1776, u2_uk_n1777, u2_uk_n1778, u2_uk_n1779, u2_uk_n1781, 
        u2_uk_n1782, u2_uk_n1783, u2_uk_n1785, u2_uk_n1786, u2_uk_n1788, u2_uk_n1789, u2_uk_n1790, u2_uk_n1791, u2_uk_n1793, 
        u2_uk_n1794, u2_uk_n1796, u2_uk_n1799, u2_uk_n1800, u2_uk_n1801, u2_uk_n1802, u2_uk_n1805, u2_uk_n1806, u2_uk_n1810, 
        u2_uk_n1811, u2_uk_n187, u2_uk_n207, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n220, u2_uk_n222, 
        u2_uk_n223, u2_uk_n230, u2_uk_n238, u2_uk_n31, u2_uk_n313, u2_uk_n363, u2_uk_n63, u2_uk_n677, u2_uk_n702, 
        u2_uk_n83, u2_uk_n92, u2_uk_n93, u2_uk_n931, u2_uk_n933, u2_uk_n94, u2_uk_n99;
  output u0_N101, u0_N104, u0_N105, u0_N108, u0_N111, u0_N112, u0_N113, u0_N115, u0_N118, 
        u0_N119, u0_N121, u0_N123, u0_N125, u0_N126, u0_N130, u0_N135, u0_N141, u0_N152, 
        u0_N320, u0_N325, u0_N329, u0_N335, u0_N339, u0_N343, u0_N345, u0_N349, u0_N450, 
        u0_N452, u0_N454, u0_N455, u0_N456, u0_N459, u0_N461, u0_N462, u0_N464, u0_N468, 
        u0_N469, u0_N470, u0_N472, u0_N474, u0_N478, u0_N479, u0_N96, u0_N97, u0_uk_n680, 
        u0_uk_n691, u0_uk_n856, u0_uk_n889, u0_uk_n989, u0_uk_n998, u1_FP_1, u1_FP_10, u1_FP_14, u1_FP_20, 
        u1_FP_25, u1_FP_26, u1_FP_3, u1_FP_8, u1_K10_10, u1_K10_11, u1_K10_13, u1_K10_14, u1_K10_15, 
        u1_K10_16, u1_K10_17, u1_K10_18, u1_K10_19, u1_K10_20, u1_K10_21, u1_K10_27, u1_K10_28, u1_K10_34, 
        u1_K10_36, u1_K11_10, u1_K11_15, u1_K11_16, u1_K11_18, u1_K11_21, u1_K11_27, u1_K11_28, u1_K11_29, 
        u1_K11_3, u1_K11_32, u1_K11_33, u1_K11_4, u1_K11_45, u1_K11_6, u1_K11_7, u1_K11_9, u1_K12_33, 
        u1_K12_34, u1_K12_39, u1_K12_40, u1_K12_45, u1_K12_46, u1_K13_16, u1_K13_33, u1_K13_34, u1_K13_39, 
        u1_K13_40, u1_K13_45, u1_K13_46, u1_K13_9, u1_K14_15, u1_K14_16, u1_K14_21, u1_K14_22, u1_K14_3, 
        u1_K14_33, u1_K14_4, u1_K15_10, u1_K15_21, u1_K15_22, u1_K15_27, u1_K15_28, u1_K15_3, u1_K15_4, 
        u1_K15_9, u1_K16_10, u1_K16_15, u1_K16_16, u1_K16_3, u1_K16_33, u1_K16_39, u1_K16_4, u1_K16_40, 
        u1_K16_45, u1_K16_46, u1_K16_9, u1_K1_15, u1_K1_16, u1_K1_28, u1_K1_29, u1_K1_31, u1_K1_34, 
        u1_K2_33, u1_K2_34, u1_K2_9, u1_K3_10, u1_K3_15, u1_K3_16, u1_K3_27, u1_K3_28, u1_K3_3, 
        u1_K3_33, u1_K3_34, u1_K3_39, u1_K3_4, u1_K3_40, u1_K3_9, u1_K4_15, u1_K4_16, u1_K4_27, 
        u1_K4_28, u1_K4_30, u1_K4_32, u1_K4_33, u1_K4_34, u1_K4_39, u1_K4_40, u1_K4_45, u1_K4_46, 
        u1_K4_9, u1_K5_10, u1_K5_15, u1_K5_16, u1_K5_21, u1_K5_28, u1_K5_3, u1_K5_39, u1_K5_4, 
        u1_K5_40, u1_K5_5, u1_K5_7, u1_K5_9, u1_K6_27, u1_K6_28, u1_K6_29, u1_K6_31, u1_K6_33, 
        u1_K6_34, u1_K6_45, u1_K6_46, u1_K7_10, u1_K7_28, u1_K7_3, u1_K7_33, u1_K7_39, u1_K7_4, 
        u1_K7_40, u1_K7_45, u1_K7_9, u1_K8_21, u1_K8_22, u1_K8_33, u1_K8_45, u1_K8_46, u1_K9_28, 
        u1_K9_3, u1_K9_34, u1_K9_4, u1_N0, u1_N1, u1_N105, u1_N11, u1_N115, u1_N12, 
        u1_N121, u1_N131, u1_N132, u1_N138, u1_N14, u1_N142, u1_N146, u1_N148, u1_N154, 
        u1_N156, u1_N16, u1_N160, u1_N165, u1_N166, u1_N168, u1_N169, u1_N17, u1_N171, 
        u1_N175, u1_N176, u1_N179, u1_N181, u1_N182, u1_N183, u1_N185, u1_N189, u1_N19, 
        u1_N190, u1_N191, u1_N192, u1_N197, u1_N20, u1_N201, u1_N207, u1_N21, u1_N211, 
        u1_N215, u1_N217, u1_N22, u1_N221, u1_N225, u1_N226, u1_N229, u1_N230, u1_N231, 
        u1_N232, u1_N235, u1_N236, u1_N237, u1_N239, u1_N240, u1_N241, u1_N245, u1_N246, 
        u1_N247, u1_N248, u1_N25, u1_N251, u1_N253, u1_N254, u1_N255, u1_N256, u1_N257, 
        u1_N26, u1_N260, u1_N261, u1_N262, u1_N265, u1_N267, u1_N268, u1_N27, u1_N270, 
        u1_N271, u1_N273, u1_N275, u1_N276, u1_N277, u1_N279, u1_N281, u1_N282, u1_N283, 
        u1_N285, u1_N287, u1_N292, u1_N296, u1_N30, u1_N302, u1_N304, u1_N308, u1_N31, 
        u1_N310, u1_N314, u1_N318, u1_N32, u1_N326, u1_N331, u1_N34, u1_N341, u1_N351, 
        u1_N352, u1_N353, u1_N354, u1_N357, u1_N359, u1_N36, u1_N361, u1_N364, u1_N365, 
        u1_N367, u1_N369, u1_N37, u1_N371, u1_N375, u1_N376, u1_N377, u1_N379, u1_N38, 
        u1_N381, u1_N384, u1_N386, u1_N39, u1_N391, u1_N392, u1_N393, u1_N397, u1_N4, 
        u1_N40, u1_N400, u1_N403, u1_N406, u1_N408, u1_N409, u1_N41, u1_N414, u1_N417, 
        u1_N418, u1_N420, u1_N422, u1_N423, u1_N427, u1_N428, u1_N429, u1_N43, u1_N430, 
        u1_N433, u1_N436, u1_N437, u1_N440, u1_N442, u1_N443, u1_N447, u1_N45, u1_N451, 
        u1_N452, u1_N453, u1_N454, u1_N458, u1_N459, u1_N46, u1_N462, u1_N463, u1_N466, 
        u1_N468, u1_N469, u1_N47, u1_N471, u1_N474, u1_N476, u1_N477, u1_N479, u1_N48, 
        u1_N51, u1_N52, u1_N53, u1_N54, u1_N55, u1_N56, u1_N57, u1_N58, u1_N6, 
        u1_N61, u1_N62, u1_N63, u1_N64, u1_N68, u1_N73, u1_N78, u1_N8, u1_N83, 
        u1_N84, u1_N89, u1_N9, u1_N90, u1_N96, u1_u0_X_13, u1_u0_X_14, u1_u0_X_17, u1_u0_X_18, 
        u1_u0_X_25, u1_u0_X_26, u1_u0_X_30, u1_u0_X_32, u1_u0_X_35, u1_u0_X_36, u1_u10_X_1, u1_u10_X_11, u1_u10_X_12, 
        u1_u10_X_13, u1_u10_X_14, u1_u10_X_2, u1_u10_X_23, u1_u10_X_24, u1_u10_X_25, u1_u10_X_26, u1_u10_X_35, u1_u10_X_36, 
        u1_u10_X_43, u1_u10_X_44, u1_u10_X_47, u1_u10_X_48, u1_u11_X_1, u1_u11_X_2, u1_u11_X_31, u1_u11_X_32, u1_u11_X_35, 
        u1_u11_X_36, u1_u11_X_37, u1_u11_X_38, u1_u11_X_41, u1_u11_X_42, u1_u11_X_43, u1_u11_X_44, u1_u11_X_47, u1_u11_X_48, 
        u1_u11_X_5, u1_u11_X_6, u1_u12_X_12, u1_u12_X_14, u1_u12_X_17, u1_u12_X_18, u1_u12_X_31, u1_u12_X_32, u1_u12_X_35, 
        u1_u12_X_36, u1_u12_X_37, u1_u12_X_38, u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_47, u1_u12_X_48, 
        u1_u12_X_7, u1_u12_X_8, u1_u13_X_1, u1_u13_X_13, u1_u13_X_14, u1_u13_X_17, u1_u13_X_18, u1_u13_X_19, u1_u13_X_2, 
        u1_u13_X_20, u1_u13_X_23, u1_u13_X_24, u1_u13_X_31, u1_u13_X_32, u1_u13_X_35, u1_u13_X_36, u1_u13_X_5, u1_u13_X_6, 
        u1_u14_X_1, u1_u14_X_11, u1_u14_X_12, u1_u14_X_19, u1_u14_X_2, u1_u14_X_20, u1_u14_X_23, u1_u14_X_24, u1_u14_X_25, 
        u1_u14_X_26, u1_u14_X_29, u1_u14_X_30, u1_u14_X_5, u1_u14_X_6, u1_u14_X_7, u1_u14_X_8, u1_u15_X_1, u1_u15_X_11, 
        u1_u15_X_12, u1_u15_X_13, u1_u15_X_14, u1_u15_X_17, u1_u15_X_18, u1_u15_X_2, u1_u15_X_31, u1_u15_X_32, u1_u15_X_35, 
        u1_u15_X_36, u1_u15_X_37, u1_u15_X_38, u1_u15_X_41, u1_u15_X_42, u1_u15_X_43, u1_u15_X_44, u1_u15_X_47, u1_u15_X_48, 
        u1_u15_X_5, u1_u15_X_6, u1_u15_X_7, u1_u15_X_8, u1_u1_X_11, u1_u1_X_12, u1_u1_X_31, u1_u1_X_32, u1_u1_X_35, 
        u1_u1_X_36, u1_u1_X_7, u1_u1_X_8, u1_u2_X_1, u1_u2_X_11, u1_u2_X_12, u1_u2_X_13, u1_u2_X_14, u1_u2_X_17, 
        u1_u2_X_18, u1_u2_X_2, u1_u2_X_25, u1_u2_X_26, u1_u2_X_29, u1_u2_X_30, u1_u2_X_31, u1_u2_X_32, u1_u2_X_35, 
        u1_u2_X_36, u1_u2_X_37, u1_u2_X_38, u1_u2_X_41, u1_u2_X_42, u1_u2_X_5, u1_u2_X_6, u1_u2_X_7, u1_u2_X_8, 
        u1_u3_X_1, u1_u3_X_11, u1_u3_X_12, u1_u3_X_13, u1_u3_X_14, u1_u3_X_17, u1_u3_X_18, u1_u3_X_2, u1_u3_X_25, 
        u1_u3_X_26, u1_u3_X_35, u1_u3_X_36, u1_u3_X_37, u1_u3_X_38, u1_u3_X_41, u1_u3_X_42, u1_u3_X_43, u1_u3_X_44, 
        u1_u3_X_47, u1_u3_X_48, u1_u3_X_5, u1_u3_X_6, u1_u3_X_7, u1_u3_X_8, u1_u4_X_1, u1_u4_X_11, u1_u4_X_12, 
        u1_u4_X_13, u1_u4_X_14, u1_u4_X_17, u1_u4_X_18, u1_u4_X_19, u1_u4_X_2, u1_u4_X_20, u1_u4_X_23, u1_u4_X_24, 
        u1_u4_X_25, u1_u4_X_26, u1_u4_X_29, u1_u4_X_30, u1_u4_X_37, u1_u4_X_38, u1_u4_X_41, u1_u4_X_42, u1_u4_X_6, 
        u1_u4_X_8, u1_u5_X_11, u1_u5_X_12, u1_u5_X_25, u1_u5_X_26, u1_u5_X_30, u1_u5_X_32, u1_u5_X_35, u1_u5_X_36, 
        u1_u5_X_43, u1_u5_X_44, u1_u5_X_47, u1_u5_X_48, u1_u5_X_7, u1_u5_X_8, u1_u6_X_1, u1_u6_X_11, u1_u6_X_12, 
        u1_u6_X_2, u1_u6_X_25, u1_u6_X_26, u1_u6_X_29, u1_u6_X_30, u1_u6_X_31, u1_u6_X_32, u1_u6_X_35, u1_u6_X_36, 
        u1_u6_X_37, u1_u6_X_38, u1_u6_X_41, u1_u6_X_42, u1_u6_X_43, u1_u6_X_44, u1_u6_X_47, u1_u6_X_48, u1_u6_X_5, 
        u1_u6_X_6, u1_u6_X_7, u1_u6_X_8, u1_u7_X_19, u1_u7_X_20, u1_u7_X_23, u1_u7_X_24, u1_u7_X_31, u1_u7_X_32, 
        u1_u7_X_35, u1_u7_X_36, u1_u7_X_43, u1_u7_X_44, u1_u7_X_47, u1_u7_X_48, u1_u8_X_1, u1_u8_X_2, u1_u8_X_25, 
        u1_u8_X_26, u1_u8_X_29, u1_u8_X_30, u1_u8_X_31, u1_u8_X_32, u1_u8_X_35, u1_u8_X_36, u1_u8_X_5, u1_u8_X_6, 
        u1_u9_X_23, u1_u9_X_24, u1_u9_X_25, u1_u9_X_26, u1_u9_X_29, u1_u9_X_30, u1_u9_X_31, u1_u9_X_32, u1_u9_X_41, 
        u1_u9_X_42, u1_u9_X_7, u1_u9_X_8, u1_uk_n1007, u1_uk_n1011, u1_uk_n1021, u1_uk_n1050, u1_uk_n1060, u1_uk_n1063, 
        u1_uk_n1065, u1_uk_n1067, u1_uk_n1074, u1_uk_n1076, u1_uk_n1088, u1_uk_n1104, u1_uk_n1115, u1_uk_n1119, u1_uk_n1124, 
        u1_uk_n1137, u1_uk_n1159, u1_uk_n1162, u1_uk_n299, u1_uk_n312, u1_uk_n349, u1_uk_n353, u1_uk_n366, u1_uk_n369, 
        u1_uk_n373, u1_uk_n375, u1_uk_n376, u1_uk_n385, u1_uk_n386, u1_uk_n391, u1_uk_n407, u1_uk_n421, u1_uk_n437, 
        u1_uk_n443, u1_uk_n468, u1_uk_n496, u1_uk_n501, u1_uk_n601, u1_uk_n656, u1_uk_n671, u1_uk_n672, u1_uk_n677, 
        u1_uk_n678, u1_uk_n955, u1_uk_n988, u2_N320, u2_N321, u2_N322, u2_N327, u2_N328, u2_N329, 
        u2_N332, u2_N333, u2_N336, u2_N337, u2_N339, u2_N342, u2_N344, u2_N345, u2_N347, 
        u2_N35, u2_N350, u2_N388, u2_N390, u2_N395, u2_N398, u2_N404, u2_N405, u2_N410, 
        u2_N415, u2_N416, u2_N417, u2_N42, u2_N420, u2_N421, u2_N422, u2_N424, u2_N425, 
        u2_N427, u2_N428, u2_N430, u2_N431, u2_N432, u2_N433, u2_N435, u2_N436, u2_N437, 
        u2_N438, u2_N439, u2_N441, u2_N442, u2_N443, u2_N445, u2_N446, u2_N447, u2_N50, 
        u2_N60, u2_uk_n1143, u2_uk_n1148, u2_uk_n1150, u2_uk_n1185;
  wire u0_K11_13, u0_K11_14, u0_K11_15, u0_K11_16, u0_K11_17, u0_K11_18, u0_K11_19, u0_K11_20, u0_K11_22, 
       u0_K11_23, u0_K11_24, u0_K15_1, u0_K15_2, u0_K15_25, u0_K15_26, u0_K15_27, u0_K15_28, u0_K15_29, 
       u0_K15_3, u0_K15_30, u0_K15_37, u0_K15_38, u0_K15_39, u0_K15_4, u0_K15_40, u0_K15_41, u0_K15_42, 
       u0_K15_43, u0_K15_44, u0_K15_45, u0_K15_46, u0_K15_48, u0_K15_5, u0_K15_6, u0_K4_1, u0_K4_10, 
       u0_K4_11, u0_K4_12, u0_K4_13, u0_K4_14, u0_K4_15, u0_K4_16, u0_K4_17, u0_K4_18, u0_K4_19, 
       u0_K4_2, u0_K4_20, u0_K4_21, u0_K4_22, u0_K4_23, u0_K4_3, u0_K4_4, u0_K4_5, u0_K4_7, 
       u0_K4_8, u0_K4_9, u0_K5_25, u0_K5_27, u0_K5_29, u0_K5_30, u0_out10_1, u0_out10_10, u0_out10_16, 
       u0_out10_20, u0_out10_24, u0_out10_26, u0_out10_30, u0_out10_6, u0_out14_12, u0_out14_14, u0_out14_15, u0_out14_17, 
       u0_out14_21, u0_out14_22, u0_out14_23, u0_out14_25, u0_out14_27, u0_out14_3, u0_out14_31, u0_out14_32, u0_out14_5, 
       u0_out14_7, u0_out14_8, u0_out14_9, u0_out3_1, u0_out3_10, u0_out3_13, u0_out3_16, u0_out3_17, u0_out3_18, 
       u0_out3_2, u0_out3_20, u0_out3_23, u0_out3_24, u0_out3_26, u0_out3_28, u0_out3_30, u0_out3_31, u0_out3_6, 
       u0_out3_9, u0_out4_14, u0_out4_25, u0_out4_3, u0_out4_8, u0_u10_X_13, u0_u10_X_14, u0_u10_X_15, u0_u10_X_16, 
       u0_u10_X_17, u0_u10_X_18, u0_u10_X_19, u0_u10_X_20, u0_u10_X_21, u0_u10_X_22, u0_u10_X_23, u0_u10_X_24, u0_u10_u2_n100, 
       u0_u10_u2_n101, u0_u10_u2_n102, u0_u10_u2_n103, u0_u10_u2_n104, u0_u10_u2_n105, u0_u10_u2_n106, u0_u10_u2_n107, u0_u10_u2_n108, u0_u10_u2_n109, 
       u0_u10_u2_n110, u0_u10_u2_n111, u0_u10_u2_n112, u0_u10_u2_n113, u0_u10_u2_n114, u0_u10_u2_n115, u0_u10_u2_n116, u0_u10_u2_n117, u0_u10_u2_n118, 
       u0_u10_u2_n119, u0_u10_u2_n120, u0_u10_u2_n121, u0_u10_u2_n122, u0_u10_u2_n123, u0_u10_u2_n124, u0_u10_u2_n125, u0_u10_u2_n126, u0_u10_u2_n127, 
       u0_u10_u2_n128, u0_u10_u2_n129, u0_u10_u2_n130, u0_u10_u2_n131, u0_u10_u2_n132, u0_u10_u2_n133, u0_u10_u2_n134, u0_u10_u2_n135, u0_u10_u2_n136, 
       u0_u10_u2_n137, u0_u10_u2_n138, u0_u10_u2_n139, u0_u10_u2_n140, u0_u10_u2_n141, u0_u10_u2_n142, u0_u10_u2_n143, u0_u10_u2_n144, u0_u10_u2_n145, 
       u0_u10_u2_n146, u0_u10_u2_n147, u0_u10_u2_n148, u0_u10_u2_n149, u0_u10_u2_n150, u0_u10_u2_n151, u0_u10_u2_n152, u0_u10_u2_n153, u0_u10_u2_n154, 
       u0_u10_u2_n155, u0_u10_u2_n156, u0_u10_u2_n157, u0_u10_u2_n158, u0_u10_u2_n159, u0_u10_u2_n160, u0_u10_u2_n161, u0_u10_u2_n162, u0_u10_u2_n163, 
       u0_u10_u2_n164, u0_u10_u2_n165, u0_u10_u2_n166, u0_u10_u2_n167, u0_u10_u2_n168, u0_u10_u2_n169, u0_u10_u2_n170, u0_u10_u2_n171, u0_u10_u2_n172, 
       u0_u10_u2_n173, u0_u10_u2_n174, u0_u10_u2_n175, u0_u10_u2_n176, u0_u10_u2_n177, u0_u10_u2_n178, u0_u10_u2_n179, u0_u10_u2_n180, u0_u10_u2_n181, 
       u0_u10_u2_n182, u0_u10_u2_n183, u0_u10_u2_n184, u0_u10_u2_n185, u0_u10_u2_n186, u0_u10_u2_n187, u0_u10_u2_n188, u0_u10_u2_n95, u0_u10_u2_n96, 
       u0_u10_u2_n97, u0_u10_u2_n98, u0_u10_u2_n99, u0_u10_u3_n100, u0_u10_u3_n101, u0_u10_u3_n102, u0_u10_u3_n103, u0_u10_u3_n104, u0_u10_u3_n105, 
       u0_u10_u3_n106, u0_u10_u3_n107, u0_u10_u3_n108, u0_u10_u3_n109, u0_u10_u3_n110, u0_u10_u3_n111, u0_u10_u3_n112, u0_u10_u3_n113, u0_u10_u3_n114, 
       u0_u10_u3_n115, u0_u10_u3_n116, u0_u10_u3_n117, u0_u10_u3_n118, u0_u10_u3_n119, u0_u10_u3_n120, u0_u10_u3_n121, u0_u10_u3_n122, u0_u10_u3_n123, 
       u0_u10_u3_n124, u0_u10_u3_n125, u0_u10_u3_n126, u0_u10_u3_n127, u0_u10_u3_n128, u0_u10_u3_n129, u0_u10_u3_n130, u0_u10_u3_n131, u0_u10_u3_n132, 
       u0_u10_u3_n133, u0_u10_u3_n134, u0_u10_u3_n135, u0_u10_u3_n136, u0_u10_u3_n137, u0_u10_u3_n138, u0_u10_u3_n139, u0_u10_u3_n140, u0_u10_u3_n141, 
       u0_u10_u3_n142, u0_u10_u3_n143, u0_u10_u3_n144, u0_u10_u3_n145, u0_u10_u3_n146, u0_u10_u3_n147, u0_u10_u3_n148, u0_u10_u3_n149, u0_u10_u3_n150, 
       u0_u10_u3_n151, u0_u10_u3_n152, u0_u10_u3_n153, u0_u10_u3_n154, u0_u10_u3_n155, u0_u10_u3_n156, u0_u10_u3_n157, u0_u10_u3_n158, u0_u10_u3_n159, 
       u0_u10_u3_n160, u0_u10_u3_n161, u0_u10_u3_n162, u0_u10_u3_n163, u0_u10_u3_n164, u0_u10_u3_n165, u0_u10_u3_n166, u0_u10_u3_n167, u0_u10_u3_n168, 
       u0_u10_u3_n169, u0_u10_u3_n170, u0_u10_u3_n171, u0_u10_u3_n172, u0_u10_u3_n173, u0_u10_u3_n174, u0_u10_u3_n175, u0_u10_u3_n176, u0_u10_u3_n177, 
       u0_u10_u3_n178, u0_u10_u3_n179, u0_u10_u3_n180, u0_u10_u3_n181, u0_u10_u3_n182, u0_u10_u3_n183, u0_u10_u3_n184, u0_u10_u3_n185, u0_u10_u3_n186, 
       u0_u10_u3_n94, u0_u10_u3_n95, u0_u10_u3_n96, u0_u10_u3_n97, u0_u10_u3_n98, u0_u10_u3_n99, u0_u14_X_1, u0_u14_X_2, u0_u14_X_25, 
       u0_u14_X_26, u0_u14_X_27, u0_u14_X_28, u0_u14_X_29, u0_u14_X_3, u0_u14_X_30, u0_u14_X_37, u0_u14_X_38, u0_u14_X_39, 
       u0_u14_X_4, u0_u14_X_40, u0_u14_X_41, u0_u14_X_42, u0_u14_X_43, u0_u14_X_44, u0_u14_X_45, u0_u14_X_46, u0_u14_X_47, 
       u0_u14_X_48, u0_u14_X_5, u0_u14_X_6, u0_u14_u0_n100, u0_u14_u0_n101, u0_u14_u0_n102, u0_u14_u0_n103, u0_u14_u0_n104, u0_u14_u0_n105, 
       u0_u14_u0_n106, u0_u14_u0_n107, u0_u14_u0_n108, u0_u14_u0_n109, u0_u14_u0_n110, u0_u14_u0_n111, u0_u14_u0_n112, u0_u14_u0_n113, u0_u14_u0_n114, 
       u0_u14_u0_n115, u0_u14_u0_n116, u0_u14_u0_n117, u0_u14_u0_n118, u0_u14_u0_n119, u0_u14_u0_n120, u0_u14_u0_n121, u0_u14_u0_n122, u0_u14_u0_n123, 
       u0_u14_u0_n124, u0_u14_u0_n125, u0_u14_u0_n126, u0_u14_u0_n127, u0_u14_u0_n128, u0_u14_u0_n129, u0_u14_u0_n130, u0_u14_u0_n131, u0_u14_u0_n132, 
       u0_u14_u0_n133, u0_u14_u0_n134, u0_u14_u0_n135, u0_u14_u0_n136, u0_u14_u0_n137, u0_u14_u0_n138, u0_u14_u0_n139, u0_u14_u0_n140, u0_u14_u0_n141, 
       u0_u14_u0_n142, u0_u14_u0_n143, u0_u14_u0_n144, u0_u14_u0_n145, u0_u14_u0_n146, u0_u14_u0_n147, u0_u14_u0_n148, u0_u14_u0_n149, u0_u14_u0_n150, 
       u0_u14_u0_n151, u0_u14_u0_n152, u0_u14_u0_n153, u0_u14_u0_n154, u0_u14_u0_n155, u0_u14_u0_n156, u0_u14_u0_n157, u0_u14_u0_n158, u0_u14_u0_n159, 
       u0_u14_u0_n160, u0_u14_u0_n161, u0_u14_u0_n162, u0_u14_u0_n163, u0_u14_u0_n164, u0_u14_u0_n165, u0_u14_u0_n166, u0_u14_u0_n167, u0_u14_u0_n168, 
       u0_u14_u0_n169, u0_u14_u0_n170, u0_u14_u0_n171, u0_u14_u0_n172, u0_u14_u0_n173, u0_u14_u0_n174, u0_u14_u0_n88, u0_u14_u0_n89, u0_u14_u0_n90, 
       u0_u14_u0_n91, u0_u14_u0_n92, u0_u14_u0_n93, u0_u14_u0_n94, u0_u14_u0_n95, u0_u14_u0_n96, u0_u14_u0_n97, u0_u14_u0_n98, u0_u14_u0_n99, 
       u0_u14_u4_n100, u0_u14_u4_n101, u0_u14_u4_n102, u0_u14_u4_n103, u0_u14_u4_n104, u0_u14_u4_n105, u0_u14_u4_n106, u0_u14_u4_n107, u0_u14_u4_n108, 
       u0_u14_u4_n109, u0_u14_u4_n110, u0_u14_u4_n111, u0_u14_u4_n112, u0_u14_u4_n113, u0_u14_u4_n114, u0_u14_u4_n115, u0_u14_u4_n116, u0_u14_u4_n117, 
       u0_u14_u4_n118, u0_u14_u4_n119, u0_u14_u4_n120, u0_u14_u4_n121, u0_u14_u4_n122, u0_u14_u4_n123, u0_u14_u4_n124, u0_u14_u4_n125, u0_u14_u4_n126, 
       u0_u14_u4_n127, u0_u14_u4_n128, u0_u14_u4_n129, u0_u14_u4_n130, u0_u14_u4_n131, u0_u14_u4_n132, u0_u14_u4_n133, u0_u14_u4_n134, u0_u14_u4_n135, 
       u0_u14_u4_n136, u0_u14_u4_n137, u0_u14_u4_n138, u0_u14_u4_n139, u0_u14_u4_n140, u0_u14_u4_n141, u0_u14_u4_n142, u0_u14_u4_n143, u0_u14_u4_n144, 
       u0_u14_u4_n145, u0_u14_u4_n146, u0_u14_u4_n147, u0_u14_u4_n148, u0_u14_u4_n149, u0_u14_u4_n150, u0_u14_u4_n151, u0_u14_u4_n152, u0_u14_u4_n153, 
       u0_u14_u4_n154, u0_u14_u4_n155, u0_u14_u4_n156, u0_u14_u4_n157, u0_u14_u4_n158, u0_u14_u4_n159, u0_u14_u4_n160, u0_u14_u4_n161, u0_u14_u4_n162, 
       u0_u14_u4_n163, u0_u14_u4_n164, u0_u14_u4_n165, u0_u14_u4_n166, u0_u14_u4_n167, u0_u14_u4_n168, u0_u14_u4_n169, u0_u14_u4_n170, u0_u14_u4_n171, 
       u0_u14_u4_n172, u0_u14_u4_n173, u0_u14_u4_n174, u0_u14_u4_n175, u0_u14_u4_n176, u0_u14_u4_n177, u0_u14_u4_n178, u0_u14_u4_n179, u0_u14_u4_n180, 
       u0_u14_u4_n181, u0_u14_u4_n182, u0_u14_u4_n183, u0_u14_u4_n184, u0_u14_u4_n185, u0_u14_u4_n186, u0_u14_u4_n94, u0_u14_u4_n95, u0_u14_u4_n96, 
       u0_u14_u4_n97, u0_u14_u4_n98, u0_u14_u4_n99, u0_u14_u6_n100, u0_u14_u6_n101, u0_u14_u6_n102, u0_u14_u6_n103, u0_u14_u6_n104, u0_u14_u6_n105, 
       u0_u14_u6_n106, u0_u14_u6_n107, u0_u14_u6_n108, u0_u14_u6_n109, u0_u14_u6_n110, u0_u14_u6_n111, u0_u14_u6_n112, u0_u14_u6_n113, u0_u14_u6_n114, 
       u0_u14_u6_n115, u0_u14_u6_n116, u0_u14_u6_n117, u0_u14_u6_n118, u0_u14_u6_n119, u0_u14_u6_n120, u0_u14_u6_n121, u0_u14_u6_n122, u0_u14_u6_n123, 
       u0_u14_u6_n124, u0_u14_u6_n125, u0_u14_u6_n126, u0_u14_u6_n127, u0_u14_u6_n128, u0_u14_u6_n129, u0_u14_u6_n130, u0_u14_u6_n131, u0_u14_u6_n132, 
       u0_u14_u6_n133, u0_u14_u6_n134, u0_u14_u6_n135, u0_u14_u6_n136, u0_u14_u6_n137, u0_u14_u6_n138, u0_u14_u6_n139, u0_u14_u6_n140, u0_u14_u6_n141, 
       u0_u14_u6_n142, u0_u14_u6_n143, u0_u14_u6_n144, u0_u14_u6_n145, u0_u14_u6_n146, u0_u14_u6_n147, u0_u14_u6_n148, u0_u14_u6_n149, u0_u14_u6_n150, 
       u0_u14_u6_n151, u0_u14_u6_n152, u0_u14_u6_n153, u0_u14_u6_n154, u0_u14_u6_n155, u0_u14_u6_n156, u0_u14_u6_n157, u0_u14_u6_n158, u0_u14_u6_n159, 
       u0_u14_u6_n160, u0_u14_u6_n161, u0_u14_u6_n162, u0_u14_u6_n163, u0_u14_u6_n164, u0_u14_u6_n165, u0_u14_u6_n166, u0_u14_u6_n167, u0_u14_u6_n168, 
       u0_u14_u6_n169, u0_u14_u6_n170, u0_u14_u6_n171, u0_u14_u6_n172, u0_u14_u6_n173, u0_u14_u6_n174, u0_u14_u6_n88, u0_u14_u6_n89, u0_u14_u6_n90, 
       u0_u14_u6_n91, u0_u14_u6_n92, u0_u14_u6_n93, u0_u14_u6_n94, u0_u14_u6_n95, u0_u14_u6_n96, u0_u14_u6_n97, u0_u14_u6_n98, u0_u14_u6_n99, 
       u0_u14_u7_n100, u0_u14_u7_n101, u0_u14_u7_n102, u0_u14_u7_n103, u0_u14_u7_n104, u0_u14_u7_n105, u0_u14_u7_n106, u0_u14_u7_n107, u0_u14_u7_n108, 
       u0_u14_u7_n109, u0_u14_u7_n110, u0_u14_u7_n111, u0_u14_u7_n112, u0_u14_u7_n113, u0_u14_u7_n114, u0_u14_u7_n115, u0_u14_u7_n116, u0_u14_u7_n117, 
       u0_u14_u7_n118, u0_u14_u7_n119, u0_u14_u7_n120, u0_u14_u7_n121, u0_u14_u7_n122, u0_u14_u7_n123, u0_u14_u7_n124, u0_u14_u7_n125, u0_u14_u7_n126, 
       u0_u14_u7_n127, u0_u14_u7_n128, u0_u14_u7_n129, u0_u14_u7_n130, u0_u14_u7_n131, u0_u14_u7_n132, u0_u14_u7_n133, u0_u14_u7_n134, u0_u14_u7_n135, 
       u0_u14_u7_n136, u0_u14_u7_n137, u0_u14_u7_n138, u0_u14_u7_n139, u0_u14_u7_n140, u0_u14_u7_n141, u0_u14_u7_n142, u0_u14_u7_n143, u0_u14_u7_n144, 
       u0_u14_u7_n145, u0_u14_u7_n146, u0_u14_u7_n147, u0_u14_u7_n148, u0_u14_u7_n149, u0_u14_u7_n150, u0_u14_u7_n151, u0_u14_u7_n152, u0_u14_u7_n153, 
       u0_u14_u7_n154, u0_u14_u7_n155, u0_u14_u7_n156, u0_u14_u7_n157, u0_u14_u7_n158, u0_u14_u7_n159, u0_u14_u7_n160, u0_u14_u7_n161, u0_u14_u7_n162, 
       u0_u14_u7_n163, u0_u14_u7_n164, u0_u14_u7_n165, u0_u14_u7_n166, u0_u14_u7_n167, u0_u14_u7_n168, u0_u14_u7_n169, u0_u14_u7_n170, u0_u14_u7_n171, 
       u0_u14_u7_n172, u0_u14_u7_n173, u0_u14_u7_n174, u0_u14_u7_n175, u0_u14_u7_n176, u0_u14_u7_n177, u0_u14_u7_n178, u0_u14_u7_n179, u0_u14_u7_n180, 
       u0_u14_u7_n91, u0_u14_u7_n92, u0_u14_u7_n93, u0_u14_u7_n94, u0_u14_u7_n95, u0_u14_u7_n96, u0_u14_u7_n97, u0_u14_u7_n98, u0_u14_u7_n99, 
       u0_u3_X_1, u0_u3_X_10, u0_u3_X_11, u0_u3_X_12, u0_u3_X_13, u0_u3_X_14, u0_u3_X_15, u0_u3_X_16, u0_u3_X_17, 
       u0_u3_X_18, u0_u3_X_19, u0_u3_X_2, u0_u3_X_20, u0_u3_X_21, u0_u3_X_22, u0_u3_X_23, u0_u3_X_24, u0_u3_X_3, 
       u0_u3_X_4, u0_u3_X_5, u0_u3_X_6, u0_u3_X_7, u0_u3_X_8, u0_u3_X_9, u0_u3_u0_n100, u0_u3_u0_n101, u0_u3_u0_n102, 
       u0_u3_u0_n103, u0_u3_u0_n104, u0_u3_u0_n105, u0_u3_u0_n106, u0_u3_u0_n107, u0_u3_u0_n108, u0_u3_u0_n109, u0_u3_u0_n110, u0_u3_u0_n111, 
       u0_u3_u0_n112, u0_u3_u0_n113, u0_u3_u0_n114, u0_u3_u0_n115, u0_u3_u0_n116, u0_u3_u0_n117, u0_u3_u0_n118, u0_u3_u0_n119, u0_u3_u0_n120, 
       u0_u3_u0_n121, u0_u3_u0_n122, u0_u3_u0_n123, u0_u3_u0_n124, u0_u3_u0_n125, u0_u3_u0_n126, u0_u3_u0_n127, u0_u3_u0_n128, u0_u3_u0_n129, 
       u0_u3_u0_n130, u0_u3_u0_n131, u0_u3_u0_n132, u0_u3_u0_n133, u0_u3_u0_n134, u0_u3_u0_n135, u0_u3_u0_n136, u0_u3_u0_n137, u0_u3_u0_n138, 
       u0_u3_u0_n139, u0_u3_u0_n140, u0_u3_u0_n141, u0_u3_u0_n142, u0_u3_u0_n143, u0_u3_u0_n144, u0_u3_u0_n145, u0_u3_u0_n146, u0_u3_u0_n147, 
       u0_u3_u0_n148, u0_u3_u0_n149, u0_u3_u0_n150, u0_u3_u0_n151, u0_u3_u0_n152, u0_u3_u0_n153, u0_u3_u0_n154, u0_u3_u0_n155, u0_u3_u0_n156, 
       u0_u3_u0_n157, u0_u3_u0_n158, u0_u3_u0_n159, u0_u3_u0_n160, u0_u3_u0_n161, u0_u3_u0_n162, u0_u3_u0_n163, u0_u3_u0_n164, u0_u3_u0_n165, 
       u0_u3_u0_n166, u0_u3_u0_n167, u0_u3_u0_n168, u0_u3_u0_n169, u0_u3_u0_n170, u0_u3_u0_n171, u0_u3_u0_n172, u0_u3_u0_n173, u0_u3_u0_n174, 
       u0_u3_u0_n175, u0_u3_u0_n176, u0_u3_u0_n88, u0_u3_u0_n89, u0_u3_u0_n90, u0_u3_u0_n91, u0_u3_u0_n92, u0_u3_u0_n93, u0_u3_u0_n94, 
       u0_u3_u0_n95, u0_u3_u0_n96, u0_u3_u0_n97, u0_u3_u0_n98, u0_u3_u0_n99, u0_u3_u1_n100, u0_u3_u1_n101, u0_u3_u1_n102, u0_u3_u1_n103, 
       u0_u3_u1_n104, u0_u3_u1_n105, u0_u3_u1_n106, u0_u3_u1_n107, u0_u3_u1_n108, u0_u3_u1_n109, u0_u3_u1_n110, u0_u3_u1_n111, u0_u3_u1_n112, 
       u0_u3_u1_n113, u0_u3_u1_n114, u0_u3_u1_n115, u0_u3_u1_n116, u0_u3_u1_n117, u0_u3_u1_n118, u0_u3_u1_n119, u0_u3_u1_n120, u0_u3_u1_n121, 
       u0_u3_u1_n122, u0_u3_u1_n123, u0_u3_u1_n124, u0_u3_u1_n125, u0_u3_u1_n126, u0_u3_u1_n127, u0_u3_u1_n128, u0_u3_u1_n129, u0_u3_u1_n130, 
       u0_u3_u1_n131, u0_u3_u1_n132, u0_u3_u1_n133, u0_u3_u1_n134, u0_u3_u1_n135, u0_u3_u1_n136, u0_u3_u1_n137, u0_u3_u1_n138, u0_u3_u1_n139, 
       u0_u3_u1_n140, u0_u3_u1_n141, u0_u3_u1_n142, u0_u3_u1_n143, u0_u3_u1_n144, u0_u3_u1_n145, u0_u3_u1_n146, u0_u3_u1_n147, u0_u3_u1_n148, 
       u0_u3_u1_n149, u0_u3_u1_n150, u0_u3_u1_n151, u0_u3_u1_n152, u0_u3_u1_n153, u0_u3_u1_n154, u0_u3_u1_n155, u0_u3_u1_n156, u0_u3_u1_n157, 
       u0_u3_u1_n158, u0_u3_u1_n159, u0_u3_u1_n160, u0_u3_u1_n161, u0_u3_u1_n162, u0_u3_u1_n163, u0_u3_u1_n164, u0_u3_u1_n165, u0_u3_u1_n166, 
       u0_u3_u1_n167, u0_u3_u1_n168, u0_u3_u1_n169, u0_u3_u1_n170, u0_u3_u1_n171, u0_u3_u1_n172, u0_u3_u1_n173, u0_u3_u1_n174, u0_u3_u1_n175, 
       u0_u3_u1_n176, u0_u3_u1_n177, u0_u3_u1_n178, u0_u3_u1_n179, u0_u3_u1_n180, u0_u3_u1_n181, u0_u3_u1_n182, u0_u3_u1_n183, u0_u3_u1_n184, 
       u0_u3_u1_n185, u0_u3_u1_n186, u0_u3_u1_n187, u0_u3_u1_n188, u0_u3_u1_n95, u0_u3_u1_n96, u0_u3_u1_n97, u0_u3_u1_n98, u0_u3_u1_n99, 
       u0_u3_u2_n100, u0_u3_u2_n101, u0_u3_u2_n102, u0_u3_u2_n103, u0_u3_u2_n104, u0_u3_u2_n105, u0_u3_u2_n106, u0_u3_u2_n107, u0_u3_u2_n108, 
       u0_u3_u2_n109, u0_u3_u2_n110, u0_u3_u2_n111, u0_u3_u2_n112, u0_u3_u2_n113, u0_u3_u2_n114, u0_u3_u2_n115, u0_u3_u2_n116, u0_u3_u2_n117, 
       u0_u3_u2_n118, u0_u3_u2_n119, u0_u3_u2_n120, u0_u3_u2_n121, u0_u3_u2_n122, u0_u3_u2_n123, u0_u3_u2_n124, u0_u3_u2_n125, u0_u3_u2_n126, 
       u0_u3_u2_n127, u0_u3_u2_n128, u0_u3_u2_n129, u0_u3_u2_n130, u0_u3_u2_n131, u0_u3_u2_n132, u0_u3_u2_n133, u0_u3_u2_n134, u0_u3_u2_n135, 
       u0_u3_u2_n136, u0_u3_u2_n137, u0_u3_u2_n138, u0_u3_u2_n139, u0_u3_u2_n140, u0_u3_u2_n141, u0_u3_u2_n142, u0_u3_u2_n143, u0_u3_u2_n144, 
       u0_u3_u2_n145, u0_u3_u2_n146, u0_u3_u2_n147, u0_u3_u2_n148, u0_u3_u2_n149, u0_u3_u2_n150, u0_u3_u2_n151, u0_u3_u2_n152, u0_u3_u2_n153, 
       u0_u3_u2_n154, u0_u3_u2_n155, u0_u3_u2_n156, u0_u3_u2_n157, u0_u3_u2_n158, u0_u3_u2_n159, u0_u3_u2_n160, u0_u3_u2_n161, u0_u3_u2_n162, 
       u0_u3_u2_n163, u0_u3_u2_n164, u0_u3_u2_n165, u0_u3_u2_n166, u0_u3_u2_n167, u0_u3_u2_n168, u0_u3_u2_n169, u0_u3_u2_n170, u0_u3_u2_n171, 
       u0_u3_u2_n172, u0_u3_u2_n173, u0_u3_u2_n174, u0_u3_u2_n175, u0_u3_u2_n176, u0_u3_u2_n177, u0_u3_u2_n178, u0_u3_u2_n179, u0_u3_u2_n180, 
       u0_u3_u2_n181, u0_u3_u2_n182, u0_u3_u2_n183, u0_u3_u2_n184, u0_u3_u2_n185, u0_u3_u2_n186, u0_u3_u2_n187, u0_u3_u2_n188, u0_u3_u2_n95, 
       u0_u3_u2_n96, u0_u3_u2_n97, u0_u3_u2_n98, u0_u3_u2_n99, u0_u3_u3_n100, u0_u3_u3_n101, u0_u3_u3_n102, u0_u3_u3_n103, u0_u3_u3_n104, 
       u0_u3_u3_n105, u0_u3_u3_n106, u0_u3_u3_n107, u0_u3_u3_n108, u0_u3_u3_n109, u0_u3_u3_n110, u0_u3_u3_n111, u0_u3_u3_n112, u0_u3_u3_n113, 
       u0_u3_u3_n114, u0_u3_u3_n115, u0_u3_u3_n116, u0_u3_u3_n117, u0_u3_u3_n118, u0_u3_u3_n119, u0_u3_u3_n120, u0_u3_u3_n121, u0_u3_u3_n122, 
       u0_u3_u3_n123, u0_u3_u3_n124, u0_u3_u3_n125, u0_u3_u3_n126, u0_u3_u3_n127, u0_u3_u3_n128, u0_u3_u3_n129, u0_u3_u3_n130, u0_u3_u3_n131, 
       u0_u3_u3_n132, u0_u3_u3_n133, u0_u3_u3_n134, u0_u3_u3_n135, u0_u3_u3_n136, u0_u3_u3_n137, u0_u3_u3_n138, u0_u3_u3_n139, u0_u3_u3_n140, 
       u0_u3_u3_n141, u0_u3_u3_n142, u0_u3_u3_n143, u0_u3_u3_n144, u0_u3_u3_n145, u0_u3_u3_n146, u0_u3_u3_n147, u0_u3_u3_n148, u0_u3_u3_n149, 
       u0_u3_u3_n150, u0_u3_u3_n151, u0_u3_u3_n152, u0_u3_u3_n153, u0_u3_u3_n154, u0_u3_u3_n155, u0_u3_u3_n156, u0_u3_u3_n157, u0_u3_u3_n158, 
       u0_u3_u3_n159, u0_u3_u3_n160, u0_u3_u3_n161, u0_u3_u3_n162, u0_u3_u3_n163, u0_u3_u3_n164, u0_u3_u3_n165, u0_u3_u3_n166, u0_u3_u3_n167, 
       u0_u3_u3_n168, u0_u3_u3_n169, u0_u3_u3_n170, u0_u3_u3_n171, u0_u3_u3_n172, u0_u3_u3_n173, u0_u3_u3_n174, u0_u3_u3_n175, u0_u3_u3_n176, 
       u0_u3_u3_n177, u0_u3_u3_n178, u0_u3_u3_n179, u0_u3_u3_n180, u0_u3_u3_n181, u0_u3_u3_n182, u0_u3_u3_n183, u0_u3_u3_n184, u0_u3_u3_n185, 
       u0_u3_u3_n186, u0_u3_u3_n94, u0_u3_u3_n95, u0_u3_u3_n96, u0_u3_u3_n97, u0_u3_u3_n98, u0_u3_u3_n99, u0_u4_X_25, u0_u4_X_26, 
       u0_u4_X_27, u0_u4_X_28, u0_u4_X_29, u0_u4_X_30, u0_u4_u4_n100, u0_u4_u4_n101, u0_u4_u4_n102, u0_u4_u4_n103, u0_u4_u4_n104, 
       u0_u4_u4_n105, u0_u4_u4_n106, u0_u4_u4_n107, u0_u4_u4_n108, u0_u4_u4_n109, u0_u4_u4_n110, u0_u4_u4_n111, u0_u4_u4_n112, u0_u4_u4_n113, 
       u0_u4_u4_n114, u0_u4_u4_n115, u0_u4_u4_n116, u0_u4_u4_n117, u0_u4_u4_n118, u0_u4_u4_n119, u0_u4_u4_n120, u0_u4_u4_n121, u0_u4_u4_n122, 
       u0_u4_u4_n123, u0_u4_u4_n124, u0_u4_u4_n125, u0_u4_u4_n126, u0_u4_u4_n127, u0_u4_u4_n128, u0_u4_u4_n129, u0_u4_u4_n130, u0_u4_u4_n131, 
       u0_u4_u4_n132, u0_u4_u4_n133, u0_u4_u4_n134, u0_u4_u4_n135, u0_u4_u4_n136, u0_u4_u4_n137, u0_u4_u4_n138, u0_u4_u4_n139, u0_u4_u4_n140, 
       u0_u4_u4_n141, u0_u4_u4_n142, u0_u4_u4_n143, u0_u4_u4_n144, u0_u4_u4_n145, u0_u4_u4_n146, u0_u4_u4_n147, u0_u4_u4_n148, u0_u4_u4_n149, 
       u0_u4_u4_n150, u0_u4_u4_n151, u0_u4_u4_n152, u0_u4_u4_n153, u0_u4_u4_n154, u0_u4_u4_n155, u0_u4_u4_n156, u0_u4_u4_n157, u0_u4_u4_n158, 
       u0_u4_u4_n159, u0_u4_u4_n160, u0_u4_u4_n161, u0_u4_u4_n162, u0_u4_u4_n163, u0_u4_u4_n164, u0_u4_u4_n165, u0_u4_u4_n166, u0_u4_u4_n167, 
       u0_u4_u4_n168, u0_u4_u4_n169, u0_u4_u4_n170, u0_u4_u4_n171, u0_u4_u4_n172, u0_u4_u4_n173, u0_u4_u4_n174, u0_u4_u4_n175, u0_u4_u4_n176, 
       u0_u4_u4_n177, u0_u4_u4_n178, u0_u4_u4_n179, u0_u4_u4_n180, u0_u4_u4_n181, u0_u4_u4_n182, u0_u4_u4_n183, u0_u4_u4_n184, u0_u4_u4_n185, 
       u0_u4_u4_n186, u0_u4_u4_n94, u0_u4_u4_n95, u0_u4_u4_n96, u0_u4_u4_n97, u0_u4_u4_n98, u0_u4_u4_n99, u0_uk_n1000, u0_uk_n814, 
       u0_uk_n819, u0_uk_n821, u0_uk_n822, u0_uk_n824, u0_uk_n828, u0_uk_n833, u0_uk_n835, u0_uk_n836, u0_uk_n837, 
       u0_uk_n838, u0_uk_n914, u0_uk_n915, u0_uk_n919, u0_uk_n920, u0_uk_n921, u0_uk_n996, u0_uk_n997, u1_K10_1, 
       u1_K10_2, u1_K10_23, u1_K10_24, u1_K10_25, u1_K10_26, u1_K10_29, u1_K10_3, u1_K10_30, u1_K10_31, 
       u1_K10_32, u1_K10_4, u1_K10_41, u1_K10_42, u1_K10_43, u1_K10_44, u1_K10_45, u1_K10_46, u1_K10_47, 
       u1_K10_48, u1_K10_5, u1_K10_6, u1_K10_7, u1_K10_8, u1_K11_1, u1_K11_11, u1_K11_12, u1_K11_13, 
       u1_K11_14, u1_K11_2, u1_K11_23, u1_K11_24, u1_K11_25, u1_K11_26, u1_K11_35, u1_K11_36, u1_K11_37, 
       u1_K11_38, u1_K11_39, u1_K11_40, u1_K11_41, u1_K11_42, u1_K11_43, u1_K11_44, u1_K11_47, u1_K11_48, 
       u1_K12_1, u1_K12_10, u1_K12_11, u1_K12_12, u1_K12_13, u1_K12_14, u1_K12_15, u1_K12_16, u1_K12_17, 
       u1_K12_18, u1_K12_19, u1_K12_2, u1_K12_20, u1_K12_21, u1_K12_22, u1_K12_23, u1_K12_24, u1_K12_25, 
       u1_K12_26, u1_K12_27, u1_K12_28, u1_K12_29, u1_K12_30, u1_K12_31, u1_K12_32, u1_K12_35, u1_K12_36, 
       u1_K12_37, u1_K12_38, u1_K12_41, u1_K12_42, u1_K12_43, u1_K12_44, u1_K12_47, u1_K12_48, u1_K12_5, 
       u1_K12_6, u1_K12_7, u1_K12_8, u1_K12_9, u1_K13_1, u1_K13_12, u1_K13_14, u1_K13_17, u1_K13_18, 
       u1_K13_19, u1_K13_2, u1_K13_20, u1_K13_21, u1_K13_22, u1_K13_23, u1_K13_24, u1_K13_25, u1_K13_26, 
       u1_K13_27, u1_K13_28, u1_K13_29, u1_K13_3, u1_K13_30, u1_K13_31, u1_K13_32, u1_K13_35, u1_K13_36, 
       u1_K13_37, u1_K13_38, u1_K13_4, u1_K13_41, u1_K13_42, u1_K13_43, u1_K13_44, u1_K13_47, u1_K13_48, 
       u1_K13_5, u1_K13_6, u1_K13_7, u1_K13_8, u1_K14_1, u1_K14_10, u1_K14_11, u1_K14_12, u1_K14_13, 
       u1_K14_14, u1_K14_17, u1_K14_18, u1_K14_19, u1_K14_2, u1_K14_20, u1_K14_23, u1_K14_24, u1_K14_25, 
       u1_K14_26, u1_K14_27, u1_K14_28, u1_K14_29, u1_K14_30, u1_K14_31, u1_K14_32, u1_K14_35, u1_K14_36, 
       u1_K14_37, u1_K14_38, u1_K14_39, u1_K14_40, u1_K14_41, u1_K14_42, u1_K14_43, u1_K14_44, u1_K14_45, 
       u1_K14_46, u1_K14_47, u1_K14_48, u1_K14_5, u1_K14_6, u1_K14_7, u1_K14_8, u1_K14_9, u1_K15_1, 
       u1_K15_11, u1_K15_12, u1_K15_13, u1_K15_14, u1_K15_15, u1_K15_16, u1_K15_17, u1_K15_18, u1_K15_19, 
       u1_K15_2, u1_K15_20, u1_K15_23, u1_K15_24, u1_K15_25, u1_K15_26, u1_K15_29, u1_K15_30, u1_K15_31, 
       u1_K15_32, u1_K15_33, u1_K15_34, u1_K15_35, u1_K15_36, u1_K15_37, u1_K15_38, u1_K15_39, u1_K15_40, 
       u1_K15_41, u1_K15_42, u1_K15_43, u1_K15_44, u1_K15_45, u1_K15_46, u1_K15_47, u1_K15_48, u1_K15_5, 
       u1_K15_6, u1_K15_7, u1_K15_8, u1_K16_1, u1_K16_11, u1_K16_12, u1_K16_13, u1_K16_14, u1_K16_17, 
       u1_K16_18, u1_K16_19, u1_K16_2, u1_K16_20, u1_K16_21, u1_K16_22, u1_K16_23, u1_K16_24, u1_K16_25, 
       u1_K16_26, u1_K16_27, u1_K16_28, u1_K16_29, u1_K16_30, u1_K16_31, u1_K16_32, u1_K16_35, u1_K16_36, 
       u1_K16_37, u1_K16_38, u1_K16_41, u1_K16_42, u1_K16_43, u1_K16_44, u1_K16_47, u1_K16_48, u1_K16_5, 
       u1_K16_6, u1_K16_7, u1_K16_8, u1_K1_1, u1_K1_10, u1_K1_11, u1_K1_12, u1_K1_13, u1_K1_14, 
       u1_K1_17, u1_K1_18, u1_K1_19, u1_K1_2, u1_K1_20, u1_K1_21, u1_K1_22, u1_K1_23, u1_K1_24, 
       u1_K1_25, u1_K1_26, u1_K1_3, u1_K1_30, u1_K1_32, u1_K1_35, u1_K1_36, u1_K1_37, u1_K1_38, 
       u1_K1_39, u1_K1_4, u1_K1_40, u1_K1_41, u1_K1_42, u1_K1_43, u1_K1_44, u1_K1_45, u1_K1_46, 
       u1_K1_47, u1_K1_48, u1_K1_5, u1_K1_6, u1_K1_7, u1_K1_8, u1_K1_9, u1_K2_1, u1_K2_11, 
       u1_K2_12, u1_K2_13, u1_K2_14, u1_K2_15, u1_K2_16, u1_K2_17, u1_K2_18, u1_K2_19, u1_K2_2, 
       u1_K2_20, u1_K2_21, u1_K2_22, u1_K2_23, u1_K2_24, u1_K2_25, u1_K2_26, u1_K2_27, u1_K2_28, 
       u1_K2_29, u1_K2_3, u1_K2_30, u1_K2_31, u1_K2_32, u1_K2_35, u1_K2_36, u1_K2_37, u1_K2_38, 
       u1_K2_39, u1_K2_4, u1_K2_40, u1_K2_41, u1_K2_42, u1_K2_43, u1_K2_44, u1_K2_45, u1_K2_46, 
       u1_K2_47, u1_K2_48, u1_K2_5, u1_K2_6, u1_K2_7, u1_K2_8, u1_K3_1, u1_K3_11, u1_K3_12, 
       u1_K3_13, u1_K3_14, u1_K3_17, u1_K3_18, u1_K3_19, u1_K3_2, u1_K3_20, u1_K3_21, u1_K3_22, 
       u1_K3_23, u1_K3_24, u1_K3_25, u1_K3_26, u1_K3_29, u1_K3_30, u1_K3_31, u1_K3_32, u1_K3_35, 
       u1_K3_36, u1_K3_37, u1_K3_38, u1_K3_41, u1_K3_42, u1_K3_43, u1_K3_44, u1_K3_45, u1_K3_46, 
       u1_K3_47, u1_K3_48, u1_K3_5, u1_K3_6, u1_K3_7, u1_K3_8, u1_K4_1, u1_K4_11, u1_K4_12, 
       u1_K4_13, u1_K4_14, u1_K4_17, u1_K4_18, u1_K4_19, u1_K4_2, u1_K4_20, u1_K4_21, u1_K4_22, 
       u1_K4_23, u1_K4_24, u1_K4_25, u1_K4_26, u1_K4_35, u1_K4_36, u1_K4_37, u1_K4_38, u1_K4_41, 
       u1_K4_42, u1_K4_43, u1_K4_44, u1_K4_47, u1_K4_48, u1_K4_5, u1_K4_6, u1_K4_7, u1_K4_8, 
       u1_K5_1, u1_K5_11, u1_K5_12, u1_K5_13, u1_K5_14, u1_K5_17, u1_K5_18, u1_K5_19, u1_K5_2, 
       u1_K5_20, u1_K5_23, u1_K5_24, u1_K5_25, u1_K5_26, u1_K5_29, u1_K5_30, u1_K5_31, u1_K5_32, 
       u1_K5_33, u1_K5_34, u1_K5_35, u1_K5_36, u1_K5_37, u1_K5_38, u1_K5_41, u1_K5_42, u1_K5_43, 
       u1_K5_44, u1_K5_45, u1_K5_46, u1_K5_47, u1_K5_48, u1_K5_6, u1_K5_8, u1_K6_1, u1_K6_11, 
       u1_K6_12, u1_K6_13, u1_K6_14, u1_K6_15, u1_K6_16, u1_K6_17, u1_K6_18, u1_K6_19, u1_K6_2, 
       u1_K6_20, u1_K6_21, u1_K6_22, u1_K6_23, u1_K6_24, u1_K6_25, u1_K6_26, u1_K6_3, u1_K6_30, 
       u1_K6_32, u1_K6_35, u1_K6_36, u1_K6_37, u1_K6_38, u1_K6_39, u1_K6_4, u1_K6_40, u1_K6_41, 
       u1_K6_42, u1_K6_43, u1_K6_44, u1_K6_47, u1_K6_48, u1_K6_5, u1_K6_6, u1_K6_7, u1_K6_8, 
       u1_K7_1, u1_K7_11, u1_K7_12, u1_K7_13, u1_K7_14, u1_K7_15, u1_K7_16, u1_K7_17, u1_K7_18, 
       u1_K7_19, u1_K7_2, u1_K7_20, u1_K7_21, u1_K7_22, u1_K7_23, u1_K7_24, u1_K7_25, u1_K7_26, 
       u1_K7_29, u1_K7_30, u1_K7_31, u1_K7_32, u1_K7_35, u1_K7_36, u1_K7_37, u1_K7_38, u1_K7_41, 
       u1_K7_42, u1_K7_43, u1_K7_44, u1_K7_47, u1_K7_48, u1_K7_5, u1_K7_6, u1_K7_7, u1_K7_8, 
       u1_K8_1, u1_K8_10, u1_K8_11, u1_K8_12, u1_K8_13, u1_K8_14, u1_K8_15, u1_K8_16, u1_K8_17, 
       u1_K8_18, u1_K8_19, u1_K8_2, u1_K8_20, u1_K8_23, u1_K8_24, u1_K8_25, u1_K8_26, u1_K8_27, 
       u1_K8_28, u1_K8_29, u1_K8_3, u1_K8_30, u1_K8_31, u1_K8_32, u1_K8_35, u1_K8_36, u1_K8_37, 
       u1_K8_38, u1_K8_39, u1_K8_4, u1_K8_40, u1_K8_41, u1_K8_42, u1_K8_43, u1_K8_44, u1_K8_47, 
       u1_K8_48, u1_K8_5, u1_K8_6, u1_K8_7, u1_K8_8, u1_K8_9, u1_K9_1, u1_K9_10, u1_K9_11, 
       u1_K9_12, u1_K9_13, u1_K9_14, u1_K9_15, u1_K9_16, u1_K9_17, u1_K9_18, u1_K9_19, u1_K9_2, 
       u1_K9_20, u1_K9_21, u1_K9_22, u1_K9_23, u1_K9_24, u1_K9_25, u1_K9_26, u1_K9_29, u1_K9_30, 
       u1_K9_31, u1_K9_32, u1_K9_35, u1_K9_36, u1_K9_37, u1_K9_38, u1_K9_39, u1_K9_40, u1_K9_41, 
       u1_K9_42, u1_K9_43, u1_K9_44, u1_K9_45, u1_K9_46, u1_K9_47, u1_K9_48, u1_K9_5, u1_K9_6, 
       u1_K9_7, u1_K9_8, u1_K9_9, u1_out0_1, u1_out0_10, u1_out0_12, u1_out0_13, u1_out0_15, u1_out0_17, 
       u1_out0_18, u1_out0_2, u1_out0_20, u1_out0_21, u1_out0_22, u1_out0_23, u1_out0_26, u1_out0_27, u1_out0_28, 
       u1_out0_31, u1_out0_32, u1_out0_5, u1_out0_7, u1_out0_9, u1_out10_12, u1_out10_22, u1_out10_32, u1_out10_7, 
       u1_out11_1, u1_out11_10, u1_out11_13, u1_out11_14, u1_out11_16, u1_out11_18, u1_out11_2, u1_out11_20, u1_out11_24, 
       u1_out11_25, u1_out11_26, u1_out11_28, u1_out11_3, u1_out11_30, u1_out11_6, u1_out11_8, u1_out12_1, u1_out12_10, 
       u1_out12_14, u1_out12_17, u1_out12_20, u1_out12_23, u1_out12_25, u1_out12_26, u1_out12_3, u1_out12_31, u1_out12_8, 
       u1_out12_9, u1_out13_12, u1_out13_13, u1_out13_14, u1_out13_15, u1_out13_18, u1_out13_2, u1_out13_21, u1_out13_22, 
       u1_out13_25, u1_out13_27, u1_out13_28, u1_out13_3, u1_out13_32, u1_out13_5, u1_out13_7, u1_out13_8, u1_out14_11, 
       u1_out14_12, u1_out14_15, u1_out14_16, u1_out14_19, u1_out14_21, u1_out14_22, u1_out14_24, u1_out14_27, u1_out14_29, 
       u1_out14_30, u1_out14_32, u1_out14_4, u1_out14_5, u1_out14_6, u1_out14_7, u1_out15_1, u1_out15_10, u1_out15_14, 
       u1_out15_20, u1_out15_25, u1_out15_26, u1_out15_3, u1_out15_8, u1_out1_1, u1_out1_10, u1_out1_12, u1_out1_14, 
       u1_out1_15, u1_out1_16, u1_out1_17, u1_out1_20, u1_out1_21, u1_out1_22, u1_out1_23, u1_out1_24, u1_out1_25, 
       u1_out1_26, u1_out1_27, u1_out1_3, u1_out1_30, u1_out1_31, u1_out1_32, u1_out1_5, u1_out1_6, u1_out1_7, 
       u1_out1_8, u1_out1_9, u1_out2_1, u1_out2_10, u1_out2_15, u1_out2_20, u1_out2_21, u1_out2_26, u1_out2_27, 
       u1_out2_5, u1_out3_1, u1_out3_10, u1_out3_20, u1_out3_26, u1_out4_11, u1_out4_15, u1_out4_19, u1_out4_21, 
       u1_out4_27, u1_out4_29, u1_out4_4, u1_out4_5, u1_out5_1, u1_out5_10, u1_out5_12, u1_out5_16, u1_out5_17, 
       u1_out5_20, u1_out5_22, u1_out5_23, u1_out5_24, u1_out5_26, u1_out5_30, u1_out5_31, u1_out5_32, u1_out5_6, 
       u1_out5_7, u1_out5_9, u1_out6_1, u1_out6_10, u1_out6_16, u1_out6_20, u1_out6_24, u1_out6_26, u1_out6_30, 
       u1_out6_6, u1_out7_12, u1_out7_13, u1_out7_14, u1_out7_16, u1_out7_17, u1_out7_18, u1_out7_2, u1_out7_22, 
       u1_out7_23, u1_out7_24, u1_out7_25, u1_out7_28, u1_out7_3, u1_out7_30, u1_out7_31, u1_out7_32, u1_out7_6, 
       u1_out7_7, u1_out7_8, u1_out7_9, u1_out8_1, u1_out8_10, u1_out8_12, u1_out8_13, u1_out8_15, u1_out8_16, 
       u1_out8_18, u1_out8_2, u1_out8_20, u1_out8_21, u1_out8_22, u1_out8_24, u1_out8_26, u1_out8_27, u1_out8_28, 
       u1_out8_30, u1_out8_32, u1_out8_5, u1_out8_6, u1_out8_7, u1_out9_15, u1_out9_17, u1_out9_21, u1_out9_23, 
       u1_out9_27, u1_out9_31, u1_out9_5, u1_out9_9, u1_u0_X_1, u1_u0_X_10, u1_u0_X_11, u1_u0_X_12, u1_u0_X_19, 
       u1_u0_X_2, u1_u0_X_20, u1_u0_X_21, u1_u0_X_22, u1_u0_X_23, u1_u0_X_24, u1_u0_X_3, u1_u0_X_37, u1_u0_X_38, 
       u1_u0_X_39, u1_u0_X_4, u1_u0_X_40, u1_u0_X_41, u1_u0_X_42, u1_u0_X_43, u1_u0_X_44, u1_u0_X_45, u1_u0_X_46, 
       u1_u0_X_47, u1_u0_X_48, u1_u0_X_5, u1_u0_X_6, u1_u0_X_7, u1_u0_X_8, u1_u0_X_9, u1_u0_u0_n100, u1_u0_u0_n101, 
       u1_u0_u0_n102, u1_u0_u0_n103, u1_u0_u0_n104, u1_u0_u0_n105, u1_u0_u0_n106, u1_u0_u0_n107, u1_u0_u0_n108, u1_u0_u0_n109, u1_u0_u0_n110, 
       u1_u0_u0_n111, u1_u0_u0_n112, u1_u0_u0_n113, u1_u0_u0_n114, u1_u0_u0_n115, u1_u0_u0_n116, u1_u0_u0_n117, u1_u0_u0_n118, u1_u0_u0_n119, 
       u1_u0_u0_n120, u1_u0_u0_n121, u1_u0_u0_n122, u1_u0_u0_n123, u1_u0_u0_n124, u1_u0_u0_n125, u1_u0_u0_n126, u1_u0_u0_n127, u1_u0_u0_n128, 
       u1_u0_u0_n129, u1_u0_u0_n130, u1_u0_u0_n131, u1_u0_u0_n132, u1_u0_u0_n133, u1_u0_u0_n134, u1_u0_u0_n135, u1_u0_u0_n136, u1_u0_u0_n137, 
       u1_u0_u0_n138, u1_u0_u0_n139, u1_u0_u0_n140, u1_u0_u0_n141, u1_u0_u0_n142, u1_u0_u0_n143, u1_u0_u0_n144, u1_u0_u0_n145, u1_u0_u0_n146, 
       u1_u0_u0_n147, u1_u0_u0_n148, u1_u0_u0_n149, u1_u0_u0_n150, u1_u0_u0_n151, u1_u0_u0_n152, u1_u0_u0_n153, u1_u0_u0_n154, u1_u0_u0_n155, 
       u1_u0_u0_n156, u1_u0_u0_n157, u1_u0_u0_n158, u1_u0_u0_n159, u1_u0_u0_n160, u1_u0_u0_n161, u1_u0_u0_n162, u1_u0_u0_n163, u1_u0_u0_n164, 
       u1_u0_u0_n165, u1_u0_u0_n166, u1_u0_u0_n167, u1_u0_u0_n168, u1_u0_u0_n169, u1_u0_u0_n170, u1_u0_u0_n171, u1_u0_u0_n172, u1_u0_u0_n173, 
       u1_u0_u0_n174, u1_u0_u0_n88, u1_u0_u0_n89, u1_u0_u0_n90, u1_u0_u0_n91, u1_u0_u0_n92, u1_u0_u0_n93, u1_u0_u0_n94, u1_u0_u0_n95, 
       u1_u0_u0_n96, u1_u0_u0_n97, u1_u0_u0_n98, u1_u0_u0_n99, u1_u0_u1_n100, u1_u0_u1_n101, u1_u0_u1_n102, u1_u0_u1_n103, u1_u0_u1_n104, 
       u1_u0_u1_n105, u1_u0_u1_n106, u1_u0_u1_n107, u1_u0_u1_n108, u1_u0_u1_n109, u1_u0_u1_n110, u1_u0_u1_n111, u1_u0_u1_n112, u1_u0_u1_n113, 
       u1_u0_u1_n114, u1_u0_u1_n115, u1_u0_u1_n116, u1_u0_u1_n117, u1_u0_u1_n118, u1_u0_u1_n119, u1_u0_u1_n120, u1_u0_u1_n121, u1_u0_u1_n122, 
       u1_u0_u1_n123, u1_u0_u1_n124, u1_u0_u1_n125, u1_u0_u1_n126, u1_u0_u1_n127, u1_u0_u1_n128, u1_u0_u1_n129, u1_u0_u1_n130, u1_u0_u1_n131, 
       u1_u0_u1_n132, u1_u0_u1_n133, u1_u0_u1_n134, u1_u0_u1_n135, u1_u0_u1_n136, u1_u0_u1_n137, u1_u0_u1_n138, u1_u0_u1_n139, u1_u0_u1_n140, 
       u1_u0_u1_n141, u1_u0_u1_n142, u1_u0_u1_n143, u1_u0_u1_n144, u1_u0_u1_n145, u1_u0_u1_n146, u1_u0_u1_n147, u1_u0_u1_n148, u1_u0_u1_n149, 
       u1_u0_u1_n150, u1_u0_u1_n151, u1_u0_u1_n152, u1_u0_u1_n153, u1_u0_u1_n154, u1_u0_u1_n155, u1_u0_u1_n156, u1_u0_u1_n157, u1_u0_u1_n158, 
       u1_u0_u1_n159, u1_u0_u1_n160, u1_u0_u1_n161, u1_u0_u1_n162, u1_u0_u1_n163, u1_u0_u1_n164, u1_u0_u1_n165, u1_u0_u1_n166, u1_u0_u1_n167, 
       u1_u0_u1_n168, u1_u0_u1_n169, u1_u0_u1_n170, u1_u0_u1_n171, u1_u0_u1_n172, u1_u0_u1_n173, u1_u0_u1_n174, u1_u0_u1_n175, u1_u0_u1_n176, 
       u1_u0_u1_n177, u1_u0_u1_n178, u1_u0_u1_n179, u1_u0_u1_n180, u1_u0_u1_n181, u1_u0_u1_n182, u1_u0_u1_n183, u1_u0_u1_n184, u1_u0_u1_n185, 
       u1_u0_u1_n186, u1_u0_u1_n187, u1_u0_u1_n188, u1_u0_u1_n95, u1_u0_u1_n96, u1_u0_u1_n97, u1_u0_u1_n98, u1_u0_u1_n99, u1_u0_u3_n100, 
       u1_u0_u3_n101, u1_u0_u3_n102, u1_u0_u3_n103, u1_u0_u3_n104, u1_u0_u3_n105, u1_u0_u3_n106, u1_u0_u3_n107, u1_u0_u3_n108, u1_u0_u3_n109, 
       u1_u0_u3_n110, u1_u0_u3_n111, u1_u0_u3_n112, u1_u0_u3_n113, u1_u0_u3_n114, u1_u0_u3_n115, u1_u0_u3_n116, u1_u0_u3_n117, u1_u0_u3_n118, 
       u1_u0_u3_n119, u1_u0_u3_n120, u1_u0_u3_n121, u1_u0_u3_n122, u1_u0_u3_n123, u1_u0_u3_n124, u1_u0_u3_n125, u1_u0_u3_n126, u1_u0_u3_n127, 
       u1_u0_u3_n128, u1_u0_u3_n129, u1_u0_u3_n130, u1_u0_u3_n131, u1_u0_u3_n132, u1_u0_u3_n133, u1_u0_u3_n134, u1_u0_u3_n135, u1_u0_u3_n136, 
       u1_u0_u3_n137, u1_u0_u3_n138, u1_u0_u3_n139, u1_u0_u3_n140, u1_u0_u3_n141, u1_u0_u3_n142, u1_u0_u3_n143, u1_u0_u3_n144, u1_u0_u3_n145, 
       u1_u0_u3_n146, u1_u0_u3_n147, u1_u0_u3_n148, u1_u0_u3_n149, u1_u0_u3_n150, u1_u0_u3_n151, u1_u0_u3_n152, u1_u0_u3_n153, u1_u0_u3_n154, 
       u1_u0_u3_n155, u1_u0_u3_n156, u1_u0_u3_n157, u1_u0_u3_n158, u1_u0_u3_n159, u1_u0_u3_n160, u1_u0_u3_n161, u1_u0_u3_n162, u1_u0_u3_n163, 
       u1_u0_u3_n164, u1_u0_u3_n165, u1_u0_u3_n166, u1_u0_u3_n167, u1_u0_u3_n168, u1_u0_u3_n169, u1_u0_u3_n170, u1_u0_u3_n171, u1_u0_u3_n172, 
       u1_u0_u3_n173, u1_u0_u3_n174, u1_u0_u3_n175, u1_u0_u3_n176, u1_u0_u3_n177, u1_u0_u3_n178, u1_u0_u3_n179, u1_u0_u3_n180, u1_u0_u3_n181, 
       u1_u0_u3_n182, u1_u0_u3_n183, u1_u0_u3_n184, u1_u0_u3_n185, u1_u0_u3_n186, u1_u0_u3_n94, u1_u0_u3_n95, u1_u0_u3_n96, u1_u0_u3_n97, 
       u1_u0_u3_n98, u1_u0_u3_n99, u1_u0_u6_n100, u1_u0_u6_n101, u1_u0_u6_n102, u1_u0_u6_n103, u1_u0_u6_n104, u1_u0_u6_n105, u1_u0_u6_n106, 
       u1_u0_u6_n107, u1_u0_u6_n108, u1_u0_u6_n109, u1_u0_u6_n110, u1_u0_u6_n111, u1_u0_u6_n112, u1_u0_u6_n113, u1_u0_u6_n114, u1_u0_u6_n115, 
       u1_u0_u6_n116, u1_u0_u6_n117, u1_u0_u6_n118, u1_u0_u6_n119, u1_u0_u6_n120, u1_u0_u6_n121, u1_u0_u6_n122, u1_u0_u6_n123, u1_u0_u6_n124, 
       u1_u0_u6_n125, u1_u0_u6_n126, u1_u0_u6_n127, u1_u0_u6_n128, u1_u0_u6_n129, u1_u0_u6_n130, u1_u0_u6_n131, u1_u0_u6_n132, u1_u0_u6_n133, 
       u1_u0_u6_n134, u1_u0_u6_n135, u1_u0_u6_n136, u1_u0_u6_n137, u1_u0_u6_n138, u1_u0_u6_n139, u1_u0_u6_n140, u1_u0_u6_n141, u1_u0_u6_n142, 
       u1_u0_u6_n143, u1_u0_u6_n144, u1_u0_u6_n145, u1_u0_u6_n146, u1_u0_u6_n147, u1_u0_u6_n148, u1_u0_u6_n149, u1_u0_u6_n150, u1_u0_u6_n151, 
       u1_u0_u6_n152, u1_u0_u6_n153, u1_u0_u6_n154, u1_u0_u6_n155, u1_u0_u6_n156, u1_u0_u6_n157, u1_u0_u6_n158, u1_u0_u6_n159, u1_u0_u6_n160, 
       u1_u0_u6_n161, u1_u0_u6_n162, u1_u0_u6_n163, u1_u0_u6_n164, u1_u0_u6_n165, u1_u0_u6_n166, u1_u0_u6_n167, u1_u0_u6_n168, u1_u0_u6_n169, 
       u1_u0_u6_n170, u1_u0_u6_n171, u1_u0_u6_n172, u1_u0_u6_n173, u1_u0_u6_n174, u1_u0_u6_n88, u1_u0_u6_n89, u1_u0_u6_n90, u1_u0_u6_n91, 
       u1_u0_u6_n92, u1_u0_u6_n93, u1_u0_u6_n94, u1_u0_u6_n95, u1_u0_u6_n96, u1_u0_u6_n97, u1_u0_u6_n98, u1_u0_u6_n99, u1_u0_u7_n100, 
       u1_u0_u7_n101, u1_u0_u7_n102, u1_u0_u7_n103, u1_u0_u7_n104, u1_u0_u7_n105, u1_u0_u7_n106, u1_u0_u7_n107, u1_u0_u7_n108, u1_u0_u7_n109, 
       u1_u0_u7_n110, u1_u0_u7_n111, u1_u0_u7_n112, u1_u0_u7_n113, u1_u0_u7_n114, u1_u0_u7_n115, u1_u0_u7_n116, u1_u0_u7_n117, u1_u0_u7_n118, 
       u1_u0_u7_n119, u1_u0_u7_n120, u1_u0_u7_n121, u1_u0_u7_n122, u1_u0_u7_n123, u1_u0_u7_n124, u1_u0_u7_n125, u1_u0_u7_n126, u1_u0_u7_n127, 
       u1_u0_u7_n128, u1_u0_u7_n129, u1_u0_u7_n130, u1_u0_u7_n131, u1_u0_u7_n132, u1_u0_u7_n133, u1_u0_u7_n134, u1_u0_u7_n135, u1_u0_u7_n136, 
       u1_u0_u7_n137, u1_u0_u7_n138, u1_u0_u7_n139, u1_u0_u7_n140, u1_u0_u7_n141, u1_u0_u7_n142, u1_u0_u7_n143, u1_u0_u7_n144, u1_u0_u7_n145, 
       u1_u0_u7_n146, u1_u0_u7_n147, u1_u0_u7_n148, u1_u0_u7_n149, u1_u0_u7_n150, u1_u0_u7_n151, u1_u0_u7_n152, u1_u0_u7_n153, u1_u0_u7_n154, 
       u1_u0_u7_n155, u1_u0_u7_n156, u1_u0_u7_n157, u1_u0_u7_n158, u1_u0_u7_n159, u1_u0_u7_n160, u1_u0_u7_n161, u1_u0_u7_n162, u1_u0_u7_n163, 
       u1_u0_u7_n164, u1_u0_u7_n165, u1_u0_u7_n166, u1_u0_u7_n167, u1_u0_u7_n168, u1_u0_u7_n169, u1_u0_u7_n170, u1_u0_u7_n171, u1_u0_u7_n172, 
       u1_u0_u7_n173, u1_u0_u7_n174, u1_u0_u7_n175, u1_u0_u7_n176, u1_u0_u7_n177, u1_u0_u7_n178, u1_u0_u7_n179, u1_u0_u7_n180, u1_u0_u7_n91, 
       u1_u0_u7_n92, u1_u0_u7_n93, u1_u0_u7_n94, u1_u0_u7_n95, u1_u0_u7_n96, u1_u0_u7_n97, u1_u0_u7_n98, u1_u0_u7_n99, u1_u10_X_37, 
       u1_u10_X_38, u1_u10_X_39, u1_u10_X_40, u1_u10_X_41, u1_u10_X_42, u1_u10_u6_n100, u1_u10_u6_n101, u1_u10_u6_n102, u1_u10_u6_n103, 
       u1_u10_u6_n104, u1_u10_u6_n105, u1_u10_u6_n106, u1_u10_u6_n107, u1_u10_u6_n108, u1_u10_u6_n109, u1_u10_u6_n110, u1_u10_u6_n111, u1_u10_u6_n112, 
       u1_u10_u6_n113, u1_u10_u6_n114, u1_u10_u6_n115, u1_u10_u6_n116, u1_u10_u6_n117, u1_u10_u6_n118, u1_u10_u6_n119, u1_u10_u6_n120, u1_u10_u6_n121, 
       u1_u10_u6_n122, u1_u10_u6_n123, u1_u10_u6_n124, u1_u10_u6_n125, u1_u10_u6_n126, u1_u10_u6_n127, u1_u10_u6_n128, u1_u10_u6_n129, u1_u10_u6_n130, 
       u1_u10_u6_n131, u1_u10_u6_n132, u1_u10_u6_n133, u1_u10_u6_n134, u1_u10_u6_n135, u1_u10_u6_n136, u1_u10_u6_n137, u1_u10_u6_n138, u1_u10_u6_n139, 
       u1_u10_u6_n140, u1_u10_u6_n141, u1_u10_u6_n142, u1_u10_u6_n143, u1_u10_u6_n144, u1_u10_u6_n145, u1_u10_u6_n146, u1_u10_u6_n147, u1_u10_u6_n148, 
       u1_u10_u6_n149, u1_u10_u6_n150, u1_u10_u6_n151, u1_u10_u6_n152, u1_u10_u6_n153, u1_u10_u6_n154, u1_u10_u6_n155, u1_u10_u6_n156, u1_u10_u6_n157, 
       u1_u10_u6_n158, u1_u10_u6_n159, u1_u10_u6_n160, u1_u10_u6_n161, u1_u10_u6_n162, u1_u10_u6_n163, u1_u10_u6_n164, u1_u10_u6_n165, u1_u10_u6_n166, 
       u1_u10_u6_n167, u1_u10_u6_n168, u1_u10_u6_n169, u1_u10_u6_n170, u1_u10_u6_n171, u1_u10_u6_n172, u1_u10_u6_n173, u1_u10_u6_n174, u1_u10_u6_n88, 
       u1_u10_u6_n89, u1_u10_u6_n90, u1_u10_u6_n91, u1_u10_u6_n92, u1_u10_u6_n93, u1_u10_u6_n94, u1_u10_u6_n95, u1_u10_u6_n96, u1_u10_u6_n97, 
       u1_u10_u6_n98, u1_u10_u6_n99, u1_u11_X_10, u1_u11_X_11, u1_u11_X_12, u1_u11_X_13, u1_u11_X_14, u1_u11_X_15, u1_u11_X_16, 
       u1_u11_X_17, u1_u11_X_18, u1_u11_X_19, u1_u11_X_20, u1_u11_X_21, u1_u11_X_22, u1_u11_X_23, u1_u11_X_24, u1_u11_X_25, 
       u1_u11_X_26, u1_u11_X_27, u1_u11_X_28, u1_u11_X_29, u1_u11_X_30, u1_u11_X_7, u1_u11_X_8, u1_u11_X_9, u1_u11_u1_n100, 
       u1_u11_u1_n101, u1_u11_u1_n102, u1_u11_u1_n103, u1_u11_u1_n104, u1_u11_u1_n105, u1_u11_u1_n106, u1_u11_u1_n107, u1_u11_u1_n108, u1_u11_u1_n109, 
       u1_u11_u1_n110, u1_u11_u1_n111, u1_u11_u1_n112, u1_u11_u1_n113, u1_u11_u1_n114, u1_u11_u1_n115, u1_u11_u1_n116, u1_u11_u1_n117, u1_u11_u1_n118, 
       u1_u11_u1_n119, u1_u11_u1_n120, u1_u11_u1_n121, u1_u11_u1_n122, u1_u11_u1_n123, u1_u11_u1_n124, u1_u11_u1_n125, u1_u11_u1_n126, u1_u11_u1_n127, 
       u1_u11_u1_n128, u1_u11_u1_n129, u1_u11_u1_n130, u1_u11_u1_n131, u1_u11_u1_n132, u1_u11_u1_n133, u1_u11_u1_n134, u1_u11_u1_n135, u1_u11_u1_n136, 
       u1_u11_u1_n137, u1_u11_u1_n138, u1_u11_u1_n139, u1_u11_u1_n140, u1_u11_u1_n141, u1_u11_u1_n142, u1_u11_u1_n143, u1_u11_u1_n144, u1_u11_u1_n145, 
       u1_u11_u1_n146, u1_u11_u1_n147, u1_u11_u1_n148, u1_u11_u1_n149, u1_u11_u1_n150, u1_u11_u1_n151, u1_u11_u1_n152, u1_u11_u1_n153, u1_u11_u1_n154, 
       u1_u11_u1_n155, u1_u11_u1_n156, u1_u11_u1_n157, u1_u11_u1_n158, u1_u11_u1_n159, u1_u11_u1_n160, u1_u11_u1_n161, u1_u11_u1_n162, u1_u11_u1_n163, 
       u1_u11_u1_n164, u1_u11_u1_n165, u1_u11_u1_n166, u1_u11_u1_n167, u1_u11_u1_n168, u1_u11_u1_n169, u1_u11_u1_n170, u1_u11_u1_n171, u1_u11_u1_n172, 
       u1_u11_u1_n173, u1_u11_u1_n174, u1_u11_u1_n175, u1_u11_u1_n176, u1_u11_u1_n177, u1_u11_u1_n178, u1_u11_u1_n179, u1_u11_u1_n180, u1_u11_u1_n181, 
       u1_u11_u1_n182, u1_u11_u1_n183, u1_u11_u1_n184, u1_u11_u1_n185, u1_u11_u1_n186, u1_u11_u1_n187, u1_u11_u1_n188, u1_u11_u1_n95, u1_u11_u1_n96, 
       u1_u11_u1_n97, u1_u11_u1_n98, u1_u11_u1_n99, u1_u11_u2_n100, u1_u11_u2_n101, u1_u11_u2_n102, u1_u11_u2_n103, u1_u11_u2_n104, u1_u11_u2_n105, 
       u1_u11_u2_n106, u1_u11_u2_n107, u1_u11_u2_n108, u1_u11_u2_n109, u1_u11_u2_n110, u1_u11_u2_n111, u1_u11_u2_n112, u1_u11_u2_n113, u1_u11_u2_n114, 
       u1_u11_u2_n115, u1_u11_u2_n116, u1_u11_u2_n117, u1_u11_u2_n118, u1_u11_u2_n119, u1_u11_u2_n120, u1_u11_u2_n121, u1_u11_u2_n122, u1_u11_u2_n123, 
       u1_u11_u2_n124, u1_u11_u2_n125, u1_u11_u2_n126, u1_u11_u2_n127, u1_u11_u2_n128, u1_u11_u2_n129, u1_u11_u2_n130, u1_u11_u2_n131, u1_u11_u2_n132, 
       u1_u11_u2_n133, u1_u11_u2_n134, u1_u11_u2_n135, u1_u11_u2_n136, u1_u11_u2_n137, u1_u11_u2_n138, u1_u11_u2_n139, u1_u11_u2_n140, u1_u11_u2_n141, 
       u1_u11_u2_n142, u1_u11_u2_n143, u1_u11_u2_n144, u1_u11_u2_n145, u1_u11_u2_n146, u1_u11_u2_n147, u1_u11_u2_n148, u1_u11_u2_n149, u1_u11_u2_n150, 
       u1_u11_u2_n151, u1_u11_u2_n152, u1_u11_u2_n153, u1_u11_u2_n154, u1_u11_u2_n155, u1_u11_u2_n156, u1_u11_u2_n157, u1_u11_u2_n158, u1_u11_u2_n159, 
       u1_u11_u2_n160, u1_u11_u2_n161, u1_u11_u2_n162, u1_u11_u2_n163, u1_u11_u2_n164, u1_u11_u2_n165, u1_u11_u2_n166, u1_u11_u2_n167, u1_u11_u2_n168, 
       u1_u11_u2_n169, u1_u11_u2_n170, u1_u11_u2_n171, u1_u11_u2_n172, u1_u11_u2_n173, u1_u11_u2_n174, u1_u11_u2_n175, u1_u11_u2_n176, u1_u11_u2_n177, 
       u1_u11_u2_n178, u1_u11_u2_n179, u1_u11_u2_n180, u1_u11_u2_n181, u1_u11_u2_n182, u1_u11_u2_n183, u1_u11_u2_n184, u1_u11_u2_n185, u1_u11_u2_n186, 
       u1_u11_u2_n187, u1_u11_u2_n188, u1_u11_u2_n95, u1_u11_u2_n96, u1_u11_u2_n97, u1_u11_u2_n98, u1_u11_u2_n99, u1_u11_u3_n100, u1_u11_u3_n101, 
       u1_u11_u3_n102, u1_u11_u3_n103, u1_u11_u3_n104, u1_u11_u3_n105, u1_u11_u3_n106, u1_u11_u3_n107, u1_u11_u3_n108, u1_u11_u3_n109, u1_u11_u3_n110, 
       u1_u11_u3_n111, u1_u11_u3_n112, u1_u11_u3_n113, u1_u11_u3_n114, u1_u11_u3_n115, u1_u11_u3_n116, u1_u11_u3_n117, u1_u11_u3_n118, u1_u11_u3_n119, 
       u1_u11_u3_n120, u1_u11_u3_n121, u1_u11_u3_n122, u1_u11_u3_n123, u1_u11_u3_n124, u1_u11_u3_n125, u1_u11_u3_n126, u1_u11_u3_n127, u1_u11_u3_n128, 
       u1_u11_u3_n129, u1_u11_u3_n130, u1_u11_u3_n131, u1_u11_u3_n132, u1_u11_u3_n133, u1_u11_u3_n134, u1_u11_u3_n135, u1_u11_u3_n136, u1_u11_u3_n137, 
       u1_u11_u3_n138, u1_u11_u3_n139, u1_u11_u3_n140, u1_u11_u3_n141, u1_u11_u3_n142, u1_u11_u3_n143, u1_u11_u3_n144, u1_u11_u3_n145, u1_u11_u3_n146, 
       u1_u11_u3_n147, u1_u11_u3_n148, u1_u11_u3_n149, u1_u11_u3_n150, u1_u11_u3_n151, u1_u11_u3_n152, u1_u11_u3_n153, u1_u11_u3_n154, u1_u11_u3_n155, 
       u1_u11_u3_n156, u1_u11_u3_n157, u1_u11_u3_n158, u1_u11_u3_n159, u1_u11_u3_n160, u1_u11_u3_n161, u1_u11_u3_n162, u1_u11_u3_n163, u1_u11_u3_n164, 
       u1_u11_u3_n165, u1_u11_u3_n166, u1_u11_u3_n167, u1_u11_u3_n168, u1_u11_u3_n169, u1_u11_u3_n170, u1_u11_u3_n171, u1_u11_u3_n172, u1_u11_u3_n173, 
       u1_u11_u3_n174, u1_u11_u3_n175, u1_u11_u3_n176, u1_u11_u3_n177, u1_u11_u3_n178, u1_u11_u3_n179, u1_u11_u3_n180, u1_u11_u3_n181, u1_u11_u3_n182, 
       u1_u11_u3_n183, u1_u11_u3_n184, u1_u11_u3_n185, u1_u11_u3_n186, u1_u11_u3_n94, u1_u11_u3_n95, u1_u11_u3_n96, u1_u11_u3_n97, u1_u11_u3_n98, 
       u1_u11_u3_n99, u1_u11_u4_n100, u1_u11_u4_n101, u1_u11_u4_n102, u1_u11_u4_n103, u1_u11_u4_n104, u1_u11_u4_n105, u1_u11_u4_n106, u1_u11_u4_n107, 
       u1_u11_u4_n108, u1_u11_u4_n109, u1_u11_u4_n110, u1_u11_u4_n111, u1_u11_u4_n112, u1_u11_u4_n113, u1_u11_u4_n114, u1_u11_u4_n115, u1_u11_u4_n116, 
       u1_u11_u4_n117, u1_u11_u4_n118, u1_u11_u4_n119, u1_u11_u4_n120, u1_u11_u4_n121, u1_u11_u4_n122, u1_u11_u4_n123, u1_u11_u4_n124, u1_u11_u4_n125, 
       u1_u11_u4_n126, u1_u11_u4_n127, u1_u11_u4_n128, u1_u11_u4_n129, u1_u11_u4_n130, u1_u11_u4_n131, u1_u11_u4_n132, u1_u11_u4_n133, u1_u11_u4_n134, 
       u1_u11_u4_n135, u1_u11_u4_n136, u1_u11_u4_n137, u1_u11_u4_n138, u1_u11_u4_n139, u1_u11_u4_n140, u1_u11_u4_n141, u1_u11_u4_n142, u1_u11_u4_n143, 
       u1_u11_u4_n144, u1_u11_u4_n145, u1_u11_u4_n146, u1_u11_u4_n147, u1_u11_u4_n148, u1_u11_u4_n149, u1_u11_u4_n150, u1_u11_u4_n151, u1_u11_u4_n152, 
       u1_u11_u4_n153, u1_u11_u4_n154, u1_u11_u4_n155, u1_u11_u4_n156, u1_u11_u4_n157, u1_u11_u4_n158, u1_u11_u4_n159, u1_u11_u4_n160, u1_u11_u4_n161, 
       u1_u11_u4_n162, u1_u11_u4_n163, u1_u11_u4_n164, u1_u11_u4_n165, u1_u11_u4_n166, u1_u11_u4_n167, u1_u11_u4_n168, u1_u11_u4_n169, u1_u11_u4_n170, 
       u1_u11_u4_n171, u1_u11_u4_n172, u1_u11_u4_n173, u1_u11_u4_n174, u1_u11_u4_n175, u1_u11_u4_n176, u1_u11_u4_n177, u1_u11_u4_n178, u1_u11_u4_n179, 
       u1_u11_u4_n180, u1_u11_u4_n181, u1_u11_u4_n182, u1_u11_u4_n183, u1_u11_u4_n184, u1_u11_u4_n185, u1_u11_u4_n186, u1_u11_u4_n94, u1_u11_u4_n95, 
       u1_u11_u4_n96, u1_u11_u4_n97, u1_u11_u4_n98, u1_u11_u4_n99, u1_u12_X_1, u1_u12_X_19, u1_u12_X_2, u1_u12_X_20, u1_u12_X_21, 
       u1_u12_X_22, u1_u12_X_23, u1_u12_X_24, u1_u12_X_25, u1_u12_X_26, u1_u12_X_27, u1_u12_X_28, u1_u12_X_29, u1_u12_X_3, 
       u1_u12_X_30, u1_u12_X_4, u1_u12_X_5, u1_u12_X_6, u1_u12_u0_n100, u1_u12_u0_n101, u1_u12_u0_n102, u1_u12_u0_n103, u1_u12_u0_n104, 
       u1_u12_u0_n105, u1_u12_u0_n106, u1_u12_u0_n107, u1_u12_u0_n108, u1_u12_u0_n109, u1_u12_u0_n110, u1_u12_u0_n111, u1_u12_u0_n112, u1_u12_u0_n113, 
       u1_u12_u0_n114, u1_u12_u0_n115, u1_u12_u0_n116, u1_u12_u0_n117, u1_u12_u0_n118, u1_u12_u0_n119, u1_u12_u0_n120, u1_u12_u0_n121, u1_u12_u0_n122, 
       u1_u12_u0_n123, u1_u12_u0_n124, u1_u12_u0_n125, u1_u12_u0_n126, u1_u12_u0_n127, u1_u12_u0_n128, u1_u12_u0_n129, u1_u12_u0_n130, u1_u12_u0_n131, 
       u1_u12_u0_n132, u1_u12_u0_n133, u1_u12_u0_n134, u1_u12_u0_n135, u1_u12_u0_n136, u1_u12_u0_n137, u1_u12_u0_n138, u1_u12_u0_n139, u1_u12_u0_n140, 
       u1_u12_u0_n141, u1_u12_u0_n142, u1_u12_u0_n143, u1_u12_u0_n144, u1_u12_u0_n145, u1_u12_u0_n146, u1_u12_u0_n147, u1_u12_u0_n148, u1_u12_u0_n149, 
       u1_u12_u0_n150, u1_u12_u0_n151, u1_u12_u0_n152, u1_u12_u0_n153, u1_u12_u0_n154, u1_u12_u0_n155, u1_u12_u0_n156, u1_u12_u0_n157, u1_u12_u0_n158, 
       u1_u12_u0_n159, u1_u12_u0_n160, u1_u12_u0_n161, u1_u12_u0_n162, u1_u12_u0_n163, u1_u12_u0_n164, u1_u12_u0_n165, u1_u12_u0_n166, u1_u12_u0_n167, 
       u1_u12_u0_n168, u1_u12_u0_n169, u1_u12_u0_n170, u1_u12_u0_n171, u1_u12_u0_n172, u1_u12_u0_n173, u1_u12_u0_n174, u1_u12_u0_n88, u1_u12_u0_n89, 
       u1_u12_u0_n90, u1_u12_u0_n91, u1_u12_u0_n92, u1_u12_u0_n93, u1_u12_u0_n94, u1_u12_u0_n95, u1_u12_u0_n96, u1_u12_u0_n97, u1_u12_u0_n98, 
       u1_u12_u0_n99, u1_u12_u3_n100, u1_u12_u3_n101, u1_u12_u3_n102, u1_u12_u3_n103, u1_u12_u3_n104, u1_u12_u3_n105, u1_u12_u3_n106, u1_u12_u3_n107, 
       u1_u12_u3_n108, u1_u12_u3_n109, u1_u12_u3_n110, u1_u12_u3_n111, u1_u12_u3_n112, u1_u12_u3_n113, u1_u12_u3_n114, u1_u12_u3_n115, u1_u12_u3_n116, 
       u1_u12_u3_n117, u1_u12_u3_n118, u1_u12_u3_n119, u1_u12_u3_n120, u1_u12_u3_n121, u1_u12_u3_n122, u1_u12_u3_n123, u1_u12_u3_n124, u1_u12_u3_n125, 
       u1_u12_u3_n126, u1_u12_u3_n127, u1_u12_u3_n128, u1_u12_u3_n129, u1_u12_u3_n130, u1_u12_u3_n131, u1_u12_u3_n132, u1_u12_u3_n133, u1_u12_u3_n134, 
       u1_u12_u3_n135, u1_u12_u3_n136, u1_u12_u3_n137, u1_u12_u3_n138, u1_u12_u3_n139, u1_u12_u3_n140, u1_u12_u3_n141, u1_u12_u3_n142, u1_u12_u3_n143, 
       u1_u12_u3_n144, u1_u12_u3_n145, u1_u12_u3_n146, u1_u12_u3_n147, u1_u12_u3_n148, u1_u12_u3_n149, u1_u12_u3_n150, u1_u12_u3_n151, u1_u12_u3_n152, 
       u1_u12_u3_n153, u1_u12_u3_n154, u1_u12_u3_n155, u1_u12_u3_n156, u1_u12_u3_n157, u1_u12_u3_n158, u1_u12_u3_n159, u1_u12_u3_n160, u1_u12_u3_n161, 
       u1_u12_u3_n162, u1_u12_u3_n163, u1_u12_u3_n164, u1_u12_u3_n165, u1_u12_u3_n166, u1_u12_u3_n167, u1_u12_u3_n168, u1_u12_u3_n169, u1_u12_u3_n170, 
       u1_u12_u3_n171, u1_u12_u3_n172, u1_u12_u3_n173, u1_u12_u3_n174, u1_u12_u3_n175, u1_u12_u3_n176, u1_u12_u3_n177, u1_u12_u3_n178, u1_u12_u3_n179, 
       u1_u12_u3_n180, u1_u12_u3_n181, u1_u12_u3_n182, u1_u12_u3_n183, u1_u12_u3_n184, u1_u12_u3_n185, u1_u12_u3_n186, u1_u12_u3_n94, u1_u12_u3_n95, 
       u1_u12_u3_n96, u1_u12_u3_n97, u1_u12_u3_n98, u1_u12_u3_n99, u1_u12_u4_n100, u1_u12_u4_n101, u1_u12_u4_n102, u1_u12_u4_n103, u1_u12_u4_n104, 
       u1_u12_u4_n105, u1_u12_u4_n106, u1_u12_u4_n107, u1_u12_u4_n108, u1_u12_u4_n109, u1_u12_u4_n110, u1_u12_u4_n111, u1_u12_u4_n112, u1_u12_u4_n113, 
       u1_u12_u4_n114, u1_u12_u4_n115, u1_u12_u4_n116, u1_u12_u4_n117, u1_u12_u4_n118, u1_u12_u4_n119, u1_u12_u4_n120, u1_u12_u4_n121, u1_u12_u4_n122, 
       u1_u12_u4_n123, u1_u12_u4_n124, u1_u12_u4_n125, u1_u12_u4_n126, u1_u12_u4_n127, u1_u12_u4_n128, u1_u12_u4_n129, u1_u12_u4_n130, u1_u12_u4_n131, 
       u1_u12_u4_n132, u1_u12_u4_n133, u1_u12_u4_n134, u1_u12_u4_n135, u1_u12_u4_n136, u1_u12_u4_n137, u1_u12_u4_n138, u1_u12_u4_n139, u1_u12_u4_n140, 
       u1_u12_u4_n141, u1_u12_u4_n142, u1_u12_u4_n143, u1_u12_u4_n144, u1_u12_u4_n145, u1_u12_u4_n146, u1_u12_u4_n147, u1_u12_u4_n148, u1_u12_u4_n149, 
       u1_u12_u4_n150, u1_u12_u4_n151, u1_u12_u4_n152, u1_u12_u4_n153, u1_u12_u4_n154, u1_u12_u4_n155, u1_u12_u4_n156, u1_u12_u4_n157, u1_u12_u4_n158, 
       u1_u12_u4_n159, u1_u12_u4_n160, u1_u12_u4_n161, u1_u12_u4_n162, u1_u12_u4_n163, u1_u12_u4_n164, u1_u12_u4_n165, u1_u12_u4_n166, u1_u12_u4_n167, 
       u1_u12_u4_n168, u1_u12_u4_n169, u1_u12_u4_n170, u1_u12_u4_n171, u1_u12_u4_n172, u1_u12_u4_n173, u1_u12_u4_n174, u1_u12_u4_n175, u1_u12_u4_n176, 
       u1_u12_u4_n177, u1_u12_u4_n178, u1_u12_u4_n179, u1_u12_u4_n180, u1_u12_u4_n181, u1_u12_u4_n182, u1_u12_u4_n183, u1_u12_u4_n184, u1_u12_u4_n185, 
       u1_u12_u4_n186, u1_u12_u4_n94, u1_u12_u4_n95, u1_u12_u4_n96, u1_u12_u4_n97, u1_u12_u4_n98, u1_u12_u4_n99, u1_u13_X_10, u1_u13_X_11, 
       u1_u13_X_12, u1_u13_X_25, u1_u13_X_26, u1_u13_X_27, u1_u13_X_28, u1_u13_X_29, u1_u13_X_30, u1_u13_X_37, u1_u13_X_38, 
       u1_u13_X_39, u1_u13_X_40, u1_u13_X_41, u1_u13_X_42, u1_u13_X_43, u1_u13_X_44, u1_u13_X_45, u1_u13_X_46, u1_u13_X_47, 
       u1_u13_X_48, u1_u13_X_7, u1_u13_X_8, u1_u13_X_9, u1_u13_u1_n100, u1_u13_u1_n101, u1_u13_u1_n102, u1_u13_u1_n103, u1_u13_u1_n104, 
       u1_u13_u1_n105, u1_u13_u1_n106, u1_u13_u1_n107, u1_u13_u1_n108, u1_u13_u1_n109, u1_u13_u1_n110, u1_u13_u1_n111, u1_u13_u1_n112, u1_u13_u1_n113, 
       u1_u13_u1_n114, u1_u13_u1_n115, u1_u13_u1_n116, u1_u13_u1_n117, u1_u13_u1_n118, u1_u13_u1_n119, u1_u13_u1_n120, u1_u13_u1_n121, u1_u13_u1_n122, 
       u1_u13_u1_n123, u1_u13_u1_n124, u1_u13_u1_n125, u1_u13_u1_n126, u1_u13_u1_n127, u1_u13_u1_n128, u1_u13_u1_n129, u1_u13_u1_n130, u1_u13_u1_n131, 
       u1_u13_u1_n132, u1_u13_u1_n133, u1_u13_u1_n134, u1_u13_u1_n135, u1_u13_u1_n136, u1_u13_u1_n137, u1_u13_u1_n138, u1_u13_u1_n139, u1_u13_u1_n140, 
       u1_u13_u1_n141, u1_u13_u1_n142, u1_u13_u1_n143, u1_u13_u1_n144, u1_u13_u1_n145, u1_u13_u1_n146, u1_u13_u1_n147, u1_u13_u1_n148, u1_u13_u1_n149, 
       u1_u13_u1_n150, u1_u13_u1_n151, u1_u13_u1_n152, u1_u13_u1_n153, u1_u13_u1_n154, u1_u13_u1_n155, u1_u13_u1_n156, u1_u13_u1_n157, u1_u13_u1_n158, 
       u1_u13_u1_n159, u1_u13_u1_n160, u1_u13_u1_n161, u1_u13_u1_n162, u1_u13_u1_n163, u1_u13_u1_n164, u1_u13_u1_n165, u1_u13_u1_n166, u1_u13_u1_n167, 
       u1_u13_u1_n168, u1_u13_u1_n169, u1_u13_u1_n170, u1_u13_u1_n171, u1_u13_u1_n172, u1_u13_u1_n173, u1_u13_u1_n174, u1_u13_u1_n175, u1_u13_u1_n176, 
       u1_u13_u1_n177, u1_u13_u1_n178, u1_u13_u1_n179, u1_u13_u1_n180, u1_u13_u1_n181, u1_u13_u1_n182, u1_u13_u1_n183, u1_u13_u1_n184, u1_u13_u1_n185, 
       u1_u13_u1_n186, u1_u13_u1_n187, u1_u13_u1_n188, u1_u13_u1_n95, u1_u13_u1_n96, u1_u13_u1_n97, u1_u13_u1_n98, u1_u13_u1_n99, u1_u13_u4_n100, 
       u1_u13_u4_n101, u1_u13_u4_n102, u1_u13_u4_n103, u1_u13_u4_n104, u1_u13_u4_n105, u1_u13_u4_n106, u1_u13_u4_n107, u1_u13_u4_n108, u1_u13_u4_n109, 
       u1_u13_u4_n110, u1_u13_u4_n111, u1_u13_u4_n112, u1_u13_u4_n113, u1_u13_u4_n114, u1_u13_u4_n115, u1_u13_u4_n116, u1_u13_u4_n117, u1_u13_u4_n118, 
       u1_u13_u4_n119, u1_u13_u4_n120, u1_u13_u4_n121, u1_u13_u4_n122, u1_u13_u4_n123, u1_u13_u4_n124, u1_u13_u4_n125, u1_u13_u4_n126, u1_u13_u4_n127, 
       u1_u13_u4_n128, u1_u13_u4_n129, u1_u13_u4_n130, u1_u13_u4_n131, u1_u13_u4_n132, u1_u13_u4_n133, u1_u13_u4_n134, u1_u13_u4_n135, u1_u13_u4_n136, 
       u1_u13_u4_n137, u1_u13_u4_n138, u1_u13_u4_n139, u1_u13_u4_n140, u1_u13_u4_n141, u1_u13_u4_n142, u1_u13_u4_n143, u1_u13_u4_n144, u1_u13_u4_n145, 
       u1_u13_u4_n146, u1_u13_u4_n147, u1_u13_u4_n148, u1_u13_u4_n149, u1_u13_u4_n150, u1_u13_u4_n151, u1_u13_u4_n152, u1_u13_u4_n153, u1_u13_u4_n154, 
       u1_u13_u4_n155, u1_u13_u4_n156, u1_u13_u4_n157, u1_u13_u4_n158, u1_u13_u4_n159, u1_u13_u4_n160, u1_u13_u4_n161, u1_u13_u4_n162, u1_u13_u4_n163, 
       u1_u13_u4_n164, u1_u13_u4_n165, u1_u13_u4_n166, u1_u13_u4_n167, u1_u13_u4_n168, u1_u13_u4_n169, u1_u13_u4_n170, u1_u13_u4_n171, u1_u13_u4_n172, 
       u1_u13_u4_n173, u1_u13_u4_n174, u1_u13_u4_n175, u1_u13_u4_n176, u1_u13_u4_n177, u1_u13_u4_n178, u1_u13_u4_n179, u1_u13_u4_n180, u1_u13_u4_n181, 
       u1_u13_u4_n182, u1_u13_u4_n183, u1_u13_u4_n184, u1_u13_u4_n185, u1_u13_u4_n186, u1_u13_u4_n94, u1_u13_u4_n95, u1_u13_u4_n96, u1_u13_u4_n97, 
       u1_u13_u4_n98, u1_u13_u4_n99, u1_u13_u6_n100, u1_u13_u6_n101, u1_u13_u6_n102, u1_u13_u6_n103, u1_u13_u6_n104, u1_u13_u6_n105, u1_u13_u6_n106, 
       u1_u13_u6_n107, u1_u13_u6_n108, u1_u13_u6_n109, u1_u13_u6_n110, u1_u13_u6_n111, u1_u13_u6_n112, u1_u13_u6_n113, u1_u13_u6_n114, u1_u13_u6_n115, 
       u1_u13_u6_n116, u1_u13_u6_n117, u1_u13_u6_n118, u1_u13_u6_n119, u1_u13_u6_n120, u1_u13_u6_n121, u1_u13_u6_n122, u1_u13_u6_n123, u1_u13_u6_n124, 
       u1_u13_u6_n125, u1_u13_u6_n126, u1_u13_u6_n127, u1_u13_u6_n128, u1_u13_u6_n129, u1_u13_u6_n130, u1_u13_u6_n131, u1_u13_u6_n132, u1_u13_u6_n133, 
       u1_u13_u6_n134, u1_u13_u6_n135, u1_u13_u6_n136, u1_u13_u6_n137, u1_u13_u6_n138, u1_u13_u6_n139, u1_u13_u6_n140, u1_u13_u6_n141, u1_u13_u6_n142, 
       u1_u13_u6_n143, u1_u13_u6_n144, u1_u13_u6_n145, u1_u13_u6_n146, u1_u13_u6_n147, u1_u13_u6_n148, u1_u13_u6_n149, u1_u13_u6_n150, u1_u13_u6_n151, 
       u1_u13_u6_n152, u1_u13_u6_n153, u1_u13_u6_n154, u1_u13_u6_n155, u1_u13_u6_n156, u1_u13_u6_n157, u1_u13_u6_n158, u1_u13_u6_n159, u1_u13_u6_n160, 
       u1_u13_u6_n161, u1_u13_u6_n162, u1_u13_u6_n163, u1_u13_u6_n164, u1_u13_u6_n165, u1_u13_u6_n166, u1_u13_u6_n167, u1_u13_u6_n168, u1_u13_u6_n169, 
       u1_u13_u6_n170, u1_u13_u6_n171, u1_u13_u6_n172, u1_u13_u6_n173, u1_u13_u6_n174, u1_u13_u6_n88, u1_u13_u6_n89, u1_u13_u6_n90, u1_u13_u6_n91, 
       u1_u13_u6_n92, u1_u13_u6_n93, u1_u13_u6_n94, u1_u13_u6_n95, u1_u13_u6_n96, u1_u13_u6_n97, u1_u13_u6_n98, u1_u13_u6_n99, u1_u13_u7_n100, 
       u1_u13_u7_n101, u1_u13_u7_n102, u1_u13_u7_n103, u1_u13_u7_n104, u1_u13_u7_n105, u1_u13_u7_n106, u1_u13_u7_n107, u1_u13_u7_n108, u1_u13_u7_n109, 
       u1_u13_u7_n110, u1_u13_u7_n111, u1_u13_u7_n112, u1_u13_u7_n113, u1_u13_u7_n114, u1_u13_u7_n115, u1_u13_u7_n116, u1_u13_u7_n117, u1_u13_u7_n118, 
       u1_u13_u7_n119, u1_u13_u7_n120, u1_u13_u7_n121, u1_u13_u7_n122, u1_u13_u7_n123, u1_u13_u7_n124, u1_u13_u7_n125, u1_u13_u7_n126, u1_u13_u7_n127, 
       u1_u13_u7_n128, u1_u13_u7_n129, u1_u13_u7_n130, u1_u13_u7_n131, u1_u13_u7_n132, u1_u13_u7_n133, u1_u13_u7_n134, u1_u13_u7_n135, u1_u13_u7_n136, 
       u1_u13_u7_n137, u1_u13_u7_n138, u1_u13_u7_n139, u1_u13_u7_n140, u1_u13_u7_n141, u1_u13_u7_n142, u1_u13_u7_n143, u1_u13_u7_n144, u1_u13_u7_n145, 
       u1_u13_u7_n146, u1_u13_u7_n147, u1_u13_u7_n148, u1_u13_u7_n149, u1_u13_u7_n150, u1_u13_u7_n151, u1_u13_u7_n152, u1_u13_u7_n153, u1_u13_u7_n154, 
       u1_u13_u7_n155, u1_u13_u7_n156, u1_u13_u7_n157, u1_u13_u7_n158, u1_u13_u7_n159, u1_u13_u7_n160, u1_u13_u7_n161, u1_u13_u7_n162, u1_u13_u7_n163, 
       u1_u13_u7_n164, u1_u13_u7_n165, u1_u13_u7_n166, u1_u13_u7_n167, u1_u13_u7_n168, u1_u13_u7_n169, u1_u13_u7_n170, u1_u13_u7_n171, u1_u13_u7_n172, 
       u1_u13_u7_n173, u1_u13_u7_n174, u1_u13_u7_n175, u1_u13_u7_n176, u1_u13_u7_n177, u1_u13_u7_n178, u1_u13_u7_n179, u1_u13_u7_n180, u1_u13_u7_n91, 
       u1_u13_u7_n92, u1_u13_u7_n93, u1_u13_u7_n94, u1_u13_u7_n95, u1_u13_u7_n96, u1_u13_u7_n97, u1_u13_u7_n98, u1_u13_u7_n99, u1_u14_X_13, 
       u1_u14_X_14, u1_u14_X_15, u1_u14_X_16, u1_u14_X_17, u1_u14_X_18, u1_u14_X_31, u1_u14_X_32, u1_u14_X_33, u1_u14_X_34, 
       u1_u14_X_35, u1_u14_X_36, u1_u14_X_37, u1_u14_X_38, u1_u14_X_39, u1_u14_X_40, u1_u14_X_41, u1_u14_X_42, u1_u14_X_43, 
       u1_u14_X_44, u1_u14_X_45, u1_u14_X_46, u1_u14_X_47, u1_u14_X_48, u1_u14_u2_n100, u1_u14_u2_n101, u1_u14_u2_n102, u1_u14_u2_n103, 
       u1_u14_u2_n104, u1_u14_u2_n105, u1_u14_u2_n106, u1_u14_u2_n107, u1_u14_u2_n108, u1_u14_u2_n109, u1_u14_u2_n110, u1_u14_u2_n111, u1_u14_u2_n112, 
       u1_u14_u2_n113, u1_u14_u2_n114, u1_u14_u2_n115, u1_u14_u2_n116, u1_u14_u2_n117, u1_u14_u2_n118, u1_u14_u2_n119, u1_u14_u2_n120, u1_u14_u2_n121, 
       u1_u14_u2_n122, u1_u14_u2_n123, u1_u14_u2_n124, u1_u14_u2_n125, u1_u14_u2_n126, u1_u14_u2_n127, u1_u14_u2_n128, u1_u14_u2_n129, u1_u14_u2_n130, 
       u1_u14_u2_n131, u1_u14_u2_n132, u1_u14_u2_n133, u1_u14_u2_n134, u1_u14_u2_n135, u1_u14_u2_n136, u1_u14_u2_n137, u1_u14_u2_n138, u1_u14_u2_n139, 
       u1_u14_u2_n140, u1_u14_u2_n141, u1_u14_u2_n142, u1_u14_u2_n143, u1_u14_u2_n144, u1_u14_u2_n145, u1_u14_u2_n146, u1_u14_u2_n147, u1_u14_u2_n148, 
       u1_u14_u2_n149, u1_u14_u2_n150, u1_u14_u2_n151, u1_u14_u2_n152, u1_u14_u2_n153, u1_u14_u2_n154, u1_u14_u2_n155, u1_u14_u2_n156, u1_u14_u2_n157, 
       u1_u14_u2_n158, u1_u14_u2_n159, u1_u14_u2_n160, u1_u14_u2_n161, u1_u14_u2_n162, u1_u14_u2_n163, u1_u14_u2_n164, u1_u14_u2_n165, u1_u14_u2_n166, 
       u1_u14_u2_n167, u1_u14_u2_n168, u1_u14_u2_n169, u1_u14_u2_n170, u1_u14_u2_n171, u1_u14_u2_n172, u1_u14_u2_n173, u1_u14_u2_n174, u1_u14_u2_n175, 
       u1_u14_u2_n176, u1_u14_u2_n177, u1_u14_u2_n178, u1_u14_u2_n179, u1_u14_u2_n180, u1_u14_u2_n181, u1_u14_u2_n182, u1_u14_u2_n183, u1_u14_u2_n184, 
       u1_u14_u2_n185, u1_u14_u2_n186, u1_u14_u2_n187, u1_u14_u2_n188, u1_u14_u2_n95, u1_u14_u2_n96, u1_u14_u2_n97, u1_u14_u2_n98, u1_u14_u2_n99, 
       u1_u14_u5_n100, u1_u14_u5_n101, u1_u14_u5_n102, u1_u14_u5_n103, u1_u14_u5_n104, u1_u14_u5_n105, u1_u14_u5_n106, u1_u14_u5_n107, u1_u14_u5_n108, 
       u1_u14_u5_n109, u1_u14_u5_n110, u1_u14_u5_n111, u1_u14_u5_n112, u1_u14_u5_n113, u1_u14_u5_n114, u1_u14_u5_n115, u1_u14_u5_n116, u1_u14_u5_n117, 
       u1_u14_u5_n118, u1_u14_u5_n119, u1_u14_u5_n120, u1_u14_u5_n121, u1_u14_u5_n122, u1_u14_u5_n123, u1_u14_u5_n124, u1_u14_u5_n125, u1_u14_u5_n126, 
       u1_u14_u5_n127, u1_u14_u5_n128, u1_u14_u5_n129, u1_u14_u5_n130, u1_u14_u5_n131, u1_u14_u5_n132, u1_u14_u5_n133, u1_u14_u5_n134, u1_u14_u5_n135, 
       u1_u14_u5_n136, u1_u14_u5_n137, u1_u14_u5_n138, u1_u14_u5_n139, u1_u14_u5_n140, u1_u14_u5_n141, u1_u14_u5_n142, u1_u14_u5_n143, u1_u14_u5_n144, 
       u1_u14_u5_n145, u1_u14_u5_n146, u1_u14_u5_n147, u1_u14_u5_n148, u1_u14_u5_n149, u1_u14_u5_n150, u1_u14_u5_n151, u1_u14_u5_n152, u1_u14_u5_n153, 
       u1_u14_u5_n154, u1_u14_u5_n155, u1_u14_u5_n156, u1_u14_u5_n157, u1_u14_u5_n158, u1_u14_u5_n159, u1_u14_u5_n160, u1_u14_u5_n161, u1_u14_u5_n162, 
       u1_u14_u5_n163, u1_u14_u5_n164, u1_u14_u5_n165, u1_u14_u5_n166, u1_u14_u5_n167, u1_u14_u5_n168, u1_u14_u5_n169, u1_u14_u5_n170, u1_u14_u5_n171, 
       u1_u14_u5_n172, u1_u14_u5_n173, u1_u14_u5_n174, u1_u14_u5_n175, u1_u14_u5_n176, u1_u14_u5_n177, u1_u14_u5_n178, u1_u14_u5_n179, u1_u14_u5_n180, 
       u1_u14_u5_n181, u1_u14_u5_n182, u1_u14_u5_n183, u1_u14_u5_n184, u1_u14_u5_n185, u1_u14_u5_n186, u1_u14_u5_n187, u1_u14_u5_n188, u1_u14_u5_n189, 
       u1_u14_u5_n190, u1_u14_u5_n191, u1_u14_u5_n192, u1_u14_u5_n193, u1_u14_u5_n194, u1_u14_u5_n195, u1_u14_u5_n196, u1_u14_u5_n99, u1_u14_u6_n100, 
       u1_u14_u6_n101, u1_u14_u6_n102, u1_u14_u6_n103, u1_u14_u6_n104, u1_u14_u6_n105, u1_u14_u6_n106, u1_u14_u6_n107, u1_u14_u6_n108, u1_u14_u6_n109, 
       u1_u14_u6_n110, u1_u14_u6_n111, u1_u14_u6_n112, u1_u14_u6_n113, u1_u14_u6_n114, u1_u14_u6_n115, u1_u14_u6_n116, u1_u14_u6_n117, u1_u14_u6_n118, 
       u1_u14_u6_n119, u1_u14_u6_n120, u1_u14_u6_n121, u1_u14_u6_n122, u1_u14_u6_n123, u1_u14_u6_n124, u1_u14_u6_n125, u1_u14_u6_n126, u1_u14_u6_n127, 
       u1_u14_u6_n128, u1_u14_u6_n129, u1_u14_u6_n130, u1_u14_u6_n131, u1_u14_u6_n132, u1_u14_u6_n133, u1_u14_u6_n134, u1_u14_u6_n135, u1_u14_u6_n136, 
       u1_u14_u6_n137, u1_u14_u6_n138, u1_u14_u6_n139, u1_u14_u6_n140, u1_u14_u6_n141, u1_u14_u6_n142, u1_u14_u6_n143, u1_u14_u6_n144, u1_u14_u6_n145, 
       u1_u14_u6_n146, u1_u14_u6_n147, u1_u14_u6_n148, u1_u14_u6_n149, u1_u14_u6_n150, u1_u14_u6_n151, u1_u14_u6_n152, u1_u14_u6_n153, u1_u14_u6_n154, 
       u1_u14_u6_n155, u1_u14_u6_n156, u1_u14_u6_n157, u1_u14_u6_n158, u1_u14_u6_n159, u1_u14_u6_n160, u1_u14_u6_n161, u1_u14_u6_n162, u1_u14_u6_n163, 
       u1_u14_u6_n164, u1_u14_u6_n165, u1_u14_u6_n166, u1_u14_u6_n167, u1_u14_u6_n168, u1_u14_u6_n169, u1_u14_u6_n170, u1_u14_u6_n171, u1_u14_u6_n172, 
       u1_u14_u6_n173, u1_u14_u6_n174, u1_u14_u6_n88, u1_u14_u6_n89, u1_u14_u6_n90, u1_u14_u6_n91, u1_u14_u6_n92, u1_u14_u6_n93, u1_u14_u6_n94, 
       u1_u14_u6_n95, u1_u14_u6_n96, u1_u14_u6_n97, u1_u14_u6_n98, u1_u14_u6_n99, u1_u14_u7_n100, u1_u14_u7_n101, u1_u14_u7_n102, u1_u14_u7_n103, 
       u1_u14_u7_n104, u1_u14_u7_n105, u1_u14_u7_n106, u1_u14_u7_n107, u1_u14_u7_n108, u1_u14_u7_n109, u1_u14_u7_n110, u1_u14_u7_n111, u1_u14_u7_n112, 
       u1_u14_u7_n113, u1_u14_u7_n114, u1_u14_u7_n115, u1_u14_u7_n116, u1_u14_u7_n117, u1_u14_u7_n118, u1_u14_u7_n119, u1_u14_u7_n120, u1_u14_u7_n121, 
       u1_u14_u7_n122, u1_u14_u7_n123, u1_u14_u7_n124, u1_u14_u7_n125, u1_u14_u7_n126, u1_u14_u7_n127, u1_u14_u7_n128, u1_u14_u7_n129, u1_u14_u7_n130, 
       u1_u14_u7_n131, u1_u14_u7_n132, u1_u14_u7_n133, u1_u14_u7_n134, u1_u14_u7_n135, u1_u14_u7_n136, u1_u14_u7_n137, u1_u14_u7_n138, u1_u14_u7_n139, 
       u1_u14_u7_n140, u1_u14_u7_n141, u1_u14_u7_n142, u1_u14_u7_n143, u1_u14_u7_n144, u1_u14_u7_n145, u1_u14_u7_n146, u1_u14_u7_n147, u1_u14_u7_n148, 
       u1_u14_u7_n149, u1_u14_u7_n150, u1_u14_u7_n151, u1_u14_u7_n152, u1_u14_u7_n153, u1_u14_u7_n154, u1_u14_u7_n155, u1_u14_u7_n156, u1_u14_u7_n157, 
       u1_u14_u7_n158, u1_u14_u7_n159, u1_u14_u7_n160, u1_u14_u7_n161, u1_u14_u7_n162, u1_u14_u7_n163, u1_u14_u7_n164, u1_u14_u7_n165, u1_u14_u7_n166, 
       u1_u14_u7_n167, u1_u14_u7_n168, u1_u14_u7_n169, u1_u14_u7_n170, u1_u14_u7_n171, u1_u14_u7_n172, u1_u14_u7_n173, u1_u14_u7_n174, u1_u14_u7_n175, 
       u1_u14_u7_n176, u1_u14_u7_n177, u1_u14_u7_n178, u1_u14_u7_n179, u1_u14_u7_n180, u1_u14_u7_n91, u1_u14_u7_n92, u1_u14_u7_n93, u1_u14_u7_n94, 
       u1_u14_u7_n95, u1_u14_u7_n96, u1_u14_u7_n97, u1_u14_u7_n98, u1_u14_u7_n99, u1_u15_X_19, u1_u15_X_20, u1_u15_X_21, u1_u15_X_22, 
       u1_u15_X_23, u1_u15_X_24, u1_u15_X_25, u1_u15_X_26, u1_u15_X_27, u1_u15_X_28, u1_u15_X_29, u1_u15_X_30, u1_u15_u3_n100, 
       u1_u15_u3_n101, u1_u15_u3_n102, u1_u15_u3_n103, u1_u15_u3_n104, u1_u15_u3_n105, u1_u15_u3_n106, u1_u15_u3_n107, u1_u15_u3_n108, u1_u15_u3_n109, 
       u1_u15_u3_n110, u1_u15_u3_n111, u1_u15_u3_n112, u1_u15_u3_n113, u1_u15_u3_n114, u1_u15_u3_n115, u1_u15_u3_n116, u1_u15_u3_n117, u1_u15_u3_n118, 
       u1_u15_u3_n119, u1_u15_u3_n120, u1_u15_u3_n121, u1_u15_u3_n122, u1_u15_u3_n123, u1_u15_u3_n124, u1_u15_u3_n125, u1_u15_u3_n126, u1_u15_u3_n127, 
       u1_u15_u3_n128, u1_u15_u3_n129, u1_u15_u3_n130, u1_u15_u3_n131, u1_u15_u3_n132, u1_u15_u3_n133, u1_u15_u3_n134, u1_u15_u3_n135, u1_u15_u3_n136, 
       u1_u15_u3_n137, u1_u15_u3_n138, u1_u15_u3_n139, u1_u15_u3_n140, u1_u15_u3_n141, u1_u15_u3_n142, u1_u15_u3_n143, u1_u15_u3_n144, u1_u15_u3_n145, 
       u1_u15_u3_n146, u1_u15_u3_n147, u1_u15_u3_n148, u1_u15_u3_n149, u1_u15_u3_n150, u1_u15_u3_n151, u1_u15_u3_n152, u1_u15_u3_n153, u1_u15_u3_n154, 
       u1_u15_u3_n155, u1_u15_u3_n156, u1_u15_u3_n157, u1_u15_u3_n158, u1_u15_u3_n159, u1_u15_u3_n160, u1_u15_u3_n161, u1_u15_u3_n162, u1_u15_u3_n163, 
       u1_u15_u3_n164, u1_u15_u3_n165, u1_u15_u3_n166, u1_u15_u3_n167, u1_u15_u3_n168, u1_u15_u3_n169, u1_u15_u3_n170, u1_u15_u3_n171, u1_u15_u3_n172, 
       u1_u15_u3_n173, u1_u15_u3_n174, u1_u15_u3_n175, u1_u15_u3_n176, u1_u15_u3_n177, u1_u15_u3_n178, u1_u15_u3_n179, u1_u15_u3_n180, u1_u15_u3_n181, 
       u1_u15_u3_n182, u1_u15_u3_n183, u1_u15_u3_n184, u1_u15_u3_n185, u1_u15_u3_n186, u1_u15_u3_n94, u1_u15_u3_n95, u1_u15_u3_n96, u1_u15_u3_n97, 
       u1_u15_u3_n98, u1_u15_u3_n99, u1_u15_u4_n100, u1_u15_u4_n101, u1_u15_u4_n102, u1_u15_u4_n103, u1_u15_u4_n104, u1_u15_u4_n105, u1_u15_u4_n106, 
       u1_u15_u4_n107, u1_u15_u4_n108, u1_u15_u4_n109, u1_u15_u4_n110, u1_u15_u4_n111, u1_u15_u4_n112, u1_u15_u4_n113, u1_u15_u4_n114, u1_u15_u4_n115, 
       u1_u15_u4_n116, u1_u15_u4_n117, u1_u15_u4_n118, u1_u15_u4_n119, u1_u15_u4_n120, u1_u15_u4_n121, u1_u15_u4_n122, u1_u15_u4_n123, u1_u15_u4_n124, 
       u1_u15_u4_n125, u1_u15_u4_n126, u1_u15_u4_n127, u1_u15_u4_n128, u1_u15_u4_n129, u1_u15_u4_n130, u1_u15_u4_n131, u1_u15_u4_n132, u1_u15_u4_n133, 
       u1_u15_u4_n134, u1_u15_u4_n135, u1_u15_u4_n136, u1_u15_u4_n137, u1_u15_u4_n138, u1_u15_u4_n139, u1_u15_u4_n140, u1_u15_u4_n141, u1_u15_u4_n142, 
       u1_u15_u4_n143, u1_u15_u4_n144, u1_u15_u4_n145, u1_u15_u4_n146, u1_u15_u4_n147, u1_u15_u4_n148, u1_u15_u4_n149, u1_u15_u4_n150, u1_u15_u4_n151, 
       u1_u15_u4_n152, u1_u15_u4_n153, u1_u15_u4_n154, u1_u15_u4_n155, u1_u15_u4_n156, u1_u15_u4_n157, u1_u15_u4_n158, u1_u15_u4_n159, u1_u15_u4_n160, 
       u1_u15_u4_n161, u1_u15_u4_n162, u1_u15_u4_n163, u1_u15_u4_n164, u1_u15_u4_n165, u1_u15_u4_n166, u1_u15_u4_n167, u1_u15_u4_n168, u1_u15_u4_n169, 
       u1_u15_u4_n170, u1_u15_u4_n171, u1_u15_u4_n172, u1_u15_u4_n173, u1_u15_u4_n174, u1_u15_u4_n175, u1_u15_u4_n176, u1_u15_u4_n177, u1_u15_u4_n178, 
       u1_u15_u4_n179, u1_u15_u4_n180, u1_u15_u4_n181, u1_u15_u4_n182, u1_u15_u4_n183, u1_u15_u4_n184, u1_u15_u4_n185, u1_u15_u4_n186, u1_u15_u4_n94, 
       u1_u15_u4_n95, u1_u15_u4_n96, u1_u15_u4_n97, u1_u15_u4_n98, u1_u15_u4_n99, u1_u1_X_1, u1_u1_X_13, u1_u1_X_14, u1_u1_X_15, 
       u1_u1_X_16, u1_u1_X_17, u1_u1_X_18, u1_u1_X_19, u1_u1_X_2, u1_u1_X_20, u1_u1_X_21, u1_u1_X_22, u1_u1_X_23, 
       u1_u1_X_24, u1_u1_X_25, u1_u1_X_26, u1_u1_X_27, u1_u1_X_28, u1_u1_X_29, u1_u1_X_3, u1_u1_X_30, u1_u1_X_37, 
       u1_u1_X_38, u1_u1_X_39, u1_u1_X_4, u1_u1_X_40, u1_u1_X_41, u1_u1_X_42, u1_u1_X_43, u1_u1_X_44, u1_u1_X_45, 
       u1_u1_X_46, u1_u1_X_47, u1_u1_X_48, u1_u1_X_5, u1_u1_X_6, u1_u1_u0_n100, u1_u1_u0_n101, u1_u1_u0_n102, u1_u1_u0_n103, 
       u1_u1_u0_n104, u1_u1_u0_n105, u1_u1_u0_n106, u1_u1_u0_n107, u1_u1_u0_n108, u1_u1_u0_n109, u1_u1_u0_n110, u1_u1_u0_n111, u1_u1_u0_n112, 
       u1_u1_u0_n113, u1_u1_u0_n114, u1_u1_u0_n115, u1_u1_u0_n116, u1_u1_u0_n117, u1_u1_u0_n118, u1_u1_u0_n119, u1_u1_u0_n120, u1_u1_u0_n121, 
       u1_u1_u0_n122, u1_u1_u0_n123, u1_u1_u0_n124, u1_u1_u0_n125, u1_u1_u0_n126, u1_u1_u0_n127, u1_u1_u0_n128, u1_u1_u0_n129, u1_u1_u0_n130, 
       u1_u1_u0_n131, u1_u1_u0_n132, u1_u1_u0_n133, u1_u1_u0_n134, u1_u1_u0_n135, u1_u1_u0_n136, u1_u1_u0_n137, u1_u1_u0_n138, u1_u1_u0_n139, 
       u1_u1_u0_n140, u1_u1_u0_n141, u1_u1_u0_n142, u1_u1_u0_n143, u1_u1_u0_n144, u1_u1_u0_n145, u1_u1_u0_n146, u1_u1_u0_n147, u1_u1_u0_n148, 
       u1_u1_u0_n149, u1_u1_u0_n150, u1_u1_u0_n151, u1_u1_u0_n152, u1_u1_u0_n153, u1_u1_u0_n154, u1_u1_u0_n155, u1_u1_u0_n156, u1_u1_u0_n157, 
       u1_u1_u0_n158, u1_u1_u0_n159, u1_u1_u0_n160, u1_u1_u0_n161, u1_u1_u0_n162, u1_u1_u0_n163, u1_u1_u0_n164, u1_u1_u0_n165, u1_u1_u0_n166, 
       u1_u1_u0_n167, u1_u1_u0_n168, u1_u1_u0_n169, u1_u1_u0_n170, u1_u1_u0_n171, u1_u1_u0_n172, u1_u1_u0_n173, u1_u1_u0_n174, u1_u1_u0_n88, 
       u1_u1_u0_n89, u1_u1_u0_n90, u1_u1_u0_n91, u1_u1_u0_n92, u1_u1_u0_n93, u1_u1_u0_n94, u1_u1_u0_n95, u1_u1_u0_n96, u1_u1_u0_n97, 
       u1_u1_u0_n98, u1_u1_u0_n99, u1_u1_u2_n100, u1_u1_u2_n101, u1_u1_u2_n102, u1_u1_u2_n103, u1_u1_u2_n104, u1_u1_u2_n105, u1_u1_u2_n106, 
       u1_u1_u2_n107, u1_u1_u2_n108, u1_u1_u2_n109, u1_u1_u2_n110, u1_u1_u2_n111, u1_u1_u2_n112, u1_u1_u2_n113, u1_u1_u2_n114, u1_u1_u2_n115, 
       u1_u1_u2_n116, u1_u1_u2_n117, u1_u1_u2_n118, u1_u1_u2_n119, u1_u1_u2_n120, u1_u1_u2_n121, u1_u1_u2_n122, u1_u1_u2_n123, u1_u1_u2_n124, 
       u1_u1_u2_n125, u1_u1_u2_n126, u1_u1_u2_n127, u1_u1_u2_n128, u1_u1_u2_n129, u1_u1_u2_n130, u1_u1_u2_n131, u1_u1_u2_n132, u1_u1_u2_n133, 
       u1_u1_u2_n134, u1_u1_u2_n135, u1_u1_u2_n136, u1_u1_u2_n137, u1_u1_u2_n138, u1_u1_u2_n139, u1_u1_u2_n140, u1_u1_u2_n141, u1_u1_u2_n142, 
       u1_u1_u2_n143, u1_u1_u2_n144, u1_u1_u2_n145, u1_u1_u2_n146, u1_u1_u2_n147, u1_u1_u2_n148, u1_u1_u2_n149, u1_u1_u2_n150, u1_u1_u2_n151, 
       u1_u1_u2_n152, u1_u1_u2_n153, u1_u1_u2_n154, u1_u1_u2_n155, u1_u1_u2_n156, u1_u1_u2_n157, u1_u1_u2_n158, u1_u1_u2_n159, u1_u1_u2_n160, 
       u1_u1_u2_n161, u1_u1_u2_n162, u1_u1_u2_n163, u1_u1_u2_n164, u1_u1_u2_n165, u1_u1_u2_n166, u1_u1_u2_n167, u1_u1_u2_n168, u1_u1_u2_n169, 
       u1_u1_u2_n170, u1_u1_u2_n171, u1_u1_u2_n172, u1_u1_u2_n173, u1_u1_u2_n174, u1_u1_u2_n175, u1_u1_u2_n176, u1_u1_u2_n177, u1_u1_u2_n178, 
       u1_u1_u2_n179, u1_u1_u2_n180, u1_u1_u2_n181, u1_u1_u2_n182, u1_u1_u2_n183, u1_u1_u2_n184, u1_u1_u2_n185, u1_u1_u2_n186, u1_u1_u2_n187, 
       u1_u1_u2_n188, u1_u1_u2_n95, u1_u1_u2_n96, u1_u1_u2_n97, u1_u1_u2_n98, u1_u1_u2_n99, u1_u1_u3_n100, u1_u1_u3_n101, u1_u1_u3_n102, 
       u1_u1_u3_n103, u1_u1_u3_n104, u1_u1_u3_n105, u1_u1_u3_n106, u1_u1_u3_n107, u1_u1_u3_n108, u1_u1_u3_n109, u1_u1_u3_n110, u1_u1_u3_n111, 
       u1_u1_u3_n112, u1_u1_u3_n113, u1_u1_u3_n114, u1_u1_u3_n115, u1_u1_u3_n116, u1_u1_u3_n117, u1_u1_u3_n118, u1_u1_u3_n119, u1_u1_u3_n120, 
       u1_u1_u3_n121, u1_u1_u3_n122, u1_u1_u3_n123, u1_u1_u3_n124, u1_u1_u3_n125, u1_u1_u3_n126, u1_u1_u3_n127, u1_u1_u3_n128, u1_u1_u3_n129, 
       u1_u1_u3_n130, u1_u1_u3_n131, u1_u1_u3_n132, u1_u1_u3_n133, u1_u1_u3_n134, u1_u1_u3_n135, u1_u1_u3_n136, u1_u1_u3_n137, u1_u1_u3_n138, 
       u1_u1_u3_n139, u1_u1_u3_n140, u1_u1_u3_n141, u1_u1_u3_n142, u1_u1_u3_n143, u1_u1_u3_n144, u1_u1_u3_n145, u1_u1_u3_n146, u1_u1_u3_n147, 
       u1_u1_u3_n148, u1_u1_u3_n149, u1_u1_u3_n150, u1_u1_u3_n151, u1_u1_u3_n152, u1_u1_u3_n153, u1_u1_u3_n154, u1_u1_u3_n155, u1_u1_u3_n156, 
       u1_u1_u3_n157, u1_u1_u3_n158, u1_u1_u3_n159, u1_u1_u3_n160, u1_u1_u3_n161, u1_u1_u3_n162, u1_u1_u3_n163, u1_u1_u3_n164, u1_u1_u3_n165, 
       u1_u1_u3_n166, u1_u1_u3_n167, u1_u1_u3_n168, u1_u1_u3_n169, u1_u1_u3_n170, u1_u1_u3_n171, u1_u1_u3_n172, u1_u1_u3_n173, u1_u1_u3_n174, 
       u1_u1_u3_n175, u1_u1_u3_n176, u1_u1_u3_n177, u1_u1_u3_n178, u1_u1_u3_n179, u1_u1_u3_n180, u1_u1_u3_n181, u1_u1_u3_n182, u1_u1_u3_n183, 
       u1_u1_u3_n184, u1_u1_u3_n185, u1_u1_u3_n186, u1_u1_u3_n94, u1_u1_u3_n95, u1_u1_u3_n96, u1_u1_u3_n97, u1_u1_u3_n98, u1_u1_u3_n99, 
       u1_u1_u4_n100, u1_u1_u4_n101, u1_u1_u4_n102, u1_u1_u4_n103, u1_u1_u4_n104, u1_u1_u4_n105, u1_u1_u4_n106, u1_u1_u4_n107, u1_u1_u4_n108, 
       u1_u1_u4_n109, u1_u1_u4_n110, u1_u1_u4_n111, u1_u1_u4_n112, u1_u1_u4_n113, u1_u1_u4_n114, u1_u1_u4_n115, u1_u1_u4_n116, u1_u1_u4_n117, 
       u1_u1_u4_n118, u1_u1_u4_n119, u1_u1_u4_n120, u1_u1_u4_n121, u1_u1_u4_n122, u1_u1_u4_n123, u1_u1_u4_n124, u1_u1_u4_n125, u1_u1_u4_n126, 
       u1_u1_u4_n127, u1_u1_u4_n128, u1_u1_u4_n129, u1_u1_u4_n130, u1_u1_u4_n131, u1_u1_u4_n132, u1_u1_u4_n133, u1_u1_u4_n134, u1_u1_u4_n135, 
       u1_u1_u4_n136, u1_u1_u4_n137, u1_u1_u4_n138, u1_u1_u4_n139, u1_u1_u4_n140, u1_u1_u4_n141, u1_u1_u4_n142, u1_u1_u4_n143, u1_u1_u4_n144, 
       u1_u1_u4_n145, u1_u1_u4_n146, u1_u1_u4_n147, u1_u1_u4_n148, u1_u1_u4_n149, u1_u1_u4_n150, u1_u1_u4_n151, u1_u1_u4_n152, u1_u1_u4_n153, 
       u1_u1_u4_n154, u1_u1_u4_n155, u1_u1_u4_n156, u1_u1_u4_n157, u1_u1_u4_n158, u1_u1_u4_n159, u1_u1_u4_n160, u1_u1_u4_n161, u1_u1_u4_n162, 
       u1_u1_u4_n163, u1_u1_u4_n164, u1_u1_u4_n165, u1_u1_u4_n166, u1_u1_u4_n167, u1_u1_u4_n168, u1_u1_u4_n169, u1_u1_u4_n170, u1_u1_u4_n171, 
       u1_u1_u4_n172, u1_u1_u4_n173, u1_u1_u4_n174, u1_u1_u4_n175, u1_u1_u4_n176, u1_u1_u4_n177, u1_u1_u4_n178, u1_u1_u4_n179, u1_u1_u4_n180, 
       u1_u1_u4_n181, u1_u1_u4_n182, u1_u1_u4_n183, u1_u1_u4_n184, u1_u1_u4_n185, u1_u1_u4_n186, u1_u1_u4_n94, u1_u1_u4_n95, u1_u1_u4_n96, 
       u1_u1_u4_n97, u1_u1_u4_n98, u1_u1_u4_n99, u1_u1_u6_n100, u1_u1_u6_n101, u1_u1_u6_n102, u1_u1_u6_n103, u1_u1_u6_n104, u1_u1_u6_n105, 
       u1_u1_u6_n106, u1_u1_u6_n107, u1_u1_u6_n108, u1_u1_u6_n109, u1_u1_u6_n110, u1_u1_u6_n111, u1_u1_u6_n112, u1_u1_u6_n113, u1_u1_u6_n114, 
       u1_u1_u6_n115, u1_u1_u6_n116, u1_u1_u6_n117, u1_u1_u6_n118, u1_u1_u6_n119, u1_u1_u6_n120, u1_u1_u6_n121, u1_u1_u6_n122, u1_u1_u6_n123, 
       u1_u1_u6_n124, u1_u1_u6_n125, u1_u1_u6_n126, u1_u1_u6_n127, u1_u1_u6_n128, u1_u1_u6_n129, u1_u1_u6_n130, u1_u1_u6_n131, u1_u1_u6_n132, 
       u1_u1_u6_n133, u1_u1_u6_n134, u1_u1_u6_n135, u1_u1_u6_n136, u1_u1_u6_n137, u1_u1_u6_n138, u1_u1_u6_n139, u1_u1_u6_n140, u1_u1_u6_n141, 
       u1_u1_u6_n142, u1_u1_u6_n143, u1_u1_u6_n144, u1_u1_u6_n145, u1_u1_u6_n146, u1_u1_u6_n147, u1_u1_u6_n148, u1_u1_u6_n149, u1_u1_u6_n150, 
       u1_u1_u6_n151, u1_u1_u6_n152, u1_u1_u6_n153, u1_u1_u6_n154, u1_u1_u6_n155, u1_u1_u6_n156, u1_u1_u6_n157, u1_u1_u6_n158, u1_u1_u6_n159, 
       u1_u1_u6_n160, u1_u1_u6_n161, u1_u1_u6_n162, u1_u1_u6_n163, u1_u1_u6_n164, u1_u1_u6_n165, u1_u1_u6_n166, u1_u1_u6_n167, u1_u1_u6_n168, 
       u1_u1_u6_n169, u1_u1_u6_n170, u1_u1_u6_n171, u1_u1_u6_n172, u1_u1_u6_n173, u1_u1_u6_n174, u1_u1_u6_n88, u1_u1_u6_n89, u1_u1_u6_n90, 
       u1_u1_u6_n91, u1_u1_u6_n92, u1_u1_u6_n93, u1_u1_u6_n94, u1_u1_u6_n95, u1_u1_u6_n96, u1_u1_u6_n97, u1_u1_u6_n98, u1_u1_u6_n99, 
       u1_u1_u7_n100, u1_u1_u7_n101, u1_u1_u7_n102, u1_u1_u7_n103, u1_u1_u7_n104, u1_u1_u7_n105, u1_u1_u7_n106, u1_u1_u7_n107, u1_u1_u7_n108, 
       u1_u1_u7_n109, u1_u1_u7_n110, u1_u1_u7_n111, u1_u1_u7_n112, u1_u1_u7_n113, u1_u1_u7_n114, u1_u1_u7_n115, u1_u1_u7_n116, u1_u1_u7_n117, 
       u1_u1_u7_n118, u1_u1_u7_n119, u1_u1_u7_n120, u1_u1_u7_n121, u1_u1_u7_n122, u1_u1_u7_n123, u1_u1_u7_n124, u1_u1_u7_n125, u1_u1_u7_n126, 
       u1_u1_u7_n127, u1_u1_u7_n128, u1_u1_u7_n129, u1_u1_u7_n130, u1_u1_u7_n131, u1_u1_u7_n132, u1_u1_u7_n133, u1_u1_u7_n134, u1_u1_u7_n135, 
       u1_u1_u7_n136, u1_u1_u7_n137, u1_u1_u7_n138, u1_u1_u7_n139, u1_u1_u7_n140, u1_u1_u7_n141, u1_u1_u7_n142, u1_u1_u7_n143, u1_u1_u7_n144, 
       u1_u1_u7_n145, u1_u1_u7_n146, u1_u1_u7_n147, u1_u1_u7_n148, u1_u1_u7_n149, u1_u1_u7_n150, u1_u1_u7_n151, u1_u1_u7_n152, u1_u1_u7_n153, 
       u1_u1_u7_n154, u1_u1_u7_n155, u1_u1_u7_n156, u1_u1_u7_n157, u1_u1_u7_n158, u1_u1_u7_n159, u1_u1_u7_n160, u1_u1_u7_n161, u1_u1_u7_n162, 
       u1_u1_u7_n163, u1_u1_u7_n164, u1_u1_u7_n165, u1_u1_u7_n166, u1_u1_u7_n167, u1_u1_u7_n168, u1_u1_u7_n169, u1_u1_u7_n170, u1_u1_u7_n171, 
       u1_u1_u7_n172, u1_u1_u7_n173, u1_u1_u7_n174, u1_u1_u7_n175, u1_u1_u7_n176, u1_u1_u7_n177, u1_u1_u7_n178, u1_u1_u7_n179, u1_u1_u7_n180, 
       u1_u1_u7_n91, u1_u1_u7_n92, u1_u1_u7_n93, u1_u1_u7_n94, u1_u1_u7_n95, u1_u1_u7_n96, u1_u1_u7_n97, u1_u1_u7_n98, u1_u1_u7_n99, 
       u1_u2_X_19, u1_u2_X_20, u1_u2_X_21, u1_u2_X_22, u1_u2_X_23, u1_u2_X_24, u1_u2_X_43, u1_u2_X_44, u1_u2_X_45, 
       u1_u2_X_46, u1_u2_X_47, u1_u2_X_48, u1_u2_u3_n100, u1_u2_u3_n101, u1_u2_u3_n102, u1_u2_u3_n103, u1_u2_u3_n104, u1_u2_u3_n105, 
       u1_u2_u3_n106, u1_u2_u3_n107, u1_u2_u3_n108, u1_u2_u3_n109, u1_u2_u3_n110, u1_u2_u3_n111, u1_u2_u3_n112, u1_u2_u3_n113, u1_u2_u3_n114, 
       u1_u2_u3_n115, u1_u2_u3_n116, u1_u2_u3_n117, u1_u2_u3_n118, u1_u2_u3_n119, u1_u2_u3_n120, u1_u2_u3_n121, u1_u2_u3_n122, u1_u2_u3_n123, 
       u1_u2_u3_n124, u1_u2_u3_n125, u1_u2_u3_n126, u1_u2_u3_n127, u1_u2_u3_n128, u1_u2_u3_n129, u1_u2_u3_n130, u1_u2_u3_n131, u1_u2_u3_n132, 
       u1_u2_u3_n133, u1_u2_u3_n134, u1_u2_u3_n135, u1_u2_u3_n136, u1_u2_u3_n137, u1_u2_u3_n138, u1_u2_u3_n139, u1_u2_u3_n140, u1_u2_u3_n141, 
       u1_u2_u3_n142, u1_u2_u3_n143, u1_u2_u3_n144, u1_u2_u3_n145, u1_u2_u3_n146, u1_u2_u3_n147, u1_u2_u3_n148, u1_u2_u3_n149, u1_u2_u3_n150, 
       u1_u2_u3_n151, u1_u2_u3_n152, u1_u2_u3_n153, u1_u2_u3_n154, u1_u2_u3_n155, u1_u2_u3_n156, u1_u2_u3_n157, u1_u2_u3_n158, u1_u2_u3_n159, 
       u1_u2_u3_n160, u1_u2_u3_n161, u1_u2_u3_n162, u1_u2_u3_n163, u1_u2_u3_n164, u1_u2_u3_n165, u1_u2_u3_n166, u1_u2_u3_n167, u1_u2_u3_n168, 
       u1_u2_u3_n169, u1_u2_u3_n170, u1_u2_u3_n171, u1_u2_u3_n172, u1_u2_u3_n173, u1_u2_u3_n174, u1_u2_u3_n175, u1_u2_u3_n176, u1_u2_u3_n177, 
       u1_u2_u3_n178, u1_u2_u3_n179, u1_u2_u3_n180, u1_u2_u3_n181, u1_u2_u3_n182, u1_u2_u3_n183, u1_u2_u3_n184, u1_u2_u3_n185, u1_u2_u3_n186, 
       u1_u2_u3_n94, u1_u2_u3_n95, u1_u2_u3_n96, u1_u2_u3_n97, u1_u2_u3_n98, u1_u2_u3_n99, u1_u2_u7_n100, u1_u2_u7_n101, u1_u2_u7_n102, 
       u1_u2_u7_n103, u1_u2_u7_n104, u1_u2_u7_n105, u1_u2_u7_n106, u1_u2_u7_n107, u1_u2_u7_n108, u1_u2_u7_n109, u1_u2_u7_n110, u1_u2_u7_n111, 
       u1_u2_u7_n112, u1_u2_u7_n113, u1_u2_u7_n114, u1_u2_u7_n115, u1_u2_u7_n116, u1_u2_u7_n117, u1_u2_u7_n118, u1_u2_u7_n119, u1_u2_u7_n120, 
       u1_u2_u7_n121, u1_u2_u7_n122, u1_u2_u7_n123, u1_u2_u7_n124, u1_u2_u7_n125, u1_u2_u7_n126, u1_u2_u7_n127, u1_u2_u7_n128, u1_u2_u7_n129, 
       u1_u2_u7_n130, u1_u2_u7_n131, u1_u2_u7_n132, u1_u2_u7_n133, u1_u2_u7_n134, u1_u2_u7_n135, u1_u2_u7_n136, u1_u2_u7_n137, u1_u2_u7_n138, 
       u1_u2_u7_n139, u1_u2_u7_n140, u1_u2_u7_n141, u1_u2_u7_n142, u1_u2_u7_n143, u1_u2_u7_n144, u1_u2_u7_n145, u1_u2_u7_n146, u1_u2_u7_n147, 
       u1_u2_u7_n148, u1_u2_u7_n149, u1_u2_u7_n150, u1_u2_u7_n151, u1_u2_u7_n152, u1_u2_u7_n153, u1_u2_u7_n154, u1_u2_u7_n155, u1_u2_u7_n156, 
       u1_u2_u7_n157, u1_u2_u7_n158, u1_u2_u7_n159, u1_u2_u7_n160, u1_u2_u7_n161, u1_u2_u7_n162, u1_u2_u7_n163, u1_u2_u7_n164, u1_u2_u7_n165, 
       u1_u2_u7_n166, u1_u2_u7_n167, u1_u2_u7_n168, u1_u2_u7_n169, u1_u2_u7_n170, u1_u2_u7_n171, u1_u2_u7_n172, u1_u2_u7_n173, u1_u2_u7_n174, 
       u1_u2_u7_n175, u1_u2_u7_n176, u1_u2_u7_n177, u1_u2_u7_n178, u1_u2_u7_n179, u1_u2_u7_n180, u1_u2_u7_n91, u1_u2_u7_n92, u1_u2_u7_n93, 
       u1_u2_u7_n94, u1_u2_u7_n95, u1_u2_u7_n96, u1_u2_u7_n97, u1_u2_u7_n98, u1_u2_u7_n99, u1_u3_X_19, u1_u3_X_20, u1_u3_X_21, 
       u1_u3_X_22, u1_u3_X_23, u1_u3_X_24, u1_u3_u3_n100, u1_u3_u3_n101, u1_u3_u3_n102, u1_u3_u3_n103, u1_u3_u3_n104, u1_u3_u3_n105, 
       u1_u3_u3_n106, u1_u3_u3_n107, u1_u3_u3_n108, u1_u3_u3_n109, u1_u3_u3_n110, u1_u3_u3_n111, u1_u3_u3_n112, u1_u3_u3_n113, u1_u3_u3_n114, 
       u1_u3_u3_n115, u1_u3_u3_n116, u1_u3_u3_n117, u1_u3_u3_n118, u1_u3_u3_n119, u1_u3_u3_n120, u1_u3_u3_n121, u1_u3_u3_n122, u1_u3_u3_n123, 
       u1_u3_u3_n124, u1_u3_u3_n125, u1_u3_u3_n126, u1_u3_u3_n127, u1_u3_u3_n128, u1_u3_u3_n129, u1_u3_u3_n130, u1_u3_u3_n131, u1_u3_u3_n132, 
       u1_u3_u3_n133, u1_u3_u3_n134, u1_u3_u3_n135, u1_u3_u3_n136, u1_u3_u3_n137, u1_u3_u3_n138, u1_u3_u3_n139, u1_u3_u3_n140, u1_u3_u3_n141, 
       u1_u3_u3_n142, u1_u3_u3_n143, u1_u3_u3_n144, u1_u3_u3_n145, u1_u3_u3_n146, u1_u3_u3_n147, u1_u3_u3_n148, u1_u3_u3_n149, u1_u3_u3_n150, 
       u1_u3_u3_n151, u1_u3_u3_n152, u1_u3_u3_n153, u1_u3_u3_n154, u1_u3_u3_n155, u1_u3_u3_n156, u1_u3_u3_n157, u1_u3_u3_n158, u1_u3_u3_n159, 
       u1_u3_u3_n160, u1_u3_u3_n161, u1_u3_u3_n162, u1_u3_u3_n163, u1_u3_u3_n164, u1_u3_u3_n165, u1_u3_u3_n166, u1_u3_u3_n167, u1_u3_u3_n168, 
       u1_u3_u3_n169, u1_u3_u3_n170, u1_u3_u3_n171, u1_u3_u3_n172, u1_u3_u3_n173, u1_u3_u3_n174, u1_u3_u3_n175, u1_u3_u3_n176, u1_u3_u3_n177, 
       u1_u3_u3_n178, u1_u3_u3_n179, u1_u3_u3_n180, u1_u3_u3_n181, u1_u3_u3_n182, u1_u3_u3_n183, u1_u3_u3_n184, u1_u3_u3_n185, u1_u3_u3_n186, 
       u1_u3_u3_n94, u1_u3_u3_n95, u1_u3_u3_n96, u1_u3_u3_n97, u1_u3_u3_n98, u1_u3_u3_n99, u1_u4_X_31, u1_u4_X_32, u1_u4_X_33, 
       u1_u4_X_34, u1_u4_X_35, u1_u4_X_36, u1_u4_X_43, u1_u4_X_44, u1_u4_X_45, u1_u4_X_46, u1_u4_X_47, u1_u4_X_48, 
       u1_u4_u5_n100, u1_u4_u5_n101, u1_u4_u5_n102, u1_u4_u5_n103, u1_u4_u5_n104, u1_u4_u5_n105, u1_u4_u5_n106, u1_u4_u5_n107, u1_u4_u5_n108, 
       u1_u4_u5_n109, u1_u4_u5_n110, u1_u4_u5_n111, u1_u4_u5_n112, u1_u4_u5_n113, u1_u4_u5_n114, u1_u4_u5_n115, u1_u4_u5_n116, u1_u4_u5_n117, 
       u1_u4_u5_n118, u1_u4_u5_n119, u1_u4_u5_n120, u1_u4_u5_n121, u1_u4_u5_n122, u1_u4_u5_n123, u1_u4_u5_n124, u1_u4_u5_n125, u1_u4_u5_n126, 
       u1_u4_u5_n127, u1_u4_u5_n128, u1_u4_u5_n129, u1_u4_u5_n130, u1_u4_u5_n131, u1_u4_u5_n132, u1_u4_u5_n133, u1_u4_u5_n134, u1_u4_u5_n135, 
       u1_u4_u5_n136, u1_u4_u5_n137, u1_u4_u5_n138, u1_u4_u5_n139, u1_u4_u5_n140, u1_u4_u5_n141, u1_u4_u5_n142, u1_u4_u5_n143, u1_u4_u5_n144, 
       u1_u4_u5_n145, u1_u4_u5_n146, u1_u4_u5_n147, u1_u4_u5_n148, u1_u4_u5_n149, u1_u4_u5_n150, u1_u4_u5_n151, u1_u4_u5_n152, u1_u4_u5_n153, 
       u1_u4_u5_n154, u1_u4_u5_n155, u1_u4_u5_n156, u1_u4_u5_n157, u1_u4_u5_n158, u1_u4_u5_n159, u1_u4_u5_n160, u1_u4_u5_n161, u1_u4_u5_n162, 
       u1_u4_u5_n163, u1_u4_u5_n164, u1_u4_u5_n165, u1_u4_u5_n166, u1_u4_u5_n167, u1_u4_u5_n168, u1_u4_u5_n169, u1_u4_u5_n170, u1_u4_u5_n171, 
       u1_u4_u5_n172, u1_u4_u5_n173, u1_u4_u5_n174, u1_u4_u5_n175, u1_u4_u5_n176, u1_u4_u5_n177, u1_u4_u5_n178, u1_u4_u5_n179, u1_u4_u5_n180, 
       u1_u4_u5_n181, u1_u4_u5_n182, u1_u4_u5_n183, u1_u4_u5_n184, u1_u4_u5_n185, u1_u4_u5_n186, u1_u4_u5_n187, u1_u4_u5_n188, u1_u4_u5_n189, 
       u1_u4_u5_n190, u1_u4_u5_n191, u1_u4_u5_n192, u1_u4_u5_n193, u1_u4_u5_n194, u1_u4_u5_n195, u1_u4_u5_n196, u1_u4_u5_n99, u1_u4_u7_n100, 
       u1_u4_u7_n101, u1_u4_u7_n102, u1_u4_u7_n103, u1_u4_u7_n104, u1_u4_u7_n105, u1_u4_u7_n106, u1_u4_u7_n107, u1_u4_u7_n108, u1_u4_u7_n109, 
       u1_u4_u7_n110, u1_u4_u7_n111, u1_u4_u7_n112, u1_u4_u7_n113, u1_u4_u7_n114, u1_u4_u7_n115, u1_u4_u7_n116, u1_u4_u7_n117, u1_u4_u7_n118, 
       u1_u4_u7_n119, u1_u4_u7_n120, u1_u4_u7_n121, u1_u4_u7_n122, u1_u4_u7_n123, u1_u4_u7_n124, u1_u4_u7_n125, u1_u4_u7_n126, u1_u4_u7_n127, 
       u1_u4_u7_n128, u1_u4_u7_n129, u1_u4_u7_n130, u1_u4_u7_n131, u1_u4_u7_n132, u1_u4_u7_n133, u1_u4_u7_n134, u1_u4_u7_n135, u1_u4_u7_n136, 
       u1_u4_u7_n137, u1_u4_u7_n138, u1_u4_u7_n139, u1_u4_u7_n140, u1_u4_u7_n141, u1_u4_u7_n142, u1_u4_u7_n143, u1_u4_u7_n144, u1_u4_u7_n145, 
       u1_u4_u7_n146, u1_u4_u7_n147, u1_u4_u7_n148, u1_u4_u7_n149, u1_u4_u7_n150, u1_u4_u7_n151, u1_u4_u7_n152, u1_u4_u7_n153, u1_u4_u7_n154, 
       u1_u4_u7_n155, u1_u4_u7_n156, u1_u4_u7_n157, u1_u4_u7_n158, u1_u4_u7_n159, u1_u4_u7_n160, u1_u4_u7_n161, u1_u4_u7_n162, u1_u4_u7_n163, 
       u1_u4_u7_n164, u1_u4_u7_n165, u1_u4_u7_n166, u1_u4_u7_n167, u1_u4_u7_n168, u1_u4_u7_n169, u1_u4_u7_n170, u1_u4_u7_n171, u1_u4_u7_n172, 
       u1_u4_u7_n173, u1_u4_u7_n174, u1_u4_u7_n175, u1_u4_u7_n176, u1_u4_u7_n177, u1_u4_u7_n178, u1_u4_u7_n179, u1_u4_u7_n180, u1_u4_u7_n91, 
       u1_u4_u7_n92, u1_u4_u7_n93, u1_u4_u7_n94, u1_u4_u7_n95, u1_u4_u7_n96, u1_u4_u7_n97, u1_u4_u7_n98, u1_u4_u7_n99, u1_u5_X_1, 
       u1_u5_X_13, u1_u5_X_14, u1_u5_X_15, u1_u5_X_16, u1_u5_X_17, u1_u5_X_18, u1_u5_X_19, u1_u5_X_2, u1_u5_X_20, 
       u1_u5_X_21, u1_u5_X_22, u1_u5_X_23, u1_u5_X_24, u1_u5_X_3, u1_u5_X_37, u1_u5_X_38, u1_u5_X_39, u1_u5_X_4, 
       u1_u5_X_40, u1_u5_X_41, u1_u5_X_42, u1_u5_X_5, u1_u5_X_6, u1_u5_u0_n100, u1_u5_u0_n101, u1_u5_u0_n102, u1_u5_u0_n103, 
       u1_u5_u0_n104, u1_u5_u0_n105, u1_u5_u0_n106, u1_u5_u0_n107, u1_u5_u0_n108, u1_u5_u0_n109, u1_u5_u0_n110, u1_u5_u0_n111, u1_u5_u0_n112, 
       u1_u5_u0_n113, u1_u5_u0_n114, u1_u5_u0_n115, u1_u5_u0_n116, u1_u5_u0_n117, u1_u5_u0_n118, u1_u5_u0_n119, u1_u5_u0_n120, u1_u5_u0_n121, 
       u1_u5_u0_n122, u1_u5_u0_n123, u1_u5_u0_n124, u1_u5_u0_n125, u1_u5_u0_n126, u1_u5_u0_n127, u1_u5_u0_n128, u1_u5_u0_n129, u1_u5_u0_n130, 
       u1_u5_u0_n131, u1_u5_u0_n132, u1_u5_u0_n133, u1_u5_u0_n134, u1_u5_u0_n135, u1_u5_u0_n136, u1_u5_u0_n137, u1_u5_u0_n138, u1_u5_u0_n139, 
       u1_u5_u0_n140, u1_u5_u0_n141, u1_u5_u0_n142, u1_u5_u0_n143, u1_u5_u0_n144, u1_u5_u0_n145, u1_u5_u0_n146, u1_u5_u0_n147, u1_u5_u0_n148, 
       u1_u5_u0_n149, u1_u5_u0_n150, u1_u5_u0_n151, u1_u5_u0_n152, u1_u5_u0_n153, u1_u5_u0_n154, u1_u5_u0_n155, u1_u5_u0_n156, u1_u5_u0_n157, 
       u1_u5_u0_n158, u1_u5_u0_n159, u1_u5_u0_n160, u1_u5_u0_n161, u1_u5_u0_n162, u1_u5_u0_n163, u1_u5_u0_n164, u1_u5_u0_n165, u1_u5_u0_n166, 
       u1_u5_u0_n167, u1_u5_u0_n168, u1_u5_u0_n169, u1_u5_u0_n170, u1_u5_u0_n171, u1_u5_u0_n172, u1_u5_u0_n173, u1_u5_u0_n174, u1_u5_u0_n88, 
       u1_u5_u0_n89, u1_u5_u0_n90, u1_u5_u0_n91, u1_u5_u0_n92, u1_u5_u0_n93, u1_u5_u0_n94, u1_u5_u0_n95, u1_u5_u0_n96, u1_u5_u0_n97, 
       u1_u5_u0_n98, u1_u5_u0_n99, u1_u5_u2_n100, u1_u5_u2_n101, u1_u5_u2_n102, u1_u5_u2_n103, u1_u5_u2_n104, u1_u5_u2_n105, u1_u5_u2_n106, 
       u1_u5_u2_n107, u1_u5_u2_n108, u1_u5_u2_n109, u1_u5_u2_n110, u1_u5_u2_n111, u1_u5_u2_n112, u1_u5_u2_n113, u1_u5_u2_n114, u1_u5_u2_n115, 
       u1_u5_u2_n116, u1_u5_u2_n117, u1_u5_u2_n118, u1_u5_u2_n119, u1_u5_u2_n120, u1_u5_u2_n121, u1_u5_u2_n122, u1_u5_u2_n123, u1_u5_u2_n124, 
       u1_u5_u2_n125, u1_u5_u2_n126, u1_u5_u2_n127, u1_u5_u2_n128, u1_u5_u2_n129, u1_u5_u2_n130, u1_u5_u2_n131, u1_u5_u2_n132, u1_u5_u2_n133, 
       u1_u5_u2_n134, u1_u5_u2_n135, u1_u5_u2_n136, u1_u5_u2_n137, u1_u5_u2_n138, u1_u5_u2_n139, u1_u5_u2_n140, u1_u5_u2_n141, u1_u5_u2_n142, 
       u1_u5_u2_n143, u1_u5_u2_n144, u1_u5_u2_n145, u1_u5_u2_n146, u1_u5_u2_n147, u1_u5_u2_n148, u1_u5_u2_n149, u1_u5_u2_n150, u1_u5_u2_n151, 
       u1_u5_u2_n152, u1_u5_u2_n153, u1_u5_u2_n154, u1_u5_u2_n155, u1_u5_u2_n156, u1_u5_u2_n157, u1_u5_u2_n158, u1_u5_u2_n159, u1_u5_u2_n160, 
       u1_u5_u2_n161, u1_u5_u2_n162, u1_u5_u2_n163, u1_u5_u2_n164, u1_u5_u2_n165, u1_u5_u2_n166, u1_u5_u2_n167, u1_u5_u2_n168, u1_u5_u2_n169, 
       u1_u5_u2_n170, u1_u5_u2_n171, u1_u5_u2_n172, u1_u5_u2_n173, u1_u5_u2_n174, u1_u5_u2_n175, u1_u5_u2_n176, u1_u5_u2_n177, u1_u5_u2_n178, 
       u1_u5_u2_n179, u1_u5_u2_n180, u1_u5_u2_n181, u1_u5_u2_n182, u1_u5_u2_n183, u1_u5_u2_n184, u1_u5_u2_n185, u1_u5_u2_n186, u1_u5_u2_n187, 
       u1_u5_u2_n188, u1_u5_u2_n95, u1_u5_u2_n96, u1_u5_u2_n97, u1_u5_u2_n98, u1_u5_u2_n99, u1_u5_u3_n100, u1_u5_u3_n101, u1_u5_u3_n102, 
       u1_u5_u3_n103, u1_u5_u3_n104, u1_u5_u3_n105, u1_u5_u3_n106, u1_u5_u3_n107, u1_u5_u3_n108, u1_u5_u3_n109, u1_u5_u3_n110, u1_u5_u3_n111, 
       u1_u5_u3_n112, u1_u5_u3_n113, u1_u5_u3_n114, u1_u5_u3_n115, u1_u5_u3_n116, u1_u5_u3_n117, u1_u5_u3_n118, u1_u5_u3_n119, u1_u5_u3_n120, 
       u1_u5_u3_n121, u1_u5_u3_n122, u1_u5_u3_n123, u1_u5_u3_n124, u1_u5_u3_n125, u1_u5_u3_n126, u1_u5_u3_n127, u1_u5_u3_n128, u1_u5_u3_n129, 
       u1_u5_u3_n130, u1_u5_u3_n131, u1_u5_u3_n132, u1_u5_u3_n133, u1_u5_u3_n134, u1_u5_u3_n135, u1_u5_u3_n136, u1_u5_u3_n137, u1_u5_u3_n138, 
       u1_u5_u3_n139, u1_u5_u3_n140, u1_u5_u3_n141, u1_u5_u3_n142, u1_u5_u3_n143, u1_u5_u3_n144, u1_u5_u3_n145, u1_u5_u3_n146, u1_u5_u3_n147, 
       u1_u5_u3_n148, u1_u5_u3_n149, u1_u5_u3_n150, u1_u5_u3_n151, u1_u5_u3_n152, u1_u5_u3_n153, u1_u5_u3_n154, u1_u5_u3_n155, u1_u5_u3_n156, 
       u1_u5_u3_n157, u1_u5_u3_n158, u1_u5_u3_n159, u1_u5_u3_n160, u1_u5_u3_n161, u1_u5_u3_n162, u1_u5_u3_n163, u1_u5_u3_n164, u1_u5_u3_n165, 
       u1_u5_u3_n166, u1_u5_u3_n167, u1_u5_u3_n168, u1_u5_u3_n169, u1_u5_u3_n170, u1_u5_u3_n171, u1_u5_u3_n172, u1_u5_u3_n173, u1_u5_u3_n174, 
       u1_u5_u3_n175, u1_u5_u3_n176, u1_u5_u3_n177, u1_u5_u3_n178, u1_u5_u3_n179, u1_u5_u3_n180, u1_u5_u3_n181, u1_u5_u3_n182, u1_u5_u3_n183, 
       u1_u5_u3_n184, u1_u5_u3_n185, u1_u5_u3_n186, u1_u5_u3_n94, u1_u5_u3_n95, u1_u5_u3_n96, u1_u5_u3_n97, u1_u5_u3_n98, u1_u5_u3_n99, 
       u1_u5_u6_n100, u1_u5_u6_n101, u1_u5_u6_n102, u1_u5_u6_n103, u1_u5_u6_n104, u1_u5_u6_n105, u1_u5_u6_n106, u1_u5_u6_n107, u1_u5_u6_n108, 
       u1_u5_u6_n109, u1_u5_u6_n110, u1_u5_u6_n111, u1_u5_u6_n112, u1_u5_u6_n113, u1_u5_u6_n114, u1_u5_u6_n115, u1_u5_u6_n116, u1_u5_u6_n117, 
       u1_u5_u6_n118, u1_u5_u6_n119, u1_u5_u6_n120, u1_u5_u6_n121, u1_u5_u6_n122, u1_u5_u6_n123, u1_u5_u6_n124, u1_u5_u6_n125, u1_u5_u6_n126, 
       u1_u5_u6_n127, u1_u5_u6_n128, u1_u5_u6_n129, u1_u5_u6_n130, u1_u5_u6_n131, u1_u5_u6_n132, u1_u5_u6_n133, u1_u5_u6_n134, u1_u5_u6_n135, 
       u1_u5_u6_n136, u1_u5_u6_n137, u1_u5_u6_n138, u1_u5_u6_n139, u1_u5_u6_n140, u1_u5_u6_n141, u1_u5_u6_n142, u1_u5_u6_n143, u1_u5_u6_n144, 
       u1_u5_u6_n145, u1_u5_u6_n146, u1_u5_u6_n147, u1_u5_u6_n148, u1_u5_u6_n149, u1_u5_u6_n150, u1_u5_u6_n151, u1_u5_u6_n152, u1_u5_u6_n153, 
       u1_u5_u6_n154, u1_u5_u6_n155, u1_u5_u6_n156, u1_u5_u6_n157, u1_u5_u6_n158, u1_u5_u6_n159, u1_u5_u6_n160, u1_u5_u6_n161, u1_u5_u6_n162, 
       u1_u5_u6_n163, u1_u5_u6_n164, u1_u5_u6_n165, u1_u5_u6_n166, u1_u5_u6_n167, u1_u5_u6_n168, u1_u5_u6_n169, u1_u5_u6_n170, u1_u5_u6_n171, 
       u1_u5_u6_n172, u1_u5_u6_n173, u1_u5_u6_n174, u1_u5_u6_n88, u1_u5_u6_n89, u1_u5_u6_n90, u1_u5_u6_n91, u1_u5_u6_n92, u1_u5_u6_n93, 
       u1_u5_u6_n94, u1_u5_u6_n95, u1_u5_u6_n96, u1_u5_u6_n97, u1_u5_u6_n98, u1_u5_u6_n99, u1_u6_X_13, u1_u6_X_14, u1_u6_X_15, 
       u1_u6_X_16, u1_u6_X_17, u1_u6_X_18, u1_u6_X_19, u1_u6_X_20, u1_u6_X_21, u1_u6_X_22, u1_u6_X_23, u1_u6_X_24, 
       u1_u6_u2_n100, u1_u6_u2_n101, u1_u6_u2_n102, u1_u6_u2_n103, u1_u6_u2_n104, u1_u6_u2_n105, u1_u6_u2_n106, u1_u6_u2_n107, u1_u6_u2_n108, 
       u1_u6_u2_n109, u1_u6_u2_n110, u1_u6_u2_n111, u1_u6_u2_n112, u1_u6_u2_n113, u1_u6_u2_n114, u1_u6_u2_n115, u1_u6_u2_n116, u1_u6_u2_n117, 
       u1_u6_u2_n118, u1_u6_u2_n119, u1_u6_u2_n120, u1_u6_u2_n121, u1_u6_u2_n122, u1_u6_u2_n123, u1_u6_u2_n124, u1_u6_u2_n125, u1_u6_u2_n126, 
       u1_u6_u2_n127, u1_u6_u2_n128, u1_u6_u2_n129, u1_u6_u2_n130, u1_u6_u2_n131, u1_u6_u2_n132, u1_u6_u2_n133, u1_u6_u2_n134, u1_u6_u2_n135, 
       u1_u6_u2_n136, u1_u6_u2_n137, u1_u6_u2_n138, u1_u6_u2_n139, u1_u6_u2_n140, u1_u6_u2_n141, u1_u6_u2_n142, u1_u6_u2_n143, u1_u6_u2_n144, 
       u1_u6_u2_n145, u1_u6_u2_n146, u1_u6_u2_n147, u1_u6_u2_n148, u1_u6_u2_n149, u1_u6_u2_n150, u1_u6_u2_n151, u1_u6_u2_n152, u1_u6_u2_n153, 
       u1_u6_u2_n154, u1_u6_u2_n155, u1_u6_u2_n156, u1_u6_u2_n157, u1_u6_u2_n158, u1_u6_u2_n159, u1_u6_u2_n160, u1_u6_u2_n161, u1_u6_u2_n162, 
       u1_u6_u2_n163, u1_u6_u2_n164, u1_u6_u2_n165, u1_u6_u2_n166, u1_u6_u2_n167, u1_u6_u2_n168, u1_u6_u2_n169, u1_u6_u2_n170, u1_u6_u2_n171, 
       u1_u6_u2_n172, u1_u6_u2_n173, u1_u6_u2_n174, u1_u6_u2_n175, u1_u6_u2_n176, u1_u6_u2_n177, u1_u6_u2_n178, u1_u6_u2_n179, u1_u6_u2_n180, 
       u1_u6_u2_n181, u1_u6_u2_n182, u1_u6_u2_n183, u1_u6_u2_n184, u1_u6_u2_n185, u1_u6_u2_n186, u1_u6_u2_n187, u1_u6_u2_n188, u1_u6_u2_n95, 
       u1_u6_u2_n96, u1_u6_u2_n97, u1_u6_u2_n98, u1_u6_u2_n99, u1_u6_u3_n100, u1_u6_u3_n101, u1_u6_u3_n102, u1_u6_u3_n103, u1_u6_u3_n104, 
       u1_u6_u3_n105, u1_u6_u3_n106, u1_u6_u3_n107, u1_u6_u3_n108, u1_u6_u3_n109, u1_u6_u3_n110, u1_u6_u3_n111, u1_u6_u3_n112, u1_u6_u3_n113, 
       u1_u6_u3_n114, u1_u6_u3_n115, u1_u6_u3_n116, u1_u6_u3_n117, u1_u6_u3_n118, u1_u6_u3_n119, u1_u6_u3_n120, u1_u6_u3_n121, u1_u6_u3_n122, 
       u1_u6_u3_n123, u1_u6_u3_n124, u1_u6_u3_n125, u1_u6_u3_n126, u1_u6_u3_n127, u1_u6_u3_n128, u1_u6_u3_n129, u1_u6_u3_n130, u1_u6_u3_n131, 
       u1_u6_u3_n132, u1_u6_u3_n133, u1_u6_u3_n134, u1_u6_u3_n135, u1_u6_u3_n136, u1_u6_u3_n137, u1_u6_u3_n138, u1_u6_u3_n139, u1_u6_u3_n140, 
       u1_u6_u3_n141, u1_u6_u3_n142, u1_u6_u3_n143, u1_u6_u3_n144, u1_u6_u3_n145, u1_u6_u3_n146, u1_u6_u3_n147, u1_u6_u3_n148, u1_u6_u3_n149, 
       u1_u6_u3_n150, u1_u6_u3_n151, u1_u6_u3_n152, u1_u6_u3_n153, u1_u6_u3_n154, u1_u6_u3_n155, u1_u6_u3_n156, u1_u6_u3_n157, u1_u6_u3_n158, 
       u1_u6_u3_n159, u1_u6_u3_n160, u1_u6_u3_n161, u1_u6_u3_n162, u1_u6_u3_n163, u1_u6_u3_n164, u1_u6_u3_n165, u1_u6_u3_n166, u1_u6_u3_n167, 
       u1_u6_u3_n168, u1_u6_u3_n169, u1_u6_u3_n170, u1_u6_u3_n171, u1_u6_u3_n172, u1_u6_u3_n173, u1_u6_u3_n174, u1_u6_u3_n175, u1_u6_u3_n176, 
       u1_u6_u3_n177, u1_u6_u3_n178, u1_u6_u3_n179, u1_u6_u3_n180, u1_u6_u3_n181, u1_u6_u3_n182, u1_u6_u3_n183, u1_u6_u3_n184, u1_u6_u3_n185, 
       u1_u6_u3_n186, u1_u6_u3_n94, u1_u6_u3_n95, u1_u6_u3_n96, u1_u6_u3_n97, u1_u6_u3_n98, u1_u6_u3_n99, u1_u7_X_1, u1_u7_X_10, 
       u1_u7_X_11, u1_u7_X_12, u1_u7_X_13, u1_u7_X_14, u1_u7_X_15, u1_u7_X_16, u1_u7_X_17, u1_u7_X_18, u1_u7_X_2, 
       u1_u7_X_25, u1_u7_X_26, u1_u7_X_27, u1_u7_X_28, u1_u7_X_29, u1_u7_X_3, u1_u7_X_30, u1_u7_X_37, u1_u7_X_38, 
       u1_u7_X_39, u1_u7_X_4, u1_u7_X_40, u1_u7_X_41, u1_u7_X_42, u1_u7_X_5, u1_u7_X_6, u1_u7_X_7, u1_u7_X_8, 
       u1_u7_X_9, u1_u7_u0_n100, u1_u7_u0_n101, u1_u7_u0_n102, u1_u7_u0_n103, u1_u7_u0_n104, u1_u7_u0_n105, u1_u7_u0_n106, u1_u7_u0_n107, 
       u1_u7_u0_n108, u1_u7_u0_n109, u1_u7_u0_n110, u1_u7_u0_n111, u1_u7_u0_n112, u1_u7_u0_n113, u1_u7_u0_n114, u1_u7_u0_n115, u1_u7_u0_n116, 
       u1_u7_u0_n117, u1_u7_u0_n118, u1_u7_u0_n119, u1_u7_u0_n120, u1_u7_u0_n121, u1_u7_u0_n122, u1_u7_u0_n123, u1_u7_u0_n124, u1_u7_u0_n125, 
       u1_u7_u0_n126, u1_u7_u0_n127, u1_u7_u0_n128, u1_u7_u0_n129, u1_u7_u0_n130, u1_u7_u0_n131, u1_u7_u0_n132, u1_u7_u0_n133, u1_u7_u0_n134, 
       u1_u7_u0_n135, u1_u7_u0_n136, u1_u7_u0_n137, u1_u7_u0_n138, u1_u7_u0_n139, u1_u7_u0_n140, u1_u7_u0_n141, u1_u7_u0_n142, u1_u7_u0_n143, 
       u1_u7_u0_n144, u1_u7_u0_n145, u1_u7_u0_n146, u1_u7_u0_n147, u1_u7_u0_n148, u1_u7_u0_n149, u1_u7_u0_n150, u1_u7_u0_n151, u1_u7_u0_n152, 
       u1_u7_u0_n153, u1_u7_u0_n154, u1_u7_u0_n155, u1_u7_u0_n156, u1_u7_u0_n157, u1_u7_u0_n158, u1_u7_u0_n159, u1_u7_u0_n160, u1_u7_u0_n161, 
       u1_u7_u0_n162, u1_u7_u0_n163, u1_u7_u0_n164, u1_u7_u0_n165, u1_u7_u0_n166, u1_u7_u0_n167, u1_u7_u0_n168, u1_u7_u0_n169, u1_u7_u0_n170, 
       u1_u7_u0_n171, u1_u7_u0_n172, u1_u7_u0_n173, u1_u7_u0_n174, u1_u7_u0_n88, u1_u7_u0_n89, u1_u7_u0_n90, u1_u7_u0_n91, u1_u7_u0_n92, 
       u1_u7_u0_n93, u1_u7_u0_n94, u1_u7_u0_n95, u1_u7_u0_n96, u1_u7_u0_n97, u1_u7_u0_n98, u1_u7_u0_n99, u1_u7_u1_n100, u1_u7_u1_n101, 
       u1_u7_u1_n102, u1_u7_u1_n103, u1_u7_u1_n104, u1_u7_u1_n105, u1_u7_u1_n106, u1_u7_u1_n107, u1_u7_u1_n108, u1_u7_u1_n109, u1_u7_u1_n110, 
       u1_u7_u1_n111, u1_u7_u1_n112, u1_u7_u1_n113, u1_u7_u1_n114, u1_u7_u1_n115, u1_u7_u1_n116, u1_u7_u1_n117, u1_u7_u1_n118, u1_u7_u1_n119, 
       u1_u7_u1_n120, u1_u7_u1_n121, u1_u7_u1_n122, u1_u7_u1_n123, u1_u7_u1_n124, u1_u7_u1_n125, u1_u7_u1_n126, u1_u7_u1_n127, u1_u7_u1_n128, 
       u1_u7_u1_n129, u1_u7_u1_n130, u1_u7_u1_n131, u1_u7_u1_n132, u1_u7_u1_n133, u1_u7_u1_n134, u1_u7_u1_n135, u1_u7_u1_n136, u1_u7_u1_n137, 
       u1_u7_u1_n138, u1_u7_u1_n139, u1_u7_u1_n140, u1_u7_u1_n141, u1_u7_u1_n142, u1_u7_u1_n143, u1_u7_u1_n144, u1_u7_u1_n145, u1_u7_u1_n146, 
       u1_u7_u1_n147, u1_u7_u1_n148, u1_u7_u1_n149, u1_u7_u1_n150, u1_u7_u1_n151, u1_u7_u1_n152, u1_u7_u1_n153, u1_u7_u1_n154, u1_u7_u1_n155, 
       u1_u7_u1_n156, u1_u7_u1_n157, u1_u7_u1_n158, u1_u7_u1_n159, u1_u7_u1_n160, u1_u7_u1_n161, u1_u7_u1_n162, u1_u7_u1_n163, u1_u7_u1_n164, 
       u1_u7_u1_n165, u1_u7_u1_n166, u1_u7_u1_n167, u1_u7_u1_n168, u1_u7_u1_n169, u1_u7_u1_n170, u1_u7_u1_n171, u1_u7_u1_n172, u1_u7_u1_n173, 
       u1_u7_u1_n174, u1_u7_u1_n175, u1_u7_u1_n176, u1_u7_u1_n177, u1_u7_u1_n178, u1_u7_u1_n179, u1_u7_u1_n180, u1_u7_u1_n181, u1_u7_u1_n182, 
       u1_u7_u1_n183, u1_u7_u1_n184, u1_u7_u1_n185, u1_u7_u1_n186, u1_u7_u1_n187, u1_u7_u1_n188, u1_u7_u1_n95, u1_u7_u1_n96, u1_u7_u1_n97, 
       u1_u7_u1_n98, u1_u7_u1_n99, u1_u7_u2_n100, u1_u7_u2_n101, u1_u7_u2_n102, u1_u7_u2_n103, u1_u7_u2_n104, u1_u7_u2_n105, u1_u7_u2_n106, 
       u1_u7_u2_n107, u1_u7_u2_n108, u1_u7_u2_n109, u1_u7_u2_n110, u1_u7_u2_n111, u1_u7_u2_n112, u1_u7_u2_n113, u1_u7_u2_n114, u1_u7_u2_n115, 
       u1_u7_u2_n116, u1_u7_u2_n117, u1_u7_u2_n118, u1_u7_u2_n119, u1_u7_u2_n120, u1_u7_u2_n121, u1_u7_u2_n122, u1_u7_u2_n123, u1_u7_u2_n124, 
       u1_u7_u2_n125, u1_u7_u2_n126, u1_u7_u2_n127, u1_u7_u2_n128, u1_u7_u2_n129, u1_u7_u2_n130, u1_u7_u2_n131, u1_u7_u2_n132, u1_u7_u2_n133, 
       u1_u7_u2_n134, u1_u7_u2_n135, u1_u7_u2_n136, u1_u7_u2_n137, u1_u7_u2_n138, u1_u7_u2_n139, u1_u7_u2_n140, u1_u7_u2_n141, u1_u7_u2_n142, 
       u1_u7_u2_n143, u1_u7_u2_n144, u1_u7_u2_n145, u1_u7_u2_n146, u1_u7_u2_n147, u1_u7_u2_n148, u1_u7_u2_n149, u1_u7_u2_n150, u1_u7_u2_n151, 
       u1_u7_u2_n152, u1_u7_u2_n153, u1_u7_u2_n154, u1_u7_u2_n155, u1_u7_u2_n156, u1_u7_u2_n157, u1_u7_u2_n158, u1_u7_u2_n159, u1_u7_u2_n160, 
       u1_u7_u2_n161, u1_u7_u2_n162, u1_u7_u2_n163, u1_u7_u2_n164, u1_u7_u2_n165, u1_u7_u2_n166, u1_u7_u2_n167, u1_u7_u2_n168, u1_u7_u2_n169, 
       u1_u7_u2_n170, u1_u7_u2_n171, u1_u7_u2_n172, u1_u7_u2_n173, u1_u7_u2_n174, u1_u7_u2_n175, u1_u7_u2_n176, u1_u7_u2_n177, u1_u7_u2_n178, 
       u1_u7_u2_n179, u1_u7_u2_n180, u1_u7_u2_n181, u1_u7_u2_n182, u1_u7_u2_n183, u1_u7_u2_n184, u1_u7_u2_n185, u1_u7_u2_n186, u1_u7_u2_n187, 
       u1_u7_u2_n188, u1_u7_u2_n95, u1_u7_u2_n96, u1_u7_u2_n97, u1_u7_u2_n98, u1_u7_u2_n99, u1_u7_u4_n100, u1_u7_u4_n101, u1_u7_u4_n102, 
       u1_u7_u4_n103, u1_u7_u4_n104, u1_u7_u4_n105, u1_u7_u4_n106, u1_u7_u4_n107, u1_u7_u4_n108, u1_u7_u4_n109, u1_u7_u4_n110, u1_u7_u4_n111, 
       u1_u7_u4_n112, u1_u7_u4_n113, u1_u7_u4_n114, u1_u7_u4_n115, u1_u7_u4_n116, u1_u7_u4_n117, u1_u7_u4_n118, u1_u7_u4_n119, u1_u7_u4_n120, 
       u1_u7_u4_n121, u1_u7_u4_n122, u1_u7_u4_n123, u1_u7_u4_n124, u1_u7_u4_n125, u1_u7_u4_n126, u1_u7_u4_n127, u1_u7_u4_n128, u1_u7_u4_n129, 
       u1_u7_u4_n130, u1_u7_u4_n131, u1_u7_u4_n132, u1_u7_u4_n133, u1_u7_u4_n134, u1_u7_u4_n135, u1_u7_u4_n136, u1_u7_u4_n137, u1_u7_u4_n138, 
       u1_u7_u4_n139, u1_u7_u4_n140, u1_u7_u4_n141, u1_u7_u4_n142, u1_u7_u4_n143, u1_u7_u4_n144, u1_u7_u4_n145, u1_u7_u4_n146, u1_u7_u4_n147, 
       u1_u7_u4_n148, u1_u7_u4_n149, u1_u7_u4_n150, u1_u7_u4_n151, u1_u7_u4_n152, u1_u7_u4_n153, u1_u7_u4_n154, u1_u7_u4_n155, u1_u7_u4_n156, 
       u1_u7_u4_n157, u1_u7_u4_n158, u1_u7_u4_n159, u1_u7_u4_n160, u1_u7_u4_n161, u1_u7_u4_n162, u1_u7_u4_n163, u1_u7_u4_n164, u1_u7_u4_n165, 
       u1_u7_u4_n166, u1_u7_u4_n167, u1_u7_u4_n168, u1_u7_u4_n169, u1_u7_u4_n170, u1_u7_u4_n171, u1_u7_u4_n172, u1_u7_u4_n173, u1_u7_u4_n174, 
       u1_u7_u4_n175, u1_u7_u4_n176, u1_u7_u4_n177, u1_u7_u4_n178, u1_u7_u4_n179, u1_u7_u4_n180, u1_u7_u4_n181, u1_u7_u4_n182, u1_u7_u4_n183, 
       u1_u7_u4_n184, u1_u7_u4_n185, u1_u7_u4_n186, u1_u7_u4_n94, u1_u7_u4_n95, u1_u7_u4_n96, u1_u7_u4_n97, u1_u7_u4_n98, u1_u7_u4_n99, 
       u1_u7_u6_n100, u1_u7_u6_n101, u1_u7_u6_n102, u1_u7_u6_n103, u1_u7_u6_n104, u1_u7_u6_n105, u1_u7_u6_n106, u1_u7_u6_n107, u1_u7_u6_n108, 
       u1_u7_u6_n109, u1_u7_u6_n110, u1_u7_u6_n111, u1_u7_u6_n112, u1_u7_u6_n113, u1_u7_u6_n114, u1_u7_u6_n115, u1_u7_u6_n116, u1_u7_u6_n117, 
       u1_u7_u6_n118, u1_u7_u6_n119, u1_u7_u6_n120, u1_u7_u6_n121, u1_u7_u6_n122, u1_u7_u6_n123, u1_u7_u6_n124, u1_u7_u6_n125, u1_u7_u6_n126, 
       u1_u7_u6_n127, u1_u7_u6_n128, u1_u7_u6_n129, u1_u7_u6_n130, u1_u7_u6_n131, u1_u7_u6_n132, u1_u7_u6_n133, u1_u7_u6_n134, u1_u7_u6_n135, 
       u1_u7_u6_n136, u1_u7_u6_n137, u1_u7_u6_n138, u1_u7_u6_n139, u1_u7_u6_n140, u1_u7_u6_n141, u1_u7_u6_n142, u1_u7_u6_n143, u1_u7_u6_n144, 
       u1_u7_u6_n145, u1_u7_u6_n146, u1_u7_u6_n147, u1_u7_u6_n148, u1_u7_u6_n149, u1_u7_u6_n150, u1_u7_u6_n151, u1_u7_u6_n152, u1_u7_u6_n153, 
       u1_u7_u6_n154, u1_u7_u6_n155, u1_u7_u6_n156, u1_u7_u6_n157, u1_u7_u6_n158, u1_u7_u6_n159, u1_u7_u6_n160, u1_u7_u6_n161, u1_u7_u6_n162, 
       u1_u7_u6_n163, u1_u7_u6_n164, u1_u7_u6_n165, u1_u7_u6_n166, u1_u7_u6_n167, u1_u7_u6_n168, u1_u7_u6_n169, u1_u7_u6_n170, u1_u7_u6_n171, 
       u1_u7_u6_n172, u1_u7_u6_n173, u1_u7_u6_n174, u1_u7_u6_n88, u1_u7_u6_n89, u1_u7_u6_n90, u1_u7_u6_n91, u1_u7_u6_n92, u1_u7_u6_n93, 
       u1_u7_u6_n94, u1_u7_u6_n95, u1_u7_u6_n96, u1_u7_u6_n97, u1_u7_u6_n98, u1_u7_u6_n99, u1_u8_X_10, u1_u8_X_11, u1_u8_X_12, 
       u1_u8_X_13, u1_u8_X_14, u1_u8_X_15, u1_u8_X_16, u1_u8_X_17, u1_u8_X_18, u1_u8_X_19, u1_u8_X_20, u1_u8_X_21, 
       u1_u8_X_22, u1_u8_X_23, u1_u8_X_24, u1_u8_X_37, u1_u8_X_38, u1_u8_X_39, u1_u8_X_40, u1_u8_X_41, u1_u8_X_42, 
       u1_u8_X_43, u1_u8_X_44, u1_u8_X_45, u1_u8_X_46, u1_u8_X_47, u1_u8_X_48, u1_u8_X_7, u1_u8_X_8, u1_u8_X_9, 
       u1_u8_u1_n100, u1_u8_u1_n101, u1_u8_u1_n102, u1_u8_u1_n103, u1_u8_u1_n104, u1_u8_u1_n105, u1_u8_u1_n106, u1_u8_u1_n107, u1_u8_u1_n108, 
       u1_u8_u1_n109, u1_u8_u1_n110, u1_u8_u1_n111, u1_u8_u1_n112, u1_u8_u1_n113, u1_u8_u1_n114, u1_u8_u1_n115, u1_u8_u1_n116, u1_u8_u1_n117, 
       u1_u8_u1_n118, u1_u8_u1_n119, u1_u8_u1_n120, u1_u8_u1_n121, u1_u8_u1_n122, u1_u8_u1_n123, u1_u8_u1_n124, u1_u8_u1_n125, u1_u8_u1_n126, 
       u1_u8_u1_n127, u1_u8_u1_n128, u1_u8_u1_n129, u1_u8_u1_n130, u1_u8_u1_n131, u1_u8_u1_n132, u1_u8_u1_n133, u1_u8_u1_n134, u1_u8_u1_n135, 
       u1_u8_u1_n136, u1_u8_u1_n137, u1_u8_u1_n138, u1_u8_u1_n139, u1_u8_u1_n140, u1_u8_u1_n141, u1_u8_u1_n142, u1_u8_u1_n143, u1_u8_u1_n144, 
       u1_u8_u1_n145, u1_u8_u1_n146, u1_u8_u1_n147, u1_u8_u1_n148, u1_u8_u1_n149, u1_u8_u1_n150, u1_u8_u1_n151, u1_u8_u1_n152, u1_u8_u1_n153, 
       u1_u8_u1_n154, u1_u8_u1_n155, u1_u8_u1_n156, u1_u8_u1_n157, u1_u8_u1_n158, u1_u8_u1_n159, u1_u8_u1_n160, u1_u8_u1_n161, u1_u8_u1_n162, 
       u1_u8_u1_n163, u1_u8_u1_n164, u1_u8_u1_n165, u1_u8_u1_n166, u1_u8_u1_n167, u1_u8_u1_n168, u1_u8_u1_n169, u1_u8_u1_n170, u1_u8_u1_n171, 
       u1_u8_u1_n172, u1_u8_u1_n173, u1_u8_u1_n174, u1_u8_u1_n175, u1_u8_u1_n176, u1_u8_u1_n177, u1_u8_u1_n178, u1_u8_u1_n179, u1_u8_u1_n180, 
       u1_u8_u1_n181, u1_u8_u1_n182, u1_u8_u1_n183, u1_u8_u1_n184, u1_u8_u1_n185, u1_u8_u1_n186, u1_u8_u1_n187, u1_u8_u1_n188, u1_u8_u1_n95, 
       u1_u8_u1_n96, u1_u8_u1_n97, u1_u8_u1_n98, u1_u8_u1_n99, u1_u8_u2_n100, u1_u8_u2_n101, u1_u8_u2_n102, u1_u8_u2_n103, u1_u8_u2_n104, 
       u1_u8_u2_n105, u1_u8_u2_n106, u1_u8_u2_n107, u1_u8_u2_n108, u1_u8_u2_n109, u1_u8_u2_n110, u1_u8_u2_n111, u1_u8_u2_n112, u1_u8_u2_n113, 
       u1_u8_u2_n114, u1_u8_u2_n115, u1_u8_u2_n116, u1_u8_u2_n117, u1_u8_u2_n118, u1_u8_u2_n119, u1_u8_u2_n120, u1_u8_u2_n121, u1_u8_u2_n122, 
       u1_u8_u2_n123, u1_u8_u2_n124, u1_u8_u2_n125, u1_u8_u2_n126, u1_u8_u2_n127, u1_u8_u2_n128, u1_u8_u2_n129, u1_u8_u2_n130, u1_u8_u2_n131, 
       u1_u8_u2_n132, u1_u8_u2_n133, u1_u8_u2_n134, u1_u8_u2_n135, u1_u8_u2_n136, u1_u8_u2_n137, u1_u8_u2_n138, u1_u8_u2_n139, u1_u8_u2_n140, 
       u1_u8_u2_n141, u1_u8_u2_n142, u1_u8_u2_n143, u1_u8_u2_n144, u1_u8_u2_n145, u1_u8_u2_n146, u1_u8_u2_n147, u1_u8_u2_n148, u1_u8_u2_n149, 
       u1_u8_u2_n150, u1_u8_u2_n151, u1_u8_u2_n152, u1_u8_u2_n153, u1_u8_u2_n154, u1_u8_u2_n155, u1_u8_u2_n156, u1_u8_u2_n157, u1_u8_u2_n158, 
       u1_u8_u2_n159, u1_u8_u2_n160, u1_u8_u2_n161, u1_u8_u2_n162, u1_u8_u2_n163, u1_u8_u2_n164, u1_u8_u2_n165, u1_u8_u2_n166, u1_u8_u2_n167, 
       u1_u8_u2_n168, u1_u8_u2_n169, u1_u8_u2_n170, u1_u8_u2_n171, u1_u8_u2_n172, u1_u8_u2_n173, u1_u8_u2_n174, u1_u8_u2_n175, u1_u8_u2_n176, 
       u1_u8_u2_n177, u1_u8_u2_n178, u1_u8_u2_n179, u1_u8_u2_n180, u1_u8_u2_n181, u1_u8_u2_n182, u1_u8_u2_n183, u1_u8_u2_n184, u1_u8_u2_n185, 
       u1_u8_u2_n186, u1_u8_u2_n187, u1_u8_u2_n188, u1_u8_u2_n95, u1_u8_u2_n96, u1_u8_u2_n97, u1_u8_u2_n98, u1_u8_u2_n99, u1_u8_u3_n100, 
       u1_u8_u3_n101, u1_u8_u3_n102, u1_u8_u3_n103, u1_u8_u3_n104, u1_u8_u3_n105, u1_u8_u3_n106, u1_u8_u3_n107, u1_u8_u3_n108, u1_u8_u3_n109, 
       u1_u8_u3_n110, u1_u8_u3_n111, u1_u8_u3_n112, u1_u8_u3_n113, u1_u8_u3_n114, u1_u8_u3_n115, u1_u8_u3_n116, u1_u8_u3_n117, u1_u8_u3_n118, 
       u1_u8_u3_n119, u1_u8_u3_n120, u1_u8_u3_n121, u1_u8_u3_n122, u1_u8_u3_n123, u1_u8_u3_n124, u1_u8_u3_n125, u1_u8_u3_n126, u1_u8_u3_n127, 
       u1_u8_u3_n128, u1_u8_u3_n129, u1_u8_u3_n130, u1_u8_u3_n131, u1_u8_u3_n132, u1_u8_u3_n133, u1_u8_u3_n134, u1_u8_u3_n135, u1_u8_u3_n136, 
       u1_u8_u3_n137, u1_u8_u3_n138, u1_u8_u3_n139, u1_u8_u3_n140, u1_u8_u3_n141, u1_u8_u3_n142, u1_u8_u3_n143, u1_u8_u3_n144, u1_u8_u3_n145, 
       u1_u8_u3_n146, u1_u8_u3_n147, u1_u8_u3_n148, u1_u8_u3_n149, u1_u8_u3_n150, u1_u8_u3_n151, u1_u8_u3_n152, u1_u8_u3_n153, u1_u8_u3_n154, 
       u1_u8_u3_n155, u1_u8_u3_n156, u1_u8_u3_n157, u1_u8_u3_n158, u1_u8_u3_n159, u1_u8_u3_n160, u1_u8_u3_n161, u1_u8_u3_n162, u1_u8_u3_n163, 
       u1_u8_u3_n164, u1_u8_u3_n165, u1_u8_u3_n166, u1_u8_u3_n167, u1_u8_u3_n168, u1_u8_u3_n169, u1_u8_u3_n170, u1_u8_u3_n171, u1_u8_u3_n172, 
       u1_u8_u3_n173, u1_u8_u3_n174, u1_u8_u3_n175, u1_u8_u3_n176, u1_u8_u3_n177, u1_u8_u3_n178, u1_u8_u3_n179, u1_u8_u3_n180, u1_u8_u3_n181, 
       u1_u8_u3_n182, u1_u8_u3_n183, u1_u8_u3_n184, u1_u8_u3_n185, u1_u8_u3_n186, u1_u8_u3_n94, u1_u8_u3_n95, u1_u8_u3_n96, u1_u8_u3_n97, 
       u1_u8_u3_n98, u1_u8_u3_n99, u1_u8_u6_n100, u1_u8_u6_n101, u1_u8_u6_n102, u1_u8_u6_n103, u1_u8_u6_n104, u1_u8_u6_n105, u1_u8_u6_n106, 
       u1_u8_u6_n107, u1_u8_u6_n108, u1_u8_u6_n109, u1_u8_u6_n110, u1_u8_u6_n111, u1_u8_u6_n112, u1_u8_u6_n113, u1_u8_u6_n114, u1_u8_u6_n115, 
       u1_u8_u6_n116, u1_u8_u6_n117, u1_u8_u6_n118, u1_u8_u6_n119, u1_u8_u6_n120, u1_u8_u6_n121, u1_u8_u6_n122, u1_u8_u6_n123, u1_u8_u6_n124, 
       u1_u8_u6_n125, u1_u8_u6_n126, u1_u8_u6_n127, u1_u8_u6_n128, u1_u8_u6_n129, u1_u8_u6_n130, u1_u8_u6_n131, u1_u8_u6_n132, u1_u8_u6_n133, 
       u1_u8_u6_n134, u1_u8_u6_n135, u1_u8_u6_n136, u1_u8_u6_n137, u1_u8_u6_n138, u1_u8_u6_n139, u1_u8_u6_n140, u1_u8_u6_n141, u1_u8_u6_n142, 
       u1_u8_u6_n143, u1_u8_u6_n144, u1_u8_u6_n145, u1_u8_u6_n146, u1_u8_u6_n147, u1_u8_u6_n148, u1_u8_u6_n149, u1_u8_u6_n150, u1_u8_u6_n151, 
       u1_u8_u6_n152, u1_u8_u6_n153, u1_u8_u6_n154, u1_u8_u6_n155, u1_u8_u6_n156, u1_u8_u6_n157, u1_u8_u6_n158, u1_u8_u6_n159, u1_u8_u6_n160, 
       u1_u8_u6_n161, u1_u8_u6_n162, u1_u8_u6_n163, u1_u8_u6_n164, u1_u8_u6_n165, u1_u8_u6_n166, u1_u8_u6_n167, u1_u8_u6_n168, u1_u8_u6_n169, 
       u1_u8_u6_n170, u1_u8_u6_n171, u1_u8_u6_n172, u1_u8_u6_n173, u1_u8_u6_n174, u1_u8_u6_n88, u1_u8_u6_n89, u1_u8_u6_n90, u1_u8_u6_n91, 
       u1_u8_u6_n92, u1_u8_u6_n93, u1_u8_u6_n94, u1_u8_u6_n95, u1_u8_u6_n96, u1_u8_u6_n97, u1_u8_u6_n98, u1_u8_u6_n99, u1_u8_u7_n100, 
       u1_u8_u7_n101, u1_u8_u7_n102, u1_u8_u7_n103, u1_u8_u7_n104, u1_u8_u7_n105, u1_u8_u7_n106, u1_u8_u7_n107, u1_u8_u7_n108, u1_u8_u7_n109, 
       u1_u8_u7_n110, u1_u8_u7_n111, u1_u8_u7_n112, u1_u8_u7_n113, u1_u8_u7_n114, u1_u8_u7_n115, u1_u8_u7_n116, u1_u8_u7_n117, u1_u8_u7_n118, 
       u1_u8_u7_n119, u1_u8_u7_n120, u1_u8_u7_n121, u1_u8_u7_n122, u1_u8_u7_n123, u1_u8_u7_n124, u1_u8_u7_n125, u1_u8_u7_n126, u1_u8_u7_n127, 
       u1_u8_u7_n128, u1_u8_u7_n129, u1_u8_u7_n130, u1_u8_u7_n131, u1_u8_u7_n132, u1_u8_u7_n133, u1_u8_u7_n134, u1_u8_u7_n135, u1_u8_u7_n136, 
       u1_u8_u7_n137, u1_u8_u7_n138, u1_u8_u7_n139, u1_u8_u7_n140, u1_u8_u7_n141, u1_u8_u7_n142, u1_u8_u7_n143, u1_u8_u7_n144, u1_u8_u7_n145, 
       u1_u8_u7_n146, u1_u8_u7_n147, u1_u8_u7_n148, u1_u8_u7_n149, u1_u8_u7_n150, u1_u8_u7_n151, u1_u8_u7_n152, u1_u8_u7_n153, u1_u8_u7_n154, 
       u1_u8_u7_n155, u1_u8_u7_n156, u1_u8_u7_n157, u1_u8_u7_n158, u1_u8_u7_n159, u1_u8_u7_n160, u1_u8_u7_n161, u1_u8_u7_n162, u1_u8_u7_n163, 
       u1_u8_u7_n164, u1_u8_u7_n165, u1_u8_u7_n166, u1_u8_u7_n167, u1_u8_u7_n168, u1_u8_u7_n169, u1_u8_u7_n170, u1_u8_u7_n171, u1_u8_u7_n172, 
       u1_u8_u7_n173, u1_u8_u7_n174, u1_u8_u7_n175, u1_u8_u7_n176, u1_u8_u7_n177, u1_u8_u7_n178, u1_u8_u7_n179, u1_u8_u7_n180, u1_u8_u7_n91, 
       u1_u8_u7_n92, u1_u8_u7_n93, u1_u8_u7_n94, u1_u8_u7_n95, u1_u8_u7_n96, u1_u8_u7_n97, u1_u8_u7_n98, u1_u8_u7_n99, u1_u9_X_1, 
       u1_u9_X_2, u1_u9_X_3, u1_u9_X_4, u1_u9_X_43, u1_u9_X_44, u1_u9_X_45, u1_u9_X_46, u1_u9_X_47, u1_u9_X_48, 
       u1_u9_X_5, u1_u9_X_6, u1_u9_u0_n100, u1_u9_u0_n101, u1_u9_u0_n102, u1_u9_u0_n103, u1_u9_u0_n104, u1_u9_u0_n105, u1_u9_u0_n106, 
       u1_u9_u0_n107, u1_u9_u0_n108, u1_u9_u0_n109, u1_u9_u0_n110, u1_u9_u0_n111, u1_u9_u0_n112, u1_u9_u0_n113, u1_u9_u0_n114, u1_u9_u0_n115, 
       u1_u9_u0_n116, u1_u9_u0_n117, u1_u9_u0_n118, u1_u9_u0_n119, u1_u9_u0_n120, u1_u9_u0_n121, u1_u9_u0_n122, u1_u9_u0_n123, u1_u9_u0_n124, 
       u1_u9_u0_n125, u1_u9_u0_n126, u1_u9_u0_n127, u1_u9_u0_n128, u1_u9_u0_n129, u1_u9_u0_n130, u1_u9_u0_n131, u1_u9_u0_n132, u1_u9_u0_n133, 
       u1_u9_u0_n134, u1_u9_u0_n135, u1_u9_u0_n136, u1_u9_u0_n137, u1_u9_u0_n138, u1_u9_u0_n139, u1_u9_u0_n140, u1_u9_u0_n141, u1_u9_u0_n142, 
       u1_u9_u0_n143, u1_u9_u0_n144, u1_u9_u0_n145, u1_u9_u0_n146, u1_u9_u0_n147, u1_u9_u0_n148, u1_u9_u0_n149, u1_u9_u0_n150, u1_u9_u0_n151, 
       u1_u9_u0_n152, u1_u9_u0_n153, u1_u9_u0_n154, u1_u9_u0_n155, u1_u9_u0_n156, u1_u9_u0_n157, u1_u9_u0_n158, u1_u9_u0_n159, u1_u9_u0_n160, 
       u1_u9_u0_n161, u1_u9_u0_n162, u1_u9_u0_n163, u1_u9_u0_n164, u1_u9_u0_n165, u1_u9_u0_n166, u1_u9_u0_n167, u1_u9_u0_n168, u1_u9_u0_n169, 
       u1_u9_u0_n170, u1_u9_u0_n171, u1_u9_u0_n172, u1_u9_u0_n173, u1_u9_u0_n174, u1_u9_u0_n88, u1_u9_u0_n89, u1_u9_u0_n90, u1_u9_u0_n91, 
       u1_u9_u0_n92, u1_u9_u0_n93, u1_u9_u0_n94, u1_u9_u0_n95, u1_u9_u0_n96, u1_u9_u0_n97, u1_u9_u0_n98, u1_u9_u0_n99, u1_u9_u7_n100, 
       u1_u9_u7_n101, u1_u9_u7_n102, u1_u9_u7_n103, u1_u9_u7_n104, u1_u9_u7_n105, u1_u9_u7_n106, u1_u9_u7_n107, u1_u9_u7_n108, u1_u9_u7_n109, 
       u1_u9_u7_n110, u1_u9_u7_n111, u1_u9_u7_n112, u1_u9_u7_n113, u1_u9_u7_n114, u1_u9_u7_n115, u1_u9_u7_n116, u1_u9_u7_n117, u1_u9_u7_n118, 
       u1_u9_u7_n119, u1_u9_u7_n120, u1_u9_u7_n121, u1_u9_u7_n122, u1_u9_u7_n123, u1_u9_u7_n124, u1_u9_u7_n125, u1_u9_u7_n126, u1_u9_u7_n127, 
       u1_u9_u7_n128, u1_u9_u7_n129, u1_u9_u7_n130, u1_u9_u7_n131, u1_u9_u7_n132, u1_u9_u7_n133, u1_u9_u7_n134, u1_u9_u7_n135, u1_u9_u7_n136, 
       u1_u9_u7_n137, u1_u9_u7_n138, u1_u9_u7_n139, u1_u9_u7_n140, u1_u9_u7_n141, u1_u9_u7_n142, u1_u9_u7_n143, u1_u9_u7_n144, u1_u9_u7_n145, 
       u1_u9_u7_n146, u1_u9_u7_n147, u1_u9_u7_n148, u1_u9_u7_n149, u1_u9_u7_n150, u1_u9_u7_n151, u1_u9_u7_n152, u1_u9_u7_n153, u1_u9_u7_n154, 
       u1_u9_u7_n155, u1_u9_u7_n156, u1_u9_u7_n157, u1_u9_u7_n158, u1_u9_u7_n159, u1_u9_u7_n160, u1_u9_u7_n161, u1_u9_u7_n162, u1_u9_u7_n163, 
       u1_u9_u7_n164, u1_u9_u7_n165, u1_u9_u7_n166, u1_u9_u7_n167, u1_u9_u7_n168, u1_u9_u7_n169, u1_u9_u7_n170, u1_u9_u7_n171, u1_u9_u7_n172, 
       u1_u9_u7_n173, u1_u9_u7_n174, u1_u9_u7_n175, u1_u9_u7_n176, u1_u9_u7_n177, u1_u9_u7_n178, u1_u9_u7_n179, u1_u9_u7_n180, u1_u9_u7_n91, 
       u1_u9_u7_n92, u1_u9_u7_n93, u1_u9_u7_n94, u1_u9_u7_n95, u1_u9_u7_n96, u1_u9_u7_n97, u1_u9_u7_n98, u1_u9_u7_n99, u1_uk_n10, 
       u1_uk_n100, u1_uk_n1000, u1_uk_n1001, u1_uk_n1002, u1_uk_n1003, u1_uk_n1004, u1_uk_n1005, u1_uk_n1006, u1_uk_n1008, 
       u1_uk_n1009, u1_uk_n1010, u1_uk_n1012, u1_uk_n1013, u1_uk_n1014, u1_uk_n1015, u1_uk_n1016, u1_uk_n1017, u1_uk_n1018, 
       u1_uk_n1019, u1_uk_n102, u1_uk_n1020, u1_uk_n1022, u1_uk_n1023, u1_uk_n1024, u1_uk_n1025, u1_uk_n1026, u1_uk_n1027, 
       u1_uk_n1028, u1_uk_n1029, u1_uk_n1030, u1_uk_n1031, u1_uk_n1032, u1_uk_n1033, u1_uk_n1034, u1_uk_n1035, u1_uk_n1036, 
       u1_uk_n1037, u1_uk_n1038, u1_uk_n1039, u1_uk_n1040, u1_uk_n1041, u1_uk_n1042, u1_uk_n1043, u1_uk_n1044, u1_uk_n1045, 
       u1_uk_n1046, u1_uk_n1047, u1_uk_n1048, u1_uk_n1049, u1_uk_n1051, u1_uk_n1052, u1_uk_n1053, u1_uk_n1054, u1_uk_n1055, 
       u1_uk_n1056, u1_uk_n1057, u1_uk_n1058, u1_uk_n1059, u1_uk_n1061, u1_uk_n1062, u1_uk_n1064, u1_uk_n1066, u1_uk_n1068, 
       u1_uk_n1069, u1_uk_n1070, u1_uk_n1071, u1_uk_n1072, u1_uk_n1073, u1_uk_n1075, u1_uk_n1077, u1_uk_n1078, u1_uk_n1079, 
       u1_uk_n1080, u1_uk_n1081, u1_uk_n1082, u1_uk_n1083, u1_uk_n1084, u1_uk_n1085, u1_uk_n1086, u1_uk_n1087, u1_uk_n1089, 
       u1_uk_n109, u1_uk_n1090, u1_uk_n1091, u1_uk_n1092, u1_uk_n1093, u1_uk_n1094, u1_uk_n1095, u1_uk_n1096, u1_uk_n1097, 
       u1_uk_n1098, u1_uk_n1099, u1_uk_n11, u1_uk_n110, u1_uk_n1100, u1_uk_n1101, u1_uk_n1102, u1_uk_n1103, u1_uk_n1105, 
       u1_uk_n1106, u1_uk_n1107, u1_uk_n1108, u1_uk_n1109, u1_uk_n1110, u1_uk_n1111, u1_uk_n1112, u1_uk_n1113, u1_uk_n1114, 
       u1_uk_n1116, u1_uk_n1117, u1_uk_n1118, u1_uk_n1120, u1_uk_n1121, u1_uk_n1122, u1_uk_n1123, u1_uk_n1125, u1_uk_n1126, 
       u1_uk_n1127, u1_uk_n1128, u1_uk_n1129, u1_uk_n1130, u1_uk_n1131, u1_uk_n1132, u1_uk_n1133, u1_uk_n1134, u1_uk_n1135, 
       u1_uk_n1136, u1_uk_n1138, u1_uk_n1139, u1_uk_n1140, u1_uk_n1141, u1_uk_n1142, u1_uk_n1143, u1_uk_n1144, u1_uk_n1145, 
       u1_uk_n1146, u1_uk_n1147, u1_uk_n1148, u1_uk_n1149, u1_uk_n1150, u1_uk_n1151, u1_uk_n1152, u1_uk_n1153, u1_uk_n1154, 
       u1_uk_n1155, u1_uk_n1156, u1_uk_n1157, u1_uk_n1158, u1_uk_n1160, u1_uk_n1161, u1_uk_n1163, u1_uk_n1164, u1_uk_n1165, 
       u1_uk_n1166, u1_uk_n1167, u1_uk_n1168, u1_uk_n1169, u1_uk_n117, u1_uk_n1170, u1_uk_n1171, u1_uk_n1172, u1_uk_n1173, 
       u1_uk_n1174, u1_uk_n1175, u1_uk_n1176, u1_uk_n1177, u1_uk_n1178, u1_uk_n1179, u1_uk_n118, u1_uk_n1180, u1_uk_n1181, 
       u1_uk_n1182, u1_uk_n1183, u1_uk_n1184, u1_uk_n1185, u1_uk_n1187, u1_uk_n1188, u1_uk_n1189, u1_uk_n1190, u1_uk_n1191, 
       u1_uk_n1192, u1_uk_n1195, u1_uk_n1197, u1_uk_n1198, u1_uk_n1201, u1_uk_n1204, u1_uk_n1205, u1_uk_n1208, u1_uk_n1209, 
       u1_uk_n1213, u1_uk_n1214, u1_uk_n1215, u1_uk_n128, u1_uk_n129, u1_uk_n141, u1_uk_n142, u1_uk_n145, u1_uk_n146, 
       u1_uk_n147, u1_uk_n148, u1_uk_n155, u1_uk_n161, u1_uk_n162, u1_uk_n163, u1_uk_n164, u1_uk_n17, u1_uk_n182, 
       u1_uk_n187, u1_uk_n188, u1_uk_n191, u1_uk_n202, u1_uk_n203, u1_uk_n207, u1_uk_n208, u1_uk_n209, u1_uk_n213, 
       u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n230, u1_uk_n231, u1_uk_n238, u1_uk_n240, 
       u1_uk_n242, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n27, u1_uk_n271, u1_uk_n277, u1_uk_n279, 
       u1_uk_n286, u1_uk_n291, u1_uk_n292, u1_uk_n294, u1_uk_n297, u1_uk_n298, u1_uk_n301, u1_uk_n305, u1_uk_n306, 
       u1_uk_n308, u1_uk_n31, u1_uk_n313, u1_uk_n319, u1_uk_n335, u1_uk_n338, u1_uk_n342, u1_uk_n346, u1_uk_n363, 
       u1_uk_n377, u1_uk_n379, u1_uk_n382, u1_uk_n395, u1_uk_n408, u1_uk_n409, u1_uk_n415, u1_uk_n454, u1_uk_n456, 
       u1_uk_n460, u1_uk_n467, u1_uk_n472, u1_uk_n500, u1_uk_n503, u1_uk_n504, u1_uk_n509, u1_uk_n515, u1_uk_n518, 
       u1_uk_n520, u1_uk_n524, u1_uk_n526, u1_uk_n551, u1_uk_n582, u1_uk_n586, u1_uk_n587, u1_uk_n590, u1_uk_n60, 
       u1_uk_n603, u1_uk_n605, u1_uk_n608, u1_uk_n63, u1_uk_n634, u1_uk_n662, u1_uk_n665, u1_uk_n676, u1_uk_n681, 
       u1_uk_n682, u1_uk_n685, u1_uk_n686, u1_uk_n688, u1_uk_n689, u1_uk_n692, u1_uk_n694, u1_uk_n695, u1_uk_n702, 
       u1_uk_n717, u1_uk_n83, u1_uk_n92, u1_uk_n93, u1_uk_n94, u1_uk_n945, u1_uk_n946, u1_uk_n947, u1_uk_n948, 
       u1_uk_n949, u1_uk_n950, u1_uk_n951, u1_uk_n952, u1_uk_n953, u1_uk_n954, u1_uk_n956, u1_uk_n957, u1_uk_n958, 
       u1_uk_n959, u1_uk_n960, u1_uk_n961, u1_uk_n962, u1_uk_n963, u1_uk_n964, u1_uk_n965, u1_uk_n966, u1_uk_n967, 
       u1_uk_n968, u1_uk_n969, u1_uk_n970, u1_uk_n971, u1_uk_n972, u1_uk_n973, u1_uk_n974, u1_uk_n975, u1_uk_n976, 
       u1_uk_n977, u1_uk_n978, u1_uk_n979, u1_uk_n980, u1_uk_n981, u1_uk_n982, u1_uk_n983, u1_uk_n984, u1_uk_n985, 
       u1_uk_n986, u1_uk_n987, u1_uk_n989, u1_uk_n99, u1_uk_n990, u1_uk_n991, u1_uk_n992, u1_uk_n993, u1_uk_n994, 
       u1_uk_n995, u1_uk_n996, u1_uk_n997, u1_uk_n998, u1_uk_n999, u2_K11_1, u2_K11_10, u2_K11_12, u2_K11_19, 
       u2_K11_2, u2_K11_20, u2_K11_22, u2_K11_23, u2_K11_24, u2_K11_25, u2_K11_26, u2_K11_27, u2_K11_28, 
       u2_K11_3, u2_K11_30, u2_K11_5, u2_K11_8, u2_K13_38, u2_K13_39, u2_K13_41, u2_K13_43, u2_K13_48, 
       u2_K14_1, u2_K14_15, u2_K14_19, u2_K14_2, u2_K14_20, u2_K14_22, u2_K14_23, u2_K14_24, u2_K14_37, 
       u2_K14_38, u2_K14_4, u2_K14_40, u2_K14_41, u2_K14_43, u2_K14_44, u2_K14_45, u2_K14_46, u2_K14_47, 
       u2_K14_48, u2_K14_5, u2_K14_7, u2_K14_9, u2_K2_31, u2_K2_32, u2_K2_33, u2_out10_1, u2_out10_10, 
       u2_out10_13, u2_out10_14, u2_out10_17, u2_out10_18, u2_out10_2, u2_out10_20, u2_out10_23, u2_out10_25, u2_out10_26, 
       u2_out10_28, u2_out10_3, u2_out10_31, u2_out10_8, u2_out10_9, u2_out12_12, u2_out12_15, u2_out12_21, u2_out12_22, 
       u2_out12_27, u2_out12_32, u2_out12_5, u2_out12_7, u2_out13_1, u2_out13_10, u2_out13_12, u2_out13_13, u2_out13_15, 
       u2_out13_16, u2_out13_17, u2_out13_18, u2_out13_2, u2_out13_20, u2_out13_21, u2_out13_22, u2_out13_23, u2_out13_24, 
       u2_out13_26, u2_out13_27, u2_out13_28, u2_out13_30, u2_out13_31, u2_out13_32, u2_out13_5, u2_out13_6, u2_out13_7, 
       u2_out13_9, u2_out1_11, u2_out1_19, u2_out1_29, u2_out1_4, u2_u10_X_1, u2_u10_X_10, u2_u10_X_11, u2_u10_X_12, 
       u2_u10_X_19, u2_u10_X_2, u2_u10_X_20, u2_u10_X_21, u2_u10_X_22, u2_u10_X_23, u2_u10_X_24, u2_u10_X_25, u2_u10_X_26, 
       u2_u10_X_27, u2_u10_X_28, u2_u10_X_29, u2_u10_X_3, u2_u10_X_30, u2_u10_X_4, u2_u10_X_5, u2_u10_X_6, u2_u10_X_7, 
       u2_u10_X_8, u2_u10_X_9, u2_u10_u0_n100, u2_u10_u0_n101, u2_u10_u0_n102, u2_u10_u0_n103, u2_u10_u0_n104, u2_u10_u0_n105, u2_u10_u0_n106, 
       u2_u10_u0_n107, u2_u10_u0_n108, u2_u10_u0_n109, u2_u10_u0_n110, u2_u10_u0_n111, u2_u10_u0_n112, u2_u10_u0_n113, u2_u10_u0_n114, u2_u10_u0_n115, 
       u2_u10_u0_n116, u2_u10_u0_n117, u2_u10_u0_n118, u2_u10_u0_n119, u2_u10_u0_n120, u2_u10_u0_n121, u2_u10_u0_n122, u2_u10_u0_n123, u2_u10_u0_n124, 
       u2_u10_u0_n125, u2_u10_u0_n126, u2_u10_u0_n127, u2_u10_u0_n128, u2_u10_u0_n129, u2_u10_u0_n130, u2_u10_u0_n131, u2_u10_u0_n132, u2_u10_u0_n133, 
       u2_u10_u0_n134, u2_u10_u0_n135, u2_u10_u0_n136, u2_u10_u0_n137, u2_u10_u0_n138, u2_u10_u0_n139, u2_u10_u0_n140, u2_u10_u0_n141, u2_u10_u0_n142, 
       u2_u10_u0_n143, u2_u10_u0_n144, u2_u10_u0_n145, u2_u10_u0_n146, u2_u10_u0_n147, u2_u10_u0_n148, u2_u10_u0_n149, u2_u10_u0_n150, u2_u10_u0_n151, 
       u2_u10_u0_n152, u2_u10_u0_n153, u2_u10_u0_n154, u2_u10_u0_n155, u2_u10_u0_n156, u2_u10_u0_n157, u2_u10_u0_n158, u2_u10_u0_n159, u2_u10_u0_n160, 
       u2_u10_u0_n161, u2_u10_u0_n162, u2_u10_u0_n163, u2_u10_u0_n164, u2_u10_u0_n165, u2_u10_u0_n166, u2_u10_u0_n167, u2_u10_u0_n168, u2_u10_u0_n169, 
       u2_u10_u0_n170, u2_u10_u0_n171, u2_u10_u0_n172, u2_u10_u0_n173, u2_u10_u0_n174, u2_u10_u0_n88, u2_u10_u0_n89, u2_u10_u0_n90, u2_u10_u0_n91, 
       u2_u10_u0_n92, u2_u10_u0_n93, u2_u10_u0_n94, u2_u10_u0_n95, u2_u10_u0_n96, u2_u10_u0_n97, u2_u10_u0_n98, u2_u10_u0_n99, u2_u10_u1_n100, 
       u2_u10_u1_n101, u2_u10_u1_n102, u2_u10_u1_n103, u2_u10_u1_n104, u2_u10_u1_n105, u2_u10_u1_n106, u2_u10_u1_n107, u2_u10_u1_n108, u2_u10_u1_n109, 
       u2_u10_u1_n110, u2_u10_u1_n111, u2_u10_u1_n112, u2_u10_u1_n113, u2_u10_u1_n114, u2_u10_u1_n115, u2_u10_u1_n116, u2_u10_u1_n117, u2_u10_u1_n118, 
       u2_u10_u1_n119, u2_u10_u1_n120, u2_u10_u1_n121, u2_u10_u1_n122, u2_u10_u1_n123, u2_u10_u1_n124, u2_u10_u1_n125, u2_u10_u1_n126, u2_u10_u1_n127, 
       u2_u10_u1_n128, u2_u10_u1_n129, u2_u10_u1_n130, u2_u10_u1_n131, u2_u10_u1_n132, u2_u10_u1_n133, u2_u10_u1_n134, u2_u10_u1_n135, u2_u10_u1_n136, 
       u2_u10_u1_n137, u2_u10_u1_n138, u2_u10_u1_n139, u2_u10_u1_n140, u2_u10_u1_n141, u2_u10_u1_n142, u2_u10_u1_n143, u2_u10_u1_n144, u2_u10_u1_n145, 
       u2_u10_u1_n146, u2_u10_u1_n147, u2_u10_u1_n148, u2_u10_u1_n149, u2_u10_u1_n150, u2_u10_u1_n151, u2_u10_u1_n152, u2_u10_u1_n153, u2_u10_u1_n154, 
       u2_u10_u1_n155, u2_u10_u1_n156, u2_u10_u1_n157, u2_u10_u1_n158, u2_u10_u1_n159, u2_u10_u1_n160, u2_u10_u1_n161, u2_u10_u1_n162, u2_u10_u1_n163, 
       u2_u10_u1_n164, u2_u10_u1_n165, u2_u10_u1_n166, u2_u10_u1_n167, u2_u10_u1_n168, u2_u10_u1_n169, u2_u10_u1_n170, u2_u10_u1_n171, u2_u10_u1_n172, 
       u2_u10_u1_n173, u2_u10_u1_n174, u2_u10_u1_n175, u2_u10_u1_n176, u2_u10_u1_n177, u2_u10_u1_n178, u2_u10_u1_n179, u2_u10_u1_n180, u2_u10_u1_n181, 
       u2_u10_u1_n182, u2_u10_u1_n183, u2_u10_u1_n184, u2_u10_u1_n185, u2_u10_u1_n186, u2_u10_u1_n187, u2_u10_u1_n188, u2_u10_u1_n95, u2_u10_u1_n96, 
       u2_u10_u1_n97, u2_u10_u1_n98, u2_u10_u1_n99, u2_u10_u3_n100, u2_u10_u3_n101, u2_u10_u3_n102, u2_u10_u3_n103, u2_u10_u3_n104, u2_u10_u3_n105, 
       u2_u10_u3_n106, u2_u10_u3_n107, u2_u10_u3_n108, u2_u10_u3_n109, u2_u10_u3_n110, u2_u10_u3_n111, u2_u10_u3_n112, u2_u10_u3_n113, u2_u10_u3_n114, 
       u2_u10_u3_n115, u2_u10_u3_n116, u2_u10_u3_n117, u2_u10_u3_n118, u2_u10_u3_n119, u2_u10_u3_n120, u2_u10_u3_n121, u2_u10_u3_n122, u2_u10_u3_n123, 
       u2_u10_u3_n124, u2_u10_u3_n125, u2_u10_u3_n126, u2_u10_u3_n127, u2_u10_u3_n128, u2_u10_u3_n129, u2_u10_u3_n130, u2_u10_u3_n131, u2_u10_u3_n132, 
       u2_u10_u3_n133, u2_u10_u3_n134, u2_u10_u3_n135, u2_u10_u3_n136, u2_u10_u3_n137, u2_u10_u3_n138, u2_u10_u3_n139, u2_u10_u3_n140, u2_u10_u3_n141, 
       u2_u10_u3_n142, u2_u10_u3_n143, u2_u10_u3_n144, u2_u10_u3_n145, u2_u10_u3_n146, u2_u10_u3_n147, u2_u10_u3_n148, u2_u10_u3_n149, u2_u10_u3_n150, 
       u2_u10_u3_n151, u2_u10_u3_n152, u2_u10_u3_n153, u2_u10_u3_n154, u2_u10_u3_n155, u2_u10_u3_n156, u2_u10_u3_n157, u2_u10_u3_n158, u2_u10_u3_n159, 
       u2_u10_u3_n160, u2_u10_u3_n161, u2_u10_u3_n162, u2_u10_u3_n163, u2_u10_u3_n164, u2_u10_u3_n165, u2_u10_u3_n166, u2_u10_u3_n167, u2_u10_u3_n168, 
       u2_u10_u3_n169, u2_u10_u3_n170, u2_u10_u3_n171, u2_u10_u3_n172, u2_u10_u3_n173, u2_u10_u3_n174, u2_u10_u3_n175, u2_u10_u3_n176, u2_u10_u3_n177, 
       u2_u10_u3_n178, u2_u10_u3_n179, u2_u10_u3_n180, u2_u10_u3_n181, u2_u10_u3_n182, u2_u10_u3_n183, u2_u10_u3_n184, u2_u10_u3_n185, u2_u10_u3_n186, 
       u2_u10_u3_n94, u2_u10_u3_n95, u2_u10_u3_n96, u2_u10_u3_n97, u2_u10_u3_n98, u2_u10_u3_n99, u2_u10_u4_n100, u2_u10_u4_n101, u2_u10_u4_n102, 
       u2_u10_u4_n103, u2_u10_u4_n104, u2_u10_u4_n105, u2_u10_u4_n106, u2_u10_u4_n107, u2_u10_u4_n108, u2_u10_u4_n109, u2_u10_u4_n110, u2_u10_u4_n111, 
       u2_u10_u4_n112, u2_u10_u4_n113, u2_u10_u4_n114, u2_u10_u4_n115, u2_u10_u4_n116, u2_u10_u4_n117, u2_u10_u4_n118, u2_u10_u4_n119, u2_u10_u4_n120, 
       u2_u10_u4_n121, u2_u10_u4_n122, u2_u10_u4_n123, u2_u10_u4_n124, u2_u10_u4_n125, u2_u10_u4_n126, u2_u10_u4_n127, u2_u10_u4_n128, u2_u10_u4_n129, 
       u2_u10_u4_n130, u2_u10_u4_n131, u2_u10_u4_n132, u2_u10_u4_n133, u2_u10_u4_n134, u2_u10_u4_n135, u2_u10_u4_n136, u2_u10_u4_n137, u2_u10_u4_n138, 
       u2_u10_u4_n139, u2_u10_u4_n140, u2_u10_u4_n141, u2_u10_u4_n142, u2_u10_u4_n143, u2_u10_u4_n144, u2_u10_u4_n145, u2_u10_u4_n146, u2_u10_u4_n147, 
       u2_u10_u4_n148, u2_u10_u4_n149, u2_u10_u4_n150, u2_u10_u4_n151, u2_u10_u4_n152, u2_u10_u4_n153, u2_u10_u4_n154, u2_u10_u4_n155, u2_u10_u4_n156, 
       u2_u10_u4_n157, u2_u10_u4_n158, u2_u10_u4_n159, u2_u10_u4_n160, u2_u10_u4_n161, u2_u10_u4_n162, u2_u10_u4_n163, u2_u10_u4_n164, u2_u10_u4_n165, 
       u2_u10_u4_n166, u2_u10_u4_n167, u2_u10_u4_n168, u2_u10_u4_n169, u2_u10_u4_n170, u2_u10_u4_n171, u2_u10_u4_n172, u2_u10_u4_n173, u2_u10_u4_n174, 
       u2_u10_u4_n175, u2_u10_u4_n176, u2_u10_u4_n177, u2_u10_u4_n178, u2_u10_u4_n179, u2_u10_u4_n180, u2_u10_u4_n181, u2_u10_u4_n182, u2_u10_u4_n183, 
       u2_u10_u4_n184, u2_u10_u4_n185, u2_u10_u4_n186, u2_u10_u4_n94, u2_u10_u4_n95, u2_u10_u4_n96, u2_u10_u4_n97, u2_u10_u4_n98, u2_u10_u4_n99, 
       u2_u12_X_37, u2_u12_X_38, u2_u12_X_39, u2_u12_X_40, u2_u12_X_41, u2_u12_X_42, u2_u12_X_43, u2_u12_X_44, u2_u12_X_45, 
       u2_u12_X_46, u2_u12_X_47, u2_u12_X_48, u2_u12_u6_n100, u2_u12_u6_n101, u2_u12_u6_n102, u2_u12_u6_n103, u2_u12_u6_n104, u2_u12_u6_n105, 
       u2_u12_u6_n106, u2_u12_u6_n107, u2_u12_u6_n108, u2_u12_u6_n109, u2_u12_u6_n110, u2_u12_u6_n111, u2_u12_u6_n112, u2_u12_u6_n113, u2_u12_u6_n114, 
       u2_u12_u6_n115, u2_u12_u6_n116, u2_u12_u6_n117, u2_u12_u6_n118, u2_u12_u6_n119, u2_u12_u6_n120, u2_u12_u6_n121, u2_u12_u6_n122, u2_u12_u6_n123, 
       u2_u12_u6_n124, u2_u12_u6_n125, u2_u12_u6_n126, u2_u12_u6_n127, u2_u12_u6_n128, u2_u12_u6_n129, u2_u12_u6_n130, u2_u12_u6_n131, u2_u12_u6_n132, 
       u2_u12_u6_n133, u2_u12_u6_n134, u2_u12_u6_n135, u2_u12_u6_n136, u2_u12_u6_n137, u2_u12_u6_n138, u2_u12_u6_n139, u2_u12_u6_n140, u2_u12_u6_n141, 
       u2_u12_u6_n142, u2_u12_u6_n143, u2_u12_u6_n144, u2_u12_u6_n145, u2_u12_u6_n146, u2_u12_u6_n147, u2_u12_u6_n148, u2_u12_u6_n149, u2_u12_u6_n150, 
       u2_u12_u6_n151, u2_u12_u6_n152, u2_u12_u6_n153, u2_u12_u6_n154, u2_u12_u6_n155, u2_u12_u6_n156, u2_u12_u6_n157, u2_u12_u6_n158, u2_u12_u6_n159, 
       u2_u12_u6_n160, u2_u12_u6_n161, u2_u12_u6_n162, u2_u12_u6_n163, u2_u12_u6_n164, u2_u12_u6_n165, u2_u12_u6_n166, u2_u12_u6_n167, u2_u12_u6_n168, 
       u2_u12_u6_n169, u2_u12_u6_n170, u2_u12_u6_n171, u2_u12_u6_n172, u2_u12_u6_n173, u2_u12_u6_n174, u2_u12_u6_n88, u2_u12_u6_n89, u2_u12_u6_n90, 
       u2_u12_u6_n91, u2_u12_u6_n92, u2_u12_u6_n93, u2_u12_u6_n94, u2_u12_u6_n95, u2_u12_u6_n96, u2_u12_u6_n97, u2_u12_u6_n98, u2_u12_u6_n99, 
       u2_u12_u7_n100, u2_u12_u7_n101, u2_u12_u7_n102, u2_u12_u7_n103, u2_u12_u7_n104, u2_u12_u7_n105, u2_u12_u7_n106, u2_u12_u7_n107, u2_u12_u7_n108, 
       u2_u12_u7_n109, u2_u12_u7_n110, u2_u12_u7_n111, u2_u12_u7_n112, u2_u12_u7_n113, u2_u12_u7_n114, u2_u12_u7_n115, u2_u12_u7_n116, u2_u12_u7_n117, 
       u2_u12_u7_n118, u2_u12_u7_n119, u2_u12_u7_n120, u2_u12_u7_n121, u2_u12_u7_n122, u2_u12_u7_n123, u2_u12_u7_n124, u2_u12_u7_n125, u2_u12_u7_n126, 
       u2_u12_u7_n127, u2_u12_u7_n128, u2_u12_u7_n129, u2_u12_u7_n130, u2_u12_u7_n131, u2_u12_u7_n132, u2_u12_u7_n133, u2_u12_u7_n134, u2_u12_u7_n135, 
       u2_u12_u7_n136, u2_u12_u7_n137, u2_u12_u7_n138, u2_u12_u7_n139, u2_u12_u7_n140, u2_u12_u7_n141, u2_u12_u7_n142, u2_u12_u7_n143, u2_u12_u7_n144, 
       u2_u12_u7_n145, u2_u12_u7_n146, u2_u12_u7_n147, u2_u12_u7_n148, u2_u12_u7_n149, u2_u12_u7_n150, u2_u12_u7_n151, u2_u12_u7_n152, u2_u12_u7_n153, 
       u2_u12_u7_n154, u2_u12_u7_n155, u2_u12_u7_n156, u2_u12_u7_n157, u2_u12_u7_n158, u2_u12_u7_n159, u2_u12_u7_n160, u2_u12_u7_n161, u2_u12_u7_n162, 
       u2_u12_u7_n163, u2_u12_u7_n164, u2_u12_u7_n165, u2_u12_u7_n166, u2_u12_u7_n167, u2_u12_u7_n168, u2_u12_u7_n169, u2_u12_u7_n170, u2_u12_u7_n171, 
       u2_u12_u7_n172, u2_u12_u7_n173, u2_u12_u7_n174, u2_u12_u7_n175, u2_u12_u7_n176, u2_u12_u7_n177, u2_u12_u7_n178, u2_u12_u7_n179, u2_u12_u7_n180, 
       u2_u12_u7_n91, u2_u12_u7_n92, u2_u12_u7_n93, u2_u12_u7_n94, u2_u12_u7_n95, u2_u12_u7_n96, u2_u12_u7_n97, u2_u12_u7_n98, u2_u12_u7_n99, 
       u2_u13_X_1, u2_u13_X_10, u2_u13_X_11, u2_u13_X_12, u2_u13_X_13, u2_u13_X_14, u2_u13_X_15, u2_u13_X_16, u2_u13_X_17, 
       u2_u13_X_18, u2_u13_X_19, u2_u13_X_2, u2_u13_X_20, u2_u13_X_21, u2_u13_X_22, u2_u13_X_23, u2_u13_X_24, u2_u13_X_3, 
       u2_u13_X_37, u2_u13_X_38, u2_u13_X_39, u2_u13_X_4, u2_u13_X_40, u2_u13_X_41, u2_u13_X_42, u2_u13_X_43, u2_u13_X_44, 
       u2_u13_X_45, u2_u13_X_46, u2_u13_X_47, u2_u13_X_48, u2_u13_X_5, u2_u13_X_6, u2_u13_X_7, u2_u13_X_8, u2_u13_X_9, 
       u2_u13_u0_n100, u2_u13_u0_n101, u2_u13_u0_n102, u2_u13_u0_n103, u2_u13_u0_n104, u2_u13_u0_n105, u2_u13_u0_n106, u2_u13_u0_n107, u2_u13_u0_n108, 
       u2_u13_u0_n109, u2_u13_u0_n110, u2_u13_u0_n111, u2_u13_u0_n112, u2_u13_u0_n113, u2_u13_u0_n114, u2_u13_u0_n115, u2_u13_u0_n116, u2_u13_u0_n117, 
       u2_u13_u0_n118, u2_u13_u0_n119, u2_u13_u0_n120, u2_u13_u0_n121, u2_u13_u0_n122, u2_u13_u0_n123, u2_u13_u0_n124, u2_u13_u0_n125, u2_u13_u0_n126, 
       u2_u13_u0_n127, u2_u13_u0_n128, u2_u13_u0_n129, u2_u13_u0_n130, u2_u13_u0_n131, u2_u13_u0_n132, u2_u13_u0_n133, u2_u13_u0_n134, u2_u13_u0_n135, 
       u2_u13_u0_n136, u2_u13_u0_n137, u2_u13_u0_n138, u2_u13_u0_n139, u2_u13_u0_n140, u2_u13_u0_n141, u2_u13_u0_n142, u2_u13_u0_n143, u2_u13_u0_n144, 
       u2_u13_u0_n145, u2_u13_u0_n146, u2_u13_u0_n147, u2_u13_u0_n148, u2_u13_u0_n149, u2_u13_u0_n150, u2_u13_u0_n151, u2_u13_u0_n152, u2_u13_u0_n153, 
       u2_u13_u0_n154, u2_u13_u0_n155, u2_u13_u0_n156, u2_u13_u0_n157, u2_u13_u0_n158, u2_u13_u0_n159, u2_u13_u0_n160, u2_u13_u0_n161, u2_u13_u0_n162, 
       u2_u13_u0_n163, u2_u13_u0_n164, u2_u13_u0_n165, u2_u13_u0_n166, u2_u13_u0_n167, u2_u13_u0_n168, u2_u13_u0_n169, u2_u13_u0_n170, u2_u13_u0_n171, 
       u2_u13_u0_n172, u2_u13_u0_n173, u2_u13_u0_n174, u2_u13_u0_n88, u2_u13_u0_n89, u2_u13_u0_n90, u2_u13_u0_n91, u2_u13_u0_n92, u2_u13_u0_n93, 
       u2_u13_u0_n94, u2_u13_u0_n95, u2_u13_u0_n96, u2_u13_u0_n97, u2_u13_u0_n98, u2_u13_u0_n99, u2_u13_u1_n100, u2_u13_u1_n101, u2_u13_u1_n102, 
       u2_u13_u1_n103, u2_u13_u1_n104, u2_u13_u1_n105, u2_u13_u1_n106, u2_u13_u1_n107, u2_u13_u1_n108, u2_u13_u1_n109, u2_u13_u1_n110, u2_u13_u1_n111, 
       u2_u13_u1_n112, u2_u13_u1_n113, u2_u13_u1_n114, u2_u13_u1_n115, u2_u13_u1_n116, u2_u13_u1_n117, u2_u13_u1_n118, u2_u13_u1_n119, u2_u13_u1_n120, 
       u2_u13_u1_n121, u2_u13_u1_n122, u2_u13_u1_n123, u2_u13_u1_n124, u2_u13_u1_n125, u2_u13_u1_n126, u2_u13_u1_n127, u2_u13_u1_n128, u2_u13_u1_n129, 
       u2_u13_u1_n130, u2_u13_u1_n131, u2_u13_u1_n132, u2_u13_u1_n133, u2_u13_u1_n134, u2_u13_u1_n135, u2_u13_u1_n136, u2_u13_u1_n137, u2_u13_u1_n138, 
       u2_u13_u1_n139, u2_u13_u1_n140, u2_u13_u1_n141, u2_u13_u1_n142, u2_u13_u1_n143, u2_u13_u1_n144, u2_u13_u1_n145, u2_u13_u1_n146, u2_u13_u1_n147, 
       u2_u13_u1_n148, u2_u13_u1_n149, u2_u13_u1_n150, u2_u13_u1_n151, u2_u13_u1_n152, u2_u13_u1_n153, u2_u13_u1_n154, u2_u13_u1_n155, u2_u13_u1_n156, 
       u2_u13_u1_n157, u2_u13_u1_n158, u2_u13_u1_n159, u2_u13_u1_n160, u2_u13_u1_n161, u2_u13_u1_n162, u2_u13_u1_n163, u2_u13_u1_n164, u2_u13_u1_n165, 
       u2_u13_u1_n166, u2_u13_u1_n167, u2_u13_u1_n168, u2_u13_u1_n169, u2_u13_u1_n170, u2_u13_u1_n171, u2_u13_u1_n172, u2_u13_u1_n173, u2_u13_u1_n174, 
       u2_u13_u1_n175, u2_u13_u1_n176, u2_u13_u1_n177, u2_u13_u1_n178, u2_u13_u1_n179, u2_u13_u1_n180, u2_u13_u1_n181, u2_u13_u1_n182, u2_u13_u1_n183, 
       u2_u13_u1_n184, u2_u13_u1_n185, u2_u13_u1_n186, u2_u13_u1_n187, u2_u13_u1_n188, u2_u13_u1_n95, u2_u13_u1_n96, u2_u13_u1_n97, u2_u13_u1_n98, 
       u2_u13_u1_n99, u2_u13_u2_n100, u2_u13_u2_n101, u2_u13_u2_n102, u2_u13_u2_n103, u2_u13_u2_n104, u2_u13_u2_n105, u2_u13_u2_n106, u2_u13_u2_n107, 
       u2_u13_u2_n108, u2_u13_u2_n109, u2_u13_u2_n110, u2_u13_u2_n111, u2_u13_u2_n112, u2_u13_u2_n113, u2_u13_u2_n114, u2_u13_u2_n115, u2_u13_u2_n116, 
       u2_u13_u2_n117, u2_u13_u2_n118, u2_u13_u2_n119, u2_u13_u2_n120, u2_u13_u2_n121, u2_u13_u2_n122, u2_u13_u2_n123, u2_u13_u2_n124, u2_u13_u2_n125, 
       u2_u13_u2_n126, u2_u13_u2_n127, u2_u13_u2_n128, u2_u13_u2_n129, u2_u13_u2_n130, u2_u13_u2_n131, u2_u13_u2_n132, u2_u13_u2_n133, u2_u13_u2_n134, 
       u2_u13_u2_n135, u2_u13_u2_n136, u2_u13_u2_n137, u2_u13_u2_n138, u2_u13_u2_n139, u2_u13_u2_n140, u2_u13_u2_n141, u2_u13_u2_n142, u2_u13_u2_n143, 
       u2_u13_u2_n144, u2_u13_u2_n145, u2_u13_u2_n146, u2_u13_u2_n147, u2_u13_u2_n148, u2_u13_u2_n149, u2_u13_u2_n150, u2_u13_u2_n151, u2_u13_u2_n152, 
       u2_u13_u2_n153, u2_u13_u2_n154, u2_u13_u2_n155, u2_u13_u2_n156, u2_u13_u2_n157, u2_u13_u2_n158, u2_u13_u2_n159, u2_u13_u2_n160, u2_u13_u2_n161, 
       u2_u13_u2_n162, u2_u13_u2_n163, u2_u13_u2_n164, u2_u13_u2_n165, u2_u13_u2_n166, u2_u13_u2_n167, u2_u13_u2_n168, u2_u13_u2_n169, u2_u13_u2_n170, 
       u2_u13_u2_n171, u2_u13_u2_n172, u2_u13_u2_n173, u2_u13_u2_n174, u2_u13_u2_n175, u2_u13_u2_n176, u2_u13_u2_n177, u2_u13_u2_n178, u2_u13_u2_n179, 
       u2_u13_u2_n180, u2_u13_u2_n181, u2_u13_u2_n182, u2_u13_u2_n183, u2_u13_u2_n184, u2_u13_u2_n185, u2_u13_u2_n186, u2_u13_u2_n187, u2_u13_u2_n188, 
       u2_u13_u2_n95, u2_u13_u2_n96, u2_u13_u2_n97, u2_u13_u2_n98, u2_u13_u2_n99, u2_u13_u3_n100, u2_u13_u3_n101, u2_u13_u3_n102, u2_u13_u3_n103, 
       u2_u13_u3_n104, u2_u13_u3_n105, u2_u13_u3_n106, u2_u13_u3_n107, u2_u13_u3_n108, u2_u13_u3_n109, u2_u13_u3_n110, u2_u13_u3_n111, u2_u13_u3_n112, 
       u2_u13_u3_n113, u2_u13_u3_n114, u2_u13_u3_n115, u2_u13_u3_n116, u2_u13_u3_n117, u2_u13_u3_n118, u2_u13_u3_n119, u2_u13_u3_n120, u2_u13_u3_n121, 
       u2_u13_u3_n122, u2_u13_u3_n123, u2_u13_u3_n124, u2_u13_u3_n125, u2_u13_u3_n126, u2_u13_u3_n127, u2_u13_u3_n128, u2_u13_u3_n129, u2_u13_u3_n130, 
       u2_u13_u3_n131, u2_u13_u3_n132, u2_u13_u3_n133, u2_u13_u3_n134, u2_u13_u3_n135, u2_u13_u3_n136, u2_u13_u3_n137, u2_u13_u3_n138, u2_u13_u3_n139, 
       u2_u13_u3_n140, u2_u13_u3_n141, u2_u13_u3_n142, u2_u13_u3_n143, u2_u13_u3_n144, u2_u13_u3_n145, u2_u13_u3_n146, u2_u13_u3_n147, u2_u13_u3_n148, 
       u2_u13_u3_n149, u2_u13_u3_n150, u2_u13_u3_n151, u2_u13_u3_n152, u2_u13_u3_n153, u2_u13_u3_n154, u2_u13_u3_n155, u2_u13_u3_n156, u2_u13_u3_n157, 
       u2_u13_u3_n158, u2_u13_u3_n159, u2_u13_u3_n160, u2_u13_u3_n161, u2_u13_u3_n162, u2_u13_u3_n163, u2_u13_u3_n164, u2_u13_u3_n165, u2_u13_u3_n166, 
       u2_u13_u3_n167, u2_u13_u3_n168, u2_u13_u3_n169, u2_u13_u3_n170, u2_u13_u3_n171, u2_u13_u3_n172, u2_u13_u3_n173, u2_u13_u3_n174, u2_u13_u3_n175, 
       u2_u13_u3_n176, u2_u13_u3_n177, u2_u13_u3_n178, u2_u13_u3_n179, u2_u13_u3_n180, u2_u13_u3_n181, u2_u13_u3_n182, u2_u13_u3_n183, u2_u13_u3_n184, 
       u2_u13_u3_n185, u2_u13_u3_n186, u2_u13_u3_n94, u2_u13_u3_n95, u2_u13_u3_n96, u2_u13_u3_n97, u2_u13_u3_n98, u2_u13_u3_n99, u2_u13_u6_n100, 
       u2_u13_u6_n101, u2_u13_u6_n102, u2_u13_u6_n103, u2_u13_u6_n104, u2_u13_u6_n105, u2_u13_u6_n106, u2_u13_u6_n107, u2_u13_u6_n108, u2_u13_u6_n109, 
       u2_u13_u6_n110, u2_u13_u6_n111, u2_u13_u6_n112, u2_u13_u6_n113, u2_u13_u6_n114, u2_u13_u6_n115, u2_u13_u6_n116, u2_u13_u6_n117, u2_u13_u6_n118, 
       u2_u13_u6_n119, u2_u13_u6_n120, u2_u13_u6_n121, u2_u13_u6_n122, u2_u13_u6_n123, u2_u13_u6_n124, u2_u13_u6_n125, u2_u13_u6_n126, u2_u13_u6_n127, 
       u2_u13_u6_n128, u2_u13_u6_n129, u2_u13_u6_n130, u2_u13_u6_n131, u2_u13_u6_n132, u2_u13_u6_n133, u2_u13_u6_n134, u2_u13_u6_n135, u2_u13_u6_n136, 
       u2_u13_u6_n137, u2_u13_u6_n138, u2_u13_u6_n139, u2_u13_u6_n140, u2_u13_u6_n141, u2_u13_u6_n142, u2_u13_u6_n143, u2_u13_u6_n144, u2_u13_u6_n145, 
       u2_u13_u6_n146, u2_u13_u6_n147, u2_u13_u6_n148, u2_u13_u6_n149, u2_u13_u6_n150, u2_u13_u6_n151, u2_u13_u6_n152, u2_u13_u6_n153, u2_u13_u6_n154, 
       u2_u13_u6_n155, u2_u13_u6_n156, u2_u13_u6_n157, u2_u13_u6_n158, u2_u13_u6_n159, u2_u13_u6_n160, u2_u13_u6_n161, u2_u13_u6_n162, u2_u13_u6_n163, 
       u2_u13_u6_n164, u2_u13_u6_n165, u2_u13_u6_n166, u2_u13_u6_n167, u2_u13_u6_n168, u2_u13_u6_n169, u2_u13_u6_n170, u2_u13_u6_n171, u2_u13_u6_n172, 
       u2_u13_u6_n173, u2_u13_u6_n174, u2_u13_u6_n88, u2_u13_u6_n89, u2_u13_u6_n90, u2_u13_u6_n91, u2_u13_u6_n92, u2_u13_u6_n93, u2_u13_u6_n94, 
       u2_u13_u6_n95, u2_u13_u6_n96, u2_u13_u6_n97, u2_u13_u6_n98, u2_u13_u6_n99, u2_u13_u7_n100, u2_u13_u7_n101, u2_u13_u7_n102, u2_u13_u7_n103, 
       u2_u13_u7_n104, u2_u13_u7_n105, u2_u13_u7_n106, u2_u13_u7_n107, u2_u13_u7_n108, u2_u13_u7_n109, u2_u13_u7_n110, u2_u13_u7_n111, u2_u13_u7_n112, 
       u2_u13_u7_n113, u2_u13_u7_n114, u2_u13_u7_n115, u2_u13_u7_n116, u2_u13_u7_n117, u2_u13_u7_n118, u2_u13_u7_n119, u2_u13_u7_n120, u2_u13_u7_n121, 
       u2_u13_u7_n122, u2_u13_u7_n123, u2_u13_u7_n124, u2_u13_u7_n125, u2_u13_u7_n126, u2_u13_u7_n127, u2_u13_u7_n128, u2_u13_u7_n129, u2_u13_u7_n130, 
       u2_u13_u7_n131, u2_u13_u7_n132, u2_u13_u7_n133, u2_u13_u7_n134, u2_u13_u7_n135, u2_u13_u7_n136, u2_u13_u7_n137, u2_u13_u7_n138, u2_u13_u7_n139, 
       u2_u13_u7_n140, u2_u13_u7_n141, u2_u13_u7_n142, u2_u13_u7_n143, u2_u13_u7_n144, u2_u13_u7_n145, u2_u13_u7_n146, u2_u13_u7_n147, u2_u13_u7_n148, 
       u2_u13_u7_n149, u2_u13_u7_n150, u2_u13_u7_n151, u2_u13_u7_n152, u2_u13_u7_n153, u2_u13_u7_n154, u2_u13_u7_n155, u2_u13_u7_n156, u2_u13_u7_n157, 
       u2_u13_u7_n158, u2_u13_u7_n159, u2_u13_u7_n160, u2_u13_u7_n161, u2_u13_u7_n162, u2_u13_u7_n163, u2_u13_u7_n164, u2_u13_u7_n165, u2_u13_u7_n166, 
       u2_u13_u7_n167, u2_u13_u7_n168, u2_u13_u7_n169, u2_u13_u7_n170, u2_u13_u7_n171, u2_u13_u7_n172, u2_u13_u7_n173, u2_u13_u7_n174, u2_u13_u7_n175, 
       u2_u13_u7_n176, u2_u13_u7_n177, u2_u13_u7_n178, u2_u13_u7_n179, u2_u13_u7_n180, u2_u13_u7_n91, u2_u13_u7_n92, u2_u13_u7_n93, u2_u13_u7_n94, 
       u2_u13_u7_n95, u2_u13_u7_n96, u2_u13_u7_n97, u2_u13_u7_n98, u2_u13_u7_n99, u2_u1_X_31, u2_u1_X_32, u2_u1_X_33, u2_u1_X_34, 
       u2_u1_X_35, u2_u1_X_36, u2_u1_u5_n100, u2_u1_u5_n101, u2_u1_u5_n102, u2_u1_u5_n103, u2_u1_u5_n104, u2_u1_u5_n105, u2_u1_u5_n106, 
       u2_u1_u5_n107, u2_u1_u5_n108, u2_u1_u5_n109, u2_u1_u5_n110, u2_u1_u5_n111, u2_u1_u5_n112, u2_u1_u5_n113, u2_u1_u5_n114, u2_u1_u5_n115, 
       u2_u1_u5_n116, u2_u1_u5_n117, u2_u1_u5_n118, u2_u1_u5_n119, u2_u1_u5_n120, u2_u1_u5_n121, u2_u1_u5_n122, u2_u1_u5_n123, u2_u1_u5_n124, 
       u2_u1_u5_n125, u2_u1_u5_n126, u2_u1_u5_n127, u2_u1_u5_n128, u2_u1_u5_n129, u2_u1_u5_n130, u2_u1_u5_n131, u2_u1_u5_n132, u2_u1_u5_n133, 
       u2_u1_u5_n134, u2_u1_u5_n135, u2_u1_u5_n136, u2_u1_u5_n137, u2_u1_u5_n138, u2_u1_u5_n139, u2_u1_u5_n140, u2_u1_u5_n141, u2_u1_u5_n142, 
       u2_u1_u5_n143, u2_u1_u5_n144, u2_u1_u5_n145, u2_u1_u5_n146, u2_u1_u5_n147, u2_u1_u5_n148, u2_u1_u5_n149, u2_u1_u5_n150, u2_u1_u5_n151, 
       u2_u1_u5_n152, u2_u1_u5_n153, u2_u1_u5_n154, u2_u1_u5_n155, u2_u1_u5_n156, u2_u1_u5_n157, u2_u1_u5_n158, u2_u1_u5_n159, u2_u1_u5_n160, 
       u2_u1_u5_n161, u2_u1_u5_n162, u2_u1_u5_n163, u2_u1_u5_n164, u2_u1_u5_n165, u2_u1_u5_n166, u2_u1_u5_n167, u2_u1_u5_n168, u2_u1_u5_n169, 
       u2_u1_u5_n170, u2_u1_u5_n171, u2_u1_u5_n172, u2_u1_u5_n173, u2_u1_u5_n174, u2_u1_u5_n175, u2_u1_u5_n176, u2_u1_u5_n177, u2_u1_u5_n178, 
       u2_u1_u5_n179, u2_u1_u5_n180, u2_u1_u5_n181, u2_u1_u5_n182, u2_u1_u5_n183, u2_u1_u5_n184, u2_u1_u5_n185, u2_u1_u5_n186, u2_u1_u5_n187, 
       u2_u1_u5_n188, u2_u1_u5_n189, u2_u1_u5_n190, u2_u1_u5_n191, u2_u1_u5_n192, u2_u1_u5_n193, u2_u1_u5_n194, u2_u1_u5_n195, u2_u1_u5_n196, 
       u2_u1_u5_n99, u2_uk_n1000, u2_uk_n312, u2_uk_n338, u2_uk_n342, u2_uk_n349, u2_uk_n353, u2_uk_n369, u2_uk_n391, 
       u2_uk_n407, u2_uk_n676, u2_uk_n685, u2_uk_n686, u2_uk_n717, u2_uk_n930, u2_uk_n932,  u2_uk_n999;
  XOR2_X1 u0_U204 (.B( u0_L9_30 ) , .Z( u0_N349 ) , .A( u0_out10_30 ) );
  XOR2_X1 u0_U208 (.B( u0_L9_26 ) , .Z( u0_N345 ) , .A( u0_out10_26 ) );
  XOR2_X1 u0_U210 (.B( u0_L9_24 ) , .Z( u0_N343 ) , .A( u0_out10_24 ) );
  XOR2_X1 u0_U215 (.B( u0_L9_20 ) , .Z( u0_N339 ) , .A( u0_out10_20 ) );
  XOR2_X1 u0_U219 (.B( u0_L9_16 ) , .Z( u0_N335 ) , .A( u0_out10_16 ) );
  XOR2_X1 u0_U226 (.B( u0_L9_10 ) , .Z( u0_N329 ) , .A( u0_out10_10 ) );
  XOR2_X1 u0_U230 (.B( u0_L9_6 ) , .Z( u0_N325 ) , .A( u0_out10_6 ) );
  XOR2_X1 u0_U235 (.B( u0_L9_1 ) , .Z( u0_N320 ) , .A( u0_out10_1 ) );
  XOR2_X1 u0_U422 (.B( u0_L3_25 ) , .Z( u0_N152 ) , .A( u0_out4_25 ) );
  XOR2_X1 u0_U434 (.B( u0_L3_14 ) , .Z( u0_N141 ) , .A( u0_out4_14 ) );
  XOR2_X1 u0_U441 (.B( u0_L3_8 ) , .Z( u0_N135 ) , .A( u0_out4_8 ) );
  XOR2_X1 u0_U446 (.B( u0_L3_3 ) , .Z( u0_N130 ) , .A( u0_out4_3 ) );
  XOR2_X1 u0_U451 (.B( u0_L2_31 ) , .Z( u0_N126 ) , .A( u0_out3_31 ) );
  XOR2_X1 u0_U452 (.B( u0_L2_30 ) , .Z( u0_N125 ) , .A( u0_out3_30 ) );
  XOR2_X1 u0_U454 (.B( u0_L2_28 ) , .Z( u0_N123 ) , .A( u0_out3_28 ) );
  XOR2_X1 u0_U456 (.B( u0_L2_26 ) , .Z( u0_N121 ) , .A( u0_out3_26 ) );
  XOR2_X1 u0_U459 (.B( u0_L2_24 ) , .Z( u0_N119 ) , .A( u0_out3_24 ) );
  XOR2_X1 u0_U460 (.B( u0_L2_23 ) , .Z( u0_N118 ) , .A( u0_out3_23 ) );
  XOR2_X1 u0_U463 (.B( u0_L2_20 ) , .Z( u0_N115 ) , .A( u0_out3_20 ) );
  XOR2_X1 u0_U465 (.B( u0_L2_18 ) , .Z( u0_N113 ) , .A( u0_out3_18 ) );
  XOR2_X1 u0_U466 (.B( u0_L2_17 ) , .Z( u0_N112 ) , .A( u0_out3_17 ) );
  XOR2_X1 u0_U467 (.B( u0_L2_16 ) , .Z( u0_N111 ) , .A( u0_out3_16 ) );
  XOR2_X1 u0_U471 (.B( u0_L2_13 ) , .Z( u0_N108 ) , .A( u0_out3_13 ) );
  XOR2_X1 u0_U474 (.B( u0_L2_10 ) , .Z( u0_N105 ) , .A( u0_out3_10 ) );
  XOR2_X1 u0_U475 (.B( u0_L2_9 ) , .Z( u0_N104 ) , .A( u0_out3_9 ) );
  XOR2_X1 u0_U478 (.B( u0_L2_6 ) , .Z( u0_N101 ) , .A( u0_out3_6 ) );
  XOR2_X1 u0_U5 (.B( u0_L2_2 ) , .Z( u0_N97 ) , .A( u0_out3_2 ) );
  XOR2_X1 u0_U6 (.B( u0_L2_1 ) , .Z( u0_N96 ) , .A( u0_out3_1 ) );
  XOR2_X1 u0_U60 (.B( u0_L13_32 ) , .Z( u0_N479 ) , .A( u0_out14_32 ) );
  XOR2_X1 u0_U61 (.B( u0_L13_31 ) , .Z( u0_N478 ) , .A( u0_out14_31 ) );
  XOR2_X1 u0_U65 (.B( u0_L13_27 ) , .Z( u0_N474 ) , .A( u0_out14_27 ) );
  XOR2_X1 u0_U67 (.B( u0_L13_25 ) , .Z( u0_N472 ) , .A( u0_out14_25 ) );
  XOR2_X1 u0_U69 (.B( u0_L13_23 ) , .Z( u0_N470 ) , .A( u0_out14_23 ) );
  XOR2_X1 u0_U71 (.B( u0_L13_22 ) , .Z( u0_N469 ) , .A( u0_out14_22 ) );
  XOR2_X1 u0_U72 (.B( u0_L13_21 ) , .Z( u0_N468 ) , .A( u0_out14_21 ) );
  XOR2_X1 u0_U76 (.B( u0_L13_17 ) , .Z( u0_N464 ) , .A( u0_out14_17 ) );
  XOR2_X1 u0_U78 (.B( u0_L13_15 ) , .Z( u0_N462 ) , .A( u0_out14_15 ) );
  XOR2_X1 u0_U79 (.B( u0_L13_14 ) , .Z( u0_N461 ) , .A( u0_out14_14 ) );
  XOR2_X1 u0_U82 (.B( u0_L13_12 ) , .Z( u0_N459 ) , .A( u0_out14_12 ) );
  XOR2_X1 u0_U85 (.B( u0_L13_9 ) , .Z( u0_N456 ) , .A( u0_out14_9 ) );
  XOR2_X1 u0_U86 (.B( u0_L13_8 ) , .Z( u0_N455 ) , .A( u0_out14_8 ) );
  XOR2_X1 u0_U87 (.B( u0_L13_7 ) , .Z( u0_N454 ) , .A( u0_out14_7 ) );
  XOR2_X1 u0_U89 (.B( u0_L13_5 ) , .Z( u0_N452 ) , .A( u0_out14_5 ) );
  XOR2_X1 u0_U91 (.B( u0_L13_3 ) , .Z( u0_N450 ) , .A( u0_out14_3 ) );
  XOR2_X1 u0_u10_U33 (.B( u0_K11_24 ) , .A( u0_R9_17 ) , .Z( u0_u10_X_24 ) );
  XOR2_X1 u0_u10_U34 (.B( u0_K11_23 ) , .A( u0_R9_16 ) , .Z( u0_u10_X_23 ) );
  XOR2_X1 u0_u10_U35 (.B( u0_K11_22 ) , .A( u0_R9_15 ) , .Z( u0_u10_X_22 ) );
  XOR2_X1 u0_u10_U36 (.B( u0_K11_21 ) , .A( u0_R9_14 ) , .Z( u0_u10_X_21 ) );
  XOR2_X1 u0_u10_U37 (.B( u0_K11_20 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_20 ) );
  XOR2_X1 u0_u10_U39 (.B( u0_K11_19 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_19 ) );
  XOR2_X1 u0_u10_U40 (.B( u0_K11_18 ) , .A( u0_R9_13 ) , .Z( u0_u10_X_18 ) );
  XOR2_X1 u0_u10_U41 (.B( u0_K11_17 ) , .A( u0_R9_12 ) , .Z( u0_u10_X_17 ) );
  XOR2_X1 u0_u10_U42 (.B( u0_K11_16 ) , .A( u0_R9_11 ) , .Z( u0_u10_X_16 ) );
  XOR2_X1 u0_u10_U43 (.B( u0_K11_15 ) , .A( u0_R9_10 ) , .Z( u0_u10_X_15 ) );
  XOR2_X1 u0_u10_U44 (.B( u0_K11_14 ) , .A( u0_R9_9 ) , .Z( u0_u10_X_14 ) );
  XOR2_X1 u0_u10_U45 (.B( u0_K11_13 ) , .A( u0_R9_8 ) , .Z( u0_u10_X_13 ) );
  OAI22_X1 u0_u10_u2_U10 (.ZN( u0_u10_u2_n109 ) , .A2( u0_u10_u2_n113 ) , .B2( u0_u10_u2_n133 ) , .B1( u0_u10_u2_n167 ) , .A1( u0_u10_u2_n168 ) );
  NAND3_X1 u0_u10_u2_U100 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n98 ) );
  OAI22_X1 u0_u10_u2_U11 (.B1( u0_u10_u2_n151 ) , .A2( u0_u10_u2_n152 ) , .A1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n160 ) , .B2( u0_u10_u2_n168 ) );
  NOR3_X1 u0_u10_u2_U12 (.A1( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n151 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U13 (.ZN( u0_u10_u2_n144 ) , .B2( u0_u10_u2_n155 ) , .A( u0_u10_u2_n172 ) , .B1( u0_u10_u2_n185 ) );
  AOI21_X1 u0_u10_u2_U14 (.B2( u0_u10_u2_n143 ) , .ZN( u0_u10_u2_n145 ) , .B1( u0_u10_u2_n152 ) , .A( u0_u10_u2_n171 ) );
  AOI21_X1 u0_u10_u2_U15 (.B2( u0_u10_u2_n120 ) , .B1( u0_u10_u2_n121 ) , .ZN( u0_u10_u2_n126 ) , .A( u0_u10_u2_n167 ) );
  INV_X1 u0_u10_u2_U16 (.A( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n171 ) );
  INV_X1 u0_u10_u2_U17 (.A( u0_u10_u2_n120 ) , .ZN( u0_u10_u2_n188 ) );
  NAND2_X1 u0_u10_u2_U18 (.A2( u0_u10_u2_n122 ) , .ZN( u0_u10_u2_n150 ) , .A1( u0_u10_u2_n152 ) );
  INV_X1 u0_u10_u2_U19 (.A( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U20 (.A( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n173 ) );
  NAND2_X1 u0_u10_u2_U21 (.A1( u0_u10_u2_n132 ) , .A2( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n157 ) );
  INV_X1 u0_u10_u2_U22 (.A( u0_u10_u2_n113 ) , .ZN( u0_u10_u2_n178 ) );
  INV_X1 u0_u10_u2_U23 (.A( u0_u10_u2_n139 ) , .ZN( u0_u10_u2_n175 ) );
  INV_X1 u0_u10_u2_U24 (.A( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n181 ) );
  INV_X1 u0_u10_u2_U25 (.A( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n177 ) );
  INV_X1 u0_u10_u2_U26 (.A( u0_u10_u2_n116 ) , .ZN( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U27 (.A( u0_u10_u2_n131 ) , .ZN( u0_u10_u2_n179 ) );
  INV_X1 u0_u10_u2_U28 (.A( u0_u10_u2_n154 ) , .ZN( u0_u10_u2_n176 ) );
  NAND2_X1 u0_u10_u2_U29 (.A2( u0_u10_u2_n116 ) , .A1( u0_u10_u2_n117 ) , .ZN( u0_u10_u2_n118 ) );
  NOR2_X1 u0_u10_u2_U3 (.ZN( u0_u10_u2_n121 ) , .A2( u0_u10_u2_n177 ) , .A1( u0_u10_u2_n180 ) );
  INV_X1 u0_u10_u2_U30 (.A( u0_u10_u2_n132 ) , .ZN( u0_u10_u2_n182 ) );
  INV_X1 u0_u10_u2_U31 (.A( u0_u10_u2_n158 ) , .ZN( u0_u10_u2_n183 ) );
  OAI21_X1 u0_u10_u2_U32 (.A( u0_u10_u2_n156 ) , .B1( u0_u10_u2_n157 ) , .ZN( u0_u10_u2_n158 ) , .B2( u0_u10_u2_n179 ) );
  NOR2_X1 u0_u10_u2_U33 (.ZN( u0_u10_u2_n156 ) , .A1( u0_u10_u2_n166 ) , .A2( u0_u10_u2_n169 ) );
  NOR2_X1 u0_u10_u2_U34 (.A2( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n140 ) );
  NOR2_X1 u0_u10_u2_U35 (.A2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n153 ) , .A1( u0_u10_u2_n156 ) );
  AOI211_X1 u0_u10_u2_U36 (.ZN( u0_u10_u2_n130 ) , .C1( u0_u10_u2_n138 ) , .C2( u0_u10_u2_n179 ) , .B( u0_u10_u2_n96 ) , .A( u0_u10_u2_n97 ) );
  OAI22_X1 u0_u10_u2_U37 (.B1( u0_u10_u2_n133 ) , .A2( u0_u10_u2_n137 ) , .A1( u0_u10_u2_n152 ) , .B2( u0_u10_u2_n168 ) , .ZN( u0_u10_u2_n97 ) );
  OAI221_X1 u0_u10_u2_U38 (.B1( u0_u10_u2_n113 ) , .C1( u0_u10_u2_n132 ) , .A( u0_u10_u2_n149 ) , .B2( u0_u10_u2_n171 ) , .C2( u0_u10_u2_n172 ) , .ZN( u0_u10_u2_n96 ) );
  OAI221_X1 u0_u10_u2_U39 (.A( u0_u10_u2_n115 ) , .C2( u0_u10_u2_n123 ) , .B2( u0_u10_u2_n143 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n163 ) , .C1( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U4 (.A( u0_u10_u2_n134 ) , .ZN( u0_u10_u2_n185 ) );
  OAI21_X1 u0_u10_u2_U40 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n115 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n178 ) );
  OAI221_X1 u0_u10_u2_U41 (.A( u0_u10_u2_n135 ) , .B2( u0_u10_u2_n136 ) , .B1( u0_u10_u2_n137 ) , .ZN( u0_u10_u2_n162 ) , .C2( u0_u10_u2_n167 ) , .C1( u0_u10_u2_n185 ) );
  AND3_X1 u0_u10_u2_U42 (.A3( u0_u10_u2_n131 ) , .A2( u0_u10_u2_n132 ) , .A1( u0_u10_u2_n133 ) , .ZN( u0_u10_u2_n136 ) );
  AOI22_X1 u0_u10_u2_U43 (.ZN( u0_u10_u2_n135 ) , .B1( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n156 ) , .B2( u0_u10_u2_n180 ) , .A2( u0_u10_u2_n188 ) );
  AOI21_X1 u0_u10_u2_U44 (.ZN( u0_u10_u2_n149 ) , .B1( u0_u10_u2_n173 ) , .B2( u0_u10_u2_n188 ) , .A( u0_u10_u2_n95 ) );
  AND3_X1 u0_u10_u2_U45 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n156 ) , .ZN( u0_u10_u2_n95 ) );
  OAI21_X1 u0_u10_u2_U46 (.A( u0_u10_u2_n141 ) , .B2( u0_u10_u2_n142 ) , .ZN( u0_u10_u2_n146 ) , .B1( u0_u10_u2_n153 ) );
  OAI21_X1 u0_u10_u2_U47 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n141 ) , .B1( u0_u10_u2_n176 ) , .B2( u0_u10_u2_n177 ) );
  NOR3_X1 u0_u10_u2_U48 (.ZN( u0_u10_u2_n142 ) , .A3( u0_u10_u2_n175 ) , .A2( u0_u10_u2_n178 ) , .A1( u0_u10_u2_n181 ) );
  OAI21_X1 u0_u10_u2_U49 (.A( u0_u10_u2_n101 ) , .B2( u0_u10_u2_n121 ) , .B1( u0_u10_u2_n153 ) , .ZN( u0_u10_u2_n164 ) );
  INV_X1 u0_u10_u2_U5 (.A( u0_u10_u2_n150 ) , .ZN( u0_u10_u2_n184 ) );
  NAND2_X1 u0_u10_u2_U50 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n155 ) );
  NAND2_X1 u0_u10_u2_U51 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n143 ) );
  NAND2_X1 u0_u10_u2_U52 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n152 ) );
  NAND2_X1 u0_u10_u2_U53 (.A1( u0_u10_u2_n100 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n132 ) );
  INV_X1 u0_u10_u2_U54 (.A( u0_u10_u2_n140 ) , .ZN( u0_u10_u2_n168 ) );
  INV_X1 u0_u10_u2_U55 (.A( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n167 ) );
  NAND2_X1 u0_u10_u2_U56 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n113 ) );
  NAND2_X1 u0_u10_u2_U57 (.A1( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n131 ) );
  NAND2_X1 u0_u10_u2_U58 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n107 ) , .ZN( u0_u10_u2_n139 ) );
  NAND2_X1 u0_u10_u2_U59 (.A1( u0_u10_u2_n103 ) , .A2( u0_u10_u2_n105 ) , .ZN( u0_u10_u2_n133 ) );
  NOR4_X1 u0_u10_u2_U6 (.A4( u0_u10_u2_n124 ) , .A3( u0_u10_u2_n125 ) , .A2( u0_u10_u2_n126 ) , .A1( u0_u10_u2_n127 ) , .ZN( u0_u10_u2_n128 ) );
  NAND2_X1 u0_u10_u2_U60 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n103 ) , .ZN( u0_u10_u2_n154 ) );
  NAND2_X1 u0_u10_u2_U61 (.A2( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n104 ) , .ZN( u0_u10_u2_n119 ) );
  NAND2_X1 u0_u10_u2_U62 (.A2( u0_u10_u2_n107 ) , .A1( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n123 ) );
  NAND2_X1 u0_u10_u2_U63 (.A1( u0_u10_u2_n104 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n122 ) );
  INV_X1 u0_u10_u2_U64 (.A( u0_u10_u2_n114 ) , .ZN( u0_u10_u2_n172 ) );
  NAND2_X1 u0_u10_u2_U65 (.A2( u0_u10_u2_n100 ) , .A1( u0_u10_u2_n102 ) , .ZN( u0_u10_u2_n116 ) );
  NAND2_X1 u0_u10_u2_U66 (.A1( u0_u10_u2_n102 ) , .A2( u0_u10_u2_n108 ) , .ZN( u0_u10_u2_n120 ) );
  NAND2_X1 u0_u10_u2_U67 (.A2( u0_u10_u2_n105 ) , .A1( u0_u10_u2_n106 ) , .ZN( u0_u10_u2_n117 ) );
  INV_X1 u0_u10_u2_U68 (.ZN( u0_u10_u2_n187 ) , .A( u0_u10_u2_n99 ) );
  OAI21_X1 u0_u10_u2_U69 (.B1( u0_u10_u2_n137 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n98 ) , .ZN( u0_u10_u2_n99 ) );
  AOI21_X1 u0_u10_u2_U7 (.ZN( u0_u10_u2_n124 ) , .B1( u0_u10_u2_n131 ) , .B2( u0_u10_u2_n143 ) , .A( u0_u10_u2_n172 ) );
  NOR2_X1 u0_u10_u2_U70 (.A2( u0_u10_X_16 ) , .ZN( u0_u10_u2_n140 ) , .A1( u0_u10_u2_n166 ) );
  NOR2_X1 u0_u10_u2_U71 (.A2( u0_u10_X_13 ) , .A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n100 ) );
  NOR2_X1 u0_u10_u2_U72 (.A2( u0_u10_X_16 ) , .A1( u0_u10_X_17 ) , .ZN( u0_u10_u2_n138 ) );
  NOR2_X1 u0_u10_u2_U73 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n104 ) );
  NOR2_X1 u0_u10_u2_U74 (.A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n103 ) , .A1( u0_u10_u2_n174 ) );
  NOR2_X1 u0_u10_u2_U75 (.A2( u0_u10_X_15 ) , .ZN( u0_u10_u2_n102 ) , .A1( u0_u10_u2_n165 ) );
  NOR2_X1 u0_u10_u2_U76 (.A2( u0_u10_X_17 ) , .ZN( u0_u10_u2_n114 ) , .A1( u0_u10_u2_n169 ) );
  AND2_X1 u0_u10_u2_U77 (.A1( u0_u10_X_15 ) , .ZN( u0_u10_u2_n105 ) , .A2( u0_u10_u2_n165 ) );
  AND2_X1 u0_u10_u2_U78 (.A2( u0_u10_X_15 ) , .A1( u0_u10_X_18 ) , .ZN( u0_u10_u2_n107 ) );
  AND2_X1 u0_u10_u2_U79 (.A1( u0_u10_X_14 ) , .ZN( u0_u10_u2_n106 ) , .A2( u0_u10_u2_n174 ) );
  AOI21_X1 u0_u10_u2_U8 (.B2( u0_u10_u2_n119 ) , .ZN( u0_u10_u2_n127 ) , .A( u0_u10_u2_n137 ) , .B1( u0_u10_u2_n155 ) );
  AND2_X1 u0_u10_u2_U80 (.A1( u0_u10_X_13 ) , .A2( u0_u10_X_14 ) , .ZN( u0_u10_u2_n108 ) );
  INV_X1 u0_u10_u2_U81 (.A( u0_u10_X_16 ) , .ZN( u0_u10_u2_n169 ) );
  INV_X1 u0_u10_u2_U82 (.A( u0_u10_X_17 ) , .ZN( u0_u10_u2_n166 ) );
  INV_X1 u0_u10_u2_U83 (.A( u0_u10_X_13 ) , .ZN( u0_u10_u2_n174 ) );
  INV_X1 u0_u10_u2_U84 (.A( u0_u10_X_18 ) , .ZN( u0_u10_u2_n165 ) );
  NAND4_X1 u0_u10_u2_U85 (.ZN( u0_out10_30 ) , .A4( u0_u10_u2_n147 ) , .A3( u0_u10_u2_n148 ) , .A2( u0_u10_u2_n149 ) , .A1( u0_u10_u2_n187 ) );
  NOR3_X1 u0_u10_u2_U86 (.A3( u0_u10_u2_n144 ) , .A2( u0_u10_u2_n145 ) , .A1( u0_u10_u2_n146 ) , .ZN( u0_u10_u2_n147 ) );
  AOI21_X1 u0_u10_u2_U87 (.B2( u0_u10_u2_n138 ) , .ZN( u0_u10_u2_n148 ) , .A( u0_u10_u2_n162 ) , .B1( u0_u10_u2_n182 ) );
  NAND4_X1 u0_u10_u2_U88 (.ZN( u0_out10_24 ) , .A4( u0_u10_u2_n111 ) , .A3( u0_u10_u2_n112 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n187 ) );
  AOI221_X1 u0_u10_u2_U89 (.A( u0_u10_u2_n109 ) , .B1( u0_u10_u2_n110 ) , .ZN( u0_u10_u2_n111 ) , .C1( u0_u10_u2_n134 ) , .C2( u0_u10_u2_n170 ) , .B2( u0_u10_u2_n173 ) );
  AOI21_X1 u0_u10_u2_U9 (.B2( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n125 ) , .A( u0_u10_u2_n171 ) , .B1( u0_u10_u2_n184 ) );
  AOI21_X1 u0_u10_u2_U90 (.ZN( u0_u10_u2_n112 ) , .B2( u0_u10_u2_n156 ) , .A( u0_u10_u2_n164 ) , .B1( u0_u10_u2_n181 ) );
  NAND4_X1 u0_u10_u2_U91 (.ZN( u0_out10_16 ) , .A4( u0_u10_u2_n128 ) , .A3( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n130 ) , .A2( u0_u10_u2_n186 ) );
  AOI22_X1 u0_u10_u2_U92 (.A2( u0_u10_u2_n118 ) , .ZN( u0_u10_u2_n129 ) , .A1( u0_u10_u2_n140 ) , .B1( u0_u10_u2_n157 ) , .B2( u0_u10_u2_n170 ) );
  INV_X1 u0_u10_u2_U93 (.A( u0_u10_u2_n163 ) , .ZN( u0_u10_u2_n186 ) );
  OR4_X1 u0_u10_u2_U94 (.ZN( u0_out10_6 ) , .A4( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n162 ) , .A2( u0_u10_u2_n163 ) , .A1( u0_u10_u2_n164 ) );
  OR3_X1 u0_u10_u2_U95 (.A2( u0_u10_u2_n159 ) , .A1( u0_u10_u2_n160 ) , .ZN( u0_u10_u2_n161 ) , .A3( u0_u10_u2_n183 ) );
  AOI21_X1 u0_u10_u2_U96 (.B2( u0_u10_u2_n154 ) , .B1( u0_u10_u2_n155 ) , .ZN( u0_u10_u2_n159 ) , .A( u0_u10_u2_n167 ) );
  NAND3_X1 u0_u10_u2_U97 (.A2( u0_u10_u2_n117 ) , .A1( u0_u10_u2_n122 ) , .A3( u0_u10_u2_n123 ) , .ZN( u0_u10_u2_n134 ) );
  NAND3_X1 u0_u10_u2_U98 (.ZN( u0_u10_u2_n110 ) , .A2( u0_u10_u2_n131 ) , .A3( u0_u10_u2_n139 ) , .A1( u0_u10_u2_n154 ) );
  NAND3_X1 u0_u10_u2_U99 (.A2( u0_u10_u2_n100 ) , .ZN( u0_u10_u2_n101 ) , .A1( u0_u10_u2_n104 ) , .A3( u0_u10_u2_n114 ) );
  OAI22_X1 u0_u10_u3_U10 (.B1( u0_u10_u3_n113 ) , .A2( u0_u10_u3_n135 ) , .A1( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n164 ) , .ZN( u0_u10_u3_n98 ) );
  OAI211_X1 u0_u10_u3_U11 (.B( u0_u10_u3_n106 ) , .ZN( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n128 ) , .C1( u0_u10_u3_n167 ) , .A( u0_u10_u3_n181 ) );
  AOI221_X1 u0_u10_u3_U12 (.C1( u0_u10_u3_n105 ) , .ZN( u0_u10_u3_n106 ) , .A( u0_u10_u3_n131 ) , .B2( u0_u10_u3_n132 ) , .C2( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n169 ) );
  INV_X1 u0_u10_u3_U13 (.ZN( u0_u10_u3_n181 ) , .A( u0_u10_u3_n98 ) );
  NAND2_X1 u0_u10_u3_U14 (.ZN( u0_u10_u3_n105 ) , .A2( u0_u10_u3_n130 ) , .A1( u0_u10_u3_n155 ) );
  AOI22_X1 u0_u10_u3_U15 (.B1( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n116 ) , .ZN( u0_u10_u3_n123 ) , .B2( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U16 (.ZN( u0_u10_u3_n116 ) , .A2( u0_u10_u3_n151 ) , .A1( u0_u10_u3_n182 ) );
  NOR2_X1 u0_u10_u3_U17 (.ZN( u0_u10_u3_n126 ) , .A2( u0_u10_u3_n150 ) , .A1( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U18 (.ZN( u0_u10_u3_n112 ) , .B2( u0_u10_u3_n146 ) , .B1( u0_u10_u3_n155 ) , .A( u0_u10_u3_n167 ) );
  NAND2_X1 u0_u10_u3_U19 (.A1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n142 ) , .A2( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U20 (.ZN( u0_u10_u3_n132 ) , .A2( u0_u10_u3_n152 ) , .A1( u0_u10_u3_n156 ) );
  AND2_X1 u0_u10_u3_U21 (.A2( u0_u10_u3_n113 ) , .A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n151 ) );
  INV_X1 u0_u10_u3_U22 (.A( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n165 ) );
  INV_X1 u0_u10_u3_U23 (.A( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n170 ) );
  NAND2_X1 u0_u10_u3_U24 (.A1( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .ZN( u0_u10_u3_n140 ) );
  NAND2_X1 u0_u10_u3_U25 (.ZN( u0_u10_u3_n117 ) , .A1( u0_u10_u3_n124 ) , .A2( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U26 (.ZN( u0_u10_u3_n143 ) , .A1( u0_u10_u3_n165 ) , .A2( u0_u10_u3_n167 ) );
  INV_X1 u0_u10_u3_U27 (.A( u0_u10_u3_n130 ) , .ZN( u0_u10_u3_n177 ) );
  INV_X1 u0_u10_u3_U28 (.A( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n176 ) );
  INV_X1 u0_u10_u3_U29 (.A( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n174 ) );
  INV_X1 u0_u10_u3_U3 (.A( u0_u10_u3_n129 ) , .ZN( u0_u10_u3_n183 ) );
  INV_X1 u0_u10_u3_U30 (.A( u0_u10_u3_n139 ) , .ZN( u0_u10_u3_n185 ) );
  NOR2_X1 u0_u10_u3_U31 (.ZN( u0_u10_u3_n135 ) , .A2( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n169 ) );
  OAI222_X1 u0_u10_u3_U32 (.C2( u0_u10_u3_n107 ) , .A2( u0_u10_u3_n108 ) , .B1( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n138 ) , .B2( u0_u10_u3_n146 ) , .C1( u0_u10_u3_n154 ) , .A1( u0_u10_u3_n164 ) );
  NOR4_X1 u0_u10_u3_U33 (.A4( u0_u10_u3_n157 ) , .A3( u0_u10_u3_n158 ) , .A2( u0_u10_u3_n159 ) , .A1( u0_u10_u3_n160 ) , .ZN( u0_u10_u3_n161 ) );
  AOI21_X1 u0_u10_u3_U34 (.B2( u0_u10_u3_n152 ) , .B1( u0_u10_u3_n153 ) , .ZN( u0_u10_u3_n158 ) , .A( u0_u10_u3_n164 ) );
  AOI21_X1 u0_u10_u3_U35 (.A( u0_u10_u3_n154 ) , .B2( u0_u10_u3_n155 ) , .B1( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n157 ) );
  AOI21_X1 u0_u10_u3_U36 (.A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n150 ) , .B1( u0_u10_u3_n151 ) , .ZN( u0_u10_u3_n159 ) );
  AOI211_X1 u0_u10_u3_U37 (.ZN( u0_u10_u3_n109 ) , .A( u0_u10_u3_n119 ) , .C2( u0_u10_u3_n129 ) , .B( u0_u10_u3_n138 ) , .C1( u0_u10_u3_n141 ) );
  AOI211_X1 u0_u10_u3_U38 (.B( u0_u10_u3_n119 ) , .A( u0_u10_u3_n120 ) , .C2( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n122 ) , .C1( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U39 (.A( u0_u10_u3_n156 ) , .ZN( u0_u10_u3_n179 ) );
  INV_X1 u0_u10_u3_U4 (.A( u0_u10_u3_n140 ) , .ZN( u0_u10_u3_n182 ) );
  OAI22_X1 u0_u10_u3_U40 (.B1( u0_u10_u3_n118 ) , .ZN( u0_u10_u3_n120 ) , .A1( u0_u10_u3_n135 ) , .B2( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n178 ) );
  AND3_X1 u0_u10_u3_U41 (.ZN( u0_u10_u3_n118 ) , .A2( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n144 ) , .A3( u0_u10_u3_n152 ) );
  INV_X1 u0_u10_u3_U42 (.A( u0_u10_u3_n121 ) , .ZN( u0_u10_u3_n164 ) );
  NAND2_X1 u0_u10_u3_U43 (.ZN( u0_u10_u3_n133 ) , .A1( u0_u10_u3_n154 ) , .A2( u0_u10_u3_n164 ) );
  OAI211_X1 u0_u10_u3_U44 (.B( u0_u10_u3_n127 ) , .ZN( u0_u10_u3_n139 ) , .C1( u0_u10_u3_n150 ) , .C2( u0_u10_u3_n154 ) , .A( u0_u10_u3_n184 ) );
  INV_X1 u0_u10_u3_U45 (.A( u0_u10_u3_n125 ) , .ZN( u0_u10_u3_n184 ) );
  AOI221_X1 u0_u10_u3_U46 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n127 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n169 ) , .B2( u0_u10_u3_n170 ) , .B1( u0_u10_u3_n174 ) );
  OAI22_X1 u0_u10_u3_U47 (.A1( u0_u10_u3_n124 ) , .ZN( u0_u10_u3_n125 ) , .B2( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n165 ) , .B1( u0_u10_u3_n167 ) );
  NOR2_X1 u0_u10_u3_U48 (.A1( u0_u10_u3_n113 ) , .ZN( u0_u10_u3_n131 ) , .A2( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U49 (.A1( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n150 ) , .A2( u0_u10_u3_n99 ) );
  INV_X1 u0_u10_u3_U5 (.A( u0_u10_u3_n117 ) , .ZN( u0_u10_u3_n178 ) );
  NAND2_X1 u0_u10_u3_U50 (.A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n155 ) , .A1( u0_u10_u3_n97 ) );
  INV_X1 u0_u10_u3_U51 (.A( u0_u10_u3_n141 ) , .ZN( u0_u10_u3_n167 ) );
  AOI21_X1 u0_u10_u3_U52 (.B2( u0_u10_u3_n114 ) , .B1( u0_u10_u3_n146 ) , .A( u0_u10_u3_n154 ) , .ZN( u0_u10_u3_n94 ) );
  AOI21_X1 u0_u10_u3_U53 (.ZN( u0_u10_u3_n110 ) , .B2( u0_u10_u3_n142 ) , .B1( u0_u10_u3_n186 ) , .A( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U54 (.A( u0_u10_u3_n145 ) , .ZN( u0_u10_u3_n186 ) );
  AOI21_X1 u0_u10_u3_U55 (.B1( u0_u10_u3_n124 ) , .A( u0_u10_u3_n149 ) , .B2( u0_u10_u3_n155 ) , .ZN( u0_u10_u3_n95 ) );
  INV_X1 u0_u10_u3_U56 (.A( u0_u10_u3_n149 ) , .ZN( u0_u10_u3_n169 ) );
  NAND2_X1 u0_u10_u3_U57 (.ZN( u0_u10_u3_n124 ) , .A1( u0_u10_u3_n96 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U58 (.A2( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n146 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U59 (.A1( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n145 ) , .A2( u0_u10_u3_n99 ) );
  AOI221_X1 u0_u10_u3_U6 (.A( u0_u10_u3_n131 ) , .C2( u0_u10_u3_n132 ) , .C1( u0_u10_u3_n133 ) , .ZN( u0_u10_u3_n134 ) , .B1( u0_u10_u3_n143 ) , .B2( u0_u10_u3_n177 ) );
  NAND2_X1 u0_u10_u3_U60 (.A1( u0_u10_u3_n100 ) , .ZN( u0_u10_u3_n156 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U61 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n148 ) );
  NAND2_X1 u0_u10_u3_U62 (.A1( u0_u10_u3_n100 ) , .A2( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n128 ) );
  NAND2_X1 u0_u10_u3_U63 (.A2( u0_u10_u3_n101 ) , .A1( u0_u10_u3_n102 ) , .ZN( u0_u10_u3_n152 ) );
  NAND2_X1 u0_u10_u3_U64 (.A2( u0_u10_u3_n101 ) , .ZN( u0_u10_u3_n114 ) , .A1( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U65 (.ZN( u0_u10_u3_n107 ) , .A1( u0_u10_u3_n97 ) , .A2( u0_u10_u3_n99 ) );
  NAND2_X1 u0_u10_u3_U66 (.A2( u0_u10_u3_n100 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n113 ) );
  NAND2_X1 u0_u10_u3_U67 (.A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n153 ) , .A2( u0_u10_u3_n97 ) );
  NAND2_X1 u0_u10_u3_U68 (.A2( u0_u10_u3_n103 ) , .A1( u0_u10_u3_n104 ) , .ZN( u0_u10_u3_n130 ) );
  NAND2_X1 u0_u10_u3_U69 (.A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n96 ) );
  OAI22_X1 u0_u10_u3_U7 (.B2( u0_u10_u3_n147 ) , .A2( u0_u10_u3_n148 ) , .ZN( u0_u10_u3_n160 ) , .B1( u0_u10_u3_n165 ) , .A1( u0_u10_u3_n168 ) );
  NAND2_X1 u0_u10_u3_U70 (.A1( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n103 ) , .ZN( u0_u10_u3_n108 ) );
  NOR2_X1 u0_u10_u3_U71 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n99 ) );
  NOR2_X1 u0_u10_u3_U72 (.A2( u0_u10_X_21 ) , .A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n103 ) );
  NOR2_X1 u0_u10_u3_U73 (.A2( u0_u10_X_24 ) , .A1( u0_u10_u3_n171 ) , .ZN( u0_u10_u3_n97 ) );
  NOR2_X1 u0_u10_u3_U74 (.A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n141 ) , .A1( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U75 (.A2( u0_u10_X_19 ) , .A1( u0_u10_u3_n172 ) , .ZN( u0_u10_u3_n96 ) );
  NAND2_X1 u0_u10_u3_U76 (.A1( u0_u10_X_22 ) , .A2( u0_u10_X_23 ) , .ZN( u0_u10_u3_n154 ) );
  NAND2_X1 u0_u10_u3_U77 (.A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n149 ) , .A2( u0_u10_u3_n166 ) );
  NOR2_X1 u0_u10_u3_U78 (.A2( u0_u10_X_22 ) , .A1( u0_u10_X_23 ) , .ZN( u0_u10_u3_n121 ) );
  AND2_X1 u0_u10_u3_U79 (.A1( u0_u10_X_24 ) , .ZN( u0_u10_u3_n101 ) , .A2( u0_u10_u3_n171 ) );
  AND3_X1 u0_u10_u3_U8 (.A3( u0_u10_u3_n144 ) , .A2( u0_u10_u3_n145 ) , .A1( u0_u10_u3_n146 ) , .ZN( u0_u10_u3_n147 ) );
  AND2_X1 u0_u10_u3_U80 (.A1( u0_u10_X_19 ) , .ZN( u0_u10_u3_n102 ) , .A2( u0_u10_u3_n172 ) );
  AND2_X1 u0_u10_u3_U81 (.A1( u0_u10_X_21 ) , .A2( u0_u10_X_24 ) , .ZN( u0_u10_u3_n100 ) );
  AND2_X1 u0_u10_u3_U82 (.A2( u0_u10_X_19 ) , .A1( u0_u10_X_20 ) , .ZN( u0_u10_u3_n104 ) );
  INV_X1 u0_u10_u3_U83 (.A( u0_u10_X_22 ) , .ZN( u0_u10_u3_n166 ) );
  INV_X1 u0_u10_u3_U84 (.A( u0_u10_X_21 ) , .ZN( u0_u10_u3_n171 ) );
  INV_X1 u0_u10_u3_U85 (.A( u0_u10_X_20 ) , .ZN( u0_u10_u3_n172 ) );
  OR4_X1 u0_u10_u3_U86 (.ZN( u0_out10_10 ) , .A4( u0_u10_u3_n136 ) , .A3( u0_u10_u3_n137 ) , .A1( u0_u10_u3_n138 ) , .A2( u0_u10_u3_n139 ) );
  OAI222_X1 u0_u10_u3_U87 (.C1( u0_u10_u3_n128 ) , .ZN( u0_u10_u3_n137 ) , .B1( u0_u10_u3_n148 ) , .A2( u0_u10_u3_n150 ) , .B2( u0_u10_u3_n154 ) , .C2( u0_u10_u3_n164 ) , .A1( u0_u10_u3_n167 ) );
  OAI221_X1 u0_u10_u3_U88 (.A( u0_u10_u3_n134 ) , .B2( u0_u10_u3_n135 ) , .ZN( u0_u10_u3_n136 ) , .C1( u0_u10_u3_n149 ) , .B1( u0_u10_u3_n151 ) , .C2( u0_u10_u3_n183 ) );
  NAND4_X1 u0_u10_u3_U89 (.ZN( u0_out10_26 ) , .A4( u0_u10_u3_n109 ) , .A3( u0_u10_u3_n110 ) , .A2( u0_u10_u3_n111 ) , .A1( u0_u10_u3_n173 ) );
  INV_X1 u0_u10_u3_U9 (.A( u0_u10_u3_n143 ) , .ZN( u0_u10_u3_n168 ) );
  INV_X1 u0_u10_u3_U90 (.ZN( u0_u10_u3_n173 ) , .A( u0_u10_u3_n94 ) );
  OAI21_X1 u0_u10_u3_U91 (.ZN( u0_u10_u3_n111 ) , .B2( u0_u10_u3_n117 ) , .A( u0_u10_u3_n133 ) , .B1( u0_u10_u3_n176 ) );
  NAND4_X1 u0_u10_u3_U92 (.ZN( u0_out10_20 ) , .A4( u0_u10_u3_n122 ) , .A3( u0_u10_u3_n123 ) , .A1( u0_u10_u3_n175 ) , .A2( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U93 (.A( u0_u10_u3_n126 ) , .ZN( u0_u10_u3_n180 ) );
  INV_X1 u0_u10_u3_U94 (.A( u0_u10_u3_n112 ) , .ZN( u0_u10_u3_n175 ) );
  NAND4_X1 u0_u10_u3_U95 (.ZN( u0_out10_1 ) , .A4( u0_u10_u3_n161 ) , .A3( u0_u10_u3_n162 ) , .A2( u0_u10_u3_n163 ) , .A1( u0_u10_u3_n185 ) );
  NAND2_X1 u0_u10_u3_U96 (.ZN( u0_u10_u3_n163 ) , .A2( u0_u10_u3_n170 ) , .A1( u0_u10_u3_n176 ) );
  AOI22_X1 u0_u10_u3_U97 (.B2( u0_u10_u3_n140 ) , .B1( u0_u10_u3_n141 ) , .A2( u0_u10_u3_n142 ) , .ZN( u0_u10_u3_n162 ) , .A1( u0_u10_u3_n177 ) );
  NAND3_X1 u0_u10_u3_U98 (.A1( u0_u10_u3_n114 ) , .ZN( u0_u10_u3_n115 ) , .A2( u0_u10_u3_n145 ) , .A3( u0_u10_u3_n153 ) );
  NAND3_X1 u0_u10_u3_U99 (.ZN( u0_u10_u3_n129 ) , .A2( u0_u10_u3_n144 ) , .A1( u0_u10_u3_n153 ) , .A3( u0_u10_u3_n182 ) );
  XOR2_X1 u0_u14_U10 (.B( u0_K15_45 ) , .A( u0_R13_30 ) , .Z( u0_u14_X_45 ) );
  XOR2_X1 u0_u14_U11 (.B( u0_K15_44 ) , .A( u0_R13_29 ) , .Z( u0_u14_X_44 ) );
  XOR2_X1 u0_u14_U12 (.B( u0_K15_43 ) , .A( u0_R13_28 ) , .Z( u0_u14_X_43 ) );
  XOR2_X1 u0_u14_U13 (.B( u0_K15_42 ) , .A( u0_R13_29 ) , .Z( u0_u14_X_42 ) );
  XOR2_X1 u0_u14_U14 (.B( u0_K15_41 ) , .A( u0_R13_28 ) , .Z( u0_u14_X_41 ) );
  XOR2_X1 u0_u14_U15 (.B( u0_K15_40 ) , .A( u0_R13_27 ) , .Z( u0_u14_X_40 ) );
  XOR2_X1 u0_u14_U16 (.B( u0_K15_3 ) , .A( u0_R13_2 ) , .Z( u0_u14_X_3 ) );
  XOR2_X1 u0_u14_U17 (.B( u0_K15_39 ) , .A( u0_R13_26 ) , .Z( u0_u14_X_39 ) );
  XOR2_X1 u0_u14_U18 (.B( u0_K15_38 ) , .A( u0_R13_25 ) , .Z( u0_u14_X_38 ) );
  XOR2_X1 u0_u14_U19 (.B( u0_K15_37 ) , .A( u0_R13_24 ) , .Z( u0_u14_X_37 ) );
  XOR2_X1 u0_u14_U26 (.B( u0_K15_30 ) , .A( u0_R13_21 ) , .Z( u0_u14_X_30 ) );
  XOR2_X1 u0_u14_U27 (.B( u0_K15_2 ) , .A( u0_R13_1 ) , .Z( u0_u14_X_2 ) );
  XOR2_X1 u0_u14_U28 (.B( u0_K15_29 ) , .A( u0_R13_20 ) , .Z( u0_u14_X_29 ) );
  XOR2_X1 u0_u14_U29 (.B( u0_K15_28 ) , .A( u0_R13_19 ) , .Z( u0_u14_X_28 ) );
  XOR2_X1 u0_u14_U30 (.B( u0_K15_27 ) , .A( u0_R13_18 ) , .Z( u0_u14_X_27 ) );
  XOR2_X1 u0_u14_U31 (.B( u0_K15_26 ) , .A( u0_R13_17 ) , .Z( u0_u14_X_26 ) );
  XOR2_X1 u0_u14_U32 (.B( u0_K15_25 ) , .A( u0_R13_16 ) , .Z( u0_u14_X_25 ) );
  XOR2_X1 u0_u14_U38 (.B( u0_K15_1 ) , .A( u0_R13_32 ) , .Z( u0_u14_X_1 ) );
  XOR2_X1 u0_u14_U4 (.B( u0_K15_6 ) , .A( u0_R13_5 ) , .Z( u0_u14_X_6 ) );
  XOR2_X1 u0_u14_U5 (.B( u0_K15_5 ) , .A( u0_R13_4 ) , .Z( u0_u14_X_5 ) );
  XOR2_X1 u0_u14_U6 (.B( u0_K15_4 ) , .A( u0_R13_3 ) , .Z( u0_u14_X_4 ) );
  XOR2_X1 u0_u14_U7 (.B( u0_K15_48 ) , .A( u0_R13_1 ) , .Z( u0_u14_X_48 ) );
  XOR2_X1 u0_u14_U8 (.B( u0_K15_47 ) , .A( u0_R13_32 ) , .Z( u0_u14_X_47 ) );
  XOR2_X1 u0_u14_U9 (.B( u0_K15_46 ) , .A( u0_R13_31 ) , .Z( u0_u14_X_46 ) );
  AND3_X1 u0_u14_u0_U10 (.A2( u0_u14_u0_n112 ) , .ZN( u0_u14_u0_n127 ) , .A3( u0_u14_u0_n130 ) , .A1( u0_u14_u0_n148 ) );
  NAND2_X1 u0_u14_u0_U11 (.ZN( u0_u14_u0_n113 ) , .A1( u0_u14_u0_n139 ) , .A2( u0_u14_u0_n149 ) );
  AND2_X1 u0_u14_u0_U12 (.ZN( u0_u14_u0_n107 ) , .A1( u0_u14_u0_n130 ) , .A2( u0_u14_u0_n140 ) );
  AND2_X1 u0_u14_u0_U13 (.A2( u0_u14_u0_n129 ) , .A1( u0_u14_u0_n130 ) , .ZN( u0_u14_u0_n151 ) );
  AND2_X1 u0_u14_u0_U14 (.A1( u0_u14_u0_n108 ) , .A2( u0_u14_u0_n125 ) , .ZN( u0_u14_u0_n145 ) );
  INV_X1 u0_u14_u0_U15 (.A( u0_u14_u0_n143 ) , .ZN( u0_u14_u0_n173 ) );
  NOR2_X1 u0_u14_u0_U16 (.A2( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n147 ) , .A1( u0_u14_u0_n160 ) );
  NOR2_X1 u0_u14_u0_U17 (.A1( u0_u14_u0_n163 ) , .A2( u0_u14_u0_n164 ) , .ZN( u0_u14_u0_n95 ) );
  AOI21_X1 u0_u14_u0_U18 (.B1( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n132 ) , .A( u0_u14_u0_n165 ) , .B2( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U19 (.A( u0_u14_u0_n142 ) , .ZN( u0_u14_u0_n165 ) );
  OAI221_X1 u0_u14_u0_U20 (.C1( u0_u14_u0_n121 ) , .ZN( u0_u14_u0_n122 ) , .B2( u0_u14_u0_n127 ) , .A( u0_u14_u0_n143 ) , .B1( u0_u14_u0_n144 ) , .C2( u0_u14_u0_n147 ) );
  OAI22_X1 u0_u14_u0_U21 (.B1( u0_u14_u0_n125 ) , .ZN( u0_u14_u0_n126 ) , .A1( u0_u14_u0_n138 ) , .A2( u0_u14_u0_n146 ) , .B2( u0_u14_u0_n147 ) );
  OAI22_X1 u0_u14_u0_U22 (.B1( u0_u14_u0_n131 ) , .A1( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n147 ) , .A2( u0_u14_u0_n90 ) , .ZN( u0_u14_u0_n91 ) );
  AND3_X1 u0_u14_u0_U23 (.A3( u0_u14_u0_n121 ) , .A2( u0_u14_u0_n125 ) , .A1( u0_u14_u0_n148 ) , .ZN( u0_u14_u0_n90 ) );
  NAND2_X1 u0_u14_u0_U24 (.A1( u0_u14_u0_n100 ) , .A2( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n125 ) );
  INV_X1 u0_u14_u0_U25 (.A( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n161 ) );
  NOR2_X1 u0_u14_u0_U26 (.A1( u0_u14_u0_n120 ) , .ZN( u0_u14_u0_n143 ) , .A2( u0_u14_u0_n167 ) );
  OAI221_X1 u0_u14_u0_U27 (.C1( u0_u14_u0_n112 ) , .ZN( u0_u14_u0_n120 ) , .B1( u0_u14_u0_n138 ) , .B2( u0_u14_u0_n141 ) , .C2( u0_u14_u0_n147 ) , .A( u0_u14_u0_n172 ) );
  AOI211_X1 u0_u14_u0_U28 (.B( u0_u14_u0_n115 ) , .A( u0_u14_u0_n116 ) , .C2( u0_u14_u0_n117 ) , .C1( u0_u14_u0_n118 ) , .ZN( u0_u14_u0_n119 ) );
  AOI22_X1 u0_u14_u0_U29 (.B2( u0_u14_u0_n109 ) , .A2( u0_u14_u0_n110 ) , .ZN( u0_u14_u0_n111 ) , .B1( u0_u14_u0_n118 ) , .A1( u0_u14_u0_n160 ) );
  INV_X1 u0_u14_u0_U3 (.A( u0_u14_u0_n113 ) , .ZN( u0_u14_u0_n166 ) );
  NAND2_X1 u0_u14_u0_U30 (.A1( u0_u14_u0_n100 ) , .ZN( u0_u14_u0_n129 ) , .A2( u0_u14_u0_n95 ) );
  INV_X1 u0_u14_u0_U31 (.A( u0_u14_u0_n118 ) , .ZN( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U32 (.ZN( u0_u14_u0_n104 ) , .B1( u0_u14_u0_n107 ) , .B2( u0_u14_u0_n141 ) , .A( u0_u14_u0_n144 ) );
  AOI21_X1 u0_u14_u0_U33 (.B1( u0_u14_u0_n127 ) , .B2( u0_u14_u0_n129 ) , .A( u0_u14_u0_n138 ) , .ZN( u0_u14_u0_n96 ) );
  AOI21_X1 u0_u14_u0_U34 (.ZN( u0_u14_u0_n116 ) , .B2( u0_u14_u0_n142 ) , .A( u0_u14_u0_n144 ) , .B1( u0_u14_u0_n166 ) );
  NAND2_X1 u0_u14_u0_U35 (.A2( u0_u14_u0_n100 ) , .A1( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n139 ) );
  NAND2_X1 u0_u14_u0_U36 (.A2( u0_u14_u0_n100 ) , .ZN( u0_u14_u0_n131 ) , .A1( u0_u14_u0_n92 ) );
  NAND2_X1 u0_u14_u0_U37 (.A1( u0_u14_u0_n101 ) , .A2( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n150 ) );
  INV_X1 u0_u14_u0_U38 (.A( u0_u14_u0_n138 ) , .ZN( u0_u14_u0_n160 ) );
  NAND2_X1 u0_u14_u0_U39 (.A1( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n128 ) , .A2( u0_u14_u0_n95 ) );
  AOI21_X1 u0_u14_u0_U4 (.B1( u0_u14_u0_n114 ) , .ZN( u0_u14_u0_n115 ) , .B2( u0_u14_u0_n129 ) , .A( u0_u14_u0_n161 ) );
  NAND2_X1 u0_u14_u0_U40 (.ZN( u0_u14_u0_n148 ) , .A1( u0_u14_u0_n93 ) , .A2( u0_u14_u0_n95 ) );
  NAND2_X1 u0_u14_u0_U41 (.A2( u0_u14_u0_n102 ) , .A1( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n149 ) );
  NAND2_X1 u0_u14_u0_U42 (.A2( u0_u14_u0_n102 ) , .ZN( u0_u14_u0_n114 ) , .A1( u0_u14_u0_n92 ) );
  NAND2_X1 u0_u14_u0_U43 (.A2( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n121 ) , .A1( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U44 (.ZN( u0_u14_u0_n172 ) , .A( u0_u14_u0_n88 ) );
  OAI222_X1 u0_u14_u0_U45 (.C1( u0_u14_u0_n108 ) , .A1( u0_u14_u0_n125 ) , .B2( u0_u14_u0_n128 ) , .B1( u0_u14_u0_n144 ) , .A2( u0_u14_u0_n158 ) , .C2( u0_u14_u0_n161 ) , .ZN( u0_u14_u0_n88 ) );
  NAND2_X1 u0_u14_u0_U46 (.ZN( u0_u14_u0_n112 ) , .A2( u0_u14_u0_n92 ) , .A1( u0_u14_u0_n93 ) );
  OR3_X1 u0_u14_u0_U47 (.A3( u0_u14_u0_n152 ) , .A2( u0_u14_u0_n153 ) , .A1( u0_u14_u0_n154 ) , .ZN( u0_u14_u0_n155 ) );
  AOI21_X1 u0_u14_u0_U48 (.B2( u0_u14_u0_n150 ) , .B1( u0_u14_u0_n151 ) , .ZN( u0_u14_u0_n152 ) , .A( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U49 (.A( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n145 ) , .B1( u0_u14_u0_n146 ) , .ZN( u0_u14_u0_n154 ) );
  AOI21_X1 u0_u14_u0_U5 (.B2( u0_u14_u0_n131 ) , .ZN( u0_u14_u0_n134 ) , .B1( u0_u14_u0_n151 ) , .A( u0_u14_u0_n158 ) );
  AOI21_X1 u0_u14_u0_U50 (.A( u0_u14_u0_n147 ) , .B2( u0_u14_u0_n148 ) , .B1( u0_u14_u0_n149 ) , .ZN( u0_u14_u0_n153 ) );
  INV_X1 u0_u14_u0_U51 (.ZN( u0_u14_u0_n171 ) , .A( u0_u14_u0_n99 ) );
  OAI211_X1 u0_u14_u0_U52 (.C2( u0_u14_u0_n140 ) , .C1( u0_u14_u0_n161 ) , .A( u0_u14_u0_n169 ) , .B( u0_u14_u0_n98 ) , .ZN( u0_u14_u0_n99 ) );
  AOI211_X1 u0_u14_u0_U53 (.C1( u0_u14_u0_n118 ) , .A( u0_u14_u0_n123 ) , .B( u0_u14_u0_n96 ) , .C2( u0_u14_u0_n97 ) , .ZN( u0_u14_u0_n98 ) );
  INV_X1 u0_u14_u0_U54 (.ZN( u0_u14_u0_n169 ) , .A( u0_u14_u0_n91 ) );
  NOR2_X1 u0_u14_u0_U55 (.A2( u0_u14_X_4 ) , .A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n118 ) );
  NOR2_X1 u0_u14_u0_U56 (.A2( u0_u14_X_2 ) , .ZN( u0_u14_u0_n103 ) , .A1( u0_u14_u0_n164 ) );
  NOR2_X1 u0_u14_u0_U57 (.A2( u0_u14_X_1 ) , .A1( u0_u14_X_2 ) , .ZN( u0_u14_u0_n92 ) );
  NOR2_X1 u0_u14_u0_U58 (.A2( u0_u14_X_1 ) , .ZN( u0_u14_u0_n101 ) , .A1( u0_u14_u0_n163 ) );
  NAND2_X1 u0_u14_u0_U59 (.A2( u0_u14_X_4 ) , .A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n144 ) );
  NOR2_X1 u0_u14_u0_U6 (.A1( u0_u14_u0_n108 ) , .ZN( u0_u14_u0_n123 ) , .A2( u0_u14_u0_n158 ) );
  NOR2_X1 u0_u14_u0_U60 (.A2( u0_u14_X_5 ) , .ZN( u0_u14_u0_n136 ) , .A1( u0_u14_u0_n159 ) );
  NAND2_X1 u0_u14_u0_U61 (.A1( u0_u14_X_5 ) , .ZN( u0_u14_u0_n138 ) , .A2( u0_u14_u0_n159 ) );
  AND2_X1 u0_u14_u0_U62 (.A2( u0_u14_X_3 ) , .A1( u0_u14_X_6 ) , .ZN( u0_u14_u0_n102 ) );
  AND2_X1 u0_u14_u0_U63 (.A1( u0_u14_X_6 ) , .A2( u0_u14_u0_n162 ) , .ZN( u0_u14_u0_n93 ) );
  INV_X1 u0_u14_u0_U64 (.A( u0_u14_X_4 ) , .ZN( u0_u14_u0_n159 ) );
  INV_X1 u0_u14_u0_U65 (.A( u0_u14_X_1 ) , .ZN( u0_u14_u0_n164 ) );
  INV_X1 u0_u14_u0_U66 (.A( u0_u14_X_2 ) , .ZN( u0_u14_u0_n163 ) );
  INV_X1 u0_u14_u0_U67 (.A( u0_u14_X_3 ) , .ZN( u0_u14_u0_n162 ) );
  INV_X1 u0_u14_u0_U68 (.A( u0_u14_u0_n126 ) , .ZN( u0_u14_u0_n168 ) );
  AOI211_X1 u0_u14_u0_U69 (.B( u0_u14_u0_n133 ) , .A( u0_u14_u0_n134 ) , .C2( u0_u14_u0_n135 ) , .C1( u0_u14_u0_n136 ) , .ZN( u0_u14_u0_n137 ) );
  OAI21_X1 u0_u14_u0_U7 (.B1( u0_u14_u0_n150 ) , .B2( u0_u14_u0_n158 ) , .A( u0_u14_u0_n172 ) , .ZN( u0_u14_u0_n89 ) );
  INV_X1 u0_u14_u0_U70 (.ZN( u0_u14_u0_n174 ) , .A( u0_u14_u0_n89 ) );
  AOI211_X1 u0_u14_u0_U71 (.B( u0_u14_u0_n104 ) , .A( u0_u14_u0_n105 ) , .ZN( u0_u14_u0_n106 ) , .C2( u0_u14_u0_n113 ) , .C1( u0_u14_u0_n160 ) );
  OR4_X1 u0_u14_u0_U72 (.ZN( u0_out14_31 ) , .A4( u0_u14_u0_n155 ) , .A2( u0_u14_u0_n156 ) , .A1( u0_u14_u0_n157 ) , .A3( u0_u14_u0_n173 ) );
  AOI21_X1 u0_u14_u0_U73 (.A( u0_u14_u0_n138 ) , .B2( u0_u14_u0_n139 ) , .B1( u0_u14_u0_n140 ) , .ZN( u0_u14_u0_n157 ) );
  AOI21_X1 u0_u14_u0_U74 (.B2( u0_u14_u0_n141 ) , .B1( u0_u14_u0_n142 ) , .ZN( u0_u14_u0_n156 ) , .A( u0_u14_u0_n161 ) );
  OR4_X1 u0_u14_u0_U75 (.ZN( u0_out14_17 ) , .A4( u0_u14_u0_n122 ) , .A2( u0_u14_u0_n123 ) , .A1( u0_u14_u0_n124 ) , .A3( u0_u14_u0_n170 ) );
  AOI21_X1 u0_u14_u0_U76 (.B2( u0_u14_u0_n107 ) , .ZN( u0_u14_u0_n124 ) , .B1( u0_u14_u0_n128 ) , .A( u0_u14_u0_n161 ) );
  INV_X1 u0_u14_u0_U77 (.A( u0_u14_u0_n111 ) , .ZN( u0_u14_u0_n170 ) );
  AOI21_X1 u0_u14_u0_U78 (.B1( u0_u14_u0_n132 ) , .ZN( u0_u14_u0_n133 ) , .A( u0_u14_u0_n144 ) , .B2( u0_u14_u0_n166 ) );
  OAI22_X1 u0_u14_u0_U79 (.ZN( u0_u14_u0_n105 ) , .A2( u0_u14_u0_n132 ) , .B1( u0_u14_u0_n146 ) , .A1( u0_u14_u0_n147 ) , .B2( u0_u14_u0_n161 ) );
  AND2_X1 u0_u14_u0_U8 (.A1( u0_u14_u0_n114 ) , .A2( u0_u14_u0_n121 ) , .ZN( u0_u14_u0_n146 ) );
  NAND2_X1 u0_u14_u0_U80 (.ZN( u0_u14_u0_n110 ) , .A2( u0_u14_u0_n132 ) , .A1( u0_u14_u0_n145 ) );
  INV_X1 u0_u14_u0_U81 (.A( u0_u14_u0_n119 ) , .ZN( u0_u14_u0_n167 ) );
  NAND2_X1 u0_u14_u0_U82 (.A2( u0_u14_u0_n103 ) , .ZN( u0_u14_u0_n140 ) , .A1( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U83 (.A1( u0_u14_u0_n101 ) , .ZN( u0_u14_u0_n130 ) , .A2( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U84 (.ZN( u0_u14_u0_n108 ) , .A1( u0_u14_u0_n92 ) , .A2( u0_u14_u0_n94 ) );
  NAND2_X1 u0_u14_u0_U85 (.ZN( u0_u14_u0_n142 ) , .A1( u0_u14_u0_n94 ) , .A2( u0_u14_u0_n95 ) );
  NOR2_X1 u0_u14_u0_U86 (.A2( u0_u14_X_6 ) , .ZN( u0_u14_u0_n100 ) , .A1( u0_u14_u0_n162 ) );
  NOR2_X1 u0_u14_u0_U87 (.A2( u0_u14_X_3 ) , .A1( u0_u14_X_6 ) , .ZN( u0_u14_u0_n94 ) );
  NAND3_X1 u0_u14_u0_U88 (.ZN( u0_out14_23 ) , .A3( u0_u14_u0_n137 ) , .A1( u0_u14_u0_n168 ) , .A2( u0_u14_u0_n171 ) );
  NAND3_X1 u0_u14_u0_U89 (.A3( u0_u14_u0_n127 ) , .A2( u0_u14_u0_n128 ) , .ZN( u0_u14_u0_n135 ) , .A1( u0_u14_u0_n150 ) );
  AND2_X1 u0_u14_u0_U9 (.A1( u0_u14_u0_n131 ) , .ZN( u0_u14_u0_n141 ) , .A2( u0_u14_u0_n150 ) );
  NAND3_X1 u0_u14_u0_U90 (.ZN( u0_u14_u0_n117 ) , .A3( u0_u14_u0_n132 ) , .A2( u0_u14_u0_n139 ) , .A1( u0_u14_u0_n148 ) );
  NAND3_X1 u0_u14_u0_U91 (.ZN( u0_u14_u0_n109 ) , .A2( u0_u14_u0_n114 ) , .A3( u0_u14_u0_n140 ) , .A1( u0_u14_u0_n149 ) );
  NAND3_X1 u0_u14_u0_U92 (.ZN( u0_out14_9 ) , .A3( u0_u14_u0_n106 ) , .A2( u0_u14_u0_n171 ) , .A1( u0_u14_u0_n174 ) );
  NAND3_X1 u0_u14_u0_U93 (.A2( u0_u14_u0_n128 ) , .A1( u0_u14_u0_n132 ) , .A3( u0_u14_u0_n146 ) , .ZN( u0_u14_u0_n97 ) );
  OAI22_X1 u0_u14_u4_U10 (.B2( u0_u14_u4_n135 ) , .ZN( u0_u14_u4_n137 ) , .B1( u0_u14_u4_n153 ) , .A1( u0_u14_u4_n155 ) , .A2( u0_u14_u4_n171 ) );
  AND3_X1 u0_u14_u4_U11 (.A2( u0_u14_u4_n134 ) , .ZN( u0_u14_u4_n135 ) , .A3( u0_u14_u4_n145 ) , .A1( u0_u14_u4_n157 ) );
  NAND2_X1 u0_u14_u4_U12 (.ZN( u0_u14_u4_n132 ) , .A2( u0_u14_u4_n170 ) , .A1( u0_u14_u4_n173 ) );
  AOI21_X1 u0_u14_u4_U13 (.B2( u0_u14_u4_n160 ) , .B1( u0_u14_u4_n161 ) , .ZN( u0_u14_u4_n162 ) , .A( u0_u14_u4_n170 ) );
  AOI21_X1 u0_u14_u4_U14 (.ZN( u0_u14_u4_n107 ) , .B2( u0_u14_u4_n143 ) , .A( u0_u14_u4_n174 ) , .B1( u0_u14_u4_n184 ) );
  AOI21_X1 u0_u14_u4_U15 (.B2( u0_u14_u4_n158 ) , .B1( u0_u14_u4_n159 ) , .ZN( u0_u14_u4_n163 ) , .A( u0_u14_u4_n174 ) );
  AOI21_X1 u0_u14_u4_U16 (.A( u0_u14_u4_n153 ) , .B2( u0_u14_u4_n154 ) , .B1( u0_u14_u4_n155 ) , .ZN( u0_u14_u4_n165 ) );
  AOI21_X1 u0_u14_u4_U17 (.A( u0_u14_u4_n156 ) , .B2( u0_u14_u4_n157 ) , .ZN( u0_u14_u4_n164 ) , .B1( u0_u14_u4_n184 ) );
  INV_X1 u0_u14_u4_U18 (.A( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n170 ) );
  AND2_X1 u0_u14_u4_U19 (.A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n155 ) , .A1( u0_u14_u4_n160 ) );
  INV_X1 u0_u14_u4_U20 (.A( u0_u14_u4_n156 ) , .ZN( u0_u14_u4_n175 ) );
  NAND2_X1 u0_u14_u4_U21 (.A2( u0_u14_u4_n118 ) , .ZN( u0_u14_u4_n131 ) , .A1( u0_u14_u4_n147 ) );
  NAND2_X1 u0_u14_u4_U22 (.A1( u0_u14_u4_n119 ) , .A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n130 ) );
  NAND2_X1 u0_u14_u4_U23 (.ZN( u0_u14_u4_n117 ) , .A2( u0_u14_u4_n118 ) , .A1( u0_u14_u4_n148 ) );
  NAND2_X1 u0_u14_u4_U24 (.ZN( u0_u14_u4_n129 ) , .A1( u0_u14_u4_n134 ) , .A2( u0_u14_u4_n148 ) );
  AND3_X1 u0_u14_u4_U25 (.A1( u0_u14_u4_n119 ) , .A2( u0_u14_u4_n143 ) , .A3( u0_u14_u4_n154 ) , .ZN( u0_u14_u4_n161 ) );
  AND2_X1 u0_u14_u4_U26 (.A1( u0_u14_u4_n145 ) , .A2( u0_u14_u4_n147 ) , .ZN( u0_u14_u4_n159 ) );
  OR3_X1 u0_u14_u4_U27 (.A3( u0_u14_u4_n114 ) , .A2( u0_u14_u4_n115 ) , .A1( u0_u14_u4_n116 ) , .ZN( u0_u14_u4_n136 ) );
  AOI21_X1 u0_u14_u4_U28 (.A( u0_u14_u4_n113 ) , .ZN( u0_u14_u4_n116 ) , .B2( u0_u14_u4_n173 ) , .B1( u0_u14_u4_n174 ) );
  AOI21_X1 u0_u14_u4_U29 (.ZN( u0_u14_u4_n115 ) , .B2( u0_u14_u4_n145 ) , .B1( u0_u14_u4_n146 ) , .A( u0_u14_u4_n156 ) );
  NOR2_X1 u0_u14_u4_U3 (.ZN( u0_u14_u4_n121 ) , .A1( u0_u14_u4_n181 ) , .A2( u0_u14_u4_n182 ) );
  OAI22_X1 u0_u14_u4_U30 (.ZN( u0_u14_u4_n114 ) , .A2( u0_u14_u4_n121 ) , .B1( u0_u14_u4_n160 ) , .B2( u0_u14_u4_n170 ) , .A1( u0_u14_u4_n171 ) );
  INV_X1 u0_u14_u4_U31 (.A( u0_u14_u4_n158 ) , .ZN( u0_u14_u4_n182 ) );
  INV_X1 u0_u14_u4_U32 (.ZN( u0_u14_u4_n181 ) , .A( u0_u14_u4_n96 ) );
  INV_X1 u0_u14_u4_U33 (.A( u0_u14_u4_n144 ) , .ZN( u0_u14_u4_n179 ) );
  INV_X1 u0_u14_u4_U34 (.A( u0_u14_u4_n157 ) , .ZN( u0_u14_u4_n178 ) );
  NAND2_X1 u0_u14_u4_U35 (.A2( u0_u14_u4_n154 ) , .A1( u0_u14_u4_n96 ) , .ZN( u0_u14_u4_n97 ) );
  INV_X1 u0_u14_u4_U36 (.ZN( u0_u14_u4_n186 ) , .A( u0_u14_u4_n95 ) );
  OAI221_X1 u0_u14_u4_U37 (.C1( u0_u14_u4_n134 ) , .B1( u0_u14_u4_n158 ) , .B2( u0_u14_u4_n171 ) , .C2( u0_u14_u4_n173 ) , .A( u0_u14_u4_n94 ) , .ZN( u0_u14_u4_n95 ) );
  AOI222_X1 u0_u14_u4_U38 (.B2( u0_u14_u4_n132 ) , .A1( u0_u14_u4_n138 ) , .C2( u0_u14_u4_n175 ) , .A2( u0_u14_u4_n179 ) , .C1( u0_u14_u4_n181 ) , .B1( u0_u14_u4_n185 ) , .ZN( u0_u14_u4_n94 ) );
  INV_X1 u0_u14_u4_U39 (.A( u0_u14_u4_n113 ) , .ZN( u0_u14_u4_n185 ) );
  INV_X1 u0_u14_u4_U4 (.A( u0_u14_u4_n117 ) , .ZN( u0_u14_u4_n184 ) );
  INV_X1 u0_u14_u4_U40 (.A( u0_u14_u4_n143 ) , .ZN( u0_u14_u4_n183 ) );
  NOR2_X1 u0_u14_u4_U41 (.ZN( u0_u14_u4_n138 ) , .A1( u0_u14_u4_n168 ) , .A2( u0_u14_u4_n169 ) );
  NOR2_X1 u0_u14_u4_U42 (.A1( u0_u14_u4_n150 ) , .A2( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n153 ) );
  NOR2_X1 u0_u14_u4_U43 (.A2( u0_u14_u4_n128 ) , .A1( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n156 ) );
  AOI22_X1 u0_u14_u4_U44 (.B2( u0_u14_u4_n122 ) , .A1( u0_u14_u4_n123 ) , .ZN( u0_u14_u4_n124 ) , .B1( u0_u14_u4_n128 ) , .A2( u0_u14_u4_n172 ) );
  INV_X1 u0_u14_u4_U45 (.A( u0_u14_u4_n153 ) , .ZN( u0_u14_u4_n172 ) );
  NAND2_X1 u0_u14_u4_U46 (.A2( u0_u14_u4_n120 ) , .ZN( u0_u14_u4_n123 ) , .A1( u0_u14_u4_n161 ) );
  AOI22_X1 u0_u14_u4_U47 (.B2( u0_u14_u4_n132 ) , .A2( u0_u14_u4_n133 ) , .ZN( u0_u14_u4_n140 ) , .A1( u0_u14_u4_n150 ) , .B1( u0_u14_u4_n179 ) );
  NAND2_X1 u0_u14_u4_U48 (.ZN( u0_u14_u4_n133 ) , .A2( u0_u14_u4_n146 ) , .A1( u0_u14_u4_n154 ) );
  NAND2_X1 u0_u14_u4_U49 (.A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n154 ) , .A2( u0_u14_u4_n98 ) );
  NOR4_X1 u0_u14_u4_U5 (.A4( u0_u14_u4_n106 ) , .A3( u0_u14_u4_n107 ) , .A2( u0_u14_u4_n108 ) , .A1( u0_u14_u4_n109 ) , .ZN( u0_u14_u4_n110 ) );
  NAND2_X1 u0_u14_u4_U50 (.A1( u0_u14_u4_n101 ) , .ZN( u0_u14_u4_n158 ) , .A2( u0_u14_u4_n99 ) );
  AOI21_X1 u0_u14_u4_U51 (.ZN( u0_u14_u4_n127 ) , .A( u0_u14_u4_n136 ) , .B2( u0_u14_u4_n150 ) , .B1( u0_u14_u4_n180 ) );
  INV_X1 u0_u14_u4_U52 (.A( u0_u14_u4_n160 ) , .ZN( u0_u14_u4_n180 ) );
  NAND2_X1 u0_u14_u4_U53 (.A2( u0_u14_u4_n104 ) , .A1( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n146 ) );
  NAND2_X1 u0_u14_u4_U54 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n160 ) );
  NAND2_X1 u0_u14_u4_U55 (.ZN( u0_u14_u4_n134 ) , .A1( u0_u14_u4_n98 ) , .A2( u0_u14_u4_n99 ) );
  NAND2_X1 u0_u14_u4_U56 (.A1( u0_u14_u4_n103 ) , .A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n143 ) );
  NAND2_X1 u0_u14_u4_U57 (.A2( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n145 ) , .A1( u0_u14_u4_n98 ) );
  NAND2_X1 u0_u14_u4_U58 (.A1( u0_u14_u4_n100 ) , .A2( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n120 ) );
  NAND2_X1 u0_u14_u4_U59 (.A1( u0_u14_u4_n102 ) , .A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n148 ) );
  AOI21_X1 u0_u14_u4_U6 (.ZN( u0_u14_u4_n106 ) , .B2( u0_u14_u4_n146 ) , .B1( u0_u14_u4_n158 ) , .A( u0_u14_u4_n170 ) );
  NAND2_X1 u0_u14_u4_U60 (.A2( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n157 ) );
  INV_X1 u0_u14_u4_U61 (.A( u0_u14_u4_n150 ) , .ZN( u0_u14_u4_n173 ) );
  INV_X1 u0_u14_u4_U62 (.A( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n171 ) );
  NAND2_X1 u0_u14_u4_U63 (.A1( u0_u14_u4_n100 ) , .ZN( u0_u14_u4_n118 ) , .A2( u0_u14_u4_n99 ) );
  NAND2_X1 u0_u14_u4_U64 (.A2( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n144 ) );
  NAND2_X1 u0_u14_u4_U65 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n105 ) , .ZN( u0_u14_u4_n96 ) );
  INV_X1 u0_u14_u4_U66 (.A( u0_u14_u4_n128 ) , .ZN( u0_u14_u4_n174 ) );
  NAND2_X1 u0_u14_u4_U67 (.A2( u0_u14_u4_n102 ) , .ZN( u0_u14_u4_n119 ) , .A1( u0_u14_u4_n98 ) );
  NAND2_X1 u0_u14_u4_U68 (.A2( u0_u14_u4_n101 ) , .A1( u0_u14_u4_n103 ) , .ZN( u0_u14_u4_n147 ) );
  NAND2_X1 u0_u14_u4_U69 (.A2( u0_u14_u4_n104 ) , .ZN( u0_u14_u4_n113 ) , .A1( u0_u14_u4_n99 ) );
  AOI21_X1 u0_u14_u4_U7 (.ZN( u0_u14_u4_n108 ) , .B2( u0_u14_u4_n134 ) , .B1( u0_u14_u4_n155 ) , .A( u0_u14_u4_n156 ) );
  NOR2_X1 u0_u14_u4_U70 (.A2( u0_u14_X_28 ) , .ZN( u0_u14_u4_n150 ) , .A1( u0_u14_u4_n168 ) );
  NOR2_X1 u0_u14_u4_U71 (.A2( u0_u14_X_29 ) , .ZN( u0_u14_u4_n152 ) , .A1( u0_u14_u4_n169 ) );
  NOR2_X1 u0_u14_u4_U72 (.A2( u0_u14_X_30 ) , .ZN( u0_u14_u4_n105 ) , .A1( u0_u14_u4_n176 ) );
  NOR2_X1 u0_u14_u4_U73 (.A2( u0_u14_X_26 ) , .ZN( u0_u14_u4_n100 ) , .A1( u0_u14_u4_n177 ) );
  NOR2_X1 u0_u14_u4_U74 (.A2( u0_u14_X_28 ) , .A1( u0_u14_X_29 ) , .ZN( u0_u14_u4_n128 ) );
  NOR2_X1 u0_u14_u4_U75 (.A2( u0_u14_X_27 ) , .A1( u0_u14_X_30 ) , .ZN( u0_u14_u4_n102 ) );
  NOR2_X1 u0_u14_u4_U76 (.A2( u0_u14_X_25 ) , .A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n98 ) );
  AND2_X1 u0_u14_u4_U77 (.A2( u0_u14_X_25 ) , .A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n104 ) );
  AND2_X1 u0_u14_u4_U78 (.A1( u0_u14_X_30 ) , .A2( u0_u14_u4_n176 ) , .ZN( u0_u14_u4_n99 ) );
  AND2_X1 u0_u14_u4_U79 (.A1( u0_u14_X_26 ) , .ZN( u0_u14_u4_n101 ) , .A2( u0_u14_u4_n177 ) );
  AOI21_X1 u0_u14_u4_U8 (.ZN( u0_u14_u4_n109 ) , .A( u0_u14_u4_n153 ) , .B1( u0_u14_u4_n159 ) , .B2( u0_u14_u4_n184 ) );
  AND2_X1 u0_u14_u4_U80 (.A1( u0_u14_X_27 ) , .A2( u0_u14_X_30 ) , .ZN( u0_u14_u4_n103 ) );
  INV_X1 u0_u14_u4_U81 (.A( u0_u14_X_28 ) , .ZN( u0_u14_u4_n169 ) );
  INV_X1 u0_u14_u4_U82 (.A( u0_u14_X_29 ) , .ZN( u0_u14_u4_n168 ) );
  INV_X1 u0_u14_u4_U83 (.A( u0_u14_X_25 ) , .ZN( u0_u14_u4_n177 ) );
  INV_X1 u0_u14_u4_U84 (.A( u0_u14_X_27 ) , .ZN( u0_u14_u4_n176 ) );
  NAND4_X1 u0_u14_u4_U85 (.ZN( u0_out14_25 ) , .A4( u0_u14_u4_n139 ) , .A3( u0_u14_u4_n140 ) , .A2( u0_u14_u4_n141 ) , .A1( u0_u14_u4_n142 ) );
  OAI21_X1 u0_u14_u4_U86 (.A( u0_u14_u4_n128 ) , .B2( u0_u14_u4_n129 ) , .B1( u0_u14_u4_n130 ) , .ZN( u0_u14_u4_n142 ) );
  OAI21_X1 u0_u14_u4_U87 (.B2( u0_u14_u4_n131 ) , .ZN( u0_u14_u4_n141 ) , .A( u0_u14_u4_n175 ) , .B1( u0_u14_u4_n183 ) );
  NAND4_X1 u0_u14_u4_U88 (.ZN( u0_out14_14 ) , .A4( u0_u14_u4_n124 ) , .A3( u0_u14_u4_n125 ) , .A2( u0_u14_u4_n126 ) , .A1( u0_u14_u4_n127 ) );
  AOI22_X1 u0_u14_u4_U89 (.B2( u0_u14_u4_n117 ) , .ZN( u0_u14_u4_n126 ) , .A1( u0_u14_u4_n129 ) , .B1( u0_u14_u4_n152 ) , .A2( u0_u14_u4_n175 ) );
  AOI211_X1 u0_u14_u4_U9 (.B( u0_u14_u4_n136 ) , .A( u0_u14_u4_n137 ) , .C2( u0_u14_u4_n138 ) , .ZN( u0_u14_u4_n139 ) , .C1( u0_u14_u4_n182 ) );
  AOI22_X1 u0_u14_u4_U90 (.ZN( u0_u14_u4_n125 ) , .B2( u0_u14_u4_n131 ) , .A2( u0_u14_u4_n132 ) , .B1( u0_u14_u4_n138 ) , .A1( u0_u14_u4_n178 ) );
  NAND4_X1 u0_u14_u4_U91 (.ZN( u0_out14_8 ) , .A4( u0_u14_u4_n110 ) , .A3( u0_u14_u4_n111 ) , .A2( u0_u14_u4_n112 ) , .A1( u0_u14_u4_n186 ) );
  NAND2_X1 u0_u14_u4_U92 (.ZN( u0_u14_u4_n112 ) , .A2( u0_u14_u4_n130 ) , .A1( u0_u14_u4_n150 ) );
  AOI22_X1 u0_u14_u4_U93 (.ZN( u0_u14_u4_n111 ) , .B2( u0_u14_u4_n132 ) , .A1( u0_u14_u4_n152 ) , .B1( u0_u14_u4_n178 ) , .A2( u0_u14_u4_n97 ) );
  AOI22_X1 u0_u14_u4_U94 (.B2( u0_u14_u4_n149 ) , .B1( u0_u14_u4_n150 ) , .A2( u0_u14_u4_n151 ) , .A1( u0_u14_u4_n152 ) , .ZN( u0_u14_u4_n167 ) );
  NOR4_X1 u0_u14_u4_U95 (.A4( u0_u14_u4_n162 ) , .A3( u0_u14_u4_n163 ) , .A2( u0_u14_u4_n164 ) , .A1( u0_u14_u4_n165 ) , .ZN( u0_u14_u4_n166 ) );
  NAND3_X1 u0_u14_u4_U96 (.ZN( u0_out14_3 ) , .A3( u0_u14_u4_n166 ) , .A1( u0_u14_u4_n167 ) , .A2( u0_u14_u4_n186 ) );
  NAND3_X1 u0_u14_u4_U97 (.A3( u0_u14_u4_n146 ) , .A2( u0_u14_u4_n147 ) , .A1( u0_u14_u4_n148 ) , .ZN( u0_u14_u4_n149 ) );
  NAND3_X1 u0_u14_u4_U98 (.A3( u0_u14_u4_n143 ) , .A2( u0_u14_u4_n144 ) , .A1( u0_u14_u4_n145 ) , .ZN( u0_u14_u4_n151 ) );
  NAND3_X1 u0_u14_u4_U99 (.A3( u0_u14_u4_n121 ) , .ZN( u0_u14_u4_n122 ) , .A2( u0_u14_u4_n144 ) , .A1( u0_u14_u4_n154 ) );
  AOI21_X1 u0_u14_u6_U10 (.ZN( u0_u14_u6_n106 ) , .A( u0_u14_u6_n142 ) , .B2( u0_u14_u6_n159 ) , .B1( u0_u14_u6_n164 ) );
  INV_X1 u0_u14_u6_U11 (.A( u0_u14_u6_n155 ) , .ZN( u0_u14_u6_n161 ) );
  INV_X1 u0_u14_u6_U12 (.A( u0_u14_u6_n128 ) , .ZN( u0_u14_u6_n164 ) );
  NAND2_X1 u0_u14_u6_U13 (.ZN( u0_u14_u6_n110 ) , .A1( u0_u14_u6_n122 ) , .A2( u0_u14_u6_n129 ) );
  NAND2_X1 u0_u14_u6_U14 (.ZN( u0_u14_u6_n124 ) , .A2( u0_u14_u6_n146 ) , .A1( u0_u14_u6_n148 ) );
  INV_X1 u0_u14_u6_U15 (.A( u0_u14_u6_n132 ) , .ZN( u0_u14_u6_n171 ) );
  AND2_X1 u0_u14_u6_U16 (.A1( u0_u14_u6_n100 ) , .ZN( u0_u14_u6_n130 ) , .A2( u0_u14_u6_n147 ) );
  INV_X1 u0_u14_u6_U17 (.A( u0_u14_u6_n127 ) , .ZN( u0_u14_u6_n173 ) );
  INV_X1 u0_u14_u6_U18 (.A( u0_u14_u6_n121 ) , .ZN( u0_u14_u6_n167 ) );
  INV_X1 u0_u14_u6_U19 (.A( u0_u14_u6_n100 ) , .ZN( u0_u14_u6_n169 ) );
  INV_X1 u0_u14_u6_U20 (.A( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n170 ) );
  INV_X1 u0_u14_u6_U21 (.A( u0_u14_u6_n113 ) , .ZN( u0_u14_u6_n168 ) );
  AND2_X1 u0_u14_u6_U22 (.A1( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n119 ) , .ZN( u0_u14_u6_n133 ) );
  AND2_X1 u0_u14_u6_U23 (.A2( u0_u14_u6_n121 ) , .A1( u0_u14_u6_n122 ) , .ZN( u0_u14_u6_n131 ) );
  AND3_X1 u0_u14_u6_U24 (.ZN( u0_u14_u6_n120 ) , .A2( u0_u14_u6_n127 ) , .A1( u0_u14_u6_n132 ) , .A3( u0_u14_u6_n145 ) );
  INV_X1 u0_u14_u6_U25 (.A( u0_u14_u6_n146 ) , .ZN( u0_u14_u6_n163 ) );
  AOI222_X1 u0_u14_u6_U26 (.ZN( u0_u14_u6_n114 ) , .A1( u0_u14_u6_n118 ) , .A2( u0_u14_u6_n126 ) , .B2( u0_u14_u6_n151 ) , .C2( u0_u14_u6_n159 ) , .C1( u0_u14_u6_n168 ) , .B1( u0_u14_u6_n169 ) );
  NOR2_X1 u0_u14_u6_U27 (.A1( u0_u14_u6_n162 ) , .A2( u0_u14_u6_n165 ) , .ZN( u0_u14_u6_n98 ) );
  AOI211_X1 u0_u14_u6_U28 (.B( u0_u14_u6_n149 ) , .A( u0_u14_u6_n150 ) , .C2( u0_u14_u6_n151 ) , .C1( u0_u14_u6_n152 ) , .ZN( u0_u14_u6_n153 ) );
  AOI21_X1 u0_u14_u6_U29 (.B2( u0_u14_u6_n147 ) , .B1( u0_u14_u6_n148 ) , .ZN( u0_u14_u6_n149 ) , .A( u0_u14_u6_n158 ) );
  INV_X1 u0_u14_u6_U3 (.A( u0_u14_u6_n110 ) , .ZN( u0_u14_u6_n166 ) );
  AOI21_X1 u0_u14_u6_U30 (.A( u0_u14_u6_n144 ) , .B2( u0_u14_u6_n145 ) , .B1( u0_u14_u6_n146 ) , .ZN( u0_u14_u6_n150 ) );
  NAND2_X1 u0_u14_u6_U31 (.A2( u0_u14_u6_n143 ) , .ZN( u0_u14_u6_n152 ) , .A1( u0_u14_u6_n166 ) );
  NAND2_X1 u0_u14_u6_U32 (.A1( u0_u14_u6_n144 ) , .ZN( u0_u14_u6_n151 ) , .A2( u0_u14_u6_n158 ) );
  NAND2_X1 u0_u14_u6_U33 (.ZN( u0_u14_u6_n132 ) , .A1( u0_u14_u6_n91 ) , .A2( u0_u14_u6_n97 ) );
  AOI22_X1 u0_u14_u6_U34 (.B2( u0_u14_u6_n110 ) , .B1( u0_u14_u6_n111 ) , .A1( u0_u14_u6_n112 ) , .ZN( u0_u14_u6_n115 ) , .A2( u0_u14_u6_n161 ) );
  NAND4_X1 u0_u14_u6_U35 (.A3( u0_u14_u6_n109 ) , .ZN( u0_u14_u6_n112 ) , .A4( u0_u14_u6_n132 ) , .A2( u0_u14_u6_n147 ) , .A1( u0_u14_u6_n166 ) );
  NOR2_X1 u0_u14_u6_U36 (.ZN( u0_u14_u6_n109 ) , .A1( u0_u14_u6_n170 ) , .A2( u0_u14_u6_n173 ) );
  NOR2_X1 u0_u14_u6_U37 (.A2( u0_u14_u6_n126 ) , .ZN( u0_u14_u6_n155 ) , .A1( u0_u14_u6_n160 ) );
  NAND2_X1 u0_u14_u6_U38 (.ZN( u0_u14_u6_n146 ) , .A2( u0_u14_u6_n94 ) , .A1( u0_u14_u6_n99 ) );
  AOI211_X1 u0_u14_u6_U39 (.B( u0_u14_u6_n134 ) , .A( u0_u14_u6_n135 ) , .C1( u0_u14_u6_n136 ) , .ZN( u0_u14_u6_n137 ) , .C2( u0_u14_u6_n151 ) );
  AOI22_X1 u0_u14_u6_U4 (.B2( u0_u14_u6_n101 ) , .A1( u0_u14_u6_n102 ) , .ZN( u0_u14_u6_n103 ) , .B1( u0_u14_u6_n160 ) , .A2( u0_u14_u6_n161 ) );
  AOI21_X1 u0_u14_u6_U40 (.B2( u0_u14_u6_n132 ) , .B1( u0_u14_u6_n133 ) , .ZN( u0_u14_u6_n134 ) , .A( u0_u14_u6_n158 ) );
  NAND4_X1 u0_u14_u6_U41 (.A4( u0_u14_u6_n127 ) , .A3( u0_u14_u6_n128 ) , .A2( u0_u14_u6_n129 ) , .A1( u0_u14_u6_n130 ) , .ZN( u0_u14_u6_n136 ) );
  AOI21_X1 u0_u14_u6_U42 (.B1( u0_u14_u6_n131 ) , .ZN( u0_u14_u6_n135 ) , .A( u0_u14_u6_n144 ) , .B2( u0_u14_u6_n146 ) );
  INV_X1 u0_u14_u6_U43 (.A( u0_u14_u6_n111 ) , .ZN( u0_u14_u6_n158 ) );
  NAND2_X1 u0_u14_u6_U44 (.ZN( u0_u14_u6_n127 ) , .A1( u0_u14_u6_n91 ) , .A2( u0_u14_u6_n92 ) );
  NAND2_X1 u0_u14_u6_U45 (.ZN( u0_u14_u6_n129 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n96 ) );
  INV_X1 u0_u14_u6_U46 (.A( u0_u14_u6_n144 ) , .ZN( u0_u14_u6_n159 ) );
  NAND2_X1 u0_u14_u6_U47 (.ZN( u0_u14_u6_n145 ) , .A2( u0_u14_u6_n97 ) , .A1( u0_u14_u6_n98 ) );
  NAND2_X1 u0_u14_u6_U48 (.ZN( u0_u14_u6_n148 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n94 ) );
  NAND2_X1 u0_u14_u6_U49 (.ZN( u0_u14_u6_n108 ) , .A2( u0_u14_u6_n139 ) , .A1( u0_u14_u6_n144 ) );
  NOR2_X1 u0_u14_u6_U5 (.A1( u0_u14_u6_n118 ) , .ZN( u0_u14_u6_n143 ) , .A2( u0_u14_u6_n168 ) );
  NAND2_X1 u0_u14_u6_U50 (.ZN( u0_u14_u6_n121 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n97 ) );
  NAND2_X1 u0_u14_u6_U51 (.ZN( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n95 ) );
  AND2_X1 u0_u14_u6_U52 (.ZN( u0_u14_u6_n118 ) , .A2( u0_u14_u6_n91 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U53 (.ZN( u0_u14_u6_n147 ) , .A2( u0_u14_u6_n98 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U54 (.ZN( u0_u14_u6_n128 ) , .A1( u0_u14_u6_n94 ) , .A2( u0_u14_u6_n96 ) );
  NAND2_X1 u0_u14_u6_U55 (.ZN( u0_u14_u6_n119 ) , .A2( u0_u14_u6_n95 ) , .A1( u0_u14_u6_n99 ) );
  NAND2_X1 u0_u14_u6_U56 (.ZN( u0_u14_u6_n123 ) , .A2( u0_u14_u6_n91 ) , .A1( u0_u14_u6_n96 ) );
  NAND2_X1 u0_u14_u6_U57 (.ZN( u0_u14_u6_n100 ) , .A2( u0_u14_u6_n92 ) , .A1( u0_u14_u6_n98 ) );
  NAND2_X1 u0_u14_u6_U58 (.ZN( u0_u14_u6_n122 ) , .A1( u0_u14_u6_n94 ) , .A2( u0_u14_u6_n97 ) );
  INV_X1 u0_u14_u6_U59 (.A( u0_u14_u6_n139 ) , .ZN( u0_u14_u6_n160 ) );
  INV_X1 u0_u14_u6_U6 (.ZN( u0_u14_u6_n172 ) , .A( u0_u14_u6_n88 ) );
  NAND2_X1 u0_u14_u6_U60 (.ZN( u0_u14_u6_n113 ) , .A1( u0_u14_u6_n96 ) , .A2( u0_u14_u6_n98 ) );
  NOR2_X1 u0_u14_u6_U61 (.A2( u0_u14_X_40 ) , .A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n126 ) );
  NOR2_X1 u0_u14_u6_U62 (.A2( u0_u14_X_39 ) , .A1( u0_u14_X_42 ) , .ZN( u0_u14_u6_n92 ) );
  NOR2_X1 u0_u14_u6_U63 (.A2( u0_u14_X_39 ) , .A1( u0_u14_u6_n156 ) , .ZN( u0_u14_u6_n97 ) );
  NOR2_X1 u0_u14_u6_U64 (.A2( u0_u14_X_38 ) , .A1( u0_u14_u6_n165 ) , .ZN( u0_u14_u6_n95 ) );
  NOR2_X1 u0_u14_u6_U65 (.A2( u0_u14_X_41 ) , .ZN( u0_u14_u6_n111 ) , .A1( u0_u14_u6_n157 ) );
  NOR2_X1 u0_u14_u6_U66 (.A2( u0_u14_X_37 ) , .A1( u0_u14_u6_n162 ) , .ZN( u0_u14_u6_n94 ) );
  NOR2_X1 u0_u14_u6_U67 (.A2( u0_u14_X_37 ) , .A1( u0_u14_X_38 ) , .ZN( u0_u14_u6_n91 ) );
  NAND2_X1 u0_u14_u6_U68 (.A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n144 ) , .A2( u0_u14_u6_n157 ) );
  NAND2_X1 u0_u14_u6_U69 (.A2( u0_u14_X_40 ) , .A1( u0_u14_X_41 ) , .ZN( u0_u14_u6_n139 ) );
  OAI21_X1 u0_u14_u6_U7 (.A( u0_u14_u6_n159 ) , .B1( u0_u14_u6_n169 ) , .B2( u0_u14_u6_n173 ) , .ZN( u0_u14_u6_n90 ) );
  AND2_X1 u0_u14_u6_U70 (.A1( u0_u14_X_39 ) , .A2( u0_u14_u6_n156 ) , .ZN( u0_u14_u6_n96 ) );
  AND2_X1 u0_u14_u6_U71 (.A1( u0_u14_X_39 ) , .A2( u0_u14_X_42 ) , .ZN( u0_u14_u6_n99 ) );
  INV_X1 u0_u14_u6_U72 (.A( u0_u14_X_40 ) , .ZN( u0_u14_u6_n157 ) );
  INV_X1 u0_u14_u6_U73 (.A( u0_u14_X_37 ) , .ZN( u0_u14_u6_n165 ) );
  INV_X1 u0_u14_u6_U74 (.A( u0_u14_X_38 ) , .ZN( u0_u14_u6_n162 ) );
  INV_X1 u0_u14_u6_U75 (.A( u0_u14_X_42 ) , .ZN( u0_u14_u6_n156 ) );
  NAND4_X1 u0_u14_u6_U76 (.ZN( u0_out14_32 ) , .A4( u0_u14_u6_n103 ) , .A3( u0_u14_u6_n104 ) , .A2( u0_u14_u6_n105 ) , .A1( u0_u14_u6_n106 ) );
  AOI22_X1 u0_u14_u6_U77 (.ZN( u0_u14_u6_n105 ) , .A2( u0_u14_u6_n108 ) , .A1( u0_u14_u6_n118 ) , .B2( u0_u14_u6_n126 ) , .B1( u0_u14_u6_n171 ) );
  AOI22_X1 u0_u14_u6_U78 (.ZN( u0_u14_u6_n104 ) , .A1( u0_u14_u6_n111 ) , .B1( u0_u14_u6_n124 ) , .B2( u0_u14_u6_n151 ) , .A2( u0_u14_u6_n93 ) );
  NAND4_X1 u0_u14_u6_U79 (.ZN( u0_out14_12 ) , .A4( u0_u14_u6_n114 ) , .A3( u0_u14_u6_n115 ) , .A2( u0_u14_u6_n116 ) , .A1( u0_u14_u6_n117 ) );
  AOI22_X1 u0_u14_u6_U8 (.A2( u0_u14_u6_n151 ) , .B2( u0_u14_u6_n161 ) , .A1( u0_u14_u6_n167 ) , .B1( u0_u14_u6_n170 ) , .ZN( u0_u14_u6_n89 ) );
  OAI22_X1 u0_u14_u6_U80 (.B2( u0_u14_u6_n111 ) , .ZN( u0_u14_u6_n116 ) , .B1( u0_u14_u6_n126 ) , .A2( u0_u14_u6_n164 ) , .A1( u0_u14_u6_n167 ) );
  OAI21_X1 u0_u14_u6_U81 (.A( u0_u14_u6_n108 ) , .ZN( u0_u14_u6_n117 ) , .B2( u0_u14_u6_n141 ) , .B1( u0_u14_u6_n163 ) );
  OAI211_X1 u0_u14_u6_U82 (.ZN( u0_out14_22 ) , .B( u0_u14_u6_n137 ) , .A( u0_u14_u6_n138 ) , .C2( u0_u14_u6_n139 ) , .C1( u0_u14_u6_n140 ) );
  AOI22_X1 u0_u14_u6_U83 (.B1( u0_u14_u6_n124 ) , .A2( u0_u14_u6_n125 ) , .A1( u0_u14_u6_n126 ) , .ZN( u0_u14_u6_n138 ) , .B2( u0_u14_u6_n161 ) );
  AND4_X1 u0_u14_u6_U84 (.A3( u0_u14_u6_n119 ) , .A1( u0_u14_u6_n120 ) , .A4( u0_u14_u6_n129 ) , .ZN( u0_u14_u6_n140 ) , .A2( u0_u14_u6_n143 ) );
  OAI211_X1 u0_u14_u6_U85 (.ZN( u0_out14_7 ) , .B( u0_u14_u6_n153 ) , .C2( u0_u14_u6_n154 ) , .C1( u0_u14_u6_n155 ) , .A( u0_u14_u6_n174 ) );
  NOR3_X1 u0_u14_u6_U86 (.A1( u0_u14_u6_n141 ) , .ZN( u0_u14_u6_n154 ) , .A3( u0_u14_u6_n164 ) , .A2( u0_u14_u6_n171 ) );
  INV_X1 u0_u14_u6_U87 (.A( u0_u14_u6_n142 ) , .ZN( u0_u14_u6_n174 ) );
  NAND3_X1 u0_u14_u6_U88 (.A2( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n125 ) , .A1( u0_u14_u6_n130 ) , .A3( u0_u14_u6_n131 ) );
  NAND3_X1 u0_u14_u6_U89 (.A3( u0_u14_u6_n133 ) , .ZN( u0_u14_u6_n141 ) , .A1( u0_u14_u6_n145 ) , .A2( u0_u14_u6_n148 ) );
  AOI21_X1 u0_u14_u6_U9 (.B1( u0_u14_u6_n107 ) , .B2( u0_u14_u6_n132 ) , .A( u0_u14_u6_n158 ) , .ZN( u0_u14_u6_n88 ) );
  NAND3_X1 u0_u14_u6_U90 (.ZN( u0_u14_u6_n101 ) , .A3( u0_u14_u6_n107 ) , .A2( u0_u14_u6_n121 ) , .A1( u0_u14_u6_n127 ) );
  NAND3_X1 u0_u14_u6_U91 (.ZN( u0_u14_u6_n102 ) , .A3( u0_u14_u6_n130 ) , .A2( u0_u14_u6_n145 ) , .A1( u0_u14_u6_n166 ) );
  NAND3_X1 u0_u14_u6_U92 (.A3( u0_u14_u6_n113 ) , .A1( u0_u14_u6_n119 ) , .A2( u0_u14_u6_n123 ) , .ZN( u0_u14_u6_n93 ) );
  NAND3_X1 u0_u14_u6_U93 (.ZN( u0_u14_u6_n142 ) , .A2( u0_u14_u6_n172 ) , .A3( u0_u14_u6_n89 ) , .A1( u0_u14_u6_n90 ) );
  AND3_X1 u0_u14_u7_U10 (.A3( u0_u14_u7_n110 ) , .A2( u0_u14_u7_n127 ) , .A1( u0_u14_u7_n132 ) , .ZN( u0_u14_u7_n92 ) );
  OAI21_X1 u0_u14_u7_U11 (.A( u0_u14_u7_n161 ) , .B1( u0_u14_u7_n168 ) , .B2( u0_u14_u7_n173 ) , .ZN( u0_u14_u7_n91 ) );
  AOI211_X1 u0_u14_u7_U12 (.A( u0_u14_u7_n117 ) , .ZN( u0_u14_u7_n118 ) , .C2( u0_u14_u7_n126 ) , .C1( u0_u14_u7_n177 ) , .B( u0_u14_u7_n180 ) );
  OAI22_X1 u0_u14_u7_U13 (.B1( u0_u14_u7_n115 ) , .ZN( u0_u14_u7_n117 ) , .A2( u0_u14_u7_n133 ) , .A1( u0_u14_u7_n137 ) , .B2( u0_u14_u7_n162 ) );
  INV_X1 u0_u14_u7_U14 (.A( u0_u14_u7_n116 ) , .ZN( u0_u14_u7_n180 ) );
  NOR3_X1 u0_u14_u7_U15 (.ZN( u0_u14_u7_n115 ) , .A3( u0_u14_u7_n145 ) , .A2( u0_u14_u7_n168 ) , .A1( u0_u14_u7_n169 ) );
  NOR3_X1 u0_u14_u7_U16 (.A2( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n135 ) , .ZN( u0_u14_u7_n136 ) , .A3( u0_u14_u7_n171 ) );
  NOR2_X1 u0_u14_u7_U17 (.A1( u0_u14_u7_n130 ) , .A2( u0_u14_u7_n134 ) , .ZN( u0_u14_u7_n153 ) );
  NOR2_X1 u0_u14_u7_U18 (.ZN( u0_u14_u7_n111 ) , .A2( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n169 ) );
  AOI21_X1 u0_u14_u7_U19 (.ZN( u0_u14_u7_n104 ) , .B2( u0_u14_u7_n112 ) , .B1( u0_u14_u7_n127 ) , .A( u0_u14_u7_n164 ) );
  AOI21_X1 u0_u14_u7_U20 (.ZN( u0_u14_u7_n106 ) , .B1( u0_u14_u7_n133 ) , .B2( u0_u14_u7_n146 ) , .A( u0_u14_u7_n162 ) );
  AOI21_X1 u0_u14_u7_U21 (.A( u0_u14_u7_n101 ) , .ZN( u0_u14_u7_n107 ) , .B2( u0_u14_u7_n128 ) , .B1( u0_u14_u7_n175 ) );
  INV_X1 u0_u14_u7_U22 (.A( u0_u14_u7_n101 ) , .ZN( u0_u14_u7_n165 ) );
  INV_X1 u0_u14_u7_U23 (.A( u0_u14_u7_n138 ) , .ZN( u0_u14_u7_n171 ) );
  INV_X1 u0_u14_u7_U24 (.A( u0_u14_u7_n131 ) , .ZN( u0_u14_u7_n177 ) );
  INV_X1 u0_u14_u7_U25 (.A( u0_u14_u7_n110 ) , .ZN( u0_u14_u7_n174 ) );
  NAND2_X1 u0_u14_u7_U26 (.A1( u0_u14_u7_n129 ) , .A2( u0_u14_u7_n132 ) , .ZN( u0_u14_u7_n149 ) );
  NAND2_X1 u0_u14_u7_U27 (.A1( u0_u14_u7_n113 ) , .A2( u0_u14_u7_n124 ) , .ZN( u0_u14_u7_n130 ) );
  INV_X1 u0_u14_u7_U28 (.A( u0_u14_u7_n128 ) , .ZN( u0_u14_u7_n168 ) );
  INV_X1 u0_u14_u7_U29 (.A( u0_u14_u7_n148 ) , .ZN( u0_u14_u7_n169 ) );
  INV_X1 u0_u14_u7_U3 (.A( u0_u14_u7_n149 ) , .ZN( u0_u14_u7_n175 ) );
  INV_X1 u0_u14_u7_U30 (.A( u0_u14_u7_n112 ) , .ZN( u0_u14_u7_n173 ) );
  INV_X1 u0_u14_u7_U31 (.A( u0_u14_u7_n127 ) , .ZN( u0_u14_u7_n179 ) );
  NOR2_X1 u0_u14_u7_U32 (.ZN( u0_u14_u7_n101 ) , .A2( u0_u14_u7_n150 ) , .A1( u0_u14_u7_n156 ) );
  AOI211_X1 u0_u14_u7_U33 (.B( u0_u14_u7_n154 ) , .A( u0_u14_u7_n155 ) , .C1( u0_u14_u7_n156 ) , .ZN( u0_u14_u7_n157 ) , .C2( u0_u14_u7_n172 ) );
  INV_X1 u0_u14_u7_U34 (.A( u0_u14_u7_n153 ) , .ZN( u0_u14_u7_n172 ) );
  AOI211_X1 u0_u14_u7_U35 (.B( u0_u14_u7_n139 ) , .A( u0_u14_u7_n140 ) , .C2( u0_u14_u7_n141 ) , .ZN( u0_u14_u7_n142 ) , .C1( u0_u14_u7_n156 ) );
  NAND4_X1 u0_u14_u7_U36 (.A3( u0_u14_u7_n127 ) , .A2( u0_u14_u7_n128 ) , .A1( u0_u14_u7_n129 ) , .ZN( u0_u14_u7_n141 ) , .A4( u0_u14_u7_n147 ) );
  AOI21_X1 u0_u14_u7_U37 (.A( u0_u14_u7_n137 ) , .B1( u0_u14_u7_n138 ) , .ZN( u0_u14_u7_n139 ) , .B2( u0_u14_u7_n146 ) );
  OAI22_X1 u0_u14_u7_U38 (.B1( u0_u14_u7_n136 ) , .ZN( u0_u14_u7_n140 ) , .A1( u0_u14_u7_n153 ) , .B2( u0_u14_u7_n162 ) , .A2( u0_u14_u7_n164 ) );
  INV_X1 u0_u14_u7_U39 (.A( u0_u14_u7_n125 ) , .ZN( u0_u14_u7_n161 ) );
  INV_X1 u0_u14_u7_U4 (.A( u0_u14_u7_n154 ) , .ZN( u0_u14_u7_n178 ) );
  AOI21_X1 u0_u14_u7_U40 (.ZN( u0_u14_u7_n123 ) , .B1( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n177 ) , .A( u0_u14_u7_n97 ) );
  AOI21_X1 u0_u14_u7_U41 (.B2( u0_u14_u7_n113 ) , .B1( u0_u14_u7_n124 ) , .A( u0_u14_u7_n125 ) , .ZN( u0_u14_u7_n97 ) );
  INV_X1 u0_u14_u7_U42 (.A( u0_u14_u7_n152 ) , .ZN( u0_u14_u7_n162 ) );
  AOI22_X1 u0_u14_u7_U43 (.A2( u0_u14_u7_n114 ) , .ZN( u0_u14_u7_n119 ) , .B1( u0_u14_u7_n130 ) , .A1( u0_u14_u7_n156 ) , .B2( u0_u14_u7_n165 ) );
  NAND2_X1 u0_u14_u7_U44 (.A2( u0_u14_u7_n112 ) , .ZN( u0_u14_u7_n114 ) , .A1( u0_u14_u7_n175 ) );
  AOI22_X1 u0_u14_u7_U45 (.B2( u0_u14_u7_n149 ) , .B1( u0_u14_u7_n150 ) , .A2( u0_u14_u7_n151 ) , .A1( u0_u14_u7_n152 ) , .ZN( u0_u14_u7_n158 ) );
  NOR2_X1 u0_u14_u7_U46 (.ZN( u0_u14_u7_n137 ) , .A1( u0_u14_u7_n150 ) , .A2( u0_u14_u7_n161 ) );
  AND2_X1 u0_u14_u7_U47 (.ZN( u0_u14_u7_n145 ) , .A2( u0_u14_u7_n98 ) , .A1( u0_u14_u7_n99 ) );
  AOI21_X1 u0_u14_u7_U48 (.ZN( u0_u14_u7_n105 ) , .B2( u0_u14_u7_n110 ) , .A( u0_u14_u7_n125 ) , .B1( u0_u14_u7_n147 ) );
  NAND2_X1 u0_u14_u7_U49 (.ZN( u0_u14_u7_n146 ) , .A1( u0_u14_u7_n95 ) , .A2( u0_u14_u7_n98 ) );
  INV_X1 u0_u14_u7_U5 (.A( u0_u14_u7_n111 ) , .ZN( u0_u14_u7_n170 ) );
  NAND2_X1 u0_u14_u7_U50 (.A2( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n147 ) , .A1( u0_u14_u7_n93 ) );
  NAND2_X1 u0_u14_u7_U51 (.A1( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n127 ) , .A2( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U52 (.A2( u0_u14_u7_n102 ) , .A1( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n133 ) );
  OR2_X1 u0_u14_u7_U53 (.ZN( u0_u14_u7_n126 ) , .A2( u0_u14_u7_n152 ) , .A1( u0_u14_u7_n156 ) );
  NAND2_X1 u0_u14_u7_U54 (.ZN( u0_u14_u7_n112 ) , .A2( u0_u14_u7_n96 ) , .A1( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U55 (.A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n128 ) , .A1( u0_u14_u7_n98 ) );
  INV_X1 u0_u14_u7_U56 (.A( u0_u14_u7_n150 ) , .ZN( u0_u14_u7_n164 ) );
  AND2_X1 u0_u14_u7_U57 (.ZN( u0_u14_u7_n134 ) , .A1( u0_u14_u7_n93 ) , .A2( u0_u14_u7_n98 ) );
  NAND2_X1 u0_u14_u7_U58 (.ZN( u0_u14_u7_n110 ) , .A1( u0_u14_u7_n95 ) , .A2( u0_u14_u7_n96 ) );
  NAND2_X1 u0_u14_u7_U59 (.A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n124 ) , .A1( u0_u14_u7_n96 ) );
  AOI211_X1 u0_u14_u7_U6 (.ZN( u0_u14_u7_n116 ) , .A( u0_u14_u7_n155 ) , .C1( u0_u14_u7_n161 ) , .C2( u0_u14_u7_n171 ) , .B( u0_u14_u7_n94 ) );
  NAND2_X1 u0_u14_u7_U60 (.ZN( u0_u14_u7_n132 ) , .A1( u0_u14_u7_n93 ) , .A2( u0_u14_u7_n96 ) );
  NAND2_X1 u0_u14_u7_U61 (.A2( u0_u14_u7_n103 ) , .ZN( u0_u14_u7_n131 ) , .A1( u0_u14_u7_n95 ) );
  NOR2_X1 u0_u14_u7_U62 (.A2( u0_u14_X_47 ) , .ZN( u0_u14_u7_n150 ) , .A1( u0_u14_u7_n163 ) );
  NOR2_X1 u0_u14_u7_U63 (.A2( u0_u14_X_43 ) , .A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n103 ) );
  NOR2_X1 u0_u14_u7_U64 (.A2( u0_u14_X_48 ) , .A1( u0_u14_u7_n166 ) , .ZN( u0_u14_u7_n95 ) );
  NOR2_X1 u0_u14_u7_U65 (.A2( u0_u14_X_44 ) , .A1( u0_u14_u7_n167 ) , .ZN( u0_u14_u7_n98 ) );
  NOR2_X1 u0_u14_u7_U66 (.A2( u0_u14_X_45 ) , .A1( u0_u14_X_48 ) , .ZN( u0_u14_u7_n99 ) );
  NOR2_X1 u0_u14_u7_U67 (.A2( u0_u14_X_46 ) , .A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n152 ) );
  AND2_X1 u0_u14_u7_U68 (.A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n156 ) , .A2( u0_u14_u7_n163 ) );
  NAND2_X1 u0_u14_u7_U69 (.A2( u0_u14_X_46 ) , .A1( u0_u14_X_47 ) , .ZN( u0_u14_u7_n125 ) );
  OAI222_X1 u0_u14_u7_U7 (.C2( u0_u14_u7_n101 ) , .B2( u0_u14_u7_n111 ) , .A1( u0_u14_u7_n113 ) , .C1( u0_u14_u7_n146 ) , .A2( u0_u14_u7_n162 ) , .B1( u0_u14_u7_n164 ) , .ZN( u0_u14_u7_n94 ) );
  AND2_X1 u0_u14_u7_U70 (.A2( u0_u14_X_43 ) , .A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n96 ) );
  AND2_X1 u0_u14_u7_U71 (.A2( u0_u14_X_45 ) , .A1( u0_u14_X_48 ) , .ZN( u0_u14_u7_n102 ) );
  AND2_X1 u0_u14_u7_U72 (.A1( u0_u14_X_48 ) , .A2( u0_u14_u7_n166 ) , .ZN( u0_u14_u7_n93 ) );
  INV_X1 u0_u14_u7_U73 (.A( u0_u14_X_46 ) , .ZN( u0_u14_u7_n163 ) );
  AND2_X1 u0_u14_u7_U74 (.A1( u0_u14_X_44 ) , .ZN( u0_u14_u7_n100 ) , .A2( u0_u14_u7_n167 ) );
  INV_X1 u0_u14_u7_U75 (.A( u0_u14_X_43 ) , .ZN( u0_u14_u7_n167 ) );
  INV_X1 u0_u14_u7_U76 (.A( u0_u14_X_45 ) , .ZN( u0_u14_u7_n166 ) );
  NAND4_X1 u0_u14_u7_U77 (.ZN( u0_out14_27 ) , .A4( u0_u14_u7_n118 ) , .A3( u0_u14_u7_n119 ) , .A2( u0_u14_u7_n120 ) , .A1( u0_u14_u7_n121 ) );
  OAI21_X1 u0_u14_u7_U78 (.ZN( u0_u14_u7_n121 ) , .B2( u0_u14_u7_n145 ) , .A( u0_u14_u7_n150 ) , .B1( u0_u14_u7_n174 ) );
  OAI21_X1 u0_u14_u7_U79 (.ZN( u0_u14_u7_n120 ) , .A( u0_u14_u7_n161 ) , .B2( u0_u14_u7_n170 ) , .B1( u0_u14_u7_n179 ) );
  INV_X1 u0_u14_u7_U8 (.A( u0_u14_u7_n133 ) , .ZN( u0_u14_u7_n176 ) );
  NAND4_X1 u0_u14_u7_U80 (.ZN( u0_out14_21 ) , .A4( u0_u14_u7_n157 ) , .A3( u0_u14_u7_n158 ) , .A2( u0_u14_u7_n159 ) , .A1( u0_u14_u7_n160 ) );
  OAI21_X1 u0_u14_u7_U81 (.B1( u0_u14_u7_n145 ) , .ZN( u0_u14_u7_n160 ) , .A( u0_u14_u7_n161 ) , .B2( u0_u14_u7_n177 ) );
  OAI21_X1 u0_u14_u7_U82 (.ZN( u0_u14_u7_n159 ) , .A( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n171 ) , .B1( u0_u14_u7_n174 ) );
  NAND4_X1 u0_u14_u7_U83 (.ZN( u0_out14_15 ) , .A4( u0_u14_u7_n142 ) , .A3( u0_u14_u7_n143 ) , .A2( u0_u14_u7_n144 ) , .A1( u0_u14_u7_n178 ) );
  OR2_X1 u0_u14_u7_U84 (.A2( u0_u14_u7_n125 ) , .A1( u0_u14_u7_n129 ) , .ZN( u0_u14_u7_n144 ) );
  AOI22_X1 u0_u14_u7_U85 (.A2( u0_u14_u7_n126 ) , .ZN( u0_u14_u7_n143 ) , .B2( u0_u14_u7_n165 ) , .B1( u0_u14_u7_n173 ) , .A1( u0_u14_u7_n174 ) );
  NAND4_X1 u0_u14_u7_U86 (.ZN( u0_out14_5 ) , .A4( u0_u14_u7_n108 ) , .A3( u0_u14_u7_n109 ) , .A1( u0_u14_u7_n116 ) , .A2( u0_u14_u7_n123 ) );
  AOI22_X1 u0_u14_u7_U87 (.ZN( u0_u14_u7_n109 ) , .A2( u0_u14_u7_n126 ) , .B2( u0_u14_u7_n145 ) , .B1( u0_u14_u7_n156 ) , .A1( u0_u14_u7_n171 ) );
  NOR4_X1 u0_u14_u7_U88 (.A4( u0_u14_u7_n104 ) , .A3( u0_u14_u7_n105 ) , .A2( u0_u14_u7_n106 ) , .A1( u0_u14_u7_n107 ) , .ZN( u0_u14_u7_n108 ) );
  NAND2_X1 u0_u14_u7_U89 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n148 ) , .A2( u0_u14_u7_n95 ) );
  OAI221_X1 u0_u14_u7_U9 (.C1( u0_u14_u7_n101 ) , .C2( u0_u14_u7_n147 ) , .ZN( u0_u14_u7_n155 ) , .B2( u0_u14_u7_n162 ) , .A( u0_u14_u7_n91 ) , .B1( u0_u14_u7_n92 ) );
  NAND2_X1 u0_u14_u7_U90 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n113 ) , .A2( u0_u14_u7_n93 ) );
  NAND2_X1 u0_u14_u7_U91 (.A1( u0_u14_u7_n100 ) , .ZN( u0_u14_u7_n138 ) , .A2( u0_u14_u7_n99 ) );
  NAND2_X1 u0_u14_u7_U92 (.A1( u0_u14_u7_n100 ) , .A2( u0_u14_u7_n102 ) , .ZN( u0_u14_u7_n129 ) );
  OAI211_X1 u0_u14_u7_U93 (.B( u0_u14_u7_n122 ) , .A( u0_u14_u7_n123 ) , .C2( u0_u14_u7_n124 ) , .ZN( u0_u14_u7_n154 ) , .C1( u0_u14_u7_n162 ) );
  AOI222_X1 u0_u14_u7_U94 (.ZN( u0_u14_u7_n122 ) , .C2( u0_u14_u7_n126 ) , .C1( u0_u14_u7_n145 ) , .B1( u0_u14_u7_n161 ) , .A2( u0_u14_u7_n165 ) , .B2( u0_u14_u7_n170 ) , .A1( u0_u14_u7_n176 ) );
  NAND3_X1 u0_u14_u7_U95 (.A3( u0_u14_u7_n146 ) , .A2( u0_u14_u7_n147 ) , .A1( u0_u14_u7_n148 ) , .ZN( u0_u14_u7_n151 ) );
  NAND3_X1 u0_u14_u7_U96 (.A3( u0_u14_u7_n131 ) , .A2( u0_u14_u7_n132 ) , .A1( u0_u14_u7_n133 ) , .ZN( u0_u14_u7_n135 ) );
  XOR2_X1 u0_u3_U1 (.B( u0_K4_9 ) , .A( u0_R2_6 ) , .Z( u0_u3_X_9 ) );
  XOR2_X1 u0_u3_U16 (.B( u0_K4_3 ) , .A( u0_R2_2 ) , .Z( u0_u3_X_3 ) );
  XOR2_X1 u0_u3_U2 (.B( u0_K4_8 ) , .A( u0_R2_5 ) , .Z( u0_u3_X_8 ) );
  XOR2_X1 u0_u3_U27 (.B( u0_K4_2 ) , .A( u0_R2_1 ) , .Z( u0_u3_X_2 ) );
  XOR2_X1 u0_u3_U3 (.B( u0_K4_7 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_7 ) );
  XOR2_X1 u0_u3_U33 (.B( u0_K4_24 ) , .A( u0_R2_17 ) , .Z( u0_u3_X_24 ) );
  XOR2_X1 u0_u3_U34 (.B( u0_K4_23 ) , .A( u0_R2_16 ) , .Z( u0_u3_X_23 ) );
  XOR2_X1 u0_u3_U35 (.B( u0_K4_22 ) , .A( u0_R2_15 ) , .Z( u0_u3_X_22 ) );
  XOR2_X1 u0_u3_U36 (.B( u0_K4_21 ) , .A( u0_R2_14 ) , .Z( u0_u3_X_21 ) );
  XOR2_X1 u0_u3_U37 (.B( u0_K4_20 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_20 ) );
  XOR2_X1 u0_u3_U38 (.B( u0_K4_1 ) , .A( u0_R2_32 ) , .Z( u0_u3_X_1 ) );
  XOR2_X1 u0_u3_U39 (.B( u0_K4_19 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_19 ) );
  XOR2_X1 u0_u3_U4 (.B( u0_K4_6 ) , .A( u0_R2_5 ) , .Z( u0_u3_X_6 ) );
  XOR2_X1 u0_u3_U40 (.B( u0_K4_18 ) , .A( u0_R2_13 ) , .Z( u0_u3_X_18 ) );
  XOR2_X1 u0_u3_U41 (.B( u0_K4_17 ) , .A( u0_R2_12 ) , .Z( u0_u3_X_17 ) );
  XOR2_X1 u0_u3_U42 (.B( u0_K4_16 ) , .A( u0_R2_11 ) , .Z( u0_u3_X_16 ) );
  XOR2_X1 u0_u3_U43 (.B( u0_K4_15 ) , .A( u0_R2_10 ) , .Z( u0_u3_X_15 ) );
  XOR2_X1 u0_u3_U44 (.B( u0_K4_14 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_14 ) );
  XOR2_X1 u0_u3_U45 (.B( u0_K4_13 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_13 ) );
  XOR2_X1 u0_u3_U46 (.B( u0_K4_12 ) , .A( u0_R2_9 ) , .Z( u0_u3_X_12 ) );
  XOR2_X1 u0_u3_U47 (.B( u0_K4_11 ) , .A( u0_R2_8 ) , .Z( u0_u3_X_11 ) );
  XOR2_X1 u0_u3_U48 (.B( u0_K4_10 ) , .A( u0_R2_7 ) , .Z( u0_u3_X_10 ) );
  XOR2_X1 u0_u3_U5 (.B( u0_K4_5 ) , .A( u0_R2_4 ) , .Z( u0_u3_X_5 ) );
  XOR2_X1 u0_u3_U6 (.B( u0_K4_4 ) , .A( u0_R2_3 ) , .Z( u0_u3_X_4 ) );
  AND2_X1 u0_u3_u0_U10 (.A1( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n143 ) , .A2( u0_u3_u0_n152 ) );
  AND2_X1 u0_u3_u0_U11 (.ZN( u0_u3_u0_n109 ) , .A1( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n142 ) );
  AND2_X1 u0_u3_u0_U12 (.A2( u0_u3_u0_n131 ) , .A1( u0_u3_u0_n132 ) , .ZN( u0_u3_u0_n153 ) );
  AND2_X1 u0_u3_u0_U13 (.A1( u0_u3_u0_n110 ) , .A2( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U14 (.A( u0_u3_u0_n145 ) , .ZN( u0_u3_u0_n175 ) );
  NOR2_X1 u0_u3_u0_U15 (.A2( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n149 ) , .A1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U16 (.B1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n134 ) , .A( u0_u3_u0_n167 ) , .B2( u0_u3_u0_n95 ) );
  OAI22_X1 u0_u3_u0_U17 (.B1( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n149 ) , .A2( u0_u3_u0_n92 ) , .ZN( u0_u3_u0_n93 ) );
  AND3_X1 u0_u3_u0_U18 (.A3( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n127 ) , .A1( u0_u3_u0_n150 ) , .ZN( u0_u3_u0_n92 ) );
  OAI22_X1 u0_u3_u0_U19 (.B1( u0_u3_u0_n127 ) , .ZN( u0_u3_u0_n128 ) , .A1( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n148 ) , .B2( u0_u3_u0_n149 ) );
  NOR2_X1 u0_u3_u0_U20 (.A1( u0_u3_u0_n165 ) , .A2( u0_u3_u0_n166 ) , .ZN( u0_u3_u0_n97 ) );
  AOI22_X1 u0_u3_u0_U21 (.B2( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n112 ) , .ZN( u0_u3_u0_n113 ) , .B1( u0_u3_u0_n120 ) , .A1( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U22 (.A2( u0_u3_u0_n104 ) , .A1( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n151 ) );
  INV_X1 u0_u3_u0_U23 (.A( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U24 (.A( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n160 ) );
  NAND2_X1 u0_u3_u0_U25 (.A2( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n133 ) , .A1( u0_u3_u0_n94 ) );
  NAND2_X1 u0_u3_u0_U26 (.ZN( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n94 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U27 (.ZN( u0_u3_u0_n106 ) , .B1( u0_u3_u0_n109 ) , .B2( u0_u3_u0_n143 ) , .A( u0_u3_u0_n146 ) );
  AOI21_X1 u0_u3_u0_U28 (.B1( u0_u3_u0_n129 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n98 ) );
  NAND2_X1 u0_u3_u0_U29 (.A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n116 ) , .A1( u0_u3_u0_n94 ) );
  INV_X1 u0_u3_u0_U3 (.A( u0_u3_u0_n115 ) , .ZN( u0_u3_u0_n168 ) );
  NOR2_X1 u0_u3_u0_U30 (.A1( u0_u3_u0_n122 ) , .ZN( u0_u3_u0_n145 ) , .A2( u0_u3_u0_n169 ) );
  OAI221_X1 u0_u3_u0_U31 (.C1( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n122 ) , .B1( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n143 ) , .C2( u0_u3_u0_n149 ) , .A( u0_u3_u0_n174 ) );
  AOI211_X1 u0_u3_u0_U32 (.B( u0_u3_u0_n117 ) , .A( u0_u3_u0_n118 ) , .C2( u0_u3_u0_n119 ) , .C1( u0_u3_u0_n120 ) , .ZN( u0_u3_u0_n121 ) );
  NAND2_X1 u0_u3_u0_U33 (.A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n96 ) );
  NAND2_X1 u0_u3_u0_U34 (.A1( u0_u3_u0_n102 ) , .A2( u0_u3_u0_n105 ) , .ZN( u0_u3_u0_n127 ) );
  NAND2_X1 u0_u3_u0_U35 (.A1( u0_u3_u0_n103 ) , .A2( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n152 ) );
  INV_X1 u0_u3_u0_U36 (.A( u0_u3_u0_n140 ) , .ZN( u0_u3_u0_n162 ) );
  NAND2_X1 u0_u3_u0_U37 (.A2( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n141 ) );
  NAND2_X1 u0_u3_u0_U38 (.ZN( u0_u3_u0_n114 ) , .A2( u0_u3_u0_n94 ) , .A1( u0_u3_u0_n95 ) );
  NAND2_X1 u0_u3_u0_U39 (.A1( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n132 ) , .A2( u0_u3_u0_n96 ) );
  AOI21_X1 u0_u3_u0_U4 (.B1( u0_u3_u0_n116 ) , .ZN( u0_u3_u0_n117 ) , .B2( u0_u3_u0_n131 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U40 (.ZN( u0_u3_u0_n174 ) , .A( u0_u3_u0_n90 ) );
  OAI222_X1 u0_u3_u0_U41 (.C1( u0_u3_u0_n110 ) , .A1( u0_u3_u0_n127 ) , .B2( u0_u3_u0_n130 ) , .B1( u0_u3_u0_n146 ) , .A2( u0_u3_u0_n160 ) , .C2( u0_u3_u0_n163 ) , .ZN( u0_u3_u0_n90 ) );
  OR3_X1 u0_u3_u0_U42 (.A3( u0_u3_u0_n154 ) , .A2( u0_u3_u0_n155 ) , .A1( u0_u3_u0_n156 ) , .ZN( u0_u3_u0_n157 ) );
  AOI21_X1 u0_u3_u0_U43 (.A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n147 ) , .B1( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n156 ) );
  AOI21_X1 u0_u3_u0_U44 (.B2( u0_u3_u0_n152 ) , .B1( u0_u3_u0_n153 ) , .ZN( u0_u3_u0_n154 ) , .A( u0_u3_u0_n160 ) );
  AOI21_X1 u0_u3_u0_U45 (.A( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n150 ) , .B1( u0_u3_u0_n151 ) , .ZN( u0_u3_u0_n155 ) );
  INV_X1 u0_u3_u0_U46 (.A( u0_u3_u0_n101 ) , .ZN( u0_u3_u0_n173 ) );
  OAI211_X1 u0_u3_u0_U47 (.B( u0_u3_u0_n100 ) , .ZN( u0_u3_u0_n101 ) , .C2( u0_u3_u0_n142 ) , .C1( u0_u3_u0_n163 ) , .A( u0_u3_u0_n171 ) );
  INV_X1 u0_u3_u0_U48 (.ZN( u0_u3_u0_n171 ) , .A( u0_u3_u0_n93 ) );
  AOI211_X1 u0_u3_u0_U49 (.ZN( u0_u3_u0_n100 ) , .C1( u0_u3_u0_n120 ) , .A( u0_u3_u0_n125 ) , .B( u0_u3_u0_n98 ) , .C2( u0_u3_u0_n99 ) );
  AOI21_X1 u0_u3_u0_U5 (.B2( u0_u3_u0_n133 ) , .ZN( u0_u3_u0_n136 ) , .B1( u0_u3_u0_n153 ) , .A( u0_u3_u0_n160 ) );
  NOR2_X1 u0_u3_u0_U50 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n120 ) );
  NOR2_X1 u0_u3_u0_U51 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n96 ) );
  NOR2_X1 u0_u3_u0_U52 (.A2( u0_u3_X_6 ) , .ZN( u0_u3_u0_n102 ) , .A1( u0_u3_u0_n164 ) );
  NOR2_X1 u0_u3_u0_U53 (.A2( u0_u3_X_1 ) , .ZN( u0_u3_u0_n103 ) , .A1( u0_u3_u0_n165 ) );
  NAND2_X1 u0_u3_u0_U54 (.A2( u0_u3_X_4 ) , .A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n146 ) );
  NOR2_X1 u0_u3_u0_U55 (.A2( u0_u3_X_5 ) , .ZN( u0_u3_u0_n138 ) , .A1( u0_u3_u0_n161 ) );
  NAND2_X1 u0_u3_u0_U56 (.A1( u0_u3_X_5 ) , .ZN( u0_u3_u0_n140 ) , .A2( u0_u3_u0_n161 ) );
  AND2_X1 u0_u3_u0_U57 (.A2( u0_u3_X_3 ) , .A1( u0_u3_X_6 ) , .ZN( u0_u3_u0_n104 ) );
  AND2_X1 u0_u3_u0_U58 (.A1( u0_u3_X_6 ) , .A2( u0_u3_u0_n164 ) , .ZN( u0_u3_u0_n95 ) );
  INV_X1 u0_u3_u0_U59 (.A( u0_u3_X_4 ) , .ZN( u0_u3_u0_n161 ) );
  NOR2_X1 u0_u3_u0_U6 (.A1( u0_u3_u0_n110 ) , .ZN( u0_u3_u0_n125 ) , .A2( u0_u3_u0_n160 ) );
  INV_X1 u0_u3_u0_U60 (.A( u0_u3_X_1 ) , .ZN( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U61 (.A( u0_u3_X_3 ) , .ZN( u0_u3_u0_n164 ) );
  INV_X1 u0_u3_u0_U62 (.A( u0_u3_u0_n128 ) , .ZN( u0_u3_u0_n170 ) );
  AOI211_X1 u0_u3_u0_U63 (.B( u0_u3_u0_n135 ) , .A( u0_u3_u0_n136 ) , .C2( u0_u3_u0_n137 ) , .C1( u0_u3_u0_n138 ) , .ZN( u0_u3_u0_n139 ) );
  OR4_X1 u0_u3_u0_U64 (.ZN( u0_out3_31 ) , .A4( u0_u3_u0_n157 ) , .A2( u0_u3_u0_n158 ) , .A1( u0_u3_u0_n159 ) , .A3( u0_u3_u0_n175 ) );
  AOI21_X1 u0_u3_u0_U65 (.A( u0_u3_u0_n140 ) , .B2( u0_u3_u0_n141 ) , .B1( u0_u3_u0_n142 ) , .ZN( u0_u3_u0_n159 ) );
  OR4_X1 u0_u3_u0_U66 (.ZN( u0_out3_17 ) , .A4( u0_u3_u0_n124 ) , .A2( u0_u3_u0_n125 ) , .A1( u0_u3_u0_n126 ) , .A3( u0_u3_u0_n172 ) );
  AOI21_X1 u0_u3_u0_U67 (.B2( u0_u3_u0_n109 ) , .ZN( u0_u3_u0_n126 ) , .B1( u0_u3_u0_n130 ) , .A( u0_u3_u0_n163 ) );
  INV_X1 u0_u3_u0_U68 (.A( u0_u3_u0_n113 ) , .ZN( u0_u3_u0_n172 ) );
  INV_X1 u0_u3_u0_U69 (.ZN( u0_u3_u0_n176 ) , .A( u0_u3_u0_n91 ) );
  OAI21_X1 u0_u3_u0_U7 (.B1( u0_u3_u0_n152 ) , .B2( u0_u3_u0_n160 ) , .A( u0_u3_u0_n174 ) , .ZN( u0_u3_u0_n91 ) );
  AOI211_X1 u0_u3_u0_U70 (.B( u0_u3_u0_n106 ) , .A( u0_u3_u0_n107 ) , .ZN( u0_u3_u0_n108 ) , .C2( u0_u3_u0_n115 ) , .C1( u0_u3_u0_n162 ) );
  AOI21_X1 u0_u3_u0_U71 (.B2( u0_u3_u0_n143 ) , .B1( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n158 ) , .A( u0_u3_u0_n163 ) );
  AOI21_X1 u0_u3_u0_U72 (.ZN( u0_u3_u0_n118 ) , .B2( u0_u3_u0_n144 ) , .A( u0_u3_u0_n146 ) , .B1( u0_u3_u0_n168 ) );
  INV_X1 u0_u3_u0_U73 (.A( u0_u3_u0_n144 ) , .ZN( u0_u3_u0_n167 ) );
  NOR2_X1 u0_u3_u0_U74 (.A2( u0_u3_X_1 ) , .A1( u0_u3_X_2 ) , .ZN( u0_u3_u0_n94 ) );
  NOR2_X1 u0_u3_u0_U75 (.A2( u0_u3_X_2 ) , .ZN( u0_u3_u0_n105 ) , .A1( u0_u3_u0_n166 ) );
  INV_X1 u0_u3_u0_U76 (.A( u0_u3_X_2 ) , .ZN( u0_u3_u0_n165 ) );
  OR2_X1 u0_u3_u0_U77 (.A2( u0_u3_u0_n129 ) , .A1( u0_u3_u0_n146 ) , .ZN( u0_u3_u0_n88 ) );
  OR2_X1 u0_u3_u0_U78 (.A1( u0_u3_u0_n123 ) , .A2( u0_u3_u0_n149 ) , .ZN( u0_u3_u0_n89 ) );
  NAND3_X1 u0_u3_u0_U79 (.ZN( u0_u3_u0_n124 ) , .A3( u0_u3_u0_n145 ) , .A1( u0_u3_u0_n88 ) , .A2( u0_u3_u0_n89 ) );
  AND2_X1 u0_u3_u0_U8 (.A1( u0_u3_u0_n116 ) , .A2( u0_u3_u0_n123 ) , .ZN( u0_u3_u0_n148 ) );
  AND3_X1 u0_u3_u0_U80 (.A2( u0_u3_u0_n114 ) , .ZN( u0_u3_u0_n129 ) , .A3( u0_u3_u0_n132 ) , .A1( u0_u3_u0_n150 ) );
  NAND2_X1 u0_u3_u0_U81 (.A2( u0_u3_u0_n103 ) , .ZN( u0_u3_u0_n123 ) , .A1( u0_u3_u0_n95 ) );
  AOI21_X1 u0_u3_u0_U82 (.B1( u0_u3_u0_n134 ) , .ZN( u0_u3_u0_n135 ) , .A( u0_u3_u0_n146 ) , .B2( u0_u3_u0_n168 ) );
  OAI22_X1 u0_u3_u0_U83 (.ZN( u0_u3_u0_n107 ) , .A2( u0_u3_u0_n134 ) , .B1( u0_u3_u0_n148 ) , .A1( u0_u3_u0_n149 ) , .B2( u0_u3_u0_n163 ) );
  NAND2_X1 u0_u3_u0_U84 (.ZN( u0_u3_u0_n112 ) , .A2( u0_u3_u0_n134 ) , .A1( u0_u3_u0_n147 ) );
  INV_X1 u0_u3_u0_U85 (.A( u0_u3_u0_n121 ) , .ZN( u0_u3_u0_n169 ) );
  NAND2_X1 u0_u3_u0_U86 (.ZN( u0_u3_u0_n150 ) , .A1( u0_u3_u0_n95 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U87 (.A1( u0_u3_u0_n102 ) , .ZN( u0_u3_u0_n131 ) , .A2( u0_u3_u0_n97 ) );
  NAND3_X1 u0_u3_u0_U88 (.ZN( u0_out3_23 ) , .A3( u0_u3_u0_n139 ) , .A1( u0_u3_u0_n170 ) , .A2( u0_u3_u0_n173 ) );
  NAND3_X1 u0_u3_u0_U89 (.A3( u0_u3_u0_n129 ) , .A2( u0_u3_u0_n130 ) , .ZN( u0_u3_u0_n137 ) , .A1( u0_u3_u0_n152 ) );
  NAND2_X1 u0_u3_u0_U9 (.ZN( u0_u3_u0_n115 ) , .A1( u0_u3_u0_n141 ) , .A2( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U90 (.ZN( u0_u3_u0_n119 ) , .A3( u0_u3_u0_n134 ) , .A2( u0_u3_u0_n141 ) , .A1( u0_u3_u0_n150 ) );
  NAND3_X1 u0_u3_u0_U91 (.ZN( u0_u3_u0_n111 ) , .A2( u0_u3_u0_n116 ) , .A3( u0_u3_u0_n142 ) , .A1( u0_u3_u0_n151 ) );
  NAND3_X1 u0_u3_u0_U92 (.ZN( u0_out3_9 ) , .A3( u0_u3_u0_n108 ) , .A2( u0_u3_u0_n173 ) , .A1( u0_u3_u0_n176 ) );
  NAND3_X1 u0_u3_u0_U93 (.A2( u0_u3_u0_n130 ) , .A1( u0_u3_u0_n134 ) , .A3( u0_u3_u0_n148 ) , .ZN( u0_u3_u0_n99 ) );
  NAND2_X1 u0_u3_u0_U94 (.A1( u0_u3_u0_n104 ) , .ZN( u0_u3_u0_n130 ) , .A2( u0_u3_u0_n97 ) );
  NAND2_X1 u0_u3_u0_U95 (.ZN( u0_u3_u0_n144 ) , .A1( u0_u3_u0_n96 ) , .A2( u0_u3_u0_n97 ) );
  NOR2_X1 u0_u3_u1_U10 (.A1( u0_u3_u1_n112 ) , .A2( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n118 ) );
  NAND3_X1 u0_u3_u1_U100 (.ZN( u0_u3_u1_n113 ) , .A1( u0_u3_u1_n120 ) , .A3( u0_u3_u1_n133 ) , .A2( u0_u3_u1_n155 ) );
  OAI21_X1 u0_u3_u1_U11 (.ZN( u0_u3_u1_n101 ) , .B1( u0_u3_u1_n141 ) , .A( u0_u3_u1_n146 ) , .B2( u0_u3_u1_n183 ) );
  AOI21_X1 u0_u3_u1_U12 (.B2( u0_u3_u1_n155 ) , .B1( u0_u3_u1_n156 ) , .ZN( u0_u3_u1_n157 ) , .A( u0_u3_u1_n174 ) );
  NAND2_X1 u0_u3_u1_U13 (.ZN( u0_u3_u1_n140 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n155 ) );
  NAND2_X1 u0_u3_u1_U14 (.A1( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n153 ) );
  INV_X1 u0_u3_u1_U15 (.A( u0_u3_u1_n139 ) , .ZN( u0_u3_u1_n174 ) );
  OR4_X1 u0_u3_u1_U16 (.A4( u0_u3_u1_n106 ) , .A3( u0_u3_u1_n107 ) , .ZN( u0_u3_u1_n108 ) , .A1( u0_u3_u1_n117 ) , .A2( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U17 (.ZN( u0_u3_u1_n106 ) , .A( u0_u3_u1_n112 ) , .B1( u0_u3_u1_n154 ) , .B2( u0_u3_u1_n156 ) );
  INV_X1 u0_u3_u1_U18 (.A( u0_u3_u1_n101 ) , .ZN( u0_u3_u1_n184 ) );
  AOI21_X1 u0_u3_u1_U19 (.ZN( u0_u3_u1_n107 ) , .B1( u0_u3_u1_n134 ) , .B2( u0_u3_u1_n149 ) , .A( u0_u3_u1_n174 ) );
  INV_X1 u0_u3_u1_U20 (.A( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n171 ) );
  NAND2_X1 u0_u3_u1_U21 (.ZN( u0_u3_u1_n141 ) , .A1( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n156 ) );
  AND2_X1 u0_u3_u1_U22 (.A1( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n161 ) );
  NAND2_X1 u0_u3_u1_U23 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n116 ) , .ZN( u0_u3_u1_n148 ) );
  NAND2_X1 u0_u3_u1_U24 (.A2( u0_u3_u1_n133 ) , .A1( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n159 ) );
  NAND2_X1 u0_u3_u1_U25 (.A2( u0_u3_u1_n115 ) , .A1( u0_u3_u1_n120 ) , .ZN( u0_u3_u1_n132 ) );
  INV_X1 u0_u3_u1_U26 (.A( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n178 ) );
  INV_X1 u0_u3_u1_U27 (.A( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n183 ) );
  AND2_X1 u0_u3_u1_U28 (.A1( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n149 ) );
  INV_X1 u0_u3_u1_U29 (.A( u0_u3_u1_n131 ) , .ZN( u0_u3_u1_n180 ) );
  INV_X1 u0_u3_u1_U3 (.A( u0_u3_u1_n159 ) , .ZN( u0_u3_u1_n182 ) );
  AOI221_X1 u0_u3_u1_U30 (.B1( u0_u3_u1_n140 ) , .ZN( u0_u3_u1_n167 ) , .B2( u0_u3_u1_n172 ) , .C2( u0_u3_u1_n175 ) , .C1( u0_u3_u1_n178 ) , .A( u0_u3_u1_n188 ) );
  INV_X1 u0_u3_u1_U31 (.ZN( u0_u3_u1_n188 ) , .A( u0_u3_u1_n97 ) );
  AOI211_X1 u0_u3_u1_U32 (.A( u0_u3_u1_n118 ) , .C1( u0_u3_u1_n132 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n96 ) , .ZN( u0_u3_u1_n97 ) );
  AOI21_X1 u0_u3_u1_U33 (.B2( u0_u3_u1_n121 ) , .B1( u0_u3_u1_n135 ) , .A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n96 ) );
  OAI221_X1 u0_u3_u1_U34 (.A( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n138 ) , .B2( u0_u3_u1_n152 ) , .C1( u0_u3_u1_n174 ) , .B1( u0_u3_u1_n187 ) );
  INV_X1 u0_u3_u1_U35 (.A( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n187 ) );
  AOI211_X1 u0_u3_u1_U36 (.B( u0_u3_u1_n117 ) , .A( u0_u3_u1_n118 ) , .ZN( u0_u3_u1_n119 ) , .C2( u0_u3_u1_n146 ) , .C1( u0_u3_u1_n159 ) );
  NOR2_X1 u0_u3_u1_U37 (.A1( u0_u3_u1_n168 ) , .A2( u0_u3_u1_n176 ) , .ZN( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U38 (.A1( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n146 ) , .A2( u0_u3_u1_n160 ) );
  NAND2_X1 u0_u3_u1_U39 (.A2( u0_u3_u1_n112 ) , .ZN( u0_u3_u1_n139 ) , .A1( u0_u3_u1_n152 ) );
  AOI221_X1 u0_u3_u1_U4 (.A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .C1( u0_u3_u1_n140 ) , .B2( u0_u3_u1_n141 ) , .ZN( u0_u3_u1_n142 ) , .B1( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U40 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n156 ) , .A2( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U41 (.ZN( u0_u3_u1_n117 ) , .A1( u0_u3_u1_n121 ) , .A2( u0_u3_u1_n160 ) );
  OAI21_X1 u0_u3_u1_U42 (.B2( u0_u3_u1_n123 ) , .ZN( u0_u3_u1_n145 ) , .B1( u0_u3_u1_n160 ) , .A( u0_u3_u1_n185 ) );
  INV_X1 u0_u3_u1_U43 (.A( u0_u3_u1_n122 ) , .ZN( u0_u3_u1_n185 ) );
  AOI21_X1 u0_u3_u1_U44 (.B2( u0_u3_u1_n120 ) , .B1( u0_u3_u1_n121 ) , .ZN( u0_u3_u1_n122 ) , .A( u0_u3_u1_n128 ) );
  AOI21_X1 u0_u3_u1_U45 (.A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n129 ) , .ZN( u0_u3_u1_n130 ) , .B1( u0_u3_u1_n150 ) );
  NAND2_X1 u0_u3_u1_U46 (.ZN( u0_u3_u1_n112 ) , .A1( u0_u3_u1_n169 ) , .A2( u0_u3_u1_n170 ) );
  NAND2_X1 u0_u3_u1_U47 (.ZN( u0_u3_u1_n129 ) , .A2( u0_u3_u1_n95 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U48 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n154 ) , .A2( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U49 (.A2( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n135 ) , .A1( u0_u3_u1_n99 ) );
  AOI211_X1 u0_u3_u1_U5 (.ZN( u0_u3_u1_n124 ) , .A( u0_u3_u1_n138 ) , .C2( u0_u3_u1_n139 ) , .B( u0_u3_u1_n145 ) , .C1( u0_u3_u1_n147 ) );
  AOI21_X1 u0_u3_u1_U50 (.A( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n153 ) , .B1( u0_u3_u1_n154 ) , .ZN( u0_u3_u1_n158 ) );
  INV_X1 u0_u3_u1_U51 (.A( u0_u3_u1_n160 ) , .ZN( u0_u3_u1_n175 ) );
  NAND2_X1 u0_u3_u1_U52 (.A1( u0_u3_u1_n100 ) , .ZN( u0_u3_u1_n116 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U53 (.A1( u0_u3_u1_n102 ) , .ZN( u0_u3_u1_n131 ) , .A2( u0_u3_u1_n95 ) );
  NAND2_X1 u0_u3_u1_U54 (.A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n121 ) , .A1( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U55 (.A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n153 ) , .A2( u0_u3_u1_n98 ) );
  NAND2_X1 u0_u3_u1_U56 (.A2( u0_u3_u1_n104 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n133 ) );
  NAND2_X1 u0_u3_u1_U57 (.ZN( u0_u3_u1_n150 ) , .A2( u0_u3_u1_n98 ) , .A1( u0_u3_u1_n99 ) );
  NAND2_X1 u0_u3_u1_U58 (.A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n155 ) , .A2( u0_u3_u1_n95 ) );
  OAI21_X1 u0_u3_u1_U59 (.ZN( u0_u3_u1_n109 ) , .B1( u0_u3_u1_n129 ) , .B2( u0_u3_u1_n160 ) , .A( u0_u3_u1_n167 ) );
  AOI22_X1 u0_u3_u1_U6 (.B2( u0_u3_u1_n113 ) , .A2( u0_u3_u1_n114 ) , .ZN( u0_u3_u1_n125 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  NAND2_X1 u0_u3_u1_U60 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n120 ) );
  NAND2_X1 u0_u3_u1_U61 (.A1( u0_u3_u1_n102 ) , .A2( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n115 ) );
  NAND2_X1 u0_u3_u1_U62 (.A2( u0_u3_u1_n100 ) , .A1( u0_u3_u1_n104 ) , .ZN( u0_u3_u1_n151 ) );
  NAND2_X1 u0_u3_u1_U63 (.A2( u0_u3_u1_n103 ) , .A1( u0_u3_u1_n105 ) , .ZN( u0_u3_u1_n161 ) );
  INV_X1 u0_u3_u1_U64 (.A( u0_u3_u1_n152 ) , .ZN( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U65 (.A( u0_u3_u1_n128 ) , .ZN( u0_u3_u1_n172 ) );
  NAND2_X1 u0_u3_u1_U66 (.A2( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n103 ) , .ZN( u0_u3_u1_n123 ) );
  AOI211_X1 u0_u3_u1_U67 (.B( u0_u3_u1_n162 ) , .A( u0_u3_u1_n163 ) , .C2( u0_u3_u1_n164 ) , .ZN( u0_u3_u1_n165 ) , .C1( u0_u3_u1_n171 ) );
  AOI21_X1 u0_u3_u1_U68 (.A( u0_u3_u1_n160 ) , .B2( u0_u3_u1_n161 ) , .ZN( u0_u3_u1_n162 ) , .B1( u0_u3_u1_n182 ) );
  OR2_X1 u0_u3_u1_U69 (.A2( u0_u3_u1_n157 ) , .A1( u0_u3_u1_n158 ) , .ZN( u0_u3_u1_n163 ) );
  NAND2_X1 u0_u3_u1_U7 (.ZN( u0_u3_u1_n114 ) , .A1( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n156 ) );
  NOR2_X1 u0_u3_u1_U70 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n95 ) );
  NOR2_X1 u0_u3_u1_U71 (.A1( u0_u3_X_12 ) , .A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n100 ) );
  NOR2_X1 u0_u3_u1_U72 (.A2( u0_u3_X_8 ) , .A1( u0_u3_u1_n177 ) , .ZN( u0_u3_u1_n99 ) );
  NOR2_X1 u0_u3_u1_U73 (.A2( u0_u3_X_12 ) , .ZN( u0_u3_u1_n102 ) , .A1( u0_u3_u1_n176 ) );
  NOR2_X1 u0_u3_u1_U74 (.A2( u0_u3_X_9 ) , .ZN( u0_u3_u1_n105 ) , .A1( u0_u3_u1_n168 ) );
  NAND2_X1 u0_u3_u1_U75 (.A1( u0_u3_X_10 ) , .ZN( u0_u3_u1_n160 ) , .A2( u0_u3_u1_n169 ) );
  NAND2_X1 u0_u3_u1_U76 (.A2( u0_u3_X_10 ) , .A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n152 ) );
  NAND2_X1 u0_u3_u1_U77 (.A1( u0_u3_X_11 ) , .ZN( u0_u3_u1_n128 ) , .A2( u0_u3_u1_n170 ) );
  AND2_X1 u0_u3_u1_U78 (.A2( u0_u3_X_7 ) , .A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n104 ) );
  AND2_X1 u0_u3_u1_U79 (.A1( u0_u3_X_8 ) , .ZN( u0_u3_u1_n103 ) , .A2( u0_u3_u1_n177 ) );
  AOI22_X1 u0_u3_u1_U8 (.B2( u0_u3_u1_n136 ) , .A2( u0_u3_u1_n137 ) , .ZN( u0_u3_u1_n143 ) , .A1( u0_u3_u1_n171 ) , .B1( u0_u3_u1_n173 ) );
  INV_X1 u0_u3_u1_U80 (.A( u0_u3_X_10 ) , .ZN( u0_u3_u1_n170 ) );
  INV_X1 u0_u3_u1_U81 (.A( u0_u3_X_9 ) , .ZN( u0_u3_u1_n176 ) );
  INV_X1 u0_u3_u1_U82 (.A( u0_u3_X_11 ) , .ZN( u0_u3_u1_n169 ) );
  INV_X1 u0_u3_u1_U83 (.A( u0_u3_X_12 ) , .ZN( u0_u3_u1_n168 ) );
  INV_X1 u0_u3_u1_U84 (.A( u0_u3_X_7 ) , .ZN( u0_u3_u1_n177 ) );
  NAND4_X1 u0_u3_u1_U85 (.ZN( u0_out3_28 ) , .A4( u0_u3_u1_n124 ) , .A3( u0_u3_u1_n125 ) , .A2( u0_u3_u1_n126 ) , .A1( u0_u3_u1_n127 ) );
  OAI21_X1 u0_u3_u1_U86 (.ZN( u0_u3_u1_n127 ) , .B2( u0_u3_u1_n139 ) , .B1( u0_u3_u1_n175 ) , .A( u0_u3_u1_n183 ) );
  OAI21_X1 u0_u3_u1_U87 (.ZN( u0_u3_u1_n126 ) , .B2( u0_u3_u1_n140 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n178 ) );
  NAND4_X1 u0_u3_u1_U88 (.ZN( u0_out3_18 ) , .A4( u0_u3_u1_n165 ) , .A3( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n167 ) , .A2( u0_u3_u1_n186 ) );
  AOI22_X1 u0_u3_u1_U89 (.B2( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n147 ) , .A2( u0_u3_u1_n148 ) , .ZN( u0_u3_u1_n166 ) , .A1( u0_u3_u1_n172 ) );
  INV_X1 u0_u3_u1_U9 (.A( u0_u3_u1_n147 ) , .ZN( u0_u3_u1_n181 ) );
  INV_X1 u0_u3_u1_U90 (.A( u0_u3_u1_n145 ) , .ZN( u0_u3_u1_n186 ) );
  NAND4_X1 u0_u3_u1_U91 (.ZN( u0_out3_2 ) , .A4( u0_u3_u1_n142 ) , .A3( u0_u3_u1_n143 ) , .A2( u0_u3_u1_n144 ) , .A1( u0_u3_u1_n179 ) );
  INV_X1 u0_u3_u1_U92 (.A( u0_u3_u1_n130 ) , .ZN( u0_u3_u1_n179 ) );
  OAI21_X1 u0_u3_u1_U93 (.B2( u0_u3_u1_n132 ) , .ZN( u0_u3_u1_n144 ) , .A( u0_u3_u1_n146 ) , .B1( u0_u3_u1_n180 ) );
  OR4_X1 u0_u3_u1_U94 (.ZN( u0_out3_13 ) , .A4( u0_u3_u1_n108 ) , .A3( u0_u3_u1_n109 ) , .A2( u0_u3_u1_n110 ) , .A1( u0_u3_u1_n111 ) );
  AOI21_X1 u0_u3_u1_U95 (.ZN( u0_u3_u1_n111 ) , .A( u0_u3_u1_n128 ) , .B2( u0_u3_u1_n131 ) , .B1( u0_u3_u1_n135 ) );
  AOI21_X1 u0_u3_u1_U96 (.ZN( u0_u3_u1_n110 ) , .A( u0_u3_u1_n116 ) , .B1( u0_u3_u1_n152 ) , .B2( u0_u3_u1_n160 ) );
  NAND3_X1 u0_u3_u1_U97 (.A3( u0_u3_u1_n149 ) , .A2( u0_u3_u1_n150 ) , .A1( u0_u3_u1_n151 ) , .ZN( u0_u3_u1_n164 ) );
  NAND3_X1 u0_u3_u1_U98 (.A3( u0_u3_u1_n134 ) , .A2( u0_u3_u1_n135 ) , .ZN( u0_u3_u1_n136 ) , .A1( u0_u3_u1_n151 ) );
  NAND3_X1 u0_u3_u1_U99 (.A1( u0_u3_u1_n133 ) , .ZN( u0_u3_u1_n137 ) , .A2( u0_u3_u1_n154 ) , .A3( u0_u3_u1_n181 ) );
  OAI22_X1 u0_u3_u2_U10 (.B1( u0_u3_u2_n151 ) , .A2( u0_u3_u2_n152 ) , .A1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n160 ) , .B2( u0_u3_u2_n168 ) );
  NAND3_X1 u0_u3_u2_U100 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n98 ) );
  NOR3_X1 u0_u3_u2_U11 (.A1( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n151 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U12 (.B2( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n125 ) , .A( u0_u3_u2_n171 ) , .B1( u0_u3_u2_n184 ) );
  INV_X1 u0_u3_u2_U13 (.A( u0_u3_u2_n150 ) , .ZN( u0_u3_u2_n184 ) );
  AOI21_X1 u0_u3_u2_U14 (.ZN( u0_u3_u2_n144 ) , .B2( u0_u3_u2_n155 ) , .A( u0_u3_u2_n172 ) , .B1( u0_u3_u2_n185 ) );
  AOI21_X1 u0_u3_u2_U15 (.B2( u0_u3_u2_n143 ) , .ZN( u0_u3_u2_n145 ) , .B1( u0_u3_u2_n152 ) , .A( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U16 (.A( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n171 ) );
  INV_X1 u0_u3_u2_U17 (.A( u0_u3_u2_n120 ) , .ZN( u0_u3_u2_n188 ) );
  NAND2_X1 u0_u3_u2_U18 (.A2( u0_u3_u2_n122 ) , .ZN( u0_u3_u2_n150 ) , .A1( u0_u3_u2_n152 ) );
  INV_X1 u0_u3_u2_U19 (.A( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n170 ) );
  INV_X1 u0_u3_u2_U20 (.A( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n173 ) );
  NAND2_X1 u0_u3_u2_U21 (.A1( u0_u3_u2_n132 ) , .A2( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n157 ) );
  INV_X1 u0_u3_u2_U22 (.A( u0_u3_u2_n113 ) , .ZN( u0_u3_u2_n178 ) );
  INV_X1 u0_u3_u2_U23 (.A( u0_u3_u2_n139 ) , .ZN( u0_u3_u2_n175 ) );
  INV_X1 u0_u3_u2_U24 (.A( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n181 ) );
  INV_X1 u0_u3_u2_U25 (.A( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n177 ) );
  INV_X1 u0_u3_u2_U26 (.A( u0_u3_u2_n116 ) , .ZN( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U27 (.A( u0_u3_u2_n131 ) , .ZN( u0_u3_u2_n179 ) );
  INV_X1 u0_u3_u2_U28 (.A( u0_u3_u2_n154 ) , .ZN( u0_u3_u2_n176 ) );
  NAND2_X1 u0_u3_u2_U29 (.A2( u0_u3_u2_n116 ) , .A1( u0_u3_u2_n117 ) , .ZN( u0_u3_u2_n118 ) );
  NOR2_X1 u0_u3_u2_U3 (.ZN( u0_u3_u2_n121 ) , .A2( u0_u3_u2_n177 ) , .A1( u0_u3_u2_n180 ) );
  INV_X1 u0_u3_u2_U30 (.A( u0_u3_u2_n132 ) , .ZN( u0_u3_u2_n182 ) );
  INV_X1 u0_u3_u2_U31 (.A( u0_u3_u2_n158 ) , .ZN( u0_u3_u2_n183 ) );
  OAI21_X1 u0_u3_u2_U32 (.A( u0_u3_u2_n156 ) , .B1( u0_u3_u2_n157 ) , .ZN( u0_u3_u2_n158 ) , .B2( u0_u3_u2_n179 ) );
  NOR2_X1 u0_u3_u2_U33 (.ZN( u0_u3_u2_n156 ) , .A1( u0_u3_u2_n166 ) , .A2( u0_u3_u2_n169 ) );
  NOR2_X1 u0_u3_u2_U34 (.A2( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n140 ) );
  NOR2_X1 u0_u3_u2_U35 (.A2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n153 ) , .A1( u0_u3_u2_n156 ) );
  AOI211_X1 u0_u3_u2_U36 (.ZN( u0_u3_u2_n130 ) , .C1( u0_u3_u2_n138 ) , .C2( u0_u3_u2_n179 ) , .B( u0_u3_u2_n96 ) , .A( u0_u3_u2_n97 ) );
  OAI22_X1 u0_u3_u2_U37 (.B1( u0_u3_u2_n133 ) , .A2( u0_u3_u2_n137 ) , .A1( u0_u3_u2_n152 ) , .B2( u0_u3_u2_n168 ) , .ZN( u0_u3_u2_n97 ) );
  OAI221_X1 u0_u3_u2_U38 (.B1( u0_u3_u2_n113 ) , .C1( u0_u3_u2_n132 ) , .A( u0_u3_u2_n149 ) , .B2( u0_u3_u2_n171 ) , .C2( u0_u3_u2_n172 ) , .ZN( u0_u3_u2_n96 ) );
  OAI221_X1 u0_u3_u2_U39 (.A( u0_u3_u2_n115 ) , .C2( u0_u3_u2_n123 ) , .B2( u0_u3_u2_n143 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n163 ) , .C1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U4 (.A( u0_u3_u2_n134 ) , .ZN( u0_u3_u2_n185 ) );
  OAI21_X1 u0_u3_u2_U40 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n115 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n178 ) );
  OAI221_X1 u0_u3_u2_U41 (.A( u0_u3_u2_n135 ) , .B2( u0_u3_u2_n136 ) , .B1( u0_u3_u2_n137 ) , .ZN( u0_u3_u2_n162 ) , .C2( u0_u3_u2_n167 ) , .C1( u0_u3_u2_n185 ) );
  AND3_X1 u0_u3_u2_U42 (.A3( u0_u3_u2_n131 ) , .A2( u0_u3_u2_n132 ) , .A1( u0_u3_u2_n133 ) , .ZN( u0_u3_u2_n136 ) );
  AOI22_X1 u0_u3_u2_U43 (.ZN( u0_u3_u2_n135 ) , .B1( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n156 ) , .B2( u0_u3_u2_n180 ) , .A2( u0_u3_u2_n188 ) );
  AOI21_X1 u0_u3_u2_U44 (.ZN( u0_u3_u2_n149 ) , .B1( u0_u3_u2_n173 ) , .B2( u0_u3_u2_n188 ) , .A( u0_u3_u2_n95 ) );
  AND3_X1 u0_u3_u2_U45 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n156 ) , .ZN( u0_u3_u2_n95 ) );
  OAI21_X1 u0_u3_u2_U46 (.A( u0_u3_u2_n141 ) , .B2( u0_u3_u2_n142 ) , .ZN( u0_u3_u2_n146 ) , .B1( u0_u3_u2_n153 ) );
  OAI21_X1 u0_u3_u2_U47 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n141 ) , .B1( u0_u3_u2_n176 ) , .B2( u0_u3_u2_n177 ) );
  NOR3_X1 u0_u3_u2_U48 (.ZN( u0_u3_u2_n142 ) , .A3( u0_u3_u2_n175 ) , .A2( u0_u3_u2_n178 ) , .A1( u0_u3_u2_n181 ) );
  OAI21_X1 u0_u3_u2_U49 (.A( u0_u3_u2_n101 ) , .B2( u0_u3_u2_n121 ) , .B1( u0_u3_u2_n153 ) , .ZN( u0_u3_u2_n164 ) );
  NOR4_X1 u0_u3_u2_U5 (.A4( u0_u3_u2_n124 ) , .A3( u0_u3_u2_n125 ) , .A2( u0_u3_u2_n126 ) , .A1( u0_u3_u2_n127 ) , .ZN( u0_u3_u2_n128 ) );
  NAND2_X1 u0_u3_u2_U50 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U51 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n143 ) );
  NAND2_X1 u0_u3_u2_U52 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n152 ) );
  NAND2_X1 u0_u3_u2_U53 (.A1( u0_u3_u2_n100 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n132 ) );
  INV_X1 u0_u3_u2_U54 (.A( u0_u3_u2_n140 ) , .ZN( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U55 (.A( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n167 ) );
  INV_X1 u0_u3_u2_U56 (.ZN( u0_u3_u2_n187 ) , .A( u0_u3_u2_n99 ) );
  OAI21_X1 u0_u3_u2_U57 (.B1( u0_u3_u2_n137 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n98 ) , .ZN( u0_u3_u2_n99 ) );
  NAND2_X1 u0_u3_u2_U58 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n113 ) );
  NAND2_X1 u0_u3_u2_U59 (.A1( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n131 ) );
  AOI21_X1 u0_u3_u2_U6 (.B2( u0_u3_u2_n119 ) , .ZN( u0_u3_u2_n127 ) , .A( u0_u3_u2_n137 ) , .B1( u0_u3_u2_n155 ) );
  NAND2_X1 u0_u3_u2_U60 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n107 ) , .ZN( u0_u3_u2_n139 ) );
  NAND2_X1 u0_u3_u2_U61 (.A1( u0_u3_u2_n103 ) , .A2( u0_u3_u2_n105 ) , .ZN( u0_u3_u2_n133 ) );
  NAND2_X1 u0_u3_u2_U62 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n103 ) , .ZN( u0_u3_u2_n154 ) );
  NAND2_X1 u0_u3_u2_U63 (.A2( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n104 ) , .ZN( u0_u3_u2_n119 ) );
  NAND2_X1 u0_u3_u2_U64 (.A2( u0_u3_u2_n107 ) , .A1( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n123 ) );
  NAND2_X1 u0_u3_u2_U65 (.A1( u0_u3_u2_n104 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n122 ) );
  INV_X1 u0_u3_u2_U66 (.A( u0_u3_u2_n114 ) , .ZN( u0_u3_u2_n172 ) );
  NAND2_X1 u0_u3_u2_U67 (.A2( u0_u3_u2_n100 ) , .A1( u0_u3_u2_n102 ) , .ZN( u0_u3_u2_n116 ) );
  NAND2_X1 u0_u3_u2_U68 (.A1( u0_u3_u2_n102 ) , .A2( u0_u3_u2_n108 ) , .ZN( u0_u3_u2_n120 ) );
  NAND2_X1 u0_u3_u2_U69 (.A2( u0_u3_u2_n105 ) , .A1( u0_u3_u2_n106 ) , .ZN( u0_u3_u2_n117 ) );
  AOI21_X1 u0_u3_u2_U7 (.ZN( u0_u3_u2_n124 ) , .B1( u0_u3_u2_n131 ) , .B2( u0_u3_u2_n143 ) , .A( u0_u3_u2_n172 ) );
  NOR2_X1 u0_u3_u2_U70 (.A2( u0_u3_X_16 ) , .ZN( u0_u3_u2_n140 ) , .A1( u0_u3_u2_n166 ) );
  NOR2_X1 u0_u3_u2_U71 (.A2( u0_u3_X_13 ) , .A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n100 ) );
  NOR2_X1 u0_u3_u2_U72 (.A2( u0_u3_X_16 ) , .A1( u0_u3_X_17 ) , .ZN( u0_u3_u2_n138 ) );
  NOR2_X1 u0_u3_u2_U73 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n104 ) );
  NOR2_X1 u0_u3_u2_U74 (.A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n103 ) , .A1( u0_u3_u2_n174 ) );
  NOR2_X1 u0_u3_u2_U75 (.A2( u0_u3_X_15 ) , .ZN( u0_u3_u2_n102 ) , .A1( u0_u3_u2_n165 ) );
  NOR2_X1 u0_u3_u2_U76 (.A2( u0_u3_X_17 ) , .ZN( u0_u3_u2_n114 ) , .A1( u0_u3_u2_n169 ) );
  AND2_X1 u0_u3_u2_U77 (.A1( u0_u3_X_15 ) , .ZN( u0_u3_u2_n105 ) , .A2( u0_u3_u2_n165 ) );
  AND2_X1 u0_u3_u2_U78 (.A2( u0_u3_X_15 ) , .A1( u0_u3_X_18 ) , .ZN( u0_u3_u2_n107 ) );
  AND2_X1 u0_u3_u2_U79 (.A1( u0_u3_X_14 ) , .ZN( u0_u3_u2_n106 ) , .A2( u0_u3_u2_n174 ) );
  AOI21_X1 u0_u3_u2_U8 (.B2( u0_u3_u2_n120 ) , .B1( u0_u3_u2_n121 ) , .ZN( u0_u3_u2_n126 ) , .A( u0_u3_u2_n167 ) );
  AND2_X1 u0_u3_u2_U80 (.A1( u0_u3_X_13 ) , .A2( u0_u3_X_14 ) , .ZN( u0_u3_u2_n108 ) );
  INV_X1 u0_u3_u2_U81 (.A( u0_u3_X_16 ) , .ZN( u0_u3_u2_n169 ) );
  INV_X1 u0_u3_u2_U82 (.A( u0_u3_X_17 ) , .ZN( u0_u3_u2_n166 ) );
  INV_X1 u0_u3_u2_U83 (.A( u0_u3_X_13 ) , .ZN( u0_u3_u2_n174 ) );
  INV_X1 u0_u3_u2_U84 (.A( u0_u3_X_18 ) , .ZN( u0_u3_u2_n165 ) );
  NAND4_X1 u0_u3_u2_U85 (.ZN( u0_out3_24 ) , .A4( u0_u3_u2_n111 ) , .A3( u0_u3_u2_n112 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n187 ) );
  AOI221_X1 u0_u3_u2_U86 (.A( u0_u3_u2_n109 ) , .B1( u0_u3_u2_n110 ) , .ZN( u0_u3_u2_n111 ) , .C1( u0_u3_u2_n134 ) , .C2( u0_u3_u2_n170 ) , .B2( u0_u3_u2_n173 ) );
  AOI21_X1 u0_u3_u2_U87 (.ZN( u0_u3_u2_n112 ) , .B2( u0_u3_u2_n156 ) , .A( u0_u3_u2_n164 ) , .B1( u0_u3_u2_n181 ) );
  NAND4_X1 u0_u3_u2_U88 (.ZN( u0_out3_16 ) , .A4( u0_u3_u2_n128 ) , .A3( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n130 ) , .A2( u0_u3_u2_n186 ) );
  AOI22_X1 u0_u3_u2_U89 (.A2( u0_u3_u2_n118 ) , .ZN( u0_u3_u2_n129 ) , .A1( u0_u3_u2_n140 ) , .B1( u0_u3_u2_n157 ) , .B2( u0_u3_u2_n170 ) );
  OAI22_X1 u0_u3_u2_U9 (.ZN( u0_u3_u2_n109 ) , .A2( u0_u3_u2_n113 ) , .B2( u0_u3_u2_n133 ) , .B1( u0_u3_u2_n167 ) , .A1( u0_u3_u2_n168 ) );
  INV_X1 u0_u3_u2_U90 (.A( u0_u3_u2_n163 ) , .ZN( u0_u3_u2_n186 ) );
  NAND4_X1 u0_u3_u2_U91 (.ZN( u0_out3_30 ) , .A4( u0_u3_u2_n147 ) , .A3( u0_u3_u2_n148 ) , .A2( u0_u3_u2_n149 ) , .A1( u0_u3_u2_n187 ) );
  AOI21_X1 u0_u3_u2_U92 (.B2( u0_u3_u2_n138 ) , .ZN( u0_u3_u2_n148 ) , .A( u0_u3_u2_n162 ) , .B1( u0_u3_u2_n182 ) );
  NOR3_X1 u0_u3_u2_U93 (.A3( u0_u3_u2_n144 ) , .A2( u0_u3_u2_n145 ) , .A1( u0_u3_u2_n146 ) , .ZN( u0_u3_u2_n147 ) );
  OR4_X1 u0_u3_u2_U94 (.ZN( u0_out3_6 ) , .A4( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n162 ) , .A2( u0_u3_u2_n163 ) , .A1( u0_u3_u2_n164 ) );
  OR3_X1 u0_u3_u2_U95 (.A2( u0_u3_u2_n159 ) , .A1( u0_u3_u2_n160 ) , .ZN( u0_u3_u2_n161 ) , .A3( u0_u3_u2_n183 ) );
  AOI21_X1 u0_u3_u2_U96 (.B2( u0_u3_u2_n154 ) , .B1( u0_u3_u2_n155 ) , .ZN( u0_u3_u2_n159 ) , .A( u0_u3_u2_n167 ) );
  NAND3_X1 u0_u3_u2_U97 (.A2( u0_u3_u2_n117 ) , .A1( u0_u3_u2_n122 ) , .A3( u0_u3_u2_n123 ) , .ZN( u0_u3_u2_n134 ) );
  NAND3_X1 u0_u3_u2_U98 (.ZN( u0_u3_u2_n110 ) , .A2( u0_u3_u2_n131 ) , .A3( u0_u3_u2_n139 ) , .A1( u0_u3_u2_n154 ) );
  NAND3_X1 u0_u3_u2_U99 (.A2( u0_u3_u2_n100 ) , .ZN( u0_u3_u2_n101 ) , .A1( u0_u3_u2_n104 ) , .A3( u0_u3_u2_n114 ) );
  OAI22_X1 u0_u3_u3_U10 (.B1( u0_u3_u3_n113 ) , .A2( u0_u3_u3_n135 ) , .A1( u0_u3_u3_n150 ) , .B2( u0_u3_u3_n164 ) , .ZN( u0_u3_u3_n98 ) );
  OAI211_X1 u0_u3_u3_U11 (.B( u0_u3_u3_n106 ) , .ZN( u0_u3_u3_n119 ) , .C2( u0_u3_u3_n128 ) , .C1( u0_u3_u3_n167 ) , .A( u0_u3_u3_n181 ) );
  AOI221_X1 u0_u3_u3_U12 (.C1( u0_u3_u3_n105 ) , .ZN( u0_u3_u3_n106 ) , .A( u0_u3_u3_n131 ) , .B2( u0_u3_u3_n132 ) , .C2( u0_u3_u3_n133 ) , .B1( u0_u3_u3_n169 ) );
  INV_X1 u0_u3_u3_U13 (.ZN( u0_u3_u3_n181 ) , .A( u0_u3_u3_n98 ) );
  NAND2_X1 u0_u3_u3_U14 (.ZN( u0_u3_u3_n105 ) , .A2( u0_u3_u3_n130 ) , .A1( u0_u3_u3_n155 ) );
  AOI22_X1 u0_u3_u3_U15 (.B1( u0_u3_u3_n115 ) , .A2( u0_u3_u3_n116 ) , .ZN( u0_u3_u3_n123 ) , .B2( u0_u3_u3_n133 ) , .A1( u0_u3_u3_n169 ) );
  NAND2_X1 u0_u3_u3_U16 (.ZN( u0_u3_u3_n116 ) , .A2( u0_u3_u3_n151 ) , .A1( u0_u3_u3_n182 ) );
  NOR2_X1 u0_u3_u3_U17 (.ZN( u0_u3_u3_n126 ) , .A2( u0_u3_u3_n150 ) , .A1( u0_u3_u3_n164 ) );
  AOI21_X1 u0_u3_u3_U18 (.ZN( u0_u3_u3_n112 ) , .B2( u0_u3_u3_n146 ) , .B1( u0_u3_u3_n155 ) , .A( u0_u3_u3_n167 ) );
  NAND2_X1 u0_u3_u3_U19 (.A1( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n142 ) , .A2( u0_u3_u3_n164 ) );
  NAND2_X1 u0_u3_u3_U20 (.ZN( u0_u3_u3_n132 ) , .A2( u0_u3_u3_n152 ) , .A1( u0_u3_u3_n156 ) );
  INV_X1 u0_u3_u3_U21 (.A( u0_u3_u3_n133 ) , .ZN( u0_u3_u3_n165 ) );
  NAND2_X1 u0_u3_u3_U22 (.ZN( u0_u3_u3_n143 ) , .A1( u0_u3_u3_n165 ) , .A2( u0_u3_u3_n167 ) );
  AND2_X1 u0_u3_u3_U23 (.A2( u0_u3_u3_n113 ) , .A1( u0_u3_u3_n114 ) , .ZN( u0_u3_u3_n151 ) );
  INV_X1 u0_u3_u3_U24 (.A( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n170 ) );
  NAND2_X1 u0_u3_u3_U25 (.A1( u0_u3_u3_n107 ) , .A2( u0_u3_u3_n108 ) , .ZN( u0_u3_u3_n140 ) );
  NAND2_X1 u0_u3_u3_U26 (.ZN( u0_u3_u3_n117 ) , .A1( u0_u3_u3_n124 ) , .A2( u0_u3_u3_n148 ) );
  INV_X1 u0_u3_u3_U27 (.A( u0_u3_u3_n130 ) , .ZN( u0_u3_u3_n177 ) );
  INV_X1 u0_u3_u3_U28 (.A( u0_u3_u3_n128 ) , .ZN( u0_u3_u3_n176 ) );
  INV_X1 u0_u3_u3_U29 (.A( u0_u3_u3_n155 ) , .ZN( u0_u3_u3_n174 ) );
  INV_X1 u0_u3_u3_U3 (.A( u0_u3_u3_n140 ) , .ZN( u0_u3_u3_n182 ) );
  INV_X1 u0_u3_u3_U30 (.A( u0_u3_u3_n139 ) , .ZN( u0_u3_u3_n185 ) );
  NOR2_X1 u0_u3_u3_U31 (.ZN( u0_u3_u3_n135 ) , .A2( u0_u3_u3_n141 ) , .A1( u0_u3_u3_n169 ) );
  INV_X1 u0_u3_u3_U32 (.A( u0_u3_u3_n156 ) , .ZN( u0_u3_u3_n179 ) );
  OAI22_X1 u0_u3_u3_U33 (.B1( u0_u3_u3_n118 ) , .ZN( u0_u3_u3_n120 ) , .A1( u0_u3_u3_n135 ) , .B2( u0_u3_u3_n154 ) , .A2( u0_u3_u3_n178 ) );
  AND3_X1 u0_u3_u3_U34 (.ZN( u0_u3_u3_n118 ) , .A2( u0_u3_u3_n124 ) , .A1( u0_u3_u3_n144 ) , .A3( u0_u3_u3_n152 ) );
  OAI222_X1 u0_u3_u3_U35 (.C2( u0_u3_u3_n107 ) , .A2( u0_u3_u3_n108 ) , .B1( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n138 ) , .B2( u0_u3_u3_n146 ) , .C1( u0_u3_u3_n154 ) , .A1( u0_u3_u3_n164 ) );
  NOR4_X1 u0_u3_u3_U36 (.A4( u0_u3_u3_n157 ) , .A3( u0_u3_u3_n158 ) , .A2( u0_u3_u3_n159 ) , .A1( u0_u3_u3_n160 ) , .ZN( u0_u3_u3_n161 ) );
  AOI21_X1 u0_u3_u3_U37 (.B2( u0_u3_u3_n152 ) , .B1( u0_u3_u3_n153 ) , .ZN( u0_u3_u3_n158 ) , .A( u0_u3_u3_n164 ) );
  AOI21_X1 u0_u3_u3_U38 (.A( u0_u3_u3_n149 ) , .B2( u0_u3_u3_n150 ) , .B1( u0_u3_u3_n151 ) , .ZN( u0_u3_u3_n159 ) );
  AOI21_X1 u0_u3_u3_U39 (.A( u0_u3_u3_n154 ) , .B2( u0_u3_u3_n155 ) , .B1( u0_u3_u3_n156 ) , .ZN( u0_u3_u3_n157 ) );
  INV_X1 u0_u3_u3_U4 (.A( u0_u3_u3_n129 ) , .ZN( u0_u3_u3_n183 ) );
  AOI211_X1 u0_u3_u3_U40 (.ZN( u0_u3_u3_n109 ) , .A( u0_u3_u3_n119 ) , .C2( u0_u3_u3_n129 ) , .B( u0_u3_u3_n138 ) , .C1( u0_u3_u3_n141 ) );
  INV_X1 u0_u3_u3_U41 (.A( u0_u3_u3_n121 ) , .ZN( u0_u3_u3_n164 ) );
  NAND2_X1 u0_u3_u3_U42 (.ZN( u0_u3_u3_n133 ) , .A1( u0_u3_u3_n154 ) , .A2( u0_u3_u3_n164 ) );
  OAI211_X1 u0_u3_u3_U43 (.B( u0_u3_u3_n127 ) , .ZN( u0_u3_u3_n139 ) , .C1( u0_u3_u3_n150 ) , .C2( u0_u3_u3_n154 ) , .A( u0_u3_u3_n184 ) );
  INV_X1 u0_u3_u3_U44 (.A( u0_u3_u3_n125 ) , .ZN( u0_u3_u3_n184 ) );
  AOI221_X1 u0_u3_u3_U45 (.A( u0_u3_u3_n126 ) , .ZN( u0_u3_u3_n127 ) , .C2( u0_u3_u3_n132 ) , .C1( u0_u3_u3_n169 ) , .B2( u0_u3_u3_n170 ) , .B1( u0_u3_u3_n174 ) );
  OAI22_X1 u0_u3_u3_U46 (.A1( u0_u3_u3_n124 ) , .ZN( u0_u3_u3_n125 ) , .B2( u0_u3_u3_n145 ) , .A2( u0_u3_u3_n165 ) , .B1( u0_u3_u3_n167 ) );
  NOR2_X1 u0_u3_u3_U47 (.A1( u0_u3_u3_n113 ) , .ZN( u0_u3_u3_n131 ) , .A2( u0_u3_u3_n154 ) );
  NAND2_X1 u0_u3_u3_U48 (.A1( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n150 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U49 (.A2( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n155 ) , .A1( u0_u3_u3_n97 ) );
  INV_X1 u0_u3_u3_U5 (.A( u0_u3_u3_n117 ) , .ZN( u0_u3_u3_n178 ) );
  INV_X1 u0_u3_u3_U50 (.A( u0_u3_u3_n141 ) , .ZN( u0_u3_u3_n167 ) );
  AOI21_X1 u0_u3_u3_U51 (.B2( u0_u3_u3_n114 ) , .B1( u0_u3_u3_n146 ) , .A( u0_u3_u3_n154 ) , .ZN( u0_u3_u3_n94 ) );
  AOI21_X1 u0_u3_u3_U52 (.ZN( u0_u3_u3_n110 ) , .B2( u0_u3_u3_n142 ) , .B1( u0_u3_u3_n186 ) , .A( u0_u3_u3_n95 ) );
  INV_X1 u0_u3_u3_U53 (.A( u0_u3_u3_n145 ) , .ZN( u0_u3_u3_n186 ) );
  AOI21_X1 u0_u3_u3_U54 (.B1( u0_u3_u3_n124 ) , .A( u0_u3_u3_n149 ) , .B2( u0_u3_u3_n155 ) , .ZN( u0_u3_u3_n95 ) );
  INV_X1 u0_u3_u3_U55 (.A( u0_u3_u3_n149 ) , .ZN( u0_u3_u3_n169 ) );
  NAND2_X1 u0_u3_u3_U56 (.ZN( u0_u3_u3_n124 ) , .A1( u0_u3_u3_n96 ) , .A2( u0_u3_u3_n97 ) );
  NAND2_X1 u0_u3_u3_U57 (.A2( u0_u3_u3_n100 ) , .ZN( u0_u3_u3_n146 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U58 (.A1( u0_u3_u3_n101 ) , .ZN( u0_u3_u3_n145 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U59 (.A1( u0_u3_u3_n100 ) , .ZN( u0_u3_u3_n156 ) , .A2( u0_u3_u3_n99 ) );
  AOI221_X1 u0_u3_u3_U6 (.A( u0_u3_u3_n131 ) , .C2( u0_u3_u3_n132 ) , .C1( u0_u3_u3_n133 ) , .ZN( u0_u3_u3_n134 ) , .B1( u0_u3_u3_n143 ) , .B2( u0_u3_u3_n177 ) );
  NAND2_X1 u0_u3_u3_U60 (.A2( u0_u3_u3_n101 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n148 ) );
  NAND2_X1 u0_u3_u3_U61 (.A1( u0_u3_u3_n100 ) , .A2( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n128 ) );
  NAND2_X1 u0_u3_u3_U62 (.A2( u0_u3_u3_n101 ) , .A1( u0_u3_u3_n102 ) , .ZN( u0_u3_u3_n152 ) );
  NAND2_X1 u0_u3_u3_U63 (.A2( u0_u3_u3_n101 ) , .ZN( u0_u3_u3_n114 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U64 (.ZN( u0_u3_u3_n107 ) , .A1( u0_u3_u3_n97 ) , .A2( u0_u3_u3_n99 ) );
  NAND2_X1 u0_u3_u3_U65 (.A2( u0_u3_u3_n100 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n113 ) );
  NAND2_X1 u0_u3_u3_U66 (.A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n153 ) , .A2( u0_u3_u3_n97 ) );
  NAND2_X1 u0_u3_u3_U67 (.A2( u0_u3_u3_n103 ) , .A1( u0_u3_u3_n104 ) , .ZN( u0_u3_u3_n130 ) );
  NAND2_X1 u0_u3_u3_U68 (.A2( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n144 ) , .A1( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U69 (.A1( u0_u3_u3_n102 ) , .A2( u0_u3_u3_n103 ) , .ZN( u0_u3_u3_n108 ) );
  OAI22_X1 u0_u3_u3_U7 (.B2( u0_u3_u3_n147 ) , .A2( u0_u3_u3_n148 ) , .ZN( u0_u3_u3_n160 ) , .B1( u0_u3_u3_n165 ) , .A1( u0_u3_u3_n168 ) );
  NOR2_X1 u0_u3_u3_U70 (.A2( u0_u3_X_19 ) , .A1( u0_u3_X_20 ) , .ZN( u0_u3_u3_n99 ) );
  NOR2_X1 u0_u3_u3_U71 (.A2( u0_u3_X_21 ) , .A1( u0_u3_X_24 ) , .ZN( u0_u3_u3_n103 ) );
  NOR2_X1 u0_u3_u3_U72 (.A2( u0_u3_X_24 ) , .A1( u0_u3_u3_n171 ) , .ZN( u0_u3_u3_n97 ) );
  NOR2_X1 u0_u3_u3_U73 (.A2( u0_u3_X_19 ) , .A1( u0_u3_u3_n172 ) , .ZN( u0_u3_u3_n96 ) );
  NAND2_X1 u0_u3_u3_U74 (.A1( u0_u3_X_22 ) , .A2( u0_u3_X_23 ) , .ZN( u0_u3_u3_n154 ) );
  AND2_X1 u0_u3_u3_U75 (.A1( u0_u3_X_24 ) , .ZN( u0_u3_u3_n101 ) , .A2( u0_u3_u3_n171 ) );
  AND2_X1 u0_u3_u3_U76 (.A1( u0_u3_X_19 ) , .ZN( u0_u3_u3_n102 ) , .A2( u0_u3_u3_n172 ) );
  AND2_X1 u0_u3_u3_U77 (.A1( u0_u3_X_21 ) , .A2( u0_u3_X_24 ) , .ZN( u0_u3_u3_n100 ) );
  AND2_X1 u0_u3_u3_U78 (.A2( u0_u3_X_19 ) , .A1( u0_u3_X_20 ) , .ZN( u0_u3_u3_n104 ) );
  INV_X1 u0_u3_u3_U79 (.A( u0_u3_X_21 ) , .ZN( u0_u3_u3_n171 ) );
  AND3_X1 u0_u3_u3_U8 (.A3( u0_u3_u3_n144 ) , .A2( u0_u3_u3_n145 ) , .A1( u0_u3_u3_n146 ) , .ZN( u0_u3_u3_n147 ) );
  INV_X1 u0_u3_u3_U80 (.A( u0_u3_X_20 ) , .ZN( u0_u3_u3_n172 ) );
  INV_X1 u0_u3_u3_U81 (.A( u0_u3_X_22 ) , .ZN( u0_u3_u3_n166 ) );
  NAND4_X1 u0_u3_u3_U82 (.ZN( u0_out3_26 ) , .A4( u0_u3_u3_n109 ) , .A3( u0_u3_u3_n110 ) , .A2( u0_u3_u3_n111 ) , .A1( u0_u3_u3_n173 ) );
  INV_X1 u0_u3_u3_U83 (.ZN( u0_u3_u3_n173 ) , .A( u0_u3_u3_n94 ) );
  OAI21_X1 u0_u3_u3_U84 (.ZN( u0_u3_u3_n111 ) , .B2( u0_u3_u3_n117 ) , .A( u0_u3_u3_n133 ) , .B1( u0_u3_u3_n176 ) );
  NAND4_X1 u0_u3_u3_U85 (.ZN( u0_out3_1 ) , .A4( u0_u3_u3_n161 ) , .A3( u0_u3_u3_n162 ) , .A2( u0_u3_u3_n163 ) , .A1( u0_u3_u3_n185 ) );
  NAND2_X1 u0_u3_u3_U86 (.ZN( u0_u3_u3_n163 ) , .A2( u0_u3_u3_n170 ) , .A1( u0_u3_u3_n176 ) );
  AOI22_X1 u0_u3_u3_U87 (.B2( u0_u3_u3_n140 ) , .B1( u0_u3_u3_n141 ) , .A2( u0_u3_u3_n142 ) , .ZN( u0_u3_u3_n162 ) , .A1( u0_u3_u3_n177 ) );
  NAND4_X1 u0_u3_u3_U88 (.ZN( u0_out3_20 ) , .A4( u0_u3_u3_n122 ) , .A3( u0_u3_u3_n123 ) , .A1( u0_u3_u3_n175 ) , .A2( u0_u3_u3_n180 ) );
  INV_X1 u0_u3_u3_U89 (.A( u0_u3_u3_n126 ) , .ZN( u0_u3_u3_n180 ) );
  INV_X1 u0_u3_u3_U9 (.A( u0_u3_u3_n143 ) , .ZN( u0_u3_u3_n168 ) );
  INV_X1 u0_u3_u3_U90 (.A( u0_u3_u3_n112 ) , .ZN( u0_u3_u3_n175 ) );
  OR4_X1 u0_u3_u3_U91 (.ZN( u0_out3_10 ) , .A4( u0_u3_u3_n136 ) , .A3( u0_u3_u3_n137 ) , .A1( u0_u3_u3_n138 ) , .A2( u0_u3_u3_n139 ) );
  OAI222_X1 u0_u3_u3_U92 (.C1( u0_u3_u3_n128 ) , .ZN( u0_u3_u3_n137 ) , .B1( u0_u3_u3_n148 ) , .A2( u0_u3_u3_n150 ) , .B2( u0_u3_u3_n154 ) , .C2( u0_u3_u3_n164 ) , .A1( u0_u3_u3_n167 ) );
  AOI211_X1 u0_u3_u3_U93 (.B( u0_u3_u3_n119 ) , .A( u0_u3_u3_n120 ) , .C2( u0_u3_u3_n121 ) , .ZN( u0_u3_u3_n122 ) , .C1( u0_u3_u3_n179 ) );
  OAI221_X1 u0_u3_u3_U94 (.A( u0_u3_u3_n134 ) , .B2( u0_u3_u3_n135 ) , .ZN( u0_u3_u3_n136 ) , .C1( u0_u3_u3_n149 ) , .B1( u0_u3_u3_n151 ) , .C2( u0_u3_u3_n183 ) );
  NOR2_X1 u0_u3_u3_U95 (.A2( u0_u3_X_23 ) , .ZN( u0_u3_u3_n141 ) , .A1( u0_u3_u3_n166 ) );
  NAND2_X1 u0_u3_u3_U96 (.A1( u0_u3_X_23 ) , .ZN( u0_u3_u3_n149 ) , .A2( u0_u3_u3_n166 ) );
  NOR2_X1 u0_u3_u3_U97 (.A2( u0_u3_X_22 ) , .A1( u0_u3_X_23 ) , .ZN( u0_u3_u3_n121 ) );
  NAND3_X1 u0_u3_u3_U98 (.A1( u0_u3_u3_n114 ) , .ZN( u0_u3_u3_n115 ) , .A2( u0_u3_u3_n145 ) , .A3( u0_u3_u3_n153 ) );
  NAND3_X1 u0_u3_u3_U99 (.ZN( u0_u3_u3_n129 ) , .A2( u0_u3_u3_n144 ) , .A1( u0_u3_u3_n153 ) , .A3( u0_u3_u3_n182 ) );
  XOR2_X1 u0_u4_U26 (.B( u0_K5_30 ) , .A( u0_R3_21 ) , .Z( u0_u4_X_30 ) );
  XOR2_X1 u0_u4_U28 (.B( u0_K5_29 ) , .A( u0_R3_20 ) , .Z( u0_u4_X_29 ) );
  XOR2_X1 u0_u4_U29 (.B( u0_K5_28 ) , .A( u0_R3_19 ) , .Z( u0_u4_X_28 ) );
  XOR2_X1 u0_u4_U30 (.B( u0_K5_27 ) , .A( u0_R3_18 ) , .Z( u0_u4_X_27 ) );
  XOR2_X1 u0_u4_U31 (.B( u0_K5_26 ) , .A( u0_R3_17 ) , .Z( u0_u4_X_26 ) );
  XOR2_X1 u0_u4_U32 (.B( u0_K5_25 ) , .A( u0_R3_16 ) , .Z( u0_u4_X_25 ) );
  OAI22_X1 u0_u4_u4_U10 (.B2( u0_u4_u4_n135 ) , .ZN( u0_u4_u4_n137 ) , .B1( u0_u4_u4_n153 ) , .A1( u0_u4_u4_n155 ) , .A2( u0_u4_u4_n171 ) );
  AND3_X1 u0_u4_u4_U11 (.A2( u0_u4_u4_n134 ) , .ZN( u0_u4_u4_n135 ) , .A3( u0_u4_u4_n145 ) , .A1( u0_u4_u4_n157 ) );
  NAND2_X1 u0_u4_u4_U12 (.ZN( u0_u4_u4_n132 ) , .A2( u0_u4_u4_n170 ) , .A1( u0_u4_u4_n173 ) );
  AOI21_X1 u0_u4_u4_U13 (.B2( u0_u4_u4_n160 ) , .B1( u0_u4_u4_n161 ) , .ZN( u0_u4_u4_n162 ) , .A( u0_u4_u4_n170 ) );
  AOI21_X1 u0_u4_u4_U14 (.ZN( u0_u4_u4_n107 ) , .B2( u0_u4_u4_n143 ) , .A( u0_u4_u4_n174 ) , .B1( u0_u4_u4_n184 ) );
  AOI21_X1 u0_u4_u4_U15 (.B2( u0_u4_u4_n158 ) , .B1( u0_u4_u4_n159 ) , .ZN( u0_u4_u4_n163 ) , .A( u0_u4_u4_n174 ) );
  AOI21_X1 u0_u4_u4_U16 (.A( u0_u4_u4_n153 ) , .B2( u0_u4_u4_n154 ) , .B1( u0_u4_u4_n155 ) , .ZN( u0_u4_u4_n165 ) );
  AOI21_X1 u0_u4_u4_U17 (.A( u0_u4_u4_n156 ) , .B2( u0_u4_u4_n157 ) , .ZN( u0_u4_u4_n164 ) , .B1( u0_u4_u4_n184 ) );
  INV_X1 u0_u4_u4_U18 (.A( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n170 ) );
  AND2_X1 u0_u4_u4_U19 (.A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n155 ) , .A1( u0_u4_u4_n160 ) );
  INV_X1 u0_u4_u4_U20 (.A( u0_u4_u4_n156 ) , .ZN( u0_u4_u4_n175 ) );
  NAND2_X1 u0_u4_u4_U21 (.A2( u0_u4_u4_n118 ) , .ZN( u0_u4_u4_n131 ) , .A1( u0_u4_u4_n147 ) );
  NAND2_X1 u0_u4_u4_U22 (.A1( u0_u4_u4_n119 ) , .A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n130 ) );
  NAND2_X1 u0_u4_u4_U23 (.ZN( u0_u4_u4_n117 ) , .A2( u0_u4_u4_n118 ) , .A1( u0_u4_u4_n148 ) );
  NAND2_X1 u0_u4_u4_U24 (.ZN( u0_u4_u4_n129 ) , .A1( u0_u4_u4_n134 ) , .A2( u0_u4_u4_n148 ) );
  AND3_X1 u0_u4_u4_U25 (.A1( u0_u4_u4_n119 ) , .A2( u0_u4_u4_n143 ) , .A3( u0_u4_u4_n154 ) , .ZN( u0_u4_u4_n161 ) );
  AND2_X1 u0_u4_u4_U26 (.A1( u0_u4_u4_n145 ) , .A2( u0_u4_u4_n147 ) , .ZN( u0_u4_u4_n159 ) );
  OR3_X1 u0_u4_u4_U27 (.A3( u0_u4_u4_n114 ) , .A2( u0_u4_u4_n115 ) , .A1( u0_u4_u4_n116 ) , .ZN( u0_u4_u4_n136 ) );
  AOI21_X1 u0_u4_u4_U28 (.A( u0_u4_u4_n113 ) , .ZN( u0_u4_u4_n116 ) , .B2( u0_u4_u4_n173 ) , .B1( u0_u4_u4_n174 ) );
  AOI21_X1 u0_u4_u4_U29 (.ZN( u0_u4_u4_n115 ) , .B2( u0_u4_u4_n145 ) , .B1( u0_u4_u4_n146 ) , .A( u0_u4_u4_n156 ) );
  NOR2_X1 u0_u4_u4_U3 (.ZN( u0_u4_u4_n121 ) , .A1( u0_u4_u4_n181 ) , .A2( u0_u4_u4_n182 ) );
  OAI22_X1 u0_u4_u4_U30 (.ZN( u0_u4_u4_n114 ) , .A2( u0_u4_u4_n121 ) , .B1( u0_u4_u4_n160 ) , .B2( u0_u4_u4_n170 ) , .A1( u0_u4_u4_n171 ) );
  INV_X1 u0_u4_u4_U31 (.A( u0_u4_u4_n158 ) , .ZN( u0_u4_u4_n182 ) );
  INV_X1 u0_u4_u4_U32 (.ZN( u0_u4_u4_n181 ) , .A( u0_u4_u4_n96 ) );
  INV_X1 u0_u4_u4_U33 (.A( u0_u4_u4_n144 ) , .ZN( u0_u4_u4_n179 ) );
  INV_X1 u0_u4_u4_U34 (.A( u0_u4_u4_n157 ) , .ZN( u0_u4_u4_n178 ) );
  NAND2_X1 u0_u4_u4_U35 (.A2( u0_u4_u4_n154 ) , .A1( u0_u4_u4_n96 ) , .ZN( u0_u4_u4_n97 ) );
  INV_X1 u0_u4_u4_U36 (.ZN( u0_u4_u4_n186 ) , .A( u0_u4_u4_n95 ) );
  OAI221_X1 u0_u4_u4_U37 (.C1( u0_u4_u4_n134 ) , .B1( u0_u4_u4_n158 ) , .B2( u0_u4_u4_n171 ) , .C2( u0_u4_u4_n173 ) , .A( u0_u4_u4_n94 ) , .ZN( u0_u4_u4_n95 ) );
  AOI222_X1 u0_u4_u4_U38 (.B2( u0_u4_u4_n132 ) , .A1( u0_u4_u4_n138 ) , .C2( u0_u4_u4_n175 ) , .A2( u0_u4_u4_n179 ) , .C1( u0_u4_u4_n181 ) , .B1( u0_u4_u4_n185 ) , .ZN( u0_u4_u4_n94 ) );
  INV_X1 u0_u4_u4_U39 (.A( u0_u4_u4_n113 ) , .ZN( u0_u4_u4_n185 ) );
  INV_X1 u0_u4_u4_U4 (.A( u0_u4_u4_n117 ) , .ZN( u0_u4_u4_n184 ) );
  INV_X1 u0_u4_u4_U40 (.A( u0_u4_u4_n143 ) , .ZN( u0_u4_u4_n183 ) );
  NOR2_X1 u0_u4_u4_U41 (.ZN( u0_u4_u4_n138 ) , .A1( u0_u4_u4_n168 ) , .A2( u0_u4_u4_n169 ) );
  NOR2_X1 u0_u4_u4_U42 (.A1( u0_u4_u4_n150 ) , .A2( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n153 ) );
  NOR2_X1 u0_u4_u4_U43 (.A2( u0_u4_u4_n128 ) , .A1( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n156 ) );
  AOI22_X1 u0_u4_u4_U44 (.B2( u0_u4_u4_n122 ) , .A1( u0_u4_u4_n123 ) , .ZN( u0_u4_u4_n124 ) , .B1( u0_u4_u4_n128 ) , .A2( u0_u4_u4_n172 ) );
  INV_X1 u0_u4_u4_U45 (.A( u0_u4_u4_n153 ) , .ZN( u0_u4_u4_n172 ) );
  NAND2_X1 u0_u4_u4_U46 (.A2( u0_u4_u4_n120 ) , .ZN( u0_u4_u4_n123 ) , .A1( u0_u4_u4_n161 ) );
  AOI22_X1 u0_u4_u4_U47 (.B2( u0_u4_u4_n132 ) , .A2( u0_u4_u4_n133 ) , .ZN( u0_u4_u4_n140 ) , .A1( u0_u4_u4_n150 ) , .B1( u0_u4_u4_n179 ) );
  NAND2_X1 u0_u4_u4_U48 (.ZN( u0_u4_u4_n133 ) , .A2( u0_u4_u4_n146 ) , .A1( u0_u4_u4_n154 ) );
  NAND2_X1 u0_u4_u4_U49 (.A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n154 ) , .A2( u0_u4_u4_n98 ) );
  NOR4_X1 u0_u4_u4_U5 (.A4( u0_u4_u4_n106 ) , .A3( u0_u4_u4_n107 ) , .A2( u0_u4_u4_n108 ) , .A1( u0_u4_u4_n109 ) , .ZN( u0_u4_u4_n110 ) );
  NAND2_X1 u0_u4_u4_U50 (.A1( u0_u4_u4_n101 ) , .ZN( u0_u4_u4_n158 ) , .A2( u0_u4_u4_n99 ) );
  AOI21_X1 u0_u4_u4_U51 (.ZN( u0_u4_u4_n127 ) , .A( u0_u4_u4_n136 ) , .B2( u0_u4_u4_n150 ) , .B1( u0_u4_u4_n180 ) );
  INV_X1 u0_u4_u4_U52 (.A( u0_u4_u4_n160 ) , .ZN( u0_u4_u4_n180 ) );
  NAND2_X1 u0_u4_u4_U53 (.A2( u0_u4_u4_n104 ) , .A1( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n146 ) );
  NAND2_X1 u0_u4_u4_U54 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n160 ) );
  NAND2_X1 u0_u4_u4_U55 (.ZN( u0_u4_u4_n134 ) , .A1( u0_u4_u4_n98 ) , .A2( u0_u4_u4_n99 ) );
  NAND2_X1 u0_u4_u4_U56 (.A1( u0_u4_u4_n103 ) , .A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n143 ) );
  NAND2_X1 u0_u4_u4_U57 (.A2( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n145 ) , .A1( u0_u4_u4_n98 ) );
  NAND2_X1 u0_u4_u4_U58 (.A1( u0_u4_u4_n100 ) , .A2( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n120 ) );
  NAND2_X1 u0_u4_u4_U59 (.A1( u0_u4_u4_n102 ) , .A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n148 ) );
  AOI21_X1 u0_u4_u4_U6 (.ZN( u0_u4_u4_n106 ) , .B2( u0_u4_u4_n146 ) , .B1( u0_u4_u4_n158 ) , .A( u0_u4_u4_n170 ) );
  NAND2_X1 u0_u4_u4_U60 (.A2( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n157 ) );
  INV_X1 u0_u4_u4_U61 (.A( u0_u4_u4_n150 ) , .ZN( u0_u4_u4_n173 ) );
  INV_X1 u0_u4_u4_U62 (.A( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n171 ) );
  NAND2_X1 u0_u4_u4_U63 (.A1( u0_u4_u4_n100 ) , .ZN( u0_u4_u4_n118 ) , .A2( u0_u4_u4_n99 ) );
  NAND2_X1 u0_u4_u4_U64 (.A2( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n144 ) );
  NAND2_X1 u0_u4_u4_U65 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n105 ) , .ZN( u0_u4_u4_n96 ) );
  INV_X1 u0_u4_u4_U66 (.A( u0_u4_u4_n128 ) , .ZN( u0_u4_u4_n174 ) );
  NAND2_X1 u0_u4_u4_U67 (.A2( u0_u4_u4_n102 ) , .ZN( u0_u4_u4_n119 ) , .A1( u0_u4_u4_n98 ) );
  NAND2_X1 u0_u4_u4_U68 (.A2( u0_u4_u4_n101 ) , .A1( u0_u4_u4_n103 ) , .ZN( u0_u4_u4_n147 ) );
  NAND2_X1 u0_u4_u4_U69 (.A2( u0_u4_u4_n104 ) , .ZN( u0_u4_u4_n113 ) , .A1( u0_u4_u4_n99 ) );
  AOI21_X1 u0_u4_u4_U7 (.ZN( u0_u4_u4_n108 ) , .B2( u0_u4_u4_n134 ) , .B1( u0_u4_u4_n155 ) , .A( u0_u4_u4_n156 ) );
  NOR2_X1 u0_u4_u4_U70 (.A2( u0_u4_X_28 ) , .ZN( u0_u4_u4_n150 ) , .A1( u0_u4_u4_n168 ) );
  NOR2_X1 u0_u4_u4_U71 (.A2( u0_u4_X_29 ) , .ZN( u0_u4_u4_n152 ) , .A1( u0_u4_u4_n169 ) );
  NOR2_X1 u0_u4_u4_U72 (.A2( u0_u4_X_30 ) , .ZN( u0_u4_u4_n105 ) , .A1( u0_u4_u4_n176 ) );
  NOR2_X1 u0_u4_u4_U73 (.A2( u0_u4_X_26 ) , .ZN( u0_u4_u4_n100 ) , .A1( u0_u4_u4_n177 ) );
  NOR2_X1 u0_u4_u4_U74 (.A2( u0_u4_X_28 ) , .A1( u0_u4_X_29 ) , .ZN( u0_u4_u4_n128 ) );
  NOR2_X1 u0_u4_u4_U75 (.A2( u0_u4_X_27 ) , .A1( u0_u4_X_30 ) , .ZN( u0_u4_u4_n102 ) );
  NOR2_X1 u0_u4_u4_U76 (.A2( u0_u4_X_25 ) , .A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n98 ) );
  AND2_X1 u0_u4_u4_U77 (.A2( u0_u4_X_25 ) , .A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n104 ) );
  AND2_X1 u0_u4_u4_U78 (.A1( u0_u4_X_30 ) , .A2( u0_u4_u4_n176 ) , .ZN( u0_u4_u4_n99 ) );
  AND2_X1 u0_u4_u4_U79 (.A1( u0_u4_X_26 ) , .ZN( u0_u4_u4_n101 ) , .A2( u0_u4_u4_n177 ) );
  AOI21_X1 u0_u4_u4_U8 (.ZN( u0_u4_u4_n109 ) , .A( u0_u4_u4_n153 ) , .B1( u0_u4_u4_n159 ) , .B2( u0_u4_u4_n184 ) );
  AND2_X1 u0_u4_u4_U80 (.A1( u0_u4_X_27 ) , .A2( u0_u4_X_30 ) , .ZN( u0_u4_u4_n103 ) );
  INV_X1 u0_u4_u4_U81 (.A( u0_u4_X_28 ) , .ZN( u0_u4_u4_n169 ) );
  INV_X1 u0_u4_u4_U82 (.A( u0_u4_X_29 ) , .ZN( u0_u4_u4_n168 ) );
  INV_X1 u0_u4_u4_U83 (.A( u0_u4_X_25 ) , .ZN( u0_u4_u4_n177 ) );
  INV_X1 u0_u4_u4_U84 (.A( u0_u4_X_27 ) , .ZN( u0_u4_u4_n176 ) );
  NAND4_X1 u0_u4_u4_U85 (.ZN( u0_out4_25 ) , .A4( u0_u4_u4_n139 ) , .A3( u0_u4_u4_n140 ) , .A2( u0_u4_u4_n141 ) , .A1( u0_u4_u4_n142 ) );
  OAI21_X1 u0_u4_u4_U86 (.B2( u0_u4_u4_n131 ) , .ZN( u0_u4_u4_n141 ) , .A( u0_u4_u4_n175 ) , .B1( u0_u4_u4_n183 ) );
  OAI21_X1 u0_u4_u4_U87 (.A( u0_u4_u4_n128 ) , .B2( u0_u4_u4_n129 ) , .B1( u0_u4_u4_n130 ) , .ZN( u0_u4_u4_n142 ) );
  NAND4_X1 u0_u4_u4_U88 (.ZN( u0_out4_14 ) , .A4( u0_u4_u4_n124 ) , .A3( u0_u4_u4_n125 ) , .A2( u0_u4_u4_n126 ) , .A1( u0_u4_u4_n127 ) );
  AOI22_X1 u0_u4_u4_U89 (.B2( u0_u4_u4_n117 ) , .ZN( u0_u4_u4_n126 ) , .A1( u0_u4_u4_n129 ) , .B1( u0_u4_u4_n152 ) , .A2( u0_u4_u4_n175 ) );
  AOI211_X1 u0_u4_u4_U9 (.B( u0_u4_u4_n136 ) , .A( u0_u4_u4_n137 ) , .C2( u0_u4_u4_n138 ) , .ZN( u0_u4_u4_n139 ) , .C1( u0_u4_u4_n182 ) );
  AOI22_X1 u0_u4_u4_U90 (.ZN( u0_u4_u4_n125 ) , .B2( u0_u4_u4_n131 ) , .A2( u0_u4_u4_n132 ) , .B1( u0_u4_u4_n138 ) , .A1( u0_u4_u4_n178 ) );
  NAND4_X1 u0_u4_u4_U91 (.ZN( u0_out4_8 ) , .A4( u0_u4_u4_n110 ) , .A3( u0_u4_u4_n111 ) , .A2( u0_u4_u4_n112 ) , .A1( u0_u4_u4_n186 ) );
  NAND2_X1 u0_u4_u4_U92 (.ZN( u0_u4_u4_n112 ) , .A2( u0_u4_u4_n130 ) , .A1( u0_u4_u4_n150 ) );
  AOI22_X1 u0_u4_u4_U93 (.ZN( u0_u4_u4_n111 ) , .B2( u0_u4_u4_n132 ) , .A1( u0_u4_u4_n152 ) , .B1( u0_u4_u4_n178 ) , .A2( u0_u4_u4_n97 ) );
  AOI22_X1 u0_u4_u4_U94 (.B2( u0_u4_u4_n149 ) , .B1( u0_u4_u4_n150 ) , .A2( u0_u4_u4_n151 ) , .A1( u0_u4_u4_n152 ) , .ZN( u0_u4_u4_n167 ) );
  NOR4_X1 u0_u4_u4_U95 (.A4( u0_u4_u4_n162 ) , .A3( u0_u4_u4_n163 ) , .A2( u0_u4_u4_n164 ) , .A1( u0_u4_u4_n165 ) , .ZN( u0_u4_u4_n166 ) );
  NAND3_X1 u0_u4_u4_U96 (.ZN( u0_out4_3 ) , .A3( u0_u4_u4_n166 ) , .A1( u0_u4_u4_n167 ) , .A2( u0_u4_u4_n186 ) );
  NAND3_X1 u0_u4_u4_U97 (.A3( u0_u4_u4_n146 ) , .A2( u0_u4_u4_n147 ) , .A1( u0_u4_u4_n148 ) , .ZN( u0_u4_u4_n149 ) );
  NAND3_X1 u0_u4_u4_U98 (.A3( u0_u4_u4_n143 ) , .A2( u0_u4_u4_n144 ) , .A1( u0_u4_u4_n145 ) , .ZN( u0_u4_u4_n151 ) );
  NAND3_X1 u0_u4_u4_U99 (.A3( u0_u4_u4_n121 ) , .ZN( u0_u4_u4_n122 ) , .A2( u0_u4_u4_n144 ) , .A1( u0_u4_u4_n154 ) );
  OAI21_X1 u0_uk_U104 (.ZN( u0_K4_5 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n502 ) , .A( u0_uk_n821 ) );
  NAND2_X1 u0_uk_U105 (.A1( u0_uk_K_r2_53 ) , .ZN( u0_uk_n821 ) , .A2( u0_uk_n99 ) );
  INV_X1 u0_uk_U1066 (.A( u0_key_r_33 ) , .ZN( u0_uk_n691 ) );
  INV_X1 u0_uk_U1135 (.ZN( u0_K4_2 ) , .A( u0_uk_n828 ) );
  AOI22_X1 u0_uk_U1136 (.B2( u0_uk_K_r2_26 ) , .A2( u0_uk_K_r2_46 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n148 ) , .ZN( u0_uk_n828 ) );
  INV_X1 u0_uk_U1137 (.ZN( u0_K4_20 ) , .A( u0_uk_n835 ) );
  AOI22_X1 u0_uk_U1138 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_33 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n208 ) , .ZN( u0_uk_n835 ) );
  NAND2_X1 u0_uk_U125 (.A1( u0_uk_K_r0_52 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n856 ) );
  OAI22_X1 u0_uk_U127 (.ZN( u0_K4_15 ) , .A1( u0_uk_n242 ) , .A2( u0_uk_n502 ) , .B2( u0_uk_n530 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U139 (.ZN( u0_K11_15 ) , .A1( u0_uk_n147 ) , .A2( u0_uk_n197 ) , .B2( u0_uk_n212 ) , .B1( u0_uk_n93 ) );
  INV_X1 u0_uk_U151 (.ZN( u0_K11_19 ) , .A( u0_uk_n1000 ) );
  AOI22_X1 u0_uk_U152 (.B2( u0_uk_K_r9_10 ) , .A2( u0_uk_K_r9_48 ) , .ZN( u0_uk_n1000 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n220 ) );
  OAI22_X1 u0_uk_U156 (.ZN( u0_K4_19 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n511 ) , .B2( u0_uk_n523 ) );
  OAI22_X1 u0_uk_U164 (.ZN( u0_K5_30 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n463 ) , .B2( u0_uk_n480 ) );
  NAND2_X1 u0_uk_U171 (.A1( u0_key_r_18 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n889 ) );
  INV_X1 u0_uk_U180 (.ZN( u0_K11_14 ) , .A( u0_uk_n1002 ) );
  INV_X1 u0_uk_U207 (.ZN( u0_K15_30 ) , .A( u0_uk_n919 ) );
  AOI22_X1 u0_uk_U208 (.B2( u0_uk_K_r13_0 ) , .A2( u0_uk_K_r13_38 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n919 ) );
  OAI22_X1 u0_uk_U236 (.ZN( u0_K15_39 ) , .A1( u0_uk_n128 ) , .B2( u0_uk_n22 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n40 ) );
  OAI22_X1 u0_uk_U244 (.ZN( u0_K15_44 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n22 ) , .A2( u0_uk_n4 ) );
  OAI21_X1 u0_uk_U245 (.ZN( u0_K15_48 ) , .B1( u0_uk_n27 ) , .B2( u0_uk_n34 ) , .A( u0_uk_n914 ) );
  NAND2_X1 u0_uk_U246 (.A1( u0_uk_K_r13_35 ) , .A2( u0_uk_n10 ) , .ZN( u0_uk_n914 ) );
  INV_X1 u0_uk_U291 (.ZN( u0_K4_8 ) , .A( u0_uk_n819 ) );
  AOI22_X1 u0_uk_U292 (.B2( u0_uk_K_r2_41 ) , .A2( u0_uk_K_r2_46 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n819 ) );
  INV_X1 u0_uk_U304 (.ZN( u0_K15_26 ) , .A( u0_uk_n920 ) );
  AOI22_X1 u0_uk_U305 (.B2( u0_uk_K_r13_38 ) , .A2( u0_uk_K_r13_44 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n920 ) );
  OAI22_X1 u0_uk_U320 (.ZN( u0_K15_46 ) , .B2( u0_uk_n13 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .A2( u0_uk_n40 ) );
  OAI22_X1 u0_uk_U337 (.ZN( u0_K15_4 ) , .A1( u0_uk_n100 ) , .B1( u0_uk_n222 ) , .B2( u0_uk_n38 ) , .A2( u0_uk_n8 ) );
  INV_X1 u0_uk_U345 (.ZN( u0_K4_4 ) , .A( u0_uk_n822 ) );
  AOI22_X1 u0_uk_U346 (.B2( u0_uk_K_r2_13 ) , .A2( u0_uk_K_r2_18 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n822 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U360 (.ZN( u0_K15_40 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n41 ) , .B2( u0_uk_n9 ) );
  OAI22_X1 u0_uk_U381 (.ZN( u0_K15_28 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n230 ) , .B2( u0_uk_n33 ) , .A2( u0_uk_n5 ) );
  OAI22_X1 u0_uk_U401 (.ZN( u0_K4_16 ) , .B1( u0_uk_n128 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n525 ) , .B2( u0_uk_n529 ) );
  OAI22_X1 u0_uk_U421 (.ZN( u0_K4_9 ) , .A1( u0_uk_n146 ) , .B1( u0_uk_n217 ) , .A2( u0_uk_n519 ) , .B2( u0_uk_n529 ) );
  OAI22_X1 u0_uk_U425 (.ZN( u0_K15_1 ) , .A2( u0_uk_n1 ) , .B2( u0_uk_n20 ) , .A1( u0_uk_n230 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U454 (.ZN( u0_K15_37 ) , .B2( u0_uk_n12 ) , .A1( u0_uk_n187 ) , .B1( u0_uk_n27 ) , .A2( u0_uk_n39 ) );
  NAND2_X1 u0_uk_U458 (.A1( u0_uk_K_r9_38 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n989 ) );
  OAI22_X1 u0_uk_U482 (.ZN( u0_K15_29 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n21 ) , .A2( u0_uk_n39 ) );
  OAI22_X1 u0_uk_U487 (.ZN( u0_K5_29 ) , .A1( u0_uk_n118 ) , .B1( u0_uk_n222 ) , .A2( u0_uk_n462 ) , .B2( u0_uk_n481 ) );
  INV_X1 u0_uk_U508 (.ZN( u0_K11_17 ) , .A( u0_uk_n1001 ) );
  OAI21_X1 u0_uk_U513 (.ZN( u0_K4_17 ) , .B1( u0_uk_n250 ) , .B2( u0_uk_n519 ) , .A( u0_uk_n838 ) );
  NAND2_X1 u0_uk_U514 (.A1( u0_uk_K_r2_27 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n838 ) );
  OAI22_X1 u0_uk_U526 (.ZN( u0_K4_12 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n161 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n517 ) );
  OAI22_X1 u0_uk_U529 (.ZN( u0_K15_2 ) , .A2( u0_uk_n1 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n30 ) );
  INV_X1 u0_uk_U562 (.ZN( u0_K15_38 ) , .A( u0_uk_n916 ) );
  INV_X1 u0_uk_U584 (.ZN( u0_K4_10 ) , .A( u0_uk_n839 ) );
  INV_X1 u0_uk_U592 (.ZN( u0_K11_22 ) , .A( u0_uk_n997 ) );
  AOI22_X1 u0_uk_U593 (.B2( u0_uk_K_r9_13 ) , .A2( u0_uk_K_r9_19 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n251 ) , .ZN( u0_uk_n997 ) );
  INV_X1 u0_uk_U643 (.ZN( u0_K4_23 ) , .A( u0_uk_n833 ) );
  AOI22_X1 u0_uk_U644 (.B2( u0_uk_K_r2_18 ) , .A2( u0_uk_K_r2_55 ) , .B1( u0_uk_n207 ) , .ZN( u0_uk_n833 ) , .A1( u0_uk_n94 ) );
  INV_X1 u0_uk_U649 (.A( u0_key_r_44 ) , .ZN( u0_uk_n680 ) );
  INV_X1 u0_uk_U660 (.ZN( u0_K15_43 ) , .A( u0_uk_n915 ) );
  AOI22_X1 u0_uk_U661 (.A2( u0_uk_K_r13_2 ) , .B2( u0_uk_K_r13_23 ) , .A1( u0_uk_n163 ) , .ZN( u0_uk_n915 ) , .B1( u0_uk_n93 ) );
  OAI22_X1 u0_uk_U684 (.ZN( u0_K4_7 ) , .B1( u0_uk_n202 ) , .B2( u0_uk_n531 ) , .A2( u0_uk_n535 ) , .A1( u0_uk_n99 ) );
  OAI21_X1 u0_uk_U686 (.ZN( u0_K15_25 ) , .B2( u0_uk_n12 ) , .B1( u0_uk_n147 ) , .A( u0_uk_n921 ) );
  NAND2_X1 u0_uk_U687 (.A1( u0_uk_K_r13_22 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n921 ) );
  OAI21_X1 u0_uk_U690 (.ZN( u0_K5_25 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n475 ) , .A( u0_uk_n814 ) );
  NAND2_X1 u0_uk_U691 (.A1( u0_uk_K_r3_35 ) , .A2( u0_uk_n128 ) , .ZN( u0_uk_n814 ) );
  INV_X1 u0_uk_U702 (.ZN( u0_K4_3 ) , .A( u0_uk_n824 ) );
  AOI22_X1 u0_uk_U703 (.A2( u0_uk_K_r2_4 ) , .B2( u0_uk_K_r2_41 ) , .A1( u0_uk_n238 ) , .ZN( u0_uk_n824 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U726 (.ZN( u0_K15_42 ) , .A1( u0_uk_n141 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n3 ) , .B2( u0_uk_n9 ) );
  OAI21_X1 u0_uk_U75 (.ZN( u0_K11_23 ) , .B2( u0_uk_n190 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n996 ) );
  OAI22_X1 u0_uk_U752 (.ZN( u0_K11_13 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n164 ) , .A2( u0_uk_n196 ) , .B2( u0_uk_n200 ) );
  NAND2_X1 u0_uk_U76 (.A1( u0_uk_K_r9_27 ) , .A2( u0_uk_n202 ) , .ZN( u0_uk_n996 ) );
  NAND2_X1 u0_uk_U763 (.A1( u0_uk_K_r9_5 ) , .A2( u0_uk_n17 ) , .ZN( u0_uk_n998 ) );
  OAI22_X1 u0_uk_U766 (.ZN( u0_K4_21 ) , .B1( u0_uk_n146 ) , .A1( u0_uk_n238 ) , .A2( u0_uk_n511 ) , .B2( u0_uk_n517 ) );
  OAI22_X1 u0_uk_U771 (.ZN( u0_K15_27 ) , .A1( u0_uk_n128 ) , .B1( u0_uk_n188 ) , .B2( u0_uk_n23 ) , .A2( u0_uk_n41 ) );
  OAI22_X1 u0_uk_U772 (.ZN( u0_K4_13 ) , .B1( u0_uk_n240 ) , .B2( u0_uk_n530 ) , .A2( u0_uk_n534 ) , .A1( u0_uk_n60 ) );
  INV_X1 u0_uk_U774 (.ZN( u0_K5_27 ) , .A( u0_uk_n813 ) );
  OAI21_X1 u0_uk_U802 (.ZN( u0_K4_1 ) , .B1( u0_uk_n252 ) , .B2( u0_uk_n535 ) , .A( u0_uk_n836 ) );
  NAND2_X1 u0_uk_U803 (.A1( u0_uk_K_r2_25 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n836 ) );
  OAI21_X1 u0_uk_U804 (.ZN( u0_K4_18 ) , .B2( u0_uk_n510 ) , .A( u0_uk_n837 ) , .B1( u0_uk_n92 ) );
  NAND2_X1 u0_uk_U805 (.A1( u0_uk_K_r2_20 ) , .A2( u0_uk_n31 ) , .ZN( u0_uk_n837 ) );
  INV_X1 u0_uk_U829 (.ZN( u0_K11_20 ) , .A( u0_uk_n999 ) );
  OAI21_X1 u0_uk_U838 (.ZN( u0_K4_22 ) , .B2( u0_uk_n531 ) , .B1( u0_uk_n60 ) , .A( u0_uk_n834 ) );
  OAI22_X1 u0_uk_U842 (.ZN( u0_K15_6 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n24 ) , .A2( u0_uk_n6 ) );
  OAI22_X1 u0_uk_U850 (.ZN( u0_K15_3 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .A2( u0_uk_n20 ) , .B2( u0_uk_n36 ) );
  OAI22_X1 u0_uk_U88 (.ZN( u0_K15_41 ) , .B1( u0_uk_n17 ) , .A1( u0_uk_n187 ) , .B2( u0_uk_n23 ) , .A2( u0_uk_n5 ) );
  OAI22_X1 u0_uk_U884 (.ZN( u0_K4_11 ) , .B1( u0_uk_n117 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n497 ) , .B2( u0_uk_n525 ) );
  OAI22_X1 u0_uk_U886 (.ZN( u0_K15_45 ) , .A1( u0_uk_n155 ) , .B1( u0_uk_n17 ) , .B2( u0_uk_n21 ) , .A2( u0_uk_n3 ) );
  OAI22_X1 u0_uk_U914 (.ZN( u0_K4_14 ) , .A1( u0_uk_n164 ) , .A2( u0_uk_n510 ) , .B2( u0_uk_n536 ) , .B1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U933 (.ZN( u0_K11_16 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n190 ) , .B2( u0_uk_n196 ) );
  OAI22_X1 u0_uk_U942 (.ZN( u0_K11_24 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n201 ) , .B2( u0_uk_n206 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U95 (.ZN( u0_K15_5 ) , .B1( u0_uk_n220 ) , .A2( u0_uk_n26 ) , .B2( u0_uk_n29 ) , .A1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U959 (.ZN( u0_K11_18 ) , .A1( u0_uk_n110 ) , .B1( u0_uk_n214 ) , .A2( u0_uk_n215 ) , .B2( u0_uk_n221 ) );
  XOR2_X1 u1_U100 (.B( u1_L12_27 ) , .Z( u1_N442 ) , .A( u1_out13_27 ) );
  XOR2_X1 u1_U102 (.B( u1_L12_25 ) , .Z( u1_N440 ) , .A( u1_out13_25 ) );
  XOR2_X1 u1_U106 (.B( u1_L12_22 ) , .Z( u1_N437 ) , .A( u1_out13_22 ) );
  XOR2_X1 u1_U107 (.B( u1_L12_21 ) , .Z( u1_N436 ) , .A( u1_out13_21 ) );
  XOR2_X1 u1_U110 (.B( u1_L12_18 ) , .Z( u1_N433 ) , .A( u1_out13_18 ) );
  XOR2_X1 u1_U113 (.B( u1_L12_15 ) , .Z( u1_N430 ) , .A( u1_out13_15 ) );
  XOR2_X1 u1_U114 (.B( u1_L0_12 ) , .Z( u1_N43 ) , .A( u1_out1_12 ) );
  XOR2_X1 u1_U115 (.B( u1_L12_14 ) , .Z( u1_N429 ) , .A( u1_out13_14 ) );
  XOR2_X1 u1_U116 (.B( u1_L12_13 ) , .Z( u1_N428 ) , .A( u1_out13_13 ) );
  XOR2_X1 u1_U117 (.B( u1_L12_12 ) , .Z( u1_N427 ) , .A( u1_out13_12 ) );
  XOR2_X1 u1_U12 (.B( u1_L1_27 ) , .Z( u1_N90 ) , .A( u1_out2_27 ) );
  XOR2_X1 u1_U121 (.B( u1_L12_8 ) , .Z( u1_N423 ) , .A( u1_out13_8 ) );
  XOR2_X1 u1_U122 (.B( u1_L12_7 ) , .Z( u1_N422 ) , .A( u1_out13_7 ) );
  XOR2_X1 u1_U124 (.B( u1_L12_5 ) , .Z( u1_N420 ) , .A( u1_out13_5 ) );
  XOR2_X1 u1_U127 (.B( u1_L12_3 ) , .Z( u1_N418 ) , .A( u1_out13_3 ) );
  XOR2_X1 u1_U128 (.B( u1_L12_2 ) , .Z( u1_N417 ) , .A( u1_out13_2 ) );
  XOR2_X1 u1_U13 (.Z( u1_N9 ) , .B( u1_desIn_r_12 ) , .A( u1_out0_10 ) );
  XOR2_X1 u1_U131 (.B( u1_L11_31 ) , .Z( u1_N414 ) , .A( u1_out12_31 ) );
  XOR2_X1 u1_U136 (.B( u1_L0_10 ) , .Z( u1_N41 ) , .A( u1_out1_10 ) );
  XOR2_X1 u1_U137 (.B( u1_L11_26 ) , .Z( u1_N409 ) , .A( u1_out12_26 ) );
  XOR2_X1 u1_U138 (.B( u1_L11_25 ) , .Z( u1_N408 ) , .A( u1_out12_25 ) );
  XOR2_X1 u1_U14 (.B( u1_L1_26 ) , .Z( u1_N89 ) , .A( u1_out2_26 ) );
  XOR2_X1 u1_U140 (.B( u1_L11_23 ) , .Z( u1_N406 ) , .A( u1_out12_23 ) );
  XOR2_X1 u1_U143 (.B( u1_L11_20 ) , .Z( u1_N403 ) , .A( u1_out12_20 ) );
  XOR2_X1 u1_U146 (.B( u1_L11_17 ) , .Z( u1_N400 ) , .A( u1_out12_17 ) );
  XOR2_X1 u1_U147 (.B( u1_L0_9 ) , .Z( u1_N40 ) , .A( u1_out1_9 ) );
  XOR2_X1 u1_U148 (.Z( u1_N4 ) , .B( u1_desIn_r_38 ) , .A( u1_out0_5 ) );
  XOR2_X1 u1_U151 (.B( u1_L11_14 ) , .Z( u1_N397 ) , .A( u1_out12_14 ) );
  XOR2_X1 u1_U155 (.B( u1_L11_10 ) , .Z( u1_N393 ) , .A( u1_out12_10 ) );
  XOR2_X1 u1_U156 (.B( u1_L11_9 ) , .Z( u1_N392 ) , .A( u1_out12_9 ) );
  XOR2_X1 u1_U157 (.B( u1_L11_8 ) , .Z( u1_N391 ) , .A( u1_out12_8 ) );
  XOR2_X1 u1_U159 (.B( u1_L0_8 ) , .Z( u1_N39 ) , .A( u1_out1_8 ) );
  XOR2_X1 u1_U163 (.B( u1_L11_3 ) , .Z( u1_N386 ) , .A( u1_out12_3 ) );
  XOR2_X1 u1_U165 (.B( u1_L11_1 ) , .Z( u1_N384 ) , .A( u1_out12_1 ) );
  XOR2_X1 u1_U168 (.B( u1_L10_30 ) , .Z( u1_N381 ) , .A( u1_out11_30 ) );
  XOR2_X1 u1_U170 (.B( u1_L0_7 ) , .Z( u1_N38 ) , .A( u1_out1_7 ) );
  XOR2_X1 u1_U171 (.B( u1_L10_28 ) , .Z( u1_N379 ) , .A( u1_out11_28 ) );
  XOR2_X1 u1_U173 (.B( u1_L10_26 ) , .Z( u1_N377 ) , .A( u1_out11_26 ) );
  XOR2_X1 u1_U174 (.B( u1_L10_25 ) , .Z( u1_N376 ) , .A( u1_out11_25 ) );
  XOR2_X1 u1_U175 (.B( u1_L10_24 ) , .Z( u1_N375 ) , .A( u1_out11_24 ) );
  XOR2_X1 u1_U179 (.B( u1_L10_20 ) , .Z( u1_N371 ) , .A( u1_out11_20 ) );
  XOR2_X1 u1_U181 (.B( u1_L0_6 ) , .Z( u1_N37 ) , .A( u1_out1_6 ) );
  XOR2_X1 u1_U182 (.B( u1_L10_18 ) , .Z( u1_N369 ) , .A( u1_out11_18 ) );
  XOR2_X1 u1_U184 (.B( u1_L10_16 ) , .Z( u1_N367 ) , .A( u1_out11_16 ) );
  XOR2_X1 u1_U186 (.B( u1_L10_14 ) , .Z( u1_N365 ) , .A( u1_out11_14 ) );
  XOR2_X1 u1_U187 (.B( u1_L10_13 ) , .Z( u1_N364 ) , .A( u1_out11_13 ) );
  XOR2_X1 u1_U19 (.B( u1_L1_21 ) , .Z( u1_N84 ) , .A( u1_out2_21 ) );
  XOR2_X1 u1_U190 (.B( u1_L10_10 ) , .Z( u1_N361 ) , .A( u1_out11_10 ) );
  XOR2_X1 u1_U192 (.B( u1_L0_5 ) , .Z( u1_N36 ) , .A( u1_out1_5 ) );
  XOR2_X1 u1_U193 (.B( u1_L10_8 ) , .Z( u1_N359 ) , .A( u1_out11_8 ) );
  XOR2_X1 u1_U195 (.B( u1_L10_6 ) , .Z( u1_N357 ) , .A( u1_out11_6 ) );
  XOR2_X1 u1_U198 (.B( u1_L10_3 ) , .Z( u1_N354 ) , .A( u1_out11_3 ) );
  XOR2_X1 u1_U199 (.B( u1_L10_2 ) , .Z( u1_N353 ) , .A( u1_out11_2 ) );
  XOR2_X1 u1_U20 (.B( u1_L1_20 ) , .Z( u1_N83 ) , .A( u1_out2_20 ) );
  XOR2_X1 u1_U200 (.B( u1_L10_1 ) , .Z( u1_N352 ) , .A( u1_out11_1 ) );
  XOR2_X1 u1_U201 (.B( u1_L9_32 ) , .Z( u1_N351 ) , .A( u1_out10_32 ) );
  XOR2_X1 u1_U212 (.B( u1_L9_22 ) , .Z( u1_N341 ) , .A( u1_out10_22 ) );
  XOR2_X1 u1_U214 (.B( u1_L0_3 ) , .Z( u1_N34 ) , .A( u1_out1_3 ) );
  XOR2_X1 u1_U223 (.B( u1_L9_12 ) , .Z( u1_N331 ) , .A( u1_out10_12 ) );
  XOR2_X1 u1_U229 (.B( u1_L9_7 ) , .Z( u1_N326 ) , .A( u1_out10_7 ) );
  XOR2_X1 u1_U236 (.B( u1_L0_1 ) , .Z( u1_N32 ) , .A( u1_out1_1 ) );
  XOR2_X1 u1_U238 (.B( u1_L8_31 ) , .Z( u1_N318 ) , .A( u1_out9_31 ) );
  XOR2_X1 u1_U24 (.Z( u1_N8 ) , .B( u1_desIn_r_4 ) , .A( u1_out0_9 ) );
  XOR2_X1 u1_U242 (.B( u1_L8_27 ) , .Z( u1_N314 ) , .A( u1_out9_27 ) );
  XOR2_X1 u1_U246 (.B( u1_L8_23 ) , .Z( u1_N310 ) , .A( u1_out9_23 ) );
  XOR2_X1 u1_U247 (.Z( u1_N31 ) , .B( u1_desIn_r_56 ) , .A( u1_out0_32 ) );
  XOR2_X1 u1_U249 (.B( u1_L8_21 ) , .Z( u1_N308 ) , .A( u1_out9_21 ) );
  XOR2_X1 u1_U253 (.B( u1_L8_17 ) , .Z( u1_N304 ) , .A( u1_out9_17 ) );
  XOR2_X1 u1_U255 (.B( u1_L8_15 ) , .Z( u1_N302 ) , .A( u1_out9_15 ) );
  XOR2_X1 u1_U258 (.Z( u1_N30 ) , .B( u1_desIn_r_48 ) , .A( u1_out0_31 ) );
  XOR2_X1 u1_U26 (.B( u1_L1_15 ) , .Z( u1_N78 ) , .A( u1_out2_15 ) );
  XOR2_X1 u1_U263 (.B( u1_L8_9 ) , .Z( u1_N296 ) , .A( u1_out9_9 ) );
  XOR2_X1 u1_U267 (.B( u1_L8_5 ) , .Z( u1_N292 ) , .A( u1_out9_5 ) );
  XOR2_X1 u1_U273 (.B( u1_L7_32 ) , .Z( u1_N287 ) , .A( u1_out8_32 ) );
  XOR2_X1 u1_U275 (.B( u1_L7_30 ) , .Z( u1_N285 ) , .A( u1_out8_30 ) );
  XOR2_X1 u1_U277 (.B( u1_L7_28 ) , .Z( u1_N283 ) , .A( u1_out8_28 ) );
  XOR2_X1 u1_U278 (.B( u1_L7_27 ) , .Z( u1_N282 ) , .A( u1_out8_27 ) );
  XOR2_X1 u1_U279 (.B( u1_L7_26 ) , .Z( u1_N281 ) , .A( u1_out8_26 ) );
  XOR2_X1 u1_U282 (.B( u1_L7_24 ) , .Z( u1_N279 ) , .A( u1_out8_24 ) );
  XOR2_X1 u1_U284 (.B( u1_L7_22 ) , .Z( u1_N277 ) , .A( u1_out8_22 ) );
  XOR2_X1 u1_U285 (.B( u1_L7_21 ) , .Z( u1_N276 ) , .A( u1_out8_21 ) );
  XOR2_X1 u1_U286 (.B( u1_L7_20 ) , .Z( u1_N275 ) , .A( u1_out8_20 ) );
  XOR2_X1 u1_U288 (.B( u1_L7_18 ) , .Z( u1_N273 ) , .A( u1_out8_18 ) );
  XOR2_X1 u1_U290 (.B( u1_L7_16 ) , .Z( u1_N271 ) , .A( u1_out8_16 ) );
  XOR2_X1 u1_U291 (.B( u1_L7_15 ) , .Z( u1_N270 ) , .A( u1_out8_15 ) );
  XOR2_X1 u1_U292 (.Z( u1_N27 ) , .B( u1_desIn_r_24 ) , .A( u1_out0_28 ) );
  XOR2_X1 u1_U294 (.B( u1_L7_13 ) , .Z( u1_N268 ) , .A( u1_out8_13 ) );
  XOR2_X1 u1_U295 (.B( u1_L7_12 ) , .Z( u1_N267 ) , .A( u1_out8_12 ) );
  XOR2_X1 u1_U297 (.B( u1_L7_10 ) , .Z( u1_N265 ) , .A( u1_out8_10 ) );
  XOR2_X1 u1_U300 (.B( u1_L7_7 ) , .Z( u1_N262 ) , .A( u1_out8_7 ) );
  XOR2_X1 u1_U301 (.B( u1_L7_6 ) , .Z( u1_N261 ) , .A( u1_out8_6 ) );
  XOR2_X1 u1_U302 (.B( u1_L7_5 ) , .Z( u1_N260 ) , .A( u1_out8_5 ) );
  XOR2_X1 u1_U303 (.Z( u1_N26 ) , .B( u1_desIn_r_16 ) , .A( u1_out0_27 ) );
  XOR2_X1 u1_U306 (.B( u1_L7_2 ) , .Z( u1_N257 ) , .A( u1_out8_2 ) );
  XOR2_X1 u1_U307 (.B( u1_L7_1 ) , .Z( u1_N256 ) , .A( u1_out8_1 ) );
  XOR2_X1 u1_U308 (.B( u1_L6_32 ) , .Z( u1_N255 ) , .A( u1_out7_32 ) );
  XOR2_X1 u1_U309 (.B( u1_L6_31 ) , .Z( u1_N254 ) , .A( u1_out7_31 ) );
  XOR2_X1 u1_U31 (.B( u1_L1_10 ) , .Z( u1_N73 ) , .A( u1_out2_10 ) );
  XOR2_X1 u1_U310 (.B( u1_L6_30 ) , .Z( u1_N253 ) , .A( u1_out7_30 ) );
  XOR2_X1 u1_U312 (.B( u1_L6_28 ) , .Z( u1_N251 ) , .A( u1_out7_28 ) );
  XOR2_X1 u1_U314 (.Z( u1_N25 ) , .B( u1_desIn_r_8 ) , .A( u1_out0_26 ) );
  XOR2_X1 u1_U316 (.B( u1_L6_25 ) , .Z( u1_N248 ) , .A( u1_out7_25 ) );
  XOR2_X1 u1_U317 (.B( u1_L6_24 ) , .Z( u1_N247 ) , .A( u1_out7_24 ) );
  XOR2_X1 u1_U318 (.B( u1_L6_23 ) , .Z( u1_N246 ) , .A( u1_out7_23 ) );
  XOR2_X1 u1_U319 (.B( u1_L6_22 ) , .Z( u1_N245 ) , .A( u1_out7_22 ) );
  XOR2_X1 u1_U323 (.B( u1_L6_18 ) , .Z( u1_N241 ) , .A( u1_out7_18 ) );
  XOR2_X1 u1_U324 (.B( u1_L6_17 ) , .Z( u1_N240 ) , .A( u1_out7_17 ) );
  XOR2_X1 u1_U326 (.B( u1_L6_16 ) , .Z( u1_N239 ) , .A( u1_out7_16 ) );
  XOR2_X1 u1_U328 (.B( u1_L6_14 ) , .Z( u1_N237 ) , .A( u1_out7_14 ) );
  XOR2_X1 u1_U329 (.B( u1_L6_13 ) , .Z( u1_N236 ) , .A( u1_out7_13 ) );
  XOR2_X1 u1_U330 (.B( u1_L6_12 ) , .Z( u1_N235 ) , .A( u1_out7_12 ) );
  XOR2_X1 u1_U333 (.B( u1_L6_9 ) , .Z( u1_N232 ) , .A( u1_out7_9 ) );
  XOR2_X1 u1_U334 (.B( u1_L6_8 ) , .Z( u1_N231 ) , .A( u1_out7_8 ) );
  XOR2_X1 u1_U335 (.B( u1_L6_7 ) , .Z( u1_N230 ) , .A( u1_out7_7 ) );
  XOR2_X1 u1_U337 (.B( u1_L6_6 ) , .Z( u1_N229 ) , .A( u1_out7_6 ) );
  XOR2_X1 u1_U340 (.B( u1_L6_3 ) , .Z( u1_N226 ) , .A( u1_out7_3 ) );
  XOR2_X1 u1_U341 (.B( u1_L6_2 ) , .Z( u1_N225 ) , .A( u1_out7_2 ) );
  XOR2_X1 u1_U345 (.B( u1_L5_30 ) , .Z( u1_N221 ) , .A( u1_out6_30 ) );
  XOR2_X1 u1_U347 (.Z( u1_N22 ) , .B( u1_desIn_r_50 ) , .A( u1_out0_23 ) );
  XOR2_X1 u1_U350 (.B( u1_L5_26 ) , .Z( u1_N217 ) , .A( u1_out6_26 ) );
  XOR2_X1 u1_U352 (.B( u1_L5_24 ) , .Z( u1_N215 ) , .A( u1_out6_24 ) );
  XOR2_X1 u1_U356 (.B( u1_L5_20 ) , .Z( u1_N211 ) , .A( u1_out6_20 ) );
  XOR2_X1 u1_U358 (.Z( u1_N21 ) , .B( u1_desIn_r_42 ) , .A( u1_out0_22 ) );
  XOR2_X1 u1_U361 (.B( u1_L5_16 ) , .Z( u1_N207 ) , .A( u1_out6_16 ) );
  XOR2_X1 u1_U367 (.B( u1_L5_10 ) , .Z( u1_N201 ) , .A( u1_out6_10 ) );
  XOR2_X1 u1_U369 (.Z( u1_N20 ) , .B( u1_desIn_r_34 ) , .A( u1_out0_21 ) );
  XOR2_X1 u1_U37 (.B( u1_L1_5 ) , .Z( u1_N68 ) , .A( u1_out2_5 ) );
  XOR2_X1 u1_U373 (.B( u1_L5_6 ) , .Z( u1_N197 ) , .A( u1_out6_6 ) );
  XOR2_X1 u1_U378 (.B( u1_L5_1 ) , .Z( u1_N192 ) , .A( u1_out6_1 ) );
  XOR2_X1 u1_U379 (.B( u1_L4_32 ) , .Z( u1_N191 ) , .A( u1_out5_32 ) );
  XOR2_X1 u1_U380 (.B( u1_L4_31 ) , .Z( u1_N190 ) , .A( u1_out5_31 ) );
  XOR2_X1 u1_U381 (.Z( u1_N19 ) , .B( u1_desIn_r_26 ) , .A( u1_out0_20 ) );
  XOR2_X1 u1_U382 (.B( u1_L4_30 ) , .Z( u1_N189 ) , .A( u1_out5_30 ) );
  XOR2_X1 u1_U386 (.B( u1_L4_26 ) , .Z( u1_N185 ) , .A( u1_out5_26 ) );
  XOR2_X1 u1_U388 (.B( u1_L4_24 ) , .Z( u1_N183 ) , .A( u1_out5_24 ) );
  XOR2_X1 u1_U389 (.B( u1_L4_23 ) , .Z( u1_N182 ) , .A( u1_out5_23 ) );
  XOR2_X1 u1_U390 (.B( u1_L4_22 ) , .Z( u1_N181 ) , .A( u1_out5_22 ) );
  XOR2_X1 u1_U393 (.B( u1_L4_20 ) , .Z( u1_N179 ) , .A( u1_out5_20 ) );
  XOR2_X1 u1_U396 (.B( u1_L4_17 ) , .Z( u1_N176 ) , .A( u1_out5_17 ) );
  XOR2_X1 u1_U397 (.B( u1_L4_16 ) , .Z( u1_N175 ) , .A( u1_out5_16 ) );
  XOR2_X1 u1_U401 (.B( u1_L4_12 ) , .Z( u1_N171 ) , .A( u1_out5_12 ) );
  XOR2_X1 u1_U403 (.Z( u1_N17 ) , .B( u1_desIn_r_10 ) , .A( u1_out0_18 ) );
  XOR2_X1 u1_U404 (.B( u1_L4_10 ) , .Z( u1_N169 ) , .A( u1_out5_10 ) );
  XOR2_X1 u1_U405 (.B( u1_L4_9 ) , .Z( u1_N168 ) , .A( u1_out5_9 ) );
  XOR2_X1 u1_U407 (.B( u1_L4_7 ) , .Z( u1_N166 ) , .A( u1_out5_7 ) );
  XOR2_X1 u1_U408 (.B( u1_L4_6 ) , .Z( u1_N165 ) , .A( u1_out5_6 ) );
  XOR2_X1 u1_U41 (.B( u1_L1_1 ) , .Z( u1_N64 ) , .A( u1_out2_1 ) );
  XOR2_X1 u1_U413 (.B( u1_L4_1 ) , .Z( u1_N160 ) , .A( u1_out5_1 ) );
  XOR2_X1 u1_U414 (.Z( u1_N16 ) , .B( u1_desIn_r_2 ) , .A( u1_out0_17 ) );
  XOR2_X1 u1_U418 (.B( u1_L3_29 ) , .Z( u1_N156 ) , .A( u1_out4_29 ) );
  XOR2_X1 u1_U42 (.B( u1_L0_32 ) , .Z( u1_N63 ) , .A( u1_out1_32 ) );
  XOR2_X1 u1_U420 (.B( u1_L3_27 ) , .Z( u1_N154 ) , .A( u1_out4_27 ) );
  XOR2_X1 u1_U427 (.B( u1_L3_21 ) , .Z( u1_N148 ) , .A( u1_out4_21 ) );
  XOR2_X1 u1_U429 (.B( u1_L3_19 ) , .Z( u1_N146 ) , .A( u1_out4_19 ) );
  XOR2_X1 u1_U43 (.B( u1_L0_31 ) , .Z( u1_N62 ) , .A( u1_out1_31 ) );
  XOR2_X1 u1_U433 (.B( u1_L3_15 ) , .Z( u1_N142 ) , .A( u1_out4_15 ) );
  XOR2_X1 u1_U436 (.Z( u1_N14 ) , .B( u1_desIn_r_52 ) , .A( u1_out0_15 ) );
  XOR2_X1 u1_U438 (.B( u1_L3_11 ) , .Z( u1_N138 ) , .A( u1_out4_11 ) );
  XOR2_X1 u1_U44 (.B( u1_L0_30 ) , .Z( u1_N61 ) , .A( u1_out1_30 ) );
  XOR2_X1 u1_U444 (.B( u1_L3_5 ) , .Z( u1_N132 ) , .A( u1_out4_5 ) );
  XOR2_X1 u1_U445 (.B( u1_L3_4 ) , .Z( u1_N131 ) , .A( u1_out4_4 ) );
  XOR2_X1 u1_U456 (.B( u1_L2_26 ) , .Z( u1_N121 ) , .A( u1_out3_26 ) );
  XOR2_X1 u1_U458 (.Z( u1_N12 ) , .B( u1_desIn_r_36 ) , .A( u1_out0_13 ) );
  XOR2_X1 u1_U46 (.Z( u1_N6 ) , .B( u1_desIn_r_54 ) , .A( u1_out0_7 ) );
  XOR2_X1 u1_U463 (.B( u1_L2_20 ) , .Z( u1_N115 ) , .A( u1_out3_20 ) );
  XOR2_X1 u1_U469 (.Z( u1_N11 ) , .B( u1_desIn_r_28 ) , .A( u1_out0_12 ) );
  XOR2_X1 u1_U474 (.B( u1_L2_10 ) , .Z( u1_N105 ) , .A( u1_out3_10 ) );
  XOR2_X1 u1_U48 (.B( u1_L0_27 ) , .Z( u1_N58 ) , .A( u1_out1_27 ) );
  XOR2_X1 u1_U481 (.Z( u1_N1 ) , .B( u1_desIn_r_14 ) , .A( u1_out0_2 ) );
  XOR2_X1 u1_U482 (.Z( u1_N0 ) , .B( u1_desIn_r_6 ) , .A( u1_out0_1 ) );
  XOR2_X1 u1_U484 (.Z( u1_FP_8 ) , .B( u1_L14_8 ) , .A( u1_out15_8 ) );
  XOR2_X1 u1_U489 (.Z( u1_FP_3 ) , .B( u1_L14_3 ) , .A( u1_out15_3 ) );
  XOR2_X1 u1_U49 (.B( u1_L0_26 ) , .Z( u1_N57 ) , .A( u1_out1_26 ) );
  XOR2_X1 u1_U497 (.Z( u1_FP_26 ) , .B( u1_L14_26 ) , .A( u1_out15_26 ) );
  XOR2_X1 u1_U498 (.Z( u1_FP_25 ) , .B( u1_L14_25 ) , .A( u1_out15_25 ) );
  XOR2_X1 u1_U50 (.B( u1_L0_25 ) , .Z( u1_N56 ) , .A( u1_out1_25 ) );
  XOR2_X1 u1_U503 (.Z( u1_FP_20 ) , .B( u1_L14_20 ) , .A( u1_out15_20 ) );
  XOR2_X1 u1_U504 (.Z( u1_FP_1 ) , .B( u1_L14_1 ) , .A( u1_out15_1 ) );
  XOR2_X1 u1_U51 (.B( u1_L0_24 ) , .Z( u1_N55 ) , .A( u1_out1_24 ) );
  XOR2_X1 u1_U510 (.Z( u1_FP_14 ) , .B( u1_L14_14 ) , .A( u1_out15_14 ) );
  XOR2_X1 u1_U514 (.Z( u1_FP_10 ) , .B( u1_L14_10 ) , .A( u1_out15_10 ) );
  XOR2_X1 u1_U52 (.B( u1_L0_23 ) , .Z( u1_N54 ) , .A( u1_out1_23 ) );
  XOR2_X1 u1_U53 (.B( u1_L0_22 ) , .Z( u1_N53 ) , .A( u1_out1_22 ) );
  XOR2_X1 u1_U54 (.B( u1_L0_21 ) , .Z( u1_N52 ) , .A( u1_out1_21 ) );
  XOR2_X1 u1_U55 (.B( u1_L0_20 ) , .Z( u1_N51 ) , .A( u1_out1_20 ) );
  XOR2_X1 u1_U59 (.B( u1_L0_17 ) , .Z( u1_N48 ) , .A( u1_out1_17 ) );
  XOR2_X1 u1_U6 (.B( u1_L2_1 ) , .Z( u1_N96 ) , .A( u1_out3_1 ) );
  XOR2_X1 u1_U60 (.B( u1_L13_32 ) , .Z( u1_N479 ) , .A( u1_out14_32 ) );
  XOR2_X1 u1_U62 (.B( u1_L13_30 ) , .Z( u1_N477 ) , .A( u1_out14_30 ) );
  XOR2_X1 u1_U63 (.B( u1_L13_29 ) , .Z( u1_N476 ) , .A( u1_out14_29 ) );
  XOR2_X1 u1_U65 (.B( u1_L13_27 ) , .Z( u1_N474 ) , .A( u1_out14_27 ) );
  XOR2_X1 u1_U68 (.B( u1_L13_24 ) , .Z( u1_N471 ) , .A( u1_out14_24 ) );
  XOR2_X1 u1_U70 (.B( u1_L0_16 ) , .Z( u1_N47 ) , .A( u1_out1_16 ) );
  XOR2_X1 u1_U71 (.B( u1_L13_22 ) , .Z( u1_N469 ) , .A( u1_out14_22 ) );
  XOR2_X1 u1_U72 (.B( u1_L13_21 ) , .Z( u1_N468 ) , .A( u1_out14_21 ) );
  XOR2_X1 u1_U74 (.B( u1_L13_19 ) , .Z( u1_N466 ) , .A( u1_out14_19 ) );
  XOR2_X1 u1_U77 (.B( u1_L13_16 ) , .Z( u1_N463 ) , .A( u1_out14_16 ) );
  XOR2_X1 u1_U78 (.B( u1_L13_15 ) , .Z( u1_N462 ) , .A( u1_out14_15 ) );
  XOR2_X1 u1_U81 (.B( u1_L0_15 ) , .Z( u1_N46 ) , .A( u1_out1_15 ) );
  XOR2_X1 u1_U82 (.B( u1_L13_12 ) , .Z( u1_N459 ) , .A( u1_out14_12 ) );
  XOR2_X1 u1_U83 (.B( u1_L13_11 ) , .Z( u1_N458 ) , .A( u1_out14_11 ) );
  XOR2_X1 u1_U87 (.B( u1_L13_7 ) , .Z( u1_N454 ) , .A( u1_out14_7 ) );
  XOR2_X1 u1_U88 (.B( u1_L13_6 ) , .Z( u1_N453 ) , .A( u1_out14_6 ) );
  XOR2_X1 u1_U89 (.B( u1_L13_5 ) , .Z( u1_N452 ) , .A( u1_out14_5 ) );
  XOR2_X1 u1_U90 (.B( u1_L13_4 ) , .Z( u1_N451 ) , .A( u1_out14_4 ) );
  XOR2_X1 u1_U92 (.B( u1_L0_14 ) , .Z( u1_N45 ) , .A( u1_out1_14 ) );
  XOR2_X1 u1_U95 (.B( u1_L12_32 ) , .Z( u1_N447 ) , .A( u1_out13_32 ) );
  XOR2_X1 u1_U99 (.B( u1_L12_28 ) , .Z( u1_N443 ) , .A( u1_out13_28 ) );
  XOR2_X1 u1_u0_U1 (.B( u1_K1_9 ) , .A( u1_desIn_r_47 ) , .Z( u1_u0_X_9 ) );
  XOR2_X1 u1_u0_U10 (.B( u1_K1_45 ) , .A( u1_desIn_r_41 ) , .Z( u1_u0_X_45 ) );
  XOR2_X1 u1_u0_U11 (.B( u1_K1_44 ) , .A( u1_desIn_r_33 ) , .Z( u1_u0_X_44 ) );
  XOR2_X1 u1_u0_U12 (.B( u1_K1_43 ) , .A( u1_desIn_r_25 ) , .Z( u1_u0_X_43 ) );
  XOR2_X1 u1_u0_U13 (.B( u1_K1_42 ) , .A( u1_desIn_r_33 ) , .Z( u1_u0_X_42 ) );
  XOR2_X1 u1_u0_U14 (.B( u1_K1_41 ) , .A( u1_desIn_r_25 ) , .Z( u1_u0_X_41 ) );
  XOR2_X1 u1_u0_U15 (.B( u1_K1_40 ) , .A( u1_desIn_r_17 ) , .Z( u1_u0_X_40 ) );
  XOR2_X1 u1_u0_U16 (.B( u1_K1_3 ) , .A( u1_desIn_r_15 ) , .Z( u1_u0_X_3 ) );
  XOR2_X1 u1_u0_U17 (.B( u1_K1_39 ) , .A( u1_desIn_r_9 ) , .Z( u1_u0_X_39 ) );
  XOR2_X1 u1_u0_U18 (.B( u1_K1_38 ) , .A( u1_desIn_r_1 ) , .Z( u1_u0_X_38 ) );
  XOR2_X1 u1_u0_U19 (.B( u1_K1_37 ) , .A( u1_desIn_r_59 ) , .Z( u1_u0_X_37 ) );
  XOR2_X1 u1_u0_U2 (.B( u1_K1_8 ) , .A( u1_desIn_r_39 ) , .Z( u1_u0_X_8 ) );
  XOR2_X1 u1_u0_U20 (.B( u1_K1_36 ) , .A( u1_desIn_r_1 ) , .Z( u1_u0_X_36 ) );
  XOR2_X1 u1_u0_U21 (.B( u1_K1_35 ) , .A( u1_desIn_r_59 ) , .Z( u1_u0_X_35 ) );
  XOR2_X1 u1_u0_U24 (.B( u1_K1_32 ) , .A( u1_desIn_r_35 ) , .Z( u1_u0_X_32 ) );
  XOR2_X1 u1_u0_U26 (.B( u1_K1_30 ) , .A( u1_desIn_r_35 ) , .Z( u1_u0_X_30 ) );
  XOR2_X1 u1_u0_U27 (.B( u1_K1_2 ) , .A( u1_desIn_r_7 ) , .Z( u1_u0_X_2 ) );
  XOR2_X1 u1_u0_U3 (.B( u1_K1_7 ) , .A( u1_desIn_r_31 ) , .Z( u1_u0_X_7 ) );
  XOR2_X1 u1_u0_U31 (.B( u1_K1_26 ) , .A( u1_desIn_r_3 ) , .Z( u1_u0_X_26 ) );
  XOR2_X1 u1_u0_U32 (.B( u1_K1_25 ) , .A( u1_desIn_r_61 ) , .Z( u1_u0_X_25 ) );
  XOR2_X1 u1_u0_U33 (.B( u1_K1_24 ) , .A( u1_desIn_r_3 ) , .Z( u1_u0_X_24 ) );
  XOR2_X1 u1_u0_U34 (.B( u1_K1_23 ) , .A( u1_desIn_r_61 ) , .Z( u1_u0_X_23 ) );
  XOR2_X1 u1_u0_U35 (.B( u1_K1_22 ) , .A( u1_desIn_r_53 ) , .Z( u1_u0_X_22 ) );
  XOR2_X1 u1_u0_U36 (.B( u1_K1_21 ) , .A( u1_desIn_r_45 ) , .Z( u1_u0_X_21 ) );
  XOR2_X1 u1_u0_U37 (.B( u1_K1_20 ) , .A( u1_desIn_r_37 ) , .Z( u1_u0_X_20 ) );
  XOR2_X1 u1_u0_U38 (.B( u1_K1_1 ) , .A( u1_desIn_r_57 ) , .Z( u1_u0_X_1 ) );
  XOR2_X1 u1_u0_U39 (.B( u1_K1_19 ) , .A( u1_desIn_r_29 ) , .Z( u1_u0_X_19 ) );
  XOR2_X1 u1_u0_U4 (.B( u1_K1_6 ) , .A( u1_desIn_r_39 ) , .Z( u1_u0_X_6 ) );
  XOR2_X1 u1_u0_U40 (.B( u1_K1_18 ) , .A( u1_desIn_r_37 ) , .Z( u1_u0_X_18 ) );
  XOR2_X1 u1_u0_U41 (.B( u1_K1_17 ) , .A( u1_desIn_r_29 ) , .Z( u1_u0_X_17 ) );
  XOR2_X1 u1_u0_U44 (.B( u1_K1_14 ) , .A( u1_desIn_r_5 ) , .Z( u1_u0_X_14 ) );
  XOR2_X1 u1_u0_U45 (.B( u1_K1_13 ) , .A( u1_desIn_r_63 ) , .Z( u1_u0_X_13 ) );
  XOR2_X1 u1_u0_U46 (.B( u1_K1_12 ) , .A( u1_desIn_r_5 ) , .Z( u1_u0_X_12 ) );
  XOR2_X1 u1_u0_U47 (.B( u1_K1_11 ) , .A( u1_desIn_r_63 ) , .Z( u1_u0_X_11 ) );
  XOR2_X1 u1_u0_U48 (.B( u1_K1_10 ) , .A( u1_desIn_r_55 ) , .Z( u1_u0_X_10 ) );
  XOR2_X1 u1_u0_U5 (.B( u1_K1_5 ) , .A( u1_desIn_r_31 ) , .Z( u1_u0_X_5 ) );
  XOR2_X1 u1_u0_U6 (.B( u1_K1_4 ) , .A( u1_desIn_r_23 ) , .Z( u1_u0_X_4 ) );
  XOR2_X1 u1_u0_U7 (.B( u1_K1_48 ) , .A( u1_desIn_r_7 ) , .Z( u1_u0_X_48 ) );
  XOR2_X1 u1_u0_U8 (.B( u1_K1_47 ) , .A( u1_desIn_r_57 ) , .Z( u1_u0_X_47 ) );
  XOR2_X1 u1_u0_U9 (.B( u1_K1_46 ) , .A( u1_desIn_r_49 ) , .Z( u1_u0_X_46 ) );
  NAND2_X1 u1_u0_u0_U10 (.ZN( u1_u0_u0_n113 ) , .A1( u1_u0_u0_n139 ) , .A2( u1_u0_u0_n149 ) );
  AND3_X1 u1_u0_u0_U11 (.A2( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n127 ) , .A3( u1_u0_u0_n130 ) , .A1( u1_u0_u0_n148 ) );
  AND2_X1 u1_u0_u0_U12 (.ZN( u1_u0_u0_n107 ) , .A1( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n140 ) );
  AND2_X1 u1_u0_u0_U13 (.A2( u1_u0_u0_n129 ) , .A1( u1_u0_u0_n130 ) , .ZN( u1_u0_u0_n151 ) );
  AND2_X1 u1_u0_u0_U14 (.A1( u1_u0_u0_n108 ) , .A2( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U15 (.A( u1_u0_u0_n143 ) , .ZN( u1_u0_u0_n173 ) );
  NOR2_X1 u1_u0_u0_U16 (.A2( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n147 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U17 (.ZN( u1_u0_u0_n172 ) , .A( u1_u0_u0_n88 ) );
  OAI222_X1 u1_u0_u0_U18 (.C1( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n125 ) , .B2( u1_u0_u0_n128 ) , .B1( u1_u0_u0_n144 ) , .A2( u1_u0_u0_n158 ) , .C2( u1_u0_u0_n161 ) , .ZN( u1_u0_u0_n88 ) );
  AOI21_X1 u1_u0_u0_U19 (.B1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n132 ) , .A( u1_u0_u0_n165 ) , .B2( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U20 (.A( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n165 ) );
  OAI22_X1 u1_u0_u0_U21 (.B1( u1_u0_u0_n125 ) , .ZN( u1_u0_u0_n126 ) , .A1( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n146 ) , .B2( u1_u0_u0_n147 ) );
  OAI22_X1 u1_u0_u0_U22 (.B1( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n147 ) , .A2( u1_u0_u0_n90 ) , .ZN( u1_u0_u0_n91 ) );
  AND3_X1 u1_u0_u0_U23 (.A3( u1_u0_u0_n121 ) , .A2( u1_u0_u0_n125 ) , .A1( u1_u0_u0_n148 ) , .ZN( u1_u0_u0_n90 ) );
  INV_X1 u1_u0_u0_U24 (.A( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n161 ) );
  AOI22_X1 u1_u0_u0_U25 (.B2( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n110 ) , .ZN( u1_u0_u0_n111 ) , .B1( u1_u0_u0_n118 ) , .A1( u1_u0_u0_n160 ) );
  INV_X1 u1_u0_u0_U26 (.A( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U27 (.B1( u1_u0_u0_n127 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n96 ) );
  AOI21_X1 u1_u0_u0_U28 (.ZN( u1_u0_u0_n104 ) , .B1( u1_u0_u0_n107 ) , .B2( u1_u0_u0_n141 ) , .A( u1_u0_u0_n144 ) );
  NAND2_X1 u1_u0_u0_U29 (.A1( u1_u0_u0_n100 ) , .A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n125 ) );
  INV_X1 u1_u0_u0_U3 (.A( u1_u0_u0_n113 ) , .ZN( u1_u0_u0_n166 ) );
  NAND2_X1 u1_u0_u0_U30 (.A2( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n131 ) , .A1( u1_u0_u0_n92 ) );
  NAND2_X1 u1_u0_u0_U31 (.A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n114 ) , .A1( u1_u0_u0_n92 ) );
  NOR2_X1 u1_u0_u0_U32 (.A1( u1_u0_u0_n120 ) , .ZN( u1_u0_u0_n143 ) , .A2( u1_u0_u0_n167 ) );
  OAI221_X1 u1_u0_u0_U33 (.C1( u1_u0_u0_n112 ) , .ZN( u1_u0_u0_n120 ) , .B1( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n141 ) , .C2( u1_u0_u0_n147 ) , .A( u1_u0_u0_n172 ) );
  AOI21_X1 u1_u0_u0_U34 (.ZN( u1_u0_u0_n116 ) , .B2( u1_u0_u0_n142 ) , .A( u1_u0_u0_n144 ) , .B1( u1_u0_u0_n166 ) );
  INV_X1 u1_u0_u0_U35 (.A( u1_u0_u0_n138 ) , .ZN( u1_u0_u0_n160 ) );
  NAND2_X1 u1_u0_u0_U36 (.A2( u1_u0_u0_n102 ) , .A1( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n149 ) );
  NAND2_X1 u1_u0_u0_U37 (.ZN( u1_u0_u0_n112 ) , .A2( u1_u0_u0_n92 ) , .A1( u1_u0_u0_n93 ) );
  OR3_X1 u1_u0_u0_U38 (.A3( u1_u0_u0_n152 ) , .A2( u1_u0_u0_n153 ) , .A1( u1_u0_u0_n154 ) , .ZN( u1_u0_u0_n155 ) );
  AOI21_X1 u1_u0_u0_U39 (.B2( u1_u0_u0_n150 ) , .B1( u1_u0_u0_n151 ) , .ZN( u1_u0_u0_n152 ) , .A( u1_u0_u0_n158 ) );
  NOR2_X1 u1_u0_u0_U4 (.A1( u1_u0_u0_n108 ) , .ZN( u1_u0_u0_n123 ) , .A2( u1_u0_u0_n158 ) );
  AOI21_X1 u1_u0_u0_U40 (.A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n145 ) , .B1( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n154 ) );
  AOI21_X1 u1_u0_u0_U41 (.A( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n148 ) , .B1( u1_u0_u0_n149 ) , .ZN( u1_u0_u0_n153 ) );
  INV_X1 u1_u0_u0_U42 (.ZN( u1_u0_u0_n171 ) , .A( u1_u0_u0_n99 ) );
  OAI211_X1 u1_u0_u0_U43 (.C2( u1_u0_u0_n140 ) , .C1( u1_u0_u0_n161 ) , .A( u1_u0_u0_n169 ) , .B( u1_u0_u0_n98 ) , .ZN( u1_u0_u0_n99 ) );
  AOI211_X1 u1_u0_u0_U44 (.C1( u1_u0_u0_n118 ) , .A( u1_u0_u0_n123 ) , .B( u1_u0_u0_n96 ) , .C2( u1_u0_u0_n97 ) , .ZN( u1_u0_u0_n98 ) );
  INV_X1 u1_u0_u0_U45 (.ZN( u1_u0_u0_n169 ) , .A( u1_u0_u0_n91 ) );
  NOR2_X1 u1_u0_u0_U46 (.A2( u1_u0_X_2 ) , .ZN( u1_u0_u0_n103 ) , .A1( u1_u0_u0_n164 ) );
  NOR2_X1 u1_u0_u0_U47 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n118 ) );
  NAND2_X1 u1_u0_u0_U48 (.A2( u1_u0_X_4 ) , .A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n144 ) );
  NOR2_X1 u1_u0_u0_U49 (.A2( u1_u0_X_5 ) , .ZN( u1_u0_u0_n136 ) , .A1( u1_u0_u0_n159 ) );
  AOI21_X1 u1_u0_u0_U5 (.B2( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n134 ) , .B1( u1_u0_u0_n151 ) , .A( u1_u0_u0_n158 ) );
  NAND2_X1 u1_u0_u0_U50 (.A1( u1_u0_X_5 ) , .ZN( u1_u0_u0_n138 ) , .A2( u1_u0_u0_n159 ) );
  AND2_X1 u1_u0_u0_U51 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n102 ) );
  AND2_X1 u1_u0_u0_U52 (.A1( u1_u0_X_6 ) , .A2( u1_u0_u0_n162 ) , .ZN( u1_u0_u0_n93 ) );
  INV_X1 u1_u0_u0_U53 (.A( u1_u0_X_4 ) , .ZN( u1_u0_u0_n159 ) );
  INV_X1 u1_u0_u0_U54 (.A( u1_u0_X_2 ) , .ZN( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U55 (.A( u1_u0_X_3 ) , .ZN( u1_u0_u0_n162 ) );
  INV_X1 u1_u0_u0_U56 (.A( u1_u0_u0_n126 ) , .ZN( u1_u0_u0_n168 ) );
  AOI211_X1 u1_u0_u0_U57 (.B( u1_u0_u0_n133 ) , .A( u1_u0_u0_n134 ) , .C2( u1_u0_u0_n135 ) , .C1( u1_u0_u0_n136 ) , .ZN( u1_u0_u0_n137 ) );
  OR4_X1 u1_u0_u0_U58 (.ZN( u1_out0_17 ) , .A4( u1_u0_u0_n122 ) , .A2( u1_u0_u0_n123 ) , .A1( u1_u0_u0_n124 ) , .A3( u1_u0_u0_n170 ) );
  AOI21_X1 u1_u0_u0_U59 (.B2( u1_u0_u0_n107 ) , .ZN( u1_u0_u0_n124 ) , .B1( u1_u0_u0_n128 ) , .A( u1_u0_u0_n161 ) );
  OAI21_X1 u1_u0_u0_U6 (.B1( u1_u0_u0_n150 ) , .B2( u1_u0_u0_n158 ) , .A( u1_u0_u0_n172 ) , .ZN( u1_u0_u0_n89 ) );
  INV_X1 u1_u0_u0_U60 (.A( u1_u0_u0_n111 ) , .ZN( u1_u0_u0_n170 ) );
  OR4_X1 u1_u0_u0_U61 (.ZN( u1_out0_31 ) , .A4( u1_u0_u0_n155 ) , .A2( u1_u0_u0_n156 ) , .A1( u1_u0_u0_n157 ) , .A3( u1_u0_u0_n173 ) );
  AOI21_X1 u1_u0_u0_U62 (.A( u1_u0_u0_n138 ) , .B2( u1_u0_u0_n139 ) , .B1( u1_u0_u0_n140 ) , .ZN( u1_u0_u0_n157 ) );
  AOI21_X1 u1_u0_u0_U63 (.B2( u1_u0_u0_n141 ) , .B1( u1_u0_u0_n142 ) , .ZN( u1_u0_u0_n156 ) , .A( u1_u0_u0_n161 ) );
  INV_X1 u1_u0_u0_U64 (.ZN( u1_u0_u0_n174 ) , .A( u1_u0_u0_n89 ) );
  AOI211_X1 u1_u0_u0_U65 (.B( u1_u0_u0_n104 ) , .A( u1_u0_u0_n105 ) , .ZN( u1_u0_u0_n106 ) , .C2( u1_u0_u0_n113 ) , .C1( u1_u0_u0_n160 ) );
  AOI211_X1 u1_u0_u0_U66 (.B( u1_u0_u0_n115 ) , .A( u1_u0_u0_n116 ) , .C2( u1_u0_u0_n117 ) , .C1( u1_u0_u0_n118 ) , .ZN( u1_u0_u0_n119 ) );
  NAND2_X1 u1_u0_u0_U67 (.A2( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n121 ) , .A1( u1_u0_u0_n93 ) );
  NAND2_X1 u1_u0_u0_U68 (.A1( u1_u0_u0_n101 ) , .A2( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n150 ) );
  NOR2_X1 u1_u0_u0_U69 (.A2( u1_u0_X_1 ) , .A1( u1_u0_X_2 ) , .ZN( u1_u0_u0_n92 ) );
  AOI21_X1 u1_u0_u0_U7 (.B1( u1_u0_u0_n114 ) , .ZN( u1_u0_u0_n115 ) , .B2( u1_u0_u0_n129 ) , .A( u1_u0_u0_n161 ) );
  NAND2_X1 u1_u0_u0_U70 (.A2( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n139 ) );
  NOR2_X1 u1_u0_u0_U71 (.A2( u1_u0_X_1 ) , .ZN( u1_u0_u0_n101 ) , .A1( u1_u0_u0_n163 ) );
  INV_X1 u1_u0_u0_U72 (.A( u1_u0_X_1 ) , .ZN( u1_u0_u0_n164 ) );
  NAND2_X1 u1_u0_u0_U73 (.A1( u1_u0_u0_n102 ) , .ZN( u1_u0_u0_n128 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U74 (.A1( u1_u0_u0_n100 ) , .ZN( u1_u0_u0_n129 ) , .A2( u1_u0_u0_n95 ) );
  NAND2_X1 u1_u0_u0_U75 (.ZN( u1_u0_u0_n148 ) , .A1( u1_u0_u0_n93 ) , .A2( u1_u0_u0_n95 ) );
  OAI221_X1 u1_u0_u0_U76 (.C1( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n122 ) , .B2( u1_u0_u0_n127 ) , .A( u1_u0_u0_n143 ) , .B1( u1_u0_u0_n144 ) , .C2( u1_u0_u0_n147 ) );
  NOR2_X1 u1_u0_u0_U77 (.A1( u1_u0_u0_n163 ) , .A2( u1_u0_u0_n164 ) , .ZN( u1_u0_u0_n95 ) );
  AOI21_X1 u1_u0_u0_U78 (.B1( u1_u0_u0_n132 ) , .ZN( u1_u0_u0_n133 ) , .A( u1_u0_u0_n144 ) , .B2( u1_u0_u0_n166 ) );
  OAI22_X1 u1_u0_u0_U79 (.ZN( u1_u0_u0_n105 ) , .A2( u1_u0_u0_n132 ) , .B1( u1_u0_u0_n146 ) , .A1( u1_u0_u0_n147 ) , .B2( u1_u0_u0_n161 ) );
  AND2_X1 u1_u0_u0_U8 (.A1( u1_u0_u0_n114 ) , .A2( u1_u0_u0_n121 ) , .ZN( u1_u0_u0_n146 ) );
  NAND2_X1 u1_u0_u0_U80 (.ZN( u1_u0_u0_n110 ) , .A2( u1_u0_u0_n132 ) , .A1( u1_u0_u0_n145 ) );
  INV_X1 u1_u0_u0_U81 (.A( u1_u0_u0_n119 ) , .ZN( u1_u0_u0_n167 ) );
  NAND2_X1 u1_u0_u0_U82 (.A2( u1_u0_u0_n103 ) , .ZN( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U83 (.A1( u1_u0_u0_n101 ) , .ZN( u1_u0_u0_n130 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U84 (.ZN( u1_u0_u0_n108 ) , .A1( u1_u0_u0_n92 ) , .A2( u1_u0_u0_n94 ) );
  NAND2_X1 u1_u0_u0_U85 (.ZN( u1_u0_u0_n142 ) , .A1( u1_u0_u0_n94 ) , .A2( u1_u0_u0_n95 ) );
  NOR2_X1 u1_u0_u0_U86 (.A2( u1_u0_X_6 ) , .ZN( u1_u0_u0_n100 ) , .A1( u1_u0_u0_n162 ) );
  NOR2_X1 u1_u0_u0_U87 (.A2( u1_u0_X_3 ) , .A1( u1_u0_X_6 ) , .ZN( u1_u0_u0_n94 ) );
  NAND3_X1 u1_u0_u0_U88 (.ZN( u1_out0_23 ) , .A3( u1_u0_u0_n137 ) , .A1( u1_u0_u0_n168 ) , .A2( u1_u0_u0_n171 ) );
  NAND3_X1 u1_u0_u0_U89 (.A3( u1_u0_u0_n127 ) , .A2( u1_u0_u0_n128 ) , .ZN( u1_u0_u0_n135 ) , .A1( u1_u0_u0_n150 ) );
  AND2_X1 u1_u0_u0_U9 (.A1( u1_u0_u0_n131 ) , .ZN( u1_u0_u0_n141 ) , .A2( u1_u0_u0_n150 ) );
  NAND3_X1 u1_u0_u0_U90 (.ZN( u1_u0_u0_n117 ) , .A3( u1_u0_u0_n132 ) , .A2( u1_u0_u0_n139 ) , .A1( u1_u0_u0_n148 ) );
  NAND3_X1 u1_u0_u0_U91 (.ZN( u1_u0_u0_n109 ) , .A2( u1_u0_u0_n114 ) , .A3( u1_u0_u0_n140 ) , .A1( u1_u0_u0_n149 ) );
  NAND3_X1 u1_u0_u0_U92 (.ZN( u1_out0_9 ) , .A3( u1_u0_u0_n106 ) , .A2( u1_u0_u0_n171 ) , .A1( u1_u0_u0_n174 ) );
  NAND3_X1 u1_u0_u0_U93 (.A2( u1_u0_u0_n128 ) , .A1( u1_u0_u0_n132 ) , .A3( u1_u0_u0_n146 ) , .ZN( u1_u0_u0_n97 ) );
  AOI21_X1 u1_u0_u1_U10 (.B2( u1_u0_u1_n155 ) , .B1( u1_u0_u1_n156 ) , .ZN( u1_u0_u1_n157 ) , .A( u1_u0_u1_n174 ) );
  NAND3_X1 u1_u0_u1_U100 (.ZN( u1_u0_u1_n113 ) , .A1( u1_u0_u1_n120 ) , .A3( u1_u0_u1_n133 ) , .A2( u1_u0_u1_n155 ) );
  NAND2_X1 u1_u0_u1_U11 (.ZN( u1_u0_u1_n140 ) , .A2( u1_u0_u1_n150 ) , .A1( u1_u0_u1_n155 ) );
  NAND2_X1 u1_u0_u1_U12 (.A1( u1_u0_u1_n131 ) , .ZN( u1_u0_u1_n147 ) , .A2( u1_u0_u1_n153 ) );
  AOI22_X1 u1_u0_u1_U13 (.B2( u1_u0_u1_n136 ) , .A2( u1_u0_u1_n137 ) , .ZN( u1_u0_u1_n143 ) , .A1( u1_u0_u1_n171 ) , .B1( u1_u0_u1_n173 ) );
  INV_X1 u1_u0_u1_U14 (.A( u1_u0_u1_n147 ) , .ZN( u1_u0_u1_n181 ) );
  INV_X1 u1_u0_u1_U15 (.A( u1_u0_u1_n139 ) , .ZN( u1_u0_u1_n174 ) );
  OR4_X1 u1_u0_u1_U16 (.A4( u1_u0_u1_n106 ) , .A3( u1_u0_u1_n107 ) , .ZN( u1_u0_u1_n108 ) , .A1( u1_u0_u1_n117 ) , .A2( u1_u0_u1_n184 ) );
  AOI21_X1 u1_u0_u1_U17 (.ZN( u1_u0_u1_n106 ) , .A( u1_u0_u1_n112 ) , .B1( u1_u0_u1_n154 ) , .B2( u1_u0_u1_n156 ) );
  AOI21_X1 u1_u0_u1_U18 (.ZN( u1_u0_u1_n107 ) , .B1( u1_u0_u1_n134 ) , .B2( u1_u0_u1_n149 ) , .A( u1_u0_u1_n174 ) );
  INV_X1 u1_u0_u1_U19 (.A( u1_u0_u1_n101 ) , .ZN( u1_u0_u1_n184 ) );
  INV_X1 u1_u0_u1_U20 (.A( u1_u0_u1_n112 ) , .ZN( u1_u0_u1_n171 ) );
  NAND2_X1 u1_u0_u1_U21 (.ZN( u1_u0_u1_n141 ) , .A1( u1_u0_u1_n153 ) , .A2( u1_u0_u1_n156 ) );
  AND2_X1 u1_u0_u1_U22 (.A1( u1_u0_u1_n123 ) , .ZN( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n161 ) );
  NAND2_X1 u1_u0_u1_U23 (.A2( u1_u0_u1_n115 ) , .A1( u1_u0_u1_n116 ) , .ZN( u1_u0_u1_n148 ) );
  NAND2_X1 u1_u0_u1_U24 (.A2( u1_u0_u1_n133 ) , .A1( u1_u0_u1_n135 ) , .ZN( u1_u0_u1_n159 ) );
  NAND2_X1 u1_u0_u1_U25 (.A2( u1_u0_u1_n115 ) , .A1( u1_u0_u1_n120 ) , .ZN( u1_u0_u1_n132 ) );
  INV_X1 u1_u0_u1_U26 (.A( u1_u0_u1_n154 ) , .ZN( u1_u0_u1_n178 ) );
  INV_X1 u1_u0_u1_U27 (.A( u1_u0_u1_n151 ) , .ZN( u1_u0_u1_n183 ) );
  AND2_X1 u1_u0_u1_U28 (.A1( u1_u0_u1_n129 ) , .A2( u1_u0_u1_n133 ) , .ZN( u1_u0_u1_n149 ) );
  INV_X1 u1_u0_u1_U29 (.A( u1_u0_u1_n131 ) , .ZN( u1_u0_u1_n180 ) );
  INV_X1 u1_u0_u1_U3 (.A( u1_u0_u1_n159 ) , .ZN( u1_u0_u1_n182 ) );
  AOI221_X1 u1_u0_u1_U30 (.B1( u1_u0_u1_n140 ) , .ZN( u1_u0_u1_n167 ) , .B2( u1_u0_u1_n172 ) , .C2( u1_u0_u1_n175 ) , .C1( u1_u0_u1_n178 ) , .A( u1_u0_u1_n188 ) );
  INV_X1 u1_u0_u1_U31 (.ZN( u1_u0_u1_n188 ) , .A( u1_u0_u1_n97 ) );
  AOI211_X1 u1_u0_u1_U32 (.A( u1_u0_u1_n118 ) , .C1( u1_u0_u1_n132 ) , .C2( u1_u0_u1_n139 ) , .B( u1_u0_u1_n96 ) , .ZN( u1_u0_u1_n97 ) );
  AOI21_X1 u1_u0_u1_U33 (.B2( u1_u0_u1_n121 ) , .B1( u1_u0_u1_n135 ) , .A( u1_u0_u1_n152 ) , .ZN( u1_u0_u1_n96 ) );
  OAI221_X1 u1_u0_u1_U34 (.A( u1_u0_u1_n119 ) , .C2( u1_u0_u1_n129 ) , .ZN( u1_u0_u1_n138 ) , .B2( u1_u0_u1_n152 ) , .C1( u1_u0_u1_n174 ) , .B1( u1_u0_u1_n187 ) );
  INV_X1 u1_u0_u1_U35 (.A( u1_u0_u1_n148 ) , .ZN( u1_u0_u1_n187 ) );
  AOI211_X1 u1_u0_u1_U36 (.B( u1_u0_u1_n117 ) , .A( u1_u0_u1_n118 ) , .ZN( u1_u0_u1_n119 ) , .C2( u1_u0_u1_n146 ) , .C1( u1_u0_u1_n159 ) );
  NOR2_X1 u1_u0_u1_U37 (.A1( u1_u0_u1_n168 ) , .A2( u1_u0_u1_n176 ) , .ZN( u1_u0_u1_n98 ) );
  AOI211_X1 u1_u0_u1_U38 (.B( u1_u0_u1_n162 ) , .A( u1_u0_u1_n163 ) , .C2( u1_u0_u1_n164 ) , .ZN( u1_u0_u1_n165 ) , .C1( u1_u0_u1_n171 ) );
  AOI21_X1 u1_u0_u1_U39 (.A( u1_u0_u1_n160 ) , .B2( u1_u0_u1_n161 ) , .ZN( u1_u0_u1_n162 ) , .B1( u1_u0_u1_n182 ) );
  AOI221_X1 u1_u0_u1_U4 (.A( u1_u0_u1_n138 ) , .C2( u1_u0_u1_n139 ) , .C1( u1_u0_u1_n140 ) , .B2( u1_u0_u1_n141 ) , .ZN( u1_u0_u1_n142 ) , .B1( u1_u0_u1_n175 ) );
  OR2_X1 u1_u0_u1_U40 (.A2( u1_u0_u1_n157 ) , .A1( u1_u0_u1_n158 ) , .ZN( u1_u0_u1_n163 ) );
  OAI21_X1 u1_u0_u1_U41 (.B2( u1_u0_u1_n123 ) , .ZN( u1_u0_u1_n145 ) , .B1( u1_u0_u1_n160 ) , .A( u1_u0_u1_n185 ) );
  INV_X1 u1_u0_u1_U42 (.A( u1_u0_u1_n122 ) , .ZN( u1_u0_u1_n185 ) );
  AOI21_X1 u1_u0_u1_U43 (.B2( u1_u0_u1_n120 ) , .B1( u1_u0_u1_n121 ) , .ZN( u1_u0_u1_n122 ) , .A( u1_u0_u1_n128 ) );
  NAND2_X1 u1_u0_u1_U44 (.A1( u1_u0_u1_n128 ) , .ZN( u1_u0_u1_n146 ) , .A2( u1_u0_u1_n160 ) );
  NAND2_X1 u1_u0_u1_U45 (.A2( u1_u0_u1_n112 ) , .ZN( u1_u0_u1_n139 ) , .A1( u1_u0_u1_n152 ) );
  NAND2_X1 u1_u0_u1_U46 (.A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n156 ) , .A2( u1_u0_u1_n99 ) );
  NOR2_X1 u1_u0_u1_U47 (.ZN( u1_u0_u1_n117 ) , .A1( u1_u0_u1_n121 ) , .A2( u1_u0_u1_n160 ) );
  AOI21_X1 u1_u0_u1_U48 (.A( u1_u0_u1_n128 ) , .B2( u1_u0_u1_n129 ) , .ZN( u1_u0_u1_n130 ) , .B1( u1_u0_u1_n150 ) );
  NAND2_X1 u1_u0_u1_U49 (.ZN( u1_u0_u1_n112 ) , .A1( u1_u0_u1_n169 ) , .A2( u1_u0_u1_n170 ) );
  AOI211_X1 u1_u0_u1_U5 (.ZN( u1_u0_u1_n124 ) , .A( u1_u0_u1_n138 ) , .C2( u1_u0_u1_n139 ) , .B( u1_u0_u1_n145 ) , .C1( u1_u0_u1_n147 ) );
  NAND2_X1 u1_u0_u1_U50 (.ZN( u1_u0_u1_n129 ) , .A2( u1_u0_u1_n95 ) , .A1( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U51 (.A1( u1_u0_u1_n102 ) , .ZN( u1_u0_u1_n154 ) , .A2( u1_u0_u1_n99 ) );
  NAND2_X1 u1_u0_u1_U52 (.A2( u1_u0_u1_n100 ) , .ZN( u1_u0_u1_n135 ) , .A1( u1_u0_u1_n99 ) );
  AOI21_X1 u1_u0_u1_U53 (.A( u1_u0_u1_n152 ) , .B2( u1_u0_u1_n153 ) , .B1( u1_u0_u1_n154 ) , .ZN( u1_u0_u1_n158 ) );
  INV_X1 u1_u0_u1_U54 (.A( u1_u0_u1_n160 ) , .ZN( u1_u0_u1_n175 ) );
  NAND2_X1 u1_u0_u1_U55 (.A1( u1_u0_u1_n100 ) , .ZN( u1_u0_u1_n116 ) , .A2( u1_u0_u1_n95 ) );
  NAND2_X1 u1_u0_u1_U56 (.A1( u1_u0_u1_n102 ) , .ZN( u1_u0_u1_n131 ) , .A2( u1_u0_u1_n95 ) );
  NAND2_X1 u1_u0_u1_U57 (.A2( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n121 ) , .A1( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U58 (.A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n153 ) , .A2( u1_u0_u1_n98 ) );
  NAND2_X1 u1_u0_u1_U59 (.A2( u1_u0_u1_n104 ) , .A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n133 ) );
  AOI22_X1 u1_u0_u1_U6 (.B2( u1_u0_u1_n113 ) , .A2( u1_u0_u1_n114 ) , .ZN( u1_u0_u1_n125 ) , .A1( u1_u0_u1_n171 ) , .B1( u1_u0_u1_n173 ) );
  NAND2_X1 u1_u0_u1_U60 (.ZN( u1_u0_u1_n150 ) , .A2( u1_u0_u1_n98 ) , .A1( u1_u0_u1_n99 ) );
  NAND2_X1 u1_u0_u1_U61 (.A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n155 ) , .A2( u1_u0_u1_n95 ) );
  OAI21_X1 u1_u0_u1_U62 (.ZN( u1_u0_u1_n109 ) , .B1( u1_u0_u1_n129 ) , .B2( u1_u0_u1_n160 ) , .A( u1_u0_u1_n167 ) );
  NAND2_X1 u1_u0_u1_U63 (.A2( u1_u0_u1_n100 ) , .A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n120 ) );
  NAND2_X1 u1_u0_u1_U64 (.A1( u1_u0_u1_n102 ) , .A2( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n115 ) );
  NAND2_X1 u1_u0_u1_U65 (.A2( u1_u0_u1_n100 ) , .A1( u1_u0_u1_n104 ) , .ZN( u1_u0_u1_n151 ) );
  NAND2_X1 u1_u0_u1_U66 (.A2( u1_u0_u1_n103 ) , .A1( u1_u0_u1_n105 ) , .ZN( u1_u0_u1_n161 ) );
  INV_X1 u1_u0_u1_U67 (.A( u1_u0_u1_n152 ) , .ZN( u1_u0_u1_n173 ) );
  INV_X1 u1_u0_u1_U68 (.A( u1_u0_u1_n128 ) , .ZN( u1_u0_u1_n172 ) );
  NAND2_X1 u1_u0_u1_U69 (.A2( u1_u0_u1_n102 ) , .A1( u1_u0_u1_n103 ) , .ZN( u1_u0_u1_n123 ) );
  NAND2_X1 u1_u0_u1_U7 (.ZN( u1_u0_u1_n114 ) , .A1( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n156 ) );
  NOR2_X1 u1_u0_u1_U70 (.A2( u1_u0_X_7 ) , .A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n95 ) );
  NOR2_X1 u1_u0_u1_U71 (.A1( u1_u0_X_12 ) , .A2( u1_u0_X_9 ) , .ZN( u1_u0_u1_n100 ) );
  NOR2_X1 u1_u0_u1_U72 (.A2( u1_u0_X_8 ) , .A1( u1_u0_u1_n177 ) , .ZN( u1_u0_u1_n99 ) );
  NOR2_X1 u1_u0_u1_U73 (.A2( u1_u0_X_12 ) , .ZN( u1_u0_u1_n102 ) , .A1( u1_u0_u1_n176 ) );
  NOR2_X1 u1_u0_u1_U74 (.A2( u1_u0_X_9 ) , .ZN( u1_u0_u1_n105 ) , .A1( u1_u0_u1_n168 ) );
  NAND2_X1 u1_u0_u1_U75 (.A1( u1_u0_X_10 ) , .ZN( u1_u0_u1_n160 ) , .A2( u1_u0_u1_n169 ) );
  NAND2_X1 u1_u0_u1_U76 (.A2( u1_u0_X_10 ) , .A1( u1_u0_X_11 ) , .ZN( u1_u0_u1_n152 ) );
  NAND2_X1 u1_u0_u1_U77 (.A1( u1_u0_X_11 ) , .ZN( u1_u0_u1_n128 ) , .A2( u1_u0_u1_n170 ) );
  AND2_X1 u1_u0_u1_U78 (.A2( u1_u0_X_7 ) , .A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n104 ) );
  AND2_X1 u1_u0_u1_U79 (.A1( u1_u0_X_8 ) , .ZN( u1_u0_u1_n103 ) , .A2( u1_u0_u1_n177 ) );
  NOR2_X1 u1_u0_u1_U8 (.A1( u1_u0_u1_n112 ) , .A2( u1_u0_u1_n116 ) , .ZN( u1_u0_u1_n118 ) );
  INV_X1 u1_u0_u1_U80 (.A( u1_u0_X_10 ) , .ZN( u1_u0_u1_n170 ) );
  INV_X1 u1_u0_u1_U81 (.A( u1_u0_X_9 ) , .ZN( u1_u0_u1_n176 ) );
  INV_X1 u1_u0_u1_U82 (.A( u1_u0_X_11 ) , .ZN( u1_u0_u1_n169 ) );
  INV_X1 u1_u0_u1_U83 (.A( u1_u0_X_12 ) , .ZN( u1_u0_u1_n168 ) );
  INV_X1 u1_u0_u1_U84 (.A( u1_u0_X_7 ) , .ZN( u1_u0_u1_n177 ) );
  NAND4_X1 u1_u0_u1_U85 (.ZN( u1_out0_28 ) , .A4( u1_u0_u1_n124 ) , .A3( u1_u0_u1_n125 ) , .A2( u1_u0_u1_n126 ) , .A1( u1_u0_u1_n127 ) );
  OAI21_X1 u1_u0_u1_U86 (.ZN( u1_u0_u1_n127 ) , .B2( u1_u0_u1_n139 ) , .B1( u1_u0_u1_n175 ) , .A( u1_u0_u1_n183 ) );
  OAI21_X1 u1_u0_u1_U87 (.ZN( u1_u0_u1_n126 ) , .B2( u1_u0_u1_n140 ) , .A( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n178 ) );
  NAND4_X1 u1_u0_u1_U88 (.ZN( u1_out0_18 ) , .A4( u1_u0_u1_n165 ) , .A3( u1_u0_u1_n166 ) , .A1( u1_u0_u1_n167 ) , .A2( u1_u0_u1_n186 ) );
  AOI22_X1 u1_u0_u1_U89 (.B2( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n147 ) , .A2( u1_u0_u1_n148 ) , .ZN( u1_u0_u1_n166 ) , .A1( u1_u0_u1_n172 ) );
  OAI21_X1 u1_u0_u1_U9 (.ZN( u1_u0_u1_n101 ) , .B1( u1_u0_u1_n141 ) , .A( u1_u0_u1_n146 ) , .B2( u1_u0_u1_n183 ) );
  INV_X1 u1_u0_u1_U90 (.A( u1_u0_u1_n145 ) , .ZN( u1_u0_u1_n186 ) );
  NAND4_X1 u1_u0_u1_U91 (.ZN( u1_out0_2 ) , .A4( u1_u0_u1_n142 ) , .A3( u1_u0_u1_n143 ) , .A2( u1_u0_u1_n144 ) , .A1( u1_u0_u1_n179 ) );
  OAI21_X1 u1_u0_u1_U92 (.B2( u1_u0_u1_n132 ) , .ZN( u1_u0_u1_n144 ) , .A( u1_u0_u1_n146 ) , .B1( u1_u0_u1_n180 ) );
  INV_X1 u1_u0_u1_U93 (.A( u1_u0_u1_n130 ) , .ZN( u1_u0_u1_n179 ) );
  OR4_X1 u1_u0_u1_U94 (.ZN( u1_out0_13 ) , .A4( u1_u0_u1_n108 ) , .A3( u1_u0_u1_n109 ) , .A2( u1_u0_u1_n110 ) , .A1( u1_u0_u1_n111 ) );
  AOI21_X1 u1_u0_u1_U95 (.ZN( u1_u0_u1_n111 ) , .A( u1_u0_u1_n128 ) , .B2( u1_u0_u1_n131 ) , .B1( u1_u0_u1_n135 ) );
  AOI21_X1 u1_u0_u1_U96 (.ZN( u1_u0_u1_n110 ) , .A( u1_u0_u1_n116 ) , .B1( u1_u0_u1_n152 ) , .B2( u1_u0_u1_n160 ) );
  NAND3_X1 u1_u0_u1_U97 (.A3( u1_u0_u1_n149 ) , .A2( u1_u0_u1_n150 ) , .A1( u1_u0_u1_n151 ) , .ZN( u1_u0_u1_n164 ) );
  NAND3_X1 u1_u0_u1_U98 (.A3( u1_u0_u1_n134 ) , .A2( u1_u0_u1_n135 ) , .ZN( u1_u0_u1_n136 ) , .A1( u1_u0_u1_n151 ) );
  NAND3_X1 u1_u0_u1_U99 (.A1( u1_u0_u1_n133 ) , .ZN( u1_u0_u1_n137 ) , .A2( u1_u0_u1_n154 ) , .A3( u1_u0_u1_n181 ) );
  OAI22_X1 u1_u0_u3_U10 (.B1( u1_u0_u3_n113 ) , .A2( u1_u0_u3_n135 ) , .A1( u1_u0_u3_n150 ) , .B2( u1_u0_u3_n164 ) , .ZN( u1_u0_u3_n98 ) );
  OAI211_X1 u1_u0_u3_U11 (.B( u1_u0_u3_n106 ) , .ZN( u1_u0_u3_n119 ) , .C2( u1_u0_u3_n128 ) , .C1( u1_u0_u3_n167 ) , .A( u1_u0_u3_n181 ) );
  AOI221_X1 u1_u0_u3_U12 (.C1( u1_u0_u3_n105 ) , .ZN( u1_u0_u3_n106 ) , .A( u1_u0_u3_n131 ) , .B2( u1_u0_u3_n132 ) , .C2( u1_u0_u3_n133 ) , .B1( u1_u0_u3_n169 ) );
  INV_X1 u1_u0_u3_U13 (.ZN( u1_u0_u3_n181 ) , .A( u1_u0_u3_n98 ) );
  NAND2_X1 u1_u0_u3_U14 (.ZN( u1_u0_u3_n105 ) , .A2( u1_u0_u3_n130 ) , .A1( u1_u0_u3_n155 ) );
  AOI22_X1 u1_u0_u3_U15 (.B1( u1_u0_u3_n115 ) , .A2( u1_u0_u3_n116 ) , .ZN( u1_u0_u3_n123 ) , .B2( u1_u0_u3_n133 ) , .A1( u1_u0_u3_n169 ) );
  NAND2_X1 u1_u0_u3_U16 (.ZN( u1_u0_u3_n116 ) , .A2( u1_u0_u3_n151 ) , .A1( u1_u0_u3_n182 ) );
  NOR2_X1 u1_u0_u3_U17 (.ZN( u1_u0_u3_n126 ) , .A2( u1_u0_u3_n150 ) , .A1( u1_u0_u3_n164 ) );
  AOI21_X1 u1_u0_u3_U18 (.ZN( u1_u0_u3_n112 ) , .B2( u1_u0_u3_n146 ) , .B1( u1_u0_u3_n155 ) , .A( u1_u0_u3_n167 ) );
  NAND2_X1 u1_u0_u3_U19 (.A1( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n142 ) , .A2( u1_u0_u3_n164 ) );
  NAND2_X1 u1_u0_u3_U20 (.ZN( u1_u0_u3_n132 ) , .A2( u1_u0_u3_n152 ) , .A1( u1_u0_u3_n156 ) );
  INV_X1 u1_u0_u3_U21 (.A( u1_u0_u3_n133 ) , .ZN( u1_u0_u3_n165 ) );
  AND2_X1 u1_u0_u3_U22 (.A2( u1_u0_u3_n113 ) , .A1( u1_u0_u3_n114 ) , .ZN( u1_u0_u3_n151 ) );
  INV_X1 u1_u0_u3_U23 (.A( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n170 ) );
  NAND2_X1 u1_u0_u3_U24 (.A1( u1_u0_u3_n107 ) , .A2( u1_u0_u3_n108 ) , .ZN( u1_u0_u3_n140 ) );
  NAND2_X1 u1_u0_u3_U25 (.ZN( u1_u0_u3_n117 ) , .A1( u1_u0_u3_n124 ) , .A2( u1_u0_u3_n148 ) );
  NAND2_X1 u1_u0_u3_U26 (.ZN( u1_u0_u3_n143 ) , .A1( u1_u0_u3_n165 ) , .A2( u1_u0_u3_n167 ) );
  INV_X1 u1_u0_u3_U27 (.A( u1_u0_u3_n130 ) , .ZN( u1_u0_u3_n177 ) );
  INV_X1 u1_u0_u3_U28 (.A( u1_u0_u3_n128 ) , .ZN( u1_u0_u3_n176 ) );
  INV_X1 u1_u0_u3_U29 (.A( u1_u0_u3_n155 ) , .ZN( u1_u0_u3_n174 ) );
  INV_X1 u1_u0_u3_U3 (.A( u1_u0_u3_n140 ) , .ZN( u1_u0_u3_n182 ) );
  INV_X1 u1_u0_u3_U30 (.A( u1_u0_u3_n139 ) , .ZN( u1_u0_u3_n185 ) );
  NOR2_X1 u1_u0_u3_U31 (.ZN( u1_u0_u3_n135 ) , .A2( u1_u0_u3_n141 ) , .A1( u1_u0_u3_n169 ) );
  OAI222_X1 u1_u0_u3_U32 (.C2( u1_u0_u3_n107 ) , .A2( u1_u0_u3_n108 ) , .B1( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n138 ) , .B2( u1_u0_u3_n146 ) , .C1( u1_u0_u3_n154 ) , .A1( u1_u0_u3_n164 ) );
  NOR4_X1 u1_u0_u3_U33 (.A4( u1_u0_u3_n157 ) , .A3( u1_u0_u3_n158 ) , .A2( u1_u0_u3_n159 ) , .A1( u1_u0_u3_n160 ) , .ZN( u1_u0_u3_n161 ) );
  AOI21_X1 u1_u0_u3_U34 (.B2( u1_u0_u3_n152 ) , .B1( u1_u0_u3_n153 ) , .ZN( u1_u0_u3_n158 ) , .A( u1_u0_u3_n164 ) );
  AOI21_X1 u1_u0_u3_U35 (.A( u1_u0_u3_n154 ) , .B2( u1_u0_u3_n155 ) , .B1( u1_u0_u3_n156 ) , .ZN( u1_u0_u3_n157 ) );
  AOI21_X1 u1_u0_u3_U36 (.A( u1_u0_u3_n149 ) , .B2( u1_u0_u3_n150 ) , .B1( u1_u0_u3_n151 ) , .ZN( u1_u0_u3_n159 ) );
  OAI211_X1 u1_u0_u3_U37 (.B( u1_u0_u3_n127 ) , .ZN( u1_u0_u3_n139 ) , .C1( u1_u0_u3_n150 ) , .C2( u1_u0_u3_n154 ) , .A( u1_u0_u3_n184 ) );
  INV_X1 u1_u0_u3_U38 (.A( u1_u0_u3_n125 ) , .ZN( u1_u0_u3_n184 ) );
  AOI221_X1 u1_u0_u3_U39 (.A( u1_u0_u3_n126 ) , .ZN( u1_u0_u3_n127 ) , .C2( u1_u0_u3_n132 ) , .C1( u1_u0_u3_n169 ) , .B2( u1_u0_u3_n170 ) , .B1( u1_u0_u3_n174 ) );
  INV_X1 u1_u0_u3_U4 (.A( u1_u0_u3_n129 ) , .ZN( u1_u0_u3_n183 ) );
  OAI22_X1 u1_u0_u3_U40 (.A1( u1_u0_u3_n124 ) , .ZN( u1_u0_u3_n125 ) , .B2( u1_u0_u3_n145 ) , .A2( u1_u0_u3_n165 ) , .B1( u1_u0_u3_n167 ) );
  AOI211_X1 u1_u0_u3_U41 (.ZN( u1_u0_u3_n109 ) , .A( u1_u0_u3_n119 ) , .C2( u1_u0_u3_n129 ) , .B( u1_u0_u3_n138 ) , .C1( u1_u0_u3_n141 ) );
  AOI211_X1 u1_u0_u3_U42 (.B( u1_u0_u3_n119 ) , .A( u1_u0_u3_n120 ) , .C2( u1_u0_u3_n121 ) , .ZN( u1_u0_u3_n122 ) , .C1( u1_u0_u3_n179 ) );
  INV_X1 u1_u0_u3_U43 (.A( u1_u0_u3_n156 ) , .ZN( u1_u0_u3_n179 ) );
  OAI22_X1 u1_u0_u3_U44 (.B1( u1_u0_u3_n118 ) , .ZN( u1_u0_u3_n120 ) , .A1( u1_u0_u3_n135 ) , .B2( u1_u0_u3_n154 ) , .A2( u1_u0_u3_n178 ) );
  AND3_X1 u1_u0_u3_U45 (.ZN( u1_u0_u3_n118 ) , .A2( u1_u0_u3_n124 ) , .A1( u1_u0_u3_n144 ) , .A3( u1_u0_u3_n152 ) );
  INV_X1 u1_u0_u3_U46 (.A( u1_u0_u3_n121 ) , .ZN( u1_u0_u3_n164 ) );
  NAND2_X1 u1_u0_u3_U47 (.ZN( u1_u0_u3_n133 ) , .A1( u1_u0_u3_n154 ) , .A2( u1_u0_u3_n164 ) );
  NOR2_X1 u1_u0_u3_U48 (.A1( u1_u0_u3_n113 ) , .ZN( u1_u0_u3_n131 ) , .A2( u1_u0_u3_n154 ) );
  NAND2_X1 u1_u0_u3_U49 (.A1( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n150 ) , .A2( u1_u0_u3_n99 ) );
  INV_X1 u1_u0_u3_U5 (.A( u1_u0_u3_n117 ) , .ZN( u1_u0_u3_n178 ) );
  NAND2_X1 u1_u0_u3_U50 (.A2( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n155 ) , .A1( u1_u0_u3_n97 ) );
  INV_X1 u1_u0_u3_U51 (.A( u1_u0_u3_n141 ) , .ZN( u1_u0_u3_n167 ) );
  AOI21_X1 u1_u0_u3_U52 (.B2( u1_u0_u3_n114 ) , .B1( u1_u0_u3_n146 ) , .A( u1_u0_u3_n154 ) , .ZN( u1_u0_u3_n94 ) );
  AOI21_X1 u1_u0_u3_U53 (.ZN( u1_u0_u3_n110 ) , .B2( u1_u0_u3_n142 ) , .B1( u1_u0_u3_n186 ) , .A( u1_u0_u3_n95 ) );
  INV_X1 u1_u0_u3_U54 (.A( u1_u0_u3_n145 ) , .ZN( u1_u0_u3_n186 ) );
  AOI21_X1 u1_u0_u3_U55 (.B1( u1_u0_u3_n124 ) , .A( u1_u0_u3_n149 ) , .B2( u1_u0_u3_n155 ) , .ZN( u1_u0_u3_n95 ) );
  INV_X1 u1_u0_u3_U56 (.A( u1_u0_u3_n149 ) , .ZN( u1_u0_u3_n169 ) );
  NAND2_X1 u1_u0_u3_U57 (.ZN( u1_u0_u3_n124 ) , .A1( u1_u0_u3_n96 ) , .A2( u1_u0_u3_n97 ) );
  NAND2_X1 u1_u0_u3_U58 (.A2( u1_u0_u3_n100 ) , .ZN( u1_u0_u3_n146 ) , .A1( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U59 (.A1( u1_u0_u3_n101 ) , .ZN( u1_u0_u3_n145 ) , .A2( u1_u0_u3_n99 ) );
  AOI221_X1 u1_u0_u3_U6 (.A( u1_u0_u3_n131 ) , .C2( u1_u0_u3_n132 ) , .C1( u1_u0_u3_n133 ) , .ZN( u1_u0_u3_n134 ) , .B1( u1_u0_u3_n143 ) , .B2( u1_u0_u3_n177 ) );
  NAND2_X1 u1_u0_u3_U60 (.A1( u1_u0_u3_n100 ) , .ZN( u1_u0_u3_n156 ) , .A2( u1_u0_u3_n99 ) );
  NAND2_X1 u1_u0_u3_U61 (.A2( u1_u0_u3_n101 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n148 ) );
  NAND2_X1 u1_u0_u3_U62 (.A1( u1_u0_u3_n100 ) , .A2( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n128 ) );
  NAND2_X1 u1_u0_u3_U63 (.A2( u1_u0_u3_n101 ) , .A1( u1_u0_u3_n102 ) , .ZN( u1_u0_u3_n152 ) );
  NAND2_X1 u1_u0_u3_U64 (.A2( u1_u0_u3_n101 ) , .ZN( u1_u0_u3_n114 ) , .A1( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U65 (.ZN( u1_u0_u3_n107 ) , .A1( u1_u0_u3_n97 ) , .A2( u1_u0_u3_n99 ) );
  NAND2_X1 u1_u0_u3_U66 (.A2( u1_u0_u3_n100 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n113 ) );
  NAND2_X1 u1_u0_u3_U67 (.A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n153 ) , .A2( u1_u0_u3_n97 ) );
  NAND2_X1 u1_u0_u3_U68 (.A2( u1_u0_u3_n103 ) , .A1( u1_u0_u3_n104 ) , .ZN( u1_u0_u3_n130 ) );
  NAND2_X1 u1_u0_u3_U69 (.A2( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n144 ) , .A1( u1_u0_u3_n96 ) );
  OAI22_X1 u1_u0_u3_U7 (.B2( u1_u0_u3_n147 ) , .A2( u1_u0_u3_n148 ) , .ZN( u1_u0_u3_n160 ) , .B1( u1_u0_u3_n165 ) , .A1( u1_u0_u3_n168 ) );
  NAND2_X1 u1_u0_u3_U70 (.A1( u1_u0_u3_n102 ) , .A2( u1_u0_u3_n103 ) , .ZN( u1_u0_u3_n108 ) );
  NOR2_X1 u1_u0_u3_U71 (.A2( u1_u0_X_19 ) , .A1( u1_u0_X_20 ) , .ZN( u1_u0_u3_n99 ) );
  NOR2_X1 u1_u0_u3_U72 (.A2( u1_u0_X_21 ) , .A1( u1_u0_X_24 ) , .ZN( u1_u0_u3_n103 ) );
  NOR2_X1 u1_u0_u3_U73 (.A2( u1_u0_X_24 ) , .A1( u1_u0_u3_n171 ) , .ZN( u1_u0_u3_n97 ) );
  NOR2_X1 u1_u0_u3_U74 (.A2( u1_u0_X_23 ) , .ZN( u1_u0_u3_n141 ) , .A1( u1_u0_u3_n166 ) );
  NOR2_X1 u1_u0_u3_U75 (.A2( u1_u0_X_19 ) , .A1( u1_u0_u3_n172 ) , .ZN( u1_u0_u3_n96 ) );
  NAND2_X1 u1_u0_u3_U76 (.A1( u1_u0_X_22 ) , .A2( u1_u0_X_23 ) , .ZN( u1_u0_u3_n154 ) );
  NAND2_X1 u1_u0_u3_U77 (.A1( u1_u0_X_23 ) , .ZN( u1_u0_u3_n149 ) , .A2( u1_u0_u3_n166 ) );
  NOR2_X1 u1_u0_u3_U78 (.A2( u1_u0_X_22 ) , .A1( u1_u0_X_23 ) , .ZN( u1_u0_u3_n121 ) );
  AND2_X1 u1_u0_u3_U79 (.A1( u1_u0_X_24 ) , .ZN( u1_u0_u3_n101 ) , .A2( u1_u0_u3_n171 ) );
  AND3_X1 u1_u0_u3_U8 (.A3( u1_u0_u3_n144 ) , .A2( u1_u0_u3_n145 ) , .A1( u1_u0_u3_n146 ) , .ZN( u1_u0_u3_n147 ) );
  AND2_X1 u1_u0_u3_U80 (.A1( u1_u0_X_19 ) , .ZN( u1_u0_u3_n102 ) , .A2( u1_u0_u3_n172 ) );
  AND2_X1 u1_u0_u3_U81 (.A1( u1_u0_X_21 ) , .A2( u1_u0_X_24 ) , .ZN( u1_u0_u3_n100 ) );
  AND2_X1 u1_u0_u3_U82 (.A2( u1_u0_X_19 ) , .A1( u1_u0_X_20 ) , .ZN( u1_u0_u3_n104 ) );
  INV_X1 u1_u0_u3_U83 (.A( u1_u0_X_22 ) , .ZN( u1_u0_u3_n166 ) );
  INV_X1 u1_u0_u3_U84 (.A( u1_u0_X_21 ) , .ZN( u1_u0_u3_n171 ) );
  INV_X1 u1_u0_u3_U85 (.A( u1_u0_X_20 ) , .ZN( u1_u0_u3_n172 ) );
  NAND4_X1 u1_u0_u3_U86 (.ZN( u1_out0_26 ) , .A4( u1_u0_u3_n109 ) , .A3( u1_u0_u3_n110 ) , .A2( u1_u0_u3_n111 ) , .A1( u1_u0_u3_n173 ) );
  INV_X1 u1_u0_u3_U87 (.ZN( u1_u0_u3_n173 ) , .A( u1_u0_u3_n94 ) );
  OAI21_X1 u1_u0_u3_U88 (.ZN( u1_u0_u3_n111 ) , .B2( u1_u0_u3_n117 ) , .A( u1_u0_u3_n133 ) , .B1( u1_u0_u3_n176 ) );
  NAND4_X1 u1_u0_u3_U89 (.ZN( u1_out0_20 ) , .A4( u1_u0_u3_n122 ) , .A3( u1_u0_u3_n123 ) , .A1( u1_u0_u3_n175 ) , .A2( u1_u0_u3_n180 ) );
  INV_X1 u1_u0_u3_U9 (.A( u1_u0_u3_n143 ) , .ZN( u1_u0_u3_n168 ) );
  INV_X1 u1_u0_u3_U90 (.A( u1_u0_u3_n126 ) , .ZN( u1_u0_u3_n180 ) );
  INV_X1 u1_u0_u3_U91 (.A( u1_u0_u3_n112 ) , .ZN( u1_u0_u3_n175 ) );
  NAND4_X1 u1_u0_u3_U92 (.ZN( u1_out0_1 ) , .A4( u1_u0_u3_n161 ) , .A3( u1_u0_u3_n162 ) , .A2( u1_u0_u3_n163 ) , .A1( u1_u0_u3_n185 ) );
  NAND2_X1 u1_u0_u3_U93 (.ZN( u1_u0_u3_n163 ) , .A2( u1_u0_u3_n170 ) , .A1( u1_u0_u3_n176 ) );
  AOI22_X1 u1_u0_u3_U94 (.B2( u1_u0_u3_n140 ) , .B1( u1_u0_u3_n141 ) , .A2( u1_u0_u3_n142 ) , .ZN( u1_u0_u3_n162 ) , .A1( u1_u0_u3_n177 ) );
  OR4_X1 u1_u0_u3_U95 (.ZN( u1_out0_10 ) , .A4( u1_u0_u3_n136 ) , .A3( u1_u0_u3_n137 ) , .A1( u1_u0_u3_n138 ) , .A2( u1_u0_u3_n139 ) );
  OAI222_X1 u1_u0_u3_U96 (.C1( u1_u0_u3_n128 ) , .ZN( u1_u0_u3_n137 ) , .B1( u1_u0_u3_n148 ) , .A2( u1_u0_u3_n150 ) , .B2( u1_u0_u3_n154 ) , .C2( u1_u0_u3_n164 ) , .A1( u1_u0_u3_n167 ) );
  OAI221_X1 u1_u0_u3_U97 (.A( u1_u0_u3_n134 ) , .B2( u1_u0_u3_n135 ) , .ZN( u1_u0_u3_n136 ) , .C1( u1_u0_u3_n149 ) , .B1( u1_u0_u3_n151 ) , .C2( u1_u0_u3_n183 ) );
  NAND3_X1 u1_u0_u3_U98 (.A1( u1_u0_u3_n114 ) , .ZN( u1_u0_u3_n115 ) , .A2( u1_u0_u3_n145 ) , .A3( u1_u0_u3_n153 ) );
  NAND3_X1 u1_u0_u3_U99 (.ZN( u1_u0_u3_n129 ) , .A2( u1_u0_u3_n144 ) , .A1( u1_u0_u3_n153 ) , .A3( u1_u0_u3_n182 ) );
  AOI22_X1 u1_u0_u6_U10 (.A2( u1_u0_u6_n151 ) , .B2( u1_u0_u6_n161 ) , .A1( u1_u0_u6_n167 ) , .B1( u1_u0_u6_n170 ) , .ZN( u1_u0_u6_n89 ) );
  AOI21_X1 u1_u0_u6_U11 (.B1( u1_u0_u6_n107 ) , .B2( u1_u0_u6_n132 ) , .A( u1_u0_u6_n158 ) , .ZN( u1_u0_u6_n88 ) );
  AOI21_X1 u1_u0_u6_U12 (.B2( u1_u0_u6_n147 ) , .B1( u1_u0_u6_n148 ) , .ZN( u1_u0_u6_n149 ) , .A( u1_u0_u6_n158 ) );
  AOI21_X1 u1_u0_u6_U13 (.ZN( u1_u0_u6_n106 ) , .A( u1_u0_u6_n142 ) , .B2( u1_u0_u6_n159 ) , .B1( u1_u0_u6_n164 ) );
  INV_X1 u1_u0_u6_U14 (.A( u1_u0_u6_n155 ) , .ZN( u1_u0_u6_n161 ) );
  INV_X1 u1_u0_u6_U15 (.A( u1_u0_u6_n128 ) , .ZN( u1_u0_u6_n164 ) );
  NAND2_X1 u1_u0_u6_U16 (.ZN( u1_u0_u6_n110 ) , .A1( u1_u0_u6_n122 ) , .A2( u1_u0_u6_n129 ) );
  NAND2_X1 u1_u0_u6_U17 (.ZN( u1_u0_u6_n124 ) , .A2( u1_u0_u6_n146 ) , .A1( u1_u0_u6_n148 ) );
  INV_X1 u1_u0_u6_U18 (.A( u1_u0_u6_n132 ) , .ZN( u1_u0_u6_n171 ) );
  AND2_X1 u1_u0_u6_U19 (.A1( u1_u0_u6_n100 ) , .ZN( u1_u0_u6_n130 ) , .A2( u1_u0_u6_n147 ) );
  INV_X1 u1_u0_u6_U20 (.A( u1_u0_u6_n127 ) , .ZN( u1_u0_u6_n173 ) );
  INV_X1 u1_u0_u6_U21 (.A( u1_u0_u6_n121 ) , .ZN( u1_u0_u6_n167 ) );
  INV_X1 u1_u0_u6_U22 (.A( u1_u0_u6_n100 ) , .ZN( u1_u0_u6_n169 ) );
  INV_X1 u1_u0_u6_U23 (.A( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n170 ) );
  INV_X1 u1_u0_u6_U24 (.A( u1_u0_u6_n113 ) , .ZN( u1_u0_u6_n168 ) );
  AND2_X1 u1_u0_u6_U25 (.A1( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n119 ) , .ZN( u1_u0_u6_n133 ) );
  AND2_X1 u1_u0_u6_U26 (.A2( u1_u0_u6_n121 ) , .A1( u1_u0_u6_n122 ) , .ZN( u1_u0_u6_n131 ) );
  AND3_X1 u1_u0_u6_U27 (.ZN( u1_u0_u6_n120 ) , .A2( u1_u0_u6_n127 ) , .A1( u1_u0_u6_n132 ) , .A3( u1_u0_u6_n145 ) );
  INV_X1 u1_u0_u6_U28 (.A( u1_u0_u6_n146 ) , .ZN( u1_u0_u6_n163 ) );
  AOI222_X1 u1_u0_u6_U29 (.ZN( u1_u0_u6_n114 ) , .A1( u1_u0_u6_n118 ) , .A2( u1_u0_u6_n126 ) , .B2( u1_u0_u6_n151 ) , .C2( u1_u0_u6_n159 ) , .C1( u1_u0_u6_n168 ) , .B1( u1_u0_u6_n169 ) );
  INV_X1 u1_u0_u6_U3 (.A( u1_u0_u6_n110 ) , .ZN( u1_u0_u6_n166 ) );
  NOR2_X1 u1_u0_u6_U30 (.A1( u1_u0_u6_n162 ) , .A2( u1_u0_u6_n165 ) , .ZN( u1_u0_u6_n98 ) );
  AOI211_X1 u1_u0_u6_U31 (.B( u1_u0_u6_n134 ) , .A( u1_u0_u6_n135 ) , .C1( u1_u0_u6_n136 ) , .ZN( u1_u0_u6_n137 ) , .C2( u1_u0_u6_n151 ) );
  AOI21_X1 u1_u0_u6_U32 (.B2( u1_u0_u6_n132 ) , .B1( u1_u0_u6_n133 ) , .ZN( u1_u0_u6_n134 ) , .A( u1_u0_u6_n158 ) );
  NAND4_X1 u1_u0_u6_U33 (.A4( u1_u0_u6_n127 ) , .A3( u1_u0_u6_n128 ) , .A2( u1_u0_u6_n129 ) , .A1( u1_u0_u6_n130 ) , .ZN( u1_u0_u6_n136 ) );
  AOI21_X1 u1_u0_u6_U34 (.B1( u1_u0_u6_n131 ) , .ZN( u1_u0_u6_n135 ) , .A( u1_u0_u6_n144 ) , .B2( u1_u0_u6_n146 ) );
  NAND2_X1 u1_u0_u6_U35 (.A1( u1_u0_u6_n144 ) , .ZN( u1_u0_u6_n151 ) , .A2( u1_u0_u6_n158 ) );
  NAND2_X1 u1_u0_u6_U36 (.ZN( u1_u0_u6_n132 ) , .A1( u1_u0_u6_n91 ) , .A2( u1_u0_u6_n97 ) );
  AOI22_X1 u1_u0_u6_U37 (.B2( u1_u0_u6_n110 ) , .B1( u1_u0_u6_n111 ) , .A1( u1_u0_u6_n112 ) , .ZN( u1_u0_u6_n115 ) , .A2( u1_u0_u6_n161 ) );
  NAND4_X1 u1_u0_u6_U38 (.A3( u1_u0_u6_n109 ) , .ZN( u1_u0_u6_n112 ) , .A4( u1_u0_u6_n132 ) , .A2( u1_u0_u6_n147 ) , .A1( u1_u0_u6_n166 ) );
  NOR2_X1 u1_u0_u6_U39 (.ZN( u1_u0_u6_n109 ) , .A1( u1_u0_u6_n170 ) , .A2( u1_u0_u6_n173 ) );
  INV_X1 u1_u0_u6_U4 (.A( u1_u0_u6_n142 ) , .ZN( u1_u0_u6_n174 ) );
  NOR2_X1 u1_u0_u6_U40 (.A2( u1_u0_u6_n126 ) , .ZN( u1_u0_u6_n155 ) , .A1( u1_u0_u6_n160 ) );
  NAND2_X1 u1_u0_u6_U41 (.ZN( u1_u0_u6_n146 ) , .A2( u1_u0_u6_n94 ) , .A1( u1_u0_u6_n99 ) );
  AOI21_X1 u1_u0_u6_U42 (.A( u1_u0_u6_n144 ) , .B2( u1_u0_u6_n145 ) , .B1( u1_u0_u6_n146 ) , .ZN( u1_u0_u6_n150 ) );
  INV_X1 u1_u0_u6_U43 (.A( u1_u0_u6_n111 ) , .ZN( u1_u0_u6_n158 ) );
  NAND2_X1 u1_u0_u6_U44 (.ZN( u1_u0_u6_n127 ) , .A1( u1_u0_u6_n91 ) , .A2( u1_u0_u6_n92 ) );
  NAND2_X1 u1_u0_u6_U45 (.ZN( u1_u0_u6_n129 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n96 ) );
  INV_X1 u1_u0_u6_U46 (.A( u1_u0_u6_n144 ) , .ZN( u1_u0_u6_n159 ) );
  NAND2_X1 u1_u0_u6_U47 (.ZN( u1_u0_u6_n145 ) , .A2( u1_u0_u6_n97 ) , .A1( u1_u0_u6_n98 ) );
  NAND2_X1 u1_u0_u6_U48 (.ZN( u1_u0_u6_n148 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n94 ) );
  NAND2_X1 u1_u0_u6_U49 (.ZN( u1_u0_u6_n108 ) , .A2( u1_u0_u6_n139 ) , .A1( u1_u0_u6_n144 ) );
  NAND2_X1 u1_u0_u6_U5 (.A2( u1_u0_u6_n143 ) , .ZN( u1_u0_u6_n152 ) , .A1( u1_u0_u6_n166 ) );
  NAND2_X1 u1_u0_u6_U50 (.ZN( u1_u0_u6_n121 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n97 ) );
  NAND2_X1 u1_u0_u6_U51 (.ZN( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n95 ) );
  AND2_X1 u1_u0_u6_U52 (.ZN( u1_u0_u6_n118 ) , .A2( u1_u0_u6_n91 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U53 (.ZN( u1_u0_u6_n147 ) , .A2( u1_u0_u6_n98 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U54 (.ZN( u1_u0_u6_n128 ) , .A1( u1_u0_u6_n94 ) , .A2( u1_u0_u6_n96 ) );
  NAND2_X1 u1_u0_u6_U55 (.ZN( u1_u0_u6_n119 ) , .A2( u1_u0_u6_n95 ) , .A1( u1_u0_u6_n99 ) );
  NAND2_X1 u1_u0_u6_U56 (.ZN( u1_u0_u6_n123 ) , .A2( u1_u0_u6_n91 ) , .A1( u1_u0_u6_n96 ) );
  NAND2_X1 u1_u0_u6_U57 (.ZN( u1_u0_u6_n100 ) , .A2( u1_u0_u6_n92 ) , .A1( u1_u0_u6_n98 ) );
  NAND2_X1 u1_u0_u6_U58 (.ZN( u1_u0_u6_n122 ) , .A1( u1_u0_u6_n94 ) , .A2( u1_u0_u6_n97 ) );
  INV_X1 u1_u0_u6_U59 (.A( u1_u0_u6_n139 ) , .ZN( u1_u0_u6_n160 ) );
  AOI22_X1 u1_u0_u6_U6 (.B2( u1_u0_u6_n101 ) , .A1( u1_u0_u6_n102 ) , .ZN( u1_u0_u6_n103 ) , .B1( u1_u0_u6_n160 ) , .A2( u1_u0_u6_n161 ) );
  NAND2_X1 u1_u0_u6_U60 (.ZN( u1_u0_u6_n113 ) , .A1( u1_u0_u6_n96 ) , .A2( u1_u0_u6_n98 ) );
  NOR2_X1 u1_u0_u6_U61 (.A2( u1_u0_X_40 ) , .A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n126 ) );
  NOR2_X1 u1_u0_u6_U62 (.A2( u1_u0_X_39 ) , .A1( u1_u0_X_42 ) , .ZN( u1_u0_u6_n92 ) );
  NOR2_X1 u1_u0_u6_U63 (.A2( u1_u0_X_39 ) , .A1( u1_u0_u6_n156 ) , .ZN( u1_u0_u6_n97 ) );
  NOR2_X1 u1_u0_u6_U64 (.A2( u1_u0_X_38 ) , .A1( u1_u0_u6_n165 ) , .ZN( u1_u0_u6_n95 ) );
  NOR2_X1 u1_u0_u6_U65 (.A2( u1_u0_X_41 ) , .ZN( u1_u0_u6_n111 ) , .A1( u1_u0_u6_n157 ) );
  NOR2_X1 u1_u0_u6_U66 (.A2( u1_u0_X_37 ) , .A1( u1_u0_u6_n162 ) , .ZN( u1_u0_u6_n94 ) );
  NOR2_X1 u1_u0_u6_U67 (.A2( u1_u0_X_37 ) , .A1( u1_u0_X_38 ) , .ZN( u1_u0_u6_n91 ) );
  NAND2_X1 u1_u0_u6_U68 (.A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n144 ) , .A2( u1_u0_u6_n157 ) );
  NAND2_X1 u1_u0_u6_U69 (.A2( u1_u0_X_40 ) , .A1( u1_u0_X_41 ) , .ZN( u1_u0_u6_n139 ) );
  NOR2_X1 u1_u0_u6_U7 (.A1( u1_u0_u6_n118 ) , .ZN( u1_u0_u6_n143 ) , .A2( u1_u0_u6_n168 ) );
  AND2_X1 u1_u0_u6_U70 (.A1( u1_u0_X_39 ) , .A2( u1_u0_u6_n156 ) , .ZN( u1_u0_u6_n96 ) );
  AND2_X1 u1_u0_u6_U71 (.A1( u1_u0_X_39 ) , .A2( u1_u0_X_42 ) , .ZN( u1_u0_u6_n99 ) );
  INV_X1 u1_u0_u6_U72 (.A( u1_u0_X_40 ) , .ZN( u1_u0_u6_n157 ) );
  INV_X1 u1_u0_u6_U73 (.A( u1_u0_X_37 ) , .ZN( u1_u0_u6_n165 ) );
  INV_X1 u1_u0_u6_U74 (.A( u1_u0_X_38 ) , .ZN( u1_u0_u6_n162 ) );
  INV_X1 u1_u0_u6_U75 (.A( u1_u0_X_42 ) , .ZN( u1_u0_u6_n156 ) );
  NAND4_X1 u1_u0_u6_U76 (.ZN( u1_out0_32 ) , .A4( u1_u0_u6_n103 ) , .A3( u1_u0_u6_n104 ) , .A2( u1_u0_u6_n105 ) , .A1( u1_u0_u6_n106 ) );
  AOI22_X1 u1_u0_u6_U77 (.ZN( u1_u0_u6_n105 ) , .A2( u1_u0_u6_n108 ) , .A1( u1_u0_u6_n118 ) , .B2( u1_u0_u6_n126 ) , .B1( u1_u0_u6_n171 ) );
  AOI22_X1 u1_u0_u6_U78 (.ZN( u1_u0_u6_n104 ) , .A1( u1_u0_u6_n111 ) , .B1( u1_u0_u6_n124 ) , .B2( u1_u0_u6_n151 ) , .A2( u1_u0_u6_n93 ) );
  NAND4_X1 u1_u0_u6_U79 (.ZN( u1_out0_12 ) , .A4( u1_u0_u6_n114 ) , .A3( u1_u0_u6_n115 ) , .A2( u1_u0_u6_n116 ) , .A1( u1_u0_u6_n117 ) );
  OAI21_X1 u1_u0_u6_U8 (.A( u1_u0_u6_n159 ) , .B1( u1_u0_u6_n169 ) , .B2( u1_u0_u6_n173 ) , .ZN( u1_u0_u6_n90 ) );
  OAI22_X1 u1_u0_u6_U80 (.B2( u1_u0_u6_n111 ) , .ZN( u1_u0_u6_n116 ) , .B1( u1_u0_u6_n126 ) , .A2( u1_u0_u6_n164 ) , .A1( u1_u0_u6_n167 ) );
  OAI21_X1 u1_u0_u6_U81 (.A( u1_u0_u6_n108 ) , .ZN( u1_u0_u6_n117 ) , .B2( u1_u0_u6_n141 ) , .B1( u1_u0_u6_n163 ) );
  OAI211_X1 u1_u0_u6_U82 (.ZN( u1_out0_7 ) , .B( u1_u0_u6_n153 ) , .C2( u1_u0_u6_n154 ) , .C1( u1_u0_u6_n155 ) , .A( u1_u0_u6_n174 ) );
  NOR3_X1 u1_u0_u6_U83 (.A1( u1_u0_u6_n141 ) , .ZN( u1_u0_u6_n154 ) , .A3( u1_u0_u6_n164 ) , .A2( u1_u0_u6_n171 ) );
  AOI211_X1 u1_u0_u6_U84 (.B( u1_u0_u6_n149 ) , .A( u1_u0_u6_n150 ) , .C2( u1_u0_u6_n151 ) , .C1( u1_u0_u6_n152 ) , .ZN( u1_u0_u6_n153 ) );
  OAI211_X1 u1_u0_u6_U85 (.ZN( u1_out0_22 ) , .B( u1_u0_u6_n137 ) , .A( u1_u0_u6_n138 ) , .C2( u1_u0_u6_n139 ) , .C1( u1_u0_u6_n140 ) );
  AOI22_X1 u1_u0_u6_U86 (.B1( u1_u0_u6_n124 ) , .A2( u1_u0_u6_n125 ) , .A1( u1_u0_u6_n126 ) , .ZN( u1_u0_u6_n138 ) , .B2( u1_u0_u6_n161 ) );
  AND4_X1 u1_u0_u6_U87 (.A3( u1_u0_u6_n119 ) , .A1( u1_u0_u6_n120 ) , .A4( u1_u0_u6_n129 ) , .ZN( u1_u0_u6_n140 ) , .A2( u1_u0_u6_n143 ) );
  NAND3_X1 u1_u0_u6_U88 (.A2( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n125 ) , .A1( u1_u0_u6_n130 ) , .A3( u1_u0_u6_n131 ) );
  NAND3_X1 u1_u0_u6_U89 (.A3( u1_u0_u6_n133 ) , .ZN( u1_u0_u6_n141 ) , .A1( u1_u0_u6_n145 ) , .A2( u1_u0_u6_n148 ) );
  INV_X1 u1_u0_u6_U9 (.ZN( u1_u0_u6_n172 ) , .A( u1_u0_u6_n88 ) );
  NAND3_X1 u1_u0_u6_U90 (.ZN( u1_u0_u6_n101 ) , .A3( u1_u0_u6_n107 ) , .A2( u1_u0_u6_n121 ) , .A1( u1_u0_u6_n127 ) );
  NAND3_X1 u1_u0_u6_U91 (.ZN( u1_u0_u6_n102 ) , .A3( u1_u0_u6_n130 ) , .A2( u1_u0_u6_n145 ) , .A1( u1_u0_u6_n166 ) );
  NAND3_X1 u1_u0_u6_U92 (.A3( u1_u0_u6_n113 ) , .A1( u1_u0_u6_n119 ) , .A2( u1_u0_u6_n123 ) , .ZN( u1_u0_u6_n93 ) );
  NAND3_X1 u1_u0_u6_U93 (.ZN( u1_u0_u6_n142 ) , .A2( u1_u0_u6_n172 ) , .A3( u1_u0_u6_n89 ) , .A1( u1_u0_u6_n90 ) );
  OAI21_X1 u1_u0_u7_U10 (.A( u1_u0_u7_n161 ) , .B1( u1_u0_u7_n168 ) , .B2( u1_u0_u7_n173 ) , .ZN( u1_u0_u7_n91 ) );
  AOI211_X1 u1_u0_u7_U11 (.A( u1_u0_u7_n117 ) , .ZN( u1_u0_u7_n118 ) , .C2( u1_u0_u7_n126 ) , .C1( u1_u0_u7_n177 ) , .B( u1_u0_u7_n180 ) );
  OAI22_X1 u1_u0_u7_U12 (.B1( u1_u0_u7_n115 ) , .ZN( u1_u0_u7_n117 ) , .A2( u1_u0_u7_n133 ) , .A1( u1_u0_u7_n137 ) , .B2( u1_u0_u7_n162 ) );
  INV_X1 u1_u0_u7_U13 (.A( u1_u0_u7_n116 ) , .ZN( u1_u0_u7_n180 ) );
  NOR3_X1 u1_u0_u7_U14 (.ZN( u1_u0_u7_n115 ) , .A3( u1_u0_u7_n145 ) , .A2( u1_u0_u7_n168 ) , .A1( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U15 (.A( u1_u0_u7_n133 ) , .ZN( u1_u0_u7_n176 ) );
  NOR3_X1 u1_u0_u7_U16 (.A2( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n135 ) , .ZN( u1_u0_u7_n136 ) , .A3( u1_u0_u7_n171 ) );
  NOR2_X1 u1_u0_u7_U17 (.A1( u1_u0_u7_n130 ) , .A2( u1_u0_u7_n134 ) , .ZN( u1_u0_u7_n153 ) );
  AOI21_X1 u1_u0_u7_U18 (.ZN( u1_u0_u7_n104 ) , .B2( u1_u0_u7_n112 ) , .B1( u1_u0_u7_n127 ) , .A( u1_u0_u7_n164 ) );
  AOI21_X1 u1_u0_u7_U19 (.ZN( u1_u0_u7_n106 ) , .B1( u1_u0_u7_n133 ) , .B2( u1_u0_u7_n146 ) , .A( u1_u0_u7_n162 ) );
  AOI21_X1 u1_u0_u7_U20 (.A( u1_u0_u7_n101 ) , .ZN( u1_u0_u7_n107 ) , .B2( u1_u0_u7_n128 ) , .B1( u1_u0_u7_n175 ) );
  INV_X1 u1_u0_u7_U21 (.A( u1_u0_u7_n101 ) , .ZN( u1_u0_u7_n165 ) );
  NOR2_X1 u1_u0_u7_U22 (.ZN( u1_u0_u7_n111 ) , .A2( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U23 (.A( u1_u0_u7_n138 ) , .ZN( u1_u0_u7_n171 ) );
  INV_X1 u1_u0_u7_U24 (.A( u1_u0_u7_n131 ) , .ZN( u1_u0_u7_n177 ) );
  INV_X1 u1_u0_u7_U25 (.A( u1_u0_u7_n110 ) , .ZN( u1_u0_u7_n174 ) );
  NAND2_X1 u1_u0_u7_U26 (.A1( u1_u0_u7_n129 ) , .A2( u1_u0_u7_n132 ) , .ZN( u1_u0_u7_n149 ) );
  NAND2_X1 u1_u0_u7_U27 (.A1( u1_u0_u7_n113 ) , .A2( u1_u0_u7_n124 ) , .ZN( u1_u0_u7_n130 ) );
  INV_X1 u1_u0_u7_U28 (.A( u1_u0_u7_n112 ) , .ZN( u1_u0_u7_n173 ) );
  INV_X1 u1_u0_u7_U29 (.A( u1_u0_u7_n128 ) , .ZN( u1_u0_u7_n168 ) );
  OAI21_X1 u1_u0_u7_U3 (.ZN( u1_u0_u7_n159 ) , .A( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n171 ) , .B1( u1_u0_u7_n174 ) );
  INV_X1 u1_u0_u7_U30 (.A( u1_u0_u7_n148 ) , .ZN( u1_u0_u7_n169 ) );
  INV_X1 u1_u0_u7_U31 (.A( u1_u0_u7_n127 ) , .ZN( u1_u0_u7_n179 ) );
  INV_X1 u1_u0_u7_U32 (.A( u1_u0_u7_n153 ) , .ZN( u1_u0_u7_n172 ) );
  NOR2_X1 u1_u0_u7_U33 (.ZN( u1_u0_u7_n101 ) , .A2( u1_u0_u7_n150 ) , .A1( u1_u0_u7_n156 ) );
  AOI211_X1 u1_u0_u7_U34 (.B( u1_u0_u7_n139 ) , .A( u1_u0_u7_n140 ) , .C2( u1_u0_u7_n141 ) , .ZN( u1_u0_u7_n142 ) , .C1( u1_u0_u7_n156 ) );
  NAND4_X1 u1_u0_u7_U35 (.A3( u1_u0_u7_n127 ) , .A2( u1_u0_u7_n128 ) , .A1( u1_u0_u7_n129 ) , .ZN( u1_u0_u7_n141 ) , .A4( u1_u0_u7_n147 ) );
  AOI21_X1 u1_u0_u7_U36 (.A( u1_u0_u7_n137 ) , .B1( u1_u0_u7_n138 ) , .ZN( u1_u0_u7_n139 ) , .B2( u1_u0_u7_n146 ) );
  OAI22_X1 u1_u0_u7_U37 (.B1( u1_u0_u7_n136 ) , .ZN( u1_u0_u7_n140 ) , .A1( u1_u0_u7_n153 ) , .B2( u1_u0_u7_n162 ) , .A2( u1_u0_u7_n164 ) );
  INV_X1 u1_u0_u7_U38 (.A( u1_u0_u7_n125 ) , .ZN( u1_u0_u7_n161 ) );
  AOI21_X1 u1_u0_u7_U39 (.ZN( u1_u0_u7_n123 ) , .B1( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n177 ) , .A( u1_u0_u7_n97 ) );
  INV_X1 u1_u0_u7_U4 (.A( u1_u0_u7_n149 ) , .ZN( u1_u0_u7_n175 ) );
  AOI21_X1 u1_u0_u7_U40 (.B2( u1_u0_u7_n113 ) , .B1( u1_u0_u7_n124 ) , .A( u1_u0_u7_n125 ) , .ZN( u1_u0_u7_n97 ) );
  INV_X1 u1_u0_u7_U41 (.A( u1_u0_u7_n152 ) , .ZN( u1_u0_u7_n162 ) );
  AOI22_X1 u1_u0_u7_U42 (.A2( u1_u0_u7_n114 ) , .ZN( u1_u0_u7_n119 ) , .B1( u1_u0_u7_n130 ) , .A1( u1_u0_u7_n156 ) , .B2( u1_u0_u7_n165 ) );
  NAND2_X1 u1_u0_u7_U43 (.A2( u1_u0_u7_n112 ) , .ZN( u1_u0_u7_n114 ) , .A1( u1_u0_u7_n175 ) );
  NOR2_X1 u1_u0_u7_U44 (.ZN( u1_u0_u7_n137 ) , .A1( u1_u0_u7_n150 ) , .A2( u1_u0_u7_n161 ) );
  AND2_X1 u1_u0_u7_U45 (.ZN( u1_u0_u7_n145 ) , .A2( u1_u0_u7_n98 ) , .A1( u1_u0_u7_n99 ) );
  AOI21_X1 u1_u0_u7_U46 (.ZN( u1_u0_u7_n105 ) , .B2( u1_u0_u7_n110 ) , .A( u1_u0_u7_n125 ) , .B1( u1_u0_u7_n147 ) );
  NAND2_X1 u1_u0_u7_U47 (.ZN( u1_u0_u7_n146 ) , .A1( u1_u0_u7_n95 ) , .A2( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U48 (.A2( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n147 ) , .A1( u1_u0_u7_n93 ) );
  NAND2_X1 u1_u0_u7_U49 (.A1( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n127 ) , .A2( u1_u0_u7_n99 ) );
  INV_X1 u1_u0_u7_U5 (.A( u1_u0_u7_n154 ) , .ZN( u1_u0_u7_n178 ) );
  NAND2_X1 u1_u0_u7_U50 (.A2( u1_u0_u7_n102 ) , .A1( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n133 ) );
  OR2_X1 u1_u0_u7_U51 (.ZN( u1_u0_u7_n126 ) , .A2( u1_u0_u7_n152 ) , .A1( u1_u0_u7_n156 ) );
  NAND2_X1 u1_u0_u7_U52 (.ZN( u1_u0_u7_n112 ) , .A2( u1_u0_u7_n96 ) , .A1( u1_u0_u7_n99 ) );
  NAND2_X1 u1_u0_u7_U53 (.A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n128 ) , .A1( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U54 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n113 ) , .A2( u1_u0_u7_n93 ) );
  NAND2_X1 u1_u0_u7_U55 (.ZN( u1_u0_u7_n110 ) , .A1( u1_u0_u7_n95 ) , .A2( u1_u0_u7_n96 ) );
  INV_X1 u1_u0_u7_U56 (.A( u1_u0_u7_n150 ) , .ZN( u1_u0_u7_n164 ) );
  AND2_X1 u1_u0_u7_U57 (.ZN( u1_u0_u7_n134 ) , .A1( u1_u0_u7_n93 ) , .A2( u1_u0_u7_n98 ) );
  NAND2_X1 u1_u0_u7_U58 (.A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n124 ) , .A1( u1_u0_u7_n96 ) );
  NAND2_X1 u1_u0_u7_U59 (.A1( u1_u0_u7_n100 ) , .A2( u1_u0_u7_n102 ) , .ZN( u1_u0_u7_n129 ) );
  AOI211_X1 u1_u0_u7_U6 (.ZN( u1_u0_u7_n116 ) , .A( u1_u0_u7_n155 ) , .C1( u1_u0_u7_n161 ) , .C2( u1_u0_u7_n171 ) , .B( u1_u0_u7_n94 ) );
  NAND2_X1 u1_u0_u7_U60 (.A2( u1_u0_u7_n103 ) , .ZN( u1_u0_u7_n131 ) , .A1( u1_u0_u7_n95 ) );
  NAND2_X1 u1_u0_u7_U61 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n138 ) , .A2( u1_u0_u7_n99 ) );
  NAND2_X1 u1_u0_u7_U62 (.ZN( u1_u0_u7_n132 ) , .A1( u1_u0_u7_n93 ) , .A2( u1_u0_u7_n96 ) );
  NAND2_X1 u1_u0_u7_U63 (.A1( u1_u0_u7_n100 ) , .ZN( u1_u0_u7_n148 ) , .A2( u1_u0_u7_n95 ) );
  NOR2_X1 u1_u0_u7_U64 (.A2( u1_u0_X_47 ) , .ZN( u1_u0_u7_n150 ) , .A1( u1_u0_u7_n163 ) );
  NOR2_X1 u1_u0_u7_U65 (.A2( u1_u0_X_43 ) , .A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n103 ) );
  NOR2_X1 u1_u0_u7_U66 (.A2( u1_u0_X_48 ) , .A1( u1_u0_u7_n166 ) , .ZN( u1_u0_u7_n95 ) );
  NOR2_X1 u1_u0_u7_U67 (.A2( u1_u0_X_45 ) , .A1( u1_u0_X_48 ) , .ZN( u1_u0_u7_n99 ) );
  NOR2_X1 u1_u0_u7_U68 (.A2( u1_u0_X_44 ) , .A1( u1_u0_u7_n167 ) , .ZN( u1_u0_u7_n98 ) );
  NOR2_X1 u1_u0_u7_U69 (.A2( u1_u0_X_46 ) , .A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n152 ) );
  OAI222_X1 u1_u0_u7_U7 (.C2( u1_u0_u7_n101 ) , .B2( u1_u0_u7_n111 ) , .A1( u1_u0_u7_n113 ) , .C1( u1_u0_u7_n146 ) , .A2( u1_u0_u7_n162 ) , .B1( u1_u0_u7_n164 ) , .ZN( u1_u0_u7_n94 ) );
  NAND2_X1 u1_u0_u7_U70 (.A2( u1_u0_X_46 ) , .A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n125 ) );
  AND2_X1 u1_u0_u7_U71 (.A1( u1_u0_X_47 ) , .ZN( u1_u0_u7_n156 ) , .A2( u1_u0_u7_n163 ) );
  AND2_X1 u1_u0_u7_U72 (.A2( u1_u0_X_45 ) , .A1( u1_u0_X_48 ) , .ZN( u1_u0_u7_n102 ) );
  AND2_X1 u1_u0_u7_U73 (.A2( u1_u0_X_43 ) , .A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n96 ) );
  AND2_X1 u1_u0_u7_U74 (.A1( u1_u0_X_44 ) , .ZN( u1_u0_u7_n100 ) , .A2( u1_u0_u7_n167 ) );
  AND2_X1 u1_u0_u7_U75 (.A1( u1_u0_X_48 ) , .A2( u1_u0_u7_n166 ) , .ZN( u1_u0_u7_n93 ) );
  INV_X1 u1_u0_u7_U76 (.A( u1_u0_X_46 ) , .ZN( u1_u0_u7_n163 ) );
  INV_X1 u1_u0_u7_U77 (.A( u1_u0_X_45 ) , .ZN( u1_u0_u7_n166 ) );
  NAND4_X1 u1_u0_u7_U78 (.ZN( u1_out0_5 ) , .A4( u1_u0_u7_n108 ) , .A3( u1_u0_u7_n109 ) , .A1( u1_u0_u7_n116 ) , .A2( u1_u0_u7_n123 ) );
  AOI22_X1 u1_u0_u7_U79 (.ZN( u1_u0_u7_n109 ) , .A2( u1_u0_u7_n126 ) , .B2( u1_u0_u7_n145 ) , .B1( u1_u0_u7_n156 ) , .A1( u1_u0_u7_n171 ) );
  OAI221_X1 u1_u0_u7_U8 (.C1( u1_u0_u7_n101 ) , .C2( u1_u0_u7_n147 ) , .ZN( u1_u0_u7_n155 ) , .B2( u1_u0_u7_n162 ) , .A( u1_u0_u7_n91 ) , .B1( u1_u0_u7_n92 ) );
  NOR4_X1 u1_u0_u7_U80 (.A4( u1_u0_u7_n104 ) , .A3( u1_u0_u7_n105 ) , .A2( u1_u0_u7_n106 ) , .A1( u1_u0_u7_n107 ) , .ZN( u1_u0_u7_n108 ) );
  NAND4_X1 u1_u0_u7_U81 (.ZN( u1_out0_27 ) , .A4( u1_u0_u7_n118 ) , .A3( u1_u0_u7_n119 ) , .A2( u1_u0_u7_n120 ) , .A1( u1_u0_u7_n121 ) );
  OAI21_X1 u1_u0_u7_U82 (.ZN( u1_u0_u7_n121 ) , .B2( u1_u0_u7_n145 ) , .A( u1_u0_u7_n150 ) , .B1( u1_u0_u7_n174 ) );
  OAI21_X1 u1_u0_u7_U83 (.ZN( u1_u0_u7_n120 ) , .A( u1_u0_u7_n161 ) , .B2( u1_u0_u7_n170 ) , .B1( u1_u0_u7_n179 ) );
  NAND4_X1 u1_u0_u7_U84 (.ZN( u1_out0_21 ) , .A4( u1_u0_u7_n157 ) , .A3( u1_u0_u7_n158 ) , .A2( u1_u0_u7_n159 ) , .A1( u1_u0_u7_n160 ) );
  OAI21_X1 u1_u0_u7_U85 (.B1( u1_u0_u7_n145 ) , .ZN( u1_u0_u7_n160 ) , .A( u1_u0_u7_n161 ) , .B2( u1_u0_u7_n177 ) );
  AOI22_X1 u1_u0_u7_U86 (.B2( u1_u0_u7_n149 ) , .B1( u1_u0_u7_n150 ) , .A2( u1_u0_u7_n151 ) , .A1( u1_u0_u7_n152 ) , .ZN( u1_u0_u7_n158 ) );
  NAND4_X1 u1_u0_u7_U87 (.ZN( u1_out0_15 ) , .A4( u1_u0_u7_n142 ) , .A3( u1_u0_u7_n143 ) , .A2( u1_u0_u7_n144 ) , .A1( u1_u0_u7_n178 ) );
  OR2_X1 u1_u0_u7_U88 (.A2( u1_u0_u7_n125 ) , .A1( u1_u0_u7_n129 ) , .ZN( u1_u0_u7_n144 ) );
  AOI22_X1 u1_u0_u7_U89 (.A2( u1_u0_u7_n126 ) , .ZN( u1_u0_u7_n143 ) , .B2( u1_u0_u7_n165 ) , .B1( u1_u0_u7_n173 ) , .A1( u1_u0_u7_n174 ) );
  AND3_X1 u1_u0_u7_U9 (.A3( u1_u0_u7_n110 ) , .A2( u1_u0_u7_n127 ) , .A1( u1_u0_u7_n132 ) , .ZN( u1_u0_u7_n92 ) );
  INV_X1 u1_u0_u7_U90 (.A( u1_u0_X_43 ) , .ZN( u1_u0_u7_n167 ) );
  AOI211_X1 u1_u0_u7_U91 (.B( u1_u0_u7_n154 ) , .A( u1_u0_u7_n155 ) , .C1( u1_u0_u7_n156 ) , .ZN( u1_u0_u7_n157 ) , .C2( u1_u0_u7_n172 ) );
  OAI211_X1 u1_u0_u7_U92 (.B( u1_u0_u7_n122 ) , .A( u1_u0_u7_n123 ) , .C2( u1_u0_u7_n124 ) , .ZN( u1_u0_u7_n154 ) , .C1( u1_u0_u7_n162 ) );
  AOI222_X1 u1_u0_u7_U93 (.ZN( u1_u0_u7_n122 ) , .C2( u1_u0_u7_n126 ) , .C1( u1_u0_u7_n145 ) , .B1( u1_u0_u7_n161 ) , .A2( u1_u0_u7_n165 ) , .B2( u1_u0_u7_n170 ) , .A1( u1_u0_u7_n176 ) );
  INV_X1 u1_u0_u7_U94 (.A( u1_u0_u7_n111 ) , .ZN( u1_u0_u7_n170 ) );
  NAND3_X1 u1_u0_u7_U95 (.A3( u1_u0_u7_n146 ) , .A2( u1_u0_u7_n147 ) , .A1( u1_u0_u7_n148 ) , .ZN( u1_u0_u7_n151 ) );
  NAND3_X1 u1_u0_u7_U96 (.A3( u1_u0_u7_n131 ) , .A2( u1_u0_u7_n132 ) , .A1( u1_u0_u7_n133 ) , .ZN( u1_u0_u7_n135 ) );
  XOR2_X1 u1_u10_U11 (.B( u1_K11_44 ) , .A( u1_R9_29 ) , .Z( u1_u10_X_44 ) );
  XOR2_X1 u1_u10_U12 (.B( u1_K11_43 ) , .A( u1_R9_28 ) , .Z( u1_u10_X_43 ) );
  XOR2_X1 u1_u10_U13 (.B( u1_K11_42 ) , .A( u1_R9_29 ) , .Z( u1_u10_X_42 ) );
  XOR2_X1 u1_u10_U14 (.B( u1_K11_41 ) , .A( u1_R9_28 ) , .Z( u1_u10_X_41 ) );
  XOR2_X1 u1_u10_U15 (.B( u1_K11_40 ) , .A( u1_R9_27 ) , .Z( u1_u10_X_40 ) );
  XOR2_X1 u1_u10_U17 (.B( u1_K11_39 ) , .A( u1_R9_26 ) , .Z( u1_u10_X_39 ) );
  XOR2_X1 u1_u10_U18 (.B( u1_K11_38 ) , .A( u1_R9_25 ) , .Z( u1_u10_X_38 ) );
  XOR2_X1 u1_u10_U19 (.B( u1_K11_37 ) , .A( u1_R9_24 ) , .Z( u1_u10_X_37 ) );
  XOR2_X1 u1_u10_U20 (.B( u1_K11_36 ) , .A( u1_R9_25 ) , .Z( u1_u10_X_36 ) );
  XOR2_X1 u1_u10_U21 (.B( u1_K11_35 ) , .A( u1_R9_24 ) , .Z( u1_u10_X_35 ) );
  XOR2_X1 u1_u10_U27 (.B( u1_K11_2 ) , .A( u1_R9_1 ) , .Z( u1_u10_X_2 ) );
  XOR2_X1 u1_u10_U31 (.B( u1_K11_26 ) , .A( u1_R9_17 ) , .Z( u1_u10_X_26 ) );
  XOR2_X1 u1_u10_U32 (.B( u1_K11_25 ) , .A( u1_R9_16 ) , .Z( u1_u10_X_25 ) );
  XOR2_X1 u1_u10_U33 (.B( u1_K11_24 ) , .A( u1_R9_17 ) , .Z( u1_u10_X_24 ) );
  XOR2_X1 u1_u10_U34 (.B( u1_K11_23 ) , .A( u1_R9_16 ) , .Z( u1_u10_X_23 ) );
  XOR2_X1 u1_u10_U38 (.B( u1_K11_1 ) , .A( u1_R9_32 ) , .Z( u1_u10_X_1 ) );
  XOR2_X1 u1_u10_U44 (.B( u1_K11_14 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_14 ) );
  XOR2_X1 u1_u10_U45 (.B( u1_K11_13 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_13 ) );
  XOR2_X1 u1_u10_U46 (.B( u1_K11_12 ) , .A( u1_R9_9 ) , .Z( u1_u10_X_12 ) );
  XOR2_X1 u1_u10_U47 (.B( u1_K11_11 ) , .A( u1_R9_8 ) , .Z( u1_u10_X_11 ) );
  XOR2_X1 u1_u10_U7 (.B( u1_K11_48 ) , .A( u1_R9_1 ) , .Z( u1_u10_X_48 ) );
  XOR2_X1 u1_u10_U8 (.B( u1_K11_47 ) , .A( u1_R9_32 ) , .Z( u1_u10_X_47 ) );
  AOI22_X1 u1_u10_u6_U10 (.A2( u1_u10_u6_n151 ) , .B2( u1_u10_u6_n161 ) , .A1( u1_u10_u6_n167 ) , .B1( u1_u10_u6_n170 ) , .ZN( u1_u10_u6_n89 ) );
  AOI21_X1 u1_u10_u6_U11 (.B1( u1_u10_u6_n107 ) , .B2( u1_u10_u6_n132 ) , .A( u1_u10_u6_n158 ) , .ZN( u1_u10_u6_n88 ) );
  AOI21_X1 u1_u10_u6_U12 (.B2( u1_u10_u6_n147 ) , .B1( u1_u10_u6_n148 ) , .ZN( u1_u10_u6_n149 ) , .A( u1_u10_u6_n158 ) );
  AOI21_X1 u1_u10_u6_U13 (.ZN( u1_u10_u6_n106 ) , .A( u1_u10_u6_n142 ) , .B2( u1_u10_u6_n159 ) , .B1( u1_u10_u6_n164 ) );
  INV_X1 u1_u10_u6_U14 (.A( u1_u10_u6_n155 ) , .ZN( u1_u10_u6_n161 ) );
  INV_X1 u1_u10_u6_U15 (.A( u1_u10_u6_n128 ) , .ZN( u1_u10_u6_n164 ) );
  NAND2_X1 u1_u10_u6_U16 (.ZN( u1_u10_u6_n110 ) , .A1( u1_u10_u6_n122 ) , .A2( u1_u10_u6_n129 ) );
  NAND2_X1 u1_u10_u6_U17 (.ZN( u1_u10_u6_n124 ) , .A2( u1_u10_u6_n146 ) , .A1( u1_u10_u6_n148 ) );
  INV_X1 u1_u10_u6_U18 (.A( u1_u10_u6_n132 ) , .ZN( u1_u10_u6_n171 ) );
  AND2_X1 u1_u10_u6_U19 (.A1( u1_u10_u6_n100 ) , .ZN( u1_u10_u6_n130 ) , .A2( u1_u10_u6_n147 ) );
  INV_X1 u1_u10_u6_U20 (.A( u1_u10_u6_n127 ) , .ZN( u1_u10_u6_n173 ) );
  INV_X1 u1_u10_u6_U21 (.A( u1_u10_u6_n121 ) , .ZN( u1_u10_u6_n167 ) );
  INV_X1 u1_u10_u6_U22 (.A( u1_u10_u6_n100 ) , .ZN( u1_u10_u6_n169 ) );
  INV_X1 u1_u10_u6_U23 (.A( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n170 ) );
  INV_X1 u1_u10_u6_U24 (.A( u1_u10_u6_n113 ) , .ZN( u1_u10_u6_n168 ) );
  AND2_X1 u1_u10_u6_U25 (.A1( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n119 ) , .ZN( u1_u10_u6_n133 ) );
  AND2_X1 u1_u10_u6_U26 (.A2( u1_u10_u6_n121 ) , .A1( u1_u10_u6_n122 ) , .ZN( u1_u10_u6_n131 ) );
  AND3_X1 u1_u10_u6_U27 (.ZN( u1_u10_u6_n120 ) , .A2( u1_u10_u6_n127 ) , .A1( u1_u10_u6_n132 ) , .A3( u1_u10_u6_n145 ) );
  INV_X1 u1_u10_u6_U28 (.A( u1_u10_u6_n146 ) , .ZN( u1_u10_u6_n163 ) );
  AOI222_X1 u1_u10_u6_U29 (.ZN( u1_u10_u6_n114 ) , .A1( u1_u10_u6_n118 ) , .A2( u1_u10_u6_n126 ) , .B2( u1_u10_u6_n151 ) , .C2( u1_u10_u6_n159 ) , .C1( u1_u10_u6_n168 ) , .B1( u1_u10_u6_n169 ) );
  INV_X1 u1_u10_u6_U3 (.A( u1_u10_u6_n110 ) , .ZN( u1_u10_u6_n166 ) );
  NOR2_X1 u1_u10_u6_U30 (.A1( u1_u10_u6_n162 ) , .A2( u1_u10_u6_n165 ) , .ZN( u1_u10_u6_n98 ) );
  AOI211_X1 u1_u10_u6_U31 (.B( u1_u10_u6_n134 ) , .A( u1_u10_u6_n135 ) , .C1( u1_u10_u6_n136 ) , .ZN( u1_u10_u6_n137 ) , .C2( u1_u10_u6_n151 ) );
  NAND4_X1 u1_u10_u6_U32 (.A4( u1_u10_u6_n127 ) , .A3( u1_u10_u6_n128 ) , .A2( u1_u10_u6_n129 ) , .A1( u1_u10_u6_n130 ) , .ZN( u1_u10_u6_n136 ) );
  AOI21_X1 u1_u10_u6_U33 (.B2( u1_u10_u6_n132 ) , .B1( u1_u10_u6_n133 ) , .ZN( u1_u10_u6_n134 ) , .A( u1_u10_u6_n158 ) );
  AOI21_X1 u1_u10_u6_U34 (.B1( u1_u10_u6_n131 ) , .ZN( u1_u10_u6_n135 ) , .A( u1_u10_u6_n144 ) , .B2( u1_u10_u6_n146 ) );
  NAND2_X1 u1_u10_u6_U35 (.A1( u1_u10_u6_n144 ) , .ZN( u1_u10_u6_n151 ) , .A2( u1_u10_u6_n158 ) );
  NAND2_X1 u1_u10_u6_U36 (.ZN( u1_u10_u6_n132 ) , .A1( u1_u10_u6_n91 ) , .A2( u1_u10_u6_n97 ) );
  AOI22_X1 u1_u10_u6_U37 (.B2( u1_u10_u6_n110 ) , .B1( u1_u10_u6_n111 ) , .A1( u1_u10_u6_n112 ) , .ZN( u1_u10_u6_n115 ) , .A2( u1_u10_u6_n161 ) );
  NAND4_X1 u1_u10_u6_U38 (.A3( u1_u10_u6_n109 ) , .ZN( u1_u10_u6_n112 ) , .A4( u1_u10_u6_n132 ) , .A2( u1_u10_u6_n147 ) , .A1( u1_u10_u6_n166 ) );
  NOR2_X1 u1_u10_u6_U39 (.ZN( u1_u10_u6_n109 ) , .A1( u1_u10_u6_n170 ) , .A2( u1_u10_u6_n173 ) );
  INV_X1 u1_u10_u6_U4 (.A( u1_u10_u6_n142 ) , .ZN( u1_u10_u6_n174 ) );
  NOR2_X1 u1_u10_u6_U40 (.A2( u1_u10_u6_n126 ) , .ZN( u1_u10_u6_n155 ) , .A1( u1_u10_u6_n160 ) );
  NAND2_X1 u1_u10_u6_U41 (.ZN( u1_u10_u6_n146 ) , .A2( u1_u10_u6_n94 ) , .A1( u1_u10_u6_n99 ) );
  AOI21_X1 u1_u10_u6_U42 (.A( u1_u10_u6_n144 ) , .B2( u1_u10_u6_n145 ) , .B1( u1_u10_u6_n146 ) , .ZN( u1_u10_u6_n150 ) );
  INV_X1 u1_u10_u6_U43 (.A( u1_u10_u6_n111 ) , .ZN( u1_u10_u6_n158 ) );
  NAND2_X1 u1_u10_u6_U44 (.ZN( u1_u10_u6_n127 ) , .A1( u1_u10_u6_n91 ) , .A2( u1_u10_u6_n92 ) );
  NAND2_X1 u1_u10_u6_U45 (.ZN( u1_u10_u6_n129 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n96 ) );
  INV_X1 u1_u10_u6_U46 (.A( u1_u10_u6_n144 ) , .ZN( u1_u10_u6_n159 ) );
  NAND2_X1 u1_u10_u6_U47 (.ZN( u1_u10_u6_n145 ) , .A2( u1_u10_u6_n97 ) , .A1( u1_u10_u6_n98 ) );
  NAND2_X1 u1_u10_u6_U48 (.ZN( u1_u10_u6_n148 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n94 ) );
  NAND2_X1 u1_u10_u6_U49 (.ZN( u1_u10_u6_n108 ) , .A2( u1_u10_u6_n139 ) , .A1( u1_u10_u6_n144 ) );
  NAND2_X1 u1_u10_u6_U5 (.A2( u1_u10_u6_n143 ) , .ZN( u1_u10_u6_n152 ) , .A1( u1_u10_u6_n166 ) );
  NAND2_X1 u1_u10_u6_U50 (.ZN( u1_u10_u6_n121 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n97 ) );
  NAND2_X1 u1_u10_u6_U51 (.ZN( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n95 ) );
  AND2_X1 u1_u10_u6_U52 (.ZN( u1_u10_u6_n118 ) , .A2( u1_u10_u6_n91 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U53 (.ZN( u1_u10_u6_n147 ) , .A2( u1_u10_u6_n98 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U54 (.ZN( u1_u10_u6_n128 ) , .A1( u1_u10_u6_n94 ) , .A2( u1_u10_u6_n96 ) );
  NAND2_X1 u1_u10_u6_U55 (.ZN( u1_u10_u6_n119 ) , .A2( u1_u10_u6_n95 ) , .A1( u1_u10_u6_n99 ) );
  NAND2_X1 u1_u10_u6_U56 (.ZN( u1_u10_u6_n123 ) , .A2( u1_u10_u6_n91 ) , .A1( u1_u10_u6_n96 ) );
  NAND2_X1 u1_u10_u6_U57 (.ZN( u1_u10_u6_n100 ) , .A2( u1_u10_u6_n92 ) , .A1( u1_u10_u6_n98 ) );
  NAND2_X1 u1_u10_u6_U58 (.ZN( u1_u10_u6_n122 ) , .A1( u1_u10_u6_n94 ) , .A2( u1_u10_u6_n97 ) );
  INV_X1 u1_u10_u6_U59 (.A( u1_u10_u6_n139 ) , .ZN( u1_u10_u6_n160 ) );
  AOI22_X1 u1_u10_u6_U6 (.B2( u1_u10_u6_n101 ) , .A1( u1_u10_u6_n102 ) , .ZN( u1_u10_u6_n103 ) , .B1( u1_u10_u6_n160 ) , .A2( u1_u10_u6_n161 ) );
  NAND2_X1 u1_u10_u6_U60 (.ZN( u1_u10_u6_n113 ) , .A1( u1_u10_u6_n96 ) , .A2( u1_u10_u6_n98 ) );
  NOR2_X1 u1_u10_u6_U61 (.A2( u1_u10_X_40 ) , .A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n126 ) );
  NOR2_X1 u1_u10_u6_U62 (.A2( u1_u10_X_39 ) , .A1( u1_u10_X_42 ) , .ZN( u1_u10_u6_n92 ) );
  NOR2_X1 u1_u10_u6_U63 (.A2( u1_u10_X_39 ) , .A1( u1_u10_u6_n156 ) , .ZN( u1_u10_u6_n97 ) );
  NOR2_X1 u1_u10_u6_U64 (.A2( u1_u10_X_38 ) , .A1( u1_u10_u6_n165 ) , .ZN( u1_u10_u6_n95 ) );
  NOR2_X1 u1_u10_u6_U65 (.A2( u1_u10_X_41 ) , .ZN( u1_u10_u6_n111 ) , .A1( u1_u10_u6_n157 ) );
  NOR2_X1 u1_u10_u6_U66 (.A2( u1_u10_X_37 ) , .A1( u1_u10_u6_n162 ) , .ZN( u1_u10_u6_n94 ) );
  NOR2_X1 u1_u10_u6_U67 (.A2( u1_u10_X_37 ) , .A1( u1_u10_X_38 ) , .ZN( u1_u10_u6_n91 ) );
  NAND2_X1 u1_u10_u6_U68 (.A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n144 ) , .A2( u1_u10_u6_n157 ) );
  NAND2_X1 u1_u10_u6_U69 (.A2( u1_u10_X_40 ) , .A1( u1_u10_X_41 ) , .ZN( u1_u10_u6_n139 ) );
  NOR2_X1 u1_u10_u6_U7 (.A1( u1_u10_u6_n118 ) , .ZN( u1_u10_u6_n143 ) , .A2( u1_u10_u6_n168 ) );
  AND2_X1 u1_u10_u6_U70 (.A1( u1_u10_X_39 ) , .A2( u1_u10_u6_n156 ) , .ZN( u1_u10_u6_n96 ) );
  AND2_X1 u1_u10_u6_U71 (.A1( u1_u10_X_39 ) , .A2( u1_u10_X_42 ) , .ZN( u1_u10_u6_n99 ) );
  INV_X1 u1_u10_u6_U72 (.A( u1_u10_X_40 ) , .ZN( u1_u10_u6_n157 ) );
  INV_X1 u1_u10_u6_U73 (.A( u1_u10_X_37 ) , .ZN( u1_u10_u6_n165 ) );
  INV_X1 u1_u10_u6_U74 (.A( u1_u10_X_38 ) , .ZN( u1_u10_u6_n162 ) );
  INV_X1 u1_u10_u6_U75 (.A( u1_u10_X_42 ) , .ZN( u1_u10_u6_n156 ) );
  NAND4_X1 u1_u10_u6_U76 (.ZN( u1_out10_32 ) , .A4( u1_u10_u6_n103 ) , .A3( u1_u10_u6_n104 ) , .A2( u1_u10_u6_n105 ) , .A1( u1_u10_u6_n106 ) );
  AOI22_X1 u1_u10_u6_U77 (.ZN( u1_u10_u6_n105 ) , .A2( u1_u10_u6_n108 ) , .A1( u1_u10_u6_n118 ) , .B2( u1_u10_u6_n126 ) , .B1( u1_u10_u6_n171 ) );
  AOI22_X1 u1_u10_u6_U78 (.ZN( u1_u10_u6_n104 ) , .A1( u1_u10_u6_n111 ) , .B1( u1_u10_u6_n124 ) , .B2( u1_u10_u6_n151 ) , .A2( u1_u10_u6_n93 ) );
  NAND4_X1 u1_u10_u6_U79 (.ZN( u1_out10_12 ) , .A4( u1_u10_u6_n114 ) , .A3( u1_u10_u6_n115 ) , .A2( u1_u10_u6_n116 ) , .A1( u1_u10_u6_n117 ) );
  INV_X1 u1_u10_u6_U8 (.ZN( u1_u10_u6_n172 ) , .A( u1_u10_u6_n88 ) );
  OAI22_X1 u1_u10_u6_U80 (.B2( u1_u10_u6_n111 ) , .ZN( u1_u10_u6_n116 ) , .B1( u1_u10_u6_n126 ) , .A2( u1_u10_u6_n164 ) , .A1( u1_u10_u6_n167 ) );
  OAI21_X1 u1_u10_u6_U81 (.A( u1_u10_u6_n108 ) , .ZN( u1_u10_u6_n117 ) , .B2( u1_u10_u6_n141 ) , .B1( u1_u10_u6_n163 ) );
  OAI211_X1 u1_u10_u6_U82 (.ZN( u1_out10_7 ) , .B( u1_u10_u6_n153 ) , .C2( u1_u10_u6_n154 ) , .C1( u1_u10_u6_n155 ) , .A( u1_u10_u6_n174 ) );
  NOR3_X1 u1_u10_u6_U83 (.A1( u1_u10_u6_n141 ) , .ZN( u1_u10_u6_n154 ) , .A3( u1_u10_u6_n164 ) , .A2( u1_u10_u6_n171 ) );
  AOI211_X1 u1_u10_u6_U84 (.B( u1_u10_u6_n149 ) , .A( u1_u10_u6_n150 ) , .C2( u1_u10_u6_n151 ) , .C1( u1_u10_u6_n152 ) , .ZN( u1_u10_u6_n153 ) );
  OAI211_X1 u1_u10_u6_U85 (.ZN( u1_out10_22 ) , .B( u1_u10_u6_n137 ) , .A( u1_u10_u6_n138 ) , .C2( u1_u10_u6_n139 ) , .C1( u1_u10_u6_n140 ) );
  AOI22_X1 u1_u10_u6_U86 (.B1( u1_u10_u6_n124 ) , .A2( u1_u10_u6_n125 ) , .A1( u1_u10_u6_n126 ) , .ZN( u1_u10_u6_n138 ) , .B2( u1_u10_u6_n161 ) );
  AND4_X1 u1_u10_u6_U87 (.A3( u1_u10_u6_n119 ) , .A1( u1_u10_u6_n120 ) , .A4( u1_u10_u6_n129 ) , .ZN( u1_u10_u6_n140 ) , .A2( u1_u10_u6_n143 ) );
  NAND3_X1 u1_u10_u6_U88 (.A2( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n125 ) , .A1( u1_u10_u6_n130 ) , .A3( u1_u10_u6_n131 ) );
  NAND3_X1 u1_u10_u6_U89 (.A3( u1_u10_u6_n133 ) , .ZN( u1_u10_u6_n141 ) , .A1( u1_u10_u6_n145 ) , .A2( u1_u10_u6_n148 ) );
  OAI21_X1 u1_u10_u6_U9 (.A( u1_u10_u6_n159 ) , .B1( u1_u10_u6_n169 ) , .B2( u1_u10_u6_n173 ) , .ZN( u1_u10_u6_n90 ) );
  NAND3_X1 u1_u10_u6_U90 (.ZN( u1_u10_u6_n101 ) , .A3( u1_u10_u6_n107 ) , .A2( u1_u10_u6_n121 ) , .A1( u1_u10_u6_n127 ) );
  NAND3_X1 u1_u10_u6_U91 (.ZN( u1_u10_u6_n102 ) , .A3( u1_u10_u6_n130 ) , .A2( u1_u10_u6_n145 ) , .A1( u1_u10_u6_n166 ) );
  NAND3_X1 u1_u10_u6_U92 (.A3( u1_u10_u6_n113 ) , .A1( u1_u10_u6_n119 ) , .A2( u1_u10_u6_n123 ) , .ZN( u1_u10_u6_n93 ) );
  NAND3_X1 u1_u10_u6_U93 (.ZN( u1_u10_u6_n142 ) , .A2( u1_u10_u6_n172 ) , .A3( u1_u10_u6_n89 ) , .A1( u1_u10_u6_n90 ) );
  XOR2_X1 u1_u11_U1 (.B( u1_K12_9 ) , .A( u1_R10_6 ) , .Z( u1_u11_X_9 ) );
  XOR2_X1 u1_u11_U11 (.B( u1_K12_44 ) , .A( u1_R10_29 ) , .Z( u1_u11_X_44 ) );
  XOR2_X1 u1_u11_U12 (.B( u1_K12_43 ) , .A( u1_R10_28 ) , .Z( u1_u11_X_43 ) );
  XOR2_X1 u1_u11_U13 (.B( u1_K12_42 ) , .A( u1_R10_29 ) , .Z( u1_u11_X_42 ) );
  XOR2_X1 u1_u11_U14 (.B( u1_K12_41 ) , .A( u1_R10_28 ) , .Z( u1_u11_X_41 ) );
  XOR2_X1 u1_u11_U18 (.B( u1_K12_38 ) , .A( u1_R10_25 ) , .Z( u1_u11_X_38 ) );
  XOR2_X1 u1_u11_U19 (.B( u1_K12_37 ) , .A( u1_R10_24 ) , .Z( u1_u11_X_37 ) );
  XOR2_X1 u1_u11_U2 (.B( u1_K12_8 ) , .A( u1_R10_5 ) , .Z( u1_u11_X_8 ) );
  XOR2_X1 u1_u11_U20 (.B( u1_K12_36 ) , .A( u1_R10_25 ) , .Z( u1_u11_X_36 ) );
  XOR2_X1 u1_u11_U21 (.B( u1_K12_35 ) , .A( u1_R10_24 ) , .Z( u1_u11_X_35 ) );
  XOR2_X1 u1_u11_U24 (.B( u1_K12_32 ) , .A( u1_R10_21 ) , .Z( u1_u11_X_32 ) );
  XOR2_X1 u1_u11_U25 (.B( u1_K12_31 ) , .A( u1_R10_20 ) , .Z( u1_u11_X_31 ) );
  XOR2_X1 u1_u11_U26 (.B( u1_K12_30 ) , .A( u1_R10_21 ) , .Z( u1_u11_X_30 ) );
  XOR2_X1 u1_u11_U27 (.B( u1_K12_2 ) , .A( u1_R10_1 ) , .Z( u1_u11_X_2 ) );
  XOR2_X1 u1_u11_U28 (.B( u1_K12_29 ) , .A( u1_R10_20 ) , .Z( u1_u11_X_29 ) );
  XOR2_X1 u1_u11_U29 (.B( u1_K12_28 ) , .A( u1_R10_19 ) , .Z( u1_u11_X_28 ) );
  XOR2_X1 u1_u11_U3 (.B( u1_K12_7 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_7 ) );
  XOR2_X1 u1_u11_U30 (.B( u1_K12_27 ) , .A( u1_R10_18 ) , .Z( u1_u11_X_27 ) );
  XOR2_X1 u1_u11_U31 (.B( u1_K12_26 ) , .A( u1_R10_17 ) , .Z( u1_u11_X_26 ) );
  XOR2_X1 u1_u11_U32 (.B( u1_K12_25 ) , .A( u1_R10_16 ) , .Z( u1_u11_X_25 ) );
  XOR2_X1 u1_u11_U33 (.B( u1_K12_24 ) , .A( u1_R10_17 ) , .Z( u1_u11_X_24 ) );
  XOR2_X1 u1_u11_U34 (.B( u1_K12_23 ) , .A( u1_R10_16 ) , .Z( u1_u11_X_23 ) );
  XOR2_X1 u1_u11_U35 (.B( u1_K12_22 ) , .A( u1_R10_15 ) , .Z( u1_u11_X_22 ) );
  XOR2_X1 u1_u11_U36 (.B( u1_K12_21 ) , .A( u1_R10_14 ) , .Z( u1_u11_X_21 ) );
  XOR2_X1 u1_u11_U37 (.B( u1_K12_20 ) , .A( u1_R10_13 ) , .Z( u1_u11_X_20 ) );
  XOR2_X1 u1_u11_U38 (.B( u1_K12_1 ) , .A( u1_R10_32 ) , .Z( u1_u11_X_1 ) );
  XOR2_X1 u1_u11_U39 (.B( u1_K12_19 ) , .A( u1_R10_12 ) , .Z( u1_u11_X_19 ) );
  XOR2_X1 u1_u11_U4 (.B( u1_K12_6 ) , .A( u1_R10_5 ) , .Z( u1_u11_X_6 ) );
  XOR2_X1 u1_u11_U40 (.B( u1_K12_18 ) , .A( u1_R10_13 ) , .Z( u1_u11_X_18 ) );
  XOR2_X1 u1_u11_U41 (.B( u1_K12_17 ) , .A( u1_R10_12 ) , .Z( u1_u11_X_17 ) );
  XOR2_X1 u1_u11_U42 (.B( u1_K12_16 ) , .A( u1_R10_11 ) , .Z( u1_u11_X_16 ) );
  XOR2_X1 u1_u11_U43 (.B( u1_K12_15 ) , .A( u1_R10_10 ) , .Z( u1_u11_X_15 ) );
  XOR2_X1 u1_u11_U44 (.B( u1_K12_14 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_14 ) );
  XOR2_X1 u1_u11_U45 (.B( u1_K12_13 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_13 ) );
  XOR2_X1 u1_u11_U46 (.B( u1_K12_12 ) , .A( u1_R10_9 ) , .Z( u1_u11_X_12 ) );
  XOR2_X1 u1_u11_U47 (.B( u1_K12_11 ) , .A( u1_R10_8 ) , .Z( u1_u11_X_11 ) );
  XOR2_X1 u1_u11_U48 (.B( u1_K12_10 ) , .A( u1_R10_7 ) , .Z( u1_u11_X_10 ) );
  XOR2_X1 u1_u11_U5 (.B( u1_K12_5 ) , .A( u1_R10_4 ) , .Z( u1_u11_X_5 ) );
  XOR2_X1 u1_u11_U7 (.B( u1_K12_48 ) , .A( u1_R10_1 ) , .Z( u1_u11_X_48 ) );
  XOR2_X1 u1_u11_U8 (.B( u1_K12_47 ) , .A( u1_R10_32 ) , .Z( u1_u11_X_47 ) );
  NOR2_X1 u1_u11_u1_U10 (.A1( u1_u11_u1_n112 ) , .A2( u1_u11_u1_n116 ) , .ZN( u1_u11_u1_n118 ) );
  NAND3_X1 u1_u11_u1_U100 (.ZN( u1_u11_u1_n113 ) , .A1( u1_u11_u1_n120 ) , .A3( u1_u11_u1_n133 ) , .A2( u1_u11_u1_n155 ) );
  OAI21_X1 u1_u11_u1_U11 (.ZN( u1_u11_u1_n101 ) , .B1( u1_u11_u1_n141 ) , .A( u1_u11_u1_n146 ) , .B2( u1_u11_u1_n183 ) );
  AOI21_X1 u1_u11_u1_U12 (.B2( u1_u11_u1_n155 ) , .B1( u1_u11_u1_n156 ) , .ZN( u1_u11_u1_n157 ) , .A( u1_u11_u1_n174 ) );
  NAND2_X1 u1_u11_u1_U13 (.ZN( u1_u11_u1_n140 ) , .A2( u1_u11_u1_n150 ) , .A1( u1_u11_u1_n155 ) );
  NAND2_X1 u1_u11_u1_U14 (.A1( u1_u11_u1_n131 ) , .ZN( u1_u11_u1_n147 ) , .A2( u1_u11_u1_n153 ) );
  INV_X1 u1_u11_u1_U15 (.A( u1_u11_u1_n139 ) , .ZN( u1_u11_u1_n174 ) );
  OR4_X1 u1_u11_u1_U16 (.A4( u1_u11_u1_n106 ) , .A3( u1_u11_u1_n107 ) , .ZN( u1_u11_u1_n108 ) , .A1( u1_u11_u1_n117 ) , .A2( u1_u11_u1_n184 ) );
  AOI21_X1 u1_u11_u1_U17 (.ZN( u1_u11_u1_n106 ) , .A( u1_u11_u1_n112 ) , .B1( u1_u11_u1_n154 ) , .B2( u1_u11_u1_n156 ) );
  AOI21_X1 u1_u11_u1_U18 (.ZN( u1_u11_u1_n107 ) , .B1( u1_u11_u1_n134 ) , .B2( u1_u11_u1_n149 ) , .A( u1_u11_u1_n174 ) );
  INV_X1 u1_u11_u1_U19 (.A( u1_u11_u1_n101 ) , .ZN( u1_u11_u1_n184 ) );
  INV_X1 u1_u11_u1_U20 (.A( u1_u11_u1_n112 ) , .ZN( u1_u11_u1_n171 ) );
  NAND2_X1 u1_u11_u1_U21 (.ZN( u1_u11_u1_n141 ) , .A1( u1_u11_u1_n153 ) , .A2( u1_u11_u1_n156 ) );
  AND2_X1 u1_u11_u1_U22 (.A1( u1_u11_u1_n123 ) , .ZN( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n161 ) );
  NAND2_X1 u1_u11_u1_U23 (.A2( u1_u11_u1_n115 ) , .A1( u1_u11_u1_n116 ) , .ZN( u1_u11_u1_n148 ) );
  NAND2_X1 u1_u11_u1_U24 (.A2( u1_u11_u1_n133 ) , .A1( u1_u11_u1_n135 ) , .ZN( u1_u11_u1_n159 ) );
  NAND2_X1 u1_u11_u1_U25 (.A2( u1_u11_u1_n115 ) , .A1( u1_u11_u1_n120 ) , .ZN( u1_u11_u1_n132 ) );
  INV_X1 u1_u11_u1_U26 (.A( u1_u11_u1_n154 ) , .ZN( u1_u11_u1_n178 ) );
  INV_X1 u1_u11_u1_U27 (.A( u1_u11_u1_n151 ) , .ZN( u1_u11_u1_n183 ) );
  AND2_X1 u1_u11_u1_U28 (.A1( u1_u11_u1_n129 ) , .A2( u1_u11_u1_n133 ) , .ZN( u1_u11_u1_n149 ) );
  INV_X1 u1_u11_u1_U29 (.A( u1_u11_u1_n131 ) , .ZN( u1_u11_u1_n180 ) );
  INV_X1 u1_u11_u1_U3 (.A( u1_u11_u1_n159 ) , .ZN( u1_u11_u1_n182 ) );
  OAI221_X1 u1_u11_u1_U30 (.A( u1_u11_u1_n119 ) , .C2( u1_u11_u1_n129 ) , .ZN( u1_u11_u1_n138 ) , .B2( u1_u11_u1_n152 ) , .C1( u1_u11_u1_n174 ) , .B1( u1_u11_u1_n187 ) );
  INV_X1 u1_u11_u1_U31 (.A( u1_u11_u1_n148 ) , .ZN( u1_u11_u1_n187 ) );
  AOI211_X1 u1_u11_u1_U32 (.B( u1_u11_u1_n117 ) , .A( u1_u11_u1_n118 ) , .ZN( u1_u11_u1_n119 ) , .C2( u1_u11_u1_n146 ) , .C1( u1_u11_u1_n159 ) );
  NOR2_X1 u1_u11_u1_U33 (.A1( u1_u11_u1_n168 ) , .A2( u1_u11_u1_n176 ) , .ZN( u1_u11_u1_n98 ) );
  AOI211_X1 u1_u11_u1_U34 (.B( u1_u11_u1_n162 ) , .A( u1_u11_u1_n163 ) , .C2( u1_u11_u1_n164 ) , .ZN( u1_u11_u1_n165 ) , .C1( u1_u11_u1_n171 ) );
  AOI21_X1 u1_u11_u1_U35 (.A( u1_u11_u1_n160 ) , .B2( u1_u11_u1_n161 ) , .ZN( u1_u11_u1_n162 ) , .B1( u1_u11_u1_n182 ) );
  OR2_X1 u1_u11_u1_U36 (.A2( u1_u11_u1_n157 ) , .A1( u1_u11_u1_n158 ) , .ZN( u1_u11_u1_n163 ) );
  NAND2_X1 u1_u11_u1_U37 (.A1( u1_u11_u1_n128 ) , .ZN( u1_u11_u1_n146 ) , .A2( u1_u11_u1_n160 ) );
  NAND2_X1 u1_u11_u1_U38 (.A2( u1_u11_u1_n112 ) , .ZN( u1_u11_u1_n139 ) , .A1( u1_u11_u1_n152 ) );
  NAND2_X1 u1_u11_u1_U39 (.A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n156 ) , .A2( u1_u11_u1_n99 ) );
  AOI221_X1 u1_u11_u1_U4 (.A( u1_u11_u1_n138 ) , .C2( u1_u11_u1_n139 ) , .C1( u1_u11_u1_n140 ) , .B2( u1_u11_u1_n141 ) , .ZN( u1_u11_u1_n142 ) , .B1( u1_u11_u1_n175 ) );
  AOI221_X1 u1_u11_u1_U40 (.B1( u1_u11_u1_n140 ) , .ZN( u1_u11_u1_n167 ) , .B2( u1_u11_u1_n172 ) , .C2( u1_u11_u1_n175 ) , .C1( u1_u11_u1_n178 ) , .A( u1_u11_u1_n188 ) );
  INV_X1 u1_u11_u1_U41 (.ZN( u1_u11_u1_n188 ) , .A( u1_u11_u1_n97 ) );
  AOI211_X1 u1_u11_u1_U42 (.A( u1_u11_u1_n118 ) , .C1( u1_u11_u1_n132 ) , .C2( u1_u11_u1_n139 ) , .B( u1_u11_u1_n96 ) , .ZN( u1_u11_u1_n97 ) );
  AOI21_X1 u1_u11_u1_U43 (.B2( u1_u11_u1_n121 ) , .B1( u1_u11_u1_n135 ) , .A( u1_u11_u1_n152 ) , .ZN( u1_u11_u1_n96 ) );
  NOR2_X1 u1_u11_u1_U44 (.ZN( u1_u11_u1_n117 ) , .A1( u1_u11_u1_n121 ) , .A2( u1_u11_u1_n160 ) );
  OAI21_X1 u1_u11_u1_U45 (.B2( u1_u11_u1_n123 ) , .ZN( u1_u11_u1_n145 ) , .B1( u1_u11_u1_n160 ) , .A( u1_u11_u1_n185 ) );
  INV_X1 u1_u11_u1_U46 (.A( u1_u11_u1_n122 ) , .ZN( u1_u11_u1_n185 ) );
  AOI21_X1 u1_u11_u1_U47 (.B2( u1_u11_u1_n120 ) , .B1( u1_u11_u1_n121 ) , .ZN( u1_u11_u1_n122 ) , .A( u1_u11_u1_n128 ) );
  AOI21_X1 u1_u11_u1_U48 (.A( u1_u11_u1_n128 ) , .B2( u1_u11_u1_n129 ) , .ZN( u1_u11_u1_n130 ) , .B1( u1_u11_u1_n150 ) );
  NAND2_X1 u1_u11_u1_U49 (.ZN( u1_u11_u1_n112 ) , .A1( u1_u11_u1_n169 ) , .A2( u1_u11_u1_n170 ) );
  AOI211_X1 u1_u11_u1_U5 (.ZN( u1_u11_u1_n124 ) , .A( u1_u11_u1_n138 ) , .C2( u1_u11_u1_n139 ) , .B( u1_u11_u1_n145 ) , .C1( u1_u11_u1_n147 ) );
  NAND2_X1 u1_u11_u1_U50 (.ZN( u1_u11_u1_n129 ) , .A2( u1_u11_u1_n95 ) , .A1( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U51 (.A1( u1_u11_u1_n102 ) , .ZN( u1_u11_u1_n154 ) , .A2( u1_u11_u1_n99 ) );
  NAND2_X1 u1_u11_u1_U52 (.A2( u1_u11_u1_n100 ) , .ZN( u1_u11_u1_n135 ) , .A1( u1_u11_u1_n99 ) );
  AOI21_X1 u1_u11_u1_U53 (.A( u1_u11_u1_n152 ) , .B2( u1_u11_u1_n153 ) , .B1( u1_u11_u1_n154 ) , .ZN( u1_u11_u1_n158 ) );
  INV_X1 u1_u11_u1_U54 (.A( u1_u11_u1_n160 ) , .ZN( u1_u11_u1_n175 ) );
  NAND2_X1 u1_u11_u1_U55 (.A1( u1_u11_u1_n100 ) , .ZN( u1_u11_u1_n116 ) , .A2( u1_u11_u1_n95 ) );
  NAND2_X1 u1_u11_u1_U56 (.A1( u1_u11_u1_n102 ) , .ZN( u1_u11_u1_n131 ) , .A2( u1_u11_u1_n95 ) );
  NAND2_X1 u1_u11_u1_U57 (.A2( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n121 ) , .A1( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U58 (.A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n153 ) , .A2( u1_u11_u1_n98 ) );
  NAND2_X1 u1_u11_u1_U59 (.A2( u1_u11_u1_n104 ) , .A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n133 ) );
  AOI22_X1 u1_u11_u1_U6 (.B2( u1_u11_u1_n113 ) , .A2( u1_u11_u1_n114 ) , .ZN( u1_u11_u1_n125 ) , .A1( u1_u11_u1_n171 ) , .B1( u1_u11_u1_n173 ) );
  NAND2_X1 u1_u11_u1_U60 (.ZN( u1_u11_u1_n150 ) , .A2( u1_u11_u1_n98 ) , .A1( u1_u11_u1_n99 ) );
  NAND2_X1 u1_u11_u1_U61 (.A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n155 ) , .A2( u1_u11_u1_n95 ) );
  OAI21_X1 u1_u11_u1_U62 (.ZN( u1_u11_u1_n109 ) , .B1( u1_u11_u1_n129 ) , .B2( u1_u11_u1_n160 ) , .A( u1_u11_u1_n167 ) );
  NAND2_X1 u1_u11_u1_U63 (.A2( u1_u11_u1_n100 ) , .A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n120 ) );
  NAND2_X1 u1_u11_u1_U64 (.A1( u1_u11_u1_n102 ) , .A2( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n115 ) );
  NAND2_X1 u1_u11_u1_U65 (.A2( u1_u11_u1_n100 ) , .A1( u1_u11_u1_n104 ) , .ZN( u1_u11_u1_n151 ) );
  NAND2_X1 u1_u11_u1_U66 (.A2( u1_u11_u1_n103 ) , .A1( u1_u11_u1_n105 ) , .ZN( u1_u11_u1_n161 ) );
  INV_X1 u1_u11_u1_U67 (.A( u1_u11_u1_n152 ) , .ZN( u1_u11_u1_n173 ) );
  INV_X1 u1_u11_u1_U68 (.A( u1_u11_u1_n128 ) , .ZN( u1_u11_u1_n172 ) );
  NAND2_X1 u1_u11_u1_U69 (.A2( u1_u11_u1_n102 ) , .A1( u1_u11_u1_n103 ) , .ZN( u1_u11_u1_n123 ) );
  NAND2_X1 u1_u11_u1_U7 (.ZN( u1_u11_u1_n114 ) , .A1( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n156 ) );
  NOR2_X1 u1_u11_u1_U70 (.A2( u1_u11_X_7 ) , .A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n95 ) );
  NOR2_X1 u1_u11_u1_U71 (.A1( u1_u11_X_12 ) , .A2( u1_u11_X_9 ) , .ZN( u1_u11_u1_n100 ) );
  NOR2_X1 u1_u11_u1_U72 (.A2( u1_u11_X_8 ) , .A1( u1_u11_u1_n177 ) , .ZN( u1_u11_u1_n99 ) );
  NOR2_X1 u1_u11_u1_U73 (.A2( u1_u11_X_12 ) , .ZN( u1_u11_u1_n102 ) , .A1( u1_u11_u1_n176 ) );
  NOR2_X1 u1_u11_u1_U74 (.A2( u1_u11_X_9 ) , .ZN( u1_u11_u1_n105 ) , .A1( u1_u11_u1_n168 ) );
  NAND2_X1 u1_u11_u1_U75 (.A1( u1_u11_X_10 ) , .ZN( u1_u11_u1_n160 ) , .A2( u1_u11_u1_n169 ) );
  NAND2_X1 u1_u11_u1_U76 (.A2( u1_u11_X_10 ) , .A1( u1_u11_X_11 ) , .ZN( u1_u11_u1_n152 ) );
  NAND2_X1 u1_u11_u1_U77 (.A1( u1_u11_X_11 ) , .ZN( u1_u11_u1_n128 ) , .A2( u1_u11_u1_n170 ) );
  AND2_X1 u1_u11_u1_U78 (.A2( u1_u11_X_7 ) , .A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n104 ) );
  AND2_X1 u1_u11_u1_U79 (.A1( u1_u11_X_8 ) , .ZN( u1_u11_u1_n103 ) , .A2( u1_u11_u1_n177 ) );
  AOI22_X1 u1_u11_u1_U8 (.B2( u1_u11_u1_n136 ) , .A2( u1_u11_u1_n137 ) , .ZN( u1_u11_u1_n143 ) , .A1( u1_u11_u1_n171 ) , .B1( u1_u11_u1_n173 ) );
  INV_X1 u1_u11_u1_U80 (.A( u1_u11_X_10 ) , .ZN( u1_u11_u1_n170 ) );
  INV_X1 u1_u11_u1_U81 (.A( u1_u11_X_9 ) , .ZN( u1_u11_u1_n176 ) );
  INV_X1 u1_u11_u1_U82 (.A( u1_u11_X_11 ) , .ZN( u1_u11_u1_n169 ) );
  INV_X1 u1_u11_u1_U83 (.A( u1_u11_X_12 ) , .ZN( u1_u11_u1_n168 ) );
  INV_X1 u1_u11_u1_U84 (.A( u1_u11_X_7 ) , .ZN( u1_u11_u1_n177 ) );
  NAND4_X1 u1_u11_u1_U85 (.ZN( u1_out11_18 ) , .A4( u1_u11_u1_n165 ) , .A3( u1_u11_u1_n166 ) , .A1( u1_u11_u1_n167 ) , .A2( u1_u11_u1_n186 ) );
  AOI22_X1 u1_u11_u1_U86 (.B2( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n147 ) , .A2( u1_u11_u1_n148 ) , .ZN( u1_u11_u1_n166 ) , .A1( u1_u11_u1_n172 ) );
  INV_X1 u1_u11_u1_U87 (.A( u1_u11_u1_n145 ) , .ZN( u1_u11_u1_n186 ) );
  NAND4_X1 u1_u11_u1_U88 (.ZN( u1_out11_2 ) , .A4( u1_u11_u1_n142 ) , .A3( u1_u11_u1_n143 ) , .A2( u1_u11_u1_n144 ) , .A1( u1_u11_u1_n179 ) );
  OAI21_X1 u1_u11_u1_U89 (.B2( u1_u11_u1_n132 ) , .ZN( u1_u11_u1_n144 ) , .A( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n180 ) );
  INV_X1 u1_u11_u1_U9 (.A( u1_u11_u1_n147 ) , .ZN( u1_u11_u1_n181 ) );
  INV_X1 u1_u11_u1_U90 (.A( u1_u11_u1_n130 ) , .ZN( u1_u11_u1_n179 ) );
  NAND4_X1 u1_u11_u1_U91 (.ZN( u1_out11_28 ) , .A4( u1_u11_u1_n124 ) , .A3( u1_u11_u1_n125 ) , .A2( u1_u11_u1_n126 ) , .A1( u1_u11_u1_n127 ) );
  OAI21_X1 u1_u11_u1_U92 (.ZN( u1_u11_u1_n127 ) , .B2( u1_u11_u1_n139 ) , .B1( u1_u11_u1_n175 ) , .A( u1_u11_u1_n183 ) );
  OAI21_X1 u1_u11_u1_U93 (.ZN( u1_u11_u1_n126 ) , .B2( u1_u11_u1_n140 ) , .A( u1_u11_u1_n146 ) , .B1( u1_u11_u1_n178 ) );
  OR4_X1 u1_u11_u1_U94 (.ZN( u1_out11_13 ) , .A4( u1_u11_u1_n108 ) , .A3( u1_u11_u1_n109 ) , .A2( u1_u11_u1_n110 ) , .A1( u1_u11_u1_n111 ) );
  AOI21_X1 u1_u11_u1_U95 (.ZN( u1_u11_u1_n111 ) , .A( u1_u11_u1_n128 ) , .B2( u1_u11_u1_n131 ) , .B1( u1_u11_u1_n135 ) );
  AOI21_X1 u1_u11_u1_U96 (.ZN( u1_u11_u1_n110 ) , .A( u1_u11_u1_n116 ) , .B1( u1_u11_u1_n152 ) , .B2( u1_u11_u1_n160 ) );
  NAND3_X1 u1_u11_u1_U97 (.A3( u1_u11_u1_n149 ) , .A2( u1_u11_u1_n150 ) , .A1( u1_u11_u1_n151 ) , .ZN( u1_u11_u1_n164 ) );
  NAND3_X1 u1_u11_u1_U98 (.A3( u1_u11_u1_n134 ) , .A2( u1_u11_u1_n135 ) , .ZN( u1_u11_u1_n136 ) , .A1( u1_u11_u1_n151 ) );
  NAND3_X1 u1_u11_u1_U99 (.A1( u1_u11_u1_n133 ) , .ZN( u1_u11_u1_n137 ) , .A2( u1_u11_u1_n154 ) , .A3( u1_u11_u1_n181 ) );
  OAI22_X1 u1_u11_u2_U10 (.ZN( u1_u11_u2_n109 ) , .A2( u1_u11_u2_n113 ) , .B2( u1_u11_u2_n133 ) , .B1( u1_u11_u2_n167 ) , .A1( u1_u11_u2_n168 ) );
  NAND3_X1 u1_u11_u2_U100 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n98 ) );
  OAI22_X1 u1_u11_u2_U11 (.B1( u1_u11_u2_n151 ) , .A2( u1_u11_u2_n152 ) , .A1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n160 ) , .B2( u1_u11_u2_n168 ) );
  NOR3_X1 u1_u11_u2_U12 (.A1( u1_u11_u2_n150 ) , .ZN( u1_u11_u2_n151 ) , .A3( u1_u11_u2_n175 ) , .A2( u1_u11_u2_n188 ) );
  AOI21_X1 u1_u11_u2_U13 (.ZN( u1_u11_u2_n144 ) , .B2( u1_u11_u2_n155 ) , .A( u1_u11_u2_n172 ) , .B1( u1_u11_u2_n185 ) );
  AOI21_X1 u1_u11_u2_U14 (.B2( u1_u11_u2_n143 ) , .ZN( u1_u11_u2_n145 ) , .B1( u1_u11_u2_n152 ) , .A( u1_u11_u2_n171 ) );
  AOI21_X1 u1_u11_u2_U15 (.B2( u1_u11_u2_n120 ) , .B1( u1_u11_u2_n121 ) , .ZN( u1_u11_u2_n126 ) , .A( u1_u11_u2_n167 ) );
  INV_X1 u1_u11_u2_U16 (.A( u1_u11_u2_n156 ) , .ZN( u1_u11_u2_n171 ) );
  INV_X1 u1_u11_u2_U17 (.A( u1_u11_u2_n120 ) , .ZN( u1_u11_u2_n188 ) );
  NAND2_X1 u1_u11_u2_U18 (.A2( u1_u11_u2_n122 ) , .ZN( u1_u11_u2_n150 ) , .A1( u1_u11_u2_n152 ) );
  INV_X1 u1_u11_u2_U19 (.A( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n170 ) );
  INV_X1 u1_u11_u2_U20 (.A( u1_u11_u2_n137 ) , .ZN( u1_u11_u2_n173 ) );
  NAND2_X1 u1_u11_u2_U21 (.A1( u1_u11_u2_n132 ) , .A2( u1_u11_u2_n139 ) , .ZN( u1_u11_u2_n157 ) );
  INV_X1 u1_u11_u2_U22 (.A( u1_u11_u2_n113 ) , .ZN( u1_u11_u2_n178 ) );
  INV_X1 u1_u11_u2_U23 (.A( u1_u11_u2_n139 ) , .ZN( u1_u11_u2_n175 ) );
  INV_X1 u1_u11_u2_U24 (.A( u1_u11_u2_n155 ) , .ZN( u1_u11_u2_n181 ) );
  INV_X1 u1_u11_u2_U25 (.A( u1_u11_u2_n119 ) , .ZN( u1_u11_u2_n177 ) );
  INV_X1 u1_u11_u2_U26 (.A( u1_u11_u2_n116 ) , .ZN( u1_u11_u2_n180 ) );
  INV_X1 u1_u11_u2_U27 (.A( u1_u11_u2_n131 ) , .ZN( u1_u11_u2_n179 ) );
  INV_X1 u1_u11_u2_U28 (.A( u1_u11_u2_n154 ) , .ZN( u1_u11_u2_n176 ) );
  NAND2_X1 u1_u11_u2_U29 (.A2( u1_u11_u2_n116 ) , .A1( u1_u11_u2_n117 ) , .ZN( u1_u11_u2_n118 ) );
  NOR2_X1 u1_u11_u2_U3 (.ZN( u1_u11_u2_n121 ) , .A2( u1_u11_u2_n177 ) , .A1( u1_u11_u2_n180 ) );
  INV_X1 u1_u11_u2_U30 (.A( u1_u11_u2_n132 ) , .ZN( u1_u11_u2_n182 ) );
  INV_X1 u1_u11_u2_U31 (.A( u1_u11_u2_n158 ) , .ZN( u1_u11_u2_n183 ) );
  OAI21_X1 u1_u11_u2_U32 (.A( u1_u11_u2_n156 ) , .B1( u1_u11_u2_n157 ) , .ZN( u1_u11_u2_n158 ) , .B2( u1_u11_u2_n179 ) );
  NOR2_X1 u1_u11_u2_U33 (.ZN( u1_u11_u2_n156 ) , .A1( u1_u11_u2_n166 ) , .A2( u1_u11_u2_n169 ) );
  NOR2_X1 u1_u11_u2_U34 (.A2( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n137 ) , .A1( u1_u11_u2_n140 ) );
  NOR2_X1 u1_u11_u2_U35 (.A2( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n153 ) , .A1( u1_u11_u2_n156 ) );
  AOI211_X1 u1_u11_u2_U36 (.ZN( u1_u11_u2_n130 ) , .C1( u1_u11_u2_n138 ) , .C2( u1_u11_u2_n179 ) , .B( u1_u11_u2_n96 ) , .A( u1_u11_u2_n97 ) );
  OAI22_X1 u1_u11_u2_U37 (.B1( u1_u11_u2_n133 ) , .A2( u1_u11_u2_n137 ) , .A1( u1_u11_u2_n152 ) , .B2( u1_u11_u2_n168 ) , .ZN( u1_u11_u2_n97 ) );
  OAI221_X1 u1_u11_u2_U38 (.B1( u1_u11_u2_n113 ) , .C1( u1_u11_u2_n132 ) , .A( u1_u11_u2_n149 ) , .B2( u1_u11_u2_n171 ) , .C2( u1_u11_u2_n172 ) , .ZN( u1_u11_u2_n96 ) );
  OAI221_X1 u1_u11_u2_U39 (.A( u1_u11_u2_n115 ) , .C2( u1_u11_u2_n123 ) , .B2( u1_u11_u2_n143 ) , .B1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n163 ) , .C1( u1_u11_u2_n168 ) );
  INV_X1 u1_u11_u2_U4 (.A( u1_u11_u2_n134 ) , .ZN( u1_u11_u2_n185 ) );
  OAI21_X1 u1_u11_u2_U40 (.A( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n115 ) , .B1( u1_u11_u2_n176 ) , .B2( u1_u11_u2_n178 ) );
  OAI221_X1 u1_u11_u2_U41 (.A( u1_u11_u2_n135 ) , .B2( u1_u11_u2_n136 ) , .B1( u1_u11_u2_n137 ) , .ZN( u1_u11_u2_n162 ) , .C2( u1_u11_u2_n167 ) , .C1( u1_u11_u2_n185 ) );
  AND3_X1 u1_u11_u2_U42 (.A3( u1_u11_u2_n131 ) , .A2( u1_u11_u2_n132 ) , .A1( u1_u11_u2_n133 ) , .ZN( u1_u11_u2_n136 ) );
  AOI22_X1 u1_u11_u2_U43 (.ZN( u1_u11_u2_n135 ) , .B1( u1_u11_u2_n140 ) , .A1( u1_u11_u2_n156 ) , .B2( u1_u11_u2_n180 ) , .A2( u1_u11_u2_n188 ) );
  AOI21_X1 u1_u11_u2_U44 (.ZN( u1_u11_u2_n149 ) , .B1( u1_u11_u2_n173 ) , .B2( u1_u11_u2_n188 ) , .A( u1_u11_u2_n95 ) );
  AND3_X1 u1_u11_u2_U45 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n156 ) , .ZN( u1_u11_u2_n95 ) );
  OAI21_X1 u1_u11_u2_U46 (.A( u1_u11_u2_n101 ) , .B2( u1_u11_u2_n121 ) , .B1( u1_u11_u2_n153 ) , .ZN( u1_u11_u2_n164 ) );
  NAND2_X1 u1_u11_u2_U47 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n155 ) );
  NAND2_X1 u1_u11_u2_U48 (.A2( u1_u11_u2_n105 ) , .A1( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n143 ) );
  NAND2_X1 u1_u11_u2_U49 (.A1( u1_u11_u2_n104 ) , .A2( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n152 ) );
  INV_X1 u1_u11_u2_U5 (.A( u1_u11_u2_n150 ) , .ZN( u1_u11_u2_n184 ) );
  NAND2_X1 u1_u11_u2_U50 (.A1( u1_u11_u2_n100 ) , .A2( u1_u11_u2_n105 ) , .ZN( u1_u11_u2_n132 ) );
  INV_X1 u1_u11_u2_U51 (.A( u1_u11_u2_n140 ) , .ZN( u1_u11_u2_n168 ) );
  INV_X1 u1_u11_u2_U52 (.A( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n167 ) );
  OAI21_X1 u1_u11_u2_U53 (.A( u1_u11_u2_n141 ) , .B2( u1_u11_u2_n142 ) , .ZN( u1_u11_u2_n146 ) , .B1( u1_u11_u2_n153 ) );
  OAI21_X1 u1_u11_u2_U54 (.A( u1_u11_u2_n140 ) , .ZN( u1_u11_u2_n141 ) , .B1( u1_u11_u2_n176 ) , .B2( u1_u11_u2_n177 ) );
  NOR3_X1 u1_u11_u2_U55 (.ZN( u1_u11_u2_n142 ) , .A3( u1_u11_u2_n175 ) , .A2( u1_u11_u2_n178 ) , .A1( u1_u11_u2_n181 ) );
  INV_X1 u1_u11_u2_U56 (.ZN( u1_u11_u2_n187 ) , .A( u1_u11_u2_n99 ) );
  OAI21_X1 u1_u11_u2_U57 (.B1( u1_u11_u2_n137 ) , .B2( u1_u11_u2_n143 ) , .A( u1_u11_u2_n98 ) , .ZN( u1_u11_u2_n99 ) );
  NAND2_X1 u1_u11_u2_U58 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n113 ) );
  NAND2_X1 u1_u11_u2_U59 (.A1( u1_u11_u2_n106 ) , .A2( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n131 ) );
  NOR4_X1 u1_u11_u2_U6 (.A4( u1_u11_u2_n124 ) , .A3( u1_u11_u2_n125 ) , .A2( u1_u11_u2_n126 ) , .A1( u1_u11_u2_n127 ) , .ZN( u1_u11_u2_n128 ) );
  NAND2_X1 u1_u11_u2_U60 (.A1( u1_u11_u2_n103 ) , .A2( u1_u11_u2_n107 ) , .ZN( u1_u11_u2_n139 ) );
  NAND2_X1 u1_u11_u2_U61 (.A1( u1_u11_u2_n103 ) , .A2( u1_u11_u2_n105 ) , .ZN( u1_u11_u2_n133 ) );
  NAND2_X1 u1_u11_u2_U62 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n103 ) , .ZN( u1_u11_u2_n154 ) );
  NAND2_X1 u1_u11_u2_U63 (.A2( u1_u11_u2_n103 ) , .A1( u1_u11_u2_n104 ) , .ZN( u1_u11_u2_n119 ) );
  NAND2_X1 u1_u11_u2_U64 (.A2( u1_u11_u2_n107 ) , .A1( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n123 ) );
  NAND2_X1 u1_u11_u2_U65 (.A1( u1_u11_u2_n104 ) , .A2( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n122 ) );
  INV_X1 u1_u11_u2_U66 (.A( u1_u11_u2_n114 ) , .ZN( u1_u11_u2_n172 ) );
  NAND2_X1 u1_u11_u2_U67 (.A2( u1_u11_u2_n100 ) , .A1( u1_u11_u2_n102 ) , .ZN( u1_u11_u2_n116 ) );
  NAND2_X1 u1_u11_u2_U68 (.A1( u1_u11_u2_n102 ) , .A2( u1_u11_u2_n108 ) , .ZN( u1_u11_u2_n120 ) );
  NAND2_X1 u1_u11_u2_U69 (.A2( u1_u11_u2_n105 ) , .A1( u1_u11_u2_n106 ) , .ZN( u1_u11_u2_n117 ) );
  AOI21_X1 u1_u11_u2_U7 (.ZN( u1_u11_u2_n124 ) , .B1( u1_u11_u2_n131 ) , .B2( u1_u11_u2_n143 ) , .A( u1_u11_u2_n172 ) );
  NOR2_X1 u1_u11_u2_U70 (.A2( u1_u11_X_16 ) , .ZN( u1_u11_u2_n140 ) , .A1( u1_u11_u2_n166 ) );
  NOR2_X1 u1_u11_u2_U71 (.A2( u1_u11_X_13 ) , .A1( u1_u11_X_14 ) , .ZN( u1_u11_u2_n100 ) );
  NOR2_X1 u1_u11_u2_U72 (.A2( u1_u11_X_16 ) , .A1( u1_u11_X_17 ) , .ZN( u1_u11_u2_n138 ) );
  NOR2_X1 u1_u11_u2_U73 (.A2( u1_u11_X_15 ) , .A1( u1_u11_X_18 ) , .ZN( u1_u11_u2_n104 ) );
  NOR2_X1 u1_u11_u2_U74 (.A2( u1_u11_X_14 ) , .ZN( u1_u11_u2_n103 ) , .A1( u1_u11_u2_n174 ) );
  NOR2_X1 u1_u11_u2_U75 (.A2( u1_u11_X_15 ) , .ZN( u1_u11_u2_n102 ) , .A1( u1_u11_u2_n165 ) );
  NOR2_X1 u1_u11_u2_U76 (.A2( u1_u11_X_17 ) , .ZN( u1_u11_u2_n114 ) , .A1( u1_u11_u2_n169 ) );
  AND2_X1 u1_u11_u2_U77 (.A1( u1_u11_X_15 ) , .ZN( u1_u11_u2_n105 ) , .A2( u1_u11_u2_n165 ) );
  AND2_X1 u1_u11_u2_U78 (.A2( u1_u11_X_15 ) , .A1( u1_u11_X_18 ) , .ZN( u1_u11_u2_n107 ) );
  AND2_X1 u1_u11_u2_U79 (.A1( u1_u11_X_14 ) , .ZN( u1_u11_u2_n106 ) , .A2( u1_u11_u2_n174 ) );
  AOI21_X1 u1_u11_u2_U8 (.B2( u1_u11_u2_n119 ) , .ZN( u1_u11_u2_n127 ) , .A( u1_u11_u2_n137 ) , .B1( u1_u11_u2_n155 ) );
  AND2_X1 u1_u11_u2_U80 (.A1( u1_u11_X_13 ) , .A2( u1_u11_X_14 ) , .ZN( u1_u11_u2_n108 ) );
  INV_X1 u1_u11_u2_U81 (.A( u1_u11_X_16 ) , .ZN( u1_u11_u2_n169 ) );
  INV_X1 u1_u11_u2_U82 (.A( u1_u11_X_17 ) , .ZN( u1_u11_u2_n166 ) );
  INV_X1 u1_u11_u2_U83 (.A( u1_u11_X_13 ) , .ZN( u1_u11_u2_n174 ) );
  INV_X1 u1_u11_u2_U84 (.A( u1_u11_X_18 ) , .ZN( u1_u11_u2_n165 ) );
  NAND4_X1 u1_u11_u2_U85 (.ZN( u1_out11_30 ) , .A4( u1_u11_u2_n147 ) , .A3( u1_u11_u2_n148 ) , .A2( u1_u11_u2_n149 ) , .A1( u1_u11_u2_n187 ) );
  NOR3_X1 u1_u11_u2_U86 (.A3( u1_u11_u2_n144 ) , .A2( u1_u11_u2_n145 ) , .A1( u1_u11_u2_n146 ) , .ZN( u1_u11_u2_n147 ) );
  AOI21_X1 u1_u11_u2_U87 (.B2( u1_u11_u2_n138 ) , .ZN( u1_u11_u2_n148 ) , .A( u1_u11_u2_n162 ) , .B1( u1_u11_u2_n182 ) );
  NAND4_X1 u1_u11_u2_U88 (.ZN( u1_out11_24 ) , .A4( u1_u11_u2_n111 ) , .A3( u1_u11_u2_n112 ) , .A1( u1_u11_u2_n130 ) , .A2( u1_u11_u2_n187 ) );
  AOI221_X1 u1_u11_u2_U89 (.A( u1_u11_u2_n109 ) , .B1( u1_u11_u2_n110 ) , .ZN( u1_u11_u2_n111 ) , .C1( u1_u11_u2_n134 ) , .C2( u1_u11_u2_n170 ) , .B2( u1_u11_u2_n173 ) );
  AOI21_X1 u1_u11_u2_U9 (.B2( u1_u11_u2_n123 ) , .ZN( u1_u11_u2_n125 ) , .A( u1_u11_u2_n171 ) , .B1( u1_u11_u2_n184 ) );
  AOI21_X1 u1_u11_u2_U90 (.ZN( u1_u11_u2_n112 ) , .B2( u1_u11_u2_n156 ) , .A( u1_u11_u2_n164 ) , .B1( u1_u11_u2_n181 ) );
  NAND4_X1 u1_u11_u2_U91 (.ZN( u1_out11_16 ) , .A4( u1_u11_u2_n128 ) , .A3( u1_u11_u2_n129 ) , .A1( u1_u11_u2_n130 ) , .A2( u1_u11_u2_n186 ) );
  AOI22_X1 u1_u11_u2_U92 (.A2( u1_u11_u2_n118 ) , .ZN( u1_u11_u2_n129 ) , .A1( u1_u11_u2_n140 ) , .B1( u1_u11_u2_n157 ) , .B2( u1_u11_u2_n170 ) );
  INV_X1 u1_u11_u2_U93 (.A( u1_u11_u2_n163 ) , .ZN( u1_u11_u2_n186 ) );
  OR4_X1 u1_u11_u2_U94 (.ZN( u1_out11_6 ) , .A4( u1_u11_u2_n161 ) , .A3( u1_u11_u2_n162 ) , .A2( u1_u11_u2_n163 ) , .A1( u1_u11_u2_n164 ) );
  OR3_X1 u1_u11_u2_U95 (.A2( u1_u11_u2_n159 ) , .A1( u1_u11_u2_n160 ) , .ZN( u1_u11_u2_n161 ) , .A3( u1_u11_u2_n183 ) );
  AOI21_X1 u1_u11_u2_U96 (.B2( u1_u11_u2_n154 ) , .B1( u1_u11_u2_n155 ) , .ZN( u1_u11_u2_n159 ) , .A( u1_u11_u2_n167 ) );
  NAND3_X1 u1_u11_u2_U97 (.A2( u1_u11_u2_n117 ) , .A1( u1_u11_u2_n122 ) , .A3( u1_u11_u2_n123 ) , .ZN( u1_u11_u2_n134 ) );
  NAND3_X1 u1_u11_u2_U98 (.ZN( u1_u11_u2_n110 ) , .A2( u1_u11_u2_n131 ) , .A3( u1_u11_u2_n139 ) , .A1( u1_u11_u2_n154 ) );
  NAND3_X1 u1_u11_u2_U99 (.A2( u1_u11_u2_n100 ) , .ZN( u1_u11_u2_n101 ) , .A1( u1_u11_u2_n104 ) , .A3( u1_u11_u2_n114 ) );
  OAI211_X1 u1_u11_u3_U10 (.B( u1_u11_u3_n106 ) , .ZN( u1_u11_u3_n119 ) , .C2( u1_u11_u3_n128 ) , .C1( u1_u11_u3_n167 ) , .A( u1_u11_u3_n181 ) );
  INV_X1 u1_u11_u3_U11 (.ZN( u1_u11_u3_n181 ) , .A( u1_u11_u3_n98 ) );
  AOI221_X1 u1_u11_u3_U12 (.C1( u1_u11_u3_n105 ) , .ZN( u1_u11_u3_n106 ) , .A( u1_u11_u3_n131 ) , .B2( u1_u11_u3_n132 ) , .C2( u1_u11_u3_n133 ) , .B1( u1_u11_u3_n169 ) );
  OAI22_X1 u1_u11_u3_U13 (.B1( u1_u11_u3_n113 ) , .A2( u1_u11_u3_n135 ) , .A1( u1_u11_u3_n150 ) , .B2( u1_u11_u3_n164 ) , .ZN( u1_u11_u3_n98 ) );
  AOI22_X1 u1_u11_u3_U14 (.B1( u1_u11_u3_n115 ) , .A2( u1_u11_u3_n116 ) , .ZN( u1_u11_u3_n123 ) , .B2( u1_u11_u3_n133 ) , .A1( u1_u11_u3_n169 ) );
  NAND2_X1 u1_u11_u3_U15 (.ZN( u1_u11_u3_n116 ) , .A2( u1_u11_u3_n151 ) , .A1( u1_u11_u3_n182 ) );
  NOR2_X1 u1_u11_u3_U16 (.ZN( u1_u11_u3_n126 ) , .A2( u1_u11_u3_n150 ) , .A1( u1_u11_u3_n164 ) );
  AOI21_X1 u1_u11_u3_U17 (.ZN( u1_u11_u3_n112 ) , .B2( u1_u11_u3_n146 ) , .B1( u1_u11_u3_n155 ) , .A( u1_u11_u3_n167 ) );
  NAND2_X1 u1_u11_u3_U18 (.A1( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n142 ) , .A2( u1_u11_u3_n164 ) );
  NAND2_X1 u1_u11_u3_U19 (.ZN( u1_u11_u3_n132 ) , .A2( u1_u11_u3_n152 ) , .A1( u1_u11_u3_n156 ) );
  INV_X1 u1_u11_u3_U20 (.A( u1_u11_u3_n133 ) , .ZN( u1_u11_u3_n165 ) );
  AND2_X1 u1_u11_u3_U21 (.A2( u1_u11_u3_n113 ) , .A1( u1_u11_u3_n114 ) , .ZN( u1_u11_u3_n151 ) );
  INV_X1 u1_u11_u3_U22 (.A( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n170 ) );
  NAND2_X1 u1_u11_u3_U23 (.A1( u1_u11_u3_n107 ) , .A2( u1_u11_u3_n108 ) , .ZN( u1_u11_u3_n140 ) );
  NAND2_X1 u1_u11_u3_U24 (.ZN( u1_u11_u3_n117 ) , .A1( u1_u11_u3_n124 ) , .A2( u1_u11_u3_n148 ) );
  NAND2_X1 u1_u11_u3_U25 (.ZN( u1_u11_u3_n143 ) , .A1( u1_u11_u3_n165 ) , .A2( u1_u11_u3_n167 ) );
  INV_X1 u1_u11_u3_U26 (.A( u1_u11_u3_n130 ) , .ZN( u1_u11_u3_n177 ) );
  INV_X1 u1_u11_u3_U27 (.A( u1_u11_u3_n128 ) , .ZN( u1_u11_u3_n176 ) );
  NAND2_X1 u1_u11_u3_U28 (.ZN( u1_u11_u3_n105 ) , .A2( u1_u11_u3_n130 ) , .A1( u1_u11_u3_n155 ) );
  INV_X1 u1_u11_u3_U29 (.A( u1_u11_u3_n155 ) , .ZN( u1_u11_u3_n174 ) );
  INV_X1 u1_u11_u3_U3 (.A( u1_u11_u3_n140 ) , .ZN( u1_u11_u3_n182 ) );
  INV_X1 u1_u11_u3_U30 (.A( u1_u11_u3_n139 ) , .ZN( u1_u11_u3_n185 ) );
  NOR2_X1 u1_u11_u3_U31 (.ZN( u1_u11_u3_n135 ) , .A2( u1_u11_u3_n141 ) , .A1( u1_u11_u3_n169 ) );
  OAI222_X1 u1_u11_u3_U32 (.C2( u1_u11_u3_n107 ) , .A2( u1_u11_u3_n108 ) , .B1( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n138 ) , .B2( u1_u11_u3_n146 ) , .C1( u1_u11_u3_n154 ) , .A1( u1_u11_u3_n164 ) );
  NOR4_X1 u1_u11_u3_U33 (.A4( u1_u11_u3_n157 ) , .A3( u1_u11_u3_n158 ) , .A2( u1_u11_u3_n159 ) , .A1( u1_u11_u3_n160 ) , .ZN( u1_u11_u3_n161 ) );
  AOI21_X1 u1_u11_u3_U34 (.B2( u1_u11_u3_n152 ) , .B1( u1_u11_u3_n153 ) , .ZN( u1_u11_u3_n158 ) , .A( u1_u11_u3_n164 ) );
  AOI21_X1 u1_u11_u3_U35 (.A( u1_u11_u3_n154 ) , .B2( u1_u11_u3_n155 ) , .B1( u1_u11_u3_n156 ) , .ZN( u1_u11_u3_n157 ) );
  AOI21_X1 u1_u11_u3_U36 (.A( u1_u11_u3_n149 ) , .B2( u1_u11_u3_n150 ) , .B1( u1_u11_u3_n151 ) , .ZN( u1_u11_u3_n159 ) );
  AOI211_X1 u1_u11_u3_U37 (.ZN( u1_u11_u3_n109 ) , .A( u1_u11_u3_n119 ) , .C2( u1_u11_u3_n129 ) , .B( u1_u11_u3_n138 ) , .C1( u1_u11_u3_n141 ) );
  AOI211_X1 u1_u11_u3_U38 (.B( u1_u11_u3_n119 ) , .A( u1_u11_u3_n120 ) , .C2( u1_u11_u3_n121 ) , .ZN( u1_u11_u3_n122 ) , .C1( u1_u11_u3_n179 ) );
  INV_X1 u1_u11_u3_U39 (.A( u1_u11_u3_n156 ) , .ZN( u1_u11_u3_n179 ) );
  INV_X1 u1_u11_u3_U4 (.A( u1_u11_u3_n129 ) , .ZN( u1_u11_u3_n183 ) );
  OAI22_X1 u1_u11_u3_U40 (.B1( u1_u11_u3_n118 ) , .ZN( u1_u11_u3_n120 ) , .A1( u1_u11_u3_n135 ) , .B2( u1_u11_u3_n154 ) , .A2( u1_u11_u3_n178 ) );
  AND3_X1 u1_u11_u3_U41 (.ZN( u1_u11_u3_n118 ) , .A2( u1_u11_u3_n124 ) , .A1( u1_u11_u3_n144 ) , .A3( u1_u11_u3_n152 ) );
  INV_X1 u1_u11_u3_U42 (.A( u1_u11_u3_n121 ) , .ZN( u1_u11_u3_n164 ) );
  NAND2_X1 u1_u11_u3_U43 (.ZN( u1_u11_u3_n133 ) , .A1( u1_u11_u3_n154 ) , .A2( u1_u11_u3_n164 ) );
  NOR2_X1 u1_u11_u3_U44 (.A1( u1_u11_u3_n113 ) , .ZN( u1_u11_u3_n131 ) , .A2( u1_u11_u3_n154 ) );
  NAND2_X1 u1_u11_u3_U45 (.A1( u1_u11_u3_n103 ) , .ZN( u1_u11_u3_n150 ) , .A2( u1_u11_u3_n99 ) );
  NAND2_X1 u1_u11_u3_U46 (.A2( u1_u11_u3_n102 ) , .ZN( u1_u11_u3_n155 ) , .A1( u1_u11_u3_n97 ) );
  OAI211_X1 u1_u11_u3_U47 (.B( u1_u11_u3_n127 ) , .ZN( u1_u11_u3_n139 ) , .C1( u1_u11_u3_n150 ) , .C2( u1_u11_u3_n154 ) , .A( u1_u11_u3_n184 ) );
  INV_X1 u1_u11_u3_U48 (.A( u1_u11_u3_n125 ) , .ZN( u1_u11_u3_n184 ) );
  AOI221_X1 u1_u11_u3_U49 (.A( u1_u11_u3_n126 ) , .ZN( u1_u11_u3_n127 ) , .C2( u1_u11_u3_n132 ) , .C1( u1_u11_u3_n169 ) , .B2( u1_u11_u3_n170 ) , .B1( u1_u11_u3_n174 ) );
  INV_X1 u1_u11_u3_U5 (.A( u1_u11_u3_n117 ) , .ZN( u1_u11_u3_n178 ) );
  OAI22_X1 u1_u11_u3_U50 (.A1( u1_u11_u3_n124 ) , .ZN( u1_u11_u3_n125 ) , .B2( u1_u11_u3_n145 ) , .A2( u1_u11_u3_n165 ) , .B1( u1_u11_u3_n167 ) );
  INV_X1 u1_u11_u3_U51 (.A( u1_u11_u3_n141 ) , .ZN( u1_u11_u3_n167 ) );
  AOI21_X1 u1_u11_u3_U52 (.B2( u1_u11_u3_n114 ) , .B1( u1_u11_u3_n146 ) , .A( u1_u11_u3_n154 ) , .ZN( u1_u11_u3_n94 ) );
  AOI21_X1 u1_u11_u3_U53 (.ZN( u1_u11_u3_n110 ) , .B2( u1_u11_u3_n142 ) , .B1( u1_u11_u3_n186 ) , .A( u1_u11_u3_n95 ) );
  INV_X1 u1_u11_u3_U54 (.A( u1_u11_u3_n145 ) , .ZN( u1_u11_u3_n186 ) );
  AOI21_X1 u1_u11_u3_U55 (.B1( u1_u11_u3_n124 ) , .A( u1_u11_u3_n149 ) , .B2( u1_u11_u3_n155 ) , .ZN( u1_u11_u3_n95 ) );
  INV_X1 u1_u11_u3_U56 (.A( u1_u11_u3_n149 ) , .ZN( u1_u11_u3_n169 ) );
  NAND2_X1 u1_u11_u3_U57 (.ZN( u1_u11_u3_n124 ) , .A1( u1_u11_u3_n96 ) , .A2( u1_u11_u3_n97 ) );
  NAND2_X1 u1_u11_u3_U58 (.A2( u1_u11_u3_n100 ) , .ZN( u1_u11_u3_n146 ) , .A1( u1_u11_u3_n96 ) );
  NAND2_X1 u1_u11_u3_U59 (.A1( u1_u11_u3_n101 ) , .ZN( u1_u11_u3_n145 ) , .A2( u1_u11_u3_n99 ) );
  AOI221_X1 u1_u11_u3_U6 (.A( u1_u11_u3_n131 ) , .C2( u1_u11_u3_n132 ) , .C1( u1_u11_u3_n133 ) , .ZN( u1_u11_u3_n134 ) , .B1( u1_u11_u3_n143 ) , .B2( u1_u11_u3_n177 ) );
  NAND2_X1 u1_u11_u3_U60 (.A1( u1_u11_u3_n100 ) , .ZN( u1_u11_u3_n156 ) , .A2( u1_u11_u3_n99 ) );
  NAND2_X1 u1_u11_u3_U61 (.A2( u1_u11_u3_n101 ) , .A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n148 ) );
  NAND2_X1 u1_u11_u3_U62 (.A1( u1_u11_u3_n100 ) , .A2( u1_u11_u3_n102 ) , .ZN( u1_u11_u3_n128 ) );
  NAND2_X1 u1_u11_u3_U63 (.A2( u1_u11_u3_n101 ) , .A1( u1_u11_u3_n102 ) , .ZN( u1_u11_u3_n152 ) );
  NAND2_X1 u1_u11_u3_U64 (.A2( u1_u11_u3_n101 ) , .ZN( u1_u11_u3_n114 ) , .A1( u1_u11_u3_n96 ) );
  NAND2_X1 u1_u11_u3_U65 (.ZN( u1_u11_u3_n107 ) , .A1( u1_u11_u3_n97 ) , .A2( u1_u11_u3_n99 ) );
  NAND2_X1 u1_u11_u3_U66 (.A2( u1_u11_u3_n100 ) , .A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n113 ) );
  NAND2_X1 u1_u11_u3_U67 (.A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n153 ) , .A2( u1_u11_u3_n97 ) );
  NAND2_X1 u1_u11_u3_U68 (.A2( u1_u11_u3_n103 ) , .A1( u1_u11_u3_n104 ) , .ZN( u1_u11_u3_n130 ) );
  NAND2_X1 u1_u11_u3_U69 (.A2( u1_u11_u3_n103 ) , .ZN( u1_u11_u3_n144 ) , .A1( u1_u11_u3_n96 ) );
  OAI22_X1 u1_u11_u3_U7 (.B2( u1_u11_u3_n147 ) , .A2( u1_u11_u3_n148 ) , .ZN( u1_u11_u3_n160 ) , .B1( u1_u11_u3_n165 ) , .A1( u1_u11_u3_n168 ) );
  NAND2_X1 u1_u11_u3_U70 (.A1( u1_u11_u3_n102 ) , .A2( u1_u11_u3_n103 ) , .ZN( u1_u11_u3_n108 ) );
  NOR2_X1 u1_u11_u3_U71 (.A2( u1_u11_X_19 ) , .A1( u1_u11_X_20 ) , .ZN( u1_u11_u3_n99 ) );
  NOR2_X1 u1_u11_u3_U72 (.A2( u1_u11_X_21 ) , .A1( u1_u11_X_24 ) , .ZN( u1_u11_u3_n103 ) );
  NOR2_X1 u1_u11_u3_U73 (.A2( u1_u11_X_24 ) , .A1( u1_u11_u3_n171 ) , .ZN( u1_u11_u3_n97 ) );
  NOR2_X1 u1_u11_u3_U74 (.A2( u1_u11_X_23 ) , .ZN( u1_u11_u3_n141 ) , .A1( u1_u11_u3_n166 ) );
  NOR2_X1 u1_u11_u3_U75 (.A2( u1_u11_X_19 ) , .A1( u1_u11_u3_n172 ) , .ZN( u1_u11_u3_n96 ) );
  NAND2_X1 u1_u11_u3_U76 (.A1( u1_u11_X_22 ) , .A2( u1_u11_X_23 ) , .ZN( u1_u11_u3_n154 ) );
  NAND2_X1 u1_u11_u3_U77 (.A1( u1_u11_X_23 ) , .ZN( u1_u11_u3_n149 ) , .A2( u1_u11_u3_n166 ) );
  NOR2_X1 u1_u11_u3_U78 (.A2( u1_u11_X_22 ) , .A1( u1_u11_X_23 ) , .ZN( u1_u11_u3_n121 ) );
  AND2_X1 u1_u11_u3_U79 (.A1( u1_u11_X_24 ) , .ZN( u1_u11_u3_n101 ) , .A2( u1_u11_u3_n171 ) );
  AND3_X1 u1_u11_u3_U8 (.A3( u1_u11_u3_n144 ) , .A2( u1_u11_u3_n145 ) , .A1( u1_u11_u3_n146 ) , .ZN( u1_u11_u3_n147 ) );
  AND2_X1 u1_u11_u3_U80 (.A1( u1_u11_X_19 ) , .ZN( u1_u11_u3_n102 ) , .A2( u1_u11_u3_n172 ) );
  AND2_X1 u1_u11_u3_U81 (.A1( u1_u11_X_21 ) , .A2( u1_u11_X_24 ) , .ZN( u1_u11_u3_n100 ) );
  AND2_X1 u1_u11_u3_U82 (.A2( u1_u11_X_19 ) , .A1( u1_u11_X_20 ) , .ZN( u1_u11_u3_n104 ) );
  INV_X1 u1_u11_u3_U83 (.A( u1_u11_X_22 ) , .ZN( u1_u11_u3_n166 ) );
  INV_X1 u1_u11_u3_U84 (.A( u1_u11_X_21 ) , .ZN( u1_u11_u3_n171 ) );
  INV_X1 u1_u11_u3_U85 (.A( u1_u11_X_20 ) , .ZN( u1_u11_u3_n172 ) );
  NAND4_X1 u1_u11_u3_U86 (.ZN( u1_out11_26 ) , .A4( u1_u11_u3_n109 ) , .A3( u1_u11_u3_n110 ) , .A2( u1_u11_u3_n111 ) , .A1( u1_u11_u3_n173 ) );
  INV_X1 u1_u11_u3_U87 (.ZN( u1_u11_u3_n173 ) , .A( u1_u11_u3_n94 ) );
  OAI21_X1 u1_u11_u3_U88 (.ZN( u1_u11_u3_n111 ) , .B2( u1_u11_u3_n117 ) , .A( u1_u11_u3_n133 ) , .B1( u1_u11_u3_n176 ) );
  NAND4_X1 u1_u11_u3_U89 (.ZN( u1_out11_20 ) , .A4( u1_u11_u3_n122 ) , .A3( u1_u11_u3_n123 ) , .A1( u1_u11_u3_n175 ) , .A2( u1_u11_u3_n180 ) );
  INV_X1 u1_u11_u3_U9 (.A( u1_u11_u3_n143 ) , .ZN( u1_u11_u3_n168 ) );
  INV_X1 u1_u11_u3_U90 (.A( u1_u11_u3_n126 ) , .ZN( u1_u11_u3_n180 ) );
  INV_X1 u1_u11_u3_U91 (.A( u1_u11_u3_n112 ) , .ZN( u1_u11_u3_n175 ) );
  OAI222_X1 u1_u11_u3_U92 (.C1( u1_u11_u3_n128 ) , .ZN( u1_u11_u3_n137 ) , .B1( u1_u11_u3_n148 ) , .A2( u1_u11_u3_n150 ) , .B2( u1_u11_u3_n154 ) , .C2( u1_u11_u3_n164 ) , .A1( u1_u11_u3_n167 ) );
  NAND4_X1 u1_u11_u3_U93 (.ZN( u1_out11_1 ) , .A4( u1_u11_u3_n161 ) , .A3( u1_u11_u3_n162 ) , .A2( u1_u11_u3_n163 ) , .A1( u1_u11_u3_n185 ) );
  NAND2_X1 u1_u11_u3_U94 (.ZN( u1_u11_u3_n163 ) , .A2( u1_u11_u3_n170 ) , .A1( u1_u11_u3_n176 ) );
  AOI22_X1 u1_u11_u3_U95 (.B2( u1_u11_u3_n140 ) , .B1( u1_u11_u3_n141 ) , .A2( u1_u11_u3_n142 ) , .ZN( u1_u11_u3_n162 ) , .A1( u1_u11_u3_n177 ) );
  OR4_X1 u1_u11_u3_U96 (.ZN( u1_out11_10 ) , .A4( u1_u11_u3_n136 ) , .A3( u1_u11_u3_n137 ) , .A1( u1_u11_u3_n138 ) , .A2( u1_u11_u3_n139 ) );
  OAI221_X1 u1_u11_u3_U97 (.A( u1_u11_u3_n134 ) , .B2( u1_u11_u3_n135 ) , .ZN( u1_u11_u3_n136 ) , .C1( u1_u11_u3_n149 ) , .B1( u1_u11_u3_n151 ) , .C2( u1_u11_u3_n183 ) );
  NAND3_X1 u1_u11_u3_U98 (.A1( u1_u11_u3_n114 ) , .ZN( u1_u11_u3_n115 ) , .A2( u1_u11_u3_n145 ) , .A3( u1_u11_u3_n153 ) );
  NAND3_X1 u1_u11_u3_U99 (.ZN( u1_u11_u3_n129 ) , .A2( u1_u11_u3_n144 ) , .A1( u1_u11_u3_n153 ) , .A3( u1_u11_u3_n182 ) );
  OAI22_X1 u1_u11_u4_U10 (.B2( u1_u11_u4_n135 ) , .ZN( u1_u11_u4_n137 ) , .B1( u1_u11_u4_n153 ) , .A1( u1_u11_u4_n155 ) , .A2( u1_u11_u4_n171 ) );
  AND3_X1 u1_u11_u4_U11 (.A2( u1_u11_u4_n134 ) , .ZN( u1_u11_u4_n135 ) , .A3( u1_u11_u4_n145 ) , .A1( u1_u11_u4_n157 ) );
  NAND2_X1 u1_u11_u4_U12 (.ZN( u1_u11_u4_n132 ) , .A2( u1_u11_u4_n170 ) , .A1( u1_u11_u4_n173 ) );
  AOI21_X1 u1_u11_u4_U13 (.B2( u1_u11_u4_n160 ) , .B1( u1_u11_u4_n161 ) , .ZN( u1_u11_u4_n162 ) , .A( u1_u11_u4_n170 ) );
  AOI21_X1 u1_u11_u4_U14 (.ZN( u1_u11_u4_n107 ) , .B2( u1_u11_u4_n143 ) , .A( u1_u11_u4_n174 ) , .B1( u1_u11_u4_n184 ) );
  AOI21_X1 u1_u11_u4_U15 (.B2( u1_u11_u4_n158 ) , .B1( u1_u11_u4_n159 ) , .ZN( u1_u11_u4_n163 ) , .A( u1_u11_u4_n174 ) );
  AOI21_X1 u1_u11_u4_U16 (.A( u1_u11_u4_n153 ) , .B2( u1_u11_u4_n154 ) , .B1( u1_u11_u4_n155 ) , .ZN( u1_u11_u4_n165 ) );
  AOI21_X1 u1_u11_u4_U17 (.A( u1_u11_u4_n156 ) , .B2( u1_u11_u4_n157 ) , .ZN( u1_u11_u4_n164 ) , .B1( u1_u11_u4_n184 ) );
  INV_X1 u1_u11_u4_U18 (.A( u1_u11_u4_n138 ) , .ZN( u1_u11_u4_n170 ) );
  AND2_X1 u1_u11_u4_U19 (.A2( u1_u11_u4_n120 ) , .ZN( u1_u11_u4_n155 ) , .A1( u1_u11_u4_n160 ) );
  INV_X1 u1_u11_u4_U20 (.A( u1_u11_u4_n156 ) , .ZN( u1_u11_u4_n175 ) );
  NAND2_X1 u1_u11_u4_U21 (.A2( u1_u11_u4_n118 ) , .ZN( u1_u11_u4_n131 ) , .A1( u1_u11_u4_n147 ) );
  NAND2_X1 u1_u11_u4_U22 (.A1( u1_u11_u4_n119 ) , .A2( u1_u11_u4_n120 ) , .ZN( u1_u11_u4_n130 ) );
  NAND2_X1 u1_u11_u4_U23 (.ZN( u1_u11_u4_n117 ) , .A2( u1_u11_u4_n118 ) , .A1( u1_u11_u4_n148 ) );
  NAND2_X1 u1_u11_u4_U24 (.ZN( u1_u11_u4_n129 ) , .A1( u1_u11_u4_n134 ) , .A2( u1_u11_u4_n148 ) );
  AND3_X1 u1_u11_u4_U25 (.A1( u1_u11_u4_n119 ) , .A2( u1_u11_u4_n143 ) , .A3( u1_u11_u4_n154 ) , .ZN( u1_u11_u4_n161 ) );
  AND2_X1 u1_u11_u4_U26 (.A1( u1_u11_u4_n145 ) , .A2( u1_u11_u4_n147 ) , .ZN( u1_u11_u4_n159 ) );
  OR3_X1 u1_u11_u4_U27 (.A3( u1_u11_u4_n114 ) , .A2( u1_u11_u4_n115 ) , .A1( u1_u11_u4_n116 ) , .ZN( u1_u11_u4_n136 ) );
  AOI21_X1 u1_u11_u4_U28 (.A( u1_u11_u4_n113 ) , .ZN( u1_u11_u4_n116 ) , .B2( u1_u11_u4_n173 ) , .B1( u1_u11_u4_n174 ) );
  AOI21_X1 u1_u11_u4_U29 (.ZN( u1_u11_u4_n115 ) , .B2( u1_u11_u4_n145 ) , .B1( u1_u11_u4_n146 ) , .A( u1_u11_u4_n156 ) );
  NOR2_X1 u1_u11_u4_U3 (.ZN( u1_u11_u4_n121 ) , .A1( u1_u11_u4_n181 ) , .A2( u1_u11_u4_n182 ) );
  OAI22_X1 u1_u11_u4_U30 (.ZN( u1_u11_u4_n114 ) , .A2( u1_u11_u4_n121 ) , .B1( u1_u11_u4_n160 ) , .B2( u1_u11_u4_n170 ) , .A1( u1_u11_u4_n171 ) );
  INV_X1 u1_u11_u4_U31 (.A( u1_u11_u4_n158 ) , .ZN( u1_u11_u4_n182 ) );
  INV_X1 u1_u11_u4_U32 (.ZN( u1_u11_u4_n181 ) , .A( u1_u11_u4_n96 ) );
  INV_X1 u1_u11_u4_U33 (.A( u1_u11_u4_n144 ) , .ZN( u1_u11_u4_n179 ) );
  INV_X1 u1_u11_u4_U34 (.A( u1_u11_u4_n157 ) , .ZN( u1_u11_u4_n178 ) );
  NAND2_X1 u1_u11_u4_U35 (.A2( u1_u11_u4_n154 ) , .A1( u1_u11_u4_n96 ) , .ZN( u1_u11_u4_n97 ) );
  INV_X1 u1_u11_u4_U36 (.ZN( u1_u11_u4_n186 ) , .A( u1_u11_u4_n95 ) );
  OAI221_X1 u1_u11_u4_U37 (.C1( u1_u11_u4_n134 ) , .B1( u1_u11_u4_n158 ) , .B2( u1_u11_u4_n171 ) , .C2( u1_u11_u4_n173 ) , .A( u1_u11_u4_n94 ) , .ZN( u1_u11_u4_n95 ) );
  AOI222_X1 u1_u11_u4_U38 (.B2( u1_u11_u4_n132 ) , .A1( u1_u11_u4_n138 ) , .C2( u1_u11_u4_n175 ) , .A2( u1_u11_u4_n179 ) , .C1( u1_u11_u4_n181 ) , .B1( u1_u11_u4_n185 ) , .ZN( u1_u11_u4_n94 ) );
  INV_X1 u1_u11_u4_U39 (.A( u1_u11_u4_n113 ) , .ZN( u1_u11_u4_n185 ) );
  INV_X1 u1_u11_u4_U4 (.A( u1_u11_u4_n117 ) , .ZN( u1_u11_u4_n184 ) );
  INV_X1 u1_u11_u4_U40 (.A( u1_u11_u4_n143 ) , .ZN( u1_u11_u4_n183 ) );
  NOR2_X1 u1_u11_u4_U41 (.ZN( u1_u11_u4_n138 ) , .A1( u1_u11_u4_n168 ) , .A2( u1_u11_u4_n169 ) );
  NOR2_X1 u1_u11_u4_U42 (.A1( u1_u11_u4_n150 ) , .A2( u1_u11_u4_n152 ) , .ZN( u1_u11_u4_n153 ) );
  NOR2_X1 u1_u11_u4_U43 (.A2( u1_u11_u4_n128 ) , .A1( u1_u11_u4_n138 ) , .ZN( u1_u11_u4_n156 ) );
  AOI22_X1 u1_u11_u4_U44 (.B2( u1_u11_u4_n122 ) , .A1( u1_u11_u4_n123 ) , .ZN( u1_u11_u4_n124 ) , .B1( u1_u11_u4_n128 ) , .A2( u1_u11_u4_n172 ) );
  INV_X1 u1_u11_u4_U45 (.A( u1_u11_u4_n153 ) , .ZN( u1_u11_u4_n172 ) );
  NAND2_X1 u1_u11_u4_U46 (.A2( u1_u11_u4_n120 ) , .ZN( u1_u11_u4_n123 ) , .A1( u1_u11_u4_n161 ) );
  AOI22_X1 u1_u11_u4_U47 (.B2( u1_u11_u4_n132 ) , .A2( u1_u11_u4_n133 ) , .ZN( u1_u11_u4_n140 ) , .A1( u1_u11_u4_n150 ) , .B1( u1_u11_u4_n179 ) );
  NAND2_X1 u1_u11_u4_U48 (.ZN( u1_u11_u4_n133 ) , .A2( u1_u11_u4_n146 ) , .A1( u1_u11_u4_n154 ) );
  NAND2_X1 u1_u11_u4_U49 (.A1( u1_u11_u4_n103 ) , .ZN( u1_u11_u4_n154 ) , .A2( u1_u11_u4_n98 ) );
  NOR4_X1 u1_u11_u4_U5 (.A4( u1_u11_u4_n106 ) , .A3( u1_u11_u4_n107 ) , .A2( u1_u11_u4_n108 ) , .A1( u1_u11_u4_n109 ) , .ZN( u1_u11_u4_n110 ) );
  NAND2_X1 u1_u11_u4_U50 (.A1( u1_u11_u4_n101 ) , .ZN( u1_u11_u4_n158 ) , .A2( u1_u11_u4_n99 ) );
  AOI21_X1 u1_u11_u4_U51 (.ZN( u1_u11_u4_n127 ) , .A( u1_u11_u4_n136 ) , .B2( u1_u11_u4_n150 ) , .B1( u1_u11_u4_n180 ) );
  INV_X1 u1_u11_u4_U52 (.A( u1_u11_u4_n160 ) , .ZN( u1_u11_u4_n180 ) );
  NAND2_X1 u1_u11_u4_U53 (.A2( u1_u11_u4_n104 ) , .A1( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n146 ) );
  NAND2_X1 u1_u11_u4_U54 (.A2( u1_u11_u4_n101 ) , .A1( u1_u11_u4_n102 ) , .ZN( u1_u11_u4_n160 ) );
  NAND2_X1 u1_u11_u4_U55 (.ZN( u1_u11_u4_n134 ) , .A1( u1_u11_u4_n98 ) , .A2( u1_u11_u4_n99 ) );
  NAND2_X1 u1_u11_u4_U56 (.A1( u1_u11_u4_n103 ) , .A2( u1_u11_u4_n104 ) , .ZN( u1_u11_u4_n143 ) );
  NAND2_X1 u1_u11_u4_U57 (.A2( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n145 ) , .A1( u1_u11_u4_n98 ) );
  NAND2_X1 u1_u11_u4_U58 (.A1( u1_u11_u4_n100 ) , .A2( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n120 ) );
  NAND2_X1 u1_u11_u4_U59 (.A1( u1_u11_u4_n102 ) , .A2( u1_u11_u4_n104 ) , .ZN( u1_u11_u4_n148 ) );
  AOI21_X1 u1_u11_u4_U6 (.ZN( u1_u11_u4_n106 ) , .B2( u1_u11_u4_n146 ) , .B1( u1_u11_u4_n158 ) , .A( u1_u11_u4_n170 ) );
  NAND2_X1 u1_u11_u4_U60 (.A2( u1_u11_u4_n100 ) , .A1( u1_u11_u4_n103 ) , .ZN( u1_u11_u4_n157 ) );
  INV_X1 u1_u11_u4_U61 (.A( u1_u11_u4_n150 ) , .ZN( u1_u11_u4_n173 ) );
  INV_X1 u1_u11_u4_U62 (.A( u1_u11_u4_n152 ) , .ZN( u1_u11_u4_n171 ) );
  NAND2_X1 u1_u11_u4_U63 (.A1( u1_u11_u4_n100 ) , .ZN( u1_u11_u4_n118 ) , .A2( u1_u11_u4_n99 ) );
  NAND2_X1 u1_u11_u4_U64 (.A2( u1_u11_u4_n100 ) , .A1( u1_u11_u4_n102 ) , .ZN( u1_u11_u4_n144 ) );
  NAND2_X1 u1_u11_u4_U65 (.A2( u1_u11_u4_n101 ) , .A1( u1_u11_u4_n105 ) , .ZN( u1_u11_u4_n96 ) );
  INV_X1 u1_u11_u4_U66 (.A( u1_u11_u4_n128 ) , .ZN( u1_u11_u4_n174 ) );
  NAND2_X1 u1_u11_u4_U67 (.A2( u1_u11_u4_n102 ) , .ZN( u1_u11_u4_n119 ) , .A1( u1_u11_u4_n98 ) );
  NAND2_X1 u1_u11_u4_U68 (.A2( u1_u11_u4_n101 ) , .A1( u1_u11_u4_n103 ) , .ZN( u1_u11_u4_n147 ) );
  NAND2_X1 u1_u11_u4_U69 (.A2( u1_u11_u4_n104 ) , .ZN( u1_u11_u4_n113 ) , .A1( u1_u11_u4_n99 ) );
  AOI21_X1 u1_u11_u4_U7 (.ZN( u1_u11_u4_n108 ) , .B2( u1_u11_u4_n134 ) , .B1( u1_u11_u4_n155 ) , .A( u1_u11_u4_n156 ) );
  NOR2_X1 u1_u11_u4_U70 (.A2( u1_u11_X_28 ) , .ZN( u1_u11_u4_n150 ) , .A1( u1_u11_u4_n168 ) );
  NOR2_X1 u1_u11_u4_U71 (.A2( u1_u11_X_29 ) , .ZN( u1_u11_u4_n152 ) , .A1( u1_u11_u4_n169 ) );
  NOR2_X1 u1_u11_u4_U72 (.A2( u1_u11_X_26 ) , .ZN( u1_u11_u4_n100 ) , .A1( u1_u11_u4_n177 ) );
  NOR2_X1 u1_u11_u4_U73 (.A2( u1_u11_X_30 ) , .ZN( u1_u11_u4_n105 ) , .A1( u1_u11_u4_n176 ) );
  NOR2_X1 u1_u11_u4_U74 (.A2( u1_u11_X_28 ) , .A1( u1_u11_X_29 ) , .ZN( u1_u11_u4_n128 ) );
  NOR2_X1 u1_u11_u4_U75 (.A2( u1_u11_X_25 ) , .A1( u1_u11_X_26 ) , .ZN( u1_u11_u4_n98 ) );
  NOR2_X1 u1_u11_u4_U76 (.A2( u1_u11_X_27 ) , .A1( u1_u11_X_30 ) , .ZN( u1_u11_u4_n102 ) );
  AND2_X1 u1_u11_u4_U77 (.A2( u1_u11_X_25 ) , .A1( u1_u11_X_26 ) , .ZN( u1_u11_u4_n104 ) );
  AND2_X1 u1_u11_u4_U78 (.A1( u1_u11_X_30 ) , .A2( u1_u11_u4_n176 ) , .ZN( u1_u11_u4_n99 ) );
  AND2_X1 u1_u11_u4_U79 (.A1( u1_u11_X_26 ) , .ZN( u1_u11_u4_n101 ) , .A2( u1_u11_u4_n177 ) );
  AOI21_X1 u1_u11_u4_U8 (.ZN( u1_u11_u4_n109 ) , .A( u1_u11_u4_n153 ) , .B1( u1_u11_u4_n159 ) , .B2( u1_u11_u4_n184 ) );
  AND2_X1 u1_u11_u4_U80 (.A1( u1_u11_X_27 ) , .A2( u1_u11_X_30 ) , .ZN( u1_u11_u4_n103 ) );
  INV_X1 u1_u11_u4_U81 (.A( u1_u11_X_28 ) , .ZN( u1_u11_u4_n169 ) );
  INV_X1 u1_u11_u4_U82 (.A( u1_u11_X_29 ) , .ZN( u1_u11_u4_n168 ) );
  INV_X1 u1_u11_u4_U83 (.A( u1_u11_X_25 ) , .ZN( u1_u11_u4_n177 ) );
  INV_X1 u1_u11_u4_U84 (.A( u1_u11_X_27 ) , .ZN( u1_u11_u4_n176 ) );
  NAND4_X1 u1_u11_u4_U85 (.ZN( u1_out11_25 ) , .A4( u1_u11_u4_n139 ) , .A3( u1_u11_u4_n140 ) , .A2( u1_u11_u4_n141 ) , .A1( u1_u11_u4_n142 ) );
  OAI21_X1 u1_u11_u4_U86 (.A( u1_u11_u4_n128 ) , .B2( u1_u11_u4_n129 ) , .B1( u1_u11_u4_n130 ) , .ZN( u1_u11_u4_n142 ) );
  OAI21_X1 u1_u11_u4_U87 (.B2( u1_u11_u4_n131 ) , .ZN( u1_u11_u4_n141 ) , .A( u1_u11_u4_n175 ) , .B1( u1_u11_u4_n183 ) );
  NAND4_X1 u1_u11_u4_U88 (.ZN( u1_out11_14 ) , .A4( u1_u11_u4_n124 ) , .A3( u1_u11_u4_n125 ) , .A2( u1_u11_u4_n126 ) , .A1( u1_u11_u4_n127 ) );
  AOI22_X1 u1_u11_u4_U89 (.B2( u1_u11_u4_n117 ) , .ZN( u1_u11_u4_n126 ) , .A1( u1_u11_u4_n129 ) , .B1( u1_u11_u4_n152 ) , .A2( u1_u11_u4_n175 ) );
  AOI211_X1 u1_u11_u4_U9 (.B( u1_u11_u4_n136 ) , .A( u1_u11_u4_n137 ) , .C2( u1_u11_u4_n138 ) , .ZN( u1_u11_u4_n139 ) , .C1( u1_u11_u4_n182 ) );
  AOI22_X1 u1_u11_u4_U90 (.ZN( u1_u11_u4_n125 ) , .B2( u1_u11_u4_n131 ) , .A2( u1_u11_u4_n132 ) , .B1( u1_u11_u4_n138 ) , .A1( u1_u11_u4_n178 ) );
  NAND4_X1 u1_u11_u4_U91 (.ZN( u1_out11_8 ) , .A4( u1_u11_u4_n110 ) , .A3( u1_u11_u4_n111 ) , .A2( u1_u11_u4_n112 ) , .A1( u1_u11_u4_n186 ) );
  NAND2_X1 u1_u11_u4_U92 (.ZN( u1_u11_u4_n112 ) , .A2( u1_u11_u4_n130 ) , .A1( u1_u11_u4_n150 ) );
  AOI22_X1 u1_u11_u4_U93 (.ZN( u1_u11_u4_n111 ) , .B2( u1_u11_u4_n132 ) , .A1( u1_u11_u4_n152 ) , .B1( u1_u11_u4_n178 ) , .A2( u1_u11_u4_n97 ) );
  AOI22_X1 u1_u11_u4_U94 (.B2( u1_u11_u4_n149 ) , .B1( u1_u11_u4_n150 ) , .A2( u1_u11_u4_n151 ) , .A1( u1_u11_u4_n152 ) , .ZN( u1_u11_u4_n167 ) );
  NOR4_X1 u1_u11_u4_U95 (.A4( u1_u11_u4_n162 ) , .A3( u1_u11_u4_n163 ) , .A2( u1_u11_u4_n164 ) , .A1( u1_u11_u4_n165 ) , .ZN( u1_u11_u4_n166 ) );
  NAND3_X1 u1_u11_u4_U96 (.ZN( u1_out11_3 ) , .A3( u1_u11_u4_n166 ) , .A1( u1_u11_u4_n167 ) , .A2( u1_u11_u4_n186 ) );
  NAND3_X1 u1_u11_u4_U97 (.A3( u1_u11_u4_n146 ) , .A2( u1_u11_u4_n147 ) , .A1( u1_u11_u4_n148 ) , .ZN( u1_u11_u4_n149 ) );
  NAND3_X1 u1_u11_u4_U98 (.A3( u1_u11_u4_n143 ) , .A2( u1_u11_u4_n144 ) , .A1( u1_u11_u4_n145 ) , .ZN( u1_u11_u4_n151 ) );
  NAND3_X1 u1_u11_u4_U99 (.A3( u1_u11_u4_n121 ) , .ZN( u1_u11_u4_n122 ) , .A2( u1_u11_u4_n144 ) , .A1( u1_u11_u4_n154 ) );
  XOR2_X1 u1_u12_U11 (.B( u1_K13_44 ) , .A( u1_R11_29 ) , .Z( u1_u12_X_44 ) );
  XOR2_X1 u1_u12_U12 (.B( u1_K13_43 ) , .A( u1_R11_28 ) , .Z( u1_u12_X_43 ) );
  XOR2_X1 u1_u12_U13 (.B( u1_K13_42 ) , .A( u1_R11_29 ) , .Z( u1_u12_X_42 ) );
  XOR2_X1 u1_u12_U14 (.B( u1_K13_41 ) , .A( u1_R11_28 ) , .Z( u1_u12_X_41 ) );
  XOR2_X1 u1_u12_U16 (.B( u1_K13_3 ) , .A( u1_R11_2 ) , .Z( u1_u12_X_3 ) );
  XOR2_X1 u1_u12_U18 (.B( u1_K13_38 ) , .A( u1_R11_25 ) , .Z( u1_u12_X_38 ) );
  XOR2_X1 u1_u12_U19 (.B( u1_K13_37 ) , .A( u1_R11_24 ) , .Z( u1_u12_X_37 ) );
  XOR2_X1 u1_u12_U2 (.B( u1_K13_8 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_8 ) );
  XOR2_X1 u1_u12_U20 (.B( u1_K13_36 ) , .A( u1_R11_25 ) , .Z( u1_u12_X_36 ) );
  XOR2_X1 u1_u12_U21 (.B( u1_K13_35 ) , .A( u1_R11_24 ) , .Z( u1_u12_X_35 ) );
  XOR2_X1 u1_u12_U24 (.B( u1_K13_32 ) , .A( u1_R11_21 ) , .Z( u1_u12_X_32 ) );
  XOR2_X1 u1_u12_U25 (.B( u1_K13_31 ) , .A( u1_R11_20 ) , .Z( u1_u12_X_31 ) );
  XOR2_X1 u1_u12_U26 (.B( u1_K13_30 ) , .A( u1_R11_21 ) , .Z( u1_u12_X_30 ) );
  XOR2_X1 u1_u12_U27 (.B( u1_K13_2 ) , .A( u1_R11_1 ) , .Z( u1_u12_X_2 ) );
  XOR2_X1 u1_u12_U28 (.B( u1_K13_29 ) , .A( u1_R11_20 ) , .Z( u1_u12_X_29 ) );
  XOR2_X1 u1_u12_U29 (.B( u1_K13_28 ) , .A( u1_R11_19 ) , .Z( u1_u12_X_28 ) );
  XOR2_X1 u1_u12_U3 (.B( u1_K13_7 ) , .A( u1_R11_4 ) , .Z( u1_u12_X_7 ) );
  XOR2_X1 u1_u12_U30 (.B( u1_K13_27 ) , .A( u1_R11_18 ) , .Z( u1_u12_X_27 ) );
  XOR2_X1 u1_u12_U31 (.B( u1_K13_26 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_26 ) );
  XOR2_X1 u1_u12_U32 (.B( u1_K13_25 ) , .A( u1_R11_16 ) , .Z( u1_u12_X_25 ) );
  XOR2_X1 u1_u12_U33 (.B( u1_K13_24 ) , .A( u1_R11_17 ) , .Z( u1_u12_X_24 ) );
  XOR2_X1 u1_u12_U34 (.B( u1_K13_23 ) , .A( u1_R11_16 ) , .Z( u1_u12_X_23 ) );
  XOR2_X1 u1_u12_U35 (.B( u1_K13_22 ) , .A( u1_R11_15 ) , .Z( u1_u12_X_22 ) );
  XOR2_X1 u1_u12_U36 (.B( u1_K13_21 ) , .A( u1_R11_14 ) , .Z( u1_u12_X_21 ) );
  XOR2_X1 u1_u12_U37 (.B( u1_K13_20 ) , .A( u1_R11_13 ) , .Z( u1_u12_X_20 ) );
  XOR2_X1 u1_u12_U38 (.B( u1_K13_1 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_1 ) );
  XOR2_X1 u1_u12_U39 (.B( u1_K13_19 ) , .A( u1_R11_12 ) , .Z( u1_u12_X_19 ) );
  XOR2_X1 u1_u12_U4 (.B( u1_K13_6 ) , .A( u1_R11_5 ) , .Z( u1_u12_X_6 ) );
  XOR2_X1 u1_u12_U40 (.B( u1_K13_18 ) , .A( u1_R11_13 ) , .Z( u1_u12_X_18 ) );
  XOR2_X1 u1_u12_U41 (.B( u1_K13_17 ) , .A( u1_R11_12 ) , .Z( u1_u12_X_17 ) );
  XOR2_X1 u1_u12_U44 (.B( u1_K13_14 ) , .A( u1_R11_9 ) , .Z( u1_u12_X_14 ) );
  XOR2_X1 u1_u12_U46 (.B( u1_K13_12 ) , .A( u1_R11_9 ) , .Z( u1_u12_X_12 ) );
  XOR2_X1 u1_u12_U5 (.B( u1_K13_5 ) , .A( u1_R11_4 ) , .Z( u1_u12_X_5 ) );
  XOR2_X1 u1_u12_U6 (.B( u1_K13_4 ) , .A( u1_R11_3 ) , .Z( u1_u12_X_4 ) );
  XOR2_X1 u1_u12_U7 (.B( u1_K13_48 ) , .A( u1_R11_1 ) , .Z( u1_u12_X_48 ) );
  XOR2_X1 u1_u12_U8 (.B( u1_K13_47 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_47 ) );
  NAND2_X1 u1_u12_u0_U10 (.ZN( u1_u12_u0_n113 ) , .A1( u1_u12_u0_n139 ) , .A2( u1_u12_u0_n149 ) );
  AND3_X1 u1_u12_u0_U11 (.A2( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n127 ) , .A3( u1_u12_u0_n130 ) , .A1( u1_u12_u0_n148 ) );
  AND2_X1 u1_u12_u0_U12 (.ZN( u1_u12_u0_n107 ) , .A1( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n140 ) );
  AND2_X1 u1_u12_u0_U13 (.A2( u1_u12_u0_n129 ) , .A1( u1_u12_u0_n130 ) , .ZN( u1_u12_u0_n151 ) );
  AND2_X1 u1_u12_u0_U14 (.A1( u1_u12_u0_n108 ) , .A2( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n145 ) );
  INV_X1 u1_u12_u0_U15 (.A( u1_u12_u0_n143 ) , .ZN( u1_u12_u0_n173 ) );
  NOR2_X1 u1_u12_u0_U16 (.A2( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n147 ) , .A1( u1_u12_u0_n160 ) );
  AOI21_X1 u1_u12_u0_U17 (.B1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n132 ) , .A( u1_u12_u0_n165 ) , .B2( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U18 (.A( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n165 ) );
  OAI22_X1 u1_u12_u0_U19 (.B1( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n147 ) , .A2( u1_u12_u0_n90 ) , .ZN( u1_u12_u0_n91 ) );
  AND3_X1 u1_u12_u0_U20 (.A3( u1_u12_u0_n121 ) , .A2( u1_u12_u0_n125 ) , .A1( u1_u12_u0_n148 ) , .ZN( u1_u12_u0_n90 ) );
  OAI22_X1 u1_u12_u0_U21 (.B1( u1_u12_u0_n125 ) , .ZN( u1_u12_u0_n126 ) , .A1( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n146 ) , .B2( u1_u12_u0_n147 ) );
  INV_X1 u1_u12_u0_U22 (.A( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n161 ) );
  AOI22_X1 u1_u12_u0_U23 (.B2( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n110 ) , .ZN( u1_u12_u0_n111 ) , .B1( u1_u12_u0_n118 ) , .A1( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U24 (.A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U25 (.A2( u1_u12_u0_n102 ) , .A1( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n149 ) );
  INV_X1 u1_u12_u0_U26 (.A( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n158 ) );
  NAND2_X1 u1_u12_u0_U27 (.A2( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n131 ) , .A1( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U28 (.ZN( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n92 ) , .A2( u1_u12_u0_n94 ) );
  AOI21_X1 u1_u12_u0_U29 (.ZN( u1_u12_u0_n104 ) , .B1( u1_u12_u0_n107 ) , .B2( u1_u12_u0_n141 ) , .A( u1_u12_u0_n144 ) );
  INV_X1 u1_u12_u0_U3 (.A( u1_u12_u0_n113 ) , .ZN( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U30 (.ZN( u1_u12_u0_n116 ) , .B2( u1_u12_u0_n142 ) , .A( u1_u12_u0_n144 ) , .B1( u1_u12_u0_n166 ) );
  AOI21_X1 u1_u12_u0_U31 (.B1( u1_u12_u0_n127 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n96 ) );
  NAND2_X1 u1_u12_u0_U32 (.A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n114 ) , .A1( u1_u12_u0_n92 ) );
  NOR2_X1 u1_u12_u0_U33 (.A1( u1_u12_u0_n120 ) , .ZN( u1_u12_u0_n143 ) , .A2( u1_u12_u0_n167 ) );
  OAI221_X1 u1_u12_u0_U34 (.C1( u1_u12_u0_n112 ) , .ZN( u1_u12_u0_n120 ) , .B1( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n141 ) , .C2( u1_u12_u0_n147 ) , .A( u1_u12_u0_n172 ) );
  AOI211_X1 u1_u12_u0_U35 (.B( u1_u12_u0_n115 ) , .A( u1_u12_u0_n116 ) , .C2( u1_u12_u0_n117 ) , .C1( u1_u12_u0_n118 ) , .ZN( u1_u12_u0_n119 ) );
  NAND2_X1 u1_u12_u0_U36 (.A1( u1_u12_u0_n100 ) , .A2( u1_u12_u0_n103 ) , .ZN( u1_u12_u0_n125 ) );
  NAND2_X1 u1_u12_u0_U37 (.A1( u1_u12_u0_n101 ) , .A2( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n150 ) );
  INV_X1 u1_u12_u0_U38 (.A( u1_u12_u0_n138 ) , .ZN( u1_u12_u0_n160 ) );
  NAND2_X1 u1_u12_u0_U39 (.A2( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n139 ) );
  AOI21_X1 u1_u12_u0_U4 (.B1( u1_u12_u0_n114 ) , .ZN( u1_u12_u0_n115 ) , .B2( u1_u12_u0_n129 ) , .A( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U40 (.A1( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n130 ) , .A2( u1_u12_u0_n94 ) );
  NAND2_X1 u1_u12_u0_U41 (.ZN( u1_u12_u0_n112 ) , .A2( u1_u12_u0_n92 ) , .A1( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U42 (.ZN( u1_u12_u0_n172 ) , .A( u1_u12_u0_n88 ) );
  OAI222_X1 u1_u12_u0_U43 (.C1( u1_u12_u0_n108 ) , .A1( u1_u12_u0_n125 ) , .B2( u1_u12_u0_n128 ) , .B1( u1_u12_u0_n144 ) , .A2( u1_u12_u0_n158 ) , .C2( u1_u12_u0_n161 ) , .ZN( u1_u12_u0_n88 ) );
  NAND2_X1 u1_u12_u0_U44 (.A2( u1_u12_u0_n101 ) , .ZN( u1_u12_u0_n121 ) , .A1( u1_u12_u0_n93 ) );
  OR3_X1 u1_u12_u0_U45 (.A3( u1_u12_u0_n152 ) , .A2( u1_u12_u0_n153 ) , .A1( u1_u12_u0_n154 ) , .ZN( u1_u12_u0_n155 ) );
  AOI21_X1 u1_u12_u0_U46 (.B2( u1_u12_u0_n150 ) , .B1( u1_u12_u0_n151 ) , .ZN( u1_u12_u0_n152 ) , .A( u1_u12_u0_n158 ) );
  AOI21_X1 u1_u12_u0_U47 (.A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n145 ) , .B1( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n154 ) );
  AOI21_X1 u1_u12_u0_U48 (.A( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n148 ) , .B1( u1_u12_u0_n149 ) , .ZN( u1_u12_u0_n153 ) );
  INV_X1 u1_u12_u0_U49 (.ZN( u1_u12_u0_n171 ) , .A( u1_u12_u0_n99 ) );
  AOI21_X1 u1_u12_u0_U5 (.B2( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n134 ) , .B1( u1_u12_u0_n151 ) , .A( u1_u12_u0_n158 ) );
  OAI211_X1 u1_u12_u0_U50 (.C2( u1_u12_u0_n140 ) , .C1( u1_u12_u0_n161 ) , .A( u1_u12_u0_n169 ) , .B( u1_u12_u0_n98 ) , .ZN( u1_u12_u0_n99 ) );
  INV_X1 u1_u12_u0_U51 (.ZN( u1_u12_u0_n169 ) , .A( u1_u12_u0_n91 ) );
  AOI211_X1 u1_u12_u0_U52 (.C1( u1_u12_u0_n118 ) , .A( u1_u12_u0_n123 ) , .B( u1_u12_u0_n96 ) , .C2( u1_u12_u0_n97 ) , .ZN( u1_u12_u0_n98 ) );
  NOR2_X1 u1_u12_u0_U53 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n118 ) );
  NOR2_X1 u1_u12_u0_U54 (.A2( u1_u12_X_1 ) , .ZN( u1_u12_u0_n101 ) , .A1( u1_u12_u0_n163 ) );
  NOR2_X1 u1_u12_u0_U55 (.A2( u1_u12_X_6 ) , .ZN( u1_u12_u0_n100 ) , .A1( u1_u12_u0_n162 ) );
  NAND2_X1 u1_u12_u0_U56 (.A2( u1_u12_X_4 ) , .A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n144 ) );
  NOR2_X1 u1_u12_u0_U57 (.A2( u1_u12_X_5 ) , .ZN( u1_u12_u0_n136 ) , .A1( u1_u12_u0_n159 ) );
  NAND2_X1 u1_u12_u0_U58 (.A1( u1_u12_X_5 ) , .ZN( u1_u12_u0_n138 ) , .A2( u1_u12_u0_n159 ) );
  AND2_X1 u1_u12_u0_U59 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n102 ) );
  NOR2_X1 u1_u12_u0_U6 (.A1( u1_u12_u0_n108 ) , .ZN( u1_u12_u0_n123 ) , .A2( u1_u12_u0_n158 ) );
  AND2_X1 u1_u12_u0_U60 (.A1( u1_u12_X_6 ) , .A2( u1_u12_u0_n162 ) , .ZN( u1_u12_u0_n93 ) );
  INV_X1 u1_u12_u0_U61 (.A( u1_u12_X_4 ) , .ZN( u1_u12_u0_n159 ) );
  INV_X1 u1_u12_u0_U62 (.A( u1_u12_X_1 ) , .ZN( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U63 (.A( u1_u12_X_3 ) , .ZN( u1_u12_u0_n162 ) );
  OR4_X1 u1_u12_u0_U64 (.ZN( u1_out12_17 ) , .A4( u1_u12_u0_n122 ) , .A2( u1_u12_u0_n123 ) , .A1( u1_u12_u0_n124 ) , .A3( u1_u12_u0_n170 ) );
  AOI21_X1 u1_u12_u0_U65 (.B2( u1_u12_u0_n107 ) , .ZN( u1_u12_u0_n124 ) , .B1( u1_u12_u0_n128 ) , .A( u1_u12_u0_n161 ) );
  INV_X1 u1_u12_u0_U66 (.A( u1_u12_u0_n111 ) , .ZN( u1_u12_u0_n170 ) );
  OR4_X1 u1_u12_u0_U67 (.ZN( u1_out12_31 ) , .A4( u1_u12_u0_n155 ) , .A2( u1_u12_u0_n156 ) , .A1( u1_u12_u0_n157 ) , .A3( u1_u12_u0_n173 ) );
  AOI21_X1 u1_u12_u0_U68 (.A( u1_u12_u0_n138 ) , .B2( u1_u12_u0_n139 ) , .B1( u1_u12_u0_n140 ) , .ZN( u1_u12_u0_n157 ) );
  AOI21_X1 u1_u12_u0_U69 (.B2( u1_u12_u0_n141 ) , .B1( u1_u12_u0_n142 ) , .ZN( u1_u12_u0_n156 ) , .A( u1_u12_u0_n161 ) );
  OAI21_X1 u1_u12_u0_U7 (.B1( u1_u12_u0_n150 ) , .B2( u1_u12_u0_n158 ) , .A( u1_u12_u0_n172 ) , .ZN( u1_u12_u0_n89 ) );
  INV_X1 u1_u12_u0_U70 (.ZN( u1_u12_u0_n174 ) , .A( u1_u12_u0_n89 ) );
  AOI211_X1 u1_u12_u0_U71 (.B( u1_u12_u0_n104 ) , .A( u1_u12_u0_n105 ) , .ZN( u1_u12_u0_n106 ) , .C2( u1_u12_u0_n113 ) , .C1( u1_u12_u0_n160 ) );
  INV_X1 u1_u12_u0_U72 (.A( u1_u12_u0_n126 ) , .ZN( u1_u12_u0_n168 ) );
  AOI211_X1 u1_u12_u0_U73 (.B( u1_u12_u0_n133 ) , .A( u1_u12_u0_n134 ) , .C2( u1_u12_u0_n135 ) , .C1( u1_u12_u0_n136 ) , .ZN( u1_u12_u0_n137 ) );
  NOR2_X1 u1_u12_u0_U74 (.A1( u1_u12_u0_n163 ) , .A2( u1_u12_u0_n164 ) , .ZN( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U75 (.A2( u1_u12_X_3 ) , .A1( u1_u12_X_6 ) , .ZN( u1_u12_u0_n94 ) );
  OAI221_X1 u1_u12_u0_U76 (.C1( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n122 ) , .B2( u1_u12_u0_n127 ) , .A( u1_u12_u0_n143 ) , .B1( u1_u12_u0_n144 ) , .C2( u1_u12_u0_n147 ) );
  AOI21_X1 u1_u12_u0_U77 (.B1( u1_u12_u0_n132 ) , .ZN( u1_u12_u0_n133 ) , .A( u1_u12_u0_n144 ) , .B2( u1_u12_u0_n166 ) );
  OAI22_X1 u1_u12_u0_U78 (.ZN( u1_u12_u0_n105 ) , .A2( u1_u12_u0_n132 ) , .B1( u1_u12_u0_n146 ) , .A1( u1_u12_u0_n147 ) , .B2( u1_u12_u0_n161 ) );
  NAND2_X1 u1_u12_u0_U79 (.ZN( u1_u12_u0_n110 ) , .A2( u1_u12_u0_n132 ) , .A1( u1_u12_u0_n145 ) );
  AND2_X1 u1_u12_u0_U8 (.A1( u1_u12_u0_n114 ) , .A2( u1_u12_u0_n121 ) , .ZN( u1_u12_u0_n146 ) );
  INV_X1 u1_u12_u0_U80 (.A( u1_u12_u0_n119 ) , .ZN( u1_u12_u0_n167 ) );
  NAND2_X1 u1_u12_u0_U81 (.ZN( u1_u12_u0_n148 ) , .A1( u1_u12_u0_n93 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U82 (.A1( u1_u12_u0_n100 ) , .ZN( u1_u12_u0_n129 ) , .A2( u1_u12_u0_n95 ) );
  NAND2_X1 u1_u12_u0_U83 (.A1( u1_u12_u0_n102 ) , .ZN( u1_u12_u0_n128 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U84 (.A2( u1_u12_X_1 ) , .A1( u1_u12_X_2 ) , .ZN( u1_u12_u0_n92 ) );
  NAND2_X1 u1_u12_u0_U85 (.ZN( u1_u12_u0_n142 ) , .A1( u1_u12_u0_n94 ) , .A2( u1_u12_u0_n95 ) );
  NOR2_X1 u1_u12_u0_U86 (.A2( u1_u12_X_2 ) , .ZN( u1_u12_u0_n103 ) , .A1( u1_u12_u0_n164 ) );
  INV_X1 u1_u12_u0_U87 (.A( u1_u12_X_2 ) , .ZN( u1_u12_u0_n163 ) );
  NAND3_X1 u1_u12_u0_U88 (.ZN( u1_out12_23 ) , .A3( u1_u12_u0_n137 ) , .A1( u1_u12_u0_n168 ) , .A2( u1_u12_u0_n171 ) );
  NAND3_X1 u1_u12_u0_U89 (.A3( u1_u12_u0_n127 ) , .A2( u1_u12_u0_n128 ) , .ZN( u1_u12_u0_n135 ) , .A1( u1_u12_u0_n150 ) );
  AND2_X1 u1_u12_u0_U9 (.A1( u1_u12_u0_n131 ) , .ZN( u1_u12_u0_n141 ) , .A2( u1_u12_u0_n150 ) );
  NAND3_X1 u1_u12_u0_U90 (.ZN( u1_u12_u0_n117 ) , .A3( u1_u12_u0_n132 ) , .A2( u1_u12_u0_n139 ) , .A1( u1_u12_u0_n148 ) );
  NAND3_X1 u1_u12_u0_U91 (.ZN( u1_u12_u0_n109 ) , .A2( u1_u12_u0_n114 ) , .A3( u1_u12_u0_n140 ) , .A1( u1_u12_u0_n149 ) );
  NAND3_X1 u1_u12_u0_U92 (.ZN( u1_out12_9 ) , .A3( u1_u12_u0_n106 ) , .A2( u1_u12_u0_n171 ) , .A1( u1_u12_u0_n174 ) );
  NAND3_X1 u1_u12_u0_U93 (.A2( u1_u12_u0_n128 ) , .A1( u1_u12_u0_n132 ) , .A3( u1_u12_u0_n146 ) , .ZN( u1_u12_u0_n97 ) );
  OAI22_X1 u1_u12_u3_U10 (.B1( u1_u12_u3_n113 ) , .A2( u1_u12_u3_n135 ) , .A1( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n164 ) , .ZN( u1_u12_u3_n98 ) );
  OAI211_X1 u1_u12_u3_U11 (.B( u1_u12_u3_n106 ) , .ZN( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n128 ) , .C1( u1_u12_u3_n167 ) , .A( u1_u12_u3_n181 ) );
  AOI221_X1 u1_u12_u3_U12 (.C1( u1_u12_u3_n105 ) , .ZN( u1_u12_u3_n106 ) , .A( u1_u12_u3_n131 ) , .B2( u1_u12_u3_n132 ) , .C2( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n169 ) );
  INV_X1 u1_u12_u3_U13 (.ZN( u1_u12_u3_n181 ) , .A( u1_u12_u3_n98 ) );
  NAND2_X1 u1_u12_u3_U14 (.ZN( u1_u12_u3_n105 ) , .A2( u1_u12_u3_n130 ) , .A1( u1_u12_u3_n155 ) );
  AOI22_X1 u1_u12_u3_U15 (.B1( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n116 ) , .ZN( u1_u12_u3_n123 ) , .B2( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U16 (.ZN( u1_u12_u3_n116 ) , .A2( u1_u12_u3_n151 ) , .A1( u1_u12_u3_n182 ) );
  NOR2_X1 u1_u12_u3_U17 (.ZN( u1_u12_u3_n126 ) , .A2( u1_u12_u3_n150 ) , .A1( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U18 (.ZN( u1_u12_u3_n112 ) , .B2( u1_u12_u3_n146 ) , .B1( u1_u12_u3_n155 ) , .A( u1_u12_u3_n167 ) );
  NAND2_X1 u1_u12_u3_U19 (.A1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n142 ) , .A2( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U20 (.ZN( u1_u12_u3_n132 ) , .A2( u1_u12_u3_n152 ) , .A1( u1_u12_u3_n156 ) );
  AND2_X1 u1_u12_u3_U21 (.A2( u1_u12_u3_n113 ) , .A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n151 ) );
  INV_X1 u1_u12_u3_U22 (.A( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n165 ) );
  INV_X1 u1_u12_u3_U23 (.A( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n170 ) );
  NAND2_X1 u1_u12_u3_U24 (.A1( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .ZN( u1_u12_u3_n140 ) );
  NAND2_X1 u1_u12_u3_U25 (.ZN( u1_u12_u3_n117 ) , .A1( u1_u12_u3_n124 ) , .A2( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U26 (.ZN( u1_u12_u3_n143 ) , .A1( u1_u12_u3_n165 ) , .A2( u1_u12_u3_n167 ) );
  INV_X1 u1_u12_u3_U27 (.A( u1_u12_u3_n130 ) , .ZN( u1_u12_u3_n177 ) );
  INV_X1 u1_u12_u3_U28 (.A( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n176 ) );
  INV_X1 u1_u12_u3_U29 (.A( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n174 ) );
  INV_X1 u1_u12_u3_U3 (.A( u1_u12_u3_n129 ) , .ZN( u1_u12_u3_n183 ) );
  INV_X1 u1_u12_u3_U30 (.A( u1_u12_u3_n139 ) , .ZN( u1_u12_u3_n185 ) );
  NOR2_X1 u1_u12_u3_U31 (.ZN( u1_u12_u3_n135 ) , .A2( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n169 ) );
  OAI222_X1 u1_u12_u3_U32 (.C2( u1_u12_u3_n107 ) , .A2( u1_u12_u3_n108 ) , .B1( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n138 ) , .B2( u1_u12_u3_n146 ) , .C1( u1_u12_u3_n154 ) , .A1( u1_u12_u3_n164 ) );
  NOR4_X1 u1_u12_u3_U33 (.A4( u1_u12_u3_n157 ) , .A3( u1_u12_u3_n158 ) , .A2( u1_u12_u3_n159 ) , .A1( u1_u12_u3_n160 ) , .ZN( u1_u12_u3_n161 ) );
  AOI21_X1 u1_u12_u3_U34 (.B2( u1_u12_u3_n152 ) , .B1( u1_u12_u3_n153 ) , .ZN( u1_u12_u3_n158 ) , .A( u1_u12_u3_n164 ) );
  AOI21_X1 u1_u12_u3_U35 (.A( u1_u12_u3_n154 ) , .B2( u1_u12_u3_n155 ) , .B1( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n157 ) );
  AOI21_X1 u1_u12_u3_U36 (.A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n150 ) , .B1( u1_u12_u3_n151 ) , .ZN( u1_u12_u3_n159 ) );
  AOI211_X1 u1_u12_u3_U37 (.ZN( u1_u12_u3_n109 ) , .A( u1_u12_u3_n119 ) , .C2( u1_u12_u3_n129 ) , .B( u1_u12_u3_n138 ) , .C1( u1_u12_u3_n141 ) );
  AOI211_X1 u1_u12_u3_U38 (.B( u1_u12_u3_n119 ) , .A( u1_u12_u3_n120 ) , .C2( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n122 ) , .C1( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U39 (.A( u1_u12_u3_n156 ) , .ZN( u1_u12_u3_n179 ) );
  INV_X1 u1_u12_u3_U4 (.A( u1_u12_u3_n140 ) , .ZN( u1_u12_u3_n182 ) );
  OAI22_X1 u1_u12_u3_U40 (.B1( u1_u12_u3_n118 ) , .ZN( u1_u12_u3_n120 ) , .A1( u1_u12_u3_n135 ) , .B2( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n178 ) );
  AND3_X1 u1_u12_u3_U41 (.ZN( u1_u12_u3_n118 ) , .A2( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n144 ) , .A3( u1_u12_u3_n152 ) );
  INV_X1 u1_u12_u3_U42 (.A( u1_u12_u3_n121 ) , .ZN( u1_u12_u3_n164 ) );
  NAND2_X1 u1_u12_u3_U43 (.ZN( u1_u12_u3_n133 ) , .A1( u1_u12_u3_n154 ) , .A2( u1_u12_u3_n164 ) );
  OAI211_X1 u1_u12_u3_U44 (.B( u1_u12_u3_n127 ) , .ZN( u1_u12_u3_n139 ) , .C1( u1_u12_u3_n150 ) , .C2( u1_u12_u3_n154 ) , .A( u1_u12_u3_n184 ) );
  INV_X1 u1_u12_u3_U45 (.A( u1_u12_u3_n125 ) , .ZN( u1_u12_u3_n184 ) );
  AOI221_X1 u1_u12_u3_U46 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n127 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n169 ) , .B2( u1_u12_u3_n170 ) , .B1( u1_u12_u3_n174 ) );
  OAI22_X1 u1_u12_u3_U47 (.A1( u1_u12_u3_n124 ) , .ZN( u1_u12_u3_n125 ) , .B2( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n165 ) , .B1( u1_u12_u3_n167 ) );
  NOR2_X1 u1_u12_u3_U48 (.A1( u1_u12_u3_n113 ) , .ZN( u1_u12_u3_n131 ) , .A2( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U49 (.A1( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n150 ) , .A2( u1_u12_u3_n99 ) );
  INV_X1 u1_u12_u3_U5 (.A( u1_u12_u3_n117 ) , .ZN( u1_u12_u3_n178 ) );
  NAND2_X1 u1_u12_u3_U50 (.A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n155 ) , .A1( u1_u12_u3_n97 ) );
  INV_X1 u1_u12_u3_U51 (.A( u1_u12_u3_n141 ) , .ZN( u1_u12_u3_n167 ) );
  AOI21_X1 u1_u12_u3_U52 (.B2( u1_u12_u3_n114 ) , .B1( u1_u12_u3_n146 ) , .A( u1_u12_u3_n154 ) , .ZN( u1_u12_u3_n94 ) );
  AOI21_X1 u1_u12_u3_U53 (.ZN( u1_u12_u3_n110 ) , .B2( u1_u12_u3_n142 ) , .B1( u1_u12_u3_n186 ) , .A( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U54 (.A( u1_u12_u3_n145 ) , .ZN( u1_u12_u3_n186 ) );
  AOI21_X1 u1_u12_u3_U55 (.B1( u1_u12_u3_n124 ) , .A( u1_u12_u3_n149 ) , .B2( u1_u12_u3_n155 ) , .ZN( u1_u12_u3_n95 ) );
  INV_X1 u1_u12_u3_U56 (.A( u1_u12_u3_n149 ) , .ZN( u1_u12_u3_n169 ) );
  NAND2_X1 u1_u12_u3_U57 (.ZN( u1_u12_u3_n124 ) , .A1( u1_u12_u3_n96 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U58 (.A2( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n146 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U59 (.A1( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n145 ) , .A2( u1_u12_u3_n99 ) );
  AOI221_X1 u1_u12_u3_U6 (.A( u1_u12_u3_n131 ) , .C2( u1_u12_u3_n132 ) , .C1( u1_u12_u3_n133 ) , .ZN( u1_u12_u3_n134 ) , .B1( u1_u12_u3_n143 ) , .B2( u1_u12_u3_n177 ) );
  NAND2_X1 u1_u12_u3_U60 (.A1( u1_u12_u3_n100 ) , .ZN( u1_u12_u3_n156 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U61 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n148 ) );
  NAND2_X1 u1_u12_u3_U62 (.A1( u1_u12_u3_n100 ) , .A2( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n128 ) );
  NAND2_X1 u1_u12_u3_U63 (.A2( u1_u12_u3_n101 ) , .A1( u1_u12_u3_n102 ) , .ZN( u1_u12_u3_n152 ) );
  NAND2_X1 u1_u12_u3_U64 (.A2( u1_u12_u3_n101 ) , .ZN( u1_u12_u3_n114 ) , .A1( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U65 (.ZN( u1_u12_u3_n107 ) , .A1( u1_u12_u3_n97 ) , .A2( u1_u12_u3_n99 ) );
  NAND2_X1 u1_u12_u3_U66 (.A2( u1_u12_u3_n100 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n113 ) );
  NAND2_X1 u1_u12_u3_U67 (.A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n153 ) , .A2( u1_u12_u3_n97 ) );
  NAND2_X1 u1_u12_u3_U68 (.A2( u1_u12_u3_n103 ) , .A1( u1_u12_u3_n104 ) , .ZN( u1_u12_u3_n130 ) );
  NAND2_X1 u1_u12_u3_U69 (.A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n96 ) );
  OAI22_X1 u1_u12_u3_U7 (.B2( u1_u12_u3_n147 ) , .A2( u1_u12_u3_n148 ) , .ZN( u1_u12_u3_n160 ) , .B1( u1_u12_u3_n165 ) , .A1( u1_u12_u3_n168 ) );
  NAND2_X1 u1_u12_u3_U70 (.A1( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n103 ) , .ZN( u1_u12_u3_n108 ) );
  NOR2_X1 u1_u12_u3_U71 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n99 ) );
  NOR2_X1 u1_u12_u3_U72 (.A2( u1_u12_X_21 ) , .A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n103 ) );
  NOR2_X1 u1_u12_u3_U73 (.A2( u1_u12_X_24 ) , .A1( u1_u12_u3_n171 ) , .ZN( u1_u12_u3_n97 ) );
  NOR2_X1 u1_u12_u3_U74 (.A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n141 ) , .A1( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U75 (.A2( u1_u12_X_19 ) , .A1( u1_u12_u3_n172 ) , .ZN( u1_u12_u3_n96 ) );
  NAND2_X1 u1_u12_u3_U76 (.A1( u1_u12_X_22 ) , .A2( u1_u12_X_23 ) , .ZN( u1_u12_u3_n154 ) );
  NAND2_X1 u1_u12_u3_U77 (.A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n149 ) , .A2( u1_u12_u3_n166 ) );
  NOR2_X1 u1_u12_u3_U78 (.A2( u1_u12_X_22 ) , .A1( u1_u12_X_23 ) , .ZN( u1_u12_u3_n121 ) );
  AND2_X1 u1_u12_u3_U79 (.A1( u1_u12_X_24 ) , .ZN( u1_u12_u3_n101 ) , .A2( u1_u12_u3_n171 ) );
  AND3_X1 u1_u12_u3_U8 (.A3( u1_u12_u3_n144 ) , .A2( u1_u12_u3_n145 ) , .A1( u1_u12_u3_n146 ) , .ZN( u1_u12_u3_n147 ) );
  AND2_X1 u1_u12_u3_U80 (.A1( u1_u12_X_19 ) , .ZN( u1_u12_u3_n102 ) , .A2( u1_u12_u3_n172 ) );
  AND2_X1 u1_u12_u3_U81 (.A1( u1_u12_X_21 ) , .A2( u1_u12_X_24 ) , .ZN( u1_u12_u3_n100 ) );
  AND2_X1 u1_u12_u3_U82 (.A2( u1_u12_X_19 ) , .A1( u1_u12_X_20 ) , .ZN( u1_u12_u3_n104 ) );
  INV_X1 u1_u12_u3_U83 (.A( u1_u12_X_22 ) , .ZN( u1_u12_u3_n166 ) );
  INV_X1 u1_u12_u3_U84 (.A( u1_u12_X_21 ) , .ZN( u1_u12_u3_n171 ) );
  INV_X1 u1_u12_u3_U85 (.A( u1_u12_X_20 ) , .ZN( u1_u12_u3_n172 ) );
  NAND4_X1 u1_u12_u3_U86 (.ZN( u1_out12_26 ) , .A4( u1_u12_u3_n109 ) , .A3( u1_u12_u3_n110 ) , .A2( u1_u12_u3_n111 ) , .A1( u1_u12_u3_n173 ) );
  INV_X1 u1_u12_u3_U87 (.ZN( u1_u12_u3_n173 ) , .A( u1_u12_u3_n94 ) );
  OAI21_X1 u1_u12_u3_U88 (.ZN( u1_u12_u3_n111 ) , .B2( u1_u12_u3_n117 ) , .A( u1_u12_u3_n133 ) , .B1( u1_u12_u3_n176 ) );
  NAND4_X1 u1_u12_u3_U89 (.ZN( u1_out12_20 ) , .A4( u1_u12_u3_n122 ) , .A3( u1_u12_u3_n123 ) , .A1( u1_u12_u3_n175 ) , .A2( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U9 (.A( u1_u12_u3_n143 ) , .ZN( u1_u12_u3_n168 ) );
  INV_X1 u1_u12_u3_U90 (.A( u1_u12_u3_n126 ) , .ZN( u1_u12_u3_n180 ) );
  INV_X1 u1_u12_u3_U91 (.A( u1_u12_u3_n112 ) , .ZN( u1_u12_u3_n175 ) );
  NAND4_X1 u1_u12_u3_U92 (.ZN( u1_out12_1 ) , .A4( u1_u12_u3_n161 ) , .A3( u1_u12_u3_n162 ) , .A2( u1_u12_u3_n163 ) , .A1( u1_u12_u3_n185 ) );
  NAND2_X1 u1_u12_u3_U93 (.ZN( u1_u12_u3_n163 ) , .A2( u1_u12_u3_n170 ) , .A1( u1_u12_u3_n176 ) );
  AOI22_X1 u1_u12_u3_U94 (.B2( u1_u12_u3_n140 ) , .B1( u1_u12_u3_n141 ) , .A2( u1_u12_u3_n142 ) , .ZN( u1_u12_u3_n162 ) , .A1( u1_u12_u3_n177 ) );
  OR4_X1 u1_u12_u3_U95 (.ZN( u1_out12_10 ) , .A4( u1_u12_u3_n136 ) , .A3( u1_u12_u3_n137 ) , .A1( u1_u12_u3_n138 ) , .A2( u1_u12_u3_n139 ) );
  OAI222_X1 u1_u12_u3_U96 (.C1( u1_u12_u3_n128 ) , .ZN( u1_u12_u3_n137 ) , .B1( u1_u12_u3_n148 ) , .A2( u1_u12_u3_n150 ) , .B2( u1_u12_u3_n154 ) , .C2( u1_u12_u3_n164 ) , .A1( u1_u12_u3_n167 ) );
  OAI221_X1 u1_u12_u3_U97 (.A( u1_u12_u3_n134 ) , .B2( u1_u12_u3_n135 ) , .ZN( u1_u12_u3_n136 ) , .C1( u1_u12_u3_n149 ) , .B1( u1_u12_u3_n151 ) , .C2( u1_u12_u3_n183 ) );
  NAND3_X1 u1_u12_u3_U98 (.A1( u1_u12_u3_n114 ) , .ZN( u1_u12_u3_n115 ) , .A2( u1_u12_u3_n145 ) , .A3( u1_u12_u3_n153 ) );
  NAND3_X1 u1_u12_u3_U99 (.ZN( u1_u12_u3_n129 ) , .A2( u1_u12_u3_n144 ) , .A1( u1_u12_u3_n153 ) , .A3( u1_u12_u3_n182 ) );
  OAI22_X1 u1_u12_u4_U10 (.B2( u1_u12_u4_n135 ) , .ZN( u1_u12_u4_n137 ) , .B1( u1_u12_u4_n153 ) , .A1( u1_u12_u4_n155 ) , .A2( u1_u12_u4_n171 ) );
  AND3_X1 u1_u12_u4_U11 (.A2( u1_u12_u4_n134 ) , .ZN( u1_u12_u4_n135 ) , .A3( u1_u12_u4_n145 ) , .A1( u1_u12_u4_n157 ) );
  NAND2_X1 u1_u12_u4_U12 (.ZN( u1_u12_u4_n132 ) , .A2( u1_u12_u4_n170 ) , .A1( u1_u12_u4_n173 ) );
  AOI21_X1 u1_u12_u4_U13 (.B2( u1_u12_u4_n160 ) , .B1( u1_u12_u4_n161 ) , .ZN( u1_u12_u4_n162 ) , .A( u1_u12_u4_n170 ) );
  AOI21_X1 u1_u12_u4_U14 (.ZN( u1_u12_u4_n107 ) , .B2( u1_u12_u4_n143 ) , .A( u1_u12_u4_n174 ) , .B1( u1_u12_u4_n184 ) );
  AOI21_X1 u1_u12_u4_U15 (.B2( u1_u12_u4_n158 ) , .B1( u1_u12_u4_n159 ) , .ZN( u1_u12_u4_n163 ) , .A( u1_u12_u4_n174 ) );
  AOI21_X1 u1_u12_u4_U16 (.A( u1_u12_u4_n153 ) , .B2( u1_u12_u4_n154 ) , .B1( u1_u12_u4_n155 ) , .ZN( u1_u12_u4_n165 ) );
  AOI21_X1 u1_u12_u4_U17 (.A( u1_u12_u4_n156 ) , .B2( u1_u12_u4_n157 ) , .ZN( u1_u12_u4_n164 ) , .B1( u1_u12_u4_n184 ) );
  INV_X1 u1_u12_u4_U18 (.A( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n170 ) );
  AND2_X1 u1_u12_u4_U19 (.A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n155 ) , .A1( u1_u12_u4_n160 ) );
  INV_X1 u1_u12_u4_U20 (.A( u1_u12_u4_n156 ) , .ZN( u1_u12_u4_n175 ) );
  NAND2_X1 u1_u12_u4_U21 (.A2( u1_u12_u4_n118 ) , .ZN( u1_u12_u4_n131 ) , .A1( u1_u12_u4_n147 ) );
  NAND2_X1 u1_u12_u4_U22 (.A1( u1_u12_u4_n119 ) , .A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n130 ) );
  NAND2_X1 u1_u12_u4_U23 (.ZN( u1_u12_u4_n117 ) , .A2( u1_u12_u4_n118 ) , .A1( u1_u12_u4_n148 ) );
  NAND2_X1 u1_u12_u4_U24 (.ZN( u1_u12_u4_n129 ) , .A1( u1_u12_u4_n134 ) , .A2( u1_u12_u4_n148 ) );
  AND3_X1 u1_u12_u4_U25 (.A1( u1_u12_u4_n119 ) , .A2( u1_u12_u4_n143 ) , .A3( u1_u12_u4_n154 ) , .ZN( u1_u12_u4_n161 ) );
  AND2_X1 u1_u12_u4_U26 (.A1( u1_u12_u4_n145 ) , .A2( u1_u12_u4_n147 ) , .ZN( u1_u12_u4_n159 ) );
  OR3_X1 u1_u12_u4_U27 (.A3( u1_u12_u4_n114 ) , .A2( u1_u12_u4_n115 ) , .A1( u1_u12_u4_n116 ) , .ZN( u1_u12_u4_n136 ) );
  AOI21_X1 u1_u12_u4_U28 (.A( u1_u12_u4_n113 ) , .ZN( u1_u12_u4_n116 ) , .B2( u1_u12_u4_n173 ) , .B1( u1_u12_u4_n174 ) );
  AOI21_X1 u1_u12_u4_U29 (.ZN( u1_u12_u4_n115 ) , .B2( u1_u12_u4_n145 ) , .B1( u1_u12_u4_n146 ) , .A( u1_u12_u4_n156 ) );
  NOR2_X1 u1_u12_u4_U3 (.ZN( u1_u12_u4_n121 ) , .A1( u1_u12_u4_n181 ) , .A2( u1_u12_u4_n182 ) );
  OAI22_X1 u1_u12_u4_U30 (.ZN( u1_u12_u4_n114 ) , .A2( u1_u12_u4_n121 ) , .B1( u1_u12_u4_n160 ) , .B2( u1_u12_u4_n170 ) , .A1( u1_u12_u4_n171 ) );
  INV_X1 u1_u12_u4_U31 (.A( u1_u12_u4_n158 ) , .ZN( u1_u12_u4_n182 ) );
  INV_X1 u1_u12_u4_U32 (.ZN( u1_u12_u4_n181 ) , .A( u1_u12_u4_n96 ) );
  INV_X1 u1_u12_u4_U33 (.A( u1_u12_u4_n144 ) , .ZN( u1_u12_u4_n179 ) );
  INV_X1 u1_u12_u4_U34 (.A( u1_u12_u4_n157 ) , .ZN( u1_u12_u4_n178 ) );
  NAND2_X1 u1_u12_u4_U35 (.A2( u1_u12_u4_n154 ) , .A1( u1_u12_u4_n96 ) , .ZN( u1_u12_u4_n97 ) );
  INV_X1 u1_u12_u4_U36 (.ZN( u1_u12_u4_n186 ) , .A( u1_u12_u4_n95 ) );
  OAI221_X1 u1_u12_u4_U37 (.C1( u1_u12_u4_n134 ) , .B1( u1_u12_u4_n158 ) , .B2( u1_u12_u4_n171 ) , .C2( u1_u12_u4_n173 ) , .A( u1_u12_u4_n94 ) , .ZN( u1_u12_u4_n95 ) );
  AOI222_X1 u1_u12_u4_U38 (.B2( u1_u12_u4_n132 ) , .A1( u1_u12_u4_n138 ) , .C2( u1_u12_u4_n175 ) , .A2( u1_u12_u4_n179 ) , .C1( u1_u12_u4_n181 ) , .B1( u1_u12_u4_n185 ) , .ZN( u1_u12_u4_n94 ) );
  INV_X1 u1_u12_u4_U39 (.A( u1_u12_u4_n113 ) , .ZN( u1_u12_u4_n185 ) );
  INV_X1 u1_u12_u4_U4 (.A( u1_u12_u4_n117 ) , .ZN( u1_u12_u4_n184 ) );
  INV_X1 u1_u12_u4_U40 (.A( u1_u12_u4_n143 ) , .ZN( u1_u12_u4_n183 ) );
  NOR2_X1 u1_u12_u4_U41 (.ZN( u1_u12_u4_n138 ) , .A1( u1_u12_u4_n168 ) , .A2( u1_u12_u4_n169 ) );
  NOR2_X1 u1_u12_u4_U42 (.A1( u1_u12_u4_n150 ) , .A2( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n153 ) );
  NOR2_X1 u1_u12_u4_U43 (.A2( u1_u12_u4_n128 ) , .A1( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n156 ) );
  AOI22_X1 u1_u12_u4_U44 (.B2( u1_u12_u4_n122 ) , .A1( u1_u12_u4_n123 ) , .ZN( u1_u12_u4_n124 ) , .B1( u1_u12_u4_n128 ) , .A2( u1_u12_u4_n172 ) );
  INV_X1 u1_u12_u4_U45 (.A( u1_u12_u4_n153 ) , .ZN( u1_u12_u4_n172 ) );
  NAND2_X1 u1_u12_u4_U46 (.A2( u1_u12_u4_n120 ) , .ZN( u1_u12_u4_n123 ) , .A1( u1_u12_u4_n161 ) );
  AOI22_X1 u1_u12_u4_U47 (.B2( u1_u12_u4_n132 ) , .A2( u1_u12_u4_n133 ) , .ZN( u1_u12_u4_n140 ) , .A1( u1_u12_u4_n150 ) , .B1( u1_u12_u4_n179 ) );
  NAND2_X1 u1_u12_u4_U48 (.ZN( u1_u12_u4_n133 ) , .A2( u1_u12_u4_n146 ) , .A1( u1_u12_u4_n154 ) );
  NAND2_X1 u1_u12_u4_U49 (.A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n154 ) , .A2( u1_u12_u4_n98 ) );
  NOR4_X1 u1_u12_u4_U5 (.A4( u1_u12_u4_n106 ) , .A3( u1_u12_u4_n107 ) , .A2( u1_u12_u4_n108 ) , .A1( u1_u12_u4_n109 ) , .ZN( u1_u12_u4_n110 ) );
  NAND2_X1 u1_u12_u4_U50 (.A1( u1_u12_u4_n101 ) , .ZN( u1_u12_u4_n158 ) , .A2( u1_u12_u4_n99 ) );
  AOI21_X1 u1_u12_u4_U51 (.ZN( u1_u12_u4_n127 ) , .A( u1_u12_u4_n136 ) , .B2( u1_u12_u4_n150 ) , .B1( u1_u12_u4_n180 ) );
  INV_X1 u1_u12_u4_U52 (.A( u1_u12_u4_n160 ) , .ZN( u1_u12_u4_n180 ) );
  NAND2_X1 u1_u12_u4_U53 (.A2( u1_u12_u4_n104 ) , .A1( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n146 ) );
  NAND2_X1 u1_u12_u4_U54 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n160 ) );
  NAND2_X1 u1_u12_u4_U55 (.ZN( u1_u12_u4_n134 ) , .A1( u1_u12_u4_n98 ) , .A2( u1_u12_u4_n99 ) );
  NAND2_X1 u1_u12_u4_U56 (.A1( u1_u12_u4_n103 ) , .A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n143 ) );
  NAND2_X1 u1_u12_u4_U57 (.A2( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n145 ) , .A1( u1_u12_u4_n98 ) );
  NAND2_X1 u1_u12_u4_U58 (.A1( u1_u12_u4_n100 ) , .A2( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n120 ) );
  NAND2_X1 u1_u12_u4_U59 (.A1( u1_u12_u4_n102 ) , .A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n148 ) );
  AOI21_X1 u1_u12_u4_U6 (.ZN( u1_u12_u4_n106 ) , .B2( u1_u12_u4_n146 ) , .B1( u1_u12_u4_n158 ) , .A( u1_u12_u4_n170 ) );
  NAND2_X1 u1_u12_u4_U60 (.A2( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n157 ) );
  INV_X1 u1_u12_u4_U61 (.A( u1_u12_u4_n150 ) , .ZN( u1_u12_u4_n173 ) );
  INV_X1 u1_u12_u4_U62 (.A( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n171 ) );
  NAND2_X1 u1_u12_u4_U63 (.A1( u1_u12_u4_n100 ) , .ZN( u1_u12_u4_n118 ) , .A2( u1_u12_u4_n99 ) );
  NAND2_X1 u1_u12_u4_U64 (.A2( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n144 ) );
  NAND2_X1 u1_u12_u4_U65 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n105 ) , .ZN( u1_u12_u4_n96 ) );
  INV_X1 u1_u12_u4_U66 (.A( u1_u12_u4_n128 ) , .ZN( u1_u12_u4_n174 ) );
  NAND2_X1 u1_u12_u4_U67 (.A2( u1_u12_u4_n102 ) , .ZN( u1_u12_u4_n119 ) , .A1( u1_u12_u4_n98 ) );
  NAND2_X1 u1_u12_u4_U68 (.A2( u1_u12_u4_n101 ) , .A1( u1_u12_u4_n103 ) , .ZN( u1_u12_u4_n147 ) );
  NAND2_X1 u1_u12_u4_U69 (.A2( u1_u12_u4_n104 ) , .ZN( u1_u12_u4_n113 ) , .A1( u1_u12_u4_n99 ) );
  AOI21_X1 u1_u12_u4_U7 (.ZN( u1_u12_u4_n108 ) , .B2( u1_u12_u4_n134 ) , .B1( u1_u12_u4_n155 ) , .A( u1_u12_u4_n156 ) );
  NOR2_X1 u1_u12_u4_U70 (.A2( u1_u12_X_28 ) , .ZN( u1_u12_u4_n150 ) , .A1( u1_u12_u4_n168 ) );
  NOR2_X1 u1_u12_u4_U71 (.A2( u1_u12_X_29 ) , .ZN( u1_u12_u4_n152 ) , .A1( u1_u12_u4_n169 ) );
  NOR2_X1 u1_u12_u4_U72 (.A2( u1_u12_X_30 ) , .ZN( u1_u12_u4_n105 ) , .A1( u1_u12_u4_n176 ) );
  NOR2_X1 u1_u12_u4_U73 (.A2( u1_u12_X_26 ) , .ZN( u1_u12_u4_n100 ) , .A1( u1_u12_u4_n177 ) );
  NOR2_X1 u1_u12_u4_U74 (.A2( u1_u12_X_28 ) , .A1( u1_u12_X_29 ) , .ZN( u1_u12_u4_n128 ) );
  NOR2_X1 u1_u12_u4_U75 (.A2( u1_u12_X_27 ) , .A1( u1_u12_X_30 ) , .ZN( u1_u12_u4_n102 ) );
  NOR2_X1 u1_u12_u4_U76 (.A2( u1_u12_X_25 ) , .A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n98 ) );
  AND2_X1 u1_u12_u4_U77 (.A2( u1_u12_X_25 ) , .A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n104 ) );
  AND2_X1 u1_u12_u4_U78 (.A1( u1_u12_X_30 ) , .A2( u1_u12_u4_n176 ) , .ZN( u1_u12_u4_n99 ) );
  AND2_X1 u1_u12_u4_U79 (.A1( u1_u12_X_26 ) , .ZN( u1_u12_u4_n101 ) , .A2( u1_u12_u4_n177 ) );
  AOI21_X1 u1_u12_u4_U8 (.ZN( u1_u12_u4_n109 ) , .A( u1_u12_u4_n153 ) , .B1( u1_u12_u4_n159 ) , .B2( u1_u12_u4_n184 ) );
  AND2_X1 u1_u12_u4_U80 (.A1( u1_u12_X_27 ) , .A2( u1_u12_X_30 ) , .ZN( u1_u12_u4_n103 ) );
  INV_X1 u1_u12_u4_U81 (.A( u1_u12_X_28 ) , .ZN( u1_u12_u4_n169 ) );
  INV_X1 u1_u12_u4_U82 (.A( u1_u12_X_29 ) , .ZN( u1_u12_u4_n168 ) );
  INV_X1 u1_u12_u4_U83 (.A( u1_u12_X_25 ) , .ZN( u1_u12_u4_n177 ) );
  INV_X1 u1_u12_u4_U84 (.A( u1_u12_X_27 ) , .ZN( u1_u12_u4_n176 ) );
  NAND4_X1 u1_u12_u4_U85 (.ZN( u1_out12_25 ) , .A4( u1_u12_u4_n139 ) , .A3( u1_u12_u4_n140 ) , .A2( u1_u12_u4_n141 ) , .A1( u1_u12_u4_n142 ) );
  OAI21_X1 u1_u12_u4_U86 (.A( u1_u12_u4_n128 ) , .B2( u1_u12_u4_n129 ) , .B1( u1_u12_u4_n130 ) , .ZN( u1_u12_u4_n142 ) );
  OAI21_X1 u1_u12_u4_U87 (.B2( u1_u12_u4_n131 ) , .ZN( u1_u12_u4_n141 ) , .A( u1_u12_u4_n175 ) , .B1( u1_u12_u4_n183 ) );
  NAND4_X1 u1_u12_u4_U88 (.ZN( u1_out12_14 ) , .A4( u1_u12_u4_n124 ) , .A3( u1_u12_u4_n125 ) , .A2( u1_u12_u4_n126 ) , .A1( u1_u12_u4_n127 ) );
  AOI22_X1 u1_u12_u4_U89 (.B2( u1_u12_u4_n117 ) , .ZN( u1_u12_u4_n126 ) , .A1( u1_u12_u4_n129 ) , .B1( u1_u12_u4_n152 ) , .A2( u1_u12_u4_n175 ) );
  AOI211_X1 u1_u12_u4_U9 (.B( u1_u12_u4_n136 ) , .A( u1_u12_u4_n137 ) , .C2( u1_u12_u4_n138 ) , .ZN( u1_u12_u4_n139 ) , .C1( u1_u12_u4_n182 ) );
  AOI22_X1 u1_u12_u4_U90 (.ZN( u1_u12_u4_n125 ) , .B2( u1_u12_u4_n131 ) , .A2( u1_u12_u4_n132 ) , .B1( u1_u12_u4_n138 ) , .A1( u1_u12_u4_n178 ) );
  NAND4_X1 u1_u12_u4_U91 (.ZN( u1_out12_8 ) , .A4( u1_u12_u4_n110 ) , .A3( u1_u12_u4_n111 ) , .A2( u1_u12_u4_n112 ) , .A1( u1_u12_u4_n186 ) );
  NAND2_X1 u1_u12_u4_U92 (.ZN( u1_u12_u4_n112 ) , .A2( u1_u12_u4_n130 ) , .A1( u1_u12_u4_n150 ) );
  AOI22_X1 u1_u12_u4_U93 (.ZN( u1_u12_u4_n111 ) , .B2( u1_u12_u4_n132 ) , .A1( u1_u12_u4_n152 ) , .B1( u1_u12_u4_n178 ) , .A2( u1_u12_u4_n97 ) );
  AOI22_X1 u1_u12_u4_U94 (.B2( u1_u12_u4_n149 ) , .B1( u1_u12_u4_n150 ) , .A2( u1_u12_u4_n151 ) , .A1( u1_u12_u4_n152 ) , .ZN( u1_u12_u4_n167 ) );
  NOR4_X1 u1_u12_u4_U95 (.A4( u1_u12_u4_n162 ) , .A3( u1_u12_u4_n163 ) , .A2( u1_u12_u4_n164 ) , .A1( u1_u12_u4_n165 ) , .ZN( u1_u12_u4_n166 ) );
  NAND3_X1 u1_u12_u4_U96 (.ZN( u1_out12_3 ) , .A3( u1_u12_u4_n166 ) , .A1( u1_u12_u4_n167 ) , .A2( u1_u12_u4_n186 ) );
  NAND3_X1 u1_u12_u4_U97 (.A3( u1_u12_u4_n146 ) , .A2( u1_u12_u4_n147 ) , .A1( u1_u12_u4_n148 ) , .ZN( u1_u12_u4_n149 ) );
  NAND3_X1 u1_u12_u4_U98 (.A3( u1_u12_u4_n143 ) , .A2( u1_u12_u4_n144 ) , .A1( u1_u12_u4_n145 ) , .ZN( u1_u12_u4_n151 ) );
  NAND3_X1 u1_u12_u4_U99 (.A3( u1_u12_u4_n121 ) , .ZN( u1_u12_u4_n122 ) , .A2( u1_u12_u4_n144 ) , .A1( u1_u12_u4_n154 ) );
  XOR2_X1 u1_u13_U1 (.B( u1_K14_9 ) , .A( u1_R12_6 ) , .Z( u1_u13_X_9 ) );
  XOR2_X1 u1_u13_U10 (.B( u1_K14_45 ) , .A( u1_R12_30 ) , .Z( u1_u13_X_45 ) );
  XOR2_X1 u1_u13_U11 (.B( u1_K14_44 ) , .A( u1_R12_29 ) , .Z( u1_u13_X_44 ) );
  XOR2_X1 u1_u13_U12 (.B( u1_K14_43 ) , .A( u1_R12_28 ) , .Z( u1_u13_X_43 ) );
  XOR2_X1 u1_u13_U13 (.B( u1_K14_42 ) , .A( u1_R12_29 ) , .Z( u1_u13_X_42 ) );
  XOR2_X1 u1_u13_U14 (.B( u1_K14_41 ) , .A( u1_R12_28 ) , .Z( u1_u13_X_41 ) );
  XOR2_X1 u1_u13_U15 (.B( u1_K14_40 ) , .A( u1_R12_27 ) , .Z( u1_u13_X_40 ) );
  XOR2_X1 u1_u13_U17 (.B( u1_K14_39 ) , .A( u1_R12_26 ) , .Z( u1_u13_X_39 ) );
  XOR2_X1 u1_u13_U18 (.B( u1_K14_38 ) , .A( u1_R12_25 ) , .Z( u1_u13_X_38 ) );
  XOR2_X1 u1_u13_U19 (.B( u1_K14_37 ) , .A( u1_R12_24 ) , .Z( u1_u13_X_37 ) );
  XOR2_X1 u1_u13_U2 (.B( u1_K14_8 ) , .A( u1_R12_5 ) , .Z( u1_u13_X_8 ) );
  XOR2_X1 u1_u13_U20 (.B( u1_K14_36 ) , .A( u1_R12_25 ) , .Z( u1_u13_X_36 ) );
  XOR2_X1 u1_u13_U21 (.B( u1_K14_35 ) , .A( u1_R12_24 ) , .Z( u1_u13_X_35 ) );
  XOR2_X1 u1_u13_U24 (.B( u1_K14_32 ) , .A( u1_R12_21 ) , .Z( u1_u13_X_32 ) );
  XOR2_X1 u1_u13_U25 (.B( u1_K14_31 ) , .A( u1_R12_20 ) , .Z( u1_u13_X_31 ) );
  XOR2_X1 u1_u13_U26 (.B( u1_K14_30 ) , .A( u1_R12_21 ) , .Z( u1_u13_X_30 ) );
  XOR2_X1 u1_u13_U27 (.B( u1_K14_2 ) , .A( u1_R12_1 ) , .Z( u1_u13_X_2 ) );
  XOR2_X1 u1_u13_U28 (.B( u1_K14_29 ) , .A( u1_R12_20 ) , .Z( u1_u13_X_29 ) );
  XOR2_X1 u1_u13_U29 (.B( u1_K14_28 ) , .A( u1_R12_19 ) , .Z( u1_u13_X_28 ) );
  XOR2_X1 u1_u13_U3 (.B( u1_K14_7 ) , .A( u1_R12_4 ) , .Z( u1_u13_X_7 ) );
  XOR2_X1 u1_u13_U30 (.B( u1_K14_27 ) , .A( u1_R12_18 ) , .Z( u1_u13_X_27 ) );
  XOR2_X1 u1_u13_U31 (.B( u1_K14_26 ) , .A( u1_R12_17 ) , .Z( u1_u13_X_26 ) );
  XOR2_X1 u1_u13_U32 (.B( u1_K14_25 ) , .A( u1_R12_16 ) , .Z( u1_u13_X_25 ) );
  XOR2_X1 u1_u13_U33 (.B( u1_K14_24 ) , .A( u1_R12_17 ) , .Z( u1_u13_X_24 ) );
  XOR2_X1 u1_u13_U34 (.B( u1_K14_23 ) , .A( u1_R12_16 ) , .Z( u1_u13_X_23 ) );
  XOR2_X1 u1_u13_U37 (.B( u1_K14_20 ) , .A( u1_R12_13 ) , .Z( u1_u13_X_20 ) );
  XOR2_X1 u1_u13_U38 (.B( u1_K14_1 ) , .A( u1_R12_32 ) , .Z( u1_u13_X_1 ) );
  XOR2_X1 u1_u13_U39 (.B( u1_K14_19 ) , .A( u1_R12_12 ) , .Z( u1_u13_X_19 ) );
  XOR2_X1 u1_u13_U4 (.B( u1_K14_6 ) , .A( u1_R12_5 ) , .Z( u1_u13_X_6 ) );
  XOR2_X1 u1_u13_U40 (.B( u1_K14_18 ) , .A( u1_R12_13 ) , .Z( u1_u13_X_18 ) );
  XOR2_X1 u1_u13_U41 (.B( u1_K14_17 ) , .A( u1_R12_12 ) , .Z( u1_u13_X_17 ) );
  XOR2_X1 u1_u13_U44 (.B( u1_K14_14 ) , .A( u1_R12_9 ) , .Z( u1_u13_X_14 ) );
  XOR2_X1 u1_u13_U45 (.B( u1_K14_13 ) , .A( u1_R12_8 ) , .Z( u1_u13_X_13 ) );
  XOR2_X1 u1_u13_U46 (.B( u1_K14_12 ) , .A( u1_R12_9 ) , .Z( u1_u13_X_12 ) );
  XOR2_X1 u1_u13_U47 (.B( u1_K14_11 ) , .A( u1_R12_8 ) , .Z( u1_u13_X_11 ) );
  XOR2_X1 u1_u13_U48 (.B( u1_K14_10 ) , .A( u1_R12_7 ) , .Z( u1_u13_X_10 ) );
  XOR2_X1 u1_u13_U5 (.B( u1_K14_5 ) , .A( u1_R12_4 ) , .Z( u1_u13_X_5 ) );
  XOR2_X1 u1_u13_U7 (.B( u1_K14_48 ) , .A( u1_R12_1 ) , .Z( u1_u13_X_48 ) );
  XOR2_X1 u1_u13_U8 (.B( u1_K14_47 ) , .A( u1_R12_32 ) , .Z( u1_u13_X_47 ) );
  XOR2_X1 u1_u13_U9 (.B( u1_K14_46 ) , .A( u1_R12_31 ) , .Z( u1_u13_X_46 ) );
  NAND2_X1 u1_u13_u1_U10 (.A1( u1_u13_u1_n131 ) , .ZN( u1_u13_u1_n147 ) , .A2( u1_u13_u1_n153 ) );
  NAND3_X1 u1_u13_u1_U100 (.ZN( u1_u13_u1_n113 ) , .A1( u1_u13_u1_n120 ) , .A3( u1_u13_u1_n133 ) , .A2( u1_u13_u1_n155 ) );
  AOI22_X1 u1_u13_u1_U11 (.B2( u1_u13_u1_n136 ) , .A2( u1_u13_u1_n137 ) , .ZN( u1_u13_u1_n143 ) , .A1( u1_u13_u1_n171 ) , .B1( u1_u13_u1_n173 ) );
  INV_X1 u1_u13_u1_U12 (.A( u1_u13_u1_n147 ) , .ZN( u1_u13_u1_n181 ) );
  INV_X1 u1_u13_u1_U13 (.A( u1_u13_u1_n139 ) , .ZN( u1_u13_u1_n174 ) );
  OR4_X1 u1_u13_u1_U14 (.A4( u1_u13_u1_n106 ) , .A3( u1_u13_u1_n107 ) , .ZN( u1_u13_u1_n108 ) , .A1( u1_u13_u1_n117 ) , .A2( u1_u13_u1_n184 ) );
  AOI21_X1 u1_u13_u1_U15 (.ZN( u1_u13_u1_n106 ) , .A( u1_u13_u1_n112 ) , .B1( u1_u13_u1_n154 ) , .B2( u1_u13_u1_n156 ) );
  AOI21_X1 u1_u13_u1_U16 (.ZN( u1_u13_u1_n107 ) , .B1( u1_u13_u1_n134 ) , .B2( u1_u13_u1_n149 ) , .A( u1_u13_u1_n174 ) );
  INV_X1 u1_u13_u1_U17 (.A( u1_u13_u1_n101 ) , .ZN( u1_u13_u1_n184 ) );
  INV_X1 u1_u13_u1_U18 (.A( u1_u13_u1_n112 ) , .ZN( u1_u13_u1_n171 ) );
  NAND2_X1 u1_u13_u1_U19 (.ZN( u1_u13_u1_n141 ) , .A1( u1_u13_u1_n153 ) , .A2( u1_u13_u1_n156 ) );
  AND2_X1 u1_u13_u1_U20 (.A1( u1_u13_u1_n123 ) , .ZN( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n161 ) );
  NAND2_X1 u1_u13_u1_U21 (.A2( u1_u13_u1_n115 ) , .A1( u1_u13_u1_n116 ) , .ZN( u1_u13_u1_n148 ) );
  NAND2_X1 u1_u13_u1_U22 (.A2( u1_u13_u1_n133 ) , .A1( u1_u13_u1_n135 ) , .ZN( u1_u13_u1_n159 ) );
  NAND2_X1 u1_u13_u1_U23 (.A2( u1_u13_u1_n115 ) , .A1( u1_u13_u1_n120 ) , .ZN( u1_u13_u1_n132 ) );
  INV_X1 u1_u13_u1_U24 (.A( u1_u13_u1_n154 ) , .ZN( u1_u13_u1_n178 ) );
  AOI22_X1 u1_u13_u1_U25 (.B2( u1_u13_u1_n113 ) , .A2( u1_u13_u1_n114 ) , .ZN( u1_u13_u1_n125 ) , .A1( u1_u13_u1_n171 ) , .B1( u1_u13_u1_n173 ) );
  NAND2_X1 u1_u13_u1_U26 (.ZN( u1_u13_u1_n114 ) , .A1( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n156 ) );
  INV_X1 u1_u13_u1_U27 (.A( u1_u13_u1_n151 ) , .ZN( u1_u13_u1_n183 ) );
  AND2_X1 u1_u13_u1_U28 (.A1( u1_u13_u1_n129 ) , .A2( u1_u13_u1_n133 ) , .ZN( u1_u13_u1_n149 ) );
  INV_X1 u1_u13_u1_U29 (.A( u1_u13_u1_n131 ) , .ZN( u1_u13_u1_n180 ) );
  INV_X1 u1_u13_u1_U3 (.A( u1_u13_u1_n159 ) , .ZN( u1_u13_u1_n182 ) );
  OAI221_X1 u1_u13_u1_U30 (.A( u1_u13_u1_n119 ) , .C2( u1_u13_u1_n129 ) , .ZN( u1_u13_u1_n138 ) , .B2( u1_u13_u1_n152 ) , .C1( u1_u13_u1_n174 ) , .B1( u1_u13_u1_n187 ) );
  INV_X1 u1_u13_u1_U31 (.A( u1_u13_u1_n148 ) , .ZN( u1_u13_u1_n187 ) );
  AOI211_X1 u1_u13_u1_U32 (.B( u1_u13_u1_n117 ) , .A( u1_u13_u1_n118 ) , .ZN( u1_u13_u1_n119 ) , .C2( u1_u13_u1_n146 ) , .C1( u1_u13_u1_n159 ) );
  NOR2_X1 u1_u13_u1_U33 (.A1( u1_u13_u1_n168 ) , .A2( u1_u13_u1_n176 ) , .ZN( u1_u13_u1_n98 ) );
  AOI211_X1 u1_u13_u1_U34 (.B( u1_u13_u1_n162 ) , .A( u1_u13_u1_n163 ) , .C2( u1_u13_u1_n164 ) , .ZN( u1_u13_u1_n165 ) , .C1( u1_u13_u1_n171 ) );
  AOI21_X1 u1_u13_u1_U35 (.A( u1_u13_u1_n160 ) , .B2( u1_u13_u1_n161 ) , .ZN( u1_u13_u1_n162 ) , .B1( u1_u13_u1_n182 ) );
  OR2_X1 u1_u13_u1_U36 (.A2( u1_u13_u1_n157 ) , .A1( u1_u13_u1_n158 ) , .ZN( u1_u13_u1_n163 ) );
  OAI21_X1 u1_u13_u1_U37 (.B2( u1_u13_u1_n123 ) , .ZN( u1_u13_u1_n145 ) , .B1( u1_u13_u1_n160 ) , .A( u1_u13_u1_n185 ) );
  INV_X1 u1_u13_u1_U38 (.A( u1_u13_u1_n122 ) , .ZN( u1_u13_u1_n185 ) );
  AOI21_X1 u1_u13_u1_U39 (.B2( u1_u13_u1_n120 ) , .B1( u1_u13_u1_n121 ) , .ZN( u1_u13_u1_n122 ) , .A( u1_u13_u1_n128 ) );
  AOI221_X1 u1_u13_u1_U4 (.A( u1_u13_u1_n138 ) , .C2( u1_u13_u1_n139 ) , .C1( u1_u13_u1_n140 ) , .B2( u1_u13_u1_n141 ) , .ZN( u1_u13_u1_n142 ) , .B1( u1_u13_u1_n175 ) );
  NAND2_X1 u1_u13_u1_U40 (.A1( u1_u13_u1_n128 ) , .ZN( u1_u13_u1_n146 ) , .A2( u1_u13_u1_n160 ) );
  NAND2_X1 u1_u13_u1_U41 (.A2( u1_u13_u1_n112 ) , .ZN( u1_u13_u1_n139 ) , .A1( u1_u13_u1_n152 ) );
  NAND2_X1 u1_u13_u1_U42 (.A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n156 ) , .A2( u1_u13_u1_n99 ) );
  AOI221_X1 u1_u13_u1_U43 (.B1( u1_u13_u1_n140 ) , .ZN( u1_u13_u1_n167 ) , .B2( u1_u13_u1_n172 ) , .C2( u1_u13_u1_n175 ) , .C1( u1_u13_u1_n178 ) , .A( u1_u13_u1_n188 ) );
  INV_X1 u1_u13_u1_U44 (.ZN( u1_u13_u1_n188 ) , .A( u1_u13_u1_n97 ) );
  AOI211_X1 u1_u13_u1_U45 (.A( u1_u13_u1_n118 ) , .C1( u1_u13_u1_n132 ) , .C2( u1_u13_u1_n139 ) , .B( u1_u13_u1_n96 ) , .ZN( u1_u13_u1_n97 ) );
  AOI21_X1 u1_u13_u1_U46 (.B2( u1_u13_u1_n121 ) , .B1( u1_u13_u1_n135 ) , .A( u1_u13_u1_n152 ) , .ZN( u1_u13_u1_n96 ) );
  NOR2_X1 u1_u13_u1_U47 (.ZN( u1_u13_u1_n117 ) , .A1( u1_u13_u1_n121 ) , .A2( u1_u13_u1_n160 ) );
  AOI21_X1 u1_u13_u1_U48 (.A( u1_u13_u1_n128 ) , .B2( u1_u13_u1_n129 ) , .ZN( u1_u13_u1_n130 ) , .B1( u1_u13_u1_n150 ) );
  NAND2_X1 u1_u13_u1_U49 (.ZN( u1_u13_u1_n112 ) , .A1( u1_u13_u1_n169 ) , .A2( u1_u13_u1_n170 ) );
  AOI211_X1 u1_u13_u1_U5 (.ZN( u1_u13_u1_n124 ) , .A( u1_u13_u1_n138 ) , .C2( u1_u13_u1_n139 ) , .B( u1_u13_u1_n145 ) , .C1( u1_u13_u1_n147 ) );
  NAND2_X1 u1_u13_u1_U50 (.ZN( u1_u13_u1_n129 ) , .A2( u1_u13_u1_n95 ) , .A1( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U51 (.A1( u1_u13_u1_n102 ) , .ZN( u1_u13_u1_n154 ) , .A2( u1_u13_u1_n99 ) );
  NAND2_X1 u1_u13_u1_U52 (.A2( u1_u13_u1_n100 ) , .ZN( u1_u13_u1_n135 ) , .A1( u1_u13_u1_n99 ) );
  AOI21_X1 u1_u13_u1_U53 (.A( u1_u13_u1_n152 ) , .B2( u1_u13_u1_n153 ) , .B1( u1_u13_u1_n154 ) , .ZN( u1_u13_u1_n158 ) );
  INV_X1 u1_u13_u1_U54 (.A( u1_u13_u1_n160 ) , .ZN( u1_u13_u1_n175 ) );
  NAND2_X1 u1_u13_u1_U55 (.A1( u1_u13_u1_n100 ) , .ZN( u1_u13_u1_n116 ) , .A2( u1_u13_u1_n95 ) );
  NAND2_X1 u1_u13_u1_U56 (.A1( u1_u13_u1_n102 ) , .ZN( u1_u13_u1_n131 ) , .A2( u1_u13_u1_n95 ) );
  NAND2_X1 u1_u13_u1_U57 (.A2( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n121 ) , .A1( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U58 (.A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n153 ) , .A2( u1_u13_u1_n98 ) );
  NAND2_X1 u1_u13_u1_U59 (.A2( u1_u13_u1_n104 ) , .A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n133 ) );
  NOR2_X1 u1_u13_u1_U6 (.A1( u1_u13_u1_n112 ) , .A2( u1_u13_u1_n116 ) , .ZN( u1_u13_u1_n118 ) );
  NAND2_X1 u1_u13_u1_U60 (.ZN( u1_u13_u1_n150 ) , .A2( u1_u13_u1_n98 ) , .A1( u1_u13_u1_n99 ) );
  NAND2_X1 u1_u13_u1_U61 (.A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n155 ) , .A2( u1_u13_u1_n95 ) );
  OAI21_X1 u1_u13_u1_U62 (.ZN( u1_u13_u1_n109 ) , .B1( u1_u13_u1_n129 ) , .B2( u1_u13_u1_n160 ) , .A( u1_u13_u1_n167 ) );
  NAND2_X1 u1_u13_u1_U63 (.A2( u1_u13_u1_n100 ) , .A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n120 ) );
  NAND2_X1 u1_u13_u1_U64 (.A1( u1_u13_u1_n102 ) , .A2( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n115 ) );
  NAND2_X1 u1_u13_u1_U65 (.A2( u1_u13_u1_n100 ) , .A1( u1_u13_u1_n104 ) , .ZN( u1_u13_u1_n151 ) );
  NAND2_X1 u1_u13_u1_U66 (.A2( u1_u13_u1_n103 ) , .A1( u1_u13_u1_n105 ) , .ZN( u1_u13_u1_n161 ) );
  INV_X1 u1_u13_u1_U67 (.A( u1_u13_u1_n152 ) , .ZN( u1_u13_u1_n173 ) );
  INV_X1 u1_u13_u1_U68 (.A( u1_u13_u1_n128 ) , .ZN( u1_u13_u1_n172 ) );
  NAND2_X1 u1_u13_u1_U69 (.A2( u1_u13_u1_n102 ) , .A1( u1_u13_u1_n103 ) , .ZN( u1_u13_u1_n123 ) );
  OAI21_X1 u1_u13_u1_U7 (.ZN( u1_u13_u1_n101 ) , .B1( u1_u13_u1_n141 ) , .A( u1_u13_u1_n146 ) , .B2( u1_u13_u1_n183 ) );
  NOR2_X1 u1_u13_u1_U70 (.A2( u1_u13_X_7 ) , .A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n95 ) );
  NOR2_X1 u1_u13_u1_U71 (.A1( u1_u13_X_12 ) , .A2( u1_u13_X_9 ) , .ZN( u1_u13_u1_n100 ) );
  NOR2_X1 u1_u13_u1_U72 (.A2( u1_u13_X_8 ) , .A1( u1_u13_u1_n177 ) , .ZN( u1_u13_u1_n99 ) );
  NOR2_X1 u1_u13_u1_U73 (.A2( u1_u13_X_12 ) , .ZN( u1_u13_u1_n102 ) , .A1( u1_u13_u1_n176 ) );
  NOR2_X1 u1_u13_u1_U74 (.A2( u1_u13_X_9 ) , .ZN( u1_u13_u1_n105 ) , .A1( u1_u13_u1_n168 ) );
  NAND2_X1 u1_u13_u1_U75 (.A1( u1_u13_X_10 ) , .ZN( u1_u13_u1_n160 ) , .A2( u1_u13_u1_n169 ) );
  NAND2_X1 u1_u13_u1_U76 (.A2( u1_u13_X_10 ) , .A1( u1_u13_X_11 ) , .ZN( u1_u13_u1_n152 ) );
  NAND2_X1 u1_u13_u1_U77 (.A1( u1_u13_X_11 ) , .ZN( u1_u13_u1_n128 ) , .A2( u1_u13_u1_n170 ) );
  AND2_X1 u1_u13_u1_U78 (.A2( u1_u13_X_7 ) , .A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n104 ) );
  AND2_X1 u1_u13_u1_U79 (.A1( u1_u13_X_8 ) , .ZN( u1_u13_u1_n103 ) , .A2( u1_u13_u1_n177 ) );
  AOI21_X1 u1_u13_u1_U8 (.B2( u1_u13_u1_n155 ) , .B1( u1_u13_u1_n156 ) , .ZN( u1_u13_u1_n157 ) , .A( u1_u13_u1_n174 ) );
  INV_X1 u1_u13_u1_U80 (.A( u1_u13_X_10 ) , .ZN( u1_u13_u1_n170 ) );
  INV_X1 u1_u13_u1_U81 (.A( u1_u13_X_9 ) , .ZN( u1_u13_u1_n176 ) );
  INV_X1 u1_u13_u1_U82 (.A( u1_u13_X_11 ) , .ZN( u1_u13_u1_n169 ) );
  INV_X1 u1_u13_u1_U83 (.A( u1_u13_X_12 ) , .ZN( u1_u13_u1_n168 ) );
  INV_X1 u1_u13_u1_U84 (.A( u1_u13_X_7 ) , .ZN( u1_u13_u1_n177 ) );
  NAND4_X1 u1_u13_u1_U85 (.ZN( u1_out13_18 ) , .A4( u1_u13_u1_n165 ) , .A3( u1_u13_u1_n166 ) , .A1( u1_u13_u1_n167 ) , .A2( u1_u13_u1_n186 ) );
  AOI22_X1 u1_u13_u1_U86 (.B2( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n147 ) , .A2( u1_u13_u1_n148 ) , .ZN( u1_u13_u1_n166 ) , .A1( u1_u13_u1_n172 ) );
  INV_X1 u1_u13_u1_U87 (.A( u1_u13_u1_n145 ) , .ZN( u1_u13_u1_n186 ) );
  NAND4_X1 u1_u13_u1_U88 (.ZN( u1_out13_2 ) , .A4( u1_u13_u1_n142 ) , .A3( u1_u13_u1_n143 ) , .A2( u1_u13_u1_n144 ) , .A1( u1_u13_u1_n179 ) );
  OAI21_X1 u1_u13_u1_U89 (.B2( u1_u13_u1_n132 ) , .ZN( u1_u13_u1_n144 ) , .A( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n180 ) );
  NAND2_X1 u1_u13_u1_U9 (.ZN( u1_u13_u1_n140 ) , .A2( u1_u13_u1_n150 ) , .A1( u1_u13_u1_n155 ) );
  INV_X1 u1_u13_u1_U90 (.A( u1_u13_u1_n130 ) , .ZN( u1_u13_u1_n179 ) );
  NAND4_X1 u1_u13_u1_U91 (.ZN( u1_out13_28 ) , .A4( u1_u13_u1_n124 ) , .A3( u1_u13_u1_n125 ) , .A2( u1_u13_u1_n126 ) , .A1( u1_u13_u1_n127 ) );
  OAI21_X1 u1_u13_u1_U92 (.ZN( u1_u13_u1_n127 ) , .B2( u1_u13_u1_n139 ) , .B1( u1_u13_u1_n175 ) , .A( u1_u13_u1_n183 ) );
  OAI21_X1 u1_u13_u1_U93 (.ZN( u1_u13_u1_n126 ) , .B2( u1_u13_u1_n140 ) , .A( u1_u13_u1_n146 ) , .B1( u1_u13_u1_n178 ) );
  OR4_X1 u1_u13_u1_U94 (.ZN( u1_out13_13 ) , .A4( u1_u13_u1_n108 ) , .A3( u1_u13_u1_n109 ) , .A2( u1_u13_u1_n110 ) , .A1( u1_u13_u1_n111 ) );
  AOI21_X1 u1_u13_u1_U95 (.ZN( u1_u13_u1_n111 ) , .A( u1_u13_u1_n128 ) , .B2( u1_u13_u1_n131 ) , .B1( u1_u13_u1_n135 ) );
  AOI21_X1 u1_u13_u1_U96 (.ZN( u1_u13_u1_n110 ) , .A( u1_u13_u1_n116 ) , .B1( u1_u13_u1_n152 ) , .B2( u1_u13_u1_n160 ) );
  NAND3_X1 u1_u13_u1_U97 (.A3( u1_u13_u1_n149 ) , .A2( u1_u13_u1_n150 ) , .A1( u1_u13_u1_n151 ) , .ZN( u1_u13_u1_n164 ) );
  NAND3_X1 u1_u13_u1_U98 (.A3( u1_u13_u1_n134 ) , .A2( u1_u13_u1_n135 ) , .ZN( u1_u13_u1_n136 ) , .A1( u1_u13_u1_n151 ) );
  NAND3_X1 u1_u13_u1_U99 (.A1( u1_u13_u1_n133 ) , .ZN( u1_u13_u1_n137 ) , .A2( u1_u13_u1_n154 ) , .A3( u1_u13_u1_n181 ) );
  OAI22_X1 u1_u13_u4_U10 (.B2( u1_u13_u4_n135 ) , .ZN( u1_u13_u4_n137 ) , .B1( u1_u13_u4_n153 ) , .A1( u1_u13_u4_n155 ) , .A2( u1_u13_u4_n171 ) );
  AND3_X1 u1_u13_u4_U11 (.A2( u1_u13_u4_n134 ) , .ZN( u1_u13_u4_n135 ) , .A3( u1_u13_u4_n145 ) , .A1( u1_u13_u4_n157 ) );
  NAND2_X1 u1_u13_u4_U12 (.ZN( u1_u13_u4_n132 ) , .A2( u1_u13_u4_n170 ) , .A1( u1_u13_u4_n173 ) );
  AOI21_X1 u1_u13_u4_U13 (.B2( u1_u13_u4_n160 ) , .B1( u1_u13_u4_n161 ) , .ZN( u1_u13_u4_n162 ) , .A( u1_u13_u4_n170 ) );
  AOI21_X1 u1_u13_u4_U14 (.ZN( u1_u13_u4_n107 ) , .B2( u1_u13_u4_n143 ) , .A( u1_u13_u4_n174 ) , .B1( u1_u13_u4_n184 ) );
  AOI21_X1 u1_u13_u4_U15 (.B2( u1_u13_u4_n158 ) , .B1( u1_u13_u4_n159 ) , .ZN( u1_u13_u4_n163 ) , .A( u1_u13_u4_n174 ) );
  AOI21_X1 u1_u13_u4_U16 (.A( u1_u13_u4_n153 ) , .B2( u1_u13_u4_n154 ) , .B1( u1_u13_u4_n155 ) , .ZN( u1_u13_u4_n165 ) );
  AOI21_X1 u1_u13_u4_U17 (.A( u1_u13_u4_n156 ) , .B2( u1_u13_u4_n157 ) , .ZN( u1_u13_u4_n164 ) , .B1( u1_u13_u4_n184 ) );
  INV_X1 u1_u13_u4_U18 (.A( u1_u13_u4_n138 ) , .ZN( u1_u13_u4_n170 ) );
  AND2_X1 u1_u13_u4_U19 (.A2( u1_u13_u4_n120 ) , .ZN( u1_u13_u4_n155 ) , .A1( u1_u13_u4_n160 ) );
  INV_X1 u1_u13_u4_U20 (.A( u1_u13_u4_n156 ) , .ZN( u1_u13_u4_n175 ) );
  NAND2_X1 u1_u13_u4_U21 (.A2( u1_u13_u4_n118 ) , .ZN( u1_u13_u4_n131 ) , .A1( u1_u13_u4_n147 ) );
  NAND2_X1 u1_u13_u4_U22 (.A1( u1_u13_u4_n119 ) , .A2( u1_u13_u4_n120 ) , .ZN( u1_u13_u4_n130 ) );
  NAND2_X1 u1_u13_u4_U23 (.ZN( u1_u13_u4_n117 ) , .A2( u1_u13_u4_n118 ) , .A1( u1_u13_u4_n148 ) );
  NAND2_X1 u1_u13_u4_U24 (.ZN( u1_u13_u4_n129 ) , .A1( u1_u13_u4_n134 ) , .A2( u1_u13_u4_n148 ) );
  AND3_X1 u1_u13_u4_U25 (.A1( u1_u13_u4_n119 ) , .A2( u1_u13_u4_n143 ) , .A3( u1_u13_u4_n154 ) , .ZN( u1_u13_u4_n161 ) );
  AND2_X1 u1_u13_u4_U26 (.A1( u1_u13_u4_n145 ) , .A2( u1_u13_u4_n147 ) , .ZN( u1_u13_u4_n159 ) );
  OR3_X1 u1_u13_u4_U27 (.A3( u1_u13_u4_n114 ) , .A2( u1_u13_u4_n115 ) , .A1( u1_u13_u4_n116 ) , .ZN( u1_u13_u4_n136 ) );
  AOI21_X1 u1_u13_u4_U28 (.A( u1_u13_u4_n113 ) , .ZN( u1_u13_u4_n116 ) , .B2( u1_u13_u4_n173 ) , .B1( u1_u13_u4_n174 ) );
  AOI21_X1 u1_u13_u4_U29 (.ZN( u1_u13_u4_n115 ) , .B2( u1_u13_u4_n145 ) , .B1( u1_u13_u4_n146 ) , .A( u1_u13_u4_n156 ) );
  NOR2_X1 u1_u13_u4_U3 (.ZN( u1_u13_u4_n121 ) , .A1( u1_u13_u4_n181 ) , .A2( u1_u13_u4_n182 ) );
  OAI22_X1 u1_u13_u4_U30 (.ZN( u1_u13_u4_n114 ) , .A2( u1_u13_u4_n121 ) , .B1( u1_u13_u4_n160 ) , .B2( u1_u13_u4_n170 ) , .A1( u1_u13_u4_n171 ) );
  INV_X1 u1_u13_u4_U31 (.A( u1_u13_u4_n158 ) , .ZN( u1_u13_u4_n182 ) );
  INV_X1 u1_u13_u4_U32 (.ZN( u1_u13_u4_n181 ) , .A( u1_u13_u4_n96 ) );
  INV_X1 u1_u13_u4_U33 (.A( u1_u13_u4_n144 ) , .ZN( u1_u13_u4_n179 ) );
  INV_X1 u1_u13_u4_U34 (.A( u1_u13_u4_n157 ) , .ZN( u1_u13_u4_n178 ) );
  NAND2_X1 u1_u13_u4_U35 (.A2( u1_u13_u4_n154 ) , .A1( u1_u13_u4_n96 ) , .ZN( u1_u13_u4_n97 ) );
  INV_X1 u1_u13_u4_U36 (.ZN( u1_u13_u4_n186 ) , .A( u1_u13_u4_n95 ) );
  OAI221_X1 u1_u13_u4_U37 (.C1( u1_u13_u4_n134 ) , .B1( u1_u13_u4_n158 ) , .B2( u1_u13_u4_n171 ) , .C2( u1_u13_u4_n173 ) , .A( u1_u13_u4_n94 ) , .ZN( u1_u13_u4_n95 ) );
  AOI222_X1 u1_u13_u4_U38 (.B2( u1_u13_u4_n132 ) , .A1( u1_u13_u4_n138 ) , .C2( u1_u13_u4_n175 ) , .A2( u1_u13_u4_n179 ) , .C1( u1_u13_u4_n181 ) , .B1( u1_u13_u4_n185 ) , .ZN( u1_u13_u4_n94 ) );
  INV_X1 u1_u13_u4_U39 (.A( u1_u13_u4_n113 ) , .ZN( u1_u13_u4_n185 ) );
  INV_X1 u1_u13_u4_U4 (.A( u1_u13_u4_n117 ) , .ZN( u1_u13_u4_n184 ) );
  INV_X1 u1_u13_u4_U40 (.A( u1_u13_u4_n143 ) , .ZN( u1_u13_u4_n183 ) );
  NOR2_X1 u1_u13_u4_U41 (.ZN( u1_u13_u4_n138 ) , .A1( u1_u13_u4_n168 ) , .A2( u1_u13_u4_n169 ) );
  NOR2_X1 u1_u13_u4_U42 (.A1( u1_u13_u4_n150 ) , .A2( u1_u13_u4_n152 ) , .ZN( u1_u13_u4_n153 ) );
  NOR2_X1 u1_u13_u4_U43 (.A2( u1_u13_u4_n128 ) , .A1( u1_u13_u4_n138 ) , .ZN( u1_u13_u4_n156 ) );
  AOI22_X1 u1_u13_u4_U44 (.B2( u1_u13_u4_n122 ) , .A1( u1_u13_u4_n123 ) , .ZN( u1_u13_u4_n124 ) , .B1( u1_u13_u4_n128 ) , .A2( u1_u13_u4_n172 ) );
  NAND2_X1 u1_u13_u4_U45 (.A2( u1_u13_u4_n120 ) , .ZN( u1_u13_u4_n123 ) , .A1( u1_u13_u4_n161 ) );
  INV_X1 u1_u13_u4_U46 (.A( u1_u13_u4_n153 ) , .ZN( u1_u13_u4_n172 ) );
  AOI22_X1 u1_u13_u4_U47 (.B2( u1_u13_u4_n132 ) , .A2( u1_u13_u4_n133 ) , .ZN( u1_u13_u4_n140 ) , .A1( u1_u13_u4_n150 ) , .B1( u1_u13_u4_n179 ) );
  NAND2_X1 u1_u13_u4_U48 (.ZN( u1_u13_u4_n133 ) , .A2( u1_u13_u4_n146 ) , .A1( u1_u13_u4_n154 ) );
  NAND2_X1 u1_u13_u4_U49 (.A1( u1_u13_u4_n103 ) , .ZN( u1_u13_u4_n154 ) , .A2( u1_u13_u4_n98 ) );
  NOR4_X1 u1_u13_u4_U5 (.A4( u1_u13_u4_n106 ) , .A3( u1_u13_u4_n107 ) , .A2( u1_u13_u4_n108 ) , .A1( u1_u13_u4_n109 ) , .ZN( u1_u13_u4_n110 ) );
  NAND2_X1 u1_u13_u4_U50 (.A1( u1_u13_u4_n101 ) , .ZN( u1_u13_u4_n158 ) , .A2( u1_u13_u4_n99 ) );
  AOI21_X1 u1_u13_u4_U51 (.ZN( u1_u13_u4_n127 ) , .A( u1_u13_u4_n136 ) , .B2( u1_u13_u4_n150 ) , .B1( u1_u13_u4_n180 ) );
  INV_X1 u1_u13_u4_U52 (.A( u1_u13_u4_n160 ) , .ZN( u1_u13_u4_n180 ) );
  NAND2_X1 u1_u13_u4_U53 (.A2( u1_u13_u4_n104 ) , .A1( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n146 ) );
  NAND2_X1 u1_u13_u4_U54 (.A2( u1_u13_u4_n101 ) , .A1( u1_u13_u4_n102 ) , .ZN( u1_u13_u4_n160 ) );
  NAND2_X1 u1_u13_u4_U55 (.ZN( u1_u13_u4_n134 ) , .A1( u1_u13_u4_n98 ) , .A2( u1_u13_u4_n99 ) );
  NAND2_X1 u1_u13_u4_U56 (.A1( u1_u13_u4_n103 ) , .A2( u1_u13_u4_n104 ) , .ZN( u1_u13_u4_n143 ) );
  NAND2_X1 u1_u13_u4_U57 (.A2( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n145 ) , .A1( u1_u13_u4_n98 ) );
  NAND2_X1 u1_u13_u4_U58 (.A1( u1_u13_u4_n100 ) , .A2( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n120 ) );
  NAND2_X1 u1_u13_u4_U59 (.A1( u1_u13_u4_n102 ) , .A2( u1_u13_u4_n104 ) , .ZN( u1_u13_u4_n148 ) );
  AOI21_X1 u1_u13_u4_U6 (.ZN( u1_u13_u4_n106 ) , .B2( u1_u13_u4_n146 ) , .B1( u1_u13_u4_n158 ) , .A( u1_u13_u4_n170 ) );
  NAND2_X1 u1_u13_u4_U60 (.A2( u1_u13_u4_n100 ) , .A1( u1_u13_u4_n103 ) , .ZN( u1_u13_u4_n157 ) );
  INV_X1 u1_u13_u4_U61 (.A( u1_u13_u4_n150 ) , .ZN( u1_u13_u4_n173 ) );
  INV_X1 u1_u13_u4_U62 (.A( u1_u13_u4_n152 ) , .ZN( u1_u13_u4_n171 ) );
  NAND2_X1 u1_u13_u4_U63 (.A1( u1_u13_u4_n100 ) , .ZN( u1_u13_u4_n118 ) , .A2( u1_u13_u4_n99 ) );
  NAND2_X1 u1_u13_u4_U64 (.A2( u1_u13_u4_n100 ) , .A1( u1_u13_u4_n102 ) , .ZN( u1_u13_u4_n144 ) );
  NAND2_X1 u1_u13_u4_U65 (.A2( u1_u13_u4_n101 ) , .A1( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n96 ) );
  INV_X1 u1_u13_u4_U66 (.A( u1_u13_u4_n128 ) , .ZN( u1_u13_u4_n174 ) );
  NAND2_X1 u1_u13_u4_U67 (.A2( u1_u13_u4_n102 ) , .ZN( u1_u13_u4_n119 ) , .A1( u1_u13_u4_n98 ) );
  NAND2_X1 u1_u13_u4_U68 (.A2( u1_u13_u4_n101 ) , .A1( u1_u13_u4_n103 ) , .ZN( u1_u13_u4_n147 ) );
  NAND2_X1 u1_u13_u4_U69 (.A2( u1_u13_u4_n104 ) , .ZN( u1_u13_u4_n113 ) , .A1( u1_u13_u4_n99 ) );
  AOI21_X1 u1_u13_u4_U7 (.ZN( u1_u13_u4_n108 ) , .B2( u1_u13_u4_n134 ) , .B1( u1_u13_u4_n155 ) , .A( u1_u13_u4_n156 ) );
  NOR2_X1 u1_u13_u4_U70 (.A2( u1_u13_X_28 ) , .ZN( u1_u13_u4_n150 ) , .A1( u1_u13_u4_n168 ) );
  NOR2_X1 u1_u13_u4_U71 (.A2( u1_u13_X_29 ) , .ZN( u1_u13_u4_n152 ) , .A1( u1_u13_u4_n169 ) );
  NOR2_X1 u1_u13_u4_U72 (.A2( u1_u13_X_30 ) , .ZN( u1_u13_u4_n105 ) , .A1( u1_u13_u4_n176 ) );
  NOR2_X1 u1_u13_u4_U73 (.A2( u1_u13_X_26 ) , .ZN( u1_u13_u4_n100 ) , .A1( u1_u13_u4_n177 ) );
  NOR2_X1 u1_u13_u4_U74 (.A2( u1_u13_X_28 ) , .A1( u1_u13_X_29 ) , .ZN( u1_u13_u4_n128 ) );
  NOR2_X1 u1_u13_u4_U75 (.A2( u1_u13_X_27 ) , .A1( u1_u13_X_30 ) , .ZN( u1_u13_u4_n102 ) );
  NOR2_X1 u1_u13_u4_U76 (.A2( u1_u13_X_25 ) , .A1( u1_u13_X_26 ) , .ZN( u1_u13_u4_n98 ) );
  AND2_X1 u1_u13_u4_U77 (.A2( u1_u13_X_25 ) , .A1( u1_u13_X_26 ) , .ZN( u1_u13_u4_n104 ) );
  AND2_X1 u1_u13_u4_U78 (.A1( u1_u13_X_30 ) , .A2( u1_u13_u4_n176 ) , .ZN( u1_u13_u4_n99 ) );
  AND2_X1 u1_u13_u4_U79 (.A1( u1_u13_X_26 ) , .ZN( u1_u13_u4_n101 ) , .A2( u1_u13_u4_n177 ) );
  AOI21_X1 u1_u13_u4_U8 (.ZN( u1_u13_u4_n109 ) , .A( u1_u13_u4_n153 ) , .B1( u1_u13_u4_n159 ) , .B2( u1_u13_u4_n184 ) );
  AND2_X1 u1_u13_u4_U80 (.A1( u1_u13_X_27 ) , .A2( u1_u13_X_30 ) , .ZN( u1_u13_u4_n103 ) );
  INV_X1 u1_u13_u4_U81 (.A( u1_u13_X_28 ) , .ZN( u1_u13_u4_n169 ) );
  INV_X1 u1_u13_u4_U82 (.A( u1_u13_X_29 ) , .ZN( u1_u13_u4_n168 ) );
  INV_X1 u1_u13_u4_U83 (.A( u1_u13_X_25 ) , .ZN( u1_u13_u4_n177 ) );
  INV_X1 u1_u13_u4_U84 (.A( u1_u13_X_27 ) , .ZN( u1_u13_u4_n176 ) );
  NAND4_X1 u1_u13_u4_U85 (.ZN( u1_out13_25 ) , .A4( u1_u13_u4_n139 ) , .A3( u1_u13_u4_n140 ) , .A2( u1_u13_u4_n141 ) , .A1( u1_u13_u4_n142 ) );
  OAI21_X1 u1_u13_u4_U86 (.A( u1_u13_u4_n128 ) , .B2( u1_u13_u4_n129 ) , .B1( u1_u13_u4_n130 ) , .ZN( u1_u13_u4_n142 ) );
  OAI21_X1 u1_u13_u4_U87 (.B2( u1_u13_u4_n131 ) , .ZN( u1_u13_u4_n141 ) , .A( u1_u13_u4_n175 ) , .B1( u1_u13_u4_n183 ) );
  NAND4_X1 u1_u13_u4_U88 (.ZN( u1_out13_14 ) , .A4( u1_u13_u4_n124 ) , .A3( u1_u13_u4_n125 ) , .A2( u1_u13_u4_n126 ) , .A1( u1_u13_u4_n127 ) );
  AOI22_X1 u1_u13_u4_U89 (.B2( u1_u13_u4_n117 ) , .ZN( u1_u13_u4_n126 ) , .A1( u1_u13_u4_n129 ) , .B1( u1_u13_u4_n152 ) , .A2( u1_u13_u4_n175 ) );
  AOI211_X1 u1_u13_u4_U9 (.B( u1_u13_u4_n136 ) , .A( u1_u13_u4_n137 ) , .C2( u1_u13_u4_n138 ) , .ZN( u1_u13_u4_n139 ) , .C1( u1_u13_u4_n182 ) );
  AOI22_X1 u1_u13_u4_U90 (.ZN( u1_u13_u4_n125 ) , .B2( u1_u13_u4_n131 ) , .A2( u1_u13_u4_n132 ) , .B1( u1_u13_u4_n138 ) , .A1( u1_u13_u4_n178 ) );
  NAND4_X1 u1_u13_u4_U91 (.ZN( u1_out13_8 ) , .A4( u1_u13_u4_n110 ) , .A3( u1_u13_u4_n111 ) , .A2( u1_u13_u4_n112 ) , .A1( u1_u13_u4_n186 ) );
  NAND2_X1 u1_u13_u4_U92 (.ZN( u1_u13_u4_n112 ) , .A2( u1_u13_u4_n130 ) , .A1( u1_u13_u4_n150 ) );
  AOI22_X1 u1_u13_u4_U93 (.ZN( u1_u13_u4_n111 ) , .B2( u1_u13_u4_n132 ) , .A1( u1_u13_u4_n152 ) , .B1( u1_u13_u4_n178 ) , .A2( u1_u13_u4_n97 ) );
  AOI22_X1 u1_u13_u4_U94 (.B2( u1_u13_u4_n149 ) , .B1( u1_u13_u4_n150 ) , .A2( u1_u13_u4_n151 ) , .A1( u1_u13_u4_n152 ) , .ZN( u1_u13_u4_n167 ) );
  NOR4_X1 u1_u13_u4_U95 (.A4( u1_u13_u4_n162 ) , .A3( u1_u13_u4_n163 ) , .A2( u1_u13_u4_n164 ) , .A1( u1_u13_u4_n165 ) , .ZN( u1_u13_u4_n166 ) );
  NAND3_X1 u1_u13_u4_U96 (.ZN( u1_out13_3 ) , .A3( u1_u13_u4_n166 ) , .A1( u1_u13_u4_n167 ) , .A2( u1_u13_u4_n186 ) );
  NAND3_X1 u1_u13_u4_U97 (.A3( u1_u13_u4_n146 ) , .A2( u1_u13_u4_n147 ) , .A1( u1_u13_u4_n148 ) , .ZN( u1_u13_u4_n149 ) );
  NAND3_X1 u1_u13_u4_U98 (.A3( u1_u13_u4_n143 ) , .A2( u1_u13_u4_n144 ) , .A1( u1_u13_u4_n145 ) , .ZN( u1_u13_u4_n151 ) );
  NAND3_X1 u1_u13_u4_U99 (.A3( u1_u13_u4_n121 ) , .ZN( u1_u13_u4_n122 ) , .A2( u1_u13_u4_n144 ) , .A1( u1_u13_u4_n154 ) );
  AOI22_X1 u1_u13_u6_U10 (.A2( u1_u13_u6_n151 ) , .B2( u1_u13_u6_n161 ) , .A1( u1_u13_u6_n167 ) , .B1( u1_u13_u6_n170 ) , .ZN( u1_u13_u6_n89 ) );
  AOI21_X1 u1_u13_u6_U11 (.B1( u1_u13_u6_n107 ) , .B2( u1_u13_u6_n132 ) , .A( u1_u13_u6_n158 ) , .ZN( u1_u13_u6_n88 ) );
  AOI21_X1 u1_u13_u6_U12 (.B2( u1_u13_u6_n147 ) , .B1( u1_u13_u6_n148 ) , .ZN( u1_u13_u6_n149 ) , .A( u1_u13_u6_n158 ) );
  AOI21_X1 u1_u13_u6_U13 (.ZN( u1_u13_u6_n106 ) , .A( u1_u13_u6_n142 ) , .B2( u1_u13_u6_n159 ) , .B1( u1_u13_u6_n164 ) );
  INV_X1 u1_u13_u6_U14 (.A( u1_u13_u6_n155 ) , .ZN( u1_u13_u6_n161 ) );
  INV_X1 u1_u13_u6_U15 (.A( u1_u13_u6_n128 ) , .ZN( u1_u13_u6_n164 ) );
  NAND2_X1 u1_u13_u6_U16 (.ZN( u1_u13_u6_n110 ) , .A1( u1_u13_u6_n122 ) , .A2( u1_u13_u6_n129 ) );
  NAND2_X1 u1_u13_u6_U17 (.ZN( u1_u13_u6_n124 ) , .A2( u1_u13_u6_n146 ) , .A1( u1_u13_u6_n148 ) );
  INV_X1 u1_u13_u6_U18 (.A( u1_u13_u6_n132 ) , .ZN( u1_u13_u6_n171 ) );
  AND2_X1 u1_u13_u6_U19 (.A1( u1_u13_u6_n100 ) , .ZN( u1_u13_u6_n130 ) , .A2( u1_u13_u6_n147 ) );
  INV_X1 u1_u13_u6_U20 (.A( u1_u13_u6_n127 ) , .ZN( u1_u13_u6_n173 ) );
  INV_X1 u1_u13_u6_U21 (.A( u1_u13_u6_n121 ) , .ZN( u1_u13_u6_n167 ) );
  INV_X1 u1_u13_u6_U22 (.A( u1_u13_u6_n100 ) , .ZN( u1_u13_u6_n169 ) );
  INV_X1 u1_u13_u6_U23 (.A( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n170 ) );
  INV_X1 u1_u13_u6_U24 (.A( u1_u13_u6_n113 ) , .ZN( u1_u13_u6_n168 ) );
  AND2_X1 u1_u13_u6_U25 (.A1( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n119 ) , .ZN( u1_u13_u6_n133 ) );
  AND2_X1 u1_u13_u6_U26 (.A2( u1_u13_u6_n121 ) , .A1( u1_u13_u6_n122 ) , .ZN( u1_u13_u6_n131 ) );
  AND3_X1 u1_u13_u6_U27 (.ZN( u1_u13_u6_n120 ) , .A2( u1_u13_u6_n127 ) , .A1( u1_u13_u6_n132 ) , .A3( u1_u13_u6_n145 ) );
  INV_X1 u1_u13_u6_U28 (.A( u1_u13_u6_n146 ) , .ZN( u1_u13_u6_n163 ) );
  AOI222_X1 u1_u13_u6_U29 (.ZN( u1_u13_u6_n114 ) , .A1( u1_u13_u6_n118 ) , .A2( u1_u13_u6_n126 ) , .B2( u1_u13_u6_n151 ) , .C2( u1_u13_u6_n159 ) , .C1( u1_u13_u6_n168 ) , .B1( u1_u13_u6_n169 ) );
  INV_X1 u1_u13_u6_U3 (.A( u1_u13_u6_n110 ) , .ZN( u1_u13_u6_n166 ) );
  NOR2_X1 u1_u13_u6_U30 (.A1( u1_u13_u6_n162 ) , .A2( u1_u13_u6_n165 ) , .ZN( u1_u13_u6_n98 ) );
  AOI211_X1 u1_u13_u6_U31 (.B( u1_u13_u6_n134 ) , .A( u1_u13_u6_n135 ) , .C1( u1_u13_u6_n136 ) , .ZN( u1_u13_u6_n137 ) , .C2( u1_u13_u6_n151 ) );
  AOI21_X1 u1_u13_u6_U32 (.B2( u1_u13_u6_n132 ) , .B1( u1_u13_u6_n133 ) , .ZN( u1_u13_u6_n134 ) , .A( u1_u13_u6_n158 ) );
  AOI21_X1 u1_u13_u6_U33 (.B1( u1_u13_u6_n131 ) , .ZN( u1_u13_u6_n135 ) , .A( u1_u13_u6_n144 ) , .B2( u1_u13_u6_n146 ) );
  NAND4_X1 u1_u13_u6_U34 (.A4( u1_u13_u6_n127 ) , .A3( u1_u13_u6_n128 ) , .A2( u1_u13_u6_n129 ) , .A1( u1_u13_u6_n130 ) , .ZN( u1_u13_u6_n136 ) );
  NAND2_X1 u1_u13_u6_U35 (.A1( u1_u13_u6_n144 ) , .ZN( u1_u13_u6_n151 ) , .A2( u1_u13_u6_n158 ) );
  NAND2_X1 u1_u13_u6_U36 (.ZN( u1_u13_u6_n132 ) , .A1( u1_u13_u6_n91 ) , .A2( u1_u13_u6_n97 ) );
  AOI22_X1 u1_u13_u6_U37 (.B2( u1_u13_u6_n110 ) , .B1( u1_u13_u6_n111 ) , .A1( u1_u13_u6_n112 ) , .ZN( u1_u13_u6_n115 ) , .A2( u1_u13_u6_n161 ) );
  NAND4_X1 u1_u13_u6_U38 (.A3( u1_u13_u6_n109 ) , .ZN( u1_u13_u6_n112 ) , .A4( u1_u13_u6_n132 ) , .A2( u1_u13_u6_n147 ) , .A1( u1_u13_u6_n166 ) );
  NOR2_X1 u1_u13_u6_U39 (.ZN( u1_u13_u6_n109 ) , .A1( u1_u13_u6_n170 ) , .A2( u1_u13_u6_n173 ) );
  INV_X1 u1_u13_u6_U4 (.A( u1_u13_u6_n142 ) , .ZN( u1_u13_u6_n174 ) );
  NOR2_X1 u1_u13_u6_U40 (.A2( u1_u13_u6_n126 ) , .ZN( u1_u13_u6_n155 ) , .A1( u1_u13_u6_n160 ) );
  NAND2_X1 u1_u13_u6_U41 (.ZN( u1_u13_u6_n146 ) , .A2( u1_u13_u6_n94 ) , .A1( u1_u13_u6_n99 ) );
  AOI21_X1 u1_u13_u6_U42 (.A( u1_u13_u6_n144 ) , .B2( u1_u13_u6_n145 ) , .B1( u1_u13_u6_n146 ) , .ZN( u1_u13_u6_n150 ) );
  INV_X1 u1_u13_u6_U43 (.A( u1_u13_u6_n111 ) , .ZN( u1_u13_u6_n158 ) );
  NAND2_X1 u1_u13_u6_U44 (.ZN( u1_u13_u6_n127 ) , .A1( u1_u13_u6_n91 ) , .A2( u1_u13_u6_n92 ) );
  NAND2_X1 u1_u13_u6_U45 (.ZN( u1_u13_u6_n129 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n96 ) );
  INV_X1 u1_u13_u6_U46 (.A( u1_u13_u6_n144 ) , .ZN( u1_u13_u6_n159 ) );
  NAND2_X1 u1_u13_u6_U47 (.ZN( u1_u13_u6_n145 ) , .A2( u1_u13_u6_n97 ) , .A1( u1_u13_u6_n98 ) );
  NAND2_X1 u1_u13_u6_U48 (.ZN( u1_u13_u6_n148 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n94 ) );
  NAND2_X1 u1_u13_u6_U49 (.ZN( u1_u13_u6_n108 ) , .A2( u1_u13_u6_n139 ) , .A1( u1_u13_u6_n144 ) );
  NAND2_X1 u1_u13_u6_U5 (.A2( u1_u13_u6_n143 ) , .ZN( u1_u13_u6_n152 ) , .A1( u1_u13_u6_n166 ) );
  NAND2_X1 u1_u13_u6_U50 (.ZN( u1_u13_u6_n121 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n97 ) );
  NAND2_X1 u1_u13_u6_U51 (.ZN( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n95 ) );
  AND2_X1 u1_u13_u6_U52 (.ZN( u1_u13_u6_n118 ) , .A2( u1_u13_u6_n91 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U53 (.ZN( u1_u13_u6_n147 ) , .A2( u1_u13_u6_n98 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U54 (.ZN( u1_u13_u6_n128 ) , .A1( u1_u13_u6_n94 ) , .A2( u1_u13_u6_n96 ) );
  NAND2_X1 u1_u13_u6_U55 (.ZN( u1_u13_u6_n119 ) , .A2( u1_u13_u6_n95 ) , .A1( u1_u13_u6_n99 ) );
  NAND2_X1 u1_u13_u6_U56 (.ZN( u1_u13_u6_n123 ) , .A2( u1_u13_u6_n91 ) , .A1( u1_u13_u6_n96 ) );
  NAND2_X1 u1_u13_u6_U57 (.ZN( u1_u13_u6_n100 ) , .A2( u1_u13_u6_n92 ) , .A1( u1_u13_u6_n98 ) );
  NAND2_X1 u1_u13_u6_U58 (.ZN( u1_u13_u6_n122 ) , .A1( u1_u13_u6_n94 ) , .A2( u1_u13_u6_n97 ) );
  INV_X1 u1_u13_u6_U59 (.A( u1_u13_u6_n139 ) , .ZN( u1_u13_u6_n160 ) );
  AOI22_X1 u1_u13_u6_U6 (.B2( u1_u13_u6_n101 ) , .A1( u1_u13_u6_n102 ) , .ZN( u1_u13_u6_n103 ) , .B1( u1_u13_u6_n160 ) , .A2( u1_u13_u6_n161 ) );
  NAND2_X1 u1_u13_u6_U60 (.ZN( u1_u13_u6_n113 ) , .A1( u1_u13_u6_n96 ) , .A2( u1_u13_u6_n98 ) );
  NOR2_X1 u1_u13_u6_U61 (.A2( u1_u13_X_40 ) , .A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n126 ) );
  NOR2_X1 u1_u13_u6_U62 (.A2( u1_u13_X_39 ) , .A1( u1_u13_X_42 ) , .ZN( u1_u13_u6_n92 ) );
  NOR2_X1 u1_u13_u6_U63 (.A2( u1_u13_X_39 ) , .A1( u1_u13_u6_n156 ) , .ZN( u1_u13_u6_n97 ) );
  NOR2_X1 u1_u13_u6_U64 (.A2( u1_u13_X_38 ) , .A1( u1_u13_u6_n165 ) , .ZN( u1_u13_u6_n95 ) );
  NOR2_X1 u1_u13_u6_U65 (.A2( u1_u13_X_41 ) , .ZN( u1_u13_u6_n111 ) , .A1( u1_u13_u6_n157 ) );
  NOR2_X1 u1_u13_u6_U66 (.A2( u1_u13_X_37 ) , .A1( u1_u13_u6_n162 ) , .ZN( u1_u13_u6_n94 ) );
  NOR2_X1 u1_u13_u6_U67 (.A2( u1_u13_X_37 ) , .A1( u1_u13_X_38 ) , .ZN( u1_u13_u6_n91 ) );
  NAND2_X1 u1_u13_u6_U68 (.A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n144 ) , .A2( u1_u13_u6_n157 ) );
  NAND2_X1 u1_u13_u6_U69 (.A2( u1_u13_X_40 ) , .A1( u1_u13_X_41 ) , .ZN( u1_u13_u6_n139 ) );
  NOR2_X1 u1_u13_u6_U7 (.A1( u1_u13_u6_n118 ) , .ZN( u1_u13_u6_n143 ) , .A2( u1_u13_u6_n168 ) );
  AND2_X1 u1_u13_u6_U70 (.A1( u1_u13_X_39 ) , .A2( u1_u13_u6_n156 ) , .ZN( u1_u13_u6_n96 ) );
  AND2_X1 u1_u13_u6_U71 (.A1( u1_u13_X_39 ) , .A2( u1_u13_X_42 ) , .ZN( u1_u13_u6_n99 ) );
  INV_X1 u1_u13_u6_U72 (.A( u1_u13_X_40 ) , .ZN( u1_u13_u6_n157 ) );
  INV_X1 u1_u13_u6_U73 (.A( u1_u13_X_37 ) , .ZN( u1_u13_u6_n165 ) );
  INV_X1 u1_u13_u6_U74 (.A( u1_u13_X_38 ) , .ZN( u1_u13_u6_n162 ) );
  INV_X1 u1_u13_u6_U75 (.A( u1_u13_X_42 ) , .ZN( u1_u13_u6_n156 ) );
  NAND4_X1 u1_u13_u6_U76 (.ZN( u1_out13_32 ) , .A4( u1_u13_u6_n103 ) , .A3( u1_u13_u6_n104 ) , .A2( u1_u13_u6_n105 ) , .A1( u1_u13_u6_n106 ) );
  AOI22_X1 u1_u13_u6_U77 (.ZN( u1_u13_u6_n105 ) , .A2( u1_u13_u6_n108 ) , .A1( u1_u13_u6_n118 ) , .B2( u1_u13_u6_n126 ) , .B1( u1_u13_u6_n171 ) );
  AOI22_X1 u1_u13_u6_U78 (.ZN( u1_u13_u6_n104 ) , .A1( u1_u13_u6_n111 ) , .B1( u1_u13_u6_n124 ) , .B2( u1_u13_u6_n151 ) , .A2( u1_u13_u6_n93 ) );
  NAND4_X1 u1_u13_u6_U79 (.ZN( u1_out13_12 ) , .A4( u1_u13_u6_n114 ) , .A3( u1_u13_u6_n115 ) , .A2( u1_u13_u6_n116 ) , .A1( u1_u13_u6_n117 ) );
  OAI21_X1 u1_u13_u6_U8 (.A( u1_u13_u6_n159 ) , .B1( u1_u13_u6_n169 ) , .B2( u1_u13_u6_n173 ) , .ZN( u1_u13_u6_n90 ) );
  OAI22_X1 u1_u13_u6_U80 (.B2( u1_u13_u6_n111 ) , .ZN( u1_u13_u6_n116 ) , .B1( u1_u13_u6_n126 ) , .A2( u1_u13_u6_n164 ) , .A1( u1_u13_u6_n167 ) );
  OAI21_X1 u1_u13_u6_U81 (.A( u1_u13_u6_n108 ) , .ZN( u1_u13_u6_n117 ) , .B2( u1_u13_u6_n141 ) , .B1( u1_u13_u6_n163 ) );
  OAI211_X1 u1_u13_u6_U82 (.ZN( u1_out13_7 ) , .B( u1_u13_u6_n153 ) , .C2( u1_u13_u6_n154 ) , .C1( u1_u13_u6_n155 ) , .A( u1_u13_u6_n174 ) );
  NOR3_X1 u1_u13_u6_U83 (.A1( u1_u13_u6_n141 ) , .ZN( u1_u13_u6_n154 ) , .A3( u1_u13_u6_n164 ) , .A2( u1_u13_u6_n171 ) );
  AOI211_X1 u1_u13_u6_U84 (.B( u1_u13_u6_n149 ) , .A( u1_u13_u6_n150 ) , .C2( u1_u13_u6_n151 ) , .C1( u1_u13_u6_n152 ) , .ZN( u1_u13_u6_n153 ) );
  OAI211_X1 u1_u13_u6_U85 (.ZN( u1_out13_22 ) , .B( u1_u13_u6_n137 ) , .A( u1_u13_u6_n138 ) , .C2( u1_u13_u6_n139 ) , .C1( u1_u13_u6_n140 ) );
  AOI22_X1 u1_u13_u6_U86 (.B1( u1_u13_u6_n124 ) , .A2( u1_u13_u6_n125 ) , .A1( u1_u13_u6_n126 ) , .ZN( u1_u13_u6_n138 ) , .B2( u1_u13_u6_n161 ) );
  AND4_X1 u1_u13_u6_U87 (.A3( u1_u13_u6_n119 ) , .A1( u1_u13_u6_n120 ) , .A4( u1_u13_u6_n129 ) , .ZN( u1_u13_u6_n140 ) , .A2( u1_u13_u6_n143 ) );
  NAND3_X1 u1_u13_u6_U88 (.A2( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n125 ) , .A1( u1_u13_u6_n130 ) , .A3( u1_u13_u6_n131 ) );
  NAND3_X1 u1_u13_u6_U89 (.A3( u1_u13_u6_n133 ) , .ZN( u1_u13_u6_n141 ) , .A1( u1_u13_u6_n145 ) , .A2( u1_u13_u6_n148 ) );
  INV_X1 u1_u13_u6_U9 (.ZN( u1_u13_u6_n172 ) , .A( u1_u13_u6_n88 ) );
  NAND3_X1 u1_u13_u6_U90 (.ZN( u1_u13_u6_n101 ) , .A3( u1_u13_u6_n107 ) , .A2( u1_u13_u6_n121 ) , .A1( u1_u13_u6_n127 ) );
  NAND3_X1 u1_u13_u6_U91 (.ZN( u1_u13_u6_n102 ) , .A3( u1_u13_u6_n130 ) , .A2( u1_u13_u6_n145 ) , .A1( u1_u13_u6_n166 ) );
  NAND3_X1 u1_u13_u6_U92 (.A3( u1_u13_u6_n113 ) , .A1( u1_u13_u6_n119 ) , .A2( u1_u13_u6_n123 ) , .ZN( u1_u13_u6_n93 ) );
  NAND3_X1 u1_u13_u6_U93 (.ZN( u1_u13_u6_n142 ) , .A2( u1_u13_u6_n172 ) , .A3( u1_u13_u6_n89 ) , .A1( u1_u13_u6_n90 ) );
  AND3_X1 u1_u13_u7_U10 (.A3( u1_u13_u7_n110 ) , .A2( u1_u13_u7_n127 ) , .A1( u1_u13_u7_n132 ) , .ZN( u1_u13_u7_n92 ) );
  OAI21_X1 u1_u13_u7_U11 (.A( u1_u13_u7_n161 ) , .B1( u1_u13_u7_n168 ) , .B2( u1_u13_u7_n173 ) , .ZN( u1_u13_u7_n91 ) );
  AOI211_X1 u1_u13_u7_U12 (.A( u1_u13_u7_n117 ) , .ZN( u1_u13_u7_n118 ) , .C2( u1_u13_u7_n126 ) , .C1( u1_u13_u7_n177 ) , .B( u1_u13_u7_n180 ) );
  OAI22_X1 u1_u13_u7_U13 (.B1( u1_u13_u7_n115 ) , .ZN( u1_u13_u7_n117 ) , .A2( u1_u13_u7_n133 ) , .A1( u1_u13_u7_n137 ) , .B2( u1_u13_u7_n162 ) );
  INV_X1 u1_u13_u7_U14 (.A( u1_u13_u7_n116 ) , .ZN( u1_u13_u7_n180 ) );
  NOR3_X1 u1_u13_u7_U15 (.ZN( u1_u13_u7_n115 ) , .A3( u1_u13_u7_n145 ) , .A2( u1_u13_u7_n168 ) , .A1( u1_u13_u7_n169 ) );
  OAI211_X1 u1_u13_u7_U16 (.B( u1_u13_u7_n122 ) , .A( u1_u13_u7_n123 ) , .C2( u1_u13_u7_n124 ) , .ZN( u1_u13_u7_n154 ) , .C1( u1_u13_u7_n162 ) );
  AOI222_X1 u1_u13_u7_U17 (.ZN( u1_u13_u7_n122 ) , .C2( u1_u13_u7_n126 ) , .C1( u1_u13_u7_n145 ) , .B1( u1_u13_u7_n161 ) , .A2( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n170 ) , .A1( u1_u13_u7_n176 ) );
  INV_X1 u1_u13_u7_U18 (.A( u1_u13_u7_n133 ) , .ZN( u1_u13_u7_n176 ) );
  NOR3_X1 u1_u13_u7_U19 (.A2( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n135 ) , .ZN( u1_u13_u7_n136 ) , .A3( u1_u13_u7_n171 ) );
  NOR2_X1 u1_u13_u7_U20 (.A1( u1_u13_u7_n130 ) , .A2( u1_u13_u7_n134 ) , .ZN( u1_u13_u7_n153 ) );
  INV_X1 u1_u13_u7_U21 (.A( u1_u13_u7_n101 ) , .ZN( u1_u13_u7_n165 ) );
  NOR2_X1 u1_u13_u7_U22 (.ZN( u1_u13_u7_n111 ) , .A2( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n169 ) );
  AOI21_X1 u1_u13_u7_U23 (.ZN( u1_u13_u7_n104 ) , .B2( u1_u13_u7_n112 ) , .B1( u1_u13_u7_n127 ) , .A( u1_u13_u7_n164 ) );
  AOI21_X1 u1_u13_u7_U24 (.ZN( u1_u13_u7_n106 ) , .B1( u1_u13_u7_n133 ) , .B2( u1_u13_u7_n146 ) , .A( u1_u13_u7_n162 ) );
  AOI21_X1 u1_u13_u7_U25 (.A( u1_u13_u7_n101 ) , .ZN( u1_u13_u7_n107 ) , .B2( u1_u13_u7_n128 ) , .B1( u1_u13_u7_n175 ) );
  INV_X1 u1_u13_u7_U26 (.A( u1_u13_u7_n138 ) , .ZN( u1_u13_u7_n171 ) );
  INV_X1 u1_u13_u7_U27 (.A( u1_u13_u7_n131 ) , .ZN( u1_u13_u7_n177 ) );
  INV_X1 u1_u13_u7_U28 (.A( u1_u13_u7_n110 ) , .ZN( u1_u13_u7_n174 ) );
  NAND2_X1 u1_u13_u7_U29 (.A1( u1_u13_u7_n129 ) , .A2( u1_u13_u7_n132 ) , .ZN( u1_u13_u7_n149 ) );
  OAI21_X1 u1_u13_u7_U3 (.ZN( u1_u13_u7_n159 ) , .A( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n171 ) , .B1( u1_u13_u7_n174 ) );
  NAND2_X1 u1_u13_u7_U30 (.A1( u1_u13_u7_n113 ) , .A2( u1_u13_u7_n124 ) , .ZN( u1_u13_u7_n130 ) );
  INV_X1 u1_u13_u7_U31 (.A( u1_u13_u7_n112 ) , .ZN( u1_u13_u7_n173 ) );
  INV_X1 u1_u13_u7_U32 (.A( u1_u13_u7_n128 ) , .ZN( u1_u13_u7_n168 ) );
  INV_X1 u1_u13_u7_U33 (.A( u1_u13_u7_n148 ) , .ZN( u1_u13_u7_n169 ) );
  INV_X1 u1_u13_u7_U34 (.A( u1_u13_u7_n127 ) , .ZN( u1_u13_u7_n179 ) );
  NOR2_X1 u1_u13_u7_U35 (.ZN( u1_u13_u7_n101 ) , .A2( u1_u13_u7_n150 ) , .A1( u1_u13_u7_n156 ) );
  AOI211_X1 u1_u13_u7_U36 (.B( u1_u13_u7_n154 ) , .A( u1_u13_u7_n155 ) , .C1( u1_u13_u7_n156 ) , .ZN( u1_u13_u7_n157 ) , .C2( u1_u13_u7_n172 ) );
  INV_X1 u1_u13_u7_U37 (.A( u1_u13_u7_n153 ) , .ZN( u1_u13_u7_n172 ) );
  AOI211_X1 u1_u13_u7_U38 (.B( u1_u13_u7_n139 ) , .A( u1_u13_u7_n140 ) , .C2( u1_u13_u7_n141 ) , .ZN( u1_u13_u7_n142 ) , .C1( u1_u13_u7_n156 ) );
  NAND4_X1 u1_u13_u7_U39 (.A3( u1_u13_u7_n127 ) , .A2( u1_u13_u7_n128 ) , .A1( u1_u13_u7_n129 ) , .ZN( u1_u13_u7_n141 ) , .A4( u1_u13_u7_n147 ) );
  INV_X1 u1_u13_u7_U4 (.A( u1_u13_u7_n111 ) , .ZN( u1_u13_u7_n170 ) );
  AOI21_X1 u1_u13_u7_U40 (.A( u1_u13_u7_n137 ) , .B1( u1_u13_u7_n138 ) , .ZN( u1_u13_u7_n139 ) , .B2( u1_u13_u7_n146 ) );
  OAI22_X1 u1_u13_u7_U41 (.B1( u1_u13_u7_n136 ) , .ZN( u1_u13_u7_n140 ) , .A1( u1_u13_u7_n153 ) , .B2( u1_u13_u7_n162 ) , .A2( u1_u13_u7_n164 ) );
  AOI21_X1 u1_u13_u7_U42 (.ZN( u1_u13_u7_n123 ) , .B1( u1_u13_u7_n165 ) , .B2( u1_u13_u7_n177 ) , .A( u1_u13_u7_n97 ) );
  AOI21_X1 u1_u13_u7_U43 (.B2( u1_u13_u7_n113 ) , .B1( u1_u13_u7_n124 ) , .A( u1_u13_u7_n125 ) , .ZN( u1_u13_u7_n97 ) );
  INV_X1 u1_u13_u7_U44 (.A( u1_u13_u7_n125 ) , .ZN( u1_u13_u7_n161 ) );
  INV_X1 u1_u13_u7_U45 (.A( u1_u13_u7_n152 ) , .ZN( u1_u13_u7_n162 ) );
  AOI22_X1 u1_u13_u7_U46 (.A2( u1_u13_u7_n114 ) , .ZN( u1_u13_u7_n119 ) , .B1( u1_u13_u7_n130 ) , .A1( u1_u13_u7_n156 ) , .B2( u1_u13_u7_n165 ) );
  NAND2_X1 u1_u13_u7_U47 (.A2( u1_u13_u7_n112 ) , .ZN( u1_u13_u7_n114 ) , .A1( u1_u13_u7_n175 ) );
  AND2_X1 u1_u13_u7_U48 (.ZN( u1_u13_u7_n145 ) , .A2( u1_u13_u7_n98 ) , .A1( u1_u13_u7_n99 ) );
  NOR2_X1 u1_u13_u7_U49 (.ZN( u1_u13_u7_n137 ) , .A1( u1_u13_u7_n150 ) , .A2( u1_u13_u7_n161 ) );
  INV_X1 u1_u13_u7_U5 (.A( u1_u13_u7_n149 ) , .ZN( u1_u13_u7_n175 ) );
  AOI21_X1 u1_u13_u7_U50 (.ZN( u1_u13_u7_n105 ) , .B2( u1_u13_u7_n110 ) , .A( u1_u13_u7_n125 ) , .B1( u1_u13_u7_n147 ) );
  NAND2_X1 u1_u13_u7_U51 (.ZN( u1_u13_u7_n146 ) , .A1( u1_u13_u7_n95 ) , .A2( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U52 (.A2( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n147 ) , .A1( u1_u13_u7_n93 ) );
  NAND2_X1 u1_u13_u7_U53 (.A1( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n127 ) , .A2( u1_u13_u7_n99 ) );
  OR2_X1 u1_u13_u7_U54 (.ZN( u1_u13_u7_n126 ) , .A2( u1_u13_u7_n152 ) , .A1( u1_u13_u7_n156 ) );
  NAND2_X1 u1_u13_u7_U55 (.A2( u1_u13_u7_n102 ) , .A1( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n133 ) );
  NAND2_X1 u1_u13_u7_U56 (.ZN( u1_u13_u7_n112 ) , .A2( u1_u13_u7_n96 ) , .A1( u1_u13_u7_n99 ) );
  NAND2_X1 u1_u13_u7_U57 (.A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n128 ) , .A1( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U58 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n113 ) , .A2( u1_u13_u7_n93 ) );
  NAND2_X1 u1_u13_u7_U59 (.A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n124 ) , .A1( u1_u13_u7_n96 ) );
  INV_X1 u1_u13_u7_U6 (.A( u1_u13_u7_n154 ) , .ZN( u1_u13_u7_n178 ) );
  NAND2_X1 u1_u13_u7_U60 (.ZN( u1_u13_u7_n110 ) , .A1( u1_u13_u7_n95 ) , .A2( u1_u13_u7_n96 ) );
  INV_X1 u1_u13_u7_U61 (.A( u1_u13_u7_n150 ) , .ZN( u1_u13_u7_n164 ) );
  AND2_X1 u1_u13_u7_U62 (.ZN( u1_u13_u7_n134 ) , .A1( u1_u13_u7_n93 ) , .A2( u1_u13_u7_n98 ) );
  NAND2_X1 u1_u13_u7_U63 (.A1( u1_u13_u7_n100 ) , .A2( u1_u13_u7_n102 ) , .ZN( u1_u13_u7_n129 ) );
  NAND2_X1 u1_u13_u7_U64 (.A2( u1_u13_u7_n103 ) , .ZN( u1_u13_u7_n131 ) , .A1( u1_u13_u7_n95 ) );
  NAND2_X1 u1_u13_u7_U65 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n138 ) , .A2( u1_u13_u7_n99 ) );
  NAND2_X1 u1_u13_u7_U66 (.ZN( u1_u13_u7_n132 ) , .A1( u1_u13_u7_n93 ) , .A2( u1_u13_u7_n96 ) );
  NAND2_X1 u1_u13_u7_U67 (.A1( u1_u13_u7_n100 ) , .ZN( u1_u13_u7_n148 ) , .A2( u1_u13_u7_n95 ) );
  NOR2_X1 u1_u13_u7_U68 (.A2( u1_u13_X_47 ) , .ZN( u1_u13_u7_n150 ) , .A1( u1_u13_u7_n163 ) );
  NOR2_X1 u1_u13_u7_U69 (.A2( u1_u13_X_43 ) , .A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n103 ) );
  AOI211_X1 u1_u13_u7_U7 (.ZN( u1_u13_u7_n116 ) , .A( u1_u13_u7_n155 ) , .C1( u1_u13_u7_n161 ) , .C2( u1_u13_u7_n171 ) , .B( u1_u13_u7_n94 ) );
  NOR2_X1 u1_u13_u7_U70 (.A2( u1_u13_X_48 ) , .A1( u1_u13_u7_n166 ) , .ZN( u1_u13_u7_n95 ) );
  NOR2_X1 u1_u13_u7_U71 (.A2( u1_u13_X_45 ) , .A1( u1_u13_X_48 ) , .ZN( u1_u13_u7_n99 ) );
  NOR2_X1 u1_u13_u7_U72 (.A2( u1_u13_X_44 ) , .A1( u1_u13_u7_n167 ) , .ZN( u1_u13_u7_n98 ) );
  NOR2_X1 u1_u13_u7_U73 (.A2( u1_u13_X_46 ) , .A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n152 ) );
  AND2_X1 u1_u13_u7_U74 (.A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n156 ) , .A2( u1_u13_u7_n163 ) );
  NAND2_X1 u1_u13_u7_U75 (.A2( u1_u13_X_46 ) , .A1( u1_u13_X_47 ) , .ZN( u1_u13_u7_n125 ) );
  AND2_X1 u1_u13_u7_U76 (.A2( u1_u13_X_45 ) , .A1( u1_u13_X_48 ) , .ZN( u1_u13_u7_n102 ) );
  AND2_X1 u1_u13_u7_U77 (.A2( u1_u13_X_43 ) , .A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n96 ) );
  AND2_X1 u1_u13_u7_U78 (.A1( u1_u13_X_44 ) , .ZN( u1_u13_u7_n100 ) , .A2( u1_u13_u7_n167 ) );
  AND2_X1 u1_u13_u7_U79 (.A1( u1_u13_X_48 ) , .A2( u1_u13_u7_n166 ) , .ZN( u1_u13_u7_n93 ) );
  OAI222_X1 u1_u13_u7_U8 (.C2( u1_u13_u7_n101 ) , .B2( u1_u13_u7_n111 ) , .A1( u1_u13_u7_n113 ) , .C1( u1_u13_u7_n146 ) , .A2( u1_u13_u7_n162 ) , .B1( u1_u13_u7_n164 ) , .ZN( u1_u13_u7_n94 ) );
  INV_X1 u1_u13_u7_U80 (.A( u1_u13_X_46 ) , .ZN( u1_u13_u7_n163 ) );
  INV_X1 u1_u13_u7_U81 (.A( u1_u13_X_43 ) , .ZN( u1_u13_u7_n167 ) );
  INV_X1 u1_u13_u7_U82 (.A( u1_u13_X_45 ) , .ZN( u1_u13_u7_n166 ) );
  NAND4_X1 u1_u13_u7_U83 (.ZN( u1_out13_5 ) , .A4( u1_u13_u7_n108 ) , .A3( u1_u13_u7_n109 ) , .A1( u1_u13_u7_n116 ) , .A2( u1_u13_u7_n123 ) );
  AOI22_X1 u1_u13_u7_U84 (.ZN( u1_u13_u7_n109 ) , .A2( u1_u13_u7_n126 ) , .B2( u1_u13_u7_n145 ) , .B1( u1_u13_u7_n156 ) , .A1( u1_u13_u7_n171 ) );
  NOR4_X1 u1_u13_u7_U85 (.A4( u1_u13_u7_n104 ) , .A3( u1_u13_u7_n105 ) , .A2( u1_u13_u7_n106 ) , .A1( u1_u13_u7_n107 ) , .ZN( u1_u13_u7_n108 ) );
  NAND4_X1 u1_u13_u7_U86 (.ZN( u1_out13_27 ) , .A4( u1_u13_u7_n118 ) , .A3( u1_u13_u7_n119 ) , .A2( u1_u13_u7_n120 ) , .A1( u1_u13_u7_n121 ) );
  OAI21_X1 u1_u13_u7_U87 (.ZN( u1_u13_u7_n121 ) , .B2( u1_u13_u7_n145 ) , .A( u1_u13_u7_n150 ) , .B1( u1_u13_u7_n174 ) );
  OAI21_X1 u1_u13_u7_U88 (.ZN( u1_u13_u7_n120 ) , .A( u1_u13_u7_n161 ) , .B2( u1_u13_u7_n170 ) , .B1( u1_u13_u7_n179 ) );
  NAND4_X1 u1_u13_u7_U89 (.ZN( u1_out13_21 ) , .A4( u1_u13_u7_n157 ) , .A3( u1_u13_u7_n158 ) , .A2( u1_u13_u7_n159 ) , .A1( u1_u13_u7_n160 ) );
  OAI221_X1 u1_u13_u7_U9 (.C1( u1_u13_u7_n101 ) , .C2( u1_u13_u7_n147 ) , .ZN( u1_u13_u7_n155 ) , .B2( u1_u13_u7_n162 ) , .A( u1_u13_u7_n91 ) , .B1( u1_u13_u7_n92 ) );
  OAI21_X1 u1_u13_u7_U90 (.B1( u1_u13_u7_n145 ) , .ZN( u1_u13_u7_n160 ) , .A( u1_u13_u7_n161 ) , .B2( u1_u13_u7_n177 ) );
  AOI22_X1 u1_u13_u7_U91 (.B2( u1_u13_u7_n149 ) , .B1( u1_u13_u7_n150 ) , .A2( u1_u13_u7_n151 ) , .A1( u1_u13_u7_n152 ) , .ZN( u1_u13_u7_n158 ) );
  NAND4_X1 u1_u13_u7_U92 (.ZN( u1_out13_15 ) , .A4( u1_u13_u7_n142 ) , .A3( u1_u13_u7_n143 ) , .A2( u1_u13_u7_n144 ) , .A1( u1_u13_u7_n178 ) );
  OR2_X1 u1_u13_u7_U93 (.A2( u1_u13_u7_n125 ) , .A1( u1_u13_u7_n129 ) , .ZN( u1_u13_u7_n144 ) );
  AOI22_X1 u1_u13_u7_U94 (.A2( u1_u13_u7_n126 ) , .ZN( u1_u13_u7_n143 ) , .B2( u1_u13_u7_n165 ) , .B1( u1_u13_u7_n173 ) , .A1( u1_u13_u7_n174 ) );
  NAND3_X1 u1_u13_u7_U95 (.A3( u1_u13_u7_n146 ) , .A2( u1_u13_u7_n147 ) , .A1( u1_u13_u7_n148 ) , .ZN( u1_u13_u7_n151 ) );
  NAND3_X1 u1_u13_u7_U96 (.A3( u1_u13_u7_n131 ) , .A2( u1_u13_u7_n132 ) , .A1( u1_u13_u7_n133 ) , .ZN( u1_u13_u7_n135 ) );
  XOR2_X1 u1_u14_U10 (.B( u1_K15_45 ) , .A( u1_R13_30 ) , .Z( u1_u14_X_45 ) );
  XOR2_X1 u1_u14_U11 (.B( u1_K15_44 ) , .A( u1_R13_29 ) , .Z( u1_u14_X_44 ) );
  XOR2_X1 u1_u14_U12 (.B( u1_K15_43 ) , .A( u1_R13_28 ) , .Z( u1_u14_X_43 ) );
  XOR2_X1 u1_u14_U13 (.B( u1_K15_42 ) , .A( u1_R13_29 ) , .Z( u1_u14_X_42 ) );
  XOR2_X1 u1_u14_U14 (.B( u1_K15_41 ) , .A( u1_R13_28 ) , .Z( u1_u14_X_41 ) );
  XOR2_X1 u1_u14_U15 (.B( u1_K15_40 ) , .A( u1_R13_27 ) , .Z( u1_u14_X_40 ) );
  XOR2_X1 u1_u14_U17 (.B( u1_K15_39 ) , .A( u1_R13_26 ) , .Z( u1_u14_X_39 ) );
  XOR2_X1 u1_u14_U18 (.B( u1_K15_38 ) , .A( u1_R13_25 ) , .Z( u1_u14_X_38 ) );
  XOR2_X1 u1_u14_U19 (.B( u1_K15_37 ) , .A( u1_R13_24 ) , .Z( u1_u14_X_37 ) );
  XOR2_X1 u1_u14_U2 (.B( u1_K15_8 ) , .A( u1_R13_5 ) , .Z( u1_u14_X_8 ) );
  XOR2_X1 u1_u14_U20 (.B( u1_K15_36 ) , .A( u1_R13_25 ) , .Z( u1_u14_X_36 ) );
  XOR2_X1 u1_u14_U21 (.B( u1_K15_35 ) , .A( u1_R13_24 ) , .Z( u1_u14_X_35 ) );
  XOR2_X1 u1_u14_U22 (.B( u1_K15_34 ) , .A( u1_R13_23 ) , .Z( u1_u14_X_34 ) );
  XOR2_X1 u1_u14_U23 (.B( u1_K15_33 ) , .A( u1_R13_22 ) , .Z( u1_u14_X_33 ) );
  XOR2_X1 u1_u14_U24 (.B( u1_K15_32 ) , .A( u1_R13_21 ) , .Z( u1_u14_X_32 ) );
  XOR2_X1 u1_u14_U25 (.B( u1_K15_31 ) , .A( u1_R13_20 ) , .Z( u1_u14_X_31 ) );
  XOR2_X1 u1_u14_U26 (.B( u1_K15_30 ) , .A( u1_R13_21 ) , .Z( u1_u14_X_30 ) );
  XOR2_X1 u1_u14_U27 (.B( u1_K15_2 ) , .A( u1_R13_1 ) , .Z( u1_u14_X_2 ) );
  XOR2_X1 u1_u14_U28 (.B( u1_K15_29 ) , .A( u1_R13_20 ) , .Z( u1_u14_X_29 ) );
  XOR2_X1 u1_u14_U3 (.B( u1_K15_7 ) , .A( u1_R13_4 ) , .Z( u1_u14_X_7 ) );
  XOR2_X1 u1_u14_U31 (.B( u1_K15_26 ) , .A( u1_R13_17 ) , .Z( u1_u14_X_26 ) );
  XOR2_X1 u1_u14_U32 (.B( u1_K15_25 ) , .A( u1_R13_16 ) , .Z( u1_u14_X_25 ) );
  XOR2_X1 u1_u14_U33 (.B( u1_K15_24 ) , .A( u1_R13_17 ) , .Z( u1_u14_X_24 ) );
  XOR2_X1 u1_u14_U34 (.B( u1_K15_23 ) , .A( u1_R13_16 ) , .Z( u1_u14_X_23 ) );
  XOR2_X1 u1_u14_U37 (.B( u1_K15_20 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_20 ) );
  XOR2_X1 u1_u14_U38 (.B( u1_K15_1 ) , .A( u1_R13_32 ) , .Z( u1_u14_X_1 ) );
  XOR2_X1 u1_u14_U39 (.B( u1_K15_19 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_19 ) );
  XOR2_X1 u1_u14_U4 (.B( u1_K15_6 ) , .A( u1_R13_5 ) , .Z( u1_u14_X_6 ) );
  XOR2_X1 u1_u14_U40 (.B( u1_K15_18 ) , .A( u1_R13_13 ) , .Z( u1_u14_X_18 ) );
  XOR2_X1 u1_u14_U41 (.B( u1_K15_17 ) , .A( u1_R13_12 ) , .Z( u1_u14_X_17 ) );
  XOR2_X1 u1_u14_U42 (.B( u1_K15_16 ) , .A( u1_R13_11 ) , .Z( u1_u14_X_16 ) );
  XOR2_X1 u1_u14_U43 (.B( u1_K15_15 ) , .A( u1_R13_10 ) , .Z( u1_u14_X_15 ) );
  XOR2_X1 u1_u14_U44 (.B( u1_K15_14 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_14 ) );
  XOR2_X1 u1_u14_U45 (.B( u1_K15_13 ) , .A( u1_R13_8 ) , .Z( u1_u14_X_13 ) );
  XOR2_X1 u1_u14_U46 (.B( u1_K15_12 ) , .A( u1_R13_9 ) , .Z( u1_u14_X_12 ) );
  XOR2_X1 u1_u14_U47 (.B( u1_K15_11 ) , .A( u1_R13_8 ) , .Z( u1_u14_X_11 ) );
  XOR2_X1 u1_u14_U5 (.B( u1_K15_5 ) , .A( u1_R13_4 ) , .Z( u1_u14_X_5 ) );
  XOR2_X1 u1_u14_U7 (.B( u1_K15_48 ) , .A( u1_R13_1 ) , .Z( u1_u14_X_48 ) );
  XOR2_X1 u1_u14_U8 (.B( u1_K15_47 ) , .A( u1_R13_32 ) , .Z( u1_u14_X_47 ) );
  XOR2_X1 u1_u14_U9 (.B( u1_K15_46 ) , .A( u1_R13_31 ) , .Z( u1_u14_X_46 ) );
  OAI22_X1 u1_u14_u2_U10 (.ZN( u1_u14_u2_n109 ) , .A2( u1_u14_u2_n113 ) , .B2( u1_u14_u2_n133 ) , .B1( u1_u14_u2_n167 ) , .A1( u1_u14_u2_n168 ) );
  NAND3_X1 u1_u14_u2_U100 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n98 ) );
  OAI22_X1 u1_u14_u2_U11 (.B1( u1_u14_u2_n151 ) , .A2( u1_u14_u2_n152 ) , .A1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n160 ) , .B2( u1_u14_u2_n168 ) );
  NOR3_X1 u1_u14_u2_U12 (.A1( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n151 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U13 (.ZN( u1_u14_u2_n144 ) , .B2( u1_u14_u2_n155 ) , .A( u1_u14_u2_n172 ) , .B1( u1_u14_u2_n185 ) );
  AOI21_X1 u1_u14_u2_U14 (.B2( u1_u14_u2_n143 ) , .ZN( u1_u14_u2_n145 ) , .B1( u1_u14_u2_n152 ) , .A( u1_u14_u2_n171 ) );
  AOI21_X1 u1_u14_u2_U15 (.B2( u1_u14_u2_n120 ) , .B1( u1_u14_u2_n121 ) , .ZN( u1_u14_u2_n126 ) , .A( u1_u14_u2_n167 ) );
  INV_X1 u1_u14_u2_U16 (.A( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n171 ) );
  INV_X1 u1_u14_u2_U17 (.A( u1_u14_u2_n120 ) , .ZN( u1_u14_u2_n188 ) );
  NAND2_X1 u1_u14_u2_U18 (.A2( u1_u14_u2_n122 ) , .ZN( u1_u14_u2_n150 ) , .A1( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U19 (.A( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U20 (.A( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n173 ) );
  NAND2_X1 u1_u14_u2_U21 (.A1( u1_u14_u2_n132 ) , .A2( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n157 ) );
  INV_X1 u1_u14_u2_U22 (.A( u1_u14_u2_n113 ) , .ZN( u1_u14_u2_n178 ) );
  INV_X1 u1_u14_u2_U23 (.A( u1_u14_u2_n139 ) , .ZN( u1_u14_u2_n175 ) );
  INV_X1 u1_u14_u2_U24 (.A( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U25 (.A( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n177 ) );
  INV_X1 u1_u14_u2_U26 (.A( u1_u14_u2_n116 ) , .ZN( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U27 (.A( u1_u14_u2_n131 ) , .ZN( u1_u14_u2_n179 ) );
  INV_X1 u1_u14_u2_U28 (.A( u1_u14_u2_n154 ) , .ZN( u1_u14_u2_n176 ) );
  NAND2_X1 u1_u14_u2_U29 (.A2( u1_u14_u2_n116 ) , .A1( u1_u14_u2_n117 ) , .ZN( u1_u14_u2_n118 ) );
  NOR2_X1 u1_u14_u2_U3 (.ZN( u1_u14_u2_n121 ) , .A2( u1_u14_u2_n177 ) , .A1( u1_u14_u2_n180 ) );
  INV_X1 u1_u14_u2_U30 (.A( u1_u14_u2_n132 ) , .ZN( u1_u14_u2_n182 ) );
  INV_X1 u1_u14_u2_U31 (.A( u1_u14_u2_n158 ) , .ZN( u1_u14_u2_n183 ) );
  OAI21_X1 u1_u14_u2_U32 (.A( u1_u14_u2_n156 ) , .B1( u1_u14_u2_n157 ) , .ZN( u1_u14_u2_n158 ) , .B2( u1_u14_u2_n179 ) );
  NOR2_X1 u1_u14_u2_U33 (.ZN( u1_u14_u2_n156 ) , .A1( u1_u14_u2_n166 ) , .A2( u1_u14_u2_n169 ) );
  NOR2_X1 u1_u14_u2_U34 (.A2( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n140 ) );
  NOR2_X1 u1_u14_u2_U35 (.A2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n153 ) , .A1( u1_u14_u2_n156 ) );
  AOI211_X1 u1_u14_u2_U36 (.ZN( u1_u14_u2_n130 ) , .C1( u1_u14_u2_n138 ) , .C2( u1_u14_u2_n179 ) , .B( u1_u14_u2_n96 ) , .A( u1_u14_u2_n97 ) );
  OAI22_X1 u1_u14_u2_U37 (.B1( u1_u14_u2_n133 ) , .A2( u1_u14_u2_n137 ) , .A1( u1_u14_u2_n152 ) , .B2( u1_u14_u2_n168 ) , .ZN( u1_u14_u2_n97 ) );
  OAI221_X1 u1_u14_u2_U38 (.B1( u1_u14_u2_n113 ) , .C1( u1_u14_u2_n132 ) , .A( u1_u14_u2_n149 ) , .B2( u1_u14_u2_n171 ) , .C2( u1_u14_u2_n172 ) , .ZN( u1_u14_u2_n96 ) );
  OAI221_X1 u1_u14_u2_U39 (.A( u1_u14_u2_n115 ) , .C2( u1_u14_u2_n123 ) , .B2( u1_u14_u2_n143 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n163 ) , .C1( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U4 (.A( u1_u14_u2_n134 ) , .ZN( u1_u14_u2_n185 ) );
  OAI21_X1 u1_u14_u2_U40 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n115 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n178 ) );
  OAI221_X1 u1_u14_u2_U41 (.A( u1_u14_u2_n135 ) , .B2( u1_u14_u2_n136 ) , .B1( u1_u14_u2_n137 ) , .ZN( u1_u14_u2_n162 ) , .C2( u1_u14_u2_n167 ) , .C1( u1_u14_u2_n185 ) );
  AND3_X1 u1_u14_u2_U42 (.A3( u1_u14_u2_n131 ) , .A2( u1_u14_u2_n132 ) , .A1( u1_u14_u2_n133 ) , .ZN( u1_u14_u2_n136 ) );
  AOI22_X1 u1_u14_u2_U43 (.ZN( u1_u14_u2_n135 ) , .B1( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n156 ) , .B2( u1_u14_u2_n180 ) , .A2( u1_u14_u2_n188 ) );
  AOI21_X1 u1_u14_u2_U44 (.ZN( u1_u14_u2_n149 ) , .B1( u1_u14_u2_n173 ) , .B2( u1_u14_u2_n188 ) , .A( u1_u14_u2_n95 ) );
  AND3_X1 u1_u14_u2_U45 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n156 ) , .ZN( u1_u14_u2_n95 ) );
  OAI21_X1 u1_u14_u2_U46 (.A( u1_u14_u2_n101 ) , .B2( u1_u14_u2_n121 ) , .B1( u1_u14_u2_n153 ) , .ZN( u1_u14_u2_n164 ) );
  NAND2_X1 u1_u14_u2_U47 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n155 ) );
  NAND2_X1 u1_u14_u2_U48 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n143 ) );
  NAND2_X1 u1_u14_u2_U49 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n152 ) );
  INV_X1 u1_u14_u2_U5 (.A( u1_u14_u2_n150 ) , .ZN( u1_u14_u2_n184 ) );
  NAND2_X1 u1_u14_u2_U50 (.A1( u1_u14_u2_n100 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n132 ) );
  INV_X1 u1_u14_u2_U51 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n168 ) );
  INV_X1 u1_u14_u2_U52 (.A( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n167 ) );
  OAI21_X1 u1_u14_u2_U53 (.A( u1_u14_u2_n141 ) , .B2( u1_u14_u2_n142 ) , .ZN( u1_u14_u2_n146 ) , .B1( u1_u14_u2_n153 ) );
  OAI21_X1 u1_u14_u2_U54 (.A( u1_u14_u2_n140 ) , .ZN( u1_u14_u2_n141 ) , .B1( u1_u14_u2_n176 ) , .B2( u1_u14_u2_n177 ) );
  NOR3_X1 u1_u14_u2_U55 (.ZN( u1_u14_u2_n142 ) , .A3( u1_u14_u2_n175 ) , .A2( u1_u14_u2_n178 ) , .A1( u1_u14_u2_n181 ) );
  INV_X1 u1_u14_u2_U56 (.ZN( u1_u14_u2_n187 ) , .A( u1_u14_u2_n99 ) );
  OAI21_X1 u1_u14_u2_U57 (.B1( u1_u14_u2_n137 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n98 ) , .ZN( u1_u14_u2_n99 ) );
  NAND2_X1 u1_u14_u2_U58 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n113 ) );
  NAND2_X1 u1_u14_u2_U59 (.A1( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n131 ) );
  NOR4_X1 u1_u14_u2_U6 (.A4( u1_u14_u2_n124 ) , .A3( u1_u14_u2_n125 ) , .A2( u1_u14_u2_n126 ) , .A1( u1_u14_u2_n127 ) , .ZN( u1_u14_u2_n128 ) );
  NAND2_X1 u1_u14_u2_U60 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n107 ) , .ZN( u1_u14_u2_n139 ) );
  NAND2_X1 u1_u14_u2_U61 (.A1( u1_u14_u2_n103 ) , .A2( u1_u14_u2_n105 ) , .ZN( u1_u14_u2_n133 ) );
  NAND2_X1 u1_u14_u2_U62 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n103 ) , .ZN( u1_u14_u2_n154 ) );
  NAND2_X1 u1_u14_u2_U63 (.A2( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n104 ) , .ZN( u1_u14_u2_n119 ) );
  NAND2_X1 u1_u14_u2_U64 (.A2( u1_u14_u2_n107 ) , .A1( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n123 ) );
  NAND2_X1 u1_u14_u2_U65 (.A1( u1_u14_u2_n104 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n122 ) );
  INV_X1 u1_u14_u2_U66 (.A( u1_u14_u2_n114 ) , .ZN( u1_u14_u2_n172 ) );
  NAND2_X1 u1_u14_u2_U67 (.A2( u1_u14_u2_n100 ) , .A1( u1_u14_u2_n102 ) , .ZN( u1_u14_u2_n116 ) );
  NAND2_X1 u1_u14_u2_U68 (.A1( u1_u14_u2_n102 ) , .A2( u1_u14_u2_n108 ) , .ZN( u1_u14_u2_n120 ) );
  NAND2_X1 u1_u14_u2_U69 (.A2( u1_u14_u2_n105 ) , .A1( u1_u14_u2_n106 ) , .ZN( u1_u14_u2_n117 ) );
  AOI21_X1 u1_u14_u2_U7 (.B2( u1_u14_u2_n119 ) , .ZN( u1_u14_u2_n127 ) , .A( u1_u14_u2_n137 ) , .B1( u1_u14_u2_n155 ) );
  NOR2_X1 u1_u14_u2_U70 (.A2( u1_u14_X_16 ) , .ZN( u1_u14_u2_n140 ) , .A1( u1_u14_u2_n166 ) );
  NOR2_X1 u1_u14_u2_U71 (.A2( u1_u14_X_13 ) , .A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n100 ) );
  NOR2_X1 u1_u14_u2_U72 (.A2( u1_u14_X_16 ) , .A1( u1_u14_X_17 ) , .ZN( u1_u14_u2_n138 ) );
  NOR2_X1 u1_u14_u2_U73 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n104 ) );
  NOR2_X1 u1_u14_u2_U74 (.A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n103 ) , .A1( u1_u14_u2_n174 ) );
  NOR2_X1 u1_u14_u2_U75 (.A2( u1_u14_X_15 ) , .ZN( u1_u14_u2_n102 ) , .A1( u1_u14_u2_n165 ) );
  NOR2_X1 u1_u14_u2_U76 (.A2( u1_u14_X_17 ) , .ZN( u1_u14_u2_n114 ) , .A1( u1_u14_u2_n169 ) );
  AND2_X1 u1_u14_u2_U77 (.A1( u1_u14_X_15 ) , .ZN( u1_u14_u2_n105 ) , .A2( u1_u14_u2_n165 ) );
  AND2_X1 u1_u14_u2_U78 (.A2( u1_u14_X_15 ) , .A1( u1_u14_X_18 ) , .ZN( u1_u14_u2_n107 ) );
  AND2_X1 u1_u14_u2_U79 (.A1( u1_u14_X_14 ) , .ZN( u1_u14_u2_n106 ) , .A2( u1_u14_u2_n174 ) );
  AOI21_X1 u1_u14_u2_U8 (.ZN( u1_u14_u2_n124 ) , .B1( u1_u14_u2_n131 ) , .B2( u1_u14_u2_n143 ) , .A( u1_u14_u2_n172 ) );
  AND2_X1 u1_u14_u2_U80 (.A1( u1_u14_X_13 ) , .A2( u1_u14_X_14 ) , .ZN( u1_u14_u2_n108 ) );
  INV_X1 u1_u14_u2_U81 (.A( u1_u14_X_16 ) , .ZN( u1_u14_u2_n169 ) );
  INV_X1 u1_u14_u2_U82 (.A( u1_u14_X_17 ) , .ZN( u1_u14_u2_n166 ) );
  INV_X1 u1_u14_u2_U83 (.A( u1_u14_X_13 ) , .ZN( u1_u14_u2_n174 ) );
  INV_X1 u1_u14_u2_U84 (.A( u1_u14_X_18 ) , .ZN( u1_u14_u2_n165 ) );
  NAND4_X1 u1_u14_u2_U85 (.ZN( u1_out14_30 ) , .A4( u1_u14_u2_n147 ) , .A3( u1_u14_u2_n148 ) , .A2( u1_u14_u2_n149 ) , .A1( u1_u14_u2_n187 ) );
  NOR3_X1 u1_u14_u2_U86 (.A3( u1_u14_u2_n144 ) , .A2( u1_u14_u2_n145 ) , .A1( u1_u14_u2_n146 ) , .ZN( u1_u14_u2_n147 ) );
  AOI21_X1 u1_u14_u2_U87 (.B2( u1_u14_u2_n138 ) , .ZN( u1_u14_u2_n148 ) , .A( u1_u14_u2_n162 ) , .B1( u1_u14_u2_n182 ) );
  NAND4_X1 u1_u14_u2_U88 (.ZN( u1_out14_24 ) , .A4( u1_u14_u2_n111 ) , .A3( u1_u14_u2_n112 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n187 ) );
  AOI221_X1 u1_u14_u2_U89 (.A( u1_u14_u2_n109 ) , .B1( u1_u14_u2_n110 ) , .ZN( u1_u14_u2_n111 ) , .C1( u1_u14_u2_n134 ) , .C2( u1_u14_u2_n170 ) , .B2( u1_u14_u2_n173 ) );
  AOI21_X1 u1_u14_u2_U9 (.B2( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n125 ) , .A( u1_u14_u2_n171 ) , .B1( u1_u14_u2_n184 ) );
  AOI21_X1 u1_u14_u2_U90 (.ZN( u1_u14_u2_n112 ) , .B2( u1_u14_u2_n156 ) , .A( u1_u14_u2_n164 ) , .B1( u1_u14_u2_n181 ) );
  NAND4_X1 u1_u14_u2_U91 (.ZN( u1_out14_16 ) , .A4( u1_u14_u2_n128 ) , .A3( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n130 ) , .A2( u1_u14_u2_n186 ) );
  AOI22_X1 u1_u14_u2_U92 (.A2( u1_u14_u2_n118 ) , .ZN( u1_u14_u2_n129 ) , .A1( u1_u14_u2_n140 ) , .B1( u1_u14_u2_n157 ) , .B2( u1_u14_u2_n170 ) );
  INV_X1 u1_u14_u2_U93 (.A( u1_u14_u2_n163 ) , .ZN( u1_u14_u2_n186 ) );
  OR4_X1 u1_u14_u2_U94 (.ZN( u1_out14_6 ) , .A4( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n162 ) , .A2( u1_u14_u2_n163 ) , .A1( u1_u14_u2_n164 ) );
  OR3_X1 u1_u14_u2_U95 (.A2( u1_u14_u2_n159 ) , .A1( u1_u14_u2_n160 ) , .ZN( u1_u14_u2_n161 ) , .A3( u1_u14_u2_n183 ) );
  AOI21_X1 u1_u14_u2_U96 (.B2( u1_u14_u2_n154 ) , .B1( u1_u14_u2_n155 ) , .ZN( u1_u14_u2_n159 ) , .A( u1_u14_u2_n167 ) );
  NAND3_X1 u1_u14_u2_U97 (.A2( u1_u14_u2_n117 ) , .A1( u1_u14_u2_n122 ) , .A3( u1_u14_u2_n123 ) , .ZN( u1_u14_u2_n134 ) );
  NAND3_X1 u1_u14_u2_U98 (.ZN( u1_u14_u2_n110 ) , .A2( u1_u14_u2_n131 ) , .A3( u1_u14_u2_n139 ) , .A1( u1_u14_u2_n154 ) );
  NAND3_X1 u1_u14_u2_U99 (.A2( u1_u14_u2_n100 ) , .ZN( u1_u14_u2_n101 ) , .A1( u1_u14_u2_n104 ) , .A3( u1_u14_u2_n114 ) );
  INV_X1 u1_u14_u5_U10 (.A( u1_u14_u5_n121 ) , .ZN( u1_u14_u5_n177 ) );
  NOR3_X1 u1_u14_u5_U100 (.A3( u1_u14_u5_n141 ) , .A1( u1_u14_u5_n142 ) , .ZN( u1_u14_u5_n143 ) , .A2( u1_u14_u5_n191 ) );
  NAND4_X1 u1_u14_u5_U101 (.ZN( u1_out14_4 ) , .A4( u1_u14_u5_n112 ) , .A2( u1_u14_u5_n113 ) , .A1( u1_u14_u5_n114 ) , .A3( u1_u14_u5_n195 ) );
  AOI211_X1 u1_u14_u5_U102 (.A( u1_u14_u5_n110 ) , .C1( u1_u14_u5_n111 ) , .ZN( u1_u14_u5_n112 ) , .B( u1_u14_u5_n118 ) , .C2( u1_u14_u5_n177 ) );
  AOI222_X1 u1_u14_u5_U103 (.ZN( u1_u14_u5_n113 ) , .A1( u1_u14_u5_n131 ) , .C1( u1_u14_u5_n148 ) , .B2( u1_u14_u5_n174 ) , .C2( u1_u14_u5_n178 ) , .A2( u1_u14_u5_n179 ) , .B1( u1_u14_u5_n99 ) );
  NAND3_X1 u1_u14_u5_U104 (.A2( u1_u14_u5_n154 ) , .A3( u1_u14_u5_n158 ) , .A1( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n99 ) );
  NOR2_X1 u1_u14_u5_U11 (.ZN( u1_u14_u5_n160 ) , .A2( u1_u14_u5_n173 ) , .A1( u1_u14_u5_n177 ) );
  INV_X1 u1_u14_u5_U12 (.A( u1_u14_u5_n150 ) , .ZN( u1_u14_u5_n174 ) );
  AOI21_X1 u1_u14_u5_U13 (.A( u1_u14_u5_n160 ) , .B2( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n162 ) , .B1( u1_u14_u5_n192 ) );
  INV_X1 u1_u14_u5_U14 (.A( u1_u14_u5_n159 ) , .ZN( u1_u14_u5_n192 ) );
  AOI21_X1 u1_u14_u5_U15 (.A( u1_u14_u5_n156 ) , .B2( u1_u14_u5_n157 ) , .B1( u1_u14_u5_n158 ) , .ZN( u1_u14_u5_n163 ) );
  AOI21_X1 u1_u14_u5_U16 (.B2( u1_u14_u5_n139 ) , .B1( u1_u14_u5_n140 ) , .ZN( u1_u14_u5_n141 ) , .A( u1_u14_u5_n150 ) );
  OAI21_X1 u1_u14_u5_U17 (.A( u1_u14_u5_n133 ) , .B2( u1_u14_u5_n134 ) , .B1( u1_u14_u5_n135 ) , .ZN( u1_u14_u5_n142 ) );
  OAI21_X1 u1_u14_u5_U18 (.ZN( u1_u14_u5_n133 ) , .B2( u1_u14_u5_n147 ) , .A( u1_u14_u5_n173 ) , .B1( u1_u14_u5_n188 ) );
  NAND2_X1 u1_u14_u5_U19 (.A2( u1_u14_u5_n119 ) , .A1( u1_u14_u5_n123 ) , .ZN( u1_u14_u5_n137 ) );
  INV_X1 u1_u14_u5_U20 (.A( u1_u14_u5_n155 ) , .ZN( u1_u14_u5_n194 ) );
  NAND2_X1 u1_u14_u5_U21 (.A1( u1_u14_u5_n121 ) , .ZN( u1_u14_u5_n132 ) , .A2( u1_u14_u5_n172 ) );
  NAND2_X1 u1_u14_u5_U22 (.A2( u1_u14_u5_n122 ) , .ZN( u1_u14_u5_n136 ) , .A1( u1_u14_u5_n154 ) );
  NAND2_X1 u1_u14_u5_U23 (.A2( u1_u14_u5_n119 ) , .A1( u1_u14_u5_n120 ) , .ZN( u1_u14_u5_n159 ) );
  INV_X1 u1_u14_u5_U24 (.A( u1_u14_u5_n156 ) , .ZN( u1_u14_u5_n175 ) );
  INV_X1 u1_u14_u5_U25 (.A( u1_u14_u5_n158 ) , .ZN( u1_u14_u5_n188 ) );
  INV_X1 u1_u14_u5_U26 (.A( u1_u14_u5_n152 ) , .ZN( u1_u14_u5_n179 ) );
  INV_X1 u1_u14_u5_U27 (.A( u1_u14_u5_n140 ) , .ZN( u1_u14_u5_n182 ) );
  INV_X1 u1_u14_u5_U28 (.A( u1_u14_u5_n151 ) , .ZN( u1_u14_u5_n183 ) );
  INV_X1 u1_u14_u5_U29 (.A( u1_u14_u5_n123 ) , .ZN( u1_u14_u5_n185 ) );
  NOR2_X1 u1_u14_u5_U3 (.ZN( u1_u14_u5_n134 ) , .A1( u1_u14_u5_n183 ) , .A2( u1_u14_u5_n190 ) );
  INV_X1 u1_u14_u5_U30 (.A( u1_u14_u5_n161 ) , .ZN( u1_u14_u5_n184 ) );
  INV_X1 u1_u14_u5_U31 (.A( u1_u14_u5_n139 ) , .ZN( u1_u14_u5_n189 ) );
  INV_X1 u1_u14_u5_U32 (.A( u1_u14_u5_n157 ) , .ZN( u1_u14_u5_n190 ) );
  INV_X1 u1_u14_u5_U33 (.A( u1_u14_u5_n120 ) , .ZN( u1_u14_u5_n193 ) );
  NAND2_X1 u1_u14_u5_U34 (.ZN( u1_u14_u5_n111 ) , .A1( u1_u14_u5_n140 ) , .A2( u1_u14_u5_n155 ) );
  INV_X1 u1_u14_u5_U35 (.A( u1_u14_u5_n117 ) , .ZN( u1_u14_u5_n196 ) );
  OAI221_X1 u1_u14_u5_U36 (.A( u1_u14_u5_n116 ) , .ZN( u1_u14_u5_n117 ) , .B2( u1_u14_u5_n119 ) , .C1( u1_u14_u5_n153 ) , .C2( u1_u14_u5_n158 ) , .B1( u1_u14_u5_n172 ) );
  AOI222_X1 u1_u14_u5_U37 (.ZN( u1_u14_u5_n116 ) , .B2( u1_u14_u5_n145 ) , .C1( u1_u14_u5_n148 ) , .A2( u1_u14_u5_n174 ) , .C2( u1_u14_u5_n177 ) , .B1( u1_u14_u5_n187 ) , .A1( u1_u14_u5_n193 ) );
  INV_X1 u1_u14_u5_U38 (.A( u1_u14_u5_n115 ) , .ZN( u1_u14_u5_n187 ) );
  NOR2_X1 u1_u14_u5_U39 (.ZN( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n170 ) , .A2( u1_u14_u5_n180 ) );
  INV_X1 u1_u14_u5_U4 (.A( u1_u14_u5_n138 ) , .ZN( u1_u14_u5_n191 ) );
  AOI22_X1 u1_u14_u5_U40 (.B2( u1_u14_u5_n131 ) , .A2( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n169 ) , .B1( u1_u14_u5_n174 ) , .A1( u1_u14_u5_n185 ) );
  NOR2_X1 u1_u14_u5_U41 (.A1( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n150 ) , .A2( u1_u14_u5_n173 ) );
  AOI21_X1 u1_u14_u5_U42 (.A( u1_u14_u5_n118 ) , .B2( u1_u14_u5_n145 ) , .ZN( u1_u14_u5_n168 ) , .B1( u1_u14_u5_n186 ) );
  INV_X1 u1_u14_u5_U43 (.A( u1_u14_u5_n122 ) , .ZN( u1_u14_u5_n186 ) );
  NOR2_X1 u1_u14_u5_U44 (.A1( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n152 ) , .A2( u1_u14_u5_n176 ) );
  NOR2_X1 u1_u14_u5_U45 (.A1( u1_u14_u5_n115 ) , .ZN( u1_u14_u5_n118 ) , .A2( u1_u14_u5_n153 ) );
  NOR2_X1 u1_u14_u5_U46 (.A2( u1_u14_u5_n145 ) , .ZN( u1_u14_u5_n156 ) , .A1( u1_u14_u5_n174 ) );
  NOR2_X1 u1_u14_u5_U47 (.ZN( u1_u14_u5_n121 ) , .A2( u1_u14_u5_n145 ) , .A1( u1_u14_u5_n176 ) );
  AOI22_X1 u1_u14_u5_U48 (.ZN( u1_u14_u5_n114 ) , .A2( u1_u14_u5_n137 ) , .A1( u1_u14_u5_n145 ) , .B2( u1_u14_u5_n175 ) , .B1( u1_u14_u5_n193 ) );
  OAI211_X1 u1_u14_u5_U49 (.B( u1_u14_u5_n124 ) , .A( u1_u14_u5_n125 ) , .C2( u1_u14_u5_n126 ) , .C1( u1_u14_u5_n127 ) , .ZN( u1_u14_u5_n128 ) );
  OAI21_X1 u1_u14_u5_U5 (.B2( u1_u14_u5_n136 ) , .B1( u1_u14_u5_n137 ) , .ZN( u1_u14_u5_n138 ) , .A( u1_u14_u5_n177 ) );
  NOR3_X1 u1_u14_u5_U50 (.ZN( u1_u14_u5_n127 ) , .A1( u1_u14_u5_n136 ) , .A3( u1_u14_u5_n148 ) , .A2( u1_u14_u5_n182 ) );
  OAI21_X1 u1_u14_u5_U51 (.ZN( u1_u14_u5_n124 ) , .A( u1_u14_u5_n177 ) , .B2( u1_u14_u5_n183 ) , .B1( u1_u14_u5_n189 ) );
  OAI21_X1 u1_u14_u5_U52 (.ZN( u1_u14_u5_n125 ) , .A( u1_u14_u5_n174 ) , .B2( u1_u14_u5_n185 ) , .B1( u1_u14_u5_n190 ) );
  AOI21_X1 u1_u14_u5_U53 (.A( u1_u14_u5_n153 ) , .B2( u1_u14_u5_n154 ) , .B1( u1_u14_u5_n155 ) , .ZN( u1_u14_u5_n164 ) );
  AOI21_X1 u1_u14_u5_U54 (.ZN( u1_u14_u5_n110 ) , .B1( u1_u14_u5_n122 ) , .B2( u1_u14_u5_n139 ) , .A( u1_u14_u5_n153 ) );
  INV_X1 u1_u14_u5_U55 (.A( u1_u14_u5_n153 ) , .ZN( u1_u14_u5_n176 ) );
  INV_X1 u1_u14_u5_U56 (.A( u1_u14_u5_n126 ) , .ZN( u1_u14_u5_n173 ) );
  AND2_X1 u1_u14_u5_U57 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n147 ) );
  AND2_X1 u1_u14_u5_U58 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n148 ) );
  NAND2_X1 u1_u14_u5_U59 (.A1( u1_u14_u5_n105 ) , .A2( u1_u14_u5_n106 ) , .ZN( u1_u14_u5_n158 ) );
  INV_X1 u1_u14_u5_U6 (.A( u1_u14_u5_n135 ) , .ZN( u1_u14_u5_n178 ) );
  NAND2_X1 u1_u14_u5_U60 (.A2( u1_u14_u5_n108 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n139 ) );
  NAND2_X1 u1_u14_u5_U61 (.A1( u1_u14_u5_n106 ) , .A2( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n119 ) );
  NAND2_X1 u1_u14_u5_U62 (.A2( u1_u14_u5_n103 ) , .A1( u1_u14_u5_n105 ) , .ZN( u1_u14_u5_n140 ) );
  NAND2_X1 u1_u14_u5_U63 (.A2( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n105 ) , .ZN( u1_u14_u5_n155 ) );
  NAND2_X1 u1_u14_u5_U64 (.A2( u1_u14_u5_n106 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n122 ) );
  NAND2_X1 u1_u14_u5_U65 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n106 ) , .ZN( u1_u14_u5_n115 ) );
  NAND2_X1 u1_u14_u5_U66 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n103 ) , .ZN( u1_u14_u5_n161 ) );
  NAND2_X1 u1_u14_u5_U67 (.A1( u1_u14_u5_n105 ) , .A2( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n154 ) );
  INV_X1 u1_u14_u5_U68 (.A( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n172 ) );
  NAND2_X1 u1_u14_u5_U69 (.A1( u1_u14_u5_n103 ) , .A2( u1_u14_u5_n108 ) , .ZN( u1_u14_u5_n123 ) );
  OAI22_X1 u1_u14_u5_U7 (.B2( u1_u14_u5_n149 ) , .B1( u1_u14_u5_n150 ) , .A2( u1_u14_u5_n151 ) , .A1( u1_u14_u5_n152 ) , .ZN( u1_u14_u5_n165 ) );
  NAND2_X1 u1_u14_u5_U70 (.A2( u1_u14_u5_n103 ) , .A1( u1_u14_u5_n107 ) , .ZN( u1_u14_u5_n151 ) );
  NAND2_X1 u1_u14_u5_U71 (.A2( u1_u14_u5_n107 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n120 ) );
  NAND2_X1 u1_u14_u5_U72 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n109 ) , .ZN( u1_u14_u5_n157 ) );
  AND2_X1 u1_u14_u5_U73 (.A2( u1_u14_u5_n100 ) , .A1( u1_u14_u5_n104 ) , .ZN( u1_u14_u5_n131 ) );
  INV_X1 u1_u14_u5_U74 (.A( u1_u14_u5_n102 ) , .ZN( u1_u14_u5_n195 ) );
  OAI221_X1 u1_u14_u5_U75 (.A( u1_u14_u5_n101 ) , .ZN( u1_u14_u5_n102 ) , .C2( u1_u14_u5_n115 ) , .C1( u1_u14_u5_n126 ) , .B1( u1_u14_u5_n134 ) , .B2( u1_u14_u5_n160 ) );
  OAI21_X1 u1_u14_u5_U76 (.ZN( u1_u14_u5_n101 ) , .B1( u1_u14_u5_n137 ) , .A( u1_u14_u5_n146 ) , .B2( u1_u14_u5_n147 ) );
  NOR2_X1 u1_u14_u5_U77 (.A2( u1_u14_X_34 ) , .A1( u1_u14_X_35 ) , .ZN( u1_u14_u5_n145 ) );
  NOR2_X1 u1_u14_u5_U78 (.A2( u1_u14_X_34 ) , .ZN( u1_u14_u5_n146 ) , .A1( u1_u14_u5_n171 ) );
  NOR2_X1 u1_u14_u5_U79 (.A2( u1_u14_X_31 ) , .A1( u1_u14_X_32 ) , .ZN( u1_u14_u5_n103 ) );
  NOR3_X1 u1_u14_u5_U8 (.A2( u1_u14_u5_n147 ) , .A1( u1_u14_u5_n148 ) , .ZN( u1_u14_u5_n149 ) , .A3( u1_u14_u5_n194 ) );
  NOR2_X1 u1_u14_u5_U80 (.A2( u1_u14_X_36 ) , .ZN( u1_u14_u5_n105 ) , .A1( u1_u14_u5_n180 ) );
  NOR2_X1 u1_u14_u5_U81 (.A2( u1_u14_X_33 ) , .ZN( u1_u14_u5_n108 ) , .A1( u1_u14_u5_n170 ) );
  NOR2_X1 u1_u14_u5_U82 (.A2( u1_u14_X_33 ) , .A1( u1_u14_X_36 ) , .ZN( u1_u14_u5_n107 ) );
  NOR2_X1 u1_u14_u5_U83 (.A2( u1_u14_X_31 ) , .ZN( u1_u14_u5_n104 ) , .A1( u1_u14_u5_n181 ) );
  NAND2_X1 u1_u14_u5_U84 (.A2( u1_u14_X_34 ) , .A1( u1_u14_X_35 ) , .ZN( u1_u14_u5_n153 ) );
  NAND2_X1 u1_u14_u5_U85 (.A1( u1_u14_X_34 ) , .ZN( u1_u14_u5_n126 ) , .A2( u1_u14_u5_n171 ) );
  AND2_X1 u1_u14_u5_U86 (.A1( u1_u14_X_31 ) , .A2( u1_u14_X_32 ) , .ZN( u1_u14_u5_n106 ) );
  AND2_X1 u1_u14_u5_U87 (.A1( u1_u14_X_31 ) , .ZN( u1_u14_u5_n109 ) , .A2( u1_u14_u5_n181 ) );
  INV_X1 u1_u14_u5_U88 (.A( u1_u14_X_33 ) , .ZN( u1_u14_u5_n180 ) );
  INV_X1 u1_u14_u5_U89 (.A( u1_u14_X_35 ) , .ZN( u1_u14_u5_n171 ) );
  NOR2_X1 u1_u14_u5_U9 (.ZN( u1_u14_u5_n135 ) , .A1( u1_u14_u5_n173 ) , .A2( u1_u14_u5_n176 ) );
  INV_X1 u1_u14_u5_U90 (.A( u1_u14_X_36 ) , .ZN( u1_u14_u5_n170 ) );
  INV_X1 u1_u14_u5_U91 (.A( u1_u14_X_32 ) , .ZN( u1_u14_u5_n181 ) );
  NAND4_X1 u1_u14_u5_U92 (.ZN( u1_out14_29 ) , .A4( u1_u14_u5_n129 ) , .A3( u1_u14_u5_n130 ) , .A2( u1_u14_u5_n168 ) , .A1( u1_u14_u5_n196 ) );
  AOI221_X1 u1_u14_u5_U93 (.A( u1_u14_u5_n128 ) , .ZN( u1_u14_u5_n129 ) , .C2( u1_u14_u5_n132 ) , .B2( u1_u14_u5_n159 ) , .B1( u1_u14_u5_n176 ) , .C1( u1_u14_u5_n184 ) );
  AOI222_X1 u1_u14_u5_U94 (.ZN( u1_u14_u5_n130 ) , .A2( u1_u14_u5_n146 ) , .B1( u1_u14_u5_n147 ) , .C2( u1_u14_u5_n175 ) , .B2( u1_u14_u5_n179 ) , .A1( u1_u14_u5_n188 ) , .C1( u1_u14_u5_n194 ) );
  NAND4_X1 u1_u14_u5_U95 (.ZN( u1_out14_19 ) , .A4( u1_u14_u5_n166 ) , .A3( u1_u14_u5_n167 ) , .A2( u1_u14_u5_n168 ) , .A1( u1_u14_u5_n169 ) );
  AOI22_X1 u1_u14_u5_U96 (.B2( u1_u14_u5_n145 ) , .A2( u1_u14_u5_n146 ) , .ZN( u1_u14_u5_n167 ) , .B1( u1_u14_u5_n182 ) , .A1( u1_u14_u5_n189 ) );
  NOR4_X1 u1_u14_u5_U97 (.A4( u1_u14_u5_n162 ) , .A3( u1_u14_u5_n163 ) , .A2( u1_u14_u5_n164 ) , .A1( u1_u14_u5_n165 ) , .ZN( u1_u14_u5_n166 ) );
  NAND4_X1 u1_u14_u5_U98 (.ZN( u1_out14_11 ) , .A4( u1_u14_u5_n143 ) , .A3( u1_u14_u5_n144 ) , .A2( u1_u14_u5_n169 ) , .A1( u1_u14_u5_n196 ) );
  AOI22_X1 u1_u14_u5_U99 (.A2( u1_u14_u5_n132 ) , .ZN( u1_u14_u5_n144 ) , .B2( u1_u14_u5_n145 ) , .B1( u1_u14_u5_n184 ) , .A1( u1_u14_u5_n194 ) );
  AOI22_X1 u1_u14_u6_U10 (.A2( u1_u14_u6_n151 ) , .B2( u1_u14_u6_n161 ) , .A1( u1_u14_u6_n167 ) , .B1( u1_u14_u6_n170 ) , .ZN( u1_u14_u6_n89 ) );
  AOI21_X1 u1_u14_u6_U11 (.B1( u1_u14_u6_n107 ) , .B2( u1_u14_u6_n132 ) , .A( u1_u14_u6_n158 ) , .ZN( u1_u14_u6_n88 ) );
  AOI21_X1 u1_u14_u6_U12 (.B2( u1_u14_u6_n147 ) , .B1( u1_u14_u6_n148 ) , .ZN( u1_u14_u6_n149 ) , .A( u1_u14_u6_n158 ) );
  AOI21_X1 u1_u14_u6_U13 (.ZN( u1_u14_u6_n106 ) , .A( u1_u14_u6_n142 ) , .B2( u1_u14_u6_n159 ) , .B1( u1_u14_u6_n164 ) );
  INV_X1 u1_u14_u6_U14 (.A( u1_u14_u6_n155 ) , .ZN( u1_u14_u6_n161 ) );
  INV_X1 u1_u14_u6_U15 (.A( u1_u14_u6_n128 ) , .ZN( u1_u14_u6_n164 ) );
  NAND2_X1 u1_u14_u6_U16 (.ZN( u1_u14_u6_n110 ) , .A1( u1_u14_u6_n122 ) , .A2( u1_u14_u6_n129 ) );
  NAND2_X1 u1_u14_u6_U17 (.ZN( u1_u14_u6_n124 ) , .A2( u1_u14_u6_n146 ) , .A1( u1_u14_u6_n148 ) );
  INV_X1 u1_u14_u6_U18 (.A( u1_u14_u6_n132 ) , .ZN( u1_u14_u6_n171 ) );
  AND2_X1 u1_u14_u6_U19 (.A1( u1_u14_u6_n100 ) , .ZN( u1_u14_u6_n130 ) , .A2( u1_u14_u6_n147 ) );
  INV_X1 u1_u14_u6_U20 (.A( u1_u14_u6_n127 ) , .ZN( u1_u14_u6_n173 ) );
  INV_X1 u1_u14_u6_U21 (.A( u1_u14_u6_n121 ) , .ZN( u1_u14_u6_n167 ) );
  INV_X1 u1_u14_u6_U22 (.A( u1_u14_u6_n100 ) , .ZN( u1_u14_u6_n169 ) );
  INV_X1 u1_u14_u6_U23 (.A( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n170 ) );
  INV_X1 u1_u14_u6_U24 (.A( u1_u14_u6_n113 ) , .ZN( u1_u14_u6_n168 ) );
  AND2_X1 u1_u14_u6_U25 (.A1( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n119 ) , .ZN( u1_u14_u6_n133 ) );
  AND2_X1 u1_u14_u6_U26 (.A2( u1_u14_u6_n121 ) , .A1( u1_u14_u6_n122 ) , .ZN( u1_u14_u6_n131 ) );
  AND3_X1 u1_u14_u6_U27 (.ZN( u1_u14_u6_n120 ) , .A2( u1_u14_u6_n127 ) , .A1( u1_u14_u6_n132 ) , .A3( u1_u14_u6_n145 ) );
  INV_X1 u1_u14_u6_U28 (.A( u1_u14_u6_n146 ) , .ZN( u1_u14_u6_n163 ) );
  AOI222_X1 u1_u14_u6_U29 (.ZN( u1_u14_u6_n114 ) , .A1( u1_u14_u6_n118 ) , .A2( u1_u14_u6_n126 ) , .B2( u1_u14_u6_n151 ) , .C2( u1_u14_u6_n159 ) , .C1( u1_u14_u6_n168 ) , .B1( u1_u14_u6_n169 ) );
  INV_X1 u1_u14_u6_U3 (.A( u1_u14_u6_n110 ) , .ZN( u1_u14_u6_n166 ) );
  NOR2_X1 u1_u14_u6_U30 (.A1( u1_u14_u6_n162 ) , .A2( u1_u14_u6_n165 ) , .ZN( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U31 (.A1( u1_u14_u6_n144 ) , .ZN( u1_u14_u6_n151 ) , .A2( u1_u14_u6_n158 ) );
  NAND2_X1 u1_u14_u6_U32 (.ZN( u1_u14_u6_n132 ) , .A1( u1_u14_u6_n91 ) , .A2( u1_u14_u6_n97 ) );
  AOI22_X1 u1_u14_u6_U33 (.B2( u1_u14_u6_n110 ) , .B1( u1_u14_u6_n111 ) , .A1( u1_u14_u6_n112 ) , .ZN( u1_u14_u6_n115 ) , .A2( u1_u14_u6_n161 ) );
  NAND4_X1 u1_u14_u6_U34 (.A3( u1_u14_u6_n109 ) , .ZN( u1_u14_u6_n112 ) , .A4( u1_u14_u6_n132 ) , .A2( u1_u14_u6_n147 ) , .A1( u1_u14_u6_n166 ) );
  NOR2_X1 u1_u14_u6_U35 (.ZN( u1_u14_u6_n109 ) , .A1( u1_u14_u6_n170 ) , .A2( u1_u14_u6_n173 ) );
  NOR2_X1 u1_u14_u6_U36 (.A2( u1_u14_u6_n126 ) , .ZN( u1_u14_u6_n155 ) , .A1( u1_u14_u6_n160 ) );
  NAND2_X1 u1_u14_u6_U37 (.ZN( u1_u14_u6_n146 ) , .A2( u1_u14_u6_n94 ) , .A1( u1_u14_u6_n99 ) );
  AOI21_X1 u1_u14_u6_U38 (.A( u1_u14_u6_n144 ) , .B2( u1_u14_u6_n145 ) , .B1( u1_u14_u6_n146 ) , .ZN( u1_u14_u6_n150 ) );
  AOI211_X1 u1_u14_u6_U39 (.B( u1_u14_u6_n134 ) , .A( u1_u14_u6_n135 ) , .C1( u1_u14_u6_n136 ) , .ZN( u1_u14_u6_n137 ) , .C2( u1_u14_u6_n151 ) );
  INV_X1 u1_u14_u6_U4 (.A( u1_u14_u6_n142 ) , .ZN( u1_u14_u6_n174 ) );
  AOI21_X1 u1_u14_u6_U40 (.B2( u1_u14_u6_n132 ) , .B1( u1_u14_u6_n133 ) , .ZN( u1_u14_u6_n134 ) , .A( u1_u14_u6_n158 ) );
  NAND4_X1 u1_u14_u6_U41 (.A4( u1_u14_u6_n127 ) , .A3( u1_u14_u6_n128 ) , .A2( u1_u14_u6_n129 ) , .A1( u1_u14_u6_n130 ) , .ZN( u1_u14_u6_n136 ) );
  AOI21_X1 u1_u14_u6_U42 (.B1( u1_u14_u6_n131 ) , .ZN( u1_u14_u6_n135 ) , .A( u1_u14_u6_n144 ) , .B2( u1_u14_u6_n146 ) );
  INV_X1 u1_u14_u6_U43 (.A( u1_u14_u6_n111 ) , .ZN( u1_u14_u6_n158 ) );
  NAND2_X1 u1_u14_u6_U44 (.ZN( u1_u14_u6_n127 ) , .A1( u1_u14_u6_n91 ) , .A2( u1_u14_u6_n92 ) );
  NAND2_X1 u1_u14_u6_U45 (.ZN( u1_u14_u6_n129 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n96 ) );
  INV_X1 u1_u14_u6_U46 (.A( u1_u14_u6_n144 ) , .ZN( u1_u14_u6_n159 ) );
  NAND2_X1 u1_u14_u6_U47 (.ZN( u1_u14_u6_n145 ) , .A2( u1_u14_u6_n97 ) , .A1( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U48 (.ZN( u1_u14_u6_n148 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n94 ) );
  NAND2_X1 u1_u14_u6_U49 (.ZN( u1_u14_u6_n108 ) , .A2( u1_u14_u6_n139 ) , .A1( u1_u14_u6_n144 ) );
  NAND2_X1 u1_u14_u6_U5 (.A2( u1_u14_u6_n143 ) , .ZN( u1_u14_u6_n152 ) , .A1( u1_u14_u6_n166 ) );
  NAND2_X1 u1_u14_u6_U50 (.ZN( u1_u14_u6_n121 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n97 ) );
  NAND2_X1 u1_u14_u6_U51 (.ZN( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n95 ) );
  AND2_X1 u1_u14_u6_U52 (.ZN( u1_u14_u6_n118 ) , .A2( u1_u14_u6_n91 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U53 (.ZN( u1_u14_u6_n147 ) , .A2( u1_u14_u6_n98 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U54 (.ZN( u1_u14_u6_n128 ) , .A1( u1_u14_u6_n94 ) , .A2( u1_u14_u6_n96 ) );
  NAND2_X1 u1_u14_u6_U55 (.ZN( u1_u14_u6_n119 ) , .A2( u1_u14_u6_n95 ) , .A1( u1_u14_u6_n99 ) );
  NAND2_X1 u1_u14_u6_U56 (.ZN( u1_u14_u6_n123 ) , .A2( u1_u14_u6_n91 ) , .A1( u1_u14_u6_n96 ) );
  NAND2_X1 u1_u14_u6_U57 (.ZN( u1_u14_u6_n100 ) , .A2( u1_u14_u6_n92 ) , .A1( u1_u14_u6_n98 ) );
  NAND2_X1 u1_u14_u6_U58 (.ZN( u1_u14_u6_n122 ) , .A1( u1_u14_u6_n94 ) , .A2( u1_u14_u6_n97 ) );
  INV_X1 u1_u14_u6_U59 (.A( u1_u14_u6_n139 ) , .ZN( u1_u14_u6_n160 ) );
  AOI22_X1 u1_u14_u6_U6 (.B2( u1_u14_u6_n101 ) , .A1( u1_u14_u6_n102 ) , .ZN( u1_u14_u6_n103 ) , .B1( u1_u14_u6_n160 ) , .A2( u1_u14_u6_n161 ) );
  NAND2_X1 u1_u14_u6_U60 (.ZN( u1_u14_u6_n113 ) , .A1( u1_u14_u6_n96 ) , .A2( u1_u14_u6_n98 ) );
  NOR2_X1 u1_u14_u6_U61 (.A2( u1_u14_X_40 ) , .A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n126 ) );
  NOR2_X1 u1_u14_u6_U62 (.A2( u1_u14_X_39 ) , .A1( u1_u14_X_42 ) , .ZN( u1_u14_u6_n92 ) );
  NOR2_X1 u1_u14_u6_U63 (.A2( u1_u14_X_39 ) , .A1( u1_u14_u6_n156 ) , .ZN( u1_u14_u6_n97 ) );
  NOR2_X1 u1_u14_u6_U64 (.A2( u1_u14_X_38 ) , .A1( u1_u14_u6_n165 ) , .ZN( u1_u14_u6_n95 ) );
  NOR2_X1 u1_u14_u6_U65 (.A2( u1_u14_X_41 ) , .ZN( u1_u14_u6_n111 ) , .A1( u1_u14_u6_n157 ) );
  NOR2_X1 u1_u14_u6_U66 (.A2( u1_u14_X_37 ) , .A1( u1_u14_u6_n162 ) , .ZN( u1_u14_u6_n94 ) );
  NOR2_X1 u1_u14_u6_U67 (.A2( u1_u14_X_37 ) , .A1( u1_u14_X_38 ) , .ZN( u1_u14_u6_n91 ) );
  NAND2_X1 u1_u14_u6_U68 (.A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n144 ) , .A2( u1_u14_u6_n157 ) );
  NAND2_X1 u1_u14_u6_U69 (.A2( u1_u14_X_40 ) , .A1( u1_u14_X_41 ) , .ZN( u1_u14_u6_n139 ) );
  NOR2_X1 u1_u14_u6_U7 (.A1( u1_u14_u6_n118 ) , .ZN( u1_u14_u6_n143 ) , .A2( u1_u14_u6_n168 ) );
  AND2_X1 u1_u14_u6_U70 (.A1( u1_u14_X_39 ) , .A2( u1_u14_u6_n156 ) , .ZN( u1_u14_u6_n96 ) );
  AND2_X1 u1_u14_u6_U71 (.A1( u1_u14_X_39 ) , .A2( u1_u14_X_42 ) , .ZN( u1_u14_u6_n99 ) );
  INV_X1 u1_u14_u6_U72 (.A( u1_u14_X_40 ) , .ZN( u1_u14_u6_n157 ) );
  INV_X1 u1_u14_u6_U73 (.A( u1_u14_X_37 ) , .ZN( u1_u14_u6_n165 ) );
  INV_X1 u1_u14_u6_U74 (.A( u1_u14_X_38 ) , .ZN( u1_u14_u6_n162 ) );
  INV_X1 u1_u14_u6_U75 (.A( u1_u14_X_42 ) , .ZN( u1_u14_u6_n156 ) );
  NAND4_X1 u1_u14_u6_U76 (.ZN( u1_out14_32 ) , .A4( u1_u14_u6_n103 ) , .A3( u1_u14_u6_n104 ) , .A2( u1_u14_u6_n105 ) , .A1( u1_u14_u6_n106 ) );
  AOI22_X1 u1_u14_u6_U77 (.ZN( u1_u14_u6_n105 ) , .A2( u1_u14_u6_n108 ) , .A1( u1_u14_u6_n118 ) , .B2( u1_u14_u6_n126 ) , .B1( u1_u14_u6_n171 ) );
  AOI22_X1 u1_u14_u6_U78 (.ZN( u1_u14_u6_n104 ) , .A1( u1_u14_u6_n111 ) , .B1( u1_u14_u6_n124 ) , .B2( u1_u14_u6_n151 ) , .A2( u1_u14_u6_n93 ) );
  NAND4_X1 u1_u14_u6_U79 (.ZN( u1_out14_12 ) , .A4( u1_u14_u6_n114 ) , .A3( u1_u14_u6_n115 ) , .A2( u1_u14_u6_n116 ) , .A1( u1_u14_u6_n117 ) );
  INV_X1 u1_u14_u6_U8 (.ZN( u1_u14_u6_n172 ) , .A( u1_u14_u6_n88 ) );
  OAI22_X1 u1_u14_u6_U80 (.B2( u1_u14_u6_n111 ) , .ZN( u1_u14_u6_n116 ) , .B1( u1_u14_u6_n126 ) , .A2( u1_u14_u6_n164 ) , .A1( u1_u14_u6_n167 ) );
  OAI21_X1 u1_u14_u6_U81 (.A( u1_u14_u6_n108 ) , .ZN( u1_u14_u6_n117 ) , .B2( u1_u14_u6_n141 ) , .B1( u1_u14_u6_n163 ) );
  OAI211_X1 u1_u14_u6_U82 (.ZN( u1_out14_22 ) , .B( u1_u14_u6_n137 ) , .A( u1_u14_u6_n138 ) , .C2( u1_u14_u6_n139 ) , .C1( u1_u14_u6_n140 ) );
  AOI22_X1 u1_u14_u6_U83 (.B1( u1_u14_u6_n124 ) , .A2( u1_u14_u6_n125 ) , .A1( u1_u14_u6_n126 ) , .ZN( u1_u14_u6_n138 ) , .B2( u1_u14_u6_n161 ) );
  AND4_X1 u1_u14_u6_U84 (.A3( u1_u14_u6_n119 ) , .A1( u1_u14_u6_n120 ) , .A4( u1_u14_u6_n129 ) , .ZN( u1_u14_u6_n140 ) , .A2( u1_u14_u6_n143 ) );
  OAI211_X1 u1_u14_u6_U85 (.ZN( u1_out14_7 ) , .B( u1_u14_u6_n153 ) , .C2( u1_u14_u6_n154 ) , .C1( u1_u14_u6_n155 ) , .A( u1_u14_u6_n174 ) );
  NOR3_X1 u1_u14_u6_U86 (.A1( u1_u14_u6_n141 ) , .ZN( u1_u14_u6_n154 ) , .A3( u1_u14_u6_n164 ) , .A2( u1_u14_u6_n171 ) );
  AOI211_X1 u1_u14_u6_U87 (.B( u1_u14_u6_n149 ) , .A( u1_u14_u6_n150 ) , .C2( u1_u14_u6_n151 ) , .C1( u1_u14_u6_n152 ) , .ZN( u1_u14_u6_n153 ) );
  NAND3_X1 u1_u14_u6_U88 (.A2( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n125 ) , .A1( u1_u14_u6_n130 ) , .A3( u1_u14_u6_n131 ) );
  NAND3_X1 u1_u14_u6_U89 (.A3( u1_u14_u6_n133 ) , .ZN( u1_u14_u6_n141 ) , .A1( u1_u14_u6_n145 ) , .A2( u1_u14_u6_n148 ) );
  OAI21_X1 u1_u14_u6_U9 (.A( u1_u14_u6_n159 ) , .B1( u1_u14_u6_n169 ) , .B2( u1_u14_u6_n173 ) , .ZN( u1_u14_u6_n90 ) );
  NAND3_X1 u1_u14_u6_U90 (.ZN( u1_u14_u6_n101 ) , .A3( u1_u14_u6_n107 ) , .A2( u1_u14_u6_n121 ) , .A1( u1_u14_u6_n127 ) );
  NAND3_X1 u1_u14_u6_U91 (.ZN( u1_u14_u6_n102 ) , .A3( u1_u14_u6_n130 ) , .A2( u1_u14_u6_n145 ) , .A1( u1_u14_u6_n166 ) );
  NAND3_X1 u1_u14_u6_U92 (.A3( u1_u14_u6_n113 ) , .A1( u1_u14_u6_n119 ) , .A2( u1_u14_u6_n123 ) , .ZN( u1_u14_u6_n93 ) );
  NAND3_X1 u1_u14_u6_U93 (.ZN( u1_u14_u6_n142 ) , .A2( u1_u14_u6_n172 ) , .A3( u1_u14_u6_n89 ) , .A1( u1_u14_u6_n90 ) );
  OAI21_X1 u1_u14_u7_U10 (.A( u1_u14_u7_n161 ) , .B1( u1_u14_u7_n168 ) , .B2( u1_u14_u7_n173 ) , .ZN( u1_u14_u7_n91 ) );
  AOI211_X1 u1_u14_u7_U11 (.A( u1_u14_u7_n117 ) , .ZN( u1_u14_u7_n118 ) , .C2( u1_u14_u7_n126 ) , .C1( u1_u14_u7_n177 ) , .B( u1_u14_u7_n180 ) );
  OAI22_X1 u1_u14_u7_U12 (.B1( u1_u14_u7_n115 ) , .ZN( u1_u14_u7_n117 ) , .A2( u1_u14_u7_n133 ) , .A1( u1_u14_u7_n137 ) , .B2( u1_u14_u7_n162 ) );
  INV_X1 u1_u14_u7_U13 (.A( u1_u14_u7_n116 ) , .ZN( u1_u14_u7_n180 ) );
  NOR3_X1 u1_u14_u7_U14 (.ZN( u1_u14_u7_n115 ) , .A3( u1_u14_u7_n145 ) , .A2( u1_u14_u7_n168 ) , .A1( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U15 (.A( u1_u14_u7_n133 ) , .ZN( u1_u14_u7_n176 ) );
  NOR3_X1 u1_u14_u7_U16 (.A2( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n135 ) , .ZN( u1_u14_u7_n136 ) , .A3( u1_u14_u7_n171 ) );
  NOR2_X1 u1_u14_u7_U17 (.A1( u1_u14_u7_n130 ) , .A2( u1_u14_u7_n134 ) , .ZN( u1_u14_u7_n153 ) );
  AOI21_X1 u1_u14_u7_U18 (.ZN( u1_u14_u7_n104 ) , .B2( u1_u14_u7_n112 ) , .B1( u1_u14_u7_n127 ) , .A( u1_u14_u7_n164 ) );
  AOI21_X1 u1_u14_u7_U19 (.ZN( u1_u14_u7_n106 ) , .B1( u1_u14_u7_n133 ) , .B2( u1_u14_u7_n146 ) , .A( u1_u14_u7_n162 ) );
  AOI21_X1 u1_u14_u7_U20 (.A( u1_u14_u7_n101 ) , .ZN( u1_u14_u7_n107 ) , .B2( u1_u14_u7_n128 ) , .B1( u1_u14_u7_n175 ) );
  INV_X1 u1_u14_u7_U21 (.A( u1_u14_u7_n101 ) , .ZN( u1_u14_u7_n165 ) );
  NOR2_X1 u1_u14_u7_U22 (.ZN( u1_u14_u7_n111 ) , .A2( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U23 (.A( u1_u14_u7_n138 ) , .ZN( u1_u14_u7_n171 ) );
  INV_X1 u1_u14_u7_U24 (.A( u1_u14_u7_n131 ) , .ZN( u1_u14_u7_n177 ) );
  INV_X1 u1_u14_u7_U25 (.A( u1_u14_u7_n110 ) , .ZN( u1_u14_u7_n174 ) );
  NAND2_X1 u1_u14_u7_U26 (.A1( u1_u14_u7_n129 ) , .A2( u1_u14_u7_n132 ) , .ZN( u1_u14_u7_n149 ) );
  NAND2_X1 u1_u14_u7_U27 (.A1( u1_u14_u7_n113 ) , .A2( u1_u14_u7_n124 ) , .ZN( u1_u14_u7_n130 ) );
  INV_X1 u1_u14_u7_U28 (.A( u1_u14_u7_n112 ) , .ZN( u1_u14_u7_n173 ) );
  INV_X1 u1_u14_u7_U29 (.A( u1_u14_u7_n128 ) , .ZN( u1_u14_u7_n168 ) );
  OAI21_X1 u1_u14_u7_U3 (.ZN( u1_u14_u7_n159 ) , .A( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n171 ) , .B1( u1_u14_u7_n174 ) );
  INV_X1 u1_u14_u7_U30 (.A( u1_u14_u7_n148 ) , .ZN( u1_u14_u7_n169 ) );
  INV_X1 u1_u14_u7_U31 (.A( u1_u14_u7_n127 ) , .ZN( u1_u14_u7_n179 ) );
  NOR2_X1 u1_u14_u7_U32 (.ZN( u1_u14_u7_n101 ) , .A2( u1_u14_u7_n150 ) , .A1( u1_u14_u7_n156 ) );
  AOI211_X1 u1_u14_u7_U33 (.B( u1_u14_u7_n139 ) , .A( u1_u14_u7_n140 ) , .C2( u1_u14_u7_n141 ) , .ZN( u1_u14_u7_n142 ) , .C1( u1_u14_u7_n156 ) );
  NAND4_X1 u1_u14_u7_U34 (.A3( u1_u14_u7_n127 ) , .A2( u1_u14_u7_n128 ) , .A1( u1_u14_u7_n129 ) , .ZN( u1_u14_u7_n141 ) , .A4( u1_u14_u7_n147 ) );
  AOI21_X1 u1_u14_u7_U35 (.A( u1_u14_u7_n137 ) , .B1( u1_u14_u7_n138 ) , .ZN( u1_u14_u7_n139 ) , .B2( u1_u14_u7_n146 ) );
  OAI22_X1 u1_u14_u7_U36 (.B1( u1_u14_u7_n136 ) , .ZN( u1_u14_u7_n140 ) , .A1( u1_u14_u7_n153 ) , .B2( u1_u14_u7_n162 ) , .A2( u1_u14_u7_n164 ) );
  INV_X1 u1_u14_u7_U37 (.A( u1_u14_u7_n125 ) , .ZN( u1_u14_u7_n161 ) );
  AOI21_X1 u1_u14_u7_U38 (.ZN( u1_u14_u7_n123 ) , .B1( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n177 ) , .A( u1_u14_u7_n97 ) );
  AOI21_X1 u1_u14_u7_U39 (.B2( u1_u14_u7_n113 ) , .B1( u1_u14_u7_n124 ) , .A( u1_u14_u7_n125 ) , .ZN( u1_u14_u7_n97 ) );
  INV_X1 u1_u14_u7_U4 (.A( u1_u14_u7_n149 ) , .ZN( u1_u14_u7_n175 ) );
  INV_X1 u1_u14_u7_U40 (.A( u1_u14_u7_n152 ) , .ZN( u1_u14_u7_n162 ) );
  AOI22_X1 u1_u14_u7_U41 (.A2( u1_u14_u7_n114 ) , .ZN( u1_u14_u7_n119 ) , .B1( u1_u14_u7_n130 ) , .A1( u1_u14_u7_n156 ) , .B2( u1_u14_u7_n165 ) );
  NAND2_X1 u1_u14_u7_U42 (.A2( u1_u14_u7_n112 ) , .ZN( u1_u14_u7_n114 ) , .A1( u1_u14_u7_n175 ) );
  NOR2_X1 u1_u14_u7_U43 (.ZN( u1_u14_u7_n137 ) , .A1( u1_u14_u7_n150 ) , .A2( u1_u14_u7_n161 ) );
  AND2_X1 u1_u14_u7_U44 (.ZN( u1_u14_u7_n145 ) , .A2( u1_u14_u7_n98 ) , .A1( u1_u14_u7_n99 ) );
  AOI21_X1 u1_u14_u7_U45 (.ZN( u1_u14_u7_n105 ) , .B2( u1_u14_u7_n110 ) , .A( u1_u14_u7_n125 ) , .B1( u1_u14_u7_n147 ) );
  NAND2_X1 u1_u14_u7_U46 (.ZN( u1_u14_u7_n146 ) , .A1( u1_u14_u7_n95 ) , .A2( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U47 (.A2( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n147 ) , .A1( u1_u14_u7_n93 ) );
  NAND2_X1 u1_u14_u7_U48 (.A1( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n127 ) , .A2( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U49 (.A2( u1_u14_u7_n102 ) , .A1( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n133 ) );
  INV_X1 u1_u14_u7_U5 (.A( u1_u14_u7_n154 ) , .ZN( u1_u14_u7_n178 ) );
  OR2_X1 u1_u14_u7_U50 (.ZN( u1_u14_u7_n126 ) , .A2( u1_u14_u7_n152 ) , .A1( u1_u14_u7_n156 ) );
  NAND2_X1 u1_u14_u7_U51 (.ZN( u1_u14_u7_n112 ) , .A2( u1_u14_u7_n96 ) , .A1( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U52 (.A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n128 ) , .A1( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U53 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n113 ) , .A2( u1_u14_u7_n93 ) );
  NAND2_X1 u1_u14_u7_U54 (.ZN( u1_u14_u7_n110 ) , .A1( u1_u14_u7_n95 ) , .A2( u1_u14_u7_n96 ) );
  INV_X1 u1_u14_u7_U55 (.A( u1_u14_u7_n150 ) , .ZN( u1_u14_u7_n164 ) );
  AND2_X1 u1_u14_u7_U56 (.ZN( u1_u14_u7_n134 ) , .A1( u1_u14_u7_n93 ) , .A2( u1_u14_u7_n98 ) );
  NAND2_X1 u1_u14_u7_U57 (.A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n124 ) , .A1( u1_u14_u7_n96 ) );
  NAND2_X1 u1_u14_u7_U58 (.A1( u1_u14_u7_n100 ) , .A2( u1_u14_u7_n102 ) , .ZN( u1_u14_u7_n129 ) );
  NAND2_X1 u1_u14_u7_U59 (.A2( u1_u14_u7_n103 ) , .ZN( u1_u14_u7_n131 ) , .A1( u1_u14_u7_n95 ) );
  AOI211_X1 u1_u14_u7_U6 (.ZN( u1_u14_u7_n116 ) , .A( u1_u14_u7_n155 ) , .C1( u1_u14_u7_n161 ) , .C2( u1_u14_u7_n171 ) , .B( u1_u14_u7_n94 ) );
  NAND2_X1 u1_u14_u7_U60 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n138 ) , .A2( u1_u14_u7_n99 ) );
  NAND2_X1 u1_u14_u7_U61 (.ZN( u1_u14_u7_n132 ) , .A1( u1_u14_u7_n93 ) , .A2( u1_u14_u7_n96 ) );
  NAND2_X1 u1_u14_u7_U62 (.A1( u1_u14_u7_n100 ) , .ZN( u1_u14_u7_n148 ) , .A2( u1_u14_u7_n95 ) );
  AOI211_X1 u1_u14_u7_U63 (.B( u1_u14_u7_n154 ) , .A( u1_u14_u7_n155 ) , .C1( u1_u14_u7_n156 ) , .ZN( u1_u14_u7_n157 ) , .C2( u1_u14_u7_n172 ) );
  INV_X1 u1_u14_u7_U64 (.A( u1_u14_u7_n153 ) , .ZN( u1_u14_u7_n172 ) );
  NOR2_X1 u1_u14_u7_U65 (.A2( u1_u14_X_47 ) , .ZN( u1_u14_u7_n150 ) , .A1( u1_u14_u7_n163 ) );
  NOR2_X1 u1_u14_u7_U66 (.A2( u1_u14_X_43 ) , .A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n103 ) );
  NOR2_X1 u1_u14_u7_U67 (.A2( u1_u14_X_48 ) , .A1( u1_u14_u7_n166 ) , .ZN( u1_u14_u7_n95 ) );
  NOR2_X1 u1_u14_u7_U68 (.A2( u1_u14_X_45 ) , .A1( u1_u14_X_48 ) , .ZN( u1_u14_u7_n99 ) );
  NOR2_X1 u1_u14_u7_U69 (.A2( u1_u14_X_44 ) , .A1( u1_u14_u7_n167 ) , .ZN( u1_u14_u7_n98 ) );
  OAI222_X1 u1_u14_u7_U7 (.C2( u1_u14_u7_n101 ) , .B2( u1_u14_u7_n111 ) , .A1( u1_u14_u7_n113 ) , .C1( u1_u14_u7_n146 ) , .A2( u1_u14_u7_n162 ) , .B1( u1_u14_u7_n164 ) , .ZN( u1_u14_u7_n94 ) );
  NOR2_X1 u1_u14_u7_U70 (.A2( u1_u14_X_46 ) , .A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n152 ) );
  NAND2_X1 u1_u14_u7_U71 (.A2( u1_u14_X_46 ) , .A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n125 ) );
  AND2_X1 u1_u14_u7_U72 (.A1( u1_u14_X_47 ) , .ZN( u1_u14_u7_n156 ) , .A2( u1_u14_u7_n163 ) );
  AND2_X1 u1_u14_u7_U73 (.A2( u1_u14_X_45 ) , .A1( u1_u14_X_48 ) , .ZN( u1_u14_u7_n102 ) );
  AND2_X1 u1_u14_u7_U74 (.A2( u1_u14_X_43 ) , .A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n96 ) );
  AND2_X1 u1_u14_u7_U75 (.A1( u1_u14_X_44 ) , .ZN( u1_u14_u7_n100 ) , .A2( u1_u14_u7_n167 ) );
  AND2_X1 u1_u14_u7_U76 (.A1( u1_u14_X_48 ) , .A2( u1_u14_u7_n166 ) , .ZN( u1_u14_u7_n93 ) );
  INV_X1 u1_u14_u7_U77 (.A( u1_u14_X_46 ) , .ZN( u1_u14_u7_n163 ) );
  INV_X1 u1_u14_u7_U78 (.A( u1_u14_X_43 ) , .ZN( u1_u14_u7_n167 ) );
  INV_X1 u1_u14_u7_U79 (.A( u1_u14_X_45 ) , .ZN( u1_u14_u7_n166 ) );
  OAI221_X1 u1_u14_u7_U8 (.C1( u1_u14_u7_n101 ) , .C2( u1_u14_u7_n147 ) , .ZN( u1_u14_u7_n155 ) , .B2( u1_u14_u7_n162 ) , .A( u1_u14_u7_n91 ) , .B1( u1_u14_u7_n92 ) );
  NAND4_X1 u1_u14_u7_U80 (.ZN( u1_out14_5 ) , .A4( u1_u14_u7_n108 ) , .A3( u1_u14_u7_n109 ) , .A1( u1_u14_u7_n116 ) , .A2( u1_u14_u7_n123 ) );
  AOI22_X1 u1_u14_u7_U81 (.ZN( u1_u14_u7_n109 ) , .A2( u1_u14_u7_n126 ) , .B2( u1_u14_u7_n145 ) , .B1( u1_u14_u7_n156 ) , .A1( u1_u14_u7_n171 ) );
  NOR4_X1 u1_u14_u7_U82 (.A4( u1_u14_u7_n104 ) , .A3( u1_u14_u7_n105 ) , .A2( u1_u14_u7_n106 ) , .A1( u1_u14_u7_n107 ) , .ZN( u1_u14_u7_n108 ) );
  NAND4_X1 u1_u14_u7_U83 (.ZN( u1_out14_27 ) , .A4( u1_u14_u7_n118 ) , .A3( u1_u14_u7_n119 ) , .A2( u1_u14_u7_n120 ) , .A1( u1_u14_u7_n121 ) );
  OAI21_X1 u1_u14_u7_U84 (.ZN( u1_u14_u7_n121 ) , .B2( u1_u14_u7_n145 ) , .A( u1_u14_u7_n150 ) , .B1( u1_u14_u7_n174 ) );
  OAI21_X1 u1_u14_u7_U85 (.ZN( u1_u14_u7_n120 ) , .A( u1_u14_u7_n161 ) , .B2( u1_u14_u7_n170 ) , .B1( u1_u14_u7_n179 ) );
  NAND4_X1 u1_u14_u7_U86 (.ZN( u1_out14_21 ) , .A4( u1_u14_u7_n157 ) , .A3( u1_u14_u7_n158 ) , .A2( u1_u14_u7_n159 ) , .A1( u1_u14_u7_n160 ) );
  OAI21_X1 u1_u14_u7_U87 (.B1( u1_u14_u7_n145 ) , .ZN( u1_u14_u7_n160 ) , .A( u1_u14_u7_n161 ) , .B2( u1_u14_u7_n177 ) );
  AOI22_X1 u1_u14_u7_U88 (.B2( u1_u14_u7_n149 ) , .B1( u1_u14_u7_n150 ) , .A2( u1_u14_u7_n151 ) , .A1( u1_u14_u7_n152 ) , .ZN( u1_u14_u7_n158 ) );
  NAND4_X1 u1_u14_u7_U89 (.ZN( u1_out14_15 ) , .A4( u1_u14_u7_n142 ) , .A3( u1_u14_u7_n143 ) , .A2( u1_u14_u7_n144 ) , .A1( u1_u14_u7_n178 ) );
  AND3_X1 u1_u14_u7_U9 (.A3( u1_u14_u7_n110 ) , .A2( u1_u14_u7_n127 ) , .A1( u1_u14_u7_n132 ) , .ZN( u1_u14_u7_n92 ) );
  OR2_X1 u1_u14_u7_U90 (.A2( u1_u14_u7_n125 ) , .A1( u1_u14_u7_n129 ) , .ZN( u1_u14_u7_n144 ) );
  AOI22_X1 u1_u14_u7_U91 (.A2( u1_u14_u7_n126 ) , .ZN( u1_u14_u7_n143 ) , .B2( u1_u14_u7_n165 ) , .B1( u1_u14_u7_n173 ) , .A1( u1_u14_u7_n174 ) );
  OAI211_X1 u1_u14_u7_U92 (.B( u1_u14_u7_n122 ) , .A( u1_u14_u7_n123 ) , .C2( u1_u14_u7_n124 ) , .ZN( u1_u14_u7_n154 ) , .C1( u1_u14_u7_n162 ) );
  AOI222_X1 u1_u14_u7_U93 (.ZN( u1_u14_u7_n122 ) , .C2( u1_u14_u7_n126 ) , .C1( u1_u14_u7_n145 ) , .B1( u1_u14_u7_n161 ) , .A2( u1_u14_u7_n165 ) , .B2( u1_u14_u7_n170 ) , .A1( u1_u14_u7_n176 ) );
  INV_X1 u1_u14_u7_U94 (.A( u1_u14_u7_n111 ) , .ZN( u1_u14_u7_n170 ) );
  NAND3_X1 u1_u14_u7_U95 (.A3( u1_u14_u7_n146 ) , .A2( u1_u14_u7_n147 ) , .A1( u1_u14_u7_n148 ) , .ZN( u1_u14_u7_n151 ) );
  NAND3_X1 u1_u14_u7_U96 (.A3( u1_u14_u7_n131 ) , .A2( u1_u14_u7_n132 ) , .A1( u1_u14_u7_n133 ) , .ZN( u1_u14_u7_n135 ) );
  XOR2_X1 u1_u15_U11 (.A( u1_FP_61 ) , .B( u1_K16_44 ) , .Z( u1_u15_X_44 ) );
  XOR2_X1 u1_u15_U12 (.A( u1_FP_60 ) , .B( u1_K16_43 ) , .Z( u1_u15_X_43 ) );
  XOR2_X1 u1_u15_U13 (.A( u1_FP_61 ) , .B( u1_K16_42 ) , .Z( u1_u15_X_42 ) );
  XOR2_X1 u1_u15_U14 (.A( u1_FP_60 ) , .B( u1_K16_41 ) , .Z( u1_u15_X_41 ) );
  XOR2_X1 u1_u15_U18 (.A( u1_FP_57 ) , .B( u1_K16_38 ) , .Z( u1_u15_X_38 ) );
  XOR2_X1 u1_u15_U19 (.A( u1_FP_56 ) , .B( u1_K16_37 ) , .Z( u1_u15_X_37 ) );
  XOR2_X1 u1_u15_U2 (.A( u1_FP_37 ) , .B( u1_K16_8 ) , .Z( u1_u15_X_8 ) );
  XOR2_X1 u1_u15_U20 (.A( u1_FP_57 ) , .B( u1_K16_36 ) , .Z( u1_u15_X_36 ) );
  XOR2_X1 u1_u15_U21 (.A( u1_FP_56 ) , .B( u1_K16_35 ) , .Z( u1_u15_X_35 ) );
  XOR2_X1 u1_u15_U24 (.A( u1_FP_53 ) , .B( u1_K16_32 ) , .Z( u1_u15_X_32 ) );
  XOR2_X1 u1_u15_U25 (.A( u1_FP_52 ) , .B( u1_K16_31 ) , .Z( u1_u15_X_31 ) );
  XOR2_X1 u1_u15_U26 (.A( u1_FP_53 ) , .B( u1_K16_30 ) , .Z( u1_u15_X_30 ) );
  XOR2_X1 u1_u15_U27 (.A( u1_FP_33 ) , .B( u1_K16_2 ) , .Z( u1_u15_X_2 ) );
  XOR2_X1 u1_u15_U28 (.A( u1_FP_52 ) , .B( u1_K16_29 ) , .Z( u1_u15_X_29 ) );
  XOR2_X1 u1_u15_U29 (.A( u1_FP_51 ) , .B( u1_K16_28 ) , .Z( u1_u15_X_28 ) );
  XOR2_X1 u1_u15_U3 (.A( u1_FP_36 ) , .B( u1_K16_7 ) , .Z( u1_u15_X_7 ) );
  XOR2_X1 u1_u15_U30 (.A( u1_FP_50 ) , .B( u1_K16_27 ) , .Z( u1_u15_X_27 ) );
  XOR2_X1 u1_u15_U31 (.A( u1_FP_49 ) , .B( u1_K16_26 ) , .Z( u1_u15_X_26 ) );
  XOR2_X1 u1_u15_U32 (.A( u1_FP_48 ) , .B( u1_K16_25 ) , .Z( u1_u15_X_25 ) );
  XOR2_X1 u1_u15_U33 (.A( u1_FP_49 ) , .B( u1_K16_24 ) , .Z( u1_u15_X_24 ) );
  XOR2_X1 u1_u15_U34 (.A( u1_FP_48 ) , .B( u1_K16_23 ) , .Z( u1_u15_X_23 ) );
  XOR2_X1 u1_u15_U35 (.A( u1_FP_47 ) , .B( u1_K16_22 ) , .Z( u1_u15_X_22 ) );
  XOR2_X1 u1_u15_U36 (.A( u1_FP_46 ) , .B( u1_K16_21 ) , .Z( u1_u15_X_21 ) );
  XOR2_X1 u1_u15_U37 (.A( u1_FP_45 ) , .B( u1_K16_20 ) , .Z( u1_u15_X_20 ) );
  XOR2_X1 u1_u15_U38 (.A( u1_FP_64 ) , .B( u1_K16_1 ) , .Z( u1_u15_X_1 ) );
  XOR2_X1 u1_u15_U39 (.A( u1_FP_44 ) , .B( u1_K16_19 ) , .Z( u1_u15_X_19 ) );
  XOR2_X1 u1_u15_U4 (.A( u1_FP_37 ) , .B( u1_K16_6 ) , .Z( u1_u15_X_6 ) );
  XOR2_X1 u1_u15_U40 (.A( u1_FP_45 ) , .B( u1_K16_18 ) , .Z( u1_u15_X_18 ) );
  XOR2_X1 u1_u15_U41 (.A( u1_FP_44 ) , .B( u1_K16_17 ) , .Z( u1_u15_X_17 ) );
  XOR2_X1 u1_u15_U44 (.A( u1_FP_41 ) , .B( u1_K16_14 ) , .Z( u1_u15_X_14 ) );
  XOR2_X1 u1_u15_U45 (.A( u1_FP_40 ) , .B( u1_K16_13 ) , .Z( u1_u15_X_13 ) );
  XOR2_X1 u1_u15_U46 (.A( u1_FP_41 ) , .B( u1_K16_12 ) , .Z( u1_u15_X_12 ) );
  XOR2_X1 u1_u15_U47 (.A( u1_FP_40 ) , .B( u1_K16_11 ) , .Z( u1_u15_X_11 ) );
  XOR2_X1 u1_u15_U5 (.A( u1_FP_36 ) , .B( u1_K16_5 ) , .Z( u1_u15_X_5 ) );
  XOR2_X1 u1_u15_U7 (.A( u1_FP_33 ) , .B( u1_K16_48 ) , .Z( u1_u15_X_48 ) );
  XOR2_X1 u1_u15_U8 (.A( u1_FP_64 ) , .B( u1_K16_47 ) , .Z( u1_u15_X_47 ) );
  OAI22_X1 u1_u15_u3_U10 (.B1( u1_u15_u3_n113 ) , .A2( u1_u15_u3_n135 ) , .A1( u1_u15_u3_n150 ) , .B2( u1_u15_u3_n164 ) , .ZN( u1_u15_u3_n98 ) );
  OAI211_X1 u1_u15_u3_U11 (.B( u1_u15_u3_n106 ) , .ZN( u1_u15_u3_n119 ) , .C2( u1_u15_u3_n128 ) , .C1( u1_u15_u3_n167 ) , .A( u1_u15_u3_n181 ) );
  AOI221_X1 u1_u15_u3_U12 (.C1( u1_u15_u3_n105 ) , .ZN( u1_u15_u3_n106 ) , .A( u1_u15_u3_n131 ) , .B2( u1_u15_u3_n132 ) , .C2( u1_u15_u3_n133 ) , .B1( u1_u15_u3_n169 ) );
  INV_X1 u1_u15_u3_U13 (.ZN( u1_u15_u3_n181 ) , .A( u1_u15_u3_n98 ) );
  NAND2_X1 u1_u15_u3_U14 (.ZN( u1_u15_u3_n105 ) , .A2( u1_u15_u3_n130 ) , .A1( u1_u15_u3_n155 ) );
  AOI22_X1 u1_u15_u3_U15 (.B1( u1_u15_u3_n115 ) , .A2( u1_u15_u3_n116 ) , .ZN( u1_u15_u3_n123 ) , .B2( u1_u15_u3_n133 ) , .A1( u1_u15_u3_n169 ) );
  NAND2_X1 u1_u15_u3_U16 (.ZN( u1_u15_u3_n116 ) , .A2( u1_u15_u3_n151 ) , .A1( u1_u15_u3_n182 ) );
  NOR2_X1 u1_u15_u3_U17 (.ZN( u1_u15_u3_n126 ) , .A2( u1_u15_u3_n150 ) , .A1( u1_u15_u3_n164 ) );
  AOI21_X1 u1_u15_u3_U18 (.ZN( u1_u15_u3_n112 ) , .B2( u1_u15_u3_n146 ) , .B1( u1_u15_u3_n155 ) , .A( u1_u15_u3_n167 ) );
  NAND2_X1 u1_u15_u3_U19 (.A1( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n142 ) , .A2( u1_u15_u3_n164 ) );
  NAND2_X1 u1_u15_u3_U20 (.ZN( u1_u15_u3_n132 ) , .A2( u1_u15_u3_n152 ) , .A1( u1_u15_u3_n156 ) );
  AND2_X1 u1_u15_u3_U21 (.A2( u1_u15_u3_n113 ) , .A1( u1_u15_u3_n114 ) , .ZN( u1_u15_u3_n151 ) );
  INV_X1 u1_u15_u3_U22 (.A( u1_u15_u3_n133 ) , .ZN( u1_u15_u3_n165 ) );
  INV_X1 u1_u15_u3_U23 (.A( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n170 ) );
  NAND2_X1 u1_u15_u3_U24 (.A1( u1_u15_u3_n107 ) , .A2( u1_u15_u3_n108 ) , .ZN( u1_u15_u3_n140 ) );
  NAND2_X1 u1_u15_u3_U25 (.ZN( u1_u15_u3_n117 ) , .A1( u1_u15_u3_n124 ) , .A2( u1_u15_u3_n148 ) );
  NAND2_X1 u1_u15_u3_U26 (.ZN( u1_u15_u3_n143 ) , .A1( u1_u15_u3_n165 ) , .A2( u1_u15_u3_n167 ) );
  INV_X1 u1_u15_u3_U27 (.A( u1_u15_u3_n130 ) , .ZN( u1_u15_u3_n177 ) );
  INV_X1 u1_u15_u3_U28 (.A( u1_u15_u3_n128 ) , .ZN( u1_u15_u3_n176 ) );
  INV_X1 u1_u15_u3_U29 (.A( u1_u15_u3_n155 ) , .ZN( u1_u15_u3_n174 ) );
  INV_X1 u1_u15_u3_U3 (.A( u1_u15_u3_n129 ) , .ZN( u1_u15_u3_n183 ) );
  INV_X1 u1_u15_u3_U30 (.A( u1_u15_u3_n139 ) , .ZN( u1_u15_u3_n185 ) );
  NOR2_X1 u1_u15_u3_U31 (.ZN( u1_u15_u3_n135 ) , .A2( u1_u15_u3_n141 ) , .A1( u1_u15_u3_n169 ) );
  OAI222_X1 u1_u15_u3_U32 (.C2( u1_u15_u3_n107 ) , .A2( u1_u15_u3_n108 ) , .B1( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n138 ) , .B2( u1_u15_u3_n146 ) , .C1( u1_u15_u3_n154 ) , .A1( u1_u15_u3_n164 ) );
  NOR4_X1 u1_u15_u3_U33 (.A4( u1_u15_u3_n157 ) , .A3( u1_u15_u3_n158 ) , .A2( u1_u15_u3_n159 ) , .A1( u1_u15_u3_n160 ) , .ZN( u1_u15_u3_n161 ) );
  AOI21_X1 u1_u15_u3_U34 (.B2( u1_u15_u3_n152 ) , .B1( u1_u15_u3_n153 ) , .ZN( u1_u15_u3_n158 ) , .A( u1_u15_u3_n164 ) );
  AOI21_X1 u1_u15_u3_U35 (.A( u1_u15_u3_n154 ) , .B2( u1_u15_u3_n155 ) , .B1( u1_u15_u3_n156 ) , .ZN( u1_u15_u3_n157 ) );
  AOI21_X1 u1_u15_u3_U36 (.A( u1_u15_u3_n149 ) , .B2( u1_u15_u3_n150 ) , .B1( u1_u15_u3_n151 ) , .ZN( u1_u15_u3_n159 ) );
  AOI211_X1 u1_u15_u3_U37 (.ZN( u1_u15_u3_n109 ) , .A( u1_u15_u3_n119 ) , .C2( u1_u15_u3_n129 ) , .B( u1_u15_u3_n138 ) , .C1( u1_u15_u3_n141 ) );
  AOI211_X1 u1_u15_u3_U38 (.B( u1_u15_u3_n119 ) , .A( u1_u15_u3_n120 ) , .C2( u1_u15_u3_n121 ) , .ZN( u1_u15_u3_n122 ) , .C1( u1_u15_u3_n179 ) );
  INV_X1 u1_u15_u3_U39 (.A( u1_u15_u3_n156 ) , .ZN( u1_u15_u3_n179 ) );
  INV_X1 u1_u15_u3_U4 (.A( u1_u15_u3_n140 ) , .ZN( u1_u15_u3_n182 ) );
  OAI22_X1 u1_u15_u3_U40 (.B1( u1_u15_u3_n118 ) , .ZN( u1_u15_u3_n120 ) , .A1( u1_u15_u3_n135 ) , .B2( u1_u15_u3_n154 ) , .A2( u1_u15_u3_n178 ) );
  AND3_X1 u1_u15_u3_U41 (.ZN( u1_u15_u3_n118 ) , .A2( u1_u15_u3_n124 ) , .A1( u1_u15_u3_n144 ) , .A3( u1_u15_u3_n152 ) );
  INV_X1 u1_u15_u3_U42 (.A( u1_u15_u3_n121 ) , .ZN( u1_u15_u3_n164 ) );
  NAND2_X1 u1_u15_u3_U43 (.ZN( u1_u15_u3_n133 ) , .A1( u1_u15_u3_n154 ) , .A2( u1_u15_u3_n164 ) );
  OAI211_X1 u1_u15_u3_U44 (.B( u1_u15_u3_n127 ) , .ZN( u1_u15_u3_n139 ) , .C1( u1_u15_u3_n150 ) , .C2( u1_u15_u3_n154 ) , .A( u1_u15_u3_n184 ) );
  INV_X1 u1_u15_u3_U45 (.A( u1_u15_u3_n125 ) , .ZN( u1_u15_u3_n184 ) );
  AOI221_X1 u1_u15_u3_U46 (.A( u1_u15_u3_n126 ) , .ZN( u1_u15_u3_n127 ) , .C2( u1_u15_u3_n132 ) , .C1( u1_u15_u3_n169 ) , .B2( u1_u15_u3_n170 ) , .B1( u1_u15_u3_n174 ) );
  OAI22_X1 u1_u15_u3_U47 (.A1( u1_u15_u3_n124 ) , .ZN( u1_u15_u3_n125 ) , .B2( u1_u15_u3_n145 ) , .A2( u1_u15_u3_n165 ) , .B1( u1_u15_u3_n167 ) );
  NOR2_X1 u1_u15_u3_U48 (.A1( u1_u15_u3_n113 ) , .ZN( u1_u15_u3_n131 ) , .A2( u1_u15_u3_n154 ) );
  NAND2_X1 u1_u15_u3_U49 (.A1( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n150 ) , .A2( u1_u15_u3_n99 ) );
  INV_X1 u1_u15_u3_U5 (.A( u1_u15_u3_n117 ) , .ZN( u1_u15_u3_n178 ) );
  NAND2_X1 u1_u15_u3_U50 (.A2( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n155 ) , .A1( u1_u15_u3_n97 ) );
  INV_X1 u1_u15_u3_U51 (.A( u1_u15_u3_n141 ) , .ZN( u1_u15_u3_n167 ) );
  AOI21_X1 u1_u15_u3_U52 (.B2( u1_u15_u3_n114 ) , .B1( u1_u15_u3_n146 ) , .A( u1_u15_u3_n154 ) , .ZN( u1_u15_u3_n94 ) );
  AOI21_X1 u1_u15_u3_U53 (.ZN( u1_u15_u3_n110 ) , .B2( u1_u15_u3_n142 ) , .B1( u1_u15_u3_n186 ) , .A( u1_u15_u3_n95 ) );
  INV_X1 u1_u15_u3_U54 (.A( u1_u15_u3_n145 ) , .ZN( u1_u15_u3_n186 ) );
  AOI21_X1 u1_u15_u3_U55 (.B1( u1_u15_u3_n124 ) , .A( u1_u15_u3_n149 ) , .B2( u1_u15_u3_n155 ) , .ZN( u1_u15_u3_n95 ) );
  INV_X1 u1_u15_u3_U56 (.A( u1_u15_u3_n149 ) , .ZN( u1_u15_u3_n169 ) );
  NAND2_X1 u1_u15_u3_U57 (.ZN( u1_u15_u3_n124 ) , .A1( u1_u15_u3_n96 ) , .A2( u1_u15_u3_n97 ) );
  NAND2_X1 u1_u15_u3_U58 (.A2( u1_u15_u3_n100 ) , .ZN( u1_u15_u3_n146 ) , .A1( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U59 (.A1( u1_u15_u3_n101 ) , .ZN( u1_u15_u3_n145 ) , .A2( u1_u15_u3_n99 ) );
  AOI221_X1 u1_u15_u3_U6 (.A( u1_u15_u3_n131 ) , .C2( u1_u15_u3_n132 ) , .C1( u1_u15_u3_n133 ) , .ZN( u1_u15_u3_n134 ) , .B1( u1_u15_u3_n143 ) , .B2( u1_u15_u3_n177 ) );
  NAND2_X1 u1_u15_u3_U60 (.A1( u1_u15_u3_n100 ) , .ZN( u1_u15_u3_n156 ) , .A2( u1_u15_u3_n99 ) );
  NAND2_X1 u1_u15_u3_U61 (.A2( u1_u15_u3_n101 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n148 ) );
  NAND2_X1 u1_u15_u3_U62 (.A1( u1_u15_u3_n100 ) , .A2( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n128 ) );
  NAND2_X1 u1_u15_u3_U63 (.A2( u1_u15_u3_n101 ) , .A1( u1_u15_u3_n102 ) , .ZN( u1_u15_u3_n152 ) );
  NAND2_X1 u1_u15_u3_U64 (.A2( u1_u15_u3_n101 ) , .ZN( u1_u15_u3_n114 ) , .A1( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U65 (.ZN( u1_u15_u3_n107 ) , .A1( u1_u15_u3_n97 ) , .A2( u1_u15_u3_n99 ) );
  NAND2_X1 u1_u15_u3_U66 (.A2( u1_u15_u3_n100 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n113 ) );
  NAND2_X1 u1_u15_u3_U67 (.A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n153 ) , .A2( u1_u15_u3_n97 ) );
  NAND2_X1 u1_u15_u3_U68 (.A2( u1_u15_u3_n103 ) , .A1( u1_u15_u3_n104 ) , .ZN( u1_u15_u3_n130 ) );
  NAND2_X1 u1_u15_u3_U69 (.A2( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n144 ) , .A1( u1_u15_u3_n96 ) );
  OAI22_X1 u1_u15_u3_U7 (.B2( u1_u15_u3_n147 ) , .A2( u1_u15_u3_n148 ) , .ZN( u1_u15_u3_n160 ) , .B1( u1_u15_u3_n165 ) , .A1( u1_u15_u3_n168 ) );
  NAND2_X1 u1_u15_u3_U70 (.A1( u1_u15_u3_n102 ) , .A2( u1_u15_u3_n103 ) , .ZN( u1_u15_u3_n108 ) );
  NOR2_X1 u1_u15_u3_U71 (.A2( u1_u15_X_19 ) , .A1( u1_u15_X_20 ) , .ZN( u1_u15_u3_n99 ) );
  NOR2_X1 u1_u15_u3_U72 (.A2( u1_u15_X_21 ) , .A1( u1_u15_X_24 ) , .ZN( u1_u15_u3_n103 ) );
  NOR2_X1 u1_u15_u3_U73 (.A2( u1_u15_X_24 ) , .A1( u1_u15_u3_n171 ) , .ZN( u1_u15_u3_n97 ) );
  NOR2_X1 u1_u15_u3_U74 (.A2( u1_u15_X_23 ) , .ZN( u1_u15_u3_n141 ) , .A1( u1_u15_u3_n166 ) );
  NOR2_X1 u1_u15_u3_U75 (.A2( u1_u15_X_19 ) , .A1( u1_u15_u3_n172 ) , .ZN( u1_u15_u3_n96 ) );
  NAND2_X1 u1_u15_u3_U76 (.A1( u1_u15_X_22 ) , .A2( u1_u15_X_23 ) , .ZN( u1_u15_u3_n154 ) );
  NAND2_X1 u1_u15_u3_U77 (.A1( u1_u15_X_23 ) , .ZN( u1_u15_u3_n149 ) , .A2( u1_u15_u3_n166 ) );
  NOR2_X1 u1_u15_u3_U78 (.A2( u1_u15_X_22 ) , .A1( u1_u15_X_23 ) , .ZN( u1_u15_u3_n121 ) );
  AND2_X1 u1_u15_u3_U79 (.A1( u1_u15_X_24 ) , .ZN( u1_u15_u3_n101 ) , .A2( u1_u15_u3_n171 ) );
  AND3_X1 u1_u15_u3_U8 (.A3( u1_u15_u3_n144 ) , .A2( u1_u15_u3_n145 ) , .A1( u1_u15_u3_n146 ) , .ZN( u1_u15_u3_n147 ) );
  AND2_X1 u1_u15_u3_U80 (.A1( u1_u15_X_19 ) , .ZN( u1_u15_u3_n102 ) , .A2( u1_u15_u3_n172 ) );
  AND2_X1 u1_u15_u3_U81 (.A1( u1_u15_X_21 ) , .A2( u1_u15_X_24 ) , .ZN( u1_u15_u3_n100 ) );
  AND2_X1 u1_u15_u3_U82 (.A2( u1_u15_X_19 ) , .A1( u1_u15_X_20 ) , .ZN( u1_u15_u3_n104 ) );
  INV_X1 u1_u15_u3_U83 (.A( u1_u15_X_22 ) , .ZN( u1_u15_u3_n166 ) );
  INV_X1 u1_u15_u3_U84 (.A( u1_u15_X_21 ) , .ZN( u1_u15_u3_n171 ) );
  INV_X1 u1_u15_u3_U85 (.A( u1_u15_X_20 ) , .ZN( u1_u15_u3_n172 ) );
  OR4_X1 u1_u15_u3_U86 (.ZN( u1_out15_10 ) , .A4( u1_u15_u3_n136 ) , .A3( u1_u15_u3_n137 ) , .A1( u1_u15_u3_n138 ) , .A2( u1_u15_u3_n139 ) );
  OAI222_X1 u1_u15_u3_U87 (.C1( u1_u15_u3_n128 ) , .ZN( u1_u15_u3_n137 ) , .B1( u1_u15_u3_n148 ) , .A2( u1_u15_u3_n150 ) , .B2( u1_u15_u3_n154 ) , .C2( u1_u15_u3_n164 ) , .A1( u1_u15_u3_n167 ) );
  OAI221_X1 u1_u15_u3_U88 (.A( u1_u15_u3_n134 ) , .B2( u1_u15_u3_n135 ) , .ZN( u1_u15_u3_n136 ) , .C1( u1_u15_u3_n149 ) , .B1( u1_u15_u3_n151 ) , .C2( u1_u15_u3_n183 ) );
  NAND4_X1 u1_u15_u3_U89 (.ZN( u1_out15_1 ) , .A4( u1_u15_u3_n161 ) , .A3( u1_u15_u3_n162 ) , .A2( u1_u15_u3_n163 ) , .A1( u1_u15_u3_n185 ) );
  INV_X1 u1_u15_u3_U9 (.A( u1_u15_u3_n143 ) , .ZN( u1_u15_u3_n168 ) );
  NAND2_X1 u1_u15_u3_U90 (.ZN( u1_u15_u3_n163 ) , .A2( u1_u15_u3_n170 ) , .A1( u1_u15_u3_n176 ) );
  AOI22_X1 u1_u15_u3_U91 (.B2( u1_u15_u3_n140 ) , .B1( u1_u15_u3_n141 ) , .A2( u1_u15_u3_n142 ) , .ZN( u1_u15_u3_n162 ) , .A1( u1_u15_u3_n177 ) );
  NAND4_X1 u1_u15_u3_U92 (.ZN( u1_out15_26 ) , .A4( u1_u15_u3_n109 ) , .A3( u1_u15_u3_n110 ) , .A2( u1_u15_u3_n111 ) , .A1( u1_u15_u3_n173 ) );
  INV_X1 u1_u15_u3_U93 (.ZN( u1_u15_u3_n173 ) , .A( u1_u15_u3_n94 ) );
  OAI21_X1 u1_u15_u3_U94 (.ZN( u1_u15_u3_n111 ) , .B2( u1_u15_u3_n117 ) , .A( u1_u15_u3_n133 ) , .B1( u1_u15_u3_n176 ) );
  NAND4_X1 u1_u15_u3_U95 (.ZN( u1_out15_20 ) , .A4( u1_u15_u3_n122 ) , .A3( u1_u15_u3_n123 ) , .A1( u1_u15_u3_n175 ) , .A2( u1_u15_u3_n180 ) );
  INV_X1 u1_u15_u3_U96 (.A( u1_u15_u3_n126 ) , .ZN( u1_u15_u3_n180 ) );
  INV_X1 u1_u15_u3_U97 (.A( u1_u15_u3_n112 ) , .ZN( u1_u15_u3_n175 ) );
  NAND3_X1 u1_u15_u3_U98 (.A1( u1_u15_u3_n114 ) , .ZN( u1_u15_u3_n115 ) , .A2( u1_u15_u3_n145 ) , .A3( u1_u15_u3_n153 ) );
  NAND3_X1 u1_u15_u3_U99 (.ZN( u1_u15_u3_n129 ) , .A2( u1_u15_u3_n144 ) , .A1( u1_u15_u3_n153 ) , .A3( u1_u15_u3_n182 ) );
  OAI22_X1 u1_u15_u4_U10 (.B2( u1_u15_u4_n135 ) , .ZN( u1_u15_u4_n137 ) , .B1( u1_u15_u4_n153 ) , .A1( u1_u15_u4_n155 ) , .A2( u1_u15_u4_n171 ) );
  AND3_X1 u1_u15_u4_U11 (.A2( u1_u15_u4_n134 ) , .ZN( u1_u15_u4_n135 ) , .A3( u1_u15_u4_n145 ) , .A1( u1_u15_u4_n157 ) );
  NAND2_X1 u1_u15_u4_U12 (.ZN( u1_u15_u4_n132 ) , .A2( u1_u15_u4_n170 ) , .A1( u1_u15_u4_n173 ) );
  AOI21_X1 u1_u15_u4_U13 (.B2( u1_u15_u4_n160 ) , .B1( u1_u15_u4_n161 ) , .ZN( u1_u15_u4_n162 ) , .A( u1_u15_u4_n170 ) );
  AOI21_X1 u1_u15_u4_U14 (.ZN( u1_u15_u4_n107 ) , .B2( u1_u15_u4_n143 ) , .A( u1_u15_u4_n174 ) , .B1( u1_u15_u4_n184 ) );
  AOI21_X1 u1_u15_u4_U15 (.B2( u1_u15_u4_n158 ) , .B1( u1_u15_u4_n159 ) , .ZN( u1_u15_u4_n163 ) , .A( u1_u15_u4_n174 ) );
  AOI21_X1 u1_u15_u4_U16 (.A( u1_u15_u4_n153 ) , .B2( u1_u15_u4_n154 ) , .B1( u1_u15_u4_n155 ) , .ZN( u1_u15_u4_n165 ) );
  AOI21_X1 u1_u15_u4_U17 (.A( u1_u15_u4_n156 ) , .B2( u1_u15_u4_n157 ) , .ZN( u1_u15_u4_n164 ) , .B1( u1_u15_u4_n184 ) );
  INV_X1 u1_u15_u4_U18 (.A( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n170 ) );
  AND2_X1 u1_u15_u4_U19 (.A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n155 ) , .A1( u1_u15_u4_n160 ) );
  INV_X1 u1_u15_u4_U20 (.A( u1_u15_u4_n156 ) , .ZN( u1_u15_u4_n175 ) );
  NAND2_X1 u1_u15_u4_U21 (.A2( u1_u15_u4_n118 ) , .ZN( u1_u15_u4_n131 ) , .A1( u1_u15_u4_n147 ) );
  NAND2_X1 u1_u15_u4_U22 (.A1( u1_u15_u4_n119 ) , .A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n130 ) );
  NAND2_X1 u1_u15_u4_U23 (.ZN( u1_u15_u4_n117 ) , .A2( u1_u15_u4_n118 ) , .A1( u1_u15_u4_n148 ) );
  NAND2_X1 u1_u15_u4_U24 (.ZN( u1_u15_u4_n129 ) , .A1( u1_u15_u4_n134 ) , .A2( u1_u15_u4_n148 ) );
  AND3_X1 u1_u15_u4_U25 (.A1( u1_u15_u4_n119 ) , .A2( u1_u15_u4_n143 ) , .A3( u1_u15_u4_n154 ) , .ZN( u1_u15_u4_n161 ) );
  AND2_X1 u1_u15_u4_U26 (.A1( u1_u15_u4_n145 ) , .A2( u1_u15_u4_n147 ) , .ZN( u1_u15_u4_n159 ) );
  OR3_X1 u1_u15_u4_U27 (.A3( u1_u15_u4_n114 ) , .A2( u1_u15_u4_n115 ) , .A1( u1_u15_u4_n116 ) , .ZN( u1_u15_u4_n136 ) );
  AOI21_X1 u1_u15_u4_U28 (.A( u1_u15_u4_n113 ) , .ZN( u1_u15_u4_n116 ) , .B2( u1_u15_u4_n173 ) , .B1( u1_u15_u4_n174 ) );
  AOI21_X1 u1_u15_u4_U29 (.ZN( u1_u15_u4_n115 ) , .B2( u1_u15_u4_n145 ) , .B1( u1_u15_u4_n146 ) , .A( u1_u15_u4_n156 ) );
  NOR2_X1 u1_u15_u4_U3 (.ZN( u1_u15_u4_n121 ) , .A1( u1_u15_u4_n181 ) , .A2( u1_u15_u4_n182 ) );
  OAI22_X1 u1_u15_u4_U30 (.ZN( u1_u15_u4_n114 ) , .A2( u1_u15_u4_n121 ) , .B1( u1_u15_u4_n160 ) , .B2( u1_u15_u4_n170 ) , .A1( u1_u15_u4_n171 ) );
  INV_X1 u1_u15_u4_U31 (.A( u1_u15_u4_n158 ) , .ZN( u1_u15_u4_n182 ) );
  INV_X1 u1_u15_u4_U32 (.ZN( u1_u15_u4_n181 ) , .A( u1_u15_u4_n96 ) );
  INV_X1 u1_u15_u4_U33 (.A( u1_u15_u4_n144 ) , .ZN( u1_u15_u4_n179 ) );
  INV_X1 u1_u15_u4_U34 (.A( u1_u15_u4_n157 ) , .ZN( u1_u15_u4_n178 ) );
  NAND2_X1 u1_u15_u4_U35 (.A2( u1_u15_u4_n154 ) , .A1( u1_u15_u4_n96 ) , .ZN( u1_u15_u4_n97 ) );
  INV_X1 u1_u15_u4_U36 (.ZN( u1_u15_u4_n186 ) , .A( u1_u15_u4_n95 ) );
  OAI221_X1 u1_u15_u4_U37 (.C1( u1_u15_u4_n134 ) , .B1( u1_u15_u4_n158 ) , .B2( u1_u15_u4_n171 ) , .C2( u1_u15_u4_n173 ) , .A( u1_u15_u4_n94 ) , .ZN( u1_u15_u4_n95 ) );
  AOI222_X1 u1_u15_u4_U38 (.B2( u1_u15_u4_n132 ) , .A1( u1_u15_u4_n138 ) , .C2( u1_u15_u4_n175 ) , .A2( u1_u15_u4_n179 ) , .C1( u1_u15_u4_n181 ) , .B1( u1_u15_u4_n185 ) , .ZN( u1_u15_u4_n94 ) );
  INV_X1 u1_u15_u4_U39 (.A( u1_u15_u4_n113 ) , .ZN( u1_u15_u4_n185 ) );
  INV_X1 u1_u15_u4_U4 (.A( u1_u15_u4_n117 ) , .ZN( u1_u15_u4_n184 ) );
  INV_X1 u1_u15_u4_U40 (.A( u1_u15_u4_n143 ) , .ZN( u1_u15_u4_n183 ) );
  NOR2_X1 u1_u15_u4_U41 (.ZN( u1_u15_u4_n138 ) , .A1( u1_u15_u4_n168 ) , .A2( u1_u15_u4_n169 ) );
  NOR2_X1 u1_u15_u4_U42 (.A1( u1_u15_u4_n150 ) , .A2( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n153 ) );
  NOR2_X1 u1_u15_u4_U43 (.A2( u1_u15_u4_n128 ) , .A1( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n156 ) );
  AOI22_X1 u1_u15_u4_U44 (.B2( u1_u15_u4_n122 ) , .A1( u1_u15_u4_n123 ) , .ZN( u1_u15_u4_n124 ) , .B1( u1_u15_u4_n128 ) , .A2( u1_u15_u4_n172 ) );
  NAND2_X1 u1_u15_u4_U45 (.A2( u1_u15_u4_n120 ) , .ZN( u1_u15_u4_n123 ) , .A1( u1_u15_u4_n161 ) );
  INV_X1 u1_u15_u4_U46 (.A( u1_u15_u4_n153 ) , .ZN( u1_u15_u4_n172 ) );
  AOI22_X1 u1_u15_u4_U47 (.B2( u1_u15_u4_n132 ) , .A2( u1_u15_u4_n133 ) , .ZN( u1_u15_u4_n140 ) , .A1( u1_u15_u4_n150 ) , .B1( u1_u15_u4_n179 ) );
  NAND2_X1 u1_u15_u4_U48 (.ZN( u1_u15_u4_n133 ) , .A2( u1_u15_u4_n146 ) , .A1( u1_u15_u4_n154 ) );
  NAND2_X1 u1_u15_u4_U49 (.A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n154 ) , .A2( u1_u15_u4_n98 ) );
  NOR4_X1 u1_u15_u4_U5 (.A4( u1_u15_u4_n106 ) , .A3( u1_u15_u4_n107 ) , .A2( u1_u15_u4_n108 ) , .A1( u1_u15_u4_n109 ) , .ZN( u1_u15_u4_n110 ) );
  NAND2_X1 u1_u15_u4_U50 (.A1( u1_u15_u4_n101 ) , .ZN( u1_u15_u4_n158 ) , .A2( u1_u15_u4_n99 ) );
  AOI21_X1 u1_u15_u4_U51 (.ZN( u1_u15_u4_n127 ) , .A( u1_u15_u4_n136 ) , .B2( u1_u15_u4_n150 ) , .B1( u1_u15_u4_n180 ) );
  INV_X1 u1_u15_u4_U52 (.A( u1_u15_u4_n160 ) , .ZN( u1_u15_u4_n180 ) );
  NAND2_X1 u1_u15_u4_U53 (.A2( u1_u15_u4_n104 ) , .A1( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n146 ) );
  NAND2_X1 u1_u15_u4_U54 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n160 ) );
  NAND2_X1 u1_u15_u4_U55 (.ZN( u1_u15_u4_n134 ) , .A1( u1_u15_u4_n98 ) , .A2( u1_u15_u4_n99 ) );
  NAND2_X1 u1_u15_u4_U56 (.A1( u1_u15_u4_n103 ) , .A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n143 ) );
  NAND2_X1 u1_u15_u4_U57 (.A2( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n145 ) , .A1( u1_u15_u4_n98 ) );
  NAND2_X1 u1_u15_u4_U58 (.A1( u1_u15_u4_n100 ) , .A2( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n120 ) );
  NAND2_X1 u1_u15_u4_U59 (.A1( u1_u15_u4_n102 ) , .A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n148 ) );
  AOI21_X1 u1_u15_u4_U6 (.ZN( u1_u15_u4_n106 ) , .B2( u1_u15_u4_n146 ) , .B1( u1_u15_u4_n158 ) , .A( u1_u15_u4_n170 ) );
  NAND2_X1 u1_u15_u4_U60 (.A2( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n157 ) );
  INV_X1 u1_u15_u4_U61 (.A( u1_u15_u4_n150 ) , .ZN( u1_u15_u4_n173 ) );
  INV_X1 u1_u15_u4_U62 (.A( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n171 ) );
  NAND2_X1 u1_u15_u4_U63 (.A1( u1_u15_u4_n100 ) , .ZN( u1_u15_u4_n118 ) , .A2( u1_u15_u4_n99 ) );
  NAND2_X1 u1_u15_u4_U64 (.A2( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n144 ) );
  NAND2_X1 u1_u15_u4_U65 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n105 ) , .ZN( u1_u15_u4_n96 ) );
  INV_X1 u1_u15_u4_U66 (.A( u1_u15_u4_n128 ) , .ZN( u1_u15_u4_n174 ) );
  NAND2_X1 u1_u15_u4_U67 (.A2( u1_u15_u4_n102 ) , .ZN( u1_u15_u4_n119 ) , .A1( u1_u15_u4_n98 ) );
  NAND2_X1 u1_u15_u4_U68 (.A2( u1_u15_u4_n101 ) , .A1( u1_u15_u4_n103 ) , .ZN( u1_u15_u4_n147 ) );
  NAND2_X1 u1_u15_u4_U69 (.A2( u1_u15_u4_n104 ) , .ZN( u1_u15_u4_n113 ) , .A1( u1_u15_u4_n99 ) );
  AOI21_X1 u1_u15_u4_U7 (.ZN( u1_u15_u4_n108 ) , .B2( u1_u15_u4_n134 ) , .B1( u1_u15_u4_n155 ) , .A( u1_u15_u4_n156 ) );
  NOR2_X1 u1_u15_u4_U70 (.A2( u1_u15_X_28 ) , .ZN( u1_u15_u4_n150 ) , .A1( u1_u15_u4_n168 ) );
  NOR2_X1 u1_u15_u4_U71 (.A2( u1_u15_X_29 ) , .ZN( u1_u15_u4_n152 ) , .A1( u1_u15_u4_n169 ) );
  NOR2_X1 u1_u15_u4_U72 (.A2( u1_u15_X_26 ) , .ZN( u1_u15_u4_n100 ) , .A1( u1_u15_u4_n177 ) );
  NOR2_X1 u1_u15_u4_U73 (.A2( u1_u15_X_30 ) , .ZN( u1_u15_u4_n105 ) , .A1( u1_u15_u4_n176 ) );
  NOR2_X1 u1_u15_u4_U74 (.A2( u1_u15_X_28 ) , .A1( u1_u15_X_29 ) , .ZN( u1_u15_u4_n128 ) );
  NOR2_X1 u1_u15_u4_U75 (.A2( u1_u15_X_25 ) , .A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n98 ) );
  NOR2_X1 u1_u15_u4_U76 (.A2( u1_u15_X_27 ) , .A1( u1_u15_X_30 ) , .ZN( u1_u15_u4_n102 ) );
  AND2_X1 u1_u15_u4_U77 (.A2( u1_u15_X_25 ) , .A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n104 ) );
  AND2_X1 u1_u15_u4_U78 (.A1( u1_u15_X_30 ) , .A2( u1_u15_u4_n176 ) , .ZN( u1_u15_u4_n99 ) );
  AND2_X1 u1_u15_u4_U79 (.A1( u1_u15_X_26 ) , .ZN( u1_u15_u4_n101 ) , .A2( u1_u15_u4_n177 ) );
  AOI21_X1 u1_u15_u4_U8 (.ZN( u1_u15_u4_n109 ) , .A( u1_u15_u4_n153 ) , .B1( u1_u15_u4_n159 ) , .B2( u1_u15_u4_n184 ) );
  AND2_X1 u1_u15_u4_U80 (.A1( u1_u15_X_27 ) , .A2( u1_u15_X_30 ) , .ZN( u1_u15_u4_n103 ) );
  INV_X1 u1_u15_u4_U81 (.A( u1_u15_X_28 ) , .ZN( u1_u15_u4_n169 ) );
  INV_X1 u1_u15_u4_U82 (.A( u1_u15_X_29 ) , .ZN( u1_u15_u4_n168 ) );
  INV_X1 u1_u15_u4_U83 (.A( u1_u15_X_25 ) , .ZN( u1_u15_u4_n177 ) );
  INV_X1 u1_u15_u4_U84 (.A( u1_u15_X_27 ) , .ZN( u1_u15_u4_n176 ) );
  NAND4_X1 u1_u15_u4_U85 (.ZN( u1_out15_25 ) , .A4( u1_u15_u4_n139 ) , .A3( u1_u15_u4_n140 ) , .A2( u1_u15_u4_n141 ) , .A1( u1_u15_u4_n142 ) );
  OAI21_X1 u1_u15_u4_U86 (.A( u1_u15_u4_n128 ) , .B2( u1_u15_u4_n129 ) , .B1( u1_u15_u4_n130 ) , .ZN( u1_u15_u4_n142 ) );
  OAI21_X1 u1_u15_u4_U87 (.B2( u1_u15_u4_n131 ) , .ZN( u1_u15_u4_n141 ) , .A( u1_u15_u4_n175 ) , .B1( u1_u15_u4_n183 ) );
  NAND4_X1 u1_u15_u4_U88 (.ZN( u1_out15_14 ) , .A4( u1_u15_u4_n124 ) , .A3( u1_u15_u4_n125 ) , .A2( u1_u15_u4_n126 ) , .A1( u1_u15_u4_n127 ) );
  AOI22_X1 u1_u15_u4_U89 (.B2( u1_u15_u4_n117 ) , .ZN( u1_u15_u4_n126 ) , .A1( u1_u15_u4_n129 ) , .B1( u1_u15_u4_n152 ) , .A2( u1_u15_u4_n175 ) );
  AOI211_X1 u1_u15_u4_U9 (.B( u1_u15_u4_n136 ) , .A( u1_u15_u4_n137 ) , .C2( u1_u15_u4_n138 ) , .ZN( u1_u15_u4_n139 ) , .C1( u1_u15_u4_n182 ) );
  AOI22_X1 u1_u15_u4_U90 (.ZN( u1_u15_u4_n125 ) , .B2( u1_u15_u4_n131 ) , .A2( u1_u15_u4_n132 ) , .B1( u1_u15_u4_n138 ) , .A1( u1_u15_u4_n178 ) );
  AOI22_X1 u1_u15_u4_U91 (.B2( u1_u15_u4_n149 ) , .B1( u1_u15_u4_n150 ) , .A2( u1_u15_u4_n151 ) , .A1( u1_u15_u4_n152 ) , .ZN( u1_u15_u4_n167 ) );
  NOR4_X1 u1_u15_u4_U92 (.A4( u1_u15_u4_n162 ) , .A3( u1_u15_u4_n163 ) , .A2( u1_u15_u4_n164 ) , .A1( u1_u15_u4_n165 ) , .ZN( u1_u15_u4_n166 ) );
  NAND4_X1 u1_u15_u4_U93 (.ZN( u1_out15_8 ) , .A4( u1_u15_u4_n110 ) , .A3( u1_u15_u4_n111 ) , .A2( u1_u15_u4_n112 ) , .A1( u1_u15_u4_n186 ) );
  NAND2_X1 u1_u15_u4_U94 (.ZN( u1_u15_u4_n112 ) , .A2( u1_u15_u4_n130 ) , .A1( u1_u15_u4_n150 ) );
  AOI22_X1 u1_u15_u4_U95 (.ZN( u1_u15_u4_n111 ) , .B2( u1_u15_u4_n132 ) , .A1( u1_u15_u4_n152 ) , .B1( u1_u15_u4_n178 ) , .A2( u1_u15_u4_n97 ) );
  NAND3_X1 u1_u15_u4_U96 (.ZN( u1_out15_3 ) , .A3( u1_u15_u4_n166 ) , .A1( u1_u15_u4_n167 ) , .A2( u1_u15_u4_n186 ) );
  NAND3_X1 u1_u15_u4_U97 (.A3( u1_u15_u4_n146 ) , .A2( u1_u15_u4_n147 ) , .A1( u1_u15_u4_n148 ) , .ZN( u1_u15_u4_n149 ) );
  NAND3_X1 u1_u15_u4_U98 (.A3( u1_u15_u4_n143 ) , .A2( u1_u15_u4_n144 ) , .A1( u1_u15_u4_n145 ) , .ZN( u1_u15_u4_n151 ) );
  NAND3_X1 u1_u15_u4_U99 (.A3( u1_u15_u4_n121 ) , .ZN( u1_u15_u4_n122 ) , .A2( u1_u15_u4_n144 ) , .A1( u1_u15_u4_n154 ) );
  XOR2_X1 u1_u1_U10 (.B( u1_K2_45 ) , .A( u1_R0_30 ) , .Z( u1_u1_X_45 ) );
  XOR2_X1 u1_u1_U11 (.B( u1_K2_44 ) , .A( u1_R0_29 ) , .Z( u1_u1_X_44 ) );
  XOR2_X1 u1_u1_U12 (.B( u1_K2_43 ) , .A( u1_R0_28 ) , .Z( u1_u1_X_43 ) );
  XOR2_X1 u1_u1_U13 (.B( u1_K2_42 ) , .A( u1_R0_29 ) , .Z( u1_u1_X_42 ) );
  XOR2_X1 u1_u1_U14 (.B( u1_K2_41 ) , .A( u1_R0_28 ) , .Z( u1_u1_X_41 ) );
  XOR2_X1 u1_u1_U15 (.B( u1_K2_40 ) , .A( u1_R0_27 ) , .Z( u1_u1_X_40 ) );
  XOR2_X1 u1_u1_U16 (.B( u1_K2_3 ) , .A( u1_R0_2 ) , .Z( u1_u1_X_3 ) );
  XOR2_X1 u1_u1_U17 (.B( u1_K2_39 ) , .A( u1_R0_26 ) , .Z( u1_u1_X_39 ) );
  XOR2_X1 u1_u1_U18 (.B( u1_K2_38 ) , .A( u1_R0_25 ) , .Z( u1_u1_X_38 ) );
  XOR2_X1 u1_u1_U19 (.B( u1_K2_37 ) , .A( u1_R0_24 ) , .Z( u1_u1_X_37 ) );
  XOR2_X1 u1_u1_U2 (.B( u1_K2_8 ) , .A( u1_R0_5 ) , .Z( u1_u1_X_8 ) );
  XOR2_X1 u1_u1_U20 (.B( u1_K2_36 ) , .A( u1_R0_25 ) , .Z( u1_u1_X_36 ) );
  XOR2_X1 u1_u1_U21 (.B( u1_K2_35 ) , .A( u1_R0_24 ) , .Z( u1_u1_X_35 ) );
  XOR2_X1 u1_u1_U24 (.B( u1_K2_32 ) , .A( u1_R0_21 ) , .Z( u1_u1_X_32 ) );
  XOR2_X1 u1_u1_U25 (.B( u1_K2_31 ) , .A( u1_R0_20 ) , .Z( u1_u1_X_31 ) );
  XOR2_X1 u1_u1_U26 (.B( u1_K2_30 ) , .A( u1_R0_21 ) , .Z( u1_u1_X_30 ) );
  XOR2_X1 u1_u1_U27 (.B( u1_K2_2 ) , .A( u1_R0_1 ) , .Z( u1_u1_X_2 ) );
  XOR2_X1 u1_u1_U28 (.B( u1_K2_29 ) , .A( u1_R0_20 ) , .Z( u1_u1_X_29 ) );
  XOR2_X1 u1_u1_U29 (.B( u1_K2_28 ) , .A( u1_R0_19 ) , .Z( u1_u1_X_28 ) );
  XOR2_X1 u1_u1_U3 (.B( u1_K2_7 ) , .A( u1_R0_4 ) , .Z( u1_u1_X_7 ) );
  XOR2_X1 u1_u1_U30 (.B( u1_K2_27 ) , .A( u1_R0_18 ) , .Z( u1_u1_X_27 ) );
  XOR2_X1 u1_u1_U31 (.B( u1_K2_26 ) , .A( u1_R0_17 ) , .Z( u1_u1_X_26 ) );
  XOR2_X1 u1_u1_U32 (.B( u1_K2_25 ) , .A( u1_R0_16 ) , .Z( u1_u1_X_25 ) );
  XOR2_X1 u1_u1_U33 (.B( u1_K2_24 ) , .A( u1_R0_17 ) , .Z( u1_u1_X_24 ) );
  XOR2_X1 u1_u1_U34 (.B( u1_K2_23 ) , .A( u1_R0_16 ) , .Z( u1_u1_X_23 ) );
  XOR2_X1 u1_u1_U35 (.B( u1_K2_22 ) , .A( u1_R0_15 ) , .Z( u1_u1_X_22 ) );
  XOR2_X1 u1_u1_U36 (.B( u1_K2_21 ) , .A( u1_R0_14 ) , .Z( u1_u1_X_21 ) );
  XOR2_X1 u1_u1_U37 (.B( u1_K2_20 ) , .A( u1_R0_13 ) , .Z( u1_u1_X_20 ) );
  XOR2_X1 u1_u1_U38 (.B( u1_K2_1 ) , .A( u1_R0_32 ) , .Z( u1_u1_X_1 ) );
  XOR2_X1 u1_u1_U39 (.B( u1_K2_19 ) , .A( u1_R0_12 ) , .Z( u1_u1_X_19 ) );
  XOR2_X1 u1_u1_U4 (.B( u1_K2_6 ) , .A( u1_R0_5 ) , .Z( u1_u1_X_6 ) );
  XOR2_X1 u1_u1_U40 (.B( u1_K2_18 ) , .A( u1_R0_13 ) , .Z( u1_u1_X_18 ) );
  XOR2_X1 u1_u1_U41 (.B( u1_K2_17 ) , .A( u1_R0_12 ) , .Z( u1_u1_X_17 ) );
  XOR2_X1 u1_u1_U42 (.B( u1_K2_16 ) , .A( u1_R0_11 ) , .Z( u1_u1_X_16 ) );
  XOR2_X1 u1_u1_U43 (.B( u1_K2_15 ) , .A( u1_R0_10 ) , .Z( u1_u1_X_15 ) );
  XOR2_X1 u1_u1_U44 (.B( u1_K2_14 ) , .A( u1_R0_9 ) , .Z( u1_u1_X_14 ) );
  XOR2_X1 u1_u1_U45 (.B( u1_K2_13 ) , .A( u1_R0_8 ) , .Z( u1_u1_X_13 ) );
  XOR2_X1 u1_u1_U46 (.B( u1_K2_12 ) , .A( u1_R0_9 ) , .Z( u1_u1_X_12 ) );
  XOR2_X1 u1_u1_U47 (.B( u1_K2_11 ) , .A( u1_R0_8 ) , .Z( u1_u1_X_11 ) );
  XOR2_X1 u1_u1_U5 (.B( u1_K2_5 ) , .A( u1_R0_4 ) , .Z( u1_u1_X_5 ) );
  XOR2_X1 u1_u1_U6 (.B( u1_K2_4 ) , .A( u1_R0_3 ) , .Z( u1_u1_X_4 ) );
  XOR2_X1 u1_u1_U7 (.B( u1_K2_48 ) , .A( u1_R0_1 ) , .Z( u1_u1_X_48 ) );
  XOR2_X1 u1_u1_U8 (.B( u1_K2_47 ) , .A( u1_R0_32 ) , .Z( u1_u1_X_47 ) );
  XOR2_X1 u1_u1_U9 (.B( u1_K2_46 ) , .A( u1_R0_31 ) , .Z( u1_u1_X_46 ) );
  AND3_X1 u1_u1_u0_U10 (.A2( u1_u1_u0_n112 ) , .ZN( u1_u1_u0_n127 ) , .A3( u1_u1_u0_n130 ) , .A1( u1_u1_u0_n148 ) );
  NAND2_X1 u1_u1_u0_U11 (.ZN( u1_u1_u0_n113 ) , .A1( u1_u1_u0_n139 ) , .A2( u1_u1_u0_n149 ) );
  AND2_X1 u1_u1_u0_U12 (.ZN( u1_u1_u0_n107 ) , .A1( u1_u1_u0_n130 ) , .A2( u1_u1_u0_n140 ) );
  AND2_X1 u1_u1_u0_U13 (.A2( u1_u1_u0_n129 ) , .A1( u1_u1_u0_n130 ) , .ZN( u1_u1_u0_n151 ) );
  AND2_X1 u1_u1_u0_U14 (.A1( u1_u1_u0_n108 ) , .A2( u1_u1_u0_n125 ) , .ZN( u1_u1_u0_n145 ) );
  INV_X1 u1_u1_u0_U15 (.A( u1_u1_u0_n143 ) , .ZN( u1_u1_u0_n173 ) );
  NOR2_X1 u1_u1_u0_U16 (.A2( u1_u1_u0_n136 ) , .ZN( u1_u1_u0_n147 ) , .A1( u1_u1_u0_n160 ) );
  NOR2_X1 u1_u1_u0_U17 (.A1( u1_u1_u0_n163 ) , .A2( u1_u1_u0_n164 ) , .ZN( u1_u1_u0_n95 ) );
  AOI21_X1 u1_u1_u0_U18 (.B1( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n132 ) , .A( u1_u1_u0_n165 ) , .B2( u1_u1_u0_n93 ) );
  INV_X1 u1_u1_u0_U19 (.A( u1_u1_u0_n142 ) , .ZN( u1_u1_u0_n165 ) );
  OAI221_X1 u1_u1_u0_U20 (.C1( u1_u1_u0_n121 ) , .ZN( u1_u1_u0_n122 ) , .B2( u1_u1_u0_n127 ) , .A( u1_u1_u0_n143 ) , .B1( u1_u1_u0_n144 ) , .C2( u1_u1_u0_n147 ) );
  OAI22_X1 u1_u1_u0_U21 (.B1( u1_u1_u0_n125 ) , .ZN( u1_u1_u0_n126 ) , .A1( u1_u1_u0_n138 ) , .A2( u1_u1_u0_n146 ) , .B2( u1_u1_u0_n147 ) );
  OAI22_X1 u1_u1_u0_U22 (.B1( u1_u1_u0_n131 ) , .A1( u1_u1_u0_n144 ) , .B2( u1_u1_u0_n147 ) , .A2( u1_u1_u0_n90 ) , .ZN( u1_u1_u0_n91 ) );
  AND3_X1 u1_u1_u0_U23 (.A3( u1_u1_u0_n121 ) , .A2( u1_u1_u0_n125 ) , .A1( u1_u1_u0_n148 ) , .ZN( u1_u1_u0_n90 ) );
  INV_X1 u1_u1_u0_U24 (.A( u1_u1_u0_n136 ) , .ZN( u1_u1_u0_n161 ) );
  NOR2_X1 u1_u1_u0_U25 (.A1( u1_u1_u0_n120 ) , .ZN( u1_u1_u0_n143 ) , .A2( u1_u1_u0_n167 ) );
  OAI221_X1 u1_u1_u0_U26 (.C1( u1_u1_u0_n112 ) , .ZN( u1_u1_u0_n120 ) , .B1( u1_u1_u0_n138 ) , .B2( u1_u1_u0_n141 ) , .C2( u1_u1_u0_n147 ) , .A( u1_u1_u0_n172 ) );
  AOI211_X1 u1_u1_u0_U27 (.B( u1_u1_u0_n115 ) , .A( u1_u1_u0_n116 ) , .C2( u1_u1_u0_n117 ) , .C1( u1_u1_u0_n118 ) , .ZN( u1_u1_u0_n119 ) );
  AOI22_X1 u1_u1_u0_U28 (.B2( u1_u1_u0_n109 ) , .A2( u1_u1_u0_n110 ) , .ZN( u1_u1_u0_n111 ) , .B1( u1_u1_u0_n118 ) , .A1( u1_u1_u0_n160 ) );
  INV_X1 u1_u1_u0_U29 (.A( u1_u1_u0_n118 ) , .ZN( u1_u1_u0_n158 ) );
  INV_X1 u1_u1_u0_U3 (.A( u1_u1_u0_n113 ) , .ZN( u1_u1_u0_n166 ) );
  AOI21_X1 u1_u1_u0_U30 (.ZN( u1_u1_u0_n104 ) , .B1( u1_u1_u0_n107 ) , .B2( u1_u1_u0_n141 ) , .A( u1_u1_u0_n144 ) );
  AOI21_X1 u1_u1_u0_U31 (.B1( u1_u1_u0_n127 ) , .B2( u1_u1_u0_n129 ) , .A( u1_u1_u0_n138 ) , .ZN( u1_u1_u0_n96 ) );
  AOI21_X1 u1_u1_u0_U32 (.ZN( u1_u1_u0_n116 ) , .B2( u1_u1_u0_n142 ) , .A( u1_u1_u0_n144 ) , .B1( u1_u1_u0_n166 ) );
  NAND2_X1 u1_u1_u0_U33 (.A1( u1_u1_u0_n100 ) , .A2( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n125 ) );
  NAND2_X1 u1_u1_u0_U34 (.A2( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n140 ) , .A1( u1_u1_u0_n94 ) );
  NAND2_X1 u1_u1_u0_U35 (.A1( u1_u1_u0_n101 ) , .A2( u1_u1_u0_n102 ) , .ZN( u1_u1_u0_n150 ) );
  INV_X1 u1_u1_u0_U36 (.A( u1_u1_u0_n138 ) , .ZN( u1_u1_u0_n160 ) );
  NAND2_X1 u1_u1_u0_U37 (.ZN( u1_u1_u0_n142 ) , .A1( u1_u1_u0_n94 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U38 (.A1( u1_u1_u0_n102 ) , .ZN( u1_u1_u0_n128 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U39 (.A2( u1_u1_u0_n102 ) , .A1( u1_u1_u0_n103 ) , .ZN( u1_u1_u0_n149 ) );
  AOI21_X1 u1_u1_u0_U4 (.B1( u1_u1_u0_n114 ) , .ZN( u1_u1_u0_n115 ) , .B2( u1_u1_u0_n129 ) , .A( u1_u1_u0_n161 ) );
  NAND2_X1 u1_u1_u0_U40 (.A1( u1_u1_u0_n100 ) , .ZN( u1_u1_u0_n129 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U41 (.A2( u1_u1_u0_n100 ) , .A1( u1_u1_u0_n101 ) , .ZN( u1_u1_u0_n139 ) );
  NAND2_X1 u1_u1_u0_U42 (.A2( u1_u1_u0_n100 ) , .ZN( u1_u1_u0_n131 ) , .A1( u1_u1_u0_n92 ) );
  NAND2_X1 u1_u1_u0_U43 (.ZN( u1_u1_u0_n108 ) , .A1( u1_u1_u0_n92 ) , .A2( u1_u1_u0_n94 ) );
  NAND2_X1 u1_u1_u0_U44 (.ZN( u1_u1_u0_n148 ) , .A1( u1_u1_u0_n93 ) , .A2( u1_u1_u0_n95 ) );
  NAND2_X1 u1_u1_u0_U45 (.A2( u1_u1_u0_n102 ) , .ZN( u1_u1_u0_n114 ) , .A1( u1_u1_u0_n92 ) );
  NAND2_X1 u1_u1_u0_U46 (.A1( u1_u1_u0_n101 ) , .ZN( u1_u1_u0_n130 ) , .A2( u1_u1_u0_n94 ) );
  NAND2_X1 u1_u1_u0_U47 (.A2( u1_u1_u0_n101 ) , .ZN( u1_u1_u0_n121 ) , .A1( u1_u1_u0_n93 ) );
  INV_X1 u1_u1_u0_U48 (.ZN( u1_u1_u0_n172 ) , .A( u1_u1_u0_n88 ) );
  OAI222_X1 u1_u1_u0_U49 (.C1( u1_u1_u0_n108 ) , .A1( u1_u1_u0_n125 ) , .B2( u1_u1_u0_n128 ) , .B1( u1_u1_u0_n144 ) , .A2( u1_u1_u0_n158 ) , .C2( u1_u1_u0_n161 ) , .ZN( u1_u1_u0_n88 ) );
  AOI21_X1 u1_u1_u0_U5 (.B2( u1_u1_u0_n131 ) , .ZN( u1_u1_u0_n134 ) , .B1( u1_u1_u0_n151 ) , .A( u1_u1_u0_n158 ) );
  NAND2_X1 u1_u1_u0_U50 (.ZN( u1_u1_u0_n112 ) , .A2( u1_u1_u0_n92 ) , .A1( u1_u1_u0_n93 ) );
  OR3_X1 u1_u1_u0_U51 (.A3( u1_u1_u0_n152 ) , .A2( u1_u1_u0_n153 ) , .A1( u1_u1_u0_n154 ) , .ZN( u1_u1_u0_n155 ) );
  AOI21_X1 u1_u1_u0_U52 (.B2( u1_u1_u0_n150 ) , .B1( u1_u1_u0_n151 ) , .ZN( u1_u1_u0_n152 ) , .A( u1_u1_u0_n158 ) );
  AOI21_X1 u1_u1_u0_U53 (.A( u1_u1_u0_n144 ) , .B2( u1_u1_u0_n145 ) , .B1( u1_u1_u0_n146 ) , .ZN( u1_u1_u0_n154 ) );
  AOI21_X1 u1_u1_u0_U54 (.A( u1_u1_u0_n147 ) , .B2( u1_u1_u0_n148 ) , .B1( u1_u1_u0_n149 ) , .ZN( u1_u1_u0_n153 ) );
  INV_X1 u1_u1_u0_U55 (.ZN( u1_u1_u0_n171 ) , .A( u1_u1_u0_n99 ) );
  OAI211_X1 u1_u1_u0_U56 (.C2( u1_u1_u0_n140 ) , .C1( u1_u1_u0_n161 ) , .A( u1_u1_u0_n169 ) , .B( u1_u1_u0_n98 ) , .ZN( u1_u1_u0_n99 ) );
  INV_X1 u1_u1_u0_U57 (.ZN( u1_u1_u0_n169 ) , .A( u1_u1_u0_n91 ) );
  AOI211_X1 u1_u1_u0_U58 (.C1( u1_u1_u0_n118 ) , .A( u1_u1_u0_n123 ) , .B( u1_u1_u0_n96 ) , .C2( u1_u1_u0_n97 ) , .ZN( u1_u1_u0_n98 ) );
  NOR2_X1 u1_u1_u0_U59 (.A2( u1_u1_X_2 ) , .ZN( u1_u1_u0_n103 ) , .A1( u1_u1_u0_n164 ) );
  NOR2_X1 u1_u1_u0_U6 (.A1( u1_u1_u0_n108 ) , .ZN( u1_u1_u0_n123 ) , .A2( u1_u1_u0_n158 ) );
  NOR2_X1 u1_u1_u0_U60 (.A2( u1_u1_X_3 ) , .A1( u1_u1_X_6 ) , .ZN( u1_u1_u0_n94 ) );
  NOR2_X1 u1_u1_u0_U61 (.A2( u1_u1_X_6 ) , .ZN( u1_u1_u0_n100 ) , .A1( u1_u1_u0_n162 ) );
  NOR2_X1 u1_u1_u0_U62 (.A2( u1_u1_X_4 ) , .A1( u1_u1_X_5 ) , .ZN( u1_u1_u0_n118 ) );
  NOR2_X1 u1_u1_u0_U63 (.A2( u1_u1_X_1 ) , .A1( u1_u1_X_2 ) , .ZN( u1_u1_u0_n92 ) );
  NOR2_X1 u1_u1_u0_U64 (.A2( u1_u1_X_1 ) , .ZN( u1_u1_u0_n101 ) , .A1( u1_u1_u0_n163 ) );
  NAND2_X1 u1_u1_u0_U65 (.A2( u1_u1_X_4 ) , .A1( u1_u1_X_5 ) , .ZN( u1_u1_u0_n144 ) );
  NOR2_X1 u1_u1_u0_U66 (.A2( u1_u1_X_5 ) , .ZN( u1_u1_u0_n136 ) , .A1( u1_u1_u0_n159 ) );
  NAND2_X1 u1_u1_u0_U67 (.A1( u1_u1_X_5 ) , .ZN( u1_u1_u0_n138 ) , .A2( u1_u1_u0_n159 ) );
  AND2_X1 u1_u1_u0_U68 (.A2( u1_u1_X_3 ) , .A1( u1_u1_X_6 ) , .ZN( u1_u1_u0_n102 ) );
  AND2_X1 u1_u1_u0_U69 (.A1( u1_u1_X_6 ) , .A2( u1_u1_u0_n162 ) , .ZN( u1_u1_u0_n93 ) );
  OAI21_X1 u1_u1_u0_U7 (.B1( u1_u1_u0_n150 ) , .B2( u1_u1_u0_n158 ) , .A( u1_u1_u0_n172 ) , .ZN( u1_u1_u0_n89 ) );
  INV_X1 u1_u1_u0_U70 (.A( u1_u1_X_4 ) , .ZN( u1_u1_u0_n159 ) );
  INV_X1 u1_u1_u0_U71 (.A( u1_u1_X_1 ) , .ZN( u1_u1_u0_n164 ) );
  INV_X1 u1_u1_u0_U72 (.A( u1_u1_X_2 ) , .ZN( u1_u1_u0_n163 ) );
  INV_X1 u1_u1_u0_U73 (.A( u1_u1_X_3 ) , .ZN( u1_u1_u0_n162 ) );
  INV_X1 u1_u1_u0_U74 (.A( u1_u1_u0_n126 ) , .ZN( u1_u1_u0_n168 ) );
  AOI211_X1 u1_u1_u0_U75 (.B( u1_u1_u0_n133 ) , .A( u1_u1_u0_n134 ) , .C2( u1_u1_u0_n135 ) , .C1( u1_u1_u0_n136 ) , .ZN( u1_u1_u0_n137 ) );
  INV_X1 u1_u1_u0_U76 (.ZN( u1_u1_u0_n174 ) , .A( u1_u1_u0_n89 ) );
  AOI211_X1 u1_u1_u0_U77 (.B( u1_u1_u0_n104 ) , .A( u1_u1_u0_n105 ) , .ZN( u1_u1_u0_n106 ) , .C2( u1_u1_u0_n113 ) , .C1( u1_u1_u0_n160 ) );
  OR4_X1 u1_u1_u0_U78 (.ZN( u1_out1_17 ) , .A4( u1_u1_u0_n122 ) , .A2( u1_u1_u0_n123 ) , .A1( u1_u1_u0_n124 ) , .A3( u1_u1_u0_n170 ) );
  AOI21_X1 u1_u1_u0_U79 (.B2( u1_u1_u0_n107 ) , .ZN( u1_u1_u0_n124 ) , .B1( u1_u1_u0_n128 ) , .A( u1_u1_u0_n161 ) );
  AND2_X1 u1_u1_u0_U8 (.A1( u1_u1_u0_n114 ) , .A2( u1_u1_u0_n121 ) , .ZN( u1_u1_u0_n146 ) );
  INV_X1 u1_u1_u0_U80 (.A( u1_u1_u0_n111 ) , .ZN( u1_u1_u0_n170 ) );
  OR4_X1 u1_u1_u0_U81 (.ZN( u1_out1_31 ) , .A4( u1_u1_u0_n155 ) , .A2( u1_u1_u0_n156 ) , .A1( u1_u1_u0_n157 ) , .A3( u1_u1_u0_n173 ) );
  AOI21_X1 u1_u1_u0_U82 (.A( u1_u1_u0_n138 ) , .B2( u1_u1_u0_n139 ) , .B1( u1_u1_u0_n140 ) , .ZN( u1_u1_u0_n157 ) );
  AOI21_X1 u1_u1_u0_U83 (.B2( u1_u1_u0_n141 ) , .B1( u1_u1_u0_n142 ) , .ZN( u1_u1_u0_n156 ) , .A( u1_u1_u0_n161 ) );
  AOI21_X1 u1_u1_u0_U84 (.B1( u1_u1_u0_n132 ) , .ZN( u1_u1_u0_n133 ) , .A( u1_u1_u0_n144 ) , .B2( u1_u1_u0_n166 ) );
  OAI22_X1 u1_u1_u0_U85 (.ZN( u1_u1_u0_n105 ) , .A2( u1_u1_u0_n132 ) , .B1( u1_u1_u0_n146 ) , .A1( u1_u1_u0_n147 ) , .B2( u1_u1_u0_n161 ) );
  NAND2_X1 u1_u1_u0_U86 (.ZN( u1_u1_u0_n110 ) , .A2( u1_u1_u0_n132 ) , .A1( u1_u1_u0_n145 ) );
  INV_X1 u1_u1_u0_U87 (.A( u1_u1_u0_n119 ) , .ZN( u1_u1_u0_n167 ) );
  NAND3_X1 u1_u1_u0_U88 (.ZN( u1_out1_23 ) , .A3( u1_u1_u0_n137 ) , .A1( u1_u1_u0_n168 ) , .A2( u1_u1_u0_n171 ) );
  NAND3_X1 u1_u1_u0_U89 (.A3( u1_u1_u0_n127 ) , .A2( u1_u1_u0_n128 ) , .ZN( u1_u1_u0_n135 ) , .A1( u1_u1_u0_n150 ) );
  AND2_X1 u1_u1_u0_U9 (.A1( u1_u1_u0_n131 ) , .ZN( u1_u1_u0_n141 ) , .A2( u1_u1_u0_n150 ) );
  NAND3_X1 u1_u1_u0_U90 (.ZN( u1_u1_u0_n117 ) , .A3( u1_u1_u0_n132 ) , .A2( u1_u1_u0_n139 ) , .A1( u1_u1_u0_n148 ) );
  NAND3_X1 u1_u1_u0_U91 (.ZN( u1_u1_u0_n109 ) , .A2( u1_u1_u0_n114 ) , .A3( u1_u1_u0_n140 ) , .A1( u1_u1_u0_n149 ) );
  NAND3_X1 u1_u1_u0_U92 (.ZN( u1_out1_9 ) , .A3( u1_u1_u0_n106 ) , .A2( u1_u1_u0_n171 ) , .A1( u1_u1_u0_n174 ) );
  NAND3_X1 u1_u1_u0_U93 (.A2( u1_u1_u0_n128 ) , .A1( u1_u1_u0_n132 ) , .A3( u1_u1_u0_n146 ) , .ZN( u1_u1_u0_n97 ) );
  OAI22_X1 u1_u1_u2_U10 (.ZN( u1_u1_u2_n109 ) , .A2( u1_u1_u2_n113 ) , .B2( u1_u1_u2_n133 ) , .B1( u1_u1_u2_n167 ) , .A1( u1_u1_u2_n168 ) );
  NAND3_X1 u1_u1_u2_U100 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n104 ) , .A3( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n98 ) );
  OAI22_X1 u1_u1_u2_U11 (.B1( u1_u1_u2_n151 ) , .A2( u1_u1_u2_n152 ) , .A1( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n160 ) , .B2( u1_u1_u2_n168 ) );
  NOR3_X1 u1_u1_u2_U12 (.A1( u1_u1_u2_n150 ) , .ZN( u1_u1_u2_n151 ) , .A3( u1_u1_u2_n175 ) , .A2( u1_u1_u2_n188 ) );
  AOI21_X1 u1_u1_u2_U13 (.ZN( u1_u1_u2_n144 ) , .B2( u1_u1_u2_n155 ) , .A( u1_u1_u2_n172 ) , .B1( u1_u1_u2_n185 ) );
  AOI21_X1 u1_u1_u2_U14 (.B2( u1_u1_u2_n143 ) , .ZN( u1_u1_u2_n145 ) , .B1( u1_u1_u2_n152 ) , .A( u1_u1_u2_n171 ) );
  AOI21_X1 u1_u1_u2_U15 (.B2( u1_u1_u2_n120 ) , .B1( u1_u1_u2_n121 ) , .ZN( u1_u1_u2_n126 ) , .A( u1_u1_u2_n167 ) );
  INV_X1 u1_u1_u2_U16 (.A( u1_u1_u2_n156 ) , .ZN( u1_u1_u2_n171 ) );
  INV_X1 u1_u1_u2_U17 (.A( u1_u1_u2_n120 ) , .ZN( u1_u1_u2_n188 ) );
  NAND2_X1 u1_u1_u2_U18 (.A2( u1_u1_u2_n122 ) , .ZN( u1_u1_u2_n150 ) , .A1( u1_u1_u2_n152 ) );
  INV_X1 u1_u1_u2_U19 (.A( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n170 ) );
  INV_X1 u1_u1_u2_U20 (.A( u1_u1_u2_n137 ) , .ZN( u1_u1_u2_n173 ) );
  NAND2_X1 u1_u1_u2_U21 (.A1( u1_u1_u2_n132 ) , .A2( u1_u1_u2_n139 ) , .ZN( u1_u1_u2_n157 ) );
  INV_X1 u1_u1_u2_U22 (.A( u1_u1_u2_n113 ) , .ZN( u1_u1_u2_n178 ) );
  INV_X1 u1_u1_u2_U23 (.A( u1_u1_u2_n139 ) , .ZN( u1_u1_u2_n175 ) );
  INV_X1 u1_u1_u2_U24 (.A( u1_u1_u2_n155 ) , .ZN( u1_u1_u2_n181 ) );
  INV_X1 u1_u1_u2_U25 (.A( u1_u1_u2_n119 ) , .ZN( u1_u1_u2_n177 ) );
  INV_X1 u1_u1_u2_U26 (.A( u1_u1_u2_n116 ) , .ZN( u1_u1_u2_n180 ) );
  INV_X1 u1_u1_u2_U27 (.A( u1_u1_u2_n131 ) , .ZN( u1_u1_u2_n179 ) );
  INV_X1 u1_u1_u2_U28 (.A( u1_u1_u2_n154 ) , .ZN( u1_u1_u2_n176 ) );
  NAND2_X1 u1_u1_u2_U29 (.A2( u1_u1_u2_n116 ) , .A1( u1_u1_u2_n117 ) , .ZN( u1_u1_u2_n118 ) );
  NOR2_X1 u1_u1_u2_U3 (.ZN( u1_u1_u2_n121 ) , .A2( u1_u1_u2_n177 ) , .A1( u1_u1_u2_n180 ) );
  INV_X1 u1_u1_u2_U30 (.A( u1_u1_u2_n132 ) , .ZN( u1_u1_u2_n182 ) );
  INV_X1 u1_u1_u2_U31 (.A( u1_u1_u2_n158 ) , .ZN( u1_u1_u2_n183 ) );
  OAI21_X1 u1_u1_u2_U32 (.A( u1_u1_u2_n156 ) , .B1( u1_u1_u2_n157 ) , .ZN( u1_u1_u2_n158 ) , .B2( u1_u1_u2_n179 ) );
  NOR2_X1 u1_u1_u2_U33 (.ZN( u1_u1_u2_n156 ) , .A1( u1_u1_u2_n166 ) , .A2( u1_u1_u2_n169 ) );
  NOR2_X1 u1_u1_u2_U34 (.A2( u1_u1_u2_n114 ) , .ZN( u1_u1_u2_n137 ) , .A1( u1_u1_u2_n140 ) );
  NOR2_X1 u1_u1_u2_U35 (.A2( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n153 ) , .A1( u1_u1_u2_n156 ) );
  AOI211_X1 u1_u1_u2_U36 (.ZN( u1_u1_u2_n130 ) , .C1( u1_u1_u2_n138 ) , .C2( u1_u1_u2_n179 ) , .B( u1_u1_u2_n96 ) , .A( u1_u1_u2_n97 ) );
  OAI22_X1 u1_u1_u2_U37 (.B1( u1_u1_u2_n133 ) , .A2( u1_u1_u2_n137 ) , .A1( u1_u1_u2_n152 ) , .B2( u1_u1_u2_n168 ) , .ZN( u1_u1_u2_n97 ) );
  OAI221_X1 u1_u1_u2_U38 (.B1( u1_u1_u2_n113 ) , .C1( u1_u1_u2_n132 ) , .A( u1_u1_u2_n149 ) , .B2( u1_u1_u2_n171 ) , .C2( u1_u1_u2_n172 ) , .ZN( u1_u1_u2_n96 ) );
  OAI221_X1 u1_u1_u2_U39 (.A( u1_u1_u2_n115 ) , .C2( u1_u1_u2_n123 ) , .B2( u1_u1_u2_n143 ) , .B1( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n163 ) , .C1( u1_u1_u2_n168 ) );
  INV_X1 u1_u1_u2_U4 (.A( u1_u1_u2_n134 ) , .ZN( u1_u1_u2_n185 ) );
  OAI21_X1 u1_u1_u2_U40 (.A( u1_u1_u2_n114 ) , .ZN( u1_u1_u2_n115 ) , .B1( u1_u1_u2_n176 ) , .B2( u1_u1_u2_n178 ) );
  OAI221_X1 u1_u1_u2_U41 (.A( u1_u1_u2_n135 ) , .B2( u1_u1_u2_n136 ) , .B1( u1_u1_u2_n137 ) , .ZN( u1_u1_u2_n162 ) , .C2( u1_u1_u2_n167 ) , .C1( u1_u1_u2_n185 ) );
  AND3_X1 u1_u1_u2_U42 (.A3( u1_u1_u2_n131 ) , .A2( u1_u1_u2_n132 ) , .A1( u1_u1_u2_n133 ) , .ZN( u1_u1_u2_n136 ) );
  AOI22_X1 u1_u1_u2_U43 (.ZN( u1_u1_u2_n135 ) , .B1( u1_u1_u2_n140 ) , .A1( u1_u1_u2_n156 ) , .B2( u1_u1_u2_n180 ) , .A2( u1_u1_u2_n188 ) );
  AOI21_X1 u1_u1_u2_U44 (.ZN( u1_u1_u2_n149 ) , .B1( u1_u1_u2_n173 ) , .B2( u1_u1_u2_n188 ) , .A( u1_u1_u2_n95 ) );
  AND3_X1 u1_u1_u2_U45 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n104 ) , .A3( u1_u1_u2_n156 ) , .ZN( u1_u1_u2_n95 ) );
  OAI21_X1 u1_u1_u2_U46 (.A( u1_u1_u2_n101 ) , .B2( u1_u1_u2_n121 ) , .B1( u1_u1_u2_n153 ) , .ZN( u1_u1_u2_n164 ) );
  NAND2_X1 u1_u1_u2_U47 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n107 ) , .ZN( u1_u1_u2_n155 ) );
  NAND2_X1 u1_u1_u2_U48 (.A2( u1_u1_u2_n105 ) , .A1( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n143 ) );
  NAND2_X1 u1_u1_u2_U49 (.A1( u1_u1_u2_n104 ) , .A2( u1_u1_u2_n106 ) , .ZN( u1_u1_u2_n152 ) );
  INV_X1 u1_u1_u2_U5 (.A( u1_u1_u2_n150 ) , .ZN( u1_u1_u2_n184 ) );
  NAND2_X1 u1_u1_u2_U50 (.A1( u1_u1_u2_n100 ) , .A2( u1_u1_u2_n105 ) , .ZN( u1_u1_u2_n132 ) );
  INV_X1 u1_u1_u2_U51 (.A( u1_u1_u2_n140 ) , .ZN( u1_u1_u2_n168 ) );
  INV_X1 u1_u1_u2_U52 (.A( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n167 ) );
  OAI21_X1 u1_u1_u2_U53 (.A( u1_u1_u2_n141 ) , .B2( u1_u1_u2_n142 ) , .ZN( u1_u1_u2_n146 ) , .B1( u1_u1_u2_n153 ) );
  OAI21_X1 u1_u1_u2_U54 (.A( u1_u1_u2_n140 ) , .ZN( u1_u1_u2_n141 ) , .B1( u1_u1_u2_n176 ) , .B2( u1_u1_u2_n177 ) );
  NOR3_X1 u1_u1_u2_U55 (.ZN( u1_u1_u2_n142 ) , .A3( u1_u1_u2_n175 ) , .A2( u1_u1_u2_n178 ) , .A1( u1_u1_u2_n181 ) );
  NAND2_X1 u1_u1_u2_U56 (.A1( u1_u1_u2_n102 ) , .A2( u1_u1_u2_n106 ) , .ZN( u1_u1_u2_n113 ) );
  NAND2_X1 u1_u1_u2_U57 (.A1( u1_u1_u2_n106 ) , .A2( u1_u1_u2_n107 ) , .ZN( u1_u1_u2_n131 ) );
  NAND2_X1 u1_u1_u2_U58 (.A1( u1_u1_u2_n103 ) , .A2( u1_u1_u2_n107 ) , .ZN( u1_u1_u2_n139 ) );
  NAND2_X1 u1_u1_u2_U59 (.A1( u1_u1_u2_n103 ) , .A2( u1_u1_u2_n105 ) , .ZN( u1_u1_u2_n133 ) );
  NOR4_X1 u1_u1_u2_U6 (.A4( u1_u1_u2_n124 ) , .A3( u1_u1_u2_n125 ) , .A2( u1_u1_u2_n126 ) , .A1( u1_u1_u2_n127 ) , .ZN( u1_u1_u2_n128 ) );
  NAND2_X1 u1_u1_u2_U60 (.A1( u1_u1_u2_n102 ) , .A2( u1_u1_u2_n103 ) , .ZN( u1_u1_u2_n154 ) );
  NAND2_X1 u1_u1_u2_U61 (.A2( u1_u1_u2_n103 ) , .A1( u1_u1_u2_n104 ) , .ZN( u1_u1_u2_n119 ) );
  NAND2_X1 u1_u1_u2_U62 (.A2( u1_u1_u2_n107 ) , .A1( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n123 ) );
  NAND2_X1 u1_u1_u2_U63 (.A1( u1_u1_u2_n104 ) , .A2( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n122 ) );
  INV_X1 u1_u1_u2_U64 (.A( u1_u1_u2_n114 ) , .ZN( u1_u1_u2_n172 ) );
  NAND2_X1 u1_u1_u2_U65 (.A2( u1_u1_u2_n100 ) , .A1( u1_u1_u2_n102 ) , .ZN( u1_u1_u2_n116 ) );
  NAND2_X1 u1_u1_u2_U66 (.A1( u1_u1_u2_n102 ) , .A2( u1_u1_u2_n108 ) , .ZN( u1_u1_u2_n120 ) );
  NAND2_X1 u1_u1_u2_U67 (.A2( u1_u1_u2_n105 ) , .A1( u1_u1_u2_n106 ) , .ZN( u1_u1_u2_n117 ) );
  INV_X1 u1_u1_u2_U68 (.ZN( u1_u1_u2_n187 ) , .A( u1_u1_u2_n99 ) );
  OAI21_X1 u1_u1_u2_U69 (.B1( u1_u1_u2_n137 ) , .B2( u1_u1_u2_n143 ) , .A( u1_u1_u2_n98 ) , .ZN( u1_u1_u2_n99 ) );
  AOI21_X1 u1_u1_u2_U7 (.B2( u1_u1_u2_n119 ) , .ZN( u1_u1_u2_n127 ) , .A( u1_u1_u2_n137 ) , .B1( u1_u1_u2_n155 ) );
  NOR2_X1 u1_u1_u2_U70 (.A2( u1_u1_X_16 ) , .ZN( u1_u1_u2_n140 ) , .A1( u1_u1_u2_n166 ) );
  NOR2_X1 u1_u1_u2_U71 (.A2( u1_u1_X_13 ) , .A1( u1_u1_X_14 ) , .ZN( u1_u1_u2_n100 ) );
  NOR2_X1 u1_u1_u2_U72 (.A2( u1_u1_X_16 ) , .A1( u1_u1_X_17 ) , .ZN( u1_u1_u2_n138 ) );
  NOR2_X1 u1_u1_u2_U73 (.A2( u1_u1_X_15 ) , .A1( u1_u1_X_18 ) , .ZN( u1_u1_u2_n104 ) );
  NOR2_X1 u1_u1_u2_U74 (.A2( u1_u1_X_14 ) , .ZN( u1_u1_u2_n103 ) , .A1( u1_u1_u2_n174 ) );
  NOR2_X1 u1_u1_u2_U75 (.A2( u1_u1_X_15 ) , .ZN( u1_u1_u2_n102 ) , .A1( u1_u1_u2_n165 ) );
  NOR2_X1 u1_u1_u2_U76 (.A2( u1_u1_X_17 ) , .ZN( u1_u1_u2_n114 ) , .A1( u1_u1_u2_n169 ) );
  AND2_X1 u1_u1_u2_U77 (.A1( u1_u1_X_15 ) , .ZN( u1_u1_u2_n105 ) , .A2( u1_u1_u2_n165 ) );
  AND2_X1 u1_u1_u2_U78 (.A2( u1_u1_X_15 ) , .A1( u1_u1_X_18 ) , .ZN( u1_u1_u2_n107 ) );
  AND2_X1 u1_u1_u2_U79 (.A1( u1_u1_X_14 ) , .ZN( u1_u1_u2_n106 ) , .A2( u1_u1_u2_n174 ) );
  AOI21_X1 u1_u1_u2_U8 (.ZN( u1_u1_u2_n124 ) , .B1( u1_u1_u2_n131 ) , .B2( u1_u1_u2_n143 ) , .A( u1_u1_u2_n172 ) );
  AND2_X1 u1_u1_u2_U80 (.A1( u1_u1_X_13 ) , .A2( u1_u1_X_14 ) , .ZN( u1_u1_u2_n108 ) );
  INV_X1 u1_u1_u2_U81 (.A( u1_u1_X_16 ) , .ZN( u1_u1_u2_n169 ) );
  INV_X1 u1_u1_u2_U82 (.A( u1_u1_X_17 ) , .ZN( u1_u1_u2_n166 ) );
  INV_X1 u1_u1_u2_U83 (.A( u1_u1_X_13 ) , .ZN( u1_u1_u2_n174 ) );
  INV_X1 u1_u1_u2_U84 (.A( u1_u1_X_18 ) , .ZN( u1_u1_u2_n165 ) );
  NAND4_X1 u1_u1_u2_U85 (.ZN( u1_out1_30 ) , .A4( u1_u1_u2_n147 ) , .A3( u1_u1_u2_n148 ) , .A2( u1_u1_u2_n149 ) , .A1( u1_u1_u2_n187 ) );
  NOR3_X1 u1_u1_u2_U86 (.A3( u1_u1_u2_n144 ) , .A2( u1_u1_u2_n145 ) , .A1( u1_u1_u2_n146 ) , .ZN( u1_u1_u2_n147 ) );
  AOI21_X1 u1_u1_u2_U87 (.B2( u1_u1_u2_n138 ) , .ZN( u1_u1_u2_n148 ) , .A( u1_u1_u2_n162 ) , .B1( u1_u1_u2_n182 ) );
  NAND4_X1 u1_u1_u2_U88 (.ZN( u1_out1_24 ) , .A4( u1_u1_u2_n111 ) , .A3( u1_u1_u2_n112 ) , .A1( u1_u1_u2_n130 ) , .A2( u1_u1_u2_n187 ) );
  AOI221_X1 u1_u1_u2_U89 (.A( u1_u1_u2_n109 ) , .B1( u1_u1_u2_n110 ) , .ZN( u1_u1_u2_n111 ) , .C1( u1_u1_u2_n134 ) , .C2( u1_u1_u2_n170 ) , .B2( u1_u1_u2_n173 ) );
  AOI21_X1 u1_u1_u2_U9 (.B2( u1_u1_u2_n123 ) , .ZN( u1_u1_u2_n125 ) , .A( u1_u1_u2_n171 ) , .B1( u1_u1_u2_n184 ) );
  AOI21_X1 u1_u1_u2_U90 (.ZN( u1_u1_u2_n112 ) , .B2( u1_u1_u2_n156 ) , .A( u1_u1_u2_n164 ) , .B1( u1_u1_u2_n181 ) );
  NAND4_X1 u1_u1_u2_U91 (.ZN( u1_out1_16 ) , .A4( u1_u1_u2_n128 ) , .A3( u1_u1_u2_n129 ) , .A1( u1_u1_u2_n130 ) , .A2( u1_u1_u2_n186 ) );
  AOI22_X1 u1_u1_u2_U92 (.A2( u1_u1_u2_n118 ) , .ZN( u1_u1_u2_n129 ) , .A1( u1_u1_u2_n140 ) , .B1( u1_u1_u2_n157 ) , .B2( u1_u1_u2_n170 ) );
  INV_X1 u1_u1_u2_U93 (.A( u1_u1_u2_n163 ) , .ZN( u1_u1_u2_n186 ) );
  OR4_X1 u1_u1_u2_U94 (.ZN( u1_out1_6 ) , .A4( u1_u1_u2_n161 ) , .A3( u1_u1_u2_n162 ) , .A2( u1_u1_u2_n163 ) , .A1( u1_u1_u2_n164 ) );
  OR3_X1 u1_u1_u2_U95 (.A2( u1_u1_u2_n159 ) , .A1( u1_u1_u2_n160 ) , .ZN( u1_u1_u2_n161 ) , .A3( u1_u1_u2_n183 ) );
  AOI21_X1 u1_u1_u2_U96 (.B2( u1_u1_u2_n154 ) , .B1( u1_u1_u2_n155 ) , .ZN( u1_u1_u2_n159 ) , .A( u1_u1_u2_n167 ) );
  NAND3_X1 u1_u1_u2_U97 (.A2( u1_u1_u2_n117 ) , .A1( u1_u1_u2_n122 ) , .A3( u1_u1_u2_n123 ) , .ZN( u1_u1_u2_n134 ) );
  NAND3_X1 u1_u1_u2_U98 (.ZN( u1_u1_u2_n110 ) , .A2( u1_u1_u2_n131 ) , .A3( u1_u1_u2_n139 ) , .A1( u1_u1_u2_n154 ) );
  NAND3_X1 u1_u1_u2_U99 (.A2( u1_u1_u2_n100 ) , .ZN( u1_u1_u2_n101 ) , .A1( u1_u1_u2_n104 ) , .A3( u1_u1_u2_n114 ) );
  OAI22_X1 u1_u1_u3_U10 (.B1( u1_u1_u3_n113 ) , .A2( u1_u1_u3_n135 ) , .A1( u1_u1_u3_n150 ) , .B2( u1_u1_u3_n164 ) , .ZN( u1_u1_u3_n98 ) );
  OAI211_X1 u1_u1_u3_U11 (.B( u1_u1_u3_n106 ) , .ZN( u1_u1_u3_n119 ) , .C2( u1_u1_u3_n128 ) , .C1( u1_u1_u3_n167 ) , .A( u1_u1_u3_n181 ) );
  AOI221_X1 u1_u1_u3_U12 (.C1( u1_u1_u3_n105 ) , .ZN( u1_u1_u3_n106 ) , .A( u1_u1_u3_n131 ) , .B2( u1_u1_u3_n132 ) , .C2( u1_u1_u3_n133 ) , .B1( u1_u1_u3_n169 ) );
  INV_X1 u1_u1_u3_U13 (.ZN( u1_u1_u3_n181 ) , .A( u1_u1_u3_n98 ) );
  NAND2_X1 u1_u1_u3_U14 (.ZN( u1_u1_u3_n105 ) , .A2( u1_u1_u3_n130 ) , .A1( u1_u1_u3_n155 ) );
  AOI22_X1 u1_u1_u3_U15 (.B1( u1_u1_u3_n115 ) , .A2( u1_u1_u3_n116 ) , .ZN( u1_u1_u3_n123 ) , .B2( u1_u1_u3_n133 ) , .A1( u1_u1_u3_n169 ) );
  NAND2_X1 u1_u1_u3_U16 (.ZN( u1_u1_u3_n116 ) , .A2( u1_u1_u3_n151 ) , .A1( u1_u1_u3_n182 ) );
  NOR2_X1 u1_u1_u3_U17 (.ZN( u1_u1_u3_n126 ) , .A2( u1_u1_u3_n150 ) , .A1( u1_u1_u3_n164 ) );
  AOI21_X1 u1_u1_u3_U18 (.ZN( u1_u1_u3_n112 ) , .B2( u1_u1_u3_n146 ) , .B1( u1_u1_u3_n155 ) , .A( u1_u1_u3_n167 ) );
  NAND2_X1 u1_u1_u3_U19 (.A1( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n142 ) , .A2( u1_u1_u3_n164 ) );
  NAND2_X1 u1_u1_u3_U20 (.ZN( u1_u1_u3_n132 ) , .A2( u1_u1_u3_n152 ) , .A1( u1_u1_u3_n156 ) );
  AND2_X1 u1_u1_u3_U21 (.A2( u1_u1_u3_n113 ) , .A1( u1_u1_u3_n114 ) , .ZN( u1_u1_u3_n151 ) );
  INV_X1 u1_u1_u3_U22 (.A( u1_u1_u3_n133 ) , .ZN( u1_u1_u3_n165 ) );
  INV_X1 u1_u1_u3_U23 (.A( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n170 ) );
  NAND2_X1 u1_u1_u3_U24 (.A1( u1_u1_u3_n107 ) , .A2( u1_u1_u3_n108 ) , .ZN( u1_u1_u3_n140 ) );
  NAND2_X1 u1_u1_u3_U25 (.ZN( u1_u1_u3_n117 ) , .A1( u1_u1_u3_n124 ) , .A2( u1_u1_u3_n148 ) );
  NAND2_X1 u1_u1_u3_U26 (.ZN( u1_u1_u3_n143 ) , .A1( u1_u1_u3_n165 ) , .A2( u1_u1_u3_n167 ) );
  INV_X1 u1_u1_u3_U27 (.A( u1_u1_u3_n130 ) , .ZN( u1_u1_u3_n177 ) );
  INV_X1 u1_u1_u3_U28 (.A( u1_u1_u3_n128 ) , .ZN( u1_u1_u3_n176 ) );
  INV_X1 u1_u1_u3_U29 (.A( u1_u1_u3_n155 ) , .ZN( u1_u1_u3_n174 ) );
  INV_X1 u1_u1_u3_U3 (.A( u1_u1_u3_n129 ) , .ZN( u1_u1_u3_n183 ) );
  INV_X1 u1_u1_u3_U30 (.A( u1_u1_u3_n139 ) , .ZN( u1_u1_u3_n185 ) );
  NOR2_X1 u1_u1_u3_U31 (.ZN( u1_u1_u3_n135 ) , .A2( u1_u1_u3_n141 ) , .A1( u1_u1_u3_n169 ) );
  OAI222_X1 u1_u1_u3_U32 (.C2( u1_u1_u3_n107 ) , .A2( u1_u1_u3_n108 ) , .B1( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n138 ) , .B2( u1_u1_u3_n146 ) , .C1( u1_u1_u3_n154 ) , .A1( u1_u1_u3_n164 ) );
  NOR4_X1 u1_u1_u3_U33 (.A4( u1_u1_u3_n157 ) , .A3( u1_u1_u3_n158 ) , .A2( u1_u1_u3_n159 ) , .A1( u1_u1_u3_n160 ) , .ZN( u1_u1_u3_n161 ) );
  AOI21_X1 u1_u1_u3_U34 (.B2( u1_u1_u3_n152 ) , .B1( u1_u1_u3_n153 ) , .ZN( u1_u1_u3_n158 ) , .A( u1_u1_u3_n164 ) );
  AOI21_X1 u1_u1_u3_U35 (.A( u1_u1_u3_n154 ) , .B2( u1_u1_u3_n155 ) , .B1( u1_u1_u3_n156 ) , .ZN( u1_u1_u3_n157 ) );
  AOI21_X1 u1_u1_u3_U36 (.A( u1_u1_u3_n149 ) , .B2( u1_u1_u3_n150 ) , .B1( u1_u1_u3_n151 ) , .ZN( u1_u1_u3_n159 ) );
  AOI211_X1 u1_u1_u3_U37 (.ZN( u1_u1_u3_n109 ) , .A( u1_u1_u3_n119 ) , .C2( u1_u1_u3_n129 ) , .B( u1_u1_u3_n138 ) , .C1( u1_u1_u3_n141 ) );
  AOI211_X1 u1_u1_u3_U38 (.B( u1_u1_u3_n119 ) , .A( u1_u1_u3_n120 ) , .C2( u1_u1_u3_n121 ) , .ZN( u1_u1_u3_n122 ) , .C1( u1_u1_u3_n179 ) );
  INV_X1 u1_u1_u3_U39 (.A( u1_u1_u3_n156 ) , .ZN( u1_u1_u3_n179 ) );
  INV_X1 u1_u1_u3_U4 (.A( u1_u1_u3_n140 ) , .ZN( u1_u1_u3_n182 ) );
  OAI22_X1 u1_u1_u3_U40 (.B1( u1_u1_u3_n118 ) , .ZN( u1_u1_u3_n120 ) , .A1( u1_u1_u3_n135 ) , .B2( u1_u1_u3_n154 ) , .A2( u1_u1_u3_n178 ) );
  AND3_X1 u1_u1_u3_U41 (.ZN( u1_u1_u3_n118 ) , .A2( u1_u1_u3_n124 ) , .A1( u1_u1_u3_n144 ) , .A3( u1_u1_u3_n152 ) );
  INV_X1 u1_u1_u3_U42 (.A( u1_u1_u3_n121 ) , .ZN( u1_u1_u3_n164 ) );
  NAND2_X1 u1_u1_u3_U43 (.ZN( u1_u1_u3_n133 ) , .A1( u1_u1_u3_n154 ) , .A2( u1_u1_u3_n164 ) );
  OAI211_X1 u1_u1_u3_U44 (.B( u1_u1_u3_n127 ) , .ZN( u1_u1_u3_n139 ) , .C1( u1_u1_u3_n150 ) , .C2( u1_u1_u3_n154 ) , .A( u1_u1_u3_n184 ) );
  INV_X1 u1_u1_u3_U45 (.A( u1_u1_u3_n125 ) , .ZN( u1_u1_u3_n184 ) );
  AOI221_X1 u1_u1_u3_U46 (.A( u1_u1_u3_n126 ) , .ZN( u1_u1_u3_n127 ) , .C2( u1_u1_u3_n132 ) , .C1( u1_u1_u3_n169 ) , .B2( u1_u1_u3_n170 ) , .B1( u1_u1_u3_n174 ) );
  OAI22_X1 u1_u1_u3_U47 (.A1( u1_u1_u3_n124 ) , .ZN( u1_u1_u3_n125 ) , .B2( u1_u1_u3_n145 ) , .A2( u1_u1_u3_n165 ) , .B1( u1_u1_u3_n167 ) );
  NOR2_X1 u1_u1_u3_U48 (.A1( u1_u1_u3_n113 ) , .ZN( u1_u1_u3_n131 ) , .A2( u1_u1_u3_n154 ) );
  NAND2_X1 u1_u1_u3_U49 (.A1( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n150 ) , .A2( u1_u1_u3_n99 ) );
  INV_X1 u1_u1_u3_U5 (.A( u1_u1_u3_n117 ) , .ZN( u1_u1_u3_n178 ) );
  NAND2_X1 u1_u1_u3_U50 (.A2( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n155 ) , .A1( u1_u1_u3_n97 ) );
  INV_X1 u1_u1_u3_U51 (.A( u1_u1_u3_n141 ) , .ZN( u1_u1_u3_n167 ) );
  AOI21_X1 u1_u1_u3_U52 (.B2( u1_u1_u3_n114 ) , .B1( u1_u1_u3_n146 ) , .A( u1_u1_u3_n154 ) , .ZN( u1_u1_u3_n94 ) );
  AOI21_X1 u1_u1_u3_U53 (.ZN( u1_u1_u3_n110 ) , .B2( u1_u1_u3_n142 ) , .B1( u1_u1_u3_n186 ) , .A( u1_u1_u3_n95 ) );
  INV_X1 u1_u1_u3_U54 (.A( u1_u1_u3_n145 ) , .ZN( u1_u1_u3_n186 ) );
  AOI21_X1 u1_u1_u3_U55 (.B1( u1_u1_u3_n124 ) , .A( u1_u1_u3_n149 ) , .B2( u1_u1_u3_n155 ) , .ZN( u1_u1_u3_n95 ) );
  INV_X1 u1_u1_u3_U56 (.A( u1_u1_u3_n149 ) , .ZN( u1_u1_u3_n169 ) );
  NAND2_X1 u1_u1_u3_U57 (.ZN( u1_u1_u3_n124 ) , .A1( u1_u1_u3_n96 ) , .A2( u1_u1_u3_n97 ) );
  NAND2_X1 u1_u1_u3_U58 (.A2( u1_u1_u3_n100 ) , .ZN( u1_u1_u3_n146 ) , .A1( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U59 (.A1( u1_u1_u3_n101 ) , .ZN( u1_u1_u3_n145 ) , .A2( u1_u1_u3_n99 ) );
  AOI221_X1 u1_u1_u3_U6 (.A( u1_u1_u3_n131 ) , .C2( u1_u1_u3_n132 ) , .C1( u1_u1_u3_n133 ) , .ZN( u1_u1_u3_n134 ) , .B1( u1_u1_u3_n143 ) , .B2( u1_u1_u3_n177 ) );
  NAND2_X1 u1_u1_u3_U60 (.A1( u1_u1_u3_n100 ) , .ZN( u1_u1_u3_n156 ) , .A2( u1_u1_u3_n99 ) );
  NAND2_X1 u1_u1_u3_U61 (.A2( u1_u1_u3_n101 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n148 ) );
  NAND2_X1 u1_u1_u3_U62 (.A1( u1_u1_u3_n100 ) , .A2( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n128 ) );
  NAND2_X1 u1_u1_u3_U63 (.A2( u1_u1_u3_n101 ) , .A1( u1_u1_u3_n102 ) , .ZN( u1_u1_u3_n152 ) );
  NAND2_X1 u1_u1_u3_U64 (.A2( u1_u1_u3_n101 ) , .ZN( u1_u1_u3_n114 ) , .A1( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U65 (.ZN( u1_u1_u3_n107 ) , .A1( u1_u1_u3_n97 ) , .A2( u1_u1_u3_n99 ) );
  NAND2_X1 u1_u1_u3_U66 (.A2( u1_u1_u3_n100 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n113 ) );
  NAND2_X1 u1_u1_u3_U67 (.A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n153 ) , .A2( u1_u1_u3_n97 ) );
  NAND2_X1 u1_u1_u3_U68 (.A2( u1_u1_u3_n103 ) , .A1( u1_u1_u3_n104 ) , .ZN( u1_u1_u3_n130 ) );
  NAND2_X1 u1_u1_u3_U69 (.A2( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n144 ) , .A1( u1_u1_u3_n96 ) );
  OAI22_X1 u1_u1_u3_U7 (.B2( u1_u1_u3_n147 ) , .A2( u1_u1_u3_n148 ) , .ZN( u1_u1_u3_n160 ) , .B1( u1_u1_u3_n165 ) , .A1( u1_u1_u3_n168 ) );
  NAND2_X1 u1_u1_u3_U70 (.A1( u1_u1_u3_n102 ) , .A2( u1_u1_u3_n103 ) , .ZN( u1_u1_u3_n108 ) );
  NOR2_X1 u1_u1_u3_U71 (.A2( u1_u1_X_19 ) , .A1( u1_u1_X_20 ) , .ZN( u1_u1_u3_n99 ) );
  NOR2_X1 u1_u1_u3_U72 (.A2( u1_u1_X_21 ) , .A1( u1_u1_X_24 ) , .ZN( u1_u1_u3_n103 ) );
  NOR2_X1 u1_u1_u3_U73 (.A2( u1_u1_X_24 ) , .A1( u1_u1_u3_n171 ) , .ZN( u1_u1_u3_n97 ) );
  NOR2_X1 u1_u1_u3_U74 (.A2( u1_u1_X_23 ) , .ZN( u1_u1_u3_n141 ) , .A1( u1_u1_u3_n166 ) );
  NOR2_X1 u1_u1_u3_U75 (.A2( u1_u1_X_19 ) , .A1( u1_u1_u3_n172 ) , .ZN( u1_u1_u3_n96 ) );
  NAND2_X1 u1_u1_u3_U76 (.A1( u1_u1_X_22 ) , .A2( u1_u1_X_23 ) , .ZN( u1_u1_u3_n154 ) );
  NAND2_X1 u1_u1_u3_U77 (.A1( u1_u1_X_23 ) , .ZN( u1_u1_u3_n149 ) , .A2( u1_u1_u3_n166 ) );
  NOR2_X1 u1_u1_u3_U78 (.A2( u1_u1_X_22 ) , .A1( u1_u1_X_23 ) , .ZN( u1_u1_u3_n121 ) );
  AND2_X1 u1_u1_u3_U79 (.A1( u1_u1_X_24 ) , .ZN( u1_u1_u3_n101 ) , .A2( u1_u1_u3_n171 ) );
  AND3_X1 u1_u1_u3_U8 (.A3( u1_u1_u3_n144 ) , .A2( u1_u1_u3_n145 ) , .A1( u1_u1_u3_n146 ) , .ZN( u1_u1_u3_n147 ) );
  AND2_X1 u1_u1_u3_U80 (.A1( u1_u1_X_19 ) , .ZN( u1_u1_u3_n102 ) , .A2( u1_u1_u3_n172 ) );
  AND2_X1 u1_u1_u3_U81 (.A1( u1_u1_X_21 ) , .A2( u1_u1_X_24 ) , .ZN( u1_u1_u3_n100 ) );
  AND2_X1 u1_u1_u3_U82 (.A2( u1_u1_X_19 ) , .A1( u1_u1_X_20 ) , .ZN( u1_u1_u3_n104 ) );
  INV_X1 u1_u1_u3_U83 (.A( u1_u1_X_22 ) , .ZN( u1_u1_u3_n166 ) );
  INV_X1 u1_u1_u3_U84 (.A( u1_u1_X_21 ) , .ZN( u1_u1_u3_n171 ) );
  INV_X1 u1_u1_u3_U85 (.A( u1_u1_X_20 ) , .ZN( u1_u1_u3_n172 ) );
  OR4_X1 u1_u1_u3_U86 (.ZN( u1_out1_10 ) , .A4( u1_u1_u3_n136 ) , .A3( u1_u1_u3_n137 ) , .A1( u1_u1_u3_n138 ) , .A2( u1_u1_u3_n139 ) );
  OAI222_X1 u1_u1_u3_U87 (.C1( u1_u1_u3_n128 ) , .ZN( u1_u1_u3_n137 ) , .B1( u1_u1_u3_n148 ) , .A2( u1_u1_u3_n150 ) , .B2( u1_u1_u3_n154 ) , .C2( u1_u1_u3_n164 ) , .A1( u1_u1_u3_n167 ) );
  OAI221_X1 u1_u1_u3_U88 (.A( u1_u1_u3_n134 ) , .B2( u1_u1_u3_n135 ) , .ZN( u1_u1_u3_n136 ) , .C1( u1_u1_u3_n149 ) , .B1( u1_u1_u3_n151 ) , .C2( u1_u1_u3_n183 ) );
  NAND4_X1 u1_u1_u3_U89 (.ZN( u1_out1_26 ) , .A4( u1_u1_u3_n109 ) , .A3( u1_u1_u3_n110 ) , .A2( u1_u1_u3_n111 ) , .A1( u1_u1_u3_n173 ) );
  INV_X1 u1_u1_u3_U9 (.A( u1_u1_u3_n143 ) , .ZN( u1_u1_u3_n168 ) );
  INV_X1 u1_u1_u3_U90 (.ZN( u1_u1_u3_n173 ) , .A( u1_u1_u3_n94 ) );
  OAI21_X1 u1_u1_u3_U91 (.ZN( u1_u1_u3_n111 ) , .B2( u1_u1_u3_n117 ) , .A( u1_u1_u3_n133 ) , .B1( u1_u1_u3_n176 ) );
  NAND4_X1 u1_u1_u3_U92 (.ZN( u1_out1_20 ) , .A4( u1_u1_u3_n122 ) , .A3( u1_u1_u3_n123 ) , .A1( u1_u1_u3_n175 ) , .A2( u1_u1_u3_n180 ) );
  INV_X1 u1_u1_u3_U93 (.A( u1_u1_u3_n112 ) , .ZN( u1_u1_u3_n175 ) );
  INV_X1 u1_u1_u3_U94 (.A( u1_u1_u3_n126 ) , .ZN( u1_u1_u3_n180 ) );
  NAND4_X1 u1_u1_u3_U95 (.ZN( u1_out1_1 ) , .A4( u1_u1_u3_n161 ) , .A3( u1_u1_u3_n162 ) , .A2( u1_u1_u3_n163 ) , .A1( u1_u1_u3_n185 ) );
  NAND2_X1 u1_u1_u3_U96 (.ZN( u1_u1_u3_n163 ) , .A2( u1_u1_u3_n170 ) , .A1( u1_u1_u3_n176 ) );
  AOI22_X1 u1_u1_u3_U97 (.B2( u1_u1_u3_n140 ) , .B1( u1_u1_u3_n141 ) , .A2( u1_u1_u3_n142 ) , .ZN( u1_u1_u3_n162 ) , .A1( u1_u1_u3_n177 ) );
  NAND3_X1 u1_u1_u3_U98 (.A1( u1_u1_u3_n114 ) , .ZN( u1_u1_u3_n115 ) , .A2( u1_u1_u3_n145 ) , .A3( u1_u1_u3_n153 ) );
  NAND3_X1 u1_u1_u3_U99 (.ZN( u1_u1_u3_n129 ) , .A2( u1_u1_u3_n144 ) , .A1( u1_u1_u3_n153 ) , .A3( u1_u1_u3_n182 ) );
  OAI22_X1 u1_u1_u4_U10 (.B2( u1_u1_u4_n135 ) , .ZN( u1_u1_u4_n137 ) , .B1( u1_u1_u4_n153 ) , .A1( u1_u1_u4_n155 ) , .A2( u1_u1_u4_n171 ) );
  AND3_X1 u1_u1_u4_U11 (.A2( u1_u1_u4_n134 ) , .ZN( u1_u1_u4_n135 ) , .A3( u1_u1_u4_n145 ) , .A1( u1_u1_u4_n157 ) );
  NAND2_X1 u1_u1_u4_U12 (.ZN( u1_u1_u4_n132 ) , .A2( u1_u1_u4_n170 ) , .A1( u1_u1_u4_n173 ) );
  AOI21_X1 u1_u1_u4_U13 (.B2( u1_u1_u4_n160 ) , .B1( u1_u1_u4_n161 ) , .ZN( u1_u1_u4_n162 ) , .A( u1_u1_u4_n170 ) );
  AOI21_X1 u1_u1_u4_U14 (.ZN( u1_u1_u4_n107 ) , .B2( u1_u1_u4_n143 ) , .A( u1_u1_u4_n174 ) , .B1( u1_u1_u4_n184 ) );
  AOI21_X1 u1_u1_u4_U15 (.B2( u1_u1_u4_n158 ) , .B1( u1_u1_u4_n159 ) , .ZN( u1_u1_u4_n163 ) , .A( u1_u1_u4_n174 ) );
  AOI21_X1 u1_u1_u4_U16 (.A( u1_u1_u4_n153 ) , .B2( u1_u1_u4_n154 ) , .B1( u1_u1_u4_n155 ) , .ZN( u1_u1_u4_n165 ) );
  AOI21_X1 u1_u1_u4_U17 (.A( u1_u1_u4_n156 ) , .B2( u1_u1_u4_n157 ) , .ZN( u1_u1_u4_n164 ) , .B1( u1_u1_u4_n184 ) );
  INV_X1 u1_u1_u4_U18 (.A( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n170 ) );
  AND2_X1 u1_u1_u4_U19 (.A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n155 ) , .A1( u1_u1_u4_n160 ) );
  INV_X1 u1_u1_u4_U20 (.A( u1_u1_u4_n156 ) , .ZN( u1_u1_u4_n175 ) );
  NAND2_X1 u1_u1_u4_U21 (.A2( u1_u1_u4_n118 ) , .ZN( u1_u1_u4_n131 ) , .A1( u1_u1_u4_n147 ) );
  NAND2_X1 u1_u1_u4_U22 (.A1( u1_u1_u4_n119 ) , .A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n130 ) );
  NAND2_X1 u1_u1_u4_U23 (.ZN( u1_u1_u4_n117 ) , .A2( u1_u1_u4_n118 ) , .A1( u1_u1_u4_n148 ) );
  NAND2_X1 u1_u1_u4_U24 (.ZN( u1_u1_u4_n129 ) , .A1( u1_u1_u4_n134 ) , .A2( u1_u1_u4_n148 ) );
  AND3_X1 u1_u1_u4_U25 (.A1( u1_u1_u4_n119 ) , .A2( u1_u1_u4_n143 ) , .A3( u1_u1_u4_n154 ) , .ZN( u1_u1_u4_n161 ) );
  AND2_X1 u1_u1_u4_U26 (.A1( u1_u1_u4_n145 ) , .A2( u1_u1_u4_n147 ) , .ZN( u1_u1_u4_n159 ) );
  OR3_X1 u1_u1_u4_U27 (.A3( u1_u1_u4_n114 ) , .A2( u1_u1_u4_n115 ) , .A1( u1_u1_u4_n116 ) , .ZN( u1_u1_u4_n136 ) );
  AOI21_X1 u1_u1_u4_U28 (.A( u1_u1_u4_n113 ) , .ZN( u1_u1_u4_n116 ) , .B2( u1_u1_u4_n173 ) , .B1( u1_u1_u4_n174 ) );
  AOI21_X1 u1_u1_u4_U29 (.ZN( u1_u1_u4_n115 ) , .B2( u1_u1_u4_n145 ) , .B1( u1_u1_u4_n146 ) , .A( u1_u1_u4_n156 ) );
  NOR2_X1 u1_u1_u4_U3 (.ZN( u1_u1_u4_n121 ) , .A1( u1_u1_u4_n181 ) , .A2( u1_u1_u4_n182 ) );
  OAI22_X1 u1_u1_u4_U30 (.ZN( u1_u1_u4_n114 ) , .A2( u1_u1_u4_n121 ) , .B1( u1_u1_u4_n160 ) , .B2( u1_u1_u4_n170 ) , .A1( u1_u1_u4_n171 ) );
  INV_X1 u1_u1_u4_U31 (.A( u1_u1_u4_n158 ) , .ZN( u1_u1_u4_n182 ) );
  INV_X1 u1_u1_u4_U32 (.ZN( u1_u1_u4_n181 ) , .A( u1_u1_u4_n96 ) );
  INV_X1 u1_u1_u4_U33 (.A( u1_u1_u4_n144 ) , .ZN( u1_u1_u4_n179 ) );
  INV_X1 u1_u1_u4_U34 (.A( u1_u1_u4_n157 ) , .ZN( u1_u1_u4_n178 ) );
  NAND2_X1 u1_u1_u4_U35 (.A2( u1_u1_u4_n154 ) , .A1( u1_u1_u4_n96 ) , .ZN( u1_u1_u4_n97 ) );
  INV_X1 u1_u1_u4_U36 (.ZN( u1_u1_u4_n186 ) , .A( u1_u1_u4_n95 ) );
  OAI221_X1 u1_u1_u4_U37 (.C1( u1_u1_u4_n134 ) , .B1( u1_u1_u4_n158 ) , .B2( u1_u1_u4_n171 ) , .C2( u1_u1_u4_n173 ) , .A( u1_u1_u4_n94 ) , .ZN( u1_u1_u4_n95 ) );
  AOI222_X1 u1_u1_u4_U38 (.B2( u1_u1_u4_n132 ) , .A1( u1_u1_u4_n138 ) , .C2( u1_u1_u4_n175 ) , .A2( u1_u1_u4_n179 ) , .C1( u1_u1_u4_n181 ) , .B1( u1_u1_u4_n185 ) , .ZN( u1_u1_u4_n94 ) );
  INV_X1 u1_u1_u4_U39 (.A( u1_u1_u4_n113 ) , .ZN( u1_u1_u4_n185 ) );
  INV_X1 u1_u1_u4_U4 (.A( u1_u1_u4_n117 ) , .ZN( u1_u1_u4_n184 ) );
  INV_X1 u1_u1_u4_U40 (.A( u1_u1_u4_n143 ) , .ZN( u1_u1_u4_n183 ) );
  NOR2_X1 u1_u1_u4_U41 (.ZN( u1_u1_u4_n138 ) , .A1( u1_u1_u4_n168 ) , .A2( u1_u1_u4_n169 ) );
  NOR2_X1 u1_u1_u4_U42 (.A1( u1_u1_u4_n150 ) , .A2( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n153 ) );
  NOR2_X1 u1_u1_u4_U43 (.A2( u1_u1_u4_n128 ) , .A1( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n156 ) );
  AOI22_X1 u1_u1_u4_U44 (.B2( u1_u1_u4_n122 ) , .A1( u1_u1_u4_n123 ) , .ZN( u1_u1_u4_n124 ) , .B1( u1_u1_u4_n128 ) , .A2( u1_u1_u4_n172 ) );
  NAND2_X1 u1_u1_u4_U45 (.A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n123 ) , .A1( u1_u1_u4_n161 ) );
  INV_X1 u1_u1_u4_U46 (.A( u1_u1_u4_n153 ) , .ZN( u1_u1_u4_n172 ) );
  AOI22_X1 u1_u1_u4_U47 (.B2( u1_u1_u4_n132 ) , .A2( u1_u1_u4_n133 ) , .ZN( u1_u1_u4_n140 ) , .A1( u1_u1_u4_n150 ) , .B1( u1_u1_u4_n179 ) );
  NAND2_X1 u1_u1_u4_U48 (.ZN( u1_u1_u4_n133 ) , .A2( u1_u1_u4_n146 ) , .A1( u1_u1_u4_n154 ) );
  NAND2_X1 u1_u1_u4_U49 (.A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n154 ) , .A2( u1_u1_u4_n98 ) );
  NOR4_X1 u1_u1_u4_U5 (.A4( u1_u1_u4_n106 ) , .A3( u1_u1_u4_n107 ) , .A2( u1_u1_u4_n108 ) , .A1( u1_u1_u4_n109 ) , .ZN( u1_u1_u4_n110 ) );
  NAND2_X1 u1_u1_u4_U50 (.A1( u1_u1_u4_n101 ) , .ZN( u1_u1_u4_n158 ) , .A2( u1_u1_u4_n99 ) );
  AOI21_X1 u1_u1_u4_U51 (.ZN( u1_u1_u4_n127 ) , .A( u1_u1_u4_n136 ) , .B2( u1_u1_u4_n150 ) , .B1( u1_u1_u4_n180 ) );
  INV_X1 u1_u1_u4_U52 (.A( u1_u1_u4_n160 ) , .ZN( u1_u1_u4_n180 ) );
  NAND2_X1 u1_u1_u4_U53 (.A2( u1_u1_u4_n104 ) , .A1( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n146 ) );
  NAND2_X1 u1_u1_u4_U54 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n160 ) );
  NAND2_X1 u1_u1_u4_U55 (.ZN( u1_u1_u4_n134 ) , .A1( u1_u1_u4_n98 ) , .A2( u1_u1_u4_n99 ) );
  NAND2_X1 u1_u1_u4_U56 (.A1( u1_u1_u4_n103 ) , .A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n143 ) );
  NAND2_X1 u1_u1_u4_U57 (.A2( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n145 ) , .A1( u1_u1_u4_n98 ) );
  NAND2_X1 u1_u1_u4_U58 (.A1( u1_u1_u4_n100 ) , .A2( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n120 ) );
  NAND2_X1 u1_u1_u4_U59 (.A1( u1_u1_u4_n102 ) , .A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n148 ) );
  AOI21_X1 u1_u1_u4_U6 (.ZN( u1_u1_u4_n106 ) , .B2( u1_u1_u4_n146 ) , .B1( u1_u1_u4_n158 ) , .A( u1_u1_u4_n170 ) );
  NAND2_X1 u1_u1_u4_U60 (.A2( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n157 ) );
  INV_X1 u1_u1_u4_U61 (.A( u1_u1_u4_n150 ) , .ZN( u1_u1_u4_n173 ) );
  INV_X1 u1_u1_u4_U62 (.A( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n171 ) );
  NAND2_X1 u1_u1_u4_U63 (.A1( u1_u1_u4_n100 ) , .ZN( u1_u1_u4_n118 ) , .A2( u1_u1_u4_n99 ) );
  NAND2_X1 u1_u1_u4_U64 (.A2( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n144 ) );
  NAND2_X1 u1_u1_u4_U65 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n96 ) );
  INV_X1 u1_u1_u4_U66 (.A( u1_u1_u4_n128 ) , .ZN( u1_u1_u4_n174 ) );
  NAND2_X1 u1_u1_u4_U67 (.A2( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n119 ) , .A1( u1_u1_u4_n98 ) );
  NAND2_X1 u1_u1_u4_U68 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n147 ) );
  NAND2_X1 u1_u1_u4_U69 (.A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n113 ) , .A1( u1_u1_u4_n99 ) );
  AOI21_X1 u1_u1_u4_U7 (.ZN( u1_u1_u4_n108 ) , .B2( u1_u1_u4_n134 ) , .B1( u1_u1_u4_n155 ) , .A( u1_u1_u4_n156 ) );
  NOR2_X1 u1_u1_u4_U70 (.A2( u1_u1_X_28 ) , .ZN( u1_u1_u4_n150 ) , .A1( u1_u1_u4_n168 ) );
  NOR2_X1 u1_u1_u4_U71 (.A2( u1_u1_X_29 ) , .ZN( u1_u1_u4_n152 ) , .A1( u1_u1_u4_n169 ) );
  NOR2_X1 u1_u1_u4_U72 (.A2( u1_u1_X_30 ) , .ZN( u1_u1_u4_n105 ) , .A1( u1_u1_u4_n176 ) );
  NOR2_X1 u1_u1_u4_U73 (.A2( u1_u1_X_26 ) , .ZN( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n177 ) );
  NOR2_X1 u1_u1_u4_U74 (.A2( u1_u1_X_28 ) , .A1( u1_u1_X_29 ) , .ZN( u1_u1_u4_n128 ) );
  NOR2_X1 u1_u1_u4_U75 (.A2( u1_u1_X_27 ) , .A1( u1_u1_X_30 ) , .ZN( u1_u1_u4_n102 ) );
  NOR2_X1 u1_u1_u4_U76 (.A2( u1_u1_X_25 ) , .A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n98 ) );
  AND2_X1 u1_u1_u4_U77 (.A2( u1_u1_X_25 ) , .A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n104 ) );
  AND2_X1 u1_u1_u4_U78 (.A1( u1_u1_X_30 ) , .A2( u1_u1_u4_n176 ) , .ZN( u1_u1_u4_n99 ) );
  AND2_X1 u1_u1_u4_U79 (.A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n101 ) , .A2( u1_u1_u4_n177 ) );
  AOI21_X1 u1_u1_u4_U8 (.ZN( u1_u1_u4_n109 ) , .A( u1_u1_u4_n153 ) , .B1( u1_u1_u4_n159 ) , .B2( u1_u1_u4_n184 ) );
  AND2_X1 u1_u1_u4_U80 (.A1( u1_u1_X_27 ) , .A2( u1_u1_X_30 ) , .ZN( u1_u1_u4_n103 ) );
  INV_X1 u1_u1_u4_U81 (.A( u1_u1_X_28 ) , .ZN( u1_u1_u4_n169 ) );
  INV_X1 u1_u1_u4_U82 (.A( u1_u1_X_29 ) , .ZN( u1_u1_u4_n168 ) );
  INV_X1 u1_u1_u4_U83 (.A( u1_u1_X_25 ) , .ZN( u1_u1_u4_n177 ) );
  INV_X1 u1_u1_u4_U84 (.A( u1_u1_X_27 ) , .ZN( u1_u1_u4_n176 ) );
  NAND4_X1 u1_u1_u4_U85 (.ZN( u1_out1_25 ) , .A4( u1_u1_u4_n139 ) , .A3( u1_u1_u4_n140 ) , .A2( u1_u1_u4_n141 ) , .A1( u1_u1_u4_n142 ) );
  OAI21_X1 u1_u1_u4_U86 (.A( u1_u1_u4_n128 ) , .B2( u1_u1_u4_n129 ) , .B1( u1_u1_u4_n130 ) , .ZN( u1_u1_u4_n142 ) );
  OAI21_X1 u1_u1_u4_U87 (.B2( u1_u1_u4_n131 ) , .ZN( u1_u1_u4_n141 ) , .A( u1_u1_u4_n175 ) , .B1( u1_u1_u4_n183 ) );
  NAND4_X1 u1_u1_u4_U88 (.ZN( u1_out1_14 ) , .A4( u1_u1_u4_n124 ) , .A3( u1_u1_u4_n125 ) , .A2( u1_u1_u4_n126 ) , .A1( u1_u1_u4_n127 ) );
  AOI22_X1 u1_u1_u4_U89 (.B2( u1_u1_u4_n117 ) , .ZN( u1_u1_u4_n126 ) , .A1( u1_u1_u4_n129 ) , .B1( u1_u1_u4_n152 ) , .A2( u1_u1_u4_n175 ) );
  AOI211_X1 u1_u1_u4_U9 (.B( u1_u1_u4_n136 ) , .A( u1_u1_u4_n137 ) , .C2( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n139 ) , .C1( u1_u1_u4_n182 ) );
  AOI22_X1 u1_u1_u4_U90 (.ZN( u1_u1_u4_n125 ) , .B2( u1_u1_u4_n131 ) , .A2( u1_u1_u4_n132 ) , .B1( u1_u1_u4_n138 ) , .A1( u1_u1_u4_n178 ) );
  NAND4_X1 u1_u1_u4_U91 (.ZN( u1_out1_8 ) , .A4( u1_u1_u4_n110 ) , .A3( u1_u1_u4_n111 ) , .A2( u1_u1_u4_n112 ) , .A1( u1_u1_u4_n186 ) );
  NAND2_X1 u1_u1_u4_U92 (.ZN( u1_u1_u4_n112 ) , .A2( u1_u1_u4_n130 ) , .A1( u1_u1_u4_n150 ) );
  AOI22_X1 u1_u1_u4_U93 (.ZN( u1_u1_u4_n111 ) , .B2( u1_u1_u4_n132 ) , .A1( u1_u1_u4_n152 ) , .B1( u1_u1_u4_n178 ) , .A2( u1_u1_u4_n97 ) );
  AOI22_X1 u1_u1_u4_U94 (.B2( u1_u1_u4_n149 ) , .B1( u1_u1_u4_n150 ) , .A2( u1_u1_u4_n151 ) , .A1( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n167 ) );
  NOR4_X1 u1_u1_u4_U95 (.A4( u1_u1_u4_n162 ) , .A3( u1_u1_u4_n163 ) , .A2( u1_u1_u4_n164 ) , .A1( u1_u1_u4_n165 ) , .ZN( u1_u1_u4_n166 ) );
  NAND3_X1 u1_u1_u4_U96 (.ZN( u1_out1_3 ) , .A3( u1_u1_u4_n166 ) , .A1( u1_u1_u4_n167 ) , .A2( u1_u1_u4_n186 ) );
  NAND3_X1 u1_u1_u4_U97 (.A3( u1_u1_u4_n146 ) , .A2( u1_u1_u4_n147 ) , .A1( u1_u1_u4_n148 ) , .ZN( u1_u1_u4_n149 ) );
  NAND3_X1 u1_u1_u4_U98 (.A3( u1_u1_u4_n143 ) , .A2( u1_u1_u4_n144 ) , .A1( u1_u1_u4_n145 ) , .ZN( u1_u1_u4_n151 ) );
  NAND3_X1 u1_u1_u4_U99 (.A3( u1_u1_u4_n121 ) , .ZN( u1_u1_u4_n122 ) , .A2( u1_u1_u4_n144 ) , .A1( u1_u1_u4_n154 ) );
  AOI22_X1 u1_u1_u6_U10 (.A2( u1_u1_u6_n151 ) , .B2( u1_u1_u6_n161 ) , .A1( u1_u1_u6_n167 ) , .B1( u1_u1_u6_n170 ) , .ZN( u1_u1_u6_n89 ) );
  AOI21_X1 u1_u1_u6_U11 (.B1( u1_u1_u6_n107 ) , .B2( u1_u1_u6_n132 ) , .A( u1_u1_u6_n158 ) , .ZN( u1_u1_u6_n88 ) );
  AOI21_X1 u1_u1_u6_U12 (.B2( u1_u1_u6_n147 ) , .B1( u1_u1_u6_n148 ) , .ZN( u1_u1_u6_n149 ) , .A( u1_u1_u6_n158 ) );
  AOI21_X1 u1_u1_u6_U13 (.ZN( u1_u1_u6_n106 ) , .A( u1_u1_u6_n142 ) , .B2( u1_u1_u6_n159 ) , .B1( u1_u1_u6_n164 ) );
  INV_X1 u1_u1_u6_U14 (.A( u1_u1_u6_n155 ) , .ZN( u1_u1_u6_n161 ) );
  INV_X1 u1_u1_u6_U15 (.A( u1_u1_u6_n128 ) , .ZN( u1_u1_u6_n164 ) );
  NAND2_X1 u1_u1_u6_U16 (.ZN( u1_u1_u6_n110 ) , .A1( u1_u1_u6_n122 ) , .A2( u1_u1_u6_n129 ) );
  NAND2_X1 u1_u1_u6_U17 (.ZN( u1_u1_u6_n124 ) , .A2( u1_u1_u6_n146 ) , .A1( u1_u1_u6_n148 ) );
  INV_X1 u1_u1_u6_U18 (.A( u1_u1_u6_n132 ) , .ZN( u1_u1_u6_n171 ) );
  AND2_X1 u1_u1_u6_U19 (.A1( u1_u1_u6_n100 ) , .ZN( u1_u1_u6_n130 ) , .A2( u1_u1_u6_n147 ) );
  INV_X1 u1_u1_u6_U20 (.A( u1_u1_u6_n127 ) , .ZN( u1_u1_u6_n173 ) );
  INV_X1 u1_u1_u6_U21 (.A( u1_u1_u6_n121 ) , .ZN( u1_u1_u6_n167 ) );
  INV_X1 u1_u1_u6_U22 (.A( u1_u1_u6_n100 ) , .ZN( u1_u1_u6_n169 ) );
  INV_X1 u1_u1_u6_U23 (.A( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n170 ) );
  INV_X1 u1_u1_u6_U24 (.A( u1_u1_u6_n113 ) , .ZN( u1_u1_u6_n168 ) );
  AND2_X1 u1_u1_u6_U25 (.A1( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n119 ) , .ZN( u1_u1_u6_n133 ) );
  AND2_X1 u1_u1_u6_U26 (.A2( u1_u1_u6_n121 ) , .A1( u1_u1_u6_n122 ) , .ZN( u1_u1_u6_n131 ) );
  AND3_X1 u1_u1_u6_U27 (.ZN( u1_u1_u6_n120 ) , .A2( u1_u1_u6_n127 ) , .A1( u1_u1_u6_n132 ) , .A3( u1_u1_u6_n145 ) );
  INV_X1 u1_u1_u6_U28 (.A( u1_u1_u6_n146 ) , .ZN( u1_u1_u6_n163 ) );
  AOI222_X1 u1_u1_u6_U29 (.ZN( u1_u1_u6_n114 ) , .A1( u1_u1_u6_n118 ) , .A2( u1_u1_u6_n126 ) , .B2( u1_u1_u6_n151 ) , .C2( u1_u1_u6_n159 ) , .C1( u1_u1_u6_n168 ) , .B1( u1_u1_u6_n169 ) );
  INV_X1 u1_u1_u6_U3 (.A( u1_u1_u6_n110 ) , .ZN( u1_u1_u6_n166 ) );
  NOR2_X1 u1_u1_u6_U30 (.A1( u1_u1_u6_n162 ) , .A2( u1_u1_u6_n165 ) , .ZN( u1_u1_u6_n98 ) );
  AOI211_X1 u1_u1_u6_U31 (.B( u1_u1_u6_n134 ) , .A( u1_u1_u6_n135 ) , .C1( u1_u1_u6_n136 ) , .ZN( u1_u1_u6_n137 ) , .C2( u1_u1_u6_n151 ) );
  AOI21_X1 u1_u1_u6_U32 (.B1( u1_u1_u6_n131 ) , .ZN( u1_u1_u6_n135 ) , .A( u1_u1_u6_n144 ) , .B2( u1_u1_u6_n146 ) );
  NAND4_X1 u1_u1_u6_U33 (.A4( u1_u1_u6_n127 ) , .A3( u1_u1_u6_n128 ) , .A2( u1_u1_u6_n129 ) , .A1( u1_u1_u6_n130 ) , .ZN( u1_u1_u6_n136 ) );
  AOI21_X1 u1_u1_u6_U34 (.B2( u1_u1_u6_n132 ) , .B1( u1_u1_u6_n133 ) , .ZN( u1_u1_u6_n134 ) , .A( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U35 (.A1( u1_u1_u6_n144 ) , .ZN( u1_u1_u6_n151 ) , .A2( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U36 (.ZN( u1_u1_u6_n132 ) , .A1( u1_u1_u6_n91 ) , .A2( u1_u1_u6_n97 ) );
  AOI22_X1 u1_u1_u6_U37 (.B2( u1_u1_u6_n110 ) , .B1( u1_u1_u6_n111 ) , .A1( u1_u1_u6_n112 ) , .ZN( u1_u1_u6_n115 ) , .A2( u1_u1_u6_n161 ) );
  NAND4_X1 u1_u1_u6_U38 (.A3( u1_u1_u6_n109 ) , .ZN( u1_u1_u6_n112 ) , .A4( u1_u1_u6_n132 ) , .A2( u1_u1_u6_n147 ) , .A1( u1_u1_u6_n166 ) );
  NOR2_X1 u1_u1_u6_U39 (.ZN( u1_u1_u6_n109 ) , .A1( u1_u1_u6_n170 ) , .A2( u1_u1_u6_n173 ) );
  INV_X1 u1_u1_u6_U4 (.A( u1_u1_u6_n142 ) , .ZN( u1_u1_u6_n174 ) );
  NOR2_X1 u1_u1_u6_U40 (.A2( u1_u1_u6_n126 ) , .ZN( u1_u1_u6_n155 ) , .A1( u1_u1_u6_n160 ) );
  NAND2_X1 u1_u1_u6_U41 (.ZN( u1_u1_u6_n146 ) , .A2( u1_u1_u6_n94 ) , .A1( u1_u1_u6_n99 ) );
  AOI21_X1 u1_u1_u6_U42 (.A( u1_u1_u6_n144 ) , .B2( u1_u1_u6_n145 ) , .B1( u1_u1_u6_n146 ) , .ZN( u1_u1_u6_n150 ) );
  INV_X1 u1_u1_u6_U43 (.A( u1_u1_u6_n111 ) , .ZN( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U44 (.ZN( u1_u1_u6_n127 ) , .A1( u1_u1_u6_n91 ) , .A2( u1_u1_u6_n92 ) );
  NAND2_X1 u1_u1_u6_U45 (.ZN( u1_u1_u6_n129 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n96 ) );
  INV_X1 u1_u1_u6_U46 (.A( u1_u1_u6_n144 ) , .ZN( u1_u1_u6_n159 ) );
  NAND2_X1 u1_u1_u6_U47 (.ZN( u1_u1_u6_n145 ) , .A2( u1_u1_u6_n97 ) , .A1( u1_u1_u6_n98 ) );
  NAND2_X1 u1_u1_u6_U48 (.ZN( u1_u1_u6_n148 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n94 ) );
  NAND2_X1 u1_u1_u6_U49 (.ZN( u1_u1_u6_n108 ) , .A2( u1_u1_u6_n139 ) , .A1( u1_u1_u6_n144 ) );
  NAND2_X1 u1_u1_u6_U5 (.A2( u1_u1_u6_n143 ) , .ZN( u1_u1_u6_n152 ) , .A1( u1_u1_u6_n166 ) );
  NAND2_X1 u1_u1_u6_U50 (.ZN( u1_u1_u6_n121 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n97 ) );
  NAND2_X1 u1_u1_u6_U51 (.ZN( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n95 ) );
  AND2_X1 u1_u1_u6_U52 (.ZN( u1_u1_u6_n118 ) , .A2( u1_u1_u6_n91 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U53 (.ZN( u1_u1_u6_n147 ) , .A2( u1_u1_u6_n98 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U54 (.ZN( u1_u1_u6_n128 ) , .A1( u1_u1_u6_n94 ) , .A2( u1_u1_u6_n96 ) );
  NAND2_X1 u1_u1_u6_U55 (.ZN( u1_u1_u6_n119 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U56 (.ZN( u1_u1_u6_n123 ) , .A2( u1_u1_u6_n91 ) , .A1( u1_u1_u6_n96 ) );
  NAND2_X1 u1_u1_u6_U57 (.ZN( u1_u1_u6_n100 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n98 ) );
  NAND2_X1 u1_u1_u6_U58 (.ZN( u1_u1_u6_n122 ) , .A1( u1_u1_u6_n94 ) , .A2( u1_u1_u6_n97 ) );
  INV_X1 u1_u1_u6_U59 (.A( u1_u1_u6_n139 ) , .ZN( u1_u1_u6_n160 ) );
  AOI22_X1 u1_u1_u6_U6 (.B2( u1_u1_u6_n101 ) , .A1( u1_u1_u6_n102 ) , .ZN( u1_u1_u6_n103 ) , .B1( u1_u1_u6_n160 ) , .A2( u1_u1_u6_n161 ) );
  NAND2_X1 u1_u1_u6_U60 (.ZN( u1_u1_u6_n113 ) , .A1( u1_u1_u6_n96 ) , .A2( u1_u1_u6_n98 ) );
  NOR2_X1 u1_u1_u6_U61 (.A2( u1_u1_X_40 ) , .A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n126 ) );
  NOR2_X1 u1_u1_u6_U62 (.A2( u1_u1_X_39 ) , .A1( u1_u1_X_42 ) , .ZN( u1_u1_u6_n92 ) );
  NOR2_X1 u1_u1_u6_U63 (.A2( u1_u1_X_39 ) , .A1( u1_u1_u6_n156 ) , .ZN( u1_u1_u6_n97 ) );
  NOR2_X1 u1_u1_u6_U64 (.A2( u1_u1_X_38 ) , .A1( u1_u1_u6_n165 ) , .ZN( u1_u1_u6_n95 ) );
  NOR2_X1 u1_u1_u6_U65 (.A2( u1_u1_X_41 ) , .ZN( u1_u1_u6_n111 ) , .A1( u1_u1_u6_n157 ) );
  NOR2_X1 u1_u1_u6_U66 (.A2( u1_u1_X_37 ) , .A1( u1_u1_u6_n162 ) , .ZN( u1_u1_u6_n94 ) );
  NOR2_X1 u1_u1_u6_U67 (.A2( u1_u1_X_37 ) , .A1( u1_u1_X_38 ) , .ZN( u1_u1_u6_n91 ) );
  NAND2_X1 u1_u1_u6_U68 (.A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n144 ) , .A2( u1_u1_u6_n157 ) );
  NAND2_X1 u1_u1_u6_U69 (.A2( u1_u1_X_40 ) , .A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n139 ) );
  NOR2_X1 u1_u1_u6_U7 (.A1( u1_u1_u6_n118 ) , .ZN( u1_u1_u6_n143 ) , .A2( u1_u1_u6_n168 ) );
  AND2_X1 u1_u1_u6_U70 (.A1( u1_u1_X_39 ) , .A2( u1_u1_u6_n156 ) , .ZN( u1_u1_u6_n96 ) );
  AND2_X1 u1_u1_u6_U71 (.A1( u1_u1_X_39 ) , .A2( u1_u1_X_42 ) , .ZN( u1_u1_u6_n99 ) );
  INV_X1 u1_u1_u6_U72 (.A( u1_u1_X_40 ) , .ZN( u1_u1_u6_n157 ) );
  INV_X1 u1_u1_u6_U73 (.A( u1_u1_X_37 ) , .ZN( u1_u1_u6_n165 ) );
  INV_X1 u1_u1_u6_U74 (.A( u1_u1_X_38 ) , .ZN( u1_u1_u6_n162 ) );
  INV_X1 u1_u1_u6_U75 (.A( u1_u1_X_42 ) , .ZN( u1_u1_u6_n156 ) );
  NAND4_X1 u1_u1_u6_U76 (.ZN( u1_out1_32 ) , .A4( u1_u1_u6_n103 ) , .A3( u1_u1_u6_n104 ) , .A2( u1_u1_u6_n105 ) , .A1( u1_u1_u6_n106 ) );
  AOI22_X1 u1_u1_u6_U77 (.ZN( u1_u1_u6_n105 ) , .A2( u1_u1_u6_n108 ) , .A1( u1_u1_u6_n118 ) , .B2( u1_u1_u6_n126 ) , .B1( u1_u1_u6_n171 ) );
  AOI22_X1 u1_u1_u6_U78 (.ZN( u1_u1_u6_n104 ) , .A1( u1_u1_u6_n111 ) , .B1( u1_u1_u6_n124 ) , .B2( u1_u1_u6_n151 ) , .A2( u1_u1_u6_n93 ) );
  NAND4_X1 u1_u1_u6_U79 (.ZN( u1_out1_12 ) , .A4( u1_u1_u6_n114 ) , .A3( u1_u1_u6_n115 ) , .A2( u1_u1_u6_n116 ) , .A1( u1_u1_u6_n117 ) );
  OAI21_X1 u1_u1_u6_U8 (.A( u1_u1_u6_n159 ) , .B1( u1_u1_u6_n169 ) , .B2( u1_u1_u6_n173 ) , .ZN( u1_u1_u6_n90 ) );
  OAI22_X1 u1_u1_u6_U80 (.B2( u1_u1_u6_n111 ) , .ZN( u1_u1_u6_n116 ) , .B1( u1_u1_u6_n126 ) , .A2( u1_u1_u6_n164 ) , .A1( u1_u1_u6_n167 ) );
  OAI21_X1 u1_u1_u6_U81 (.A( u1_u1_u6_n108 ) , .ZN( u1_u1_u6_n117 ) , .B2( u1_u1_u6_n141 ) , .B1( u1_u1_u6_n163 ) );
  OAI211_X1 u1_u1_u6_U82 (.ZN( u1_out1_7 ) , .B( u1_u1_u6_n153 ) , .C2( u1_u1_u6_n154 ) , .C1( u1_u1_u6_n155 ) , .A( u1_u1_u6_n174 ) );
  NOR3_X1 u1_u1_u6_U83 (.A1( u1_u1_u6_n141 ) , .ZN( u1_u1_u6_n154 ) , .A3( u1_u1_u6_n164 ) , .A2( u1_u1_u6_n171 ) );
  AOI211_X1 u1_u1_u6_U84 (.B( u1_u1_u6_n149 ) , .A( u1_u1_u6_n150 ) , .C2( u1_u1_u6_n151 ) , .C1( u1_u1_u6_n152 ) , .ZN( u1_u1_u6_n153 ) );
  OAI211_X1 u1_u1_u6_U85 (.ZN( u1_out1_22 ) , .B( u1_u1_u6_n137 ) , .A( u1_u1_u6_n138 ) , .C2( u1_u1_u6_n139 ) , .C1( u1_u1_u6_n140 ) );
  AND4_X1 u1_u1_u6_U86 (.A3( u1_u1_u6_n119 ) , .A1( u1_u1_u6_n120 ) , .A4( u1_u1_u6_n129 ) , .ZN( u1_u1_u6_n140 ) , .A2( u1_u1_u6_n143 ) );
  AOI22_X1 u1_u1_u6_U87 (.B1( u1_u1_u6_n124 ) , .A2( u1_u1_u6_n125 ) , .A1( u1_u1_u6_n126 ) , .ZN( u1_u1_u6_n138 ) , .B2( u1_u1_u6_n161 ) );
  NAND3_X1 u1_u1_u6_U88 (.A2( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n125 ) , .A1( u1_u1_u6_n130 ) , .A3( u1_u1_u6_n131 ) );
  NAND3_X1 u1_u1_u6_U89 (.A3( u1_u1_u6_n133 ) , .ZN( u1_u1_u6_n141 ) , .A1( u1_u1_u6_n145 ) , .A2( u1_u1_u6_n148 ) );
  INV_X1 u1_u1_u6_U9 (.ZN( u1_u1_u6_n172 ) , .A( u1_u1_u6_n88 ) );
  NAND3_X1 u1_u1_u6_U90 (.ZN( u1_u1_u6_n101 ) , .A3( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n121 ) , .A1( u1_u1_u6_n127 ) );
  NAND3_X1 u1_u1_u6_U91 (.ZN( u1_u1_u6_n102 ) , .A3( u1_u1_u6_n130 ) , .A2( u1_u1_u6_n145 ) , .A1( u1_u1_u6_n166 ) );
  NAND3_X1 u1_u1_u6_U92 (.A3( u1_u1_u6_n113 ) , .A1( u1_u1_u6_n119 ) , .A2( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n93 ) );
  NAND3_X1 u1_u1_u6_U93 (.ZN( u1_u1_u6_n142 ) , .A2( u1_u1_u6_n172 ) , .A3( u1_u1_u6_n89 ) , .A1( u1_u1_u6_n90 ) );
  AND3_X1 u1_u1_u7_U10 (.A3( u1_u1_u7_n110 ) , .A2( u1_u1_u7_n127 ) , .A1( u1_u1_u7_n132 ) , .ZN( u1_u1_u7_n92 ) );
  OAI21_X1 u1_u1_u7_U11 (.A( u1_u1_u7_n161 ) , .B1( u1_u1_u7_n168 ) , .B2( u1_u1_u7_n173 ) , .ZN( u1_u1_u7_n91 ) );
  AOI211_X1 u1_u1_u7_U12 (.A( u1_u1_u7_n117 ) , .ZN( u1_u1_u7_n118 ) , .C2( u1_u1_u7_n126 ) , .C1( u1_u1_u7_n177 ) , .B( u1_u1_u7_n180 ) );
  OAI22_X1 u1_u1_u7_U13 (.B1( u1_u1_u7_n115 ) , .ZN( u1_u1_u7_n117 ) , .A2( u1_u1_u7_n133 ) , .A1( u1_u1_u7_n137 ) , .B2( u1_u1_u7_n162 ) );
  INV_X1 u1_u1_u7_U14 (.A( u1_u1_u7_n116 ) , .ZN( u1_u1_u7_n180 ) );
  NOR3_X1 u1_u1_u7_U15 (.ZN( u1_u1_u7_n115 ) , .A3( u1_u1_u7_n145 ) , .A2( u1_u1_u7_n168 ) , .A1( u1_u1_u7_n169 ) );
  OAI211_X1 u1_u1_u7_U16 (.B( u1_u1_u7_n122 ) , .A( u1_u1_u7_n123 ) , .C2( u1_u1_u7_n124 ) , .ZN( u1_u1_u7_n154 ) , .C1( u1_u1_u7_n162 ) );
  AOI222_X1 u1_u1_u7_U17 (.ZN( u1_u1_u7_n122 ) , .C2( u1_u1_u7_n126 ) , .C1( u1_u1_u7_n145 ) , .B1( u1_u1_u7_n161 ) , .A2( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n170 ) , .A1( u1_u1_u7_n176 ) );
  INV_X1 u1_u1_u7_U18 (.A( u1_u1_u7_n133 ) , .ZN( u1_u1_u7_n176 ) );
  NOR3_X1 u1_u1_u7_U19 (.A2( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n135 ) , .ZN( u1_u1_u7_n136 ) , .A3( u1_u1_u7_n171 ) );
  NOR2_X1 u1_u1_u7_U20 (.A1( u1_u1_u7_n130 ) , .A2( u1_u1_u7_n134 ) , .ZN( u1_u1_u7_n153 ) );
  INV_X1 u1_u1_u7_U21 (.A( u1_u1_u7_n101 ) , .ZN( u1_u1_u7_n165 ) );
  NOR2_X1 u1_u1_u7_U22 (.ZN( u1_u1_u7_n111 ) , .A2( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n169 ) );
  AOI21_X1 u1_u1_u7_U23 (.ZN( u1_u1_u7_n104 ) , .B2( u1_u1_u7_n112 ) , .B1( u1_u1_u7_n127 ) , .A( u1_u1_u7_n164 ) );
  AOI21_X1 u1_u1_u7_U24 (.ZN( u1_u1_u7_n106 ) , .B1( u1_u1_u7_n133 ) , .B2( u1_u1_u7_n146 ) , .A( u1_u1_u7_n162 ) );
  AOI21_X1 u1_u1_u7_U25 (.A( u1_u1_u7_n101 ) , .ZN( u1_u1_u7_n107 ) , .B2( u1_u1_u7_n128 ) , .B1( u1_u1_u7_n175 ) );
  INV_X1 u1_u1_u7_U26 (.A( u1_u1_u7_n138 ) , .ZN( u1_u1_u7_n171 ) );
  INV_X1 u1_u1_u7_U27 (.A( u1_u1_u7_n131 ) , .ZN( u1_u1_u7_n177 ) );
  INV_X1 u1_u1_u7_U28 (.A( u1_u1_u7_n110 ) , .ZN( u1_u1_u7_n174 ) );
  NAND2_X1 u1_u1_u7_U29 (.A1( u1_u1_u7_n129 ) , .A2( u1_u1_u7_n132 ) , .ZN( u1_u1_u7_n149 ) );
  OAI21_X1 u1_u1_u7_U3 (.ZN( u1_u1_u7_n159 ) , .A( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n171 ) , .B1( u1_u1_u7_n174 ) );
  NAND2_X1 u1_u1_u7_U30 (.A1( u1_u1_u7_n113 ) , .A2( u1_u1_u7_n124 ) , .ZN( u1_u1_u7_n130 ) );
  INV_X1 u1_u1_u7_U31 (.A( u1_u1_u7_n112 ) , .ZN( u1_u1_u7_n173 ) );
  INV_X1 u1_u1_u7_U32 (.A( u1_u1_u7_n128 ) , .ZN( u1_u1_u7_n168 ) );
  INV_X1 u1_u1_u7_U33 (.A( u1_u1_u7_n148 ) , .ZN( u1_u1_u7_n169 ) );
  INV_X1 u1_u1_u7_U34 (.A( u1_u1_u7_n127 ) , .ZN( u1_u1_u7_n179 ) );
  NOR2_X1 u1_u1_u7_U35 (.ZN( u1_u1_u7_n101 ) , .A2( u1_u1_u7_n150 ) , .A1( u1_u1_u7_n156 ) );
  AOI211_X1 u1_u1_u7_U36 (.B( u1_u1_u7_n154 ) , .A( u1_u1_u7_n155 ) , .C1( u1_u1_u7_n156 ) , .ZN( u1_u1_u7_n157 ) , .C2( u1_u1_u7_n172 ) );
  INV_X1 u1_u1_u7_U37 (.A( u1_u1_u7_n153 ) , .ZN( u1_u1_u7_n172 ) );
  AOI211_X1 u1_u1_u7_U38 (.B( u1_u1_u7_n139 ) , .A( u1_u1_u7_n140 ) , .C2( u1_u1_u7_n141 ) , .ZN( u1_u1_u7_n142 ) , .C1( u1_u1_u7_n156 ) );
  NAND4_X1 u1_u1_u7_U39 (.A3( u1_u1_u7_n127 ) , .A2( u1_u1_u7_n128 ) , .A1( u1_u1_u7_n129 ) , .ZN( u1_u1_u7_n141 ) , .A4( u1_u1_u7_n147 ) );
  INV_X1 u1_u1_u7_U4 (.A( u1_u1_u7_n111 ) , .ZN( u1_u1_u7_n170 ) );
  AOI21_X1 u1_u1_u7_U40 (.A( u1_u1_u7_n137 ) , .B1( u1_u1_u7_n138 ) , .ZN( u1_u1_u7_n139 ) , .B2( u1_u1_u7_n146 ) );
  OAI22_X1 u1_u1_u7_U41 (.B1( u1_u1_u7_n136 ) , .ZN( u1_u1_u7_n140 ) , .A1( u1_u1_u7_n153 ) , .B2( u1_u1_u7_n162 ) , .A2( u1_u1_u7_n164 ) );
  AOI21_X1 u1_u1_u7_U42 (.ZN( u1_u1_u7_n123 ) , .B1( u1_u1_u7_n165 ) , .B2( u1_u1_u7_n177 ) , .A( u1_u1_u7_n97 ) );
  AOI21_X1 u1_u1_u7_U43 (.B2( u1_u1_u7_n113 ) , .B1( u1_u1_u7_n124 ) , .A( u1_u1_u7_n125 ) , .ZN( u1_u1_u7_n97 ) );
  INV_X1 u1_u1_u7_U44 (.A( u1_u1_u7_n125 ) , .ZN( u1_u1_u7_n161 ) );
  INV_X1 u1_u1_u7_U45 (.A( u1_u1_u7_n152 ) , .ZN( u1_u1_u7_n162 ) );
  AOI22_X1 u1_u1_u7_U46 (.A2( u1_u1_u7_n114 ) , .ZN( u1_u1_u7_n119 ) , .B1( u1_u1_u7_n130 ) , .A1( u1_u1_u7_n156 ) , .B2( u1_u1_u7_n165 ) );
  NAND2_X1 u1_u1_u7_U47 (.A2( u1_u1_u7_n112 ) , .ZN( u1_u1_u7_n114 ) , .A1( u1_u1_u7_n175 ) );
  AND2_X1 u1_u1_u7_U48 (.ZN( u1_u1_u7_n145 ) , .A2( u1_u1_u7_n98 ) , .A1( u1_u1_u7_n99 ) );
  NOR2_X1 u1_u1_u7_U49 (.ZN( u1_u1_u7_n137 ) , .A1( u1_u1_u7_n150 ) , .A2( u1_u1_u7_n161 ) );
  INV_X1 u1_u1_u7_U5 (.A( u1_u1_u7_n149 ) , .ZN( u1_u1_u7_n175 ) );
  AOI21_X1 u1_u1_u7_U50 (.ZN( u1_u1_u7_n105 ) , .B2( u1_u1_u7_n110 ) , .A( u1_u1_u7_n125 ) , .B1( u1_u1_u7_n147 ) );
  NAND2_X1 u1_u1_u7_U51 (.ZN( u1_u1_u7_n146 ) , .A1( u1_u1_u7_n95 ) , .A2( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U52 (.A2( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n147 ) , .A1( u1_u1_u7_n93 ) );
  NAND2_X1 u1_u1_u7_U53 (.A1( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n127 ) , .A2( u1_u1_u7_n99 ) );
  OR2_X1 u1_u1_u7_U54 (.ZN( u1_u1_u7_n126 ) , .A2( u1_u1_u7_n152 ) , .A1( u1_u1_u7_n156 ) );
  NAND2_X1 u1_u1_u7_U55 (.A2( u1_u1_u7_n102 ) , .A1( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n133 ) );
  NAND2_X1 u1_u1_u7_U56 (.ZN( u1_u1_u7_n112 ) , .A2( u1_u1_u7_n96 ) , .A1( u1_u1_u7_n99 ) );
  NAND2_X1 u1_u1_u7_U57 (.A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n128 ) , .A1( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U58 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n113 ) , .A2( u1_u1_u7_n93 ) );
  NAND2_X1 u1_u1_u7_U59 (.A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n124 ) , .A1( u1_u1_u7_n96 ) );
  INV_X1 u1_u1_u7_U6 (.A( u1_u1_u7_n154 ) , .ZN( u1_u1_u7_n178 ) );
  NAND2_X1 u1_u1_u7_U60 (.ZN( u1_u1_u7_n110 ) , .A1( u1_u1_u7_n95 ) , .A2( u1_u1_u7_n96 ) );
  INV_X1 u1_u1_u7_U61 (.A( u1_u1_u7_n150 ) , .ZN( u1_u1_u7_n164 ) );
  AND2_X1 u1_u1_u7_U62 (.ZN( u1_u1_u7_n134 ) , .A1( u1_u1_u7_n93 ) , .A2( u1_u1_u7_n98 ) );
  NAND2_X1 u1_u1_u7_U63 (.A1( u1_u1_u7_n100 ) , .A2( u1_u1_u7_n102 ) , .ZN( u1_u1_u7_n129 ) );
  NAND2_X1 u1_u1_u7_U64 (.A2( u1_u1_u7_n103 ) , .ZN( u1_u1_u7_n131 ) , .A1( u1_u1_u7_n95 ) );
  NAND2_X1 u1_u1_u7_U65 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n138 ) , .A2( u1_u1_u7_n99 ) );
  NAND2_X1 u1_u1_u7_U66 (.ZN( u1_u1_u7_n132 ) , .A1( u1_u1_u7_n93 ) , .A2( u1_u1_u7_n96 ) );
  NAND2_X1 u1_u1_u7_U67 (.A1( u1_u1_u7_n100 ) , .ZN( u1_u1_u7_n148 ) , .A2( u1_u1_u7_n95 ) );
  NOR2_X1 u1_u1_u7_U68 (.A2( u1_u1_X_47 ) , .ZN( u1_u1_u7_n150 ) , .A1( u1_u1_u7_n163 ) );
  NOR2_X1 u1_u1_u7_U69 (.A2( u1_u1_X_43 ) , .A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n103 ) );
  AOI211_X1 u1_u1_u7_U7 (.ZN( u1_u1_u7_n116 ) , .A( u1_u1_u7_n155 ) , .C1( u1_u1_u7_n161 ) , .C2( u1_u1_u7_n171 ) , .B( u1_u1_u7_n94 ) );
  NOR2_X1 u1_u1_u7_U70 (.A2( u1_u1_X_48 ) , .A1( u1_u1_u7_n166 ) , .ZN( u1_u1_u7_n95 ) );
  NOR2_X1 u1_u1_u7_U71 (.A2( u1_u1_X_45 ) , .A1( u1_u1_X_48 ) , .ZN( u1_u1_u7_n99 ) );
  NOR2_X1 u1_u1_u7_U72 (.A2( u1_u1_X_44 ) , .A1( u1_u1_u7_n167 ) , .ZN( u1_u1_u7_n98 ) );
  NOR2_X1 u1_u1_u7_U73 (.A2( u1_u1_X_46 ) , .A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n152 ) );
  AND2_X1 u1_u1_u7_U74 (.A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n156 ) , .A2( u1_u1_u7_n163 ) );
  NAND2_X1 u1_u1_u7_U75 (.A2( u1_u1_X_46 ) , .A1( u1_u1_X_47 ) , .ZN( u1_u1_u7_n125 ) );
  AND2_X1 u1_u1_u7_U76 (.A2( u1_u1_X_45 ) , .A1( u1_u1_X_48 ) , .ZN( u1_u1_u7_n102 ) );
  AND2_X1 u1_u1_u7_U77 (.A2( u1_u1_X_43 ) , .A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n96 ) );
  AND2_X1 u1_u1_u7_U78 (.A1( u1_u1_X_44 ) , .ZN( u1_u1_u7_n100 ) , .A2( u1_u1_u7_n167 ) );
  AND2_X1 u1_u1_u7_U79 (.A1( u1_u1_X_48 ) , .A2( u1_u1_u7_n166 ) , .ZN( u1_u1_u7_n93 ) );
  OAI222_X1 u1_u1_u7_U8 (.C2( u1_u1_u7_n101 ) , .B2( u1_u1_u7_n111 ) , .A1( u1_u1_u7_n113 ) , .C1( u1_u1_u7_n146 ) , .A2( u1_u1_u7_n162 ) , .B1( u1_u1_u7_n164 ) , .ZN( u1_u1_u7_n94 ) );
  INV_X1 u1_u1_u7_U80 (.A( u1_u1_X_46 ) , .ZN( u1_u1_u7_n163 ) );
  INV_X1 u1_u1_u7_U81 (.A( u1_u1_X_43 ) , .ZN( u1_u1_u7_n167 ) );
  INV_X1 u1_u1_u7_U82 (.A( u1_u1_X_45 ) , .ZN( u1_u1_u7_n166 ) );
  NAND4_X1 u1_u1_u7_U83 (.ZN( u1_out1_5 ) , .A4( u1_u1_u7_n108 ) , .A3( u1_u1_u7_n109 ) , .A1( u1_u1_u7_n116 ) , .A2( u1_u1_u7_n123 ) );
  AOI22_X1 u1_u1_u7_U84 (.ZN( u1_u1_u7_n109 ) , .A2( u1_u1_u7_n126 ) , .B2( u1_u1_u7_n145 ) , .B1( u1_u1_u7_n156 ) , .A1( u1_u1_u7_n171 ) );
  NOR4_X1 u1_u1_u7_U85 (.A4( u1_u1_u7_n104 ) , .A3( u1_u1_u7_n105 ) , .A2( u1_u1_u7_n106 ) , .A1( u1_u1_u7_n107 ) , .ZN( u1_u1_u7_n108 ) );
  NAND4_X1 u1_u1_u7_U86 (.ZN( u1_out1_27 ) , .A4( u1_u1_u7_n118 ) , .A3( u1_u1_u7_n119 ) , .A2( u1_u1_u7_n120 ) , .A1( u1_u1_u7_n121 ) );
  OAI21_X1 u1_u1_u7_U87 (.ZN( u1_u1_u7_n121 ) , .B2( u1_u1_u7_n145 ) , .A( u1_u1_u7_n150 ) , .B1( u1_u1_u7_n174 ) );
  OAI21_X1 u1_u1_u7_U88 (.ZN( u1_u1_u7_n120 ) , .A( u1_u1_u7_n161 ) , .B2( u1_u1_u7_n170 ) , .B1( u1_u1_u7_n179 ) );
  NAND4_X1 u1_u1_u7_U89 (.ZN( u1_out1_21 ) , .A4( u1_u1_u7_n157 ) , .A3( u1_u1_u7_n158 ) , .A2( u1_u1_u7_n159 ) , .A1( u1_u1_u7_n160 ) );
  OAI221_X1 u1_u1_u7_U9 (.C1( u1_u1_u7_n101 ) , .C2( u1_u1_u7_n147 ) , .ZN( u1_u1_u7_n155 ) , .B2( u1_u1_u7_n162 ) , .A( u1_u1_u7_n91 ) , .B1( u1_u1_u7_n92 ) );
  OAI21_X1 u1_u1_u7_U90 (.B1( u1_u1_u7_n145 ) , .ZN( u1_u1_u7_n160 ) , .A( u1_u1_u7_n161 ) , .B2( u1_u1_u7_n177 ) );
  AOI22_X1 u1_u1_u7_U91 (.B2( u1_u1_u7_n149 ) , .B1( u1_u1_u7_n150 ) , .A2( u1_u1_u7_n151 ) , .A1( u1_u1_u7_n152 ) , .ZN( u1_u1_u7_n158 ) );
  NAND4_X1 u1_u1_u7_U92 (.ZN( u1_out1_15 ) , .A4( u1_u1_u7_n142 ) , .A3( u1_u1_u7_n143 ) , .A2( u1_u1_u7_n144 ) , .A1( u1_u1_u7_n178 ) );
  OR2_X1 u1_u1_u7_U93 (.A2( u1_u1_u7_n125 ) , .A1( u1_u1_u7_n129 ) , .ZN( u1_u1_u7_n144 ) );
  AOI22_X1 u1_u1_u7_U94 (.A2( u1_u1_u7_n126 ) , .ZN( u1_u1_u7_n143 ) , .B2( u1_u1_u7_n165 ) , .B1( u1_u1_u7_n173 ) , .A1( u1_u1_u7_n174 ) );
  NAND3_X1 u1_u1_u7_U95 (.A3( u1_u1_u7_n146 ) , .A2( u1_u1_u7_n147 ) , .A1( u1_u1_u7_n148 ) , .ZN( u1_u1_u7_n151 ) );
  NAND3_X1 u1_u1_u7_U96 (.A3( u1_u1_u7_n131 ) , .A2( u1_u1_u7_n132 ) , .A1( u1_u1_u7_n133 ) , .ZN( u1_u1_u7_n135 ) );
  XOR2_X1 u1_u2_U10 (.B( u1_K3_45 ) , .A( u1_R1_30 ) , .Z( u1_u2_X_45 ) );
  XOR2_X1 u1_u2_U11 (.B( u1_K3_44 ) , .A( u1_R1_29 ) , .Z( u1_u2_X_44 ) );
  XOR2_X1 u1_u2_U12 (.B( u1_K3_43 ) , .A( u1_R1_28 ) , .Z( u1_u2_X_43 ) );
  XOR2_X1 u1_u2_U13 (.B( u1_K3_42 ) , .A( u1_R1_29 ) , .Z( u1_u2_X_42 ) );
  XOR2_X1 u1_u2_U14 (.B( u1_K3_41 ) , .A( u1_R1_28 ) , .Z( u1_u2_X_41 ) );
  XOR2_X1 u1_u2_U18 (.B( u1_K3_38 ) , .A( u1_R1_25 ) , .Z( u1_u2_X_38 ) );
  XOR2_X1 u1_u2_U19 (.B( u1_K3_37 ) , .A( u1_R1_24 ) , .Z( u1_u2_X_37 ) );
  XOR2_X1 u1_u2_U2 (.B( u1_K3_8 ) , .A( u1_R1_5 ) , .Z( u1_u2_X_8 ) );
  XOR2_X1 u1_u2_U20 (.B( u1_K3_36 ) , .A( u1_R1_25 ) , .Z( u1_u2_X_36 ) );
  XOR2_X1 u1_u2_U21 (.B( u1_K3_35 ) , .A( u1_R1_24 ) , .Z( u1_u2_X_35 ) );
  XOR2_X1 u1_u2_U24 (.B( u1_K3_32 ) , .A( u1_R1_21 ) , .Z( u1_u2_X_32 ) );
  XOR2_X1 u1_u2_U25 (.B( u1_K3_31 ) , .A( u1_R1_20 ) , .Z( u1_u2_X_31 ) );
  XOR2_X1 u1_u2_U26 (.B( u1_K3_30 ) , .A( u1_R1_21 ) , .Z( u1_u2_X_30 ) );
  XOR2_X1 u1_u2_U27 (.B( u1_K3_2 ) , .A( u1_R1_1 ) , .Z( u1_u2_X_2 ) );
  XOR2_X1 u1_u2_U28 (.B( u1_K3_29 ) , .A( u1_R1_20 ) , .Z( u1_u2_X_29 ) );
  XOR2_X1 u1_u2_U3 (.B( u1_K3_7 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_7 ) );
  XOR2_X1 u1_u2_U31 (.B( u1_K3_26 ) , .A( u1_R1_17 ) , .Z( u1_u2_X_26 ) );
  XOR2_X1 u1_u2_U32 (.B( u1_K3_25 ) , .A( u1_R1_16 ) , .Z( u1_u2_X_25 ) );
  XOR2_X1 u1_u2_U33 (.B( u1_K3_24 ) , .A( u1_R1_17 ) , .Z( u1_u2_X_24 ) );
  XOR2_X1 u1_u2_U34 (.B( u1_K3_23 ) , .A( u1_R1_16 ) , .Z( u1_u2_X_23 ) );
  XOR2_X1 u1_u2_U35 (.B( u1_K3_22 ) , .A( u1_R1_15 ) , .Z( u1_u2_X_22 ) );
  XOR2_X1 u1_u2_U36 (.B( u1_K3_21 ) , .A( u1_R1_14 ) , .Z( u1_u2_X_21 ) );
  XOR2_X1 u1_u2_U37 (.B( u1_K3_20 ) , .A( u1_R1_13 ) , .Z( u1_u2_X_20 ) );
  XOR2_X1 u1_u2_U38 (.B( u1_K3_1 ) , .A( u1_R1_32 ) , .Z( u1_u2_X_1 ) );
  XOR2_X1 u1_u2_U39 (.B( u1_K3_19 ) , .A( u1_R1_12 ) , .Z( u1_u2_X_19 ) );
  XOR2_X1 u1_u2_U4 (.B( u1_K3_6 ) , .A( u1_R1_5 ) , .Z( u1_u2_X_6 ) );
  XOR2_X1 u1_u2_U40 (.B( u1_K3_18 ) , .A( u1_R1_13 ) , .Z( u1_u2_X_18 ) );
  XOR2_X1 u1_u2_U41 (.B( u1_K3_17 ) , .A( u1_R1_12 ) , .Z( u1_u2_X_17 ) );
  XOR2_X1 u1_u2_U44 (.B( u1_K3_14 ) , .A( u1_R1_9 ) , .Z( u1_u2_X_14 ) );
  XOR2_X1 u1_u2_U45 (.B( u1_K3_13 ) , .A( u1_R1_8 ) , .Z( u1_u2_X_13 ) );
  XOR2_X1 u1_u2_U46 (.B( u1_K3_12 ) , .A( u1_R1_9 ) , .Z( u1_u2_X_12 ) );
  XOR2_X1 u1_u2_U47 (.B( u1_K3_11 ) , .A( u1_R1_8 ) , .Z( u1_u2_X_11 ) );
  XOR2_X1 u1_u2_U5 (.B( u1_K3_5 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_5 ) );
  XOR2_X1 u1_u2_U7 (.B( u1_K3_48 ) , .A( u1_R1_1 ) , .Z( u1_u2_X_48 ) );
  XOR2_X1 u1_u2_U8 (.B( u1_K3_47 ) , .A( u1_R1_32 ) , .Z( u1_u2_X_47 ) );
  XOR2_X1 u1_u2_U9 (.B( u1_K3_46 ) , .A( u1_R1_31 ) , .Z( u1_u2_X_46 ) );
  OAI22_X1 u1_u2_u3_U10 (.B1( u1_u2_u3_n113 ) , .A2( u1_u2_u3_n135 ) , .A1( u1_u2_u3_n150 ) , .B2( u1_u2_u3_n164 ) , .ZN( u1_u2_u3_n98 ) );
  OAI211_X1 u1_u2_u3_U11 (.B( u1_u2_u3_n106 ) , .ZN( u1_u2_u3_n119 ) , .C2( u1_u2_u3_n128 ) , .C1( u1_u2_u3_n167 ) , .A( u1_u2_u3_n181 ) );
  AOI221_X1 u1_u2_u3_U12 (.C1( u1_u2_u3_n105 ) , .ZN( u1_u2_u3_n106 ) , .A( u1_u2_u3_n131 ) , .B2( u1_u2_u3_n132 ) , .C2( u1_u2_u3_n133 ) , .B1( u1_u2_u3_n169 ) );
  INV_X1 u1_u2_u3_U13 (.ZN( u1_u2_u3_n181 ) , .A( u1_u2_u3_n98 ) );
  NAND2_X1 u1_u2_u3_U14 (.ZN( u1_u2_u3_n105 ) , .A2( u1_u2_u3_n130 ) , .A1( u1_u2_u3_n155 ) );
  AOI22_X1 u1_u2_u3_U15 (.B1( u1_u2_u3_n115 ) , .A2( u1_u2_u3_n116 ) , .ZN( u1_u2_u3_n123 ) , .B2( u1_u2_u3_n133 ) , .A1( u1_u2_u3_n169 ) );
  NAND2_X1 u1_u2_u3_U16 (.ZN( u1_u2_u3_n116 ) , .A2( u1_u2_u3_n151 ) , .A1( u1_u2_u3_n182 ) );
  NOR2_X1 u1_u2_u3_U17 (.ZN( u1_u2_u3_n126 ) , .A2( u1_u2_u3_n150 ) , .A1( u1_u2_u3_n164 ) );
  AOI21_X1 u1_u2_u3_U18 (.ZN( u1_u2_u3_n112 ) , .B2( u1_u2_u3_n146 ) , .B1( u1_u2_u3_n155 ) , .A( u1_u2_u3_n167 ) );
  NAND2_X1 u1_u2_u3_U19 (.A1( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n142 ) , .A2( u1_u2_u3_n164 ) );
  NAND2_X1 u1_u2_u3_U20 (.ZN( u1_u2_u3_n132 ) , .A2( u1_u2_u3_n152 ) , .A1( u1_u2_u3_n156 ) );
  AND2_X1 u1_u2_u3_U21 (.A2( u1_u2_u3_n113 ) , .A1( u1_u2_u3_n114 ) , .ZN( u1_u2_u3_n151 ) );
  INV_X1 u1_u2_u3_U22 (.A( u1_u2_u3_n133 ) , .ZN( u1_u2_u3_n165 ) );
  INV_X1 u1_u2_u3_U23 (.A( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n170 ) );
  NAND2_X1 u1_u2_u3_U24 (.A1( u1_u2_u3_n107 ) , .A2( u1_u2_u3_n108 ) , .ZN( u1_u2_u3_n140 ) );
  NAND2_X1 u1_u2_u3_U25 (.ZN( u1_u2_u3_n117 ) , .A1( u1_u2_u3_n124 ) , .A2( u1_u2_u3_n148 ) );
  NAND2_X1 u1_u2_u3_U26 (.ZN( u1_u2_u3_n143 ) , .A1( u1_u2_u3_n165 ) , .A2( u1_u2_u3_n167 ) );
  INV_X1 u1_u2_u3_U27 (.A( u1_u2_u3_n130 ) , .ZN( u1_u2_u3_n177 ) );
  INV_X1 u1_u2_u3_U28 (.A( u1_u2_u3_n128 ) , .ZN( u1_u2_u3_n176 ) );
  INV_X1 u1_u2_u3_U29 (.A( u1_u2_u3_n155 ) , .ZN( u1_u2_u3_n174 ) );
  INV_X1 u1_u2_u3_U3 (.A( u1_u2_u3_n129 ) , .ZN( u1_u2_u3_n183 ) );
  INV_X1 u1_u2_u3_U30 (.A( u1_u2_u3_n139 ) , .ZN( u1_u2_u3_n185 ) );
  NOR2_X1 u1_u2_u3_U31 (.ZN( u1_u2_u3_n135 ) , .A2( u1_u2_u3_n141 ) , .A1( u1_u2_u3_n169 ) );
  OAI222_X1 u1_u2_u3_U32 (.C2( u1_u2_u3_n107 ) , .A2( u1_u2_u3_n108 ) , .B1( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n138 ) , .B2( u1_u2_u3_n146 ) , .C1( u1_u2_u3_n154 ) , .A1( u1_u2_u3_n164 ) );
  NOR4_X1 u1_u2_u3_U33 (.A4( u1_u2_u3_n157 ) , .A3( u1_u2_u3_n158 ) , .A2( u1_u2_u3_n159 ) , .A1( u1_u2_u3_n160 ) , .ZN( u1_u2_u3_n161 ) );
  AOI21_X1 u1_u2_u3_U34 (.B2( u1_u2_u3_n152 ) , .B1( u1_u2_u3_n153 ) , .ZN( u1_u2_u3_n158 ) , .A( u1_u2_u3_n164 ) );
  AOI21_X1 u1_u2_u3_U35 (.A( u1_u2_u3_n154 ) , .B2( u1_u2_u3_n155 ) , .B1( u1_u2_u3_n156 ) , .ZN( u1_u2_u3_n157 ) );
  AOI21_X1 u1_u2_u3_U36 (.A( u1_u2_u3_n149 ) , .B2( u1_u2_u3_n150 ) , .B1( u1_u2_u3_n151 ) , .ZN( u1_u2_u3_n159 ) );
  AOI211_X1 u1_u2_u3_U37 (.ZN( u1_u2_u3_n109 ) , .A( u1_u2_u3_n119 ) , .C2( u1_u2_u3_n129 ) , .B( u1_u2_u3_n138 ) , .C1( u1_u2_u3_n141 ) );
  AOI211_X1 u1_u2_u3_U38 (.B( u1_u2_u3_n119 ) , .A( u1_u2_u3_n120 ) , .C2( u1_u2_u3_n121 ) , .ZN( u1_u2_u3_n122 ) , .C1( u1_u2_u3_n179 ) );
  INV_X1 u1_u2_u3_U39 (.A( u1_u2_u3_n156 ) , .ZN( u1_u2_u3_n179 ) );
  INV_X1 u1_u2_u3_U4 (.A( u1_u2_u3_n140 ) , .ZN( u1_u2_u3_n182 ) );
  OAI22_X1 u1_u2_u3_U40 (.B1( u1_u2_u3_n118 ) , .ZN( u1_u2_u3_n120 ) , .A1( u1_u2_u3_n135 ) , .B2( u1_u2_u3_n154 ) , .A2( u1_u2_u3_n178 ) );
  AND3_X1 u1_u2_u3_U41 (.ZN( u1_u2_u3_n118 ) , .A2( u1_u2_u3_n124 ) , .A1( u1_u2_u3_n144 ) , .A3( u1_u2_u3_n152 ) );
  INV_X1 u1_u2_u3_U42 (.A( u1_u2_u3_n121 ) , .ZN( u1_u2_u3_n164 ) );
  NAND2_X1 u1_u2_u3_U43 (.ZN( u1_u2_u3_n133 ) , .A1( u1_u2_u3_n154 ) , .A2( u1_u2_u3_n164 ) );
  OAI211_X1 u1_u2_u3_U44 (.B( u1_u2_u3_n127 ) , .ZN( u1_u2_u3_n139 ) , .C1( u1_u2_u3_n150 ) , .C2( u1_u2_u3_n154 ) , .A( u1_u2_u3_n184 ) );
  INV_X1 u1_u2_u3_U45 (.A( u1_u2_u3_n125 ) , .ZN( u1_u2_u3_n184 ) );
  AOI221_X1 u1_u2_u3_U46 (.A( u1_u2_u3_n126 ) , .ZN( u1_u2_u3_n127 ) , .C2( u1_u2_u3_n132 ) , .C1( u1_u2_u3_n169 ) , .B2( u1_u2_u3_n170 ) , .B1( u1_u2_u3_n174 ) );
  OAI22_X1 u1_u2_u3_U47 (.A1( u1_u2_u3_n124 ) , .ZN( u1_u2_u3_n125 ) , .B2( u1_u2_u3_n145 ) , .A2( u1_u2_u3_n165 ) , .B1( u1_u2_u3_n167 ) );
  NOR2_X1 u1_u2_u3_U48 (.A1( u1_u2_u3_n113 ) , .ZN( u1_u2_u3_n131 ) , .A2( u1_u2_u3_n154 ) );
  NAND2_X1 u1_u2_u3_U49 (.A1( u1_u2_u3_n103 ) , .ZN( u1_u2_u3_n150 ) , .A2( u1_u2_u3_n99 ) );
  INV_X1 u1_u2_u3_U5 (.A( u1_u2_u3_n117 ) , .ZN( u1_u2_u3_n178 ) );
  NAND2_X1 u1_u2_u3_U50 (.A2( u1_u2_u3_n102 ) , .ZN( u1_u2_u3_n155 ) , .A1( u1_u2_u3_n97 ) );
  INV_X1 u1_u2_u3_U51 (.A( u1_u2_u3_n141 ) , .ZN( u1_u2_u3_n167 ) );
  AOI21_X1 u1_u2_u3_U52 (.B2( u1_u2_u3_n114 ) , .B1( u1_u2_u3_n146 ) , .A( u1_u2_u3_n154 ) , .ZN( u1_u2_u3_n94 ) );
  AOI21_X1 u1_u2_u3_U53 (.ZN( u1_u2_u3_n110 ) , .B2( u1_u2_u3_n142 ) , .B1( u1_u2_u3_n186 ) , .A( u1_u2_u3_n95 ) );
  INV_X1 u1_u2_u3_U54 (.A( u1_u2_u3_n145 ) , .ZN( u1_u2_u3_n186 ) );
  AOI21_X1 u1_u2_u3_U55 (.B1( u1_u2_u3_n124 ) , .A( u1_u2_u3_n149 ) , .B2( u1_u2_u3_n155 ) , .ZN( u1_u2_u3_n95 ) );
  INV_X1 u1_u2_u3_U56 (.A( u1_u2_u3_n149 ) , .ZN( u1_u2_u3_n169 ) );
  NAND2_X1 u1_u2_u3_U57 (.ZN( u1_u2_u3_n124 ) , .A1( u1_u2_u3_n96 ) , .A2( u1_u2_u3_n97 ) );
  NAND2_X1 u1_u2_u3_U58 (.A2( u1_u2_u3_n100 ) , .ZN( u1_u2_u3_n146 ) , .A1( u1_u2_u3_n96 ) );
  NAND2_X1 u1_u2_u3_U59 (.A1( u1_u2_u3_n101 ) , .ZN( u1_u2_u3_n145 ) , .A2( u1_u2_u3_n99 ) );
  AOI221_X1 u1_u2_u3_U6 (.A( u1_u2_u3_n131 ) , .C2( u1_u2_u3_n132 ) , .C1( u1_u2_u3_n133 ) , .ZN( u1_u2_u3_n134 ) , .B1( u1_u2_u3_n143 ) , .B2( u1_u2_u3_n177 ) );
  NAND2_X1 u1_u2_u3_U60 (.A1( u1_u2_u3_n100 ) , .ZN( u1_u2_u3_n156 ) , .A2( u1_u2_u3_n99 ) );
  NAND2_X1 u1_u2_u3_U61 (.A2( u1_u2_u3_n101 ) , .A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n148 ) );
  NAND2_X1 u1_u2_u3_U62 (.A1( u1_u2_u3_n100 ) , .A2( u1_u2_u3_n102 ) , .ZN( u1_u2_u3_n128 ) );
  NAND2_X1 u1_u2_u3_U63 (.A2( u1_u2_u3_n101 ) , .A1( u1_u2_u3_n102 ) , .ZN( u1_u2_u3_n152 ) );
  NAND2_X1 u1_u2_u3_U64 (.A2( u1_u2_u3_n101 ) , .ZN( u1_u2_u3_n114 ) , .A1( u1_u2_u3_n96 ) );
  NAND2_X1 u1_u2_u3_U65 (.ZN( u1_u2_u3_n107 ) , .A1( u1_u2_u3_n97 ) , .A2( u1_u2_u3_n99 ) );
  NAND2_X1 u1_u2_u3_U66 (.A2( u1_u2_u3_n100 ) , .A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n113 ) );
  NAND2_X1 u1_u2_u3_U67 (.A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n153 ) , .A2( u1_u2_u3_n97 ) );
  NAND2_X1 u1_u2_u3_U68 (.A2( u1_u2_u3_n103 ) , .A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n130 ) );
  NAND2_X1 u1_u2_u3_U69 (.A2( u1_u2_u3_n103 ) , .ZN( u1_u2_u3_n144 ) , .A1( u1_u2_u3_n96 ) );
  OAI22_X1 u1_u2_u3_U7 (.B2( u1_u2_u3_n147 ) , .A2( u1_u2_u3_n148 ) , .ZN( u1_u2_u3_n160 ) , .B1( u1_u2_u3_n165 ) , .A1( u1_u2_u3_n168 ) );
  NAND2_X1 u1_u2_u3_U70 (.A1( u1_u2_u3_n102 ) , .A2( u1_u2_u3_n103 ) , .ZN( u1_u2_u3_n108 ) );
  NOR2_X1 u1_u2_u3_U71 (.A2( u1_u2_X_19 ) , .A1( u1_u2_X_20 ) , .ZN( u1_u2_u3_n99 ) );
  NOR2_X1 u1_u2_u3_U72 (.A2( u1_u2_X_21 ) , .A1( u1_u2_X_24 ) , .ZN( u1_u2_u3_n103 ) );
  NOR2_X1 u1_u2_u3_U73 (.A2( u1_u2_X_24 ) , .A1( u1_u2_u3_n171 ) , .ZN( u1_u2_u3_n97 ) );
  NOR2_X1 u1_u2_u3_U74 (.A2( u1_u2_X_23 ) , .ZN( u1_u2_u3_n141 ) , .A1( u1_u2_u3_n166 ) );
  NOR2_X1 u1_u2_u3_U75 (.A2( u1_u2_X_19 ) , .A1( u1_u2_u3_n172 ) , .ZN( u1_u2_u3_n96 ) );
  NAND2_X1 u1_u2_u3_U76 (.A1( u1_u2_X_22 ) , .A2( u1_u2_X_23 ) , .ZN( u1_u2_u3_n154 ) );
  NAND2_X1 u1_u2_u3_U77 (.A1( u1_u2_X_23 ) , .ZN( u1_u2_u3_n149 ) , .A2( u1_u2_u3_n166 ) );
  NOR2_X1 u1_u2_u3_U78 (.A2( u1_u2_X_22 ) , .A1( u1_u2_X_23 ) , .ZN( u1_u2_u3_n121 ) );
  AND2_X1 u1_u2_u3_U79 (.A1( u1_u2_X_24 ) , .ZN( u1_u2_u3_n101 ) , .A2( u1_u2_u3_n171 ) );
  AND3_X1 u1_u2_u3_U8 (.A3( u1_u2_u3_n144 ) , .A2( u1_u2_u3_n145 ) , .A1( u1_u2_u3_n146 ) , .ZN( u1_u2_u3_n147 ) );
  AND2_X1 u1_u2_u3_U80 (.A1( u1_u2_X_19 ) , .ZN( u1_u2_u3_n102 ) , .A2( u1_u2_u3_n172 ) );
  AND2_X1 u1_u2_u3_U81 (.A1( u1_u2_X_21 ) , .A2( u1_u2_X_24 ) , .ZN( u1_u2_u3_n100 ) );
  AND2_X1 u1_u2_u3_U82 (.A2( u1_u2_X_19 ) , .A1( u1_u2_X_20 ) , .ZN( u1_u2_u3_n104 ) );
  INV_X1 u1_u2_u3_U83 (.A( u1_u2_X_22 ) , .ZN( u1_u2_u3_n166 ) );
  INV_X1 u1_u2_u3_U84 (.A( u1_u2_X_21 ) , .ZN( u1_u2_u3_n171 ) );
  INV_X1 u1_u2_u3_U85 (.A( u1_u2_X_20 ) , .ZN( u1_u2_u3_n172 ) );
  OR4_X1 u1_u2_u3_U86 (.ZN( u1_out2_10 ) , .A4( u1_u2_u3_n136 ) , .A3( u1_u2_u3_n137 ) , .A1( u1_u2_u3_n138 ) , .A2( u1_u2_u3_n139 ) );
  OAI222_X1 u1_u2_u3_U87 (.C1( u1_u2_u3_n128 ) , .ZN( u1_u2_u3_n137 ) , .B1( u1_u2_u3_n148 ) , .A2( u1_u2_u3_n150 ) , .B2( u1_u2_u3_n154 ) , .C2( u1_u2_u3_n164 ) , .A1( u1_u2_u3_n167 ) );
  OAI221_X1 u1_u2_u3_U88 (.A( u1_u2_u3_n134 ) , .B2( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n136 ) , .C1( u1_u2_u3_n149 ) , .B1( u1_u2_u3_n151 ) , .C2( u1_u2_u3_n183 ) );
  NAND4_X1 u1_u2_u3_U89 (.ZN( u1_out2_26 ) , .A4( u1_u2_u3_n109 ) , .A3( u1_u2_u3_n110 ) , .A2( u1_u2_u3_n111 ) , .A1( u1_u2_u3_n173 ) );
  INV_X1 u1_u2_u3_U9 (.A( u1_u2_u3_n143 ) , .ZN( u1_u2_u3_n168 ) );
  INV_X1 u1_u2_u3_U90 (.ZN( u1_u2_u3_n173 ) , .A( u1_u2_u3_n94 ) );
  OAI21_X1 u1_u2_u3_U91 (.ZN( u1_u2_u3_n111 ) , .B2( u1_u2_u3_n117 ) , .A( u1_u2_u3_n133 ) , .B1( u1_u2_u3_n176 ) );
  NAND4_X1 u1_u2_u3_U92 (.ZN( u1_out2_20 ) , .A4( u1_u2_u3_n122 ) , .A3( u1_u2_u3_n123 ) , .A1( u1_u2_u3_n175 ) , .A2( u1_u2_u3_n180 ) );
  INV_X1 u1_u2_u3_U93 (.A( u1_u2_u3_n112 ) , .ZN( u1_u2_u3_n175 ) );
  INV_X1 u1_u2_u3_U94 (.A( u1_u2_u3_n126 ) , .ZN( u1_u2_u3_n180 ) );
  NAND4_X1 u1_u2_u3_U95 (.ZN( u1_out2_1 ) , .A4( u1_u2_u3_n161 ) , .A3( u1_u2_u3_n162 ) , .A2( u1_u2_u3_n163 ) , .A1( u1_u2_u3_n185 ) );
  NAND2_X1 u1_u2_u3_U96 (.ZN( u1_u2_u3_n163 ) , .A2( u1_u2_u3_n170 ) , .A1( u1_u2_u3_n176 ) );
  AOI22_X1 u1_u2_u3_U97 (.B2( u1_u2_u3_n140 ) , .B1( u1_u2_u3_n141 ) , .A2( u1_u2_u3_n142 ) , .ZN( u1_u2_u3_n162 ) , .A1( u1_u2_u3_n177 ) );
  NAND3_X1 u1_u2_u3_U98 (.A1( u1_u2_u3_n114 ) , .ZN( u1_u2_u3_n115 ) , .A2( u1_u2_u3_n145 ) , .A3( u1_u2_u3_n153 ) );
  NAND3_X1 u1_u2_u3_U99 (.ZN( u1_u2_u3_n129 ) , .A2( u1_u2_u3_n144 ) , .A1( u1_u2_u3_n153 ) , .A3( u1_u2_u3_n182 ) );
  AND3_X1 u1_u2_u7_U10 (.A3( u1_u2_u7_n110 ) , .A2( u1_u2_u7_n127 ) , .A1( u1_u2_u7_n132 ) , .ZN( u1_u2_u7_n92 ) );
  OAI21_X1 u1_u2_u7_U11 (.A( u1_u2_u7_n161 ) , .B1( u1_u2_u7_n168 ) , .B2( u1_u2_u7_n173 ) , .ZN( u1_u2_u7_n91 ) );
  AOI211_X1 u1_u2_u7_U12 (.A( u1_u2_u7_n117 ) , .ZN( u1_u2_u7_n118 ) , .C2( u1_u2_u7_n126 ) , .C1( u1_u2_u7_n177 ) , .B( u1_u2_u7_n180 ) );
  OAI22_X1 u1_u2_u7_U13 (.B1( u1_u2_u7_n115 ) , .ZN( u1_u2_u7_n117 ) , .A2( u1_u2_u7_n133 ) , .A1( u1_u2_u7_n137 ) , .B2( u1_u2_u7_n162 ) );
  INV_X1 u1_u2_u7_U14 (.A( u1_u2_u7_n116 ) , .ZN( u1_u2_u7_n180 ) );
  NOR3_X1 u1_u2_u7_U15 (.ZN( u1_u2_u7_n115 ) , .A3( u1_u2_u7_n145 ) , .A2( u1_u2_u7_n168 ) , .A1( u1_u2_u7_n169 ) );
  OAI211_X1 u1_u2_u7_U16 (.B( u1_u2_u7_n122 ) , .A( u1_u2_u7_n123 ) , .C2( u1_u2_u7_n124 ) , .ZN( u1_u2_u7_n154 ) , .C1( u1_u2_u7_n162 ) );
  AOI222_X1 u1_u2_u7_U17 (.ZN( u1_u2_u7_n122 ) , .C2( u1_u2_u7_n126 ) , .C1( u1_u2_u7_n145 ) , .B1( u1_u2_u7_n161 ) , .A2( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n170 ) , .A1( u1_u2_u7_n176 ) );
  INV_X1 u1_u2_u7_U18 (.A( u1_u2_u7_n133 ) , .ZN( u1_u2_u7_n176 ) );
  NOR3_X1 u1_u2_u7_U19 (.A2( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n135 ) , .ZN( u1_u2_u7_n136 ) , .A3( u1_u2_u7_n171 ) );
  NOR2_X1 u1_u2_u7_U20 (.A1( u1_u2_u7_n130 ) , .A2( u1_u2_u7_n134 ) , .ZN( u1_u2_u7_n153 ) );
  INV_X1 u1_u2_u7_U21 (.A( u1_u2_u7_n101 ) , .ZN( u1_u2_u7_n165 ) );
  NOR2_X1 u1_u2_u7_U22 (.ZN( u1_u2_u7_n111 ) , .A2( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n169 ) );
  AOI21_X1 u1_u2_u7_U23 (.ZN( u1_u2_u7_n104 ) , .B2( u1_u2_u7_n112 ) , .B1( u1_u2_u7_n127 ) , .A( u1_u2_u7_n164 ) );
  AOI21_X1 u1_u2_u7_U24 (.ZN( u1_u2_u7_n106 ) , .B1( u1_u2_u7_n133 ) , .B2( u1_u2_u7_n146 ) , .A( u1_u2_u7_n162 ) );
  AOI21_X1 u1_u2_u7_U25 (.A( u1_u2_u7_n101 ) , .ZN( u1_u2_u7_n107 ) , .B2( u1_u2_u7_n128 ) , .B1( u1_u2_u7_n175 ) );
  INV_X1 u1_u2_u7_U26 (.A( u1_u2_u7_n138 ) , .ZN( u1_u2_u7_n171 ) );
  INV_X1 u1_u2_u7_U27 (.A( u1_u2_u7_n131 ) , .ZN( u1_u2_u7_n177 ) );
  INV_X1 u1_u2_u7_U28 (.A( u1_u2_u7_n110 ) , .ZN( u1_u2_u7_n174 ) );
  NAND2_X1 u1_u2_u7_U29 (.A1( u1_u2_u7_n129 ) , .A2( u1_u2_u7_n132 ) , .ZN( u1_u2_u7_n149 ) );
  OAI21_X1 u1_u2_u7_U3 (.ZN( u1_u2_u7_n159 ) , .A( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n171 ) , .B1( u1_u2_u7_n174 ) );
  NAND2_X1 u1_u2_u7_U30 (.A1( u1_u2_u7_n113 ) , .A2( u1_u2_u7_n124 ) , .ZN( u1_u2_u7_n130 ) );
  INV_X1 u1_u2_u7_U31 (.A( u1_u2_u7_n112 ) , .ZN( u1_u2_u7_n173 ) );
  INV_X1 u1_u2_u7_U32 (.A( u1_u2_u7_n128 ) , .ZN( u1_u2_u7_n168 ) );
  INV_X1 u1_u2_u7_U33 (.A( u1_u2_u7_n148 ) , .ZN( u1_u2_u7_n169 ) );
  INV_X1 u1_u2_u7_U34 (.A( u1_u2_u7_n127 ) , .ZN( u1_u2_u7_n179 ) );
  NOR2_X1 u1_u2_u7_U35 (.ZN( u1_u2_u7_n101 ) , .A2( u1_u2_u7_n150 ) , .A1( u1_u2_u7_n156 ) );
  AOI211_X1 u1_u2_u7_U36 (.B( u1_u2_u7_n154 ) , .A( u1_u2_u7_n155 ) , .C1( u1_u2_u7_n156 ) , .ZN( u1_u2_u7_n157 ) , .C2( u1_u2_u7_n172 ) );
  INV_X1 u1_u2_u7_U37 (.A( u1_u2_u7_n153 ) , .ZN( u1_u2_u7_n172 ) );
  AOI211_X1 u1_u2_u7_U38 (.B( u1_u2_u7_n139 ) , .A( u1_u2_u7_n140 ) , .C2( u1_u2_u7_n141 ) , .ZN( u1_u2_u7_n142 ) , .C1( u1_u2_u7_n156 ) );
  NAND4_X1 u1_u2_u7_U39 (.A3( u1_u2_u7_n127 ) , .A2( u1_u2_u7_n128 ) , .A1( u1_u2_u7_n129 ) , .ZN( u1_u2_u7_n141 ) , .A4( u1_u2_u7_n147 ) );
  INV_X1 u1_u2_u7_U4 (.A( u1_u2_u7_n111 ) , .ZN( u1_u2_u7_n170 ) );
  AOI21_X1 u1_u2_u7_U40 (.A( u1_u2_u7_n137 ) , .B1( u1_u2_u7_n138 ) , .ZN( u1_u2_u7_n139 ) , .B2( u1_u2_u7_n146 ) );
  OAI22_X1 u1_u2_u7_U41 (.B1( u1_u2_u7_n136 ) , .ZN( u1_u2_u7_n140 ) , .A1( u1_u2_u7_n153 ) , .B2( u1_u2_u7_n162 ) , .A2( u1_u2_u7_n164 ) );
  AOI21_X1 u1_u2_u7_U42 (.ZN( u1_u2_u7_n123 ) , .B1( u1_u2_u7_n165 ) , .B2( u1_u2_u7_n177 ) , .A( u1_u2_u7_n97 ) );
  AOI21_X1 u1_u2_u7_U43 (.B2( u1_u2_u7_n113 ) , .B1( u1_u2_u7_n124 ) , .A( u1_u2_u7_n125 ) , .ZN( u1_u2_u7_n97 ) );
  INV_X1 u1_u2_u7_U44 (.A( u1_u2_u7_n125 ) , .ZN( u1_u2_u7_n161 ) );
  INV_X1 u1_u2_u7_U45 (.A( u1_u2_u7_n152 ) , .ZN( u1_u2_u7_n162 ) );
  AOI22_X1 u1_u2_u7_U46 (.A2( u1_u2_u7_n114 ) , .ZN( u1_u2_u7_n119 ) , .B1( u1_u2_u7_n130 ) , .A1( u1_u2_u7_n156 ) , .B2( u1_u2_u7_n165 ) );
  NAND2_X1 u1_u2_u7_U47 (.A2( u1_u2_u7_n112 ) , .ZN( u1_u2_u7_n114 ) , .A1( u1_u2_u7_n175 ) );
  AND2_X1 u1_u2_u7_U48 (.ZN( u1_u2_u7_n145 ) , .A2( u1_u2_u7_n98 ) , .A1( u1_u2_u7_n99 ) );
  NOR2_X1 u1_u2_u7_U49 (.ZN( u1_u2_u7_n137 ) , .A1( u1_u2_u7_n150 ) , .A2( u1_u2_u7_n161 ) );
  INV_X1 u1_u2_u7_U5 (.A( u1_u2_u7_n149 ) , .ZN( u1_u2_u7_n175 ) );
  AOI21_X1 u1_u2_u7_U50 (.ZN( u1_u2_u7_n105 ) , .B2( u1_u2_u7_n110 ) , .A( u1_u2_u7_n125 ) , .B1( u1_u2_u7_n147 ) );
  NAND2_X1 u1_u2_u7_U51 (.ZN( u1_u2_u7_n146 ) , .A1( u1_u2_u7_n95 ) , .A2( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U52 (.A2( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n147 ) , .A1( u1_u2_u7_n93 ) );
  NAND2_X1 u1_u2_u7_U53 (.A1( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n127 ) , .A2( u1_u2_u7_n99 ) );
  OR2_X1 u1_u2_u7_U54 (.ZN( u1_u2_u7_n126 ) , .A2( u1_u2_u7_n152 ) , .A1( u1_u2_u7_n156 ) );
  NAND2_X1 u1_u2_u7_U55 (.A2( u1_u2_u7_n102 ) , .A1( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n133 ) );
  NAND2_X1 u1_u2_u7_U56 (.ZN( u1_u2_u7_n112 ) , .A2( u1_u2_u7_n96 ) , .A1( u1_u2_u7_n99 ) );
  NAND2_X1 u1_u2_u7_U57 (.A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n128 ) , .A1( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U58 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n113 ) , .A2( u1_u2_u7_n93 ) );
  NAND2_X1 u1_u2_u7_U59 (.A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n124 ) , .A1( u1_u2_u7_n96 ) );
  INV_X1 u1_u2_u7_U6 (.A( u1_u2_u7_n154 ) , .ZN( u1_u2_u7_n178 ) );
  NAND2_X1 u1_u2_u7_U60 (.ZN( u1_u2_u7_n110 ) , .A1( u1_u2_u7_n95 ) , .A2( u1_u2_u7_n96 ) );
  INV_X1 u1_u2_u7_U61 (.A( u1_u2_u7_n150 ) , .ZN( u1_u2_u7_n164 ) );
  AND2_X1 u1_u2_u7_U62 (.ZN( u1_u2_u7_n134 ) , .A1( u1_u2_u7_n93 ) , .A2( u1_u2_u7_n98 ) );
  NAND2_X1 u1_u2_u7_U63 (.A1( u1_u2_u7_n100 ) , .A2( u1_u2_u7_n102 ) , .ZN( u1_u2_u7_n129 ) );
  NAND2_X1 u1_u2_u7_U64 (.A2( u1_u2_u7_n103 ) , .ZN( u1_u2_u7_n131 ) , .A1( u1_u2_u7_n95 ) );
  NAND2_X1 u1_u2_u7_U65 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n138 ) , .A2( u1_u2_u7_n99 ) );
  NAND2_X1 u1_u2_u7_U66 (.ZN( u1_u2_u7_n132 ) , .A1( u1_u2_u7_n93 ) , .A2( u1_u2_u7_n96 ) );
  NAND2_X1 u1_u2_u7_U67 (.A1( u1_u2_u7_n100 ) , .ZN( u1_u2_u7_n148 ) , .A2( u1_u2_u7_n95 ) );
  NOR2_X1 u1_u2_u7_U68 (.A2( u1_u2_X_47 ) , .ZN( u1_u2_u7_n150 ) , .A1( u1_u2_u7_n163 ) );
  NOR2_X1 u1_u2_u7_U69 (.A2( u1_u2_X_43 ) , .A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n103 ) );
  AOI211_X1 u1_u2_u7_U7 (.ZN( u1_u2_u7_n116 ) , .A( u1_u2_u7_n155 ) , .C1( u1_u2_u7_n161 ) , .C2( u1_u2_u7_n171 ) , .B( u1_u2_u7_n94 ) );
  NOR2_X1 u1_u2_u7_U70 (.A2( u1_u2_X_48 ) , .A1( u1_u2_u7_n166 ) , .ZN( u1_u2_u7_n95 ) );
  NOR2_X1 u1_u2_u7_U71 (.A2( u1_u2_X_45 ) , .A1( u1_u2_X_48 ) , .ZN( u1_u2_u7_n99 ) );
  NOR2_X1 u1_u2_u7_U72 (.A2( u1_u2_X_44 ) , .A1( u1_u2_u7_n167 ) , .ZN( u1_u2_u7_n98 ) );
  NOR2_X1 u1_u2_u7_U73 (.A2( u1_u2_X_46 ) , .A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n152 ) );
  AND2_X1 u1_u2_u7_U74 (.A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n156 ) , .A2( u1_u2_u7_n163 ) );
  NAND2_X1 u1_u2_u7_U75 (.A2( u1_u2_X_46 ) , .A1( u1_u2_X_47 ) , .ZN( u1_u2_u7_n125 ) );
  AND2_X1 u1_u2_u7_U76 (.A2( u1_u2_X_45 ) , .A1( u1_u2_X_48 ) , .ZN( u1_u2_u7_n102 ) );
  AND2_X1 u1_u2_u7_U77 (.A2( u1_u2_X_43 ) , .A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n96 ) );
  AND2_X1 u1_u2_u7_U78 (.A1( u1_u2_X_44 ) , .ZN( u1_u2_u7_n100 ) , .A2( u1_u2_u7_n167 ) );
  AND2_X1 u1_u2_u7_U79 (.A1( u1_u2_X_48 ) , .A2( u1_u2_u7_n166 ) , .ZN( u1_u2_u7_n93 ) );
  OAI222_X1 u1_u2_u7_U8 (.C2( u1_u2_u7_n101 ) , .B2( u1_u2_u7_n111 ) , .A1( u1_u2_u7_n113 ) , .C1( u1_u2_u7_n146 ) , .A2( u1_u2_u7_n162 ) , .B1( u1_u2_u7_n164 ) , .ZN( u1_u2_u7_n94 ) );
  INV_X1 u1_u2_u7_U80 (.A( u1_u2_X_46 ) , .ZN( u1_u2_u7_n163 ) );
  INV_X1 u1_u2_u7_U81 (.A( u1_u2_X_43 ) , .ZN( u1_u2_u7_n167 ) );
  INV_X1 u1_u2_u7_U82 (.A( u1_u2_X_45 ) , .ZN( u1_u2_u7_n166 ) );
  NAND4_X1 u1_u2_u7_U83 (.ZN( u1_out2_5 ) , .A4( u1_u2_u7_n108 ) , .A3( u1_u2_u7_n109 ) , .A1( u1_u2_u7_n116 ) , .A2( u1_u2_u7_n123 ) );
  AOI22_X1 u1_u2_u7_U84 (.ZN( u1_u2_u7_n109 ) , .A2( u1_u2_u7_n126 ) , .B2( u1_u2_u7_n145 ) , .B1( u1_u2_u7_n156 ) , .A1( u1_u2_u7_n171 ) );
  NOR4_X1 u1_u2_u7_U85 (.A4( u1_u2_u7_n104 ) , .A3( u1_u2_u7_n105 ) , .A2( u1_u2_u7_n106 ) , .A1( u1_u2_u7_n107 ) , .ZN( u1_u2_u7_n108 ) );
  NAND4_X1 u1_u2_u7_U86 (.ZN( u1_out2_27 ) , .A4( u1_u2_u7_n118 ) , .A3( u1_u2_u7_n119 ) , .A2( u1_u2_u7_n120 ) , .A1( u1_u2_u7_n121 ) );
  OAI21_X1 u1_u2_u7_U87 (.ZN( u1_u2_u7_n121 ) , .B2( u1_u2_u7_n145 ) , .A( u1_u2_u7_n150 ) , .B1( u1_u2_u7_n174 ) );
  OAI21_X1 u1_u2_u7_U88 (.ZN( u1_u2_u7_n120 ) , .A( u1_u2_u7_n161 ) , .B2( u1_u2_u7_n170 ) , .B1( u1_u2_u7_n179 ) );
  NAND4_X1 u1_u2_u7_U89 (.ZN( u1_out2_21 ) , .A4( u1_u2_u7_n157 ) , .A3( u1_u2_u7_n158 ) , .A2( u1_u2_u7_n159 ) , .A1( u1_u2_u7_n160 ) );
  OAI221_X1 u1_u2_u7_U9 (.C1( u1_u2_u7_n101 ) , .C2( u1_u2_u7_n147 ) , .ZN( u1_u2_u7_n155 ) , .B2( u1_u2_u7_n162 ) , .A( u1_u2_u7_n91 ) , .B1( u1_u2_u7_n92 ) );
  OAI21_X1 u1_u2_u7_U90 (.B1( u1_u2_u7_n145 ) , .ZN( u1_u2_u7_n160 ) , .A( u1_u2_u7_n161 ) , .B2( u1_u2_u7_n177 ) );
  AOI22_X1 u1_u2_u7_U91 (.B2( u1_u2_u7_n149 ) , .B1( u1_u2_u7_n150 ) , .A2( u1_u2_u7_n151 ) , .A1( u1_u2_u7_n152 ) , .ZN( u1_u2_u7_n158 ) );
  NAND4_X1 u1_u2_u7_U92 (.ZN( u1_out2_15 ) , .A4( u1_u2_u7_n142 ) , .A3( u1_u2_u7_n143 ) , .A2( u1_u2_u7_n144 ) , .A1( u1_u2_u7_n178 ) );
  OR2_X1 u1_u2_u7_U93 (.A2( u1_u2_u7_n125 ) , .A1( u1_u2_u7_n129 ) , .ZN( u1_u2_u7_n144 ) );
  AOI22_X1 u1_u2_u7_U94 (.A2( u1_u2_u7_n126 ) , .ZN( u1_u2_u7_n143 ) , .B2( u1_u2_u7_n165 ) , .B1( u1_u2_u7_n173 ) , .A1( u1_u2_u7_n174 ) );
  NAND3_X1 u1_u2_u7_U95 (.A3( u1_u2_u7_n146 ) , .A2( u1_u2_u7_n147 ) , .A1( u1_u2_u7_n148 ) , .ZN( u1_u2_u7_n151 ) );
  NAND3_X1 u1_u2_u7_U96 (.A3( u1_u2_u7_n131 ) , .A2( u1_u2_u7_n132 ) , .A1( u1_u2_u7_n133 ) , .ZN( u1_u2_u7_n135 ) );
  XOR2_X1 u1_u3_U11 (.B( u1_K4_44 ) , .A( u1_R2_29 ) , .Z( u1_u3_X_44 ) );
  XOR2_X1 u1_u3_U12 (.B( u1_K4_43 ) , .A( u1_R2_28 ) , .Z( u1_u3_X_43 ) );
  XOR2_X1 u1_u3_U13 (.B( u1_K4_42 ) , .A( u1_R2_29 ) , .Z( u1_u3_X_42 ) );
  XOR2_X1 u1_u3_U14 (.B( u1_K4_41 ) , .A( u1_R2_28 ) , .Z( u1_u3_X_41 ) );
  XOR2_X1 u1_u3_U18 (.B( u1_K4_38 ) , .A( u1_R2_25 ) , .Z( u1_u3_X_38 ) );
  XOR2_X1 u1_u3_U19 (.B( u1_K4_37 ) , .A( u1_R2_24 ) , .Z( u1_u3_X_37 ) );
  XOR2_X1 u1_u3_U2 (.B( u1_K4_8 ) , .A( u1_R2_5 ) , .Z( u1_u3_X_8 ) );
  XOR2_X1 u1_u3_U20 (.B( u1_K4_36 ) , .A( u1_R2_25 ) , .Z( u1_u3_X_36 ) );
  XOR2_X1 u1_u3_U21 (.B( u1_K4_35 ) , .A( u1_R2_24 ) , .Z( u1_u3_X_35 ) );
  XOR2_X1 u1_u3_U27 (.B( u1_K4_2 ) , .A( u1_R2_1 ) , .Z( u1_u3_X_2 ) );
  XOR2_X1 u1_u3_U3 (.B( u1_K4_7 ) , .A( u1_R2_4 ) , .Z( u1_u3_X_7 ) );
  XOR2_X1 u1_u3_U31 (.B( u1_K4_26 ) , .A( u1_R2_17 ) , .Z( u1_u3_X_26 ) );
  XOR2_X1 u1_u3_U32 (.B( u1_K4_25 ) , .A( u1_R2_16 ) , .Z( u1_u3_X_25 ) );
  XOR2_X1 u1_u3_U33 (.B( u1_K4_24 ) , .A( u1_R2_17 ) , .Z( u1_u3_X_24 ) );
  XOR2_X1 u1_u3_U34 (.B( u1_K4_23 ) , .A( u1_R2_16 ) , .Z( u1_u3_X_23 ) );
  XOR2_X1 u1_u3_U35 (.B( u1_K4_22 ) , .A( u1_R2_15 ) , .Z( u1_u3_X_22 ) );
  XOR2_X1 u1_u3_U36 (.B( u1_K4_21 ) , .A( u1_R2_14 ) , .Z( u1_u3_X_21 ) );
  XOR2_X1 u1_u3_U37 (.B( u1_K4_20 ) , .A( u1_R2_13 ) , .Z( u1_u3_X_20 ) );
  XOR2_X1 u1_u3_U38 (.B( u1_K4_1 ) , .A( u1_R2_32 ) , .Z( u1_u3_X_1 ) );
  XOR2_X1 u1_u3_U39 (.B( u1_K4_19 ) , .A( u1_R2_12 ) , .Z( u1_u3_X_19 ) );
  XOR2_X1 u1_u3_U4 (.B( u1_K4_6 ) , .A( u1_R2_5 ) , .Z( u1_u3_X_6 ) );
  XOR2_X1 u1_u3_U40 (.B( u1_K4_18 ) , .A( u1_R2_13 ) , .Z( u1_u3_X_18 ) );
  XOR2_X1 u1_u3_U41 (.B( u1_K4_17 ) , .A( u1_R2_12 ) , .Z( u1_u3_X_17 ) );
  XOR2_X1 u1_u3_U44 (.B( u1_K4_14 ) , .A( u1_R2_9 ) , .Z( u1_u3_X_14 ) );
  XOR2_X1 u1_u3_U45 (.B( u1_K4_13 ) , .A( u1_R2_8 ) , .Z( u1_u3_X_13 ) );
  XOR2_X1 u1_u3_U46 (.B( u1_K4_12 ) , .A( u1_R2_9 ) , .Z( u1_u3_X_12 ) );
  XOR2_X1 u1_u3_U47 (.B( u1_K4_11 ) , .A( u1_R2_8 ) , .Z( u1_u3_X_11 ) );
  XOR2_X1 u1_u3_U5 (.B( u1_K4_5 ) , .A( u1_R2_4 ) , .Z( u1_u3_X_5 ) );
  XOR2_X1 u1_u3_U7 (.B( u1_K4_48 ) , .A( u1_R2_1 ) , .Z( u1_u3_X_48 ) );
  XOR2_X1 u1_u3_U8 (.B( u1_K4_47 ) , .A( u1_R2_32 ) , .Z( u1_u3_X_47 ) );
  OAI22_X1 u1_u3_u3_U10 (.B1( u1_u3_u3_n113 ) , .A2( u1_u3_u3_n135 ) , .A1( u1_u3_u3_n150 ) , .B2( u1_u3_u3_n164 ) , .ZN( u1_u3_u3_n98 ) );
  OAI211_X1 u1_u3_u3_U11 (.B( u1_u3_u3_n106 ) , .ZN( u1_u3_u3_n119 ) , .C2( u1_u3_u3_n128 ) , .C1( u1_u3_u3_n167 ) , .A( u1_u3_u3_n181 ) );
  AOI221_X1 u1_u3_u3_U12 (.C1( u1_u3_u3_n105 ) , .ZN( u1_u3_u3_n106 ) , .A( u1_u3_u3_n131 ) , .B2( u1_u3_u3_n132 ) , .C2( u1_u3_u3_n133 ) , .B1( u1_u3_u3_n169 ) );
  INV_X1 u1_u3_u3_U13 (.ZN( u1_u3_u3_n181 ) , .A( u1_u3_u3_n98 ) );
  NAND2_X1 u1_u3_u3_U14 (.ZN( u1_u3_u3_n105 ) , .A2( u1_u3_u3_n130 ) , .A1( u1_u3_u3_n155 ) );
  AOI22_X1 u1_u3_u3_U15 (.B1( u1_u3_u3_n115 ) , .A2( u1_u3_u3_n116 ) , .ZN( u1_u3_u3_n123 ) , .B2( u1_u3_u3_n133 ) , .A1( u1_u3_u3_n169 ) );
  NAND2_X1 u1_u3_u3_U16 (.ZN( u1_u3_u3_n116 ) , .A2( u1_u3_u3_n151 ) , .A1( u1_u3_u3_n182 ) );
  NOR2_X1 u1_u3_u3_U17 (.ZN( u1_u3_u3_n126 ) , .A2( u1_u3_u3_n150 ) , .A1( u1_u3_u3_n164 ) );
  AOI21_X1 u1_u3_u3_U18 (.ZN( u1_u3_u3_n112 ) , .B2( u1_u3_u3_n146 ) , .B1( u1_u3_u3_n155 ) , .A( u1_u3_u3_n167 ) );
  NAND2_X1 u1_u3_u3_U19 (.A1( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n142 ) , .A2( u1_u3_u3_n164 ) );
  NAND2_X1 u1_u3_u3_U20 (.ZN( u1_u3_u3_n132 ) , .A2( u1_u3_u3_n152 ) , .A1( u1_u3_u3_n156 ) );
  INV_X1 u1_u3_u3_U21 (.A( u1_u3_u3_n133 ) , .ZN( u1_u3_u3_n165 ) );
  NAND2_X1 u1_u3_u3_U22 (.ZN( u1_u3_u3_n143 ) , .A1( u1_u3_u3_n165 ) , .A2( u1_u3_u3_n167 ) );
  AND2_X1 u1_u3_u3_U23 (.A2( u1_u3_u3_n113 ) , .A1( u1_u3_u3_n114 ) , .ZN( u1_u3_u3_n151 ) );
  INV_X1 u1_u3_u3_U24 (.A( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n170 ) );
  NAND2_X1 u1_u3_u3_U25 (.A1( u1_u3_u3_n107 ) , .A2( u1_u3_u3_n108 ) , .ZN( u1_u3_u3_n140 ) );
  NAND2_X1 u1_u3_u3_U26 (.ZN( u1_u3_u3_n117 ) , .A1( u1_u3_u3_n124 ) , .A2( u1_u3_u3_n148 ) );
  INV_X1 u1_u3_u3_U27 (.A( u1_u3_u3_n130 ) , .ZN( u1_u3_u3_n177 ) );
  INV_X1 u1_u3_u3_U28 (.A( u1_u3_u3_n128 ) , .ZN( u1_u3_u3_n176 ) );
  INV_X1 u1_u3_u3_U29 (.A( u1_u3_u3_n155 ) , .ZN( u1_u3_u3_n174 ) );
  INV_X1 u1_u3_u3_U3 (.A( u1_u3_u3_n140 ) , .ZN( u1_u3_u3_n182 ) );
  INV_X1 u1_u3_u3_U30 (.A( u1_u3_u3_n139 ) , .ZN( u1_u3_u3_n185 ) );
  NOR2_X1 u1_u3_u3_U31 (.ZN( u1_u3_u3_n135 ) , .A2( u1_u3_u3_n141 ) , .A1( u1_u3_u3_n169 ) );
  INV_X1 u1_u3_u3_U32 (.A( u1_u3_u3_n156 ) , .ZN( u1_u3_u3_n179 ) );
  OAI22_X1 u1_u3_u3_U33 (.B1( u1_u3_u3_n118 ) , .ZN( u1_u3_u3_n120 ) , .A1( u1_u3_u3_n135 ) , .B2( u1_u3_u3_n154 ) , .A2( u1_u3_u3_n178 ) );
  AND3_X1 u1_u3_u3_U34 (.ZN( u1_u3_u3_n118 ) , .A2( u1_u3_u3_n124 ) , .A1( u1_u3_u3_n144 ) , .A3( u1_u3_u3_n152 ) );
  OAI222_X1 u1_u3_u3_U35 (.C2( u1_u3_u3_n107 ) , .A2( u1_u3_u3_n108 ) , .B1( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n138 ) , .B2( u1_u3_u3_n146 ) , .C1( u1_u3_u3_n154 ) , .A1( u1_u3_u3_n164 ) );
  NOR4_X1 u1_u3_u3_U36 (.A4( u1_u3_u3_n157 ) , .A3( u1_u3_u3_n158 ) , .A2( u1_u3_u3_n159 ) , .A1( u1_u3_u3_n160 ) , .ZN( u1_u3_u3_n161 ) );
  AOI21_X1 u1_u3_u3_U37 (.B2( u1_u3_u3_n152 ) , .B1( u1_u3_u3_n153 ) , .ZN( u1_u3_u3_n158 ) , .A( u1_u3_u3_n164 ) );
  AOI21_X1 u1_u3_u3_U38 (.A( u1_u3_u3_n149 ) , .B2( u1_u3_u3_n150 ) , .B1( u1_u3_u3_n151 ) , .ZN( u1_u3_u3_n159 ) );
  AOI21_X1 u1_u3_u3_U39 (.A( u1_u3_u3_n154 ) , .B2( u1_u3_u3_n155 ) , .B1( u1_u3_u3_n156 ) , .ZN( u1_u3_u3_n157 ) );
  INV_X1 u1_u3_u3_U4 (.A( u1_u3_u3_n129 ) , .ZN( u1_u3_u3_n183 ) );
  AOI211_X1 u1_u3_u3_U40 (.ZN( u1_u3_u3_n109 ) , .A( u1_u3_u3_n119 ) , .C2( u1_u3_u3_n129 ) , .B( u1_u3_u3_n138 ) , .C1( u1_u3_u3_n141 ) );
  INV_X1 u1_u3_u3_U41 (.A( u1_u3_u3_n121 ) , .ZN( u1_u3_u3_n164 ) );
  NAND2_X1 u1_u3_u3_U42 (.ZN( u1_u3_u3_n133 ) , .A1( u1_u3_u3_n154 ) , .A2( u1_u3_u3_n164 ) );
  OAI211_X1 u1_u3_u3_U43 (.B( u1_u3_u3_n127 ) , .ZN( u1_u3_u3_n139 ) , .C1( u1_u3_u3_n150 ) , .C2( u1_u3_u3_n154 ) , .A( u1_u3_u3_n184 ) );
  INV_X1 u1_u3_u3_U44 (.A( u1_u3_u3_n125 ) , .ZN( u1_u3_u3_n184 ) );
  AOI221_X1 u1_u3_u3_U45 (.A( u1_u3_u3_n126 ) , .ZN( u1_u3_u3_n127 ) , .C2( u1_u3_u3_n132 ) , .C1( u1_u3_u3_n169 ) , .B2( u1_u3_u3_n170 ) , .B1( u1_u3_u3_n174 ) );
  OAI22_X1 u1_u3_u3_U46 (.A1( u1_u3_u3_n124 ) , .ZN( u1_u3_u3_n125 ) , .B2( u1_u3_u3_n145 ) , .A2( u1_u3_u3_n165 ) , .B1( u1_u3_u3_n167 ) );
  NOR2_X1 u1_u3_u3_U47 (.A1( u1_u3_u3_n113 ) , .ZN( u1_u3_u3_n131 ) , .A2( u1_u3_u3_n154 ) );
  NAND2_X1 u1_u3_u3_U48 (.A1( u1_u3_u3_n103 ) , .ZN( u1_u3_u3_n150 ) , .A2( u1_u3_u3_n99 ) );
  NAND2_X1 u1_u3_u3_U49 (.A2( u1_u3_u3_n102 ) , .ZN( u1_u3_u3_n155 ) , .A1( u1_u3_u3_n97 ) );
  INV_X1 u1_u3_u3_U5 (.A( u1_u3_u3_n117 ) , .ZN( u1_u3_u3_n178 ) );
  INV_X1 u1_u3_u3_U50 (.A( u1_u3_u3_n141 ) , .ZN( u1_u3_u3_n167 ) );
  AOI21_X1 u1_u3_u3_U51 (.B2( u1_u3_u3_n114 ) , .B1( u1_u3_u3_n146 ) , .A( u1_u3_u3_n154 ) , .ZN( u1_u3_u3_n94 ) );
  AOI21_X1 u1_u3_u3_U52 (.ZN( u1_u3_u3_n110 ) , .B2( u1_u3_u3_n142 ) , .B1( u1_u3_u3_n186 ) , .A( u1_u3_u3_n95 ) );
  INV_X1 u1_u3_u3_U53 (.A( u1_u3_u3_n145 ) , .ZN( u1_u3_u3_n186 ) );
  AOI21_X1 u1_u3_u3_U54 (.B1( u1_u3_u3_n124 ) , .A( u1_u3_u3_n149 ) , .B2( u1_u3_u3_n155 ) , .ZN( u1_u3_u3_n95 ) );
  INV_X1 u1_u3_u3_U55 (.A( u1_u3_u3_n149 ) , .ZN( u1_u3_u3_n169 ) );
  NAND2_X1 u1_u3_u3_U56 (.ZN( u1_u3_u3_n124 ) , .A1( u1_u3_u3_n96 ) , .A2( u1_u3_u3_n97 ) );
  NAND2_X1 u1_u3_u3_U57 (.A2( u1_u3_u3_n100 ) , .ZN( u1_u3_u3_n146 ) , .A1( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U58 (.A1( u1_u3_u3_n101 ) , .ZN( u1_u3_u3_n145 ) , .A2( u1_u3_u3_n99 ) );
  NAND2_X1 u1_u3_u3_U59 (.A1( u1_u3_u3_n100 ) , .ZN( u1_u3_u3_n156 ) , .A2( u1_u3_u3_n99 ) );
  AOI221_X1 u1_u3_u3_U6 (.A( u1_u3_u3_n131 ) , .C2( u1_u3_u3_n132 ) , .C1( u1_u3_u3_n133 ) , .ZN( u1_u3_u3_n134 ) , .B1( u1_u3_u3_n143 ) , .B2( u1_u3_u3_n177 ) );
  NAND2_X1 u1_u3_u3_U60 (.A2( u1_u3_u3_n101 ) , .A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n148 ) );
  NAND2_X1 u1_u3_u3_U61 (.A1( u1_u3_u3_n100 ) , .A2( u1_u3_u3_n102 ) , .ZN( u1_u3_u3_n128 ) );
  NAND2_X1 u1_u3_u3_U62 (.A2( u1_u3_u3_n101 ) , .A1( u1_u3_u3_n102 ) , .ZN( u1_u3_u3_n152 ) );
  NAND2_X1 u1_u3_u3_U63 (.A2( u1_u3_u3_n101 ) , .ZN( u1_u3_u3_n114 ) , .A1( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U64 (.ZN( u1_u3_u3_n107 ) , .A1( u1_u3_u3_n97 ) , .A2( u1_u3_u3_n99 ) );
  NAND2_X1 u1_u3_u3_U65 (.A2( u1_u3_u3_n100 ) , .A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n113 ) );
  NAND2_X1 u1_u3_u3_U66 (.A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n153 ) , .A2( u1_u3_u3_n97 ) );
  NAND2_X1 u1_u3_u3_U67 (.A2( u1_u3_u3_n103 ) , .A1( u1_u3_u3_n104 ) , .ZN( u1_u3_u3_n130 ) );
  NAND2_X1 u1_u3_u3_U68 (.A2( u1_u3_u3_n103 ) , .ZN( u1_u3_u3_n144 ) , .A1( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U69 (.A1( u1_u3_u3_n102 ) , .A2( u1_u3_u3_n103 ) , .ZN( u1_u3_u3_n108 ) );
  OAI22_X1 u1_u3_u3_U7 (.B2( u1_u3_u3_n147 ) , .A2( u1_u3_u3_n148 ) , .ZN( u1_u3_u3_n160 ) , .B1( u1_u3_u3_n165 ) , .A1( u1_u3_u3_n168 ) );
  NOR2_X1 u1_u3_u3_U70 (.A2( u1_u3_X_19 ) , .A1( u1_u3_X_20 ) , .ZN( u1_u3_u3_n99 ) );
  NOR2_X1 u1_u3_u3_U71 (.A2( u1_u3_X_21 ) , .A1( u1_u3_X_24 ) , .ZN( u1_u3_u3_n103 ) );
  NOR2_X1 u1_u3_u3_U72 (.A2( u1_u3_X_24 ) , .A1( u1_u3_u3_n171 ) , .ZN( u1_u3_u3_n97 ) );
  NOR2_X1 u1_u3_u3_U73 (.A2( u1_u3_X_19 ) , .A1( u1_u3_u3_n172 ) , .ZN( u1_u3_u3_n96 ) );
  NAND2_X1 u1_u3_u3_U74 (.A1( u1_u3_X_22 ) , .A2( u1_u3_X_23 ) , .ZN( u1_u3_u3_n154 ) );
  AND2_X1 u1_u3_u3_U75 (.A1( u1_u3_X_24 ) , .ZN( u1_u3_u3_n101 ) , .A2( u1_u3_u3_n171 ) );
  AND2_X1 u1_u3_u3_U76 (.A1( u1_u3_X_19 ) , .ZN( u1_u3_u3_n102 ) , .A2( u1_u3_u3_n172 ) );
  AND2_X1 u1_u3_u3_U77 (.A1( u1_u3_X_21 ) , .A2( u1_u3_X_24 ) , .ZN( u1_u3_u3_n100 ) );
  AND2_X1 u1_u3_u3_U78 (.A2( u1_u3_X_19 ) , .A1( u1_u3_X_20 ) , .ZN( u1_u3_u3_n104 ) );
  INV_X1 u1_u3_u3_U79 (.A( u1_u3_X_21 ) , .ZN( u1_u3_u3_n171 ) );
  AND3_X1 u1_u3_u3_U8 (.A3( u1_u3_u3_n144 ) , .A2( u1_u3_u3_n145 ) , .A1( u1_u3_u3_n146 ) , .ZN( u1_u3_u3_n147 ) );
  INV_X1 u1_u3_u3_U80 (.A( u1_u3_X_20 ) , .ZN( u1_u3_u3_n172 ) );
  INV_X1 u1_u3_u3_U81 (.A( u1_u3_X_22 ) , .ZN( u1_u3_u3_n166 ) );
  NAND4_X1 u1_u3_u3_U82 (.ZN( u1_out3_26 ) , .A4( u1_u3_u3_n109 ) , .A3( u1_u3_u3_n110 ) , .A2( u1_u3_u3_n111 ) , .A1( u1_u3_u3_n173 ) );
  INV_X1 u1_u3_u3_U83 (.ZN( u1_u3_u3_n173 ) , .A( u1_u3_u3_n94 ) );
  OAI21_X1 u1_u3_u3_U84 (.ZN( u1_u3_u3_n111 ) , .B2( u1_u3_u3_n117 ) , .A( u1_u3_u3_n133 ) , .B1( u1_u3_u3_n176 ) );
  NAND4_X1 u1_u3_u3_U85 (.ZN( u1_out3_1 ) , .A4( u1_u3_u3_n161 ) , .A3( u1_u3_u3_n162 ) , .A2( u1_u3_u3_n163 ) , .A1( u1_u3_u3_n185 ) );
  NAND2_X1 u1_u3_u3_U86 (.ZN( u1_u3_u3_n163 ) , .A2( u1_u3_u3_n170 ) , .A1( u1_u3_u3_n176 ) );
  AOI22_X1 u1_u3_u3_U87 (.B2( u1_u3_u3_n140 ) , .B1( u1_u3_u3_n141 ) , .A2( u1_u3_u3_n142 ) , .ZN( u1_u3_u3_n162 ) , .A1( u1_u3_u3_n177 ) );
  NAND4_X1 u1_u3_u3_U88 (.ZN( u1_out3_20 ) , .A4( u1_u3_u3_n122 ) , .A3( u1_u3_u3_n123 ) , .A1( u1_u3_u3_n175 ) , .A2( u1_u3_u3_n180 ) );
  INV_X1 u1_u3_u3_U89 (.A( u1_u3_u3_n126 ) , .ZN( u1_u3_u3_n180 ) );
  INV_X1 u1_u3_u3_U9 (.A( u1_u3_u3_n143 ) , .ZN( u1_u3_u3_n168 ) );
  INV_X1 u1_u3_u3_U90 (.A( u1_u3_u3_n112 ) , .ZN( u1_u3_u3_n175 ) );
  OR4_X1 u1_u3_u3_U91 (.ZN( u1_out3_10 ) , .A4( u1_u3_u3_n136 ) , .A3( u1_u3_u3_n137 ) , .A1( u1_u3_u3_n138 ) , .A2( u1_u3_u3_n139 ) );
  OAI222_X1 u1_u3_u3_U92 (.C1( u1_u3_u3_n128 ) , .ZN( u1_u3_u3_n137 ) , .B1( u1_u3_u3_n148 ) , .A2( u1_u3_u3_n150 ) , .B2( u1_u3_u3_n154 ) , .C2( u1_u3_u3_n164 ) , .A1( u1_u3_u3_n167 ) );
  AOI211_X1 u1_u3_u3_U93 (.B( u1_u3_u3_n119 ) , .A( u1_u3_u3_n120 ) , .C2( u1_u3_u3_n121 ) , .ZN( u1_u3_u3_n122 ) , .C1( u1_u3_u3_n179 ) );
  OAI221_X1 u1_u3_u3_U94 (.A( u1_u3_u3_n134 ) , .B2( u1_u3_u3_n135 ) , .ZN( u1_u3_u3_n136 ) , .C1( u1_u3_u3_n149 ) , .B1( u1_u3_u3_n151 ) , .C2( u1_u3_u3_n183 ) );
  NOR2_X1 u1_u3_u3_U95 (.A2( u1_u3_X_23 ) , .ZN( u1_u3_u3_n141 ) , .A1( u1_u3_u3_n166 ) );
  NAND2_X1 u1_u3_u3_U96 (.A1( u1_u3_X_23 ) , .ZN( u1_u3_u3_n149 ) , .A2( u1_u3_u3_n166 ) );
  NOR2_X1 u1_u3_u3_U97 (.A2( u1_u3_X_22 ) , .A1( u1_u3_X_23 ) , .ZN( u1_u3_u3_n121 ) );
  NAND3_X1 u1_u3_u3_U98 (.A1( u1_u3_u3_n114 ) , .ZN( u1_u3_u3_n115 ) , .A2( u1_u3_u3_n145 ) , .A3( u1_u3_u3_n153 ) );
  NAND3_X1 u1_u3_u3_U99 (.ZN( u1_u3_u3_n129 ) , .A2( u1_u3_u3_n144 ) , .A1( u1_u3_u3_n153 ) , .A3( u1_u3_u3_n182 ) );
  XOR2_X1 u1_u4_U10 (.B( u1_K5_45 ) , .A( u1_R3_30 ) , .Z( u1_u4_X_45 ) );
  XOR2_X1 u1_u4_U11 (.B( u1_K5_44 ) , .A( u1_R3_29 ) , .Z( u1_u4_X_44 ) );
  XOR2_X1 u1_u4_U12 (.B( u1_K5_43 ) , .A( u1_R3_28 ) , .Z( u1_u4_X_43 ) );
  XOR2_X1 u1_u4_U13 (.B( u1_K5_42 ) , .A( u1_R3_29 ) , .Z( u1_u4_X_42 ) );
  XOR2_X1 u1_u4_U14 (.B( u1_K5_41 ) , .A( u1_R3_28 ) , .Z( u1_u4_X_41 ) );
  XOR2_X1 u1_u4_U18 (.B( u1_K5_38 ) , .A( u1_R3_25 ) , .Z( u1_u4_X_38 ) );
  XOR2_X1 u1_u4_U19 (.B( u1_K5_37 ) , .A( u1_R3_24 ) , .Z( u1_u4_X_37 ) );
  XOR2_X1 u1_u4_U2 (.B( u1_K5_8 ) , .A( u1_R3_5 ) , .Z( u1_u4_X_8 ) );
  XOR2_X1 u1_u4_U20 (.B( u1_K5_36 ) , .A( u1_R3_25 ) , .Z( u1_u4_X_36 ) );
  XOR2_X1 u1_u4_U21 (.B( u1_K5_35 ) , .A( u1_R3_24 ) , .Z( u1_u4_X_35 ) );
  XOR2_X1 u1_u4_U22 (.B( u1_K5_34 ) , .A( u1_R3_23 ) , .Z( u1_u4_X_34 ) );
  XOR2_X1 u1_u4_U23 (.B( u1_K5_33 ) , .A( u1_R3_22 ) , .Z( u1_u4_X_33 ) );
  XOR2_X1 u1_u4_U24 (.B( u1_K5_32 ) , .A( u1_R3_21 ) , .Z( u1_u4_X_32 ) );
  XOR2_X1 u1_u4_U25 (.B( u1_K5_31 ) , .A( u1_R3_20 ) , .Z( u1_u4_X_31 ) );
  XOR2_X1 u1_u4_U26 (.B( u1_K5_30 ) , .A( u1_R3_21 ) , .Z( u1_u4_X_30 ) );
  XOR2_X1 u1_u4_U27 (.B( u1_K5_2 ) , .A( u1_R3_1 ) , .Z( u1_u4_X_2 ) );
  XOR2_X1 u1_u4_U28 (.B( u1_K5_29 ) , .A( u1_R3_20 ) , .Z( u1_u4_X_29 ) );
  XOR2_X1 u1_u4_U31 (.B( u1_K5_26 ) , .A( u1_R3_17 ) , .Z( u1_u4_X_26 ) );
  XOR2_X1 u1_u4_U32 (.B( u1_K5_25 ) , .A( u1_R3_16 ) , .Z( u1_u4_X_25 ) );
  XOR2_X1 u1_u4_U33 (.B( u1_K5_24 ) , .A( u1_R3_17 ) , .Z( u1_u4_X_24 ) );
  XOR2_X1 u1_u4_U34 (.B( u1_K5_23 ) , .A( u1_R3_16 ) , .Z( u1_u4_X_23 ) );
  XOR2_X1 u1_u4_U37 (.B( u1_K5_20 ) , .A( u1_R3_13 ) , .Z( u1_u4_X_20 ) );
  XOR2_X1 u1_u4_U38 (.B( u1_K5_1 ) , .A( u1_R3_32 ) , .Z( u1_u4_X_1 ) );
  XOR2_X1 u1_u4_U39 (.B( u1_K5_19 ) , .A( u1_R3_12 ) , .Z( u1_u4_X_19 ) );
  XOR2_X1 u1_u4_U4 (.B( u1_K5_6 ) , .A( u1_R3_5 ) , .Z( u1_u4_X_6 ) );
  XOR2_X1 u1_u4_U40 (.B( u1_K5_18 ) , .A( u1_R3_13 ) , .Z( u1_u4_X_18 ) );
  XOR2_X1 u1_u4_U41 (.B( u1_K5_17 ) , .A( u1_R3_12 ) , .Z( u1_u4_X_17 ) );
  XOR2_X1 u1_u4_U44 (.B( u1_K5_14 ) , .A( u1_R3_9 ) , .Z( u1_u4_X_14 ) );
  XOR2_X1 u1_u4_U45 (.B( u1_K5_13 ) , .A( u1_R3_8 ) , .Z( u1_u4_X_13 ) );
  XOR2_X1 u1_u4_U46 (.B( u1_K5_12 ) , .A( u1_R3_9 ) , .Z( u1_u4_X_12 ) );
  XOR2_X1 u1_u4_U47 (.B( u1_K5_11 ) , .A( u1_R3_8 ) , .Z( u1_u4_X_11 ) );
  XOR2_X1 u1_u4_U7 (.B( u1_K5_48 ) , .A( u1_R3_1 ) , .Z( u1_u4_X_48 ) );
  XOR2_X1 u1_u4_U8 (.B( u1_K5_47 ) , .A( u1_R3_32 ) , .Z( u1_u4_X_47 ) );
  XOR2_X1 u1_u4_U9 (.B( u1_K5_46 ) , .A( u1_R3_31 ) , .Z( u1_u4_X_46 ) );
  NOR2_X1 u1_u4_u5_U10 (.ZN( u1_u4_u5_n135 ) , .A1( u1_u4_u5_n173 ) , .A2( u1_u4_u5_n176 ) );
  NOR3_X1 u1_u4_u5_U100 (.A3( u1_u4_u5_n141 ) , .A1( u1_u4_u5_n142 ) , .ZN( u1_u4_u5_n143 ) , .A2( u1_u4_u5_n191 ) );
  NAND4_X1 u1_u4_u5_U101 (.ZN( u1_out4_4 ) , .A4( u1_u4_u5_n112 ) , .A2( u1_u4_u5_n113 ) , .A1( u1_u4_u5_n114 ) , .A3( u1_u4_u5_n195 ) );
  AOI211_X1 u1_u4_u5_U102 (.A( u1_u4_u5_n110 ) , .C1( u1_u4_u5_n111 ) , .ZN( u1_u4_u5_n112 ) , .B( u1_u4_u5_n118 ) , .C2( u1_u4_u5_n177 ) );
  INV_X1 u1_u4_u5_U103 (.A( u1_u4_u5_n102 ) , .ZN( u1_u4_u5_n195 ) );
  NAND3_X1 u1_u4_u5_U104 (.A2( u1_u4_u5_n154 ) , .A3( u1_u4_u5_n158 ) , .A1( u1_u4_u5_n161 ) , .ZN( u1_u4_u5_n99 ) );
  INV_X1 u1_u4_u5_U11 (.A( u1_u4_u5_n121 ) , .ZN( u1_u4_u5_n177 ) );
  NOR2_X1 u1_u4_u5_U12 (.ZN( u1_u4_u5_n160 ) , .A2( u1_u4_u5_n173 ) , .A1( u1_u4_u5_n177 ) );
  INV_X1 u1_u4_u5_U13 (.A( u1_u4_u5_n150 ) , .ZN( u1_u4_u5_n174 ) );
  AOI21_X1 u1_u4_u5_U14 (.A( u1_u4_u5_n160 ) , .B2( u1_u4_u5_n161 ) , .ZN( u1_u4_u5_n162 ) , .B1( u1_u4_u5_n192 ) );
  INV_X1 u1_u4_u5_U15 (.A( u1_u4_u5_n159 ) , .ZN( u1_u4_u5_n192 ) );
  AOI21_X1 u1_u4_u5_U16 (.A( u1_u4_u5_n156 ) , .B2( u1_u4_u5_n157 ) , .B1( u1_u4_u5_n158 ) , .ZN( u1_u4_u5_n163 ) );
  AOI21_X1 u1_u4_u5_U17 (.B2( u1_u4_u5_n139 ) , .B1( u1_u4_u5_n140 ) , .ZN( u1_u4_u5_n141 ) , .A( u1_u4_u5_n150 ) );
  OAI21_X1 u1_u4_u5_U18 (.A( u1_u4_u5_n133 ) , .B2( u1_u4_u5_n134 ) , .B1( u1_u4_u5_n135 ) , .ZN( u1_u4_u5_n142 ) );
  OAI21_X1 u1_u4_u5_U19 (.ZN( u1_u4_u5_n133 ) , .B2( u1_u4_u5_n147 ) , .A( u1_u4_u5_n173 ) , .B1( u1_u4_u5_n188 ) );
  NAND2_X1 u1_u4_u5_U20 (.A2( u1_u4_u5_n119 ) , .A1( u1_u4_u5_n123 ) , .ZN( u1_u4_u5_n137 ) );
  INV_X1 u1_u4_u5_U21 (.A( u1_u4_u5_n155 ) , .ZN( u1_u4_u5_n194 ) );
  NAND2_X1 u1_u4_u5_U22 (.A1( u1_u4_u5_n121 ) , .ZN( u1_u4_u5_n132 ) , .A2( u1_u4_u5_n172 ) );
  NAND2_X1 u1_u4_u5_U23 (.A2( u1_u4_u5_n122 ) , .ZN( u1_u4_u5_n136 ) , .A1( u1_u4_u5_n154 ) );
  NAND2_X1 u1_u4_u5_U24 (.A2( u1_u4_u5_n119 ) , .A1( u1_u4_u5_n120 ) , .ZN( u1_u4_u5_n159 ) );
  INV_X1 u1_u4_u5_U25 (.A( u1_u4_u5_n156 ) , .ZN( u1_u4_u5_n175 ) );
  INV_X1 u1_u4_u5_U26 (.A( u1_u4_u5_n158 ) , .ZN( u1_u4_u5_n188 ) );
  INV_X1 u1_u4_u5_U27 (.A( u1_u4_u5_n152 ) , .ZN( u1_u4_u5_n179 ) );
  INV_X1 u1_u4_u5_U28 (.A( u1_u4_u5_n140 ) , .ZN( u1_u4_u5_n182 ) );
  INV_X1 u1_u4_u5_U29 (.A( u1_u4_u5_n151 ) , .ZN( u1_u4_u5_n183 ) );
  NOR2_X1 u1_u4_u5_U3 (.ZN( u1_u4_u5_n134 ) , .A1( u1_u4_u5_n183 ) , .A2( u1_u4_u5_n190 ) );
  INV_X1 u1_u4_u5_U30 (.A( u1_u4_u5_n123 ) , .ZN( u1_u4_u5_n185 ) );
  INV_X1 u1_u4_u5_U31 (.A( u1_u4_u5_n161 ) , .ZN( u1_u4_u5_n184 ) );
  INV_X1 u1_u4_u5_U32 (.A( u1_u4_u5_n139 ) , .ZN( u1_u4_u5_n189 ) );
  INV_X1 u1_u4_u5_U33 (.A( u1_u4_u5_n157 ) , .ZN( u1_u4_u5_n190 ) );
  INV_X1 u1_u4_u5_U34 (.A( u1_u4_u5_n120 ) , .ZN( u1_u4_u5_n193 ) );
  NAND2_X1 u1_u4_u5_U35 (.ZN( u1_u4_u5_n111 ) , .A1( u1_u4_u5_n140 ) , .A2( u1_u4_u5_n155 ) );
  INV_X1 u1_u4_u5_U36 (.A( u1_u4_u5_n117 ) , .ZN( u1_u4_u5_n196 ) );
  OAI221_X1 u1_u4_u5_U37 (.A( u1_u4_u5_n116 ) , .ZN( u1_u4_u5_n117 ) , .B2( u1_u4_u5_n119 ) , .C1( u1_u4_u5_n153 ) , .C2( u1_u4_u5_n158 ) , .B1( u1_u4_u5_n172 ) );
  AOI222_X1 u1_u4_u5_U38 (.ZN( u1_u4_u5_n116 ) , .B2( u1_u4_u5_n145 ) , .C1( u1_u4_u5_n148 ) , .A2( u1_u4_u5_n174 ) , .C2( u1_u4_u5_n177 ) , .B1( u1_u4_u5_n187 ) , .A1( u1_u4_u5_n193 ) );
  INV_X1 u1_u4_u5_U39 (.A( u1_u4_u5_n115 ) , .ZN( u1_u4_u5_n187 ) );
  INV_X1 u1_u4_u5_U4 (.A( u1_u4_u5_n138 ) , .ZN( u1_u4_u5_n191 ) );
  NOR2_X1 u1_u4_u5_U40 (.ZN( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n170 ) , .A2( u1_u4_u5_n180 ) );
  OAI221_X1 u1_u4_u5_U41 (.A( u1_u4_u5_n101 ) , .ZN( u1_u4_u5_n102 ) , .C2( u1_u4_u5_n115 ) , .C1( u1_u4_u5_n126 ) , .B1( u1_u4_u5_n134 ) , .B2( u1_u4_u5_n160 ) );
  OAI21_X1 u1_u4_u5_U42 (.ZN( u1_u4_u5_n101 ) , .B1( u1_u4_u5_n137 ) , .A( u1_u4_u5_n146 ) , .B2( u1_u4_u5_n147 ) );
  AOI22_X1 u1_u4_u5_U43 (.B2( u1_u4_u5_n131 ) , .A2( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n169 ) , .B1( u1_u4_u5_n174 ) , .A1( u1_u4_u5_n185 ) );
  NOR2_X1 u1_u4_u5_U44 (.A1( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n150 ) , .A2( u1_u4_u5_n173 ) );
  AOI21_X1 u1_u4_u5_U45 (.A( u1_u4_u5_n118 ) , .B2( u1_u4_u5_n145 ) , .ZN( u1_u4_u5_n168 ) , .B1( u1_u4_u5_n186 ) );
  INV_X1 u1_u4_u5_U46 (.A( u1_u4_u5_n122 ) , .ZN( u1_u4_u5_n186 ) );
  NOR2_X1 u1_u4_u5_U47 (.A1( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n152 ) , .A2( u1_u4_u5_n176 ) );
  NOR2_X1 u1_u4_u5_U48 (.A1( u1_u4_u5_n115 ) , .ZN( u1_u4_u5_n118 ) , .A2( u1_u4_u5_n153 ) );
  NOR2_X1 u1_u4_u5_U49 (.A2( u1_u4_u5_n145 ) , .ZN( u1_u4_u5_n156 ) , .A1( u1_u4_u5_n174 ) );
  OAI21_X1 u1_u4_u5_U5 (.B2( u1_u4_u5_n136 ) , .B1( u1_u4_u5_n137 ) , .ZN( u1_u4_u5_n138 ) , .A( u1_u4_u5_n177 ) );
  NOR2_X1 u1_u4_u5_U50 (.ZN( u1_u4_u5_n121 ) , .A2( u1_u4_u5_n145 ) , .A1( u1_u4_u5_n176 ) );
  AOI22_X1 u1_u4_u5_U51 (.ZN( u1_u4_u5_n114 ) , .A2( u1_u4_u5_n137 ) , .A1( u1_u4_u5_n145 ) , .B2( u1_u4_u5_n175 ) , .B1( u1_u4_u5_n193 ) );
  OAI211_X1 u1_u4_u5_U52 (.B( u1_u4_u5_n124 ) , .A( u1_u4_u5_n125 ) , .C2( u1_u4_u5_n126 ) , .C1( u1_u4_u5_n127 ) , .ZN( u1_u4_u5_n128 ) );
  NOR3_X1 u1_u4_u5_U53 (.ZN( u1_u4_u5_n127 ) , .A1( u1_u4_u5_n136 ) , .A3( u1_u4_u5_n148 ) , .A2( u1_u4_u5_n182 ) );
  OAI21_X1 u1_u4_u5_U54 (.ZN( u1_u4_u5_n124 ) , .A( u1_u4_u5_n177 ) , .B2( u1_u4_u5_n183 ) , .B1( u1_u4_u5_n189 ) );
  OAI21_X1 u1_u4_u5_U55 (.ZN( u1_u4_u5_n125 ) , .A( u1_u4_u5_n174 ) , .B2( u1_u4_u5_n185 ) , .B1( u1_u4_u5_n190 ) );
  AOI21_X1 u1_u4_u5_U56 (.A( u1_u4_u5_n153 ) , .B2( u1_u4_u5_n154 ) , .B1( u1_u4_u5_n155 ) , .ZN( u1_u4_u5_n164 ) );
  AOI21_X1 u1_u4_u5_U57 (.ZN( u1_u4_u5_n110 ) , .B1( u1_u4_u5_n122 ) , .B2( u1_u4_u5_n139 ) , .A( u1_u4_u5_n153 ) );
  INV_X1 u1_u4_u5_U58 (.A( u1_u4_u5_n153 ) , .ZN( u1_u4_u5_n176 ) );
  INV_X1 u1_u4_u5_U59 (.A( u1_u4_u5_n126 ) , .ZN( u1_u4_u5_n173 ) );
  AOI222_X1 u1_u4_u5_U6 (.ZN( u1_u4_u5_n113 ) , .A1( u1_u4_u5_n131 ) , .C1( u1_u4_u5_n148 ) , .B2( u1_u4_u5_n174 ) , .C2( u1_u4_u5_n178 ) , .A2( u1_u4_u5_n179 ) , .B1( u1_u4_u5_n99 ) );
  AND2_X1 u1_u4_u5_U60 (.A2( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n107 ) , .ZN( u1_u4_u5_n147 ) );
  AND2_X1 u1_u4_u5_U61 (.A2( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n108 ) , .ZN( u1_u4_u5_n148 ) );
  NAND2_X1 u1_u4_u5_U62 (.A1( u1_u4_u5_n105 ) , .A2( u1_u4_u5_n106 ) , .ZN( u1_u4_u5_n158 ) );
  NAND2_X1 u1_u4_u5_U63 (.A2( u1_u4_u5_n108 ) , .A1( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n139 ) );
  NAND2_X1 u1_u4_u5_U64 (.A1( u1_u4_u5_n106 ) , .A2( u1_u4_u5_n108 ) , .ZN( u1_u4_u5_n119 ) );
  NAND2_X1 u1_u4_u5_U65 (.A2( u1_u4_u5_n103 ) , .A1( u1_u4_u5_n105 ) , .ZN( u1_u4_u5_n140 ) );
  NAND2_X1 u1_u4_u5_U66 (.A2( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n105 ) , .ZN( u1_u4_u5_n155 ) );
  NAND2_X1 u1_u4_u5_U67 (.A2( u1_u4_u5_n106 ) , .A1( u1_u4_u5_n107 ) , .ZN( u1_u4_u5_n122 ) );
  NAND2_X1 u1_u4_u5_U68 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n106 ) , .ZN( u1_u4_u5_n115 ) );
  NAND2_X1 u1_u4_u5_U69 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n103 ) , .ZN( u1_u4_u5_n161 ) );
  INV_X1 u1_u4_u5_U7 (.A( u1_u4_u5_n135 ) , .ZN( u1_u4_u5_n178 ) );
  NAND2_X1 u1_u4_u5_U70 (.A1( u1_u4_u5_n105 ) , .A2( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n154 ) );
  INV_X1 u1_u4_u5_U71 (.A( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n172 ) );
  NAND2_X1 u1_u4_u5_U72 (.A1( u1_u4_u5_n103 ) , .A2( u1_u4_u5_n108 ) , .ZN( u1_u4_u5_n123 ) );
  NAND2_X1 u1_u4_u5_U73 (.A2( u1_u4_u5_n103 ) , .A1( u1_u4_u5_n107 ) , .ZN( u1_u4_u5_n151 ) );
  NAND2_X1 u1_u4_u5_U74 (.A2( u1_u4_u5_n107 ) , .A1( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n120 ) );
  NAND2_X1 u1_u4_u5_U75 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n109 ) , .ZN( u1_u4_u5_n157 ) );
  AND2_X1 u1_u4_u5_U76 (.A2( u1_u4_u5_n100 ) , .A1( u1_u4_u5_n104 ) , .ZN( u1_u4_u5_n131 ) );
  NOR2_X1 u1_u4_u5_U77 (.A2( u1_u4_X_34 ) , .A1( u1_u4_X_35 ) , .ZN( u1_u4_u5_n145 ) );
  NOR2_X1 u1_u4_u5_U78 (.A2( u1_u4_X_34 ) , .ZN( u1_u4_u5_n146 ) , .A1( u1_u4_u5_n171 ) );
  NOR2_X1 u1_u4_u5_U79 (.A2( u1_u4_X_31 ) , .A1( u1_u4_X_32 ) , .ZN( u1_u4_u5_n103 ) );
  OAI22_X1 u1_u4_u5_U8 (.B2( u1_u4_u5_n149 ) , .B1( u1_u4_u5_n150 ) , .A2( u1_u4_u5_n151 ) , .A1( u1_u4_u5_n152 ) , .ZN( u1_u4_u5_n165 ) );
  NOR2_X1 u1_u4_u5_U80 (.A2( u1_u4_X_36 ) , .ZN( u1_u4_u5_n105 ) , .A1( u1_u4_u5_n180 ) );
  NOR2_X1 u1_u4_u5_U81 (.A2( u1_u4_X_33 ) , .ZN( u1_u4_u5_n108 ) , .A1( u1_u4_u5_n170 ) );
  NOR2_X1 u1_u4_u5_U82 (.A2( u1_u4_X_33 ) , .A1( u1_u4_X_36 ) , .ZN( u1_u4_u5_n107 ) );
  NOR2_X1 u1_u4_u5_U83 (.A2( u1_u4_X_31 ) , .ZN( u1_u4_u5_n104 ) , .A1( u1_u4_u5_n181 ) );
  NAND2_X1 u1_u4_u5_U84 (.A2( u1_u4_X_34 ) , .A1( u1_u4_X_35 ) , .ZN( u1_u4_u5_n153 ) );
  NAND2_X1 u1_u4_u5_U85 (.A1( u1_u4_X_34 ) , .ZN( u1_u4_u5_n126 ) , .A2( u1_u4_u5_n171 ) );
  AND2_X1 u1_u4_u5_U86 (.A1( u1_u4_X_31 ) , .A2( u1_u4_X_32 ) , .ZN( u1_u4_u5_n106 ) );
  AND2_X1 u1_u4_u5_U87 (.A1( u1_u4_X_31 ) , .ZN( u1_u4_u5_n109 ) , .A2( u1_u4_u5_n181 ) );
  INV_X1 u1_u4_u5_U88 (.A( u1_u4_X_33 ) , .ZN( u1_u4_u5_n180 ) );
  INV_X1 u1_u4_u5_U89 (.A( u1_u4_X_35 ) , .ZN( u1_u4_u5_n171 ) );
  NOR3_X1 u1_u4_u5_U9 (.A2( u1_u4_u5_n147 ) , .A1( u1_u4_u5_n148 ) , .ZN( u1_u4_u5_n149 ) , .A3( u1_u4_u5_n194 ) );
  INV_X1 u1_u4_u5_U90 (.A( u1_u4_X_36 ) , .ZN( u1_u4_u5_n170 ) );
  INV_X1 u1_u4_u5_U91 (.A( u1_u4_X_32 ) , .ZN( u1_u4_u5_n181 ) );
  NAND4_X1 u1_u4_u5_U92 (.ZN( u1_out4_29 ) , .A4( u1_u4_u5_n129 ) , .A3( u1_u4_u5_n130 ) , .A2( u1_u4_u5_n168 ) , .A1( u1_u4_u5_n196 ) );
  AOI221_X1 u1_u4_u5_U93 (.A( u1_u4_u5_n128 ) , .ZN( u1_u4_u5_n129 ) , .C2( u1_u4_u5_n132 ) , .B2( u1_u4_u5_n159 ) , .B1( u1_u4_u5_n176 ) , .C1( u1_u4_u5_n184 ) );
  AOI222_X1 u1_u4_u5_U94 (.ZN( u1_u4_u5_n130 ) , .A2( u1_u4_u5_n146 ) , .B1( u1_u4_u5_n147 ) , .C2( u1_u4_u5_n175 ) , .B2( u1_u4_u5_n179 ) , .A1( u1_u4_u5_n188 ) , .C1( u1_u4_u5_n194 ) );
  NAND4_X1 u1_u4_u5_U95 (.ZN( u1_out4_19 ) , .A4( u1_u4_u5_n166 ) , .A3( u1_u4_u5_n167 ) , .A2( u1_u4_u5_n168 ) , .A1( u1_u4_u5_n169 ) );
  AOI22_X1 u1_u4_u5_U96 (.B2( u1_u4_u5_n145 ) , .A2( u1_u4_u5_n146 ) , .ZN( u1_u4_u5_n167 ) , .B1( u1_u4_u5_n182 ) , .A1( u1_u4_u5_n189 ) );
  NOR4_X1 u1_u4_u5_U97 (.A4( u1_u4_u5_n162 ) , .A3( u1_u4_u5_n163 ) , .A2( u1_u4_u5_n164 ) , .A1( u1_u4_u5_n165 ) , .ZN( u1_u4_u5_n166 ) );
  NAND4_X1 u1_u4_u5_U98 (.ZN( u1_out4_11 ) , .A4( u1_u4_u5_n143 ) , .A3( u1_u4_u5_n144 ) , .A2( u1_u4_u5_n169 ) , .A1( u1_u4_u5_n196 ) );
  AOI22_X1 u1_u4_u5_U99 (.A2( u1_u4_u5_n132 ) , .ZN( u1_u4_u5_n144 ) , .B2( u1_u4_u5_n145 ) , .B1( u1_u4_u5_n184 ) , .A1( u1_u4_u5_n194 ) );
  AND3_X1 u1_u4_u7_U10 (.A3( u1_u4_u7_n110 ) , .A2( u1_u4_u7_n127 ) , .A1( u1_u4_u7_n132 ) , .ZN( u1_u4_u7_n92 ) );
  OAI21_X1 u1_u4_u7_U11 (.A( u1_u4_u7_n161 ) , .B1( u1_u4_u7_n168 ) , .B2( u1_u4_u7_n173 ) , .ZN( u1_u4_u7_n91 ) );
  AOI211_X1 u1_u4_u7_U12 (.A( u1_u4_u7_n117 ) , .ZN( u1_u4_u7_n118 ) , .C2( u1_u4_u7_n126 ) , .C1( u1_u4_u7_n177 ) , .B( u1_u4_u7_n180 ) );
  OAI22_X1 u1_u4_u7_U13 (.B1( u1_u4_u7_n115 ) , .ZN( u1_u4_u7_n117 ) , .A2( u1_u4_u7_n133 ) , .A1( u1_u4_u7_n137 ) , .B2( u1_u4_u7_n162 ) );
  INV_X1 u1_u4_u7_U14 (.A( u1_u4_u7_n116 ) , .ZN( u1_u4_u7_n180 ) );
  NOR3_X1 u1_u4_u7_U15 (.ZN( u1_u4_u7_n115 ) , .A3( u1_u4_u7_n145 ) , .A2( u1_u4_u7_n168 ) , .A1( u1_u4_u7_n169 ) );
  NOR3_X1 u1_u4_u7_U16 (.A2( u1_u4_u7_n134 ) , .A1( u1_u4_u7_n135 ) , .ZN( u1_u4_u7_n136 ) , .A3( u1_u4_u7_n171 ) );
  NOR2_X1 u1_u4_u7_U17 (.A1( u1_u4_u7_n130 ) , .A2( u1_u4_u7_n134 ) , .ZN( u1_u4_u7_n153 ) );
  NOR2_X1 u1_u4_u7_U18 (.ZN( u1_u4_u7_n111 ) , .A2( u1_u4_u7_n134 ) , .A1( u1_u4_u7_n169 ) );
  AOI21_X1 u1_u4_u7_U19 (.ZN( u1_u4_u7_n104 ) , .B2( u1_u4_u7_n112 ) , .B1( u1_u4_u7_n127 ) , .A( u1_u4_u7_n164 ) );
  AOI21_X1 u1_u4_u7_U20 (.ZN( u1_u4_u7_n106 ) , .B1( u1_u4_u7_n133 ) , .B2( u1_u4_u7_n146 ) , .A( u1_u4_u7_n162 ) );
  AOI21_X1 u1_u4_u7_U21 (.A( u1_u4_u7_n101 ) , .ZN( u1_u4_u7_n107 ) , .B2( u1_u4_u7_n128 ) , .B1( u1_u4_u7_n175 ) );
  INV_X1 u1_u4_u7_U22 (.A( u1_u4_u7_n101 ) , .ZN( u1_u4_u7_n165 ) );
  INV_X1 u1_u4_u7_U23 (.A( u1_u4_u7_n138 ) , .ZN( u1_u4_u7_n171 ) );
  INV_X1 u1_u4_u7_U24 (.A( u1_u4_u7_n131 ) , .ZN( u1_u4_u7_n177 ) );
  INV_X1 u1_u4_u7_U25 (.A( u1_u4_u7_n110 ) , .ZN( u1_u4_u7_n174 ) );
  NAND2_X1 u1_u4_u7_U26 (.A1( u1_u4_u7_n129 ) , .A2( u1_u4_u7_n132 ) , .ZN( u1_u4_u7_n149 ) );
  NAND2_X1 u1_u4_u7_U27 (.A1( u1_u4_u7_n113 ) , .A2( u1_u4_u7_n124 ) , .ZN( u1_u4_u7_n130 ) );
  INV_X1 u1_u4_u7_U28 (.A( u1_u4_u7_n128 ) , .ZN( u1_u4_u7_n168 ) );
  INV_X1 u1_u4_u7_U29 (.A( u1_u4_u7_n148 ) , .ZN( u1_u4_u7_n169 ) );
  INV_X1 u1_u4_u7_U3 (.A( u1_u4_u7_n149 ) , .ZN( u1_u4_u7_n175 ) );
  INV_X1 u1_u4_u7_U30 (.A( u1_u4_u7_n112 ) , .ZN( u1_u4_u7_n173 ) );
  INV_X1 u1_u4_u7_U31 (.A( u1_u4_u7_n127 ) , .ZN( u1_u4_u7_n179 ) );
  NOR2_X1 u1_u4_u7_U32 (.ZN( u1_u4_u7_n101 ) , .A2( u1_u4_u7_n150 ) , .A1( u1_u4_u7_n156 ) );
  AOI211_X1 u1_u4_u7_U33 (.B( u1_u4_u7_n154 ) , .A( u1_u4_u7_n155 ) , .C1( u1_u4_u7_n156 ) , .ZN( u1_u4_u7_n157 ) , .C2( u1_u4_u7_n172 ) );
  INV_X1 u1_u4_u7_U34 (.A( u1_u4_u7_n153 ) , .ZN( u1_u4_u7_n172 ) );
  AOI211_X1 u1_u4_u7_U35 (.B( u1_u4_u7_n139 ) , .A( u1_u4_u7_n140 ) , .C2( u1_u4_u7_n141 ) , .ZN( u1_u4_u7_n142 ) , .C1( u1_u4_u7_n156 ) );
  NAND4_X1 u1_u4_u7_U36 (.A3( u1_u4_u7_n127 ) , .A2( u1_u4_u7_n128 ) , .A1( u1_u4_u7_n129 ) , .ZN( u1_u4_u7_n141 ) , .A4( u1_u4_u7_n147 ) );
  AOI21_X1 u1_u4_u7_U37 (.A( u1_u4_u7_n137 ) , .B1( u1_u4_u7_n138 ) , .ZN( u1_u4_u7_n139 ) , .B2( u1_u4_u7_n146 ) );
  OAI22_X1 u1_u4_u7_U38 (.B1( u1_u4_u7_n136 ) , .ZN( u1_u4_u7_n140 ) , .A1( u1_u4_u7_n153 ) , .B2( u1_u4_u7_n162 ) , .A2( u1_u4_u7_n164 ) );
  INV_X1 u1_u4_u7_U39 (.A( u1_u4_u7_n125 ) , .ZN( u1_u4_u7_n161 ) );
  INV_X1 u1_u4_u7_U4 (.A( u1_u4_u7_n154 ) , .ZN( u1_u4_u7_n178 ) );
  AOI21_X1 u1_u4_u7_U40 (.ZN( u1_u4_u7_n123 ) , .B1( u1_u4_u7_n165 ) , .B2( u1_u4_u7_n177 ) , .A( u1_u4_u7_n97 ) );
  AOI21_X1 u1_u4_u7_U41 (.B2( u1_u4_u7_n113 ) , .B1( u1_u4_u7_n124 ) , .A( u1_u4_u7_n125 ) , .ZN( u1_u4_u7_n97 ) );
  INV_X1 u1_u4_u7_U42 (.A( u1_u4_u7_n152 ) , .ZN( u1_u4_u7_n162 ) );
  AOI22_X1 u1_u4_u7_U43 (.A2( u1_u4_u7_n114 ) , .ZN( u1_u4_u7_n119 ) , .B1( u1_u4_u7_n130 ) , .A1( u1_u4_u7_n156 ) , .B2( u1_u4_u7_n165 ) );
  NAND2_X1 u1_u4_u7_U44 (.A2( u1_u4_u7_n112 ) , .ZN( u1_u4_u7_n114 ) , .A1( u1_u4_u7_n175 ) );
  AOI22_X1 u1_u4_u7_U45 (.B2( u1_u4_u7_n149 ) , .B1( u1_u4_u7_n150 ) , .A2( u1_u4_u7_n151 ) , .A1( u1_u4_u7_n152 ) , .ZN( u1_u4_u7_n158 ) );
  NOR2_X1 u1_u4_u7_U46 (.ZN( u1_u4_u7_n137 ) , .A1( u1_u4_u7_n150 ) , .A2( u1_u4_u7_n161 ) );
  AND2_X1 u1_u4_u7_U47 (.ZN( u1_u4_u7_n145 ) , .A2( u1_u4_u7_n98 ) , .A1( u1_u4_u7_n99 ) );
  AOI21_X1 u1_u4_u7_U48 (.ZN( u1_u4_u7_n105 ) , .B2( u1_u4_u7_n110 ) , .A( u1_u4_u7_n125 ) , .B1( u1_u4_u7_n147 ) );
  NAND2_X1 u1_u4_u7_U49 (.ZN( u1_u4_u7_n146 ) , .A1( u1_u4_u7_n95 ) , .A2( u1_u4_u7_n98 ) );
  INV_X1 u1_u4_u7_U5 (.A( u1_u4_u7_n111 ) , .ZN( u1_u4_u7_n170 ) );
  NAND2_X1 u1_u4_u7_U50 (.A2( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n147 ) , .A1( u1_u4_u7_n93 ) );
  NAND2_X1 u1_u4_u7_U51 (.A1( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n127 ) , .A2( u1_u4_u7_n99 ) );
  NAND2_X1 u1_u4_u7_U52 (.A2( u1_u4_u7_n102 ) , .A1( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n133 ) );
  OR2_X1 u1_u4_u7_U53 (.ZN( u1_u4_u7_n126 ) , .A2( u1_u4_u7_n152 ) , .A1( u1_u4_u7_n156 ) );
  NAND2_X1 u1_u4_u7_U54 (.ZN( u1_u4_u7_n112 ) , .A2( u1_u4_u7_n96 ) , .A1( u1_u4_u7_n99 ) );
  NAND2_X1 u1_u4_u7_U55 (.A2( u1_u4_u7_n102 ) , .ZN( u1_u4_u7_n128 ) , .A1( u1_u4_u7_n98 ) );
  INV_X1 u1_u4_u7_U56 (.A( u1_u4_u7_n150 ) , .ZN( u1_u4_u7_n164 ) );
  AND2_X1 u1_u4_u7_U57 (.ZN( u1_u4_u7_n134 ) , .A1( u1_u4_u7_n93 ) , .A2( u1_u4_u7_n98 ) );
  NAND2_X1 u1_u4_u7_U58 (.ZN( u1_u4_u7_n110 ) , .A1( u1_u4_u7_n95 ) , .A2( u1_u4_u7_n96 ) );
  NAND2_X1 u1_u4_u7_U59 (.A2( u1_u4_u7_n102 ) , .ZN( u1_u4_u7_n124 ) , .A1( u1_u4_u7_n96 ) );
  AOI211_X1 u1_u4_u7_U6 (.ZN( u1_u4_u7_n116 ) , .A( u1_u4_u7_n155 ) , .C1( u1_u4_u7_n161 ) , .C2( u1_u4_u7_n171 ) , .B( u1_u4_u7_n94 ) );
  NAND2_X1 u1_u4_u7_U60 (.ZN( u1_u4_u7_n132 ) , .A1( u1_u4_u7_n93 ) , .A2( u1_u4_u7_n96 ) );
  NAND2_X1 u1_u4_u7_U61 (.A2( u1_u4_u7_n103 ) , .ZN( u1_u4_u7_n131 ) , .A1( u1_u4_u7_n95 ) );
  NOR2_X1 u1_u4_u7_U62 (.A2( u1_u4_X_47 ) , .ZN( u1_u4_u7_n150 ) , .A1( u1_u4_u7_n163 ) );
  NOR2_X1 u1_u4_u7_U63 (.A2( u1_u4_X_43 ) , .A1( u1_u4_X_44 ) , .ZN( u1_u4_u7_n103 ) );
  NOR2_X1 u1_u4_u7_U64 (.A2( u1_u4_X_48 ) , .A1( u1_u4_u7_n166 ) , .ZN( u1_u4_u7_n95 ) );
  NOR2_X1 u1_u4_u7_U65 (.A2( u1_u4_X_44 ) , .A1( u1_u4_u7_n167 ) , .ZN( u1_u4_u7_n98 ) );
  NOR2_X1 u1_u4_u7_U66 (.A2( u1_u4_X_45 ) , .A1( u1_u4_X_48 ) , .ZN( u1_u4_u7_n99 ) );
  NOR2_X1 u1_u4_u7_U67 (.A2( u1_u4_X_46 ) , .A1( u1_u4_X_47 ) , .ZN( u1_u4_u7_n152 ) );
  AND2_X1 u1_u4_u7_U68 (.A1( u1_u4_X_47 ) , .ZN( u1_u4_u7_n156 ) , .A2( u1_u4_u7_n163 ) );
  NAND2_X1 u1_u4_u7_U69 (.A2( u1_u4_X_46 ) , .A1( u1_u4_X_47 ) , .ZN( u1_u4_u7_n125 ) );
  OAI222_X1 u1_u4_u7_U7 (.C2( u1_u4_u7_n101 ) , .B2( u1_u4_u7_n111 ) , .A1( u1_u4_u7_n113 ) , .C1( u1_u4_u7_n146 ) , .A2( u1_u4_u7_n162 ) , .B1( u1_u4_u7_n164 ) , .ZN( u1_u4_u7_n94 ) );
  AND2_X1 u1_u4_u7_U70 (.A2( u1_u4_X_43 ) , .A1( u1_u4_X_44 ) , .ZN( u1_u4_u7_n96 ) );
  AND2_X1 u1_u4_u7_U71 (.A2( u1_u4_X_45 ) , .A1( u1_u4_X_48 ) , .ZN( u1_u4_u7_n102 ) );
  AND2_X1 u1_u4_u7_U72 (.A1( u1_u4_X_48 ) , .A2( u1_u4_u7_n166 ) , .ZN( u1_u4_u7_n93 ) );
  INV_X1 u1_u4_u7_U73 (.A( u1_u4_X_46 ) , .ZN( u1_u4_u7_n163 ) );
  AND2_X1 u1_u4_u7_U74 (.A1( u1_u4_X_44 ) , .ZN( u1_u4_u7_n100 ) , .A2( u1_u4_u7_n167 ) );
  INV_X1 u1_u4_u7_U75 (.A( u1_u4_X_45 ) , .ZN( u1_u4_u7_n166 ) );
  INV_X1 u1_u4_u7_U76 (.A( u1_u4_X_43 ) , .ZN( u1_u4_u7_n167 ) );
  NAND4_X1 u1_u4_u7_U77 (.ZN( u1_out4_5 ) , .A4( u1_u4_u7_n108 ) , .A3( u1_u4_u7_n109 ) , .A1( u1_u4_u7_n116 ) , .A2( u1_u4_u7_n123 ) );
  AOI22_X1 u1_u4_u7_U78 (.ZN( u1_u4_u7_n109 ) , .A2( u1_u4_u7_n126 ) , .B2( u1_u4_u7_n145 ) , .B1( u1_u4_u7_n156 ) , .A1( u1_u4_u7_n171 ) );
  NOR4_X1 u1_u4_u7_U79 (.A4( u1_u4_u7_n104 ) , .A3( u1_u4_u7_n105 ) , .A2( u1_u4_u7_n106 ) , .A1( u1_u4_u7_n107 ) , .ZN( u1_u4_u7_n108 ) );
  INV_X1 u1_u4_u7_U8 (.A( u1_u4_u7_n133 ) , .ZN( u1_u4_u7_n176 ) );
  NAND4_X1 u1_u4_u7_U80 (.ZN( u1_out4_27 ) , .A4( u1_u4_u7_n118 ) , .A3( u1_u4_u7_n119 ) , .A2( u1_u4_u7_n120 ) , .A1( u1_u4_u7_n121 ) );
  OAI21_X1 u1_u4_u7_U81 (.ZN( u1_u4_u7_n121 ) , .B2( u1_u4_u7_n145 ) , .A( u1_u4_u7_n150 ) , .B1( u1_u4_u7_n174 ) );
  OAI21_X1 u1_u4_u7_U82 (.ZN( u1_u4_u7_n120 ) , .A( u1_u4_u7_n161 ) , .B2( u1_u4_u7_n170 ) , .B1( u1_u4_u7_n179 ) );
  NAND4_X1 u1_u4_u7_U83 (.ZN( u1_out4_21 ) , .A4( u1_u4_u7_n157 ) , .A3( u1_u4_u7_n158 ) , .A2( u1_u4_u7_n159 ) , .A1( u1_u4_u7_n160 ) );
  OAI21_X1 u1_u4_u7_U84 (.B1( u1_u4_u7_n145 ) , .ZN( u1_u4_u7_n160 ) , .A( u1_u4_u7_n161 ) , .B2( u1_u4_u7_n177 ) );
  OAI21_X1 u1_u4_u7_U85 (.ZN( u1_u4_u7_n159 ) , .A( u1_u4_u7_n165 ) , .B2( u1_u4_u7_n171 ) , .B1( u1_u4_u7_n174 ) );
  NAND4_X1 u1_u4_u7_U86 (.ZN( u1_out4_15 ) , .A4( u1_u4_u7_n142 ) , .A3( u1_u4_u7_n143 ) , .A2( u1_u4_u7_n144 ) , .A1( u1_u4_u7_n178 ) );
  OR2_X1 u1_u4_u7_U87 (.A2( u1_u4_u7_n125 ) , .A1( u1_u4_u7_n129 ) , .ZN( u1_u4_u7_n144 ) );
  AOI22_X1 u1_u4_u7_U88 (.A2( u1_u4_u7_n126 ) , .ZN( u1_u4_u7_n143 ) , .B2( u1_u4_u7_n165 ) , .B1( u1_u4_u7_n173 ) , .A1( u1_u4_u7_n174 ) );
  NAND2_X1 u1_u4_u7_U89 (.A1( u1_u4_u7_n100 ) , .ZN( u1_u4_u7_n148 ) , .A2( u1_u4_u7_n95 ) );
  OAI221_X1 u1_u4_u7_U9 (.C1( u1_u4_u7_n101 ) , .C2( u1_u4_u7_n147 ) , .ZN( u1_u4_u7_n155 ) , .B2( u1_u4_u7_n162 ) , .A( u1_u4_u7_n91 ) , .B1( u1_u4_u7_n92 ) );
  NAND2_X1 u1_u4_u7_U90 (.A1( u1_u4_u7_n100 ) , .ZN( u1_u4_u7_n113 ) , .A2( u1_u4_u7_n93 ) );
  NAND2_X1 u1_u4_u7_U91 (.A1( u1_u4_u7_n100 ) , .ZN( u1_u4_u7_n138 ) , .A2( u1_u4_u7_n99 ) );
  NAND2_X1 u1_u4_u7_U92 (.A1( u1_u4_u7_n100 ) , .A2( u1_u4_u7_n102 ) , .ZN( u1_u4_u7_n129 ) );
  OAI211_X1 u1_u4_u7_U93 (.B( u1_u4_u7_n122 ) , .A( u1_u4_u7_n123 ) , .C2( u1_u4_u7_n124 ) , .ZN( u1_u4_u7_n154 ) , .C1( u1_u4_u7_n162 ) );
  AOI222_X1 u1_u4_u7_U94 (.ZN( u1_u4_u7_n122 ) , .C2( u1_u4_u7_n126 ) , .C1( u1_u4_u7_n145 ) , .B1( u1_u4_u7_n161 ) , .A2( u1_u4_u7_n165 ) , .B2( u1_u4_u7_n170 ) , .A1( u1_u4_u7_n176 ) );
  NAND3_X1 u1_u4_u7_U95 (.A3( u1_u4_u7_n146 ) , .A2( u1_u4_u7_n147 ) , .A1( u1_u4_u7_n148 ) , .ZN( u1_u4_u7_n151 ) );
  NAND3_X1 u1_u4_u7_U96 (.A3( u1_u4_u7_n131 ) , .A2( u1_u4_u7_n132 ) , .A1( u1_u4_u7_n133 ) , .ZN( u1_u4_u7_n135 ) );
  XOR2_X1 u1_u5_U11 (.B( u1_K6_44 ) , .A( u1_R4_29 ) , .Z( u1_u5_X_44 ) );
  XOR2_X1 u1_u5_U12 (.B( u1_K6_43 ) , .A( u1_R4_28 ) , .Z( u1_u5_X_43 ) );
  XOR2_X1 u1_u5_U13 (.B( u1_K6_42 ) , .A( u1_R4_29 ) , .Z( u1_u5_X_42 ) );
  XOR2_X1 u1_u5_U14 (.B( u1_K6_41 ) , .A( u1_R4_28 ) , .Z( u1_u5_X_41 ) );
  XOR2_X1 u1_u5_U15 (.B( u1_K6_40 ) , .A( u1_R4_27 ) , .Z( u1_u5_X_40 ) );
  XOR2_X1 u1_u5_U16 (.B( u1_K6_3 ) , .A( u1_R4_2 ) , .Z( u1_u5_X_3 ) );
  XOR2_X1 u1_u5_U17 (.B( u1_K6_39 ) , .A( u1_R4_26 ) , .Z( u1_u5_X_39 ) );
  XOR2_X1 u1_u5_U18 (.B( u1_K6_38 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_38 ) );
  XOR2_X1 u1_u5_U19 (.B( u1_K6_37 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_37 ) );
  XOR2_X1 u1_u5_U2 (.B( u1_K6_8 ) , .A( u1_R4_5 ) , .Z( u1_u5_X_8 ) );
  XOR2_X1 u1_u5_U20 (.B( u1_K6_36 ) , .A( u1_R4_25 ) , .Z( u1_u5_X_36 ) );
  XOR2_X1 u1_u5_U21 (.B( u1_K6_35 ) , .A( u1_R4_24 ) , .Z( u1_u5_X_35 ) );
  XOR2_X1 u1_u5_U24 (.B( u1_K6_32 ) , .A( u1_R4_21 ) , .Z( u1_u5_X_32 ) );
  XOR2_X1 u1_u5_U26 (.B( u1_K6_30 ) , .A( u1_R4_21 ) , .Z( u1_u5_X_30 ) );
  XOR2_X1 u1_u5_U27 (.B( u1_K6_2 ) , .A( u1_R4_1 ) , .Z( u1_u5_X_2 ) );
  XOR2_X1 u1_u5_U3 (.B( u1_K6_7 ) , .A( u1_R4_4 ) , .Z( u1_u5_X_7 ) );
  XOR2_X1 u1_u5_U31 (.B( u1_K6_26 ) , .A( u1_R4_17 ) , .Z( u1_u5_X_26 ) );
  XOR2_X1 u1_u5_U32 (.B( u1_K6_25 ) , .A( u1_R4_16 ) , .Z( u1_u5_X_25 ) );
  XOR2_X1 u1_u5_U33 (.B( u1_K6_24 ) , .A( u1_R4_17 ) , .Z( u1_u5_X_24 ) );
  XOR2_X1 u1_u5_U34 (.B( u1_K6_23 ) , .A( u1_R4_16 ) , .Z( u1_u5_X_23 ) );
  XOR2_X1 u1_u5_U35 (.B( u1_K6_22 ) , .A( u1_R4_15 ) , .Z( u1_u5_X_22 ) );
  XOR2_X1 u1_u5_U36 (.B( u1_K6_21 ) , .A( u1_R4_14 ) , .Z( u1_u5_X_21 ) );
  XOR2_X1 u1_u5_U37 (.B( u1_K6_20 ) , .A( u1_R4_13 ) , .Z( u1_u5_X_20 ) );
  XOR2_X1 u1_u5_U38 (.B( u1_K6_1 ) , .A( u1_R4_32 ) , .Z( u1_u5_X_1 ) );
  XOR2_X1 u1_u5_U39 (.B( u1_K6_19 ) , .A( u1_R4_12 ) , .Z( u1_u5_X_19 ) );
  XOR2_X1 u1_u5_U4 (.B( u1_K6_6 ) , .A( u1_R4_5 ) , .Z( u1_u5_X_6 ) );
  XOR2_X1 u1_u5_U40 (.B( u1_K6_18 ) , .A( u1_R4_13 ) , .Z( u1_u5_X_18 ) );
  XOR2_X1 u1_u5_U41 (.B( u1_K6_17 ) , .A( u1_R4_12 ) , .Z( u1_u5_X_17 ) );
  XOR2_X1 u1_u5_U42 (.B( u1_K6_16 ) , .A( u1_R4_11 ) , .Z( u1_u5_X_16 ) );
  XOR2_X1 u1_u5_U43 (.B( u1_K6_15 ) , .A( u1_R4_10 ) , .Z( u1_u5_X_15 ) );
  XOR2_X1 u1_u5_U44 (.B( u1_K6_14 ) , .A( u1_R4_9 ) , .Z( u1_u5_X_14 ) );
  XOR2_X1 u1_u5_U45 (.B( u1_K6_13 ) , .A( u1_R4_8 ) , .Z( u1_u5_X_13 ) );
  XOR2_X1 u1_u5_U46 (.B( u1_K6_12 ) , .A( u1_R4_9 ) , .Z( u1_u5_X_12 ) );
  XOR2_X1 u1_u5_U47 (.B( u1_K6_11 ) , .A( u1_R4_8 ) , .Z( u1_u5_X_11 ) );
  XOR2_X1 u1_u5_U5 (.B( u1_K6_5 ) , .A( u1_R4_4 ) , .Z( u1_u5_X_5 ) );
  XOR2_X1 u1_u5_U6 (.B( u1_K6_4 ) , .A( u1_R4_3 ) , .Z( u1_u5_X_4 ) );
  XOR2_X1 u1_u5_U7 (.B( u1_K6_48 ) , .A( u1_R4_1 ) , .Z( u1_u5_X_48 ) );
  XOR2_X1 u1_u5_U8 (.B( u1_K6_47 ) , .A( u1_R4_32 ) , .Z( u1_u5_X_47 ) );
  NAND2_X1 u1_u5_u0_U10 (.ZN( u1_u5_u0_n113 ) , .A1( u1_u5_u0_n139 ) , .A2( u1_u5_u0_n149 ) );
  AND3_X1 u1_u5_u0_U11 (.A2( u1_u5_u0_n112 ) , .ZN( u1_u5_u0_n127 ) , .A3( u1_u5_u0_n130 ) , .A1( u1_u5_u0_n148 ) );
  AND2_X1 u1_u5_u0_U12 (.ZN( u1_u5_u0_n107 ) , .A1( u1_u5_u0_n130 ) , .A2( u1_u5_u0_n140 ) );
  AND2_X1 u1_u5_u0_U13 (.A2( u1_u5_u0_n129 ) , .A1( u1_u5_u0_n130 ) , .ZN( u1_u5_u0_n151 ) );
  AND2_X1 u1_u5_u0_U14 (.A1( u1_u5_u0_n108 ) , .A2( u1_u5_u0_n125 ) , .ZN( u1_u5_u0_n145 ) );
  INV_X1 u1_u5_u0_U15 (.A( u1_u5_u0_n143 ) , .ZN( u1_u5_u0_n173 ) );
  NOR2_X1 u1_u5_u0_U16 (.A2( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n147 ) , .A1( u1_u5_u0_n160 ) );
  AOI21_X1 u1_u5_u0_U17 (.B1( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n132 ) , .A( u1_u5_u0_n165 ) , .B2( u1_u5_u0_n93 ) );
  INV_X1 u1_u5_u0_U18 (.A( u1_u5_u0_n142 ) , .ZN( u1_u5_u0_n165 ) );
  OAI22_X1 u1_u5_u0_U19 (.B1( u1_u5_u0_n131 ) , .A1( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n147 ) , .A2( u1_u5_u0_n90 ) , .ZN( u1_u5_u0_n91 ) );
  AND3_X1 u1_u5_u0_U20 (.A3( u1_u5_u0_n121 ) , .A2( u1_u5_u0_n125 ) , .A1( u1_u5_u0_n148 ) , .ZN( u1_u5_u0_n90 ) );
  OAI22_X1 u1_u5_u0_U21 (.B1( u1_u5_u0_n125 ) , .ZN( u1_u5_u0_n126 ) , .A1( u1_u5_u0_n138 ) , .A2( u1_u5_u0_n146 ) , .B2( u1_u5_u0_n147 ) );
  NOR2_X1 u1_u5_u0_U22 (.A1( u1_u5_u0_n163 ) , .A2( u1_u5_u0_n164 ) , .ZN( u1_u5_u0_n95 ) );
  INV_X1 u1_u5_u0_U23 (.A( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n161 ) );
  AOI22_X1 u1_u5_u0_U24 (.B2( u1_u5_u0_n109 ) , .A2( u1_u5_u0_n110 ) , .ZN( u1_u5_u0_n111 ) , .B1( u1_u5_u0_n118 ) , .A1( u1_u5_u0_n160 ) );
  NAND2_X1 u1_u5_u0_U25 (.A2( u1_u5_u0_n102 ) , .A1( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n149 ) );
  INV_X1 u1_u5_u0_U26 (.A( u1_u5_u0_n118 ) , .ZN( u1_u5_u0_n158 ) );
  NAND2_X1 u1_u5_u0_U27 (.A2( u1_u5_u0_n100 ) , .ZN( u1_u5_u0_n131 ) , .A1( u1_u5_u0_n92 ) );
  NAND2_X1 u1_u5_u0_U28 (.ZN( u1_u5_u0_n108 ) , .A1( u1_u5_u0_n92 ) , .A2( u1_u5_u0_n94 ) );
  AOI21_X1 u1_u5_u0_U29 (.ZN( u1_u5_u0_n104 ) , .B1( u1_u5_u0_n107 ) , .B2( u1_u5_u0_n141 ) , .A( u1_u5_u0_n144 ) );
  INV_X1 u1_u5_u0_U3 (.A( u1_u5_u0_n113 ) , .ZN( u1_u5_u0_n166 ) );
  AOI21_X1 u1_u5_u0_U30 (.B1( u1_u5_u0_n127 ) , .B2( u1_u5_u0_n129 ) , .A( u1_u5_u0_n138 ) , .ZN( u1_u5_u0_n96 ) );
  NAND2_X1 u1_u5_u0_U31 (.A2( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n114 ) , .A1( u1_u5_u0_n92 ) );
  AOI21_X1 u1_u5_u0_U32 (.ZN( u1_u5_u0_n116 ) , .B2( u1_u5_u0_n142 ) , .A( u1_u5_u0_n144 ) , .B1( u1_u5_u0_n166 ) );
  NOR2_X1 u1_u5_u0_U33 (.A1( u1_u5_u0_n120 ) , .ZN( u1_u5_u0_n143 ) , .A2( u1_u5_u0_n167 ) );
  OAI221_X1 u1_u5_u0_U34 (.C1( u1_u5_u0_n112 ) , .ZN( u1_u5_u0_n120 ) , .B1( u1_u5_u0_n138 ) , .B2( u1_u5_u0_n141 ) , .C2( u1_u5_u0_n147 ) , .A( u1_u5_u0_n172 ) );
  AOI211_X1 u1_u5_u0_U35 (.B( u1_u5_u0_n115 ) , .A( u1_u5_u0_n116 ) , .C2( u1_u5_u0_n117 ) , .C1( u1_u5_u0_n118 ) , .ZN( u1_u5_u0_n119 ) );
  NAND2_X1 u1_u5_u0_U36 (.A2( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n140 ) , .A1( u1_u5_u0_n94 ) );
  NAND2_X1 u1_u5_u0_U37 (.A1( u1_u5_u0_n100 ) , .A2( u1_u5_u0_n103 ) , .ZN( u1_u5_u0_n125 ) );
  NAND2_X1 u1_u5_u0_U38 (.A1( u1_u5_u0_n101 ) , .A2( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n150 ) );
  INV_X1 u1_u5_u0_U39 (.A( u1_u5_u0_n138 ) , .ZN( u1_u5_u0_n160 ) );
  AOI21_X1 u1_u5_u0_U4 (.B1( u1_u5_u0_n114 ) , .ZN( u1_u5_u0_n115 ) , .B2( u1_u5_u0_n129 ) , .A( u1_u5_u0_n161 ) );
  NAND2_X1 u1_u5_u0_U40 (.A2( u1_u5_u0_n100 ) , .A1( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n139 ) );
  NAND2_X1 u1_u5_u0_U41 (.ZN( u1_u5_u0_n112 ) , .A2( u1_u5_u0_n92 ) , .A1( u1_u5_u0_n93 ) );
  NAND2_X1 u1_u5_u0_U42 (.A1( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n130 ) , .A2( u1_u5_u0_n94 ) );
  INV_X1 u1_u5_u0_U43 (.ZN( u1_u5_u0_n172 ) , .A( u1_u5_u0_n88 ) );
  OAI222_X1 u1_u5_u0_U44 (.C1( u1_u5_u0_n108 ) , .A1( u1_u5_u0_n125 ) , .B2( u1_u5_u0_n128 ) , .B1( u1_u5_u0_n144 ) , .A2( u1_u5_u0_n158 ) , .C2( u1_u5_u0_n161 ) , .ZN( u1_u5_u0_n88 ) );
  NAND2_X1 u1_u5_u0_U45 (.A2( u1_u5_u0_n101 ) , .ZN( u1_u5_u0_n121 ) , .A1( u1_u5_u0_n93 ) );
  OR3_X1 u1_u5_u0_U46 (.A3( u1_u5_u0_n152 ) , .A2( u1_u5_u0_n153 ) , .A1( u1_u5_u0_n154 ) , .ZN( u1_u5_u0_n155 ) );
  AOI21_X1 u1_u5_u0_U47 (.A( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n145 ) , .B1( u1_u5_u0_n146 ) , .ZN( u1_u5_u0_n154 ) );
  AOI21_X1 u1_u5_u0_U48 (.B2( u1_u5_u0_n150 ) , .B1( u1_u5_u0_n151 ) , .ZN( u1_u5_u0_n152 ) , .A( u1_u5_u0_n158 ) );
  AOI21_X1 u1_u5_u0_U49 (.A( u1_u5_u0_n147 ) , .B2( u1_u5_u0_n148 ) , .B1( u1_u5_u0_n149 ) , .ZN( u1_u5_u0_n153 ) );
  AOI21_X1 u1_u5_u0_U5 (.B2( u1_u5_u0_n131 ) , .ZN( u1_u5_u0_n134 ) , .B1( u1_u5_u0_n151 ) , .A( u1_u5_u0_n158 ) );
  INV_X1 u1_u5_u0_U50 (.ZN( u1_u5_u0_n171 ) , .A( u1_u5_u0_n99 ) );
  OAI211_X1 u1_u5_u0_U51 (.C2( u1_u5_u0_n140 ) , .C1( u1_u5_u0_n161 ) , .A( u1_u5_u0_n169 ) , .B( u1_u5_u0_n98 ) , .ZN( u1_u5_u0_n99 ) );
  INV_X1 u1_u5_u0_U52 (.ZN( u1_u5_u0_n169 ) , .A( u1_u5_u0_n91 ) );
  AOI211_X1 u1_u5_u0_U53 (.C1( u1_u5_u0_n118 ) , .A( u1_u5_u0_n123 ) , .B( u1_u5_u0_n96 ) , .C2( u1_u5_u0_n97 ) , .ZN( u1_u5_u0_n98 ) );
  NOR2_X1 u1_u5_u0_U54 (.A2( u1_u5_X_4 ) , .A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n118 ) );
  NOR2_X1 u1_u5_u0_U55 (.A2( u1_u5_X_1 ) , .ZN( u1_u5_u0_n101 ) , .A1( u1_u5_u0_n163 ) );
  NOR2_X1 u1_u5_u0_U56 (.A2( u1_u5_X_3 ) , .A1( u1_u5_X_6 ) , .ZN( u1_u5_u0_n94 ) );
  NOR2_X1 u1_u5_u0_U57 (.A2( u1_u5_X_6 ) , .ZN( u1_u5_u0_n100 ) , .A1( u1_u5_u0_n162 ) );
  NAND2_X1 u1_u5_u0_U58 (.A2( u1_u5_X_4 ) , .A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n144 ) );
  NOR2_X1 u1_u5_u0_U59 (.A2( u1_u5_X_5 ) , .ZN( u1_u5_u0_n136 ) , .A1( u1_u5_u0_n159 ) );
  NOR2_X1 u1_u5_u0_U6 (.A1( u1_u5_u0_n108 ) , .ZN( u1_u5_u0_n123 ) , .A2( u1_u5_u0_n158 ) );
  NAND2_X1 u1_u5_u0_U60 (.A1( u1_u5_X_5 ) , .ZN( u1_u5_u0_n138 ) , .A2( u1_u5_u0_n159 ) );
  AND2_X1 u1_u5_u0_U61 (.A2( u1_u5_X_3 ) , .A1( u1_u5_X_6 ) , .ZN( u1_u5_u0_n102 ) );
  AND2_X1 u1_u5_u0_U62 (.A1( u1_u5_X_6 ) , .A2( u1_u5_u0_n162 ) , .ZN( u1_u5_u0_n93 ) );
  INV_X1 u1_u5_u0_U63 (.A( u1_u5_X_4 ) , .ZN( u1_u5_u0_n159 ) );
  INV_X1 u1_u5_u0_U64 (.A( u1_u5_X_1 ) , .ZN( u1_u5_u0_n164 ) );
  INV_X1 u1_u5_u0_U65 (.A( u1_u5_X_3 ) , .ZN( u1_u5_u0_n162 ) );
  INV_X1 u1_u5_u0_U66 (.A( u1_u5_u0_n126 ) , .ZN( u1_u5_u0_n168 ) );
  AOI211_X1 u1_u5_u0_U67 (.B( u1_u5_u0_n133 ) , .A( u1_u5_u0_n134 ) , .C2( u1_u5_u0_n135 ) , .C1( u1_u5_u0_n136 ) , .ZN( u1_u5_u0_n137 ) );
  OR4_X1 u1_u5_u0_U68 (.ZN( u1_out5_17 ) , .A1( u1_u5_u0_n122 ) , .A2( u1_u5_u0_n123 ) , .A4( u1_u5_u0_n124 ) , .A3( u1_u5_u0_n170 ) );
  AOI21_X1 u1_u5_u0_U69 (.B2( u1_u5_u0_n107 ) , .ZN( u1_u5_u0_n124 ) , .B1( u1_u5_u0_n128 ) , .A( u1_u5_u0_n161 ) );
  OAI21_X1 u1_u5_u0_U7 (.B1( u1_u5_u0_n150 ) , .B2( u1_u5_u0_n158 ) , .A( u1_u5_u0_n172 ) , .ZN( u1_u5_u0_n89 ) );
  INV_X1 u1_u5_u0_U70 (.A( u1_u5_u0_n111 ) , .ZN( u1_u5_u0_n170 ) );
  OR4_X1 u1_u5_u0_U71 (.ZN( u1_out5_31 ) , .A4( u1_u5_u0_n155 ) , .A2( u1_u5_u0_n156 ) , .A1( u1_u5_u0_n157 ) , .A3( u1_u5_u0_n173 ) );
  AOI21_X1 u1_u5_u0_U72 (.A( u1_u5_u0_n138 ) , .B2( u1_u5_u0_n139 ) , .B1( u1_u5_u0_n140 ) , .ZN( u1_u5_u0_n157 ) );
  AOI21_X1 u1_u5_u0_U73 (.B2( u1_u5_u0_n141 ) , .B1( u1_u5_u0_n142 ) , .ZN( u1_u5_u0_n156 ) , .A( u1_u5_u0_n161 ) );
  INV_X1 u1_u5_u0_U74 (.ZN( u1_u5_u0_n174 ) , .A( u1_u5_u0_n89 ) );
  AOI211_X1 u1_u5_u0_U75 (.B( u1_u5_u0_n104 ) , .A( u1_u5_u0_n105 ) , .ZN( u1_u5_u0_n106 ) , .C2( u1_u5_u0_n113 ) , .C1( u1_u5_u0_n160 ) );
  OAI221_X1 u1_u5_u0_U76 (.C1( u1_u5_u0_n121 ) , .ZN( u1_u5_u0_n122 ) , .B2( u1_u5_u0_n127 ) , .A( u1_u5_u0_n143 ) , .B1( u1_u5_u0_n144 ) , .C2( u1_u5_u0_n147 ) );
  AOI21_X1 u1_u5_u0_U77 (.B1( u1_u5_u0_n132 ) , .ZN( u1_u5_u0_n133 ) , .A( u1_u5_u0_n144 ) , .B2( u1_u5_u0_n166 ) );
  OAI22_X1 u1_u5_u0_U78 (.ZN( u1_u5_u0_n105 ) , .A2( u1_u5_u0_n132 ) , .B1( u1_u5_u0_n146 ) , .A1( u1_u5_u0_n147 ) , .B2( u1_u5_u0_n161 ) );
  NAND2_X1 u1_u5_u0_U79 (.ZN( u1_u5_u0_n110 ) , .A2( u1_u5_u0_n132 ) , .A1( u1_u5_u0_n145 ) );
  AND2_X1 u1_u5_u0_U8 (.A1( u1_u5_u0_n114 ) , .A2( u1_u5_u0_n121 ) , .ZN( u1_u5_u0_n146 ) );
  INV_X1 u1_u5_u0_U80 (.A( u1_u5_u0_n119 ) , .ZN( u1_u5_u0_n167 ) );
  NAND2_X1 u1_u5_u0_U81 (.ZN( u1_u5_u0_n148 ) , .A1( u1_u5_u0_n93 ) , .A2( u1_u5_u0_n95 ) );
  NAND2_X1 u1_u5_u0_U82 (.A1( u1_u5_u0_n100 ) , .ZN( u1_u5_u0_n129 ) , .A2( u1_u5_u0_n95 ) );
  NAND2_X1 u1_u5_u0_U83 (.A1( u1_u5_u0_n102 ) , .ZN( u1_u5_u0_n128 ) , .A2( u1_u5_u0_n95 ) );
  NOR2_X1 u1_u5_u0_U84 (.A2( u1_u5_X_1 ) , .A1( u1_u5_X_2 ) , .ZN( u1_u5_u0_n92 ) );
  NAND2_X1 u1_u5_u0_U85 (.ZN( u1_u5_u0_n142 ) , .A1( u1_u5_u0_n94 ) , .A2( u1_u5_u0_n95 ) );
  NOR2_X1 u1_u5_u0_U86 (.A2( u1_u5_X_2 ) , .ZN( u1_u5_u0_n103 ) , .A1( u1_u5_u0_n164 ) );
  INV_X1 u1_u5_u0_U87 (.A( u1_u5_X_2 ) , .ZN( u1_u5_u0_n163 ) );
  NAND3_X1 u1_u5_u0_U88 (.ZN( u1_out5_23 ) , .A3( u1_u5_u0_n137 ) , .A1( u1_u5_u0_n168 ) , .A2( u1_u5_u0_n171 ) );
  NAND3_X1 u1_u5_u0_U89 (.A3( u1_u5_u0_n127 ) , .A2( u1_u5_u0_n128 ) , .ZN( u1_u5_u0_n135 ) , .A1( u1_u5_u0_n150 ) );
  AND2_X1 u1_u5_u0_U9 (.A1( u1_u5_u0_n131 ) , .ZN( u1_u5_u0_n141 ) , .A2( u1_u5_u0_n150 ) );
  NAND3_X1 u1_u5_u0_U90 (.ZN( u1_u5_u0_n117 ) , .A3( u1_u5_u0_n132 ) , .A2( u1_u5_u0_n139 ) , .A1( u1_u5_u0_n148 ) );
  NAND3_X1 u1_u5_u0_U91 (.ZN( u1_u5_u0_n109 ) , .A2( u1_u5_u0_n114 ) , .A3( u1_u5_u0_n140 ) , .A1( u1_u5_u0_n149 ) );
  NAND3_X1 u1_u5_u0_U92 (.ZN( u1_out5_9 ) , .A3( u1_u5_u0_n106 ) , .A2( u1_u5_u0_n171 ) , .A1( u1_u5_u0_n174 ) );
  NAND3_X1 u1_u5_u0_U93 (.A2( u1_u5_u0_n128 ) , .A1( u1_u5_u0_n132 ) , .A3( u1_u5_u0_n146 ) , .ZN( u1_u5_u0_n97 ) );
  OAI22_X1 u1_u5_u2_U10 (.ZN( u1_u5_u2_n109 ) , .A2( u1_u5_u2_n113 ) , .B2( u1_u5_u2_n133 ) , .B1( u1_u5_u2_n167 ) , .A1( u1_u5_u2_n168 ) );
  NAND3_X1 u1_u5_u2_U100 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n104 ) , .A3( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n98 ) );
  OAI22_X1 u1_u5_u2_U11 (.B1( u1_u5_u2_n151 ) , .A2( u1_u5_u2_n152 ) , .A1( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n160 ) , .B2( u1_u5_u2_n168 ) );
  NOR3_X1 u1_u5_u2_U12 (.A1( u1_u5_u2_n150 ) , .ZN( u1_u5_u2_n151 ) , .A3( u1_u5_u2_n175 ) , .A2( u1_u5_u2_n188 ) );
  AOI21_X1 u1_u5_u2_U13 (.ZN( u1_u5_u2_n144 ) , .B2( u1_u5_u2_n155 ) , .A( u1_u5_u2_n172 ) , .B1( u1_u5_u2_n185 ) );
  AOI21_X1 u1_u5_u2_U14 (.B2( u1_u5_u2_n143 ) , .ZN( u1_u5_u2_n145 ) , .B1( u1_u5_u2_n152 ) , .A( u1_u5_u2_n171 ) );
  AOI21_X1 u1_u5_u2_U15 (.B2( u1_u5_u2_n120 ) , .B1( u1_u5_u2_n121 ) , .ZN( u1_u5_u2_n126 ) , .A( u1_u5_u2_n167 ) );
  INV_X1 u1_u5_u2_U16 (.A( u1_u5_u2_n156 ) , .ZN( u1_u5_u2_n171 ) );
  INV_X1 u1_u5_u2_U17 (.A( u1_u5_u2_n120 ) , .ZN( u1_u5_u2_n188 ) );
  NAND2_X1 u1_u5_u2_U18 (.A2( u1_u5_u2_n122 ) , .ZN( u1_u5_u2_n150 ) , .A1( u1_u5_u2_n152 ) );
  INV_X1 u1_u5_u2_U19 (.A( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n170 ) );
  INV_X1 u1_u5_u2_U20 (.A( u1_u5_u2_n137 ) , .ZN( u1_u5_u2_n173 ) );
  NAND2_X1 u1_u5_u2_U21 (.A1( u1_u5_u2_n132 ) , .A2( u1_u5_u2_n139 ) , .ZN( u1_u5_u2_n157 ) );
  INV_X1 u1_u5_u2_U22 (.A( u1_u5_u2_n113 ) , .ZN( u1_u5_u2_n178 ) );
  INV_X1 u1_u5_u2_U23 (.A( u1_u5_u2_n139 ) , .ZN( u1_u5_u2_n175 ) );
  INV_X1 u1_u5_u2_U24 (.A( u1_u5_u2_n155 ) , .ZN( u1_u5_u2_n181 ) );
  INV_X1 u1_u5_u2_U25 (.A( u1_u5_u2_n119 ) , .ZN( u1_u5_u2_n177 ) );
  INV_X1 u1_u5_u2_U26 (.A( u1_u5_u2_n116 ) , .ZN( u1_u5_u2_n180 ) );
  INV_X1 u1_u5_u2_U27 (.A( u1_u5_u2_n131 ) , .ZN( u1_u5_u2_n179 ) );
  INV_X1 u1_u5_u2_U28 (.A( u1_u5_u2_n154 ) , .ZN( u1_u5_u2_n176 ) );
  NAND2_X1 u1_u5_u2_U29 (.A2( u1_u5_u2_n116 ) , .A1( u1_u5_u2_n117 ) , .ZN( u1_u5_u2_n118 ) );
  NOR2_X1 u1_u5_u2_U3 (.ZN( u1_u5_u2_n121 ) , .A2( u1_u5_u2_n177 ) , .A1( u1_u5_u2_n180 ) );
  INV_X1 u1_u5_u2_U30 (.A( u1_u5_u2_n132 ) , .ZN( u1_u5_u2_n182 ) );
  INV_X1 u1_u5_u2_U31 (.A( u1_u5_u2_n158 ) , .ZN( u1_u5_u2_n183 ) );
  OAI21_X1 u1_u5_u2_U32 (.A( u1_u5_u2_n156 ) , .B1( u1_u5_u2_n157 ) , .ZN( u1_u5_u2_n158 ) , .B2( u1_u5_u2_n179 ) );
  NOR2_X1 u1_u5_u2_U33 (.ZN( u1_u5_u2_n156 ) , .A1( u1_u5_u2_n166 ) , .A2( u1_u5_u2_n169 ) );
  NOR2_X1 u1_u5_u2_U34 (.A2( u1_u5_u2_n114 ) , .ZN( u1_u5_u2_n137 ) , .A1( u1_u5_u2_n140 ) );
  NOR2_X1 u1_u5_u2_U35 (.A2( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n153 ) , .A1( u1_u5_u2_n156 ) );
  AOI211_X1 u1_u5_u2_U36 (.ZN( u1_u5_u2_n130 ) , .C1( u1_u5_u2_n138 ) , .C2( u1_u5_u2_n179 ) , .B( u1_u5_u2_n96 ) , .A( u1_u5_u2_n97 ) );
  OAI22_X1 u1_u5_u2_U37 (.B1( u1_u5_u2_n133 ) , .A2( u1_u5_u2_n137 ) , .A1( u1_u5_u2_n152 ) , .B2( u1_u5_u2_n168 ) , .ZN( u1_u5_u2_n97 ) );
  OAI221_X1 u1_u5_u2_U38 (.B1( u1_u5_u2_n113 ) , .C1( u1_u5_u2_n132 ) , .A( u1_u5_u2_n149 ) , .B2( u1_u5_u2_n171 ) , .C2( u1_u5_u2_n172 ) , .ZN( u1_u5_u2_n96 ) );
  OAI221_X1 u1_u5_u2_U39 (.A( u1_u5_u2_n115 ) , .C2( u1_u5_u2_n123 ) , .B2( u1_u5_u2_n143 ) , .B1( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n163 ) , .C1( u1_u5_u2_n168 ) );
  INV_X1 u1_u5_u2_U4 (.A( u1_u5_u2_n134 ) , .ZN( u1_u5_u2_n185 ) );
  OAI21_X1 u1_u5_u2_U40 (.A( u1_u5_u2_n114 ) , .ZN( u1_u5_u2_n115 ) , .B1( u1_u5_u2_n176 ) , .B2( u1_u5_u2_n178 ) );
  OAI221_X1 u1_u5_u2_U41 (.A( u1_u5_u2_n135 ) , .B2( u1_u5_u2_n136 ) , .B1( u1_u5_u2_n137 ) , .ZN( u1_u5_u2_n162 ) , .C2( u1_u5_u2_n167 ) , .C1( u1_u5_u2_n185 ) );
  AND3_X1 u1_u5_u2_U42 (.A3( u1_u5_u2_n131 ) , .A2( u1_u5_u2_n132 ) , .A1( u1_u5_u2_n133 ) , .ZN( u1_u5_u2_n136 ) );
  AOI22_X1 u1_u5_u2_U43 (.ZN( u1_u5_u2_n135 ) , .B1( u1_u5_u2_n140 ) , .A1( u1_u5_u2_n156 ) , .B2( u1_u5_u2_n180 ) , .A2( u1_u5_u2_n188 ) );
  AOI21_X1 u1_u5_u2_U44 (.ZN( u1_u5_u2_n149 ) , .B1( u1_u5_u2_n173 ) , .B2( u1_u5_u2_n188 ) , .A( u1_u5_u2_n95 ) );
  AND3_X1 u1_u5_u2_U45 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n104 ) , .A3( u1_u5_u2_n156 ) , .ZN( u1_u5_u2_n95 ) );
  OAI21_X1 u1_u5_u2_U46 (.A( u1_u5_u2_n101 ) , .B2( u1_u5_u2_n121 ) , .B1( u1_u5_u2_n153 ) , .ZN( u1_u5_u2_n164 ) );
  NAND2_X1 u1_u5_u2_U47 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n107 ) , .ZN( u1_u5_u2_n155 ) );
  NAND2_X1 u1_u5_u2_U48 (.A2( u1_u5_u2_n105 ) , .A1( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n143 ) );
  NAND2_X1 u1_u5_u2_U49 (.A1( u1_u5_u2_n104 ) , .A2( u1_u5_u2_n106 ) , .ZN( u1_u5_u2_n152 ) );
  INV_X1 u1_u5_u2_U5 (.A( u1_u5_u2_n150 ) , .ZN( u1_u5_u2_n184 ) );
  NAND2_X1 u1_u5_u2_U50 (.A1( u1_u5_u2_n100 ) , .A2( u1_u5_u2_n105 ) , .ZN( u1_u5_u2_n132 ) );
  INV_X1 u1_u5_u2_U51 (.A( u1_u5_u2_n140 ) , .ZN( u1_u5_u2_n168 ) );
  INV_X1 u1_u5_u2_U52 (.A( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n167 ) );
  OAI21_X1 u1_u5_u2_U53 (.A( u1_u5_u2_n141 ) , .B2( u1_u5_u2_n142 ) , .ZN( u1_u5_u2_n146 ) , .B1( u1_u5_u2_n153 ) );
  OAI21_X1 u1_u5_u2_U54 (.A( u1_u5_u2_n140 ) , .ZN( u1_u5_u2_n141 ) , .B1( u1_u5_u2_n176 ) , .B2( u1_u5_u2_n177 ) );
  NOR3_X1 u1_u5_u2_U55 (.ZN( u1_u5_u2_n142 ) , .A3( u1_u5_u2_n175 ) , .A2( u1_u5_u2_n178 ) , .A1( u1_u5_u2_n181 ) );
  INV_X1 u1_u5_u2_U56 (.ZN( u1_u5_u2_n187 ) , .A( u1_u5_u2_n99 ) );
  OAI21_X1 u1_u5_u2_U57 (.B1( u1_u5_u2_n137 ) , .B2( u1_u5_u2_n143 ) , .A( u1_u5_u2_n98 ) , .ZN( u1_u5_u2_n99 ) );
  NAND2_X1 u1_u5_u2_U58 (.A1( u1_u5_u2_n102 ) , .A2( u1_u5_u2_n106 ) , .ZN( u1_u5_u2_n113 ) );
  NAND2_X1 u1_u5_u2_U59 (.A1( u1_u5_u2_n106 ) , .A2( u1_u5_u2_n107 ) , .ZN( u1_u5_u2_n131 ) );
  NOR4_X1 u1_u5_u2_U6 (.A4( u1_u5_u2_n124 ) , .A3( u1_u5_u2_n125 ) , .A2( u1_u5_u2_n126 ) , .A1( u1_u5_u2_n127 ) , .ZN( u1_u5_u2_n128 ) );
  NAND2_X1 u1_u5_u2_U60 (.A1( u1_u5_u2_n103 ) , .A2( u1_u5_u2_n107 ) , .ZN( u1_u5_u2_n139 ) );
  NAND2_X1 u1_u5_u2_U61 (.A1( u1_u5_u2_n103 ) , .A2( u1_u5_u2_n105 ) , .ZN( u1_u5_u2_n133 ) );
  NAND2_X1 u1_u5_u2_U62 (.A1( u1_u5_u2_n102 ) , .A2( u1_u5_u2_n103 ) , .ZN( u1_u5_u2_n154 ) );
  NAND2_X1 u1_u5_u2_U63 (.A2( u1_u5_u2_n103 ) , .A1( u1_u5_u2_n104 ) , .ZN( u1_u5_u2_n119 ) );
  NAND2_X1 u1_u5_u2_U64 (.A2( u1_u5_u2_n107 ) , .A1( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n123 ) );
  NAND2_X1 u1_u5_u2_U65 (.A1( u1_u5_u2_n104 ) , .A2( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n122 ) );
  INV_X1 u1_u5_u2_U66 (.A( u1_u5_u2_n114 ) , .ZN( u1_u5_u2_n172 ) );
  NAND2_X1 u1_u5_u2_U67 (.A2( u1_u5_u2_n100 ) , .A1( u1_u5_u2_n102 ) , .ZN( u1_u5_u2_n116 ) );
  NAND2_X1 u1_u5_u2_U68 (.A1( u1_u5_u2_n102 ) , .A2( u1_u5_u2_n108 ) , .ZN( u1_u5_u2_n120 ) );
  NAND2_X1 u1_u5_u2_U69 (.A2( u1_u5_u2_n105 ) , .A1( u1_u5_u2_n106 ) , .ZN( u1_u5_u2_n117 ) );
  AOI21_X1 u1_u5_u2_U7 (.B2( u1_u5_u2_n119 ) , .ZN( u1_u5_u2_n127 ) , .A( u1_u5_u2_n137 ) , .B1( u1_u5_u2_n155 ) );
  NOR2_X1 u1_u5_u2_U70 (.A2( u1_u5_X_16 ) , .ZN( u1_u5_u2_n140 ) , .A1( u1_u5_u2_n166 ) );
  NOR2_X1 u1_u5_u2_U71 (.A2( u1_u5_X_13 ) , .A1( u1_u5_X_14 ) , .ZN( u1_u5_u2_n100 ) );
  NOR2_X1 u1_u5_u2_U72 (.A2( u1_u5_X_16 ) , .A1( u1_u5_X_17 ) , .ZN( u1_u5_u2_n138 ) );
  NOR2_X1 u1_u5_u2_U73 (.A2( u1_u5_X_15 ) , .A1( u1_u5_X_18 ) , .ZN( u1_u5_u2_n104 ) );
  NOR2_X1 u1_u5_u2_U74 (.A2( u1_u5_X_14 ) , .ZN( u1_u5_u2_n103 ) , .A1( u1_u5_u2_n174 ) );
  NOR2_X1 u1_u5_u2_U75 (.A2( u1_u5_X_15 ) , .ZN( u1_u5_u2_n102 ) , .A1( u1_u5_u2_n165 ) );
  NOR2_X1 u1_u5_u2_U76 (.A2( u1_u5_X_17 ) , .ZN( u1_u5_u2_n114 ) , .A1( u1_u5_u2_n169 ) );
  AND2_X1 u1_u5_u2_U77 (.A1( u1_u5_X_15 ) , .ZN( u1_u5_u2_n105 ) , .A2( u1_u5_u2_n165 ) );
  AND2_X1 u1_u5_u2_U78 (.A2( u1_u5_X_15 ) , .A1( u1_u5_X_18 ) , .ZN( u1_u5_u2_n107 ) );
  AND2_X1 u1_u5_u2_U79 (.A1( u1_u5_X_14 ) , .ZN( u1_u5_u2_n106 ) , .A2( u1_u5_u2_n174 ) );
  AOI21_X1 u1_u5_u2_U8 (.ZN( u1_u5_u2_n124 ) , .B1( u1_u5_u2_n131 ) , .B2( u1_u5_u2_n143 ) , .A( u1_u5_u2_n172 ) );
  AND2_X1 u1_u5_u2_U80 (.A1( u1_u5_X_13 ) , .A2( u1_u5_X_14 ) , .ZN( u1_u5_u2_n108 ) );
  INV_X1 u1_u5_u2_U81 (.A( u1_u5_X_16 ) , .ZN( u1_u5_u2_n169 ) );
  INV_X1 u1_u5_u2_U82 (.A( u1_u5_X_17 ) , .ZN( u1_u5_u2_n166 ) );
  INV_X1 u1_u5_u2_U83 (.A( u1_u5_X_13 ) , .ZN( u1_u5_u2_n174 ) );
  INV_X1 u1_u5_u2_U84 (.A( u1_u5_X_18 ) , .ZN( u1_u5_u2_n165 ) );
  NAND4_X1 u1_u5_u2_U85 (.ZN( u1_out5_30 ) , .A4( u1_u5_u2_n147 ) , .A3( u1_u5_u2_n148 ) , .A2( u1_u5_u2_n149 ) , .A1( u1_u5_u2_n187 ) );
  NOR3_X1 u1_u5_u2_U86 (.A3( u1_u5_u2_n144 ) , .A2( u1_u5_u2_n145 ) , .A1( u1_u5_u2_n146 ) , .ZN( u1_u5_u2_n147 ) );
  AOI21_X1 u1_u5_u2_U87 (.B2( u1_u5_u2_n138 ) , .ZN( u1_u5_u2_n148 ) , .A( u1_u5_u2_n162 ) , .B1( u1_u5_u2_n182 ) );
  NAND4_X1 u1_u5_u2_U88 (.ZN( u1_out5_24 ) , .A4( u1_u5_u2_n111 ) , .A3( u1_u5_u2_n112 ) , .A1( u1_u5_u2_n130 ) , .A2( u1_u5_u2_n187 ) );
  AOI221_X1 u1_u5_u2_U89 (.A( u1_u5_u2_n109 ) , .B1( u1_u5_u2_n110 ) , .ZN( u1_u5_u2_n111 ) , .C1( u1_u5_u2_n134 ) , .C2( u1_u5_u2_n170 ) , .B2( u1_u5_u2_n173 ) );
  AOI21_X1 u1_u5_u2_U9 (.B2( u1_u5_u2_n123 ) , .ZN( u1_u5_u2_n125 ) , .A( u1_u5_u2_n171 ) , .B1( u1_u5_u2_n184 ) );
  AOI21_X1 u1_u5_u2_U90 (.ZN( u1_u5_u2_n112 ) , .B2( u1_u5_u2_n156 ) , .A( u1_u5_u2_n164 ) , .B1( u1_u5_u2_n181 ) );
  NAND4_X1 u1_u5_u2_U91 (.ZN( u1_out5_16 ) , .A4( u1_u5_u2_n128 ) , .A3( u1_u5_u2_n129 ) , .A1( u1_u5_u2_n130 ) , .A2( u1_u5_u2_n186 ) );
  AOI22_X1 u1_u5_u2_U92 (.A2( u1_u5_u2_n118 ) , .ZN( u1_u5_u2_n129 ) , .A1( u1_u5_u2_n140 ) , .B1( u1_u5_u2_n157 ) , .B2( u1_u5_u2_n170 ) );
  INV_X1 u1_u5_u2_U93 (.A( u1_u5_u2_n163 ) , .ZN( u1_u5_u2_n186 ) );
  OR4_X1 u1_u5_u2_U94 (.ZN( u1_out5_6 ) , .A4( u1_u5_u2_n161 ) , .A3( u1_u5_u2_n162 ) , .A2( u1_u5_u2_n163 ) , .A1( u1_u5_u2_n164 ) );
  OR3_X1 u1_u5_u2_U95 (.A2( u1_u5_u2_n159 ) , .A1( u1_u5_u2_n160 ) , .ZN( u1_u5_u2_n161 ) , .A3( u1_u5_u2_n183 ) );
  AOI21_X1 u1_u5_u2_U96 (.B2( u1_u5_u2_n154 ) , .B1( u1_u5_u2_n155 ) , .ZN( u1_u5_u2_n159 ) , .A( u1_u5_u2_n167 ) );
  NAND3_X1 u1_u5_u2_U97 (.A2( u1_u5_u2_n117 ) , .A1( u1_u5_u2_n122 ) , .A3( u1_u5_u2_n123 ) , .ZN( u1_u5_u2_n134 ) );
  NAND3_X1 u1_u5_u2_U98 (.ZN( u1_u5_u2_n110 ) , .A2( u1_u5_u2_n131 ) , .A3( u1_u5_u2_n139 ) , .A1( u1_u5_u2_n154 ) );
  NAND3_X1 u1_u5_u2_U99 (.A2( u1_u5_u2_n100 ) , .ZN( u1_u5_u2_n101 ) , .A1( u1_u5_u2_n104 ) , .A3( u1_u5_u2_n114 ) );
  OAI22_X1 u1_u5_u3_U10 (.B1( u1_u5_u3_n113 ) , .A2( u1_u5_u3_n135 ) , .A1( u1_u5_u3_n150 ) , .B2( u1_u5_u3_n164 ) , .ZN( u1_u5_u3_n98 ) );
  OAI211_X1 u1_u5_u3_U11 (.B( u1_u5_u3_n106 ) , .ZN( u1_u5_u3_n119 ) , .C2( u1_u5_u3_n128 ) , .C1( u1_u5_u3_n167 ) , .A( u1_u5_u3_n181 ) );
  AOI221_X1 u1_u5_u3_U12 (.C1( u1_u5_u3_n105 ) , .ZN( u1_u5_u3_n106 ) , .A( u1_u5_u3_n131 ) , .B2( u1_u5_u3_n132 ) , .C2( u1_u5_u3_n133 ) , .B1( u1_u5_u3_n169 ) );
  INV_X1 u1_u5_u3_U13 (.ZN( u1_u5_u3_n181 ) , .A( u1_u5_u3_n98 ) );
  NAND2_X1 u1_u5_u3_U14 (.ZN( u1_u5_u3_n105 ) , .A2( u1_u5_u3_n130 ) , .A1( u1_u5_u3_n155 ) );
  AOI22_X1 u1_u5_u3_U15 (.B1( u1_u5_u3_n115 ) , .A2( u1_u5_u3_n116 ) , .ZN( u1_u5_u3_n123 ) , .B2( u1_u5_u3_n133 ) , .A1( u1_u5_u3_n169 ) );
  NAND2_X1 u1_u5_u3_U16 (.ZN( u1_u5_u3_n116 ) , .A2( u1_u5_u3_n151 ) , .A1( u1_u5_u3_n182 ) );
  NOR2_X1 u1_u5_u3_U17 (.ZN( u1_u5_u3_n126 ) , .A2( u1_u5_u3_n150 ) , .A1( u1_u5_u3_n164 ) );
  AOI21_X1 u1_u5_u3_U18 (.ZN( u1_u5_u3_n112 ) , .B2( u1_u5_u3_n146 ) , .B1( u1_u5_u3_n155 ) , .A( u1_u5_u3_n167 ) );
  NAND2_X1 u1_u5_u3_U19 (.A1( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n142 ) , .A2( u1_u5_u3_n164 ) );
  NAND2_X1 u1_u5_u3_U20 (.ZN( u1_u5_u3_n132 ) , .A2( u1_u5_u3_n152 ) , .A1( u1_u5_u3_n156 ) );
  AND2_X1 u1_u5_u3_U21 (.A2( u1_u5_u3_n113 ) , .A1( u1_u5_u3_n114 ) , .ZN( u1_u5_u3_n151 ) );
  INV_X1 u1_u5_u3_U22 (.A( u1_u5_u3_n133 ) , .ZN( u1_u5_u3_n165 ) );
  INV_X1 u1_u5_u3_U23 (.A( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n170 ) );
  NAND2_X1 u1_u5_u3_U24 (.A1( u1_u5_u3_n107 ) , .A2( u1_u5_u3_n108 ) , .ZN( u1_u5_u3_n140 ) );
  NAND2_X1 u1_u5_u3_U25 (.ZN( u1_u5_u3_n117 ) , .A1( u1_u5_u3_n124 ) , .A2( u1_u5_u3_n148 ) );
  NAND2_X1 u1_u5_u3_U26 (.ZN( u1_u5_u3_n143 ) , .A1( u1_u5_u3_n165 ) , .A2( u1_u5_u3_n167 ) );
  INV_X1 u1_u5_u3_U27 (.A( u1_u5_u3_n130 ) , .ZN( u1_u5_u3_n177 ) );
  INV_X1 u1_u5_u3_U28 (.A( u1_u5_u3_n128 ) , .ZN( u1_u5_u3_n176 ) );
  INV_X1 u1_u5_u3_U29 (.A( u1_u5_u3_n155 ) , .ZN( u1_u5_u3_n174 ) );
  INV_X1 u1_u5_u3_U3 (.A( u1_u5_u3_n129 ) , .ZN( u1_u5_u3_n183 ) );
  INV_X1 u1_u5_u3_U30 (.A( u1_u5_u3_n139 ) , .ZN( u1_u5_u3_n185 ) );
  NOR2_X1 u1_u5_u3_U31 (.ZN( u1_u5_u3_n135 ) , .A2( u1_u5_u3_n141 ) , .A1( u1_u5_u3_n169 ) );
  OAI222_X1 u1_u5_u3_U32 (.C2( u1_u5_u3_n107 ) , .A2( u1_u5_u3_n108 ) , .B1( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n138 ) , .B2( u1_u5_u3_n146 ) , .C1( u1_u5_u3_n154 ) , .A1( u1_u5_u3_n164 ) );
  NOR4_X1 u1_u5_u3_U33 (.A4( u1_u5_u3_n157 ) , .A3( u1_u5_u3_n158 ) , .A2( u1_u5_u3_n159 ) , .A1( u1_u5_u3_n160 ) , .ZN( u1_u5_u3_n161 ) );
  AOI21_X1 u1_u5_u3_U34 (.B2( u1_u5_u3_n152 ) , .B1( u1_u5_u3_n153 ) , .ZN( u1_u5_u3_n158 ) , .A( u1_u5_u3_n164 ) );
  AOI21_X1 u1_u5_u3_U35 (.A( u1_u5_u3_n154 ) , .B2( u1_u5_u3_n155 ) , .B1( u1_u5_u3_n156 ) , .ZN( u1_u5_u3_n157 ) );
  AOI21_X1 u1_u5_u3_U36 (.A( u1_u5_u3_n149 ) , .B2( u1_u5_u3_n150 ) , .B1( u1_u5_u3_n151 ) , .ZN( u1_u5_u3_n159 ) );
  AOI211_X1 u1_u5_u3_U37 (.ZN( u1_u5_u3_n109 ) , .A( u1_u5_u3_n119 ) , .C2( u1_u5_u3_n129 ) , .B( u1_u5_u3_n138 ) , .C1( u1_u5_u3_n141 ) );
  AOI211_X1 u1_u5_u3_U38 (.B( u1_u5_u3_n119 ) , .A( u1_u5_u3_n120 ) , .C2( u1_u5_u3_n121 ) , .ZN( u1_u5_u3_n122 ) , .C1( u1_u5_u3_n179 ) );
  INV_X1 u1_u5_u3_U39 (.A( u1_u5_u3_n156 ) , .ZN( u1_u5_u3_n179 ) );
  INV_X1 u1_u5_u3_U4 (.A( u1_u5_u3_n140 ) , .ZN( u1_u5_u3_n182 ) );
  OAI22_X1 u1_u5_u3_U40 (.B1( u1_u5_u3_n118 ) , .ZN( u1_u5_u3_n120 ) , .A1( u1_u5_u3_n135 ) , .B2( u1_u5_u3_n154 ) , .A2( u1_u5_u3_n178 ) );
  AND3_X1 u1_u5_u3_U41 (.ZN( u1_u5_u3_n118 ) , .A2( u1_u5_u3_n124 ) , .A1( u1_u5_u3_n144 ) , .A3( u1_u5_u3_n152 ) );
  INV_X1 u1_u5_u3_U42 (.A( u1_u5_u3_n121 ) , .ZN( u1_u5_u3_n164 ) );
  NAND2_X1 u1_u5_u3_U43 (.ZN( u1_u5_u3_n133 ) , .A1( u1_u5_u3_n154 ) , .A2( u1_u5_u3_n164 ) );
  OAI211_X1 u1_u5_u3_U44 (.B( u1_u5_u3_n127 ) , .ZN( u1_u5_u3_n139 ) , .C1( u1_u5_u3_n150 ) , .C2( u1_u5_u3_n154 ) , .A( u1_u5_u3_n184 ) );
  INV_X1 u1_u5_u3_U45 (.A( u1_u5_u3_n125 ) , .ZN( u1_u5_u3_n184 ) );
  AOI221_X1 u1_u5_u3_U46 (.A( u1_u5_u3_n126 ) , .ZN( u1_u5_u3_n127 ) , .C2( u1_u5_u3_n132 ) , .C1( u1_u5_u3_n169 ) , .B2( u1_u5_u3_n170 ) , .B1( u1_u5_u3_n174 ) );
  OAI22_X1 u1_u5_u3_U47 (.A1( u1_u5_u3_n124 ) , .ZN( u1_u5_u3_n125 ) , .B2( u1_u5_u3_n145 ) , .A2( u1_u5_u3_n165 ) , .B1( u1_u5_u3_n167 ) );
  NOR2_X1 u1_u5_u3_U48 (.A1( u1_u5_u3_n113 ) , .ZN( u1_u5_u3_n131 ) , .A2( u1_u5_u3_n154 ) );
  NAND2_X1 u1_u5_u3_U49 (.A1( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n150 ) , .A2( u1_u5_u3_n99 ) );
  INV_X1 u1_u5_u3_U5 (.A( u1_u5_u3_n117 ) , .ZN( u1_u5_u3_n178 ) );
  NAND2_X1 u1_u5_u3_U50 (.A2( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n155 ) , .A1( u1_u5_u3_n97 ) );
  INV_X1 u1_u5_u3_U51 (.A( u1_u5_u3_n141 ) , .ZN( u1_u5_u3_n167 ) );
  AOI21_X1 u1_u5_u3_U52 (.B2( u1_u5_u3_n114 ) , .B1( u1_u5_u3_n146 ) , .A( u1_u5_u3_n154 ) , .ZN( u1_u5_u3_n94 ) );
  AOI21_X1 u1_u5_u3_U53 (.ZN( u1_u5_u3_n110 ) , .B2( u1_u5_u3_n142 ) , .B1( u1_u5_u3_n186 ) , .A( u1_u5_u3_n95 ) );
  INV_X1 u1_u5_u3_U54 (.A( u1_u5_u3_n145 ) , .ZN( u1_u5_u3_n186 ) );
  AOI21_X1 u1_u5_u3_U55 (.B1( u1_u5_u3_n124 ) , .A( u1_u5_u3_n149 ) , .B2( u1_u5_u3_n155 ) , .ZN( u1_u5_u3_n95 ) );
  INV_X1 u1_u5_u3_U56 (.A( u1_u5_u3_n149 ) , .ZN( u1_u5_u3_n169 ) );
  NAND2_X1 u1_u5_u3_U57 (.ZN( u1_u5_u3_n124 ) , .A1( u1_u5_u3_n96 ) , .A2( u1_u5_u3_n97 ) );
  NAND2_X1 u1_u5_u3_U58 (.A2( u1_u5_u3_n100 ) , .ZN( u1_u5_u3_n146 ) , .A1( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U59 (.A1( u1_u5_u3_n101 ) , .ZN( u1_u5_u3_n145 ) , .A2( u1_u5_u3_n99 ) );
  AOI221_X1 u1_u5_u3_U6 (.A( u1_u5_u3_n131 ) , .C2( u1_u5_u3_n132 ) , .C1( u1_u5_u3_n133 ) , .ZN( u1_u5_u3_n134 ) , .B1( u1_u5_u3_n143 ) , .B2( u1_u5_u3_n177 ) );
  NAND2_X1 u1_u5_u3_U60 (.A1( u1_u5_u3_n100 ) , .ZN( u1_u5_u3_n156 ) , .A2( u1_u5_u3_n99 ) );
  NAND2_X1 u1_u5_u3_U61 (.A2( u1_u5_u3_n101 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n148 ) );
  NAND2_X1 u1_u5_u3_U62 (.A1( u1_u5_u3_n100 ) , .A2( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n128 ) );
  NAND2_X1 u1_u5_u3_U63 (.A2( u1_u5_u3_n101 ) , .A1( u1_u5_u3_n102 ) , .ZN( u1_u5_u3_n152 ) );
  NAND2_X1 u1_u5_u3_U64 (.A2( u1_u5_u3_n101 ) , .ZN( u1_u5_u3_n114 ) , .A1( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U65 (.ZN( u1_u5_u3_n107 ) , .A1( u1_u5_u3_n97 ) , .A2( u1_u5_u3_n99 ) );
  NAND2_X1 u1_u5_u3_U66 (.A2( u1_u5_u3_n100 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n113 ) );
  NAND2_X1 u1_u5_u3_U67 (.A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n153 ) , .A2( u1_u5_u3_n97 ) );
  NAND2_X1 u1_u5_u3_U68 (.A2( u1_u5_u3_n103 ) , .A1( u1_u5_u3_n104 ) , .ZN( u1_u5_u3_n130 ) );
  NAND2_X1 u1_u5_u3_U69 (.A2( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n144 ) , .A1( u1_u5_u3_n96 ) );
  OAI22_X1 u1_u5_u3_U7 (.B2( u1_u5_u3_n147 ) , .A2( u1_u5_u3_n148 ) , .ZN( u1_u5_u3_n160 ) , .B1( u1_u5_u3_n165 ) , .A1( u1_u5_u3_n168 ) );
  NAND2_X1 u1_u5_u3_U70 (.A1( u1_u5_u3_n102 ) , .A2( u1_u5_u3_n103 ) , .ZN( u1_u5_u3_n108 ) );
  NOR2_X1 u1_u5_u3_U71 (.A2( u1_u5_X_19 ) , .A1( u1_u5_X_20 ) , .ZN( u1_u5_u3_n99 ) );
  NOR2_X1 u1_u5_u3_U72 (.A2( u1_u5_X_21 ) , .A1( u1_u5_X_24 ) , .ZN( u1_u5_u3_n103 ) );
  NOR2_X1 u1_u5_u3_U73 (.A2( u1_u5_X_24 ) , .A1( u1_u5_u3_n171 ) , .ZN( u1_u5_u3_n97 ) );
  NOR2_X1 u1_u5_u3_U74 (.A2( u1_u5_X_23 ) , .ZN( u1_u5_u3_n141 ) , .A1( u1_u5_u3_n166 ) );
  NOR2_X1 u1_u5_u3_U75 (.A2( u1_u5_X_19 ) , .A1( u1_u5_u3_n172 ) , .ZN( u1_u5_u3_n96 ) );
  NAND2_X1 u1_u5_u3_U76 (.A1( u1_u5_X_22 ) , .A2( u1_u5_X_23 ) , .ZN( u1_u5_u3_n154 ) );
  NAND2_X1 u1_u5_u3_U77 (.A1( u1_u5_X_23 ) , .ZN( u1_u5_u3_n149 ) , .A2( u1_u5_u3_n166 ) );
  NOR2_X1 u1_u5_u3_U78 (.A2( u1_u5_X_22 ) , .A1( u1_u5_X_23 ) , .ZN( u1_u5_u3_n121 ) );
  AND2_X1 u1_u5_u3_U79 (.A1( u1_u5_X_24 ) , .ZN( u1_u5_u3_n101 ) , .A2( u1_u5_u3_n171 ) );
  AND3_X1 u1_u5_u3_U8 (.A3( u1_u5_u3_n144 ) , .A2( u1_u5_u3_n145 ) , .A1( u1_u5_u3_n146 ) , .ZN( u1_u5_u3_n147 ) );
  AND2_X1 u1_u5_u3_U80 (.A1( u1_u5_X_19 ) , .ZN( u1_u5_u3_n102 ) , .A2( u1_u5_u3_n172 ) );
  AND2_X1 u1_u5_u3_U81 (.A1( u1_u5_X_21 ) , .A2( u1_u5_X_24 ) , .ZN( u1_u5_u3_n100 ) );
  AND2_X1 u1_u5_u3_U82 (.A2( u1_u5_X_19 ) , .A1( u1_u5_X_20 ) , .ZN( u1_u5_u3_n104 ) );
  INV_X1 u1_u5_u3_U83 (.A( u1_u5_X_22 ) , .ZN( u1_u5_u3_n166 ) );
  INV_X1 u1_u5_u3_U84 (.A( u1_u5_X_21 ) , .ZN( u1_u5_u3_n171 ) );
  INV_X1 u1_u5_u3_U85 (.A( u1_u5_X_20 ) , .ZN( u1_u5_u3_n172 ) );
  NAND4_X1 u1_u5_u3_U86 (.ZN( u1_out5_26 ) , .A4( u1_u5_u3_n109 ) , .A3( u1_u5_u3_n110 ) , .A2( u1_u5_u3_n111 ) , .A1( u1_u5_u3_n173 ) );
  INV_X1 u1_u5_u3_U87 (.ZN( u1_u5_u3_n173 ) , .A( u1_u5_u3_n94 ) );
  OAI21_X1 u1_u5_u3_U88 (.ZN( u1_u5_u3_n111 ) , .B2( u1_u5_u3_n117 ) , .A( u1_u5_u3_n133 ) , .B1( u1_u5_u3_n176 ) );
  NAND4_X1 u1_u5_u3_U89 (.ZN( u1_out5_20 ) , .A4( u1_u5_u3_n122 ) , .A3( u1_u5_u3_n123 ) , .A1( u1_u5_u3_n175 ) , .A2( u1_u5_u3_n180 ) );
  INV_X1 u1_u5_u3_U9 (.A( u1_u5_u3_n143 ) , .ZN( u1_u5_u3_n168 ) );
  INV_X1 u1_u5_u3_U90 (.A( u1_u5_u3_n126 ) , .ZN( u1_u5_u3_n180 ) );
  INV_X1 u1_u5_u3_U91 (.A( u1_u5_u3_n112 ) , .ZN( u1_u5_u3_n175 ) );
  OR4_X1 u1_u5_u3_U92 (.ZN( u1_out5_10 ) , .A4( u1_u5_u3_n136 ) , .A3( u1_u5_u3_n137 ) , .A1( u1_u5_u3_n138 ) , .A2( u1_u5_u3_n139 ) );
  OAI222_X1 u1_u5_u3_U93 (.C1( u1_u5_u3_n128 ) , .ZN( u1_u5_u3_n137 ) , .B1( u1_u5_u3_n148 ) , .A2( u1_u5_u3_n150 ) , .B2( u1_u5_u3_n154 ) , .C2( u1_u5_u3_n164 ) , .A1( u1_u5_u3_n167 ) );
  OAI221_X1 u1_u5_u3_U94 (.A( u1_u5_u3_n134 ) , .B2( u1_u5_u3_n135 ) , .ZN( u1_u5_u3_n136 ) , .C1( u1_u5_u3_n149 ) , .B1( u1_u5_u3_n151 ) , .C2( u1_u5_u3_n183 ) );
  NAND4_X1 u1_u5_u3_U95 (.ZN( u1_out5_1 ) , .A4( u1_u5_u3_n161 ) , .A3( u1_u5_u3_n162 ) , .A2( u1_u5_u3_n163 ) , .A1( u1_u5_u3_n185 ) );
  NAND2_X1 u1_u5_u3_U96 (.ZN( u1_u5_u3_n163 ) , .A2( u1_u5_u3_n170 ) , .A1( u1_u5_u3_n176 ) );
  AOI22_X1 u1_u5_u3_U97 (.B2( u1_u5_u3_n140 ) , .B1( u1_u5_u3_n141 ) , .A2( u1_u5_u3_n142 ) , .ZN( u1_u5_u3_n162 ) , .A1( u1_u5_u3_n177 ) );
  NAND3_X1 u1_u5_u3_U98 (.A1( u1_u5_u3_n114 ) , .ZN( u1_u5_u3_n115 ) , .A2( u1_u5_u3_n145 ) , .A3( u1_u5_u3_n153 ) );
  NAND3_X1 u1_u5_u3_U99 (.ZN( u1_u5_u3_n129 ) , .A2( u1_u5_u3_n144 ) , .A1( u1_u5_u3_n153 ) , .A3( u1_u5_u3_n182 ) );
  OAI21_X1 u1_u5_u6_U10 (.A( u1_u5_u6_n159 ) , .B1( u1_u5_u6_n169 ) , .B2( u1_u5_u6_n173 ) , .ZN( u1_u5_u6_n90 ) );
  INV_X1 u1_u5_u6_U11 (.ZN( u1_u5_u6_n172 ) , .A( u1_u5_u6_n88 ) );
  AOI22_X1 u1_u5_u6_U12 (.A2( u1_u5_u6_n151 ) , .B2( u1_u5_u6_n161 ) , .A1( u1_u5_u6_n167 ) , .B1( u1_u5_u6_n170 ) , .ZN( u1_u5_u6_n89 ) );
  AOI21_X1 u1_u5_u6_U13 (.ZN( u1_u5_u6_n106 ) , .A( u1_u5_u6_n142 ) , .B2( u1_u5_u6_n159 ) , .B1( u1_u5_u6_n164 ) );
  INV_X1 u1_u5_u6_U14 (.A( u1_u5_u6_n155 ) , .ZN( u1_u5_u6_n161 ) );
  INV_X1 u1_u5_u6_U15 (.A( u1_u5_u6_n128 ) , .ZN( u1_u5_u6_n164 ) );
  NAND2_X1 u1_u5_u6_U16 (.ZN( u1_u5_u6_n110 ) , .A1( u1_u5_u6_n122 ) , .A2( u1_u5_u6_n129 ) );
  NAND2_X1 u1_u5_u6_U17 (.ZN( u1_u5_u6_n124 ) , .A2( u1_u5_u6_n146 ) , .A1( u1_u5_u6_n148 ) );
  INV_X1 u1_u5_u6_U18 (.A( u1_u5_u6_n132 ) , .ZN( u1_u5_u6_n171 ) );
  AND2_X1 u1_u5_u6_U19 (.A1( u1_u5_u6_n100 ) , .ZN( u1_u5_u6_n130 ) , .A2( u1_u5_u6_n147 ) );
  INV_X1 u1_u5_u6_U20 (.A( u1_u5_u6_n127 ) , .ZN( u1_u5_u6_n173 ) );
  INV_X1 u1_u5_u6_U21 (.A( u1_u5_u6_n121 ) , .ZN( u1_u5_u6_n167 ) );
  INV_X1 u1_u5_u6_U22 (.A( u1_u5_u6_n100 ) , .ZN( u1_u5_u6_n169 ) );
  INV_X1 u1_u5_u6_U23 (.A( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n170 ) );
  INV_X1 u1_u5_u6_U24 (.A( u1_u5_u6_n113 ) , .ZN( u1_u5_u6_n168 ) );
  AND2_X1 u1_u5_u6_U25 (.A1( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n119 ) , .ZN( u1_u5_u6_n133 ) );
  AND2_X1 u1_u5_u6_U26 (.A2( u1_u5_u6_n121 ) , .A1( u1_u5_u6_n122 ) , .ZN( u1_u5_u6_n131 ) );
  AND3_X1 u1_u5_u6_U27 (.ZN( u1_u5_u6_n120 ) , .A2( u1_u5_u6_n127 ) , .A1( u1_u5_u6_n132 ) , .A3( u1_u5_u6_n145 ) );
  INV_X1 u1_u5_u6_U28 (.A( u1_u5_u6_n146 ) , .ZN( u1_u5_u6_n163 ) );
  AOI222_X1 u1_u5_u6_U29 (.ZN( u1_u5_u6_n114 ) , .A1( u1_u5_u6_n118 ) , .A2( u1_u5_u6_n126 ) , .B2( u1_u5_u6_n151 ) , .C2( u1_u5_u6_n159 ) , .C1( u1_u5_u6_n168 ) , .B1( u1_u5_u6_n169 ) );
  INV_X1 u1_u5_u6_U3 (.A( u1_u5_u6_n110 ) , .ZN( u1_u5_u6_n166 ) );
  NOR2_X1 u1_u5_u6_U30 (.A1( u1_u5_u6_n162 ) , .A2( u1_u5_u6_n165 ) , .ZN( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U31 (.A1( u1_u5_u6_n144 ) , .ZN( u1_u5_u6_n151 ) , .A2( u1_u5_u6_n158 ) );
  NAND2_X1 u1_u5_u6_U32 (.ZN( u1_u5_u6_n132 ) , .A1( u1_u5_u6_n91 ) , .A2( u1_u5_u6_n97 ) );
  NOR2_X1 u1_u5_u6_U33 (.A2( u1_u5_u6_n126 ) , .ZN( u1_u5_u6_n155 ) , .A1( u1_u5_u6_n160 ) );
  NAND2_X1 u1_u5_u6_U34 (.ZN( u1_u5_u6_n146 ) , .A2( u1_u5_u6_n94 ) , .A1( u1_u5_u6_n99 ) );
  AOI21_X1 u1_u5_u6_U35 (.A( u1_u5_u6_n144 ) , .B2( u1_u5_u6_n145 ) , .B1( u1_u5_u6_n146 ) , .ZN( u1_u5_u6_n150 ) );
  INV_X1 u1_u5_u6_U36 (.A( u1_u5_u6_n111 ) , .ZN( u1_u5_u6_n158 ) );
  NAND2_X1 u1_u5_u6_U37 (.ZN( u1_u5_u6_n127 ) , .A1( u1_u5_u6_n91 ) , .A2( u1_u5_u6_n92 ) );
  NAND2_X1 u1_u5_u6_U38 (.ZN( u1_u5_u6_n129 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n96 ) );
  INV_X1 u1_u5_u6_U39 (.A( u1_u5_u6_n144 ) , .ZN( u1_u5_u6_n159 ) );
  INV_X1 u1_u5_u6_U4 (.A( u1_u5_u6_n142 ) , .ZN( u1_u5_u6_n174 ) );
  NAND2_X1 u1_u5_u6_U40 (.ZN( u1_u5_u6_n145 ) , .A2( u1_u5_u6_n97 ) , .A1( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U41 (.ZN( u1_u5_u6_n148 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n94 ) );
  NAND2_X1 u1_u5_u6_U42 (.ZN( u1_u5_u6_n108 ) , .A2( u1_u5_u6_n139 ) , .A1( u1_u5_u6_n144 ) );
  NAND2_X1 u1_u5_u6_U43 (.ZN( u1_u5_u6_n121 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n97 ) );
  NAND2_X1 u1_u5_u6_U44 (.ZN( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n95 ) );
  AND2_X1 u1_u5_u6_U45 (.ZN( u1_u5_u6_n118 ) , .A2( u1_u5_u6_n91 ) , .A1( u1_u5_u6_n99 ) );
  AOI22_X1 u1_u5_u6_U46 (.B2( u1_u5_u6_n110 ) , .B1( u1_u5_u6_n111 ) , .A1( u1_u5_u6_n112 ) , .ZN( u1_u5_u6_n115 ) , .A2( u1_u5_u6_n161 ) );
  NAND4_X1 u1_u5_u6_U47 (.A3( u1_u5_u6_n109 ) , .ZN( u1_u5_u6_n112 ) , .A4( u1_u5_u6_n132 ) , .A2( u1_u5_u6_n147 ) , .A1( u1_u5_u6_n166 ) );
  NOR2_X1 u1_u5_u6_U48 (.ZN( u1_u5_u6_n109 ) , .A1( u1_u5_u6_n170 ) , .A2( u1_u5_u6_n173 ) );
  NAND2_X1 u1_u5_u6_U49 (.ZN( u1_u5_u6_n147 ) , .A2( u1_u5_u6_n98 ) , .A1( u1_u5_u6_n99 ) );
  NAND2_X1 u1_u5_u6_U5 (.A2( u1_u5_u6_n143 ) , .ZN( u1_u5_u6_n152 ) , .A1( u1_u5_u6_n166 ) );
  NAND2_X1 u1_u5_u6_U50 (.ZN( u1_u5_u6_n128 ) , .A1( u1_u5_u6_n94 ) , .A2( u1_u5_u6_n96 ) );
  AOI211_X1 u1_u5_u6_U51 (.B( u1_u5_u6_n134 ) , .A( u1_u5_u6_n135 ) , .C1( u1_u5_u6_n136 ) , .ZN( u1_u5_u6_n137 ) , .C2( u1_u5_u6_n151 ) );
  AOI21_X1 u1_u5_u6_U52 (.B2( u1_u5_u6_n132 ) , .B1( u1_u5_u6_n133 ) , .ZN( u1_u5_u6_n134 ) , .A( u1_u5_u6_n158 ) );
  AOI21_X1 u1_u5_u6_U53 (.B1( u1_u5_u6_n131 ) , .ZN( u1_u5_u6_n135 ) , .A( u1_u5_u6_n144 ) , .B2( u1_u5_u6_n146 ) );
  NAND4_X1 u1_u5_u6_U54 (.A4( u1_u5_u6_n127 ) , .A3( u1_u5_u6_n128 ) , .A2( u1_u5_u6_n129 ) , .A1( u1_u5_u6_n130 ) , .ZN( u1_u5_u6_n136 ) );
  NAND2_X1 u1_u5_u6_U55 (.ZN( u1_u5_u6_n119 ) , .A2( u1_u5_u6_n95 ) , .A1( u1_u5_u6_n99 ) );
  NAND2_X1 u1_u5_u6_U56 (.ZN( u1_u5_u6_n123 ) , .A2( u1_u5_u6_n91 ) , .A1( u1_u5_u6_n96 ) );
  NAND2_X1 u1_u5_u6_U57 (.ZN( u1_u5_u6_n100 ) , .A2( u1_u5_u6_n92 ) , .A1( u1_u5_u6_n98 ) );
  NAND2_X1 u1_u5_u6_U58 (.ZN( u1_u5_u6_n122 ) , .A1( u1_u5_u6_n94 ) , .A2( u1_u5_u6_n97 ) );
  INV_X1 u1_u5_u6_U59 (.A( u1_u5_u6_n139 ) , .ZN( u1_u5_u6_n160 ) );
  AOI22_X1 u1_u5_u6_U6 (.B2( u1_u5_u6_n101 ) , .A1( u1_u5_u6_n102 ) , .ZN( u1_u5_u6_n103 ) , .B1( u1_u5_u6_n160 ) , .A2( u1_u5_u6_n161 ) );
  NAND2_X1 u1_u5_u6_U60 (.ZN( u1_u5_u6_n113 ) , .A1( u1_u5_u6_n96 ) , .A2( u1_u5_u6_n98 ) );
  NOR2_X1 u1_u5_u6_U61 (.A2( u1_u5_X_40 ) , .A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n126 ) );
  NOR2_X1 u1_u5_u6_U62 (.A2( u1_u5_X_39 ) , .A1( u1_u5_X_42 ) , .ZN( u1_u5_u6_n92 ) );
  NOR2_X1 u1_u5_u6_U63 (.A2( u1_u5_X_39 ) , .A1( u1_u5_u6_n156 ) , .ZN( u1_u5_u6_n97 ) );
  NOR2_X1 u1_u5_u6_U64 (.A2( u1_u5_X_38 ) , .A1( u1_u5_u6_n165 ) , .ZN( u1_u5_u6_n95 ) );
  NOR2_X1 u1_u5_u6_U65 (.A2( u1_u5_X_41 ) , .ZN( u1_u5_u6_n111 ) , .A1( u1_u5_u6_n157 ) );
  NOR2_X1 u1_u5_u6_U66 (.A2( u1_u5_X_37 ) , .A1( u1_u5_u6_n162 ) , .ZN( u1_u5_u6_n94 ) );
  NOR2_X1 u1_u5_u6_U67 (.A2( u1_u5_X_37 ) , .A1( u1_u5_X_38 ) , .ZN( u1_u5_u6_n91 ) );
  NAND2_X1 u1_u5_u6_U68 (.A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n144 ) , .A2( u1_u5_u6_n157 ) );
  NAND2_X1 u1_u5_u6_U69 (.A2( u1_u5_X_40 ) , .A1( u1_u5_X_41 ) , .ZN( u1_u5_u6_n139 ) );
  NOR2_X1 u1_u5_u6_U7 (.A1( u1_u5_u6_n118 ) , .ZN( u1_u5_u6_n143 ) , .A2( u1_u5_u6_n168 ) );
  AND2_X1 u1_u5_u6_U70 (.A1( u1_u5_X_39 ) , .A2( u1_u5_u6_n156 ) , .ZN( u1_u5_u6_n96 ) );
  AND2_X1 u1_u5_u6_U71 (.A1( u1_u5_X_39 ) , .A2( u1_u5_X_42 ) , .ZN( u1_u5_u6_n99 ) );
  INV_X1 u1_u5_u6_U72 (.A( u1_u5_X_40 ) , .ZN( u1_u5_u6_n157 ) );
  INV_X1 u1_u5_u6_U73 (.A( u1_u5_X_37 ) , .ZN( u1_u5_u6_n165 ) );
  INV_X1 u1_u5_u6_U74 (.A( u1_u5_X_38 ) , .ZN( u1_u5_u6_n162 ) );
  INV_X1 u1_u5_u6_U75 (.A( u1_u5_X_42 ) , .ZN( u1_u5_u6_n156 ) );
  NAND4_X1 u1_u5_u6_U76 (.ZN( u1_out5_32 ) , .A4( u1_u5_u6_n103 ) , .A3( u1_u5_u6_n104 ) , .A2( u1_u5_u6_n105 ) , .A1( u1_u5_u6_n106 ) );
  AOI22_X1 u1_u5_u6_U77 (.ZN( u1_u5_u6_n105 ) , .A2( u1_u5_u6_n108 ) , .A1( u1_u5_u6_n118 ) , .B2( u1_u5_u6_n126 ) , .B1( u1_u5_u6_n171 ) );
  AOI22_X1 u1_u5_u6_U78 (.ZN( u1_u5_u6_n104 ) , .A1( u1_u5_u6_n111 ) , .B1( u1_u5_u6_n124 ) , .B2( u1_u5_u6_n151 ) , .A2( u1_u5_u6_n93 ) );
  NAND4_X1 u1_u5_u6_U79 (.ZN( u1_out5_12 ) , .A4( u1_u5_u6_n114 ) , .A3( u1_u5_u6_n115 ) , .A2( u1_u5_u6_n116 ) , .A1( u1_u5_u6_n117 ) );
  AOI21_X1 u1_u5_u6_U8 (.B1( u1_u5_u6_n107 ) , .B2( u1_u5_u6_n132 ) , .A( u1_u5_u6_n158 ) , .ZN( u1_u5_u6_n88 ) );
  OAI22_X1 u1_u5_u6_U80 (.B2( u1_u5_u6_n111 ) , .ZN( u1_u5_u6_n116 ) , .B1( u1_u5_u6_n126 ) , .A2( u1_u5_u6_n164 ) , .A1( u1_u5_u6_n167 ) );
  OAI21_X1 u1_u5_u6_U81 (.A( u1_u5_u6_n108 ) , .ZN( u1_u5_u6_n117 ) , .B2( u1_u5_u6_n141 ) , .B1( u1_u5_u6_n163 ) );
  OAI211_X1 u1_u5_u6_U82 (.ZN( u1_out5_7 ) , .B( u1_u5_u6_n153 ) , .C2( u1_u5_u6_n154 ) , .C1( u1_u5_u6_n155 ) , .A( u1_u5_u6_n174 ) );
  NOR3_X1 u1_u5_u6_U83 (.A1( u1_u5_u6_n141 ) , .ZN( u1_u5_u6_n154 ) , .A3( u1_u5_u6_n164 ) , .A2( u1_u5_u6_n171 ) );
  AOI211_X1 u1_u5_u6_U84 (.B( u1_u5_u6_n149 ) , .A( u1_u5_u6_n150 ) , .C2( u1_u5_u6_n151 ) , .C1( u1_u5_u6_n152 ) , .ZN( u1_u5_u6_n153 ) );
  OAI211_X1 u1_u5_u6_U85 (.ZN( u1_out5_22 ) , .B( u1_u5_u6_n137 ) , .A( u1_u5_u6_n138 ) , .C2( u1_u5_u6_n139 ) , .C1( u1_u5_u6_n140 ) );
  AOI22_X1 u1_u5_u6_U86 (.B1( u1_u5_u6_n124 ) , .A2( u1_u5_u6_n125 ) , .A1( u1_u5_u6_n126 ) , .ZN( u1_u5_u6_n138 ) , .B2( u1_u5_u6_n161 ) );
  AND4_X1 u1_u5_u6_U87 (.A3( u1_u5_u6_n119 ) , .A1( u1_u5_u6_n120 ) , .A4( u1_u5_u6_n129 ) , .ZN( u1_u5_u6_n140 ) , .A2( u1_u5_u6_n143 ) );
  NAND3_X1 u1_u5_u6_U88 (.A2( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n125 ) , .A1( u1_u5_u6_n130 ) , .A3( u1_u5_u6_n131 ) );
  NAND3_X1 u1_u5_u6_U89 (.A3( u1_u5_u6_n133 ) , .ZN( u1_u5_u6_n141 ) , .A1( u1_u5_u6_n145 ) , .A2( u1_u5_u6_n148 ) );
  AOI21_X1 u1_u5_u6_U9 (.B2( u1_u5_u6_n147 ) , .B1( u1_u5_u6_n148 ) , .ZN( u1_u5_u6_n149 ) , .A( u1_u5_u6_n158 ) );
  NAND3_X1 u1_u5_u6_U90 (.ZN( u1_u5_u6_n101 ) , .A3( u1_u5_u6_n107 ) , .A2( u1_u5_u6_n121 ) , .A1( u1_u5_u6_n127 ) );
  NAND3_X1 u1_u5_u6_U91 (.ZN( u1_u5_u6_n102 ) , .A3( u1_u5_u6_n130 ) , .A2( u1_u5_u6_n145 ) , .A1( u1_u5_u6_n166 ) );
  NAND3_X1 u1_u5_u6_U92 (.A3( u1_u5_u6_n113 ) , .A1( u1_u5_u6_n119 ) , .A2( u1_u5_u6_n123 ) , .ZN( u1_u5_u6_n93 ) );
  NAND3_X1 u1_u5_u6_U93 (.ZN( u1_u5_u6_n142 ) , .A2( u1_u5_u6_n172 ) , .A3( u1_u5_u6_n89 ) , .A1( u1_u5_u6_n90 ) );
  XOR2_X1 u1_u6_U11 (.B( u1_K7_44 ) , .A( u1_R5_29 ) , .Z( u1_u6_X_44 ) );
  XOR2_X1 u1_u6_U12 (.B( u1_K7_43 ) , .A( u1_R5_28 ) , .Z( u1_u6_X_43 ) );
  XOR2_X1 u1_u6_U13 (.B( u1_K7_42 ) , .A( u1_R5_29 ) , .Z( u1_u6_X_42 ) );
  XOR2_X1 u1_u6_U14 (.B( u1_K7_41 ) , .A( u1_R5_28 ) , .Z( u1_u6_X_41 ) );
  XOR2_X1 u1_u6_U18 (.B( u1_K7_38 ) , .A( u1_R5_25 ) , .Z( u1_u6_X_38 ) );
  XOR2_X1 u1_u6_U19 (.B( u1_K7_37 ) , .A( u1_R5_24 ) , .Z( u1_u6_X_37 ) );
  XOR2_X1 u1_u6_U2 (.B( u1_K7_8 ) , .A( u1_R5_5 ) , .Z( u1_u6_X_8 ) );
  XOR2_X1 u1_u6_U20 (.B( u1_K7_36 ) , .A( u1_R5_25 ) , .Z( u1_u6_X_36 ) );
  XOR2_X1 u1_u6_U21 (.B( u1_K7_35 ) , .A( u1_R5_24 ) , .Z( u1_u6_X_35 ) );
  XOR2_X1 u1_u6_U24 (.B( u1_K7_32 ) , .A( u1_R5_21 ) , .Z( u1_u6_X_32 ) );
  XOR2_X1 u1_u6_U25 (.B( u1_K7_31 ) , .A( u1_R5_20 ) , .Z( u1_u6_X_31 ) );
  XOR2_X1 u1_u6_U26 (.B( u1_K7_30 ) , .A( u1_R5_21 ) , .Z( u1_u6_X_30 ) );
  XOR2_X1 u1_u6_U27 (.B( u1_K7_2 ) , .A( u1_R5_1 ) , .Z( u1_u6_X_2 ) );
  XOR2_X1 u1_u6_U28 (.B( u1_K7_29 ) , .A( u1_R5_20 ) , .Z( u1_u6_X_29 ) );
  XOR2_X1 u1_u6_U3 (.B( u1_K7_7 ) , .A( u1_R5_4 ) , .Z( u1_u6_X_7 ) );
  XOR2_X1 u1_u6_U31 (.B( u1_K7_26 ) , .A( u1_R5_17 ) , .Z( u1_u6_X_26 ) );
  XOR2_X1 u1_u6_U32 (.B( u1_K7_25 ) , .A( u1_R5_16 ) , .Z( u1_u6_X_25 ) );
  XOR2_X1 u1_u6_U33 (.B( u1_K7_24 ) , .A( u1_R5_17 ) , .Z( u1_u6_X_24 ) );
  XOR2_X1 u1_u6_U34 (.B( u1_K7_23 ) , .A( u1_R5_16 ) , .Z( u1_u6_X_23 ) );
  XOR2_X1 u1_u6_U35 (.B( u1_K7_22 ) , .A( u1_R5_15 ) , .Z( u1_u6_X_22 ) );
  XOR2_X1 u1_u6_U36 (.B( u1_K7_21 ) , .A( u1_R5_14 ) , .Z( u1_u6_X_21 ) );
  XOR2_X1 u1_u6_U37 (.B( u1_K7_20 ) , .A( u1_R5_13 ) , .Z( u1_u6_X_20 ) );
  XOR2_X1 u1_u6_U38 (.B( u1_K7_1 ) , .A( u1_R5_32 ) , .Z( u1_u6_X_1 ) );
  XOR2_X1 u1_u6_U39 (.B( u1_K7_19 ) , .A( u1_R5_12 ) , .Z( u1_u6_X_19 ) );
  XOR2_X1 u1_u6_U4 (.B( u1_K7_6 ) , .A( u1_R5_5 ) , .Z( u1_u6_X_6 ) );
  XOR2_X1 u1_u6_U40 (.B( u1_K7_18 ) , .A( u1_R5_13 ) , .Z( u1_u6_X_18 ) );
  XOR2_X1 u1_u6_U41 (.B( u1_K7_17 ) , .A( u1_R5_12 ) , .Z( u1_u6_X_17 ) );
  XOR2_X1 u1_u6_U42 (.B( u1_K7_16 ) , .A( u1_R5_11 ) , .Z( u1_u6_X_16 ) );
  XOR2_X1 u1_u6_U43 (.B( u1_K7_15 ) , .A( u1_R5_10 ) , .Z( u1_u6_X_15 ) );
  XOR2_X1 u1_u6_U44 (.B( u1_K7_14 ) , .A( u1_R5_9 ) , .Z( u1_u6_X_14 ) );
  XOR2_X1 u1_u6_U45 (.B( u1_K7_13 ) , .A( u1_R5_8 ) , .Z( u1_u6_X_13 ) );
  XOR2_X1 u1_u6_U46 (.B( u1_K7_12 ) , .A( u1_R5_9 ) , .Z( u1_u6_X_12 ) );
  XOR2_X1 u1_u6_U47 (.B( u1_K7_11 ) , .A( u1_R5_8 ) , .Z( u1_u6_X_11 ) );
  XOR2_X1 u1_u6_U5 (.B( u1_K7_5 ) , .A( u1_R5_4 ) , .Z( u1_u6_X_5 ) );
  XOR2_X1 u1_u6_U7 (.B( u1_K7_48 ) , .A( u1_R5_1 ) , .Z( u1_u6_X_48 ) );
  XOR2_X1 u1_u6_U8 (.B( u1_K7_47 ) , .A( u1_R5_32 ) , .Z( u1_u6_X_47 ) );
  OAI22_X1 u1_u6_u2_U10 (.B1( u1_u6_u2_n151 ) , .A2( u1_u6_u2_n152 ) , .A1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n160 ) , .B2( u1_u6_u2_n168 ) );
  NAND3_X1 u1_u6_u2_U100 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n98 ) );
  NOR3_X1 u1_u6_u2_U11 (.A1( u1_u6_u2_n150 ) , .ZN( u1_u6_u2_n151 ) , .A3( u1_u6_u2_n175 ) , .A2( u1_u6_u2_n188 ) );
  AOI21_X1 u1_u6_u2_U12 (.B2( u1_u6_u2_n123 ) , .ZN( u1_u6_u2_n125 ) , .A( u1_u6_u2_n171 ) , .B1( u1_u6_u2_n184 ) );
  INV_X1 u1_u6_u2_U13 (.A( u1_u6_u2_n150 ) , .ZN( u1_u6_u2_n184 ) );
  AOI21_X1 u1_u6_u2_U14 (.ZN( u1_u6_u2_n144 ) , .B2( u1_u6_u2_n155 ) , .A( u1_u6_u2_n172 ) , .B1( u1_u6_u2_n185 ) );
  AOI21_X1 u1_u6_u2_U15 (.B2( u1_u6_u2_n143 ) , .ZN( u1_u6_u2_n145 ) , .B1( u1_u6_u2_n152 ) , .A( u1_u6_u2_n171 ) );
  INV_X1 u1_u6_u2_U16 (.A( u1_u6_u2_n156 ) , .ZN( u1_u6_u2_n171 ) );
  INV_X1 u1_u6_u2_U17 (.A( u1_u6_u2_n120 ) , .ZN( u1_u6_u2_n188 ) );
  NAND2_X1 u1_u6_u2_U18 (.A2( u1_u6_u2_n122 ) , .ZN( u1_u6_u2_n150 ) , .A1( u1_u6_u2_n152 ) );
  INV_X1 u1_u6_u2_U19 (.A( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n170 ) );
  INV_X1 u1_u6_u2_U20 (.A( u1_u6_u2_n137 ) , .ZN( u1_u6_u2_n173 ) );
  NAND2_X1 u1_u6_u2_U21 (.A1( u1_u6_u2_n132 ) , .A2( u1_u6_u2_n139 ) , .ZN( u1_u6_u2_n157 ) );
  INV_X1 u1_u6_u2_U22 (.A( u1_u6_u2_n113 ) , .ZN( u1_u6_u2_n178 ) );
  INV_X1 u1_u6_u2_U23 (.A( u1_u6_u2_n139 ) , .ZN( u1_u6_u2_n175 ) );
  INV_X1 u1_u6_u2_U24 (.A( u1_u6_u2_n155 ) , .ZN( u1_u6_u2_n181 ) );
  INV_X1 u1_u6_u2_U25 (.A( u1_u6_u2_n119 ) , .ZN( u1_u6_u2_n177 ) );
  INV_X1 u1_u6_u2_U26 (.A( u1_u6_u2_n116 ) , .ZN( u1_u6_u2_n180 ) );
  INV_X1 u1_u6_u2_U27 (.A( u1_u6_u2_n131 ) , .ZN( u1_u6_u2_n179 ) );
  INV_X1 u1_u6_u2_U28 (.A( u1_u6_u2_n154 ) , .ZN( u1_u6_u2_n176 ) );
  NAND2_X1 u1_u6_u2_U29 (.A2( u1_u6_u2_n116 ) , .A1( u1_u6_u2_n117 ) , .ZN( u1_u6_u2_n118 ) );
  NOR2_X1 u1_u6_u2_U3 (.ZN( u1_u6_u2_n121 ) , .A2( u1_u6_u2_n177 ) , .A1( u1_u6_u2_n180 ) );
  INV_X1 u1_u6_u2_U30 (.A( u1_u6_u2_n132 ) , .ZN( u1_u6_u2_n182 ) );
  INV_X1 u1_u6_u2_U31 (.A( u1_u6_u2_n158 ) , .ZN( u1_u6_u2_n183 ) );
  OAI21_X1 u1_u6_u2_U32 (.A( u1_u6_u2_n156 ) , .B1( u1_u6_u2_n157 ) , .ZN( u1_u6_u2_n158 ) , .B2( u1_u6_u2_n179 ) );
  NOR2_X1 u1_u6_u2_U33 (.ZN( u1_u6_u2_n156 ) , .A1( u1_u6_u2_n166 ) , .A2( u1_u6_u2_n169 ) );
  NOR2_X1 u1_u6_u2_U34 (.A2( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n137 ) , .A1( u1_u6_u2_n140 ) );
  NOR2_X1 u1_u6_u2_U35 (.A2( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n153 ) , .A1( u1_u6_u2_n156 ) );
  AOI211_X1 u1_u6_u2_U36 (.ZN( u1_u6_u2_n130 ) , .C1( u1_u6_u2_n138 ) , .C2( u1_u6_u2_n179 ) , .B( u1_u6_u2_n96 ) , .A( u1_u6_u2_n97 ) );
  OAI22_X1 u1_u6_u2_U37 (.B1( u1_u6_u2_n133 ) , .A2( u1_u6_u2_n137 ) , .A1( u1_u6_u2_n152 ) , .B2( u1_u6_u2_n168 ) , .ZN( u1_u6_u2_n97 ) );
  OAI221_X1 u1_u6_u2_U38 (.B1( u1_u6_u2_n113 ) , .C1( u1_u6_u2_n132 ) , .A( u1_u6_u2_n149 ) , .B2( u1_u6_u2_n171 ) , .C2( u1_u6_u2_n172 ) , .ZN( u1_u6_u2_n96 ) );
  OAI221_X1 u1_u6_u2_U39 (.A( u1_u6_u2_n115 ) , .C2( u1_u6_u2_n123 ) , .B2( u1_u6_u2_n143 ) , .B1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n163 ) , .C1( u1_u6_u2_n168 ) );
  INV_X1 u1_u6_u2_U4 (.A( u1_u6_u2_n134 ) , .ZN( u1_u6_u2_n185 ) );
  OAI21_X1 u1_u6_u2_U40 (.A( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n115 ) , .B1( u1_u6_u2_n176 ) , .B2( u1_u6_u2_n178 ) );
  OAI221_X1 u1_u6_u2_U41 (.A( u1_u6_u2_n135 ) , .B2( u1_u6_u2_n136 ) , .B1( u1_u6_u2_n137 ) , .ZN( u1_u6_u2_n162 ) , .C2( u1_u6_u2_n167 ) , .C1( u1_u6_u2_n185 ) );
  AND3_X1 u1_u6_u2_U42 (.A3( u1_u6_u2_n131 ) , .A2( u1_u6_u2_n132 ) , .A1( u1_u6_u2_n133 ) , .ZN( u1_u6_u2_n136 ) );
  AOI22_X1 u1_u6_u2_U43 (.ZN( u1_u6_u2_n135 ) , .B1( u1_u6_u2_n140 ) , .A1( u1_u6_u2_n156 ) , .B2( u1_u6_u2_n180 ) , .A2( u1_u6_u2_n188 ) );
  AOI21_X1 u1_u6_u2_U44 (.ZN( u1_u6_u2_n149 ) , .B1( u1_u6_u2_n173 ) , .B2( u1_u6_u2_n188 ) , .A( u1_u6_u2_n95 ) );
  AND3_X1 u1_u6_u2_U45 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n156 ) , .ZN( u1_u6_u2_n95 ) );
  OAI21_X1 u1_u6_u2_U46 (.A( u1_u6_u2_n101 ) , .B2( u1_u6_u2_n121 ) , .B1( u1_u6_u2_n153 ) , .ZN( u1_u6_u2_n164 ) );
  NAND2_X1 u1_u6_u2_U47 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n155 ) );
  NAND2_X1 u1_u6_u2_U48 (.A2( u1_u6_u2_n105 ) , .A1( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n143 ) );
  NAND2_X1 u1_u6_u2_U49 (.A1( u1_u6_u2_n104 ) , .A2( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n152 ) );
  NOR4_X1 u1_u6_u2_U5 (.A4( u1_u6_u2_n124 ) , .A3( u1_u6_u2_n125 ) , .A2( u1_u6_u2_n126 ) , .A1( u1_u6_u2_n127 ) , .ZN( u1_u6_u2_n128 ) );
  NAND2_X1 u1_u6_u2_U50 (.A1( u1_u6_u2_n100 ) , .A2( u1_u6_u2_n105 ) , .ZN( u1_u6_u2_n132 ) );
  INV_X1 u1_u6_u2_U51 (.A( u1_u6_u2_n140 ) , .ZN( u1_u6_u2_n168 ) );
  INV_X1 u1_u6_u2_U52 (.A( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n167 ) );
  OAI21_X1 u1_u6_u2_U53 (.A( u1_u6_u2_n141 ) , .B2( u1_u6_u2_n142 ) , .ZN( u1_u6_u2_n146 ) , .B1( u1_u6_u2_n153 ) );
  OAI21_X1 u1_u6_u2_U54 (.A( u1_u6_u2_n140 ) , .ZN( u1_u6_u2_n141 ) , .B1( u1_u6_u2_n176 ) , .B2( u1_u6_u2_n177 ) );
  NOR3_X1 u1_u6_u2_U55 (.ZN( u1_u6_u2_n142 ) , .A3( u1_u6_u2_n175 ) , .A2( u1_u6_u2_n178 ) , .A1( u1_u6_u2_n181 ) );
  NAND2_X1 u1_u6_u2_U56 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n113 ) );
  NAND2_X1 u1_u6_u2_U57 (.A1( u1_u6_u2_n106 ) , .A2( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n131 ) );
  NAND2_X1 u1_u6_u2_U58 (.A1( u1_u6_u2_n103 ) , .A2( u1_u6_u2_n107 ) , .ZN( u1_u6_u2_n139 ) );
  NAND2_X1 u1_u6_u2_U59 (.A1( u1_u6_u2_n103 ) , .A2( u1_u6_u2_n105 ) , .ZN( u1_u6_u2_n133 ) );
  AOI21_X1 u1_u6_u2_U6 (.B2( u1_u6_u2_n119 ) , .ZN( u1_u6_u2_n127 ) , .A( u1_u6_u2_n137 ) , .B1( u1_u6_u2_n155 ) );
  NAND2_X1 u1_u6_u2_U60 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n103 ) , .ZN( u1_u6_u2_n154 ) );
  NAND2_X1 u1_u6_u2_U61 (.A2( u1_u6_u2_n103 ) , .A1( u1_u6_u2_n104 ) , .ZN( u1_u6_u2_n119 ) );
  NAND2_X1 u1_u6_u2_U62 (.A2( u1_u6_u2_n107 ) , .A1( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n123 ) );
  NAND2_X1 u1_u6_u2_U63 (.A1( u1_u6_u2_n104 ) , .A2( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n122 ) );
  INV_X1 u1_u6_u2_U64 (.A( u1_u6_u2_n114 ) , .ZN( u1_u6_u2_n172 ) );
  NAND2_X1 u1_u6_u2_U65 (.A2( u1_u6_u2_n100 ) , .A1( u1_u6_u2_n102 ) , .ZN( u1_u6_u2_n116 ) );
  NAND2_X1 u1_u6_u2_U66 (.A1( u1_u6_u2_n102 ) , .A2( u1_u6_u2_n108 ) , .ZN( u1_u6_u2_n120 ) );
  NAND2_X1 u1_u6_u2_U67 (.A2( u1_u6_u2_n105 ) , .A1( u1_u6_u2_n106 ) , .ZN( u1_u6_u2_n117 ) );
  INV_X1 u1_u6_u2_U68 (.ZN( u1_u6_u2_n187 ) , .A( u1_u6_u2_n99 ) );
  OAI21_X1 u1_u6_u2_U69 (.B1( u1_u6_u2_n137 ) , .B2( u1_u6_u2_n143 ) , .A( u1_u6_u2_n98 ) , .ZN( u1_u6_u2_n99 ) );
  AOI21_X1 u1_u6_u2_U7 (.ZN( u1_u6_u2_n124 ) , .B1( u1_u6_u2_n131 ) , .B2( u1_u6_u2_n143 ) , .A( u1_u6_u2_n172 ) );
  NOR2_X1 u1_u6_u2_U70 (.A2( u1_u6_X_16 ) , .ZN( u1_u6_u2_n140 ) , .A1( u1_u6_u2_n166 ) );
  NOR2_X1 u1_u6_u2_U71 (.A2( u1_u6_X_13 ) , .A1( u1_u6_X_14 ) , .ZN( u1_u6_u2_n100 ) );
  NOR2_X1 u1_u6_u2_U72 (.A2( u1_u6_X_16 ) , .A1( u1_u6_X_17 ) , .ZN( u1_u6_u2_n138 ) );
  NOR2_X1 u1_u6_u2_U73 (.A2( u1_u6_X_15 ) , .A1( u1_u6_X_18 ) , .ZN( u1_u6_u2_n104 ) );
  NOR2_X1 u1_u6_u2_U74 (.A2( u1_u6_X_14 ) , .ZN( u1_u6_u2_n103 ) , .A1( u1_u6_u2_n174 ) );
  NOR2_X1 u1_u6_u2_U75 (.A2( u1_u6_X_15 ) , .ZN( u1_u6_u2_n102 ) , .A1( u1_u6_u2_n165 ) );
  NOR2_X1 u1_u6_u2_U76 (.A2( u1_u6_X_17 ) , .ZN( u1_u6_u2_n114 ) , .A1( u1_u6_u2_n169 ) );
  AND2_X1 u1_u6_u2_U77 (.A1( u1_u6_X_15 ) , .ZN( u1_u6_u2_n105 ) , .A2( u1_u6_u2_n165 ) );
  AND2_X1 u1_u6_u2_U78 (.A2( u1_u6_X_15 ) , .A1( u1_u6_X_18 ) , .ZN( u1_u6_u2_n107 ) );
  AND2_X1 u1_u6_u2_U79 (.A1( u1_u6_X_14 ) , .ZN( u1_u6_u2_n106 ) , .A2( u1_u6_u2_n174 ) );
  AOI21_X1 u1_u6_u2_U8 (.B2( u1_u6_u2_n120 ) , .B1( u1_u6_u2_n121 ) , .ZN( u1_u6_u2_n126 ) , .A( u1_u6_u2_n167 ) );
  AND2_X1 u1_u6_u2_U80 (.A1( u1_u6_X_13 ) , .A2( u1_u6_X_14 ) , .ZN( u1_u6_u2_n108 ) );
  INV_X1 u1_u6_u2_U81 (.A( u1_u6_X_16 ) , .ZN( u1_u6_u2_n169 ) );
  INV_X1 u1_u6_u2_U82 (.A( u1_u6_X_17 ) , .ZN( u1_u6_u2_n166 ) );
  INV_X1 u1_u6_u2_U83 (.A( u1_u6_X_13 ) , .ZN( u1_u6_u2_n174 ) );
  INV_X1 u1_u6_u2_U84 (.A( u1_u6_X_18 ) , .ZN( u1_u6_u2_n165 ) );
  NAND4_X1 u1_u6_u2_U85 (.ZN( u1_out6_16 ) , .A4( u1_u6_u2_n128 ) , .A3( u1_u6_u2_n129 ) , .A1( u1_u6_u2_n130 ) , .A2( u1_u6_u2_n186 ) );
  AOI22_X1 u1_u6_u2_U86 (.A2( u1_u6_u2_n118 ) , .ZN( u1_u6_u2_n129 ) , .A1( u1_u6_u2_n140 ) , .B1( u1_u6_u2_n157 ) , .B2( u1_u6_u2_n170 ) );
  INV_X1 u1_u6_u2_U87 (.A( u1_u6_u2_n163 ) , .ZN( u1_u6_u2_n186 ) );
  NAND4_X1 u1_u6_u2_U88 (.ZN( u1_out6_24 ) , .A4( u1_u6_u2_n111 ) , .A3( u1_u6_u2_n112 ) , .A1( u1_u6_u2_n130 ) , .A2( u1_u6_u2_n187 ) );
  AOI221_X1 u1_u6_u2_U89 (.A( u1_u6_u2_n109 ) , .B1( u1_u6_u2_n110 ) , .ZN( u1_u6_u2_n111 ) , .C1( u1_u6_u2_n134 ) , .C2( u1_u6_u2_n170 ) , .B2( u1_u6_u2_n173 ) );
  OAI22_X1 u1_u6_u2_U9 (.ZN( u1_u6_u2_n109 ) , .A2( u1_u6_u2_n113 ) , .B2( u1_u6_u2_n133 ) , .B1( u1_u6_u2_n167 ) , .A1( u1_u6_u2_n168 ) );
  AOI21_X1 u1_u6_u2_U90 (.ZN( u1_u6_u2_n112 ) , .B2( u1_u6_u2_n156 ) , .A( u1_u6_u2_n164 ) , .B1( u1_u6_u2_n181 ) );
  NAND4_X1 u1_u6_u2_U91 (.ZN( u1_out6_30 ) , .A4( u1_u6_u2_n147 ) , .A3( u1_u6_u2_n148 ) , .A2( u1_u6_u2_n149 ) , .A1( u1_u6_u2_n187 ) );
  AOI21_X1 u1_u6_u2_U92 (.B2( u1_u6_u2_n138 ) , .ZN( u1_u6_u2_n148 ) , .A( u1_u6_u2_n162 ) , .B1( u1_u6_u2_n182 ) );
  NOR3_X1 u1_u6_u2_U93 (.A3( u1_u6_u2_n144 ) , .A2( u1_u6_u2_n145 ) , .A1( u1_u6_u2_n146 ) , .ZN( u1_u6_u2_n147 ) );
  OR4_X1 u1_u6_u2_U94 (.ZN( u1_out6_6 ) , .A4( u1_u6_u2_n161 ) , .A3( u1_u6_u2_n162 ) , .A2( u1_u6_u2_n163 ) , .A1( u1_u6_u2_n164 ) );
  OR3_X1 u1_u6_u2_U95 (.A2( u1_u6_u2_n159 ) , .A1( u1_u6_u2_n160 ) , .ZN( u1_u6_u2_n161 ) , .A3( u1_u6_u2_n183 ) );
  AOI21_X1 u1_u6_u2_U96 (.B2( u1_u6_u2_n154 ) , .B1( u1_u6_u2_n155 ) , .ZN( u1_u6_u2_n159 ) , .A( u1_u6_u2_n167 ) );
  NAND3_X1 u1_u6_u2_U97 (.A2( u1_u6_u2_n117 ) , .A1( u1_u6_u2_n122 ) , .A3( u1_u6_u2_n123 ) , .ZN( u1_u6_u2_n134 ) );
  NAND3_X1 u1_u6_u2_U98 (.ZN( u1_u6_u2_n110 ) , .A2( u1_u6_u2_n131 ) , .A3( u1_u6_u2_n139 ) , .A1( u1_u6_u2_n154 ) );
  NAND3_X1 u1_u6_u2_U99 (.A2( u1_u6_u2_n100 ) , .ZN( u1_u6_u2_n101 ) , .A1( u1_u6_u2_n104 ) , .A3( u1_u6_u2_n114 ) );
  OAI22_X1 u1_u6_u3_U10 (.B1( u1_u6_u3_n113 ) , .A2( u1_u6_u3_n135 ) , .A1( u1_u6_u3_n150 ) , .B2( u1_u6_u3_n164 ) , .ZN( u1_u6_u3_n98 ) );
  OAI211_X1 u1_u6_u3_U11 (.B( u1_u6_u3_n106 ) , .ZN( u1_u6_u3_n119 ) , .C2( u1_u6_u3_n128 ) , .C1( u1_u6_u3_n167 ) , .A( u1_u6_u3_n181 ) );
  AOI221_X1 u1_u6_u3_U12 (.C1( u1_u6_u3_n105 ) , .ZN( u1_u6_u3_n106 ) , .A( u1_u6_u3_n131 ) , .B2( u1_u6_u3_n132 ) , .C2( u1_u6_u3_n133 ) , .B1( u1_u6_u3_n169 ) );
  INV_X1 u1_u6_u3_U13 (.ZN( u1_u6_u3_n181 ) , .A( u1_u6_u3_n98 ) );
  NAND2_X1 u1_u6_u3_U14 (.ZN( u1_u6_u3_n105 ) , .A2( u1_u6_u3_n130 ) , .A1( u1_u6_u3_n155 ) );
  AOI22_X1 u1_u6_u3_U15 (.B1( u1_u6_u3_n115 ) , .A2( u1_u6_u3_n116 ) , .ZN( u1_u6_u3_n123 ) , .B2( u1_u6_u3_n133 ) , .A1( u1_u6_u3_n169 ) );
  NAND2_X1 u1_u6_u3_U16 (.ZN( u1_u6_u3_n116 ) , .A2( u1_u6_u3_n151 ) , .A1( u1_u6_u3_n182 ) );
  NOR2_X1 u1_u6_u3_U17 (.ZN( u1_u6_u3_n126 ) , .A2( u1_u6_u3_n150 ) , .A1( u1_u6_u3_n164 ) );
  AOI21_X1 u1_u6_u3_U18 (.ZN( u1_u6_u3_n112 ) , .B2( u1_u6_u3_n146 ) , .B1( u1_u6_u3_n155 ) , .A( u1_u6_u3_n167 ) );
  NAND2_X1 u1_u6_u3_U19 (.A1( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n142 ) , .A2( u1_u6_u3_n164 ) );
  NAND2_X1 u1_u6_u3_U20 (.ZN( u1_u6_u3_n132 ) , .A2( u1_u6_u3_n152 ) , .A1( u1_u6_u3_n156 ) );
  AND2_X1 u1_u6_u3_U21 (.A2( u1_u6_u3_n113 ) , .A1( u1_u6_u3_n114 ) , .ZN( u1_u6_u3_n151 ) );
  INV_X1 u1_u6_u3_U22 (.A( u1_u6_u3_n133 ) , .ZN( u1_u6_u3_n165 ) );
  INV_X1 u1_u6_u3_U23 (.A( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n170 ) );
  NAND2_X1 u1_u6_u3_U24 (.A1( u1_u6_u3_n107 ) , .A2( u1_u6_u3_n108 ) , .ZN( u1_u6_u3_n140 ) );
  NAND2_X1 u1_u6_u3_U25 (.ZN( u1_u6_u3_n117 ) , .A1( u1_u6_u3_n124 ) , .A2( u1_u6_u3_n148 ) );
  NAND2_X1 u1_u6_u3_U26 (.ZN( u1_u6_u3_n143 ) , .A1( u1_u6_u3_n165 ) , .A2( u1_u6_u3_n167 ) );
  INV_X1 u1_u6_u3_U27 (.A( u1_u6_u3_n130 ) , .ZN( u1_u6_u3_n177 ) );
  INV_X1 u1_u6_u3_U28 (.A( u1_u6_u3_n128 ) , .ZN( u1_u6_u3_n176 ) );
  INV_X1 u1_u6_u3_U29 (.A( u1_u6_u3_n155 ) , .ZN( u1_u6_u3_n174 ) );
  INV_X1 u1_u6_u3_U3 (.A( u1_u6_u3_n129 ) , .ZN( u1_u6_u3_n183 ) );
  INV_X1 u1_u6_u3_U30 (.A( u1_u6_u3_n139 ) , .ZN( u1_u6_u3_n185 ) );
  NOR2_X1 u1_u6_u3_U31 (.ZN( u1_u6_u3_n135 ) , .A2( u1_u6_u3_n141 ) , .A1( u1_u6_u3_n169 ) );
  OAI222_X1 u1_u6_u3_U32 (.C2( u1_u6_u3_n107 ) , .A2( u1_u6_u3_n108 ) , .B1( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n138 ) , .B2( u1_u6_u3_n146 ) , .C1( u1_u6_u3_n154 ) , .A1( u1_u6_u3_n164 ) );
  NOR4_X1 u1_u6_u3_U33 (.A4( u1_u6_u3_n157 ) , .A3( u1_u6_u3_n158 ) , .A2( u1_u6_u3_n159 ) , .A1( u1_u6_u3_n160 ) , .ZN( u1_u6_u3_n161 ) );
  AOI21_X1 u1_u6_u3_U34 (.B2( u1_u6_u3_n152 ) , .B1( u1_u6_u3_n153 ) , .ZN( u1_u6_u3_n158 ) , .A( u1_u6_u3_n164 ) );
  AOI21_X1 u1_u6_u3_U35 (.A( u1_u6_u3_n154 ) , .B2( u1_u6_u3_n155 ) , .B1( u1_u6_u3_n156 ) , .ZN( u1_u6_u3_n157 ) );
  AOI21_X1 u1_u6_u3_U36 (.A( u1_u6_u3_n149 ) , .B2( u1_u6_u3_n150 ) , .B1( u1_u6_u3_n151 ) , .ZN( u1_u6_u3_n159 ) );
  AOI211_X1 u1_u6_u3_U37 (.ZN( u1_u6_u3_n109 ) , .A( u1_u6_u3_n119 ) , .C2( u1_u6_u3_n129 ) , .B( u1_u6_u3_n138 ) , .C1( u1_u6_u3_n141 ) );
  AOI211_X1 u1_u6_u3_U38 (.B( u1_u6_u3_n119 ) , .A( u1_u6_u3_n120 ) , .C2( u1_u6_u3_n121 ) , .ZN( u1_u6_u3_n122 ) , .C1( u1_u6_u3_n179 ) );
  INV_X1 u1_u6_u3_U39 (.A( u1_u6_u3_n156 ) , .ZN( u1_u6_u3_n179 ) );
  INV_X1 u1_u6_u3_U4 (.A( u1_u6_u3_n140 ) , .ZN( u1_u6_u3_n182 ) );
  OAI22_X1 u1_u6_u3_U40 (.B1( u1_u6_u3_n118 ) , .ZN( u1_u6_u3_n120 ) , .A1( u1_u6_u3_n135 ) , .B2( u1_u6_u3_n154 ) , .A2( u1_u6_u3_n178 ) );
  AND3_X1 u1_u6_u3_U41 (.ZN( u1_u6_u3_n118 ) , .A2( u1_u6_u3_n124 ) , .A1( u1_u6_u3_n144 ) , .A3( u1_u6_u3_n152 ) );
  INV_X1 u1_u6_u3_U42 (.A( u1_u6_u3_n121 ) , .ZN( u1_u6_u3_n164 ) );
  NAND2_X1 u1_u6_u3_U43 (.ZN( u1_u6_u3_n133 ) , .A1( u1_u6_u3_n154 ) , .A2( u1_u6_u3_n164 ) );
  OAI211_X1 u1_u6_u3_U44 (.B( u1_u6_u3_n127 ) , .ZN( u1_u6_u3_n139 ) , .C1( u1_u6_u3_n150 ) , .C2( u1_u6_u3_n154 ) , .A( u1_u6_u3_n184 ) );
  INV_X1 u1_u6_u3_U45 (.A( u1_u6_u3_n125 ) , .ZN( u1_u6_u3_n184 ) );
  AOI221_X1 u1_u6_u3_U46 (.A( u1_u6_u3_n126 ) , .ZN( u1_u6_u3_n127 ) , .C2( u1_u6_u3_n132 ) , .C1( u1_u6_u3_n169 ) , .B2( u1_u6_u3_n170 ) , .B1( u1_u6_u3_n174 ) );
  OAI22_X1 u1_u6_u3_U47 (.A1( u1_u6_u3_n124 ) , .ZN( u1_u6_u3_n125 ) , .B2( u1_u6_u3_n145 ) , .A2( u1_u6_u3_n165 ) , .B1( u1_u6_u3_n167 ) );
  NOR2_X1 u1_u6_u3_U48 (.A1( u1_u6_u3_n113 ) , .ZN( u1_u6_u3_n131 ) , .A2( u1_u6_u3_n154 ) );
  NAND2_X1 u1_u6_u3_U49 (.A1( u1_u6_u3_n103 ) , .ZN( u1_u6_u3_n150 ) , .A2( u1_u6_u3_n99 ) );
  INV_X1 u1_u6_u3_U5 (.A( u1_u6_u3_n117 ) , .ZN( u1_u6_u3_n178 ) );
  NAND2_X1 u1_u6_u3_U50 (.A2( u1_u6_u3_n102 ) , .ZN( u1_u6_u3_n155 ) , .A1( u1_u6_u3_n97 ) );
  INV_X1 u1_u6_u3_U51 (.A( u1_u6_u3_n141 ) , .ZN( u1_u6_u3_n167 ) );
  AOI21_X1 u1_u6_u3_U52 (.B2( u1_u6_u3_n114 ) , .B1( u1_u6_u3_n146 ) , .A( u1_u6_u3_n154 ) , .ZN( u1_u6_u3_n94 ) );
  AOI21_X1 u1_u6_u3_U53 (.ZN( u1_u6_u3_n110 ) , .B2( u1_u6_u3_n142 ) , .B1( u1_u6_u3_n186 ) , .A( u1_u6_u3_n95 ) );
  INV_X1 u1_u6_u3_U54 (.A( u1_u6_u3_n145 ) , .ZN( u1_u6_u3_n186 ) );
  AOI21_X1 u1_u6_u3_U55 (.B1( u1_u6_u3_n124 ) , .A( u1_u6_u3_n149 ) , .B2( u1_u6_u3_n155 ) , .ZN( u1_u6_u3_n95 ) );
  INV_X1 u1_u6_u3_U56 (.A( u1_u6_u3_n149 ) , .ZN( u1_u6_u3_n169 ) );
  NAND2_X1 u1_u6_u3_U57 (.ZN( u1_u6_u3_n124 ) , .A1( u1_u6_u3_n96 ) , .A2( u1_u6_u3_n97 ) );
  NAND2_X1 u1_u6_u3_U58 (.A2( u1_u6_u3_n100 ) , .ZN( u1_u6_u3_n146 ) , .A1( u1_u6_u3_n96 ) );
  NAND2_X1 u1_u6_u3_U59 (.A1( u1_u6_u3_n101 ) , .ZN( u1_u6_u3_n145 ) , .A2( u1_u6_u3_n99 ) );
  AOI221_X1 u1_u6_u3_U6 (.A( u1_u6_u3_n131 ) , .C2( u1_u6_u3_n132 ) , .C1( u1_u6_u3_n133 ) , .ZN( u1_u6_u3_n134 ) , .B1( u1_u6_u3_n143 ) , .B2( u1_u6_u3_n177 ) );
  NAND2_X1 u1_u6_u3_U60 (.A1( u1_u6_u3_n100 ) , .ZN( u1_u6_u3_n156 ) , .A2( u1_u6_u3_n99 ) );
  NAND2_X1 u1_u6_u3_U61 (.A2( u1_u6_u3_n101 ) , .A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n148 ) );
  NAND2_X1 u1_u6_u3_U62 (.A1( u1_u6_u3_n100 ) , .A2( u1_u6_u3_n102 ) , .ZN( u1_u6_u3_n128 ) );
  NAND2_X1 u1_u6_u3_U63 (.A2( u1_u6_u3_n101 ) , .A1( u1_u6_u3_n102 ) , .ZN( u1_u6_u3_n152 ) );
  NAND2_X1 u1_u6_u3_U64 (.A2( u1_u6_u3_n101 ) , .ZN( u1_u6_u3_n114 ) , .A1( u1_u6_u3_n96 ) );
  NAND2_X1 u1_u6_u3_U65 (.ZN( u1_u6_u3_n107 ) , .A1( u1_u6_u3_n97 ) , .A2( u1_u6_u3_n99 ) );
  NAND2_X1 u1_u6_u3_U66 (.A2( u1_u6_u3_n100 ) , .A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n113 ) );
  NAND2_X1 u1_u6_u3_U67 (.A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n153 ) , .A2( u1_u6_u3_n97 ) );
  NAND2_X1 u1_u6_u3_U68 (.A2( u1_u6_u3_n103 ) , .A1( u1_u6_u3_n104 ) , .ZN( u1_u6_u3_n130 ) );
  NAND2_X1 u1_u6_u3_U69 (.A2( u1_u6_u3_n103 ) , .ZN( u1_u6_u3_n144 ) , .A1( u1_u6_u3_n96 ) );
  OAI22_X1 u1_u6_u3_U7 (.B2( u1_u6_u3_n147 ) , .A2( u1_u6_u3_n148 ) , .ZN( u1_u6_u3_n160 ) , .B1( u1_u6_u3_n165 ) , .A1( u1_u6_u3_n168 ) );
  NAND2_X1 u1_u6_u3_U70 (.A1( u1_u6_u3_n102 ) , .A2( u1_u6_u3_n103 ) , .ZN( u1_u6_u3_n108 ) );
  NOR2_X1 u1_u6_u3_U71 (.A2( u1_u6_X_19 ) , .A1( u1_u6_X_20 ) , .ZN( u1_u6_u3_n99 ) );
  NOR2_X1 u1_u6_u3_U72 (.A2( u1_u6_X_21 ) , .A1( u1_u6_X_24 ) , .ZN( u1_u6_u3_n103 ) );
  NOR2_X1 u1_u6_u3_U73 (.A2( u1_u6_X_24 ) , .A1( u1_u6_u3_n171 ) , .ZN( u1_u6_u3_n97 ) );
  NOR2_X1 u1_u6_u3_U74 (.A2( u1_u6_X_23 ) , .ZN( u1_u6_u3_n141 ) , .A1( u1_u6_u3_n166 ) );
  NOR2_X1 u1_u6_u3_U75 (.A2( u1_u6_X_19 ) , .A1( u1_u6_u3_n172 ) , .ZN( u1_u6_u3_n96 ) );
  NAND2_X1 u1_u6_u3_U76 (.A1( u1_u6_X_22 ) , .A2( u1_u6_X_23 ) , .ZN( u1_u6_u3_n154 ) );
  NAND2_X1 u1_u6_u3_U77 (.A1( u1_u6_X_23 ) , .ZN( u1_u6_u3_n149 ) , .A2( u1_u6_u3_n166 ) );
  NOR2_X1 u1_u6_u3_U78 (.A2( u1_u6_X_22 ) , .A1( u1_u6_X_23 ) , .ZN( u1_u6_u3_n121 ) );
  AND2_X1 u1_u6_u3_U79 (.A1( u1_u6_X_24 ) , .ZN( u1_u6_u3_n101 ) , .A2( u1_u6_u3_n171 ) );
  AND3_X1 u1_u6_u3_U8 (.A3( u1_u6_u3_n144 ) , .A2( u1_u6_u3_n145 ) , .A1( u1_u6_u3_n146 ) , .ZN( u1_u6_u3_n147 ) );
  AND2_X1 u1_u6_u3_U80 (.A1( u1_u6_X_19 ) , .ZN( u1_u6_u3_n102 ) , .A2( u1_u6_u3_n172 ) );
  AND2_X1 u1_u6_u3_U81 (.A1( u1_u6_X_21 ) , .A2( u1_u6_X_24 ) , .ZN( u1_u6_u3_n100 ) );
  AND2_X1 u1_u6_u3_U82 (.A2( u1_u6_X_19 ) , .A1( u1_u6_X_20 ) , .ZN( u1_u6_u3_n104 ) );
  INV_X1 u1_u6_u3_U83 (.A( u1_u6_X_22 ) , .ZN( u1_u6_u3_n166 ) );
  INV_X1 u1_u6_u3_U84 (.A( u1_u6_X_21 ) , .ZN( u1_u6_u3_n171 ) );
  INV_X1 u1_u6_u3_U85 (.A( u1_u6_X_20 ) , .ZN( u1_u6_u3_n172 ) );
  NAND4_X1 u1_u6_u3_U86 (.ZN( u1_out6_20 ) , .A4( u1_u6_u3_n122 ) , .A3( u1_u6_u3_n123 ) , .A1( u1_u6_u3_n175 ) , .A2( u1_u6_u3_n180 ) );
  INV_X1 u1_u6_u3_U87 (.A( u1_u6_u3_n126 ) , .ZN( u1_u6_u3_n180 ) );
  INV_X1 u1_u6_u3_U88 (.A( u1_u6_u3_n112 ) , .ZN( u1_u6_u3_n175 ) );
  NAND4_X1 u1_u6_u3_U89 (.ZN( u1_out6_26 ) , .A4( u1_u6_u3_n109 ) , .A3( u1_u6_u3_n110 ) , .A2( u1_u6_u3_n111 ) , .A1( u1_u6_u3_n173 ) );
  INV_X1 u1_u6_u3_U9 (.A( u1_u6_u3_n143 ) , .ZN( u1_u6_u3_n168 ) );
  INV_X1 u1_u6_u3_U90 (.ZN( u1_u6_u3_n173 ) , .A( u1_u6_u3_n94 ) );
  OAI21_X1 u1_u6_u3_U91 (.ZN( u1_u6_u3_n111 ) , .B2( u1_u6_u3_n117 ) , .A( u1_u6_u3_n133 ) , .B1( u1_u6_u3_n176 ) );
  NAND4_X1 u1_u6_u3_U92 (.ZN( u1_out6_1 ) , .A4( u1_u6_u3_n161 ) , .A3( u1_u6_u3_n162 ) , .A2( u1_u6_u3_n163 ) , .A1( u1_u6_u3_n185 ) );
  NAND2_X1 u1_u6_u3_U93 (.ZN( u1_u6_u3_n163 ) , .A2( u1_u6_u3_n170 ) , .A1( u1_u6_u3_n176 ) );
  AOI22_X1 u1_u6_u3_U94 (.B2( u1_u6_u3_n140 ) , .B1( u1_u6_u3_n141 ) , .A2( u1_u6_u3_n142 ) , .ZN( u1_u6_u3_n162 ) , .A1( u1_u6_u3_n177 ) );
  OR4_X1 u1_u6_u3_U95 (.ZN( u1_out6_10 ) , .A4( u1_u6_u3_n136 ) , .A3( u1_u6_u3_n137 ) , .A1( u1_u6_u3_n138 ) , .A2( u1_u6_u3_n139 ) );
  OAI222_X1 u1_u6_u3_U96 (.C1( u1_u6_u3_n128 ) , .ZN( u1_u6_u3_n137 ) , .B1( u1_u6_u3_n148 ) , .A2( u1_u6_u3_n150 ) , .B2( u1_u6_u3_n154 ) , .C2( u1_u6_u3_n164 ) , .A1( u1_u6_u3_n167 ) );
  OAI221_X1 u1_u6_u3_U97 (.A( u1_u6_u3_n134 ) , .B2( u1_u6_u3_n135 ) , .ZN( u1_u6_u3_n136 ) , .C1( u1_u6_u3_n149 ) , .B1( u1_u6_u3_n151 ) , .C2( u1_u6_u3_n183 ) );
  NAND3_X1 u1_u6_u3_U98 (.A1( u1_u6_u3_n114 ) , .ZN( u1_u6_u3_n115 ) , .A2( u1_u6_u3_n145 ) , .A3( u1_u6_u3_n153 ) );
  NAND3_X1 u1_u6_u3_U99 (.ZN( u1_u6_u3_n129 ) , .A2( u1_u6_u3_n144 ) , .A1( u1_u6_u3_n153 ) , .A3( u1_u6_u3_n182 ) );
  XOR2_X1 u1_u7_U1 (.B( u1_K8_9 ) , .A( u1_R6_6 ) , .Z( u1_u7_X_9 ) );
  XOR2_X1 u1_u7_U11 (.B( u1_K8_44 ) , .A( u1_R6_29 ) , .Z( u1_u7_X_44 ) );
  XOR2_X1 u1_u7_U12 (.B( u1_K8_43 ) , .A( u1_R6_28 ) , .Z( u1_u7_X_43 ) );
  XOR2_X1 u1_u7_U13 (.B( u1_K8_42 ) , .A( u1_R6_29 ) , .Z( u1_u7_X_42 ) );
  XOR2_X1 u1_u7_U14 (.B( u1_K8_41 ) , .A( u1_R6_28 ) , .Z( u1_u7_X_41 ) );
  XOR2_X1 u1_u7_U15 (.B( u1_K8_40 ) , .A( u1_R6_27 ) , .Z( u1_u7_X_40 ) );
  XOR2_X1 u1_u7_U16 (.B( u1_K8_3 ) , .A( u1_R6_2 ) , .Z( u1_u7_X_3 ) );
  XOR2_X1 u1_u7_U17 (.B( u1_K8_39 ) , .A( u1_R6_26 ) , .Z( u1_u7_X_39 ) );
  XOR2_X1 u1_u7_U18 (.B( u1_K8_38 ) , .A( u1_R6_25 ) , .Z( u1_u7_X_38 ) );
  XOR2_X1 u1_u7_U19 (.B( u1_K8_37 ) , .A( u1_R6_24 ) , .Z( u1_u7_X_37 ) );
  XOR2_X1 u1_u7_U2 (.B( u1_K8_8 ) , .A( u1_R6_5 ) , .Z( u1_u7_X_8 ) );
  XOR2_X1 u1_u7_U20 (.B( u1_K8_36 ) , .A( u1_R6_25 ) , .Z( u1_u7_X_36 ) );
  XOR2_X1 u1_u7_U21 (.B( u1_K8_35 ) , .A( u1_R6_24 ) , .Z( u1_u7_X_35 ) );
  XOR2_X1 u1_u7_U24 (.B( u1_K8_32 ) , .A( u1_R6_21 ) , .Z( u1_u7_X_32 ) );
  XOR2_X1 u1_u7_U25 (.B( u1_K8_31 ) , .A( u1_R6_20 ) , .Z( u1_u7_X_31 ) );
  XOR2_X1 u1_u7_U26 (.B( u1_K8_30 ) , .A( u1_R6_21 ) , .Z( u1_u7_X_30 ) );
  XOR2_X1 u1_u7_U27 (.B( u1_K8_2 ) , .A( u1_R6_1 ) , .Z( u1_u7_X_2 ) );
  XOR2_X1 u1_u7_U28 (.B( u1_K8_29 ) , .A( u1_R6_20 ) , .Z( u1_u7_X_29 ) );
  XOR2_X1 u1_u7_U29 (.B( u1_K8_28 ) , .A( u1_R6_19 ) , .Z( u1_u7_X_28 ) );
  XOR2_X1 u1_u7_U3 (.B( u1_K8_7 ) , .A( u1_R6_4 ) , .Z( u1_u7_X_7 ) );
  XOR2_X1 u1_u7_U30 (.B( u1_K8_27 ) , .A( u1_R6_18 ) , .Z( u1_u7_X_27 ) );
  XOR2_X1 u1_u7_U31 (.B( u1_K8_26 ) , .A( u1_R6_17 ) , .Z( u1_u7_X_26 ) );
  XOR2_X1 u1_u7_U32 (.B( u1_K8_25 ) , .A( u1_R6_16 ) , .Z( u1_u7_X_25 ) );
  XOR2_X1 u1_u7_U33 (.B( u1_K8_24 ) , .A( u1_R6_17 ) , .Z( u1_u7_X_24 ) );
  XOR2_X1 u1_u7_U34 (.B( u1_K8_23 ) , .A( u1_R6_16 ) , .Z( u1_u7_X_23 ) );
  XOR2_X1 u1_u7_U37 (.B( u1_K8_20 ) , .A( u1_R6_13 ) , .Z( u1_u7_X_20 ) );
  XOR2_X1 u1_u7_U38 (.B( u1_K8_1 ) , .A( u1_R6_32 ) , .Z( u1_u7_X_1 ) );
  XOR2_X1 u1_u7_U39 (.B( u1_K8_19 ) , .A( u1_R6_12 ) , .Z( u1_u7_X_19 ) );
  XOR2_X1 u1_u7_U4 (.B( u1_K8_6 ) , .A( u1_R6_5 ) , .Z( u1_u7_X_6 ) );
  XOR2_X1 u1_u7_U40 (.B( u1_K8_18 ) , .A( u1_R6_13 ) , .Z( u1_u7_X_18 ) );
  XOR2_X1 u1_u7_U41 (.B( u1_K8_17 ) , .A( u1_R6_12 ) , .Z( u1_u7_X_17 ) );
  XOR2_X1 u1_u7_U42 (.B( u1_K8_16 ) , .A( u1_R6_11 ) , .Z( u1_u7_X_16 ) );
  XOR2_X1 u1_u7_U43 (.B( u1_K8_15 ) , .A( u1_R6_10 ) , .Z( u1_u7_X_15 ) );
  XOR2_X1 u1_u7_U44 (.B( u1_K8_14 ) , .A( u1_R6_9 ) , .Z( u1_u7_X_14 ) );
  XOR2_X1 u1_u7_U45 (.B( u1_K8_13 ) , .A( u1_R6_8 ) , .Z( u1_u7_X_13 ) );
  XOR2_X1 u1_u7_U46 (.B( u1_K8_12 ) , .A( u1_R6_9 ) , .Z( u1_u7_X_12 ) );
  XOR2_X1 u1_u7_U47 (.B( u1_K8_11 ) , .A( u1_R6_8 ) , .Z( u1_u7_X_11 ) );
  XOR2_X1 u1_u7_U48 (.B( u1_K8_10 ) , .A( u1_R6_7 ) , .Z( u1_u7_X_10 ) );
  XOR2_X1 u1_u7_U5 (.B( u1_K8_5 ) , .A( u1_R6_4 ) , .Z( u1_u7_X_5 ) );
  XOR2_X1 u1_u7_U6 (.B( u1_K8_4 ) , .A( u1_R6_3 ) , .Z( u1_u7_X_4 ) );
  XOR2_X1 u1_u7_U7 (.B( u1_K8_48 ) , .A( u1_R6_1 ) , .Z( u1_u7_X_48 ) );
  XOR2_X1 u1_u7_U8 (.B( u1_K8_47 ) , .A( u1_R6_32 ) , .Z( u1_u7_X_47 ) );
  AND3_X1 u1_u7_u0_U10 (.A2( u1_u7_u0_n112 ) , .ZN( u1_u7_u0_n127 ) , .A3( u1_u7_u0_n130 ) , .A1( u1_u7_u0_n148 ) );
  NAND2_X1 u1_u7_u0_U11 (.ZN( u1_u7_u0_n113 ) , .A1( u1_u7_u0_n139 ) , .A2( u1_u7_u0_n149 ) );
  AND2_X1 u1_u7_u0_U12 (.ZN( u1_u7_u0_n107 ) , .A1( u1_u7_u0_n130 ) , .A2( u1_u7_u0_n140 ) );
  AND2_X1 u1_u7_u0_U13 (.A2( u1_u7_u0_n129 ) , .A1( u1_u7_u0_n130 ) , .ZN( u1_u7_u0_n151 ) );
  AND2_X1 u1_u7_u0_U14 (.A1( u1_u7_u0_n108 ) , .A2( u1_u7_u0_n125 ) , .ZN( u1_u7_u0_n145 ) );
  INV_X1 u1_u7_u0_U15 (.A( u1_u7_u0_n143 ) , .ZN( u1_u7_u0_n173 ) );
  NOR2_X1 u1_u7_u0_U16 (.A2( u1_u7_u0_n136 ) , .ZN( u1_u7_u0_n147 ) , .A1( u1_u7_u0_n160 ) );
  NOR2_X1 u1_u7_u0_U17 (.A1( u1_u7_u0_n163 ) , .A2( u1_u7_u0_n164 ) , .ZN( u1_u7_u0_n95 ) );
  AOI21_X1 u1_u7_u0_U18 (.B1( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n132 ) , .A( u1_u7_u0_n165 ) , .B2( u1_u7_u0_n93 ) );
  INV_X1 u1_u7_u0_U19 (.A( u1_u7_u0_n142 ) , .ZN( u1_u7_u0_n165 ) );
  OAI22_X1 u1_u7_u0_U20 (.B1( u1_u7_u0_n125 ) , .ZN( u1_u7_u0_n126 ) , .A1( u1_u7_u0_n138 ) , .A2( u1_u7_u0_n146 ) , .B2( u1_u7_u0_n147 ) );
  OAI22_X1 u1_u7_u0_U21 (.B1( u1_u7_u0_n131 ) , .A1( u1_u7_u0_n144 ) , .B2( u1_u7_u0_n147 ) , .A2( u1_u7_u0_n90 ) , .ZN( u1_u7_u0_n91 ) );
  AND3_X1 u1_u7_u0_U22 (.A3( u1_u7_u0_n121 ) , .A2( u1_u7_u0_n125 ) , .A1( u1_u7_u0_n148 ) , .ZN( u1_u7_u0_n90 ) );
  INV_X1 u1_u7_u0_U23 (.A( u1_u7_u0_n136 ) , .ZN( u1_u7_u0_n161 ) );
  AOI22_X1 u1_u7_u0_U24 (.B2( u1_u7_u0_n109 ) , .A2( u1_u7_u0_n110 ) , .ZN( u1_u7_u0_n111 ) , .B1( u1_u7_u0_n118 ) , .A1( u1_u7_u0_n160 ) );
  INV_X1 u1_u7_u0_U25 (.A( u1_u7_u0_n118 ) , .ZN( u1_u7_u0_n158 ) );
  AOI21_X1 u1_u7_u0_U26 (.ZN( u1_u7_u0_n104 ) , .B1( u1_u7_u0_n107 ) , .B2( u1_u7_u0_n141 ) , .A( u1_u7_u0_n144 ) );
  AOI21_X1 u1_u7_u0_U27 (.B1( u1_u7_u0_n127 ) , .B2( u1_u7_u0_n129 ) , .A( u1_u7_u0_n138 ) , .ZN( u1_u7_u0_n96 ) );
  AOI21_X1 u1_u7_u0_U28 (.ZN( u1_u7_u0_n116 ) , .B2( u1_u7_u0_n142 ) , .A( u1_u7_u0_n144 ) , .B1( u1_u7_u0_n166 ) );
  NOR2_X1 u1_u7_u0_U29 (.A1( u1_u7_u0_n120 ) , .ZN( u1_u7_u0_n143 ) , .A2( u1_u7_u0_n167 ) );
  INV_X1 u1_u7_u0_U3 (.A( u1_u7_u0_n113 ) , .ZN( u1_u7_u0_n166 ) );
  OAI221_X1 u1_u7_u0_U30 (.C1( u1_u7_u0_n112 ) , .ZN( u1_u7_u0_n120 ) , .B1( u1_u7_u0_n138 ) , .B2( u1_u7_u0_n141 ) , .C2( u1_u7_u0_n147 ) , .A( u1_u7_u0_n172 ) );
  AOI211_X1 u1_u7_u0_U31 (.B( u1_u7_u0_n115 ) , .A( u1_u7_u0_n116 ) , .C2( u1_u7_u0_n117 ) , .C1( u1_u7_u0_n118 ) , .ZN( u1_u7_u0_n119 ) );
  NAND2_X1 u1_u7_u0_U32 (.A1( u1_u7_u0_n100 ) , .A2( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n125 ) );
  NAND2_X1 u1_u7_u0_U33 (.A1( u1_u7_u0_n101 ) , .A2( u1_u7_u0_n102 ) , .ZN( u1_u7_u0_n150 ) );
  INV_X1 u1_u7_u0_U34 (.A( u1_u7_u0_n138 ) , .ZN( u1_u7_u0_n160 ) );
  NAND2_X1 u1_u7_u0_U35 (.A1( u1_u7_u0_n102 ) , .ZN( u1_u7_u0_n128 ) , .A2( u1_u7_u0_n95 ) );
  NAND2_X1 u1_u7_u0_U36 (.A1( u1_u7_u0_n100 ) , .ZN( u1_u7_u0_n129 ) , .A2( u1_u7_u0_n95 ) );
  NAND2_X1 u1_u7_u0_U37 (.A2( u1_u7_u0_n100 ) , .ZN( u1_u7_u0_n131 ) , .A1( u1_u7_u0_n92 ) );
  NAND2_X1 u1_u7_u0_U38 (.A2( u1_u7_u0_n100 ) , .A1( u1_u7_u0_n101 ) , .ZN( u1_u7_u0_n139 ) );
  NAND2_X1 u1_u7_u0_U39 (.ZN( u1_u7_u0_n148 ) , .A1( u1_u7_u0_n93 ) , .A2( u1_u7_u0_n95 ) );
  AOI21_X1 u1_u7_u0_U4 (.B1( u1_u7_u0_n114 ) , .ZN( u1_u7_u0_n115 ) , .B2( u1_u7_u0_n129 ) , .A( u1_u7_u0_n161 ) );
  NAND2_X1 u1_u7_u0_U40 (.A2( u1_u7_u0_n102 ) , .A1( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n149 ) );
  NAND2_X1 u1_u7_u0_U41 (.A2( u1_u7_u0_n102 ) , .ZN( u1_u7_u0_n114 ) , .A1( u1_u7_u0_n92 ) );
  NAND2_X1 u1_u7_u0_U42 (.A2( u1_u7_u0_n101 ) , .ZN( u1_u7_u0_n121 ) , .A1( u1_u7_u0_n93 ) );
  INV_X1 u1_u7_u0_U43 (.ZN( u1_u7_u0_n172 ) , .A( u1_u7_u0_n88 ) );
  OAI222_X1 u1_u7_u0_U44 (.C1( u1_u7_u0_n108 ) , .A1( u1_u7_u0_n125 ) , .B2( u1_u7_u0_n128 ) , .B1( u1_u7_u0_n144 ) , .A2( u1_u7_u0_n158 ) , .C2( u1_u7_u0_n161 ) , .ZN( u1_u7_u0_n88 ) );
  NAND2_X1 u1_u7_u0_U45 (.ZN( u1_u7_u0_n112 ) , .A2( u1_u7_u0_n92 ) , .A1( u1_u7_u0_n93 ) );
  OR3_X1 u1_u7_u0_U46 (.A3( u1_u7_u0_n152 ) , .A2( u1_u7_u0_n153 ) , .A1( u1_u7_u0_n154 ) , .ZN( u1_u7_u0_n155 ) );
  AOI21_X1 u1_u7_u0_U47 (.A( u1_u7_u0_n144 ) , .B2( u1_u7_u0_n145 ) , .B1( u1_u7_u0_n146 ) , .ZN( u1_u7_u0_n154 ) );
  AOI21_X1 u1_u7_u0_U48 (.B2( u1_u7_u0_n150 ) , .B1( u1_u7_u0_n151 ) , .ZN( u1_u7_u0_n152 ) , .A( u1_u7_u0_n158 ) );
  AOI21_X1 u1_u7_u0_U49 (.A( u1_u7_u0_n147 ) , .B2( u1_u7_u0_n148 ) , .B1( u1_u7_u0_n149 ) , .ZN( u1_u7_u0_n153 ) );
  AOI21_X1 u1_u7_u0_U5 (.B2( u1_u7_u0_n131 ) , .ZN( u1_u7_u0_n134 ) , .B1( u1_u7_u0_n151 ) , .A( u1_u7_u0_n158 ) );
  INV_X1 u1_u7_u0_U50 (.ZN( u1_u7_u0_n171 ) , .A( u1_u7_u0_n99 ) );
  OAI211_X1 u1_u7_u0_U51 (.C2( u1_u7_u0_n140 ) , .C1( u1_u7_u0_n161 ) , .A( u1_u7_u0_n169 ) , .B( u1_u7_u0_n98 ) , .ZN( u1_u7_u0_n99 ) );
  INV_X1 u1_u7_u0_U52 (.ZN( u1_u7_u0_n169 ) , .A( u1_u7_u0_n91 ) );
  AOI211_X1 u1_u7_u0_U53 (.C1( u1_u7_u0_n118 ) , .A( u1_u7_u0_n123 ) , .B( u1_u7_u0_n96 ) , .C2( u1_u7_u0_n97 ) , .ZN( u1_u7_u0_n98 ) );
  NOR2_X1 u1_u7_u0_U54 (.A2( u1_u7_X_6 ) , .ZN( u1_u7_u0_n100 ) , .A1( u1_u7_u0_n162 ) );
  NOR2_X1 u1_u7_u0_U55 (.A2( u1_u7_X_4 ) , .A1( u1_u7_X_5 ) , .ZN( u1_u7_u0_n118 ) );
  NOR2_X1 u1_u7_u0_U56 (.A2( u1_u7_X_2 ) , .ZN( u1_u7_u0_n103 ) , .A1( u1_u7_u0_n164 ) );
  NOR2_X1 u1_u7_u0_U57 (.A2( u1_u7_X_1 ) , .A1( u1_u7_X_2 ) , .ZN( u1_u7_u0_n92 ) );
  NOR2_X1 u1_u7_u0_U58 (.A2( u1_u7_X_1 ) , .ZN( u1_u7_u0_n101 ) , .A1( u1_u7_u0_n163 ) );
  NAND2_X1 u1_u7_u0_U59 (.A2( u1_u7_X_4 ) , .A1( u1_u7_X_5 ) , .ZN( u1_u7_u0_n144 ) );
  NOR2_X1 u1_u7_u0_U6 (.A1( u1_u7_u0_n108 ) , .ZN( u1_u7_u0_n123 ) , .A2( u1_u7_u0_n158 ) );
  NOR2_X1 u1_u7_u0_U60 (.A2( u1_u7_X_5 ) , .ZN( u1_u7_u0_n136 ) , .A1( u1_u7_u0_n159 ) );
  NAND2_X1 u1_u7_u0_U61 (.A1( u1_u7_X_5 ) , .ZN( u1_u7_u0_n138 ) , .A2( u1_u7_u0_n159 ) );
  NOR2_X1 u1_u7_u0_U62 (.A2( u1_u7_X_3 ) , .A1( u1_u7_X_6 ) , .ZN( u1_u7_u0_n94 ) );
  AND2_X1 u1_u7_u0_U63 (.A2( u1_u7_X_3 ) , .A1( u1_u7_X_6 ) , .ZN( u1_u7_u0_n102 ) );
  AND2_X1 u1_u7_u0_U64 (.A1( u1_u7_X_6 ) , .A2( u1_u7_u0_n162 ) , .ZN( u1_u7_u0_n93 ) );
  INV_X1 u1_u7_u0_U65 (.A( u1_u7_X_4 ) , .ZN( u1_u7_u0_n159 ) );
  INV_X1 u1_u7_u0_U66 (.A( u1_u7_X_1 ) , .ZN( u1_u7_u0_n164 ) );
  INV_X1 u1_u7_u0_U67 (.A( u1_u7_X_2 ) , .ZN( u1_u7_u0_n163 ) );
  INV_X1 u1_u7_u0_U68 (.A( u1_u7_X_3 ) , .ZN( u1_u7_u0_n162 ) );
  INV_X1 u1_u7_u0_U69 (.A( u1_u7_u0_n126 ) , .ZN( u1_u7_u0_n168 ) );
  OAI21_X1 u1_u7_u0_U7 (.B1( u1_u7_u0_n150 ) , .B2( u1_u7_u0_n158 ) , .A( u1_u7_u0_n172 ) , .ZN( u1_u7_u0_n89 ) );
  AOI211_X1 u1_u7_u0_U70 (.B( u1_u7_u0_n133 ) , .A( u1_u7_u0_n134 ) , .C2( u1_u7_u0_n135 ) , .C1( u1_u7_u0_n136 ) , .ZN( u1_u7_u0_n137 ) );
  OR4_X1 u1_u7_u0_U71 (.ZN( u1_out7_17 ) , .A1( u1_u7_u0_n122 ) , .A2( u1_u7_u0_n123 ) , .A4( u1_u7_u0_n124 ) , .A3( u1_u7_u0_n170 ) );
  AOI21_X1 u1_u7_u0_U72 (.B2( u1_u7_u0_n107 ) , .ZN( u1_u7_u0_n124 ) , .B1( u1_u7_u0_n128 ) , .A( u1_u7_u0_n161 ) );
  INV_X1 u1_u7_u0_U73 (.A( u1_u7_u0_n111 ) , .ZN( u1_u7_u0_n170 ) );
  OR4_X1 u1_u7_u0_U74 (.ZN( u1_out7_31 ) , .A4( u1_u7_u0_n155 ) , .A2( u1_u7_u0_n156 ) , .A1( u1_u7_u0_n157 ) , .A3( u1_u7_u0_n173 ) );
  AOI21_X1 u1_u7_u0_U75 (.A( u1_u7_u0_n138 ) , .B2( u1_u7_u0_n139 ) , .B1( u1_u7_u0_n140 ) , .ZN( u1_u7_u0_n157 ) );
  AOI21_X1 u1_u7_u0_U76 (.B2( u1_u7_u0_n141 ) , .B1( u1_u7_u0_n142 ) , .ZN( u1_u7_u0_n156 ) , .A( u1_u7_u0_n161 ) );
  INV_X1 u1_u7_u0_U77 (.ZN( u1_u7_u0_n174 ) , .A( u1_u7_u0_n89 ) );
  AOI211_X1 u1_u7_u0_U78 (.B( u1_u7_u0_n104 ) , .A( u1_u7_u0_n105 ) , .ZN( u1_u7_u0_n106 ) , .C2( u1_u7_u0_n113 ) , .C1( u1_u7_u0_n160 ) );
  OAI221_X1 u1_u7_u0_U79 (.C1( u1_u7_u0_n121 ) , .ZN( u1_u7_u0_n122 ) , .B2( u1_u7_u0_n127 ) , .A( u1_u7_u0_n143 ) , .B1( u1_u7_u0_n144 ) , .C2( u1_u7_u0_n147 ) );
  AND2_X1 u1_u7_u0_U8 (.A1( u1_u7_u0_n114 ) , .A2( u1_u7_u0_n121 ) , .ZN( u1_u7_u0_n146 ) );
  AOI21_X1 u1_u7_u0_U80 (.B1( u1_u7_u0_n132 ) , .ZN( u1_u7_u0_n133 ) , .A( u1_u7_u0_n144 ) , .B2( u1_u7_u0_n166 ) );
  OAI22_X1 u1_u7_u0_U81 (.ZN( u1_u7_u0_n105 ) , .A2( u1_u7_u0_n132 ) , .B1( u1_u7_u0_n146 ) , .A1( u1_u7_u0_n147 ) , .B2( u1_u7_u0_n161 ) );
  NAND2_X1 u1_u7_u0_U82 (.ZN( u1_u7_u0_n110 ) , .A2( u1_u7_u0_n132 ) , .A1( u1_u7_u0_n145 ) );
  INV_X1 u1_u7_u0_U83 (.A( u1_u7_u0_n119 ) , .ZN( u1_u7_u0_n167 ) );
  NAND2_X1 u1_u7_u0_U84 (.A2( u1_u7_u0_n103 ) , .ZN( u1_u7_u0_n140 ) , .A1( u1_u7_u0_n94 ) );
  NAND2_X1 u1_u7_u0_U85 (.A1( u1_u7_u0_n101 ) , .ZN( u1_u7_u0_n130 ) , .A2( u1_u7_u0_n94 ) );
  NAND2_X1 u1_u7_u0_U86 (.ZN( u1_u7_u0_n108 ) , .A1( u1_u7_u0_n92 ) , .A2( u1_u7_u0_n94 ) );
  NAND2_X1 u1_u7_u0_U87 (.ZN( u1_u7_u0_n142 ) , .A1( u1_u7_u0_n94 ) , .A2( u1_u7_u0_n95 ) );
  NAND3_X1 u1_u7_u0_U88 (.ZN( u1_out7_23 ) , .A3( u1_u7_u0_n137 ) , .A1( u1_u7_u0_n168 ) , .A2( u1_u7_u0_n171 ) );
  NAND3_X1 u1_u7_u0_U89 (.A3( u1_u7_u0_n127 ) , .A2( u1_u7_u0_n128 ) , .ZN( u1_u7_u0_n135 ) , .A1( u1_u7_u0_n150 ) );
  AND2_X1 u1_u7_u0_U9 (.A1( u1_u7_u0_n131 ) , .ZN( u1_u7_u0_n141 ) , .A2( u1_u7_u0_n150 ) );
  NAND3_X1 u1_u7_u0_U90 (.ZN( u1_u7_u0_n117 ) , .A3( u1_u7_u0_n132 ) , .A2( u1_u7_u0_n139 ) , .A1( u1_u7_u0_n148 ) );
  NAND3_X1 u1_u7_u0_U91 (.ZN( u1_u7_u0_n109 ) , .A2( u1_u7_u0_n114 ) , .A3( u1_u7_u0_n140 ) , .A1( u1_u7_u0_n149 ) );
  NAND3_X1 u1_u7_u0_U92 (.ZN( u1_out7_9 ) , .A3( u1_u7_u0_n106 ) , .A2( u1_u7_u0_n171 ) , .A1( u1_u7_u0_n174 ) );
  NAND3_X1 u1_u7_u0_U93 (.A2( u1_u7_u0_n128 ) , .A1( u1_u7_u0_n132 ) , .A3( u1_u7_u0_n146 ) , .ZN( u1_u7_u0_n97 ) );
  AOI21_X1 u1_u7_u1_U10 (.B2( u1_u7_u1_n155 ) , .B1( u1_u7_u1_n156 ) , .ZN( u1_u7_u1_n157 ) , .A( u1_u7_u1_n174 ) );
  NAND3_X1 u1_u7_u1_U100 (.ZN( u1_u7_u1_n113 ) , .A1( u1_u7_u1_n120 ) , .A3( u1_u7_u1_n133 ) , .A2( u1_u7_u1_n155 ) );
  NAND2_X1 u1_u7_u1_U11 (.ZN( u1_u7_u1_n140 ) , .A2( u1_u7_u1_n150 ) , .A1( u1_u7_u1_n155 ) );
  NAND2_X1 u1_u7_u1_U12 (.A1( u1_u7_u1_n131 ) , .ZN( u1_u7_u1_n147 ) , .A2( u1_u7_u1_n153 ) );
  AOI22_X1 u1_u7_u1_U13 (.B2( u1_u7_u1_n136 ) , .A2( u1_u7_u1_n137 ) , .ZN( u1_u7_u1_n143 ) , .A1( u1_u7_u1_n171 ) , .B1( u1_u7_u1_n173 ) );
  INV_X1 u1_u7_u1_U14 (.A( u1_u7_u1_n147 ) , .ZN( u1_u7_u1_n181 ) );
  INV_X1 u1_u7_u1_U15 (.A( u1_u7_u1_n139 ) , .ZN( u1_u7_u1_n174 ) );
  OR4_X1 u1_u7_u1_U16 (.A4( u1_u7_u1_n106 ) , .A3( u1_u7_u1_n107 ) , .ZN( u1_u7_u1_n108 ) , .A1( u1_u7_u1_n117 ) , .A2( u1_u7_u1_n184 ) );
  AOI21_X1 u1_u7_u1_U17 (.ZN( u1_u7_u1_n106 ) , .A( u1_u7_u1_n112 ) , .B1( u1_u7_u1_n154 ) , .B2( u1_u7_u1_n156 ) );
  AOI21_X1 u1_u7_u1_U18 (.ZN( u1_u7_u1_n107 ) , .B1( u1_u7_u1_n134 ) , .B2( u1_u7_u1_n149 ) , .A( u1_u7_u1_n174 ) );
  INV_X1 u1_u7_u1_U19 (.A( u1_u7_u1_n101 ) , .ZN( u1_u7_u1_n184 ) );
  INV_X1 u1_u7_u1_U20 (.A( u1_u7_u1_n112 ) , .ZN( u1_u7_u1_n171 ) );
  NAND2_X1 u1_u7_u1_U21 (.ZN( u1_u7_u1_n141 ) , .A1( u1_u7_u1_n153 ) , .A2( u1_u7_u1_n156 ) );
  AND2_X1 u1_u7_u1_U22 (.A1( u1_u7_u1_n123 ) , .ZN( u1_u7_u1_n134 ) , .A2( u1_u7_u1_n161 ) );
  NAND2_X1 u1_u7_u1_U23 (.A2( u1_u7_u1_n115 ) , .A1( u1_u7_u1_n116 ) , .ZN( u1_u7_u1_n148 ) );
  NAND2_X1 u1_u7_u1_U24 (.A2( u1_u7_u1_n133 ) , .A1( u1_u7_u1_n135 ) , .ZN( u1_u7_u1_n159 ) );
  NAND2_X1 u1_u7_u1_U25 (.A2( u1_u7_u1_n115 ) , .A1( u1_u7_u1_n120 ) , .ZN( u1_u7_u1_n132 ) );
  INV_X1 u1_u7_u1_U26 (.A( u1_u7_u1_n154 ) , .ZN( u1_u7_u1_n178 ) );
  INV_X1 u1_u7_u1_U27 (.A( u1_u7_u1_n151 ) , .ZN( u1_u7_u1_n183 ) );
  AND2_X1 u1_u7_u1_U28 (.A1( u1_u7_u1_n129 ) , .A2( u1_u7_u1_n133 ) , .ZN( u1_u7_u1_n149 ) );
  INV_X1 u1_u7_u1_U29 (.A( u1_u7_u1_n131 ) , .ZN( u1_u7_u1_n180 ) );
  INV_X1 u1_u7_u1_U3 (.A( u1_u7_u1_n159 ) , .ZN( u1_u7_u1_n182 ) );
  OAI221_X1 u1_u7_u1_U30 (.A( u1_u7_u1_n119 ) , .C2( u1_u7_u1_n129 ) , .ZN( u1_u7_u1_n138 ) , .B2( u1_u7_u1_n152 ) , .C1( u1_u7_u1_n174 ) , .B1( u1_u7_u1_n187 ) );
  INV_X1 u1_u7_u1_U31 (.A( u1_u7_u1_n148 ) , .ZN( u1_u7_u1_n187 ) );
  AOI211_X1 u1_u7_u1_U32 (.B( u1_u7_u1_n117 ) , .A( u1_u7_u1_n118 ) , .ZN( u1_u7_u1_n119 ) , .C2( u1_u7_u1_n146 ) , .C1( u1_u7_u1_n159 ) );
  NOR2_X1 u1_u7_u1_U33 (.A1( u1_u7_u1_n168 ) , .A2( u1_u7_u1_n176 ) , .ZN( u1_u7_u1_n98 ) );
  AOI211_X1 u1_u7_u1_U34 (.B( u1_u7_u1_n162 ) , .A( u1_u7_u1_n163 ) , .C2( u1_u7_u1_n164 ) , .ZN( u1_u7_u1_n165 ) , .C1( u1_u7_u1_n171 ) );
  AOI21_X1 u1_u7_u1_U35 (.A( u1_u7_u1_n160 ) , .B2( u1_u7_u1_n161 ) , .ZN( u1_u7_u1_n162 ) , .B1( u1_u7_u1_n182 ) );
  OR2_X1 u1_u7_u1_U36 (.A2( u1_u7_u1_n157 ) , .A1( u1_u7_u1_n158 ) , .ZN( u1_u7_u1_n163 ) );
  NAND2_X1 u1_u7_u1_U37 (.A1( u1_u7_u1_n128 ) , .ZN( u1_u7_u1_n146 ) , .A2( u1_u7_u1_n160 ) );
  NAND2_X1 u1_u7_u1_U38 (.A2( u1_u7_u1_n112 ) , .ZN( u1_u7_u1_n139 ) , .A1( u1_u7_u1_n152 ) );
  NAND2_X1 u1_u7_u1_U39 (.A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n156 ) , .A2( u1_u7_u1_n99 ) );
  AOI221_X1 u1_u7_u1_U4 (.A( u1_u7_u1_n138 ) , .C2( u1_u7_u1_n139 ) , .C1( u1_u7_u1_n140 ) , .B2( u1_u7_u1_n141 ) , .ZN( u1_u7_u1_n142 ) , .B1( u1_u7_u1_n175 ) );
  AOI221_X1 u1_u7_u1_U40 (.B1( u1_u7_u1_n140 ) , .ZN( u1_u7_u1_n167 ) , .B2( u1_u7_u1_n172 ) , .C2( u1_u7_u1_n175 ) , .C1( u1_u7_u1_n178 ) , .A( u1_u7_u1_n188 ) );
  INV_X1 u1_u7_u1_U41 (.ZN( u1_u7_u1_n188 ) , .A( u1_u7_u1_n97 ) );
  AOI211_X1 u1_u7_u1_U42 (.A( u1_u7_u1_n118 ) , .C1( u1_u7_u1_n132 ) , .C2( u1_u7_u1_n139 ) , .B( u1_u7_u1_n96 ) , .ZN( u1_u7_u1_n97 ) );
  AOI21_X1 u1_u7_u1_U43 (.B2( u1_u7_u1_n121 ) , .B1( u1_u7_u1_n135 ) , .A( u1_u7_u1_n152 ) , .ZN( u1_u7_u1_n96 ) );
  NOR2_X1 u1_u7_u1_U44 (.ZN( u1_u7_u1_n117 ) , .A1( u1_u7_u1_n121 ) , .A2( u1_u7_u1_n160 ) );
  OAI21_X1 u1_u7_u1_U45 (.B2( u1_u7_u1_n123 ) , .ZN( u1_u7_u1_n145 ) , .B1( u1_u7_u1_n160 ) , .A( u1_u7_u1_n185 ) );
  INV_X1 u1_u7_u1_U46 (.A( u1_u7_u1_n122 ) , .ZN( u1_u7_u1_n185 ) );
  AOI21_X1 u1_u7_u1_U47 (.B2( u1_u7_u1_n120 ) , .B1( u1_u7_u1_n121 ) , .ZN( u1_u7_u1_n122 ) , .A( u1_u7_u1_n128 ) );
  AOI21_X1 u1_u7_u1_U48 (.A( u1_u7_u1_n128 ) , .B2( u1_u7_u1_n129 ) , .ZN( u1_u7_u1_n130 ) , .B1( u1_u7_u1_n150 ) );
  NAND2_X1 u1_u7_u1_U49 (.ZN( u1_u7_u1_n112 ) , .A1( u1_u7_u1_n169 ) , .A2( u1_u7_u1_n170 ) );
  AOI211_X1 u1_u7_u1_U5 (.ZN( u1_u7_u1_n124 ) , .A( u1_u7_u1_n138 ) , .C2( u1_u7_u1_n139 ) , .B( u1_u7_u1_n145 ) , .C1( u1_u7_u1_n147 ) );
  NAND2_X1 u1_u7_u1_U50 (.ZN( u1_u7_u1_n129 ) , .A2( u1_u7_u1_n95 ) , .A1( u1_u7_u1_n98 ) );
  NAND2_X1 u1_u7_u1_U51 (.A1( u1_u7_u1_n102 ) , .ZN( u1_u7_u1_n154 ) , .A2( u1_u7_u1_n99 ) );
  NAND2_X1 u1_u7_u1_U52 (.A2( u1_u7_u1_n100 ) , .ZN( u1_u7_u1_n135 ) , .A1( u1_u7_u1_n99 ) );
  AOI21_X1 u1_u7_u1_U53 (.A( u1_u7_u1_n152 ) , .B2( u1_u7_u1_n153 ) , .B1( u1_u7_u1_n154 ) , .ZN( u1_u7_u1_n158 ) );
  INV_X1 u1_u7_u1_U54 (.A( u1_u7_u1_n160 ) , .ZN( u1_u7_u1_n175 ) );
  NAND2_X1 u1_u7_u1_U55 (.A1( u1_u7_u1_n100 ) , .ZN( u1_u7_u1_n116 ) , .A2( u1_u7_u1_n95 ) );
  NAND2_X1 u1_u7_u1_U56 (.A1( u1_u7_u1_n102 ) , .ZN( u1_u7_u1_n131 ) , .A2( u1_u7_u1_n95 ) );
  NAND2_X1 u1_u7_u1_U57 (.A2( u1_u7_u1_n104 ) , .ZN( u1_u7_u1_n121 ) , .A1( u1_u7_u1_n98 ) );
  NAND2_X1 u1_u7_u1_U58 (.A1( u1_u7_u1_n103 ) , .ZN( u1_u7_u1_n153 ) , .A2( u1_u7_u1_n98 ) );
  NAND2_X1 u1_u7_u1_U59 (.A2( u1_u7_u1_n104 ) , .A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n133 ) );
  AOI22_X1 u1_u7_u1_U6 (.B2( u1_u7_u1_n113 ) , .A2( u1_u7_u1_n114 ) , .ZN( u1_u7_u1_n125 ) , .A1( u1_u7_u1_n171 ) , .B1( u1_u7_u1_n173 ) );
  NAND2_X1 u1_u7_u1_U60 (.ZN( u1_u7_u1_n150 ) , .A2( u1_u7_u1_n98 ) , .A1( u1_u7_u1_n99 ) );
  NAND2_X1 u1_u7_u1_U61 (.A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n155 ) , .A2( u1_u7_u1_n95 ) );
  OAI21_X1 u1_u7_u1_U62 (.ZN( u1_u7_u1_n109 ) , .B1( u1_u7_u1_n129 ) , .B2( u1_u7_u1_n160 ) , .A( u1_u7_u1_n167 ) );
  NAND2_X1 u1_u7_u1_U63 (.A2( u1_u7_u1_n100 ) , .A1( u1_u7_u1_n103 ) , .ZN( u1_u7_u1_n120 ) );
  NAND2_X1 u1_u7_u1_U64 (.A1( u1_u7_u1_n102 ) , .A2( u1_u7_u1_n104 ) , .ZN( u1_u7_u1_n115 ) );
  NAND2_X1 u1_u7_u1_U65 (.A2( u1_u7_u1_n100 ) , .A1( u1_u7_u1_n104 ) , .ZN( u1_u7_u1_n151 ) );
  NAND2_X1 u1_u7_u1_U66 (.A2( u1_u7_u1_n103 ) , .A1( u1_u7_u1_n105 ) , .ZN( u1_u7_u1_n161 ) );
  INV_X1 u1_u7_u1_U67 (.A( u1_u7_u1_n152 ) , .ZN( u1_u7_u1_n173 ) );
  INV_X1 u1_u7_u1_U68 (.A( u1_u7_u1_n128 ) , .ZN( u1_u7_u1_n172 ) );
  NAND2_X1 u1_u7_u1_U69 (.A2( u1_u7_u1_n102 ) , .A1( u1_u7_u1_n103 ) , .ZN( u1_u7_u1_n123 ) );
  NAND2_X1 u1_u7_u1_U7 (.ZN( u1_u7_u1_n114 ) , .A1( u1_u7_u1_n134 ) , .A2( u1_u7_u1_n156 ) );
  NOR2_X1 u1_u7_u1_U70 (.A2( u1_u7_X_7 ) , .A1( u1_u7_X_8 ) , .ZN( u1_u7_u1_n95 ) );
  NOR2_X1 u1_u7_u1_U71 (.A1( u1_u7_X_12 ) , .A2( u1_u7_X_9 ) , .ZN( u1_u7_u1_n100 ) );
  NOR2_X1 u1_u7_u1_U72 (.A2( u1_u7_X_8 ) , .A1( u1_u7_u1_n177 ) , .ZN( u1_u7_u1_n99 ) );
  NOR2_X1 u1_u7_u1_U73 (.A2( u1_u7_X_12 ) , .ZN( u1_u7_u1_n102 ) , .A1( u1_u7_u1_n176 ) );
  NOR2_X1 u1_u7_u1_U74 (.A2( u1_u7_X_9 ) , .ZN( u1_u7_u1_n105 ) , .A1( u1_u7_u1_n168 ) );
  NAND2_X1 u1_u7_u1_U75 (.A1( u1_u7_X_10 ) , .ZN( u1_u7_u1_n160 ) , .A2( u1_u7_u1_n169 ) );
  NAND2_X1 u1_u7_u1_U76 (.A2( u1_u7_X_10 ) , .A1( u1_u7_X_11 ) , .ZN( u1_u7_u1_n152 ) );
  NAND2_X1 u1_u7_u1_U77 (.A1( u1_u7_X_11 ) , .ZN( u1_u7_u1_n128 ) , .A2( u1_u7_u1_n170 ) );
  AND2_X1 u1_u7_u1_U78 (.A2( u1_u7_X_7 ) , .A1( u1_u7_X_8 ) , .ZN( u1_u7_u1_n104 ) );
  AND2_X1 u1_u7_u1_U79 (.A1( u1_u7_X_8 ) , .ZN( u1_u7_u1_n103 ) , .A2( u1_u7_u1_n177 ) );
  NOR2_X1 u1_u7_u1_U8 (.A1( u1_u7_u1_n112 ) , .A2( u1_u7_u1_n116 ) , .ZN( u1_u7_u1_n118 ) );
  INV_X1 u1_u7_u1_U80 (.A( u1_u7_X_10 ) , .ZN( u1_u7_u1_n170 ) );
  INV_X1 u1_u7_u1_U81 (.A( u1_u7_X_9 ) , .ZN( u1_u7_u1_n176 ) );
  INV_X1 u1_u7_u1_U82 (.A( u1_u7_X_11 ) , .ZN( u1_u7_u1_n169 ) );
  INV_X1 u1_u7_u1_U83 (.A( u1_u7_X_12 ) , .ZN( u1_u7_u1_n168 ) );
  INV_X1 u1_u7_u1_U84 (.A( u1_u7_X_7 ) , .ZN( u1_u7_u1_n177 ) );
  NAND4_X1 u1_u7_u1_U85 (.ZN( u1_out7_18 ) , .A4( u1_u7_u1_n165 ) , .A3( u1_u7_u1_n166 ) , .A1( u1_u7_u1_n167 ) , .A2( u1_u7_u1_n186 ) );
  AOI22_X1 u1_u7_u1_U86 (.B2( u1_u7_u1_n146 ) , .B1( u1_u7_u1_n147 ) , .A2( u1_u7_u1_n148 ) , .ZN( u1_u7_u1_n166 ) , .A1( u1_u7_u1_n172 ) );
  INV_X1 u1_u7_u1_U87 (.A( u1_u7_u1_n145 ) , .ZN( u1_u7_u1_n186 ) );
  NAND4_X1 u1_u7_u1_U88 (.ZN( u1_out7_2 ) , .A4( u1_u7_u1_n142 ) , .A3( u1_u7_u1_n143 ) , .A2( u1_u7_u1_n144 ) , .A1( u1_u7_u1_n179 ) );
  OAI21_X1 u1_u7_u1_U89 (.B2( u1_u7_u1_n132 ) , .ZN( u1_u7_u1_n144 ) , .A( u1_u7_u1_n146 ) , .B1( u1_u7_u1_n180 ) );
  OAI21_X1 u1_u7_u1_U9 (.ZN( u1_u7_u1_n101 ) , .B1( u1_u7_u1_n141 ) , .A( u1_u7_u1_n146 ) , .B2( u1_u7_u1_n183 ) );
  INV_X1 u1_u7_u1_U90 (.A( u1_u7_u1_n130 ) , .ZN( u1_u7_u1_n179 ) );
  NAND4_X1 u1_u7_u1_U91 (.ZN( u1_out7_28 ) , .A4( u1_u7_u1_n124 ) , .A3( u1_u7_u1_n125 ) , .A2( u1_u7_u1_n126 ) , .A1( u1_u7_u1_n127 ) );
  OAI21_X1 u1_u7_u1_U92 (.ZN( u1_u7_u1_n127 ) , .B2( u1_u7_u1_n139 ) , .B1( u1_u7_u1_n175 ) , .A( u1_u7_u1_n183 ) );
  OAI21_X1 u1_u7_u1_U93 (.ZN( u1_u7_u1_n126 ) , .B2( u1_u7_u1_n140 ) , .A( u1_u7_u1_n146 ) , .B1( u1_u7_u1_n178 ) );
  OR4_X1 u1_u7_u1_U94 (.ZN( u1_out7_13 ) , .A4( u1_u7_u1_n108 ) , .A3( u1_u7_u1_n109 ) , .A2( u1_u7_u1_n110 ) , .A1( u1_u7_u1_n111 ) );
  AOI21_X1 u1_u7_u1_U95 (.ZN( u1_u7_u1_n111 ) , .A( u1_u7_u1_n128 ) , .B2( u1_u7_u1_n131 ) , .B1( u1_u7_u1_n135 ) );
  AOI21_X1 u1_u7_u1_U96 (.ZN( u1_u7_u1_n110 ) , .A( u1_u7_u1_n116 ) , .B1( u1_u7_u1_n152 ) , .B2( u1_u7_u1_n160 ) );
  NAND3_X1 u1_u7_u1_U97 (.A3( u1_u7_u1_n149 ) , .A2( u1_u7_u1_n150 ) , .A1( u1_u7_u1_n151 ) , .ZN( u1_u7_u1_n164 ) );
  NAND3_X1 u1_u7_u1_U98 (.A3( u1_u7_u1_n134 ) , .A2( u1_u7_u1_n135 ) , .ZN( u1_u7_u1_n136 ) , .A1( u1_u7_u1_n151 ) );
  NAND3_X1 u1_u7_u1_U99 (.A1( u1_u7_u1_n133 ) , .ZN( u1_u7_u1_n137 ) , .A2( u1_u7_u1_n154 ) , .A3( u1_u7_u1_n181 ) );
  OAI22_X1 u1_u7_u2_U10 (.ZN( u1_u7_u2_n109 ) , .A2( u1_u7_u2_n113 ) , .B2( u1_u7_u2_n133 ) , .B1( u1_u7_u2_n167 ) , .A1( u1_u7_u2_n168 ) );
  NAND3_X1 u1_u7_u2_U100 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n104 ) , .A3( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n98 ) );
  OAI22_X1 u1_u7_u2_U11 (.B1( u1_u7_u2_n151 ) , .A2( u1_u7_u2_n152 ) , .A1( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n160 ) , .B2( u1_u7_u2_n168 ) );
  NOR3_X1 u1_u7_u2_U12 (.A1( u1_u7_u2_n150 ) , .ZN( u1_u7_u2_n151 ) , .A3( u1_u7_u2_n175 ) , .A2( u1_u7_u2_n188 ) );
  AOI21_X1 u1_u7_u2_U13 (.ZN( u1_u7_u2_n144 ) , .B2( u1_u7_u2_n155 ) , .A( u1_u7_u2_n172 ) , .B1( u1_u7_u2_n185 ) );
  AOI21_X1 u1_u7_u2_U14 (.B2( u1_u7_u2_n143 ) , .ZN( u1_u7_u2_n145 ) , .B1( u1_u7_u2_n152 ) , .A( u1_u7_u2_n171 ) );
  AOI21_X1 u1_u7_u2_U15 (.B2( u1_u7_u2_n120 ) , .B1( u1_u7_u2_n121 ) , .ZN( u1_u7_u2_n126 ) , .A( u1_u7_u2_n167 ) );
  INV_X1 u1_u7_u2_U16 (.A( u1_u7_u2_n156 ) , .ZN( u1_u7_u2_n171 ) );
  INV_X1 u1_u7_u2_U17 (.A( u1_u7_u2_n120 ) , .ZN( u1_u7_u2_n188 ) );
  NAND2_X1 u1_u7_u2_U18 (.A2( u1_u7_u2_n122 ) , .ZN( u1_u7_u2_n150 ) , .A1( u1_u7_u2_n152 ) );
  INV_X1 u1_u7_u2_U19 (.A( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n170 ) );
  INV_X1 u1_u7_u2_U20 (.A( u1_u7_u2_n137 ) , .ZN( u1_u7_u2_n173 ) );
  NAND2_X1 u1_u7_u2_U21 (.A1( u1_u7_u2_n132 ) , .A2( u1_u7_u2_n139 ) , .ZN( u1_u7_u2_n157 ) );
  INV_X1 u1_u7_u2_U22 (.A( u1_u7_u2_n113 ) , .ZN( u1_u7_u2_n178 ) );
  INV_X1 u1_u7_u2_U23 (.A( u1_u7_u2_n139 ) , .ZN( u1_u7_u2_n175 ) );
  INV_X1 u1_u7_u2_U24 (.A( u1_u7_u2_n155 ) , .ZN( u1_u7_u2_n181 ) );
  INV_X1 u1_u7_u2_U25 (.A( u1_u7_u2_n119 ) , .ZN( u1_u7_u2_n177 ) );
  INV_X1 u1_u7_u2_U26 (.A( u1_u7_u2_n116 ) , .ZN( u1_u7_u2_n180 ) );
  INV_X1 u1_u7_u2_U27 (.A( u1_u7_u2_n131 ) , .ZN( u1_u7_u2_n179 ) );
  INV_X1 u1_u7_u2_U28 (.A( u1_u7_u2_n154 ) , .ZN( u1_u7_u2_n176 ) );
  NAND2_X1 u1_u7_u2_U29 (.A2( u1_u7_u2_n116 ) , .A1( u1_u7_u2_n117 ) , .ZN( u1_u7_u2_n118 ) );
  NOR2_X1 u1_u7_u2_U3 (.ZN( u1_u7_u2_n121 ) , .A2( u1_u7_u2_n177 ) , .A1( u1_u7_u2_n180 ) );
  INV_X1 u1_u7_u2_U30 (.A( u1_u7_u2_n132 ) , .ZN( u1_u7_u2_n182 ) );
  INV_X1 u1_u7_u2_U31 (.A( u1_u7_u2_n158 ) , .ZN( u1_u7_u2_n183 ) );
  OAI21_X1 u1_u7_u2_U32 (.A( u1_u7_u2_n156 ) , .B1( u1_u7_u2_n157 ) , .ZN( u1_u7_u2_n158 ) , .B2( u1_u7_u2_n179 ) );
  NOR2_X1 u1_u7_u2_U33 (.ZN( u1_u7_u2_n156 ) , .A1( u1_u7_u2_n166 ) , .A2( u1_u7_u2_n169 ) );
  NOR2_X1 u1_u7_u2_U34 (.A2( u1_u7_u2_n114 ) , .ZN( u1_u7_u2_n137 ) , .A1( u1_u7_u2_n140 ) );
  NOR2_X1 u1_u7_u2_U35 (.A2( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n153 ) , .A1( u1_u7_u2_n156 ) );
  AOI211_X1 u1_u7_u2_U36 (.ZN( u1_u7_u2_n130 ) , .C1( u1_u7_u2_n138 ) , .C2( u1_u7_u2_n179 ) , .B( u1_u7_u2_n96 ) , .A( u1_u7_u2_n97 ) );
  OAI22_X1 u1_u7_u2_U37 (.B1( u1_u7_u2_n133 ) , .A2( u1_u7_u2_n137 ) , .A1( u1_u7_u2_n152 ) , .B2( u1_u7_u2_n168 ) , .ZN( u1_u7_u2_n97 ) );
  OAI221_X1 u1_u7_u2_U38 (.B1( u1_u7_u2_n113 ) , .C1( u1_u7_u2_n132 ) , .A( u1_u7_u2_n149 ) , .B2( u1_u7_u2_n171 ) , .C2( u1_u7_u2_n172 ) , .ZN( u1_u7_u2_n96 ) );
  OAI221_X1 u1_u7_u2_U39 (.A( u1_u7_u2_n115 ) , .C2( u1_u7_u2_n123 ) , .B2( u1_u7_u2_n143 ) , .B1( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n163 ) , .C1( u1_u7_u2_n168 ) );
  INV_X1 u1_u7_u2_U4 (.A( u1_u7_u2_n134 ) , .ZN( u1_u7_u2_n185 ) );
  OAI21_X1 u1_u7_u2_U40 (.A( u1_u7_u2_n114 ) , .ZN( u1_u7_u2_n115 ) , .B1( u1_u7_u2_n176 ) , .B2( u1_u7_u2_n178 ) );
  OAI221_X1 u1_u7_u2_U41 (.A( u1_u7_u2_n135 ) , .B2( u1_u7_u2_n136 ) , .B1( u1_u7_u2_n137 ) , .ZN( u1_u7_u2_n162 ) , .C2( u1_u7_u2_n167 ) , .C1( u1_u7_u2_n185 ) );
  AND3_X1 u1_u7_u2_U42 (.A3( u1_u7_u2_n131 ) , .A2( u1_u7_u2_n132 ) , .A1( u1_u7_u2_n133 ) , .ZN( u1_u7_u2_n136 ) );
  AOI22_X1 u1_u7_u2_U43 (.ZN( u1_u7_u2_n135 ) , .B1( u1_u7_u2_n140 ) , .A1( u1_u7_u2_n156 ) , .B2( u1_u7_u2_n180 ) , .A2( u1_u7_u2_n188 ) );
  AOI21_X1 u1_u7_u2_U44 (.ZN( u1_u7_u2_n149 ) , .B1( u1_u7_u2_n173 ) , .B2( u1_u7_u2_n188 ) , .A( u1_u7_u2_n95 ) );
  AND3_X1 u1_u7_u2_U45 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n104 ) , .A3( u1_u7_u2_n156 ) , .ZN( u1_u7_u2_n95 ) );
  OAI21_X1 u1_u7_u2_U46 (.A( u1_u7_u2_n101 ) , .B2( u1_u7_u2_n121 ) , .B1( u1_u7_u2_n153 ) , .ZN( u1_u7_u2_n164 ) );
  NAND2_X1 u1_u7_u2_U47 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n107 ) , .ZN( u1_u7_u2_n155 ) );
  NAND2_X1 u1_u7_u2_U48 (.A2( u1_u7_u2_n105 ) , .A1( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n143 ) );
  NAND2_X1 u1_u7_u2_U49 (.A1( u1_u7_u2_n104 ) , .A2( u1_u7_u2_n106 ) , .ZN( u1_u7_u2_n152 ) );
  INV_X1 u1_u7_u2_U5 (.A( u1_u7_u2_n150 ) , .ZN( u1_u7_u2_n184 ) );
  NAND2_X1 u1_u7_u2_U50 (.A1( u1_u7_u2_n100 ) , .A2( u1_u7_u2_n105 ) , .ZN( u1_u7_u2_n132 ) );
  INV_X1 u1_u7_u2_U51 (.A( u1_u7_u2_n140 ) , .ZN( u1_u7_u2_n168 ) );
  INV_X1 u1_u7_u2_U52 (.A( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n167 ) );
  OAI21_X1 u1_u7_u2_U53 (.A( u1_u7_u2_n141 ) , .B2( u1_u7_u2_n142 ) , .ZN( u1_u7_u2_n146 ) , .B1( u1_u7_u2_n153 ) );
  OAI21_X1 u1_u7_u2_U54 (.A( u1_u7_u2_n140 ) , .ZN( u1_u7_u2_n141 ) , .B1( u1_u7_u2_n176 ) , .B2( u1_u7_u2_n177 ) );
  NOR3_X1 u1_u7_u2_U55 (.ZN( u1_u7_u2_n142 ) , .A3( u1_u7_u2_n175 ) , .A2( u1_u7_u2_n178 ) , .A1( u1_u7_u2_n181 ) );
  INV_X1 u1_u7_u2_U56 (.ZN( u1_u7_u2_n187 ) , .A( u1_u7_u2_n99 ) );
  OAI21_X1 u1_u7_u2_U57 (.B1( u1_u7_u2_n137 ) , .B2( u1_u7_u2_n143 ) , .A( u1_u7_u2_n98 ) , .ZN( u1_u7_u2_n99 ) );
  NAND2_X1 u1_u7_u2_U58 (.A1( u1_u7_u2_n102 ) , .A2( u1_u7_u2_n106 ) , .ZN( u1_u7_u2_n113 ) );
  NAND2_X1 u1_u7_u2_U59 (.A1( u1_u7_u2_n106 ) , .A2( u1_u7_u2_n107 ) , .ZN( u1_u7_u2_n131 ) );
  NOR4_X1 u1_u7_u2_U6 (.A4( u1_u7_u2_n124 ) , .A3( u1_u7_u2_n125 ) , .A2( u1_u7_u2_n126 ) , .A1( u1_u7_u2_n127 ) , .ZN( u1_u7_u2_n128 ) );
  NAND2_X1 u1_u7_u2_U60 (.A1( u1_u7_u2_n103 ) , .A2( u1_u7_u2_n107 ) , .ZN( u1_u7_u2_n139 ) );
  NAND2_X1 u1_u7_u2_U61 (.A1( u1_u7_u2_n103 ) , .A2( u1_u7_u2_n105 ) , .ZN( u1_u7_u2_n133 ) );
  NAND2_X1 u1_u7_u2_U62 (.A1( u1_u7_u2_n102 ) , .A2( u1_u7_u2_n103 ) , .ZN( u1_u7_u2_n154 ) );
  NAND2_X1 u1_u7_u2_U63 (.A2( u1_u7_u2_n103 ) , .A1( u1_u7_u2_n104 ) , .ZN( u1_u7_u2_n119 ) );
  NAND2_X1 u1_u7_u2_U64 (.A2( u1_u7_u2_n107 ) , .A1( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n123 ) );
  NAND2_X1 u1_u7_u2_U65 (.A1( u1_u7_u2_n104 ) , .A2( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n122 ) );
  INV_X1 u1_u7_u2_U66 (.A( u1_u7_u2_n114 ) , .ZN( u1_u7_u2_n172 ) );
  NAND2_X1 u1_u7_u2_U67 (.A2( u1_u7_u2_n100 ) , .A1( u1_u7_u2_n102 ) , .ZN( u1_u7_u2_n116 ) );
  NAND2_X1 u1_u7_u2_U68 (.A1( u1_u7_u2_n102 ) , .A2( u1_u7_u2_n108 ) , .ZN( u1_u7_u2_n120 ) );
  NAND2_X1 u1_u7_u2_U69 (.A2( u1_u7_u2_n105 ) , .A1( u1_u7_u2_n106 ) , .ZN( u1_u7_u2_n117 ) );
  AOI21_X1 u1_u7_u2_U7 (.B2( u1_u7_u2_n119 ) , .ZN( u1_u7_u2_n127 ) , .A( u1_u7_u2_n137 ) , .B1( u1_u7_u2_n155 ) );
  NOR2_X1 u1_u7_u2_U70 (.A2( u1_u7_X_16 ) , .ZN( u1_u7_u2_n140 ) , .A1( u1_u7_u2_n166 ) );
  NOR2_X1 u1_u7_u2_U71 (.A2( u1_u7_X_13 ) , .A1( u1_u7_X_14 ) , .ZN( u1_u7_u2_n100 ) );
  NOR2_X1 u1_u7_u2_U72 (.A2( u1_u7_X_16 ) , .A1( u1_u7_X_17 ) , .ZN( u1_u7_u2_n138 ) );
  NOR2_X1 u1_u7_u2_U73 (.A2( u1_u7_X_15 ) , .A1( u1_u7_X_18 ) , .ZN( u1_u7_u2_n104 ) );
  NOR2_X1 u1_u7_u2_U74 (.A2( u1_u7_X_14 ) , .ZN( u1_u7_u2_n103 ) , .A1( u1_u7_u2_n174 ) );
  NOR2_X1 u1_u7_u2_U75 (.A2( u1_u7_X_15 ) , .ZN( u1_u7_u2_n102 ) , .A1( u1_u7_u2_n165 ) );
  NOR2_X1 u1_u7_u2_U76 (.A2( u1_u7_X_17 ) , .ZN( u1_u7_u2_n114 ) , .A1( u1_u7_u2_n169 ) );
  AND2_X1 u1_u7_u2_U77 (.A1( u1_u7_X_15 ) , .ZN( u1_u7_u2_n105 ) , .A2( u1_u7_u2_n165 ) );
  AND2_X1 u1_u7_u2_U78 (.A2( u1_u7_X_15 ) , .A1( u1_u7_X_18 ) , .ZN( u1_u7_u2_n107 ) );
  AND2_X1 u1_u7_u2_U79 (.A1( u1_u7_X_14 ) , .ZN( u1_u7_u2_n106 ) , .A2( u1_u7_u2_n174 ) );
  AOI21_X1 u1_u7_u2_U8 (.ZN( u1_u7_u2_n124 ) , .B1( u1_u7_u2_n131 ) , .B2( u1_u7_u2_n143 ) , .A( u1_u7_u2_n172 ) );
  AND2_X1 u1_u7_u2_U80 (.A1( u1_u7_X_13 ) , .A2( u1_u7_X_14 ) , .ZN( u1_u7_u2_n108 ) );
  INV_X1 u1_u7_u2_U81 (.A( u1_u7_X_16 ) , .ZN( u1_u7_u2_n169 ) );
  INV_X1 u1_u7_u2_U82 (.A( u1_u7_X_17 ) , .ZN( u1_u7_u2_n166 ) );
  INV_X1 u1_u7_u2_U83 (.A( u1_u7_X_13 ) , .ZN( u1_u7_u2_n174 ) );
  INV_X1 u1_u7_u2_U84 (.A( u1_u7_X_18 ) , .ZN( u1_u7_u2_n165 ) );
  NAND4_X1 u1_u7_u2_U85 (.ZN( u1_out7_24 ) , .A4( u1_u7_u2_n111 ) , .A3( u1_u7_u2_n112 ) , .A1( u1_u7_u2_n130 ) , .A2( u1_u7_u2_n187 ) );
  AOI221_X1 u1_u7_u2_U86 (.A( u1_u7_u2_n109 ) , .B1( u1_u7_u2_n110 ) , .ZN( u1_u7_u2_n111 ) , .C1( u1_u7_u2_n134 ) , .C2( u1_u7_u2_n170 ) , .B2( u1_u7_u2_n173 ) );
  AOI21_X1 u1_u7_u2_U87 (.ZN( u1_u7_u2_n112 ) , .B2( u1_u7_u2_n156 ) , .A( u1_u7_u2_n164 ) , .B1( u1_u7_u2_n181 ) );
  NAND4_X1 u1_u7_u2_U88 (.ZN( u1_out7_30 ) , .A4( u1_u7_u2_n147 ) , .A3( u1_u7_u2_n148 ) , .A2( u1_u7_u2_n149 ) , .A1( u1_u7_u2_n187 ) );
  NOR3_X1 u1_u7_u2_U89 (.A3( u1_u7_u2_n144 ) , .A2( u1_u7_u2_n145 ) , .A1( u1_u7_u2_n146 ) , .ZN( u1_u7_u2_n147 ) );
  AOI21_X1 u1_u7_u2_U9 (.B2( u1_u7_u2_n123 ) , .ZN( u1_u7_u2_n125 ) , .A( u1_u7_u2_n171 ) , .B1( u1_u7_u2_n184 ) );
  AOI21_X1 u1_u7_u2_U90 (.B2( u1_u7_u2_n138 ) , .ZN( u1_u7_u2_n148 ) , .A( u1_u7_u2_n162 ) , .B1( u1_u7_u2_n182 ) );
  NAND4_X1 u1_u7_u2_U91 (.ZN( u1_out7_16 ) , .A4( u1_u7_u2_n128 ) , .A3( u1_u7_u2_n129 ) , .A1( u1_u7_u2_n130 ) , .A2( u1_u7_u2_n186 ) );
  AOI22_X1 u1_u7_u2_U92 (.A2( u1_u7_u2_n118 ) , .ZN( u1_u7_u2_n129 ) , .A1( u1_u7_u2_n140 ) , .B1( u1_u7_u2_n157 ) , .B2( u1_u7_u2_n170 ) );
  INV_X1 u1_u7_u2_U93 (.A( u1_u7_u2_n163 ) , .ZN( u1_u7_u2_n186 ) );
  OR4_X1 u1_u7_u2_U94 (.ZN( u1_out7_6 ) , .A4( u1_u7_u2_n161 ) , .A3( u1_u7_u2_n162 ) , .A2( u1_u7_u2_n163 ) , .A1( u1_u7_u2_n164 ) );
  OR3_X1 u1_u7_u2_U95 (.A2( u1_u7_u2_n159 ) , .A1( u1_u7_u2_n160 ) , .ZN( u1_u7_u2_n161 ) , .A3( u1_u7_u2_n183 ) );
  AOI21_X1 u1_u7_u2_U96 (.B2( u1_u7_u2_n154 ) , .B1( u1_u7_u2_n155 ) , .ZN( u1_u7_u2_n159 ) , .A( u1_u7_u2_n167 ) );
  NAND3_X1 u1_u7_u2_U97 (.A2( u1_u7_u2_n117 ) , .A1( u1_u7_u2_n122 ) , .A3( u1_u7_u2_n123 ) , .ZN( u1_u7_u2_n134 ) );
  NAND3_X1 u1_u7_u2_U98 (.ZN( u1_u7_u2_n110 ) , .A2( u1_u7_u2_n131 ) , .A3( u1_u7_u2_n139 ) , .A1( u1_u7_u2_n154 ) );
  NAND3_X1 u1_u7_u2_U99 (.A2( u1_u7_u2_n100 ) , .ZN( u1_u7_u2_n101 ) , .A1( u1_u7_u2_n104 ) , .A3( u1_u7_u2_n114 ) );
  OAI22_X1 u1_u7_u4_U10 (.B2( u1_u7_u4_n135 ) , .ZN( u1_u7_u4_n137 ) , .B1( u1_u7_u4_n153 ) , .A1( u1_u7_u4_n155 ) , .A2( u1_u7_u4_n171 ) );
  AND3_X1 u1_u7_u4_U11 (.A2( u1_u7_u4_n134 ) , .ZN( u1_u7_u4_n135 ) , .A3( u1_u7_u4_n145 ) , .A1( u1_u7_u4_n157 ) );
  NAND2_X1 u1_u7_u4_U12 (.ZN( u1_u7_u4_n132 ) , .A2( u1_u7_u4_n170 ) , .A1( u1_u7_u4_n173 ) );
  AOI21_X1 u1_u7_u4_U13 (.B2( u1_u7_u4_n160 ) , .B1( u1_u7_u4_n161 ) , .ZN( u1_u7_u4_n162 ) , .A( u1_u7_u4_n170 ) );
  AOI21_X1 u1_u7_u4_U14 (.ZN( u1_u7_u4_n107 ) , .B2( u1_u7_u4_n143 ) , .A( u1_u7_u4_n174 ) , .B1( u1_u7_u4_n184 ) );
  AOI21_X1 u1_u7_u4_U15 (.B2( u1_u7_u4_n158 ) , .B1( u1_u7_u4_n159 ) , .ZN( u1_u7_u4_n163 ) , .A( u1_u7_u4_n174 ) );
  AOI21_X1 u1_u7_u4_U16 (.A( u1_u7_u4_n153 ) , .B2( u1_u7_u4_n154 ) , .B1( u1_u7_u4_n155 ) , .ZN( u1_u7_u4_n165 ) );
  AOI21_X1 u1_u7_u4_U17 (.A( u1_u7_u4_n156 ) , .B2( u1_u7_u4_n157 ) , .ZN( u1_u7_u4_n164 ) , .B1( u1_u7_u4_n184 ) );
  INV_X1 u1_u7_u4_U18 (.A( u1_u7_u4_n138 ) , .ZN( u1_u7_u4_n170 ) );
  AND2_X1 u1_u7_u4_U19 (.A2( u1_u7_u4_n120 ) , .ZN( u1_u7_u4_n155 ) , .A1( u1_u7_u4_n160 ) );
  INV_X1 u1_u7_u4_U20 (.A( u1_u7_u4_n156 ) , .ZN( u1_u7_u4_n175 ) );
  NAND2_X1 u1_u7_u4_U21 (.A2( u1_u7_u4_n118 ) , .ZN( u1_u7_u4_n131 ) , .A1( u1_u7_u4_n147 ) );
  NAND2_X1 u1_u7_u4_U22 (.A1( u1_u7_u4_n119 ) , .A2( u1_u7_u4_n120 ) , .ZN( u1_u7_u4_n130 ) );
  NAND2_X1 u1_u7_u4_U23 (.ZN( u1_u7_u4_n117 ) , .A2( u1_u7_u4_n118 ) , .A1( u1_u7_u4_n148 ) );
  NAND2_X1 u1_u7_u4_U24 (.ZN( u1_u7_u4_n129 ) , .A1( u1_u7_u4_n134 ) , .A2( u1_u7_u4_n148 ) );
  AND3_X1 u1_u7_u4_U25 (.A1( u1_u7_u4_n119 ) , .A2( u1_u7_u4_n143 ) , .A3( u1_u7_u4_n154 ) , .ZN( u1_u7_u4_n161 ) );
  AND2_X1 u1_u7_u4_U26 (.A1( u1_u7_u4_n145 ) , .A2( u1_u7_u4_n147 ) , .ZN( u1_u7_u4_n159 ) );
  OR3_X1 u1_u7_u4_U27 (.A3( u1_u7_u4_n114 ) , .A2( u1_u7_u4_n115 ) , .A1( u1_u7_u4_n116 ) , .ZN( u1_u7_u4_n136 ) );
  AOI21_X1 u1_u7_u4_U28 (.A( u1_u7_u4_n113 ) , .ZN( u1_u7_u4_n116 ) , .B2( u1_u7_u4_n173 ) , .B1( u1_u7_u4_n174 ) );
  AOI21_X1 u1_u7_u4_U29 (.ZN( u1_u7_u4_n115 ) , .B2( u1_u7_u4_n145 ) , .B1( u1_u7_u4_n146 ) , .A( u1_u7_u4_n156 ) );
  NOR2_X1 u1_u7_u4_U3 (.ZN( u1_u7_u4_n121 ) , .A1( u1_u7_u4_n181 ) , .A2( u1_u7_u4_n182 ) );
  OAI22_X1 u1_u7_u4_U30 (.ZN( u1_u7_u4_n114 ) , .A2( u1_u7_u4_n121 ) , .B1( u1_u7_u4_n160 ) , .B2( u1_u7_u4_n170 ) , .A1( u1_u7_u4_n171 ) );
  INV_X1 u1_u7_u4_U31 (.A( u1_u7_u4_n158 ) , .ZN( u1_u7_u4_n182 ) );
  INV_X1 u1_u7_u4_U32 (.ZN( u1_u7_u4_n181 ) , .A( u1_u7_u4_n96 ) );
  INV_X1 u1_u7_u4_U33 (.A( u1_u7_u4_n144 ) , .ZN( u1_u7_u4_n179 ) );
  INV_X1 u1_u7_u4_U34 (.A( u1_u7_u4_n157 ) , .ZN( u1_u7_u4_n178 ) );
  NAND2_X1 u1_u7_u4_U35 (.A2( u1_u7_u4_n154 ) , .A1( u1_u7_u4_n96 ) , .ZN( u1_u7_u4_n97 ) );
  INV_X1 u1_u7_u4_U36 (.ZN( u1_u7_u4_n186 ) , .A( u1_u7_u4_n95 ) );
  OAI221_X1 u1_u7_u4_U37 (.C1( u1_u7_u4_n134 ) , .B1( u1_u7_u4_n158 ) , .B2( u1_u7_u4_n171 ) , .C2( u1_u7_u4_n173 ) , .A( u1_u7_u4_n94 ) , .ZN( u1_u7_u4_n95 ) );
  AOI222_X1 u1_u7_u4_U38 (.B2( u1_u7_u4_n132 ) , .A1( u1_u7_u4_n138 ) , .C2( u1_u7_u4_n175 ) , .A2( u1_u7_u4_n179 ) , .C1( u1_u7_u4_n181 ) , .B1( u1_u7_u4_n185 ) , .ZN( u1_u7_u4_n94 ) );
  INV_X1 u1_u7_u4_U39 (.A( u1_u7_u4_n113 ) , .ZN( u1_u7_u4_n185 ) );
  INV_X1 u1_u7_u4_U4 (.A( u1_u7_u4_n117 ) , .ZN( u1_u7_u4_n184 ) );
  INV_X1 u1_u7_u4_U40 (.A( u1_u7_u4_n143 ) , .ZN( u1_u7_u4_n183 ) );
  NOR2_X1 u1_u7_u4_U41 (.ZN( u1_u7_u4_n138 ) , .A1( u1_u7_u4_n168 ) , .A2( u1_u7_u4_n169 ) );
  NOR2_X1 u1_u7_u4_U42 (.A1( u1_u7_u4_n150 ) , .A2( u1_u7_u4_n152 ) , .ZN( u1_u7_u4_n153 ) );
  NOR2_X1 u1_u7_u4_U43 (.A2( u1_u7_u4_n128 ) , .A1( u1_u7_u4_n138 ) , .ZN( u1_u7_u4_n156 ) );
  AOI22_X1 u1_u7_u4_U44 (.B2( u1_u7_u4_n122 ) , .A1( u1_u7_u4_n123 ) , .ZN( u1_u7_u4_n124 ) , .B1( u1_u7_u4_n128 ) , .A2( u1_u7_u4_n172 ) );
  NAND2_X1 u1_u7_u4_U45 (.A2( u1_u7_u4_n120 ) , .ZN( u1_u7_u4_n123 ) , .A1( u1_u7_u4_n161 ) );
  INV_X1 u1_u7_u4_U46 (.A( u1_u7_u4_n153 ) , .ZN( u1_u7_u4_n172 ) );
  AOI22_X1 u1_u7_u4_U47 (.B2( u1_u7_u4_n132 ) , .A2( u1_u7_u4_n133 ) , .ZN( u1_u7_u4_n140 ) , .A1( u1_u7_u4_n150 ) , .B1( u1_u7_u4_n179 ) );
  NAND2_X1 u1_u7_u4_U48 (.ZN( u1_u7_u4_n133 ) , .A2( u1_u7_u4_n146 ) , .A1( u1_u7_u4_n154 ) );
  NAND2_X1 u1_u7_u4_U49 (.A1( u1_u7_u4_n103 ) , .ZN( u1_u7_u4_n154 ) , .A2( u1_u7_u4_n98 ) );
  NOR4_X1 u1_u7_u4_U5 (.A4( u1_u7_u4_n106 ) , .A3( u1_u7_u4_n107 ) , .A2( u1_u7_u4_n108 ) , .A1( u1_u7_u4_n109 ) , .ZN( u1_u7_u4_n110 ) );
  NAND2_X1 u1_u7_u4_U50 (.A1( u1_u7_u4_n101 ) , .ZN( u1_u7_u4_n158 ) , .A2( u1_u7_u4_n99 ) );
  AOI21_X1 u1_u7_u4_U51 (.ZN( u1_u7_u4_n127 ) , .A( u1_u7_u4_n136 ) , .B2( u1_u7_u4_n150 ) , .B1( u1_u7_u4_n180 ) );
  INV_X1 u1_u7_u4_U52 (.A( u1_u7_u4_n160 ) , .ZN( u1_u7_u4_n180 ) );
  NAND2_X1 u1_u7_u4_U53 (.A2( u1_u7_u4_n104 ) , .A1( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n146 ) );
  NAND2_X1 u1_u7_u4_U54 (.A2( u1_u7_u4_n101 ) , .A1( u1_u7_u4_n102 ) , .ZN( u1_u7_u4_n160 ) );
  NAND2_X1 u1_u7_u4_U55 (.ZN( u1_u7_u4_n134 ) , .A1( u1_u7_u4_n98 ) , .A2( u1_u7_u4_n99 ) );
  NAND2_X1 u1_u7_u4_U56 (.A1( u1_u7_u4_n103 ) , .A2( u1_u7_u4_n104 ) , .ZN( u1_u7_u4_n143 ) );
  NAND2_X1 u1_u7_u4_U57 (.A2( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n145 ) , .A1( u1_u7_u4_n98 ) );
  NAND2_X1 u1_u7_u4_U58 (.A1( u1_u7_u4_n100 ) , .A2( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n120 ) );
  NAND2_X1 u1_u7_u4_U59 (.A1( u1_u7_u4_n102 ) , .A2( u1_u7_u4_n104 ) , .ZN( u1_u7_u4_n148 ) );
  AOI21_X1 u1_u7_u4_U6 (.ZN( u1_u7_u4_n106 ) , .B2( u1_u7_u4_n146 ) , .B1( u1_u7_u4_n158 ) , .A( u1_u7_u4_n170 ) );
  NAND2_X1 u1_u7_u4_U60 (.A2( u1_u7_u4_n100 ) , .A1( u1_u7_u4_n103 ) , .ZN( u1_u7_u4_n157 ) );
  INV_X1 u1_u7_u4_U61 (.A( u1_u7_u4_n150 ) , .ZN( u1_u7_u4_n173 ) );
  INV_X1 u1_u7_u4_U62 (.A( u1_u7_u4_n152 ) , .ZN( u1_u7_u4_n171 ) );
  NAND2_X1 u1_u7_u4_U63 (.A1( u1_u7_u4_n100 ) , .ZN( u1_u7_u4_n118 ) , .A2( u1_u7_u4_n99 ) );
  NAND2_X1 u1_u7_u4_U64 (.A2( u1_u7_u4_n100 ) , .A1( u1_u7_u4_n102 ) , .ZN( u1_u7_u4_n144 ) );
  NAND2_X1 u1_u7_u4_U65 (.A2( u1_u7_u4_n101 ) , .A1( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n96 ) );
  INV_X1 u1_u7_u4_U66 (.A( u1_u7_u4_n128 ) , .ZN( u1_u7_u4_n174 ) );
  NAND2_X1 u1_u7_u4_U67 (.A2( u1_u7_u4_n102 ) , .ZN( u1_u7_u4_n119 ) , .A1( u1_u7_u4_n98 ) );
  NAND2_X1 u1_u7_u4_U68 (.A2( u1_u7_u4_n101 ) , .A1( u1_u7_u4_n103 ) , .ZN( u1_u7_u4_n147 ) );
  NAND2_X1 u1_u7_u4_U69 (.A2( u1_u7_u4_n104 ) , .ZN( u1_u7_u4_n113 ) , .A1( u1_u7_u4_n99 ) );
  AOI21_X1 u1_u7_u4_U7 (.ZN( u1_u7_u4_n108 ) , .B2( u1_u7_u4_n134 ) , .B1( u1_u7_u4_n155 ) , .A( u1_u7_u4_n156 ) );
  NOR2_X1 u1_u7_u4_U70 (.A2( u1_u7_X_28 ) , .ZN( u1_u7_u4_n150 ) , .A1( u1_u7_u4_n168 ) );
  NOR2_X1 u1_u7_u4_U71 (.A2( u1_u7_X_29 ) , .ZN( u1_u7_u4_n152 ) , .A1( u1_u7_u4_n169 ) );
  NOR2_X1 u1_u7_u4_U72 (.A2( u1_u7_X_26 ) , .ZN( u1_u7_u4_n100 ) , .A1( u1_u7_u4_n177 ) );
  NOR2_X1 u1_u7_u4_U73 (.A2( u1_u7_X_30 ) , .ZN( u1_u7_u4_n105 ) , .A1( u1_u7_u4_n176 ) );
  NOR2_X1 u1_u7_u4_U74 (.A2( u1_u7_X_28 ) , .A1( u1_u7_X_29 ) , .ZN( u1_u7_u4_n128 ) );
  NOR2_X1 u1_u7_u4_U75 (.A2( u1_u7_X_25 ) , .A1( u1_u7_X_26 ) , .ZN( u1_u7_u4_n98 ) );
  NOR2_X1 u1_u7_u4_U76 (.A2( u1_u7_X_27 ) , .A1( u1_u7_X_30 ) , .ZN( u1_u7_u4_n102 ) );
  AND2_X1 u1_u7_u4_U77 (.A2( u1_u7_X_25 ) , .A1( u1_u7_X_26 ) , .ZN( u1_u7_u4_n104 ) );
  AND2_X1 u1_u7_u4_U78 (.A1( u1_u7_X_30 ) , .A2( u1_u7_u4_n176 ) , .ZN( u1_u7_u4_n99 ) );
  AND2_X1 u1_u7_u4_U79 (.A1( u1_u7_X_26 ) , .ZN( u1_u7_u4_n101 ) , .A2( u1_u7_u4_n177 ) );
  AOI21_X1 u1_u7_u4_U8 (.ZN( u1_u7_u4_n109 ) , .A( u1_u7_u4_n153 ) , .B1( u1_u7_u4_n159 ) , .B2( u1_u7_u4_n184 ) );
  AND2_X1 u1_u7_u4_U80 (.A1( u1_u7_X_27 ) , .A2( u1_u7_X_30 ) , .ZN( u1_u7_u4_n103 ) );
  INV_X1 u1_u7_u4_U81 (.A( u1_u7_X_28 ) , .ZN( u1_u7_u4_n169 ) );
  INV_X1 u1_u7_u4_U82 (.A( u1_u7_X_29 ) , .ZN( u1_u7_u4_n168 ) );
  INV_X1 u1_u7_u4_U83 (.A( u1_u7_X_25 ) , .ZN( u1_u7_u4_n177 ) );
  INV_X1 u1_u7_u4_U84 (.A( u1_u7_X_27 ) , .ZN( u1_u7_u4_n176 ) );
  NAND4_X1 u1_u7_u4_U85 (.ZN( u1_out7_25 ) , .A4( u1_u7_u4_n139 ) , .A3( u1_u7_u4_n140 ) , .A2( u1_u7_u4_n141 ) , .A1( u1_u7_u4_n142 ) );
  OAI21_X1 u1_u7_u4_U86 (.A( u1_u7_u4_n128 ) , .B2( u1_u7_u4_n129 ) , .B1( u1_u7_u4_n130 ) , .ZN( u1_u7_u4_n142 ) );
  OAI21_X1 u1_u7_u4_U87 (.B2( u1_u7_u4_n131 ) , .ZN( u1_u7_u4_n141 ) , .A( u1_u7_u4_n175 ) , .B1( u1_u7_u4_n183 ) );
  NAND4_X1 u1_u7_u4_U88 (.ZN( u1_out7_14 ) , .A4( u1_u7_u4_n124 ) , .A3( u1_u7_u4_n125 ) , .A2( u1_u7_u4_n126 ) , .A1( u1_u7_u4_n127 ) );
  AOI22_X1 u1_u7_u4_U89 (.B2( u1_u7_u4_n117 ) , .ZN( u1_u7_u4_n126 ) , .A1( u1_u7_u4_n129 ) , .B1( u1_u7_u4_n152 ) , .A2( u1_u7_u4_n175 ) );
  AOI211_X1 u1_u7_u4_U9 (.B( u1_u7_u4_n136 ) , .A( u1_u7_u4_n137 ) , .C2( u1_u7_u4_n138 ) , .ZN( u1_u7_u4_n139 ) , .C1( u1_u7_u4_n182 ) );
  AOI22_X1 u1_u7_u4_U90 (.ZN( u1_u7_u4_n125 ) , .B2( u1_u7_u4_n131 ) , .A2( u1_u7_u4_n132 ) , .B1( u1_u7_u4_n138 ) , .A1( u1_u7_u4_n178 ) );
  NAND4_X1 u1_u7_u4_U91 (.ZN( u1_out7_8 ) , .A4( u1_u7_u4_n110 ) , .A3( u1_u7_u4_n111 ) , .A2( u1_u7_u4_n112 ) , .A1( u1_u7_u4_n186 ) );
  NAND2_X1 u1_u7_u4_U92 (.ZN( u1_u7_u4_n112 ) , .A2( u1_u7_u4_n130 ) , .A1( u1_u7_u4_n150 ) );
  AOI22_X1 u1_u7_u4_U93 (.ZN( u1_u7_u4_n111 ) , .B2( u1_u7_u4_n132 ) , .A1( u1_u7_u4_n152 ) , .B1( u1_u7_u4_n178 ) , .A2( u1_u7_u4_n97 ) );
  AOI22_X1 u1_u7_u4_U94 (.B2( u1_u7_u4_n149 ) , .B1( u1_u7_u4_n150 ) , .A2( u1_u7_u4_n151 ) , .A1( u1_u7_u4_n152 ) , .ZN( u1_u7_u4_n167 ) );
  NOR4_X1 u1_u7_u4_U95 (.A4( u1_u7_u4_n162 ) , .A3( u1_u7_u4_n163 ) , .A2( u1_u7_u4_n164 ) , .A1( u1_u7_u4_n165 ) , .ZN( u1_u7_u4_n166 ) );
  NAND3_X1 u1_u7_u4_U96 (.ZN( u1_out7_3 ) , .A3( u1_u7_u4_n166 ) , .A1( u1_u7_u4_n167 ) , .A2( u1_u7_u4_n186 ) );
  NAND3_X1 u1_u7_u4_U97 (.A3( u1_u7_u4_n146 ) , .A2( u1_u7_u4_n147 ) , .A1( u1_u7_u4_n148 ) , .ZN( u1_u7_u4_n149 ) );
  NAND3_X1 u1_u7_u4_U98 (.A3( u1_u7_u4_n143 ) , .A2( u1_u7_u4_n144 ) , .A1( u1_u7_u4_n145 ) , .ZN( u1_u7_u4_n151 ) );
  NAND3_X1 u1_u7_u4_U99 (.A3( u1_u7_u4_n121 ) , .ZN( u1_u7_u4_n122 ) , .A2( u1_u7_u4_n144 ) , .A1( u1_u7_u4_n154 ) );
  INV_X1 u1_u7_u6_U10 (.ZN( u1_u7_u6_n172 ) , .A( u1_u7_u6_n88 ) );
  OAI21_X1 u1_u7_u6_U11 (.A( u1_u7_u6_n159 ) , .B1( u1_u7_u6_n169 ) , .B2( u1_u7_u6_n173 ) , .ZN( u1_u7_u6_n90 ) );
  AOI22_X1 u1_u7_u6_U12 (.A2( u1_u7_u6_n151 ) , .B2( u1_u7_u6_n161 ) , .A1( u1_u7_u6_n167 ) , .B1( u1_u7_u6_n170 ) , .ZN( u1_u7_u6_n89 ) );
  AOI21_X1 u1_u7_u6_U13 (.ZN( u1_u7_u6_n106 ) , .A( u1_u7_u6_n142 ) , .B2( u1_u7_u6_n159 ) , .B1( u1_u7_u6_n164 ) );
  INV_X1 u1_u7_u6_U14 (.A( u1_u7_u6_n155 ) , .ZN( u1_u7_u6_n161 ) );
  INV_X1 u1_u7_u6_U15 (.A( u1_u7_u6_n128 ) , .ZN( u1_u7_u6_n164 ) );
  NAND2_X1 u1_u7_u6_U16 (.ZN( u1_u7_u6_n110 ) , .A1( u1_u7_u6_n122 ) , .A2( u1_u7_u6_n129 ) );
  NAND2_X1 u1_u7_u6_U17 (.ZN( u1_u7_u6_n124 ) , .A2( u1_u7_u6_n146 ) , .A1( u1_u7_u6_n148 ) );
  INV_X1 u1_u7_u6_U18 (.A( u1_u7_u6_n132 ) , .ZN( u1_u7_u6_n171 ) );
  AND2_X1 u1_u7_u6_U19 (.A1( u1_u7_u6_n100 ) , .ZN( u1_u7_u6_n130 ) , .A2( u1_u7_u6_n147 ) );
  INV_X1 u1_u7_u6_U20 (.A( u1_u7_u6_n127 ) , .ZN( u1_u7_u6_n173 ) );
  INV_X1 u1_u7_u6_U21 (.A( u1_u7_u6_n121 ) , .ZN( u1_u7_u6_n167 ) );
  INV_X1 u1_u7_u6_U22 (.A( u1_u7_u6_n100 ) , .ZN( u1_u7_u6_n169 ) );
  INV_X1 u1_u7_u6_U23 (.A( u1_u7_u6_n123 ) , .ZN( u1_u7_u6_n170 ) );
  INV_X1 u1_u7_u6_U24 (.A( u1_u7_u6_n113 ) , .ZN( u1_u7_u6_n168 ) );
  AND2_X1 u1_u7_u6_U25 (.A1( u1_u7_u6_n107 ) , .A2( u1_u7_u6_n119 ) , .ZN( u1_u7_u6_n133 ) );
  AND2_X1 u1_u7_u6_U26 (.A2( u1_u7_u6_n121 ) , .A1( u1_u7_u6_n122 ) , .ZN( u1_u7_u6_n131 ) );
  AND3_X1 u1_u7_u6_U27 (.ZN( u1_u7_u6_n120 ) , .A2( u1_u7_u6_n127 ) , .A1( u1_u7_u6_n132 ) , .A3( u1_u7_u6_n145 ) );
  INV_X1 u1_u7_u6_U28 (.A( u1_u7_u6_n146 ) , .ZN( u1_u7_u6_n163 ) );
  AOI222_X1 u1_u7_u6_U29 (.ZN( u1_u7_u6_n114 ) , .A1( u1_u7_u6_n118 ) , .A2( u1_u7_u6_n126 ) , .B2( u1_u7_u6_n151 ) , .C2( u1_u7_u6_n159 ) , .C1( u1_u7_u6_n168 ) , .B1( u1_u7_u6_n169 ) );
  INV_X1 u1_u7_u6_U3 (.A( u1_u7_u6_n110 ) , .ZN( u1_u7_u6_n166 ) );
  NOR2_X1 u1_u7_u6_U30 (.A1( u1_u7_u6_n162 ) , .A2( u1_u7_u6_n165 ) , .ZN( u1_u7_u6_n98 ) );
  NAND2_X1 u1_u7_u6_U31 (.A1( u1_u7_u6_n144 ) , .ZN( u1_u7_u6_n151 ) , .A2( u1_u7_u6_n158 ) );
  NAND2_X1 u1_u7_u6_U32 (.ZN( u1_u7_u6_n132 ) , .A1( u1_u7_u6_n91 ) , .A2( u1_u7_u6_n97 ) );
  AOI22_X1 u1_u7_u6_U33 (.B2( u1_u7_u6_n110 ) , .B1( u1_u7_u6_n111 ) , .A1( u1_u7_u6_n112 ) , .ZN( u1_u7_u6_n115 ) , .A2( u1_u7_u6_n161 ) );
  NAND4_X1 u1_u7_u6_U34 (.A3( u1_u7_u6_n109 ) , .ZN( u1_u7_u6_n112 ) , .A4( u1_u7_u6_n132 ) , .A2( u1_u7_u6_n147 ) , .A1( u1_u7_u6_n166 ) );
  NOR2_X1 u1_u7_u6_U35 (.ZN( u1_u7_u6_n109 ) , .A1( u1_u7_u6_n170 ) , .A2( u1_u7_u6_n173 ) );
  NOR2_X1 u1_u7_u6_U36 (.A2( u1_u7_u6_n126 ) , .ZN( u1_u7_u6_n155 ) , .A1( u1_u7_u6_n160 ) );
  NAND2_X1 u1_u7_u6_U37 (.ZN( u1_u7_u6_n146 ) , .A2( u1_u7_u6_n94 ) , .A1( u1_u7_u6_n99 ) );
  AOI21_X1 u1_u7_u6_U38 (.A( u1_u7_u6_n144 ) , .B2( u1_u7_u6_n145 ) , .B1( u1_u7_u6_n146 ) , .ZN( u1_u7_u6_n150 ) );
  AOI211_X1 u1_u7_u6_U39 (.B( u1_u7_u6_n134 ) , .A( u1_u7_u6_n135 ) , .C1( u1_u7_u6_n136 ) , .ZN( u1_u7_u6_n137 ) , .C2( u1_u7_u6_n151 ) );
  INV_X1 u1_u7_u6_U4 (.A( u1_u7_u6_n142 ) , .ZN( u1_u7_u6_n174 ) );
  NAND4_X1 u1_u7_u6_U40 (.A4( u1_u7_u6_n127 ) , .A3( u1_u7_u6_n128 ) , .A2( u1_u7_u6_n129 ) , .A1( u1_u7_u6_n130 ) , .ZN( u1_u7_u6_n136 ) );
  AOI21_X1 u1_u7_u6_U41 (.B2( u1_u7_u6_n132 ) , .B1( u1_u7_u6_n133 ) , .ZN( u1_u7_u6_n134 ) , .A( u1_u7_u6_n158 ) );
  AOI21_X1 u1_u7_u6_U42 (.B1( u1_u7_u6_n131 ) , .ZN( u1_u7_u6_n135 ) , .A( u1_u7_u6_n144 ) , .B2( u1_u7_u6_n146 ) );
  INV_X1 u1_u7_u6_U43 (.A( u1_u7_u6_n111 ) , .ZN( u1_u7_u6_n158 ) );
  NAND2_X1 u1_u7_u6_U44 (.ZN( u1_u7_u6_n127 ) , .A1( u1_u7_u6_n91 ) , .A2( u1_u7_u6_n92 ) );
  NAND2_X1 u1_u7_u6_U45 (.ZN( u1_u7_u6_n129 ) , .A2( u1_u7_u6_n95 ) , .A1( u1_u7_u6_n96 ) );
  INV_X1 u1_u7_u6_U46 (.A( u1_u7_u6_n144 ) , .ZN( u1_u7_u6_n159 ) );
  NAND2_X1 u1_u7_u6_U47 (.ZN( u1_u7_u6_n145 ) , .A2( u1_u7_u6_n97 ) , .A1( u1_u7_u6_n98 ) );
  NAND2_X1 u1_u7_u6_U48 (.ZN( u1_u7_u6_n148 ) , .A2( u1_u7_u6_n92 ) , .A1( u1_u7_u6_n94 ) );
  NAND2_X1 u1_u7_u6_U49 (.ZN( u1_u7_u6_n108 ) , .A2( u1_u7_u6_n139 ) , .A1( u1_u7_u6_n144 ) );
  NAND2_X1 u1_u7_u6_U5 (.A2( u1_u7_u6_n143 ) , .ZN( u1_u7_u6_n152 ) , .A1( u1_u7_u6_n166 ) );
  NAND2_X1 u1_u7_u6_U50 (.ZN( u1_u7_u6_n121 ) , .A2( u1_u7_u6_n95 ) , .A1( u1_u7_u6_n97 ) );
  NAND2_X1 u1_u7_u6_U51 (.ZN( u1_u7_u6_n107 ) , .A2( u1_u7_u6_n92 ) , .A1( u1_u7_u6_n95 ) );
  AND2_X1 u1_u7_u6_U52 (.ZN( u1_u7_u6_n118 ) , .A2( u1_u7_u6_n91 ) , .A1( u1_u7_u6_n99 ) );
  NAND2_X1 u1_u7_u6_U53 (.ZN( u1_u7_u6_n147 ) , .A2( u1_u7_u6_n98 ) , .A1( u1_u7_u6_n99 ) );
  NAND2_X1 u1_u7_u6_U54 (.ZN( u1_u7_u6_n128 ) , .A1( u1_u7_u6_n94 ) , .A2( u1_u7_u6_n96 ) );
  NAND2_X1 u1_u7_u6_U55 (.ZN( u1_u7_u6_n119 ) , .A2( u1_u7_u6_n95 ) , .A1( u1_u7_u6_n99 ) );
  NAND2_X1 u1_u7_u6_U56 (.ZN( u1_u7_u6_n123 ) , .A2( u1_u7_u6_n91 ) , .A1( u1_u7_u6_n96 ) );
  NAND2_X1 u1_u7_u6_U57 (.ZN( u1_u7_u6_n100 ) , .A2( u1_u7_u6_n92 ) , .A1( u1_u7_u6_n98 ) );
  NAND2_X1 u1_u7_u6_U58 (.ZN( u1_u7_u6_n122 ) , .A1( u1_u7_u6_n94 ) , .A2( u1_u7_u6_n97 ) );
  INV_X1 u1_u7_u6_U59 (.A( u1_u7_u6_n139 ) , .ZN( u1_u7_u6_n160 ) );
  AOI22_X1 u1_u7_u6_U6 (.B2( u1_u7_u6_n101 ) , .A1( u1_u7_u6_n102 ) , .ZN( u1_u7_u6_n103 ) , .B1( u1_u7_u6_n160 ) , .A2( u1_u7_u6_n161 ) );
  NAND2_X1 u1_u7_u6_U60 (.ZN( u1_u7_u6_n113 ) , .A1( u1_u7_u6_n96 ) , .A2( u1_u7_u6_n98 ) );
  NOR2_X1 u1_u7_u6_U61 (.A2( u1_u7_X_40 ) , .A1( u1_u7_X_41 ) , .ZN( u1_u7_u6_n126 ) );
  NOR2_X1 u1_u7_u6_U62 (.A2( u1_u7_X_39 ) , .A1( u1_u7_X_42 ) , .ZN( u1_u7_u6_n92 ) );
  NOR2_X1 u1_u7_u6_U63 (.A2( u1_u7_X_39 ) , .A1( u1_u7_u6_n156 ) , .ZN( u1_u7_u6_n97 ) );
  NOR2_X1 u1_u7_u6_U64 (.A2( u1_u7_X_38 ) , .A1( u1_u7_u6_n165 ) , .ZN( u1_u7_u6_n95 ) );
  NOR2_X1 u1_u7_u6_U65 (.A2( u1_u7_X_41 ) , .ZN( u1_u7_u6_n111 ) , .A1( u1_u7_u6_n157 ) );
  NOR2_X1 u1_u7_u6_U66 (.A2( u1_u7_X_37 ) , .A1( u1_u7_u6_n162 ) , .ZN( u1_u7_u6_n94 ) );
  NOR2_X1 u1_u7_u6_U67 (.A2( u1_u7_X_37 ) , .A1( u1_u7_X_38 ) , .ZN( u1_u7_u6_n91 ) );
  NAND2_X1 u1_u7_u6_U68 (.A1( u1_u7_X_41 ) , .ZN( u1_u7_u6_n144 ) , .A2( u1_u7_u6_n157 ) );
  NAND2_X1 u1_u7_u6_U69 (.A2( u1_u7_X_40 ) , .A1( u1_u7_X_41 ) , .ZN( u1_u7_u6_n139 ) );
  NOR2_X1 u1_u7_u6_U7 (.A1( u1_u7_u6_n118 ) , .ZN( u1_u7_u6_n143 ) , .A2( u1_u7_u6_n168 ) );
  AND2_X1 u1_u7_u6_U70 (.A1( u1_u7_X_39 ) , .A2( u1_u7_u6_n156 ) , .ZN( u1_u7_u6_n96 ) );
  AND2_X1 u1_u7_u6_U71 (.A1( u1_u7_X_39 ) , .A2( u1_u7_X_42 ) , .ZN( u1_u7_u6_n99 ) );
  INV_X1 u1_u7_u6_U72 (.A( u1_u7_X_40 ) , .ZN( u1_u7_u6_n157 ) );
  INV_X1 u1_u7_u6_U73 (.A( u1_u7_X_37 ) , .ZN( u1_u7_u6_n165 ) );
  INV_X1 u1_u7_u6_U74 (.A( u1_u7_X_38 ) , .ZN( u1_u7_u6_n162 ) );
  INV_X1 u1_u7_u6_U75 (.A( u1_u7_X_42 ) , .ZN( u1_u7_u6_n156 ) );
  NAND4_X1 u1_u7_u6_U76 (.ZN( u1_out7_12 ) , .A4( u1_u7_u6_n114 ) , .A3( u1_u7_u6_n115 ) , .A2( u1_u7_u6_n116 ) , .A1( u1_u7_u6_n117 ) );
  OAI22_X1 u1_u7_u6_U77 (.B2( u1_u7_u6_n111 ) , .ZN( u1_u7_u6_n116 ) , .B1( u1_u7_u6_n126 ) , .A2( u1_u7_u6_n164 ) , .A1( u1_u7_u6_n167 ) );
  OAI21_X1 u1_u7_u6_U78 (.A( u1_u7_u6_n108 ) , .ZN( u1_u7_u6_n117 ) , .B2( u1_u7_u6_n141 ) , .B1( u1_u7_u6_n163 ) );
  NAND4_X1 u1_u7_u6_U79 (.ZN( u1_out7_32 ) , .A4( u1_u7_u6_n103 ) , .A3( u1_u7_u6_n104 ) , .A2( u1_u7_u6_n105 ) , .A1( u1_u7_u6_n106 ) );
  AOI21_X1 u1_u7_u6_U8 (.B1( u1_u7_u6_n107 ) , .B2( u1_u7_u6_n132 ) , .A( u1_u7_u6_n158 ) , .ZN( u1_u7_u6_n88 ) );
  AOI22_X1 u1_u7_u6_U80 (.ZN( u1_u7_u6_n105 ) , .A2( u1_u7_u6_n108 ) , .A1( u1_u7_u6_n118 ) , .B2( u1_u7_u6_n126 ) , .B1( u1_u7_u6_n171 ) );
  AOI22_X1 u1_u7_u6_U81 (.ZN( u1_u7_u6_n104 ) , .A1( u1_u7_u6_n111 ) , .B1( u1_u7_u6_n124 ) , .B2( u1_u7_u6_n151 ) , .A2( u1_u7_u6_n93 ) );
  OAI211_X1 u1_u7_u6_U82 (.ZN( u1_out7_7 ) , .B( u1_u7_u6_n153 ) , .C2( u1_u7_u6_n154 ) , .C1( u1_u7_u6_n155 ) , .A( u1_u7_u6_n174 ) );
  NOR3_X1 u1_u7_u6_U83 (.A1( u1_u7_u6_n141 ) , .ZN( u1_u7_u6_n154 ) , .A3( u1_u7_u6_n164 ) , .A2( u1_u7_u6_n171 ) );
  AOI211_X1 u1_u7_u6_U84 (.B( u1_u7_u6_n149 ) , .A( u1_u7_u6_n150 ) , .C2( u1_u7_u6_n151 ) , .C1( u1_u7_u6_n152 ) , .ZN( u1_u7_u6_n153 ) );
  OAI211_X1 u1_u7_u6_U85 (.ZN( u1_out7_22 ) , .B( u1_u7_u6_n137 ) , .A( u1_u7_u6_n138 ) , .C2( u1_u7_u6_n139 ) , .C1( u1_u7_u6_n140 ) );
  AOI22_X1 u1_u7_u6_U86 (.B1( u1_u7_u6_n124 ) , .A2( u1_u7_u6_n125 ) , .A1( u1_u7_u6_n126 ) , .ZN( u1_u7_u6_n138 ) , .B2( u1_u7_u6_n161 ) );
  AND4_X1 u1_u7_u6_U87 (.A3( u1_u7_u6_n119 ) , .A1( u1_u7_u6_n120 ) , .A4( u1_u7_u6_n129 ) , .ZN( u1_u7_u6_n140 ) , .A2( u1_u7_u6_n143 ) );
  NAND3_X1 u1_u7_u6_U88 (.A2( u1_u7_u6_n123 ) , .ZN( u1_u7_u6_n125 ) , .A1( u1_u7_u6_n130 ) , .A3( u1_u7_u6_n131 ) );
  NAND3_X1 u1_u7_u6_U89 (.A3( u1_u7_u6_n133 ) , .ZN( u1_u7_u6_n141 ) , .A1( u1_u7_u6_n145 ) , .A2( u1_u7_u6_n148 ) );
  AOI21_X1 u1_u7_u6_U9 (.B2( u1_u7_u6_n147 ) , .B1( u1_u7_u6_n148 ) , .ZN( u1_u7_u6_n149 ) , .A( u1_u7_u6_n158 ) );
  NAND3_X1 u1_u7_u6_U90 (.ZN( u1_u7_u6_n101 ) , .A3( u1_u7_u6_n107 ) , .A2( u1_u7_u6_n121 ) , .A1( u1_u7_u6_n127 ) );
  NAND3_X1 u1_u7_u6_U91 (.ZN( u1_u7_u6_n102 ) , .A3( u1_u7_u6_n130 ) , .A2( u1_u7_u6_n145 ) , .A1( u1_u7_u6_n166 ) );
  NAND3_X1 u1_u7_u6_U92 (.A3( u1_u7_u6_n113 ) , .A1( u1_u7_u6_n119 ) , .A2( u1_u7_u6_n123 ) , .ZN( u1_u7_u6_n93 ) );
  NAND3_X1 u1_u7_u6_U93 (.ZN( u1_u7_u6_n142 ) , .A2( u1_u7_u6_n172 ) , .A3( u1_u7_u6_n89 ) , .A1( u1_u7_u6_n90 ) );
  XOR2_X1 u1_u8_U1 (.B( u1_K9_9 ) , .A( u1_R7_6 ) , .Z( u1_u8_X_9 ) );
  XOR2_X1 u1_u8_U10 (.B( u1_K9_45 ) , .A( u1_R7_30 ) , .Z( u1_u8_X_45 ) );
  XOR2_X1 u1_u8_U11 (.B( u1_K9_44 ) , .A( u1_R7_29 ) , .Z( u1_u8_X_44 ) );
  XOR2_X1 u1_u8_U12 (.B( u1_K9_43 ) , .A( u1_R7_28 ) , .Z( u1_u8_X_43 ) );
  XOR2_X1 u1_u8_U13 (.B( u1_K9_42 ) , .A( u1_R7_29 ) , .Z( u1_u8_X_42 ) );
  XOR2_X1 u1_u8_U14 (.B( u1_K9_41 ) , .A( u1_R7_28 ) , .Z( u1_u8_X_41 ) );
  XOR2_X1 u1_u8_U15 (.B( u1_K9_40 ) , .A( u1_R7_27 ) , .Z( u1_u8_X_40 ) );
  XOR2_X1 u1_u8_U17 (.B( u1_K9_39 ) , .A( u1_R7_26 ) , .Z( u1_u8_X_39 ) );
  XOR2_X1 u1_u8_U18 (.B( u1_K9_38 ) , .A( u1_R7_25 ) , .Z( u1_u8_X_38 ) );
  XOR2_X1 u1_u8_U19 (.B( u1_K9_37 ) , .A( u1_R7_24 ) , .Z( u1_u8_X_37 ) );
  XOR2_X1 u1_u8_U2 (.B( u1_K9_8 ) , .A( u1_R7_5 ) , .Z( u1_u8_X_8 ) );
  XOR2_X1 u1_u8_U20 (.B( u1_K9_36 ) , .A( u1_R7_25 ) , .Z( u1_u8_X_36 ) );
  XOR2_X1 u1_u8_U21 (.B( u1_K9_35 ) , .A( u1_R7_24 ) , .Z( u1_u8_X_35 ) );
  XOR2_X1 u1_u8_U24 (.B( u1_K9_32 ) , .A( u1_R7_21 ) , .Z( u1_u8_X_32 ) );
  XOR2_X1 u1_u8_U25 (.B( u1_K9_31 ) , .A( u1_R7_20 ) , .Z( u1_u8_X_31 ) );
  XOR2_X1 u1_u8_U26 (.B( u1_K9_30 ) , .A( u1_R7_21 ) , .Z( u1_u8_X_30 ) );
  XOR2_X1 u1_u8_U27 (.B( u1_K9_2 ) , .A( u1_R7_1 ) , .Z( u1_u8_X_2 ) );
  XOR2_X1 u1_u8_U28 (.B( u1_K9_29 ) , .A( u1_R7_20 ) , .Z( u1_u8_X_29 ) );
  XOR2_X1 u1_u8_U3 (.B( u1_K9_7 ) , .A( u1_R7_4 ) , .Z( u1_u8_X_7 ) );
  XOR2_X1 u1_u8_U31 (.B( u1_K9_26 ) , .A( u1_R7_17 ) , .Z( u1_u8_X_26 ) );
  XOR2_X1 u1_u8_U32 (.B( u1_K9_25 ) , .A( u1_R7_16 ) , .Z( u1_u8_X_25 ) );
  XOR2_X1 u1_u8_U33 (.B( u1_K9_24 ) , .A( u1_R7_17 ) , .Z( u1_u8_X_24 ) );
  XOR2_X1 u1_u8_U34 (.B( u1_K9_23 ) , .A( u1_R7_16 ) , .Z( u1_u8_X_23 ) );
  XOR2_X1 u1_u8_U35 (.B( u1_K9_22 ) , .A( u1_R7_15 ) , .Z( u1_u8_X_22 ) );
  XOR2_X1 u1_u8_U36 (.B( u1_K9_21 ) , .A( u1_R7_14 ) , .Z( u1_u8_X_21 ) );
  XOR2_X1 u1_u8_U37 (.B( u1_K9_20 ) , .A( u1_R7_13 ) , .Z( u1_u8_X_20 ) );
  XOR2_X1 u1_u8_U38 (.B( u1_K9_1 ) , .A( u1_R7_32 ) , .Z( u1_u8_X_1 ) );
  XOR2_X1 u1_u8_U39 (.B( u1_K9_19 ) , .A( u1_R7_12 ) , .Z( u1_u8_X_19 ) );
  XOR2_X1 u1_u8_U4 (.B( u1_K9_6 ) , .A( u1_R7_5 ) , .Z( u1_u8_X_6 ) );
  XOR2_X1 u1_u8_U40 (.B( u1_K9_18 ) , .A( u1_R7_13 ) , .Z( u1_u8_X_18 ) );
  XOR2_X1 u1_u8_U41 (.B( u1_K9_17 ) , .A( u1_R7_12 ) , .Z( u1_u8_X_17 ) );
  XOR2_X1 u1_u8_U42 (.B( u1_K9_16 ) , .A( u1_R7_11 ) , .Z( u1_u8_X_16 ) );
  XOR2_X1 u1_u8_U43 (.B( u1_K9_15 ) , .A( u1_R7_10 ) , .Z( u1_u8_X_15 ) );
  XOR2_X1 u1_u8_U44 (.B( u1_K9_14 ) , .A( u1_R7_9 ) , .Z( u1_u8_X_14 ) );
  XOR2_X1 u1_u8_U45 (.B( u1_K9_13 ) , .A( u1_R7_8 ) , .Z( u1_u8_X_13 ) );
  XOR2_X1 u1_u8_U46 (.B( u1_K9_12 ) , .A( u1_R7_9 ) , .Z( u1_u8_X_12 ) );
  XOR2_X1 u1_u8_U47 (.B( u1_K9_11 ) , .A( u1_R7_8 ) , .Z( u1_u8_X_11 ) );
  XOR2_X1 u1_u8_U48 (.B( u1_K9_10 ) , .A( u1_R7_7 ) , .Z( u1_u8_X_10 ) );
  XOR2_X1 u1_u8_U5 (.B( u1_K9_5 ) , .A( u1_R7_4 ) , .Z( u1_u8_X_5 ) );
  XOR2_X1 u1_u8_U7 (.B( u1_K9_48 ) , .A( u1_R7_1 ) , .Z( u1_u8_X_48 ) );
  XOR2_X1 u1_u8_U8 (.B( u1_K9_47 ) , .A( u1_R7_32 ) , .Z( u1_u8_X_47 ) );
  XOR2_X1 u1_u8_U9 (.B( u1_K9_46 ) , .A( u1_R7_31 ) , .Z( u1_u8_X_46 ) );
  AOI21_X1 u1_u8_u1_U10 (.B2( u1_u8_u1_n155 ) , .B1( u1_u8_u1_n156 ) , .ZN( u1_u8_u1_n157 ) , .A( u1_u8_u1_n174 ) );
  NAND3_X1 u1_u8_u1_U100 (.ZN( u1_u8_u1_n113 ) , .A1( u1_u8_u1_n120 ) , .A3( u1_u8_u1_n133 ) , .A2( u1_u8_u1_n155 ) );
  NAND2_X1 u1_u8_u1_U11 (.ZN( u1_u8_u1_n140 ) , .A2( u1_u8_u1_n150 ) , .A1( u1_u8_u1_n155 ) );
  NAND2_X1 u1_u8_u1_U12 (.A1( u1_u8_u1_n131 ) , .ZN( u1_u8_u1_n147 ) , .A2( u1_u8_u1_n153 ) );
  AOI22_X1 u1_u8_u1_U13 (.B2( u1_u8_u1_n136 ) , .A2( u1_u8_u1_n137 ) , .ZN( u1_u8_u1_n143 ) , .A1( u1_u8_u1_n171 ) , .B1( u1_u8_u1_n173 ) );
  INV_X1 u1_u8_u1_U14 (.A( u1_u8_u1_n147 ) , .ZN( u1_u8_u1_n181 ) );
  INV_X1 u1_u8_u1_U15 (.A( u1_u8_u1_n139 ) , .ZN( u1_u8_u1_n174 ) );
  INV_X1 u1_u8_u1_U16 (.A( u1_u8_u1_n112 ) , .ZN( u1_u8_u1_n171 ) );
  NAND2_X1 u1_u8_u1_U17 (.ZN( u1_u8_u1_n141 ) , .A1( u1_u8_u1_n153 ) , .A2( u1_u8_u1_n156 ) );
  AND2_X1 u1_u8_u1_U18 (.A1( u1_u8_u1_n123 ) , .ZN( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n161 ) );
  NAND2_X1 u1_u8_u1_U19 (.A2( u1_u8_u1_n115 ) , .A1( u1_u8_u1_n116 ) , .ZN( u1_u8_u1_n148 ) );
  NAND2_X1 u1_u8_u1_U20 (.A2( u1_u8_u1_n133 ) , .A1( u1_u8_u1_n135 ) , .ZN( u1_u8_u1_n159 ) );
  NAND2_X1 u1_u8_u1_U21 (.A2( u1_u8_u1_n115 ) , .A1( u1_u8_u1_n120 ) , .ZN( u1_u8_u1_n132 ) );
  INV_X1 u1_u8_u1_U22 (.A( u1_u8_u1_n154 ) , .ZN( u1_u8_u1_n178 ) );
  INV_X1 u1_u8_u1_U23 (.A( u1_u8_u1_n151 ) , .ZN( u1_u8_u1_n183 ) );
  AND2_X1 u1_u8_u1_U24 (.A1( u1_u8_u1_n129 ) , .A2( u1_u8_u1_n133 ) , .ZN( u1_u8_u1_n149 ) );
  INV_X1 u1_u8_u1_U25 (.A( u1_u8_u1_n131 ) , .ZN( u1_u8_u1_n180 ) );
  OR4_X1 u1_u8_u1_U26 (.A4( u1_u8_u1_n106 ) , .A3( u1_u8_u1_n107 ) , .ZN( u1_u8_u1_n108 ) , .A1( u1_u8_u1_n117 ) , .A2( u1_u8_u1_n184 ) );
  AOI21_X1 u1_u8_u1_U27 (.ZN( u1_u8_u1_n106 ) , .A( u1_u8_u1_n112 ) , .B1( u1_u8_u1_n154 ) , .B2( u1_u8_u1_n156 ) );
  AOI21_X1 u1_u8_u1_U28 (.ZN( u1_u8_u1_n107 ) , .B1( u1_u8_u1_n134 ) , .B2( u1_u8_u1_n149 ) , .A( u1_u8_u1_n174 ) );
  INV_X1 u1_u8_u1_U29 (.A( u1_u8_u1_n101 ) , .ZN( u1_u8_u1_n184 ) );
  INV_X1 u1_u8_u1_U3 (.A( u1_u8_u1_n159 ) , .ZN( u1_u8_u1_n182 ) );
  AOI221_X1 u1_u8_u1_U30 (.B1( u1_u8_u1_n140 ) , .ZN( u1_u8_u1_n167 ) , .B2( u1_u8_u1_n172 ) , .C2( u1_u8_u1_n175 ) , .C1( u1_u8_u1_n178 ) , .A( u1_u8_u1_n188 ) );
  INV_X1 u1_u8_u1_U31 (.ZN( u1_u8_u1_n188 ) , .A( u1_u8_u1_n97 ) );
  AOI211_X1 u1_u8_u1_U32 (.A( u1_u8_u1_n118 ) , .C1( u1_u8_u1_n132 ) , .C2( u1_u8_u1_n139 ) , .B( u1_u8_u1_n96 ) , .ZN( u1_u8_u1_n97 ) );
  AOI21_X1 u1_u8_u1_U33 (.B2( u1_u8_u1_n121 ) , .B1( u1_u8_u1_n135 ) , .A( u1_u8_u1_n152 ) , .ZN( u1_u8_u1_n96 ) );
  OAI221_X1 u1_u8_u1_U34 (.A( u1_u8_u1_n119 ) , .C2( u1_u8_u1_n129 ) , .ZN( u1_u8_u1_n138 ) , .B2( u1_u8_u1_n152 ) , .C1( u1_u8_u1_n174 ) , .B1( u1_u8_u1_n187 ) );
  INV_X1 u1_u8_u1_U35 (.A( u1_u8_u1_n148 ) , .ZN( u1_u8_u1_n187 ) );
  AOI211_X1 u1_u8_u1_U36 (.B( u1_u8_u1_n117 ) , .A( u1_u8_u1_n118 ) , .ZN( u1_u8_u1_n119 ) , .C2( u1_u8_u1_n146 ) , .C1( u1_u8_u1_n159 ) );
  NOR2_X1 u1_u8_u1_U37 (.A1( u1_u8_u1_n168 ) , .A2( u1_u8_u1_n176 ) , .ZN( u1_u8_u1_n98 ) );
  AOI211_X1 u1_u8_u1_U38 (.B( u1_u8_u1_n162 ) , .A( u1_u8_u1_n163 ) , .C2( u1_u8_u1_n164 ) , .ZN( u1_u8_u1_n165 ) , .C1( u1_u8_u1_n171 ) );
  AOI21_X1 u1_u8_u1_U39 (.A( u1_u8_u1_n160 ) , .B2( u1_u8_u1_n161 ) , .ZN( u1_u8_u1_n162 ) , .B1( u1_u8_u1_n182 ) );
  AOI221_X1 u1_u8_u1_U4 (.A( u1_u8_u1_n138 ) , .C2( u1_u8_u1_n139 ) , .C1( u1_u8_u1_n140 ) , .B2( u1_u8_u1_n141 ) , .ZN( u1_u8_u1_n142 ) , .B1( u1_u8_u1_n175 ) );
  OR2_X1 u1_u8_u1_U40 (.A2( u1_u8_u1_n157 ) , .A1( u1_u8_u1_n158 ) , .ZN( u1_u8_u1_n163 ) );
  NAND2_X1 u1_u8_u1_U41 (.A1( u1_u8_u1_n128 ) , .ZN( u1_u8_u1_n146 ) , .A2( u1_u8_u1_n160 ) );
  NAND2_X1 u1_u8_u1_U42 (.A2( u1_u8_u1_n112 ) , .ZN( u1_u8_u1_n139 ) , .A1( u1_u8_u1_n152 ) );
  NAND2_X1 u1_u8_u1_U43 (.A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n156 ) , .A2( u1_u8_u1_n99 ) );
  NOR2_X1 u1_u8_u1_U44 (.ZN( u1_u8_u1_n117 ) , .A1( u1_u8_u1_n121 ) , .A2( u1_u8_u1_n160 ) );
  OAI21_X1 u1_u8_u1_U45 (.B2( u1_u8_u1_n123 ) , .ZN( u1_u8_u1_n145 ) , .B1( u1_u8_u1_n160 ) , .A( u1_u8_u1_n185 ) );
  INV_X1 u1_u8_u1_U46 (.A( u1_u8_u1_n122 ) , .ZN( u1_u8_u1_n185 ) );
  AOI21_X1 u1_u8_u1_U47 (.B2( u1_u8_u1_n120 ) , .B1( u1_u8_u1_n121 ) , .ZN( u1_u8_u1_n122 ) , .A( u1_u8_u1_n128 ) );
  AOI21_X1 u1_u8_u1_U48 (.A( u1_u8_u1_n128 ) , .B2( u1_u8_u1_n129 ) , .ZN( u1_u8_u1_n130 ) , .B1( u1_u8_u1_n150 ) );
  NAND2_X1 u1_u8_u1_U49 (.ZN( u1_u8_u1_n112 ) , .A1( u1_u8_u1_n169 ) , .A2( u1_u8_u1_n170 ) );
  AOI211_X1 u1_u8_u1_U5 (.ZN( u1_u8_u1_n124 ) , .A( u1_u8_u1_n138 ) , .C2( u1_u8_u1_n139 ) , .B( u1_u8_u1_n145 ) , .C1( u1_u8_u1_n147 ) );
  NAND2_X1 u1_u8_u1_U50 (.ZN( u1_u8_u1_n129 ) , .A2( u1_u8_u1_n95 ) , .A1( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U51 (.A1( u1_u8_u1_n102 ) , .ZN( u1_u8_u1_n154 ) , .A2( u1_u8_u1_n99 ) );
  NAND2_X1 u1_u8_u1_U52 (.A2( u1_u8_u1_n100 ) , .ZN( u1_u8_u1_n135 ) , .A1( u1_u8_u1_n99 ) );
  AOI21_X1 u1_u8_u1_U53 (.A( u1_u8_u1_n152 ) , .B2( u1_u8_u1_n153 ) , .B1( u1_u8_u1_n154 ) , .ZN( u1_u8_u1_n158 ) );
  INV_X1 u1_u8_u1_U54 (.A( u1_u8_u1_n160 ) , .ZN( u1_u8_u1_n175 ) );
  NAND2_X1 u1_u8_u1_U55 (.A1( u1_u8_u1_n100 ) , .ZN( u1_u8_u1_n116 ) , .A2( u1_u8_u1_n95 ) );
  NAND2_X1 u1_u8_u1_U56 (.A1( u1_u8_u1_n102 ) , .ZN( u1_u8_u1_n131 ) , .A2( u1_u8_u1_n95 ) );
  NAND2_X1 u1_u8_u1_U57 (.A2( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n121 ) , .A1( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U58 (.A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n153 ) , .A2( u1_u8_u1_n98 ) );
  NAND2_X1 u1_u8_u1_U59 (.A2( u1_u8_u1_n104 ) , .A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n133 ) );
  AOI22_X1 u1_u8_u1_U6 (.B2( u1_u8_u1_n113 ) , .A2( u1_u8_u1_n114 ) , .ZN( u1_u8_u1_n125 ) , .A1( u1_u8_u1_n171 ) , .B1( u1_u8_u1_n173 ) );
  NAND2_X1 u1_u8_u1_U60 (.ZN( u1_u8_u1_n150 ) , .A2( u1_u8_u1_n98 ) , .A1( u1_u8_u1_n99 ) );
  NAND2_X1 u1_u8_u1_U61 (.A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n155 ) , .A2( u1_u8_u1_n95 ) );
  OAI21_X1 u1_u8_u1_U62 (.ZN( u1_u8_u1_n109 ) , .B1( u1_u8_u1_n129 ) , .B2( u1_u8_u1_n160 ) , .A( u1_u8_u1_n167 ) );
  NAND2_X1 u1_u8_u1_U63 (.A2( u1_u8_u1_n100 ) , .A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n120 ) );
  NAND2_X1 u1_u8_u1_U64 (.A1( u1_u8_u1_n102 ) , .A2( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n115 ) );
  NAND2_X1 u1_u8_u1_U65 (.A2( u1_u8_u1_n100 ) , .A1( u1_u8_u1_n104 ) , .ZN( u1_u8_u1_n151 ) );
  NAND2_X1 u1_u8_u1_U66 (.A2( u1_u8_u1_n103 ) , .A1( u1_u8_u1_n105 ) , .ZN( u1_u8_u1_n161 ) );
  INV_X1 u1_u8_u1_U67 (.A( u1_u8_u1_n152 ) , .ZN( u1_u8_u1_n173 ) );
  INV_X1 u1_u8_u1_U68 (.A( u1_u8_u1_n128 ) , .ZN( u1_u8_u1_n172 ) );
  NAND2_X1 u1_u8_u1_U69 (.A2( u1_u8_u1_n102 ) , .A1( u1_u8_u1_n103 ) , .ZN( u1_u8_u1_n123 ) );
  NAND2_X1 u1_u8_u1_U7 (.ZN( u1_u8_u1_n114 ) , .A1( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n156 ) );
  NOR2_X1 u1_u8_u1_U70 (.A2( u1_u8_X_7 ) , .A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n95 ) );
  NOR2_X1 u1_u8_u1_U71 (.A1( u1_u8_X_12 ) , .A2( u1_u8_X_9 ) , .ZN( u1_u8_u1_n100 ) );
  NOR2_X1 u1_u8_u1_U72 (.A2( u1_u8_X_8 ) , .A1( u1_u8_u1_n177 ) , .ZN( u1_u8_u1_n99 ) );
  NOR2_X1 u1_u8_u1_U73 (.A2( u1_u8_X_12 ) , .ZN( u1_u8_u1_n102 ) , .A1( u1_u8_u1_n176 ) );
  NOR2_X1 u1_u8_u1_U74 (.A2( u1_u8_X_9 ) , .ZN( u1_u8_u1_n105 ) , .A1( u1_u8_u1_n168 ) );
  NAND2_X1 u1_u8_u1_U75 (.A1( u1_u8_X_10 ) , .ZN( u1_u8_u1_n160 ) , .A2( u1_u8_u1_n169 ) );
  NAND2_X1 u1_u8_u1_U76 (.A2( u1_u8_X_10 ) , .A1( u1_u8_X_11 ) , .ZN( u1_u8_u1_n152 ) );
  NAND2_X1 u1_u8_u1_U77 (.A1( u1_u8_X_11 ) , .ZN( u1_u8_u1_n128 ) , .A2( u1_u8_u1_n170 ) );
  AND2_X1 u1_u8_u1_U78 (.A2( u1_u8_X_7 ) , .A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n104 ) );
  AND2_X1 u1_u8_u1_U79 (.A1( u1_u8_X_8 ) , .ZN( u1_u8_u1_n103 ) , .A2( u1_u8_u1_n177 ) );
  NOR2_X1 u1_u8_u1_U8 (.A1( u1_u8_u1_n112 ) , .A2( u1_u8_u1_n116 ) , .ZN( u1_u8_u1_n118 ) );
  INV_X1 u1_u8_u1_U80 (.A( u1_u8_X_10 ) , .ZN( u1_u8_u1_n170 ) );
  INV_X1 u1_u8_u1_U81 (.A( u1_u8_X_9 ) , .ZN( u1_u8_u1_n176 ) );
  INV_X1 u1_u8_u1_U82 (.A( u1_u8_X_11 ) , .ZN( u1_u8_u1_n169 ) );
  INV_X1 u1_u8_u1_U83 (.A( u1_u8_X_12 ) , .ZN( u1_u8_u1_n168 ) );
  INV_X1 u1_u8_u1_U84 (.A( u1_u8_X_7 ) , .ZN( u1_u8_u1_n177 ) );
  NAND4_X1 u1_u8_u1_U85 (.ZN( u1_out8_28 ) , .A4( u1_u8_u1_n124 ) , .A3( u1_u8_u1_n125 ) , .A2( u1_u8_u1_n126 ) , .A1( u1_u8_u1_n127 ) );
  OAI21_X1 u1_u8_u1_U86 (.ZN( u1_u8_u1_n127 ) , .B2( u1_u8_u1_n139 ) , .B1( u1_u8_u1_n175 ) , .A( u1_u8_u1_n183 ) );
  OAI21_X1 u1_u8_u1_U87 (.ZN( u1_u8_u1_n126 ) , .B2( u1_u8_u1_n140 ) , .A( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n178 ) );
  NAND4_X1 u1_u8_u1_U88 (.ZN( u1_out8_18 ) , .A4( u1_u8_u1_n165 ) , .A3( u1_u8_u1_n166 ) , .A1( u1_u8_u1_n167 ) , .A2( u1_u8_u1_n186 ) );
  AOI22_X1 u1_u8_u1_U89 (.B2( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n147 ) , .A2( u1_u8_u1_n148 ) , .ZN( u1_u8_u1_n166 ) , .A1( u1_u8_u1_n172 ) );
  OAI21_X1 u1_u8_u1_U9 (.ZN( u1_u8_u1_n101 ) , .B1( u1_u8_u1_n141 ) , .A( u1_u8_u1_n146 ) , .B2( u1_u8_u1_n183 ) );
  INV_X1 u1_u8_u1_U90 (.A( u1_u8_u1_n145 ) , .ZN( u1_u8_u1_n186 ) );
  NAND4_X1 u1_u8_u1_U91 (.ZN( u1_out8_2 ) , .A4( u1_u8_u1_n142 ) , .A3( u1_u8_u1_n143 ) , .A2( u1_u8_u1_n144 ) , .A1( u1_u8_u1_n179 ) );
  OAI21_X1 u1_u8_u1_U92 (.B2( u1_u8_u1_n132 ) , .ZN( u1_u8_u1_n144 ) , .A( u1_u8_u1_n146 ) , .B1( u1_u8_u1_n180 ) );
  INV_X1 u1_u8_u1_U93 (.A( u1_u8_u1_n130 ) , .ZN( u1_u8_u1_n179 ) );
  OR4_X1 u1_u8_u1_U94 (.ZN( u1_out8_13 ) , .A4( u1_u8_u1_n108 ) , .A3( u1_u8_u1_n109 ) , .A2( u1_u8_u1_n110 ) , .A1( u1_u8_u1_n111 ) );
  AOI21_X1 u1_u8_u1_U95 (.ZN( u1_u8_u1_n111 ) , .A( u1_u8_u1_n128 ) , .B2( u1_u8_u1_n131 ) , .B1( u1_u8_u1_n135 ) );
  AOI21_X1 u1_u8_u1_U96 (.ZN( u1_u8_u1_n110 ) , .A( u1_u8_u1_n116 ) , .B1( u1_u8_u1_n152 ) , .B2( u1_u8_u1_n160 ) );
  NAND3_X1 u1_u8_u1_U97 (.A3( u1_u8_u1_n149 ) , .A2( u1_u8_u1_n150 ) , .A1( u1_u8_u1_n151 ) , .ZN( u1_u8_u1_n164 ) );
  NAND3_X1 u1_u8_u1_U98 (.A3( u1_u8_u1_n134 ) , .A2( u1_u8_u1_n135 ) , .ZN( u1_u8_u1_n136 ) , .A1( u1_u8_u1_n151 ) );
  NAND3_X1 u1_u8_u1_U99 (.A1( u1_u8_u1_n133 ) , .ZN( u1_u8_u1_n137 ) , .A2( u1_u8_u1_n154 ) , .A3( u1_u8_u1_n181 ) );
  OAI22_X1 u1_u8_u2_U10 (.B1( u1_u8_u2_n151 ) , .A2( u1_u8_u2_n152 ) , .A1( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n160 ) , .B2( u1_u8_u2_n168 ) );
  NAND3_X1 u1_u8_u2_U100 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n104 ) , .A3( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n98 ) );
  NOR3_X1 u1_u8_u2_U11 (.A1( u1_u8_u2_n150 ) , .ZN( u1_u8_u2_n151 ) , .A3( u1_u8_u2_n175 ) , .A2( u1_u8_u2_n188 ) );
  AOI21_X1 u1_u8_u2_U12 (.B2( u1_u8_u2_n123 ) , .ZN( u1_u8_u2_n125 ) , .A( u1_u8_u2_n171 ) , .B1( u1_u8_u2_n184 ) );
  INV_X1 u1_u8_u2_U13 (.A( u1_u8_u2_n150 ) , .ZN( u1_u8_u2_n184 ) );
  AOI21_X1 u1_u8_u2_U14 (.ZN( u1_u8_u2_n144 ) , .B2( u1_u8_u2_n155 ) , .A( u1_u8_u2_n172 ) , .B1( u1_u8_u2_n185 ) );
  AOI21_X1 u1_u8_u2_U15 (.B2( u1_u8_u2_n143 ) , .ZN( u1_u8_u2_n145 ) , .B1( u1_u8_u2_n152 ) , .A( u1_u8_u2_n171 ) );
  INV_X1 u1_u8_u2_U16 (.A( u1_u8_u2_n156 ) , .ZN( u1_u8_u2_n171 ) );
  INV_X1 u1_u8_u2_U17 (.A( u1_u8_u2_n120 ) , .ZN( u1_u8_u2_n188 ) );
  NAND2_X1 u1_u8_u2_U18 (.A2( u1_u8_u2_n122 ) , .ZN( u1_u8_u2_n150 ) , .A1( u1_u8_u2_n152 ) );
  INV_X1 u1_u8_u2_U19 (.A( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n170 ) );
  INV_X1 u1_u8_u2_U20 (.A( u1_u8_u2_n137 ) , .ZN( u1_u8_u2_n173 ) );
  NAND2_X1 u1_u8_u2_U21 (.A1( u1_u8_u2_n132 ) , .A2( u1_u8_u2_n139 ) , .ZN( u1_u8_u2_n157 ) );
  INV_X1 u1_u8_u2_U22 (.A( u1_u8_u2_n113 ) , .ZN( u1_u8_u2_n178 ) );
  INV_X1 u1_u8_u2_U23 (.A( u1_u8_u2_n139 ) , .ZN( u1_u8_u2_n175 ) );
  INV_X1 u1_u8_u2_U24 (.A( u1_u8_u2_n155 ) , .ZN( u1_u8_u2_n181 ) );
  INV_X1 u1_u8_u2_U25 (.A( u1_u8_u2_n119 ) , .ZN( u1_u8_u2_n177 ) );
  INV_X1 u1_u8_u2_U26 (.A( u1_u8_u2_n116 ) , .ZN( u1_u8_u2_n180 ) );
  INV_X1 u1_u8_u2_U27 (.A( u1_u8_u2_n131 ) , .ZN( u1_u8_u2_n179 ) );
  INV_X1 u1_u8_u2_U28 (.A( u1_u8_u2_n154 ) , .ZN( u1_u8_u2_n176 ) );
  NAND2_X1 u1_u8_u2_U29 (.A2( u1_u8_u2_n116 ) , .A1( u1_u8_u2_n117 ) , .ZN( u1_u8_u2_n118 ) );
  NOR2_X1 u1_u8_u2_U3 (.ZN( u1_u8_u2_n121 ) , .A2( u1_u8_u2_n177 ) , .A1( u1_u8_u2_n180 ) );
  INV_X1 u1_u8_u2_U30 (.A( u1_u8_u2_n132 ) , .ZN( u1_u8_u2_n182 ) );
  INV_X1 u1_u8_u2_U31 (.A( u1_u8_u2_n158 ) , .ZN( u1_u8_u2_n183 ) );
  OAI21_X1 u1_u8_u2_U32 (.A( u1_u8_u2_n156 ) , .B1( u1_u8_u2_n157 ) , .ZN( u1_u8_u2_n158 ) , .B2( u1_u8_u2_n179 ) );
  NOR2_X1 u1_u8_u2_U33 (.ZN( u1_u8_u2_n156 ) , .A1( u1_u8_u2_n166 ) , .A2( u1_u8_u2_n169 ) );
  NOR2_X1 u1_u8_u2_U34 (.A2( u1_u8_u2_n114 ) , .ZN( u1_u8_u2_n137 ) , .A1( u1_u8_u2_n140 ) );
  NOR2_X1 u1_u8_u2_U35 (.A2( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n153 ) , .A1( u1_u8_u2_n156 ) );
  AOI211_X1 u1_u8_u2_U36 (.ZN( u1_u8_u2_n130 ) , .C1( u1_u8_u2_n138 ) , .C2( u1_u8_u2_n179 ) , .B( u1_u8_u2_n96 ) , .A( u1_u8_u2_n97 ) );
  OAI22_X1 u1_u8_u2_U37 (.B1( u1_u8_u2_n133 ) , .A2( u1_u8_u2_n137 ) , .A1( u1_u8_u2_n152 ) , .B2( u1_u8_u2_n168 ) , .ZN( u1_u8_u2_n97 ) );
  OAI221_X1 u1_u8_u2_U38 (.B1( u1_u8_u2_n113 ) , .C1( u1_u8_u2_n132 ) , .A( u1_u8_u2_n149 ) , .B2( u1_u8_u2_n171 ) , .C2( u1_u8_u2_n172 ) , .ZN( u1_u8_u2_n96 ) );
  OAI221_X1 u1_u8_u2_U39 (.A( u1_u8_u2_n115 ) , .C2( u1_u8_u2_n123 ) , .B2( u1_u8_u2_n143 ) , .B1( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n163 ) , .C1( u1_u8_u2_n168 ) );
  INV_X1 u1_u8_u2_U4 (.A( u1_u8_u2_n134 ) , .ZN( u1_u8_u2_n185 ) );
  OAI21_X1 u1_u8_u2_U40 (.A( u1_u8_u2_n114 ) , .ZN( u1_u8_u2_n115 ) , .B1( u1_u8_u2_n176 ) , .B2( u1_u8_u2_n178 ) );
  OAI221_X1 u1_u8_u2_U41 (.A( u1_u8_u2_n135 ) , .B2( u1_u8_u2_n136 ) , .B1( u1_u8_u2_n137 ) , .ZN( u1_u8_u2_n162 ) , .C2( u1_u8_u2_n167 ) , .C1( u1_u8_u2_n185 ) );
  AND3_X1 u1_u8_u2_U42 (.A3( u1_u8_u2_n131 ) , .A2( u1_u8_u2_n132 ) , .A1( u1_u8_u2_n133 ) , .ZN( u1_u8_u2_n136 ) );
  AOI22_X1 u1_u8_u2_U43 (.ZN( u1_u8_u2_n135 ) , .B1( u1_u8_u2_n140 ) , .A1( u1_u8_u2_n156 ) , .B2( u1_u8_u2_n180 ) , .A2( u1_u8_u2_n188 ) );
  AOI21_X1 u1_u8_u2_U44 (.ZN( u1_u8_u2_n149 ) , .B1( u1_u8_u2_n173 ) , .B2( u1_u8_u2_n188 ) , .A( u1_u8_u2_n95 ) );
  AND3_X1 u1_u8_u2_U45 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n104 ) , .A3( u1_u8_u2_n156 ) , .ZN( u1_u8_u2_n95 ) );
  OAI21_X1 u1_u8_u2_U46 (.A( u1_u8_u2_n101 ) , .B2( u1_u8_u2_n121 ) , .B1( u1_u8_u2_n153 ) , .ZN( u1_u8_u2_n164 ) );
  NAND2_X1 u1_u8_u2_U47 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n107 ) , .ZN( u1_u8_u2_n155 ) );
  NAND2_X1 u1_u8_u2_U48 (.A2( u1_u8_u2_n105 ) , .A1( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n143 ) );
  NAND2_X1 u1_u8_u2_U49 (.A1( u1_u8_u2_n104 ) , .A2( u1_u8_u2_n106 ) , .ZN( u1_u8_u2_n152 ) );
  NOR4_X1 u1_u8_u2_U5 (.A4( u1_u8_u2_n124 ) , .A3( u1_u8_u2_n125 ) , .A2( u1_u8_u2_n126 ) , .A1( u1_u8_u2_n127 ) , .ZN( u1_u8_u2_n128 ) );
  NAND2_X1 u1_u8_u2_U50 (.A1( u1_u8_u2_n100 ) , .A2( u1_u8_u2_n105 ) , .ZN( u1_u8_u2_n132 ) );
  INV_X1 u1_u8_u2_U51 (.A( u1_u8_u2_n140 ) , .ZN( u1_u8_u2_n168 ) );
  INV_X1 u1_u8_u2_U52 (.A( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n167 ) );
  OAI21_X1 u1_u8_u2_U53 (.A( u1_u8_u2_n141 ) , .B2( u1_u8_u2_n142 ) , .ZN( u1_u8_u2_n146 ) , .B1( u1_u8_u2_n153 ) );
  OAI21_X1 u1_u8_u2_U54 (.A( u1_u8_u2_n140 ) , .ZN( u1_u8_u2_n141 ) , .B1( u1_u8_u2_n176 ) , .B2( u1_u8_u2_n177 ) );
  NOR3_X1 u1_u8_u2_U55 (.ZN( u1_u8_u2_n142 ) , .A3( u1_u8_u2_n175 ) , .A2( u1_u8_u2_n178 ) , .A1( u1_u8_u2_n181 ) );
  NAND2_X1 u1_u8_u2_U56 (.A1( u1_u8_u2_n102 ) , .A2( u1_u8_u2_n106 ) , .ZN( u1_u8_u2_n113 ) );
  NAND2_X1 u1_u8_u2_U57 (.A1( u1_u8_u2_n106 ) , .A2( u1_u8_u2_n107 ) , .ZN( u1_u8_u2_n131 ) );
  NAND2_X1 u1_u8_u2_U58 (.A1( u1_u8_u2_n103 ) , .A2( u1_u8_u2_n107 ) , .ZN( u1_u8_u2_n139 ) );
  NAND2_X1 u1_u8_u2_U59 (.A1( u1_u8_u2_n103 ) , .A2( u1_u8_u2_n105 ) , .ZN( u1_u8_u2_n133 ) );
  AOI21_X1 u1_u8_u2_U6 (.B2( u1_u8_u2_n119 ) , .ZN( u1_u8_u2_n127 ) , .A( u1_u8_u2_n137 ) , .B1( u1_u8_u2_n155 ) );
  NAND2_X1 u1_u8_u2_U60 (.A1( u1_u8_u2_n102 ) , .A2( u1_u8_u2_n103 ) , .ZN( u1_u8_u2_n154 ) );
  NAND2_X1 u1_u8_u2_U61 (.A2( u1_u8_u2_n103 ) , .A1( u1_u8_u2_n104 ) , .ZN( u1_u8_u2_n119 ) );
  NAND2_X1 u1_u8_u2_U62 (.A2( u1_u8_u2_n107 ) , .A1( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n123 ) );
  NAND2_X1 u1_u8_u2_U63 (.A1( u1_u8_u2_n104 ) , .A2( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n122 ) );
  INV_X1 u1_u8_u2_U64 (.A( u1_u8_u2_n114 ) , .ZN( u1_u8_u2_n172 ) );
  NAND2_X1 u1_u8_u2_U65 (.A2( u1_u8_u2_n100 ) , .A1( u1_u8_u2_n102 ) , .ZN( u1_u8_u2_n116 ) );
  NAND2_X1 u1_u8_u2_U66 (.A1( u1_u8_u2_n102 ) , .A2( u1_u8_u2_n108 ) , .ZN( u1_u8_u2_n120 ) );
  NAND2_X1 u1_u8_u2_U67 (.A2( u1_u8_u2_n105 ) , .A1( u1_u8_u2_n106 ) , .ZN( u1_u8_u2_n117 ) );
  INV_X1 u1_u8_u2_U68 (.ZN( u1_u8_u2_n187 ) , .A( u1_u8_u2_n99 ) );
  OAI21_X1 u1_u8_u2_U69 (.B1( u1_u8_u2_n137 ) , .B2( u1_u8_u2_n143 ) , .A( u1_u8_u2_n98 ) , .ZN( u1_u8_u2_n99 ) );
  AOI21_X1 u1_u8_u2_U7 (.ZN( u1_u8_u2_n124 ) , .B1( u1_u8_u2_n131 ) , .B2( u1_u8_u2_n143 ) , .A( u1_u8_u2_n172 ) );
  NOR2_X1 u1_u8_u2_U70 (.A2( u1_u8_X_16 ) , .ZN( u1_u8_u2_n140 ) , .A1( u1_u8_u2_n166 ) );
  NOR2_X1 u1_u8_u2_U71 (.A2( u1_u8_X_13 ) , .A1( u1_u8_X_14 ) , .ZN( u1_u8_u2_n100 ) );
  NOR2_X1 u1_u8_u2_U72 (.A2( u1_u8_X_16 ) , .A1( u1_u8_X_17 ) , .ZN( u1_u8_u2_n138 ) );
  NOR2_X1 u1_u8_u2_U73 (.A2( u1_u8_X_15 ) , .A1( u1_u8_X_18 ) , .ZN( u1_u8_u2_n104 ) );
  NOR2_X1 u1_u8_u2_U74 (.A2( u1_u8_X_14 ) , .ZN( u1_u8_u2_n103 ) , .A1( u1_u8_u2_n174 ) );
  NOR2_X1 u1_u8_u2_U75 (.A2( u1_u8_X_15 ) , .ZN( u1_u8_u2_n102 ) , .A1( u1_u8_u2_n165 ) );
  NOR2_X1 u1_u8_u2_U76 (.A2( u1_u8_X_17 ) , .ZN( u1_u8_u2_n114 ) , .A1( u1_u8_u2_n169 ) );
  AND2_X1 u1_u8_u2_U77 (.A1( u1_u8_X_15 ) , .ZN( u1_u8_u2_n105 ) , .A2( u1_u8_u2_n165 ) );
  AND2_X1 u1_u8_u2_U78 (.A2( u1_u8_X_15 ) , .A1( u1_u8_X_18 ) , .ZN( u1_u8_u2_n107 ) );
  AND2_X1 u1_u8_u2_U79 (.A1( u1_u8_X_14 ) , .ZN( u1_u8_u2_n106 ) , .A2( u1_u8_u2_n174 ) );
  AOI21_X1 u1_u8_u2_U8 (.B2( u1_u8_u2_n120 ) , .B1( u1_u8_u2_n121 ) , .ZN( u1_u8_u2_n126 ) , .A( u1_u8_u2_n167 ) );
  AND2_X1 u1_u8_u2_U80 (.A1( u1_u8_X_13 ) , .A2( u1_u8_X_14 ) , .ZN( u1_u8_u2_n108 ) );
  INV_X1 u1_u8_u2_U81 (.A( u1_u8_X_16 ) , .ZN( u1_u8_u2_n169 ) );
  INV_X1 u1_u8_u2_U82 (.A( u1_u8_X_17 ) , .ZN( u1_u8_u2_n166 ) );
  INV_X1 u1_u8_u2_U83 (.A( u1_u8_X_13 ) , .ZN( u1_u8_u2_n174 ) );
  INV_X1 u1_u8_u2_U84 (.A( u1_u8_X_18 ) , .ZN( u1_u8_u2_n165 ) );
  NAND4_X1 u1_u8_u2_U85 (.ZN( u1_out8_30 ) , .A4( u1_u8_u2_n147 ) , .A3( u1_u8_u2_n148 ) , .A2( u1_u8_u2_n149 ) , .A1( u1_u8_u2_n187 ) );
  NOR3_X1 u1_u8_u2_U86 (.A3( u1_u8_u2_n144 ) , .A2( u1_u8_u2_n145 ) , .A1( u1_u8_u2_n146 ) , .ZN( u1_u8_u2_n147 ) );
  AOI21_X1 u1_u8_u2_U87 (.B2( u1_u8_u2_n138 ) , .ZN( u1_u8_u2_n148 ) , .A( u1_u8_u2_n162 ) , .B1( u1_u8_u2_n182 ) );
  NAND4_X1 u1_u8_u2_U88 (.ZN( u1_out8_24 ) , .A4( u1_u8_u2_n111 ) , .A3( u1_u8_u2_n112 ) , .A1( u1_u8_u2_n130 ) , .A2( u1_u8_u2_n187 ) );
  AOI221_X1 u1_u8_u2_U89 (.A( u1_u8_u2_n109 ) , .B1( u1_u8_u2_n110 ) , .ZN( u1_u8_u2_n111 ) , .C1( u1_u8_u2_n134 ) , .C2( u1_u8_u2_n170 ) , .B2( u1_u8_u2_n173 ) );
  OAI22_X1 u1_u8_u2_U9 (.ZN( u1_u8_u2_n109 ) , .A2( u1_u8_u2_n113 ) , .B2( u1_u8_u2_n133 ) , .B1( u1_u8_u2_n167 ) , .A1( u1_u8_u2_n168 ) );
  AOI21_X1 u1_u8_u2_U90 (.ZN( u1_u8_u2_n112 ) , .B2( u1_u8_u2_n156 ) , .A( u1_u8_u2_n164 ) , .B1( u1_u8_u2_n181 ) );
  NAND4_X1 u1_u8_u2_U91 (.ZN( u1_out8_16 ) , .A4( u1_u8_u2_n128 ) , .A3( u1_u8_u2_n129 ) , .A1( u1_u8_u2_n130 ) , .A2( u1_u8_u2_n186 ) );
  AOI22_X1 u1_u8_u2_U92 (.A2( u1_u8_u2_n118 ) , .ZN( u1_u8_u2_n129 ) , .A1( u1_u8_u2_n140 ) , .B1( u1_u8_u2_n157 ) , .B2( u1_u8_u2_n170 ) );
  INV_X1 u1_u8_u2_U93 (.A( u1_u8_u2_n163 ) , .ZN( u1_u8_u2_n186 ) );
  OR4_X1 u1_u8_u2_U94 (.ZN( u1_out8_6 ) , .A4( u1_u8_u2_n161 ) , .A3( u1_u8_u2_n162 ) , .A2( u1_u8_u2_n163 ) , .A1( u1_u8_u2_n164 ) );
  OR3_X1 u1_u8_u2_U95 (.A2( u1_u8_u2_n159 ) , .A1( u1_u8_u2_n160 ) , .ZN( u1_u8_u2_n161 ) , .A3( u1_u8_u2_n183 ) );
  AOI21_X1 u1_u8_u2_U96 (.B2( u1_u8_u2_n154 ) , .B1( u1_u8_u2_n155 ) , .ZN( u1_u8_u2_n159 ) , .A( u1_u8_u2_n167 ) );
  NAND3_X1 u1_u8_u2_U97 (.A2( u1_u8_u2_n117 ) , .A1( u1_u8_u2_n122 ) , .A3( u1_u8_u2_n123 ) , .ZN( u1_u8_u2_n134 ) );
  NAND3_X1 u1_u8_u2_U98 (.ZN( u1_u8_u2_n110 ) , .A2( u1_u8_u2_n131 ) , .A3( u1_u8_u2_n139 ) , .A1( u1_u8_u2_n154 ) );
  NAND3_X1 u1_u8_u2_U99 (.A2( u1_u8_u2_n100 ) , .ZN( u1_u8_u2_n101 ) , .A1( u1_u8_u2_n104 ) , .A3( u1_u8_u2_n114 ) );
  OAI22_X1 u1_u8_u3_U10 (.B1( u1_u8_u3_n113 ) , .A2( u1_u8_u3_n135 ) , .A1( u1_u8_u3_n150 ) , .B2( u1_u8_u3_n164 ) , .ZN( u1_u8_u3_n98 ) );
  OAI211_X1 u1_u8_u3_U11 (.B( u1_u8_u3_n106 ) , .ZN( u1_u8_u3_n119 ) , .C2( u1_u8_u3_n128 ) , .C1( u1_u8_u3_n167 ) , .A( u1_u8_u3_n181 ) );
  AOI221_X1 u1_u8_u3_U12 (.C1( u1_u8_u3_n105 ) , .ZN( u1_u8_u3_n106 ) , .A( u1_u8_u3_n131 ) , .B2( u1_u8_u3_n132 ) , .C2( u1_u8_u3_n133 ) , .B1( u1_u8_u3_n169 ) );
  INV_X1 u1_u8_u3_U13 (.ZN( u1_u8_u3_n181 ) , .A( u1_u8_u3_n98 ) );
  NAND2_X1 u1_u8_u3_U14 (.ZN( u1_u8_u3_n105 ) , .A2( u1_u8_u3_n130 ) , .A1( u1_u8_u3_n155 ) );
  AOI22_X1 u1_u8_u3_U15 (.B1( u1_u8_u3_n115 ) , .A2( u1_u8_u3_n116 ) , .ZN( u1_u8_u3_n123 ) , .B2( u1_u8_u3_n133 ) , .A1( u1_u8_u3_n169 ) );
  NAND2_X1 u1_u8_u3_U16 (.ZN( u1_u8_u3_n116 ) , .A2( u1_u8_u3_n151 ) , .A1( u1_u8_u3_n182 ) );
  NOR2_X1 u1_u8_u3_U17 (.ZN( u1_u8_u3_n126 ) , .A2( u1_u8_u3_n150 ) , .A1( u1_u8_u3_n164 ) );
  AOI21_X1 u1_u8_u3_U18 (.ZN( u1_u8_u3_n112 ) , .B2( u1_u8_u3_n146 ) , .B1( u1_u8_u3_n155 ) , .A( u1_u8_u3_n167 ) );
  NAND2_X1 u1_u8_u3_U19 (.A1( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n142 ) , .A2( u1_u8_u3_n164 ) );
  NAND2_X1 u1_u8_u3_U20 (.ZN( u1_u8_u3_n132 ) , .A2( u1_u8_u3_n152 ) , .A1( u1_u8_u3_n156 ) );
  AND2_X1 u1_u8_u3_U21 (.A2( u1_u8_u3_n113 ) , .A1( u1_u8_u3_n114 ) , .ZN( u1_u8_u3_n151 ) );
  INV_X1 u1_u8_u3_U22 (.A( u1_u8_u3_n133 ) , .ZN( u1_u8_u3_n165 ) );
  INV_X1 u1_u8_u3_U23 (.A( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n170 ) );
  NAND2_X1 u1_u8_u3_U24 (.A1( u1_u8_u3_n107 ) , .A2( u1_u8_u3_n108 ) , .ZN( u1_u8_u3_n140 ) );
  NAND2_X1 u1_u8_u3_U25 (.ZN( u1_u8_u3_n117 ) , .A1( u1_u8_u3_n124 ) , .A2( u1_u8_u3_n148 ) );
  NAND2_X1 u1_u8_u3_U26 (.ZN( u1_u8_u3_n143 ) , .A1( u1_u8_u3_n165 ) , .A2( u1_u8_u3_n167 ) );
  INV_X1 u1_u8_u3_U27 (.A( u1_u8_u3_n130 ) , .ZN( u1_u8_u3_n177 ) );
  INV_X1 u1_u8_u3_U28 (.A( u1_u8_u3_n128 ) , .ZN( u1_u8_u3_n176 ) );
  INV_X1 u1_u8_u3_U29 (.A( u1_u8_u3_n155 ) , .ZN( u1_u8_u3_n174 ) );
  INV_X1 u1_u8_u3_U3 (.A( u1_u8_u3_n129 ) , .ZN( u1_u8_u3_n183 ) );
  INV_X1 u1_u8_u3_U30 (.A( u1_u8_u3_n139 ) , .ZN( u1_u8_u3_n185 ) );
  NOR2_X1 u1_u8_u3_U31 (.ZN( u1_u8_u3_n135 ) , .A2( u1_u8_u3_n141 ) , .A1( u1_u8_u3_n169 ) );
  OAI222_X1 u1_u8_u3_U32 (.C2( u1_u8_u3_n107 ) , .A2( u1_u8_u3_n108 ) , .B1( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n138 ) , .B2( u1_u8_u3_n146 ) , .C1( u1_u8_u3_n154 ) , .A1( u1_u8_u3_n164 ) );
  NOR4_X1 u1_u8_u3_U33 (.A4( u1_u8_u3_n157 ) , .A3( u1_u8_u3_n158 ) , .A2( u1_u8_u3_n159 ) , .A1( u1_u8_u3_n160 ) , .ZN( u1_u8_u3_n161 ) );
  AOI21_X1 u1_u8_u3_U34 (.B2( u1_u8_u3_n152 ) , .B1( u1_u8_u3_n153 ) , .ZN( u1_u8_u3_n158 ) , .A( u1_u8_u3_n164 ) );
  AOI21_X1 u1_u8_u3_U35 (.A( u1_u8_u3_n149 ) , .B2( u1_u8_u3_n150 ) , .B1( u1_u8_u3_n151 ) , .ZN( u1_u8_u3_n159 ) );
  AOI21_X1 u1_u8_u3_U36 (.A( u1_u8_u3_n154 ) , .B2( u1_u8_u3_n155 ) , .B1( u1_u8_u3_n156 ) , .ZN( u1_u8_u3_n157 ) );
  AOI211_X1 u1_u8_u3_U37 (.ZN( u1_u8_u3_n109 ) , .A( u1_u8_u3_n119 ) , .C2( u1_u8_u3_n129 ) , .B( u1_u8_u3_n138 ) , .C1( u1_u8_u3_n141 ) );
  AOI211_X1 u1_u8_u3_U38 (.B( u1_u8_u3_n119 ) , .A( u1_u8_u3_n120 ) , .C2( u1_u8_u3_n121 ) , .ZN( u1_u8_u3_n122 ) , .C1( u1_u8_u3_n179 ) );
  INV_X1 u1_u8_u3_U39 (.A( u1_u8_u3_n156 ) , .ZN( u1_u8_u3_n179 ) );
  INV_X1 u1_u8_u3_U4 (.A( u1_u8_u3_n140 ) , .ZN( u1_u8_u3_n182 ) );
  OAI22_X1 u1_u8_u3_U40 (.B1( u1_u8_u3_n118 ) , .ZN( u1_u8_u3_n120 ) , .A1( u1_u8_u3_n135 ) , .B2( u1_u8_u3_n154 ) , .A2( u1_u8_u3_n178 ) );
  AND3_X1 u1_u8_u3_U41 (.ZN( u1_u8_u3_n118 ) , .A2( u1_u8_u3_n124 ) , .A1( u1_u8_u3_n144 ) , .A3( u1_u8_u3_n152 ) );
  INV_X1 u1_u8_u3_U42 (.A( u1_u8_u3_n121 ) , .ZN( u1_u8_u3_n164 ) );
  NAND2_X1 u1_u8_u3_U43 (.ZN( u1_u8_u3_n133 ) , .A1( u1_u8_u3_n154 ) , .A2( u1_u8_u3_n164 ) );
  OAI211_X1 u1_u8_u3_U44 (.B( u1_u8_u3_n127 ) , .ZN( u1_u8_u3_n139 ) , .C1( u1_u8_u3_n150 ) , .C2( u1_u8_u3_n154 ) , .A( u1_u8_u3_n184 ) );
  INV_X1 u1_u8_u3_U45 (.A( u1_u8_u3_n125 ) , .ZN( u1_u8_u3_n184 ) );
  AOI221_X1 u1_u8_u3_U46 (.A( u1_u8_u3_n126 ) , .ZN( u1_u8_u3_n127 ) , .C2( u1_u8_u3_n132 ) , .C1( u1_u8_u3_n169 ) , .B2( u1_u8_u3_n170 ) , .B1( u1_u8_u3_n174 ) );
  OAI22_X1 u1_u8_u3_U47 (.A1( u1_u8_u3_n124 ) , .ZN( u1_u8_u3_n125 ) , .B2( u1_u8_u3_n145 ) , .A2( u1_u8_u3_n165 ) , .B1( u1_u8_u3_n167 ) );
  NOR2_X1 u1_u8_u3_U48 (.A1( u1_u8_u3_n113 ) , .ZN( u1_u8_u3_n131 ) , .A2( u1_u8_u3_n154 ) );
  NAND2_X1 u1_u8_u3_U49 (.A1( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n150 ) , .A2( u1_u8_u3_n99 ) );
  INV_X1 u1_u8_u3_U5 (.A( u1_u8_u3_n117 ) , .ZN( u1_u8_u3_n178 ) );
  NAND2_X1 u1_u8_u3_U50 (.A2( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n155 ) , .A1( u1_u8_u3_n97 ) );
  INV_X1 u1_u8_u3_U51 (.A( u1_u8_u3_n141 ) , .ZN( u1_u8_u3_n167 ) );
  AOI21_X1 u1_u8_u3_U52 (.B2( u1_u8_u3_n114 ) , .B1( u1_u8_u3_n146 ) , .A( u1_u8_u3_n154 ) , .ZN( u1_u8_u3_n94 ) );
  AOI21_X1 u1_u8_u3_U53 (.ZN( u1_u8_u3_n110 ) , .B2( u1_u8_u3_n142 ) , .B1( u1_u8_u3_n186 ) , .A( u1_u8_u3_n95 ) );
  INV_X1 u1_u8_u3_U54 (.A( u1_u8_u3_n145 ) , .ZN( u1_u8_u3_n186 ) );
  AOI21_X1 u1_u8_u3_U55 (.B1( u1_u8_u3_n124 ) , .A( u1_u8_u3_n149 ) , .B2( u1_u8_u3_n155 ) , .ZN( u1_u8_u3_n95 ) );
  INV_X1 u1_u8_u3_U56 (.A( u1_u8_u3_n149 ) , .ZN( u1_u8_u3_n169 ) );
  NAND2_X1 u1_u8_u3_U57 (.ZN( u1_u8_u3_n124 ) , .A1( u1_u8_u3_n96 ) , .A2( u1_u8_u3_n97 ) );
  NAND2_X1 u1_u8_u3_U58 (.A2( u1_u8_u3_n100 ) , .ZN( u1_u8_u3_n146 ) , .A1( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U59 (.A1( u1_u8_u3_n101 ) , .ZN( u1_u8_u3_n145 ) , .A2( u1_u8_u3_n99 ) );
  AOI221_X1 u1_u8_u3_U6 (.A( u1_u8_u3_n131 ) , .C2( u1_u8_u3_n132 ) , .C1( u1_u8_u3_n133 ) , .ZN( u1_u8_u3_n134 ) , .B1( u1_u8_u3_n143 ) , .B2( u1_u8_u3_n177 ) );
  NAND2_X1 u1_u8_u3_U60 (.A1( u1_u8_u3_n100 ) , .ZN( u1_u8_u3_n156 ) , .A2( u1_u8_u3_n99 ) );
  NAND2_X1 u1_u8_u3_U61 (.A2( u1_u8_u3_n101 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n148 ) );
  NAND2_X1 u1_u8_u3_U62 (.A1( u1_u8_u3_n100 ) , .A2( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n128 ) );
  NAND2_X1 u1_u8_u3_U63 (.A2( u1_u8_u3_n101 ) , .A1( u1_u8_u3_n102 ) , .ZN( u1_u8_u3_n152 ) );
  NAND2_X1 u1_u8_u3_U64 (.A2( u1_u8_u3_n101 ) , .ZN( u1_u8_u3_n114 ) , .A1( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U65 (.ZN( u1_u8_u3_n107 ) , .A1( u1_u8_u3_n97 ) , .A2( u1_u8_u3_n99 ) );
  NAND2_X1 u1_u8_u3_U66 (.A2( u1_u8_u3_n100 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n113 ) );
  NAND2_X1 u1_u8_u3_U67 (.A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n153 ) , .A2( u1_u8_u3_n97 ) );
  NAND2_X1 u1_u8_u3_U68 (.A2( u1_u8_u3_n103 ) , .A1( u1_u8_u3_n104 ) , .ZN( u1_u8_u3_n130 ) );
  NAND2_X1 u1_u8_u3_U69 (.A2( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n144 ) , .A1( u1_u8_u3_n96 ) );
  OAI22_X1 u1_u8_u3_U7 (.B2( u1_u8_u3_n147 ) , .A2( u1_u8_u3_n148 ) , .ZN( u1_u8_u3_n160 ) , .B1( u1_u8_u3_n165 ) , .A1( u1_u8_u3_n168 ) );
  NAND2_X1 u1_u8_u3_U70 (.A1( u1_u8_u3_n102 ) , .A2( u1_u8_u3_n103 ) , .ZN( u1_u8_u3_n108 ) );
  NOR2_X1 u1_u8_u3_U71 (.A2( u1_u8_X_19 ) , .A1( u1_u8_X_20 ) , .ZN( u1_u8_u3_n99 ) );
  NOR2_X1 u1_u8_u3_U72 (.A2( u1_u8_X_21 ) , .A1( u1_u8_X_24 ) , .ZN( u1_u8_u3_n103 ) );
  NOR2_X1 u1_u8_u3_U73 (.A2( u1_u8_X_24 ) , .A1( u1_u8_u3_n171 ) , .ZN( u1_u8_u3_n97 ) );
  NOR2_X1 u1_u8_u3_U74 (.A2( u1_u8_X_23 ) , .ZN( u1_u8_u3_n141 ) , .A1( u1_u8_u3_n166 ) );
  NOR2_X1 u1_u8_u3_U75 (.A2( u1_u8_X_19 ) , .A1( u1_u8_u3_n172 ) , .ZN( u1_u8_u3_n96 ) );
  NAND2_X1 u1_u8_u3_U76 (.A1( u1_u8_X_22 ) , .A2( u1_u8_X_23 ) , .ZN( u1_u8_u3_n154 ) );
  NAND2_X1 u1_u8_u3_U77 (.A1( u1_u8_X_23 ) , .ZN( u1_u8_u3_n149 ) , .A2( u1_u8_u3_n166 ) );
  NOR2_X1 u1_u8_u3_U78 (.A2( u1_u8_X_22 ) , .A1( u1_u8_X_23 ) , .ZN( u1_u8_u3_n121 ) );
  AND2_X1 u1_u8_u3_U79 (.A1( u1_u8_X_24 ) , .ZN( u1_u8_u3_n101 ) , .A2( u1_u8_u3_n171 ) );
  AND3_X1 u1_u8_u3_U8 (.A3( u1_u8_u3_n144 ) , .A2( u1_u8_u3_n145 ) , .A1( u1_u8_u3_n146 ) , .ZN( u1_u8_u3_n147 ) );
  AND2_X1 u1_u8_u3_U80 (.A1( u1_u8_X_19 ) , .ZN( u1_u8_u3_n102 ) , .A2( u1_u8_u3_n172 ) );
  AND2_X1 u1_u8_u3_U81 (.A1( u1_u8_X_21 ) , .A2( u1_u8_X_24 ) , .ZN( u1_u8_u3_n100 ) );
  AND2_X1 u1_u8_u3_U82 (.A2( u1_u8_X_19 ) , .A1( u1_u8_X_20 ) , .ZN( u1_u8_u3_n104 ) );
  INV_X1 u1_u8_u3_U83 (.A( u1_u8_X_22 ) , .ZN( u1_u8_u3_n166 ) );
  INV_X1 u1_u8_u3_U84 (.A( u1_u8_X_21 ) , .ZN( u1_u8_u3_n171 ) );
  INV_X1 u1_u8_u3_U85 (.A( u1_u8_X_20 ) , .ZN( u1_u8_u3_n172 ) );
  OR4_X1 u1_u8_u3_U86 (.ZN( u1_out8_10 ) , .A4( u1_u8_u3_n136 ) , .A3( u1_u8_u3_n137 ) , .A1( u1_u8_u3_n138 ) , .A2( u1_u8_u3_n139 ) );
  OAI222_X1 u1_u8_u3_U87 (.C1( u1_u8_u3_n128 ) , .ZN( u1_u8_u3_n137 ) , .B1( u1_u8_u3_n148 ) , .A2( u1_u8_u3_n150 ) , .B2( u1_u8_u3_n154 ) , .C2( u1_u8_u3_n164 ) , .A1( u1_u8_u3_n167 ) );
  OAI221_X1 u1_u8_u3_U88 (.A( u1_u8_u3_n134 ) , .B2( u1_u8_u3_n135 ) , .ZN( u1_u8_u3_n136 ) , .C1( u1_u8_u3_n149 ) , .B1( u1_u8_u3_n151 ) , .C2( u1_u8_u3_n183 ) );
  NAND4_X1 u1_u8_u3_U89 (.ZN( u1_out8_26 ) , .A4( u1_u8_u3_n109 ) , .A3( u1_u8_u3_n110 ) , .A2( u1_u8_u3_n111 ) , .A1( u1_u8_u3_n173 ) );
  INV_X1 u1_u8_u3_U9 (.A( u1_u8_u3_n143 ) , .ZN( u1_u8_u3_n168 ) );
  INV_X1 u1_u8_u3_U90 (.ZN( u1_u8_u3_n173 ) , .A( u1_u8_u3_n94 ) );
  OAI21_X1 u1_u8_u3_U91 (.ZN( u1_u8_u3_n111 ) , .B2( u1_u8_u3_n117 ) , .A( u1_u8_u3_n133 ) , .B1( u1_u8_u3_n176 ) );
  NAND4_X1 u1_u8_u3_U92 (.ZN( u1_out8_20 ) , .A4( u1_u8_u3_n122 ) , .A3( u1_u8_u3_n123 ) , .A1( u1_u8_u3_n175 ) , .A2( u1_u8_u3_n180 ) );
  INV_X1 u1_u8_u3_U93 (.A( u1_u8_u3_n126 ) , .ZN( u1_u8_u3_n180 ) );
  INV_X1 u1_u8_u3_U94 (.A( u1_u8_u3_n112 ) , .ZN( u1_u8_u3_n175 ) );
  NAND4_X1 u1_u8_u3_U95 (.ZN( u1_out8_1 ) , .A4( u1_u8_u3_n161 ) , .A3( u1_u8_u3_n162 ) , .A2( u1_u8_u3_n163 ) , .A1( u1_u8_u3_n185 ) );
  NAND2_X1 u1_u8_u3_U96 (.ZN( u1_u8_u3_n163 ) , .A2( u1_u8_u3_n170 ) , .A1( u1_u8_u3_n176 ) );
  AOI22_X1 u1_u8_u3_U97 (.B2( u1_u8_u3_n140 ) , .B1( u1_u8_u3_n141 ) , .A2( u1_u8_u3_n142 ) , .ZN( u1_u8_u3_n162 ) , .A1( u1_u8_u3_n177 ) );
  NAND3_X1 u1_u8_u3_U98 (.A1( u1_u8_u3_n114 ) , .ZN( u1_u8_u3_n115 ) , .A2( u1_u8_u3_n145 ) , .A3( u1_u8_u3_n153 ) );
  NAND3_X1 u1_u8_u3_U99 (.ZN( u1_u8_u3_n129 ) , .A2( u1_u8_u3_n144 ) , .A1( u1_u8_u3_n153 ) , .A3( u1_u8_u3_n182 ) );
  AOI22_X1 u1_u8_u6_U10 (.A2( u1_u8_u6_n151 ) , .B2( u1_u8_u6_n161 ) , .A1( u1_u8_u6_n167 ) , .B1( u1_u8_u6_n170 ) , .ZN( u1_u8_u6_n89 ) );
  AOI21_X1 u1_u8_u6_U11 (.B1( u1_u8_u6_n107 ) , .B2( u1_u8_u6_n132 ) , .A( u1_u8_u6_n158 ) , .ZN( u1_u8_u6_n88 ) );
  AOI21_X1 u1_u8_u6_U12 (.B2( u1_u8_u6_n147 ) , .B1( u1_u8_u6_n148 ) , .ZN( u1_u8_u6_n149 ) , .A( u1_u8_u6_n158 ) );
  AOI21_X1 u1_u8_u6_U13 (.ZN( u1_u8_u6_n106 ) , .A( u1_u8_u6_n142 ) , .B2( u1_u8_u6_n159 ) , .B1( u1_u8_u6_n164 ) );
  INV_X1 u1_u8_u6_U14 (.A( u1_u8_u6_n155 ) , .ZN( u1_u8_u6_n161 ) );
  INV_X1 u1_u8_u6_U15 (.A( u1_u8_u6_n128 ) , .ZN( u1_u8_u6_n164 ) );
  NAND2_X1 u1_u8_u6_U16 (.ZN( u1_u8_u6_n110 ) , .A1( u1_u8_u6_n122 ) , .A2( u1_u8_u6_n129 ) );
  NAND2_X1 u1_u8_u6_U17 (.ZN( u1_u8_u6_n124 ) , .A2( u1_u8_u6_n146 ) , .A1( u1_u8_u6_n148 ) );
  INV_X1 u1_u8_u6_U18 (.A( u1_u8_u6_n132 ) , .ZN( u1_u8_u6_n171 ) );
  AND2_X1 u1_u8_u6_U19 (.A1( u1_u8_u6_n100 ) , .ZN( u1_u8_u6_n130 ) , .A2( u1_u8_u6_n147 ) );
  INV_X1 u1_u8_u6_U20 (.A( u1_u8_u6_n127 ) , .ZN( u1_u8_u6_n173 ) );
  INV_X1 u1_u8_u6_U21 (.A( u1_u8_u6_n121 ) , .ZN( u1_u8_u6_n167 ) );
  INV_X1 u1_u8_u6_U22 (.A( u1_u8_u6_n100 ) , .ZN( u1_u8_u6_n169 ) );
  INV_X1 u1_u8_u6_U23 (.A( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n170 ) );
  INV_X1 u1_u8_u6_U24 (.A( u1_u8_u6_n113 ) , .ZN( u1_u8_u6_n168 ) );
  AND2_X1 u1_u8_u6_U25 (.A1( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n119 ) , .ZN( u1_u8_u6_n133 ) );
  AND2_X1 u1_u8_u6_U26 (.A2( u1_u8_u6_n121 ) , .A1( u1_u8_u6_n122 ) , .ZN( u1_u8_u6_n131 ) );
  AND3_X1 u1_u8_u6_U27 (.ZN( u1_u8_u6_n120 ) , .A2( u1_u8_u6_n127 ) , .A1( u1_u8_u6_n132 ) , .A3( u1_u8_u6_n145 ) );
  INV_X1 u1_u8_u6_U28 (.A( u1_u8_u6_n146 ) , .ZN( u1_u8_u6_n163 ) );
  AOI222_X1 u1_u8_u6_U29 (.ZN( u1_u8_u6_n114 ) , .A1( u1_u8_u6_n118 ) , .A2( u1_u8_u6_n126 ) , .B2( u1_u8_u6_n151 ) , .C2( u1_u8_u6_n159 ) , .C1( u1_u8_u6_n168 ) , .B1( u1_u8_u6_n169 ) );
  INV_X1 u1_u8_u6_U3 (.A( u1_u8_u6_n110 ) , .ZN( u1_u8_u6_n166 ) );
  NOR2_X1 u1_u8_u6_U30 (.A1( u1_u8_u6_n162 ) , .A2( u1_u8_u6_n165 ) , .ZN( u1_u8_u6_n98 ) );
  AOI211_X1 u1_u8_u6_U31 (.B( u1_u8_u6_n134 ) , .A( u1_u8_u6_n135 ) , .C1( u1_u8_u6_n136 ) , .ZN( u1_u8_u6_n137 ) , .C2( u1_u8_u6_n151 ) );
  AOI21_X1 u1_u8_u6_U32 (.B2( u1_u8_u6_n132 ) , .B1( u1_u8_u6_n133 ) , .ZN( u1_u8_u6_n134 ) , .A( u1_u8_u6_n158 ) );
  NAND4_X1 u1_u8_u6_U33 (.A4( u1_u8_u6_n127 ) , .A3( u1_u8_u6_n128 ) , .A2( u1_u8_u6_n129 ) , .A1( u1_u8_u6_n130 ) , .ZN( u1_u8_u6_n136 ) );
  AOI21_X1 u1_u8_u6_U34 (.B1( u1_u8_u6_n131 ) , .ZN( u1_u8_u6_n135 ) , .A( u1_u8_u6_n144 ) , .B2( u1_u8_u6_n146 ) );
  NAND2_X1 u1_u8_u6_U35 (.A1( u1_u8_u6_n144 ) , .ZN( u1_u8_u6_n151 ) , .A2( u1_u8_u6_n158 ) );
  NAND2_X1 u1_u8_u6_U36 (.ZN( u1_u8_u6_n132 ) , .A1( u1_u8_u6_n91 ) , .A2( u1_u8_u6_n97 ) );
  AOI22_X1 u1_u8_u6_U37 (.B2( u1_u8_u6_n110 ) , .B1( u1_u8_u6_n111 ) , .A1( u1_u8_u6_n112 ) , .ZN( u1_u8_u6_n115 ) , .A2( u1_u8_u6_n161 ) );
  NAND4_X1 u1_u8_u6_U38 (.A3( u1_u8_u6_n109 ) , .ZN( u1_u8_u6_n112 ) , .A4( u1_u8_u6_n132 ) , .A2( u1_u8_u6_n147 ) , .A1( u1_u8_u6_n166 ) );
  NOR2_X1 u1_u8_u6_U39 (.ZN( u1_u8_u6_n109 ) , .A1( u1_u8_u6_n170 ) , .A2( u1_u8_u6_n173 ) );
  INV_X1 u1_u8_u6_U4 (.A( u1_u8_u6_n142 ) , .ZN( u1_u8_u6_n174 ) );
  NOR2_X1 u1_u8_u6_U40 (.A2( u1_u8_u6_n126 ) , .ZN( u1_u8_u6_n155 ) , .A1( u1_u8_u6_n160 ) );
  NAND2_X1 u1_u8_u6_U41 (.ZN( u1_u8_u6_n146 ) , .A2( u1_u8_u6_n94 ) , .A1( u1_u8_u6_n99 ) );
  AOI21_X1 u1_u8_u6_U42 (.A( u1_u8_u6_n144 ) , .B2( u1_u8_u6_n145 ) , .B1( u1_u8_u6_n146 ) , .ZN( u1_u8_u6_n150 ) );
  INV_X1 u1_u8_u6_U43 (.A( u1_u8_u6_n111 ) , .ZN( u1_u8_u6_n158 ) );
  NAND2_X1 u1_u8_u6_U44 (.ZN( u1_u8_u6_n127 ) , .A1( u1_u8_u6_n91 ) , .A2( u1_u8_u6_n92 ) );
  NAND2_X1 u1_u8_u6_U45 (.ZN( u1_u8_u6_n129 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n96 ) );
  INV_X1 u1_u8_u6_U46 (.A( u1_u8_u6_n144 ) , .ZN( u1_u8_u6_n159 ) );
  NAND2_X1 u1_u8_u6_U47 (.ZN( u1_u8_u6_n145 ) , .A2( u1_u8_u6_n97 ) , .A1( u1_u8_u6_n98 ) );
  NAND2_X1 u1_u8_u6_U48 (.ZN( u1_u8_u6_n148 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n94 ) );
  NAND2_X1 u1_u8_u6_U49 (.ZN( u1_u8_u6_n108 ) , .A2( u1_u8_u6_n139 ) , .A1( u1_u8_u6_n144 ) );
  NAND2_X1 u1_u8_u6_U5 (.A2( u1_u8_u6_n143 ) , .ZN( u1_u8_u6_n152 ) , .A1( u1_u8_u6_n166 ) );
  NAND2_X1 u1_u8_u6_U50 (.ZN( u1_u8_u6_n121 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n97 ) );
  NAND2_X1 u1_u8_u6_U51 (.ZN( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n95 ) );
  AND2_X1 u1_u8_u6_U52 (.ZN( u1_u8_u6_n118 ) , .A2( u1_u8_u6_n91 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U53 (.ZN( u1_u8_u6_n147 ) , .A2( u1_u8_u6_n98 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U54 (.ZN( u1_u8_u6_n128 ) , .A1( u1_u8_u6_n94 ) , .A2( u1_u8_u6_n96 ) );
  NAND2_X1 u1_u8_u6_U55 (.ZN( u1_u8_u6_n119 ) , .A2( u1_u8_u6_n95 ) , .A1( u1_u8_u6_n99 ) );
  NAND2_X1 u1_u8_u6_U56 (.ZN( u1_u8_u6_n123 ) , .A2( u1_u8_u6_n91 ) , .A1( u1_u8_u6_n96 ) );
  NAND2_X1 u1_u8_u6_U57 (.ZN( u1_u8_u6_n100 ) , .A2( u1_u8_u6_n92 ) , .A1( u1_u8_u6_n98 ) );
  NAND2_X1 u1_u8_u6_U58 (.ZN( u1_u8_u6_n122 ) , .A1( u1_u8_u6_n94 ) , .A2( u1_u8_u6_n97 ) );
  INV_X1 u1_u8_u6_U59 (.A( u1_u8_u6_n139 ) , .ZN( u1_u8_u6_n160 ) );
  AOI22_X1 u1_u8_u6_U6 (.B2( u1_u8_u6_n101 ) , .A1( u1_u8_u6_n102 ) , .ZN( u1_u8_u6_n103 ) , .B1( u1_u8_u6_n160 ) , .A2( u1_u8_u6_n161 ) );
  NAND2_X1 u1_u8_u6_U60 (.ZN( u1_u8_u6_n113 ) , .A1( u1_u8_u6_n96 ) , .A2( u1_u8_u6_n98 ) );
  NOR2_X1 u1_u8_u6_U61 (.A2( u1_u8_X_40 ) , .A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n126 ) );
  NOR2_X1 u1_u8_u6_U62 (.A2( u1_u8_X_39 ) , .A1( u1_u8_X_42 ) , .ZN( u1_u8_u6_n92 ) );
  NOR2_X1 u1_u8_u6_U63 (.A2( u1_u8_X_39 ) , .A1( u1_u8_u6_n156 ) , .ZN( u1_u8_u6_n97 ) );
  NOR2_X1 u1_u8_u6_U64 (.A2( u1_u8_X_38 ) , .A1( u1_u8_u6_n165 ) , .ZN( u1_u8_u6_n95 ) );
  NOR2_X1 u1_u8_u6_U65 (.A2( u1_u8_X_41 ) , .ZN( u1_u8_u6_n111 ) , .A1( u1_u8_u6_n157 ) );
  NOR2_X1 u1_u8_u6_U66 (.A2( u1_u8_X_37 ) , .A1( u1_u8_u6_n162 ) , .ZN( u1_u8_u6_n94 ) );
  NOR2_X1 u1_u8_u6_U67 (.A2( u1_u8_X_37 ) , .A1( u1_u8_X_38 ) , .ZN( u1_u8_u6_n91 ) );
  NAND2_X1 u1_u8_u6_U68 (.A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n144 ) , .A2( u1_u8_u6_n157 ) );
  NAND2_X1 u1_u8_u6_U69 (.A2( u1_u8_X_40 ) , .A1( u1_u8_X_41 ) , .ZN( u1_u8_u6_n139 ) );
  NOR2_X1 u1_u8_u6_U7 (.A1( u1_u8_u6_n118 ) , .ZN( u1_u8_u6_n143 ) , .A2( u1_u8_u6_n168 ) );
  AND2_X1 u1_u8_u6_U70 (.A1( u1_u8_X_39 ) , .A2( u1_u8_u6_n156 ) , .ZN( u1_u8_u6_n96 ) );
  AND2_X1 u1_u8_u6_U71 (.A1( u1_u8_X_39 ) , .A2( u1_u8_X_42 ) , .ZN( u1_u8_u6_n99 ) );
  INV_X1 u1_u8_u6_U72 (.A( u1_u8_X_40 ) , .ZN( u1_u8_u6_n157 ) );
  INV_X1 u1_u8_u6_U73 (.A( u1_u8_X_37 ) , .ZN( u1_u8_u6_n165 ) );
  INV_X1 u1_u8_u6_U74 (.A( u1_u8_X_38 ) , .ZN( u1_u8_u6_n162 ) );
  INV_X1 u1_u8_u6_U75 (.A( u1_u8_X_42 ) , .ZN( u1_u8_u6_n156 ) );
  NAND4_X1 u1_u8_u6_U76 (.ZN( u1_out8_12 ) , .A4( u1_u8_u6_n114 ) , .A3( u1_u8_u6_n115 ) , .A2( u1_u8_u6_n116 ) , .A1( u1_u8_u6_n117 ) );
  OAI22_X1 u1_u8_u6_U77 (.B2( u1_u8_u6_n111 ) , .ZN( u1_u8_u6_n116 ) , .B1( u1_u8_u6_n126 ) , .A2( u1_u8_u6_n164 ) , .A1( u1_u8_u6_n167 ) );
  OAI21_X1 u1_u8_u6_U78 (.A( u1_u8_u6_n108 ) , .ZN( u1_u8_u6_n117 ) , .B2( u1_u8_u6_n141 ) , .B1( u1_u8_u6_n163 ) );
  NAND4_X1 u1_u8_u6_U79 (.ZN( u1_out8_32 ) , .A4( u1_u8_u6_n103 ) , .A3( u1_u8_u6_n104 ) , .A2( u1_u8_u6_n105 ) , .A1( u1_u8_u6_n106 ) );
  OAI21_X1 u1_u8_u6_U8 (.A( u1_u8_u6_n159 ) , .B1( u1_u8_u6_n169 ) , .B2( u1_u8_u6_n173 ) , .ZN( u1_u8_u6_n90 ) );
  AOI22_X1 u1_u8_u6_U80 (.ZN( u1_u8_u6_n105 ) , .A2( u1_u8_u6_n108 ) , .A1( u1_u8_u6_n118 ) , .B2( u1_u8_u6_n126 ) , .B1( u1_u8_u6_n171 ) );
  AOI22_X1 u1_u8_u6_U81 (.ZN( u1_u8_u6_n104 ) , .A1( u1_u8_u6_n111 ) , .B1( u1_u8_u6_n124 ) , .B2( u1_u8_u6_n151 ) , .A2( u1_u8_u6_n93 ) );
  OAI211_X1 u1_u8_u6_U82 (.ZN( u1_out8_7 ) , .B( u1_u8_u6_n153 ) , .C2( u1_u8_u6_n154 ) , .C1( u1_u8_u6_n155 ) , .A( u1_u8_u6_n174 ) );
  NOR3_X1 u1_u8_u6_U83 (.A1( u1_u8_u6_n141 ) , .ZN( u1_u8_u6_n154 ) , .A3( u1_u8_u6_n164 ) , .A2( u1_u8_u6_n171 ) );
  AOI211_X1 u1_u8_u6_U84 (.B( u1_u8_u6_n149 ) , .A( u1_u8_u6_n150 ) , .C2( u1_u8_u6_n151 ) , .C1( u1_u8_u6_n152 ) , .ZN( u1_u8_u6_n153 ) );
  OAI211_X1 u1_u8_u6_U85 (.ZN( u1_out8_22 ) , .B( u1_u8_u6_n137 ) , .A( u1_u8_u6_n138 ) , .C2( u1_u8_u6_n139 ) , .C1( u1_u8_u6_n140 ) );
  AOI22_X1 u1_u8_u6_U86 (.B1( u1_u8_u6_n124 ) , .A2( u1_u8_u6_n125 ) , .A1( u1_u8_u6_n126 ) , .ZN( u1_u8_u6_n138 ) , .B2( u1_u8_u6_n161 ) );
  AND4_X1 u1_u8_u6_U87 (.A3( u1_u8_u6_n119 ) , .A1( u1_u8_u6_n120 ) , .A4( u1_u8_u6_n129 ) , .ZN( u1_u8_u6_n140 ) , .A2( u1_u8_u6_n143 ) );
  NAND3_X1 u1_u8_u6_U88 (.A2( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n125 ) , .A1( u1_u8_u6_n130 ) , .A3( u1_u8_u6_n131 ) );
  NAND3_X1 u1_u8_u6_U89 (.A3( u1_u8_u6_n133 ) , .ZN( u1_u8_u6_n141 ) , .A1( u1_u8_u6_n145 ) , .A2( u1_u8_u6_n148 ) );
  INV_X1 u1_u8_u6_U9 (.ZN( u1_u8_u6_n172 ) , .A( u1_u8_u6_n88 ) );
  NAND3_X1 u1_u8_u6_U90 (.ZN( u1_u8_u6_n101 ) , .A3( u1_u8_u6_n107 ) , .A2( u1_u8_u6_n121 ) , .A1( u1_u8_u6_n127 ) );
  NAND3_X1 u1_u8_u6_U91 (.ZN( u1_u8_u6_n102 ) , .A3( u1_u8_u6_n130 ) , .A2( u1_u8_u6_n145 ) , .A1( u1_u8_u6_n166 ) );
  NAND3_X1 u1_u8_u6_U92 (.A3( u1_u8_u6_n113 ) , .A1( u1_u8_u6_n119 ) , .A2( u1_u8_u6_n123 ) , .ZN( u1_u8_u6_n93 ) );
  NAND3_X1 u1_u8_u6_U93 (.ZN( u1_u8_u6_n142 ) , .A2( u1_u8_u6_n172 ) , .A3( u1_u8_u6_n89 ) , .A1( u1_u8_u6_n90 ) );
  AND3_X1 u1_u8_u7_U10 (.A3( u1_u8_u7_n110 ) , .A2( u1_u8_u7_n127 ) , .A1( u1_u8_u7_n132 ) , .ZN( u1_u8_u7_n92 ) );
  OAI21_X1 u1_u8_u7_U11 (.A( u1_u8_u7_n161 ) , .B1( u1_u8_u7_n168 ) , .B2( u1_u8_u7_n173 ) , .ZN( u1_u8_u7_n91 ) );
  AOI211_X1 u1_u8_u7_U12 (.A( u1_u8_u7_n117 ) , .ZN( u1_u8_u7_n118 ) , .C2( u1_u8_u7_n126 ) , .C1( u1_u8_u7_n177 ) , .B( u1_u8_u7_n180 ) );
  OAI22_X1 u1_u8_u7_U13 (.B1( u1_u8_u7_n115 ) , .ZN( u1_u8_u7_n117 ) , .A2( u1_u8_u7_n133 ) , .A1( u1_u8_u7_n137 ) , .B2( u1_u8_u7_n162 ) );
  INV_X1 u1_u8_u7_U14 (.A( u1_u8_u7_n116 ) , .ZN( u1_u8_u7_n180 ) );
  NOR3_X1 u1_u8_u7_U15 (.ZN( u1_u8_u7_n115 ) , .A3( u1_u8_u7_n145 ) , .A2( u1_u8_u7_n168 ) , .A1( u1_u8_u7_n169 ) );
  OAI211_X1 u1_u8_u7_U16 (.B( u1_u8_u7_n122 ) , .A( u1_u8_u7_n123 ) , .C2( u1_u8_u7_n124 ) , .ZN( u1_u8_u7_n154 ) , .C1( u1_u8_u7_n162 ) );
  AOI222_X1 u1_u8_u7_U17 (.ZN( u1_u8_u7_n122 ) , .C2( u1_u8_u7_n126 ) , .C1( u1_u8_u7_n145 ) , .B1( u1_u8_u7_n161 ) , .A2( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n170 ) , .A1( u1_u8_u7_n176 ) );
  INV_X1 u1_u8_u7_U18 (.A( u1_u8_u7_n133 ) , .ZN( u1_u8_u7_n176 ) );
  NOR3_X1 u1_u8_u7_U19 (.A2( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n135 ) , .ZN( u1_u8_u7_n136 ) , .A3( u1_u8_u7_n171 ) );
  NOR2_X1 u1_u8_u7_U20 (.A1( u1_u8_u7_n130 ) , .A2( u1_u8_u7_n134 ) , .ZN( u1_u8_u7_n153 ) );
  INV_X1 u1_u8_u7_U21 (.A( u1_u8_u7_n101 ) , .ZN( u1_u8_u7_n165 ) );
  NOR2_X1 u1_u8_u7_U22 (.ZN( u1_u8_u7_n111 ) , .A2( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n169 ) );
  AOI21_X1 u1_u8_u7_U23 (.ZN( u1_u8_u7_n104 ) , .B2( u1_u8_u7_n112 ) , .B1( u1_u8_u7_n127 ) , .A( u1_u8_u7_n164 ) );
  AOI21_X1 u1_u8_u7_U24 (.ZN( u1_u8_u7_n106 ) , .B1( u1_u8_u7_n133 ) , .B2( u1_u8_u7_n146 ) , .A( u1_u8_u7_n162 ) );
  AOI21_X1 u1_u8_u7_U25 (.A( u1_u8_u7_n101 ) , .ZN( u1_u8_u7_n107 ) , .B2( u1_u8_u7_n128 ) , .B1( u1_u8_u7_n175 ) );
  INV_X1 u1_u8_u7_U26 (.A( u1_u8_u7_n138 ) , .ZN( u1_u8_u7_n171 ) );
  INV_X1 u1_u8_u7_U27 (.A( u1_u8_u7_n131 ) , .ZN( u1_u8_u7_n177 ) );
  INV_X1 u1_u8_u7_U28 (.A( u1_u8_u7_n110 ) , .ZN( u1_u8_u7_n174 ) );
  NAND2_X1 u1_u8_u7_U29 (.A1( u1_u8_u7_n129 ) , .A2( u1_u8_u7_n132 ) , .ZN( u1_u8_u7_n149 ) );
  OAI21_X1 u1_u8_u7_U3 (.ZN( u1_u8_u7_n159 ) , .A( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n171 ) , .B1( u1_u8_u7_n174 ) );
  NAND2_X1 u1_u8_u7_U30 (.A1( u1_u8_u7_n113 ) , .A2( u1_u8_u7_n124 ) , .ZN( u1_u8_u7_n130 ) );
  INV_X1 u1_u8_u7_U31 (.A( u1_u8_u7_n112 ) , .ZN( u1_u8_u7_n173 ) );
  INV_X1 u1_u8_u7_U32 (.A( u1_u8_u7_n128 ) , .ZN( u1_u8_u7_n168 ) );
  INV_X1 u1_u8_u7_U33 (.A( u1_u8_u7_n148 ) , .ZN( u1_u8_u7_n169 ) );
  INV_X1 u1_u8_u7_U34 (.A( u1_u8_u7_n127 ) , .ZN( u1_u8_u7_n179 ) );
  NOR2_X1 u1_u8_u7_U35 (.ZN( u1_u8_u7_n101 ) , .A2( u1_u8_u7_n150 ) , .A1( u1_u8_u7_n156 ) );
  AOI211_X1 u1_u8_u7_U36 (.B( u1_u8_u7_n154 ) , .A( u1_u8_u7_n155 ) , .C1( u1_u8_u7_n156 ) , .ZN( u1_u8_u7_n157 ) , .C2( u1_u8_u7_n172 ) );
  INV_X1 u1_u8_u7_U37 (.A( u1_u8_u7_n153 ) , .ZN( u1_u8_u7_n172 ) );
  AOI211_X1 u1_u8_u7_U38 (.B( u1_u8_u7_n139 ) , .A( u1_u8_u7_n140 ) , .C2( u1_u8_u7_n141 ) , .ZN( u1_u8_u7_n142 ) , .C1( u1_u8_u7_n156 ) );
  NAND4_X1 u1_u8_u7_U39 (.A3( u1_u8_u7_n127 ) , .A2( u1_u8_u7_n128 ) , .A1( u1_u8_u7_n129 ) , .ZN( u1_u8_u7_n141 ) , .A4( u1_u8_u7_n147 ) );
  INV_X1 u1_u8_u7_U4 (.A( u1_u8_u7_n111 ) , .ZN( u1_u8_u7_n170 ) );
  AOI21_X1 u1_u8_u7_U40 (.A( u1_u8_u7_n137 ) , .B1( u1_u8_u7_n138 ) , .ZN( u1_u8_u7_n139 ) , .B2( u1_u8_u7_n146 ) );
  OAI22_X1 u1_u8_u7_U41 (.B1( u1_u8_u7_n136 ) , .ZN( u1_u8_u7_n140 ) , .A1( u1_u8_u7_n153 ) , .B2( u1_u8_u7_n162 ) , .A2( u1_u8_u7_n164 ) );
  AOI21_X1 u1_u8_u7_U42 (.ZN( u1_u8_u7_n123 ) , .B1( u1_u8_u7_n165 ) , .B2( u1_u8_u7_n177 ) , .A( u1_u8_u7_n97 ) );
  AOI21_X1 u1_u8_u7_U43 (.B2( u1_u8_u7_n113 ) , .B1( u1_u8_u7_n124 ) , .A( u1_u8_u7_n125 ) , .ZN( u1_u8_u7_n97 ) );
  INV_X1 u1_u8_u7_U44 (.A( u1_u8_u7_n125 ) , .ZN( u1_u8_u7_n161 ) );
  INV_X1 u1_u8_u7_U45 (.A( u1_u8_u7_n152 ) , .ZN( u1_u8_u7_n162 ) );
  AOI22_X1 u1_u8_u7_U46 (.A2( u1_u8_u7_n114 ) , .ZN( u1_u8_u7_n119 ) , .B1( u1_u8_u7_n130 ) , .A1( u1_u8_u7_n156 ) , .B2( u1_u8_u7_n165 ) );
  NAND2_X1 u1_u8_u7_U47 (.A2( u1_u8_u7_n112 ) , .ZN( u1_u8_u7_n114 ) , .A1( u1_u8_u7_n175 ) );
  AND2_X1 u1_u8_u7_U48 (.ZN( u1_u8_u7_n145 ) , .A2( u1_u8_u7_n98 ) , .A1( u1_u8_u7_n99 ) );
  NOR2_X1 u1_u8_u7_U49 (.ZN( u1_u8_u7_n137 ) , .A1( u1_u8_u7_n150 ) , .A2( u1_u8_u7_n161 ) );
  INV_X1 u1_u8_u7_U5 (.A( u1_u8_u7_n149 ) , .ZN( u1_u8_u7_n175 ) );
  AOI21_X1 u1_u8_u7_U50 (.ZN( u1_u8_u7_n105 ) , .B2( u1_u8_u7_n110 ) , .A( u1_u8_u7_n125 ) , .B1( u1_u8_u7_n147 ) );
  NAND2_X1 u1_u8_u7_U51 (.ZN( u1_u8_u7_n146 ) , .A1( u1_u8_u7_n95 ) , .A2( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U52 (.A2( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n147 ) , .A1( u1_u8_u7_n93 ) );
  NAND2_X1 u1_u8_u7_U53 (.A1( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n127 ) , .A2( u1_u8_u7_n99 ) );
  OR2_X1 u1_u8_u7_U54 (.ZN( u1_u8_u7_n126 ) , .A2( u1_u8_u7_n152 ) , .A1( u1_u8_u7_n156 ) );
  NAND2_X1 u1_u8_u7_U55 (.A2( u1_u8_u7_n102 ) , .A1( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n133 ) );
  NAND2_X1 u1_u8_u7_U56 (.ZN( u1_u8_u7_n112 ) , .A2( u1_u8_u7_n96 ) , .A1( u1_u8_u7_n99 ) );
  NAND2_X1 u1_u8_u7_U57 (.A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n128 ) , .A1( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U58 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n113 ) , .A2( u1_u8_u7_n93 ) );
  NAND2_X1 u1_u8_u7_U59 (.A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n124 ) , .A1( u1_u8_u7_n96 ) );
  INV_X1 u1_u8_u7_U6 (.A( u1_u8_u7_n154 ) , .ZN( u1_u8_u7_n178 ) );
  NAND2_X1 u1_u8_u7_U60 (.ZN( u1_u8_u7_n110 ) , .A1( u1_u8_u7_n95 ) , .A2( u1_u8_u7_n96 ) );
  INV_X1 u1_u8_u7_U61 (.A( u1_u8_u7_n150 ) , .ZN( u1_u8_u7_n164 ) );
  AND2_X1 u1_u8_u7_U62 (.ZN( u1_u8_u7_n134 ) , .A1( u1_u8_u7_n93 ) , .A2( u1_u8_u7_n98 ) );
  NAND2_X1 u1_u8_u7_U63 (.A1( u1_u8_u7_n100 ) , .A2( u1_u8_u7_n102 ) , .ZN( u1_u8_u7_n129 ) );
  NAND2_X1 u1_u8_u7_U64 (.A2( u1_u8_u7_n103 ) , .ZN( u1_u8_u7_n131 ) , .A1( u1_u8_u7_n95 ) );
  NAND2_X1 u1_u8_u7_U65 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n138 ) , .A2( u1_u8_u7_n99 ) );
  NAND2_X1 u1_u8_u7_U66 (.ZN( u1_u8_u7_n132 ) , .A1( u1_u8_u7_n93 ) , .A2( u1_u8_u7_n96 ) );
  NAND2_X1 u1_u8_u7_U67 (.A1( u1_u8_u7_n100 ) , .ZN( u1_u8_u7_n148 ) , .A2( u1_u8_u7_n95 ) );
  NOR2_X1 u1_u8_u7_U68 (.A2( u1_u8_X_47 ) , .ZN( u1_u8_u7_n150 ) , .A1( u1_u8_u7_n163 ) );
  NOR2_X1 u1_u8_u7_U69 (.A2( u1_u8_X_43 ) , .A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n103 ) );
  AOI211_X1 u1_u8_u7_U7 (.ZN( u1_u8_u7_n116 ) , .A( u1_u8_u7_n155 ) , .C1( u1_u8_u7_n161 ) , .C2( u1_u8_u7_n171 ) , .B( u1_u8_u7_n94 ) );
  NOR2_X1 u1_u8_u7_U70 (.A2( u1_u8_X_48 ) , .A1( u1_u8_u7_n166 ) , .ZN( u1_u8_u7_n95 ) );
  NOR2_X1 u1_u8_u7_U71 (.A2( u1_u8_X_45 ) , .A1( u1_u8_X_48 ) , .ZN( u1_u8_u7_n99 ) );
  NOR2_X1 u1_u8_u7_U72 (.A2( u1_u8_X_44 ) , .A1( u1_u8_u7_n167 ) , .ZN( u1_u8_u7_n98 ) );
  NOR2_X1 u1_u8_u7_U73 (.A2( u1_u8_X_46 ) , .A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n152 ) );
  AND2_X1 u1_u8_u7_U74 (.A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n156 ) , .A2( u1_u8_u7_n163 ) );
  NAND2_X1 u1_u8_u7_U75 (.A2( u1_u8_X_46 ) , .A1( u1_u8_X_47 ) , .ZN( u1_u8_u7_n125 ) );
  AND2_X1 u1_u8_u7_U76 (.A2( u1_u8_X_45 ) , .A1( u1_u8_X_48 ) , .ZN( u1_u8_u7_n102 ) );
  AND2_X1 u1_u8_u7_U77 (.A2( u1_u8_X_43 ) , .A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n96 ) );
  AND2_X1 u1_u8_u7_U78 (.A1( u1_u8_X_44 ) , .ZN( u1_u8_u7_n100 ) , .A2( u1_u8_u7_n167 ) );
  AND2_X1 u1_u8_u7_U79 (.A1( u1_u8_X_48 ) , .A2( u1_u8_u7_n166 ) , .ZN( u1_u8_u7_n93 ) );
  OAI222_X1 u1_u8_u7_U8 (.C2( u1_u8_u7_n101 ) , .B2( u1_u8_u7_n111 ) , .A1( u1_u8_u7_n113 ) , .C1( u1_u8_u7_n146 ) , .A2( u1_u8_u7_n162 ) , .B1( u1_u8_u7_n164 ) , .ZN( u1_u8_u7_n94 ) );
  INV_X1 u1_u8_u7_U80 (.A( u1_u8_X_46 ) , .ZN( u1_u8_u7_n163 ) );
  INV_X1 u1_u8_u7_U81 (.A( u1_u8_X_43 ) , .ZN( u1_u8_u7_n167 ) );
  INV_X1 u1_u8_u7_U82 (.A( u1_u8_X_45 ) , .ZN( u1_u8_u7_n166 ) );
  NAND4_X1 u1_u8_u7_U83 (.ZN( u1_out8_5 ) , .A4( u1_u8_u7_n108 ) , .A3( u1_u8_u7_n109 ) , .A1( u1_u8_u7_n116 ) , .A2( u1_u8_u7_n123 ) );
  AOI22_X1 u1_u8_u7_U84 (.ZN( u1_u8_u7_n109 ) , .A2( u1_u8_u7_n126 ) , .B2( u1_u8_u7_n145 ) , .B1( u1_u8_u7_n156 ) , .A1( u1_u8_u7_n171 ) );
  NOR4_X1 u1_u8_u7_U85 (.A4( u1_u8_u7_n104 ) , .A3( u1_u8_u7_n105 ) , .A2( u1_u8_u7_n106 ) , .A1( u1_u8_u7_n107 ) , .ZN( u1_u8_u7_n108 ) );
  NAND4_X1 u1_u8_u7_U86 (.ZN( u1_out8_27 ) , .A4( u1_u8_u7_n118 ) , .A3( u1_u8_u7_n119 ) , .A2( u1_u8_u7_n120 ) , .A1( u1_u8_u7_n121 ) );
  OAI21_X1 u1_u8_u7_U87 (.ZN( u1_u8_u7_n121 ) , .B2( u1_u8_u7_n145 ) , .A( u1_u8_u7_n150 ) , .B1( u1_u8_u7_n174 ) );
  OAI21_X1 u1_u8_u7_U88 (.ZN( u1_u8_u7_n120 ) , .A( u1_u8_u7_n161 ) , .B2( u1_u8_u7_n170 ) , .B1( u1_u8_u7_n179 ) );
  NAND4_X1 u1_u8_u7_U89 (.ZN( u1_out8_21 ) , .A4( u1_u8_u7_n157 ) , .A3( u1_u8_u7_n158 ) , .A2( u1_u8_u7_n159 ) , .A1( u1_u8_u7_n160 ) );
  OAI221_X1 u1_u8_u7_U9 (.C1( u1_u8_u7_n101 ) , .C2( u1_u8_u7_n147 ) , .ZN( u1_u8_u7_n155 ) , .B2( u1_u8_u7_n162 ) , .A( u1_u8_u7_n91 ) , .B1( u1_u8_u7_n92 ) );
  OAI21_X1 u1_u8_u7_U90 (.B1( u1_u8_u7_n145 ) , .ZN( u1_u8_u7_n160 ) , .A( u1_u8_u7_n161 ) , .B2( u1_u8_u7_n177 ) );
  AOI22_X1 u1_u8_u7_U91 (.B2( u1_u8_u7_n149 ) , .B1( u1_u8_u7_n150 ) , .A2( u1_u8_u7_n151 ) , .A1( u1_u8_u7_n152 ) , .ZN( u1_u8_u7_n158 ) );
  NAND4_X1 u1_u8_u7_U92 (.ZN( u1_out8_15 ) , .A4( u1_u8_u7_n142 ) , .A3( u1_u8_u7_n143 ) , .A2( u1_u8_u7_n144 ) , .A1( u1_u8_u7_n178 ) );
  OR2_X1 u1_u8_u7_U93 (.A2( u1_u8_u7_n125 ) , .A1( u1_u8_u7_n129 ) , .ZN( u1_u8_u7_n144 ) );
  AOI22_X1 u1_u8_u7_U94 (.A2( u1_u8_u7_n126 ) , .ZN( u1_u8_u7_n143 ) , .B2( u1_u8_u7_n165 ) , .B1( u1_u8_u7_n173 ) , .A1( u1_u8_u7_n174 ) );
  NAND3_X1 u1_u8_u7_U95 (.A3( u1_u8_u7_n146 ) , .A2( u1_u8_u7_n147 ) , .A1( u1_u8_u7_n148 ) , .ZN( u1_u8_u7_n151 ) );
  NAND3_X1 u1_u8_u7_U96 (.A3( u1_u8_u7_n131 ) , .A2( u1_u8_u7_n132 ) , .A1( u1_u8_u7_n133 ) , .ZN( u1_u8_u7_n135 ) );
  XOR2_X1 u1_u9_U10 (.B( u1_K10_45 ) , .A( u1_R8_30 ) , .Z( u1_u9_X_45 ) );
  XOR2_X1 u1_u9_U11 (.B( u1_K10_44 ) , .A( u1_R8_29 ) , .Z( u1_u9_X_44 ) );
  XOR2_X1 u1_u9_U12 (.B( u1_K10_43 ) , .A( u1_R8_28 ) , .Z( u1_u9_X_43 ) );
  XOR2_X1 u1_u9_U13 (.B( u1_K10_42 ) , .A( u1_R8_29 ) , .Z( u1_u9_X_42 ) );
  XOR2_X1 u1_u9_U14 (.B( u1_K10_41 ) , .A( u1_R8_28 ) , .Z( u1_u9_X_41 ) );
  XOR2_X1 u1_u9_U16 (.B( u1_K10_3 ) , .A( u1_R8_2 ) , .Z( u1_u9_X_3 ) );
  XOR2_X1 u1_u9_U2 (.B( u1_K10_8 ) , .A( u1_R8_5 ) , .Z( u1_u9_X_8 ) );
  XOR2_X1 u1_u9_U24 (.B( u1_K10_32 ) , .A( u1_R8_21 ) , .Z( u1_u9_X_32 ) );
  XOR2_X1 u1_u9_U25 (.B( u1_K10_31 ) , .A( u1_R8_20 ) , .Z( u1_u9_X_31 ) );
  XOR2_X1 u1_u9_U26 (.B( u1_K10_30 ) , .A( u1_R8_21 ) , .Z( u1_u9_X_30 ) );
  XOR2_X1 u1_u9_U27 (.B( u1_K10_2 ) , .A( u1_R8_1 ) , .Z( u1_u9_X_2 ) );
  XOR2_X1 u1_u9_U28 (.B( u1_K10_29 ) , .A( u1_R8_20 ) , .Z( u1_u9_X_29 ) );
  XOR2_X1 u1_u9_U3 (.B( u1_K10_7 ) , .A( u1_R8_4 ) , .Z( u1_u9_X_7 ) );
  XOR2_X1 u1_u9_U31 (.B( u1_K10_26 ) , .A( u1_R8_17 ) , .Z( u1_u9_X_26 ) );
  XOR2_X1 u1_u9_U32 (.B( u1_K10_25 ) , .A( u1_R8_16 ) , .Z( u1_u9_X_25 ) );
  XOR2_X1 u1_u9_U33 (.B( u1_K10_24 ) , .A( u1_R8_17 ) , .Z( u1_u9_X_24 ) );
  XOR2_X1 u1_u9_U34 (.B( u1_K10_23 ) , .A( u1_R8_16 ) , .Z( u1_u9_X_23 ) );
  XOR2_X1 u1_u9_U38 (.B( u1_K10_1 ) , .A( u1_R8_32 ) , .Z( u1_u9_X_1 ) );
  XOR2_X1 u1_u9_U4 (.B( u1_K10_6 ) , .A( u1_R8_5 ) , .Z( u1_u9_X_6 ) );
  XOR2_X1 u1_u9_U5 (.B( u1_K10_5 ) , .A( u1_R8_4 ) , .Z( u1_u9_X_5 ) );
  XOR2_X1 u1_u9_U6 (.B( u1_K10_4 ) , .A( u1_R8_3 ) , .Z( u1_u9_X_4 ) );
  XOR2_X1 u1_u9_U7 (.B( u1_K10_48 ) , .A( u1_R8_1 ) , .Z( u1_u9_X_48 ) );
  XOR2_X1 u1_u9_U8 (.B( u1_K10_47 ) , .A( u1_R8_32 ) , .Z( u1_u9_X_47 ) );
  XOR2_X1 u1_u9_U9 (.B( u1_K10_46 ) , .A( u1_R8_31 ) , .Z( u1_u9_X_46 ) );
  AND3_X1 u1_u9_u0_U10 (.A2( u1_u9_u0_n112 ) , .ZN( u1_u9_u0_n127 ) , .A3( u1_u9_u0_n130 ) , .A1( u1_u9_u0_n148 ) );
  NAND2_X1 u1_u9_u0_U11 (.ZN( u1_u9_u0_n113 ) , .A1( u1_u9_u0_n139 ) , .A2( u1_u9_u0_n149 ) );
  AND2_X1 u1_u9_u0_U12 (.ZN( u1_u9_u0_n107 ) , .A1( u1_u9_u0_n130 ) , .A2( u1_u9_u0_n140 ) );
  AND2_X1 u1_u9_u0_U13 (.A2( u1_u9_u0_n129 ) , .A1( u1_u9_u0_n130 ) , .ZN( u1_u9_u0_n151 ) );
  AND2_X1 u1_u9_u0_U14 (.A1( u1_u9_u0_n108 ) , .A2( u1_u9_u0_n125 ) , .ZN( u1_u9_u0_n145 ) );
  INV_X1 u1_u9_u0_U15 (.A( u1_u9_u0_n143 ) , .ZN( u1_u9_u0_n173 ) );
  NOR2_X1 u1_u9_u0_U16 (.A2( u1_u9_u0_n136 ) , .ZN( u1_u9_u0_n147 ) , .A1( u1_u9_u0_n160 ) );
  AOI21_X1 u1_u9_u0_U17 (.B1( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n132 ) , .A( u1_u9_u0_n165 ) , .B2( u1_u9_u0_n93 ) );
  INV_X1 u1_u9_u0_U18 (.A( u1_u9_u0_n142 ) , .ZN( u1_u9_u0_n165 ) );
  OAI221_X1 u1_u9_u0_U19 (.C1( u1_u9_u0_n121 ) , .ZN( u1_u9_u0_n122 ) , .B2( u1_u9_u0_n127 ) , .A( u1_u9_u0_n143 ) , .B1( u1_u9_u0_n144 ) , .C2( u1_u9_u0_n147 ) );
  OAI22_X1 u1_u9_u0_U20 (.B1( u1_u9_u0_n131 ) , .A1( u1_u9_u0_n144 ) , .B2( u1_u9_u0_n147 ) , .A2( u1_u9_u0_n90 ) , .ZN( u1_u9_u0_n91 ) );
  AND3_X1 u1_u9_u0_U21 (.A3( u1_u9_u0_n121 ) , .A2( u1_u9_u0_n125 ) , .A1( u1_u9_u0_n148 ) , .ZN( u1_u9_u0_n90 ) );
  OAI22_X1 u1_u9_u0_U22 (.B1( u1_u9_u0_n125 ) , .ZN( u1_u9_u0_n126 ) , .A1( u1_u9_u0_n138 ) , .A2( u1_u9_u0_n146 ) , .B2( u1_u9_u0_n147 ) );
  NOR2_X1 u1_u9_u0_U23 (.A1( u1_u9_u0_n163 ) , .A2( u1_u9_u0_n164 ) , .ZN( u1_u9_u0_n95 ) );
  INV_X1 u1_u9_u0_U24 (.A( u1_u9_u0_n136 ) , .ZN( u1_u9_u0_n161 ) );
  NOR2_X1 u1_u9_u0_U25 (.A1( u1_u9_u0_n120 ) , .ZN( u1_u9_u0_n143 ) , .A2( u1_u9_u0_n167 ) );
  OAI221_X1 u1_u9_u0_U26 (.C1( u1_u9_u0_n112 ) , .ZN( u1_u9_u0_n120 ) , .B1( u1_u9_u0_n138 ) , .B2( u1_u9_u0_n141 ) , .C2( u1_u9_u0_n147 ) , .A( u1_u9_u0_n172 ) );
  AOI211_X1 u1_u9_u0_U27 (.B( u1_u9_u0_n115 ) , .A( u1_u9_u0_n116 ) , .C2( u1_u9_u0_n117 ) , .C1( u1_u9_u0_n118 ) , .ZN( u1_u9_u0_n119 ) );
  NAND2_X1 u1_u9_u0_U28 (.A1( u1_u9_u0_n101 ) , .A2( u1_u9_u0_n102 ) , .ZN( u1_u9_u0_n150 ) );
  AOI22_X1 u1_u9_u0_U29 (.B2( u1_u9_u0_n109 ) , .A2( u1_u9_u0_n110 ) , .ZN( u1_u9_u0_n111 ) , .B1( u1_u9_u0_n118 ) , .A1( u1_u9_u0_n160 ) );
  INV_X1 u1_u9_u0_U3 (.A( u1_u9_u0_n113 ) , .ZN( u1_u9_u0_n166 ) );
  INV_X1 u1_u9_u0_U30 (.A( u1_u9_u0_n118 ) , .ZN( u1_u9_u0_n158 ) );
  NAND2_X1 u1_u9_u0_U31 (.A2( u1_u9_u0_n100 ) , .A1( u1_u9_u0_n101 ) , .ZN( u1_u9_u0_n139 ) );
  NAND2_X1 u1_u9_u0_U32 (.A2( u1_u9_u0_n100 ) , .ZN( u1_u9_u0_n131 ) , .A1( u1_u9_u0_n92 ) );
  NAND2_X1 u1_u9_u0_U33 (.ZN( u1_u9_u0_n108 ) , .A1( u1_u9_u0_n92 ) , .A2( u1_u9_u0_n94 ) );
  AOI21_X1 u1_u9_u0_U34 (.ZN( u1_u9_u0_n104 ) , .B1( u1_u9_u0_n107 ) , .B2( u1_u9_u0_n141 ) , .A( u1_u9_u0_n144 ) );
  AOI21_X1 u1_u9_u0_U35 (.B1( u1_u9_u0_n127 ) , .B2( u1_u9_u0_n129 ) , .A( u1_u9_u0_n138 ) , .ZN( u1_u9_u0_n96 ) );
  NAND2_X1 u1_u9_u0_U36 (.A2( u1_u9_u0_n102 ) , .ZN( u1_u9_u0_n114 ) , .A1( u1_u9_u0_n92 ) );
  AOI21_X1 u1_u9_u0_U37 (.ZN( u1_u9_u0_n116 ) , .B2( u1_u9_u0_n142 ) , .A( u1_u9_u0_n144 ) , .B1( u1_u9_u0_n166 ) );
  NAND2_X1 u1_u9_u0_U38 (.A1( u1_u9_u0_n101 ) , .ZN( u1_u9_u0_n130 ) , .A2( u1_u9_u0_n94 ) );
  NAND2_X1 u1_u9_u0_U39 (.A1( u1_u9_u0_n100 ) , .A2( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n125 ) );
  AOI21_X1 u1_u9_u0_U4 (.B1( u1_u9_u0_n114 ) , .ZN( u1_u9_u0_n115 ) , .B2( u1_u9_u0_n129 ) , .A( u1_u9_u0_n161 ) );
  NAND2_X1 u1_u9_u0_U40 (.A2( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n140 ) , .A1( u1_u9_u0_n94 ) );
  INV_X1 u1_u9_u0_U41 (.A( u1_u9_u0_n138 ) , .ZN( u1_u9_u0_n160 ) );
  NAND2_X1 u1_u9_u0_U42 (.A2( u1_u9_u0_n102 ) , .A1( u1_u9_u0_n103 ) , .ZN( u1_u9_u0_n149 ) );
  NAND2_X1 u1_u9_u0_U43 (.A2( u1_u9_u0_n101 ) , .ZN( u1_u9_u0_n121 ) , .A1( u1_u9_u0_n93 ) );
  NAND2_X1 u1_u9_u0_U44 (.ZN( u1_u9_u0_n112 ) , .A2( u1_u9_u0_n92 ) , .A1( u1_u9_u0_n93 ) );
  INV_X1 u1_u9_u0_U45 (.ZN( u1_u9_u0_n172 ) , .A( u1_u9_u0_n88 ) );
  OAI222_X1 u1_u9_u0_U46 (.C1( u1_u9_u0_n108 ) , .A1( u1_u9_u0_n125 ) , .B2( u1_u9_u0_n128 ) , .B1( u1_u9_u0_n144 ) , .A2( u1_u9_u0_n158 ) , .C2( u1_u9_u0_n161 ) , .ZN( u1_u9_u0_n88 ) );
  OR3_X1 u1_u9_u0_U47 (.A3( u1_u9_u0_n152 ) , .A2( u1_u9_u0_n153 ) , .A1( u1_u9_u0_n154 ) , .ZN( u1_u9_u0_n155 ) );
  AOI21_X1 u1_u9_u0_U48 (.A( u1_u9_u0_n144 ) , .B2( u1_u9_u0_n145 ) , .B1( u1_u9_u0_n146 ) , .ZN( u1_u9_u0_n154 ) );
  AOI21_X1 u1_u9_u0_U49 (.B2( u1_u9_u0_n150 ) , .B1( u1_u9_u0_n151 ) , .ZN( u1_u9_u0_n152 ) , .A( u1_u9_u0_n158 ) );
  AOI21_X1 u1_u9_u0_U5 (.B2( u1_u9_u0_n131 ) , .ZN( u1_u9_u0_n134 ) , .B1( u1_u9_u0_n151 ) , .A( u1_u9_u0_n158 ) );
  AOI21_X1 u1_u9_u0_U50 (.A( u1_u9_u0_n147 ) , .B2( u1_u9_u0_n148 ) , .B1( u1_u9_u0_n149 ) , .ZN( u1_u9_u0_n153 ) );
  INV_X1 u1_u9_u0_U51 (.ZN( u1_u9_u0_n171 ) , .A( u1_u9_u0_n99 ) );
  OAI211_X1 u1_u9_u0_U52 (.C2( u1_u9_u0_n140 ) , .C1( u1_u9_u0_n161 ) , .A( u1_u9_u0_n169 ) , .B( u1_u9_u0_n98 ) , .ZN( u1_u9_u0_n99 ) );
  INV_X1 u1_u9_u0_U53 (.ZN( u1_u9_u0_n169 ) , .A( u1_u9_u0_n91 ) );
  AOI211_X1 u1_u9_u0_U54 (.C1( u1_u9_u0_n118 ) , .A( u1_u9_u0_n123 ) , .B( u1_u9_u0_n96 ) , .C2( u1_u9_u0_n97 ) , .ZN( u1_u9_u0_n98 ) );
  NOR2_X1 u1_u9_u0_U55 (.A2( u1_u9_X_2 ) , .ZN( u1_u9_u0_n103 ) , .A1( u1_u9_u0_n164 ) );
  NOR2_X1 u1_u9_u0_U56 (.A2( u1_u9_X_4 ) , .A1( u1_u9_X_5 ) , .ZN( u1_u9_u0_n118 ) );
  NOR2_X1 u1_u9_u0_U57 (.A2( u1_u9_X_3 ) , .A1( u1_u9_X_6 ) , .ZN( u1_u9_u0_n94 ) );
  NOR2_X1 u1_u9_u0_U58 (.A2( u1_u9_X_6 ) , .ZN( u1_u9_u0_n100 ) , .A1( u1_u9_u0_n162 ) );
  NAND2_X1 u1_u9_u0_U59 (.A2( u1_u9_X_4 ) , .A1( u1_u9_X_5 ) , .ZN( u1_u9_u0_n144 ) );
  NOR2_X1 u1_u9_u0_U6 (.A1( u1_u9_u0_n108 ) , .ZN( u1_u9_u0_n123 ) , .A2( u1_u9_u0_n158 ) );
  NOR2_X1 u1_u9_u0_U60 (.A2( u1_u9_X_5 ) , .ZN( u1_u9_u0_n136 ) , .A1( u1_u9_u0_n159 ) );
  NAND2_X1 u1_u9_u0_U61 (.A1( u1_u9_X_5 ) , .ZN( u1_u9_u0_n138 ) , .A2( u1_u9_u0_n159 ) );
  AND2_X1 u1_u9_u0_U62 (.A2( u1_u9_X_3 ) , .A1( u1_u9_X_6 ) , .ZN( u1_u9_u0_n102 ) );
  AND2_X1 u1_u9_u0_U63 (.A1( u1_u9_X_6 ) , .A2( u1_u9_u0_n162 ) , .ZN( u1_u9_u0_n93 ) );
  INV_X1 u1_u9_u0_U64 (.A( u1_u9_X_4 ) , .ZN( u1_u9_u0_n159 ) );
  INV_X1 u1_u9_u0_U65 (.A( u1_u9_X_3 ) , .ZN( u1_u9_u0_n162 ) );
  INV_X1 u1_u9_u0_U66 (.A( u1_u9_X_2 ) , .ZN( u1_u9_u0_n163 ) );
  INV_X1 u1_u9_u0_U67 (.A( u1_u9_u0_n126 ) , .ZN( u1_u9_u0_n168 ) );
  AOI211_X1 u1_u9_u0_U68 (.B( u1_u9_u0_n133 ) , .A( u1_u9_u0_n134 ) , .C2( u1_u9_u0_n135 ) , .C1( u1_u9_u0_n136 ) , .ZN( u1_u9_u0_n137 ) );
  INV_X1 u1_u9_u0_U69 (.ZN( u1_u9_u0_n174 ) , .A( u1_u9_u0_n89 ) );
  OAI21_X1 u1_u9_u0_U7 (.B1( u1_u9_u0_n150 ) , .B2( u1_u9_u0_n158 ) , .A( u1_u9_u0_n172 ) , .ZN( u1_u9_u0_n89 ) );
  AOI211_X1 u1_u9_u0_U70 (.B( u1_u9_u0_n104 ) , .A( u1_u9_u0_n105 ) , .ZN( u1_u9_u0_n106 ) , .C2( u1_u9_u0_n113 ) , .C1( u1_u9_u0_n160 ) );
  OR4_X1 u1_u9_u0_U71 (.ZN( u1_out9_17 ) , .A4( u1_u9_u0_n122 ) , .A2( u1_u9_u0_n123 ) , .A1( u1_u9_u0_n124 ) , .A3( u1_u9_u0_n170 ) );
  AOI21_X1 u1_u9_u0_U72 (.B2( u1_u9_u0_n107 ) , .ZN( u1_u9_u0_n124 ) , .B1( u1_u9_u0_n128 ) , .A( u1_u9_u0_n161 ) );
  INV_X1 u1_u9_u0_U73 (.A( u1_u9_u0_n111 ) , .ZN( u1_u9_u0_n170 ) );
  OR4_X1 u1_u9_u0_U74 (.ZN( u1_out9_31 ) , .A4( u1_u9_u0_n155 ) , .A2( u1_u9_u0_n156 ) , .A1( u1_u9_u0_n157 ) , .A3( u1_u9_u0_n173 ) );
  AOI21_X1 u1_u9_u0_U75 (.A( u1_u9_u0_n138 ) , .B2( u1_u9_u0_n139 ) , .B1( u1_u9_u0_n140 ) , .ZN( u1_u9_u0_n157 ) );
  AOI21_X1 u1_u9_u0_U76 (.B2( u1_u9_u0_n141 ) , .B1( u1_u9_u0_n142 ) , .ZN( u1_u9_u0_n156 ) , .A( u1_u9_u0_n161 ) );
  AOI21_X1 u1_u9_u0_U77 (.B1( u1_u9_u0_n132 ) , .ZN( u1_u9_u0_n133 ) , .A( u1_u9_u0_n144 ) , .B2( u1_u9_u0_n166 ) );
  OAI22_X1 u1_u9_u0_U78 (.ZN( u1_u9_u0_n105 ) , .A2( u1_u9_u0_n132 ) , .B1( u1_u9_u0_n146 ) , .A1( u1_u9_u0_n147 ) , .B2( u1_u9_u0_n161 ) );
  NAND2_X1 u1_u9_u0_U79 (.ZN( u1_u9_u0_n110 ) , .A2( u1_u9_u0_n132 ) , .A1( u1_u9_u0_n145 ) );
  AND2_X1 u1_u9_u0_U8 (.A1( u1_u9_u0_n114 ) , .A2( u1_u9_u0_n121 ) , .ZN( u1_u9_u0_n146 ) );
  INV_X1 u1_u9_u0_U80 (.A( u1_u9_u0_n119 ) , .ZN( u1_u9_u0_n167 ) );
  NAND2_X1 u1_u9_u0_U81 (.ZN( u1_u9_u0_n148 ) , .A1( u1_u9_u0_n93 ) , .A2( u1_u9_u0_n95 ) );
  NAND2_X1 u1_u9_u0_U82 (.A1( u1_u9_u0_n100 ) , .ZN( u1_u9_u0_n129 ) , .A2( u1_u9_u0_n95 ) );
  NAND2_X1 u1_u9_u0_U83 (.A1( u1_u9_u0_n102 ) , .ZN( u1_u9_u0_n128 ) , .A2( u1_u9_u0_n95 ) );
  NOR2_X1 u1_u9_u0_U84 (.A2( u1_u9_X_1 ) , .A1( u1_u9_X_2 ) , .ZN( u1_u9_u0_n92 ) );
  NAND2_X1 u1_u9_u0_U85 (.ZN( u1_u9_u0_n142 ) , .A1( u1_u9_u0_n94 ) , .A2( u1_u9_u0_n95 ) );
  NOR2_X1 u1_u9_u0_U86 (.A2( u1_u9_X_1 ) , .ZN( u1_u9_u0_n101 ) , .A1( u1_u9_u0_n163 ) );
  INV_X1 u1_u9_u0_U87 (.A( u1_u9_X_1 ) , .ZN( u1_u9_u0_n164 ) );
  NAND3_X1 u1_u9_u0_U88 (.ZN( u1_out9_23 ) , .A3( u1_u9_u0_n137 ) , .A1( u1_u9_u0_n168 ) , .A2( u1_u9_u0_n171 ) );
  NAND3_X1 u1_u9_u0_U89 (.A3( u1_u9_u0_n127 ) , .A2( u1_u9_u0_n128 ) , .ZN( u1_u9_u0_n135 ) , .A1( u1_u9_u0_n150 ) );
  AND2_X1 u1_u9_u0_U9 (.A1( u1_u9_u0_n131 ) , .ZN( u1_u9_u0_n141 ) , .A2( u1_u9_u0_n150 ) );
  NAND3_X1 u1_u9_u0_U90 (.ZN( u1_u9_u0_n117 ) , .A3( u1_u9_u0_n132 ) , .A2( u1_u9_u0_n139 ) , .A1( u1_u9_u0_n148 ) );
  NAND3_X1 u1_u9_u0_U91 (.ZN( u1_u9_u0_n109 ) , .A2( u1_u9_u0_n114 ) , .A3( u1_u9_u0_n140 ) , .A1( u1_u9_u0_n149 ) );
  NAND3_X1 u1_u9_u0_U92 (.ZN( u1_out9_9 ) , .A3( u1_u9_u0_n106 ) , .A2( u1_u9_u0_n171 ) , .A1( u1_u9_u0_n174 ) );
  NAND3_X1 u1_u9_u0_U93 (.A2( u1_u9_u0_n128 ) , .A1( u1_u9_u0_n132 ) , .A3( u1_u9_u0_n146 ) , .ZN( u1_u9_u0_n97 ) );
  AND3_X1 u1_u9_u7_U10 (.A3( u1_u9_u7_n110 ) , .A2( u1_u9_u7_n127 ) , .A1( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U11 (.A( u1_u9_u7_n161 ) , .B1( u1_u9_u7_n168 ) , .B2( u1_u9_u7_n173 ) , .ZN( u1_u9_u7_n91 ) );
  AOI211_X1 u1_u9_u7_U12 (.A( u1_u9_u7_n117 ) , .ZN( u1_u9_u7_n118 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n177 ) , .B( u1_u9_u7_n180 ) );
  OAI22_X1 u1_u9_u7_U13 (.B1( u1_u9_u7_n115 ) , .ZN( u1_u9_u7_n117 ) , .A2( u1_u9_u7_n133 ) , .A1( u1_u9_u7_n137 ) , .B2( u1_u9_u7_n162 ) );
  INV_X1 u1_u9_u7_U14 (.A( u1_u9_u7_n116 ) , .ZN( u1_u9_u7_n180 ) );
  NOR3_X1 u1_u9_u7_U15 (.ZN( u1_u9_u7_n115 ) , .A3( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n168 ) , .A1( u1_u9_u7_n169 ) );
  OAI211_X1 u1_u9_u7_U16 (.B( u1_u9_u7_n122 ) , .A( u1_u9_u7_n123 ) , .C2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n154 ) , .C1( u1_u9_u7_n162 ) );
  AOI222_X1 u1_u9_u7_U17 (.ZN( u1_u9_u7_n122 ) , .C2( u1_u9_u7_n126 ) , .C1( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n161 ) , .A2( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n170 ) , .A1( u1_u9_u7_n176 ) );
  INV_X1 u1_u9_u7_U18 (.A( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n176 ) );
  NOR3_X1 u1_u9_u7_U19 (.A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n135 ) , .ZN( u1_u9_u7_n136 ) , .A3( u1_u9_u7_n171 ) );
  NOR2_X1 u1_u9_u7_U20 (.A1( u1_u9_u7_n130 ) , .A2( u1_u9_u7_n134 ) , .ZN( u1_u9_u7_n153 ) );
  INV_X1 u1_u9_u7_U21 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n165 ) );
  NOR2_X1 u1_u9_u7_U22 (.ZN( u1_u9_u7_n111 ) , .A2( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n169 ) );
  AOI21_X1 u1_u9_u7_U23 (.ZN( u1_u9_u7_n104 ) , .B2( u1_u9_u7_n112 ) , .B1( u1_u9_u7_n127 ) , .A( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U24 (.ZN( u1_u9_u7_n106 ) , .B1( u1_u9_u7_n133 ) , .B2( u1_u9_u7_n146 ) , .A( u1_u9_u7_n162 ) );
  AOI21_X1 u1_u9_u7_U25 (.A( u1_u9_u7_n101 ) , .ZN( u1_u9_u7_n107 ) , .B2( u1_u9_u7_n128 ) , .B1( u1_u9_u7_n175 ) );
  INV_X1 u1_u9_u7_U26 (.A( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n171 ) );
  INV_X1 u1_u9_u7_U27 (.A( u1_u9_u7_n131 ) , .ZN( u1_u9_u7_n177 ) );
  INV_X1 u1_u9_u7_U28 (.A( u1_u9_u7_n110 ) , .ZN( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U29 (.A1( u1_u9_u7_n129 ) , .A2( u1_u9_u7_n132 ) , .ZN( u1_u9_u7_n149 ) );
  OAI21_X1 u1_u9_u7_U3 (.ZN( u1_u9_u7_n159 ) , .A( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n171 ) , .B1( u1_u9_u7_n174 ) );
  NAND2_X1 u1_u9_u7_U30 (.A1( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n124 ) , .ZN( u1_u9_u7_n130 ) );
  INV_X1 u1_u9_u7_U31 (.A( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n173 ) );
  INV_X1 u1_u9_u7_U32 (.A( u1_u9_u7_n128 ) , .ZN( u1_u9_u7_n168 ) );
  INV_X1 u1_u9_u7_U33 (.A( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n169 ) );
  INV_X1 u1_u9_u7_U34 (.A( u1_u9_u7_n127 ) , .ZN( u1_u9_u7_n179 ) );
  NOR2_X1 u1_u9_u7_U35 (.ZN( u1_u9_u7_n101 ) , .A2( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n156 ) );
  AOI211_X1 u1_u9_u7_U36 (.B( u1_u9_u7_n154 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n156 ) , .ZN( u1_u9_u7_n157 ) , .C2( u1_u9_u7_n172 ) );
  INV_X1 u1_u9_u7_U37 (.A( u1_u9_u7_n153 ) , .ZN( u1_u9_u7_n172 ) );
  AOI211_X1 u1_u9_u7_U38 (.B( u1_u9_u7_n139 ) , .A( u1_u9_u7_n140 ) , .C2( u1_u9_u7_n141 ) , .ZN( u1_u9_u7_n142 ) , .C1( u1_u9_u7_n156 ) );
  NAND4_X1 u1_u9_u7_U39 (.A3( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n141 ) , .A4( u1_u9_u7_n147 ) );
  INV_X1 u1_u9_u7_U4 (.A( u1_u9_u7_n111 ) , .ZN( u1_u9_u7_n170 ) );
  AOI21_X1 u1_u9_u7_U40 (.A( u1_u9_u7_n137 ) , .B1( u1_u9_u7_n138 ) , .ZN( u1_u9_u7_n139 ) , .B2( u1_u9_u7_n146 ) );
  OAI22_X1 u1_u9_u7_U41 (.B1( u1_u9_u7_n136 ) , .ZN( u1_u9_u7_n140 ) , .A1( u1_u9_u7_n153 ) , .B2( u1_u9_u7_n162 ) , .A2( u1_u9_u7_n164 ) );
  AOI21_X1 u1_u9_u7_U42 (.ZN( u1_u9_u7_n123 ) , .B1( u1_u9_u7_n165 ) , .B2( u1_u9_u7_n177 ) , .A( u1_u9_u7_n97 ) );
  AOI21_X1 u1_u9_u7_U43 (.B2( u1_u9_u7_n113 ) , .B1( u1_u9_u7_n124 ) , .A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n97 ) );
  INV_X1 u1_u9_u7_U44 (.A( u1_u9_u7_n125 ) , .ZN( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U45 (.A( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n162 ) );
  AOI22_X1 u1_u9_u7_U46 (.A2( u1_u9_u7_n114 ) , .ZN( u1_u9_u7_n119 ) , .B1( u1_u9_u7_n130 ) , .A1( u1_u9_u7_n156 ) , .B2( u1_u9_u7_n165 ) );
  NAND2_X1 u1_u9_u7_U47 (.A2( u1_u9_u7_n112 ) , .ZN( u1_u9_u7_n114 ) , .A1( u1_u9_u7_n175 ) );
  AND2_X1 u1_u9_u7_U48 (.ZN( u1_u9_u7_n145 ) , .A2( u1_u9_u7_n98 ) , .A1( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U49 (.ZN( u1_u9_u7_n137 ) , .A1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n161 ) );
  INV_X1 u1_u9_u7_U5 (.A( u1_u9_u7_n149 ) , .ZN( u1_u9_u7_n175 ) );
  AOI21_X1 u1_u9_u7_U50 (.ZN( u1_u9_u7_n105 ) , .B2( u1_u9_u7_n110 ) , .A( u1_u9_u7_n125 ) , .B1( u1_u9_u7_n147 ) );
  NAND2_X1 u1_u9_u7_U51 (.ZN( u1_u9_u7_n146 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U52 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U53 (.A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n127 ) , .A2( u1_u9_u7_n99 ) );
  OR2_X1 u1_u9_u7_U54 (.ZN( u1_u9_u7_n126 ) , .A2( u1_u9_u7_n152 ) , .A1( u1_u9_u7_n156 ) );
  NAND2_X1 u1_u9_u7_U55 (.A2( u1_u9_u7_n102 ) , .A1( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n133 ) );
  NAND2_X1 u1_u9_u7_U56 (.ZN( u1_u9_u7_n112 ) , .A2( u1_u9_u7_n96 ) , .A1( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U57 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n128 ) , .A1( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U58 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n113 ) , .A2( u1_u9_u7_n93 ) );
  NAND2_X1 u1_u9_u7_U59 (.A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n124 ) , .A1( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U6 (.A( u1_u9_u7_n154 ) , .ZN( u1_u9_u7_n178 ) );
  NAND2_X1 u1_u9_u7_U60 (.ZN( u1_u9_u7_n110 ) , .A1( u1_u9_u7_n95 ) , .A2( u1_u9_u7_n96 ) );
  INV_X1 u1_u9_u7_U61 (.A( u1_u9_u7_n150 ) , .ZN( u1_u9_u7_n164 ) );
  AND2_X1 u1_u9_u7_U62 (.ZN( u1_u9_u7_n134 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n98 ) );
  NAND2_X1 u1_u9_u7_U63 (.A1( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n102 ) , .ZN( u1_u9_u7_n129 ) );
  NAND2_X1 u1_u9_u7_U64 (.A2( u1_u9_u7_n103 ) , .ZN( u1_u9_u7_n131 ) , .A1( u1_u9_u7_n95 ) );
  NAND2_X1 u1_u9_u7_U65 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n138 ) , .A2( u1_u9_u7_n99 ) );
  NAND2_X1 u1_u9_u7_U66 (.ZN( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n93 ) , .A2( u1_u9_u7_n96 ) );
  NAND2_X1 u1_u9_u7_U67 (.A1( u1_u9_u7_n100 ) , .ZN( u1_u9_u7_n148 ) , .A2( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U68 (.A2( u1_u9_X_47 ) , .ZN( u1_u9_u7_n150 ) , .A1( u1_u9_u7_n163 ) );
  NOR2_X1 u1_u9_u7_U69 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n103 ) );
  AOI211_X1 u1_u9_u7_U7 (.ZN( u1_u9_u7_n116 ) , .A( u1_u9_u7_n155 ) , .C1( u1_u9_u7_n161 ) , .C2( u1_u9_u7_n171 ) , .B( u1_u9_u7_n94 ) );
  NOR2_X1 u1_u9_u7_U70 (.A2( u1_u9_X_48 ) , .A1( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n95 ) );
  NOR2_X1 u1_u9_u7_U71 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n99 ) );
  NOR2_X1 u1_u9_u7_U72 (.A2( u1_u9_X_44 ) , .A1( u1_u9_u7_n167 ) , .ZN( u1_u9_u7_n98 ) );
  NOR2_X1 u1_u9_u7_U73 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n152 ) );
  AND2_X1 u1_u9_u7_U74 (.A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n156 ) , .A2( u1_u9_u7_n163 ) );
  NAND2_X1 u1_u9_u7_U75 (.A2( u1_u9_X_46 ) , .A1( u1_u9_X_47 ) , .ZN( u1_u9_u7_n125 ) );
  AND2_X1 u1_u9_u7_U76 (.A2( u1_u9_X_45 ) , .A1( u1_u9_X_48 ) , .ZN( u1_u9_u7_n102 ) );
  AND2_X1 u1_u9_u7_U77 (.A2( u1_u9_X_43 ) , .A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n96 ) );
  AND2_X1 u1_u9_u7_U78 (.A1( u1_u9_X_44 ) , .ZN( u1_u9_u7_n100 ) , .A2( u1_u9_u7_n167 ) );
  AND2_X1 u1_u9_u7_U79 (.A1( u1_u9_X_48 ) , .A2( u1_u9_u7_n166 ) , .ZN( u1_u9_u7_n93 ) );
  OAI222_X1 u1_u9_u7_U8 (.C2( u1_u9_u7_n101 ) , .B2( u1_u9_u7_n111 ) , .A1( u1_u9_u7_n113 ) , .C1( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n162 ) , .B1( u1_u9_u7_n164 ) , .ZN( u1_u9_u7_n94 ) );
  INV_X1 u1_u9_u7_U80 (.A( u1_u9_X_46 ) , .ZN( u1_u9_u7_n163 ) );
  INV_X1 u1_u9_u7_U81 (.A( u1_u9_X_43 ) , .ZN( u1_u9_u7_n167 ) );
  INV_X1 u1_u9_u7_U82 (.A( u1_u9_X_45 ) , .ZN( u1_u9_u7_n166 ) );
  NAND4_X1 u1_u9_u7_U83 (.ZN( u1_out9_5 ) , .A4( u1_u9_u7_n108 ) , .A3( u1_u9_u7_n109 ) , .A1( u1_u9_u7_n116 ) , .A2( u1_u9_u7_n123 ) );
  AOI22_X1 u1_u9_u7_U84 (.ZN( u1_u9_u7_n109 ) , .A2( u1_u9_u7_n126 ) , .B2( u1_u9_u7_n145 ) , .B1( u1_u9_u7_n156 ) , .A1( u1_u9_u7_n171 ) );
  NOR4_X1 u1_u9_u7_U85 (.A4( u1_u9_u7_n104 ) , .A3( u1_u9_u7_n105 ) , .A2( u1_u9_u7_n106 ) , .A1( u1_u9_u7_n107 ) , .ZN( u1_u9_u7_n108 ) );
  NAND4_X1 u1_u9_u7_U86 (.ZN( u1_out9_27 ) , .A4( u1_u9_u7_n118 ) , .A3( u1_u9_u7_n119 ) , .A2( u1_u9_u7_n120 ) , .A1( u1_u9_u7_n121 ) );
  OAI21_X1 u1_u9_u7_U87 (.ZN( u1_u9_u7_n121 ) , .B2( u1_u9_u7_n145 ) , .A( u1_u9_u7_n150 ) , .B1( u1_u9_u7_n174 ) );
  OAI21_X1 u1_u9_u7_U88 (.ZN( u1_u9_u7_n120 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n170 ) , .B1( u1_u9_u7_n179 ) );
  NAND4_X1 u1_u9_u7_U89 (.ZN( u1_out9_21 ) , .A4( u1_u9_u7_n157 ) , .A3( u1_u9_u7_n158 ) , .A2( u1_u9_u7_n159 ) , .A1( u1_u9_u7_n160 ) );
  OAI221_X1 u1_u9_u7_U9 (.C1( u1_u9_u7_n101 ) , .C2( u1_u9_u7_n147 ) , .ZN( u1_u9_u7_n155 ) , .B2( u1_u9_u7_n162 ) , .A( u1_u9_u7_n91 ) , .B1( u1_u9_u7_n92 ) );
  OAI21_X1 u1_u9_u7_U90 (.B1( u1_u9_u7_n145 ) , .ZN( u1_u9_u7_n160 ) , .A( u1_u9_u7_n161 ) , .B2( u1_u9_u7_n177 ) );
  AOI22_X1 u1_u9_u7_U91 (.B2( u1_u9_u7_n149 ) , .B1( u1_u9_u7_n150 ) , .A2( u1_u9_u7_n151 ) , .A1( u1_u9_u7_n152 ) , .ZN( u1_u9_u7_n158 ) );
  NAND4_X1 u1_u9_u7_U92 (.ZN( u1_out9_15 ) , .A4( u1_u9_u7_n142 ) , .A3( u1_u9_u7_n143 ) , .A2( u1_u9_u7_n144 ) , .A1( u1_u9_u7_n178 ) );
  OR2_X1 u1_u9_u7_U93 (.A2( u1_u9_u7_n125 ) , .A1( u1_u9_u7_n129 ) , .ZN( u1_u9_u7_n144 ) );
  AOI22_X1 u1_u9_u7_U94 (.A2( u1_u9_u7_n126 ) , .ZN( u1_u9_u7_n143 ) , .B2( u1_u9_u7_n165 ) , .B1( u1_u9_u7_n173 ) , .A1( u1_u9_u7_n174 ) );
  NAND3_X1 u1_u9_u7_U95 (.A3( u1_u9_u7_n146 ) , .A2( u1_u9_u7_n147 ) , .A1( u1_u9_u7_n148 ) , .ZN( u1_u9_u7_n151 ) );
  NAND3_X1 u1_u9_u7_U96 (.A3( u1_u9_u7_n131 ) , .A2( u1_u9_u7_n132 ) , .A1( u1_u9_u7_n133 ) , .ZN( u1_u9_u7_n135 ) );
  INV_X1 u1_uk_U10 (.A( u1_uk_n209 ) , .ZN( u1_uk_n83 ) );
  AOI22_X1 u1_uk_U100 (.B2( u1_uk_K_r0_28 ) , .A2( u1_uk_K_r0_49 ) , .ZN( u1_uk_n1031 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1000 (.ZN( u1_K6_23 ) , .A( u1_uk_n1093 ) , .B2( u1_uk_n1472 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1001 (.A1( u1_uk_K_r4_27 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1093 ) );
  OAI21_X1 u1_uk_U1002 (.ZN( u1_K3_35 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1042 ) , .B2( u1_uk_n1308 ) );
  NAND2_X1 u1_uk_U1003 (.A1( u1_uk_K_r1_7 ) , .ZN( u1_uk_n1042 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U1004 (.ZN( u1_K14_46 ) , .B2( u1_uk_n1820 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n961 ) );
  NAND2_X1 u1_uk_U1005 (.A1( u1_uk_K_r12_22 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n961 ) );
  OAI21_X1 u1_uk_U1006 (.ZN( u1_K16_4 ) , .B2( u1_uk_n1257 ) , .B1( u1_uk_n99 ) , .A( u1_uk_n995 ) );
  NAND2_X1 u1_uk_U1007 (.A1( u1_uk_K_r14_3 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n995 ) );
  OAI21_X1 u1_uk_U1008 (.ZN( u1_K8_4 ) , .A( u1_uk_n1146 ) , .B2( u1_uk_n1537 ) , .B1( u1_uk_n17 ) );
  NAND2_X1 u1_uk_U1009 (.A1( u1_uk_K_r6_19 ) , .ZN( u1_uk_n1146 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U101 (.ZN( u1_K15_41 ) , .B2( u1_uk_n1865 ) , .A2( u1_uk_n1883 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1010 (.ZN( u1_K5_4 ) , .A( u1_uk_n1085 ) , .B2( u1_uk_n1411 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1011 (.A1( u1_uk_K_r3_4 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1085 ) );
  OAI21_X1 u1_uk_U1012 (.ZN( u1_K4_5 ) , .A( u1_uk_n1068 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1386 ) );
  NAND2_X1 u1_uk_U1013 (.A1( u1_uk_K_r2_53 ) , .ZN( u1_uk_n1068 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1014 (.ZN( u1_K3_5 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1048 ) , .B2( u1_uk_n1332 ) );
  NAND2_X1 u1_uk_U1015 (.A1( u1_uk_K_r1_10 ) , .ZN( u1_uk_n1048 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1016 (.ZN( u1_K5_45 ) , .A( u1_uk_n1084 ) , .B2( u1_uk_n1400 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1017 (.A1( u1_uk_K_r3_43 ) , .ZN( u1_uk_n1084 ) , .A2( u1_uk_n11 ) );
  OAI21_X1 u1_uk_U1018 (.ZN( u1_K3_45 ) , .A( u1_uk_n1046 ) , .B2( u1_uk_n1335 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U1019 (.A1( u1_uk_K_r1_16 ) , .ZN( u1_uk_n1046 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U102 (.ZN( u1_K13_41 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1753 ) , .A2( u1_uk_n1768 ) , .A1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U1020 (.ZN( u1_K1_13 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1214 ) , .A( u1_uk_n999 ) );
  NAND2_X1 u1_uk_U1021 (.A1( u1_key_r_46 ) , .A2( u1_uk_n146 ) , .ZN( u1_uk_n999 ) );
  OAI21_X1 u1_uk_U1022 (.ZN( u1_K1_17 ) , .A( u1_uk_n1001 ) , .B2( u1_uk_n1183 ) , .B1( u1_uk_n129 ) );
  NAND2_X1 u1_uk_U1023 (.A1( u1_key_r_10 ) , .ZN( u1_uk_n1001 ) , .A2( u1_uk_n187 ) );
  OAI21_X1 u1_uk_U1024 (.ZN( u1_K10_21 ) , .B2( u1_uk_n1660 ) , .A( u1_uk_n308 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1025 (.A1( u1_uk_K_r8_19 ) , .ZN( u1_uk_n308 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1026 (.ZN( u1_K1_37 ) , .A( u1_uk_n1013 ) , .B2( u1_uk_n1174 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U1027 (.A1( u1_key_r_50 ) , .ZN( u1_uk_n1013 ) , .A2( u1_uk_n162 ) );
  OAI21_X1 u1_uk_U1028 (.ZN( u1_K9_39 ) , .A( u1_uk_n1165 ) , .B2( u1_uk_n1601 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1029 (.A1( u1_uk_K_r7_31 ) , .ZN( u1_uk_n1165 ) , .A2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U103 (.ZN( u1_K7_41 ) , .A2( u1_uk_n1486 ) , .B2( u1_uk_n1516 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U1030 (.ZN( u1_K14_44 ) , .B2( u1_uk_n1807 ) , .B1( u1_uk_n251 ) , .A( u1_uk_n959 ) );
  NAND2_X1 u1_uk_U1031 (.A1( u1_uk_K_r12_15 ) , .A2( u1_uk_n279 ) , .ZN( u1_uk_n959 ) );
  OAI21_X1 u1_uk_U1032 (.ZN( u1_K9_44 ) , .A( u1_uk_n1168 ) , .B2( u1_uk_n1615 ) , .B1( u1_uk_n223 ) );
  NAND2_X1 u1_uk_U1033 (.A1( u1_uk_K_r7_0 ) , .ZN( u1_uk_n1168 ) , .A2( u1_uk_n207 ) );
  OAI21_X1 u1_uk_U1034 (.ZN( u1_K12_6 ) , .B2( u1_uk_n1732 ) , .B1( u1_uk_n230 ) , .A( u1_uk_n662 ) );
  NAND2_X1 u1_uk_U1035 (.A1( u1_uk_K_r10_10 ) , .A2( u1_uk_n251 ) , .ZN( u1_uk_n662 ) );
  OAI21_X1 u1_uk_U1036 (.ZN( u1_K8_46 ) , .A( u1_uk_n1145 ) , .B2( u1_uk_n1562 ) , .B1( u1_uk_n188 ) );
  NAND2_X1 u1_uk_U1037 (.A1( u1_uk_K_r6_37 ) , .ZN( u1_uk_n1145 ) , .A2( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U1038 (.ZN( u1_K10_13 ) , .B2( u1_uk_n1635 ) , .A( u1_uk_n301 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1039 (.A1( u1_uk_K_r8_48 ) , .ZN( u1_uk_n301 ) , .A2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U104 (.ZN( u1_K4_41 ) , .B2( u1_uk_n1349 ) , .A2( u1_uk_n1366 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U1040 (.ZN( u1_K12_36 ) , .B2( u1_uk_n1728 ) , .A( u1_uk_n587 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1041 (.A1( u1_uk_K_r10_52 ) , .A2( u1_uk_n110 ) , .ZN( u1_uk_n587 ) );
  OAI21_X1 u1_uk_U1042 (.ZN( u1_K16_41 ) , .B2( u1_uk_n1245 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n991 ) );
  NAND2_X1 u1_uk_U1043 (.A1( u1_uk_K_r14_42 ) , .A2( u1_uk_n141 ) , .ZN( u1_uk_n991 ) );
  OAI21_X1 u1_uk_U1044 (.ZN( u1_K8_41 ) , .A( u1_uk_n1141 ) , .B2( u1_uk_n1547 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U1045 (.A1( u1_uk_K_r6_30 ) , .ZN( u1_uk_n1141 ) , .A2( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U1046 (.ZN( u1_K6_41 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1099 ) , .B2( u1_uk_n1475 ) );
  NAND2_X1 u1_uk_U1047 (.A1( u1_uk_K_r4_31 ) , .ZN( u1_uk_n1099 ) , .A2( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U1048 (.ZN( u1_K16_28 ) , .B2( u1_uk_n1219 ) , .A( u1_uk_n984 ) , .B1( u1_uk_n99 ) );
  NAND2_X1 u1_uk_U1049 (.A1( u1_uk_K_r14_8 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n984 ) );
  OAI21_X1 u1_uk_U1050 (.ZN( u1_K8_28 ) , .A( u1_uk_n1133 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1562 ) );
  NAND2_X1 u1_uk_U1051 (.A1( u1_uk_K_r6_51 ) , .ZN( u1_uk_n1133 ) , .A2( u1_uk_n145 ) );
  OAI21_X1 u1_uk_U1052 (.ZN( u1_K4_28 ) , .A( u1_uk_n1059 ) , .B2( u1_uk_n1381 ) , .B1( u1_uk_n148 ) );
  NAND2_X1 u1_uk_U1053 (.A1( u1_uk_K_r2_21 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1059 ) );
  OAI21_X1 u1_uk_U1054 (.ZN( u1_K9_14 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1151 ) , .B2( u1_uk_n1604 ) );
  NAND2_X1 u1_uk_U1055 (.A1( u1_uk_K_r7_34 ) , .A2( u1_uk_n100 ) , .ZN( u1_uk_n1151 ) );
  OAI21_X1 u1_uk_U1056 (.ZN( u1_K7_31 ) , .A( u1_uk_n1117 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1508 ) );
  NAND2_X1 u1_uk_U1057 (.A1( u1_uk_K_r5_16 ) , .ZN( u1_uk_n1117 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1058 (.ZN( u1_K14_40 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1823 ) , .A( u1_uk_n958 ) );
  NAND2_X1 u1_uk_U1059 (.A1( u1_uk_K_r12_21 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n958 ) );
  AOI22_X1 u1_uk_U106 (.B2( u1_uk_K_r9_19 ) , .A2( u1_uk_K_r9_25 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n250 ) , .ZN( u1_uk_n496 ) );
  OAI21_X1 u1_uk_U1060 (.ZN( u1_K12_40 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1729 ) , .A( u1_uk_n603 ) );
  NAND2_X1 u1_uk_U1061 (.A1( u1_uk_K_r10_49 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n603 ) );
  OAI21_X1 u1_uk_U1062 (.ZN( u1_K15_14 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1851 ) , .A( u1_uk_n966 ) );
  NAND2_X1 u1_uk_U1063 (.A1( u1_uk_K_r13_32 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n966 ) );
  OAI21_X1 u1_uk_U1064 (.ZN( u1_K10_32 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1618 ) , .A( u1_uk_n346 ) );
  NAND2_X1 u1_uk_U1065 (.A1( u1_uk_K_r8_51 ) , .A2( u1_uk_n142 ) , .ZN( u1_uk_n346 ) );
  OAI21_X1 u1_uk_U1066 (.ZN( u1_K15_32 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1855 ) , .A( u1_uk_n971 ) );
  NAND2_X1 u1_uk_U1067 (.A1( u1_uk_K_r13_36 ) , .A2( u1_uk_n147 ) , .ZN( u1_uk_n971 ) );
  OAI21_X1 u1_uk_U1068 (.ZN( u1_K16_42 ) , .B2( u1_uk_n1241 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n992 ) );
  NAND2_X1 u1_uk_U1069 (.A1( u1_uk_K_r14_38 ) , .A2( u1_uk_n31 ) , .ZN( u1_uk_n992 ) );
  OAI22_X1 u1_uk_U107 (.ZN( u1_K1_5 ) , .A2( u1_uk_n1176 ) , .B2( u1_uk_n1180 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U1070 (.ZN( u1_K8_42 ) , .A( u1_uk_n1142 ) , .B2( u1_uk_n1540 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U1071 (.A1( u1_uk_K_r6_22 ) , .ZN( u1_uk_n1142 ) , .A2( u1_uk_n117 ) );
  OAI21_X1 u1_uk_U1072 (.ZN( u1_K7_38 ) , .A( u1_uk_n1122 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1499 ) );
  NAND2_X1 u1_uk_U1073 (.A1( u1_uk_K_r5_8 ) , .ZN( u1_uk_n1122 ) , .A2( u1_uk_n17 ) );
  OAI21_X1 u1_uk_U1074 (.ZN( u1_K5_42 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1082 ) , .B2( u1_uk_n1412 ) );
  NAND2_X1 u1_uk_U1075 (.A1( u1_uk_K_r3_9 ) , .ZN( u1_uk_n1082 ) , .A2( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1076 (.ZN( u1_K4_38 ) , .A( u1_uk_n1064 ) , .B2( u1_uk_n1383 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U1077 (.A1( u1_uk_K_r2_50 ) , .ZN( u1_uk_n1064 ) , .A2( u1_uk_n155 ) );
  INV_X1 u1_uk_U1078 (.A( u1_key_r_9 ) , .ZN( u1_uk_n1179 ) );
  INV_X1 u1_uk_U1079 (.A( u1_key_r_7 ) , .ZN( u1_uk_n1177 ) );
  OAI22_X1 u1_uk_U108 (.ZN( u1_K16_5 ) , .A2( u1_uk_n1221 ) , .B2( u1_uk_n1224 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n294 ) );
  INV_X1 u1_uk_U1080 (.A( u1_key_r_6 ) , .ZN( u1_uk_n1176 ) );
  INV_X1 u1_uk_U1081 (.A( u1_key_r_54 ) , .ZN( u1_uk_n1215 ) );
  INV_X1 u1_uk_U1082 (.A( u1_key_r_33 ) , .ZN( u1_uk_n1197 ) );
  INV_X1 u1_uk_U1083 (.A( u1_key_r_23 ) , .ZN( u1_uk_n1188 ) );
  INV_X1 u1_uk_U1084 (.A( u1_key_r_26 ) , .ZN( u1_uk_n1191 ) );
  INV_X1 u1_uk_U1085 (.A( u1_key_r_40 ) , .ZN( u1_uk_n1204 ) );
  INV_X1 u1_uk_U1086 (.A( u1_key_r_30 ) , .ZN( u1_uk_n1195 ) );
  INV_X1 u1_uk_U1087 (.A( u1_key_r_47 ) , .ZN( u1_uk_n1209 ) );
  INV_X1 u1_uk_U1088 (.A( u1_key_r_34 ) , .ZN( u1_uk_n1198 ) );
  INV_X1 u1_uk_U1089 (.A( u1_key_r_27 ) , .ZN( u1_uk_n1192 ) );
  OAI22_X1 u1_uk_U109 (.ZN( u1_K15_5 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1859 ) , .A2( u1_uk_n1862 ) , .B1( u1_uk_n217 ) );
  INV_X1 u1_uk_U1090 (.A( u1_key_r_24 ) , .ZN( u1_uk_n1189 ) );
  INV_X1 u1_uk_U1091 (.A( u1_key_r_20 ) , .ZN( u1_uk_n1185 ) );
  INV_X1 u1_uk_U1092 (.A( u1_key_r_37 ) , .ZN( u1_uk_n1201 ) );
  INV_X1 u1_uk_U1093 (.A( u1_key_r_52 ) , .ZN( u1_uk_n1213 ) );
  INV_X1 u1_uk_U1094 (.A( u1_key_r_0 ) , .ZN( u1_uk_n1172 ) );
  INV_X1 u1_uk_U1095 (.A( u1_key_r_16 ) , .ZN( u1_uk_n1182 ) );
  INV_X1 u1_uk_U1096 (.A( u1_key_r_13 ) , .ZN( u1_uk_n1180 ) );
  INV_X1 u1_uk_U1097 (.A( u1_key_r_1 ) , .ZN( u1_uk_n1173 ) );
  INV_X1 u1_uk_U1098 (.A( u1_key_r_2 ) , .ZN( u1_uk_n1174 ) );
  INV_X1 u1_uk_U1099 (.A( u1_key_r_19 ) , .ZN( u1_uk_n1184 ) );
  INV_X1 u1_uk_U11 (.A( u1_uk_n298 ) , .ZN( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U110 (.ZN( u1_K14_5 ) , .B2( u1_uk_n1826 ) , .B1( u1_uk_n250 ) , .A( u1_uk_n962 ) );
  INV_X1 u1_uk_U1100 (.A( u1_key_r_4 ) , .ZN( u1_uk_n1175 ) );
  INV_X1 u1_uk_U1101 (.A( u1_key_r_17 ) , .ZN( u1_uk_n1183 ) );
  INV_X1 u1_uk_U1102 (.A( u1_key_r_53 ) , .ZN( u1_uk_n1214 ) );
  OAI21_X1 u1_uk_U1103 (.ZN( u1_K13_28 ) , .B2( u1_uk_n1783 ) , .B1( u1_uk_n230 ) , .A( u1_uk_n695 ) );
  NAND2_X1 u1_uk_U1104 (.A1( u1_uk_K_r11_21 ) , .A2( u1_uk_n277 ) , .ZN( u1_uk_n695 ) );
  OAI21_X1 u1_uk_U1105 (.ZN( u1_K8_14 ) , .A( u1_uk_n1129 ) , .B2( u1_uk_n1559 ) , .B1( u1_uk_n203 ) );
  NAND2_X1 u1_uk_U1106 (.A1( u1_uk_K_r6_34 ) , .ZN( u1_uk_n1129 ) , .A2( u1_uk_n291 ) );
  OAI21_X1 u1_uk_U1107 (.ZN( u1_K16_14 ) , .B2( u1_uk_n1235 ) , .B1( u1_uk_n252 ) , .A( u1_uk_n981 ) );
  NAND2_X1 u1_uk_U1108 (.A1( u1_uk_K_r14_18 ) , .A2( u1_uk_n291 ) , .ZN( u1_uk_n981 ) );
  OAI21_X1 u1_uk_U1109 (.ZN( u1_K3_40 ) , .A( u1_uk_n1044 ) , .B2( u1_uk_n1330 ) , .B1( u1_uk_n209 ) );
  NAND2_X1 u1_uk_U111 (.A1( u1_uk_K_r12_10 ) , .A2( u1_uk_n298 ) , .ZN( u1_uk_n962 ) );
  NAND2_X1 u1_uk_U1110 (.A1( u1_uk_K_r1_21 ) , .ZN( u1_uk_n1044 ) , .A2( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U1111 (.ZN( u1_K16_39 ) , .B2( u1_uk_n1231 ) , .B1( u1_uk_n291 ) , .A( u1_uk_n990 ) );
  NAND2_X1 u1_uk_U1112 (.A1( u1_uk_K_r14_15 ) , .A2( u1_uk_n214 ) , .ZN( u1_uk_n990 ) );
  OAI21_X1 u1_uk_U1113 (.ZN( u1_K8_39 ) , .A( u1_uk_n1139 ) , .B2( u1_uk_n1556 ) , .B1( u1_uk_n203 ) );
  NAND2_X1 u1_uk_U1114 (.A1( u1_uk_K_r6_31 ) , .ZN( u1_uk_n1139 ) , .A2( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U1115 (.ZN( u1_K5_39 ) , .A( u1_uk_n1081 ) , .B2( u1_uk_n1406 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U1116 (.A1( u1_uk_K_r3_16 ) , .ZN( u1_uk_n1081 ) , .A2( u1_uk_n242 ) );
  AOI22_X1 u1_uk_U1118 (.B2( u1_uk_K_r11_26 ) , .A2( u1_uk_K_r11_6 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n203 ) , .ZN( u1_uk_n671 ) );
  INV_X1 u1_uk_U1119 (.ZN( u1_K9_11 ) , .A( u1_uk_n1148 ) );
  INV_X1 u1_uk_U112 (.ZN( u1_K13_5 ) , .A( u1_uk_n948 ) );
  AOI22_X1 u1_uk_U1120 (.B2( u1_uk_K_r7_48 ) , .A2( u1_uk_K_r7_55 ) , .B1( u1_uk_n109 ) , .ZN( u1_uk_n1148 ) , .A1( u1_uk_n220 ) );
  AOI22_X1 u1_uk_U1122 (.B2( u1_uk_K_r0_34 ) , .A2( u1_uk_K_r0_55 ) , .ZN( u1_uk_n1021 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) );
  INV_X1 u1_uk_U1123 (.ZN( u1_K1_11 ) , .A( u1_uk_n997 ) );
  AOI22_X1 u1_uk_U1124 (.B2( u1_key_r_32 ) , .A2( u1_key_r_39 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n277 ) , .ZN( u1_uk_n997 ) );
  INV_X1 u1_uk_U1125 (.ZN( u1_K1_18 ) , .A( u1_uk_n1002 ) );
  AOI22_X1 u1_uk_U1126 (.A2( u1_key_r_5 ) , .B2( u1_key_r_55 ) , .ZN( u1_uk_n1002 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n294 ) );
  INV_X1 u1_uk_U1127 (.ZN( u1_K1_41 ) , .A( u1_uk_n1015 ) );
  AOI22_X1 u1_uk_U1128 (.B2( u1_key_r_35 ) , .A2( u1_key_r_42 ) , .ZN( u1_uk_n1015 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n298 ) );
  AOI22_X1 u1_uk_U113 (.B2( u1_uk_K_r11_48 ) , .A2( u1_uk_K_r11_53 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n223 ) , .ZN( u1_uk_n948 ) );
  AOI22_X1 u1_uk_U1130 (.B2( u1_uk_K_r9_12 ) , .A2( u1_uk_K_r9_18 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n501 ) );
  INV_X1 u1_uk_U1131 (.ZN( u1_K11_12 ) , .A( u1_uk_n379 ) );
  AOI22_X1 u1_uk_U1132 (.B2( u1_uk_K_r9_25 ) , .A2( u1_uk_K_r9_6 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n291 ) , .ZN( u1_uk_n379 ) );
  INV_X1 u1_uk_U1133 (.ZN( u1_K8_12 ) , .A( u1_uk_n1128 ) );
  AOI22_X1 u1_uk_U1134 (.B2( u1_uk_K_r6_3 ) , .A2( u1_uk_K_r6_53 ) , .ZN( u1_uk_n1128 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) );
  INV_X1 u1_uk_U1135 (.ZN( u1_K2_7 ) , .A( u1_uk_n1034 ) );
  AOI22_X1 u1_uk_U1136 (.B2( u1_uk_K_r0_13 ) , .A2( u1_uk_K_r0_34 ) , .ZN( u1_uk_n1034 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n27 ) );
  INV_X1 u1_uk_U1137 (.ZN( u1_K1_20 ) , .A( u1_uk_n1003 ) );
  AOI22_X1 u1_uk_U1138 (.B2( u1_key_r_48 ) , .A2( u1_key_r_55 ) , .ZN( u1_uk_n1003 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U114 (.ZN( u1_K12_5 ) , .A2( u1_uk_n1712 ) , .B2( u1_uk_n1738 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n99 ) );
  AOI22_X1 u1_uk_U1140 (.B2( u1_uk_K_r9_1 ) , .A2( u1_uk_K_r9_9 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n421 ) );
  INV_X1 u1_uk_U1141 (.ZN( u1_K12_32 ) , .A( u1_uk_n582 ) );
  AOI22_X1 u1_uk_U1142 (.B2( u1_uk_K_r10_23 ) , .A2( u1_uk_K_r10_28 ) , .B1( u1_uk_n10 ) , .A1( u1_uk_n294 ) , .ZN( u1_uk_n582 ) );
  INV_X1 u1_uk_U1143 (.ZN( u1_K2_32 ) , .A( u1_uk_n1029 ) );
  AOI22_X1 u1_uk_U1144 (.B2( u1_uk_K_r0_15 ) , .A2( u1_uk_K_r0_36 ) , .ZN( u1_uk_n1029 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n271 ) );
  INV_X1 u1_uk_U1145 (.ZN( u1_K9_20 ) , .A( u1_uk_n1156 ) );
  AOI22_X1 u1_uk_U1146 (.B2( u1_uk_K_r7_32 ) , .A2( u1_uk_K_r7_39 ) , .B1( u1_uk_n11 ) , .ZN( u1_uk_n1156 ) , .A1( u1_uk_n294 ) );
  INV_X1 u1_uk_U1147 (.ZN( u1_K4_20 ) , .A( u1_uk_n1054 ) );
  AOI22_X1 u1_uk_U1148 (.B2( u1_uk_K_r2_13 ) , .A2( u1_uk_K_r2_33 ) , .ZN( u1_uk_n1054 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n207 ) );
  INV_X1 u1_uk_U1149 (.ZN( u1_K7_13 ) , .A( u1_uk_n1106 ) );
  OAI22_X1 u1_uk_U115 (.ZN( u1_K9_5 ) , .B2( u1_uk_n1610 ) , .A2( u1_uk_n1616 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n188 ) );
  AOI22_X1 u1_uk_U1150 (.B2( u1_uk_K_r5_26 ) , .A2( u1_uk_K_r5_48 ) , .ZN( u1_uk_n1106 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n217 ) );
  INV_X1 u1_uk_U1151 (.ZN( u1_K1_32 ) , .A( u1_uk_n1010 ) );
  AOI22_X1 u1_uk_U1152 (.B2( u1_key_r_22 ) , .A2( u1_key_r_29 ) , .ZN( u1_uk_n1010 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) );
  INV_X1 u1_uk_U1153 (.ZN( u1_K7_32 ) , .A( u1_uk_n1118 ) );
  AOI22_X1 u1_uk_U1154 (.B2( u1_uk_K_r5_0 ) , .A2( u1_uk_K_r5_51 ) , .ZN( u1_uk_n1118 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n222 ) );
  INV_X1 u1_uk_U1155 (.ZN( u1_K6_2 ) , .A( u1_uk_n1096 ) );
  AOI22_X1 u1_uk_U1156 (.B2( u1_uk_K_r4_17 ) , .A2( u1_uk_K_r4_55 ) , .ZN( u1_uk_n1096 ) , .B1( u1_uk_n257 ) , .A1( u1_uk_n27 ) );
  AOI22_X1 u1_uk_U1158 (.B2( u1_uk_K_r8_17 ) , .A2( u1_uk_K_r8_39 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n297 ) , .ZN( u1_uk_n299 ) );
  INV_X1 u1_uk_U1159 (.ZN( u1_K8_15 ) , .A( u1_uk_n1130 ) );
  OAI22_X1 u1_uk_U116 (.ZN( u1_K7_5 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1487 ) , .A2( u1_uk_n1504 ) , .B1( u1_uk_n242 ) );
  AOI22_X1 u1_uk_U1160 (.B2( u1_uk_K_r6_10 ) , .A2( u1_uk_K_r6_17 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1130 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U1161 (.ZN( u1_K7_25 ) , .A( u1_uk_n1114 ) );
  AOI22_X1 u1_uk_U1162 (.B2( u1_uk_K_r5_31 ) , .A2( u1_uk_K_r5_7 ) , .A1( u1_uk_n10 ) , .ZN( u1_uk_n1114 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U1163 (.ZN( u1_K13_12 ) , .A( u1_uk_n676 ) );
  AOI22_X1 u1_uk_U1164 (.B2( u1_uk_K_r11_34 ) , .A2( u1_uk_K_r11_54 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n252 ) , .ZN( u1_uk_n676 ) );
  AOI22_X1 u1_uk_U1165 (.B1( n116 ) , .A2( u1_uk_K_r13_2 ) , .B2( u1_uk_K_r13_23 ) , .A1( u1_uk_n286 ) , .ZN( u1_uk_n974 ) );
  INV_X1 u1_uk_U1166 (.ZN( u1_K15_43 ) , .A( u1_uk_n974 ) );
  AOI22_X1 u1_uk_U1167 (.B2( u1_uk_K_r11_26 ) , .A2( u1_uk_K_r11_46 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n27 ) , .ZN( u1_uk_n702 ) );
  INV_X1 u1_uk_U1168 (.ZN( u1_K13_2 ) , .A( u1_uk_n702 ) );
  INV_X1 u1_uk_U1169 (.ZN( u1_K12_1 ) , .A( u1_uk_n515 ) );
  OAI22_X1 u1_uk_U117 (.ZN( u1_K5_5 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1398 ) , .B2( u1_uk_n1422 ) , .B1( u1_uk_n242 ) );
  INV_X1 u1_uk_U1170 (.ZN( u1_K9_2 ) , .A( u1_uk_n1160 ) );
  INV_X1 u1_uk_U1171 (.ZN( u1_K4_2 ) , .A( u1_uk_n1061 ) );
  INV_X1 u1_uk_U1172 (.ZN( u1_K13_6 ) , .A( u1_uk_n949 ) );
  OAI22_X1 u1_uk_U118 (.ZN( u1_K2_5 ) , .B2( u1_uk_n1274 ) , .A2( u1_uk_n1277 ) , .A1( u1_uk_n291 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U119 (.ZN( u1_K10_41 ) , .A2( u1_uk_n1624 ) , .B2( u1_uk_n1652 ) , .A1( u1_uk_n223 ) , .B1( u1_uk_n31 ) );
  INV_X1 u1_uk_U12 (.A( u1_uk_n208 ) , .ZN( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U120 (.ZN( u1_K14_41 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1806 ) , .B2( u1_uk_n1811 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U121 (.ZN( u1_K12_41 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1735 ) , .A2( u1_uk_n1744 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U122 (.ZN( u1_K3_41 ) , .A2( u1_uk_n1313 ) , .B2( u1_uk_n1318 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U123 (.ZN( u1_K16_47 ) , .B2( u1_uk_n1218 ) , .A2( u1_uk_n1222 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U124 (.ZN( u1_K13_47 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1782 ) , .A2( u1_uk_n1792 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U125 (.ZN( u1_K12_47 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1709 ) , .A2( u1_uk_n1736 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U126 (.ZN( u1_K11_47 ) , .A( u1_uk_n472 ) );
  AOI22_X1 u1_uk_U127 (.B2( u1_uk_K_r9_15 ) , .A2( u1_uk_K_r9_23 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n223 ) , .ZN( u1_uk_n472 ) );
  OAI22_X1 u1_uk_U128 (.ZN( u1_K10_47 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1624 ) , .B2( u1_uk_n1639 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U129 (.ZN( u1_K8_47 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1561 ) , .A2( u1_uk_n1567 ) , .A1( u1_uk_n294 ) );
  INV_X1 u1_uk_U13 (.A( u1_uk_n222 ) , .ZN( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U130 (.ZN( u1_K7_47 ) , .A2( u1_uk_n1486 ) , .B2( u1_uk_n1500 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U131 (.ZN( u1_K6_47 ) , .A( u1_uk_n1100 ) , .B1( u1_uk_n142 ) , .B2( u1_uk_n1449 ) );
  NAND2_X1 u1_uk_U132 (.A1( u1_uk_K_r4_23 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1100 ) );
  OAI22_X1 u1_uk_U133 (.ZN( u1_K5_47 ) , .B2( u1_uk_n1395 ) , .A2( u1_uk_n1419 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U134 (.ZN( u1_K4_47 ) , .B2( u1_uk_n1380 ) , .A2( u1_uk_n1389 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U135 (.ZN( u1_K2_47 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1033 ) , .B2( u1_uk_n1271 ) );
  NAND2_X1 u1_uk_U136 (.A1( u1_uk_K_r0_52 ) , .ZN( u1_uk_n1033 ) , .A2( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U137 (.ZN( u1_K1_15 ) , .B2( u1_uk_n1191 ) , .A2( u1_uk_n1197 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U138 (.ZN( u1_K4_15 ) , .B2( u1_uk_n1358 ) , .A2( u1_uk_n1386 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U139 (.ZN( u1_K5_15 ) , .A( u1_uk_n1072 ) , .B2( u1_uk_n1409 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U14 (.ZN( u1_uk_n100 ) , .A( u1_uk_n213 ) );
  NAND2_X1 u1_uk_U140 (.A1( u1_uk_K_r3_34 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1072 ) );
  AOI22_X1 u1_uk_U142 (.B2( u1_uk_K_r11_11 ) , .A2( u1_uk_K_r11_48 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n678 ) );
  OAI22_X1 u1_uk_U143 (.ZN( u1_K7_15 ) , .A2( u1_uk_n1484 ) , .B2( u1_uk_n1524 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n92 ) );
  INV_X1 u1_uk_U144 (.ZN( u1_K12_15 ) , .A( u1_uk_n504 ) );
  AOI22_X1 u1_uk_U145 (.B2( u1_uk_K_r10_25 ) , .A2( u1_uk_K_r10_34 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n252 ) , .ZN( u1_uk_n504 ) );
  OAI22_X1 u1_uk_U146 (.ZN( u1_K3_15 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1312 ) , .B2( u1_uk_n1347 ) , .A1( u1_uk_n286 ) );
  INV_X1 u1_uk_U147 (.ZN( u1_K13_19 ) , .A( u1_uk_n685 ) );
  AOI22_X1 u1_uk_U148 (.B2( u1_uk_K_r11_19 ) , .A2( u1_uk_K_r11_39 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n252 ) , .ZN( u1_uk_n685 ) );
  OAI22_X1 u1_uk_U149 (.ZN( u1_K11_15 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1676 ) , .A2( u1_uk_n1691 ) , .A1( u1_uk_n297 ) );
  INV_X1 u1_uk_U15 (.A( u1_uk_n188 ) , .ZN( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U150 (.ZN( u1_K6_19 ) , .A( u1_uk_n1091 ) , .B2( u1_uk_n1444 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U151 (.A1( u1_uk_K_r4_48 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1091 ) );
  OAI21_X1 u1_uk_U152 (.ZN( u1_K2_15 ) , .A( u1_uk_n1024 ) , .B2( u1_uk_n1291 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U153 (.A1( u1_uk_K_r0_19 ) , .ZN( u1_uk_n1024 ) , .A2( u1_uk_n118 ) );
  OAI22_X1 u1_uk_U154 (.ZN( u1_K1_19 ) , .B2( u1_uk_n1175 ) , .A2( u1_uk_n1215 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U155 (.ZN( u1_K16_15 ) , .B2( u1_uk_n1236 ) , .A2( u1_uk_n1243 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U156 (.ZN( u1_K10_15 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1622 ) , .B2( u1_uk_n1659 ) , .B1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U157 (.ZN( u1_K15_15 ) , .B2( u1_uk_n1873 ) , .B1( u1_uk_n222 ) , .A( u1_uk_n967 ) );
  NAND2_X1 u1_uk_U158 (.A1( u1_uk_K_r13_19 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n967 ) );
  INV_X1 u1_uk_U159 (.ZN( u1_K14_19 ) , .A( u1_uk_n951 ) );
  INV_X1 u1_uk_U16 (.ZN( u1_uk_n109 ) , .A( u1_uk_n231 ) );
  AOI22_X1 u1_uk_U160 (.B2( u1_uk_K_r12_25 ) , .A2( u1_uk_K_r12_33 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n951 ) );
  AOI22_X1 u1_uk_U162 (.B2( u1_uk_K_r9_10 ) , .A2( u1_uk_K_r9_48 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n222 ) , .ZN( u1_uk_n386 ) );
  INV_X1 u1_uk_U163 (.ZN( u1_K9_19 ) , .A( u1_uk_n1154 ) );
  AOI22_X1 u1_uk_U164 (.B1( u1_uk_K_r7_13 ) , .A2( u1_uk_K_r7_20 ) , .ZN( u1_uk_n1154 ) , .A1( u1_uk_n291 ) , .B2( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U165 (.ZN( u1_K7_19 ) , .B2( u1_uk_n1495 ) , .A2( u1_uk_n1505 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U166 (.ZN( u1_K4_19 ) , .B2( u1_uk_n1365 ) , .A2( u1_uk_n1377 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U167 (.ZN( u1_K3_19 ) , .A( u1_uk_n1037 ) , .B2( u1_uk_n1324 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U168 (.A1( u1_uk_K_r1_33 ) , .ZN( u1_uk_n1037 ) , .A2( u1_uk_n63 ) );
  INV_X1 u1_uk_U169 (.ZN( u1_K2_19 ) , .A( u1_uk_n1025 ) );
  INV_X1 u1_uk_U17 (.ZN( u1_uk_n110 ) , .A( u1_uk_n209 ) );
  AOI22_X1 u1_uk_U170 (.B2( u1_uk_K_r0_11 ) , .A2( u1_uk_K_r0_47 ) , .ZN( u1_uk_n1025 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U171 (.ZN( u1_K14_15 ) , .A1( u1_uk_n146 ) , .A2( u1_uk_n1803 ) , .B2( u1_uk_n1841 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U172 (.ZN( u1_K8_19 ) , .B2( u1_uk_n1538 ) , .A2( u1_uk_n1545 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U173 (.ZN( u1_K10_19 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1633 ) , .A2( u1_uk_n1643 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U174 (.ZN( u1_K5_30 ) , .B2( u1_uk_n1408 ) , .A2( u1_uk_n1425 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U175 (.ZN( u1_K2_30 ) , .B2( u1_uk_n1260 ) , .A2( u1_uk_n1289 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U176 (.ZN( u1_K14_30 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1811 ) , .A2( u1_uk_n1838 ) , .B1( u1_uk_n223 ) );
  INV_X1 u1_uk_U177 (.ZN( u1_K12_30 ) , .A( u1_uk_n526 ) );
  AOI22_X1 u1_uk_U178 (.B2( u1_uk_K_r10_23 ) , .A2( u1_uk_K_r10_42 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n271 ) , .ZN( u1_uk_n526 ) );
  OAI22_X1 u1_uk_U179 (.ZN( u1_K10_30 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1628 ) , .A2( u1_uk_n1656 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U18 (.ZN( u1_uk_n118 ) , .A( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U180 (.ZN( u1_K12_24 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1716 ) , .A2( u1_uk_n1745 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U181 (.ZN( u1_K1_14 ) , .A( u1_uk_n1000 ) , .B2( u1_uk_n1190 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U182 (.A1( u1_key_r_18 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1000 ) );
  INV_X1 u1_uk_U183 (.A( u1_key_r_25 ) , .ZN( u1_uk_n1190 ) );
  OAI21_X1 u1_uk_U184 (.ZN( u1_K8_30 ) , .A( u1_uk_n1136 ) , .B2( u1_uk_n1555 ) , .B1( u1_uk_n207 ) );
  NAND2_X1 u1_uk_U185 (.A1( u1_uk_K_r6_29 ) , .ZN( u1_uk_n1136 ) , .A2( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U186 (.ZN( u1_K16_30 ) , .B2( u1_uk_n1256 ) , .B1( u1_uk_n222 ) , .A( u1_uk_n987 ) );
  NAND2_X1 u1_uk_U187 (.A1( u1_uk_K_r14_45 ) , .A2( u1_uk_n279 ) , .ZN( u1_uk_n987 ) );
  OAI22_X1 u1_uk_U188 (.ZN( u1_K13_14 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1756 ) , .A2( u1_uk_n1780 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U189 (.ZN( u1_K12_14 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1718 ) , .A2( u1_uk_n1723 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U19 (.ZN( u1_uk_n141 ) , .A( u1_uk_n238 ) );
  INV_X1 u1_uk_U190 (.ZN( u1_K11_14 ) , .A( u1_uk_n382 ) );
  AOI22_X1 u1_uk_U191 (.B2( u1_uk_K_r9_12 ) , .A2( u1_uk_K_r9_6 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n207 ) , .ZN( u1_uk_n382 ) );
  OAI21_X1 u1_uk_U192 (.ZN( u1_K10_24 ) , .B2( u1_uk_n1629 ) , .B1( u1_uk_n17 ) , .A( u1_uk_n319 ) );
  NAND2_X1 u1_uk_U193 (.A1( u1_uk_K_r8_40 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n319 ) );
  OAI22_X1 u1_uk_U194 (.ZN( u1_K6_14 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1440 ) , .B2( u1_uk_n1446 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U195 (.ZN( u1_K2_14 ) , .A( u1_uk_n1023 ) );
  AOI22_X1 u1_uk_U196 (.B2( u1_uk_K_r0_11 ) , .A2( u1_uk_K_r0_32 ) , .ZN( u1_uk_n1023 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U197 (.ZN( u1_K1_24 ) , .B2( u1_uk_n1180 ) , .A2( u1_uk_n1185 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U198 (.ZN( u1_K10_14 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1630 ) , .A2( u1_uk_n1661 ) , .B1( u1_uk_n213 ) );
  OAI21_X1 u1_uk_U199 (.ZN( u1_K13_30 ) , .B2( u1_uk_n1776 ) , .A( u1_uk_n717 ) , .B1( u1_uk_n83 ) );
  INV_X1 u1_uk_U20 (.ZN( u1_uk_n142 ) , .A( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U200 (.A1( u1_uk_K_r11_28 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n717 ) );
  OAI21_X1 u1_uk_U201 (.ZN( u1_K14_24 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1812 ) , .A( u1_uk_n952 ) );
  NAND2_X1 u1_uk_U202 (.A1( u1_uk_K_r12_41 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n952 ) );
  INV_X1 u1_uk_U203 (.ZN( u1_K7_24 ) , .A( u1_uk_n1113 ) );
  AOI22_X1 u1_uk_U204 (.B2( u1_uk_K_r5_18 ) , .A2( u1_uk_K_r5_40 ) , .ZN( u1_uk_n1113 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U205 (.ZN( u1_K4_24 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1352 ) , .A2( u1_uk_n1393 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U206 (.ZN( u1_K3_24 ) , .A( u1_uk_n1038 ) );
  AOI22_X1 u1_uk_U207 (.B2( u1_uk_K_r1_17 ) , .A2( u1_uk_K_r1_41 ) , .ZN( u1_uk_n1038 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U208 (.ZN( u1_K15_24 ) , .A1( u1_uk_n146 ) , .A2( u1_uk_n1846 ) , .B2( u1_uk_n1864 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U209 (.ZN( u1_K1_30 ) , .A( u1_uk_n1009 ) , .B2( u1_uk_n1213 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U21 (.ZN( u1_uk_n128 ) , .A( u1_uk_n297 ) );
  NAND2_X1 u1_uk_U210 (.A1( u1_key_r_45 ) , .ZN( u1_uk_n1009 ) , .A2( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U211 (.ZN( u1_K9_30 ) , .A( u1_uk_n1161 ) , .B2( u1_uk_n1600 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U212 (.A1( u1_uk_K_r7_29 ) , .ZN( u1_uk_n1161 ) , .A2( u1_uk_n187 ) );
  OAI21_X1 u1_uk_U213 (.ZN( u1_K4_30 ) , .A( u1_uk_n1062 ) , .B2( u1_uk_n1375 ) , .B1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U214 (.A1( u1_uk_K_r2_28 ) , .ZN( u1_uk_n1062 ) , .A2( u1_uk_n230 ) );
  INV_X1 u1_uk_U215 (.ZN( u1_K15_30 ) , .A( u1_uk_n970 ) );
  AOI22_X1 u1_uk_U216 (.B2( u1_uk_K_r13_0 ) , .A2( u1_uk_K_r13_38 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n970 ) );
  OAI22_X1 u1_uk_U217 (.ZN( u1_K3_14 ) , .B2( u1_uk_n1340 ) , .A2( u1_uk_n1347 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n31 ) );
  AOI22_X1 u1_uk_U219 (.B2( u1_uk_K_r2_31 ) , .A2( u1_uk_K_r2_49 ) , .ZN( u1_uk_n1063 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U22 (.ZN( u1_uk_n147 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U220 (.ZN( u1_K1_31 ) , .A2( u1_uk_n1177 ) , .B2( u1_uk_n1181 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U221 (.A( u1_key_r_14 ) , .ZN( u1_uk_n1181 ) );
  OAI22_X1 u1_uk_U222 (.ZN( u1_K16_31 ) , .A2( u1_uk_n1222 ) , .B2( u1_uk_n1225 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U223 (.ZN( u1_K8_31 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1529 ) , .A2( u1_uk_n1567 ) , .B1( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U224 (.ZN( u1_K12_31 ) , .B2( u1_uk_n1715 ) , .B1( u1_uk_n207 ) , .A( u1_uk_n551 ) );
  NAND2_X1 u1_uk_U225 (.A1( u1_uk_K_r10_44 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n551 ) );
  AOI22_X1 u1_uk_U227 (.B2( u1_uk_K_r9_22 ) , .A2( u1_uk_K_r9_30 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n251 ) , .ZN( u1_uk_n437 ) );
  OAI22_X1 u1_uk_U228 (.ZN( u1_K2_31 ) , .B2( u1_uk_n1260 ) , .A2( u1_uk_n1275 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n220 ) );
  INV_X1 u1_uk_U229 (.ZN( u1_K11_39 ) , .A( u1_uk_n460 ) );
  INV_X1 u1_uk_U23 (.ZN( u1_uk_n117 ) , .A( u1_uk_n277 ) );
  AOI22_X1 u1_uk_U230 (.B2( u1_uk_K_r9_30 ) , .A2( u1_uk_K_r9_7 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n292 ) , .ZN( u1_uk_n460 ) );
  AOI22_X1 u1_uk_U232 (.B2( u1_uk_K_r8_44 ) , .A2( u1_uk_K_r8_52 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n209 ) , .ZN( u1_uk_n373 ) );
  OAI22_X1 u1_uk_U233 (.ZN( u1_K13_31 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1772 ) , .A2( u1_uk_n1790 ) , .A1( u1_uk_n207 ) );
  OAI21_X1 u1_uk_U234 (.ZN( u1_K10_31 ) , .B2( u1_uk_n1645 ) , .B1( u1_uk_n298 ) , .A( u1_uk_n342 ) );
  NAND2_X1 u1_uk_U235 (.A1( u1_uk_K_r8_16 ) , .A2( u1_uk_n277 ) , .ZN( u1_uk_n342 ) );
  OAI22_X1 u1_uk_U236 (.ZN( u1_K6_31 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1455 ) , .A2( u1_uk_n1460 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U237 (.ZN( u1_K3_31 ) , .B2( u1_uk_n1333 ) , .A2( u1_uk_n1339 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U238 (.ZN( u1_K5_31 ) , .B1( u1_uk_n100 ) , .A( u1_uk_n1077 ) , .B2( u1_uk_n1401 ) );
  NAND2_X1 u1_uk_U239 (.A1( u1_uk_K_r3_44 ) , .ZN( u1_uk_n1077 ) , .A2( u1_uk_n27 ) );
  INV_X1 u1_uk_U24 (.ZN( u1_uk_n129 ) , .A( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U240 (.ZN( u1_K15_31 ) , .B2( u1_uk_n1843 ) , .A2( u1_uk_n1860 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U241 (.ZN( u1_K1_39 ) , .A( u1_uk_n1014 ) , .B2( u1_uk_n1187 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U242 (.A1( u1_key_r_15 ) , .ZN( u1_uk_n1014 ) , .A2( u1_uk_n155 ) );
  INV_X1 u1_uk_U243 (.A( u1_key_r_22 ) , .ZN( u1_uk_n1187 ) );
  OAI22_X1 u1_uk_U244 (.ZN( u1_K14_31 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1827 ) , .A2( u1_uk_n1833 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U245 (.ZN( u1_K9_31 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1572 ) , .A2( u1_uk_n1613 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U246 (.ZN( u1_K15_39 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1848 ) , .B2( u1_uk_n1866 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U247 (.ZN( u1_K14_39 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1832 ) , .A2( u1_uk_n1836 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U248 (.ZN( u1_K13_39 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1755 ) , .A2( u1_uk_n1774 ) , .B1( u1_uk_n240 ) );
  OAI21_X1 u1_uk_U249 (.ZN( u1_K12_39 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1720 ) , .A( u1_uk_n590 ) );
  INV_X1 u1_uk_U25 (.ZN( u1_uk_n146 ) , .A( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U250 (.A1( u1_uk_K_r10_16 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n590 ) );
  OAI22_X1 u1_uk_U251 (.ZN( u1_K16_48 ) , .B2( u1_uk_n1230 ) , .A2( u1_uk_n1238 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U252 (.ZN( u1_K16_44 ) , .B2( u1_uk_n1246 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n994 ) );
  NAND2_X1 u1_uk_U253 (.A1( u1_uk_K_r14_43 ) , .A2( u1_uk_n94 ) , .ZN( u1_uk_n994 ) );
  OAI21_X1 u1_uk_U254 (.ZN( u1_K8_44 ) , .A( u1_uk_n1144 ) , .B1( u1_uk_n141 ) , .B2( u1_uk_n1568 ) );
  NAND2_X1 u1_uk_U255 (.A1( u1_uk_K_r6_0 ) , .ZN( u1_uk_n1144 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U256 (.ZN( u1_K8_48 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1534 ) , .B2( u1_uk_n1541 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U257 (.ZN( u1_K5_44 ) , .B2( u1_uk_n1419 ) , .A2( u1_uk_n1425 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U258 (.ZN( u1_K5_48 ) , .B2( u1_uk_n1407 ) , .A2( u1_uk_n1414 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U259 (.ZN( u1_K1_48 ) , .A( u1_uk_n1019 ) );
  INV_X1 u1_uk_U26 (.ZN( u1_uk_n145 ) , .A( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U260 (.B2( u1_key_r_21 ) , .A2( u1_key_r_28 ) , .ZN( u1_uk_n1019 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n291 ) );
  INV_X1 u1_uk_U261 (.ZN( u1_K1_44 ) , .A( u1_uk_n1017 ) );
  AOI22_X1 u1_uk_U262 (.B2( u1_key_r_36 ) , .A2( u1_key_r_43 ) , .ZN( u1_uk_n1017 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U263 (.ZN( u1_K15_44 ) , .B2( u1_uk_n1866 ) , .A2( u1_uk_n1884 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U264 (.ZN( u1_K15_48 ) , .B1( u1_uk_n10 ) , .B2( u1_uk_n1854 ) , .A( u1_uk_n975 ) );
  NAND2_X1 u1_uk_U265 (.A1( u1_uk_K_r13_35 ) , .A2( u1_uk_n148 ) , .ZN( u1_uk_n975 ) );
  OAI22_X1 u1_uk_U266 (.ZN( u1_K14_48 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1798 ) , .A2( u1_uk_n1836 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U267 (.ZN( u1_K13_44 ) , .B2( u1_uk_n1754 ) , .A2( u1_uk_n1769 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U268 (.ZN( u1_K13_48 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1785 ) , .A( u1_uk_n947 ) );
  NAND2_X1 u1_uk_U269 (.A1( u1_uk_K_r11_8 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n947 ) );
  INV_X1 u1_uk_U27 (.ZN( u1_uk_n148 ) , .A( u1_uk_n214 ) );
  INV_X1 u1_uk_U270 (.ZN( u1_K12_44 ) , .A( u1_uk_n608 ) );
  AOI22_X1 u1_uk_U271 (.B2( u1_uk_K_r10_37 ) , .A2( u1_uk_K_r10_42 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n271 ) , .ZN( u1_uk_n608 ) );
  OAI22_X1 u1_uk_U272 (.ZN( u1_K12_48 ) , .B2( u1_uk_n1721 ) , .A2( u1_uk_n1730 ) , .B1( u1_uk_n207 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U273 (.ZN( u1_K11_44 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1683 ) , .A2( u1_uk_n1703 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U274 (.ZN( u1_K10_44 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1627 ) , .A2( u1_uk_n1647 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U275 (.ZN( u1_K10_48 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1640 ) , .A2( u1_uk_n1656 ) , .A1( u1_uk_n240 ) );
  INV_X1 u1_uk_U276 (.ZN( u1_K9_48 ) , .A( u1_uk_n1170 ) );
  AOI22_X1 u1_uk_U277 (.B2( u1_uk_K_r7_16 ) , .A2( u1_uk_K_r7_9 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1170 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U278 (.ZN( u1_K7_44 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1489 ) , .A2( u1_uk_n1510 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U279 (.ZN( u1_K7_48 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1501 ) , .A2( u1_uk_n1521 ) , .B1( u1_uk_n291 ) );
  INV_X1 u1_uk_U28 (.A( u1_uk_n202 ) , .ZN( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U280 (.ZN( u1_K6_44 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1458 ) , .A2( u1_uk_n1476 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U281 (.ZN( u1_K6_48 ) , .B2( u1_uk_n1463 ) , .A2( u1_uk_n1470 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U282 (.ZN( u1_K4_44 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1350 ) , .A2( u1_uk_n1367 ) , .B1( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U283 (.ZN( u1_K3_44 ) , .A( u1_uk_n1045 ) , .B2( u1_uk_n1314 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U284 (.A1( u1_uk_K_r1_15 ) , .ZN( u1_uk_n1045 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U285 (.ZN( u1_K3_48 ) , .B2( u1_uk_n1307 ) , .A2( u1_uk_n1342 ) , .A1( u1_uk_n148 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U286 (.ZN( u1_K2_44 ) , .B2( u1_uk_n1281 ) , .A2( u1_uk_n1303 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U287 (.ZN( u1_K16_6 ) , .B2( u1_uk_n1244 ) , .A2( u1_uk_n1249 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U288 (.ZN( u1_K10_6 ) , .B1( u1_uk_n129 ) , .A2( u1_uk_n1621 ) , .B2( u1_uk_n1649 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U289 (.ZN( u1_K8_6 ) , .B2( u1_uk_n1544 ) , .A2( u1_uk_n1549 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n92 ) );
  INV_X1 u1_uk_U29 (.ZN( u1_uk_n10 ) , .A( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U290 (.ZN( u1_K6_6 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1474 ) , .A2( u1_uk_n1478 ) , .A1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U291 (.ZN( u1_K6_8 ) , .A( u1_uk_n1103 ) , .B2( u1_uk_n1446 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U292 (.A1( u1_uk_K_r4_18 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1103 ) );
  OAI21_X1 u1_uk_U293 (.ZN( u1_K5_6 ) , .A( u1_uk_n1086 ) , .B2( u1_uk_n1417 ) , .B1( u1_uk_n93 ) );
  NAND2_X1 u1_uk_U294 (.A1( u1_uk_K_r3_10 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1086 ) );
  OAI21_X1 u1_uk_U295 (.ZN( u1_K4_6 ) , .A( u1_uk_n1069 ) , .B2( u1_uk_n1365 ) , .B1( u1_uk_n83 ) );
  NAND2_X1 u1_uk_U296 (.A1( u1_uk_K_r2_24 ) , .ZN( u1_uk_n1069 ) , .A2( u1_uk_n145 ) );
  OAI22_X1 u1_uk_U297 (.ZN( u1_K2_6 ) , .B2( u1_uk_n1279 ) , .A2( u1_uk_n1300 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U298 (.ZN( u1_K1_8 ) , .A1( u1_uk_n100 ) , .A2( u1_uk_n1176 ) , .B2( u1_uk_n1189 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U299 (.ZN( u1_K15_8 ) , .A( u1_uk_n976 ) );
  INV_X1 u1_uk_U3 (.A( u1_uk_n191 ) , .ZN( u1_uk_n31 ) );
  INV_X1 u1_uk_U30 (.ZN( u1_uk_n17 ) , .A( u1_uk_n214 ) );
  AOI22_X1 u1_uk_U300 (.B2( u1_uk_K_r13_13 ) , .A2( u1_uk_K_r13_17 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n976 ) );
  OAI22_X1 u1_uk_U301 (.ZN( u1_K12_8 ) , .B2( u1_uk_n1731 ) , .A2( u1_uk_n1752 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U302 (.ZN( u1_K8_8 ) , .B2( u1_uk_n1558 ) , .A2( u1_uk_n1564 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n94 ) );
  INV_X1 u1_uk_U303 (.ZN( u1_K7_8 ) , .A( u1_uk_n1126 ) );
  AOI22_X1 u1_uk_U304 (.B2( u1_uk_K_r5_26 ) , .A2( u1_uk_K_r5_4 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1126 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U305 (.ZN( u1_K5_8 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1415 ) , .A2( u1_uk_n1437 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U306 (.ZN( u1_K4_8 ) , .A( u1_uk_n1070 ) );
  AOI22_X1 u1_uk_U307 (.B2( u1_uk_K_r2_41 ) , .A2( u1_uk_K_r2_46 ) , .ZN( u1_uk_n1070 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U308 (.ZN( u1_K3_8 ) , .A2( u1_uk_n1310 ) , .B2( u1_uk_n1326 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U309 (.ZN( u1_K2_8 ) , .A( u1_uk_n1035 ) , .B2( u1_uk_n1270 ) , .B1( u1_uk_n148 ) );
  INV_X1 u1_uk_U31 (.ZN( u1_uk_n11 ) , .A( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U310 (.A1( u1_uk_K_r0_17 ) , .ZN( u1_uk_n1035 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U311 (.ZN( u1_K7_26 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1500 ) , .A2( u1_uk_n1520 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U312 (.ZN( u1_K1_26 ) , .A( u1_uk_n1006 ) );
  AOI22_X1 u1_uk_U313 (.B2( u1_key_r_31 ) , .A2( u1_key_r_51 ) , .ZN( u1_uk_n1006 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U314 (.ZN( u1_K16_8 ) , .A2( u1_uk_n1221 ) , .B2( u1_uk_n1234 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n60 ) );
  INV_X1 u1_uk_U315 (.ZN( u1_K9_26 ) , .A( u1_uk_n1158 ) );
  AOI22_X1 u1_uk_U316 (.B2( u1_uk_K_r7_15 ) , .A2( u1_uk_K_r7_8 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1158 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U317 (.ZN( u1_K4_26 ) , .A( u1_uk_n1058 ) );
  AOI22_X1 u1_uk_U318 (.B2( u1_uk_K_r2_16 ) , .A2( u1_uk_K_r2_7 ) , .ZN( u1_uk_n1058 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n207 ) );
  INV_X1 u1_uk_U319 (.ZN( u1_K15_26 ) , .A( u1_uk_n969 ) );
  INV_X1 u1_uk_U32 (.ZN( u1_uk_n155 ) , .A( u1_uk_n271 ) );
  AOI22_X1 u1_uk_U320 (.B2( u1_uk_K_r13_38 ) , .A2( u1_uk_K_r13_44 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n291 ) , .ZN( u1_uk_n969 ) );
  OAI21_X1 u1_uk_U321 (.ZN( u1_K6_26 ) , .A( u1_uk_n1094 ) , .B2( u1_uk_n1469 ) , .B1( u1_uk_n251 ) );
  NAND2_X1 u1_uk_U322 (.A1( u1_uk_K_r4_35 ) , .ZN( u1_uk_n1094 ) , .A2( u1_uk_n297 ) );
  OAI21_X1 u1_uk_U323 (.ZN( u1_K11_26 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1695 ) , .A( u1_uk_n409 ) );
  NAND2_X1 u1_uk_U324 (.A1( u1_uk_K_r9_35 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n409 ) );
  OAI21_X1 u1_uk_U325 (.ZN( u1_K13_26 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1765 ) , .A( u1_uk_n694 ) );
  NAND2_X1 u1_uk_U326 (.A1( u1_uk_K_r11_7 ) , .A2( u1_uk_n31 ) , .ZN( u1_uk_n694 ) );
  OAI22_X1 u1_uk_U327 (.ZN( u1_K5_26 ) , .A2( u1_uk_n1396 ) , .B2( u1_uk_n1406 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U328 (.ZN( u1_K2_26 ) , .B2( u1_uk_n1289 ) , .A2( u1_uk_n1295 ) , .A1( u1_uk_n214 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U329 (.ZN( u1_K16_26 ) , .B2( u1_uk_n1241 ) , .A2( u1_uk_n1255 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n279 ) );
  INV_X1 u1_uk_U33 (.ZN( u1_uk_n161 ) , .A( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U330 (.ZN( u1_K14_26 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1822 ) , .A2( u1_uk_n1839 ) , .A1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U331 (.ZN( u1_K12_26 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1710 ) , .B2( u1_uk_n1720 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U332 (.ZN( u1_K10_26 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1639 ) , .A2( u1_uk_n1655 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U333 (.ZN( u1_K8_26 ) , .A1( u1_uk_n10 ) , .A2( u1_uk_n1533 ) , .B2( u1_uk_n1540 ) , .B1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U334 (.ZN( u1_K3_26 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1329 ) , .A2( u1_uk_n1345 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U335 (.ZN( u1_K5_46 ) , .B2( u1_uk_n1394 ) , .A1( u1_uk_n141 ) , .A2( u1_uk_n1431 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U336 (.ZN( u1_K15_46 ) , .A2( u1_uk_n1848 ) , .B2( u1_uk_n1875 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U337 (.ZN( u1_K13_46 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1763 ) , .A2( u1_uk_n1775 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U338 (.ZN( u1_K12_46 ) , .B2( u1_uk_n1708 ) , .A2( u1_uk_n1748 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U339 (.ZN( u1_K4_46 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1360 ) , .A2( u1_uk_n1374 ) , .B1( u1_uk_n257 ) );
  INV_X1 u1_uk_U34 (.ZN( u1_uk_n162 ) , .A( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U340 (.ZN( u1_K3_46 ) , .A( u1_uk_n1047 ) , .B2( u1_uk_n1327 ) , .B1( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U341 (.A1( u1_uk_K_r1_22 ) , .ZN( u1_uk_n1047 ) , .A2( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U342 (.ZN( u1_K2_46 ) , .A2( u1_uk_n1266 ) , .B2( u1_uk_n1293 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U343 (.ZN( u1_K1_46 ) , .A( u1_uk_n1018 ) , .B2( u1_uk_n1173 ) , .B1( u1_uk_n17 ) );
  NAND2_X1 u1_uk_U344 (.A1( u1_key_r_49 ) , .ZN( u1_uk_n1018 ) , .A2( u1_uk_n142 ) );
  OAI22_X1 u1_uk_U345 (.ZN( u1_K11_4 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1693 ) , .A2( u1_uk_n1699 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U346 (.ZN( u1_K15_4 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1850 ) , .A2( u1_uk_n1880 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U347 (.ZN( u1_K14_4 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1816 ) , .A2( u1_uk_n1824 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U348 (.ZN( u1_K7_4 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1504 ) , .A2( u1_uk_n1527 ) , .B1( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U349 (.ZN( u1_K1_4 ) , .A( u1_uk_n1020 ) , .B2( u1_uk_n1214 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U35 (.ZN( u1_uk_n187 ) , .A( u1_uk_n213 ) );
  NAND2_X1 u1_uk_U350 (.A1( u1_key_r_3 ) , .ZN( u1_uk_n1020 ) , .A2( u1_uk_n223 ) );
  INV_X1 u1_uk_U351 (.ZN( u1_K6_4 ) , .A( u1_uk_n1101 ) );
  AOI22_X1 u1_uk_U352 (.B2( u1_uk_K_r4_41 ) , .A2( u1_uk_K_r4_47 ) , .ZN( u1_uk_n1101 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n297 ) );
  AOI22_X1 u1_uk_U354 (.B2( u1_uk_K_r2_13 ) , .A2( u1_uk_K_r2_18 ) , .ZN( u1_uk_n1067 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U355 (.ZN( u1_K3_4 ) , .B2( u1_uk_n1323 ) , .A2( u1_uk_n1331 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U356 (.ZN( u1_K2_4 ) , .B2( u1_uk_n1268 ) , .A2( u1_uk_n1297 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U357 (.ZN( u1_K1_40 ) , .B2( u1_uk_n1172 ) , .A2( u1_uk_n1213 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U358 (.ZN( u1_K16_40 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1218 ) , .A2( u1_uk_n1256 ) , .B1( u1_uk_n257 ) );
  BUF_X1 u1_uk_U36 (.Z( u1_uk_n230 ) , .A( u1_uk_n277 ) );
  AOI22_X1 u1_uk_U360 (.B2( u1_uk_K_r10_27 ) , .A2( u1_uk_K_r10_4 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n31 ) , .ZN( u1_uk_n656 ) );
  OAI22_X1 u1_uk_U361 (.ZN( u1_K10_4 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1642 ) , .A2( u1_uk_n1661 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U362 (.ZN( u1_K15_40 ) , .A2( u1_uk_n1847 ) , .B2( u1_uk_n1879 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U363 (.ZN( u1_K13_40 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1774 ) , .A2( u1_uk_n1784 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U364 (.ZN( u1_K6_40 ) , .A2( u1_uk_n1442 ) , .B2( u1_uk_n1450 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n240 ) );
  AOI22_X1 u1_uk_U366 (.B2( u1_uk_K_r9_45 ) , .A2( u1_uk_K_r9_9 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n292 ) , .ZN( u1_uk_n468 ) );
  OAI21_X1 u1_uk_U367 (.ZN( u1_K9_46 ) , .B1( u1_uk_n11 ) , .A( u1_uk_n1169 ) , .B2( u1_uk_n1607 ) );
  NAND2_X1 u1_uk_U368 (.A1( u1_uk_K_r7_37 ) , .ZN( u1_uk_n1169 ) , .A2( u1_uk_n31 ) );
  BUF_X1 u1_uk_U37 (.Z( u1_uk_n213 ) , .A( u1_uk_n286 ) );
  AOI22_X1 u1_uk_U370 (.B2( u1_uk_K_r5_23 ) , .A2( u1_uk_K_r5_31 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1124 ) , .B1( u1_uk_n208 ) );
  AOI22_X1 u1_uk_U372 (.A2( u1_uk_K_r8_2 ) , .B2( u1_uk_K_r8_22 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n250 ) , .ZN( u1_uk_n375 ) );
  OAI22_X1 u1_uk_U373 (.ZN( u1_K11_40 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1664 ) , .B2( u1_uk_n1672 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U374 (.ZN( u1_K8_40 ) , .B2( u1_uk_n1555 ) , .A2( u1_uk_n1561 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U375 (.ZN( u1_K7_40 ) , .A2( u1_uk_n1482 ) , .B2( u1_uk_n1494 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U376 (.ZN( u1_K4_40 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1372 ) , .A2( u1_uk_n1382 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U377 (.ZN( u1_K2_40 ) , .A2( u1_uk_n1265 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1296 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U378 (.ZN( u1_K15_33 ) , .B2( u1_uk_n1870 ) , .B1( u1_uk_n83 ) , .A( u1_uk_n972 ) );
  NAND2_X1 u1_uk_U379 (.A1( u1_uk_K_r13_31 ) , .A2( u1_uk_n60 ) , .ZN( u1_uk_n972 ) );
  BUF_X1 u1_uk_U38 (.Z( u1_uk_n208 ) , .A( u1_uk_n291 ) );
  OAI21_X1 u1_uk_U380 (.ZN( u1_K2_33 ) , .A( u1_uk_n1030 ) , .B2( u1_uk_n1288 ) , .B1( u1_uk_n223 ) );
  NAND2_X1 u1_uk_U381 (.A1( u1_uk_K_r0_31 ) , .ZN( u1_uk_n1030 ) , .A2( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U382 (.ZN( u1_K1_28 ) , .B2( u1_uk_n1173 ) , .A2( u1_uk_n1178 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n238 ) );
  INV_X1 u1_uk_U383 (.A( u1_key_r_8 ) , .ZN( u1_uk_n1178 ) );
  OAI22_X1 u1_uk_U384 (.ZN( u1_K14_28 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1821 ) , .A2( u1_uk_n1827 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U385 (.ZN( u1_K11_28 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1672 ) , .A2( u1_uk_n1704 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U386 (.ZN( u1_K6_28 ) , .B2( u1_uk_n1450 ) , .A2( u1_uk_n1477 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U387 (.ZN( u1_K3_28 ) , .B2( u1_uk_n1328 ) , .A2( u1_uk_n1333 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U388 (.ZN( u1_K5_33 ) , .A( u1_uk_n1078 ) , .B2( u1_uk_n1431 ) , .B1( u1_uk_n214 ) );
  NAND2_X1 u1_uk_U389 (.A1( u1_uk_K_r3_14 ) , .ZN( u1_uk_n1078 ) , .A2( u1_uk_n252 ) );
  BUF_X1 u1_uk_U39 (.Z( u1_uk_n202 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U390 (.ZN( u1_K15_28 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1855 ) , .A2( u1_uk_n1883 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U391 (.ZN( u1_K12_28 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1710 ) , .A2( u1_uk_n1714 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U392 (.ZN( u1_K10_28 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1640 ) , .A2( u1_uk_n1647 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U393 (.ZN( u1_K9_28 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1607 ) , .A2( u1_uk_n1614 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U394 (.ZN( u1_K7_28 ) , .B2( u1_uk_n1501 ) , .A2( u1_uk_n1510 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U395 (.ZN( u1_K5_28 ) , .B2( u1_uk_n1396 ) , .A2( u1_uk_n1400 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U396 (.ZN( u1_K14_1 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1808 ) , .A2( u1_uk_n1813 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U397 (.ZN( u1_K11_1 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1688 ) , .A2( u1_uk_n1705 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U398 (.ZN( u1_K3_1 ) , .B2( u1_uk_n1315 ) , .A2( u1_uk_n1320 ) , .A1( u1_uk_n279 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U399 (.ZN( u1_K2_1 ) , .B2( u1_uk_n1284 ) , .A2( u1_uk_n1305 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U4 (.ZN( u1_uk_n164 ) , .A( u1_uk_n203 ) );
  BUF_X1 u1_uk_U40 (.Z( u1_uk_n209 ) , .A( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U400 (.ZN( u1_K7_1 ) , .A( u1_uk_n1108 ) , .B2( u1_uk_n1492 ) , .B1( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U401 (.A1( u1_uk_K_r5_10 ) , .ZN( u1_uk_n1108 ) , .A2( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U402 (.ZN( u1_K5_1 ) , .B2( u1_uk_n1422 ) , .A2( u1_uk_n1429 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U403 (.ZN( u1_K1_9 ) , .B2( u1_uk_n1209 ) , .A2( u1_uk_n1215 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U404 (.ZN( u1_K13_16 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1761 ) , .A2( u1_uk_n1766 ) , .B1( u1_uk_n202 ) );
  OAI21_X1 u1_uk_U405 (.ZN( u1_K10_16 ) , .B2( u1_uk_n1660 ) , .B1( u1_uk_n286 ) , .A( u1_uk_n305 ) );
  NAND2_X1 u1_uk_U406 (.A1( u1_uk_K_r8_32 ) , .A2( u1_uk_n203 ) , .ZN( u1_uk_n305 ) );
  OAI22_X1 u1_uk_U407 (.ZN( u1_K9_16 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1578 ) , .A2( u1_uk_n1585 ) , .B1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U408 (.ZN( u1_K8_16 ) , .B2( u1_uk_n1536 ) , .A2( u1_uk_n1544 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U409 (.ZN( u1_K7_16 ) , .A( u1_uk_n1107 ) , .B2( u1_uk_n1526 ) , .B1( u1_uk_n161 ) );
  BUF_X1 u1_uk_U41 (.Z( u1_uk_n203 ) , .A( u1_uk_n291 ) );
  NAND2_X1 u1_uk_U410 (.A1( u1_uk_K_r5_32 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1107 ) );
  OAI22_X1 u1_uk_U411 (.ZN( u1_K6_16 ) , .B2( u1_uk_n1466 ) , .A2( u1_uk_n1472 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U412 (.ZN( u1_K4_16 ) , .B2( u1_uk_n1359 ) , .A2( u1_uk_n1363 ) , .B1( u1_uk_n145 ) , .A1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U413 (.ZN( u1_K3_16 ) , .A( u1_uk_n1036 ) , .B2( u1_uk_n1348 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U414 (.A1( u1_uk_K_r1_6 ) , .ZN( u1_uk_n1036 ) , .A2( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U415 (.ZN( u1_K1_16 ) , .B2( u1_uk_n1192 ) , .A2( u1_uk_n1198 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U416 (.ZN( u1_K15_9 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1873 ) , .A( u1_uk_n977 ) );
  NAND2_X1 u1_uk_U417 (.A1( u1_uk_K_r13_4 ) , .A2( u1_uk_n63 ) , .ZN( u1_uk_n977 ) );
  OAI21_X1 u1_uk_U418 (.ZN( u1_K14_9 ) , .B2( u1_uk_n1818 ) , .B1( u1_uk_n83 ) , .A( u1_uk_n963 ) );
  NAND2_X1 u1_uk_U419 (.A1( u1_uk_K_r12_18 ) , .ZN( u1_uk_n963 ) , .A2( u1_uk_n99 ) );
  BUF_X1 u1_uk_U42 (.Z( u1_uk_n242 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U420 (.ZN( u1_K13_9 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1761 ) , .A2( u1_uk_n1773 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U421 (.ZN( u1_K12_9 ) , .A1( u1_uk_n10 ) , .B2( u1_uk_n1745 ) , .A2( u1_uk_n1752 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U422 (.ZN( u1_K11_9 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1663 ) , .A2( u1_uk_n1693 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U423 (.ZN( u1_K8_9 ) , .A1( u1_uk_n109 ) , .A2( u1_uk_n1532 ) , .B2( u1_uk_n1538 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U424 (.ZN( u1_K5_9 ) , .B2( u1_uk_n1427 ) , .A2( u1_uk_n1437 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U425 (.ZN( u1_K4_9 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1359 ) , .A2( u1_uk_n1369 ) , .B1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U426 (.ZN( u1_K3_9 ) , .A( u1_uk_n1049 ) , .B2( u1_uk_n1325 ) , .B1( u1_uk_n277 ) );
  NAND2_X1 u1_uk_U427 (.A1( u1_uk_K_r1_18 ) , .ZN( u1_uk_n1049 ) , .A2( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U428 (.ZN( u1_K2_9 ) , .A2( u1_uk_n1262 ) , .B2( u1_uk_n1291 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U429 (.ZN( u1_K16_9 ) , .B2( u1_uk_n1251 ) , .A2( u1_uk_n1258 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n60 ) );
  BUF_X1 u1_uk_U43 (.Z( u1_uk_n220 ) , .A( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U430 (.ZN( u1_K12_33 ) , .B2( u1_uk_n1748 ) , .A( u1_uk_n586 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U431 (.A1( u1_uk_K_r10_14 ) , .A2( u1_uk_n117 ) , .ZN( u1_uk_n586 ) );
  OAI22_X1 u1_uk_U432 (.ZN( u1_K16_16 ) , .B2( u1_uk_n1237 ) , .A2( u1_uk_n1244 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U433 (.ZN( u1_K15_16 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1859 ) , .A2( u1_uk_n1874 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U434 (.ZN( u1_K5_16 ) , .B1( u1_uk_n129 ) , .A2( u1_uk_n1397 ) , .B2( u1_uk_n1410 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U435 (.ZN( u1_K2_16 ) , .B2( u1_uk_n1274 ) , .A2( u1_uk_n1292 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U436 (.ZN( u1_K2_28 ) , .A( u1_uk_n1028 ) );
  AOI22_X1 u1_uk_U437 (.B2( u1_uk_K_r0_15 ) , .A2( u1_uk_K_r0_49 ) , .ZN( u1_uk_n1028 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U438 (.ZN( u1_K14_37 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1815 ) , .A2( u1_uk_n1821 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U439 (.ZN( u1_K5_37 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1395 ) , .A2( u1_uk_n1433 ) , .B1( u1_uk_n257 ) );
  BUF_X1 u1_uk_U44 (.Z( u1_uk_n214 ) , .A( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U440 (.ZN( u1_K4_37 ) , .B2( u1_uk_n1361 ) , .A2( u1_uk_n1375 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n209 ) );
  AOI22_X1 u1_uk_U442 (.B2( u1_uk_K_r8_28 ) , .A2( u1_uk_K_r8_52 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n208 ) , .ZN( u1_uk_n366 ) );
  INV_X1 u1_uk_U443 (.ZN( u1_K8_37 ) , .A( u1_uk_n1138 ) );
  AOI22_X1 u1_uk_U444 (.B2( u1_uk_K_r6_14 ) , .A2( u1_uk_K_r6_7 ) , .ZN( u1_uk_n1138 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n203 ) );
  AOI22_X1 u1_uk_U446 (.B2( u1_uk_K_r8_17 ) , .A2( u1_uk_K_r8_27 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n297 ) , .ZN( u1_uk_n376 ) );
  INV_X1 u1_uk_U447 (.ZN( u1_K9_9 ) , .A( u1_uk_n1171 ) );
  AOI22_X1 u1_uk_U448 (.B2( u1_uk_K_r7_13 ) , .A1( u1_uk_K_r7_6 ) , .ZN( u1_uk_n1171 ) , .A2( u1_uk_n148 ) , .B1( u1_uk_n207 ) );
  BUF_X1 u1_uk_U45 (.Z( u1_uk_n240 ) , .A( u1_uk_n271 ) );
  AOI22_X1 u1_uk_U450 (.B2( u1_uk_K_r4_3 ) , .A2( u1_uk_K_r4_41 ) , .ZN( u1_uk_n1104 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U451 (.ZN( u1_K7_9 ) , .B2( u1_uk_n1491 ) , .A2( u1_uk_n1498 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U452 (.ZN( u1_K15_1 ) , .B2( u1_uk_n1868 ) , .A2( u1_uk_n1887 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n99 ) );
  INV_X1 u1_uk_U453 (.ZN( u1_K16_37 ) , .A( u1_uk_n989 ) );
  AOI22_X1 u1_uk_U454 (.B2( u1_uk_K_r14_2 ) , .A2( u1_uk_K_r14_50 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n989 ) );
  OAI22_X1 u1_uk_U455 (.ZN( u1_K16_33 ) , .B2( u1_uk_n1250 ) , .A2( u1_uk_n1255 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U456 (.ZN( u1_K14_33 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1815 ) , .A2( u1_uk_n1833 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U457 (.ZN( u1_K13_33 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1753 ) , .A2( u1_uk_n1758 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U458 (.ZN( u1_K11_33 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1683 ) , .A2( u1_uk_n1689 ) , .B1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U459 (.ZN( u1_K7_33 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1494 ) , .A2( u1_uk_n1514 ) , .B1( u1_uk_n279 ) );
  BUF_X1 u1_uk_U46 (.Z( u1_uk_n238 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U460 (.ZN( u1_K3_33 ) , .B2( u1_uk_n1322 ) , .A2( u1_uk_n1339 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n203 ) );
  AOI22_X1 u1_uk_U462 (.B2( u1_uk_K_r7_1 ) , .A2( u1_uk_K_r7_8 ) , .ZN( u1_uk_n1162 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n286 ) );
  AOI22_X1 u1_uk_U464 (.B2( u1_uk_K_r8_22 ) , .A2( u1_uk_K_r8_42 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n297 ) , .ZN( u1_uk_n349 ) );
  AOI22_X1 u1_uk_U466 (.B2( u1_key_r_44 ) , .A2( u1_key_r_51 ) , .ZN( u1_uk_n1011 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U467 (.ZN( u1_K8_33 ) , .B2( u1_uk_n1528 ) , .A2( u1_uk_n1533 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U468 (.ZN( u1_K6_33 ) , .B2( u1_uk_n1458 ) , .A2( u1_uk_n1463 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U469 (.ZN( u1_K4_33 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1349 ) , .A2( u1_uk_n1356 ) , .A1( u1_uk_n250 ) );
  BUF_X1 u1_uk_U47 (.Z( u1_uk_n217 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U470 (.ZN( u1_K15_37 ) , .A2( u1_uk_n1849 ) , .B2( u1_uk_n1876 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U471 (.ZN( u1_K13_37 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1764 ) , .A2( u1_uk_n1776 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U472 (.ZN( u1_K12_37 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1709 ) , .A2( u1_uk_n1749 ) , .A1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U473 (.ZN( u1_K11_37 ) , .B2( u1_uk_n1694 ) , .A( u1_uk_n456 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U474 (.A1( u1_uk_K_r9_38 ) , .ZN( u1_uk_n456 ) , .A2( u1_uk_n63 ) );
  OAI21_X1 u1_uk_U475 (.ZN( u1_K9_37 ) , .A( u1_uk_n1164 ) , .B2( u1_uk_n1581 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U476 (.A1( u1_uk_K_r7_7 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n1164 ) );
  OAI21_X1 u1_uk_U477 (.ZN( u1_K6_37 ) , .A( u1_uk_n1098 ) , .B2( u1_uk_n1468 ) , .B1( u1_uk_n271 ) );
  NAND2_X1 u1_uk_U478 (.A1( u1_uk_K_r4_38 ) , .ZN( u1_uk_n1098 ) , .A2( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U479 (.ZN( u1_K3_37 ) , .B2( u1_uk_n1322 ) , .A2( u1_uk_n1328 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n94 ) );
  BUF_X1 u1_uk_U48 (.Z( u1_uk_n223 ) , .A( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U480 (.ZN( u1_K1_29 ) , .B2( u1_uk_n1182 ) , .A2( u1_uk_n1188 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U481 (.ZN( u1_K10_36 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1619 ) , .A( u1_uk_n363 ) );
  NAND2_X1 u1_uk_U482 (.A1( u1_uk_K_r8_21 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n363 ) );
  OAI21_X1 u1_uk_U483 (.ZN( u1_K14_29 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1837 ) , .A( u1_uk_n954 ) );
  NAND2_X1 u1_uk_U484 (.A1( u1_uk_K_r12_44 ) , .A2( u1_uk_n164 ) , .ZN( u1_uk_n954 ) );
  OAI22_X1 u1_uk_U485 (.ZN( u1_K13_29 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1772 ) , .A2( u1_uk_n1775 ) , .B1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U486 (.ZN( u1_K11_29 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1664 ) , .A( u1_uk_n415 ) );
  NAND2_X1 u1_uk_U487 (.A1( u1_uk_K_r9_0 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n415 ) );
  OAI21_X1 u1_uk_U488 (.ZN( u1_K3_29 ) , .A( u1_uk_n1040 ) , .B2( u1_uk_n1343 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U489 (.A1( u1_uk_K_r1_44 ) , .ZN( u1_uk_n1040 ) , .A2( u1_uk_n294 ) );
  BUF_X1 u1_uk_U49 (.Z( u1_uk_n231 ) , .A( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U490 (.ZN( u1_K2_29 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1267 ) , .B2( u1_uk_n1282 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U491 (.ZN( u1_K15_29 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1849 ) , .B2( u1_uk_n1867 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U492 (.ZN( u1_K10_29 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1627 ) , .A2( u1_uk_n1655 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U493 (.ZN( u1_K9_29 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1595 ) , .A2( u1_uk_n1599 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U494 (.ZN( u1_K5_29 ) , .B2( u1_uk_n1407 ) , .A1( u1_uk_n142 ) , .A2( u1_uk_n1426 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U495 (.ZN( u1_K16_29 ) , .A( u1_uk_n985 ) );
  AOI22_X1 u1_uk_U496 (.B2( u1_uk_K_r14_16 ) , .A2( u1_uk_K_r14_23 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n277 ) , .ZN( u1_uk_n985 ) );
  INV_X1 u1_uk_U497 (.ZN( u1_K8_29 ) , .A( u1_uk_n1134 ) );
  AOI22_X1 u1_uk_U498 (.B2( u1_uk_K_r6_28 ) , .A2( u1_uk_K_r6_35 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1134 ) , .B1( u1_uk_n230 ) );
  OAI21_X1 u1_uk_U499 (.ZN( u1_K6_29 ) , .A( u1_uk_n1095 ) , .B2( u1_uk_n1442 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U5 (.ZN( u1_uk_n163 ) , .A( u1_uk_n202 ) );
  BUF_X1 u1_uk_U50 (.Z( u1_uk_n191 ) , .A( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U500 (.A1( u1_uk_K_r4_0 ) , .ZN( u1_uk_n1095 ) , .A2( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U502 (.B2( u1_uk_K_r2_31 ) , .A2( u1_uk_K_r2_36 ) , .ZN( u1_uk_n1060 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U503 (.ZN( u1_K12_29 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1721 ) , .A2( u1_uk_n1744 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U504 (.ZN( u1_K7_29 ) , .B2( u1_uk_n1489 ) , .A2( u1_uk_n1520 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U505 (.ZN( u1_K14_2 ) , .A1( u1_uk_n182 ) , .B2( u1_uk_n1824 ) , .A2( u1_uk_n1831 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U506 (.ZN( u1_K11_2 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1673 ) , .A2( u1_uk_n1707 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U507 (.ZN( u1_K3_2 ) , .B2( u1_uk_n1331 ) , .A2( u1_uk_n1336 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U508 (.ZN( u1_K2_2 ) , .B2( u1_uk_n1273 ) , .A2( u1_uk_n1305 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U509 (.ZN( u1_K8_2 ) , .A( u1_uk_n1135 ) , .B2( u1_uk_n1545 ) , .B1( u1_uk_n155 ) );
  BUF_X1 u1_uk_U51 (.Z( u1_uk_n207 ) , .A( u1_uk_n291 ) );
  NAND2_X1 u1_uk_U510 (.A1( u1_uk_K_r6_27 ) , .ZN( u1_uk_n1135 ) , .A2( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U511 (.ZN( u1_K7_2 ) , .A( u1_uk_n1116 ) , .B2( u1_uk_n1484 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U512 (.A1( u1_uk_K_r5_41 ) , .ZN( u1_uk_n1116 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U513 (.ZN( u1_K5_2 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1397 ) , .B2( u1_uk_n1402 ) , .B1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U514 (.ZN( u1_K9_12 ) , .A( u1_uk_n1149 ) , .B2( u1_uk_n1573 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U515 (.A1( u1_uk_K_r7_53 ) , .ZN( u1_uk_n1149 ) , .A2( u1_uk_n142 ) );
  OAI21_X1 u1_uk_U516 (.ZN( u1_K1_12 ) , .B2( u1_uk_n1184 ) , .B1( u1_uk_n148 ) , .A( u1_uk_n998 ) );
  NAND2_X1 u1_uk_U517 (.A1( u1_key_r_12 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n998 ) );
  OAI21_X1 u1_uk_U518 (.ZN( u1_K13_17 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1773 ) , .A( u1_uk_n681 ) );
  NAND2_X1 u1_uk_U519 (.A1( u1_uk_K_r11_27 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n681 ) );
  BUF_X1 u1_uk_U52 (.Z( u1_uk_n222 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U520 (.ZN( u1_K10_17 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1626 ) , .A2( u1_uk_n1654 ) , .B1( u1_uk_n251 ) );
  OAI21_X1 u1_uk_U521 (.ZN( u1_K9_17 ) , .B1( u1_uk_n10 ) , .A( u1_uk_n1152 ) , .B2( u1_uk_n1598 ) );
  NAND2_X1 u1_uk_U522 (.A1( u1_uk_K_r7_26 ) , .ZN( u1_uk_n1152 ) , .A2( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U523 (.ZN( u1_K8_17 ) , .A( u1_uk_n1131 ) , .B2( u1_uk_n1552 ) , .B1( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U524 (.A1( u1_uk_K_r6_26 ) , .ZN( u1_uk_n1131 ) , .A2( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U525 (.ZN( u1_K7_17 ) , .B2( u1_uk_n1488 ) , .A2( u1_uk_n1518 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U526 (.ZN( u1_K4_17 ) , .A( u1_uk_n1051 ) , .B2( u1_uk_n1369 ) , .B1( u1_uk_n292 ) );
  NAND2_X1 u1_uk_U527 (.A1( u1_uk_K_r2_27 ) , .ZN( u1_uk_n1051 ) , .A2( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U528 (.ZN( u1_K3_17 ) , .B2( u1_uk_n1317 ) , .A2( u1_uk_n1340 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U529 (.ZN( u1_K15_12 ) , .A1( u1_uk_n147 ) , .A2( u1_uk_n1845 ) , .B2( u1_uk_n1863 ) , .B1( u1_uk_n240 ) );
  BUF_X1 u1_uk_U53 (.Z( u1_uk_n188 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U530 (.ZN( u1_K14_12 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1831 ) , .A2( u1_uk_n1835 ) , .B1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U531 (.ZN( u1_K12_12 ) , .B2( u1_uk_n1719 ) , .A( u1_uk_n503 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U532 (.A1( u1_uk_K_r10_11 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n503 ) );
  OAI22_X1 u1_uk_U533 (.ZN( u1_K15_2 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1858 ) , .A2( u1_uk_n1887 ) , .B1( u1_uk_n213 ) );
  INV_X1 u1_uk_U534 (.ZN( u1_K12_17 ) , .A( u1_uk_n509 ) );
  AOI22_X1 u1_uk_U535 (.B2( u1_uk_K_r10_18 ) , .A2( u1_uk_K_r10_41 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n257 ) , .ZN( u1_uk_n509 ) );
  AOI22_X1 u1_uk_U537 (.B2( u1_uk_K_r9_4 ) , .A2( u1_uk_K_r9_55 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n188 ) , .ZN( u1_uk_n385 ) );
  INV_X1 u1_uk_U538 (.ZN( u1_K7_12 ) , .A( u1_uk_n1105 ) );
  AOI22_X1 u1_uk_U539 (.B2( u1_uk_K_r5_17 ) , .A2( u1_uk_K_r5_39 ) , .ZN( u1_uk_n1105 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n242 ) );
  BUF_X1 u1_uk_U54 (.Z( u1_uk_n250 ) , .A( u1_uk_n257 ) );
  OAI21_X1 u1_uk_U540 (.ZN( u1_K5_12 ) , .A( u1_uk_n1071 ) , .B2( u1_uk_n1405 ) , .B1( u1_uk_n230 ) );
  NAND2_X1 u1_uk_U541 (.A1( u1_uk_K_r3_11 ) , .ZN( u1_uk_n1071 ) , .A2( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U542 (.ZN( u1_K4_12 ) , .B2( u1_uk_n1371 ) , .A2( u1_uk_n1391 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U543 (.ZN( u1_K3_12 ) , .B2( u1_uk_n1336 ) , .A2( u1_uk_n1341 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U544 (.ZN( u1_K2_12 ) , .A2( u1_uk_n1263 ) , .B2( u1_uk_n1278 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U545 (.ZN( u1_K1_36 ) , .B2( u1_uk_n1188 ) , .A2( u1_uk_n1195 ) , .A1( u1_uk_n148 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U546 (.ZN( u1_K16_12 ) , .B2( u1_uk_n1228 ) , .B1( u1_uk_n223 ) , .A( u1_uk_n979 ) );
  NAND2_X1 u1_uk_U547 (.A1( u1_uk_K_r14_12 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n979 ) );
  OAI21_X1 u1_uk_U548 (.ZN( u1_K16_17 ) , .B2( u1_uk_n1227 ) , .B1( u1_uk_n202 ) , .A( u1_uk_n982 ) );
  NAND2_X1 u1_uk_U549 (.A1( u1_uk_K_r14_10 ) , .A2( u1_uk_n257 ) , .ZN( u1_uk_n982 ) );
  BUF_X1 u1_uk_U55 (.Z( u1_uk_n251 ) , .A( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U550 (.ZN( u1_K9_36 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1599 ) , .A2( u1_uk_n1605 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U551 (.ZN( u1_K15_17 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1844 ) , .B2( u1_uk_n1862 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U552 (.ZN( u1_K14_17 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1810 ) , .A2( u1_uk_n1834 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U553 (.ZN( u1_K5_17 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1404 ) , .A2( u1_uk_n1424 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U554 (.ZN( u1_K6_17 ) , .A( u1_uk_n1089 ) );
  AOI22_X1 u1_uk_U555 (.B2( u1_uk_K_r4_4 ) , .A2( u1_uk_K_r4_55 ) , .ZN( u1_uk_n1089 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U556 (.ZN( u1_K15_36 ) , .B2( u1_uk_n1856 ) , .A2( u1_uk_n1870 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U557 (.ZN( u1_K14_36 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1800 ) , .A2( u1_uk_n1838 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U558 (.ZN( u1_K13_36 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1777 ) , .A2( u1_uk_n1783 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U559 (.ZN( u1_K3_36 ) , .B2( u1_uk_n1309 ) , .A2( u1_uk_n1344 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n203 ) );
  BUF_X1 u1_uk_U56 (.A( u1_uk_n251 ) , .Z( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U560 (.ZN( u1_K2_36 ) , .B2( u1_uk_n1272 ) , .A2( u1_uk_n1288 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U561 (.ZN( u1_K1_38 ) , .B2( u1_uk_n1195 ) , .A2( u1_uk_n1201 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U562 (.ZN( u1_K16_36 ) , .B2( u1_uk_n1233 ) , .A2( u1_uk_n1240 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U563 (.ZN( u1_K12_38 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1708 ) , .A2( u1_uk_n1735 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U564 (.ZN( u1_K11_38 ) , .B2( u1_uk_n1670 ) , .A2( u1_uk_n1678 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U565 (.ZN( u1_K9_38 ) , .B2( u1_uk_n1605 ) , .A2( u1_uk_n1612 ) , .B1( u1_uk_n214 ) , .A1( u1_uk_n92 ) );
  INV_X1 u1_uk_U566 (.ZN( u1_K7_36 ) , .A( u1_uk_n1121 ) );
  AOI22_X1 u1_uk_U567 (.B2( u1_uk_K_r5_1 ) , .A2( u1_uk_K_r5_21 ) , .ZN( u1_uk_n1121 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n220 ) );
  INV_X1 u1_uk_U568 (.ZN( u1_K11_36 ) , .A( u1_uk_n454 ) );
  AOI22_X1 u1_uk_U569 (.B2( u1_uk_K_r9_15 ) , .A2( u1_uk_K_r9_7 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n202 ) , .ZN( u1_uk_n454 ) );
  BUF_X1 u1_uk_U57 (.Z( u1_uk_n286 ) , .A( u1_uk_n294 ) );
  INV_X1 u1_uk_U570 (.ZN( u1_K5_36 ) , .A( u1_uk_n1080 ) );
  AOI22_X1 u1_uk_U571 (.B2( u1_uk_K_r3_29 ) , .A2( u1_uk_K_r3_52 ) , .ZN( u1_uk_n1080 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U572 (.ZN( u1_K15_38 ) , .A( u1_uk_n973 ) );
  AOI22_X1 u1_uk_U573 (.B2( u1_uk_K_r13_23 ) , .A2( u1_uk_K_r13_44 ) , .A1( u1_uk_n110 ) , .B1( u1_uk_n220 ) , .ZN( u1_uk_n973 ) );
  AOI22_X1 u1_uk_U575 (.B2( u1_uk_K_r8_28 ) , .A2( u1_uk_K_r8_8 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n369 ) );
  OAI22_X1 u1_uk_U576 (.ZN( u1_K8_36 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1554 ) , .A2( u1_uk_n1560 ) , .A1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U577 (.ZN( u1_K6_38 ) , .B2( u1_uk_n1448 ) , .B1( u1_uk_n145 ) , .A2( u1_uk_n1455 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U578 (.ZN( u1_K5_38 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1394 ) , .A2( u1_uk_n1418 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U579 (.ZN( u1_K16_10 ) , .B2( u1_uk_n1249 ) , .A2( u1_uk_n1252 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n83 ) );
  BUF_X1 u1_uk_U58 (.Z( u1_uk_n291 ) , .A( u1_uk_n294 ) );
  OAI21_X1 u1_uk_U580 (.ZN( u1_K15_10 ) , .B2( u1_uk_n1869 ) , .B1( u1_uk_n94 ) , .A( u1_uk_n964 ) );
  NAND2_X1 u1_uk_U581 (.A1( u1_uk_K_r13_55 ) , .A2( u1_uk_n92 ) , .ZN( u1_uk_n964 ) );
  OAI22_X1 u1_uk_U582 (.ZN( u1_K14_10 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1809 ) , .A2( u1_uk_n1814 ) , .B1( u1_uk_n213 ) );
  OAI21_X1 u1_uk_U583 (.ZN( u1_K11_10 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1663 ) , .A( u1_uk_n377 ) );
  NAND2_X1 u1_uk_U584 (.A1( u1_uk_K_r9_54 ) , .A2( u1_uk_n17 ) , .ZN( u1_uk_n377 ) );
  OAI22_X1 u1_uk_U585 (.ZN( u1_K10_10 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1625 ) , .A2( u1_uk_n1653 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U586 (.ZN( u1_K5_10 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1403 ) , .A2( u1_uk_n1423 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U587 (.ZN( u1_K9_10 ) , .A( u1_uk_n1147 ) );
  AOI22_X1 u1_uk_U588 (.B1( n116 ) , .B2( u1_uk_K_r7_25 ) , .A2( u1_uk_K_r7_32 ) , .ZN( u1_uk_n1147 ) , .A1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U589 (.ZN( u1_K8_10 ) , .B2( u1_uk_n1549 ) , .A2( u1_uk_n1551 ) , .A1( u1_uk_n277 ) , .B1( u1_uk_n92 ) );
  BUF_X1 u1_uk_U59 (.Z( u1_uk_n279 ) , .A( u1_uk_n297 ) );
  AOI22_X1 u1_uk_U591 (.B2( u1_uk_K_r4_3 ) , .A2( u1_uk_K_r4_54 ) , .ZN( u1_uk_n1088 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n208 ) );
  AOI22_X1 u1_uk_U593 (.B2( u1_uk_K_r2_26 ) , .A2( u1_uk_K_r2_6 ) , .ZN( u1_uk_n1050 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U594 (.ZN( u1_K1_10 ) , .A( u1_uk_n996 ) );
  AOI22_X1 u1_uk_U595 (.B2( u1_key_r_41 ) , .A2( u1_key_r_48 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n298 ) , .ZN( u1_uk_n996 ) );
  OAI22_X1 u1_uk_U596 (.ZN( u1_K16_22 ) , .B2( u1_uk_n1235 ) , .A2( u1_uk_n1242 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U597 (.ZN( u1_K12_22 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1722 ) , .A2( u1_uk_n1732 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U598 (.ZN( u1_K3_22 ) , .B2( u1_uk_n1311 ) , .A2( u1_uk_n1346 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n191 ) );
  INV_X1 u1_uk_U599 (.ZN( u1_K13_22 ) , .A( u1_uk_n692 ) );
  INV_X1 u1_uk_U6 (.ZN( u1_uk_n182 ) , .A( u1_uk_n223 ) );
  BUF_X1 u1_uk_U60 (.Z( u1_uk_n271 ) , .A( u1_uk_n297 ) );
  AOI22_X1 u1_uk_U600 (.B2( u1_uk_K_r11_10 ) , .A2( u1_uk_K_r11_47 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n238 ) , .ZN( u1_uk_n692 ) );
  AOI22_X1 u1_uk_U602 (.B2( u1_uk_K_r9_13 ) , .A2( u1_uk_K_r9_19 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n230 ) , .ZN( u1_uk_n407 ) );
  AOI22_X1 u1_uk_U604 (.B2( u1_uk_K_r8_27 ) , .A2( u1_uk_K_r8_5 ) , .B1( u1_uk_n148 ) , .A1( u1_uk_n279 ) , .ZN( u1_uk_n312 ) );
  INV_X1 u1_uk_U605 (.ZN( u1_K9_22 ) , .A( u1_uk_n1157 ) );
  AOI22_X1 u1_uk_U606 (.B2( u1_uk_K_r7_41 ) , .A2( u1_uk_K_r7_48 ) , .ZN( u1_uk_n1157 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U607 (.ZN( u1_K8_22 ) , .B2( u1_uk_n1559 ) , .A2( u1_uk_n1565 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n60 ) );
  AOI22_X1 u1_uk_U609 (.B2( u1_uk_K_r3_24 ) , .A2( u1_uk_K_r3_33 ) , .ZN( u1_uk_n1074 ) , .B1( u1_uk_n222 ) , .A1( u1_uk_n31 ) );
  BUF_X1 u1_uk_U61 (.Z( u1_uk_n277 ) , .A( u1_uk_n297 ) );
  INV_X1 u1_uk_U610 (.ZN( u1_K1_22 ) , .A( u1_uk_n1004 ) );
  AOI22_X1 u1_uk_U611 (.B2( u1_key_r_25 ) , .A2( u1_key_r_32 ) , .ZN( u1_uk_n1004 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U612 (.ZN( u1_K16_35 ) , .B2( u1_uk_n1238 ) , .A2( u1_uk_n1245 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U613 (.ZN( u1_K11_35 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1695 ) , .A2( u1_uk_n1703 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U614 (.ZN( u1_K8_35 ) , .B2( u1_uk_n1541 ) , .A2( u1_uk_n1547 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U615 (.ZN( u1_K7_35 ) , .A( u1_uk_n1120 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1482 ) );
  NAND2_X1 u1_uk_U616 (.A1( u1_uk_K_r5_37 ) , .ZN( u1_uk_n1120 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U617 (.ZN( u1_K15_35 ) , .B2( u1_uk_n1860 ) , .A2( u1_uk_n1875 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U618 (.ZN( u1_K13_35 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1764 ) , .A2( u1_uk_n1793 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U619 (.ZN( u1_K12_35 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1728 ) , .A2( u1_uk_n1737 ) , .B1( u1_uk_n213 ) );
  BUF_X1 u1_uk_U62 (.Z( u1_uk_n292 ) , .A( u1_uk_n294 ) );
  INV_X1 u1_uk_U620 (.ZN( u1_K14_35 ) , .A( u1_uk_n956 ) );
  AOI22_X1 u1_uk_U621 (.B2( u1_uk_K_r12_1 ) , .A2( u1_uk_K_r12_7 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n242 ) , .ZN( u1_uk_n956 ) );
  AOI22_X1 u1_uk_U623 (.B2( u1_uk_K_r8_2 ) , .A2( u1_uk_K_r8_37 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n252 ) , .ZN( u1_uk_n353 ) );
  INV_X1 u1_uk_U624 (.ZN( u1_K9_35 ) , .A( u1_uk_n1163 ) );
  AOI22_X1 u1_uk_U625 (.B2( u1_uk_K_r7_16 ) , .A2( u1_uk_K_r7_23 ) , .ZN( u1_uk_n1163 ) , .B1( u1_uk_n129 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U626 (.ZN( u1_K6_35 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1469 ) , .A2( u1_uk_n1476 ) , .A1( u1_uk_n203 ) );
  INV_X1 u1_uk_U627 (.ZN( u1_K5_35 ) , .A( u1_uk_n1079 ) );
  AOI22_X1 u1_uk_U628 (.B2( u1_uk_K_r3_29 ) , .A2( u1_uk_K_r3_38 ) , .ZN( u1_uk_n1079 ) , .B1( u1_uk_n251 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U629 (.ZN( u1_K4_35 ) , .B2( u1_uk_n1361 ) , .A2( u1_uk_n1390 ) , .B1( u1_uk_n142 ) , .A1( u1_uk_n271 ) );
  BUF_X1 u1_uk_U63 (.Z( u1_uk_n257 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U630 (.ZN( u1_K2_35 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1275 ) , .A2( u1_uk_n1293 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U631 (.ZN( u1_K1_35 ) , .A( u1_uk_n1012 ) );
  AOI22_X1 u1_uk_U632 (.B2( u1_key_r_28 ) , .A2( u1_key_r_35 ) , .ZN( u1_uk_n1012 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U633 (.ZN( u1_K16_11 ) , .B2( u1_uk_n1242 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n978 ) );
  NAND2_X1 u1_uk_U634 (.A1( u1_uk_K_r14_39 ) , .A2( u1_uk_n94 ) , .ZN( u1_uk_n978 ) );
  OAI21_X1 u1_uk_U635 (.ZN( u1_K15_11 ) , .B2( u1_uk_n1880 ) , .B1( u1_uk_n250 ) , .A( u1_uk_n965 ) );
  NAND2_X1 u1_uk_U636 (.A1( u1_uk_K_r13_25 ) , .A2( u1_uk_n230 ) , .ZN( u1_uk_n965 ) );
  OAI22_X1 u1_uk_U637 (.ZN( u1_K14_11 ) , .A2( u1_uk_n1801 ) , .B2( u1_uk_n1808 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U638 (.ZN( u1_K11_11 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1676 ) , .A2( u1_uk_n1682 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U639 (.ZN( u1_K3_11 ) , .A2( u1_uk_n1310 ) , .B2( u1_uk_n1315 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n191 ) );
  BUF_X1 u1_uk_U64 (.Z( u1_uk_n294 ) , .A( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U640 (.ZN( u1_K2_11 ) , .A( u1_uk_n1022 ) , .B2( u1_uk_n1297 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U641 (.A1( u1_uk_K_r0_25 ) , .ZN( u1_uk_n1022 ) , .A2( u1_uk_n141 ) );
  AOI22_X1 u1_uk_U643 (.B2( u1_uk_K_r11_17 ) , .A2( u1_uk_K_r11_54 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n191 ) , .ZN( u1_uk_n672 ) );
  OAI22_X1 u1_uk_U644 (.ZN( u1_K10_11 ) , .B2( u1_uk_n1626 ) , .A2( u1_uk_n1643 ) , .A1( u1_uk_n214 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U645 (.ZN( u1_K8_11 ) , .A( u1_uk_n1127 ) , .B2( u1_uk_n1565 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U646 (.A1( u1_uk_K_r6_55 ) , .ZN( u1_uk_n1127 ) , .A2( u1_uk_n147 ) );
  OAI22_X1 u1_uk_U647 (.ZN( u1_K7_11 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1488 ) , .A2( u1_uk_n1505 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U648 (.ZN( u1_K6_11 ) , .B2( u1_uk_n1453 ) , .A2( u1_uk_n1457 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U649 (.ZN( u1_K5_11 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1399 ) , .B2( u1_uk_n1423 ) , .B1( u1_uk_n220 ) );
  BUF_X1 u1_uk_U65 (.Z( u1_uk_n297 ) , .A( u1_uk_n298 ) );
  INV_X1 u1_uk_U650 (.ZN( u1_K4_23 ) , .A( u1_uk_n1056 ) );
  AOI22_X1 u1_uk_U651 (.B2( u1_uk_K_r2_18 ) , .A2( u1_uk_K_r2_55 ) , .ZN( u1_uk_n1056 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U652 (.ZN( u1_K16_45 ) , .B2( u1_uk_n1247 ) , .A2( u1_uk_n1250 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U653 (.ZN( u1_K1_45 ) , .B2( u1_uk_n1201 ) , .A2( u1_uk_n1208 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n242 ) );
  INV_X1 u1_uk_U654 (.A( u1_key_r_44 ) , .ZN( u1_uk_n1208 ) );
  OAI22_X1 u1_uk_U655 (.ZN( u1_K14_43 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1829 ) , .A2( u1_uk_n1832 ) , .B1( u1_uk_n231 ) );
  OAI21_X1 u1_uk_U656 (.ZN( u1_K4_43 ) , .A( u1_uk_n1066 ) , .B2( u1_uk_n1389 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U657 (.A1( u1_uk_K_r2_29 ) , .ZN( u1_uk_n1066 ) , .A2( u1_uk_n128 ) );
  OAI22_X1 u1_uk_U658 (.ZN( u1_K3_43 ) , .B2( u1_uk_n1334 ) , .A2( u1_uk_n1338 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U659 (.ZN( u1_K2_43 ) , .A( u1_uk_n1032 ) , .B2( u1_uk_n1276 ) , .B1( u1_uk_n162 ) );
  INV_X1 u1_uk_U66 (.A( n116 ) , .ZN( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U660 (.A1( u1_uk_K_r0_2 ) , .ZN( u1_uk_n1032 ) , .A2( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U661 (.ZN( u1_K11_3 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1669 ) , .A2( u1_uk_n1687 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U662 (.ZN( u1_K1_7 ) , .B2( u1_uk_n1185 ) , .A2( u1_uk_n1192 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U663 (.ZN( u1_K4_7 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1353 ) , .B2( u1_uk_n1357 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U664 (.ZN( u1_K9_25 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1608 ) , .A2( u1_uk_n1615 ) , .B1( u1_uk_n292 ) );
  INV_X1 u1_uk_U665 (.ZN( u1_K16_43 ) , .A( u1_uk_n993 ) );
  AOI22_X1 u1_uk_U666 (.B2( u1_uk_K_r14_16 ) , .A2( u1_uk_K_r14_9 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) , .ZN( u1_uk_n993 ) );
  INV_X1 u1_uk_U667 (.ZN( u1_K5_43 ) , .A( u1_uk_n1083 ) );
  AOI22_X1 u1_uk_U668 (.B2( u1_uk_K_r3_15 ) , .A2( u1_uk_K_r3_38 ) , .ZN( u1_uk_n1083 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U669 (.ZN( u1_K14_45 ) , .B2( u1_uk_n1830 ) , .B1( u1_uk_n251 ) , .A( u1_uk_n960 ) );
  NAND2_X1 u1_uk_U670 (.A1( u1_uk_K_r12_16 ) , .A2( u1_uk_n292 ) , .ZN( u1_uk_n960 ) );
  OAI21_X1 u1_uk_U671 (.ZN( u1_K13_43 ) , .B2( u1_uk_n1792 ) , .B1( u1_uk_n191 ) , .A( u1_uk_n946 ) );
  NAND2_X1 u1_uk_U672 (.A1( u1_uk_K_r11_29 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n946 ) );
  OAI21_X1 u1_uk_U673 (.ZN( u1_K12_45 ) , .B2( u1_uk_n1714 ) , .B1( u1_uk_n191 ) , .A( u1_uk_n634 ) );
  NAND2_X1 u1_uk_U674 (.A1( u1_uk_K_r10_43 ) , .A2( u1_uk_n214 ) , .ZN( u1_uk_n634 ) );
  OAI22_X1 u1_uk_U675 (.ZN( u1_K11_43 ) , .B1( u1_uk_n146 ) , .B2( u1_uk_n1662 ) , .A2( u1_uk_n1704 ) , .A1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U676 (.ZN( u1_K10_43 ) , .A2( u1_uk_n1623 ) , .B2( u1_uk_n1651 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U677 (.ZN( u1_K10_45 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1628 ) , .A2( u1_uk_n1644 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U678 (.ZN( u1_K9_43 ) , .A1( u1_uk_n11 ) , .B2( u1_uk_n1588 ) , .A2( u1_uk_n1595 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U679 (.ZN( u1_K9_45 ) , .B2( u1_uk_n1571 ) , .A2( u1_uk_n1612 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U68 (.A1( n116 ) , .B2( u1_uk_K_r14_2 ) , .A2( u1_uk_K_r14_9 ) , .B1( u1_uk_n213 ) , .ZN( u1_uk_n988 ) );
  OAI22_X1 u1_uk_U680 (.ZN( u1_K7_43 ) , .A1( u1_uk_n141 ) , .A2( u1_uk_n1485 ) , .B2( u1_uk_n1514 ) , .B1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U681 (.ZN( u1_K10_7 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1634 ) , .A2( u1_uk_n1654 ) , .A1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U682 (.ZN( u1_K6_7 ) , .A( u1_uk_n1102 ) , .B2( u1_uk_n1465 ) , .B1( u1_uk_n222 ) );
  NAND2_X1 u1_uk_U683 (.A1( u1_uk_K_r4_33 ) , .ZN( u1_uk_n1102 ) , .A2( u1_uk_n208 ) );
  OAI21_X1 u1_uk_U684 (.ZN( u1_K12_7 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1750 ) , .A( u1_uk_n665 ) );
  NAND2_X1 u1_uk_U685 (.A1( u1_uk_K_r10_19 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n665 ) );
  OAI21_X1 u1_uk_U686 (.ZN( u1_K11_7 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1691 ) , .A( u1_uk_n500 ) );
  NAND2_X1 u1_uk_U687 (.A1( u1_uk_K_r9_33 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n500 ) );
  OAI21_X1 u1_uk_U688 (.ZN( u1_K15_25 ) , .B2( u1_uk_n1876 ) , .B1( u1_uk_n223 ) , .A( u1_uk_n968 ) );
  NAND2_X1 u1_uk_U689 (.A1( u1_uk_K_r13_22 ) , .A2( u1_uk_n213 ) , .ZN( u1_uk_n968 ) );
  OAI22_X1 u1_uk_U690 (.ZN( u1_K11_25 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1677 ) , .A2( u1_uk_n1696 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U691 (.ZN( u1_K13_25 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1765 ) , .A2( u1_uk_n1790 ) , .B1( u1_uk_n191 ) );
  OAI21_X1 u1_uk_U692 (.ZN( u1_K2_25 ) , .A( u1_uk_n1026 ) , .B2( u1_uk_n1294 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U693 (.A1( u1_uk_K_r0_22 ) , .ZN( u1_uk_n1026 ) , .A2( u1_uk_n109 ) );
  OAI22_X1 u1_uk_U694 (.ZN( u1_K16_25 ) , .B2( u1_uk_n1239 ) , .A2( u1_uk_n1246 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U695 (.ZN( u1_K12_25 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1729 ) , .A2( u1_uk_n1734 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U696 (.ZN( u1_K10_25 ) , .A1( u1_uk_n109 ) , .A2( u1_uk_n1623 ) , .B2( u1_uk_n1641 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U697 (.ZN( u1_K8_25 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1563 ) , .A2( u1_uk_n1568 ) , .A1( u1_uk_n214 ) );
  INV_X1 u1_uk_U698 (.ZN( u1_K8_43 ) , .A( u1_uk_n1143 ) );
  AOI22_X1 u1_uk_U699 (.B2( u1_uk_K_r6_21 ) , .A2( u1_uk_K_r6_28 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1143 ) , .B1( u1_uk_n277 ) );
  INV_X1 u1_uk_U7 (.ZN( u1_uk_n102 ) , .A( u1_uk_n230 ) );
  AOI22_X1 u1_uk_U70 (.B2( u1_uk_K_r9_45 ) , .A2( u1_uk_K_r9_49 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n443 ) );
  OAI22_X1 u1_uk_U700 (.ZN( u1_K16_3 ) , .B2( u1_uk_n1228 ) , .A2( u1_uk_n1236 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U701 (.ZN( u1_K15_7 ) , .B2( u1_uk_n1853 ) , .A2( u1_uk_n1869 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U702 (.ZN( u1_K16_7 ) , .B2( u1_uk_n1229 ) , .A2( u1_uk_n1237 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n60 ) );
  AOI22_X1 u1_uk_U704 (.B2( u1_uk_K_r10_18 ) , .A2( u1_uk_K_r10_27 ) , .B1( u1_uk_n129 ) , .A1( u1_uk_n231 ) , .ZN( u1_uk_n601 ) );
  INV_X1 u1_uk_U705 (.ZN( u1_K8_3 ) , .A( u1_uk_n1140 ) );
  AOI22_X1 u1_uk_U706 (.B2( u1_uk_K_r6_10 ) , .A2( u1_uk_K_r6_3 ) , .ZN( u1_uk_n1140 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n294 ) );
  AOI22_X1 u1_uk_U708 (.A2( u1_uk_K_r2_4 ) , .B2( u1_uk_K_r2_41 ) , .ZN( u1_uk_n1065 ) , .B1( u1_uk_n161 ) , .A1( u1_uk_n188 ) );
  INV_X1 u1_uk_U709 (.ZN( u1_K13_7 ) , .A( u1_uk_n950 ) );
  AOI22_X1 u1_uk_U710 (.B2( u1_uk_K_r11_10 ) , .A2( u1_uk_K_r11_5 ) , .B1( u1_uk_n207 ) , .A1( u1_uk_n93 ) , .ZN( u1_uk_n950 ) );
  OAI21_X1 u1_uk_U711 (.ZN( u1_K5_7 ) , .A( u1_uk_n1087 ) , .B2( u1_uk_n1435 ) , .B1( u1_uk_n250 ) );
  NAND2_X1 u1_uk_U712 (.A1( u1_uk_K_r3_19 ) , .ZN( u1_uk_n1087 ) , .A2( u1_uk_n188 ) );
  INV_X1 u1_uk_U713 (.ZN( u1_K1_25 ) , .A( u1_uk_n1005 ) );
  AOI22_X1 u1_uk_U714 (.B2( u1_key_r_29 ) , .A2( u1_key_r_36 ) , .ZN( u1_uk_n1005 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n250 ) );
  INV_X1 u1_uk_U715 (.ZN( u1_K4_25 ) , .A( u1_uk_n1057 ) );
  AOI22_X1 u1_uk_U716 (.B2( u1_uk_K_r2_16 ) , .A2( u1_uk_K_r2_49 ) , .ZN( u1_uk_n1057 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U717 (.ZN( u1_K12_2 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1711 ) , .B2( u1_uk_n1716 ) , .A1( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U718 (.ZN( u1_K10_2 ) , .B2( u1_uk_n1622 ) , .B1( u1_uk_n257 ) , .A( u1_uk_n338 ) );
  NAND2_X1 u1_uk_U719 (.A1( u1_uk_K_r8_41 ) , .A2( u1_uk_n188 ) , .ZN( u1_uk_n338 ) );
  AOI22_X1 u1_uk_U72 (.B2( u1_uk_K_r6_14 ) , .A2( u1_uk_K_r6_21 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1137 ) , .B1( u1_uk_n214 ) );
  OAI21_X1 u1_uk_U720 (.ZN( u1_K1_2 ) , .A( u1_uk_n1008 ) , .B2( u1_uk_n1175 ) , .B1( u1_uk_n242 ) );
  NAND2_X1 u1_uk_U721 (.A1( u1_key_r_11 ) , .ZN( u1_uk_n1008 ) , .A2( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U722 (.ZN( u1_K4_32 ) , .A1( u1_uk_n110 ) , .A2( u1_uk_n1356 ) , .B2( u1_uk_n1380 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U723 (.ZN( u1_K16_32 ) , .B2( u1_uk_n1231 ) , .A2( u1_uk_n1239 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U724 (.ZN( u1_K8_32 ) , .B2( u1_uk_n1556 ) , .A2( u1_uk_n1563 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U725 (.ZN( u1_K11_32 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1670 ) , .A2( u1_uk_n1690 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U726 (.ZN( u1_K13_32 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1758 ) , .B2( u1_uk_n1782 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U727 (.ZN( u1_K6_32 ) , .B2( u1_uk_n1448 ) , .A2( u1_uk_n1464 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U728 (.ZN( u1_K3_32 ) , .B2( u1_uk_n1308 ) , .A2( u1_uk_n1343 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U729 (.ZN( u1_K5_32 ) , .B2( u1_uk_n1408 ) , .A2( u1_uk_n1412 ) , .B1( u1_uk_n147 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U730 (.ZN( u1_K14_32 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1799 ) , .A2( u1_uk_n1837 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U731 (.ZN( u1_K9_32 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1601 ) , .A2( u1_uk_n1608 ) , .B1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U732 (.ZN( u1_K15_42 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1879 ) , .A2( u1_uk_n1885 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U733 (.ZN( u1_K14_42 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1798 ) , .A2( u1_uk_n1829 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U734 (.ZN( u1_K13_42 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1763 ) , .A2( u1_uk_n1769 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U735 (.ZN( u1_K11_42 ) , .A1( u1_uk_n164 ) , .B2( u1_uk_n1694 ) , .A2( u1_uk_n1702 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U736 (.ZN( u1_K10_42 ) , .B2( u1_uk_n1619 ) , .A1( u1_uk_n162 ) , .A2( u1_uk_n1645 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U737 (.ZN( u1_K4_42 ) , .B2( u1_uk_n1360 ) , .A2( u1_uk_n1367 ) , .B1( u1_uk_n141 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U738 (.ZN( u1_K3_42 ) , .B2( u1_uk_n1307 ) , .A2( u1_uk_n1334 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U739 (.ZN( u1_K2_42 ) , .B2( u1_uk_n1296 ) , .A2( u1_uk_n1304 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U74 (.B2( u1_uk_K_r5_0 ) , .A2( u1_uk_K_r5_35 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1119 ) , .B1( u1_uk_n209 ) );
  INV_X1 u1_uk_U740 (.ZN( u1_K12_42 ) , .A( u1_uk_n605 ) );
  AOI22_X1 u1_uk_U741 (.B2( u1_uk_K_r10_28 ) , .A2( u1_uk_K_r10_9 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n294 ) , .ZN( u1_uk_n605 ) );
  INV_X1 u1_uk_U742 (.ZN( u1_K9_42 ) , .A( u1_uk_n1167 ) );
  AOI22_X1 u1_uk_U743 (.B2( u1_uk_K_r7_15 ) , .A2( u1_uk_K_r7_22 ) , .ZN( u1_uk_n1167 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n291 ) );
  INV_X1 u1_uk_U744 (.ZN( u1_K7_42 ) , .A( u1_uk_n1123 ) );
  AOI22_X1 u1_uk_U745 (.B2( u1_uk_K_r5_1 ) , .A2( u1_uk_K_r5_36 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1123 ) , .B1( u1_uk_n297 ) );
  INV_X1 u1_uk_U746 (.ZN( u1_K1_42 ) , .A( u1_uk_n1016 ) );
  AOI22_X1 u1_uk_U747 (.B2( u1_key_r_31 ) , .A2( u1_key_r_38 ) , .ZN( u1_uk_n1016 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U748 (.ZN( u1_K14_27 ) , .B2( u1_uk_n1839 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n953 ) );
  NAND2_X1 u1_uk_U749 (.A1( u1_uk_K_r12_42 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n953 ) );
  OAI22_X1 u1_uk_U75 (.ZN( u1_K15_34 ) , .A1( u1_uk_n148 ) , .B2( u1_uk_n1856 ) , .A2( u1_uk_n1884 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U750 (.ZN( u1_K12_27 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1717 ) , .A2( u1_uk_n1749 ) , .B1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U751 (.ZN( u1_K10_27 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1632 ) , .A( u1_uk_n335 ) );
  NAND2_X1 u1_uk_U752 (.A1( u1_uk_K_r8_43 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n335 ) );
  OAI22_X1 u1_uk_U753 (.ZN( u1_K8_27 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1529 ) , .A2( u1_uk_n1534 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U754 (.ZN( u1_K16_27 ) , .B2( u1_uk_n1225 ) , .A2( u1_uk_n1230 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U755 (.ZN( u1_K12_13 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1719 ) , .A2( u1_uk_n1751 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U756 (.ZN( u1_K11_13 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1688 ) , .A2( u1_uk_n1692 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U757 (.ZN( u1_K8_13 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1531 ) , .B2( u1_uk_n1537 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U758 (.ZN( u1_K6_13 ) , .B2( u1_uk_n1462 ) , .A2( u1_uk_n1466 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U759 (.ZN( u1_K2_13 ) , .A2( u1_uk_n1261 ) , .B2( u1_uk_n1290 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U760 (.ZN( u1_K1_21 ) , .B2( u1_uk_n1183 ) , .A2( u1_uk_n1189 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n222 ) );
  OAI21_X1 u1_uk_U761 (.ZN( u1_K9_13 ) , .A( u1_uk_n1150 ) , .B2( u1_uk_n1579 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U762 (.A1( u1_uk_K_r7_5 ) , .ZN( u1_uk_n1150 ) , .A2( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U763 (.ZN( u1_K11_27 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1684 ) , .A2( u1_uk_n1690 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U764 (.ZN( u1_K13_27 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1754 ) , .A2( u1_uk_n1777 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U765 (.ZN( u1_K14_21 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1814 ) , .A2( u1_uk_n1840 ) , .B1( u1_uk_n220 ) );
  OAI21_X1 u1_uk_U766 (.ZN( u1_K11_21 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1667 ) , .A( u1_uk_n395 ) );
  NAND2_X1 u1_uk_U767 (.A1( u1_uk_K_r9_5 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n395 ) );
  OAI22_X1 u1_uk_U768 (.ZN( u1_K9_21 ) , .B2( u1_uk_n1598 ) , .A2( u1_uk_n1603 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U769 (.ZN( u1_K5_21 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1409 ) , .A2( u1_uk_n1429 ) , .B1( u1_uk_n202 ) );
  AOI22_X1 u1_uk_U77 (.B2( u1_uk_K_r12_30 ) , .A2( u1_uk_K_r12_36 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n279 ) , .ZN( u1_uk_n955 ) );
  OAI22_X1 u1_uk_U770 (.ZN( u1_K2_21 ) , .A2( u1_uk_n1264 ) , .B2( u1_uk_n1268 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n223 ) );
  OAI21_X1 u1_uk_U771 (.ZN( u1_K7_21 ) , .A( u1_uk_n1110 ) , .B2( u1_uk_n1526 ) , .B1( u1_uk_n271 ) );
  NAND2_X1 u1_uk_U772 (.A1( u1_uk_K_r5_19 ) , .ZN( u1_uk_n1110 ) , .A2( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U773 (.ZN( u1_K4_21 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1371 ) , .A2( u1_uk_n1377 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U774 (.ZN( u1_K15_21 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1846 ) , .B2( u1_uk_n1850 ) , .A1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U775 (.ZN( u1_K14_13 ) , .B2( u1_uk_n1812 ) , .A2( u1_uk_n1817 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U776 (.ZN( u1_K4_27 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1350 ) , .A2( u1_uk_n1376 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U777 (.ZN( u1_K15_27 ) , .A1( u1_uk_n148 ) , .A2( u1_uk_n1847 ) , .B2( u1_uk_n1865 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U778 (.ZN( u1_K4_13 ) , .A2( u1_uk_n1354 ) , .B2( u1_uk_n1358 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n209 ) );
  INV_X1 u1_uk_U779 (.ZN( u1_K12_21 ) , .A( u1_uk_n520 ) );
  OAI22_X1 u1_uk_U78 (.ZN( u1_K12_34 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1715 ) , .B2( u1_uk_n1730 ) , .B1( u1_uk_n213 ) );
  AOI22_X1 u1_uk_U780 (.B2( u1_uk_K_r10_25 ) , .A2( u1_uk_K_r10_48 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n250 ) , .ZN( u1_uk_n520 ) );
  AOI22_X1 u1_uk_U782 (.B2( u1_uk_K_r11_11 ) , .A2( u1_uk_K_r11_6 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n240 ) , .ZN( u1_uk_n677 ) );
  INV_X1 u1_uk_U783 (.ZN( u1_K13_21 ) , .A( u1_uk_n689 ) );
  AOI22_X1 u1_uk_U784 (.B2( u1_uk_K_r11_34 ) , .A2( u1_uk_K_r11_39 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n230 ) , .ZN( u1_uk_n689 ) );
  INV_X1 u1_uk_U785 (.ZN( u1_K6_21 ) , .A( u1_uk_n1092 ) );
  AOI22_X1 u1_uk_U786 (.B2( u1_uk_K_r4_11 ) , .A2( u1_uk_K_r4_5 ) , .ZN( u1_uk_n1092 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n298 ) );
  OAI21_X1 u1_uk_U787 (.ZN( u1_K16_13 ) , .B2( u1_uk_n1257 ) , .B1( u1_uk_n297 ) , .A( u1_uk_n980 ) );
  NAND2_X1 u1_uk_U788 (.A1( u1_uk_K_r14_46 ) , .A2( u1_uk_n242 ) , .ZN( u1_uk_n980 ) );
  OAI22_X1 u1_uk_U789 (.ZN( u1_K6_27 ) , .B2( u1_uk_n1459 ) , .A2( u1_uk_n1464 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n93 ) );
  OAI21_X1 u1_uk_U79 (.ZN( u1_K6_34 ) , .A( u1_uk_n1097 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1471 ) );
  AOI22_X1 u1_uk_U791 (.B2( u1_uk_K_r3_15 ) , .A2( u1_uk_K_r3_51 ) , .ZN( u1_uk_n1076 ) , .B1( u1_uk_n240 ) , .A1( u1_uk_n83 ) );
  INV_X1 u1_uk_U792 (.ZN( u1_K2_27 ) , .A( u1_uk_n1027 ) );
  AOI22_X1 u1_uk_U793 (.B2( u1_uk_K_r0_28 ) , .A2( u1_uk_K_r0_7 ) , .ZN( u1_uk_n1027 ) , .A1( u1_uk_n129 ) , .B1( u1_uk_n252 ) );
  OAI21_X1 u1_uk_U794 (.ZN( u1_K3_27 ) , .A( u1_uk_n1039 ) , .B2( u1_uk_n1345 ) , .B1( u1_uk_n231 ) );
  NAND2_X1 u1_uk_U795 (.A1( u1_uk_K_r1_42 ) , .ZN( u1_uk_n1039 ) , .A2( u1_uk_n298 ) );
  AOI22_X1 u1_uk_U797 (.B2( u1_uk_K_r5_23 ) , .A2( u1_uk_K_r5_43 ) , .ZN( u1_uk_n1115 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n203 ) );
  AOI22_X1 u1_uk_U799 (.B2( u1_key_r_14 ) , .A2( u1_key_r_21 ) , .ZN( u1_uk_n1007 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n257 ) );
  INV_X1 u1_uk_U8 (.A( u1_uk_n203 ) , .ZN( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U80 (.A1( u1_uk_K_r4_49 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1097 ) );
  AOI22_X1 u1_uk_U801 (.B2( u1_uk_K_r7_2 ) , .A2( u1_uk_K_r7_9 ) , .B1( u1_uk_n100 ) , .ZN( u1_uk_n1159 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U802 (.ZN( u1_K16_1 ) , .B2( u1_uk_n1248 ) , .A2( u1_uk_n1251 ) , .A1( u1_uk_n220 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U803 (.ZN( u1_K13_1 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1757 ) , .A( u1_uk_n686 ) );
  NAND2_X1 u1_uk_U804 (.A1( u1_uk_K_r11_25 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n686 ) );
  OAI22_X1 u1_uk_U805 (.ZN( u1_K6_1 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1462 ) , .A2( u1_uk_n1478 ) , .B1( u1_uk_n188 ) );
  INV_X1 u1_uk_U806 (.ZN( u1_K9_1 ) , .A( u1_uk_n1155 ) );
  AOI22_X1 u1_uk_U807 (.B2( u1_uk_K_r7_24 ) , .A2( u1_uk_K_r7_6 ) , .ZN( u1_uk_n1155 ) , .B1( u1_uk_n155 ) , .A1( u1_uk_n250 ) );
  OAI21_X1 u1_uk_U808 (.ZN( u1_K4_1 ) , .A( u1_uk_n1053 ) , .B2( u1_uk_n1353 ) , .B1( u1_uk_n252 ) );
  NAND2_X1 u1_uk_U809 (.A1( u1_uk_K_r2_25 ) , .ZN( u1_uk_n1053 ) , .A2( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U81 (.ZN( u1_K4_34 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1366 ) , .A2( u1_uk_n1382 ) , .B1( u1_uk_n202 ) );
  OAI21_X1 u1_uk_U810 (.ZN( u1_K4_18 ) , .A( u1_uk_n1052 ) , .B2( u1_uk_n1378 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U811 (.A1( u1_uk_K_r2_20 ) , .ZN( u1_uk_n1052 ) , .A2( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U812 (.ZN( u1_K5_18 ) , .A2( u1_uk_n1399 ) , .B2( u1_uk_n1436 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U813 (.ZN( u1_K13_20 ) , .B1( u1_uk_n128 ) , .B2( u1_uk_n1762 ) , .A( u1_uk_n688 ) );
  NAND2_X1 u1_uk_U814 (.A1( u1_uk_K_r11_33 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n688 ) );
  OAI21_X1 u1_uk_U815 (.ZN( u1_K13_18 ) , .B2( u1_uk_n1780 ) , .B1( u1_uk_n231 ) , .A( u1_uk_n682 ) );
  NAND2_X1 u1_uk_U816 (.A1( u1_uk_K_r11_20 ) , .A2( u1_uk_n291 ) , .ZN( u1_uk_n682 ) );
  OAI22_X1 u1_uk_U817 (.ZN( u1_K7_18 ) , .A2( u1_uk_n1483 ) , .B2( u1_uk_n1496 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n92 ) );
  OAI21_X1 u1_uk_U818 (.ZN( u1_K8_18 ) , .A( u1_uk_n1132 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1557 ) );
  NAND2_X1 u1_uk_U819 (.A1( u1_uk_K_r6_46 ) , .ZN( u1_uk_n1132 ) , .A2( u1_uk_n146 ) );
  OAI21_X1 u1_uk_U82 (.ZN( u1_K3_34 ) , .B1( u1_uk_n100 ) , .A( u1_uk_n1041 ) , .B2( u1_uk_n1329 ) );
  OAI22_X1 u1_uk_U820 (.ZN( u1_K2_18 ) , .B2( u1_uk_n1269 ) , .A2( u1_uk_n1300 ) , .A1( u1_uk_n252 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U821 (.ZN( u1_K16_18 ) , .B2( u1_uk_n1259 ) , .B1( u1_uk_n94 ) , .A( u1_uk_n983 ) );
  NAND2_X1 u1_uk_U822 (.A1( u1_uk_K_r14_5 ) , .A2( u1_uk_n118 ) , .ZN( u1_uk_n983 ) );
  OAI22_X1 u1_uk_U823 (.ZN( u1_K10_18 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1620 ) , .B2( u1_uk_n1634 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U824 (.ZN( u1_K15_18 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1852 ) , .A2( u1_uk_n1882 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U825 (.ZN( u1_K3_20 ) , .B2( u1_uk_n1320 ) , .A2( u1_uk_n1326 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U826 (.ZN( u1_K12_20 ) , .B1( u1_uk_n162 ) , .B2( u1_uk_n1722 ) , .A( u1_uk_n518 ) );
  NAND2_X1 u1_uk_U827 (.A1( u1_uk_K_r10_47 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n518 ) );
  OAI22_X1 u1_uk_U828 (.ZN( u1_K16_20 ) , .B2( u1_uk_n1252 ) , .A2( u1_uk_n1259 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U829 (.ZN( u1_K15_20 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1845 ) , .B2( u1_uk_n1874 ) , .A1( u1_uk_n298 ) );
  NAND2_X1 u1_uk_U83 (.A1( u1_uk_K_r1_36 ) , .ZN( u1_uk_n1041 ) , .A2( u1_uk_n27 ) );
  OAI22_X1 u1_uk_U830 (.ZN( u1_K8_20 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1551 ) , .A2( u1_uk_n1557 ) , .A1( u1_uk_n222 ) );
  INV_X1 u1_uk_U831 (.ZN( u1_K9_18 ) , .A( u1_uk_n1153 ) );
  AOI22_X1 u1_uk_U832 (.B2( u1_uk_K_r7_39 ) , .A2( u1_uk_K_r7_46 ) , .ZN( u1_uk_n1153 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n230 ) );
  INV_X1 u1_uk_U833 (.ZN( u1_K6_18 ) , .A( u1_uk_n1090 ) );
  AOI22_X1 u1_uk_U834 (.B2( u1_uk_K_r4_11 ) , .A2( u1_uk_K_r4_17 ) , .ZN( u1_uk_n1090 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n252 ) );
  AOI22_X1 u1_uk_U836 (.B2( u1_uk_K_r9_10 ) , .A2( u1_uk_K_r9_4 ) , .A1( u1_uk_n100 ) , .B1( u1_uk_n292 ) , .ZN( u1_uk_n391 ) );
  INV_X1 u1_uk_U837 (.ZN( u1_K7_20 ) , .A( u1_uk_n1109 ) );
  AOI22_X1 u1_uk_U838 (.B2( u1_uk_K_r5_18 ) , .A2( u1_uk_K_r5_53 ) , .A1( u1_uk_n11 ) , .ZN( u1_uk_n1109 ) , .B1( u1_uk_n207 ) );
  INV_X1 u1_uk_U839 (.ZN( u1_K5_20 ) , .A( u1_uk_n1073 ) );
  OAI22_X1 u1_uk_U84 (.ZN( u1_K2_34 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1272 ) , .A2( u1_uk_n1303 ) , .A1( u1_uk_n217 ) );
  AOI22_X1 u1_uk_U840 (.B2( u1_uk_K_r3_24 ) , .A2( u1_uk_K_r3_47 ) , .ZN( u1_uk_n1073 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n83 ) );
  OAI21_X1 u1_uk_U841 (.ZN( u1_K4_22 ) , .A( u1_uk_n1055 ) , .B2( u1_uk_n1357 ) , .B1( u1_uk_n161 ) );
  NAND2_X1 u1_uk_U842 (.A1( u1_uk_K_r2_47 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n1055 ) );
  OAI22_X1 u1_uk_U843 (.ZN( u1_K1_6 ) , .B2( u1_uk_n1198 ) , .A2( u1_uk_n1205 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n240 ) );
  INV_X1 u1_uk_U844 (.A( u1_key_r_41 ) , .ZN( u1_uk_n1205 ) );
  OAI22_X1 u1_uk_U845 (.ZN( u1_K15_6 ) , .B2( u1_uk_n1864 ) , .A2( u1_uk_n1882 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U846 (.ZN( u1_K1_43 ) , .A2( u1_uk_n1179 ) , .B2( u1_uk_n1182 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n60 ) );
  OAI21_X1 u1_uk_U847 (.ZN( u1_K13_3 ) , .B2( u1_uk_n1781 ) , .B1( u1_uk_n27 ) , .A( u1_uk_n945 ) );
  NAND2_X1 u1_uk_U848 (.A1( u1_uk_K_r11_4 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n945 ) );
  OAI22_X1 u1_uk_U849 (.ZN( u1_K7_3 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1495 ) , .A2( u1_uk_n1517 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U85 (.ZN( u1_K16_23 ) , .B2( u1_uk_n1243 ) , .A2( u1_uk_n1248 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U850 (.ZN( u1_K15_3 ) , .B2( u1_uk_n1852 ) , .A2( u1_uk_n1868 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n83 ) );
  INV_X1 u1_uk_U851 (.ZN( u1_K7_6 ) , .A( u1_uk_n1125 ) );
  AOI22_X1 u1_uk_U852 (.B2( u1_uk_K_r5_39 ) , .A2( u1_uk_K_r5_4 ) , .ZN( u1_uk_n1125 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U853 (.ZN( u1_K14_3 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1842 ) , .A( u1_uk_n957 ) );
  NAND2_X1 u1_uk_U854 (.A1( u1_uk_K_r12_47 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n957 ) );
  OAI21_X1 u1_uk_U855 (.ZN( u1_K3_3 ) , .A( u1_uk_n1043 ) , .B2( u1_uk_n1348 ) , .B1( u1_uk_n242 ) );
  NAND2_X1 u1_uk_U856 (.A1( u1_uk_K_r1_47 ) , .ZN( u1_uk_n1043 ) , .A2( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U857 (.ZN( u1_K16_2 ) , .B2( u1_uk_n1220 ) , .B1( u1_uk_n155 ) , .A( u1_uk_n986 ) );
  NAND2_X1 u1_uk_U858 (.A1( u1_uk_K_r14_11 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n986 ) );
  AOI22_X1 u1_uk_U859 (.B2( u1_uk_K_r7_20 ) , .A2( u1_uk_K_r7_27 ) , .ZN( u1_uk_n1160 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n286 ) );
  INV_X1 u1_uk_U86 (.ZN( u1_K12_23 ) , .A( u1_uk_n524 ) );
  AOI22_X1 u1_uk_U860 (.B2( u1_uk_K_r2_26 ) , .A2( u1_uk_K_r2_46 ) , .ZN( u1_uk_n1061 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n279 ) );
  OAI21_X1 u1_uk_U861 (.ZN( u1_K10_1 ) , .B2( u1_uk_n1630 ) , .A( u1_uk_n306 ) , .B1( u1_uk_n31 ) );
  NAND2_X1 u1_uk_U862 (.A1( u1_uk_K_r8_10 ) , .A2( u1_uk_n118 ) , .ZN( u1_uk_n306 ) );
  OAI22_X1 u1_uk_U863 (.ZN( u1_K1_1 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1204 ) , .A2( u1_uk_n1209 ) , .B1( u1_uk_n240 ) );
  AOI22_X1 u1_uk_U864 (.B2( u1_uk_K_r10_39 ) , .A2( u1_uk_K_r10_48 ) , .B1( u1_uk_n155 ) , .A1( u1_uk_n213 ) , .ZN( u1_uk_n515 ) );
  AOI22_X1 u1_uk_U865 (.B2( u1_uk_K_r11_19 ) , .A2( u1_uk_K_r11_24 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n220 ) , .ZN( u1_uk_n949 ) );
  OAI22_X1 u1_uk_U866 (.ZN( u1_K3_18 ) , .B2( u1_uk_n1325 ) , .A2( u1_uk_n1332 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U867 (.ZN( u1_K14_22 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1802 ) , .A2( u1_uk_n1840 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U868 (.ZN( u1_K10_5 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1625 ) , .A2( u1_uk_n1642 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U869 (.ZN( u1_K5_41 ) , .B2( u1_uk_n1418 ) , .A2( u1_uk_n1426 ) , .A1( u1_uk_n238 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U87 (.B2( u1_uk_K_r10_32 ) , .A2( u1_uk_K_r10_41 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n238 ) , .ZN( u1_uk_n524 ) );
  OAI22_X1 u1_uk_U870 (.ZN( u1_K15_22 ) , .B2( u1_uk_n1858 ) , .A2( u1_uk_n1872 ) , .A1( u1_uk_n209 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U871 (.ZN( u1_K6_22 ) , .B2( u1_uk_n1447 ) , .A2( u1_uk_n1452 ) , .A1( u1_uk_n294 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U872 (.ZN( u1_K15_23 ) , .B2( u1_uk_n1863 ) , .A2( u1_uk_n1881 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U873 (.ZN( u1_K14_23 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1802 ) , .B2( u1_uk_n1809 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U874 (.ZN( u1_K5_23 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1415 ) , .A2( u1_uk_n1424 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U875 (.ZN( u1_K13_34 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1768 ) , .A2( u1_uk_n1784 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U876 (.ZN( u1_K5_34 ) , .B1( u1_uk_n118 ) , .A2( u1_uk_n1401 ) , .B2( u1_uk_n1414 ) , .A1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U877 (.ZN( u1_K3_47 ) , .B2( u1_uk_n1327 ) , .A2( u1_uk_n1335 ) , .A1( u1_uk_n251 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U878 (.ZN( u1_K8_5 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1564 ) , .A2( u1_uk_n1570 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U879 (.ZN( u1_K6_5 ) , .B2( u1_uk_n1452 ) , .A2( u1_uk_n1456 ) , .A1( u1_uk_n188 ) , .B1( u1_uk_n27 ) );
  OAI21_X1 u1_uk_U88 (.ZN( u1_K11_23 ) , .B2( u1_uk_n1698 ) , .B1( u1_uk_n292 ) , .A( u1_uk_n408 ) );
  OAI22_X1 u1_uk_U880 (.ZN( u1_K12_10 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1718 ) , .A2( u1_uk_n1739 ) , .A1( u1_uk_n207 ) );
  OAI22_X1 u1_uk_U881 (.ZN( u1_K12_11 ) , .B1( u1_uk_n102 ) , .A2( u1_uk_n1713 ) , .B2( u1_uk_n1739 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U882 (.ZN( u1_K7_10 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1487 ) , .A2( u1_uk_n1517 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U883 (.B1( n116 ) , .ZN( u1_K4_11 ) , .B2( u1_uk_n1363 ) , .A2( u1_uk_n1391 ) , .A1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U884 (.ZN( u1_K3_10 ) , .B2( u1_uk_n1316 ) , .A2( u1_uk_n1321 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U885 (.ZN( u1_K15_45 ) , .B2( u1_uk_n1867 ) , .A2( u1_uk_n1885 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U886 (.ZN( u1_K13_45 ) , .B1( u1_uk_n162 ) , .B2( u1_uk_n1755 ) , .A2( u1_uk_n1793 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U887 (.ZN( u1_K12_43 ) , .B2( u1_uk_n1717 ) , .A2( u1_uk_n1737 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U888 (.ZN( u1_K6_45 ) , .B2( u1_uk_n1454 ) , .A2( u1_uk_n1459 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U889 (.ZN( u1_K3_30 ) , .B2( u1_uk_n1318 ) , .A2( u1_uk_n1344 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n94 ) );
  NAND2_X1 u1_uk_U89 (.A1( u1_uk_K_r9_27 ) , .A2( u1_uk_n298 ) , .ZN( u1_uk_n408 ) );
  OAI22_X1 u1_uk_U890 (.ZN( u1_K8_1 ) , .B1( u1_uk_n146 ) , .A2( u1_uk_n1532 ) , .B2( u1_uk_n1548 ) , .A1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U891 (.ZN( u1_K14_6 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1803 ) , .B2( u1_uk_n1810 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U892 (.ZN( u1_K10_3 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1633 ) , .A2( u1_uk_n1653 ) , .A1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U893 (.ZN( u1_K9_3 ) , .B1( u1_uk_n147 ) , .A2( u1_uk_n1573 ) , .B2( u1_uk_n1577 ) , .A1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U894 (.ZN( u1_K9_7 ) , .B1( u1_uk_n146 ) , .A2( u1_uk_n1574 ) , .B2( u1_uk_n1578 ) , .A1( u1_uk_n188 ) );
  OAI22_X1 u1_uk_U895 (.ZN( u1_K6_12 ) , .A2( u1_uk_n1440 ) , .B2( u1_uk_n1456 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U896 (.ZN( u1_K5_3 ) , .B2( u1_uk_n1404 ) , .A2( u1_uk_n1411 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U897 (.ZN( u1_K7_14 ) , .B2( u1_uk_n1492 ) , .A2( u1_uk_n1527 ) , .A1( u1_uk_n202 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U898 (.ZN( u1_K14_7 ) , .B2( u1_uk_n1816 ) , .A2( u1_uk_n1835 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U899 (.ZN( u1_K13_24 ) , .B2( u1_uk_n1756 ) , .A2( u1_uk_n1797 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n99 ) );
  INV_X1 u1_uk_U9 (.A( u1_uk_n209 ) , .ZN( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U90 (.ZN( u1_K10_23 ) , .B2( u1_uk_n1620 ) , .B1( u1_uk_n294 ) , .A( u1_uk_n313 ) );
  OAI22_X1 u1_uk_U900 (.ZN( u1_K6_24 ) , .B2( u1_uk_n1457 ) , .A2( u1_uk_n1461 ) , .A1( u1_uk_n286 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U901 (.ZN( u1_K15_13 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1844 ) , .B2( u1_uk_n1872 ) , .A1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U902 (.ZN( u1_K3_21 ) , .B2( u1_uk_n1321 ) , .A2( u1_uk_n1346 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U903 (.ZN( u1_K9_24 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1574 ) , .A2( u1_uk_n1616 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U904 (.ZN( u1_K5_19 ) , .A2( u1_uk_n1398 ) , .B2( u1_uk_n1435 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U905 (.ZN( u1_K5_24 ) , .B2( u1_uk_n1402 ) , .A2( u1_uk_n1427 ) , .B1( u1_uk_n145 ) , .A1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U906 (.ZN( u1_K2_24 ) , .A2( u1_uk_n1264 ) , .B2( u1_uk_n1279 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U907 (.ZN( u1_K16_21 ) , .B2( u1_uk_n1227 ) , .A2( u1_uk_n1234 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U908 (.ZN( u1_K8_21 ) , .B2( u1_uk_n1552 ) , .A2( u1_uk_n1558 ) , .B1( u1_uk_n17 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U909 (.ZN( u1_K16_24 ) , .B2( u1_uk_n1224 ) , .A2( u1_uk_n1229 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n63 ) );
  NAND2_X1 u1_uk_U91 (.A1( u1_uk_K_r8_13 ) , .A2( u1_uk_n271 ) , .ZN( u1_uk_n313 ) );
  OAI22_X1 u1_uk_U910 (.ZN( u1_K7_30 ) , .B2( u1_uk_n1490 ) , .A2( u1_uk_n1521 ) , .A1( u1_uk_n213 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U911 (.ZN( u1_K5_13 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1405 ) , .A2( u1_uk_n1436 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U912 (.ZN( u1_K5_14 ) , .B2( u1_uk_n1403 ) , .B1( u1_uk_n141 ) , .A2( u1_uk_n1410 ) , .A1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U913 (.ZN( u1_K4_14 ) , .B1( u1_uk_n110 ) , .B2( u1_uk_n1352 ) , .A2( u1_uk_n1378 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U914 (.ZN( u1_K3_13 ) , .B2( u1_uk_n1319 ) , .A2( u1_uk_n1324 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U915 (.ZN( u1_K4_36 ) , .B2( u1_uk_n1376 ) , .A2( u1_uk_n1381 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U916 (.ZN( u1_K2_17 ) , .A2( u1_uk_n1261 ) , .B2( u1_uk_n1277 ) , .A1( u1_uk_n291 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U917 (.ZN( u1_K6_30 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1438 ) , .A2( u1_uk_n1443 ) , .A1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U918 (.ZN( u1_K3_25 ) , .B2( u1_uk_n1309 ) , .A2( u1_uk_n1313 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U919 (.ZN( u1_K16_38 ) , .B2( u1_uk_n1240 ) , .A2( u1_uk_n1247 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U92 (.ZN( u1_K8_23 ) , .B2( u1_uk_n1543 ) , .A2( u1_uk_n1548 ) , .A1( u1_uk_n279 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U920 (.ZN( u1_K8_38 ) , .B1( u1_uk_n145 ) , .B2( u1_uk_n1560 ) , .A2( u1_uk_n1566 ) , .A1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U921 (.ZN( u1_K7_39 ) , .B2( u1_uk_n1516 ) , .A2( u1_uk_n1523 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n92 ) );
  OAI22_X1 u1_uk_U922 (.ZN( u1_K6_42 ) , .B1( u1_uk_n118 ) , .B2( u1_uk_n1468 ) , .A2( u1_uk_n1475 ) , .A1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U923 (.ZN( u1_K6_39 ) , .A2( u1_uk_n1441 ) , .B2( u1_uk_n1460 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U924 (.ZN( u1_K4_39 ) , .B2( u1_uk_n1351 ) , .A2( u1_uk_n1372 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n257 ) );
  OAI22_X1 u1_uk_U925 (.ZN( u1_K3_38 ) , .A2( u1_uk_n1314 ) , .B2( u1_uk_n1330 ) , .A1( u1_uk_n207 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U926 (.ZN( u1_K3_39 ) , .B2( u1_uk_n1338 ) , .A2( u1_uk_n1342 ) , .A1( u1_uk_n203 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U927 (.ZN( u1_K2_39 ) , .A2( u1_uk_n1266 ) , .B2( u1_uk_n1281 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U928 (.ZN( u1_K13_23 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1767 ) , .A2( u1_uk_n1797 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U929 (.ZN( u1_K9_23 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1584 ) , .A2( u1_uk_n1592 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U93 (.ZN( u1_K3_23 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1311 ) , .B2( u1_uk_n1316 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U930 (.ZN( u1_K9_47 ) , .B2( u1_uk_n1606 ) , .A2( u1_uk_n1613 ) , .A1( u1_uk_n163 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U931 (.ZN( u1_K12_16 ) , .A2( u1_uk_n1711 ) , .B2( u1_uk_n1723 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U932 (.ZN( u1_K11_16 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1692 ) , .A2( u1_uk_n1698 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U933 (.ZN( u1_K11_48 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1689 ) , .A2( u1_uk_n1696 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U934 (.ZN( u1_K11_6 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1699 ) , .A2( u1_uk_n1705 ) , .B1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U935 (.ZN( u1_K9_6 ) , .B2( u1_uk_n1585 ) , .A2( u1_uk_n1593 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U936 (.ZN( u1_K9_8 ) , .B2( u1_uk_n1603 ) , .A2( u1_uk_n1610 ) , .A1( u1_uk_n187 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U937 (.ZN( u1_K14_8 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1801 ) , .B2( u1_uk_n1819 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U938 (.ZN( u1_K12_18 ) , .A1( u1_uk_n164 ) , .A2( u1_uk_n1713 ) , .B2( u1_uk_n1751 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U939 (.ZN( u1_K14_20 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1813 ) , .A2( u1_uk_n1819 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U94 (.ZN( u1_K2_23 ) , .B2( u1_uk_n1278 ) , .A2( u1_uk_n1299 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U940 (.ZN( u1_K2_20 ) , .A2( u1_uk_n1263 ) , .B2( u1_uk_n1292 ) , .A1( u1_uk_n142 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U941 (.ZN( u1_K11_24 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1682 ) , .A2( u1_uk_n1687 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U942 (.ZN( u1_K14_14 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1834 ) , .A2( u1_uk_n1841 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U943 (.ZN( u1_K8_24 ) , .B2( u1_uk_n1530 ) , .A1( u1_uk_n155 ) , .A2( u1_uk_n1570 ) , .B1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U944 (.ZN( u1_K16_46 ) , .B2( u1_uk_n1219 ) , .A2( u1_uk_n1253 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U945 (.ZN( u1_K15_47 ) , .B2( u1_uk_n1854 ) , .A2( u1_uk_n1886 ) , .B1( u1_uk_n208 ) , .A1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U946 (.ZN( u1_K14_47 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1820 ) , .A2( u1_uk_n1830 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U947 (.ZN( u1_K10_46 ) , .B2( u1_uk_n1632 ) , .A2( u1_uk_n1641 ) , .B1( u1_uk_n279 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U948 (.ZN( u1_K10_34 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1618 ) , .A2( u1_uk_n1644 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U949 (.ZN( u1_K9_34 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1581 ) , .A2( u1_uk_n1588 ) , .B1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U95 (.ZN( u1_K11_41 ) , .B2( u1_uk_n1702 ) , .B1( u1_uk_n217 ) , .A( u1_uk_n467 ) );
  OAI22_X1 u1_uk_U950 (.ZN( u1_K6_46 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1443 ) , .B2( u1_uk_n1471 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U951 (.ZN( u1_K13_4 ) , .A1( u1_uk_n155 ) , .B2( u1_uk_n1762 ) , .A2( u1_uk_n1767 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U952 (.ZN( u1_K9_4 ) , .A1( u1_uk_n10 ) , .B2( u1_uk_n1579 ) , .A2( u1_uk_n1586 ) , .B1( u1_uk_n298 ) );
  OAI22_X1 u1_uk_U953 (.ZN( u1_K4_48 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1355 ) , .B2( u1_uk_n1383 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U954 (.ZN( u1_K2_48 ) , .B2( u1_uk_n1271 ) , .A2( u1_uk_n1286 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U955 (.ZN( u1_K10_8 ) , .A1( u1_uk_n129 ) , .A2( u1_uk_n1621 ) , .B2( u1_uk_n1635 ) , .B1( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U956 (.ZN( u1_K13_8 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1781 ) , .A2( u1_uk_n1787 ) , .B1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U957 (.ZN( u1_K6_20 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1439 ) , .B2( u1_uk_n1444 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U958 (.ZN( u1_K11_18 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1667 ) , .A2( u1_uk_n1673 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U959 (.ZN( u1_K14_18 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1818 ) , .A2( u1_uk_n1826 ) , .B1( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U96 (.A1( u1_uk_K_r9_31 ) , .A2( u1_uk_n203 ) , .ZN( u1_uk_n467 ) );
  OAI22_X1 u1_uk_U960 (.ZN( u1_K12_19 ) , .A1( u1_uk_n110 ) , .A2( u1_uk_n1712 ) , .B2( u1_uk_n1750 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U961 (.ZN( u1_K16_19 ) , .B2( u1_uk_n1220 ) , .A2( u1_uk_n1258 ) , .A1( u1_uk_n141 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U962 (.ZN( u1_K15_19 ) , .A1( u1_uk_n163 ) , .B2( u1_uk_n1851 ) , .A2( u1_uk_n1881 ) , .B1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U963 (.ZN( u1_K10_20 ) , .B2( u1_uk_n1629 ) , .A1( u1_uk_n163 ) , .A2( u1_uk_n1659 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U964 (.ZN( u1_K14_16 ) , .A1( u1_uk_n142 ) , .A2( u1_uk_n1804 ) , .B2( u1_uk_n1842 ) , .B1( u1_uk_n217 ) );
  OAI22_X1 u1_uk_U965 (.ZN( u1_K6_36 ) , .A1( u1_uk_n11 ) , .A2( u1_uk_n1441 ) , .B2( u1_uk_n1449 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U966 (.ZN( u1_K14_38 ) , .A2( u1_uk_n1807 ) , .B2( u1_uk_n1823 ) , .B1( u1_uk_n230 ) , .A1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U967 (.ZN( u1_K13_38 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1785 ) , .A2( u1_uk_n1791 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U968 (.ZN( u1_K2_38 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1276 ) , .A2( u1_uk_n1295 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U969 (.ZN( u1_K7_37 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1499 ) , .A2( u1_uk_n1523 ) , .B1( u1_uk_n250 ) );
  INV_X1 u1_uk_U97 (.ZN( u1_K9_41 ) , .A( u1_uk_n1166 ) );
  OAI22_X1 u1_uk_U970 (.ZN( u1_K2_37 ) , .A2( u1_uk_n1267 ) , .B2( u1_uk_n1294 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U971 (.ZN( u1_K9_40 ) , .B2( u1_uk_n1600 ) , .A2( u1_uk_n1606 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U972 (.ZN( u1_K5_40 ) , .B2( u1_uk_n1413 ) , .A2( u1_uk_n1430 ) , .A1( u1_uk_n162 ) , .B1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U973 (.ZN( u1_K2_22 ) , .B2( u1_uk_n1273 ) , .A2( u1_uk_n1290 ) , .B1( u1_uk_n222 ) , .A1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U974 (.ZN( u1_K8_45 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1528 ) , .A2( u1_uk_n1566 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U975 (.ZN( u1_K11_45 ) , .A1( u1_uk_n161 ) , .B2( u1_uk_n1677 ) , .A2( u1_uk_n1684 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U976 (.ZN( u1_K7_45 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1490 ) , .A2( u1_uk_n1507 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U977 (.ZN( u1_K6_43 ) , .A1( u1_uk_n129 ) , .B2( u1_uk_n1438 ) , .A2( u1_uk_n1477 ) , .B1( u1_uk_n203 ) );
  OAI22_X1 u1_uk_U978 (.ZN( u1_K4_45 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1351 ) , .A2( u1_uk_n1390 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U979 (.ZN( u1_K2_45 ) , .B2( u1_uk_n1282 ) , .A2( u1_uk_n1304 ) , .A1( u1_uk_n145 ) , .B1( u1_uk_n191 ) );
  AOI22_X1 u1_uk_U98 (.B2( u1_uk_K_r7_23 ) , .A2( u1_uk_K_r7_30 ) , .ZN( u1_uk_n1166 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U980 (.ZN( u1_K2_3 ) , .B2( u1_uk_n1269 ) , .A2( u1_uk_n1284 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U981 (.ZN( u1_K6_3 ) , .B2( u1_uk_n1447 ) , .A2( u1_uk_n1461 ) , .A1( u1_uk_n161 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U982 (.ZN( u1_K3_6 ) , .A2( u1_uk_n1312 ) , .B2( u1_uk_n1317 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U983 (.ZN( u1_K8_7 ) , .A2( u1_uk_n1530 ) , .B2( u1_uk_n1536 ) , .A1( u1_uk_n155 ) , .B1( u1_uk_n230 ) );
  OAI22_X1 u1_uk_U984 (.ZN( u1_K7_7 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1496 ) , .A2( u1_uk_n1518 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U985 (.ZN( u1_K3_7 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1323 ) , .A2( u1_uk_n1341 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U986 (.ZN( u1_K9_15 ) , .B2( u1_uk_n1577 ) , .A2( u1_uk_n1584 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U987 (.ZN( u1_K6_15 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1453 ) , .A2( u1_uk_n1465 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U988 (.ZN( u1_K6_25 ) , .B2( u1_uk_n1454 ) , .A2( u1_uk_n1470 ) , .A1( u1_uk_n17 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U989 (.ZN( u1_K14_25 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1800 ) , .A2( u1_uk_n1806 ) , .B1( u1_uk_n222 ) );
  INV_X1 u1_uk_U99 (.ZN( u1_K2_41 ) , .A( u1_uk_n1031 ) );
  OAI22_X1 u1_uk_U990 (.ZN( u1_K1_23 ) , .B2( u1_uk_n1197 ) , .A2( u1_uk_n1204 ) , .A1( u1_uk_n128 ) , .B1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U991 (.ZN( u1_K1_34 ) , .B2( u1_uk_n1174 ) , .A2( u1_uk_n1179 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n213 ) );
  OAI22_X1 u1_uk_U992 (.ZN( u1_K1_47 ) , .B2( u1_uk_n1172 ) , .A2( u1_uk_n1177 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U993 (.ZN( u1_K1_3 ) , .B2( u1_uk_n1184 ) , .A2( u1_uk_n1191 ) , .A1( u1_uk_n128 ) , .B1( u1_uk_n238 ) );
  OAI21_X1 u1_uk_U994 (.ZN( u1_K5_25 ) , .A( u1_uk_n1075 ) , .B2( u1_uk_n1413 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U995 (.A1( u1_uk_K_r3_35 ) , .ZN( u1_uk_n1075 ) , .A2( u1_uk_n63 ) );
  OAI21_X1 u1_uk_U996 (.ZN( u1_K7_22 ) , .A( u1_uk_n1111 ) , .B2( u1_uk_n1498 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U997 (.A1( u1_uk_K_r5_5 ) , .A2( u1_uk_n11 ) , .ZN( u1_uk_n1111 ) );
  OAI21_X1 u1_uk_U998 (.ZN( u1_K7_23 ) , .A( u1_uk_n1112 ) , .B2( u1_uk_n1483 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U999 (.A1( u1_uk_K_r5_13 ) , .ZN( u1_uk_n1112 ) , .A2( u1_uk_n17 ) );
  XOR2_X1 u2_U100 (.B( u2_L12_27 ) , .Z( u2_N442 ) , .A( u2_out13_27 ) );
  XOR2_X1 u2_U101 (.B( u2_L12_26 ) , .Z( u2_N441 ) , .A( u2_out13_26 ) );
  XOR2_X1 u2_U104 (.B( u2_L12_24 ) , .Z( u2_N439 ) , .A( u2_out13_24 ) );
  XOR2_X1 u2_U105 (.B( u2_L12_23 ) , .Z( u2_N438 ) , .A( u2_out13_23 ) );
  XOR2_X1 u2_U106 (.B( u2_L12_22 ) , .Z( u2_N437 ) , .A( u2_out13_22 ) );
  XOR2_X1 u2_U107 (.B( u2_L12_21 ) , .Z( u2_N436 ) , .A( u2_out13_21 ) );
  XOR2_X1 u2_U108 (.B( u2_L12_20 ) , .Z( u2_N435 ) , .A( u2_out13_20 ) );
  XOR2_X1 u2_U110 (.B( u2_L12_18 ) , .Z( u2_N433 ) , .A( u2_out13_18 ) );
  XOR2_X1 u2_U111 (.B( u2_L12_17 ) , .Z( u2_N432 ) , .A( u2_out13_17 ) );
  XOR2_X1 u2_U112 (.B( u2_L12_16 ) , .Z( u2_N431 ) , .A( u2_out13_16 ) );
  XOR2_X1 u2_U113 (.B( u2_L12_15 ) , .Z( u2_N430 ) , .A( u2_out13_15 ) );
  XOR2_X1 u2_U116 (.B( u2_L12_13 ) , .Z( u2_N428 ) , .A( u2_out13_13 ) );
  XOR2_X1 u2_U117 (.B( u2_L12_12 ) , .Z( u2_N427 ) , .A( u2_out13_12 ) );
  XOR2_X1 u2_U119 (.B( u2_L12_10 ) , .Z( u2_N425 ) , .A( u2_out13_10 ) );
  XOR2_X1 u2_U120 (.B( u2_L12_9 ) , .Z( u2_N424 ) , .A( u2_out13_9 ) );
  XOR2_X1 u2_U122 (.B( u2_L12_7 ) , .Z( u2_N422 ) , .A( u2_out13_7 ) );
  XOR2_X1 u2_U123 (.B( u2_L12_6 ) , .Z( u2_N421 ) , .A( u2_out13_6 ) );
  XOR2_X1 u2_U124 (.B( u2_L12_5 ) , .Z( u2_N420 ) , .A( u2_out13_5 ) );
  XOR2_X1 u2_U125 (.B( u2_L0_11 ) , .Z( u2_N42 ) , .A( u2_out1_11 ) );
  XOR2_X1 u2_U128 (.B( u2_L12_2 ) , .Z( u2_N417 ) , .A( u2_out13_2 ) );
  XOR2_X1 u2_U129 (.B( u2_L12_1 ) , .Z( u2_N416 ) , .A( u2_out13_1 ) );
  XOR2_X1 u2_U130 (.B( u2_L11_32 ) , .Z( u2_N415 ) , .A( u2_out12_32 ) );
  XOR2_X1 u2_U135 (.B( u2_L11_27 ) , .Z( u2_N410 ) , .A( u2_out12_27 ) );
  XOR2_X1 u2_U141 (.B( u2_L11_22 ) , .Z( u2_N405 ) , .A( u2_out12_22 ) );
  XOR2_X1 u2_U142 (.B( u2_L11_21 ) , .Z( u2_N404 ) , .A( u2_out12_21 ) );
  XOR2_X1 u2_U150 (.B( u2_L11_15 ) , .Z( u2_N398 ) , .A( u2_out12_15 ) );
  XOR2_X1 u2_U153 (.B( u2_L11_12 ) , .Z( u2_N395 ) , .A( u2_out12_12 ) );
  XOR2_X1 u2_U158 (.B( u2_L11_7 ) , .Z( u2_N390 ) , .A( u2_out12_7 ) );
  XOR2_X1 u2_U161 (.B( u2_L11_5 ) , .Z( u2_N388 ) , .A( u2_out12_5 ) );
  XOR2_X1 u2_U202 (.B( u2_L9_31 ) , .Z( u2_N350 ) , .A( u2_out10_31 ) );
  XOR2_X1 u2_U203 (.B( u2_L0_4 ) , .Z( u2_N35 ) , .A( u2_out1_4 ) );
  XOR2_X1 u2_U206 (.B( u2_L9_28 ) , .Z( u2_N347 ) , .A( u2_out10_28 ) );
  XOR2_X1 u2_U208 (.B( u2_L9_26 ) , .Z( u2_N345 ) , .A( u2_out10_26 ) );
  XOR2_X1 u2_U209 (.B( u2_L9_25 ) , .Z( u2_N344 ) , .A( u2_out10_25 ) );
  XOR2_X1 u2_U211 (.B( u2_L9_23 ) , .Z( u2_N342 ) , .A( u2_out10_23 ) );
  XOR2_X1 u2_U215 (.B( u2_L9_20 ) , .Z( u2_N339 ) , .A( u2_out10_20 ) );
  XOR2_X1 u2_U217 (.B( u2_L9_18 ) , .Z( u2_N337 ) , .A( u2_out10_18 ) );
  XOR2_X1 u2_U218 (.B( u2_L9_17 ) , .Z( u2_N336 ) , .A( u2_out10_17 ) );
  XOR2_X1 u2_U221 (.B( u2_L9_14 ) , .Z( u2_N333 ) , .A( u2_out10_14 ) );
  XOR2_X1 u2_U222 (.B( u2_L9_13 ) , .Z( u2_N332 ) , .A( u2_out10_13 ) );
  XOR2_X1 u2_U226 (.B( u2_L9_10 ) , .Z( u2_N329 ) , .A( u2_out10_10 ) );
  XOR2_X1 u2_U227 (.B( u2_L9_9 ) , .Z( u2_N328 ) , .A( u2_out10_9 ) );
  XOR2_X1 u2_U228 (.B( u2_L9_8 ) , .Z( u2_N327 ) , .A( u2_out10_8 ) );
  XOR2_X1 u2_U233 (.B( u2_L9_3 ) , .Z( u2_N322 ) , .A( u2_out10_3 ) );
  XOR2_X1 u2_U234 (.B( u2_L9_2 ) , .Z( u2_N321 ) , .A( u2_out10_2 ) );
  XOR2_X1 u2_U235 (.B( u2_L9_1 ) , .Z( u2_N320 ) , .A( u2_out10_1 ) );
  XOR2_X1 u2_U45 (.B( u2_L0_29 ) , .Z( u2_N60 ) , .A( u2_out1_29 ) );
  XOR2_X1 u2_U56 (.B( u2_L0_19 ) , .Z( u2_N50 ) , .A( u2_out1_19 ) );
  XOR2_X1 u2_U95 (.B( u2_L12_32 ) , .Z( u2_N447 ) , .A( u2_out13_32 ) );
  XOR2_X1 u2_U96 (.B( u2_L12_31 ) , .Z( u2_N446 ) , .A( u2_out13_31 ) );
  XOR2_X1 u2_U97 (.B( u2_L12_30 ) , .Z( u2_N445 ) , .A( u2_out13_30 ) );
  XOR2_X1 u2_U99 (.B( u2_L12_28 ) , .Z( u2_N443 ) , .A( u2_out13_28 ) );
  XOR2_X1 u2_u10_U1 (.B( u2_K11_9 ) , .A( u2_R9_6 ) , .Z( u2_u10_X_9 ) );
  XOR2_X1 u2_u10_U16 (.B( u2_K11_3 ) , .A( u2_R9_2 ) , .Z( u2_u10_X_3 ) );
  XOR2_X1 u2_u10_U2 (.B( u2_K11_8 ) , .A( u2_R9_5 ) , .Z( u2_u10_X_8 ) );
  XOR2_X1 u2_u10_U26 (.B( u2_K11_30 ) , .A( u2_R9_21 ) , .Z( u2_u10_X_30 ) );
  XOR2_X1 u2_u10_U27 (.B( u2_K11_2 ) , .A( u2_R9_1 ) , .Z( u2_u10_X_2 ) );
  XOR2_X1 u2_u10_U28 (.B( u2_K11_29 ) , .A( u2_R9_20 ) , .Z( u2_u10_X_29 ) );
  XOR2_X1 u2_u10_U29 (.B( u2_K11_28 ) , .A( u2_R9_19 ) , .Z( u2_u10_X_28 ) );
  XOR2_X1 u2_u10_U3 (.B( u2_K11_7 ) , .A( u2_R9_4 ) , .Z( u2_u10_X_7 ) );
  XOR2_X1 u2_u10_U30 (.B( u2_K11_27 ) , .A( u2_R9_18 ) , .Z( u2_u10_X_27 ) );
  XOR2_X1 u2_u10_U31 (.B( u2_K11_26 ) , .A( u2_R9_17 ) , .Z( u2_u10_X_26 ) );
  XOR2_X1 u2_u10_U32 (.B( u2_K11_25 ) , .A( u2_R9_16 ) , .Z( u2_u10_X_25 ) );
  XOR2_X1 u2_u10_U33 (.B( u2_K11_24 ) , .A( u2_R9_17 ) , .Z( u2_u10_X_24 ) );
  XOR2_X1 u2_u10_U34 (.B( u2_K11_23 ) , .A( u2_R9_16 ) , .Z( u2_u10_X_23 ) );
  XOR2_X1 u2_u10_U35 (.B( u2_K11_22 ) , .A( u2_R9_15 ) , .Z( u2_u10_X_22 ) );
  XOR2_X1 u2_u10_U36 (.B( u2_K11_21 ) , .A( u2_R9_14 ) , .Z( u2_u10_X_21 ) );
  XOR2_X1 u2_u10_U37 (.B( u2_K11_20 ) , .A( u2_R9_13 ) , .Z( u2_u10_X_20 ) );
  XOR2_X1 u2_u10_U38 (.B( u2_K11_1 ) , .A( u2_R9_32 ) , .Z( u2_u10_X_1 ) );
  XOR2_X1 u2_u10_U39 (.B( u2_K11_19 ) , .A( u2_R9_12 ) , .Z( u2_u10_X_19 ) );
  XOR2_X1 u2_u10_U4 (.B( u2_K11_6 ) , .A( u2_R9_5 ) , .Z( u2_u10_X_6 ) );
  XOR2_X1 u2_u10_U46 (.B( u2_K11_12 ) , .A( u2_R9_9 ) , .Z( u2_u10_X_12 ) );
  XOR2_X1 u2_u10_U47 (.B( u2_K11_11 ) , .A( u2_R9_8 ) , .Z( u2_u10_X_11 ) );
  XOR2_X1 u2_u10_U48 (.B( u2_K11_10 ) , .A( u2_R9_7 ) , .Z( u2_u10_X_10 ) );
  XOR2_X1 u2_u10_U5 (.B( u2_K11_5 ) , .A( u2_R9_4 ) , .Z( u2_u10_X_5 ) );
  XOR2_X1 u2_u10_U6 (.B( u2_K11_4 ) , .A( u2_R9_3 ) , .Z( u2_u10_X_4 ) );
  AND3_X1 u2_u10_u0_U10 (.A2( u2_u10_u0_n112 ) , .ZN( u2_u10_u0_n127 ) , .A3( u2_u10_u0_n130 ) , .A1( u2_u10_u0_n148 ) );
  NAND2_X1 u2_u10_u0_U11 (.ZN( u2_u10_u0_n113 ) , .A1( u2_u10_u0_n139 ) , .A2( u2_u10_u0_n149 ) );
  AND2_X1 u2_u10_u0_U12 (.ZN( u2_u10_u0_n107 ) , .A1( u2_u10_u0_n130 ) , .A2( u2_u10_u0_n140 ) );
  AND2_X1 u2_u10_u0_U13 (.A2( u2_u10_u0_n129 ) , .A1( u2_u10_u0_n130 ) , .ZN( u2_u10_u0_n151 ) );
  AND2_X1 u2_u10_u0_U14 (.A1( u2_u10_u0_n108 ) , .A2( u2_u10_u0_n125 ) , .ZN( u2_u10_u0_n145 ) );
  INV_X1 u2_u10_u0_U15 (.A( u2_u10_u0_n143 ) , .ZN( u2_u10_u0_n173 ) );
  NOR2_X1 u2_u10_u0_U16 (.A2( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n147 ) , .A1( u2_u10_u0_n160 ) );
  NOR2_X1 u2_u10_u0_U17 (.A1( u2_u10_u0_n163 ) , .A2( u2_u10_u0_n164 ) , .ZN( u2_u10_u0_n95 ) );
  AOI21_X1 u2_u10_u0_U18 (.B1( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n132 ) , .A( u2_u10_u0_n165 ) , .B2( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U19 (.A( u2_u10_u0_n142 ) , .ZN( u2_u10_u0_n165 ) );
  OAI221_X1 u2_u10_u0_U20 (.C1( u2_u10_u0_n121 ) , .ZN( u2_u10_u0_n122 ) , .B2( u2_u10_u0_n127 ) , .A( u2_u10_u0_n143 ) , .B1( u2_u10_u0_n144 ) , .C2( u2_u10_u0_n147 ) );
  OAI22_X1 u2_u10_u0_U21 (.B1( u2_u10_u0_n125 ) , .ZN( u2_u10_u0_n126 ) , .A1( u2_u10_u0_n138 ) , .A2( u2_u10_u0_n146 ) , .B2( u2_u10_u0_n147 ) );
  OAI22_X1 u2_u10_u0_U22 (.B1( u2_u10_u0_n131 ) , .A1( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n147 ) , .A2( u2_u10_u0_n90 ) , .ZN( u2_u10_u0_n91 ) );
  AND3_X1 u2_u10_u0_U23 (.A3( u2_u10_u0_n121 ) , .A2( u2_u10_u0_n125 ) , .A1( u2_u10_u0_n148 ) , .ZN( u2_u10_u0_n90 ) );
  NAND2_X1 u2_u10_u0_U24 (.A1( u2_u10_u0_n100 ) , .A2( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n125 ) );
  INV_X1 u2_u10_u0_U25 (.A( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n161 ) );
  NOR2_X1 u2_u10_u0_U26 (.A1( u2_u10_u0_n120 ) , .ZN( u2_u10_u0_n143 ) , .A2( u2_u10_u0_n167 ) );
  OAI221_X1 u2_u10_u0_U27 (.C1( u2_u10_u0_n112 ) , .ZN( u2_u10_u0_n120 ) , .B1( u2_u10_u0_n138 ) , .B2( u2_u10_u0_n141 ) , .C2( u2_u10_u0_n147 ) , .A( u2_u10_u0_n172 ) );
  AOI211_X1 u2_u10_u0_U28 (.B( u2_u10_u0_n115 ) , .A( u2_u10_u0_n116 ) , .C2( u2_u10_u0_n117 ) , .C1( u2_u10_u0_n118 ) , .ZN( u2_u10_u0_n119 ) );
  AOI22_X1 u2_u10_u0_U29 (.B2( u2_u10_u0_n109 ) , .A2( u2_u10_u0_n110 ) , .ZN( u2_u10_u0_n111 ) , .B1( u2_u10_u0_n118 ) , .A1( u2_u10_u0_n160 ) );
  INV_X1 u2_u10_u0_U3 (.A( u2_u10_u0_n113 ) , .ZN( u2_u10_u0_n166 ) );
  NAND2_X1 u2_u10_u0_U30 (.A1( u2_u10_u0_n100 ) , .ZN( u2_u10_u0_n129 ) , .A2( u2_u10_u0_n95 ) );
  INV_X1 u2_u10_u0_U31 (.A( u2_u10_u0_n118 ) , .ZN( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U32 (.ZN( u2_u10_u0_n104 ) , .B1( u2_u10_u0_n107 ) , .B2( u2_u10_u0_n141 ) , .A( u2_u10_u0_n144 ) );
  AOI21_X1 u2_u10_u0_U33 (.B1( u2_u10_u0_n127 ) , .B2( u2_u10_u0_n129 ) , .A( u2_u10_u0_n138 ) , .ZN( u2_u10_u0_n96 ) );
  AOI21_X1 u2_u10_u0_U34 (.ZN( u2_u10_u0_n116 ) , .B2( u2_u10_u0_n142 ) , .A( u2_u10_u0_n144 ) , .B1( u2_u10_u0_n166 ) );
  NAND2_X1 u2_u10_u0_U35 (.A2( u2_u10_u0_n100 ) , .A1( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n139 ) );
  NAND2_X1 u2_u10_u0_U36 (.A2( u2_u10_u0_n100 ) , .ZN( u2_u10_u0_n131 ) , .A1( u2_u10_u0_n92 ) );
  NAND2_X1 u2_u10_u0_U37 (.A1( u2_u10_u0_n101 ) , .A2( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n150 ) );
  INV_X1 u2_u10_u0_U38 (.A( u2_u10_u0_n138 ) , .ZN( u2_u10_u0_n160 ) );
  NAND2_X1 u2_u10_u0_U39 (.A1( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n128 ) , .A2( u2_u10_u0_n95 ) );
  AOI21_X1 u2_u10_u0_U4 (.B1( u2_u10_u0_n114 ) , .ZN( u2_u10_u0_n115 ) , .B2( u2_u10_u0_n129 ) , .A( u2_u10_u0_n161 ) );
  NAND2_X1 u2_u10_u0_U40 (.ZN( u2_u10_u0_n148 ) , .A1( u2_u10_u0_n93 ) , .A2( u2_u10_u0_n95 ) );
  NAND2_X1 u2_u10_u0_U41 (.A2( u2_u10_u0_n102 ) , .A1( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n149 ) );
  NAND2_X1 u2_u10_u0_U42 (.A2( u2_u10_u0_n102 ) , .ZN( u2_u10_u0_n114 ) , .A1( u2_u10_u0_n92 ) );
  NAND2_X1 u2_u10_u0_U43 (.A2( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n121 ) , .A1( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U44 (.ZN( u2_u10_u0_n172 ) , .A( u2_u10_u0_n88 ) );
  OAI222_X1 u2_u10_u0_U45 (.C1( u2_u10_u0_n108 ) , .A1( u2_u10_u0_n125 ) , .B2( u2_u10_u0_n128 ) , .B1( u2_u10_u0_n144 ) , .A2( u2_u10_u0_n158 ) , .C2( u2_u10_u0_n161 ) , .ZN( u2_u10_u0_n88 ) );
  NAND2_X1 u2_u10_u0_U46 (.ZN( u2_u10_u0_n112 ) , .A2( u2_u10_u0_n92 ) , .A1( u2_u10_u0_n93 ) );
  OR3_X1 u2_u10_u0_U47 (.A3( u2_u10_u0_n152 ) , .A2( u2_u10_u0_n153 ) , .A1( u2_u10_u0_n154 ) , .ZN( u2_u10_u0_n155 ) );
  AOI21_X1 u2_u10_u0_U48 (.A( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n145 ) , .B1( u2_u10_u0_n146 ) , .ZN( u2_u10_u0_n154 ) );
  AOI21_X1 u2_u10_u0_U49 (.B2( u2_u10_u0_n150 ) , .B1( u2_u10_u0_n151 ) , .ZN( u2_u10_u0_n152 ) , .A( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U5 (.B2( u2_u10_u0_n131 ) , .ZN( u2_u10_u0_n134 ) , .B1( u2_u10_u0_n151 ) , .A( u2_u10_u0_n158 ) );
  AOI21_X1 u2_u10_u0_U50 (.A( u2_u10_u0_n147 ) , .B2( u2_u10_u0_n148 ) , .B1( u2_u10_u0_n149 ) , .ZN( u2_u10_u0_n153 ) );
  INV_X1 u2_u10_u0_U51 (.ZN( u2_u10_u0_n171 ) , .A( u2_u10_u0_n99 ) );
  OAI211_X1 u2_u10_u0_U52 (.C2( u2_u10_u0_n140 ) , .C1( u2_u10_u0_n161 ) , .A( u2_u10_u0_n169 ) , .B( u2_u10_u0_n98 ) , .ZN( u2_u10_u0_n99 ) );
  AOI211_X1 u2_u10_u0_U53 (.C1( u2_u10_u0_n118 ) , .A( u2_u10_u0_n123 ) , .B( u2_u10_u0_n96 ) , .C2( u2_u10_u0_n97 ) , .ZN( u2_u10_u0_n98 ) );
  INV_X1 u2_u10_u0_U54 (.ZN( u2_u10_u0_n169 ) , .A( u2_u10_u0_n91 ) );
  NOR2_X1 u2_u10_u0_U55 (.A2( u2_u10_X_4 ) , .A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n118 ) );
  NOR2_X1 u2_u10_u0_U56 (.A2( u2_u10_X_2 ) , .ZN( u2_u10_u0_n103 ) , .A1( u2_u10_u0_n164 ) );
  NOR2_X1 u2_u10_u0_U57 (.A2( u2_u10_X_1 ) , .A1( u2_u10_X_2 ) , .ZN( u2_u10_u0_n92 ) );
  NOR2_X1 u2_u10_u0_U58 (.A2( u2_u10_X_1 ) , .ZN( u2_u10_u0_n101 ) , .A1( u2_u10_u0_n163 ) );
  NAND2_X1 u2_u10_u0_U59 (.A2( u2_u10_X_4 ) , .A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n144 ) );
  NOR2_X1 u2_u10_u0_U6 (.A1( u2_u10_u0_n108 ) , .ZN( u2_u10_u0_n123 ) , .A2( u2_u10_u0_n158 ) );
  NOR2_X1 u2_u10_u0_U60 (.A2( u2_u10_X_5 ) , .ZN( u2_u10_u0_n136 ) , .A1( u2_u10_u0_n159 ) );
  NAND2_X1 u2_u10_u0_U61 (.A1( u2_u10_X_5 ) , .ZN( u2_u10_u0_n138 ) , .A2( u2_u10_u0_n159 ) );
  AND2_X1 u2_u10_u0_U62 (.A2( u2_u10_X_3 ) , .A1( u2_u10_X_6 ) , .ZN( u2_u10_u0_n102 ) );
  AND2_X1 u2_u10_u0_U63 (.A1( u2_u10_X_6 ) , .A2( u2_u10_u0_n162 ) , .ZN( u2_u10_u0_n93 ) );
  INV_X1 u2_u10_u0_U64 (.A( u2_u10_X_4 ) , .ZN( u2_u10_u0_n159 ) );
  INV_X1 u2_u10_u0_U65 (.A( u2_u10_X_1 ) , .ZN( u2_u10_u0_n164 ) );
  INV_X1 u2_u10_u0_U66 (.A( u2_u10_X_2 ) , .ZN( u2_u10_u0_n163 ) );
  INV_X1 u2_u10_u0_U67 (.A( u2_u10_X_3 ) , .ZN( u2_u10_u0_n162 ) );
  INV_X1 u2_u10_u0_U68 (.A( u2_u10_u0_n126 ) , .ZN( u2_u10_u0_n168 ) );
  AOI211_X1 u2_u10_u0_U69 (.B( u2_u10_u0_n133 ) , .A( u2_u10_u0_n134 ) , .C2( u2_u10_u0_n135 ) , .C1( u2_u10_u0_n136 ) , .ZN( u2_u10_u0_n137 ) );
  OAI21_X1 u2_u10_u0_U7 (.B1( u2_u10_u0_n150 ) , .B2( u2_u10_u0_n158 ) , .A( u2_u10_u0_n172 ) , .ZN( u2_u10_u0_n89 ) );
  INV_X1 u2_u10_u0_U70 (.ZN( u2_u10_u0_n174 ) , .A( u2_u10_u0_n89 ) );
  AOI211_X1 u2_u10_u0_U71 (.B( u2_u10_u0_n104 ) , .A( u2_u10_u0_n105 ) , .ZN( u2_u10_u0_n106 ) , .C2( u2_u10_u0_n113 ) , .C1( u2_u10_u0_n160 ) );
  OR4_X1 u2_u10_u0_U72 (.ZN( u2_out10_17 ) , .A4( u2_u10_u0_n122 ) , .A2( u2_u10_u0_n123 ) , .A1( u2_u10_u0_n124 ) , .A3( u2_u10_u0_n170 ) );
  AOI21_X1 u2_u10_u0_U73 (.B2( u2_u10_u0_n107 ) , .ZN( u2_u10_u0_n124 ) , .B1( u2_u10_u0_n128 ) , .A( u2_u10_u0_n161 ) );
  INV_X1 u2_u10_u0_U74 (.A( u2_u10_u0_n111 ) , .ZN( u2_u10_u0_n170 ) );
  OR4_X1 u2_u10_u0_U75 (.ZN( u2_out10_31 ) , .A4( u2_u10_u0_n155 ) , .A2( u2_u10_u0_n156 ) , .A1( u2_u10_u0_n157 ) , .A3( u2_u10_u0_n173 ) );
  AOI21_X1 u2_u10_u0_U76 (.A( u2_u10_u0_n138 ) , .B2( u2_u10_u0_n139 ) , .B1( u2_u10_u0_n140 ) , .ZN( u2_u10_u0_n157 ) );
  AOI21_X1 u2_u10_u0_U77 (.B2( u2_u10_u0_n141 ) , .B1( u2_u10_u0_n142 ) , .ZN( u2_u10_u0_n156 ) , .A( u2_u10_u0_n161 ) );
  AOI21_X1 u2_u10_u0_U78 (.B1( u2_u10_u0_n132 ) , .ZN( u2_u10_u0_n133 ) , .A( u2_u10_u0_n144 ) , .B2( u2_u10_u0_n166 ) );
  OAI22_X1 u2_u10_u0_U79 (.ZN( u2_u10_u0_n105 ) , .A2( u2_u10_u0_n132 ) , .B1( u2_u10_u0_n146 ) , .A1( u2_u10_u0_n147 ) , .B2( u2_u10_u0_n161 ) );
  AND2_X1 u2_u10_u0_U8 (.A1( u2_u10_u0_n114 ) , .A2( u2_u10_u0_n121 ) , .ZN( u2_u10_u0_n146 ) );
  NAND2_X1 u2_u10_u0_U80 (.ZN( u2_u10_u0_n110 ) , .A2( u2_u10_u0_n132 ) , .A1( u2_u10_u0_n145 ) );
  INV_X1 u2_u10_u0_U81 (.A( u2_u10_u0_n119 ) , .ZN( u2_u10_u0_n167 ) );
  NAND2_X1 u2_u10_u0_U82 (.A2( u2_u10_u0_n103 ) , .ZN( u2_u10_u0_n140 ) , .A1( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U83 (.A1( u2_u10_u0_n101 ) , .ZN( u2_u10_u0_n130 ) , .A2( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U84 (.ZN( u2_u10_u0_n108 ) , .A1( u2_u10_u0_n92 ) , .A2( u2_u10_u0_n94 ) );
  NAND2_X1 u2_u10_u0_U85 (.ZN( u2_u10_u0_n142 ) , .A1( u2_u10_u0_n94 ) , .A2( u2_u10_u0_n95 ) );
  NOR2_X1 u2_u10_u0_U86 (.A2( u2_u10_X_6 ) , .ZN( u2_u10_u0_n100 ) , .A1( u2_u10_u0_n162 ) );
  NOR2_X1 u2_u10_u0_U87 (.A2( u2_u10_X_3 ) , .A1( u2_u10_X_6 ) , .ZN( u2_u10_u0_n94 ) );
  NAND3_X1 u2_u10_u0_U88 (.ZN( u2_out10_23 ) , .A3( u2_u10_u0_n137 ) , .A1( u2_u10_u0_n168 ) , .A2( u2_u10_u0_n171 ) );
  NAND3_X1 u2_u10_u0_U89 (.A3( u2_u10_u0_n127 ) , .A2( u2_u10_u0_n128 ) , .ZN( u2_u10_u0_n135 ) , .A1( u2_u10_u0_n150 ) );
  AND2_X1 u2_u10_u0_U9 (.A1( u2_u10_u0_n131 ) , .ZN( u2_u10_u0_n141 ) , .A2( u2_u10_u0_n150 ) );
  NAND3_X1 u2_u10_u0_U90 (.ZN( u2_u10_u0_n117 ) , .A3( u2_u10_u0_n132 ) , .A2( u2_u10_u0_n139 ) , .A1( u2_u10_u0_n148 ) );
  NAND3_X1 u2_u10_u0_U91 (.ZN( u2_u10_u0_n109 ) , .A2( u2_u10_u0_n114 ) , .A3( u2_u10_u0_n140 ) , .A1( u2_u10_u0_n149 ) );
  NAND3_X1 u2_u10_u0_U92 (.ZN( u2_out10_9 ) , .A3( u2_u10_u0_n106 ) , .A2( u2_u10_u0_n171 ) , .A1( u2_u10_u0_n174 ) );
  NAND3_X1 u2_u10_u0_U93 (.A2( u2_u10_u0_n128 ) , .A1( u2_u10_u0_n132 ) , .A3( u2_u10_u0_n146 ) , .ZN( u2_u10_u0_n97 ) );
  AOI21_X1 u2_u10_u1_U10 (.B2( u2_u10_u1_n155 ) , .B1( u2_u10_u1_n156 ) , .ZN( u2_u10_u1_n157 ) , .A( u2_u10_u1_n174 ) );
  NAND3_X1 u2_u10_u1_U100 (.ZN( u2_u10_u1_n113 ) , .A1( u2_u10_u1_n120 ) , .A3( u2_u10_u1_n133 ) , .A2( u2_u10_u1_n155 ) );
  NAND2_X1 u2_u10_u1_U11 (.ZN( u2_u10_u1_n140 ) , .A2( u2_u10_u1_n150 ) , .A1( u2_u10_u1_n155 ) );
  NAND2_X1 u2_u10_u1_U12 (.A1( u2_u10_u1_n131 ) , .ZN( u2_u10_u1_n147 ) , .A2( u2_u10_u1_n153 ) );
  AOI22_X1 u2_u10_u1_U13 (.B2( u2_u10_u1_n136 ) , .A2( u2_u10_u1_n137 ) , .ZN( u2_u10_u1_n143 ) , .A1( u2_u10_u1_n171 ) , .B1( u2_u10_u1_n173 ) );
  INV_X1 u2_u10_u1_U14 (.A( u2_u10_u1_n147 ) , .ZN( u2_u10_u1_n181 ) );
  INV_X1 u2_u10_u1_U15 (.A( u2_u10_u1_n139 ) , .ZN( u2_u10_u1_n174 ) );
  OR4_X1 u2_u10_u1_U16 (.A4( u2_u10_u1_n106 ) , .A3( u2_u10_u1_n107 ) , .ZN( u2_u10_u1_n108 ) , .A1( u2_u10_u1_n117 ) , .A2( u2_u10_u1_n184 ) );
  AOI21_X1 u2_u10_u1_U17 (.ZN( u2_u10_u1_n106 ) , .A( u2_u10_u1_n112 ) , .B1( u2_u10_u1_n154 ) , .B2( u2_u10_u1_n156 ) );
  AOI21_X1 u2_u10_u1_U18 (.ZN( u2_u10_u1_n107 ) , .B1( u2_u10_u1_n134 ) , .B2( u2_u10_u1_n149 ) , .A( u2_u10_u1_n174 ) );
  INV_X1 u2_u10_u1_U19 (.A( u2_u10_u1_n101 ) , .ZN( u2_u10_u1_n184 ) );
  INV_X1 u2_u10_u1_U20 (.A( u2_u10_u1_n112 ) , .ZN( u2_u10_u1_n171 ) );
  NAND2_X1 u2_u10_u1_U21 (.ZN( u2_u10_u1_n141 ) , .A1( u2_u10_u1_n153 ) , .A2( u2_u10_u1_n156 ) );
  AND2_X1 u2_u10_u1_U22 (.A1( u2_u10_u1_n123 ) , .ZN( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n161 ) );
  NAND2_X1 u2_u10_u1_U23 (.A2( u2_u10_u1_n115 ) , .A1( u2_u10_u1_n116 ) , .ZN( u2_u10_u1_n148 ) );
  NAND2_X1 u2_u10_u1_U24 (.A2( u2_u10_u1_n133 ) , .A1( u2_u10_u1_n135 ) , .ZN( u2_u10_u1_n159 ) );
  NAND2_X1 u2_u10_u1_U25 (.A2( u2_u10_u1_n115 ) , .A1( u2_u10_u1_n120 ) , .ZN( u2_u10_u1_n132 ) );
  INV_X1 u2_u10_u1_U26 (.A( u2_u10_u1_n154 ) , .ZN( u2_u10_u1_n178 ) );
  INV_X1 u2_u10_u1_U27 (.A( u2_u10_u1_n151 ) , .ZN( u2_u10_u1_n183 ) );
  AND2_X1 u2_u10_u1_U28 (.A1( u2_u10_u1_n129 ) , .A2( u2_u10_u1_n133 ) , .ZN( u2_u10_u1_n149 ) );
  INV_X1 u2_u10_u1_U29 (.A( u2_u10_u1_n131 ) , .ZN( u2_u10_u1_n180 ) );
  INV_X1 u2_u10_u1_U3 (.A( u2_u10_u1_n159 ) , .ZN( u2_u10_u1_n182 ) );
  OAI221_X1 u2_u10_u1_U30 (.A( u2_u10_u1_n119 ) , .C2( u2_u10_u1_n129 ) , .ZN( u2_u10_u1_n138 ) , .B2( u2_u10_u1_n152 ) , .C1( u2_u10_u1_n174 ) , .B1( u2_u10_u1_n187 ) );
  INV_X1 u2_u10_u1_U31 (.A( u2_u10_u1_n148 ) , .ZN( u2_u10_u1_n187 ) );
  AOI211_X1 u2_u10_u1_U32 (.B( u2_u10_u1_n117 ) , .A( u2_u10_u1_n118 ) , .ZN( u2_u10_u1_n119 ) , .C2( u2_u10_u1_n146 ) , .C1( u2_u10_u1_n159 ) );
  NOR2_X1 u2_u10_u1_U33 (.A1( u2_u10_u1_n168 ) , .A2( u2_u10_u1_n176 ) , .ZN( u2_u10_u1_n98 ) );
  OAI21_X1 u2_u10_u1_U34 (.B2( u2_u10_u1_n123 ) , .ZN( u2_u10_u1_n145 ) , .B1( u2_u10_u1_n160 ) , .A( u2_u10_u1_n185 ) );
  INV_X1 u2_u10_u1_U35 (.A( u2_u10_u1_n122 ) , .ZN( u2_u10_u1_n185 ) );
  AOI21_X1 u2_u10_u1_U36 (.B2( u2_u10_u1_n120 ) , .B1( u2_u10_u1_n121 ) , .ZN( u2_u10_u1_n122 ) , .A( u2_u10_u1_n128 ) );
  NAND2_X1 u2_u10_u1_U37 (.A1( u2_u10_u1_n128 ) , .ZN( u2_u10_u1_n146 ) , .A2( u2_u10_u1_n160 ) );
  NAND2_X1 u2_u10_u1_U38 (.A2( u2_u10_u1_n112 ) , .ZN( u2_u10_u1_n139 ) , .A1( u2_u10_u1_n152 ) );
  NAND2_X1 u2_u10_u1_U39 (.A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n156 ) , .A2( u2_u10_u1_n99 ) );
  AOI221_X1 u2_u10_u1_U4 (.A( u2_u10_u1_n138 ) , .C2( u2_u10_u1_n139 ) , .C1( u2_u10_u1_n140 ) , .B2( u2_u10_u1_n141 ) , .ZN( u2_u10_u1_n142 ) , .B1( u2_u10_u1_n175 ) );
  AOI221_X1 u2_u10_u1_U40 (.B1( u2_u10_u1_n140 ) , .ZN( u2_u10_u1_n167 ) , .B2( u2_u10_u1_n172 ) , .C2( u2_u10_u1_n175 ) , .C1( u2_u10_u1_n178 ) , .A( u2_u10_u1_n188 ) );
  INV_X1 u2_u10_u1_U41 (.ZN( u2_u10_u1_n188 ) , .A( u2_u10_u1_n97 ) );
  AOI211_X1 u2_u10_u1_U42 (.A( u2_u10_u1_n118 ) , .C1( u2_u10_u1_n132 ) , .C2( u2_u10_u1_n139 ) , .B( u2_u10_u1_n96 ) , .ZN( u2_u10_u1_n97 ) );
  AOI21_X1 u2_u10_u1_U43 (.B2( u2_u10_u1_n121 ) , .B1( u2_u10_u1_n135 ) , .A( u2_u10_u1_n152 ) , .ZN( u2_u10_u1_n96 ) );
  NOR2_X1 u2_u10_u1_U44 (.ZN( u2_u10_u1_n117 ) , .A1( u2_u10_u1_n121 ) , .A2( u2_u10_u1_n160 ) );
  AOI21_X1 u2_u10_u1_U45 (.A( u2_u10_u1_n128 ) , .B2( u2_u10_u1_n129 ) , .ZN( u2_u10_u1_n130 ) , .B1( u2_u10_u1_n150 ) );
  NAND2_X1 u2_u10_u1_U46 (.ZN( u2_u10_u1_n112 ) , .A1( u2_u10_u1_n169 ) , .A2( u2_u10_u1_n170 ) );
  NAND2_X1 u2_u10_u1_U47 (.ZN( u2_u10_u1_n129 ) , .A2( u2_u10_u1_n95 ) , .A1( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U48 (.A1( u2_u10_u1_n102 ) , .ZN( u2_u10_u1_n154 ) , .A2( u2_u10_u1_n99 ) );
  NAND2_X1 u2_u10_u1_U49 (.A2( u2_u10_u1_n100 ) , .ZN( u2_u10_u1_n135 ) , .A1( u2_u10_u1_n99 ) );
  AOI211_X1 u2_u10_u1_U5 (.ZN( u2_u10_u1_n124 ) , .A( u2_u10_u1_n138 ) , .C2( u2_u10_u1_n139 ) , .B( u2_u10_u1_n145 ) , .C1( u2_u10_u1_n147 ) );
  AOI21_X1 u2_u10_u1_U50 (.A( u2_u10_u1_n152 ) , .B2( u2_u10_u1_n153 ) , .B1( u2_u10_u1_n154 ) , .ZN( u2_u10_u1_n158 ) );
  INV_X1 u2_u10_u1_U51 (.A( u2_u10_u1_n160 ) , .ZN( u2_u10_u1_n175 ) );
  NAND2_X1 u2_u10_u1_U52 (.A1( u2_u10_u1_n100 ) , .ZN( u2_u10_u1_n116 ) , .A2( u2_u10_u1_n95 ) );
  NAND2_X1 u2_u10_u1_U53 (.A1( u2_u10_u1_n102 ) , .ZN( u2_u10_u1_n131 ) , .A2( u2_u10_u1_n95 ) );
  NAND2_X1 u2_u10_u1_U54 (.A2( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n121 ) , .A1( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U55 (.A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n153 ) , .A2( u2_u10_u1_n98 ) );
  NAND2_X1 u2_u10_u1_U56 (.A2( u2_u10_u1_n104 ) , .A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n133 ) );
  NAND2_X1 u2_u10_u1_U57 (.ZN( u2_u10_u1_n150 ) , .A2( u2_u10_u1_n98 ) , .A1( u2_u10_u1_n99 ) );
  NAND2_X1 u2_u10_u1_U58 (.A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n155 ) , .A2( u2_u10_u1_n95 ) );
  OAI21_X1 u2_u10_u1_U59 (.ZN( u2_u10_u1_n109 ) , .B1( u2_u10_u1_n129 ) , .B2( u2_u10_u1_n160 ) , .A( u2_u10_u1_n167 ) );
  AOI22_X1 u2_u10_u1_U6 (.B2( u2_u10_u1_n113 ) , .A2( u2_u10_u1_n114 ) , .ZN( u2_u10_u1_n125 ) , .A1( u2_u10_u1_n171 ) , .B1( u2_u10_u1_n173 ) );
  NAND2_X1 u2_u10_u1_U60 (.A2( u2_u10_u1_n100 ) , .A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n120 ) );
  NAND2_X1 u2_u10_u1_U61 (.A1( u2_u10_u1_n102 ) , .A2( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n115 ) );
  NAND2_X1 u2_u10_u1_U62 (.A2( u2_u10_u1_n100 ) , .A1( u2_u10_u1_n104 ) , .ZN( u2_u10_u1_n151 ) );
  NAND2_X1 u2_u10_u1_U63 (.A2( u2_u10_u1_n103 ) , .A1( u2_u10_u1_n105 ) , .ZN( u2_u10_u1_n161 ) );
  INV_X1 u2_u10_u1_U64 (.A( u2_u10_u1_n152 ) , .ZN( u2_u10_u1_n173 ) );
  INV_X1 u2_u10_u1_U65 (.A( u2_u10_u1_n128 ) , .ZN( u2_u10_u1_n172 ) );
  NAND2_X1 u2_u10_u1_U66 (.A2( u2_u10_u1_n102 ) , .A1( u2_u10_u1_n103 ) , .ZN( u2_u10_u1_n123 ) );
  AOI211_X1 u2_u10_u1_U67 (.B( u2_u10_u1_n162 ) , .A( u2_u10_u1_n163 ) , .C2( u2_u10_u1_n164 ) , .ZN( u2_u10_u1_n165 ) , .C1( u2_u10_u1_n171 ) );
  AOI21_X1 u2_u10_u1_U68 (.A( u2_u10_u1_n160 ) , .B2( u2_u10_u1_n161 ) , .ZN( u2_u10_u1_n162 ) , .B1( u2_u10_u1_n182 ) );
  OR2_X1 u2_u10_u1_U69 (.A2( u2_u10_u1_n157 ) , .A1( u2_u10_u1_n158 ) , .ZN( u2_u10_u1_n163 ) );
  NAND2_X1 u2_u10_u1_U7 (.ZN( u2_u10_u1_n114 ) , .A1( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n156 ) );
  NOR2_X1 u2_u10_u1_U70 (.A2( u2_u10_X_7 ) , .A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n95 ) );
  NOR2_X1 u2_u10_u1_U71 (.A1( u2_u10_X_12 ) , .A2( u2_u10_X_9 ) , .ZN( u2_u10_u1_n100 ) );
  NOR2_X1 u2_u10_u1_U72 (.A2( u2_u10_X_8 ) , .A1( u2_u10_u1_n177 ) , .ZN( u2_u10_u1_n99 ) );
  NOR2_X1 u2_u10_u1_U73 (.A2( u2_u10_X_12 ) , .ZN( u2_u10_u1_n102 ) , .A1( u2_u10_u1_n176 ) );
  NOR2_X1 u2_u10_u1_U74 (.A2( u2_u10_X_9 ) , .ZN( u2_u10_u1_n105 ) , .A1( u2_u10_u1_n168 ) );
  NAND2_X1 u2_u10_u1_U75 (.A1( u2_u10_X_10 ) , .ZN( u2_u10_u1_n160 ) , .A2( u2_u10_u1_n169 ) );
  NAND2_X1 u2_u10_u1_U76 (.A2( u2_u10_X_10 ) , .A1( u2_u10_X_11 ) , .ZN( u2_u10_u1_n152 ) );
  NAND2_X1 u2_u10_u1_U77 (.A1( u2_u10_X_11 ) , .ZN( u2_u10_u1_n128 ) , .A2( u2_u10_u1_n170 ) );
  AND2_X1 u2_u10_u1_U78 (.A2( u2_u10_X_7 ) , .A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n104 ) );
  AND2_X1 u2_u10_u1_U79 (.A1( u2_u10_X_8 ) , .ZN( u2_u10_u1_n103 ) , .A2( u2_u10_u1_n177 ) );
  NOR2_X1 u2_u10_u1_U8 (.A1( u2_u10_u1_n112 ) , .A2( u2_u10_u1_n116 ) , .ZN( u2_u10_u1_n118 ) );
  INV_X1 u2_u10_u1_U80 (.A( u2_u10_X_10 ) , .ZN( u2_u10_u1_n170 ) );
  INV_X1 u2_u10_u1_U81 (.A( u2_u10_X_9 ) , .ZN( u2_u10_u1_n176 ) );
  INV_X1 u2_u10_u1_U82 (.A( u2_u10_X_11 ) , .ZN( u2_u10_u1_n169 ) );
  INV_X1 u2_u10_u1_U83 (.A( u2_u10_X_12 ) , .ZN( u2_u10_u1_n168 ) );
  INV_X1 u2_u10_u1_U84 (.A( u2_u10_X_7 ) , .ZN( u2_u10_u1_n177 ) );
  NAND4_X1 u2_u10_u1_U85 (.ZN( u2_out10_28 ) , .A4( u2_u10_u1_n124 ) , .A3( u2_u10_u1_n125 ) , .A2( u2_u10_u1_n126 ) , .A1( u2_u10_u1_n127 ) );
  OAI21_X1 u2_u10_u1_U86 (.ZN( u2_u10_u1_n127 ) , .B2( u2_u10_u1_n139 ) , .B1( u2_u10_u1_n175 ) , .A( u2_u10_u1_n183 ) );
  OAI21_X1 u2_u10_u1_U87 (.ZN( u2_u10_u1_n126 ) , .B2( u2_u10_u1_n140 ) , .A( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n178 ) );
  NAND4_X1 u2_u10_u1_U88 (.ZN( u2_out10_18 ) , .A4( u2_u10_u1_n165 ) , .A3( u2_u10_u1_n166 ) , .A1( u2_u10_u1_n167 ) , .A2( u2_u10_u1_n186 ) );
  AOI22_X1 u2_u10_u1_U89 (.B2( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n147 ) , .A2( u2_u10_u1_n148 ) , .ZN( u2_u10_u1_n166 ) , .A1( u2_u10_u1_n172 ) );
  OAI21_X1 u2_u10_u1_U9 (.ZN( u2_u10_u1_n101 ) , .B1( u2_u10_u1_n141 ) , .A( u2_u10_u1_n146 ) , .B2( u2_u10_u1_n183 ) );
  INV_X1 u2_u10_u1_U90 (.A( u2_u10_u1_n145 ) , .ZN( u2_u10_u1_n186 ) );
  NAND4_X1 u2_u10_u1_U91 (.ZN( u2_out10_2 ) , .A4( u2_u10_u1_n142 ) , .A3( u2_u10_u1_n143 ) , .A2( u2_u10_u1_n144 ) , .A1( u2_u10_u1_n179 ) );
  OAI21_X1 u2_u10_u1_U92 (.B2( u2_u10_u1_n132 ) , .ZN( u2_u10_u1_n144 ) , .A( u2_u10_u1_n146 ) , .B1( u2_u10_u1_n180 ) );
  INV_X1 u2_u10_u1_U93 (.A( u2_u10_u1_n130 ) , .ZN( u2_u10_u1_n179 ) );
  OR4_X1 u2_u10_u1_U94 (.ZN( u2_out10_13 ) , .A4( u2_u10_u1_n108 ) , .A3( u2_u10_u1_n109 ) , .A2( u2_u10_u1_n110 ) , .A1( u2_u10_u1_n111 ) );
  AOI21_X1 u2_u10_u1_U95 (.ZN( u2_u10_u1_n111 ) , .A( u2_u10_u1_n128 ) , .B2( u2_u10_u1_n131 ) , .B1( u2_u10_u1_n135 ) );
  AOI21_X1 u2_u10_u1_U96 (.ZN( u2_u10_u1_n110 ) , .A( u2_u10_u1_n116 ) , .B1( u2_u10_u1_n152 ) , .B2( u2_u10_u1_n160 ) );
  NAND3_X1 u2_u10_u1_U97 (.A3( u2_u10_u1_n149 ) , .A2( u2_u10_u1_n150 ) , .A1( u2_u10_u1_n151 ) , .ZN( u2_u10_u1_n164 ) );
  NAND3_X1 u2_u10_u1_U98 (.A3( u2_u10_u1_n134 ) , .A2( u2_u10_u1_n135 ) , .ZN( u2_u10_u1_n136 ) , .A1( u2_u10_u1_n151 ) );
  NAND3_X1 u2_u10_u1_U99 (.A1( u2_u10_u1_n133 ) , .ZN( u2_u10_u1_n137 ) , .A2( u2_u10_u1_n154 ) , .A3( u2_u10_u1_n181 ) );
  OAI22_X1 u2_u10_u3_U10 (.B1( u2_u10_u3_n113 ) , .A2( u2_u10_u3_n135 ) , .A1( u2_u10_u3_n150 ) , .B2( u2_u10_u3_n164 ) , .ZN( u2_u10_u3_n98 ) );
  OAI211_X1 u2_u10_u3_U11 (.B( u2_u10_u3_n106 ) , .ZN( u2_u10_u3_n119 ) , .C2( u2_u10_u3_n128 ) , .C1( u2_u10_u3_n167 ) , .A( u2_u10_u3_n181 ) );
  AOI221_X1 u2_u10_u3_U12 (.C1( u2_u10_u3_n105 ) , .ZN( u2_u10_u3_n106 ) , .A( u2_u10_u3_n131 ) , .B2( u2_u10_u3_n132 ) , .C2( u2_u10_u3_n133 ) , .B1( u2_u10_u3_n169 ) );
  INV_X1 u2_u10_u3_U13 (.ZN( u2_u10_u3_n181 ) , .A( u2_u10_u3_n98 ) );
  NAND2_X1 u2_u10_u3_U14 (.ZN( u2_u10_u3_n105 ) , .A2( u2_u10_u3_n130 ) , .A1( u2_u10_u3_n155 ) );
  AOI22_X1 u2_u10_u3_U15 (.B1( u2_u10_u3_n115 ) , .A2( u2_u10_u3_n116 ) , .ZN( u2_u10_u3_n123 ) , .B2( u2_u10_u3_n133 ) , .A1( u2_u10_u3_n169 ) );
  NAND2_X1 u2_u10_u3_U16 (.ZN( u2_u10_u3_n116 ) , .A2( u2_u10_u3_n151 ) , .A1( u2_u10_u3_n182 ) );
  NOR2_X1 u2_u10_u3_U17 (.ZN( u2_u10_u3_n126 ) , .A2( u2_u10_u3_n150 ) , .A1( u2_u10_u3_n164 ) );
  AOI21_X1 u2_u10_u3_U18 (.ZN( u2_u10_u3_n112 ) , .B2( u2_u10_u3_n146 ) , .B1( u2_u10_u3_n155 ) , .A( u2_u10_u3_n167 ) );
  NAND2_X1 u2_u10_u3_U19 (.A1( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n142 ) , .A2( u2_u10_u3_n164 ) );
  NAND2_X1 u2_u10_u3_U20 (.ZN( u2_u10_u3_n132 ) , .A2( u2_u10_u3_n152 ) , .A1( u2_u10_u3_n156 ) );
  AND2_X1 u2_u10_u3_U21 (.A2( u2_u10_u3_n113 ) , .A1( u2_u10_u3_n114 ) , .ZN( u2_u10_u3_n151 ) );
  INV_X1 u2_u10_u3_U22 (.A( u2_u10_u3_n133 ) , .ZN( u2_u10_u3_n165 ) );
  INV_X1 u2_u10_u3_U23 (.A( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n170 ) );
  NAND2_X1 u2_u10_u3_U24 (.A1( u2_u10_u3_n107 ) , .A2( u2_u10_u3_n108 ) , .ZN( u2_u10_u3_n140 ) );
  NAND2_X1 u2_u10_u3_U25 (.ZN( u2_u10_u3_n117 ) , .A1( u2_u10_u3_n124 ) , .A2( u2_u10_u3_n148 ) );
  NAND2_X1 u2_u10_u3_U26 (.ZN( u2_u10_u3_n143 ) , .A1( u2_u10_u3_n165 ) , .A2( u2_u10_u3_n167 ) );
  INV_X1 u2_u10_u3_U27 (.A( u2_u10_u3_n130 ) , .ZN( u2_u10_u3_n177 ) );
  INV_X1 u2_u10_u3_U28 (.A( u2_u10_u3_n128 ) , .ZN( u2_u10_u3_n176 ) );
  INV_X1 u2_u10_u3_U29 (.A( u2_u10_u3_n155 ) , .ZN( u2_u10_u3_n174 ) );
  INV_X1 u2_u10_u3_U3 (.A( u2_u10_u3_n129 ) , .ZN( u2_u10_u3_n183 ) );
  INV_X1 u2_u10_u3_U30 (.A( u2_u10_u3_n139 ) , .ZN( u2_u10_u3_n185 ) );
  NOR2_X1 u2_u10_u3_U31 (.ZN( u2_u10_u3_n135 ) , .A2( u2_u10_u3_n141 ) , .A1( u2_u10_u3_n169 ) );
  OAI222_X1 u2_u10_u3_U32 (.C2( u2_u10_u3_n107 ) , .A2( u2_u10_u3_n108 ) , .B1( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n138 ) , .B2( u2_u10_u3_n146 ) , .C1( u2_u10_u3_n154 ) , .A1( u2_u10_u3_n164 ) );
  NOR4_X1 u2_u10_u3_U33 (.A4( u2_u10_u3_n157 ) , .A3( u2_u10_u3_n158 ) , .A2( u2_u10_u3_n159 ) , .A1( u2_u10_u3_n160 ) , .ZN( u2_u10_u3_n161 ) );
  AOI21_X1 u2_u10_u3_U34 (.B2( u2_u10_u3_n152 ) , .B1( u2_u10_u3_n153 ) , .ZN( u2_u10_u3_n158 ) , .A( u2_u10_u3_n164 ) );
  AOI21_X1 u2_u10_u3_U35 (.A( u2_u10_u3_n154 ) , .B2( u2_u10_u3_n155 ) , .B1( u2_u10_u3_n156 ) , .ZN( u2_u10_u3_n157 ) );
  AOI21_X1 u2_u10_u3_U36 (.A( u2_u10_u3_n149 ) , .B2( u2_u10_u3_n150 ) , .B1( u2_u10_u3_n151 ) , .ZN( u2_u10_u3_n159 ) );
  AOI211_X1 u2_u10_u3_U37 (.ZN( u2_u10_u3_n109 ) , .A( u2_u10_u3_n119 ) , .C2( u2_u10_u3_n129 ) , .B( u2_u10_u3_n138 ) , .C1( u2_u10_u3_n141 ) );
  AOI211_X1 u2_u10_u3_U38 (.B( u2_u10_u3_n119 ) , .A( u2_u10_u3_n120 ) , .C2( u2_u10_u3_n121 ) , .ZN( u2_u10_u3_n122 ) , .C1( u2_u10_u3_n179 ) );
  INV_X1 u2_u10_u3_U39 (.A( u2_u10_u3_n156 ) , .ZN( u2_u10_u3_n179 ) );
  INV_X1 u2_u10_u3_U4 (.A( u2_u10_u3_n140 ) , .ZN( u2_u10_u3_n182 ) );
  OAI22_X1 u2_u10_u3_U40 (.B1( u2_u10_u3_n118 ) , .ZN( u2_u10_u3_n120 ) , .A1( u2_u10_u3_n135 ) , .B2( u2_u10_u3_n154 ) , .A2( u2_u10_u3_n178 ) );
  AND3_X1 u2_u10_u3_U41 (.ZN( u2_u10_u3_n118 ) , .A2( u2_u10_u3_n124 ) , .A1( u2_u10_u3_n144 ) , .A3( u2_u10_u3_n152 ) );
  INV_X1 u2_u10_u3_U42 (.A( u2_u10_u3_n121 ) , .ZN( u2_u10_u3_n164 ) );
  NAND2_X1 u2_u10_u3_U43 (.ZN( u2_u10_u3_n133 ) , .A1( u2_u10_u3_n154 ) , .A2( u2_u10_u3_n164 ) );
  OAI211_X1 u2_u10_u3_U44 (.B( u2_u10_u3_n127 ) , .ZN( u2_u10_u3_n139 ) , .C1( u2_u10_u3_n150 ) , .C2( u2_u10_u3_n154 ) , .A( u2_u10_u3_n184 ) );
  INV_X1 u2_u10_u3_U45 (.A( u2_u10_u3_n125 ) , .ZN( u2_u10_u3_n184 ) );
  AOI221_X1 u2_u10_u3_U46 (.A( u2_u10_u3_n126 ) , .ZN( u2_u10_u3_n127 ) , .C2( u2_u10_u3_n132 ) , .C1( u2_u10_u3_n169 ) , .B2( u2_u10_u3_n170 ) , .B1( u2_u10_u3_n174 ) );
  OAI22_X1 u2_u10_u3_U47 (.A1( u2_u10_u3_n124 ) , .ZN( u2_u10_u3_n125 ) , .B2( u2_u10_u3_n145 ) , .A2( u2_u10_u3_n165 ) , .B1( u2_u10_u3_n167 ) );
  NOR2_X1 u2_u10_u3_U48 (.A1( u2_u10_u3_n113 ) , .ZN( u2_u10_u3_n131 ) , .A2( u2_u10_u3_n154 ) );
  NAND2_X1 u2_u10_u3_U49 (.A1( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n150 ) , .A2( u2_u10_u3_n99 ) );
  INV_X1 u2_u10_u3_U5 (.A( u2_u10_u3_n117 ) , .ZN( u2_u10_u3_n178 ) );
  NAND2_X1 u2_u10_u3_U50 (.A2( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n155 ) , .A1( u2_u10_u3_n97 ) );
  INV_X1 u2_u10_u3_U51 (.A( u2_u10_u3_n141 ) , .ZN( u2_u10_u3_n167 ) );
  AOI21_X1 u2_u10_u3_U52 (.B2( u2_u10_u3_n114 ) , .B1( u2_u10_u3_n146 ) , .A( u2_u10_u3_n154 ) , .ZN( u2_u10_u3_n94 ) );
  AOI21_X1 u2_u10_u3_U53 (.ZN( u2_u10_u3_n110 ) , .B2( u2_u10_u3_n142 ) , .B1( u2_u10_u3_n186 ) , .A( u2_u10_u3_n95 ) );
  INV_X1 u2_u10_u3_U54 (.A( u2_u10_u3_n145 ) , .ZN( u2_u10_u3_n186 ) );
  AOI21_X1 u2_u10_u3_U55 (.B1( u2_u10_u3_n124 ) , .A( u2_u10_u3_n149 ) , .B2( u2_u10_u3_n155 ) , .ZN( u2_u10_u3_n95 ) );
  INV_X1 u2_u10_u3_U56 (.A( u2_u10_u3_n149 ) , .ZN( u2_u10_u3_n169 ) );
  NAND2_X1 u2_u10_u3_U57 (.ZN( u2_u10_u3_n124 ) , .A1( u2_u10_u3_n96 ) , .A2( u2_u10_u3_n97 ) );
  NAND2_X1 u2_u10_u3_U58 (.A2( u2_u10_u3_n100 ) , .ZN( u2_u10_u3_n146 ) , .A1( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U59 (.A1( u2_u10_u3_n101 ) , .ZN( u2_u10_u3_n145 ) , .A2( u2_u10_u3_n99 ) );
  AOI221_X1 u2_u10_u3_U6 (.A( u2_u10_u3_n131 ) , .C2( u2_u10_u3_n132 ) , .C1( u2_u10_u3_n133 ) , .ZN( u2_u10_u3_n134 ) , .B1( u2_u10_u3_n143 ) , .B2( u2_u10_u3_n177 ) );
  NAND2_X1 u2_u10_u3_U60 (.A1( u2_u10_u3_n100 ) , .ZN( u2_u10_u3_n156 ) , .A2( u2_u10_u3_n99 ) );
  NAND2_X1 u2_u10_u3_U61 (.A2( u2_u10_u3_n101 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n148 ) );
  NAND2_X1 u2_u10_u3_U62 (.A1( u2_u10_u3_n100 ) , .A2( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n128 ) );
  NAND2_X1 u2_u10_u3_U63 (.A2( u2_u10_u3_n101 ) , .A1( u2_u10_u3_n102 ) , .ZN( u2_u10_u3_n152 ) );
  NAND2_X1 u2_u10_u3_U64 (.A2( u2_u10_u3_n101 ) , .ZN( u2_u10_u3_n114 ) , .A1( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U65 (.ZN( u2_u10_u3_n107 ) , .A1( u2_u10_u3_n97 ) , .A2( u2_u10_u3_n99 ) );
  NAND2_X1 u2_u10_u3_U66 (.A2( u2_u10_u3_n100 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n113 ) );
  NAND2_X1 u2_u10_u3_U67 (.A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n153 ) , .A2( u2_u10_u3_n97 ) );
  NAND2_X1 u2_u10_u3_U68 (.A2( u2_u10_u3_n103 ) , .A1( u2_u10_u3_n104 ) , .ZN( u2_u10_u3_n130 ) );
  NAND2_X1 u2_u10_u3_U69 (.A2( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n144 ) , .A1( u2_u10_u3_n96 ) );
  OAI22_X1 u2_u10_u3_U7 (.B2( u2_u10_u3_n147 ) , .A2( u2_u10_u3_n148 ) , .ZN( u2_u10_u3_n160 ) , .B1( u2_u10_u3_n165 ) , .A1( u2_u10_u3_n168 ) );
  NAND2_X1 u2_u10_u3_U70 (.A1( u2_u10_u3_n102 ) , .A2( u2_u10_u3_n103 ) , .ZN( u2_u10_u3_n108 ) );
  NOR2_X1 u2_u10_u3_U71 (.A2( u2_u10_X_19 ) , .A1( u2_u10_X_20 ) , .ZN( u2_u10_u3_n99 ) );
  NOR2_X1 u2_u10_u3_U72 (.A2( u2_u10_X_21 ) , .A1( u2_u10_X_24 ) , .ZN( u2_u10_u3_n103 ) );
  NOR2_X1 u2_u10_u3_U73 (.A2( u2_u10_X_24 ) , .A1( u2_u10_u3_n171 ) , .ZN( u2_u10_u3_n97 ) );
  NOR2_X1 u2_u10_u3_U74 (.A2( u2_u10_X_23 ) , .ZN( u2_u10_u3_n141 ) , .A1( u2_u10_u3_n166 ) );
  NOR2_X1 u2_u10_u3_U75 (.A2( u2_u10_X_19 ) , .A1( u2_u10_u3_n172 ) , .ZN( u2_u10_u3_n96 ) );
  NAND2_X1 u2_u10_u3_U76 (.A1( u2_u10_X_22 ) , .A2( u2_u10_X_23 ) , .ZN( u2_u10_u3_n154 ) );
  NAND2_X1 u2_u10_u3_U77 (.A1( u2_u10_X_23 ) , .ZN( u2_u10_u3_n149 ) , .A2( u2_u10_u3_n166 ) );
  NOR2_X1 u2_u10_u3_U78 (.A2( u2_u10_X_22 ) , .A1( u2_u10_X_23 ) , .ZN( u2_u10_u3_n121 ) );
  AND2_X1 u2_u10_u3_U79 (.A1( u2_u10_X_24 ) , .ZN( u2_u10_u3_n101 ) , .A2( u2_u10_u3_n171 ) );
  AND3_X1 u2_u10_u3_U8 (.A3( u2_u10_u3_n144 ) , .A2( u2_u10_u3_n145 ) , .A1( u2_u10_u3_n146 ) , .ZN( u2_u10_u3_n147 ) );
  AND2_X1 u2_u10_u3_U80 (.A1( u2_u10_X_19 ) , .ZN( u2_u10_u3_n102 ) , .A2( u2_u10_u3_n172 ) );
  AND2_X1 u2_u10_u3_U81 (.A1( u2_u10_X_21 ) , .A2( u2_u10_X_24 ) , .ZN( u2_u10_u3_n100 ) );
  AND2_X1 u2_u10_u3_U82 (.A2( u2_u10_X_19 ) , .A1( u2_u10_X_20 ) , .ZN( u2_u10_u3_n104 ) );
  INV_X1 u2_u10_u3_U83 (.A( u2_u10_X_22 ) , .ZN( u2_u10_u3_n166 ) );
  INV_X1 u2_u10_u3_U84 (.A( u2_u10_X_21 ) , .ZN( u2_u10_u3_n171 ) );
  INV_X1 u2_u10_u3_U85 (.A( u2_u10_X_20 ) , .ZN( u2_u10_u3_n172 ) );
  OR4_X1 u2_u10_u3_U86 (.ZN( u2_out10_10 ) , .A4( u2_u10_u3_n136 ) , .A3( u2_u10_u3_n137 ) , .A1( u2_u10_u3_n138 ) , .A2( u2_u10_u3_n139 ) );
  OAI222_X1 u2_u10_u3_U87 (.C1( u2_u10_u3_n128 ) , .ZN( u2_u10_u3_n137 ) , .B1( u2_u10_u3_n148 ) , .A2( u2_u10_u3_n150 ) , .B2( u2_u10_u3_n154 ) , .C2( u2_u10_u3_n164 ) , .A1( u2_u10_u3_n167 ) );
  OAI221_X1 u2_u10_u3_U88 (.A( u2_u10_u3_n134 ) , .B2( u2_u10_u3_n135 ) , .ZN( u2_u10_u3_n136 ) , .C1( u2_u10_u3_n149 ) , .B1( u2_u10_u3_n151 ) , .C2( u2_u10_u3_n183 ) );
  NAND4_X1 u2_u10_u3_U89 (.ZN( u2_out10_26 ) , .A4( u2_u10_u3_n109 ) , .A3( u2_u10_u3_n110 ) , .A2( u2_u10_u3_n111 ) , .A1( u2_u10_u3_n173 ) );
  INV_X1 u2_u10_u3_U9 (.A( u2_u10_u3_n143 ) , .ZN( u2_u10_u3_n168 ) );
  INV_X1 u2_u10_u3_U90 (.ZN( u2_u10_u3_n173 ) , .A( u2_u10_u3_n94 ) );
  OAI21_X1 u2_u10_u3_U91 (.ZN( u2_u10_u3_n111 ) , .B2( u2_u10_u3_n117 ) , .A( u2_u10_u3_n133 ) , .B1( u2_u10_u3_n176 ) );
  NAND4_X1 u2_u10_u3_U92 (.ZN( u2_out10_20 ) , .A4( u2_u10_u3_n122 ) , .A3( u2_u10_u3_n123 ) , .A1( u2_u10_u3_n175 ) , .A2( u2_u10_u3_n180 ) );
  INV_X1 u2_u10_u3_U93 (.A( u2_u10_u3_n126 ) , .ZN( u2_u10_u3_n180 ) );
  INV_X1 u2_u10_u3_U94 (.A( u2_u10_u3_n112 ) , .ZN( u2_u10_u3_n175 ) );
  NAND4_X1 u2_u10_u3_U95 (.ZN( u2_out10_1 ) , .A4( u2_u10_u3_n161 ) , .A3( u2_u10_u3_n162 ) , .A2( u2_u10_u3_n163 ) , .A1( u2_u10_u3_n185 ) );
  NAND2_X1 u2_u10_u3_U96 (.ZN( u2_u10_u3_n163 ) , .A2( u2_u10_u3_n170 ) , .A1( u2_u10_u3_n176 ) );
  AOI22_X1 u2_u10_u3_U97 (.B2( u2_u10_u3_n140 ) , .B1( u2_u10_u3_n141 ) , .A2( u2_u10_u3_n142 ) , .ZN( u2_u10_u3_n162 ) , .A1( u2_u10_u3_n177 ) );
  NAND3_X1 u2_u10_u3_U98 (.A1( u2_u10_u3_n114 ) , .ZN( u2_u10_u3_n115 ) , .A2( u2_u10_u3_n145 ) , .A3( u2_u10_u3_n153 ) );
  NAND3_X1 u2_u10_u3_U99 (.ZN( u2_u10_u3_n129 ) , .A2( u2_u10_u3_n144 ) , .A1( u2_u10_u3_n153 ) , .A3( u2_u10_u3_n182 ) );
  AOI21_X1 u2_u10_u4_U10 (.ZN( u2_u10_u4_n106 ) , .B2( u2_u10_u4_n146 ) , .B1( u2_u10_u4_n158 ) , .A( u2_u10_u4_n170 ) );
  AOI21_X1 u2_u10_u4_U11 (.ZN( u2_u10_u4_n108 ) , .B2( u2_u10_u4_n134 ) , .B1( u2_u10_u4_n155 ) , .A( u2_u10_u4_n156 ) );
  AOI21_X1 u2_u10_u4_U12 (.ZN( u2_u10_u4_n109 ) , .A( u2_u10_u4_n153 ) , .B1( u2_u10_u4_n159 ) , .B2( u2_u10_u4_n184 ) );
  AOI211_X1 u2_u10_u4_U13 (.B( u2_u10_u4_n136 ) , .A( u2_u10_u4_n137 ) , .C2( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n139 ) , .C1( u2_u10_u4_n182 ) );
  OAI22_X1 u2_u10_u4_U14 (.B2( u2_u10_u4_n135 ) , .ZN( u2_u10_u4_n137 ) , .B1( u2_u10_u4_n153 ) , .A1( u2_u10_u4_n155 ) , .A2( u2_u10_u4_n171 ) );
  AND3_X1 u2_u10_u4_U15 (.A2( u2_u10_u4_n134 ) , .ZN( u2_u10_u4_n135 ) , .A3( u2_u10_u4_n145 ) , .A1( u2_u10_u4_n157 ) );
  NAND2_X1 u2_u10_u4_U16 (.ZN( u2_u10_u4_n132 ) , .A2( u2_u10_u4_n170 ) , .A1( u2_u10_u4_n173 ) );
  AOI21_X1 u2_u10_u4_U17 (.B2( u2_u10_u4_n160 ) , .B1( u2_u10_u4_n161 ) , .ZN( u2_u10_u4_n162 ) , .A( u2_u10_u4_n170 ) );
  AOI21_X1 u2_u10_u4_U18 (.ZN( u2_u10_u4_n107 ) , .B2( u2_u10_u4_n143 ) , .A( u2_u10_u4_n174 ) , .B1( u2_u10_u4_n184 ) );
  AOI21_X1 u2_u10_u4_U19 (.B2( u2_u10_u4_n158 ) , .B1( u2_u10_u4_n159 ) , .ZN( u2_u10_u4_n163 ) , .A( u2_u10_u4_n174 ) );
  AOI21_X1 u2_u10_u4_U20 (.A( u2_u10_u4_n153 ) , .B2( u2_u10_u4_n154 ) , .B1( u2_u10_u4_n155 ) , .ZN( u2_u10_u4_n165 ) );
  AOI21_X1 u2_u10_u4_U21 (.A( u2_u10_u4_n156 ) , .B2( u2_u10_u4_n157 ) , .ZN( u2_u10_u4_n164 ) , .B1( u2_u10_u4_n184 ) );
  INV_X1 u2_u10_u4_U22 (.A( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n170 ) );
  AND2_X1 u2_u10_u4_U23 (.A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n155 ) , .A1( u2_u10_u4_n160 ) );
  INV_X1 u2_u10_u4_U24 (.A( u2_u10_u4_n156 ) , .ZN( u2_u10_u4_n175 ) );
  NAND2_X1 u2_u10_u4_U25 (.A2( u2_u10_u4_n118 ) , .ZN( u2_u10_u4_n131 ) , .A1( u2_u10_u4_n147 ) );
  NAND2_X1 u2_u10_u4_U26 (.A1( u2_u10_u4_n119 ) , .A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n130 ) );
  NAND2_X1 u2_u10_u4_U27 (.ZN( u2_u10_u4_n117 ) , .A2( u2_u10_u4_n118 ) , .A1( u2_u10_u4_n148 ) );
  NAND2_X1 u2_u10_u4_U28 (.ZN( u2_u10_u4_n129 ) , .A1( u2_u10_u4_n134 ) , .A2( u2_u10_u4_n148 ) );
  AND3_X1 u2_u10_u4_U29 (.A1( u2_u10_u4_n119 ) , .A2( u2_u10_u4_n143 ) , .A3( u2_u10_u4_n154 ) , .ZN( u2_u10_u4_n161 ) );
  NOR2_X1 u2_u10_u4_U3 (.ZN( u2_u10_u4_n121 ) , .A1( u2_u10_u4_n181 ) , .A2( u2_u10_u4_n182 ) );
  AND2_X1 u2_u10_u4_U30 (.A1( u2_u10_u4_n145 ) , .A2( u2_u10_u4_n147 ) , .ZN( u2_u10_u4_n159 ) );
  OR3_X1 u2_u10_u4_U31 (.A3( u2_u10_u4_n114 ) , .A2( u2_u10_u4_n115 ) , .A1( u2_u10_u4_n116 ) , .ZN( u2_u10_u4_n136 ) );
  AOI21_X1 u2_u10_u4_U32 (.A( u2_u10_u4_n113 ) , .ZN( u2_u10_u4_n116 ) , .B2( u2_u10_u4_n173 ) , .B1( u2_u10_u4_n174 ) );
  AOI21_X1 u2_u10_u4_U33 (.ZN( u2_u10_u4_n115 ) , .B2( u2_u10_u4_n145 ) , .B1( u2_u10_u4_n146 ) , .A( u2_u10_u4_n156 ) );
  OAI22_X1 u2_u10_u4_U34 (.ZN( u2_u10_u4_n114 ) , .A2( u2_u10_u4_n121 ) , .B1( u2_u10_u4_n160 ) , .B2( u2_u10_u4_n170 ) , .A1( u2_u10_u4_n171 ) );
  INV_X1 u2_u10_u4_U35 (.A( u2_u10_u4_n158 ) , .ZN( u2_u10_u4_n182 ) );
  INV_X1 u2_u10_u4_U36 (.ZN( u2_u10_u4_n181 ) , .A( u2_u10_u4_n96 ) );
  INV_X1 u2_u10_u4_U37 (.A( u2_u10_u4_n144 ) , .ZN( u2_u10_u4_n179 ) );
  INV_X1 u2_u10_u4_U38 (.A( u2_u10_u4_n157 ) , .ZN( u2_u10_u4_n178 ) );
  NAND2_X1 u2_u10_u4_U39 (.A2( u2_u10_u4_n154 ) , .A1( u2_u10_u4_n96 ) , .ZN( u2_u10_u4_n97 ) );
  INV_X1 u2_u10_u4_U4 (.A( u2_u10_u4_n117 ) , .ZN( u2_u10_u4_n184 ) );
  INV_X1 u2_u10_u4_U40 (.A( u2_u10_u4_n143 ) , .ZN( u2_u10_u4_n183 ) );
  NOR2_X1 u2_u10_u4_U41 (.ZN( u2_u10_u4_n138 ) , .A1( u2_u10_u4_n168 ) , .A2( u2_u10_u4_n169 ) );
  NOR2_X1 u2_u10_u4_U42 (.A1( u2_u10_u4_n150 ) , .A2( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n153 ) );
  NOR2_X1 u2_u10_u4_U43 (.A2( u2_u10_u4_n128 ) , .A1( u2_u10_u4_n138 ) , .ZN( u2_u10_u4_n156 ) );
  AOI22_X1 u2_u10_u4_U44 (.B2( u2_u10_u4_n122 ) , .A1( u2_u10_u4_n123 ) , .ZN( u2_u10_u4_n124 ) , .B1( u2_u10_u4_n128 ) , .A2( u2_u10_u4_n172 ) );
  INV_X1 u2_u10_u4_U45 (.A( u2_u10_u4_n153 ) , .ZN( u2_u10_u4_n172 ) );
  NAND2_X1 u2_u10_u4_U46 (.A2( u2_u10_u4_n120 ) , .ZN( u2_u10_u4_n123 ) , .A1( u2_u10_u4_n161 ) );
  AOI22_X1 u2_u10_u4_U47 (.B2( u2_u10_u4_n132 ) , .A2( u2_u10_u4_n133 ) , .ZN( u2_u10_u4_n140 ) , .A1( u2_u10_u4_n150 ) , .B1( u2_u10_u4_n179 ) );
  NAND2_X1 u2_u10_u4_U48 (.ZN( u2_u10_u4_n133 ) , .A2( u2_u10_u4_n146 ) , .A1( u2_u10_u4_n154 ) );
  NAND2_X1 u2_u10_u4_U49 (.A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n154 ) , .A2( u2_u10_u4_n98 ) );
  INV_X1 u2_u10_u4_U5 (.ZN( u2_u10_u4_n186 ) , .A( u2_u10_u4_n95 ) );
  NAND2_X1 u2_u10_u4_U50 (.A1( u2_u10_u4_n101 ) , .ZN( u2_u10_u4_n158 ) , .A2( u2_u10_u4_n99 ) );
  AOI21_X1 u2_u10_u4_U51 (.ZN( u2_u10_u4_n127 ) , .A( u2_u10_u4_n136 ) , .B2( u2_u10_u4_n150 ) , .B1( u2_u10_u4_n180 ) );
  INV_X1 u2_u10_u4_U52 (.A( u2_u10_u4_n160 ) , .ZN( u2_u10_u4_n180 ) );
  NAND2_X1 u2_u10_u4_U53 (.A2( u2_u10_u4_n104 ) , .A1( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n146 ) );
  NAND2_X1 u2_u10_u4_U54 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n160 ) );
  NAND2_X1 u2_u10_u4_U55 (.ZN( u2_u10_u4_n134 ) , .A1( u2_u10_u4_n98 ) , .A2( u2_u10_u4_n99 ) );
  NAND2_X1 u2_u10_u4_U56 (.A1( u2_u10_u4_n103 ) , .A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n143 ) );
  NAND2_X1 u2_u10_u4_U57 (.A2( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n145 ) , .A1( u2_u10_u4_n98 ) );
  NAND2_X1 u2_u10_u4_U58 (.A1( u2_u10_u4_n100 ) , .A2( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n120 ) );
  NAND2_X1 u2_u10_u4_U59 (.A1( u2_u10_u4_n102 ) , .A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n148 ) );
  OAI221_X1 u2_u10_u4_U6 (.C1( u2_u10_u4_n134 ) , .B1( u2_u10_u4_n158 ) , .B2( u2_u10_u4_n171 ) , .C2( u2_u10_u4_n173 ) , .A( u2_u10_u4_n94 ) , .ZN( u2_u10_u4_n95 ) );
  NAND2_X1 u2_u10_u4_U60 (.A2( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n157 ) );
  INV_X1 u2_u10_u4_U61 (.A( u2_u10_u4_n150 ) , .ZN( u2_u10_u4_n173 ) );
  INV_X1 u2_u10_u4_U62 (.A( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n171 ) );
  NAND2_X1 u2_u10_u4_U63 (.A1( u2_u10_u4_n100 ) , .ZN( u2_u10_u4_n118 ) , .A2( u2_u10_u4_n99 ) );
  NAND2_X1 u2_u10_u4_U64 (.A2( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n144 ) );
  NAND2_X1 u2_u10_u4_U65 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n105 ) , .ZN( u2_u10_u4_n96 ) );
  INV_X1 u2_u10_u4_U66 (.A( u2_u10_u4_n128 ) , .ZN( u2_u10_u4_n174 ) );
  NAND2_X1 u2_u10_u4_U67 (.A2( u2_u10_u4_n102 ) , .ZN( u2_u10_u4_n119 ) , .A1( u2_u10_u4_n98 ) );
  NAND2_X1 u2_u10_u4_U68 (.A2( u2_u10_u4_n101 ) , .A1( u2_u10_u4_n103 ) , .ZN( u2_u10_u4_n147 ) );
  NAND2_X1 u2_u10_u4_U69 (.A2( u2_u10_u4_n104 ) , .ZN( u2_u10_u4_n113 ) , .A1( u2_u10_u4_n99 ) );
  AOI222_X1 u2_u10_u4_U7 (.B2( u2_u10_u4_n132 ) , .A1( u2_u10_u4_n138 ) , .C2( u2_u10_u4_n175 ) , .A2( u2_u10_u4_n179 ) , .C1( u2_u10_u4_n181 ) , .B1( u2_u10_u4_n185 ) , .ZN( u2_u10_u4_n94 ) );
  NOR2_X1 u2_u10_u4_U70 (.A2( u2_u10_X_28 ) , .ZN( u2_u10_u4_n150 ) , .A1( u2_u10_u4_n168 ) );
  NOR2_X1 u2_u10_u4_U71 (.A2( u2_u10_X_29 ) , .ZN( u2_u10_u4_n152 ) , .A1( u2_u10_u4_n169 ) );
  NOR2_X1 u2_u10_u4_U72 (.A2( u2_u10_X_30 ) , .ZN( u2_u10_u4_n105 ) , .A1( u2_u10_u4_n176 ) );
  NOR2_X1 u2_u10_u4_U73 (.A2( u2_u10_X_26 ) , .ZN( u2_u10_u4_n100 ) , .A1( u2_u10_u4_n177 ) );
  NOR2_X1 u2_u10_u4_U74 (.A2( u2_u10_X_28 ) , .A1( u2_u10_X_29 ) , .ZN( u2_u10_u4_n128 ) );
  NOR2_X1 u2_u10_u4_U75 (.A2( u2_u10_X_27 ) , .A1( u2_u10_X_30 ) , .ZN( u2_u10_u4_n102 ) );
  NOR2_X1 u2_u10_u4_U76 (.A2( u2_u10_X_25 ) , .A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n98 ) );
  AND2_X1 u2_u10_u4_U77 (.A2( u2_u10_X_25 ) , .A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n104 ) );
  AND2_X1 u2_u10_u4_U78 (.A1( u2_u10_X_30 ) , .A2( u2_u10_u4_n176 ) , .ZN( u2_u10_u4_n99 ) );
  AND2_X1 u2_u10_u4_U79 (.A1( u2_u10_X_26 ) , .ZN( u2_u10_u4_n101 ) , .A2( u2_u10_u4_n177 ) );
  INV_X1 u2_u10_u4_U8 (.A( u2_u10_u4_n113 ) , .ZN( u2_u10_u4_n185 ) );
  AND2_X1 u2_u10_u4_U80 (.A1( u2_u10_X_27 ) , .A2( u2_u10_X_30 ) , .ZN( u2_u10_u4_n103 ) );
  INV_X1 u2_u10_u4_U81 (.A( u2_u10_X_28 ) , .ZN( u2_u10_u4_n169 ) );
  INV_X1 u2_u10_u4_U82 (.A( u2_u10_X_29 ) , .ZN( u2_u10_u4_n168 ) );
  INV_X1 u2_u10_u4_U83 (.A( u2_u10_X_25 ) , .ZN( u2_u10_u4_n177 ) );
  INV_X1 u2_u10_u4_U84 (.A( u2_u10_X_27 ) , .ZN( u2_u10_u4_n176 ) );
  NAND4_X1 u2_u10_u4_U85 (.ZN( u2_out10_25 ) , .A4( u2_u10_u4_n139 ) , .A3( u2_u10_u4_n140 ) , .A2( u2_u10_u4_n141 ) , .A1( u2_u10_u4_n142 ) );
  OAI21_X1 u2_u10_u4_U86 (.A( u2_u10_u4_n128 ) , .B2( u2_u10_u4_n129 ) , .B1( u2_u10_u4_n130 ) , .ZN( u2_u10_u4_n142 ) );
  OAI21_X1 u2_u10_u4_U87 (.B2( u2_u10_u4_n131 ) , .ZN( u2_u10_u4_n141 ) , .A( u2_u10_u4_n175 ) , .B1( u2_u10_u4_n183 ) );
  NAND4_X1 u2_u10_u4_U88 (.ZN( u2_out10_14 ) , .A4( u2_u10_u4_n124 ) , .A3( u2_u10_u4_n125 ) , .A2( u2_u10_u4_n126 ) , .A1( u2_u10_u4_n127 ) );
  AOI22_X1 u2_u10_u4_U89 (.B2( u2_u10_u4_n117 ) , .ZN( u2_u10_u4_n126 ) , .A1( u2_u10_u4_n129 ) , .B1( u2_u10_u4_n152 ) , .A2( u2_u10_u4_n175 ) );
  NOR4_X1 u2_u10_u4_U9 (.A4( u2_u10_u4_n106 ) , .A3( u2_u10_u4_n107 ) , .A2( u2_u10_u4_n108 ) , .A1( u2_u10_u4_n109 ) , .ZN( u2_u10_u4_n110 ) );
  AOI22_X1 u2_u10_u4_U90 (.ZN( u2_u10_u4_n125 ) , .B2( u2_u10_u4_n131 ) , .A2( u2_u10_u4_n132 ) , .B1( u2_u10_u4_n138 ) , .A1( u2_u10_u4_n178 ) );
  NAND4_X1 u2_u10_u4_U91 (.ZN( u2_out10_8 ) , .A4( u2_u10_u4_n110 ) , .A3( u2_u10_u4_n111 ) , .A2( u2_u10_u4_n112 ) , .A1( u2_u10_u4_n186 ) );
  NAND2_X1 u2_u10_u4_U92 (.ZN( u2_u10_u4_n112 ) , .A2( u2_u10_u4_n130 ) , .A1( u2_u10_u4_n150 ) );
  AOI22_X1 u2_u10_u4_U93 (.ZN( u2_u10_u4_n111 ) , .B2( u2_u10_u4_n132 ) , .A1( u2_u10_u4_n152 ) , .B1( u2_u10_u4_n178 ) , .A2( u2_u10_u4_n97 ) );
  AOI22_X1 u2_u10_u4_U94 (.B2( u2_u10_u4_n149 ) , .B1( u2_u10_u4_n150 ) , .A2( u2_u10_u4_n151 ) , .A1( u2_u10_u4_n152 ) , .ZN( u2_u10_u4_n167 ) );
  NOR4_X1 u2_u10_u4_U95 (.A4( u2_u10_u4_n162 ) , .A3( u2_u10_u4_n163 ) , .A2( u2_u10_u4_n164 ) , .A1( u2_u10_u4_n165 ) , .ZN( u2_u10_u4_n166 ) );
  NAND3_X1 u2_u10_u4_U96 (.ZN( u2_out10_3 ) , .A3( u2_u10_u4_n166 ) , .A1( u2_u10_u4_n167 ) , .A2( u2_u10_u4_n186 ) );
  NAND3_X1 u2_u10_u4_U97 (.A3( u2_u10_u4_n146 ) , .A2( u2_u10_u4_n147 ) , .A1( u2_u10_u4_n148 ) , .ZN( u2_u10_u4_n149 ) );
  NAND3_X1 u2_u10_u4_U98 (.A3( u2_u10_u4_n143 ) , .A2( u2_u10_u4_n144 ) , .A1( u2_u10_u4_n145 ) , .ZN( u2_u10_u4_n151 ) );
  NAND3_X1 u2_u10_u4_U99 (.A3( u2_u10_u4_n121 ) , .ZN( u2_u10_u4_n122 ) , .A2( u2_u10_u4_n144 ) , .A1( u2_u10_u4_n154 ) );
  XOR2_X1 u2_u12_U10 (.B( u2_K13_45 ) , .A( u2_R11_30 ) , .Z( u2_u12_X_45 ) );
  XOR2_X1 u2_u12_U11 (.B( u2_K13_44 ) , .A( u2_R11_29 ) , .Z( u2_u12_X_44 ) );
  XOR2_X1 u2_u12_U12 (.B( u2_K13_43 ) , .A( u2_R11_28 ) , .Z( u2_u12_X_43 ) );
  XOR2_X1 u2_u12_U13 (.B( u2_K13_42 ) , .A( u2_R11_29 ) , .Z( u2_u12_X_42 ) );
  XOR2_X1 u2_u12_U14 (.B( u2_K13_41 ) , .A( u2_R11_28 ) , .Z( u2_u12_X_41 ) );
  XOR2_X1 u2_u12_U15 (.B( u2_K13_40 ) , .A( u2_R11_27 ) , .Z( u2_u12_X_40 ) );
  XOR2_X1 u2_u12_U17 (.B( u2_K13_39 ) , .A( u2_R11_26 ) , .Z( u2_u12_X_39 ) );
  XOR2_X1 u2_u12_U18 (.B( u2_K13_38 ) , .A( u2_R11_25 ) , .Z( u2_u12_X_38 ) );
  XOR2_X1 u2_u12_U19 (.B( u2_K13_37 ) , .A( u2_R11_24 ) , .Z( u2_u12_X_37 ) );
  XOR2_X1 u2_u12_U7 (.B( u2_K13_48 ) , .A( u2_R11_1 ) , .Z( u2_u12_X_48 ) );
  XOR2_X1 u2_u12_U8 (.B( u2_K13_47 ) , .A( u2_R11_32 ) , .Z( u2_u12_X_47 ) );
  XOR2_X1 u2_u12_U9 (.B( u2_K13_46 ) , .A( u2_R11_31 ) , .Z( u2_u12_X_46 ) );
  AOI22_X1 u2_u12_u6_U10 (.A2( u2_u12_u6_n151 ) , .B2( u2_u12_u6_n161 ) , .A1( u2_u12_u6_n167 ) , .B1( u2_u12_u6_n170 ) , .ZN( u2_u12_u6_n89 ) );
  AOI21_X1 u2_u12_u6_U11 (.B1( u2_u12_u6_n107 ) , .B2( u2_u12_u6_n132 ) , .A( u2_u12_u6_n158 ) , .ZN( u2_u12_u6_n88 ) );
  AOI21_X1 u2_u12_u6_U12 (.B2( u2_u12_u6_n147 ) , .B1( u2_u12_u6_n148 ) , .ZN( u2_u12_u6_n149 ) , .A( u2_u12_u6_n158 ) );
  AOI21_X1 u2_u12_u6_U13 (.ZN( u2_u12_u6_n106 ) , .A( u2_u12_u6_n142 ) , .B2( u2_u12_u6_n159 ) , .B1( u2_u12_u6_n164 ) );
  INV_X1 u2_u12_u6_U14 (.A( u2_u12_u6_n155 ) , .ZN( u2_u12_u6_n161 ) );
  INV_X1 u2_u12_u6_U15 (.A( u2_u12_u6_n128 ) , .ZN( u2_u12_u6_n164 ) );
  NAND2_X1 u2_u12_u6_U16 (.ZN( u2_u12_u6_n110 ) , .A1( u2_u12_u6_n122 ) , .A2( u2_u12_u6_n129 ) );
  NAND2_X1 u2_u12_u6_U17 (.ZN( u2_u12_u6_n124 ) , .A2( u2_u12_u6_n146 ) , .A1( u2_u12_u6_n148 ) );
  INV_X1 u2_u12_u6_U18 (.A( u2_u12_u6_n132 ) , .ZN( u2_u12_u6_n171 ) );
  AND2_X1 u2_u12_u6_U19 (.A1( u2_u12_u6_n100 ) , .ZN( u2_u12_u6_n130 ) , .A2( u2_u12_u6_n147 ) );
  INV_X1 u2_u12_u6_U20 (.A( u2_u12_u6_n127 ) , .ZN( u2_u12_u6_n173 ) );
  INV_X1 u2_u12_u6_U21 (.A( u2_u12_u6_n121 ) , .ZN( u2_u12_u6_n167 ) );
  INV_X1 u2_u12_u6_U22 (.A( u2_u12_u6_n100 ) , .ZN( u2_u12_u6_n169 ) );
  INV_X1 u2_u12_u6_U23 (.A( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n170 ) );
  INV_X1 u2_u12_u6_U24 (.A( u2_u12_u6_n113 ) , .ZN( u2_u12_u6_n168 ) );
  AND2_X1 u2_u12_u6_U25 (.A1( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n119 ) , .ZN( u2_u12_u6_n133 ) );
  AND2_X1 u2_u12_u6_U26 (.A2( u2_u12_u6_n121 ) , .A1( u2_u12_u6_n122 ) , .ZN( u2_u12_u6_n131 ) );
  AND3_X1 u2_u12_u6_U27 (.ZN( u2_u12_u6_n120 ) , .A2( u2_u12_u6_n127 ) , .A1( u2_u12_u6_n132 ) , .A3( u2_u12_u6_n145 ) );
  INV_X1 u2_u12_u6_U28 (.A( u2_u12_u6_n146 ) , .ZN( u2_u12_u6_n163 ) );
  AOI222_X1 u2_u12_u6_U29 (.ZN( u2_u12_u6_n114 ) , .A1( u2_u12_u6_n118 ) , .A2( u2_u12_u6_n126 ) , .B2( u2_u12_u6_n151 ) , .C2( u2_u12_u6_n159 ) , .C1( u2_u12_u6_n168 ) , .B1( u2_u12_u6_n169 ) );
  INV_X1 u2_u12_u6_U3 (.A( u2_u12_u6_n110 ) , .ZN( u2_u12_u6_n166 ) );
  NOR2_X1 u2_u12_u6_U30 (.A1( u2_u12_u6_n162 ) , .A2( u2_u12_u6_n165 ) , .ZN( u2_u12_u6_n98 ) );
  AOI211_X1 u2_u12_u6_U31 (.B( u2_u12_u6_n134 ) , .A( u2_u12_u6_n135 ) , .C1( u2_u12_u6_n136 ) , .ZN( u2_u12_u6_n137 ) , .C2( u2_u12_u6_n151 ) );
  AOI21_X1 u2_u12_u6_U32 (.B2( u2_u12_u6_n132 ) , .B1( u2_u12_u6_n133 ) , .ZN( u2_u12_u6_n134 ) , .A( u2_u12_u6_n158 ) );
  AOI21_X1 u2_u12_u6_U33 (.B1( u2_u12_u6_n131 ) , .ZN( u2_u12_u6_n135 ) , .A( u2_u12_u6_n144 ) , .B2( u2_u12_u6_n146 ) );
  NAND4_X1 u2_u12_u6_U34 (.A4( u2_u12_u6_n127 ) , .A3( u2_u12_u6_n128 ) , .A2( u2_u12_u6_n129 ) , .A1( u2_u12_u6_n130 ) , .ZN( u2_u12_u6_n136 ) );
  NAND2_X1 u2_u12_u6_U35 (.A1( u2_u12_u6_n144 ) , .ZN( u2_u12_u6_n151 ) , .A2( u2_u12_u6_n158 ) );
  NAND2_X1 u2_u12_u6_U36 (.ZN( u2_u12_u6_n132 ) , .A1( u2_u12_u6_n91 ) , .A2( u2_u12_u6_n97 ) );
  AOI22_X1 u2_u12_u6_U37 (.B2( u2_u12_u6_n110 ) , .B1( u2_u12_u6_n111 ) , .A1( u2_u12_u6_n112 ) , .ZN( u2_u12_u6_n115 ) , .A2( u2_u12_u6_n161 ) );
  NAND4_X1 u2_u12_u6_U38 (.A3( u2_u12_u6_n109 ) , .ZN( u2_u12_u6_n112 ) , .A4( u2_u12_u6_n132 ) , .A2( u2_u12_u6_n147 ) , .A1( u2_u12_u6_n166 ) );
  NOR2_X1 u2_u12_u6_U39 (.ZN( u2_u12_u6_n109 ) , .A1( u2_u12_u6_n170 ) , .A2( u2_u12_u6_n173 ) );
  INV_X1 u2_u12_u6_U4 (.A( u2_u12_u6_n142 ) , .ZN( u2_u12_u6_n174 ) );
  NOR2_X1 u2_u12_u6_U40 (.A2( u2_u12_u6_n126 ) , .ZN( u2_u12_u6_n155 ) , .A1( u2_u12_u6_n160 ) );
  NAND2_X1 u2_u12_u6_U41 (.ZN( u2_u12_u6_n146 ) , .A2( u2_u12_u6_n94 ) , .A1( u2_u12_u6_n99 ) );
  AOI21_X1 u2_u12_u6_U42 (.A( u2_u12_u6_n144 ) , .B2( u2_u12_u6_n145 ) , .B1( u2_u12_u6_n146 ) , .ZN( u2_u12_u6_n150 ) );
  INV_X1 u2_u12_u6_U43 (.A( u2_u12_u6_n111 ) , .ZN( u2_u12_u6_n158 ) );
  NAND2_X1 u2_u12_u6_U44 (.ZN( u2_u12_u6_n127 ) , .A1( u2_u12_u6_n91 ) , .A2( u2_u12_u6_n92 ) );
  NAND2_X1 u2_u12_u6_U45 (.ZN( u2_u12_u6_n129 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n96 ) );
  INV_X1 u2_u12_u6_U46 (.A( u2_u12_u6_n144 ) , .ZN( u2_u12_u6_n159 ) );
  NAND2_X1 u2_u12_u6_U47 (.ZN( u2_u12_u6_n145 ) , .A2( u2_u12_u6_n97 ) , .A1( u2_u12_u6_n98 ) );
  NAND2_X1 u2_u12_u6_U48 (.ZN( u2_u12_u6_n148 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n94 ) );
  NAND2_X1 u2_u12_u6_U49 (.ZN( u2_u12_u6_n108 ) , .A2( u2_u12_u6_n139 ) , .A1( u2_u12_u6_n144 ) );
  NAND2_X1 u2_u12_u6_U5 (.A2( u2_u12_u6_n143 ) , .ZN( u2_u12_u6_n152 ) , .A1( u2_u12_u6_n166 ) );
  NAND2_X1 u2_u12_u6_U50 (.ZN( u2_u12_u6_n121 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n97 ) );
  NAND2_X1 u2_u12_u6_U51 (.ZN( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n95 ) );
  AND2_X1 u2_u12_u6_U52 (.ZN( u2_u12_u6_n118 ) , .A2( u2_u12_u6_n91 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U53 (.ZN( u2_u12_u6_n147 ) , .A2( u2_u12_u6_n98 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U54 (.ZN( u2_u12_u6_n128 ) , .A1( u2_u12_u6_n94 ) , .A2( u2_u12_u6_n96 ) );
  NAND2_X1 u2_u12_u6_U55 (.ZN( u2_u12_u6_n119 ) , .A2( u2_u12_u6_n95 ) , .A1( u2_u12_u6_n99 ) );
  NAND2_X1 u2_u12_u6_U56 (.ZN( u2_u12_u6_n123 ) , .A2( u2_u12_u6_n91 ) , .A1( u2_u12_u6_n96 ) );
  NAND2_X1 u2_u12_u6_U57 (.ZN( u2_u12_u6_n100 ) , .A2( u2_u12_u6_n92 ) , .A1( u2_u12_u6_n98 ) );
  NAND2_X1 u2_u12_u6_U58 (.ZN( u2_u12_u6_n122 ) , .A1( u2_u12_u6_n94 ) , .A2( u2_u12_u6_n97 ) );
  INV_X1 u2_u12_u6_U59 (.A( u2_u12_u6_n139 ) , .ZN( u2_u12_u6_n160 ) );
  AOI22_X1 u2_u12_u6_U6 (.B2( u2_u12_u6_n101 ) , .A1( u2_u12_u6_n102 ) , .ZN( u2_u12_u6_n103 ) , .B1( u2_u12_u6_n160 ) , .A2( u2_u12_u6_n161 ) );
  NAND2_X1 u2_u12_u6_U60 (.ZN( u2_u12_u6_n113 ) , .A1( u2_u12_u6_n96 ) , .A2( u2_u12_u6_n98 ) );
  NOR2_X1 u2_u12_u6_U61 (.A2( u2_u12_X_40 ) , .A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n126 ) );
  NOR2_X1 u2_u12_u6_U62 (.A2( u2_u12_X_39 ) , .A1( u2_u12_X_42 ) , .ZN( u2_u12_u6_n92 ) );
  NOR2_X1 u2_u12_u6_U63 (.A2( u2_u12_X_39 ) , .A1( u2_u12_u6_n156 ) , .ZN( u2_u12_u6_n97 ) );
  NOR2_X1 u2_u12_u6_U64 (.A2( u2_u12_X_38 ) , .A1( u2_u12_u6_n165 ) , .ZN( u2_u12_u6_n95 ) );
  NOR2_X1 u2_u12_u6_U65 (.A2( u2_u12_X_41 ) , .ZN( u2_u12_u6_n111 ) , .A1( u2_u12_u6_n157 ) );
  NOR2_X1 u2_u12_u6_U66 (.A2( u2_u12_X_37 ) , .A1( u2_u12_u6_n162 ) , .ZN( u2_u12_u6_n94 ) );
  NOR2_X1 u2_u12_u6_U67 (.A2( u2_u12_X_37 ) , .A1( u2_u12_X_38 ) , .ZN( u2_u12_u6_n91 ) );
  NAND2_X1 u2_u12_u6_U68 (.A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n144 ) , .A2( u2_u12_u6_n157 ) );
  NAND2_X1 u2_u12_u6_U69 (.A2( u2_u12_X_40 ) , .A1( u2_u12_X_41 ) , .ZN( u2_u12_u6_n139 ) );
  NOR2_X1 u2_u12_u6_U7 (.A1( u2_u12_u6_n118 ) , .ZN( u2_u12_u6_n143 ) , .A2( u2_u12_u6_n168 ) );
  AND2_X1 u2_u12_u6_U70 (.A1( u2_u12_X_39 ) , .A2( u2_u12_u6_n156 ) , .ZN( u2_u12_u6_n96 ) );
  AND2_X1 u2_u12_u6_U71 (.A1( u2_u12_X_39 ) , .A2( u2_u12_X_42 ) , .ZN( u2_u12_u6_n99 ) );
  INV_X1 u2_u12_u6_U72 (.A( u2_u12_X_40 ) , .ZN( u2_u12_u6_n157 ) );
  INV_X1 u2_u12_u6_U73 (.A( u2_u12_X_37 ) , .ZN( u2_u12_u6_n165 ) );
  INV_X1 u2_u12_u6_U74 (.A( u2_u12_X_38 ) , .ZN( u2_u12_u6_n162 ) );
  INV_X1 u2_u12_u6_U75 (.A( u2_u12_X_42 ) , .ZN( u2_u12_u6_n156 ) );
  NAND4_X1 u2_u12_u6_U76 (.ZN( u2_out12_32 ) , .A4( u2_u12_u6_n103 ) , .A3( u2_u12_u6_n104 ) , .A2( u2_u12_u6_n105 ) , .A1( u2_u12_u6_n106 ) );
  AOI22_X1 u2_u12_u6_U77 (.ZN( u2_u12_u6_n105 ) , .A2( u2_u12_u6_n108 ) , .A1( u2_u12_u6_n118 ) , .B2( u2_u12_u6_n126 ) , .B1( u2_u12_u6_n171 ) );
  AOI22_X1 u2_u12_u6_U78 (.ZN( u2_u12_u6_n104 ) , .A1( u2_u12_u6_n111 ) , .B1( u2_u12_u6_n124 ) , .B2( u2_u12_u6_n151 ) , .A2( u2_u12_u6_n93 ) );
  NAND4_X1 u2_u12_u6_U79 (.ZN( u2_out12_12 ) , .A4( u2_u12_u6_n114 ) , .A3( u2_u12_u6_n115 ) , .A2( u2_u12_u6_n116 ) , .A1( u2_u12_u6_n117 ) );
  INV_X1 u2_u12_u6_U8 (.ZN( u2_u12_u6_n172 ) , .A( u2_u12_u6_n88 ) );
  OAI22_X1 u2_u12_u6_U80 (.B2( u2_u12_u6_n111 ) , .ZN( u2_u12_u6_n116 ) , .B1( u2_u12_u6_n126 ) , .A2( u2_u12_u6_n164 ) , .A1( u2_u12_u6_n167 ) );
  OAI21_X1 u2_u12_u6_U81 (.A( u2_u12_u6_n108 ) , .ZN( u2_u12_u6_n117 ) , .B2( u2_u12_u6_n141 ) , .B1( u2_u12_u6_n163 ) );
  OAI211_X1 u2_u12_u6_U82 (.ZN( u2_out12_22 ) , .B( u2_u12_u6_n137 ) , .A( u2_u12_u6_n138 ) , .C2( u2_u12_u6_n139 ) , .C1( u2_u12_u6_n140 ) );
  AOI22_X1 u2_u12_u6_U83 (.B1( u2_u12_u6_n124 ) , .A2( u2_u12_u6_n125 ) , .A1( u2_u12_u6_n126 ) , .ZN( u2_u12_u6_n138 ) , .B2( u2_u12_u6_n161 ) );
  AND4_X1 u2_u12_u6_U84 (.A3( u2_u12_u6_n119 ) , .A1( u2_u12_u6_n120 ) , .A4( u2_u12_u6_n129 ) , .ZN( u2_u12_u6_n140 ) , .A2( u2_u12_u6_n143 ) );
  OAI211_X1 u2_u12_u6_U85 (.ZN( u2_out12_7 ) , .B( u2_u12_u6_n153 ) , .C2( u2_u12_u6_n154 ) , .C1( u2_u12_u6_n155 ) , .A( u2_u12_u6_n174 ) );
  NOR3_X1 u2_u12_u6_U86 (.A1( u2_u12_u6_n141 ) , .ZN( u2_u12_u6_n154 ) , .A3( u2_u12_u6_n164 ) , .A2( u2_u12_u6_n171 ) );
  AOI211_X1 u2_u12_u6_U87 (.B( u2_u12_u6_n149 ) , .A( u2_u12_u6_n150 ) , .C2( u2_u12_u6_n151 ) , .C1( u2_u12_u6_n152 ) , .ZN( u2_u12_u6_n153 ) );
  NAND3_X1 u2_u12_u6_U88 (.A2( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n125 ) , .A1( u2_u12_u6_n130 ) , .A3( u2_u12_u6_n131 ) );
  NAND3_X1 u2_u12_u6_U89 (.A3( u2_u12_u6_n133 ) , .ZN( u2_u12_u6_n141 ) , .A1( u2_u12_u6_n145 ) , .A2( u2_u12_u6_n148 ) );
  OAI21_X1 u2_u12_u6_U9 (.A( u2_u12_u6_n159 ) , .B1( u2_u12_u6_n169 ) , .B2( u2_u12_u6_n173 ) , .ZN( u2_u12_u6_n90 ) );
  NAND3_X1 u2_u12_u6_U90 (.ZN( u2_u12_u6_n101 ) , .A3( u2_u12_u6_n107 ) , .A2( u2_u12_u6_n121 ) , .A1( u2_u12_u6_n127 ) );
  NAND3_X1 u2_u12_u6_U91 (.ZN( u2_u12_u6_n102 ) , .A3( u2_u12_u6_n130 ) , .A2( u2_u12_u6_n145 ) , .A1( u2_u12_u6_n166 ) );
  NAND3_X1 u2_u12_u6_U92 (.A3( u2_u12_u6_n113 ) , .A1( u2_u12_u6_n119 ) , .A2( u2_u12_u6_n123 ) , .ZN( u2_u12_u6_n93 ) );
  NAND3_X1 u2_u12_u6_U93 (.ZN( u2_u12_u6_n142 ) , .A2( u2_u12_u6_n172 ) , .A3( u2_u12_u6_n89 ) , .A1( u2_u12_u6_n90 ) );
  AND3_X1 u2_u12_u7_U10 (.A3( u2_u12_u7_n110 ) , .A2( u2_u12_u7_n127 ) , .A1( u2_u12_u7_n132 ) , .ZN( u2_u12_u7_n92 ) );
  OAI21_X1 u2_u12_u7_U11 (.A( u2_u12_u7_n161 ) , .B1( u2_u12_u7_n168 ) , .B2( u2_u12_u7_n173 ) , .ZN( u2_u12_u7_n91 ) );
  AOI211_X1 u2_u12_u7_U12 (.A( u2_u12_u7_n117 ) , .ZN( u2_u12_u7_n118 ) , .C2( u2_u12_u7_n126 ) , .C1( u2_u12_u7_n177 ) , .B( u2_u12_u7_n180 ) );
  OAI22_X1 u2_u12_u7_U13 (.B1( u2_u12_u7_n115 ) , .ZN( u2_u12_u7_n117 ) , .A2( u2_u12_u7_n133 ) , .A1( u2_u12_u7_n137 ) , .B2( u2_u12_u7_n162 ) );
  INV_X1 u2_u12_u7_U14 (.A( u2_u12_u7_n116 ) , .ZN( u2_u12_u7_n180 ) );
  NOR3_X1 u2_u12_u7_U15 (.ZN( u2_u12_u7_n115 ) , .A3( u2_u12_u7_n145 ) , .A2( u2_u12_u7_n168 ) , .A1( u2_u12_u7_n169 ) );
  OAI211_X1 u2_u12_u7_U16 (.B( u2_u12_u7_n122 ) , .A( u2_u12_u7_n123 ) , .C2( u2_u12_u7_n124 ) , .ZN( u2_u12_u7_n154 ) , .C1( u2_u12_u7_n162 ) );
  AOI222_X1 u2_u12_u7_U17 (.ZN( u2_u12_u7_n122 ) , .C2( u2_u12_u7_n126 ) , .C1( u2_u12_u7_n145 ) , .B1( u2_u12_u7_n161 ) , .A2( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n170 ) , .A1( u2_u12_u7_n176 ) );
  INV_X1 u2_u12_u7_U18 (.A( u2_u12_u7_n133 ) , .ZN( u2_u12_u7_n176 ) );
  NOR3_X1 u2_u12_u7_U19 (.A2( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n135 ) , .ZN( u2_u12_u7_n136 ) , .A3( u2_u12_u7_n171 ) );
  NOR2_X1 u2_u12_u7_U20 (.A1( u2_u12_u7_n130 ) , .A2( u2_u12_u7_n134 ) , .ZN( u2_u12_u7_n153 ) );
  INV_X1 u2_u12_u7_U21 (.A( u2_u12_u7_n101 ) , .ZN( u2_u12_u7_n165 ) );
  NOR2_X1 u2_u12_u7_U22 (.ZN( u2_u12_u7_n111 ) , .A2( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n169 ) );
  AOI21_X1 u2_u12_u7_U23 (.ZN( u2_u12_u7_n104 ) , .B2( u2_u12_u7_n112 ) , .B1( u2_u12_u7_n127 ) , .A( u2_u12_u7_n164 ) );
  AOI21_X1 u2_u12_u7_U24 (.ZN( u2_u12_u7_n106 ) , .B1( u2_u12_u7_n133 ) , .B2( u2_u12_u7_n146 ) , .A( u2_u12_u7_n162 ) );
  AOI21_X1 u2_u12_u7_U25 (.A( u2_u12_u7_n101 ) , .ZN( u2_u12_u7_n107 ) , .B2( u2_u12_u7_n128 ) , .B1( u2_u12_u7_n175 ) );
  INV_X1 u2_u12_u7_U26 (.A( u2_u12_u7_n138 ) , .ZN( u2_u12_u7_n171 ) );
  INV_X1 u2_u12_u7_U27 (.A( u2_u12_u7_n131 ) , .ZN( u2_u12_u7_n177 ) );
  INV_X1 u2_u12_u7_U28 (.A( u2_u12_u7_n110 ) , .ZN( u2_u12_u7_n174 ) );
  NAND2_X1 u2_u12_u7_U29 (.A1( u2_u12_u7_n129 ) , .A2( u2_u12_u7_n132 ) , .ZN( u2_u12_u7_n149 ) );
  OAI21_X1 u2_u12_u7_U3 (.ZN( u2_u12_u7_n159 ) , .A( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n171 ) , .B1( u2_u12_u7_n174 ) );
  NAND2_X1 u2_u12_u7_U30 (.A1( u2_u12_u7_n113 ) , .A2( u2_u12_u7_n124 ) , .ZN( u2_u12_u7_n130 ) );
  INV_X1 u2_u12_u7_U31 (.A( u2_u12_u7_n112 ) , .ZN( u2_u12_u7_n173 ) );
  INV_X1 u2_u12_u7_U32 (.A( u2_u12_u7_n128 ) , .ZN( u2_u12_u7_n168 ) );
  INV_X1 u2_u12_u7_U33 (.A( u2_u12_u7_n148 ) , .ZN( u2_u12_u7_n169 ) );
  INV_X1 u2_u12_u7_U34 (.A( u2_u12_u7_n127 ) , .ZN( u2_u12_u7_n179 ) );
  NOR2_X1 u2_u12_u7_U35 (.ZN( u2_u12_u7_n101 ) , .A2( u2_u12_u7_n150 ) , .A1( u2_u12_u7_n156 ) );
  AOI211_X1 u2_u12_u7_U36 (.B( u2_u12_u7_n154 ) , .A( u2_u12_u7_n155 ) , .C1( u2_u12_u7_n156 ) , .ZN( u2_u12_u7_n157 ) , .C2( u2_u12_u7_n172 ) );
  INV_X1 u2_u12_u7_U37 (.A( u2_u12_u7_n153 ) , .ZN( u2_u12_u7_n172 ) );
  AOI211_X1 u2_u12_u7_U38 (.B( u2_u12_u7_n139 ) , .A( u2_u12_u7_n140 ) , .C2( u2_u12_u7_n141 ) , .ZN( u2_u12_u7_n142 ) , .C1( u2_u12_u7_n156 ) );
  NAND4_X1 u2_u12_u7_U39 (.A3( u2_u12_u7_n127 ) , .A2( u2_u12_u7_n128 ) , .A1( u2_u12_u7_n129 ) , .ZN( u2_u12_u7_n141 ) , .A4( u2_u12_u7_n147 ) );
  INV_X1 u2_u12_u7_U4 (.A( u2_u12_u7_n111 ) , .ZN( u2_u12_u7_n170 ) );
  AOI21_X1 u2_u12_u7_U40 (.A( u2_u12_u7_n137 ) , .B1( u2_u12_u7_n138 ) , .ZN( u2_u12_u7_n139 ) , .B2( u2_u12_u7_n146 ) );
  OAI22_X1 u2_u12_u7_U41 (.B1( u2_u12_u7_n136 ) , .ZN( u2_u12_u7_n140 ) , .A1( u2_u12_u7_n153 ) , .B2( u2_u12_u7_n162 ) , .A2( u2_u12_u7_n164 ) );
  AOI21_X1 u2_u12_u7_U42 (.ZN( u2_u12_u7_n123 ) , .B1( u2_u12_u7_n165 ) , .B2( u2_u12_u7_n177 ) , .A( u2_u12_u7_n97 ) );
  AOI21_X1 u2_u12_u7_U43 (.B2( u2_u12_u7_n113 ) , .B1( u2_u12_u7_n124 ) , .A( u2_u12_u7_n125 ) , .ZN( u2_u12_u7_n97 ) );
  INV_X1 u2_u12_u7_U44 (.A( u2_u12_u7_n125 ) , .ZN( u2_u12_u7_n161 ) );
  INV_X1 u2_u12_u7_U45 (.A( u2_u12_u7_n152 ) , .ZN( u2_u12_u7_n162 ) );
  AOI22_X1 u2_u12_u7_U46 (.A2( u2_u12_u7_n114 ) , .ZN( u2_u12_u7_n119 ) , .B1( u2_u12_u7_n130 ) , .A1( u2_u12_u7_n156 ) , .B2( u2_u12_u7_n165 ) );
  NAND2_X1 u2_u12_u7_U47 (.A2( u2_u12_u7_n112 ) , .ZN( u2_u12_u7_n114 ) , .A1( u2_u12_u7_n175 ) );
  AND2_X1 u2_u12_u7_U48 (.ZN( u2_u12_u7_n145 ) , .A2( u2_u12_u7_n98 ) , .A1( u2_u12_u7_n99 ) );
  NOR2_X1 u2_u12_u7_U49 (.ZN( u2_u12_u7_n137 ) , .A1( u2_u12_u7_n150 ) , .A2( u2_u12_u7_n161 ) );
  INV_X1 u2_u12_u7_U5 (.A( u2_u12_u7_n149 ) , .ZN( u2_u12_u7_n175 ) );
  AOI21_X1 u2_u12_u7_U50 (.ZN( u2_u12_u7_n105 ) , .B2( u2_u12_u7_n110 ) , .A( u2_u12_u7_n125 ) , .B1( u2_u12_u7_n147 ) );
  NAND2_X1 u2_u12_u7_U51 (.ZN( u2_u12_u7_n146 ) , .A1( u2_u12_u7_n95 ) , .A2( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U52 (.A2( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n147 ) , .A1( u2_u12_u7_n93 ) );
  NAND2_X1 u2_u12_u7_U53 (.A1( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n127 ) , .A2( u2_u12_u7_n99 ) );
  OR2_X1 u2_u12_u7_U54 (.ZN( u2_u12_u7_n126 ) , .A2( u2_u12_u7_n152 ) , .A1( u2_u12_u7_n156 ) );
  NAND2_X1 u2_u12_u7_U55 (.A2( u2_u12_u7_n102 ) , .A1( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n133 ) );
  NAND2_X1 u2_u12_u7_U56 (.ZN( u2_u12_u7_n112 ) , .A2( u2_u12_u7_n96 ) , .A1( u2_u12_u7_n99 ) );
  NAND2_X1 u2_u12_u7_U57 (.A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n128 ) , .A1( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U58 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n113 ) , .A2( u2_u12_u7_n93 ) );
  NAND2_X1 u2_u12_u7_U59 (.A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n124 ) , .A1( u2_u12_u7_n96 ) );
  INV_X1 u2_u12_u7_U6 (.A( u2_u12_u7_n154 ) , .ZN( u2_u12_u7_n178 ) );
  NAND2_X1 u2_u12_u7_U60 (.ZN( u2_u12_u7_n110 ) , .A1( u2_u12_u7_n95 ) , .A2( u2_u12_u7_n96 ) );
  INV_X1 u2_u12_u7_U61 (.A( u2_u12_u7_n150 ) , .ZN( u2_u12_u7_n164 ) );
  AND2_X1 u2_u12_u7_U62 (.ZN( u2_u12_u7_n134 ) , .A1( u2_u12_u7_n93 ) , .A2( u2_u12_u7_n98 ) );
  NAND2_X1 u2_u12_u7_U63 (.A1( u2_u12_u7_n100 ) , .A2( u2_u12_u7_n102 ) , .ZN( u2_u12_u7_n129 ) );
  NAND2_X1 u2_u12_u7_U64 (.A2( u2_u12_u7_n103 ) , .ZN( u2_u12_u7_n131 ) , .A1( u2_u12_u7_n95 ) );
  NAND2_X1 u2_u12_u7_U65 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n138 ) , .A2( u2_u12_u7_n99 ) );
  NAND2_X1 u2_u12_u7_U66 (.ZN( u2_u12_u7_n132 ) , .A1( u2_u12_u7_n93 ) , .A2( u2_u12_u7_n96 ) );
  NAND2_X1 u2_u12_u7_U67 (.A1( u2_u12_u7_n100 ) , .ZN( u2_u12_u7_n148 ) , .A2( u2_u12_u7_n95 ) );
  NOR2_X1 u2_u12_u7_U68 (.A2( u2_u12_X_47 ) , .ZN( u2_u12_u7_n150 ) , .A1( u2_u12_u7_n163 ) );
  NOR2_X1 u2_u12_u7_U69 (.A2( u2_u12_X_43 ) , .A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n103 ) );
  AOI211_X1 u2_u12_u7_U7 (.ZN( u2_u12_u7_n116 ) , .A( u2_u12_u7_n155 ) , .C1( u2_u12_u7_n161 ) , .C2( u2_u12_u7_n171 ) , .B( u2_u12_u7_n94 ) );
  NOR2_X1 u2_u12_u7_U70 (.A2( u2_u12_X_48 ) , .A1( u2_u12_u7_n166 ) , .ZN( u2_u12_u7_n95 ) );
  NOR2_X1 u2_u12_u7_U71 (.A2( u2_u12_X_45 ) , .A1( u2_u12_X_48 ) , .ZN( u2_u12_u7_n99 ) );
  NOR2_X1 u2_u12_u7_U72 (.A2( u2_u12_X_44 ) , .A1( u2_u12_u7_n167 ) , .ZN( u2_u12_u7_n98 ) );
  NOR2_X1 u2_u12_u7_U73 (.A2( u2_u12_X_46 ) , .A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n152 ) );
  AND2_X1 u2_u12_u7_U74 (.A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n156 ) , .A2( u2_u12_u7_n163 ) );
  NAND2_X1 u2_u12_u7_U75 (.A2( u2_u12_X_46 ) , .A1( u2_u12_X_47 ) , .ZN( u2_u12_u7_n125 ) );
  AND2_X1 u2_u12_u7_U76 (.A2( u2_u12_X_45 ) , .A1( u2_u12_X_48 ) , .ZN( u2_u12_u7_n102 ) );
  AND2_X1 u2_u12_u7_U77 (.A2( u2_u12_X_43 ) , .A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n96 ) );
  AND2_X1 u2_u12_u7_U78 (.A1( u2_u12_X_44 ) , .ZN( u2_u12_u7_n100 ) , .A2( u2_u12_u7_n167 ) );
  AND2_X1 u2_u12_u7_U79 (.A1( u2_u12_X_48 ) , .A2( u2_u12_u7_n166 ) , .ZN( u2_u12_u7_n93 ) );
  OAI222_X1 u2_u12_u7_U8 (.C2( u2_u12_u7_n101 ) , .B2( u2_u12_u7_n111 ) , .A1( u2_u12_u7_n113 ) , .C1( u2_u12_u7_n146 ) , .A2( u2_u12_u7_n162 ) , .B1( u2_u12_u7_n164 ) , .ZN( u2_u12_u7_n94 ) );
  INV_X1 u2_u12_u7_U80 (.A( u2_u12_X_46 ) , .ZN( u2_u12_u7_n163 ) );
  INV_X1 u2_u12_u7_U81 (.A( u2_u12_X_43 ) , .ZN( u2_u12_u7_n167 ) );
  INV_X1 u2_u12_u7_U82 (.A( u2_u12_X_45 ) , .ZN( u2_u12_u7_n166 ) );
  NAND4_X1 u2_u12_u7_U83 (.ZN( u2_out12_27 ) , .A4( u2_u12_u7_n118 ) , .A3( u2_u12_u7_n119 ) , .A2( u2_u12_u7_n120 ) , .A1( u2_u12_u7_n121 ) );
  OAI21_X1 u2_u12_u7_U84 (.ZN( u2_u12_u7_n121 ) , .B2( u2_u12_u7_n145 ) , .A( u2_u12_u7_n150 ) , .B1( u2_u12_u7_n174 ) );
  OAI21_X1 u2_u12_u7_U85 (.ZN( u2_u12_u7_n120 ) , .A( u2_u12_u7_n161 ) , .B2( u2_u12_u7_n170 ) , .B1( u2_u12_u7_n179 ) );
  NAND4_X1 u2_u12_u7_U86 (.ZN( u2_out12_21 ) , .A4( u2_u12_u7_n157 ) , .A3( u2_u12_u7_n158 ) , .A2( u2_u12_u7_n159 ) , .A1( u2_u12_u7_n160 ) );
  OAI21_X1 u2_u12_u7_U87 (.B1( u2_u12_u7_n145 ) , .ZN( u2_u12_u7_n160 ) , .A( u2_u12_u7_n161 ) , .B2( u2_u12_u7_n177 ) );
  AOI22_X1 u2_u12_u7_U88 (.B2( u2_u12_u7_n149 ) , .B1( u2_u12_u7_n150 ) , .A2( u2_u12_u7_n151 ) , .A1( u2_u12_u7_n152 ) , .ZN( u2_u12_u7_n158 ) );
  NAND4_X1 u2_u12_u7_U89 (.ZN( u2_out12_15 ) , .A4( u2_u12_u7_n142 ) , .A3( u2_u12_u7_n143 ) , .A2( u2_u12_u7_n144 ) , .A1( u2_u12_u7_n178 ) );
  OAI221_X1 u2_u12_u7_U9 (.C1( u2_u12_u7_n101 ) , .C2( u2_u12_u7_n147 ) , .ZN( u2_u12_u7_n155 ) , .B2( u2_u12_u7_n162 ) , .A( u2_u12_u7_n91 ) , .B1( u2_u12_u7_n92 ) );
  OR2_X1 u2_u12_u7_U90 (.A2( u2_u12_u7_n125 ) , .A1( u2_u12_u7_n129 ) , .ZN( u2_u12_u7_n144 ) );
  AOI22_X1 u2_u12_u7_U91 (.A2( u2_u12_u7_n126 ) , .ZN( u2_u12_u7_n143 ) , .B2( u2_u12_u7_n165 ) , .B1( u2_u12_u7_n173 ) , .A1( u2_u12_u7_n174 ) );
  NAND4_X1 u2_u12_u7_U92 (.ZN( u2_out12_5 ) , .A4( u2_u12_u7_n108 ) , .A3( u2_u12_u7_n109 ) , .A1( u2_u12_u7_n116 ) , .A2( u2_u12_u7_n123 ) );
  AOI22_X1 u2_u12_u7_U93 (.ZN( u2_u12_u7_n109 ) , .A2( u2_u12_u7_n126 ) , .B2( u2_u12_u7_n145 ) , .B1( u2_u12_u7_n156 ) , .A1( u2_u12_u7_n171 ) );
  NOR4_X1 u2_u12_u7_U94 (.A4( u2_u12_u7_n104 ) , .A3( u2_u12_u7_n105 ) , .A2( u2_u12_u7_n106 ) , .A1( u2_u12_u7_n107 ) , .ZN( u2_u12_u7_n108 ) );
  NAND3_X1 u2_u12_u7_U95 (.A3( u2_u12_u7_n146 ) , .A2( u2_u12_u7_n147 ) , .A1( u2_u12_u7_n148 ) , .ZN( u2_u12_u7_n151 ) );
  NAND3_X1 u2_u12_u7_U96 (.A3( u2_u12_u7_n131 ) , .A2( u2_u12_u7_n132 ) , .A1( u2_u12_u7_n133 ) , .ZN( u2_u12_u7_n135 ) );
  XOR2_X1 u2_u13_U1 (.B( u2_K14_9 ) , .A( u2_R12_6 ) , .Z( u2_u13_X_9 ) );
  XOR2_X1 u2_u13_U10 (.B( u2_K14_45 ) , .A( u2_R12_30 ) , .Z( u2_u13_X_45 ) );
  XOR2_X1 u2_u13_U11 (.B( u2_K14_44 ) , .A( u2_R12_29 ) , .Z( u2_u13_X_44 ) );
  XOR2_X1 u2_u13_U12 (.B( u2_K14_43 ) , .A( u2_R12_28 ) , .Z( u2_u13_X_43 ) );
  XOR2_X1 u2_u13_U13 (.B( u2_K14_42 ) , .A( u2_R12_29 ) , .Z( u2_u13_X_42 ) );
  XOR2_X1 u2_u13_U14 (.B( u2_K14_41 ) , .A( u2_R12_28 ) , .Z( u2_u13_X_41 ) );
  XOR2_X1 u2_u13_U15 (.B( u2_K14_40 ) , .A( u2_R12_27 ) , .Z( u2_u13_X_40 ) );
  XOR2_X1 u2_u13_U16 (.B( u2_K14_3 ) , .A( u2_R12_2 ) , .Z( u2_u13_X_3 ) );
  XOR2_X1 u2_u13_U17 (.B( u2_K14_39 ) , .A( u2_R12_26 ) , .Z( u2_u13_X_39 ) );
  XOR2_X1 u2_u13_U18 (.B( u2_K14_38 ) , .A( u2_R12_25 ) , .Z( u2_u13_X_38 ) );
  XOR2_X1 u2_u13_U19 (.B( u2_K14_37 ) , .A( u2_R12_24 ) , .Z( u2_u13_X_37 ) );
  XOR2_X1 u2_u13_U2 (.B( u2_K14_8 ) , .A( u2_R12_5 ) , .Z( u2_u13_X_8 ) );
  XOR2_X1 u2_u13_U27 (.B( u2_K14_2 ) , .A( u2_R12_1 ) , .Z( u2_u13_X_2 ) );
  XOR2_X1 u2_u13_U3 (.B( u2_K14_7 ) , .A( u2_R12_4 ) , .Z( u2_u13_X_7 ) );
  XOR2_X1 u2_u13_U33 (.B( u2_K14_24 ) , .A( u2_R12_17 ) , .Z( u2_u13_X_24 ) );
  XOR2_X1 u2_u13_U34 (.B( u2_K14_23 ) , .A( u2_R12_16 ) , .Z( u2_u13_X_23 ) );
  XOR2_X1 u2_u13_U35 (.B( u2_K14_22 ) , .A( u2_R12_15 ) , .Z( u2_u13_X_22 ) );
  XOR2_X1 u2_u13_U36 (.B( u2_K14_21 ) , .A( u2_R12_14 ) , .Z( u2_u13_X_21 ) );
  XOR2_X1 u2_u13_U37 (.B( u2_K14_20 ) , .A( u2_R12_13 ) , .Z( u2_u13_X_20 ) );
  XOR2_X1 u2_u13_U38 (.B( u2_K14_1 ) , .A( u2_R12_32 ) , .Z( u2_u13_X_1 ) );
  XOR2_X1 u2_u13_U39 (.B( u2_K14_19 ) , .A( u2_R12_12 ) , .Z( u2_u13_X_19 ) );
  XOR2_X1 u2_u13_U4 (.B( u2_K14_6 ) , .A( u2_R12_5 ) , .Z( u2_u13_X_6 ) );
  XOR2_X1 u2_u13_U40 (.B( u2_K14_18 ) , .A( u2_R12_13 ) , .Z( u2_u13_X_18 ) );
  XOR2_X1 u2_u13_U41 (.B( u2_K14_17 ) , .A( u2_R12_12 ) , .Z( u2_u13_X_17 ) );
  XOR2_X1 u2_u13_U42 (.B( u2_K14_16 ) , .A( u2_R12_11 ) , .Z( u2_u13_X_16 ) );
  XOR2_X1 u2_u13_U43 (.B( u2_K14_15 ) , .A( u2_R12_10 ) , .Z( u2_u13_X_15 ) );
  XOR2_X1 u2_u13_U44 (.B( u2_K14_14 ) , .A( u2_R12_9 ) , .Z( u2_u13_X_14 ) );
  XOR2_X1 u2_u13_U45 (.B( u2_K14_13 ) , .A( u2_R12_8 ) , .Z( u2_u13_X_13 ) );
  XOR2_X1 u2_u13_U46 (.B( u2_K14_12 ) , .A( u2_R12_9 ) , .Z( u2_u13_X_12 ) );
  XOR2_X1 u2_u13_U47 (.B( u2_K14_11 ) , .A( u2_R12_8 ) , .Z( u2_u13_X_11 ) );
  XOR2_X1 u2_u13_U48 (.B( u2_K14_10 ) , .A( u2_R12_7 ) , .Z( u2_u13_X_10 ) );
  XOR2_X1 u2_u13_U5 (.B( u2_K14_5 ) , .A( u2_R12_4 ) , .Z( u2_u13_X_5 ) );
  XOR2_X1 u2_u13_U6 (.B( u2_K14_4 ) , .A( u2_R12_3 ) , .Z( u2_u13_X_4 ) );
  XOR2_X1 u2_u13_U7 (.B( u2_K14_48 ) , .A( u2_R12_1 ) , .Z( u2_u13_X_48 ) );
  XOR2_X1 u2_u13_U8 (.B( u2_K14_47 ) , .A( u2_R12_32 ) , .Z( u2_u13_X_47 ) );
  XOR2_X1 u2_u13_U9 (.B( u2_K14_46 ) , .A( u2_R12_31 ) , .Z( u2_u13_X_46 ) );
  AND3_X1 u2_u13_u0_U10 (.A2( u2_u13_u0_n112 ) , .ZN( u2_u13_u0_n127 ) , .A3( u2_u13_u0_n130 ) , .A1( u2_u13_u0_n148 ) );
  NAND2_X1 u2_u13_u0_U11 (.ZN( u2_u13_u0_n113 ) , .A1( u2_u13_u0_n139 ) , .A2( u2_u13_u0_n149 ) );
  AND2_X1 u2_u13_u0_U12 (.ZN( u2_u13_u0_n107 ) , .A1( u2_u13_u0_n130 ) , .A2( u2_u13_u0_n140 ) );
  AND2_X1 u2_u13_u0_U13 (.A2( u2_u13_u0_n129 ) , .A1( u2_u13_u0_n130 ) , .ZN( u2_u13_u0_n151 ) );
  AND2_X1 u2_u13_u0_U14 (.A1( u2_u13_u0_n108 ) , .A2( u2_u13_u0_n125 ) , .ZN( u2_u13_u0_n145 ) );
  INV_X1 u2_u13_u0_U15 (.A( u2_u13_u0_n143 ) , .ZN( u2_u13_u0_n173 ) );
  NOR2_X1 u2_u13_u0_U16 (.A2( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n147 ) , .A1( u2_u13_u0_n160 ) );
  INV_X1 u2_u13_u0_U17 (.ZN( u2_u13_u0_n172 ) , .A( u2_u13_u0_n88 ) );
  OAI222_X1 u2_u13_u0_U18 (.C1( u2_u13_u0_n108 ) , .A1( u2_u13_u0_n125 ) , .B2( u2_u13_u0_n128 ) , .B1( u2_u13_u0_n144 ) , .A2( u2_u13_u0_n158 ) , .C2( u2_u13_u0_n161 ) , .ZN( u2_u13_u0_n88 ) );
  NOR2_X1 u2_u13_u0_U19 (.A1( u2_u13_u0_n163 ) , .A2( u2_u13_u0_n164 ) , .ZN( u2_u13_u0_n95 ) );
  AOI21_X1 u2_u13_u0_U20 (.B1( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n132 ) , .A( u2_u13_u0_n165 ) , .B2( u2_u13_u0_n93 ) );
  INV_X1 u2_u13_u0_U21 (.A( u2_u13_u0_n142 ) , .ZN( u2_u13_u0_n165 ) );
  OAI221_X1 u2_u13_u0_U22 (.C1( u2_u13_u0_n121 ) , .ZN( u2_u13_u0_n122 ) , .B2( u2_u13_u0_n127 ) , .A( u2_u13_u0_n143 ) , .B1( u2_u13_u0_n144 ) , .C2( u2_u13_u0_n147 ) );
  OAI22_X1 u2_u13_u0_U23 (.B1( u2_u13_u0_n125 ) , .ZN( u2_u13_u0_n126 ) , .A1( u2_u13_u0_n138 ) , .A2( u2_u13_u0_n146 ) , .B2( u2_u13_u0_n147 ) );
  OAI22_X1 u2_u13_u0_U24 (.B1( u2_u13_u0_n131 ) , .A1( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n147 ) , .A2( u2_u13_u0_n90 ) , .ZN( u2_u13_u0_n91 ) );
  AND3_X1 u2_u13_u0_U25 (.A3( u2_u13_u0_n121 ) , .A2( u2_u13_u0_n125 ) , .A1( u2_u13_u0_n148 ) , .ZN( u2_u13_u0_n90 ) );
  INV_X1 u2_u13_u0_U26 (.A( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n161 ) );
  NOR2_X1 u2_u13_u0_U27 (.A1( u2_u13_u0_n120 ) , .ZN( u2_u13_u0_n143 ) , .A2( u2_u13_u0_n167 ) );
  OAI221_X1 u2_u13_u0_U28 (.C1( u2_u13_u0_n112 ) , .ZN( u2_u13_u0_n120 ) , .B1( u2_u13_u0_n138 ) , .B2( u2_u13_u0_n141 ) , .C2( u2_u13_u0_n147 ) , .A( u2_u13_u0_n172 ) );
  AOI211_X1 u2_u13_u0_U29 (.B( u2_u13_u0_n115 ) , .A( u2_u13_u0_n116 ) , .C2( u2_u13_u0_n117 ) , .C1( u2_u13_u0_n118 ) , .ZN( u2_u13_u0_n119 ) );
  INV_X1 u2_u13_u0_U3 (.A( u2_u13_u0_n113 ) , .ZN( u2_u13_u0_n166 ) );
  AOI22_X1 u2_u13_u0_U30 (.B2( u2_u13_u0_n109 ) , .A2( u2_u13_u0_n110 ) , .ZN( u2_u13_u0_n111 ) , .B1( u2_u13_u0_n118 ) , .A1( u2_u13_u0_n160 ) );
  INV_X1 u2_u13_u0_U31 (.A( u2_u13_u0_n118 ) , .ZN( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U32 (.ZN( u2_u13_u0_n104 ) , .B1( u2_u13_u0_n107 ) , .B2( u2_u13_u0_n141 ) , .A( u2_u13_u0_n144 ) );
  AOI21_X1 u2_u13_u0_U33 (.B1( u2_u13_u0_n127 ) , .B2( u2_u13_u0_n129 ) , .A( u2_u13_u0_n138 ) , .ZN( u2_u13_u0_n96 ) );
  AOI21_X1 u2_u13_u0_U34 (.ZN( u2_u13_u0_n116 ) , .B2( u2_u13_u0_n142 ) , .A( u2_u13_u0_n144 ) , .B1( u2_u13_u0_n166 ) );
  NAND2_X1 u2_u13_u0_U35 (.A1( u2_u13_u0_n100 ) , .A2( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n125 ) );
  NAND2_X1 u2_u13_u0_U36 (.A1( u2_u13_u0_n101 ) , .A2( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n150 ) );
  INV_X1 u2_u13_u0_U37 (.A( u2_u13_u0_n138 ) , .ZN( u2_u13_u0_n160 ) );
  NAND2_X1 u2_u13_u0_U38 (.A1( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n128 ) , .A2( u2_u13_u0_n95 ) );
  NAND2_X1 u2_u13_u0_U39 (.A1( u2_u13_u0_n100 ) , .ZN( u2_u13_u0_n129 ) , .A2( u2_u13_u0_n95 ) );
  AOI21_X1 u2_u13_u0_U4 (.B1( u2_u13_u0_n114 ) , .ZN( u2_u13_u0_n115 ) , .B2( u2_u13_u0_n129 ) , .A( u2_u13_u0_n161 ) );
  NAND2_X1 u2_u13_u0_U40 (.A2( u2_u13_u0_n100 ) , .ZN( u2_u13_u0_n131 ) , .A1( u2_u13_u0_n92 ) );
  NAND2_X1 u2_u13_u0_U41 (.A2( u2_u13_u0_n100 ) , .A1( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n139 ) );
  NAND2_X1 u2_u13_u0_U42 (.ZN( u2_u13_u0_n148 ) , .A1( u2_u13_u0_n93 ) , .A2( u2_u13_u0_n95 ) );
  NAND2_X1 u2_u13_u0_U43 (.A2( u2_u13_u0_n102 ) , .A1( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n149 ) );
  NAND2_X1 u2_u13_u0_U44 (.A2( u2_u13_u0_n102 ) , .ZN( u2_u13_u0_n114 ) , .A1( u2_u13_u0_n92 ) );
  NAND2_X1 u2_u13_u0_U45 (.A2( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n121 ) , .A1( u2_u13_u0_n93 ) );
  NAND2_X1 u2_u13_u0_U46 (.ZN( u2_u13_u0_n112 ) , .A2( u2_u13_u0_n92 ) , .A1( u2_u13_u0_n93 ) );
  OR3_X1 u2_u13_u0_U47 (.A3( u2_u13_u0_n152 ) , .A2( u2_u13_u0_n153 ) , .A1( u2_u13_u0_n154 ) , .ZN( u2_u13_u0_n155 ) );
  AOI21_X1 u2_u13_u0_U48 (.B2( u2_u13_u0_n150 ) , .B1( u2_u13_u0_n151 ) , .ZN( u2_u13_u0_n152 ) , .A( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U49 (.A( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n145 ) , .B1( u2_u13_u0_n146 ) , .ZN( u2_u13_u0_n154 ) );
  AOI21_X1 u2_u13_u0_U5 (.B2( u2_u13_u0_n131 ) , .ZN( u2_u13_u0_n134 ) , .B1( u2_u13_u0_n151 ) , .A( u2_u13_u0_n158 ) );
  AOI21_X1 u2_u13_u0_U50 (.A( u2_u13_u0_n147 ) , .B2( u2_u13_u0_n148 ) , .B1( u2_u13_u0_n149 ) , .ZN( u2_u13_u0_n153 ) );
  INV_X1 u2_u13_u0_U51 (.ZN( u2_u13_u0_n171 ) , .A( u2_u13_u0_n99 ) );
  OAI211_X1 u2_u13_u0_U52 (.C2( u2_u13_u0_n140 ) , .C1( u2_u13_u0_n161 ) , .A( u2_u13_u0_n169 ) , .B( u2_u13_u0_n98 ) , .ZN( u2_u13_u0_n99 ) );
  INV_X1 u2_u13_u0_U53 (.ZN( u2_u13_u0_n169 ) , .A( u2_u13_u0_n91 ) );
  AOI211_X1 u2_u13_u0_U54 (.C1( u2_u13_u0_n118 ) , .A( u2_u13_u0_n123 ) , .B( u2_u13_u0_n96 ) , .C2( u2_u13_u0_n97 ) , .ZN( u2_u13_u0_n98 ) );
  NOR2_X1 u2_u13_u0_U55 (.A2( u2_u13_X_6 ) , .ZN( u2_u13_u0_n100 ) , .A1( u2_u13_u0_n162 ) );
  NOR2_X1 u2_u13_u0_U56 (.A2( u2_u13_X_4 ) , .A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n118 ) );
  NOR2_X1 u2_u13_u0_U57 (.A2( u2_u13_X_2 ) , .ZN( u2_u13_u0_n103 ) , .A1( u2_u13_u0_n164 ) );
  NOR2_X1 u2_u13_u0_U58 (.A2( u2_u13_X_1 ) , .A1( u2_u13_X_2 ) , .ZN( u2_u13_u0_n92 ) );
  NOR2_X1 u2_u13_u0_U59 (.A2( u2_u13_X_1 ) , .ZN( u2_u13_u0_n101 ) , .A1( u2_u13_u0_n163 ) );
  NOR2_X1 u2_u13_u0_U6 (.A1( u2_u13_u0_n108 ) , .ZN( u2_u13_u0_n123 ) , .A2( u2_u13_u0_n158 ) );
  NAND2_X1 u2_u13_u0_U60 (.A2( u2_u13_X_4 ) , .A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n144 ) );
  NOR2_X1 u2_u13_u0_U61 (.A2( u2_u13_X_5 ) , .ZN( u2_u13_u0_n136 ) , .A1( u2_u13_u0_n159 ) );
  NAND2_X1 u2_u13_u0_U62 (.A1( u2_u13_X_5 ) , .ZN( u2_u13_u0_n138 ) , .A2( u2_u13_u0_n159 ) );
  NOR2_X1 u2_u13_u0_U63 (.A2( u2_u13_X_3 ) , .A1( u2_u13_X_6 ) , .ZN( u2_u13_u0_n94 ) );
  AND2_X1 u2_u13_u0_U64 (.A2( u2_u13_X_3 ) , .A1( u2_u13_X_6 ) , .ZN( u2_u13_u0_n102 ) );
  AND2_X1 u2_u13_u0_U65 (.A1( u2_u13_X_6 ) , .A2( u2_u13_u0_n162 ) , .ZN( u2_u13_u0_n93 ) );
  INV_X1 u2_u13_u0_U66 (.A( u2_u13_X_4 ) , .ZN( u2_u13_u0_n159 ) );
  INV_X1 u2_u13_u0_U67 (.A( u2_u13_X_1 ) , .ZN( u2_u13_u0_n164 ) );
  INV_X1 u2_u13_u0_U68 (.A( u2_u13_X_2 ) , .ZN( u2_u13_u0_n163 ) );
  INV_X1 u2_u13_u0_U69 (.A( u2_u13_X_3 ) , .ZN( u2_u13_u0_n162 ) );
  OAI21_X1 u2_u13_u0_U7 (.B1( u2_u13_u0_n150 ) , .B2( u2_u13_u0_n158 ) , .A( u2_u13_u0_n172 ) , .ZN( u2_u13_u0_n89 ) );
  INV_X1 u2_u13_u0_U70 (.A( u2_u13_u0_n126 ) , .ZN( u2_u13_u0_n168 ) );
  AOI211_X1 u2_u13_u0_U71 (.B( u2_u13_u0_n133 ) , .A( u2_u13_u0_n134 ) , .C2( u2_u13_u0_n135 ) , .C1( u2_u13_u0_n136 ) , .ZN( u2_u13_u0_n137 ) );
  INV_X1 u2_u13_u0_U72 (.ZN( u2_u13_u0_n174 ) , .A( u2_u13_u0_n89 ) );
  AOI211_X1 u2_u13_u0_U73 (.B( u2_u13_u0_n104 ) , .A( u2_u13_u0_n105 ) , .ZN( u2_u13_u0_n106 ) , .C2( u2_u13_u0_n113 ) , .C1( u2_u13_u0_n160 ) );
  OR4_X1 u2_u13_u0_U74 (.ZN( u2_out13_17 ) , .A4( u2_u13_u0_n122 ) , .A2( u2_u13_u0_n123 ) , .A1( u2_u13_u0_n124 ) , .A3( u2_u13_u0_n170 ) );
  AOI21_X1 u2_u13_u0_U75 (.B2( u2_u13_u0_n107 ) , .ZN( u2_u13_u0_n124 ) , .B1( u2_u13_u0_n128 ) , .A( u2_u13_u0_n161 ) );
  INV_X1 u2_u13_u0_U76 (.A( u2_u13_u0_n111 ) , .ZN( u2_u13_u0_n170 ) );
  OR4_X1 u2_u13_u0_U77 (.ZN( u2_out13_31 ) , .A4( u2_u13_u0_n155 ) , .A2( u2_u13_u0_n156 ) , .A1( u2_u13_u0_n157 ) , .A3( u2_u13_u0_n173 ) );
  AOI21_X1 u2_u13_u0_U78 (.A( u2_u13_u0_n138 ) , .B2( u2_u13_u0_n139 ) , .B1( u2_u13_u0_n140 ) , .ZN( u2_u13_u0_n157 ) );
  AOI21_X1 u2_u13_u0_U79 (.B2( u2_u13_u0_n141 ) , .B1( u2_u13_u0_n142 ) , .ZN( u2_u13_u0_n156 ) , .A( u2_u13_u0_n161 ) );
  AND2_X1 u2_u13_u0_U8 (.A1( u2_u13_u0_n114 ) , .A2( u2_u13_u0_n121 ) , .ZN( u2_u13_u0_n146 ) );
  AOI21_X1 u2_u13_u0_U80 (.B1( u2_u13_u0_n132 ) , .ZN( u2_u13_u0_n133 ) , .A( u2_u13_u0_n144 ) , .B2( u2_u13_u0_n166 ) );
  OAI22_X1 u2_u13_u0_U81 (.ZN( u2_u13_u0_n105 ) , .A2( u2_u13_u0_n132 ) , .B1( u2_u13_u0_n146 ) , .A1( u2_u13_u0_n147 ) , .B2( u2_u13_u0_n161 ) );
  NAND2_X1 u2_u13_u0_U82 (.ZN( u2_u13_u0_n110 ) , .A2( u2_u13_u0_n132 ) , .A1( u2_u13_u0_n145 ) );
  INV_X1 u2_u13_u0_U83 (.A( u2_u13_u0_n119 ) , .ZN( u2_u13_u0_n167 ) );
  NAND2_X1 u2_u13_u0_U84 (.A2( u2_u13_u0_n103 ) , .ZN( u2_u13_u0_n140 ) , .A1( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U85 (.A1( u2_u13_u0_n101 ) , .ZN( u2_u13_u0_n130 ) , .A2( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U86 (.ZN( u2_u13_u0_n108 ) , .A1( u2_u13_u0_n92 ) , .A2( u2_u13_u0_n94 ) );
  NAND2_X1 u2_u13_u0_U87 (.ZN( u2_u13_u0_n142 ) , .A1( u2_u13_u0_n94 ) , .A2( u2_u13_u0_n95 ) );
  NAND3_X1 u2_u13_u0_U88 (.ZN( u2_out13_23 ) , .A3( u2_u13_u0_n137 ) , .A1( u2_u13_u0_n168 ) , .A2( u2_u13_u0_n171 ) );
  NAND3_X1 u2_u13_u0_U89 (.A3( u2_u13_u0_n127 ) , .A2( u2_u13_u0_n128 ) , .ZN( u2_u13_u0_n135 ) , .A1( u2_u13_u0_n150 ) );
  AND2_X1 u2_u13_u0_U9 (.A1( u2_u13_u0_n131 ) , .ZN( u2_u13_u0_n141 ) , .A2( u2_u13_u0_n150 ) );
  NAND3_X1 u2_u13_u0_U90 (.ZN( u2_u13_u0_n117 ) , .A3( u2_u13_u0_n132 ) , .A2( u2_u13_u0_n139 ) , .A1( u2_u13_u0_n148 ) );
  NAND3_X1 u2_u13_u0_U91 (.ZN( u2_u13_u0_n109 ) , .A2( u2_u13_u0_n114 ) , .A3( u2_u13_u0_n140 ) , .A1( u2_u13_u0_n149 ) );
  NAND3_X1 u2_u13_u0_U92 (.ZN( u2_out13_9 ) , .A3( u2_u13_u0_n106 ) , .A2( u2_u13_u0_n171 ) , .A1( u2_u13_u0_n174 ) );
  NAND3_X1 u2_u13_u0_U93 (.A2( u2_u13_u0_n128 ) , .A1( u2_u13_u0_n132 ) , .A3( u2_u13_u0_n146 ) , .ZN( u2_u13_u0_n97 ) );
  AOI21_X1 u2_u13_u1_U10 (.B2( u2_u13_u1_n155 ) , .B1( u2_u13_u1_n156 ) , .ZN( u2_u13_u1_n157 ) , .A( u2_u13_u1_n174 ) );
  NAND3_X1 u2_u13_u1_U100 (.ZN( u2_u13_u1_n113 ) , .A1( u2_u13_u1_n120 ) , .A3( u2_u13_u1_n133 ) , .A2( u2_u13_u1_n155 ) );
  NAND2_X1 u2_u13_u1_U11 (.ZN( u2_u13_u1_n140 ) , .A2( u2_u13_u1_n150 ) , .A1( u2_u13_u1_n155 ) );
  NAND2_X1 u2_u13_u1_U12 (.A1( u2_u13_u1_n131 ) , .ZN( u2_u13_u1_n147 ) , .A2( u2_u13_u1_n153 ) );
  INV_X1 u2_u13_u1_U13 (.A( u2_u13_u1_n139 ) , .ZN( u2_u13_u1_n174 ) );
  OR4_X1 u2_u13_u1_U14 (.A4( u2_u13_u1_n106 ) , .A3( u2_u13_u1_n107 ) , .ZN( u2_u13_u1_n108 ) , .A1( u2_u13_u1_n117 ) , .A2( u2_u13_u1_n184 ) );
  AOI21_X1 u2_u13_u1_U15 (.ZN( u2_u13_u1_n106 ) , .A( u2_u13_u1_n112 ) , .B1( u2_u13_u1_n154 ) , .B2( u2_u13_u1_n156 ) );
  AOI21_X1 u2_u13_u1_U16 (.ZN( u2_u13_u1_n107 ) , .B1( u2_u13_u1_n134 ) , .B2( u2_u13_u1_n149 ) , .A( u2_u13_u1_n174 ) );
  INV_X1 u2_u13_u1_U17 (.A( u2_u13_u1_n101 ) , .ZN( u2_u13_u1_n184 ) );
  INV_X1 u2_u13_u1_U18 (.A( u2_u13_u1_n112 ) , .ZN( u2_u13_u1_n171 ) );
  NAND2_X1 u2_u13_u1_U19 (.ZN( u2_u13_u1_n141 ) , .A1( u2_u13_u1_n153 ) , .A2( u2_u13_u1_n156 ) );
  AND2_X1 u2_u13_u1_U20 (.A1( u2_u13_u1_n123 ) , .ZN( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n161 ) );
  NAND2_X1 u2_u13_u1_U21 (.A2( u2_u13_u1_n115 ) , .A1( u2_u13_u1_n116 ) , .ZN( u2_u13_u1_n148 ) );
  NAND2_X1 u2_u13_u1_U22 (.A2( u2_u13_u1_n133 ) , .A1( u2_u13_u1_n135 ) , .ZN( u2_u13_u1_n159 ) );
  NAND2_X1 u2_u13_u1_U23 (.A2( u2_u13_u1_n115 ) , .A1( u2_u13_u1_n120 ) , .ZN( u2_u13_u1_n132 ) );
  INV_X1 u2_u13_u1_U24 (.A( u2_u13_u1_n154 ) , .ZN( u2_u13_u1_n178 ) );
  AOI22_X1 u2_u13_u1_U25 (.B2( u2_u13_u1_n113 ) , .A2( u2_u13_u1_n114 ) , .ZN( u2_u13_u1_n125 ) , .A1( u2_u13_u1_n171 ) , .B1( u2_u13_u1_n173 ) );
  NAND2_X1 u2_u13_u1_U26 (.ZN( u2_u13_u1_n114 ) , .A1( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n156 ) );
  INV_X1 u2_u13_u1_U27 (.A( u2_u13_u1_n151 ) , .ZN( u2_u13_u1_n183 ) );
  AND2_X1 u2_u13_u1_U28 (.A1( u2_u13_u1_n129 ) , .A2( u2_u13_u1_n133 ) , .ZN( u2_u13_u1_n149 ) );
  INV_X1 u2_u13_u1_U29 (.A( u2_u13_u1_n131 ) , .ZN( u2_u13_u1_n180 ) );
  INV_X1 u2_u13_u1_U3 (.A( u2_u13_u1_n159 ) , .ZN( u2_u13_u1_n182 ) );
  OAI221_X1 u2_u13_u1_U30 (.A( u2_u13_u1_n119 ) , .C2( u2_u13_u1_n129 ) , .ZN( u2_u13_u1_n138 ) , .B2( u2_u13_u1_n152 ) , .C1( u2_u13_u1_n174 ) , .B1( u2_u13_u1_n187 ) );
  INV_X1 u2_u13_u1_U31 (.A( u2_u13_u1_n148 ) , .ZN( u2_u13_u1_n187 ) );
  AOI211_X1 u2_u13_u1_U32 (.B( u2_u13_u1_n117 ) , .A( u2_u13_u1_n118 ) , .ZN( u2_u13_u1_n119 ) , .C2( u2_u13_u1_n146 ) , .C1( u2_u13_u1_n159 ) );
  NOR2_X1 u2_u13_u1_U33 (.A1( u2_u13_u1_n168 ) , .A2( u2_u13_u1_n176 ) , .ZN( u2_u13_u1_n98 ) );
  AOI211_X1 u2_u13_u1_U34 (.B( u2_u13_u1_n162 ) , .A( u2_u13_u1_n163 ) , .C2( u2_u13_u1_n164 ) , .ZN( u2_u13_u1_n165 ) , .C1( u2_u13_u1_n171 ) );
  AOI21_X1 u2_u13_u1_U35 (.A( u2_u13_u1_n160 ) , .B2( u2_u13_u1_n161 ) , .ZN( u2_u13_u1_n162 ) , .B1( u2_u13_u1_n182 ) );
  OR2_X1 u2_u13_u1_U36 (.A2( u2_u13_u1_n157 ) , .A1( u2_u13_u1_n158 ) , .ZN( u2_u13_u1_n163 ) );
  OAI21_X1 u2_u13_u1_U37 (.B2( u2_u13_u1_n123 ) , .ZN( u2_u13_u1_n145 ) , .B1( u2_u13_u1_n160 ) , .A( u2_u13_u1_n185 ) );
  INV_X1 u2_u13_u1_U38 (.A( u2_u13_u1_n122 ) , .ZN( u2_u13_u1_n185 ) );
  AOI21_X1 u2_u13_u1_U39 (.B2( u2_u13_u1_n120 ) , .B1( u2_u13_u1_n121 ) , .ZN( u2_u13_u1_n122 ) , .A( u2_u13_u1_n128 ) );
  AOI221_X1 u2_u13_u1_U4 (.A( u2_u13_u1_n138 ) , .C2( u2_u13_u1_n139 ) , .C1( u2_u13_u1_n140 ) , .B2( u2_u13_u1_n141 ) , .ZN( u2_u13_u1_n142 ) , .B1( u2_u13_u1_n175 ) );
  NAND2_X1 u2_u13_u1_U40 (.A1( u2_u13_u1_n128 ) , .ZN( u2_u13_u1_n146 ) , .A2( u2_u13_u1_n160 ) );
  NAND2_X1 u2_u13_u1_U41 (.A2( u2_u13_u1_n112 ) , .ZN( u2_u13_u1_n139 ) , .A1( u2_u13_u1_n152 ) );
  NAND2_X1 u2_u13_u1_U42 (.A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n156 ) , .A2( u2_u13_u1_n99 ) );
  AOI221_X1 u2_u13_u1_U43 (.B1( u2_u13_u1_n140 ) , .ZN( u2_u13_u1_n167 ) , .B2( u2_u13_u1_n172 ) , .C2( u2_u13_u1_n175 ) , .C1( u2_u13_u1_n178 ) , .A( u2_u13_u1_n188 ) );
  INV_X1 u2_u13_u1_U44 (.ZN( u2_u13_u1_n188 ) , .A( u2_u13_u1_n97 ) );
  AOI211_X1 u2_u13_u1_U45 (.A( u2_u13_u1_n118 ) , .C1( u2_u13_u1_n132 ) , .C2( u2_u13_u1_n139 ) , .B( u2_u13_u1_n96 ) , .ZN( u2_u13_u1_n97 ) );
  AOI21_X1 u2_u13_u1_U46 (.B2( u2_u13_u1_n121 ) , .B1( u2_u13_u1_n135 ) , .A( u2_u13_u1_n152 ) , .ZN( u2_u13_u1_n96 ) );
  NOR2_X1 u2_u13_u1_U47 (.ZN( u2_u13_u1_n117 ) , .A1( u2_u13_u1_n121 ) , .A2( u2_u13_u1_n160 ) );
  AOI21_X1 u2_u13_u1_U48 (.A( u2_u13_u1_n128 ) , .B2( u2_u13_u1_n129 ) , .ZN( u2_u13_u1_n130 ) , .B1( u2_u13_u1_n150 ) );
  NAND2_X1 u2_u13_u1_U49 (.ZN( u2_u13_u1_n112 ) , .A1( u2_u13_u1_n169 ) , .A2( u2_u13_u1_n170 ) );
  AOI211_X1 u2_u13_u1_U5 (.ZN( u2_u13_u1_n124 ) , .A( u2_u13_u1_n138 ) , .C2( u2_u13_u1_n139 ) , .B( u2_u13_u1_n145 ) , .C1( u2_u13_u1_n147 ) );
  NAND2_X1 u2_u13_u1_U50 (.ZN( u2_u13_u1_n129 ) , .A2( u2_u13_u1_n95 ) , .A1( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U51 (.A1( u2_u13_u1_n102 ) , .ZN( u2_u13_u1_n154 ) , .A2( u2_u13_u1_n99 ) );
  NAND2_X1 u2_u13_u1_U52 (.A2( u2_u13_u1_n100 ) , .ZN( u2_u13_u1_n135 ) , .A1( u2_u13_u1_n99 ) );
  AOI21_X1 u2_u13_u1_U53 (.A( u2_u13_u1_n152 ) , .B2( u2_u13_u1_n153 ) , .B1( u2_u13_u1_n154 ) , .ZN( u2_u13_u1_n158 ) );
  INV_X1 u2_u13_u1_U54 (.A( u2_u13_u1_n160 ) , .ZN( u2_u13_u1_n175 ) );
  NAND2_X1 u2_u13_u1_U55 (.A1( u2_u13_u1_n100 ) , .ZN( u2_u13_u1_n116 ) , .A2( u2_u13_u1_n95 ) );
  NAND2_X1 u2_u13_u1_U56 (.A1( u2_u13_u1_n102 ) , .ZN( u2_u13_u1_n131 ) , .A2( u2_u13_u1_n95 ) );
  NAND2_X1 u2_u13_u1_U57 (.A2( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n121 ) , .A1( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U58 (.A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n153 ) , .A2( u2_u13_u1_n98 ) );
  NAND2_X1 u2_u13_u1_U59 (.A2( u2_u13_u1_n104 ) , .A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n133 ) );
  AOI22_X1 u2_u13_u1_U6 (.B2( u2_u13_u1_n136 ) , .A2( u2_u13_u1_n137 ) , .ZN( u2_u13_u1_n143 ) , .A1( u2_u13_u1_n171 ) , .B1( u2_u13_u1_n173 ) );
  NAND2_X1 u2_u13_u1_U60 (.ZN( u2_u13_u1_n150 ) , .A2( u2_u13_u1_n98 ) , .A1( u2_u13_u1_n99 ) );
  NAND2_X1 u2_u13_u1_U61 (.A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n155 ) , .A2( u2_u13_u1_n95 ) );
  OAI21_X1 u2_u13_u1_U62 (.ZN( u2_u13_u1_n109 ) , .B1( u2_u13_u1_n129 ) , .B2( u2_u13_u1_n160 ) , .A( u2_u13_u1_n167 ) );
  NAND2_X1 u2_u13_u1_U63 (.A2( u2_u13_u1_n100 ) , .A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n120 ) );
  NAND2_X1 u2_u13_u1_U64 (.A1( u2_u13_u1_n102 ) , .A2( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n115 ) );
  NAND2_X1 u2_u13_u1_U65 (.A2( u2_u13_u1_n100 ) , .A1( u2_u13_u1_n104 ) , .ZN( u2_u13_u1_n151 ) );
  NAND2_X1 u2_u13_u1_U66 (.A2( u2_u13_u1_n103 ) , .A1( u2_u13_u1_n105 ) , .ZN( u2_u13_u1_n161 ) );
  INV_X1 u2_u13_u1_U67 (.A( u2_u13_u1_n152 ) , .ZN( u2_u13_u1_n173 ) );
  INV_X1 u2_u13_u1_U68 (.A( u2_u13_u1_n128 ) , .ZN( u2_u13_u1_n172 ) );
  NAND2_X1 u2_u13_u1_U69 (.A2( u2_u13_u1_n102 ) , .A1( u2_u13_u1_n103 ) , .ZN( u2_u13_u1_n123 ) );
  INV_X1 u2_u13_u1_U7 (.A( u2_u13_u1_n147 ) , .ZN( u2_u13_u1_n181 ) );
  NOR2_X1 u2_u13_u1_U70 (.A2( u2_u13_X_7 ) , .A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n95 ) );
  NOR2_X1 u2_u13_u1_U71 (.A1( u2_u13_X_12 ) , .A2( u2_u13_X_9 ) , .ZN( u2_u13_u1_n100 ) );
  NOR2_X1 u2_u13_u1_U72 (.A2( u2_u13_X_8 ) , .A1( u2_u13_u1_n177 ) , .ZN( u2_u13_u1_n99 ) );
  NOR2_X1 u2_u13_u1_U73 (.A2( u2_u13_X_12 ) , .ZN( u2_u13_u1_n102 ) , .A1( u2_u13_u1_n176 ) );
  NOR2_X1 u2_u13_u1_U74 (.A2( u2_u13_X_9 ) , .ZN( u2_u13_u1_n105 ) , .A1( u2_u13_u1_n168 ) );
  NAND2_X1 u2_u13_u1_U75 (.A1( u2_u13_X_10 ) , .ZN( u2_u13_u1_n160 ) , .A2( u2_u13_u1_n169 ) );
  NAND2_X1 u2_u13_u1_U76 (.A2( u2_u13_X_10 ) , .A1( u2_u13_X_11 ) , .ZN( u2_u13_u1_n152 ) );
  NAND2_X1 u2_u13_u1_U77 (.A1( u2_u13_X_11 ) , .ZN( u2_u13_u1_n128 ) , .A2( u2_u13_u1_n170 ) );
  AND2_X1 u2_u13_u1_U78 (.A2( u2_u13_X_7 ) , .A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n104 ) );
  AND2_X1 u2_u13_u1_U79 (.A1( u2_u13_X_8 ) , .ZN( u2_u13_u1_n103 ) , .A2( u2_u13_u1_n177 ) );
  NOR2_X1 u2_u13_u1_U8 (.A1( u2_u13_u1_n112 ) , .A2( u2_u13_u1_n116 ) , .ZN( u2_u13_u1_n118 ) );
  INV_X1 u2_u13_u1_U80 (.A( u2_u13_X_10 ) , .ZN( u2_u13_u1_n170 ) );
  INV_X1 u2_u13_u1_U81 (.A( u2_u13_X_9 ) , .ZN( u2_u13_u1_n176 ) );
  INV_X1 u2_u13_u1_U82 (.A( u2_u13_X_11 ) , .ZN( u2_u13_u1_n169 ) );
  INV_X1 u2_u13_u1_U83 (.A( u2_u13_X_12 ) , .ZN( u2_u13_u1_n168 ) );
  INV_X1 u2_u13_u1_U84 (.A( u2_u13_X_7 ) , .ZN( u2_u13_u1_n177 ) );
  NAND4_X1 u2_u13_u1_U85 (.ZN( u2_out13_28 ) , .A4( u2_u13_u1_n124 ) , .A3( u2_u13_u1_n125 ) , .A2( u2_u13_u1_n126 ) , .A1( u2_u13_u1_n127 ) );
  OAI21_X1 u2_u13_u1_U86 (.ZN( u2_u13_u1_n127 ) , .B2( u2_u13_u1_n139 ) , .B1( u2_u13_u1_n175 ) , .A( u2_u13_u1_n183 ) );
  OAI21_X1 u2_u13_u1_U87 (.ZN( u2_u13_u1_n126 ) , .B2( u2_u13_u1_n140 ) , .A( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n178 ) );
  NAND4_X1 u2_u13_u1_U88 (.ZN( u2_out13_18 ) , .A4( u2_u13_u1_n165 ) , .A3( u2_u13_u1_n166 ) , .A1( u2_u13_u1_n167 ) , .A2( u2_u13_u1_n186 ) );
  AOI22_X1 u2_u13_u1_U89 (.B2( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n147 ) , .A2( u2_u13_u1_n148 ) , .ZN( u2_u13_u1_n166 ) , .A1( u2_u13_u1_n172 ) );
  OAI21_X1 u2_u13_u1_U9 (.ZN( u2_u13_u1_n101 ) , .B1( u2_u13_u1_n141 ) , .A( u2_u13_u1_n146 ) , .B2( u2_u13_u1_n183 ) );
  INV_X1 u2_u13_u1_U90 (.A( u2_u13_u1_n145 ) , .ZN( u2_u13_u1_n186 ) );
  NAND4_X1 u2_u13_u1_U91 (.ZN( u2_out13_2 ) , .A4( u2_u13_u1_n142 ) , .A3( u2_u13_u1_n143 ) , .A2( u2_u13_u1_n144 ) , .A1( u2_u13_u1_n179 ) );
  OAI21_X1 u2_u13_u1_U92 (.B2( u2_u13_u1_n132 ) , .ZN( u2_u13_u1_n144 ) , .A( u2_u13_u1_n146 ) , .B1( u2_u13_u1_n180 ) );
  INV_X1 u2_u13_u1_U93 (.A( u2_u13_u1_n130 ) , .ZN( u2_u13_u1_n179 ) );
  OR4_X1 u2_u13_u1_U94 (.ZN( u2_out13_13 ) , .A4( u2_u13_u1_n108 ) , .A3( u2_u13_u1_n109 ) , .A2( u2_u13_u1_n110 ) , .A1( u2_u13_u1_n111 ) );
  AOI21_X1 u2_u13_u1_U95 (.ZN( u2_u13_u1_n111 ) , .A( u2_u13_u1_n128 ) , .B2( u2_u13_u1_n131 ) , .B1( u2_u13_u1_n135 ) );
  AOI21_X1 u2_u13_u1_U96 (.ZN( u2_u13_u1_n110 ) , .A( u2_u13_u1_n116 ) , .B1( u2_u13_u1_n152 ) , .B2( u2_u13_u1_n160 ) );
  NAND3_X1 u2_u13_u1_U97 (.A3( u2_u13_u1_n149 ) , .A2( u2_u13_u1_n150 ) , .A1( u2_u13_u1_n151 ) , .ZN( u2_u13_u1_n164 ) );
  NAND3_X1 u2_u13_u1_U98 (.A3( u2_u13_u1_n134 ) , .A2( u2_u13_u1_n135 ) , .ZN( u2_u13_u1_n136 ) , .A1( u2_u13_u1_n151 ) );
  NAND3_X1 u2_u13_u1_U99 (.A1( u2_u13_u1_n133 ) , .ZN( u2_u13_u1_n137 ) , .A2( u2_u13_u1_n154 ) , .A3( u2_u13_u1_n181 ) );
  OAI22_X1 u2_u13_u2_U10 (.B1( u2_u13_u2_n151 ) , .A2( u2_u13_u2_n152 ) , .A1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n160 ) , .B2( u2_u13_u2_n168 ) );
  NAND3_X1 u2_u13_u2_U100 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n98 ) );
  NOR3_X1 u2_u13_u2_U11 (.A1( u2_u13_u2_n150 ) , .ZN( u2_u13_u2_n151 ) , .A3( u2_u13_u2_n175 ) , .A2( u2_u13_u2_n188 ) );
  AOI21_X1 u2_u13_u2_U12 (.B2( u2_u13_u2_n123 ) , .ZN( u2_u13_u2_n125 ) , .A( u2_u13_u2_n171 ) , .B1( u2_u13_u2_n184 ) );
  INV_X1 u2_u13_u2_U13 (.A( u2_u13_u2_n150 ) , .ZN( u2_u13_u2_n184 ) );
  AOI21_X1 u2_u13_u2_U14 (.ZN( u2_u13_u2_n144 ) , .B2( u2_u13_u2_n155 ) , .A( u2_u13_u2_n172 ) , .B1( u2_u13_u2_n185 ) );
  AOI21_X1 u2_u13_u2_U15 (.B2( u2_u13_u2_n143 ) , .ZN( u2_u13_u2_n145 ) , .B1( u2_u13_u2_n152 ) , .A( u2_u13_u2_n171 ) );
  INV_X1 u2_u13_u2_U16 (.A( u2_u13_u2_n156 ) , .ZN( u2_u13_u2_n171 ) );
  INV_X1 u2_u13_u2_U17 (.A( u2_u13_u2_n120 ) , .ZN( u2_u13_u2_n188 ) );
  NAND2_X1 u2_u13_u2_U18 (.A2( u2_u13_u2_n122 ) , .ZN( u2_u13_u2_n150 ) , .A1( u2_u13_u2_n152 ) );
  INV_X1 u2_u13_u2_U19 (.A( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n170 ) );
  INV_X1 u2_u13_u2_U20 (.A( u2_u13_u2_n137 ) , .ZN( u2_u13_u2_n173 ) );
  NAND2_X1 u2_u13_u2_U21 (.A1( u2_u13_u2_n132 ) , .A2( u2_u13_u2_n139 ) , .ZN( u2_u13_u2_n157 ) );
  INV_X1 u2_u13_u2_U22 (.A( u2_u13_u2_n113 ) , .ZN( u2_u13_u2_n178 ) );
  INV_X1 u2_u13_u2_U23 (.A( u2_u13_u2_n139 ) , .ZN( u2_u13_u2_n175 ) );
  INV_X1 u2_u13_u2_U24 (.A( u2_u13_u2_n155 ) , .ZN( u2_u13_u2_n181 ) );
  INV_X1 u2_u13_u2_U25 (.A( u2_u13_u2_n119 ) , .ZN( u2_u13_u2_n177 ) );
  INV_X1 u2_u13_u2_U26 (.A( u2_u13_u2_n116 ) , .ZN( u2_u13_u2_n180 ) );
  INV_X1 u2_u13_u2_U27 (.A( u2_u13_u2_n131 ) , .ZN( u2_u13_u2_n179 ) );
  INV_X1 u2_u13_u2_U28 (.A( u2_u13_u2_n154 ) , .ZN( u2_u13_u2_n176 ) );
  NAND2_X1 u2_u13_u2_U29 (.A2( u2_u13_u2_n116 ) , .A1( u2_u13_u2_n117 ) , .ZN( u2_u13_u2_n118 ) );
  NOR2_X1 u2_u13_u2_U3 (.ZN( u2_u13_u2_n121 ) , .A2( u2_u13_u2_n177 ) , .A1( u2_u13_u2_n180 ) );
  INV_X1 u2_u13_u2_U30 (.A( u2_u13_u2_n132 ) , .ZN( u2_u13_u2_n182 ) );
  INV_X1 u2_u13_u2_U31 (.A( u2_u13_u2_n158 ) , .ZN( u2_u13_u2_n183 ) );
  OAI21_X1 u2_u13_u2_U32 (.A( u2_u13_u2_n156 ) , .B1( u2_u13_u2_n157 ) , .ZN( u2_u13_u2_n158 ) , .B2( u2_u13_u2_n179 ) );
  NOR2_X1 u2_u13_u2_U33 (.ZN( u2_u13_u2_n156 ) , .A1( u2_u13_u2_n166 ) , .A2( u2_u13_u2_n169 ) );
  NOR2_X1 u2_u13_u2_U34 (.A2( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n137 ) , .A1( u2_u13_u2_n140 ) );
  NOR2_X1 u2_u13_u2_U35 (.A2( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n153 ) , .A1( u2_u13_u2_n156 ) );
  AOI211_X1 u2_u13_u2_U36 (.ZN( u2_u13_u2_n130 ) , .C1( u2_u13_u2_n138 ) , .C2( u2_u13_u2_n179 ) , .B( u2_u13_u2_n96 ) , .A( u2_u13_u2_n97 ) );
  OAI22_X1 u2_u13_u2_U37 (.B1( u2_u13_u2_n133 ) , .A2( u2_u13_u2_n137 ) , .A1( u2_u13_u2_n152 ) , .B2( u2_u13_u2_n168 ) , .ZN( u2_u13_u2_n97 ) );
  OAI221_X1 u2_u13_u2_U38 (.B1( u2_u13_u2_n113 ) , .C1( u2_u13_u2_n132 ) , .A( u2_u13_u2_n149 ) , .B2( u2_u13_u2_n171 ) , .C2( u2_u13_u2_n172 ) , .ZN( u2_u13_u2_n96 ) );
  OAI221_X1 u2_u13_u2_U39 (.A( u2_u13_u2_n115 ) , .C2( u2_u13_u2_n123 ) , .B2( u2_u13_u2_n143 ) , .B1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n163 ) , .C1( u2_u13_u2_n168 ) );
  INV_X1 u2_u13_u2_U4 (.A( u2_u13_u2_n134 ) , .ZN( u2_u13_u2_n185 ) );
  OAI21_X1 u2_u13_u2_U40 (.A( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n115 ) , .B1( u2_u13_u2_n176 ) , .B2( u2_u13_u2_n178 ) );
  OAI221_X1 u2_u13_u2_U41 (.A( u2_u13_u2_n135 ) , .B2( u2_u13_u2_n136 ) , .B1( u2_u13_u2_n137 ) , .ZN( u2_u13_u2_n162 ) , .C2( u2_u13_u2_n167 ) , .C1( u2_u13_u2_n185 ) );
  AND3_X1 u2_u13_u2_U42 (.A3( u2_u13_u2_n131 ) , .A2( u2_u13_u2_n132 ) , .A1( u2_u13_u2_n133 ) , .ZN( u2_u13_u2_n136 ) );
  AOI22_X1 u2_u13_u2_U43 (.ZN( u2_u13_u2_n135 ) , .B1( u2_u13_u2_n140 ) , .A1( u2_u13_u2_n156 ) , .B2( u2_u13_u2_n180 ) , .A2( u2_u13_u2_n188 ) );
  AOI21_X1 u2_u13_u2_U44 (.ZN( u2_u13_u2_n149 ) , .B1( u2_u13_u2_n173 ) , .B2( u2_u13_u2_n188 ) , .A( u2_u13_u2_n95 ) );
  AND3_X1 u2_u13_u2_U45 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n156 ) , .ZN( u2_u13_u2_n95 ) );
  OAI21_X1 u2_u13_u2_U46 (.A( u2_u13_u2_n141 ) , .B2( u2_u13_u2_n142 ) , .ZN( u2_u13_u2_n146 ) , .B1( u2_u13_u2_n153 ) );
  OAI21_X1 u2_u13_u2_U47 (.A( u2_u13_u2_n140 ) , .ZN( u2_u13_u2_n141 ) , .B1( u2_u13_u2_n176 ) , .B2( u2_u13_u2_n177 ) );
  NOR3_X1 u2_u13_u2_U48 (.ZN( u2_u13_u2_n142 ) , .A3( u2_u13_u2_n175 ) , .A2( u2_u13_u2_n178 ) , .A1( u2_u13_u2_n181 ) );
  OAI21_X1 u2_u13_u2_U49 (.A( u2_u13_u2_n101 ) , .B2( u2_u13_u2_n121 ) , .B1( u2_u13_u2_n153 ) , .ZN( u2_u13_u2_n164 ) );
  NOR4_X1 u2_u13_u2_U5 (.A4( u2_u13_u2_n124 ) , .A3( u2_u13_u2_n125 ) , .A2( u2_u13_u2_n126 ) , .A1( u2_u13_u2_n127 ) , .ZN( u2_u13_u2_n128 ) );
  NAND2_X1 u2_u13_u2_U50 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n155 ) );
  NAND2_X1 u2_u13_u2_U51 (.A2( u2_u13_u2_n105 ) , .A1( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n143 ) );
  NAND2_X1 u2_u13_u2_U52 (.A1( u2_u13_u2_n104 ) , .A2( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n152 ) );
  NAND2_X1 u2_u13_u2_U53 (.A1( u2_u13_u2_n100 ) , .A2( u2_u13_u2_n105 ) , .ZN( u2_u13_u2_n132 ) );
  INV_X1 u2_u13_u2_U54 (.A( u2_u13_u2_n140 ) , .ZN( u2_u13_u2_n168 ) );
  INV_X1 u2_u13_u2_U55 (.A( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n167 ) );
  NAND2_X1 u2_u13_u2_U56 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n113 ) );
  NAND2_X1 u2_u13_u2_U57 (.A1( u2_u13_u2_n106 ) , .A2( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n131 ) );
  NAND2_X1 u2_u13_u2_U58 (.A1( u2_u13_u2_n103 ) , .A2( u2_u13_u2_n107 ) , .ZN( u2_u13_u2_n139 ) );
  NAND2_X1 u2_u13_u2_U59 (.A1( u2_u13_u2_n103 ) , .A2( u2_u13_u2_n105 ) , .ZN( u2_u13_u2_n133 ) );
  AOI21_X1 u2_u13_u2_U6 (.B2( u2_u13_u2_n119 ) , .ZN( u2_u13_u2_n127 ) , .A( u2_u13_u2_n137 ) , .B1( u2_u13_u2_n155 ) );
  NAND2_X1 u2_u13_u2_U60 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n103 ) , .ZN( u2_u13_u2_n154 ) );
  NAND2_X1 u2_u13_u2_U61 (.A2( u2_u13_u2_n103 ) , .A1( u2_u13_u2_n104 ) , .ZN( u2_u13_u2_n119 ) );
  NAND2_X1 u2_u13_u2_U62 (.A2( u2_u13_u2_n107 ) , .A1( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n123 ) );
  NAND2_X1 u2_u13_u2_U63 (.A1( u2_u13_u2_n104 ) , .A2( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n122 ) );
  INV_X1 u2_u13_u2_U64 (.A( u2_u13_u2_n114 ) , .ZN( u2_u13_u2_n172 ) );
  NAND2_X1 u2_u13_u2_U65 (.A2( u2_u13_u2_n100 ) , .A1( u2_u13_u2_n102 ) , .ZN( u2_u13_u2_n116 ) );
  NAND2_X1 u2_u13_u2_U66 (.A1( u2_u13_u2_n102 ) , .A2( u2_u13_u2_n108 ) , .ZN( u2_u13_u2_n120 ) );
  NAND2_X1 u2_u13_u2_U67 (.A2( u2_u13_u2_n105 ) , .A1( u2_u13_u2_n106 ) , .ZN( u2_u13_u2_n117 ) );
  INV_X1 u2_u13_u2_U68 (.ZN( u2_u13_u2_n187 ) , .A( u2_u13_u2_n99 ) );
  OAI21_X1 u2_u13_u2_U69 (.B1( u2_u13_u2_n137 ) , .B2( u2_u13_u2_n143 ) , .A( u2_u13_u2_n98 ) , .ZN( u2_u13_u2_n99 ) );
  AOI21_X1 u2_u13_u2_U7 (.ZN( u2_u13_u2_n124 ) , .B1( u2_u13_u2_n131 ) , .B2( u2_u13_u2_n143 ) , .A( u2_u13_u2_n172 ) );
  NOR2_X1 u2_u13_u2_U70 (.A2( u2_u13_X_16 ) , .ZN( u2_u13_u2_n140 ) , .A1( u2_u13_u2_n166 ) );
  NOR2_X1 u2_u13_u2_U71 (.A2( u2_u13_X_13 ) , .A1( u2_u13_X_14 ) , .ZN( u2_u13_u2_n100 ) );
  NOR2_X1 u2_u13_u2_U72 (.A2( u2_u13_X_16 ) , .A1( u2_u13_X_17 ) , .ZN( u2_u13_u2_n138 ) );
  NOR2_X1 u2_u13_u2_U73 (.A2( u2_u13_X_15 ) , .A1( u2_u13_X_18 ) , .ZN( u2_u13_u2_n104 ) );
  NOR2_X1 u2_u13_u2_U74 (.A2( u2_u13_X_14 ) , .ZN( u2_u13_u2_n103 ) , .A1( u2_u13_u2_n174 ) );
  NOR2_X1 u2_u13_u2_U75 (.A2( u2_u13_X_15 ) , .ZN( u2_u13_u2_n102 ) , .A1( u2_u13_u2_n165 ) );
  NOR2_X1 u2_u13_u2_U76 (.A2( u2_u13_X_17 ) , .ZN( u2_u13_u2_n114 ) , .A1( u2_u13_u2_n169 ) );
  AND2_X1 u2_u13_u2_U77 (.A1( u2_u13_X_15 ) , .ZN( u2_u13_u2_n105 ) , .A2( u2_u13_u2_n165 ) );
  AND2_X1 u2_u13_u2_U78 (.A2( u2_u13_X_15 ) , .A1( u2_u13_X_18 ) , .ZN( u2_u13_u2_n107 ) );
  AND2_X1 u2_u13_u2_U79 (.A1( u2_u13_X_14 ) , .ZN( u2_u13_u2_n106 ) , .A2( u2_u13_u2_n174 ) );
  AOI21_X1 u2_u13_u2_U8 (.B2( u2_u13_u2_n120 ) , .B1( u2_u13_u2_n121 ) , .ZN( u2_u13_u2_n126 ) , .A( u2_u13_u2_n167 ) );
  AND2_X1 u2_u13_u2_U80 (.A1( u2_u13_X_13 ) , .A2( u2_u13_X_14 ) , .ZN( u2_u13_u2_n108 ) );
  INV_X1 u2_u13_u2_U81 (.A( u2_u13_X_16 ) , .ZN( u2_u13_u2_n169 ) );
  INV_X1 u2_u13_u2_U82 (.A( u2_u13_X_17 ) , .ZN( u2_u13_u2_n166 ) );
  INV_X1 u2_u13_u2_U83 (.A( u2_u13_X_13 ) , .ZN( u2_u13_u2_n174 ) );
  INV_X1 u2_u13_u2_U84 (.A( u2_u13_X_18 ) , .ZN( u2_u13_u2_n165 ) );
  NAND4_X1 u2_u13_u2_U85 (.ZN( u2_out13_30 ) , .A4( u2_u13_u2_n147 ) , .A3( u2_u13_u2_n148 ) , .A2( u2_u13_u2_n149 ) , .A1( u2_u13_u2_n187 ) );
  AOI21_X1 u2_u13_u2_U86 (.B2( u2_u13_u2_n138 ) , .ZN( u2_u13_u2_n148 ) , .A( u2_u13_u2_n162 ) , .B1( u2_u13_u2_n182 ) );
  NOR3_X1 u2_u13_u2_U87 (.A3( u2_u13_u2_n144 ) , .A2( u2_u13_u2_n145 ) , .A1( u2_u13_u2_n146 ) , .ZN( u2_u13_u2_n147 ) );
  NAND4_X1 u2_u13_u2_U88 (.ZN( u2_out13_24 ) , .A4( u2_u13_u2_n111 ) , .A3( u2_u13_u2_n112 ) , .A1( u2_u13_u2_n130 ) , .A2( u2_u13_u2_n187 ) );
  AOI221_X1 u2_u13_u2_U89 (.A( u2_u13_u2_n109 ) , .B1( u2_u13_u2_n110 ) , .ZN( u2_u13_u2_n111 ) , .C1( u2_u13_u2_n134 ) , .C2( u2_u13_u2_n170 ) , .B2( u2_u13_u2_n173 ) );
  OAI22_X1 u2_u13_u2_U9 (.ZN( u2_u13_u2_n109 ) , .A2( u2_u13_u2_n113 ) , .B2( u2_u13_u2_n133 ) , .B1( u2_u13_u2_n167 ) , .A1( u2_u13_u2_n168 ) );
  AOI21_X1 u2_u13_u2_U90 (.ZN( u2_u13_u2_n112 ) , .B2( u2_u13_u2_n156 ) , .A( u2_u13_u2_n164 ) , .B1( u2_u13_u2_n181 ) );
  NAND4_X1 u2_u13_u2_U91 (.ZN( u2_out13_16 ) , .A4( u2_u13_u2_n128 ) , .A3( u2_u13_u2_n129 ) , .A1( u2_u13_u2_n130 ) , .A2( u2_u13_u2_n186 ) );
  AOI22_X1 u2_u13_u2_U92 (.A2( u2_u13_u2_n118 ) , .ZN( u2_u13_u2_n129 ) , .A1( u2_u13_u2_n140 ) , .B1( u2_u13_u2_n157 ) , .B2( u2_u13_u2_n170 ) );
  INV_X1 u2_u13_u2_U93 (.A( u2_u13_u2_n163 ) , .ZN( u2_u13_u2_n186 ) );
  OR4_X1 u2_u13_u2_U94 (.ZN( u2_out13_6 ) , .A4( u2_u13_u2_n161 ) , .A3( u2_u13_u2_n162 ) , .A2( u2_u13_u2_n163 ) , .A1( u2_u13_u2_n164 ) );
  OR3_X1 u2_u13_u2_U95 (.A2( u2_u13_u2_n159 ) , .A1( u2_u13_u2_n160 ) , .ZN( u2_u13_u2_n161 ) , .A3( u2_u13_u2_n183 ) );
  AOI21_X1 u2_u13_u2_U96 (.B2( u2_u13_u2_n154 ) , .B1( u2_u13_u2_n155 ) , .ZN( u2_u13_u2_n159 ) , .A( u2_u13_u2_n167 ) );
  NAND3_X1 u2_u13_u2_U97 (.A2( u2_u13_u2_n117 ) , .A1( u2_u13_u2_n122 ) , .A3( u2_u13_u2_n123 ) , .ZN( u2_u13_u2_n134 ) );
  NAND3_X1 u2_u13_u2_U98 (.ZN( u2_u13_u2_n110 ) , .A2( u2_u13_u2_n131 ) , .A3( u2_u13_u2_n139 ) , .A1( u2_u13_u2_n154 ) );
  NAND3_X1 u2_u13_u2_U99 (.A2( u2_u13_u2_n100 ) , .ZN( u2_u13_u2_n101 ) , .A1( u2_u13_u2_n104 ) , .A3( u2_u13_u2_n114 ) );
  OAI22_X1 u2_u13_u3_U10 (.B1( u2_u13_u3_n113 ) , .A2( u2_u13_u3_n135 ) , .A1( u2_u13_u3_n150 ) , .B2( u2_u13_u3_n164 ) , .ZN( u2_u13_u3_n98 ) );
  OAI211_X1 u2_u13_u3_U11 (.B( u2_u13_u3_n106 ) , .ZN( u2_u13_u3_n119 ) , .C2( u2_u13_u3_n128 ) , .C1( u2_u13_u3_n167 ) , .A( u2_u13_u3_n181 ) );
  AOI221_X1 u2_u13_u3_U12 (.C1( u2_u13_u3_n105 ) , .ZN( u2_u13_u3_n106 ) , .A( u2_u13_u3_n131 ) , .B2( u2_u13_u3_n132 ) , .C2( u2_u13_u3_n133 ) , .B1( u2_u13_u3_n169 ) );
  INV_X1 u2_u13_u3_U13 (.ZN( u2_u13_u3_n181 ) , .A( u2_u13_u3_n98 ) );
  NAND2_X1 u2_u13_u3_U14 (.ZN( u2_u13_u3_n105 ) , .A2( u2_u13_u3_n130 ) , .A1( u2_u13_u3_n155 ) );
  AOI22_X1 u2_u13_u3_U15 (.B1( u2_u13_u3_n115 ) , .A2( u2_u13_u3_n116 ) , .ZN( u2_u13_u3_n123 ) , .B2( u2_u13_u3_n133 ) , .A1( u2_u13_u3_n169 ) );
  NAND2_X1 u2_u13_u3_U16 (.ZN( u2_u13_u3_n116 ) , .A2( u2_u13_u3_n151 ) , .A1( u2_u13_u3_n182 ) );
  NOR2_X1 u2_u13_u3_U17 (.ZN( u2_u13_u3_n126 ) , .A2( u2_u13_u3_n150 ) , .A1( u2_u13_u3_n164 ) );
  AOI21_X1 u2_u13_u3_U18 (.ZN( u2_u13_u3_n112 ) , .B2( u2_u13_u3_n146 ) , .B1( u2_u13_u3_n155 ) , .A( u2_u13_u3_n167 ) );
  NAND2_X1 u2_u13_u3_U19 (.A1( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n142 ) , .A2( u2_u13_u3_n164 ) );
  NAND2_X1 u2_u13_u3_U20 (.ZN( u2_u13_u3_n132 ) , .A2( u2_u13_u3_n152 ) , .A1( u2_u13_u3_n156 ) );
  AND2_X1 u2_u13_u3_U21 (.A2( u2_u13_u3_n113 ) , .A1( u2_u13_u3_n114 ) , .ZN( u2_u13_u3_n151 ) );
  INV_X1 u2_u13_u3_U22 (.A( u2_u13_u3_n133 ) , .ZN( u2_u13_u3_n165 ) );
  INV_X1 u2_u13_u3_U23 (.A( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n170 ) );
  NAND2_X1 u2_u13_u3_U24 (.A1( u2_u13_u3_n107 ) , .A2( u2_u13_u3_n108 ) , .ZN( u2_u13_u3_n140 ) );
  NAND2_X1 u2_u13_u3_U25 (.ZN( u2_u13_u3_n117 ) , .A1( u2_u13_u3_n124 ) , .A2( u2_u13_u3_n148 ) );
  NAND2_X1 u2_u13_u3_U26 (.ZN( u2_u13_u3_n143 ) , .A1( u2_u13_u3_n165 ) , .A2( u2_u13_u3_n167 ) );
  INV_X1 u2_u13_u3_U27 (.A( u2_u13_u3_n130 ) , .ZN( u2_u13_u3_n177 ) );
  INV_X1 u2_u13_u3_U28 (.A( u2_u13_u3_n128 ) , .ZN( u2_u13_u3_n176 ) );
  INV_X1 u2_u13_u3_U29 (.A( u2_u13_u3_n155 ) , .ZN( u2_u13_u3_n174 ) );
  INV_X1 u2_u13_u3_U3 (.A( u2_u13_u3_n129 ) , .ZN( u2_u13_u3_n183 ) );
  INV_X1 u2_u13_u3_U30 (.A( u2_u13_u3_n139 ) , .ZN( u2_u13_u3_n185 ) );
  NOR2_X1 u2_u13_u3_U31 (.ZN( u2_u13_u3_n135 ) , .A2( u2_u13_u3_n141 ) , .A1( u2_u13_u3_n169 ) );
  OAI222_X1 u2_u13_u3_U32 (.C2( u2_u13_u3_n107 ) , .A2( u2_u13_u3_n108 ) , .B1( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n138 ) , .B2( u2_u13_u3_n146 ) , .C1( u2_u13_u3_n154 ) , .A1( u2_u13_u3_n164 ) );
  NOR4_X1 u2_u13_u3_U33 (.A4( u2_u13_u3_n157 ) , .A3( u2_u13_u3_n158 ) , .A2( u2_u13_u3_n159 ) , .A1( u2_u13_u3_n160 ) , .ZN( u2_u13_u3_n161 ) );
  AOI21_X1 u2_u13_u3_U34 (.B2( u2_u13_u3_n152 ) , .B1( u2_u13_u3_n153 ) , .ZN( u2_u13_u3_n158 ) , .A( u2_u13_u3_n164 ) );
  AOI21_X1 u2_u13_u3_U35 (.A( u2_u13_u3_n154 ) , .B2( u2_u13_u3_n155 ) , .B1( u2_u13_u3_n156 ) , .ZN( u2_u13_u3_n157 ) );
  AOI21_X1 u2_u13_u3_U36 (.A( u2_u13_u3_n149 ) , .B2( u2_u13_u3_n150 ) , .B1( u2_u13_u3_n151 ) , .ZN( u2_u13_u3_n159 ) );
  AOI211_X1 u2_u13_u3_U37 (.ZN( u2_u13_u3_n109 ) , .A( u2_u13_u3_n119 ) , .C2( u2_u13_u3_n129 ) , .B( u2_u13_u3_n138 ) , .C1( u2_u13_u3_n141 ) );
  AOI211_X1 u2_u13_u3_U38 (.B( u2_u13_u3_n119 ) , .A( u2_u13_u3_n120 ) , .C2( u2_u13_u3_n121 ) , .ZN( u2_u13_u3_n122 ) , .C1( u2_u13_u3_n179 ) );
  INV_X1 u2_u13_u3_U39 (.A( u2_u13_u3_n156 ) , .ZN( u2_u13_u3_n179 ) );
  INV_X1 u2_u13_u3_U4 (.A( u2_u13_u3_n140 ) , .ZN( u2_u13_u3_n182 ) );
  OAI22_X1 u2_u13_u3_U40 (.B1( u2_u13_u3_n118 ) , .ZN( u2_u13_u3_n120 ) , .A1( u2_u13_u3_n135 ) , .B2( u2_u13_u3_n154 ) , .A2( u2_u13_u3_n178 ) );
  AND3_X1 u2_u13_u3_U41 (.ZN( u2_u13_u3_n118 ) , .A2( u2_u13_u3_n124 ) , .A1( u2_u13_u3_n144 ) , .A3( u2_u13_u3_n152 ) );
  INV_X1 u2_u13_u3_U42 (.A( u2_u13_u3_n121 ) , .ZN( u2_u13_u3_n164 ) );
  NAND2_X1 u2_u13_u3_U43 (.ZN( u2_u13_u3_n133 ) , .A1( u2_u13_u3_n154 ) , .A2( u2_u13_u3_n164 ) );
  OAI211_X1 u2_u13_u3_U44 (.B( u2_u13_u3_n127 ) , .ZN( u2_u13_u3_n139 ) , .C1( u2_u13_u3_n150 ) , .C2( u2_u13_u3_n154 ) , .A( u2_u13_u3_n184 ) );
  INV_X1 u2_u13_u3_U45 (.A( u2_u13_u3_n125 ) , .ZN( u2_u13_u3_n184 ) );
  AOI221_X1 u2_u13_u3_U46 (.A( u2_u13_u3_n126 ) , .ZN( u2_u13_u3_n127 ) , .C2( u2_u13_u3_n132 ) , .C1( u2_u13_u3_n169 ) , .B2( u2_u13_u3_n170 ) , .B1( u2_u13_u3_n174 ) );
  OAI22_X1 u2_u13_u3_U47 (.A1( u2_u13_u3_n124 ) , .ZN( u2_u13_u3_n125 ) , .B2( u2_u13_u3_n145 ) , .A2( u2_u13_u3_n165 ) , .B1( u2_u13_u3_n167 ) );
  NOR2_X1 u2_u13_u3_U48 (.A1( u2_u13_u3_n113 ) , .ZN( u2_u13_u3_n131 ) , .A2( u2_u13_u3_n154 ) );
  NAND2_X1 u2_u13_u3_U49 (.A1( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n150 ) , .A2( u2_u13_u3_n99 ) );
  INV_X1 u2_u13_u3_U5 (.A( u2_u13_u3_n117 ) , .ZN( u2_u13_u3_n178 ) );
  NAND2_X1 u2_u13_u3_U50 (.A2( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n155 ) , .A1( u2_u13_u3_n97 ) );
  INV_X1 u2_u13_u3_U51 (.A( u2_u13_u3_n141 ) , .ZN( u2_u13_u3_n167 ) );
  AOI21_X1 u2_u13_u3_U52 (.B2( u2_u13_u3_n114 ) , .B1( u2_u13_u3_n146 ) , .A( u2_u13_u3_n154 ) , .ZN( u2_u13_u3_n94 ) );
  AOI21_X1 u2_u13_u3_U53 (.ZN( u2_u13_u3_n110 ) , .B2( u2_u13_u3_n142 ) , .B1( u2_u13_u3_n186 ) , .A( u2_u13_u3_n95 ) );
  INV_X1 u2_u13_u3_U54 (.A( u2_u13_u3_n145 ) , .ZN( u2_u13_u3_n186 ) );
  AOI21_X1 u2_u13_u3_U55 (.B1( u2_u13_u3_n124 ) , .A( u2_u13_u3_n149 ) , .B2( u2_u13_u3_n155 ) , .ZN( u2_u13_u3_n95 ) );
  INV_X1 u2_u13_u3_U56 (.A( u2_u13_u3_n149 ) , .ZN( u2_u13_u3_n169 ) );
  NAND2_X1 u2_u13_u3_U57 (.ZN( u2_u13_u3_n124 ) , .A1( u2_u13_u3_n96 ) , .A2( u2_u13_u3_n97 ) );
  NAND2_X1 u2_u13_u3_U58 (.A2( u2_u13_u3_n100 ) , .ZN( u2_u13_u3_n146 ) , .A1( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U59 (.A1( u2_u13_u3_n101 ) , .ZN( u2_u13_u3_n145 ) , .A2( u2_u13_u3_n99 ) );
  AOI221_X1 u2_u13_u3_U6 (.A( u2_u13_u3_n131 ) , .C2( u2_u13_u3_n132 ) , .C1( u2_u13_u3_n133 ) , .ZN( u2_u13_u3_n134 ) , .B1( u2_u13_u3_n143 ) , .B2( u2_u13_u3_n177 ) );
  NAND2_X1 u2_u13_u3_U60 (.A1( u2_u13_u3_n100 ) , .ZN( u2_u13_u3_n156 ) , .A2( u2_u13_u3_n99 ) );
  NAND2_X1 u2_u13_u3_U61 (.A2( u2_u13_u3_n101 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n148 ) );
  NAND2_X1 u2_u13_u3_U62 (.A1( u2_u13_u3_n100 ) , .A2( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n128 ) );
  NAND2_X1 u2_u13_u3_U63 (.A2( u2_u13_u3_n101 ) , .A1( u2_u13_u3_n102 ) , .ZN( u2_u13_u3_n152 ) );
  NAND2_X1 u2_u13_u3_U64 (.A2( u2_u13_u3_n101 ) , .ZN( u2_u13_u3_n114 ) , .A1( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U65 (.ZN( u2_u13_u3_n107 ) , .A1( u2_u13_u3_n97 ) , .A2( u2_u13_u3_n99 ) );
  NAND2_X1 u2_u13_u3_U66 (.A2( u2_u13_u3_n100 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n113 ) );
  NAND2_X1 u2_u13_u3_U67 (.A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n153 ) , .A2( u2_u13_u3_n97 ) );
  NAND2_X1 u2_u13_u3_U68 (.A2( u2_u13_u3_n103 ) , .A1( u2_u13_u3_n104 ) , .ZN( u2_u13_u3_n130 ) );
  NAND2_X1 u2_u13_u3_U69 (.A2( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n144 ) , .A1( u2_u13_u3_n96 ) );
  OAI22_X1 u2_u13_u3_U7 (.B2( u2_u13_u3_n147 ) , .A2( u2_u13_u3_n148 ) , .ZN( u2_u13_u3_n160 ) , .B1( u2_u13_u3_n165 ) , .A1( u2_u13_u3_n168 ) );
  NAND2_X1 u2_u13_u3_U70 (.A1( u2_u13_u3_n102 ) , .A2( u2_u13_u3_n103 ) , .ZN( u2_u13_u3_n108 ) );
  NOR2_X1 u2_u13_u3_U71 (.A2( u2_u13_X_19 ) , .A1( u2_u13_X_20 ) , .ZN( u2_u13_u3_n99 ) );
  NOR2_X1 u2_u13_u3_U72 (.A2( u2_u13_X_21 ) , .A1( u2_u13_X_24 ) , .ZN( u2_u13_u3_n103 ) );
  NOR2_X1 u2_u13_u3_U73 (.A2( u2_u13_X_24 ) , .A1( u2_u13_u3_n171 ) , .ZN( u2_u13_u3_n97 ) );
  NOR2_X1 u2_u13_u3_U74 (.A2( u2_u13_X_23 ) , .ZN( u2_u13_u3_n141 ) , .A1( u2_u13_u3_n166 ) );
  NOR2_X1 u2_u13_u3_U75 (.A2( u2_u13_X_19 ) , .A1( u2_u13_u3_n172 ) , .ZN( u2_u13_u3_n96 ) );
  NAND2_X1 u2_u13_u3_U76 (.A1( u2_u13_X_22 ) , .A2( u2_u13_X_23 ) , .ZN( u2_u13_u3_n154 ) );
  NAND2_X1 u2_u13_u3_U77 (.A1( u2_u13_X_23 ) , .ZN( u2_u13_u3_n149 ) , .A2( u2_u13_u3_n166 ) );
  NOR2_X1 u2_u13_u3_U78 (.A2( u2_u13_X_22 ) , .A1( u2_u13_X_23 ) , .ZN( u2_u13_u3_n121 ) );
  AND2_X1 u2_u13_u3_U79 (.A1( u2_u13_X_24 ) , .ZN( u2_u13_u3_n101 ) , .A2( u2_u13_u3_n171 ) );
  AND3_X1 u2_u13_u3_U8 (.A3( u2_u13_u3_n144 ) , .A2( u2_u13_u3_n145 ) , .A1( u2_u13_u3_n146 ) , .ZN( u2_u13_u3_n147 ) );
  AND2_X1 u2_u13_u3_U80 (.A1( u2_u13_X_19 ) , .ZN( u2_u13_u3_n102 ) , .A2( u2_u13_u3_n172 ) );
  AND2_X1 u2_u13_u3_U81 (.A1( u2_u13_X_21 ) , .A2( u2_u13_X_24 ) , .ZN( u2_u13_u3_n100 ) );
  AND2_X1 u2_u13_u3_U82 (.A2( u2_u13_X_19 ) , .A1( u2_u13_X_20 ) , .ZN( u2_u13_u3_n104 ) );
  INV_X1 u2_u13_u3_U83 (.A( u2_u13_X_22 ) , .ZN( u2_u13_u3_n166 ) );
  INV_X1 u2_u13_u3_U84 (.A( u2_u13_X_21 ) , .ZN( u2_u13_u3_n171 ) );
  INV_X1 u2_u13_u3_U85 (.A( u2_u13_X_20 ) , .ZN( u2_u13_u3_n172 ) );
  NAND4_X1 u2_u13_u3_U86 (.ZN( u2_out13_26 ) , .A4( u2_u13_u3_n109 ) , .A3( u2_u13_u3_n110 ) , .A2( u2_u13_u3_n111 ) , .A1( u2_u13_u3_n173 ) );
  INV_X1 u2_u13_u3_U87 (.ZN( u2_u13_u3_n173 ) , .A( u2_u13_u3_n94 ) );
  OAI21_X1 u2_u13_u3_U88 (.ZN( u2_u13_u3_n111 ) , .B2( u2_u13_u3_n117 ) , .A( u2_u13_u3_n133 ) , .B1( u2_u13_u3_n176 ) );
  NAND4_X1 u2_u13_u3_U89 (.ZN( u2_out13_20 ) , .A4( u2_u13_u3_n122 ) , .A3( u2_u13_u3_n123 ) , .A1( u2_u13_u3_n175 ) , .A2( u2_u13_u3_n180 ) );
  INV_X1 u2_u13_u3_U9 (.A( u2_u13_u3_n143 ) , .ZN( u2_u13_u3_n168 ) );
  INV_X1 u2_u13_u3_U90 (.A( u2_u13_u3_n112 ) , .ZN( u2_u13_u3_n175 ) );
  INV_X1 u2_u13_u3_U91 (.A( u2_u13_u3_n126 ) , .ZN( u2_u13_u3_n180 ) );
  NAND4_X1 u2_u13_u3_U92 (.ZN( u2_out13_1 ) , .A4( u2_u13_u3_n161 ) , .A3( u2_u13_u3_n162 ) , .A2( u2_u13_u3_n163 ) , .A1( u2_u13_u3_n185 ) );
  NAND2_X1 u2_u13_u3_U93 (.ZN( u2_u13_u3_n163 ) , .A2( u2_u13_u3_n170 ) , .A1( u2_u13_u3_n176 ) );
  AOI22_X1 u2_u13_u3_U94 (.B2( u2_u13_u3_n140 ) , .B1( u2_u13_u3_n141 ) , .A2( u2_u13_u3_n142 ) , .ZN( u2_u13_u3_n162 ) , .A1( u2_u13_u3_n177 ) );
  OR4_X1 u2_u13_u3_U95 (.ZN( u2_out13_10 ) , .A4( u2_u13_u3_n136 ) , .A3( u2_u13_u3_n137 ) , .A1( u2_u13_u3_n138 ) , .A2( u2_u13_u3_n139 ) );
  OAI222_X1 u2_u13_u3_U96 (.C1( u2_u13_u3_n128 ) , .ZN( u2_u13_u3_n137 ) , .B1( u2_u13_u3_n148 ) , .A2( u2_u13_u3_n150 ) , .B2( u2_u13_u3_n154 ) , .C2( u2_u13_u3_n164 ) , .A1( u2_u13_u3_n167 ) );
  OAI221_X1 u2_u13_u3_U97 (.A( u2_u13_u3_n134 ) , .B2( u2_u13_u3_n135 ) , .ZN( u2_u13_u3_n136 ) , .C1( u2_u13_u3_n149 ) , .B1( u2_u13_u3_n151 ) , .C2( u2_u13_u3_n183 ) );
  NAND3_X1 u2_u13_u3_U98 (.A1( u2_u13_u3_n114 ) , .ZN( u2_u13_u3_n115 ) , .A2( u2_u13_u3_n145 ) , .A3( u2_u13_u3_n153 ) );
  NAND3_X1 u2_u13_u3_U99 (.ZN( u2_u13_u3_n129 ) , .A2( u2_u13_u3_n144 ) , .A1( u2_u13_u3_n153 ) , .A3( u2_u13_u3_n182 ) );
  AOI22_X1 u2_u13_u6_U10 (.A2( u2_u13_u6_n151 ) , .B2( u2_u13_u6_n161 ) , .A1( u2_u13_u6_n167 ) , .B1( u2_u13_u6_n170 ) , .ZN( u2_u13_u6_n89 ) );
  AOI21_X1 u2_u13_u6_U11 (.B1( u2_u13_u6_n107 ) , .B2( u2_u13_u6_n132 ) , .A( u2_u13_u6_n158 ) , .ZN( u2_u13_u6_n88 ) );
  AOI21_X1 u2_u13_u6_U12 (.B2( u2_u13_u6_n147 ) , .B1( u2_u13_u6_n148 ) , .ZN( u2_u13_u6_n149 ) , .A( u2_u13_u6_n158 ) );
  AOI21_X1 u2_u13_u6_U13 (.ZN( u2_u13_u6_n106 ) , .A( u2_u13_u6_n142 ) , .B2( u2_u13_u6_n159 ) , .B1( u2_u13_u6_n164 ) );
  INV_X1 u2_u13_u6_U14 (.A( u2_u13_u6_n155 ) , .ZN( u2_u13_u6_n161 ) );
  INV_X1 u2_u13_u6_U15 (.A( u2_u13_u6_n128 ) , .ZN( u2_u13_u6_n164 ) );
  NAND2_X1 u2_u13_u6_U16 (.ZN( u2_u13_u6_n110 ) , .A1( u2_u13_u6_n122 ) , .A2( u2_u13_u6_n129 ) );
  NAND2_X1 u2_u13_u6_U17 (.ZN( u2_u13_u6_n124 ) , .A2( u2_u13_u6_n146 ) , .A1( u2_u13_u6_n148 ) );
  INV_X1 u2_u13_u6_U18 (.A( u2_u13_u6_n132 ) , .ZN( u2_u13_u6_n171 ) );
  AND2_X1 u2_u13_u6_U19 (.A1( u2_u13_u6_n100 ) , .ZN( u2_u13_u6_n130 ) , .A2( u2_u13_u6_n147 ) );
  INV_X1 u2_u13_u6_U20 (.A( u2_u13_u6_n127 ) , .ZN( u2_u13_u6_n173 ) );
  INV_X1 u2_u13_u6_U21 (.A( u2_u13_u6_n121 ) , .ZN( u2_u13_u6_n167 ) );
  INV_X1 u2_u13_u6_U22 (.A( u2_u13_u6_n100 ) , .ZN( u2_u13_u6_n169 ) );
  INV_X1 u2_u13_u6_U23 (.A( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n170 ) );
  INV_X1 u2_u13_u6_U24 (.A( u2_u13_u6_n113 ) , .ZN( u2_u13_u6_n168 ) );
  AND2_X1 u2_u13_u6_U25 (.A1( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n119 ) , .ZN( u2_u13_u6_n133 ) );
  AND2_X1 u2_u13_u6_U26 (.A2( u2_u13_u6_n121 ) , .A1( u2_u13_u6_n122 ) , .ZN( u2_u13_u6_n131 ) );
  AND3_X1 u2_u13_u6_U27 (.ZN( u2_u13_u6_n120 ) , .A2( u2_u13_u6_n127 ) , .A1( u2_u13_u6_n132 ) , .A3( u2_u13_u6_n145 ) );
  INV_X1 u2_u13_u6_U28 (.A( u2_u13_u6_n146 ) , .ZN( u2_u13_u6_n163 ) );
  AOI222_X1 u2_u13_u6_U29 (.ZN( u2_u13_u6_n114 ) , .A1( u2_u13_u6_n118 ) , .A2( u2_u13_u6_n126 ) , .B2( u2_u13_u6_n151 ) , .C2( u2_u13_u6_n159 ) , .C1( u2_u13_u6_n168 ) , .B1( u2_u13_u6_n169 ) );
  INV_X1 u2_u13_u6_U3 (.A( u2_u13_u6_n110 ) , .ZN( u2_u13_u6_n166 ) );
  NOR2_X1 u2_u13_u6_U30 (.A1( u2_u13_u6_n162 ) , .A2( u2_u13_u6_n165 ) , .ZN( u2_u13_u6_n98 ) );
  AOI211_X1 u2_u13_u6_U31 (.B( u2_u13_u6_n134 ) , .A( u2_u13_u6_n135 ) , .C1( u2_u13_u6_n136 ) , .ZN( u2_u13_u6_n137 ) , .C2( u2_u13_u6_n151 ) );
  AOI21_X1 u2_u13_u6_U32 (.B2( u2_u13_u6_n132 ) , .B1( u2_u13_u6_n133 ) , .ZN( u2_u13_u6_n134 ) , .A( u2_u13_u6_n158 ) );
  AOI21_X1 u2_u13_u6_U33 (.B1( u2_u13_u6_n131 ) , .ZN( u2_u13_u6_n135 ) , .A( u2_u13_u6_n144 ) , .B2( u2_u13_u6_n146 ) );
  NAND4_X1 u2_u13_u6_U34 (.A4( u2_u13_u6_n127 ) , .A3( u2_u13_u6_n128 ) , .A2( u2_u13_u6_n129 ) , .A1( u2_u13_u6_n130 ) , .ZN( u2_u13_u6_n136 ) );
  NAND2_X1 u2_u13_u6_U35 (.A1( u2_u13_u6_n144 ) , .ZN( u2_u13_u6_n151 ) , .A2( u2_u13_u6_n158 ) );
  NAND2_X1 u2_u13_u6_U36 (.ZN( u2_u13_u6_n132 ) , .A1( u2_u13_u6_n91 ) , .A2( u2_u13_u6_n97 ) );
  AOI22_X1 u2_u13_u6_U37 (.B2( u2_u13_u6_n110 ) , .B1( u2_u13_u6_n111 ) , .A1( u2_u13_u6_n112 ) , .ZN( u2_u13_u6_n115 ) , .A2( u2_u13_u6_n161 ) );
  NAND4_X1 u2_u13_u6_U38 (.A3( u2_u13_u6_n109 ) , .ZN( u2_u13_u6_n112 ) , .A4( u2_u13_u6_n132 ) , .A2( u2_u13_u6_n147 ) , .A1( u2_u13_u6_n166 ) );
  NOR2_X1 u2_u13_u6_U39 (.ZN( u2_u13_u6_n109 ) , .A1( u2_u13_u6_n170 ) , .A2( u2_u13_u6_n173 ) );
  INV_X1 u2_u13_u6_U4 (.A( u2_u13_u6_n142 ) , .ZN( u2_u13_u6_n174 ) );
  NOR2_X1 u2_u13_u6_U40 (.A2( u2_u13_u6_n126 ) , .ZN( u2_u13_u6_n155 ) , .A1( u2_u13_u6_n160 ) );
  NAND2_X1 u2_u13_u6_U41 (.ZN( u2_u13_u6_n146 ) , .A2( u2_u13_u6_n94 ) , .A1( u2_u13_u6_n99 ) );
  AOI21_X1 u2_u13_u6_U42 (.A( u2_u13_u6_n144 ) , .B2( u2_u13_u6_n145 ) , .B1( u2_u13_u6_n146 ) , .ZN( u2_u13_u6_n150 ) );
  INV_X1 u2_u13_u6_U43 (.A( u2_u13_u6_n111 ) , .ZN( u2_u13_u6_n158 ) );
  NAND2_X1 u2_u13_u6_U44 (.ZN( u2_u13_u6_n127 ) , .A1( u2_u13_u6_n91 ) , .A2( u2_u13_u6_n92 ) );
  NAND2_X1 u2_u13_u6_U45 (.ZN( u2_u13_u6_n129 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n96 ) );
  INV_X1 u2_u13_u6_U46 (.A( u2_u13_u6_n144 ) , .ZN( u2_u13_u6_n159 ) );
  NAND2_X1 u2_u13_u6_U47 (.ZN( u2_u13_u6_n145 ) , .A2( u2_u13_u6_n97 ) , .A1( u2_u13_u6_n98 ) );
  NAND2_X1 u2_u13_u6_U48 (.ZN( u2_u13_u6_n148 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n94 ) );
  NAND2_X1 u2_u13_u6_U49 (.ZN( u2_u13_u6_n108 ) , .A2( u2_u13_u6_n139 ) , .A1( u2_u13_u6_n144 ) );
  NAND2_X1 u2_u13_u6_U5 (.A2( u2_u13_u6_n143 ) , .ZN( u2_u13_u6_n152 ) , .A1( u2_u13_u6_n166 ) );
  NAND2_X1 u2_u13_u6_U50 (.ZN( u2_u13_u6_n121 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n97 ) );
  NAND2_X1 u2_u13_u6_U51 (.ZN( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n95 ) );
  AND2_X1 u2_u13_u6_U52 (.ZN( u2_u13_u6_n118 ) , .A2( u2_u13_u6_n91 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U53 (.ZN( u2_u13_u6_n147 ) , .A2( u2_u13_u6_n98 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U54 (.ZN( u2_u13_u6_n128 ) , .A1( u2_u13_u6_n94 ) , .A2( u2_u13_u6_n96 ) );
  NAND2_X1 u2_u13_u6_U55 (.ZN( u2_u13_u6_n119 ) , .A2( u2_u13_u6_n95 ) , .A1( u2_u13_u6_n99 ) );
  NAND2_X1 u2_u13_u6_U56 (.ZN( u2_u13_u6_n123 ) , .A2( u2_u13_u6_n91 ) , .A1( u2_u13_u6_n96 ) );
  NAND2_X1 u2_u13_u6_U57 (.ZN( u2_u13_u6_n100 ) , .A2( u2_u13_u6_n92 ) , .A1( u2_u13_u6_n98 ) );
  NAND2_X1 u2_u13_u6_U58 (.ZN( u2_u13_u6_n122 ) , .A1( u2_u13_u6_n94 ) , .A2( u2_u13_u6_n97 ) );
  INV_X1 u2_u13_u6_U59 (.A( u2_u13_u6_n139 ) , .ZN( u2_u13_u6_n160 ) );
  AOI22_X1 u2_u13_u6_U6 (.B2( u2_u13_u6_n101 ) , .A1( u2_u13_u6_n102 ) , .ZN( u2_u13_u6_n103 ) , .B1( u2_u13_u6_n160 ) , .A2( u2_u13_u6_n161 ) );
  NAND2_X1 u2_u13_u6_U60 (.ZN( u2_u13_u6_n113 ) , .A1( u2_u13_u6_n96 ) , .A2( u2_u13_u6_n98 ) );
  NOR2_X1 u2_u13_u6_U61 (.A2( u2_u13_X_40 ) , .A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n126 ) );
  NOR2_X1 u2_u13_u6_U62 (.A2( u2_u13_X_39 ) , .A1( u2_u13_X_42 ) , .ZN( u2_u13_u6_n92 ) );
  NOR2_X1 u2_u13_u6_U63 (.A2( u2_u13_X_39 ) , .A1( u2_u13_u6_n156 ) , .ZN( u2_u13_u6_n97 ) );
  NOR2_X1 u2_u13_u6_U64 (.A2( u2_u13_X_38 ) , .A1( u2_u13_u6_n165 ) , .ZN( u2_u13_u6_n95 ) );
  NOR2_X1 u2_u13_u6_U65 (.A2( u2_u13_X_41 ) , .ZN( u2_u13_u6_n111 ) , .A1( u2_u13_u6_n157 ) );
  NOR2_X1 u2_u13_u6_U66 (.A2( u2_u13_X_37 ) , .A1( u2_u13_u6_n162 ) , .ZN( u2_u13_u6_n94 ) );
  NOR2_X1 u2_u13_u6_U67 (.A2( u2_u13_X_37 ) , .A1( u2_u13_X_38 ) , .ZN( u2_u13_u6_n91 ) );
  NAND2_X1 u2_u13_u6_U68 (.A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n144 ) , .A2( u2_u13_u6_n157 ) );
  NAND2_X1 u2_u13_u6_U69 (.A2( u2_u13_X_40 ) , .A1( u2_u13_X_41 ) , .ZN( u2_u13_u6_n139 ) );
  NOR2_X1 u2_u13_u6_U7 (.A1( u2_u13_u6_n118 ) , .ZN( u2_u13_u6_n143 ) , .A2( u2_u13_u6_n168 ) );
  AND2_X1 u2_u13_u6_U70 (.A1( u2_u13_X_39 ) , .A2( u2_u13_u6_n156 ) , .ZN( u2_u13_u6_n96 ) );
  AND2_X1 u2_u13_u6_U71 (.A1( u2_u13_X_39 ) , .A2( u2_u13_X_42 ) , .ZN( u2_u13_u6_n99 ) );
  INV_X1 u2_u13_u6_U72 (.A( u2_u13_X_40 ) , .ZN( u2_u13_u6_n157 ) );
  INV_X1 u2_u13_u6_U73 (.A( u2_u13_X_37 ) , .ZN( u2_u13_u6_n165 ) );
  INV_X1 u2_u13_u6_U74 (.A( u2_u13_X_38 ) , .ZN( u2_u13_u6_n162 ) );
  INV_X1 u2_u13_u6_U75 (.A( u2_u13_X_42 ) , .ZN( u2_u13_u6_n156 ) );
  NAND4_X1 u2_u13_u6_U76 (.ZN( u2_out13_32 ) , .A4( u2_u13_u6_n103 ) , .A3( u2_u13_u6_n104 ) , .A2( u2_u13_u6_n105 ) , .A1( u2_u13_u6_n106 ) );
  AOI22_X1 u2_u13_u6_U77 (.ZN( u2_u13_u6_n105 ) , .A2( u2_u13_u6_n108 ) , .A1( u2_u13_u6_n118 ) , .B2( u2_u13_u6_n126 ) , .B1( u2_u13_u6_n171 ) );
  AOI22_X1 u2_u13_u6_U78 (.ZN( u2_u13_u6_n104 ) , .A1( u2_u13_u6_n111 ) , .B1( u2_u13_u6_n124 ) , .B2( u2_u13_u6_n151 ) , .A2( u2_u13_u6_n93 ) );
  NAND4_X1 u2_u13_u6_U79 (.ZN( u2_out13_12 ) , .A4( u2_u13_u6_n114 ) , .A3( u2_u13_u6_n115 ) , .A2( u2_u13_u6_n116 ) , .A1( u2_u13_u6_n117 ) );
  OAI21_X1 u2_u13_u6_U8 (.A( u2_u13_u6_n159 ) , .B1( u2_u13_u6_n169 ) , .B2( u2_u13_u6_n173 ) , .ZN( u2_u13_u6_n90 ) );
  OAI22_X1 u2_u13_u6_U80 (.B2( u2_u13_u6_n111 ) , .ZN( u2_u13_u6_n116 ) , .B1( u2_u13_u6_n126 ) , .A2( u2_u13_u6_n164 ) , .A1( u2_u13_u6_n167 ) );
  OAI21_X1 u2_u13_u6_U81 (.A( u2_u13_u6_n108 ) , .ZN( u2_u13_u6_n117 ) , .B2( u2_u13_u6_n141 ) , .B1( u2_u13_u6_n163 ) );
  OAI211_X1 u2_u13_u6_U82 (.ZN( u2_out13_7 ) , .B( u2_u13_u6_n153 ) , .C2( u2_u13_u6_n154 ) , .C1( u2_u13_u6_n155 ) , .A( u2_u13_u6_n174 ) );
  NOR3_X1 u2_u13_u6_U83 (.A1( u2_u13_u6_n141 ) , .ZN( u2_u13_u6_n154 ) , .A3( u2_u13_u6_n164 ) , .A2( u2_u13_u6_n171 ) );
  AOI211_X1 u2_u13_u6_U84 (.B( u2_u13_u6_n149 ) , .A( u2_u13_u6_n150 ) , .C2( u2_u13_u6_n151 ) , .C1( u2_u13_u6_n152 ) , .ZN( u2_u13_u6_n153 ) );
  OAI211_X1 u2_u13_u6_U85 (.ZN( u2_out13_22 ) , .B( u2_u13_u6_n137 ) , .A( u2_u13_u6_n138 ) , .C2( u2_u13_u6_n139 ) , .C1( u2_u13_u6_n140 ) );
  AOI22_X1 u2_u13_u6_U86 (.B1( u2_u13_u6_n124 ) , .A2( u2_u13_u6_n125 ) , .A1( u2_u13_u6_n126 ) , .ZN( u2_u13_u6_n138 ) , .B2( u2_u13_u6_n161 ) );
  AND4_X1 u2_u13_u6_U87 (.A3( u2_u13_u6_n119 ) , .A1( u2_u13_u6_n120 ) , .A4( u2_u13_u6_n129 ) , .ZN( u2_u13_u6_n140 ) , .A2( u2_u13_u6_n143 ) );
  NAND3_X1 u2_u13_u6_U88 (.A2( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n125 ) , .A1( u2_u13_u6_n130 ) , .A3( u2_u13_u6_n131 ) );
  NAND3_X1 u2_u13_u6_U89 (.A3( u2_u13_u6_n133 ) , .ZN( u2_u13_u6_n141 ) , .A1( u2_u13_u6_n145 ) , .A2( u2_u13_u6_n148 ) );
  INV_X1 u2_u13_u6_U9 (.ZN( u2_u13_u6_n172 ) , .A( u2_u13_u6_n88 ) );
  NAND3_X1 u2_u13_u6_U90 (.ZN( u2_u13_u6_n101 ) , .A3( u2_u13_u6_n107 ) , .A2( u2_u13_u6_n121 ) , .A1( u2_u13_u6_n127 ) );
  NAND3_X1 u2_u13_u6_U91 (.ZN( u2_u13_u6_n102 ) , .A3( u2_u13_u6_n130 ) , .A2( u2_u13_u6_n145 ) , .A1( u2_u13_u6_n166 ) );
  NAND3_X1 u2_u13_u6_U92 (.A3( u2_u13_u6_n113 ) , .A1( u2_u13_u6_n119 ) , .A2( u2_u13_u6_n123 ) , .ZN( u2_u13_u6_n93 ) );
  NAND3_X1 u2_u13_u6_U93 (.ZN( u2_u13_u6_n142 ) , .A2( u2_u13_u6_n172 ) , .A3( u2_u13_u6_n89 ) , .A1( u2_u13_u6_n90 ) );
  AND3_X1 u2_u13_u7_U10 (.A3( u2_u13_u7_n110 ) , .A2( u2_u13_u7_n127 ) , .A1( u2_u13_u7_n132 ) , .ZN( u2_u13_u7_n92 ) );
  OAI21_X1 u2_u13_u7_U11 (.A( u2_u13_u7_n161 ) , .B1( u2_u13_u7_n168 ) , .B2( u2_u13_u7_n173 ) , .ZN( u2_u13_u7_n91 ) );
  AOI211_X1 u2_u13_u7_U12 (.A( u2_u13_u7_n117 ) , .ZN( u2_u13_u7_n118 ) , .C2( u2_u13_u7_n126 ) , .C1( u2_u13_u7_n177 ) , .B( u2_u13_u7_n180 ) );
  OAI22_X1 u2_u13_u7_U13 (.B1( u2_u13_u7_n115 ) , .ZN( u2_u13_u7_n117 ) , .A2( u2_u13_u7_n133 ) , .A1( u2_u13_u7_n137 ) , .B2( u2_u13_u7_n162 ) );
  INV_X1 u2_u13_u7_U14 (.A( u2_u13_u7_n116 ) , .ZN( u2_u13_u7_n180 ) );
  NOR3_X1 u2_u13_u7_U15 (.ZN( u2_u13_u7_n115 ) , .A3( u2_u13_u7_n145 ) , .A2( u2_u13_u7_n168 ) , .A1( u2_u13_u7_n169 ) );
  OAI211_X1 u2_u13_u7_U16 (.B( u2_u13_u7_n122 ) , .A( u2_u13_u7_n123 ) , .C2( u2_u13_u7_n124 ) , .ZN( u2_u13_u7_n154 ) , .C1( u2_u13_u7_n162 ) );
  AOI222_X1 u2_u13_u7_U17 (.ZN( u2_u13_u7_n122 ) , .C2( u2_u13_u7_n126 ) , .C1( u2_u13_u7_n145 ) , .B1( u2_u13_u7_n161 ) , .A2( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n170 ) , .A1( u2_u13_u7_n176 ) );
  INV_X1 u2_u13_u7_U18 (.A( u2_u13_u7_n133 ) , .ZN( u2_u13_u7_n176 ) );
  NOR3_X1 u2_u13_u7_U19 (.A2( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n135 ) , .ZN( u2_u13_u7_n136 ) , .A3( u2_u13_u7_n171 ) );
  NOR2_X1 u2_u13_u7_U20 (.A1( u2_u13_u7_n130 ) , .A2( u2_u13_u7_n134 ) , .ZN( u2_u13_u7_n153 ) );
  INV_X1 u2_u13_u7_U21 (.A( u2_u13_u7_n101 ) , .ZN( u2_u13_u7_n165 ) );
  NOR2_X1 u2_u13_u7_U22 (.ZN( u2_u13_u7_n111 ) , .A2( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n169 ) );
  AOI21_X1 u2_u13_u7_U23 (.ZN( u2_u13_u7_n104 ) , .B2( u2_u13_u7_n112 ) , .B1( u2_u13_u7_n127 ) , .A( u2_u13_u7_n164 ) );
  AOI21_X1 u2_u13_u7_U24 (.ZN( u2_u13_u7_n106 ) , .B1( u2_u13_u7_n133 ) , .B2( u2_u13_u7_n146 ) , .A( u2_u13_u7_n162 ) );
  AOI21_X1 u2_u13_u7_U25 (.A( u2_u13_u7_n101 ) , .ZN( u2_u13_u7_n107 ) , .B2( u2_u13_u7_n128 ) , .B1( u2_u13_u7_n175 ) );
  INV_X1 u2_u13_u7_U26 (.A( u2_u13_u7_n138 ) , .ZN( u2_u13_u7_n171 ) );
  INV_X1 u2_u13_u7_U27 (.A( u2_u13_u7_n131 ) , .ZN( u2_u13_u7_n177 ) );
  INV_X1 u2_u13_u7_U28 (.A( u2_u13_u7_n110 ) , .ZN( u2_u13_u7_n174 ) );
  NAND2_X1 u2_u13_u7_U29 (.A1( u2_u13_u7_n129 ) , .A2( u2_u13_u7_n132 ) , .ZN( u2_u13_u7_n149 ) );
  OAI21_X1 u2_u13_u7_U3 (.ZN( u2_u13_u7_n159 ) , .A( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n171 ) , .B1( u2_u13_u7_n174 ) );
  NAND2_X1 u2_u13_u7_U30 (.A1( u2_u13_u7_n113 ) , .A2( u2_u13_u7_n124 ) , .ZN( u2_u13_u7_n130 ) );
  INV_X1 u2_u13_u7_U31 (.A( u2_u13_u7_n112 ) , .ZN( u2_u13_u7_n173 ) );
  INV_X1 u2_u13_u7_U32 (.A( u2_u13_u7_n128 ) , .ZN( u2_u13_u7_n168 ) );
  INV_X1 u2_u13_u7_U33 (.A( u2_u13_u7_n148 ) , .ZN( u2_u13_u7_n169 ) );
  INV_X1 u2_u13_u7_U34 (.A( u2_u13_u7_n127 ) , .ZN( u2_u13_u7_n179 ) );
  NOR2_X1 u2_u13_u7_U35 (.ZN( u2_u13_u7_n101 ) , .A2( u2_u13_u7_n150 ) , .A1( u2_u13_u7_n156 ) );
  AOI211_X1 u2_u13_u7_U36 (.B( u2_u13_u7_n154 ) , .A( u2_u13_u7_n155 ) , .C1( u2_u13_u7_n156 ) , .ZN( u2_u13_u7_n157 ) , .C2( u2_u13_u7_n172 ) );
  INV_X1 u2_u13_u7_U37 (.A( u2_u13_u7_n153 ) , .ZN( u2_u13_u7_n172 ) );
  AOI211_X1 u2_u13_u7_U38 (.B( u2_u13_u7_n139 ) , .A( u2_u13_u7_n140 ) , .C2( u2_u13_u7_n141 ) , .ZN( u2_u13_u7_n142 ) , .C1( u2_u13_u7_n156 ) );
  NAND4_X1 u2_u13_u7_U39 (.A3( u2_u13_u7_n127 ) , .A2( u2_u13_u7_n128 ) , .A1( u2_u13_u7_n129 ) , .ZN( u2_u13_u7_n141 ) , .A4( u2_u13_u7_n147 ) );
  INV_X1 u2_u13_u7_U4 (.A( u2_u13_u7_n111 ) , .ZN( u2_u13_u7_n170 ) );
  AOI21_X1 u2_u13_u7_U40 (.A( u2_u13_u7_n137 ) , .B1( u2_u13_u7_n138 ) , .ZN( u2_u13_u7_n139 ) , .B2( u2_u13_u7_n146 ) );
  OAI22_X1 u2_u13_u7_U41 (.B1( u2_u13_u7_n136 ) , .ZN( u2_u13_u7_n140 ) , .A1( u2_u13_u7_n153 ) , .B2( u2_u13_u7_n162 ) , .A2( u2_u13_u7_n164 ) );
  AOI21_X1 u2_u13_u7_U42 (.ZN( u2_u13_u7_n123 ) , .B1( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n177 ) , .A( u2_u13_u7_n97 ) );
  AOI21_X1 u2_u13_u7_U43 (.B2( u2_u13_u7_n113 ) , .B1( u2_u13_u7_n124 ) , .A( u2_u13_u7_n125 ) , .ZN( u2_u13_u7_n97 ) );
  INV_X1 u2_u13_u7_U44 (.A( u2_u13_u7_n125 ) , .ZN( u2_u13_u7_n161 ) );
  INV_X1 u2_u13_u7_U45 (.A( u2_u13_u7_n152 ) , .ZN( u2_u13_u7_n162 ) );
  AOI22_X1 u2_u13_u7_U46 (.A2( u2_u13_u7_n114 ) , .ZN( u2_u13_u7_n119 ) , .B1( u2_u13_u7_n130 ) , .A1( u2_u13_u7_n156 ) , .B2( u2_u13_u7_n165 ) );
  NAND2_X1 u2_u13_u7_U47 (.A2( u2_u13_u7_n112 ) , .ZN( u2_u13_u7_n114 ) , .A1( u2_u13_u7_n175 ) );
  AND2_X1 u2_u13_u7_U48 (.ZN( u2_u13_u7_n145 ) , .A2( u2_u13_u7_n98 ) , .A1( u2_u13_u7_n99 ) );
  NOR2_X1 u2_u13_u7_U49 (.ZN( u2_u13_u7_n137 ) , .A1( u2_u13_u7_n150 ) , .A2( u2_u13_u7_n161 ) );
  INV_X1 u2_u13_u7_U5 (.A( u2_u13_u7_n149 ) , .ZN( u2_u13_u7_n175 ) );
  AOI21_X1 u2_u13_u7_U50 (.ZN( u2_u13_u7_n105 ) , .B2( u2_u13_u7_n110 ) , .A( u2_u13_u7_n125 ) , .B1( u2_u13_u7_n147 ) );
  NAND2_X1 u2_u13_u7_U51 (.ZN( u2_u13_u7_n146 ) , .A1( u2_u13_u7_n95 ) , .A2( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U52 (.A2( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n147 ) , .A1( u2_u13_u7_n93 ) );
  NAND2_X1 u2_u13_u7_U53 (.A1( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n127 ) , .A2( u2_u13_u7_n99 ) );
  OR2_X1 u2_u13_u7_U54 (.ZN( u2_u13_u7_n126 ) , .A2( u2_u13_u7_n152 ) , .A1( u2_u13_u7_n156 ) );
  NAND2_X1 u2_u13_u7_U55 (.A2( u2_u13_u7_n102 ) , .A1( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n133 ) );
  NAND2_X1 u2_u13_u7_U56 (.ZN( u2_u13_u7_n112 ) , .A2( u2_u13_u7_n96 ) , .A1( u2_u13_u7_n99 ) );
  NAND2_X1 u2_u13_u7_U57 (.A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n128 ) , .A1( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U58 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n113 ) , .A2( u2_u13_u7_n93 ) );
  NAND2_X1 u2_u13_u7_U59 (.A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n124 ) , .A1( u2_u13_u7_n96 ) );
  INV_X1 u2_u13_u7_U6 (.A( u2_u13_u7_n154 ) , .ZN( u2_u13_u7_n178 ) );
  NAND2_X1 u2_u13_u7_U60 (.ZN( u2_u13_u7_n110 ) , .A1( u2_u13_u7_n95 ) , .A2( u2_u13_u7_n96 ) );
  INV_X1 u2_u13_u7_U61 (.A( u2_u13_u7_n150 ) , .ZN( u2_u13_u7_n164 ) );
  AND2_X1 u2_u13_u7_U62 (.ZN( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n93 ) , .A2( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U63 (.A1( u2_u13_u7_n100 ) , .A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n129 ) );
  NAND2_X1 u2_u13_u7_U64 (.A2( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n131 ) , .A1( u2_u13_u7_n95 ) );
  NAND2_X1 u2_u13_u7_U65 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n138 ) , .A2( u2_u13_u7_n99 ) );
  NAND2_X1 u2_u13_u7_U66 (.ZN( u2_u13_u7_n132 ) , .A1( u2_u13_u7_n93 ) , .A2( u2_u13_u7_n96 ) );
  NAND2_X1 u2_u13_u7_U67 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n148 ) , .A2( u2_u13_u7_n95 ) );
  NOR2_X1 u2_u13_u7_U68 (.A2( u2_u13_X_47 ) , .ZN( u2_u13_u7_n150 ) , .A1( u2_u13_u7_n163 ) );
  NOR2_X1 u2_u13_u7_U69 (.A2( u2_u13_X_43 ) , .A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n103 ) );
  AOI211_X1 u2_u13_u7_U7 (.ZN( u2_u13_u7_n116 ) , .A( u2_u13_u7_n155 ) , .C1( u2_u13_u7_n161 ) , .C2( u2_u13_u7_n171 ) , .B( u2_u13_u7_n94 ) );
  NOR2_X1 u2_u13_u7_U70 (.A2( u2_u13_X_48 ) , .A1( u2_u13_u7_n166 ) , .ZN( u2_u13_u7_n95 ) );
  NOR2_X1 u2_u13_u7_U71 (.A2( u2_u13_X_45 ) , .A1( u2_u13_X_48 ) , .ZN( u2_u13_u7_n99 ) );
  NOR2_X1 u2_u13_u7_U72 (.A2( u2_u13_X_44 ) , .A1( u2_u13_u7_n167 ) , .ZN( u2_u13_u7_n98 ) );
  NOR2_X1 u2_u13_u7_U73 (.A2( u2_u13_X_46 ) , .A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n152 ) );
  AND2_X1 u2_u13_u7_U74 (.A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n156 ) , .A2( u2_u13_u7_n163 ) );
  NAND2_X1 u2_u13_u7_U75 (.A2( u2_u13_X_46 ) , .A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n125 ) );
  AND2_X1 u2_u13_u7_U76 (.A2( u2_u13_X_45 ) , .A1( u2_u13_X_48 ) , .ZN( u2_u13_u7_n102 ) );
  AND2_X1 u2_u13_u7_U77 (.A2( u2_u13_X_43 ) , .A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n96 ) );
  AND2_X1 u2_u13_u7_U78 (.A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n100 ) , .A2( u2_u13_u7_n167 ) );
  AND2_X1 u2_u13_u7_U79 (.A1( u2_u13_X_48 ) , .A2( u2_u13_u7_n166 ) , .ZN( u2_u13_u7_n93 ) );
  OAI222_X1 u2_u13_u7_U8 (.C2( u2_u13_u7_n101 ) , .B2( u2_u13_u7_n111 ) , .A1( u2_u13_u7_n113 ) , .C1( u2_u13_u7_n146 ) , .A2( u2_u13_u7_n162 ) , .B1( u2_u13_u7_n164 ) , .ZN( u2_u13_u7_n94 ) );
  INV_X1 u2_u13_u7_U80 (.A( u2_u13_X_46 ) , .ZN( u2_u13_u7_n163 ) );
  INV_X1 u2_u13_u7_U81 (.A( u2_u13_X_43 ) , .ZN( u2_u13_u7_n167 ) );
  INV_X1 u2_u13_u7_U82 (.A( u2_u13_X_45 ) , .ZN( u2_u13_u7_n166 ) );
  NAND4_X1 u2_u13_u7_U83 (.ZN( u2_out13_27 ) , .A4( u2_u13_u7_n118 ) , .A3( u2_u13_u7_n119 ) , .A2( u2_u13_u7_n120 ) , .A1( u2_u13_u7_n121 ) );
  OAI21_X1 u2_u13_u7_U84 (.ZN( u2_u13_u7_n121 ) , .B2( u2_u13_u7_n145 ) , .A( u2_u13_u7_n150 ) , .B1( u2_u13_u7_n174 ) );
  OAI21_X1 u2_u13_u7_U85 (.ZN( u2_u13_u7_n120 ) , .A( u2_u13_u7_n161 ) , .B2( u2_u13_u7_n170 ) , .B1( u2_u13_u7_n179 ) );
  NAND4_X1 u2_u13_u7_U86 (.ZN( u2_out13_21 ) , .A4( u2_u13_u7_n157 ) , .A3( u2_u13_u7_n158 ) , .A2( u2_u13_u7_n159 ) , .A1( u2_u13_u7_n160 ) );
  OAI21_X1 u2_u13_u7_U87 (.B1( u2_u13_u7_n145 ) , .ZN( u2_u13_u7_n160 ) , .A( u2_u13_u7_n161 ) , .B2( u2_u13_u7_n177 ) );
  AOI22_X1 u2_u13_u7_U88 (.B2( u2_u13_u7_n149 ) , .B1( u2_u13_u7_n150 ) , .A2( u2_u13_u7_n151 ) , .A1( u2_u13_u7_n152 ) , .ZN( u2_u13_u7_n158 ) );
  NAND4_X1 u2_u13_u7_U89 (.ZN( u2_out13_15 ) , .A4( u2_u13_u7_n142 ) , .A3( u2_u13_u7_n143 ) , .A2( u2_u13_u7_n144 ) , .A1( u2_u13_u7_n178 ) );
  OAI221_X1 u2_u13_u7_U9 (.C1( u2_u13_u7_n101 ) , .C2( u2_u13_u7_n147 ) , .ZN( u2_u13_u7_n155 ) , .B2( u2_u13_u7_n162 ) , .A( u2_u13_u7_n91 ) , .B1( u2_u13_u7_n92 ) );
  OR2_X1 u2_u13_u7_U90 (.A2( u2_u13_u7_n125 ) , .A1( u2_u13_u7_n129 ) , .ZN( u2_u13_u7_n144 ) );
  AOI22_X1 u2_u13_u7_U91 (.A2( u2_u13_u7_n126 ) , .ZN( u2_u13_u7_n143 ) , .B2( u2_u13_u7_n165 ) , .B1( u2_u13_u7_n173 ) , .A1( u2_u13_u7_n174 ) );
  NAND4_X1 u2_u13_u7_U92 (.ZN( u2_out13_5 ) , .A4( u2_u13_u7_n108 ) , .A3( u2_u13_u7_n109 ) , .A1( u2_u13_u7_n116 ) , .A2( u2_u13_u7_n123 ) );
  AOI22_X1 u2_u13_u7_U93 (.ZN( u2_u13_u7_n109 ) , .A2( u2_u13_u7_n126 ) , .B2( u2_u13_u7_n145 ) , .B1( u2_u13_u7_n156 ) , .A1( u2_u13_u7_n171 ) );
  NOR4_X1 u2_u13_u7_U94 (.A4( u2_u13_u7_n104 ) , .A3( u2_u13_u7_n105 ) , .A2( u2_u13_u7_n106 ) , .A1( u2_u13_u7_n107 ) , .ZN( u2_u13_u7_n108 ) );
  NAND3_X1 u2_u13_u7_U95 (.A3( u2_u13_u7_n146 ) , .A2( u2_u13_u7_n147 ) , .A1( u2_u13_u7_n148 ) , .ZN( u2_u13_u7_n151 ) );
  NAND3_X1 u2_u13_u7_U96 (.A3( u2_u13_u7_n131 ) , .A2( u2_u13_u7_n132 ) , .A1( u2_u13_u7_n133 ) , .ZN( u2_u13_u7_n135 ) );
  XOR2_X1 u2_u1_U20 (.B( u2_K2_36 ) , .A( u2_R0_25 ) , .Z( u2_u1_X_36 ) );
  XOR2_X1 u2_u1_U21 (.B( u2_K2_35 ) , .A( u2_R0_24 ) , .Z( u2_u1_X_35 ) );
  XOR2_X1 u2_u1_U22 (.B( u2_K2_34 ) , .A( u2_R0_23 ) , .Z( u2_u1_X_34 ) );
  XOR2_X1 u2_u1_U23 (.B( u2_K2_33 ) , .A( u2_R0_22 ) , .Z( u2_u1_X_33 ) );
  XOR2_X1 u2_u1_U24 (.B( u2_K2_32 ) , .A( u2_R0_21 ) , .Z( u2_u1_X_32 ) );
  XOR2_X1 u2_u1_U25 (.B( u2_K2_31 ) , .A( u2_R0_20 ) , .Z( u2_u1_X_31 ) );
  INV_X1 u2_u1_u5_U10 (.A( u2_u1_u5_n121 ) , .ZN( u2_u1_u5_n177 ) );
  NOR3_X1 u2_u1_u5_U100 (.A3( u2_u1_u5_n141 ) , .A1( u2_u1_u5_n142 ) , .ZN( u2_u1_u5_n143 ) , .A2( u2_u1_u5_n191 ) );
  NAND4_X1 u2_u1_u5_U101 (.ZN( u2_out1_4 ) , .A4( u2_u1_u5_n112 ) , .A2( u2_u1_u5_n113 ) , .A1( u2_u1_u5_n114 ) , .A3( u2_u1_u5_n195 ) );
  AOI211_X1 u2_u1_u5_U102 (.A( u2_u1_u5_n110 ) , .C1( u2_u1_u5_n111 ) , .ZN( u2_u1_u5_n112 ) , .B( u2_u1_u5_n118 ) , .C2( u2_u1_u5_n177 ) );
  AOI222_X1 u2_u1_u5_U103 (.ZN( u2_u1_u5_n113 ) , .A1( u2_u1_u5_n131 ) , .C1( u2_u1_u5_n148 ) , .B2( u2_u1_u5_n174 ) , .C2( u2_u1_u5_n178 ) , .A2( u2_u1_u5_n179 ) , .B1( u2_u1_u5_n99 ) );
  NAND3_X1 u2_u1_u5_U104 (.A2( u2_u1_u5_n154 ) , .A3( u2_u1_u5_n158 ) , .A1( u2_u1_u5_n161 ) , .ZN( u2_u1_u5_n99 ) );
  NOR2_X1 u2_u1_u5_U11 (.ZN( u2_u1_u5_n160 ) , .A2( u2_u1_u5_n173 ) , .A1( u2_u1_u5_n177 ) );
  INV_X1 u2_u1_u5_U12 (.A( u2_u1_u5_n150 ) , .ZN( u2_u1_u5_n174 ) );
  AOI21_X1 u2_u1_u5_U13 (.A( u2_u1_u5_n160 ) , .B2( u2_u1_u5_n161 ) , .ZN( u2_u1_u5_n162 ) , .B1( u2_u1_u5_n192 ) );
  INV_X1 u2_u1_u5_U14 (.A( u2_u1_u5_n159 ) , .ZN( u2_u1_u5_n192 ) );
  AOI21_X1 u2_u1_u5_U15 (.A( u2_u1_u5_n156 ) , .B2( u2_u1_u5_n157 ) , .B1( u2_u1_u5_n158 ) , .ZN( u2_u1_u5_n163 ) );
  AOI21_X1 u2_u1_u5_U16 (.B2( u2_u1_u5_n139 ) , .B1( u2_u1_u5_n140 ) , .ZN( u2_u1_u5_n141 ) , .A( u2_u1_u5_n150 ) );
  OAI21_X1 u2_u1_u5_U17 (.A( u2_u1_u5_n133 ) , .B2( u2_u1_u5_n134 ) , .B1( u2_u1_u5_n135 ) , .ZN( u2_u1_u5_n142 ) );
  OAI21_X1 u2_u1_u5_U18 (.ZN( u2_u1_u5_n133 ) , .B2( u2_u1_u5_n147 ) , .A( u2_u1_u5_n173 ) , .B1( u2_u1_u5_n188 ) );
  NAND2_X1 u2_u1_u5_U19 (.A2( u2_u1_u5_n119 ) , .A1( u2_u1_u5_n123 ) , .ZN( u2_u1_u5_n137 ) );
  INV_X1 u2_u1_u5_U20 (.A( u2_u1_u5_n155 ) , .ZN( u2_u1_u5_n194 ) );
  NAND2_X1 u2_u1_u5_U21 (.A1( u2_u1_u5_n121 ) , .ZN( u2_u1_u5_n132 ) , .A2( u2_u1_u5_n172 ) );
  NAND2_X1 u2_u1_u5_U22 (.A2( u2_u1_u5_n122 ) , .ZN( u2_u1_u5_n136 ) , .A1( u2_u1_u5_n154 ) );
  NAND2_X1 u2_u1_u5_U23 (.A2( u2_u1_u5_n119 ) , .A1( u2_u1_u5_n120 ) , .ZN( u2_u1_u5_n159 ) );
  INV_X1 u2_u1_u5_U24 (.A( u2_u1_u5_n156 ) , .ZN( u2_u1_u5_n175 ) );
  INV_X1 u2_u1_u5_U25 (.A( u2_u1_u5_n158 ) , .ZN( u2_u1_u5_n188 ) );
  INV_X1 u2_u1_u5_U26 (.A( u2_u1_u5_n152 ) , .ZN( u2_u1_u5_n179 ) );
  INV_X1 u2_u1_u5_U27 (.A( u2_u1_u5_n140 ) , .ZN( u2_u1_u5_n182 ) );
  INV_X1 u2_u1_u5_U28 (.A( u2_u1_u5_n151 ) , .ZN( u2_u1_u5_n183 ) );
  INV_X1 u2_u1_u5_U29 (.A( u2_u1_u5_n123 ) , .ZN( u2_u1_u5_n185 ) );
  NOR2_X1 u2_u1_u5_U3 (.ZN( u2_u1_u5_n134 ) , .A1( u2_u1_u5_n183 ) , .A2( u2_u1_u5_n190 ) );
  INV_X1 u2_u1_u5_U30 (.A( u2_u1_u5_n161 ) , .ZN( u2_u1_u5_n184 ) );
  INV_X1 u2_u1_u5_U31 (.A( u2_u1_u5_n139 ) , .ZN( u2_u1_u5_n189 ) );
  INV_X1 u2_u1_u5_U32 (.A( u2_u1_u5_n157 ) , .ZN( u2_u1_u5_n190 ) );
  INV_X1 u2_u1_u5_U33 (.A( u2_u1_u5_n120 ) , .ZN( u2_u1_u5_n193 ) );
  NAND2_X1 u2_u1_u5_U34 (.ZN( u2_u1_u5_n111 ) , .A1( u2_u1_u5_n140 ) , .A2( u2_u1_u5_n155 ) );
  INV_X1 u2_u1_u5_U35 (.A( u2_u1_u5_n117 ) , .ZN( u2_u1_u5_n196 ) );
  OAI221_X1 u2_u1_u5_U36 (.A( u2_u1_u5_n116 ) , .ZN( u2_u1_u5_n117 ) , .B2( u2_u1_u5_n119 ) , .C1( u2_u1_u5_n153 ) , .C2( u2_u1_u5_n158 ) , .B1( u2_u1_u5_n172 ) );
  AOI222_X1 u2_u1_u5_U37 (.ZN( u2_u1_u5_n116 ) , .B2( u2_u1_u5_n145 ) , .C1( u2_u1_u5_n148 ) , .A2( u2_u1_u5_n174 ) , .C2( u2_u1_u5_n177 ) , .B1( u2_u1_u5_n187 ) , .A1( u2_u1_u5_n193 ) );
  INV_X1 u2_u1_u5_U38 (.A( u2_u1_u5_n115 ) , .ZN( u2_u1_u5_n187 ) );
  NOR2_X1 u2_u1_u5_U39 (.ZN( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n170 ) , .A2( u2_u1_u5_n180 ) );
  INV_X1 u2_u1_u5_U4 (.A( u2_u1_u5_n138 ) , .ZN( u2_u1_u5_n191 ) );
  AOI22_X1 u2_u1_u5_U40 (.B2( u2_u1_u5_n131 ) , .A2( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n169 ) , .B1( u2_u1_u5_n174 ) , .A1( u2_u1_u5_n185 ) );
  NOR2_X1 u2_u1_u5_U41 (.A1( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n150 ) , .A2( u2_u1_u5_n173 ) );
  AOI21_X1 u2_u1_u5_U42 (.A( u2_u1_u5_n118 ) , .B2( u2_u1_u5_n145 ) , .ZN( u2_u1_u5_n168 ) , .B1( u2_u1_u5_n186 ) );
  INV_X1 u2_u1_u5_U43 (.A( u2_u1_u5_n122 ) , .ZN( u2_u1_u5_n186 ) );
  NOR2_X1 u2_u1_u5_U44 (.A1( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n152 ) , .A2( u2_u1_u5_n176 ) );
  NOR2_X1 u2_u1_u5_U45 (.A1( u2_u1_u5_n115 ) , .ZN( u2_u1_u5_n118 ) , .A2( u2_u1_u5_n153 ) );
  NOR2_X1 u2_u1_u5_U46 (.A2( u2_u1_u5_n145 ) , .ZN( u2_u1_u5_n156 ) , .A1( u2_u1_u5_n174 ) );
  NOR2_X1 u2_u1_u5_U47 (.ZN( u2_u1_u5_n121 ) , .A2( u2_u1_u5_n145 ) , .A1( u2_u1_u5_n176 ) );
  AOI22_X1 u2_u1_u5_U48 (.ZN( u2_u1_u5_n114 ) , .A2( u2_u1_u5_n137 ) , .A1( u2_u1_u5_n145 ) , .B2( u2_u1_u5_n175 ) , .B1( u2_u1_u5_n193 ) );
  OAI211_X1 u2_u1_u5_U49 (.B( u2_u1_u5_n124 ) , .A( u2_u1_u5_n125 ) , .C2( u2_u1_u5_n126 ) , .C1( u2_u1_u5_n127 ) , .ZN( u2_u1_u5_n128 ) );
  OAI21_X1 u2_u1_u5_U5 (.B2( u2_u1_u5_n136 ) , .B1( u2_u1_u5_n137 ) , .ZN( u2_u1_u5_n138 ) , .A( u2_u1_u5_n177 ) );
  OAI21_X1 u2_u1_u5_U50 (.ZN( u2_u1_u5_n124 ) , .A( u2_u1_u5_n177 ) , .B2( u2_u1_u5_n183 ) , .B1( u2_u1_u5_n189 ) );
  NOR3_X1 u2_u1_u5_U51 (.ZN( u2_u1_u5_n127 ) , .A1( u2_u1_u5_n136 ) , .A3( u2_u1_u5_n148 ) , .A2( u2_u1_u5_n182 ) );
  OAI21_X1 u2_u1_u5_U52 (.ZN( u2_u1_u5_n125 ) , .A( u2_u1_u5_n174 ) , .B2( u2_u1_u5_n185 ) , .B1( u2_u1_u5_n190 ) );
  AOI21_X1 u2_u1_u5_U53 (.A( u2_u1_u5_n153 ) , .B2( u2_u1_u5_n154 ) , .B1( u2_u1_u5_n155 ) , .ZN( u2_u1_u5_n164 ) );
  AOI21_X1 u2_u1_u5_U54 (.ZN( u2_u1_u5_n110 ) , .B1( u2_u1_u5_n122 ) , .B2( u2_u1_u5_n139 ) , .A( u2_u1_u5_n153 ) );
  INV_X1 u2_u1_u5_U55 (.A( u2_u1_u5_n153 ) , .ZN( u2_u1_u5_n176 ) );
  INV_X1 u2_u1_u5_U56 (.A( u2_u1_u5_n126 ) , .ZN( u2_u1_u5_n173 ) );
  AND2_X1 u2_u1_u5_U57 (.A2( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n107 ) , .ZN( u2_u1_u5_n147 ) );
  AND2_X1 u2_u1_u5_U58 (.A2( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n108 ) , .ZN( u2_u1_u5_n148 ) );
  NAND2_X1 u2_u1_u5_U59 (.A1( u2_u1_u5_n105 ) , .A2( u2_u1_u5_n106 ) , .ZN( u2_u1_u5_n158 ) );
  INV_X1 u2_u1_u5_U6 (.A( u2_u1_u5_n135 ) , .ZN( u2_u1_u5_n178 ) );
  NAND2_X1 u2_u1_u5_U60 (.A2( u2_u1_u5_n108 ) , .A1( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n139 ) );
  NAND2_X1 u2_u1_u5_U61 (.A1( u2_u1_u5_n106 ) , .A2( u2_u1_u5_n108 ) , .ZN( u2_u1_u5_n119 ) );
  NAND2_X1 u2_u1_u5_U62 (.A2( u2_u1_u5_n103 ) , .A1( u2_u1_u5_n105 ) , .ZN( u2_u1_u5_n140 ) );
  NAND2_X1 u2_u1_u5_U63 (.A2( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n105 ) , .ZN( u2_u1_u5_n155 ) );
  NAND2_X1 u2_u1_u5_U64 (.A2( u2_u1_u5_n106 ) , .A1( u2_u1_u5_n107 ) , .ZN( u2_u1_u5_n122 ) );
  NAND2_X1 u2_u1_u5_U65 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n106 ) , .ZN( u2_u1_u5_n115 ) );
  NAND2_X1 u2_u1_u5_U66 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n103 ) , .ZN( u2_u1_u5_n161 ) );
  NAND2_X1 u2_u1_u5_U67 (.A1( u2_u1_u5_n105 ) , .A2( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n154 ) );
  INV_X1 u2_u1_u5_U68 (.A( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n172 ) );
  NAND2_X1 u2_u1_u5_U69 (.A1( u2_u1_u5_n103 ) , .A2( u2_u1_u5_n108 ) , .ZN( u2_u1_u5_n123 ) );
  OAI22_X1 u2_u1_u5_U7 (.B2( u2_u1_u5_n149 ) , .B1( u2_u1_u5_n150 ) , .A2( u2_u1_u5_n151 ) , .A1( u2_u1_u5_n152 ) , .ZN( u2_u1_u5_n165 ) );
  NAND2_X1 u2_u1_u5_U70 (.A2( u2_u1_u5_n103 ) , .A1( u2_u1_u5_n107 ) , .ZN( u2_u1_u5_n151 ) );
  NAND2_X1 u2_u1_u5_U71 (.A2( u2_u1_u5_n107 ) , .A1( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n120 ) );
  NAND2_X1 u2_u1_u5_U72 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n157 ) );
  AND2_X1 u2_u1_u5_U73 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n104 ) , .ZN( u2_u1_u5_n131 ) );
  INV_X1 u2_u1_u5_U74 (.A( u2_u1_u5_n102 ) , .ZN( u2_u1_u5_n195 ) );
  OAI221_X1 u2_u1_u5_U75 (.A( u2_u1_u5_n101 ) , .ZN( u2_u1_u5_n102 ) , .C2( u2_u1_u5_n115 ) , .C1( u2_u1_u5_n126 ) , .B1( u2_u1_u5_n134 ) , .B2( u2_u1_u5_n160 ) );
  OAI21_X1 u2_u1_u5_U76 (.ZN( u2_u1_u5_n101 ) , .B1( u2_u1_u5_n137 ) , .A( u2_u1_u5_n146 ) , .B2( u2_u1_u5_n147 ) );
  NOR2_X1 u2_u1_u5_U77 (.A2( u2_u1_X_34 ) , .A1( u2_u1_X_35 ) , .ZN( u2_u1_u5_n145 ) );
  NOR2_X1 u2_u1_u5_U78 (.A2( u2_u1_X_34 ) , .ZN( u2_u1_u5_n146 ) , .A1( u2_u1_u5_n171 ) );
  NOR2_X1 u2_u1_u5_U79 (.A2( u2_u1_X_31 ) , .A1( u2_u1_X_32 ) , .ZN( u2_u1_u5_n103 ) );
  NOR3_X1 u2_u1_u5_U8 (.A2( u2_u1_u5_n147 ) , .A1( u2_u1_u5_n148 ) , .ZN( u2_u1_u5_n149 ) , .A3( u2_u1_u5_n194 ) );
  NOR2_X1 u2_u1_u5_U80 (.A2( u2_u1_X_36 ) , .ZN( u2_u1_u5_n105 ) , .A1( u2_u1_u5_n180 ) );
  NOR2_X1 u2_u1_u5_U81 (.A2( u2_u1_X_33 ) , .ZN( u2_u1_u5_n108 ) , .A1( u2_u1_u5_n170 ) );
  NOR2_X1 u2_u1_u5_U82 (.A2( u2_u1_X_33 ) , .A1( u2_u1_X_36 ) , .ZN( u2_u1_u5_n107 ) );
  NOR2_X1 u2_u1_u5_U83 (.A2( u2_u1_X_31 ) , .ZN( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n181 ) );
  NAND2_X1 u2_u1_u5_U84 (.A2( u2_u1_X_34 ) , .A1( u2_u1_X_35 ) , .ZN( u2_u1_u5_n153 ) );
  NAND2_X1 u2_u1_u5_U85 (.A1( u2_u1_X_34 ) , .ZN( u2_u1_u5_n126 ) , .A2( u2_u1_u5_n171 ) );
  AND2_X1 u2_u1_u5_U86 (.A1( u2_u1_X_31 ) , .A2( u2_u1_X_32 ) , .ZN( u2_u1_u5_n106 ) );
  AND2_X1 u2_u1_u5_U87 (.A1( u2_u1_X_31 ) , .ZN( u2_u1_u5_n109 ) , .A2( u2_u1_u5_n181 ) );
  INV_X1 u2_u1_u5_U88 (.A( u2_u1_X_33 ) , .ZN( u2_u1_u5_n180 ) );
  INV_X1 u2_u1_u5_U89 (.A( u2_u1_X_35 ) , .ZN( u2_u1_u5_n171 ) );
  NOR2_X1 u2_u1_u5_U9 (.ZN( u2_u1_u5_n135 ) , .A1( u2_u1_u5_n173 ) , .A2( u2_u1_u5_n176 ) );
  INV_X1 u2_u1_u5_U90 (.A( u2_u1_X_36 ) , .ZN( u2_u1_u5_n170 ) );
  INV_X1 u2_u1_u5_U91 (.A( u2_u1_X_32 ) , .ZN( u2_u1_u5_n181 ) );
  NAND4_X1 u2_u1_u5_U92 (.ZN( u2_out1_29 ) , .A4( u2_u1_u5_n129 ) , .A3( u2_u1_u5_n130 ) , .A2( u2_u1_u5_n168 ) , .A1( u2_u1_u5_n196 ) );
  AOI221_X1 u2_u1_u5_U93 (.A( u2_u1_u5_n128 ) , .ZN( u2_u1_u5_n129 ) , .C2( u2_u1_u5_n132 ) , .B2( u2_u1_u5_n159 ) , .B1( u2_u1_u5_n176 ) , .C1( u2_u1_u5_n184 ) );
  AOI222_X1 u2_u1_u5_U94 (.ZN( u2_u1_u5_n130 ) , .A2( u2_u1_u5_n146 ) , .B1( u2_u1_u5_n147 ) , .C2( u2_u1_u5_n175 ) , .B2( u2_u1_u5_n179 ) , .A1( u2_u1_u5_n188 ) , .C1( u2_u1_u5_n194 ) );
  NAND4_X1 u2_u1_u5_U95 (.ZN( u2_out1_19 ) , .A4( u2_u1_u5_n166 ) , .A3( u2_u1_u5_n167 ) , .A2( u2_u1_u5_n168 ) , .A1( u2_u1_u5_n169 ) );
  AOI22_X1 u2_u1_u5_U96 (.B2( u2_u1_u5_n145 ) , .A2( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n167 ) , .B1( u2_u1_u5_n182 ) , .A1( u2_u1_u5_n189 ) );
  NOR4_X1 u2_u1_u5_U97 (.A4( u2_u1_u5_n162 ) , .A3( u2_u1_u5_n163 ) , .A2( u2_u1_u5_n164 ) , .A1( u2_u1_u5_n165 ) , .ZN( u2_u1_u5_n166 ) );
  NAND4_X1 u2_u1_u5_U98 (.ZN( u2_out1_11 ) , .A4( u2_u1_u5_n143 ) , .A3( u2_u1_u5_n144 ) , .A2( u2_u1_u5_n169 ) , .A1( u2_u1_u5_n196 ) );
  AOI22_X1 u2_u1_u5_U99 (.A2( u2_u1_u5_n132 ) , .ZN( u2_u1_u5_n144 ) , .B2( u2_u1_u5_n145 ) , .B1( u2_u1_u5_n184 ) , .A1( u2_u1_u5_n194 ) );
  AOI22_X1 u2_uk_U100 (.B2( u2_uk_K_r9_19 ) , .A2( u2_uk_K_r9_25 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n142 ) , .ZN( u2_uk_n391 ) );
  OAI21_X1 u2_uk_U1011 (.ZN( u2_K14_44 ) , .B2( u2_uk_n1777 ) , .B1( u2_uk_n238 ) , .A( u2_uk_n717 ) );
  NAND2_X1 u2_uk_U1012 (.A1( u2_uk_K_r12_15 ) , .A2( u2_uk_n214 ) , .ZN( u2_uk_n717 ) );
  INV_X1 u2_uk_U1046 (.A( u2_key_r_54 ) , .ZN( u2_uk_n1185 ) );
  INV_X1 u2_uk_U1059 (.A( u2_key_r_13 ) , .ZN( u2_uk_n1150 ) );
  INV_X1 u2_uk_U1060 (.A( u2_key_r_1 ) , .ZN( u2_uk_n1143 ) );
  OAI22_X1 u2_uk_U107 (.ZN( u2_K14_41 ) , .A1( u2_uk_n147 ) , .A2( u2_uk_n1776 ) , .B2( u2_uk_n1781 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1094 (.ZN( u2_K11_8 ) , .A( u2_uk_n407 ) );
  AOI22_X1 u2_uk_U1095 (.B2( u2_uk_K_r9_12 ) , .A2( u2_uk_K_r9_18 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n230 ) , .ZN( u2_uk_n407 ) );
  INV_X1 u2_uk_U1096 (.ZN( u2_K11_12 ) , .A( u2_uk_n313 ) );
  INV_X1 u2_uk_U1102 (.ZN( u2_K2_32 ) , .A( u2_uk_n999 ) );
  AOI22_X1 u2_uk_U1103 (.B2( u2_uk_K_r0_15 ) , .A2( u2_uk_K_r0_36 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n155 ) , .ZN( u2_uk_n999 ) );
  OAI22_X1 u2_uk_U146 (.ZN( u2_K14_15 ) , .A2( u2_uk_n1773 ) , .B2( u2_uk_n1811 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n99 ) );
  INV_X1 u2_uk_U147 (.ZN( u2_K14_19 ) , .A( u2_uk_n685 ) );
  AOI22_X1 u2_uk_U148 (.B2( u2_uk_K_r12_25 ) , .A2( u2_uk_K_r12_33 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n685 ) );
  INV_X1 u2_uk_U149 (.ZN( u2_K11_19 ) , .A( u2_uk_n338 ) );
  AOI22_X1 u2_uk_U150 (.B2( u2_uk_K_r9_10 ) , .A2( u2_uk_K_r9_48 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n338 ) );
  INV_X1 u2_uk_U187 (.ZN( u2_K11_30 ) , .A( u2_uk_n369 ) );
  AOI22_X1 u2_uk_U188 (.B2( u2_uk_K_r9_1 ) , .A2( u2_uk_K_r9_9 ) , .B1( u2_uk_n110 ) , .A1( u2_uk_n213 ) , .ZN( u2_uk_n369 ) );
  OAI21_X1 u2_uk_U192 (.ZN( u2_K14_24 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1782 ) , .A( u2_uk_n686 ) );
  NAND2_X1 u2_uk_U193 (.A1( u2_uk_K_r12_41 ) , .A2( u2_uk_n17 ) , .ZN( u2_uk_n686 ) );
  OAI22_X1 u2_uk_U219 (.ZN( u2_K2_31 ) , .B2( u2_uk_n1230 ) , .A2( u2_uk_n1245 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U239 (.ZN( u2_K13_39 ) , .B1( u2_uk_n161 ) , .B2( u2_uk_n1725 ) , .A2( u2_uk_n1744 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U252 (.ZN( u2_K14_48 ) , .B2( u2_uk_n1768 ) , .A2( u2_uk_n1806 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U254 (.ZN( u2_K13_48 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1755 ) , .A( u2_uk_n677 ) );
  OAI21_X1 u2_uk_U309 (.ZN( u2_K11_26 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1665 ) , .A( u2_uk_n363 ) );
  OAI22_X1 u2_uk_U332 (.ZN( u2_K14_4 ) , .B2( u2_uk_n1786 ) , .A2( u2_uk_n1794 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U352 (.ZN( u2_K14_40 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1793 ) , .A( u2_uk_n702 ) );
  OAI21_X1 u2_uk_U364 (.ZN( u2_K2_33 ) , .A( u2_uk_n1000 ) , .B2( u2_uk_n1258 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U365 (.A1( u2_uk_K_r0_31 ) , .ZN( u2_uk_n1000 ) , .A2( u2_uk_n147 ) );
  INV_X1 u2_uk_U367 (.A( u2_key_r_8 ) , .ZN( u2_uk_n1148 ) );
  OAI22_X1 u2_uk_U371 (.ZN( u2_K11_28 ) , .B1( u2_uk_n148 ) , .B2( u2_uk_n1642 ) , .A2( u2_uk_n1674 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U383 (.ZN( u2_K14_1 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1778 ) , .A2( u2_uk_n1783 ) );
  OAI21_X1 u2_uk_U409 (.ZN( u2_K14_9 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1788 ) , .A( u2_uk_n933 ) );
  OAI22_X1 u2_uk_U431 (.ZN( u2_K11_1 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1658 ) , .A2( u2_uk_n1675 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U461 (.ZN( u2_K14_37 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1785 ) , .A2( u2_uk_n1791 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U496 (.ZN( u2_K14_2 ) , .B2( u2_uk_n1794 ) , .A2( u2_uk_n1801 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U520 (.ZN( u2_K11_2 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1643 ) , .A2( u2_uk_n1677 ) , .A1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U574 (.ZN( u2_K11_10 ) , .B2( u2_uk_n1633 ) , .A( u2_uk_n312 ) , .B1( u2_uk_n83 ) );
  NAND2_X1 u2_uk_U575 (.A1( u2_uk_K_r9_54 ) , .A2( u2_uk_n31 ) , .ZN( u2_uk_n312 ) );
  INV_X1 u2_uk_U591 (.ZN( u2_K11_22 ) , .A( u2_uk_n349 ) );
  AOI22_X1 u2_uk_U592 (.B2( u2_uk_K_r9_13 ) , .A2( u2_uk_K_r9_19 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n349 ) );
  OAI22_X1 u2_uk_U651 (.ZN( u2_K14_43 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1799 ) , .A2( u2_uk_n1802 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U665 (.ZN( u2_K14_45 ) , .B2( u2_uk_n1800 ) , .B1( u2_uk_n238 ) , .A( u2_uk_n930 ) );
  NAND2_X1 u2_uk_U666 (.A1( u2_uk_K_r12_16 ) , .A2( u2_uk_n220 ) , .ZN( u2_uk_n930 ) );
  OAI21_X1 u2_uk_U667 (.ZN( u2_K13_43 ) , .B2( u2_uk_n1762 ) , .B1( u2_uk_n187 ) , .A( u2_uk_n676 ) );
  NAND2_X1 u2_uk_U668 (.A1( u2_uk_K_r11_29 ) , .A2( u2_uk_n147 ) , .ZN( u2_uk_n676 ) );
  OAI22_X1 u2_uk_U688 (.ZN( u2_K11_25 ) , .A1( u2_uk_n163 ) , .B2( u2_uk_n1647 ) , .A2( u2_uk_n1666 ) , .B1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U71 (.ZN( u2_K11_23 ) , .B1( u2_uk_n164 ) , .B2( u2_uk_n1668 ) , .A( u2_uk_n353 ) );
  NAND2_X1 u2_uk_U72 (.A1( u2_uk_K_r9_27 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n353 ) );
  OAI22_X1 u2_uk_U756 (.ZN( u2_K11_27 ) , .B1( u2_uk_n146 ) , .B2( u2_uk_n1654 ) , .A2( u2_uk_n1660 ) , .A1( u2_uk_n93 ) );
  INV_X1 u2_uk_U824 (.ZN( u2_K11_20 ) , .A( u2_uk_n342 ) );
  AOI22_X1 u2_uk_U825 (.B2( u2_uk_K_r9_10 ) , .A2( u2_uk_K_r9_4 ) , .A1( u2_uk_n110 ) , .B1( u2_uk_n162 ) , .ZN( u2_uk_n342 ) );
  OAI22_X1 u2_uk_U837 (.ZN( u2_K11_3 ) , .B2( u2_uk_n1639 ) , .A2( u2_uk_n1657 ) , .A1( u2_uk_n207 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U846 (.ZN( u2_K14_22 ) , .A1( u2_uk_n162 ) , .B2( u2_uk_n1772 ) , .A2( u2_uk_n1810 ) , .B1( u2_uk_n83 ) );
  OAI22_X1 u2_uk_U852 (.ZN( u2_K14_23 ) , .A1( u2_uk_n163 ) , .A2( u2_uk_n1772 ) , .B2( u2_uk_n1779 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U876 (.ZN( u2_K14_7 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n146 ) , .B2( u2_uk_n1786 ) , .A2( u2_uk_n1805 ) );
  OAI22_X1 u2_uk_U89 (.ZN( u2_K13_41 ) , .A1( u2_uk_n129 ) , .B2( u2_uk_n1723 ) , .A2( u2_uk_n1738 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U917 (.ZN( u2_K14_20 ) , .B1( u2_uk_n141 ) , .B2( u2_uk_n1783 ) , .A2( u2_uk_n1789 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U920 (.ZN( u2_K11_24 ) , .B1( u2_uk_n147 ) , .B2( u2_uk_n1652 ) , .A2( u2_uk_n1657 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U924 (.ZN( u2_K14_47 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1790 ) , .A2( u2_uk_n1800 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U94 (.ZN( u2_K14_5 ) , .B2( u2_uk_n1796 ) , .B1( u2_uk_n209 ) , .A( u2_uk_n932 ) );
  OAI22_X1 u2_uk_U943 (.ZN( u2_K14_38 ) , .B1( u2_uk_n145 ) , .A2( u2_uk_n1777 ) , .B2( u2_uk_n1793 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U944 (.ZN( u2_K13_38 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1755 ) , .A2( u2_uk_n1761 ) , .A1( u2_uk_n99 ) );
  NAND2_X1 u2_uk_U95 (.A1( u2_uk_K_r12_10 ) , .A2( u2_uk_n223 ) , .ZN( u2_uk_n932 ) );
  OAI21_X1 u2_uk_U983 (.ZN( u2_K14_46 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1790 ) , .A( u2_uk_n931 ) );
  INV_X1 u2_uk_U99 (.ZN( u2_K11_5 ) , .A( u2_uk_n391 ) );
endmodule

